`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3zzvviuV0lrvGoHE6xd+hg/t1hxkyrSY0s9zyes3R6Mvxay9MmwCGqW75JWiN4/
+aZXXD3QAd8o+GYmV0alDehjb50je4592J6ieGyqAI73dBKqJYZLZfRb2gUSw8Vz
RO8+FErARiHJJ59m3ATRKatvG8pFCnSApbmLJPVNnUdRP9jAxGEg0rq9mI2YQRls
TXMLwGUy/ieLUzsM1AvZuAwZAUlwydGyPwhT+bCUFojPaGAO4ojDSyHMOi6r2wvm
MBnoFCHQdESSgPSHid2vIw==
`protect END_PROTECTED
