`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XINRSOsMP3NwF3SX0pbQSDEX8p6jdWKqfsbbF9HeJHxjxBgu+4aTU6OZwuzrqqQ2
4RAgZHqOEsjy8Ucyj1+U2MUjH/rdG/g7akMinopLkWy7YrBSNK3H8Q3ylo4gC8hk
H57p4VQjPMtywMGpxGg57oAuWcl9DgpHcblP3mOtUu25IPmGRyhGd4s4oQBC1Vp6
7amjOCymDOGUoBY9ZsQSayG5mgaM6JJvZZ2q7oPBbsgPJMLjEDo+EfIxo1P0zXUK
pSLds8/xPn4ziKzoicYDCJAWNamI6Oxur/DaW/uiKeMZrmGhu5D6yZky5I94JO7o
CgjKig1h6lEhMf7IFq0qPH35YNEgzAFe64UF92zrTUL0x/HrRO1Th1lsSYr56sBK
aadNesy6LrYYzHmpv+tY7zIR5NFDJuM1e/irKfo+R4K9Lfy44/OiVILaPG5zpzHP
EAQWExp8W2lOXXBfw5rKy2K47KEYYi+UaIJ07/d1+sxI+SyNykIH+yxEJpTHzJ+D
`protect END_PROTECTED
