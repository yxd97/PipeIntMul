`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gg6tAjmY38vfqTK7CDlfkwe7Q1Adl1EbPElvib6RKA1pkEtuzDD9USXAszV1KSCd
dKV9sfDYcLE/Awp+aRcSnRnd9EGlzi5odQzjThiO9oBi8K2KsuSWwSxnqX+NrVlT
VsLzMGsj6bx12nTk3HN4sqjbMaGKVN+dDugJB87TenF6zEoSIVVYhfT7MiKIN9V3
Dvj7wR6BaIyIqTjLlsX9WPR94iqdWSj0G5szjVTpDHG5fTmCPZ71+/FHuDNQb0B8
478WYrzH59iDCtKlv4CkkRJrNx0HOpldZ55ZQXILRF5j6Yw0yDRIK9N60oN0rjgB
ReOtiOakub9pA0tDAsDlM83T/tHrPGco5YDlxVZQphdvrPheXpm12CBZflgWDIns
`protect END_PROTECTED
