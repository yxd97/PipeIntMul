`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+CS/IYLFbHfZLHRTLeo0pEOo47wlujmTKEi3V3YE+hjKoJP0bDqTISbeVArE2m6
GeDCccy8Nk8Nr574Te2eCJ4LPxL44tkHlv8C3YUKxTm01VejvFbxtWWhuS6s+cUq
ICgKPR2IEuZYgycAHfPSYvfSHxDI6QEeqXZp6+2CzZhqLKyrRleNbdx+V+6Apekz
wacGrpPHFlNtvHvzL/uzSKNUh/RpxveHPLBJiUnRISSxQ3nsdKRGEzsJaGoji6dz
egYobbSPb+hnHQ9MXNl9adan/77lvfIt0K0eMU1W0bEqWZtUMCmE5djstppRM6xU
OtO14Z1KKc7qtRs650B/PHnvjhLupe21nV3aUQvlPO5uTkGh9L6AsQtpXbgppbP6
Mg2VV2a1ranFr0WhNcKkhnO9bByLcZiIAI2FzGViqEjNv56/sXcOlEcshvwOtUxy
iMX6wYX3gm4duaB68ATMNAIk4wOEggM+4dl9dKTHR58JtqJSoOrVUlX8B7dGrHpb
NYAF8pCz5HlLalssq0rnMkr7x72YT8AdML97e40eTRcqOU4jXST1o8wK7m5dwmQj
/B8jCEkJxaWx3A6K3Q7w5aYXs9G0x+HVBcJqkx8zSdbzxMPgxksBio0xLCbvOpgJ
Fj4QMc8qvaH9sOmGmENK/NWNLIwVbXNsfQ6WzjdgyNZckfvOFRYNE52zxYLsPFM4
y4HQCbTLQW9+t9FZNX+p40fJKz4NE/ujegxAdAs2OGla4t8CCXmzgaishZpBS4dQ
2M4pOtDHGh41+ajTYNkbIMYfwGhnUO0Ae32D2tgW3E1A357QVo5bGdxK9gTAlrjb
jpgvrI0yELIGi29WYhTNZ7lDfq4qIRfchnQIPfa3KtAz6rCxAl/dZPVND2d59BXX
`protect END_PROTECTED
