`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lrErVjo8+Kesq/0eV/qGJ2BV/hsEHTyI1lvU3o//NgvE6G6KxIbymU+0x1zqCpOU
0KWB0UI58iJXUUQR2PZPuQ5ThixAVlwSSS0shDhPWd6ynquQxL1vZisOmBiPq7FY
hzonRnrfpvrsAsqGgJV6npZTJocsdARMLcvWaN8XtJxiZ8+//yny3rgPPbBrd5lI
KrLeARG7oxCi/J8s4Dm3/QXlC9+7Wuvyofyt5NbDW3wdfZkX2gsII2QWSC+8Gi8q
u6hDXpr5SONXUfDRfOzcJ+gxL1RevK0UaIz6iH/lq9Nt0y88gJY+FVOcOA6zGW6F
wsiAHo3Re7Hz9QQI7niwzbXzs6wbNz/wzFZqlt2laEZgJXCU0SJBzvs7PKorgoGk
50WpQE9kBVVw+J1rGseRFVq7Hy7v36DFddZYTtTcPpLeGZy51oMJEIKNHu6zdYGK
Wx/UOXg/STD2XtGmeFnALrxbv/hNNxpVcgt5HCXy09t1Ms27W+dGq8Bjtee3eP3U
q5TUstKgdN8GWuW1rQiP4SnqsUaknk+AHwJ7O2izoGhFrtV269UgPxATCG3xfYoK
2emtMrfqlwA8ydnACL85YyjjZagmFao7JZn3RRIIEVFOaxGfXpTKkvoU2zcTdXQz
ig7n7QJSwtMUPqpOYdg1aRPqTOuFW/FOUAymm9FVRHIKjBgqOQOh5vI9pelsPf8i
DCu4S8pfaJkv0FTVpDvCMwI6Jitbb43lXJwepwwkEb1fzQ9uKeuciH4UtHnJuBcf
g7DUXO4pDm/UqfZ9i1J4JbI62svoLzitM2sbUeXyw+Blo+Grx8/WvAuY35uU75GX
H6yVu4WaZTocI21rn5+g69EtBJ+s7caqbwO2jFB5tMsu9b2cEY2Adr4Q5aT4MlUQ
gKEn8UZZnTJFjkOryTlfgQc2nEUGGCuPgnwdvurf53Uy5TTLfmcoV7SAbIJ7MABU
gBD48gkYJzGxuJCvRbhxGZYxd49bCiuHq78I1KZXxd+K6IINSlWHF8+NivirTjSV
p2TQUnPsDys1T+X+FnqGEYlsXMN/o65H380c1ANBQNlW+mW4o3iLtvPbxEmucr/i
WyVGcvLkE4415H+R9IhJN673Fb8qWf8lIXpDIqQxawIkhpKVgJmdwebNgfFKYnH9
t3Otwv4QOUkbAo94aDADXhqJEnf2ZSBzjSEk75t3gBkvLZDII430lw/QBmUIJYil
jvWYkhy3A7yP2A4ElI6M2kN8FSrYeVux1LouD/f1TG2PgbUgZlZQmdjJ0I+NbQCZ
H3thwV6eDrYeyWS81IahKzARmy/L3wM9eDOj4qX4iLdi0s+nht9o8CmacBtqZZOe
bxETGCnVfEQXgUqgqpVFcZuQWcdQ9VlsiV5qPtixWyjz6vsmd9m++t4yOVc9aW7e
epy3g59hO7jtssZa2CljtE0byM/S/zPTgP8sMIh+PvpEadLVahvHg49hBrzZ2bnG
Johp0rh+rgk6Iuntfj2aVnKhRngjCS9FVThuNfTQO9oZ3HC+UINrsQwfp7fIn4tK
8Xi33FqwPlWFfICh03/4I5CdhVaU5LQ7bQz/8xCHkjOm8b1oBN4m9JHOia1sDRSk
cjXZFk31ZOZMOc8MziccfyLiVzeKw6c+/JKstLl3qoV/mootSJUZq10D+EHqCaIQ
KCAw2o5oJrE7bkO4+9do5SeKEDBIjfYOszL6MJvysVwXjtFLUZmZGnMP+BpWZXgi
xquWErWCUXdepR7XoZFPn/naKikg7xHcqzRCQX/J9QDQUuTyHOhV8pr3ogKvhAnn
SNKlFfN6jNn/FhUhS/RnprtRdR8rj6lylEFwMm8Nqi6YzFvn7BZ2AVkMyXS28kSV
TnUy/iSbcKDXwaScYUAOOQlgMn4nhqK1blqhoJaEBSg6lVMtZJ11H+ddcvH+RvYh
5gg3ARRuxCSPGhhtl4i1nwNa+n7wZeBSjzbMT2NQRNolYanPeCIvhgZmawXaZPoC
olQLjrAvIap83zVahOtlStos8fqxiabMjptWQAY59YOCSnun2O4XP4WLhYBkctOB
27pyzRvkpPjjDufvRx82i/vFqyFUZBbwRVlfAdppJDtQUJ43ZNS+cyAwMKOGe0mP
DvQgH6Rwl5QeVU+D4RXHsOmXP+nO6IyXXAgWMFkhErWpHkIEjgG62G5Op8Mvj//H
RpG3Fggu5x5Ak2ms38ThRKtGe97Hc1jngV4t0SgxB1BM/0GXw2fiWh5zJYssTjNf
b7xPLNYgMWqqvYA1uT3gl2UTnjJBN+o3Q2/exaueip2XJqDSp55Zv4Fm8Z5adrFL
SUWZAFgudjBzZbhgc8/2FS+gsLTd6qSK5VcFlSgNqmWIIj6nhfvSoE2JBTPZtwar
/G/2Yw+MLYWv4uQWXDT7qBuux4YC3cKtn+/+mcRpH6zfchY8PBIsv1JyIcydqvdl
z9lUQKqTHZq8EOuC87pnKU5A8EFAubp/1i93H7SexyWpgMR39CkNYRQgVLVEBAPc
gwhQxLKqP8qaz5t50GSw6F1LvUvbleYzrUaQOvk28KAHrG9XJ9QlYugSELFQG4kg
GK2IY+936kx1I3FLY+lSpA2UNYrBEIWBjvZUwjUIKUXZGdxX9WwYoAeaw1xIh+vN
Js1SEykjl6lSlE61SFjuFLclcYrBpFwYH993V3hDuvjsVdkdmgMoackmNvT3vB3j
BSbJ4cFHKG3WLja5SaiYKEGE14tbBxYI9RwpEcjqWA3zG0b97uyK9t1A+wq7Bq7y
YcS+cGWGW0jx49/EIDIcKu9LmAIVYeY3kHAFncc+nn0TZPM7H+CThG8sFShsA5K6
Gk50z4MzQinp2r4zrNDxTJ2qlCIPbDmC2iwZEUpeGRnddWyuPty+oSzZ23ERwx09
LtZmAvRNb+xjcbDleJ/T7/9SY6zWRRD6Z8QQXY9C7KczFkS9M1f9hIBJ5CqrQ62T
KVgoBvyUZiCL8id1JcZCR8lTnpHIDZZ6pE2S/Evi0iUGUSIj3gSkVyQ9ieVXlLVe
q4+d101Rw/YlpFEhOglZn6biVw1vBoqa7osjzyyjlUGj4gjkEqf6kgUBQZ8McYpn
tLUPyuwoqPopAs92YKvGyuKEkc/LcX+HrMotbaXBxYofJLoL2+YbY00HcFCPhNYw
q/ZXzilLqx6aftEi6eFjwAJUWwT2xXoZMZRfm3jIbc7cjiBQNDPBrk/7fbWl8pKi
EZyz3TYsb5UUFklSyu7ZpXbD05TPT6q4o/FZPQz7YhU/PqJ/upHoTkmWx3U6Ypz3
gMf4Wf7y3LWEX8HrG+N3g8oZw/+8NdNBcAOxTmRJzDmnEzRhHyO3p4zPunJ8YStB
55kkb1NwotzSHsNsle3KmWJHBF/+btk8o4+gwjnvV+VQaattgLKXMdIElzE4zGZm
HRp7cMcE2/gt8KciUAJVYQv/fKQ1yf7jXmKJdzUJx31rfbaN8sxlrryGVUUBCoWh
pfSZSLXPSdZMw2aU2rb05d6bsV2oqRmMwtEb5Tot3By/Bz7gm5FtFJ61P9L3T8OA
S4Pqq3NSCkLlS8k8v5iO7Paig2kCnqwy0cIJEd2N5q+ep7FlIOylfWwrHn6WpIZx
hQnIddu5ju3QUv+ax/Augh5TTmdxaMoKmPjKxXePKKk4vP2KtIKGBCl1GqWmC1Zl
RwKZcUy3YxpFkhwMyKH+qc5CM67hVncN1bf7C5NKjRKpOm/qr5lrZ1HFZESDnE6P
pZh2Ge41D5Sz93YlEM+WaBkqYwCNyJQYmZqdYNrp0+b29vAi0J4aP+oOVLAITJc6
zWMShIe9VQYH9IZ/WGrOH3uAhb8VaTWxjVnk5kEhO1GYmI02o3iG9SmlzRHF6YBx
BXjDGrvBP6fWIW4b7mjfWU43+3uPT7V656I0GeBed71zXOIL1y0bH63JpeJ7ksxY
1JkW3Dormjg65CQ8ggn2bM0omSIKaYWV66zWHTTvuunbbfjW3LfcvAfjvfwdUCHK
/AvTIUiUb+pgWU5YsLDHTjjybq8PCiGHkrdX8u8TyQ5i90pXzwW1JN8Tmj7nsX8w
709eKvxQDXXk3aLtfWWOHiojwXuZPmiXwTd3aZzIH0VSyptmU/objejvY344VrOp
0lX6Omf78OStuyuoKsf5ajZfZ9n12FvKpkUNnEejeyohs0uiD8oTgtQxS7gwF/kz
B9TvMrrS3J1xBbo7lxU/3TvtwjlLF/8v/1d4qke0iEp7iy2Tr0DQgdWYinfUrVau
1qUMcVXsOoXkIIs2vSpXGJV1v1dSYzDQg37JViYcXWN9gvFiEaZbQYChsu8B3wt/
FG8N+Mc4XR3GXi/f5LHbgQL6W9JfMAo+n6kLlbFO9MwiB6XFSXv8BdLrnLqZdblq
0LJBRM8o8OE4ioFFGBcUi3HWU+wxOUz0i4m3EbODuWG1Ue4qOrAhosoj2X1K/CdH
R6Q8aTFtVhWwUkf0SCkE74dM6SgZ9TNW+DiuUQuqeZ6PPD9o5oA6+IZTTBLS3NTP
RQJoG/zvTPTFBhxL+yl+/RKUchmJFM08iHQMJcnTjKteCZEY0yKwBaSFP88AH56T
7jYotY0GKsp33RLrg7jzM0Dz0OFI+GuSMpCiYzSEqxb0MwtgBdJP2R40x6UXhX8c
duaHcNz1H6T72kNY2hVlt0UrtLR6DqoKwjrNQXKYK4TABf9THtIABpKklF6a+H1+
Iau8kQMULZKfQb+tqbHtFMqBQvwGC0lS/9QrdcOUDz9NzbHeYRsCujVBYlhTCWCj
Xl+ECi7PpMHlS6tcIIY04oM+0YtG2U1xtjwRI/duE3FWTrt2lSaNtxCum22vjmAc
ktAyTFOVQZ+YVAaaLlZmIGrE/y+phdyhGzINNfqjymJJVRN0O+6ORXnFvsyzXEu2
+fQTDIGUmHEWsR1WWkIFVEkBimw8bTycuVJ+6z9lHNK1MmIrfXsP0flCPZec0eum
pLwTdRr9J1QgcOzKW8WgtlPPvkmSPzKk0qbjioTKgzWksiImzC4B2Ru7Lu3Qk6Dq
U1/CyzSaIrgQRVj06PybplAnRmtchYrAt7UDCEkiNdU54/rTxfDrRk0R9w4i6vC+
JTe1XRDtA2erN7Wl+IwYDzcdEZpVnl2G9fW/YvyuFVXddGAGPX4VRGy9eVIDvyuC
qhzcNYP4mVO1tG4siFu6VXI8hnRbg+jmUgO19w1fWuVryMD4+3CHsiqYBJdFeZET
1VWtOdBjEg8bVFuu9Ktc9Q==
`protect END_PROTECTED
