`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLx76lEagA5WH8ygFF2+H6kCtVyoSBd5TuMojHT2aY0UCNDDEKnPI06s9CsvS9qP
Bywh+BmWPw22zRtX6BUbIN0fcoXVvvcL4CnCs7J6ON6mTrgwiHnps9jS3GtY3F4G
VVSl9KrKMZhLDP0If5sRfoNweROzRmfSfsLPaDdd3N5EhsV0c6HuJEHaVyO31RHy
0lQR2ZuLvL+2NUhyGQXjDyg48I6LzJm11pvH++LPGZVZ1Yg3xBp+Uqjm7sjx9ZNk
egu4HBqAgrEZJ7qR2EsfAwCwRDh7qT3sWLmAcpJBI6X0DMviyC1+HBgNmx5YEmHy
7k9S+A6bMG4Ab8A857OAmq9ylGMZD9TPlTpAHNCCGW/PYipUyOrt17KiKit4ARNS
XSPQPI6q3BE7pA0Pqa9WGXEIoxNwszzvQh7vdAyJJ9e9XQ6Q6yFQeXcGCzA6iT2/
5fhjhtUsX6NAkZY7cLfSmX1JMC7y2aloG2l8EPt0TZc=
`protect END_PROTECTED
