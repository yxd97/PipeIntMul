`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nGrhPi8p26n/TmSFqQKBYv5dijHJmf2K3Z7a4fBJchC1mrxw+3uUnkT2DDgVYO8U
xN191rjcUPm6BH3LNSdCzyLr5PGzWmiQwR+57Skj4UpqCLZogUm5IFgcX9SmP7RD
Th/NqQzSlVC0DMkeSgJ5PplpxImwaBvvnn5mXcaqMm7S4ZhHSscsaWD5lNmoG9I+
eG0LaSmOAXxpnsFAXqxFsZW7hMbrrhnt+4sZ532E6I2DECBoiQk+iJ5dsENykn9j
PKjAL4GrwoQB6KUwY1xAamThRZSMfZiZMwJMpfbUsZklpcT8P2U8a8PsTi14J3S3
YFGOZwcqYWPszXm75SUUJElP2Aei6Nv+W6+X6g3GuluuE42Vyd7ufJuzkHxUB+rE
lvHM9IJ2Zjw73bbx38F7VAwnWZTfDBgc4RI7W/kv6bIRgjHz6SdOR4JBP8QmlaBZ
aSa/nxcDdYY93R10d2ltH1j6lUD8aUcSnINLu4UI1WiwSLytD26OLYjs1dw++Dzr
UR1+tuS82QCi2AtD9JKR0XQMjf10J7k3zP+XaSjANnKQZA3PM0QtIyulPMC9ZeYh
yVKskPVQfTDb5dtxNclIzQ==
`protect END_PROTECTED
