`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WUqODBs4bSFHT2AjjeuXWmHaJoJMGPLWuKZur35Y3Vkud+EMyKgUkH2iCJ3oJPWk
5fXkq0+AFS5yHX/9+DEkvppccX0nIPMQgPHIWSPPwA0W4L3klnjAi53qKRg87yEN
SWMC9aFJALmFZUFWIrLORXl42u36M4VTWwmirRNvo9UrLARYaeUCSykhswawed2a
nGz+fZzzmSQnJAEZVo4ClZygPkXREPDm9CNLA+yTnYNcYmFPhEQpIR4c00GJ2lRQ
Zfbr4IByQ4JIHw/EOacIkAdUY8qYGlFOdStyGQs3xRM=
`protect END_PROTECTED
