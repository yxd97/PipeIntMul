`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ME7QPJaUR3rBXiPQnGtiPo2dbzJHXdADTEXNGEfonZFMDbHhe340dbPoeMhy1lEc
FauF6fDuIcRk3/zU+WpDWrSjc4iJajMqux8uTafBCp+aA+X2j3PJdf7CLF9Htzpu
exbLwFhy24u05tBXlUvSskwjpAyMCLyYrihtyD6Yqk0Zre4vKFwS2sdxZ4Df4GRF
y+zvTN4Jc5AOx1+C3hPNDA25Ve5qSt9BShad7FeY54OEXReXldzNb9aWB7yTY3zU
qXZLjqLGnA9cpPqCHfSk6OAwLmzq1N32HA2ThvLsKiiOdmU4SJsJzc4BHkcrjnG5
JDFGl70IRb719AYmhSpTwJDvZ3VsFtMPtja880OXO2ZZfLS23i8F/UcPqzy1ysJu
aAxgjaaZo/tyEnS7nO1ETzkeg6KfIde2nph2mcy/2W7KiotGpwerQ0CWJ9mWxq3X
AaqhcSb/8R+fpKJY/ghCHnz3Hb5cQRDuxKwegHnMwajnK3ZboVrW2Zlfu13O0ors
pvquvgbfJrO9VZa87TEUnGJ9Lm7QKeNyo8C/b+bW7t/8i8KwZOSlW2RJQf1rB98i
gCWsfAIuKelWcveJhuKp63sa/1Jlj8dQffEkgMmpxmfUIeuSRo5wcMMpnQMGDSZD
XKYG/WwnHDx/+A3mN5ZQvLLgRmXkDYje/ubvc5xFeks8OYuMCkgAqVXtk/wh6F2U
N1pnrLPmVRB650YYcP9BF342vXU1Kij9nPEB2ZY1VS0WjbtrJudSR7dRpmhsY1mg
mIa1xfaIczKjfcFxiXL18RgGY0rT+lq5+M0/FRG0Ah9GHe1TicZ+mhgirmCgv6El
bgXpEjyyyalC+0AViWZmhBLblr/9E7DaAQt3Hu6dXdfxR/qJJnj+8J4ITytg1WkO
2vDIaoSJzoqcsbQ2lYCmPrM3//NiMfUnZaCfTg3gEAZemcZGRXXAfVWDpGnYOOSW
13UlDO3iFGxvIftxQ+YcA3JdBAbKCWpZCBEE0ZnpFEa9OsxFr5jLzUO9RppBv++8
XI0vE+tdiRmgQTnuNBFvwC9LSAG54YdnV4CtsoO39V+HPDW1pusNo1xtskpPMdYO
38nvAO43q8tO6m4Y/7x40CTzl5ZNkXMgEbaZakDPa0G6Yjf7AKVuE0ZecqFGxrZv
8YAMYvmP5wDL4cbIL6v7iy5QtDTa5sUT3+jmKQO6Fu1TFoNe2zkHM4RXHJ8LS9Tb
yR9TSCy3BKRekb6V33cUGm5G5jmF/6Z6O/EdGMZFJAigeucwBYL+3xicZINESWSs
gLj/teBjIL2GqnthN5I3dc1dirYHf5KxSlUMkNh8sFFnwIEujOhBpz6gi3/D6BwD
CRQidNrApbmf3OqF1gZUbXz6pnznjU5/isv8YN/Il8OFERzoaS/fLGlDmFMHPxFB
vJqHLWhSHVG0WzCQiFe9Bk9ivzlYehdmGvBMvICx44rwFcTTOBA/FwAkEB74MMVu
iTBG/epHyEqI7axOz7Q6+noiOAvXkzeHgQ0yzatmUorNgLLFdtidWW4C0dNLH1DI
g+S3AXCIb9RWOZo3jxQD1wWyNVPAOQ4ryE3L6lIqOyLXob/Yd3MYlRInhw4N6/8Z
SedAltvipznnm/bBw3DU3ePiNHTm4KXjBCg2oa5jrScJZBlpPsHaFlQT1IZgfVBc
uVJMqE2YGcsIZTE8nsu+haFFpYKvvm7MmZpDsXh3yUEtfjY0jLzk63lA9GsFo6da
aa9egxDYwJyaW2bBne7p9en2wweCvB5NF1n19VLRe0Rzp0rSOst2EyCO0pLzRWie
LvumwkX4ngae9dsOLLbeWc+oM9ruYsjvUM9cxnJN0QlAXfLfwUy0u5/7mtW1BRjc
Y4aGdle+ozlkaBi4Cr4qZJoKyHBeuNb0c4gRKyJHHbKcG0n/u+oBESu940LE3Y3n
6v6R6upPkJTKzydzSXFuLIgR4rIGIGXysgXfig1Ji8noendrcixgR4rElCpXRCK1
OeV3jOJbFqmFp6zjDw3tbAC//1CHgwHyu14jrqq2353KspPCkRQd/himaeKeLtrs
BgIZi7VvnkIJXophGZRRhv/2+fA3PfOrjutQuJoiJ8LMMuoVYtYqv+T7/XHbZuER
bWf42fAzSOkvHswmGsJdIggWJ9tP/RHDEaEPePENfvJSHCuy1CH7YbASCwvY5vxj
4Pb3oT5JqPtTgnPRLHtI9brzG3WV4kmjxfC1mJW75i6Y/ovCB6h8A7epxtq8Exx/
F4t/E4ubgVjqXxEiZa42+tXy+qnlyXJ5nATa5JWVjnUIe/7m1ypYBxbD26AXvVmR
v0tEFxrWtTz01U5fw06FJW46I290CYV5V8Qa1QssSd3kn5EYWNIkiU5FoVwtd8WP
SAhYDg8DrDWdKC52QIzZzPtZhBCpPjzUOfNxldE/sHx/0v/i8w7k7wX3RS+H7oy0
IGDgCJ4uEU1q/N2DOhfCPQpro23dZ0pRaULBMwzPP8nS6nUVLuu9u+40vMgRjBZD
jbSqmL4EvmY7S1jDFiY2OegUBfEXhZ4ltk/u/aTWnvBAvotTGbKat5KIP6Ue7rw3
adeI7SlusRdI+aeao1lRg6ZKbrAiS8VNxuB8LVVpfABUG5W+R7FeD17R7rAgSu4x
7Xipvx+UvUj2b3jSGjTduQLuMcriiowtwkT6iEDxriRMOGRSZBADaHCcRvHk8g3Q
2sT99MrBY7+yDWClVCDAl0B8cfDI3fcJJBEz9KIE3sq0OeYoL4urN0lY9i8UyF6k
60ojz6S1Q5k2Ssaeiw5pKwMtVoOXSxgB05B6GXkJOqjhJm3y/IWNGK0CGu4gqoJ0
O3Xe8LD9PJRV2UKdEqMse0ImzK5M4EN9iRWfTirJbj/gQjlxrWwJo1AOtGSMRtDi
FZ45zZAnGkAtsYl0m8p2c4z64y8ACurWCjcdg8pvV2FAkza91JIQTOY5+x6AGqja
hNBGCvXNc/K+45ksxeeAglRF6j2WAvieJCwjsIq3mPyS8ZrydXg9oA5OSLJedzrG
9B46sJ5Slgh/Y7c6uhE0e52TNPEnm4ANq0qkDCaPd6GBNCO3s5UvVsgkVlKKE23W
5ZNSgOB2LBLy3UoIcXcMpSEp9QZJdSoXg9ia9XIMj19nHsIxIEU5cMXKjuXS0sVt
aPrAiiYomRzi0xZ551INxTiHnsXIp7RfFEJeLIi0cwizZJcJq9hiyRJBzBlnINru
IItGUN/A3UW2WcYvGA7zkJKiW+vhuNL6nS8e64eVFdAF5qib/zQbzfV/Gb9WtWjP
ncFioJ/GxcjF2rtVMPvt2HJhn+q93xOEl4A2aSvsm6BC4Pfed7UBvimjVAI9hb1s
SSZ1aXwZ2gIR3JtR7nPSgOP1GJD5mIR/fxjoxzjxku4ZJP/DEtLkrAwebUNG0C1H
aEc7OzEVw+NpBsUsc7/QhAhoqUefMd76Vywkqs/5RpG5NL0NldlXFnWcpei1cQmb
6cDP4HhlhxwI2Lli6mc5DXTtMuQzytTRwdfFHVdxpbu64zpiOnW6raYh3eMmy5do
MNpIXjve2d7H6K0JZJl6d66pky/Yl9VBydwEj0jli0h8bJY5J85UVJWZ8z1NBmJ+
hqCGnbbMk6fNKYuLy6vVRK3FPJrt+r6dEsAdLM+64bJbYOj/WSrjMWZ7oRjoRtg+
3dffLOlyb4z6XdyGxw8AGQAaWp2JA8qwfdPQR3p1nZ6pV7qiGpNiyRWbqAzExj4J
hoK9tmWU3ZycZV+UNxroqVo6UMr0QElBiXBXllElnIC0EqtULtFonG61M4wjA5nO
Aer4lljUg1y803jW16Wa2CRipHeqZ343WfALFOni/j7rn+QAspFgq9hBPqhJ3v1F
ehqKS0Mk99bDUdiqaLAcvF2hSAJFf91JWONzqAEfTXrU1uyjL+cupPFk9VgS1op4
u5RRSyzAO2einTNtbK8rma05azYGIXM4rg6Ti9SK/oS1JmyK2+2NAGmTxmXzu50x
Ow0AwSzLK7TnsnwD1XTynzgyZbf7JFqnhcIAAHSaewsjKNNV+RRqaxjmb9uxLFDm
7q2ClIczYM90vOmaa8LXp1r5Dcx3JKlfyMrqHASCT9ryExw4PU6BJqq/knP6vt/9
JqKPcrCfV54Wk8jDOOBb4ZdfXBkr8WxFu9nwt4klvPrCAhwfzdUUnYyu3I6a6Qzy
vDPWc/zlpFjD6tRHO3ULasFI2gRpGyHUyfxqdnsqjQRprWPygzzusIDsGyHWt84b
ZPeenGI/WTHqseXbqeF4fUwq8kN8rW4zN9UJAspmFJpf0aUwcSluKJWD8n2flpmn
MuAaunATf0QnYJQ0fOiAjq5iJ0LaHb8q7AQYdG4GoUA41jrL4BC8PQ3hZnCvxvHc
X3Z1PcqUAc7/guA6SL5BmwXrvvZm6oyIvqh4jsRILpiph79n4gVNvnww730i4dD7
a7gmBjG0S4H6DX56u0zlKADRErsv9XiQu1UsiEG5s+wnhrIFmPG+NyPrf8mAuAjo
LsfD+MV5AFoA6Uuvcn3K8OInIcvUC9V4Uu7LkyFUvXm4k+MpxxHRyLcsIdw1++1z
5aHP9CIa1ZwiLEX/nxdHMRb1YkMcwiNfg9FNzgt9S2RxS3WLSHy5NlxjGTY4fqos
/Sr2y+rQyAgtynLSwyTTP4ZZZu7UfFRznEjJaIAQkqyQe3C/MYAAZ4IwYHZ3Eh25
B/eTAokCZisJt1ti9CJrYrYRd2yl2fIVU0N6/nJs1nF1PJrOs0FLLGcvZCHkQIAo
t01TsztvFDnMDMeXoURXPz6kTQQvqx/liGW8ybziO7jTVFBkeeNqE7Acz5nXB6uk
Dkgmy1KgFP/mmw/Y5T3i8Jyzn+2zsOw+gte7DR5btU+8MUP0Oof3N7NVl6Xiitic
bqdyuqR6HwNgu0WX+rVC+eIJKNLpDVUXkkyuGCWvj13R8Yn6TnNOBnut/0dtPCXc
zv0O6CtD7HgsgN3IFO98tKmYAWh7nGFCLMTLCldVPDJ5mLTEz+uWLuCVc3ml0Gdi
m848ueuV7eW4lZ1gGYQDoPKqHHXewUm7lGf6JNdOZeY/odEaB0wMOjJmheeUIdKh
Jw274eb6U3mxQ2EpCDllC1h5Kkf2PgbY5qml/jYBhzXIHSbzyLviQk156VbE3oHx
jq1+FnGsMBmHrsLBricaxeGuN2MYxVkcaMazT3N2/lXnuoqk4ekPklFYxPYWGTcQ
Ua41VBf3HZ4kxFkgTPLEUV13Rb45lEAJ2UzRjY82V8yLdJvSCpK714giqYwGvm/Q
tasY7RKkt7H2jZz7hzOKxHXCccdbXJmuyRZ8Fc8pNEJAq6j+6yMQS9DSdc/2oKLK
6EYUCG6xCVGZWwohCTyteQQDNDQTjj0jPygD6kZPzDFPomVgnHy6FBbErmUWh4c0
XKKdIRFcg/sAtUXUse3ta+xH3aqWQd3Pdu8HnIHcgtKakIAUzUOteHg915LKlNOe
CsHjzGBZYrEtse6jN6YzJx9wf05R0QsKD8b9TXHOcJ8pAbQ5u9bq3jziNuK2OnTY
kxHKSAoXLKuKCi3+Sqovq7p9UgypU8Afz01A5V1NSIDJY6Nss2+70BL+f4QGAagU
sG5swRCcwu1v7d4DB7TfQJLTw/AYmFVMtaf+YvLX1kSSZtsID/LKnzTew5OIMZOV
mNNg8lN2bax5qdFk4T52xCK2OPS+Mp6rk2mKDyDeztGoYx5kImYWUoUszlH92Ijv
dfK4bIEsMBNa9WHfA/M7G4K6qRSAiH28ITdY7JDe/SCys7Q4x+Dk4aYKREnuQWEv
BbxfaqE1dGLogW56X69oLdCBZoFv6KnJEor6ZgR/1CM05o8F4kOlyWX0WZldKkef
+purk5ui29/aKYslK9XTdPx3tAHkukidKrvNKJnMvdBynVIahUSYarqsIjOz8N2i
pjSjxVM9aF0NY+ye2mLPyax2kUalZCZHT7YWYbKybrW9MJv5YbW9KYsRwLcvgXlk
bcKhbqyxU6IQ/w5SCFoQBD0ar9S0ZsVocv6wAE2bxxDT8C04e86CVvSPDBzlE9HD
fmgG04PGlD9Ioa6fisZwFEoOjyvIduivVgWwUJ/n6aYaeRT4jzClEvM9yfGju/6z
Xzjb3PmY6AS9TuxIeNn9ZiY2YzQ8JoPCgSsgy+ppfDnQmZsoZU8EjtDONZqpMxks
C4AybsXr2Ip31HZ5yVuYfcY4R/RgvbAHQ4W44KXlX9qItiflgKksIq7FlBzxWIHC
KshcHCjM7EI0M5WjeFAmIdDKcq9GD0iwp7BPqkbpvKqUg1O/9/+Q3eVuRfDo0/3P
YwrWWJnsB0FpbS/wiM6NkDyFLmPRFAac9gMp6moM4chEgaihBw9vg6kaq+2WvQJZ
JF4hPxhoahmgezMoVt0WAI26OACRPfyLi3bRYs+SdQ7uozvHHA7Ov6avG0xb2kcZ
86/hx1+BYD6hkr1R3o5zKWxTrzfIPcIU+l1as5sxDXCRRe9arJXwzuC+LABaq6Kt
JQ4cBP+XjIK9iZvt77pp5lzfCe8GT9Ey51VkpzeMPGfW292B2vM9BZphKRNWiUI3
Ol88sbxG3GDx6Bbjw5urCpwO+P+ZK3ll+YNgjP0WjZJY15jDOiiXIshS8/QzKlV7
R3UHa8veuL3F70pZN/aMobUrCcCvWscsdJQVx5obnQNvWzfbCC9wmb+sGslliOQS
O5C1zqXRHiO90qLmniwAPWt5t795b7m/0rTQ82Ul4dG8Q19MUCKH4TZ0tLUzO4rw
eMNoXXSXY6QgL3v/I4WfaLoZtO74CUZrAPwg0ErYcIfGQ0TUVdyXKM4e2F/EtTh5
lA1IRPGAHCp/A0rwKB+7f0m4FGmKH7gMA3tNf+lBVDk4mf0e2sw89jzFrmorhTS6
HjloVgnI8RnOpNsPPKcP8NyvffR5wqoXM3DZZUbyTvbeTuXDSZcIRbpvXHYLVjxr
cjE+uygsA8zscuKT4ocsofstEi9H4wyPwUszHGlaQnHSO+XkzHAXX4j4psD/IQ0a
SR+8Z3RMePJEbUDnmCLaYKt9QWjZWqHBCEaibjo8sXeCDZUfgJ3ncfOHSNILP0JH
ZSMUbwrei5whdNoEtxuAnp01YxLOLN6M2Sf5Zzjf9KppWbq6o5Xs0AsU4Tdq/8Ip
QYng+1QLGE1gCWHtVxinOp4hCsSDiJnp+sdBjjx8PuAeJiogDRatQrV2Yq6m62Q+
4EwGtkFv3j7+RuoQYx2NSmC2+EpgXj9M4a5ZuWnA4uf/QXhLZdO+Vu3/x39FLwd+
Lm6xQayjrX8ELTQxRnTeoVgrzf16kenvOZsmCb+3WfnP0pPwsHAIknJU9uAIrS8E
Fv8/bMd8TJE0X1Ji1h1kleoikNb/YED1u9os3Ov4eJ/Nnmuq/MAigtCdJzsecsq6
VaG65fL0WEJlGboJD0v4vzCBouz6CkbpCMYS4ONjW6Q0i/yfv3sPF5CWD22Zcw2R
T4KZh/hNeXcFnFQb1MtknzLKZzfbvfGywyQJU6R76BvlYTR1sAq4xbWpDFjlMnlB
jj2G3XUQtWHwK+ybwCN5jKvX3XHYt7VYmM7zBTw9vK7Vcih7/kc4xYBVMVYet27Q
1yHeRHoeqHUdLsIvvjlhXd+YVaXyXEejf1apGCRGtG2tOAS2OJuLkKEgfN+JPTW4
Xe/Fj3iEfepW27Dskw4e3c2w6i54UKTA6pTWlsUWSsLK+M2MnS+IcmzX4XhR2/JO
ypwh/oHBVXczFAwW6k6pl4RxCF42DWQ8LA6cOBPqsCBKLiDePNuaNelX06Z5L60d
W3TCca9ZRSsF6gzvqE3Xxy0Ll4pmJNkX2Qb1vZyRLekOyohJUJfIJas4xS6Ni6WP
mWBO21Lfg+40U5Mf++LKetuyZfflu0VLwxwFFHhq/5+olyw+a5PT0y/RIkv0+VPa
BIXh7XWqgAU1w4BGSLUHFbHZhhQorJNV/kQRFjl6T4/SsPc3FZDeItyI9O9ii9ZP
p+aY41J+WfqiEzDvQXj2gZrRynh/a4AsBasg48W8aPRrFbVYBiZoxhUY/TgRVd5X
alCg2sOWw294erjAlu87kFSnwV2OP4fSN2D6HaVPJQLcnl6xRThTfnInrni5aVC8
KMwLJFoLinni3kMrqD7h+97EKHssc/KD1UxScH2cLE0ruYbVCJ9nNbGGOyXFg4OL
aylzdzGh8OZLEzefH/iNQAX8aXUFqoMEF3TGJPg6rQg=
`protect END_PROTECTED
