`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4MT/iaO0u/oJECEomJ5HnuPHF+cxcZ44ljjRWjo7jIbSxPSoJpCi/XhrHBObHEVT
yVwSLDcR460aoK8A5HBjYB3dne1PN/G6JVsMmDqLSs5YPmdmfVrBMoj9lmqpxNsO
RIToP7cyzGWyf/J750VseqhnKym1Yk17EPzfAf2Ew2F7TrjTpPNM9OK+4+XQHh/G
LehqeQ7hhuQzfLPuGq3U2c3fI+AgYgnXJE6vBvqNAKDBCLT6ZN3xITExtoQ6z7cs
66p0Nj4Zh4FxlBnzbIVZxg9Imdxr2IErfDT1zVqFwHNAOnFdPQLWbt9wjo6Ypbdm
a2TOnu6VD8OE57mgpBLPN1rmjsK/k9H3yB0+7FpC6tnn0UaddL5K8RLuyGgYBTWB
QpirkI7++qLDJVorq02c5ZZRan16G4y88pxx26+rwNBDwG7DFVKff/rmOtxsB/Eh
tMnuMZTX35/tV5/YVjTDk8YPe2lm2ygRjyoQGgQ8b47KKLB+arQSaJFqaxTml584
PvVhBHjfSmCAzamVXA8fS/j8hUzzGusLZhSMJ7OvNR/oF1cYhqGVBwj3jsZC+S2z
hGmce3cxvATjudhtjLRkGwcZae9sAjjORbaKAZHOuNSm722tOcq8hLCK6K0PrKOQ
sF5Jhr8sQJ2AhmkZj3snUf0tzNwAExVKEdO0pYuMmUfi9F0zcdFGctZOjXIu5Wyz
bXKH+5VO5qSQQjFsr0oxTIVZY7ZTMATV3RFbAqXWuyl36KkzL18dyn88vZ6dXvcj
pNFx6blykLs4A1qtqKTf9N6ME2ydLvruGPAwHSdwwfnCo5uSueFRz2lhy/pLqCYC
zz5taoQLU4ezNmgS3GoRJoctX3HoEhKxij8g1lDYSP/vlMs9N1aFkALra9VZBcfZ
+Ovx3fxC38kev86QD7V65lITU2aC7PzLL5CMH6a4brFRoK/I6VmxiMV4fBTL58bc
PjUAawwyywC+MzwmgJ6U20Chod8wnW7V8jvNoxJqcr84mDvsBq24ZEmEBii5e/gz
B0Qdi3Rm7jWLQlmjeLaQ8IRW8BcpMioIJfBD8W+DuXVoUT54Oi2MeUPBJYyU+Rpa
mapQhlLlQjIKqV7x4Zc8WV1WDWrQn1voElAv1/ui6GG8nztzf9HXe0rB2B9X9Adg
LftLdGNcqGKK2o5nG558jBYUyylRhLsCS5dl3daEX5aH0c21a2z3JGe9+vv6/Azm
mXvOyX12tUxGwefM4qToonbnpDouQtKesehKx/zPO0IDFTMcNbdE7PniieZAPpIo
EtVw9hthQh/CLwQB2SHn6WcRAkYKIhmKXjbCURV5p21qkUcH5GW8n23BHILZAHct
ZzV/zI+XtdiIUTJ1yvZZo9ivwD3voHQYv32nsIDx78rPaz6ZHetzYJQ0yMv8OEWb
lxB+bLo+W5qCKfeXWIaAaRAVtB8B5/oyaPZ7TQvYM5NjURLqPOQh2KacP0+RDpdf
dtk5alrAUARsu3WlHx6gyxle9rYOg7EjqNwd3oUss0ZRBX9mSAgJuG3vIotjagLz
PDZZoets93mBIMwSeTNp6O6vqczdQkk1mqXsTvG/qKeqyj6nEIJYc3ZrIcwLww20
CRpGLusx0Pv6UTmyfuQ+Bg0wYaIJkv+1VV4JZWhxJjA9fVkKWZb6Xeze9YPxUAwf
n9K+4ZSPAM5G+0Ecul7ERS2ANbos7RxBoai3/yxd802Y8XxvLsjgy5TYKNimjUnb
ApYJJqXPFHJKynQKqtcLJBPz/9j5kJtjjGYoRhcv7TJpWha6zj3xDnHeW72EnmRm
fw1W0iJhTBibZaNplkaW5upkzJ5ZUl68Dno0GndL2gmvIZKoVx1sNi0AVYRF1L3I
dQDAAEz5n2o+9nyPvzMq6N6VMqY3kGvVDyChPW7APJ7kp1MK4z2LX63m3d45cBvr
qrnZaN9DJ6dXW5CNDwdoEmzEfDtP8HobHs5gULYpUVz2ve9X97DjH1Zy1efMA7F5
XAXw0TJqKP3srv1x3YA4UMQjBpJKk/VvpzVg2ijAVY6wBW12mPWsphB/ZJnTuP9F
u/kNIlc4wY8t0fvDZ1/LMF7tAez7U7lQ48qGs4VCFOpFNDTwe8KjIdMA/bWJQn+f
EGkVjGknYklFwQBJahsvfunga404m6h8fvmV7hSoAr4+UuaOl9bJ19RlsWbVm5SJ
rj7G480gw3kJs6qJ7YM0creaQk27EO6HSbZnC0D56IpYxJjUaoskwD4tpsTfJprU
3C6njemMDEU0ZTlXhmarTj3vQdefJ2Dx3DSAoi1ZEc6KKbjdohRxKh1JGoLk7R3g
GYMRur+dBABV84tteeSqfeWwMvcAlbVw/naRmjizM8B6uzHihxwJRjXVqNHJHcEn
QgJ07leuOlXCqUXUBe8HlmxVoEiNPLD8EJVxFIJ9RXDGqdMBUr3GhBxHN2YN0boA
V9tCNuTXTfEhhVO+0qkuhiBJhJwTfYvelKmHOAuVpv4e0aM0alXLgMa5vPVNaJYK
lHIy8xo9iP5d+7Iad0IrdV57oZJxua0gJaiSH7KsuTjCNbx6PQm016XNSdKGgNA3
XRfp7w7MESPzzGwki0txJNC87wnMbbS5tF3ptqe+mhcMcMcrFUktiv1HFu/OPw1h
ho48UkzFm+G5Mop7EeMC+6N8CViV15khhfFhQh8Ytq4I7jta76JmVOfgF7Tk04CT
Zuor4iNT02qyhnDO+dux7Ru5KbjHDnTZBoOkPTVG0sgDFEregpfi5diDsv19e1Jq
XynU05ZSD5YyMEKO0noStg==
`protect END_PROTECTED
