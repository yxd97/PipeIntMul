`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yWQFKZmFJHxoNkJLC9k+MDYqrAcB1aIDV8d9JuX5dvwk0B351ZOuUFb0XTVlECd
YU0xzSa0kA/fskn91D3VmsrbW/KYc2Q9Zyp03gh5QtagwlsMPIOMC2tMiAL4pNWM
upanixpP9AuL2tkIunScRcROwLsDyU4OAqp4nbsVAlrh1HTKZMt3wD0vc+WWnpPM
J2PrmkhOSrcFpHj21FrNzutDR3KlSAihLyehG/Yg+EvsVLL/l3CtZzSuy43Hd/2V
5QRx3Dnd60l0W9/lunrJRfGMF2aNY2jST6MBCc3ZmD/aUQuw93j9FK6Yza6GNQMV
2ijk6LxM9kHoOvR5CRR7Ww==
`protect END_PROTECTED
