`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hojKTbOUY3vNL9IIqYoIpb0bMSi8fVEioOLpsgNABClGDe+NIwGJ8BVZRlJ8AEn2
Qhewa3y70jlcerkIq+HFxAD3Ey98nosph1qTRKhd95LhOHAwYxQpck6ZMCjJyN99
G320lCCbOEKpKpC1oe83t9ZlkthmjZvZj6hktCAXG4evc/GBIh3EiY5k45Xmx04g
qJ8OKKgsAn0NvPSAmpDmtuHzmce14mH8cEWDlZUrCYXm8dz0vlmU5XMrqfwKRGOd
8b4HizeeNuuNmVFVNYMNzViPrD7pDkI0tynUm32EGpY=
`protect END_PROTECTED
