`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
drZRGucekkswjVTLmb/b97kRQi5aMHEFD8iiLfzTZJYt8VgHfTTq+lOjz7jZq9BZ
KWbwMvJi3YhSy87rVAOkRa6IIYn0uwRUYk4idsj8g3cTuIi8/cavlaBoGwSvSZbX
ZLSrt7UHeHZSmoJlSB4udFDa9DuV9K2qqt6trrdbHMF0abfCt4GvN5MMDElgYfSS
8GHAylS2+KlLdn+JCMx7Gof4266PtFPuJbAMq1twc+p525VRVaV8xK1xFqfkq5qK
tLUsW9wBVZiUG+y8ZOAXaJJawO/Qeeq6jwF6e4i2rxLYxaNEztGieJR+mvCczIsS
rI9XA1sCj/C0hoLbE6hQ74Cv//cgHMXxCdpgrQB0PhcxanRCaQtjWOhlArEwRGHF
VLZ4IrrciKN16zNU9fW4RPfKf75xshvGSybsXH2geW/w/MCnDdtZ0d6etDnN/KJu
6LkNqniiOWG1Kjx5OA+0Q3pV3wXjPrWsSWOmyg13Aob96O/9JXvUs2AqCM6e/ISf
m6L7TS6p5QSzxTwxe1/jSrIKChfoEuEXCbsatuvUdGAsjBRKci37RlVkLm9cpPxK
ymbQFJChKdWzNzZa9Swa8R5dDkKZxOB0mkYvPKpF9IUQj8I6Ccq5tcs4YvTdHHT4
McIQ+tUZ2A8oZfFbaeswGiCQsttk2K6YKZAIJZbPXes7neJx/F0k6CLxcMyeBDDh
v0TLD274b2x5/rrDXfn/49hZq3JN6bZwJW53T6VRg89R8ibxuRiiw3dHxbZmdZ19
OG0ykhNAVgMNZ/MZYGJ0cLfqFSw15SzO/87ypo7c5d0ENbAVk6Mr+Q19XT4TdgaY
Ts0TP5PEAm1+pZ4l0pfywkitbyYWCNB32lecBdYjUlzx9Vpj0y0Q0e0Tg3DnLwDV
/3hNSAoNYm6SkxsTFr3abzLRiaiakH6TTmMtBH8b1kE8ReDP5HUcqpHwL/CfP0uv
3HG0BzVdDTmz+pOyO+WmhMItH74js+JEY9/jI5X50hhEO0fojA6nK0iKpNwPKFtq
KxHsL3W+eeRvKFNvNIyunGg+0Gu2G9PKbxufcrfgC/pSKRkPc6jmxHT3PEfX8zqe
xGnpMaBjV2gP6KarQDp2n3i5Yh4QQ///iEmOLYoh2Kjg+p7JrRd5wThy8ltmiB6N
tROL0Qh6jz3bkgt/dkjnRmCp9hVBe/o5mZhZoq5d9tXvBIHX9Oe0SfNNKhuXYNuz
pmLyY62PfPljXNK2ymVtvy6uF825kM9ThQTMBIoEdM3MJRLXQplUg7pHsvDZ2RLD
5JUmR2fPEBYuAJXs86Z1Y3c8zI8jGWDtdY/kgYRCjsNpqmj+MWl5U2T/p5I7RAMf
GgJyA53paYuUybnbxDfd7zRlvIDwF8Awg6zQFjr3DareCAIabvMecnp0oDEDHb/1
hcNkhvcFJ9vEJlEAtZHd2WUbI8kE4Dv0d1PQ/mi6daUWj2XgSMUPnuLk9X5/15rs
5i8cpOILGV83jMcs3bl0XQvKlq0LCwXEhR6Xy1Xcpl45NQ8fGcxgub9GodPxHrq7
Y4ebFFTQD2yxPy6qQrXHbFs9jZMuPH+noindU2DgQtaeTXcceFSRSKy5DplGYip1
exgbtiXI46HHflQqVm7qxZs+AsDUi5VCaXU9uHCS+E6dZ3KNJdRLrmo4rmj4P877
N1F0faYlP0BhhtoDc+tQl/dS3x0PBmWPpnjrxOrvpWu0QcVRzIICdr9k9QOiuI+Y
JV9W+vFQutWG63L/qWV3Z1FZfgWXWCKVoTsj7/0j/pZyfHy2H9CyttREVWurVm+M
+d6mf/DknZiyr6Hwx5T/EGaETCcf1C4mdOkls51/uAf3q2uVPh2ZENA8H5/dKvuA
IJj+oJFW9lOIwmPWaBOtgKx/LzAR/hft66xL44DhZDSpKMVJxfbwtcazAFBttnRs
6UUWaQk4KDMaoKq01ywTp0QpIt8MFKJb4YsXCdsBq+nu5j6j0otUZh45/NdZod89
cVciSW6FuChFQJzoug4PJ0J5dwI3H1DzN3gFr6E6XymTiHFaycP4W62Qc39hjGZ4
2Af+vl95TbF2un0kI6PXI9DT+SZ2y8QM3L9XDQf7ZZMUUbpVTtzXVbmF5iPaNJRy
p1UiI/RtgcTr/XKQE/wPZIyfgwIXPnpc3H5DbKPnooEnsFpfjplUWqmnrj2hReiJ
PgEQu5EndxdNYrp/U2e43cT6omHinQ/mcld0WEDilQlyZyToymARCCDY9dTngPli
K17cQNP2VFeUqZVz1CZo7dOLxh54kEKli0hwbCqzu0HyNP182p7hppg07dDp0KnD
Chj26yqV4iU+YmHzDi86ZE7cBFHO7dArUuROros6wQagyaC/yhMsWRjiyebsYH23
D25X/QV0FWJakujBBWBaEM5yLYbU36gnBfoZYN5iF4Vxx5ljyTtQZON7Pg4S4AyW
h9PiTSDAPT/1McS4EeJHLa9AXADubZuSSg7xcqyq4Lj2Sp1yvN3j4239cUwWk5G2
jelQJxg/iIoChB2xplJkKHfLxEeNpZ4y+pLGp4GX1If7BPb3og/AhqDUdlVNUhCh
HeENTbc9VNKq63cD3z37emYgkjiX7aJWARo2ewLsdZd6AzqJydTphaiAH/L3934G
/1isBwFoPOJpNU0yDWXh/xsFcUNQLxLqYikvEYyE/6NpeE371N0CcgOzJZfI/84/
QC/xW5rdAO3lN5g/OMt/eoR1jHA5f4SLZJr4rlPHWXMf6O4nWXfTaAYMyyYat/Ek
0ufGgvp0z/gaxj3SpvxiQKIx8377hO9WKMosGp1NNrNOWpBLIUu1rk25Cwu/yd3S
LTfoindt+yiqEKZbYzAYDvBuNzjjfvSBoIQzYNya4abFjKzuPT23vt1+qCKWoxmu
SxrtgdHPIsJ6sICjNS5on0Rb+7CzCwcrF5kuwZLvs3Cek4qMDDA+RpYMTUg3eRxs
f846z0TFJPpStnNb/N4b0ddZ4MFFu9ANBC2OJWWMQwzcoG17zF5mwyBlGFN/Z+qM
aqo5JdEyIJKWxlM0SHdsAA4GPAvh4VQsyCSD1RQU+dnYrKtuj3vDwug2kt3Vtr8C
Axyy9kIY4W+eJX1r2ZmVYDs5WPvIVNrwVXqUNyXmxT2+sRQ88xBOcwG2jTGuM7Y7
UkMzM4S0CL+24CV13WHEUw+Bmu3mN3e3jx2T20rJLA7zTe4UoqtulclwJ0atm8At
Y93eyUuEtPpimVDmUEFrzNUbpXQd5eFj8ylNq9SgfO5l2iLqB1ZmxegjzmhFQn5n
M6KTOeHaqk26pU3oDjjK39w4iCtr5AsGOTGkBBmOAeyoCfve3biebuK/OKjFnnTM
SP/78Cu3uZW3o6zjfcH/KcYU3g+IF+3wlf+ZD9UP+uoKTbbW0Cw4uvMNMaGRNWii
sQ7z3EMn2XVW/1R6EmZY92DT3kM+cpFV/jFl3J7/N5ZjNlBYFTXIjRIX6K7iLbRe
unlq1i9m0Aj3FNPRplD4qn/s/dZCXt+KTNjgqK3IJ9IptripoFlTubnFsdsKrCNu
ntssZPKMGFS39tfUGUV2msqoTUnN7zBQntGG/2/Rak6aKJkNwOrvAaYtkVwo7qtU
5YBhuTX23us/rJ+XxjsAj3MhW269UkPomTF6uWZ0jEXkwJEaYnzyWQYU8PJ/avuC
FCvIwYVTSE4zK/DW1Ret/HJmgCNiDzb/iFelFO2YBkjmNf9ZrLUSzmdU6El4BJ6p
PyUlGBR6cpsrzKqIb5E+xjPQCATTMFQK6cU1tS+w+qe1UookMMhLF+2438nQKKyO
kPukT6hubZUQzP6b9JRt/uWXMwPNotsdbFCBLi+35ui1U/P8BEfRvTNFcWv9NUyg
w1SDapDpP6r204gbCMKxSADL77yJ8eOu/tPlAcP4VkMTsObP0UFZW1UxdM4gvSnk
jlPd8XMZqwxZfQ0B+qSdIOgvJ67msNAMdMl42qY4/kdd5Y1e9om16nw0NJvr2NuP
qoEQZT7GUN961GMfb4F6QZFiVvXCS8MxQIXU8p5n7N1X/yjkw7BhWQ291WiDR/h6
+kXeRlWUPsIdXmh3MUNUlz8djHDDvFbSEuI+WqPDKpDtKJAXbqA3zLovqawwdp2r
QLTLPiU1fOfMcW+VBT1T39Dev1yoD3ppIN8aOP1sAW+sjrxuuPDIZJu/Lf0XFGkW
vGt5yV3yrTxeLX7AVzRQp2MRu5u2eBWzgu76GhVUQY8VTdP5LCzqitacV/FXFkcA
dzLAAduilqFfcFt1gJWmIaxzZyvtuArT5rQ8N3xgqBE=
`protect END_PROTECTED
