`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZc7GB86OmZ3OPH/gNQNUOJw9k/4edBZeAc2K6LpCvj0bHGKX5shXccS9TMTlkdz
sjHeW/Ox92AyIYefrbZeHLun0HJYj/hH+QC6VSr06SaYxm0yBCXMZU+BcqRVEISB
GsbNHFrJjT228YZF8Nr8BjUQW6+NAI4dzyNHgYEAbYczHsKRdHvtT6sIhkwn5P6s
i+GZNF/ATo54Z+3c8KKS8WdiK9IcMHUymGgarbFfwNOBUHB6EknhZec9R47KOD7q
j0xaVZkcJyAR4a9DicCTGMFwuVXF9SyCfcSTjdHUFISZi5mVf7h8ku8aVAad8Usa
ZKg6SseFyUSz0dVcXXN9DbdukJw8GJnbCjMYxSQM7eU/tkmvCtjcAu4t6Fs9N+yr
6YoN0dIYDDsV5AC6OGO22W8bJgDGqCthUsxYZyIOFHnkjrnRNGD57iV1XWuTpoE7
crxVk/9jCBK+5Jw4Rqq0ulO3G27kyUEW+OxAMDd1/5+oQ5UxM/e5OxWKBZWQFGKK
4PjqhKSevZcr+06oKG2DddZU3z2daCZIsjrcpoY8M+srXRpdJJXSNdQYraxEYW+3
2vDPzOBOUiLrLUoe3c4IygoDzsZS0XdWHGt0Ip9XSlo=
`protect END_PROTECTED
