`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3fnJnkVAyWb4RVUS9ghz9GitSaVL+SwvejkJsVEh0rD4Jyj+T6moupfzERR9gFSW
ZCFt7xoSKi5hd2uHEeYuRp7ezdv+rBcST/UeJZRsZGhPUDyAxAZqOqFofMyprLHr
t25446wHw95BOCFPeokCI9/PjgqcZHkC7l22h0Dwx8oChmPvvRB6DE3ZaiNJyU17
4EXQcmTxbY/UuGBcSkQtNmnv77PAgG/N+6JzZVpEj5Si251VErnTUVOMvikWza7n
ASTzYg7DkbpL+40Oyj4bl5RvZsmVlywTdMUgsAh/f0wcbrVELJneikGMkqEOncKw
9AZCj/uyuBSJCkB/oJ6EFgRkzfJXVLA9gFif5U0y2VBAXPPbMqqnQi6TceMO7HBp
xB7ohg55ZzzXKTfyncXMCsDGWHrDsINjRtQ6SPfvrt8PQ6Q6gqqS25W8BWZXlhXa
xA8+RPp7YfFjl/cdhqmIVc7YY1T3q80Mu0EktA/ot7XuOMsOpeKQxJf6eqRRROhs
F5ZZmcOPwTrZ3L1gLmv+6eiF9Ul2JGDU3z1vFKL0gcZGmcTzfemZ9sFBTfBVr1l8
qkZgrAZ49sBCRLe2EgDFp9CCmKNXrw5ZrN70aKhPAxyOG90xZTYKUAuZ1CjINUAE
o2LSmz/4+jTsLx21VFUjIRtrHcEKKmMcAdEXCinrCPlOaOA8uqgKBGpEmXJiyovb
XS8tscRAVwa3ESnLlcppUkJqeEtceKv9gMIgEpGs0gnPJ5THKbm0mvZtvhS//bP9
sLSN1s+doQwSj41HNhyBTQ==
`protect END_PROTECTED
