`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bny+WMdug/WRwU2vw6ceTpTKcCyFbPVFRd0byxSPpdUVkEJONxDGyYQleisDzL+K
cvSiLdjvAuZ/G9l1Ne6UIhkCw/TA2+5AGEpLg/qgNR3+JfzEWSq3hU/9p3ZMCguu
kmGER/oefPaFwJEeEjPIJIMOB2jMiw4KkKwhLoGHw0P6Y/9U3z7sdkf7xCsbrFLe
XOVFmXJpGJpiMbczvBOIdnmmxk10beq0LVRQC3AcI+U8KHnsuKoiMQN0rhqgdYHt
2Hb/1KpLdPTM0kUce5iARggJMdtZ0OSJi3Vq5nDSkgIqPwh5rpBCDv0E3rcWDMNE
A+boprirD/I3C9+lQRoMdtkG6fDb5YfNv3RfrmbcQf3vebLQ6clLonQGgeJSTo2B
txy+mm55DEr1qj1pBgnvV0SsSzh00paAmblUOyKxPXU1egPS+wtJokBmUU4Xs8PT
v1BOfAtkrdrOeP4Dx3Szvd6ENLI2tCDc1z9GY8csx8nxMJ5BPeMI1mnimIKC9j4Y
PSHOMmWmOpdZuHtBER4/KjAdBxdHtW8qyfXUFsVTlNOSfHXFrUigPn0U1uDkSZqc
W0myr7IAXloBVj/O2F73XEbJJ/hDLMHihjbATfAEJ9Pny4bB+HvIFlVm6L7eRk2j
NtbEb4aQBnDHhE1q86zGLHiveSeJWYx9k2lskFmt6k0dodlGXa9Lx0rcSFUOltUr
K2lpiacCDYOegliA9a0E2srG+rglfbR0Y6iRIjCqp6RWALRhJi2MdxK0JoBhve/f
4eNegh0I8lEGK04J4sX1itqEqRm3hkWjgNKtwcASiMF9LX4TvPAbQk0cB7qg7P/+
WpDuFAY9l7YMNLqW45Wd5PJ0s2s24ctO79Qvj/6etm9FhzZNsG6s5RmUBP3jnzja
DccTA4sV++tBIoKVmTuowaKgMUwlRKcjK6ecPfR2A7Zqx9xpNf3vEHr3TX9W3HzY
`protect END_PROTECTED
