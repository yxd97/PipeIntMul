`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDts5wIzvPFP2EPkaU0NQWU9B0bsqH6g9+QovJyqxdZkLQi4J4nkSzEu+82g7f1k
iL7/pd4KNry06RhChNWuSmyaIjg8wIENOSAX3FvZsgnKpH6LN8Lut04FA4mNPxa0
PB7IzF213huayr+x8Vpn5fECAYQZ2vEmrxtCPWdMEv1zQyvl2lcb0PxMEjNzlh85
ZuTlfSAPB9YRTNvoZUYS1rAyQbIrmTAHPOZ5oKQXw7pK3BWIKWhvTEqfCGOPCVra
nOStuI99kn8H1VkMb0gH9g==
`protect END_PROTECTED
