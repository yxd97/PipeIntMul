`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ktoSg9exb1VkXokZ5tTyccaHVH/WZuj9AlY2Qc5G1chyKiz19LV2jntJXGVM1TgS
SBi/0d2SA9QgSS8bE9IXsH9hd/qnTuyaYiYzC7NBNtZTbzOPPUKvcIlXAApFETKR
/TON6FBGPpMHmnhNKN0SG4GxyX3SHyO0Flu0897vk1ObSHz5zGOhnNi6EYKJ7JdK
IDKrivk0PCgN/oBX7rDbKZIxUsZyxWyYaJRwwo31TgK18B9Ld+6jbYNhv78DvtvJ
xRrL9K5KxC/0+T2oy3NBf6YaHmhAIkg+GoaxRhlVZfXp+Fg3eWEiybFRMp1NEea3
aZcYYrDiDqj5pIDvc/8KD/gjDmDqCO0nRj2iDT+FVRbxvOH26tiPWvVLszKCceyQ
k/r1v1Lo22vH48c4qGyl+RRIw1sLazoif7o22OrgI18POC41FPyBg+Ee5JQewXFv
Q4fDQOsZCfiNYFxbHrJuJ3ebaWzFHTlsRsS/jSJbpTBE4eaoDTbdMu2L+f4ZXYp3
T26WN8DSdPE2jVKHhML8/lTRg/kXlPQGuLvGFV9l/Lf8RAPFfUiXcD7aDWDaECoo
Ou1WrJ0X1Odq+VxndAnaRBTC9YZmxLpXDWhWHFDz/Zc=
`protect END_PROTECTED
