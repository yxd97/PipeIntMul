`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOAdyXcc/iRvqLvRUBGBw+k8F9r6uvBjoJ9Lg6hIdmFoXz+cUIlaZKrWKaObTwrn
NATfsl5S1U7+0J7FaBUFr9gWmb3tkrBesW2ILHokEnGf5gQowneILKVLnYgzaqWB
L1h5x59KOC7QajCHFlD80G33vxqK631kTz7dh+nReq59zcwmgFedjlDZRBMJ4M2H
GgpziVx9krz+iDXXHGsSprxfGQD93sVC+8hTcxzbUNU8E9jcCkEs1tA6KsE381D7
pz7Ly4YFa5lvPqagg79aRBxkAnj9v2DdT+FYOaCP8v6Ldc1Brl0KnRbVIsbiEQAf
qrVEyw5T5U0HlkNvXsnyw5sNr3ClDbwmuSaMTT1THVInTFfI3uVV1R7b4mgnxMTE
UH+oF1v0y3boWyaobrrUtJNWTzm8VYVBidugjE1vYAJAJ1Ujhakpell4Lc+qMviu
qGd3lcbdGsc0uuEiDMlbNp/zZkAUTaAwfOWvMTFCK/sAZ6/SVnpdKHTuRyFCIJ7e
7cdbTlXv1WqnCQwfzaRc1q7N6kt3XLmB3C1eNWh7N7T7s8YcGH5ydgb+U0oQzCC0
W8FPbwv6jgKgEcOHcK1icA==
`protect END_PROTECTED
