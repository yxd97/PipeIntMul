`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CN4KaOZvQh2AUmWqgli0iREgLpBtMsQzSRGAor58xJ/5pTIGNgvJ6t6WTm4j/T8P
t8ydoW/x4gWRd+mHwDcsTIekq5PezLE3gvsC7hASAw+Hzi/ERRUBNJT+FCLKRrWU
6KG05L7ux4MXBuj8EVCOi66GRaEy/1PBeVZ2wf3HvmcaiGdtpajkk4kqBqcRzSo/
nG4RUvnFPwPYTkNRa+eY5JIamCFRGzWIPa1s5gbdRxXxUPd8hbX/652Q8sTBL2Td
XjnPChah6AzXKqGslMLbuSmq+Rh1B6uIJmvqna/k+FvRHMkJH03D9UqNjli0jMTX
In4bpkYnuAwZFx9opmupQFBk5vnMYKBm3cWSdIc9G51q+v6BJpw7neUyNUUdZ3DQ
ujW3K+dl5KbYNJLxFOcW+7YKL8EjeRJ34s1wjvXX7LxCbSzZiwR/hhx2Nn9FzpAr
buxy1YKmImj7Lyy/w8pWM/HjiVzgfCnfTCm7GmyBYojN6+CwRdA4iZoqyy7d87qw
mWBpN7nIifbCFn9y16W22/AwJDRiL1G1vVL5Cdp2gB8=
`protect END_PROTECTED
