`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S4/79h/pC0+JBmdH2uk49dDjYQ5TkYeCVIgnpgFdur72Fk020JpA+sB8gZwigwte
2zy7M9zcMdFtfGmiuVl310E9JSAn3v6jW6Y0Vcib4x0GYwtBqLBUGL0UUcJB8hx3
sdthCAMa8syhadP+yZ/a+YmAwFfO8dxz/Q/AjhW3s+P5Vne9dONhoIVbouQshr6X
p1tLsSGxRhMWqJoR/Ru3teLEx+xsU23PwjLpk1fplA8vNhh6VWTdB7m5dlZxc9i9
TyhXNNXoAHE1C7gXdccahloU52cEYw1uKsWyImPKwt0KGYJvVNIzFofyqwmro8Hq
8hFw3X6I3GNZfI9MGXGjHYw23j0ag22RXdHwNXhOuBz+DkJVDmBs3QT7HDaWM422
fHe5ZJaQZGqJXXDY9REBvf2zCwogA3lRD0axScrThVNxngXHe8YbKB/C22Jjv1M8
7rucfd0zz6RPcny4HyWEn0fIuWAuRQvw75gaNeKzzSiGFYiGKVP8skHscQIhWmN5
`protect END_PROTECTED
