`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFHbRuHfaUW1YHda2jJVPd/N3ZgAgXuOHAKZ6lP84auGVQSstzuAJ5A3hq/XJDpT
eVyWe+Eo+1G1Vv5/WAnyMF2j0FgrjX38hwR7/B//Jn3xpxBXKZ+TkDBjXyAb08Ta
wrC/ZacldjNdpPXXbSHSEiHKAPOyyfyWlWCLA41RmtuXDWiC6eFWqSGgEJopuAoJ
hXji2uVFCJRsDKk1I5TN7NofXAloALm5TEYa3+yLV7eY16pKiWA6VY9CchwJXpqj
Uo9sDXLAMmubGiWywY3LIeDiNafv61MewcEUeWnvvXM=
`protect END_PROTECTED
