`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmdA1yUk9mRLyUpYMjuFaAtRzJ9xK2/KYCxbjVeOmGsZNh3oNDVpWQniQ3xG/ZF3
X6oL65JOozyDTI2/IQUlkp1QRL6QmiN+JKWs+232Qpifyt8sJOu49BrFwe67cDF+
Wk7G+Yxr5Ab0DlFskhg1gzSm78b1GhF7Mld3dHJIczoJzlwc+2Gli8FA1p4nH1DV
8Uqzp/O0n44wreiPSYMzMzZtM4G7DWt+Fl9L7/aR7rwQV0+mVcoaYbkVN+HqjHR+
958XcQaXTNyndD3ch1CY5b2ZqGtcB9ZYh0oy2YcD6yC26Uff9J7z97KFFqPC7Lne
le9Zp2OmLxCJHnZtnpvfsPQinpNEIs5b0DXo+WLWP7jHWMK62SAAoXyQCwU8Vb4+
xW5HUpHYJStIo+01TLQtdsA+K/a9vO9rH2MLWrKwtUdNg8IuGXCb7eRyRmNTD6lM
edKQ+7yCOhIxvH7Rf7+qhHUAZDpHmcKpmAcYfCoMd+jVFzhfH4Ku97/gSsw8Llb4
LI/ip6g3ubLncRi1Vz1myBiIiRzxXHUqNuEsh5sLWxlPpZsCC31ZFkn2qSL46a8F
pc/Is6RPyRnk2ak9PGEbpaXP6Jk1aQM4gRGuiw5vJmu9qfKdtAo7pPuPSThNsBub
P91BZSSckxsQRpjIfQaITA0e2Lfs9biUX5F0aHJ3A50C0X021jxKmh7fIpRYRYCz
2U9YAke0HE9sWhxzS/ayjY/r30uzrr8utnicrwjJcF3gEDGxt14tlJ9lgzqpvr/X
mfI48uofgEY/cXg9W/x1WWvmqBhMJjc6mZb8q6K3qZfy56CaoIKnKpEtoq66fBbl
aO7qn6asWky5N9SPJjhHsmdGCqC5WM71spfTP+jqp7TjhBxjNm4av+zwMqgQap0F
sQqzI66ke2MZBhCWSHfBDUa0EWxwUCXXCu+8wkct3gv8ccJdskrcb0JUx099L6BY
xrqHP28IJLiWY1MnYq6nxztz27UnllXTfNl9MMu062FOs4XhZ7feAXAyJM+erhju
H5UjgF/PSEa4XjEwKiKph6nRaHHD/wPG7Vr1iUQWTc0pAPD//fa29z+Patvtt66/
l6UUrtBJhuzRoCTf75soqUeTRiC+oRWtDm7hfZdKF1Vouz/r3jN2sbO8EhaCTYWP
xw2lUhLtp6u2XP5pZPU7Clsv9Bd42Us2jyXDFQw2NFTO0lv7Aau634oyEwFmQsOk
xr4V4iq36FbPyCTJXYPkFsJc9oiCi9rGwXeppYqHH4EeM8ve+yVOki6kxSyelVlm
YDYEZH+e54obYNiqoi45HUveVPRKElDMO6My87z1ph74H5q7NI4RJVdUH2YnxyIF
LElcfgH84E93tDoYdLPs2tW/WqP/xXgyEbxS8d1BStPwmcLbprailV78RKjhi5KR
Y7/xSnHTM0r0xipcaXdEqLUw3lxZ66G2Wysqzz1ZyVMTiqZD0ekX2JAd5axK4Qzw
BUZbneKF73PSatS+q68JZwo8m5Mc41vZgAPby6Laf3NUgg8pd+IZCjWMiyr2iYRg
NqlmjG8aSU4zJswEkoEbLCv6kNzHaUmLfdqKBZ7Ez+TViz943TZicnAj13CI/pT0
Gj0xC+Zap77QCKVysOC6MASlSyqd1jl92DkRtK9J7vZMT0tCaE831Ub7abLyn+I8
w35p0VLt/zkU9+AjFS4aJBgWkXI3iKHgJHlgtQAYDbQkWf7OEq00TwL4UmASj7Wo
kS6sn9Pr0qNi3AAmNJeQJgMLeXZooGzG/P5X3eDRussWx/sBYf28Q6g6bdj4gHb+
HOfD4WmZiLoZOK9K24Kc4CyNIdRQrdZ0Mh1IQwlWlBKPBkz5MyvccWU/gHoUnPAN
5UqXkD7L+1gbi+FZwqBIWCkDGBgkF/rlWvq2X/hnLh4t8quxiP3jK7VBcGgT6ChN
islq5ht1ReQ8tXKrom2EGneLxWhoUL0++QX6ve8H0zvZ9nH/nPSVYRYBBp6KCk8z
zJE6R7HCzLZ1G8r1rLHM7c5na9Z1XJhhXVMT3CfLxi7e4WcNqYFM+hfSa4QxtOlo
16b0QWTyvnM9RtTah1+VoksiYBcSrrrcNzprUvbaJuKZL4xicTyXwl/15oEAI6dl
81kh3BWi0wmeVANeD0f7moF4s2WUrg9Ss0ALkH3ePIBLy59a8xgbkLcK2+f4Q+uB
yl0AYlaQVMKfzMwLmeCMl6IyILvQ3PhUA7JV3Vq9+STl7TpGRH+ZuXh2wZ0Vnnm8
Pj+F7OkeUAQNBDsky455TmcRW0ufLbTC/GaweCoCYv+AtCOt9mJO5B2LjWZXzOq8
BX0kG16PZRjKfGE/x6YmjpmmGjMBpui98jNZgIdb/d7xRZImZpGSDYn8UsVEbOk8
joCu6Hix3CahS8z/M08fYByK6vmi0IG74ohfdCQ7g4Yd1Q5tNHQ6BPX6WskKXz6I
gwOsZhLFvBtfGp053vlNqobPETdrMRCsRbFvt/GbwrcbXXm8J9qRe6SxoqpWdJ08
gnsm6BBc2Pi2tkrbv9cQSzlRv883MBhPrvIsC9AKztEiRwA4+5EGexx2SHejVh22
iYRxDcAF3yteMAKrqnb8XJrxzZFlgp+CXK1Conov+Gopvmny+Vt87bnRXHugo7++
yKHLP7RvmRzoM8FUYQU1fAf5Jve6dANYmfDuHLORy1UeBErXS5253Gd9sSqPFZzz
H0NQIhnhOC4bHa7cLyW0s4pg3gQVJqlLfssBAbqBG8eXjwzPdp6FFIPCbpdIx52R
JCQA8SydiO8C3QWiY3TJ9c19Kgt/70pbAWRznlXWMUnlJKzwTY+YrBMlzlUEskxl
tE20jz46o+BgGrmzCZE3ejs5B5jycvM/EVdnjNC6XtJL+rljr8bNXReWDxsDJSrc
pgvMZCIQwa3DPIs8Id5EclH48WdiXbeckGu1WDzx25MkuC5E8QpVjkCTyPv6s2cK
OyFYORyQN8ooRMOWdRDfNKCKVHgz3yQBKXxsfPJH+gGYy5JcDxORzjfNQAfqZeUC
ujs1wTvgL0i4lPMqeKkE0wni7lCFB5uVIcRGs4s7j8DWY0rzXtxkgKXVUVn+wERd
zJdP2i38nNWDf9PMrLppOXkMEthowPndbguTxHTPtlOfbwUKb3q/AI/hNC4zmcMy
u75BWluwxG2TRYM9D58xneTwTCpxdXkdPHJjF4FExVSX2WKUdv2k2iOMkxKl5IYU
y8jZZo0881W4Oc44AloJENyHyrW/g/rk2HSy7CqS9XJk1CIm7QDwmQDp39wHmC/j
CEFHMH/8g8FFR9j73HwD2DTbxMUj4u8tV7yL++5poVUbxZoaXqrFNywZ1kUSuGPQ
K9nKbuePL/B52o3q2zR5/EHgr9SKIezPx2mMjnW80ulpqdLO2RkLNy4vDY/VCXgb
a8is+lQbrgFfwEeJPvhsg/wFoMjWYyi2FuOktONDXM7iDSko+ZjwcfgoJc1XYtZu
wdszDOvGrSJligaY9F4xbTNVbiLEMLmPqLVfWY5STObrKnqBWW6mxv/1IlXW2w1M
/sjdR3Et5zAJ6I4HmpL5PNwwL++OdBOod42n/3JrRfBGfbml0dtu08zDC3dJvEFT
x0WSMc7+veIETYjnP2O5voyYU4dhLrw3bXvymLHyxV7zt4/3bjqYKNlswCTWHZRo
c+qTPRHj5M9lKaSoUn5c43DJ9qspBYK5yi/Qf+1ZgDZWcMrBNpDiNVsELJQPUJfj
+tJ5HwUz+TgWH2/XktEVyxAssk9dGMvf6JIDTFIXg+Dfv+m28bcCvJGH/3/gvV5E
YAZ6YL+3HlUOb+3KiJHNiNK0woRi2Ml1HyExX+o3jvTCIPNxlAiV2riM0VGpWr5L
PGNg31WA3fqoSMJ7V5PjvoU3Vwb9bXYqnP+6Dh2NcblWanbVcUC5Xrqxp6RbLXTQ
2rYwE22i3McAUFP3TbIbBy+0sOLprf7UOa8qOpxoGoPHvVUniM+xoMdlC0MSa7/z
bze9IbDPGtkcRAQLnPbFPdp9HkAq87fpA0uPT6EFpVNdnbDQBnjyPiY0f1yRoyjF
3mmAD7VyVLuYlmDB0hl8KvtrU4Hr1phFblHNnjLlJVHqM+rgXRVkj1BwUqQqD/Yt
pd8yVKJbNOCu/HPKu6RcqVKAd87hktlBQS12g2RKraNNAwgyMZHPn4rTK2llDrmB
wBjHjJtk8q8/KiDCFANDfb/kGZ6BOmdZKq9Co/buwk78qfTcZkrJSVdKiyM7+dZS
OEBlXlyBsCtPuN4v8cIqV5W9PM4pKMXnJvU0kwMXTTDMUOWhcDsjqpLFLf8VHATw
ha/mMrP7tBEjnsexXTlZHPG9mFDjHYaOq861Xy3S67h+nVuj83+xU/bM48mKqN8Y
dm1+SPUUawEaozqLDoGwqA1BIHXHuSXGZt/Ibb9XQBgJ0mF1u93LoYhR2Jz/koKV
cNp8mWVTCta2kIQs3m/gyrLNkDL3H+H1leVQy9yeT34gspHwdDOCvUjAYRZqDuwR
5Fwv/eV13dt90GgVzaOsSwY74M3whBNg1LbMUKzP9kbnXuVkTfsw0rUslZ/OAsuP
1zHGk7goQGHZa7pdOT2OuKzPqlqkTHFLXqDpYKhTtp+VQ/JpdbgzEWB+Cy46D1UW
NygH+gq6iLtslBami4veKQ==
`protect END_PROTECTED
