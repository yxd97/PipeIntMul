`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZBhIVtbtDgMGEhcr8u1WmF32viElr/ahzAjNS29UYYsDVXNfaqvapYCnV5OoRb1G
LXmnSZWRm8Jd2XJOovhHd0C4Bcum5UhVIDFdooLjzS1uJvaF5XYbP28UDsVLWxRN
HFPB/Wy1wLum2vWdoKjE7j3FeqPbv9ILz6LZ09D553dxVW/CMf3wXXty0rA+0TaS
/jXN1IYov8E+L5Ue4BcHRcEnerfOIoDCTfRkQKPnPrdEMf2gOxZrwSNY6/XRVM/b
+N8UpD7HCD7cTkJbI/alMjH+No4RthnLOiyFlzuUxdAdi3ux5UQYG0doqhRrT/9e
5Ff8K2LV5BR7Dku2IiHtNdxs4d3/uzS1qzq0YT+xN5YKUv/pXhGBhl/KHQIe8wbW
/qDi54ScdsBNMQiuC9gTdxAMLymmigwmHHqFkXrWZ83ZXeCV2z7td6gMDKhlmFJf
zz2qafzJgp14I9DiBQUPK2/+AcZ5oKQRDIRMJjjzX91hNSUQHREJ8/1KOXDnmjrQ
rSpdOeNBDi+Hu/cIkCuUNEL/bqLcEC7VLl+s0m5dg6gd+QvRr1zDP9t8qo9DLjfl
JT7D2QGP3TOPFqpTVa0Uh1CDrKCKb/NEJRqQJ9KiOp2rehJHKGHZ3FpjrpgOUeJg
wZSYaB0fRjqjzZH6gHC2/jeWB56jjm8nAcxDnGY68uNXbWRGyLkj9riYrqXWdERD
eA3H75k4SFRpzFma6+jNGaAI9N4Q1VjqxN/gLXsh/+Fz+qskO09YpRe1qZ/+lRLL
7gCy+SlUdKhqYBGZzJDDfNt7qxQRHwiHmDyv7Wsv52dVTvICPpTnVPho7ILJJSdK
U8mRFjh+Cr3ucS5us8YJpk8Qwvey/TMnHKlBD/rkIXD3VqEggfdT/in8f7zetuIe
PdSKt81l2kAMFz9Emj79cW8dXq2Q65d8+bE7FCZwAlLeeOKoCz+LAG+tvMV1UyI3
DVann6rBh9efdet0ChZOoPVawLlVPUJajtkC92ss6ryT4QZJuD4hvNZtr5IyXGQ2
kvbImpv1Jsb6qsf6ddYjYutwM4z3p6zHc860KiiHDK0z4ENzKB4x421t8ZeeesqX
hB//+aRCuBWuwERVQQ/IYTrAwtOS5a1lOWKgJqBpSG6x7mwqwd5V2Ydkn5r5n3n3
JFQQ58QVRiKTWEHOBqcTqoTqhNl+3+oyWwZHOjgq3CWQ9q7E0yGIaiJP2P5GBQDf
4ATBABLIPDJb56+NJqiNxBAuHT+pIs5XYJWeBQHug2LAxrKRoSpbfEj0H0ChI6By
cubj4k09thwSFfNJmO3ms8AlCAWIop86OGgSltdQV6ys18zLnXDM8nNXyWisYX5U
W19U0jyBaUZTwJ5JpPGAqdF4nF4If3i3LWyuqoPsEkxsIJj+1AIcqkg3XVDjAOhn
ZxfH5ZMkxFh2BDHIhtpC7TCgxxsa1oedtnfIDoGKNMX/3miz36rS7SMgfU/gqwxN
4sPfmu4kRwK0tjMLLG+ZPb0flG+EIrAthbzQ+SjuR1E=
`protect END_PROTECTED
