`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fHGo+gT79NWDDiHtzyOTcgpkk1d3YyMYr69iqGYuVZgrHHrJQMl6cL55Eo0+kzAV
T4IyV0SSNzqE/29kJmVibsidcIA05+mNK06SJQe+jx+NI5mPE6zYjYIb4vAHuBMt
kios4qCPITn4ZUd9XMdYJUQwxQDg9blll6JJiz4hp/gw1w2DwJhDtjL/i4+LcJ+k
AyGLpSe2ugrrM5B7J5RqEyzguAY5TvCUT4U4sd3v3W9sJrrvd/mGDkElcHMRgnN/
riXC/F+6q1H1gX/kGKVXUvTt7L/0zDhR3EI9EoYcs9EI4QfFB3OZzddKPb8W9YNM
Hhh6bi5OMCnkf9vTKnGvNXltwMjmPx8h8lUPw5Eyxd8B3JCIky8yZZiKFUT54MMx
hjjsoBDxqiJzT8YwjEP8Rw==
`protect END_PROTECTED
