`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44YPldktOA/sF40MXQ2GTlT24NwSgioa9+CPuTFozliutPVa1QqqzkdA2e/PjMJA
cZrmIaikA8MMfD5eiC4/a7YNdyOWjGOYdGeJbKHWVD5PZmuYk5yaqAeTfDD4WmdR
yWgMvVpWqydxdjw66cwFGInmleC9VNlP12IyGLLzVHnhSiciZVzK4lRPtGfDf5TM
/vk2evTWKAhI8+MpJpc9lLynZQS5MNf9OnnLfmuT/Lild7EQ5qnUrENBL1UWLA+9
To6kDbE85OzFI0VNpGaXDg2RL6cmPMGuLEYA6eXu1DlGHMie4VKNFmN/eNoyzd9S
tDhQSrQxY8tCszQaEbin5Glby8eklrNOKSFKrAudsORPcg2XlOzbDEJFEijZrBOT
jJngEIMb0cQyYi+JJ2QjokNpCYxyTAgjJ8Eh6lGvDYqIp19PSbgbZeEi9vtm4Jv5
pq7q0ZtBrUkrnxobSuEJCAvRbAdGTj/s1LRVuE328jPEk65Ju1OYDykbJTV7rf5J
+xTUTP9IOPlMb1iikVxkLGQGCSRtHIjk9eBcmKzhqdoHdgBD3XR+B0y3mUZKf8Zb
l6ae8dbD3KLaI9GSXFCIQiigcNi799tOznUmIaHXzgKujgE9NXMPfY2ptvAFZgce
9ilgTpwQQteYUZwKUpa1l3mZhiVjYiGWi8kJL2kd2xYxIiPPlqLM6ebtVN6YeGmS
Xg+cajM5rloSumNxQYmHn9uD/jLaLGCotncA6s+KQO6pM/fMzonE70B3NZYFbzmV
AhPDTqGhDdAb824XYLMt9/P08zPTkz3CuYh/cM/GU2hi0PhwL/TtlrXd8HiDCyTP
upPbueOB/4uv9Rn/iHeHfsBnmH1DIHVGWFduyNUY7lK6Kak3I/kGAm6YE4Q1NkrE
qkubOUQqpd/AzpvIkM3ZkCtVntX4Q5ft+ZrEFY971cIORhGmCHjybi3ccRQxSzLi
74aYD+mdCMOVDAVFaqxNLWJ60TlVm7LsN+813ktOXUU=
`protect END_PROTECTED
