`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqk6BVz7gZRWhcBCqJIqGMFG1XmbraH0SaR3H8CPRmPO/2UqC+cSQM3hmRY05FYG
J8/5OnsbcJgxyImFGALGRi0n5wLuh8qlgG4FpYLdOs84CokgukLe4R2/MrwRWOyN
bqw/yGClAkQc2WPmvgslb4OczvFT1hRPAQNxamolrp0PMOuitYmvbV8UUVLk1mdF
2ediXxNAXwAMef5mS8y9t67+XCoGw9U8Jd7hMhy6L/UkueHYeJkhek9tG9K2+MqF
EVangNkgE7Gnzp2mmhg6IeWlogSb4rQ7F+hq5JLUqk6k6R5Wb/wfE8S04PNifvlB
XeyJSQKv5JisCvNcBGnOsA84HljjAykfJY38hsxKlg+s957Hu2ctIzfqkJb93uDm
YN71FLdaM/F7TLf+ulQRJm4ZaiIlQ8VhIVkJwDcIWO8fuOVTFMyWGcgAdO36EPTU
8WNN+40CwqIPGvgdckLd/l3FehdMFAmvqVvHzo7fXR8kvNClmyCvxWoopppdGDwB
RVQQkxPU+BvFIxDUpOVgu0iNmkj3WpxuaEFfN+eSP6RWwM1jgXx97giGimvUgQtx
vDVFtgZy/d5CE3Q5K+bjpMHTutaI/Vg4JseCuEfkedC0vuLWsLWChQ10M7QxrJBH
FIGRVUzSGkunGqErvncT3TRlcJEgUNFcapRtHdRJarZeWFSEqmTK/pvgOx3BxSpD
aC061qwpz8JxLHkUbSgl5EWJpUv4u4zFqBFLyEf2r3/KdHZVDptam9OpYiveY3f6
eHDwbxjgE5A9lmZBhVKVFICN9D9e7z/L1B0D0Kohhb2iI1FriguM+NSjoIYPsXq+
EEQIC0ArxOGkCyehVbZhKB/YMdmPP8sQj4FD+9Bu522B28aNDlkopkXuzalzA187
fcAtsSHgYj9WPFvHXif+OcbEJUy2PsG93A/M3FZ5hhO77Xl9NaATNT3b8yLOaB3r
sx63fL5FjmFmAFjiQbAmuBmsMnK+A4VUKiN72G3vVXbuGtZ4UetZLBvzsRiZYsU9
YF+vPothMHCdtjxxW7dElsjhqcvtiRHa5xNwdPD5hMTf/Cal0XJ4QgPX3PdqZ+GW
6M1BbfIbqFXWJBVcNSENk2rSwvLwAOcLbYcvZ7hCdpHIAfbwKw2NGVpkpeMX1qdC
`protect END_PROTECTED
