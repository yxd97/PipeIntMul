`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nF4ld5ju7FoOVLiNH8E/2z4eEjfEmHtVH0J2OFhA+EM3kHIr4tuZ5Kf2QmJbASZf
XU4zfFSHljjDNoc1h7eUJ0CsBLARtoA1LTGGQdHJ58Qrjy9UdTuQjb5poISmdA/V
zSm1e2QZ+1BtdSPnwXuKetWYvESdERmh0rAdXFfM3c3cSSSI/v6cpiEhGcwIUmwQ
wp6HO+HWPrNwJYC6RlBNet0L6ar2R1tTuvrwVbBJubyrJ/h4CVRXfJqOxKVaqThP
hgUnEY/PrMQ2piaG8T8lPlMeWHwvuO28MAYtsI3Yv+hmDBNxTVTWDOxUMlcubQwR
sa888imBD5EMEeAIIlJnYQ==
`protect END_PROTECTED
