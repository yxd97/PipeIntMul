`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhj32SF9DywHjAhDQHt88vWw2P16X3Lbs1pxlLzobHreGIm7VYk9lIJZycuwtkio
lnBk4OyvxqtirsyuUD2VMUqAWY1XBp8NF5rnhqah6awqSj46QhyimmYrpO0fOsno
5n2zMaOUkvZggXopDpXKSU0XEi+3KdKI6LDtmFNXt9bsbuqvOf+POYpo+R+2NcSy
/p3ql6bf15do3zrrCwmpcV4vOq0IyO9h+HwJMKtdlu6D7+YgWwg+V5/B/7LSIYYm
DzhajvLtML6KNEQ3md7h/w==
`protect END_PROTECTED
