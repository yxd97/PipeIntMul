`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iUxX68LLePQRsoAokws471OEkx4UJsoDhzAMbz/MtEJTG0xLK2eB7T9iy74j+tt
E/TEpfnIC1mrxuKFBSybFUi0a9jqYhWeyf8Ix0DAvz3NKhCUvlUrHAAkQn80nSFp
HHtfFQ+O3lBA/eFs+wf/ffbty5SXzQUC2iudvbKFZJCtRPVv59nf0vgf8ByTsn4M
JA9lScbWUGXUynwRxs4vXulYlqdeux6wL0LUDwT546q4FcoBv+49J4/NbD1qt7jT
SKlrs4C92UaE9UL/xGTZRxru4dHgMSDol+JkystQEcr+8XSUwUvQemK6rRWWufk6
1m60sO0+9nrfG/O8AZNmNlfOPq+PeiXNX0gEmJqLw5uCdEjdiBiii6z2OS31+utQ
3h1dbxi0lQb5QKo26qkBC0EWx50JVVznTDSp5CEBC488diNfWS6o2+SaAJAapFN5
IjvZgS5Y+yFRjFWq2a23n3y+FyFIRQBw6CFkf1v1okp8YB226qcLAwdcOoMwpn32
nIpN1F8BS6p+v9Kyi+W4m5MNbp1w6SWIKW3cxE/BfZvoN9F1t+cGmE7iw3TlU/0e
kAPxd70ZTPgEf2eXdjX8aipo37iAxAhNbi8uVSbfG9QWMt8k7lCQ9NaaZkA9R7eC
I5rQF03ZGnEmwm5G+GXlSc8FKFu5/AvGQAeFSdG3jPHWdDJV4OQKdRdq+rKdKseW
tAPAvMWePdS4UdPGHVTpqg0ggYh6BQ3mWxqIIAw4HQHbFfy/MWHELD/RTYl7XrQX
x0O+af3qfUuLklkIA5RaHMghulxDWevBzQmuyofjN1/ioii1ZTj0a0+58M0IF5Pu
9s0uVuM3CvyJrtB9IhA4ahxC6eKs+S+nkktgcNRQkcu5ybBNiYG4KJbllZSIqTIy
z59G9zJGcFBMrtgY4NmL4ON0+KomY1Ymip49QbXE6nrMTDemNVa4tjH6jmbcTldw
h5A7Vs1HH5WyUhwZM4c+vS2HQu+zJJ6Y3L1OenEqTrP0TryE5dRzXhuHIg2ZOcNb
hp7rZUZ+mhNyXWDKDtwj/2di6IcfoSIs8mD1Zp4R4gQZMGDj36F7DiSTpsOFp+i4
sHNDxOKc5m8m3fNdynNPKohCWqqSDnsbnSyCGOaPTy5MfW6zu2S6pbckF33PkIHU
Q1j1BuhBs2PWaOLnOWSNWx761AHWywwbztpM/466ZEt1AueT33gOZCjrK/XZ9aUz
gKzkYW0LhCgvK0puL6uL9Wq+Z/ub5JYZOSjvBJqaTBW1ZgQhMk9bDcjAz5/truQT
`protect END_PROTECTED
