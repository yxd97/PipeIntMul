`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gy4mRa+Jamilfvzr50sgShR4Fdg1TRt+259OKIVgKGiqySh1KOYT7SvcIUI/QywD
gzY75Pb9G14SvbikbqjF4nRYanSsaTEm6o7ligJuPxW4cdNcgSdLHID0RCkveZlH
XZA8N/vHEtAxPJ6bHvKw7YOpDTXXORpglOEb5GKYjplxOmlrIL+QWGB/mKCgpzu+
ZixSyXPDEWfyC3G0OW/DQ6fBH+8KngdCMZh5y08UETP9lkgDY0bwUF/U+B/eKCO0
31nbZudvcMqqkCUnbpdXt9eWvv/7Gf8mUSVO0LIvQtMX8LrlNPXtbkskzegD40LC
pvczZskIhhpTNYpVtWwM/w4HIUWxCm4l30vk1dEQAcLfuIxxPBNmj4kKFhqCaMi3
VMEfl4bXzkNBzWD7MEo1hPAa2UbKggkphIzVJbc53RuvxeXS2XC9t4/kXLsm6wwW
TaP3ccWmdMlkOEnmhaeMDz7wVdzLGk4WnSZR4tMBNLTtb/LNPYxiudd0EWT22Ayu
QJAmtZAwxheNk6bW5VxfUB4oqrwE2YmX3cOXSF6X6ZyXFs3AvfUuwra8/7JAbxQV
HSEtaZIE+JHQL9x6HZHFTnTR16tFFh/X3J5gXIAjrj3NiKgSdT97Ez+qiJd7P9EU
PcLoZvnc7CdcB3PvyqN86kSV9QcLr2/atnJ3G0It3ua+dCfZo7D8Jr7b/eOXu9wb
`protect END_PROTECTED
