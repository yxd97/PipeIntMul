`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Caaz7nV6O6CwQ8iew70QFyutdsbxpee9w8gg9mBoA17z9h0gWpcPX/foRdstxZ3K
U2NoiQXs+bH9jGdLiHHbcQuW9HarBPb1o3aSvHtM7E7Yyt7OmN5N5Yoijdi/NDp5
38VZlVoDUtzIoe5Wz6Jhaw3fkcdqwWEfN0R92pp0pnq/A+kUyvXmbE3adbjRlQvX
x1EC8B8MnA9MoUt77Jdp4sjVemt8orA6CuXvvy6Ze6T4iaiDQzIDV0xfV6crc7ie
N76/b2YXm3jcGcWJgPKY6wDGByChvUyB6pAJ/MtaXlqTqmXO1rcGbyt66fY+zuXA
sXlwo5838C9Wcj7TOmq/YsHQ/rW2JbksjEPef/ASrjcxo/kwC1W9dR4MtXZhkpoT
DPzTx4I6LPRg2Y3ZFsyvQH6IfD8d7shuTSxmNZzO19Y+KQTp1g+1IUqICLngE3u4
a+3aXUr9FCOHq3zNFzrew/AXCWAc3rhUrD0HQALk5YBHwyfMAaemdZ0CpbKUK+ZD
lBjI9GyoIbjO/6QweTOUKaLDnnDGUYQsk++wY/OAldQS+3dCm7P2/FHnN3/QWRnE
XNDTYx81IBwCEk2RdaINpPmRr/uhSpTuvlDlihPGT8cN04SCbLa+TaGxiJd7yNXH
WjZCpHqQnQDbbKwQabvbYgkWo+EOOM/Aq2ZYEHJKU0I1Hus50I94ovho8PEa18UH
Ab/+NOz0/0iYj8gZJlHeMdoIXHBEQRaQDXEFeCuKbDEtFicj+gxGWMXQ8BPiwzP7
9hFXCS53orH32rybP0Opo30VsaCK0dNWcy/4rGD6PuQ0//9RFHgB+55b6wSaw5V5
XhVfQmdIHi7EarOzXEg6ybxuzAwb5q7U3R2/UUKMnTWqL8pfkeJc3ZzU2yiUUlml
gAx6SgNZ0Hqz4XyL8+VhWpOP0zZ41SkG9X/k+wm/tg0vsn5LNnQJzr7sZ3dmeWXu
zAv9YqkurWuG1Pm58qMbc8c5DILO9mNR0S6UGm0lHTHZEUWgTq47NlMQBwnbo3Yi
8oRevwOSu3X5xb6ojlACo6ep/nhd1tc500Iy7jO2WdRPzyEHRo8GreSDbYVd0r0h
cycrI90TCqx2V3FzjCirgMokMj7ag5Ka3epC1Nmx/3JX9jRyhA3ERAKz4/ZHF+yE
`protect END_PROTECTED
