`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chzfsXiHFgoyoATyEOcTSHiKBQ5hDR+FuFBDk1KOQAQUyt8+FmOKDKVYEP39dAdx
HL1KY9/CBV/ne4mFjaxstTu0UEK1clEYlcyVVKhljOAzsjtZ9vHjaDuc9chfAuFe
hwQ9DMcDBrnpv8ZCHGQo6D3Yk8Xhi6lz4omCcsl+AtTl4WU3HSvy72V1MRAqcreX
rS5X/+SP5bRrydM6f9YGzdCBb7/MDwxx8zMJgXAI1GW2TmPvOvKQ0Mm0L33VQ06V
fNIIOKdatRvdG7m01p0lCbcG0q6J6npKEr3Mw5b4jj+WeUucTPcpcVg9CcJb6Q0U
Tzdk5iIjYAUIFZoPnSQsDuAh2neFwIb3TeehYxN9sYhMTlrTUTXWi2+GFhAOZCkI
0h3KQJ2SfwlrcgWzmK9wEClyoXaIxQ1wx6/eutN0cdmcHoHEcs9ajGhbiEzhgIx5
YoHzF4BNGcsd8gXZjRiNNwiJPGB8CZnqmrgrYvh59jDiX4SA+r95vSlV2iqoB177
1wEUh7Ec2m9vVa9Y+Ib2sENGumn6BhD/yTcBuzLViL/4E60YoE9J4B1yHBSuPHLH
h4LWV8ozvpdK7/KyN9tFnklT+2SN08vkh6CV/17FNRi27qk5rncZCw808giptkV7
vNAYOewBDSLxLmiYQkeu7XwuhtUjvcVrnLKbwO49My5q54PdjBAB/RJQ4Q45+hsA
XcrRR16sEX+yMxwdpAq+kVF+WI1dI4tM9Ys5nfHGrDjHfU2TpCLewc98p86Nj6/q
/CrtBJEqhF387kER+S7XIg==
`protect END_PROTECTED
