`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h3pNd3BDCahDoNDpIA7RDQ9Elkde0LIhZqZsts+u6RI+S3Gc6LQLEnOqkPFSnC9O
d3n+Tph8HxpBOo0hILBCP9O+ixz0qWvp37wGLE+sSgjOSNU+2z7GFVe7MaToXTYt
Y0qkYhsNzWyqBgfzKGRQ4e9vImVvCN513+UIeJV5Eg+XKMJovlv4POkxQZDqESI9
S9lAQKQDqJ9gVfjPNDn0S+AKxiLDbFGQp4hXSGigZAxILtfykeLwVuhSLJisgSya
/8X8Ep+WZGJj8jFLVeTPMUK/KYeD09IiKRgR2JeaIsqMKca83m1kM+yRgtWXqahf
0bkJPBrlWRsX/WZXnR97U8VUONOrwuzGtvICu7OuW/2rscWuJlufLXk70IZ27xQ7
wIFVhyzEzPqGBKVSl+5FDwo2Ps5Vk3rS22LnGs0+RnGcqPHuvGxItNG2tLB1BWyY
2KeGenZbLsPHyI6yF2opm+m03AbXWm5Om6EU5RV7AdDK4TtCdPmJ4VjY9EzSlloR
`protect END_PROTECTED
