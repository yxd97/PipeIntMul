`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuBUXpee/hmHz8YR6Xa7waG6t+rlqvAz5bAMI6uVDgA5qv78cdfmF3pp0VbEda6n
gHyK6na9N6srvYBOP3XR6eXC1oPvwnrYwq/TWYVl0UXdynCE1gbVazbZ2bf7tSUu
QG1Jt8fxC6p7QgbpFxmx0KlPHWe5c2ECG5BX4olIrIXO2JjAa36KxQIX9aqQ/9yY
yQddjHujWoSKeXK3ek8M5xXVh31GqSAVJZYirb/Tlo9b+9NnaSYMnX0YEAwifiVD
KtEhmWq8CbtPqIGPOoPB7MhK2EsxVDa/4LnR7rfPMr0R6LAZH8fy7/i6Er95bAkU
Q1aOVR3nZtE+gNRN/LenoWTs8rlsrjgyLEIAvyZlQqYSpykXBEjyewu4ILDYlN9W
`protect END_PROTECTED
