`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tpI6hSq08M6H/6l2tgV9+361ijchtE5Wix29ggqud9u4YEPOo/PdhKMhS0jPemSY
8GJxtEaiqITTb+DIaZdOgE/f7Mi1tbMFgIWeSBHKAM13s9JEknflZmlKaWXkiAuk
ciXKm2BHcVGdspEd/KVHP3z3dzdQC/4Kpyc0nrPQnBqDycjYlY9f29YcIud0S9MQ
O2aO5N08ANIy5WuTfZXMpVTaSRQr+23yIa2JpbF1wo8H9kHk5oeH4CjjY0UyaXC8
SM9TpHVtFHBLkJudj4sEsJxyaVkbN7PmMhr5AIz4/jdcYIqIbVfWCmfnDJUqVOe3
SSoucnDJVbRs0ZmIWYzVgBSrWJisGarnliQpqIpKZ8SOl5+8Oki8AmBqEGa+RDqC
r/0P/ZI0TlYsffCPWB6wMc5/bbHnFOdAaPxkt3Y2W4Q=
`protect END_PROTECTED
