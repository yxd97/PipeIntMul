`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0uzz3tleIxxdP2JtOtxEfapV3O+bp3GXkFzbkn7bteI+3vp9qQqACEty1K94hTD
zMdAaGaX2qo4B/mNahsmJ7ZTnhd5EpE/vU3w0p1mCAB8c+MwwPZVgcRhe7pVjQ0G
SOqbiuH13TMqC8n19730l7JJkEybo67VzSvH0x76otvqjXRfJnz54JPZaVVGsBt5
I6Ie7Zo9vDsywofkRB7rFDMh4WLBdsW8GEmG5NP7U1+6CPNzj8ynVSbTRoEOPGF4
euXO3p+nGTpWSQPUltAz0FZRXz7+tVlsmwX6fBZP/5+aMpqORLVZXIrVPnlLc55I
C7smMX6due/pEm/8IpbGb32hwgNFLeVp90UgQtTzJZ8mKwMenP1mvvKx6z3+iAM0
xHeBJQRbI8FKCygzqpuvt3nA+bEnRh8fnEo6Fn5TRyFOfaoW+rVHjKTNnIWZBWfz
RcuNRCplKaC8FLLBj4hkyQe9oZdgEdqGQeSNDmKm4LBeTF3YqVPkMJMPAXuflIX0
+qPqRJfLSQECcX0FghuhsQ7qn4MFmfaYmU2CVf73Bd+/OtcGcTsKOo8LF4TkSNoQ
38b1AkdRkeKv1gIF5KhVr0vm31TO5E5LcKfDX2k6rA8A7shNbfOcnr/MMPmi3jEX
KmQA//dycgcTBYHujxh3zNI48guB9dfUU80d2+hKL0RY2fgJFWm65gqLuFssb4ms
E+4U74FyJNw2ZgmjSSdms5YdKeR7CB1NFMNwH5l4VXSt/0ni/nMxDFzPyYsdBIZ5
NmVxkZIoPKrK+OTf0pmvXrDuiRGYrya134UK2vnexU2gQXtHM99uaO/YKYqm5Cl4
QBNogVMH3wp9U5GBVEAR7Op7omlERobzx83oteaMjuV8MeTIrjpQsmBy2vVaFBPp
SEQD/bh8UBW/spzxy7RH4Rc/kkTMReioj3IHgRx3IMYctZzQY4/wblSTcupKmz0D
vjU9H/JVdz9MA5l/Rqhj54agblPY6dcy2YwYzYzAoqMDuN2c4DW6Dt1RI6LsjTqZ
/eikT6uMXKi+2Fblyy0VycGMXjaohI7LcIaj2H5UNGV7rJALRqIwasx5PdQP72+y
GAoROlfG3xsgmwEwfBT+aYDPrU+xab8Qz1lILH5j1rEih5h/0x8NrlTpTX0TFTsp
LZtYnOmdecOBKRDiER+JHWyjJ5YNBEov04+SCORWDcNx+F33rY3x9H1RJSu/2gq8
VQ+5gKCuTAXrhwSjwjCtlxlLjpCOc1x3mwsNtf+7EbSTQLmvpcddo8Tbz+9jTQ2W
6OcETfqnjlBLqJ77rhxkRMbDLL9F4tVxc/4nUIPYMFGtOtKlS+OuVjJDzYgCpE5w
V6RU7hgMCPzfFRc0RBDT59lCqq02Hu9+SmlH9q66tLw2pbEqRlMMHl1arvZeTV8Y
7i/dJLlGOJBNElCq8zeqGO1GBnbK02w4sXfR+423tHsKTYBszzGW8DcumqLjSA7D
GvFvRN/M9rbnsijmXfIj+Kq0YxfQ/spJ53g9H31+B8Dlq6RKUgmoNJJ2VbYVtZoQ
MjzFWhpZX4+CU/8bckB/Bk+kFyYJsW8cRGQVB3H+t86vhZLxOE+boM7sN7WWAfYu
TBBu3niyRMT3/UN0ROBNBMTr0AITmSVUVmqhYcX4DYMGesmS+kr1TNLpQIJW/b1L
dx+YrwWqYYgwC8fK0U5SRdmP5bTas+V9XG9Cm7VSKYHLKOTIU3PSdurIP8oqsy3g
zEAuyqpY2hDKlmDaWjqZ9FZPduP+5YFPH/WR/XcPbDkEASN6+eGSQTyUyPR65Fa7
mQdJT8tB0g4QRK6iJL+yD2ujWwqyTxdwBc3zmfp9G+tvbrOZyYp8So26o1Khe/qD
vA7y+2gk9wHm6l7EAxEHY+0EsR+14Al/UNaQHc1wpKRLqm3remd2u1oWVl31w4Zk
I7hK7blaLYdFHRbIzw2grdcqaggS2U5F66dLhrUu8oVwjgB80zCPj/n6wS2fnOCh
Rh1itgBD8s8Jp1M8N2bR9CI+3dowsLRm1pKiwulTg/czHOJ8DeEDDtfSDRKk4CnX
E5VtR65HFoHsaXG5PqWc/7rcZ1hdmd71oJlxgXAYkGQou/nPumDZei8RKHDqtrSv
Eh9Pig7TX6pfGcvRCmWprR+pALUmdPCKlKf8aHLJcy4yTALO0yjjvL5oXh/9lwJ8
JJ08PSzw7qtLD/DSyC46v9/cc08kDCxBV1EJ88HjDDMd6uai/kFJRfCmsouVIZzf
88+pD2CTa3VXugjxlfh6FADP3Pm3maoW2bV0tT5QJoKXl4DTIYSZ22zJjZvkUMYY
ZpyM043XLwWyUrVWa1hVs5GHWEtyAZfCR2ZCSsIsWQUb43SsOSeQ+LU9yotY+sVv
h5+j727noTbz02+73Sw4R3z6rjSAJUxwUv08SCUQr+uH/RRh1moJr4hWLLJB81Z0
Z/RRcG68NTsQhHiPMYBiEq/iXWZRqraNRM3/FD1ArrrMZXjH1RN8OIF++jC66npS
Rq7ddyZi4uDVGCLBWC93o7ZKuCnVecwX94hBFBCX9cpWitfK8Wtn05j9pa5GLo4z
w9SBnG2wkN57ijzz4GbA7K9rlVJ02bmooTUoUhGoeprIhJeQBXoCDuEga7yGhiHr
Dw+6P6ftXaTC9FqflPv/6P9Jq6EJYKKVb3/HDCxnNZZH2M/uAbYlcN5vXocppgY2
P/IWPoF/Urn28UD9fRY+br90uscLlpRmO2A/E6ntpaLZHlyepmBobq/+LSlXYA13
0Rjkh4GsOXuXjdM9/knmtm20zfyRYTjWhO4sb2GwcUusTDSlw/eePlq4Y8G20hMp
pDR2nu6QOZGhY4A3Rgva1itqtqE23Ym384YkWM7VFB0xato9ZVS0L2AXVmfvfp6Q
M5TBwa0r62M2G4Y/jV8V8/XMYMbsyM67s94Ba046g9qP0gj4UtFjIVein5vRneXb
E8QqkNdyVuba7h8u+r1poth/GrWiTy+r1BUN4xI0M8HxOLpEGlkyywozYyqFz4s4
eN7zyV6FEuPxQcgb6N+KaZFakq7DgA9nDdsUDoJXSsVulp2os1esBdbEsYQIMXlj
ZKHaPO8PQMyiOCxQyOJY3aOEY2XoJXk185E6cq13rVhPZErpS7MxmK1K+D3gn0VN
/20jzk1uZRbMIIPLm+6UAmuCCDvM6ZVWL7Sl8AxaDa7t3cBzl1Z7XvglumRrRTic
41ixDuJdbZFpAq1j2TltUxEkzB5jvGApKACChmTu7HayDF6EmCL6K0n/bUIuu1oT
a3j+vr/qlJbd7m6mvy96hIJMT1N12iq+Y9HiJjzgjkCWjCO9g2fVuXtRHFiCQRHV
ckUKkgWpToCaZor6upa1zpJgjiNuQsMMtUeY/1hz73KR1mSBjCYTaQvbKrJtMmBN
3tTa/Bpf9bMiA8R/e3BAe5pQ1uVT1WNFByAKSGAJMBSFjetl4Tqa9Idb2HNBorUa
gWqrDLicPAOkwUDqiGnJnrBJbhsCwpNyG/5b2W0WLleozoUUP9qwryqqlZVOcMGu
aN+8ofWtAGaxJGZtMp2rdqfUn/XMsB3mxoqNFPv+dor+vVVZod6SqScJ+9oiZjWM
UNLkO6UpZH8sXQ/8MAan8h2zcdJz+lxxOul3tIYEpl6mBDn7rR2lvcKVqpC1PeDt
qOhmDHxSnbVXXNtkR7yFLsAUiQ1g07/QzTfX2WPPrESShHPPFB4sVl4KVOtIitW5
lgq9BTNpAmYOd7Fwc3hfZCc8BEWiul51kbDQxxxCk4LSu28AvnbYfFzEPxCwbu5e
l+uW7fv3qXfTN++184pajDJYtoigt2BnWbw8mZRICZvJ2xyUZJI774HQ+/TUK3p2
E//ubEyRBPo5vR1wAfwWuuFpaCNxkh7jUGLTX4qdFSDuzjPJ/9FQELGEWPV11wTo
CxHAzb8PT3MTmXIGKkadkx5J9iyI5UjjrWWh0qnI95Uc172QAndT8jHKVYIbvk/v
Y3qop0ZrEDTx+DbFQKOCJgGGlcL2TN6LcpWByD+pbBxTUZ/tSjyswn04HSxJEWMD
SGq4Af+Rg1lyqhUn1HCDz4eVQaem1IXtMTDyiyY5J3N+fmaFGxWxUc0fk66aD1Xt
JzK6ZCXq+MJHopRG11YQqWWVRjqwSoWKTGcrzxyBoMyFe4943UOyE5BZRv+VIalL
5Y6WOrLAPD6S07HgJ8sgu94Us1hvDYBoAurZ+psHT0vVUeS7xRI9eIC5nAX5IS5e
C+GEl0XQR28RiVVNrEBD+Co1LC74023CvVMxu5kWngqZ8rOYbEDLhzlwF5UGluuU
ig7Q6Z/rmAYhRGGitgZ76q+CUy0PhWqgO9OKJVTZ2c+JcDilEySFpIobW1G7dO9k
dVY4szTWfwcBqZ0mP6HAZaSUVYRQ40BSXBSuoGiCtMZAv11vRXMYlQyCDv+RtxPY
aPZrfSK5giYWYM0zL2r70CGSUBiFEBqjS5c4LDcHyc2Cd9R7OBkrzc8xJuDQxnzd
iPYSpwSjMePRTv5fN95c9r1juED/5x1Mpkq3BxC1eChKaKBnNbs5NP3w4226L++d
qzRy7ARONqo/Rlc11rAsI7fFR3zcJE7lL+TiAMXK8y54L28WSwTjygeyad13Ox0C
zwQZFHXle8wPZZV5ZQYAtJO0Mik/1rbugpILIFIAg/RLMLNDlIlVOXnSKZcnJx6v
BIpq1n6eGVQxTqm/fOw3N4NyWn5yeQyCkZP7lzLRsmE=
`protect END_PROTECTED
