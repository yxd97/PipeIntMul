`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KylBfklu2R1yVkxfj37WkqdYzubNGi3p0t2SYwOYKHIe9Sq+No34+YpqxQ8kIttf
ygM7xgDgZ9G1N8embW9FQyzEIQ52tBry2H24cnkFeC6MULE7i4bv4gh5T2MVBjRR
OX8D4J9txVvHGhwWqEdByN5o5ez/AI+twA+GTAIgjHhFwaWOWtduxLBG1nfXSjal
bGMQPpNZ0UVKHb95GBFGy2uWZYsECksl7Wwqj2AO233lyKrNRQ0/cOq6wTMQopwC
+xm/9Sd+K3l3EZEHXJQNMJe1WiFUGz1KLctSdQ+BdaUfKdC6YrRv7DQLsKy7jt+s
`protect END_PROTECTED
