`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6SXIJ8zmx4cm841pTWkiVszyhu9TqB8FjbIxKoQ56V4wMS51fpY9BKhNosCry2g
DL1VjkRgK1XBJU+Yiy2OILrgmr/yxDtC1gafXL6PaHPAwgqKFS2iGxub9ahmHuuv
rDKh8Q1Wy96JCsCtucbUOP7tTQcVVJxScfCwb0b/LdkxyTn3byArexRisb0QT/2K
i0WPkjqP0pNfHGNDPGUxrOSzdmFaAdp2ErndXE/gGY32MF27DFdeM3o+2pEvqEUr
kEYnTzHALwoIK/2a+HTTSosI/leKfRkieVlYIhqLPF5E1iNvQLtQNnPBtuxRWmpx
NsEHs/TfNOpRRD5TIVBgY84OE5pZmEFa4xmgdgwms7993vymVADySUck1uunAd5c
Rp7DbpuMBLuEETMf9PGNatTkYeEdrhPHZ28rx1hNRY+eZosgVXdV26ydmRmlB6IY
rhfFKv5SHH7Lq0WplcWAENV3jhE3Hdv17NWhaK83FtLJOObnuPiGQvBkXWJVGRon
WJcAzAGa8BXFOZEvaId5f/zemKw+eYR7YUZ4OcXoK/wMv+b78//VQiBcR2tD+AJF
2bre5phtojhnuhPT/npfTs4CGHnnRMi00s5mq2Y5IfRBBNilPhvMftoJXYxSo7qE
sw/g4iIXuINxCl2kXCEyKZ+xJ3sLGXvDFZ+e8r/1wbFqhvh1xiwsJ6hzWtcDLtSn
xXLlj2JVIWtoajii9OESKOV1MJ3hL8Xc/4JJigLSx8QYxhuWLzNdwOhT8Wjr+9Fx
TpedWUDWFNAq1Snm8XxLaw==
`protect END_PROTECTED
