`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJNWb3EJzd09NqdTx0dAc/7lGCijkCUYV5sdNb+K0oIHtYQBD/0LZiRab2FWhoGG
y7Oa72LkXDUhCAOybfVNyAzZX/QiuIxtZJtMNOYZJ35SHewMwqv5NHliswa2JSh8
8tHj+HgkuGaJn2TFe4DcWikGmQrdzYsydxyuREYy4h/86GRknAjxnUtGGElrcXiz
X0ChhyM56+anLpwFdS0LSVasDXnzmKEDa+W7rEHkPq8cmMtwlqvIm5GCjgyMJNsU
JW9bxtsx+ChTuizvrF8W4TfhoCFYBlUV3NaXdQ5WjfK2/6fCNhCW5nF3xeLWidvR
XToJnKc3Z5VdDdQndKiztXd4UNyJo5qX1ITw1IkTTYUD8Wrf5byGxpfMl83RMPKy
tfrm+rfAXK8llhdhln5RbiSiYrw0fv2s9ucLuZFthFF9LUXMVBepcxhE/THzibLE
sB/+rMDPKj9MVjrSZeO1jYXhmK8wWnvtdA0JAZCVrfw=
`protect END_PROTECTED
