`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+aWlE3eZqH6NOrvf1yOm1Is4BKVr2OP02wyj/coPDGA8ZwHA4sOKiU+4gUqGcoO
JJkA74vL1xs/teDegX0VG2d6LcoBFjjGVhW4LgMTh8Qlvwu7fVfJUW5Egh/TVmly
3/gjlJ3vA8B/VZKm2sV4wFo2i/uFaHqHZrRdymT0XG+MU6DT+hvlYYVHmkMtX6IP
vpfMugjvhX+AqYUh6mojFoCj/CKh0VxuADCet27eMSrlK0BCYgA0Kf6bYo8yE4Dz
QVkBwIlRNlNY3lkAj8jkmPR2fFlgrZXS/vVdG51epD3r7H/wjEXF7dsFnkEcQIY2
3faWD2d+Qu2a9VvpyhjF+o9/RO00rfC9pGePk1xcgwKcKQbyWQUZqZadUHOK12SH
fP2uoHKRx5tMcmumuLxrCYTArOY9vrniNKg8EDe4JhvbZCczzWSqqV9DUeFPTk1n
w9fEyowbNvMgg8kSYbHcbV2ZsEi4OS74d/XDfg6v0Yg=
`protect END_PROTECTED
