`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNyeCirOqXixQe34ecddxDyr8NkV1NE3dyR35k5JZfiFPO/Wm/KePrFOzd5PwQxt
E8rZv+REmGOuy9PxCZdLtnCPwnxf2aKXFcerG11TI7SMq4nF42mQfYzMuvxPJKyJ
JlwtJUfSBWNUPIF7YVNUqkjztxfBhRoLd95Lwp1q5WkWR/0uAdQKJ1vozWFPS7vi
6FSNEgehw7KgApw4r9GP28jHA08ghCjjw79gRqUlZy4AY7+T1DpXIxyOUwL/PWZn
KOmjKCxPtiDVHQ5Ev9utgZcNT4V+fAg3KbMf3WTptRmNfrAL/1ZS+ZyxprSHrEHh
1oYMBFt+OFCXIt70lQcsI4EXdTBvqcVIFmdPZ3NOX6ADyqAywWuzwzZLfTZ+5QEy
ooDEqcxUmCS0UlaW2wkhiwz3F5PHxWA55Iq4b8vor5dfUNXPuboltL4G0q2VkNcK
6Sr/8ktY/y7IufG4wyZil1yaGWYap1liUG9TfPqlHFABpqxfydYMqGqR2Y5T1ltc
XURuIu1PbjQ41iiGSD0Jig==
`protect END_PROTECTED
