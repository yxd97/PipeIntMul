`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISqZDg25AVa+VGQ/VNdw5WgUBGnp1j2JEYTyTqwxVBBL9Hk+PMPmoPVrcAgHX8v2
ZZ3ZrCDayGyGlqr6/um5tXfJfmoZHpOCXzoC4rpfYjsC50GREbWt9XCRetXOXj8b
SRmApIaoNSIR45HDtEqOSr4HGA4+RwEyw7G6yyXZueMnE2LSMtM6GWGlCBmlocvW
D+F7lDFt4yW2hwy33A3pKiSY5GeOw+MfqwqDqigFTsA2J7+tnrUZDa8PcSiYwH3o
D8xnxyW0SI08UD+Y5ZQHuhO4OLkzguRwrZzuvcST4VBr24WqaKq0UImckKi2WTjP
kvEKnD0tj8RegqQXBM+DqXPSuyUcQEhSt95ldS5u3yGbCQHqfFYee5z47Updt9ek
ovzRNg3ItJMgVrITxNP0CQx8h3i4H/o/9utvufXx2Jcx7PcaER3Cv86o4F3BS37f
ZYz8rF6ap5+Z+5nfgl8Y84f9CKVp2zULMO2N9utH4YvU5tPdQp7Nkv7cp8ttX+US
`protect END_PROTECTED
