`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIqjvBKvOfgQtcRmel/HrqKDYTlu3wPhu7v2vU963mC1dqdlJ9uNYCRSuL0OOy75
62+3wworzvcp/Npqe8YpT0LMuKYDCKVWIepK3nJkv+5Jva6eo891O/1YFdAoIyC4
AxmgHSsmgtHNGMY+H8PrMthsiFJKv/DLnLk8cJxE6kVTk8rafidHUqaqwk3qmobN
1Hv/c7bPWa8R597sxSigZsl+xS7Ra5IWkpFooC/RHTuiH+HPEzUmYiV3e8WzwtsU
teLfUd8S4Jjxolu9m5l6vS7zzHoboFxfT3T5fFX6dTxhdbwvG2xJ/RZam1LRKZq/
72LU3E5kyHKFzO3Ox8SIIn5QXNzWcnm7dRqtkqvgYlLCIU0BcHlm8QrJ/n04B5sy
C1YldEl1BczzYn7zu5GSWQYD5T+ZkPOfP617JGq2v4UrS2GjegdQ4TNXLiTos6Tb
/KC125X9n5sV8CA+XIzrKa7RhATP48jD63OsA4hf3GocYWUhOFU7AYuYYS8y5d3j
C3pNEONWjs4KQJgrGo4FyZtPaAFqdnfNfQzjrAHMuPyTk0BcH0S+UgcSZvins3fh
77Db9Bb2QZWRY+awy+U+fxNm0+3ZnwdgGEZUHS8p0E/1/gGUPjWccHce61IF1Bee
//XQkODLDcqOC3278b6pMrkOHEiubGL6wX/Q9oMjmRnxJEB+QdnUNVphoVT9Mmiy
twRuX1FYpqda3bs3QOZu5Q==
`protect END_PROTECTED
