`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7/KNc5G9hXUvml1Y2Q9dNWULV4B+jaYyUBQ7L5OygGj/cTByPaztJFLnknGx0jl
MD7dyjmYB2fO8G07og9FJr3z7OCOqoPkkapBjPiVAAF/OrSxejnZciqevGw3+2rB
4UU/HHNSoV9IyxXkbOU3RtMgbZbxCqn+/GeH6TQEhQecVvUkdwHj+3ng5u9bPr1y
wTkdcAddMRHZYHenZZL61SW18gtrc0A/QbCXQYg3ucpu1AVTAfnLKQeLtVQbJOXD
H0Rk/g+72Z99jIHlwe4vx7h963DQ8HwG3FiniqImotYqiwgrsk523gjDZwZee17W
IyggZ6Nb1w7S2ysKzbMK8k2WCfg2Tzd+wdwsXltIjw2d/zpow2yWxe1GcLZ+eKFB
y0bVh85VKc27VqypyxHKPDi7XoGZB7yY6veB7yOkRWHt2IEqtlYHhaFsaj3OPhzq
ok6HJLFVpvZuteR+nqzxTKOmftT/Hp351DtoDzbpS1DmAO8j0D9RNTzJ+Lc1aJiu
0SyqDfctJac2bivIZiGUauI9KVT5O1sxchi5XqMxTiVDF5Dpkg432eTW3EahP+pK
wrb+LxdHHWMzpmXqRB43uI9ItK5Tu1c5cKt7m7FnYXoYvkWGKkD97nCCN/g8+DDr
d2MVTZxBDOTUxAMW17fgcA==
`protect END_PROTECTED
