`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USevLBeEstmcTP0JkY2RU+CgnjdzhCkejNTjef48AvFubd+4GlnRTKV60Zgdjnru
oe1q2kgKstWHDYmzBU/Rlrtg7FBwNDYUyox3gVfIiQdfTJ89HSj3MzlCino3p92/
WTDLMAlNZs2HgBr4ItcN6tVzbGJAZFgwwFvaKOL2dgB4mUcd5Z9ORgDYUG/pIag1
ZDtKxwwaReNrrt5eYCo2A7Pnhag20s6RIZ1ysk3/DKS69kvrCMsNOL4YjnwNo8nd
Qy2ShmGwC6b23i/6yG0lbdjVNc5VVYonXz7EVluigrM0g1O3KD/sPmDqfDaTwkbr
PQFhCNGKmPrMcZEZPwTqiI4SFcqrh/Q5m5csmzpgotEsu1cjdwX4f2Z9KM4K77Pz
0+jfbejmMWX2Cwm8SYSRqK4ha1nv6sJE3XgVG4izU1sPReuet2WTAG2GUxn3n90a
LfnN9AwwMA5ccfoBRYl2RDqwKiQtfqQyIJ+8tXRa3ZoV4ncEwkbvVo98ACXpYswc
`protect END_PROTECTED
