`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAlQbcUrsPtncCPpFcEo7dqAagCCTDh2zMMc5NGYQz8+KZcWZNtKvhm4kTyk6dDz
QTvmkWMJVNLoRdXYmu967bG6XOhLGIXzLMjKEjEQ7qEkJelsXRt0PRPPrDCt7pDY
/hdZCDAXdQr46G0gP4thYpKgOqcrSDEkDMgV0AdNZWK1UULO7LElbXuVrEezrgAJ
R4PLtKniV18cHOve+/Q61P6tfrgHBgsIlupdp/APMT7eMyiDmOV8ZuzkailqZa0o
CXfv3HBAzMQOyNuDJJRItx7x5aKH63VsDyc4mdUlPY18lydoelmhgMLgzR0AYdrd
WsH1wzgjV37vh3PyMSsTmE4xMPTJnrcH5vVOYcBiSZFv7S9DWHaT/GpCwSVm4ZiH
dF8uJ0gGcKQMOKnAJqF3KORRxVWbYv3GNhOy/OHJHtwyjj4Rj6JdP6lJnHw/w7+4
8iVfY8+4KX5/CnyNuItF3aW/C0imymCAKG2MCkStxkb/bhjmJMYm1HaqYqkwQy53
vWjJPtvE/kX0S1kbH3wvPyPdhPgCsm7HVmUiQ9+7TgTib3ZOGCv+vKS6teAW9G5k
UUTB3zLuXYXeUiPhLtLrC1ApoNz+6rMTI6cc4l1UdRhfiqOORkuS3rYLTsJQ1Mew
Cva4VNvMkeQZ7lOjxWS7BTEX5/BBct/QmsZJnrGS7UjV8fRWcgYCKasgDvR6K/Hi
OvLNVgbS0ab9TENRMLlXGyocRdfU5olF+wWboT59n6zJK3AoN6DlEhl/CosO1OCd
Mjgr+OxN4iV8NGdG71mifxlxcCXeYUpsEqHTBLcRhwgwrjAOs38FuIdag2v1yac+
I/v0qtLVr+DR8f2B5ZGcCBwHw5o6rhJ5enwrHXQ0VNxNzes2Yv+aIfkhKjLsmZC1
VjXz4QLHOBG786FYRBae+94+RCZHiXDba5+smHQwVhMdPAq+f0D6V78MhY8YTTlK
FBZO/h1p82AvsTfq4W1gJh8vFPiDUPrgQQydn1RX3XyFYR28sctlNlbI1AeKWhH7
L+ufa18A55WVW9H1rB74rg==
`protect END_PROTECTED
