`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzPTQ/r66X0snmPlcXV6K9/Q9rLiVCxWznt4urlcx2vqyKjsHcLrhjBIV3PqkhUp
G3+SacCefYQ8euXInAbXfTfdxSsolmauXpqGBd8KBohrm/vbh50hZQSh+Wmw6dS7
gF4LQfUXrVq/bisLYdQSN4r6KvIoELT5MKFmVtRKGEx3QPIQM81wSkQNIpySHrqa
6y9H5Q5J5gAXN5uSMlu3sNK1GQ8fi9PiDgEOC9HjRVOLpgLTwT+SDc6Gnc2YZ+u7
nBVU5M2c69lv27paAVi4x2xKzoYvMwkA5IoPtm3rVlnyU/H8sTfOYHxUAdvamqyU
dLQOhEMz36yKgfnPW3p06g==
`protect END_PROTECTED
