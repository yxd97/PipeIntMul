`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44HaGyCgoNQGIJaASj1FZLS/tU0dEhU5jKglHb6ddOrYGqox+jNsDp1nN+R6MwOJ
tJrxZS9WVt/E7otmJBIq5UkYNpwRy7zYNHB29C4KuckNaTr0AIMG+H5Jak3TMq4x
eKLe9BbrA0tIZk1qK9TzBkdtMPZVwAHi4wOUW6B0Q/tmZ3GgDcLOWcBuXHEX+rzm
NjL2cXfPC0zgkHQ9fCitMgJI7qj8wrvnN9XG9Tv5ML3XZySwVaODfGItvRmlQari
rd3m/0OTUdNaqoO6NWgb6dwYPoBMKtqOlJ/PA1j9uf0wUm68HfqkxSa2Rta8i8to
G9iajSDil08GkbPxfxRJOkjvG1Iqth5QSd2GRPTKBnA=
`protect END_PROTECTED
