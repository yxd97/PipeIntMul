`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Beqwgj3jzSYF/1QLZmeFL6DwSk3nsfoXtDbo7eobkTpbALojPzRSGHwdiT1DeNxG
WIMl3T4yAkyA5gm5TcY4Q9McBl8O04Qgz4PrkNJKjg7jhUmtMDGKwpNrqVtofy0g
YuqrrIb2Ow4vKCk8ru2rrMxSkLixJRiPJe9CsLkBc7Ie3hIre0VbPB8sQ9aSfYuL
qMdJZaEnWXCRpZ6mtNO7/mYTAgGwz7raSK/zSi7nnlR+QGZizBe/9//2HtkOA8ds
zhbx3Ul0+ox4lvO2KPYoYxJvek398Vn/GMlBAnCiNy9tlxJVjcE4yfLjBdw+H39T
kDcbcXyJFRT4FkwFv8UZ86JVzF8cOwydqMguS/EuoCbeN5HKrK0m64gkCClOWfAb
FW32z3h9tbEy02OSvNdZiXA9sdeX6Z1e1s12LipRJvgFHOEzrdb6WMAw89NBMelb
p647Aav8ffSsS2dSHh0ROml6dGIlYfGsuDo9WMSWXBU=
`protect END_PROTECTED
