`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt8SzRZ18rUX+GXf53nr+JqZ6k2Ns8tnMdSro4+pbaiwJkMXQk68LdbzxAp9nyxT
tBWyIQBgLafzjZslVSbAXo6qaopJfxPtHf4v/ARqkGNhaHYeIxM4jheUl4f0hKiI
sH5PG4CfMTgCZLSAnKkVR6GizqBTLRw7v2Di1etOoYrX3AQcl6eNbj8o6146u/6u
Uo9aKyM4M95LaSqXwl7ZQjmUGP3h15N6gyRoJJP5ubzmPwiSYUEbwJGvrGuObTCj
LikorfPgseHAtxGA1+O8aiHbnzDuzEcsiWa9K/1BDB7s/5CGAqV3lp2GKK15KWGo
q0Al1uNTvJ942/ORSo5QjkDMa2DSvPHoMrAf47ieLrMpnGrVGc2ZHCzKIm59GyY1
fQNWwFaqwPFDTrN9xvqjmGGoijH/qzu/UioMNZeEIldvVxkeBlVVreJGB/fTXsKf
7ixmrOyd4iM3muUQ8xcDmbBJq/YMGqKpT946ZOs0B9iEolIq6JGNZ2lujG4dG/Qo
j+V+Sqtb2CNpLTyHwTj8RW/PjDtBi5zf7RxiB+DksnLKA56VfzaZ5s9+PIdGfAA2
to9zClGEsLcRkIM20f/R0dHHwYf2Z0hE4m32XXnhz9Msze/O6nyo07dvrepBq/gQ
QGWCsyLJDLaPl2BuabCmoSL8daZs+4Pr11frnHgQVuxAXAGzkx1FzfkwFHZpEOML
4dcyO6enWZQgT8VH8pNBiLAPagFMaqYBGJRPpa3+IsiGIL5gRDx2wTFT43kkOrWY
Lk0l8wE6X5ih3cKCqANNuSQJOg6uFrpSFTEc2bBDeKEVWZlpRr/VnRi39pIlT29Y
miyWreFwBrnCPxQeMa3V1dRn/F4ci9yZwg91zbA/NKqiukGJJNkRdYDr/7NgNV9D
zo1WhP005put13o/mZ49v6vsC4Hzd1sL40VnUO8lFxyR3Q21aJloRNv8BJW7YEmK
XouIg8/1xyoONbe6u0D6Erzt1rH1Lgeu7kp/YRLl52KSs3NUYc+DFGpgI/aTeuGL
dQz3h2UFszECYNOiU2KzvNeW8U/R8YKQtlgQRj1UYVRdFAqUp9bGcHiUeP5r4WAi
4spEvFgtV2IqohyjvotNBb+U287o3ZFSJRf9L3PCfK8=
`protect END_PROTECTED
