`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrj5zU5MRL443S1Pr1Zfbllx3zEwIQtNIyjcUMGzHzQvx+UCwD+8tHNgLt2CH0rn
MJLv9CtnPRrhVVx7hLXquSKgoDAOZ7B0iq0O/yMZyUevZ0GqdUadhuk/ElSVqFgP
HBPSiLixyW1aw9KqnvhZTupnWbq8BURYI0va3QA7jt2mC+RkoZQ9ZS0Echrv+NNM
vNt/kE3Y5Dhtmg0zOjV8ZvxortzSpDoJJrdyLbiQtq3WpGPVtcbmzGK2iTDF49xq
Fc4St+yW6TIOlOAg47EkvCkqKlHVT/bHP+fsQQ3HgnML3qbU1E0iyA9jfL4TU/Oh
j497ZjuZe4mJHlTGFVJrUjz9GHIoa4KgjUq0Jbr3iwc4cqvGQh9FS31iadex2IEu
+kuqwQTVpMEAIHxhLOv05B3DrGOVz578GyVrnimYlIrDLAZCTN24GmBMrAZea9bK
Pg6nlEvuUtNjNsiKhZFhmBd/nXi+AXbCYZa8NnDuKyIIRWuqzT1IR0cScz2uuoJc
179nKTw9muls44IW0ijIdnLJ2GZW7ayx0d9ZgK03w84CemJ59TODjBxXkbKxzUSK
SxTRP7PDC/oGH0eBfMOXE0Uoan6mop0uTckkwwUH/yMMo8mVSFf5mghaB/gbeF58
jotr4u6NPBTc5xij+23QDDSBmrQdDQbMfh3wCWg/Mdh1nNs5C3vW9lq414lPzOnj
LO+i17NuXYy0lugIsm5AUQZHLefTUQnKIeV3iZeS63XqhmcN+DIS20oWUXv24au7
yHH9Tk13QOWrLJUIi7wvrOyLCyq3sIDAjgUdySBl1L2OJCUx39FfhwMvdnZbUf4y
XmVUUOduCl3kTuLohh0XV+6htw6hipaQzeBFtl6yUriEIBEEiWYiLwLjSFW/n2ZE
2Sr6n8oiroDRPdhlEcnwO0lYZFHElVfCeZd6oMH248egwAW0LTA8p9HXkfvW5TWK
s8pMd5Py4BFR1+5cyv+eiepxPGmTyOYabiuc6hago8JVms7Krl1F9/zkU3RB5b8g
TE43OPMiLJeo042JXqFicuLojIb3lPtZ9E9E9Zalo8l4MblPqo6c8xSJLJMzCtGX
`protect END_PROTECTED
