`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2cx1TeoOFI93TPmwsbl/Wui8VxQ+P2YF0LgpF6jVTkOCeQ71TLsGatQ8ScrHGlWs
EolsDZt4dqxU+51DB72t7pv5gWJxdlFOqrwcjd99YvFIdEmd/p7m7i3S70vcgQhO
pyTruC/EGDjMscqU/m68XbAbFQhwgvbe62wKQwd0fAeCW8g+0unxyrmZ3kEFNlSN
8J7Yhad+jI3jak+pWfJ61g5qolbYcYAVeKPR0mzOR9YSpof8dw19i/lF/rZNSNmH
HCJZdCsIKnLeJODsCl1a+K4ZyO1GhMJb/Ke426nIlKNlvXVb8tbGS7exxQdCBB5+
8/Fm/HUuDwfXSXGZ0U55zw11r9eWn5eFs5Xf/Kx5nNJPCp9tD9m/2z9RQHpGAQvi
`protect END_PROTECTED
