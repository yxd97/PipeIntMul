`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJspuBckWgCneJZopL3sZ60NaOZJPFKQ4nu2uVi3e5AzEobZI8g4xVIzhIhgcXs9
ziKpbBiJWfKs65nubhzUZoutFaeLOr+IBbcga2DvAcGjw1HHgMfM0grnJ+2NWhUf
Iq0diKb4JPceDIyqilOthC0hKM9jaXDBHDLBgGx+vEwBVXOCEjpvllHFc8zFT6cT
YCsv/RO5ziljhXS7n3eXNTJAcNGnKeGz/XzAXi2+2/m1we66rXWVpZ5ZIXwuJ/j1
DKjAB+LhoL44et9QVz5XfdvpsbcruN1aU2BxtbV6PTN4HeSx23CT6VCdVMfJ8+aq
yXjskGbp8nrCd8SUjni9c/JaKagtqYGli+uDOKFTCVCQ5AbOR7puiXmzPUM/Nhm8
BrdJIOlbfCV6e8rRLdbzVRrjuaRBIuN94iRV05LtO5u0JFzg0WeuKupcQOU8uu6n
Vr9CHeyRVrZj/ous1L1FtA==
`protect END_PROTECTED
