`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66b42rIqT2pxUFCMK4Bmm/MRfQZMabLSgC2A1LL3n7ZUywEmhK5diEiLYjeNm6Ms
jkQiVwDga/vOGtUychGAWLUuHnyK2WMvSZuaYVKuKXU1TTgg/ePcLGhqq2oVYAap
r8p/MXeG7WJoHGP9a7BHASpmvX8mMBRh0b6bBJ9CWoecZqC6NDRro4yaYHjOXfwv
8y90WTdCp/K/Ni7IAGk2jeJhi3vpL3qwSlMDkH5ML6+DcdFJFavurGl5QE1kCDXx
k9kTATk1SRtqgNblWwnE+w==
`protect END_PROTECTED
