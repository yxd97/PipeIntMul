`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gL7dUdGp8LjM41P/Yzh9MIvkc59j9h6I0uCz8Tzn0p+uLi46qH+MH37e2FI39NEp
0M8AFMiVJx2YMkc8AuiQtArMc1AtVLShh+zaq9zj0H9LrKumkXwEOkTQd6j1Idv4
PAY/B4CyIF4whSEPAxSB7e6F88b+SxWnRa/mQpE7oZkkhCpjWwGKm/viI3KF2pvw
xyBesrZ/+VGVn0Q2rXXwszQ02tWCCYbXTTFaIpsTGPY9ldtTVYccNXQtcVyFnz4Y
ljcozW6WV/Xb6Y1aJKS8E5bunBdtDeL5OnLlkeE1s5BX1gTIXUcVNGysqc7MwJjP
uvma4GLkoZVkDZMehRjKI8DMdFz6lepvZHxnInr+HkbRvlEUr1u87S/Q5EjSHL4i
8RUig6sNnPWGYPm0P56Go78vkFdibGbd9adWA3bXFq7HOTt2oXZN210YBqZ7j7iH
VPPdM0sDLjjGqjTQ4TYRYlH+KV+z+QQa0trPMO4whSIhHQb2HPZcKpN4DilPUXXi
c9EZik/4XZx1BxiMAy350oapTa+a7d9GPNqVynZNhY8=
`protect END_PROTECTED
