`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+As3pmJmcnAxZSZi8M/9inue3O31bVIAZLgx6r5H/7DwLtl+0lnM+8M318p3BrjM
98uCbp7asoxzcnZKnkIf45lCHGoDJyQKQe8GjGuyNX4v0UrJbA5Thg0E+NQ2TB9h
De2m2zVEKty3/fl6gHfgXVxN2kSE7G0QLUa8tDakZ77B8TtB/ECUaFnk11TWD+jq
WvXDMp6Vv+hxZF4sjQDZTOG5p4PzHWdqmxsHG2V1havOGRMBOZEfVZX1JbFa6fEs
YAdGz0bsWy2+SPFUCAJutfFSlcd3WMhyLWrw6AzTWYA/VCxYpRNy5H9EhLc4+ge4
u2qFGAXKEjKhOWA87AGrjJ23DmliMeqnfCAzfyKInJvpfGwXy3M8F+GOJaEFE6r5
zqQhTYfjWDVsu7G5/Zrvxs7dyKG2k34IBbFiPqmXe3RheW+qmwILn/FG0QBJ+zwO
DQmiyDY7OpD+M6XmfaV3MwNqLi79fJCt2H0psHJhLd22eEnYwDbFyrkNxSLFumcd
vxHMNgbxhI2AUfgEZktq7xThsOB8Q7AtGcog6QpwsU6DNv+hq1PfPOTOWTs1KKoP
tAkDcRDYP0nAfeO+qmgZ5uS+liz0d9R+6j/Fp8K0jRKDzcj1tmG1+NrnzeGQdGA1
JrWNASd8jgetULHzlhgrpFBoFzer32IJKKq3VdcSGFeiEAxTySo+iq7oY18/dytG
Tw9Or2v4+q9hMwMNebgZzqJAjj9gjQnHhLuS+a5UileqVIpFTMbgWX7hpl4S6PLZ
hkio7eARiaEmZXbkmQCtGfomgsZwgd2kiD1rmrVsbvApLok/TFWa37GydOPlE9kI
c6+FTQpyWkpD04Aml3AtVtequvryW9RgpGAmD2ACGQ99az9ovIxMdcpmQcTTOFJi
vRdtR3c9kU2QOjoE2WCLAZEKNfZieyvazlnTD+lSEX91HrZBhMlzGyS08omsxwQ+
ECDtCAh48eqCzm+IaL9m0vb8a+gq32EjVMVkC6XcQmKGT+PFRAp8jjywpNvYqTAR
Mnya1LoIOsR5IsmuV0L80vDu94IqAyc+jMd6osooSKWtRufhyntulAG2QK326x8Y
13XpD0ozQIydM9+z0zax4gRtWf5WvReIO1JpBQ7y05T1y9A1Wd34p+N6LTBKBIHj
Qk41wfeM953NtHWg7dBZiHVQICq8Oi7UYTWDniT4tVS2rCZPwY3AAB07fzXvkidU
RKv33CeGX5K9k70dHaNBDicjPFoEXNTeangxz7aYKOzZY6f0CCA7lfabs73qVXj1
M+QshkR4CsFAW8PwcJ5qw+e6VwX9BH1NJa3w8nByZuLJEh5T9y7Z7n/uWZz+6JPV
NOl3hrQWBJu0kfjBo2at0A==
`protect END_PROTECTED
