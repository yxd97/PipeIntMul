`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dngroHHb+km8SV/1o1PIKsMB5Dl2IzNLP3iooPOA78/3Md52/8OzDp0nrayhxN5U
Fe5ujSeundMsTPwFs8soTtPToLj8lAnR1dbRZGDUBb50Te8BdBXXN/POrDWX/DdY
sXALxr0a/C4N7TMazCvMeNiPi1eiEILbwNXSKj0353b5Zxocv3p02osc6YX3gt20
H1uB4Tyr1g5hWjp4qZ+OIJXsIW6K1LrmZRQoKr600oLmKXAVJtb0qrHJFqcT/iH5
Dad4PbEyBqPMzkwU+1cm+z+yqMFffwt+ttDtOI20M/0+jg7FRD6sluDU0hoO6/d7
wb5hXEQZqgsSoXj184jAwAE1Dxgx7lDHfpSy6ckY0DmqqngOyAjohGillkIbuPUU
rFkK1VhQcL6JDPOWvjugTjlkp/snjN0A0xEF/3c1Rhw1eNdc8D0mMDPtAyrZ3tH4
pofbKIy6n/MwAvvDxTZMIN1Zw3IPDhKCa01FpzKOd7kMG4UBWNWH9C7iAdFondJz
+mb/JQHI7sbGYsgfleQBJCjI/oafFnh3FIX3kxNbn8mfgI/MYrVoeHogVwNKxMiB
rxAesaqNSu/J/WgMlZLu/Y3c/Dfl/+H1M4Bii9RX58Ti3XufmDfZEi0O51mIgyRM
fi3t7+q2YKWHlUpfLdjwa1Jh9+8AoQfk+gXWrq/WTiOlJ8UAEymUGzexaun8bHkv
fMxKTZrQoU/HxoXMnPNoDE7ePHIS5kcqEFNTHGrR0gsGxbVrhDNYHW84jf2O4kzR
JFgnvGvI/jM6m+kMoJ5idg4lGL5V7G53GJlOG8bcjgJC2Hf7GSvNMobhb3NF1rmk
QSKauQFlFQXbGTETrZotP3yZmAIMRTtdYNPFl2LbdRcifoWfwyOgARtHl7de/Rl/
NMWQStJ0UwAJKttzY8i18wVeI4Xn1HsN2u2p+rljIm37VgqtIpBFUVqYpSbhyRfO
BXgkyRPwTwC6r6Wixoz7bA==
`protect END_PROTECTED
