`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vm7nMOuGyIhGlmxds90hRJiPf7bJW98zLhJv9o7u26nxAteKh4dGmA6A0Vv2KfMM
5b94kIJijqS/hljNUfCZS43uPDFrYhIPdg0v5l3Vzm95YNr2S6hOxndycGw8yp8S
Ut64P9OG/qH4slCXbUJBG9geZv22D9PSObbxUI/uM1jhAbWuazOZ0gmhjzjbZug/
+aOgsp1+/dDPvpocLpImwpyJ41IQFz0Ue5xIWp3v3C49UI8So0zWwOrdiii2O9mo
NGtajyyHGVN2DoaFh9PPUwfQNBHNCCw+QDq+i+u7HhUwXFp0Y/v9M/gKMDPS5FRj
llsyBRwQx0VIwP0gQ+FFnG86WI76ijg9wqinKgUnO/yPnB0SEKTEUsm2OCI1f5JN
K5tCXVN9s4YxzRzXW5HggyL6c97tlKubbUnP2SqeQbJSasb3kRfcRbiaGjSVsyty
W+f4ma2hFgExY22yJVGNaRQo+q0afZciF7k5pDDciABhsppNxzjqf/ZIVfqk/6q9
ldkqAaaRtxReb6BqJetxpkE6tZ64RSVZff3u1g4NyIQ=
`protect END_PROTECTED
