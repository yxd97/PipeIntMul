`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aoJ7rydUewLp+3WeM+ycOjIMZfmBWhc5BZkrH3bcfkk33UgaH04vFvxeQ1VywunA
6W4U97NtyGKtYPPumz0HOQ+DUFc2Ns+5umeIVDJMSL7izsW5V43ANeR9wQbU84vY
Dp+2EDFEPDYV2/hfZ95atx33XKN1uINjTEp+YVkB0gjR5TtQGANfKz97RJV/rEqu
VuvUitEVr1l2rC+Pppa4nsGTMnLZZJ2iSgAC5D3gBcqZd2KH20+MdLsr248QeBtx
aRkVkyg3vAuKhxVJB6n4wMnAKgTJ2Ndpv38QVaXLqUeoJjmZOkGP/kM4eYbiE+/h
BR1w0Jei3g9864k8A3g0ue++TrwEGZKAbRxbeGn8lgoTmc9UfmzGwdqw2awPMial
CT8r2frFofAekpgr1MkcE2Rr4ToEztgTy10/K+xFiC1Lt6Rs1MHmlbnxiEV/TgJJ
Z96hveujCSGsZIUHSkcuDPu7uTQ1I5J4xqQ+WihIRYwzjO7YI5b9UdwcQxGpmGsE
iBl0Yp9Ws5wduTNIeHMQ46Nua4zEuhZlKTmILuR7G3AdnfyUolNaucZBFVmXl7xt
4mjGgHur1OA5QQR7jo82P+n9+ja7luJeIGFQ2XhiW8rwOfRwm6dBoEpPz7b0voLe
LlQ+z1D8SToTg2+Vktpo9R0efVTOLRDcrhSpmAR36kmNO3clLwEqZzYtdG/eatEF
dtTMuIwvYoLJifkP/+SW2eWTaodyzjPbzzxJVEsLNt9DZJ6C2scAcCE8juvLckEP
ZPhPM6xkSxVtLSZqqpj/uLRXLtO+riTJHz5WClCI4jwJew9f9kJT9FZkoF0Iz6IN
RDhD9dhXZMaDTYYCCC3m4H3Qa21IaoIoCXB4IIv5S2PNN5uf5/RHIZilpwnlF5mt
GOlWQfbx92xaROja5AaX8h4m4putHC0z7amHuxX9ff5UmMsjSS+OTdAhcM5RGTh6
`protect END_PROTECTED
