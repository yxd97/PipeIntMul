`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8jVMIyu62r7SyhGd8hzbj7xUCEP47+WfXLQ7fT+ySyGRf6+LuuDO7YdtxyhHvjG
8ps2NMQ/2Vl86ZIvQIwk/xItsm5SX/mAd3M3DF0iLh+LJgLirSw5urgVY+uTr6nk
LFJ+ZgUmqPRVlSR33nV2jkt3aDvC2TR5yfCqwYFeD6b1+dtAFbqNOXgLIuKWjkMp
qE0TwsAxeiYbTd86SPrbcU6DIxYTnj2e/fTeCQEHS5+VZkkxHdmhwOAy0S09YSPN
tg9u1KD/+9t7U60/frcWCmbcNuu/YPDzCqewJ8yecQnSJ9GtYF2Hrdvbt0d+1lEA
T8PVo7mTGsZo39wW06rUcAcDGV3Of3WvlsLGcLFmuNhLOXm8xy101w2ES2Hnrw0j
6fC/jRSWSEmkOAoQJxmf6pwduqou4Fbh63fxhgHfDWvkW6sZzcbI7wIwBJBgIfGV
MOL+xBF12T0QxQX/O3JN94g8nkf0pZQaUpsjaVwtzAX+DrxKtnJdR4WeQRvaK6qF
DxuHAMe5DfxDFr5Kia+/mwKsAAeZgYstml3U55hqRdUXUxv9UBpQSK8UG2u4pAmo
mZpw4UiVNXeZfDc0snORESvztPwD6/5+elewtFJXRLuVetPkBB913hCVTx1qf5Lq
1zXFP74wfl+2N3ZXLc6+gK7rcBdqFN4SMBI7ZGeM98IhXUfZIvYHlNYozjydoV5v
DSWxYBOlCc9FwKCQ3CJJS5Kt9rXKq0MiZknrXpxrBI7oamRMMy4kDInIVPbIjkhF
`protect END_PROTECTED
