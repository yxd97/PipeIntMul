`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LyafO8r35s5/OwUpKwDJhoECcIrUDB4+ggFpmpZlGdWIspoC/UE+8ZhZ40wxs3Cl
YPN/uOhXp39Vwf1J46PaUKUwoi43DG3Z3ojD3a6BfUNtTMxeVxGMgqr8BUbggjel
Ct1wkdBBIA/ZuR7hnX84SSkxcB7f3OvCfVILFi325cndA7db0XB7flofQB/WeKpy
QsszvnL0wAkNMpOzsjBOo20GUqUM+H0YB+EKSN28SXtuEAQToCXkPlTOH5yJw7tx
JWx5qT+uherlu5an2Yz1oYykBrb2xHOVWzDV2T8UbUVKttxIz87xVSx/m01xKs54
PPQICUa5BLqn3cvuKCH1smyU5xBeRkd/ROGt/Bu4D1EVmg0bzpZFUe96Up7pHpzg
+q3+NBvXqGOj8wDiXKCUPwbmmfnZPyxXsBvztXpR3qFcgBUPu86aFl6REd/WqYHN
ruqqpRTsqsHlAz/WmMuME1pR7yjg4IcsF+PpZWPwMWXB7liYyN2MP7EsUafVIjxN
pUu8KQdSHvzDQpn+6DyFAVBds3L9L5dpswo4CVOIOWTc9Ovo2FvyVdpetcFdZAOu
CxW8Vuo8hde+y4bH2bjWRy0mAc7YruUFN80HiJFXc7Grqzqxd3S0o3g2ElCuIefq
o75GEs0euM7qlJN1P8fUiFTks0f4buCfpu1sIXa4ynwjRcT12qD35IpDEhSbikiB
1S/UsN5w7SfOoMP41g1OCGZZhb8lWewj6zw6VwhT4fEbAZeDq8rWZ59wiQn5mMoa
OKYu3VTLZ2HlcqqrhgNNtX9lKdwuy2sWp7X7fCDkkrwKkuWWYmFQJj9kXJJxqxrm
cG9K2yyFAyzb2Sb8U99myz20ZFxtVOc2Ibr7hjRtS8YbpjQ8Etn1PvpqsFb3yzB7
jPMTxa/mdGIIo11onD3Z9z3++dxztj6nHUknX8jcE7NnzNqMUNgih9kn8iY+qOke
UsXpaKYpsMTKPoWYS8UKXITM2N6LG/8DR5WjcaOmvGdn7YUzlDTzQ0UqyCc0kvfX
kUZ7mUSTeAcc60ps6ND8tKz0EBsr46DD/FIkWiTS3Qfin6s6/22lU50tsZRsaTCy
k11p+GzlzGi2ibxM+vKETPGyiIGD6m5h5WsKk9rgO907QTX2ocm8zqhFerfn53/6
huntyU5bIN7FISw6Drs2ckLUHsMiRtC43VCEMSP9b7c2tYg9ZxijWeUYw7uLhL76
oEwn0Tp5WTq6F2uvYO79sZzzGoeWzZ6Lpo9l3W0By8+BxBFSggU1WTyisp2Zsz8n
WMAULMemgwhpEefpTUYXqUhgxfx1X/fh7gn/4q4GEZPiimbCYLr0CCbxrAnl+Qdc
Mzf5RZMZV8E9Za1+5GCpcQ6khFh2a6jdZm2MIy+pbCDh4ymMgS8QBM8F4VMFRgxr
rY1EwTnwLX4a2LYcROqqK+mHk6DDy9up7EZdMptFR1GH8xVow3LPVHOA7f7fy5zt
iuPMH5/7zRS2qOsyrF1t/giOSYWl3+uC1thV/OEIp6V3W8nsItrD+ScXJdCw6GA0
1oi4rHc2QFhwZJ8v808uwTo4Tabr0Ssn5DmNBKYCs6r8VyEUB20noBIeZJ0R0WZv
`protect END_PROTECTED
