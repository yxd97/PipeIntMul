`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HnhTMIGFM3MrnjcMW4d3QT3D4x7TKIXF91ltWpM9j28meq+83HFOqLHCPB7U9+Hf
MDTEAzk3Y7G3i9Vqh/ACvHPd/k8aWG+P58OZFiHHT7WKUbtAu19eplH7v6gDp6Aq
HIYeSw97+tXZ1RF9g+SI9fFPoOephhXUmd8zIKnu76YU3wxpf37MqOEpsK2GHs3c
gLHdQsSOtoiH4OIRVjo7RlZUF+WvWMZLfhONn/ccsjmgU1Sgjgx9W2Z8C7qrl/Mq
dRlE7asLq+vO7KbSlgBW1XYHXJYnlYyEOOkLPvFQkkhZZQK6BkunzvP2kBiHONwN
/eP0TbFwkFmyRpCeKEU1CGHVbeeItC64dUKyFkhLRjC47mxvY+cq9n+NCPjlnHaM
nd+98J6a6PelSUihKSpWQ9fSLiNEg/0Mc4I7UU1m42imK5ky1FQJo29eCFWKbx/r
iNpjcvkQwflIMlBSn6pFF9UyYGtzJNBrzlTXJnr++sFFYHb5SN8qdBqJ6hbBaVzg
E5lTpftXhnfmQ04OLn/gbFmFP0SPgAfpYUx0ob5zqTuiFew2Km/33R+anC1QpkBO
BGTNmKe61/Ty+KOkyEaJ7hF/1s+8KuBNKVRwpuprSm+PJBEzPbKTwUwJzwolZckb
Wm97SOdrzRtA2NhhIVk89YQCOMiieEBgk01+Gz+51PmgUD8XCrMQnvfc8acuXckA
an4MSc78tE9ZlRJLaawMfUuLewQ5I1uxrXLbdSmxvHclAF4+y4NL5QuFYjjKuDM+
ya2ge+pMufzsKqxhZuqyK1hDo1SgrAvILleFCKHBoY+Oq7ri82Z+Ts4r6QvySmgm
J8OnycMCqS52QzH+2Puq7+q6fS9VAXnkWy72Wq/chDJ2dwweZ/RB7Mv8avkH6Nw8
dLsJV8n7DrFtR5QgcgQi4UZAiUGBeOta6jB9gjIsE/lZOMnthS5lxWjEbAnLa9Tl
QAJO7+acQpnCg8sWLKBz2znuapZWEum8wAiDCmuHeOykQIKlPla8RsNHpGmZC/lb
5vDfwNoZSMCA/LI/USWe96nxOZOLc7wbjmfbMgvewN6lU5uJ8ou5uLPt+B6gxZXo
8WLuDk47eAuJSEkJsZcQrjnENYkjFSVcMqdMRqefuYDmfplqS/xam/r7px4s0Tx8
BxFEVpa05NjpkChOpW9tq56m8ANpIIcukzJAfGohqilV19rxEtrVT1cCXSWmshPF
sNq0d7ZMunNw5dI3i7tnT49MwBd192tq7DuRNlpon82iEdC+TX7buhmrBxkxG+e+
Bb0Od3h15LtRo/bPo5wB7P5zuFRaszRPp/ZrqLGOFr0XBU5JvpQJGE1eIsE6SqNw
YCYCTyfUjM9a7qdTfkNKJyca/7zB+fCvGrZ4+nVKgcqX3/QMcvy68f38mVBE+WHc
AU1kBfPuVpV3C++jh1NkrqNvXC5/ux3Mdvky2kfAvOaYUaadrFPPOxCZooqqcCHz
AykLf8k0aooP7jAg3/1xTrrHY8CHJ4nAz/jDsa7qUUk55LRmsXIrfrsosqvteocl
d+vrKVbB8ksMtljVUESrSpUAmjpPcPGQsQRx8LudjkAHqO9JLIL0OK6zSD8yjsj4
VMosonxzo2XuuloecokJ08VQhiOkJJ1ftnG4negeLH660gNOv92kooVAICMLeEHv
b/e+pQCfQMyxLoAE2nKClnf4d68gMcK5lXrVcUW7qRX9nfy97JT3KLGlOatfPne6
zPrzVyJi0JwVPf66dRb3o86vLRokSrAw+9I5xb+xdwQiMawN7Qwj+SqlofuDjKtZ
Y0fHWTNF56/wVB5SFoF0TqG11NiB69xMIQ3wxCvpaxdx34faRmeDXvuLwyzFWIFZ
9X9ZkeLIQl0qSVURASdHjHZ19bKcR0B88Iog89Wp72TyT+ayfIc8Pb+IKU3ytrb3
NagIfElVmBUoqft7//jUTTG/Fi3r3E418hAlakPLuRxYRwkOqZ/W1GYv1ywuGgQg
K2vAFcLUbw0eB1U50hN0H9H4q9PrXUdxMtMz6xgy4R6SRkPT03UloDVba7Qlg7F5
0wA6P6qArQ7I6G/QAVqk67lhboBsq2vyDZ/vflhqsImomkRFqqgxU50YizxzzVW4
giCIboAihRx1YbGUtFoX0IfFmWikVzXZu4hofd/NCrHmPa53gRF/CjEEp6mwe66W
Zm8DGcoMCR/KNOpt3Uopn5SSExtCH6ShLPeHTKiZeFJAaCN8ByT+Nb8gglg3yY2K
BYFNxsTtrm3ZR8/HZ+4r6/wv0Q0AYkBJvzg77+9HuhyiYnaLdL6QyaElA/P3xN1w
cMYDK06kXOJEUxDPcmALL+LxMIj+8VsbrvGhd+05WutgsxFAshzFus6ATD9cAFux
/Rl4mpB5Ady7POnaU9tvoz0sQRm3syDB5ams7k1/69t1/gKWoHu5ei5DwdOqN74c
i7CkUcvMXkYcWFwNr5NJSRY/ibq4cTJTEQYi0ExaWNMXKlD5MUgIz4HUIkkGS0NS
5UCwKRalmAvL8GE1J4QhkRuF3ENfkUwbICbnys7DLUS84PEgNmilxW2nzOaGsS9F
V/IeaD8wk3Qa5EzEWr+E3C34MUmFzJKL5HR76asFBn7CIRvuEfSNLaej4TSZRUji
Kn1eeGuh8jRnfyB7NxlgsWPt6b80OojSNUyB2oDm8g9p/OU3QwpxHS1Cjx/OUMBF
iMLwkdzGiO8VJuxym4ORWog6XNIxoo7NQ8rxU5zuZRdnsQBquvFCRT3YyEq3QZ+D
k+Er7AoK+jgLDgkgtiZ92g==
`protect END_PROTECTED
