`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E7xXQMjySsg0NBmHzscylzWE/HI+Zu1QEAo9IB7CNBBmTwx10sbrgrR3fkh+4bNj
wywc6HfIuBsAViPkxktVlP0PR4/SG9efaEdXa2pAalY+cURGoNykAQKmys5FHAq0
0AxKLjXBcCrccY3voD+P0aSigxKviZsAm3Pc3Ampa6rN9WrCPraXj1AbXyc1YMd5
NmalOWOlBEcT+/BOlx/glB+Kj1iDPAOU4LSjkPVwVDTP8OVJiwc+KHOc9y3ernaz
7LTjPvGjwCUN0h1pdIKBt1JJd1LmDWgqA1EgeD/GT8bHyenHF7+L1KysgSFsai0l
HwgXWJgacjDC2hfL+F2xrtqN3M6RPjnqfbU85aF/wf9SczFgvbL7ezaPeYHxc7TQ
o0+Wlrmt0Qg1MFy8ARu/EppSHgIfaJdCeGBkpFgoX/H2BkjdtBEGci2OiCR9vbGR
Iro+b2SQzCJVcvG7r2/vZUmHLiBQVX43JXvRvoG+Mh2jw1/NcsIKTFz3QSOQv9sa
U3xLJ/Lk6FF86sFM3iBI4i1TeEppe/hKjVlN+dicLXY4P/J4o3u1+wi2oIf9LX+I
JZF9yyu94c4RQz6sJktXUShtlSyCkOMQbMWOJF2n7fIkogJc5nk1L3YqNEoKUvEC
o8ftKZivEXavRgi6XyDpr2aDrvPeeV6G5GaRaYOXKkQrgMGf+1aT1cYUAuRJ3PkQ
S/P2+OQ2KYTpHWGFEhUeh1lD+mu78THM2bgaaDQAlkGQMircxGuSrr+ydH/3NIqE
+2tockOMwVbGmnuslBCfDAkFTJUgawGN7Ymslyk1tDzi7lok5nR5uIsBZ/bbLgYF
Xnsg/Zh0fxuQgvQNuarEnGPb6mt2IQ4jOkKRetc2uQGS2uKDhxjWGTBifPJ4ZaZy
DvaQPl/HxSq7Fgu02L07R7sjMsnA7m54cNmEXXHcMAltdr/KeLmqXmeO7cHwohHh
yFjm5DO1T+sz5F5s7g9q1HmtJ1/4YTbv8f7mvu/V8x7sbkjg0udjGLsi93Z+ujSB
uS167S7ddrvX4yTRpl1Xne+sshX1on8Cw8OSHTUYZIuLCmvAKArJ6UHB5svWYvLQ
z57j6Lx9fwegbPbCcjGryjgE1plCk3+T6LX1lyIM9z9KmTaT+i54N08LVtTh5X3W
owBBkE4ohQ01Z5i1AP0T+dbbzA4sI+axLoBgyVOqVThE7EkSubDEmQylMDf9N7+W
XFvQ32IeGdhwbh91lHaANrb+pOsL2KJYZATfYCuJbZvZMtf2YZ6Nu0TydD/pgeu2
Acuie/Mwdb13UEklPee19fRnjNTsMvD3Ujps9p8icYGUePkKwLInGo6TOC9yVRTC
AekwcIu9YqL3a8zmFleOLVCjFPIhr9Mv58ALlXSgxLeThqDi6QycJHUknYZ8jsVf
Va8hVhPP+P2GMYchVZO7yse8C5cVO6QP5e8Xr2FJxQqQ2oUd71gZq3teZmLNjfNS
`protect END_PROTECTED
