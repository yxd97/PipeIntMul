`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zgA+rHudN0A1mvKDW7/qIqjoKx5TDNN8rq/JCbtSE6i2s6sU9jQlh7/zRw+VkJ9d
YVzS8axTwI8xBfpHiN7VXrS5/mqW6VP+oeDJcQQ4LOyDyCLfFz5DvWWnVMUp84Dl
B8yf6wUyrIDGrh5h5W4cmPcK1ERJXgfrADvytwG6uEQqJzMu5bmjk9rQZoJ7MGaQ
mUjAs0NsQMZmvpKDYxh2q5Fbr1kgCq5E5DxM4fJJi3gPbV7oKHFMxEHXIH1wYoJY
ibKw+eYlrAHxtHfTs7o/EO29mKaPIYADqMgt6GBKtexp0y9xV27nr9VJAuwLl/Yh
T7esYBfxNqg3ZoYnb1akRg4LBulq9PBQvDeRKE9uFp6hjtF/u61iP/O8UKqYozNf
oz/mQjusAL/Rh83VO4iB4gZPA0zb2TkbeXO6TiRIqLqVTsycJh2toYpfq4Xde+IH
wyR6G1hw2PqDCGiqdm5toV3g7V7o+fS3UEvoxl+h6oihMQx4Y9C6WGi/NZVBlT0N
Cs4+AT7wmkfQzyOQAm3yAg7BzXa+jZMLTVZ3nWVsfHRDUhL1OdXntIDbwmiiLb51
dBke9+KnU/G4PMPrRmgsyrDhLJYc2uRuFg9u8bh+V3gvBJUsyv0hiHHinCApNIlA
QkRJQ6KfRQU98vCQUMKsH2GT7toO9AGAzK7ypUqQ3ohSPL8sjVSCFssUqegOd89x
lwe2wiaJvt2wfdXvbT/glU6jzrYg+tooEEeeDIkpaU9QFy+5zgPtlqEjceHt58D0
lCMOK9j5nKzvER6FiTuA7s1B/fmhEyfSQEVWRKBoTrideWitI9xB+DV//HhQdetJ
Xko4fqqotWR5k95g6E/ZpJ4rHbZnW5mJRPiC0EmeGZCRAcpBvdLedRKvxhVqPUUO
JBPl3Vr1PDJE1d3/dNgnx+RFaHwgwWS2lgC691j0SO7eVMOeRzWGlW8JfBC/CnOs
GxQDfr949Ext36O2Wgs4B6wIRPszpfmpFOJU2OVugBI43ZMD7dBUAQxa3XcigluB
EIgHAQs7vSC3KvkO4XXvkDCJkSFM7wcHuxN1t0SEkEuRCgGwdZUUn85+YGIkJhkP
xBamqQArc1byHS3gFuVMfta5+/dj+4f7P9SEb9SnIzqWOLqA9fHAmUqy42eimB+c
kyq2xIVKTueJdA+Dolqnr2TIAHPWr6NkWZHv5AcjoTouAR80fMyZ0fX4zaXN1eb0
F0ZTF11cFTohTQ83jBcdQem09mXaks9nNLoeORHtp7dY1nREu+qProYM2lqlJkrv
qTjP6Cl4A9IvyD2CkuwzLmpV5nq4Iier0A4OIXFBiiUUfnrH4pLZCPQLj+KmGlbe
NED4BJL++UG53+Bq4Mkv+F5lfXa6+ivJznxnFkQ8AEwlPoaSGa5cO+tQk7+pdSxX
jsSAIo4RhyYS0uev910cc5sDWZW3XLD2gj9bq9uz7UuusbExKj0eJzkgV3N7jgME
xie3BFpi3mYFyHnQ5jz7hn9Lt6d7T7mO6mVCmU9ooYohMkjfOuFuun7cQ9e6xmYD
3NmbM+4IxklTZWmEwWwdFQ2tZaeUTZ4GPNs55r022SVPSlT34oU30zn4TWSJomrr
8nFcEXrQsg7R2gZlvUYN72jMJQwJFl8cYlo0k2RvE+X55F5/zbPR90uWI+V8cl3j
hJf9KTqGX2GKo4qtxrSuaVxUdYwjLfpL6ph4O5itySkCO5+M4A6kr1veKlkK92kH
yWeYskECQ9NIPOe5FcZ5UC4jS4t3mmzIdpbdLG8Xn42s8UDgmVPCjfPt9QU6U+Gz
JtzvASuQ1Eo83HcS2DfgSDOMyTsTBu4QIX0SljB3y/QtaYpC11bPeF1RnC3DRtf1
2TT5yIxNzvqlFfvr+o7Hp/+umsUxz9HV/6xxuQcji04QrvJulMeCMuO5EpEdP37E
JODl03tCVvamerNqKm0jGgEqpjf0ZcVJBiJUwp36eX4gBWs7w4wGO4umLwwHNFlp
tSnGQAU7/kS0jOKKAp5OpdJR68nSdzl1+/vTbe1vdkZ0vL8kCJVnXflOEja7xOdj
4s6VEhUS4CCXgLVa5ys23A6kOHUCaAxcRv2sHTG+juZQa/SQUTXBovTQxF6BxTFg
UkyCOgOi2UekEHfK/CpKt8BLqZsPA5fpNFSx2BMqhCJLm+popY33mCPe7wSAJrdt
skdL590EALQdkfTkSLNLgBgTCF38N6YIYVHaqolpbT2AxJNb7oGCQcVmqLVuEQEb
QOVmEE57vcsiTA2y+KkYS4Mb/CUKncDk5M4Y7roCj+dJQQAa9hjI9i+XXsek4d4m
1FkUD4evlwEbBNMBZvWHNceutOx/LdNoK5jG3L/0BZ3lbMcMJh5i0327WVuPPXlm
GzsooYGVr4Cwc5RAUz/MTyvqjll1vC56bzGXS+G/H71hfIkY66gn8OxobcqMdftX
cFe8L7epGCN1Nm5uke8dKuJLyPpuVDOeYOcU3j3G8ojqyLHCRwCjIktsmJPjG/V2
sSMFRhtLCwQLgA6hnYg7WF5r8JIMxyZFcWixEBGwLfx6Pfqqcr4PiiCjRWbxUceI
M9QbRmLLUqYW/iupdyH3A3ByuUFHyZZFDdjS68ixeTUozwg4spZXv/1fz/WQi2Xr
HUxD4m5hj9pD2pzuw8oBVV52Xeq7kIu13Jb8xqIkxwBn5htnUHPVWcHz2ijnFZXR
E1FFUyuXQUwJmaQ3UUZUc6i2vNjohnA9TCzYQvuyboSV62r5/Hmn3RtJXq9B26Z2
7rmEDc9Hw8WDLTO10Js/dcSbdxRvTo5WE/s8vyBsR90AA8kpCe9HJJdpWlo6LLdB
MNMq9q6iFMAqbLXqDTNqptbmUlzsW4fPYieTRN1g66NO9LJdfK1jgdMST5IHV4Wg
Y4XKqN4+ee58oomH1uMPgFmfmTr9dp9in4fi7Ja6XSxo9im9Dfjwt2NmSgY8um3g
3uz3POfre0+G37Eoih/StsWGeNjA/22f8iHyYb4BPp2wvAkeg9KI6dXq9Hu5TI71
iXtkkwyMAP5WgnNfjvy68httc7Rnm3T2DaMGCAtrlJh//VGeKjc43g4QiVvF3296
SdStzJDsqiure+HhHLZTj1tgozUtbnxKOxjvV18Vad4Z5/1iYLwuLJfigROXe2il
pLmzpsK4XR45dc+7sAIS91TBLVmipU3T0KZFRQeiW77LEB4Wn6e9FLbD+1GOUN0R
3jfNaWTt1ZSMkC1WBJK6IdoHj4WpThTK3j1ZPN1mWwTopP0jhAAphWiyZ2Sj4zTo
KO9skbCiMWkA9ocKvJ/ZbJwc4rbU7HckRDAd/Qar/jBolvfdF7/T0MqWf13hRsE2
GYRKr8pceJKnjJZGUtMTV8ifJRunYfx+rIAh5oKPFu9u1WjbOyEVjG3/t8YvO329
9/pIyYCUWqZ7dsir3+y2LvKS8tnJZYMf0E8DwmBAxc8OHPwyEwSRUtzmg1YvHIXH
VlRAZ240wSb1aC6zsX9MPhFJl8WymRcpcazJM7d6fRShGGngfEC+mN9XP9lbT8Zz
jGiorCD2bq/UjyFUANNo8rZIVggIMIcau3nO1bn5op0Xb1TlHtcIIDnthhohqu1a
CjS48/q4QpfovsznrOjpkQgGhVxRORGol/VJsY8vKAmCsWORy1f/vRZImXCBXlo/
i7c6P3NTZFrlBXe7kKCXqPN6j3v3SbeJZU6IgZtnmm04U1Ual2ds4LVjiTYh85a5
HMX/savl5ewojeNo1zZeJSTpLBBYwQV3S+OUppyUJb2JeQVWky7xu8jT59EBcg6N
a3e7bm3a2hW8C6Ha7xdUcbRgtzcxNsvO8Dtxy/EY/rJdptOxY52CUKvSi+GkB8iw
z1YIwowrsZjtIwGAcGcNgJkS7PhIUcxm3rP4FICUgLNBcA6tGwXmaZH07SqUvlXu
mwe9LqcvSIWMqDd5McnNFPPvjccLgCAWJmBOnqJ6ei+1xJrpmrOfnJQjJdT8zaa+
QDKfwfCFqp5ChZOPL+EnKw3Wd4ALV/5OJQGvraxh+YbupJ5v+nSIDQ7ANQVds7a3
4zKLvG2IMpbtXEl+5Dn4fTxGoIe9WGEGO66FX7S3UlWmde6Wbeju6wg6dkZvyYti
1DJE32yrFsELOb6A+lmFDY++gLHrBvM3Am+LjkJBGjT2+oYzI+NHT223vOUZcmL4
miqVDYaBgozZIozuc8nE6VhF9tPyidUxWSy9nWSz6YeM5kHd5D75ELoJpian6MJ2
g+phK9FwIEWAszw7uYfiZ4mqGGj5kyd0qmmNwh59LukWSfutE8pRWMn/1QQB2Ubu
LCxa/eEXaNUste65AXJU4AyrchIAcMHcsMgm3Fo6BLafzorTFwbiDme2HQBrRaPq
IwBaZ2U5/eBD3cMmmh6RWCmDZFEULvlpZ12jLO05BmTYHCIaxyzrCUEAtqNfT1g4
CqkYAWCnDEfJX1/lUvfiMWVAB3yTH+yVWBTy5/jWkcr/btr1zQtcyNHzvYpDPqtQ
XbtrTDqnk8KKa18oh86sEI+vSleba5f9XPLpbUd4QvFDGclYazjYV1vlNNvjZO0y
T1cEcNqv0vsrTITijtivWZRm4Dp0SgYMgC5Po+ArRyCcj9+pFaG/gv3xIH+bRH1W
2V0Bby5xQ/T0ZikASk5byrBhvGrV7fr8YD/FyiHkztSqrb0gCuxdwNqErtuIGLS4
0m2ujghead+D+sc8LFxqaUH55V1Nx01A+FzIY9QJNOUc+eH9SH8Alosume3grZui
i2ROtl/lJvJbSeeOZa3xukEbH4WooMiqRWlBzAecalBmL3XJPL2chrYmuEP0uQg1
9pALQcNpmtIDa47tfCMy5dIHNV2c/3ojUB84ggaxm3knC592XPIv1SyfuPh07v5R
ZfI5JkGTQ5TaK/NAVgign51RAL4SCLWtAA/cbH3fHH71I0J4qwqCz4mhxteGkNSJ
TyUtvVrDU2AGo/nMNW5HC4mJ5DZCGYi8YB+JM4+DkYs7az4P13QN5cp2rpZrzpZ7
ZpmqtMgH3PDxA74jAA5bOW3+tLDbI2QODTfSaClRqZAW5w/YQ3xnfMX926YH00yZ
8MiHBDBS56JuZ05gnQSD2QdKnQAa5NyoGjMXbYXXgBuFGLqvaN/FVh3zhCZ7wBln
t+WJ52y3rUxT5xCkxoWIzvN/8L63LUQpBMPmjbP2eBIBNDGfSHJ7EXRP2mvrSEdq
AVfpiAHQQZdXAT46bLBkK8U8iQVbGQMFJhOFpEHUkRS2p17+CEYrEYI6jRBaZ20C
E4qTdAwaKQrKKfdPTynTgnwu0VJottIx+kwp4F+MdORfBIMqtTK7DNCnqWos1x5q
tUpghVeiTz3jQuy2VbbMF0jNvTzOLZR8q/x0vGIBofTNWOoJohs5bC8DP3qZFvcS
aAiTSJXTluc2Q2NMIBT/nR4mQbS1seeyNTP9U8gsOO4XafBHqvSN2LgL0eKVrpQi
c8VEjRlMTFMl3AGrJ0C5WH8XP6ROpwboFuk38p58KZXvPLDLNVOjQUhWuVINketz
4VXJpgxMv9oj6f+edmL8ZiErKsTqF3/FyAiQO7MqUlP5h1WY0m1Noc7+X4xaDtgy
4ljY/3N+vYP9DFFSVYIH1HYhAMLe0lpXaU5GxHf0Pza5NBnWTK3xoKBw5ChUnnVO
S07AAdt6BIuaDbX4gFR/AY6gA3neZZVlDjQpsaR/SzfQ29Q4fvShbjr94/YEoXP2
0x0o3wHYmyWTCCjWZByXsIu2F7IKY6VKox6bAe6WJZjr6R84ryZ2aLS1N6UMFtYo
yzzA/NrxbzmXYWC2wsJ8wCkuUkS+TeCkKQyrYJVq3tkq7bHAFT0a7Eh2re7Z9gR+
l8Szi4onfz8vZSR5yU1vHmFrzghN4kcUDu+8zYLhZ+h6W0ovT8/sZ6DlertkFfG9
qnJOYB1BHQgftspfllh/ATlb+VKs2Yfb9GlNFGCfBQU=
`protect END_PROTECTED
