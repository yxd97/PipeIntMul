`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w0bykYPqNyRkyr7StbQfx6URUkQ0sO30P0chUBfxrRy/4Otk4Oczu6Lh31c/60/o
vcC0d8sRYe6KvZ6UI8cF4UyxDyXmNiIFtqxJNctMZDSMKOFGe/z5pOPiT5bP6MxK
Jqn02VHvRfQ4A7XNJYsIHrr4h7aMcbItAS1KmJwVsvI13biQNwTEu5kRuEqkylfr
HwGy68ybspLmila6n2qUY5R3xlmP8CDgMXA0prnmnzhlTsBCR1dqdy3jz9ld6r0I
zZPh4BWtrQSANsX9UlqJLIeYcoHwqFhTmCPUVRByQFGysqoL2iwBI6saUpwElv/W
F5G5Nc+wANX1zCOUvtab3henvCISQ75GLk//ac83YYOx1aeHuZRNAivOQsmIrDT0
22W0cUO3RxrL1dJmC5SJdrmphw644nBRgsCCOOTYVss=
`protect END_PROTECTED
