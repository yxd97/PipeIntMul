`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ma4/qS1Jq70qzpXWI3tGzjH5Da4FwFLbpHls4+/FgcAFEsqt0w4fEXoZvXBxySmU
7xP/koZYv8dwGtv+3IdqxLvoVceaNfsgToIOj0bOVf8JOB6h0VhFmnO7JV4Z+6u8
CFEHsJqmFbBq4pa7nym16cQ2QUAfaPYfR0YjeXwI4elaTjo/MjUseBPAm/zrNqYs
kTbwPg1h4LkUddSRdBXjFHF7e5NpBdlgAwT1Rn6oIIVBaj0OEEDoZO7dGpbvn54Z
kccuKWSoV+apwAtU1rWXTm+XbfNYgtBvBoIWDgLrvfzd1cX+RPtCfNHTmszis7Mg
/M7KTJGbr2+c/KyVpAxTw96qPY8juMKTXHtxjMVA3FMKev3+S7J6avxcg6duSfMx
VTVxC1KMjHa9cUKbgfxBOZR6gVVrmGQ5ySn8HhIiXFr8wBYf1oEKJZ6/ure70dQc
RYD3fRhUgG3SqdCZKla8DXSrxSWBG+frBc+vvT/AA+HWxCyXqkCmnZIF0C8HCIvR
WqSGgRu06unWLnGx1FRqtw==
`protect END_PROTECTED
