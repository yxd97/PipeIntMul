`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vDvvDGX96Iwf5ZG55SdyzdSUpnh51NIVdf+butocBLqo54T03+4csjPJ2DKEp01J
yEmY+GXwR/HalqD2klsawETMZBUgyc6sq/iNw7rUzytBNAHY/JoXeetru2wgcEKa
jopwnP2wC3nIa+fsP5qDeFWApQmg2cnwQWVX38re8yFi+HqW379fsErMcLfU3cxG
RcID2VbHRKxZbStkfF3aLX951sjg++QlPls6w/sgDVpdpKQdcWaMNf26CnYb8tsH
DP4xaRiDrtLfNaMFV9aAd97FNuB6KIvny/xXMWNfKPs=
`protect END_PROTECTED
