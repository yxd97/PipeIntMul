`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNPFG/255Hn8pIaWcyucspubTpxiwhSiXd9YHyGLzw/45mnJYUq0kwZAtO8XVzX9
haljAd7X3RgzFTFIW8mID/FEfojGovgibbKBnEUjjRGf4OPHrQI5pBSYCV7a/G3o
0LQZgNmWyGQ7psPnT5xxMi/Ix1uoYy29+grBRM1MSSR/g2YziY6c8yMhy0DOoxwY
HFxiF3wyJ2H3aXkHGJvgmp3S0rZZVPb3hZ9IgHsuEFlyk6O2ezevoQfZCQIKXjQ3
ksw5KkeOvqOJ5QFCtBAu9LTtLiNrdOdpnOdybkvntKEK5BGbE3Q0DlIL77aFmQJV
zi03rhhzOyqzcW3rBDBgmZB0/T3m5PVNFyDyhoNV5yD+Yqqg0wh6we/d8+A9USjq
KR7kwKFSNX5UgD1sm49p2CkTb0ddq+8vWry9MUocGcY=
`protect END_PROTECTED
