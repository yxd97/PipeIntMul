`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEu9rYM2wHaQHW05mlAOlHZgHdqlsZfn2YAh1rKtndIBHddQhJg97Jukj1BZ9v5K
uTcr+PE5/Leuo+eWbUKdmAZjTvKyZLVGudWzO/ZmBz/XovONik3nkEIjk6Id8EBX
hDVFYYSSwCcH2o4NJRws5rWntPaaV044jyQIh+Asyh0+8gR9cqG5MGKEusAHm+I+
uYzSCkznkTNfhhB6W2EozAJT74/v0aWO9s13/yF/79S5E2HkqdACyZD3MWW5eBKe
X+BkTfffnT9eDJiSswvNaz9zBJPhhsDpjgM6YD3TuV3XLEd/2oskmHrwIGVpXx2f
Bn3IkHzo5Dyb1rHU4Ih8IEQ1kR4rGmgStg04hDRj8zMwW2SO3NjfvD/g1Q5Tk383
6ENtS9gagwpGFAsX3t732wolQI6FWSrvOkjO5bOllWkzAkDsM7e+xSfMszIvBp8B
01ai5MP5IpPZLOeszHp79sAEuA7v49vll1w9qyOcbNUYe7yysGZqK2EER2hnuKi2
`protect END_PROTECTED
