`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nxxi6VLVuhorJd7z/ktMpjnqDGv6KHuSfCwiItyn8x/qLwiV/anRk+DGJzciv9IW
XF9PNr1s4Axmy8NHpEapxcKOPOWzuBoEf2mSLg6BGhd8YbyjoQCitU5VQWCVBHw6
B65j8U+afeY6zX0krjoH1UCSK8OVhv5feJC1+WgwtQH9nYd5UqASLJafRv5T4374
cOrBnistqPYMDhXwPFEt5NUdcyPtLi4l4B4aC+K4QvjK5NSOz51lkPzPXwhqaIm+
WKt/ervMlXBY/i1JhE3slqkYuANEx1wChizI+dyyaHUkwHK7rsp8jti+gXfihSq+
anJyU/7wNKcotJpG8qLXMgWNaVw6QDXFXnc1rh3YBNBreS/aDP1xZfja4nlZm3aQ
iMyFri0YQZeotLUFmrTYyvuWoGNviPt9rPQ/aHTiFog=
`protect END_PROTECTED
