`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5E2kAEFsxB2FY2pjt/8fQy1BcQwqPJVEPgjff89BBedOICrb8YV7XniZUbJ/ctFN
NNzok1hiiIepRkJ6nKYEOkAIBM2r79PRhHaH7XgqqCjhjxz/Kkg80hvewjpobqeG
/gzt+7vW5O61+wTbvMYpubIG4DX3Muh3csmaoeiFidDgseAeJPwp8M3SWlYt9kpj
nuLEC43CNvZ8sKV9sMfvl/9vpMsN16n/+eTqjxdCSaJQLPo0RWBN4LjabGYZr2X5
ivFFd987OR3t1mTgKGwVQO+k/BNQCVmiOL8ve/k86tunIO9vLc0ttHOjK9RCXb9H
Z15zQfBSJYsmFHeqabtu/law/dOa8EtLwQSLYl23fVC3QRO6BZp6gQ+4FsB9SUzi
q8vDySpWK0WLkBji9SMKG1LNBMZnMLyQPkGEPEoq7w4bczMsK5u6a4AvLmIXJKnQ
4yd6aI9Gg0x7DDyziMuLb49lCnGE9vh9F+oino2cgHU9juptTKu9vj1lmwiVcVU8
guLWFYWYrDZ3552HYeUWrjoJrrUN3Y0+TwgwQv67+GxqwTqIJy2QGu8gN2BvFq61
31zgI1+EZP1sVOzgbv6U8kHkMLDnFtiuBUNGakx364AbOwetX0VgPJCDR/q0PdVk
vD4YMlkzQnF1MIoBxRJkQJR5NVJq9CH2FSxQ7Nf7uVvk40oYYykjCS2dbMq50PMI
CVBPME17xVOOYuvYX/v3ToFqZoz8cuQwSGk52FyRiel/AeAoBUIUC1C3FZJykLv2
HqHoBNavTM1xvw3bhtn5g5kayBMXXs7RTBzOOUD1VbgTDk78uBQW17sHPwk4YdWW
z0xzMxR1dNycRkSZvaQCwx7h22rSMNhkEkoI045/I3Ff4ZkGorTDU6plEGJAUx36
i7ikIveSjpOlcazmgOEsGaM9HEr9sOc9Uww9XqArjf5VrUZN+mObLHTIrgJwmVA8
XDkjwHZLQLJ6Ng6FWRD0etS9gowxWJmVH87K/LrN23ZKKM/+N6FplZEU65m6e2dc
B/NZo4ru2s7mvm1QT6mQpo2Rn6Ynk7AGCP8+T9eT2m4K+gijAGfLo2/WTKlQuq8j
OVUMRdtisN83KGPwRIdP4tRqEhpHReUNor7Cjd9PRUzcHdMiNTZ+j3/XtIN8GL4H
e9fKRy/KqETBuce1zJFc54yM5Oq54Jd17TLz10Qr0zoi7AF4VB+7dNLwAJOv4ht5
NLmajlIS90UNSi2L1T+MeSafQLbof233oIe2HLk9bmLX/PQZThyvzGtj71KB4M13
rNn3ov87Bpx7JDDioFAqVaNhAdkC/EeInb0mAURr2PuqjWGTF6Tof4/l4pflEvMO
0DJt1Zykbs6MVUbmubt26ZODvzdMaEBrvVKETA2xpE2GUCAVvj3bQUS6SWjW7mHu
knwO0ZMI+/ECphCYWdJce/WJZCIy2r7+Tq6iGQf065W2vFWqgFG3qcnexVa9IMFv
1PTH2CeSOqWTH1yhpX6dyLMLZ8sKyebBwsTPlVQtYPJ+i5R3EwefkI6HP8hWmvf6
W/A1ytzMQGaVUxijPo5ixp/enRYW31P4wGHEnowmpvI0b7OuB8Ms7re3yUWffbRq
Mvw005R/NEv8VwGwok+eEeJIZ4Iw7emnCAzMYzdYh4i6+TFLMpFZaPEZlAJjlAda
hkEUvwEQsbkW/xlXVSk4/N2I/2z6zBRuyxUqOL6BB9UJcpXx+Au2qhufQupYFrHu
orBHMNUS6fBBwPrjbEmya61RSK/C/ThmHt6Zl16eFdOuAgSU+BLmGgl1wKoi1CYK
PdU1T5XJcqHmEIYPnz6fDAdd+ytID3hyI86F3hSL2uxC72+MqC5+fLQs20+pQwZi
N+Pp9p2BDUA+HQ+vOqxr40OFRjDDG9aHdFrHVEHUTgsVG9KtlnfH/IL0DKZTt5hI
SDNiWJ+JsGDoekl05WYO5Wr8l3DkVgJ1LovEcrSKRZ9AyxaEasCSyqk9qEDewsVJ
NjEsVw0sHmxgmPSMRBrY+clatk5oy4KzwoYPw/rlPmvokJWvJ9CGohoEj+ZYr7fl
cxMpeS6Frr9S2rU+2bG6RqeDsN1ba4RrXMdN3HMzSnFnXIPcm9+hAQIaC7tsQJ8O
JTTZTPfqIL942ZdeILxvdXxJQoAjM0Dja/K4gF9MPRigQWiJOsKgNsHhe8j0f8dT
OMhzVnb5uECitxAuq5Cr3MEsiClnTTNbLrZgFbgajslDvcLc7S9Ig3LjSQLFntvN
+Rm75GOrLE4X2RgCyl+/3Q4FG80KMVR1fMCbP59HmaHmc2h5X3Ib7f58zsvfgy9/
0aurKSY2UsTXpiI1+UWuHkE+/LewNUzfC5kqRtYqbIO8SpAy4x/wH5ihtiLXQ4qt
IIKA6iZelbhlTpL2jBYC0jiHHaiXvjK3KCHYEiImMnVS4vSWL2foqd9QBFXDmQNI
WmR4fZyP/maDkxnm5FZLBCKWTm91cslZNPlKCdo5bPHTR3BZSupabJS5kkUsFUxO
rIDof34FqEedn7MKAjjPKcSO3rHfZj4sNWNRLRQvn3Spu42y/fCeqM2b/N1A6JM5
RSP8XwWvVm1KWhxDkmCmqnV0tRFM/VDVL4BP0rUHnkoWCw8X53c1uJvuJQB8EWlj
BYm7Xl0QKoZJ2adGh/R9iWgeAlMddbR6/tUR2FAgHv7QbwJkbIYnCX955HpLqWKh
opfk7i/zz/m2WxKkruJEObXofWt33grEk00HnGpiYbmdA7MQzYW4iN2Dp5b5zmQz
slVmFEFGrn8LA6CyD8UY2oxXN7FQW+igrWmIDsmSuCw2UuNf8fq3dqtVsMbUGEud
XiPF3nZtJNw/rksUv9/uKzEEUNpzDXg8yAtwB0QJwVfnPEwTif/aUYfvTaECTlN2
gHTFUTwTEkDVQ/5clqRKqaShhQdtQ23O0Dz/BrIxy7DUy866dMWrsZ1utM0QIsP4
YI8RhgGD6PKdB3g1XhqffNqMMVolQtRyLFySVkZP+TWIvipGHLdARrWD/kOgDBpZ
zQv8aeq9a3DAH67wJA4FwNZR8FJ/tiNuoQ/e42XGz9Vs3qKF/TNh80zG5lS3OCTk
A6sPm/aHyiPX5sw9ChZBK9RoVCnwvykDS6YjqHXW5pp1pEIEO6e6mX4No3lFfiO7
QQrcVQUr5L9eagQGHrtE6ACx8Pee86GLd05zViJeozAJ5iyzjcNcKmEgzATqthw6
NOUFmurZH+naHogk7/ghfIJxkuSDqBHqRGIDPND/a6oFB/0ZgH3/rV3Tqeydo/6e
`protect END_PROTECTED
