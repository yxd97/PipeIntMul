`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VI9k7GwnQX/NKqI/E/8IpLrPpahV3Z5aDNIO2qqCGqWgC+oAkqrqTTC9Wmozj+yc
xBYpdk+m+Ed16jgT9s6wPnKkgycvcNDOOgfOB+I9nrFJCoK6asJpdXmXFjV5vlfj
Qqda1UdEw/3gEJjP5ANaCEChxM4ILJrrZ3z22Mv8+iSoKBDyWydg14TbEIU2YT/5
FEytEAWCWUA/OiBFS9XM2YWYHScNtYyhOP1lvedmxnSyve7PBUgQ1AWi20zbtN6f
m2X9kY9PlbEroayGV1PCv/WZMQmQQmJr8zXg/f8koOBjZPVN7wUJgIo4c8HIpiXl
DtdH9QWyC/v1RZEDi+M9vzAum4EaiCgC3j2tnBN+GtL1U4YHEUN77rH7BxU+JJT8
sZ8/KhfjUYLARbPw6gfrI8/mBf19Vg0O/PkPLBpZJR3LIWjCetdqjM21xvVb8pJP
rKC8OFW687yD4RL6QWCPrU4psQhT8fDLl7W0+MZwWhxjbId8BHXPGlaC4MPS25Pc
8G89Z2onnVaPHnUgeWyF36S5JbhNu9MIRhJwm2E/JdbrI43QW+ayrJEE2GdOeT/d
0uABU7Uu/5Z/o3etM1jFY4IA7lITNg6sZvUEw8QroBU+5T4vE+Y8WMyDFIK8ApSC
SEoIC5FDqGSnOr/1CKxQCVd1GabEcX906YUdkUzpZbq8e/0DAp/VqmpQ+Gtzr7oU
FKwr501rKmfEKrYsQlK1wD8QDzLeF5nzFl+42hVdNXnb/zxBHulNgc/TJ5kXnPa6
MD/MUm488WgCiJqx5xnW/AK5vx5OwMpjE6vchaLuuIfHmjrxEjd2blITZ2g72vYj
WLRMl3/JHm7fBzkZ/pyq1m9v/WiCjY/Jy/3ZlXBBo3vRYS7Q5JnbBmSeNl3sqjZu
mKiPVByBW39Bq5a7V21dPqAbnpaf83IqiWqBRHXJC95qCVErNdKw6gW7ZBzIjv8i
sRDg6EvPhn5xMVAYNBOLwOmiLeeKtj4jHwar6AHubFTmkINLtClG0icm+awjrosW
3xxruwhaRwAvMGEII6hfhxf9SvfbFNXelSxdqN3+4Kst6Uonc48Lm1/HZe0hMFPv
ocdXdoBn+RmlC86R8Y7hnPWLD+IJm6omTO9zZMCJn22wBWKcCC2w1W3zbDIvhm3e
3zCeAlk0kiHQ1CzOJI0HODD18Bz4ekRCuSlFfD3k+WeKifp7d0j7hMb+QPHORFrQ
wxUq491dgyrhC8JYToPv024LXzWrtzTjQsFWe++JO58F780brebgwvoRthmb6CqC
5RTKPh5hDMEZW9xMtNp29jBgMf4bStBIE5b3xWf7alWwxUlcCaxMfscwqxGByHRC
sdngnGHjRM6oZxrxEWMJ3R/0eDlsHdeYzevMjeXIuYA/k3QMsafi8aZsyKsb/UV3
XDjrC7u+ZsrCBAWkNmzGXNbTsZOsjMLMroZTDRW6RIt9+YA0d3Oow/IH50c42ej5
OPuGTAQgWGZzS0a23RkLHAPIuNmRqVJCkArMH7+8kNup+N44Pv9ZB980HqVeiqSW
P0mR+3ezApSKZQTUyvK6GEJqgVSZGB+GTo97leA4kTXO8wiR1mXCOQSQDFdq0YeK
oNv35LWo2I7/RYwQ7c44c0rDGypksOq3tMehR7SS8Nqh2efwLmL6n6yfVaAOpXTz
gKZTXodAUdwT2NQy8vVHFCES3p2jzyp6nrIgd1PGBc8msgmg2G58kzZxiq8uUv59
l8IbNUnk1+P2+BYDRaDiJoKmxYcV1zUUL2en92oobTd83IceN1mY0B780MJfWABT
+HWirxra43F8ci7XnXRlUZfO3A3piEryryP2bCTQyaiw4k3aM7sAmjqon/Pse/bZ
BH5CVecYykn50ycmf9sooQAamFm19/QWAVsMZl7QvpgOBhw/HlBcFEz66u8DstTU
Jbtwjbn5GgqCut3PuhHiruE1syWuiBtEe6SuVK6ISSwLVfyx1KHkBzMV6j40ccv1
jPdlCFK05wDvPrd9711GmRjlL7XgtjPfSSAXVOIz/0pqUHv+58tacUwsPvbP2fUO
I0Tmrb3SppG7DvPDNMfhUK4CD7tt1y1tmP8vhxmp0RZq7AK37SG4fr3aeMG10y9+
7mDDjU+9Hgxei58yWg4nQdJulmSwf5Gx23l8+fRvLsKZ14/NB3+KyHk7vIF//fRl
25FF7vnNJ3OFniW+dPXaeez7USP/s+eS/snQV8n5PzaNH1Nzgy/Z7YxPUG/3HxUu
4gg3jMVA/r1GZ14Vs2y/UF9J77ZGmqwX4igxqg3ta3KsfzzzQ2EyQuM7F+fmcKOL
/W5qf9gM/1fnWmN8LvPvGGWu/0cnJ3uSlbt3SkKr6t7s3i1vVbIDDbnsHhTQez2h
UgHIkOvoMD44cOr3wvoS1sPHRaYKVu1zB+tRA3VvWbhgrT3Ha8o/Vv3f1r9JBKxk
BvsF/84Bk2RNfaZqiFhcNjes/eHUhjKZMHHp7yI0Fgl6K57KAJ0PSIMSswC/+7hG
e77O+5ytfcPxkWUnRs0Ik5SqN4YAdQJAltv3//tu/p2U85rYs+hhSECSJLxysUNq
cGi7hPkvsy14jBD1zfKb9kSddvk2IaDOU9ICRDZ+WaoBptfDN7u+pp+I7zAIptHW
jAi28Zx4JHy/qYa2BvwppFTvbbTwQ4/jOIPB+VmRAkP9PleI+9hrgjGKPeluou8h
1/coJi1HN+p+xhI5z9n094mcyH/GRWlhyH1Ia9b5LzIBRbfjB3MYWAovJtBZ+eRL
JG8pIzziQgZExQTxousvgSGgoraBCKehBK9i5GN+KsvzfDe6R9h0Mu0XWTF+BE1t
XPOr9iRxA9qyJKK53oMVZKd7WYnIgRpMvTJdqRa4LqIy5FUFdkpc2g034RILwCcU
6CPJ05dNGv6gVgQjNizbrIAgEfXTthNmklR0QZID+2jvJ7r60ZuQIWwfeRlo7fWw
ur3DWlExI3XtAiRFsHl1Os6TK2euL9vvPW9bOig5hO0fH7jQKdU/oCv4nQI+dsW9
SJxshbvhbwpuLpl7kfqXufS+sYCXerBInE+WuHR3vx/It1pbMN+CPfuGNW5Rheli
cUOFzjsJUPHPI+sAUrCYG+MSTM2w/EgY+HivNk8foCdpHky5Cyo3PDTMNt5n/NYd
1r6aVKkK9tG5KG0R0n4ig+Uceb+SIgfNgDMwsl3XitNmtOoZfvL/qR8uLxUxZGUW
L6aE3FYBMuWscK9VeOpNlAMVRx8LJJ4DjwcMhL1p8ZZ7j/AydcnGW+iD/USOrp0F
8/qx9qDIKA6KqznSbhxv/0pqWHTBEtXsmq0cRvhENZc9h0FEfiI4Xgz14F4yiNl5
gLDYoQPOlBGJcKAH+cV6xQnoMBPkoAV4p4M2t35+d2riPiogJl2hxKpa+WcJmXwR
8AJwtx3ykO0HB27t8FwqqfopnYcurUh4v0dlTqnteRQV1gJiJ39oOayFmwp1sFwv
MY/ftedcrXeQfqi9Qzwbpx1y1VsMr2hMnHpLp7XD4yo3217DkEuu8oFQt1C3MzPN
qJ58OdAp0zzNlpUwfgw0iZcx1R7bK1qPLi24cab61C9sbf/Phpz511WfXVXEuU4N
eV53hzzVLdvkW9SJs0sW2WwcsSRwDMH6t4iW3mq1iv80tPjY8/nYDhQ+p+DplNs6
+86s1CVUxTV5OKZM9OPgWNsSip0PYXtO0x1gADRcCKjO6tZnbOcdscYfd0obkz3u
phI6khqNL1C0omboBPITFheZvvMvogcWWngIY692LNM2wpRryKOX7ow3FMZW1SLx
5rbquxeP5P2HaSqfKW5z1zJo45Ikg6/IOUnG3aGbscnKqt0YsGeFR69E0uWKfQRG
M2enbhFYpLSzslDNSSc1LWtCz7YK+0vkXZvBsb5d9Ig7aDAh1Ff+9fb6yxMf65Kk
Mfm3iDPdp4SIOn/oubeEJ25A3stSAu557kao0lRICVeZIXH0+Szl+HFI4s1H01Hy
M1lrpf5TymgnoZcYtrdTSAmc848NzTXx1HHuf7h5LQ3MNkykJTUab/suMxRRWh54
xwHN6lT0UzgyYhQ8YTyW+bu9gp+UFlBU11pYL4N0Q7tYT1hTtyXzy55oJYmO+7DF
mqmPz0Cw7uFLhHxVf4Df3/6uLfwt4cWUghY1lum6GVPuMkFvoJrA5u3UD0H+jtN2
co35/p0m9RCaK9fDHAaA2sw7vtkbLv25gKy3plF5G+fnx78+DUvEtvzUwMO+TkNR
dmZZQLBkfYwMy+aQmF6g0jqlmi5N2/GvgG87wWTvatLiZ+XpguIpyamXK5ba90H3
1EGRCG14nZGnqI+6l9xOwnJH6vD7wfg1+LnjqCC6kvXsntpFx/VddvI5rTa8eDyw
5i4+skf2veG6Evu3563OWNZ3R/g92TorH0XkwTh+igg6Qfwpwc0HfKNIoU1WdM6w
bcDQQNF8NOcoLl25NhGPlH4fNN700Uvu1ib/XAr/K9z/nf32FkeQYpANPKQ9hsQY
uzkodFkAXZztIlMaKC2/sqmG4eqIKo5opxILrHlJMNZzPG5nvjQHfkNzcZ7k4mhz
O/R/8nFRvDo8e6OC0qYApvKG0FJNugbarfrfk+M5vK9YXl771bqhI+tibOKGBh81
4JW18kWIRgJVLWjZKpXetKePr+dvZHBcTTwBfsh0NTrKYFdOJ3UaWm0vDKvbRe6+
hHlvm5rVAxjrXD7gKAY/nvvj54guKXIjRWkGHIGYcipDb2ifB/OLV27GfmGmNMwh
8G4D0xIiDWrPVpwuBglHynNoSWDkcr/obkVgRF/J84aEG0tb1dpOWV2UB6/o82n9
qwnlscs7w7uh4UFlF8DG/qEOag/F69qCb5F/Y3msxmz3UMt+LY6I+v4SOQpdg2JQ
hTBMVCXzd7+gEXoXDfLQRXkerjJ0QdpY/vQp0jvCIetML4CWc6h5h2uNV74riPxc
AmKTHwhvkAUWfsqgFsAQbJhPTpPW6rMHApzCWC/tUSrLoOROHSolOxl0E8GxwT58
kcRLdx3Qk36rmNhhTbYnrWcDRqm1e42CwA8i88P1VtW2cMIzgV/v9KiGeS+isA9r
ELgo9lKFG85uH+EU/4k9WflMWAuBdRiQ96ycWDUlkQ55g0paHyf9EhluJR1HQAqN
RBRpyz6zI8BST+FiPU+Tqip/c35lAr+i45R86PWBAnZq0hbGn/4DBDfixacPvO+I
xdOL1AcIxoIJHxwk42Y12jGQkbZs3vOEmEgUxG5to2D+bw86JHaWwwXkeZhPDoPb
QDwKGJKAtYfMp6IMnkUImxbFe+Ep1gBgHI8XMeamCc2s8hW5PlWFAH/zPNPBE26c
/qxTEc7oQy20yx9teXd/cAS1tMQtnqi415RZ6t0jIqR/3cdQDPJSjQdfozBYCcKa
YumQZ2I61FoP2fGGv0Gu6q8fQZLpCEBEC77itrA9d9Sgkg2gVz0gV3qLdVlYcTit
O0B86/5awOuE/Z9PdIYr6AwlnoYELrk0qhGxuUddIViXuTtm+lzI1rbcVhlBWVZt
Xdl3Br3qK9mDkTFABYLqNJlVvJP8axJAkBbC+W6M69d6viu9KXTjNJKaU2kGR56E
79yIhCTskJGsu9eVh3QZBsG9r0i6BNNmD7DvUgnBObNwpA0ymO7dZZj2I30l+SC5
6WXhLZ736FMPTRLK+r3SoEg353k/RLPHIzjX+AtVhQ8wX0vypIgqO/jJu7jGO2Y9
fBFLPAvRf5AAVzhMqn97NpyeGGw0MDxJZb/wQZEnysFoo80zBjaiPuYJV/oruiE1
+ompf95gjp8uzHowQrZgTd3Ye/6mIpHfo7i/j691Obirzs+d+HM6gCI/qLkPpo6J
j8RA2YrLqskJZ8xM3XGhl/xntIO4lcOsDHk8kf1jogyLrUD/LO57rgI8OYvelHRO
LdcfKjb6/u46ATH6zawMtrvqoWAdQrmWnlz6YSL/r2Dw50D7GM9W4wOxtPIeUURn
cUYGibnJqMRM1upzbl6O36mMECeXlFQ/f1Z6nHhPY2tQG7WzEDObSkQwU9xdiUGx
FIQEjEPSTCt1i0sxhh3PLVogocsGN2MkwkOsjMKDKaAZvGbSVdy9O27pU4jwQR8x
+oy/h7sqLsSvOk9AALg6rqBNkAfVTkkELfyOHBr2d5gZDjZTdWiW4KA1L2006snQ
36MGUmW6WCGC6CgOTs1VQgEhrAx9dAgQj9ZdTLV3n+HziDq08uiJngQHaabcG/h9
QBDEkzivtCNP1dEH/setVNLiXqmk5T2rsO6uvMUnIQ6mCPEUateGbP8u1qd5Z4X6
Ho4Z5rJ9y4Zr9pfICgO6UIjqDqPJIJLbuSfRwpin+Zk+Mp4MIYI62bs93sxH2Tfw
TBZVcSNn0cj0PPd7mQZD7KynAiEDtAk7BmIqcjE2dycAbYR5uFlqKYh7bRpPEoKN
pvy7r40ND/cN2FX9w83hkBOfv1brOzR7vonuRBA8KJBj6IhUQ/XXz7wYoiiMEYek
fcSV4/LqC1iZXm7t0euEWVXOBHQITYWB9Cp6dxTUuXiSJm31jwRBT5ziHoVDmuPh
lTpJp/2F8A3dUaw6ig+2d3YJgxHqZ2hBkUtDvFGJhqbpf1Z/Okdpj85A43DmC21J
a6TOR33JsBnKq49eHOwgj8dZN6u0dyZ6lt5tXWL48DRS+l4sCemrbRrGs9JB8Gzt
HwpGheVkUMlyyC84ZuREtA8gaZKDPnJR3+0gc1WI9CauXr3MSmKcV3vPWWPamazc
NKdmpTD6j6Bk7R/b4bZWvkk5HMUpAKNhTD8uyDtThHijA/W9GZp0tsrl9HKeSyHZ
62zvHcdZ4Km9v/N+X/UmBMrTQ3dt3unO0Hn1/+j1WusTtvl+u+oB6YirvWqP0Cde
XgcuVzmGAh11uxgR4rRIzGlSmXvQ8ATrCkpWEzWRNNDnUlOiUcm6M+TAzwMjd3lT
Bc5SI2+QZunCSHPIKN4fOFWllWTwhLRGDFaAt/cO6z+mQWPiPlXfqB1k85SQ4UZH
tY3Av+hbvVQGiIqhyhvZJapHuJyIKj6Rj1xLLAIAVLkqwPqptVB0cf8j2rY4T3QH
D0stOlqXuiR8LthMbxsUW7GYsJY3C1nTaGF/Q+itcbambQRjgwQivsAWj/J/ICJV
9KgAlkLJfeHFY6rk7mLVptTTEDimM7ceG3yE7jhmYDRLAIPDLXylMtxSnYKAtK+q
cr5mqX8nhQd2ONx07fD7q0v5sYmIWnzSV6QI9xxZAme/X5mAMiCkfjY1d4Ea50Vy
S3W/xV0sEt791TvD4uojUiqkwwnDeiPZ8sIsMTByqgnLGEMkFzrlewMlhMoLX/sq
IHvUDoDIcrGSn0Nhm9bOMOqOJ8lrDtVmW3JlfJcVz8JC3ZdwDkfsekyaEsX9vaBs
L2ApKUpmJfpPBLZn2FewapsAVGGW68TbLMNDdCpD8kx6vYZwu2b2dLrzR5+fyltG
p6nfnmZa2rXlOOygU9KjLvkmAkMnYFCtz+wrZS9/sI49QfIh78v+HUNFN012GsWU
2vqj5ZuPOgAESlZ0Kakz2g/m5rjDFkykaO/AUVcexywv/cCNgkC3iM72JTSSluKv
MfGLhn+ODU4LdyK35a6NY3SlcAgpQuqEH/rXCdckAs1rC0QDxXughKr05iyrptLK
I6Q6TzCGcUvyXWNX0y3Sqrb9JyZ/hCskQdhLGAslOKpAKRkSqOXkY45Auu1LEXzx
M/26HFgV3W1gw/lp5voERJX+cgOMvxRcViZMde+FZqZdxvBBhGnFCKdVMxgN0q16
mE3LuRyLOGiWMmBtG7O2/EPyskhE2zFs2+8QMTtEkDIuy9G9D4BOQqI6mXP+Fn3B
+iAnPQGDIEjxyEDZVKvYwCMffcPBgcQNkco3awVS1Re1c6hKbMJWBpzEQw58VM2G
uQDIZ5m7nI0geGmbpdOBYaqhj6T145npyqOGXrLb7ocJAH7EWEkOgxagd6Lb9lap
zW0s808oqaI+9ENmZ7OOLtzwTb3sayxInkgDgaLI+uWwJlOnnFu6R17LVfyuGAJd
+JZnyP2JpSDTxUdQCRp0EGNFFskQX57AwUfbIzu2RrlI1Ph7fFXtUlvv3+P1kAK4
E/iQruoxhQLJx9wHUqfgBcMvK24PAClHRoWzIZwA0SYKqEe2kb5+veeooM8Nw6hV
9gPA7abZkXTI+gHTJSYvu1KFab+kAsti/R1qnuIA4J4/4njduPMEJP3CsVKjE8VC
nc4in9EzuljTN8UGk8C/QBufvZEwJB4gnbbLn+VUiHMD72727MNtd6xC+AxO3dCu
SmHmxEsqUbQN2NVfF9GRbe8c316v8IG+2W0hyapyXVhT8d7sGMoYmTLlZTLotKh7
6a5wn88Ovj3zvhMb0gajZ+fshdZ2Fh2NEVjF2Xj3PJJzM2xgWcmyjqxKQQVrSGR2
uvl4K/W6RgHgLa3wr9RZpxfuTSYICEqnhK17kjxYV/DlxZQ9AI0QLBcQoBjo0sZ/
ctYD97YXYu4VNlPTt0ZKJYwxHBMZb/XqT5XV63/ohfd7X7MQ9tCecR3I6V2gGfMb
qOwysTmUcU7bZxx9CwCrQakJK5VKKdLtfMjqaeIwQKJY4BfmVkBNe2oPwNpm2GiT
jHTgcimGomOs7+q0Qqw9Xo6j2tK+IiCfRCsNgk/QtWaXJxIVAkWKchrcRDGJMhzy
+pZAK7sE1eA0hVOhQao9E2Y9to0aeHuAgp6u/dTFA2hKIu3bwQUma+gYsjSvMHXD
fYVo+SY/qGIFgR6/dKxhuofGiRaDVb7lUSirqJLOU7CVUubRSozueW3MGXGhncsf
OMpUseXd4y3RPd3qrSgUK6xcwNSb+mhntYmWUMDJEdeCCcP2lKS2X6RFRnkmIxau
TPV+nL4ytgRYoM5SIivUKg+6qUIsycLO2H5dO808NnVqsVVW3upCB/kpsHh3Q5bc
SoONQoSM+FiGuDyBXQV4yHtd6WTwDMFYnh17E7To7u1P4aE30lkd+sggGoL7yA89
feOxaP2co3TDNJ7TSqm23m3FOynfcRTQA1xb9/BZvPQ5fmlZp3etNYuqLacw7kmN
wQrj5SXzFahFZDLokjykD/7ijpeHvMWZfNZZS1IdWxehPbalcz6WpBFK2dRN2l39
oXm2O6Ua/C/zHPZejuVhkWGpCpNLn2MlkjTtoTJZStmfxQ8X5BokzjFqQZKx85LI
Ax1pGNXCy3+lpxZdoIM1juT8zLAtKzqz2c3qNevd3yQd5eTfztWT13wfYX715STg
mPO+yHHZWPdXA9HXYXTYZl4SONsvAwiR1ICAe473Lj62o9yXVyNlTqwkLyN9SH0q
P24GgPqGiubw5SqI0KWIWH7PGctJ10nG514UV04osoyN1TL0w+vyUPkJrr0hGlfG
3tkWtRZG2uxkjkSe25ns+GgGXKR0uZVXpfNcLxgQdLwx4+5WbE/pPItMhVBqEN0j
GCywxRnKOpa9DC2/78Sj213WFpUTwJKO+AzQ5ZDdc+P/LC4hx0/TeZC7mLa3y9fs
it2bZ3qqBvkynxR3LPD2+M30ZwKzHBqjq9geNOaYfTz4ufs9US7JsXe+vpVCO0o4
gqUIncRP+G2LWkEm5Ib1OCPNsAugOX+wNvcn4LRPf/O4FmiNFdelB/WPcfDlSMb9
UNd/fwU3kiZq9SwJgyzYIXM+4flTL2VMN1np47/moQ0QK1vJcMfZ3Sm0Yco61es8
iYec0OdNbv5WTxQ84AURIVh/D0bxZ0HXluCOqNOgqxFdc/AUQNGkoElQgquRPolq
uo2daryZQZQe3NMVVW8XhIYr71nANSdbnoVG0PiHTDTWSiby6u8nehr75F6+pyuR
mhq8bMtO4J6ckrkDw2zyP9MVARkkpu4AN8E5p3tzYy0xU2ynCPb/ma0PpaxxPuPd
MyZvy+QK801Yt/9tWRiVlLENULfL3Bl6OEMIVgs7/8xllG3QLADCHDhozXLEljMs
V6S9zEmLkwyVfKTNomLUEfyFLsfqbWlNkQvphOqK40nAjDCovR4Dlst0tQFIX+hJ
uZcQ5P2HPbFs/POF0KAtcXYN9nLQf+KtloUHOiY6BGzCHUYZ6z/kHPBYTKPrx7yT
4fmriJ2g4Bc86OjQlRRusuunKeY0mfEfb6YYLbTr0nGJ/jQQDah3IHiF9biQgWCX
Jz+UpSUlm7FaUxBP3AX7LCNwCtdBWOYzPqabNNvCpOIUes2/tLa7V++di5rHQJt8
u3krcnSg6rHoryjhkDGMhDOOxJ4sK0AMOjhPNCJ+u3ca7FfgBbvjvwSOeY5tl2+C
37G9/77L+V58jCTE6u3h6bOeZJ7B1w9py0vxgd85LH9P0/H7AEOxKZyFY7caaxka
mYD6RKHg834B1KVJHi7yCjwHt3nDXXtCuqVTlRd1BxS/0yYVbKfsUS3ET9eKB5lK
VXjSSAb7QIKrCBzliOyUMSi9rOI97JD6AaZQ5EqBO75/aElSHfY9F+22TSCLCQgi
sMhDOX+55Jb5c+atR2XY+fl6rUxwugL9Jy9lxVKaYP2ejQH6cqEP6mxNSjIz+JQm
Zn4h7T1mPjV9ICsH2UF7k6NAg2ooetCsyrvxGQNVXZqVPYN+mp5urqVhQ9mz2c79
Duhkh7AJGQOUCnDxSUa8JRnRoTCmK1fTZ8KCxDWiRp34NTpxnsBKOzL/hmweReqH
PA8UKLXJ0nQ+XSy19tgElYNA8tFoNmJnde83UNmDV/iw9dcqAO/2sBPPWBUZq+J2
C/ZPqzCoqU4J9vB8jevc0dFC9TtSNuThiT92W//yvvKSfELmek0N7jEGHxcUQiLo
O7hauC882d3GlD74x1c8uas7pZf4QNXpngW2gJ9Iekvw0L0FelYdIg+eKFf7KcEY
lgEQUgS2LGeO3Q0jfpLEyHIrU+tqJQqw1aCMBCA/JLR1srFKEkby8kV4nXC1g14y
rQ6XU724HuzAxPeznRSeRlymc7BS8pT4OGC5GquTEcJsoKQ3uK/2Y5qY0qJBczrk
Ze8m8aytG55lY6KxqjF9vWnEeRhpAT7swdNoU88nSQyjUUPFtXE9yaXVeqFUH6ac
1t//aWz2zX9Msi8bhyClF0qk947BFz3MWPJl+/0ZIzcKZZMdYu2GKKLHkPUe7sl0
b8PBXHBKbgco8ETLpY1On7/C0osU0QacjL9lciZxl1QDCMKw28ApxYxJDkHZgjOg
91rlz1j9Gr8Inhs759VftixnkzaLeFvxmTEGBcnsdt5n2LEs7bDVr8roBmLyvrZb
9DynzEd7181uD8bgJk7sVjQcgzam3at02iFKWQp9EC6i5OOMD121aX72QqCgRUjB
TzFC85NcHuSHTIc0ZReOBTn9EN03VI5m9FvIsXEbTjsZvTWHsVTj7ZVA1eH22voh
8ngkFp1zo+yYKUckDay+b3DaZ5vMRWRsFQhYCx+gh8oQuOQszx03mHojEW5wtSvE
KDoKZstlSEQwWpRATmlzbd7AxLttEYH8OYh+pnddahzxrdnFoIZepAV1VdwP7i/I
CS02/B82JM9HrYcNzyArU55J5jKtsP9SbPVvAxD3O8EeVmeGKSLd9ztQMMlnCc7e
XhgTpe+1tFU6vTgUr8b9WWZ0z37gr3k99XWcSnPObWlPzKsC6d1gvskFJ6rSje5A
AVicAQZ1IBzfmn9fcbKHXqhjv7fH0j8QkwKMPiZw3Dw/HTTyrsbyS3zg7t7LEdTE
tU9+NG6q6g8jrcbEv1VMhrKvpbW8nyEMRj2Y+XnOhGEUxqMZK21WD10eShzj1opy
BjDK+A7cWvS4zsI/St2FGQaR8xZVTDncloS8G4hJOVTha5xVKjWOyPFiFK6cO4Xn
q7efu2jr6BF6G6mPStSTiYQO+b9gahVA17yr9afvZ9H2eC84QgQtpvqK6z3niF4F
vEWBLyjZxS4pD0b4rDZ6y/JnjQwm/lhIRz3hQh3JCbtVCY+BSwI2VbZHpyqZPdaQ
tZjLBF1MHBH8nDXzVr7jLsvZR7OztS+K0yhnV0aVuEBxtilxHxJsgVr0kf8wOLSC
G2kq1m+ZHQsnoNEKmwBEvjwLC0j+WXx525yMvqLkCXEklQS/JvawcuyfKu2CpmbR
+LasB3Er/Iliz2JtkxW/U5SvsfHEsqy+USqr4lsMU7KpdyACy2phArzOb8bAKnp6
QrrevFS8bO04ytLMeFOemtVmo8U8oJewG8SgL4k0pWrYGYaznzuMXuZE7Bwz9heg
gIeSyMRGMCi2NWWti9f7zM60jTyt5xij0xr8N9dnPai/cZfZc8z5iimSwJqOXSzr
MjBTTzq9Ji1CgDDe5GOUxVlgH2+dGTysB3zKbpqg5Z/RSF8eaR8LQROgWuNfE7jy
UI0d+rlHF4X9XvEi4QpA3BVlXn7yJe8uC1MFaiA1nAKawGxtKMjAOQmfwbJT7t6C
0cS5QvwdWWYLp48VdAw7O9a1uo/zNSlbjhrpu/X+9aBQLlr5xxkF8YVeC6JYCbrw
tvOP0GtHeQex2nNuEyYqn6gXZ9SiPq/kp8ke/X31Ka+Z95Ogw84BsInlRejPJDF6
4+xN8DQ7u64f0Wrcccl8UKYNtCr1eeL2zFVk9EXtMHjyYJpGtO0dFTgR9x58/U1M
ZJ0dBbST/KT3idOMqCa/M2IlJ6qryZFhcYjAGxt3y22bV9kFBaApwT2eFNVfDfdD
2EnORJmfKoMjvsbkRs0sQDqaf3o+KDI8eNt01160wvQyxoOrFecs7tuogTU642N+
I4C7dNvsb7eM/TUOLbRLhyhhkffqzy4CupIZ+bzX6PC89jGjMWC77MBKQmeaiOpC
csARNYx+keOCmj+MYQgBVjDmAKq/JT/gCmH8IQon0L+F6NrAAQVdToh/3bURLpbq
sbH3dYhsP2drFQZ+h1umT7bsrBMHiPQpeNn+XhEkJjBpFu6v2COfTLp/9s94/Sqm
ZBmIA0tPMlzbNVCRW8S7ZRjTYpCE1YZUaiarPPhyPU+d0Da4CgRMrw7IQCXNGGXb
hXsNtPLD3k2m5L868PbfHmsPlZFXAkZNotkB/36GQYADR501y1Dmx2AqisAK5GQR
rQWoMqCdyJqjGSfN3H7tREWvaI+Lik1O7yvpLMh4wampbf/phBUETzriy756r/Nf
G0y4EY8no4CtqlzGUqHBaNuBoIjAl3o3QgXkAiIjvZ8jPrG0qCU0BspddFjlI0eY
V064V1M0mxm/fr8uvxEPjLYADjHwXi1h5UD36X09ktCILhhAh6crt4II652umfkI
gx7Kp53Q1y0S9XU3JMSqCC7dLnSUTCmfYDFSji79QQdIPNdxNtpEJuKnannMjIxj
YEwlmJHablqN94pDFNirNP7x2mu7SbheCQgV2qnANJX4MSG1aP4D78lbQuxadglC
5lXRDO2hIdbamQ75wHBRJsmcQy/IcdH0cbEESy112yD5r0a/SEX/HRJav7dbfAQj
98yDeZKJitcyxx8JzKvglgT4h441nGguiLQt+q7NXO90MaINdfEoksO3ADNfy4ow
/ZXI1N03x67YniZWGtlUP2Lz/q/OE31SrecrqK4FHYRyxWNoiYkfz4KZPa73rL0x
YGL9QkwD6LVzkI231jJLAHMthZiSh6mZW1Ngupjwn6zZCFBG8QEKK+h2mp1cAcRU
ZTaLCs1IqQBmAC3z4Aguv+GdF4jLP0ix8viNME3u/RCS47/yuu2PLLvUp2uzmIEs
K1U6rL6/YmBm0RSmJKK5MOQ/DucbXcNmIj2F0K9zOi1cgWo0C7ba8HzDQ8pcoNxV
Ed1oCnR33S0egMU1gdM06aLVutZNSPPw7J38e/ksBAUQIijl/qBnH/Yl4E9mOoL/
3UVl2BO1mPtJs4iEP+YX4CVgT+lXj38vZ9lIgF0DaCXbsHTUqB7YPvp4F1EG6LoW
QiGjehHzhpqy40cwDmeQ0tJFZq6nvNwB6RyqO8mmSyXFxHGBIfAgpJoy9G3eRHuH
16W2kcmurJdcv+PaFZPOTW+BvZ87nxEpTUqC4UpY7XZyx99zS6XtGbo/YIIqPJn7
VwfmVcoIwaBhmwj/h7nvVyr+YpTL9ZV3lUB4VncndeOojo/V7x8QiZG7SCp1nHAw
VLEJVXvu2hitIdimXGHtI71t+obsw7r+XYlcKgZ/T3ihuLmIhAslrUvqtZv1fREF
jo2+hnJFy/wM0HnRGcz3Qz089LvD2kg6dhfe9qgY1Dmtpqo2M0AfHnQ0OoQXgUuH
RPozH4UdDmp/RFFhcCKj/nUKcaDgtSlxubW6AI+9FqAE9euF6hoMAD6iKa2siAvE
lUWY4CZWaiUuSebUNdkWzFPu6tYXCvP8541eXECoVwprLn/K2eos8x9qQqZLzRG8
laIwpGytx9lcQV/He4XBdPIEZCT3jjJrZY8RBzcD03tjngYzaer9M92vDnEMPir1
BGm9oLLbaVg4ihEZNx2ZQNyhg4a0wcXYVARel68VL8heC6XA9cpOYrmh42UuIL0L
pzEWvsY17IOoMDhHU2ath+/XOhV3EYFnwCmWl3nLZKEkxI7VXedNR+YXa8c8zBxI
4s7c/FeEAikUN/TFOwXNNHUnZEMoL+lhj/pINeGfKMrbyQ0k7Ayxw6bX8gBq++g9
2IGnX3JQ0sRfLq01hQNbM/iE4FYNbcxSYubf6xIIF80Rv6Z8kyFNkX+Dx0KyoYXo
W8Pftev0FWm0YSO5r/NdKPqDQQRb57CNOR8ny6ZbeelJSvWCcuOAad1PkifjYSOq
ie4RE6A8T4otG46KtgLu6+cWuV+2Suenlpoow3GbM0z6VBuokXh/XivZm8SQG0z9
xqwzfb7+FQYkVv6f4iqIyeZV02xG2qalaKtqJEli1Hk5IRxZvfYiE9FFITqOyKGC
BcyCk2gp3JBxhc2Y4NvP5pXPkQZdo1oFP8KsPSyH5YZiX+7UDxErBkVttMWSp92Y
RysaBhDRBcVnTNKARbXTzRPqmOLcwDuJ8MvQhueQdKQDp3HYm67RqandU7xg9iMI
VK0fDZSm7RJs4gng9jLny/SXPVRvGwxzGesPCwsHtQJFRXKlqnYoBofsGjbtHJo3
qk9411Y7u4iBe0lfJ4aKyHNDsmhTHJDBEFNlpsb4xNKVwY1feMRz494E36bvTJfg
VnULv785Phbj1JrxVJ7FusMi5l5BvcYdj1iVWKjSeYtmPBrQN/c9mb0gjlxJEMc+
QO8eNbS/Q0ypwxejLgxwFuExmjjtBz8EON825VzKDXmAQ1DjQ78kopyS1jbR0bxz
ViR7zFhp6JdJ8F/6a1uGJhyUwvx6ylFzmTWqv4LRpyYZhQqoe1AtyiqCts+jKSJA
dpIixzN3HMdcAZGrvtVoyIe3t8W0gW2BTKZuNBGzIe3vFQWFxPIiqpxZ7wI/LrPX
wKT4BmyfJ2zRxh9nh2nF9A6HUft9rIeHbfQ+Lkmpds3eiLuxIPi9dg7diwgp7pUy
TtSuISz0AoNdLwksQbf4HQ8Q7xEgS+MsmD/JkWdCzYdPAU37XHD9Mb2GKpY+byvY
P6+OYGyMXAmcYfVSqM9qO0J1cjbcfbpT56V4xrDH34yrdyJvI7juMDNNTafP44lW
b5n+5L/i7o9tPBgaexha+dGXiH1Gbfo3rFaivGh5oErINbamV2TV671T/hygE0uW
bGFdYbAg/uvNnJcPTMPJNcLLuk9b96vL2DP7Dc0iovcoMJKhucZKLC5xzwnEi0Ok
KEV23wmxD8/NZtlijH6pLFWKDz/WOT3bqHry4y5o3RxqIBeU02ARYxKvzeJzV6Xn
iVCbqQtPCjmP0BcDynOG9ucjxOCMgPdSMGZdhqr15cvQ4rporVEQ5+YI3It3YmQt
EWMpxTHyjdeF9HRrQu2wu8skm1ljI1iwxN/00UabHGLrJAswFdQdaWyPnOr27nRY
VDeHVg2Nm9GKaBttSuWtOhVt+FgoRrpAOml5VrFg7wYiE76U3EIG8We87UvTPX4r
9SCwp7060Z9+ib/E+Y6x4nJG9aW1vz7Iv29KmTJE7E6+ByQT6Z/ftq2Uy34w+LWZ
GGgh1DTXB3o054yXTyZ1FcZ10hoVKTeylL262U6EKwF/bDnzWNTRsZlwDpgxWOaD
inIkWTCbWWeogRNMV9RYq/9P8QlYvS/idHzOO5HNudli6VtfsznsBcEQkdaiv3dk
nhfKJfngC+W5k3XfGZLaacsz5qdziGbrFnEViWew1vDlDwFW442BtxATSj+zwRio
ewEYNL1DAYmgnFzP2ic9BY3zHjawBsB7WJMAjSi2/1F5/Mra4dE8rQZJBGC8Y7br
y1b/bqW8h5RGAeG3ZQht/FqHtJWAB7s0AEnW3oqG7yhdIlGWIVs4f6fsG16XuqXO
VUKeQT9kC1wRzF73hf2PNXxhX+oW9DHSQQEP4PwIUF/ExaNtUktHJA6KyVRRb9cV
BdMqZIvQN0adiPaBJxWAy2xmxsBMIpjr9MHdAa7irTspioIaFYZis4kXS6iZi19N
u/goZq9neXb9atcCQ6aINDiyjtFLIdji19TFFnN5UbljZxuEkuBzyp+VHvk2jns2
DHJM+D4a6XRbhOurngxNVnBL1urqpXASq1IRpJfw+i9zfRqjNNLOiy9FvIDxA4nd
sIsBPSzNviaiTjXxAukhEOFPM87nnfgdRmM+6/mHQBamY9HAhRsm1njBWDSo6/bj
inmrOc9SbL4o903+/JVeqiSyltuXO2G6Cxw/S/L43JKO82lYzFQrOsd03le/S5NK
L1TGZ8oXBpH+TRNHC8ofagviMjjEGVigqWXFMNdnhN1AfgkvX6SnC3VQCPL1mhZl
yNR/Rdxt8y0Qy5C6SjJcRzTWJ3zbLCI18gDW727fLdxl7Vzx+6b/nd99FD+slLng
GbefH/Hxb5p/OG9z/JQfGkE7D0yGMRxcqK2sGwEGCoZxwSP1tSxpmUkgbi5lVcg9
MXoO7DstB+/xz/F3FatBep5lXjqQln2p6Z4bilQX8NnE2SdZLSHWQZjOffo9S0xC
plit6Vgan3FIZT2LVPrTJWYbfLWp6U18MAXAdpk0Do7eqLsMAKW5knkyQ89YqMyb
YY6VddHBqh/LwnqmDMqEwl83iEU3Wv7vQXMdQFzq3SAKGRRuxZzoEWWHuCl7HXti
qoGPh6QwrsuX2ogzPBgs9s0foJq8ru4Nyu/tw22baHwvH7+eEN6iHiReBAmLCKrP
a7ms8iFVzVuHmY/O+kETn15wqfbuc8VJjDNYdtBS7+43wT0SNa/Hi0Ei6+9qOgix
RShzvHwLSG9zhP43M1RW9QEXwvuOzPZHdqvGTo4VXN5OxjB3QRF5tJCgZyvPo23I
oKLiqv3Y/udWo/jbXHXB3dNZI4dFuE4J7FJGEfh/LyXzYoT/xdqlBSM3aukIQhdp
smHUFfqYPxLyXz7g3/O6RDIc60XzYLazhJxEanXWMIre+AEjXAkB6LRIZEN8jjOA
MeiLnzgoof+K8g4Xue4un311bzEQOBc8+qC4C77QAw/ABdYlWqRW0eaBXW/ucMwI
r3PjFf74nDcY5TGMvSPuRZ9oKnIZ3rpAuzpL41H4Y6aj6uyBnh9Q03RkwYc722D8
/VHmr9CkOwAou+PmPq7HUHvnClf4J/Pysi86v4F1E0983zTQvqTt7Z9n5ex4G6g+
aDS4ka4NH1CbSBPUvVzoVHeCDXxgymjA4RfY61R8iq47Ntoh6vNPc7ypcidl7kSW
MXN2Ws7WdEAujjai1x3eQ58iWCnc8lM3fayxttxq+58C8n14zvi1Yxzc5eli8aoV
X6ZZS5SdgivVDq1T6ufMw7n9toUMKWEE/ID3dqB/npTYSQbUdo4am34yxW1iELPN
d/ilDHfhmA5eAp/GhSj9MA4vXmKjrd75WVLWfsT7/ruR4Kywar0hBY7LjkTa+8p9
d0iJ361hIsh+V4WsiAP44yIykJlIxzWO5MOaakbCZG2r/UcdXDdD09zpl8MbN25+
NPpZoJT8/XkUpe3/KEJrmX3igo6RIE5VdbnLRGrldcawmTg822eEdi3VlcdRR36s
/7+HIZvHf2JpaeO/neScpfRzZM7Uw3XyKuk4aUB6L6eiuO9egUK9to4KYivMhPb3
qlRUhV2f4CCl57YIjiYhD0SVg2//uZcCY5Zjjpj2Io7MqPKQanKSRDvDTygilMhG
DDNF+VHZ4CR3MXS5Q42dJOvwTTsDGhLHQD1u1+h4nMfrfD/IigmMeDEiZjmMs30t
6mthoClu9UxTkGooDocqqHfYXTC6AAIPlbw1GolqjMyrwN/Vgp++C6lyTZ416QE+
ue+jlq/GscVzczeZkJch4y9XyJesO7ORLRrd7tPerjasao4bLyFWdz0FipSh2RMD
b9T6Lj1no6GOR6n/rvljE4OXojopDVJUQ/ojtGaZ4o0iBm0xfS4FeRjsoesvK/g1
rB65Vmw9cPBRkPYmMsSPhdAsnsC/HZ9mnBUp2JIxkRisYviQlAuMf6dzi7cEetGH
s4XTWEJUgNWoLoEESGAk6FuB/oY4bwG4mD7d64T/znctpmvcXIpqqwxhu8L+mzPR
A8Ssd5SKUrIEYRggi7crOeYe7HKIoTxj92grSA4pqMbTapu5kee8hHYgJDHAqmpp
k5ya98rT5NF9HmwEawXOvuR85Q3Ya4mEw0DPtcp8HpwmMXacmvuNU/Y2y5oP9Lf+
x358KTYz6SSKmgQEHkeDlwmbdaASdyAvpW7scGqCiVXiCCREcG+ba5DMt04+R6Ro
erVB/4UC9ASe3u599+iHpAVmgABo8BDh6MTmO1pLLFiZ6/Y/QR3ppLU1cL0mkVEE
6MjPs6C4iBnjncWX+sGLuF/LXtYsXITTRzMZYLoi7Yp+D2moKGgKGaY7EB7ke42l
otYR5Ufi+VYie+/2n0Dj2ESQr5lva2XYeXJrc1GuWQXwSY8Agd9N1/4JJZSaj47M
Z5aLt+nhnMJkrWghLBaO4MqI2WAQgFtSP32zMrGIEfWEuusHUIDS87lOBSlTl0JG
6T5UQeZIsBYlO4ssWFO/dTyo9QC8g3DxAzT/Hm1uiZaa/55RrZq248Eq0G7ry7zP
741Hn8adoybK5t50pEb5tPTLFuqy+dQA2zCi92dBVvl4TxI1TgJWnS/r2FyX5I8G
eg1Is0VvkVJFAKXtSU4OLvN9tupkmxD92M0HpsVtSutxdi4F7XC98eUKVARwlDuU
/DwZtNNVkjP5ZKjhd+tu/qwbkK9ixLgRTGK0T7uyo4osmc79G+3DAhpTUlDxxBKU
uCq+/dbPhwKBMcT78h30DAC8iGiTV78fIBnjpS35cKXTGJmMGSHuSoJhc/Ly9ron
m7TYXFHleIVPwQQt3Hag+SO63lVtHQldofTWdpzVQ0iBgVyMNKzQmRx6J/UL53Ln
4wH158UbqzSSrn9qrAbECs9l4o34W97cHriMtiSKqMgEyX3Um2afXfgRoRcyBBcx
a1O4GqRQI7QRjHYCqlyx9CqaNcJmw4UoVcoMRdyVf+e9Kl2kIwHV1acBAJpyLUfp
jDqJqdYy+AGRBqmLwHuWB3NdbIbZmkvN//FXiMH/Ib8Tl0jx40n99Xv7NK9nzV82
aqPS9Dgn4sTfsLICeT78jaWlOgNMxe/8WjU/uEqvznxCUxKyKMYZqa0OLeU9PFrh
Vasi9MtX1g5SLtcVq6Bw09dbxITa/C7Ers0Qi1pGp77uUyQzVt7WVrXIIKoUxITk
ZBA9rkhexxCFEXWVV/UKQiLC1WhZFEky2OdI7xuDVO6MSg4twDy0l6EwzGp7q/QF
5vzneoK8Cl5XmkN2ivxDcoQSbout767YqpQWcVk8xtD0+Up8o6CRCmyJA8CXk1KL
oPrjQhWtPoMhoW1dNab2TPWRBGEikMgkD/vWlxenzPZbon7c2Uv/muzu6gd1gjZ9
c+In8AciSopnpqSazfFPQtxSD0qNCBbjTk6oLCJe8TOJu72viZ7VA6oE9tES2ZA6
0w7fDNBOxh2n8b9P0Doc4L9td9k8AVVN5LJZQOFX+XPl2GojAdVqOxJ1w5kdd1NN
cWoSLibFyvb+zg+5keMKtLZRUhNf46jWfwHkyWxkD1UIVjKjTjwlMaureTPRdSd2
4vpk6OC2RG/sGC6jJpi7xDhpv8j1NN4/22+EznbTn3THVwd4fBuR6evP6K1artKO
HwL21y368TFcnbuc8CFL1H+Otn+vRzwyXymIGB685Ft+w68izXb6yHpZm1TVeIqf
dwYRxfx7YLgLj/MX2X0w1AAVl8vN6U2HeetPJpYmLno8PRs4+BnaxjFIPHLfXzZ6
r3jU7AMmKWqe8nRdFMjA9F5ZYZsVl5Gnw1uXgXzYFYuxi8pwov8QJge59sYohPll
b1mUUjaZjIodsiJ5jglN9c2cvUXuCJdH6UBxCH3msJ6/NqmF2Hq23yV9nXkHZPMT
9eKOyaqWUQ2gs8dqYuCf0Hny0jVKxRmim5n6LtiYPwB3dBo+u072vagq0irJMFHQ
TI0klyitBLEoXre0jwIjGvE9tBz4lCS8VfRZCxpW9WXpyYwX3pSFImA2xvkMU+DP
5mNSWQQer7nTRkmKEfp0Bo8/ufIoirCeMjVN+wexHHMSqu5RE+O65Ynif5YDUihj
PCne8WYqz+It2UhsoQXLBE0lNQ2a3k5EqrdUb2QgP90kXMkkQOYhGPzwQ43Pabq3
TPxSJTYX5RH26tTiwYgRiTHU91F5yLWODcXHSXuTdBjtVSyUDaj2Fkx3UT4VxWwV
8vyPSB8xMMZd6dDHMk/i8MKmQZKzyaVQlRDi/QM/Rww8p1YQLVa10J6RM2nwusj1
pQD8Rn+KsNY6Rl8C3BGuRYC0zaHSYNmrrZU5cJTmRey3Q/nzWpF45aHUsdUIanLT
hKbvn5ogBmRP4B01+G9sqe6SOcmccbrxG521tAbwqTjwof5NMT2arxv5A93u4rEE
RVg700q2SGbB2tZRnxF3AfzVZP1pxmZVnErWwypvlkltAEHpmIfU3qwX5sfx31aw
tuMtVi42QS321RiVC/CISVZRHn1nT+XhXGiEdfIpI+u93bIqSfoZbFmBN1d5NUaJ
wrA68oPrqgWgDD3JdHsdMGg0kZk/Zo6veVlAvmFGYjwVtf87oWOigqpadWkgtlE3
SPpdZfXQKJuk1zWsAaERjpffJjfXFmpalDvHktO7sN3AtSGY9oH7DCIujVPrWIVK
6HjDsdI84WRFA229WeLNZAuxIvf8axKmZao2EZV3q9O2eQRnfl+AgKd1CkgIr9XZ
CjAgzzXyHSwCbZg2psY/2JIIDeM29xY8ThleUOW0MZX8VlGkpFnkvUIGS0exV5kR
j8OLpT1Xz2m/02yMxb8KpJpKcA5xGiSV1Hk4CS1kPoq2rw3kMlV0wzu+t29AFAws
n+DdiFoqoUITyETY+bgh+GmuDfUmHVIvTstQlzn4yasxU0Sf0Oie52c20N3nTH2S
Z+/KhKnsaMM5bZIl7sUKGzWJq2ODqASPnKUP05GNHtyRQ6EmCW/xJSVOUtV/XT2+
XowZXhGJrFIKUuZJGte9JoChyU5q8kLQeWgFrW2pyBaWWuGIiMinfsD7pBRuX/zS
6p22Z38cK25i2dU1cChR0x+1ZJFpK7yJ1l+YChw1do2Wxg4/zpnkXwv2ahT3htqL
TRVA4tW7NGd1Kh2cy8tO68HIxNdYducKNmzovhwxH72OZEx7QwIjX88bxj6Q6Q9E
71CBOecpvM/aH1NMLzEtNutobmxn8Jv2SXaeC/YW4LrI/vdXUQ1rGkrTB5PB7WTu
/erZmkWTFgJ0Pji543v+BqKAmDNCYwjZDd+VpNXIxvPCm9330r353z5Q3aYj7meC
vsbs1Y2NgJsfO1E6dU39x7I1uOVZqR1EZx3sKZiKx3JuIFCuXO45a5HPOY/fEs4C
4sEyZ9H2lGIkIKsemtql04y/OrleZsLvLp0N3uQrNPQ24J45/OSxmCqIXu6tU5lt
qHnS+jxqVwB3t1KCwQkRQ6Z5poDPbakAmOxNqq3ZKd5VbimNBKeVdzhSbqlpvBkP
kdpYcwsWGOc8AJiJvST90YIGbZgjaSzwbyip6bKhtVYYn/YPpSXYQTT3rIERHIQ7
UqAriBthYCdlzpAFQdG3EqzuYQUYpY9wJ+hnc4NMI01a+1H8WLTnugptvOLQTWX5
0L1gm+9ZqO0dUTBjJjInZWPyfHVYyXvid7h5CMMUI9D5OOtcALIOdSdG7HdZ/vDY
k/qYVrnYTz3hvH7dmg+7yIwe1PJiB5nwMfatQyFAu8chbVWlDRxYqSvAfZCd7spN
+qngtACF51rX5ENaNDCG6SRpqlEB9ksi6HkHflSRL+SBuDb5+Y3yTHB/Q+sDh+tQ
bjZ6Lk+NjeRUH3sm+CLzTRj67HYV3pBRpGq5/Ni21Wizp/ZVUbll67SFKrEnjFVx
fg0Xcr2B7K+RQzu78dcMNs5NbrFAW0E199ERTts5/8ci0x6DNw9KmhhJAIRpxGLA
Hatwp7AsKgb8awmP7I11jfDdCm0Fq+/ygrU4gUJfkNpP7TbkBMI2qVu5nAn5oJR3
t50XXBngjsTiW0Wr/Mw4xyWtrp9l+kLtqVU35ybmtkVI3+v9PjFfkLW+bPZhhKco
butVPg+RVl7Q5I/Ayfv7zsMGhMdBPJxsugRxYPESyc5fPjorIOn6zvnLqGE9Nd2E
fWYMEiP/nWxMeh4vDGA1fBGToiWdTZ+p3TUeZj6MJh/WwIyZd2e0w/k8OqglTw0w
Hv+x6bnNMiKhZ5CPgLBUyptRVJkNn6zi4VjfJQiQOQ4jZstCh7DSmefXCBCsLy5D
UxP+OVg9ipaDJL8tGvIrj/sXIDeBNPOdyY51lXa5Y5i8DI3RGkMbrhxNW3jr7oK/
ZW8SPGio75GmDiLKGwsCvJqssLKb0/5T5NyPl5oPlq/kQb72Jtbkf0ac4lIl4s5p
RFOOVjFsTerZKCYXhxOM3tvpTIg2k+S1VIht9a6kZPWWjYvMCiLziBmvTmhbKrE0
XQojwOOKn/4W9FUErLWbWwAJS3Sn85jIPCtHncs72431RHqz/eygJSi9pyvs8dUF
xMfBuozxUvAgNREtuxZi3bMhc8UtTNkjqxK7i3MA8Z8dk+9dJzlFMUxZcy+9kEUB
VU2SHfKpfg0qJOflZ+Vwz978spo1konZ+7ES8bBI0MP/FzxFfA7NYqZXYunZCNGC
CJlcLWkcNPk00KdzeW1jGJ5ishMBo8p7Mdy5Au+KE5YvRKOFpCnir6S8wSC1nd/I
7Q/aIvpvjgESgjTYH8zpJBs+4Cm04MRH51HLEohff2fpyrBAwgNQVVrZi/B76wUj
Ixkc/PazR5J4vNRcYsjRkT2bS3OcD9dxeFQiVSxqUBEKwrL3RWfH5ia5UP1NXL9d
jRpbQOF0IMKIJLbK8QAy90aLcmrja82AyYTVEnsDWMfmA83DPa6YhM55LNenf4pI
KB31K1C6phlsBdlRrCHE4/JHOhQrceGe39GTAy9zrHCL4wmkwZL65Y/ecp56jrps
keA7k+H1NH315KLbU0giLM/aV/+4OA/0APo2SjDI7wefDDTiaoT5L0ZLZvp3lWuV
m41t5ePndxx94NK3B2eSO6YtZ7asiXS/xp9exfXHVLDB521CSIpuGD4e9zuDrnV4
s8pTFVF/VUeT5aqN+Hu20T29jQmuAYxupuV2F+bE5upi3ot0z7Ey3yobVnbKoUAq
ch07PvDwfvX5N82tgmAuZfc6xIr50o58LQQiiw8o0PIIA81BUnDbtiXv9/VQDBXz
3wE2bY45dcJp83xNaP+pq+PfrZDbc6Q24Wr+/+gDofuBuveUcK76NNW7DJh8r10z
/54V7jxU2sx2rtr2GUAU/oFik8hEwXUWq1lQPdutsBXYbiVrZ4C7wLxSPM6AOAW6
PuKE/l73O5P9ertll37Quium9cA4hN4xs5LTez3pDeQsqwhfSyQLBuBV7y2WLGsi
JfKoSOfP+8djfMwyWiPbMOlFajTdsUxeWEhXNFJ0n1RaYIIYBU5Rkylj4KtJJAkK
4PSb70679ucz6mazbci652qFgE6N+yYpmOfV1WqYt9EMe1CvnDoS7lmfKQQE6AYQ
xvgMHYtcQdJloN31W6NAkVRRWBa4+kso9gJuOA3NjuvNCU83DaIxDwJCenGeAQVK
GC94F7uIGEJ21eoHGK/WX9jM1D2AZEY6hs4pGmSowKJqENrGGq8kRowM0JrhSgw6
RkamvPoNr/l4dKvQLHZwcrkkyJ+y0A7eAOqU8VI/tC+hXA4sZY8bbSRuU7W/OV25
FJLtK7DtlJBS+h5GAFFiCCswfVVyAZKslG3OSgk5jRy1gEXMuWnUcWhwgZwhwY6y
FZQLq0AifbszJieCs6y8ZXHl71pUK1AWz3b/bVTtbwfudQEMe6wcgdTGbTT6FRbW
P/AIcHMccSQxHJcCENnXXlqscL6aMWQyvmMS1ORhfpvG6aA2uBY52H2u8A1erLSA
5pr0sNX8hr9sifzXFS4ihCBto/qSRO2y4bRYFw+Ucmc3FQmsIZCxWo0U1trteBJ4
Pq1ZwZPJZ/QJJEZbgkBdR1IkQU6KdK+FUKS6sh1S2TyENJgHV1LR3SCcyBBO/Tak
U1Ku8O4ToMVFPo10KB8lsXpkqznaDl2doDmq1GnqlISHHryoKc8m2Fa4JRlHFoDK
a/2+ux5xvtiDwNYbwoF1dN1jUeQJLKrZwVHgC8erH2rm7Y5gHFMHiLO6/3jnNjaQ
xze4LdV5hJ+p915oDKtiHJid8mf7OaMPqmVeylA6VlO5fzFMrb2m+D0hEdL2bSlC
PYGei918b947jTsYPcg8MCrX2yrhT79yjLClu1k6TVqh6p16RFaEZy+jw4+/fvn+
z9J+Yrt84P+3WZrStHb4PZKqLsKjw6ROR1pAGRUbJSXdfyttb6XNlmHlV91K3f03
lllN5DAE7LXSUDQwPE0bAx2z0gNrcUE8l0dNp7Uor/albyWPcf61AfZQNJ7Ch2wp
GWVi8t/O4XUURQha8WBOsVdOIeC1bgWI60QRsh+4AL+wBs6S+2DO9KG9FqzhI8nn
SfTTDLpJSdGslBLXeLJCO0gcqMMh2uSwC4tVmlNzU7POUyWtfXOi7jTgmQUO8nUq
nWr0rQ93AJ+FsSXzYG1CVKVwalAZawZI9ry3RdTX0qRRLixrARy5ZuGAyK3d9scR
EaH1o1xTsz2/iAF9TCXwnak98wcpLa9yMWxB6bPOtICZ3C/LfMZAMAySchtRnmgk
0BaE+5jN3IVRr4nMF03YvrUySQEKn3U/taThwqOQ/0S9QTtPTRtVbfS1s++R+UKf
XSmweEoUx7dh6fDYE4e18I4fdRK0HTutq/PnTJ9Nfd7hA0bJ6G4uCmykLlA4Hkry
++f83hmVIzi2aH59C2t95D2z9dDJTmvW0PzZeEn2m94LrhGTQCR/FVo5k503zctq
88ReRXvLvy1RspA0oPBXcrOnq99cLfCwn6BLoznhMrfEN/Tr3GwzVCQrnYwYG8g8
eK1ekfQi50inUtQnNIxbh1hJkuI2LARM2D/NIH7mgvscP74F0rzkfokCfK+8i992
CndMtvbxfc52cj5l38RHxkbU8YLEVXK/p+jUC8vCHbcwQDppiTg0OzFgxwNGOk5A
J+oVGpdWF5mJNwvDAkPrVASBNrbeJ6xQA7BkzxjdHeN54/bZaWqwOE9gBeNADnwP
CprFJutJQqc1HQJlaBwzXafMK5lDb/m63vRacmnSd0pHRkqVEy16+2cO2vqBOjnO
tlpDQDkssGvx1yYysVkL8WWI1kfqGEvHG0x0T0XB0OkTuvfiO3UFCbheWK8hQ3cs
v2hSSN7gnAfLQ65q9s25DiCBk7wVUn2W94BsCL6Po4s2o69W9GNpdayM/OCR3j5x
JlajwIgoaC3/S3cx/PGEFthHxwRFtqf6QCDVvWbWAS4WG8ZKTFkzfkCKs7QL1N4y
cwQwgEh26jpJdu+O0hted03rqptX4CkpUthaZHh7pvDhXgi5IvmGzxxEtS1HD9uH
LeTG9d0iChZILMgALdHG0eC85SGxov6DNUanOg2c8dXHT66kded+RtPBaGVAkwPL
kT52Qyc1D7Du/USvxPTBcezVur1RgCzWYnqNyrxZoJAfepV2Un56uRvQYMqfUpxm
E65WmkZVjMe8Yb26TAO9A2u9rcTrdFC4f0w2l1EujMC2XI5D1c2Zparb+hGUVibG
5nObYp2GkmhJOFI2TrqscJB5EbQe2yaTSFIfo86sXZvsHFXdLx4ypSoizWrw6WZK
+geA8IPyhJrTn7aYeXoM58pn/5txoUihXiSCEKBXi9Dh2Or7sK9p38/2cRvxpvUU
J2KYmqvmw1ixIkrPmDYxHWfMF2qjLxDeNJWgjqPBKCNUSlPWT15zWKdcDPVfF4tm
toRrH3Y3OuUg/krTJp9JqStNEiwQLOjWWD+7suhELIjVAyAKH1r/uCyJnvVUed0o
bduHROsg4WvRMbgX/IZqWKwd8nK/LN+HxWzL6a9JtosvrbkRP4b0QwLEKWG5AcG9
UyuKK+rUItg22frkkXzc6leyEVXazoH2V+44WAqUE7KvGRAaNSQ7fvnlX5Mofey+
MkdRz77ehCfiYDob2CRqPX/smi/X9KpYpg/s1JUz5CbtJb8u8jc+2C2vMDl0QHrF
r74hl5WsRBEwY7NEmJHeT4MdMh56ps/kriP0hScrvVA4drLiJYPq1nUGgQD9345J
ZfT80jDtoEPzb80i2/FWg4sCCxIPoaqDg1924wnIz2JE6wrRyIS3vGsHUHpDSJy9
o51ecAz8kCjP7T+dgP0/L3kv7s0ndCL3K99CzeIkRB9ZGePgo8XPYeRDx62/7mPi
q6M3eC0sSARF8LTk8sh/2S1t5yxFnadgIwNT5R5TVy4LCe66xJJdnEaBvolpabBk
MT0cfyWPk/B2/ZOHSduCJqf15QuTPqKRwhNzDe9EKSmBtTWTNSbIxZ8URnchBleb
pGSSX6m5TkBd0Plh+7RLwSVR+RcD9JL+lCHIClAztLSkZdHdsGbwLMX7LNiVZKYu
L8fbOTg5UniwL+06d4TI/q1bmDLFfE1iOKvK01dAtYAESlwg/hpjTs7Pqyi0UqP6
z65jVEPtSt5VN70AEddOc9wr97fArH2W4AwdvQf31lqzaCS9BubydHKsh/mxmssJ
anmzvtituxE0PZO+hu+8kzEjyzciINYnn+nnO/O31RIjRKUuHS0qhuA1M55r40hl
v1c4rrbob1Ey1HOGrAMOY0Ri6i/5cU3MWx25jSCuLzSLMM6bHJupcI1N3HfQ0/TM
nJMRPetGgAo9n08oPQYW7mInYrk/7miBjQqMXe5a//0dNsxstWVRuEtlaHqzoZtS
u0NxaacvsQ5HBKqfUa6+rsyqAKaF4rY7bR+0424v61kJq5KV960RxJURhk9IaKyL
0yGY8JsNf09PIu8u550ccK4JJ7vU366ajQj3IxpJDFu8QcRJ97CJbRKEstBai3cn
aaF3r37KaYPnC0eeqNRB1FLUnIxZ2f6zdMhyg7orow9rAAFO+7aVU/UTRWsjJdGa
9SkAhBryFaiKX89mNsBLck5wrgGuTm3Zh++oRPMbIkFmy1hIpya5yXMRbi0V7h9V
SNHzxdXMg5jgl3nIXMLEE+XUmBYAfaDmZb6ycDWTbxD209fgkfoaG0awnMuEIg2D
OLCrHdI3TndeNAUFvcPYiLu+sLnPc3CZ/CePAXHvpLYefOkvV0Q4+SBn+WOLcApb
C1NkJne5kalAtSKoUIyDR3zFm2xtL99aibGX7xR2F8mDK4vepOo3CwbMcJF2v1m5
BOgAS3q5dFn4GXv+ETNRyAI2nxStdmpzemx+ZHOS0tiVrpa3a+BK4nT7SSDnPb0z
sikoxGf0JWaXH/t/n9q8EoFDTKP7d0zacortZ4ZJSlPU9cfWYZwiA2pKavCzOeeB
dxZpzDlf1JRpMIfVg/YFGgTaeKEt6KnUYuIK5MNLK3v4eK85EAv1Or+ag0Ud8ffh
4dY+ZSR9z0wnKp3DJ9A4jzdeA6NUyRrAMSpc7IVp8xpMzpRDiDR9TEvlrtfN3e8o
0s3GEhtRgfCSw8qs43Cixijm/SlPA+kkW3XE6gfuVdR7AvZNudrd+fMS0h6YjBWs
5JMpVgyfBrkQuZC3t6wnIW/gDS1REHZYQiPAuLznrkEiT/Fh9LBGkLr6+m3KNrzO
qnwwRkAv0+TaJ6u8T868JNDYpZOINeLeDe6j9ultK8CW59crBlTr0a7ZW+m2iqzK
dVd5Ld2FvtXXM/OH3/QDeiSMXQ8GYm99gFDruvZKmTNLFPTY2mxm6nCx5BzDfuTz
AsQbPet8XsuACEi1kGpne5HCnKin1LKDjzFvfIEQ064qJLAuG+xWACgXzwvKzMQV
OWWhDjCJZ7p2MU5kxYm7BADAkibh4Z8lsdDYATBbwoSVBriFEJ+hMhPGEbi78Vf4
MtheUlqDGJbqkK7nS43E6XsWIHtSE/4xYqJqUL2m08sEdza6djwvybAL0G5It9me
CVwylTwObKfCdY4YqU4IejuTf56dtTIFT5Hhvno+ikdvTw4tHE9Zg6xIPmjOA4ye
yXtKf+GVaV+5mCp0x3b1S0cDh3S202KOShfSIy/Y68lN4H88SZxdbJu0lxCJ6pS2
2/YWiW/YJBjcxyLhu4mbJJPsEcr9UtwC4PpUE74AXU8VcuBV1ay3cCDub6hyM90a
ygpWseA8h29g7+CGfyg5FvSZMs/pmycrX7drtCtKRca+9Kj5EDHmeJFn/5FyO9G7
v2w6BR5dtePPCdZhuUMmyTqnJUZZ6OOkjkR0FFyfD5Ukb2LUtAjwxdWWJZtQ8mfy
ebZIk/+LfmOggofRismcLf9fRPR4RAUAmCjw+Akl5vV6zbA3i3JiwZqojG1aviLH
A2hn6fNsOQqil+I61GRtzBHsrQ1vJcb7qi60+MIXp5F2JNlahMDGiSwp8tiDWvGw
fZh+PB/2lRh2xy94eF8jgK8nbL3R85Gw59twB9eGs6mLGMjbEES9l41Sh3VVtwJx
zJ5IQPpBmseZa4nrpeZ6Xd9wQKuFd9pxiu2mGB8o5PlWM4czkgEl2JCctjPR+bAi
krPnRKrRZ7MUEmfm1kMJwjC3toHJG757AuIoTavmUid+ZUdTcaoU5F6ROeqt/7Yb
ZgYLzIKYm6BjxxuXbGjlZt2AMGND9HPOUVfc0Npq0EFU5+saqdyiam7u0xcwo9E+
a9ZlCVblhRn5nhNDt1soYkKBu/uRf2C0ZKJ5j9DRxKiOYen2G+j8nntx9vlwY+MY
g7/9KHaiFaAM23Dv1elXvHaHkEIdbj+M+htR94N57msYQ4lAyW4oCFbXJbcV6ZQm
JRccVmVc8Q6PbY6R23zFHOhGpnc+F48glVXjlfcXeCypB7dBD4frG+R0YeVhOpTk
swuWD9YTkThmzqD+AR1dIIO7lX+tBKCnbWDpT0XJkgUfscSXbbNrswCwfUerbJGI
W++Jrew/sbmszGPOZCpnpNJ/nvNXA4qaTFsznOp9TrHBndgosSyVFAWdvbzRYJb2
9h2vMUD1/dztrCHDF+W62q5vBOusArQy+hPtU7NZOUsIgXihBkkog/AzkhuiuYR5
s/ePw+YcIaFZYcd4HgnHNEoy/yDYaDLs6Y0PkTRVQKIjLvHaTGC7OFqO74l4+yN9
ntVVk78u1rzQF0lNWyrEpwCFXgjGOjSu7lB4QzDxeHtT/j/9USGqrD/JIQ5xpcm+
NR/2Bal2VmR3LUkZyjPwIMYzo7J/mz48/OMTaXDDtKtNFBKDSve/cXmxLnLIz5z8
lBc2CMhCGgUKp7SARwCnj1kob7vIAGIP28T20NK+28XaSUZs8qJ3dxfy4m9vM2nR
QaOBHcWqWBqehd2SaeLU8bkZDSGthHOWH405OKIDP3NYHUunKesmNie2+RDJNUJU
1EdN1S5w3lHa1Jov7s/Hc2cAPq5x8fXUz4osJiQBNJV6hDqF+KG41aqmxz/O0ZZt
IsnWM5pqU9v7RLqdF4gQ4vLxNG/6mvmQsVv2idds5034maISfYbeoIBE9ip5z5jy
4qDzbMfPC+IGBrOMyQgSAsOKjr8O3tscsGfWwh9DbgbLUHmDtpUbH/IWNDRtqdk/
kDQQRM6ydTmW848RWsztSf0fGlIrGAe+wSgv+o+D57sZl5m3Ovgj10KhXwGVxKuH
FWPb5fwu22Jg+E8SCwVblTRhH/uULfXiugUJRiucZEJkZJm2J3YfyiqdyrIfD5vR
jvNJt4950VkQNFwAAeHFqOZh03WpbOQOSFFdC8nlDgjcTr2PEpCoFEwVQjzODhqa
XO8qxsFrixQ0vo1qSJnBmEP+y5nw/TX2g4j357b1Rmxu5e2i1TksmTFfPIyo78pX
LzB8gBNh3HV+OhbEexp7KR27Otg5ThmKf+dGMZ0hpSgAnYayQUhWvr699bQ19eHa
B5k7TeWwcuMm2LQlmkQhmW8T4zDRcoNPkfSvlfudWjVlW6kt1Z75RPMHWnfC6VZ+
0vLj2hftYALSWz83UcQAC0tRSis5V+lSoPNEpzdeOu0+tArELmd0slT4rQZSn+jL
VeF1tOUfnZixWOCgJfV+z1WifEKs2ecvojntiLv2Ta/RiosnVyywhCZBLZl9v4f9
3/wY0N4psK4WXb0N3d+Hu5RR58gYSXP3ek5Boh3kudsYqah4e8p+999ezeIfh07h
dPYKkjNj0u0u1L3meW/tTvfFYByrUWtvnsZUN6NJ0UxGu8Wag7Mn/4pGsUB/WVov
IJC3Rfkofw+uHBAhFvxjK6+O76ccmINVkisIExnHzxwVQu6xBjuzanjYzvWSph2r
PLNbvRDMO4yiMGTqbDR/k4QhnzxfVL3AYAaANfDJ0ABI3L26NWWQafwUG3nBHt60
Lt90z51v8msUU3hL2bjix5ugFjJDOc1biba3wGzYuvi8dLd1ytBuDzfWWh+gaP7p
/umQky6piD8/pPSoNeuNzvVexmtXlQdxrkpJlxI8CxGTU8MRnqC7iG6rwtX36lWM
h0ZWd1MpJ5BeVZRSjmwiKCqSKGbyJYbTuOfGOrTQ6vkacJTDN7WkSOxYnFciqnjU
p2RM0qiBDGUcMPYQSNMgQP0ZKfCA7prZxffs8YLymgLKspq4nDZOvxCYW7Tp0kKa
eVUDWRIYEYsguO8qlzV6yNfooA1QuLZ0rwmr/P0MqBvRrk9S/GYC+iREOGhpL95N
Nmyt3xH7szOVe6IMjld0EY1dczOWs+xRDsgEDzxDJ7kaJXj+Ifcu1689/if7YXxZ
8wZJKPASlZ1ZHCrahGjkW4sda4aR2be3WIDjt05rYJeb68B2Ana3JXoHzAR/N9/j
faBN1aVHOhziGvlhrk5EDUGPZxAxeZEBQohU1gHWd2pp4C74SdD2m72v3GvpWzL8
RBYZGaeWh+n1ll+DszmSmP05M5JiA2Met0BlipIcSCW5yCQnsp92MoPGxO0DsGjq
k5LE4PM/N7UGLp6EhYx+iBRJES9CiWKsii9OOv5Joq71EV37Bsv91KcbH525T2g8
QOkiqCNUkzZJCc6xYTPCXIDtsbwhd9sEg1j5OFxHHhLLp4/tw8uRethxwtyDum63
cjm7mFX+4eEGYD6+astJSvc4F0UsyPRjeag+3vbEBeoU8UYxVYLER9At7laJQAKZ
eJGtcdZ5zFTc6oqB551F1LkYkeiqCZ05SArDYiXN1y14K47WlRjUwbzSjtug8UAV
/lZx6Rb43cwwEgfoIF9E7CnsJg6lOPWJbSE+I6Hl9BF2Y5US9zN+Px2FrLA5Qbdw
N/rrNAVZDxRgj+mluc/jBhXteIKy/TdSFXTIJA2PUcxbhqBXlpg3m2Wy3zjnTwKY
svdZY/4gw+l3lfIB2ZLr5odjp4us+is4Ye/mEH/DhYZcgpTkwdyClp5WmKuKSDn7
uH7Em1CqseRvfnofZfz2/PXNB3OoRZMo8h48XcRvYvR2NTCGDQrJSOp2WDLQ5flZ
q/DJUg966sVBmNnfnDfZUObZTAqqz5RJ1G7a+CxeoORqzS9Ie7QUne4kFD01CPD7
hZYg+cow8ZgKq+WWVJn258aMSmuY/b8YXq7xzvo3e8Dfm1um+IkpzYugkyhWXJ5H
KJDztDZwdlpItMNu85Vt7cR/J9v18yngWLI5+AQXxlIzrqYXCveRMCaKG5BfP8D3
fAXxLRXaioQqXFsP269QGhyciucDw9IprvUOljkTZiTK/KlHG67qVqVr/88rA5KJ
rQ+75mYr05b3FV/EvB9IJm8Uet2PRpxgyEZBbVZs2hIF3YBMKR10aasZ6X2Xk07w
VoGY8e4DoNNIW1pyMi3hLdh7Z7LUwrRGCLibsebhCLsrrWG/8Kpa0X/6k13qZ+d8
Q23KGyPcPXpogfKLIPZk2E13DFeC5439ek0oEEiwepPk+kilZadSKY8iEi8SCoo9
i3Gkl/r4+ElAMllGhBsdQwIwCqoltXReORWZ8o6iSW806ATg6NZXAhzJPpj4SR9m
+hY3lbzK9Kao2K6PnedrGnjP9BN0tO8LCGDGvG9IHXDjkevgypqXIy4x1lZFiy9S
4ur7ZSlF/zRzQO5K61w5tgTmhHmkeHXv9cKSnF222CxoOoacko/FIYK1F1enoj5g
o5KK6NInL7jySXXM1v3SR+E2S8J0zQ7xEAa/jYwZs2jKqQZreX+I1TOzuA2Yrf1h
iI1f3igMzMR0mY795Wzq5XV+oypmF3oVewg45wUT/bb2KoXBJGbbRIJFfXDVmBEL
cuFHWrvYJOROyKnEPm4KALUn3ix17pDaUlpkDLcADAVGCrx/3Bt31IPaD/WRX93i
hFqTvn18J3hRrxtYiFxW/hsYrCG9WaPxYtkg1mehV4hcEYJ5aiqpeANjcPUTW9W6
rlwwrTSPvj1kzwmF/Ca8qw05nNnetTWCU/kfZMz59wm+BVL/ZWRSyCLPbIEA9yhJ
ibNP61BLZxLgaaQeqEt6noZQcsm8TtQY58U6UwnJ5qKLnIz54RjgfdvF5+VX6ORt
e5Gykbv2e7K9Iajleyu/pAaDCQGeRsK30vvEC8TghhryCk6n2BjW9Cf0t4JFMmhV
qcrzYUE0QmDjBs8HghiXvwj3atuptCEOd6Sm2IwHsbRur96p62dS2Tdah9sQUuyz
oL86CaAp89XPDuri1xE3VA==
`protect END_PROTECTED
