`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYpshJ+Kjn7cx9LVbmeAPNz+iYHTA6K3RfUflfShT1BT6yP8STtWHVq5nJZuiXDR
3FY+16OwDmGWFiixugtbOp89MNrlcwLxoAywGph203hWmKDw6fcz41GPLxhNI+d+
gVfXPtqa3c1SE+tzCY8dT05xjfpGl8E8KNvrXdHiOP5o1efz9OBnoF0KcqahxqaU
ybRD97trjrJ5ixwAK3goztczDHbJI1vxbQQ8ys6+YRaWyWYMtc/4NOzFxlwLRQUe
ThycORwYzXdLEXSVMbVZ7w==
`protect END_PROTECTED
