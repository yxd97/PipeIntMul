`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fqlGbomxyavuBpKZ6KpawO2fAdBfjrozchLmM3L9p8qfNIfqRTyW7dYuYFZS40U
dX3Ecf5ymTvQ9oOhjQ5JH/rMwsZuQcE8iPVXSsCpp6ym4zJSn0y5IyzH+YWUgkiA
xV+Vc9OFiIdDJz54YFd3fMGsMywYiBkBVz2O2vjar7WxfsyC4FvIHFrf6vHRWfzQ
74vzjvrSm3x+P2B+QtGcXCBSjxBiz7LsZeVcFkF2uPkZsxNDbmlkleQgCOSYjw2P
`protect END_PROTECTED
