`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tUGKi5NgYszX4Rk8bacw32CuTqEInnjR0Oowgm8JvHdiQA2HkWqORgRLkEx+gChv
fL+s+nwwmER9g0K9RjOPaUDGR9Q2VnBswZB1EirO2ahH4HFQFWf1DgsqPsuXQ0JG
lo2IA0aNF53fAalEqx3SOhWGEjwjgyQPX73vCY7PLSsxFQI6fCQZJH63Pgj2az01
o2qkGWpPEgt/uojOpIxb5/x7wm3EFHJBk3dFBEq5AN+1Z7NVHNicV0SghfIVsfoq
3UCMTO48DkAv6Ly1M5oTPi55FmnOYLT8HvQXS5x2/ushj7GYQXg0+yvN91ejwhw+
YHWYjvTBaQz6fhUJ0DAPMZEwmKstMPKz6rRLLJOkcmimzdVkleDSvTPh2mOsmkPy
3BO/zU2xQgOWCcNt5n+iZwHJirzMyA2kPmkp7JSzG1/AZBtYKws6P6xzqDa4zp08
6+RsBdjjUgqysmgXXleMes2twROV5daHzO4LyIMSHcitnQrk3q64yWR4ulgMedDO
Z1ov7zG80zVlraQvXPqd0Q976Bd8U+sDuPeOTc4T4LJE9IRTJUMYbMfItov4cQWv
DnkiQmdZSV0gv2eG1mjT3Si8VR00oCF3yVT8QFHoJIrDJ05+m9mzWMdzzMNg8niF
q2hyT4lUPKuROhrj9XveCAdrg2k2wVuxJvbBLCeyFLRsfznBmAOLzrRUkt/O+sji
ywfQFj6HUnYsx5+lmcfpt7ycAX4uTLnM50082hL6kXkAlv4+7g6jVVf143RS0bNc
r7VueJ1lacmCJb/bWS0fQ3Zw3u8gCm4wiq+ITS2xHq1qUPc6F6YhWaS2F4SJRucz
nejbgOkrW0F/3PGCdOsa7o1EcAkArxrF7GmN4rQ5mQnOVXGigNFJYkpO1nil6mqi
zuRh6dHxuII5ygYFhLFWPX5krq4/96kwF91nYPXXLPj70C5bMDpFVKJ/vI3ofxU+
PPEP9Mv3xAtfBs6tFmCweIdlRGTrkeQSiAuvN8IhDsKAcbnSJgesZBR2J9XzYFl6
OdqY5a/hXVb53knOJPvWZ1A759DPByEho6abg8D2lCfQfiLASvqpnGnzeBXnPjTj
RD6YiLsGmd6W7Xe1ce8zT/T7T0FxJr4VWKwet4HqVcM1jHJCoq7yk6CiEF7if4zb
EhIxQcoy86q1FMqwNmdUprf40cSJmKSsPDIW2ERM79bzpC9w8C5hcLOHLO32aOVD
r+46hIKnVp4wEK9Tftu7tiH0oqnqHbXua0gVxFIXuK+Jb7jQ6/jBuIrW/YpSmhA2
oBhFYqejYEaLCKib60EfEczYQI1h1Jpb5tYuLlEi4PLbg8pYLeEsHpUPT/FRJQnG
F5x4F+cgSRIHt1J69/frbYhX4VIJE+ir3IDv1/KUZywDI5i/rfj7ARr0Spj2mMXa
yMJw5Iv95jlRwMal425TFAzyVBVtro0pG2aUT/fCbc4Fd9w6PXkFBoEBFH0QrPzW
PkObU+eVc9BvytsvqJSuxt1nL+pZlZlMBi+szp5FQXUFIkGTuWe2H4M4EV5ZzSG2
23rbX2S9svBASmOZKXSqSA2Hucaf75X8ml+2OC4XnN1eOd9NHnct5+LIGYUOHUum
rVcVtKlQjfJOR5I1D/JEf5hsB4VTHq/kdmQ2/oGLJJA/xT2H7PIyKXaTaqISi4AZ
oHHr0J0Ar4pArSFOx+9C2i7oi9VNDQVdb3k92kjLT18osZHeUGAfDAtA47OO+c0+
mD6Gu8hOQL3bDHIDfojg9TJ54aiGnbE7JSjkn5LiZiTTSVGRwR657+EjxSkC+ice
9eWceDa8GaGwJI8RYpUqJgS29RFmaUZ6QrU76+W3ZqWDw03M/rGfDu4fugpoYuu7
ulwgTKD21F7wzolIU4s7hwC66bQ7+VSwOrErVPskfCpcQg8lARI3KA4ne944dsfm
+oJTffnhuipcDFw6qudqErJhdt+9YVoDEueylzihX2xtGGUacIu7Xol2BNwYuWKU
VQyvcIKEWXyNRTQ4lw1RhubpOiqha9fAGMKAGay//BxdqmtrM+1vp02RmzBzVJhK
ZybMC1Gu4ijuO4ESmzuk4fHe3Uu7sGdgcZLiu7BcEiErJ5V3lSrpycJOsBchOuvJ
ynuDBhoZuQatWRd7XY2WnGckp9r/Tu6NAxRG5q+ZRnupF57aR2Yc4vuP6LCE3DfI
CpZSOZpdLDXNSb9H285dC8gqEYCToaVQXsnt1LMNzglvO9NZghkRNdLtYWI7dJoF
PlleI81+ml/ZliVOEzIN2eIdFatP3b7905Ussf6n+8zeIW2+Zy5PJnJj69MEAlzf
8+EnPaqqDl/xhjHuD6/yUzyc4UJ05rnSIFHFoBBHS9ksaayRg8OC2LlGw/IwZ2yR
zw6onMdCcaggJp6n2zuE3BC3RWqkWwvzFMkaMSRXQDMwNaXHQeR5h4rS3SbHsjnt
UdDPr18H48GI57+DrtCxByUqT16T5ERYjTHREQk3x15QNWYfeWPpfJUjw2oifnkJ
ZX5NC+b8QQDXsTHAQb5y0i0JAm+uXfHRCA8RmBpOJM7etUX5JmjBOAxE2/TiOJQl
4f9TORzpYwAB0I6Lj1Knmhpd9zndVtUMXCPHgvj7pWAl7F2Uxg0aVYgLlxY8Ya2X
RLzvjjhSbFyMbwSh4p1ah6C/5pgV1V3I334tm0B2jMbrZcJEx2WAXYeXCIvmBkLF
e6SFYPWCBu30uES6a9viSfWPjYaEBU2cXg7IqbcNC1x7VGD9evRp2DSZ1Diyzdw8
RbAm6at1aqGeROT73rr8g/w7I2Ww4l5A6kj0dvD0iv3CR/p1Rk7vveM/SB8J5HRu
TpVk4omGs/Wi3bezCNhFNr5+3RPNdOrbRh5geoF4iBD+VvWxPgyiuUYaVxWkDDFL
IlOyV7raxbDIahChZJGsXI3P49HeQEJ2sdJ6ca/E6ELpIbfx4NGNP79VM2KdcZAx
jah2imKF7PjmyqkeeZge8YhGjNVXkbM7VPSqztXCP3d2R1pYqSv9MQcP/fxfeCCt
G0qXFqVytUy8bi88Luq2U8mC6gl7iLlN0MxcaR3u6N7IKMFOLrBthZLYHdDDvNWE
+p2LSgt3JuzbuxDmIgsFBSdJsz6w9V6JGwSNupjwmUI69/1TST8+KH+whZ4V0Gyp
SP1jkUnNAGhNBSmDlqIxC1dBwzGhYHLepZH62JCeG/r8NYK1/NxHY/HUdnyuXyBF
f/R43fCrw/veQL1yqqanm09UXsGPSUZQu77g/MOurLC3i94WT7mrL2wyEoiuB4wh
S0FXUj/cSib0PEveWbpsi3JdZ60fm/mV6yaDU4P0x9ZCkK72wKHiU3snuvKbq88V
WKbpLQq2rVOeU9nhzYhnGwxBtEgg8yi82du0dTApIBq7wVAcQ8daqkbFgmJ0zDRI
Q/7R4BTfaHzxzchu139lDHf7Z19AfmR6xNP9J3V92/ipS76uL7ymu1d98siYhDi1
+wKdlQRHvfhIERfIFcWnG+XxVF6eXGE+TnNt1WJUULEQlKoPLGIoWf/iyu+Mq6NT
9Kz/5ebiV5f30ShmvNZXmXXFG+SXgh1+c9UO68rfS4Dpx6U17VVjIn57PdnfHnL0
cOeCJMI/ujys+FkmPM8w+ZYerHL/IsZJoKWFHQX5MMQftKynpvpg0C+D11tUlG5O
T4tZTECgeZqJydnAvhmVsli8IYpCQslNmS7SBsEmsFCpGqkbNIjYb6btegU4WBFr
b+byW3tgunFz7LeJAsAG6F/oc60yWNmrkZq8Kt+Eg303rVl9pPppUqpoNJOvQsTy
YZODCADg+a7Q24WfHX/gSEY1nNfLTpSruLZvmgHKpr5e4Snw7QIIIEYJhXcdHMeo
Ba9UwnaKvlcWPfnBygLcami5Jw/skMC8t4oNZ+L4ZOmW/b82au5y3w6o3jFxCdmR
uYGDeobitgQgRuiOFWbXfLngvSqoJ8u6fdSTZjZ6uR5EQ8JqjpnwmnXvN6WPM+KT
50a730KwvYGlq9RsIlH/vrhmYVcVHq/ev5TRfZ8+Gbm6MsgGpF+gcyFrXVvSrbGk
FhjKO7tGCHMTIS/ix1be3h4BfBdTyoot1wKuyefPMHv6rMl1eJAcc4UzmcjnCtUX
jw5ztaEwwkXtrR1OLm3XLJaXwCX5QLpPPbC6t9LuvNGtNptnVcnPdgUGvvWyXT9I
ykTmXNIxTWnNYO6RCQ1/fsixMMIUNXkG/rdlUmgw7//exeQMvB0TPtMqbBlY3tM0
oil4AbRzgs6k+SevTA5Y2mruK/oO0YncUjLfYZ9L0+bFq31N9G8k6GBb7/8oxEjV
RAiZ6eq6ZJT9u0QSiYRifrfKigMJFKl8pTI9SPLUkdNy3f/3H2l6XIeKwm9Ei1Wm
qKHlN2FI9MKI4CYGI90u6YlHkGsyR7aIZ/G+MOpcP7nTYi2kmt6AhKRHAQ5i2Vl4
OUhfY4QkcgLkgriTJLjlHAU8zMxIQALJ+veP2lUot3ACKmCKrQ5SfCUvwpdpoyo8
hAomDAqMg1N41xdAmKp0sQ6B7+oETsFoZtMR6X3/3IP5SFPWqDJQJpLGyp7UIobF
9oMs8/8767tTnHsgB0SuevPdH5CW6g6nTTA2a73KFwiSicw+UaPMX2z0tCN7HAQk
Gt9v+DqK3US2eCVY78Q46wykUJKxbbwkYJmExzpDKDoORZAwbYGLEFrLJxrsSB4c
xUkNDiYOzb3VrnSAdhUktpGV96H6ezCSwd9IxYguQO7TASSWjmdBqWXQWhJ5q8gw
b0blsErgImb+MksOD42gFl5OaLoUtSrO3kFCpQaIOFIqBRSBLGcRmvw3xIoEq2vn
h6Aenky36P3jXTAamaqV/Uj08nBpuSstdvSvcjZLdh8YDmNMDre0+acZ1kZbti6r
Z993TDbdSBIxy/tztjEG2mLMe9fVHNv2lsCAxiDoT5yBMjSXQwCvQnn+VB+Nkceu
umIKEN3ZeyJKEeMZb9xIF3ImQJ2KU3dHUFQ/3cE8SbSEy48sI+LkkZ4dk+NXlGpV
CjRxsybLt3w9CtYlSdSbl4YjF/Qsweo32eI5h5Pgt1qBGttp6DGL+NBMWGj1Ycv5
qzvRzSSkT6bYfkJV0rq/h4ZOfqg8JxMGK7p7q42Tf1SmFwRyLiyGOjdTEyE5b3ru
WmE9eZRxWfn6ijgWYWgdDv+g2LLy9UiOwP5ZFUhIcLSB/JuRrf4OVR0fwTQtPxCe
BeMAdarlSqIl7/ZPiyBoj+DhTVu7KIVs0RGdB7K/vPUlFIU7KTjUJ53yGJUhacGs
bkiSmf15RCnD1oZwuBmm6md4cyLfpPtKYiny/70dhgnLWi4w6SiwfOp5ESClKGn8
CvxkMWOw58A33ZpnHnRjC2nwZuzDfm8Q965bq/0httaIt6aGyvB9ikkRT3gbhI6l
w8AmJ2taYeAIqPWK6tAVVxqCa0QxhVYfyr3FFwkIcCtJjA+Vmr2N74Ay4EIDI+kO
2WUSdEvdMAaRm1Ce89uY81L2P/JRAem+PwINGkb32t0FPj4rRjakGAtNRYQzUwrc
j7WHw5Dojl8+xLNvMQeQoVXP0YlBzUviF4Uzx7+jBRXVS6LBGsE5fDfv/yQcS8zI
OUjrEPeLXQSIHaBlyskGViwGp63LoBRiJZ56K3LmokYZ/3nhmZQktZSY5MsQKqsD
5ZNxwxqMetOZHXi+QzYSDqvkgLkNb3TMpHQBrOh0laZ04Tux4iERjqxic4gwi12M
XSK7xswzR1KIXyVo8Y+gB56B9U6uEeq5CrXl96C+cYrkS+j9GSap7Q6KLjZHAM+u
yT86vCdfOKu6cep6WC0kIqnjaANzd2LwkC/+vw4AQ9I3Y+1a6q3CZUX8lADBkamw
nFm0ANEIheqlvICq+8InGMFwqRPSjybBXA6wWIG/XX821gE2dB4JsnqP9RTZUcDq
qwtVi7XhnshWHlVenmzPR2gtv1tXaTgThTXp5Y5D5gLzq6As+ObBlpf+u4Br0kud
Jfloa96qm3WaGZfWITmMPepE78VRWma0kL7o5pa396XW3qZSKKb17OnKPOGJxai2
Qg4nNsYsCTKa0eVq73neq5aPXT3ChHSQ9A1MDEKlOPU4S06RMdCaiZKFxXWMtAR7
2b/V2eHzj1567rtJjlAd/PvDhOY3Zo5wjcOkd4uvCFy2+wkOdxRcZHAJWEpz7mvj
yQB00kVGxL90++tCYeVSpmsAcEQCwjXjH+Ak8XvmGGEjgccqivwI2jwtCLGfHPEx
DOlb+mp0RCRec0wB/Td2U1GcGv1c9u8qAOBpfX2FmYEzhhQ9pm2aM5nWtPkEplRp
EBYUJP9uUxhjh6b1DJnMYrVy7c6XfNK1VbiuFMcrf10zoZVHGTVsfHFOWTGsDvY3
RtmVBmXIoSlt4x9qT2nwE2Si9f3i/VREeNIxvikEinvOXkzaV3KKQ671lG9T22pp
3YS6/QIjlEu9BLX8cO1/gGyN4Gq0OQmiSJ7SPnQPPuBLBRSzjp7mEv10UsXMnUzC
SKay/byFBmBFpFldn9jok8nf8B0tFoNcPYu3gfyeZP0i/zSyfDvaGfNwPAFkVDvM
oSc496OMPTGQ/3htWr8qh5hnYWuR/xZhB4ne9xn3io8GvK059fjw8VT0RFUnaRfW
PhgJvfNQYMD5570IDG6GB7iMI5wxSQpJF6DEO1jduOtEsHy3j6KMz3tVBSrpxru9
H5BYKmEdVbAZ/K1RilsZrM2zF6prge+tV59m/pZIgJTgPMBar1s1kuZPkniRmPPg
vNL1PjVKe7Qk/G7dYmLTWVc0D75fgoqEIwDUqDxPPTDsXY31B0/FrsEZsm83arMm
FQ1TeqUY5A686KyUYwZmCgvEASn9gYF+QCaQr96x550yiNQb4Wc2BxI9XFIM/bg5
gD+KSX+4JdYc84T00+YcZWb5jZVV6UvAoEfSwfT+k/7ml0HcLVSq3huJKh+RvY45
de3kRS/BzM5Ay6tc/MXdoEUEvN0af5YyBbr0E49+jLqM2k43p9JkdwECtoILCZ2l
rOqnf0bXB9e8nvBxY1OjmM1/ZniHzpM5s2I5ZY6AAua03gDK6jvdc0nbfQaK9k7+
Br8F5X9UxEO0MmIFT/rkpLpoXOdjjXVklqmE7IMri3ZJ1+9negRbsb96mGMOkfdx
+ZrlXnov87xscMq8ktwCoxaKA3apvhu6VcQN22J5dOISeUgUsdSnlxHN15Y9mTuz
6Th90LzkHjjoxELu6uvUEhbqsvVxaTMqyQ8lBP7BfjQo6NmvfmtvaRSjDvyQNzfe
RAJ9pA+CLF7odYfjZZCRPy+6+CYkjdccVJjA0kFYLWgHcob2IMJGjwhv1QS6WepE
8ROZQrr79YeMYnRx2H7qcTUhkBo0pdrYoWISJdIw3JZKMkizlYt1oD6v63PAMIJZ
P+4JDgSNFU/ESQI6mhFMkObrvZHP45UtqAB8bH/1gQsPzsYQnrT0LuFmuVtr/qPI
TUd1jxxO/TM1bK9QJICgbOn+ktT4dYOACl2yGV6R0m5H4pi7Nu8wbPLIgZHiuNZl
LOIjv3oqI2LxNYADDPynI0B6jx4CaT2AlNjkOFqjdY4kqpm59zuGxvvL+iSRuO0e
bKXb2Q/g6DKURwV3lvcLYQBbp2bPzVoqI633GFuiIrapmodINfHzsmxnKp2mpy/Q
xKCVyyJp5RwkeyHkj1oinzd2crFymwX8g5/Arxfm2H4DqgYegvnH+/NlAqRbaIP0
Jc9fOzH7GuNMnHXx27TKsaSHqReDu8ol6KA+kkjnaA1FwoC7+gg8w/NWXA1mm76B
OkFwzlmGzFy75L/kFAiEyq+/w1ybxkVeWUPtV17dlMDeiyGzduO217kQZEmHSwmF
fRVHDNEtIzX2JVI3RXBeoCygoOM3VoBT2pcoBtGEv1kcPtH1IaQ5VZSdnyaFi9Nz
03Q+zhpZtMgC/WcSXpOjiHRv61XNRJZcPEoil849p/Ul/GOWRE/6N4Z6mrGn6NXR
jLX2ZZtg4LocwPuYraSSQcYly3oiYGTP6NnUZC9BZ+HOfdcj18ZS/u4kz+9Q4F8W
hxyEFyuO8cQWDsg2+/FfXcQHWCGnY/djtdpnX4GVQ0OzQXJS6jmvWmUTEYxx+HhW
bo//l3PO+xLiCmIXlyK0D8xOZB29ovKx09vDpkKlikBD0qw2sF9Xg42Pg02Db55P
UEz5vzYUmZCruDsn9sKpsCkyp/MxNL6qMbTUcPY4DXkUWIH6Qvw2hGM/FZOQnYTh
Tr4GIMsLakHGGMZIG03RIAIbW6K+afH+3T6lU6OkdQtI/6L3KEN7i9pOXH0+0ygM
jol1l+IV8Mej8Fw3npzQqwGgAoBbzgDsUD2o8cuhJCIwKHApPnRyc5seFR6Q26zH
i9Uz/SeoN6PIMu/J52t/+6Bl+uIU21kqnLiOsa/cxrvpHxnWjznjINfnXmHBYtNv
e2i7jQT7z8daNqxPXtvgkYmdpuCSiGwQQsHWJnsP5PujGYNeT5Tx8KIJr8It5ag9
tnH4Bc+DT+8Krm6aIQbEvMVFSQFCjGjsF0GWLKHtkqqPCpWV8Tg3QQwNi1IsxWIM
LcdrnoI0NzB1NOHt8SejQbaf05QPlMu9tpHqOlsxmsUOQqWVtCOEMxYvyh35hFOp
Kz48CXIpy5RNp1ms10uAKW/puqdSzruyaKAObqZ+tanjboe0L1v4E/lTv8CiHGIa
OdVutkp0hdBr8iVibo5qNfG7i10+vFbDbZdk1+FzSPYMgiEtbPESbFsBe0PqXY6N
JU1yGGMjCdMGNu32/nIb5XuTMTImKntHm/Gkqo/N8FzXkDyb+plOYl5Fl4h0O+cM
CUIqUkRNgSjhVMlp2AMfZTl3fiaTqa5rgfVmwU0sRygVrcnkS+1lESaOkotKgwu4
WIpOTi868165PSSEXKXFFk3biNbzAsheT0xtjdbkfXhKYKffbPi0DyQpQQSYYclV
E/lpJealyHFvOdzpJ2fnah+1ANQu6d23I03jU5EkHeml5ehiaXj8yrxM1oYcePiv
SnaMl+XX5AZFrHBg82g4y2M3L2t/lC0Jwn6qyqBhQsxaOI+INo+r/Wd1FdM+IpVU
8WSaVRKIU/KsryIwnkq/hXpMLByYX0cmUhkD4irGmLlmr7MIqn+S9m6SW0ZI/w8t
kL4rlDO2MfTMoLs0u2U6YuCcRJkOH7FLmpA0jnLN4kv+XX5bCrcpESYn8axHgS2U
Rwg3xq2wAzDkb6au2CgipJyMvVwW5tCAYUfr8XFcSzYv9DioDXb+a6NlKQ5rwNCx
9ddxulvN/VfjP58MIGbO0AhCFaHtfAqNaBTayGRABIMJ7lbPO7u59CecB/xVCrD9
JeyjykZvxIzBpRloRQHijtUHAdiYb5/0PVGojqidvxBTL6bxx0IaPZxAY+XBwraB
oWkI5f17lqh06Wrmyd/zIh44AvF05h1NoVLwod0+9cco1Qdm9SagbJaUVSpRQ+wb
HRKeKZ6VOyRQqAkgiHkW+IBnFpd90eLu5v/nGIeaPhRIYeWEDVjkvUAZGPzF/IKi
Sl0rKJuTpz15s71FtAe8Qp8LoMBpoUKFCZAF38TOXpnTiXcH/x2ThttjxIxBZIlb
CvgEjwnseUHwxu5wVa3DloiyHFBYCIjEvMI1DMzJyrhdrMVJs49SqUmXUtBLbrXu
r7ip5rkHcnp3rJ/97aW4CTWbGxrYXvQRFwyruDQkaC8tM3fGOiwSk++b3zoqMuh6
260ukpw2vt5LpZtMGvTfQGQVcPxedrsOC4ZSlmKVRG4WKTxvsghjOXtQPqaeL38V
kD0eyQjQy2lwMCrBjq4sDfXRSWkCSFbelpu2gyNlArjX5YxMMKIIqvhxkm8molnr
vxN4AznfNsfXhvL4Ronf1pzWM3F98j2ARf24djU9gjoUyu1/cyT14WaQ5xEIwAuj
wiQGX8srkoYMcwnhH/hXnyjo1R3iG5dJLWP8X7Mo2LRBT/4VdMpp3grKAME2c6Py
7oq4BS2nLOpO04W2tuBCwsvcu1y6QOd8R4q9Gatj2f/5tWsRApMvOesJLfC7DKNf
H0ijCI+MeJ/kLxWw+ixouCl7nLkwLgAjT2tHQtQSFHWCqa/T+V9jR5tlPDi1x2Hz
TrixFhOKJpdWGQfLdWvBQrYuQ2e0R3BsWTJva1g4t457TNs6BARl228Ymv84FGfH
sxzZ9f1mvKJnnmOSLXllRZo0Hpt5ekTmLiwDg/PDdkrkT4WVu4drQxNYuoQfoHP5
FhCqXhdzGk+b+BJXhQSL8xIlajUL7xX9RWoD4IfE28NY/VS3Du2xWB66PXI+OsIV
ncn7+nR6bkG8TmQDFwoJBdIy2o7nf2GSjN5UbZOF4so4TlgI1auSSlUb48KkymWT
fAfX8BQqDZr4x3/I+OcptpI5UI7i1wpw+/EmJJwaprNZQEYMVfiqAR90lW2N+WAi
QKbWVNV9RaWqqUzUyUMuu/KSlgRo1mARgugts4mnD8gXjEywLzlyZ8NNlLNFKAHB
qouaS8Bp77Buj/baVja+0HLbV3gAfw4RqvrZMfjlKohKR6+wqknTAVctFoMMYgV4
9Vykg6nmMc5BXyAqcoLB5JAMHQMMi0an695Uv+2sUvEE+lzVQmDJy9Ra8kRDFn6q
uNzCZJqMVLaAU8tsuyWepgpIsuBNagI5WXWtoqtmsDQ1owoajeHlqf8uzjDYMWb/
0OpZphlrie5NWxVx9QA2oCoRVPmiC+kHQf+iut6hhP+WHwcI/dbFdJTzZGxQKOg5
Zu2FvNpmYkJCIo9lgJFbcj9sJQ/KHqNuEhOFYrvbZZ6yzdGam5HS2cdqIjshqCaq
BZzsTxie5eVckXvGnfdRihKUwwyB2ACZAq0Tl+xPExdNDQbXe0PBb2mdkrb0vEek
K+Kc+Omu7mkKI/rZmVxq7Om1j2KhLtlHV9fHsxRObY9CBmIAB7DPdRVZwiY6oKAD
ffSiw3sA7tPLHp0YyI2ZK+Rb73kB9WnxA8QeJXFDEJg4e97T+pjdzpWF6lh3Jgr6
Fmc5vMhAiauw4dfAQU7uzHutTK56+PLSi1VY0G7c08FhEzNGvjgK7wjugtQXpWez
Rk7FsWztsqG+5/D87IFBTfkkQw5B1ZQPClAOIlw2x+Tmq0ArulQIjcmV60WgZQ4I
IGgTyOpEvvFnCbMCroxeHimE9hNn6lSbSRzdgOulm5WbD8AW3KrC9NL9QA2mftKp
Di/MdAjy3y6bvmMrhajPtAC9c8RMEJ0ebOLNyTE44WQIxqZreHtOXIH2rFHqP+ZC
p5WR9yw6hPVCWm5Oo7E4qDYi+t0AOO0ypfFYbN9sSxF0WjwPqbc/kvAcEBV5/BlR
C+gETON9ffpLJvqVH/hzfv67VIZci7RgAhibcIA6JcXKC/7ldBphrQus4+MY6OGL
3M0Z590pyEPwOUWEE06JEWi+WRUdhQciOyNgtcAJy+Q/FOyCHI8ZAx8OgzREN487
5lhbHiTibFK/qn5ojMxxZl0EZ2t2IyfaFWTyMTpYmvxfMAqeAFKs1yVllrIvRdw8
Oo4r0DRHcr9HrS1BaHluIedwf+8kMbtHwRrVyNURbkoxUD9vfpzywNXvJb09pmpv
7idYBIC0q+lAVaW6YMIKPnSQhf0Q4fEh5j6avomJGCsbrBpBI1oOWmz/raFzLjsU
PvaEx+OhgJDYxNmkKlEiVOM/u2fiphvtndrutrDnT8VmXGqnBIy3zTB7jykQ6ir0
bQg7wwJPVh5nNpNYF7r7ehNxIHOsQQcrYeyS6h81F29fM4zcrtptSmS3HlzWSPnT
TDqwpcXWAkSsnwCG3HyZTMy/sVmmucJi2qMBMsj1e30M3o11OTkZfTJf6Ojc8hjd
m7WaDOWte+lw3jtzmvxJS4DK2N6WTox7AL5+W273sf2YVnEVZA61Nz9aRnEACMdJ
xQ/+R82swyk5GifpYYeg0GVXAZC/UC2q+1d6jXi+x/OsPUXy6MVi1jTwyt+NoaTo
GVycpCxSCBlGvB7TDogetsWmZlidmTa99oLB5nXxQsaieVJL1p2EL/XFJvImPyZa
a/7ehjcZ9/2/sB8NHqzGc3XUj1DCVL262Xjp4iWc6OHE2ZCmGvejhxiWye6HjF1G
a5BiaLp4lKYsxJFRwKVycmZmKQGQTaLm7td6p9zG5fPVWuKx0Q/lW4m9/tCfufd3
jqpCtKZkQ9ccvRiF5dzierTa6Kd0O5WemtX7ye8ywncDksQ+gUWoQvzDUWgHCv7K
JKoq2C0qVM55vVPnrbULMe4wTlUwJ589HHFe3bzVLaDKm+pAeCfdj/S38lSQDuWG
jlw6n3Nb5XZyLq4zUbtM6oEmlhuu6k/Qo4CjbcmqpvHPWKhRs69fr5J0KhrhsF92
n9kt5jAGtivutwHcUIcPEpaHwVVv5K0Zu4/JPXwA/0urBfy2jnq/usEihf9rtkZg
jrF/0RDzGLgv+r+R2lM+AUtFZpMWeuPaYwrWSraAO3Yv3/AIOWlOBrQylBkumTVl
M+Yu0YYWO5dQw3mUxwAbP2WwsdseVKWL18N1j2WZgoMp2v3xUsdMMPSF7n5shkRH
RT7fmo8YxeXA/rd4pGhxbkkUI2vRuyess9p+xl/UXm+UnN/KxVgX5PnakbY3xgCv
zjLUqT1TY9bJdkyi06QI+9PP1545hcxy2no3hBqM+R9tCHXh6e7+mrrOwCtuGBGl
B7EHz1RBddyQppGklZI681c14r1i+XCjBX6ifpwSldCXCpEfkZswx++txBKccHha
3+K/KHmxk/XV0tnEDgkkimmTyDNUZp/dpSNNF3WIuAd+4gr9YxT8Rto5vmekDtQl
2jShkMoOo2pA9i38KTtGyPdbASwatPP2einbPBauendrtTkmX7ZDfN3ucheRFJE8
0EigRAzSHFK6GkxqDd2kC08HEsCxQ43pVbcoQvt645+KtO0krlb7vjXQOPUc1i8Z
UGiftWNmmd5CQOBuKgM5QcMjMiCwJJvZo/HY6HPfM+tmTjwGe4NezIJbpGyh+MdJ
pd+RnH2C3U06zVHrw4f5jwRofY3LjelGO3YDETOhkODSD58Yfi6MdHATFNFlnZsp
x44HGT5xswvsKoZ/6Ko9A5frz6XY3Pv9hc+BlSKcZlXolCWQ3F4lDe+rkIEILwPW
dennL2AllTb5/sUZrKbGJjzjlz2GwDhYDFmXatiyWxKfQf4XYVqgkyFNRd2WgNqi
dDP5/ok5SF0PRlZqa6qmn5uZ1uNu+EKSd0lTSG+LKKjqgf9qQ3X0S7cY5R69b9WE
RU5RRyiejN11cXIA2XKbm7q9qJXIdt+K3M1/TodVEy1M+Fm8uqaXFStSqjXk4tM9
YEZ5NSN8W6PTsO1wwenwkuSQhYw1AxVUQQGs+qiwCM2rNsnPoR0+4f/mEGRZIaeb
ukxCS+kd3iBtKbPTAws4cgjCwLneN6la3vgJWiGyx1SFHPi11CWkgxorUpqAHUad
1Vc7NlFvlixBFSJ1Fm5G8uOQGUfdIV2ktX8hMJItM+Fg1mkfN/boQh0qJpU+dLcW
aF83RihMEITFYB6r4aa8GAVV9VkcmpnzyowudHYjTouTHwFjaE/YRfwlCl3YhHUl
LSZXgu9jF8DGXe6bJiwhlWD9gWZo3SeuNWZfdJvS6j+S+nDGs98D8lGa8pLV+Fa+
Kc/Khm1dBl5du4N2jAhmAZVmRzHb8r+RWV/xA60+KDjsWk2e9fX3o4PV3lbMkQFU
A9wiFX7rPdLKz3Iin3WUOfdkfDeNUT5EyhqHNIwRTr6W0SPYWedweMGDqWfy6lTj
QtDCfCedzYuQr0H/82nNnV5H/xaend9MZmIRQMxWeG9pRYE6nfuPr9V/HdqaMCwY
/8u7x+1zgdF640v8OdoodGkrpFMezOoDfdb8OQSKGpkhMvrd9QuDt1hrNnOM10wW
6maIrYdnISaF2iYvO/INGphxMWqZjP4ekdlwMCJs3LRm1c8jNvWwIRkRx+QdQN3L
YIsTp0WxAKbgAyoBnPaSTJU+TuYXr2iBNy3PV2Rtkf3Tq98uCGWRFFjmyePPFySe
w6EjurCEi4vBP5vr+KWZUGIFVFaxkIJkxXobWPB4qAavnXJZcIsNLc2oXR0qzi1N
wqt5/3FRmfJ50MHn3T895eTkz4+An+8eOJSLDGhImQ88nV7ZT5I7pS10Zst1vI7r
YkWS1qpwM1IlDlUCZ5WmVOUXwLf4fo4WzEmvs/tu9D+ZZimyEOBh4HC3us1FKh5g
Zg3NzfMUGd5ORddi5Y0tSfGQ+NxxNuuqfj36zZ9j1g0u9y44uNaP6zxmnFgck8iz
UrWQUF3/en9wb1B1Dskf/AjzVFttlo8p98SbRY0pFIAUQX8Mxq+gRn13G5gLbdVf
JwcrIQdEDRPIprIFxpRdjBlSIz+rzCtLzeRCn1xkwfvCb8TyQEwHuC6rvSwXaWXA
GodVF89T1P1syTgVUnlZjcgK5z5/ynzOaL+zHdwjucAyjPjDlon8a7DgcaiOfkAi
CyjI4y+kvN5fdu/mqoutFyFkCXHJCAvPHgOdXN1rCrjHlo1Ks8m2mW6TjhsZgohZ
sbpyDmBXcfpe9gpEHPLwneLvxmxirq4hOgZxW+dbLHCQ/ejHWitUlbckSnbwBn49
mggpDPARHEBUQUMIbyffNjyVpwkpohePbvanPdDEDNRSfijPFihHjylDX4xA18wz
KeJ3pNlVfC6C0x8Y6nfoqIqPjxcpFMb506te34tPGKAQePjsFgHohbl/IVVioKKv
nLXUhqeWwgQX6R83SWnXImaZHHAJajW7w9YHVGaPxirVXxYq1iBg+zbww93QiqFE
KXNb/GIPLaN4GRX9lcIac3F8fk4dKatEMjpV0LNsplpIW5ntVTBWuchzQDbq/e6p
vJbKEJnWUlS1LsI5ZusPdaaq6T09knY8zH3SLOEoX7C8U5EMpJZrkg+1fC/Mw7pt
zYDr9UVL/3lVL2aJvvQw5EFAL9+fhoIJvwpm0AFyp0BEe4eJQNuCHj564digPluR
D9NJUd9mx8GOE9k/CJ47prxsPD5ScAICEWqR8EjQs4Ip/iMbSX5YrF2rKAoXlNoj
GWAmddu4AenHjx+pDq2BTf70svi+x7kJ8UmIX1Zn3B2u1eQ6lCzqp2ZaEcGVkwRF
N3c85UdUbd0T+ps1pYWhYDmVtwU7aqiBh/qcjOwvc4paGhMyccwI+2Vf5JIk0MLa
1IBRCsjJfR3z+a1RaHyGTeNz9h0cYfQW+pY5/y5Vd80l+5GuZ6r1biDYd0VBh8+i
bl6GnCutsTou6WfnMBugPY/WpZsRlPi7S2ibJO0ZM0M/58W58SmXJgWxZrNAgml+
t7fPk2PZMXt8l+EkFVK5KAtBMLPx0t8klsaMTk1tBhicbfftX5sshZ4liaJF9Oay
6V3Jy1VvSo7jiJNJD6k+aFgDXC4TSCDQvLQ4vy1rfoCfKQUXO05gDT9EwGefZ3vj
+PUdKDwFj/Vwlad7qNiR1ePYh4jJEC+RtFuNRaP+VSdAkcC9Vdw7ULHSQ2RRqUNF
6KK6Q5Bh+0PqywmSCwtqA/5sFHw1sa5vm+AZMX8sDaotO1M/c2L6nIS08R5K6zah
8IzzNDwOhqqCwphGpNAbwfSB4TFMGNowucuQmIIropoS6qrrhxaz19Az8Uf0vZOG
v9tuVaI+6GHboRWkc+h0pEhSxHv1LCfrG/DzsBAkPX2+UPVyEg6bG0cNY7rIDlW2
lovXgAjVhf18as5mmeuRrgyXOcLde+Qgy33vWmN5W0DhVgubeakOGU+3fR4Zk28q
dI2lhRgpDSrF29mH4Z9Qd1vcu38fcsiDjiVmcVtHNFzRLAdp9m9BTFdyeryYQCtY
ap4nxPPIBWkEC1TLvi7Yzx7/m0wTa8Q8WZpzeW7qHWJOg/fwCToZ63pZaFQCx6T2
CDiw6T8y6CZ4UGlkMEqq40VnewDyXMKlCydIqHcNLNmlrQZ9ZVpwUVSAtytY2mE8
BROYZB/NJ97UfHFfS6xH5+ZysajanzCFA59UZfdivc9o3FhUldaF7POv65sXnJdR
VY6tQeifxohPFaftCU8zUpiJ+53sU3Th20rw8U5gDwaMN0QjzWP0slDIwXTd8XaI
k85IYurOSJTeceS0YXnnYZE5zsQ+LxdfKLUI3afBsOy4yYj8sSKBDY4l4sGGFxnY
52+yOCe4vDmFAK3QCqNHTwQBU+2I4d/awsN9GwBEyxphHANW+s7EFftIwjzbgfmM
T+K0SIdDC5o0SNzrnahdgAC1XY3sqbd2ovt4Sl4ztK1QKNqFdzJIMMbjc1JOvg1Q
US20NuUbEwurVt+9vuvxwK3pQCYRBY1jjyrb0dEB+CRDTDhx6dvz1FbVMq9vW8Yd
99e+Z6Ybu9XNgETPS6mI7OggvsMdDVNm8sSgwYQN4xAACpxBi3Npq05r1Bj34r7w
vdQrWUFHpsN9YH4NcmByagSbfwiZMt9SDIU8tXHMa8F2EZ/sLUwkATNqVH9p0xVM
Sp9yBuSqTRGORooh/V3ig0SENJLqG/63CsfXM5ca+gNIlEIrPNqgJiLmFY2toDWs
/kz+9SzlngSz2WNMXoXNdV2UdK0l1KKHkR3VQz/s8zCZdyUURgAuBqBuByDBiEvw
z6jSF02pm2NzRb+kW+pLNUYir7ySWGDhojzHeAJcJI3fpufM8/SCLH8NFOPXexrM
xedsMNEZ3WSFsoK10BzlhWR12SWEX/jJNRCApTwAuKNhHFNHfs3XVWKHQ2jdRptW
j2P/6Qxz/wi6aoeVhWbA0w0vrxoC76lTp3KmQa6QgH57k1GtwTPe0JKpTkMo9C0y
IlU2dfR91Y2i8GhaRqPJ2duN12AD134VXgyjkcbjQRAxy8Oa1re9VJGry7Ct6Oao
GDfA2hT5pdPKyl/6ffmg7u1lEj8Zqr7NZsKR4k5IkIocae9ZMyrHWwkcsnItfBja
ic+VelFY7gYngt3s7Bh9hSB8jAMYmHyzSfKqOt87kItoC2ATxKgS0Lz4sOttTN3c
l3XJDYaVpmOynM0FueEQGjSmuMc61jKjpAn49ZqcbAB6P0haYUavSacHlbwwnbj3
quCJL0FqDyomiY53T88MFlPvm+4xQEuCBpVHFCTp3GSrZ8F4/kEtjNK3ckOMPGxl
rC7IMriDqpTEz83n3/HH26XpZRpRI/46zxcLO4z+DKAvDKxLZEVpEqyXYhA26OI4
9AqCQ1/iQjFzzzl4NS68UFMp7WyYwbRA4urn07nqkbsgO76gZJ5zQIkoMT+BSKOF
lO/5ZLiYZZRYCqJsDfVji9IjeEAdF2UINMxVhgxfxSGjSsZUF9tHZGh2FiULVHHd
PDDFlW9si788WTTTkWqx1evzw2b2AWVCyRaKveA57bVouRLPywECatcJ/8udARGk
utHBvAHGdguN+2K52LKinmZR8ldzy26/Mx7mRzI21PLqGPFoytBSaPt9Mz3c4hNj
3dKMZxl9aSHcZIGPnhXAf4txQTiGsiwOmidEXUvVSptDdlXmrVYPq8mOF8mDq3AE
m5l1dl5s80xnusq7FIf0NXw4O3kWDM4CzlaqaAOGyU9XmGx4RtLzzdqIsZCwuSZK
pWehLHveMACiBraj74ruvOVErmuSHJ2/jSQKu9D+QEISXfG5fsfHfqKMeZkC0+b5
P2bX8/weQLFunUF81sORNOtd+IFlm6grhbb9tn2Gni8fB4H9P6vOQuJzc/sy1yxH
GXd4cIqwFduCpFV3tpUZNW1f4e6sN6TOMQb/kddoJq5vKwWwMasOBg7AIfFuOgp1
sVqP7YUDGXeckCMd3nPYy2ePSEyFx+KPfYOlgsn0VZrTZ3Te0XOedrE0B2HsQT28
KvtkYhppHGXNsOZAqE6/6dW82XKYQ3ZPYfSEjpFzuvYzq8mt5Y+gD5AL1FFsLFXC
4VWWNIuj6ZZGEewqiXH4rbiYQaVaxKEVEwm0RHM/AjACKLvbwRfUWN/OjD0hpfGf
iphIWT5cMOB02XPpvc7ej70aEEY5UlnPzcNWbk66Zvkpyk4Ies0zMyis7uyoXMI6
CTc660IIA/sFAR6/mmpS0pxy9VyGTn/dwYZcamZ84mI3fXhkn3Mt21zq4hwxTgk3
KO3NWwwtUDydQ9B4FCVgdAPeMg6hT23P3vpI4sLBQvz4Ir2ruLfLIR0D5tPFlINy
6MbwgRXLc8jPAl6KOyMU4P8GNhWyh6u2d94HoEUOZJpuCMumWKFfcmpMJRQ0qm1d
pE4Ad/MZbwSUWwRxqdpJd05Tn+UBi8YihtyF+AK3ZRBKtqliF/WrB7TE+GWyl+/7
tq0W0DryT+/5e+cD7EXfZkEDXDO7GRVbUlrm6TWdidXjR9LrESF1VPJrDtEG5ECj
Sc6MT7V1RDXCfSJPs53GFCuLLtBerkIYzXOFaHPz4cm7tUr35WLI2TiRPQllQPHA
wZwVkXU80Zx2f5SkUnGfNH/EZp7aBdSn9xZ2DLPWgxHGBN040D132FeAKrYeUmOy
iNmndW+YCyS2fdIhTIvigwNwaw6Q4vwamAOI4FBbxEHoxptpJYrB30zSRvNc+YN/
iAl6nq958Iexp72NkNesBxf2GXYliHf5t2p/xtYj7g0rG+DCfiCYq93BXvZYvoE5
2gky4w2RwMoNIJJ6JzUK9m1gRwRnWy2IquGAlQS3BdGOb04LpiA15aI751HYmNmd
Fm42R4x+KzWS3Z4du1QrLcvkfHwpJpvrJHv+ls1SKGWDW3pVsQUo00COY2w7ba4l
VTPN6ewDmNcHQkmf7c2f2j9n1CCTt81XiFUyBc67RBNkrmyLvVpDgcm9gcG6pIvZ
jfdsI27EWb3jyNA7M9IXzlRLgfuM2PvLfjayCVN2gB3ErWfCXtT8A5yabTtIL1Po
eGHj5rsV+ONumrw+1RFLftXNZRU+AQnLRZ064KG9VAGsGQmeqmYqYdAGlxXG4c/5
n8lcSBd/EHg5pA3vn5BseAuN+WHs6GOcGKJNepm6WwtG7jbyebsklhJWrUzSyI4c
2ldEg5SA+rBZul/ORmQ+JEsnv2za7t1TK0VdMtXAn/fUvZVXdIfwiO/r7S5xrdvf
w4KamCOxH3i00mSntqEiYH4jwNnw75KCKfkOqcMaKcFPakgT97/Kq8ReeLm8mpVZ
XCpZkN5NZ5arRymL2TFiRrFnSDnqa+/xMvyxz9hGmKeLqS1oTD7xjo4TBn38G8T4
QPzdpnitQzxw6mOQyuQLUT7DEJZl9eb5LbvluCxf959FB9GnY/yQO487FiNzSCZb
wE3T+frkuPZQeEewVc0jgWRVKYkC3vDsKev8uGwddSmUjYQAsESxMTrvyxTxEnwP
vBCkHzBIhelvYO7D7JLW/w2kFBGh1htHvuQZjdk/EwrGMNibItWPYA9IyEg9Osg3
LZ3JQCCpp7OpCAgXQbDgQ7/BTNpyDaJGa8nBl/5H/memhR/5yFEJmuzcvQJXIpzB
LifqIqXiEkrcA2NQ8Nmypla0gCpVC/hEzAg12dAvp89uRgrO6ja7cHykdJ5wOxQR
syLLUynTqsvXVFCLc4hwPJ7FdHPIFJNOzwoy63UATNe25GIlHbZCO8Xjp0OqgU8T
hbHGSLG2mAMQK3h82XPyiIsQD3j4ht+LVPotU1KgnkSaVo5P1vb6OXMMbuQnGbfd
YrF032g//UY8nWo9UUyCVKJORO53rHKVvmWBbScMsPk5is870bh2diKbmkcGJSbi
Z32vBscKVXRrgzxVCY0HpHmGvBtrVR/v+kfWWCsg2CF5jB8x6pmj3FqJdAsmYB19
KUVQek8OHZSF9EULFlPKVSIcgRBEJsQapsm40gwmTuLcY4jHuys9HqbIU7vWoWP2
JF/MDs7EZg3+7J0w6Ai19+x/BUpZcAySb4x4CIrDbSWDq6isDv8NHrsrvomAXDNc
iX+6+cVqGmk72gVAQLCosxmFs+Ad4qa59IeszhIaPL2KUX7FPMUPHOC321LgKtVD
smeP19tlRrubVzaYZooUMOmcToXI91Cqd2mEFffRTqTkSOX782EvFbXHBz5XjlC0
/qEZmsJRIA1CPoyDE0jDwqNIBl26Ew1ydzMe8DAUpjiSJwNomiQIV4bVP56y4IOG
jxtfgWwraNiGMz1UyUwxbdW7Rts/AsygwQWEdH6CFazFrLqwPGNeLAVYthODJHU9
6WvFWoUtlK3pEFI3WjW7Q8DCgRTKayx2Asj+PFYzTxYHEUeaFYCckqlpLKV4aVry
09i96K4O+5NehshGEULHx0fvOmGX0G7EE/y+95zbC71QpkYeG9idKHajqkW1hGx7
oA0J5duA58cIdTMzEc6/mFkwXhS060/o/gfpA5igl6EoAPsujSuLigIH3tDDzAdj
oYRdKfSFM5Z50B/B9YkcPSuKvfVc0KR+92eim8is42Zda82tluWS+NYHZQzs4gn6
uVQdQSv8OnEe1K3tTrpjsGsKWkbQJDAA7F8T8Tilsdbv5BfdTBd7ac08CV3lpM/B
kJNi1GeOv65JOGVkUsPGFO4PxPE1TdcnhdUExO9dRuRtUwtYCiJNWWsuusE3lkar
FLbyVlc9RPr5AEihvr97k2634DnS+ZHGuoTzSnJG9Z7/U7bu7+p9YtyJEYpm7K+p
5XH5A3GEZIZuXIDWSdsglrMNfdoNLzrFRiB/V87wCrsv7qo7NhUBsVYNQrxdQSod
vuNX05cMQBZ2tXAhjAP+cfjzbnGmQ1VAqK5Uy6Vxz5n02DLwLHmYDpeqJ31wgGpy
4cYSE08lv/1L8Lh2Rneox5QQipkEb57X0Ry5H0blpcqkhG+0lHGk9rihf9bXlcK5
kn9wv01IMU1miY64sUGEwWABNWnWo6ONsJW3JJZsNw+4pqXW0IkLtHfoWYFcJO31
FHy0DL4tJ90Gwp+rCDiv/C+6eHYcWj4N654xBwTvkEyfHlnbnGDaq2NOagCu4bWQ
xBhQOP7jwpsDypwQuSo3s7YO9PtePoZYrOwPs8tfac8c/HXd3kzEEV25Rgnvs3VX
3OUJkAeAP/4V0/t7Sp0z6KBbM2ZI68FPy4C9aG40a9X0CnfOe+s2UsUIFg8XfwmC
6jxeyQGPt4Mnuy7MJjJAHTvLgBcEsYSxYQndkK/DL22E30OH/j067UHb0iYLDRdQ
a2Es1j7PqHKqZ1Wr7JhGG0OZT3Wj/bYr9/fS3DMn0xSqRN5iJCBIgCi7o130pD9O
KwXHQ6kFMgsK0CooIW+sOw+ozpqodA1vlRwuu+/CCigtWRrse5FFRb+FuaaWmyo8
IGnSAZbFSM9aMJ+x1vLdxulC5lpv2TRku+tG7Gx5i4o3LPjr6f3bqCH/A68hySrW
qjBOUM8SmNZFS0YgnWDdbH8QbWuDkZVAnvcTzaKiKs2t/eeb5J3QY9eHXsC7F/ce
Mcrpnw/r7I5wjMNCsVpiiDmeYdLpypGVlwPbijEUehjmmlVAkxWKaEeUCaLlyRxq
JZIMIxQ02APavn8+3T8MBzFfsz03WkHHmwvOmnzY+MRyGvds34ChY8I7RZPod+Aj
AHLIMx+FWvD7SC+c6PJBsO7pfNCkrxqmcnxgb8f9wwyXBv8u+1At8OywBCAp1KBl
kd5R0lNFs9HN8ZKqRTLKTVcBgO6krVmoaXWueseZw5a2GYPAKsCEKq0OsHi+mXKn
y++fq92PK4P0Lbs8myHtSaRpkCv8cFG5yQtDdLIeyj9hiZlvssnDkc7icktk2GPu
saBTbSf6tGgOSh3Wq+WBzwq+Sjx4euU6Nk7waok8gIO2bLUme+ygAU/mz/Pm+obu
0+vSnymhTwK1XbqrXaMbv8+t43ceaT1BHUYqdNjsjr1OT94ZkzP6hAAetCAuhmcD
e5KgYK4H2HhEB17faxf/OYlPMwK0AxjpSfDQhyqcVIMPAk9hfrpc62ZJoy/l0c8J
+PuOmFhQMyBys3FBGz1yWCR1nW84KES5XCjcvUWZ1NG2iEL4uSKc4ZZ+KIUPe0Wx
GZ15UBOXOZDO279c1sQtEe0gnL8AesICJEn0XR6xfNjrRSmcfSZpwXIuHTVfb2Zl
WGEWmXWD2tlsjD94dfPuMK9VB/yxhefgIMULqPtnGrUhFL6QB2+dKN/xSJ0p68AQ
YjrT56XVefm8LAtshdIfh/htF+33nIyc3fDqLnWiFX2L8ipx/72YdyugpA7WiEgh
hnsOdLL0b7SvQmhKLWcfDGD8ckSEPO1rZWzWaUV+r7KLNqJXe4V1GoXv5NAc3+hq
2p1DLjLNNZqrteeCBRDbmZoAlGeND12uGcNmxhvFuxTEQ+Oy9heYl4QT7q4451bL
KiJAzgOlgEpX1M5W4yCVKNexJV2zBNMKFNsV+W3yjHSc7oiosyZrcA+iL7/7PCqi
iwtdLle0QBuSS92tXM3Vt0YbxFbh6tGL3SJMggVSNmmTcPlrdQ6uM8bMMlSE2jH3
9gGE5CONhCerG72cRtbLbyk8OMBsW/SZVDmLpJ+hP6UR0Uud5mTjbcgXxZSeSN50
LkTf23mX5sj2OB0DUVC+KuJDbokUQkfyGHQMsWB5+ph4GpsnXuXiwerIXtnBukJs
qyQlHxqQVWWG1xwJSY8LD8F9GaWCjI32iZo34mNb0BMJzO8iC4NVI5QbriFLdOmj
y/fxnIv8scaxJCYD49NhJBw7oA5eZcM4Tziipggpy3mHPDg8PgvevzQnq/vhtS9m
ilfR52ctyXNPJRb3JbB/yXjxYb7j1fYSUnCo27jMIOq/FyxyOaOwckFa729/5yB+
f//2TvQAnOPm2JETOOpCXzS6qaI644vViB13YRA0oKQbkwMqimVkI4hgs3F2Rpm2
OZV7tDJAsnriS9wO9gU2ztTp9+28hlu0u5EL8Dm00fRXXrog7e7p6YYpeB2x+TT5
RSuHSAQeRx0RPQ0mF2bbFIZsQfH4ME7/iRzbNuweifHBVZ8n5sFQcFI6B7Eb+ffY
Kcx0IJlek8lORVSpro51daVz/ag20jGUSz7vt92+qM1QqKzdD1FUBdBI4fWQ+czi
b2EX+EUt3NL8U5I8Zo/GTEFMwp4gOKnuMGuKd/2KZak1Z2h1LUaRpiESD2Uzk119
/cPfIqn80zto8pbzRGQBvvghKqVvzhpggMbOtYGaBw+0+rv3lVv96XWM61SUsefe
EvMEzAxFRv85rPe10S0Agx3sPo7hlDZBwW20xAQx9P0+UQVNLSFihiOX8JFj8urY
RqgsBIjF/76waJ5od+lBeV09mbQFZLBa6DaDWrNKrdry1C6S5pLqNGzDNSAPpnvJ
Gt6vR4cD89yId7UOwBgGCgR7judIk5RAIVLDGtsOyUZAr9k7k3d5GJXnlCJbvmX6
D2dwAuUopYsYNX8KsH8clo4rA96jSKBpoaUJZfnwcgmjJZ/v05HWxdXN5xCY4I5/
BGQgdZD/7BQkfO/J6chLyiESTqHKt9As816sA1JaAktyDZS+ipRj7wthTRW9rmbJ
m4KxJQSTz4NvsHda48WDO4Pm39xg0hm6qhCYMmwVlEMcSvmONYvJCkARvi6b166m
/a/iRBAnKYILZFd6ZqV4XBLlr0yHixv4sNssq+MeEMDcg+XL5IPvq7yIRWZw4HBu
MJelEoOGtyRoYMqSDYMsVQRg/Lpuao5QiVK4/C/U2XLgokSHKXIR7cWklbgFQkmD
xNOJbfM9ZGqRRwAplEsKQ58/YYd+cHa9Gkkl8SZx3eHRq98rLFmbhOX+f/mwuGlX
Y/t8XkDMjkO0EtRxbPiTIzqZpB78TbQGn/NFMNZ+KL9r5/7djijOL5Sm+rcWLnEX
GefCDMlJmaBz/b5RF6Xg+89UY8oRlrL5478csAsH5YQ1qetBHkCOs8ihXZBGfxI4
FVzEijLSSDzlU/txu3fdRdM+9ix89ouB4MGau8oF85ELOvhbgpnKCVGwCW2rTqZb
HgJqSfsSi2F+w2TRxA4PaxIHNE517bqPjH1lpq3M+PRBVsl4sKkZpiG9Kv3M5x2A
2q6aqsZiOHYz4LW5kzd4xbqf113xXAlciSrW+2AdCAhNFovQBwdp80g3s1lz/PXi
ApMbJIk3gPUS/uocbDuyTzlnZd2KQWcZsR5FE9OgFGntvJtyXkBs73Z+O1fAdsrY
XWAHmy42bAzFY/dw0RRLCevsWy6RcqYPAHcZOrS2OXWJbhIPBOPbAo00FICUIujt
tOfK1YR6Hpg4FKnC0+e+38T2L9+beLyD70Xx9A4ipGsf7V6jkKT7rC+MR5MGrddo
ehOf/ZKWDqVZRRzbVwWhAkvrxS9DgG/tP9O2nC2H0cOpIUwKjVPsLUi08uzDysIb
wPc3m7syORcfpnGccBXykQgncclWEiC++p2sFIvxw9TBCR3+kvw9Dx7fRsgtM9tN
OKNxbCTUfVCgfikWKZNiwUNEp+N0+fryDegGIV5n9bSICsVlED7iFjxSXyTB4con
Vn2daIDTUxNOy6NWAUb7gcfOxkcsN4/aaU9U6TrnRZ+1+5wBDtCqF7VSddDBOza0
yEcNKC2NdUL6KECbAfzpk2wpGGsK+Huj7Cem29ogChHBzP5qMcE+JMRv5EeEVd6d
QtBq8wANxwV5Iqg/MbWLy/Sbi83iukszgMD4AmO6xgeaUfH96mHpFpoke3xfZ+lI
jJhh2PWyHYhN3yx/sQq3/NgfCV2lqpPsCJDzsqhjsWMOAATsmBPCRlszC+olj26D
blzCyFzptgnb4FZZzCHEdUNUoZSc1RIOeWFdkiuS8N29kqgVVLfC7rnwEQIrHMHN
USeyZPt5RhvJuVBFyG+dlj148EEL1EWsvfuyp8Ztp5lnNQcaTDu/kOdI1ZP+lgLD
LzpRBlXhzLo3kLnPMNB23N2oXtk3jtLkKKOVrgB3GYjw+9Vi8a2MFeMdm6X1jm+l
1LlvGC2iP03qSOnQ0tn8gNHtFRSBNfv/B67fGCDRsfi7N3HClxHgFyFrE+hZyUZp
NrrXfDHy5P//kJyA2jWexgSE9hokvIQJtFF9quQ1zkEYQi+4ZwA3kTvhnmDbmSUg
YpEyyjUSrrFpKWq8GfFcy+LvRXyZztCU3E4ViCzUUeWNwE5Jn8SRRAMKST/ERJ/4
8yZbVNdGZ560Phvvnbo2Z/aCVeqjY4kilFnmLSAWP8XSEzqjZJLNMhufFCwfeIf8
rB5bUtpm48hq/QHG4jPb5I+KG0buXJ3AnevkqNfERwzgF+jZKUNkvYVRkoPNEGOe
HeASO43KQBejqNm/GBuoPHcW7r2fcNWygtNjreMokW+ZwWlEgXdbo+l41Q77ECzL
w95y730JLhtSWhz1LGaEDVBCz6q3lI+CK2dEiNqKKZ4xkfsjQS1Ae3PJdUIkbo3j
ospQAZrTOKq5Zyd1aOBWzm4Pip4A2UZtI1LpdDhQhrYJ7TsPm8arrmY0rmywDlFq
cDf8ek4/bSnvZ9GyLi2u2xvBzF/66PsiYnCpHV24365uObsEr2RYm1vcp8LX/vZU
gwqsYtoEk7rQLGdTlXPcBkDnfZfHlw03NI3dfLDO1BrsqWqJ1v8OSptaW5F/tZMJ
lDVspKdXe7C9POxtmh/YD4yaW1NAhaaThbLMd2ps3UbEweAonk+Z4slvwmtq3tsY
JcDKhF+Iv95fe/ACheOf0+FmJhTQAn1XUYN3GeNDpTtk+s8N5sRuglzz8Y2MukC0
e1ax5oEKlreFouYeMYGVq0YHO62tP4+A4q6Vnyv3iGrKo0mbgBGnoPw+XlGWp5JL
RrNQ4gUu9ibPakEljGWtZ6RbyP83pJL7uW207ZhmEpvAKumh2HMBD+fQkGeeEZb3
T6k8r+Eqy0dezLCFQ+PsB6PrmIP3rStHYP077ypMJGKB050A5lZ2s9Q++MZej9IP
DE4O+rJabMaHrglHBg4MSu3E+QhCA1Zp4EOp46q2MZM9Jp6aXx+dQu+tj3SHF4+E
e2AquDIPCpEG2fQ9lplqP9kZE4zSODj4/mSZTPlOgqWD/OvzrZcd6vEnWSJbbwoj
HvrQ4p0hJkHuISiD5rXSnpV/om/kZ7PK2dsHMuRnPUs9r1uhcX07Dqzxp2kherEQ
0TML+BB+mmu1mRdLIAyTRh7+pVQmFbi5L9yYh1H5eSlEW5fkq95A5llNuy93W+Is
E1gq6VyOy4JPoDoFB0g6VoN7NK26jbER6l/TKrGH6GzgrbM8YqMQB2QfCS4ifauB
BXGZ7JdVhGi2k1ajh5WwFCsjQEGbh3j1+aNVdFsLk2cw5ylxY3mGQ8eh0KdVZ16y
Dhf32Ng2Uk1k4hNMlmkoUa+M2qLkS1jmo+9H3nsTkAgJ+lEciFg/lIRyozAF1j7h
K7nQwqxc9Sp5x72JzM99HnXfBde1ANYYcPnFrc+FO60vMflVGdB3XrbIdmPOQFRP
uZyY05OtdGLb3CIjy/qSTdSs8feidrkrVjJSV2aqnA/csmbFkgHe1FqrKHW81Tqn
Ale542VhRLWQAHGfveQVqAV6m5x5Ll1k1nxJ6RWzk4wbGy2PEWR5/g85D5gM+9iX
sUkR0csMrlTb3wsPnOMwDoSo/oo7vzw4WCCl0VNsrzFb4jR7TSlwUM8PajPnLwVa
dLs7dV9bwMl1Dc61or3kOmQsT+2vM5W4iNs0Weo+bpJ3YvlrrY7npe1353c4AAfJ
Bi1y2k7sWME42zPOsAbefvZoAXbXvXhlAcTRaNGwtDiQ6buPJl9+z4NORbBdYkJ1
QbjCcvPSqWQ1r7tXfPdbPmc3J26Dpk91L9fcIcIoERJAE7auTdg1vYC68cXDtlnT
eosrfc3fXc0GJVNAQ5NGsAJFgTQIHqrNBk9RHeIE74goj1FbPxMFGQVtm+Viy+X6
8SRmDLfkBHcXs28Pa93QLgy392o9XuXbsXK8/gvu6IqSSmFjEl90oST2GMFKV7zJ
bougZ3uwhrs7x8DrbSyWiuTifuT6H0J1OSPiSBWb5p0/m5lVKRZnL1zjFp0agtwN
STJwuZi88v9tSeKZtFRjP25tlwT0KncXmT9hYhyVhjsTE2EHQEV3K519SQy//RMX
xpwQ+p4nV763/lQs/eLbjZ1gzn6jwzFuCi2dczE8l/EqyCUT3go0zzIHg/z/s+Ln
SxdVTZ6nFxJfvZ7lMqqCfs81CbkMFYF6mmM3FrHoGvmVk8ULDHuJP5YvhJrBK+sY
DUy7u4dchmuHkBq9ymE1xSrsJTgTO22VjdaUZg4aDvrkgrO1RS5RrNTDQizep4Le
djnnvumr4M76bAp2kzi3+EOr8/yOnEv+iLiFHaBhu3tWU4C6c+KoswUzC43so7E/
F+htXPjbLccQsoHzRejXkzrF5rWmPqUh9a22yXjBjeUiCfkVGg2V6YOQ4dX0JOUn
Tg2fH6/0AHujAbq+8Qle2jorjRgwXsc6/3kgit477JIprpjl0eoe0g0vy1NtCOWQ
IctSYPG6epivptmPJGxxKhTuTL0g2TXnZwqQnU/shLnjOc48GP6OOuB6sC4fX7fs
Gn6LNZX20t2+aeUxC59MN6mBQ3HGOCWzLeGa53/j6/iFXxf228NFVlHdEn+CyMxu
n5WwOazhpCyns/xh/XooDnCuWnmGq3YdsZlrgzIcC8KaOCQklBuod6avVbB9pb18
cZjhtKbUzvLj/rKC2DGhvTDxcsBpT+a3QJV6o2Kkc3Afksdads+o/sVbraVvLt/I
DnnlM9CbKRt7aQBjhzIkDoRbzID5JG5dJY5qsvUwF28GDPGCydseFyy0ZTzi48So
1Rh1uKqeGjsoJ9Xab9EAMeHjOcDJyB0EZXu4HCEkmRPHzLfxzJWMhRHicF7dmqSB
SQ86bQNfCEzazGaD7S8h7GLeyw170Gos86L4TLULxIdxHzATAIidU6RAwjy+dhQD
JAiLQGhboPymRcdI0jFeh0rpUeNWrtZMe1o39NYizGT3bxV82A3KqTTPQ51YEZ1c
pkLwr3DwJ+Mg2naATKC45KrEouny5pkQnOwOiPszgCOnoiBTWIr0n8fIV5p4e/D7
KMLaccJ9edcot4rZItjXsxDV8GUI+aE3NjVo07RiBYh+hXdhZbQuPP2nKHtcbtQz
Wt6aTqfYidd5Ynzndp0D6KmnC5mGpvn/6F33r5D2tfDXerFgzTEPw/pXwO1wRlac
q5VtqGJWpdwApaqKQqC46ITUPrI48C9Hv6lpJibe8IoSTbLEJ2U695y4EfB9xCjS
3ZPGuDFGgC+HbRTpaevZn3PujaLIOkmGH7Z/13Urmdf0LOtul7nlrZ1uKD4GjwXb
Wszm445bETSanDo4h9m1WIhSZlFV7JZUk2/u+v0uOtoKJGYrpmq9n80JjuDDNvhg
chvfONqqNvFaAc236EGiQOwX+LuglMspp6qQm0sr3JDTD945ZfUEDS8zeUZQ0dSw
l7otu6EmUnuWdgTihCMLNo1HQ2EMetitw1aEkOsKSyOgqTXLnIPlxGOL6MY+EA0W
qoPQZXt1O0y6xbk9sRo8AK/y2W8zV15eS4kWkjqMswcRBBEqHdgF6mbYWNssvOuO
gmIqXuRNv3ibGkITchmiFGDeCc/qhCRn+uGkS2W08riboOm9nH3e5SPiTk7XcYrB
MSFF0mXBvKHboBG6DNIbcQpU8Q/jtcRwlZOPHxel+dfvYMm1bdsuRci4j4K4GBAR
0DEzC6dhgRlwuaniAe2jRvLfBV2gmjIt2lw9rLEI/MCaIr16Rk8l8b7MOHzv9M9r
eO7H3HVjFCPnnABSSO9HltAhx4gJfLWWxvvNE0lhUIGoK01Fp3xIsaGisOtSdS5c
LkafZgdgALRreyvkRV4D83Bjn4dMWQc+SJlBdmM7QAF3ZhQXxV+ykc64foc1a9tE
jqhKOp3r/5KYfI9b8rxib7tWXpumkCzmQEMhgsgf4OKXYWkZ22YULNBw+YKJXkJ9
QdA9LpZGUcUxvms8Jctya40ZjGqdHQPdu+yvozJNkwZxpTwdsHIJdtKLO9hrk2bd
0wYHGH01uVcdOwRUmKpPnebK90LQU2XYhe9a7ZOrssbO2K0k6H9Sqz5kxmwy3oW1
sDk1uRYavEv5YBU5sGpT5lRQlkY4QlpU6LUKwn6gHphNhvhjprvmDEYOZnYl5jQs
S7dL9o7Ye0mFRCf+ZyJBYpu7l2wpKGZdqpQEt4Xt9dOYqnCiEBUMlupb6DOVfYYP
AcOyxl08BrM7Yxx3f6Tsv4esm6a8JMDGlFTmLw80XSJVAGSupTNEDgoR/QSOP6rN
XjIxe+/vxyp/NzgBrDCFpD4n/wIO7RVWRmDG7yIGKorq/wdzZaeywPm6z6vfWxVW
2ZaoFrLHySZiJ/j2VtILnvuIB7lboqsHYelCEqBL2AL/jxFt8gKNjlYCrb3j8O3F
7j3bwEwrAyflxETAjLQgkDGzRyPiT02O3DGIgSUF9+3gE4UAV4jY6KfNM7yrw+Xx
Dxm0gfDH4XWDcql97yjQ6BPi8OVXpQ740GvtosBN3c8FCs1ghjT6y4D0syFnfni6
D5/q+lo6PdDXdWawdSuGigo3RGhcPEAEQsHUU86Hq7zMqn9zgm+4hyANvH7ZIUDq
gPZAxtAhqkxhtJYMbybZEwUuP5bkrl1zUqM7wr4nDb1nedNiqHoeaaBxBioxB9TU
aCo1qbEi6SuBe/TgYwZ+xdfUm3jwqEAj+x41epB7BSeC69QW7VQiS7VrBZDnZ7yJ
hccp2Y3pCijkglOLp0126FIXTx50/Atw1vpxnFTOKf0JAmmVqybwXlei2rgU1n/f
ZiMPbhKEmU06SU7GdSgssQUMtorqmZJX1+tu6iOQh7MKdLfXq1voDQq81knmTTRY
XvePLLJvRwFrbc1P1FQSZs4BLL+6QJlfXrwYSrZZ8yiI5Ny/7csALsZiYuNygMHx
oeKay5eRw73pqYALLCIoD4yujSdzpssM0L5XOGRaE9abJQWnNSr2hVxUyMbU+pKi
dAFhng821xcmvKPRfXLGDftSdqI4xvv6mLCDChZvqIWpRT76Sp96HLtM41Ju5Qw5
/FLGmwynLZw+ji66xsjpnQpC47YBBfkdsUtMhdhzvZh3/I3ufT56S02av/l26ZB7
w790GD0kjJPTaddq5CCPzUnxzzSefpA5fOKI/1j11rqA1Igf6OlptRTUbVLVVNEZ
T1wz0029ls02uNEbTZM5sgYN1KU6x97gcqzQXRh98f9J7DDA/L5N3YE62OTwr7V1
xbxas5FhssqGivTWDR1zkkVHLmjqbMF9Hof765JNT/w/WgzI8GrcVU+kGAgVCvot
MdgxpwscuadOGNpnxNv2Ug==
`protect END_PROTECTED
