`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kuaHGIr+0b53kudazYNmG2qEpViQW8uDxkQ3lctpAbkGiTZOkDFiKMhjM7JckLGA
MZv21wkXyNA3aU0alrM2YmuAoyhMKs6AIb6LOdL+dNLL5i0f0OgxH1N6Jse07Rku
5oRW6f5TI8b6/3Ld+PjWLf04TD/EkcmDqC7GPwNr+Xi1AN68xmnj8gAqd/MrTobv
RXIjFQPA6WB/VLp+A5Y3LmDogQl3WK4FfFdAK6Q7VkcVg8pvAbp9AkG3TGTNAs5U
NHHQuASCoXCmpq3/IdJDVK/96AqZ1pZM9hvd0P/FtjDiKOw5Lloy4FuvqjlEnC+i
SWa6zvwQ1nVmX9/ohyrTbFaE94k2hs8V2YU54m3oYxthtzczz9zc4eYzOPqAW01l
bA+3+GYCxMEVV3RBSnEcLpc3/gSRNc2P4b3oE0ZybdyCeYpoICs/zmJYnca1FIyI
pW560BO15XiHC1l7pen/lIt6Lo6wwPXYPx3Z9uiAjUHDOKScNpqo404ulzSALsJt
`protect END_PROTECTED
