`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XzmiZA5D3vuU/HUZEzWIoUOnLuCHs41t+IBvWz+HbKpUu8upBmchAp2zdmfn/Dku
PfCyYbCq3TMGaFQLyvgnRIuryTF5f/rNjRTjubH94LD0cfu8CQHnN3eGUacUFgbe
X7V0bwwWDWIsbOC/dGyuus3fEtt2PUtj0ggaFX1mAEo+CWAoeE1KECrGcw3q4O9H
ZvCivFsx7C4hNAW6jH+ybA==
`protect END_PROTECTED
