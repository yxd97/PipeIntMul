`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3AZmd4+wM2YUX2Cw+BXtoBP4oaXwgbmNhYbpqVJOpAporkauvTDRfCmvxJl0ULs
Kku/P5klmPFcovj/6SyyP0Q2N4DPfhd6KNJaziCL07oO2bTKmpSvgyEJvwtHi3rS
foCCOCUiAETdvXw65pN6eTtaXHG52kcGQbMax0ev0ygQV6LH8WOUxUBFPxDkkb9W
DS/0DwK+Xlu+OYvtgaMj3lrr22yHs73fSeqYfhD2rMlCqIcCT7ZhyFq01S1kRUH3
6wExo0lsCmVT7NrmkrMf1d9P2ZgePB345W8/7Meu1cmg4vWnn3qJuRfzqnORLRSW
BHmuanCl2UOsSS5fq2+oF/z/iKfOWtQlsFnVjyo382QgCPfbUC+0XAvvEmyr68c9
MDNPMw9blKwAAIW3pT4f6ji38G9Y8sTYkJhpzeMPUCVPcfDdfkV6GQQTURokDyBy
6+G/BovqadyAzhopcbJAWUmhvdzfITTJ97Sds0pK3uidmfjFtpsxptJi8EwoKTN6
Iy8d4Ajlr+2J5yDteZ68Sr96Y/HpLhuNn8xHYPmEL9o=
`protect END_PROTECTED
