`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EyGzJxJDtPUGLsiaz4aHgw1QpPp8r1rXcoI3Utc1LPzRRjhhvQ1YQLsvn2aao9QI
lxooAdO7QFtAf1Du1BSR9Hxdq/wwqCdPP4zRnWUT2yc1PVUoOvtyQp8RhgfQ4jwy
R3t8+gzNrh9qedG90MZsTjPn9szX1hisoiQxMeP9v+EO6jm4MVLgHwYOShp/Nfwh
MrC1ydnotR0XMaFM/8J47TPFBCop2TBUOtHp4BfkphuqSSjBFO854i2/5z/A3+Wf
5fiDcYID4vo3QRCK9Fn14Ro9qPiZuVm7f3ipAIumwAP6E96QG5nGSI735lYm5yi6
GxtD7XkYsXxeA5AI8zq66WaUmyW6cdc9drjYj/1YOmEI5lWQ/yTYs/8b7SeoqgrV
Pm/VbVRjIIyIvprtt8UK8pUvyxDDAObHMnozEXtq2r5uuSBboS9aE0uWdJWJeFjM
zQDiZlEJNmSD6WCjvJKIE6aZHdAuuTe919jCqm8DevNw6fVjfACl0JVpcHBVzo9g
sC1g+7mrUWo/mJASAGQn6Yd26v4LRnCmNlbcbE+252VblqidfIZqnzcmNUAJ+oQY
j8XPZoi3G/KIGdjSsnD8AT93F39dx2UlwJxcvQOJjrcE/+BYjhSThyzrNg5/4vtg
5t+p7i/vjcscA0fVzc3eeOAXgl7imXbjFf0OC5N15EDB4Wzn33kYReT/aPughqug
Os4smNSN9sKcrWtNSamZgSHSty3dR3Quc9o3O/2jU/wvnzkH7EjTwd2ZJeUTXnd+
5ukgMaFpjeBqFbD1McgT6thBgtBasWaxWaxvPJ+tRf95G25w17JAO2PlLtjK0puP
G8OaZEzxu9zSDKME9LWkOyAZbmdEiuEeYUYjx4G1LW5MbfhSonVRN/i5kqjcOPgf
1auUeeWtTYbsfTzmjFYxLM+8d19nCAkEEkARGOoOwsgbj1cylHzl9DcoEL5IfQNv
PMU0AzIpThiTgOICkA+iIo3Y6crwTmWlvTYzwFR6HwtXH7vTDTeJqgs6SWvBumJr
A4BG91djVnUiZuisDmgUAn+1uGHCuRZ2g4m+2ob1v3A20aQqmDoQmwTs8GmiJ5Gh
XRfZduzEQWACSSWpABDLH9eX6yXx+NEu2nTRw4GCOmJGYaCVH1Xqt65SAx2KFUmu
1o5be4M1AFZ47bQGzeQlpNhvWO8ZzMz5tSKoG0nZJssKIkrDddwnbyo4c/XMZrP8
sukSk+zVXK+wOPoblS5M9Cwq0HnBvGlJZ5yRu/XePW5unvw+jzldw033RVuRXiil
OSWKMXJWMnJc9yg+oNL92bgwkBYr7u6iIc39Jf3Wk2ldOHjHcg+4DWfnbwPDGYIr
g7qpgXhHYEixhYYQXy9YIXafSecjhzY7cF4fUqiaCSsqQccpCnr25cYi6ukIeqHq
t+nVDxE8Q6gF6FJTbRtyl0dVm01ArDOrQDiBlCAQtpi1BVE5Ve8+Phlvm+LECxFm
7/YjXX3L5NIsUGA1ncltBg==
`protect END_PROTECTED
