`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKLCQ5Mw94hQRaS7+PL5w4B8+MaLWx7sLUn+/7O67AudUsYcdiS1VXvn/NeSNurE
vX/t6J3tZBBd48idelPHhVpddBsXmpdyxKKXFR9tvo+7EbA1Ch5avNXPUdw+wNR+
UFL4Be4xk7mFtwEB79WGtuW2CvIEXhLPiy90SB64fXEC7Ru7Kn8rjt2hC9KXhLm1
UnOhbaCsQqrsLGppt1nSVT3JbCmVl2WGp77itviWDwm+VW4mWD8i0tEIrQz2nOl2
SvNm24PiEXcdZETVTXE7MHqmwH0IcJPXBKpMxDpRTyMlogr6MergQccutve/hoS4
PIBLzjcHQY/hykUroxW/NMC5XhR6+Olb+UYpAd7f2oJNjGjlSrQ3L0l4Kl1wrmAn
IO7avvHRHGdUMex15oAZpAGFNMc45foN98736J9/Bq+Vuyy9Lzisrv0pLpSgSVgQ
2NlswWk3xSJbU9Jtl7Ihm8b3YABcYvRZP9tpYLlKcH4EV4bBUNNI9bl9BJ+s2dYV
AKRPnb1yD/9o/GPfLXIa1Nl+6f1Xg67GMYHmhaRkkotXqVZvFwKu4ukx3nEMMvrG
eC2xUi4thx1jbilPPRKfG+CUhSF4Q1vjQV6cSiqyGpDexYDOOHpGDs17xJZCIsTq
`protect END_PROTECTED
