`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K6+W5A/pgvAWz9YaSG/3Wo/+7oLyi1m2yVJBe1xPSBnhfEvroew4S30xvpMriCtq
7P+7zxAuxNcuIePW6dJoUyGlxUYcEd+csbNBhG3j1PxYoGcipCa3u3phFZ8MR8OG
Ek5pAiOLk7pZtSmHOE2UepEqQmOCjIqgbIQbKVkxWj34BGp4Ts8P7C/UMinCiqDs
b4E5PFw6rMMHuJxgMlthJM+f8cA2h97FtdJLLMaTzGvcvdE/jQTK5gFStcq2TbjW
PCtR0s6m0UwsbUQhL/TYLWphKPyJjswOd8JR1E+BYOe0MwLsMkTkzSCCEwlr/imz
Jmljz8nH+U415t5PLvrNGI+QKbikal/B3KNmMGjFQwSdOknaa8ztjuBjUqL9YpZp
YhGIg+tuRiZryfJPmf+gZgUKt1RiAzZ09TRC7gc6LrIZOBptwlDe9OtV54UXaP09
PMj/C/PisAwCV3wpCJ6YZC7zk31aAodevUYBhhEjcvpDqVTD+A8S7lwNRwKuseWd
ILztampHdGKhCJ8qmrXw2nJvKsutn0wRQTJQfXs3ik/EjznDxzaPLifa0VGUREdu
pPZ/usiWdO2HStvYgsthoNLuStafvy8aD4iCaaq78+uDET9Nio7cx2kXZgvZnRC7
9BkPXBIbLpYLboJTmTV27T0lCdhAEiYzOVhMMGGBCrd1co4k+T7op3BHsKOt8KSI
eHpyBzRdhqEZlXHHKFxAKVnNYwmYtJ9e/lG50m3mFQk=
`protect END_PROTECTED
