`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
onnD36vJ7LieQFDlKOWemzekN2bmndKY0w3ZOgE8J4my16SZMRbpRJ1Be0WVQtwE
Y5WsveypmVaLydLcMbixuljoCx2AgxVId/1DQSDexhgOoB7UxbBWWOkXqfBfUcDY
ivwmg8ZrJr4pOs3xGPc6pNZHcenr7W6bjsUvZfMOxhJHMKmOh7irsRI7AXz5iL6B
P83Yc2EiXp7DzgMiX/jDeY3E6e9Wfj4aB2eFB5kzZVQxgkWFJsjckHvNuPdATFKE
raA76CopntEWzndJ82Gjk6q/aDODDTqn1okZ1pUiClkM3roBn2jr+j66Pn9j19ZW
YHfAEwSr0jdl8VSZmXzKy55yPej07Ate0EkqlGGwb7g=
`protect END_PROTECTED
