`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SY1theNCDinxM/2wLd47HDAeE64xCYhHL4K9gs9JZ6U6H8DzKMYX3kXxsPjh7xaf
uCW3c8EOjWRIKDHZUgZza5i/TVi7814FZyWr8CTZ0U8rJare4xWlxHQcW/ubNysD
1H6KF2r0uU5C0hGc0sb95+G0TqP6Deuqf+iFDVtJueei4QhbMbj6tFip7ZjHWjB8
wRqe3dFTZ0DzIFt4+Tc2iPTgsUpt0rDjfUGLWyydQ8/SlDTmKk4BKB7KeQICRZaq
2x0UpcKIHkCccgfYL08kz5cg84R09rD7NzANX/fZVyPc+6BEnino7jv08S/Lnn/f
zpPqugdwsoIgTJcyIRNt7EKZMqzc5us0s3Ap3puLMVW4uQJdlgP9zSKUZhZ6UZfH
ScOXojc/PxciU8Xsoq2AxIxR534cMBSg/HiPM7apSSG54P8Jng94NSAdcAWREH+g
LCEH6h5amWBmSwddE4H/gYsFll/LxrvBt1dg7eGY8ml/pLiSEP8rIbyBlNbZ0Hna
3aoWwnj3QZTImp1SC91YdzMEKhEk06Woc5AhVcwassUBioDIR3VuXKCMCM9FXw+0
I8mjChNZ43e8YWWevu0tJfz3nztSzwoySEx87ARvAQwagC0CULMnkfPcLvcc6r/Y
CogZk0tNxHtC0UJ1BRncSgXz2UDIQvsZYdVUqkND2ULibwOeefKcLML1F75IOz50
rDmD16ug58ORRhN+W5NaHLw1dDCCMdH98cti3jhelNakfXkin1Fu95AFwtnfmVaT
EH8Wuo3lskLwojqOuQ49lav09ZHB8hMzvoH8XIhJDneefuORCu/tTchafGRdKdiQ
uGfawojpBQQQAIBq702AkHdqWsm+TdlZLhFaBwfte3t28BQU2Yfs3hiAtAn61XMC
ocwCDZE8xjHbnSpCHbWoIpSpmXUOEUaDxsdocTTpjaNbPOiNiE5+P69WD7C2PHcx
`protect END_PROTECTED
