`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ojn5SwqbXPEFOVs7E42fOcycFvUtr045upIznjosvhrgJpg8O7/DHTYNITHFYJWM
QsETO3bpTD6Y7pSapkDcM9PXcl+evVvEQft4xcvBPp1fK0DTZK5TDjLOkutT9ANX
H6PdDW1+Y/dmDJNn/OO744eGZzcLue0zdvWQVo6KAqIZPdRadIK3SglOW7P9tf5O
gRfAh711/6zXkVV4iEMpjqxAo4zqrOlbSi9eDNoTNJw9VahrOy+t/ogNS5mPjrz3
qOELddDk4pqIA7mUUtWK9x4pTaI828E1os7Ect73nNDL6ZdRMaR7w3leb/+YlJlX
maxrz5K7pQS7GU0RCVdMOlwNnLESVZ9v91z17cJmyKERc0wuqVdc1DTz/NQYxxSR
FH6uBpCDfVt0sTli5epdMmAhEmQ8AmIVzB5eqQXd5VE8NZPdjCSk+JsqTGdNjtog
iZpNO0i1Kr0xUwGoP5DiQxVXy5FyHgBKQrowK5S8RzCZIYqoNVUH7ex+nz1Wf3w/
jskSss7dUFIvs8Z3gAMpHsN0ZXWtTBkq7Tu+P4S6ptREr9h1Ipanq3XbXuWmfz8E
bZqUl/vEfGl1b3GsAYFT6wlSzUuqiJ85CKqZgG5cxQbwt87YfX8eD5H4FBjmPVth
FNuwtN5akK/cld/J9KhTtfX59flW8yDpHTQ8LMsNAktmLQ76sdWkZGYs9iFs0orB
gtaG5nn0uf3oB1GdHfXopw3uGFn1h5XvqZF2ojCSdiNtiDEJyBTCz1NgenTDmfRL
rVAMY1UgUpjd/dh1PbFxFJt6qN7c6Vpgi/zkaTc/iP2Z3GCVIec8s6QLJYnQmI41
/X6hePQAUZJXdysJULSpWkCnzGFwxTACQPhjT5kWPAiu1Elbr/xRzuXqhCh178w8
NdkCyL435de3LokopBgV4zE6FezXwpjokWMgXCYl4yg=
`protect END_PROTECTED
