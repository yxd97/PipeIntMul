`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OUVr5rp8w1LsMzqpekHihVNe+qgcbVWf+6q4Et1Api6vIEAUes01O174ZcNDw2hJ
KOWErmuIrZAWbzIlx7vTCjd5Dnmf7MSDfYDRVKOD9mvu2p6M1VBElNTXP7Ki9Xso
PU3y68/pR0/lMtVuxqXTB+cV+XnCvkWUpo3B4tXYWCg3aZkYND0M+d3uksB9vu3I
/1t1/ehbSIN9TbRRotaSj3oL6Sr6SH/VGIfAr5u9BvcfHr9YLvM98T3pfvS04CvC
M3Fb86ZPQ1M9BqCrq9bARjYmFQLAc9i4gQQ95M/TP3bUkbfX85+4ImJ3yHtWSRNi
6EFUVk9YLEWFsB2stzjtNh5qcSERq4c1bSy2jaHnjtWt/CdUXB3rzbHFYYaEGga5
P8zIOrwcZfMaU81EpVuiviheTBrmwxJrHyDXNXbNuHNNXz8bQ4Bfzw1tD5SG1xXV
UsedVYfAvhOzp3zajYiCm8mIFEkdbK4QSizqNyGpXLgEcAOnbnGSBwz7EVgdNPvw
R5F9uGm1RDGbPedX46eEoAQuox5EiybeLqh6CB2pg5/xtEhPilYKOl3u7mEJJOuF
1JLn40zfgDRaZcdrFteMocygdR8aaKJc+OdCfoaS2CmfotJ3ur09GwrefzUa7ZDA
G9W8RUX4On8sP1eq1gTc76dnpM7vzrogkVY0PqeMnJQV7ZSp1JvE0QiK00ZMjMvM
8SruMAUtX/9gZRsPv3GMUf8QUgXwjhCNleCA3RhX0Nm6YgxweySJY8P5o5A4rj4D
ApiwneFCj0Bf6VHzKA4hK2hR/oXBBv7NdQuyH2mJWx8wLf/2xYCmaHh9MNIsxPNX
pHGH+7Bi6nHOyQ3DSKcJCEWid3gZRzO5u9rfktUxMZvRGuC52+AiaZMwzjoB/2BR
AEtJQ5pLR0brXDlNK5gR5QOa0RYiqkc41IwvncN8x788x44yjlupajys71/I9H6n
6zz9ut07UFVqRm1kOYIeeYq4MJu0KInFbg8/Q3Qpu3nEsqVf31MdVRBDQ/f0X6+c
G6ZvhIbt4E/UFgQgfSgmwWgHJqJBST/Y2H5kzcrH3VKCjuL7cD6Z3NRKrBKZXDDW
22BdRzSYSei12C8asTz8zbg4eTnE60ijJnyk+98Ueun7o19PK4q4eJCyTZf4UB8L
JKnro7WBj57f263MivkX9xXawkHh77VaGzgnUush0P8qA0CCCYqwkF6TvFYtqTMX
sIDuS1CfWoQZ9OFg3+LBPa/9HSsXjyN2AYPl/T63M7vgYJr3yD4qPqhWjkmyhUZr
oQtqHhfct8myTnsO7cuZGXsVHJNwhWWTGSKjyDqMvuknPDIcfTpdqFIRcGTeT3yO
B2ZGZJpc0zVvzxgW2TYiks8uXDJak94YKWnmpZDWA4NNbTE8EFj56khniXmw9qM1
vHDKVe5grXIcCjFJ41WjgE3YiAQm0mE3etU3bAr0KT6rrOL1lXLeFv6uFHjLWhaO
OBy+vx+eAJtXLBOVd7xhbJuCMRy4l4V7t9rLj10SX4eurqFClM7XrkttmEEUXQKG
TD8ujF7L2CY2J6DojUIvw+pxbYk4ef3z4kD8d3x5YVmTk3RmPMred48+uoMuW4mg
n+AJf4r2lP3bGCk2hwBK+b8UhVCRW1k1ovpo2zK9wOjd76rl8V0kH4ax2HbB+IL9
JqAB5VsAYswzDSxNKHmoJfS2VwkBpHM6uK2sbakqsDuCJPnRK2xiGOT6qDSY8RYd
HMYSVJmI+PqgMcZnZJx6kh75jkczQ97/pJfnVfsj1QGL55+H9uPIXbmxwOSBrFyW
dM1nWasMVoqJx25ZjbgeIfn3fM8wlK7tnuUOB3NvePk/LEgITXSWgcwzPSI6hVRX
`protect END_PROTECTED
