`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0R/OE65suCr9pWvytdi/hidBUSGzt6lJurlRQHWlJbaeil2cKRhoDqd3NYOostf
QSZiyrDv7B3zrK1iWKuLDdxh/Xujv56a/T0JEXY5JLHned77NIYtKYJekCIKzaYy
XUroq3NzDklLOOYsUWc4YyAdp9mXy6Wd2xJqVNquIwE8qXQLp/bAFrgeIefjYrLX
iK1zOwqlxFF20rTlWrwGRfSDvTsaegkGumVajdsQab9a3r1MKexRiQpnQgzpDwVl
slZVHMi830q9r5wzBNK1NPspo04vEOXoJqqtRweQXWYfQnM7vfzWEYsx/cLhIN/2
uQNOrUnjUJc1MpM+pnnKqT7YLCfnGNMRCpm/V7NIP+Py0nD0XZZRyopvalP3nPMT
mQ9vy2V1xM7I4GMMkZNOWOSmUDiFfGNUjeGP/5yIvhXx3MiNH/IW7S0TIFZbqyol
769siEHYtFmi5Y8drrLE+fVrjlXjJm7QCCqD7eoR452omZddq9mRwHQWvU94fxDO
wQG2QFYAURP8v5SFa/sPBdr5YarFw61y2zZog3onBpRzNLZmGUV6DtDHVK9Zxh8Q
aOFt2KEURxV+W2Oi1hQ+kKiUWIgK3QQJiX1PKMweC+hgwjOCQ4+S6Ae9KyLLWIzS
MHAw0EMu9W0DmudA7GvO8vm0a4u105vq0T7rnj56xp9QRb2msZ5+57Bumg8mP4Kj
CUvF16PFEOxvlym8+xACGQ2rjUStd6b4aKdnh1EdAQ0=
`protect END_PROTECTED
