`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKHp4/MYNZtPLAcUkLZK4EEOr8NzUB+wGrfh0dsJHDyGetE6O9kcsL6CTdeW7DZH
9kR1xzrF79B40eLs6cJ1glyQxO53ulI9EZxvpv0ig0AwRGuGoQBN+BtnDolCvUIG
JttHaqZi7Zsw9uSMgX/a2XeinxhDTz3OYpv/geqrvr76fEY28qZ6g/HDe9VQ4skg
qVhoFEkNa0UFv5AVKO0vQoGEgByjCZ8eifIyGcVe0WidxjNPOCY3HrhtsgvrN8ot
pamfxRFO5J9FFLQmZo/CKQ==
`protect END_PROTECTED
