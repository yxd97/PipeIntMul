`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D4sIJXzxH/h+YI1Z425sOgwcYLy/QBB0dfj3WiU3WQv39UJpLKED/dOVlAJ8mGU3
PzUcxLOcl5Nz1VikJSSrtG1t8wJeUjXxpDcU1GTEvjoV0W05BfK2MECcdtyFXxT4
uv9S4AeZY/Z4/MR4Tmm7xSlyyNGpGr6osKzyxcDEkhvRnQsBgMbm4pW02MklLqoF
f7uDUXrDYzHLGPJhxziE1VAOmA18XKX/F9Tr3UOF6qDO6vUcmyDOE0kgUsBa6NNu
UwxlEiQtP39/CaYZPe21OXAAaID9oQrGMv4HbJXxSklOqWK0GwTbrnhAcOeVaOBj
KTCLUug4lGSzDaOIcGpTt/7CRcC9JcnZJovwL9FrqOoaassmdpc1wZT7ErYVLKZA
PzUqXa5IRvRZsCM7PBPTSF/8YZiu7nvs+cPn9bCQYlmC39XmYqWAOAhw320cyIE6
iYAfjd62ejtQKRGwUhIR6j73r404XP5ieSGb3y75foBtLu2AcsqWW6pFNpUau/7S
G+mL1pM+mNprns78/o7N0KsMJHOWFPHwjwJimZ4kTI8ElXvPR2AMKAWUUMH+9v0B
+vSaWAn4/qkrQwgyLfWvnhv6vOxEc/aCJ46Vh6R7IldzaW8fy86+dP0JV7tCii2u
/OUcRXluXrQMjN6eCGyQ2xRU8jxE94K2aBWkLo3YXmZoBw5SX7JZ7CnPT1jUYmkN
L5+vM2XUDKQNMIjusIzYKhqzDS9Qe9gl4QQoU+fDnNpxr1NXlXuid3RFByEkB5l7
bTrhVotgiNXoH93HGpEfvfGPv2kIRm/4L3kM4o5c8zhUeUT+762Mkk+Wf8pMTaDy
JiM4YYCHDdoYbbKdyJ8r7Yzq1WgFgMXz82Bn3PccjMHCKPQZhx+YuOo8YYkuCr8P
4u/4uvYkIiZ5WfiGpYCJLTHnGE7/Qpv+Ca3hozUmnNkhwmQHXGZ0AtviwYJ889Z1
N/Wch4mrogsWPzN2iSsfvNhPm12lo+G2dtBW9jKWGdDBE/pkWZ7Q3Lh6Mhclxm0s
kEolKGMVu+7GOz8boJa2CiooQRyvETnx+lVx5MUUiuragdNoVotzG8EkWii6ryul
Na8MPTt+xS0FIcJzlMATHY7m057GxRkTiKz1kFJ9ZWB2ds3j+ft8cAHw8Mm5voCO
1KkAduV2POZeRHT8dTtSsOM901ZTl6FM41s7v0msqau+aR6TqS4ib5YH4VZ4OPu8
6HcZ+X63Jgpqk2MvI/eGZDcaIBILvo4aRyNb0xy4Dvs=
`protect END_PROTECTED
