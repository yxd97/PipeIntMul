`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kXE1D3QRnv5Fb/5nVLG0lVlecuvjgmzaQSkZD+BYSNdYkabjJdcy47ehmTvy0dkT
HvRsSGfhbiB3EsHVIGpcV4CAKVb6/M4wIbB04zVcidCLrjl/hAGKjc3qdj4cmmR4
UKis9vV3rSveEbML+lmv4nNZH6nuIa0CmOPhP7T5s9h/otoe/Sj/Ga8MrDmdWWM0
F87mQQaYfHAygn148J13tKxEKalzivQYEvHlcBt0nS7jpQ5s5/2LGHOTdrrY8601
2cdVMb8of+Xb1ZaTlskrP1K2Uzr4yY2sJMYt5iLk4iEpb0GFGQs+kuuwiz7pbs4S
h6kjY1h22v+OHAkvZR43kg==
`protect END_PROTECTED
