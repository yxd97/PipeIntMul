`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1yoKjGltJyRltiUrK5BJtV/9FtdgZlmXTgR55IT9hPs0BDuGp/BEYb45fGn1WLqA
l+M+mVH3bqmPrL3gXQc24fzMr/l9TZ282l0Rwuy/S6ZOx6D2rGMxGmWXbiLoeije
d+8qN08QRzt50jh0z/gjrihxnEm35AN0jpz0q9pLK3ytoPZ4xvG4zsC1/YOyEBJn
WKC7TuglQnDPOQeRd2xA1a91gLQMHutSrQLMTAE1dhnpVX1h2WcRPUeWyqcE6Sbo
NYhmGnLRNKuRJT9h2ZhXuCOx2oEb1fFLtnfMJXCWIhd3wFo4K6x5CctAV3r2SBYi
giiAXIRQiSG25ntcQ2dY+rMkyq0UBE+oJj7Bh27djVljHfcMYpEXyH2XldVaGu/C
7jitXJDGowi5/Ka+mGxM/dbCmSflMMqZYQiwgho3eq8=
`protect END_PROTECTED
