`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQAoKvdoqT0Gn/uIabeUvyFIANQvTnTCGpKElODfNRn3Z0tAqx96LbeS4croWE1B
LlnHkR3/gV7208QmGeNfXDXO5DefmDK0uH0+Z7WeUiOZ2AmBX6KLg2JQlJ3UlxvC
tfddOI6K8R95SHT4qXVdc5JzuMG51VWX2Uic8+EuWafVJsRkmDfiurCAfLRC06Ll
oDnxLe3REIl0V2L7G380X8hvhRo7FqWHRjKWK5OfnBJ/wDrsV+P3E5OZis7z3nSL
yw/RKyMb08dX/WyzGEVDXBGcxWn40twDM6+WCrKadBOuFYbo6XBb0IBA6Hrbk5S2
61pxsQLyTmOx1TwzCJIpt0UCEqXG+m+vjbL5C1hsZYnfZnGDouUIOwrCDiwDvPGd
cJhjhxw3DdBsPiyh+tk0FFVQjRHtyvLodtI6D5wd7Pzn7Pa7BEfSzRLVi33Zry9O
7tvWRM1fWN0y1/y1Euzx+sfuYv/mZ8TE2PTyUGk4KfiQsvbcvPOKDrdiUej6LBBI
6KOvLW2JOveRXcOPZBe3O8k2qLtOL2U3td/Lmxya08NGhUFbNBXWtG03O1ZH99iS
xcPpPGrDuLxW/bSXsQ5kzw==
`protect END_PROTECTED
