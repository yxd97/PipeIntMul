`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5mTg2mN0pJO3meZ9srkEqwCOD31U73Ms80EM5rvqC5NRmFPDIbv5A80XBlKL6i1q
fqe31kTmzFuX71QeU61FrByvN/nZ0w2TiYaODiYwQevdh6UpcwCNTGFb8/+8uYXV
oRYrbZHMlULeIqbt6pxetnQ8P2OQAdsQPoW5AiUz2i1vK1aPz4u0f6JtzmlQqkNi
lUNSvBITS5nb3Ht0OYTgf0okGt52tsNMYG6xPdhsF9wDzUTqi24B8sUHxP5Qmbtb
fYLvFhuMzQOuKysxEoiB1mbkTCjl22lE2RUj8PccI9yQBOAKCO8kfor807+Xw18M
oUumm3Uh3d4NtZ6M3rh/In19tnHPYz6NpNX4b1XxdCwbWdLd1y01Skj70fntNKMt
65AhuOBLU5mIAdE8HJQlQPr80snE3siKsfFibGW/tJ6G+C2CnmKallm7+aL2x/sz
`protect END_PROTECTED
