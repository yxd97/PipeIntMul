`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qd+kG7D638CfXlakz/V5rjWrjOGztvVQfT1iSDm3Eu/VAqSWf/6GH9DOnmvEZJ7O
goUEy99dv8LFqMwSr5cjRUVY8LKji0d6plHUTvod61Loawp7vAqDxJKcTLXZbbHM
5i4qtmZiN+/kVvgH1GZ7wxreTuxcAWy5aeufIfs/ruWMcnfRT2UstwEXLGs6tgxT
A/xnzt8eVGI7T8eCrlZE3TEaR712FojNgS1+TvwbyrVO7HVuXraJtA/auLG3q2hi
X37AKdyhMqVHpCnFlifx/jtOyHQomNrBLs5caQOVMjyTkXFb9Vlnz/yJ0ZPAmV2Z
9OzHyjOBtxaIBzlyvs2+QjZo7qBDYNu1S5yv8yCVjyKXCBgtark1AVdEWWdJGvrr
Ny/VYzTXtb+ZU73zqyeyTaIG5V/PzLE5LPkZwwNdMzFlhSthnS/uP6lreMGJriT7
ExOPuwJbf2CpvhZFLtqK7J4JUdvAg/BDeTJN2CRlH7C0P2lz0aKWdr8k55bYjALq
/0Gmzo+5XVJJsX3N7gdqWBkXIzfdPZPd3E56y2ztyN30QQ/2nHUpHP05inoHY7dV
ewRWJwUkwfxnze6Q1ClG+m/0+Mn8LC9b8tjf2uLw0xQ=
`protect END_PROTECTED
