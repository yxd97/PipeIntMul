`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A28bZ/CHwXPbpgkI4xT8yT5GUMUy9EuLss9pnI3jPLuFUJ9lBYL2/lweIf/NUnf9
aZd+nZ5kIEDGfjaCtQDB5Y9pyeKvR9k1bMOBcAPv5o9GRF+1tFFxGtVCywlxuMkl
LJDno/Wn4sDksCvZzXaRQt+cZt6Re7fGVXcH9G9p3fe2FE4+cnQtb0j5oKzvHaOR
phw6IeEyn4i3XcWXoZSFtL3VMXjZrp2MYOUWFFdDjJT1xn18jx6KpNI1oyCazxgy
+b//Wx69BC3eGAf2IIjqTTCbAg8KJsvCmKYiM7z2H0Hi0pGo+pCHj+sOSdplJXmJ
RpZ+TLl8REOdkSK9MjCjX4+Cwj1gx8qal1197W+dZoAmkyadfeL/tBN22ZWobwfc
hZJOLDFrpi3CVVCe1iBSMVT6U2qk/FRWcFWrjyKH28IIkcWYBHjK0SLmgnsQwWOM
POpqU+7eMxozPsZmooAQdaeOpww/MULBdwChNT/aZJ7uG/iOKvQNRaT/c5s+milp
mqtPMNtir1OKSuG/lRsF3tuDRDUWPhttaDW3/GlI0wbYgGFSzfm00AetWcrOnKP5
ZNnITAZsbq0xcM/r17+WB+mkVSH/yFun6+5YnxBIhq1QxfTSeSa4a39UrfMz+kB7
sEIckIQGfxC0VgrzRyFMBg==
`protect END_PROTECTED
