`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwYclpyUHybITtbpPNiWcqbGPiBMYI8SeuC62h9SU2V9GIiKn06vhpoSJ5y5opBY
aAHLzDWoXCUSZFRhwmLYKj5IvLkpDaXPz/j0bfIg9Tyot6eQml5WGvgeLYYEaPOp
BcFsgDToYtLD0qNEJ7a3FAxD66+HupXnQzG7ai3/STkJqeB0sHNM0kYBW0cJmPTw
OtzK13EtT6Jhf88SpXWwVGLOL+L8r5EWkvJKmYv6ryhN0WkEJDySNEIvC3tD/8xx
GiOhCZpmiQC4tCu2ZanQ0tOUBAYzdDz81Z8wXF+zOVLB1+CFFU4fvBgrAbQnqblA
QjQdW3KLv9lfH7UeLrNOfx0pgrZ4e0HAToBO7O3YswWAQINmg4PW39Pc7LNvZwI5
+VgM1G0WjlVl/WfPD/Ls2g9MMmSIYVIULNnqliPGlLOQOoc++Lw5YmKMU0Pk5O8A
0XF8vNnR9q9rxXOGzqyDWLNL2wan6dTOicoKA87G/EZ3i7lh3Zdzb/YeRUWU2Im3
arDqT3dbUsP3MW6/u3JTHMeztu7fHZ0TmnFHsDTkU/XBC9S3KxyY54juxmTRea50
bcczQHnxS+ejmbDe8Qb7Gg2YfNwWhaQjPo9D2aJ0hYC5PsuCBQMYJmeqppZ1pmgw
cQBkwhzrkJDKZnfCA+coKp60wjTFfbTTTFWHHeGqGnacUdW0KmSACAZVXHLlgGUc
4cGyYpx8xmvqdpQ1lm7LaweVkVwbLlj2OnQ1vnPnckwQhNqUxpXqMVVrPpF54c6L
3D/xPYB0UZ6Tr6AD7suHSa2bMNV1Q5RqWr2yEeL3M+hpceAXPg74O0f/SA/PyHIT
C0KFJPhTXZbt7KqVxxpT1iG1Hxfi8EQieJD905rYPNx8PK2CQv1gdQyNef20x5xW
jmeYQXtRcugec8AToJtDRtVeOZy/XR5MUW66R+nnJhkANRwcd5oCVpN9/onqjnKD
DuKXH3PHSxoRKAVBnqRxXCMuFOu035R8ODyxc2aaSoxurnfIwD7QYt4TLIelkjGZ
eiKCLsLcFCZ9lPHc/+6cf7rCKI2QMtgyhsIYph6Y5H7Q/0xGKEnEF1OyybbA5yHS
P4Wday7dUKBeWEY/q3Z3Gl9lP4/JYZ+uWYR9VdxaaiVRq/E2Y7XxMwztmhjJTU3D
ROjeuCUI3FTAT1WWbEPrn+4BMOpGaIzzgJTVH3FlCMx5qQksyNmQy6CpzUtZPQ9I
fNhhtqB5RdeLXnEDX2f/H1l4IpMHKibb6awkHX3HaoY1/AGgAGGD3zi2oVEHXPUC
bSAppbB7Yr3a/Zi/W2e+9b9jpzIKIoSdusYCYkyuo1P0zOjIjQH2c7/7u2vVrYYW
UANXssIQXx1KvCseJjSV0S2EO4ugQo3OwbW2GKCYHj/qfv4d5o6VPHM9RJ5bxJPt
kWeFobJ3K2hlG+wKlTcq7FyFEmyayE9A6THQ5PgGQ5sL2vDxlRzA+6wAU3bgmUmr
wAVQRwBhCZ1ERzftODfWIGjUCmKKxEr+aEf/IR93Y3Kk0n7rczC4sXzPBWW+tugO
I3sbY521jupzVa5d+F2+KlUX3+VSPT3kTEyPYAjMpkG5ZZGO8IqlBd7BicnDTRNT
mcAtrBKChaXs158UAS9KitY1Moq/gH2a3ij1qc5BhOGaSoIu08zErsx6mxeF60ny
/djHtpV1bVzyhp/zoHq3mPbW6QoYqHal3KeHXsysDStgUazplK1eWu5xDt0bEREs
mjl7BtWb9JOIRsnrWfOpZ7MgtEiubgTzzpGm8rml2RHYyxfiUFnt7KEYdphJw4/D
BPzWMDYKkpCSnX9M0TVvZLmS8/T60HF3pqgYILyAGGtP9hv7ahKlSwq30qM0YeyH
eeOg/356n7GUXZN4nS5jGvorGyz2UEyYU2b/bgcD8RoDjH+VOVxH97VXyZMqapFq
DDWLMxnhqKd1XNbWIgG+duu+pXpzzymo88gzi4cEWl5rLjI2FZlrHieQFr7roG0L
Cud8IqZVxz9CsZtWLOvNuNJN5ONo0tSz0KnC5lOLF/DHUCpRxeYO0gFBAPUWwE6L
k4+aDjA259B3icQhGz8aw2OqId9aW5lxRp1fwkJeMfAObbTRkzwHhj5dg3PSafFQ
faIHwTDw0fFTUenFs+I/Zy8NvQl/1fJunNaTPD4scWlgqXm22fzbYeqe8opbXnTo
vvgTSRRxnMLgScMQ12qtIdtnmLAdO2nkQWMpqUWSax3S28GPYhIrWly74RS/ccYY
0mt/f8c3zbV22D7z4d3I42v4Ov0yK0Ysgq53mc26uIMVdDnTWT3S25JkoFSZNIY9
AEZJTVLwQoqVcmc5F5lL8Q==
`protect END_PROTECTED
