`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dnGxxLiCoM7NCnXwLhVwJnPI9uZYrTZLorPt+PCoF1NrZO7fD7Zfc7cY8uz6DHh/
0aVn75a4hgmbHKq3yctTCNbyJEqzC16kXZffHmqmoUAhOp3fK3qXsxhbFOi804tl
gmzeTSFlHeQWPmjxbqYXRGWRpKSqcl4k7nMqhLk9fZ45NvOMM3VgU2vpLBkv9N6Z
kamZOwXUzbp29Sjl/n3fTGAghusPWFTlr/y6v6tUUL6XKxm80G1/yKU4dsiqaNpX
ZkbsNf8duOvpvkJiOr8t08cFXhJoGtEdN34/LbV+uSw=
`protect END_PROTECTED
