`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nlpzPjcLGWZuFmG13310YY9WLcELJllbALPel7IYDFEgZqEoi8zlQpS2GsQxEe3a
0LYGt3NjmGsOV7zmEJQ3no7fPcvu/bTo1m/KNi/Hq+eeyVTUOBveb5S5MuKIVgw3
757cwyFNAOn5Axqqg11tCiaViyrt6lpE28Kg0Qq7akAIx1dB1kScgeotDenFWdZe
Yx91MPgfRHsdQZDgIfbohhqblCmc9QnPWqH8Wtoo+W8WiqrtxUqnAuNXZV7mkWcs
thf9KPmn/H8D2LAkXGU9+UR/W8CNJSHFoGsaNYuYoY7i9lKEdVzX3sAXAmdFTpP5
daYc4mMP3X3oKkP70KN2VA8YgVWhSpBHDUdTrgYpTcFrOmW0b9gD/R25WjU43Z28
2t1yUXa/vwxYRE0/itkkTbx22i0AyohjIqupOFWr81UJmnBGz+r9ueYFVkzkjbHS
W+SSGDlbdzjeCrV0tq002Dr72qxXN1p3ceEBVXN+sVS2oRp0X/svun9qvyZxbh9z
tO6dGWcmUVJ/ePHma/SFxkcayLMfDLLIPaU+wN1vTHzV3SZEERXkveGcaivV2C2N
2BkFoSyqbCrQSAd90ccfHsCrLik2rvOkXYqDt/0OjQweYS4am/JyL3OVJ7CSlyti
n1fYHviq+Yr02jsddnI9gFDd53u/iBFJpphH33wbsWjyE69TMVlina5grgkeim+r
BgBuAIQ0t/IZjALDhqOTQiHKTUHmWIJdW7+UxvxWXl3sDI7wGfCadzr7V3qpVxe9
4Nc/6I4cIKoS/yrBf6PVhcz/mr+IPO0v8dXJ5rvwAYNY5wxzWVIDdI+9+dwtMZ7m
kzoy+jkQ3M4k4Sje4IGzrUg6Soo5mK6rgyBVaOmGk18zOQT2h5hvybOfGJOl0F/n
qX+WqLuk5cw68A+j/CU3Ng==
`protect END_PROTECTED
