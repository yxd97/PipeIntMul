`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kif2QzSOBty6LFUVNo8keR9p2P7b7TLfHEZ6x/FWed5QGCZbZh6tQUirA+Dnz72
OJD1k+ZxIOEzlyNbbO5/0znu8JJlBFU+3hYZfsCGcxgQNzbAkLI68+9xks/eQJgF
W4V2X5OdAe0A6dOGbF43XQq5BLZVpK4myJHd5+i6dUZZW/qPJhKp0r8/a41QTCIK
G27XZEBQoeOvmDYlcmx3Rcx2/uoC9BWnSazFLQ6oMlTnb2L22w94kTb2+SdIwUmz
wOuBF1Vp5CaNx06wZuc86/mYnPr5nCYduqqV9t4ADMTiml9ctpoFZDaCzuZAeihJ
wNTMifaW+32WF76UlQi94weruPbIrlBF/KQMB43/3LqpNWVIl7cCDvkUqebtuwzn
Od8JHgWfaBLqi6eyeoh7lv7duhePvuydEiPWQ4rnXxGFLcnur60OFj2RMQBVDnWk
oL8eANrXLovWVfVtEesEPSBHl4PzPNXf27LEILWeqFNERf7ZuvqHzkzkUXwDjBvS
5ciGZH2uTR7wQ91UwEPa+FyUJS2aFRNLs4RfT8uEkVTdJZb31yUUyCGys+OZx9rO
WlsU1tTzuN37UjLoeYAkzWaqe1Aj3ILOlZ3dnqCbbU+3CUBdbjMlYbxfbDMT3sOQ
93+8k7j5Xj0FQfUL4M5D+Mv4YT0KxIqNDtyIR+LNdmY=
`protect END_PROTECTED
