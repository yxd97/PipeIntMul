`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdiKUKLLJa4dZfkJQv+GAnTtLUZgIZQVEOAinwsK3Gk6ebiLOiQjV+sgIDmJWLz0
auj9eh1qkAlKcY18vQsWfKFaBLe88qZvh+GKav16F5dRNl0erFYEgHs81nKmoS5U
yk9Yw6m9wNDIDGpmG+CXu9lotRSBzzlVooOB/h4efSAlqZIbow7NREbp9U/KewRi
Iyb6zCEvS/9XTmEi+5vjn8dyiH0CUNbfJtfoxVoHRDtL/0GkRN2kppP3PMrEAftq
nXctXfINuJPaBDWlhUiukELzeKptqyTfaqVR2bGNQ65RwAMHHQpW+b0llbX+98H/
ae9K3eAQxWZxdoU5MbOWGnWhMTsr2DG11IGUJJHJlNUOrNr87C7zAXnywHVlIgnY
/OoT2asvELI0Mmj2SRK86RzZ1ytblvy7pt5LLE5Mo99zYS6+a2XkqCmnffkoCKFx
g1t6eLtPu083FCFgz+NljsJB9AGmH1VrtKIS0HtMObXxloDywAKuWaGCO+d2BiKZ
djNnJ8vSAJHJC98T92jpYeHfCdwHfqHd2OF7VCY9zLFwb3vjplPpHgL53Qcj5YyL
eFmInpoakN5zGg3Dcb+Enlcfr1xYLmnV/jbDHeeDKAO3lqrHK9QHVKO/Wn0E0WXm
Idh4atpYDayopBBBUYxNnKmrAFpMTi3y9xFY7U/Mz6Q=
`protect END_PROTECTED
