`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zc+aDP44jZoLMEN36N2/bTUJcf3FVMAtZpUifUtv4kGzuiDMPsKWWLptmsQQZAfb
HyDMeSsU73C2I5OkzbTNq2OGH0p+903c34gs6fquTj64IWY7hhN0JuaEWe0+m0e1
Euwi6PUV86WlG0xHbqc5JvWdaTp10HU70nt1aM/BIAFIrFoILDgTVHyH/pDerJP4
zEMB360k0hB4j+LdY5Z5bMlL0YBG2mEBIJ0ywG6iCYy62FUYEkmVNJjdj6meONwK
JQLaayMhT1MmdFiV1Gycnq//SiSW7ex0xYEdJekFLGI6INC6pobEVNgfrvVQ3Cua
SoYBJN3g8KVdeQfxpFhugat+7lB7qOvE9njX2W9J6iCN4twJ1SlasXJEKobEBnuU
KfAXnp9HlXsoVysvKoOhPcyOl95N0kNRSU3s3r2nPSROIPqWHykONoo0iTzkaiQ1
kh4T5mxiXcwDvGHEB8N0Ldg1zrkqSwZiZNoA6eQsXbLDMJKUSyI3CagbZERP78tK
r+HfBuqgvNe77etloKp8Phk3lMVRg4UM2j7MUQjPkcmcFfl+E+4nSioS+m03ZEHy
cpFC/t4ezea1vF7rKcS98jQKl+xtnXXKrxrbNdFCxjGypS93FQ5GrxyHhfIYxTSY
UlD72t5MG+JveOY19neFLg==
`protect END_PROTECTED
