`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K19geURWmz8yRs8ZqIPZaYRu/x6av+CyatT1q3I0ubIHj4LoDZ6t2FgKF9RoNzFV
nGR5OfCmwScvgz+j9tnMzxeznVHu4mIFHIEGJeyJBf14vNbwl5E2U77k6fUlqlKe
25eBGkRW0CMsxWHF+Dx46CSkBvXwrdY8a7x8gTMrZGRXROz77lb5gNwGUXWNS18w
uSavFlytPDlUYx6DX++S9dnhTi2etZSk23zmWRHf5tUpebCr/lCwiItuBNN0Sv6f
MoFu1/Tfi+ahbPN9prvvhUPrxaHbZMWBHTHtm0584g2TSldEJecS5jilbE76ttsW
NDWiUWs7470UFzXUrudISwsef05r8G/wp8FCxBAC0//uiG5Bv4EWc3nO0hEs/ZdT
gOR+swcHk6auVch6IceH6ZSszWwYFP3WK4Vbb9YEX0LB7An31QE7HulL06JpPjWn
wdteNk1wM4Elt7JEi9/lRemKUZ3geSCcitGu9/70oczSX7w2nAe9mMuMknzfICtv
plSpcYkIDeMgWabXWP9lhRU64478MZwW79P4HKyCkPC5xnow/7EeDhEfYr/ld+qg
rZn2TOoWH0CsWS4PoagyUcA7dffSLYapSxsjbJGHI7nByreGy0E7YlA9yorQWYCP
EYv8b2uiMmjfLoTVfCxfUV+l3uVtzXvJsgXHqHHfGUFCyogjWfbi5OUbaH8UyYjt
LyXqZtfR9TxI3SMyu0Go2EgZhOWNT8ZmLUrwm6S4f+/xWCioJ1sWDfuFURR/OE0p
wvin2iw0nx7EPwbvQNp+fQ==
`protect END_PROTECTED
