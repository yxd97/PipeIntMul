`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C2ogOBz4F/MjGHtdhuYaliYkdR8CAeITAS+XIt9QQ+E7fhd398FYLSHZ+vrJaVmN
yecApeox+Jan8Boe6Gh3WDn1IVsA36onXDoz6C/7AyEPh0f26xO23hy/dFAYVqhM
VHeoFp+BZIoWcIdXNpCWDGTgXvcvgy1xVP1oTgCAINnYA56AZ166GXUwbPy5557s
WFGokxkvZK+Q4gxQuAuBakhEkeROvE0E1YhT0zWw6n1CnHnq5Vdqp2lph0nOkulb
KOUaEzFXQISdLWh+lx3PKPs/tdKjLuA+nVMR1uf/KM2Ok2HE0ow18ODefEvHo7ca
Q5HzjFSmXwgto77HvzEG5t5IJisvAOJc61PFItean3wZKcSg6J15xfyL6doPquQR
70Rnmz6dIUYaf++jOD5xmBhetUG3JFsBdOBKh/nBRH6/gApWMoQzJ/2mL66RXVmJ
xU9EfzoHCc2W2QiWxQ4+dXtL+qLFMhEsHzPnUQm78jC76Z0ObneUKOPnuGaxDJTQ
tUbfXhMn7RwULGpn66BPdnhX6920708/p0Q5B9Na3wIvd0ZcQQJw6j0onYzNugUi
`protect END_PROTECTED
