`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ll22dGLz1SCL45MMJtaT0x77xijTRrR7kMDu61Biv3MClGl+jZ5uBdJYy81z06Ne
ynkl+vWg69ebgizUK+7G/g+/xmYDVxQHr2pxhE71ezqgL2vRU9oseafkuonMlWZJ
NMbliEk7J16HienNQtTscs/ki7Zkq5tiatgwav1n8mqm6yeimdeQk70bts7YJ7Cw
mTDWTRdQniwS9q5Q9NamROgqMoKtIDENuzjFOB3wkJvoWX25xb2F0686zvANev4t
u3cJ5EG6PYZABjDcakxbUcKZ0r5O6gX6UxTq18/rChMhtYahM/BaEVVdpnRlog2a
iwsSDbEUSFWuLu6y2FXDr9eQn/s0X0u/11k+uMYn3D60C9o9qj+TvE1hFr52a8z3
FqtFcyt7+si0PRGVssVtXUbWv11fYnwxniw+0i7R7hqosrv08bPCWPx7OL0NRo+T
YjQ1nrq4xNty5rfmhVUGsP/jiApTf1fDn8DqIfOWH/5hrYg2NrVETrv3mtbPYofm
cP3kcyqKO4bFglM3jk0U2Nw7Bd0svxub1iRNgNt6CkqcSClozOVwQ/NWQMXyfXiW
d3AgtTjGyTJNjqK1US61zwze6tfd7IZPNgtjddSr69awZlgFwWfvZGzfke5D2rPL
XBwoGghlYJeReQJLyWuHezgkh8RHdhREFejj2+bp8/5E5G5uL4/h3OmHzNlkDDcN
VnZ0TIgLAAUNBuQQG8XTeg==
`protect END_PROTECTED
