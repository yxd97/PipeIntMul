`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VgJY0DSyNZt7dxbzXAP5R9pkseJWW/VIaudG6Q6HsXa+JCQDRhDjxYKkd4/OsWgy
UL6x3T7LdhLf7cBf7jU2vC5C9zde7kO5XBkNz2h2GSw9rT/bUVnTlQrhihHp4x3R
KlVo+LSJbDoikl42EpuKyV16Oo3g03iesd1ypYTbq74RJdgW7PbseqY8IEkkNxE2
Y2HaVCogrlCdDBb9CKssjVifrk6V/Mrp5llBfxN0nfiLDwQYzRIvP8TAL0pAeA2+
29XCnZpqODcmZIDPkEBspYvVnAFnPxRfSqsX59YmPkhs+c3O6AJImC8ZnuqrS/Dh
vEsE4Knn/PUxUhen9yF1LA==
`protect END_PROTECTED
