`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xLj4AVPPogreOZtz8wnNg2YVdbFH6zqWi37hLXNU7v0nHucOv9pTHC4k89xMIduq
f7SVB6x8PksBIKVkwmQkVyLVI0gleogW0y3bgaWQNsDyc4VPniJwPNmkB47StoqO
p5vHIpxJwyoq3o08FTffyyCZ0N29903mMBSvDNTKAbywr6DNUe+D9iIk7g35/u01
tx8m6FWCU3wK5m5oSEti9aBMXwpry6BgAulMWiNNmkgm5IbuNsN19LkdOQHE5CWh
vghrYUtVo2Zl/vbhK+aDHm1h7TXLs1nMkwZW2l28oLkFy1gOaFqFUHJdNmUbFZ+Z
TTUrD7Id9ibnGrei0XqNAo49XlDHlYJ3tNuAwaDi0EfXMJ9qRmOkZn69eJe3e2JF
`protect END_PROTECTED
