`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9buNiT1o1AWTa/sSYokTvx3BrvQEl9fvWFlSzW6pqlR/RI1E7HOWOhQ9nGsWft5/
mCX+lof79LzzfEDFJCgeKy3Wp76Rk2EFosSp0eSSSvU51hzplfwfkn5GJGSTZ3Ov
EJLBq9vrR447Xi10nkxjwVcG9bIstd4EksnG27xZ7pmsjL9C26MNJhfzEhaJQSLu
b4vfPZFqoPCv9F2QhXtjOKZPHeudoZYDhEGu9raE+ae3h8hWWCgO2RqfQEAYvvV6
VPQqtwZiHn2uS+sL+CLelvYKoM8VS6LDa8idzmfDOujaQCR8yLXdAlqVTl1FSLTf
DL9o5nLbga/fjRFCGEFGfSapaSkeU/W6pTkmviq6FciAAnODaQ0nrEoQC0zMnOGo
iVoAjtu+J8ulsq/tr2WkyX2wcI208fioOwLdFj1F5nKLlDhlChRA+vTz59I/0RZz
9aIMq/dUCfY5mWKAwnhoJG1hEfpMEqmT5tn/oBE1TRXDnrGTqYJ4zGVtU1bDvRUN
`protect END_PROTECTED
