`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdilDnPIPq5sRl0TQmOEXHSsv+wd96QhpUhK3knsFBJRITHO7HFleL/zZvRxjXQh
QQjIlcVzeFpxf/ZUWFP6FYb6KdyRjNJzqKDlvNQyVwKneWWdT0Y/7M9PTXmy/xfQ
vuIIZNffynYuMlF4L3bCeAtEnT2/C0y0JW82qvDQiGk/ifPFrBU1tsfvOwyBkbl8
wzNqSWIWFBaNpprjAkdhb7R7a4ZlqdYjUPS60rAm9FHA2BBr8peQaGqL3GVISBAN
ESgboAEreqBG0UiutodZocKeME29YlBrzztp1oNK6nHxuxAxE6/fiUDFFAJ+UksZ
vvtwJGfANqXx5ax9aU12YhpWjW06U9B7I+PXv8+QYIIG89iubLQ45Hia3Hd+Wa6n
`protect END_PROTECTED
