`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/OLBEti/hoZUXjPL/NW3xf9I+uhyG4me08qWvvpRuEsBfdQkd//10TV6+9wqjREI
1i6TsDxZEmJo/GuKLHa63EVAUNN0rasMaRgzJ9IqBKKaB2jrRCCZ49F22Cwm3NKP
NbCmacwcMXLoJh0BpC4oXZ+Q4pWD0O8UUyUoCy9vEdzNSgDsMb2jY0lGx1VQf0h1
MLUGucDaDo64Q7rLEr6wI2qesCreGGhzu2Uxwppq0gSJmsVQG21ehIzMbdvMYU+r
PWZ97bc5IEbwLu6a25U/JlzQtoLQcS6vw6pqI97tR/mW2MGZK/XvNDPTpsdGc+ai
/PWtiMUKH70Cx8bO7mNH+jZ75a2tBurIF5OnZHorzTJCYY0HboV8G0FCGgfgFdwt
aKwQ4VCgpjyp01dA//ohnA42yprkLkoBzfEMBvhfAHo=
`protect END_PROTECTED
