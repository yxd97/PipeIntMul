`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y+HlwypNlvhCoX4v51XfpovmchgS6HfUMfhby8RyiqJ8LYuLhhFKg5MbsNPOL4w3
AnPMwy2oCQTxtppyW8JOxr3N+t2NZLC0PGRFJgW9CVTLAvT/U4PM09pWInDE43LR
V8XFu+45Sj+RbjCThU5uxTtZZVracgWvfTkhqLLyIUCasmIvb0NL9uIGVQ24fKJ9
PA80ufo2d5ehgRCLRiFQuH+arLXhKqs9MJqSZKt4QMXKzKRqO/RxQXCOydUxjdYU
7uk3f98Is7I48hfT33OSjdjnOueIhA7V5V31qEYsrMG+HYNpBHeOl3tfxhAKZUII
ElH0GSJBBobS3xP4ZAsvXksSgA111TDWUIFXtIoPU9Xv9T4Y3ZoDhiMUEBoAtMYW
zEL1/SthU46l7pM4nBD+vIEapHJpRgMRilazp318m6Pb0RhF88FFiP89OoMwpzoP
OV93fEZc5fpOAzqmk/pi8Rx9enQEkH0cy+/Psv5Z4jT2YLRBxDLubmyw13rCdYUN
bPypWXklUpI8LG1gzBVhk4iDBnPkVPDR/qbe35s7QYgkPcgy3HAQwFgRtlgIQEB/
cpfyCyIA6f09uafmexU838mIFP3dTJhCmnMDvgIYwlR6lHN3CG9OFSeNlpVlzJhz
ZkzjQRvylDk1ilTT6/8Yvg==
`protect END_PROTECTED
