`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mc0+ikuHh5hB2bv4rN7AehZhwfKPRrVvmVz15VUm3ylAURZmf3o7S6JHHzwU+Wss
s6pFkzgRbesi2+jDp+TMpLu+tcZamwyhXetEykQT3QE8BcO5vC1gIKgYH3Gv5IWb
AzNjSJ1uR45yQ/yTunp7e4C25/Kamy6TBHHLOaroXNK9ASnoUY1qSMH149pO34B/
S7hkeX46KdgR+8H5CFQTth1RZm+/06GUXqBTWc02QquvAxBPW5OTiqGwMjIrGu8B
8hkeValp/4krGDHDjdej2FvnEtsWVdeODmhydKFn3Mux/e8eXFWOWu/Ho7CMi49V
vLG7UAMqAaucvkAj8r7TyTlq5CrJCreP8suNCs5N+2oTVHGyPbTwOCZRNY5xP/e3
`protect END_PROTECTED
