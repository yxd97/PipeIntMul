`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WT9Y5csQ9U4IsEmT5L6avUMtjU+tou/xfyykHOa5IF+9ekFtLRuHs4MAfzgVz5UB
b8xnxU2Y4/fuHeIGclbJUkYfVMVeT4h4/VvgNVoBmWcBJVX0HAC3j8Osqeqpr7WG
cHhAfxPV3E9Gkc1yyUVQwgL40u4vmG+73HBMui0oLaG2BGqGgzH29CGCA2ZrzALG
3GWXZB5wopiM/Rc2QK3IaZmE/fS7wleU9YI0S+XN+6LctMFbqakcyK7w0cHrTfsl
3qzx/2kBZ1c8v1pyI5LgxlRHVWHcpAMMAXlTGAyc85QcYFX+Ni6BN3rYWfvZy3I5
49Z4TEoco+dOkKqXzKY8PwoQmpppaDVz87zgpzXO+lOWL26BznTD6JPvTnOnRfsM
LJbh/EbQtah6kW1X7cJkMs0Yb5tsXJb4Akr6RkaxIhYXC7KxxxcYVZ3/QW0tC/Ov
lKHMt2wYO5MjKJiwI1Jici6zaoz0yVYpC0rjLGVhPu6HgAvDSustM+ng/sivzO6w
T67fESoVik498+CDW+Hv53u0EGrza/vzCF98JwpbMccF20g8toprvw9b1lKp16j4
4MwS78LS2RT6G6grwsPcoKYqwi21rPpLCa/iE2C3k7lkFB8Faj32StvEpYCkc8Cn
3ca/UDGtkFd2c0TO91jRiIjPIw2VRf3lCwozjx4kNUYQ7qXtgO8mQKR3epTMUlg1
8wZ41W2qTfYId6gemJR2Rh8XL6+xlE1MBzULSNGO7Nqc5saljPwx3LmNlCNCqyL9
UnMIVJtp0F4dW5ERE3ts10Ada0WpAScS+1KLaMhQ7NyAy/2JcCHa54sm3ab++kjn
l1QoeNoAkS/SraFXkxINSezfBUoOs00gPZNjjOOzCkA39ZKWI4keFOAeOnEp3FfQ
wE98BQO5Y2sXcBI50ZQRkCymxRIYZ/BtVBzE1Kbeq5dSDBp8L5xkLzSQ451fJmPI
`protect END_PROTECTED
