`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neKJhqp1U4Goitf4uJ9AQa7nKBP1egVm5FCDumrUm9B9sipv9m9Udgre90Xp7hP0
eknl/D1ZkVxXUXDelP8CCwj8ZdhaDPiAP0wOxmqS4VpEAQxRb02SZCYqsDtAVYTE
gwiazSTH/x9hdV9XJyVOJPINBEAZutV/VlkbIHivaaAxrP90ctDeFI0mqq65Xrxo
YlzI2gU+Ha9JTgOEr8ToYxDfSpwRrnsKJYotVkZTZXevU9jcqKRLuh0oJbOGl7Nl
`protect END_PROTECTED
