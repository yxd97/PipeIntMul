`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aBNO+QIcYuiNlaG9Id3wZlj799ZBUzd3HXoZpCva6aqnqx7ljuRY9gbvIQEsOEzj
1BZkdt+1TKaniIR2A2F9SyWisVZF76MJ1XSr4SW54COIy5uVqzTT4Cz3riEIfx2r
gwOZsa8YlncC/eWlEUN231IugnvfphB4KFDaI04xMaVzxlLTg3rWugbAq/0hL5AA
qd5UpsnMk+EJNr50/SoSHwD6xn4GwiSZiJfqkRIEStsSGmznn1WBVBIIIMTrk/hO
yuLxx9JKsdc5/p/GyEEqnlutn50++maL/wZsD8ScPise+EvZja0eGOwbvF27Rws8
x2fcS24DGGfTUAm83c4SfUiGt3xJ7U6bgQL4kkBwFCK74v+G3DAjU5x9GWqIIbf1
SDs+KbUKZ3i4KyqGUwb6MJ9/7A5I25vboc5KZO6hlT2+m0+hHZH3QWLhcYZYgKoX
`protect END_PROTECTED
