`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94TYbhipZdeqYrcCRYUX9rWXx5V+9o23ptsmIt47BGL6GlW1euACio/AuUumjCk5
+t3eyQFHHDC6oHxlHBRhWmgnXCqLehyCQwgmiWsyMOFaOB4KzaUBquyBa0WZQr48
s6g7Rea6gJ17qjuJ8C8enY15G7jWOqQka04DrVawFNi6rBHtbU7H80gpSdms0B27
xUu/g81ZOiKrmu5uFt3qvGXvLnTOe2Laq+GbOrlu9H0u13WgTcrPT3SrjoG68vqj
QDcYDhxr2DA7Kangk6edrQ==
`protect END_PROTECTED
