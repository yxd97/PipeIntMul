`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kDACcO6lUmla8GGAm++CEP3FZoSE33eiv+0wqBo2548DB8zclGJLA81cnPsgyYxw
qA7iZx22TjhwG7U2r+D8YIdWwjA8D3MtIa6NuMGrT+AyXVHrKCw1mpik8Map72zT
Oa5JUzY4zgzkDUH5UFfZYw3RopT80gJ8MKOzQPCJcEt7yVdP114dOgPCqXWdp/mv
zvRPlPPREpdKMCFrJVgACRcgvion501e9POquRWWD/LIsjIogpfNcXlsdXqOopC5
5A/A6v9SZXZXerPUMYORJJgVdMx0Nlp6nc+DYcEJSgO8gEvCo3b0mQEwCGS64oUe
9L6CShjxlzB30hQebKIP13I2CO0M6Gom0fMl4NvKSrYpcYWw9qqyFoKle8JxoGdN
RpkDILPTDgbzwb7azlB6V/uDEKV3FIalFZz+p56au+qv4i+82DjDPVP5FYIexl+l
MkhhG4obY4sziAuk6J+LLKdqObvVUxaJCf6I/310bpGwOLnfSlsZyOEb/Qho/F43
axeTfi/r7uqYdXSDEpeIUE+ZHpBoVgCEGcNVh7aVoj/zE+0XQD+sQRunTlriVp8x
d7vsF/jVovDMt8DGE6xsHzJqXzM7HFTRrYlfEQAMtUWlazwzWk6DEy7ClmTFDMx2
imXudEN5B6MeUqm0AXijCo9NByMcPAQGkc5IE6JipsRlQxoRGeaWtSNulPiQ2GFK
HmRbuMMkGK5enXNwDg5xVTN/R3bWdP4aCpI6/1aG0tHpXUk6jghjJcRosDJSn/T6
erUWub7pEGDTRJeNNUyqNSOGe/UMo8Z1ZeEXFxdUJHPv4RE3JkTcEWlS3XTBr3uL
IkvtJQkWxiEXmJ5sr4/KREQaFIZmcT9hmMEaNcN/lNT0cl03t4FI2eMNiIdD5TYF
q1bIcNaEqpqTtYPD/OYOl1beCZts4UoTCm6scH1UHaiiApcIBEGAjhmFfAXiDqAh
WFkkxL9pEZfR21Q69w6L/CpewISZxVrNgKfpIJhvA+36BXj+HS7L0TqWktQoVizL
Gt8so8jCgXDCdQSNX5C/K9P2GTDFBTJ4suBYfnvUbf73DcDMlAtf7qjU8LO406rA
elibK3nq6x/R2qQJdADtGGJneVpM3dhBVL5JRrqKHw77ReWrMCy4LsNqCqAv5UWF
NKrQ3g+X8ZOcWSsdzi5HtXgZ2GpJAlr88r+HbGSFJ7Ey6eSLsHlEnHRrPzPFg+wN
aQ0CjmuApLI/DBcDfBO+6OF9qH66TeDf754eZJHiBGg000oEQswadShWXHscuEnL
BIuMnwUwCNIzsUbwjZIuz6pYvEJu+cFFtA/TtRZoXW73QOJEl0jAI5OvvTYHQykH
YWVd2YQCTXNAr6DtRzX9fRLrCOxFZo0qES7sIEe2MHNNiHo25e4FxPtp6utbFbed
XhrGLPq9HbJWg3xHEL2ZOcYhi1HjHlnm0FSkDV7QpW3ihPxJb4y6D6C9MNq8s4OE
5XdOZf4dyqBbe172eZfZEqK2Narji2K3sYg40Kdtjp6Ju+Hr0Z8bjgN8d9Ifn6K7
9UfNmHu+J1mY4TRa9vV7RA4+wU1ZAXkFFOPi2Fq+GQZTQLfBcOtfulLAyhPYyiSV
eRQUEMOJ9JsrmgLKpzMGivYfCXUkmg2j52KvMUDWbbB22+YK4Rr9ddMWPYMAL6j6
AZDRswhcxJ2VVMfuFC/8PqiuRvA8KPVEwMceD6yXDCz5xkBWuqaJjzWmjh+yp5Fh
LxiBiryjkvkdvQov8MdRLUS2hX3n8RxLT8P7mLH97LBX6tJTElZCucRSqCBhCjak
E2X0NcLcwXTNFm7JE/Cp8iz10zn0DtLavZt6nWXSlkfRES7nJj6OochOFQaWSJAa
af1b93Ib9WT08it9wtENcER3uWemg2YhWV6RajVRlKCDtPjjuCauBeaePK/wEwqP
U4wH65yRopzR913ZAc4zS1JVQZD0JvmnXhVByZTRQsBvVx2wBDXIYeEvOJs/NWvX
o/xP5gfirDr+pjk+Y8m0LYR2614fJyiCyJ3O7OXaPWqub23J4IXUzygdcmEts1RQ
KSESewC/hg6WAtuHW7SxgmXND7iYZzUcH6TfqXX1vrvFI4RG8AgtdgrUmE2gHGSB
BejHxGiK5b8RJ1znZ6WTqh0YrEyKdUMPhmw343rRwYI=
`protect END_PROTECTED
