`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgALlTeWbFqB/niK+hi8RLlYs+47aWAbBFXkzg44xuyKWBWn7OUGDlTtLigU7kuj
3XjXimV1oqZeyxB2nsJk+DWVQDn7ZPGJvL3auD1zZy4G4BKgAVj+cNqMIkZhWJKQ
3TqabxBkx+r3TsG6vc3OdSK2AnWbUIVWj+EcsjKFcoCm9GibtO3wKp5ABH8Cv8NF
fTd235qGNj3gRe0Wt10Sjk30Brb4XsKgTTrvC6ahvye1SQgDa0uSt54uOlJicXeM
GCVfIpga6/QOX2fQ3SqO7kPVJP3hUHkMDN5c1xtqqj9dkuHGjCwhHOylE+J3nHFx
gKLn+42KInwaVE/W/i48wD8A9vJaHQiz4iua+WdHtxQL2cXzn0d4lDYfiFE0uS9h
BkBzKbnrIYg69yyzTpIRt0ySE3Qv9admYJCXA1b9Sy8=
`protect END_PROTECTED
