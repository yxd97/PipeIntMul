`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98RlsEwvc1opky+xNIbLpzkBw7L4LdmZuPDOY/lPqcjRhv5KHwkCHusBZ6uijcwb
4QepbYyEHPN8nPTwtm8Yqvt4eHE9658oxQpDccMvI5tnh33rSszJkfgGDK6E9ck+
Emh48DGS4rnk7evVlqHUkN85yk5LbUDoYnfNxW0VYaoRTTpts15lB6mcNuslJ41z
gVsjedc96CBKBoE7GmDjMLpnLZsJI/YCLoe+q3G2cvPWKWckG7RQzYk15VARdzCL
WPqXJr+3zJJhfS9AhYLioJ6MlVBM/twEEgsC70SfqpoL1tKbVdIPiQjrMPg19+wS
bR8d/GnvjscIBjYIHFR4X/MEb//Q31Z8goozhM7t0PaX71zn7sPww/fbI1FAc974
+5u4MYJcAayPl6NVwrQaCJTSlkdaY56h0UWhViaXlKJsgHhFBUx7ynlHnQSlhF3A
QJCeML+d8sdpzhDLush2U7aR2N6AtKJntTvLfDiyXAoDKZalGtixFf/tJy7W7QT+
/HXv61Vpz/+bNZw0QoZjYLDWqWyPgibK5LqzL2YHwU1GPFT9w/2wsj5ZTzyvW1XR
ubSbwqXNMHZFLaDXhxZDTQ==
`protect END_PROTECTED
