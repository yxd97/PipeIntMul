`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9H+/S6e+xlxTqfHTVVSZ/rQ2mAH0lwYxb3puR6Ie2oz0fuEIESadeYi9+I9qPbIs
NxaY8Lz3eRFwYcd8mFnfcgDemEcjlvRa0W6oRC3ERcZ2O5dh71F+atb1LBS1vn3Q
CD3KN74FADflD0ReG0PoYWY0WE77JykJYch0O0tKvM0zvVmLCpg7UHV7DEnMOT6T
lkUz9DpxNOjFfG8tdJNovCNg1QBN8I75ifDs00Mdf8ibQuR525Kwa2ESNycqHs8d
F3A9UET1gbE/3/EoqvCQQjNBmGXlDFIZpZ3xL18AJA9LWuSck8mjZC6v6V4TQcZo
XJOJesZ6SBbsFpwnXTc2E+yuYWoHrqqt5E0/3BoQ3InKvBPxtiIZYFHkIpMgjslT
T37Vtsg5UmvIqvKQxM39olR0rwivKfwliGRGImp39D/+PMcHQL58VX5LAF4Tybhw
7TPkt3vg6Yg4hkN8CRgByyHIsyyoyedorn3RYrtPapMyEyjTfXGxbLxebkgOvcFP
JnTV9jYYY76ur+jRQYqWMTP8WlEN6WMwkFW8veiy0NjTZk0FRWbeD+ZqMk56/qs+
8GPqu9qy4khaRJElUhJKeRq4ZMhEySD6lxAmaqfyncQ=
`protect END_PROTECTED
