`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpiEWxLEwRqWAvg1/HWwaGpKOSEGbrtcjpxuZCNYS+gD35gR6e3tuiTFwoRPDhu1
LAURG0v8CEoOAJdz1VuG93mgL7pZlQiA0sjdNpuG3VkoaOKXHaosq5TbBzDZEKlh
CLz5L3lb78yh0DFQyvakNHrABfv+o/I/Jomc4FcXRqKDiS1dg6pWDtOsW4QNSB0F
tViz126Hz1LxhrlcLwwAwl2Dwx8kOHrfkRcexhK0kHWVXSxLTsWBr5ZyaW/iY6Ob
wDfAFM2GIE3vPiXTuewMd4VLyLn/X833nD/GgzrIxabX/j6G/0kUgWGLJq6M3x1T
aLINJwU/h6nN8mWZ1MhDa4gFkTZAtWzZl0og5waLiliI1D7Q9W4yViqrwQYBq4fq
Tcd/p9E0YDuJkXD4xqBNSv1LGFc8WnwbXJjPj9PDlCE0bIBXAE1nh+Y9bS6M5AG9
ua6B08bGnptNVLkmDnpARp4LB0dAq4IV2PhqYcek6oStECi3wonmz41jUVb5mU7+
s9Ml7rzy+DqWRFKZ4SfdtOv3uJxQEltOXJkwUyysKZ/UFFbodJqOGNhttwv3hJPE
FfZPbJcqYDfz0Av4Klbrxm4/U0VGMXvjx9j2ZzD03JF5hTNmHoaL68c3JiX8K5ys
XWYQrY4NgEswJ0Q6tFGKOCPZ/9x8k7rv4MB/HPREDKfU9SyuMAMHjp26uWgHq7za
cTxQsSxmnMVfAPeIn4VyJm3v3ll81VoqJut+Uxo6Sb6tVzOI/ckF7NvsMpME6Cwu
XDXo35dfBUfsFctLUgDZWKjCj+RWgHSySSkkXk4W3f1KnFgUXYBTJGG3N6XKAN7L
vCFOONZGq6vwQpX6ZwmPmRdrHI6nCWF3rRHyhdY6LKuvBjEEs5bnvMl3i+TDR73B
LaqOLyTBckzEPiMlv8zabKTWXtY/4tJfujX7xpcSE9carRsICHc6+8+zShF9gAqC
cbZsYe+v/5Os+YhXMeCSQLTNBgi2yyzVcy1g6Ftf6400QbRD+v4M1NWyWCvQjd58
`protect END_PROTECTED
