`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BEoPyDLlMkQh7gC8djTo7WBdVomyxzIdNDLcIvcBvgKyw7s2sliQCz8NceAuej0T
cRz0BMXgdF3YTHNbsEWhWCiimWCiCFlcvR32QVjWGDlyTZC1pN6oGv4ZCmM5WO3E
mFjkPdMIn5Z0L8vITT8DwT7oLphgwkBAcYWuH+NPEVaCbYyGZo7xLDGF6gfnHQ4V
P79McpckW6nD2mNCJD8YYhzOIuKoOxxxri855Ct51kG3liZJQF8CaAVh/oRw9CAJ
dc50IxFN7CIfcssenp3BtP5TjEKPcQC5XeyF354uEoKB2de8LQrRYK62Ys3I5aBW
ia/Y6M9gcuUi8PJQXeodiKepiQKgdOCNuymeN92Zalu/EQYOwaJdxttloxh2JRIp
NB7F+M04QQSoWAjntitRVQjrScmZsj4bQC0goQmGRlROUvf7KYwUaXqysXKR4vpP
/JqDn2x9VRyBSvg4/JPMCl8NHhCHck704BcWCr5Eh6eoSsGmoatV4TIGk0l6MnjO
Oho2TPxJv5pgdV1hOWafLBYmbYqQP1KqZW5+LDAmqWrgDl9hJ8zhxZfplnILXXMa
fVmVUbwHc33Wm6tDJJPathEXZr98zhk91Yz/jGOC7J9AXz7TwpBOUW7uofp8nOSs
5thZifRXMyYcWacy5d0m1CQCR+zubOzlwrZfs7VMIJv/Tn903oH7/zF2piSffKok
MGE+HFGGyZ75FFSRyQzPwa3axL8ylB9QIhs66Jv8K8CDdtF3ty+k6G9K1bxZakNd
g2XYTkr/LPCeGVuTLcYx8JJJmGc9sTxy7FfrbHPiCh1VHJA5iKXH/RP++c7UsAs/
5pSq14qhzYnAyIrk2J0vUW7H/R4HQlF7LWcWbO0Y8vmrYFOTdj+caSHtHDDKL/J+
rkjP99X95WjLbNxDJYdjPDKBXAmKCs/a+lfB5vbyX0YhXLI595OTR5R/iCsipe2N
aH81KU6atSsGgCAG14JNKVa/97Z4u+VlhhAcSSzuJzB+5TOCM/K6M4UTiuSQ7/qv
`protect END_PROTECTED
