`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lnPtY0P36iR6zEAKOsHbNwIEX9UJI5Pqx6Ni+kZqJ4jPIx8gRYYMTzxMLryzLo1k
Xh33qNwk8fdvZrFzJ4vj3dXubKH+mXpD6GOydXRTuSiyhZ5iPKPcxH7C+aTGUYXY
azFyznZhwMRlv8M6kxcw3FQxhvbkRV+BBUqM7WRhC3Etg0z5Pcn+Vrb9fo3M44eT
fqXCwRn6s5SsO+JYI0MUmEGOIdSTS4XFjsCTUMbRCse0Q5QrYdiluaF1PwAmKJfL
ffak6fscjnNqUeirw9NDX9uxvZhSepRjB+NySd3/xy3bkVUo98oMe7Ns7bCfaoxr
e5sCLj3aB1PakpTu30+pUC9Yqoee0oDVxIDzvIpGYiuWwvGXoq9sPsBm02uhyaSj
nfkRKeLUePCQS7hu7KDk8qQvL9sSkklDydCU15h2YhmAtxsRgBxmmGHFW4a07Jj/
Nt9BW3QdUh+OJIKBG372lkYVG5J4pI+c2oF8vUPw/R5gIvpWGYHxTbvxShGh0NK3
Hq0LeWoJfDAxTzzj7UGpnJcYlUu1l4NkE2C23iKqe4fpi7yfeX/af7g1rSrzBPcV
vbc4vmX+tXcdM07VR/NERH40e2+nCDgVfDfNvBAwQN3Z/oo3Tv8iWPkedLY/dX79
YOWxrCVBOlkSFtH+m8fpazq0nwu7ry3UQ6sy4lXmwZtHcADi5afLGBi2S5aGrfH+
A7BwHqCSroQ45B55YFcAdu89Zj1Rx9j4wBcYFs8PbQI=
`protect END_PROTECTED
