`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k4l6obgsOnle1hgTMrrRgqNLSMdLF924JOjnd/FV/j2o8y/w81fHSoYsUuR03prq
6qN7NsElA73gjsQuW/z6RwUsJtb77uiRrLqrgWeUr4HbHofekduUZNN8vmeuEy1o
Cdj5H+ZC+8ZXNUbUllB6Kq1e0PRkwHIHJuezBHzmtxqZssKDiO2OAVoWGYUsstvC
GpybWtpnbW3m6syqTsfRsE5Yr2D3OwXt7iD+PYmcVnSd4/NLox8hzZm7Kni8ICCZ
GgfuWtvvyGNbwSg7tJQJ9mEkdfJT5zvKJYEM0ZDsAW4etlqGmgMlZipNzdfk6MWe
383X8H9aIfEzOaDIBMBq3YPtpKz143yJq7D1U8QZwDJkMndMNagwm7wdDgXytfYw
78wm6lTQH7Xmxf/u1X01teDEwMH/pdjSjkoG1j6F9mzQOJaAhtPNTcoKAXoSsnxV
HZSsWoRhkKrcOenQ2VhskChSkqGvHxnmCOxD1TgOdRt0kOAzwFZgEJG0un7hY8HC
`protect END_PROTECTED
