`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0T4KqrN5YugTQnLpi2cyHacArxKFIYMEwQb6ESP3NUskhr/8Iie1ulF9SL0uFcL
hd+qlw8AIrAxHdeAA/kMY4LQnjDwtLUXev7HabThZplo677kzNuGsbc7NX2p4MXE
zvdbSp5MVDBlBsWr2WZ7pQn1mleIkEjfV0J8jPkMtSlh5rCod/PSVXBNXdl88qRi
kLtKJBKOT+wVIo2lPE9Kjrw8UC6FyderL3IU3+kgvVm20W94y03uYnEpyMhGTGMY
8bFNEKoSDHKaP9lEFU5z7IXLq5SPfunS9k/4SHe2Q6AImLGJpFXX5JLlCPXlHu7k
BVpn8fNIiEUQjDvh2OF+kbilKN3GQiikQZWRtq3wxXrl9LE/kV5dL3ycS+6zONM+
QWrFdKUmCX6kTKMuz7g++Qlu+v6s0w5Tl7TEc3W/c8ouuohtHB2QdhN0xKwGrTKY
Dtflsqf2w0qp6EtjRSI3f5FDODq6RuhXfUqgyeNlBf8fsfRO3cKMZ4H80LxG7JJh
CowBC8tEKNB90BdYkAPAYl309c95+lCTrS5rZj4WeMcf3k7DLh3c5uJ4mc14clN+
V+hCbXX+p+BQqkTfkslARQ==
`protect END_PROTECTED
