`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8VRij84y61v+13GTWryaeKKzfUA2VjQsfJJzjHGMPV5GS3qAplGFzE/C2+uHAD8W
T4GNfIWozc6YSAyZRIBKEpVjAj5xf1rn6XcUMNMMc13E0Ka8ixdTaSRBGehv3EOD
R7kjlLu8ZpWBpAex/3Ko6kfHds9No3E1HzP9zZhfF1uReIx67qE2vc84fTNty3Xz
YWJlCy/XnAYQTpgHLJ1Sg8B79VInYf8JRldft5ODIX51fXfrYV+pwjz0Tih5M13p
x/yaiMCKJi/zbpI/fTR5kQUIXR38UirTHGjLNV+gpGC31GENfN4CVVeNZpu2Z0bQ
aSDypNAO+Vergc0oJlHsDX9+l9pa4W21PP6/W8XO5NzG0sytkLtfXN/nT35+z53K
bwybW1Mb5US7f0romuIEpw==
`protect END_PROTECTED
