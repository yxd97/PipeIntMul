`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qoG6PbeR33bvjrtckm55OpDJUg0nBOML7QF/C6uwwHAZrghQsDeZJ1S/cORAU6O
/1aPhE7RhNmEEsUQZHzH6x/qaguSt6SviyNHr62yLU5fpXn7mLXtCt+UrJTvdhXv
rPVGbMNYFaxi4V7dhsqBjYafimADV5J6I2GmhYN6VszOi8JzJ7BKbN21CFgoC3Uj
+UddW951ymGRfCa/Ph9EzRuODYu3aBX/3SUi4kGyNQcJqbvT3YVc+WqitCt43bTd
M3YJKWfgLJFfSvocXB1JQS1XMlJ/wP9rgL6cARzJyrmHqoKLznSJxIpW5fuE1ecB
H88ntC2WsqJDCsV2vzVkrI0JGSdGnriHLT5Q//+BvYivC2ZiMWVBETwm6ovhED8j
njOTMeG5kvprkhcQ7jFR8GAuDr5q5N1sK7cvxsBGZHkUM7K8b9VFb4aX1a0MqgPE
Q9QQjv1Mdp2NuIXgULVRVeZ/cRu5WWPeDgYkgbJR6VzNf9yLOCLJNKOKIi7YwzUX
bJqtuVMeGeUStP2b+cSDwKTQ5x6R3Leok48oLVUp4OcCcwJ8Rj5TV796PjIVejZe
aYcLQNjBrEWmDN6I8+AEa99KdeeV0/83NRhJxcnqfyqxqbF6DGogKytL4IAfhIXQ
EcmB2LKtPab5Xjc75z1fxluHFxkOD7IECqlSMNuuKk/km3vwCNXeBWW2ItfSKTb7
Mol3SAD5cEj3YJ/VH1gRDJdraixyMhFU+C0uK2mI6vmTcBSbfum+kiIZ+1GdrxSt
y3HWhqyCB8n40JbHRzHlJ4RV1lxpowrdUhkL0cw6Oa+StfdoaeO+EbY+Ohh+cMss
xfrDY8MG9j1Dw1+m1ODEscjXq0RReefh4tF+KRemuxX5cY+MBI3cKX2fO4jhRarS
2TKpXO3CappxKQe/pBC5xFI6XTaN52i6mZ318w7O+lu7GOBh88WUFiB3nbht9Bs0
jX7tGS7LDV3qx4ksaO+EZrTpnYVLJw/m2KWQUe1Z4hRG/3/GqKBUPrm64rjWa97H
XeIeRSzlKzYTBvPhRUt6M/4j5wnDv2wMBZmgcQY/w9MkyDKRj76limfVLSSzBMiK
0iU/kFgpIS5AahnF4cVrCk89By+p0XQcj0WovGNO2FT5JTlMMbEi2md4d0Cl5rNf
u/MehtmaQZUaPrWiHwkTEPiWuVQyYBMx8cQlXLeAhJSiU6HtdY+bt6mpoZFH1bU3
iLWr8R7sz08poN1SRXtTR05W37j3Gg9DP9T56iGxVA9kS8MidJxrDMpIOii5ruUn
lTa5D6H13WNRcfLYltTuVB1a2f1YajFYbppicyyKynpuJQ+6pRF89YFSjQhb+6wH
ALjo63NPC59EN9mLguQzMHv2/6jO9sS7kPMixI7N6JJQG84aOWvMFmiWR4uqcR6k
ZUlLkeZAUrYRELuVC2WFTzqXclt4UM8+ILhVSvJtY7ezoFjFfoE4rQyPGfcz+jo3
Dmfizw42HDjPr6xiVoPPZ5Bft6lV7IfHMam1O5F0DujrpOkMPcMQL7P4pnXP8oXl
dFGH/fbef01I9i7HuHddKyGetwxuYE8rG10v7fBB28v7rSm9RFsfYub6H34oavyS
wDWW6nuY65OJy88kpbIiA/JW72A5sYDDF5VPxBgKSvooTVKGRv1Fq9K5nKDsAE1S
mK3SLuJz1Thrz3k8X1SYE4ZIxUIsuQ8pKV9GNATmwuDgqJcQ5baLQeqEkDLQH9qe
4sEdD1xXhX5K4Y0TxT3Fc9y8a4mFcXAwEf+/45UbA3QgTjpQ+eN0hkspvrs5OqpI
UxLSFDRKH6Vpx3r4Op1XpfTT9PeSs5/eA8rkqLNJ3XLWKlRrgbTUYZj0iQEZVp70
zG/4WvSFd2kqRpM6Ou2s6t61aiWXlJrleC1XGL5SdbbBr7qqY6Np1sxRKo7HyL8L
fyT8W/+1//gy3Ew50Jr//5LWA0h8sWCe3rbHcgSZlOU=
`protect END_PROTECTED
