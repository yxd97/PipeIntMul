`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6VZ0nuUoc0ObXGM28DeTVldzD9UhqMbvMoy08Kp8uHgWcb8i6m51x/EELlYXZhxR
RFC4jupkQREA2CNmpe5apVMeEaqiH/yHEUvV6In8VzWSy8JLd4OL4K42H4O9YacH
cDALF+3+ZvaKGCm+UrY5hhI9zl8wnZaW2ssOkgbdWhT+zn970BFXNp1YzbLyGTgc
z8puLHrVt/49fu/h7p7kJj88IXo6bMBIgf+ZrHdex2cLMov74W7atLJ4tLeBvNgD
TFrG52m73lxekesRmnAyYg==
`protect END_PROTECTED
