`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SIhuCMMWOz6eEfeQgrY2+7ErSZ621h5WGPZBZPIcptPg1zZqUSZRNPHwos8RLzmS
jRtL7wZUhLWS1b+8vfiSa6kYDEnk9ly4jEO7N0p6TVx8ZokCQzeVqDYWdP58/jcR
63KTNotq9YTdby0qgdCxWv67KRwRlNWjIEk8tu2pPN1HAYwKLLKCDH+eP2U+SOY4
vA8yvDYoJpOgge8kZSF4Jdq4Ny+5x8OoQxEnzgVY/HqkQIyar72jQjYUDhWfY68C
K+89SNEvYA2ojsfxuwEMJ8bUxO5K+jOhGxY67sMZKG9Uxr4IDCTMA5Agp2qOShMB
HbZO1qlzqxjbHbGU9Lny6rI9dmotP0/j6hHyAUicu7z9n+uc0rPNwHG0Ms2hgWi2
dgJ6w4EqR2El8VDZ0RQxhHOOzbn+jV2nYz72Oyv+nMh2GvzDybwN1+CuY316O2lR
EA2nu3RfveyjbuZEpljd0bgjE2L4g1mpgZcEKRiLkLcfUU+QCe7OYfurodrrU1Pm
J2xHCClFTypj+fm5u1P+/8lyZJrxr2iql08TSzeRUsyHHJpPTYfLi99KrPCzhNYp
kPIw1p1S3tuwLKcIgZY4iodkYBZxi9a1gP9mIUystTK+ue/N46Ws5jRIHS4wLVpb
89YKq/geN5DWBqU9jcI2corWDR6ZdmAW32A/opkepxc=
`protect END_PROTECTED
