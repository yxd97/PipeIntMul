`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D0Tp/C3/hXXCl4zLBZf2IAi/i1ISQbUsyrHN+mayJs8cKD1f0w071WGAf4nX85Xp
VZDJxcd0SzLnIXoULV4qfRonNSW27kIOFvHdpLgEtRNTE0iHjDK8we5clvbiHhXT
8MaiBy9SEm5aSxUFo981DliZS2ENTrHbdfq6v+QyayJN8BzEt0LNNp8dNNWE+AHI
6c5Ev0Mkx76Ucks1zqavUEm2rU/cWB09bmOm5EtP7/iO45fLeBgxeDwTzlBJ/Oq2
2wlllSGJn7ugtKcUXiwJIy7CkvEEFQpCqJETOAtAZcdIl5Sc9j+oCVoavI7HMrPe
TKwFE8v2flilwBdItghbnQ==
`protect END_PROTECTED
