`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOqsfHKGsmj9DD2micwtUW534ve53Razg9tvkOm/qbB/JBo0jz9/V1sp3W97obHN
2VXxNzvvtiS/nDAJcta09uIU3iezmnwjGMkwjKx/IMREP96GO+6xGit1bNuP7NZU
a7nJADdBXxIAiIrzFvGQI3lNCEul5UGpQTE5Y2T3mBCoeDbgfOvE4DqM/dqgqdS0
xQyOxYbXcjdlEg6RbvLocLJQkvWOQjD7cKivFGibFRyAfvP9DmJxwwuxYbhOc+0V
LG5KtjgCx44yeZvMsDiPr8cGxF7qobPjwfW4CWpzNA5s1g5SsHH69mAKUChthGPG
jY1H4lIvMUDSIhT1Y52QtLW/zIlH+4uQkeJoDEnLCNNCThSt4X0dO3XyHhs3kKjp
lmBY3HRrTfipI75xZgJfFgPZ3yPRIMzibwRJXuZ7xu6xIlDp/DRYJ0oe1FJKwxSN
ka4XfhYfUzjA6VUeeGkDvKvO6FWO6/vP5MPbBN2NmN4LxcyraI/hmk5t/X4fNpMf
WBRByWx2/hfs7ZFb40glh5/RwXqtVvh4vmo55nQ0tkPaQyZXAiDSJWxLjlfe1XzA
gjsPKdOtXexDfTnn+uMasgR+IzNhGXpFtCW8LZZuVrA=
`protect END_PROTECTED
