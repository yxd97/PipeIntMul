`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s0tnH3vMwo+E+IA3O9zz9HSP+UKVGURc5PQmRC+6FlaKw6AmA84N0f4Lnh05Z9aK
jNkDKkMKh+llPjMhLlpcxkW2cbUVn6C4UKEePI+eZtRyRARgwfhUdOh7FsNkDGzo
JhJNNKhC00i2s7p+SdCBLryJcmfyXzxaC7uOw0GIjjUj4t/SLl3/d+nOilm/a0Ma
wDM2qkxZkBKgCT1fOuuZ7xV609e5QZdAqknhzriBgKX5PwLV50Rz7XHslR1nXbMH
w9bz97gMGv25XqMSB7e/qJUUBJMGa2agAFUL767es6L2vIdh9PcsLU3nRn+z5xwa
ZKOfuqOGJzOJWVCERHzD345udSakcwZ/Aty1naQ4nt8DH6cS6n/xykM8aqJHPJYP
DReWkPRTaxadnUCJ0E02fSyTjNpVMsePVnFdsyqfolbNy+ehG8MKnzyoEz2EFgGa
paeCuhhXHVNIaN4HrfTxEiw//eSxGsq4T7dmPPdiUVry3FjGt4RomXRvSmiECGov
`protect END_PROTECTED
