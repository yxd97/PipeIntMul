`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YOwAO7vGYqO1f90aQV9YgGx5QXgYf0GXGbwLBLGliC6xDRuY8nphfDnIA+bpt+53
rRMMW+TjVQpzboN2dwYMHj+/fiQEz4PRzYXjc1bnVAAQHOKMoXK0E5RAsJZCYKSl
TW7jkIjOk0boFkUci0dHf3IaAI+U+7CRJWHUrfSDOeUXsUZ8cqbVkxsfVwYc8l06
M1mtVn4TOIhVcTfIJHiaP+zMUqr2DmKjsGVZm9tX4pt1R7sh0D3hbFkXZ5J7BujO
nxSyvqpdIz4vDzPCFpLkUbrf+/eV9Lzuj8wEd3JIgK7kZB12LCJ5nPiOI5BoHNSU
6AWECjJMM9wOmX0M23oxCJ+DoAExk5gfq9VJWpkzF67eCtu9LAIEduCLeebvNqRv
NFbDDtx6W2N/9Sd1IAJnSMep48UZuTzTWH4c1gckAu5RK6flN4OV755CpTJmozID
`protect END_PROTECTED
