`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D3NrV5g27oODG70TNIm4+qMrtm6bRJ86GPpvCveqtRy2rGHKjBK61MppKEg8lzOA
iSgVJViXJYUzAC7vbjsn1yh4nDO1gR0TqXBHvN1ubjwVpJz9K6sfJVAP7CbVdbCJ
Y2tNr+O24xuCFmhti/vUiKnCKXDvTVmYkhCSoBMUczitpcxGdh+QlSKvqbxYLR9w
zdNZC81jefiaXgq4EZGkmpcFypbiyuY+lD6MmxpXWajH/gwvrsnw/TV7o/Xjpt67
SZ47eOBZvQTrlsm/fk99ETG9kO6JwXqS86uVkaMz2k/bU+BnQHEbrQhne0Gz/HVR
rB71c8+q67N6FmKJhPu9LoKFpShp+Tpjr6sW8eHZ38aQwxCiNvxp3NeIPZw7nYKa
jkWJiDKkKiEQLyBrguwQfSAIyKAXReMAlItbXK78QdYO1auMUXYnSAaugOZu+KOr
XpAeEBb2llcWou8KBV/uFoXhMSsBkA6tMJ/IGh7wWDYa8f6DHtyBRtPn9Ss+ORnb
GQj8GfypI+yfDDMoafpmtwUVP9iM0i7IBnetsObMY0NBJ/mQt+OcMSBf92MXUW87
fkQc/bGWdbo9dQN5nyLvaP6pQpd3yGbyTcSbd+ENZI5+kXGRXcs58ypNysr17sYO
BXsSYWrSZC4x+lsYlE0myi3ccTVnTmcqcQRN/KBQCBUUw6NoAt78sZ4sFvjmyiLB
`protect END_PROTECTED
