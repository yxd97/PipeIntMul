`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fldEXZbtNOVaJgsMT2/PlSM1pI9OrZ8RlFzb/zPthihX+ynLoMsqnjR8350Jpky/
qx8+SGF/el3pP4FqT7JrP59+LOBAbU3zwZsGwHTuJcvtVlSTxinBgnbk89rRVXlD
cwMK4p9K6IT8xFQiuTjzEvxHtHYbzK1JuC8rsBsJ0SOZ4DlflQYxdklyzVFl8k2P
LXcw1kqjDsl65xaCYKXlw2Izbm3C85yUIf8G3tZaBVHMML5yt3sLPvTciSWw77Ij
C4V8Xi6G5j0DjgB8veHh4/gVysBwn7Gpo2udHr1c7O4tUA0n4olshKhNY9crtWoJ
SggD4ciRL+CgUsBrTBCJ/wFfNMaVhzBzsbZiQ8+HN0brngp+btx2Wm+hVyxUumyc
8X+MD5iB18QANiDyRCmlS0JPR7xjeCYP/iQPeWrZlOnFOG0+x8mKIyq3EL0RJF5C
FWKcFg2lfWFv1CMtL1TvSOImaZoIvC5f2FjTtM8jK/dhht3fTva1a5wKeDGy51tZ
neQDGdLZYqKmdly93WzacCDOIzSSFmon6UfY8mci8Fk=
`protect END_PROTECTED
