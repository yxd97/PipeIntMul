`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xwr+l9Zwn9Xcdq2LlzyDIz1DGn6+8wFfYu8Gu4fz6yU5BTdH+mjjwebWyboQSW5h
xK41BQ6X82zzj9d20/if8xmhluEFAOkrmodTTbHymI6Y9h9KOOnJm3+jqlesNBas
xyo4EJRGolInzcUb9p8PeHIlXRYnRT9HuJkZbcF0tHHR8XIUc/uJdC82Z/yr1bFj
50gFH9kIo6McxhDScehMcVAVRaOFqr81qOghEBKnM81ytdvmc/Rut/z8OvSjU71h
hyzexev6aWZ/qF75yiNNPcZ8h+lnSS3rsn5BHLzP68E=
`protect END_PROTECTED
