`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pJeDMyRaEU1HNkUT0XHe30sWvOBr6g0gTXViMnJlx0m2gbpyyQUwvORMi+My4eAZ
udCQS21aXCUb+wQXaetJS/JPWewwrkc1jdapwM3wDM8EaiOnDk7fB0p82+f2Qr/i
PuL8d3/pOoS6weNwODkWwzpmfN1tVcoxjgwOBdKM3JsUh2WMyqrvsAmhQVvKNgb/
Xo1CIAd6ZgCdrMxKdJpR9wgTY9s+KTH5LP1ITJkaTMSOI2UKuatrhGiTpm8Xw+bk
KS1sPvUvOIodSNTWl5s3KlGh3/0Q+P6+qQ3krivq3pMF0/HxK/iIvE5Ha9IMuHTD
`protect END_PROTECTED
