`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvrdJ915/A1X0XYUzLqWJJDj8scbtGmavwNvdB+PSMNAke170JIoA3AfpvrmWafP
ecrv03cwNa1KtDHsE2MWC2a29lcB105UkEDFwRTaxy2jK6QxpZ1WDyxHAJwYUjzV
4dmGgsox3Cifho88vxGhoBBTNAjvo4x8dXu8/Fy+tgX2MYWOOopLYeWkK3zPCdnD
xaKmdYdDHNDx9DPgncDniXwNuq+xionS2Nk7i4H4IwBudI21wRD2xJD9pBGo2obu
b0bFZPoexytyTpOLA+0ayvcGQYtP7ADJLXk9xwpHdh61iL8LWVji10fz3hSsigmA
w8mgA9Q5IHY/h4HDVzd/wkJTKVnQxQGkiuDyWvuMpmANvI8ITD1xnya36TgpMBxq
`protect END_PROTECTED
