`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OWu0bhge2HuOtp7k357G8QPgl7sH8cPyJU1m70soLJpIoK+ClX8Gfdy5rR22XXP9
13dv8IrXtKW9q1pz2b8Ann9e7QJSEShndUBPk9VL6yGlnJIaMIZIXeoFUCDQzfqM
JIkc1sbsMsYJ4VrZeWS9mGfulvi6A6zJqZsV/1J0aw/oeqXEcpMw91859PnB+Mfs
cvVndQGdFB/7SpWEmUhp1N5nVW8IpckbGL3qRRnpPvX8C43nCYhuNdqkuq/wmaO9
RRc9zLY9ZNqvjdy6lMiFeQ==
`protect END_PROTECTED
