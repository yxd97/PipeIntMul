`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ma1BKZI7nO1gSgyj035YdrnHYoF2t3Vzdd4oyI42n7Z62lCCIRp0+5Pu4Ide+vN4
ZT70Uxrqtlq3OT4+gFu4ZK8bWhoBc8DazFG6kSu4iBGhYTrel3p4kkFHxP2M4LGo
Gbez6sF2UgiQ9bWYFMdeN/esb76lovwznK7kw+n82mcifPBN8Nd9ArCaZ7xBWCK6
qXWdVhKUmjjA5183QY/ldWn3vu5FOX7dC0DDHOuMVwgf0kK9Aanj2F8MwcBErO50
`protect END_PROTECTED
