`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tphbNwJQE3T8j0rH9NaDtN1ivSL/pVkeKgjaRi+4IVYLsusRuDT86WY9fl8MAg0n
GaMyKNRVhph/mDgrLScRag+BSX8jvajihZ/PCeupKKNu4FOqBiuKJkYn2lVc00OJ
/EL+M/DEMLY1RFpqZjm7I2PvqO6xzo9KbpiABFRHB4hpJmnUg28lYTwS9BKxecot
Dgs1+EwW4K8bTqsIdG5DvObK4+cuUOUbUEbc1KXazPJgxSDQ5xz9rxf8cunmZVBn
iS+YTZsVL7XEaC9XeRbVGfaPJTx5zcqg7UEVo+mQdC3lqsRShvd3twg+Ja6pSLEG
lFGmRW4bgyeokOvL4TeojlW13b7kKod+gMe5j59SotfUK1AGRbMuIYlDpSOD3aC9
MSBDkfk/QEVGFlUb84YvF1QEjU1L1PBIhQvUOs3Eugk=
`protect END_PROTECTED
