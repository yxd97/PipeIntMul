`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MU2DOHvVIp8Q0hHzOvkJkntabl9HL71Meli1wVgLtT4r3hbi+wqUQjgKzv0kA0r7
Y+yE6I5UD/IMDhH9WzXMqMdXyk31016FROdzCZz23H4aMGjNwXI2893ezcOkwxaW
GzeFtZURL4d6swn71gt5RlZTwiU2XNr7CL/gqU6MmKDw0pqlxzhxEgxOwF2BBA+f
kx1AFsgofRvbM/zqPaJlQyE9EQf5inSQEEotuRlD35W16+M0TOdmzswCK+qIT+Sa
PMiS3kOAO0sDgxIPmXrWlm7tZOcdwr4lW2TUXJ0pp5QiUTIGeqcfXQ35N8fYgVuk
VfS6o/phZ9iGQmhelFPNCAznPu3ffL/IlsBF2jeQNgm9boXYx5Bdr9jkOlmutUru
0JWUgfkG2g/CTplxq/cLwAOwN7KMO8rsaOOuNWaM3QZ7DFOFiCOqtxtiGbtq5XFM
AMi0Oi0sIg5azaG2D2kG2Nj5QY8Jb5dEObuaGpihhkMZ7biZpcnjnX1LmPkOhbY2
`protect END_PROTECTED
