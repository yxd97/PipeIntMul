`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K4VsioNqBAxWTyFsUu91PMjPj/aD/tKWOdf+dxNNt0AZY5riqb6KrKdSpiseKPa4
f0+iKGRj8Z556pTRZG7xr+FpPKysA3HQe1qfE1Ynl8pwo8pyrGslrL3ckxYBdtyB
BikPxeVRYsU7kLWrIL4RQ22bTahpbGLiRfY7JH/1T/dJSS71olrROcRFasvcyUi9
V67V8kI91/6mcZq4cjKJThQXiRKQDlY8xKUPyCVe2By/lrqfSX2FXLbwuxR6HoAo
u0a03yH4/T4PMAQ4VMcKuUuWCnZYrHf49St/1+aIfUC5Iy+cVvPY7K9Ui1QBz7pn
p871GF8Fun2K0YjZYSVihmYNCv23ilFiSq9Lz5BVkKrurlYAUz6MiX7R9egt4YmE
w/vIOkA+exsnjhxYh+NWd5j9w9Fh4W7AZhLjumYwL6hVHVudoA19D9FxMhDF4QQF
XH76++cI6ryopUFxMMuKKldQZ3n45Q3v+9jKy9m7SsXgbYJMD/oIW1V/+nc9ugA2
Z/nlpxTc6abJs3OEvr0uPiNdnx5gNHEe5cQoT8WDfSbiacSziBV0DE9nVBqEGW5a
OfmmboXpzkgOwl+zKCqrGIErCHjFRyo07VujT0tX4WjlHEDHM9JXqnaPX/IZxTC+
imxdY8RhkXYw7zha81IdWrVQXXTDE3FCOAzKESaeCrQ=
`protect END_PROTECTED
