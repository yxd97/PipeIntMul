`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+lNTX4yePVe03mS8Fgk/OQazxjGh4D1Z6YilUFZu7Pmuhz226q1eytwDqum5j3mm
RVW/Oh4yqj3xZjEbRJUA5kK53/zR6UpVfngX+jKMGHBLsa0RzqsKvwDZTZXNbl5+
NuTRS5SL7TbCB5p2jTtDJBsVyKU/U9HGVo1FfapkPuT2yb9u/EWzwdV56SC8eu76
zodxGF0ZqNHpNgO6UQnxVHkOsxvt/i0pZabq8X6v/WcyA0Ruf2vtLPYAq5SoA4xK
DE3MJ/BR0HWoCLiZEJjlcpA3L5ieRWPQWyKc2UUFvpD7GupN3c6tA//eY76L3CxN
OUh8gICvdyPZX8fARwNIyrlTdgrIfU28/rChpEtlcoA4hR05ExaxpP7GmybGEyOV
n/B9U08TTcLNM5LdfEfxBXYYDrh++EjHwpt1VbbXPTiuArvaInNFR0/v2cVYA45x
MPIg1ep0XTCf7eONh3c8dWK9FtxBo02DzUhQ53+PZt8=
`protect END_PROTECTED
