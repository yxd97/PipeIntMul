`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qcgRX062/o0xu0aV3sRP3855eeKzFfrF2tubV2ea87MyyTKVIoOWXAqzGS1CUXjm
Thk65qpKz2PXHSdELzkRvmOD3lTTcARqh1xMZ50Ei+W1YQH+w9uEaWbKKdZMixrD
lqsvK0fN3em3xp1iObZZkbSypDWPbumpUci39wBGQ75YiTneIZ4ATaL7ttywggGd
Iz2Edh0jpWIswTfHjDK4REBXaoyq6a7iFWIlZSDrPxk8LxX2abfI3cbcCde2v/5B
uZZssHs9u3XzJKTKo9m8mblrZA+FxdXk4IVSlp8dU3luLbvKXC2YLPCgxysbheXR
fwuSsL3NHdzz7T7S9Xt2AUrOR9t7S3Bia/56CflKv275DZ3vna3Ai4H/pDrwXrLP
9FXDhzSGkzyNaqvVRD7z2GKthqZiQlAkHs+s9Rkx4/gY2jL0pUKugDzMO6yMuZn0
1XLpfYS3vuUJJSLlxYkyIV2nigId++vYg402Iq5B1U43nrqA6oxl1uwFrxPEzyP/
IDHnkm/ucaMRFZcgq2N3al3kFc9emVD2VKm+6CrQIZ6gDk0dVU8gdZbHdeeQE6DS
UE6OlNQ6vBL9xa6a829pbCmzVsv9mCN48A2nBNmSDGjoXXhp0T/HrBfUDrziHL57
FhTqgaWXBsEXNo52fXfjcIQpUodQIWrcmmUPqg9hZ/qr7ontmWYOz1l3Ybk5NFpO
34bCxltOjzHgyjt3pXylQBaBQN/3Ex1PcPJ8NjxF8eThM+OqPftzrSgyU7W6DhLR
Gla4+v1lA8bBM17j7LiLTdsNZHEN5zLFEi7rmyoUcqvDfglqZrPAXj0S/Gf5k0xU
roN+wCdlrjoE4sPTcJ/40iHFKSknxkBJg/gXAE/p7In2S6Ynt8kkigASv/z0R94W
0CfFEXhd6lpEnZr2KRukWdOxBry+hG7nvSQ5CfdxaNsfjxQArWgX27K+p0eqnWYC
uhTG8cwhDLMmjmSKUPlxkgdzFHj+wqZ0sN/RNIecZXli0Pl87gIzASE5eQLTIlp2
bxPZcFa3MMsodKlYpJMPmQaq6gEEbNnhxFLxSuAHzAUDbsImVwe3euu3Q9DYCeJ6
hdJegN6/Y9KCIDaki9XMQfP/MXSj2vGEIweOFBJ2WiIyutUBZKOS+BsVocWYUArp
0L66UVRk5PnQcZZGcie0ihh9gGakKeUWafjoAN94U35AtXq/Oh+2G7n0HWo8KwXO
tb/LAhB3+huxeU0p8iJjlRGiDebAMM015hFPzEL5bi/NE96zRLs5+Cjhsx5P/gwf
wNpVks3XwpvTVsM5dR+FK7Z2LztAF8ZN1oStQFQsSvgOcR/2YpPrDAK5ysroTw31
88U7r+ZUwUUJVRMy5mC5bXz/bAFUdG//NbSeoUzy66NWAidGBxxOqhUrE5nLJJXM
+7iPwHMCkbCR+cqWSmxqKbGIn/s5gioKXA3fnjWP1FxEvZBrADH56mj+A4CYFktk
dYZXngV2RY4EZOXpWYoqtFYdQDZ1GH3/jMxHotJLHWSsTWEx//DImzl9YP0EiK3O
niZgnfZihCnEO+4WMxTKqa/EDxDW3oElNm8sfzq747tdu4P84Dk0lAtd8CFrwUF6
du7+aON1K1Wpfq/FSynnDqdNEOF+OJhwj72XG8d+rD0BiZ/tJ7Dl3GQmrACM81Vv
QW5eoXAxk7T+eI3C5VN8793vYekNNEzAGc9PaTQ/uJCP/3OUHkaz707WiYius0Zw
rHkwmG5pJbgN8e38LKXLW9IyEY4IQaf6D//HmvYTuyKQKpXJRAg+O70nELFGBfxy
ViZWxWrlsnvh2pIvFms8BOjLiOIlIR0zrnbH90QvuDTdMYyeevxsUUtbfrXYUunj
Jm/+QFcbl6QlTdbDw8l6+INO+JTMCxR1fABRMSoQb9XVEcrOajwYcpS9Hh/oKMIf
jK9+bCvUdPS51tRZJb4Rqf/YbSOEb7q5Bj/LSh0NwIM6lZE94NBMavg3IpKCUvKc
QxwmZT6WU6JyC0frs1yC45ZCScC+pZeqIEeAwTs+hlZr/4rOLAT0jnAr0maEjczq
GzW85IqbJ4X9hSURYt8ywyF7/lcD6HLWWnRMmrpDPrp841Q9DsKolxyG/PDpHkqF
PQMbgqrJyVPByPUZApVpFSe4+wFOVKTb95TR7LB71Qby5eEK3anX9Hzf7jB1ItV8
Aq9eNOMGEWL55VhKopmK8myJjlv78JUAlrz1LJj963mLiBqe0Zj0spDJfEbxjBOI
1ywnIRvSKUaZHG2CZiFNik2GCWa+6a9N28iKINUacLbB9I1w835HTIXKjK3AsqAl
/J0I5A+vIQE9KYvsiR4EYolhT1ld46C/7rlw/SzWtPm0F7mX5x/GnDRF7BKU1Qgy
rCTP7lL2p8c7eTeKPwNMty5e/3oWX+QHwNfwL5hi8cu3kM+9Gj8V+xp+cPUhdgXa
Hjz8zhLieGMDZshyPOb6m0KbMhW8WhvYNMJKo8tPeQrX8ZMbHxNepVmj5ygbHjjA
V+60kSrSNkTzSutEowIxz6wr3Ok33E5RXaj4SueU/5mh5kZxA2hktZzX9NTjWSdx
9WaevvJbkmJjkUzJqwRoufXjJBTDyrYoIOEwMPwnQflgB4D6AmXVQaW3re1+Fsv9
iVmgQ1hE3L4zGVHBGXMifqyLM4Xa0vJmIFjBHJFbZfGpiUsgcDGTqu7oqSZyazNb
PFRmLp3JJPm7INdr71KFnF+riHB/7cInes4V2DKMwEaEem6YENnX1hmXNsatDIWo
WYPk+6oDR1HWxlM17+PXAski2h9vk5ZcYVpqYbmzcACpQ9tpSIfqBAYfgttlAb+K
HzmTzfh8eYcRgN08igA/XbOYDUduzBXDbJA21tknH/ocQ4ftV52y7C/0SfAdQMHv
X/wwm+7bZKvQzUnjKp+dXnY5yC46OtNzHZ9jIOi2K4S7h4hA8cadDb13V3t6hk5q
hvrnp1/hK6OHRhO47HO2fTL+Er2MXmnb9mtWzkCPySt1Qshx08jqaDQfDmgMGMVN
l4TqTrULGh0VaFIQ1RUxsNRsjsJCkMRTk6tVLvBVEKc4IHh0B1QoCyavLjmxkXe3
K/FLX/vssDcfxbQbMFPGsAIhcI2pwljdkVU2RglBDNFk5xj/UKi/VgOKyYQ7jS5K
KQSbyZ1zdbD1YbU94H1JPb9IudbYro7MiYBZtyJNgfraRjqn1gL4A3F7yUwmLVBt
k7JvytmBI+2Nf3B0YHYpqaWZF+zMhCGyo4DCrRECmY64rkP/DICsdpmxjebVLgys
2/dr9kquyp05xNVX7qVIKklEwzt9uzKtb/QgMHxPkmRXg8RHbA0IQUNd4xuV/sMG
RRjs8r5FEEsqJackC/QGj9Q8Zy2OyV64IdSqb6A1GnNEQHqkJDNi0hOMXkyeStrM
Td79Vt8WWlyv9WBPUqNxvHpFGOoVjgdrMOoqXVPAl//jMu+fVLKBL1cknBgMMFRo
WKLpf6gL9MfxtNFEmUV1oHgibh0CrzxJ0kJAnjGuB/WEf6kdMes99ybBwbl2Nziw
l+N7eP0GliYm/0plV1bK4yIm7DxejpzXudQeej4egeHDA15MQ4OPKEYS+Q8i2xD9
cOZNldUGP9tBL9kSV9Ke4aSA5ht7pZS0cpu5ZmUAZ2z/sUHx8Cxc8j3zwi4VyjmX
oBANhjD8xSiROq7dCVT3pTwknQt++LjHzJSIcHD3jEKWeHU7iT0Lkq8sz5w373No
JRWwprUqUyURYYVxg2mFCOa4mx5zIAnllfhWf4n76kPNSyaXmNidTOCikWWkq8Fv
EB3QjwEMzQQRhug82dAIqWRMKCGSKxK0dvGNf/2oPD2NQ/ZiNax0d9npewp79DoH
mXcO0R0YWdJuYQ20qeZdhuajCPAlXaKYefjvrtld7ciFqTdmpXvgythk9yhFQ/60
I9JBJr81SVdidxD08n9zM7ldHQCqgq6ZeQ5bg5hXDRQtLZsmeoEZxgnTm9DcWL8y
LW56n0Ml2971fqrUXUBXFsblcfAB/3QuJRngkcDZwXh/GYtVGlvKQmvXxRODSVbc
8QbD2cD6Nd1nFUOqg+K0NKzZx6NlCqwflUhWlu74O75+puGYbRzHROOhsotWAa30
eOK92z+AJt1Uj882Tdv2lb2iJZ1RiFqel7KOdQSTigdci0SJD783t8wzwC1emO5L
4+qampvqLoXIr0kTlvFCbz88vHKNqE4ur6ASQpFG6i22PP+S4j53CRNIjhz8aZvF
E8pIE8X13cS99HHiVYo3UXu1+O0xP96n0vlX8gR1WBB/+z90sLJPD/y5h95dTJH7
iqaYRP1pHiw0N5gyMTHQ5FP/OdVN1vDwT9A0bTdetcAg+sEbt2D7y5XdfgEtg/s+
6Xsp7q1KZrRkGCdzxR8cp1GhOd1hzY4QTPTE1UrUNKlOeqQcYb0Tcv1w1u6H3Wyq
5ULO0NiLHjTXdw9ueNwcc3Fm9cl8g36Kfdzzpid1pmql9HfViSvRsgEw8zuLLxLc
D/hoDZow41cE5NiYXBxQHK82UbKS9ukYyF4U/Y4GQFyByWKpBhmlWjhHYMcxpD3e
+c6rbYyC+f2i0QyVHst1xpAaONn/FjjkaKnSduAEgdBhctGaUwvch54uUyrXGLYx
kKr7GGoDskuMeOAKnJBXu/AcpN5zoISy65BlrS+TvnOvwNlndPnOWXhVymIRIfjg
iEDtmgF3mcmOmdNfi+KeuUP2oMpEEQ0noYU5xb753PAQKXjG+Yri9hJEXg6PpLro
rKsFxPA/hIFezFa1kKaSIobO3UHnvgDOpwiHKJv0BQpGbCPY3VaovigC3P3W6oee
WqhSxaHNleMEqei+tGhENrjECIK7TyM0mVb20LNnHAO/hZV6T+4gcdyrNMRdCoAY
5wawi5cL6GM5SBkQ5RA27mUKM4jy0lFmHmPXnKA3otbK/D7Bl1/PGShCD8Imo+4s
6C/pHCBt+17T4BFuZeai8I6r/Gko39+TKxZzoMAfZtdHv/5AF/4W+Y7gpmegRoZk
+RRVOpfCaGiwdA+Cz/St+l59Zp8kGzvlZC5Se2A4HldTSO4ch3fm7S/vewKHaUxM
kV88d54oKFTq4lHRHWA0AhUUoQui7VeLwAcClD6hlT8SirY+/sbirFILl/sYTBV0
KuR7Bpnu6STlEuT07pIBJzsmRN62VZQeUG+i3P3tZP2TOqcAzQgkSiVmbi0AWWVx
kpd0jevIqqyh77ogSPZDUl3CinpJVnp9ORIHV7Y3vaOxQrDek2rSyQvWQDUnJYS8
9L8ZQODgp4/U9t4k/giBBqdy97PMuroynjU06curGwJexK9tqwnqVtmd5vUE7K/R
W1BfMXaLmqWrOUfe28hNO8Ez9REmQGiVCt+0NHOZiXJm3MyGG0YZzZVl8Sz2CJy3
nq0kMtT4C47pSTHTfMUpEAWUZRPiAbG5vG0YCK/IENvgjrMOYN+4jTv6ZoDXFQWc
5S6lMwYeOEHjD6mkvJmJjVkrvFPbaYkPaP4EoBmrJPAx/H+MSUTUZZpLxc3+/duw
ehPWAUfoAEryE+SZhgFAPB6fk/KEQYRCZmm0q3N54BUqYAJChioA6baxEU+1T3IO
nOpEXlORQcmOF1cMJkNHAqkIcEEtKnR8Qknaif9C3VIvXARAPSP+V+ZSns6tT+Qs
eaGg+YuE/aHuH8hv6uH83bBO4SJF2tmSTrKYe8+GiKgBWZixUH9IKdnPrkMgqiHk
hmjGB0SZlgSls2EGM0eQzYZah4shFrQ2MjWRgNJQ3i2HKCqfMzdYeD6HBxERLHOw
mFcaRqMZkE/5KP8s9IU/X0/sTx9jGFYPmFLy6wA9YYc8k6Bswucwoqh/UjwurkEV
7tqExj14bk0sQQnx12YDw1xkOqN0bbsctl9VLXYrNYQzMNp4EmZDKRp2ppOWLebJ
t7PCFEJD8CTt72ajaEth8FeO/Zdv8mOkLUBeKGslU7mif2K+JZLkSkDLPAEI6h98
6xzOAddvFoPYwfKyg1R3JYuBrdsrSjHBd2ULZmVGH3ttjHYJU+RV2shMutN66ubn
672xlaMrw8nyYZL/ncZ63xYF4rXradoKENoHLYweEa6KhPkQJTBAitdU3GEP80zs
2OuOl8ogP6cWDm5qC+Y44pZo4U5wUIMWok5mbXJDpUOcj9DEZd6gpnx/bcGl3Fsx
dqqsbikCu6qr6w+MscuRyTcP12DTduY2XguS5//doX8P3J3L8Q0/MSv/pLE5mnAe
8wWQ9mr2QlHjJ+nu9w+drLRdgNXLj/M1waKvCE9eQI3uODrhA2/CmIb8nlSoN1eK
fijR/8lkjUBwke/g8mUG0DJwQ6sE1ADgsOC6SKhKW/4q2YYC6/O4DzwkeQR03ltH
f8C/I03G9KsjnrqWJ6sTOLTThyaKJQ2dmEHsR4SRO7NQTK6DfUukjfqo166J+Pea
OXDoL8+X6HfWzbmOrY8YG1Q/kHbcVF0s0QpfZCN8p1Tv/eWSCkbzX5At3DhhKXxt
Ah9kYU1vPY19KQruRAsn3sFPG96549gjkv+rZinjve4JxQH1ggJe80K4mn23H9w3
WFKJu6LKzTaTUSraBAMzVGNfpBtXlehVPjyp5AvwTzD1Wv+MCo8+SM1qX1y9q6MZ
8nB5bMsGfwx4REH7cSVcT7SkdM3dScdTAb3xQeS6n8U+eF8f7WFkvaXVmUOdPkyy
iEv8rnpOOzlepdfULnzQ4LeTwVXav4Ag4erVy7rhvjs02D5Bz/kdlgecWZlmnK6B
rjPB+GN8n1Y76U2lIoEMhL/FafVGEmNYA30XcsP9FshZ5Wk/33nTZEEn5WEGLIrr
sepGe0qaj8vV7cBFB2Gq6xMwucFuZhT1pLJmBu1I1/X+1WDT97l9Kc0hU+7MOpWh
+8QYtE1+bmpxv0YDDxwBPG9d/peqiuZz7/xx++hKGYn6FY5CecqXst/F1uR+ZbOo
r0decsAzao3aOMPDPd85QdjP939GBHDLqoDRoF9a0vjSnr4qQr6+3hfojzYwvchT
w6Y6MJrWugGejYJi8rcFSadi2xDKLrFizyBU5P1t2GPINtWLDyv+UB3/5Up/Kpmy
1yU4awLSnjGTIFxoqcAoOAPVDn0Mnhknbu/yIpEKtjHbY+SIhbijLkCNs3hlftJe
LHYtaFEupsfVGl6Q6yuvw5pxELtEgVpsj/IZvFOQYT8fgXpOXVmCEsFEDOLhGhfw
AeC7UVHyeYkq3zFWCjVejjOsc/4pwrGNzrfdu7HLYx+PIpc5Aau9cW9ds1YZrrwq
O+jad61O620lrn1Zs316hQRF0SySlKT/kLgNzroNJRGS5UtQXma77gQlEjQzS6Nc
3kuTfY3Yy5VZEW3tt0IXwmZziwDh+0q9uZcD5xj00A37ZbBunNmV05AzBEKSIQ8n
BSW/d5LaE/p8GvbDCXd9DHx/p99D6X4h58bR8PjIORZYe0SR1KY5mLPUrGSfUA3A
5gBcsP182S3cRVTKI9hdD2Q+ftPOMYDEtPmUN+3R/SlpmuEL4vI3jdY1YtA2G/E8
QiEijBi2Hz1vvyu0zvaic0R8rx8l2Vxtfw+OzKR0HEw85rW8/nBggq+YAVNv1FPZ
f4aFjai0PzJIbDAmqIbHpU/vPpv+OlVzz4OkKN78E7tF+Xg3p6yI3S2AcE0ymWHA
XMnu8xu7nKZGNgWSbK9cJe5eE1+bQA2nvxtWW659fsqsQJPdHiQUO5tmk9i5Il6U
WZLxcv/ivk1im7ap4KuqX2br4p3xlYQTaWA6fW4f0H9Fhn2nK++bR7Zot2qgHwVp
4CmG0rqg4rWo599UHmFRtWrYXTEMjYbpNtgHvXyyejuNDhJ1dJ4Qq7/8U9gHDd7t
qi0qObMOA07nsB7sOSQGx5JX15jCvwTKIqyDcW0VkRnmKbZAIZys3OWomtiKELqE
jc5gNOe1sGEQP1ChaDnZSI2mLzVoGjtLfTHLCbw7/lFZNTvzm+Pk/HIk+ARmuCDk
ZKFe6Lz2wcWHehVxPoRRVfm322++6rHxvfifRJes4yBaR0xMsTfSuJ/cz9RLGVgs
7pCxsFTsXHISaIk6ya1edim1GNwhYf7NWeDW+oe4UAI4RP+gFwh2FtpfSfU+JD3j
UNbhb/78/G6exu7iGBmLFRp6MGD59H7xCE3gYMTJfsB/OGi4FxAZzW2tH/GxIygG
bBqePw/kSVs6tnXlGUI9+aPDhWOQYefsj8qNAlZzRvXw8Zd+dZxUgYyo/zkYTcJw
XL0LXkqFvOAfAXbMzUm5PeMNLxBBYiOHJnk6C3TrzD1kIbxjWLkRrW2O3DfK97YG
EbZ1x8hqKiqtwXn+jUIEYkKPkIz1Ku6mmoRsMYVSQv1dImK1Rhgmr5qSgPetArf9
IJp6uGvRfSIK5UwzpSpfa/omaBHP8TmH4oY8WpghU3nY2N5CWJ0PlfnmuQl996n1
2jjWaCV78uwHnyNddOHGdr19Scrrs9gh2d2/44/FnQXtRgQ31ExTahNpenBPSrt7
lAnDvR0sAPjyMc0emIgiJGzUVEdEUapklMqAu4rVpwRBjMMAnnUliTxVbBJHSNGF
LBB6TD3/l1h21ZouRjMr6jP10bBEnWPoYlGGmyNvjD/rqeTtvZ4r8YUUGvanzP/z
+KaQNpzMJ3pgyTZ75eslcYNOhfnP8Wq6qxHTx1fV7QwrERHy4cNDn0lPEUrU7fRi
wZyWOFVIPMbOaVEcJVCEKsZq1Pj7tKiyl3j73G3TdFHBP6dB1q9Iz8yZuOOy07cc
C9dd65qy7kB/nCKljcfiB/6pHC/QbAsERQ3gqrO0n68NrXUTDuh5R1aT0Cfev2ok
jMfpYXzps0EhZ6sWy2s8SJrN/H5iZcLAEV8/+Ms8sSwAJL+vIT0wRupli4qLPfTv
RH3X+ggz7BmP/bI6lb0lexJXu6lGYZY5Vm0d49Y14TA6XNwaMSmaYYMlpNqmz6lZ
BYVY3ZT9PI0fok/RGUapNr1of/2mQ+BlN3jMqpTvYnUW22+WXlgt/vB03CosoKxI
BoqOxfQZ5hxzDqNrZhN60BwStLOiwAmx/w7cFpJ1IBVv5Qo7D/uvkYxpPKWznMzh
nGA+8h9Bq0zsus9VNp/0qKFlTHYeOPYleJTRvm1ZH2Xpn1QFkPw5r+webs/STVFi
Ypjs3Z2aZTDdOXetQKAor19hbuiUnRc/jQRHuHs3maa/wrmLm43xwg/PIMwlyszx
8luqJwIfpH9ToeZs07R4UI7mJKm9vc8zTzkklgTOt62Ajm/hVMfmZIUrucYOvNIh
d5Sg6sn4/Il349KrL8LX0By+j9oCBinYpJCrLCqbI/QiD8Qt+kI1NqxzfS4iNis6
1t0uuYlxAV7UKI8vps7xSy4RMhHIA0/wa/4TvL875VXdBucy6B640ibDefUoOFF5
JdnI7AdmVHeLj+Ot/HNkOrw2l6o4FF1K+LxJOFmqsC3oO/VfQsxtk8fcfZe0GHZV
EKr1GyyGf7FHjWln4Sjgyjp0U0bU7Xm8iTZsLwz0baSTkoilaCTTpHLyy7y178yy
yMGxbNlTGL3xXqV0HmrUsucfuMlRLTwu3Jt4oFEGqpgWaE3qRPlU+bALxFZ9T+wV
A7EJMYkhmMREucayZzcy8zo0tMUHEFHP0AY003yTVG9MZRLTYTfTlncxWski46/B
ObMbTgIL8CoZTWeAabThwTCPgyV+PNer9Iz1SG55ugdXeaXg5AUyouaLt/ObKmiJ
lFOWFvoZMROosWcnOYUIfMXV5jgZe+SM2orLoTVMUwnHUtFGOBj0+h/ZUbc5B601
`protect END_PROTECTED
