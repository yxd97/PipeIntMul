`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JYwFOc+2IMpt2a76V0Is0sy83VunkivCYLZfDtAERAzeRAWecxDUScUCA4R2JXrp
o68jnqsFthNFKn8d6mbZsuVc5XtHCaiIGhiKOOh3yU4t7MDjKT6BvSl3xPqGSRfq
j29Kd3+q+sSDAE0uK8MLNbGlCg8Z2RHpVsZNXtR2T7X6oGOm5iBk73XupWIXCQFo
Qx5nh1BSfDZlmaF7x7xYG/4bdmGVemNRQQocTPnEpIacwtwAxN1EVFDyo0EokkEd
94XSAZmBgukDSIMQjbzvLW1FjGBXmdfLWQ+tpuViMVEr7WzIxJmP6m5KVNA2f52M
mcajf26rAnXUUK690XHtL6KTrv54v744d7NZ3iZIaAu55PG7RQQODHfvTrPUQDjP
9Fr7+Rp6dyvuJ8ZvSV/QKWFV6iin4nYC/vdubp5MIAgb4UhcCpXmJLqaKYfXPREd
Cs4stfKSRaNLvVN/z1k6EKahKY4H6OGBPm8zsVu9QAkl5zfJtvXjAiOYK8DxsXQx
LsU4xMyHBzdqlndPCnJDoTQb36EvdJB9UdC7Ib6C9n3v+hiPUjmQosdby3USy83a
oDrH9xnjB41LicCJ0gK2SKlz/gXQW5BDjRnIqE6012U=
`protect END_PROTECTED
