`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNN/9FXiLG54NSChZl6mvJ0SAy3OVRtQkemLYZgGtpPwrj3CATCkw/aUX6xPIFwJ
mEUvw5Qd6xzc7QfiKp4DNZm44WL2XJhypa5vxKV73pbPVOwZ/ftxHMfkQzAl18nU
qPbfmeKS0GEGi9bbkcFHKEUexI6UWea6X7Ycp0sa9NuwdUPVSkTgEq4NeKydsA3P
+gODRuc1IN9AqzmIa3eCV2pFRT4wXBOMzcELL/gx30r18vzTPJRxybjhmsbe4HPj
cmiSkHBgiiB3FUaahrc66A==
`protect END_PROTECTED
