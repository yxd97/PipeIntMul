`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFeKJuVEDfVZwYSVxPFhemX/JElKEYz5gx8zZlpC43oetStlrhcmFf0Ojdm2xNar
I5t65Haast/RMFlf8Nr/rptY3lmEqVs3AIzhtPN2r7sGwMQk7CZbhVa6FTIqzVo6
XWlNQxKC2b80NJ31MZf2uwGSQkQ+v2jeHczY+3eADBsmv05nY2wLx632j9yqUPAQ
H5omIpLn6evbBdU1oBeWryX5sRDzEqbG412qUXWqcPYmXdtYqafWn3wUT1BT1gCr
RWFiAWnH8BNjJNt3tvz2ncmIqwkMQZQCuGHrXJCivLGCL8nuheb7oP0+CjY077Ph
`protect END_PROTECTED
