`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fLHeRp8jQMES6DnQPbSDL2hPyAjZPM6Hy1Q48jEBX29hmN2AFpOBGeLKh5GWgi9V
cdCL7Mym96zzaDtHgjpY7MNx3pxjR7xg9rovbBTQwzuDDcarYYgbpLFBuCw8XM6I
FZELat8LJPy+HSGG2nC3li4DxngZ36sQ03aTlp0QHjET1N2wRGZSVulSw+tVHHSa
wv3q5O1ozsY+hrVFt0ti29uWhgHA5dbmEFiqX0FUbGEURZweP+fL8SUt9tYl1bt1
FiWm7eo7tZC00bKyz8n8yJ3jwcEvch7b6nYoJNG3GtqKu+SPN3M7lddGDTopMUbG
nJ/9A19zUYYmo/9E9lIGwg==
`protect END_PROTECTED
