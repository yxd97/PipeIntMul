`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2DFBYkBe/OcKrfdfq17DAIaU1McqbGeTf+idIMIxDM+mPD+XGUk4QvZ17mbbhxu
XCZkwrla2aM8f33cWLj+eGP8BQXW4+X4QwnUvqdBkfNlD7lstVbHJrWTr6PNf7Ug
ufDMak0kxppZs5QUqLRkPqHagRPfddRx913G9dUKVx57l7WkKFFpbv5FO2sTprkz
v6ONuCo1CHge/DacEG/mRB7aHYqz7m02vKLq7hBz7pIqdhdMKhbKEznIQdqp8hUN
GcBt08McAJ0TsRyrvvi76dliM2O90jmJIgutQlbVPXQrtmm14YbX6m+LzEpvtTCO
J9GuLhloPSoW9c+k2usbVu1Zb0PZosx5iRH6pMhWxr40l66TOhWyyjKeY0XHL8t4
lHkTaoqpP9/Qrh17bFJtuF2DN0Q+TYDD0XYJDlL/T/Jd19xhz5Z9+1oF9qFoaaHE
qr/Bc49vmwRvTWqc+8X1AuiKuKUPNZXj8HqS0L++V1UQRrghXSvLV0q/Im/f/cWS
ubCX3xSfF/mooqr9AsOrx4g2WFfZJeZt2S0a8eg/e4fPgyfVp9V+o8zFWTmQSLo8
3PhfF49iYpDAm6Rz7t0XfgqVb/4EGlo7hEii5OiU3sdLWqUflwHwWzhv6AxFjAB/
tFrLgZonqx/iNGOEs+YszugDI7dWNBNIgde0xD4e88uetdIEzAUZT0qVrknygXhX
pxxb/DHe/MVfYH75pHTTm8wH47Nmc89TPPF4Ak37QbFFwIH+voPdYGVSZSR2hGIn
UCuQXstCLjHH8IdW4w6nHdnQukwK8gJ68Ab0Bb32VnPKG4PswPa44Wp8OaEztDqn
lH4MMkpGrjNA5GwdKeblOpp0NnSINcylmx3ycJdh2AuMvq1mG+a13+25foXH9ZdP
kOPkMEg2wJbgeGkJ7Snv8NOjwMBfK+9ie8/ti788Uf2V/VYQ5JccNvb6WQp6Reyh
yrfCJ34uJ7hMfAax0Ht18QvMlujq6YqOZ3nSZulJNxwgHnBFCHXBaaiQYdR9Cd0/
/ykbjs594SD2+AYFhBgO5DYEE9+xW/i6vNcUYaF5xFktLSEAfebnZPQaVhV7BSv0
ctcdLsdxrKiuLigIMi5TzeT2bMkUYx9lpW3ZO3JkcbjC5i13UuGzNasgjZqIdrms
BEmwSfxENs0NgtijQITd3m9mWWquzmiqIW3jvBGkXlFPMN5wr8NhsKdbcQabJuuA
i0nnSw+oilmJXNFLpQpUC0KT9iLUXBzrv7xJf2P2oqTcxo8OITFw61q3nRNwN2X9
IjcmtO2MUMedafDRrzSMtSMEmX/4XpTbT7wtW7LVbARsr+SLrWV5Bs0uO1J9knt7
//UFE5ylVcoM+AV9E84jNnQaF6gXE/xoSMqMIukX/IVOIjH4dcAGzzjUqwURAoWT
`protect END_PROTECTED
