`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XAulHs8dKrW8VxhnZThdsekdnJmxnYrJsRHTTjeNoA8rFQL0lyrBDGiJqMM+Vz9B
KYfmUQJ3q++j/1JQvvnkNzhu9HH72kwLveKO/7Yxdg1v5lLhnNyEOvRJbwSERyLK
jIFp7iH7Iyjy6PoNT2/3td17jVhPlswntvdP7ggZjs0P8clj0J3m09cY5qoxjz+E
K43oYxzvaVMWpzHboOyD2hEIy2en/b1Sgx4iVpPF1gzkEmDtsDAGdnBME8T93laD
0fTY3UEbHprQ2ZDk2hLs55f5z6q+ffUYslrbfLYBolhutGl3TADKPuJpJ/zPYuJE
zhR4iDPp4l+V+kmmeVzwgt5k4HDADVMD9qm8p7xNzogJOercuaTJyapOa0ypexiT
8jvzoxcucsJxEhl4RtxM2CYgwpDMuNVHoisp9EZozrJ//O49Ow/MXTeQOPSDW15p
GUV4QElCMNq5k6foc1Bo9sQukPQbItPULG/zZ14cRgSFWOSuYIYhQa2TgAH8GgXH
O1auXczhfpXiYlaM5IQckGZLob24alpwwVp/55se7N6GbpHJHuzEW3FFOVfSLHNS
1Q85e5lLwj2FI4tcJ42SYQ==
`protect END_PROTECTED
