`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHr67BqHfhV/fyl7OFgaHEkjHvuX+5E7GyRTM8mWH9RkwJjzM4e4vdxCSqhyYjaT
xOvXhvV8EYDJYZP0WK/QGDq/jVcs/BX17jrsVMq42mP9JPfqxKIJCpGyRxr/Zyn7
iOMTK5dTCyzZlpx0FmKtLhROp70q5LdJMCKBn87M7XSljHYGkK5iziuJ84x/DZJW
hkx5Gdqmo+Qel3rUtqqsu04WjMKC6y1agrB5edrTNpNdAcyfLs6MpHmtpBpFBsu8
Ggh7Y2ZE5c1n9Af3Oilcw8aCHh4Lj9+JRW+ajf6dkbASs8brKKJoFKAfEev6xKdk
ff837Czwt7VDalYwmjEeqVjP3ykPAGte+YhPnDblYE9N+QMRmZ1xHHOyXSoIdurh
4Pgi/Od5F3+LPZBfRvkKhQRczZQSZyfpz0gqdl7Jyl9+rwKeiHfYYez2oeIvV1L9
NsMacZ3DJwI4DX5kLAReJAl0ezQfcxCwffb+bCwCHEo=
`protect END_PROTECTED
