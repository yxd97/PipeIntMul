`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i/RSyoVDjGm+SBL5QiZ5tq6pdwJCkhRrzGYDwB+ZwlPXUbFWNSyAKUtYfFjht6xd
na6lUwsbGLUnX/l09e0HsMc7C5OmTZxaS22/KmGufj+2k6Fh8bJQilpJ5FfUD3LU
8e9fba0onkrQwJI3CCrZW3rbrNZ4bMcNZladIMBdLc5cTO76IWUls2ncDLS44qRV
iYN7bLKwmAgWOJ0M48+V6C61dleOhHpohfWsR4upXYrAK7a0MKh1NdZOyaUGTP7D
4yMueZz1cVg6zWV6GEqLDDs9L3PM/N4SWwRpGMChH0BtLfHareK2NS/lu68Pc02T
QoAO+ES145rhGlN8GrN7NKBy/oqIyhHiu6YbggWpHA1dBH7nzBVJTJrO+Sl9rmB8
FUehqoyknzP/2hiwVxF+UQThhqypDh5iNEI7l+DdTWbuCqwJTbw1i/Vt/DiuaOxy
KUDiK03kwWQXux+xTit4zizBsoPl/CyHYf0EKLP/AQ4HYClfD5qTcIkLO0OYKT3A
2XNa2IhejYm0kHBJGFxghj3hN7uKQnTUfg62nuILeFmXA3BehRi0K0/zHVAXUuIS
nyp4lxGxYvKzMTR1xOAXYDWs/q5T56DPCeFpxTs+8s2bY9piKm1/1dgDTTOem/No
+Q5Rrz9M5sfgBc0XCXTsccusQ5ll0Qpank1NhGpFbKtng6YxecjtE/Sien8GXj2c
irvi/WQ4xLlt/GLkG9cCHEPU7waNfDjB+JO3sJiMxXEeyxZCYgzi3s/LVv8rwXFD
MsRIv04YHIzKU80z09Hl3TULMZiRUvruJOYot4yfnPNQGcoYukqV1ucGtcXGwr68
IjsdunoJ/+ln3Rm2zituyMm/qVsm3rzMtbUVTI1RAJiqzY4iRdLA6zoL4OmlekmL
QOszeg0GMCv7/5fKYb/rAOjLnNKWh5GsvlJ9w53TzCdyMh9xrZh/xmJLasCJbyEt
Pb2IK+aRy+2YkQPrXkFzavIRsy9QDfVtv3qID0HbDfRSffutv7drXzjlZuYUQkLc
VvHV6MvrOf+a/pjSJc05CAkfTHxe+YOt03uW7UKOlkAAG3Cv/t30D/Nhn52zqTfA
HVz/1x/zV9/tExlrVsWIjzvSmQfZxKIiT9C+QF8244YOQcQitEAAmyNQpfvpAQkG
aB+lhuflq3KN9tCkSILlMm/RF/Fzs3nJfN7oxtnj3ISD4h6vOceFVU/0TrVYfUhT
j0+ohxkzl7Q8diolI+WkEwJxC0xmuRLPvXllf7fz+SljF8OscMWz9afiDJTp6Fwf
IOtJz1fgq5aqWFGIBx6oJ/FiVrA2BAvTIt+O7al6OaT2AbCUPTbu3aBnTAWsBs34
W9jluIeGvaX3hrJfIcz5G8wBdDzmZRRkkJKrWIh2rRjUyFpsQ4eMfHV0l4QDc87Z
DCbnJDq/CiCbYRBWOjQag3putnrozLZykTDKhoJ++zTx2bmDx15bAarbH43FABmA
ZMPDY6SaLXgCgQoOO6fxpj8nFIhFcuB8MWzPo36hYEyyJroY574jMYwGqLGAGjjE
Py2zoQsETPh5UKOAphuNiLXuK8MY+6Jn6jV12gNNkUOeQUykOu9Mf+f6FmriHm9C
LgGrhhn2TZN/N1ni0diE+/BfjYCjC8EwzfcZZFLYKCiyI78EwG3dtn0Fj1aLrsVp
LnQzFZmF2IspQ/DUuMdrkUk1GRAyjH8S4CKKZSKTWN/lajUfkl6kXLrA6HoKNTYc
N80LQ1lnr/gdIQMj0DBRMJIKeAijU5cdwkODGavhsIps66PlKxx1LMWAOO5VYbyb
LCV6BERwf2dof03ysMX26plipRHBU+XKsYrTBaQ1/ww7HGpnEd+4kGvge4I5YR6r
4M2hxeblkr5Q9vK9roC27zz/4VYLIfRSsOTFn7dkKIEhVGRI0EhHunJtLfLYnnYx
J41y9Ygb2+kwSrMciQ6RB1jibPY2tHM4Fg2/BYQNOb4T5sTT98qfJxSVoGke1xBz
juK6jX4aDk3KxI3yT/kfgTpXNWrWv/WtHssE8iF0qVi7zVuoRJL/oZ+OORhx4Jnc
rSXDUT/84Bdx/xMVF5LMCHbgt41zHJ6qjwmm5VJAvSNFLFZX+t/0mLCo/7fVjzf0
DGVGaAmrwFMM0AERcMJ+eO8X/5u2ppK4titRra+qiSAMv8+csppozkIKCUEwaIu3
QYrQ2rfVdxTL/Gj+dNoiJjCu0DAYvvSHs2xrMLk4OBxoSABBP6SdoxS4qsbWZw7V
MqR9GZ0z6dXHQWAqFPQVsD4e6ygaDpWnF8PQmxbp/V3OMzZ82RiLRNgxZGSgRT28
ysblVnMFQqzzsdiCqcYgb7sWFPP2pgaOxRPEhHQgGuukORGCulIbWgnlU5BTAMMh
2b4XX6uZNv5rK+wOxHdGnrP9eJDvo0z1xY/J/ON207aDWuJbjWNPv72BU5yMe9fZ
tf3bujkXH/wfgiUHEwUzSzlBEOS4IdO/4Z8V6a6HJ1L7p8B3yj2EWzXbDv5rIegg
H7bNV00T/uY97bsQt4JmPABNvbI1e5eEFv1rKBo0BwXflqlPf20QGJgPnCKRJSdf
GoNQQo95Oen6WcQj6G1QA810qnYVIKiDyOZllCDSY5cruH9PcmGPkmOElKA1bdh7
oae3B0sjhX3uPJx8ZrWFOND3aOi2Fs9xWBJ7cRQ26SGhH/Iht4TXJLR1pJTYZOfl
yel7g68RH8/cyFPgINY8fOyxR2E3jZ6nNf7DYfYKSDU=
`protect END_PROTECTED
