`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K2ZNsqndniWssf/u1TzRhIdW+3MhTKWgwjE3/nUdbTWHsuGBMOUoEH6c8slLOX+3
p8kzJG9snKzH7qOgIpRBX30F/5qSx0p9pWpr5LOFvIoOXGse0bDUoFK4slG8wAXb
an+e2JCghJ+jQpUUHJjh79u2cQpVaA1lVRBuQ0+k8ghf0b3fJho9M0w1BTL3WxUT
XyWyEuEObcBWSjsJ80vIleXsT4wuXj0ADxVIvHbeF5bbsHjqyeKTlW/E+hMV06n7
1QCi1EyFKp2AFU0di4/we/+PtivB2RViYHFH5tUiJs5zr+ZjqfKPpXFzaOJCT4mN
4i9ZFAyC5/49wd+7w9kYNDS66+6u9opI4G6cmNQT985K4VU3iY2fOXiTzEvxpXlb
LArfqm3PbNlFHYXwlM39DsGlUbQZWSb/ydZPGQC0iT116+HODP7zh41vbJgayBOi
fyH5uSxnsn+bhZ3LjPphsEnSTzuKR3ZOLZdKwU/pYMYWmARQF+5y9qu64ox/AkEx
Xu/p8ATL8HtIsg+oiv4V86FrOi6u9FHQc/cHREbJ2i8Sn3y40nN6zGzoY5rCpJaa
tNV4cHd52YNj3/YFyul3bjVbxy3kTnYVI0gfYkwXwyUHSrXGnNRRfuYxpBAPmlnj
uIp02DTK8wm+aF3VrziZIyu/hlOiE9E3mdOpYGYWvNzBn0gE3iuxAWUd6qTQvMgu
IkHyb621/GHg+d3i3WtJ1Gg/+M+SFKez6GCMO2Ot+Zg=
`protect END_PROTECTED
