`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8GKHoIfRfQCWQQE6yHlhc2CLSZ2gkz3GvcbyH7fhA1TnE8YTK8te+RA4V8kETl9
a/um/Zl8f4BcHmd7wlYSzEtEeQmh7Oh/wdkIKs6cn1lSFTh9pld7uymJBBNTPgaG
ytP1yPtKOy7q/NeZ9dacetxXbTnbn1wH1BhsLHCkGVcPTCrjI5/41Hc18T7kuNil
Mg3J3xzOp51eG86pCmJiHLteOl7O1CqFIAwsFHmLs2fov9IUu44xBHeUcHSpPsrX
r1MQgTRA75CYKu5eNesvp1yoBkMW3fgXNYRst6ggE6RuR2QAJPuVfYsQOC6HhOei
7OH080gGhbhnxs9SB4tbMw==
`protect END_PROTECTED
