`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UynOsvsHNgWFwWT99jsgStUTQ76I7f2iV3aO/yyapXQSN/NowXjC/BtR8XcW0AvD
JOq6nlb6se9tMbJYZqljUxptX0fICyz9tDm2ZkKUDI3Q8P9OdZHawFVAzoPzFjBG
3Iou6GOcKedhpkXkG26IrbsJiu9HWiLcywc9Lxjy7jL6nLkSNj2ki7HeERjEHxnt
go43cR410bmbgf62hWmNJawX9iM30qcHXJXgPPO6F0fSzUssYttOMmeAjbmKga4f
n8iP575VTZ5MuOmcDnKFleSFBCTBXSzhhjigefaSfRboYrV22fdpkRpITWcj9AB/
iYwlnbzdVp5+p4S6QVjzxzar0Y6h+PqpexxenC97YBto5gOFABLUA4laK8lX0j+l
08NVa7mzr6oEJ2axLfzzX69S/70dTjB2CyV3AYoo0wfONXfVnpIvot44bw2wFHS+
BnEgUCb/Wlki61GcVqDZeawfx78IllyRXdvZt0FVAR5EthyNPMuSYD5HfjfBjil2
9KBSsc5fIN81wxBUHHhZzqQ3O6tOAS1Tb9PTOvDU601l3zkXFJopCgT9fcYt6pBr
mmUnhjBE/yVma9C7OJ/i+2rUaSBn0hfLAIY6O5dYDiMGRlIa9CFDe87l8GnLQ2gN
KJpnXw/UV66O3NSJ1bVd7eAOSkwp/PBDiQvRD8tUBkVmwwJZBnbD19hm6nkkHnxR
nZO+Y48YeDLe52dBbdjcQVxEiHoQ59J4o2HByjDUI4aDOpWkeO5jbwvRBT3FlD4z
+NciubT12m8EOgMhHQQPWViebEh10UHf7dxcaOrSyTQ=
`protect END_PROTECTED
