`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UT+1R0cGIcGAMPotc8F5glps2OBfE0oqgZiZv2/NKeiF94uWlQDuyj0Kyc/JPzT1
fjSmFCnMe8arp8OnrKLazlkGZUdkllpe87KJdE9Zi8p7x6oHoHfz5m/G24rePdWP
v2uLciGTo5UVGTs1gWFzUL+gkV65MAvBkfJRG1qAVQ5fZGsSiW9BM6RC3bp1+vKB
4vmF1nQ+FlDFUGFH4INbvG9xjyPGP0SLOtcEPouMjieJD7FyxoNemmUcks+VtBeb
Q8PNnXGO1QUFiBbifkw0IcTvIS0bMv3DFfilKasA9r664GJw+KGMkW45WSNDSr+o
WqGVsHYeVMm0sJPw8/oH1QK79h7dMA3vDfiW9zqQIS5KLwGY9cNR3Hl6+guDIso/
w9+nfxjkrVKeYNBMoymDpQ==
`protect END_PROTECTED
