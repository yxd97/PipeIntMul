`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCaboKlvWTDjuGaWWPvTgkGZtJl0jciVNvGgnPxWww2S7kvyKaaFAEXov4qSkKwi
Whqcd9XzG0rAn9el8VIjr5moRXbtSzjiHcEDHKi++My2IeZRCRCS4O+B4IsM/Fpu
YfORSNvFsM5zlwzrZyuWd6SO77W+gXmsdjlZh9/9BQ4t9G2LHWd37Dgvov2agVTA
Tql5m2Jme5FJjBEG3JjEYwTztY5Bj0aiSYGsA+MVmTeCQEICCgPOFSMAWoppRNHE
FSqtc6dtp6Ue3veN65UPgw==
`protect END_PROTECTED
