`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKqpfdloQgFfAg8bQqjg/TjqS3cEU/BikqvePrlIBZp/CPSXwr7XyAHHVZXcmRft
pMMDYUm3MU3TYzskmf6/r7PkzT/Vef5O8uHsCCfocttw+kJ9OBMg67yd1nmgzuum
BBjBIcKFufNX0zuXJIFbMTuu7aASWTIehq8eZ+ZUXn2J3DbrqaAuOuj16aHJ2Vsi
FRN2R9oVPlyNe01ysi/U5ZFj5X6Sy1uDiZWoIuc8jBYOHxi2Eo0TImxgzfeTd26f
38M/qqPVdZrCEBL61+g7W665Q+86IJNMb1cP9QPOT9fNkT18PiOdePhfyI+w7dP5
OkUBzYf7Yi1kM1BhOXOZ/ew8KQkzT1/cHhJdH0Ii4xCyjz5buTPz9nhbXeBnrQmN
jHL3mtErSjmI2+ePxWOvWAscZWDb0FJW3+fQYViEwhR7cCcpfMCFX7vSS3Xvogdo
1mIXT7oJQgnlTJSPKaROWJwz1n9yjRSaAOipzd71SEkHTgCnjJEChPaFdqkrK6PB
r8uQH9jH06wK07BE7eMilYy1yGYqFYroTXoLUNpaHod+kSBLXZhtkH+Twvyas+XU
FZHEBRyOxi9tYMjKvr6x8A==
`protect END_PROTECTED
