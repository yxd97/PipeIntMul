`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0aFFp7+GnD6q7IBr3RrBaeGVGCJmmH8JUmUQV6e1bWilD3do7CIqyjRXZNtROmqD
K0898WvRmqjtzbGIAgaDehrMDQPOuyd3NQ5BfjbZlW2VVQ/y9aDw87FUoeoeCk53
LYBg+bGpWJeYyLUBteBtfhuxbTQkkcltkPsoqAa3RB3pGBue2AGLuSONsbMSmwC0
3EObJwIgLYJOanVHbmVIcpuZKrk1owesw1qU5MJjt/qhtDl9rnPVUdN+gyOSiIkZ
rvF+WX7/a4mkZqHYmhw0ePvK54LchgcOL1bwlOP5uzeKJNgR7EE8KyNwt2jR4oK5
JkeYoXajPaNiNMs8XQP5DtgZDFzuXDhNYc1java5HMg/k7woOALWl7r4ASMKI3eo
TdAtseEiS/u1fy0FKHRfsD/EsCZFHwxsFEg6Pfra46ddIkqF2ubfozttCIj7PvOR
v2DgPb1tIr6d7aL4ELzQkHyOwJ+4J/ai1Xrz58wguHNJ0xcLNYOmMAIuCbyvAPxh
UYkEC6O1y4sL43az6lWYv917ClzVVQ+Wm8BnDtEwS5shIgee6rTOZjGSdCN3lKwb
+W4HtJ3ASe6QnmZihJIV+jEyMEA5oX8/WC5YRZNr5YDTZgpOaMRofv0H1AXyfFhp
XRvOu1aKgpQ3Wn32YDx5QCB3PhDyqiWt2V7fTRTLfjZueG3iZAqf/uwz7PAnM6VG
T8Ib0KvtGZYep0VbOev1cRHUonOkXWpdI7SmdtOxs9uCYG1QbJy8DTsG8PlDf2eh
iMKJ/Vk4F4G4p5mGEe0xx8sBLuEYMtcPpvTeNEgk5dNWkDlw7h7frsQ/u50JjEkz
+CdI+zs9aTEP8V9WNxkop2Puw+uF4mjdm4QIZAQOA6ZdBEvymPiS0xObzXsi5n49
JRRFvQnbWaF4/t5aCS5s/FbGTfFPlJfyxlBkLsWLYt9Gc9+L85BZplxedX9Zo9BB
`protect END_PROTECTED
