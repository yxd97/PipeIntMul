`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Tf8MvMXNk7t2XIhqXfKn/MR6b5TrfZPQvLmBM+4sqIClzUbKdJPdCMXUGhBsheq
g/UNQGsVwotzf+Akc+okQOXZfrqKfuuqjdRnja+DIaWbej2pblBfmKdGvhaDCut3
dVV4gtKRaoHduZ/ebavVdbuu/PIFWywDK6m6hA4FxbWneu1O/7GxR1vLk4wTko2x
8CDFGxBsYzG0e1WVf9EZxgUj9ZcV0Ejc437sgnZSmNhr5jyOHKKDdK5Reu4lAMKj
M+2mtgpfLcpQK4watXj41Jm6vo2QkH+frZMYzCHMeiFB/aqyR/UwFyQSU5HczLpi
seyQ4SVJdzGqHjByycLabkwHk3X4RvboDNukLbXHdF1EycKyEj+R9RFWAju0GfOh
QqkkPg0Y3egayXRm8QB/FrojPiFgiGQ40CqAupi68XOQXJqYNxDGzayx3GWO2eSz
yF5kS7t+lEPTi+B+WhU9angJtoXtdQqCzUBV0xzq8Bd+rUVkqoUx0c4oqmjqzUxN
kTJ7n/zHwLRHkToIrqoE+fHjBD838in/hjqSaQcswqABTbiDBpbFtUNDpXoCoXDQ
v/RjeT9pbuoQTsATlRZCYw==
`protect END_PROTECTED
