`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yolT+2sd3TUZVGcQBY0FvzUK4PDAxnWRWHpGiCCgyZQBa/8TdQcBWXqltTaAjRTJ
aOvPOuDeonO3a8wGQUv+C2NfUlb4xUU6H8y1y71sWmBDuaLUf048fXq3sfVEGA+g
fU392QybJ9JORmW+2HOTnPQ42KDoaZHNfY1NFVH/amoGLHtH/a2oy82tfV027RD9
xOEc8jJvOSulN+YxYvo8FeUrgwUlTk3/3QPhILbXOpOSc+Udzb++B0uGimvNtHZO
cXD6odMvkAu1qCXbuG3Hwg==
`protect END_PROTECTED
