`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r+iB77Z66LGcTKdmPPnzkJAAZJPtXMZzipgC1D1fI8pYeIWCAqwhGsqgdCZ06KQj
X1QNNWontx6NPmwvVYUYD7KUNj2vFw8FqNP2hfQMKxle+HmX1W6betCUQodarr8Y
8zV0heXmIko0U2uwB/9YT65DfzjBAB1cfzgiHvipsAJCddkxs2BGHstz3dgFc+km
AfROO9n0Pxtz581Gsas5U49vO5lnJDlnLcA8A4j0RnzVvf0phQs/XspEwu1xnCoZ
kj24cgrrTcm8plQ+JcYcqyoWOXa3gYIy7fa/820t5YeeTbTE6L02s7Mc76V6N3SR
H2/7Jf6B7oU6j02lt0AQ/N8wldvYJd4T5lQUADVwArbpId1ItRiYKMJP6bsmeJc0
K4l74+cazsRAVfIguZGX3K8KtSK4HdcX2AMwxyoe/kkQa2bz1UI8bByCZLRCgAgo
ZchQik9WVOHXbfCKhMsInFHVAmkDCLjdlOY50MOEFYJDPkVk4W8Ld8aeEh0JlBAh
`protect END_PROTECTED
