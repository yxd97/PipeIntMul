`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zsB51Yej/fLnrfGjQTrlw4Hpo/nYSkNNtExwswSB9abzDmVCaWpvlnz6SVxqvzWJ
eDYEobEElOmDDG7sM0KSfoPydVzkJZTDwYGTUpWeZzDNPyj5W+VI+SwOFrG77vkC
BiCV1Lm9VP255H78RJekPl05AGO2HhpbkvPFvsW4qCzDpjqpAzlCsNdeszh2+nBX
yFq5XQVdF49/Yq/Th+lbJBu7iE9bF81qPkJ8DaVWXv3SuLML+I+8g0eac339HQn6
w3DW5sP0JVXEjZMsaYqCb6baf3C7Gy+U91CTy9e4l2pQMi+BHZbPkemTJlMdsPbK
fBAlRMXlEawlFXTBUS2guAFul7isMWJ37dEZnJQM/D3kgHT8QmVH87JwqkjvVCre
vTX+0i73V2SKlJ53YhJZB/6VaOAgJKjJ4of+1ebYDBAhfMVi3V7kUxOmAeB3OgCJ
ErFj8VCM3iITy7KkRSrPPMK0tp/Wt+t6MPmhN7fk8jPjZDLsfo73LUN9VML7wJRD
wY/rf+tvn7I6WoeCkDZEFD+MohG+t0vfv5iwhnrElKs7Vcf8gj7FI06tg4YbGxVp
/7cE5NMJGE6f3lFSW5eI2Iaj3FPzv6xcOJe9LO1x4LudBDtB/Vaks2D8oijDPHud
Qj/dxGRwGLdxFX3R1rrA7g==
`protect END_PROTECTED
