`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFXzReg1d25NEdr9u/Pz+WRX9EVZVAvYkAFMyEVvlyUVG6j+6ea9JHI6byPezl/0
XaUEoEEeaWRqKJtWhxjsa3QjkKAfO/nH2X7qNufoS3YwhZncULkZbsxgDgu2lfsP
DQ6/LlGBpWpDGsTOm7hjHkuRQVF5yjcSTemptdhXQtaXzdkh8R31/qFUQfjbNfg4
QBxWLMY4gP8rK5ctuUUMtdoLg/iTdJq8/Lv0y34i7Vqp+ylZNr8mNAac63KB77t5
uKJB8tz87gh1ObksMf3KYeduPIFXYX5EnJuO/XeCon7udnmukRYVe6JX8Hxg/qY9
tN8bqi6N64OYizGuqWAByo8AXnjnRYyfWPjiQ8v+td+7hUpLXrb/p4qdkv1ukCUW
VrNZB43JyLZr2fx0z/cVmbrFrMMk5E+zXqJD6NXHifTlYqmrRo78ErqGH9OHUwhl
+qvRifFpj/D2aKqKC+IccdHrWfh1D1AVOP8sikUaedhQtHlgjuh2rDddFOqfRr9U
PBfkZ/qysdwQQa2Q2lD7cIkWhAiWBjMTT2Ngb31O/nRJDEVjhBo4i5X+Pl0urMQI
zmkVtwduxk9eEizkOeVN2/s2UzfiFOwdBGB9AI6FACpkdqJkOIhU54xz4pegMtT/
bfiVaOQJ4eSlIucxQWRA2wrq3ljVVHRB6GWCOuIWmzw8e7BVayGj3L04m6Tc1fnO
5xInGKENg/HTQ/cHC2WofQreXOTMMoeE9pjTRFAH3BQIvcJfQH7rIp4iXqNsNyEf
zFuRYFDiIKseAqbgrYfc1m/FIhNNBmSKOg7k4UQyFXBanVELcmigVWKGYhF0G+Dk
WgvOowrkqaAITN5OBTFno06I1Aj2nnhMI+8jCFkrB5FMnAr18Qm3C2vSokogYvSS
olavcahQyvZF5xrJhXWvgQMK5Ct3/6lknlb5ijNM3YHW5vMUKvde1NwtU33IB5D8
j5CdROzpVAe3/B336vm5ah4/3RK8s233zb+vnqE9UMvjPAvRD/Qj6+YTlK7Bepog
AnG+Qya0YH7f/+XyaefILh/YkfZpi4JfhhnIbp4IjoULOCHvMLUopaZnuL6Na2/I
VofqbjNkGAyLmw/yLhKKfhH9F4+Pc+FInTn725Kjo9swB1oTgBiH6alC8jgCCJrt
rnr4SNI2yBd1YLtVpoefXZR5Mvw3c7wm9ERWa3zI4qtui1sT70YH8wHXacmzaWy9
jRz4e504FT+htSG7fFSpiPMcOzNiM8CdtZ6XUjT3WFOAZxkXipjcS0j85Q8LKvRv
IUGIdKrF2SnrqBM1nIox0a07x0sVwHbJaNgouQs0p9Zu0+XfDLHrGKVfmjNj703F
zYIReOMHg5CPN+skwPY3T5FbPCcVlN0civdFzovNST/H7c288kkVuXIk4c+6STqb
GSq2xRB0uIKrBup8QAbPGXOxT/HwdWvIAJmZ2v8Xpqc+3eqdHRElVwtY1ESEkuU9
4qWAl/XPQWv+nCW5WgDHYTZpEQShoXxTQrv2893XhXyEGo0ZBtWCrGqkC7kpEsKS
fpW4ZFkAwn/C0GXfV5V+grhqWTFRCEfOaBXB4MD6xZAnGvR2dWtIm2PnoAbP89dK
TOCR2e3d+EM911vf2wCugOk2Ls9JBqBg45XLnrk5iaaQZ1AOB708b0BpE/BP0sQy
IIIeAaQp9iUneQRZmKUgxMkxXN0C5gHPu3l8wLmYzPYJ05r7iCz3MfypHcQhwasf
czjqtKHNsj0Hjw2Du4zfSxuOBHffLWqxRr/f9AAHuHZtJuseVrbXohadfH5mVmmK
6hSmcEfQ9nIKBA157Gtltr0rD24dlZp5fOpKgWqOPPOmMOWIXHeok62nQb0WRXAo
G3tucfTZ9hLOnv7L/fz6MAFrS/y25Qh6FdUtwHWeNotOpionp5oj7a0wnaCLmZPc
3IYYpNRj4IvbihQgswIl5vxRtUHGXU/QB2PvJNHUmfMO1v7SOnQhlPgfmhPZgu2L
V1IL8ha0iX6Vt5PuVc4BjhNBAHWPbilzjv0NiUi8MOPjF6AbjBkbd4HwneeS5i9k
XZmEULYPn3Q4nVthAh+X5hmRk5op/4L8M6nYjEfug0rZaIXdF2KkI4zTKwTioLaA
q94j+CiG2e63GjMCwyK+suXHbRm4xmgLsduJ1PeG9zVz9ZcJYAdErOy8TMv2MZ1v
VdknINb1P+tXap95ORm5hmefvUeHORYG0C0/bD1NAUYaB8NaLtsDWEAbAGv3vwRd
d3EcmHREQhiQsHysneGYD9KY7AwLuvRMOitwvR0VwQDRt1XRVfGNJeP1hqzqshdQ
jFmBiYAw3/jO+Q00xFafcRj23WUT2KHKHNzHhuzOR7TWes2qSbUBoOzBvspLZWHs
CZCzQIZRSftC7pcG/qFU77t6lzFf6r50yQeL0cXSn0UNRaP+R04TWib/Sz1p8SgH
E4TsWUre5SiCtxMwbRRXawqnQ1F5W5kELqZ4pfUMqKUnfezxAcsGtWfdKs9EwwMU
5gpi4fGS8F1oBt7yyqhrmUv5DrtIM3lA3lW/+oCgrHcgWv2AM+C5kQ868mG7tPbZ
05EAovAuK+NW5UXqFmK9C7upDAGF4Z+guel0LVGjvyHft6E+pMW7H2HXKYvej8hn
UWO3HfZdY+U47Y0uXvJ4aWA7Nlne16HQkuW0bzNQjXkTeLPKVCT5As4U+1YlzAWG
eIoAagSNlA8VAx/1P7Lb2NpeuaSbgCnJdbSIKJFXZy6OR7kguIG8nXbX8BRiZA9Z
4rr0cOt8UQq+GXydgm72qRJV8KXpyMJi1itdFZ9PvdUA7K6mYyrTLHqq6OCHfBuU
b4Crn11bdd3S2vfssKeKvxol3EStk3XFxOLLvZSEDBLSeeVXLSa6+wLMM70b7fjA
+PMes0OqeecHLnZguj8xEH+kOrEprs6/ONefUUHnimaQc9uAHaX/WlVYqrKq83T2
cW4vqgcmRVTTsVYd7zNndCg0iGMlC3ululx8vh/TvQ8Wf0SbcdklKWPnbzC7BiWv
MaVKAFf7tfpPpeBxg5id1fNzn20iDgPOsBfkbavGC8Sn2OYWaF3DBleRHjn5I4bW
mETpSHS6QAhkhSj2GoCjGUx/SJv0N28sBmKvxPKEKiQtbGb/gtFCD337tyGD2WFt
rv7lc93wNoOLidBqhVSmgP5muRYijjWWVv5rkFjg0EZA3J4iOL8B4ZSeqIZqA2oB
Ni6eTqMFkshIE8ndmMCJLn0b1q0Dotm7u5hUf5mf+Cxbu7mS6hgylwjPaahc7cNy
LoSdQsnNXwe5z/y1N4CTIAL7QeFbK0q43FXiy1Dg16fIlVvg6LxwHPeYz59Uae7A
eIKg9s0QrJVkp1TcrKbp0jBaW+Ygy3ZwQiL39hYwpUyzneAu6pI/Y1MPmWPY+xDc
KTIDUNgxLt07otI45vYUSUBTIg0tM32qrHXqo30UhhomSrB6DPKbWrPZh7VemuzW
cxAG/w1H4P3/NGau5q6IKWVdkMhZYl4tvuQ3VFZ0DTWNsZ4fivlBhx+GZCXwy0cE
I4CWirBtGNEVuZmHWK2iVjS1ZUEiLCJPgP0E++zhhURnfTt00RqGeAqDyG76K2bq
bV6J+kPul0VypfZx4uzOxuwHDZtxzz+peOtL2k6RAmLtdW2TvAqGcvZ+vPq9Bd/f
o9fksHNnQQ1qIQnIhxjdSqIQn2zStzWM0tbi+i+Y0lhEa6RgfOB9ZxhOQYb3DsVS
OxeCCt4YNyblOSSFehwz0tCd0oFM0R/8VYwaF7J+vTc7pjcETe5pqfRovkErwxia
wa7tDyy+xlh8+88sWzuPYYHRivRmP8aoQ6BZGxO/y7eXx+9Fyo5EXfBOIoF4lqV2
yacdL55VevK2Yn5p+AEfGoRwb0dWNuahwhbhh5N/p4Rny70AYNcwZMCYM51AnR9E
EviaJq+VBg2yq+emMsU0xQFhdeJLu4jK6FzzWNCsItg6+zYpB5e7jWmI0eLQo98E
U/ens702EbN+51EpEGnBAYzXjRE9Xb3H4N17Bff04bJuu0ZNpDdHTmmHIDfsB8BS
wwKIOIA+4yDRzpCVcjrXRtx8MJWOgnrhcH5o/9gicebSxxAUsZu/1kzS3tC0M6Hx
lXSbJbkNjVZsooSPCqB8YSkORt+8EJ+2dgvCY014dpgVjVfU9C0rZIacFi0qo4y8
+tIQYnlgyqrMVpSj5ngByYJpkRSGNVWpdTnkAgk2+Dc5Xc0LIfi245OtRUVGUMY8
ZOfDzDjc2ChSSt51kiW3H1pE1neB/dKJmvmLvIVTcR1qx6KzM2/RAUEl27X6SF2M
VgT39SkgIb8qYdXN+MkTtTj60VNVf5QS8nDrJwmWp+Ntq5WNNjGfuYuxOfdgSgEM
JA2PwJ2cZxxQ6OTnG3hS3rjO1fDFv6nZO9Un1Yy8A0nIH6ksyr2N/TEQJdm2uqMg
CwepGCAzFkpMZrC83kyvuPdE0ppS7HbTRe2w5MFOFroR6RO0pLS/Ok+1wpnxk8c0
FT9+pJA2VfL0DhTw9Al6inFZ+7IQ1rfpXbIjf2/T6SfeHYYw8yCQgn5S7KNBWoFV
KgTS+WpHcpdt5ZzNl8ANkv7Gog3jWlecrJn+mtrV44yprz9+R//i53q/zuYvLSW0
qdH9wqoZ1KHpGDV7LjfPpRqhNI72DJqAq+V+XSGPcgV3U+w+i5S1uifhdpD4yIP6
0OIlcGxyqojwAS1xyIbk5KhdMh/6RCG5kc+98Zxj/geUmPWlVXY7PO3nuGjv6aVD
1ljbacphAZbIyaw0037WeVXEIBLl33TYbSI0GDBN0Bo4EnOa2QG01ErQ6mIVqV4+
mdGMrVRKy56spIRDSTheI/EbVNkO8QAokPCuRAEjkYCjfnwem3yBzwFPihb2bmEM
I16t8gYKVKZFDNGkP0zGjSOulKH+ZVrdYJHRBGABLLwJk8uQZdVXgJnVrZ6JOBJK
x4tEk0AanuZZU+1DEHGQyGm42NChXha5ueHmhk5ZkJYf4J2ZOCIcmx8OWWCUhVx0
71CErKOHNDawo4ESvzD+/z/ct/D/zUMP3QiIjc/drrpr5I0rSGHFb6FspiAiacxN
4VDWqAILhobFEo0OA9TX48eaCYhUIpPm98loeejSJ+Thqj0VFQsYR8ZvIOl8OKwz
WSMtJN8Fg4LuBooqRga2uElPrdxEWtXPVUOkTeFxcJYnp6VTjFAXuGBUxgxbxL6f
yjc5Dj/vG1RjUI40WdJYZzuQ1XxWN7apYVLXKBz6EG5YQ6ip6JB/0cvqsX0sYjUz
1vyxyt4FUlz3ngaEh0/mIRaoGXA2E9cF/RJOnAKJrgH6q+3Ckn26TEIKpDZS7wJm
ldecSQt9APjqQtHCVNAvtc5m6HhpUc/G4/2RpY86kd/8MUFLQxeoq6Ww4s87XUjC
iVoNd5RvATbblHYW6nwXpNVCHtqNgMenQLMjusljEEb+8b3j+fNM4B9ntfOw5JCL
LXP8dz454UzMyMEjUJPHcRuvrk3ymstU17x8zyq7IsFZAGhoeNhZXob2RM25oG+0
w7mGqoh7BNFptMFf2dhaJDePLs6KK/KE1qHo3TsePmJytYAnHqqRq+HCkPXiMxqR
405UX6WDYwRYznPhaJXcMVHMjAWcoFU+ODslJHM8WukseJiEbAxWtyFYOKrQQ9SJ
sgPvLZdL1kVJGAk9MDxODW8Sca5GsZpOuMb7RW/Mfw1XATo4Rpg102JzDizTcx6O
deTPJcSAnVfbZIku38o75vAAcUNsLOIKIfyqFyjI6AcJ393eCbJDZOv/nL3JcHf5
B8G3sdNGpKQFcj1BL49n/6CDWsIMqsu4SiLPaUjpQvmP8trXpKIqtr+3HwWXdEkp
AtGWcbYbfiU/O1zg/WCZu8vzYC/qdfNrCNV5KBC3F/ASFc8Lv/6QvMmrgC6SdA9O
M9H1cpgmVTUxu2xqTHds7aYNSJ78IvGUW2PvCiNviwXyKxvCyldwM2PLU7uaAXEk
LmyVlX49zLmC+SU0o/L4ZjPWka1ShBuoISN6hX+rLcDjV/zQ8dilVVUxjLmDny7n
XSqErvpC1C21YFDwI5ya1cZ98SD8dXx1pUUEZ4nZavRxGWpN0tHEanGH2rQKMq8d
IJ7GFnSqBbN0N6t41QheJaFZ3WXNF/aH8JiZSC4eD0TkAQ7kk+JnpPZPiY/RealX
m4CRPYUrWr3+3HSzhCNBrxsActdGUeHM+j9pwg/g3Mgca99NvtLQPBZkttGrqhhz
aipLLOqbWWswQl1mhyDe/8LOAUT3LGyE6eDqysbYHmLGFdbOVby2g204I6wXnuYQ
yvGL/z0goWyuyauhl4ruEmu+9Ul4DWKwskuOD1Imwnghmp0HJj5MuNUoiu5+oDYo
dnitR0c2lEynx1YeN/7RcKIfedP7jXnzE+f6A2LrkQNBlD3JEkuh7Eo9RQXm49DG
nR4IiG2GZUmzOPQ814pu4M9mPBAtuatA0Koig7sc6i6tstXwVBCvPsr4m1ZMSlmj
vJa6KjeRU09m/RieGXJVj+okcV2H34ulvK6sCGiBNulIDGRAivrKKiC75r2nItei
L23qrKyckTAC0r0bv6GxmF5eVVziwk6gYikmTrq9n8V5UqevKQRPc5HobiyfUnEZ
3QVqYDLA07M8ho2FR9raX3KB3P4OLPKKNa2ZI+rEZaV6hFp/l9TEvxFcSat+SFd4
+seL0SOgReqHckSUQawvVMTC/hX77G676VezKNgELIuY3a3gc5F0v1wPI+kOcuOL
sPSAt6my3NEdGZTqKqCPR0xdc3s1AhIPJxQaU5mEGN0TazrPfIqP5O46duMt7k+/
4ebrHhP+iRTcBBa8RWS5C0yXQJTARk5ehC/mjyIOksB5ZUrQoUrHqNvM00sarL1Y
qhsK54Hoi8nixulGrG80BK7owEx0DXBrrBEeJtrHvNAYSKm53cvK6z+sAJxlvmYh
VlPL7tGXT29sFxB5NE7W30lWdSCSpnKyfunKFDrtt/ANDe81bUUkBIJpEyMR9YdN
pvniJO3CBnsTkU4ooCN687nzaXpo7iotdOUfJBZGDiIkaL+I1D7hLBI0MAXFH7zI
akZGlFVmvChTp/lr33F7sIP7n9FYG6iq69EXPBLbieMdoziPvlYLBbjzNDDhMoHZ
n/Y+CzLAChuV0zuYTTWCj6nfwXX1VaVDBLVyUeGyC/zN8wkC7JgZuacnGrFTDTcO
ET69Dfu9EN5nZWTsXPQ7w+GOrsBRFTPHZKIAeqFTNzTJBS5ZHM4quNL7FVXRT8pb
YQHucsUSgIsrXWV9TqOhVkKbRECmAuQDyaxta8h+o6HQAnlcNE5rP5Ay9BX3wn0Q
rPc7wtpKY2TxAAPAh++MkwcHAMx8dfDocwqF/t8s2rd7HQL62a2tizgFOk038cwK
R7IAA+4xt2zpejQ29AUI6tW3bl3fWhORA0fElSHNWKoI4T5qkZVARmRQcQtUhE+F
6UnJhQ0Gox5h/Q5WuQPhd449mqn7ZfQJrxu4qQboWWxupRrjOYtUXwwkPuSIzP2m
thi4KFJTQM5GEjJNLjIFl5mnf6CNZF3z07tUjv0AkXCZ1EM9ZkYomTRCxqpHysJH
BoRCroHdAUgX9hJkp2NMGyg/Mwe043Z2lEOZno7fFkiqrp4GwJj5UVWnGq2wEhOI
oq6QjUcX70/ioYMyP0e2FOUd07GWzi7Sbr2fYqjcI00To8kAY2xuKO/ZMGMeuxNk
qKYXPq77x3yCUXLjQmwANLSZd2bZU4Td3ScRhGw50PpWagAskZuKjaN3D5HBj9At
3fQXXuCq/uRvm+oI5AysDmX6lTuWlD5EdrbY9M6avWniWGy2zPCpIzuJE7WqeFEy
P9jDlD51kdVRC6URIqdRA7B4ckoEtwJ9qP0B3yC5YTZwrlLJoPvGkghcYSuOwTvD
9dmi/FxdNpEbvKSxWddT8+n4XrOr53aYu2g2S4RcvdsoZrvb45xEKV8h6rTHlru1
7Uz17W/0u14FNEfTwUbEW8mksqU+BDKEfHwIwdap2ndUaBB514gzEyejOpkEO7zx
435EVYDWIb0FmJdq4JwJjbYmwcar56xnxo60dEl5RChtW3sdmgr/c5mUVHdAADyI
ICP/6q8wnV6DT36eIa11rP1fyLe/KUiNEOqkvj+WkbSEGYo0BQztfhOTTTO0cWM4
+HOux+Ewc8p5H89cE6Fr502vZiEtBzf4WpXHkH8IMNJkRhM1mvT4+NxbbbOt7MXR
`protect END_PROTECTED
