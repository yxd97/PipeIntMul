`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3cbNWyUU/4B3D9ZqDBpV2OTfhU+PEBYoXsEOOGPZ+zYDSjs9AJ9+ilE0dN2/NdO
2eaTChQ4Dd0Jw4+oCEULVcNcmyu1urNAiOXf775YEyUCptiCI+HpyZpckEVT68ju
5FFMe+FH7kDFtNh46FnT1N18VwZBWmIvhWlfdWPD2zpHbR2CQqJ+bj+5JhDSGC8i
zAeAYliwYvZCp+eWYPYq04yvwjtyy6kzA5JS4qrSUQlJZhJXGqMpqmRfs66GCQRu
knnHcRCns9mrBIWG7OKfzwT3g7slfsTw8m9V4xixCbfTmyg3Q9zPQLgoypYd5idU
`protect END_PROTECTED
