`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZAW4s46KHmQgOXIHpQ8xjoKaxdxRfVSTF3cNFx2ee0anB5qI8EWTwdD6ckuE57Y
/CN0eFfWYeI9FWLf4yN3DzKahnysYh4jScZHqv/Kjh0LtTh66c+HdJkLDSKrIe7S
zvk80IgEgb1QXYx6YMQZG8yJ98xhtWgCSpG9kYvOe8xFLRZ4+uyYpQCXCUKh0Chq
9dTle+yXdN+uLi5ehZ6O2JUk/ot0B0LOZzb+URdoXCVoVGrxudUce/uMspjl3Cy+
Bz/pTeKU7OXywOw19Fye7uGLPhq0c4EIpQ5kIWEEQrs7gPxpai1tTy13fbaGH3SX
ac1E6ml9kskenuBE4DS0nmcRwrP0UsivJS6HCl74lnk=
`protect END_PROTECTED
