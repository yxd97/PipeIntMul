`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hyJHnMVEbcrFIuStMWZnHJgvN2QXJOX+6I9HUPhLDHad+3we9FdPzqxNG1g9c2/V
UDbJbttreD6pX/6b/DCZySlzswrjD8XUeYOkXdIEnL0fkp/QIeKAxgTRdNntaGOO
nnCndV4dfPH8/l1VvoQbR17gagPcRxO4AZG1u+VDeyS/vnsvgvrkUVHMSrinl4sO
FzMcf4obad2txdn+dTAfpWL1KIYXYNUtQnH505ixA3AlAWbg/Pd+8g2hrBSCR1qh
ZUqqddYTA6lNYkl7hLXW8pO+0BKeYjwTYl8Khf7gpY4YyjgvVw9ei2VzMgI8ssLI
WxtbFfgWFP6rlI0ThTvK3Adog0uiCk4fq3YU/buOgU4aNN1FUbhmGr6rDFoRsqCG
Q58i5HHis9WkZ2VPx9X/A3TPJb8evmBJY/gqFeak1UXUVL7tWTVD1AF2Nk/MegSK
uE8iE6y9yhQsiyI/jhUqKb1P15JhFpW47sP1IqYmd2oX37eXnSSlUDJYC13uiXlC
vEeecf57ZdcP2wq8/cN+IVm0U9/IGersc/RZ16j/EMbZ8Zx2qNSEYa8595LUCyEo
3z43bGB8EOrwRoK8UYAXtblMc7zqLJcatVFyE/ViI1Qja/6STkvfM5czdw7YAc0T
tC7CyT46QRVJTWtuyx7nrUC+1kfLMnj8QfNYpEPzR1Yva9FYl0mHZJ5BJEvzbC1H
+bHXe/FSINr8mAqijAVoSxEdFijAEQUI9bjaqctbozEugjzaUFZES3hpnuPYGdXj
4+9QQapFDxjYj3cWcQ93J0L1GqfU7HJ6epztOYwnWB3iMrIYqLVvdKDDEMnOwflt
u+y+aka3989gc8PQkW2xLc6Fa0tK8BBFhNQVWEvN5XTBbsJL7/yJ8JHkKIdTAOI8
UwVtgyXAtmTXgrLBhRB8OZMzIYhrWxwqsLpN+7n6yay72kLEC6W/XvkiysdLx2cK
XNcWalNy+6b74e3DmHd5XL7l9pRr1PcE/tKXgu5Izw8313t3qfUNTgbmvsOVIFNO
jqz76ay7fS+i8Ix3v6fp8DYDAmKUsgMintOTvRZBzaA/EMAollHn3eyZwXgQgw6t
scEmHlrtt7HwtdZGrdpDetQMXZebAx8foLr+qul59wFXVugf5nOpqBx3hQsklI3Q
yV1t/H625pAqr0OOdqXMj6oH6pab0ZAgXgg6Q8TfktD//SoOkcgQLav4EX0AN4nQ
3r2R4OOJEXTS7e/E2/oKv8IQ8VVDH1ujjpLnEQ1hKHzytgP72qt3paPkB1MnhqWl
RV2cIMevWSqX37AICwaeiBXXktgST0BHnCbE4xpzBuCvbU5PBU63M3z58KMFT2qu
jD5Fz9SW0K4EI05oy3ws3mniJEXSX9huMfCjF4cdJEXRsPoqdSBGZfwwEr7WWBHA
+DptyfitVqtI5yHD8PWP/K10gucLxJa+YAl21utR7IxiM4fUuwYq8yTl8VDsge0Y
0nl+0a1V/+1DhhJEUPUmD6WWDSi6807+rANa8vO4OLSfzKHaksSBnuvJFJUO/Rds
UNPwt/j9YtG6pGYmflbFWkkVdSKME40+tEXnhg12Mb+CpMmCN/5AHPkfacP1exio
gV64AslN/y4g3Hos4BjPC8ucWQHn4Ysv/4ghQ8TINHb+wtwEHYkMqIwBONlZTnIA
UjgzTtImSz0CTnKFb11dwdtyPMshZ8HkoFJOVm4yZpnrh/+i3oxrfXFICfA+h0Xg
8BpuqH22T0h+sPgu0B97AwqCQl6LBtJ6v2Kw/H+Fan38qBRqIb3zmMVNceYntxJ8
a2adQ4W5KofV4e3ZUmLcyGCJy3bepQAFGm6biCMFmPoDPjX1h19kekWPTc5osiFi
hZhdpAB3z9St4jPBF2GHcMn6Aw9xqoL9W49YHEJKR7GGrug7n1p4jwbYb9lfopQ9
+i6oRwEXoLVShBt26PGtDgf/mMlQsZPQJrq6yawpWyqYGwIDmtQuOyjWG6PJc7pB
U/8xsK+cIk8RZNgDNr+m+RlkPqorZijTaa9uXiVoRNqfPm79mEb+DDz2c3HJEcY6
EcOhbK4qZVS0i+DvUeKQq/yfemqtzsFVMm5Xp8uc/EkgwP1x7c4Oji8fyki47dyH
ffpTCgkiRCdzr0jna+U9AQ5I5LI0s1qO5V/vrPBx1k9v6ulmmFdB31VKxnF+HmAC
u/lIhI/xX/1qlBXi7Xt69HO8YJTVn8hKDdw6PJjDHGCgl+ZsZEmEkwkpipXejVAA
QJ+8lNWa6bPcq5dgru/siXNlwtqlkMwUfjqQio+iGsVcWqmrjCwkWIQZbIRiyNg+
htTuW3fJIKMP0ILaBSKTf7jo730AUDmrv2h0nBRCJvkH0TPoCrAv1LJV6sq3wLLS
OGWYWaj6uUCjFi8FGzbma3KXMwuNkHx35kA59sDc4D1Tvgr6mPbqqCdoSWmzFhTW
qlWd1pQuUfn5q9IKWvJ7RJnzEn8XF+W4z/oeuXxfSxxZGlWtuEphmp/gx7/ubWJG
cvqYuj1LPZR/MHrNSnRotuKX+qn0UZXRpUP8roBno+9Ml1wH58uLscpN1VTeROtb
8/8mWKSoTrZVW9keprZ3uSIt19dTqfiK3Yw1dOGjV9Ar/Mz2Yf2hNqsNMpLTTNTB
L4eQJi7rJu/smMSZy5j1LwTJefTmrMtuoOrJC96YJzS8QnrPTDqTn8MnahfqQ4Vm
qKqsCCAiFahKd2eRsbp9N+jz5g9VRPpcWGAWZ18wzCxkiCBP6piXOPJ9zZD8nGWs
r+SP6nR9Pr4vr813YrSVQQ8RexExem9Zy65DQ4c3Kuum417xBgIA9vHRf5aQG8pa
rUceBRn9JP54R98azaHh31e5O3bfWnfLFqQzO5yaCIdGdMQ5PnC+MaE3eKqHGltf
DZPWKrcHy8n9OgDb8cFpytDBk4IrUDaw2VwGIC+2RTLaGLfdvqJFfRcHakSoiw94
JIvHjnka4bTPBzfBpuxAULpq9YOcwTgF+GfVpMNvg869DZIN1i4X5KZPjogfjlCa
ZyukGir4NpY+f2vbylyBFoRQYJPq+JYbzNEzh/9LBFOn/vnRC34lL/iRdNi1Yy61
MPZd/nzGkArZrGhqUYl/YdNGmZRIUoSNb73qSZRQQJVF8C7IhnH1Z7mJGlPZUxGC
K9aUq96HA2HUXvxzIZpbm8BkwN4aP8Bhj2EyZCkICabaUYZeVICUWwHXRgjkCL6i
mJ4qDaqAMr2j/TeefDp2sDYd30u1dp+xCXk+4BOP6oY7KFKo7vztwesI6XYot+JX
hMA5YHmpdLpiAS03LbGrTKQ7VL7BpW419ckVFZGyVvxntuDX3+wlAuYu5f7ULQVt
RStp7jHo3VpKTiFwhsHGXPdvj6wek7VnfvF0zuiki5repjJtk6sk98LVTUf+6Eiw
FvqZjGJPPFJb4DIzuUweNzNxrw/EO5wqCGm4mTXJ1YfvRMD3MhFHoQbvq8F+cV9y
Tueaj3/Se5rcTpIaCmAB88ezmiXo6z+wLD+lMIkzMlAAljKOOp0wKmCmW8mcv1XM
YT1q0xtfhgtBFLPdn0XgTKIhl5NoL08IfkHkPPFqNZC7qLgC1TkZwD1EhB8lSDbv
aURJQKt5WcrdnGhitQv0jX0OHPzdXtP+opfY64h3ysVVxMHm5X6yjHyFjYdS7JbJ
7NZiA/tXUCDvTjtpsyWNeymrmcOyk8s43lrykl5v/hdwFlwPF8TYEYq+6hPgkQ6h
Z6ii5ryh9cTim83sDc/9TqHMyz5FWCD/i2PNFRGQeMlSnBBPfaxSZO79wxQTVGKR
H36IOSywznjbKoJTH1Tq8QLGeyi9H2mzDIEAA20RYSnlVlWSHpgXJQLdwRADI8va
nor76j59zOykAP1Yn/XXsQWzTQUUAMRbpHEyBOhEZbWZRwLT9mfkVYPCb5u4fksy
CKgm1gySA8Ndgetelwf989CPm9P1A1nlcbqypLbzE3sewX13ql8ymapdfs6ehRU+
csFtY7oLzcUjr5N9tPLDfvwlZRbXYOHV/W2bICUdCknslUn+Hkw6OEVK/+a/LFW3
ho9a73vzp1oHAaD7Vtsa3GkQ/L4eePlE2aK/k5oLwURA2NldoLE4TFz5VS3qWaIS
M16May92iq7pkOtdNzOFEJxGzx3V+ne0dNfQFAyu50OMZ0CH21TRLT7fQxT5HWP3
dqANlF+7f1GpvsQXOmG1c5RWXbqpP6jBnySYHLeOBO+m6qILOEixNZ3iWoGGJNkN
dXNy2AcLsM9wWmsosbw5hvAvq1A2W0GKyotyKwqiDRmkwnepa5XhbWJNz4INxk8Z
Mdu8LC7Jvi0iy+N4cPk43ijG7qbgRE7OXd6Tu0ZcDWC2ZdbHHD2Jwq5tEfqQc/07
afK4bdWtK4oWdOA6kqzYHZWamCcTx4A3k55tUYKsccaOdj8jcaa4TrzsM9qSndSQ
/1RYXjB2Npe1Ks32d+x3+3AbMIV6UCAAnZcRBOF0a+I/UyE8JVOByzXlMOiLf6wO
+IHLEd68A7487FFVN6UAXG9S6lhLPFCGCX+8mYzeoAqNvd6+K4MDy61AAKQO/EbN
hsVl2i6HQHRsKU5VPKIovji5pEVxQYTbRTraJsr2L6UUBzKex8xw1MdjweaFjkL9
tKOskAWBQSl3cU2Y+P68fcpPqxt3WWdxcF2JUqjXrbuLbCHe4xe7GAFsDgdkmAGR
yMZB/nvhb3bRnwsNtKj/kS56sF2mw03k1RgGFkk+XRu4CUWvIgeST5SSGqfRYT9T
P+yi83YlTc7++vDeVeEvGOzRfIMrLkHNyUNB5b5w6PfuxBFrzd0A+G7ybYmD32yE
RxWnL3/onvp/oPKpYfNegtILHywTbA0in0nhC7VthnBjkWAcE0XWU6xeOczQ/Mue
dOqze3FrCHAmLsF7WMj4WQ5IldY7dJwtwRPXPgSmk3l8uYm0qzgIRnzRv+dqjO35
bPYPFniLpRCa+pUV2BsmPstoybpXSFDL4iqWthTZ17yCXTkMK6AXDzJ5RM+ZX1zo
kdm7bLdjceUVbzY5tqxpL1dBnykEqB0u1KekFJCKoBbMRokBWwtH8pYkHnXVERz3
ihDDyiKLtOEIDNfVYPIExZJtbqd9To1CYaDiLMPBU2wAj/UQ63BR1/gwCFJvzVVH
6lZlAWCGGmIb2pjTjRuN0tEc0yxpm1x621L52w3knBGmHtF6c4NJ9WzULB7xNS1I
PsZlYWKgcPraLWS7HfGQABOI4OK4KtQjUlANKP0Kgmt6mF3OdW8/MTcIJ1R4t1so
qxpVqmRcge/3bPAQDKN3LK/ynFgtBSbor+o3lcmo2gqBpJugcAWi8NYKvMj5xCfR
GCNR70uDBx2ChHH1fOYknkklvPvF2jZg0JNNVpMax9WnE95WPSlEK+lw/YIIywxe
eh4U1hmLatUS3FaoIuy3/QR9+SVWh1XW/clb6IzNjoJaFD8Mx11XwJG6CWGrwfIE
RCfKxgU5+CqmnR3qVQv1tE1TRotD+4dftXMb3begcOCu6NCiSycrbM2lsliZEX/9
W5WBmb8NvmzAfi8XPJRCKRrYMIyVVeB/bsYs//zmFhJmRkSmmdYWhB37b6NCkhKQ
RwjmmsX1tvwZttQZPsN55eenF49RzpVLKnAQrRrNXY6S8vj1/jjk7y2N9gZgEbRd
gXlbBxQ+Z2BxOoPYvZa1+sOaHgsFqNVtCQsh8AvahR3VPPTeDCgMhkG8E3AhVzXh
kRPc41JVcimi6c8dPG+U/D2etaVWTTgy3rryGSAYkCQGSpBGxsTOmuMCyFjqHzA8
4KEB/IVD0pR32AgajXZiwDNRtz5A+5dx6l4PARm3/j4eaZOUqxD0pGIinKzP1kwH
FNqF1taFnSAAktf2dxJxaGZvTB0gjXs4YgnXCSyNcmqbYBVtOdKjHEqJXqn9IEK9
X39iwCww6159Og0M/EwyGFn8b7fSVbmwKxw3f+SNKNQCHhgEAFV0QJdRSP4a7FVJ
sv0+9T6CSuRAKsnaodvEcSJP/Cr//ftKd2AO+c9l7dLa+caegLfMw7gNlXE7VTWm
gr0qQ/KVufJ9LgXun5H8HaMBhfD8YjxA5KG8dDy8w/WDWI/WI6MVYla+NjrpqdlT
V6i2LN1KXuTaV/TrEHuWZyxTa921akcrvYUBTJhwt2EiwpX8Ejlmul36VPFDEjgB
irq0MhaElUx4ZvQSNPVPQ3cYGSokMKhoUDA2LSzJ4cKHmaLy3hwodfn70Nj7Wtso
T6dFJBzTa7KzUaSWX0FwbAQTlJpTWwZ/HeMAhadaaC+vy2WQNKnwTxtvtbYlqxiw
GnThOJ6tKZ7pll/AAOfLtfJsB/dBcCSRg8MX9uOjADPsqzOrA6Sk3TRFbMmELL30
C+iiJZ5DggifI6fhfn57zZEhCohXQ3xM4lLQ0J67X0b+gFy+rGgUliw10URHGqfV
kTDMigq0ICqp+up5JdcmC4qOX5Yax4FlMyg7WaRAYbR1Hnr8B1vwQOpfW5hXbYaS
NCKch6HJTT2ebuFEU2pDRSNeJfRhfoFsC5ig3IVyroJOdm/C2CSCdYc1U+jVMtaD
mRWnNexejq31mAJW62W9QQAwNTDKXmhwePjM2tYKpLsOINPs4X96jsMLBOs0enq9
FmyItq7xxMJ31cgQ/lVlDV7bS7iL3dxrb3WDbRl7JiL+pEBhMST3ziee0ITEERGh
4r0/m40I9CPH3jiXINUG1HBOJWRa0YMWUWJKJlESzB2eLECHjufBsgPtSlyNi+au
USjD4GMyZBv36Ld1xGm+P2FXDn0KlVAfjzG35K7Oj8WonLgnWns70jxPaVLkwBNm
aSVddY/YmMI1TyQR4fohGVXdgD++v7aw79NKK76sjS7Xb6HWWH/cvsVuu/kY2rEG
1NMxOFRP+NEaPgb6WSF0kEh/e0bRUda0CGrzvJjUeWfEBmxADgpPeWLg7WzDtK8a
mmD4l0wrYbw4v+R3Y4wDKl7w7nBSyCC678DEnz+Hr0mmxul4NmGlByGnkwXnkg4/
vYbbrqAftP/Xi8XRZRkMahWlxUEZEIAj5zo0DIf64Zr3kUmR0x52LjfmmqqlZFyX
Op2MT/jvnzhR6QHkDWLzp8rUpKYEcDPncmrMkY0jrwrxnc2+/XFtdYeElCaNqsf3
8K4c3VhftazF4zaCKNMU8w==
`protect END_PROTECTED
