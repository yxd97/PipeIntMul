`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAczraFlknWayooxB7bt7Kdvbei1IZ0Kjd6OD3zl3OYkGmHsi3hmAUW+JuPlQJv4
TvT2KhwuOl4FqXD8HrlNy5o0PRJh8UX4/oPmHVYzimXgjfxA47BsLDss5Nx1ZaXR
mwVBaaLRmaBle/FnCqySECLaKod+VANe/ahsZb6jiHPA+Z9RyB+SVzNO+mFn8UIb
Z6aFn14MQLzE/2Zr2YRGYppq5D/GdbnhpmsXWa3CMIXGfzFajBD8ctuWrJQN8d8x
XIvmqlCEPyIchjXgBnD5cFkXRpsvDmBgYW7vcZjxP3Hl+NVUJc0PibciqPSI8umA
KIBx01HZAqnys4zfks5QpDllpljSmkwNVtoPD29EETbVYWuw1hir9y5W9eSsEaAW
JAzUFo5rZzNOGSsWKgY1dCxJNgAVjD0ku0s3CnwIpAZQNpPe20FzYAfhxXGI4ovj
KsDqZAug2PX/E1LKSO3aPqYWh8gNpqGjZ6iPHTXJa82ifRasiEpv8Ddc80Mw+G0t
+M+UxM3Nbwv9vP1+kPt+Vg4m5EagkU/K0ErMji0XIBVt2OQ+BWFEko0las2ThUgV
IhizZFeFVeeLBZLVwamzObqZYp2gMkZgyz15vjRKZHiKNvdA+10slZTP3n6UVMJW
6GSJs+nVRZ2kzKN7avEze9apYn/1JZQKS1XZhdIR18rHSEu+5+9Nd0+04Nu92CFf
`protect END_PROTECTED
