`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZ8Gmty0VAAn40bNS4JjTFjGbhXvfGpb3ioVajTxjEPC+viB8Z8lvn65oguyzgrQ
1kUqmX3fUP0OxtZBDAA7sXNXH0I4BX6LolzDUw9X1/vUaPUCHiMkZiMTXPTWNr/J
/kcsZ5N3d8AVv07vuffGHdwjoSSJjGGGbD9fwJ1lXOlbJCQ+sOfkQRye9Z0zP735
I7yiF9hYF8tgx0mPr9b8yl1OGJCcA3HG527vDgbyN/gz/ae0ftwrvX5ofKH7//Cn
zj4ZiPpv2MyfZWuHBFc9m5rRhCT5blUnuSrvKLs2R0eXHW+yp8fbCrbv9EC0V27l
Oql++Pr2rLGhjPLvAWS2YJaPBHJiRUrnQlXoOgyRwOZbYQThEria5za+r4RmGr02
5ubHHcYyDuY7ZAuOeZhhZw==
`protect END_PROTECTED
