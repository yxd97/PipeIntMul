`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XixSF7i6zQ1pzcmQOR3qsA4aBOFLLdWOIFv2tHcvq2hYa8nUVN1h85kOQS1POvsR
XfWgwBuoqLMWDfoS0L13ske06GgU2Pls/6gkW6XR3p4k7jhArjQyp+ZSrrJgXqzg
FSsglMEPsXPjqu+Ww4EIp3ciPSuvs0fQVxAicEiSKu9+PAxC3uscwdHahmtLOVm5
gzeoAZJh5uyu2i7LyEGUwbs3KJjGKpxfVYruZYJ5NMiM9WoOznpZTAgCRLNUIgxR
KqQEAfcvNb8bhDJOfdPSHehiT+Qhb9x/kbEyy7sZ6pCN4+5FGiOyptzKxNnpYykP
0bYj5yadKGUMSjKKr8lc74FJ11lw6NVDJTlUbG6uB+oyrsWl603uvwcC6iBStDVa
`protect END_PROTECTED
