`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bAtWI/d9QOnCLzTxItcYZ1Qvl1t33d1NVTOCasgMkClBvY2a3kZEn8AtgkEuFQr0
egRg0Uq8LpJRUUtZHFWx/94ioDwdb4MMazWsNpZkqAyynFg1BhEwUp4etDwZQOvQ
oNY+4PibTA2CuuelX7Gk3vnEcIt2PmtsUXxPdODSs71JmfyE/PdqGs5hs45USTbD
7U2h0iWgv1Iv4K4GU1NbUe+GsEuaBgAqjTe6fVmKEBylDvYMlQZTK0eyUIkzW3Rk
PqjtVIzfjb4faNH0jp9vLg==
`protect END_PROTECTED
