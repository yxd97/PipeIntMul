`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ws/YpQkux1jBpYLRLz80B4lDACpNLuPhNshd+YoYYXcP9b6R6js8fdWB8I6ZHOoR
PCy0IgA26q8ZIZN59syaBj4Vq+hbafwGUCJUDtai2ih0ZmNwis6kZ/XhWimyxLBn
YBj0ehnTQ4WlRTzrU3qBt+swpjm0PrIzoU8NCVzo/Seluxqe1YLZq32sg0Fs2WBo
Ih/kPlGe6+TrFCfsW1tv91g5FW+ovT9V6Oas6dlPrO6k5l6VvClaR8rq4n3GqWfq
mqhQU28ley85myCPSJ9C1UVYjnay3RXcxn3QkfXwbI3IaVd8OkPI4lW4vyoDP2E9
W2utb8ERCKJ803gL7Aeo/8VAZQXBKrWoUerEg0wgfcwZfrygjg4QQa/Ac4QdKsB8
2GIaFEiq5epw0e89bnIFvVKc4mA4RpvNMkVGWtFUS2wL1xxa3dIS0EtlbFdKRgiS
N2X15MDPE6GMPr/2uCKZ+z/ybchuimCZjLc/JyaqLbuqYQbR0/B5iFhGNTTfz395
3qK6YsGtY/HSceTV24NJNt+tuDkQgagd0IdaP0ab/dBzSvLIzdE7gz8BBDNzNI7u
aXVQ3EyzCaYcKakhi2ifNJ96nYDFlJfRDmEOgHZBVKp1kPuiqPydX95auwgIiihv
X6jW9sXWhrhvvtJOBLhVRo3CHPyM681n73BqnLTEhVD2D2kB6RSPRECPUhhIwu0F
j+b+B6J7Mfri4N+iZa9npYogmcY2eMGY33EN5PnLSlNFKrd9PmojY9ChoRiENngV
+s+nUjDYz2uXMCmGZ4k8lAy51UZXpHslw+q+XWcr785GeNUTGPWvxIdt1sqizzP9
ujvtLZBiTQZiwUa57WGDxWC1OI54M+VHB3gymFxZX7sWDDipAIelsCO6Anu5k3Nb
pa2oR6ub2kh+7M3BviCKarpgB0N96EMG//Y6wI1qHfyLauFul4nDfTFyYVrtHwvv
yyLh9QooaWgnNtbf1A87NAPcTYyHEFMjlB79hjBZ6g9yhJ/a5B+oJEvVoW2FtDpC
vZPPA3iwMPRfUDD0pPNIOYUwozNrx94YaS0XaQlGJWOyfj4vqXpyz32RFaRXRbN8
ZVKMAARnHHZBs9fbF4xGFBAbb0tLN7Iwq7W7eo4ptWC7Au0BkZDB66yayh2g/Dw9
VEeyFfEDvKBmVJ5EQcH/X+INTi4ZAU0QMjPoMT+Lp/LvFUIo8y5d82DKva1NYvDi
tbGmTtqMsCbFrRCzhZ+Q3fFDH6UzQ6D/i5bNzQ8lTn79VknLRupHi2GnA/TLCixj
on9dLuv25gfH0fT8t5c1P+OULTcyuWARNgJWk9B/j1MpomNDMZoSE+nDkQrC3Hlp
C+FfqOEN2bJ/kIxY+qqHLhGOYHqNmfL7eCis6Rq/ye0w7QjaAf0e2V6an1exwzzT
4YuDZ3tnR+mHODqV5vs+SM/2ja9+bfFbnvc4ZSDBmLF7yumu+HjyW4zTeNEzhAmK
bbTnkcCRwZq8j6O2yomjLz8dy9jbz8wCqZZXSgoypHknGaHSImGacZDC7x/RfP/H
yla6adSsGdkqkwotpa/xC+leB7g2thswPwwiACWHDHfqYCd5WQ0uUd96ahM8qQpD
nVoQhoQE89jub3y4hNtQ17niZtDpb8Y0WeZSeqRw1wte1XY1AQTiBOTRoYcQ6LJS
xYgbdD9758s4esv7xDpFDgHWb1qkpTgoPpKvFl9TbQzaYvKkZRqmoTqjRNpMXFBZ
kbCRUFsoFQGI+33xNAeCrBPsZswz53fI6Qw2p/EZOXe4Js9usuARG4zHcF2vS4xI
vfdTVXw64K5PKzQqW6wnAXQpB/TMsK66fbkUK0aH0lA1op+fEZiLqJHROaJsGbxr
rwQjEof1gWiieoL/uPcOhgmmTGKjTftoS5GkWND9x0BN/4AjGVqehLCm/ysFRKOJ
IJiVDucuigEUH/J5xkx+HiEmwtfqTLxqw64jDjj70wZE39lyjTqmqNLTTNKjKZ/W
qOdWMdkH1pXb+NPzVzROiS8pAnlT+QGtsJML0ABxaJ3oJwU9CxHew8bHi7KocOFN
GEdpzp6tSGrwStYvVtWm3HRwA2WoWlu3Ts3q72REIqPVlI26cL3hhUU+6uxdbzka
iFCd3WxxeXF6EK38N6m2+4jz4IUQtYDt9s6HiFdG8d7iRoFC0BiSgfqr5kF8ZpVL
DgOrDfS5AvwJUMGncATqITm8yEYCtsxuvtqOv36o0Wyie+ebRCgocMCnaB5NAweS
z1R0SC6eRogO2VCPGYuCCpFqj0PCZpRIxl/q85RZnhu2Jzq7wXkXm7ZRD0v/+FoH
tZzEgnKjNqnNdMLB3K6Wp8DSGIC+N5xgCP6VWgY0M6bAmpf3B2cpUbw2ZaqVd1vI
Te0wUoxZBGMwyRcrs3s6Kk3bJrP/gdswovCg1xapPnEAKC+s93+IAkCwJO77+T8h
AL1pY8xVQInWNXwoBEv+6vYs2TZObqXLK1xz3wsQOu2Of4NK9XBjk25QChNQ07FE
z43CUnGwErUJocqLQQZBlvQCCUI53RiSkwwOu0iFs0w5xV7gDMdj4fy0K+nfc91U
SK5ujaaknUVGE4/cCqSZRU0sh5R3VHNYXOXm+quVurArX+KZ+yesx+lk1zqRsui2
D8F8tp9Ag63kStW5z2i0aaGGzHhmykTJ34yWfLNlS+fuSBcoqWvuYDFZ/7fkTAG0
YUyYQxY5OWzVCOwv6b+GvvC3NgMhl08Kz32bqotvhAICwP2RkFBcn2l1nz/Rf/e8
Re1sy2L0xnKbZswO3dCF6Ca2NtsEevDsaGlwRHZDxdEIAxkZEG6b3pZ1VJDMkyAg
NFmFIPqHZe3KiMoVIbu83Rtvd5mZ90Osk3Y6KpG8DUeoe8EwO8nIOpg4QdxZ44ii
0e8Hb/7qH/WxEmiofcqvy9Bfy/gO6M17RGK3hZOuzIUv1lPSKj9QkT6uidOGpDAh
AcsiNt8w6kLiDLDirDn8/mVlqR2GxBFrQnMhXitsHTTCbeAyeuwkNnuji2PzjSd4
tlKo1KsIH31u+UaWNkdAcGj6McHqFMRNLQsKHFcGQH7UnLH3tWoenUz8jnJdRfiV
HqSc/dPsYe8ep0y2V/V/EKxxMmFS/cG1mjzZ3nBFfJUYsFzYK83e9NQBkiHqegqA
tbyEHbD4j7PAqD+Wmq5o87Z8Vff1xEuX1DCL4MVWiGqif9/OxWHRTfa8ShwjfvVq
yJ3XMm2vR2qjkBbKlXGlBjijX3VS/tucVGcRHn6jbJS9NnHBXdSd/CqLT+vS8nSW
RLpeklB7OpGy9WnzEM64ZkpAX8+pJ+tkaTae/FfuhQbIp+RBElrBnwtTxaWuTpij
E0OsaCMFi1YinLGOGBcyQKA//THmF0Y/Rt5a5sbReqUU9rpMWNt5z+CpBieldN/R
AP4cKa+vTn5uWlfVI1tV60kC9m9kl4jis3EcvS6VuRPa7IJaxcDwIDeJn1wq5aU1
feLUzKJXyPvnMB6Y1T6FN0INjb4+oOvcLkeQnA+axAk9NjMQyFsz7rXVvRZYEb7z
eUzRYPzD9aemqJBF7dkTFrQRs37K1Vbca1mIHnJ71QNnORwCHRm2ajjvtCPzcL7N
Rw7zkeSqSxUwjHFYbCTYku+S8sAUChS7JLthemwlCNBbkm1huaIZW3/TDcO5fmdZ
eqFpNJoT5E8fiuCF6/7iq2Wsql8p8TxchaO5lGDHwbR2LfIoRHYXkFBuoehwJGqs
472lCzh9F8d1e9yLWTAXT4CmEq4GcBArcEyPljmMELKK1FTqp+jVdccKDeTPkTJz
W24r/+LyC9+SSE0wnb2OMliYbmLVin6Y/SbdV+opai6OdEaW50CT0phviNMA9Olo
02dOpgtoaDu4seMuqLdn6dj4YQjYUgQbxT9t2ml2FJ4k2UsoGeF+Pq9mrUw5sgLd
K6co3X3WCbPU4uvLbyUzrCLqw7bSQuPH7dmh4EvpQLF5OOaFw2SEUiBU82vBMAHp
dQq1z3eXe+fgeu+ybltZYHHFFEMJKrECWPXBIBZ+fdxhyt3e9XspjHPsY8wSHM1z
5pXAFWicGKqZX6fmX3x1gABfH9ot9O9R9K907bB+1T0UxILbEa5OUviVNmyTN9m/
7i2tEy8j2SI1fpOOvG9d7iH7iWd+rmX64Fv7PEsecQhOluGDGb2WfZiQprpvcFS0
6KSy7Ot9RiCSeYbZF8tV9LJIhf+KchmhJXWrk5m5GJd7R73VXH6HRisSBcoY+jvd
WXhTUuea4aevIxnFk/HFtEqC8PYm3hVF/yKO/jsX0NVcd2b3yahTvIQt7CrDq1Mh
HBh+xwmk0sqYtgIky11Dai2eJnlG/jgx5iDNEzJx6LroQAREebe4XLCRvt6l8d5I
Jc5pQv9YgNq1IzLzMdqEEi8/u1gCOAW9ESNCGgCbqx8vieic56qlr2vcm7gO38LJ
WRhWXI0nNFOxxvzmKeaIvzc1m1kxcYAavWrO1S+VO31SvUz0UvqP/haZ5jWb8Mj/
7CYOk+zNEcmcuur5QaIK1GKTkpqVYCWmAGI75Rqroc48954b7cwmcAg5aE4rueCJ
a9uwQqyVxcdHv60LjzGvDALjjkmvobqjm4LF0Pqtx/qvBMsblmEq/y1lXpMAtjWL
JXJIJSpGtkVJmk7LeQA9nmDPeQGExucItoTflwIwqXoedWZueQ8JosVAs03Z1qOB
81aJnhLcl6UyuAQiFdZg4cuyUiVK2xYcwRmR4NMn0lpRFchz7g62AdkxhEB6Z/ha
nyVtiGVZUvYpfiXvJvyr/XuSCYe5N1Grhmagzkcpp0lqZXvj6Hu8tvofjOQFFlXf
LhmUmc/rXyobskjRqoxrSngCQ3EW9x3ONcBqupp+C0QF9fOPvWJcy8Vu6q6MNlaD
VmzXQFztkxV4ASPC6ncisLpuYtJqB98HRb0V2enu9d2QJeGGBOHdm05CfcHEqFC9
N/eTqawFX02Izz+90uKS3RrvxC+/RnTVnUItGTHEz21wCUlM1oR8055F96tsBRG5
gGQwMet0wYKavAgY+OIIHEWrYvgP9UKPWWkPVTSUyqZAuRGgL7zwJ8icn9iEtLQX
wl730i2tB1PItTRqPJCRrn2aGqdDfcFoJ7kfOzFo1TRPeMUXegj3reJK+f5uzjbX
1QyxUcjc0MMQyWvoZY0vfA==
`protect END_PROTECTED
