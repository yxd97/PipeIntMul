`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmksFnI1qn7uI8MC5efOiH3HE/OIisLPQ5Ik79aslrF+fYCEsAP32JohrCVhOK9c
3D3l6l3ErWyvmBtPb/FXLRjhz7KpD9DSdPy998+7z9/Ab386hRtcstu3rpZwqOLG
J4rnz6Rsm2+1EKWFeo9bEZsxSrWfaQTg4LnpVymMoUm8vyL26GjCLgT8f6z8j9ln
aN/nY9cz7Ebdc8vx8B+78R9hfJy2CxZjUWx9cd9NsRzgB63vQg9NowF5KfnjE/Vh
ohFCU4iIjVPb8HOpSdshKmlZbBh71eBLvZmslhRUPHCrjcam2L4L8EnhIR53FsGm
9UN7g+VhyjTKhmE0oqqjhruWMnT5SxuxRkqqqgQd4KjM4h3RSJ8LyobmekLfFV7R
LjQDYqBu+ulbwyfq6+dqbUAtYLq4IQN+4AFW48iMgAJ4O/f/bzPOoToYd8QCWIn5
J7sVwlOoD2UT4ycsJenAqHyItS7usj7GReWA9q0VHJYxWKlSjkGYCVPpF6Et2tmG
vYP/79F9iKquhrxMrV8PN6MnvFQRgYi6R1J35iqJpOorQOPN5Pflklf4nI1l73Mh
9g3jJH9Qxt4+fbfEnOhPEa/6eTdOTuqaL68IGpATMQP8eN45blbKljKhBiBV9DhZ
JS+uE3lQ5hb1Ntrg6UGvfoMXQiHSuMU8ibOxi6/UcvQDyGeZlt2j3rfYvvBFv8FD
PU3ynpCIhT+KpvoYuL1TojJULhnyf2apw9jU0GuPr12tDxB+k1XosLse4OingQFj
RM7+kEyyZxoKczzAdnwhZzVR8Y7X4TrkALSXnkFzW3joeoOxiAxWPvXcRVbEHscl
RQHBBktLm7EfRr/NDMRLls8YYKyYJ3SRlkUE++pL37jm58thSyzrjtDg19/sxYhv
8ggAPxN3XGK51nKvyGcOghp8f2/zLV6fUVkumoo0pMYq5vBoT+0ix0xbPJb7YWs6
00Gf+FVxy57XcN3StVuZ21MeLJu/pBt0yIr1A1cHa2GqbAju6pQMTArICNrOp7Hz
uOgS5NwVO/qEzIXnkXXzmHER3LDc7UJnGeqQ38gEIzmh0mjpvNjbDOiv/q/8qjkj
FKf+qzTqDDEZGuSipbq5wCj/grtkw7ZtxdeHKP+26K1cS5tuhL7lCeWbi9IuOchJ
qsuhmGPqCPBFrU46yh90n/Deun9FVEeQz8XwLyEW6Ptaz2JjAoTmlaY8eutkyxH5
AgNRsxsZTzCaPRucCfKmSnD/8nDg3IHVuLymLuchqLELm0yu/j1qu+qHMXVC/dhV
9knu9ejdS/Q2OPGbHMOP3jRA211prTNOSLzyOxvxRcaVlJizFjyaMiFr4CVlb/lk
1n4LRa8mkzFXUkz3anivCWl/e+9OnO4B26hSkB63fGOmQoAEY/1Xp5KyecJlEmKC
E70KWfzfnbtevqnTsdYrgnUGeXTM2j1evcWqQ8BIE/aX0BOl7PKRmbUG9nFHQpr3
5hgaFM5XzpRY48Ex+I2eGn50kiEAbk1m874psNyjJcQBzzIZDCZvPgzsy0Qe0ZNT
Y72D0Ytt/HgBkwYGGYD1seLDzCbZheHtJiMfWDFkaxdcv+qhxqbgPTjnEeknFZ4i
Pd1mavFsnUE0UWCmOzeR4J46AyJyQRwQRqw6yHMPvOLLGxFEZ500NcB4TH3+gOB2
vgVZbjYmOTRNKuZBx1KE41L827m/retRFn5husmBD9Buh4uTcaFGP4xZtkDdm99k
G4/7vp0estcuAYHqMooCABkIHJ8c0NDsXlrkn9FymL91/9x1RM89veIlDcPxMIvR
1rN20QRsGe8iYGCWAzQ3V+fd3wwROkFaYq96bIne4JLmesGjR6pgKLmO/RxaJVKp
tlm88Lz6Irm1K5o8yMkC8srpjElYDm9HeWPXiuh0aR2tBTapBiPoGPRbNfRpS7rw
uXEXo+Ta+ZpKR9CIB3bj7yoZkAHYIOa5yOZ9vJHJOM2z4pnOC7a4ufvQE4SvVNZ+
HdzDiTNIEp59jduzBa9G6cdZEqlgKeKoRqSivdvIwr1EtU1QDkpff+u4CHDATej/
ZWNuJABe+t1b2cB9GzvGdkb+AWNc5HJyERihijKfDhyVudk5Xq8QgeEuHwuJBJ0h
S9BvE+mjf3ftiz1P/FWI72vNuute6i/zES6GvXckCRR9By4nC28pbAf2rJwb+DLb
lf7tbUCtL8k8oxHKbT7alfuiPkxD8yM46jQtE2XeLvoIb1mSCQhlLrt7GlVTtLBb
Q6WTPYTvsXxB8tVF23/kFSx9BWOLJMmukRG8AXaTIsotOgg7Pg/h6lFze4yx6I/A
kSoFCjYjY7WqQrerZoh72354lF+f58cNJe963zctuCnCoDC6OZetYfKUVxfE3zmK
iFV+qukS1IXlbrZ/VzUWSh9JMwVrFpSm9jZbg+WLSHFpBY9+GIwC/ntfMj56UszS
1vya0/oHFEF/QiVgDReJlcSq8cZbnjlgdN6zWwboPqy45uEUoc163qqa8SgUvMI+
u6/JaLGqy7NozjxezyGoFSMdvbDZBkPRFlvhksrZK1RT5A/gOqvrL6kw/JKZNY30
XTGIM6WHNAVvCFqFFEA+lNPcAHtrBUrFnSt/zyIcWiiBHnxEJvhOCS39Rxrjddf2
k8/YItQHFMZFwR39WD+Vg9lRaMuX8aPxGMr1HP5fTylRI/HRtml8xAg6YZb7TTDD
uIWpdV5tTY1OLOJAoKnd3PGjFVydoj231J68cl2iqjeW1npUcFifidLWOJRxbSo4
H3zirCO35244oh6keMZvriqO7tLkyB7+67G4vgYPeTtE5pyrGXTMp2nmJHs6Dn/2
UghPSyhJRawCi4V2bo+AjfCchpN0mS2U8gxqlNt7tWmR/FK7j1JoRPp3GNHxU/CO
kKATK5ITX4J0/qINgl9vZRivofzwQcN50i0CartHYneMCrcWrqDj0r192e8KRFjt
D08zW41YCh0vFjPJ9Bk8JLh6PYwBtrXVqIBmBv2gEGz+143zbyLBBky3FvR3w5C9
3z3yRTdPKEHlf9VYgjcOJw0xe6ZoVafNMfnMunh8yNrZVVcPVO7GOveOWvxG3it7
PbC4hxc9wKKazPWK2KOWKHD/d2Rz7m/+QB/orAyg5GLc2SnmK5bXOfmkhmnAcq/F
PvPFNZqx/805HzMtEKvBFamCCnENL2pXUCI8M799TeyVx1FU6nmURTD+P0mHxyC9
94bafMIMmyn5fyyLS9bSXxQrVYjr6uN/tFEKS71rme9JtGPtGtYssuCwAL2uB6p6
4bmyhyU6ZNU7dAG0JZxRSWcgF2oWgmk6nI2M5dimszHT783I7M7m6DNvmPqxQE/i
sWplVOj7s8YP+V7aLqQt2UTr1ZUk0WQlMCrMWvlaw6Y2AQhJFG87KQmNsPoy7Ck7
U0lVou5SKpvgFwRCGTa25bJc17AEOsJtfgkh9qH7okeH0WowOi2Ce/UQMYUXtBYy
b1iRrIbpu6U5olO7MPqiAK9QYaSXqH4v1qTahj8OqQ0Z7pW6pabqgDPxejUb3URy
nk10K+vQzs10LHQv2mwi7Ze6K8cHpfmAultRYHynHa1HjvVZ8uVSxTJeJhCi1Dsz
qPJwhKCuVfnnEwINPB5qb5A4YOg9a1rasjXo+s3MBIGXvQ/9AvRxzHvvsUFhSMQq
kM2kIFEHhuwf+CF/11+JwnJWWEdbs2z1gslob+RlHDYSLEHxUado8d31gtf+QvPD
DdKFW1v3acf/dY1dnrPQa//tqLY/YqVNhuuGRYpqiLAgvmvzHSsZzL+27AADPa9D
K4/NjQ95x8N1WsfEnVJBWSTYgs/Av56LteuG5p/O2/s35tgKG39rQEhPlYCvJpwo
7o6PluhFFGBLjIymjKtOJCpsLlpQZgnpaWwfrkAxBbT97v3cTCRVq+rDXQ20fhGW
hcTijkSeLXV2p9pEpr8EKb5EwnZ6sSLiQrGhoeSh/RFItcknilnPErdbFijGFUxQ
8DJ37tdZjA2OpQjQkLM3zagEzATc8DddQ5O+F31+9n6xXJyvgdzPZLrDeDdXIcSi
69ko0Knj56ZXj24Lopt4oNTJOcyvJAccQEdSRhvFEHrNpdwHZ9aOOHaVV/v3X0tr
T2RhpG1iJ9qVAq2DVZBs63ldTkjzE2bALcnVCdn6v1cBjwIuuJALGyDmRu3pNHny
WADhOxBILG3xS4qaYvk01dXVRmJqAZfBt2Enjeq3cqAzK6OaTN2QWicRJ/HSiuS2
AK0iltHE6HDauMeYdyfD6pzfBtRYg58wChyPSEE2D4O9UXv0MmBqRL3qlCBt3tpx
1ksB3JpFEc8dyYEze27BsIbgFjq4mSXGVZU/3bixj52q/q/b1CtHIuDSFD39vXPd
osSzXPTigUwUadWH7l1Z5gZQjjwyyVtgbHufBflKT7wQdYAAjDh5+Tmnjo5EmU7D
LoHf0A88yoN9ay1Tl4FD5hq6ulZeQVN5S2Pw4Ph0h+hzvG7mOoH1Uvx593BrjySO
cqIw1nThG6Q9Dwlj5vRbtbPPDLU/QM8vB5Mh0Syk18RHYrQH//k3yHVNvtWNfTHY
VCAU1CtcQ3+thF08cyfL7IyFNxoLIx0s/raPNrOdElIBRwigM7oJwXN9pPxPXdzV
1FFAQP2EMqgz+XxNS+rwwbBV60c2Jj87BsxRb+f5lzwVAnn6VBkFfUnQdhoCWLWA
uO3N4WQ5VxsDq4zfPz2/esX2ydKY2O4xSYHlfV54cZRO5wzCfjbG0TXz49D5Z4Wy
HMLOr/4U8w09NaOHY+t3LQo2iSfjjhRiKFO3Cm5uS7J5ABRPGlYMchcgcY7n0uJs
E0jX+a+4gySgvxv61vgLkqPGnvc59GjuC9LnXlVhcqLHJUs1qRoip/KgjL5oyolM
2qTeDdko0XKYHEp8BKr9Yuve1yyNeEfVv0QZOk5NJWKCFty5BSNpEFg6j2iELs2y
BtsMi4HQl5x1s/pZvoH95u5v0PANLF0tMYP7IPiVmH9GUp/OyLGCqTPkGYG9rbO6
uiVtp+WrxDku4FgUGPSuPo8+u2+d8rQWVbpVj+Tet9Q2nABIF6BiGAs6uMOm2/DC
L4kjD6bXYLebdu5ICmG4THVpEaXqXLL8V7JN4dxR83+ozXhMneGhj2O0Y2udYtyv
OEABYGLZGfAZcLLDliIRnPQJjfXboiGUc+RIjPTWHUfMbZJrc/XUNDFNKqu4bx3/
uk98cyHyKLKyarvt2ddXI3phPHWxTzdsV9QuLMPb+Ol3m03gpBr7arQ6QiFrd0aC
n0nmXsRpqUM0CUmrgnlNFcSp3og6ON3P9E4AwCd3i8awYeMyb3IjXoTnjuXUa1g9
/jJSDsvIA0p87QcgvJpxc0mRwNlnDqsgPTpJA8S4ggYT8xicFNQqCCHaorLkxTsc
74ha23F/RPe5l8bU25bEQ4QdQG0CMPYs7i3k0PYn2s/z3BF67oEh2m/0vw8i6bY5
tvuW8Pj7nWQd4+e9qAHEMIGm1dEtpRLCxkYhnIJ8ZBtvhuG2pzjgwyi1BHs5EV2i
wllNV1Ubt7rofwUugr1SoV7gwWNtmMmePHLdOrW3Tig97w4ikHQ8TlmbViCesuNz
lah3gdbebkFD4lwmwJO2OIRxC3wqLznLBLWsaC1G3LFsxkIdf3F0LgtDMxWcD5Ft
sQcfl25Nl5cc12EiqF3klUAp+hP1VqApihWoW9TtSJWMfS7t/QOV2PsYyPWH3I6g
7d/3PVspKfEjdB4dQ+UWvvgNJLTPsY4s1n0sWq5Z5ZHNyJROW60DZaO1PddNajnU
A0soR09Tbm4E33RdWTgHDND6cOUaNRazGpztTNAtfCpbxTeb6odwqjDm9P/I//9+
rIZIZxy/xqyrQQ5lsGqqQ5dm+ccZ7MUwai1WY8glhwmFqVYzs6mvFNoIusr5rufI
WmD6kq2jXjKpast/SGEP0yhwcjpxXg+NmL3cYCrqGsTNPbwR7W2E1yUTy9KfzQ5n
0nLuXi0RihGXSjahC/Vk0JbMjpy327TTlA38X6lrXoBR3QyGA/OT8BWVg26dG70L
mGz5MQtCugA9YZwiEmmwGTRu8+1Gg0Vu2B4fgkjG8GZ0t+8nTQ5NdP4q+1Hv8C4s
N8GjYAf5vGjFcDCOgbkOCXwVDMKqB5xeQBuaN5M34rH4/hHh2qlTZrmCmkm3Rc9e
Ghk2Jl7UcCRF7KQUAoJnCNs1DNBV3gxd84c+Nx1+mOCeWLHVm3zTPH7M4zhIN7qk
YGy+hcGVPKYT9UleawLZrMGJZwarGWuguneX/xWaY4uUTzChggKv1dk0g0zZHJgf
72Wpr28+IzukIVrECNmlGebHaSK59XEWe10kFPcId/YvEVfHyTkazx77rag9m07D
q8Rb9S5Q2C6UT4kRulrR4PxAzFwY/pcyrp0oT1dgqsy+dcmWnZ1BGzm+q1YXvZVO
Tr5IuLkLY89+8PSahCOQjHy1r5MOuxzsYkYqIMNPGBgQRfLwVQj4ZJsFaaTAwJVG
xS2H5cgJuyUkJ5qvQrafHckGK2CujtxwKRpSFOkHw6Pf/zrphxYVAYOtEtwmvNyB
hWDmm83Cwf3ZUO0V4YgWHwYNIn0r8xfDPQInCnutYF+HvqKw+PG/q4RmHLUayXmJ
1wfOUyr54foIC/JrudrgWa6TEqYjsg+KnadoPm+u2zRWtOmJQqM8eFlB0qBBlxWM
9yf269BJxYXIEnzKG4ymVda1Z4FgVCL7xUTofM9vx7nPqQ/xNzF0qT5Ke1GAIGsg
XER+Fv6GpYyQEusa5QwyHW+12tH78E7xJMgutBOzX1Y9SLP8WXRra8V/5Jt+ZQrF
bS7y6OJbAltscAEuAtO8ljHFkMatjhQBs3M7DQ6SOCu0Su7rX9Lo+Fsg+z2QHDGW
Ih+Y6uCjLBpaW6QXRFN8D17uDdYACnHZ7hjwzFst2AZ/8xfcEcAThS+G3fhntzp+
VpyoGkFfj/OzhXu4DL0yG4/G2LSV3rjew+Wr7xD//5sdD9Grtxbh0U75ccD+HUBv
EjW7PfGPBkPMttgBKZ0bNSyt428DpWWCkcsLae8QizKw7CYT/MkL2pJjJTIUCymh
tppJEV5zpj6UztWj10jr4ezGBxVOor12hDdp2iPmrI3B1oX0f2t2snf4TSpmVuC3
S8mn5KiIsqjUIVQyPT3dnWB5l0Jj/KdAbb5yAqjkD1ZqBsOHaSUaoy6CSn/lzmu1
Lb0Vs4h1DQW4j9Pz44gc+xPwtVCSNrbRSDLe2iAiQFYUvxp5CD/ZmEPaQ6IstrMY
1kjLZapJQSZtQNGFARF2ptGVbNbMD4P3/l68zdyVwInYwTi0+uiZBNgMY1Qdb3ks
NGtRpBK2hfHxpaF8VrpbGQNCWMyj6yvcWWNohGiHhUU1yxZZaSlsOtQQKVftup1e
+q41KWUa441iJLkBsWALK7NBsJU5bdrMqrIRNbpPcyVYjCjr14gZAMfu7M0bygRu
dCjnCHm4d3Ob7CjsnHgf0D5hJ6O0j8qgir6tBTuH3QbKTjj8/qCMlZS5vE+VkxLa
dJpbWxwzx0fuw7BWoBjH9U0t3orjI1t9M+cqGtJyMI/B07Ao6Bsboy5BUsEoACBY
10wzWCNGPe9WdvDjdjTgW//jvIALtk2KTmwuhQo+uJLqxi8Ua6ayfj3NnF2Ige52
ODgn+QhYrHZJwZ+L4wNmTXRtszbxNGZ03shwa/Lcx7UdnMDH2OU3+h4sjrACnwcJ
S0pE2XuYGLjEwzafBsS36H7R8MEW8eOrx8L0UD2InZwmfI0nfbp/JcXru8gODKLw
0m0CLeQVjIA0vxuHy58D6+j1PqLPMpGzei/YkzHXsqnzKrBRXO56a+PSc8X7Pwf6
/gz/dVu/vksrQzhQX13e+YPLF6tkZJRc1Bc1JXUA8t4/xh+UNPAueV6p2kJz2M8w
+dy6IeAKGbRCC95Rm1SHx9d4/0of5dp2b4jBcN+TJDI3CURudkvv0I+9qEN6SXaY
r3bvWqj8HvONpCbvEJEvhB9KQFdpkXSOdJvePtbkGmNec7kNneVUZAoZP28qyPfJ
qJyDSSC/PNN1EmVq2Km8RPI2IbBxHAt3EXPlDAtS8IjuRq9Z57RTqmz3eigPF1sC
/rau5+ret/M7nizdpwg13KWXftja1DdtPGt/6eEFTMbd5GiVq2m+ol1tnQejzjvO
C0IDqM46SUFkL5dBdDRCnpZ/538yfXeMP8STDsq1ZD864tVUKyX94lPet0IZeQBZ
9UpYOPWr/qLdnDYrqOmvDhGG8+KzArQXkK8rBhkImsnQ40977AXWcR+YlbIaeva/
Lo2XlPPtBLAGQ8nBZu9HgIPeybNmspIBlz8nqoSdjIquOHB1ZuXDipu+jMYq3Pi0
WWiX2+Y7SiZJM5tQtYtYClgPdua3BOd+iI9avgJzWdxSnjFBD6P49Ra3EQsj7Z1h
Xml3rv6w5GbTWDjN+daVV3sZLSg90JKbYmsjcc5ytfYh7ucbiH1nkmYWSWzJP4g3
qJPYGewMRtFNCfx+VJM8Aqyq1T4whh7rW3FzeChxa6iQ8/GI7cIvZ/ZIJLUpYDrf
lLQ8hzBJJIKl81dXj31c1soM6GOT4NnP3orfuJxFsOivIIE12QXW7MleY8MuPnSv
eZviKQcv90FI0v1IZb6f2fDCJpvTr2RVY8ylrl1Ut+I3FmkkNZoXaDws2cXnPqCl
tzPtmEihg8KVRcm6N5Tw49CnpqLC9eaAWKdAW8q9YGCI14MC8vLBM4697+/CQ+Qg
ZhmZ5QwEYO8DhX+R/OzH8XhrlnN5+Y0ZvAzugzjDBUevesooe0x49Szh48Ef4JXq
GtsnkUC1ACOo8gNi3yOS5JGWnBMzMIGE/JVTCJV73MKQCb4gGAX5r9WwV23YMCEl
PUld/sQOiWYMPCt9ZOMZUFfvwZmdM36BYlxyUQjvAm2QywtSkPjr05lNoAablQML
AOAWZC0FMG4nhfsj/Knzed4UXJcxD5GPcwB6DeEIe5JoITfx4dR8WfTHzeHjvXPU
YKW0Q8xIgNikdjzptzRGysbFP4vWVYRzznnTsKv0k7bGQyDRy+j0IIX9IvbSK7zL
B9nAcVq0Bghahw0RB39PmJcgQywzqdKzMRJw4Uk1zZ5qnViRaz+MUwPAobvbxfBS
I8oi/M2wFs6+3UA0GEqaxYvZH1YDlHy+ED3ahazrrZQ0Q3iyFUVdE4sZeyEsQDl8
FCMYi/60z2EV+G5fmG03Rk4LQJy2V58tlptLkR8GAB/eZItUGB77DHHzTdBmhh0I
uX2l+2YdBLLLOEA7ZG58GC5IDUWHJlu4DRK/91fk635G4B1XgcRUpwqQsnYpSpwA
TTsc6ws9Pc2Dpyy6bl9TVIoTXsfJbj/Jfo1qo0P9f7xFwTLfaoE5E8xaeYTXG0mp
/kx46izq0zQh27Kp4Wc0V4FpiFfJCq1X+1xcnVRP+rsCoZ6dh0yFn/8aHHSe02KF
aPrMCiBJp1laDPtSMPN1uvPsJoA607GuP9LUaPRAwu/Gz0kO04/9998mLFAARQjb
IF/mzLG4RCJaSqVgzkNMWp5WCiydvSwawb66FV0sdpHSCBzobNj2q5LmLXJD6wcX
kB8PAoJjC7B40d9duKQ23fywnNAcnRa7yk+1uH7JwSEYo2bI4QDZPBS7xenLZrhw
H/RAHMvYqOhJ1XWpDNmVkcRJeOsve/OiuBxHkjZN6MaL1nMX/901/XGWANcrVnd3
tXQYVbtpSt08BP9YN7i5xbk8ytcq+K8hZ8ATiLwyiZl3tl3gak8aE6QlswSWeWH1
Xwr44Wnq1ChU35gRLJgZNAgMmosqsbJYLtfJsZB8QGDBAC7b7Mq5H8Tp6mYkyHVF
Eay+g01TjkmBuCBA3DESX6e+3IkfoOQ8r/8NGvDqZwG+8+1Yyy9V8NWbsH+eHL96
l4ZSBvhn4YBTQ1fYclbOWgH7aHMEkH0cu2tM17+tmFJIhMLSFo1E/42qqtDA5891
QcLPVuN/pTHHrCV0aKuHT9aVbSdICLiagrJxE7k6BQh3xgbx2BL+yU8nQVyw1OS3
aIDDNeUINGAuQw0UfUOG6FzSX0+KB6/nptUmx3DDeftRR7FtmyTBT7D6mVUHouEy
GWDqDL/O9OrexhCoFgkkG7JsqstOoeTcngV+EHR0AyXImAeaF7JtqvgsMebJo3e2
1bQ8T7Wm8fhoczTYEcIRikelyypK0VnrzEJarTOeaZpIeKZ83jLvVc4RygjOFk4I
HTmeAYya8sgwQgfGMM8FKhOTwYXcTCVzcxq5VfFVOEBmpV1WkqXF2XcxNBnU6Ckk
ZJFwIfVSN7P1oRhooSM2LFwlWimXic1SL8+22tG3DaoqIMBHOjF6MttkRjHdXQ8g
d4xdT+QTxb25mcCQh6dwqBBbY6BKPW+zSlluwChQShAYmAh2ocYBrSUQMsUTIthB
Zuk1jpj9cMJ8w2dZH9wkKNhrz4exxfG/meAdH/WGzK7p50fL0sFIKgCgyUR4L/Qk
ZF1VR5Bc/ClQw++Nbop7Z1bW/Sx+bJG9+f6LNzRWfZmLXvN8chSSJtZfzPjjm02u
oZDq0w/7cr0PyFIU8ynAVqe7qNMHiBF9iq5KAzYBCPbq8DqEsIKq82aidqasQBjn
VJzfzD4knBq3s1drgs29n9vE6UX1NkmI59ss6UAey1lm9eaTvtLNj5l11QGWCkGt
jlQVs5jr2AWbl3xaGl1QSsDVL6zpu6S52JGHQlDMTqExPyCtL7H8Z2oAHz4Sn+lp
uW1UN+LLDr6imyy49YP44bKnfTzys/KoJO0ert7trWXgo3YcAF9KQt9oMqxKsovX
ihUstec/hhwwycxnqqEPp/VC+1SAvFPhXA2qXFGQK1UBGF9Ha/qQ7wRwcY0co2Na
MvwMAZ6D2fDZ6NYSy07U875/WQXpIYr/gAjZWpjeKaqiHZQaY6b1QE9j33WmZ8hf
qVrNGEdx09O9aa893T0n6h/HU/JLXNwWf1T1wf6pZeBRQenDzvlvC6NnQmBJaSEf
fJzwd/qTs5K8C4qzxtMuYbtaYXnG4wfVuhAGjn1Rb7oW/ONi/5z0Uqliq4nzwYfR
iDq1qE+g2gCxge/VHZ0eYXo3LeYLwMM3ZTE7G/MJTPC1sIuVvexhtuYsp0rDsB7x
4Yig8HTE2u4a2wuOnMo/mwbWF8oHYjqMlrYiX1Mm/P8wFz1s6OjM/db+uo3Uj1Zv
hiUIM5WhwMHTCWdX2CICaOYYLqdLvqBiQZZ4eEHB12BI80czxi20gHVZHkvptLpp
mKwpJek5vhUcAL0l8ee7iYZgjNnDsDL9BZwSAFq7aeMy5LXG3Cykqb+czhRU0Zj7
lVm1OS2wjg92Wnahd8iHP93+Q0nzSFEC7mk1mdXXpfiWwPAQ27NM27FtGzANZlXZ
GiLeGvj4jnKpWoIZRY98B+YwsisPyk+rxWju9oYAg2abuz1hFdIJdBINKWHsOSr8
d8irJt2WL/DccmvrFIi8Cwv72GKmeaVDuPHESVP9kGKJXdSH7d5++kANNv4PUjeJ
ild1/Hctmejy45JRguTIWWO+5EunHhobsj/BAnJPhL0DLy4c6aSOMRd/Gfy/rTuT
5L7E31r7L6Lw1S+rMbJ2oCOHBTCkNY7zovYoO+ExiklfuFETbbEtHzz4nNLdb99Z
52rjKrJvWmWy5irL6ZnUqKgrp95IatqDKfXrm4Q+PsJdIiIUOJKz0MRjKSitzK85
+FzxzjSt/5EmD7xGXPPQynKi+WZ9UZwjdozHUWYcMwF6BNpI9hjNE+R+jz10UuXi
x4JxA5znBF1m5VE91em6tIstW3/1h/A4G3OEjms1C5FfYQ/0TKZk5MLD9Z4x2NpB
ZptR25Y8qkCXuBTBTqmuySPRGi9NaGXh57CCXSkhJr24znr1WnO5rPv68sQqv5Sm
6Y6Vt/BDnVPuepxTpsJwHUydvmzHmWnn2MGk0RnLgE4agbKaEchKtZexfWTAHta8
cRXBWX4Tr8mlltdmO4RkVMmdEmQJcC7sOAQCkQP7lX8MP1KBmoAAbZh3GvDEfHku
fxsVFaMNCIU4DE952ZQ8zyqgdZ5Yyd5B6GCjTFwIbl8gXGtOZ2lfEOQYzhRUasa0
1Q27D90WB1O3KA53Bh5FVRczK4gKwfjbV3Y1XKmYJynHvZxHWHX4GlvmwR8HwreS
YvbyovaJgyZVXcJqfXk/WxB1AvU2upRh3U9skLAOXAGGtw7Mr09VX9QExf+qnyD7
jzaJo/Xf5ixS+qF4315L3WwaAWupZ99PUjoJNNKUJrDgKPUuzxhTLV9K24QeaQZ8
CQpNZiyNbQz+OTOXZwnwcFPIICRUP+IsAHwcmsoM+RqgdC8h1US3VSmkhM6bkI7t
e7htztxoFMTuC1iPJKJJB4/sJsKfh8io7VqnnFQjX8Ce6olGl5DdYGEt9NJmVl7x
S/PxQRFMZcMvLXlRIDQsHdIKlC5+rW7YgbDZahEF5Xm9gRo5Qhs3PGSqo/p+ssio
rr0yVQU6K5YStCrpunS9tpZdC1E4Co12lLRsRuwEauD2kZiMXGjJg3LgOR/+5QzR
1dwiru4poKBR9Jbx4vwXRk+iYsesQrgItU58UFp69jle+u/KQG3UOvF3XEIBWv0N
CQSsw2oueUfuHt9wfsG6Sfp/Gz+FovhiefDgBwVIS1lrVZ6DviCBr6HlcZxQKmiJ
IybRwsYDVLuvbW7hizNvXgWB8Ab8DylMGTloNDCcse64BgtiZQVBx7j5GkM6AKNq
7MfWM5ivyN35z6kUDaNcOXEQ76j9scRsvEpBZDhJ43EiNPEmOW6HqePmYrWZYN6i
yRHRqyW4QBrOM16/sWaT4VXGT6Z4UUyiM+vrU/rnFgl/t0+X4kWk+4lqS3glk90Z
qBXQOn1GBmHcTo+O+tRytvNPDufexx94mR+UUghiBgAz5QVtyKqP3WZsoulANBrh
vinPuRytZpfWENqnalHPnpPth4G6fhE9H41sr1GT3o4IjZhfPDU4UPfDpeVfl/pb
sUr1C3bl3LLIGEz0DTRGTn+W1vcwdBQqha6x9bsk5K1Ica/dpL4MEPxTMhruo2JY
4cLgrMoPo/gPy189Mo/sTmOkw+JH7GLhScznwPNriXaRAoifhh0X+EJa6vAwf5h3
I1kHdaYDovCmgkHHFcTVhK2h8eEzGmqkBFE52DYfML1Z7HgdwegpJ0JL2TAsMPSQ
vXprofjyQZs/mUEt7XYotyg6HmKaSa/1q++SuhJoxfo1VIZIfZsB/6ONlzdPnCw8
HrF14Gyj/FINu3qSbham8mZveFWdX80zEZo3p7LlgyS894BVRwFSRsg51BVzgUGU
Fq1CY4CiMuXHBkdhzsQOu1NYILVEtUiLBWRLurJVYO3Ul+RknSqNKiLQ5QWtXbHo
aWMfN/MHXBInTg93TP8R3cOAu+Zi+TasIXidj47j1XrGupLcT674nEd0mHSgfob4
OoflH9eRWmAc1qCBga19/DXyLqkdKZrOf+/lksjRlxAVQBkH3FNK7VwLvHgcqcRg
+Z/Q8/pIBGfQf/yVwJpe5DAgQBh43TKVWCqpBFw9iYiKd/fWadELtsWMhKPErfSJ
aZIcelprVHLqMTsBqnsFYLxYE7b6CMnIs7z2FdG6cWzAnBUyGg77GrgrEOa6wsrF
AP0W5dTD9EB22b82cTPhdJeZmqYk6lBWNZKEI7fDcBrZks5KeVoaDrIX4837Sw3v
bJuH+dXfGRC21ZB90EyBO/WCVjhWu2pcZKbD7czSi9rVOAAec5T3HbpXRlivtaYd
TkT76dkBK2SDUr9fffkD2FhGK7tNieitYejLBIWJJy7kQsXPUNiYzCDXIr+jbUpJ
Ib2I5yTn7aunGv5sONf2diqKUbusw/Iz1itNMRqdoD0/heuFKZ2DEG+bbCrV3Zt7
A6vDW4w72pW5PJBfh1qGb5HW/SN9OvDBQghYEdFkaWYumIx+dyx3UHyeLtTDD+AC
g0y8GgVewkYXf7sto5c36qSy4PX390xeUnxu/eMjYF2yudhOv//Q6CvL4kLZ4KJa
wbKwbkIbu+9TLxjmnzVuqD7B0B721YBS6CKOFV2tTaQs8lt/8476AAOp4Y4qCkwr
M0X6bQJHydrR7sWhdqojJs6S3ps1cPPFQMuqmWDezMe4+1l0L7wuyUdt35B2LR6/
5lBrzBIFArkz4mFsn6GzhsEwnOOfzaPeed+39xTBbN9sLD9u9h2xR3/dMhlakq7t
3ZulNOdzXetW6oJPY8LSIYFwGxFPXQg7RmXPh0zWM2hlJi1RJK0WwMEez2A3yYhM
FJoRnF9I7FQPGgPjZSxZeAE80B2ugiH27G8d9hQoLgkU2ubKW73UN3kDwnlbXbg9
NqJekVmTvx5E/VqopoS8L5iPU9LVAwgfLm3IZYpRTXQ6hfgWlMl1r51lswmx+in9
uivaUDzSifGsYEttoQckbkScO8KW4jzf1UrTW+Wf2+C8Rm7XssZAh8IMlTqF2gwa
xyOaCtp7n7ZjepAdovWQkfM37VwL0V5BaWT3Lc2XwH2Mq8zOcZLu3GxKR7ble4Bo
Fbou5apnwDd8x0U+bsYVXUQQfM8dgGYdsFLYsmviZZRM/0DkwulE63yyLYD5PBAv
SoFdZEmhWBMx0hjN56+318kKbqy+05i/bdlRMH7jsuAToSR1pxuRmnI7b2T5vFHB
sbYuPXVFm5PwFMRQwKb7W5B1pAX4DeHZ1NSLHj41znXG7iryC8Tv9QcPk1kALx15
1mQaOJra1HbHA3SNhyB5Jrj0q4i3iHGV+ZPvOUneUv9TSVuyyqsWqLZYGBaH7K5s
qr3MtfaDNqUfyTN6y8TAkON1kV9Liox98utWt19DFoNESKavqf30jcGz10uZAinH
VgK7w27zmpz1hEbdOP7UIvpzwBqQBw4yHqEKpLtMFSTfryGGUiz0QKlKKoSiS4AZ
R6CkXprZ+seK8AnzoUZpdaKWhEZzZaVEThndTrklDGG0rdg4av1wC/EUST3iOPy1
sR7ZFLFDqbz/9BHikOV6q0jVFBVlXq8qi2lwtxEdAtxVRS0HAZBHD3sLPZsP9yN4
Mp1ceTJ7lfz46bKl9us1w9Dyz210Gc27y2NyBJdrGwmMtyqK96Mob2E36mODJzf7
I8dWZPYK/chJfKnhemjUoCl1u06Yk9NASk3vdcrEL9ktXpZnrAompXO/4exzVuA7
vfcNKVAwHVHJczXkU5G9vBGWhQrEQe1oYQ02p0Ka+rv8h2zBChcqwWDGhaXXVT6W
vCuTG4ayfSX9kah1aFDExEPYvJGHr91XT4LvmqDb+24kz6xExoLmWl+eG6NuFV3k
ZvVQVQW73jDbhiJVow8vhZA3ky48uCEA5DhC40fC5DDAlCdIzI8nKvydCRoSqwpE
1KX/SDgvW5K5Otoh5qXufJkbpnGLD2SYWMSGGQYDFKc7uk/Ng/MQBRw1CHAhcfJy
2liwWfiZlXYgI7FR1EizNmvMzP/Cx5qkwvw8XGXllImucYWHl8MbtCIl+Ftj9opa
x4y9CKhAL1ky8cG7gmL91heHNXLyVVa/VCectiLyus2fHxzQGpyq4S/CKV6RJgJ5
6M8kdB7jQCe8xgj692bcN5YZxgh7A+qEvxPdOosSqDqtb05xPzzUu+KiH4IwwGgh
o2izBJPAL9QkeyMFkvJAMb3Ubat+yffon0bPV4azh57vDERlBgu1E586ivjBl11U
+vL+Cgl4QFe3K+I9PCdbOmXffJ2n/Sj6yFMya76EpNocu3TFrNUbE8bqUahTRBmP
dCgQesfC0X1/HqIY+hdFALa/yVyaDvIEs91U2YBjC/AZ+QU369Bw8x7z55lysXBl
ZisxvX1lwSsQBVXowUATuDX68LqK6WyHdbVECWfMNKSX3QpmofwPKkeq7RzeT36R
HyGcZ9amVLTV+8Kpipe3nyiYqJLbYKoWo2McLNfCgRTi0NTkpbGsdL1k1gj510bf
h+NEMbNig8tcTsRXZrMMK1sGvob6Xzk5bKl8EgN0USLThpMbiFVGqMPQlOJ1oVOy
nN1Ml6etXW2/HDM4E3Zn18AkTP+V6k5Tkv3iJE0wJlevmfh61NjVLbUBgBGSVln7
x3FSgLv53b5dCg0WhZgVQHqFkZAamNajrvFKjC87deo+7lirlp6qmY4atYqTgWv1
kjirovuJqNtgP9kvLFY01TSeUm1oxBv2G86eh3C1VQlJwzPntZfGDwzLrSGgImHW
bjKcsU+ErgGpmJWWSXzZPlKx8okK7Kv26oC4iGRUhp817KYtx8F8XfyOeXwvuV3U
0EvZcOOG7lsipbPWuoztR3utQa695BUVbJZ3dQPDpc7VuPyXoLOY7IEC/Oceh9r9
DcDa0ckQCziKkDoVJ1EbxrjSs3Ufp1TDyMsyf6+BYQSZpEBLMQ4Htsp6V5h08Drb
zcrqb6etAEjQZTO4N5VoecyvNn5PUGL0fxsN61r+ddguqB7BSJSRNzkQcowEB9m1
miDAYhWGt1H4n/9CoJ8he81Yi7FXF2Nr0AXJlUTvFYkEyRopKC6f/zk879DMXS6z
Hm6rGiD1ZYaZUF52K0c5Xpl2uQp55Ed4IDKWzinLNFfRWeqCqfReFHIPrE7E3gg5
02RzX6X8kLwZJNQQ6MRYH3IY7Q4oybRCs31NwWx1ZwgQuriY1fOaKl8mlACKbnFx
dK9GrwvgjqeoZ3yytQceFcwy334doQiUdMAn5kUnlLjhhKt6rVPp8sUm4wxEisjl
cHv2wi/nRr8ySgZe+HDkksJLAuphtWlKyDaCO2qs+5EtE3mtkzmFmswuuFskfgvN
vB1y72LW5RNss/K3L39ISzzvcKK9Rlj5p/TX+tS3v0Yb4HGPb5Gt9KgDqnpRLT3Q
+VN8MSBWstvSNl9VLoZZRbzho4IP58Jf7x62iPYTthpuzIcu2oBG29K0CBKSkI4Q
aL8FVfXSNSFDeQx5yVUq/aySkjiVlI5+G9kfWsB7HVFaodt+k3/gwnDbnydiBnwh
6dxqN3ufwIpg0/74nOzOMqReVgQI8TF1POBJtm/K6TMj9JdtANe/y+T/J2lvefno
6mYKf/v8M7Ob0REGTGxyJ5mbnKoYDu6Wf0psz/64tc1Bd/BleEoP/+cJ9zRnRuwM
0e8mDKjE8JGLgTqqy3Weylle3u4tmiBeiapwL7rDVfG9AklrCXgRJgQwm+PZLfzx
jwGsRPYVg8JvRFKoM+6YqEWFtYtkqFBAQH0yvbFpDjPBQILZ39pjW7dk8nU1NPmh
7Ieu3Lby2Z3AuIesKhgmRUS86hvkGiih6bBMZ2L853F/pju5+7/ovm/nwbp073zQ
PrQKRWvTUp3LggCl8HpgRW8xq2wqf1Ba8xqJ+wAmmpAF7tmDn9rFmXCz2K/2qD9+
x7KOidN4Za+aL9m3m9CIKHjF6PtzGUE1p0J/xOel9BsixTvViY2Fri1+H8nh4Prs
jiUf7UJOclNKn8L18Bj/37BEvwspCfWxPn8oX9Co1NGoYsqYei17fZnvhOUH2uiU
vM70eU+6eS3MsP/H97vxpCadTgg7U2udOmZJOKdEGnStgTjHOXMnccIfX1M7ARia
Wqxr3nmfIM9QrnFDls53spRjdZXnX1mM/cRgzuDzsYmx2dBbRWHD549qK7KAkRCv
a+PdeQ9F+4K93gQy7hJITyT8oduOF8IhNM6kSLNyk/kV96wVfWhNpu7qKpKIf5ON
9ebflnNZdH8Ri+UatO+KJ6aIx+nB36vLqaXYMiZYDsCNFb7YkO94Jik79pMpRlbF
XOJ6L2mdeInIv5GIeu173tYw9imAksaZCI1okakjvkXuc9+GRxZahINVf52BmBkq
4TMCnWtd87lEpHNf/Fc1VpO2LqJ0tsuUFV3MLsMc3qyJwvHQYHKvyzZseX3FWrLW
gEHenx8fHnBs1PNhKdoQEri8ktl8dnY2G8dnT5Olo+blxuWPibtg+VT9wsY+ovD+
m4hCXAfJ/VX6k6FJfirPuVK6dBYU6oauKCWm0f1+owlboFMiaewG+8sL80+2XVuc
F6wRfQkY7iZ0kMlpF7A5YBsIcyizYaOb2WQRvDb2JrHb7bN21TT6Vt+vXlrBRPv8
JHCwSc1ts917WUMn43nInA==
`protect END_PROTECTED
