`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZCeSq4M63O7xz7Po73NVvGz//s0J6vEEmdHWQ366Ox51XTLFjdykU5/WFW2xFbRM
Q5wy2/JFzF4wZ2vHn6etQCV70+2yihGpfA2FyD/0QODgESDmHwsOFcTOyj+BPC/n
7LIIrqK6ku25wDDad8x+wB5IUUGmdpeWDsgX4twaVPUuyOxNkSPUTpaVqURBDH+R
mOVeUxqWGbq2obmmPYonP37CmxXYXqn0iUQ9EZ2hdoCMlLBNpf5VBrEthtQB+WEU
C66+vt+HthXt3NnQVwsjvDaFGW6PnhMa/kywDgpyn3u3luaPylNoEhDYVGiXJkbI
5vadh4qH+8hBExB0HKM5mFnY7BfLyPFh/kJfzBZ6t7wq/t331t64DUHPejI9Q5Nn
+iNKGxAx3LNUDVV9RE8DONgCC9Z37yzY8CsEMN4uVfARFLJKah0cAZAHuurjCr97
cUT4tCVEMmulIX1rlqphjYR5zD5hFCiH37c4QJ8JhR+Z7BmRpmnRw/YH9sC4jFRO
fMw7BLBfZt/QA6tOVwBr/zHYxtd4SONRlJGc9Odtbe5N+CQCupHZOXL+uia2P7KL
VTeBU+/LL1jugkc39RpRTw==
`protect END_PROTECTED
