`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7FPxUzrf+lEkDoDBXd7xmWjLjtSk0AmiqbqkW1gswDStvGrZIgiPw3RUn2T3IWVb
97nIrJruKKfz1R3V84HYxvgSQP/y4byYa4/qCOV0poVJzrLi7d2wmkzsEv9iHvuf
HuS/fGOiTmWaMoOZDRw+WjfqIcLw1Wia+ZM3xgDieor264NJ+n2Y/lEvLsgnCerz
93jT2/wGOQPsEPpW+n8GN1CP7Em+Rhxx1UJ15cfrdAFGS0flji02eH1euDqp17Zm
GOFmGp2Cr9PvOgg5aOj6mpkqtB/39G0aykepFD+YfKjqSGyCJ6/aly3UTm5CTnyj
Lowo8iVaBm5tBSI+4HLgumCF65ukVT3tajvRBMmQ+ciy+w2vOMR6Reap1EF8Hht5
CzEbJfqPBaIm9LkRcMHDcvKhhUFkwPv++fdH/3rgWpli/az0oTj2jNlCgXRWUpmT
TO7qhwqg6wEk2vRlVztrD0hgE5Hj7NvcC5xAavmBcv35vsyUoI69Vr1mxXYA79le
SVJRbTFqk3QtySSCFj9iPIvMPvk2lcBUwy+myrSiHpCPPohKfqrqON6CsYgj5sy8
1oVVKQamjDYp+aB9bAL5knOb6HQWTVeroRFhuwdS3vrqVEbxfzZFPQC4yQxh/Wu1
bi1eOHuwG2BTs+urHIhVXrIkLDK5vMawdMFe+j+bd8xca4xtqxsEI3Jl7UMa3hbu
yAlYT13qAg+2e0BKnGlZLa+XAIxWzqqVpVH20waN0eTo9l4eQ7dIK8I5xKDd6Ezb
H24FepbHTQbU8IuI6JMR59OmQMCpSZR5qShPLzgHFMtW6WjYZwkgHoZ2h80CTxG1
7b64nb3lMDquUQ4bb6EWvMsqn7NEv9qTtJ0tDL/RqRUuCf9xgGFjoeltnNKZkDnW
4HJw2twoo5Reg468IHaB4IwzT2xxHYgtgrmRQDi8iqNOf8xd5N9x1YLkaqwtKuzi
iMWsC9JHlkds6QkEBmFsd/E0pAn8EWdQrrslwpRkw7hL13qfzDND3HGzqaztV0dt
24nc69PH4LG/Ah1uwJFjljIwjFsd1h1XRVt9G/acotsw3hiTmTnoY9MJ3MLM64um
UbMyjwRtlqGvjZNHo+ldnLLAzHFjQZfyUf3VxbVDci+51XHiWJiB8uxwJ00huajc
kociwqQFyAgPCDoMjZ4489tGukml19WavgJwyP2oiTZQ8hxZmZYUAXQ5tXHBHWH2
tp3goke3xT4XTX0kcFku5Si/ujKIKuJhNOTBNiWDFEvKOjOWjvVssfaouTCOKDIy
m13xuYBwAIWycqhy8yyuwcvjByJFPVIM1qhqc6nRnmPn2bUauQiEZBfP9kyu9eH7
eFFjQRBb62mXUmLSvnBdFW3xN4kPFORfWx7fOhS8Opv4e3CelyoHuku9z7lRoY4H
zGcuIRlHJteb7S9RmEww8Xw8Z6mmRjWjwK2Ksxrh92Tgb0a0Bfi6HMg2R+EkoNPI
0R3tpRsEYhuMucbSVeYqoCXb4slJ9EfeSVAYIuv2dfrhFTOAr5/LGdhlRJW0vEBb
RnlKv2+/r3VLx+zjhpNQpe0vmcKTaoQEoE+vVUb1IuiAt3979EfRxUc480t9LR1B
u8NykVfSO4YsdX+eNwcYYefpaxgU5EnUdB7J7o1DsKWhu/8uE/i1hxTjDGx1JUFH
7mDLX/I13w5mVXvOeHhW4mihA46BVQoLxima8Jy6zPi8fk8QJrS1sQLAtthCvM3D
AcTRAvF9zDgAHz1SpE5FNT3LTyoyfF3KiFElAH60pvaOfwnw7za+n5fh/Msiu5Tb
8hLadUeTf0dHaWPYrv0nWuMxMAuA9sVlY+gOoqe97ewWJQTxQAO+REEw8IB2RB9z
Ut26+Zn1XUXdY9zwuE16EbzVRJXN6RJXqm2lmbiZt3o12nj8xgvu8quFANmp81dF
U+YZB+Ij3smHgh4P0j0GoiQw4XItMKpyePSwjWS7tr/UtQfjXjBZCYUovJwtbd8U
sRKHwegCIlYKwElCrOTNZA==
`protect END_PROTECTED
