`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eb5B3K5lfjIaNWKYA7O+/adzG8l2djmVX+BJneor18IYmu+rJI37+tBvVK5zMkwq
SoExkQ3Pv/ZMVtWWas3emQsk7j5UjFtGoj05WXZh8kyc7yTg8Siste9DHPW3o/Fm
RSxFcS7tF1+EwlNtOdCbsFNUEWOKYn8Vwprkl8G2EI/73odDDwxfgNC97ha5HmCY
1ms18DZ/cmfjmFfcYH1XBlj5Z8nBKrp3twxAKIPBBRTcTdzszNDOS8HWBRySSv3U
JJctjHQJG1tZAfi2cN9qPQjZqPUEvyzH7d7FCfjw81kF3de4xemnpSRHg4d/difR
yrFEF7frN7sbcF7APm0M5y9G7PVvXLJvrwpBqPWMnEEzdSmJtGmHJd0Ms25GH7mR
LtiWPF74gDEPu4Eo7FzZMmC4bzlCZ5z4PUUa4N1rGoIGbtFRpf3EQL1s1wH2eGVQ
3SQA0NOGy1k2v5aqF3MUTwM+Bz+kFVXGgRhZNQPVv24WiXwRylpaZHkWsKrgx9pg
vzHWN3w0rRsERzAPej62SdO0EEVG6gUKm0WKPQmirpX7HsAIzSRx0lvflXt/1FDB
G3B4l/c65Lio/I4LokTjZtN2ObX2KCJZ1FqIwRkF0cezSeV21VhRWHiy2Avzzfmq
NN6pA4U1aL2gTz0ZItFNBgr5bWK04VxPirT9cYlvovWJ0OLFxx1ttPoX/tDSM5N/
9PxTc08WWQVjUtEwsk+Pb4kmOfWQFsvU291jwTI1BrB73yqpbuIS76HuhHQ4eMUz
22iGSURX0yvmLBnCf8zTf/YiIXdTVUr0R4BJuiLDy3o1Rjeu7unN4cPdt1hG8p29
7Rp95I/PBEnwpT8nXuIgD4EnuA/baUvW2wVmzLp62mDiV8RHXSdTt/puRwGSu6OA
LqhKsZjD0JGioIkc7SekLRrHsuPFCUbmw0hjnd37zx42vxqNN0U7dV2iSheFcH7c
j63/Jr+HfoPExpqYoj9Dz2284WLsMMhAoYRDPSIZuhbZH0zMLq5xOBtVsstUE2vV
AWu4DMURVdPAd/2foHRyPM+DMmtVngMm4WoljfOO3A+/m2k309prue1ZuU7jjIAN
Y2tDRzf1m2YyzE9E/fD59XIk2sJFVKsFVbS7K1jGpBBBvXoYkFEd0m6HksxuGJ2L
Xlt4w3GFEEQQjaIBxS+hpmzhLyiniz6abL4TOYxAZysM+Jx4zIybQAjRSC48JmA/
X010r4yCLhfNxFu01VSToqxT1o+hH7SwcH4Wr/O+84Z7AQd1+Deu2BGykeK+Lu2a
ffJm2TCs+mvJCngnV9iA0HbJAgywtteH134BwtybKEybRm2DkncdA52Q/saII4R4
YjTsBdxcct3OseZ6irGF4I0Kf26xjH8VFl6pVdpiMvN3ChZ7TTkGs2kMnlSIItlW
2uuqXp5egvaEY+r4ofaNtSnKr6867SZtVm0/K1e1trXSv0aOzS43a/qWOGSPo4OL
gQoC34+9qRq+tT4TRWQPeI7sE9q/yoIo06vdhklSpxxmx3T65EXeK4X/wak20DBm
UogjohPPD26iE5BePrj9lFJaQrEQmMjm6HuF6ja7BU8KcSm4cSnFKBDd07mREHY3
p76t5dnnlwFGZxNU80qJ1BM1IidNPf1gasfnpendSGSmDBsYPy5GyAt5sf9T+Wfx
yKKqlvgLHYcFHam0BUxSazeN7M2CgaMop2CPe92grMY7duJyqlQ/ESgR2Ehpcu0T
LU4FaLgm6Mn/Aky71PXT+32oUnqtmf3EPlJXfhSJHoNW7JgUZ6Zh+clehgGn5L6i
DjqU98eVFKAgCmrAsdYZEKMGBWYi8Jyeor6RJ02AaESPyYm3OpiTHYcTtRh3F5FT
/kZIG0XMa6wnKruo+Pt04RArY8ee+n9dmiW/eapZQAHiwWbHvVtEVpEDTYwS+rpI
ACv7ss5LdFgSDuGfJD9pxLUCSoDzs3zmv7MJ67kUhh6Tsdn5pYMUWrznO8ifBDrQ
5hmOHY1yesQS2jBWfzjkhJZ3GJ+9ZFJ4p9p1cDRaEn5NVuxYCq72B2GHF82k/UYj
l9J1G+2xMndfLgshD1gK9618bjkUJUOp8sAUb3EvgBiAf/rnnimnQdRfQMF+/i6s
bFtx6Sa1KvCusshgk5mR1cJmPTm7Emn3I17bhvsjLezw1DhaeXSPuA9y/lDcniLu
ldL9RHPY6ht3ieUWx/HUSZJ02rs3jUobdL2PArcEB/nBeFmI/K8wlFpG9rg2YwDQ
GxOYYDkf7QO5nGnJEJvzd3h7x55aHCTG9KV3OzNKpuxsouMyT2ca2WNYLTqpPk4I
vAarPeLSFYJIN7jZzp5G+X+bnhGPpl26mfrAzZ8VIl4mXalx0CXXiTzMxLXIwo9I
rud+wiux81QAub21eLhfXTNMC1Ojy7AL0H4G8t5Hmsg2q1jqRks5EzFi+woTLhVi
zYWUCc2m5MWKnYNWP27V7Q8dO28l9EyvdZOkawQ3B19xwC8OZ8NWx85IkVaHJiuA
YDsQfdNnzj8kpAVzvr1OzatiWixiiPYcvYnp/4Eyqu2z6Yh2Xfh84pIfu+Mmb7o5
5ZmgOf3919rvtHvnyPb8U+R6QXBKrey/jX62hpkjojXl4yk66a4mHdD7iT3gx3m7
6lhVUXMcWX3/ghWdynXtiJytB2RwlRhkuwEyy+HVZZY34tPIOtha42lHnF6HhnWT
a4NOtawVynoic7riz5p8B27+3pGDc+nRF4QYDhaW6+f1YvoYu4ae7tDKk9gutdA4
n2mRezSxXYh/qBgDilba5QvY4HYSWlSPkOre3sQGZxImmvw7rXsEMSFdvPmcXPrQ
Ha/6Wksx+BeUXiRjy9hek7k1frTTjkNtrZ/RxhFdxd1YVWbuQPmlJGWwugw3/c5D
4R7A7eHCtyje8YuCuH0THEvitQ9AlUnRvopngmBLAgvvWC4nyw0yP4pqJWVfUX4A
nOjxGyV3+00IBoHHIpYx9pcfv8krsfekFVjNpZI2eH5pyZShaLWc1yJCjVnGfNUs
zMHVHcqWZ+PsU3yVuQBBPUxtwITbOtwOUYTQp+N4QM2Ju8VrZlvN175eXX52uTDK
GVE3Ewcdon4aNtKq+0/lhy7yo3lVWExc2yEItvp43w9u1hWNUFc03fjFiSOhHlR2
dXmlc8vevJxeH/9/lmrA5imr1lvdFYx9FJiIRn7VjAlYXHPHd5VSyDosOQgFSFBt
rvJ1pjOggl8d6Dr9aeY/vDWzMtuI/CxoOTyjmsR722SX5s+Y+2TgPYBzEwwgnBUV
WPiOGCkPAFt8mdRpORl2JraIr3Ict/husyakzc9EjJ9zIrQpptrggy6NIwtoo9hl
76oxQcNDndF/rR3ElsoMETvNSVz8vv6Pw3gvEEIR57hlaNanO8wVIBo4Kgu7frI4
WyE3C1NTgdbp8SzsFa+ftosfo8RV0QhSP14NnlsImL7cSdmx0FvIYyCFlvG1WnRG
Q6LprS2gCdo2/ZQ8jPXaUpSVCz1aPq+aVx5TgzJALN2579lQlnYgZeW0ZacaZdGs
OC8EjFPvdt/QdId34k7jaMZvA6avSWGnSlP092eQUSEHcdgugqTK6Homlcj2kLSp
kFiaUSfQq7SjKef9vIMH8re3nTeNvPqyabeGJfS0YdxB4IL+bA1ZNtuOhc1JroKQ
ejkdR/ba3daupi4z6mzJ/84nYx5kiJ6sjgn4onLEFAuJTfziixJ73yByy9LHFkry
gRS7VLb82O3X7epP9cmVuF1xSDjAqNPSbyjErp83o95dhbjBWzq5Fg++ME0BftsH
9rfByGkl8x/JL3nPPA49VC89bm3N4DtmyiHl9TVnaV+REOd6I2ue3MwrWt8opp9f
Jlt+zJX+OYINHu2GnWn0d00Q+Odp6zsPRgYLSjr7QE9fJr0CcNF7rseFzQvuI3SS
bmhGDJTte/JWIuhMWKKYB50z9XY1kto/NQ6v763mQspa4W0v0mB33BHc3yNoJ24Q
FHEe18m31TxtyTwiANQHWXgAa33vkyGALViBHfwRMaunnMWyuOlUYsWBOrtFpE01
G7PoDjGlYfNqyqbWB53rPjQPgH42gH1sHWyg11GOOyLovWgGFiYXPdBKTG2lK9jT
oHdjF7OnLKx+RsmI5QUcEbLVW4FdtSsQ11rcRWren2W9g+p64F1a5gxuIyQBPOt2
qXdpJI2f122WiMR1oI7M00aREGweSW47fgMhAxwiidfHL9ejTgVxbjyTyLXKE7uJ
WmvpR1FrQQzHSBs2fdwSmqYHsd2+1wY8A4OWfUBPwoMFTAeE3RjjlRXK03A2FlCj
ktv7JHDvZ8mCYshvcyeRW8kBOAhl2mpbcvNB+pft3QJZjEjAq/v+lIxy5V6jLupv
L9yv1QxlhN3nkXfk6FzzXPurwStSPycIYhti9suDike55HjPckpau6Nl+AWqyyCW
DoTpY3hFg85ge1WyCrIgtXPSvtScUwHICP/Di3KGtUuHnIr9xAMPgZAwohSr1IRK
0aIFGWyC1PpIJ0KGufEDk+3dS75Pg0mXusQIa/WIa63tAKwK/0x4ADXxxJc/VSU9
k137yOPuriiAhqi0l/PtQ9MZ0T5C9B+wG+YseT2eIB6EM9Er5L4tI3az2uZ11WFl
cw2bzWYwtiwAReftVbYSzJbq3TtDQE5H/Xpdew4eRgbAMXlcP3uyR8IC+K+TpK02
eVlsD6lO8p6RpjgZ1nPaOrbJVHeiyblMwW+GgGPB8eIKvfgnJ7Il04TBp6V+5xdl
V3OoFqs/ZoR+ipQkpkvY9uSBNlBWqY5gHfBoeUC1bnXfHN2Ar/joTJdnGOY/Tf8g
KxX1u2K0GheyRYZVnjXrDQ/Ttd/+4fSlW9+GH8/lG9VBUx4LgF1YwD86BNaOpvao
/3JH4MQ1f4+/2DGATYeMycuaZC+Tch/t+03xIGkQ2FERojATCmF25F/tDTUtRIDj
uV3zWKxAfU7mV98U9uNBNz8xfx7wmJ5eE2QUEJU+VguJx3n9aG3pUVmoZvNUKtWO
gxEbJ3VYNnF5J729GdXSvkbp/hPvoqEZ+X1j/Fah4zz0GhrQo7G+zkcYj22U7y0U
gfjdSyV4yfZ/E37ONaYDptaSnDXfFNmC348UA7JOHT57re8cnmFLgL1Vq6LwAcj1
nDrfQxzrlLskwNeS+3O8lm0gu26JcK4jmXH/QadApwMB9tqYijLnyRGZeRpcuMDc
bwzJPrlvrdLWQJWNqrp0CS9F/X1C/U+KVMghFx1ITkYAkwqYlmh9NwE+AJTsPJ3S
4j40l0TDWVTR/vx+PTYOla5Cb81ARujMMliket0OBVSFx777fkTWg/TaVMQOUn4D
8Qior3v7EYoGsz5vv5yXKvGUWtfJsS1H5RjMWFeRwRW7bxBBgo7IW93s8zB8TakO
583ejPhAuISpkQ+mqGvbzEJJgP6KMwtWXMtrmHw2m8SSRy2NtR9sjaWuy3dQg1Wz
B5AAfed4F8fEt7at4HLp8a0MKIpOSv9L7FOoBqBGgI5IzinUzPecZ5HpX/0Z5N8w
b/bAs/WSxLtjTELB321e73L46kbLChLKnkrAyp6IaRVsullhPSSPMI0pJpwnDhS+
XyHb9qtiZa3ZL7j06EPfXhhemmM3zCcNLkHsNZaTql+wD2aTWYTGONoIxQKa5nlI
NsPbRW+XeZJP81Y+SFA5/AtS7ZclmDzZ+2DOkXBeuWY6yXm5Q5xVQOPQJFuYu6M6
WfLgDb+HQGucp3oNMQ65RVthscqHVqaZclj+/DPl2Cy2EOfUntj4Dqoznl6LxWmQ
O2bbyVk8mJjtFcvhmv0qk5EK2p/84Ba3oyuFY58wV86kJlo/NDJbdgLv9+ZmYmdW
lv/S9obshHgfL4fCsCuxiEd4n474IbxRcZeCH1My69N7DDRxPOBe59/A+E1crq2d
MRtonx5sJkeCSbCX9lgwnuonb56ICuSSmxwvmuiQU7CqdiGcyRGVQzqcwZtDRcGg
Fe5C07H47ytgDEy/YcdOymByXpKCS+ymBFrovWRFVTSY60mkviJdNJqbG/Iwejsl
6Dmdgi/7kszEXFtOpHrAJWkH8dgpVbSA//q5AnCeEE76PwjRSipU+7TNI/dB+sTu
zRxLNQOj2J6YtvgeXOWRpix5EpS9V4xipzSyYcm96U649D70RaukuZoGMQqxEtQa
OVtsWAtCGsYlM1buMiyVQ0jjnTwPPJW9cQpuEIwtdh/4lbrEn8lYWLT4pwOgYynz
mbVdOfPXdGIDmqdIpriXW6Xw/4HoLiLFe3MKWFq5j7f2TQ5TClUHw+j3bE/R9L4y
AiyUOlwl9oSltbN1HqYC6Nigvp/Qgds8u+3MPa9b134gQVjR3ywAJrQs/RNlR7qH
DuIP7XjRgxO5ViqksSPppnYqDZsggJ4tfq/OW2PauxUi/HBU/lmNSnfHcaeO46mz
HTVKITiGH0BwH7tVIiLN8k98tPFhkEkx+0tbtbDQdUZCWJjdSRef4oli5FJ9R9Ic
mLcXu79N4U/Gx9rtet/KWY11TeMYRTukiRLIc/z7FX8DdFWBCrh21VfjmIRsuWut
KVt3lfMeiw323XM4gjtAr3dwi6QwLHP0IkAjTwLDnqXQvTlhZzYfkswy/z8dW5fE
BMcXxQbM/Z2K37a0lbAMlw66LFYihMt+awlRYSl5EeG+kaECSG9D+2bs1N4/OLMN
H8kI88KeU1B32sdT2iY6etxoFNWbb7g4v7agMTkkIhPPaExlZw/5jslros/nVa27
U1ZNd6LUX6oTTbxrE66hZojyvYrRaRsySMq20HQ0sHm9id7tfqIAN4/mtVayUUMj
nxpsYuQHJsJzsYZ6h3HZlUOvA2j3ld5SL/+cyI5RDGZtEooMyWsEzS4uLtydqDSI
x6napRRoWIUg6XvLqgaTwRximpyNvqnicqmBptquD2wTT+pYXVvY+UyKGIw6gM2I
aHOvZDqy1t7bVbPhPzVdYqEmCXzaqMjUFvjQP038uTcADQz6kXHSQN0Vinbw/4qe
DyoWUrYU5YwFWrPIlKaIl4aF/VUCZ+eaZyampKzLRlLcpwSk7T3UpoEQQ3SJOCBJ
5CxL0xLvfCenW+P+lUWCQuSMTwr+HQNWe04eaqU9bM+aQkkADzRq9hHVIjP9UbkS
BLE7aIkUPtxn/Ia8Ce388tiwktvm8bTKyHVmWi2rNgQkn3WjjmaybLQDpnf5GNpt
KsvxPeZjYBgacMQYCTLWFV53vXdhMKfR+B3Umz+5DiyTQeKm4WgPwXeZZ9jDkBNZ
492koWs5o54/hrZ00ZuwYW5OYx3obIItwdZnkIx3M2u38aMx2q6+vQScL1omfxmj
Z8M5S58n+YSTiiDUd/y+SP+LcaMh2fkBzY9EhhnCuAsAsV9+xUKh4lmZv7zS9hbZ
7VkHq48HNNqaAbZyorb6zPJgzkprbBNNbH0EhnoADjuFkgw6vLnFOiBcg1uBbKCA
Ka0n8291tffYFmvDtP6+cie2uL4RnGSgBA9wkPoVtDS17T0igcNvppLFUJnltBJZ
SRMpkSjsmfiyNfM5/V8CtgskvNYNgJcCpATwfXduwBNO5nedrV4rKVDSirEVtaU4
xuvOBSnsdRYqORbntpTp1aQ0nwHT4nO3aORFZZNOoMPHcYRdOtoc6/ocvIEIv+wF
OsmfokkiN7/5gYojQjCxljN1jp241hAOk+oG3iPAF7ky2HrQh6vkQSEBL0ZmPu4i
21gufwdjq0kALx+cjlb3n0ktkXmO/JVdoixrfB2YmL2vjd8CAPauPaJnciR2e+/A
clFfs6B2ADDE6MnGLO5Nd6ReHcvhs1QXm/WdeMEPfdkiHL+yPt/EJOVdEVA9kIrm
x0xD/fdFiULl+KOyZpEH8CuXiTNTUdNDqNNhKbOcouqvdiY5QvMknbR8fIOxPXDC
kJwJJCBvKE/g1z9dAV4JqJzSDjFB125cwb/mwkw4h7mL25s77/Ejv8oAuOfZftEK
FFBRp1CwWrrjiw5QhMgvOQ8Vdm/DWoGsTGev8lk93ImCSHACvs0Vn0BEtAsToWdz
JRtiqX491zNFEnO8gQF0Z1+f0Eqnqa3IGsCJhr0lJIDLFUkCz/NwRObNSo3lSRz9
LWOBdInr2QKGFzT6Ng5kD6dWj4EhYnmjthXgqUS9Nc/u58hPyQe39onTAecZ1GXY
wnlgN0BwHFvLThoSigbTba3Qz+cF1iqUBv8EoNWGhxocjlVODrUgaaLhm+ZXS7Vu
rY6z5n6t7Ui1N+pkUtJsxmCmRMeMux5v2mIHf3lPTzSuYXfeSP4fZMRHT+Wn1/I9
q9jtwwGeEm/UJcYPCGLRE+yZoctBEcXIXhF+GPbLJrejxWpDgimgK640j31P5qAU
HGZfqQzxXA/qM3CqxYQItSQjV0ZJ2BUheahKKTRCGYb3pQzu0zoAFDTXeHDUehZA
JBhP8tRH9fNBkD7gppxtZ1RwZXQ7qkzW6RgYwfF/LIkZThPJpH7iH4ShedU6cdhV
UXpkoy3A7VvJ/irm4pjs2YLPokHTSOcwbXhknSMFfMA2PofkDdy+Ueu+i265GVXf
+TUTWZB/R+Kwu3JgEMOF1IulJsF+DCGT+RlRU0FfAgI18RgyMSqqnM7ViyYr/YPv
aKaXqXLG81wO0SfdiSorUYvHjzpqw5/H5UwEPUVCxeciH+Su8/MfCNEiqyf2OFwt
3kU2rsMCUQcI2tvetF/b2839m7wMNMEuCDGGyIusls6pNvHHVO04YuMavtP1wSMI
7Eur+YT7WH3p8bss6nzOWgo54otuEfnjgjOIpO15cbYsJ2hdN4nuyXMncBOJ85xO
JEUrKqa977/6JlImsgjwWGv1qLIQ6mDv1pbZWzrY+SiRJ6HwFxlPClC8TK/eU2z2
XQmKbjCy74o6aWTPwIYljEw/mMSloy2WKm+Z8xo18KONM8KC4S2tqvW9yrRnUL9a
n5lnqIsR+YbmRWmYasD02dzCPVNucM9g0h97n6PvEokgaeDaudBNZlHTBGjYiQcw
BGFM5++VWC14QRGJnfZXpv3EX2el2+ybNwfwQNEIIzB16e+ZQIhb9Lb+C8T9IJAU
Gufy9T22iK2Uz0YjMNflOuXwm1nuf+JXa6m2V+fzY/h+nLMvWA20gylZWpwMqN3E
E6QTRiMcAjbfXKvEr5pRK1AxBqBU0n3qQzu66w6VOKmcWR16hfv8nwtKRFc/mSpp
odSsySz/m94EWlJkEeII6CcK+hveWXo+84Q/Nv3AGHymzwHQXAwaWwYKAHTlqo41
9r8HwgD5+wvov9gprl7REK2XhlzR6Rc6TnNm59iPRBvZQXDhDgcdUNTYyI9vxJK+
RLzcEi7cIV/S7zdijzjghEHkNL2SMZKWZZvrCLfVxm7Gw3+HfSW3afel/WmSj4Oo
W6TlEtwxeGyq1IZkQR1bqNq7UxUCj7eVi8lsv5IMKWW3quJf3g6WbW5nEPFu22QO
DuIz6RxS67w2UZUNP9Uzp3AoTsj2p2mcZ/yF6wuwJSHzXl9o5ornqFQsI33TYEV3
AUFj/A+bs9fCBcRYJCLdrLh4fB5/9Dltbhk7LjPmwZt9W/Wwr7lO8cOod50eOK31
OflpaWyJQsPme9kypsgPfLOMTRRSZlx+0CXqW6LoaCdjJBNr/ml3D61cVoLtccqr
jKYmFP1AbFs9fM57p7JG1Yd3NNFPZRynaAyLB9mUGT9v7M9ZzIAA52Z0kQLPwA0A
aGjtI29vK1l0mG7GaV+kEMW26lnNJ8n4m2Rbo/xQcbAXGeyOJWHG1VrVAwfT61BM
EloyZGIws/f9g9e44XjkPt4KQAqKn2rRxrScq+cnAL345dug1dvF6RIJjPb9P2Qn
1N0UBFYjiQSjvK1zEtZkYxfpvw+Hf/ufJUqxS54XhHuoDpPNp4tJytWSir71pJVE
O3ae4vgnTaN6yQwVTvPTItRh6N0s+Fs0/gB82mjT7K5T9xDNv+zN65z0F7oBqp2B
XLBzuFZoQm6n6f+0RFgMQHnWRCicXEhjhPN1pWRHpRH1dMqcbrXCjf91pN36/7gy
aaAKNr3vKbmDMeWBllBaN9P2w/1q8GRpfI9HKoEINpT4iSRF00IH8oKp+5lzpkQM
Z5Dmi8AbYnsyD6G7BZxTVI8Vx6NBCUXCVmHs+CowhTduugPM+4alawElnQwYGwXR
cKQ/ZPMcWwE8p0lgd3eLxSrpRz0RJnKs5UPCUJaIoEbY3e7EeRu7n3pe2GN6RyNt
kaGnQ3LBjtVCBP9IaZ/qLwvl+VNrRI4I3sNSTZ0B6QU782IhFCmv+eMP5yh7LRzI
pYN7BG7YRAT5X9ngiD6pVMG2CALejzEArGcY6lhrqBchm1BxZeyGDaoxfSrf6CsZ
2f6MFRhTiP7BhXrLjP29hPL6uzTQlKrM5lPxt69BG2TaEflPCQoAgoT0WTbpHLe1
FpA+XfmzLsR9I89wYQ8OyHkUuOSt/L2EZ8Rl3kX5fThf9rM2RuTjn4WKXHyfjeFX
ErM2LB9AsCU7wqJ0BaJaaMSpPhACv/8NqrYAVrVHX8sFGKqi227BVfZ4DWBaxUf8
ESB0c54+6Eg82XsX+YJ0opNHWoji5nOGrbk+5gUjiQ1NEK3nBH1A3zkLW2bK59yi
Sw/Dxkx/tfSY3R+mUE2GnAgVFzAA+SXQzldOPwwgsmAdn7fz+e49opE3ioPtsxUW
QUu0WVdTGhXSEHOeqQPv+mUJhW16aDSCZOvIIsOA5obdpsGfWsbWWpXZlhBMjNIA
cvE754YO2hi4zYfQAkLQxT+5f/P/0Hk8bwzFknExskBvLRDFh9HrBijaG06Lvhzx
IfANe06D8NpbIJTLQrwNA4yiAGnDljFvNk3uj1ofibqiWdOzJn8cdMC9SssALGI2
oVUbvOUN/BD1jHPOqoXn4orsd7B2D2BdhQfdjxAveFuRLM2d2n7I261MVYBGMIJ3
ZEeJjwP6NIuMYGpkZJY3qqTAUKM+ht3wj40ud9/oaaslTdRyiXUQmdzZNvCCoIhH
By+/VXl7lhu4EMPUP4SxM77Y5y/34HfV2zXDZawwvE6tP0vUligE+nT/aNe6dPwX
yVUQxZjrMIDFVFbeuHqTbCY8De8RY0HyMr1vU/kMAa2sSBktizHV+B2Vl88SagAr
USE3KNHwtLjh+C9lanKLS62q9lRptNF6HCw4tRs1IPWLlSM8Qme7UTA20UqUMgqQ
C9ZppQ1tTZUS+0kdXw0+ajdek99x2liu6HyodGVVj+W7KWx17L6nZOyE/QbO97u9
rnklWKusd7IxCC0aKlR5tsVK/SNwVBenX8fsuv0EOXMXKiBU/JirVYXkBunUn3jL
aT6L25IeDX7sZwuMLar3/M23MBZShOxLgp9C0vtY8z4lx6ZPgm3EM4N8FmDhhbUH
QwWbWcdjaWG9ZNyz6svBmxCpb8GJSXruHzQTeORUGwdEMOPt8LRlbHawSIgA8PO2
fI0sQaMm5WR9X23rdFHjw122Bcew23WFnPteXazZ6riW8ys6jgrkNZlRmE5Jnbbk
CVnA0mnOBgclmKgoN+yNkg+2pQsXZZMlP07kGpPHSbsUZWKT12xD7uz3dr8lcoRl
MtN8Lzs6dTJcleYcboFLFpVX/v5pz/5YfUCTKuBYInHi/d44ApxHILVAFHJGRK9h
8W3dI3gG9lsWI10Z2u/QLzTGHfpjCREe3lHQqjF06DNpJ1TDs5xE1cpQGuJGroWU
ReX1TT5csXigQnKAPM2d1a19/6KkEOeT49y7sqlyCYcrjy8NA7zEcDEYLTmN9u1t
sFoMiK1TYj2GJUuCqOMz1gfn0e5Yr+4lna+/7GtGaiokpI6vuCa/cW3Dhn0a3z58
C6pix5FRlN13tb+C1Xdo82j54/zNhFIKl6S5W0f7G3Aeg8Q1VTkmenL8kMhuROT8
i+08qDJf4RLHlFyOvt6eEIZ4XNzp2OQIwviueRKvMb6gkNIhw7ymA6RgxCjTi8TN
iV/mn+vyVrcb8YLWqFK0VVDsfFaLblDDhGhryvX6bJUVODfgpixibIQN3yhAvkJd
w3naqtq7eWTkqHPtIC2wSgt3oqDoFKp00nzrDpeKdCvPg2UJd55qZ+GBq3di1Trq
uEZdp8N316K6yWWek6fkwHyrbBBP27nBQC0oV89p9IQFBiN53FDn5IG4H16nFAvr
FYBfhvUP7CUGkOkBfk1/fNtzTimvzF06msVYfBzKjA3JirrdagI/YAv8uwgNHnMF
N3uBYgW2JZp930Kfm/Vs/3F2CjJPaT7Ml4Yg1eTluB1FDFr1paL0GY2YjfMuuld5
qH4dl/Ri9dYsbhck8zOx1AtdOPyy8eK6UIPUelfgNozqBtma6/w+Ujb1K0yhOw3p
lob7UBrBoJKqo0TVdlZDAdt+ZYJMFIL+nb648stL+Y6/hTPZTvKKhPlITWD6d8ze
DrfL5w6DgGfzXc8CigI/jG5cTit+xniDDonk3R/wmLp/7Q92ZH7nTs9qlQ0YMtlb
zi9qd24lHba2QQIa0xA6xzRuBg9UZ/19uxFbIT7I3KGh6d9mGCxjM8DeEFlOMKSB
da1DehR/aJXzgC9gpDU2MgA1ARXUbEocFTC7s07lT+Xyd2ZU6jz80LVT0linWsYU
+fnufZGZOp/KAq/L9ZOQ/9+Hp49XgQrs0DKpKRi/j36N1hQlCktgRbgYpCUo3OjP
KgafMv02F8IceJyfO0BG0Az9qAMQwmIWy0SKk3rVe1qkYA+dmv0Zk22EnIE6JKwt
vwsgNQhvXWpXrOQ5+7jeoPxLpNNMQt/VjShu1AjRdeJMint9JQUgau6hOlTLzTQU
rlEzEJ3O7g2w5GPSw0Eld36yjIw4ZS80zoXuUDIyDjKVFhZUVL3xziVMhe5aEpWk
6FUm/4n9fE5VUbGpeYeIyuNW++oy/SIRv3n6scvTzDfgXG2ZJOU6wG7OzNDyvQhp
LjeHI1i6pVerBmM2ssQbZ5B77I9FHFfBQ1x5oDvljxzVJKHS6klkv/11HYgNPFik
FGM96OexCPp8fhhNeGbarsFJGVJt+lCYrk5P3NB9ab3g2JIxWXZ2p3v64gTj1tyX
fRR1EDXMVzlER7GwXsrG5JiP858g4wxzPYxKPDX0T7hkyRx6y7VFyw2lWx3Orwd7
6DVT8TMOz/+yxuMBzkoOiovRJ+IkJJKhZvbZY4iF0NRDDUkZKvYZn7XFrwHzEzTF
xG2jHGB6Lv9bt0F6xva2O+QV9m1Uf5JVAxYN4WkUJWzUjms7wvDF49mXWxXVH/T3
piQA4X8mUQyVRKDkg3t/XYfDSr7BsQTYfctlWvyzV1ERMxtDeKVH9G763IsqgPVy
ILy5BNZWLO5ezPdvZU20wasqzvdfQ9sgsJQIQrX/v6LRvDDBJvXzj0BQ+707HFV7
YUGcnjsOBPszuc9r2AniifinUzrkPfgp+MbmvEOhpLKYDJcqUG3U+z7K08JmHRDa
CygUssG9FAswWBnw3gQL0qy0aJrs5VdaxXhbms0y545AI+slJ5Jl1c/6K9/Ry+aj
tOdWB6gyW4MbYy9PrPQ/e8+qIlwaTf0nyooClkFbjEcsSPQrJBao8f0MBUnqkMui
5gcrEdFJximRXrXOFsBjdekn0VlZyBDKFoOaWsOOxoM8inbbl90V5rRe/RWcEqEz
gEcDyL+MLxKFp6wlVLYeiRjKuekw8vomvVIb1+iGsS29CLlCI7hlqidZq+Poo1NA
mNIs9jl2LlGsilb0EqUMprTOK6aw4skujdJ964IauNIEICmlo6bkL69jOwS5pVND
p3pXlTVeQVSORf3Vw/dRRfe4wwr4BR9PF8fJS9gX1HQxCjiK2qAzEP6fT1lKY2r8
CnzariMgYOOkuS+mR4lQnJ3uGkoaMHwucf2j+E6w+AWCGsuY43IBGSu3VF518QJw
R7JvMWnkmCnXcgEBLftpMG1KNSCo+sdgkREcbpyNC00wrsNTt0VkYmhFfWckbZ4e
lVq0a2jizL5AogCLrqoh4EtvYr59ku7rHkKsG+zRn83IYwee92h2mfGSHfQx0BEN
508CySBVgFtY6IRtcaLeIAov12ExE+MHRS99qloio64cKCAgSKULVYuxGy/0Zhah
gixKmLQpM5UAMOqBMNLfVY2kTylymicAQkRTJyrznR8BMiONguNsL0dL3VT0p0Zo
Md2vKSQyOXMsOqux8HMz0nFXQxVJi4c9Cn9cITQ86ib7EotK+36lFZ7w8ost7Ki5
jWK03gImd4qP0FLeFl+/b5GgGpBv/LkULVsA3HeE4QGb/v9651NKvpWuvXqFRTDP
Lsi80lIiZBdZcWf0PcsxjyFPhRq0bP514ZU4RjA42fHotl5hztXu8gOT+YvBWzbp
H6foHmSRuDCNOosdxmYS+BUsRNuz5ZjlvC9DlzzHm2xxuBIo/9NuLO8X8YRvaSeW
0rz1wrPWrOlOyrImbPyckSF0r/UM6SbqJji7stPj+10UNvcXcwJ5E1LS9XG8d90M
Gke3jIuk8e8Ff0xafbxjpPVGVhpsTbsYE9NMtRxSyXv+hJEb/vOGidGWAwPmMZuv
a2rqYitL7mf0/rFbhaAJM8MPgKZl2KhPLMFdGMKhkdO622sDcEx/Qd2sfJAtmG5r
9XnztjVwQyxmXBUY3ziaKoRbyJH1PUMQ8hgtRtH96gtsQsZRzNhf3rD1JGwrF9+1
dUMhjoabIKz6GmWfWS+Sz8coiBXq85prVpc6tuzXvUsvNrpVsAXS3Rn+tcel9xZ2
w4LfjS1LmrjCx0GEKlSRcDuNYDvMTjFrzXwT9JoynfH9dXmnMEPbvy5M9vveGtR7
9Qvy+gP5DDRXIsE7AeRreB34du4Tu7qL87B3zRvQ+4PVeThhzbSPCPG6pgY2TOxy
CG3qkRcQ9OFBcfHxdiXfnkjBkcO3lucKgZOCfkoUMpJA+tA8aczA2dDHdO1hPcDQ
gtd9tHJHedtKOztx7ogglHYKYK71z3jasUyVlz1mSWNWgJ5oHfUJgO1m3FycPf4A
lbaCMViL6Y7+ZxOqKb5cLJ13duAUmMalnc1Jw/vs1zcfCOZ/ZcpIB6Lw6WVY3Ozj
zbq+6Qc59wSeBlAp/bf6OTp7V3eFjmHkBkEcQl06V7NDNj/nMLjOTTH5GAbmjvqk
iuec/PDogcOMS5QjqHQJMS1GkaJbyZmsI9JBz9qJjgjK8HX9B89F5TwiDqMWo/CT
05m4AuZmcBMp6WRFQ17nuTaRBk8u/5KMtP65YejM++uasQg8zdsMoUQGbuiHiVqk
t/gZbMQhisbfwEm2hm7t7FA2lr85XbNv6MM2I/yc04LU57zaR79NEoMvf7lGzFGw
oX+XEoYzY5oJsAEqo2OObiSSSoAnIIJmS64WP5JCJw4AfRvOnxnztEK8cZAmOEt1
x4rDxYcV/9A7hBwIUi0cGmT3Hm9a4kr7SkAs4mT7WKmileIzazeO16Zx3WfujaKv
TK6T3cjVJzyLjzxj+84cwHYzTDbc2ec2yAWisORKc49KyyhNAWxRPZDNpL53Pn3C
PaZfEdsaTQelRRsODYxPUhC9we7i4w72v0/UDK3BWN5JpiGN1/BgEE2iCujOyAHu
D5IVcQoSynkbAuJk5+iIgT2DopfFgG8BliUPlW3+wmN5U+Zz2dY+5JT8OdPBhRCA
bM2syZcD3LfO+Mwtyvh0GSx0Nyv64NYi2lMIa6/LVQxOuDQD+k9ZLNJSErwCWUs6
CRlOQdgL0dut50eo/ksMzIzCrDRCT7xGRT4z+FqNM6skPTOXrBpm8dIuLrIDRZLv
CkhYE3HRdl6fnNMMp8+bO/TM3G8T8F2Kqf/d7Ycyq3d3jQdc1sw5gi7eaY9AWoQ9
oH0Pb60Z5KdAyWeqDG6qYx4OxRC5mjeal75LXgJW5YtvD8iuSt/e3UTCtXLjxhpb
kUreOaZH1pUwrY7qLsKOhYK1bpktFWW3yaqDCMgP+t/lGlYgizXSy5tsglKvsJdH
CHjRFYconMgl8YKpO13Xwn7L2wvV4GbEsQo5ZmEfs/ryCElgkcJCl2zWk86YWrR0
pyT444nXXxZvcxGkhk2neArD4asDWcztnbf3vvbcBenunPOAIRAWC4TdrLpVxwlT
HJ2CuneAGljnqx9Xj1se6AwZDXxHw2YqhV7L8gPCo51w+Q9bm3UYSayMh+WoVCzJ
FNt59rGKzYjsiDPaGHgLL50llFJhTJ0veuR0MUtTzu5d6UPXmMJzRIU6Pfd4KneF
14wVZrd/orQpfuZY/NsbZwBYWOzNx0l//B3RRvUkLOifGoRHYp7vWzDgPImWu2+U
FUBpljVhOTnUwB0JMMZHHbsasu0oakllBoWKchcWkbivaL7tN0aXLThwVNQEhZBW
Yo1jNNm1dVAlwN95UNTZ8Q6Z46MjpZwtpQqSqUQB1Jhsr64IF3SlvLp8lQBdzk8s
mONyEhKOb/UOgs8uFdr8IKTgU1dOFU1bcvQMCIUshglTn8Gp6+s0CLqIcB+aUv8e
hov3YbFwFL3OMH54m+z9H6eW9sHbNOZbdXDKvBfeHWDZZQzppweFW7U4tNKzY+h8
zYC2+CNUAQ3kim87Mz0bURdaSfYFTzFxxHWuCFtEhXYQG2y7WhaYcjFFjeJ/Fxn2
+B4gy9ZInyAyBCmCNUVH0EShfuCqQb+ZmvARoMrqWgqp1fIWcr8PQDIl3oxo+/GJ
g0M0UUWxJFRTJW9fJ8GhQPNwRlSDvKNdRc0d9brxLnJrKfl+5GK4SgzbyEFkMsuK
+C+YhXPs6TvUhY7ej+Bth07+XG80uEXJQZstGJA1jg/VOIdbjjQBGJxw+iMcxXVG
jiL1q2jhmPJ8VuDlT2PAWJZeFvthL9lRy3f0t/oRhSTMluXln6pSrrrKZ9tcRoi9
H5DYcFYP5wYJ+mZwW90YssRHt4P7WsgYsQFTrKJFTX2kM7D/KIBh79aPJ4DuNIlP
efXJWQ5fJ5h6nSEz4JkZNROk70NNBTFJYCftZpzZFWkMvnUHHcFQ1fzf883Zk89S
s4Dj6+7vGZKp225CgXVQNOpko3Gu0hhs8OWzEfj5bQ3qsmLHYJtaoCmo25MuJ3h8
YaIfC6q9U1GAH1cnLL+yq9sVlFSZWu9M7g3OtBMzZjp7d5EaavWmaUhA+X9NhvsW
r/9vIrSl4AAnaDxMgj+lCW4qaPMIERDLv9HAPIGE59AKJlUN4j4C+pCQG5LbDvC8
NVe30oCXMdMMyr4h7G0IPttWhPqD52eMWY/IYilw0V91EaNUBeMqgfYNa+wf2FOl
2j0Tb5oGjux33h9Q+wNTxNRQQ0Wekp77lImOdohjNQwN0S33taEC0h5oPixxY0p9
vI6v3R2adWgBckxrQdeQjjtiomyO2LIVIK4256yGGGWWo6chcuRUcfYCN1JTF060
mbOOXHBz7o1NttW6Z1wCibto+wevdQpFuC3HEIXVdARUQAwVOu2+MyaSw1P3voZr
UTT2QnW/H/5QcYFYSrLKk9IyfofRihMljsn/WbL+mBLu8ihp+E61WvoRnko8jCZX
+lyAJhQpNu5ikSrGJt3WTBvpKG0g6++xcJMU0dpnxQmO6CLyhuBqRCSiNZPgh4Rc
WTPQQJSjeaJccFLahRo5JFYtNLtTnLxZDaKQJPONUQ5zXreBbtXOeF+lChoid7Tj
kIhE15QYgZv0qQMeUgROCFLhdWfoG12Ke2j/5ILAEr3rSlFMRs0Cuh2FSqpqQMPl
HuGnrGWDHAO6AqqcG57IjqynZS/nNrYZwl1b30rY9a/BeBAf6NRH8TqjcYc+Hifv
vqRM0ZEqczvAi0xbSbUdN9U7qVNyuk2yInmeoJv1/nfENi4IGTaXPXlXj7xYbunf
ucBr2mpAB3/ciiUqXMvE6WO85d3W7FUq2TaIItRsxe3Cl+2YfXp9dGPKIgRLhF3d
e28yEL3oqFk6GM7CRJayHPcGaobFYNvMxzeqUVRi6mx9Ye9GTX0fGgC/ZFEQXLfP
i5ggC4WYPZ5klQTRSoJ6XfWon0YIjby6f20cW0I01aqTcIuC2rcONzZqLIH65JXa
LfQbIngHw0MRcazeCZp1ZjO0dhvzg55KUfhuNY29HV7pdg1cTZmOipKRb5wJIuax
333OCZJzoWruM7/uh2Z2BiAmRd0poYF1tj2PC8veBjH0JPEspCNBu9svtQVsaq4u
Xn63ISJqNZdJ2TYLuhg851/QZWvtDGXFsZJbu0XqmxVHQLGXnR3TfGx0gD5oBkLw
O83sPneHts9GH/VG47i1KEKd19AylLwNbd5AZf0pU4tMbfXZpWW0Jxnz6FV4RhbL
aT/v85JK4Vc6xg+d5cUxqYWg+dYDtFGgCgcdwq+apNNPPBsf+RD0Q/1Bxww7LSg7
Um5hIrM1FM2OBHI8tQH6+VrEdK+KxysSG+jlKm8DiOZa9Pi9Mn+zclJHH8yEFiq3
S6ClcgWVAwhrPdX9SNMOb70relbwM/cfXh4DXnRMQ7NWEFFCROFdV0DYXi/y7MzB
6ypPR0rWDYXsranJUCwCNy9/TQ5y1EvWAooBe0vzJcIMxZSu9iEbWuO2F5i+F1yo
CJaZsVvzj8HG9bvK4HvIHNyQhJlpAsi2zCrXQtBofejbno1AGFTjeS4p9mD9mcxA
0x3Tp/DMnyaVU+yLvdWgCQl2jmT7UHo3qnioDmk3waFdz/T3kDGRX/x5FiNEuuSd
Wm2PGM59o277nZKjJyqunLmVXaJ2d6jpaGzCkAGeXxCShvMdaUjQtoeZBXt+HPLE
3HXukv9SFmDywHiwAJB8LRQlVd9rx01nEQd1aJWwe2EgJW+B9qtloSnQKcOqDYiH
14kkGMfC/NX/xURg8aUrWtKUJrJLvb4CfgYbGN4zd96MFIZHUHDqaPatS+o3LpgE
NC3Kr8oVkNtBoCh0zwCXRIOb8dnRvwZtxYoJsuRTP2628qaPIY4sbfDQ4q7WnDuQ
PPcN0kkanTQfKNE/Bwh/HNjH/km72nJC7DL76MXPd0eMSdE7A9CLb5qRHeburuZd
wrnTUej0jd96eF+k5fZ4kn75w5evgYnR6BOfjJ8EyQ1czdp/QjWzfagd96S80BHx
UOtd58SzEaqSH2/5Hn5xxPVTfkljuBbgsu8U1B90MvJFVu/QtLZ97K6uUCiBMBCn
ArjSL8AiQpdrl8dL31L79Pcq3PmoChh9bh7efQ+XmX91C7WILYV0b6znYH9JIVLb
d1Zr/J2uUXzJxu9+yWXkw7Ow+WlRd8/KCh3Xjry/VV4AIiyHUxdvChT1kphwAb1i
6DuiFHJIYfyrS1qk2RFZaegZYgt0YHEWddty1iY5N6SsF9uSST9p0voki3EduU2u
VH0QOjdOVtwkUiKP7bzdH1FtVMoaKiUluR76vDsZk+R5tDu+w5xc4ldLIWXqw5Kb
gsEylXu6kg7ZROVuBIANR71H8d7/tdllndGeBw2qgv4VsdV+msXsePNd8zjk2W+5
7uD0KCIaGfZhhIfiMecipVY+RP6fUl+b3F5ytJikR4sPBIYU9uJZ+cm7SpQ3B0RG
ffgL51QWGTHo01+afC2k3MRgwb1i1lAULxfH0VNm+L8edCiZbsyHj3xZ6l7PAxZ2
3L+48RCS16O2+JLSWV8ixnraNAMk/HjWnzJME1bAYcKqlNHwaheLV91Cr7R5/75u
WgnGOihMTp81mb7kLnV0qrhRK/bY8ey1AU9mq4SDNGBGL87PAiYK3hPFuY9cYXcR
ojxwPO7p1vP843vBwyUTxfshiHEYcc3frAQSE6D+bKg7TPAO7wdcLJUt8dRoBUzx
Ca52bs5g0TbLRlZu+nVOK2cTIoB7mjVYaQ5KTNThWTV26K/pp4V4M4YQYJqSnQnl
owvCWUNR7XuIhBLS4FfPKFmudUezSDu5CQhfLwTgVQd5+Lt4BYX7TwmXUCDBSn9w
2nvLmFNA+RO/0yApf1g9RawTsBZZ7PirWj9U0RS2+0vqYM+G8Ino+cmVNU5XzlNr
vVU94W9Pers2vxC4PjZeejZ/q/Ld/cjV8+7G4dOFJJbP3szQqbpDrRmB2mncQvs1
ODFsDN7woHVI+5ROInSm5ymLVst9Wf7/9ZK/WRcuMiWf4V/Bavcv/RHHgOEs8aiS
JC5MmKANNoWylH9LulS8YtGsWlOq/ZweUUyyp7hz0DpBNYE067pspNvh+q9iLJQN
Jr8VaRsYdduAXX5gs0wseqL3psFFKDcdysPEFoESKci0Hs40BFwWgl+TVu+P7TTh
TrrSsp7NhJ0/fJ89ZRxGkwi/z0IWSsULa2AfM5n5LL2qBfv9+fquK5rvZyiCjrfG
EhjVtIJLbve1di5KzSVrzFrK7gqYYtdc7TOAhYHoL4eMLYZ64KyD4IRMY6aNidDP
uS7k/6RGFPGLbNgLfyPrY0WnZuM8L/3E0cGW+bP6U0LAvGv9ourcOqm5No7K9MCS
iY6jf+uFdKNkgpNjmBQHyrcdL0jmXYWfmtEmX7vKSsLNqlmPHL66yhIUxmN/qVSZ
ufQWIkJ+tDfsXbBUNo1lLu3ySGX3hExwDB4MAOJwgKLR5nCEHDFBZsVRuvSaU4dO
jtkr4L70hoL5dTwrUmMO4qgJm6tpp8hOYflwrwZVVixsnh3eHgIuW/J4ypoUw7ZJ
cY+B4F9Mtnz7tCAb6JKuEi3rmpv+LFPt5krbGTrjmcYCVC3LALbd9NYlTGUkrqc9
Eu4SorPShEbOkPwv/DmTOqbK7WvT8AywCL08svlkprYoWzDqQPVUk1whcNNFg/j8
XRAtgRsvrR2dvVgCCzd7+12Qf4tJExSOZokZ4xNlKvuGBy90PjMHLqHvSTV1109B
DdAWgdn6UXNLmqWDAGQ9twpB6aF6wDQBKiJWZJgHNp5CdPKa636zzy2MQxelFuZV
OzfjKy3CILk8jMp5eyjpl0eyawrLUTM/CcrBstOnkPhAVGvBYrMuXP0sV7OczfEx
RRknuSPC338Ve5Gj1F8p5Rg++ixwuIwVWFmHEVyOhE42/9GvgLXTFzelRQ07PZ9P
4atHV7RQq7XDjproRGjDGOjSZeSBhCdc2m+f8lb1Hwn5d2GfCon2mccKaLUPplsZ
QSvssGvsrEED10w13f6hprcLkGpkgAg5mf8g5nInHy16ELyVPQtUnBJh69+8Acu3
r6gMHwQ82HT5YvjM6gfDOuGcMFLr3N5QO4rSeH9Ff5aveUDa0NQ4JKpHLhsfZZBm
25v6daApBghCclnHxoEOMdBZ9qz83oJXnJ5q2JM6QJHeTHOu+Sfp0X4gzBeAyHHS
cb242NIMyc1Qb0uTEy5RqYhGS3kkXUD7HntBCTv5ylB7vPPflexuGcRXf0pYqTXa
1SAQHCJoU+JDtWCS5+HCsz7jxFx2/SU8c+KraVYOZMNSxyE15hYcoyV7OlsZrwT9
jyWUd1wNdQuJAoWf7e/yvbmLAhePZF88bVMNh8bUl0ys9xfcLT+xnpc6zuviJr05
DB0fscxCELxj3Bz9uDw6i2fjGHx2bIQolMnKdq1I6j4BAm2XZVPhr7EIme2QwT5j
kn6a/idXhZAcFBkejEwkEdmvnOiF8RzkGVHo5tL2tw/s3HSMHUXtsDzRbhFx3LFo
oFGSyuA2XI3T37yeuwmPMUHxUT1ODA6Z0FWYyoivrlSFoEaEQNauqxp/r9lXLZQG
QaRXVbGqCFUkRsrAx3vTs0bwj9GBxklcErUYWbCDmOkg5MFBAjjSCKA0CCti6M1B
Zq3qwjtHFxg27GZ5HEpnZw/6VyqLQFUXPJAr5/0sFjwO3vi9PLhcUQ07kYF9ScCm
u6pLUua0GBgyX+6VBkiSlfwvkoosgbXLj+BLoKe2dFwGa6hocj6Y9XWAfuPrMIzv
GftoLigevgBrRVOCG9sxsmHNoH1yJAYE5HFvKb5JYQcewGJ62jAlIMIqyGR+T48X
7tJnx7gkKF6nacvC+8zn5ipoZsEVXyOtWtB336gtF2oia3777G9arZOLGjeuBTSw
3aQhe1fzHrqjeizesUKMlBilvqSgssMBv+Ettrm2IsulalfBhzH74F08wl0aE4C1
HjQa2g1ib++6H902rVB7fWK+WZ0iKDlT0nycSeO9i7QzE3Fc/weQgX4cZk5XFMrH
No2hbzeAH+L3uaiS4N4qZGtYhFuWNDgv/Ft3f5z2r4apY1X5GCIuWM/plnmocCbS
8H09lghohxTAyyIfosxZGuz0mcrcFEqY1xXM4QNfz8qDw4D5gGT8YRL0S3yzvfBi
9eNY4nTlGE9b9CYZshWMwIZw7r1qYdjtm940poENcjCtEopBxSbdKcJpm2W+I+Gg
wGUuwAc3wacMPqBfwNCxgEHQcrYMgXcbmHSIe0p2kmFBzmFq6oaHuu3aMOxAeaT/
t8z49WNIQqkhWWeiFbufi8NnSK1V2x02ZDmirZlweHG25XXaLw2fCX4CGy2U2HFb
4bTnE4ek/fn0XAa9kmkcjGZ7BKNCdRtlZ91inmqzKH2btopvlVNRqmBT9zT42kID
Ql3sdMGbc8rNylcrQyljgmkAqsrHrtODC0ajCTpmaVY9a+Xl7Ht3AT9J5PhnYQwP
JsthoGcaQiOXtQxsKW6OidLF9TPF7rUB/ZY02+URVZXNakS9Vu0q9nwUv8ZjacE9
IoQeQr/51mJEkUHbgiiR16PydVCYPlCzA48IsRN/mhJQEiEUP1+DupvQsDaSeHnw
frww7WS4Ba7iOIFAV3rv1zgCYZrZH7ypfVBPSdkpD2s3aS1aIdkpxBWkn+ewei9d
fUlLLW4/oSnhk8VsiVj8nSB7oEnZoWVj3UvR7QYJjvKi/txz2L5SAcPC8EcqBGfZ
F8jhxZc73brhNYDxc3QTbWDN8tFNv3VEJEIElGM75d/SguBf/t3TV9NJ/3TRVkCt
iNXrvwPzWNB6cZXS0lslEDhbRvaHJDWQBxAI3UzDDe1jWcN9ZQheJNoEiQY6J0Hy
OJJXPTGpfmNIs4nSYgXEW7m8aDwd3YVGz0cQVOAn82B00CwBqI5SRGI1MkGGJjux
kL/VyiGGtZRQbcgDOy7jLHky0Bp0I+1miHbVbdTJzbRZ83jEI9lXwv9hPmpw/96T
sM85JeniSbu8svgJnpiLKEfTh77aWNL+hYkKdoXl0ZwgRMyYRNALYBmmwQxar9Gm
2Nz3L3FUamN4VxOHOje7IRgTp/+7QA2VECy+PLrDNHptJe+2yCHV2DDiFsU4rklv
HB0lM4ZXQOHzOKzmTUo9g0fWH3MeshEPyKGqPcQ476lRhUkbGCABcpgjzHJfHWtW
5n7mpKiBU5pWr6Wrg7xKEwX9gAjCeTN2boLk6rO0DfBp2qREJypmPoAJYZWbAaaa
MdZmsei2YoJ7wjqbswPBtvFQqN5idS/Ynpsebos27akBKq5803CctyGGGSySNVn7
/F+Ql6xgow303yG48vxVjnbPr7xyiI+TmVAp3f+Y1KQPb/wSV3JeEEfxNtp5Yseu
stCZOS6Lc6EtfLQ94zxeWZAQ/TMuGd5VhFGd8J/xj9/lmaHN01VdDSRFKfMd/hjT
NoCp9pJ0+7LJrJfFoDKUWykUsySjEXz6LY3wvD5FO2UxPi3IKVlpIqIcqsrJVRbP
q5zBfu+hgwpfgu9Fb9PpYstXMPqBzrIhJWwbalEQkoIDQNFj38RlndKMa0zFChrp
By7asXRNH3p6xVZ61YjeRY+6wTcNK+Pz6oNE8f/6gvyCM+InLkrQSP9ZfomMX1Q6
TXgr+tmwcPH8w4/kdl7N8Fr2VcucwZ+2+zY/XegOnwZS0BWbmOUdtlSsXeD8ry1Y
gsOGKXKq+BrX3F/b0oSJrImx/PYbBellp+ysyY8Owva2ccR9NyxjQVPxoqMoAEwF
FyL66JV9IqGNyPfNVB1uSdE5SAIOWVsmktbgIy7e7+i9PLEf8y8v9P8lLULEEHtE
Jx8S+g9R8LXuo3Kj/q8Ytq0hdPazD3GRnSebMdi1Dfj9y2B4zHwnkqU8Rq1BSPz0
xN+eiWwYDQ76NAYx+waAPrmtR3UHW7Ae+hdxMJVT1Eb7pSbsXpRmGFGmVp0hbS/A
5Fn9rfBm6Zo5G2WlmsHyZOZs0rtTmby82AnqxL9ybhPJ5E2/AedyaVBJBC9ceU67
GYGhsGS2JIThrkGHknafeQxyeDvzMwCMpYDQFtMfwJawuPeH79RgKJ7XUx9dmjF9
EWZ4osfoLW1/A0dVb8qWwHjT65TeGPW4AbhE56fuUenF7PkQN2YPIp4EWH4pnabq
c7jJbXPQeumhHhknQJCdhv34ONX2FMqHk6RVleWrpoXy3pzObqVAk7sEwwdfq1Xe
Wc2MC+hlBvyKShEcLdE86MbAorKD079T5Jj8vfQfyRlSiv4ejMokwtFXTjqmeDeD
mzhO/agSBmZ7RQqbvmbOmIUnN11lM3mJtYcQ95t4cE2fSSLuoh2FKzeLJjAXhPek
nrAxekn5LCoNAuy4j2KpqT10rZKEcvbkZm1ldq0lBXQArFwcgvR+QuthieRPuNBS
FZLJzrbOmaCcFInkrTi9fCrGXr5F5CFjQJdB7utjqPFUrC099kYP5fAGv0wgBi+D
Oc7wtYkHGlUPxrDr41ETVWoPShjbml++5ztsSS7WZbshCjrFk6uw+KADT+phR8LH
vGH3Rcp1HEyZgWKsN0I6FEpuotESXy0vbab94axCq/1SqIPNlBv08enOqbeIdhj0
14vtMJ98Khssko/2EhXhDc796siDyI1aYFOAFbqikzO8Fp1jPX0E4mzl09dYma52
0j2AASEnswUtejTvlvD7wIz8whOZhECTPIlCS7SgbLmLnW+y6QuTaWPLE5J5RTqO
kTCjhoEkXdOBeDHEm6G/DYQBlQZ7OmMuiBTEn7bK38sK4UPXSVDarLfyoXkjYzfB
xMKMWJU+njlTO9Iln0w6D8rGvizqHtIkxuezPu+3SZXu8AK6v7ImtyvfkyG9emoR
cVRtmZdBgMe4hnh3coXl0Vxgn+YrV0DFgkVYymrEAQiimFCRkR9tsGmmCledt3K8
nIDiarAWcsQ3Qc1l7Mf357REYRJnnBnJ/dPb4Dg2x2W5pkmGqLb+7MU3nJOBq0/G
q863hsyNT2UVKIrU5FPCUOPLuWWv/68m+34k+1hRQlYQQSNBI7RBwUumUcnmasR/
PNfn+EzfJLP7b7Fw6UGuO8rYlN6LdEjeH6GYl0ysZQ7q01UW8Q18aCJPpGOIZS5T
Tp9T+XGTs34B2bkPw948jGdPUPcT3THopk23eJH9iD/puuwLyEDwlHEw0NA70ASE
taxhtkl+bXZnSSkPQZC+vg2gmL0xQVovARi23RxVLRWwND4BPm/C/cK38YDfMsuz
uLrWpZGcgXi07s9cSTOdQg7/V45cyRTgkeoUvUjrMFXufjlJjfprT3E2nOUJ04Aj
MH9HAWjIR9cjLwvKbbs0hyHwHEFoSdtmJ4mRnCewSPgEi/Z2s7OQWnHdNrufBmEE
PSTb0r2xGZrIKkLWAlMHuOcUd14Uq/WtBmOosC/rt+a+zYcV9f6mje9+KwbbzHs7
YUMRcX6n70t+/z4L2huuD4wYZ7RoRaXVR1kGEQPxsG7bwpvqIzlKHU5UZyxAjv/U
OdrxxY6lB6pu+QMP1nO0MppD21wN3W14U5MHHneu5ABGMpJruX9a+/5M+g4x8cZF
m/Coo/AqMLpKAJwCsRg5hSPp/vY4HRDHo6DtbQAEM9jj5EDvK40s666Cxy8Tpp/O
Z8akQOiItI0uE0EHhCwozqEs+K/1Gdg4WNUIXyA8fmr7jlXop9wZdKGkMCUDGDui
xy52qs1PS5V4sj2GMAYq+AJJqw2aBgl38hqhJ7qcCx7cXRLIal5G1o1eWSz7JswA
bWzvHT+cQePna/vy6M8sv67++Leyo99t7JUM3l5r30I1oHRv9umGmyiN106b3AKR
KV3lDDv6Ymrrs0vIvy0ChzFsidHTm+OHGEaDp3WbMwiKFeSV7yFzhdb6IqcPix66
WuO8aMdN1k14cW59vkjc/5Hg57GFAhv0VVCHpe4KuoZQ3D/8sHKSnv4JiSFqeSKq
vd2erBUx9XU4euTHwvzal2PmNNso5Va9mPBM6XMm4PzOk7QyQJIqaNEZn5qEdTYZ
BhX/oy2PFYWHWp3z+s5Micw1B0bYAwYqbocLAjzsRZsA3l0gxr1CN+wg2U820Kmm
Dhy8qkeX8Y0d7dVDBJEtVJFTE4+y4rVaw+4Oolq+bXYtg9IDD+huIuCAIkANf+sD
Y/MFrCpXh+nbNdqbVWYRT4aT5bBOka5i2eGb1/64g6CE3GM8gkzrdJlORIfCokke
pM0skT7ZBHWRPsb1EQadwRp5ySoevQPTUCcFsc+rDsoJqlNqPIreiK3rQu+LeNbM
u3Zmd0VA/i3SwHIifiN6lUWMkf8WinBjsctWo97JkuIno7T7JR3Pe+ezxIRS56Xm
ok1SiYfFv6IQgMpGoZ9g8aiMakXTpuJVNiVcAMcwloLWn0+JpTMOJy04cu14H4RH
KRjcsr7kMoeQoQZeHWQ6SUHeUni8niCBkXUFJYxtci6cKZQGRImhtCXEN04OXIYg
Si27d9e07/wZonYTU0bRdyoW3pVRVrJyfhRuyaE//7EQp+gi8/e4qiXKsM3dRN+h
vpEJnuVj3ioFBeaWkz5sQ3ivacgWo4txLYOv727t8s7y31/t0+HfL5opu1KbrlT+
8o0qzBAXHA2QefoRL95kotISs9NmslQ8T9P+RGQpNo4qLk7ggdg8SXGWQXTkV7R1
m4RUF9+R1xRJmoZ9/qdo5WzRm0+2i2wVCI5p/Eq0XCx28olIWeuJZkY8i7btCpqj
2dPPJeiRMUyFcR5k/2DrCDGzTDGgWePwpFuvLQn7uPM7czn9ReeI2WAexaPdPHof
7tbqFLL5eNwMtbSmz6tTek40/88k6mrYXfLaYfyKn6i6EXvJSRMLgHR9QZdwq150
wasLiZDoyHyROJGtgYxm3e385NWQHo1SO62fwaKkrMqvhuwLPU/MGNYmrfLIWsrk
yOY4VSebfBR7aHop/709lmmTzR9beSqY4EhqVRWs3TPwypXB43pCZH86xwncQkWH
d4L1UTLVVretuyAyw2zH0ovDRRXCfkZDvB1VtMoKA3hgsmyAQqIxzB/AfwE8Cb0B
nJMSWjcNeT8eRcVUoSoYH5mVt8TpWUCuekogDfoSydXlW0L2dEPvxy9mhqwHetkA
7DCOUeHrCte63ZqMlezvvdBnYA1gtsSJo2JGKBMTyD1614lshDxJ5JNF5qYlLGfs
QzAMuQx+qnTnr5LDhbWf16y8H85KhoU6nwKaLS09hrwcRysHtQEFFR3U3Zoq7Cy4
2xuBo//PYjYHgaIdcDwe5Wn7fBdBbT+eXPGTxGpDYNr7gwgPeIjUuTV3eW2CgZvQ
H8HKJKeVtVFpECtg65xAhn5mlyHaNtCVnCKFG68XEhYdpuuo95oY1W8qPv8K+bCE
izFeniAeemHKprcON5/q/Rqk8HJpZeL+rYJfWx0MOvj+uVWI8criBeEtNdn1EWI9
GB3yqN8ALodJyv5vxiMWOmyARfcGvlnd6IwHaj2MVx7IZe3HtmlcRxbBih0e1DUd
sVfTnyAwOecBMYFODwXsiuk4HPb/kRkP+fqe9RlR2us63ptB4Dr85bqicaDlrs7X
OzFXn8spc9MOp6G4BWtVOqbJMvKRBMWMSg2SfFiXPIzpfpte8yJoAXF0bEgnUlPt
Xfx6xmdqIs7BTVZbcepZxsUXKSZaSt9w+lnQfcVhzjM9zEhMYCCmxSz8AiIM4LoK
VJPTDdEiFjobFO7gIj0AV8/kGY3Zkdp3tu6nbOAut0RnY5yHVbMoaqPagigbNIts
SNA7KpJBE3KIJDvuEAsXHwAQ5+o9/a0CVPnR+iind41PHSqTiKJWZQngxEYEq3Lg
GodaHt6oRLD/Nh5HE8sKB527Qgtwg0sCaUMCwHpA0Ts2A0gZhPzqyOEGE75STdTH
/VpnmiKD6zvTI74Zw048RXM26yTfdJ+ECPyTbknXa28j2IVR+8BEPjsY6svao/jH
Y9T1H13dDsQUU3UNE8SJBehXEmhUfsZZSD4Zi4OT8yvHJ8IfZ8Vc3ey7XZiBmUKx
/XuTIKYkmCEFvGiFWpGxG+649NGajLPI4tCmfjpJ9tXWrKM3MHGUl7HXh6hv3Hqq
YjGZik7goxODv0tjA9tJuQ6emw+2FRprfIYoGEz/UphwVj8E0WDA9Djp48otf71x
M8sGtXwH4ElVWVpKTLQJX8Z7vTIXwz6Lm0qsqv1B6HBt/XRZBAlDv3cM/+OROgVg
Z54WOoTPtlNtFMhRuWT7AUdedaIDtgaT9UpccfKfinWqSdyv2y983Ky2On+LkXzY
T1yZoe1j+GSczZmgmpmG/bZIaJ3338J3VPC6doN4aJ5fyFjvNGZEM9CBCC6Nmgvm
0R5hdT5+Qr3scclZuSJ0e/8qMcNFQuTrh53I4zH6p6Mjg1+O2MalOSptWXAjNh1o
4jqffCXzvmg/nB5rryg9em0I44Br+Fx/FbBqFmUPVF2rMuHYmlpqaqxkisw9SU7o
FEoIILg4Sqpih+5s/IDtkUc6ZDkzW76HF6DLA4RpFeKqLF1EkxacUZNsNf3D3dQ5
QTbu1tihEAAWqP4WXbDdUi/Ihn0NWFefPlSDUsaJL8LVqZ4wJio650zTTOeCAiyr
ZiPT33bstqa7qDpqIsZGGGmdyuQHKF2cDP73+KthkTvDhgm7AmRPrRiKpWI0blOW
Ryyf0Zm64unVDq247chZcrSZivr0pAN6z+YEDgcSadmD1tYP/2OwJ037FLqyn11e
mvamPnMLWrHbzoXphVdN0Q3GbLqlD2z+jwEtIwhfqg2+ay04V5FP7+R1yMwZV84C
ywPZeR4aCgf6EW8e/WGgjlZRFsVizTxWjOMErHW5ITnWnR0jQ1nIRCp+1V1G7wlk
PRcmZFoYYc8L1bYBYm+26ZmaUrLy5ojiTcOBnJ9FjlPFgOpMgrli8wfuipYtV/kC
sODKu/LZXglJp+iNqisFKmxDe4JiU6bsRAAKJygHBnZW5W4umRlda5MpZHExSsuU
aI/bf5OACDdutrFuiiPDT10VyW2rVyg89qo/2TBSoDAP7vkO8LwHhExE0f/pieNG
lMTxjoPnIypGxxLJ1xsHVPjXCZcj1vz5lqWf2/ysGfVcBZbU7bLxM2moEu9SOAL9
PJHQrfxNS1XoLmKxYv6GqP3oOF6QTCzHqjSYp0a7tSOaqVatb5ZFjUJAmyZyE/Pu
k0y9FC1BXyCnOJ+fJVEq9+GfwIrDv6lhK1EPyuo+J/WaIdKEli/Ib3uOqSqjwIKv
Wq1ZgwokeNlklkpKVAv6y25b5IJo7HUtHYeeGuTVuyWT2J0/0BpjnZIh7C+xTs0r
3cgnEs3xWkxlFcuZfZYTSotewem4xrFfTnCkpta7yr/FR7NWo4Z+cwBSFcrc0DnN
KhhLRT+dRqyC4/Uff9LUXl62mhSVkbTk2cBbtRuj2Ky6MRqHVBxI2TN8O4jYR1Ox
y9OWjOxAsohOO57cUWukvpLUQmO8dqvSzH5x4b6THj4W3sl+fXGXaUjM/dnJJ8ed
j4uRtaJp2Tsbk3gA1CF2Bo4LfHauzo6ETRR075oun+Xp8ld4IaHSIPNs8pUsapYc
T2DHMjQKmMtEAHwgGi3OTXZB3wqf6dSsUVn7/aaplCnSx5Vjd+0x4YPCIGvwClPL
H8NuGHhBOsOBlB4dYD6ypF3sVF3wnX82vYcTVAWgDzzyzcKqK6dXPiRusP9tKa5s
mKVEu9VeMC/m9/Wa5Eucf2FxQDToiZbnyVPOkBcWADBTJyjvuEG1xWek/+VvbPpf
JCCkuM7SapumRTklJEuzyhuHBH+TO5ZfiyXSBzg/UsOyxn3uXox/6bta3ay6GFeI
v6CfVClBnnOJJqXZdENYpiS0KwNC7x1lJXS52BVOejHHC/SuM5rA2sWTPaAQW8aC
3sfUaXU7qgKc/3ZdAw2RSnxkACUgv0Bxff2unddpP42S9JnVLkpvR9zuzPuV5h8S
UuDQ2UHeGou+d0D703dtEP6O2YTb1zTGjdZzHrVPzUk=
`protect END_PROTECTED
