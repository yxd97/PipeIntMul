`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rNSgWYOmRVJxvSOCO5LOzo01C7niefbSsQsAQ746zBRbYncSgPNeJmFa0/5D4ega
x8UF/XpeffM1jDXEgj3t0CUVdr5p1DhjR4ePtpjOh9ETmDtctcgcLjLH1mm0o1Bf
+Jr7z6qpa3tQ9CTPdyLDV3De7FZZ3k8CUlmxKtMJ8gN1mdW2dFduExE/znlkTpi9
Iacc/qHnOCLTDVGA996r/G29XTpVJs5/k50lD75V/KpelV7oG3sGRRaZujlIfJ25
dtNlBvvrNNC7tElBqnKvUsf6HzySzfpdTpdcZpBIgPOAedNvL3H1tEZ/8oIDagRG
oQQhSMECAVWETJdghiC87ZBUbBa1o4R2w2RjUi3H5SX42SQEGXMgLS5AfPWaiGbT
Se24d7LnrIznSzQiZHUQ+sWNLy7DdtU18yZfgt0AjqZT5F45FReguy7itwMsHKgV
snb5qEv64NxfzVRjeWjl1oQt0VFflifmKzin4Y6lzh+niR1JBhEzTXSjxc90kKuI
OLtA0NWwvsFZm4MoAHj2iYA3UnXJMUJxIuNuCEucm4T9vNpUTuYiMStij88OlBnY
0oARRw4Hvj+LS4O5y2rVBZ4cs2yXx49z9Rq0lbZichN59nuCd+BAiUibeySnV1ID
hoBirOBwyB4u+oZRYYHy4tfbJHrw/CJDHzIrLVd+N2O0K/ZV4X+z4ihKEqeZNUos
6FIouSPKxFMy2Jh3kgbLS69lBCrrdFVzNKLPj+XIdduOjlU+iivtXrIywze/Zl4W
ocmFmXDkqeQcHl5GQhSyb9YjutMDjTe1Lroe6TiQZv+rRIbM6B3SU5quymdnEaVy
MMUzJSVrc1Twb+cml2HbAr1vzGCv5zGomwggaV7xXN1lyZkTk56S4gZl0zMCKqn3
Ul37cnO6yQekyZofGEWJ/Q3R1Cb4KhVQ5YEAk39KRmdJwcNh8MXsM/EC3DEZmiXD
t2Z2RKE/dyOHbIt3HBgehLvnNuZfe6daFbYJDhRu1d42Ow2nmdKL79MYq2TxTxbG
`protect END_PROTECTED
