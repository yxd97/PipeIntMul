`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYzh8ajpTdrvLrBjRCSsENS6JuwgzDOLwiiFxzKiY+3okABsetYrPm7o1s2f2pdA
hR2OaWlwbQuDXCBIt8PzPa2TTnelPppNzXaOtoQhEthv3pb7ofBbPrsZAMN2j9ig
l1gZZLXIcX+r+Go7wdh2YCcDYun+BY0A9l9INM30013/FpJFVRiM0Kz/BeWckqhW
mUZryq81Y1NfFMG7AomuGAqpSe7AQZ0pEUWFTD81gc54JMD50PKexw9mjQJp0id1
xEuty/V2x5lIU1+AoeXZIQ==
`protect END_PROTECTED
