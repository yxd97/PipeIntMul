`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+wyakJMF0eG8+RDCW8hxliMoQA46KXJr7yr1lCHiUaDBuTYExJ643seeRZjfw1H3
k4GhAn3mzst4Ev2fSnBHQqHFXddVX+KXb+spEAaEhc4PQKfi2AeNFxtLwRUffP3s
JYzOZGggL7Ul6jwGT4piyxtEMdo8Gb2aCcFi97x2LzFF36gkTyWiSK+QZRfR//eV
veUapxpJiZlm4HZcpu3/EwzOAMaQuoTl4E64/Uz7/SGmElJS+7YZ7UhjbMz19DU+
yK1+aYFpOmA2nZXMwfxSl2JurE8fax7SaABQc7YYikb3JA1hSsTrYqPd3iw1DVRx
MNZ28bbCNg8HJ5D790t08JhtwXbUrk+Fqx3duRyrxVt3YllaEmPjUinYdxaUFCQb
3vKUOsAMy22hmciyFHLRcMIl9/BomXx8x4rnSnJcRwhCbCvqT8Oxoq+XpJUe45/a
NH0ePkZTh+RMTM5TSD2VaV3w/m5tqXVBum2PQbAEZYIJqU+Jb8oCA0WuS/mRyV9X
`protect END_PROTECTED
