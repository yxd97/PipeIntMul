`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VDySAr03zzoG1n05qSgpfU9xVHplsmyEaDjp5GZkHfmHUdB3rSbK0I1ws0XhjIcF
PwuxMfTGyCuARI0gct1h2IY4iGPvxRmWS4MYqEStQ1BOjrc0j5526k9G8Xl73LOZ
yLmn0Iewf5TBVnzRAhCzC4XDqtZACCDREcr/3AqdWBff4gI+6e88pDvcH8ycpZT9
1Fw7RBFcXGaFmGyFIdTKOhFgBzWIww1bVrRl5PIk645qTHXDBL9QchLiFKHVhkpX
qYiHMvuzU6hZ3egrOK/zs5FtxMb4XXER6ZbDHW1hITVKDsybU4YCkvmG4DfbuBMs
hdOFLAgQ8w1QcviIlgi9RbVpk0IRGwR3maYODOE0WiUcEvKdTgQs8pM+/VjUAbg0
+0CgALF1i4uprw0hrqNoh3HjQTcfSL8ggXXyJoRYpNYLyIUiUb/Wn+gGpX/lLv5F
0DN3QYUE5wIr1h01tiobDieP8E+gJsHPX59ebRSwW+KG0gFMtd062ZDzgzMhlhq8
v3/W+p72lwpoK88/VKhwUe0S6fj7SgDPknmTFej496H45wlROP8+c4PfD8OHnJw+
DOEJ3J47ft2e3Oxe5CMMtdeNrFdOoIoEIsbBLF2MLijGykmc7xWZQUc6sSphzWZS
Go2Aca+JCQjWL84sltCKWeWBTaq4DR/PGKiHj2KAvSiM72cPA5aRtd6NaELpYtxq
f/d+4AwFVeJrOk/9zPLFMSXk8GEGMsmAWJ7BEHqcjs4=
`protect END_PROTECTED
