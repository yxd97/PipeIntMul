`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPpwGaWLFx4LiHSXjgw8X+cPCBAtn0sCHOLTIwYtC2UlZjd+A7agieU0U4WxM+xS
RZs8JdBcQ6SMZeOaX5MKTAn4G9XWYeS6TdCX3IknNHDmjM8rBOzzxA3RVN55NNDt
h7NoWL05socZL3csembGsJ6R2Jf01yHQvrG1rPUgNKfQRMKGtypNl7k1zX+9QKbS
nZE8chdowpeRbRbSyX5YOatbn7JCtjZ6oz9UVELwkNlGwRuYsfTEELwSNi4HN6xA
UD1wL+EJDL+bCOxsaipPfGuLXjhTABsR/HzQrhpXiGozyFha3lryAbf6iBqPZfqy
1lu1fS+ahzfaWOCVN1FlTA+nHU7J/n1zukLL80MsLvLjYcvOUXyCpqB2lzxjJUad
Du/amGtSRdGpW1Zb0yYEzXQMjt0IWGWrl6/hecT/MR7G/0JhWTDZUeN4No9tGN5B
09mrBs5ig58Sg2XLl3CNmUvC1pRbStV5gyemZhAAmx3LIHpKd2GZa1lkzmxQH5/+
81IRxoWzgw0Z0TqRdjOHXRb0IGpgeXtodA+Q6MGAZwtuuy6lQ1jhPxHjYJrI8Chx
PlzH+Jof+OoXVOuGdPblTL5BEKd2FtCnuxvhoSj8whPuxXc458EIVIm5rxJWgljU
tSbG7xdVSrBr5DvF/c3jZGTDhYIVZvQ4qHAN0OMMMk1zTMgYcJQQ5hPI5w1g1pq7
krDrDo3YoSaQPoHdWI4VKSy1GQDLJaXQH0seOXyzRJQ4X3nNDUeq1o5yLUyAIkbS
fynZcipL8YAorCg20AYVLOenTxY1TTOwGNOsN239074aclmNqQQYiWr1QL1xR4ov
aEOrX2AX1ef6sjL4otnDgN1/ItdkmQWOFO1WKnpUaMZD1LBrY/fMo7lt8MnDps5d
w/dDHC62MLbFu8ZlrpDkXfocSa+S9QFu7rrDZ7pAg/efOFdz6eW985vpeWvv95gP
3TkVve1JKDQGXchBuH5q5Qs5FG7//FGuRh+GgfwbpiXLN+u3ZLZh/q7d3HKR7dt6
Z/xpqeLzWZZJAkhoehV5AThCRdyZ/0p96RuIB/0kLgJkzusRiiNG3cx7HQGcD0LI
8T9WdhVyiRxINqHk8fbtbA4nxhD8J+7fwSai6goZSAjlKtGI7stCVrmX5raW3ZAD
kMNZAxkIIl9x68St55VAPO51fY4VmgHnlxFyKZZgyghmCI77r3VxOb0wSpAyXt5D
QwjMXTbsw5bZPH2cDmMOWcS+OyQt50QTwsX23jr28XCdIaxFHcNW99WzvyHh2ybq
3PCGAU715qPS6qr1pwuSDgw64HCeF047t58CSIStapvJAakfk4Cc5p8MbsZCvzP/
9MRB0xvAhfPeKtZQX46RA0M7J6y9JFCndI2aGXfLr5mXJWl8xV3xpo4CLYUgX08x
69FAFYNVS0BKHA3GHk7qbRvt1S13qL4tFUMNTSFO9ayLxW5dmfz+gbZuv0F9eFXc
Ig9raczkIuEA+FA6cXCWmSTSuLiVbhNFJRoc3MKyWNbNAspDseQD1qnX76DKXZ4B
Mizfwf3+KfFYP1ZF+7e2PZEG3z2VMBghcxE5OuWP1y6nigoWNqw8IXNOh80BVHpz
2HoEVd8ScWIDc2qpPPO1daZXvBgLQMbVg+4BOcquPr89yJXaKYiZghnFNpboBpBK
2cvrd+Qhf6ZqirK5tsHjqluANxgVAy5vc5rJ/ZwQi4Qzx4x2mKsIzrO7zIX+rPG3
uOCpOs0FPExz+uqNcbF9raD0xxeeiaRP6s7Jd0TXWr4G3a5uuEW5vumF2E0d24Zs
LO4DvAiduxaggsQffepAIaBG2jOksiWrUmmA1M9OlTWa6YHaWMEw/dGVSdI+dzCe
6hhnF1nDQMs4lLli9wc7jFvrKxQtuwXXtMhw/CbtYFO5Mdfh5P4hJiOjW5x7kp8J
WfOcFfQ73H4ai0ePKzosXYuEWLmVc2qpWigJleZuKRWwgZQDaYnZ4NurYwrkGn3S
5WIeIQgSj+4sem0KaWmhbAW1T9oQDCFIJbllexzJhqXSTCgLzrYHuXv5v6/IhP1p
Si37EYfiGxBsHxmfGC7mZ9RaSpJGrw9NFoDr6ilRDH6T+AQqQvjpVUSegGAq7R/9
nbXrRRAhXkyZKjApjXxU+sS16A4uMbdHrZO3v1LV5Xnhd4TQ0DkZvvKymxGsd01u
c/s0A331Vy/dzcGJOemj0AcKqVQwcoEpa/t4bPwv4NGBl2DRX5q2+QfVaFIZSdrN
wdMMAdbYHItinXSWRdRgxqPMk10ZymUbnzdydCwEfB71aLLDzZG0cMumf89vF6VV
U9FRvWON8MgJLsGrLnt+0gCIKwFyWGuqUUC4COKhdROqvksAeGmSLxiLWxTkzswK
FUYdyWlEUtarkxrvfv+EJRy0h5XWX7SgLE+Hq2ag9VfeZI8EoSOL3Hs15hxcnqII
a/6zJFBJqksFIlktJwzxYmvMbVae4R3QV8ZYuttsktyhZAXogoBFXF0Btd/TlS4w
6E4sGANkMeRersf3H0zVxCx73Gt4CewQxYANpuj4BII39JDj8nGCpTnvUWjdDYkS
BeW068q6X0RX2U+z4VFZZ5kV2lftf7NagV5zwrMHi71ePG0kzl0igOZQZsYhKFqh
Kf7YFB5z6le8d55cmAL4StsgkQNty3htvmxROGB0pF7jPtdi+TDHqk5DVCw+i6Ro
KgG6hTvr+AS2l791cgERUZhe7q4GRyELLV+A1GdPj3y0XTeSt46U6nyvqmj5YtKU
5dSca4kRdF9iZTyThzQSMPkQJJPcnp3Ml5y61xlkzdeiRnDC/yI45CGb+jL0iJFy
8+oPQcx65DXZajeOkabbms6oobpaJ2gvAq+RudBOP5UzZMUgG0bmxP23j91iRqRC
h07wtWpCQln/EJcH/vqMnlnJNAFWRYdCO7qdUQ2VseAt9N2g/lBE8h8jXXGeSEP3
imbhkOtzj0WGTPu3dsW+NzlPgba07kscqWCycc9+XyOVCP8sF8NcBJeItgLOS+6U
50kcZ1mvOv+LUy8iJWdqMwYmKQfNjbPAsRteg6QwGBURZXNJ2LBTqui4ET0fWuin
FMaala78Z7CSlzvTKL9HK44suwtD85IQbg2m7M8djaxxcvDhakdtMIoHcI1nr9uY
qEFe23GtetT2xk14odS3m7k2Dc5g2WL/XBH+75MYTTFBrVp/3gYy7ookSvhxXGJO
ux90AW63zHwXwhtDBjJPSb01bbqW4RfhdK9GQHKS2Z4cxsB/gXV1cNhvS9+4pBTh
INl54yKTL/zvJ9K5CT6ldX28/gtmlkKLrpRZoGEULSVS52MUcPvN6EZyMGoZzD3+
+LiK8NiE46y/XJ7gP8/AHIaZbrUTCRZxexCyM7tfj3cLKSUNSFsbM8t2kwnmDueK
v/cxE8SLwlmMojPFQNl0NO/RgLYk8p2ALGCyeukM5YxyN1QsOkCMAG+dodwqL3Do
bnXGpbQ6G+axBjI8xT7O1cC3ZGkDGyQyHgZ/fYeTMan5l9PLTlcvL28I0QdL9zlg
Wte/tC0EkeENJPAKuJ8ww29vvs/Gvo+J0Hh5wJOYSunRvr77zFF9dYTUv67oO1y9
0MIG9RfslqcqPAJTPhD0ZU0CsYcNyo5FnYN6nE00/ZD5KiZqV94ympH9jManWorw
0rxkL/BfZHSHDoOkqS3AlphbrobfsqGJ1gsQzpL0eLzjvhCB12aN1TykpA71Pzou
FD8hTUNu3/F2qC74XabW9DMkPO20dgOVIDhhP8QoyXAnFjwWnt31JloSMNrWQtuR
kXX9aSAjEtczPLp1xr94yjdElyvV7AMVgWL6qYiTxX8C50oW7E6duQ/pXhDLYAmc
Xv/SlXBGtCGRrDkM41EcKmOqkokmWhlVY+2f4alGBg630ZALyAjMSLoCENGWSsvT
BREzxIo3TuuF5IELHik4m6vXakDSUDKxN8rE4+tTQJJXkpDLr20+3zekPzuR0O45
CMgw7emptNHzYd0ZMWn4D8+XJWQ07iBto1MmiyjQRyt+StA/FtwtnbbMGxZ+gSxs
FShRMOcfYj8P3kWTd2SknibK229+zqmDS/T3cu+di0XSfvM4Mna5DhlSmyCLuJdW
LREaZ67kkT49JHAAgKdckfOnp8gw+VdL/lFVBtLRaTtFigWOk7JoQhLooiuWLS8q
dfl9rBDMuVBy/CFEOile65RxjBqmuwonHYGyFAnSMfRTAb+mRj1GMTu9E3jjKOQC
qXLCnHUh4JxzGxlA5uexn3siYmCP15FDEqpGNEzdlfhbf284AwA+Ug8VmlR25NVa
ft7ug1TDJtZXHLWuZEYe9TOTT50jLHHLEnV4/oRDgCUsftLsgGGbwWamrDjX0tBz
k8DSlQllp6eTrlv4g3x37Tp4vfY1MAMKA9C6z8UhO4v/w62hc2uPmAi18qVqfcK+
7LYE1JRWPToiV8rnjlqrGm0LMPoz2OuRS/NGDw7CtNEWB/rxmIY5+oE/r24C59Jt
tHaOog8xE3joy0D0FLWZxPLfS0AZSzQ+IL6/anOZ97CGRIW9Rlk7HwmJxwxd1nJ6
uvt0k2JKZZgT+47aOI6Cz1PSdWphJ2bDlH8Df3NanZTR/hT4G2naE7llcMCt/B9q
OMOICz8jK7jHJ16WbxjlTZFcicuRkjitgfApdeSHLwQJ7JjEsv+CSFQMdT2Vbmwt
8b3DpJmNwiI3c/ttSic0j4nhX3PP7UlsV9Wfw2xCWSHrk3bTc1k7rkK5c7xpVXmn
megFyJD++uiAOZVecRZYdnAGU4gQIpHw4ioDCUZqoellypiiKz5BSWcEJV92GfTt
mV7a27PBff62ezESXp0nrVZ4ZG7zdXz64emFWXtZAcaKtShRZy7HqgN+KWMezPF9
E7U5l5NmS5OKbPds7fxjP1nk1tSUuW8LezSV0sLPy2/poqleMdcMyrYoqTUwIiPd
BJ61SNyc86VHS38lVoE2VCY/jdWtRxvUHcEOPZZa8t09NJ5lxQbJo7bDoqsnCIQu
i8DZneKGFKbrzHAdD3OIrMrDwHxygL+ndfaoAh7E+y6ktiaIfJn5CJJQ2R11qZmd
WeFqhhPCoPvhDs64rpI7ZrAt02KtddvYCB/VCrcE61JDyfqx0heghP8RPOwsy9DX
aiuEBGFVkkwbLq0WQOKk3sYPPsBGxKCrFYYjMJmhixrMlQCJ6iyVez2gRhUngnnB
oaWchmchFOuBvuTshSAgWHUmunVBzQrjMDIPQctL0dvLEr0Fd8G0jRBEq1KYAJ32
HslPbOgMYQcE62+CIeFgiTOfFg/5mWtsGZWlxRWvhG3UoF4jf6TeExmk65TUJ2RD
Z55CUmOZRLb0JKKZSaWcvJ/fg9PNC/oX6uhsHni4II5zk0XyAhiiMGcAWUDS8y4S
xRlnmiGFIyJZJ7VmJ8ZecMPpRUjvN0ntNfvLOnsi94BWNj+Ki4UE8CrcscqpT5T8
RnRx/Y/5Vl9R2UwMGe9i+uGWXMiPOFy9Jaw+LwSIllWhuiLw2IAOaignuPVEeZYg
Wd/+GiL0PMNyeh4c0FP8GQG3DJaLLvZfoglJlNuyiCYQXq20x6tSNwG+a8df6cX2
z43vlsWboJ1DVowXlXN5KaFbjUKNVsKGpHV5BTunvPYOwHhgDT8YBULUIe67OY7P
`protect END_PROTECTED
