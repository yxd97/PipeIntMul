`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+g/R2JsLmAxMXyimWJarfkyphFXX3aTmpWY4yfdR9B0WYHKoX6WJ989qh0K8q7o
MqJt4bsS5W4Tj1O6G2YvCHFmlarpbOaIf5PVNLjbx5oRgtIMyUjh0wZP2gJq5w1h
MFVrYGZrkoIDucgnNBr+Upn/ABtzS7nFDQCm9U74HYh4WNhG/OD1EO1XpXGMd5hm
vjuJoyV87v8K/pauummcPWEU0j1Otmt+c/9v4oDs1pjLdp//Sh/h0jqiTq+2EbHJ
veE/c5ZyU1FbO3oqmgnFudAT5uXtaZyHyliRVY7xbLZmkVQ5JlvVjQn2sbCH7jJE
eft21MzpaTNGo/Wb1eSBzH0rCAVZHB4nPc+4tZtpQM4rL91Y6XgDkuHNQdWSkGK3
Gn3MYNb9sXfHPFWteic2GIPJPQxrJ2saJXRfD33MHVpYFYR8l3jYwLIIp1wY7f16
Id1EkV4lI0yOF7tVmB1R8OAC5N6E0zNkP40kSVhxlfw6xsVL6zkfBSYWUbOklSJS
V3jHFSPSzGPld7zAXujr4FhmxGU/QbUQ9EPUWgo8Zq/zT79Hb/rC56Zwmp4pq+z4
9jdA8Jnk/cuTqYBYU/8zAVP+Z28Z8GVrfgpegHH/beQPz4jVIGo6AgTawQ/Z6wIg
28+dAQtHkRGtXXjw0xG0m4HCI+6J6goIB39mfJey0A25iR4w4ymtEv6921v53lCJ
jl2h8HiGPPqVnoRLb1hkm7kCbheK116DkmMrj5yzioIsw9Kca0bFj6cRzW0uI1SI
JLkzOMB7Iu4t+I6hGkyPQUbIisOoImD2v+KYItpD/B+CuQfHJmWUR3mnKka5iJzb
k4Dc1Iau9xKBMEyhQIEvDuJ0v/DyrmR5hS+gla2jk4ExtD2YMKG2//7GcgPnWmgp
6ceCKuoGicJKwOdK9m7A1QbKjGbXrfd2kBD/sRl09DH1OL+NlRLT3vpPqPWYi+9f
fdWhitCuP2PFZnuSZvj/LOfndDr5mcOZrBhQINEMStLyfAGlyYLsLg90qrB7a+jx
WYD8PpKtVaBMZ1KJjV6ozbgix3sCzG5O2X/ZA5MFYORTctSF0P8FmzNsQfkxpSLw
LXs9nx/yUaJjVl8tO77fa+6nzVRbGABRoF0i2ZR0xH20J546s5yWIuHrpZZ5EgTg
BwIr3TbCa/5BSb/7P0BDJQetg4zWZsuzc2iVAypumIId4HDumn4eL9AiMuRUuXr2
AXqMw8ioL1cyZjuoX1lWIPQjPt8/dDm+tHGXdajMnrWSiB59h3QffdTKm7rTFzH9
Uk2OlObYe8exOMacJhcqDPgNpOdwDHzyz0rRNORCGU+cgIV5kskBhbIbrLM/ZGGj
qPQAdQZjxNJaOQNMot4E91bOKcsQIZyjuoNWIxCLSMHbCsAdej2X5y4BC9MaewU1
tQeCT2ttpRYtdDF4QuXl6HjhbYZ0ph/QeXsCwluX89P3Us2IhdixyI/Rq8XSmUmK
OaPE+mLu6nDXQunLefBdduVSy7DbRNeMkexFpiyNR47GORCdKPR/vXmPeQRgOEk0
`protect END_PROTECTED
