`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ERSQ4GfawK80lagvJ5VtwAMIopkS39+nrkiviGkbi8xLBUlCMnew+olRkpTtjUTV
aZjL6SB1iqKxyeEoxQwXwhKyhePFacd5bjjKygigs71HatAcMNUUgyfwoUuou5jg
ekWZ3vM28CTac5puZSaqa3r7UZKd69tErzsjMLD+ZhgQGIL73+/VZnKvpMRxtNAy
n2GLPcShVBYTAqLzAPfchMRYTny+r923VBN9oAzXz0JpysO6YYwCgiyR1dklenLY
DH++D9aH2DmYHlp/MnQ8T3DTDm8PTzlMTXYrYQKm04Wbx56FHcjOhg36alluWjfb
4Ylcj0fHfzRnP9srdTQ9Mkf66hsCGVAQCAy0YZDfkPG2HX8ccu5KHvp07LJ8QvQw
c6yWplu6jJAcSv0P1qmMqriux0h1UZwmDitIYfzc4kLVcP37pTDi3lgEqCPeXYsJ
/ARswGL5yoDEL29RQ4LNKMxierVGaYlNyK+1SO/7/+flj5RVHHqzt70hbITOur69
YZGPgjL5FTN5tQhAbUW1oof68IxVP7Pe/xoBM38yPok+8g0nMulEbQnu+HaZeL33
9MAAIBJjrCQChxiOPO3L4g==
`protect END_PROTECTED
