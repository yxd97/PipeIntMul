`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qyzOCzgYJJrK0aglSOjuEygvgtYDS7p/ceu/CHQ5Zthj5f4uJzZ5zkFWWY3zvDAS
km5oFG9hwvueFjRKA1V7dA2c/9Gojol5wKamfCBqS/BgVmlLk6r4zmiKXwn2FojM
QwjkLUdJ6PvaUU3I7357BnLPRYATaxjD4kJKNmxpESW6vFlWh/JuL5YIOAIfO56f
LFas0/XZF8LxQarLwCgVImymxe7b99jdY2IxTL+MR9yEnVzzV1lK7JFqY2940uvE
j43NrAYwwrnbsvbjuatrsqaOI1xBgMIgRBH8TKb3HvcNK6T8aZgxUDGKoDnoL/fj
MucnKhV2qnebqVY51ftaDEf6VwZcLGN/YlyDDKwWJIdal70xUfN5QRllC3/YJd4K
vJNudiKC2ldR/K6QQRlzuAFC3U6l00gO0fEYNz5+CLeJ3EPunYn5IWiWjlp8kaS7
CcPgkjv/GBr9+w00/jAjA3R7voNMQZmvMqdRaLirlrflhxsC1CTQqbZ4XYSOXlwu
wEdNID70Rvv3k8+7YJHC0sJlXQvW8W0G+66t/v1IVZwzaXKn9C0AuDLrra2WBF2C
SQT1C414qc6d6HHKSGk4m7FG5oTpUxN08v3Ku/5bmNmElBxS4YZthEwp/8iaH5/D
o/dn3fYKp4wjbVGmsTeFoOmrldpEQu1aVxWaWgxdhK4I+B04rfOwIgwytHvfyRfn
pg/HictjrQpR9Li90gfp2DKMzAVxp2jm2CZK+yPn8Xk575GiuQ2yuEK3TvaQYss+
ua1hJNiHjTEiIFtIab9z90DAWPC/10KXxICQL+w88Z4798vp7z8oYxP2xn8nZgNc
t8NeZjE+N9XiU4S6QvURz+/3ozh2JEcTi+YS9gqBoAB+YejcIvSz+X5j5Neymv+h
MFH3K6pX0rXxTQ1k3QH7gw==
`protect END_PROTECTED
