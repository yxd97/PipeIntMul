`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qtQNNt9ZBxyDoLb3OOxVKecTxxwZxknxxmSNSw9nSXJHA2WLptT6DCbAB4gvYVk8
C1T5U10DNX7P3r7V2s+z5xV1JiqnEnFPVZkA/tql8RAs1BSf/Y5dAl1Uuz+LCjhr
32iRFILyz9XPkzc3/UL1nT0lOaBM74tq37VSsm2/67LyxlviOy4C40YnoRjAuL53
GQxxRZHtbZDLipS0yNgomhvElb9QWBpKBiYE86VltKkVsRspSZIrRpXla2YKSN2u
b1MJ4ZSv+yzAsrnu4uS/fg==
`protect END_PROTECTED
