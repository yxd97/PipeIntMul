`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQ4LafZoBZVfZ+Y9MYl+odFj2i86E+aP078Du/e1DjemctXqWTSmSzwZOfnuS76V
TOwAwW1as9WI35c/AMCt+RVfU+Bb3MNdIg2ecENcWKDYDdJvx1TUGyCfv+kfcC0A
qkKMtU8aOoDQG/t3Rcx8s9d5BLVQNChVLSojmcag5QavxGYNM9jjKTcmQ8SwKn5T
6dZwnp0zSSGy77zc2mcz5Rc0pQJQ/caPHEIJeddHZeDtmcV80Mv+EBl5wKC+s+jA
oFAHfpGZwYrfktqOqaHKiao1bYyHO0JT+As/fA6c4W4ciKx4ZkGMhpnUNY9B/U6G
W5lroRU7IrFkr5OruCKbDARCYknZtJEQ9+3bnrRvYrbDzx6ejr2f8GdkOE0lGwPr
5WQQenQbKr68AhhMUDRtIRtik/8QE9LmD98GdfBA76cexkxOPi5k+UqmlwALP2Kp
IBgJPHZDEQWjiA4CHjQGk2O7FWNyJAKO3c7Q9nA2ZauW1tviCSRvLjHkStL5YOK+
qj68J+qaA6+AW5BtfyWcmXV7YjEf88qPRprTmIRoGJF/xeHhKu6FnpPtV3g31vhn
7n8kXEPyKq+5iKeYrmsQlzjz5m3YoHXWgP/FNijrSfqMWbcaZnpHULdTmrUi5TLt
3HwpPS2kv/MKYG1ehXxPBTocF+vtufncA1WyqzGOS6H4OFG+lXUE5Gehyd2KnlDg
PG3Q9WE3yFaW/tRaKEklkr3HDRvsaf/rtCSez2ZVV/a/vRhAebobX6WzBmOiIG3b
`protect END_PROTECTED
