`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjfWb+PknYLh1jt79zA38t+nlwMBtoy2G7lGwNgsyCtZw3FXIHaDjcSDTjOCDSgx
SP/PcjfB0XkKU5PcsLFBwaEtNJrq0LeGuM7iQPfL4EcIZlH9bkPVcXrkE9GTlmQ+
mtKYZAsPHdEVTmyy9fP6IVNLnTB+Bq5mOQnavOj5rxmyh6wBa9ugJItqpVZq7a2P
HSEcaY10ELOUzkgHvRoTIZOLmhpFbyHvGwzdiTB9Z4MLi7k8ND6TQe0+sX3RWaVL
yMW7vLe+9IVu9RdAFVnxlQCKPzrWQBvx/U1eO8WIiZO9RoLL2ohw8CX5NKiV2pOZ
v1iXu8vtU+JWA0lzbi55rypvbLFUeb5UeEdqqM2AbhYKyCzQ3EBEcpLC7yyTLlNB
3YayBxKhQ9FYwzHs8DvA7jsu99xrbmfrx6F6QkpE5Bwbwh1RP6drRlqdW2KCooXp
gh2AQvzBbGVLHWu6VuLc34r0kmUjivFghwAFbmsVTexR4B7uUzVi+7cJYJR/m9gP
6FxwAysnxCaivnrCdyc3zvdhqz2mC9WDGQ7W/k2GOw8=
`protect END_PROTECTED
