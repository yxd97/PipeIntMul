`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSnpr0wsY9vny55JuGqvnbscBg0CGMXBT9Jx4FRDsNsy4KVcsuLzw3KLBMfppMIj
/80YRssmly3nLp2N4J6u96yjiWCl2/BZOF0peflG5lQL17EyEZtQcxvKv/VAazlX
d+plimPXfsbORJVTyxsKWlzDN8O25UN3Det5CSbwq2uJAI/uUWjljzPeav4sAHih
eBATvpG48LCGBVlE06gGe3Gm1ki75Q9QH3m7U9X0wPFouoxAuuJqHaGTmd0s06QD
bM3/SoLiMkzVGy06sJ3ifREcUF8TWtbwe7FHrqALWcSjVDlCEhJot9rtbQCN9vLH
zgzYx2l34fmrO2ri6hMmzY3COsH2sh28hPCYkjc8T+UWmAUviaO4qXh0WqL8xHHv
TtbCxGsFyP3AsL5p68u9O7cv6mJOG45pSaHhsdcbdeJbfhkxjqqS55Ef9gC1+/ug
tCGZewGozHdxJhhrH1sog4lJJ4zxxS5NDvvpFmtMvFqyLd145uVr3lry9N6VJqdI
7/B8AeYlDsW0+IQGn5pDTJWQ894T+PMTy1Jv5bISth/0SJB7pDzzvir6jTckdIHt
vO9epI3rDLy8SmSIsKbL8szsk/QolBxSiJ8g2OmAKs8MYCoXIYJrGAHW2I4iGwlA
d/2WI6PoypATjaYp3m9Bnw==
`protect END_PROTECTED
