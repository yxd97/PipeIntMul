`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xri+qI1OmIdNXdH7gGT69esrq0iAuqIg7lN1IShzQZMdAVekh7ZS3dacTDqDz3Pq
8KyS+jUhh3YTqvitUYPpAHJ7NlKmgQ/xsQsC9Z8cltBOouRjHzAgLTY6eHnqKW4I
sFJ0siOKu94m/5OSTPmzlvko3yemP9A6MtUlj3DsyJ7XKvoB0O48sjddAb3KZ2XF
t7vKfRP+7wauWjSLdSotBxpXPuzDA5jtgobENwPk+JMmATu4lzQdt7huyqFuuEGq
vsrDMg7RIeVIvEhRSzPRnV3mm27f7791bX32zkxGm2uaMfXUqsLGK/MMk7fHXxXa
ykVWc7DH7Oe5tnTVhSx693GiJUycLlhyNsc4bv3dGYM5JKIm5vG9dkbArMzlmPAG
o0xK3aUnzMjmu5xJKGSnFt4MuAt44vBCdGThH8A0d5VODZ3uweY+UuVsP5RzIqOS
Hm01rpQlWEFR/LkmCiR/9o44xY6B0dl7KD4/tX0a0989sILXgWzJEKdZs+8SuIaS
1F2BWFGt0dmJHjQ3iSBBAm0ue28gW3ctwC0ZNtc89wU=
`protect END_PROTECTED
