`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ach3VjulDyYH2wFyoWncSbjswG13R6/ZnJ4p1JGKlepqD2x1vY9EID8CJNRNHqRk
EbzeslvYAaxroFISsIM7y3WEv8z7NmdNuBffcUFOHQ1IDVCz6i6L8UnACvWbzquv
YEKvTtSuhLIQYV4AhFwZpmIznJCV5ABVzwwbsDIl7/iYkemNToeAEdYRJBoYNFbs
YOS0h7VSD1o+H+pIsyhO3aDv8jZQ+sivf7PuR3YK+IQjgFkoKUWhHznovFBX8U7E
yaHysxdM/T4R8d3JTOh+7WAiEWYgzNQs3ggURfNzPs/bUK9tnsshcwSuUpdlNYLF
6BeCOhOMRjSD86RTDawVJ6SjM6Jzj7w1TCEksxNYh4Gwk9Dv4eIWfFIxcBzKA+J8
JKsIpUXoeVvmrLAP2vRuff0uqziVkUNgffYDzBOsBzw03yP8dAOgOjn4lhdn5p2n
zuZ/tiBqeYQZVMhCQpu6Jw==
`protect END_PROTECTED
