`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riEwKNhKpsD3QXs6ByeW2WwtfGrNndbAcpz/gHaRq7F6qO4LXr4fmsA1BD0zszgU
KFzRpNmSd3RaPDFeurbqJuxLN+Fh6I/yqKyqkZJBaJWyqPQZ/kwKAWaRzVdycKtA
G0yymxj7dIKoQgg0Uu8lr81ZpmYpGMgluGNp44oyhN8JrhJTuUyzf1nQicokXtro
DVBr0qoaYggw6VThc71SoWdgbERZ5pD7jwlrrRNXl5qkRcLOjwMiuRBwcIZE3zXX
w7IKE97mzpiDx+t0f2qOJWQGKysmIkfMU5X1c6w8k7WGE6pICQJTVSfpYPB+M5Mp
QhhfLj2pUg7n59yhEcV1k2qEVO+UmjM2xKbVvFgmjQblONwCJ62icCGGKchLzAcZ
kevN+YZJCkH8zBCH18d5xg==
`protect END_PROTECTED
