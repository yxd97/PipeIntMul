library verilog;
use verilog.vl_types.all;
entity X_DSP48E1 is
    generic(
        ACASCREG        : integer := 1;
        ADREG           : integer := 1;
        ALUMODEREG      : integer := 1;
        AREG            : integer := 1;
        AUTORESET_PATDET: string  := "NO_RESET";
        A_INPUT         : string  := "DIRECT";
        BCASCREG        : integer := 1;
        BREG            : integer := 1;
        B_INPUT         : string  := "DIRECT";
        CARRYINREG      : integer := 1;
        CARRYINSELREG   : integer := 1;
        CREG            : integer := 1;
        DREG            : integer := 1;
        INMODEREG       : integer := 1;
        MASK            : vl_logic_vector(0 to 47) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        MREG            : integer := 1;
        OPMODEREG       : integer := 1;
        PATTERN         : vl_logic_vector(0 to 47) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PREG            : integer := 1;
        SEL_MASK        : string  := "MASK";
        SEL_PATTERN     : string  := "PATTERN";
        USE_DPORT       : string  := "FALSE";
        USE_MULT        : string  := "MULTIPLY";
        USE_PATTERN_DETECT: string  := "NO_PATDET";
        USE_SIMD        : string  := "ONE48";
        LOC             : string  := "UNPLACED"
    );
    port(
        ACOUT           : out    vl_logic_vector(29 downto 0);
        BCOUT           : out    vl_logic_vector(17 downto 0);
        CARRYCASCOUT    : out    vl_logic;
        CARRYOUT        : out    vl_logic_vector(3 downto 0);
        MULTSIGNOUT     : out    vl_logic;
        OVERFLOW        : out    vl_logic;
        P               : out    vl_logic_vector(47 downto 0);
        PATTERNBDETECT  : out    vl_logic;
        PATTERNDETECT   : out    vl_logic;
        PCOUT           : out    vl_logic_vector(47 downto 0);
        UNDERFLOW       : out    vl_logic;
        A               : in     vl_logic_vector(29 downto 0);
        ACIN            : in     vl_logic_vector(29 downto 0);
        ALUMODE         : in     vl_logic_vector(3 downto 0);
        B               : in     vl_logic_vector(17 downto 0);
        BCIN            : in     vl_logic_vector(17 downto 0);
        C               : in     vl_logic_vector(47 downto 0);
        CARRYCASCIN     : in     vl_logic;
        CARRYIN         : in     vl_logic;
        CARRYINSEL      : in     vl_logic_vector(2 downto 0);
        CEA1            : in     vl_logic;
        CEA2            : in     vl_logic;
        CEAD            : in     vl_logic;
        CEALUMODE       : in     vl_logic;
        CEB1            : in     vl_logic;
        CEB2            : in     vl_logic;
        CEC             : in     vl_logic;
        CECARRYIN       : in     vl_logic;
        CECTRL          : in     vl_logic;
        CED             : in     vl_logic;
        CEINMODE        : in     vl_logic;
        CEM             : in     vl_logic;
        CEP             : in     vl_logic;
        CLK             : in     vl_logic;
        D               : in     vl_logic_vector(24 downto 0);
        INMODE          : in     vl_logic_vector(4 downto 0);
        MULTSIGNIN      : in     vl_logic;
        OPMODE          : in     vl_logic_vector(6 downto 0);
        PCIN            : in     vl_logic_vector(47 downto 0);
        RSTA            : in     vl_logic;
        RSTALLCARRYIN   : in     vl_logic;
        RSTALUMODE      : in     vl_logic;
        RSTB            : in     vl_logic;
        RSTC            : in     vl_logic;
        RSTCTRL         : in     vl_logic;
        RSTD            : in     vl_logic;
        RSTINMODE       : in     vl_logic;
        RSTM            : in     vl_logic;
        RSTP            : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ACASCREG : constant is 2;
    attribute mti_svvh_generic_type of ADREG : constant is 2;
    attribute mti_svvh_generic_type of ALUMODEREG : constant is 2;
    attribute mti_svvh_generic_type of AREG : constant is 2;
    attribute mti_svvh_generic_type of AUTORESET_PATDET : constant is 1;
    attribute mti_svvh_generic_type of A_INPUT : constant is 1;
    attribute mti_svvh_generic_type of BCASCREG : constant is 2;
    attribute mti_svvh_generic_type of BREG : constant is 2;
    attribute mti_svvh_generic_type of B_INPUT : constant is 1;
    attribute mti_svvh_generic_type of CARRYINREG : constant is 2;
    attribute mti_svvh_generic_type of CARRYINSELREG : constant is 2;
    attribute mti_svvh_generic_type of CREG : constant is 2;
    attribute mti_svvh_generic_type of DREG : constant is 2;
    attribute mti_svvh_generic_type of INMODEREG : constant is 2;
    attribute mti_svvh_generic_type of MASK : constant is 1;
    attribute mti_svvh_generic_type of MREG : constant is 2;
    attribute mti_svvh_generic_type of OPMODEREG : constant is 2;
    attribute mti_svvh_generic_type of PATTERN : constant is 1;
    attribute mti_svvh_generic_type of PREG : constant is 2;
    attribute mti_svvh_generic_type of SEL_MASK : constant is 1;
    attribute mti_svvh_generic_type of SEL_PATTERN : constant is 1;
    attribute mti_svvh_generic_type of USE_DPORT : constant is 1;
    attribute mti_svvh_generic_type of USE_MULT : constant is 1;
    attribute mti_svvh_generic_type of USE_PATTERN_DETECT : constant is 1;
    attribute mti_svvh_generic_type of USE_SIMD : constant is 1;
    attribute mti_svvh_generic_type of LOC : constant is 1;
end X_DSP48E1;
