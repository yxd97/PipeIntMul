`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jgLoPL6oaSAHfonoW0A0fNUqr+RVDaaTfg4523EzM0A+FiAR4yqseP5pPs8tzsxA
4KWG24m1B6Gggg+HbUIWT6LhLR8PAY0hgYMChQNwXpcOleb66U1icyLKUYJ/KjR6
XvQLqLTJv5Bh7ahE+Qt6WF6mJmZQbRElls1qBuY9CIdMeBi7HZRGCiD/gRoFquWE
7MkWgsL7u19oevG3h++zfRi+zxdket3ClYA0AfLZoVyoxwGM7PdYkLf4Xgebts7J
0IP4XDTzJ0eAWCv2xupB0anfVB760owtAHJz0mO8MwB1jt4eqK5ZTDBC6QGskdp9
LZVXuafSk0WuC6RAH6uYBA==
`protect END_PROTECTED
