`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TXULGWJylPrUEWOT9nmUm+3J7PxdC6uicKvjVOR5Eg4+oP8W8JMjRg63c3PmR2G4
obD//J/ki2XUrzW/rOWf5JD4SSJBtOI/BXtBN0POXcbDGEnTs+T7wT+7K/cEcAQO
XixywK1WS34A+7GI1wJE4KeHkDgkkrRRxfSWXfyLsiQN6bWVaMCX1qm7dU14F50l
nLQIo7xXY/MYQrO1n0xX8ql7stCAKogVBC3IO9JH2RaqTcyln++uPM3VY0kl7Y08
CEsfd6v6M2AwwkAMQ7UdS8H7xQ5x7efO6ggqg67v2JRa1yaTHDd4lE5bPoyYLAEF
uQh1rqiUKAzfj/YQWAcW9J3UWbBFZlmXijDMB+NyNq54bcGKQnYX63qkt+L5hOtF
`protect END_PROTECTED
