`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IewMnmthxi3SG80oqDE47ZkibacD0ei5v83m/uxjiJg+1Az9eIRbriKcmgfSnqBe
R9G0XKu+OUqcRp5qJPg3faX9kXnePcHPppecL2sUmprhW1Dgh8Zw0v+oe13WFFpe
wrA7iZiViXUi5vQ6elPReCRt000/pyUaXjDYZBk0XzeFbZ1UbIv5f8M2aOWNrgYe
XCgAjwbZPKJE1taXxsRrH+KsSEwVsWN3SlVRitDtQRedXwdZkZDrIOV5xV1DDr7N
Bx+V/mxPCIZ2KiJodry5lIkdSLxfmZOo+LTGxDQwwYJDai2AqkRLfln6Bp0nKJry
ZqUGfv9AZ9tb7GJZrBKU2i+dnVwOWtHiB8+jopA2nWnYwrMrVsBkladEUrM0fmYh
7wa3JzUVTC0CG2FnS7AH1IAu6pnvfsxgJXT7XJoj2UTmezktLyqNS1syUlUuHCKM
mNq9Mxz+GYy3WOPzqU4Ukd3hoOtr6ltdYc5vlmfLd+Y3zMZ/vdPJueNuThFz0x4A
RhTRdGoy8NGhPRKTcFctpZ1XGchfEu+Ql39MJkNTeUuxWf9mqX0l8xVn+Muxphi8
y/nRP/fGnabxksNYGIx3i3ICqY530OSIEcmeNdofFAU=
`protect END_PROTECTED
