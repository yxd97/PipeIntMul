`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zb5RInaTTgMqkP6bldVNZnYIuzwdmb+TDxM+OXi11c3tYo6LlhYzpZKnEKnSpRum
LCmt9XbAcE5+4JFisYnMUMcWCoYj0yheeAQmolow0vSogvegCZq455DzRvl40w6m
t653Fry0Joc/KzXPgw26JfhlCXzC+Xb3ZCjwTnePwkoGvapREvmVCsDZkKKFJYLF
A36LgGQE/2Eo/NnVY/ahvMgrSMiAuRG5qEXMmfFkT5lj1aBIPgs6eE0N50obetcg
SVcZ+eVSoxwqJ1tiIq48vvh3rNPrGE1CNZYHdEdG3MLmg10ZSyK4KvClhuX69rwT
UX3pgXTwRknVEGqab7cHDGFTwD05g97nd/VYi/tpkHjtzGWwIngHutA0kb5D66Yz
4y/qMcBI2hujNLntOY8M1TKNWMrVC5UKbfy8URPpOjKWF/zhkhA30G8xLYCpwlWg
7sRB480nYLEbqemz609Pc4Rtx7XjC5THKA3lPFe7inxntZ6/GW9nXRiRKqfQlf1x
rF18sc4e7Wj8k9+tLxohv1tF3a57Tl8q58FUh1FSs1r427FCid8fgEbgEne+BHnK
`protect END_PROTECTED
