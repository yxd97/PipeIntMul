`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2HxS3W3Gpo6kZU2TP+IHinjleMHJelcp9mcLkMNe4/DnpXMhd4p2QbxexDJKAoA
mRFE7d9eEXIodidtopfChqIM01r1XgksAem58te7DQwFaSCSyHAUvMv6lOLMl89q
TjRYRApvhsNbGnSKrToLkYh1exITMH/7wg/8xktdr9Byp7IRe23hHfBuih4lMS7X
lgE8bazmUXaAUiwMrpJq7p8yMryV39J9kvcra6Nzx6zHLn+2ZbCMYmYmAqRfjCc3
h1thg+XLJP0txBwboZR1TY1umriessk8inAyoWwPTRFCs3hiKRxL2/q3zBnslwoE
uhH/oHV+8V7D9n0tAolfg5TAiS2wvvDnNfAVpo8UFYIrgIo8TT602nMoi4J8htMN
lUeUAtEcc4P1fbTi+Og6XI58Ewc0zneZxU4dPEIbseTrheRfHFPN/7dSp19S4Iv5
Y6/zMJ7zNAPuPDbxv3INCHW7nvQPb6CANiAkwhDBKm2DCR6kp3v9sjuu5N5QPNfo
uSQu/gx3TfZNKC3uEX+Oe4IXBvyb78FIRvzThOuZo4CayFfWT7wg4nUKtcjCD3f8
8SOGYHiPMJw+s/4FTqfPGyTpj2vM8awqU2Rk2Iu5t9XF5dSeRufVTRKDL8I6Y/aI
SpmLlpdxnJPduFwzHDYXgJiUEzbPP4wbPga2tRA5LBw7fIe/669kCTmcF7MHxq5v
Ga1QUaI0lUNhIMl1maFh30WWz/h+qHlHJECgR6DFpN/KnCtoO/c0XVM7J6WizJ5c
bjvc5U3nQByk89aQFfu1DcL6cCvAFKFyikPD6IlJI61iExhrVmVqof0WVpGYph11
DKjcEl1qPhtSkWhEFt+fJP0i35bT757Bb0fe3kh6BgENRJMARVqJX/Mk9dmw1nGn
5TbZFd24XNrm2W1sXo3rD6Aol4KtGKlPDAAvrHotfK/iHCjSOYXLNcgo7z5XuMBt
3/0BxKU4ESKsXjmZbkJaBv+Ws5EcRqTpl/4O6/t9xRp4iMm4K0KXCzVE/U7JejsZ
21L0huP91IIy2uysriaig2DnZNNtUIiEV5QSVvr9LfTGBA+a5vj7oOHUOsBuknDZ
X2e9M/NGY7DE8DNS2Z9jtvYuvCFYcisud84Rj+VaLcbhh/mH1aW8MrcvNWI+5pgu
RLGDamE+xQQ2YZMnKL4IFZDZaIW3tmjTLFL3Pq9syhcar/ARcBfhI8y7EDzqxBBr
9qkXiv7mQwQxPo3fFlwJ51BEnl2Ll41McbJ3jz2ttTq02JasHBjCA4x3EWHXzzgz
n+9HeuQHe0ntTPyy+Ofqy74y1L53hXnhQH8YPgtNoLc6vWnNkmO+W0qlW2ad+0Uo
GXiUuURuB+YiOVNoRdcNk3/FIZ72dZLYqgaqWAorLu0xIpyL4nclePZ7CWwSjq5s
f9AVbZn8mlZyet5FDk1RxuNvwRYYs3aKJjDaviy8+3V5w6+kFVzUpUsRgP+KIW1G
x4JEuSZT7YgMEPBjSjVrOiUnBiGQ+xzQBuE7JtSYhc/V2LAJNUjIboLrkizn45jB
BXKK/XTTWz/xoSzpXqdqHhIz6zLc5lcaOgYOKXq2lrL9NVFMezH4lm85G8i/hyxh
LCWVorBmmDAAc512znPhwekHE3oLaOJpHc2mBubLWNvFVfqPt/8unJe9NPZEwGmB
pJAy//LMt7DskjpCAWmS0kCzmaTBowzLlDH4Xp8LZTraAdNIdG5C0OUCbRFGEwbm
vZRVAz+R96CzV1pr0MUQ+c0uAkeXeVQkIhhp1OUnZEng9j6K7RwZSCGz0O31cOE1
w03KYjWeLb9yvIVsUEDBKKqKWgPOfw9je+sKa9zYteDf/zj5rhJKvDVzhn8puBMG
8nwpgFho1z5Kp9IpCafSQPwSHvoIDiCpGoUAJvOdL8TlK1Ba/EBtrNmooUSjcjCY
jQVK0iIk9W+oGTzoXOKVC50Tc9jngIAePL4p8ORLKWA9gnlR1oR/8c0HLctPXCgD
nJuUXr/Sd7ExOMn8p+l7Lhz3RiEv4/oLiUnPfvJyevtx68RT8HLNKbBNO2SXnVav
/OIQD2HRElpXG5zjN2cKe/nClJYN4tRX8F19QXxYWYOXjqJIzj58/vtGpvqto7mE
fTOyiudDBZblQpVwZBE/zAfVx6bCEb9tift5cDkXuPBgV8M7Jb0kYHPaksfN51Rp
a64mKVCdtoaiBl55vrBnd+dMcE+M1LGpOhYbQpf+K/bMQtD4hi/QdmDjy4vg5LBu
hivaaZh3p7bgDFPS4/MZU1szQVkWIqoV2ShlOpQh0ndX3e+cIvhrEBk61O2s9aP3
n55VjeLcDLyQIu6mWVeReo9N12xUdLM6EFVNvaX8ph4qvx/igk831EB1VP/iEwuM
i7/ogyHCGUGsDyJaH8QafKJAl/zcHEXMmaRcx+atl5aAI0p45wgbGaSGz2JBQ7+5
HlCNGb90QwK6W1JBwhgWLCK81qYKFPXtJj2ONc73LvKl9qO2oHQxwPmCjRcymoRI
pSkvNOIp6lna2u3xKYaawHOMLP8o/tG7JLK863E11AHEzVW5qTm62M7DWPZWc8gH
0BBcYlDPAEF53mdjCIc4eHxSy4+wBdjUtwHIWw11c69qkA0Rp78sH+Qtwn308CD1
uiofdqwKErdwe+tu9bUCKNp3dIH45AziC5tITP0vm+3K7xozi5YX4qoSgnixYY5r
kFEhhlHOFBJsb8FV0uwmGuK8ClSgmiHfVKmWKOpDggLrKD/HKKQRrDc2yC93Z9Ds
VwGg6NOtz6sBq2kji8aY6N4mpqdTq2QgJHEJeHQ5aWFcxvyCbpvB7BEPhvDV3oRE
OokCkSUtuoOK9rfqnQenqzcn5nfoTHaS4vS7MJYyTAUimwVHQvRZKAp476A6hSkF
I9g/JAHL3O/MI+wOQaUbgnVZjmgWmTUMVr5BgpwWGpvUHVr3aRCtlTmqgH2vNNnf
BawdoLI+GJ891fWnwxwsAkbB+4TgiBA3+heBJRw8Z0Q82XuSbUFJeHpY05vVsR6d
nhUKjX+C9yseK/mmEAYnsnvxQtgBf8Wwa0uMlUijdFucuVb9G8b6fdyPJXQr0iDQ
Ku/bJn5wQ/FNNMzjh1TD9p25+b3ji7x9UrtfMvGvwQcMp8ys7XqG5kXPTHQYSDxy
bsL7EMEW2kV8xkrOjwbvWgaArdtCxwdR8AWZJsP7tXXWadBRdfc6peUhHpMLz4oX
hYM2F4sE3fguTFqH6hJ6KpttF0SY49ksnBdmwJsFIZno/eGqhmOI937PZiWVbZTm
mV+vLPYTBTl3e9UQ64qL8nAZODwLPuMRfYkngG5gKvJYPRlQ8nyEX2sN4Nn//eO+
MAmsw1xE3Vv6pQ3kelhoKALIjQAPn0gLlNm2EbBWs2JeLMjxp3cawDR6zNuI10hV
Q/FoEUA/h47GNflgWWIA+FMNQauXuihECJvUyco0bRyoVF+682pb1FERnIKfUNJD
wW505M9jIE0CJhAEJv5jIuxgLInLIUt7PFSUbkd1uERFxAnzpGoRbRDTqOFiBn9s
WoHSdxxNP6+5Wc3gLxd+sKHocCaiuz+L/DpUWkWZfcWSsXy/IyBBY80bTAuQ0WxH
5btViEWLMBKrP/f+dBHTfBGURU53PpmXQWpJuj1192UNrBnpF3mOMU+8UaOF3zdL
DgLDblWKnagcqhKewsJXwLljQVG0epCG0ZDMzAnYaIxjaWO15RJwF1omKmWKQ5Ai
J/LFrOaG9FxsWSNhVZ07fAQrm3bCktInmZrHnQqj8iUp8I9PuZw/Mi1IMch1gMNP
ozluml9nLYQuuuv5Ppmci8V1aJMPFNteDRXROawUUV34x4oezrEVeeI/qn88Hchl
qAlRnNMMAMoA54D82NDuQHueO/OE1sDmzdy/lWCaKA6kb4RohjRPe4X9ZqJ4BuoN
Lv60dS8PzOIdEI+SATZKphl6Q85VrVCMp4cXusASDOtv/mCsPiVWGc6GeiIPqbkr
WKpfQyhuwmzzaCekV+732EvTdl5Nh7E+HG7Jzovq6rmmCTw+OqRC/PWVA7hDF7Ih
VO5N0UanyY5QhWaXR5HCw6p7ZIAUaDGaBxOuiAJpKUNt11tZTq3vZ3+d7bPPa9+l
WS1LcpaxoOqrGjYsC5t4qNBXc5m07j9ydKz7EqG+EYemZSeEe0iG+aUCjvpz+9hH
zfCSXLzMb/d1FP1nM/StFqmXA8fYK83LvuvegnSF5jprcRSqyzJNdjh85Jn9fAwV
4WtLgLZ4wT1sKrVhmbtl3oKf45pu5WtqHWVlOJbUaVbC8hrxWcxvUawUen/2peyN
B5FnNrhvLkwxPfyosgFJvK7M5jwqnW2en11hkLidgC3vzbaH4NtOIreBQmupMHVF
iCnQpkf4nsClg8box8sxeWCYsvX6iPJXm2VGt7g2z7b05dp9/98VuI15/QbljNRi
r023uYshl+VMOQtioD3vkjGvAbaR6XtRNvF5Kn0X6cdGNQo5s34up5LAlAyQ3ufT
ZOlaYiGWn5MTHOmlHjGvFOtjErtKb9cvQkaWkuPYNLAh7PoNC1mSEufRYkyiib1m
CqkT5f5W/p3qIdJai7/GLRc2xxgEBDG+l46koXES7AL2sA7YFgyG+ZgdQPq+mDm3
9EzjjJklK2L0obVIuuI33rLTwdYUU23YycGEDl+I+qIjEpzLNIBCubNwxND6CiRv
hCnlirmb5hHpKXy56jQ9CdX6ZUUGP0N/kALUhM3o8cdTE0+0FQmQrJDXXswVSs5f
BAOoSKec15qSi0bIw4LvohLwd/PnWS+zilplheAihDyFx9dxQslR2UzeEtdIutbB
ZrV3IN2YIqkyZm6ijSlfw38uw10/nqyyI1DzlPP9oZur8xv32l+FKlzXISwYAxVs
01dxNg5jmEb5qQfOgNy4TD/81wP36YVEB+dvs7q0nVz7XBQ6wsvQ9e9RFrywCLbN
h7XmmMPan8sw5+bOIhKtIB3EC+hrmW0CPQaR1QrQxIfle0zpP1cJHkh5cniQxS9U
m0AviCJium7OnXVavjXV49O1M74M3zSaRUcsyEEM4chXC7mCrN0G9IJB7ENuryLR
2tI3ylr1T7x1IIzhp073ofnJD4qN9p+skXiCrjD7Xvm8KqUe0vLYEah+RkLWs3+Q
6SP+HlXKBaIlzCFW14U7omlUZa/OVeYXB4jz1oz8TAsfMpc3hJ4V7gMCZ7jfUjbD
FFUCuFNYm1gIDC7Wx9E+YTJO5I6yCwoi+aifBWkFGwpB9sJ91CHiVjltXP9UbqCz
gml1nBnjGWLywVhCO4DgDI1s2Xrh109+RRIKO6QGQIOcD1dulYpFxNpSJM/KOOSB
4cmkIAiTnqiwExoCgCRNlWOo82a8QYoxZQmSiwepraIEWupUxCJXkXj7l95TKZsS
0c/m2ihTey3kmkItW+SIbPaK4EaQ0QkmdrsImrxK6VImDys86+btu+VIDkmPVU8G
I1OP7d6t5FKsd4inTgAaAZ6chirsuDdYbiZyuJK36WJGp2xomAMgomjJ0C1BnB36
M4CBikRd64qJHSKmeFbS+NpLvwbnL858AYZZhEdbyCotZ7uIIcL762niWF7bGs4C
lAgforUFXILuiJGcLI2yuFfjYQabXfwDLS+r5NzvEFKwiWiOmgq+7maXYEy+6gkM
DhPnyZbhYU9lTLmNGxydEeSvUAfWSWE084LxXnSVgjZ9dCAx0OPT/CxcNTF8Dt/+
VFkWZslcpSuQkN/kkM/iuSuWW3UEcsmwwSxXf8teBKaQbNRgsCbOaYhSYWXN1tNB
HNfB9M/Ybc9MMbhN60CZfiINlC1u77y/CFzC5hJOMxTy6mUxQFwcLH6/OXzH0MVE
bT9Bl8Nb7ncqTfCt64ZdCHswKcrwMR9aPL5oGmp4Go/XIOQF3tQ5Z6xPq053jPXH
gn0A66YZyixTX5yJvGtMiaPlnsBXT/wvL6oxYp+wovgF0rzL/mOc/ZqzQ5WFytY6
nVuNp4egHgNg4gn3NU++aczCOf6F7o5lf7xIuxXcg5gJ8+RDOFl5mQL5zL8CLi5w
UdePe6PkahvJYSHlvK04gbNBOPjLIQB55uF2E410h6m/EoneIQznJLNIzH9nTIVv
paEpmpU8nsr0EpCjYZEOCVkGgBq1ka7K87ocPDJJ3wlzHQjiUGx5rc7hrmOV7aVS
KoJtogtpExVGYEDhouqcRC752A5IbqGN9QXO/dt/5B5rbUubt+KUp31GuQidI9vZ
EO1HNFjBzPQ62VlTUV4CAaDbb35N7sTV7O3xq40OnbSxP9R/uqmvnZmplZGyTyAw
G3DMxwuyyJlr0yEfh5zoK3XgrxUhPr6FS/vCEwK2Se07/i6lePvzN8tchuwCV8WS
4kA10eBZc+ExA8AGkOc9cGjdW2Bw9cneaLz1qUB2AKrILvpeYxUse9GIEzjI1so2
loV8q9lLE6wY7zj3Hof9/DbbuB4iH2cf4SC2d5Slirw8PM1F9PFxsfhPql5eVhiR
lptvn9KOLSj7b5RJNtFiD79e4yqguu3reVwP4kznD/J9RfxGEBM9K1cpzO23jEVC
eFE2Efz+mrh3f0jWxtXHVUjrti2KX2QTOF+mB3WoaE+/Zb7W+6eWce36aI+uAXDS
yVr8XTIpZiZL0U9TYqs3X2EFcTKUERXTTB2XBoRu43faTxGnDS0M/FAqg05qm/gV
1kVAJFI21+SvHNgzWbeMWZGuoIGKz/jco4deAJ2VRHIb9N6q42af8PEZyYR/TQ5J
lhoKDSqaU3P4T9KLzvw73Gti/84v6qBGZUKDqHRwUAHxrUwGb9c7kx6331qO0Mke
MkBP9OAoTpVyQZ2e7u9y4L2vSC/Fk6kI92ygedakKH2DCtaIV9izCDbfQt82gSFQ
u4+QoAaTIauMxnGlN0/OwCdGScXnbmSAu7KRJIfC5RdXL7Q1LHbtjkiFNcDvl06H
uPvlV9tQY8ytgVrFhj/EXcEfE1SptM1aHN4/ZMWiDvH1hLjmZygmdDaU0o/40NBl
ujpPsAheOoofONGoem3AMic3dXXMEgcbcC+nkI3jjJJ8uTJRCG0FaQ/9/Ipwpvm6
mlSu+XFOnTR8rofAD7Qn7San7NJgC+u74XVc4sradPTR5bsdn/7KKBDrKOyy9rYy
P9yM3f1pGF1PlLQ96628P/pW/Zr+K20ooXKQ7fEBJYOBpYluMOUs5vdtoiMdcRG4
B5O+FMuPnrDi0nu0BJ9ym+dsVLqEl3iQCrTDmHPbtOZG78e53vZzU0KT2J2yDY14
q1bsCa9FUajpFm7/3UfgJ4NxTrpQWh1aWSreaJbWZePlI25ppqYCdlKCI5pjSD+Z
NHRQTLBgRtYyjdVeVJDkPYiGtF4TH/YzGtWlU0ePrEwd6gDgrKc1l0pIp+KriQ4g
AETxnfk1NKr5FWPl4iiT3tTiJUu36qyr5RA31oS9sWSnNBkcZd9Zmg/D5PdudHRQ
vllPazLZRh5fIfrkfD2jbZKyKXnSngkZRGYrCtbucvhM2JNWF10cdI5fJVrf1+zv
JtmYOHlwxZJPfsU6vsTva5o24qgdN1sldWWPi8DNPqZg4ZciZcn/8jIT0EoaLD5H
Av993VNJ1TNyy6xVOQ5iTetLrwhr6JGax8q6M+tZgWd9XOQ5rLhwpV8f8xSqzaRn
+e+0wgp30HchBvjGHMduI7Yv0FxnCqZ/tymrZT0cc0HE2XSN/ljxhJutknP0AwTy
KuW2d9uvWMpFYBd7iAvXhkBt2er4khAhytPhaG52ZW0NZ4jkm5mxPusOc1/772SV
Cz65fDfLYq2HwF1WKhHcw6GHEKUCPIrskFm4aqt6yHa6yxihDifyGqtgcxULnMr1
7lEIE4om/ez+sMmSBigdouLyALQeK4X2nY1LnxMy1iePYV1NfGB9eWpLDk8n+M2/
3hdBJiqxESyOcCTSNWlBl/sqyQXzik4Jd8/gqSz1GFTNlCnNFQPzoK7yyvxEHDyR
ynGX8nYvsAFOlrGVNUi6WmdSPT2igGBGLseSc1JBHWbWtN1AtKD7jafu/DVxs7TE
/FsfBIQHyiQMQh1IdwPir9wWy20kvCIXe6e0o+bt2E0egfFZw46VmAwAcKq+sBG+
N2zmszgUiBMNN8cg0C7y0twuqcdRw4q8Krk5HeZQOwm7NEQWy1K4ffQO8HC4Y+I7
wxCl0QP92KXYD7lf8LDhX5ak17qqZYdEVJ04SYGCAPf71iWUT/zDA9LxSsm3Leo2
1lR0g/uN39Ll4GJmX7uZW/PskVUigNk47FCc/x4N8Q8KP6PY8DKW0gqof06V8+TM
Q31zKQPPcluem9Z79/xg9v+hGNohWhtOFA3nRsy9cTuDP+Cyn1HVIREWqikeNEM+
oSssnmMQtwaufqXHEwCaEgMlqEFeZmef/Qb0KCqtEy0AU00oBgZXKDNdCaLyVk4I
QsvraBkHThetIYRhQCtdJqYE66HhoFnC7LlFprVagBtY9AfZZzRHCxt/0gHb3pgI
k4CixqqLcC+CBQ9Ru6f7jW7NMOhnr2LXilk5m9NyI2UZN199AgHwpURZLp4lXRpH
SQrfsoJpXqHMoU92K203aOayKH5T5bzSrvZXzE0H2dKHiquWv31po4YdqKBIqCLO
rPJrAeGmQSyFbUWuJZPgAPCkKDPzG0UWEEhxMuvzSWZf0kT39/pZHZVJ+UOzZhSi
xXdAp60/KGYo3pW4I/3SPQFq1Da1Wpyd3bqDmLBNOvKEmS2NmujNFR6zbwz0ysY0
syzO7KrQuB2myqWKfTbRgIcPLvsPw112pil1O4i0u3GoyXGGwHrBVRdsQolNhIik
JyQ3HTTwF2TobX4EuAV/GiYx2UVKBf7EfKTHq8Doia/G0TK6Eel1xlMYOPXeDpFc
MO6aJQIcscsaN0Q8LLx7qsXN8VfGLqYGe3sIjMxHlwctRBKJ4iBek+fVtXkYqrl8
5hAXhLgNsl6xSn4V5q/om780wi+o15gJAkBzRErdzYw3tYsWcWSsZ9UQZYi3eb1s
LMCYu1ZY3YC3KP1J4U0UDRu02r0T5trJvF8atISLGKicWt49praKUpQqeLDzN9Qx
LH4Bm7TcxYJ28dgBs4X0WuT5Uzv2CLRm0z1Ob8c6lkb01a9HQdbpag85tucMqU8f
zlFqURodUJlflu052JguJt5xafjzgj4t64pfzeYYyjDTyvca0zTvh8vqXUfYhjbC
mY39jHufEDBDw/sL2TgZ1Pi9HERk+x2nvR5lMD+B1DhmzgeOO3HXpgR8s6bxKCtg
tEipxvYA1P1ynpZha3zlkp8sVEfWlsnM24WSPzMN/ACZT/2J9pTwBQiXXYTeDrC2
fnbBQHLmnkAGpYl7XD/gs3lDe2Pqkrwr3vz76HJW2gK1f5ipVuX1JXBmCcivzsUH
1/UwKf54iQNDyoR4HwxjrZAod6lpF13maCiVU7QQBiBH0VR/NGJE4Fnfzhdyw31H
p9NByi4ezegS7ZqM1GBF7kbzG/hxz5GYsXv44vwNn1TRUqsqy8In9H8WH1TbUlh+
ufDOMejSeIq0wXQLRex3MK5dSKkgq4FBVcR/3+LpnojLmWb80NzB36ksOoLPIHFM
pgd/d5BDTE9ZqxMZmcst0bZRKYwXC3+cF/R5aimBOh++UclMS6KovtC9p9NUtq79
UN+5I5o0dZSK1ZqmE4CqS4Oce3J3BYdGBA0eT821rMtcvd2w6NyU3ovhAZEzWZTq
FRb/YeHHT7P+ZswRRiNL2M7DpoQVQk0cSXlgM6uVcDMgZdiAqS4cCak3PFo1uT8b
7wrpLqyWU5pZIy2tP8/V1cEtDoXKYNgK3AvQLnJv1j25KqCudP9eTzyYgLFzlnfr
aSbyc4Ghd6zLkXwsTb7kEmCI6wqny7OUFQ2QGIhT9QRadGF7XRdryjY7S/YpO+F8
3RPZxM1P789Y7BunN2L5sfxJsYXfkpOYCL6o2vGiwdI7ehsewg+IoNivf/XKogi0
32DKUbEL2GDdCk72UikJkCGEaBKAqaWuxP/GSm+N59Cc9+u44Roxe/qk6bjeONT/
qbixETuLPbh01qBh9FLFCwED1yzWJJ5ZyOJireaV7cGlljjECQ3gqvm3JSq1zoj4
8UDeEG0aKFPnKr9IvXpNqvLyT25w4ZmVN/oXAPzIIRXsl5gQGGUl8cHlGkM5AvRL
U7+/oJvzeyaw9ztcQFbsVNvKbBXiGfJikEVMMXMNPRsLYPGs9L2Q7Qy0FVcf9tDd
PXmOdgqrVG+YvRxTK2aiaJk8zwxb025ezKg18P+v45E8kvZbN2SH5L8PLBU4+JqS
C6vpEgzqRM+sKm5EUyIY5IvCRuI5TT2tgB9BBXXEZ0aKTtP6wRXU/C+IDe7JCb4V
xSQ12bzyaI+0zB0si8eOmZIUQYpqU+T2WpXXdFjkqt2no52C9YbCvgXXjtpntdNz
Pk+Q70leWGw9XoTk3fJ5VZRhpLUF3bNVaRoOw4cgnnVTY4fYSH4c5fW+q6Hz9k1i
N4827/b4t0YnrRGjSo2m5upFHq5hHzfW4rhc2Ng5d9CMsH/2bKB/MrJwdP6OpJKE
s8N1o9a0PVzD+w4eK9Qhoi9buexxwego2Q1Dbujo1aLKHJE+9blIKhdSRCtrFAaw
Dmbno0dfdbyGDy2to0dSJmxD8wTg14RJXihISeBDb32BlQ5BbFJVp3bt/I0rrqak
EkpIUNT+T/RzUFPNkm+eVMkAO6116zx4vvGnTuKCuTGPjqDy4cp/KGG7Dj1dgQlX
PJ+d1FEyKgqrq3iiLjXgA5CgHPWAsRrVYK7MtH9brgRWp151yo/IjhJJJ3hMNYPo
srI4ZxYafGQ7lJHccqxvqmJ1b2sywD9nqtqeqALBTiNiarWgg5PGInM/rDKjcmY7
qGq4WP+FZovsfiVuD21QuQ3XQmdoMgBYDGF3Z0yrPmviomzWYucsf0t4Wq/9HeQ6
TzGp8QCUDytHHy3ydY803fqqtEvQkeuuCL2vn+nizrN57MBru/Qf5M2BTBZwiL/O
EY2aVuMEEE/lXq2yr0kvwy/OvDPPa+LqImMpkkTnbcd2dtpKDRUKX5pMxIV0KqCJ
znCTG88kNf0i7zWze0imL5/DUL2aDCxU4k1rv448x/tX56uAA8Ds42sam5gmvjHH
5x27UqhW+ugU5LiBKEWqb8WxPeOGgSRbF0Ul8QgB58Zwkv1oOb6lHsymseU9V9jn
um7zFH8ADBikI2vUE/DD0pIjnSGJXKyU03tOKhGHF4B7Drf8726I6S5H2WZyhanP
2aZK04k0jctrwC2Rk0JxUpQ6LHBhcvQKCVwn4eIyfRCFj7l1xPwOzK2aM8z937uy
hTj/El48l9ZTkxQeiWKWC3ZGa0+sOlsJRtvYO6TY/NqGhx549WI8qMg7QG9qrN32
pjicZB0UhDxW42fBgpSKL0BXb1NDAaqyCPX+OHoF2/2YklqMYTsU9uUx6L8fB7YC
WVD6wC3nf0UUjYjfYIHmBoxANKjzClgUOPFo7rfOg7Jy1hsBOppRMyzHRsS4v0VM
GuQwBQA9PVCUjXD9zdLUxi2yLUA0LMzkf/4Lojoyh+dzMWXoe03UWd4Z1eXfWbyR
D4Pc6x/k2rsNM/RlL9QzZEfQJdXeNcGTjJROCxe/BRz85ICGKNZUFDKcvcuDPRXC
6/vcHkCAOAQgIZf8bV32gA+dam4ULybdoQxmLMmLKRGG0dUcfTTTUH2balygmejx
rJhFdvtt5xVl07H48EnOgJQGe5MeY73vu6Nqq7V4LzeUPXJYq35Xo6NEIQCZWdNq
OZWgXd7UTTwQxzlzEJkBunD0JyOxMZruyx3JiiT1VeFy/ynFMjSc7wkqnhMa6hAI
8olrz4ww9/Xi2t0yziLNR7Ufl4ldmokOwC8fDjdm5UdVE7qnVfwyMk1FgkOZayK8
Ffc/BlPUjT1K2UOp9d8JPFLSl4ZuriYFqRBVRzcqI89AQe0dbFZwJXPpdD8fRPWg
v3X/Sns0Pd1ISHm9Xz3abRu2KfjQ88XZBLvvUIk/e/FP9xEXoaG+tlrricpXeCEo
iPSqxf/KI+TbnglqGpYn6WDEtnK7QDoq0+oDj3gG+HKPDoYrM5Z6alloQ+tB0k3I
UyGA42/04VpftmM3DCkmPgiAXLJoq73FOhXN0bGZwTRWPiISUb7C0wPfPbLiM64v
pakvuxjoLS4jjfAv3AWMZdYhOD7pMIBJWOMpmQlsAEkSzVqIv3sMecC7lNaxksW0
eynzyr7Ktav9HblbIujnOaaUxofjO1YGSY6cVvH0O2DmYXzFVhrBzmqQA1Oi6Ih3
1M4+szVp0ISRNg+BItXPHq2h+me36FUgAnq4M49IY9a22HYhQHaO8S/bWS+ZpFeJ
mjrGwTTcQtLICYjuS58u5xZkNWXeDh4WDq4Qc31vnXLUd3f7YYYzQj8ClqFUTLq3
d0JJGLN4zj85uwy01UxJVOdHCNSPR/vThVX0X0HBmvKhjNQNoO2eSMUQEcHNr5JG
R4MNX3hny9hVcBPgIWVrJsac832JIXvu9vvGsLny9dC0UIC08xdyz4QsqtZBRlAk
wQPJjENXGbMQVABm4Ggc0IxSYII48uGWqiYCzWDbdG/3DsMaZRZSBGayLF2UPvY+
/fUXNpPw9iOkBlvjmDsOrE2l8Adf6bkQ9Ot0NIPSxL+aP0Azpr6/YIDr7gej4kc8
lGIenWolIZrcVD5kOJ49SX2C1zhGW1blWCLZUUo6Abr6YXlgZtnqbhtGJXx2kbkO
6xVlaoRqLTC6Vy7noDc6Gz0wOiz6d6t3IEZ6GTvXzllCQcCEhgjjvKlsbg+i/fj7
I51eZLoHjRUGe32bfwROn7Tar2RxYhJcksXbehalBOoIrJnh+xjXvLJPO+MiCwtW
XMP+TtpyJ026u07av3UnJkDC7dO6ZQNPP53DU60/hlVHMObIAZXfrIkwLMr7k3dt
JT8XAIN0OpsUMHbkuf3P5tZySQtVK7HshgSM3Bz7ook+MvVvM5wJvg614bq13aAa
bntg8YnVkTCR1/cf85lUyWFI/XU0HfH2xKwBtF4Icvr711yjeU10QfwQuVfVtKPv
6BaClZKnCFRAdNbhBALNdLQDnspeFIWrt6JFdmuiib9qR7SKn8WqZ0+MvBzuCBus
ov81b4b00nC6xFoz1T1etgalyrZXXnP5bJZ5X9MBZw9FGair8yjn8rHt6XmSKiBJ
raOKbbJejE5imisJaOxd3ftptOLeHDn8TO+3eJj7Ndtzm5TvajmbonI+8pwZhCMe
aMGRwphft5L4A5mG/QLi+CURcOQCOJmSIq2bQoReQ9VoVV1OtWXzrxEOzFC29jiW
zRcye6+RYe0dStBGCS3/c1EdwRmkvaqgYMCEL8zI8etN00rinFDbUHMbclqzHJo/
A+AfydXWlL2XzuUYakn24biExBLWUs15NC0w+cLYdMI=
`protect END_PROTECTED
