`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VVSQ5EFht1dAKOeXaVcw62xOLLvSeOgpJOeVodDG2qSw8DajtlkErM1dJNuSWCq
OES4g33d9XddUKph+WxkY12fRrty/FR8rKsswyrdDFeSRdBTitFqdQxhhptQ8JtV
+VaZTnGc0JdIAs+/OLSSZWMnjp7HtF8vW9IGe+dAuh32eDzjJ+az8kSCulItPpdL
B7Q5xlh9dJV2IUjzuw53m032kNqHPMIJFRB0hquzd6vqWqeFsxVLD/14YphFNj04
SVwz8nBTuECQ3ZVQL3x70ZkROeIlV0tiy+VClhVd8i0FzaZOPe1Up3PMkwWyYKjN
pu4vlALPnkEJWJ/25CRz7Rj2rjFUuRT9p3mPxknxkz7pQs3GgvOJf4OOQHyoara7
T92bUyFFb9ssDdAUnMJ6ycgxlep1EDiU/LzKwWI1qWT8zKj/BfjkwE5fKaXMZwbB
rHC0hnCiueWct7xRdzBZZUmQ1rJ7uHJSSMwmS0FOHahDfDO+/qrep1LeM5b9FDzS
FAEoLDX0hyuk7Tyiz1D1XAlWQanS03pcZZFWcZSyFZuqL7zBuvg8IEv+5gXgZ9fK
ZjzC53+2KnPIJ+a5lFJ/ikpw/58/EPL4t7DxvreixXpfyAo6JCRH/oQZjeMLH40F
C1hx5WdIwslwYa/hyEsjDP6v+XhNNL1pVZEMWHLXO8S3/PGenlGAeO+f5CdyPxJU
Zo6XhPpDl83psP+KgW7nv/6CheAqc6iS56k6qor3pYyKlqd0UfZj3ACoQAuVEURb
BN/tR9e4Ci100rrF+frgM/0vpV7nsvXT2sZyN0vxVo/Jns9ms/HGF/y/ZCHv0Q3S
3dXYb7qodjDGKil7xTacHhyXY2QDHKey8MU1DZSYq0jh/Y8kJNf4svwseUfOwsGo
CxsIeZ2dRvNAUgD+JiRAc4jmiLEkUqc1toLqAwZqar9iFXnloAqUookMIVQTpsPx
ievUNYfoDpJf/yR77sl1lEUrgrOwZjFKgoLnOukqxAqYcKp87V64BVK9HkZ6JtU0
g/q3TIo5kbS3u5X12Tnbj4LqSIKCJc97s/CHWstuYpkjIhwC9JaCp+jSiH3Vk2Iq
`protect END_PROTECTED
