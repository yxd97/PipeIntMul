`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6u3nLlJ5H/2E7McCsqerWtBGGEJVTbSkcQazFQfd/SRB/R6uOXtrI9W/eiloWIL8
VkY6krhVWBFCuf2luDGxZzJkj9kvYKHmZXMaJ0cYt4OzH9NHx7kZ+RbuMgBbZ2S1
PGtJRiRUTFjjQy+Z87xHnKlZ6RTRDwzO3bT45RcLhTfcaDnwB3B/YxJ0wZ964k+Y
j9hHUch6xz7eNJuuj7521o0BZwlYe2yQxxd8Or7qmXvdGN2rMdvpSxVQNZEu90aZ
SfaP6gUCeQS4XakEEP+88Jb7MdiGD0JOZrEzOQqDnO6hpAd4kvMBdybzC0Bp1/rM
7xdF4CD1p8WD1XgC9JsSfBn1K/gVHSAwYU5ddx8J3Qs/aJNpnS8mV99Xvy6uIFCv
nIf4vIXxCfhxce4GrKL91Yhe6Srq4jkXjEC3tID1I3+Vwj/kwwZif7RhDYHMw6z8
I6S8TIdwSu6UJhadUq7vmx1+RfaBD57EvzFiNKErqnRa2hle/4j0YDJTTbm5tXhF
`protect END_PROTECTED
