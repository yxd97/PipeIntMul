`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDRyl5GqDbL05Zgm2W49kgJcoruy0V5FzfSKcsx95WkOzFVt3MJC5uiM03tkfFrk
guzuL8qQjZzDEXUveTm+RrlVoFOIfhQeL7XtONtfTscTOe8yPhzgDNtcdcpt6rIB
Fceg7c5enXrFJGJ0MEeRHJAE3ajxU3U7m1qvWtaVkp6pBj36FM6CtTj7gYE19bbt
v2DZgy1Il/JzTDIEAkySHU0pczBkm9OeGs+TYdTpqE/rCjVH1thHHxaBFXYkyq3J
jOi2MEB74M8wBjKJurGlAd/hchoGc3lexocOTzSogIMa56LyPcxiGn5zy12HT+sX
VbKW2KqftA8CjO7OaJ0HhhSfZwobLGytUaCBbghPhAyUekD4RJPFaj4M+faN0qz/
Z/i/cFe+tm/Bu7GKtN9jbliebgSJrEyschls+ILkaiWcd0hVpkyDycY5Xgqf5sop
aWh7hj2v5gZ1fVYskh1RL8h1R19QAthwMtCzJSouWqg7+pPbHak4NIHb7BaQ9rcF
oEnSss+0LD8VqQ6PaMontgdsrxR1Jkfp47V3vVFTSzefNgBC08FFe/B+zUb+Uhcc
DVohEQjnkAv8b/YhTcS1+Qr1jPGHwqx5+mZbUcqeGGTR9+Cr0zFdX2EifU0+8zDa
oLwSWNn7yALk5272aKAV1SZ6R2Yi1ba9xmyFIDGJz78=
`protect END_PROTECTED
