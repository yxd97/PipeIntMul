`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LCMzogXBsZ+tHJP9q1YsfTHRNZtKvm3JM3hY9zv8vSeEy/4BsLFp5HBq84CTB+r8
0fSYz1iPife3lGYpwPgEHN4lLbTgivqouvci51eEfg969URpTYJVK9XnZkKa3Nau
Faac3+aZCv0olJG+Wclxjq2x3dsEla8E6YBLGoqFD6WvtzHNSp79F+9Zvgx9L1ab
3pf1jqA5F2Q1IALvAOmttudfjyZVQhDJw1IvexCLICApMlfktcKi28j37mWIqb1x
zc+dbXlVI7QFgeV/yyMBPapWq+rc44witeBPYdT60G1oxwmtibS1HE3ou/zblL3H
tgGRR2Mn6BR7JWKdSejq4Gaw57OkrbvOa63o0JPf8M+Sduw8asLIB1FZVEX6juiO
FIcDOZRFTGOZsUMK7JHEnQhuNJSmrcAms9mqM5UWQrgaKr8IUPHfSOgayqDj0U4z
JmkJ275Zw71C2OCpngioL451JT1lYEwZ5FgPD+1a/VwtiLmPT2sTfMg71HHO9TOc
VWf/V3OOBzrVT20srUOJI+uwiWRMKOaF/QAWh3YO0AFntYDCtkrRjOhhvMuwjyMb
yLBPsIKuLq0AnER/qh4BZ3qxFMBcxtHTh0L0YseWkfmb/uCRzEXBFXHN4rCoDPaT
OPcdhPv9UDG26yhClnW8NlerWPyqVGWtbI5DvVsusUHfeAZRJB/QpFQMYDobKApX
IS46zCfkxbwH5nBKwlbcyfykAEAy3YFDqeI96HHQN8onKklLMW+H385NbFFCh3e9
fGTPZ0PREoA0YqKCTfCJWmtlvDRPDiJ7gFNElnykylGw0OvpppCNvF0OhQ/imMCh
rnW4R7T8P/DLHG5im1Pbd/y3xhbMM+IIWyclajBQ6xTE9hP7qxwz4WxmSfd66sZx
bykrooexFIRgjiiHKd80z2yjPoyRMgRSu6d0yXe2/TjSlMBVDEK/4c57zG4Db+x/
`protect END_PROTECTED
