`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0jzrOx1ALRfyx+mW6IzjihuX3G/9DJb9u3xdNEb1rLlGgN39gIY3GZS6ZrfXzFR
buVU8YjqPrJ0Aw5z+Tzmminf06GvJpSd03nLNqP/Rqhrtp2Mp63yuDWh3jdu8ldc
R4YFeZI4dfzYhZUWgVH/0LecTCTic1eDhlMXcQv0Nmn1NFbbLgvnfsal5W4HG6K7
OF5uzPVWj4uWHS1cmewUssp4UXIx4umyK+xJQX3Im5KNsNru/AOY39UeKTSi01zU
ZbRy7VWhSKM5JGfCICEu4NiVK9CACL6jP9uob1mm8nIcXJ/kJW30p1tGHmkjbbz8
vHSooTqxMkLERZ6BCpxvjw3K2UAp2OyELKwFsE9W7M39waMkuEoirgq2BhsMfJQH
ADJEg5Yn2WVepLJSjE0mZur3WVCvWrdLsu5HNqDj0zfdU6zCcU/a4rTYwywd/ily
HfGCv2gGFXorqiu7tDRuKYNVvNJkVdAx8gisOP6unhbkJJPz+IjHkWGjuFr1LG5t
cM2hkOzJYvwb5CQ3TGKT1EG9NnXh7M8OJdC0njN6JLp7RKUkywgUsEDghCm7Dwhe
LU2B2gNQSXumqfAe+sOzFvfjRjUArEcNirP9apvTQHnX2pGf+KLyc29Nz7bVPH6q
s2gN8jE3SrATcLEyFKncwJIUpC8jYDx/tlxU7TmOXSCkCf2d2kEG7D6vh8wFZUW6
SwI2c2xKTeUqt3QROSUwPt09jWw3JBV29hOP6/yh56silas7Sxrf9P+yGC4FVSB+
O1OBibfJcKHa67CvOpnjHQ==
`protect END_PROTECTED
