library verilog;
use verilog.vl_types.all;
entity TBLOCK is
end TBLOCK;
