`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yuioc6pIVPQVSVgiZTaj7Gpu7xIbzU4TOIaUgJjIbS9XLhnuI1JUybXKP2pn3gHs
IkoIPa5oZ+2WpP6fd9WMlB35dFDrm36O9WHjoWgTTvGDoZMFTMywxK7nRhmFpmZB
O6oPIXnuazBhU21rZCvGnthrI9ha3dcHIRxhiJRu+MPr0eUU57ZFjIZZyS86NJi2
yTKBaOlI+USah6+RxmmwQgqvSpkFwhKiiNnPUb6Q54Ca9dgIDWa5ofh1iuPAoLZM
JkM/tK3/ZzKj/IJ0/dnWzM1qRgzkLrfey9R8IIV24NJVM50TQpfuSOy3+K4/EJ4+
JjoKleNmuZvVHTHe2Q1Fz4E1xRgd9+FAeX455XI9uNgJbJq9jxK/G5AfndKoiy96
xVkVEOr2ecEmcGuot8HW6IZHFzXLrgsWLX/8u5sJIkhjM2TON5tGxMPsHPwqoA0P
P5uqwfD9wlo3O/vuTzvdizOzZG8ukBtQOVQNrKGkemB0QvcZqZZTfenPxPxbYpEA
kFgydMXmiLtEeOHU9cRnardazZkv2DgxV2yxU2L9uwSsGoEB7IoNZAdRHaCGMA6s
Tq1qqAY8JS2FLyWBB7NQ12c62DoByVlG6BJhpkROEfHZT3W0p8iKMEVkKQKkCd4b
KJBWAnIhhZ80R3P/GmPV2MSQ7f86AHZrYODQK62MfbGyZ8DGISJy0Tyttdbb+bHP
FkIz2LETellzIl4IsyThVTnK0BUxKoYPQ+3UuDaEp0UZdE52+MCbY8h01huIKXjK
QFYlq7sL2COgiUlDaD9WpUXascYAevFDpd00WMOQDQAF+kEQ3wBZFwtJkrMb6yR2
epe89D0Jivij3QZAkcn+KXgw2jEpZ8UlO/+eIRCbcLIm1MZLSTuyYLbWfBx+pd6n
2FgkaDN0Y8aIQTVE5FBJtS+CweJxF0C2oqjzNbEItn8zz/KfvIDxmH87FzCV9Bni
+8UTOGGbV8NoAXrv25zq1O2/VQc6FCb8hNX7mrnPlmIGze237Dn/bk0SiLTiAJ7i
W0uO8DzC5NtjzzI9qXGgn9Nk0wtXkeaWrasTRzBQHmEzjS+j0vTBJXm3/gJ0NSXv
nBkTD5ZZ2eKQN30nTXklL4h8K7gahpuBBslfaWQnEV6q+42UY8+1eVV1fx0Hc/r/
6mte9hr8CTXaDbfPWBPvvVucCtqsg+e6SdRub6YLXAJZWuCT7RmL72HmmHYS3dy1
srN2ilKo4O4WwYBNAGAahETjiZHunhnifZYfb6MTh13IQV36WWPYAOLA4yQJtf/S
yMC0+/xgbVZJPPQLfM5H4VYwnsQ4GnFudgnzsMzZ0Hj8WPbT40kk789qHjsYQaRI
2vqrbrz9FD73SrwFcNVryQPa479J7b/ikEoyndYoMeDCWt81B5kjYnScwZCyVKAH
45yatfE7b53qIV8V5dS49SByDxR/Teby4JPr5QQnyW3iYeSpwYEUkZNrp72u2KNj
u+CwvfMAEDLvSh4eC0nt2P1zIY2h4RLiZzkeOcl+vUXhwniqI8SlNtLRZDSKLxpY
67NyJtQ3iQEFXDOvTIjuwqoQec3E11TVJaunGRHCo2bOHr4gUi4ONxU+CcnERaI7
JeQMlSrJcOw4Ef3H6hlLl7PmTXpbdGa0GhWVUSgh6+6I3xNlCQOD7JY9Si5WV9AR
nm6aZ40p6tEDuLAZBrUjun1q5UJ57MpXu+o2wUO0v01xawzPKsa/0zYEk7ZizcYF
qahMJcVfYpxUjhnHGskhLtgjGhxvz+bVjqRFd4MLJ1vgmOhhDwKb+1VoSexqOxJw
WzN2+xJsoen9uWcAT/wEU4H+vW2q8LopzpSobARS4ztrH7JnGuSoGx/oS0T3a0iR
5wIsz5WL6DtPN4NcM7QJWA==
`protect END_PROTECTED
