`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K03j0qufZSJf4epMhYJkEa4uyOvPlCyiRX3acr4FrVVR3AYHvmYwaIz6st77lAMe
s2AuYpxXiinlGhjMwlmw11c7w3TEIMKhnt75/ejygsoqlxJ5AxfkmQFhgsZCGXpd
iQt2CKJ2xc3hPp0m6rI9urglW+7uZ4OntUuY3Tk3IM5I/pkGTdzZs2mnZJehA0YE
/QYRkDxdJd7waaxSj1rYMd1i6DkKIvadhFRZw4y7rn96RS0Eh9HZ1Hmk0XWmDl8k
+eKN4hs9drKMM90yegrAyihznsaB2oeRnnT5SHygPQF5M2hvjuuQ7Z/klyxQ0T8r
kIgX9rOpAAK+hFKInOXNdbNQSTs6sLTtzuIu+LpbSL4qxx96oYc0r3lJID+84xan
kGWjSnC+arlPXkTQVcfNhbTECKfOz3Re+LmE7F++4f6Vq+8kzCv4zVXxUUuXBy4l
HwBuf0OGLJdJZgRwxrVhiALJByesCeGIYJc0DBfLoIREo02ezZJLWhyEf821YIy5
oBRwTtM+KjO5WsuTuZYSCXSNMZ2etqXqrziliO6ReMvsaiSzyGByjxL2dCrVlyTR
`protect END_PROTECTED
