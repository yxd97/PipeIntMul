`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M4lu1a/c6IAiFBCL7t3rL1RXd4Mn6fLWi2UvjkwqebgYyDPwl4S14KCikAABa6Y
xX3H355onAZjIe2DEtbL9y2hw9cb1LXViybivX2vQMJjsq4ZWDvT/mZZ5zH6+OqB
5hsWuk8RcS3HcTUYbW3rBRLop7xDv3FIKndTRBfQY7BS8XSVl7X7zoAQjf4s4k+Z
hk+5JbLJGwzT6FkU7D5f8he0A63oTbbBxPY4L7zAdc77k5SbQ7p3X02fo7csNANI
Na+nGEi7Fc+Ofmh1SnApYaUs8QR9f/RMNXcJnYcKqsD7wxxyufNyM0k/xiQCO6DO
pGkLzyCplJvGKOWmhOyckbYk+ar50hHy4VRp3KFZoO259+U6SND2NQ6GAo81b2ms
PEBtC2Z9Si8/F6iTodFBJsyZrDZnyEZGpwqI7pTtLXSnbiI33/F52ubKKdl2AT8b
i38YwQJMnR+ibBotnblzcbRrXbzmnbC/R/JNmH+5ne+MYl4u5nwf1cSY3qFk/bxP
WWjePTQtIa/cwU/t/cGc1c2MaLGQ+fNCSeukna+FamTexbKoPL96C088PDQv1aFE
FuRiZ5hgQDFsWo1DCj0lcxEdbDrloePooUlQUPXWPiUncciUjeptPPVYD9N17wQS
vDpYiGkufO6ed9GJ6EezU11NkgWVV4C99MTkWzhCkU4=
`protect END_PROTECTED
