`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/FlvMUki9ImVFdrZm1EOQJ4u40xHbcpJtxOSP+AaeV338fU9SFZY1BpMl6SB0Gzb
sLL3cZpQvrRQvfUdUiO41ZgGVpuql7473fA4pM+arZ/Wjoc//9FLG1cjh/j7JRQb
0aAwvH1qLEty1Ds9UJSuVde3sRSLwVrxAj8M4GB/K/9DPzp/7tOlM18WW6AKbnRn
qeFH3YpIlvOlcHv2ndCnwjR6Rb1GA49R1NbZxn6rvRGdph0uFZUbnwhZUT/sQuDx
zd5o1Hv6lzSnHSljm6Y18O7f66UJ66WtP9i/Qow5fCwEv58/NX+6TZk+ji+roVtL
a9WIG9SYq6sRIA3yQd0U+6/L8Tb+fnJ6nz9jmo1rToBv/D8g9PXMJEtOgpCtIFoE
8mag0EOwFnincRnUIiegU1owxvKQGk/vxh2LnGhg2x5vbolFByTUuBtjIXceBsyn
+AJcawlVkac7tEYNbGHKZY12pDA1sTl+bj7PSM1YNH2leDgfRfwiBnTCsc3QTTpd
Fna6yMlr8EJpLs4BJPD8JhyuVegVdOhgrbNWXUPmShYjQTWDoP4hQ81wWIzEorEq
ik1QTsWsd1j2PaNyKd8i40Wt+Xh6xFcf0hivBZnHlGYVPYS/iKtuhrQc8pfumkUc
Up7ckEzWnwknHSK02wnEGzKvpnykO0Gbga1LPNmdkScQzZhNRBthWs0LmOJyeUDR
cx/DY4Td3je2A13cI8CLxj+jO7ucQIM3GkSCZPTiKC76ccz+nm87o5E4zoZqxplP
mPgFdqmIZ+3gzoO9qbuqZi6Fd15wk/sk5hHW3/cSArUyamWhU1mSBPH/HrjLOAc1
oldyO2jDTudjt9kgOkeeH/R1OiW+7BJfX4/lVWBXRZPRNfh3rKvmPt0QJwb1PqNV
mFn3kR/ZoY5MCWuOqJBG+13vul0MrzOOCPjPykpHh9wjhc6wPowO+fIhS8s5Irna
vt3XfnfZM7KTckiuL4btg7SJBP3gnoEj0UEhCkRArVG/RrUwnktHTq4ddTPj+aIi
HhWbttB67kG8yvNI2HU9w9ojfFNPTlwHm6W6tedDbpPMhvMIQqTshc5j2qa44Nr3
EVBD28T2pLLKXksLE6tIzXlI8n+38OLFzFN9ES+edkNVB7Mc+NJ/iDhhmBBEh978
BWWIZIgubepJLPItdTjybFmCNSZOjBE116VNrlmEpmwyxO/arUNS8tFGS1ruwwYS
3zMg+QruI8ZKk449T6ztLpzXqdD+6fR6Ec4E/S+vGcVuPFHpX6qIctaT3qqaEsK4
ErsJtIhVyAoOgbsRLjeD7sX4X9pyl+L+NYwJE0d/U3VMTxBXc3Sp6az3U0ih2KoP
OyauHqaBKsSC30a4odEA7TxwM1AalU5cUj+2rpzy0/Dgp8N0ADTA6OYVwpslS8qr
R1ztMgB/t7GWZAS/qqc/1uNxNdPWZf0oVzYMNjCzuKsEpJ9mXP8FzRoQPF8l/J96
YUtXNIPxh1qcb9bZ1ChoJFPhlX+KgwYFlAprk+fJ4MfND9TcZgTuGFetRBrS5epa
KXNt9aCsryTkq93iwIDWcVi+1rcM2EM/rxs9cq8a710DMi049fNbqzs0aWsXSIDa
H3Zos3ksmJvKjr/r5qdov/JCq6uR0t3e6C3WrV+kB5C/NS92+S6Xf4whdKSK9Fpv
33YPYDLMrnx0uUctMjWF+5NafqdS16FKhMkKillXrIBRbcH2xSRR8IGVPfJcf1VV
G2ThEyJifcvnVjEY7RfFoOfz2bRZoNDKsBbzuNI6v2Qyto7YDtMtUtTQJ2WMT1vo
qTnejrrCm1Mh1KS7oEUb5TEXNz1XsJRs2WH7uGm8Gjo=
`protect END_PROTECTED
