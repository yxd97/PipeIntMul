`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwdWVmuT4JioL6ST9cLkC5V40M/ZKWBtRY4iusCOx22GUxat7JtAmSuO98coIg8r
7UJ4cc3bGIHJ7FTJIeQqMVszxBwzlybDDrVFR1Bydfz1JRv0SOKo3n1/nOXO5/C+
LYuchxIYcKvavx7xyHJPEcsasxlj3BwCu8AtBNiNz+nwye2gjWt+hsDtSL/M+tB3
D3z20n8unMpuSLzYc/B/UaU47m7mO5znV8r5dTYmWarVkPL1cBbTAUjOgOwlEaN3
95t2NbytD2aR3wJFMXpTkR2XYVEoysHxbtDdxQQEVDG6caImgep7dBUg0gYkn3JU
z9+6Jc9Rg1Sz23dQF+gaRPIRoNAxoC/Qi6qqZZ8iiTsaF8dSNSeEvMgdcKnHUKDo
LkHX1b9GwefqFTlsfgVu91NJM8LAyOX20krUQJNCBRIwnAQ+9b1JueuBThN9hltD
`protect END_PROTECTED
