`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Ie9RM4fzsgXZOO3fhISe6s2qmuXw6lncd+oIjpdCGyjqtlhpjqvqRvFP6JBw6gv
aue9WYuud5do7Roq2JEIAXbySw7L1bt7QRv/apPNTN7pHoRNsM+Ig7KUhXY0J1Pk
Ub/ElSJkETOsri3GtI2Lab4wzBt0f5E7NEvufXjEmyZ2HPlC9CCYsqe2f5RCxy1L
XlA18QBNB3rY8BQzCYXLpYRmMFxvc24sG/a8qTqZzhXd8aO0y2zSgB95xfoGYAyu
pQ431ppgP8vZsP5R7JEYbcYPzOjTEfDJwO1VQJNPW761vU7fJ0LvsxDuh1a0xFzX
`protect END_PROTECTED
