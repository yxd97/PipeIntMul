`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qpMQAZCysMWKdlPmhb+u5k8c9DpWXFbeEEOYafi6hP4/79uNdvw4mqg3S5KP9SQo
sciG889uPfU+W/IdYmt5tid6qeoTorQ+TxMRqcZ554LN5LTLbhuOyGsm5jgEoy+0
Y2SygYS0lC/cpC8rsZEXaCkJ0ZF6hfc8INRWrC4swW7s9fx6QPvY1j2A2hDcbcJ/
ADgxm1RUTuSNBeyt85ftvMIFVNh+hgOdnxJ58TIyhA+caoy9DnMi8J1eyrI1BAKT
OXTwlOVuGA6w7aRm/CbHu8lru+Z1PEsqOC9myYPOBGRWuPSrBedG3gqmgCGmDcnv
JufC5wd+QiCzyKly/IBEBDgVkVt3a1Cs0ju83R6mK9norc8QwXRjOn4t9b33wdlE
c2tkbDXynua+S9suiD5WRAGsOOJaT7OzewYS09C67a41/rxkxO2rEAVYmk91OsGu
mB8gQfJiOBHrcj23Aw3wTUzkTf5UquYWfBozAP3HXxMuXiJ/KUfidnwaXCe/yAp6
H30+/jUpz/7Vh+fIMoT/vpTogc2zF6e4m+WVgjI/HDCsSeKESuezOT2TqWGF6EKm
ObhRukvPYEbcdUFiY0SogGnKpNGE7xdZeVPgivVohZy3s1Da9WZP5iMSntFUQUHw
A34Tm6dwJruzp93OOUnmNA==
`protect END_PROTECTED
