`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbyits7pWubrqxF7qAjDmkpCNQNIE8ALNUlu3JPBeCkVzWmwLemx8HxOD6dzfPjZ
Ul0qnK1RSP/d3IpGMr/dBvoAQrqgs+g0UVvkPmGjFTKWu0XikxwI8MAtM7PJ1Cgp
VELNjKT3PutB4R/ahVdlPhvq1px//cfuz+VoumHnFG6ww6EnCTTvJ3c7NowSJCiL
K6DVY9OMRyedYEUneN2F/qUb/TAJ98CVxg8FJ/rlmE7/RKRXLRxgHUCxwlWmSWEg
OHYlZ8Gu9D33o/BxyqdmEaRBoBcraTK/fJpSO6Jw7WHk1l5YhLuT3LQ7VIK4+j/j
UyOGVFkEsKJHgu6sqN9jQ1IPGlVu9WMA2tWF01QDSEubNr9cR+Pnyx7J0fNpI0Ul
GxH7spwZBcqACHq8tfCildfibALwQqkd7SKpba29hgRMxI+Lerc/ny06ZcxcNRsr
p00GxnEBD22zeEkRbuoUqIwHqKCx/e93LKTDgnaAcFw0CLA/thaIqEyRLntPUu5I
iUyhXiFxNHCOGO+KTFZorDCL5LszT0zl0sG4vsCrOD3YS98lp1sYrBtjJNmnbeLE
OHX7cAQpQ8dMqWWEbBH2Mg==
`protect END_PROTECTED
