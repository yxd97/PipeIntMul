`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XF+kYTbT1qffMAVQne8F9FL0hcOfGZ+ty46TcmzhJQADqGhAJHqdSJNLE8HDmJmE
+Gj0P1q0lbNGXYCV56cvlbyIj1OZUKkSg7zmgFBS/xyLOwX2A1LZ5fWtGL8QJVXd
MK9xTWP14RClvHZ6LQRIHmeJ0Hdzh6bMjPg7X3s5vJPg+RUifiQfZWGZECKwwaA1
nVc2zF66H7V2lPPGGpKhOpCQ4EhY6iZx63ai4eAxSErm/kzwrZnyGoS1PwRWXyEJ
qpspaJCf4H0I4foIJP7E8w==
`protect END_PROTECTED
