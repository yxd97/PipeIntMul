`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qF1fo10GaEzzvkzpy5bhJQ7ZS2g8wGC4JTMCY80xGRXrXNTKCUDkro+40jYw8bDX
3dJnmmt//cmzbMIfcSO4uY7a7k24QwobEKHbTMKt/pkY0F34agoRA3W3YQXt4XTY
djyVDyD9pNJKpNe/4WyOriny+78rofGwXPXil6mm8nfA8nQKWk1bQXiZ9tj2j3Sk
SfppqJZ9TMfJmb4CS2Bm9KJJ78NoqUWUh/nXqmt7M09ZA3j6DW1fAAjneUXdLJV/
f5+nrk9g9HlQDuogzYLmoYO79CMzacUU7voOZGYenyhyHorOPYfLtNFD3U15fCaJ
6rADEVTM9bgjPKrWQHCqNYn6uBGZcGb+KkOVlnSD1Qp+7XxUG6APP/stOhkLXl3i
okg+Qzy2gVZF9JtO+nCxCjZy5wwLlH2dyEzH0DCL7zPYn/xkzKc9FcWyqYrd97XL
OJ3AcattNHC/rMRFb21EvQ==
`protect END_PROTECTED
