`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HZMsMteGlhigyTKpeF8Kju/TTjlk/CFWNJBccLzZ55eQyO5bkgTOAe7VzIfskEtM
VCyaT30ZpuFO64aOxQ8Hvyvk6muLA6nkltgwmq1w2M4+dm7t95Jgy3aeDT6D0sHY
q5QU84wqD0EQPeruQniV0qxJTZMVAdZsmfHXIY+MOlx/ZzeRwhu4H6Z2nlAFKs6Q
Mzbk8AG33rzmaMo6RLwsUc5myxgfoNvjFGbIC/Nw4YhgsRNdx3yfsCjX/W/tNMix
aaToTcc+15aDRYAGsNC9RsHMYxDIK3ru+eLu6zTO3MFNwyIyIARNZg1tp8isysTY
GKb+y3m6fQLR8pIsPbk51gIxF3QKS7oSfbdt1EQsPCLHUTp7nHByfyqtbhGFGw8u
QTm/ltDHE4InD+isavrJ9QvAcAK4kKyZ4wJ89FU/CdnN+6Hkxbq8kS3z9/7tAErt
boehvcHeHulpr+h7d84a3eKvg35pmiimV3oxPEW6CCpoLCfxGgYQfGp40bOanf9P
skoQONRVcubkb77fz7NRyIo8J51ZF6q3xoz73TCHIUdiZy8Q52db3jgydyftMoFC
Z8IczTXuJzNM6XqiVrXg/1I4McqBv8OAJdMLBw+vCcpWqoRpRcydK4RJbRNwbflB
ZOocVZpZEM0LFZoQX24qEPBsmfqTIwIOV8i9X7aukdc0es7ARk6cWPfXjiQdl4eO
8QcxbXiZpmkzXIWESmXgrCKcyF6+0dPkUCcgo6YCTwwsRu986C2uY++osBSOc9+8
NG3oHoLhrS7ZpC730NqrnKyoTx+vxPcx72oh/vWFevmJ/jdKEPKN+wvSJI39pyx/
ArmHwPKRESRU76rbqnQbIJ2P3gdvuEjNerBOtb+jdpbXdgt47hldCQyzrH5HyLuo
LCdnAWlY8a1cT+9J5k2CZ/YerlW6KllsOrZKfI6hOcB7Vph75Jrk2PdgVf/WT8s9
ljk+6ZH6L//YIdHPfqpfCMgjZP9JtuAs4hZmx7ptjrR6tnektul5VSnMD0Jd02IB
`protect END_PROTECTED
