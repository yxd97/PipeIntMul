`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDDDfVkkRJ98KDE3+xFwKTNT/IrE9ghywi09T0H9T/0ScuOUBKC+9IOZ3HLY2kOy
OmEAtDN725gWY4PYM4yc/tcyJ9ZGbcHoDld47qBHWZ3XyB6/btjnMk8ajMSplckJ
59pk/1FoEYTZ8ucxqqE1L+uWT4UCWt8j9DrbRBCf5j5du2xR4kz+6HZvvtz+hJYF
LgZztoUOsQG7q39mDVJnGxyVAEVOCxIlR+UkGaTRuPtzeeCWnPl35X+xV/gNMIts
yX/VtIfDkesADkFlcjKB1ZQRuWvI7fPzQXk+iG9DfwVREckGcTUI3xNLS4bMQSes
mHC8AgK6tAr+pb5HxMmQ0zT720u6RjMGCYTQySfXQ8GVojQvCD+wyE1iwBbO1dJS
ZHtV/U77aI3SYKtsKybny1A75oO9Vo7a1m4t9//S9UPfAZOuk98+B5BSKP9vnehi
/A9RESuxCUnoWtLbPRK5TiHdmfj2Lyj6mtqYkkGGv1o1pktPXSpmhmRT5nDsTRF3
wH4uq+EWMbfGHJ7kn16ly+zoBtpw4yrCC0q4MWxEfwIwJ/BDMy8w0VX9BKPJAa6Z
5dEYS1XqiylUEMTEFmB9F48UmmwZRhcgoV2kud0iMZJn2JfgWtyRRbe9RIvpJUYL
mKiHS7bN9oq7UWPjKfNEaHpAePEw2JuJ9u2hfycZOJ6CW7KGUeEgCR/r5vIgcvue
WIDuv4A7MLvfHlT3n5rcBJayP4w34OstbrPV2NXhYzwDKUBx7EbjEi9ZyW45NJgJ
uVK6dM2BGIf42EV5kBEV1NjvVDSzEc/4kbcmfKgzQ8RR6trB1xY3zb7imN0nL0EU
ZKKcGHchgG1JA26kuVN9OOngmwZg6upiTY6b8At+AMnAwiU8SQTCVEl0oQvfcl3Q
hOoclsdDrB0k9phdBRxpayYUWlCX8A5J2Iu0xUGzEAZnAz/qfVf9wmFbC6RNBRUV
bCG77i8ZuawApA/sonnzZItAzD5WbmTnIr0IgALEnKyq67ldHa3TUbiUz69Hz3ud
yEz1cBOScdaX2+MEfJdxGdxWuFiJy57DwmUD9gCet+yYFwM+33urzXVvAjgS7q0A
P0q4tndgZSKO+5r0DxvXhfnOn25JZ3i5iWwqJdFj/oOTmiUur0qdipt88BYOy36o
/8I2ZcIPyp7GDbTIm5o8sf3+3T0RAPTmeKeBeb1wYlBJ+1+nXvoT68ka7UnPnKXZ
0kacst+eicjCBcWdJgRmgp9nzDgPZQTDbCmlpmGqHztmMzdmAJvwoF+Auxf/Loo6
CvNupDMHbW+wKWdIg9igXYh7AnaElNRZHe/QG0MpbFE2OT2N3+GnAxlpMIXKItDX
LU/rYItlT94iTyD4PyiyKim4LIB0jfXNywQv6r78O95olY63btvrLgFm+vE8rhM/
PNOK3Mir8zJT569JMiop8QN+M38ca+iksSeqZ3X2DAJLdve4hXt04FyfRzFpvrju
eJpyh9aksq+PEN0hdmbdrvOYAvp83n3Wc8AExeRSoCvVNLHZ5lVGZ5yxCHQUeVah
thB6nBAiL12TtgQ7MaPd+sgfMiI3xeZyJCYTcMplJBHv34ugdTWoKWgugIh3oydY
tZ/DrmF1O5QzJ/T6Cmmu6s70JHDH84z89sCwJgneX50MjIzWFyTguS654A9q95Pr
K5Zefk/gA6oyItgqmQ/Qa/a23WOkNaacKQkwtESVFHN6E+7NCD6NWNoSlj3877v/
G1O6SobFxmSOxll/lQQi5JoVECIzpnrDr9rrA2lift7o/kFp7vlpsdws9S/XVmi3
wF2v3A7BA6Ze1VZRnddMKvE7VaDWF/bwvpnCWkAbverVbvs76cUR69QsFDbiQezm
BtGakm9gwiFDW01QH/c06dRP7JG0Zuwri+J0bThPFFyXZs5B3FHruKgi7o2qfnLF
ZPTRa0ICaXDv3tdlPVj5mxnf1iIY0ThpsRBc6jtbbyeYy9TDeUTpzQOpS0cFQqsd
nfMgI1Ffys+/dSv4JeGDi5q1OcDyHz7gmEIprTX4y19r5COk6vOnwHZgu1coM1ED
lXkYfcaNLk0kXwVU6R1DD7jciFOOdKSJrEz/kNNrCeKPb3nUr6RAEnXGt9BsfFrz
`protect END_PROTECTED
