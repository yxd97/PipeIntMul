`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VguwxSClxWJoJ1kQhlFDDtcvXn5aTNY4SGOLQD/LgDupbWQ50tujwDdptoqKF9Ym
H8lvjDqeCbA+HxzceWo0BLgybWujRyQdSF97Kyq9tJOCsluQ5Hx3spjxijPge7H+
E90Hk2tl4F/kY6vIKTD6RLDmoe1DmrtiWN9YtUdXFo0VoxQp9Eyg7ha97U52DWcz
PN0khxikZ36AmDw+aF5/E/lttY0NmneL1Dvi73F+iPXyPhYm5K1RvgXCFbiuDpQG
23fRPNpm4MF5jAzLcWNrRwiSH6jkbwRjLCNvFkq3XEoq7tiustQZUoupxDTmzs9u
xhPfjzLmcTTIjGRB7g4fgQ==
`protect END_PROTECTED
