`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3M39jKJdkyON/t6/aU/YsiXUJcfcIKoqpn8cajqJh38udh1UTc0uFOXEqQ6tvaKW
FHyhO+taV6pVXQBMzCA04DJjqgvXQtM9aA1Xt9XVrLDejIgyZcfB0UlCkNKZ1Htg
FNP6jhX/eQldtX7SleRfTGR0rOjjua/Efka4KK4dliUV0dQUOHC69jn7JKKiIZK0
X6xw3eTZiU8+PNCnvwV1TcPsY+UcpJ10o+V1CFGVw743IucW4kOcJqkUUO+irmFO
PYi1XxbqOnKF3/PAVnXaL7/rPQJeA/vA/YNKQsLGY9AIMwtnkzLuzmRJObXiBaOQ
MY3lz3zT8KINxTMioZ8GYXbJAF3OVZe1jzHMH5V1QakuDaYqJH9k+g40QXnrBkLw
fV2LiYWk2CwxUDHRK9W3Y6s4RQ5FOIgUDJpKpmy+rNgsZxd4OIgzClUAK+QvfLrF
`protect END_PROTECTED
