`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vVPiHrR+GwRUy1VJL5Q0ZdCReixHdhamXrhls7ArSjVi5KG2haMcjCaoR1s1PY35
1IbTGgSCi+YhBygmoe31XuVDQoSZLbq0dV7E6CxWEy0lT14DcYZv7wZj11GK0QjR
yWVMtb1RsnqTGmidrx6qKAhuvq40Ge39y1btMc5j15HfXzTO/0kKpArRVCrxhHQR
5wWtW/p4z3LpIs1lLltFm2RJ7p6YDXaml+hbFMfSuygpHffV5SrGWmAy3Aep7nWK
fY4JezGGoRKgajP6bG8L3zlGxtP3ciVc/yAfYM2cxKL3KHPIrXDSTCj7ov927D9/
Rv0+0GKVhJxZBNUerp2hprn+oHc49H3SLBlvIytTeyTTSW0LtVBAffzvjaDDzIJ9
lEnZdzRj4Ua1+6gyESQcgpko5o/yUMejKIvsvnN+Gb6fyBQ4bjUHNhsgZIXrPz8X
BHTeoZQ+SgtPvbqEnGGyFfRoqgpv+ia6KcMWfciJI4TDtAwUjOWLuI90tE+7ucGq
fjO8mmWPlboKQIfxGbuwU18lH2qvmJMCtnDD9uS3hPWJrhirZXaVzmiSeJpt4JY4
TDV/UMCIg0AquAHJ4iPu6GkDseWrkHYboFnxF6p9vVYPz9d0ud4NAJt13C0GGVKB
J5SBXZaYYx7lbgdpUVZ9PDZF+ttrrQkOcwKkhHkwf0nZs5YIZ7UfqKa+AWsKAm/F
qio5tS17v9bEkNQLTc0yK5BDH/FPBxyIPHoMQHqXJ56AC0o/8YYr4niWdGyE9BcA
9NDe8JRGLWTGDOfQfpbJr2wdHwEwUHPo6NrXZx4gCi2SGBUlSlJdFFM3tjnT7Omb
mbWPA7yTHE9E2FovB4MqNVqOXszPLXs5pzD3tgN/s3lcOyiLxl6jNRyiu886UUV+
dpulNKJQAznpvCtn1otET9BzBJgc24fiZyNwOQVOPTx3gOAoUTyUNb96DrN9ktQ+
t22RVL4nd2S6gSItldNIlJKjLueu/piF7L3vGrVHFvmJcfgdGZ3wqQ2QlN+woOjz
tGtzQyf/0xujwANTtyB7ikO8MH5hGEkywNCMWvzHlkUVnhQllZhUhx2GU+X7L1G1
8MEC0mGh8HbE+JrEc73OP28JYRuRsnPmci1UfgalMQFJcPqiSHfSMKoIro+LIxWj
Rplvg7Eqa0q3B9Rwti761gcnysVQa8C9yHW+N6zWlytXW49u14RRr20WH1x7m/aX
u/Ng/8hpPZwAw5g3puj94vQ+CBKz2yjzYpr7AFr4J5JPdGhms/0M82yJdshNqB9t
deYbrjQq7YWvB4CEy9+HLmGlJk+9y0E2bthOTXwy18Kesyuy0XaX/9UiYEqkiQhQ
1sGTr8nk+y5sfv9rex1xlttZdyz25iNkvFuvFce3VY2LG2T3eArarTjAlSrEHT2P
/ls93HfVm2xHhgfPdE82YFj33v0PvH1qVcq4GDEqeCCK34hhjRseZboh01ZhJsQ2
HQmIAtCQcHTKcLO4xJBTOh/tWN9C7tkrWUbvHV9TmhiDQmL0BPIcNpKx2/Y5rfag
E5SrQMLHbPjKaJKSvE2n7UzcI22E3Wa5xIrcTgp3f6INNJ6hLrFIn7G3nsdlYJNS
GJ85aNSlR+/3mjymZ/mZNsN9QTT19HuMoZ4akhhcynxnK/pLmvA88HI1hxWHbJ5M
XpjXqJfPOi+GwfPklYXvShLtq4qlAL8aYKl6NTSbU6yMsFbzFEmSXiViSwqrNbRe
sXOFce1jgxA8tPwX7bNuiqmmQtgWd4Szaa+oZeaXAeSffIuRSTO930/ALIjw5GAC
r99vTkmWhrNbNynUY0o2gzb+de0UgQp7pHe3xO8YRfo73a04ZI136h+0JLporUFH
EHy9keD6RNrAB2y8txwikrMRXm4Xp6ICE5LDOwOV1sjvX2CfgGGa/VnhaVWeEwjn
BUbGRsuVTWVT1vWNFbtJlJ9pyAektIK55URp2aV57bo4EnPJ+vdSqb3gubty96c3
zj9EFoWdZ+D5DDUqpwWm4E26jFf/ETEeecjG6ebkiIpNmip7923lkww9S3bsHXP/
LP8WlX2tqZ01Q1sPu8+9WoEfcRwQNYgnpIwQKi/Hi4kcOKdI4rtrTnRe0lcEl4zd
UB4TL99u0AGP5Rt130Wnqa7dgwAhntMTk++7pI16J6V4rXEj19nc7nnjmeoxj5rP
S9aSSf3Mgp6mCpbzfbJFXGvekz4sWeT6pry1M53Hdeb3hSy+ID5fAbJSlxcbL0Oz
FJJeS7tnOWlxj30c26cQlWEBBt/uqg67zo8zPf5GgWSAgNM+PStU4pUsYSV+hLb3
qoHUDLcqCfTQNkeRAvkYu762+8UIC4poiTcLo7eoyPKDO1S52axFtFb1v9hP8LyB
xTYvcaQAH5NDxVqIx2jZZfC76kVu2VK926oV1sbSSfN3FESDrBzY/wliCS/B+t3Q
pnJKffsQneAQDQw5N/J0uO733yU/ZyZx82J25OylY8zppwQ251Ry7r30gIGWpI2e
bKPfw/qOFSOFCaHU4p0bZKmXBt9qCHdXHTmdb5Jm2EmbhAuGeeMaedDXC00NWmuS
CdNDPxcnXCQTUR8d08UKt9ymhNQAYgl7V5sHGm/06pfl0+L7tWmroBOyXBqe6u94
YXV9yAghW4LjZ/JlJeQXhNB8HgmLaMAOzVN1/B+Z09w8jkzIhvcOHpw+X0eK+QPn
SODZXsQ3k7vf8SM9yJuDiDk06a5yqvs8KCf36rD8VT41bTU0G9xGmAvvQHaYr58T
0bvGvtZZqX4AwxpYab2VTU9Qdjyu7gxj3vGh7pzjF/caW0IloBy8BGOqOhafYCTi
oOT1sANs8afY70ggRQTSoskQTO0EDWIwbS4CGtGf17VmKD2SWKaXC9JiatUqx+WQ
LXmks5fQ+Sew5cd0/zuOsF1wp7M23VcDSH3DIcbH1gWzlUhwgbL5Elxi4SGy/Xnr
84KB/a9EITxbFnaD/TaWCGJ8x/hrh16w23+mcdkC9GFtmpapLQ/yVgXeB0O4RRhz
NiW9+2u6iWUKOVmIfSsARCynTN60fMwpSK3Xl+W+XBWBZQVcyCxnQlDp5W+ehfYx
QGdIdrBqaH3Q3P6kv5KZH73gJb0wfHJJTR0n/AaQR462PZmYqIQmDjV9//CCEqdK
z0Pf6O2LOlh5i1Chp/2Acs8XeKYY3oEHNlpriwBSgfllDEijDJYW3ocLEddcavs/
gNMZCQBHxe1HNy9hG4vSa5JvZG0WHZHb+SQDUkuHvbJGvSWj1bJZ5cYt+cYLJHL2
bv04JgF8ridY9aS8bt7tt/pEqS5UysXy/RygT1qcaQdwan2hDrEKD2Md692eTxSA
RAJMPohSsL1j6/jGdyHuxg/DGceBYzirWallhlQpGjSTLyO8r5a9tgpk023gD/VV
XxYAoF51jqg8PHQ/4Zz62vceomcimuighb2cyFWvvxzYLt/v58z5YyedDHL3ccWM
gWGvscGf9nzxgZWZ0DHfEaXKmbyOgE8hfNOE1UT9h5tmhMnXJ7Mo2ETIDG6xgy1f
KY6z7iQA6jG21EfApuiD6naf+FuJMdCGbTJb4cVUHZbT6GinQO0KLP3opzZE6/x4
C4nPrXeCEbSJC1WhEWDaLOY7Gg1S6qFz2Oz5l9Jge3NxPgVpNOjvB+4eSjmU0tB/
dj3eAFM0jUn2A4/qaC4zUXaCTI2hrRd49nXMYOLriW25qI81ya3IOxyOMuv/s57e
ODmSeFREZKI2bTcN7jvmSda+3iVnuFiUV5eIx5Ow/reLOPcPr51/T3oZr7g0AELi
X4hH9B81KO4Lf/u7G3tmw+GqEzcvlG6UGc06fPjCeTMFGnKq5FKNrtxedRj4DXPN
9rtrW1fHHdQMEJU5gkMgd8oVnpTLNapDSvJ1KuMqvWDc4WZyz85h8lyqJbh8ENAS
AA1Cc9P+U4Zf3aGSwFVjf1rC+KghuLtmUOjDo3ftYu4Jz1RGbr10js/v8aSr/WDq
juOEMYBeix6HKBBwfeVH13To8C2P1iq6/BP9PLMS2+dBa4XPJsgqXXEuyAx1RuiE
KAjQM+296frgsuCzS25TgWjQV6CpGgzILcONp2Uuzx9IxAoKr9RUzolw9xTVnCwW
PCPnwAp/kF17SJugYPCRIjufFIPmPRAySFM5/0wto2lbz7zRdBklKi9oei4kmffg
1Iv8KJRW9hOgfiQP8CeB5ZlqiTzMJ0nYrbOThP54Y0QBW6XH7eq0cLwPcBUrWkmv
/nSOna7uapBdh16P9wdLE/9gCeqQCRSP9xgFmtAE+OqHVaMfGOoO1T36GZ74N9fZ
+vGMznyvCtoV9AsCLvsOmMvJJXgbaRYn/HuqcR15AM0B/xw+ylc/XapUeQoYHlIF
MTEQSDiE7tplyaqUpKcaVwYov7i/hEAuMSJmaPmrXlnrlO3M0k1RG9HkrWLkviFB
H732cBQd3VyclZ1m0YdMPS3SaIAk+JFtqJQ3t8mYyeqwH42AmKCas08WcEXdUbsV
LOZVCyn9WrDHBHZMpHjFDGUQStzWQpuCA0st6lefcre5HiZk4SYcug3+SBQJNb6q
5XkL/4+p5J0eV40Vv2C7S/FLz6s4njXS2FXi8dxa7xMFE+DMgH434I+OZxTAbR5d
xvRjKWzBhxnsS11jWPO73RsV8Qx6XeWWCikdPf4j5jA8OCQUaoKMqIxNcFUtOjVC
dRb77yv1yG7yIKS1Ll0dIioDZwTefMnfbnSPNI7FXkJuiK319cnBpYNbJ2Kf1q2o
zgkEK+Ocolm5BiwQ3EYURkfS+DPWtz+m+OjESom/iJiDmzvnwhQSrM2IYsnywJfK
JuWvsUjLAytjAWcJekLFGMhAuNOhaCvHxgkOzWvvfGljeQUhi+FhRC1/JlTAbI0s
oRdMN+B7B/YiwYn+ZOjWGo+Witj8BebRLtQ4gb2UuKl8GOOgd9yTPDCRS+09ca1A
pcPwuD8ajyXMrx0+AXsKKcxi65cfNB4kp1PaOsyP1ftHeugYfW90t0BIp90F2+KT
34nOVOFdkm3h2at3AoW8fpKmarHyouhS6vd2dSkz7SsuxCuNi7azOjPekKYr9xGt
cI24jnTlcmrP3z5IoowGhdTTGoIuYv+zk6ieJmpk+4TwuR0aM7kwYlYQ6oEj5Afh
BvGC56Ti3XC50FxndPu4Ob3xJD06AX36bjvLuYJmympM7yMpxRb75G3hV2eN3JvE
OnyXFhCUQeNuaSlJizi/KLmiV1NmY3BLWXaDHhmDTxt2C66tsqWjo4oTgK22LF4Y
l06+p0fh73YYEOZCJrMHLJmcXbuCDDSF64XjxEHcRQnxj3VUu1FAgBwOEJ1SlmmU
xoCkOt/L8a6NkaZKO+rbZ4mRvw2g/URXmXNmtOdjgH8/aDnRTTDTTZHwvvK0UMMk
lkrfjDMf9I2hXSCFOoBMqbkAkf0ksUftrPog/L+wP4vyW03dW5PtcLk7jUfueC7i
uu9GuxWanwrtIgRmGnfActHsn1MTFrnQneKu3d67YX5NE13zaDjy5LbIqvhTQ9bx
vf26as9Q9Z/ObXuw+yVz/ico/iJ3M+OyVZ2H7oh5xOJcjIOG8GYoFvO8+IF2Kws0
h6kVI7M5mHDYmTdVqiRQS81jV6YbAtquU3PSI6KuNoHRhNgCXpMjFxLgg63SZxlL
AdKqqAmStP7oiEqO98tT0BIBvCLC6cRXR3R4Cf8O64SGjff3o/h159MZh0YfTcfD
Lyt+aOv5fq5eH1eaLRiPMZ9fsykQcbn8HzwClVG7hwNnQMvlgRy9n4kUVBgZpF21
p5Sz+nrPkqujDUopBoEANZEZmsQCaK5hqcbYtORYXycpNUn7aJXaurRC3T5cFc+T
Pz5chShLetK1y6ogeLez4EXbfEiDk8XaSxSXPOBrPvqEXlhhRPXTpVJ0nD387eYj
iaVyUThINzatBsXUFDGzaIDR3Xi0lodWTI+5sUePI4qlJap+IMZ9sPxm5swZ33Xh
w25Cyqm33O01y1f3IieRKpxtlz74HLaqGjps3xVp4rNacnWH4UrkQJSwpZXMxua5
idfPzUaELzICzctxpPYOf/MpYD1nBNA3QdrgUz+GpgV3uSEqtTpk8VS/McNjjJZW
aiqJGendgFxAOpCJzkZdQVI9bPmZkuIOjyhxZPu7U3ywUYYYdzgromB63PljNGqJ
eKO4cX3YXoO7y0NzvoeKl6or7vhpgyFWhfM36Wfnvx5Gn/cCkWXMQtLm04miRXSK
+cNafb9xddIYwmQMXhzpSVwhkq2ScM8/ABZBosPcyiW48QRmuritoQNlhxXkV/bs
aRF8028WhhsR1WvdC2X9NXUvCuYM5B7epm1FRsomKOT8Kj6GMBKRRIVkfloMreM+
C+q9EPXwP1XFenxlpv0e0jBpVgCeCNsRFEW7ChKueXIivtRNAuCvJumei8hR7Qva
cPouSOcIMD3MXTffE9Y98rX5tTRlfuyLQOzUU/c9TOuqDOHqwgewqDzKc1fzrcyX
y48PavdG3s/YLNBz6mbpfJrBvPYx51uNEmlmDoZ1ET5bcnJo4eu+0DAC6P/yQm6N
rP7V7Hr7JJbjEuG1IfbnfinSfegLIT0KvKlEMak6MVy+2NJeuIOgopbOiqn5qwMk
gncBt0iE+8EjgMEo9ytLTZbA2dL4zJ8aH0TcNZlu7DoscFSshIQMD507PjE//GKk
6xOtYJ2M3FOMxiBiuffLnJy0o4rIePUePK4gsvSQ/3/X+aC2K6nqSJta0ECOACfY
9+fFVU+P2JSh3dpHCp1S1b1CDhp4fCGOQfaJty71loxLgvxuaptoADHgQwhnjCBS
gDsQFbjO1f/7Afh8b1iwX+xUXrBjp0TZEsEtmK0cqKqoBcv1AP+HfrQ9sv8e0OE2
6xDQdF9fFWs8IzMaDZqHYam2v/q/AxrOXoqxzXviyT5hjMf0is9zWBa/NJjlhsK9
Bxnnv//9/v9F0J5LnYU2Ikj/3hTdxBmG1zj/SaqhHoi0y/i4d+02oAoHKJASODWM
aVy8JZZIi1yabfhF4PLXtOa4zuc+mjaC/Eh8D0Btx5o65+oDjZWj7tq0/k886I1L
sr4epswu0PGiBErYmGR29NWVoPTvWYtWcBaTrp8v9DsjVZZ0uFdVaUyCGIOsDhcx
4+UzzwVtoE04TvOoogP0DguNtKxGuBhFuyhK2bQOtA/+bibUOAZ/58xpDU8o87Bj
Imn2uWP3BAD2Mg7haR1XuY9dt6/DuwHLoCLV1vhEsT42+6sBoOEm/TtJOEbZNnBH
i+oYO9a3myp/Qr6w6s61aeszoK9tAIPkyQy6YasyWFQVRD4pi4ypSRF+H/5+5oM7
/QJXdJNJt5BfywdFleIT7oFTTZCISFHDDpcZUQJZw7PdoX9LC6KFsAwL/NnN7+tl
8s46Gtb+VIhKqv3+sS0LIBw5j64bI8OFApu3lEji86Ksgd6HoQJ7akeEtUvHDxv6
QvL49JqbeORzEDF5taSxWPSM4uA+AEMbwGrQuNk1QOHbV5Ke89KFSFbcWmxxggax
jiWdzQecaFDisyY/VWKfTVaCzPkqbrNRhbF9bzZqXS8IbTJirHiKltx7L1eNDi7Z
L80+x7FrNrKKVUl1ljfDI5uDYWkA/P2dXNxeUuFlLOcvRW0MTidoWP01dv8ESCqC
HasQHsxDBm3g3kCiCQh0WLKGktIfsx6D4gAvc2rKeU0atSKeRvBC6m0UjWAr72a4
WisfxioKmr9ToHMp0nLPX1zx6RT9L6l6Xc5Rlf4iJzebGrEHOKRhzuRCoYdXAxUZ
fJ+/VaQJaZUDj9k5usD/4lSwLwAE1YC6S3Zk0r+Cql/wQ2rivVjbxD0PD0P95kXI
RiQvU6oMZMV11mWq/UnnygRv4Vu1jRQn6NlIT5Q51BgrSy3doJdDM2WX2PghpNQV
/ua08NCtgSFLfVf+bxSgs6XXzu5hh5wvYdyFRhRMGeamuh/iVIriRnoCkXJF97sh
p3Tqthd3lews4ZXrT5xxveLF/bFqJH4GPK1dS4uGcwERs8pD/kXFCEDPtq3c0xBe
aTQYnBt2NkLI1jf+9ozRllueeSxeEQGuCFQQDW7t+6UsIQJWJTEybhuPhwHWnSbq
Qq/pNIYfB/otbP37GCC9rNwOof4VwiLspGUj3f6WZMQYZNQzAy4CiAd588sHDBlQ
DQ1dAnYXFVrXuW6WGpfBmh6mdWR7Bi/sjKmyxKm4vDssX2wiTu5oDOosw7rhQPS2
w5HInvWC9yCJvhZNgsvC2gZ/bsbEoByVv6+fp0NXPlNX36s921rw3uLICiOiPEew
X1EaVtTMVEdKmsmAd/TbO56kJm/raQHUAzMwV7BQcJMDZFMGFyJhBoAdGCme+Cxh
tFa6cUQ1zLQ6y4etWNzNYu+01zaIm6kBZciUpht3ptjxePO9l+37P2hEL80EUSGT
mnyV9WWKB+8FS8fTmcdaBDiFLv2MEufheB2N+yCkeOtIXuzz/R6/t++d7j6hiknL
5i+sdzTRFyOSQ607MEzwOk61PYbabXLCrnBW2di4PbOc4tARHP8RoVbz20Zb6mXZ
3nd/g8W3vISln3dG50/BudEqzr1bRwpm2wFHo9jZGXa511MJENawDvYYYZCJvZoy
w+LzbX0XDfQLWW0gznb8HH3y8m0yGLCKkPVj4t8qvaw+mLvXci/4ZZGJvUSb8cNk
FmEMZywmNGoutN8xL8/x/4+h4ZYscm3GoDk0Nmaw37ZN22twtPZLMr4sQA313Gc/
IBo0gZRvB/tHI2Tg/WcQXpyGNiBJVbJjx88PPVz2NcerUcsWvrEH+2hw+V8ndCvm
DrT1kGAUq36Sc0qLjmKeq25x5UjHpzFRwxwYBdlfz8N5QkcXCOUqglRfD8BXrEPy
3+KJXfKzbOC4Wza3H9kI+ujDYJJKq0TDqKQ/wXvfCFlUapAgKuCKjvaN4eXBi6WU
I/fRSjkH4dKOLSy/39Hie1M+E1cMXb/cUModpkzYt19I3TaRLz96QFzeHY0ASSt/
xXR00ex5m+a/0L/fWC8mRNkNZtoAESngO3dlyHD2tW6bfCplvS3u7ba6rBpZ4nIY
5WuiY2DbCAEHph0WCH9m84jMD2eaVqPg1fGO5H9VFfjXtaxArCUnWk6QyKF0xfhK
xpL1Wme1/qg622RFHRK1tkxwGK+yxuJcgMorW7WkaJG+UocGI9m95IXU3zTThA42
Qr9xapaJqm9Pb6R8F3xYK6/ZopRvDkIpjLUCRwNMRu7mxrlmoGRpUwKf6f1fH9nv
aCRUSMBiCq4zouDCMfC/Dcct1oSpzMqHm7luqDdkqzXX3NxDGThkFDxkhQ6g2dgA
6vlAoocCMiqlWWbDxn/WTukJpyehY2VnNDXNJy9+Xx0kJDlQSe9uwXR/fVU4LDdX
Vo/OTFLHIH79PifGzYY5cysK3Ia669KCgXqmtte0OpE9ubtknUs5mpifWWJIl2X+
SLWm5vZmBxME+2ZTdV2o9uSPRoT0nzd78INkWWiQ6DdEJPcIT20ci5NpUij18Upi
c4Ao9omIuCw7UVOfgbNR49VOmN3G8ZIjAQB7WqJ4vsbpr/D6hZ/s4Cdtc/89jJOZ
oBlwiVV5QdYPHvZurSml2oIAQPH3tDYKYBSscvuSUOjjWWUFsfv6MJWpsUIsokXI
cQo6o4+eAikFdBhtezZFTr/UTAlS9zn2IXwnQteEOZ94V4uYZN9CLwJzGG7IxAfH
KB0Vy1r47HbKBS/NqLIb3M5uwTZOYxp46Ntg0YBD4/5xoGIhqUNG23ggqk7Lb6l5
cnPUMHhx/p8qXmYuQFelpJfY5UmhqA2sN6QIx85EHxU0H9lOSiw/IE5crarnsM2n
E/u9cO95APutG5S0kMj7pWuc2VUoCGqNrYYeqTyJpGwbIj/cZ3+HXn8n5Ufv+Jyt
qXRvQErMu9OMj/LWlEN1dY6dgNjj2rZ+/WUVFO1fa/vXdiB7JlOSVIJnPlJ0Kr9E
Q932dWjD/cba5To6CaE8OdHYWWWlCW1A23E+UQ8HVRenJwGC+kr0XWUXIOThgtZD
I3DTytBcwsrXJZTQ+qgxWM/Leb2b9DfZbztBO9KJBqYPCyx2mrwRIxGXWoCrr7tR
bmtq6bDkaTEo92xQasiupsFWPz00AFaARDnoANxe4m3/fdFyJCszg2SuIASX1orT
aoPbENtP5jVagNO73yiF/bFp+k78FQAi7flFLVPmu4mdqIvLw+x2d8caGxbaT54F
uE+WtPW3xKyTCg+lBqR5zcVFVqmbvnABeRuL7MgbTviCBIl5isXrqEAUih6Zfp0C
LsnC2+NWMVcDtK0ER+BPRrE172DlaYurzK5DB6QdHn9uaSW7udnHEQHn/YC2U9us
Jr25MWwd9XOHTvpQV95tT5xlY+R7DpGD8UwZPGnqjr48qGBMQhFHBe6clCErGgC5
c4upJf73Gmmq7DixfwMWsyCdYTm3LXKGd1axLWRbXxd/hdDcvVKR4IEEFoM4oiGz
INEmRok07+MqRzBCnF9aTvglk/9d2PnbU5Go8x9qPlB44oNpmayn92b6/xWUkBac
BLsVjvt3u8QJrnf/uoFGeVH3POu6aaqKpfuqCUJXYE/khgdbqdvwULLOqXp3Vd7J
c6u9eRK0vdwcDx6+Yvz9hUHY9tJwqM4hY7cVNXxQWayAOu9Gh7baevw72wRFs8uB
LdrssTK7Y6ANymdq0pWiMnZSV8UeehWr+9fpv4T9QcwjD7ODaoyYO8DRuV0LUt3M
dnUM2Su6qtFrVrOsMga84SRMw+8r2+dH9pZb/vg9/XTD2cQyS1rUyXa/qY/A9DEm
0hagLIvR15Ns6AY7VqWcsZkf+lQdI2oY5X05e0knHkVkcmSat2ezF+QaLLrps7of
DH0VSivNveWiSHe9HJqydLfYHq0RNFT7L1c3NKmZI/cmSTG3aSiWAuMe426exBWi
wQhP2d/ijQ64K7SA2N3yV+vcTr+R++Hgbl3dYeFaHQEIE5h8UwaLk3aq+tpDUXJd
7LPVMGCJYJ1GYqjD1GXeK8YXW7yDK91wgXjnHR3SY795q+KSF7NYoYW+NDzKlt7C
g7eFxZRLx+JAanQK/P9uz9UMVSqc5YK+QqhckDHM7H01bXnFjFM9gM4q2Ruq/40Y
DPjFzfE68foXjQfmgKA6kYftTn+JUSglrIFqONhFllttMn4cHMPvTVuEno9iObFD
iiI5r5XqXm7fEH0dNEfjSB2Lx6AxcJgGFg7tCwqqeyoSOTZaGjW4V93wJ95dPcMB
rKMYpRNjMu8zl3Qtl02YYuZyXHVTt9e8L5btVH7KifbCFUiSU7LCgrKK8PscywxU
pVn2/eZQSGwW0jvXQgiIGSoiX/i0mauKjcL8ruPtbkMPseEfj7XNlaNWW3l71LUd
DE0NuT0+KqLgyZNgviFKgA+NJYFjAhnhETpw8fuxq2BVBSqtVkLNJvM9QANdmTkM
kwUnzaSisER0L7cgaEyy7DUG+VeWjbT5cdV4DPYAloDEM7w5EZasenWrB8QNW7kS
PeHawIUDADFD4rhRgfgGXvS+QAhAxvrLo2NAf3DgNssc/b59WGWGG6jWsuEoMkYt
/gJmZaHM/gV/N3ugVWKDRXJUn3eih/1nLlA8XUq75nQFuM1b2/zcL3Dz8/aVIU46
jWPR0aCoUR5R6gj+pJhCfWwOEJjQXnn7uT31vffwFbq4ykoGJgJxJTbaND2q5BNj
kuxy9s0FXuRi1c2GSVAhxFZgnUPPSVLYY7Y9Qdp8Gy0yW7WRO82evvXC/g/ZO9UB
Blp7TaNQNHvbIXumfU8h5V76sHbG45kR6OjPw8zJ7rL0qHr6dGuIMVsmm7c6IMs+
A902h0ILp3QvT99gzn16m2LMIVHCSAqNZaQeV6+ta35vx2W6S4hfLydM3MfdtTlA
JpjluuDX1PzFQdnymTyHBAPVC5uw2IdVgXkJvEzpMKGl2/y7s42u+WeQhSckDy5l
FlY1TSBN4Jl5UdbJfkh0nVptbO8qnwTO4HiIwspZavub0lvv+1zjTG7Q03yodrKu
OEVIWnKb3qjMDzw/iMihWGMTpx5hQ54ZdDlaR1IYSb7fM2ZAkfib0COxB8BZTj2B
vUcTmVfWhczg6qpH3LDAaum43P5l2xcYL3+lmt+W/mEcPSjo68IQRAXt2dKXjpFp
QRokE/FJBEb5A+rTG7bdcmu+cdCN9+31+LzcBIlZYCO5rbZJ6oJ94irbVasUgyiN
NCTTDjVE48dFoXTW1WOoF5TPxQNidsAT+R3tDApuR4UpRlhPvMOKu6ddZnELvGsr
I+IL9olEQRiXWFrIv6j4UGUxxwpRTxmeCw0SbHF5IyVxkbd7f068wJqvbpeT58sY
zE/Mb1gNNktYdHgTvFVw1X1gux5m0rvGCh2KzemCJaUXO3xN6vlUoVy9h9r4Otoa
QurdDxm3SHA0Ic8oHAqgniHkqEvK/o64GKWQh/urBTN+B+U18LO9ff8Ux414IWsG
qV5zRcROMiWA35wviB2fObWmYhisgIiHxkTTHTqbyteMK2KNEPFOp3qSAxGSBJwK
cBJA4TQGOm6rrei60UpL8FbKAF8COFsBR0sPWdGfAUxTBN1FpyrZkOj0qz8O5+Mt
2unMQRaVRT9jfDzd6Bo4HIb6e09eacS0dmoQM0NpgWA/lgJ67p5cKlAamLfozPif
ozkkJ7rzVQfIsMlvf30jBiW/+rjZzRJK7vyq9Ec/7hUty5+ulrAxpSNxj+jZzcLE
HgHspdLOxWHIeMzzb+/E9zIecIyLNDubQ7RurGn/v5ZSVcu8NPO5Snulv+yAheSN
CfRyFOjfRRIZ4HSnhq7M/k0LgUzydZ5h1Y/OIq28amVGtzoohks0jowFb8jQRUKb
MgE6K5GLZ8cTzNMQwULzX1Mafo2HUrVzvhSvld/LB4cFFgWS1mHou6T+569qcQ4Q
Cq3aHggR1ZS6NJO0wmMs1pOxWw3/BkrvD0rR5GlJdeuO2ZLTnzI3MGflz9fLS/l2
bmdotMLVVf1M73BfTl/+wkwEraN6uqsdQl69pZ8MoKLVeUm5NvlD+om4oTWJMUn+
hsJ6Ish/uBnzKGzXhLFNIDxRD1p3c5mDxiVE9FEyWna6q0UIkuIjk+/zhfNc819f
UU5VdVc0QKbYkdCOzkNcp0Xy0bJNnPv4xYWyj8M2Yl1LWTfx7acwktn5vHGUkzQp
LP2q3/jBwpmVs/d5tDwyt0TawGRRlcwSTukL9T3X9pG4r4WuQH4D5BZEjLRhrsFm
Ye+SvH1Pfxd1cGKZsCtV7yv6IgnRYXzGlEifznzDiyyRPy8K1REICygT4IlwjV8y
D0HrKcKXQsL2SpyvmfwB0JFM3xymmef6kDt7+2V+8ZjITgNoEpfvGA9oWdNnrh7R
VHAYlvbNPI+bmiYuAjNKqdCLBliK9Vx6eXohK7pHDqgWUzPnoexJ06av/BPvKi0Y
sAxnykJT4ynxlQQA0tD1E+8x87rEsEpsrMxDtCZ7lgKP2iZo0ennx1TGIqUI4Eey
AoHFqL6qxxpxOYzHEjB/5MQAvzj886ntYgvd/5F3pzrJO97wE4nZY9qrArh0zM45
mqN45n1O+/uv2D2oCtbQpyMmhxPu51fOGPx7kzJhfsAGqoUN+jIAWsMh2dHYM8XU
jvEU/I1OobzM6JWV89srUpWzro/rSXGScDSnp4SbBq2kv1lZQEmTI0aI65vjJs3O
XpjdhNYLzM4FUmOnLB9cTQo5LPyyJueLzRZVJNQ5SZFIt0JNZK+b3/EM/9BFo5jB
+6Z5oEGMrtb8U9Zfu157/i0yRIJ+y6LyeUMbDwtZ3VbL6Xi5JYaIBgm3aBjt27jH
OITwcPyq/Srts/GOyW3er7XfN25SdXjvSJGAfxKmumuSa2F259Oq5K8tFGaJMswE
gEmb3yiirBNk1gKcx1qe3Hhu9CtJq2vvYoOXZzSw7Fv6Qb31OaySLIDg6/mtgp49
NRB6ObQxxbraFVtHk4t3aJ0vgTaaDQr1hVwL1MpC8oo0yhCOVMMbBNEnCQBwBoVu
koe4oC3fALVefnIRk4iwmBDyHxQgeriZ/pp4Id1x+rFgZTyI4mFf8gv45Ht7wAui
Ye9Rtd0z7cyePCEW+5BlkyQwNeyZoX9wqyTf6EafOVXY5bYvLVjPmAvW6A0yDkE5
v+8T+phzCS34t1FAO2+d43/55FXFR+TfbGM+0lgP8bhnwSAVDfTqzv8+sDMW6MCb
58lI4eBViefZCdzWRo9eZWoU3d0uYDRi5/ZUhYrbiLasW8fkKpd7iHnKdtog9Cs8
ufQ/Os4nmlJkVKay7lcPllCqnbL33GrC8d4qRnItYspIhwh1HkDJKg6kKq+1hQxy
XkkL1H8jZOQb+RQWaVhPaByKbIdZeP+QA/OUfBdlzxM0Zki9t89L1S9+GVrHeONR
OkmHeSzR+fHFXljgPXI1V6yaD5NBbE5f+Y0DFibCPsaFfJaxFtwAL5dOFlNFN8A8
zvG+BGhuKICSmZ9f2NfZVlx7r6zC4sl37rHaQVMU1O+u12ZbpJJ/jA1WA6aexq5l
iBkcknfGK5cTlneL0Gl+TzYEFA805xRGbke0X1XN4GspbknhGtUvZ5p1H49eBEoU
OA35HyNkE1jkKSuFdh/Et3M3Ki/IPzvUCHkAxacDmiKMQ0MMOBjQEH2v3UrQ2pue
lxmAwVYsXibUh76nazNFHuF4JDEMYfxqvZaJfsk/HIEWUzy2MkrryhryVFQhHaoT
DU+nB4SQWt7yEWQ9sFGnI1Fad7SKxnh8b6Az2MZ/r4xFhwoklBm+On55tuy8l3mV
MrWV7aUqBEOYp5WHx4w7lpAT/JvHo6Ce3lEV3sUqvoPKRV9Zs8y8Kgqad3z9ImQQ
VXaJDqE+4dGjgEAQPPWohNU1WGVIr/hPgFJR8mJrjlZfxNrF2XgPHFiyOmNcAeQR
ShfLvM3uHsONWCZ7F4hDI92PB+u8feckjdH0oqEAEugYWXDAEC1JaXM5T9CaDVFe
/8kZiSW/9FLWG73FiVJ0v0nIzTpIno0UQDB0FU6gG5WFzdCYiSeXyGVCnCGMIUaA
cN6Cgbb7Ypbf3sZpEf0NX2ai/JTzc4WEpRlzxZllT3TlkqH6788t0b+04rfdQhb4
x4jiyqJ5Bt5kBCSY1t6/9axLhKD9+DknJ2oXr6AO89zxZyIJ5pxflOstJ5eKWjqn
NndPhYoEcCyzT+MoSJUm8H52rkt18dFaEhlVCVwJ7imCV70jFSTKF0g4LxorcD6r
2Ypi/3forSBbZWSFX3drn0lkdW1w7NYOIbyFTi/HSqesjWhIqNP0eEDNGDM3s25o
Rlgy+xIzZtOILykMnQT3zbvJ9wIOGgwrag1e+RbtCcYlEByzSS0qJhu5wl8Rk9c5
jff24z8PkdATCXpzPjIpvktXbYWn/b8wWUzJY676vBfR1Y+CAW4gIcxhLaSp5Je7
nOcMuvVgOHlMZ3sO7/CUfoR94MIofE4yIh4hdB5wTfSeTSK9tmyjVmm/8Qwt9UqX
F6U++5w99KMQj5+c5XSa+7aBSmMMJS8c92q0qql8gkYNHblOVIBUr+U8FSlhvPEk
3PVC1L9xJsDCdNS96NKolSxw+x6vJK7dPbpCFmCgAwpx7mE+pLk20uYtIFT0u2+H
EcubLlIL9FhC/gh2WBpfsS95Br9eR1L5feTaGcyc6tx61HN1xYsyR/iUDTYzv2Vz
ciL0FDy5KxWzwuVFPiG+H1rfttkPWOCaS3i1PxMbyQN/bd+tArFQ+g3FegYmSEYu
ljGs+xxKSK3/MlUg+glxPut1dmCbW2JM4hdJJin5wFLkBSgEPwh0oKdWO1KFOO+X
NfOrKcKUNdSwQTTuXKRh9uqbHMT6nbl61pdv4lypc5X0SgnXQXV/W5n5Xh6r8Kh1
Npm+tdzZcZPHnEK7+NURdx8SerHZ9Ii1788IWR1O1fxyBZtxUhed7JlQcuFpGrA2
RILQ9rYM2wrtkPbDOSqTGAQ1hr1V0wYAk01Siyvm/dS0eiwM1byqUzziJRCwyg/V
Snl1CLKZiBLWwdfHYVT3uwy7UsHBpNJp1RR/Psd+FCHVW5ciMLmPjeMpNiQnMVzP
NHQhCd7MJu3U8WMHZe5UkLLoz9K98294M0mfB6NCPI52uoCKueIf5rYE+R/TYkGk
Uf/yqAY9JGK9irirNCDNdqTjbHg882MgEh+Do95lnMMzbFoMfcZCf0PGs67IUPKh
n1IRLxwXCQ09pH4w5b9uUKVjs96FS3NYdSXPoboh4QqfS7EbMOQGcvk8gQoHktcI
YYEVNPjEJVJMuKOACM7sNbTPaaqNv0xsU7WnzUS4cTjyQXUQUpE+IsmPy6LafNX2
em9Opy/ctMZ3g5MH5wcAH+h3erlIVfcvK/Ji+p89nBDU0KRFYth0g+hOrvvT72/q
qBFvrzREokCJqDtbTPLXU87OAEaKpN5mYMP/gEZhYH6Inf5zQZNntFPBBhZXgCrl
9s/xXxQt9WPeBTp9HVEhSD5bADl9lJNo2egIV+hSr66vNGPUFo6oRT5BzDydmMcH
ae4YNWXFsbSnBOytE/c3XNUXcLQXM/ORMQ7Ri5t9jk3zWQdcEch8wts5g3Rh1yPH
GGQGZSZ7O/WsqRVwCsLMHhj3Wn0xW7QTAKFWtJQSSO3YEXfQ6FiSKhYFZ3mZml2O
aCj1vM1+fMuYAQQt9X+8utJ/ep4XJzCLlPh07UV8egjybt8TEeJueqs+fGXee5mV
5Y1kiRhYAJ4FBtK1RJgr8LmYeZqL+LBnJfF1LYy7RANgnOk8ZNJVtRBXV97GWUEK
18FSzKvJL4yI1nExXxStOYwSfRwPEgbUMR2p0SIRSGMQeSsk/3ja5gzmSu3JoO7i
9arnCvoKCUhF5Ok4csiTpM93jAuCE/KoHOSx3fB0pVEXV+TKIjXjRCLa+1jmwUiw
`protect END_PROTECTED
