`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dcW9VT8LDDk7FEBtUHFdjm6ytK4aG/Hf616Eo91nS5YUZ6mAe53TUNzfbWrkeX2a
IeKWItTEvKQ5UU3eJ1Fss8V3+LSvLIvd9OZaFwJ3N3Q9pJC/dG9SBUUxFxtsZUnS
YYa0hdZhg4R7WmIgn1C39Pk4IVtIftikZs2MgR5ia9z+oQz8hGdImGw9pNvLSmGA
vluISkUq6AmcNn/pNIStPnBzUYVsO/t+57GKumZcLqQkbEHvAf5m2/n7DvaLN3b8
TxIsI/SFB8eeCv3t2Mj4el6AfT1N0GqXfuLOIJJmNHbWJxsdm3lYAvW2008aaEU8
jBBR01yDb3Oki183L9xJQPazAtGGHlBiKHikCzaybe+xIfvFJJdXMPPPrpSg3NH1
5JODdLAkPydZWYEfq7zTJwI4gyJu1ubeEFA5jo8Fd5Xk6+JoU88jd8vl/D0yjUAv
EyyWHWVHYMsXXxEyilMAYv2eQVeRJeQNA8bw7LcDulLQYIePB+qUtJDTobsSHahk
Z5OSarCNFJXvx2AE7m37UG/A+Em1zFXZ/F9kwOFJYn3PbH5PxKoF3qRrtefqnmnK
fNeFQQKeZk5HITkhVzJa2J8mQU9/ukFEIzdlR8yI24nQHTcpxORT9jXL0LGDLWBc
9KAJJPtcd6zDCQuQcsfRhjGNQuQ7kBD+WCqy9N48k6Jg5gZG1x/DSBaqmvecQKAL
jONA4jX4f1JbWU66WSBrCKpXMmzzRKF4vIwqQAU82GMSydk2AGKW7JuKwWmQhByC
N6sxM/3Dj9Z4B+U+CzsuS6dcXTTVMAAgkvvCJJmdathiJYdDtu+cKxZlWZvVUy5y
H7b59dVxezqxKu+pQGwOJHXc9xb9lfXGPfbbLMpD4XxVdNy0VgAV1lsp8y0jDqM3
C2MSwEyxRafCwVlaE2xx8NaKOud1xfbHn95QPN7Xg1SGC4VjP5UqTP7BiycPWKZV
Ar9LxXwoO5UGhdE/ya53k2acdTO44SGVo2xRziInIOpuW38jj8YMM8m1wSObpxH+
`protect END_PROTECTED
