`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lXWSx9NY/QVe6GgwZ3HiBaUpfX5wFdezoqYVz00spkgvcZO2psrFi5RWKmYSwfJd
fFkATXYemY8rOEFWfosMOcRATsKFqnvkmaGLhlraTHXVyRX1FQFqlCzVYTqbdJd1
IV5BLQacsH7/nUGdoM8P9pJ6aafWje7km0EJc+CCqWG0YIYLmE52xKzfHEQqyPKt
jNed75KJtPOCPQSfSDCTdGM+LaRsFXoIf8xTh7bv8ymewMLTNl+ONjKY6Fy27cWq
Fh+AyNSu/DBJpRUlCc8xFMhIs4Z9l6Zkvwavez9Bio9zgf5nbX+PMDDnn9xM5prF
AEbvgcBWVE0dgJhG+N4z0zwB3xiUWKAvqnI2SEHIbeELWhqg/n57/hLwZeoJkDuX
b5boZv142fYgrfMd+HWnrt3wS4EusVa6VjobvsuraFTt7nbZ2Xo346PswsxpgIN5
FFDApaz7Rciqk4v4hPEha+QzbKdbAnWDti8tfSSo3sviiCZ8Q902mAKe43+OFyQz
`protect END_PROTECTED
