`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZzajOpb3raUlS3WMBxHkhTmy8OQpHjWyb/CI6mKxumxeGykhZR1H5pQ5xh4a5EC
lsCLSThRqjdiJrOe/PCooBxPrFq2Z1jO1v4wPWtz6DqfqmhWKcISuc/X9GQPsSpv
NMqIiVDBxjg8bDBYd6fmVGxIjrx1WAiymR1smldfBQ2uboXCqOOxqpZsZTnLTzmV
pltE9JalQFB70UeDUjOWOj3uLOzOO1Vuk5J509CTsObpuFuPBNSObA8dRItyAgOy
yyaXLeHnarb3o1M83hAmSNhPRLAR85RKbK7l/I/afZPRuD4t1aQ1T2AA5C5AV8zN
IdA0dwdbgdO2n5gniHnxrA==
`protect END_PROTECTED
