`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vffWmGrkf+YOabbfVxOAtXTOpTU4ziDRG3qeF3ANnFfY1pIPT7jaPepnhlnRg3Ag
CqoD/r8yoRjqDGxsGeX0jHZJ1ZwXAxwXnBl5HvKQmP2+UMH+AyHFmDZXTOVVBiaS
zZwPw7f2ktdLpcHDzw8zZG79SskkSO2q7wqA6o+BVn2A/NQqqGRS/D2ABBFrGIE7
VtZAWC+NKXQbKnTmHgImv+MAHxIHBQBoXrENi+70uOGtcKahjJwuTcbv7X5JYOP2
D7M8YNnBOJIPIuVzI/Ubj5VxIL8egoB0Z7V2eEfgGkk=
`protect END_PROTECTED
