`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rtn6BskW/NlTjHuZHg75lsHSZnXlBrH4LUMCvBs+KHAWUPgo32i0VulPb6O0lddz
XsG9LAdpQCNFRg7eAg3+U1kMdCWkJWSzOZPQq6vsxQFFauN5rkdx9SOEXtFTwlDM
ezadFScMsf0TrzrpTNipVLpZwQy+PQiXA6IxpUIP5sAiuUPWs+ppsBJ+GENZIS+l
uNksIT7pGnC0Ns/+UuG1FwefoQdzOiQSKs84Kuf7Z76L1UggbNTAd6yMlT4erIvy
Ql6E+OIM7hKeSVQXGVmi+TwO0yPtoQky/vTzMWnoAyi2F35PxzqyFYYwUu/FjcPY
Wa4qf4EPgNmmUUrGIFkDwGAHIrDU9in/iRcgTDwnDQgu7XPWWUpC/FCVGWlsvcTI
dSkSM2xughj50tuWp4MK5JoHZgOh7wLttNILzalG2Qrtgx5nNPVNKXqYtAm7Vxws
IeIDYmKKStVMPB2lrxi04ge2DipvTSTsL30wWQOY/wKmUNo0dOkAoJyYhyOWZUCN
8nZF2xOCdIVvsKS/qm1kLPwbaJJ2/K93082NDuPeAdcH3H1ZXae9xso4BeiOcMLJ
afeyr1Pn9pSCbLEpgER+XjnCN6SNvwgglYT7b34mm7psDZrNbR7lCPb3PS4J4/GU
WSTRc89dG1EB5xRGf0aqu+TzmxTFz9BvzEuMbNH+9cYY4SBm+4gvj5fGM8qaIoUe
yGF7fNObOegEYigQCMSTNyRYpIjB6GFaU74CYx60AIOzzTaphrUY0H5ukiUckljd
hYRKJ7Xp2eXsH8PKpLl54D0IzusGdLXqWOwrXymw1Hm0LV8DU45H4U6HmScpa61a
TxqWuhpCjE3pRoE0/RXuq9eo9C8lthkkwkw7Nw+ZPG0FIt1heEwsNnxbWyqP9Yps
HH5/VambhnScdjHcsaJo3mgpcUf63d6fW4TN/eRrjG4MLFDSL171iLyUmTMCnoF8
eeUfRA5CKQvOsU1aVJ6lKmWU/5pVvRqLTSP+eZknfBs=
`protect END_PROTECTED
