`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mz4RBP+I3B0QWnHi5B1fR+GhVBfXC+q9/4MkIPZR7PMPa4DLv0CE5TLU9+rb5AA4
nG398hDhK5Q7XYtjKzhLs5KHOnmdQQXVOwt80UgInx7C6ZGyKmibxxN8GjCgNQX3
cUxasmF6P4Qt9OMnV3pSoPJccvgs4B4jlh7dRCiBx4Wxz8cRxMX8akXQJ/ZTBISl
sKswUQE5rPLyXUfcdQrlonPv9cpUkv4YoVFkkedwPgrYWNb2HUXssO879HaeIQ8D
ozCYIHmpfUg3o08UWuM4sBHsvIXxdBfJJDIjOtUuvRgQMovsOXoZpmXzwngMCID6
1F+mU69f635Bgn5edggur7OCMLRx6NSzU0MwaHLA7P689mQ+Is7aIsbg/9TSCHkd
5OqKY2lbUZu5fU+b+Ue9GA==
`protect END_PROTECTED
