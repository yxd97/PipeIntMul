`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3Lr27PgT60ahRczbs2Y6sB2eHa1FcQzLSAo2MtyWvlcH/tGpKUY5XPuzsm7s+7x
THnAPJX58WC0VuvK9AakZSVgCdW6Dj2Ab8mG4gDB57MeCcjXmXyMNsVrVzoOU2WH
ab0WFKr9Jk+O9FUHw6+v6lEbo22DQZ1XTiFcA+BRRnPjDjPI+caz2nN9RT0t7FJi
0zukoqZGPOyOGrOxUNkzfj1ilH3DEd3CDykj52+b4wxT9uY6/6VTKvzv6Ag8J1Z4
x/ln2s6tS6OZUCg+5HJLjA==
`protect END_PROTECTED
