`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0XoDg5VDYKhD1NIm7mtHujbcdca0JqLtEtFvluS6b84igjVyf7MFonjeaqjEuNT/
4aS/SXLebscWf3tohXN0cS0Sb2+4fA/Xcd2QGYQVQ812fobtF0SrVTOaHOSGdN1Y
7Ll3888NyM4KYd23kYKyINCUVOeN1uPyH1ZrkO3loIxeapMRFT1qcVE3baazfa2Q
Ewt9nP49ToBXf8LfA/LSMA5/PkE2Oaa6iOv3oaNWKYr33emW8wy0IJMWEtrHX851
vjTzKjpyTFj/gmfMXiDX4UKUfd2QtiPA16a/3ffv7LwklXyDTL2DBLG5J6kg/tDt
6udq11vS9zJ62+H4ZilxCjfmT1FL41Dy95SW3TEqa+zfneiy7dfDwOWmhPdKplFz
1hzVfmVNmBLFGk17c+Hw92uwdtHVFQgJYvmBk90LfQAP/M3AcmD4Z/Wt6+m5LtZf
mUi3ZPukU2nQ61EiXuAipvdLFrXskoWY0bwI685E2FNmu8Tp8N49xt6Lj/ltWxfw
MneZbxhGXUqjZHI1aQiixUiyv2f5S+zrHBXikmuAoAMuKsGl3SgpnB/e6Zb7vdoj
tOvIXFZsodnNDfTyP7IbO+DZikQzreT9sJDXOV022pr8rQrKJubzgqfN2EtlJE+K
OShVOTVlk8IKnSGx/3Kx7erKq68uiliFMapk7TnxUhuENddbwR2U6sh6MlFBWedI
u/GC3CNDqJw/3IcVL6u9FCVtc88HEwzcIgUrJ9XPYyb+PTzDJUxBCpcmOO97HE/L
7Xxjk7hkX/qR8yIGCQ/2sxmZ9WZB8pjW9BnZSCA6N5pWYBNiAw6MPxZR8OlsRpYq
Xt/J3iUn+VJQNDG5AcOSgCzc5VYTK9X1Y1wMXIhcFPztkUQybq/KFe+8R4uMilOi
8Itdc3i49usQKWBtttoyeyJAMltPhsI2BEvTwa4vtp8DgQ2FqGefY6ZyeT+lMq6q
AAqYQeFeMPWbpAzMlYmyV09G0TvOu7GScgAY9U/9vP6ycgSkhrJ0BIggTlzXbsXw
WhKkJfdfQPJokKzCZaKG26ySwKlNXnwU84CUW53yM6vKQ8IxxXXNXmvPbJiJXbR3
uJQko5Og7vBY5rNKmXfJ4yDxgRYwPgBYyKrJ4X3Ja/jIU6QzVED/7/3PMutnq0nQ
GAF1RplbWI7MRXkqWF52l0SR8f0mw8LieN5WnSpDuRkxc4Pk4z9NC8RU/x0YjWWh
ICudTkORj+KHp6HWgosCf3JlRSf0W9TgEvaAy+uy6Q/2SIwhgOHmFB6KkGwH5KYZ
w1aZQqfQoiWm+aSXVWKpCPVEhfKsV0T0EMEYXcdfpPw3aeOMawTaJwjWI80dYy8+
t4jJGXILEB8lGsgUaio4hroB9MOPHJFTO2htLDxW/RagrQO5ppercO+V+4vQ+3u+
bogiwrL/7C1wnit3cI9LiFzBCQvPjtcLW5nZZHPahDt2SYeYf34mC1EJPDCpjS0q
+mw23H3W8vf0E3o97ssjjJY7NlAWfiKmI3rQ4tDhsxjTm2VTke7JygdCLm/YYCeL
aWzLX+ZZ6o4vCuNzSoJdJZctt/Ko864xmtpICXytXAv5EWTqqFyZ0/4SdG3BgmJV
CWyetFUQLIzkdmJvYXhQeqR5GQCFv3V3ESrEEnOWtz8z8SuFvYSVZRchG4nA8ROY
8ZE79H4+9bHxc2lY4XJepeZN8HB584XHH2Mk4MUlxMrDMB22oPqpSmggL2h4qomq
ZyuvU8rfvlEkvaXPP3uPo3sJT+8fD1mJyPGEwsxIJzZiJii79yZYugQFOjoMeWm1
jhTehhGpLzW8bfvN7g48O9Cu98hmKT+0V0fUClQQxqyjDJmA8kFzX1TnjtA+L/AD
CdzRWQozh81sz6vf4vrQc02xq6Yp+LO8nQQfU90jM4JPV3tUpZ2Y6nCsYD1/yywN
WClEDidbQj+D4wXtVCsBBGsX2XXJHP0NQfwu7XqBmfVbYI6YGMraEJg8ewJYrKEz
Mg0hjDXRJ4+TbENlKhUwVkySwu1uCOVdaLFpZ9zbpthMVZjakLqRf2TmOTktIzlx
BlyiM1NMs4gDvurXlK+0vH6Bz14RQdiqr4DTV1F1QuQBR92TgSDYE5S4plX3NmN4
ZrJNKuZLZGODShZljQtqZkFwbD1Adt7u69Y1RZ+Z1bNvqjWdUHGvSIEDLI8Zu2B6
IrizSBS0hGuUUjFweSolZrquoujYEfpywa6EuM2XWPkRaDwbIuHuUGyG+O5jY+SM
gMnBwAn4g+8QbP5qms2kooqYYmIKK6KzWJf8KWftqWFvK2O9KJCgLAOlM1w6NJv6
YxoONIWjlKNRNiRXILYszhHUveQ3Nbwh9tR0cyG680QOp8/GhZrxME+H0Q/84/uJ
y+JLz/886WDdc7y7d6JOUW7FARlycMPvSh5mzpOBWBiKWYWaRL22BycRrgKw2LVd
WizWhwHbLt3JfSy7koiKvoy6b9oGNDpBo7ANGLiZ7t4JpTKtw3TOsS5IX4YoCnhg
/YOyph7ZrcDyFf38CHM2H6+xN/n3QP71oeIpJ44Er4pJJ5tQeWo22F4qTnUBJT0A
aScRfjruFHl56zXyajvX/0w1JKwwWPgY4+ETBtcz7EGUq+CfGOSzlwns7fV6ro2W
HHr2Z9ZIXuOzld8iVnvngs+yrLYxQ/ZZRWOApBxoALCg+ni41pVYmySxNWbev3ky
Pq4ohx3J4JQWj2Yb0K2o0baTTEZfNnLQgG0+vJFfaCSXPqN684WPEP/QH0aKG/4w
ZSao+9lrfaIntrhJKfKTdhqpsv4E9TqrpC1Ligg7F68hT+0O16PVzj7amFIRqm51
R+G8MZXZzoJBZDwde5sdXTdb3PP7Ec9OkGk8J94Lfbup3fGK1ABgwNe02YOroOUL
YGhqYmmBw8solSiKx2hYLezJ+hhnbc54+5RMCUSvZXdYqkggnfCTxxBIzY8xYkW9
1iL24iFf2QKIub9OVKH0cz3If56AyF9tQJlqAr6pcbg=
`protect END_PROTECTED
