`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mpICsEH6PQ0Y0PUm7g9NXgKAhFfKMTKi920f9dRSPwffSOar4yqQ2CBgDti/17eL
I/GAbMeH6BzVuYjFkXxKAQm99OMY4osWTSMDI0DYirPKSa/AqWABf7KmJVGWMmGj
rGWH85c40gj4tS6Mix6Lww23IoQHaLUFE0y//rDeaDFLPTt4dVOOEkYRLXun6ToF
NHjuT6stlTp7lYFCBLybYEBjMITd1U6y6mSijWHA22ka6DLkCrEsYS/NoCNGygv9
BOlPUu16Sy/hrS9HQVJwFTw9B+OIjs3Ms3bc6EQ5OMU6LDi5vOT8NQVgB9y2CY/G
u6cfQCvdXEBRJnBU6R4kmafiV9hjfDPVBBG8Z3n3xBW0BMKl730ZHVo215fdrwsR
raQSmgfwUEiq7WyUl1z3mRMcWzgD4xkjqjAU2tOpgdoOk+yobVvkPMAIedoQFyzd
GZi9ESjTtMg81bPO2nxUNjtpIVf1YwfValBDMdiWQlCLugQRgU+WQXUjmI6RDSyI
gvfkXB9tNa/kSPJCt1kKC7b7VxHvVhEg2ZbhGTjDj/wWSa6CUMNCJk0MCqCpHjk6
oJzkUojHEr8WOmMp3un6dRFWMICzkYTstsv+09RYRHUzG/4XL/4UFnQ+NfgRLgUI
A5djeSJIYdOZyeIbB4HCfg==
`protect END_PROTECTED
