`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nFsEQAKZY2BkwrH3ycWkpGx+VNLRzF+qhIHobd4IzufrMfVNkHpfqfMHjLBaqyrj
2KjrlVnkP+/MPOK8d6LTpT/U4ez86KfRHS9ARPPeEyqNae1A0iOQwSkvPws5T3Hf
ypzQ7XwV6hNIxcysilUSj3N3wqb3b5E6eeGVdPFAEwuMt5rqO9qhg1L7Bhtwl6sO
p6N1xyQPruAV61JhCXp6rF4RQ839C6Zg88y5d4CHz3IqcQf091DckH3N6ITKzTdT
Hw0gTxQbx1lh5F9FDIRkXtYh/5uNNtDaL8M01p1gr7JHmYsEvz0/0g3fBOdEnEyY
Rr7KauS0sRN9J9spvC5Nx6Nli13T/94+jpw+Ekqh0cSFfyHGQVyYCRLu0pZsEuxW
PEv3L1GugypQM/75FiXTeFMkMIn8W3vzF35vYkVsRNLItT8sxK0j6kpvjbkqhRY0
UEteokbbnQGI6MbsGjHMeXpk5kM2kOw5SKOpiK7ElRS275vz1w5x2dZXEobYWvFT
MRfR4naAVmMjpRaTRGpWdG8kh7mFwM9E2pWiFhs58SqRoD8Y19u3z5Od0tJTwJES
wGMS8h4R0Ny9VCCWbDEA02ZJo2BPdjeYLjNDX6H+xbRl8WHjI4mEXGA+NjpB9LU1
ZuEzohrWYeTGErTCWILMLQ==
`protect END_PROTECTED
