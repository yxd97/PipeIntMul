`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsZ/uxoLP9bsoru3J4qFCnx++uV1S+PT9rwamJLXe3LGA6D896s0YPQe18G7DGO0
+LvYDRHqcf3brudkn03KU0QYOT83h4xKQDYNS6mk5hqN71aqfViH8AcatNAveX7y
I9nC1Rxz4QvWjpUCbE6aUCISiS2iE9MljkZ0v4mzwBXqsIb2bEYJwuUrvSaSkVQC
dQbL3YXFgKBPpIdcyOsz9pueZGmUwjdvMmii/liRV4Nz7gavn8Z+9S0j7Z7xIctq
BO/0L5B9wiP/m4h6IN+Hj2EAmGu5wyeP91CLr2ZzI+CK4N6YYSFa/M32Z1MLC4Q8
+j2FJavnirysqMLs+zNmaC92wkSah/A8mtBqRVT/n3qD/nK5Ar6JhWroLPyeuQfl
pHbMJEKlQiwte37oeLspkKxk89G1dNfKQoIDgOCpOUXKS5MksID7ZB77IVP/UWAf
ROkKM79msPSv+TIy2JQjG0lbtQrnR2YfJUsSd7GJEIZXkWxiSMUZENvXwNZ2VoK6
VMxgy4FCvRz+9EQ5O2whxGh9YXoDYAa7cH3oRw9O4kuvQUp+SMmE5j+tX2Dx/gCI
IDdwo74kCVvgFpC6hJHLH/JQukkuMvqMIIAhGdf90scCgJosbMk3fEFjW5dNjpyf
7r91CZH/mJBQl0I4WFqDur7J3OSQhkTVEvVZKwN9bNlmN7JEXaytADQ0EZeBRUcM
TDpaRnBYphe3Re3rtSz7V098g5qUS+0kcK7wOSjQZ4gvkQeV/9w6Z4BaZnNymJ45
5ECJbwp3Z7IjidCKOh418w==
`protect END_PROTECTED
