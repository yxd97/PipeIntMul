`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zPUzjPQ+pL94KmQOuM03gUjkgAzlVwTAUYVcp0chs1jFLh5afB1fBMWioZ0GX5+T
uw2qQ9P9wKTdfEPHic3l+wUEzGG+1X/oUYRVyT7B56KKYVLkpqDnXJ/OhHlQXjd7
1v+WRWatCOFZrIZIs+chNApS2jo5GNfrzQOA/VKZEMKpTso9py93Fkgz2CqUyVgU
S2a67YmEqJaaF84Qkf9EekH5kKHan8aWn05ESYMZb+uHWa4CuXESI9RE14pdD7Bk
C2Ncyw4mi50+CQNg9/iSHzdhXC66KW4zDnmS+7PFlUBmpRzjUsqx/CPRRDpHkR5l
ZSgvMnPGY2avOJDo/E2iM4kJqw1cokJIkrtjbMfF/Nqh5qCr0k26k53UUwP/Amdh
y61fIiJkif7NY4vAoROLAC3WLoJBnr/xCOOVk8pZl2YSNYO7ayFDevNvY3vcAydf
ywFmuoG5ByMG9vsn2A3m5+uyLBPf6Z+AMMd6AR+RLK0uYYFgwYICXHsbv5duCzw/
oKq0J46XBEn3qvWFzyjBgjit1itBwEv/uh1JJ2aP4vKX4EIlMMTJ3/JmKASJ28ls
8wHyaqxb0EETEI5tQgfJH2foyLzltAfl6NMWbtzw7d32yAqv4fwo/smNXjZRIzAV
cFIA2ohx4HTPJzYXu1WFl3a2zrWdYXYveiW15wky2c4AY7cKOt4jmTWrr+bR5Pxg
zvCX807mDEqjwIVLcyCjoHLnKmvQH4PuFuky6wpE8i3t7jV+OGAWwFt0BTX7OCXn
bX+O9+MDoK26HTQJchL+EonbXFXvLZBkPq0DiegXLw5twLJW1UU0BftLw19T6/vQ
1jAwWCgdQXj6V0uTUuuzljMwliwZh6mqDM7i4S707/Awxfh7qd/Hc+N1Yuke3Vy3
66IDoEZR135mu/hMdqPjDIeKpO5UzznGZW36pZJ7HgKCmfEM0j81JXDGJjCgpJh5
j1APbiGwGFCiXFZ1qWxl/ZKaIUbrVKnBzMq+irVDoRmaGbPfmwCma9i8yK3ePQkU
8UxVP3gGuTIvQn7BHi02X4YQlQyGEFsx99ChMEMKUaFBFYvSuUqXMBGQKarCM5bo
w4UkhsdAIVdP8+yXIugMdteek84h9eSwPqVVRqVZirx/N6TzKHEzEayztEuDHmeF
F0rbPJd0fvmFVnLLwMzBqZXcBgyl+KtUOujywuKw+ickyinTJCvI7EaMGNNS63b/
CyoSkuvFxkjDQsWeXcomK0viVw7UJe/6koB2iOBjxEpGnh+a2yRRcfcXQWo4uOIe
1w2rBtxV4b9gTjj9PP940yBTlDCThtujWGjBozVdw3eEbOhn/S5OcdfQJA5exqMV
OxQlafcFewoTj8f93pWHg+WYh3LvphLpk6r12dzro3xOFH0GYDkAN55V6vIdTfuK
npsT9r2uMR+XOgJoYdWpIwjUmBwbcvGGx3u6wjGbRuOAGGrlOGcXwOTU0IdTxW2B
GDvpesQNwByrNLydOqYWoIRtrTgtwIZ8mltvMfHPjizO4IDRp/Ruf0zHmGV5c6FU
0GidYIQAAgpsUWAQ78VaczkmnMXwQa1CmPIwpw5uqPsz533CTw18O8MRrvVln5Zu
mpEov0VsGFe6bFN0RnZ+RWpPbS67hkCggGMuN9b2TFB4kUyzivFOm1WNn52l4sFt
NrJZzwlJqS32vflKFCtzlMCvm5sdmkDZ3TKwPgEOfUfTvB21fOtpbxmXN1S/dOy6
yM2cu2a3nIOSMg922hXfon1hRN29j642ItDuwfX2uTx6E3WoMhrI1lgnt0ZAfOq5
612bSo+ak20doODdfieSyltdjOkQlQ3RgevrUmlEzjhRFWXJ5/LTtl3ms8yaZoCW
TtBIeYgdSf6izEHp3CiElIHb9dbEsw/DUULQTcD6WItsinWreL/ow83DBpzSzXZB
ExKVf0zRk8a27YO2YoKuqIr8I2Te3bd9OvlGqPcH/cGEgl/DTf1E1D3TOHEoPsww
erTYnFlUHpyiJr63dBLhrqO6pQHxijIigUCcgEs3Lfs=
`protect END_PROTECTED
