`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zpJWUhlnaWdakEU09m9z7r36evAStL1uvq/jn0QeT7gBwvsdTYfhAxM7knkvy7g/
UvAGKrgqcih9S7hrCLdqZg6T9GUi/AD6fpU3Zk1v4ZhEh4Y1p0ZUyhq43c2OOl29
3hCphClkjS7BrNG+HEbJdWlU+i8tko7d2PKyQxpJQHT/G1KyviXSekmQiHRfQlZ6
zJlA/l5Db44uQf4TK/J7SqKWCdqtNFErX+aRp2V0kl/XLxMm2k9dF9wdF/ByLE7t
6n2Tlviqx7G5WhyCRn4eKQYzgr0ZFRMHwCvjDtabAKvup/uN3yifFq6JgyNqZyNq
TXdNSnE1Urzz8qfgoXr7cVN2gYWwVIpqEcb3k2Pj1uo=
`protect END_PROTECTED
