`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I1ENem2T4rAP4C5dN2af0RCWqYv0SWApRuuCcOcOQAc6rsNedyvtLk23EGl48kyG
xa3Iu1H0EAeUzDMDgT6kO1TAABUxySKuJZCCtcwiQegwtxkK+0Z2RRXvl0ya/0cy
6Qm0PPZXVWWr92tWmgExW64B8ecTqKpYk8/OoDij8sPkC8pO2HsKRTLzP+svP7GG
MiI5cCTnSNC3sJJVhxmRQDPbvaJfksSV5IZUV4AQEukar5+yxIXdr2KuJ9ZgzbN+
HjFUZQAF8rdjmMkTbsRw9jPSbgIuLwERWdmBpmEIcLuyrFJwca5MWznbQ5KKgPE+
3vMm1HWn7lXoYS1sdHWbq8aU0PZF0VuNFHPEGll9U+Q83GDSPCxSyqPg9BVTAIMz
7aVlb70aNd1/quBL+CRLWB+f0DumchFBKoijtBiRxQYMcH2li6Bj2+J8mSDkFQ1W
u5wTEoxGQJRctfwu/4eBHBHnGpIMnuQ8dDw6ozZJunI5ComcCrE2fdf+qvgEg3Q3
Wof/9klTXg9nC7eGtF8aJts8DzPmvB6GCxTyNhc64TruVJSB/kMIXaDFoLNPpF9u
yn9aCin9WHtK0rAM8/3T4r9S9GQ9qSNHje2NlUsG6VbNzYWv1h1S8qefblMNRZRT
tL9PCJvxFqFeyjzs1o0yLwOLuSGeKtn32ZArRfdx3Z/adfu6aEO1HNnl8RqkOsPV
/rfR8Yqu0tgc3wXTPXfS5tX7ehoQBqXAFZOQZSuKnIF+VoMLzHxJDf+jrPfK/rL6
Me9RTm4stDUkXssGQgSOhgcW6Ilt0Qm2NLqxIFnHgNN9dKQf3sFLi7izkfjnqNgK
fiRJcltgwm6zXDSDFLvySEQgZKY7pkWY+axase6/Mvun8RagmpVmBD9wJ9nhjl1i
82jZwbNk7C3sbVPslyE4sGXUYrj9iitfrVcgYL+l41oGgSJ3VAxBhfJYLO1ttZ/v
MpkUAbOIDDkLuIWGmSsKFJBNludjsAdwM85ebumGVS7eLmPaj1FbmalgYh4hLouL
N46kQ2zuc2tOWTKiUcAa3Fc97iOfv37z8PJWeIIcnWLjmkSlwNdkqZO/NJPyO8JH
qPQXV1jM6Su2HeeLzjHR1Wexazlk6HMJIc1AuacbpR7duNciIYoUohN1snk0qowY
KBUDnbp9eao1xeDAgoEJjNpN0tn3Kt8UG2C+84VdINntT2r7Pe8bz/fe4h5wjHi5
SDcN98YGLgiYF7zHUTtsl4lolWGZg1bTEpXJLT0iMYINfCu+bX7sbGNePCKhIv60
gWSEULT3VgcOMukULSZCSLoqoLPXUamHpEjwQRCaDd6E047wpoNw/K6GcAvwKDN2
N4Q+6dfPI9gat5tY6OzBbiinqUbUzA1U+z+X/qEiioyDvsLmifaw03wxsDDFwiRC
EhXgi3iyEieRUCJA46RBUbfln6LQEtn6NP+LIaYuz7R/s3NWJ5Q51T171nLQlgp2
JkYGRk50xAvTnhs5vJL9OBYtn0HvzWsjqp38c/i8e1+nuRqn0Jxx2p4DFHBD72eg
kdp4GYsayEhsUfam+8g+wMIBEe671Ady/3RshuoPZ6N5pC2AY7ifaMcccE0sxn0B
aXUe484NOxRx4Hz0ggVBjdatHeJDQHaoqgXM2hizcRilwVbjU5vOqAiJkZsxuBth
lAoIg3wCQ/GMZJpwZVCsuYAkjr2SKZVM5e6/m0baSIOiri5ythOdvv51Ii7YBhZV
W1j0LbUwTQMZ0JHY8nfmYfzlZA12yFKPTNaK+wtg4YT8ZuWWIQoq8GUfKWvw8bwd
s0FBxkPX+b8vFhM1xz1Z5qEA2tBAgCn9PLaeeTxj+GN64e30yvJkf96i+haEXAcb
KtI1d1GhI8aEmkwsl8bKYC844oLGdifPTgCGyMPW4AXUFpxWPiZOjlajSmnu4qjD
BNzv1rHMEcrsvyjDWvAAS1WzEegNWVhUY4FQHjSWkwqwYAEo+DNKrOap0SEMqxWu
bIYHarOO//bZ3iYltWYrZn9G/ntzDj2qyIslPKpTYDwxEWZXYFnEaC6GsOK9c/OT
AqwPymzTPrc0WFJROzdz+6gON9aYZ8B9nDXbmzFev7Mj1tm1zEXNcWtwPNnpbPaG
ru7ehw79M4NQ/nM/LEz59VX7Zsyob4pNCsv7bLd9FzxULHz4xncsm6WkHjXS9hBV
n/nkAGjbn8q3okEZ7TFPV2CHOI+Kjk4ylzvno1+GR9+WLZknCdW11kdw69qb8CWj
3TdjekLbdJUfhZ9ktkc5FDmsjzu6xjUGTwDHpdkUOaWXNyTzLue1hIB5VRzgqyc1
tA3S/3G3E/SFvo37u0KyRVXbCLY9c2a21w7LXd8Vq51XE+IDBrOUDjO7zMXR64H5
ync8UcdBMZDuzVTyaSk3eV8758OUCJQ8xjgsh30exxWW+TIrWCt9/KnwaICRmL5A
SsBUPQ5CrkOtu1tjmoUI3d4MUR1sYrPjeWRGiX9F72/ifT05Nx1jgIkxPZ4DoL+q
bc8k8cHwYQTaTXHQLKlwZ4I/XxOhMRpdC6mkasgOPy+kb4IqmmR9U6uGoIX94i0y
gTpUqq+tpHn4gWx3kTIkMwThJJD+jiBoMljdl1h85z72mIpoHj5cVudHb4HecE/4
/J/qrfiTbRgPak1HaBbjYyF4N2E1m/583swSnYP6DlJ09X+U5QtT+3Z33i0ZRrCG
tMmp/ux4lHKkdL4nHNKZZtOql0qhm0QKTRpOfmJlH6ZvsDdX1Tw80joNw/RjqBX7
iLgK0nAb+owjsiHxG8fpDr75WCH/8TmihSabI/pFbTETap7eW+qPaV2wzotmSDWE
tLxZKg+oJSzWbp5IsxJ32NFTV2S6N87CS19MLdMmhorpqiVQDgL4h+xIfvvQrQjy
bqB/kEnBpuq7oLZ/+32QSSbZreVGs70AnlvO8MYzNpp0IYF1v0wzjOKb9yOKSBJx
C8a+930Vd3VkswODr6SqYJiyO2FrSuvULEjxTkhjLzANCGL9SG/R0m0LBtMzArSt
ioD+N48WexsQG46q0v7DRKEuyVJP2Bb+3Yndeu4WEXGIMPDeIaJ0CoPNb9kk3Plq
/+Ktwr/AcpIuPjk2RpHO8hNA1ei9ez9gKKNjoGhjssauNYTWrX4dWwb5yq9CggYS
1UXOPgPeCy24gBs8MDiPH+8CekzHK0R1hY6+XCLEKMNy/Y7xhLQ/TTd+rSKd/7QJ
zFFT+5X5NEFFUPWEHiz9b6cs3b4Rt/nIJa1MvEvvb0soiMQAZGNChM9r0xnLbl34
CkZgX6uCEdltPXwmJO46PxCGGzh1UmnVSln0S+dunSg4T7+LXF4JVFisvDKBkeA9
CuZJiCZPIXmfovFNfh+COWfgwKgyhabqvQePuK5V9Z/weeUUsMuTjuYVMXgflmG6
tKdnY5Qq10W9wzSz7qmNRjB0jCLL0HrAbfdVZAEJSy/Dqv7Mj2OqTn3Pp4+NUIDH
A0aZOe35mmm/n47EMto/43IfDmodDw+SmdHXyhetYpuVZ7ofZXxj4EncJMr4mWik
r9LZL2ABurjQJAg3Xyv9JCv+ChBX1AMVblPIF+ivP7KDRpQ7Dl5yUlKCiNZcYtuD
SB/aOBiR987EJ3zNcSXFWAFr0rEvCfYNG5ixfJdMFpb+3F/PdZQbClpgPtX4lqcd
drX4HpdS2z5DnMKKXBm6qP8kjLGOXLsdFSEKI+j3RasqeyBvDn2auEa140FJKdgN
UyvwtlzfwpsLdanjLIAhOFWXigmM+PKWIwYuVxgKJHQTj8tPszMKGlfITCygLO99
TgArhNaDA9oKEpifLbyd7Jw35H/zUaieVDANcR5mwYSeKf6Z5Vax06SFqYtVpscg
euZXFmbnKOtLxbu0g3P7Ebr110P1H0j6FPIOtDAEPXDmlQ2agF5Z+yhRmxo3wV2t
OjbKC6KZ1iJWwnfqH+Q2nHgYMuTD07qD6UNwyVqRnF6OV4yKweW5vNZ3kZ4V2EnE
qhvY5Bc0QU6uYzWcyI5NRAnQ2pXfs9lBoI3L2eRGgLlUsTdYUcFhJYWwirvWhT9D
zcnwuhyxoyv3UPKJIFPvCx5lV+r9rFLZNh787+BmaC2d67xU3ZpxT7y2uhggRGdD
1vwU2e6NS9uCUpGdA+dnFkSlT6XlT3/R6b5QQV2HIhNct0H/K+1xShYjBPGhEwXX
14b4BOON4AoVByfLAek0GRMvlGcjJVX0z7yQbKqxGuRY2egM8f9iskP0LuRo7JYC
vQuCS2G0ZDiImmrwW1Erp/blaHh+TJ2iQo5r/AC6LuRlDYEn+kpu7tqVLXdg+zAc
BQDOuIpR1IvxholDE/WQTNdXt6Uynq0n5jJs4qk96ew9pTx1taS1ABxRjCiwbnhS
EYfyhFXUhQ/lEgG9Zs+uwyUOMnLHAQy8dv7wh5jvFXwaHGOxET+kK1A81qKLGBYe
TdbxyyaakbBHRMwC89lll1WG2dvFBG4ygtXUevy0oBo3JjlDagCAaCWlzcFbJkRX
fpPMCdSZ8rerNQKdJj+lJXS31bGPQ4dHWhXRampFtdXMYQVuVqYbLflgv6BYTSmf
aZo5UG6sS9TXt+1GFPh3CEjl0K8F4Wl/V0Ur7iSLRT4tg3f///ibdCwhUNyBL9i3
VMJ+t/dWCPFpjaTdpq5uCZjbsmav6SI/32Yms68iOChpoM/LRht9NyAAKEHJX2+C
Li9uLB43ZAFtouxieww3/kfIdY9kKBoLBrSpFjgRrmj/S3130v7IyIzgyz4+9Kbj
c+OFMiODOZJ+3GpWTtm1VlK+pTl1Bu7XY6HZocGcMPAD8HIrpVagMOaNT6LSZXHe
rpGY7QzR3jYIdLB+Peb1Y4ltqmKs1de1IgVP+y7WfrchUB0GZY3h753JFUjJ6sOa
zKluHo/6Bv73R2eJT4kATwmBRjfFHv8k3Vd26cidtb2x8den4E3myM3+zRlgsXIK
YCznZqASuiS4ua7i0oWSZKbdN0xmyBZSaw2bPOALlMZyrGuVmrAkPdwTluuL5TS+
QGMeEur3gKPhTB9s33fiyr/s41u1G5f30DmZ8f/KDRStEyPhw7Auxi4xgEFt3zj+
GGl7cXAkLJQ277ktDhNUiM9Sq0wuXR1LUhFZopYgkAYF0TLKdmd+XnkO2yggWU4h
m+s9XTIiN6hmODH3GRuZq/pzR+vO73DD9XLj3RDAseq/eI9/TEc3nMZTJ3HHK/6Q
rEWca6qZT3xKbm5rjJYoltp30MnR2O517n1AMB58VKHiPNzJ8a8rin5Bou2VvzD4
z2hjBndZoxO595qiCPOGqVJJEkU58QKZyDEnXSqSOY/mKTDT/NYvPQ1kjWuxrmBn
IGBqvcVYf8bFeV6bmqDEFfSKO60YC2GlT7hBrC3MNeMK31xgk38ex6vO22JKuMx8
YudJC+Aty8QRvv+FxHcNFomUyOKPYNlgZheAb0C/G8UN6gz+se8TO0LfQ+1shY0C
6lNVsdrp5rk/RVRx8gl2bEOCeZiwMpJXWOSWJDcraPHdkttfiSzreIXz9bkepdfF
XYZPBoeq+QlkHdS6WTv3RSYL3snWmBvH6dx/PvI5J5FjLLx6w09swA3iN4H8VjKA
K2xrQIt4OSel69PRmgbXFPQVJr9eA5X/yolIbsGrbuAhjIvlS75kOE3fBQ03yeMy
+V1aON+/S8OPgYZfy98ry+f+xwZr+m7xEs+g4agyFjqAII36zWJ5e42wNXSOseM2
gCxcS/sfg9y40ggnEFxe14Bif6+9Co7wXrpIJ17ufySAOn3riUH6IjVBSKbO5s+g
APTCm/QwnaJC4SsVRB4R9bR/Krkp7tRw16+EfZ6aBOGdnMvinmjKehr9lwoxYN4l
U/eGjhQXYLV8yciSyrDJjzHaK2unbRlOkZb42LUnVeM35WtDjOpDveM8Nwd9V876
+K7q2zcy+SvmfT1POpE514116wiucBnYkocSblZIwtP7ZKB9Dj5dh58QvEKnwx0M
krHx1yf2iDb/2o2qhVX6qKBrrGWVFOL48jP+2OOMrCV73LSr6/LmUEyZWKo8NIeo
zag+jz5zIbAU3uCwCH6H8J6WDHDD1d9mUNqtmOspTrgDJgymAblaqv8STp53z+dG
Yyu56ip78yfQ16fNLpH39Eg/gsX+BFavp7zqkeZUl/Hp5juWT4/ZneoVcTi91p4Y
TRlGt1fo5j8qNIqQEdgmU6GfifcFWWyq5K7/rp6ui8YhOyKEEIsImIuoGPOVQoHj
eXsm6I8Rh84NuVSgg4OcH1pSF24QRQ5rAlUtTOLOuH+uJbZ1JtFeJ71kHVS5fQqD
JqCw9FvJ9sRdGj4ihdCrvPwpRWnRGKkuZBMbtoB696VWjUdxJKaZAv3G/neVlVoK
e9HEe5DKzRHGPzZuvt0MHOPlq9jMsaDc35C59hcBccfK5MDnDNGOa3aatOGM/C2t
qvA0EBQff7YOtHyqcQ2ARidDzlA6mNsi86FGWfgtRn5UqROClSFefGYv6h8bkpF2
Zj3k1WgnCGInHtAtozpg5jj7LBQw/t5eEDQTJn6h9I/UX3SVUMtIXPOSPBICyhLy
6FVDVYJhNUHuWPxwuPowlpM3VvMatBSAKTvux/dR8y0sTGyIH9dNxKRC2BhKl2bI
SN5d1KW9XMR8Ecd3uFoNuhQA10DXOsQWkNjiDGqAkGqiPLBQNXZxeD4joueEn9lx
WpQhAb0MOk8Id7XycNkh1m4FGUuBNfVq5aZ67B+PGRfMQNdvyRJQQKCShU6GPT3h
ll0/Bjo3ftwd6K2JDcsSVKOLYFEnc6fwXOvFxsVzh95a1Q4KwoVkyzs3pGfgxt0Q
UPSQD6NL3toSvk5VubuQ298DhcpDtuG6bL4sNsC2eox3ppb6yCx4fu3dVZP82ISW
r04MNwEUKxXGC0VVaomf6sdBjqdafb7EhorsyEIPGu2tMHS51EwiaxQ99pTVPCmC
51n7shHLGZ8O5A+W8DTw/bRVJvzINoz0GGII+Hl3W8I9tw0WPZhfviJqliLs+1WE
icZN/ypB2dRo/m0/rp+UTrDVI6dq0TKxldtxPd3mUA89XIX6lYjljNWdyrV7UGaa
xLA6amN/C/zKK6fbgWdxIMk4TDH9mylnpyiWEdsWhqck4rfpnG7XcSsmfsvbvLFn
enPgtuYT8IoSyZ5XViVX/UudiJ3e/VpinrlsGtYyE63ZpGSPbWrCUrQlt0rU6QEU
W109p7A57IuHR/24YZqhnDA2rv2EXu0Hj75RcLGvnXyY0hzQiURzIAXDDENG8qbx
II/t78jhNYsUquEJuPMjmyjzg+AB2UI1T7l/2CJCR6mkaPuRwovvnGCObDxXgk8h
43aTgSU1m2AMdb5nnIqUF9096tMnCgW0anSCOQXbYa+OKaMTdyQ7FlbHmZ8nutOz
0v6USTZxCNNxaMl+tl3nR0iqDe7z83yXewTTS7G3exWg4UkvnMD4XCf2N71h47Qb
E8rppVP6Mc5vZaND9UhDulpuDZG9OynC/M7PXnk99AvL4EhiIs7nmyRBV8F3CSKJ
EEORugKyJf+2kd2YapDo//JZsR0rKqLyAPhNQaKV1JlXWIxmTgcBsoZsMD5a0QYb
Bg/OpILezqI7eIqP24pDLnz/ZrmmjReYyDb5n3xW+JFvsYUEWqgvpN2J0i4WMVvq
rxWaJI3pKUkD6LRhtOZTos5d0rlgLOE68FiiCF9ObgYTQcbJdQrRbuMNbq30tN7d
TYw8jmLRkO5mOIXmyRio0qh9paWGr+/qyWy4HFr0MtwRb8FSOd0D2zMySREdn4dN
F8CEXwyHgoVm3bqrDOFBYSl1SGTlW9j6EW0j0xJDJMBKDzV+crqCQz6Hvofgnayf
V6nJ/0mtaFGMVjanQTzcrxOXpXQKmUvDm9jmCdMr3Pz9F/RDj5Rr4zM3mPaCi6P7
LlWuZ9MW/Y16NeIToiVjsQSroDmzcvANXpcfuyL+ogkfLACVpg0/ARwZarxHLH7r
gwww+LPkX4eGZ5joS0v2oV2o/fyZLidoYe14f7lDWwgInuNJ3D68/vdRADZFgQC0
GE9atMoI953/LP6jN2tcFLSCkwNEzDwkOmd619ukVXqD+vM5KYPhl6t6md3tlKQz
c66CuJBAZ5fyRBuq4ONrlaCQMrgElvjwZd1LYeLRnkl9k8V0IMvbhOl46Y/OoU/a
sgXmV9m6p9uXFlocQzPXV6NNNJiYNNg0AEBdbXfzp6nfTF2wacHZfgopwMuwuIC+
eFtx+GPeowBBOohDixQAHyMmhEFOT0kkx+rYk1r14sXLw5fuPTsm7jZqUsqcAMNj
Bz9AD/JBWcfDVIDsp/7FKRmsHJtRF0FUng93q8P0CHleF3qOGQMOuLpY7bZ+ih9X
FyEDesDjmZYQifDKZtO80S/IcoRY11Lvx5OAUocgZ5Qmzd+i14438id3qm4Dgw+J
WLlIafhqMGAj60NIt7zY40Kc/+kiON9YrTMN8f2HRLpjIlF3Ewgq3de/Ga8w4gB6
J0r/pTSQDhY9RkQ2NGeetnYNb0yv3a+SK+DIA4TQn2PNAeH9fkeswKsjXnqlnzUy
Fza4OTuO9WNZ9fb9N3nmIq7b6an4xYvVO/M8Zt9ANt8ODIAfNheL3MizvpRDd2Lo
/SwGh2yv3C/w5cKIj+hwB6RuNdspdjT4UuZw17nzReVTrkFSfCeHNeqkpUczIyGC
R/IQAQ0WATK5VPPjoAiIhMAhvIU0wVGTnHI9Oe7e/ZPgLTdCrx42SW5TgyeCr7yx
kg2Ig61tVGKldzDEHqEHIbcjNM3AujNmlS1YwKB94QQAqz/N1m7kIAqNfZgVx7X+
PC9Zml4D0nXeTlItpnrqT/usLfUyVmxekZl3EIKNhjc2FN1Dy42gqSw2O+5U95dw
uZtYTjiVRqSMCbtRZb9Do+A3tCmsvpjsvL4iWHzBtrk2ny+1JvCJH9j9g1cnLkOd
HiV4NKvdcBurRBI+UcBVGTiUEGJErbwBaVHfbr2+WhL8RU3jqvY6iviP3i0h+o7J
WDJ7fGXO7XkBKfX8NbHWj0unpLc13wSsEIF+RYgsi499xTpEposiOx+exrUZFDJv
91l+OvbO4DKHWo+lDsGKxsVDldUQ2wRce6DaFicf2rtDBPrlP3lVewg6csSMDik/
Ty6dkLuiirpWzMBaAeUw9CiNKNv0+kZ0GZBcFDYYF0MdEwlbjVTWEOdqd0JXd+Zo
u9g3XbaUmVRUiVmtpe318fu0rx2DQPPdaMKjm/UHMloNzwSGUbHMgiwq8nohvaY7
2Dk9QIvHaWEXliJSZ3g1JbRNYouZOzUvs0scJTrBnRnxrf5CWa+FrZmCmNBmuBgb
Pf9aB/I2j9+xTXyg0QELa+etXIO51BF8/KaepyXi+/VWHMw1R1396EgPTnDFcr9J
WsRiLQ/Z2RaAfUjzHONwyMLHMSWFyrk77GKJMk7/pnTi7HNiptm9J1eI9PNj85V6
6FH/deY6qYo03FsMCtRuoXR3k2G2k5Xlt/TgABXTvLem78fr1ZhnWrP3+Fcijuxa
+mN5aW1dZFTKhOugGm46KofpLqvlYS3gTedVmjaqd4jlRj8ZZmSCEY2MJgMdJ5fd
wcssRpOkomjTFTX+eOY1Dyr+jpkJbf8IQDvRAragq2KTXzu8kJgChqtn3ynmJ2Yu
7erh0s1n1QSgKRaMpn72W2QtyHmdJ1adOXBdDovVNUnnYjYw64nR1vahAkUxMYD0
I7Tu2JXk7Zkcc/yt+flhE7YpuI8WbQmDGByE5u/UA4q/jA/AfwtM9TVhl+RS5pR0
clWAy2EG5RmLqXrjr2UXTAU0V+epcRTgIfPGCiDNt3McxnfFrryjiLNOr6nnNv79
1Rcr7xGBx0o7E8v9CbBbLwHqjwx/6i7cwvxHPA9wdPFa19xWuZu4XTq3N11rajJv
m1hJEW8iUgc5HNMCx4hXS5bWr6LxhqWKZhxjGmFZh525m5md+EWnDszSgTv4hIvk
LkWpnH38aVj5ufPSJG+nWJKZ22Sm7reijQjyp97ofgXdVFpPB30E2f1IsG+YGRhW
573dCEoFMNsX51Syd/Auu3blSuu+sTqFCfCtwyJGPxQi7LGLprpQEvp28QJOcwBj
lcLWj2x4x6eZEypmm0nNe1jS6H2C867+dd55Wlu8hzv9OboFkItPtVn+ZUsdCbpJ
Awr20wM0WUMHeRZU1oMatkxOkZL/QTKZgxy6VX+/E4dU+qzNQZg7S2f7mtvoXclk
hMicLsD+VDuQlFRAtxsNJtn75o5ZdIcylDJtH1a1JvzX2EOONdBbF7LmSrV5/kW0
ofcYSoXJtJLEInEnKoyJi8HoGMGvNFNBJ4urziT1t0wIlvqSXTc6HQkoBWMtjE9e
r1jqZUSr8mwa0exjBU78M4OzQ7e5cExcorC7xkK0de6Kkw071M4ha7/8pm1RmiWM
Zcmx6xs7qE9u8+6pq1dSkAVkMJDr9Ut69ukjUM7/3IiR14mY62dCNrJRdSkS9dMy
nlfvIouEZmI4m3ZFkD03SDJVoLnRj40xn1W4idxudrawfWAIoXObyt1IXisnQdun
O5fhFaD0+jSTXbjnYwo4JbF1zNtnz6caLjXs5AnhUSx9GXQxou5vaxyUwTHTE4qI
7Pz8rhdJ3VrOi/EUjkdjmH17oYG9Kcaa2r8nGJygLJkjz6zxbpGLt3co9CyCK7L4
38ZK4w4ZfAZC19MTC7XmgvS/DKgv1brpGHwKpQ1wLbdH8zBx34Pl5qz8hGJpaibX
d3qKIdFobrl86Fm2TnzAyFNZoeBdij83/ROEX0bAkezFFUqmt3hIWsIPL160AP29
cGdGi+dESxy/0nb7iDOiInlaRNLcXcd88E6debia6KNZQj3QlfjLaN3+VPB+Evh+
R1kpsC1Ulaw3HCM+mUcRNz5v/RfwJ6P8wk5pCLh8Ou9w8Qg8JfBjGf3tdN/Peegf
Bt9XECzL9w1mbZGja9Q3g0E6l5kdfvQd0pY4M5T7tomTSvb/z1afmdVRRLLRwXg6
17+Cl/gUKJ+nSBc57YcQMmqI2dCJjBghVUBt/AeYnkOJ9YzfBOpA7abd8LnGDmI2
Q+G0N2VvnsF+VCGX2sDqCbwxIoYrTgsqIUE308SjtgWuEy4+APwRi/ZII4lX/mNP
N5L0MA8wMKiAAGp5DygxYnu3kKGx5J/eNp2390G5/wlQQVnAU2U5mK4p7Bsu9H9Q
d2tHH6VjYjhFAZjDRLRXdmkygRwSkJekLF9/BFPTzLphc5eg4RKGQ7KuezfjdDPK
h09ndY0+w0Xu13BJjPlpuDzGbdmHGgZRh5JWoc8RdPqUkx3VQLeob+bWh1BkhtcD
4nzc8+WyfA2G7LUICpCoFteOF3rKLwYM8SC4BayqC2KTur0uhrfqmbUyNLik8oby
+bpHBDg8bNMwEKQzk3y+arKOX7Yw70xhMpeTrlEH5ZcbIFKskzM8S2ZqX0oluKl2
uswxikCtvHfAUXWQHmfQpnyY0lHrcLBbaTIgxSPQDPJAel0WSZ4a0d+plqu35STR
CS0OUdYywiD+plXK9x4eCEw3oxx5ezbJJ3Jb0sxAj4dQTMggYTvQUPTGoNiYP1l2
wmzo1DR6GbaRS6Y07uKtpSzyGZn7VYMRdEtNH4igUq6Kt9+xwKgtukSu078QEwXo
EIqk7MGY1gOXnhba+o9OY664MnXnqZ8T/5m3e+SLKiSADf8dceU1C8YU3h8D+83R
p3DhQboAsRvDrckYRlxyV3wyaP1mt/+w9DsP+CJ/GVJizWcuWbhzplXYMohHzfJn
3M+xsGnI93GqhAoatX6L2AcgmljUt4yod6xclpBZKUUTvrY+cIIfLHAXKJCndHwu
0z3BN0lMbhpr3vDFzDjzPOPIxKUTJ0ERob38BWBgH0IMy5zBdRHhlFE1qJU7drEO
OsR/LaTrr/gq8Hx6a9veL0G7a5M8oSOjDW//08oS63rmkF/XgBzbHMTnhJ7GCjyb
bIry28YyAqu/0KT5hNiMSlQdGXzY/zgVC4LXSdmmBgx2+hMr7jLwuZ97qKxCEcPc
lJ5TdqZ9/3fQ7hCyaFE6EdJxYkvSyCoLVV7jaSJTLXgAYKLr5N88cyAoQGaLt/Ft
fq9RHATB2Dxgh1bR2078/DWWOSGTeZbLm7e2X1TN3e2z/ydaG6nR9hIWKGTQoa/C
CEqw/qmKJCC4zGiZ+S5NtbcByvAP+LJ7lpFFs+JfelMHDpF0MMLQ9DKxhm1HWxCM
Eh1WaPQmBbx4rNLz72z6KNBMUcrEnwawdURLmj9qBoiO1tjAzhOxWpp/4JaptLmU
MIjYHXeE/vD1QOowbEo7ZVdSe68uamkm+VJFtSGl8UjabOL6Z/gUnQcT3NE7eWsF
/WEriPkSufn2BaE8n+0Tei9WTxSdy8qsQzDKLRhNPYuLQQZUI6FQa1e2MUDCUL+o
lOkBqtEqHCONwNz7VgAJkgSCIn64EUzYeQMPuUPqGKn66rQ7t0TM3+/sjk1CJ6KI
GJAZD3UtHWgYYXVrOgyR98wZeoPBAVXvZPO0UFagSk9b/EtVm3J8CWYS+Mai661A
QTC4YJD6GSYRkXhRK+mMGSr0l6f32wWv5QdDP0YWHWiZC++YIhlv3lL+jB3QN2aG
mJP3K5jWabdLXzf0KAfBrqVezzJcoQVODTmDAgRghnVA+QxAWlvLNNreGzGMmFF8
jWYUB2192AHtVEZNiuf0QWDfOuu2tDmKnIzohB1P4c+krqCcqnrRYK7L8vjDuA0K
EBUhHLRz4m5XSr+KbYpQuZig/89poDU/W128nx+d54g1+HG5f903at5PTieFx0Gd
ppa41qSVM3reXfoke8MUFg8fRv4y4y1tcx3O+SGprGNgthXlG0WRdePyjHY2IFcJ
T3FDJ7DCTWnlxM4r6nqMpgQYAx+zq99w6urWKn1701jKTI8JUWCWyC8BWjcO/Xip
BPDPd/ekT90KGjJOHjTwb/rvYjrk3a5rJhQ4kTliJlvJUTVo5d3Kcy2ONgqdYQkg
5n46tTyKHPOV1RN+7aOZC+j8XsdZHT7p0TVCfe3XttzI9HKDknMJLw5RERPxZojL
oI/orFkL6ug5D7jdCDU4AC2khEaaIkKrdFry4GcIoag1/3mNTRRFam2H0RFHStOv
MStmOEKJBkq1DmVpuAjgfo0PPZUvKA4G0KlSwTacrN02AjHpV8UH2vIQCFE5apEf
ZQjhoAKFaojB22tDE5K4VzjRO0uEeVAAkZDCnWDFW2q9GN+JAScV7FF/ABrt2dlQ
oHl0lGXCZGrZUrccg1vetYXAZSDicT0KcN1eYv0m5vP/XX2YiLFa5D/16IS5lnBy
pEtDp7O9uSKHsYZ6dY/8NOXdiAv2M9+rvteME0xJNZRLOHYvWaj8Gi863PH01Bbh
xTdpmI6PQAJhcCcA/AgS7lYN59HRnFC8cN8OlWPB3r4Xh72zp8ndNO7vxbPTdX86
iJ/ciFsrM//oi4T+98Unn7/RLncQms5JyE6vpMkMZrAHsl1hjSBEfu4FVjb7abg8
urTTgs70qJCp20MAc+qC30vU6vnnRkEwoHWtGSj8vN5lsSZySKDjF5rH/eQUCGkc
0czoO7hQc9wOcld4v5URsdocmpnZxv2j3chu7z3H1f+F/ej3tdXoP8/Oor2iJ3vH
9KdOmYuLN4VpylcS/wbOvscfAa00KSEKcCgO9UuTxCG7OfQF6rdCtixlKZjYMKMA
X8VaZhHQs/rswWywdtZR/L7Ew/FvCS7PCgdCZglw27JSAZbZJ6HAEHifkGV0tI6n
6YcMH2CrNA6mZkQfG5EXs6zsxXeP4aNlPFTY0vSuIT6vFMlJ4iWwBgkvIYby+yUE
7TpVWCoDcufM/X2/bRfLE9YA3TKmlm36lONMnjld76RPgCa/iwNPU44OfUG+eLv9
OEF4kmFxjDOmaVJHmQahdFqApSgv2p6aIfkU0x32EmBQZNq2mNSS8NvUwWp8CNDi
NhFM9rbFILmxxMD8rmJCeRZgcm27sn6GCmuqa1wv9ERWslEpvs1nr/kjHBYn3Q/w
bpsVYrei2cbTYFuApP+IW//XkGf4x7/ngBeqKFo0rjhMKEw+cDmB+94EY8FRPAyE
NkzNZKP2hwbJWSIEgJvCzdxbM56dED8TcO1797KHJUXQoWNXFD6/Il2bV73mskTe
7aU+6mWF73EXJ+x6qKMCyos/F5Z3Ym52KOufrVLIdLrU2fWq1eWqLWLCardRFqi0
6ZoI6ZEQGKUdqW3//6I/tjvWlQFBQUWx0iQrK1OtmskcVFkQ2EfhdIFxY6aJuqDg
NfPe6IW8REpg7sMYUe8PHTwvq++tri4sgd2HjI/U6qQv5Oi3gHX0KilZ5nkdi/l3
CUhEbmKngyyuZeh8LYt3mTRQOt3CJE9D64BmKsY2ingZLteJJ8b+YDodaA3lHbB6
gygLWKqzFWxmMUHktZttuZGAt7MovYrZh6CVYsUiCyoWOvzqZZqWfJQcuZQLIeDx
Q9/Y6TpeEnq1VMxZm5aojKCSD/JTJskH7Hjx7eMr0C1Oona6g5ow/Fzp+qVMNFlW
fxRkL5IUAKt3kPM93svOiCWew53puCLpukSls4BJCkBAVYjVkaPLJQu0eiBAzOK0
qb74OWnWtZqLnxAnpAbtfLyNsOqk1Ve1t+bL/0ca0pQKXuN5I+X+dH24mUexuZxX
eZTCKiKISti0BwJWBVyqiFi3sHfVmsIeUPji1vmEqyEcfVoZE4tNoTf9dmJWZMiI
tQaA71qoMTL1a3FqGMlDFLYkgXMs2xCaddBBitI0IvJpRRgXKa0jOr/ZTqTAPNRv
CfAr/F+N30M1YkHhlxgQ7n6q/zV/G593hOqKfTSx4qYGyIOHtUbKGWkJVMKmfmc3
GBOi6erB1DU3OmH/htpiP1YOX4pmjIV4+6U4UmvRzxiaOgf28bMusRbtqGhvJ99N
yOdBwg/q7yldNVEq6hg74+97L55ArvD+yUT1CcJBogPIOoPLYBNq/H8xQ+dajlnU
o8EVrmoO0hRdQ6ogMA3OACHz/hmSHQKYuVx6+L3KpzXN8DyOUz79eZNb7GPcmdpf
w12WhG48r+nFs6Plgbu13i6x4HL4QqANP2lQ+6yRrskeRHBdxPqdvUvz3uTkuEzY
H+eFRwaq64PwGuT8O8B3K6t3OYDkrB8CtFE/k0iyFmZL1WtYj6NQ1DiN9HmS4puQ
YT7E03QqhgOSsEPdktEejYGU372pgb/svqyDd21ymS4L4k+dP/vAgzliF993E1Rw
GdmZatKo1ucm66gomBimspP0WSFm35creys2q/jgd3R8SJZB1fSneFCP9rpYjCZE
pHIbYZt8Rq3DPwpoL4PVPdH5ZO9Q2bMfWulfs4zk0FLeIjWj3S4TM9vlfRZdWM5F
HRdEdA9tdTfHtp25Z1vHlEAyYkaiyyXmy/Sl7564eN2+jFcry5J+Pyslzfr4Gj6m
QiymMHE3Sx8Y1/v4RmZdsKXGlCdx1ovL2XZ0ftXG17Ci6Es1fUs+VntadrpOwds9
g7tpTUwhm4itLPWLadxRLt8DXLCuqLaH7LnM55EeHwSron9W1bhxbjm6v7MV8kiM
brYLHLYlXEH7mQXQxemKXZ8LlupW01LGrjdZvCCDQicmD40koC2yU3TqzfDKXknf
MXm2g+NvLQnmC+1PDcIpfZUcO4tLpJ+qWJk5YuAfk3XvLWquTrMnkRvMWsAPlgAB
u81BH5fQ76QSNrKHo8G2pA7HKm6HKImPx6QctFwminpouIH8zSqtaiNRKMARx85t
eO/vJOFL30sZ4iSSQX75j2OoL0ntdxhb4rUp1NBFRHan/FF2VjuzWV9WDINF7S/7
WYJ6UxNI/M8HjUeIhyIlrc/bbvPGCX3eFECevaV177e19Aon+gEzSGHeZyq+Rotm
5fUMfCiJqF/KqonRX5eCfHUiErjRsyZscbsTEi3H3HxB37tqTfTYvqAptAcUyG+b
EWJhr5fnEl+Xm1UROM5GUTFJDl9Qu6GjB1qUqS9oDD7MUxyarcnx0aiOdNqQgEcV
wBKSM0eU+hPVdO0iqMPJF723D1W7XOqxkAJoLdrQSeeug/gb8uLhe687NXx5kpyk
Wj/1g/S69Xxdsn42lnKRLddYlcbuM2tuF7eQBGxQbLIy485w2f2A7qqFeuuxX5+e
zIYob+8GwqfPKJYgZ2qH/Cw4EEvF6ytS4wBN84eA1/NK5C7D8ClXUveipNwJG/LN
hn50iCBg5KQ1E3c9grtNeYADYQQjmgJvp7P7Vr1EHv0LCWevRedzHICzK1nCNcUF
Y2sm5iZ7OSHsuGdMoIIJaTH9Yo+Ee6a/fFmzsrsFfjZS8d4p+UDgwhkSfGiqBBOV
w0VpTw1fkE0EZZeZub4KFvKRykjegM3h62xkFlmrp3JUCJqK5g5vDtcAzOwXnc5f
VLIg2hn9a9QO/cfubmuuUVrglXxub1jXZ/NeIpMcKa3/5fm3rJ0oUSHE0d9Xlv+Y
DOOrg4wzFAf0o1bfEScYauTuuFnNS8NlP8RXwsWHA9IZTF7TeuHVWLAuirzWv8m4
FZHkNqlfe1NDCHditGlLqGxX5fDNXAMDBiKejqX/f2+R7AlwGH60yvSrT1SZCE6g
QVtZxDsGwdKG8vLD0X4u2wMv150zsKJTd5UI/uCfCaCuXIrTkCRhWK04igC7rImC
EZuFKJjNVHdEnDaM5+HsW6cfdi4e7kjBtidc4PIyDCmC8f3zKENW+RBEMAoYe9UT
BKzlBO+cWSxZ1Vb5DIiyMgsZHebDTn0RmQk3t0jSahnyOihHZNvPIQcA/p1q4mTG
HpeEMcyHj+ApM4r4KsQVPIL3c26r3jA9Uw7X1hknq2Gv7+FNt8fP75zaZBlMlUad
o7Yvtd8NDp5+JZ//1Zhp4hQBwJ+kjU9kXQnLUWJk0v7UVTUEEXv6NHzYF4BRU6MA
p0peDqQywYv6ARAne757thUsgYHpE9Cw1WCd5MTJxkskv6PStsbzibWzgOme4Lvx
wbNkZMJBeMLzrPf3844aNod7h/U8ruQZDuCZxO6ma9XIA6nJzZf6cleTdMu2rKsX
uLy39LT5NFAGOVHBm7q+zKSNFvGGCnugKJzwjNd7FgBwhJMeNJ+m/Ks1LIkvolcZ
4oTS80a4UMH8dUcNznGvS55TOP0nQ5OY+BPV3HRX7nz2nHVrSGhZ4/crNToHskNU
dbjpv7BEwDRzSfvNFb44cwj5fJyI3J7Z9IRVICSEH9JkIPKiQ6Kfd3AkDsKhYXY0
ptg38CLk/I8AIdZuggUUW2ir6Ze7POR9lqcDsypUVxoM2BXzwqMq478ciuMCP2LE
LO99nXHYPfwefjp4jmwOxorK7l6CfjVCVHz5pLhXl1NppCoPJCrTyd9TiNPo4Vap
f2H3ZUN6FAd9JnzDWGMHUkJ60kK2bM5E/5YzqSkqNNjsQkTaiwJ0YrZ2Zu+oVmf7
E7elR260woxiGhS7Vxy79OP44koH9bCxYTceRgkUEa9w7arp/k1reg6USbfsMl+/
eF2BtGIUad/oa7rzvetkoC19rb9FayCXhzT6fvsxNksh39pMV5DUNNsBJY2k55Ca
f938/rmvpG/g/jHP1KAJ+5bzjBFdK5/2Cp/ZfLdCRUOMc2mC5X6vMOZez+Jj/t/7
CgpfQXuFBYh3sXVU29o+g6eZC8PVWCsN8exesyVBHZpeIZkVFmnbXqloHGx+SYaQ
aqtuyBohLtd/kK9yYiaI4OlEipxzqfJW58L03m1R2C1Ctc8gXoSz03FljRF/ydAu
aVKQ6hAgVee7g9KZxysktrdSxH3fok64MSjNdrt00uUHIQJNRPkGQcVqAyDberp7
kQ2EptfVobKIpYzL5E5xjuWCUfDoHT80jXnQjMH7z1bCD311VoN00VRzloBmPnUk
22Cgz3nwOMH2QWMLYhxGE+jaGwOx0PfJ9Z6Rn6mENT9FQgwf9Ec25ZjvIbYFZfj1
p7HdUfQ1gONVOyCRCaVEdg44O15Ajx9p0lTDDm7Jo1HQp312FEPKdmwvLk05+ifi
WdGoSm6Czx0rD6uflgApHuHiPO1enH4fLzdv44jVWqdTUhW7Rg7dyUCrsAcqOsWs
YK8xW4589IvVJ60dlHUj0nol0xnLZhCPj6FDLCK8rhTULSAnKokmJZQVv/BluFCr
DjhkHbYz3dtfX5XjyBFBohVVQQeJT1RNiUjAgESOFFUd4Iu6xiJ3ug9hgoAaPO5B
sQxxDhbvPdRetVC14FY17oHr5qWKNTdfcYbmkhSZAkR3C9xCyhJIPq+EGAZe0Qxu
49RlONzTfHXoYol1aufiqXLv/MoO/spNgPl8s+k/2F/p7RGsig6AJvVu11a87lHs
rVecsEMh+VsKI3rH5fOlIk5tbSoLbxN0ubZ4RMFaX/AX4Q8TehPbvyjrkxnmpCJQ
kIldN5rlyvgtMqQnuw9fcEI1AdnxMReL3A0kVqcOsoHKvpNXMyflnMt+VDSUVERh
G2Wz/lEFEPMKgWd/pYzZaFFvZSFftj2BEkjiTZ+UvO1V6A/yCfRpr3Hc/VqC1mSi
COPCMU86niA3OKVNFtdM6gFZ+VposPLEZuBpByMau1R9Pmx55yuLLqo3bwfvLOQU
EfUl1Ol7CU2n4GN1zQeWLj7pc8tkjzBq4fZFSoNbxQjikhEumj0tUidRWkb4z8cm
W2xg/yAXc1gepJ95JH31S0T0NEy3ktiHaYUb2Y9AwoLeb4gBT2ToMvKqCL+LYUqW
OVVERD1SA/dDHdT66DUC5+Vm0e6YSZ/NH4jClHVa5dFF/PJ6Ci85sLcS2PQNI2Cf
smpWpnRozd6u2mwuSnZ2H3om8zB2aeko7+dL+gK5eGLfzeT8r+MDhb5t/qABKqq1
v0hA6khnaWsqDGR8NExaXH0f92pgY7baxZ6otoOONo6JIsibvWQ5Jshf223KTSsC
WCM1jRr4XwzsTsa1OHhF4jF1MBczst7L6DONFA1fWQ4S7y6QNba8uJQ/6bpYN4ik
ckOHdWA39LsMQlwLdc0vtajzkyeqfb9SpM5gqQfchR5TRhkcEQBCy+twOgyU06jw
huE1UjcafRC2S8ZFj5hbq3Dy1Thac77ZBkqqdb/ljPMsFNLkAwOyCavS8GIz9GRc
i0Iuk5XOrxlPAOHpeO6qyEKjNfLlFD+qUD3LvNzDh7lxcSx59hKCf2VXfjHj/AxR
6Ug8XvhKgg54i45HJMJN6nYLxF4n9jd3raB2iLNr8qRS5yDS9cV/awZdeq2l+0VC
aFMz8M2yz3FpXwYSwtKbvAtH6cz2D7rEJ5b2+s+O2g9c1ng8SlQX2nrwWpjwkdiE
iCkCPy2GdHz2YiBGivIcN9p5TPwi0WQoD3ukIVxSf0gWewEG3nev/YayxPdW6zEr
73/RFmRfzBjLRuLQPrnZDGalcw3OjgmxzzSEVZFu/My8e+HjC3iR/C3DrbIOo2gy
pNAD/2ch8JexjuLmRNWgqX25icmABRVfXT25GrxZA2ZZOf6mW6dwgppuV5w774Ir
QTS6/OoXjArEvYbSQCBpU9x+xHvOMlSGhdLCFV3HUZk39CG6qTy3aF+NHDkLQTyK
P0R/yGZRAgXUR0cIANuzNQJ57fLrjEDuP20qFJjGSFULDGhcYRH42fgpHexqJrBQ
i0h9gXjrXJamCPC94j9fF4jcrCusH/ykEQnjqhJvPLeRY8YwMuptgttb6uGWTyUr
UuUGjb1pIqIS8EoBYL79Yjz2C9qyoF+bD/EhVVHV2RQ63nye3U2YTiqkQiaNwoL3
nNhgnuLvNFDS2IVtkaKeLgwTIbQc8EhkO0gvTBQfNx4yFlSKwRGKyHSrt/ZAsix+
TR2/7nlCdK8n1RK7YJtktRjFH7kAW+0E6jdLRIOiTqQbm54XSJxaA3by2h/i4GSb
lP/Srd44roK/HJfNE/4TbAB1U51yplbiY46S3BLHJasO6/f611Q6eZ4oPfgfalG1
yQJa0Z34YCTC33IlzZhg2OCCs1ZLdQ53qk26DDX+i/fqi84vd+BOOZYI+nrg3Rht
rAicVGiqcPuZYiTedeL7eRmdX1fzlf0FrfagQIYgBPrJDcJ9zX+PLobtd09hMlJA
a15HqnddV2WzOYue9+QbxmwhrnA2g42nOJhf70y9Bx9VgzOMZAkc6zpMNgm6Ggue
EW2LRbCn9UdPIyropIWzfnaTyu+f1C9T7Q0IqH9Cgg3tByoSNrejAp+YC8Xd+lND
MB6I31FhtNegTtgCO4oqfGD3Qxhvds6hSHY2BU9Du2iPclIwQDoZAMq+3XxxhMJl
tg9JuWD06nrxB2sv3R9enuIohFrhFRuT4IxEgmqZCcdiHt3hlonxkL6Q8jp5jOHK
Cm5ZEvMwvvYfKMJT4ATbVNd+ny2LKjIU+OWnTmBMm3ZFIk9aBTYQ8WKzJeJjQATe
Ph6gm6Kg/oAwnM5jCnv5sZPMzLLzFLwIAGfmHboKn/HHDSnVq0QsqcmxkfJx03s8
k/t78pztSTnU2Hh2+qDtzYVS9gHF/qeKSI7zpf/qLFauNCs0S14WAuBHOCW6CKWl
nAImnoWVM8o6F8KllPjn8BoKlpACfhRySUfooMB0hb7tl03kkV98+PF5BFJGV0g3
1P3SDQIa1bJ18YnofJ8288XS1I2WGDlYDfqCF3RR4RZNiKnbbIWDjkcIG1Sd3RQg
hkYMnFEUoyJA1ktpD8JC7lZFkdLhyYqUJ8qVvr9RHZBsNAIAAkr/RJAdC9QZ9pNC
ok37whmSKsjVbZZdwltDM08YVlV6KVF+qdGiojCzS9Rychq+4fgzKJu5qm1rC2Na
FouZUDi53+rRnZC3SSd3dOHGLWrsM+DVvBh5DvFIW7AnmrldN9pi6ykj8bu9qkNf
XezjbTb5iRkUA5eRZLnny2ixgfGVoKBEW4g0+uBY2n28JvdPsuOuFJyB9lavz0EY
+OkpkhG4UKP4uK7QTnZ5S0hIWzjuyIwy5ZTS2u55xzrFtoHRlAAdI7EW1AoavCmG
SdEcoJX4R+7eY9zNqHDIZOQx1eLR15/nZRlo59FIzvPbN1VvpXKSYknUmGsylbWu
qIf7wbDgyXHeUL1PPRh05gZiNgBICwDPYTNm4JHmICum3a0YaI7aj/zdn8wrFAXR
/W3XIuhUxTYe+b3uAlbV05Ym2qdvj4J7YdK8uhOv4DIo0R3zbmjllewI8LfUvNcf
k+ZhAWEYoRAVoro6ZUu1XYPVAuSRro/rw5a+XTsVIkhi1A0kzOfl8JiWOEyW0yHm
L0zThLYGt8ky7+n36WyxYffFME+JQnQW7xP//NQ1kkGRzK2Kneqnamp6ANsdNVgz
6KqpAeo87/tNy5iHNJCGagYtL+4QSz15P2bODvjbl/hdh5CkPdrC4NR4PFKHm1Kk
D15ByHJvIDyjgPqewFw4tDooOMyMRuLf9FyLo6dAutIIhkHh3u+n/Yb/yBinvNbi
v8ln8qZRMnXioEaI409aVjINBJYoiHAN3+i/EktWf/a6q/p8scPHo+1M0Cf27LBt
wCs1l96gSRZh5H1VxFRzLTDhKf42tK33oTvVzdwpL+5U9JYuijy7UZ+ZZLKwyL2H
jm4/9lOBLoJVeGolop8Q0A4uandTL9mwNo82VXvNzuqRWUMOVShygZY/axDDf9HJ
v4fYJlc/WYLDL+TppikGX0DNCNcJXbHbCcMG8T93WjoNUD+YYlkfxOFwIF7JG3He
SVbSqXWvqvrRosPILK4NjnbsGQHIf6cAHtUCgwQC9RZNS6gl8p90mdFldR8rz/BL
402qdqAaDFg3jIz41DpZVmhS6pwFimkPAYiucvXI+7e8+SHNjQsnp9TjblDTEG3i
oXe0h+YuwYKXRT3e2Q5AC9APQ+78kEWiFIQzTxn/oar0257AVYuq/I98cDsAJzdD
62rpLMIamxK9SIWgDyCV4sjLFjiPa5O6RsVMhghityjlD8ICHDfzcs5dJtXw8N8M
36oWuGz1r0Vxex/TfaGiss4Ro8mtritdQOTeM2Eu+z2KsU2UzbxDDX8IQHY5O3fp
shLK+7tYVQkKPNph82YOkeY1vt+NgZTNVuxyxjZ9Uk3PP0n6r63vAZjANtNhFLrS
iiNwxY7D5TYNqwMAcoth6iv5mg6oarKyZWyA5LFZAPD7ymWIY3+NdSqveKGW8MqM
oPjVKqNPCP0mcD16FvT6Atf90PAV+s/pbN0GiMhyclr9zuiTOQQbYtIMQymQBzda
HleRi1blHux/q7tEvESwi0cRTASdgrW51kE2jjTZGzDg+sBDpuTUfdK6Bd8I1QqH
z12JTjPpmTWdXfIEiHjaYJUOL1yF/jX8mrKlr1tJ9WBiqe8bhd9+0jb37uUe8pMO
ShIwyw28taQiGctpLCsdRvXl3+jOfrv5jDbhomrx6qyW4kCNzIgbyUjUXlCy91Sx
X3IbP5D4qM1RL8oS30BpOhVnrOXj0clRT+zPzWX+I1FNOXqOPFpOhpEzQ1dTD2Id
CI1mtZyKcjw5aWWXKCBDBe4ew00GLQF+mid+H/Hzmx/ylI8SHEVNEVXfCYTg351u
aR0kbUnlFM+cYMJXEDMOz2czpaNuI09DWwMQnTYBCWfMQd+RxuiuEsyzmmHyb/d9
hu6vfgTM75VNCaNNxvWNNIjWqddAkXT5m/lRQeUvWISdxAGsBEX9iT358gBSUEMf
58Z3prrwHCxZ2teBEX49SBRWB7YB/K1PzsJW7idAbtjq0bJb/dlQegvwUDP3YIit
gcO3vKcKz+FxMbXin+s6aYiPU/StyUxEnaSGuhr4b+6uCCBl3FY5lq5QfmuHAjXq
cvRThY8QNsf7wfNkokM8YnVGdu8AAbKkA1IEbHMbPhbMY+do1rjs1AhWjgo9wc+x
ggX1GEPU3LbHnwnGcLKRFhABt4MNziUfmW8czWLLyn8wCvoaU9pf5xb9atTYbvOY
ZH9oUE0Q4GSYZKtbb7Vms3h0njZ3SVAh9CRFMC8h5dEKY7C7SFz46h6/dkc9LCha
Pakqb1hD1rLHbAB3qU3pUizldM/A7+qAI9eCNM5JRMIfXTnMhjNNaqTuuPojkmuk
GUlEf/odZ+3vbcS0nxYaKJdkjXKVKEOTic7Q4FCUyU/TRyYlXDOInNr7s5JGoRhl
kQPpAMTnYaxYPMC9CtkAa8uyxYPVmiOn+geCnPqrzgG1g5JaLWeZ7geDGBfoF8Vx
x97wTjRJ/Cf2BpjjPekc87CG/OyP5mRFAtTqhozOMZtd8npV5TnUn8w9pUl8pXuz
FjUN6einmhtWtTvvoViyVRKbGmTlTTh90osOGmjSUFfy/yFYgqxCAryzS8zMZ2ak
E0Vn7qsV/GV4VBnW75oFfnBMiPKX2q2J0b+tUuYfxUb5vd76TipGWovNuJQSLeLq
ic1N7Hv6+0561XqtUZVbtBzUZEN1vfncJz90NacuAoJxd7d21rj0rnYJIqPvJ/3O
C5VtBHfvVo9zjniFV9oLwyhGLmmtIvw/84vFJwzD2G9loSj2nFITQIr28Jfl9wVK
xFc3K+CZBS7QEjXALjrUBhkiGnP6u0yLDqGyHUOircvRlKMeIF/jiIiU+Nl2a4rM
nizUBPhi310uFbClZH4g7j2bvl6FrjMsK1B+itc5TJ9P4rXsClIrq979+C18pDwK
Vjie3ZYWNx2cuhAvOUaxtkUEDkmg0TxPRwGq9S7USWguoj9DES5VjbtPyrt+UgOO
wY1oow767atfhuK1Sy9NbRlHIdrVUZ/cM4hmOvBaXenyzIe4n+GdGpRR2aheZXQ2
9KJVFqV7OXWJ5su8QIa6txkkqaAYopeBCIAY0aThvrQ2WBq3Tj1jaq744OmF6OQf
tp6wJ3Scv5f4NlzFz4NpPqXgaAuRASzR9UR9bjefXr7h6xKX6NO9O0GWMoSA9Aq6
B9FAE8BuViWFF2so3YkUtGsEecakebyV67fhA2u4J05sd8lYDsYiUZNRZQ9qEOVU
XnerBPSNhxn03vT29RM33nPyUECVg5ZhjXIo4MHHqLvnZd+7OHyxmiCrucrOr+LZ
Ib8zDTMAmH2ZCLOTIiCXgXwvaGWFW5p5YlmnyyllFEJAS9HEgBf0F91jwO5SMOtb
D/YanXVi8q6y0PuMRNizEY19ClEHuR9UxV5D1Fhxmez7m6MzqXYhKwgi5JGOjZtS
qBl2hrmAMcZryzydqlMbsW9lSBSlcyz2FqNNT9fAiRWFd2uR+RmdlGAWgJwj5Unn
buezRFsL21zOwCu+8fgWf+V5NizbSvNMpCNAaGB07of6T+nIPjjHV9IdnPRP3Hey
lT8wjLz3yeQadtS2292UgfI7ITEEkw5n73/WkOuL4fHrZKTy8NDnO3ShLlBQhVA/
jDjK5JfTNTUPZAJ7jSP3XNPad30feGXJ/lfW00N+4RSfSrf10DfrX1y+DlrN+RVG
7QuLpxCfcvJgOVfxM4zC5xnrn9xFBC+9yfg//a9Ns0E6LKzW3XQjHb+FF6Q3SOuV
u+4WBka1fDEE+h30xkDkINMgQAzLh35PsI3cO55asAlRPq9LeAaRePxDiMtQlbdl
LC+OSYhwhVM5p3lXxLf1k9eNZTW5gO0qiE83Ar2taxK7McxETpuDNG3xfhMBiyqo
2ptJIRE+G9Cny4FIVfrQFrOxhCwD/PZ/6dY4/soNvlIy4OVWIsdKIylz0JtkpfxN
OhP+r2mTQ11GMFVEdon5pVUb6pL1qQeqDsTVdw/vP+c6eKoqge0FSua78pFNvInW
D8KOUSvZf0ZKLGk9I6/lN2Vz2gDA3+5EoaIYH8sFtvMor5vahNq8yuuE62xyjnF1
9Fk4TUKEy4ebcYROJGtxMWpRtZmmwshqtGvd/CV1VcxF1v60RoB/UZV98m51RhXM
jqQt+DHk1OMmA5LYvs1M0zvp+t++scGx5FpWjrHSwKZ803O59AM1RaoC9PxuAEf7
MkdaEboON+ndhJipV/TWMSqrzbfDyfU3L+ljufkPb261JWJiUtGxPWUbBcsUgGyq
V6PtprIULg8EWmt0nb4fkLecsoXgyWJeJq1Ancf/i3cWUuYKjUYPQgPbFoRW9vPi
AGPt7jPPAj7g4KHu0Xeq0PyHlKUI0bEaC6i/EaGrghKMHFpHHL0v1OLAlFSQ8FC8
6KsZKUrIKayGE0R9UlBdLm9Yee3rEeT9Fr/JBF3qZY4GAO9Mt79XqoGtHxU3RE3a
t3NdlTD4McyHQa0j7xQRHchpztYTwpQrofslfSYeM1xfZF6wgtrPZAjonDnzEqJj
cU+as6oQiAmQfyjCfj3Kjc6RU9He3vxyWlXrf9UFTPqwJvtaGWwj3RlrlqNRODjU
QZ5Sipln+aQbQ+yn1sSTVJhvUbz9OZxMSI/f0y9t5GqzCRiTNzKeZSxVmFXoNvou
8l7oX4/7U07wTgExOMxLS9qRPfDaETowdlnYRKVETAwF7nycB4H6OfG5ZwmHbibJ
hxEZkUT1fAz3X/AZjO341d1NgguyjKF5g53ttklQlOb/bRHDV/gPVUH0qTBIPGIv
vpL5umUzx5sTWGtHjZk1GUiF4VHIPzbwwVGHExj5gvDFHoT42l6xhdHu2Dqcdaw+
/vxmitccyPIToVrpRJWV86aWEr4BN1w2suLQ/xWw7fHKs3/+7Ej5rwIP5hH62yBQ
azxF5S9f/p0Z2vuRIrI5Sfid+EscSCrk3uLFxAQ/gQQslQhTuhOLnimUEo/wj8by
KCkUo9qTkoC+54XeqDjpd6kB4owyaI8RPSg7IYZzMbnPGlRyaxWGYYbun8WYGvhI
DibwGFdPFJV4DVDEJYE3WmL1JIVIMzRrO5FAOuEFxCERGKl08PtItjAlfA+Z06G4
JPHpz9AsSBjFh/kfJH4Zr12jS0R7f5oFPAzIQLOp+7DBt1rSr86kmCdHj8tOo2dF
sxDlWAXaRPaEV5hIbVlHX/giAq+BVPYQtwaYmB0zVtsirFO0nXnSL/zawTf9D6tQ
nR158uvoDT3QKwVjnET6nuSYb7BICyqOIPt/E6sWWnl+kWn/OxaC6c1nXBuMzqcz
ZPUe7qfw6TZGRT2h2l+0fs2u5+QdK4Bwr9dGmFm2zMa6EOKb1d7lP/FgkYcYPl9j
rvY9aeKihferLov6x/Qnd1qhdVuC1YFZczQndkA7XJ8gu6ZB2NU6kFRnmrITsDRt
EzaeQ6SXCmyQ3bupJliXQHtH1gKOCJ/MpYxfkhP6Ph2sftIBeG6/kYHGCRJ13d71
KZ+u2edh52Kn9oBrQqw7Z40j9KVYBN54h7NhdVdxgHw6ybyt1yuFqTrV7oS9hZZ1
+fYJEnN8ZvopDjTWVzkXqoiTDJAl6pxCuTth96oR4GCH/qUtlYbrbWwnMa/1Fbaj
jgnqKX8kyaKQtETPEMqyWRl3RXQTU9fsAsRTGbwZ6kdUOaPi0VAj3nn6JvvXvDdQ
KWb51QA51Fdned7DgTeSROHBsEyoxlmgkUNnvKx+f2ols8NgUS2dJRW0Ls38/ADt
2H3wSjieVYj6JW5Nli6F1zZ0ujABUb0JXTdlf5w9i79rR/AQH0ZYYHtC/8SFCIJA
QIpW+oVXt3tpF2LXnlWoeVTrJQYChWhSVh+kblaf8WrS5dLgAtjRB+imahKlpzBU
n2QtlQRMhtEMJmpenrsg5Wiri2RUXOlnKbx5O0ZAetXf5hLqyMHOqhY2tkXH+WQi
T2743M5UfK9BYiFJulK1cz16o62i/IKY1rAtvXWqJoH+1vqzYt0FNIANHmgZVlLn
dSXPbhIyKNIC1Eapyl4lxzQ80FeIMFU5WC42J+wgIT3prMbxqSC0gQYdFVcCOKVx
f2BVYuxiglY67XYT1zkJ7qxZKYh5IU4CHL6N8Q0LrS+iDinZ9A/CGsZ/GMUW1Or+
1vP/YQGxP+WZQt4cE5/zkMDEB1aaXqQ8gaEOxqt4Ur7p6gmKbYylluwKlcHUzXWw
bAhii5PKMbvLKNyOzSe2lYakplB22N+5G9AOdhfVGSQFPvY1ibo+YRvSJJhnETdz
vrO2TIhcfpEV4jaG2w+UvBEwOOz+Amv7l1QgSHeuN1SexbNn3wICZx93N/anwphi
mw006iIN15S4CzRerCXB3WiuJe5hwcArcDOHjrRVuO53LB/3wAyMQGre58tj8GIO
ylN2W4yh7ehOIW5MAntihkN0E0vewh5+n4n91FvvXTJOPRYuKeilc92m/k7IdIaV
1nOaLl0zjHpXtefwdhFO0jWhOOCYOHZ6Wc5ag3h76i6iCEvcsx7T136APJ1qS2Pu
x1vvCZ2SB+LxJ12tJphzZtOY/+lrHm2J1ll+As+dNVgRA82RL6FU/oSaeH6/VU3F
R9Vyit+WTt7OwVQOdVnhs5drxB9uMgLGcWqWSXswI9uP4sqWxsmdsW6f2o8JJ1xH
3HV7sOmcpypIRPRj9ubXppUpCl5HuZVoUeSgLcMNIDpw66skz+BMKeq6xOyu45a8
UaaocAQBF9PuKNRMBbj90zBJHLtMce5WPh+wA+7GH4YU/kgy4ah6mFP5CQpnBl/U
SMp2rbVgKQ2lSOk5iR9X/Px9j+t3ei2LGcth11hhi5QNwb8ji80jwGOy7s7HypJh
XL23yFU3YCqad1DgBhzYAXv8UgSTlGzzJW6uTXHLuSh9rI+joOdTUq8P7xWhGuF0
er9ZTYw1lDrMgfvwff4HPy30SKj4RHjTM9rtxC3phD6T8l8UJF+zXdnjFmrkL+zM
USwrW2tdVwggBe+ol997pSDypo/OGhoZuYc5BOIiaCDmcly4aZmUUG1bx8Rcu9Y+
RP1axWSSzhwvcIb6fVY+dJ3hxXmH80XNiPd+HDIAl88lBVfc7++pwfW8kvABmmPk
CyolBCFRWpbEebdPiI8Jb2fSUPdUdCebdM0Y5fg/EcMzbeAs26Hjh0HTeYTic/vY
h36XE3ruYnQrKRwBSSOv3WLkdwf1yfZRuznwIc16bf3OBxIMEJwHXacDpJD23wap
mkTrFIlVJORunkdOzj0mf1wYkVY+yiFpnhH5QJw9QHlU4Wx0R6SmSj8t3g+e7+dk
tHMhcko2l+VH/JIEmEPxDYb4QKAUG98pELRHGKeG4e7NYKe1Q+pIgYTRHsM0q46s
0K+lXT8qDGGMhq8Wudi4S7Gr9P84SBN1AZiT0w5koh8oQt8NauMr6GYhYt8Xpbf1
Lzq+D22KaoMg4RfEASoH405DzLF7wo/SN33gzo6u6+EbuQhRtmbxyxaNALFvObL+
pj3OA9AlpBIV8RfWjQP5MiTba2ZCHibr0e38cKAtfcJjYyBwD2R0j2jBssEgwspR
JG2Fy2Ex0uTDy/hDSFh89lrXD0bZszAbbwPQc2o+jefLTgRoMnKR0V5AdCgEA+5Q
ZOe1WTVUoN8HP12RCT4Uc6hPkTKTVP6ATKh80QqslViyGL5C/nmO0ux73etJSGPl
E30ZNSvXpz8abrVX1nAyKo5sSi8zy9Kof0HG2hf4AWMmULZXTYzENb6OeKFvRHiK
pWdci+Zc8vXsjeXO2E3ipbXnSYTlZWhUa1JZAFFg4YE4zfob0hMZkmY4JofU5bai
AvFWtuXSiRxOHqiMHy+DWJilHHO1YQfUeISThIxV97TIimv7XrhUpzKKPQyYRUWZ
z3VTOzY/e+pobkkME/vAURQYXk6d19f+w9jGW/GS4zY=
`protect END_PROTECTED
