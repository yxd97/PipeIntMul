`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ovekUe7+HHRenOrPummJSzesErUKAssCX5Ql7uIB5ffOJkcpw1FHioWqzzHc90TI
+zEE9q5aGnWELQa6X4yBjh1CoDIP13ExnM3jU80nIa3/5WIVzbsudM3uI+x3tO0N
MywBjh8xWavOwRhscTgPmr+gCGyXU3wY1r4oox6mEBaTtfK6+K0BmKQeSVw0cx5h
H2ueDU+vXqomJ4gfMcC96BZDAUt0DDhNKusM5R983jbP0ygpOHf2M64x3ZMWVj8h
4D7x3T8mXq0htHiUhi87vjv2YNeCG+dl6HbrtIEMa5hHptf2pnAU6luAaIKYpWol
kV+GQMXBX6tOMDMX2IjaSnUDvIsR40KC0TgSrVijPKaA70vFPWUP3dLdIztIhBT/
c4zbWyebbfQ4BbFasKJdYYtrVHsTgkgAKjd1zE4k5tbB43xvw0Y79Ln0vJMcKolj
Ha/9O9sjStV8QYFfO6dR2CWn3EteFKOQ7yLc8Gyhgd485jEaAttbZ1iqqOe4adm5
WIOV+05sKtJZy6syxhV0hC3zUjrYVyWOp6o2eTCeTOY9SXKR+5N0j+q1kgUvltvh
e2tWFFO5ZjvsD0rMISUEpiEDSBRo8CEVG62gtJxvayRIDULMlLRuZ21aZhMf+4y7
gcAxy/pfUiCIzrvLbi1FiNRj9cLDkBdfjVeY0AZ5M1nQxD8NnDhPi5DoyYGIxKFe
fDC4EQ6c4MoxUE3FGEjYYgGzKkjzQluIsMlyos/YqNU=
`protect END_PROTECTED
