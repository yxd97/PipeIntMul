`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GI2XqoLtZ27xqIFnawJj8+crqdDWsBF+phjLdOUCAe7IQmlYFQoIjxE4v36tTyL
iF/sa7mdeW4E/Ql3g1ZVfX4B1G3cxFXQRvSTwfddiwGbaiKtUG9bB63t/6sHDwWw
30fIQzAsM+LPnQLaRQ6kSIH/QNBLjDRP/3inKHcAlArZojx3MOWF02gs5qFGUuXx
nIt94inxTdhYTz8GqZ4Eiccs5VtQA3nMdVzao9mL0ICiYoFaCNb3mY3AcXpZCPT/
44iuGccp2bSaxWoms9gMk8I7rM/WgCMu2y+6A/HcXF8d8zs9N3xbAhayqJSGnA2h
zxfYui4DkPcAISlOWtRceheq4l4YgswgAx9hZ6fjzimGu4SEX33j4gPesXroA8ub
`protect END_PROTECTED
