`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nS9JAcxsQlw/C75pi+IHnTFTF9xUHlIyPIIY2ni7I3QDxn7zk4wX8RhmYghWVJoD
oXYLX/kEeJ97cHwznnpQVGnd87NhhMYC7DJwwpfKWQw9QNgUOOuA8l3d0hmiSy5X
kygvMx2Vu8eEvkYx4VIwPTgUMkzLIZk56KiNKRtWtbXf9CuBXMF7+YvEfrISssXd
1g3YjAnB0EdW7Vlu5CYYTK3OKeeyZa3InwunnPbH6RjTSlmdyUE+aPTiP2FR46uy
LbOnC7f0jTkB70mIoX71qHpifvxJzA8WIPSEOl7JuK9KXlea7Adj4+Eb90FpQOzR
pXyfpdMCLcJ6Z7EGLoPmTBXFD6SSqcDIC9lXFCfSuiQlF8MCrUz184kPunDTlzCR
eh36w5v67r4L4v8r3M2luPfLTbC5/7YRC4R2lYXETCnWxiFP0gEd6OLFnoDY+JK/
WZQV2bV26KA4Ce0XugV0wIHSOm4y2qRczx3xqMgnfltBqoVlxIYyIuqyYJsAznoW
IYfVLA4d9XPoMHwW7tjTQZTwEroP2iYJcAGeYsP6GL4IXkNkY3v6fo2Lds32ERu9
g2G0Jo4xesu32H5SHtzJkeP7GRZzw9tPz2RTw+FS3VZ0zgCzw/3LrnJeMw5tkirf
uijGL2VwteFRmIY4PB7R7nqJzm7Ln61BX1maOv5WUxHDUaUCguSfTltQ5OcqarQQ
xTWgfTmEeA3X6FhNvOd1hnFjx8or7y6bXvsbyDs1tp7qZwHpj9XIeHlaQkRdCxeu
NRPu0cXCuSqTVgpwE0xXvmzGMB6eN0pcfqbAvagaq5GXfXdOYyY9vOHSpqZ2h7On
ynCy9P0c3CGhM9w4NLAKwv1lrYRz6Q+bi+/jnqSoNq6hMTRYehk1d9HDgar3gfUh
Dp2pe+ZM3BtFLantVgUopE1JV4lZnFkX4yBIMtEUYsNwOOqZq+0D0QVZBgAe4O3A
rp+2EhrQFCxu03LNlLEO7xsZbVRPulU6uvkzPFxt2G00OW03ZChelgnoJ4skp7OA
bpIxzsz2oFGpxZAYHyaOG7Y7MR4NmoMDTj5dIdVwDbS12DYoO52ctTGc0wuKoF2K
HJvLZqL6RkNjRWZxf8Tp2F2oBLWMqQ8IVw90fIj42GC+51rscyp28WR69ZG5eea0
N3HUpUdHgFkUJ2C3c74Ull+KGDbqmIDbTm7SknWhmJz1PN6V01/JfU04oXFTXAkL
N+0HMEuHwjj9BWs4Uch8TADh+O+ytTD9PhKHs1ag+9t8Y0COfCW9u4JFeavgWAm+
zS1CiLfCsi68n/Ch6lwWyesC/kWlH9Y1cXeS6rWZMHKr6kyLjeWriZBkjNmzSwc2
k2NVCJLy5YFxmfIH2mZeN3PUjZYCcQXJrp1IpfEeed7x0YY8B6UOxTSFEZnXuEmP
Y/je+6UPyGtXFogMYbya+TJm0PIBdJ2ph7RX7twNCGSKzsSO2oUAkqSDfNSr3Dvn
RvnGLnqWlDlJ1ojFRBAXjKFVKi1D9xkWCBtx3OCO81hpX7MajOPZLTcHnF3NH56R
JhgilUXP47K39hF25k/43yXzQR79cjucIo8jKkfCQyvDyZ2AvXOo35Lxu6/FqI/C
4UObxfMC6HZ1R1z1jQesNXzf6z0dh36W6B8h9sp9ctTWHesvVCFJkWuDPoPDnlDs
TIUcTPHFFFFUnhsSK23xRLKLkXZno9UhNpl8AEF66+uCWsrW2/joLWb+SATeDlA6
xojWRHwZD87tsWIJTJ4nCJwtsU1qfMDVW1qaBb8oWEnqpQ2FrkrKJCAwC64RC4gH
FiXALEh8LGNscnizjfchzGmnVEXRTumZNnuG56IMFoHVqiEkCxHoSX0MvAVLLRsl
Lns//eOL9LaN7uhTx6UEft4rcwonN4sD65jZD1GiBcX0bXqfpIWUSb3TC50rDUii
agQdExOW/kDTnjg4WWPX6EpI1hYISpP50Eqi9Rt4M/NjIepBrt+h4dZXw5bxa/fN
TVjOwlIBYUe02t2FuO0k3t2OIYy7UIzSoDVUQcgQu1y50NT/CEzkA7LrXvubbspv
nh+nv+gYpqchotuxPFIeLjFFUY/l5klmcbkxYznVwNtm4lo2lsvfIhf8CnLublwQ
K6rEoNHok/smXFxJZHzV3mHA901HU2UKUGHDGcLztQDqF/Iemca2mdCcKlI1ItlH
MmYO+jrq9eeMFhOzDDldyAytQAoldj1MLp10e5WdrsD042lGeaNY/bgnjUCDDuGG
wcHLP60PHw+iIoZB83o2owOxVbdGSuxXPT0Ly2NQI97BT47I2GXz/aiEpKyBAwBq
PAplKlk9G8UwOS93s0Aj7pInzXiOXZ6qPW5EhhnLdCl38OTkM0+mA0fUj7tRVrcU
T/5aeEN2u2KKHdbMfsDO1w9vM6pBoovzNQyTS29QD7kwouKQhIZR8qVn8eNtgOzA
aUD6t6dL6FacdPGRxu/cm1Om9vtY+l2ON15SCBEEWUdTTAtP6brYzxvmERJTk0O9
VXPFjXYbTFoPEZggH+bFHWMiGf0VtXBFImGYOjzp2gX9v6BM5o95UNmojOR+Z9+3
TeM5uOvdabf2KZ0oXcpmzpWQCMeyqSyyudJxTnO2SBcXFRg0tkpEfFW7Wylg6UVJ
WTNAHSpwKMKHyemXNDTn4kWmvty1DzLWZE0OTweGY+zMbzutNlvFm82oweZDEO/W
ph1eSE7Ril8O1mUgRHtZ+UczF4J7Cg6aqQWhJOTFNcCSkOpQQs3ZkH3lNe/n723F
8lMr6jOaoFlB3/GVaQVq5f/UZseoFxKQoiJtUwEiSgegMHg4OyOK1OWM7ykxO2gy
yGkPL+X+ITFCFcLvPd90/WkHVX1yYF6kHr+b8vn/TMV+zQqdn70M/4Ftxm84spVI
qODeE5hdp86IPYjwF+B3kIjX6Gkl7HDgnTkdeSJi3vxOzGpxPwzD2HpM65vzsbC5
j4/gc2zVFTBd8+k3pBC5UmG/J0xOQRU6nbMv3o9j3iW52qIXVF3hAd3CvnppKH+u
SGEcXY5ym3CFxriV2KV/IuguoIysxlzewrVAgYBjcPVo7zVMCKSE7vp1HOh1l2WO
qznzcerOgKGwILwWrr+ZC53OkVkyf9edz0D128l5yqc9Udf1wGE7oIwN/VY7Il+0
rvaanW3rcpQO5nwhdreEQbpQOs+iAZOagHhgqU9nJQ/yr6HjwTCyg+n7nz3Gs5GX
31+j62/cDpo2d8/hnaOoX/72ouOSTyc1Q30nz7svNHCZSDA0/WH0nAnN/r1ySdH4
pqjm9iPH+o7vwjg1ovxnQxPm3TfdYAGlMy/RskjG/IDxPzScL54nhPwkJUuiE8JB
CHp5vCd8Thu9Gx3crwjOCx29iheb2mJwIv6pLPo1RboRjAaHVdFJH4Na8rejdLhv
cNrV56E7t8vBfEN/h2/TPFXhOzfLIHTgvXzvg3OJiXrIRif0fhga37bhO4nTdJxM
Db1Xhey866Km2rS0cdJCyrx+kUN3hnK4NQ2ScROtCVgV56So6W0IyoP+77Cx5/SW
Fu+Wo6Rec1l0bg/nsvCzmArXjR8ZuNpZiqYGW/TJAdcqEYL2SQyWRmyKnefg7A+8
/rudnsjR0Ow5NpoePpUKlZqXGwv7pPi5t9/kiom9/feeujMv6iSxNPMUK9W3vudm
2Wn6ucflBoa7ZAZOOJ2gCD0sbry8YTNJY/Nuk1qxLgJNiyHhrBoZdbtOJTnoZ8GT
dQyT2B63kS1BCJOpW3bOBQo0Vjm9eJ7UQpBtjYrnpuC7FANWmEmgJ6RDxmMR9Pj1
iRCkvUy1C8ASpuT2FwsjO2OzqOlLwIxmC9PTyG3kStzE60L8kRatwWXASBI4sRnA
7RLSOsIFLuo4qQcIi33HNcsHN7IvAxB/TNM5A4DloEjDaIqZbOXCHCjdfFdgOfGL
Um3od+azK3TskdP82SHK3pRJuF2wUnNGEONB2+SxCpq7I3O23V/LsoL6nnL3NJ46
la2ZTErRTnR58Cy9m7NTP7VKSgNUR+aU/Wmau4jP01eIN4nz4aoWWbeEgWkvJ16W
mVqz+STGKoiiRt+DC372fvTSGrL7iVKb4hnxeCoxnTisOkjMtI4G2VC1zPFl0t6S
VJBoj95/hyety68bhA+AcMrg1VTh9kgZ8wvxnpyWwrAtJm5kfRrpmcepGYfK3AgU
scct6wmUccv6dX0F9r5AFuNYB2pGW0EOL+llCg0R21CYU3oBxl1fWRF8IKzcz/Ob
ELNMDtACR3EZjIkJcqhQEWSl4ooK7B8Um21uZ08Bq2HXBv6ymY9hDva6gFbyGJb1
uUtKIWZtTZoeG9MkH8bgHtpQMzYadiYiN/qbfm7ShlAA80JNuFgUYPMASXumsLz4
v36/w3oGSDuP9yXkLapjrkIzNQZthLL4ZOo5pjgwUdynG4srGKFrDKHIZ9ytTdid
Kn6Wq7z9ifaTBInMlfZ8RaZffeg3bQeHawodr2Nl6HYWlAiSpWdyrVyU55Z7THzi
xwPC3QzlYx9krgUpvehQ8O3+wFwrsxZJSYJxeZHySw+Vo//lLThaO8tlXV46PVaT
vrpNofmMRmGoujPPF5+ZiAIi8qHdU8kihQmBvc0804djbWd4D3kwIFoMT10KiBAn
uQNepEk+JDuZq6+Lh5QOGXT9OTyLZ8kmvlewtXSVhShvSQsXJjznBvuAWsdZEFfv
BH/12SUIgMMhyDgH48hLIEF4OMlZV+cK3BMRo4UwmZZVv41yQ+l2tBMhujQP4xwJ
FL9euXdfpqtT4pTYnwtnah9Hs1/LGupJlQrZmOE1IWx1RYInFEiPqEBqO+Tkcqzx
ODrrTqh+RBrvtpYzbDSqdIt9Lxj8kZrhHCmE8Jn3+TfTdsJ32yWA+3KluJIJNxEo
OxuZk41QdnjS3A73iPfvwBzJaZ89pfbrQQWMKrCT7rZk2HNFpPpWIdcjibMEEWl9
DASQFMr0gAdX0CNAWsjKf4kZoUkHz9CJ+o0/rzBOTc1Ods5a9XBC3m3L2EZU3blR
Ntw4itkpPbI7FKDiIoH2CFhLPZUSRMNDt8zETQPh4bAr6j5tZQoIuGKj5pQheBFS
r/+02f8k91Xy2ZpO8N5dMEsuEOJvvIfSfhT5/QY7LyyXuwOBg9J/wpzWF/C4ewQD
KHgqgM/SAWpBcJ9xnaphaB0kiDOa+fETTodhEzz6+WfwYhnD4Vt69tqns6BYxJU1
UUXjItsOin4vtnpmVfxH5bcu2MiADKmcTtah17CuknDFoDNQ/HyyrDZB9/W4+Ogk
tLJv7GKFn1JSdp9KQCYAEKOt6p/3l8852Kc2eaQCVXJCzRmoMxcdjodO39fEHAt7
zH5ildNIOuN0CjG4WsCrEq+WWCfvvmhgyG0KmWSQH4+/k2QLwiTTX2FPMT/v0Ufl
KtJrtiD2BmMPnJszJBIYQ8jzKwZm8xBx0RE1WnCdtartOlepA1kMSLHhrr9V5f8n
SmQovrZ3wZpGMzS9KTPIuSlCQp8zEr9qeebeTKccxrMcXGFTqVJKpqjrKOqp3Yet
TFXWoweNL5jI3ZMNam+wgZg442gKmhBz4lbOY/XbQhawTopjxanhi8gyHLPN2k7x
pFUNuQeR3NfS+4eTsoThxcu1+Ugf8IFj7NFPba+IyML/lMtPdX9m49SM2HoCgWcz
0DRXQ1woQ9rcquiU5AuP+AMUI4fBS3UcF8UUZyEvKOoP3mgOiwGb3jAXIIn+ldyc
9/GRoWg+fMwRgwzS5W7/3HW5ENJ0W5QGqveh4+dckm/2IFnCjK6fYZw7UB/8ElLb
rkJeJ1/qHk4rHIXG11OFkZJR0pOmZlRz7FoHBkqQ5ZRDAnv0pDx5DytPVE48B90j
0NuFHUDJclxcFr3VSAehD4HiwAjbsD5rh1xHEbPb+7m6Rbd7GBmsMe6fv96ZsewW
7m7CvK6AlwdV+INV0831cJhcLxMHk0fqhBNzJSSW//6uWP6ecBg1u8D+P+/13inD
8yC9T28q7m+tI47M5jPMnSb2nt9UQPyuzg/xEVaH7WTzfjajA7oK/R1pC9hj5XSi
cgAV4k3tKGCaTbziaQD7XJFOhfOTSUCZXgAP8jASkUxS1wxkus0d9iZAX+tf8rFz
227pNKs0TB9608Ssjb3ewjGg8nBF05puLXp7MZXEkzTTaz2g4olPlE9qMyZ3eLDU
DEKigIo53RmDT2nEnWfVcIvQ2O13U5QHWbaTGCIZy2dWTKwHnASdlBoeIw9w87/E
7npEVvdbn7Una16v9mzylESqbSfnxyyGl0gZqbDItqt5yhSJduqs7lk63vqRuW2q
Ce7lYlm13lRNOoxPkaQz+4FphzTMThvq6yDObl+G4g0J5hesEazvB56+8/0ir1RB
R8TzAl1jYRq2OW4IEv22TsAVjt4Ebj1bNSLQPjuce53iakDOF5WcNDVtSXUJF8Kl
BjNsgySqS9WDP/BP4F2OMF4kRppprJS/SZAp3FTxWrkz8F/6X5mTmjfoWSUQGfXj
4pl0YrhuDg29Cyd5BFldJMKtaaQKGrhzhPcakp+NUageWwVzc7xiwmBgqJybcbQT
1jzxaylc9wvoDqV5RbX3w2ivRbgPl23er8ZPhesTk2JX6TPlobGMHcE6ZMB3zgsk
obabZaRC6EAZaF+9Z3wYt5wthpyHsktDxXtCXmtKY0iLNyGLXDwOqLedefLDuXhq
y/hoOOPnBnEI/u3LvKtjWsXMJpbbF/ZueMhT/PPZtXCB1z+lLWlcbbChJyanlTQm
5b0MuNppxb8TfFXUROnABx3F89NOOgRK92Ywx3gGfdwNQPsXgMkBbV8VqdgUGsFb
x5Z6EeuQySW/b+Q4klHHjShNr6nFjIOQYwZ2r0Skgt4vNEybOMUYkcb2M1cPCRAJ
r9Hf0SVvgH5sNDwuw8tM1PhcIhk0jx2FOKx7UtftjDsgeqHSuGTtULcMSZeY9u8f
IruGh337Kgkq803TFpQkuxPj8bZSR4cpXcJkchufP6oI6OnUEaO6oK/aBXNQ/H6s
fujJKcLfpeEThtzI+Ms8hSiFP2Plw2quNMSQOAKdlvw040dUbAqjDPlTnpDYm3F7
1OThr/pJ4zc15gG+Mtmc6BSbBrcreE2dzowOVaNqGXNW0VcfnTUGiE94Cx+sIAZz
ycRE8Jfl9blDhv4JoB/Bs3sF9KUZwyHiWWYAYQGLITPbkoVTmJzid5d/CiSyKsIO
Mvv+J0VV15oa7jZY5habVWAKA5Jvp71isWytPnsokOeNIrDmshkYbtjHNrrL/d87
kh3qqhGJSWgwT47u4IRwgNV4SKCiw/g4oC/1tlWRLDU8jCVr71bf1hAFuqivCorY
RoMJGxSvGlGevePe8fTzm0mhse7iobj4mrXg9OkTQWmfgp8pY6+6AUk/PNLHluU6
Lyf6EudznYYnC/9/UzlSVAbMi46BclHETGgDYG+/eOrTsG5d6Rf6f79H0RLl14Vp
t3pTJBfM7xqcbfhjyS29FawCmB2tbNZRZxCGoAQ9RWccIY0lP66VYTxw/jwmIf18
d6bhd3dhBMkuVvnG5quPQ0vRZ2+CglFEXRgPAf2zB5pnz19no37FEf/7PVMy3uf1
kU7ys8YPzvJh/jfatB21xkp43Ng+IuEqR5tIVD6/cvVO2TiLzQ4+dSL/JfpzqmWv
Jg7jHGKo1N7UCRy6L0CWHJkIYN9DPHwvhsjdaAhoLysJetOxP7rE/A9CXGf5Pvnj
Q8uFdnBoA78HSteWwi7lzyApmAmM81YsCPZds6TN5IJAX+94NVGLBmQDYdoBTosM
o9EDvm2phKjhX8Q5YsGolkDWRKHGPjK/J4TQXgsac9TeEgfG7oi2nwcdFDf+DL0z
FA+/Ye99j/oJYOgcSozZl/M9WnE61iUE/EhMsHfBp7c/DCeV5zMfr1TXJ7/QGr/E
R5RG0PPLJrm3iks4tyFaTxuGz6R/ru4IoM1jvxbOr87QXZt40ZzrScEibtohanTM
68EHZEAbZGPZZBfp/HphzijkdUrhtMdt8L/selysOflOJT+lyuw6wNp7Q3YlFZvL
pJXg7RxxMZ6BxXZ4Y27bxqH0aMVIXg0ZrlAkolmkF10wZLgHojmeIFwF+xeBxXjn
hA8nIY6dHKJpUlDSBIF1SDIza1fZNH53ddWLMPkv9E1nmbiJbNnaRTqq77G8zaIj
Rjf/K3j2aNWYHypNiT4SIzgwY4olhUHelJPnza9/W5ny5o5KIXOdGgxXN6TNwXRG
2HdyNN3rg/bKc4P1JchHR3q5N51KSkwSAqXUYWTET4cC7KkQKKUKTEWqbk0yeqNI
oVmyhPSEBUBXOj42cBmwqX/VIHOjNOZt6V/6cDfMugoDvH0TR7HuU/JJxVlovAve
MfkBzpE0p2y4J6svgLovb1WDnromt6tnNy+EX5N6GKwE2qFzx3axAsNGcfbBtmL9
jz+YPU+Z76bPbQBphUK8PFBDEuHbCFA2slqIcAFvWob8OudWLB0GHoCNSLqW8yKY
cV5rLzUzT9Cj/uWnRT/5fKYriIo606pS2t5PlwMnZlffQM9tPhgVd/dnAUu9nliV
jx/2YzdUlbN6zim6CzDS14fyCRpcO1vLFtRjex7e4kY/vySJOBcuRKjgSQagqB9z
DflE5y9kz3M9aNc4+C27ukW2b5AshlpmvyXqMPs2elakjEx22ssjRJQSkN0L3HxW
lTSS5d8bRlczb3haRpuUNXwaMPgJkcTFYrPXVPib5HB6eeChczWdVCsH1ayq7pyw
JfHYvoub/bUeuUoL2akZMQO0/swZ871qZz+x8p8VRE/ZqLVkpO6jK1p9zz0fDBK8
QtCxD0CJ+EmBVAdLzK/9EEHtA1zQX58ffxjH6qBFuodMv7nwb/Ty1IHn+484xhe5
5+q8+dAAYDZcAEC7RXXWt9YCf29WboDd0eY/ZWWFmkAf0hAkBTJMqOgLHOzK00bp
oqjC54B7AHrR4e6VFQialbVWMjKrEsl7URt7jS022fdFspOLOMZCrqCTL04FusWY
UYbXcd4fHcB4km6Qecvf2Z7MX3mvxNNYxNW58VhtRWxE02dkZSi3Sj87NjUdxsfp
pTyQhkKrLlWlXtaq4QnWzkMcSn49STSr0yvSo7VK0TS/5sbAiu+pFUD/B82fheKp
KQF/SAn0CqU2MyE9Ej+g9zLjTSMpr/sObHeAEKhI+Tu3EkwpdLlmpkGStOClrgIW
kMdauXqds3cPw9JBX6CB1VeYKPpi+y0LZoHS1YS7yCTkOTuysPlJL5yvWAFUuPCW
qKPKLtJTo1Dx/dUjMt6CK1RiW8LJYsGLSNzcCx7wkctGhR6V55KG4TvHGm98DgnB
deBD49BWYo5s+JXL/RYjJy8RRvKmlXn2YHP5UbZje6bsH2ZfM6RJoDDooj9i794q
apgGWRBOw09DbI9oCo7LElBTF3FbPhmQzbsqG95rxVfTbbiauuFc16RvVJhtl17M
eTjxOz8O2dbI893VHanTz5BRb3NQhUe2AkdQWgSapliPzqv6i6Y3ViEPqlUYjOfs
o0ZHaFZAYGjEPLXezCzh6llHouLzZKnwR5SuA1kEw2vZOIQerBy3ZNUcLSWvEy6P
niDFMoP2HrqsryrnUleMhlfirp96tSBmXoPXS6G9+qa2hafJnkh+ERjoytbNfzIO
oYlqKdljJA36Cr4ICwLer2ng5YOtU3UJzQb4g2t7xMf5EEK6VPqCEIEaIFGXzjYq
pfe7gUEgehuB4KXtazlAb44IUlrKmG6EY8VW7fwx+0OaNIDb0hYsmxwYrjuE3J6b
ju6+ZXqLxNIsGGVS0m+hVsOb7w0ye78qzZglwqXYDfkjkfi2RxzPvP5jGo4ztlFN
MQM596rISpH7GM0FB7hJs8FWU9WZ5Kq9s41lu+4ebENqaaR1vT5wJMs4SOmapFhn
HM0SbVNnXDCF7Cju23vlcJITHqFSKbgNI62DizHWVOaNAVHId/AIYlRpKaO0TJeC
4JQlAarYX8B0h0yJO1+0PpBNzR0BcM9RPtQR+1nF6Z+XAGjpNkJsAas7sN8aLNXg
ADHlbwQmgdnYM1pRs9Fxjw4q/PXIMfRSytevWEOEQofNyOKD8bhYgKJVvp4Znpk+
1SYPIFqj1/Hrm2PyixKXhpgbs+GABi5MiPbTiI21Hbk9okjx6SKdlcmKZ2MqyU5z
D+tnxKBmP9Pex5LoHkGl/jPXqbytvfyJL/nnlcR/yL3o8gnYLBHfdCPPG2dVeMe1
xzy4Ylu8xcnI0FUbV5H+y2AclAhoFqkAvPGJm9T79erDzZwUv5RlS+2SsYh0wD9P
Tdo1eLQLQmY67KKl0OwtlstyNjBjAkyoW1S5fvwUszNWCMFuS/1Z1zAm3ta50+H4
pOi3P9z660NdnIJ4LtRZoS6LnWUGsl7Kp2UFmsviqYecYSpwzlZyzT2KPmQUa7Tg
I72rktkwv9PBHlvNXuhsj51k8gCCEm/8sY2cRmitSBXBmjZhJR6jaBpdtdnjz2mF
MBB32RCnfX9RaY2e8tiAKsXHOBhXLJTD3cyLgNxP54FYda4sC5yvrwTzxtvxGxD9
1n8uPhVIbJv33LeVAt55gxP7vfbEZQykJNiw2skIsWOP1+gP2ZgPuAOV+1aMfMBw
xsuiU4gFGG829ubTGL+rsyJjIDIT11pgapkpxbCfH1jJZWyEBT5H7y2Atnx4lolM
Tv0wFhYlKukTdXCjF1F82D4y/XygQBZnZDa0ZyQE2ygUNZUMKzHI/8kO0YSvdpRk
kq+N0+d9glum34LHyslI1lymuAOxIJRai+7ETkjX9kr2cBpQPrDjnmrinSevB540
oLyG4glUScXez+bnwxwordbkV355UP92v/BinwBf99KE/QEnluAR7bHOOGMYAk6t
nH7PYMKN3XJNpWMJdh/aYhzCDhgNBypBgEvbbYBucqlyt9nLPDYiBG0HHWwbyC1D
smvIv/puMe5qZ+k6OsYjz5DkBLI0Jo6z526ppTd//GUJpk85lemoFxSXvn/7XT7a
g39P66WIYPeEy5m6H9i2D2eTTwYoPNWnFsB3a2VBbSaVFo/7bZxj9G2YLIcs/BQK
7Rw3votF1mXJckeIpNgCs5iH5DUUmjzoBXh9I4BIXsJUB1W2w0W+Hnpx9flrLXvb
g/yovEmTwH8Gkm0u21bWbM+FNq+UX4kHjMu1U4Lt24f6tShwsMEuBcMNBPol4sdT
pT0VIeq1Xqge2jPuRssTPe5zf8SIr+vGYQiY2zdx7aYcpsQV8rkUh0Yyh1hct85T
27EijrLf9HiMWap2v3M7ll3G2TQ0hs0JSvXEQb30lKq+A0xvuTostpWCUOSz+aUU
W7Baa2RBxxbUFjUGXY2QidnzF9w0YjnsjeaxgSWrjZPCkPWKs1Pjxui2yO/BIZOP
6zdvd9+H4pxCj6t+xfgAvaLiTSlpd3freMyilhJByHHcgfojV/o2+P0QX4IE8eAH
/iTzpos5pSxKg0DTOmQCgWEyPzh5BFY0eXmIeVvOEposFd8YuIrYwOhnGn8Y/HAD
qbZ0Zk7DGJ/ExW5vVqJw+Uql1JlpI5znzTDVx95NeC70NKCEiz2NLkSb9j0Q3YCj
4GXt8slH45uTCbmPSVBBhAnpEBbw6Q+fK8m6z0fVGvZQqV5xCM8oCo3UKVgG3bBU
Zy0BNLvJWNJ0COThqrodfosBzCrBGdUYxNQWM2SFQ0JYamAT82kgenfzEw+src0R
BQdd1fiGX37tBIoWmOzfbMmJSi8qthVD7nL8+MPLzUBPf0PcKoCPx88QT+/DVtzB
w6d3hXUjznPrkAA4RDmWxsdQWcTjxIJTn9UdEuaA0nCJsIYWYt0fXw8tUi8DDR37
pwFq2bIa5BTSJ2t+3/2FIekv4kYQsfn4ERvy7sgqFRcm3XMfYdkogfyGDDKi08Ez
OoR5D258pMQQ9LwMmjMoC8Jpb/YYxf7yCe/3LzNzLjLu4UydtHyAK+0/aKTiyfr+
QPUoP9KwxhwgJEskKpHqs7XdcZsdygmM/sDWViHicSdIz7IRIIQNRnLYCiZ0yjM7
PVB6zomb6dM9VwqRaAXfHhAfbRmj3O16gDvQ/BZR898jfF2S0B66uDF3r3i35PYi
8plExHhMJyivJSF+JH53OK79gdUcFqPA4ziSoms4TjNfxLLnMU9SSmLiTZdff2rq
Y/5AFzTFsjEU31qfTWs7QcOB00DiDnoVnx3xBkSiiwIm8Tbil/bHcym9do+mZIgf
3hlPQL4QVQ8zr2Vq/xyZfBIo+MdYZFYbHNLuKau4lk4tTlhLhwibPppFgMMDJ/ZU
PNIQlxzpcqF74X+sgLVQFgG5iRcDwtHDGtqm6Yg/ri7DNEJtu87NT1IjmifzZsYx
oN0TXsd/1dQPTwhIal7HDoE4hsZiar+/WOdtzSmbzhZLVj65395UoSIDwqEjTi7p
7pF6CrEKqs40Tv5/ewHusAI+U9TpND/SMXd1sIkiTYB72cjlzqYn88ly0hITFtD3
0t2i9WZAw98jDY5OBvJuTumqcICZpBNI4uxUpEz39YL1G3m7ph6X1KSbSMt5k/fn
SwHLNVGQY9+z3qAxwlZjlzApDx5qnxDPX0BEr+HjppS4wOwnwj1By1IFz3WmXCbo
ulMouycNu4SM5WK2w9UF/BhkhM4msNNGTWyjjNMskEL79OeE3gHLFsr8s7GsSM1+
KnzdZ1MHNdIfBsZegzuQlaCkv0VYMsjtl7D7KuGIjgRZJqHQXAF6QYZGT8vl1ckr
w4moIwNOVS39+U7jPLev+GmyDB3ESbfHNz7ZxVLmJ7zf/BIz6mValCZfvXz4hW7s
3QvJQ345bK/Tyyh6WI8ZDX7v8gKZLGZL9EGWHkbE8knIwourlH8d/LP1mkwZve1O
Qarq/ql/TdJWo4+Gj4MyK5Ek1WZMuDGCDYwlyYWGsMxgmPxbeZjAjSeR5lFMIZW5
Y3w7+oVmtDEPoS9OA/Seuy31IxzkhakjRQuss4EI8vmdoOvj3jc2Pqnukzf0oriu
AgfIzLpzwvnLajSgg3y4cWoFVMhesHgWm2/Y1tVJZsp1RhIpCwibFiXIT6qG2cem
6oZm68+ofL8zB3FOoPEvJJ9ESdyqxEYALaPRnjfB6+iW8cKqTQWI2HKLKkj9S6lT
S2uu9dMI8hgbkhEQZTA3dUPg0ZAPvHKcqECJzHnENxV/Kok1L/139REUup6u+Nnd
f33DBum6MG56TdVzLq6Mp8vFLlAAthI54gBcF7KSA8TfNqeumkMHgRFdg01s4wom
WLujgGkUUtCIXYCh/SWE2kqAgfqZTkZBFr9zZ2+yRKJ1yZob4YQshDHGWzQV9dQZ
F+LQv/j0VftY4iPkns/6rtQajd7cfUYCBH6EYr02e2toAEG1DW4eGS/z0pb/42sw
pnVObRrrXfIUYJFnMn6csX+c8Q3hlZKBloGTbGLPrKbrGTyQkcON+PPxsp6vWt8W
InS8w0VkhARgyN16iucvSq189onxDvD6NNCu0oF8Xvzz4caKp/q7b0If1IB7qJ96
HIg12ACTg9KrQXc74HWu3wA2XFvMBdpHtTDiNdtvIcPHq/YNgvfbYZQwX8kLgQuN
wKUb9t/42NXxdJx7PSx7kBr0s7zwqhi9dfIZafj8w/1znTuH7puL6aiMWPejyg0w
1FjrqvGw5MMWnk7AQbDyp5wztYgjEkrdev3PAqjdkAOgSpLgM1wX+9NZPZ8cQu+v
4tYnXObFDFYvIzGG+vNHX458K0Te1WcM87E5FFNV+Bm9KGn5SulkmMDOYYLjvdUe
Uv9zv0LKcAOIT21vmov5x7tBz1qf85VNH/BLgcEvZ5aJ5SJZb2FliKCaEvV2W8Lg
AHR787+bXWn3GqhSEoFX8DoINYcoV+kLIqj1CD/28tZJITPTitoyKcB+CAk8y+Nh
ULD+QQ9O6QByK/MEW/bMIgBGdeAnPY/EvK1c2xJsl7mhYnEDzEwjjPoAWFS+aV/h
qb0xsqdrzvAsF2Tn8HKS7OUU2yW0wkVAVdOGpOZJE7yaMhEH9+qUVM6OJq4XYBA5
7bME7jbTx9Hsr+bzNChAP1Pupzv4f96Ka9r87AazPgrn9pD8J7VSAlYqnT+QUS5W
TiF4mSJPeFR5SLWExc1CU3ZVBrBSuotOUZiAdTia3JjGMBJDC67oyXUO7VQKbaNz
Owyt6FjAvMiewM/d4kRcGsI6d3LjGhnxBftFEpYbLdiT7OML+4mfm8joVSaWeoXE
eqf2FyXPMgmtGWT5SRFeyBxhr+FPU9TjgViU3TQkA090x5KVzFHWMBIWJBwrsu1o
JlzxJepJiOvcwq2RqfqD5keKM5ZKlC0Vb0Y4mfSWwssca5oWSq8saxmXAUOTBcNw
erwEImwxjQdX7fAX5BHYGcIA4MCEXQV6MoZsjPsi1JKu1RF6Q4Hhq++xyqE1TV6C
7til8e0piIyxslcgc2SxAE+tqlegt1FcNp2HCSF3vQ1amDc6HSB8LlANMySCWlph
4Y5cM1tckBMZYHiRvrLy72lEOADfQWbRDfKsJ7YZCq+RNKs1UHcmUOEfNCR1AZbq
AEGiMeJ2N27ay956u6kE375QmKni8Q57FJYv7EUsi/QhOqswA+glnilLBcz/24Dq
8D81N0yQFE59VE1UeQFYUe074WInSawlIRDIjuk+dhwnbMwqzbhWK0worQFw0Rmw
EyChNd5gn/lji3WOX0Jvvn+Ie/fMXS1D+fEoinWap+Ppv2QmGsOwzsZ/rmZpeYhP
HVddxFiXL0D31jzMxeNQ5BJWCs0yLB1SR2CpP29lDCFDvDxqicg3UIV1cBlipwGu
1py3wH3c8aBHQkHeDdCoq/mBlwrdp7o5LPar5ltvHQjlR5bfNwuMALU3/8sfktgx
ddmVndW22y4rQhV+2U0F6QfXmn5DGFQ9ZMTabPxJ4LLtt5pBzwbcu77d2eA+Vv2F
KQedpjpTrlU5n63wset1QQe2KUsZFTL2w9hosSabD62d+skzFh+1mne5WojIA0zr
3cFiCtj0n9Rc5Igza0nLCiH7RLUc533Jqmui24IcVl0dFcKdreBlOQwRxQZkXHpX
ZbRWgRp2JD6IW3m1eKyAbWGhaGWXVJOcuuR5psLRZ4gwszHFWrKYqr25vkN3z+QY
+g8zDFjTOy7dE4q+Ka8U6oneOHcTCBfoTKb9AgjL+XEuo8a6xcYhX2bUapz1T/yW
s+fE/lSCvyJm943j/YjCoPbbSTzDjwgM4p8p6bRcAAO5dqjhvVpfPGiGeZfAvAyc
kTYVukn/8SsWTaZdWs27MkIxvMJMmtYWhR5iahtpFPd8R8GnDVexo+Aw6+wEiEux
f+D8HgWcLfUeNf7nQddncOrX9JJeFqFkHp5uib7HSqJSI0Htu9ZZEnk3mfK611GY
lfWOypOM6rCcvCSiXX0a5vgzKIx6fJuBweSlgWwuAdsicDZf/ODCZbV2skeERDDh
b6a4ZwULWI5MlLoSf1+JbZQ85h9gE+8y2OC2cs8xa+Lld+uR40RNlzMe/ula6TeL
tX9zwhDxFFUe/ujg+Vi4EemKBtzNyWh/s533lbfq+H4UM/Flo0N+G6kldKM2MC3h
cVxvwAfdWN5G5KTwsbbiVwR4xGt+NUAV5UX/ETZur4o64c6OjSxaq0RjcznKVQA0
BTMkCxWfAo7u7ydddDFzQx/cGl8rZkAJti8NjsNRh1laWEoGOR6pHApnsg2g2RLH
7fWartOGw1R91t3r0G+NXOjjKukb/gkzrnBGazq0WQBa4gTUQt51JNnWrFvljHbi
/xt4QjsvuLmiWIKmdPh6SIYJiOOqFMYMgfs1DWQFM8ByVsCbhpojojKEl0pT+Dgc
wl/mwULbAMPsiMniUgsSAs6ri+nl2nRhGwHvqy255btWPfD4lGbia31+X7mMuAgy
46YXvrjcQNiFXsFoegrXmLn0LorsqT40NDoMjjCWDxd5b5A8n3gPtpCKaAac1YIz
VjVm8BO504wmovYwu3qratvogSZ2VbOP40aqhc1afINYwfu6zsLYZAVaRHAcuK3h
W5U8n7dzx+N1YNhoYy8Hs66XAFsFkZtrOv4kc/s5LOIYfFnnb1ZoK/BjUerOk13c
Ec4iXj/NARNahACqdmWsn5dq0Emvj1tRUMI50olkdE+KelRAX3+9FEOIGQcV1ox7
q+7y66W563fomIOdaSy5esN+3VXK2k6Zfj5vfVBvUDd1DIMNFgFsGsLbPmbkAsnm
z+VJ91MQG3tAPUyonL/F84aMPvzDzDHrvW8Qqmdv+cK/KCIDveT4otdMTQ97JY71
8mejbN0an04pudnL3NzUhRESnNmnCF7yB5ofIGjLwz7LdTWzK/xguIvRMVZSwbnS
lCDIlmqhawiyVlPdSopULjBTAAOXBXDxZaQz304uYIS+aXpdkdkvJg83R2bY+YTd
mL7DFOWmqq+fOOPMX7Y8TqW9TTUamfylXNAq5kwkJTOojAkjZTTM9RgmMkl+7Wjy
eQhUPJj3fDVjIVdMYuGhTvFbtO2+KcGUZ6rDDllDjK691Ph7+jr60fJ/uLsWHmyL
oWk2Lvutgi0MelJVlYINDyMonaV7e+TdV1ekW9kpDv/baIb415Ov5saaaffEH76u
RQ7+n6cqZT9jyyg5TlMXohn19rcWdWISkMUSi9GQxsl/oquSFT5LSJPu9j92ZMJI
hzmrHFKr/1wBsAUb4ivP+aih6UDSuE7AdObXh0Yx9ZhypyMpFmHUmTC6RfG4wx6y
taJkObEy4ujntwTDTtvFjF+aNTZW79myliKMs6CPxspWPa+RCzxMUsJKdkZcBdLF
tG+DMOpPKJZSYsApqscefspp7gTamPYhSWB5bvLAZgnOBBSmGcOQo7lXL4XU0O+s
2WFQsi10NBjH5p65ae9+Pkt9AccmY4qAalCAgM3ZrWohgdez+iXrxLEKk2mtNV4n
K5HM7VbdPysgF+jtwzBne7azA2gCXIpSJn/PXTEYvCBY8zQIt9x1BnTY+af5bkTY
QiBMgrHKdUv9afvD6Pz+lR9aj420AUnDZFuqF8P0Q62bDLDe7dtznc30gtLjh2yx
AzUrPYjpFX25R+iNk/VW+apXwghUR/ZfBaATIuDXdsWxRnnofd0S2tAtizgSs2wL
LyGNrBDduTdQphCy5J1iSzSRTqrSs3frVIDxwtNc9yyIa6yPmWms62XBts0Ddm28
eZoOspND83e/IxE5O0rqPsW/jAI2m0cfvhtXbShgUvCwbo7/0VzQMjhoNEg+ZdUw
8JsZjVz7dIJsyieivhm3IQb82xYA0EZAm/J9YmiPI2EiuNaH9rwfl0veSQGVgbjw
1bqGp6pK3oyhoXb7nTqlfuRF55WxFRtC9AVvR/XqYmczjLluhAx0ubU60Sww8odl
RLxKJ7ZXl9AbVLW/uDneoZqrXPojgItXgh0y7TzjmOFrjYLCfMnL5S3eQQ4/JncC
6REHm/oq0FtnIyld6Kdf3Gyjn+KfIUR7a5e5djglCTN71E12ptV3B75LXs/cMZCN
l8g37RK6DP7acqRywzwxJ1feQbHIlVOamGQ/H8R/27IdWPQhRjNxexUHmNxte+0b
a3eetHdME7sNMcMcjoSLwH45joh18Y/NzWHRvvGdttlAc+hDSjmAaicAKNLtE73r
3MEWv7xtLnNzvD0NViUeDuMblLmsFAnj4WbKe3KrReSGuDy67DO6XKAUFzKJY5mV
mJW129CdN92JyZivpChPELGJqQ0yMRxjHxHkn/G3Ke6u+W6/Bk962hD33BKhOIpB
2qv+lul2OESLOtL6gktC0mu7IA4K9I3Ecfshl4T/zSELBXhonBafMwju9fzIDLck
UBBGBF+tt9lSrUMojAh/qMAT3glHVXBkY/fS9Da/4zNf80I9zTMwo26fbL3w2CMI
jiJeiCMQwXPyjHlZHk/VIqmmOKxiqJeKB8hvAHCRRXN31g3L30Tsl6gx5rEFhluS
lwu7VmF2sTkHN0wp5TqXoNI/WjyCCTokgpMp6F7nskjnQ92ytZA8+IygaSYaWTpX
7KnV5tJvhSRP/WXmeNwrzRWTvPtpAQDuDJIue9LT2Lvr6wRMuFLKY5C6LG0n6/3R
NzYjZP9xfVEzVyimu6xyeJyk6JI0/ihjiF5MvW56ilt5Ia1dJWBK9XxmGe30EGua
Oe/5m3TVv/Q9V3RzCIVo3reK3PiOtcroCDQmKLes1WRQoNzVQHUoE2lr+a6lRS9V
xkYKj1In5zlp0Qiwh9cSShoxS9RgE59T4oD8dMd4gcE8/MVVDtLXZ1Qu76BIVjfh
oftoRvd1foGembkjiEpb3SSJbpQt1HnCaiVOkUPJM5deeGlCqCuUWHZo7SJhj9Go
QYPV82mDSG1RB1+pDxGovO0BCsmhEjVSUVzoThqhu4Pc8xndtHocD2TTe3B+499s
nByF/ELRdI9SceOO2eomhjRNA4ixKHEV/9cNAy4n1Bj1WC46h2rDM8KgfxklvsO+
9fpbw94q42amLc/QKvWCjSpRZVF9x2ERSFJF5+vvled4Mh7gHCTYwIfWxOLm/Kau
neeEhSjCui6XTRI67HsmdjXeWgtlwhmc9+T+lxCGHVy+NN6dyIgVXB2JDRVlonna
uhh3O5NFKwXg/CzadHRT2YFeBJ8TJb/MyY7E+hRR/cJMlt+948htZyPQkvuHKiwG
7McGtQiaoJOJeCROI8gwb+/ztvHpCrIYlu3r114pZsodPmEJPjxdHCyicofLMFej
rLJZQ8qsxq8YFLFAs4PJQjhh5yUuPItnGKX3TKKO2XsJhWh2KJ7HX+Tli7Appt3p
2y6IVKsjAiBIrt4qArjHarTWmGopx4mVC3lBw5hefl/L2Ue4rqxnILFROENpokzo
yDaSWmMian0D7ji8T1IUDIM6dYi6qP9scCiLrn23yJlq6lgdL+NykZEbAiYUe5Jj
ITff+Kz0dLSfVteEGxwuy/0ff+d60pr3hyGlpCCIaabNR2fROKTc0n6M3vXejHqB
3/X6FwO4Ggb5LFiUBI271BotCJJdrR2rkvDxTCXtEBc8ZGp/Y/vHNP/SEgFhNk6P
q1rBqDkC3fTY44lPOAynQoZEok1bBRM7dMrz9ZNlZuDUvV3qpAvKJopQwFuGemMD
/MYsgx3cGzMHzYcGZoIgU0+uFYP0ys/MO6Bl9bwVbZK8aoC8xlDLJkV/L5TnPShG
VJLKx0eX5RFn+iYT3diu825YSBg06l+XStUtxMO+i6CxpWmwPB+m89N2RFFs+wFI
28X7sWp01zLFximKqaWln54VKNxq765lsSowMABeP1jjEHHokYZndJDPR5PJ8hQ6
+UZ2HOjGdmnmKtZU/q7MtgRELtSPbrSCGyGOY//BxrtgL3aux/MEDW7Bftu/Yd58
ngEN2ges8EoUsGbqU3f3KXyT9Szt0bf7Csy1jnKqCdAXyMrdOsmNQnaEy5+HsqLs
pZjEx47sReBalyM5rlwjvoMJxSKfchLgRkdLj9RHWXUUBlwZR+6BI5FsXNfdK4lx
wz8ESE239jiUPftHzju/TQNUyrJMH/wZMdujdilcuI1r0drgNNKbSxj3akEXNEtC
ehy5h7+yp0bpt7jFg2a7ceAHdnTeruJCk2Tp5A5iyLkrb4TQ5a3H30JXP7xy+LXA
jPYHx+YynRzB+itR+4qtrUwZdzVbY/iPLcJ2hX2fBrAt3aarKD9EtXDp2Af519LW
2f8eTGb0rrEjtk1+2xtAsi+Vx9L/K/PraKp6f9C9cKteqd9GIiGOF8qj3ar9I4c3
zhjf7/IkZbN1/pQ2ECztEcswSDzURt0G0np2DRAdPqIkXePdqov2ZFuBO4O1WKUf
AhHuVoWC3aK8Q5Ur2FnTU1QgYnnts/1RbrTKtVHJHHZ3+zyXuKg9t5nnOaOnIaJV
YJc7P30ocn34QVC1870BeLfOJh3KbldXnmttTPXM9btDLLxTzRf6yqRKqe+hO2ot
fZGakeAXzsDrmCYiiTHGBZ18wpOhyOpaKDSIxyQ6ZYX+rb6LUHTq6GNp5KqGukQC
vCIaNVlRv7RxT5w9FaqbodtypgHlz6MA3r/A7//IPHPyR8f5v50uzu7v5rbOqIgR
h5mcJhHrn5D2Or6+4Cx2kw3v71gKTlgaxFjx66vvv/f11/vVykDItrZr+1QOQJ7j
LjwqwiGRe3dFhASh6ZaER1sGXEQpV4CrYYyDfUvYktS2oE5h0uINhS79fQOqoNiP
J7zgdm6ZenF4rlamD13JMrj49M+oBBq0tG+OEEWj+8TDhOhfsplO462Bn8uTPktq
OEtvKW6OtPCudrqQXuyg/tWZB3Q2IOOfHSvrwsb/dOHAQBlRBFC9t7LXBhKZDVjI
IqpESPl2cHmbKFRzHDY8RpPXlGlQio0McIpKGAdrFoFBUqYwcHDokxewzmuhQE10
gfrzoKTfgCfnlitbaLPeDRdXXylBm7QhFU5gUyMgW+v1bKbsKYVFBQUuQJ4viL9N
BqyIpY6NQHoi0Ezes2ooCeGZruR6n5X/YMxrlrBMaPtZ29XVexX+3yf/tHzvRvLm
ZnkjoM4zVuqVbkX9H+YMfKegbZntK2zZhIjggRDNSMiAJulz28vobs3IehmhUXs5
jt8IcREf3Ac0X6WCVrXkYTJ2edP8no6yncMvdGdVCr4wB4nl7mlpCkTY2ChaDH6L
ywAm+EUtOZqnVatkknmv7rQ/HqIooF6SJiJ8QpqBaOAt2HwPSnyKmuIzEwQaEe5W
ARY053kGD2wDC6sCbb4V1RpJXrexLCglJFbP1MfObkrqXVXzcS3I1Qcg2IEAwzoZ
vpJGfAUqKkeiBLiH0O7vNnUrK2R/ZK5u6G8j7BzZrr5XJvIB6fSpUc8ErVthpCtA
bTQQph334eioHpfcCTwfpVH89ThOg9MRC0CvvvwJ/p9cOKG4JlSdiupVFiIvgN0K
+qquN1LVyjjPiVDH2DcViWJr3gLveJyS6oCXPYA2JXf1l9a6BDLDFI3z2ko4kPVI
dZx+cX/sNcyDUlOtNT+TjGYTiludS00/nYXUmis8FSR90Gn2FolEPyk2CmJVrtrK
X+oVg2VzffBLDHgWxECrXqHmSQQrECYiDk4WCcHtMyzThw3Ktk3/mdo+4a+IJySi
EGJxMPM/8IvvO5uL6a0Eyl5wUXhjb5CHAp23lzIRWv+m6E2lurVmuLR9PRs7OUft
Ayc57DSRH21B9lv1o9S3su1+3ny3Gm/4DAn5GVnIHkOCveRCXlajkdw/jbplg9Z1
S0oIGD1KzJl8YXH5Pq+K99WJV6N/LiPP0slKLhy/sBUg6Xp27gI1pW2ZoV4CFpy1
MprhbPfyd5H4xbbOn5+zj4LCXa3QhFvqgdjXxS8fY2k/M8as3bkJqHlJKNg59amH
6pyn3q2xG1nGXygKfER9/0Zi1ts04z/rkr0LF9N68sr7ie8mgaWeERyi9YlQknEG
SfbhEu3jVOE3cetI2jaItscnwAoj70c5egpye4qPyZU+X2wm10U1RIqx6F99+cp2
Mj8AiPullS/aGW6bhj3M2IFNDbGE7a2M4nlNlkS61n5gD9+1FvZdsgPA8517TByX
XZbxb4VdJ7DnqR0iQJao1+ro4YS3SyDmLyzdiM3Yv+5aX8w2vLdMSGLPCR4US0Qn
3iQrd0IR0BvmPMYxq43RPJe8bCvN7wSfQLWg0kGDRw8MU1TdaGqw100wVSouq1Nl
1PLkQK0tJ3tEVNVCNHNBeQEanl95kRn/NrF9ymdg8H9jKDRYL6YBaOzPTGDCWas6
gD/9AUhlexmuATCpIbij1fXR600ovTJSR3i/gOZ2ODohPW6LMGshFEED10kY99OJ
+0IX94oAGgx2FIpkVh3qWz9QcNKH0U6kxgBfal161IAsJraPRLL7JlEliQx/xfVg
49oxT47yqaiIkp8YCV19UFuJmbxy5AJk2ChM9WdnlKijKOFdadakyiBFyU2qc83a
Im+yOXaR0f3mSLWzu7atZ2BvF/IG8JTtOfWEfGgdSkfq7R8q8TNzXmirf3bIYW3/
9LNdOwX15AsHYCoroop4gwfCNwnotGjBumZZnf4/Y64+VYlr8LoGH8sfHqAszB++
k/vCHTuS/eB25cPd0uzhl/OxxkvjFZWx//Ydm96pR/EQpfCVSdAz+MJCODxIK+A3
7UvM0fpjsg6E+9F2EpSiZwKwRByTfWiGEGwBlWI5kjB6AqPWViaX46K41VJ1EFn8
hElAn1qA3xyHPXREdD/lBt/zV3KEv/xUm4c0jA2nf/vxDHpMdYdXxLSAe/Hbr4YE
7KtTuxueX2XLWpFzooLeWFA5gz0XKKJAF2qcuvTO29Yn/H1udJCnfn0QU7U/S/17
LYKRtWpqhtEY4X109sZW10/Za70TSJXTZ2WC+2zPIi2NvMOLd92yn4F6+TZqchDI
+IsVFF77Uv4VQxO+bg9dW6ZiJE0smPpUJ/bHmFH1Qbgkfh6XbjTqaNOSIFT3Wvc2
1wM3exSq8ny+9VgeobmCxeR7X68ADH6qTCxAbiVvDCfaXNI+nX1WTwPeeHNtpIr0
gyafHN5RTi5Q6PBiiYPvc/X75JHuLinSh6H9NaZrvBsT+IvZN8sIa40jrUx3eML1
X5d+DzpzhyJLrqIIX4TxhryxpmLxEdUazbQzSefYr5JYe6UACrdUVH9IzqcI4JMn
bWWyAUsI534tgrAvo/QIhKMO16NN7wsYKfW9yt7GPWOC84qdFAfXPcFcEu/0wt5U
Sx+W5Kcx903iZ8LIJdJjzYFjqzjf67jIkCKDjAjCTsOZYmnODIi+GzkuDzTvaiar
LEfhe1ZT+RIotWscCoqSy5+n7tjzJ+ea7MpSzImn2v7NeDQ2S9lgbrrvLFB7fNgj
ma8R78vijOKOlofkG9IA1hfJLwhgCt6sDDuLSoECFkzKO+7jcXK4z1FEDC4nx0DD
NM0GI7/w6QWScQBOnFtsmG6aPqLFETlrheVRmUfg7oytvjiemOUv7OCuN1C3se6/
wI2Uhsr28dSOI4ef7IZl1lr3amFhojaEr1UuUuUS4NIv/w5KgPqSoJrSrCrUuJdn
SLCf9Jny2J6mnVgBGZiY12i1mSMKGskgYXOehT6bDzpTQcbfhvFdhXN9iEXlOKGk
LdugiZiNCZTCnsa6Oy/vwiIn1BgwOYRETYnGfbPgmsP2Akz4HYohtRZ18/NkCcOB
5bYz7+MJeZ0KEKBEassrkic2yVpTP58j1mSfSZWxETnLgnbEkyEbvdQFqxwAxZ0a
pmMa3D+nnzkZfhfXkCiwRgUeBWIdr+gjiWQUNVC5CywpOMJlAr34YIttDNGIhxNJ
e1rev1EKou8uBJ/XeWsSu+EboWmVkGlYBkItMgPEYDziU7bwcpqL44PxFf4DtVo0
2x/dTv6kTzZqszqdH68w/DYbVKGdXq1aHgCfG7FBPoEM4npVvecP0Z+3JKI5sIEn
huekKHC1LtarAcJl7KDm4SFUYWa3P7s2Rt8nEtlEwKOk8F9FflIGmPWAbx+YnIT7
LLvDJg9ANcDkgWYlyjhS0Uz00iFs7S40iUnubRjggEj3D4K5YX54Q0sXEaETvP5u
BYb25yKaja86EsBP8P2wpBdM+1rHmEnSSsEJfayJQtvFlLX0p9Xg3sKJhLjG2NGL
pNMLRfkq9tTXihoyKXzamGACfHm2Z178jnMk1RaChyAitURP3TTNYvk6FXE9WWwK
oAaD3Ki0naPwdfiCUDdIFOY+W/WQnGCK+Lcp8PVqYKO5PvH6szXF269Rqz4Z8EbV
2UEJUsGXk4CyLJTpuUGzj3FvSakifBlFn8Lr7FOQx4mRU7KuEoePeBSYvO8cf4bO
1EoBKbxvB7eoO3Ijs7+uRsGIgI6GPETpD3vbRa8uk1AOqHnVtv3OuiVKV1sS1Wi/
zFj22CapeWZQY2esapxPWVmN6XFegM4jNNTdft8w2FLkpqlrrAum5pCz77aIhr5t
gnpRT52u4GMwnHS2v3lQAqTd57O+C+ZV+htodHYD99mnaWslSy238kXospA4I+ul
xbXDfSGaItV6dZDEMjJzqhWDi1urQ5E5iIEeJP95JPdmhihw6rs5TgbN/iIxW+3P
X1snsl+4u0Vk7zAg4RAQcI6h+/G8VsyGCZs+IUysFyk1v3QwcmYDUiZx51K2zzhz
SiADsRT/f/ioMABI3pgRU45AUCA54Vz6UtdpqxX4OxHcRmVQDo6aPcMAohQzx8GY
1TGsgA+JOA8QyP32O1kyNiClG5wOm/tVzx2b0lgPeisClryJiADC4+RpnQfp6i7H
lO+UZVEK/ZTQQw1pIONmVd1JRhbHgnbsh2IeuMzx0f07yvPA/0TtyvXZhinnXeY/
gkb2z6WSVXNlVOEv1itCmibaSCr1mjFroi4r5WcoDVkax6CcL6fRmn/5+czIm80x
t5S06l9+LRiyG0Zt7maBoGHkoFZOk/D18i7qrizoGOGL3KlgzuQRZuqenVjd+TAt
l4GuRNa6xYiTKiSKyXZvRHMz7wklmTHuxUrSCEYlgTgQQpLZnH/h6cTyglatFS4l
Xc+zUmJ7I+8dXwdJSjo0UzoXpJPD1MstIqN8Vrxm2+0oJucbvo6RlSS8hc9ySuk6
w3Pyl9m4dMdJzruVXIxEoxMUe4V/9eF/5WPH0ATPvdSLwSZoF9VOw/yCMEOVn+58
LMPXzD3mDwaE9y/KGicUMGCcjuYlHZWO7TO/Iw6VhWI6j8wCe5hhL0rShZlJwSi/
PhuJEoHEHWmqjBhnMEJoFuVuW9b5ftI/R4pH9MCFYHAQrssda0WerBUp3x1cJcZw
Ozm9AZQaQ+2YENty/q8plB34eI9OElOVgwaXJiv6S/iYxxmDM5xgmN+XTHJWlGyE
EHu7zSvsZO83J/g/GSgcxvIxE8p6TLIvn527+SUecof4r8A1DFUsmXv0ExcxpgqD
1eBwVlYyUDiax7NsOq+aR6P18j8IisHEWt1R559TGkPx4xhy8R4zEBzewVhb1InQ
Ve4bQEDeoMDNZCbUjYLbFbCTeJapIYQGe4rba14KzPW1ul5fOAo2o0r8QlDbKi1/
R+kaAI/UWo+B1l8OU6SSY7/pq4mHLWUVudagQeeUsgx0kcUX8ihOCkaHzef0WUOb
xS7LPkYSu0EiN4nvn/sG2wpI7g5rNDH+b+eXQT0fEmbvXmdg7UvNLH5CkJ5lWD67
AvdEDHWJN1ujoleTa1Q5WTZJ3UpYQEIz+3XWybhhon+kiU2RasNJEXW8ja9ZhB16
KJlCtuzDhshqdoSSezYjuLHOuIjftUnEaG73ICSEI+fDppX2zr5K0zc4COdfFX29
j80Ik4w3qsCgxYIzDBPoaE/x6rJYpucHH6FG2yUiy6/OGUqyL72SBVWcgwuOoc+1
zo5ImxVpAM/Uk3C7uwSlOA56Xh4LHjNUc1XV18qqh221AiU8a7vVpEw9JCQWAb//
/AL54gVFk+JcDJCnKW/t6THWvzbLOZeB4VJ9egrpmLgfx/MwkpWi5/B51w+bP1Ue
2FJx0PunoKVfSM3O8VrLTM+lSSQd3V5DrbGghg/HZObQR1m+KVX+MnMvr5vKqowa
aCBIbNsLWR4dmBCeD87ABg0s5DIMGRjtrI9LK1Lfz02oC8JBrA7tHUvDrM2hvFqH
WavTiHqPKKtf/ozijcU/ashMa/21sB+2bEVIyCtOWFFH3OEsBQ81B6AblHGv7Ztv
XG0ffUsv7+5hUwdGCqL9L0KvQZ19gfz1JyWrDJn20UmIKyVHd23G1LFUN5NTK4ho
g28QB4QCHCjk8Xr13gLCTpU43vqkomOrwejrWLymidRkMwC/cPdbFZRVV35/D+j8
vB7bu9QNDX8ilRL4Rcvxbroo7EnSKGeOHAWV3enT580fmDP5qplTRJQg/SoPN0lB
unRjmcUF7zI7xdtxtwRD6y7Fi0KfZrsNo8wjGrAzzfxfKnvL+uIy+4iXl1nZaI/+
sB0O/5C1rg6I1L9vkEISXZmT5zWc8QYuhc3KMXxx3hxuzNQgB0Z5DGCBRSKBrARF
6LazQ/XvEg9KfcyQTw688Vw9L6ZTewIQIHvzptIG7E2C7PKysoEbuImXamp1JOv4
eIxY7hUszYMPdXEXMZWFM5f23iuysBtm9HMqy36Gy1Ek3GLjLXCT4XqEcvWjo1eA
ph8BmLhfYlP/6hD/IYOKMHroaJCwlNNMnUx4XugQisboFyYyPnHsJN1s0VE3yZVm
LmHhzGdqeyCM0tbnGIc19XsfieCxlhZMNxFtxfB2SP4vR8yZjUicp4q/tyDunLK1
XDR/Je6xpxdlW/pikwOOg+Ma/P1qL7v7ZuYyqvvswj2QS85nlokb/U/G2xri1IsP
JbXLdmS2XciuqlHXk4OEgbVTMozbapEiFI9PYupWxOrVaHA+ktaITEI2kXcgbzw0
eljI7HGTyvDKJFzq6akZLWocAxpJWHNtMzTSs00AbIxlCHcP7OLx5czG2chivdPG
isy7si01POF0ecatEmT3/ARJHZnQPC55dThje0y8GqzHefpHWoRdnVc440Qkt6Db
aazChIGXaRCYLRptfE8f/8iwL5++qbIq+MCoY1tOxcK+o3HRuACt7v3vDu4v8g1m
FyJg6TklZyWgDM3njnTNhGiLk86ejO++NK7GhNQmek8/6sCnzNStSKLw/VfBo14r
lSuGTvpCZVhSKnZnfm8Q/xXJovQtf9huZ6HifGOBVXo26NLIE/rpyXE9QngQKUje
bSJbWw5+ANMhywfSAHyeNKFngvyPNN2gdrpPb3X4TN3S2sLuesHduCo8VqpCpdrp
IVw9dq/msE906T3sQ7eF+lCGMTEc7Cxmqq03tVUPCHYaYdcHu6eoYITXow9yd9qJ
Xo7Y8Kp0yV+C/Q8Xrbq14PCYEIUzwWSY6CY02DQtEcFgeD1bmDuqVTluekgPUYsp
5mXKOO9M18+Tp7VdLFBNKh1A+81v86E+GgPh8gJzUICCSiMXqhMC+KwEi4bD+SGR
3mNHlwAA7O1YS8ymYGkgUYZElkx+ecQHwB+3AC/X4zWMJphdRVdV+A/1WN1Ujwsq
bSW/KeKrKDv0xxg9HbU/IEne9Fs835RBUjNBBLtDTiB0kmbJEcEVhSa4A8u0aPNi
E2756s0wWR+9eK634oaJQNIXRr2IYYuzVCqX8T4m8EmVn/gtOkteUaHd/vfMxg9F
oOVbpTZkfpsKNplvIm537yHNgHZr5uan8PXkOfHxDTv3uOQBhJGLl16GjFbcP9Cz
WLaGmOnhYGQ/gh7YGcLOH3WLmm8RRWFkIh/Ar70C5Iw+7eUgT8SGg4bnW1/dTYN7
Y/Pb013bbd4paM7rzUP+Q4v1ndfQBr8MxJRF8sP6CnqJb3UOz/6QpHrKxd6BuVUT
hH4FXi8an3eUGPSWImdQ57gEJKh1/hCEQok7KVbYJrUOOcE3M9NMJ/6XC8Ze6zJq
gUDpyx24wqoI1CHSMEg0Qlw28nd0Quvp43lRWkplV9fYrOK3TYcV8uM2aRpWD+F8
l9Gspsjt7H0SXAIAZdnVFruQRUJxgEGekgIro/hWDczMDa3zPuhau/K7Xt/JyYaD
cuDTaG20a1oJhC80YHZvqA5kEMeniYQLM/FVfmMxfe4VNSHneemHsj48pYSihx/o
AL/VGpXATtEVlcyWewNb87MdCPWDwxEUY6xLq4IoOoWj2fzWSvf3o7SKLQBqj6hl
tpH5VgcABGGgOXNOBtEzpU/++YAruxihB/mH59SsICWOgFUad1YUJHKAzQJGize2
38m5OCYYPnCFkh77xyDJJCwwKz5NadbSrZ54/OAhAYwbSIK6jKbPecAnmVKt6YPJ
5D/qKShooUEqIXoTJFbgZrFt5Ga7MtlYCGGOy9Zg2upuIKDy2cI9qjHUxJEoAS7G
ZdOBtimjt1a5KoMrjVK/cRJ3NpFrixF5Ib+C3dW5BertejUlGn6SrSzGPSwPEXDL
YB3gLf4DLj9OeZRUuiGV2F+Xy2VXKUGcLksyMv/NDb9V3Br5gYSQUE+JLGeTqjtC
n8vzoH3MTgddaFTBubGAmOhBjY0iL6QNHZ2AFua2Vlz1csd2ELRQdahv4xmURHRi
g5zYFun8zW3AWXNI+3phSOdzBoz2w+EdLbGZWvsi5v6WRlH7IobKI0RN80A4KMcQ
hs7hAjs4FQszEB67/ZPebufxyinJh6b2T+XgaZW0qQrD5Rq948S39xMYAdN02FqI
ZCnL4neynJoxmFI8X1YiQv7jjAobr36XwMF/n8KIo9yoHgswboe4nXH2pRVw9xcX
UoK5Pp2c8TR6LTey735zMDgqovpqnQYYICgitUaiP8MuOpV9aqlUqylVDAvFT9zu
YdiPmUf1N3Zun/JHMK2hbuGaOwSDJEaagduifT70XVnIiAIKDIoSG/Gz8H2BtLSA
1D4Zi/dIKHky/HKMgJk9WiIDSj75lRs4kgXH11dU14OkUYrs/psWN6PNxwnRcTQQ
9flOcDfl5y25XMeZjOn6a+8zxn2UFAGZ3Ge/RHZbMcHRFEKWrSKMI2RD1yppfg9H
FrJ1jPPpnrIloCLN9WgrDX+BICygYqdRxVUdmWXh8T6X0kA9g60SueJbbEjmpjE9
Fn9BJgYk1jS7a/CoHW9ddDUJ7dDRbvBKzT3nZnu7HXvjN6ht/QKDuO69xbbIBxC3
4e70YGRNRiLKRKp+VBBI5/ZZUOWrtVBZC6ogUVVhdQP1aM5UvYNok+xmg3hwRlW1
YdWCsQSqGV9XOCTuQ0Pdw8ukmn8g49KhKAWlH7c0fwqltE4f2gFJLpbRzM0JkN7D
LLk2uLjtshhJmlsAC3ErSgO+coZKHP8DksW/6sOe+zNuvTFTrqvssuOoj+I1Nmth
PFMpKV4PsWQnpAPeLMSJMjkA3UQFc6i41To2qrbT7YSjyDK6NFcdVrCECv1hyEBG
urGoHA9hij4grvSiE3uuyJ7THnROIflQzLzE07ICeydj9UWWUxxMeybckXTlynVU
Q7IAq556EEo8+8gbT9+Kz74Mt0WGnZgT6zO7K5j0fACnHOfPcww3bnOPeFXaqqku
W5yZ18VGHKJGsZPchyqV0Mp2Ffd6dQ6lK9EFMCb8T2iQWRKILKtXB3NDQck3Nalb
n46tc/a2kGamA/kAldPs00h0UsAQ9Ma/zRFurlxFgSoyEk+RU43rVT7PREcOD/tR
xNY9cirhGq/hxFDjHm4GwRjzCYjKlutGgycmN6D1wCU3KgDgbqLqhMCO7bdT6dSr
diGVQ2hU6ogjkgk3WkLJLhrqncgUJN554kmCDUnOeNKEieSIFZ5t42GDbvUjjhma
LG83XEJ9Hlf7dc67AYZWv6nrnpVjCp8A+16XAXJAFXZebGhQIHyN/GndXzhy5xLJ
yr7V9EQUSAMw8TdDiqBCBntvl3W1Z096rzWbN0eKiynt2YqdL2gFyVH5xPAbzXN7
QJgAjn2KsAwL/bwFb3boJBprRIjgADuBUlLzhBR/Jat2N2hVcADeOHCy3Gq0/+uG
rj6jxGXOvgV0zWUk/nUFyIDjUAj6S4FHVWWKTXumomDMmENlHX8z7ip7fU06xjSx
WUrTOqcAnFD3H7PZouQPMPgKRs8j83XURcNUakThAl7RTosrNwwzHu+qFBodSxDs
aQdNFx8l3mldWE+58GthF/+3MDv/7plvOKFRuaNBTE4vEoHq5IR5wQWJRH0j6RZK
1dQjh7tvqq2aWPO0dVaQlh9MBht4Vcz7JHqTXXpYxqS9mo8iLc70HctzKmH5ntnw
viiPNep9Ug3BdLb8rr64BO80IIOVSpkmp5ksEUTaSevFfU7TKH+mI86DOFiyZYpy
IqreL3TjYReOG3BHZt25unl1n/4s+f72Vi9B0a53itCe4lGxgw8U1B4Xa4c4YjDB
aSUacorZ9CgiTk7tulZAB4bmHNlnWBPPNnSMgYY2JSwJCZjIkuUCnw34rMr7VGM6
yEQO7rQW7PS6XHFyofZYr28kh2jAGye1zLceR9ibrk6mLJag3CSx+3HwWJrWZAO3
/YB+0VIh1+bdJf8ZNpWjnYqPRuGnV91FY1kR2fOxgaDx5kfa0RsrfArGMpOH+t9O
Y4/iTQMkKql7c6b3APWcJnCRczbR4U4+IvXmhvX2L6ZYAIRzmjXv6lkdpB6xXvq7
cmAYpQbVbjvDRTe+Bn7Gwstw3TTPGQLXVH8txzB+BJoCq/g6yxxflENl1qyW+TQw
3Pri27kd1vdrnPucuwPaEtUNWxM6Fk+nZCp0+uAY/HS4Tg33QMgahM7PxQAoL0C/
cyOsvRBKeIewvYXwHZmYH0AXaezRxKPrN2hYtK9tWpMC2EpCK6+Srz0/qC7sj84d
E5y6d3Sv7DAqAqdpGmSq+cGnFRgEWHMLP93Jw9XLqqHU7mbav/Ux2aYY/KV+Y5HO
nIgATWjxOPylv3CMgFNltOfa9/aplGz72FkH1jLjyT2GdYLPlUYijAe6Tk+d1CfB
3E4cF0SMYE0MKTCLMTbguI2427kedrmJk1chUlJAtpMxTFseKAUFx8mw/jmjy0Tb
BZKO60RNoE8jiN1sFZcaNqgA3q0aRpHCztnLXNTVhkJqiuYP/1haFzWeXU9uJ2kK
e8Ojj9gQ+czsYydmLPDE3A3fJ3pB0wlrUh4g8EDVLqWlNsTwrz8AX9C7Scdg/TLl
bVL/0ejEqQeRZULQAYgducfimWxjqem7aS4zk9Y1u5IcIY/QsGBRq+vri89fDFAt
cxsmYB0vd23VvZ2O0tUszQW/1kzG/nIX/NyVUURaYhr68q7hKaRqQ1GItpP+PqcP
P9yvXJIFrFIWn2ZZx0z9C79wkas5026iowXT3yVJKDw77Dmpfh6ValRDN3Od/9cb
L33Fpru5O/UlO3XMu7rJIMNUYfgAosViDIe3aKRKh0D+xjeRrFWCnJe+22is+FuI
SAKyB7ZmcpH9bSwnCdxVh3aVSdYCooKUmGvbRRDNaZOTS4/iXXBwLSqoCscUnlb7
JlBcUQuTz5fCEvg8trXfH2m2A/Yd+yAl+8GC9gY+g7DlrFq6uk7b6Xpyu1Ptsaen
`protect END_PROTECTED
