`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zMOl7M6blxDbYpc262SGjH8uVDAkcEZrJiL83K8HHhsObLu0Dx5djVGyjAlpVz2p
bg1E9Df6UZKE8b9IXYX7C2wfvRIelczc/4+pW8IrXUksQtmc5968mSVoMD1UP7b3
Q608ggoYL2thW4mXbhAySeIfJyyCJARCy+MkCBB6BUk7oszfXz6sByzfBWxQxKZc
6xm1Al83DNsy8SU7kI6rxOudW97U/D7bx0j5ZVPpiFn5cHs/qCoxyzDwy2lVZMnP
8fqIVjrDI9zV2ubewuwGw+gVXM8rL/bmaVoEhSla3KyuPd40s4snSVRI1Obfvi3B
n5vBToNtJCXtUud//jzAmAOpJuzY2zjtss5vJ3gwWsHhS0mMoV/kXHCnd/6HfY1o
DH6b/vJT/tLRQN9zWoqtw84h6JRPwtUth55V3zdNWO2Mg1KsAmgC3e9yRy6GEzKr
/fMy0tRSAKVk6ouz/F/Ed8AddtNxfsA2a3CjXprrGk8uHImQO0A5dESMYw45fV9v
DISiNa8siigEpR33N9LDvIsbW8RK91KxgJuU96NNzx6lHCjErDkdk4ptJ8MB0YLa
3vi+ZfMFpodN2qljz5pMrA==
`protect END_PROTECTED
