`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zi4MBZQcUMzhyLO3uaEQxCL3HvjVbOygWDJLy9itzfW/fmvZiTC9eKyLhn1Q8C2I
dnu47zTTbaaeZ8KgC8bVEClsbOvc29e6MbcnLf8Pfo/HMAcmjaau6g3jaqEVjCFy
ZSP7AEAa8TqSCiHOz1zerCAtkMdZV19oClRdDNb4+7H4m2n2KxI6CnpgsmFn9l0H
VH/OlkDa81/FGMWeLE0ujtLWMAVY/1enrXSV+2yLT1yS5pBV8QyBcaCMJz/I2Ct4
uBlMgr4bcmmz810i3R+QAg==
`protect END_PROTECTED
