`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDKGXl07Svssz9qeHygpcvggffWEDyuH6OFdo3Dl9dxiFLz788ckUizUSIavXjqp
4mMjIbuTDVP7DEqgrMfQ/A6FX8gdxzx92xtA3VAKJbMl7TiF7HNpD9/TYxfjNUDx
zM1qBW7/mrjhCqHgIK/Q6NaYtMwYVk28O5IUhhpuTCKlpyEL7tjLd46m/cz9o42q
XG4xFgo7IqVemnlo81E0Pt9ZGadgKUXZHA7u8uIWZL3obA2+gZctYgveC14mjCiF
u7AoFu4t3grGT9kQMDm4qO7TQUTwXN8z/0Mj4ZmMLbCeatanUBlg4sOs0P/gLxBR
5rCJEf72G4U6ihSwqaozYQ==
`protect END_PROTECTED
