`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiimY0dtSYngJXKOa8z4M19QE22lFwTt5aV4CMtv5pt6opzuR+V1KReoZCatr8uu
xOd9GvBzjSbmQ6V1kASRywMxFuWZ5RQwMZ19hFVfZhUb9nBGQ2K5FBccN2Ffuhye
/dzsWlzLQOcNhugM8oANLpT/Fj0QLhRg//O0Ah1rmgEZop9E/SBirrR/isz05ZyA
qM0GVBwPg7C17SvFeTXXQWgKGzW7VELahaIRDUWSaStHG4rg8s5K09nwjmkV2XeK
D/SxzSp+uMFD4YycnxhKw9de0mg1UQmbJ85uHLv+I+h/+bpqUaGd063VMc+RRY/k
pGAU63bDumi2niMm3/dMMXRysSuZoZIx7sQ+TLuHi9XNk+QsFalG8UCxkxzNuFCX
qeX1/xRs47G34miF/PsImmP2LFAOMxv4scyco0quPAIG5/MRduK1JOrnBbg7TaIN
JvBil0MEGqG4sCArmtPkNggjHeBrhYNlCRreG5IvVgn1fCr1Ikly1FcqnKCeYts5
kLJEcXBdw+nncuOKwNT6B9dn1PSOYYxGFEovFmXDEFNMsxVkNDsefaaYefVPNuq8
p86uKlB3nNDfR2FkNGhoqzqEd+T68icEWGEF9X4vL14yFrjsdRxY3RPCiOfACYsS
/14UXrQhxFq9pCRhVoihWRdJkKSGDJG1E9ZgnQcYUlfXGS7jrqAgGgq1Xi1ZLdBy
tqITVkmdMNxz4BijhEw+F17xhofg7xjDFK9hL4eOc4Yu/H369BFrUesubWb9C5yT
ILGY8pBi+iadJQ+697blZZt17ESKYIctQeWHNWwMtNQ49ZO8gNw8kjMYdypQOrij
62Gwn8p/kxznrjms0F8keIJ0Ne29hMwR4h2vqjvspgi4qNcDgqSU3SuFU5M2+aMW
Kan32ginRjDiHeuDneEssb61IIECXe8bop4p25xQfwBz8kY10PwTiBZzxkxCTA3b
V6dK7a1siyfFeKklL8ZaDYxqJFF8zS7gVK/Wi+uuXTGpMBZg9/aqFHvZbrszxeZ3
rHTMpzEz2xA2ney242SigATXDSGlWaLKqa5uUvs3gG5+3kwZJkNBb6gX0hB/J1dJ
XH6mImrUSOfoylUhi3jP+3rXjgs1rmH0scOP4/I8j9vaPqAyFkd+44dRmdV/WHQu
wfTfnDR2ZUkVrbsqh3VJzFh4StK60tq3S9KakkRz8WprKPgbWvt3jsK71MEzq1x8
gRx7eIJeQxlc7H2/eLUO1RO1TUAgz8EESI6ngnMPw08XvZJ69j1HFDYvetcw+LXu
/LblvxaUgWhu4+id/pdaLaely5XCDKd31WFeZW/qUyTILwuWyRx6cPfBsBxr362Q
SGInhbzLsZ7QEvPLyGSQfPhQGWhPC80CcRGeESlRVgdvKOmYbbUhhUQ8odGeHyXL
8cOhcRqNxwzCUlNHAk/YN1nycz5C0eMh/Nu50xX20rrpOc5F9RDwJVS0zfAwmKUi
bVkPFSqIRABgb5Rg2bUxEakcEm958mh1LBK/e3fBeGYUZYkcczJ+8cUkXbusUitP
mdkoqh3iGjdjRU2EGj0B9lBXqqCUj+bqgaEiRoIsZany42MlO6vH5U1xBP421Utl
8g0HQ4069hwRW303GG6bgiiWHyg5O7RCALTb0Ff4UWvsx0FpY8jb7pa9nWFausVn
OQLPg3C+hBjil4r3bXbu7bbA+aLE3Y6MD3pts4aNf4q1Fmkzn31tNT5gzLmsQiWv
BbU2dNVm4NFFndAyqXRQU5BOLAe4+bcylyCHr4c9b1bgMEKTayIYKYbUoLyE9H3P
khk6Iw1wM/6B2a8at14lmA53xRvlR63UM5pSqcX5ALXMOT/wXcyeGUmTQmnhG3Rm
9+a5pZqaP6gwyFmnjZFEejQv0BIb6ONHOZHNt/WLEeZQoFY5wKSJPD/R3QBpupG6
m82bf5uxRt09TA+cDlX2ko5WBZbSVAJ53f7Tg12e0tGeAv4aZxIFPCwCeclbEE35
1op2VVDkmnfyPQdhUySb5Cjs4sq+mEouKjqRjVecW0BWiowQNrwEXBOU6+ZxoS/I
xxl+hEgPFqIo0naIKos60n+HzYm8wOeWIIX2yBuIhErTuBYxCsJEISdyJRZGRNDb
ywp0L1dhV/1k3dA5rQgqyrD67/fvHlbB+n3EKPzvTEMySdqT/gQeSmuXASJikjnt
M900hl9tKVHdHAHInI8zUVydxXarPp2EJXdEUwlzUmbno0VWS7ETbaLWD7t1MiKe
egdrPmapoQ0dejUaMib5QQyPJFKUPAmb4N7Pyhx0q8Omo0s/d4SVp9xxCryGRk9x
ocbs0OfEimwO6ZvA7TD3I0H3h0RA7wBISa3YDPdj8YRnIHdcP1NUFuj17nKTUNfn
Y2/H7V2WjZaheoEuyh6gyPBPTJ//XerLYOKdkUVcWIaOchuCTVaM0dpiTs3eGIHQ
uprUqXQy8q2Md54k553obYziQkxn7aN5MRShnoUA1eLjQw8/xDViy23FW/7N3/gH
Jm9aGKedZuAyJ0VIVuqxzhku3RMUreplUEc5Lyny+K3aX8DmdpbsMTTk3F/Ay5u6
deNO9+6cRUhK9BYK+Grmt8JrxJv+yJ90CWi35qlrRv6YugOCVo0+LVuqzot1ehs8
lvER9DfZSxu3W3GRqqAP+KJgNonqPUVhO98AbQw9K8mPY/++KRhY8g0E18F4D2y8
ubvVFVfLQaYNQPy53kwT/pcO8dEPzasphKCz2JyI/Rlw3Npjbvmdv3IcVtc1Gut0
bj2QTLGD+hMiW12vdzB6kmm4Zs274MFYEKagd0pcleNtZgmCjzt1yYxrc7q735Ab
lLRoIwZ9jKuDrkTtPmEzcX+CJbwfVe5b1KjbpdOBVU+UO+1iUxASqFzwGP6hP220
w2uXa1Yx2OInUbRe5c6mlIy+RAH1OveoyCoF1f5rhd+g1o1LO3gVGltZSor1B1eo
PRZtPwwKDxmEYfQC+j90xW3j4Fjavxhwg1fQ5XwUskfsDZuIjdJoz3SaNtJ0MHIc
9L/4XD1NT8pWcpoS75Fh02AnqJ21yI9gQXTBjz/w7bLn2/xioXyXYftTyqUXrjg6
X7UcQ2aUVbzQxAMU2aDcixF9nuD7zHioEoN+d1UewwKwsfRB0aXzgYIHJ8EJilAY
90Ka9U9m9zONc4u2YPBRo6jpCIrp/Kd11Gc+rsVaaqHagHVRmnPF9rRUbEmlTaTA
DrK5M2rT9DENCO3AiAiNPioju1PkR8Ooe9FVjyn6xoC/gLoOZbt2xOKi8Ik91uzN
IyUARLkW+7Ck+J0AD3/Cfo/VD7RCU0BdDT+y8MUh1yx1rVX8HpC6yq0nSchT7GAw
dV6yANPgnycvbLqB/AEMSUQEJZpf+GLlP1ZXUhQerUSG4Qgu/jk275dlE7ZpHKPg
AWYxNodQx2ljBfl8iVz/XPQT3olAVUbcYMWGu92EOOig3kbci+75awY0npnvyRQW
iPs5lLFWTuXDCCT9RmUn9F+F6DnzZXsmCy+z4tuIQr3lIXZwLX6xNZoDESdAdbRj
JyhBhgzRNY7tQU5AVeLHuRRHnkkHqPRjp4kzcNhByE1EkORXtAWRsXFSrT90J2sF
L3e8ZU7Nr4mZHkRoxoBcZw==
`protect END_PROTECTED
