`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YO9gFIXxzk9UGmadU7w/vRHXAfRZJBIUwpDDLpFppDUpB6xp8PGkfkjaQlDwCdO0
xyCgNutN1v98d0Tomcg4ANt8h6Vo24ra8F60cRVnGGjSwC13Bs0H1bny73XUwElv
7Q1cEvqOcd5Bb/IR1MrEkjn2kra98fQw+0QPto5+UbtgHKatGGZ555vypEP+aR5V
yFDx3HMGZXZ/fET/ad97DeSJzdhbyxm730hmJDO4c5vmHUV3aGfjRN7F2l97owqT
Zklg7UAWV0G07QQ6sjf9qjCay8zqj+c1QDluzsHReNZE7unqdo35Mm8JJERoRzJB
7XO+Gro8kJRF5opHzH6wAt2E2j75DZMFLWYm7Bf2U8IyR5Q7VQvvyDSksTCVTscU
RowhpukYm8W2w8WhqBT4iEXRqccjwg/V/HBv3tmneYdRUmMTvcDNZldJOAmiJ9AH
wYvB87HDSz3fbuIH4PnR4Kx4o03nf5zEe7JL+FSTluqe5lay4rZT5boD+AVQMCgr
D/wXxuxeBRaSYN7Z2wCrJvNr6deDg1SaYnrRh/T3ku2kNmCy6gFFjMPWZDTtx0HW
vm6IMBnDbIKb08bML30/E3T84cApQZvedjiMzVZWUw7bajMH/1BoWpIxYXXD0/e7
1oGARNccyeaZfZZbT/rk7kWbh28u6GqZEvKGeyaV4tlLlHcFmOZbjvCCY8CB8QwJ
VfRxgjKj6r7nyZXEJckFFzsq4+nQ0Mhdv/5O1VhWNlY=
`protect END_PROTECTED
