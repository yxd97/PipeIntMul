`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PUHFnzu3kXVdjQvs0p4GRW963tsUyEcW+aKo6sG5/2/dF39mXVwV5IcTtBYNPEST
zQMVx9jgEwYUfNUqQGV7ugRHNWmMVcr0qeSaCRm38oA36q3dh5sjm5lDdZwqfNNS
ralA6DpUtvSexmGLqUlcErtKh0RpUclDPnklcJcON+wvbbk4lX20FdHJnAkDne20
mcMyb8SOOjw7fpoVWW18/ekV4qcQna/wiROrbu54dkjI+nYfTzxzRuqJ1uoLDnfq
FhUFTnVE03q8pidT8klgC2+FgpFsRQqMj17DzxhIyPs97ceiNGgOy88BS66lwa0i
+eXitvlSuqaDY7CiTJ3FpY2L2AVRRsXaqyk7y9a1RNVzn+8VI9klbidoF929D2+1
PJ3oFUr+t67Ep9332/vXKxywUCMfbMYLf3KJI8qKUOraN1IHszVMduCytPIMY4yw
kNzkOPzupZw6CLVJOLRundFGoorh884wy8cSadxjCHs=
`protect END_PROTECTED
