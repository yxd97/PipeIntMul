`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3kSmPEfuVjLTGKRgrjAbUAwO6HDFb3TjNT5a4rArBZyu7s32G5Mo0ORfxcldvMkG
dCPfD8v/OjbDVgT5R5l1aeSD69YqXS2y25BJsxdNlvJ/W1RT2g16zIJ2b5hmWx8+
D6QegSmNpYmSR1jePyMsqf//sZ3ZS8irHba7Fvae0o2yal7ReC2D9PNPa2F5u1JQ
JoH91H4rWHYtpAB9rVep19NUmPMLtn35SZyYgBn5mgtZ44hkHjR1dDDFaNyRTGgx
hPbBTCduvySX6jUsiVXW/mDieavKDRdjW0h8STcViN6qMnZkLVh829MZmRtgeFb2
DQOhNZq3MGE9RteGKIlwGcckY3N3C8huGpeUuxH83hrGK9YE3MkZ8DeqaIDxxtnC
crRkwlbFNfjs+xeC5yqUZrCLfTzVoF0ZUpfcV/TrKh44TrQhFapdeheHgtVMwAu9
iljhiKbztBOWApHm9MUmZ9JMTQ2FJ1wULcRXtbEn1Bs=
`protect END_PROTECTED
