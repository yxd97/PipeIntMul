`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X8NV0xrxNtNeIC4OaSVP5P/+ulXUO1UcInoPSZMkq2BfjU/aGiwop5VvHnLbQkos
AjfrzlmEUPctBcc9DBycbuiaoy3CP2KiSE+GPyrsFYwDPf3xKgFtiVFw5c4UZmjr
jIRT9bBd8lGXfYLIbfgscI3Uvd9Idu6kNq6IZIX9kc0WyW43+heJwXs1cFN7OqPj
nYY/rtuAbRIQnjaMe7k7U36S7Z1VURAL3PmkcTN51CJWyN65hlbop0uPdDGq1s1+
lpewgRk7BjlGeT5ZuxeKxpFAnBLhlC28sqLPojO7W3nCJCkHH4a4KPr8m65njE73
N+dp4eNk5/2XzCXKisRv6Y0GIBD8q+s8XrEC1ttZwAt/ENX5zigRwVozX6UKSiUt
MTIvCV6fPrzoOzN/T4nD4RN7+tq6pecZvMOEegH0whkQperZiS7C8hRuoYxK5584
YWWXT39IyRGQMd5B/3ZROxy1boXvQMiK347dtbgtZtem+mHgWLIQuqDltOeXuiPM
+pvXG6urAfeTkQUf50+hwsZeJcytGbnx6vtdLxPcn02iY6sX83TjrlYKGSfeyc3V
OPmOB5NZ0rj9CZ3N3mEgrVrcaTgY5/PqbYtLBRj0HC14LRlCUVX2VvHiIpFPxj4i
K9Us4rOgvp6dQDtC84V60h4eibZYDjrRVT12omk43LlyssMOwzUyiOaApVvwoh2y
0t8sareZ3SbMLsY3cd/SCG9/l95LwhB+9OQcUuJv8kzADDUBDwFXfuwWFMvjpu28
kI928aCjuAcicbYZHGBBrusLutamJ9c9lSlFMSL/y5YIKfL17zbKOE4BDV6vyEna
dutiicpFWPYb6FbC76vHEeO27htyQcd8vr2sn7g+cnkRfZ9CRbC9qGpHJJxqak5b
BD9+i+HhCsvXctMOY9GLxVwIlBuvAoYAY8t9frbFxDVD6voMNpF19RS41BmhvB0N
ug12B5LL0V2fLS1/bDc0Goxl4x9zHcQXo8KmOlB5GCH+ZGrriQnde6+Z5m46JQh1
85wk1YzqvyWBiRImN92KZXSUbYp/ylIT0YHo9tKI9RNnQzlIMfNOZSxWHrCnLLm8
BNUaH/QNfensI7ManiLDswj15+5taXrAOA0XDILYt6Q0MdjC+VXwmdCZbw5eMm+B
2bjnZ0k/rFpQqZlQBsAfdoFW4G6zPatP5ac7ySyNCefQbZFroyHE5iilpDP2dad9
YgUCI1Z5QeS7X7BtptcnyViYbZuscHl83xMpqP8a+2BW/jyUODYn/ZvYIn6+Fd9v
o++icoALFtipjmXePRUDka7zFi3tjqMPjwl4ePoyVNilKWUMlUQDaJ66JKXxz5kX
siwkqjFasUzMikc3Dw39RqguAPjULeCVjYf0EvycCQ1C98IsTYPfE2NY5+Wpa5db
IsmqFZxXSrJQwuilOkoYw4b1Ye6tlYYxmuxkRG2ApRq3K3pSNaBw1JEn5wG1UMql
Ezaa+QSGC19E6Uyw1YHjyRZVfr49Kvpx0pd5/15dbIu+i+X0jSGZ/gMqcdfmYnLk
9ZIrUhuAFwFMoWE/1y6FrTR7P3/B4I/eKe3JqhOHa2XTZaGCHxJBdN6zjg3meH1W
P48LatvXpxE+ybBZWtzZak8cvCY0MoZe8i2kTuvqifj0j3ojCvNOYZXEBuAXNThM
Zl/N74MLumQIwoAW62jRe+hYwqQFQxbzpkBWI1cD4erfMuCfgI6LcnEZG6sZPPiJ
w/jzwvhI83sdoOiSKprDkQ==
`protect END_PROTECTED
