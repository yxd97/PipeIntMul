`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pfjzZNJOltJXFBhl1niGTkIfMgCH+b82+RheLzE3HkbX2FBVGwQXRks/blHGjznM
XbZIwyhVVwhJXJN8FlxTtjdu8mwyPYRd0pSOAd6YmfveNMuwykrWOEVVSTZXvUV8
jDdNGjVK8kx88mayaMNG65dG2JVOTCQ31miXJ9PYmCx9gTWgyV7/FMYHYxQOBwn2
z+1Jx4zLPxxzVSozLn5Hfd7qZN9kuXhni2BTs0zSdYCTdyaR8flylZF5rqnLPUMp
fX2OoeFCd7lROQewqhrbERFqm53mpSbKAtW9cGyE1PWgwkIy66SUYBEphmCwdvn8
Em2NIeqcpcbNMXwX+HzmER00YJCOHwnnex4+ZrtWhrM0nhV8GtgFOd7fOSSoJs2c
FtwDdtlPZt/VF1Yuv9/OpYDbGfbxuk4g0BWv8NUwXSa4zOAMv4fvLf70+ootarrN
/ovzuAoq8FX3xyB3JLr5+sHGO9sB22x0MnX16sv70Dog7apqCHmmTQc/dlGP+YnD
1jBPKYUhWt4BTVxBm18N8E71MALT/Vu67Flw0rliOxgaWqaPEXW0SnEovJhVd+oy
AbS0QlEUyLi0cnK0TEC8Z3odlr8fuB0R+2NEgqvvN1XTXU46CLhKZSKzcSMOYCdd
egGMt6jBfjjhc55jTP8zTw==
`protect END_PROTECTED
