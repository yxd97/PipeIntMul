`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kPVFpap83Xk29PWsJF30Nw6E2Mb0H0rIJEBmtkpc0p8Y35CkAeU/JmfvtwhiMyj6
l53KcaD6Mr2sR02xgYTvywTCbTyFHjw1QpbqFAMCU1KYkEvQzXpVsmOSjFKM40Kg
dJSOJSXePZZA1wewFxDsEik8wFbj9+xDFTPCDovWAMju9wANqWC+xdtDVtgYmUhO
fKjr+tlwCsv91kfPGEk5nGlLt4XdBWS+l7mxwh4Lr5SsGLiIBBXseQh78qMN5cGb
4dDd5bB0/bESDamRdiPWb3IrJLFLZwwU5RGsA+DnJ6Y0QZ/TbA9KcJxgW7+Bhe5W
FrcSL9miDyCX1lNEwZTvSA==
`protect END_PROTECTED
