`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9AzSaWMV+An8NRkHel7YW0wrGjEZ9bRpM2MvjrhpViNnYe00mpz6IdaC8oAplPBP
aP93p9ZjBOypMldtybTv1mgjVOrOvotGN3RaRsqGx+/9FHn5Wx3Rqwo/HRdAkZrZ
X6TjYnoGxVoy57txl/LjdhYLZgvbd8eCta+z2oFd+BpBeAmZ6hSiQt3ZjrJoE0eH
rBcaou8I676pLdeumBMa8xrics2JFDJFlGGc+ssnJpfR8Zi7QsBntbACynQbpVeZ
9x2cOTDB5Upy5J59K3JeLrUnjBjrY3G+3h5FhOGlDGbClKMbQgTRLierviGNQbh8
xwPkFS/kdXxR/9747YxmPkoxlNJh1btx0zElIQaNmN4f6d/zJ0eGG7MvV+vJWdIt
Qo+LrC1/U+oPL0HxW5BkuPtNLHZIfj7uCtuQX8CYm+18P/1mXu/Fs27m9Ful2fVY
w37c33toly83GdpP9Elq+sMewvKXdyUtxfE76URFrLpQk1DA9UsWEq6P9tfRc5iK
pvHlZ0umqjrbEGe/QM0BPwhIX+pkEPeEiiZ0vM7XL6EtBn8LBfmV/jIpWneidRAK
p3fanS+Rawk4ubSeAb4qJ0A5hIWDembjnSyJRCn1i1mDOQweuPWeK98qKqCKz11E
Pc77eR8F8xbVgxR2Y1EvMIzLn89KtTLcKx3rJCNfdlq1UFA7imoKzDNATBPjHQDB
D2P0Wogvvx2XAyFY5KHaDsXPqR46KjVHmfEgpobkT/m4/nRhkdhOEpo3phWgBTBY
gBkXEok8u6KtouyPGMZyF1Vis1T9fH+Y6ORnlux5gG2ZtWXJyvpwSCwV5kjhHSoE
Lb+XCpPpEZHGGTX7C+XIU+trtJqPbQ+HX+1MK/vHwU1iIedIA7OolGDZmzieR/sC
ZMQxe0zZ8znyJrVA4yYYKzVIle/5MJJR2dJqBPSD1jyzQbKGPUdIiSfjCadIRGgH
JIkStVnWma/08ywQmCxQEZUzow33/aRuOf836nyeIGZLC+AQz8V+61oQa/f76gSh
NpQFhCOLccK2n8w9yqRIs39+GsQ0XjZno1FoUw4VuK2Wgjdwj6oC9lWE7dcHe3PC
+s79v8y3snyT2brmgLMUwbZNdVaIKyyw9XykZaak5d65idh2sPm84VcqSvbBUngJ
CDluaOrmjRlpeYvZ2+FnnLwL+eWsCD0YqBGDmnnBBCRi3ZtKthXgUYqeBwQAhhiN
drTHns9PJvGcAVD4/Ve+JaHDCZdW1XLROrnND6n2PURExtWYLZc6v7zCdtKT+KFZ
8Nt1WXYsPZbsGKlhHPU4fmXr5SbQaFqJ9sWgyFN4LkThGKCvYYM9UYa2kiXAyVY8
uiRZTH1tizVDLC5mkhwJiQr9fV8ubk3NcSYrnI5uC6Dig7pRehM1FgphtLBlyq5f
DWKrym6kQD91wfUUg5l7TlY/EtvF3iz+HH1TatM5Z1U01o9al6n5LX6xhQ9B/vJS
aQGgoNA7mUigjMjs8a8wmmvYDKQjBCWAJSRklo4eFkwQxZ0+vApFZLI+ee+S7w2N
rpWsr2C3RPlJIV51SaR/MVuzhFRSbOGSNBOB4342ft+CSW47us0RCevNpytvAcVE
NMWXxPWLKwO6rtjFav3c1kVjSYQuFiF/ZyXSakbDr34Zwi5B88MQP4pBEV+QNyDr
+37bGTioKYPftcnVr99vBfeubpJjjnXZsnJYEtJwiidPmoRxcJaEHCpU8qLMf6lf
wMpGlXNRLJ5ryM0hvIFHpKziR5/NIJH1eVS8iakTD3QEd5Ze0BFTv6tSILxILjZw
Trj5WR2DHCdy79RdY7AWJRGdsHDOc/IbEnRZAhBHhF0=
`protect END_PROTECTED
