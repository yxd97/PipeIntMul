`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHuUNJRD+msuAVSjzwF/UkMIkrTPUrpPgCucjxp5FbzLaVHK8ZXoA3L6PDs04rfA
YW3n5y8svUVIetlHK9iWfPnr7zLz5cC291WoVhAybERhENhl+d7hrJiTx7M+Spur
PU2BdJ4rFGa2XFICFj3RJ1yB6ihS9YBmu2K6R6O2H+GTFWVQacansy1jdlS+olCc
dXoD9ej95ByPAI5fIqGSWi/YeBcVdwk/W/GHB4thNmM2ZBK5U9RsmJ2m06NvPQWr
yrFcjURKh+cYWtfCE72JmhSSOx7LP/3yM3Tnb8XJIZD9znogG9yCG+nnBYQcDGn2
SIpQd7snIVyPbFYPm1dCRByrDlDYw/xRYqxkdLq64yjHmtVNqkwOqdSY14rKN94s
GUvJniJNtvg91OzAEia+Nhk936+63wxTQxyz0n+n+GbIXB3fgylZwbFq2FDGcf9n
Ex8BBM+ctrTknyot5TblJInCCcYcPt7THlY0xvRY/W20ggeI1MR0yhRL2nGCBdhO
PZNczBDTZFVOJvvqPTjLWsTIWJF+H/RGOcuT+NpR9nExqUGCUw7+lULWRMkkaXIm
3h+fg7IQFTED3FMV1FEN85YWlt7tMF3mrTnIoPnBfA2dXNrblAfpU6dOzPYfQCR1
eSmVzp4CXRrwXZi6Cl9eWZpUbG8hqlkO1KnifxgzIDhrABiK5j9EP3ZQFWeThEy1
9cIByre2b0BN0HXLkEGA5ROjSFaPs7uk7MkF8P8322f68fg+eKhifQtXgU04d9/0
moB/MfsgLXzwsK6ga60Hq4LzNM5gqNyZ/uLSYfp+WDg=
`protect END_PROTECTED
