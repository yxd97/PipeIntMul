`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5Vy9yvYJ2n+L8mPCoC5WmVAJfKQpvGKEyv4pylyO93bBQ+kk2tKrO8kfNohVo6h
L0n2GazLeqQWjlMlZGRuHsq1SeqH8nZsW8Oz4vbJfdxqfDDiYsfHzhnaskDDzX8A
EwFDKjjjrPXivxknyi+iUUQcPIPs3m8gcDw7PW3SruxxzcV7kA+n2L4Nn+65D0QX
2eOQRh07leVgMVjaICX5VzBzct1PPjTsMiqhbhAMocCWdkDiJyyhmQ8ebk0mLWds
4Q2tb25RM2hyd+qUHWoTZoJWXRMoDJOLUfSdIqgFLGWdu8/RHTFjT7YKZ7qqVSIJ
O4f4MK4NlfUve08zsFW5PBbvPV5uP5/KonzRLG7aVYcFgVQL+Hbx0SbgmrZoYLJq
U0PW7C6bXtCFIWX9Ywkd0Q==
`protect END_PROTECTED
