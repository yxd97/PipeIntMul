`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fEtKemg9tqs0/IXuJgfMHPWtuOJiPY5MsSldEVOXmZHJ12DMzizijz25MqhdBD/
YHu5RgDmwORxoD0TlDd4SicVTC7mAlWC5KVKSyYtlKXS8VI/08/8jktmLdHAuawa
wR6GjvvFNKaO4yXq/cgmNrpIWEkonzEMHVkg1GScggIkwvW/s3In4jJg5zP9WrBj
Tfj5O70KSANVFvd5clyg3meGZdDEx/HxcexnY7kCUmK77nrFrgK3vyph4V7waP8L
Wf6hbtV5NxsNL5PztlRGTvvumKQjMG77LS/gqvp7OmsURP7rh4xSt9xEi1B492uN
lJCa35TVbMuW1fDeLp52xSBEyin6qvX2m5+9JrcI9Wd1dQfyQ3c1AHJ9RxK+LT9N
6ngiGIVdlD9hGk/wiqRb6bW2I5dfS2kwReZnWUG0CCspQDjMJ5YPRzbanWG1CBZJ
rPfEIvJLs5yZhiR+9qZa6KcMXpGM10xPo0YILVJak9zTG7Z934+hCeiCA2o6RbHO
o4/LPaz2/R1uMybEpKrbVhZxTzU3ZgYixbeUe31j9yDaTJHWHAPVxP0HG9os0NfY
NieZlcE46uKeIVsJky0xvNR4xC1WfFD51CIfI5afl2RmdAmGMBOMV3ZLZFYLtV8F
Db1L/+Qc3yRPuJeQdroNhmfQN2lit6Bowm4vdWqlhggR6s0m8DUU6og+JH1lZEKU
FEwyLi6z1N8VUHCEmpGBd/7NmhjLwBp4WpnY9L/sPc9EwTIyWFMh5qBRM1i2CLBj
R8EOmwzQA5qmscyVD+Cu7+M313FfbiQo/rlOofwwfGO//KDReHm9jsEECI8mvfd3
ziCFkd3tx6KU2idzULrtPZaiFQ1+Wpr+zIN+nQ9QdDr+J6YYGiVME6GeS91bbp56
b6nhzty7DSvSQPcIB47wBChj1aLrU1SBQH3jJKKBOZVLXzVqzHmkRzU/0yPU2gsi
LrSxcBMtI2OHhf4o/URwxhgmPOo3ODYFuln93ZX/yi3gpqoluHaPVfOEXjVZYFCS
0Gzo2a0p4cQgn/5kibZ036jrfhK+vZhO6NEzQXzEx41HAlM9wwf3hbOTCQNm811H
B4VmwNu/GCcLXm7ZQXV3ofEvY2TPKCkLh0hl/VKOqZ0OfN9QcjxuwTRArEWCHY2r
wXFAhMCYT9apriUHBtI/4bLGxD/0wtnYdL0D2nQO3Qb1frt8ZAU2ZiPY9c3P8sDX
AsqgbEHlyPPdiRwSNezxBeCrhQVk79J8icjWUl65/RB984OdmskDGwZJaz2diAXr
vEEKmJeOC4EWvitdFjKaUxeVzeNcscuh4zPW+JnmwEbSy08f7D7QW6LAg7hpyhoZ
42dEHYQ6PZZZX2uMSx6Mh3AYL2maajJy47CFrxR0bSKs2SXl8JxRAH9xljye0qb2
/toRkrlE9Z0afgvAMqQhbIcOuk4fiwUwbD+YbATe7W8qfUVkyIVV8v35UNzGuawu
NqLr7Tj9P9O4hIK+tZUbUlQXxBK2eAjUXntmB9Y09eOFRn72tpU2STvpkdVFkfEL
9/ZnZrWXEuEyMSKRzoro7j22cETYmBHVrXOkn2q8XDbq4/h4AHtq8codarrqPqec
kjNzLq3B4otslXs1yXpD+J84UIbA2zIDF13Le8OhaSx54MPQzNJLifCTVFFZNdYe
91ZOqAXbTxQX1NFcBt0VdMc/wbDmLLn7HJIqFJFQgV2JvQ9TGxAkmb0Uv7T9Puj6
co2/EoZrckNhr0lnZsIREPmRkCiLawS83l44wWO+vfgM2KOCOoCM8IRCz7HimBoT
s+XJKGbZhJqCP0oxz7N6FFXu4pBrWLvy4pn76k0ecNmgwY5QuK5YGENZJhsyOQu0
aDfthmMUX83zUh4W+EiRzlN6EdqAMPJE+ClaKkZKwX2lTjjw7CVPNgd8k9hcKJid
23NvrDx5ikaRqUaHLAde4U9xayx4eLC+4t8rSyob1HUrlbHevwvuN+37N3v30BzC
O5gS7SKrgQMRR4ze7AZ2qkC67va8NF4VEZh1ymwXkw3F3BaUWDAkccrCAc+jmB1h
`protect END_PROTECTED
