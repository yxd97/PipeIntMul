`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yz6hyXzsCoqBaah1FgIzhproscQKYQ/biRg/adhmLVwqJh8Tx+d7U7lD3ibw0YaH
2VZE1pHsvZ/NH0R20jP99BCe2u4mYleKc7baA5VF7csv3TrcN4yaBNHwpd+podIS
2zlIqqEGmogggPLh/FukcJ3cPXYcsuviQITc+9aEiuhA4tAX5X4jW4v0iMQUJ3Ew
etuXu/fbgC0JPgBn8oif2cj/OWWcP7glP8+IQTS7l10Yi3QqZRqpdRam2iW+3Bua
qWJbxFRUu6m88Mei/zfaTuzOfh90ov0DKQ025gWYgABgKyIP1U+q8pHB+4Bhoufi
VSLTttl+TtcKKZtilPC3aTtIA5cTD98/0WpSjA/3Lz7PLh/uLMo05iL/RDXmemHE
ojJcIWnzWAaHIu+pMe/ZumgVdn8XNVNq/XJ1+04DKJXk5ni0OtANEcIwoLhAl5Ab
f0ofSqqkr22wLElvES+95YRxxgAnUbWlBqRzRcrQijgzdUSdXUBqOhQ+dbJEIL64
Xo+LZ1i6yEo3bUx91VsocRLquek6ebci1GQZZ20ZdU4lk+jhBVSAyFK7WHbttXQR
76YSTA41bVIVBnW3wmsn9wchi7YQaPUbbhX7g0PYsq5SjuhLUfa+MV/QsDUSVIQ0
b7Kfb8taUdf9bymoRff8oyYA+8nBtEU4e8t1vT72OaPuwidsy565KjJS/IxCcquY
nzMb6W7f+PLR1lbzYaftx3vMjN1stpHsHhDYexCh6kH52C4kONYTzw5yenkQKZNk
WHlUXxFJD3OVkxlPoMLTj3E2aI21u95e3VWtkK+7szhBzMbAN26/A2LHX7Ixy7Bi
wnikF2MPQQ6z6VNyDyvFIVxMQfRtVtRNZLS8N3SVXVfYPGMPW94UusVr+FPeDJD0
wizhHRDj+EUgz18E6quTnR8V2LDBcWHx/2fvC5SgrsliQuTnk5r7i1A7pLD5lf4M
xU+j0n82yaUgKCzX5KEJjdA+5Lt1hfTr6cVfCKMMo91uoP7wHdl3tS8wxtjbvIiH
1v7yCfu4pw3zXasEF06G3bJwebVi7fDIfk9jZTzY12ebrgjOPzvyJNxuEZVMIxCD
7GKIc+aOKEK6jYAKKt/NeHKZBcro3wi3f2PHoCh1wC34uFD15pfiSCMOlBn6vAHa
Hq75NVitIPtWEz6OdTpdjqAKlP515yiOwK27q7lTJw9/l7mQTlypFKxXNWkPzeUA
Z9kb1PJa0Pxv6T2RCGXHPXXwtqAMWCzozTBpXsiGqr+U1xbdRrzthWZi7KWFsyGz
2e/ofuNYa5cyRL3UAzddmWgEGPy5CcFJ+50TgtHlFfmWVYIVjjFfQygiq5X1yB6N
wOSnckFCNvForNOUD095BxKDSI8pxfMgkRjY5WQlRavpOKUpUTEZx5Q9ztlAPMEo
ItaUdRg+5WutNshhUiVeE5JgeiOkJKjYnBGY4vjXIkqODQW0M0rtrkiM+fvYRz0P
azqkjiY94yE+d57Ll4YbHR4ho1Gc6z3438/Gz8oxDXiktlaWZxMIlZt/yaL1VqM+
ChHuPrHgEpVXdylzouzW+mNsmXTd+C+KLncF6WIAa1QftgIi31Q2YAY3J5EuzUV+
43HiGOUuEvnMmKC4QuEQzeCESeHYofAHq9g2xP1Nk2QG+ytPC2UupEryMxmUvFIV
Pj8k/FFq1YueaqO0dpcYRziVGgE9OkO4D2ZmmsIYPR4WTPoEKr4HA50osdS0CWDC
eGSgBvAopaOg0wTrGiYFYQWEKzmNbAppAGUhqP0sVZtq9zP0/ogD2w8iifQ89H1a
eiXlxpN6pZ/TzuJno/S2dcnqTRoadO4iljNno9xekuygyPobGgJaFsTwmyyAmqm4
UlXwLxuiFUyc7d/Q19Swi56UyCZtcBiYQM02Da/PwadgACz0PjhEYslPvlz2rsNv
pc2GQYUHFZTXHlfkgRuEycfIg61nnZ3PWjQL4qTXdxFXxIUTGpx3UYROWH1nXYPY
d1J3mR63Cpk1360Fm5Ec6SpJ/w61B/HQsSjQQazwedq3Y9eMUhhwOmJHsy9EgDKh
u6AndLJEdkxkJu4UYoJ/dmpXi7rPQTaQJWCWykMm6VQcrFSbzOy5wUY+6i9F/DoL
VTWcyEF5fM5pF6qgu+Ej1WJplSEtKxwwxc7no9ZpaBllWUv+b5X6dtvjZL2BbD0B
y7v6sp7nwFdv9PFflapeFxNyZduxkc6JtxDPTKqIsvdozY7OFh51hT4EeodJ0NoP
FSDuwFaLe1bUQC8ytiNRqpbAm7CcPZmdVFIwnzBtkNmn+gD9CFfnLQ54NAaaHH00
5KGQE3kGRPbL3MVsY5RN0nUpXm6zUVPC3x4TbtWClwhOoiartXMwuQGdhF/ja7Jp
xoTOaGGHKlnH2JRZ0XC4sk8CSCpL3WsjePwLGWIn8G6H6SyXyFBZ2ZJpdDGJvwoX
7jLYeE+eu1wNjvAR44UkxU0JoipnIHs20zDf1DMHQCFK51NGGvdkgpGMuorT+oMR
fyN4sriHQRZYaEGVzxC1FqGGbO1ovpTcc9cQ0eTBkHYBKtlQruX7jq/IVeA8Q6Ft
3KpHVwdfXaUBynbdq0HveBkXxB3cyTPMlCwyU6r0ZFGw626bqG1VRZCS+lHrGdYl
CYviII3+Qt7mUJlANa4Il//ygIR8wS+4C/wYT0pMMEI3FjNbveHO2bxIeSd/V8qo
1z1b13T1m6xUgEuSoRLQPb3YT/DRvsKRYLPA1MyIJuRG+xlCg+FoOYAddUmQ8kZq
saf1jJF/L5wyU7DFAxLIdJaPpBQc0dUqmzkc0cSLotft/qRYV2eSc/xTj6Zn8gst
LWpVoX+NKHlNQeBsUf1DLesjt+DkbJzXJCkJ7mGMK3wBJsroSeBIOCnNvuFOQQX5
D3Ct6LpvziVSy1hWZkZb5ccQOv2eJ4xH87wg/mfPq001jfOnL7ST3hpiDP8U0fBn
6OaCTyJFb8fCm738bXVD7BCppuB/CN/4fwf6/dE5o7I/waEQ4x65YvtgXN4pFhex
yIvPWyGOcM0ugu2U2XxGiT4teUlhInJ75OAM99eWQIB0KXRUXVHE1wiWPG5MrK8n
KlSdl8t1Qv188uw01N09Y0AtwDxtH78PkWan296kBqkKfEMott/+5NcfB1igPeoq
xr8IW8mQu1WrlWqdFQssaMVn00p1fmQMCQtmkiqP6gDQ+9bchM5q5cqyfxQnBS5j
qHf+0/TM9TDmoZHeth2BkFTkU056DcXYKJdE8kx6AICr58YijAQEdQrQ0f0tcM1v
+JHt3zFzobZY9JkOhk++wCoxHFwWjWiK4x3FM4OXXT3CJsGphnV2qnEeKnWWgE0H
u3iFt5IgcfMEA5VQafoYkIvZYEhRwqegW1rcrIPLXAXeYmGnvIX/JWdzLpU9ztZB
PyDSigApogEtNzBcbx7B8NLrEJeQ9d7GqU6He4NWiR1pUeINg0J+EZp3zLg9K+AQ
XgQT9rmTRK1ywXWtRHx5up7UUfNIr5wQCqUTsqMl7TQd5M2ipWCEmUBvXzFQu4bO
pG8lPdF5QFZN2hq2aEhnJtS9cAMMXXCmIygLE4yuO1bacwBpVeHULjSVbQJ+QoKJ
AGM700N164DikdHDZKySvuexXRJJJzEZSbJK3w8udibSfqrz2MSSkt4nshpJ60XO
pEdZYAYd4k3KZJr9jLv2sEllNaQlMR62K4fuyFaogGXj9KPBlXHBxdS2bRmPpixQ
dq7qxOldRnDVZoonrsO47VGxaaePTUPpjzfjlQtVLwDwBrqAsOrZLz+XSDfCsVHm
GqATpb3jqdB3rg8/KcZjV2YkYo7fvdnRAw9XGgaQCnsKfsgfOjjtr4qp3nX8sk4/
WeL1P2HRazKeYByfjORWuAthrRWGIl2qX4x/JM98XXt27FwcKmY4rcbcthq7+zPd
znhTVQy7CmYhxdfs46fz3znKfIPC8x+ur5vkB5rfFmyVEyYsDo4Qbd3MDZTE7CdE
O1X+A9kWJYE93Bbwz9u5sd2O/YPk0dap45mplK+0NrVxmoBtJbzpIpAJeSvy4rUh
217m4h/9XOBZ1bAwKsofb0WVpDni1n73KOa0e4hDgIHJw5ewGN8O+ICfKLR+YX2o
jQ90rIV9b7xyXl0WLLGpH3QneRGRa0I5LK0gvMz+xk6V1/nBxu2jbsq6SYS7kJp/
Ebvy4LTSPt5hXJ5QgIiuVvasN4yKdtMLB5tww+e5a25Ww0VtEkGZ2Im6z5R6aKzq
dr/cZXkVu+3D+MB87eMWJ707vsDYS0EnUqARatr+VmnQqzk6mpo2O73lUcTI6KMz
`protect END_PROTECTED
