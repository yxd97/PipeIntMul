`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1NH5ytvk9bmxdLFlkgLKk+jfsWNd21ZE/jlwaX4D/HenR4cAzphgpM5WDmTHVvcj
RFe5jBJyTujyHlDDMIENerhFNaqw5JSGogukUv2dS9vKJlO8OwGtVHJDrIMELKnp
igjF5dhGvA6l+43BktCCiELNuKX5PghWX2RfBdvwSOq/3D6mpEKDRLN9MulfOS3N
WkViwlrIEEzsy4G8+qIGvQ2CC5I0k+HJeSKGRRHqC+Vm0xLrzG+5mMjlO9cXmYv5
xmmZNHTMmQULDU8r6AFHWpJU/UG2HvfqewZugBVJT5YVkEd3bhlmlZHSSGtXCeBt
94/6WVoGCXuOysokb+cGCP+9TZsUlSyexZgsXg7VM0zycvO+83iTqa/1lbrdUikE
3qHnh+/xbxxvuoc8aL0mapKSEmxIGAMSxclqYdB/1qcsHYtMEhqdwO9ZioF96TQr
TyuCHuAbdMgXoGOCbhFvVPOStBEnotNG/njG8C+MnjNt1iJ9sL8TupTqpP6ALTA7
1Dn3GSUKtj9ZaMKowXfCvg4uCu23CKT3/kffOyvibbMC+gKuQ2n1RxdcgUMsmpRM
xi4jrlIkk7TZ2RIzki1bDbtMTsIMEwCjxLiusu5Y98ajLeKCHSYaVcYU8+s3VFYC
XVns3IEGHTQ7DGOcITN5nnGWiiwOfYiNqXayDWtUM/NnQHThF6EEu9uVSxFB2hfQ
opIS1SMP2xon3mlMT51F2A==
`protect END_PROTECTED
