`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xwogpXmlInUQ9HsHlydAlb8/LttlvFY8YB67jy2KIQRkxjaBhNmP9TabtVh43ZzJ
EPcvqLJSAJaCTpLt3Fe6lkzFurU1/nEDt+1Dilops0zWit3Ahn6pMhQaIE5u7bYT
wOEz2fYPp3bpebfq1w4ECb8m4IzARkUHgliJG3IxETJj8L4YrPf2Am8Tfk5+kZcu
J1zqKooeD/cxvn6iPex4vpPNZLdU/EF1hqK5LP4ntbrajeGRf0Q2B9KW9GlPFGJG
CS9i06T69dVEBKdKzMXhR95rFZfiHxv6PrxxWpo/j8o=
`protect END_PROTECTED
