`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rUPoBAbLEw//oT2P7lCA8QjJ/6V5WvQmASNy1XVTpUdkGZ6osERk8r0yDESI9gdU
8QpWMk8Y5bn3RmzaQhw9XSpWtthN90eMTyT/YFIviqc0VlwSsN1bg4bgR+jpYWFE
9NJF1rqdTCYJ7NMFYoVZZY8ncGomw/3qTQtOwblo1xbLNkkogAAKNP0k/Yu4MlnD
xzTxtHXU9q2VAjuOm3FWCwd2gIxm61VHp7rwudRtfqGGdhYLD1sWr1/G+t8CBoz/
5IasmLxllihFO93ajBqUr9YclByMtCAr9CoXJ8HHskuEl3f4VSV4AuaHx4fJJ0Im
3fPyfo0MZibjw/0uyroBxRNumRT1mVxHHqvECZhYBeeVuXYf/YKmxGMDlFEGUvyF
YBtcMJeXnCD7r1uzxaaleNatAGkiWdy1nWPkHlnG9C9SuulYzUjCZLY2//qlPoJw
puG6gvz6mZgvulM7koDFEOPrW7packKZu2iqHvYHRPks6OePXivWH6iOehb+qotY
W3izFypgXJZy6sV2abXStomqCYNSCQM86n6aTN/FgMF/CwzlIgG/BZf0dA4iFJfU
38BSk+O0hpLIoz5+MpPZSw==
`protect END_PROTECTED
