`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hankjC8OWaFslh3kjotIKaTU4wdXMaF4Fy5xPGBTl0RWjhjdHcAUP7CKrEG3d2X
j3R2Wptq6G+xAaHjkNApz18Zn2gq+gLp2uv9qv84BIZJ+69GK0wFXfTqMH3z3FYW
PATlYIgawap87zppLcM8nLzriCkcf9yKlXiBU5KjKkFkHqSFCvgMBYqJa/iQXfAf
h24oahmzVGllqN9w5cfXv2EZy6nLwmNdDLVe79x2kE0teT4n40g96fp59/viayP+
yHk6eci2yakhWLceCu8aZAp7WAgy/5LxrtJ+QmsrknyMaheh1zSlZMqxKea6lTBv
p+pQReQPG7riuvXIM5XyT9BoxAILZBygdKNWVra9ZxOywClXvdMyDWK+cgKs4fD4
ZATTLBep5zRqwmmlqr/s0aiyJalfU77yLavxzi5BWpuCiGENd2MCceiBrRBr25p5
EQz/4JoQYDh39b69PgCPlXvhjruHTH5oZ7AjqPbCFdSfoEtsqxEZ2MWXydAxXhiQ
8aNsQkZlF7RIygBtd2UnmjicdSea2iYxKZoJDXFvkY1wlQzOh2ymnmoXcniPHqz0
c4cNLwT5Sd3AuHhYn4cXi9H7EyK1Qhn62GEo/gqNwy4UrxaL6GzCmFJ/W3TkHg65
G7wzGiS/lqZ07aFtcsnPujYevjIIYw09tB9tibdS2RybKuCCommqr6kRVG9AIEMH
DXLshpar/DonPr3QURa8hIU6ZpST0PIi5Gcy/oLk4sXmH3VHMAjDCp+dGmlKtAvo
7SmI86h0cgnlGY+qOyV2FZ41bP0gHCtY4m4iJLrE4pegipO1IaiJIpYMIQWGI4zz
1LzdafOucK/oJVGmK+2vWkHq0+X8DXpjVzT40HhZQ/ULt0ul92tJVCW8nonNFX2n
6yW8MHiXS0qxZHhDjzTKNxz/TJYtBTDIwHHC0je9SH/j9nIn0ePGBm5vah+06IN2
HLVjDLGWnnexgGrFhj+BFcV9SWqacRlmvXNDG7y7eZ6Zonhi3aKKVDc0mNTxXoyY
7eEGFg5nTRvz8bQbMk/F/RffxRHKJXqPfskgCbrJLniCmeiRHS/SzihactpkrDbL
`protect END_PROTECTED
