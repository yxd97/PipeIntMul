`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDZBDMSR467vTMq4viLF+GqQRWuo9WT5vhSvMcDLGj4l6+JuOMKU4RliHN60mTJ3
oFhvzSogmi76HXdcZCaQkb7lb80f6TeARIyRKQ5p3gidNNPI1CTcyQ9REb0w0CD5
bGYtUIfyn2I8UN399yCl6n1RPPsdQRtLPndzvPcIf1OgB8UYceIBPa0vqOZjkk+u
vTyOI8TnMVoBEQJz9yCXl6ICtVsvowoC7uaIxxCY3g9p/E8exMq0rrrMZNeVCmzs
59lfpfFYKo2UgOxv+Nd7ZPrqIk+nJ21ylF3BC5vjFtv2YQrezi60ICGdiQ+1o1zK
2rNtnGcFnJf46NgAy4/gQUnzS29SLzKgDcHcljJueHzhfYmLzebyFYmGj0pPdDa7
zDcQ0N/sXNU38tiF7WSVeA==
`protect END_PROTECTED
