`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hGiRMExaMkLuBy/0A0md1UMcNrWpg4eovR5BDJJApkQL488fiIUSOGZtMb8zxU48
FYQrZCD2hfzlx3jiInB3t3pcCicEDhCFZcLNZBmxSFPUTMxlcS2MzG5ApM4zxSOh
5IfAcPnWJt++z8Bq3ZcCsa6GvrP0PB1qrVispJJttYC2Um64yrCeLuA9ieXBRE7I
prgwgiV9VM+feesGrLPPb7DOOboO5gs78lGr/QEysvU8F4ShpvEh9SBEYqw3TZ78
FIz/QG2LrQkLMUYiBGqQPpLRz1Ji6jcBMbJ0McIs1/5vWLvlabzWCsTpQuMkeFGX
lFFMekPZGzyHUCuB6F9jGlsaZrEeQnbA5TR0HRWF0sOMII5f9vzPV+NeZAZjc/rc
WfDeIulr5+H9MYxqCa85IlX50eh0gT/kWd4FkBTaVGwIYYZhSZynYNhRtH+/dl7y
5gY61FdFsbTA0B2xlXiKTsAHhoWTeYkpN5w/o54fTxoG5j13PFMdA5cbVS1Zv4zK
`protect END_PROTECTED
