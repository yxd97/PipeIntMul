`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvyVnbjaLkRVrgPzq/Vo386S61nD90rgsRm8i3746NTHsI5eDyUGk0nUAPPhm6cQ
GZV+/RTvW2ez5YwiQDnhHBddh9VBImQAbk/fDl3++THBddwpug0BjRldJIk3vLf9
gMhFQUEIxA5eJvk9mciXbRWJy6et1PExwW/fiyImhrPI1n+nPNzZBOpvIhcwMbk5
25EKW6ri1INiLr7qzGXU8SU1C5zbiXB1sjDwvru8GLBKHhttch1X48PLUHvk5h6u
y3wARrTQxTRA4uNoDJsXiDgALU8rW90wfb/eqJyaRqLbiurX2U0xn/Z4zr37J0Rr
Z8M/lFIdfAUZrK0tTmOXIrs68CBb/dx3s1793imo6zCwA+KIlAx8Rq3RY8Jmjzsn
cO2cqNbsvkc2U45KBw8dAfgnxr9ZD9G9ehkaEfAjQIeIuq7KZtpTEVMR2EHdbv9r
Jv9BZ5HL/zMRjAIIz+roydHlnWtrv6e3Wy+FIcCI9cYfQe08mS5CucVCkX695lej
9DMemhJFMe28luv43xwisHAnk2/987rASu+Bc+4+TOf5s9dFxKTQF9/7xwG0wSNI
9n3CV23BCAzSzPR6jTXic7TIaFmmPrgrYfJNrwbXaqCf5lFdzQSNA/YUFuIGAEOG
UrFMfwkyvNkz1JtuDsxHb8WJl9BtG6Uev9JqjgldQ1ha4aR30ZTPS64g6rKSKpwD
44KlywIimBBdOlAq/wqeZwx5X957SUDryrMFdIZbr6N3myMqunV49mmRaaFPjwEm
z9RMPjcX4qcs+i3iD/9+CDScXWHy/UTlbZ6Tj9OunC9zKDijifYT2N9VgP405fDq
8bU7ZvTG3tp5fZ+dgt84dtyUmr6OBxhU6LOgvDQAQKWCOIwctE7fDQyS1or55PDB
`protect END_PROTECTED
