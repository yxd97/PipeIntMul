`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7bob5eEox41gIADt5GAjJ8zNA6EWG0FnNsWB1DIsA0S0KinSJFxGQgmhHvW8pw5z
Rzs0hW+xPiRX0Uqlu/duyw+EVop5Cis3n4xQAW8Cr2NAHa0k67ISXWMHn+aZFTQZ
uD3120tXnL+4LqgirbGkUdmDT8qTKOnpWBPJcgyZofZIF2Mofggzd/sbc34dDfBf
+BkfCVoeCPXb9GEnwJVIX7YFiqrK5IeZrg60iLp1e90Z684INsVfBZCmyaXqHuZJ
RnZT3A0pBoj1rNrLF1zcEFIvtt9+BHzZ4b4aqvdWlmN0v2ZjWURlgzuMAfAcaTxr
uDaybtqayhLS9l0lbL8XDn9SpBFweSifF3TPrGwSccpEjM7bQDgdSBuVK03EsDIW
qSLYpRKETypW6bLmrE21KBpAqo/gQPfBhbGVrTrsj1cQEay9bv8I78Fsx8XLT+Au
0cOeRtkKzfGuctsoS7kHrboKfqREwMpqemq8SVz/YZ8fTPmXf2GcTfogoSa+cFj+
PlEVpAYL6CFdMT675BawuUeW7FsduqpD+zb78/2UXQQUqb7c/a1iT93hMjMni7+w
K6yrrVtb9w0ZoefebNtLWsVrwelHXer/nni4NI00PI/nj1RayFxI52Z7IHb9c2CL
arQLZLniDTmKxYDN33wxnBfGMpa0uZTu9u0EPUBAwVsf8siFKYvE7adBV1XE+KM9
qG9i49KPjB1W1jKiG7d6m6GrII0VT8xLuA60+ld76CE=
`protect END_PROTECTED
