`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TTk6VVuVpqaBpAx7mi0zIbtqlj+PXr7Ix2qxlYS6iTeIwZYVfRpKfVLQiY7SokPK
2XDgSgCj2y55lsiRoHrTxCm5UlL05us6/7by/xBVUYVg+KXekDKUb8la5Ma/Rdc/
SNIrPuTqVDr8Qi2GGdZ688D2Uy+fPWg56X/VGc/qTX2++CfxfW0MUBxP0fLB2WfT
BMXOnrC3E/7zph1tgCJnqRZksGu6nx63CmdcYPIO/dzS2wf3ZoZQlqTPmmEoQJfB
XhBZ8QDl/f4j3t6CFFoGC3XXkbghCv6kiNhRuauxmQJ8dBEi8HYDzICnqDq2q161
TTJX00KPDyoNzi2p68BbV7/6petMsV4VgmbbyoWQ8ydfedEnspsUqHyZlFB83s0l
QokGhlP8wspBSxs0MhWOLK7Y592BNHpJnHNePuOGp5rjw4InBdJTyTq0iPyVKvZ/
O86liOs0N8BXAtEPoZYR8B/RjqCn90xj8cvKFnDHjq7G8pkDRez7SMUrhXjVuteS
fhrwveOSXWYNIKgoAUsQvyHDo8nfKYoWm45eW8s891Mb08pT/EMVtkctkiarAQlL
RQlEhAa3tWWDnoY+4VLZmTEgvMmot7Q5fq8xogg1loaajTNx9rNANKROR+hGnr78
Ov6eS4JJytVSQ3cjM/3drEVg3H3nuitBXzr3XQNpHXAbiJU8utUojCPTchsOG7oV
bJKrvulmEvVuF4xCgGHoYFgTEZyyzoiaI8T108wIh+WEhs9MOJpSLiFIGe4C0jdM
msAJ0L7DJ4l13psl29GpCQ==
`protect END_PROTECTED
