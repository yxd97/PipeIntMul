`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZwugyoD/D9OKBcFTkMM7Ls9LPalqEHObbEYMRg1OrXrssqksLEEesmK3qRkEpVR
1lSJhBavfZB3feLJM7bLrKZts/yMyN9/kc9aojh8kqPeAIFl3sxSACvQI56C0QPn
1L0lmC9UsYNUKe+Ee6RTR/nPmg5uGX4RQIx2UQEFMLnni/kaQHpOBWF6BTvn/LRA
UCrW78G9V2HYJIH5Gx3f+aIbAXb3nd3Xn4N5oQI/T4qb04WeoYJfA9ze1JxsjysU
DuDcDAbAeCAgwtILPl4XTEXzBIXec9ugg4nElKtcQ/1lEBNAODAFaeJqxMnUVLio
jRlhTmhtu58UdDRpdbnv/0sfrbbBZKJcHpCkCa9ZaGNVRJUxou56kbreTByVld8A
MZlh67GTDFbZzJvQBYuk0w==
`protect END_PROTECTED
