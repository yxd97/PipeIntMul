`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSrma71lXq6EAhQ7kuVtI/T/75CvHwqqFIcgq4oupDmdaI7ET0BlaUn/CxnF8+M8
Ey/N82VHhbus8fZcU4EK20FHRP+nwajogtgamJpywVAPg4lqksFB2RfVGBbuKHR1
Zx1YdlcDtOyvzEXheUBYfYY3Xw0fPKYLmgql9PuhOv5zd1tIPK7/mZbq7HFQrReB
S0i1oJwNrL9JfrZjurkH4b0gKsQmO5RzNIFWN3WsUn30gB0Yd2LPq3hyOXnc1HNi
ltbPw0S9SMKyJLf9KsPeDRgJf+MT7dRYMiXzXgJwfmuREa3Wac0W4ZY9XFeTL/gs
rBq4zl2dJXeN2OMcK+o6h5D9Zn2B9w8EUKfJCS5omEPlCjCHpoixSMDmdD7WmXU9
eLw5s8yEg2NUgonyRH3fhf93Heq5H/gFZNwWs2YBt/2Mx2FUPqzIQabatJB6oARU
vteascfXtbPjgnnJMvv3n9Nkh+qsCqq/7f5yoyosgYckMil0Q4BcU5dVbLjh8mId
4GL0Ib6r1XTniL3pJnOQPP6MdM6CNdzy9kUedvTT/jeGovkT1VeNUEPYp9AG9ZsW
yq2kF6aRsINW9a56DHHhCgEBrESzHEdq4QkqPaaBZj2GFfnhdBQrytZ1pPxNjymc
UFpxRnVUhfh7+C86NYo2O4Z51tvrQn7xLQWI45PjyiHg1KsF79xfrYcmQtfNQF4y
Fu/OkOp6/Xb2vY2obLQxgp+UxvRTi3qHTWZbFI5wCLta9m5uy5QZ5FPsiyJl+uis
sCYXBYX4F0tINWAHOUi35Q==
`protect END_PROTECTED
