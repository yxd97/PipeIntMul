`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VziFXUtCpuExxGZ4nxqOzMytPrQko50cy76GdxEn3uZ9xAP25oQZY6KQfJZEc6kG
VOMqahZbvyjMg47HmXgRlkJroOyCL1P3nPKXZD+vmXQvVbbcyuGpp1+bh5WDRPkM
ZT4tDX/fsMwllFm5Qp5GESlleCncX7g7w1U9Vyr5b15S9BzNeXNhlRl3H+tOl1pI
V9yBm07IHS2KKojMOq9gGWiM3Hv2z6+uG5VnU5/9Rb0Ho/wX8yAjy0PWJX53MFeH
643tLC3ffKALTE6aI/9dKnrw3kGZa1Om58Rf2R4bUMK3uOjKPeWIdPeS2i1AXv1w
lo7FijDuThJQqyhMZFro7kqCe2lr3yEtEQw3M4nLgemgAK/TPuJFpIk1B6zspk/I
pCrM+RHVjdDpQce/RS4S91HeyfI9vXJQWggAls4sa5PaiTLUpocFA7gTNfuukulN
nrvhAJDaLyYvMS/Pb+/wqmBBqXWqasnzd/HZxOT+xi4QtIKZ89sjgvYbWQuqrnzn
zzYoy4s7I4GsQeRNZMmcHe12v5Y16luxJbmJkyRlMSN48TfGUV3glSPDMCPjQy9L
dHubTu02QyPHJfD2vFTKysibw4lahh5B0sKsgOo4yrfYQrHGTyIGU11bA3ZsJV9y
CZ7k4aG+X7KHqkVo5KszRQ==
`protect END_PROTECTED
