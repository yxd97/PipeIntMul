`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BHOe0MCwn7TBhtsVVaPmK1SfKq6LkzOFPQtbgN2+08KD6SH30TUKGzoHMxbOLA29
1EAVebBffsa/fYyO0j1pfCWUBaq8/rYrR6i3fciQz2JH4JxYRb/DYu8i0/prIpnI
UiwgjKsuHdmsoVqT4CBzPoE1vimQdlBRPw3LqUjWlXjx1AlQM0RnGfKVo4eR9n6r
ksPWod7DBe9syvFq62i6+RBWdxOvyPEqXGtCGRuxdJl/942lUSMlErr43nR90X9m
8oB5aKUrgDvvEqBZtHnk5+ln9lxOmFDxT4VNBkMohm5fF5nQZhk29oXkh/N9C6SB
i30USJI24zrKeFqoFezrRQ==
`protect END_PROTECTED
