`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJhYaPcH6fcWy0dJN/Z/qh5CRAadkAl8z+k09EH5wzw2vrRoyU+IHEcYfIk6yS1L
0dDWQSeDRxJccZy3nf4Hdw5vwz5gey+KhS6X/h+yXTpJXqtYwsHTvH4+i97+3GRk
yEJFTjraoRsbXaDpO9n3fFCIiAk8VzBGt+nAY7p7J6HpFhZ5f0WIWzJQ/hcgya1N
r7ZWsdHmBWaEFzBkKo+0QDVUA1wV/upjWzdiNPRyYtZ9iOiJpPhjuIo7Q2DW0T9W
DyAZrUR8JbLk6ilTb3Nh5MIC9WivIOUVaa7tpJ/O14hCXBeTsioNr5sVDUq5+VqX
W4btFoERRvQhNbvk/s9Nup/RigXz5uCoTykMRXVUtx3I8kF1zuMfGlzGJ+4sFpxL
AXwlk4itL2jUdh4qJgNofeRgK4zfxU3X5SUpcIuaikm5eYWej9tBcSvLyrsWO/9M
CgSLMSU9jeiP4wCMB9AN2AGeVNjB+VyTcOvFLujKchztqxm8ltAsLMHyFJBrA8Sk
020NObyiGgLbr6IUeX/tgHU6WhSKtVrx38O9fmIawBMIwn4Bp7sKBzv6gdP7R7Ho
fl216a6x4d1eUBHmhvsCb0Bevd/Lexhx6EZ8VfVdWhWeVDVV/GhzTBc8FHlH4o9N
7lHHgnC5qRjFyPjYZv1e9PI6Lfz11WXJQYzvMWW/0SG9+3njgmR+2+zpANyzyZ5r
ocJJpA/k6U0uCumUr9lZmxUufVORhHyg9mkakX77E/8/655T1W3cr6GKdZl2mitv
pxlb3OVbZUhIJ46Jk2xeW3Qux2/QsOmfCPc7Pekxk2jEQpHogd8vlSHIEdicRf0j
FdVlqk/zOtba4HYMnYLqry05QsuR3kkhDa7+5l93lVGoTJvl+ZYf/ljPqDULAdmZ
p9IDDwuP35VaqNAE/XhEiwATCPJdbCoe8won9CAt2T9aTZmbAVUMT1U/HQU+PNQx
548hVvbbFnuXJNuuo7kIpv1uJveniM7+DMxfbZWevCo5CiB4kf15HvStmg4POeT6
a//lKW/KUKJH0Jr8LqT5aj4DxbSyArqDfKYUq4Jl7ujFNH8usrBJ0B9s4mZqcd2x
DRzfQtGX1QPAieuK6NaNo/JhnWF4kcwRlP27ahr67qnfIM+tMrOOuhvQ6L2AhQZt
xbbgr34+V1AbtiXS5uLOvYsln2wX25OI6C8PAz3btlMwNoNloMyGDquUeo+3KIrN
BJYH51DC+KIIuOM9SRvzvyzL9CBAQITQBBMyDE2C5ILrImWpPbenqC0Ej7nxOUp+
1xkaLhDtkQLoAXo/6Aggmh/6CbACs0lNJ4CPcQnEKlZgAJ+vr9WXC3Hi6U1vrdbO
do+Z3mAH+ZqsY5yeyPCVUTUYTNvwpmG4TPUrnWur9VyKzPHb9gNrGqVsFaRLrw0P
pJmrCob/0sQdRLk+wG0gdMb2GGGTENXemBmyqWL26OgVHlnrPgWic3Ogf0JPqrOE
QlBfnm3JK8L8A94yBT4lGxnZvxhpETz1f9HiyqkLj0ZmkhBL7xEo5sH+G89Tivli
`protect END_PROTECTED
