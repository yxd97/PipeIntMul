`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T75qu08t7lhXGSY+Pc/Efq6P75qvr5mhg+Wb9X8PVppRIt7P+yYLvdDgyTWwUNo7
/EqzLSwCPTXr3iTgJ9IXfChCEphfXnrP/2NZ9APhLKXwzao8TPQVzKloJ2m4aZu0
6dxgWc3czvC/B9qxMYUrmgZs8K7/5RZFvjRaY7A9YelLWaKr7LxjwpYpS5WFZDXi
F3ib65yyICTimuETUWFBcCsoH8UahZx/l/q/U8QOyYbjXsW9zZ+npHRTJxSCaWix
rd/ewPaGan3EkVxwhAOhg7FmrzJn88dFGHxnf/J7omPONlov7WhEU19kXtqvuxGH
Y2+yv3C31TvTSsC/qYjv4Q==
`protect END_PROTECTED
