`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vhj6xZrsM4eq7mGhHijTqt+jFpVYdBmfmw/XZOMXIH7A7aNlohGrS9jEgRy54Bn5
EI3yW2P/gxTJviU7MycGmiuznJeEtcOZXM5kpXXJzg7UlGaYpvMZJun7DdCg6xxc
f81rtmWFLDlNhkTLwAVrhWbWp662I11geRWolhx1sCFgSVLqyeYBISxdhiBUO8PF
p42hQD4142iy2rBuP8/a9HEQrWxwT5bgVirYZ0uAXTt/m4DAivH6NiFDWt7GGSLP
5Qnph27n7mGID7cDU0qs5w==
`protect END_PROTECTED
