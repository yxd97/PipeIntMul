`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aLZvHjb2Wa+Z4eHYhNypztLkbwwYudKA06zUyPzzOrZf2RT1vZqtFXoHZbXAoaA8
e1xa/qb1SA0QjQ21qlD7jBNfk12fCGoNZy5MF5Yutm6PtXYjtOEUbcjFcMP66dE3
iiThpschEf94z0309y8Ztpea9od8ORjdLm7+l23vyO0MbmqA+FhZTAZ+thm5Ni2Y
ly60SNDV4z/FWo0LJgWzy/OVZqUrZFFV8KArMecHg0WxOgWJ5JRXTlKRyenF0/ar
F4pC8Cys4yHQYkuP3tGRfU2CXNubHnRVtrCGRAQ7xFlVMar/MUi9jXtXdbxEks0o
Hw3DrdUVuvSHUDJJyImsUQ==
`protect END_PROTECTED
