`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bucWZvQclNc6+kP5xP2r1LLm7k+xpYOOu+PnhRRAF1YmDgwZ1nihIsESPfcvI+F
lVMHfjnIaN60BuXNRg6Vy7MK4aCySC+1nACgJyhj+HDlacO7kLbQWqT5tOt1MdTN
kTQ2NahlQNtQdZaYo0rKmGX7i0zNtcAVfdCpsbbphKCWieWYBqjBP/2m8EIQzTyL
IOS+j0a44fowBztFZJrioTKmjyF899jmY5i5/wPHsBd3EjW0srxOHZcPzh7cWXSI
jKFZbJC/cFv87qkVbaw/xrw1mSjZtRZMmvsMjzUSsKJGL4zZyakGJic59JkSkTyc
vHPht1c3qMw4qmH1miVRFH+DokpVy8M4pX0iqCxDAoqud8hQsl4TBIuhswo47Prw
rGH+AOZblFhvc8JfbTwjdm4uZsR7mY7uY8zlgqbrDWrUBEAjnPJyBxTcoORa4KPo
sLQgWbF68BCwOv5CaLEv5tDppN3isqtzGISS9+6vYtzsJWf7whfwD0fjg5SxS77Y
/BKcfJfobGvvDM3f77zzYnMiiRkUsCmmXxAGfr/KYNOROqzCunlAG2FRT8U+dUsU
`protect END_PROTECTED
