`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wEMW9l/NSsPODz7HT2qUlZ+HlvjqvprKofKwxp1kNfXQCgzbq6Tu53k6njwGAAN1
O2Vw3R37ft0elwblNWRIweZcQXh/eDBsNRelu4AR4wjRvfeTjzWn8MiyoRZ961dV
5UZZIHIM5gNqnB7Cow2VMuzOAuLWAeVn2dYGw+Hb19VHw1U2aGh93VKpZZZgaAvz
R9xV6vZZiwrkPS9xP0L6DAwiQ+MWwHLH5TQN48BX7qhagveqXCrsunjz9EdBxSZR
zbQnzcPSunt0Mxv7H9pM8kQMj41d0EzA4iLcGoYMVmeyfRyRHO5aQhPLMgcFEEy4
M+unzPMoTM1vJD8YBlubfUSa3hCkh/cMwVzKHEqaE2UYcPjobg7uwAGFWJbI/E+P
ZL1ua9bZ2u80GWeSRfDIoP4aEtpYXZfiOCiUbtF+WrQhGxgWRr51yUUFP4oUYGmX
nOBGdPglT77RGyAsDL6RzZ+zPqRzew4iyXQNZnwdj6rwFA+BmiM6WVTgoNNlOo5M
0OPTwTnLnkbrtlobxhvYfmq4JvxMjeO5LnvxDb55ooqYnT0yVoSivjXSKUzBNTWo
EkeMTkqsXSaPICml6x4Vg7hwojcPId5MznyuCdieIkQQMl/jrMQNq1xxafSuoJoE
0zaXeQUMcEx2efy2Zbd8A6i5CRSlIieNtR5TVrm+vUSI3CToKO+MsQN0I5oiaZVy
w2sHkoshgP12ESd+IZRKPd/NWNVZekHKH9hDsz8f7g0EY5NKr2qqqoPIXwFDHuLZ
K5Zz9FyklRoi4H9DeCDDoA8wNDji8y6hSW0gYLWC8T53845tPj/U0D683oVINdTO
iJKKeJoq8vtA6U9XnSltipl8ZZNAYteQsc+eDKP1khyN0YOA10fSxIoobPH/n/Ta
CJTrCOa0qKKhgUzIzAVPcGGrl7Vgyd3GUXhfSiE0+o6oluThk3lsYP7CmTdLKYO3
3rEe/Z44JbUApAqtQL/AcXnCtBAQzeZB/Tk2W962MO43LiuF91ZORCpk8Rrz5nZH
73/phPLh9qxovA0uv+Wi50PLvMONeDbSR1C2Z9AsqS96zwJxZbM+G0UhUK9lHOth
ydu5AXkfmrk2l76VPevNt4jviTJrFDLHm4yPK9oBHHEMI+j8rTZkx1b7PQKC75zb
z2AHIT87VAD/ml4eEc6Vxz+OAfooxotBx74DID+HDP+yIhxAPb1ZtBJ4Xov7mtrX
9zksLNWp6V6/AZAnQEqwaTNA8is2LZC/OqOG0miV844sjQ9wTuxRgTyQ3Hsjh4ry
7szVu81XcIKZLNxVxydhDpOAL8SWwiVxBnF2NHX6ARufPwlcEJfQFp2xvxMb2ksD
FPn68f2lOlGXu0kAagdAGWoIytJVajKX7QwhcIFh9XR4KKzRiNSPQb/OQTbFGbze
MvTf8gMN8f2oVLvY4Ef3ZNoB8OxQRhmoAjcRH8CIn7dZCWnuxFsqfRpIwCm10u5Q
waGEiNo2nI6RqfOqRLNElerNN1uBQDcmVrswSvvp5wjJRQ50/eaAyoz58aR2WGxr
zO02+VGaxyPrI04d4zkfANKyDuYUsipQiXHLuMbBCemvCf/AyMwXYcVIld/7trEy
oH0mXUybTRHULXapk0dEdLM8RD/NieqSShZ5OcaSxo06lv8tRd4anM1gpEktWkzO
zhViAG+ZCpWgPiTH4rS344Pq+01vLGi9ckaLz1C/1cRVcl6+vJtvE2OEiPV9euOv
uKheCAESAskw0sGyzvzp1oZtMOH1wfjyYo6Cz2BsaKyQ5UnAlh/NGe7o1uo3ERae
ubEW75xcQb4N0Iuj7TF2Am+pwjsYXgQ/UiexA+kQIR4O00xBiN+0/FjI40IGMcqb
A7ekGvmUBzXMWKPmBZduIqDgbZszP0Yr1/m09TzMGr17jekPw6Owf+LWQjxUmWXL
Ic3cTnvVW2Po9QdNjjGJAOUAt6c34TksUQHcEY70O9Yd1Uq2T3bDBsdZyT7WvbGv
RwOjSqN3eq+OMKB2wjJYtiw1GQIVEeMOUElg6jYCgPsQtKPFdQTI7B6Kid/Erhmk
8b77s0wTnZVTqtrfcsEkDQfr9+6zskBG9Uem1FkLupAFfKqGGls+l24vClG3rUxU
WltDQiXWVkmbZAWYjRthm0WuPGUWTsHhfDkO0Jv3oQtR/jlCuweRsiqb2C+bnuo7
PDpYluvVs1LN6OSI37sZ+YtNqYIRvjja3g58xFKROwf9GZ2wqPK0GLdTmZnfHW+o
POM1+VyWg45ukfw+9YaYnT2VQTfQvYBdXXy1R/ij/Aq1duoxgigYAQiU8fiKEiQN
tHkDAt/W8V7U6fHoCWBiCt7ScUm905PZnwDmC3v5mJCo4IQL6jKtOcKmIwfrD3sJ
5Os25on5bE4hm4geHXxe/M1eF886DljGQUisqfT1WkN8UB0fT9VOCY6ZO59OJaTh
OJu2yQw8yvansh74R6pfXUdExaeh1GdtmdNB3IPg3B8o22ChAtx8ASlhnnzN7HxL
+fiy+6fpM5NBbCs7rlZSesJmyHvLqxqGeR5skMEDL1//rSU6I/2Czy3s6YkEjc4+
PmABy3609c+KjdkQgvWnA4c67TD4hK0EJhpgNtiTz6psGTgaDKm5OTu6j9t1TH5q
tsVUuIwady1pD6rawbYoHVE2ViIBAVx47Kiwz54KN05PqvY3Am/TZrDARCDKAvDG
s/7Rx407UIFbUPIth6OJfSK+a9AExD7496cIxaShsS7IXL9Ep5DHI21kH9PHZV/8
xLOTAE+CFzwERtiQ+sOLGNM/5fItcEEh2tDrkt7p8AJvrRl/TBXdRD9ilB6FXnXw
GcvuxG9jEuQEjiB96zgfGg8px95yBBHqKuMkApQrxttCim6PqUZLj/mhv3Fy50N7
aNYesidahrsLSoL9X2s7QAYTXjlHGYrdKGKoA9Bu5/C6nkbCmoRHE05NU3gWREoT
scwWG/MDx7/zwGwdoa2IUQ+iVgmqVb5r54YpEprpldYlzb2+aEGick7C2N+95Sz/
qlL1EuNJ7z9FjTtvm4M2Zr7TsEf87fVK+jTkbLOUroEUoWvPGwmR2ktsc78MG7gu
yK94RsWhvs135oD8Dy/LdnuJLxtCk7VLAww67TwxLlM+8nOz8ZjtcV4QDOJGdKin
hdfrp7Z9oeErU51zTUlAvgEHOgkqS2SwW1svz+EmMSarcN1XI3y7ntzbw9yLZgIm
CZdgMceBp7GxIcLt94CXR4eoFgoTEBKhXit4T7VTEhRk3/Ial/unyRtgug93H1D/
y/uwP8xIvenbvZ3TVPT1y7WTmKNmqlm0mTKfgDN6k6sN1jbXeAMyMMWWorUkpQYW
Qh1qkbEheUpz4Ju69MvVrvmZtoavUWWhRxAXlUaZI0fWWcxMR0CS2y6OnjH2y6/v
rQYmlf+4a/Vc05WQjmCl0DOJuLdHdZb321Q7hM6IkUjyGTjxRDAZEvC4eTG+9n2b
bRHUYID9FMyE/PFVeRPW63zBr9hKXqXnzlbA/m3dzTFFjP2rMVWvQLewLzOmapD6
TdnAPX+IUpvFaQ36Isq/rbRpkNjofIBd0euAafQlRXPuUCvsprZyqMZyRll4JCmp
AvY/eoQhq9IjgcHiBAozj5Brp/lu95hn82yjcoPkH5N05vRL4Mh6rd5BaV/JdRbh
O/hfP6aojtWz2bs+6/2UqQbMz3nYUJEBaN1n5xyLuDsjXxxmJ5Ol0MjyZRJE72eM
ciN7HxKuFw+uoSq9E1MkMRexloVBem4Bt9HOzWM8wqhEH1RR1ZQ/ArWYmamADXuC
rkT8EqrmY3khjYX/4acI0xIrk128TEb1+E6qhpZTQh+okhOfZi1VhfXlgALJzcOz
18b6HF2flRyhcDid7jfKmah+TaHX9rOb5a1SUEx2M/RbzJ8gngqE8V/KMKXFU+vT
WKd1gc+4igZPwrG5Y30j2MJzNOjv1D4uJe+LLQoLs2DfeayPdH5tXzD+yOSGSVYW
iXr5NCdYi8yKo2Bj46cMq2mCUIlpKQngeFXUl5VN/gbl3E+YRPSo8xsiLFwNnztP
d2/0ECumJNFtYzvVxm2a4yI1dM7W3afXGg6bHWNDZLYnhcd6ZxKosIQ7kOuZspTm
OM9PWPcODjpNO+SICsik0XK9dMFhdC6Pz/6ta1xW78NhQCdZrB4oepLQn8eqjewF
MdGH+iDD5bJ0HWNmtd9/zSR1cumIc/pxAJ0KWAYauh5oHLy1QDd6PN2uWnNFajku
nM1t4b4qvn8ncbF2ok/C/VpILRrfLHd1TOWrCVG73F4WzyJEjxeadOvv+UuMWM+c
aArNJRV3YhcK6nash/56ItM+9/wIbQ4u9LkBxQ8ycvHxORaxLABG0aAsrmVTgUPq
pj8GRFgNW9GzImp5V7FQnVTwuC06FfBl6XUR0VynCcLdAq/DFoycNE/UHnWRue4M
AGOe6VI/cgywLfGYUg03azFt4rkD24urJu/aThpecm3yumNcmDjbjzog+pKib1zh
QA2lwvsQbhzUZNFAYewBKPN3shvB/TmX90Pgb0vZ7p3XATYl0wuLycEJQ1nlUdm1
Ueac9hSU+FhRRoeLSdZc1qv8uhW/zL1Fupv6RW/MBfdLSW3hlbn7wS94o9YA3idh
RcSfBK6hKYM590M6SpBtQxDYqnjl2mqF1IMXIBK51zK7GFRpGXgZaZBEKuGNeTcX
urWtuSIzSK1zeA0/a82a6H3VM+SmLxRCOrc95Q7MFCOZWEUKFY419ykZhzsInWxE
DJEAGIikyW7q3G+YNWAGaXyN564cdPzRGbn2sR8H+4WY4NwN/WS0UjDcrYj5f24S
//l9vv6P22k55GbXUT/E6OrwLwtIylICegx9qo8UWpFDTn3qdr2dgW2XYIs2Q4Fi
56ZEu6pl2pEfyjt8rcoQnd6bqkza0LIJS56FzE++69D00fH5mVM2M/68Ai3HbBnu
x27vGkz9ZCFYNvI+/zz/rfZJCOeFV+Ks3Sbm4XFYJNrj5HjtUAdXXHCf/y8/burW
pt9WO5V6bsf9H6bOiX5x2jhCxtNgdoLWosbgpQjtUGfO9ZTCgLVgmdAiNWjpbVwY
cBypl/tYmwGjFwbZYfQcSqjuj4uMSCTowW2U8+ZFoHOLQ1qo04GcTDcee9harkqw
7HKkmCiPRSE4/hcBhtOUiSzDneOQb0NX6hDlIAj1l6vMfdJpO3CNgCXvUq3o8QYd
Z5qPuUtIkEMe+iZVJ2GT7MQU83M0m0SCsFtw+krC33pJscz24It99Yvkc/Al2qJE
+fno7GTA3qWK5rtuSGidZ7WpxPO6SeZVPGIbKrq11jn/WpxEw5QQHHjl816cM0bG
4imSscEeiT4GNirC8sa9bIeJbwjEVHMZAkD9VsD1hMzV6sFtCD+oLZJwsV8Baz3E
pT5DdsxPqvkloMvVPye13nGDTSOwSXMYr73OOouZy18q1DPo5Q3EqtUX/H2Ej2v+
/goOi06foCNmpduIV7L7p7NOoetgm8+D34VbQ2h5P/ba2X3Dqa1v8IWmWxOl0rKX
u9v7Yabc5eCXjD/CtjU4TcIPH+gTcoet7uTwlSZZVorzYQprBywDCvlnHFXGNJPi
CrMfcajVw0fDBXERdkiha2CgqLxPkw44/NlHhMg0lbEJzije5BijjXMSAxYkmnA/
OWvSUXCNVq65dCIPJI8RS1UOW5qtL7B0lLR/UaavxdPByBGj9ScOzZhjCXMxtUbG
Ly4PqjvPRfe2LwtPqkQ8cevxCUpR0fQGScYr//aWhV5beVJzhb1oUnvU8ZOj82zp
y4gJHtOd8gmld1uql8y6IHVmirStTfdKNX8z9EfYdz9UxaVVKYKMAZzalJscmYMI
Dx/CFydewQNLUD6GURoTjUmkYz0UEMdEbcLMVRtlrc6u/OuLPBYVa5jPrqjrLeJe
JJV8wxIXXYKiEnz9v+1T0BzfrWW0GshOc8FxMYdfEhZEosd1ukFOc2Fq5sk7s51v
n9RSC7jxR1jdd/+dy+4jiHWfsFva5EAyvzGSkmC8u99uYBYn1FcKBM6palEJ+Qbs
HX2d5qPexMrci0cnQ/BAaoM50SugFXg8gHw/l/jYcS0aQuCQrWLMr/dJoz0mIV0T
HESGyTRRyqHoQxc6v+35DaVzOnC2GNtPY5JzOLIIqcmlromzL1qPckIAYHNXdfGm
2RElR9TEP2TKgD6eIP3FYsdg6QEQh/r0ABl2dQYlW/5fUyA9745Yo8Qymnzz7rLY
EpobH+igAgWbyFhD/ZQ9ZMW56BMPbVIYO9An1dmtxCpK5+BviyuJVtTO6W/o9eBk
1FoVw8j4r62ct54STatqfD/PbKH6K/bx+cj1VWuzMtDnnttWMXzFn7oazDvZTi7Z
vlzG6ysc1MIMKwL4NkMVhslBJiqkpxr3+ovLOVkF86lOIMicgMDvz+kDjES4GFRg
dOzEYA2xYnMr1V2SLyPSt1/N9hdcnPMijEDpJoRBvpim6DaWp/CtudA2Q2rjzgNz
uu1ogDSsjTbOOC/lM433mAFNlK6TKU0iOtjkQPPHKgsCSz7Wy2Lu3lfvjb1yiA8/
LnRMXlqVxA4pSvpbIVxir6+ZLBCA0bMad24Fbe4DHV6inATgacQ1Go3CDWe68TXe
VV5SM9t6g62q+1PztOcAAPeNLksHS6hqRgQDkjRsjUU2oTVSctb9VagVgA9bNsQl
l7U8UADeuK33mwu/oC0kWZXbA2Eco4dwZQ7ul/7oHBnwlvUEa/gIpDZ/Exysul7i
RXHM8HyhtAgPmmsk7AdgMQ+DBhZhdS6hoVtRLpUIHIyTTgRhEfbO/AYMzJDw5xj4
OFJjF6eAgs0zLs0Z/8iWJMKLNduLLvQFF+QrtknBVl7CsDXh4DjD3MaPFs+YTPj1
KOkZbQORQ4fLAE0O+MJ/F3vljvyac93e1fZ2RQD1179Bin04oqItlFyc2CqWlx5C
xFWuKIlKwA9ysK1KWsU+y/1WpTYQSnAX6CCT8NxTYXjU23U+USHvx8OhXDNwNa4U
ehFmWjLMmed2Xsp1ifXOISp8sTImSFq+F7zQgbj03nya+iMMbgL72tFUpDbx1MkO
OfyahEZiJ/nGnn5xR+5+MZRrk5jdOYS83aBT9yWxl/+Uy17tjL5D1FUa6WMglex8
/hamNDgB85ULKzOArxrRxUYXM54cmv9dzopijmkmfesGheJJAZmsODic0/LU38IA
AUoebYAOvAfXtqH5ElohlEulkLF1T9s3dvnYfe+lxuUgzf/Adv6ipUu6m4jescOT
EBLw0iJqdBT0Rh6GjU8j1m6Ddo09OHVgXhtsoZv1JT/HNeClM1mrC+SudWCbgDxV
VTTc4K8i5YBvjhtvNja/Fn5xbkb9bqQHmnuZFSERsm6e3dMzLPA91psLLoZu1X4+
z0/fjzCNqsO0uLN0gZj9VLmFxqR2Yg4eODvV48FSih+M5kXQDfnCH38dbcTb6uL8
gyNHB3gZesNWLqyVBUE41TsvrfpjJIEgFRRkZTGwnoes3/74jtB38Rboan0tc/yh
3Y7Vt93XlYf7pFe5IWbvK5GwRbzAMDNYh6CxnGyjv2xp85YhZDqcJ2UgMX8LOPai
7IgvuyzLvfRqjNgTIZZ6u6dpTHsTmha12wKvX75mO+pG6szJT+wAqp47VSP0SEyk
px96EMuUOSXGZQWKVdj7OfLpL/yLWfSkg9AblIYZTERHO4GPmggu/bE07NVlzj0a
ANWNisnCyJ/IbimFrj+gBawf9IQJAH71VuTA2fpMYIPotzBuXoU+TGnslmV0KFlf
xgkcYLZQ+HfolwbaZp6IPxNffLv8R4uv8lN/yFPBlvlV097jlEz519kKUhl7x+ce
Ns4nRWBSV/hbtbtKxXzOpoqCvaW0s2OkBybBJKhU/km7Zd+Jxe14iFAQWaSirjM9
HShFbMqEMUY20J5F5qms1yKcmXrrAIY8KOBvuY7SlrMqqMCeu8I+GvFThzZp4afQ
xxjJ0Y4MkFpLF4l8Xl6cIdhsYYaaS590IaTmzHY97aBEbHn3Z9LAPbBUrB4vDzrX
6kvV2ghur/Y3eFLuKjNpB3pv3M87Th8fbCoJGiDXvIaTIUYmezZCJP5DkcHwGepD
L+1IDMMpoyRFpltYZ131SDXj0FFLrOTFy7gbRyX1MczY6z2aUdbOt4ZNEyaFkMUL
209ddy39GgedDurpTlkv8+8k6f8kal+59r+UItoznf5K5qIzhEeNgDlXkGn14/84
6RvYBJAh4uiebHk6A31s8PZnBK8gcrwuiRcSvYO3whfiponkG4w/57n0yT7ruvtN
UNa41uvl/bOV1bVmO3i5y0Wvjo9djRo6BVYfRO3VF2wQXFNWnoVGNjddWyO82zHD
84Id29+cALNeUHS9puHTPrlsmxLR3YuMNOfnJkW3xHIRe5mUJFWZqVPo8QHh/lLx
W4grzKqJWThXSNvqXrueuJtsL1AZOSa3jBhpiLCaeHkpvJIVPN8ONMcLq/lVXt+S
PpFiHSyNTqgkjyFS8+qCIe6M7+uNMcEI/gv/j1rLWVjzqyuLvJzK5Jze/iRzFyBJ
K03Lva+8DBJ6UcCIAP9qrP4eCkskrTZtRu84Yy4eAsN0PKARV9Sj9GGx8mYaLNPN
u0vtdPjwwcw/FoTP3h4HF9TlZGugS5Z7N1cANlp3ae6pBLYJblnzHo3F6qWIs7Pq
07K9PKMYTy6KfJv6ZsySwTaMBcClWEaxvLMiSodQR7T57nIf1AEu64f8pTvBEisk
x2QMQzlE/vInoPqZWzrYPK9h1blz+iX+THuA/VHSndIUuCFu/EfMfsLQzEL+wDHv
O5tkO8taay6EL3OBZzeHuX1tCJQEfknmCheny5RSyOBU3BmAI8ifxQnZnGyIq+ha
YAOk6STNjNe+iZcOeohBpfe9TdyBf0RhStbfxK9oXCUyeHsYKrgdXa9UdP71dE7x
0rgf0XGALlgsKDO43lG3+t/XPyM5an1yPVdM5SCkdMYPl4WQHjF7ZDEI2MHS5IyW
5PI/wKfY1zs1uVIrJxbQTd/kYiLQLPZucbCe4OLQA3eIsbVVTS54xmgw0VTHgsUX
rkrU9gq3X92tyvAYgsx4DZffAyhXPczw80yl5pEcqLj09BCey+81eB7jUsYErF1i
Lwg/9M1MAzvnTZzCdnZdzNLVruQpdvPQ9cLpntkG7Ufji5TungyFj5lKqL6HM8AG
j9j4w/pRLhxkFs9NOxMkJFCJuYABVO8fkhX414pQDkuJEeZr8bEr5lgyg6DpEgl1
a61ia1SuSKJSfr+uQ3XJ+KFCN6p37bE+nwre7XUsXa65Xm2yjuAQIUfWHAMmElVA
akpiiXc3o3zUAE5zBYr+8d8ntmx7Z0CYSsU67X/PJCC00zHhtaJUfGMwj3Bkbbhr
/LM9+Mw6zcan3NHM1mjlZWDJdv27G7MRSVWleJ6XPNwyCLRoWReaOIajEM21tgEC
T4Jdpl+gjYRqyXVopOs6ArrqLaUZ9tHtwNQt3RG8WbtWzRihtF1/zJbg+lVliNqL
u+gszq1p0urpQYRXgq9wstgEmyLw7GTLmE/FQWQjJPFi/bDVjRBYZ1ehdom50wBk
vBi6IJRLHrSuMn/to6KogkIsqxSTlGMidQRAha0bY2s3TkR0Gw3SpwILYs1PqFZf
tLEZsCTaEvL+Kq7YeRs2LAzO6paS04ZojCrL1Ke/HP/cuZscLCbsDR5GRqlYY8en
HT+RWKbUhAsScqQELBdwEK8lhLIXQCDEfozkOuCo/m7SL2E/IERQ3dBFRqJqpucu
1hGfyM2xlMd27mLl9rNlf0YDKUuWR+apYLD2ddaRV5boXfPZtsj+b09+XbPcqxqW
EwXEdXz51UnCpYt7otIwtK3o6e/5IEP8fd5RCF19wd8dggQaVa6PKQFmbA2pKrE/
QWk1oJalLTh51c0xkBmM8wpKBC/0fDCpVKvc9kaeb3fmcCFmOG9ogipMz/pETcPs
R+P9NPV4yIGSb3miK2xt+/uK1Od/im2nHtc5YJ7k04oDsahGCeP9rdSJdPGAS+A4
w+cJF6V5riIZKFsn5JkULbPcYHFabyKe0vTdfN9quThfOxoCNi1I7HgMFN7Jfh91
7uI4i0D5pojaZL49lVcWxYLOlUoU2zwVOkARCnc4II1MywVjXfMKihUPaBFj31LH
UDWI7vfTa3WJ+yyWt5/yWyP9a0iH2jt3kX+kkuMw40HMhdvbGaaFSCKCo81Z6G8+
aD8LnqCzIhXCASzgZfH7eCyMuzH6/6MZwFJS3LFQLWAg9PL4wZhvYW24MSw18w65
1/GSFu438Mknj5a3v58ijVf8FsTwNRz6656s0tsKKEVao8dKeDsPPT7kazrEpUWD
tEVwMtFTlHSnbfdObT549PKNWuNze6ZXWJ19dEcZckg8lggL16KWdo8UelqPYHgV
jZ0iBIhcHOgHMCGQKd+VZZXn0GuiU1UxgHmSoAOR2QM/Tf9UvgZ5HOdA7L+Qesph
wv4IPv6Uh+BdUFebWMwxb5l2+Cuxb5/yM94zUPjlBv/d4/UzCLe+EIQaN75dSuKw
iUs8Su+fQuIVcdoeuLsCH1hGa8PXMwgRdJzobAoWrPtTAvL2ZbrL6IDEZEqc4pK2
ScFA9u8nRKQ5TNDRXpeM43My3VOyzgmGjBmO2lom0p0+z1bl0vQI3+9LusCY1cQJ
zdY84vAeawfv1QNXPb6YX/ip0/G9ZJErMKjiMUKOVHw34qTp3F0UrHTaSc9R5jLe
ZMiTYo4es8ZVQQbQggg1paLvVPd2FBgM0O1WJgm5ffRuOLhUJSbcxpKmJFlP/60E
XeoZg/ecS3jqB24wAD/CNwGt9ycWSg97c4TKUNijXtSziZTGRZFkg+yqR96m6nC2
DN4Oz6WGB7evtNBuDrCFspBcKXaLsknQTdMasEqNAvQfWOQSwDW8OFKG87pcW5yB
rTgWv4DVIonJyLTyH1cRGJzBc8kHC3VrNgxGXRA71iaEV10qJ/6wFTNuFKhw3spS
6IkaS51Gv/jZApgbOH8uvjMtbQ79BepFFIjOqT8Tg8qEpxwd33I96auHhWZqBE+K
csyhF/kdIHYjiH0YcEUTVCDbDBlh9wLuarZatOH22NYqH/P448JJvmltY+kl8NXr
86SXNqduQEkY+Cy2a/AI5m01qduNLR6Ryj4epTZ2MVix/0RKy8/wNnI9x/vjkayD
rEVs3z5Jpno2J51FPJrcvik2uf4hwM16jwo/aRtxn/CeaDC4VDwZ4jLZjxsKs3K2
poIoXsagdO/LXf2QmJ8yVDqWU4qvXGwNngJlIdB0hMEov/5g4H6M2TOJjb+3GO+O
SBxzU0iD4Z5met0znyKqlndpYuoQVYpd2MBJUfEvTPEPyRZAoIMC/YIFxOu7NLZu
Dq3sYfDYVQpal8py4BE6/MygbCfzXLzWNmrPJVcc3juo05MfX3MPHZgUXegY5DU/
mAOTwYmz+2aLOhBxSzIJiJN++y0aiYH5XTfxUw+P5oBtZYXNiic3f7CcdsZOO7nQ
LRKyBJIlZQt7ElMNhlvefJ9yhIq3JqNQF/IggzeAEysKpst9Fg8TW5RS9MY7FNxa
6izwwCh+bMkcpBZ5PWBXONVbimpy65Jc96/rp1W6N9n1Pn6gbwt9wCLIZ62jn1Bs
3OpecDfi3t4usZOyYf85xOG4I17xpPTEhfeW/2A6KeRkOCPb7FMlJK2XWdl+jsZ2
fx+Y3yHloJSmRXPJpiri7g+EpGnvAbnjs/3a0q26IVgTzR6hJzfHp2EsbIk1sDA+
6ShYUV49SXVt9NJVaitqum8OCh3IZOIMgVeorFKUdtO+qwJ9XdALbpFjyyhjxnX0
Xs4g5Kb/5I5NvZfq16dbdj2gpGIq1wKt94IDpbF7n7s4Ny538vTohHc68bFRm8MN
39R6d86NnACerjVGXQ7pliM5dM16T4tlFOand/D1o9lb7ID9nRapFHbrovz62/6j
7rqTzkbLIFrAweX7ePBSNiWIedcS+FyzfoimPIdK9H7Z/uU5i8fkc9q8Y3SVabcw
PSkRH8rqk6ho+LSIgiYDI+NL7LhkMBNKaOQGHrWZs1SQ0fkkWQH5+SkgFKzxJO4t
S9SnyS/R7SmvSreDdKkdZWaHjqN8GN2g9/Od3nH3RAonVoJG8N/+Q5foC7RrIwem
LlryfCVXfSDx4wraYHJPsjVGTmxrysXLhKtaH97N8mTXuxlYGoArwqlwPOLUiAj9
ufdrvaIkFy6WqwKK898f50OPrSGEQF2snE5OVHrLH2KLI6gfehbyiZBdpvgtVJsu
TL4L+ptkZScrDPg7D67lIQYNOA/iOw0CGGp01xfVg+pHTMHY5BCVrxMbu21mwJEN
owXPjf9b/nKAXkAerd6eaq7tCayqA37qh8jU7fP/P6WLtxhvAmKQOH3itm3w8KCO
jmhh5PT2zNu5RqJ20GrXn6I1F4zTQih8gWPWXakuOy6HJblnVw682k2NQfVSTIt2
gdTg5ZrxkLBV9eLZbNIVRyQKmt7fXPSdj5ACRvjCDZcvY4OrqmVykCQQP61a1Cck
FiNf5gP2XGakRvgVw2ZOqURu6HVniMEdKCrHHpPE69G1j94pKj50YALC8QiAIutj
IT4xBiMHlW/GqwfJGtINQe7tTsOFj49syAmp6Ba/gfacxXmx2+8pe78I05+CufqA
cn2xktXEK/xRsduz1TAWf6TpTpaioV6kuukO/WjOcPWH6LgBuSD6Ya7TvDo2ko0t
7WKtdgquZGtkY5Y5Eg9ZykrkHgb1BPsOBYeHZXw/TFhmmlEkSBAdDKPEjjg8Vk6L
2uiCGhH6MBGJTDTZJwj5msU2tlfqsJ2NPKZPcVpS2iw/pRPE9eT4B2ozg+li3a5d
lqdhRpgH6CqfApA9J8DURCLYxzijkUR4ZAN8IBfTgiT29gacfhtqLYdIvmk6vUYs
n6T+guKomIeM7FQ6Uk/VRjeEzwd8jKexvh2hZAwDT4bBGy+pAMpCT8ykNuqGpRxL
RDTCdS9AEb1nhFKgLe0yC9JTIDNBuMJ3tbFgh4A9y5SRldUL0Fz1eL1wPrgOKqCT
3vG9MmmoWWulceGI0hF7OK0zPClc1V0RxRX8K4ttmED5mPZ7W28fvB7zN7PND6T+
pv9r7gbUOUnjlASG71IsR0oN61dpy+3Xho6u2XLUDF0yaDmsbMKXP4/n1PFM+Pm3
uY4ab2ZMEXA5gbM+98AuDvHCSgG2y7bDAw6xsx6+vdtpV7FnvZkJRgbBP6zS4Mkh
Ov/+4AehkCuXtJn0PLAZMy+Sjf9T+BFPvJxnMmoFNBrNI4JwHBRI0WA5S76cKBTa
2hQumum6/N71B5mutWPYqdoD08bVlN0hfLWn5yelLawoXukgEeSlfy+OoYjyZGBW
V1f0ecUB66Ri4oCI0LuSPNqdKaXpiaDQos8SDpbYhOlxuAKttINsMRSoNNI0eo4E
fS8DJVdsBvnrQVnrFeig0fPic2SdXYoWp9yYMBsu+/QzGtGmr/d4Hj/NQNanWzV8
vXkkYvEZELTkL0ilEQUJJdDylRfYpjzZH6IxrHqcODssocxErGUNfhG+81treVuI
EhloMN3ACt0mqRZtSJfvOd+mNUb7OBFazG2ZyyvVEFr0l9B2WOm3tetTIlOWG2Wu
rj6ZpIqPcg5PLa+6cUzhoYAHT8UEQUaHpeeTjLQGdH/+Xvei43fyjsRRM17WeUc5
AI64diDD/9gL30FAuSLi7PB4KcFEsH0s6BW2K7OoVFV6aHxTgjqM/qPKVPu+XKUR
6ngOZDO7DGmsv6BhN6pPvLnPJ1FisSRhgJ77lMvbtHmptctigqyeYtaTtSDggwTC
kSRac1Q3N8ql1QI7JNb6r/gw1jruK0vOgPa9FgYLPfyMW4DhZmUMTDGN7fKn+B/V
ynMexSmFVjVc9hsZH0Wt9auosljxXS9xE1pHM72qy0J09pt4YGZ3he2jPet93iIB
Ez5ZfGWJOr0rMcT9FaB4cylCZ/JVo0xf/e6QQUEWElzj+G28lVNYnwNjse8GuE2D
gteCPGyJUY+QlD60X5e6MfREfX5yrIocn7/8Hg26nFq1veJlSjYghicYTgww25pX
e+hBw1ycQBjB8dkb+mHDpBsFyF21iAf/NkDCa3Y5/dKm0BPtMCkBPDkUyD1fObaQ
pcb1PXcNfSW7N5cb8zpHEfB0IjuhOFO9LHJO+tFf+T9Qb0XOrZhgw3f6yMMjl1Vd
cMO+x+amQNVXdKpbMOes9qyNzY/QAIQ734UN3O7E2ucG6VpuyE20m6NpGdTyfCBj
iI7qc3CJYJKB3ugCjb5VE5eZ6NfolPGT3QUCi81UuDHkG4b/kcD/ytX6k5CHV3dj
EwNfaN+Il7RtNvWo6lP0FH6AUYdcC9HXOLV0CrFPHihM5RHXZ4LKm4jOdbRYLjFn
1wDPRyk8FT/JEatJs+eVr3eXKJUo+rrsEj3PCQHjRxJ5auFNtp8yST8jWt4MRucO
KrgK6YO0a66n1P/JBFywgRj9do17BPeTYn9HqTsz6nLeIJFqblYjZX1OdDX3ZY72
FxMWNVMOTIaxefUCZBmFmzLGNIYDvdXr08R6VaQL7wd4XfRqji4VcadohSGd+mN4
4dM0rKP9LOz3qUf3Cwzwij3TQzf2wr8wNpYnOtdQoO32BmypjFlGaYumT5jD2rGw
8QpHtelArBuU0fXm1tF8CggcULy7+3yMPpt6TW5O2LfrUKEggEjTiNMKgWGjvfmd
+K5cojHq6ctC133KtfX9x4scmiQXcxVNLzekA5VpX0ngjvsXjby72PFfiDvEbg2/
bFTvcKiyOG9vaYQ0nnE74JazxHjIqB/eKzx7GzsHE0to0R98SJnXxlHaDRcwZp+I
YXXrAIMQDvqoRjfxhhTinBr5ljEjc4cxyW8YOhVeftUCK/VgeL4hIExDJsLZ4Wrp
FkccXEQmrPuET9DXZyqaRoq2lLIkc5Ds3Xfm4pHnX/ikDCL+KUCSoHK95XhkeMa2
Z2TMSSsuLqIRGpiClPcbfWgu9eMR5FM6lbA0Ln8lGStrqf4Nkfm7G1Iodo8S4coM
vLFRXvBmxxuzGDS+txSttY08Zr0h9HPBz5dbk/C6IiM35es+GQyUHdtPUXlFapqA
CpEuwS3uCu1qRvSuA4ArrHj2ZoHb6/IIBIkkC2ZQSwHYFQWTBZZRK+6aFVJRY0/O
KXqtrKGpl/mnz+x1d7cIE1LfviF0gvqLhXKzLmCaty9AN5bx8YYCqW8AI60AQmiz
PKbCNOi/ucIb79GTWdDzbKbSZYM9ZASboqo4IeM3mbNrzlyZO9dIB9GvQAIaFjXn
5qUbX9E+q7PExXd/WxtOkqLimy2jZsnrg6zNH8EOstlTjzG831O5p779XPHQdS1Z
fKbWa4J53VJ4q7GNiK3N1bJ74sI0wXNlzvfZahWzGd2uouQ7VK3TK1GpaYeS7iDf
RcpH0cAJY8a/VJL31ma6CN6fpQEUPPBt9NI8ZfeU+n/GBVytLEYaMynn5L8PyQX1
yXTzZvxSWE5qgI4nf4tomwgxbLs54HZFGS8T7123hc6FmIQSFmHB+afjYgR0WxDi
iux6mdKQ3ffrSSKla5NbbzNUO1gWrevBOmfRPQPgABCKRfXEBisV9xIdW7LxJjGg
YQYKCn4/Gxi870UfxCzKfzkBHtPVx+q8YfC+xwdXDwYBAfC4R+pXlg0+a4UXBZZp
J4a1+hgp01U97I3LLROFHxazSgKbvD82FdOjMk0o+DoqzDcxaftpG9h4SAhOJczK
kIHbyskdAClXwOba1ZyJVKKaYdOjlHmDqHbtJdjTDhlCD0MxOp0Xv1kjMjqeL9X5
r3I3rfdkkikNpVr2lejlZsFYuGY3YnIEbbzUr68CFqzOCv/hBSV3UvUvx6v22qr5
CNkspNXh6Puor+cjE7sckWK2IC28Sj9QyxpcMOrxhgKxysjxbiYBU6KYWMMfEVrg
t8f3mi/27DTZdEadf2GyGy4Xt2a5C8wdugXfL3nNpd/tssVZ6E05t4UZathG/MD+
bVNuT2kZn4pJQuGEULr5w57thlBOEa+f3mjAoIPo7KEW47En1aATBdKancJAMGlL
eeXLTP/lAo3C46gOwjSpGGmWYJBE8YG3+8POQxUVRwObuifMd4oDClvInWvJttHF
pc1dQNq+DcSHp9wqkWuEQDGcuhfM37s7rgBolQSi3dK9jCp48AjqttsQoLt9tZxw
J7GRJN+JRUkJD+VczNccUeQXFGmJf34Zi6HxcGEhndnSWPAO+b8hM6d1ALpyPBib
RJLsvafp1MKRqBCxJQTKaMXXDg6nkj6H7jHK6P+KwW5Xg/kbLwkZzUEeJVxj3ahz
WsoJJnJZm8Ws17E2CZyMceg57R55NjuDArDyiDgx9C3pGfEuZIlHyjZf6wM+EKE6
AAAzo9wv8gDjCKgWEHKLcYY0kZwCIQks5RGufAEtxvJMoE5qt5bdLxtMtTWmvzOP
GYKuMqoYvkU+zWSYqZusk7T3M03/bRCztO/xZRO/AvNSannevPcIZsvnl/luvw/d
0smuU9OLhZvBTdhjBPJELxKdpuIZTIha1KJL6UGquaQZtQuqj8oe5o+j/3OT/YUd
eAtwNg71jFb8EDDYGNTp3TpUiSXaDowK1Qzld9x6CLV5LMEh06tjBiqB0WCOC6tp
akB0BPW5QSVTzFm42UG9TiJqq5y+WC7JW6F8b43pKRg9kZkM5dCJt5fyt5KmWxQE
B3LCvBGlQCg7mxx0SUYugSyN8IztqhnibpLrxVC39PW5Ap/iHfzga8By1waHMqBI
iTHrhQUIcZZpQcb/2/Ey+O6imKqghEihdcIe+BN6x3jpWXTRBwzdCz6daK7TFjp0
yVokRFAnnkMaOFxRemnx3jMkJ1RLAp/YSYcCaGBR2des4uY59nERs8ewixbCSYGN
7neFC5qITuwyA6SEJDG4Lk1aXcf0UIfvquCs/+KKbwa/Ntmpks2WSgpZDdY97HaL
XLGk8ovB0hQNDJUBTCc8cveQ4+YWkg2hnllhsC9AbC3tjAiVInLmBK406mklGXzQ
A7uanTDDR6N0KTC6zOeW3lSNxL1xuY4DWPWAj4H1Zy3nHOQjpEjV7toid7GkrEjc
o8xwE+R+Q57PaJJtCNCunmEezdafyEM48VWZ+e5JHxkaOx6MROoc39VIDRLKyKyI
naHgZPa401rhLrAiVJhSUo+O/5LzJEcaajAxuyxA9FkXB9YidZIsuO/DysDoKZsr
0SvUhnTet+wtMJjbyZQ9oNrZpS3Gy9uDaa52kDCze93vCbzs/2QJINeMyykgdbri
L4nzZZttqk4pvCCQ0Gnb2a6yJY6t1BEqaT+C0aDn8XU1cksvjO/sWFWO/q+UJ8py
0bOFugmdm9bWn5qCnGB52wAZf2MvJNjNJ9r5kYkL8lzgHoKx1WfgozevAlotxI5I
G7EtlbAwhYGnjnSZP7cNfNOhLCpcuQ65xN10hHQT4aezjIsA3ZW4NyslZK+L9iz5
8ix0B4OH3UaDPIWUAx/IkcKUy/zsAQCVsMedroJRwTqVM7e5wVrM02WcmdJQXrgP
62ltmsphr8XQA00D0FZA4B6SMbEeZt0BWz8MFzFoJ5fSpfKmT1vjCigJm2JlEIXd
NJJk3Ik3xTfsDcgO/r9JBjTEcvH0zNplzmDb1N9cWrPNmcWXan7uAXdviMuKg+MR
RaFtsijnnoaE6eCmbwophMPPNZsS+apCr/FeMMsVZEZwxIfmoWsJpXO1M2q3CZ6k
dZhTfdSj3NQGh+ICdB3LYbE+1GAbHMDH3PoUOSpjxXHcdfIbhXvtBVKOu4cjh6iH
60nYx+7WXSn2rj/aArQnM9jNReGDK19LaZnwSGuKuksaNMfIt3lc/sIdxAt/++RJ
uVs4gT83Q5e8iPvc2R/1xMouSrCM/6szihTzEMM/SpR84cQqIJw62xePaxldR2Bv
c/tiz2apuzyHTKAk0hc0QVSV3EN+1yRBqcsF0JIqaCrKegAMejtNn3VytIpC/mJp
XpIBuTI5GexEbfEIaAgpOK2+U6Z0SjaCcSMrtC6hcy1vS9FRbUr00gzMTxiOLtx/
Q8zVCXfE0e4463x4VeWs3HfKP7sgnnxR33GbmyHRO8Gb9yYBLYmvBrJT3K2rmglJ
JZh3pdyWIG3pBaP9mESTw10OhlzrD+6eCe252EdO5ffiC9ibtXFFA8m76omPiTNO
Dxq2iPtw9VjHgOCnRMtsEX7Krk8CNUR3H0WMAIvBMcJzgOTPTioT6ZGtfbBbBQOH
oo2lFSrlxWe0l/gPGYXzQ3xf60Wfc3MDNAGZlVr7sDOy2IjlolzIBUF4zHJ0bxA4
46k1lLnzUxfkrrHl7768kYqN7Soadipvbo4nyJ8v+HOR0NYa8QlFbgSJfqQ4rSKa
X+9HUfpwGK82D+nEAdMU3M6B0EHhggVzB4w+YuWYmdAXhZfQYOQqwvXzHp7j+KCQ
QnEf29yZ2hZav6z8dB4ZGRocx5o0uy95BkvpnlzbGfA1fQ7T9iGuF4LdqYyT8A7s
S3Gu9DbDnBhr7fijwZ8SrV28z8brFtIaV0RBuWfdCvcwbBhzcGoTb2PPst+y52Gg
ZfeK+04jC3hinoIACglegP86aL59MpDo3XgKTz36AT5VrYPGMcJPoxM9GRerso0N
DVQ56vvc4Pht7vUuTW6RLuz+X9nP9prTiu8es7m7F0XaGj6VMUTW9IYOzJPqEubO
KYbzR+tTgGsCUwZcSDdfl1mlglIv0ZsL0CVtamHyo8utMMReloC7gcTzEGsu0HAb
9QvxgHAnP0usbF7NtuSmZ52XMTHIXh9A96s7tPDYmha5HRprsVjgKCsz4DhXlfJ5
CNChAh9kffJBbb3Rv4K/TLm+Vk13lkkSJyQM4gHkAeXsjPY0mkHuF9R3y93WP7F1
jfQXe1K4sP+GVodpBhdxJ3QM29sxtnpOMzGQMDhXAalvMJuoHFULxRUw/tv2nOZh
hCd6XFXAoWkWZ0xOYWu+/swnRJXVojvPzQBSDdTg0MPriToFX+RO41UBynrhvxyd
4JT+Mi6vRO9lK4gExS6JDtdwtlf6Gyblx49pyQZoUaj98WDAPeAlh0MYHtEOSd0z
E3jIJvQ+O7lG/MTy/X7VzRqHC8i309wJjkn60hST05duNV1v7xGdmHZLrVqmloHd
PvHOfb6lBXtJKOjrvoU/0BmRCP+N4YgZyJzWpl0x0ZDSrHpTaFUIbb7g2OSZDrJu
Xfgkkh6K7skAx6JmgSdiqIi1+8IIL07tvduSR8vM6K1JZUtfGINiJExYs769DXmI
glEf0+8MjXrpT5KZ5utXy4p3zTYrC/bbHyv+bkOfuIs8KFKjkO725/jsOk0lzIlW
k8MV48ljXKQZytdUyfO+lsWwNyHi6VlBblJbiUd5qXB90KfIVsswgouB2w8Uc4+0
DRNmfyEI0c6lT8CaaZVCEQC3sEzRYl0wqocw3OZcYcLB4InQSMe5FDafQ3rtF2qM
2a1AydTsuFBmUbX1sp1SotxTURhS5LWD7u+q0wXq4erKdl9za1Wra2zmcttrHQNx
kM/mNjuveOrGNCNBIJe8jNGDWfQkf681yw/Eio+JghsZIf+ynoCLq+zflUx6JoC/
D/7A/AMDcD+JZzutqKX+KtO4goA6ZAOYYxj4rB9+Uj0J3ko2dGP+k2caz3idK+I5
woJQ74xBFvke8klacRCmI+kWe4erCjkmQJDUchW6ekyWbOlm1MTCvxGAJpj+JfWW
e8w1/UABYGZAdPCYhSQ4T003u9nKNls7gOAxtRw7Yva97IkrN4jmw62as9iufX8R
erBGDaPrvs5NMSXQAGHE3bZ4wBT2Q29JR3O81l3yVwQNZyya6S6u4Jh/GWtPIUre
Wn5B/oOtUCbo0VvkPhU+aR+ypZdsdDqroWqLydFYgBgKWyngR4azdBiMTYp2zss+
8CDE6cQuby7pryydH9muRdSmJecHXDmMw+JT0MmBtzzP/d3qRVmYw3/PpWb3MuE6
aipBI/87J+kGl5uWsW/e5aY64zVAtEEtGZuTSSYTD6CGV2qh2eyon89yb1s9aZKB
ZIaUH/Xr3UKVvzdbkdME+a9t8h2mk5y6gtsBsqwLWlxfUMTnYMy3n369YjKemjzT
SgkOXu/4pQXYi5xPEEf8hLdjwvbyWGSe2VVWor0GtXC/A87AWbviMxaHSX1doV5/
rmWaevwcxeImTbEpD9tEsSAzOI1ru0RCCOlcGYBzSVttAT8MEAaINppbV1nvAzE9
5/ChHH8VIGAQDWC0azlnHuZw8r0KpJ1q4cMslFaoFiFh5lANPntFJc07g1xXblwG
eFNulucKJ3ZhcWsCpeiS5FZbPGUPN6O3FzUdMR/h/d7Mn7FEEGnelqH4ftUl06wF
Mln0Bu59qe15fcstKaFnteH5cZM2xoe1Q5wMheABn3snwzmO9CjSmgup7FidGaYs
+wOLQV26gpORYJh/H9XxcHuSqk4ne2M9q75wvJdtK9jOwrend4dgM04nfsD5JFnQ
L7G9IlFK95Ia8IOGnaa8Q/6Yk3vXJXv05iBY9svH7knt5d5gDXpws5TE9BRa9UwA
AglmJr9l8EwwpJHB/Mqd4EUkwnMrqbESkV+8ZmvzrKOfU4lqANHrHwiRBl5FPpqw
XSVEgb68MGj1KgQzJz4EgRUqlOlPB89oe5rw97ApZ/0Qgvcyb1Pu2PdJX2wsgzTW
Y87L8j7xL6ZazLVBgI4PTkTzRSooDJ55ACTYTTY1kyR8Pqg32MtQgG5RBGkX+DcU
A8gOvDAoGMDKiJ7UrE8eUQ5WplpieZunGph4x1a5uO0nEl6Q2zcStt/1XVJjdF8d
yZ6daQDYe8yYDLVjutnGsA+76y4QSKmjqDbr1p0m5GLXlmlHfSTQ7vMvW8dqGB7l
t775T3wJPslY8+rtXZKGOksyVWefRCpP9OfwwDoIFwF3aU4zTSyZ6UV/5nbaENz4
zt0+gx2yndsGJY2n3ZJlm9cL/XEApzIPoW+bz1X3bIWMCPLppBmKdjeHL44CW8qx
Fa4FvaD91q2GE1MrucbvKajvl4ZT4zTQdluXedpBse2BtBPUVxkcY+uk2UFx6Occ
YryiTm/0MqAAmdz1To1Oudu7aDZeFfzTZwCNNNrDLCudjUKHlFZVKeX6Ticyj7E2
Mg+NPQBLF+QJbY3zwCH2Ew8ONnzDEnA+MKrZtBiYS1mYN2pqJ6bSAG+Y63WXLQL+
CW/N86zeKYSUvQi4UgrrmgEo8cUuqEeCgFkZyLe7fZamJsfL3Nwi4hRfMBHHGXdw
KoNClYM8Csqzs8qCFQ6CSI+5L+yZ0f4P8TeQs/St/MVQEb3o2OcKuyDbMEZOfM40
7NvvAMR+wLLn0cpVuu01x9jbsP3+h2Dla36j3GQHhKxsMDvhygRdh1bAJQTlV42o
JseBhXhsOTQ+smyOxkOdhJda/5eqXN2d5CeLZvTnr1J4m3rmpvInWFiMCScBdHrY
z09KagykDYB5KVMC6l1PwbTqteXVjFb58fr4nzX4sp5Uet8YGwxmwqjNHDQZkoxA
53shlYVBj521mKNBKuhm4pXVd6ymC7BC0F6dHsA7YzbnCBYM3gtHzwEVcgfI7N1/
gfxOV35bDWLySIR3tbJzGSVc0hC1+pTt4Es8v7iiGOuskv0gdYqloBoUpHLFnSpi
1kWPRv+GNzdL6gn4IjrYNqAJF01l0HUUYoCqKL/3WBJx5kLfWu5+4P1ODSn1w8+L
3+OKjODDDDBFPtUVtIJS7j6denRdAoT5XlAiZaG76mupCx+p7vK2F8du3q1DjgCS
1bPC91D8jgAXCqIA7Xg6Zf7u6SWgwQmnbxSQq+1zFz1ppNX1uCu4DhPREUeF1YZT
yalnksgz93QksnxbeC31X2q0kLn7/b1W+1zYYECTkBCmeqOEBTDYKh+foXdIep2+
RqlDQNrI1qabG+aI38tzSOc/QlhH+ArvHPqBFJxOOwPn/wx3UbHGDf5AqgVN8Fof
FxVKfZMu8tV67nrZEHks87+cpKXdtBTEjcYR92YUMKb3vqPe+GYga0d47vje7R6W
vgYvlxJQ/hS/PJjpweNgyew9ynEs2WNswsuc9tq0vp+bmu3uAxuwVRA7RhR+LFAC
DtzVE7mU2YDU5hv8KHRVy7GU8tgRhf6Uco4FKPrmBXAg3EoxReErg6UI8YDCWlTD
F77UYnRqVslu0iaeAC5NoYlsMJuiUEPhQ1o9cmQQLDqjkkx/if1VT4pQIGVq604j
sUV9LPVnBNJvSofflc25RFJNEVjiiPfNJ1wpit5KgNoToVc48OtIdQEG8/nTYEc/
TS1OcnmzawtVc/9CNyIfsEMA+BSdmwLQYz6RnbZ24YgTMt6wJhnluhPhnaxnlpVE
EzrR8a2y8DeIpC50yLqHpnLI13sZLa90cQgT0uOlYjYgbtmWfCkUfh2hYpwC9VyB
NSP8gpjrWEFenq/li+ymR8n7CJNO88mwXAlJ0nHUt2AcjqSAHLldZH32uU5nX2Ga
KSNy4xVvpuXPgTUg0w+cigGUpQnQqf+nEqgIFLD+bqt6Uts+dLi/+3I3fgbrnZW7
x6sX8i0G6GoMFzcR1Pl7xm9dGTzxXHrCNl9ZR2AUK3vorVdAW3vlGvur8PLsA+QL
FdWbJaATGgezeYLdjnWnOYecY8QxoQL1Jxs08zqpdmSVIdUBLvcwZj413oF1Y0Oz
BWb1j7sE7xtlIDZm+PoR94ztuj2u11AWiDoSZjZvDzTNGou1/Fd+nRW+uihy11bs
88QSyJGFZJOqC99pO/Vn5XqY+5NkKkUcRgGPrbES7d7U3hRw0BAL3teVWGrGXmkj
iTsvej5OER2bMg0hcCO4iaajLsduPH2VmXmLsQ980llBCZ7b90NAthz/4GMlqWrz
LFFPJzcIQPrglwhe9ILxHvzS6g0OoymkxRFSzrLMfL793eCPC0YPOD8OBwWmqJhC
n6eJsPx+PhGZi/nhWExhzXuxv46tPVSplX0YowKT5CNQ64cJXYA68ZNKigQ2IjvP
wZLdIh5d4OOWY14wD8x39IymEjR1QQpuZF+u4ZBXFdVHDrCBnFoTS2q41bQFd1rO
2acVoHKuRSVB96zmjt4/RDMo+iE+uZ6D99PZ2886gtWPQ4qzAY7T6yT5BJ4TxgFv
KXop+dbXaSJK4rpVHyJ0adcY5NItL50lKMOXuEZM+Yv7+DOYEcHmYNv90oQYDrlZ
ZSOrc/hKYMskut+M3k0SUnaSEv1XSH0SY8GAznaO+j5Ta/vUsGEpDpdoRiGzrpeB
MPL2Fqh7+6KROp4uJ3mVtPSAqetzzPmTC+74jlM1hknLbqOclWN3SRwvMcyedQES
G/gjOq+zDISo5vZLsuMYSX4xi5jNEEaPWJxt9ixrn61wVmogVmK0UKh3tNw4lDyU
++jrFG/8HK6zwrrnVrXRpBH2amZuWwkEpSySIAPFwJ+BjH2Tm8+RTVPROPk1CLFf
Dt2QVBOCGRAiPx0IIlnX98VCNDzXzpV9hFsyGW6yFcxrZ3d08BGbKvBoIuSpFF81
Rg8AuaAZV/4/rb6S1t/QCL/6+WiK5k4C1rqZC/aTKnVd15d7hGUmGhRi+SurVfMZ
a2K/umFvzTEXdYEeUsk7dl8YwW/LY7xlaYQkCZDviHaOoKFyMLVSQ7y6w2UdxdXD
N5+1kPVjvmcXZ26Dve493eg5Ylh+qtRjW7bi17ss9eQmcJ4PY6DXWFTf+yOxPdoN
RyRPbR3iqEhKi9n9LeRSte/vguuCupMq0/4/Rfvs/IsEvy2p+EQ5SzUIAGSGDu1v
zjTD611P+fhJbYXvLFCgXCiIOXmE8zGPowfaSOOgjwgo7cKyU7lHsQdAsEElA8g4
wdc2eEax0ncCRgMyqbOABWEiNgT33XhWkYiQfUZNPSCD/BeBhKeTY21xwNjZRhXD
XUmm+7De6z3ZJ1Wo8eXlHKyqhgaBSeUehF5r8Py2O0ZF6oK5Kq/4D+I9UCOyL5w8
V921ejH14am2IP9afTOVcV3QzP7/f/mBGxvB4ZRJVtzyqnmdcnKag8HRWMgd4FPh
44FUQsTFUTP64yDhvIqKuuh53t7kYswwT2rTxK4JG+17/x/OdsAk1X2og+MaMklT
WLWoadXmszAZW/7xggEgcLAH8Hshzhm5Fa0KNgv5wehPNPtwQvyoTPLEMfDlf+od
h9X+mfCmlnEQ2kH8ZzZloMTeRbmLNBl8saMSWTIHLawlZg6ks1zVCKKQL4ZbWUod
VRs6dC66aOgR0AWwaeUiOyQr18H2jzwlG4dZvCHG4j7mRPlJudg9JTojNm1EXTqU
z/VrxZvl0qv5I6y4i35cbQkIbQLcXEutXHNo9jXm8niMYRDHne3ImXt2QB7wFqeU
7PNmbVfesssf4D7L6SheDvxPO6X8Xnk3cgFzaLTsg+WGKsfyWTG5sSze6PPwLXVA
MpisCVbGIXtFccqNV6NkXNKHynLi52HtecHcVykuyG9p13W+5FJWAN1q7j/7WStv
OHuhgc4+ysuP9T9jqC7oujU0iJ338tTT+9qty4oVGKW+uhgg6jpNDl+Sp7FoVxXB
RUxFG0Pq9l/1VNVSX3GIB25+rCjcJvn0qDFrRXIiL+wHfmDf+tdb71jh4itadfSC
nMilSxLUc5Ylyhxpd6GsSOJQh0/s4dRX3/EZ2AOj9M7sOvKDLxPWonUjeNEI9Y0K
yxeOXH7Uc2zKT1OBpay3870n+/xUd/hZ56z20AO5A1t1b5Wdqtf0+fGqg+nbgGog
tZEjkyw+eAlob6IbUliTS5nKK+v0rzlr6XPed+Oi1yCGeeodusFNeAFn0OIwF662
F8zBL5UKEryEeODtWFP5hr4S6bStznG+Orax8ap0wCMhx7INsUEb/OYOfc2hjVSr
mTM/ymq5GMWE7UaOTJKambAJ0bkQgiKRYi2rMlanqW0sqHwREJXcADsJ4asfyss8
RC280s3ByCwUViB7lVDZ3ya0QmGaZmwlrFfzHf0F1N9BSvl4t1I2MS86thD0KviH
eUnmlPHfjTssvl0cpxTgzxcJAXaVj/+fRhbOBn0uSONAcEFOxP94UTlbAGi8JU2A
C0/nqoKfT7tl/lFBSCDq5RSAy0ElXJgLSCMGw+daq20LYv8x9aSphuQbHDDuTZ33
Dvy7WPY9FEHmUk6QHEzSeE/9eTs+TA6zGmbrnDVztkpR8IKVbbPbxNEyhfZNOwPy
SpQYwk1hRCMWoRcoLkEruwNLT0iX87LUQpewBoQOeyG/QOr1vkWmRfgdjgL532Je
37S8tb36kR4V8tbCda8dI1pUK+r5xjIe8aAEfNedsfwfT/abyYnJ7g+3TZZt9NBB
sSBPAGEO9zvnqTGJzHS568oNCHUecNLXVPkK6iyLXl2gDR2WuoxKunY/Dn12/JZ5
7svRYeyMPxuf1DIvCRq9xa/ElnM9CSGNOX2fVgAYjTKfFqRLhXWC87BbYJUC6eTn
arPj6+iPFYbZAGXwiwx5Pm3oTo0ltBEUShsouqvn7K4Az40abav6J6R8kDeDVSU+
GkfhiHs6tZKViqeigkooBsNrC4YdreMtJxkciW1MHQuX6lIr8jOY9uAceOXGKig4
R0XynK+fhR+6Gm0QvlCeVRN6d7xZVwkrXtUVrHIXY8BTy/gfslkOPD4kCEqrm3v8
xWcyzv+0Gn+NjMRKh/oFsuX7iRRGZSYZhg5VAoe/S8MghytlDR8qmtBbEgbIxZhg
VLr1F7KuofyU7es/pKf+TCRJy5ZH+Sg20d7wlEfCBEzMD9HINNUojEIQuepq1FKe
IxBVk3yJc+irU0s1fwxyIwTD6B5r0glS8vkvGTSq+QdOkX9kuZKkIADGMz0HXYKp
qaepoxyrLq9qBmsILRJcg7NihBKdd38OMaxxw4WOQjkqy60RNgzlIH84xO3dsd+G
EhxOiaAVpMjEEhUIZbd6KdCqrwiXDoUI5EqjeUVFFPKvU17nwgcuYK54CiDFRif/
aSf6f0OfvJYjd4OAq7zzuGC0V5lCj6gi/dW5VLPRG4n5xR+Zjqw2lywppeWLjY1P
EE+gINgBdy567ZDGPTECgSKmdDBDKH1HSNy4UbpNnbl9SZ4PBi9nP4FFry7nJFZy
E6yzrSk8/Rt0CrJesg6H17h8GJXjkayhQULdaENR0X3DGF6Zl45p1UMiRJK2akaQ
rc9KlgcJzCzLUPBHgcCToumuNYvYe9tjtOq7Nz0ajFFMrNizSanVQHDGaBKlxc7P
cADTgZiUEcvsSmtlLgeIrpo+TXFIH6axL3mmr24fCO28bct41vmBSzRDmhE2p6V4
IQz8XjdrC+7HQyOlzery672XVep6oK2WlQk0Lo/FMIlw1VwtCgVwLihI/pJL1AgR
4c7H1Ny0CMcvLE3VPe+TVbLNkZmSI+9LH2MUoH+H4lPukvKbNW+kB3tl5uJ1S8ss
0p63tZJKrbym6EITXevsfpH2pJfpW5i6edY5CzPvtH6ZL+hGmA/2avW2Uh8d40+/
qIJ9d1MS7CgaZ2VThzj2WnoDcMs/gygzeRFl3WCCU9Vt5D/CE/RJX6mQ5TpDJqnP
5DheY4UOLJS0rieOt8RorSbZnN2rZbBehJ5c94aykOUbYSMi8S/jeHtCw54Nq8qs
ZK0ggJVT4Al26qNRBCxU7qEw4BE6dokO6K9jGMporDpGlFo1J+GjNkHPPoz9kXot
JVToAz7R5aYvj1jkz1yaV/kX4t2NyoD40ACoIvBJ/xsKxnHy2bi/B6tTEkqHi9h5
EcW4qxh3EoR6bzTZ0fTSYDTbrj9p73mf0L8NphPosu0WtToKoaysCOFPNmua17FE
oHCX7d75yd4ISdrZwwBOYvaBCgFDRn7lmGE0YlxebC8Q+H8fT3F4TWt3vFZEKu5J
rqre1CWLxV5BgQkB/rAULP4A6PfsKUOWLKz8oxlvuG41CEMFNw0DAwZ62ddVIs2t
yILcLOdpnKZWejcqqPauVMw/aZgXSWHbBhGpn+xG4OJlJyqQv363OWhJ1JudnJIY
Sz6mrk0oyEQNQMnVIomeKDpNsOYp1+aEhRWBp3+Ky+6qE5r9f3GUZmOG4YI3pyA6
5RsaRvgohs7hw3MHPfKuL/7dAEfH6laRGoGV3R+iYI4txqnwaKI8bL7cmaGEXXjU
PJQeeBWBOen9SulQE9FTSAvjsC0SNq2vmgySnaa2bF/l1OyUm5b8Nf3WrynD2WMe
hk9bwe7fLlvL6Htvw4ifAAjldGqvoRI/I/fx39qD9ZIdoQXgiQTjpnt5T+l60Wbf
2XBoWerqoMwWJ+KYUWHV2/79emNzRq+t7DknxPDYkJkVlWOE4pePFcT5dRlWy96L
/ejAslKpyxww0/k4WcuK6yS1rwCSvwAKRfE5ivcxkrwUp+Tp9wC2bewFSO9SAKvN
djDag14v6Y6/DL5cpu9JB3jsgknwFyPTMV+0mJ/n8keCymNv7IVxQ0VVzvzSF1d0
4gOeXKnSkmGz1U9qy7iAqYRYZwhOqbp14yg2tdLb0cKGqPAsa9HgpY7bEmZBy9FD
VUr/wnc58aZKN0C3vb1v6tTNouejYmyQ2EFuUqzbWxGgdx58SccyCche782AY1X9
J+JK5s4NZA163qpqE1oGP8rhUCL+Oid6hw3QQiOemHUe4saEkEVmAWa0gNyafrqM
tBDqRINdZ6msk3qcNSTBK7v5XPbfaSubI0fUi2pvFr2j0Z9qlKaUdbi8IJqtYFP8
6faRxj9LJN4ZxaiF3nxrLngEAVa84hm8gqTqSduP5/HF8Nzk1fnSnGV6Ex95hFNL
2eLP4fcwW0zEeOlFikx0d+vEe8JI5cnn745pKkCU3Gw8G7Uc7/vTlJnP1RSJZeGB
aqPNZ8r+3vua08Xw96xigo0k6oIy0SKE0sGMXVoR/wJFrsBSeMSHOGGFPGS5Vmx3
gMQ4rVrxHu6VfoFFLasrks6JeQ1hayke7wxf09JOswHhunGOL8jVQep0CbFnizzt
d+55dtj4mdjLagixwDfm6+l9zfJnpszg+DSA29XenmhH2iElUMscJBQEOPrCSp9l
E5NLd3wUEX4QW6kShMa/YSaNyMA1Sh/BVEjsVObsCeZmfnhFCV2wUCXZc2RJ+aCl
+j9EaItFMEe0Twk8v/ISUpOgr0Vnp0PWcpwgtxQXb5rh9d7XVRhv6fHddAZsthyh
FYVxiQR4sXynTXKBak6h1MJsPpz5Z3+TBIIIV2vDucqgj03b3k7t9RzW8EJ0HdKM
7RR9+90zRI26vvIiklwj26CvwNidIQYsbLbpNkybNBK2GqOhvYe69eol8HW8XsZM
Ff8PEeaxgQGW2eQogILkOnIz7H2oWbMLJ3SSFtLvexsp204bWMj3FfYANnYDmb2q
FWuQ2wj1uv8GyCthcmT4jPF7yZkjXhzZrEvr3tf/r+AjusycaVzN/ZBFDQVpl5bC
pkzTNNHf9CfVwXo6P6qqzNYiPYH7K5w3f/sDnDzCWdUf8W5nabPnZzRN5synlIbx
wUxVq6i46L9sXWjGQcsmlNA7VTYe54ztLuY1ZNp76aymhlrofqloKCk3Qta/WfRy
2ouzgRcSrtb3IuZw3g+EPBSqjSz0qJrLhl9ZUDVnD9yd9uTxpm7v4b+/ydtObQa4
qV3oS7Mnj5HbGGO0BxEEF7Mjy2+o9y6d/eXYqhwu3gSwpwAlv8ad3+c+AbMtX5Ck
rwGBgsOWDq+NPXSi24E8pwqZVIkaXbACZzSkAbStE5ZJ3XzrGgEK5A4muq3Ga9SX
qKqvH0hIdNCYF/MrMe0Dm0/jgBJ3UDv1aXcEo7W1UqrHXpzjdePmi86/wG2s1nkQ
vlPWu0Sr/c3QFemMSzCManAZPoxBJcL+VPNJ7WOBwx/mmbClZutD+N4RkNrUCHAm
nKAPuM4Unv/nt6BKF5tp81RQcBuUDXZz/VzpVGveoATHXXzLN78vj2vpoJA3JOOl
rZTFSD0xaqeIFCvz04KbD4Lh+9xDmUjsvMkdcgVLcIB9prfXC7i8iDXzyFgi3mOu
+92410xQkAT87v2UxIOkOJJOSuV4FJDwXLnNg5FZk8ymte4L9ARuSlV46CEO9XeJ
RaTXiLeAe4fMS6ENvKTjMyPJgNnLVwo195Pi7PERBiyvhe9gzKmuVHiz/rKXD3JB
GaWXjZvLmMMR6KJ8LDMJ0NKdee05UuFBamJNukDhQIcbBWCDdZAbgIUjtrJ2ZwN+
GdsjY/NURcKWzwSYrl+zQEiNK1bgzF3+0CZPN1jaARdYjgOSOgukFqnsE8SF8nMp
+pX5Eyo9A4g25WWEnqP8B0eD19rhaC+Pp6EEcZUurX+H2PUHHCt6akChPMxf4YcR
n+Z67EuHBaRZJrEuhKkR1TF7sJ29arSWq9okVpBt6B7kzdX14wq7cCof2FZg7ejO
3sd5tRATengOs3XjLcUUn2nx0Q+xGxD7g7PVo9zmT3p70x3e5fOxlw4IZ41eSv/W
Xs4y/qEgBnREvU0P/DuIsrXIQ6usUIg2he5PdxY/Zm3a0cookDFqOdhF8tp/HCr+
ZmBgxeChrwgxRJGLKSOLaaXcsuhSYuRbVjJoyeVQQoGcJPfT4ymcehwg/tYrULoe
dOP0lIlIuLyzDP2DDH11MOoWv7mOTRuD+S8OmCcqH/wn2AVoLFEUXHc7m1Seb38m
0HX8cKsBdAZzs9DZH0bOz/8n++u9nXL17JvyLgusbi4auXjsmGBFrzdMVi6Ufa1z
ETdVDcfRhz7Nwefj/gaI8axrtikWca4YKkei261GWylxLP7WC0Q9jtPNEamlgfkT
YOodAXVlVDMV2N3+f/h/okw8xTZYbQAhevwNYuc9yIGkRg5Co+b+8J0q+Nifji/A
kPcFkzxnQkNoVnvxx+sV4jqXs/O9DNLc77tb7fnXf8P7tX98FBx3idjjXf1ThigV
jJNnuuQuJJyLJi+qajvgx6/ZuosznynnBJpNyHwgtIjb/aT6yuPmY29wRrcYtdWW
d1eq3twQmw2UMt5TGnES3XcJnPwHz0DgXwE5SSop7ZGpTH+VrfXrSuEF4/cnf+3h
vz0t+FfesoKaB9Vqlg0vS/UmfOtz2l0GmFX/zs+KH7ThJVobmPQgjagpG0Juj+6m
+sLcxrNAd+B/qbiGLEARSha2m1MT9ibEaunZRF8n+CVPH4kCWI4M+KnHp/YOg+j7
Y/LVAHxK7kYLtck/LULIf5gMQpDnYaWIlJtzfQ66WiY+TEmAwiOMxK5NTAUV7pcM
na5N5M6RxBYLkOBddLdQxjs7WMi8PM2dl7D1sts7lA3WpGS7I1klj1/aIi/ko5Fz
6D4brYBgzGLUmHgBleJ8tcdLa+LX3C/fFQE68OpvC3H0ywdUceoYHgNkK/xIgCoQ
TobcPZgfykV2c1AXIX+wU1UAZ5F2XfS9EGY7kUwYwAJwXuwRkGlos+Ulejv1DGt9
OHwP2R1D9FQprPPCetPceQPfwWLBk2M0mqhZPWtl4MLQxEXBW/qAvO7qQWM+aYhO
L9aSGGw0M7CVv71fOI/3qJ0/FUncPltqnKCy+eNZQgxzOkyDtWj1pOTCI0XB7U8F
dAPuRtT7qrZ1M9oyXFpe7NJvAFXn4mHI2jQM/UD4VHXwdvt9ihxmqa21xDmqiAeS
0X+qXInmui/kBmC8GvgZo1SE41XvYDE/Q3vFoF6bEhlXWchzQfoYCr/AY9C7zYae
sm/lU1qzEJFfAjfwgDhtuGhv+8+UylDOebEhRYYORhjv4zTVusUxc/Co69ryDXsB
ulV43SOizg7BD+SG3wJ0nClBF74/w7JPmYR0Zz1QSvkPf/++r4Xd6D19OoYH1pML
KTCAVEJjjwkapm8h4DuryPA6nGSGkucuHyEqt9k7vtoBBCJ+ZcKhsL7juSR8QJpO
f+LrDPoFB+AE7g5C5P3m6a56k1j+X7lbhdG2M56k4P+i36viwGo3f+Y/j54dIquy
lsbYX82x52kvGH1xIg7j/l0ClmLRVaNmbxF0SVCN6PtUWUYK5UB/v1T8jW/DRA5s
kj9Upq6m9iL/uZOtG/6ISIaz3PSYnk4uB6sGBD+gHlcjf9xgkd+BG339UuW8Nqi4
PkrJY02fz9+Uoa4nw/S3QUfnbpIhiLZPLNBLNfi0PTB30jAKPWu9y7ZqqPJxPu29
YE+YI7E0LNAqMa+JARUXWi5tlqbuf8pbyBb0aZraxPjRB65DAn20n3g57AaobwTr
wGVUKA9gRlAaWSJVMHTMXzCsCYm4yvOC9t+gvAqV/Uy7mMC+a3tnw1cQtCtpNXCV
YqN+9DMuh28qZ3ll3U5G/xGsn0/kDRgpZ3jO9FQ68dV38Ayrr1C0Sb/brYaHi4j7
GKAUSPvbE3gddbfiBdj5KSgHcsWezUH34JKeY2LRm5gMroOlNNEbd3PNV+1Vqn/D
wGGu3cRXMwVbsGQduOsPQYQsYnbC12rMJvGZ15P2qBSwT/zAZ4oHAKYit8aOXVnn
kZd4Pq2PFIgUuCanZUI/RsoK7q8NOpyD1tdlMenUM0NEoZ6hXtn84q6Ab5CfOujC
ntWm/WRGwFcP4HFAiy+0paAEhlbR1RciBmFPEnzGCThlpvVoI39t8RZ876z9e//m
0Noqc99eYy8+h6QYVcvfV9xvEufzE8Ztjqry2FMbVV6W1qYP5Z5p2S0IvqAzpTiE
+0Pfb2WfFPTuCSZqepmkZoyRFxcO8FGe1hS8++vZabHgPdwROwXxSlN/B6Aiui4j
DVT9Ob5L9YXgM4XYuaCvgUkJtxI4Ccs2kIQ0eCS4Ta+4n0ImCqSHJ5WUvfo/0OaV
wl8bkQuXjxfZWZK4nIEnmIR/xboFmit2BDQ6qaLASmU1094Q9VfOgZYl08ChHHzK
VJan0p054oTENlim7bUcAgSRXb+BV6fq8h4X6m8JSuVrgYHfUN0IsN1GggQWqZjh
RkvBSygIXXY8Ay+hBqqpOsFaAoLcsI7n7llEl76GXvOfkF8xy1f0S1siu+jKQbJY
KTeiOyF+KC4d/5yjyD87knbyJM3mEVP2l9k8QFpU9brunEbT5Kdyn4NPcKRjZXJf
icGoftldkG9gJ6YG2HWvTOYLzIG+WLgogcjHKiHkwbkOB91I9cOGvHMakE0tAjtU
KmtAY9Y1yZxRuuKW+AJzItmh4HeUT0wnYLncBCcFgCK94G0MnPLfaBEUS5/sD7G1
BN2ZPIym2/VC0eC/buG1fCsojLCOh1Yx5iS6xA4feGPnHs5cJQguFJTGrqaBpKyX
H7U0V5AeAYgKDl02mWILe8ms1mcntmMufpWBZqDwf5hG0XmAmY8JlW6Um9Ve4gNh
4D33nklHwFLhss8Xsu8w/AN+Y2FkfHve87qSWOp9jA3xIu4AIKTXbazXRHuvsuTm
zME28WVBLViex/SdX1N8/tlWz+ew7giK2vFhT8qrLjdUNCvugOImvEhcwxIvxNch
zHs/ew0z/ajc2nLYOUXGRVn0Olle2J3N6H7fh5LtHbMhZhnpNHrlgqroteXRTaio
1djHPMV72G33wKd6cUH026JCaH6h98uyP7T/VF1XY+BjlNz0YNDmwbWJnv5I0RDG
x8sN3/OyfeCVQik2tz53fL1QkHBC2EVU6QS4ML5qBRLL2HsrFvag2XiwSYyeEV7r
2BvkhSRTMWUc4wTZ4SBGkyvJPNziVQHVPWqsv+6YVJet7ImTgrZykPqC9SMTF3+5
yF8MuH8N0Q5LlEca8v4aXg7ybr6S++JALk7AjBPfWXNTMZZNImRJiE4uwY9xiLnW
75dDnK5Dq41k678gJji0Lfgn4IRUFlWTi7NCRef9bkbVNlDA8WVr99rTwy5l0FNk
PZOAk2gK9eD19BilCFkf2iLzWgfRlgPERnZw2UI1prSZN3UBY3NMD7vwcsY7TMBD
QWMMy7H6HzwoiBKTnv2pJ7WGuye5ijMUP1/0DD0x9N5wZ6etI01keXxhNdqV1cXp
lEOzgsg7r1pBRR+pvUTw9co8iALrMRGpiktJIcmlDKOcnXZEGA+QQczlvS00yxd5
PWaFWw8I0K+F5j2H4XcyxLwVMu0Ps89IT0l16YIFUBf+yQO12ZwiAgnkrexLxWMR
V8rt4DifUUhsOrxnUMyy/HHVaQeokSP/zeV7/y/m0j1Rqw8EqcmqVVFytx9Dun+m
BUHvGsdmJpyGq/FvJFauMOsje1jQkKcrdX6isK1cdgyCQdChh7N3KBzVJPCdR0Xu
7020yDYCMy43Fm2pelQIRugfsRhbV4PWjTm1cCMfnmblVAp93CEhmte3S1Emba1k
hfSl4PpkbLBNK0H6g//KMJVtLHoNWs9BLwIMw6MRoh4qp6K8ZSJfWanPTyOsVAUZ
MDgQakTiBPz7/FakCQBCyZZyb7IG69C1VimEyHrBMcbVl5VqEw5Jk4yjihMCBYEq
LGdUr7sl7m6Qy+xIs1vUU2iEflgFguM6iK0CTtFFSHOAsNX66LMc80euvaNUfw19
0qU9CIMr60k0wCtBwsgchQ28v4RoVQmag5/Mbpi+Ta4yyVC1XmQdm8swQ2oc6zvA
0n/g1euug4NEg8/9kbjsR27l6Ao2zmyf1KoOOGkmKJI5/IPwkZPmgGTw4w6V70pq
E1pOIpFPPI14yFk7PtlB/cf0UFOWEBmdpQyIO7HeG385kIrpsFtNLroLMKn3b/2K
0vO4qa9IUxbX+a++9wZT9HuyBYVuz+tQSKbOOEx5QU9WDyv6LGvM1ayp85qBDSlQ
pzdcSgOhqF8a+Fh6QzepCBXmJZP9isRrYWJbgTBZFJ3RizO7xPSZwp/qjR6EwU8D
qasA0k+fvPNTpQ8qEF/JPOZ2ox/3PaHcnob6ah1rr1X9gse458kT2PHiFkj26IHR
i7TbvGaC/ETUbZc6x+vmJ+MMqcDIVhW+I3tecdR8boODltWzjHA/9FRafpvzwooV
7Pmt23G5wQ9f8ndaMnugw0V9b0rhBpPdHmsfpQP+Fg+ZY7lVVd2L+czCrAuG6EGu
NXSfmZMrN0Pglh0UxFMPRwCJxWA63YVx5iRAPMdqDF3xHTbP89EvMFHX3p1GIU7O
Ye7Dn1kHN4jUYpUJuv7eMLwJH6129WFoQKfdjW1LI0m/0QZ0E78jZ7jv0Q4h3q3v
er52Oz9v4xPpzxasDsc05LqkaU1Dcz08Ryki34DraF6mAZesSL7B6oyv+WBQ8pyx
rkcKnGeDdkXunZ+Jtq2Ja1vrsv3gpHKEsJFyk0s39c/5Xbi50THW/SdVdmH0J/TO
hmlXRFCGBzGvVBbzvmOrKR/HKVRT5ONDGChLZTL8mpnfqangh9Ocb3R2YM9YIgi5
dmkrPAUYlb35OUNYKvDPrtZJ+x5IGjsuA1F63SDalklhnec10hd809MZ2hdgH3nC
lNCsJ8IAE/+te0JGZoancBmtNE7vJZvAOdKzBzkZrvz+ObJL57y0wbUT+EkKdg2p
bcvD/MeNROhUqmcRB6MyXlCy/hBIyDQB0Xsi3C8TGh6WKb2evmp1L01jiTaXgqWW
eiOmFNxtagrzhG5uZ9zX0UlrNw9/3Nef/JeJYMdX9IrivUbe+Ks0OOioe38ZBwPB
//FBUxW+JMMBpSB8aN+0FVJr9hVBwvdbDiUcHbWSNnZ9hxLe/HB57aH8+5i9fCzp
NTU+nHlS5AU0feC4f2CWySJd5PFfls4f30fsyO+GNROBGPw8v///OTmFsOds5EeZ
cmslXP6McFwkDB+3qD75NE7DNR04N5aq4ztva2XFFE9LeMYrOBgqSC8Zws5aXef8
0262FfTdtq9UZVoovcfrdZSyZ+SPuKGLi45howRq6bRTyWVuC+Z8stXdcagQMGVX
GIkwrq08s3lPdDKXB7pGbFP4Qbpq1zqUoJo7Qjp/nNcXxbBZlTjCjowi4OfUb7NN
QxNGoq9VFrpWj33ZvMBzyQKn/b2ajfY7LgTocJzRlmJzXbc/HMnNt9zttD7EW4P2
u+QvXqhMDpvPs4lNX1y4x92fqLxYV1EGJqiUsBRn845v58Tr/SCKF7NxKeaEor2H
m5IWjKVgwtEq9TAEf2b4K0rS3hEJFCOFU0QZWmW08frPyx/qAMAB2KWYS30jOeRP
sFY9RHXGgRORwo1HYw8NHE1ZITYtTO8goQw6ocnGPPKa1m9R3eUaTjWRLZRtBdfq
Mg/fsfrdFpPHuTaf6bDBrbAxMrZrEII8ArznJNiDbuxzMNJw+4PEEC2eYOsrLwwW
YybGZ/4KaTh54YuRng48WQFdYulyI2Wt7WIsLu4RtrXz/AoQb627qNxBW5m4IkDr
rGU0O2rCggSiVJnFHEHbjgp7scNQap6GskqnlCbjeKq+TF7V4xzSGsPasuvDra92
sRMQt7Q4H58/ralHBlw4PcD5jswO56cR7tjlNbckq6WWEruFIydyK+uL46F+OK+n
BGFvGNs+7gvnAkNR9SP/zfYDGyb6ydc8QTZfduP6knw8eJHIx2fiU0oBhLo/dhEQ
SENmuDh/LlNPOniequNSAl8NmFAJEX+v22G/VKkkrGXCUIJOh3kRBF9oBhDsi6Rf
HRVFXWqT2THV20LLBxxQYiq4JrQn9FgHHbHyaNIm4npjWRs/7ODU+gVIh4Xt+5vR
fC5zscAclcnlfMju6TMpFvQI9/KwV/aG4l6Tl++7gfqEwkHFo5jPCkRjlkJX70Os
sYy2530wD7WZZ37JldRAvspzNQOWIQO7B9G0ozM/qWDv6g3hixVjHMEaXGARmwYH
cp96ruHMa7E28vLtHopbgdv9xK83lwgErPGT4v6ZLJa1F53Ul+M6g+sri26zMox9
5kLafK7+sKrQG3sXUaitEryeY90LDRXsLaFM6qPuAVl6re/CoxQOyEIPgFtgxTdo
/gM7o+kV8OaNU9LU0dG2dK8ZKTV0iOqPcixOtgR8Tg02D1qdxZATIWKIdF2edS/k
s5mqdI+rn+/GW37ObRqA33IMC0OAJ2TnBpxSRY/Cf1xSSoxmhvGzjYhaxIq1nbJk
n1FklW3oylE7Zft7zYJIfHgaLxewnQTXUw/z53az5BwWJ0eLoHjR96+zUz2Ncgwh
Josuh34h3IE0N1ZOlIL5sqiodkISXEM8WiHr3ecEMc0l/9p6HvAVCjsisovC5WnP
YjCA9k3f9Ye4CP/pda0pepnwvUvqDl+FPGRhBMLnDVhz2UOOn0B2w2eUP1eH0OCR
gat8+Kshhvy1NJtd8qR79SfNRn7JIOt3mCpLacHIw88N3KZl6lXO1xFmquYm1woK
Ee0Mga++6LsjXhs4QEJZVR7sFCZ0jypPqPMzKWPYcRdxgCBqrbM42nP1vxeuKKyN
sk3m6nKpfAlJFAP6OkG75vXq5xy7YhiSTTSNdVlT6qGbykVhvDQgbI8XcG6tNaR3
Xbl0XYftQfQzFq6Cy6L5vqt3c3H+TtJfFluZ/F0vyFQ1XMMMQe6Hm+XrNNH4OWAo
HEFJlGNW0qJyz1Nh/UZjg1d55ZgjDpym31D8CSSp3oTWJ3Rp7PLDkCaoqrhGezdC
zHnjZiTSxBqJR15FEtou3oBEUfAAPLkicP+6OmQ/u/OauOSNBwk1qCfLPbA1FW5b
e6nmMOZNap+GkTQAbezrgoA8uNHvKeeDUua9DXAYwB9y+nHeYrZNvx5ywYgKcW29
TuuJ0JldjrqTL2ibX1EX77HDm6PcxGg3tJbgjyN/G88M75VokSud6FvDHaPVb19Z
DZxpbUCEd7G2O7e5Vc34krVnXgu8YlnadOHe9xtvSxN0wve4CWKYtrPtMHlzyYlN
GVXYu47JWbs43NrqfldvF+kjQ85Gp3KIUz+Umk+hIQbBeqZMJ+brqPm6L28Ik3cO
YQTJmA5Ac9UsQtAPy0VjvztEu/Neo7fs8d8EUklo4hT4opIwzxR17riLrzbOLHLB
lseQYS5yBhz/XdkF8yHQ7qofEMfLpNncCESYclDh1Wsj9tYLoDo45Q2Y0GH69peW
Sor0VGsnTg9U7BObgUsVZyM3Il/9Lz99PcMWRJOd+Gl1IeSsrvtqVFCfx1dxsOf4
vWNrVxV0ETyV2KzibpAzHHWkAHQF6IRb6U9j/oZg8AKgcctcBXrECwqLhKVLa/4A
p2nw1AHUNAbMdN5/DKUt5Ciew17M5pyD5p3vB1+OfM9NyLKSko2/3vT1Wgly9QIG
bUZa3YtTw2H+K3Dx4ww4FkG8AHHVGkPXeWjdgv32wDXcZVZytNHOtf3WZgIc9uRp
YDrlqba44JD7XF/+2UCjUOHaNkzLWLbizE2AuJNNAdg9vI1QejptVkyKyG0xP77j
70AtG7WKXs5Y0vCnFkO5o0bqqaemOSuCq5RXC0rrjG19lBnLJsdVkh/U9b1LFka6
9dSUUgG7Hk/jVeC765vjuA9L26dJm61/FjGzwTOAjppiyEs6Fs21FUgVor3vngkd
BnI8kZHf/xBUGfn57zlRAMNsufLEF4B3l3iFLTDg5SkRY5507WrZfBWdTYzXOcFG
bkiNw3jVegDdCWWAB7PDL/HTxrz8A33+RUTUYx5LOHqN9mE/EV3HrfDao1dlw6WV
i+jI/zdsxno1sZhn+BW3TsbDlOU3YT6BPAN6Jl/leMAmgZKfNJtsMPHkUbMAyaL7
`protect END_PROTECTED
