`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98WWHwUGb7QaHf4b03gb3EQwZ4Ac4l0GBo/MeScWD2+QQxBQ8lvClnT/3MqqqYsB
Bo8mNmPjs9PEhOWt4sEqnFZQq77jOROyYPLXWvyTVDqkU3DuH30V3jPGRO2JKBlJ
fCDt1UYhHta2Jw4EcEqt11rNRIfbUY1Jb0v/SJ1qVl6obWeWNM4Al4xRPLfon124
es8jqwZSoAEpTSSoL6PkSdlu5iWCP88Kd3oz7e9fhhYVfWeIJERnqGLoBO6E/Ukf
kvI0DZmtw5CfTLfvqOWIdG9qYG7um4jvjoc8KDzQMtgTNQvEnhCmem3c2JTTXsQy
nzhNnUzwhbPgMcZUnEJnGTvfUlWlH6fgUSm/mIfA1hy+GYIbTXXCvve+ZZgOpF+w
G7lYmZbRq4xmVvA1e28gNIJ1z/cOSIzoscx2zssZhCx1kwUQSGiLGDB8+k8PO/pz
eGxTYtNhS++OsYyg8FHmgZ0lnTHZXgKuruZR6E+vFtkuXnUWP1fExsqYNidwhOPu
1dYVDZ4TamjMrdKsKwhmm9pPs+3ZT/coW1xI2jOwI/Uc0zodmlx3PcY6aT/een9G
6mpJPQmkO9fjw+OEZzYSne255WY0RNOc9g8lwHrNNWBKFDHWnMZu31CS9ZuTTO0C
Wa1W8ftvs09cOGizxFOG1LgrxMViriQL1sq+s06q7/X35wgdJo+gTmDt1w+iSNhZ
1C3/RMdW8TnWhvdexPBkiSIB1VBeMYH3yWd+6QIH8rvipQ1qOi5RHK5i5U+em1Pl
9VE7LCZww8V2MdrU6Vem0Uz1g2ty6AgbTFbUGO5QMgAMp72nqdD1b+bPl/C2EyEj
ZwbMy6YmkXdfFUvl+IdbDlThBzumrfyTk+Tmdlfx/Sl5Yaonapbq1gCLeVm2io+U
CgxwrQxQMtV7xfAeod0gwoAxPesybA6Tu2Zr082nuIerAURd4OD0z8x7eeBG+fmX
q0es0dovi6iYF2ZPqgOhpt7mVHsm5m0VFw08xNrKlj7KC7MZlqQ2ViNnGdPu++6V
b/Qy/V221RamCNZr5F5ykfWbI/kqfr2P3ljQu0AgWkcxplmdr1dzvxjASLRz7jRC
auKPXUGXk3AtsRo6v5fdyGhS8jb1jUGNu7zjwZWzfyvV/uE2B8SMp077Qo1QZH7+
498W92NrZheM5jEocFOtxmG5Eivbdr4h5oc4IAN8NFHDVupstn9mnuK99ZI/r/4X
OEaKX+GN5woF551earAVgsadVlTcdTyo4ZZVG+mXDjDYq7l9jMbe1T/N/Whi6v+R
WxMI3WnZU9SH8ZIeQT0iGGMFsk5TqUWsNd2+h6Uew4BvOSGxbm9//jqmQaQkGAfA
v7Znmg/yPw8G2NVDeMIvv2lUN+2/Yla3cNfW8d0qgFEkQjEc62lYhJD1qlCZt6YI
lt7g+1PS8gpYDQ3w9JXCsEPLVjsF49JoOGnf6m1YR9kwoXACjUecuH2VU9E6W9pG
kytbxoyjra0NeULint60vzhfWniX1rhd61TQUqkl1BkyLzkeRup0SLHJCSk3k+oI
68h/n9Q7KknIjODaso1md99nIHMoG8BrjN9iyKAl6z0spxgOcNqiX6HJSyH7/xve
JKMUARpfYrrNv2gLKvf05ElEhycsA1cdW6g/ida+70YE2md91sQtDNgXwpvvx/RW
Hhnp1/duarUG6IxtMba6sTNzjiAmQ1L5Wneas8WCiU2umgrJ+9TIm4WKXVZyCjtZ
jQiVrEQdIdHJ+0Sx1BttGfFB6dCt6eBtjQuIpm5oE/jtoajUkzuu6oEDUm/cPTse
3pzQmIBgk+umPj7R71uT8rdnLMlf5XJDgAbR/lGA++E1cMT11p/AVwpwE6j8kYj0
+Y8m/eeNrU0fK9IWCPwa0GeGap9MeuVcgQPd/ucl3Qq19JZ8uTQI7Qht8FnZVqId
iBUwn4Gc+wEalWBoG2OwGmZ3DaGXht1PrUGHruEFBCj5nzbWEHsFblJrIs3dEuXu
`protect END_PROTECTED
