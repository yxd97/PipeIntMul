`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zoNZe35fiOD+OBdcfvKIbfaAqUIJu282zXmMfWK1K93xL71TCb8puyUj4p6hmjYM
OE4H0b5k+EV1IEjgPIMElirXIV/Ewq3CFBcWYAE6R1JZpnYA9+dsulsdLRsXlAai
sAVYxxKfKh4peyJIOuaqfP+hoXgROudbM1jNAtIq91Mzqmm6TQrEVyYmZPfyBfuS
/uv84ZTLXWUR6ht+3AL/exY3cH7qgCiUuXUlBZdka+NAtCb/8qF58jwb1IRPwqaO
frpkIgHv0+7lcxfS0jqOdYg4BdgoGrdAKjZoy0VSbWvFSQ91HGSwJUmXfKIr96ho
`protect END_PROTECTED
