`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KppXYpB+zVJJIr2G7g04dljcFLNsb5QUEZ04JTbvKe6NZTxkxkA5j05Bxsb3Ry0U
W3EeLASshj/cGMMaNJT47f6GA0WBZi7Op8Tbd/Y4aMaEWtF5WB/YSe/kYUyFkhMC
lwyxdG86yGpXDH3iAj/PlSTbECZ1a6YclZ4G7YvVCKc47MywTcQ/jl2X+QKUjLsf
vq/o5AyyfL7299D7vvSN4ZlecDpfofMzShnLSSvitymhJpxAx29K1xREdDIvgACd
0Zax5s4Lt1GR1qD4vwrZyenVnrCzf6NRoguNhzo19Rh3emw5HrsdtHS1prHsUKkb
RAWZbOu4TLwtTnqkReUkJLfbDrMUvlFqxzZFfj20Zak8AY5//o4g6USwS4N7OH6N
xxrKhOH2XD70UIEeK/TAzg==
`protect END_PROTECTED
