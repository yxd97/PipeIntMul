`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3djqKXdrW+lk4khFAUH/Jub/kxzQqtADg8/X8WSsdjPiRtYrEQvsKSUF+4+i1r+X
eloCgsTS1GF4GIPy7qL4tFWqgnl7Ja/oHBtX+efKyyWtDtrdhGPNxO4khK/9+PAp
X0ic3CllCiGupiz1jDQd01xV3sLSM4PAIzRGxiM2XoP6X1Krtdw23br6LRZaezI8
BzBFiR+/0VBSC7hUtiRqEdEiX60blxL1zPrWhuJlxStygEjoRZssn/WFJjnZBScb
uW8Em0HgSlpwR1xrMBl+HSeE7VIOa+02y+f8zLS/zjzSydY2FmZx8r37f6qyYy2/
nuCNF3ADWHh3YTJZsM+G5nFiYUajDBo7K7nmp6usQlA0bQ3pORlzwiFflCesqGLN
4abFcnTAikA3N577D6AainhpwALvHXFRSZpnzpmu9n7o2c34Q+yjvXa6mYI4mEHm
AMq4nOcZMstulwHC3PyqFO5tk7eCCCOFYtBUtDzRH1D0nq5KhOLn3PjRO4aCS+St
hC4WqeElF/1W87eIR2i53GoIwbnkcLL0yXPQs1mY+zLRAMJDuX6p+IZj0RtNBVGo
X8jLM9tFrwD6u3WkdHU0rBe7eUHCIRmg/w3yM3Su7Gzgise7a+Okd0qH2LFOdZiE
mfpSZYOYl+fp0wSlZF0QKMFsCSMJXkknwsqQXnMdn2HcV8h5Iy5LzuoSgYxkMsiu
`protect END_PROTECTED
