`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODppJdISi/PX2IR8UZ8pHpJ7dQ5P5xwVZiuMXGF6DlzyxHGydUkm00I8PHuQ8HcN
i/pr+HgnbOwna/32xs6YdzW86yDWFHnKF5CQNdXm+J+5c/RDpFoskdlIx+hvLaUv
ZdcVF6uDli1mtktJ/6W+VuOrYe2G15LVgKidSJXlo/KRho5btl72XY/hpVNIX+OW
wa9K0Am6XEbStkIYKMyRxIlx0LrKg1huB5fxVnv9lXe9c9+lblQC+wzUnIWTyUNo
w9aEYmbqE928mj02/rUdt3S3dFpA2k7/y5q8m2kkaT5AQcVnVHWNwh6dX2Hhh4YI
szGiiuE83P2ElzIT20P0a8fkVbtdMMZ2azJutL/0Hob1ES4n5MDQNB6fo97nFdP+
//WokzJ+lOn3uExy4uuN/3kQ8Q02Ex2kZ4OaJNLico0=
`protect END_PROTECTED
