`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkBnWXPDixqcr0Se+W+AYO/F8ZUh736txqdcV5MolW1GS5qWyMfrj2QkJqSaisjs
qzM++AI8xSXS5jVXu+6HMtYKy+i3D7cKDr7ntm3+5vt65IuBBpno9JBdcE3qFuQc
KyTbHxC0ZZj6N7iAxHZdWJV8+2BCaTmhkiGQLNcchE8ad2XifP33821KBbi71xn8
+kDqPepDaxGWK61oWr8KISD4vFHQ+DIm6VfO1O8+/rKl2pc7mV8vHJ1h9jrwLUgG
YaBTWWOSFRlLvchXfEWcdxZorMkEiQzjSCRs/oUncEMiGsUvN2hd23+YAF58RhyN
e3044+3WhqHVn3FGFvdOYRRVtiWY2tFpWrx00SZNxZsIbGY+rQ8wLRpoiMUeBKNy
nHc51c81VPYtJ/mJ1bTR3YEKFTul26gzWgPM9b9IwIhgdlU0nCuZYC1Z9qf0KjvW
fNHpJN3huCo+KbL8Pqyf917uI3phEt3lqKBVsA4c96wQymOZ4Vj4HW+n6VwW8vER
4Zrm7Zs7cMdQG57PKmYZHvjC4SpFXuSlaX68y0GzreI=
`protect END_PROTECTED
