`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/InvY8qMGaYujNTXA6d2I1df4km/4uXcnmPMIV3Xn51cyWncI8J7MFKWkIDAYDCf
9m9e4jDAd75z+mF9gwkwZH0Zbkm16l0v0Q257V/r2A+e4jn36SbHJB74+i4wg5e4
iLkrAnHISBa13TwlSVffBNUHF1CRRr06NX3Iwv6MiQQ6Sbt0qoBX+vDizR2BabsF
PqJZS+ADaMjIGz35fU3/0Qp3EcU3c2ccigKFL0miwBE1eaoVBBP0rSVIYdnzE3fU
suW7iL0ASjZwUHqGQSRX5YttI727/Y4PjhQx/zd/Sjc3+IKTKhctQG2M7htt2BKa
4e1Z84GbTMQkl7azi2QRYfUjbadqiRTxqqdEiDrJWseExZ+ri8NN3VN6jp3m/pQs
bZj+S2+sGK+AK9lB1hkBXTj9P7yw8eoH5mQ/SnwcYHYs/kDCd3PyeapJRjFxeCBw
bIuKFugRGDYeADeIuw93oWA2bbX4kLWiiwdmSXCYj7dA7raa7HPeI3hGYwnUFf/z
c6vbJtPHk4mttaZfan7Mf2VL6sGMdb84ODR3NAxNo5gCC9xdfv+Z5+YQgvrYfFxN
yFrLzbuUJsyUmrdYksIrOOBRwXAoKJoJarc8M3aDSAr64F+YIQMvhc+Qn9KE+rKk
W0T+EWEhZhXGyl7r6tn0DNcn/3cE0ek668DlGBu1OUbV2FIawu/KUhvBqn2wvXQX
SQhdgl0p2YMHj3MB6JNQWw==
`protect END_PROTECTED
