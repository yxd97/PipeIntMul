`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NJfIK9pqbXE5Lo5/nv/weRjYjC/uTcwKFHzIA5A2GKmpJZNFVxCrP8/lSG+wvD6K
QgVxVxA+XQpu+vvJgoINfwyBgiamDFQn5eHkGp/uRm9WKEO6i+juGLTM5NGbyoOc
oed/cavzqTsPiK+lMvuUNPgtO4zPRUxkAaSJc3zA5fvqlZ4vFIjmPa/o6XsewN+W
3SLwTpYQtdOk2PsbOxRKZtRFI4Kt5fSd82dayaqda7M3h0ucJVxYIE7bbLOPjRsP
TlJzJ4knLcalJLxBoClKodd5kZcYJ+qlC/s41fIIX5HroEoO/r3hpCrmXgvVXcsW
ZJqBToVSsQ5/dwPkhQ6EEZ6vjbllKOyCMh0DUhAdg/kjbJpzjY6VlOL6+g93CMl8
OhrmvRA0PiVtjkp5iPUIlYar25CtDNuZRvV12f6y3vGPWzQq0Yq3agfyJQ6CKR7C
A1G3CI4KaurzYQdZGXCD5sZcLL8M36FI9erQErfY4AGu7FF2muI1faQDpxhP7fce
zhX7ZH/XjaQH50kolLhOMNJqaloUYoNMZO6THEP4U/7gdggJe9J/El2TEAEYvU5A
Nt1yJB1sOAriwFHW4TOVCJpRUI/q0IGrwdpqQrI+JlIRot/WdLCa93wAGxLxWhYB
Oe4c5HAc0S5m6CmQi/FH9l+YPoAPf2TO2dkPZzjzcq+0w8EnSUVUrz9NlR/wePyR
nZwoZ4vHAn7JgtEdpysjd/hADK0kZrD4s/zT15CYJV562HqUkjdnUP6lIqPaZSAJ
BNFkld7hgn+RkRpMw1OENjddIWj5Htb9I+mlY0KpQoaxDwZ+09ungizQrIAsCBEB
APNtdbDQU217OHjSs5km2deVcTnYM2t0QfWaIhohA0U=
`protect END_PROTECTED
