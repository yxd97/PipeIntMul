`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yakOVseWm4LrKKTIbpAB5DPtTHWTWNglSVjlGSY9KmNs8g38vOskLBaebhlNLILN
/5pYmX/5cD040AxQ66W0t/jMesRgSq5f/H1l0uFIJkUH4nMT4bGKV3LyIvbpClhm
tXcDNBFnX/mvL7/nYwnGTKX8f3iF9ryyR5cBq8gyFBdZ5g8edteYPe0abBF+h3/V
WCz/0ixENUatFp/sx6CIdEUZXcxzSoSAkiPelvXLeFHF3RDQyXEG0OuGkLg0lOzJ
qkN13PuLMGaAxkYKD5aIqWSTYx84on1GPhXGZIDblQYS93J/oM4sFA6UqZFSobKg
eNou2Fi4TZlqpNZz7rl+ugLCZQ4s/KdTj1kbB/S5HTH7bIqN65NOR+A+hvqEI+Yb
6MG/OSqlHTWsnPzk6xw3px/92nN9C5IMMtpID2NGg7E=
`protect END_PROTECTED
