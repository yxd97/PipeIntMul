`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNJBgk4XmfYImCaKLkiIvvYIOoUeaEaVXn1Abf8fuWxhqv+xVPpvnSJ1qv6Ig9z5
TXRg5PUDM0O3VUDy4zlGhcmmUzlPUihFwOpwqEKBMp5rNwTQXUTx8gs55kMXZzbb
JjEmkjJ7aLsepGjBKCIZtklqhfqpEanzZQurg5p4Qnt5V7ZDvJoWw8bKR3gEjArb
Xvep27FXHiWZPhzN2alR4csvU2QXB9YmbzdAjy82P0Zi4IV3bmt/U/lF4XEa/crm
dCaTBTpoHZSgUpXBsixKmAOW101YJVOvsZKyljwU6FjCyibdXgD3ucqFoDmMg5/y
AbeIdp4YDEy09xS1cWeTzXth68IweaTPSroORS/o6/MHReTLh4FgHpMXmu1XGMtf
LYetXUnDc84iIVRzxEhHiy0PHe+QMW1Yt4VKThu6zxGLVbn9+N0jBCRiF2fuFsSl
72mlKciNmfhIDk74Fgo7SaQmYur1Z4SK5bNE8ZlUaf4=
`protect END_PROTECTED
