`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuEeOGnLqxaXsz2CU8Mhbp/4JooBVDTlVFRe8muZZZ85t8Gho0N3xF2+07Mi/Huv
9smrFJlOh3bIO6jb/JWW8AaF0ebzt3/N1LhVrkwjNKJbeKkmsMCdMEwcZ/Q/oiyu
FLZrZ8rW2dTwqEADAjyBESi1XmL5KJyeExuF3ZcfpPChwd3AJiW7GsrqZ8EEtDl6
iT1Wo5x90Aw1dsQpyOdpc0zbSXQ0yZthGGjUB9Mlgbo9j5SVJMzAA31qn5m1FAs2
8ZDhA7WJcJi+pQyvBh2ZK1x7h2c8Y6vM3ul/5cHrYABWP7B0hnGZOBuBlVaHp35N
TMz0/gwkvYPU2NOuLvSq6vuQhn3PFpev8OKg4nBhupr32W5IE6tFZ3nW6uPtEANQ
`protect END_PROTECTED
