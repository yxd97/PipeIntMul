`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aZyL0YrkkulalzKBrKMc9TZruTTf9INni386KU1qhMn9bTnljA+zEnwSnJcW3YwV
vkN65kHxrsT4PAV+JZTtAJPgZLOgzLB1ZT+letdBB4Qw3Rg4mi8Ow5Wp41FBi50J
MfbDEX5ZM7WckEILiSICMC2qw7HWpmwq+Ivwe5gNsfYF84nho7G1RGgxRWcQfWlO
yf44SZKdAcgpN6xCURticpGWI0GTabBCpTL2xfj83VYJOF5kQ14f5lxh9SDvrDaC
W+0EqvVgsDjyN71TrkdkCkoYaq+NZgeA4xK+wIPk3PQLWDtP3PXt8FstIj2jAGwG
bRXWhRHlnXSaSRk2cTdbC8UpPEtHe87l4BKhMTEbhtE2s+pnk2/K312v+AmeUwXB
lzZawRkhulAya03QK7BOMxx2oia+yUESddoGiEsc4EDNwOGHwhtpUezNHxey5CFl
Wt6kbO81MrBau0xi+cZq4PO8ypg0NZ4h2Yy+xMB1KD6CvnRRB2oqL4hnuTXKgGjL
m5kFqgd2QMY+XqIc+HYWa5U2zHxLAObPz7b8LRTj4iZmpuEhJ4Ko5QcvCFDv/JZK
KDCxUEmNH/P4t1uFXlZHQ+htctAkfERg0PrtvQYpIayx2FYo55pLUz4xacTEDURg
23KtqOFaPCHm6YZE/8/P+CtVGD+GYxSWm0Zg2efGEklfjz9lWfDxfy3g5Eb4Gh1v
kEgklmQG7KlzabbS33WkXDFDgNHXZ05Ilm2NqkgN2cfwP/MfO30Q15bXa0Y2vbmi
v2FmHjRzLFmxluIytP363G0EFwXm0UKR4oD+iG+2h5/eNWnLgy8L+rIk/n3r7a35
jAGadiP1Lrph+bsqoI6T+zhbfjxedMmSS1iAtOzqLKpdg91zhddABWHofOzjYzBU
ha3H9paK/eWwJzSWFx1ZQGhAjlkzbH3fhNa/hxEBG6QoUYBRqJV135GLDsLtMnac
YfJw661LjtaSgY2FUfMBoqZn+5g5FgDhNMaFt5CTrIPPV4sr4bkgd7Mgccgis2IF
SFTYWEoZIQbQwG3WT2xCadBBJGV3XVyU5I+jh7DOzYPKkEzco0J8pkzb+PtxCV89
24NS3GJ4CKWElhdAK55BsA==
`protect END_PROTECTED
