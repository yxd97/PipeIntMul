`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYqj9axlutMvmurGRFj6aSVGXuxE+Ox9bsn1veDbJErGugWFesFRQByTCjHSY04I
7QTf5B2YoRwohpiAer46mdBweXjg7cmZ/mS3EJJ/k95p+TcQnK++8p380vACXs26
VoAdSjTrfaAT3jRANrvMXg3suFZonndkFWwMv1xQE/tthg9Fjk/EDGYlomLKbrkx
w+myENWmkIQQIgZgXQEXhQ8SEmvLpgiGGL0HgDeofpIgH8ppGAGxgBQe2t5WNbLw
33hEjsFFU+Z6a/g4fMtiKmnDpY5zHkapKyXhrqR1Q1W3PSkKAtuYYkvrI8h00Bub
Dxp2AEZ2AeAiZoLnnnxESRcxlo5Sz4EyDN/AMOUOsF0hzHn9aVKnjWPz39NPQznF
04T0yYYBv2MBfMtgmNHOliUMyQKov77l8dBgqVMpCtXNAp5BT6lwxm7GlbmFMXFZ
yPMClqBUlyS7JhRXDY1lKA==
`protect END_PROTECTED
