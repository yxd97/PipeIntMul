`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8vg+smO1HWWmWN4AfFEtQvDQOmUV7HDpAM80Cb6AbgoVbrWGampeoXo7wIAWKFUy
Qfi019Ky8UhDD4nEVy8vshekS65pqbs8ZudJrEhQj6kPyvpJYz6KSmVzp98WyXJj
qfQo2uqIjzuBIgvIsFSUwW9vYe2n1GWGo8iz3VC1Bf5Qhc+UgKvBGEuPej2cmtLY
jN/qnpnKfRPbSedfqnAMa9vUSv8W2b1Tfl5fsJqp53/Apzm1rKnJDFDtbBcQ0UUh
gbTGUNEbtrxONmUGDlTWa7Y9EW/jY+fnQR7E1pUTBtSRBRv5lA6OstmmJusWF5sn
dYxHq0U+Wnsgegks403s/3aeX89LGPeZYOb4MFx6qOxBgXlmGMHuyMDm8v6KHbXV
rrDhRSs1x9gfzt8hyE/IWTLbSC4G81frF2z45VgH6nlCBWnH1bgNi8RNgGFxWKr1
POyLjF+Emgyy+FDJ+AaauU1Xgg/kuW/yGT3dM1sMiidcNfFk+ObdLlbBKwu3WlH7
+fgoMrGkz3ygMQePgsxkEMyUX8FDV+ftSd0a0R9efQtE8DH2zLZf/pp4wh8tqJes
N10UZNWLwW8msouVrNiyzG2IgGbWfbxGRVFVmUkJ8lI81mjW2GjtMWQUZJvH5gW9
f8yiRYeEDzrCBDZ0CNhWIhZEMioQKYlrj5T6Tpaiyxbv5IxM+PNKPi/xQnhwO3th
dy0rd3Xta+k7+gzoIHo2rHl2Y30g2PF7rsWclqTnV4g5pdzdtYyM61UTxTuZWxau
q7MP2/kZlxn30fMxA2hmiqrLxmBJSlbO7p88tjUT3ey9jJjQ4LLDojnLptI7U+Ou
CBJIgUX7NWduzoNg2Znu2PKcTs/M9/Ae6a4mmqaJHntNtrOulQvMzDpxoM/2ik1T
RJ75sQCx+2Sl0udxpaIhG373qPK/115xiLvB/I3FVv7Nugn+AvPZJbauEeTOvi2R
2tcPR8n58P6rPXRHWK8LLPzbsBcxy/RLP5YJWiaFWyz+0UTN7HA13XxYS12gPyVI
u1kifmao6HWb3nFLIqb6G8h98EAASlJvCjpNIrli00cO+XitLfVsawAPSYAvOkLa
ZnIFYQGv1oQw0q73dHCfBrWEBWelbwIYLOt1QgAEKCG/tT/y7PBiHclwM8LY2ZqZ
dUua8spD7q9pDcGtzQWWcaVu24Cjq5xyikfFKAaN1X+IffvbHN1q5BWAmzZ6sNMX
1cFSrqtpnfRJTrtcycbVEl3mFTFql/rPdlJv1QnDVUTwBOLg4iduJpQyET04rmwo
Nwl8NSwf8TMiUBAggXCF5LfbKPime+ALHGMw4HMZN3jpZ/kO+WhQTpCGJL2e6v4p
aFLAJJO5da0PUgJp1A83klH1rpa4V7pOI59fTFN5YKG2TrJwk8cy+5ZYGMmgd5N0
CEcUfjZZjPl7RQEASihl6jFhW8JuIpkfV5bt7lyA3AMskgZ2AphO5mEC7b7hTI9O
PWX2L25HmxJkw5RIhdukQUxBQ5WzEOWuJMzUCWnmnpGeDn5avKh8FMGjquni5JKF
LbMWU2Of1rzfv8DOCKPlx1Eo5J+8WMF6dFnjwTNWgnJG73HASuUsngMCHR8upmTS
Zj5vq8yhKEnP2j7t1HOQFAwDR+EaXTlcu6AfBzlnnCjOe/1N0POb3lySzLg83oQM
HnaY0I1YgDy6yMic4Zz62KuwK6bZaj1LLjRF0iY6wVwAaS1zrWX8SG4HdFktjcpo
7GWJb5XNp0ukzA4cXVK09dW+g/ZLqHIoVmzGdpkzeXSfHeUsnAB5Ed2uxcSLCwx2
Lv/+lHtDfYvILwqX/Dka7wMmYTM0iAX5qgPtX/y5gkTziXCsvwS57UUhUt8MVijq
oou353DE6xhQNPOF4B0I+OgKZUA3oZBwQM2Ev7nAjhqIOAw05h3/T31E65r7fPUS
uQbMQ1XwgaicmO4imBQZbkv3ctlwI90LbaKOKDLCsjdo2spXnfC2MPJHMOcC+XZn
6px5onHJ145YT4G0mQU/DeTuPnk/b4THRiNVyf68vw6Wte0WP7lLbwCUrskc4v2S
R4ag0JF/Pxw7EGubx89GhJWkw3F92PW1p42E+bjbY+DZdjrVF1hjm4GWkZCuAu2T
H0aB8tGuWlJTxxj1pPOGorWWbqLXzHdlekYlU1e0pqPjvDFrCK1msxghn4Eb/KDr
zz83+7s2xDvNz4bGxxBnCy59d97Jui7WIpGC6KLuY+kF4CqShbQimwnnterETVwC
Jx9AjWICQaC8NbRdcdtp2fPvx23cd9TvUtKAceETq9YJz0bc8rC2TKcFVkVPPL2N
EIbtA4dxZ45t2xnnc91z+v4EeJCOQLI32/CvpK+PoguKdV0+q/EK6qRR8XulKzaO
/Qdrx6eb7ficiLwrksr96wSpGEPQSpzyyVT6rALg3ylhTeeRjMHdb4AMWVZjGE6Z
WUuRnEUB9wmAGZ56DxnPDxKKLQHPRXVTD8M1JLj4Ni9motQCU7AJCptNyoximi20
7Tgr4ggxxjhtFOGOW/vFHZl/xNcPHe16qcQRGaS58FRyzEszhKrY5KShelRfKVrz
5INbzTtCV4XD9nniuWWtZ+bMFjHbsrhwomtmWWT56Txp0E4pYBK2ybGtqMNhwSFU
FN3SXGI4GMrCvMxo3VS3oM+tmX5ma9Fc1tfAC5lFrcxd92Bce3JjexX/OWH3MFEB
Y7DVnvwYPwbyDfDbKPWPLLnQz9NObjwRMfq/hFDZC9I2Bl8bKA/fSJK0AkVBALfX
iRUfWJuADmcITDanuKi9Awlla+SbXRZsy4U8nT3GaCg+nbkHYNaR1JzT2+Rirv/0
lI6CvxodifysSrUyH5xsIY+tJDRErUpmJdKc9ZwQnTIB4+WwmOmFmD8/8Z+RamVy
Jcs1RFJ7w+RSAQNzFVwEpNZ6Fro8/6F1vGBcnsNiTAbovX+s0X9q0km4UFUnZDTz
cXL3a28+g7zenbB5BVw3MHlts+3tdycfr8pWgK8Jy6Q8z4X0gRuQPQFwKvPHO0rT
yxIvFxQSFVYreK9wxJMH5291VeYYecT6EeNdrwZHo5XUZmQ1+g2VQFKweEEpsLg/
X47184BLxSpLL084s1G1h+WrSMyV2lhFLrNIj3im04rvt1AtfEF/ZxqEz/q8Vwxk
lrKOi2Bi5q4OcgLRHc2T4j8JWydfYlnqeuxjvhawhIg4VTfawmbugJv/4wbAb02+
+3pu2OIk2ufhAT4UGGMTAFzBnrTCoA/zuzh14YLGRfFcWIfyL8RRf8JIlcRGZ0Nz
bycGarb5SOnY3KqibsJG2MzQi7U6StDjcaW0PeeGElxZdKkaeSvUICWOGYX8Qic4
L613sfauY0zo90wSkbWiT+GbMxu9mR3j59RVVTJBVwe768FO0dedgHNVMhQYaunY
5it86zCpNqcdGODPwSo+/A0caJjvwU7jYNGzzsDZo6izxMGaxfxMhWcU+81i0qK6
pl5p6fuUfv1Msh7g98OxY8hXCVCM4VXf4/OjfS7vg7wEBskOvcKljjlHFaU30CAc
vsTdphNXRi8oWeSW18SAwSc0GDHrmBaTxBTN4mLcEoinzKOrqaDhx1ub37NYQ6ni
c6RJXKgs+FgM3Bg5J8vY9/ZJWBtCuFJhmuzZix0n7jfS1y3rSY92wdZ8qEjL1H0P
TGhxR6zsT5LyEeS/2L/0eVHv+jJm4wY6MGj27YmkC/lw204asjAeW2ZKjr4nMb1N
77WetEm9dA3ljQ8MG9rl819gDBNZSZe0KAWfaF5WlmFVz6848iZIHNXIZHJeyemv
hz5+4VWow6/2mv7b51H0iJ+MIvmxUw8mSgXU8KgPgiWPG889vL7IV8XSpl0XG8eS
/bc1hXTG13nRLG8bu2oMjnWmwjDv0yxujkyNS9xfxUklP8iQl9eBjxX29MVXLz73
44jj26NfUBnaz1pK6xRdut1IEfsCLsa77so8QLTo4Td2kWGwIw+ucUTeu0wwCzIw
+ldAY71pAJqMMr+/mQaC0DugFm6vhHFqhoYR3t/wh3AmTTu0085MZloadle4pwkE
p9UhPGqIxIXbIZUCpK2DYBcVvY+U1+5hP6Gf/NgZQAdWRwgZfSYyT7+jiC+xrqaQ
kqE2SW381l8zG+j2kvDdkqwhFbwCos8bRiUQkwZh7K8zSGgSQrhonQFXktalWo3q
GbEyPTYJaYSWYHeLszhu0cu+TBsbzHZR3uO5hwv6XIvZSR4CvY8XncgaAT+OfLHn
wBFGMNgjuJo70qhalz2Bh+I1PJr/cFIK5OpuNrR7awUJIevGqjoyVpcJOntpCP4k
vJJaoTuE/dCxhRgeTNAhCMCtlQDPrVNbVP1UZFy4pHDeZS+CDe0SLlrbZb3k2TAn
ZPEZmW6DV3OjSjKwk23lXGNS38DvKVoe7eM2OgCYkvw67p06f5uZFBDlWlp4aWc6
mqhGNn3yBtG1JNTJMEl3VHX8KdjV/0zTWUSav+EwYHx/oE3HpVuNozdejdv6dPlh
nGMWVYb4Vf7OV7/ib0vXsWM+Y84uephkUrfIv0vyMGwIADIelBbg8O6M0KQxvLwE
8XAJIalNuCq2QbJI6c0I6+R2VakyHQNOiRyVj0uJ83ncLGVlYIaNy2ChrGLzckvZ
G7qHkT2BHgq4HwAJGHVkpvBlL/151t4jkEOXOoElBxepDtnxJBWPU9Ybev8xkbmr
pepJXwsRsu9wK46tk6s8uHVjKuBlra555Pi2BeKRGIi+ElTeSLHheZde/qnnrT40
0bg/F6RkthHtVxNZyoVmnKPSaClETuliK7hCQIaUNnd0IjjibUxcmSxN2u6pfgzx
Ex3Xt8IVgvZozv/ZlcplDsTEpfV+7Too392STUN7qWToQDBg20vNBOsRn+MsW5Ns
XwU++OF/1wxEQD3qLrHU3bOB2ssTCLN0VVSc9NLQu+T0fBTVo6ltWD9mavwVFLuS
NW5yv0Y12p7cyCq/7eci+Z+x9V8TDNVBg72YeMMZHOSvcqJrvvK6cYtOMFfx76Sg
qXqxZk4j79mfmDjYqVxu3zx7cU91ZxEQDmNWQwsCwqfxHcBdIaz7Qpo8+ALoy99x
0iOuLlgyh0lU4eqEBP1A4pl4PvKiUknGdGFm0urcQ8pFiPq20Lb5Ni5/RNNLNQe2
7xF/Yduq+ssqVRxQxTtAFqaxePms3zthvUy2UFA+X4kkZsCb9S0ZFfodzITAuR3j
/jrQ28C9ahndxc3WfagsmRcxfobkOydJ7rXiW1ZpSMTPdhbi92KotnK5MYejs3Ss
NBbXCvD9e7uUM0JlnDUa/WFJisob7BvOfabCd47xPr21HLruaq6927UivKivHoYP
VWuoLnVR49iWPKOrkBjnfB+p07FbZBRijj0dJ5oXfLQ0qLUdqnH9GldIg83kVHoB
rcC73J1ZNqFVDKX7IB04aK2eJoVKE7O/XeU2KWsYVkFtH+j7J5LDHI5Xorz0/q8Z
zYoJC9bFioRutYEwObhsjzzmeEaGd+QM5jqnBk8WYuKj0juGVBMErvkVIlkXipP5
r84wy+pSAFZbWxB5oXEjZEPqrlMaOYHp9Cn21zDkyF0IFc1GGclK6EQlLfjY+NSO
ZbQZ1bxjJT+0b1jzJH2nKyR6z4cD4ZSRcsUBGQ/2MELgRN2vC/0o5keXplPdngxQ
U4i2yt+RibkaNiTbXxLvBVlr+M5/J4LpbhbHgMB/m9HQNXcNN9svRiS4TL9KyYMX
u8zOcaFU7n30/FUkM5tEvXcJha4pzA0Ru60EM2kk9+GFUUvxD7j9ydpH75BpHhSe
/3uJFHRWc45MRnPEbZGucPNSFjFCJPae+JW6/VDRLoC5H37LDuFktW6F1dvm8AUM
YBWNgK7hJ1mEMOmmFZVLQ3nUBgwXGwo4tMLFCiR4D5FTOAe0ttN1s1eprdSTIRjF
vPtlA0meqz7k2qBocu2xE2LoRUyJgvJRauwFZa4uok69DOlGiwFkcmzGtWhzDpPi
OPDiBW12LZtXIsKBz14UmUz1wxL4jBjTvwSE8iUqCFZqnw7FRoe+J6CZ0l1qRo/i
M1BbvGa4c+JoczAN3xJXec5IeMtRsh294bBtMn6eRnGS6ax66hmeGgml08z34rmm
nzYadd6CklCdgNJXbm1srzYoHYm8hbQ2/4H7Ikgrj2EfCFMdUozQ/pb5SJLCirGd
vrgEPBd564Qp2ndfJToGX9BCGmMEVbcgcXOuH4AhxpMPG1lwUTStS8hf4QG8rqPE
/hSsdTXREU/RCdKo2WOdIF52j9xs5/xWXt/Regy9W5H0uuHaQEfjsRbZOvrp1dFE
AZlCrTQG3CUEbZFByaVGjUxwMgMLGOIFtA9AWVRa7ql7QWnze6lEMKPMye79RJQc
K4S+Z2uXvnfsbIjFOsjqxqGbr9OUS2HvsXNKQFfRMvrfcbnj3ILXulKWEPlr0e3b
IgRIhTzfiD0RRvMUNzphZPsnB+ycbBtM+YeMJra3tuifE84V6RKFPGizWrf9NO4s
4tnGdavecfYs8XGP36tOQLHLTZo2sLMkf8Th5/OPA7DTaPAHvifPJYZF3TLVNFAA
TwHbcCjWvlMPZjYizGKUjZWHcmzeWWy/jCuMo8TwoCqy15B0buvI6wTWgDv+0aKf
RcJRKzgH+Ciu6BRk3nzIOz1uFcWB8uF1zUuQMLDinpijtN8J3KpAsKersLlgMHkD
q3SiciEekLkGs7e641eazj1RC6fP51YrMZenzIXgGVMLfhh55k+y4HXtoWk8MVnk
5ys+Pl7GtvhWgTwR7jp175QB7kbMAhfJ/00hbHIFXMCreCmoCS2v+7RJVm1RPTXW
l1FRMaAfGVmOJCd0KfgDyjOR/1KCKL6y6IY1JNlFnCwVcJENQ44+DEVpn92fffza
WsN6YIuXf3Vs95R7NHbHCGmFxblb8PRez2OHPjHeAfcQoj29Srg/rg++b9rOCnpB
iFYz+Pp1ZLDm6CqpvAO7/g4FpNwFvREDkltnKVCVFC+ao5ZDr8DLz21vF1Q/GHPp
SJuxB+hcM+uZ5iMAJKEMpPIMXaxlC6Jh8IHKVAaLTcXX1RHiMbVqugtCIYNlvg0+
3TPlm9LuIfEzC2DFkFG1k/GsAAltFp1aqyc/i3BOfM174FGan+uQi9gszhJrnggq
HF2qldhP+9UbeUjxInea+3Yod4qA8y5dJAq2FUprOpM2WVpDsRxtYYslzq4eXhkf
Q2Ma6rnghxximniR2xnu7uClFZHSyW3eanMUK/LBE8fQeqkrn4xmRZh3jY3++mlX
uV2SFm1iO0AzGYdfp8Qe+pMkPJpwg0TqMLq60PVY4RFlCKb/d+FbJFU7/4r1XT42
KGMhEMOY5xbqudCdO/kwBsaMTQAPqUAV9Njc3XZnwZtz6Xd8y3E9yGWsSGUA8ZC2
vkABjG5ryMx4U9TJjdnrNz7koS5KETgaahbcDMHmJVqNOiueM4Kn4xWFrQIyalHM
9KHd8gZbB4U/97EeBxukYz+w0vJ+DM9LMcwOm8QMZiednNzBHqYWH7fpSEfzH5UJ
LSHeHzRjiudCYSdYALO//ugfA340B1Fl3mYC8BUXU+MqjGrVPLWCzKKA0OK9eb61
bIzqEuicGO3j2keAWIDcNiZt8chBDS1jR3TQTYsjHjtTMVmwvFofed3Rq4pBpcrH
H80oEnJS2BQ5BZJoRfaF0uJeTiuagpsZWwYyjfI/3gFLRaVHWtezlg9ijQk7Bwq5
z6TmOo/bbUaW24tqbFyvn2KPwOgji/2RpYmCmTTSHY0bU3sozYqoDLTWscVrz5+O
1EvLd+y6XtezCApCJ0Xxu15Dp8hatPVy/Jvf6X0lmTYXqFtMct5UxkRW7uIkG8Zi
WG/+ccEcFpw95kSX7rqyrk0GYloL6qdoriZSgrF1BWao0W7W+qBabg6JlNQvDC8R
fBUd/Lf/tR39khRiiVWe5Ek+dxwnHnZzKNUNpPAeDfI3yOXAGK3h9QksOEVYV0AM
ECyE7VIwZZcVjxsvaPcwpwzOmVjvwkA0JZN5GA1xIpRdwwBFmjDcFCZFXrx0911h
aVZHcK/p/BL+RWzBulehZUJ/+g0nBRkbSM9FpKRX6t8SGbaLDIT3M8fppIlghNvD
G6RBXVZZc8uYMDbaWuRURcc1nAEZX/h8zuSmMfTxcy8+zgkeyn163ksa8dnanIvb
z043Lzxpz6ecQsup2ioIkRIuX+zHKtU7PDDBvMuQhkFJ2me3m6UcauISpRSrl8tP
wEByFIulDzGyCq1UzGDSmM+AahRjL03mtVQ1qSdPL1r00RGtijldaFHEUMFlEpmz
K/atnLrFx9FuSCrPxA7FfAWqMhPDvbLyx/C3wLHVxRz5E/ybehdjQsErMndb9doO
ibt0C1fSsQDEd3F/Gn+JXE/7Wkv0baH0AkbyPqwdxSe82EXri+0jybqOnfLHm8iZ
Oy3wKLm9EcA/dRptNSAdsbcj7R2/qiWNnwRz5YzovWnCru4jcspPaAnbnmunoaLD
MDenJCrSdDFgsR5aRusTttm3aW5sg6CiAQk4A1BASpHMO9Id9E+4TAXKW2kwwtyq
89v7JzcKXkItyXqBV6EDhvK7weL34w7DziUVI1qraq7U+P6Fh0M1Rl+yt+sM5Ihp
pkBEEhJ+qH6y5Z412+JHmNbrnvgHO2W+eJocTlWAT+r/xFE0x8PTw1/XzOipOdZY
ksxbDL91k73vuqtUlR7Cb1WboztivFCXiZzrdXTGT7N8NLxI8Mai4bXPk/AAwWi3
Fcu60yaFb5RzF0YUPwdikCf3Cgwu/p9Hy4PVlOg6kroDnUo9A3yZpOZIBqg15cjE
0B+6wUXhNB9dPqL8gLGOaAtkvciNkvmC6zWAtkTF8LeSEz3N9qV9qcoyiI3t8ANz
JQiuMWtWIG88l6a4Qqh46frIANAshz00+NJ6D1HMZSQX+rWY9Iio+234pHcrr/PC
abCHsCYU68wHCVhpON4dF7dIU/hNPVeB39zU0H3hlhPNVHWUv8STwch9xjstE9Oz
wUsXjsOAG/7YTIN1lcVsLQK1jKu7tbpBshAGVlsB4V5nP2V+2jPiaRhViRVpjlEV
2K6hKKG+NwASLmPyuswwf6SXv+5BmGhgpaIhY/5qjLGg/3zVh9VA549tYlRc/Ga7
Jq+7mlfhjtBqvfWEGNNfot5/vs3kqWXXRXZbMc/KoKEKYbZe2snaMxmc8RqGj0bi
SvVOpU2vVgiD2dQHZv4/3sWgIhvzepMkV5R9PFjqAvLmb/Th0XBk5IprNnO2iYmc
byElw/DmzXOKe7R/rEaXdOPU0KviCV81JWJtJd9iewRvL7MxBxS4qoPWcwiUmmMH
+o2z4eYBBnp6HUU+Ad71pXGSls0LZjIOlqcqth8AjAut40slnH9aaERP2UkEMxTk
0mKpoMdPVvoIn1NUalVWKXqJjjDNubqR858e4CYIq5jhi+nH0yFpYUB3vMCqQ9lJ
7X6oQQFAbQAM/csUhurTNajIPxRs8x3yM4Pa/+weEPmqcoROJsTid3eVABcmB2ma
M3SkSuwBDINjfDVfRl9NcEn4F3Vt152spVTjjb0jPeHM7A3r8q9xdLA73ZwO69Qp
k26/BOw2YzJ8lU9qNE4Wj6fGIM2WZ2DH2iOmbmwNl2gjHE56o7oaVK5EN5pZ6idn
+zfpTss8TB4N9LPGRKn0XbvzMYOhYjtrE/VB4PJwP5HnBDStSzEB5wluCiMaTuuM
ow0r3oNc+wILqJIRiLMs9sFvmKxoNhwqL4rEY0K1I0riZxiy31f85ewuFHT53jEa
096gUVE9IXf0ywSVlLSJsPvz6JJqks2m0LNLpvL9ufBKxUklcVxor74c6nr+N+7H
5FVBx/xVYm7rGIp7F366Y4ctKtHY3W12ceqhgs/d1SAXLJDrWhXf4eM68XPYeYmb
8l+tokgj9JVp8cuJkR2etRj2h9//OQhj1Ap0uCWS1MoWQGsY+wzLz6dOWf1GlQOw
3CTScWPpdSDqbFsyz77Lu7UPP8mWW2gtecqX/1fUVAWZ6S5MlMxwqP6D61AkiEXq
aM/K/RhVkUgLAZc6NdfDOw+nfojacgLhyYfVFd2FBNhL3e0TCtdxlcZV6iYUn3Ln
qH61l+gDF1xn2ikVAsujzfZQhrT6IGFYENxazaSwOiLCt/FyNki4Xkxau/dc4RJA
rA6bgKdKQAu1Uuk6BIdPGIexxEBy3s2SwQBNAgUZTDtkDYXofxmD0JTWpzXiyRvf
ZRajRmibMVfh+fF4PCM7HDqn/gEiCRDuOX5QiuIhKkKPQzosrYXJk2x/Jl3E173J
ivokVCtNDj0O04e5a/1aUz89TOsB5hvDw7ii7gMCzPwCYRJwRDFDzy0q0KmmWMg8
d8crYX4oAEgGA8bvVxdWXHV1nTkSS10ZsefpQYLhF6U8kghFMXoofpfZNXHFDcgw
vYVRTv96lxe6ueLJKis9pwAPG2dz0xcR9itw96LUiKcjkClPVdts8oqNSNiwvN/B
T5uXvtEu6QKmvXMqWS1c3pslvpiALsJ5TgY4iopgmQBWQHm8WqrTsvR9ZUrZVibZ
sL4AR7r19HhQ4T0OlFfUr9MGNT1qtYlhRmfMRaF4Zk47H/4HRCeF46hVAQIJQeOA
2CWrVElboitPhIXu0oioK8UGNODTPgKfltTpOvHfAHaKfc+sqEQ1he6XfBrWXoEX
VN0SShSzF5SCdNSanmsJSwoKTUtMwCUnSFydWTevJdIc5dyLMFpS+hGLnDAt4g2+
SCMivcJ6WvC2iztZxfoNZnPhYWdjBWJFAS7MLP4ua243kmLrN0TpMUduEKOmSvQC
1C3LVul+z696z0UUFQyoiuYQz0GTACRnGm08qNxeyZ/WacK/XYDBorc/kJyqklrz
8F6b9VNWWB9qnJ5v9vjQqFX4/z9zhXe9XlgB6sZBofonKREtJlrw78l1yNK9b+ga
pSsYyDtjbezCE1nMaqpwDnpl23G7oHRC1dHuvP/zFw4uyLweJddoKUPWFEjTrkjS
aMYexBBnDuC3P2D10287KVzXVuZ2hI4IvbzNEgr/A+vRYPOeby+MO8xmwi3QnBuS
kUzleFwIdQG4McEjyAZ105X5pDFXL1/ehvVdRHEojt8EiaQ/evV9RjW8q2+qrsN9
bwQOR7C1lJKtky6OvYP5lIevrvPLf8wVsl9fEUfdR6UtSwhGdLlt/tQbKa4ftj5k
xAc2ALPU/BlUvwionMtD19UrVieSHx/YhiqjCUBBQjSHtK6GsZMd2dk5m+oTjfl1
3uwbwP4u++Z9P/idQ83ECSUfcpz5bIRnLnZUqHH1lEZBblY0TpEalM3orbR5oXu+
iz67FW46/qa4u+VD9K5Z4c351ukoGzR3gGh7H9SCbGrU1rB+whrx/f5BP3otlkgl
INw0IlwZc3l/xa2ww4TC1vgRLUXXoILXnoaatMIn3d8YCFU5UN+1QYJ0TnBLnfrL
7t/5l2HK9cu3AG/5TVHTg9tlzYXPQ2lkDP5Yz7Rlz8Jiz1dnD3H2HTt2n4L5QSug
sGaIxYlA2O0OciU+oIzvUnqa3j+gtDqSlL6pI24/jdL3BAnRpN+VrFhI0uduE9jF
XtOA2qYjiB4InhZngAL8mMu5ZumU5DTKU56xqTc4zeadSPBbDT8rNnBv8Rz1f0Ej
f6LEYzxPSPCOpUVluNEwBgfR80+TMdiMDAoHpex/TfnFP04YO2sDibg43yNbha5u
+U7vpSk2BvAa1u8/v2QFlIV0JkrmIZIDl4S/RVNQsxW5BqekuDYKDgFWJQ1NR0QR
H5H9gAwGlkaeOdmyHtRMX5rsVadbKt4j3IVUnfXd2kDTdiuVvc+fXkQ/yRB/dPRV
dtH+UZHOK1qZBvswSCd8C/sapHn9QWikqfAU6j7LreV10i6URB6XPtMJaYPYRb7e
f3teVpnn7yVzrVkEaOaUSNy/L0D33qEGliuqrDDvs4RIdGDDIewoTvrf+LCHgABF
XTfYe6S5DAo9wQTcHhfM5PdOhKzREBQ1h3RWMni5eiyw99VzqnjeuKYlLH4QgTeF
/rtRKvjX4gKix2tN82bJtU5fOgE5V0tkOUxx1Pelc/32JeVbx5+0nE90fEZjLupF
IyeJTM2YUNyxHlCCCTIS1T5TFRNqjpPX+eFHhEJRC6AVEhE57BBiTEhuuBrXveSm
aMcSxhbT7fnNl6Bn8AVcC2juTDQFFgH3xJU2HNgaLtpR+fbX0OUNHA/iFTanGoNj
LLSx0a5ZslsyZU8NEmb9vCxRwu/iixL/MmZUfPcsszaE5wOFgBW3av0HD6yiPReU
B+2FnJYrRFx22q6DQIUoLCDN+zLz4a+wDwuuN0sI3zOIukwmVDd7Y9R9KaBkfhbm
7lYOT6/83tTKye5mI/rl7TvI+JZpwbPnU2SUAIBWfBBEJ28tCeULBNabMrGKYRbq
kLC7Vh7pwjTMRG2VlwT0panl0P7z+sOynXHuKGdPV9zMKr/7avreqFKkVkOjH5uX
5W0o+1OMI6Vx0NAgl2o2oQdG/bINfAt4zfoqWB+bhh95/Hx6sKTj1vpIeChq6nEs
Yji4C0h6ARkkarRb2+2rXJg2+YlW6nuMbUDde0xmzI/gGLE4tTIjOS/YKy1xlssb
mVdK39jGrMCwRaCgLYrJQCPIYm0rhfBLdlCkQtMkdwrPNTngMm6RVjaSbhGEYFS9
yBGBs3HT7czxl5vA7bI7xcY8CDT0ArEyWTO6jW4IupPDKwhhuOtJPsyiRY09SI/8
K9U0CFi00ZynJ9fyAbEfmyHuxgTb2ws8VRilHmhPuZjjTU0UyF+pWdMsrzRo/HS1
bMmT0RoJb48pegiB0hX6CC68cwxzOy1/XSfyflBPIl7/DfUzaTbOD4zFsBy4LpmZ
wnOMmq9pjjxGn2PVDJv628tHZbclON41B4+98Yc1qn+GZ6Bgfj74DKPka0axLOLd
IOXAuKDOr77EdLK7XRh/ROOyL9rmZzdZTSITlOEDJMlWQrjbdmH0tvwF246WJdms
TTllyZzDXNzwcqhcWhjU6Cyn6OpvLziHq7Uu0bHsyvYmep1yj2aDQPmHPUjIxNHM
MWMLmL/mb84N6g9faCNrcCwGsnlLLsHEYf38B4+WAEPRirNhuGzgVDGajRFPp29i
rhafMn+2q5BAPoL0qlvd/vN7/xgbkrItfdlVePAB1PmHBokbUugK/qXzbQ5XCDRe
rVcXU6R+jXxxfXT31mCJLk52RGa7lWEbuVwmDDR7gEjC3Udtht+8YjZMWNIUuu2P
MB8nVTYV3O2J2yi70niJLnB+H20X83ANwYnKMJAILjVmdMg4FbjH2p13ujNeyCv9
BtBg6Q0kai7ZD7sHKskOIxfiqsMj2wL9Qdh0w2w9bdkecucNM/YVsPpTMlSJ/8xI
enQ12zf3h5CnqtuBb3qW6Y6kvDp5mPvoPGNK8QE2RAo3QkgHffr5llhLBiu2NDqR
aaWiX8L0KGm2/P9gJzBNJZPGQqJcdD0nz4eh0mrHCSL5hMv3kO22QnrBKdrVL7kF
hlS0YFR04FZaOvrrbNVtMMCNEIm0iOl5RIttC1RBOutwVAjxOyL8xUnjBoXbO/hV
3+UXL35KPcr5Ir/OwhtvFJuy1A3OeQ4IPC8sxhqCTtqxOXMMWBJ5AvFDaa1wQSnm
TBVmuuWURkuHxHwQ1clvXUHxXKECUkRbAdDPkdZjdL6kOnvzgs/G6Lkfp8rg7NYe
L+6iECgHV542Gr0+aIIRQK8f098Lyfe17DbmGNGxL6at76JJtRENCtarZTYyz6Ef
qe/P+urgW6R44bpXqReBEJHYOXgDXv9xDqQU9CGyCt4rKwjdE+9soBKfLyFCefwg
fog167YrPZfqDRE8qL2geurxg4FxfdGMjP48CzAg2y0nKBDNMb2EAM/IGEhXhs1b
EP5F/1WPo4BbqpXewq+NrHWdi9A3q36+tTqqKE5r4kPaNP16E6fDkx/l1+mFMmNm
XqRo/oESdNGgKvn/Vp0E8P9ofHL4ml0eqvRx2MDtNVjuETvoz8CuUn6J5Gl199ez
6CpS8e6fZzNwYha6srR8YO7oYR38VzzK4Ofs8hQgjbz4QbrdIOndQZJxuu/Ty+1q
+tctl3TSMYv9BY6FxegwYKpADe1xwGjvpuYKK/zdbp2xV8kmoif8/UKHx7NJi8Ly
Ibn3wk88ivgFsW0KqCeOdgJZ++QPUWNEM3jVLAd+MALMCOekZil39Ey3N7mFcGq9
Sf8j8obAmqst6fHBlDz6hh+yxLyTVMJdCxJlsFLhCRhN7FM20Vo9tcpk2qHBLDPy
3R0GCeaG84FB2SpRrAfcSFX+lHejEj/gcCa0oBxLb4NtPb+BaPINeQX99wHjWFBD
jz1Qv5gBYnQ7LOjNrl8nKxQfW+t1LkK0ZrmY83mPWmyCENA6jwn5ssG8+qkr84CQ
Z5LFESWWesW13VTjyRKeZglbD4zP91kHS4wRQBh28Wy5jwj8N7NagH034Ml8+uR/
D6KIBR4wrjf6xDWbI9g5du2KWdyIKQj6CeobpmU0VNuIpQaI9t0BQHlwBVkaLaPU
5JVPkQo2Uv8yN0Cyf/MpiLOeVOmh0Q0bxMrVzmKwLSRFGUAZBvOfeG1/KSjCw4YX
yn+CmNYatUEWja7Vsokk1cZw2KSCt0m2Eieu//dcD1J5EySQ1Bc425UVlJh7T3pl
KLmG8h0Kn9gH12iV8qX1IioEIG6dco+/5A4cc7/O27HGznrIaH5mQcjqRjATwc0/
j4b2S7dtfmv0uEibhjqun3zAal6VFjpIQfEq7LDWnKb5W9Pk08aPgBHItWgRkKH+
RLbkSG+aNeex7jDkjdsiPWZIEmi7lL+p/YnuGyBGDpC6+9xnK79MbnjhP0jPkUGX
gdQ+lBZiM7GT7b8KIqBuJGHGihuthfbMmUR04Ks5YWYcStCzW/cX94bFy2rTFAGN
kuu3JONPfKINr0mrhshZ9STDMlgoVDuqVXAHVRDLfvUfHLGhtPObd/LDjkILTdht
wSWiGYV8gBAl0OadsSNqiUgEfNMZBEXCZ/vQpcWAHLbc9MgakbtBsYAA5Yl587QB
jt1MpBEe5WJhqL643vHiqvKAzVj0IuwSA0bMbrg9vh+XdGFIIxh3w3kQ8tw+bL9z
dQC5ss96A+GA0+xXjEMbzCyCnxu7msiZ3jHybYcNfaXhzHaar2ripZBh9HC1mDlf
qpOSMGSMi5Z9hoxpzcq3+wExWCPXas1957w7zVRphN9WNDW0rEyZY5CK/bAC3BBl
hXNgZSZxgyhzFS+Mg3Andfvsx2CgBDOOxsMmIylYaptUXca5ZTS6r067XKq7yID5
cqHX6SJrcuPSJdDm6n2I6SDUfr+jbsbjpeS3yUu7/EIKOtwdCRzmzYuQnpV2TNRx
Nxs/hsB6rolz5VVZVdBlJiDm6KGoJayqoyNeT4NVUzXIApgx7sEQdtlGkwfP5Jph
7fbUWqZZUtbzMXmz+k8XWxnKhpDIhPDyyOw/C0IIirvH73pgSbKbSBx5ufAsq9eD
QYkqB3KKZI8KWRBtEMdr0khz0nJcjwgggMs30R6Tw0/Un9VYi2ebTSwz/2kP/Utm
hTAyjFwUq7VeR4qHfors8OAYhPhsHxHsPE+ubGB0ipIKv4x1ZRYIsL+o9rtRJyvx
`protect END_PROTECTED
