`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tj/a4rEPyK+zmkh+df/NfrDDMjWNlCcs+6UW0oZ4gxboJ4REmcQI5d+notX57JOQ
3EQmUiFN3HFlL4Sx7Omjx+I9CR6R+12eNBWPMQ2g+58V5YlrBJYQnRM+hA7eGVFZ
fU98uAFJwPh8lkWA8EXXfIIcOggIpRHF1jPL7q2BsYFSjzW7uE7s91uAjYhWrnDX
JM2vD+5UbeaW77wzo9sQAvvnkOVz67+n8B56xrQTmU7csNrGD5iwfiSbeSTQ9Y+t
JoI2kbsprSnU5Kx0J9VWPr8mif7qnz/yKBjmpIErYmGOIUtc2O/+82cMGxzCc0XS
Ta+e1NuUFc00M1uoTc7L6V0Vm+MwsdQj3pmKm9QHvuj4Ii6iuoFt41K4NKkdK9tb
SgZOT67u0CPWOIdPFH0H3jMZzDUc3QHnh3HDLsLvXqEsXIyRl5VWSA5n5cocs8wF
7tTu61nJZohMAR6MTaZxsEOOk99wYCzB0sHF0zAkjPIpJ4tLt25VaeiuREJfsOtJ
Ae8/KMtcxHYljwBiTl9dpWWEOqwciDWTDXedYt1W8rgGaQKAe9mgQ5umYVj5wsnL
aNZwrkWRME3m4c001bAdi4CQK/N3+jfNU3bkcccLeVui55F6/c90FQNY8IS93X4A
Uuo2k0gcnwxZUjMDXbj1n+iE+VJGOEMA6lIxg0tLVDY1F2PLu4Bi9YND7Ti5YWzZ
y0w6EOZ6JHP1tRdP1UY8ljBckTKwBo/nLNysQpmXDAxM+KryVrle6JM8dyQVvHCD
8uEA7mrkBzcNhwvRfSnLqY8Qyx8y+dpkrkH6oeyh+4AdZp5l6E/czfcMANqOh3jv
SSEEVQM049HqvbUqc+NlaNx/oCIudDAB5vMjomgl5a/iB5pAAne3zGFVLyHNMRZb
7Vs8FFKo/TVieatYZtydfxX+Cyl/jJY7JnLlccyvt+hk/6o325gWIn91rPp4C+Fr
`protect END_PROTECTED
