`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4U4fyBHycLfNmPYGUq9oagGcyteo/5DOb46e/3AByqFSENKpPcOI7vZBMwF1rdo
hzTwZQRa9dKpi+ZeAruCa1BnZanUkYkZMw57EjDGsWlmHenfWbpHcXIfe+iPXgzv
eP57fUnbtTYcTL4R9XLL7PWdVuTcsHpYT0xbAUoMTu22PSjI8cR4eS1A45kBRJ6i
4gDo3J4115tSujeCrNvq1KhQ0+Y+Rihoio8VsnIzTh7lZixFz9FsVeBcC/Op7org
EUDq3PfMzuQDTWubzHKy7fd3ySvk3Is740pIyVOVYgwUsmdWrePSdX/6NbAKvA/K
SLYnxtr62j4ip4iefUKr/qenufPIOyfdlOWeGABILJFpyMkzsfxPqtkqqG91/qYM
TDyrVmgehFBkVmYPqHBydHRfV98Z0oEYAvsuCoipsgjBGZ0RcWWhYMuVxtvuJkcQ
MGtpaq5ZUHPfynBCqs6ICEGfcwJzVR7PQDX6pziAAiN4lufG99kjRnERKEcyHfCC
nt2/PC2hrCKclhzCbItTuFEp9Xl1kmq2Ig5fL4TEF9KTWF59Ca9piemj90OBdpEo
ywhq5cCVcBOKciyY5eWi5MVOYmpO3xPRTegHUHPnG6vqrXKuZi1sq9pjHwshLnCx
rzwGHFWAiT1U2TzaXwQZg1IDJ4H84qFiu779JszfXEPpYy7Bkd3fj+1JFsPNGg6W
fOxBxD0/TL2oSCVsnGdIAzf2E+mR7PqddNVVbWQHTP5KjhbZvGAwxXofWXny8kFs
`protect END_PROTECTED
