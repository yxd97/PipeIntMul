`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYITbcdZoRvJcs6l0PE754PZg/JkA3GmOPQiQmssADSQJM5G2C2/SDe3UIzkKK3M
8D5J5M28lRn/qUQ8fcPwejBquz701mB9+NQq57u+PxS6RifdiiUYyA36dsO+LWv2
N8OGpm3q90yd3xlyPEsg++nMLa6MtfyO2WQruxd0E2tTiohb18VtsA8Yh/1KQpgZ
rfxUe58RTAMGiFVu2eutN49wNQWxyv7oc87gaTYPG5IvxUHv+2LIvQSQBgnkXb07
r1+YIjppAScaB/wm8Ri317zOTIhruKblimYC8MNsfALxcsfC+NEmq4NJj6B+W+fe
y8/M2b9y2nSw2j63mNHucngoE5bf5CBep06QBx/H7I47PMO1XjjSjMDqCEmDGH8I
/if4fXZrA2q78F9P12sanEJl6RvLEQd9MrDlYhj0ANk5A8Q9sfxgfcY7y0VA5Kxm
GQ83zOUX0jGU256LVw8D5OVHbq8tuKNoHDtKkAeV3DRebI//GiiyBh+3VQ8M+v2b
4M7BY4YMQlRbYBZOYpbPPCuvWNDPfdk47P7rk5mxGlOiE+vCQEPsYYyisG96X1m4
IXsRMtUWDTAAI/ewIvNSFuSqTYO7+VcvmGqFxu54fTJHEmBNvdUPj6jak7wYbUt1
dwxPVTwTnGJ89I2MbtCb6LzcJL1bU4ejHlKsOILm4bJqp6uDiu6QIJamJLsmYLZ6
IAm+VG7CdFTE5OEMMFzMbLe87exC5IP6YEiPAQ1KbGC6fHEvTB5WCqSg+le9TzuR
Nou81GieYz7vtS+t2FArKNcsRuoGGh+4VJG3cJJKTCnvbQV4DgFP0eGRmVvK5RaP
5j5ZRLLTtYJgIzIjdMHqagPqusVZVd4Gimt9ZiHiqK8MfhM9HstWucrwHDZhAXi9
ZsJudfQT44e2VvXEHephPbUViVcna3vfZBzT56VZUzMwp0qYs/m2xHCEsUDiPNyp
uHQ31TlIeLv4K1VjnDPf8WE7+bF3qx+A2qjN0R1UCoLvRdqN5HpR3jBbRfBMup6T
u/oJ7x7GRDOAIApOhVSjt/+EB01yCHoOZsscbCr6WY6nQOTblHEu63Agj6rqwe5K
x3KxP+QWVIG5Q+Q0XRqw+byQ14PLjk812akzFCjGKhknW6/VA/rf/2HIURlDapLW
vZnDDCVa0N+XQ3klc+3fGRNW2z+ni1L/WObuagkGXhkSmJppC3Pc8IMHepnvnxIU
nQe/mTkoiRzeWJVc/r57lvPUNcxTacvVIqFx+T9CJo68e8xQ8rwdnB0VlN27f5/n
3ejKrnWYFw4FpiuAf8Lpj9chDnB0TmdVswAgU4YQ8keK8yz6FVrTAUNQAKBiHsU1
9RBi7qVOHKanwT1x4NLQRJZ/su5tDJUoTSm+le8ZzmgSGWUZkx93SwOHWM95qR2Z
PJwNj61hIMieClKx2+h4HP/3x7bSURDJTnWLwvKJtWqw9k4GT5A/r45Ngg4a2epL
d70L3DOx3YWJdA3VbTnyEXPjsXAGBAVeFU5sqFdl/uX322F4laqN4cvI7C7NerXc
mw/nmHJOU15J/m3bp1YrphX1c8tm7Jtfzcz7gLM4gG86cAG8chGIB3B6uoG632bt
6U1JYlfPyA7/3Npz1Yo8Zr9w1f+J0gDXqhC8SHZyHuYzNEOk//30pMJQKHks49l/
KyZCyMKqz+0nYXROc8E5j9uo4VOMjhNASY955Wra5hk1qLYlkex+C22KuKaEtvI3
Bp0HL0wBd5TFOL3E2E+7wTfy356cZoix/Fd6qSMwHqq5G0mTI3owXUZkAmit3gfh
CsOVXTiYhkfyvrDC/DigpZ3JojQFmQka4O/S3ZCy7b61ULIAA5Uwe+FFuVl9tkEF
XaQH/CPxtsTb83eaMLrOd2XudvFdB3Q9iPQYXBsAzK3aLbckbi7tUALTGjHwvAp5
YQSu0RVd/Qb87yG+ZsP1siPhekBmB8dRIUgWb9273RK6tN9xf2x5DVxwqAcc1krN
mNbbRU7EBnwxosRGd7Gf63q3u0zlqUXJkHnZ1zBm5XKubrQXXdIfodbKFVVTfvm5
j9/aLW8JjE44WHT2UApi5nyktfpkcTZo0a9Yn7k4cmM=
`protect END_PROTECTED
