`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjNfsabuCUak5AIRHUuvsFeQxyP5QNyF12DMlSSccNNYHeH96Eq0E9jwq3OmYm4t
f9SSbZuUEhZ2LranB3zZFA5g44hp/rAHQI7MnrfNQCSUygfvy+0FnthRXC3I2XgV
iwThXW+h66I5MJiD5c3aUGyzYKUxyabOJHyy3+bnIusS44LCn674eOH5BYLz8n8g
g7pSBFFKxF6o462FtIpSm+rLIoYURxmiIG+dq5sFHovrHyBWn7x64f+8YqTGBLyy
7W+FuRLAId/QzW1dgCr/6qoeQilZOF8yn52skzttavyr8X+IVurvqebujSUaRO1E
Y/hywCqCVboUfyNdNFZJRE9TZ2xXX2bifRbk0itX0ZKlkT3Z85qGN2lB3hB+KlgH
zs4fuVNx2npONWPqKNi1tb0IxHL/XqYXephuepnBvyMvB0EpbJ7arwhmKmAgk9yK
24krOiqAVa5zWBi2uIQTXap2DORnEvcutCWEO6E7VMrIxa4FvaMMqDMpwjiUh+NN
QPkpsXEW7nrKLg1ugqU25shQT5p248Tvjw+wyPTXiVXp3hYUC23aqfyTiNXglQms
zohw+ssuJodEYCCgMdFNcR0BfFsI/26YXpz7H/4hKntbJuXv7no4l+Ws/erQAIZ8
UyzeNwgawDBx4o7FMLmoRRM4B7cUAouJ0Na30fMEnY4=
`protect END_PROTECTED
