`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QsZhY7GyR9bTfkHTsmgO39tvKIseSof1Hd5+Ftoy77oIZVP0JYtQODEzCkYx4tnZ
qwhsPsfh/jrdtJxn9nAz/fJ1oQ7P3vbksrSpHGEUx9QYwd26+IwbHZzZoxTRx7of
Q0j7174F2a39vw8XKrKHbiEWbpwWEFHB0AT3uwTxWTyoF5XSBlZU++eUr0kkZ2VB
BGHV/YBB70MCyOogfRng51RCZI2DyAo/NZ3Szv9LXhTOoxnT6hoOuFS+B/TsJ+NS
zk5ml8aVeE38viNm4mlM4Q==
`protect END_PROTECTED
