`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4I+sIpOtQ1UfCzowUr9paaZja2YsGW3WyeikGcxSUP/+57dmTjhAmDDs383RJiA+
g9p8RqTsomck+ZpKak+p+auYExU51001iGCMhfonhVZtKFC+V6piLPhjSEwYCOtr
G9PCm0SCGcjKuapmCYBtxUBkU9Vo+Nn0wa1L15McbChxYKiOxbOvSbrbGajvBER0
GE00sA7qV3+gbsrCyjSv5AQtg5BurzyqdEhi3RfDL3KxaCjgiZOnltWx98AbY9QX
auBiAkeV+rMuGewNudY7pib7k4veCUStHN5j9uROQnrUVvqgJXQbx0j691HKLUwY
WNVMXBZw34ywcv0gswli412rC+nIlr+WBIIZVZal/kk=
`protect END_PROTECTED
