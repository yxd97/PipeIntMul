`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tgg7TRTmm0JKr0EmtHvNQ4YWBXMy7D3jQkLmEGxyEwUOg+OS5xPql8zhCqk0CFl1
RfVZIy3IYetyIB5zSmJbcH5dIwa6qWGG+tjmD+8Q8nrV8VNyHHedYoU/oAnEPHER
K0GqgB4fflbrIRUjFx2p8QOyPCZRxqvkK48ger6F1q9yt7N/vbffi7N7pmHhmEoz
Wu8BUXmURG1jmrvjpu3g84Ou1J6XgeLLmb41nj6KT9itiDFVWH1Pg7nin5Hl3yME
y7PxrCoeB9WQw6eOPYzt83Zn16p22LuE/D8RWt9Y9Uz7/qfuw4yXIoRfEjygeKGy
CZUQy6vF+l6YM83qlsfmqRigRIFcBg1fS7E4J/jGZTzXBSUgIcqX6gSS+BLAjkqu
fw4tBdgtTdDEJKqcWvo+sf3vzpzrLpFGOWZgsa6ryCz6nbFK/ZY65Gfh6xx5QyRd
O9j8fo3tG3Nkt3FL5ST55ysI9gm2XV07iYCOxd2BrEDDYFlcCwV/kXkM5TGKwHDD
3J6ShfeSCpFKmhMyYGFig9mBkAZvH9b4+x5hYj1blUgYEjRb/jXkLQ8tk1dr+RYF
BesX8Fvg3p0amkFczFVd1aHC7VRBbcD06FYJs4HAWLAUzfntrKKsClmHww40h5Zr
hd/nc0Ixu4EOpiWrr8f9uzdkDbf1duj9TdIlFCOTindVUJSNBegUOZUGxEplYyxD
GDPh21qT+41KRgrBt1/670XuSVmTwIbe/o20QknAMkSUOg9sGhopv0DKYArqeMR8
16cu5WTI/CcAfQ08NT6xzppMkvBF6XHLVrORQ3NqljHNuq2X6L6rx3YTENw6O5Em
MOwD2vf6lAIOnQfe5HpGGlQwrD4WV2RqEz3NDslcgCI8fMyFOweoGklcdtUeXuKW
Zqrn1WKY4yHBEzL0NFJJDmchUTGCtu/VMpBWsVmSmhBw6rtrwJ8YkJ2Y49FUTEK/
`protect END_PROTECTED
