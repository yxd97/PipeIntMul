`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hLFX+12v2H0Kx+JZJyvQ5F6XfyLcGWq1gBVdKqOlSg3khjhfpRxZYxY6XUV9azxh
IOmEgjl5o0hyem/3LfLx5VHhGsEllSdbLvMWBzYE5j35TcupasFBeEM7P5mtmWW+
dyV6pktpIG0hF9XjGp/0EGSd2P63ybRXU7juqGTVMGqwdeq9sqHAwYk1Jd2uHQOL
UD1nI/DdYJccrksWdxlLO57I9IaWo8KOHbOPtX6NEG7KSHp2g0QuiuCjcfGsI6lO
VVXMf7KGw1JjoI2isIsDZ0GTUtCegB5zKa8eVWXHaCQ601CUha1tXiXCVR8lcV3y
dRwsbdIsas4hvQwYbnfsBOrNrjoMgC1MwUOoCtyH+4o=
`protect END_PROTECTED
