`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GXC3lvYVlp7KpKPH+/TDIt4n8N9gYCREoEvTYRkh9St8Z8ePHZri4CwrR9hLYIZl
2M4sDFi/AossbNay6Y+3KjyvX3sglBKAvJt1rxCmWBCf4tJXy07JQO7TltQcXi0s
op+lMarwHfanc6FG/FXZUsj2IqUXruUpUnB3PKqBKLQkpJGIezKdzA7N3hfAjyoX
yFRTvMeuo0EPbEKti9F2MZyL7RO9fpCzUjZo1P7AtrV5eQ/JRz5f84JRSzC7BWUP
EhnlBZiLa0Lq0gDtBJ4rgaSKq1x5QnJ6MLrBrr+eQwo//mjRkIjjXe10w2Zv9beK
cJbjbQVK/xCfpwmXHdGLPLcJFEYdbICb9kTxoaoKONThjX8tJZSbWmHQHj4pz+m7
XZK9v2yWwlr5QjtIefDFgoh9q16URLetQGzMWI0bSs8Z1WyC2F3fY96/keEhyNyx
A0sDyhbTn/gUXNvJ4tPegWALjXcit3cXmsi80weIWadBbDGa4EYyAgfidq6Wup/7
ozbmQ/y9nZyXA6+uvPVT2p//IR2Eij4GSvAEozLQgq3l7XYSDG/Ilm5fQ3PkYUT2
AgD9OvOtucXyiQmnXbVNgqlbDFIalkdw9Q6/QlNxEE8tKGBfVqRD3NiJ6SsKgwqy
xtqMeZLg52EeXSLtAipC+MSkDNpHcqlCXnrmKGNkwFWwLKjxGdGAqeddqibd6TWZ
wteF8ha/i6TvBsk2/hK3hKFw7eg3xvs00jLED7yLUF1xigYWP8T8/WWhbeAfJSlM
dUs8UkICdZwMqQj1D0L9mfeBqwG/sAT+JMZXBJiztyOrICI34cwRjvm7xBqyB3zM
f764ctryGMPw1HayrYFkY4j+BIVw1TAOnmeLX8F4E+S8Dh6odpJu9zu6Anj9oIbS
3hg+2otGFNbQNNyu7sLRgQ==
`protect END_PROTECTED
