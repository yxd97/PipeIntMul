`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFV1xG1+0Mob2mudxk9kXJ5y9yf7ZGbY2IA7EH+4NDC1RWbADujxUU/4+o08+Amy
92D5C/c/7532e3MUCBaPjUpzfTTWtQDeq1rCZZr7IC6zNaT3P+FuR38qNjXL6f8/
u6xAg2wotpYgmAfws7r0VbHxq2/i7V3MUrk0nc0agpeut+e0VKa0uOpmFBSfy+9E
zbccIs3f/f9/iXIwpv9GMol70Pa5G+h7Y91ioJJSLCE7m1YcBRpsRUwanZtXOy0k
LbVkpMJ0MaXf9eUEece5jme07EncN4GtdQLqE8gRWh9+evuATKDcPUDM/q/dHB0H
SaZRsfP3IqtRRnHaEmMflh06xcSbwfukUC4XzmkYVHjgBwRJMRqhp7PMmxD7mrDz
ysjBu5z1oudeq+N2Hik6GWCbIPfuXBytRayw+C5hYyE=
`protect END_PROTECTED
