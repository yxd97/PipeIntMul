`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k/dKaRjDJRFR6kjsiKSwzvd3DihyoCvCICU7WyMp17uajOHXXeXYet2ag7LInCpW
XxdRJX9d4r3N5dNNFtx+q5QXmz6M0FhTt3cMg4Jt5lXpySege85gu9v/4lkDEATA
mQ2mH1rzn3AdmJDXgkBQzWZD0mg/6GsSbkE6XKS257aFMMPNTo5GIJM5Omc2zjra
xP/hj4SvtWh/aMvfN1Mx6J14qa8Rdr5vOwzdFuX7ZAnyVtvnIk/9tb5NhCSbZvho
qtEq+4M0EOvNFR9GbvsBEFAZNOJ6FMsFYxMObU/YhIwULEQAYazidU9ZhuZdUdLn
rWT3rVIO4IqCqUZ9TDh+2C9KLUSBtEJL2BNRh1iCUft2PBocToLE+3ewvubhomaW
x8Khyylbs37GVJPfe36TjF68pz2ip7DBNRX8aBfNMO5StBKT1dg1KDaWZ9WGGAYJ
lFQADYPjKLwC9ANAnkW4zh0avih5rIGQDZM+v8pb4LTXGHVsfFpewIrGvT8XhvLP
XSj6H0roPm5G9YrBXEw86BsxEDPD7vLRSI85H6YqXno0ZuXin3AOsPtqO1zYhJCI
9BlO4WQhkhUickMEJgBUXVuUaqbjoDnred1HkEKdX9A=
`protect END_PROTECTED
