`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TkiBLddhxU4KQqxHN+mUrDYl3Cfl0rsaJWUvdkFUOKYAL8XfeQN4dwZQ4YPllX9H
onrXpjYPot6HIfSjHuUqBjwhLYDCU9llLCaGZ7fddEYVgOon1FhhatCipC7l2T0v
8CmJ2OtiJkCaJUPtHzFDtMYOfIZxTKdccxsDGAEEJMUYbRQ/syDU2xGYxwvuSyLt
HIp7BkHlNXi6rxsnQGUaEL1Kk39yQMu5s6F6uGoJHlg/WXzsxSbAknUVD3zXyrMG
/yqDq6B1whdBVv8Y+UrEPW/r08OT7V9kgtiJDywhsGfHja8GuDE/x7W1/Joedn2Y
XAtLib1BJrDYNGtRAEK7UikG2JWohfiQAVwo9usILzxm0dCmIdJ9figcYJXsAMhx
MGIQ/s5tT4oj7ubvRbpkWJzn7Sujj1MYAry+WVUsb35CxKB2m4e3g+YfucA9/kan
FZRGgJOjk4gmLqqYkRhXf4M0LfrecPKgH+YxCPZRRHcFHGaNU9P/0rFwF/0oSALH
QyuZePgx52I+6CMuDKV6MfenbNvWaG97Ge7XPtv85SE8mV9Apagse2AHCLryRdXc
6O1CvSrOxUiH1UbGg7qiVpIWRRpm35imVw0pEkzYUwagvHG8QmFwoM3Fj8a1gL89
hPwlP45wG31/fBNsDSrP/b45fP/saAVoOZ0+fJ91t0mGY1oWB3Xqyp4q5YRd0Ywq
/nXRYPn+i9Zvs824mJ+n1pZ0Mclshex/Sm/RksTqnuEqjJsKIcTMUOayowllila3
7/vGgcsqAiI83dFP200RnlyzvRPZEXXGyKNUPA9zp5az91LbViCyQa7CldnnWyJ7
tAHK5vmoCpJL1sMz/h+G1Q==
`protect END_PROTECTED
