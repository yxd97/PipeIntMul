`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9aeTGXm+i0ObDYyC7VB3E2X6vCmPeSVU9LO0aQGIkHAvY/SoSO8weM/CHiXFoxms
g9Wdar5uvNmlxp8Ut+a7eoQJ4qs9tSzhcg9Z57IocThYtUTBu4OxWnGzSy54PzRt
ZFSf3hU/CYcV/Loa0F0+K9JXcguwMrvaEHy5GBqA+xwEcd4zmvv3/VDIzzX8Gx/t
bUknCVJ5ptzFqPBcm/wdTXJWkFbhzjCv25CNpAmCkcJfkwlW404DD1zkMlUQbc7h
f1bjlmkain/IsMbJlUU/2AG/LFzRr6hfhymjtwR3tMius+pWOW+8KiPmot8Opy4D
eVRmxb1Kh8Qj3WLP6llXARc2Z5tfqUo/VFnka7St2JEe4v4zY9sOXW44zsv0izRp
`protect END_PROTECTED
