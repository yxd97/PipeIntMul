`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCvz3mi6qELuJgWHD9oYik7k4idV4oeGseTMJaTCbtmiPV5jpyPCfffU0TssRtgj
diLzeQDa7aq5UVKKUNdWnp+fS4xof+KxICco9sdjdO4Is8ca8wSMbbDgKNPnqlUK
671nYnGZtZudfvFhEkfzLvXwOsGynHxBgcYzwGUU8pqnGEw/+l7l2oUk8SsZhTgl
PVOCcLY4g10vPNfqGz5ZzEdB6djURd8Ukeb1R0Ja+jRE9DITUMcTE1AAuxq5KDW0
zdQ9S8Q950WkmliSIGS12jknPvsNOjE8rfHuGwXVTdGCuwl1XHHnc2m7LajdxRWX
YVOv+JIaq5ER9AIGTG+K59V1ltjoLgFafwO6spteCdeT6xvF+LzfruGwcMYikCjR
Fb4tQlsBNq9dHYXf+llx2BJuqBUUH8ZaCQPEfEgtMOK+HZ0oPe3X/wqQLqF1VM79
7xb1rvdv2x9exQZ788p0FzUyiHpQaQrv60zI3xE2w3W1eV432EG2zJvDJv+vGT5s
sgUFNDIKIfFkkKareICABQrY6DsYJqwT3zepww6R/0pTVG8YcL0Ezgo4bP8enHOX
uuGmbbc98FHL6cIxbi4rS/UEUbM6aQPl2MkwycBJPVpET5i2P+BHJxt8HCoMgGU6
2mdqlYGEx9pFcCqtbZsA85DM6oneTRwilUQ2eJJePAYH9JytHtYR9AKBJ22siBkU
imJ71Y0gLA0PIB4m0/edGiFOAQggVaz+AbKSMVkVrO4E0Jqc1M08gSBc8HMnP1fb
gCSw/Mc+KKejQ8+5NTmVytwIeHQ4DKcdfNZQhspsnpKBXWK2VIQIs0i9fU6b1Po2
w9VZZzrsrsLKtISaxGMZ9YX+WVSLpY8Z2tzuQiJHckmp7Xi5MSwAnNbLCRMBQCh0
tRU0gxtDgXJMo/+hSAy9vrq+mZbHCUafRzQ7Tw9URCN1Gcsdt4Gi3YNB2Z1h2NLr
INBQaKcZdceGq7uRlf+ZRCd8/g0o8VaQaDivh/cpzAQNyaqsV+0jce3UeU8VqdCs
qHBwHW9FFNKcZx/LRpAhG9aSHfB7VuSXJuEL8IG1qNNzBQmBIHBiKguoTyaJqCOq
C3oILnTCpFW7iUq+P7OiR4aAQzJkEjwugHqVmaFfpVAfsVaNZpeUsvKxn9GC6GhO
4n+bdLX/9UxJuyjbDjHeT3MEzeKcp5e1UuClWtdzubwwiFegYGo+9l+gbNEC01eC
oUKK/ZcvVUK5y8BROhxfY6pvoxAg+qZS5SvxuvgxJnHHWgzZP7PaOlToIu36qqam
sVupcq0zAeIAosoF6flyViJ64OuJJWtI+f5VrZKMZO9s9TO5lucnAeHw9w+2no1E
nCgv9hA1DSb58Q2+3tYLkmKWwUgGyCEP0R3jFNEDgweoLsZROHgksZXEd0Vz5a8c
AXnziKmS6kR+19VnILb93kABTiQ95HGPZ3rVYKyAt01pQT3BKQCdxYXiM/40jWAF
z9u5RFL1K6JpIvqEY+MnEWZQH6Gtg4COoRtdZb2wKhoZlLQpB94r+u+Am4Qk2uza
V05/E0v9TzkTAyyYjoQhgPeAQ3pmJij+XInSU2M5PV6NFce9hcU2fYTPlSSVInwU
mvabNu0W4pn/cA/r0cIuHPdf/TdlLmNkaqhJ+yfGGFjVOc9Y742YISJQpV7+vwwn
SnqSO1qslKI98EXEDS9/Sei+WCw5hn9l1GYIS2xyE733fYdeNl/m+1JydzddIyTg
B1j3TTphGtbQ5VU0ND4KGt6zezFLNCEpN8hibqIYifRiNrKNfF+bTh4xHMfmRbxi
nOlietUbMsSn0biHyUpQAeZSNQrZEc26+Uloi9pCZkqCj5STHuHkls1SAZTta749
GfpVk+U5fxyGxB9KAs0I+I36W+FDC35yqVu5wsWb1iYsmmpEqJiJhsNfYDMp3b4r
rWIXU1qN60TUI1gHE0FwH+djKrdCfmU0QQCGFgpQMpj57Foedo1S1IbP91rcTG2o
OmHz2a4+Q1Uz7fjqZkF6lUYoZXZ4gpctTJxornw5OEgei9wnWiTXFrbW7+pVqIxx
VLAnqSouIMG4W6+ObI+bjwVvQmeH4eOZHP1CoRJC+AGX3XffOy4DVdKdnBr3141z
dBRFBvHnetb2M/PnQxn0xRxB+u0OdbTPvkjoc+iaHH0/YbMKKJvm5xOUADUHJJxz
ujyGYEglYw15agqD8qF6UQ+UIZgCahF4SLFldscERWkUpmpnI9fhVHE37In+eVIQ
pBZ+1XhdnXD02R/v+HOEKJ2/L9ru7TE+FWFH+fDF9lUyBU+Xd/n1nS3pm00jhFlV
h1agUqe9ZscqtsTDh952cvIOn5s1+cXHL7LQPyafjGQC4jEYUE4+uKLfyuwovbHr
Hx/GrY4sHC7eKO87FuxYxbYzup2muaV7AJGiFPiqUJ/7pBWGJtlMD57YG+dLB6H7
4whZ/wTgwG4HHkZjGOSZ+CYrsioQoyw190XcL6SD77gDSFZDgzRAg3jtwyVAL+n8
Xevvqovm469jfMDEAfaYRyQBJEwfFU6reWc4AP1PZsk04r35JmfYXZN8SF60Ixyk
JiDc/H445Tqbj4Vl8NPu2VlDOBpQTU3/FOHfg1Q4Nkb6q/2JXwj7atZewLjew6dR
qwGPUkR2/HIer30Q2OczJx2Y2bSw6PV7PgrMq5Q2Xhd8XlYmV6c/kwZe8rqqa2en
VVlbD+4kxTFiqP9R1HF4SLmS+eJYCRSOwceY1okadCtrOR/Jwlo+qsKh7gYVhWLL
fq3gGncv0UxZgkoiShAF86+U2MbUgAfyMObvsBOabfM9XOOh5qG7xyjdJxYauIc6
z6P9You7bG6nA3FNBzbLVbzhRBVH1mAhdu3o/AOKx4lkEiyC2LIUpJguu5tf6k27
HfOZiLurOqfzx5Hyj2/2ninE7Inp5AazkY4T/pV7WjzbX9rdfDCNuCYwL5WBOOd+
lilM2aM0uCGCWrE+06i8utRii4Z+SkhKueINVGSVJT24V96hiRC1+OMKruxHa5uS
x5RmhbFMBu4HNNjjtD6BSNriJ8jNgHZsBEoDsewlWpbuX8JRv95/NgvuCtOwi+ds
9cuAbrBWtq7kZXSMSojSgH9sdHEdbQhSEJN/xYuc11YmIOd246iXArhynjFgFAvh
zgXulcehnEuSpFuaLzSXQIVzb7N1Z6xINL6pFwVUUEJLPHkP6kjGZhhE3XSOgPeQ
lFrHGCY4cGTlQSBN2AspGXPqS82/mHmGyHm+7kRVbiWO8bwCzBxD6vhsM9qyTu/n
seLcPEAE0wxXSbuJ1HkUaewt8pFwr1YW2XWtK4+n2u5ZqtYXD9F7RLADAY4Bj8EF
4ksU4q0Ab3Bi76uwG5u5mCG5KM3imy0ETEvestbHqjklTlpjtOoKpZN44uoJR8YJ
ZmwTnYXsO5I/MElFjkn9asxOmPWYbUSxfHQ0aZb6ZUhEI3SpE4yAeZensZl15iMG
7g+WPfctcEKxqwoWcXlyDtuTvhWc4vmyhUHBNd802nJvxxGIlXMIhLdCaKshZDzh
NCUGqMt9GfpT+7dWoQ5D4aCeUEzILLJPoIKqlzZr1R6iv+8BgKuIIhhm3aMm5l2H
BHNI8jCXgGf/e0dd1lRtg2DeQJou/ali+/1BNh33AF2GwKKERrE+syeAPEOm9Azs
Yu8EO2OpZC9gVljqekzcpXeRQ/9hCjVj5wpwKJZy4ETMDLqFZz9LVSoXmAYImm0+
P+ettk4dVnGaxdjLj4hFcFKgKTz3S0xudcAkjogfOSSNpfhSImDj9thh2EsoMt9R
iI2XxH7PiVXsRMrGmCW13iMKyejPywO0Y1QkXSQYOhWEEAhl4YQjeyN6JIjUoWpo
pMFVMNc8c3ev0dAY6nOCjQ==
`protect END_PROTECTED
