`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCY3LHbCwdN6mT+E9N/4FeHe83dllh892PK+A9ip2ZW7vOOJT80ioeQHKvUBADdc
1aOfPezpoc5KQ9SFjNc946g8LYOziPLRX0+UTYSIFcG8FsV5PD93+4RXYTywZ9ww
co2B2hnX75O1T8/+XfYK28mv3ITXBG96GQcLkrXxdwInyZRmPfKFvXxtknXMb5/e
4JzUvO4zyBCBH7Fe2QXL0KuJ3KwapLG3Ne1I1azLeKbgVzAUYl2GoCxsq02YVfJs
SVnIWchv9LDpv5sVlpIU5naEw3VoBKqU3Wp0o6kBTN9HhCPX1im+jALjlrDXfS+f
uC7226s/sshZAqq7Ay5Hat+vKRSuuG9LtLule+q5ao2z7BRl+J7y/1PhGkGzH4z2
JQz5zsjXP7zQG3aPBcdC94pDPhzzQA7s6PDuIb3zwc3Da+Gn7tQiwqkLo56bFmb2
cCDfQ9VefxaXrkoas6sjV9JodPuZP0P1UYVipdD3ReM=
`protect END_PROTECTED
