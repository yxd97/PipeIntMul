`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tdbat5ISk5nPhhmaPfd1YosZ0OSLH5jFyewf7FE2VbPgxJW1KBUdslVCWeQhKBlM
mdw4uqmvJY9H2Ci76h3eB5JwBRWqGOe8MAXuSGbvqAZDSCrvw+Y/PCObb9rhB6q7
k7OvCDV2n7LtNWNaTsoHLC3Tn7t4DG/QJKMKJWcZZbkVWQGnCKNUv+k0Vd845rw5
vqLoURLJ9uOX6j8DceAs3bsKqdjKhBfAeJPmWe6xP9CNjssQohJlGwmRl+l0nLfH
jr2XYSbQRUU3ZaYuyVphE+bT3co+QDgMMmJhYZX3nf5SQEFUm3IhWijJcOtWmLZ1
lklBHz8Lf6eDixlaGozQUy1f7vPo8AKPqMudIJQ0qMZI9W79xr7EaQ48vt26GwxY
lu6J++4hSzPU9dFlbQC0HcoORSCKbKw1nInkWMRiOvnClA9facaA8p3Dm1IqlXcy
hcBeEXqlNACX9uDnyphLKF6oBWSrmQfGDSOCDO5F/Ljk8K47kTakCYkF2+xpb3il
c1I8XoP3aA65P1DHg/bEFmxfZYXyp4F2UiIk6KbdYr4LWc/9uDrdHRzn3rwrALBA
uccBwXW7avVtGPyFJI5fYlVx4BR58gmR9DhTppaQ+5lMrXy+Kpn3MQBx/Sf4onD2
hIUDZDF2SH6WIa+lgcWu7ppn+uTc794BB/Ti/LMK1CrF6TLkdo5fU5aqoVXClN42
Cn0GXV5XqVmdG6FpywyIy2tswsIUaFA7wyH1JEThi3zjk9sbR47TBMgDA0Lsd50y
`protect END_PROTECTED
