`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QKuna1QDC+wTp3N+xurPP+7bOgtTMVbqZg64jUaD7HCbmHZImrlXccgLAAWAbj+O
6PdqPQMhmXDgpU4Exn32/dFS8Icy1NGoF1zsLRbmbKpx5VSTv5dYvCdPhp0vJZ9O
mnYNhfoAUjpsaZlu5YiKXi1fJblQndB/LKIwjq8JSk6Tj2BzYg2LdFuFHX4pUp6m
UwYrey2FAGCJhyVRnWXt6ae8+ujnYLXZEt7YbBw+ODGdCHeRW/6c38CGtCuqYbrW
vpmNM4wNHF2I24CFt8lGJWO96fl+IfM48Kj5YYUQ3BhEgn7XO3W7ntU1LSp8k6wd
z8CKERqaZDDvySg+6ER4XvOWVbtIPHVyMb+6iiAmLGKi1gxJbXovDXHbkXz1b0jS
wmPmaLxbUbi0JUAz3jTCWCnBpZvMlJIfgfjnSGKw1LIJ8A7x0BYwahXt8Zqb1ND1
ocwnqQitbis5+P6IoK7tUHuKHYa508iE+D6dJzxGgloTGYcGwM0iCfuwcTO5ytbg
f0U7ydnI83Z1ux4JLoCRIYIHTI4TfkBqy8bclMIdJ7OgNz2do0+3AGCDrPmC4Jpx
J/B3QHpFsz5NUCtru+JNtv2pTUVprZvI+RjTG3bUr0v1LXP0+odH6CNr6Kmjg1Pl
yV/dbW0sXZVQ3zMgWFpmbDk9MDO0UXC9TSo88RaHGPyOwENGHLQuRxMoF0b/8wdm
+z2oUkoZjdDnayYLvA7S11/4r3hEvjBa6hW6yYSRqrMQvOwhWH/qsOjT85TbxNw4
RhnVcDrwg1ccrewUhp5DWxDlP2XUPq3iM77Rviy3lW/XQ1dYtpre7duD4ZShlOa6
TYc6Xm8fdQywfSw8VBhZyC7jSQiAI6Yre3QNA6DFGIV2h7IIN92S4REZh0bNEQIq
5eRHn1z8IRLIY4fXANMEP/zldKD8q9Bybz1lQ5GP1p3Ul6fSy+DFqWxdQ9lx/BnY
x6t9H5+NZudr7bvns+rDqcrLWb9UJGkqKaZ1oSBoJAK3YS1PZnMCVH0RIkcUOcXt
7ZkE44VHj/IN5xcpnPQfWhjPmRT0S1kqi+y5GxMcRnMtR6UVT6lcf1fT5B/hXAV/
t+9bmq0gB65Yj+sg1s2A5c8XLeBUph+lAY+Ka+WlRLyB0wYBG1u4nAhnYCZD+hmZ
tYVq7pAuA3tXtZheb2d8dMpirRUq2wtrrzgp12qQH95pXq40YxQ62RyDkqSyOvOD
Ed+qmiurZPcriW/mzh7vNuLU8g4pDM5UyK9ovbGgn7YtIHj978/GsWRWlkpHA4j3
/fGDBScuwgvNuEBuenT9lH+EUkzTCGatAtv9TPjx8yxr/6f4K087dGnm3I/9OgpO
ij1zhh4hyRKa+ZavSOEdEpIHuvzq+cqzQadwGVKSLkyjm+m/zkstNUrvE6gz1QNm
H441sPSCmbZb6zgCnqlQQ+n4tDD+t4zVB6xGOLU/YU/ewQkJRx1T625er0Wo0+iY
mYJ6DyeqIJHwrrBX29bUFomik1w0SFEfxFD+mXAZhd71hHnK2WT9mTKfjMiAKC/4
SJgluuAUfxu5c4Ow8z8hjbcP+lRSk8XvXws3FXzGYcM4xP3UYrmYJaHZvjXfvMDI
NO7TsErT0ZGr4wZQVcuVFNxI75H5B4z78cUBLFBT0uQr5PEss5MmO87lw+2tu/p8
g2A7CpYA/uR4yHMqRQrxbMCE03GH5mW4dxMw1Bug8JfkVH7VQDDDROxYsaHlstsz
EMIMPC13E9Kv1SUYi1jce6ZUPQQwVYMbu9PI9SgAwrDNS3Fv11RjVfqqj27fjhMV
kaNO8n1oW/ZZ8qpZZ8hX/udzhwPYraXvy6l/iKk8fCGuUe/M+ngf7jV7jkugjIhR
S8U1psnV064mF0DuZaJKEiGbkjxXykBbDqCqV5Opq48N2te+0Y1Sf3AoFx/abB2m
RrJq6e5SfDFWwfs0C8tMNhtwIbOe91+opHKi4sTJgbh8dQ5Fx7eKURuC+XpyW1c/
5wOAhu8jdJTbbT0KxPqNiphf9SzgjLbF0uAx7h5p1c8=
`protect END_PROTECTED
