`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbCqSmR1HCWztxpd96/VKnCzUsA2LxSI8vFJd0tb+FWpDm0T/DYCi9+Os9udsM4Z
9Uj/qRQWxC8s9d5/GAQtdm+U70r7RK4wayw6uc6w/3KUUJCxbd9pcRyJgZD0koj8
l946jlhI9Rc7ecpKbCDn0Oqp55rA3QTfAsOuTbSzPiqUaorQrs1DMqnI2dGIp4yV
PQGfMa4KPStvSDgtVpRKZYPEeVf4g+YKudMrNvBaXVRiS6zsLTbF6oCws8Zl0K5K
FHXatnKjXtvZDzOA1zoK/p8QywfYlB/VOwg74AclQWkvm4mAXbQYYRP7eDsjp2Wq
YQt2MP4k+qGspplCBi1HsA==
`protect END_PROTECTED
