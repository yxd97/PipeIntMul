`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vX8FqnRa3XNDWRSpXijSUPOw2qGteuxIGdJL217KRh8HjfKd8l4Jz2ukVr/SK66Z
1vKZyadqLOxuzBVx3aHAkoKXI38XOlzGkau4ic0+Id6PG2iTljQu65YdcKJY+sq9
F7ZjNzRzeGEveQ0Vt9Bic8WsSNFtFJkgXWD9lVrzl6TGqHbnMHyzi+d1b/VzETLy
PWiorFLuRICyZkpuHdKzE1CJMjybvBIKDoM50NDjgLclPZPIzRwvqZmuwJxPEDum
pu8LWwWgBbOS8qQ+1cYZhhDy91kSxeRxwZWWiIQO5YHzcl6XK1/8XzqGlwIxOS/B
igwmI+XStbZadyxNj1MEeY5i1NL7GiGhIpDrA6waQHvsmzN6HRFvDZJZoHL0Q9wm
Nh2+xzbXQgZkyYOWwqNFUTKD5gPT3GW/h2j73YeaKH8tZsRgREjNjN6C2EaOMnTE
kBy2Ld807h+i9HvK96hJ33Pf9XLcbT9hMWOLkXiJHdmWZCSBXPFBu2UA9vfKeelk
XerUBBXatbk1SmrCInuCOrNWQsncIug8/M2uX0zPSMmHiovT7gJYgs5qx8+uDL/x
ASITDixJOqNLzSm+QGZfYCWFAfF1z8DCG5c0mFfF2+LyRe/PL9rnKC4bIcbRMFQj
442lqWvzg458oKjYXDyjNsgD34BLRSJ74xc6sDauRmfnhsjTe5ZBds8PbbKveKxo
jUZyum2DCphGLFaoW0WGmHu/sJ+nyaVrfunp7q/XWpwHVRlQlP43cH1YThy+TOXx
WTg8OMWknwxAS/3NvHQUYvsXdyCZXcToNqyCu+RGAN6f9OxkCqUN+pBISOa9XWtX
kYl5gbv+zF9gnZDV9mjMBmuiZxokBQZIPLH5sMrM0gllavrbWsyRR9xXVqFuw9oh
ctTfI28FrI6y9B93pCdYJy/QoqXRD5NLfgowIBA7yq4=
`protect END_PROTECTED
