`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+bHsdPawsawfvxNV9yNvSRv8JnWcyphcekArtbrTerIg+CcmrI7/ZxR+kh+fotC
RH5sEzqqRgdGz/3wVbWbMD6w0FklEV8NC/jA6bfKDcK0zoGj1H8+m7q+NFPhycba
FhBpASCATndiqrAVa1vsBad7vF/Cp1jf4Jc97HWtl/sXKIMIBD6yUmlox5HOy/bM
URrIbuUgL0/2HDtK6bx2Rj+tZ+nR46yK/W0F34etbqFhey19J5raSd1i8eRJIrdD
uga3WSJ2Dp3BxggQRMMwGTppD0cDybkWX1ImLSnpt6ONLBv/BRkleMgDQoe2XJMc
02KTYFt1G8LllcTUhbzXfprf2whU4buqHByJmv+5LOAMoLvkD1+gyvmMAh5f0sf5
iwYZjiNQOTKHnT4Jo3BJ1P00I+1BzahPLusuJCKslpr9e1tZOK/gUPDdthRa9aLm
17q+02FtX8Q45V9s4C4LzN/B3HtSaNwCqdEC71SPE72Ne6JW9H30qeie0+4PuayW
MKyj5b2/FIpvso6TSpx47d1slo0wY/wlZFoPP9HeRoKPEH98kSMjLCPAaj8KNVK4
xgfu8vu03m57Xg3tgS39Qo986dcv3p3Pn5AaW5/cvrgX1hODxu3JmkcI+SlWJ2Qm
kztH4WsNYhYnEqT2rcqp2zRp9hUZQZKvhxs0vK1F+WX16oqUbppl2JZMhFkzj8Vk
EVoIjugCcvZ8diMVJ2FlWRGxmL1XuODunwHyrzO5Gj0vPnrE3SzoqTybioxqGlJu
OO2XOah7sMdI7EbzKSanZCkAbN4X7ON/uN/Jg/6SbDwFfftMAly0OpxemUTEALGP
OtKhOkDkekWv33qJNZgDjzlO59pK5A5IN1NbY+jBTAZXIxFPglW2rIjPLUnM5H9I
UE+60kuROnF4wBdm8JYca0AEhfgOA7ApjBV/928GYUGLT835B80481vuzmLmA5aS
pfhjIcobYv+ui9jBqjY9H3xtODtg5w8Q4sf7VxyDLTaMJs2vuf1okulLyS52hkQ4
T6ANjxa0b99fzD1AkDSjEYCZEcU7jn+OTNn7umpah2Vci7jPnm+JqRoLIcCM7+vT
3V0FFahNbzf4Yt5smiv4NWswkakqIsxzYDiR+7sifL4joil5f73RnQP8Glsrc/3E
YNS7mcz3pcI/9p24HNiXTMrzB2r7vibzDNYuOPMiexsphN+M3N1fjsSBg31Scj1Z
6WJenLAS+YDXCpnYmgEBxeQEFND4Vdd0fjLth1KEC/Tnw47FoR0jW8WXdbn8tpRI
aNVXfG0GRT6UexmH+p08Q5emcHLANUqBEJCJOoBYzbhe04Y96mT2EveBWOCORgYq
Gi2sqVGOhlb2oO98OAC+66tL8mcCS0AXYhUT2xd2feaXs43ZAMIJHZK1FFCffTJi
Fybl8JnZ0sqM9xYvNOjRerleGirP7dHNQa/i/KunfF8wEvjUDllMXRPZPgPT4aiD
KxxE9ll60VPnz262MkiIikqJXuoAOK2vvyewNjyfkvnc97qic94YeSAf/x4VqKZ9
c1gUpo3+IGEs7BSTF8ZJXaZc9/g4RITL6ihmNkMDJBkemiMEpHnbC52WEPgUaijc
d0guuUg5+UlrvOPs22eG7qR//i5ErxMoVRsML1KTlk4rhTQy0ai4oBnLvEL7B3lC
1cjdyrs7DHGWKKo5jy/0p1rUYcK3hyHbDy5r6xdrL3Ze8xoaKdfYSNsZLRhZSI7O
wS7A6wct+VXigFYxwbEBFW7sdIW1GOZqX+Xc737PCLqW3ZrWhd3LHfnZ/2hA+JA7
5vISysDzy6QkmodAiJ/f2yVLetl0X8Ss/SVSnMp3fqy4AGXkaOiy6sbTbo6muzhc
10lgU1oy4qzWOnYvXcN+fQIyJCbtQjNq6twvzgm9nVsVvj2ipMAkWMmoiOaN1Yjg
o9F3BUN8QQiUhlGaANoVUepD0FHuo1KYZLCXkrWf8aG0nFLWyuleaga+GHQtkMFq
k8gQf5HrHErFmg9xRk88+OdaGuUqQsrVKEZXzllhn3AdATQw0OWIHH1zhyDsS/c2
SeiYUPIiFpixDH6AWfV+pC3bvMwjnM1dsnITaVEP6I0okqvU5i4qSynhaZguH6xB
2gJjvx5Km9ilSd6JTDlVfCE7Wp8+GDFvRPGXPita1jrrWVGmK01qLWlz7uhl1ZUi
uwvrxXsu4H4qwaTVPQzolw==
`protect END_PROTECTED
