`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nRvdulnbcumFITnMoIw9uaHnVcz8hYXiWFDZrZHMUctCyOL5TqOKyQtt1yhxSy/2
S57cbAfJFw0OgAa9Wa2vzZq4ht33/uRV6YX6TUz/fLN45TLZm2dtbFOXwLp4ONex
VPQrG2+544UGgKNORYFG6aH7QgoFJ1yGlHy49dAIAQxPj4QSGsvL6nVCm2d//Hlp
CzzQZThvgJ4lIgubNZUV6N3cfWv+CV56rc6t42nhAhpHyLHoC/l5JvGCOVQPvveM
8w9sWNFd8Kl//x+Gy+q4zHzurWPszJSYYL7PVywWpMpV7xuD+Y7/FLTPaXiHRqON
RSQ8T/YZ+sbEYDTpBi5edVMYzHuNLByEfRAjDqkKOT07nmdH0YycZZF3MZUutqaU
ayOGLUH3NvaeL10wIVdI8JW5iZpeXes87mNiAhNDRk8bN2xM4hTcG9a0OCwe12BW
VzNl1hntFXHegg5uMTHW2wv8Q3fELsUITz6F3JlI3Zdep1FcDqesEnaCGYF9GnJD
7ZzjAWfcFWtTvpgpmGcXWPOD3DAGy2jghTNx5TmW+Di88DYyqotPpbtA+YyMBrTS
77PsECFMjy0Fh0Rp8nhZ3Q==
`protect END_PROTECTED
