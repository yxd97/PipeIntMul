`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u8k6f+DCyAX/otY5DLGdQ0umE/xq8Z9yIwNKlyreVznEnax2oN9oQrsirAnOxlo6
tSw23qVspr2UuUYSPNUar4v3FPdUhBjCnWay2nA+Nthj/wwFAR/kMkEePO6IplJu
rrIbVVARNouo2zGUVWY/DuUj/zk/gHv9RZz75cY5TPdyksUGnq/Mkuqss13XCxt8
y7WxnY72ELOT9kT5JKmwuKPgDETWpCvQfZrgtSP65Mg7EnBc0DnJUzCUz5Ctl9hJ
p2Wdm8NcJ/WLKlEj1TeL2tzVIMhHTd06GwuB6W5qzJR0w3NsIs89Wu/KTboDAGa4
FiFvUB5hG0WdAjgzwAr28w062HemXPPDua5MWIVPAbF2KENuMliRvIl+DZps8Td6
gN1c1I5J3b88mSPF5Wbw44DFUlFrrCDrZhp9X3MeA6SSezD0XhhV0fdPXqmq9tZy
az+WHNWpkYKt3K4Aj7M7CFoz9O/xAKm8scjuwkLsVevQj0Jo+lFSDB8q1h8nD7Wq
JkQ4S7JN6exbZLcOIbWs+CptjXXb1bWdo7d2VgBTRBusKhBooqKxZyfyGyBocPCf
NnfboGfn127SfraIeBZmS/PugggcuThMYri84r++dYJoto5ktFeBZsdYoiR3/j4L
8CauaRB/T0AdPXVNTwOn3qLRoksfDPM/ZbriJAF0+gXkVY4zUCmPWG96l0SWq7pl
0Y8S9jRUAnjUdRsLb7aEckGJOADboIxhrrPIZRJu5IsbBUNaq1rb50WvsWXkwPuE
rEsafJqZ1kUmdDUKpIkARBL5CX4Ll7Wya9Iglc0fzf3gpli9+zIta887rUW/DBWd
pR8kRrOa06eY4A3BisWRfdnuWUL2l2rT73vGJ4fqMJ/n30QTaEZHlp2QZRDl9zbr
AfNF4nHaPY8RzZKiE7QfeaO/fyVcMYG5o8S1iAbtyZtp3UQGx9XnlPHZWzn8I3eR
og0ca0VsMLfGQRzSM+jSlbfAidFcSdoooP63i7o6lGo/0S+QJJplAiqyAfxObEMz
/n8/MbamqUVubpY8LQfYxqbgSpPTLJBH0qt89QtA+CdrmeznOW6Mv30/ExkXv1Yq
g/wifP6IYC8Lv9opCHN27r8Jngle8xD87Ki/FPgmA37ATJuTMIxSfyPVrUoki1QE
Lbv84T4iI5oORR8eIxkm/j0rrZ9GegW2XbhQ3V2x6uTahI0FNlyeFVOK+9s/JtxG
i/rJasV/C8ayhxWn/p7Tce9DWxkeOyAWKrQRyvIE+pTkm3bGVhb+66rLeRRLriBJ
6ruupUN3ihhR7tFi7XxnCKExsPlnl1bcMrZlS3EfpZIIGCJqh2qvZF6NQRgwmB6y
+n80LcNdiNhaQ7Yv/b40OThaMgpxuq446mBVZigqyJlwoyD9VCZFuZLAZqsZacFk
X/MhkSs/S/TDOmuYNJ6ZHhagAzC7mNIedMB6Ql/6BdW29kWMh3EijdX8o50c/pGz
94cc65kEI9ohzIIEwe/1TI1/jHipJljfOMsZ2b25m1/EvEJXX4CcdKPWihX9W/MS
Ggb4OBpOPxBg/hnJLAK4Vq/Hf40ZZkG5qFA+nYSCVDr+rJBwNpf76K8ytdono9wk
FNJ+Rwj+Jn2QXgewbbn+Hw+22ZP9Kyq+mFiKy9IcC3DJlSoL0i2P+0pPYC+Jv01y
UGJuSipKhiI2AdXyTYs915Oh79TgADppJ+icCOZ5L6vUKs13CCWv95lZoJ/aIU0j
3AmTPgLZgsBkZk6qOqTgGougZlM2FAG59qpGFG2bh7p0ZW4jORRyj2eOBanYISzl
q53PMPHbJibc0ZuCndwkuncO5ot+z0STQg7Gl9Ua7xnTMdxqFJUQBhkC5cl0nlR3
PX38EAfPbApEhPIbq6QdzYJejSjtJb/neWed4i2CJJIljem6EzNN5CAepToiwPv9
6iIEA85bXHvLvEujePfVpXd0tmvhoLn+2JsQW439CXz0hgxDj8pH8Z9fdcudhhC1
m4VXaWKBNUVbz8OJ5vbik58EUPflFTwsfazt7uR5kH85bDPcBUG0H7EjIQ29Ja5Z
W0LawBFvb4A25x2gGTVZBNaVz9d8OVsI90pWLGRRJFy6HTqzHXzNguZFI57H/Ues
VEJFJQO14Us8K5tBYlewhmo1nbPmvbW3rUyv9VPQ7OVCOHPXHay5mFCT4TR8VkOF
pUkBoPoNuOBCYr2mwI04eFevMEBHZNfACz4cg5yj+Htkaf6Ke/nG0OFJcH1iQCL8
q8vMRLLjyDdAIlIV8wTPsGkTb8wYJpNwnZq5SmrMoc9PlqSSjtfni4d1Dmxj3eQr
dW8s0fu66h7Wd6C3a0Xx05lOhdZpF/bw/LWTJ2GQoN5ranO4es1bIRQ1v66WyFST
E0yEaOj84+9znTyWUU2D+WOj6O4lvv6A4D5IR1smiESaAZZHELVkSpBJAESzmL7H
UDn5EkskZg6YkH0ZQvNYheMLCwsC8wsNl5MHzdKvyPG0w+T9fHcswIWD+SRCZe/y
BE6J5rDEa/y0ABm7uxk8NPP3Cua3wdgph2Jfl3Hj6mX8mBnQ89Kh/TR4j5uLv9IZ
4U9gE6digBphFlHHwUKFXuJHcNZ0NdJfLAfws0iQK0V6LFshDpxzMnRo4Jo9paJq
Q2tS1EuRC68dPAkgL9nUoW+BTAEkiI/kPFe/DO1x3RHvmWUFPCnMhP9MRsC2YbZr
7msyYNfNbvafVcfaUjHjb7iADsSJby9PoIGezpx8yCkRg/insyY3vjQ7K6UpYbl5
EBY6InqUQBGn1GHQpWNM7ZV0kVTYKTOHVvTEWbfVKlnQOqIJzHDtbu9zuIv1s3yT
msqUvMo1jl0j4xCL/OinP9nYEO2wn4lfFPKb0iUqESp+AzqM5JzYyqUzpltLHwfk
TmaF4XA0UtbNI21MzbebtEJg/p3haVeEOvbjRJ3WQA8Vd3ijuS5IYIkPVdT+Xtf5
9fQCvBcCbrYSXYCgSwphmWmEhlR9ljgruIaLWSIUbTeyMNcSAarNiyv0LfXvABOT
R4cH5EKjkzOHdhiN2BiTYg==
`protect END_PROTECTED
