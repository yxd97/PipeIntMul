`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YzsZP+4ZTI2HkGnRqbUnxYcxiH43l8CYc7hPRVQtqMH1b2hJ50hEOdVHPo2aUCs/
OLKlTQhEa+qTJm1oBAhkt0b4vVcsViEtEFItAMvKJrydMrgrRr1Hin2PpiohM1Qi
lwkPvq3J1zOauxYbevWeeuo75C+J6NLg74Qu05JN8KyUWk5Chn7NKyJjVTzMIcXi
BZx9c+B/NsazIfVe0hU+Ozi1r/2+4pu/7mrdEAhSHcssNsG2xP2D2h0Bv1aP4KXq
k3zFPbDPVL2UujfPkvb2RqdN2nYp6alZ3FPNENfoaFxpVID8n58FH5Q/U7TjiRz3
2Wvw/uKxD2baZccAxG01BQ==
`protect END_PROTECTED
