`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqJAlj2cQMewNVQHItsuDIYZX7v/pDKblk3+mg/drkmKfQxyUpONN1D1PoHZYGB4
THaN8/51srwrhOEFUuX+yvuhmlqQecvrQ3JjrZLsch2Z0kmqy5+6PDbJ17KPTQpW
AZcahWlBYSIB73joP9qjt9u2ZV91oCidIWeYiqCHKO9Vao5+g7YRkTZPPrDB35zT
7TyPGasr4Ng6RHFUwVlXa6lR7ZKMaMlD4X/7QUWvSKN6W9PuFbkdsa9gUI2ZLhk+
kxAgvZVKnb0t2dITB+Qh0UPN07fq6gf+SP2IlkazahpTe9OucNFQgtLp0GugXG1w
irlS1mhuIbtrZXFGlEOAIA==
`protect END_PROTECTED
