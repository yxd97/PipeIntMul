`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lBd+46p+ZK9PTR9cOUeKBM/JSKHPrTGoY4NVOzy/58/t/oiMvVw/7sHj+Xe2CMnq
5EiRxxWI8lwNWeDmscowIkxz11LqDAOpkPVpzROCh2IymfFkmjF2GtjQnYLI0LrH
3EdzleVafI6xhR/TwydTVx9c0mNyiEHSw0w1Kcg2EI3HN625fjiQ57TOkMiO77mV
3HPEL+sLGzkEqhT+ENmet1dy+4o2BmR07dJGLTQ7S5WkhIW61idAu2kwt6T2NP3s
HJPhP2xmSCyAzWnQ/G1dgppsJhvLMCBl6Z6kQURncdHK32ghvxPiWoyiseuwIFWU
QIrmpiSoVWLq7ikdTYK/xKiow83rwihGIJDPeSz2pO2FThII/7HkkwK7PFSC0dJ+
tnUKYYTt9Iw1+NjwYLz5WxNrj+aUHGWW7wXUS8IIMAXkTK/UqtF2nWia2mrHOURl
dtOkkOhP4UHUpO1sjN2sNfNx11HHEXoRdkIESYmb09K/GFdRc4kcsrYqDL4Z1Qj9
`protect END_PROTECTED
