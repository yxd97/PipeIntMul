`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kP9iBimAPEYB4HLyC5uvzzpyMrMRNzEODJRRggT8GZsK1YsUDaIrRTsHP0qHS8+c
ExpH9jS38EMH5fOaOrygT9C1P1rppZWlSqwAhsApBterRFrgyNInIH6N0pYgbSoM
jzM+JiSOZLa1A1Zc3q7wE783mWv/jJBHPQ4hFOkBXp9nhczWYQtbEe/GCDjFWALI
i9vvpc41/WJhv9CJSXxuLJZmrEQZQx6vj5Ag5H+Z40Cre9iGR+GpRkBai+I7baE6
MawrislnLxz+GLVi7X0zlPcWlZbTfyCdKsq5Wh83dEezvMkGheMMQz5uHxhA2dgZ
3t4enKosmmeSOYlNlStofCxSUSSULptfASyv8j3tW2aPSfq3qXwUh+omJwCsAvaj
U+UOPCBJ65Ml7gTc7kBOLmmRHnGNDGXNSrR2UUVBsIIgahP6tjOEMMHRn6LJ/TIA
6qotACwE/eUsGaUqBKj3P6SxPo61Sg7jgEfYTcS81S6XQGzU3GhzlsrupA9DeHSJ
qlqJxFK+tlyx3SKBkmDlAF45QfhBVMgMiYodWz6u1fY=
`protect END_PROTECTED
