`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AztpjDwm8bC2tRE5DWN0elabecmBkgjL0xxiIXhglkUK+Uv1qFHnnsiuYFShHMDQ
NAkae2vhVik5+6wf6M2W+4jaEvIvWBaK2s+YV+gCNRw0QQt12km+Q5/jMjhJ7MTT
a7uk4cGd4WLYoSuMpTp6+JRIRC6F4I94EIaBFpdW3w36gOLD4oY2syJv53pJMABr
hXGtv7cMMLgYshB06NMogr/U0BE6YTpraGStFHLiFZ9ZClS6TRPDFMx9aJKmrkD0
u5T2nrsjfPi2xQppnjl1q0TtJHhiGup/h4AChh3v9cnOdVuFN51f4KhfUPtOWJx9
BSl5eSIjbW2yqBpS0iEgTeClg8fhvUrDWLi642ewW0dYv2JvXBiIJ8U3UbT8bsat
0YV0eBMzH4Jnu2mtmz+UkBx7qct0x8gXBG6kmMTo8yWoTp+JpPE7PBu9Wsra/O+k
`protect END_PROTECTED
