`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXpLVJIB5KK2DvJybtK7PKLqZl5mEmtRqtXQG5j4po5JZnbuqBqAOa6yvDesr7L1
AmRV1vkaKz9uVPHEq0e1aF5vXLyho6AdQzrjlzcIgjY82cR52rge8R81oVzIOYX8
DpCzGPQLthf7UqiBb++WuIzDaqH9/Z1bai0QNWeqHGB/BWu/Rc/1Jj4RSe9wR6xF
j6beOSDjnfv319v4/UQWQTZED3UmGyhoaBUIxsD0uWRyW2DG0aiRx8BhyZlol9N/
AZQMZuh1QK22SW0HVIXtKEhZh9bKkODxRsD5AGj5Thod0IWV448Ad4SzWAAKicM/
1Hs9pXS3Xb7h/J7u0cAAdc3ikgNj+5HlvySc3jDC3fKk0gT7rRSo5RywvAUXJVcl
516/z/lFcZflv440gleGSh/voYFtKBy5CpY5craP/KLprH2lYysAjmQz8qQg1Z8E
`protect END_PROTECTED
