`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwZMC9HMkcbpLX6MOPi2z/K9hGydKfE2QR/DomB6Y0hoztuIAEZ3FM+lG6rCf7Tg
/O1VroRgr3yQ8ZVafZ/LohtCMDti5aGcCiyUbLIOyWC2fH0M+Lo/lleWQBy7Wiid
Hp14SiU3r/Jk5/NUxGJXG2Dcps2IF2HvfSgME61YmrUTA1RwV054+R1bJm29ujun
KyQYkSSfIetKOExvSlgXP6yHHR06tODfokOfT61/yRrHTxlVPIJXr3aXs+RtwgyE
qDn5ATCdnxtGe2kDpTT8oQ==
`protect END_PROTECTED
