`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5cAeQm6VVv9VaWBbEznqaGEO0CK6X0jNOxD7B4E/JCVW2ikG80nP7UOHMyiPHAg
bVWSI80NehzBC5IJEBfjfUv/0aniB3KIP73Dwk+sY4fSFPtKVvXIBgqo9akySwv1
6KUR0toxTb1aCPA5RFFsxymjMGrijN9nVbMB5xymKiboH3Ape/o+rTSxnH7Ceg+L
OEWdeFrCLTtmPi541NCrRvzluldwrdB7MYSeB/WvmtscYD0yGcUyHOG55xthZ57s
v+fRub+2DZ4sm235vPmuCKzJrszCqaj+qK66l9KHmaLNxZEp/q8xjxf9wlOY+IgY
kPDxXXT7YNCswD+MZWIFeJytFGGsUUcKrVyslNun6zuHZyfdTjSZcU74aqz2BDMe
OYL2JkRB6RrU0nFh21fTjYKl7zBlNt/fsV7i73JI9cDh98xeq0nUIFB9lLWMN11A
pvda1BVdTUNxQSS2SllAgwEO+Ctz0s6fTkHwo1coDokkrGzrr9JMktTwvq+ApE4V
P1irMI9p7owpC/a4Up72yGFKtXUuqdsjUdwmp5u0apF6ddpMxd5x+LqldYVKENDE
Va1GamYQTodnTDKi5rIymM0eEsb2Jj6YruZa0XJ2kY5BgIVstRntk4h1kwwBhv27
Kt68IrBc1V0xA8cBSYGF/nJSyde01XwXCG/M+gmk5rKZiYXgsmmBedAMYaj/HIe8
46VZXICZVwuZj+e7iq4Cdr3qNs2Hk9I4MmriHhRWJqnpILhrYzJMgWr062W3j9KE
zA12krp9PETO3zRf9eLvS/IcwfyUA98+ixODbXjUKnM6HGHgD60XlL8SPtHJA9WE
6w8PCBo2pJ2tJsiZslRuGtEGMLQJw6+sKTsKYRqV1WYWBu6cNYrY+FK4qrNfKMBK
oDBdZizoTqeZ3u7lo/69ziVr+XsINFZFlePnhE3OxKLYXfoM0+QJblq/yTrnQTYW
dJvRB5/Hn2UiZgJ1BBIoavSfFY9jvGKyycFmAQRThCuQXGaQRTOae/U80VupBk7y
tWB1Mt0Bdl0RXKIGwn+czDaQ6k731Jp/h6JX9ozJtE071qe3Zv9ma9MsJvDU18m8
mW52pC0ntBgu8YTmjfY+g1qfsUbXGPtktj7TsS339JacGUttILdbdWmnO10V2dBu
+q3T3KLCYFh5Fd45hSxFYRGrH+S+Dh/O6Lm3fqtDCyIXdt2mulB4rArVLr5JDfc3
etivqZHU9hCC7NPKDaGXLfEdCudZcHmMNjCZD2cqjuqrjIqfH1+WOgefgaSmuezo
ybIqzdp/EbFV/p4dOMMJLJMi0VgH1hHK8z9xvXIpGaYcvNVUKonzQdG+Dhf4mjRS
JdaIKCOM6ClX5oZgu+sSd4unh3wnuTIzhx3AlLmo5iOFOA2DRRfRCQruag/4oToq
ARWzSWwDHcQEnugjxRHCnTDUlfyinVm2zjm0hayl6/2LdErclX5K3jb31hO8W2Qj
fFacfvFt26AkHLlKpsCbtU2CXDRia4hZv6tybg0MOq9SwAZbFcCxBIwxOU1XehI5
qWYZgwUH7SQw0eXHWkYBdcDB/Vzvd4AnQiX17A7A0bgxNPa2del0UntggKKN6u2/
6bt+XZb05H28Qc8HSfG2xBKWU5NWEssPPtmgMRzTlLQPj4kpYXtfPZWz+BBFmGbz
6jcsKojO3DuVfEDPbP7w3yIDB/XNtwz8dB5j1cWjbEIbEXAoKD88SPh4FJfmPuoW
BXvxVpiiJmMluIcKfL711iw/vmM2cDbSsHeNb44io1C3t5XitzvVJlOLKVxUdyLh
/JBZtWlJ236fXWrouqKFzZpEGfkFy9NAiMpLQ68ItxVOsxou7iUArtSflfDUPD7t
0kjBnrMUrCBEB+lMMdLMrwP0cko3en/rCAb7YbHeW6IBZD19Nng1t9reoOcKccja
mqGqAqK3ivB6YZmaNdSxT/xqlCJ2wvXHZUeJEWOGGfOY3FlsiPhcSGe9cDCZKK0u
fOLyajxaN5lSzxernKfIjULzKmlKDW+mNY+PFwd8y37oNa5VbMIlY+Ubm3a2dy6q
0XDmbrhABwkPiz2w3FAD7Z437Tpt7VtuVOu5fi3JuzZu52q1tWLKhQe5qag+AH+w
F3rmU8WZ0mFy58HTsI4F6b1YlDCWGkIGO8g3tTXYOt1AJNEsL4xxoFBNR806BJiG
7s/9iuBmNsm8o0jxVwBtBeLjesdsjCz0m+D2skJakjUBu9vfcZ6YxPXY7Vs4gnHz
6KrPlldBO09Z/AxaktmYqna6A/dvamXQ7G77ajJAwDEahOx5mu4ijU9v1hyirytu
GBkJ/QqA/Bphi3TpI6bpBFXWm13B3ofsxBBd031qpBTjiZM6oVPwPlYORlasrb6t
sh2PnfZshl1mDMME4EV8kyUAmxudgokcCWHPLDZHAKYtGSbUJrTDDi332agFM3XW
Y1PgTQETddDWCXY+WA+tD6UJSgEwBh+QLU/ueekwz2730AclMzQXia/lzhBHtjl+
wWNZ8RReTmK/yis1sFYDrtJ8+8UboYygCXEO+uOHUA44HwjVYQQ3fOfX6OmKcaDD
PumEAkPyUX71SSAxkrbFJKtEstfgU0Ec7dWJz/AudimV9LZV3WSCwzddCBbafOIo
u+LWvsVvnydxawiiV0aFRI/DpM+5xONP3+Ak3zz1DJ91TbpZKcX8hkBj/cisx0jw
7/MsogfWupRYsetY44yNHkdykhqIm51lFFGWGTsJwrSYBtLFDeW9raEqbcdrNZ4s
6afOTG/R1LNbabPdPlH2V9JvlSdO3ZNtXz/qt59IhLlfzCbT3/yBDIBVW9sttgpF
advmz4XE+OrwmtKM2yfzSX18C4ONhj8yaxUFp9hgGpszIEp53H9CbgL3R5D68uXw
um9RgVRoxen7JrdneVzARXtTwOpG1N6gDr9dsLVipYslkRX8uEWr4GNX/j0C+b0o
l7FPSvkBfqOZ34Dmj6tyuarPxjhBDdvhuPfAz6LHXyMip6klrRvLuKU6ppzl06rd
I5CkAhKB4CE8OKNcvnta7MQqAqr/XT6GdMoxwqCF6AbqkpfZL+0sSP+KHLWjU7jq
TfvVJ7JTVxgxKqU1eYOYlmtVTykDyL5FYyncaaqE5BYTK7EZOyWw8M/klvtwjV+Z
Z6Inw6CcE/sIo/NxqCwcjnapgd39Q1V0eQD5UEAxjGx1Qy27gY4aY3nNEOHlCEss
1mLCUp45GaMV/ZR/Xlzuh4MBgCFpD7f5bF6XAs8RYe2uA61hxUmh9rdJcnYkGany
I3jf120hArypBYlYulZwhO/E51dEBPAcbMAkUERNNWmUy/OF7RrZFXXGwEaVRsow
8U/FJLnM2EthaJTA4j8f1JZWXUPb0vmjIYYbYLiPjKuooB3lWaINQLAcXOzD1BL8
k1Zx5oFdQ5GCVO6trOJ1lifBWAZBhX8Ta3FeOgroilgAGsM5WGcra34SLfTwHhyL
hx8YtGXxUFrX9EkLDz55Pcoc4IQ4TVkSbNIkiZj3+Ccrd1yx3WB+2kfaPhZJfyOk
KXOsu8QaklgKpRH7nTx7cQmkBLFTb2KdDhH9qzbNdwzs5MegDkgpoHarbIG5LDZq
m3m+7ZRxHeNFEw63c/P9VBgRPBycFH99WAB/axgwQDBgyD1FHoMQb+F6OuRU9n7c
E0yajjyeTJ83aqoOgmAC9owd8+Aj1twROeveZSjzP7K8hQ6YYgWyE2Ssqpt8nd8f
elFdA8k1fP14kGCWNeNd0BzfOSG1iTdQ1QPuWJiqdDDTXdXrBzKFRRLokB7NtlAI
tCjlSmwWxgiR+WbzDKPmx1lb4uKgQyTE0tptW2+UWRxIBATwwedKV0oJLj4mk5O/
YFwqBIVofq9HkNtWTpt77JCXw3iFUUkEOR8N1HFwlikZN5E9RiqrN9s8Ruk25acQ
7JCNw96RrREZ5xJaHYZkRU0W09FcqAVhjTp60hWYEiPcGHXbhFajhNqbuVUnGIJ1
dP2mdrQf/OqXjTyzDI8xFYYSftfepj8KXiTDcJxrLNEVE/D8lpQyGGsIWYDmoqcQ
fip/Lg2jOrWHRVPNc06EQSoQ3j4BsG+VtN52TIjHpHV0VWVZHst+JaWgza8vfHvi
7T+M5i2PV1y/RZJKFyWS+97CF7P3E2Ms9jgmrKF+eG4xzzOgTKsBJU8+/K2YmpJj
4Pmh+UDeTi9L7ZeUr/ui/Aq4wFUTv8Qgl3yrR+TdJLLxARF+mUK9NMiKl53gLC3g
ro228bLmpig4XeWgqeb/qIscp0JHrj/9hXyX331o+F2QXIIN2m9Zb73hG50lvR6w
jnxFR6FcxBjDO2tI3UNv369z+5TwO9LTCQcKSNGyH/qKagjQhPSHt+bAOtgKijza
Wu5mitss4RYXzHS7ttWXAmlpoB+IZyKlaJzE2wIJ8fOv+khez09GS1kPVGd4m3vW
s42EySrcHltA0PKkf3cl3LsWIvDk4y0yVcVGhM2R7jwUrcASXPe617jwMoKkX/2H
ZxPqidgxQtU5Ve+omZHi8lQyBuC+i8hBkDd7jQbLiwsWPoWvvyaIchKQtUfeKFOk
VU1va9ibZn0iKwaO3XFcihQk2PT5uzjM6bkS1JmIQ1e76PcLvdYFVACAOJYlEXGd
u2kT058qqDodxWVmnx6tlKXUvAlrkS83r1T8EkHhIY0oeu/L+02gZDxvQqfsh1Pt
BWin+TbOB/Zr9xVNf3TVNcCIuBelAk46Xb3Q6/C4mtyo0luUcrGy2hSEeL5Lgz/V
IbxsGN6Zq2ecG1RTi5ZI9vURS3Hi6LoMytz4WSd/kjfeNzoTNTwTBhcscHhs6IqZ
ef8cxbbeL8z2Ubd2kkaXQw==
`protect END_PROTECTED
