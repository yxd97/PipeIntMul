`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZNynXFCFcp4kp1WZuMNs2+V1ibdLvYkvZdngAGVsX/hwIIzGcdkAYHapIJi4541Z
YNnmm59cceb/tod1Bh3ogh6bHVmVXPzIVPoRxeH8VlQ52MTKc0id22dDJaxgHLHn
VZky5vN0eOFJB+skXB+qtYGNHkcVPmGx21PkQ5SlZ7LnwJKPolu6Y7k0taWBiLiy
C8nSIyXHuxhs7bjyKFnt1Fn0mjx0C26cmrDkiWycDlQlQgbKyM4mtyGJiBAjc2AC
DtTSzqvlCdgUAFXmxhlMcNf9iD1ooCd1HbkTQPaAonwaJyIIQy2bLgWM0was87s6
gk3GR6UZkM0pg0o41UNnp0SJAM20yJMe3u+0rtsF5TQqp+4RS0DnzwP/imnSaB5O
SutkeAcE3mzhk+RDUlzZaWUS6YDY4nL8nUBrB04P6tRMXh6snuAY8gvOV/57rup3
Ab2RG+DjiOo3eooBc+TWR2FboLvvuIHwRWpZBO6QFoQp75mt51KzkeHzykD4AiF+
beEpu3UKB7Nl1k6gPqNYAYWwFiqVxjxl8YuVtCZqMipT5FSoRipo2P4uIRpOx7jQ
bkVonjwulhsjU48+dfFqXyCo1gJuU/+Bo8M5EtXzx/dHFJrxV+AgETX8ehQH4Yrf
MePIbVI5E/xvf7N72q5mapeef+G7MtYPLRrzFPf3g2nLWff4ApdGTA+IhkBa6Awd
2MHnkaJIOgEGQVU9HAirGpczyKWtLVWIpNi5GwAQFzsNuNg5LtTHw1fwZWDOuYTq
QMCI8Ok7VzuXE9o+DZINxF5x8hQpv5WUU9owiVIvCauiuI1IcfbIlGtcdVrwXBy1
W0RZCPswmjlyhwwEnrZ+TaeG8PgjCIoVFd0C8ejB8u+mPrpmRGqrR1iwDXPpTFMy
wGVMVPcgGdgDpWgfOukV3GOdTAyLAGNcfTnlwMXQNa2wdkSh2JO7NPnj5l6fbSx1
4rTFQ1QgPchmuOG5ZaxgOBsQqzSiNuEpCh/Uxx1QSvelwf0s25wsf28opZ3NZCk4
vyZWIvPj5fbhi+vqgjg8tmwjdnD6XW4kaQ2hD9JjDBMElB11poNlJPx3lGKjpTeV
uX6nfrGzkEHuE0BkWGljMSUyB7lIv2cqoPbLckTx8EfaylZFS8tQhidJYLkG0SQf
RVZIYOlxmvhSbgYfD8Mde/6sOFKHiY49ikREs0TzgRHlNnjfCmmcAzKCZOtC+XwC
O5yLAmXACp28ZOPcPqNCLic5ArbZTiZ2iV4MaC6yw3hXLXSb4SysZxRqlxyv9xR6
3JWNT25RAa9h481yvkHhkyoHjqPh3/+MVCgbtRg0i8lG5qaYXp+hKBzJVbtISIdq
syj4hIXVZro25SDP7VBGj5I54XnaUv5kbAaYhQvgFWVzDVs4gxYIRwXOjDfs39e8
XrMWm4WkSHygUkHtZfm2uA==
`protect END_PROTECTED
