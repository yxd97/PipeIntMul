`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1MmcsMBd/lp4EXroCyN9tBWs7PW5WL07gZW0PzNsVMu/1ztGD6iNAPq0nNxV18XS
pgVRCWzWrc0n5+hgc1pi03xV88Q+LTXdxWS0ipMs0rk75B/hRUQ1dqMdX1g7KSkR
hu9fKkGH/r1R4cik7jXvUBmioD+rpsGBlLqq7zHU4LZAYCZ2qA6PUdUT02RgLrTR
EzhHs83EOBf7eHhYrXsgNTy5TnJdK1wISzWNi9d4586CCN+yAIGAi3CoS1eC6ZqA
USlYM0VPlw3jjEijMe3BicUjOb3r0r8b8NPyC6dYDfbHntHaZ1uST2Grx8p2/nzF
sYMWr3nchPz4JVdqSp/dxvPTRrzi+fgmcGSryygbnKuiQDCUPKiuBIpv5IfpEZpM
S0MAwYhqvv+KsjrE+72bTHVpS7XwHnRKIz2PDSDhgYwocalAEday964i+MYIYy3l
`protect END_PROTECTED
