`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UAv+MMB0M2V5Uos1AkHeCWSzzK8ZnJpZ8anqFIkdCNfzM23S6fZDFYM10yxqeE/+
WsnIbOL6VQpgAlXWUYDAyC1t0QbvzXkaFYLtata4Ulv0KEqIDQma4itcJkBZ1rXs
OpJN9CXLkFmIxTxCkY2KW8fm4oQdAyL7hcs/xjuVtaq2RPL8haMP+oQxGBrqvB9J
B64+430bkGGOmoPDbkystmGLHZy26JCa85evlcfT77nP34yYygc+SAgDuPUuFcnA
ysaIeMhji4p5hmHpgDWjXmlgblE6hGoZqHI0XvCmFrmqOrodG2N7+STtqj/26jzW
eoQr1UQJ7mLXpbUpMB9VEYq1DcO4yphMTCdexB2JH5yPdot8yOHMG7YA5soO1fIZ
Cm7vmvN2vDLsUntVLkEw1am0g604RsO80ovTY4nWaiIx8zdAxm4pZ0mKRqrO3584
s/4ALbtbz7VxTWMowCz/16gnAFOFgA4c3RqCVK1frWx/lRifOjAnbw0IL1u7Pk92
FgIX45pv7VH2FkdYE74NiE7aVw/w3YhHf47H5I1feolPaakJMBCv9sFp1U4igf6N
`protect END_PROTECTED
