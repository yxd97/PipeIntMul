`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8xbwBOhQvqspHSNwHTTHUF+3k/tJxJhG/1PIOgjJGS8X9/jsOUc/rdKuMsBTkWUd
NT5qexUkE2H4aajGqVX/5Vy2/xBDaUN3d71vhbMfYROrVAjsr1WaIUJjS91b6mZN
a8D8k1xy6bqr/m4Yu03mK1QqAUcRzbFXU+HMSYKsJZIqAVjYSEgqtYL9tmsG3Olu
DkWAb5x/PycUP28dmDcHggZmypTNnXehHJi8Q6bRzKEg07xeNSTlKF99DIfYhvZx
JINl0UiRf6tKr6aLVjUcy5g80DmqM5sFnIod1VMm+HVcHfkbDoL5ZMh3bCVgbnew
DgexhqmUEi/C6drtOtHg9uarmVMkqVo2Y0RbZ0+iQ2udFXwEmUZvPTcKBIBQQiAL
m3//IX9B+92+k7b0ab47Tdm8tNc1lqfAKBvHvOINvzcBKf0D1H5IeY/jSETEQWeP
aNJGrSGeJKUvFvzJqXujvLNDYAspe5yMkx0e+2uXrolfI67X0QL4HIwp8oqYaCV2
`protect END_PROTECTED
