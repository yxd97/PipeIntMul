`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P0Wpn/0Eu1liBdv6NFFZcuLpSG50uIu9pnnaz5w2mevXD/o9RzJQDYf6O2PE2V1z
p6IyPpKNmfVbp4yRzNocOU1vZp3AD+tuxb5k/DbekcKDy+hWF0IxODH4duFtDrwZ
l69tu9H++HNzyik0cl0KLmcYpzQ6cfMwvSVn56l3paIa6Z5auYG4kaaIRCy/ut2p
FXTEk1bmR9Kp/uSgIL5K3xfS8YHi3D3JqzV8zyVUY+/GIM4Xk9wkywenkURMQjL3
c+nCcyfGRA9LF3gguq0F3hPuotDnPM7nDs6Jbke/sII2RC6/0IKvZkKIM/DPvGaT
TkvAWNIOqPb/KlNS9fHRr37TrqAqzBTPcvwwv+xXij/JbQfDjEGo6Nm4XyqKkzmt
kJUbUHJt4QT7umRMskmKkGnrqrWQxBsgFhasVVZL/7Q7HZZU6jzu9ytxvaiR2T0t
6Dgg5+D7icSJk18/zLrWAhN9AKvuaVgOZfsItUdl5LOnazx1joRab8f7ZjC/k4+1
mogXvSyIDetcy8x5TjzPigsQmRjmzG91b1dufZi0i2QMhLN74ODQmhbHPtk69Fhe
7ZWxEoAcQf2wxANnggDzp8VCkYfiMNwZoildX8tpv2vE3oLM7LG5xLEiZ2Zn/f1b
m83EEfhde2AHiGVTbyfx4E7I0OMGlW7a4F/Ok6OclWGsWAudMXa+ZmNJWt3qklMg
Mjd/C9fg6FRZE3pBXOBUpg16zMrh36XcGXfqwT03Iagz5UnZ2JP5gM0bJmBW2LyS
a7raq17M4Q2RU75XttfB7WHulGhBxvzGjlHcgfidlkxhpCTZcaBLvurlK2RPrd8i
49fNny/jGTgW3hftF5VcHpdfSwO6XX64Wz8uvFt3a8ln6E3zliS6YqH1+iINHCN7
MVQn6H5Rwi/iSHXrj+RbGRigR4IjdOpH46wT6iRz3sLFCjOiXUmtd00M5ldeOHMl
grpKoEcroD1nSUfNHOpJCLePt5AQD/iZQOtKgx/y3OYBT5r5npQQSc4A7Vx4+R73
gRIe+YO47Zy/YNgd0J55mJkIxZg6EN7KZqrQk3aNld/6U8gT/syoANeDOcYtFcoP
V8/5o7zEyp9BgFuUq27qFXdXvNb0meEfx4p3tM60n2s2WuAUXcv7FPC+iLUsBEdy
LPDcwGAVgXiOVd08tsCx1NFey3EexsmWSGupVrjrqAZeq10zECrykjt+WoXE6xZ4
YGEhRBDBHCfctnNPrN/m5IMD0XxORdSEF5e7Js37J58=
`protect END_PROTECTED
