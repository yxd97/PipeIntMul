`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TmC5mB52OLwJpBxPJHxFTixjDCluTk2wQsCcXpMI6XMAcKFWOKyCqohHRLYktXGs
c7NeSfMYlFfr5VjmG6Gl75R8Vxp8dEVtoSFMMjh8WN7QD/kSizOK3jjBmlSErsON
BXAT+PNDUVy92ByhXdo224beLVeXG2pwN1vMGWNasfnv+BYL4HzA9e9P/1Z/z8J9
Y4fR2c7NFFPssRZwN6SP5MC035b5v06jRRksD1t7YH7RiNh2iT4yQslp4nEYq0tz
`protect END_PROTECTED
