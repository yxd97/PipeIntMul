`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oAqmmtglBiRIz64uX0hjIKvV/DIsSABD6BssCjqlxtR7rWY4o6HrvDV1x6wnPFuF
xHBicL+e1TQo4S2PirOXkO6u8mBtwMN97D5dChg+2Y5wKWAEt7O1/YvNu64wdjD3
CoXSAYjSbxGTxuuulaRYoZ5Cg++MY+AFw4tPg8ZPaRYZgAoi7Hg8jkX1lr8hFUkx
pVqzCfJ0kJsEoHKhNPdigkCzUez3mJxzQAYz0NHVrwAWkV2hSOL+eNP+9O3ptXjQ
jGh9S7kN5zGS96kPgJtbPBS3U37BmSk7WTEmKSP72RQxU3FSz2X2pCM9XvGfCO0I
a79HD37ieVjgLB41rnXvO9/fnBznX6R3r+amgqmg3h7wvVAlJKymgdteRArnWDiA
cJZRBta7746LcHDUEB2SsD6am0PfeBatVineCyAQXuBlrzUE4SHg/nBaHjeyPBvq
NRPOPrX2Nj3G5NNIMHLUSkx34Ktf9p/eXxy56Wnnz9w=
`protect END_PROTECTED
