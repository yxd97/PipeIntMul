`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vhZZjmyHI4t8l0NgdlmIXujbSOGRd4cieO6HWH1LVhA03ZuLYFo5/RMTUdt/Mpgw
/TZNjjm3CawyS5UxBBdbGJaTjal5nk1ys5or6JhO8kTnNUh6T3OvV3CgoArxCLKY
U0NfDJ+K4VHdC1zwTLiD8qI3K75eYo7FF/uYYGjBvwNwin6rr7M2AIcpiUTwG9z9
DeRIVi49ZZNH4Ykz+MzwLFWHJutnHp7Na6sXJtt+fRaPNcuU4Ns1VajjqCuH3qZv
fCUdzjvYWbqHXNzKjDH5qGVMqySKM3OKpeo8pHqHFlq4uA6MGQxEaGfNfAKXNhrS
qABuaeLhxD5RtbIWEYy4gsYeTdGPmqpzg5zO/S+ygY7+UWsZ/yjIi3pFAhJbW8XU
mTldz2/RM0UeznFaZ2FQgLeY5GLPUkwoOrkyaKxZW5+5Jvh3NsQXArZhEDC6wqDk
/Ae9Bxi89+zgsShzv77QEevEdlJplsLGUBuUwawK+6i8lucjSQFHdnq2hl/fUSM4
/xbzcREKo5LaWkd4AMx0ueLxujx8fLuC/85jX56TqIF81XezWeelmNIqKrHdta3e
pRYeoFTeWIXcXTYluNRzfiDUmVjeBcpua+h4UIiqalRLoX8xDbe2P9UyUjCOOp89
QLFF3/jTsGyK1LvQM0h5WE+DX+PDAkNux/s3oH28r8VvyyRBC3YIBXHiNZMxJKT4
`protect END_PROTECTED
