`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ekBuEE5Y0riUCoeWylVQSe2oxheXF3hU1xxgLwjTQpm6lK2k8LXr0ZQnYmkieHNF
NxEXXNCag/8DV+U3PECyXvog9RycYwYa8z/iJQnn6tGVSIYbm0nQ+xm4fZN+9tWY
BX7vGe3QtYHOlP0qu1pqLqu01Ko3Rf5K8V94qFYs46i2KpW48jLyXiBVeyQHsBEG
6Ss8nievGBXFPNNKyMq/kgzVCg37RdIZLUz5qsAtdigGQEHpmB+NiuKloZc/p+hW
ZWknbNxEfGfKVuiJjtr1Oqbh7tT3yZVtvVixgWsT0H+8cLKhbQtlP2y3VZMLf1Uu
jfohOuKCJnrIpBoB2e6xgT+9+FFLwMKYl2IPGQFyKls=
`protect END_PROTECTED
