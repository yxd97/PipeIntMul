`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xmjC2G9ykKqa5eIKKT47x218yfaAUx0s2+bwb+lSj//1MECNIr/IcPW6fHfqhrf
y+WTjTWdzZ+jygjEG63j85ApSkTMQqW5ABCRp+QN/VjBacNUibV5vV14J34C2Qpk
5ZyHakjcgBHvT0U/k16heIF4I2EOHSqazgdDw70tcghqST6qTV9h8J0JcB940Cjr
fmNzObDMMQjqMCiJ9b7kKQ4zkciAXAmuOYzgVlQSdzY53AdcMjQuG42Oj4AcMj+s
wKtQ59duJW8iQuSZibT8tzmSi8MKSaapKnopKr6aL2jzoP4SmBAbFbFYTi6GffHP
3LsiBg+KKI7pRQY4v3mqQbkXXQeRzLmpIpw+ULTTndJc/n0FuRRHEeKJhcnFb7Ks
rQ9KcK33BmdOB2ybCkAge5ITRA9yfbL0pY83uyQXi29AJlR6s7qsiB+iQveIfEqn
ZL7+yxKxKFr+l9ua1ue3Ral1P2Zm9/c4vBYjh/i99kmioeviLaPC6o29CnG4X9vB
ZUkiK8BJaARwa5h3TeWhTzl8QOkckwjJj0BhzYltZw4JcNH3VhahPRJEocN4aCLF
69RcFCTu4h6LLQYCWtuYJA==
`protect END_PROTECTED
