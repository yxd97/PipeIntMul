`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMQ5Qc60bJsasVy6fOLLBSsuxa4ZJ8yrrkiyjMR9hbCX7LqBmS+8sQSXpdjvzERa
xMtix04hxXEk59OteQAbEmyWkkQrJ5/bRKkcDzCUOgoQpoJusb3uaEHTRNZ53uKq
AS2J7IaKebvilhXj6qgDy65t8Hyq5vwnV/3QN4MkpJbfmZ3rqZE1TbEARP1Y6hLv
pZZ55b+CAxyLzTyC/BsXTGRwOaFhze5mUV+dAuVEm3D0wf3XtF/1ncdqnRjnGg9U
i4UYqsoF5/OXYPGHcQOTo56651TKQgsZ7tJbfmlfQ6ojFFbWPaSeBCJYidhqtGGk
MLx7ft167CaDXYH3lAuHQfRAkUIlkffJhMXlA3YtbIWrXJKj1CJIFkbbgAir2O2b
9eQ8ui8NjgmlnZbM/sIzTzx07ApnE5i05nE8AJeiy8aXfGs09rOIWKjD7Tt8eRuv
A5TNZjc9hki4Cxg12chafQ==
`protect END_PROTECTED
