`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GB2PYRqzWT3MkV/eaXlpgjYnlliC+CW5GYXlrzZ5GuEyFmncBNNjgc1SCVE6kJGv
sLOcUGdlGCd9cGFsuN5kUrltjGzDtYESXOI0D+vjHzKsQPjZv0Bm5wHM2jLeiVu/
y++QtUrRPciYf0b4avE6eThKG9kZHoycIq8IfOcY+UfgvL7+BfT7ZCDQ8jhH0EDE
quz3Dka8Ruj+YMYGsKD0FKLJ44tEP/ZRKEYee5oPBJ496o2Psa0RV4RehyXqu/nu
Oe6WYgJibEXdyf/vW+hNUzlI7CUopJY3j+hheyoDmvZfV3nd7iQPJ4sQZhVPtwrN
ExoiHflZEmGlGf9DahjtUlOO3TE1dZxi7WMlpKvtNM1Dgp8ZkKFWThnCHxBqhCcD
pzoXSuQZM29dBBDLYf9fB5pnttnsGNdpoDL/ey9gt41V89X9fk0MromKS4WyxH31
BmduhjSpG4uEF0K0wSSsjg/zmBeps9E6W6kzU8W1bARqbtkwhZ9doan9qUlJ4v2r
rtmjYCJ1FyziO4Z36mmpYGZn+rOLdT8mtPEhour8+fJx+Yr4FVPPbzyY5JO89S9g
qGwyx++PPjAwayoBvq9wqxEoXuPqXOjdZwkZp4Ef4uiREvlGk0O5ETEc3JDrEk9v
wNvq1u0X2ewTguhOLO5fh8eZxF91QrN0PTmOPQzIvbxfhpX+WFWG5nVKhpoTINdu
1oJ+gkv+kUdFQFdBt8Tehd+gBlv4hZj/eag0kRJerxWgIKP5QRHT58h3MPOPCABD
jeMrDcSp0ZJ0GkvzTETH6Q==
`protect END_PROTECTED
