`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CqaulBeSWZbENe29r7WCt57M9EhYaH6s2w30dIWYF7+i0U0lkAqqvVQyUJXl3ArD
Z/cnt1m2je6MK+xCeN7CxZjhkFMU8Fn3EMUwfgq30nSM34KdPGAi+rVmu5zrPBOV
0KWDDzcgYIx1IAQZOeN2Sso7UskwSnA87cVjN/zen/vEYE3RFxGr2qDZIEoEDlc6
xR3wgjRuU77ZUYSaQqJg2LBrgK5a1Ikame0V56wamsU2JJcp6rKMOe7uJVNWdoqg
DhK3r7gavo3TQusuxKfmL+mVWFSOg0TQnZZJxT/1y32RMacW9vJoOvo0BYGVCZs7
+zgWeng/rw5CR/qdiXl7mdJHqqvl1gqEHJJjvYTtRB0Ijw2GfdLaUbeD+YjIcIBS
Pem2GNPeMbk42dGKDQIGbEjSmmFkbaiZ+SkncSh5rtypQr3KNZAXLlncP6186Sh8
Aq3v3/PNe+YbpGCLfgMo66Kq5c5hN9+cvL43hz46ltUL2HvANvUmt4YdluyvCIlA
5azOuTUF8rtG4VQtYAvoGCwInHsA3uEApyEny+B/Idd0teQZNfpbsm2u+yL04iMo
xTs4BUMERF0uiTQ/hFEWCtj5k5z5r6xxJ1/aYz5bumZ4N/Vs36XptoklBwj+YgXj
IWYsmIslxfqlQ3hkbjgwZWT4RhYNSrmUcYGOiH2uUKxNF0GMy9h2ltFitO1ufNON
`protect END_PROTECTED
