`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HfVQr0Y3ChNaBU1hSPfJ0is+s+lBpdUEq9P6NlOQm5y7nYtlU2oNqOLyBgI+jDte
tHDvDd31ngkPfF3ZR3o+YynpOiNP+g4OjPVuxMzdjtLx6P4DUhWThKDJh+0bqemy
ZdvKhXrSl2r4DixU0KdIG+f5DII3hlsG6KpVoyWSua6UTg6laDzQQWxGbkx0PH6Q
bI+O73BoKcegURjJRjPkRw7oHeMsZwxXODPvTCl/n2De8IN8w9y5LCQvNRPGPIyX
zi7DLxYXPdM8txeGR+4PhHSU33uqQPW2bP21b2YX/ZhxO5p5zFu32h1bWxD1PB99
BmwWcJk8fK6EqBIDije0eFwzmO587EBtGmfjRuW6QSAtaOONOHCtEmrkp0NBsYgP
jmF1RW5qpCIK0s3QW7PbHswV/Rcs+sa3KjQtNmDm2RsaNr3q6OHg4BjtwI13FUUs
ChrurYlXwo6q02+NfX3+IdpWuQZs+PyrWhctF43uFvI4SxGMYKbmJYIKuiddPw7V
AvugwHPXFAVAaYCB5+kEgcHtHedxoVY8NDzeBe8AvKmlGHhHUQ8UO9BFEsX9YzxC
gCtNwHozq+uWG2w7up7p5/V4D67v/kmXh1cuSqkNp9eqfXfPy0wuy679+G1v/7Js
+pJAqGb/7pjCuYFeu53oMTmL4iwagRzmtNNazKWoIHWHtyWt67CMkwER+eCCS1vJ
15xySyRivbaT0JGxoRMlqyfvrXaFAu1zGQ+jxMsNMcgajS/sfx/kojQV/ugTahQX
YpTGBOhLHZTiQmCQL8WtL1B9s3D7G57uV0RkzzU1Fm5Nicbx3eU3qVrOIMiRu0h2
WU33U681XUmigeSa6ROLNZ8usxwGxF02wuFBPeQSQIY7i2ZmZ74razRnzRcTY3fl
HdoANils0oo1uIZexpVIfPhDqt24gVb4joe027L+QBpOTViT8pBU1MKlw0mFOo/l
nGcQMJstybkApO4Uli1J4OLk/H7qunv7WmCjCx9qkxMzP5btzl49piijj1Xw7/vu
zOi2tVlLlu0KxbuqnTl8tRAB1aU8xjkxpmhn9LwE7Y81kXp2gs3KH0YXCry2M9kU
WmmbitBAkGDW1VuomjHXlv8EKZnsDlJlsUNiQ7xF5L/YiNdneFtsH042hpgOXaDf
O56Q8ijmfJoZWR3E59/EJ0uGOi4ziheCmM2vctx7vjPDnrtDG0cQrndJPuabvEPD
QQbovsQ4+dgeri9Snh+W7Hz/kI3SYI0IIoy823bND+k+KtzWOyiMQkXkGGWEw4Om
sxa4g0lXI9rkbakiJ9+PBsHu3PMUQarI5JpGwUTrZSgZAY4giogBjG1/4eLAkBA+
6NXGnm+mAR5GPy2mjExDHoX6JbmygJF4FFgfgSpxms8fQIWGO9jkOJg3/VNAypmH
axyV216iR7/BY6uXfA5p6bJHZr4ZNyh39wxYQKdoty5/ntM6urcNa8ZEcSHd29A3
Oa9SShJWfS9PE+cCj5WWbV4bWjPxXGFBe/9cOrdsX1Z0Rue2HjZLQYeTjmkWeGPz
Sr8Z8vdCZYLo7LAsAxovuDUBpSpa2N1111Bk4EqrqId/rZCzXjeTWhYeQYj0aNRd
nL87k9DiWyTrvjOJATIUuOwqHqfvxEoIw6HceXChGG4KVxFWKeaiDgoYTwyvQ71q
rFxjNfoZKZ+rWcTWTCOCJuZ+/t7TXOUCrigPfUydiBp1sRXQjF4NZXBhLC1gRUmR
IJIrz7DwsYARNuwYfU+cgtf045hjZwbpZPSOSETfjf/vTWTZkCPL/9drgMko2KaT
FiYx5SszLr6vSbvYAoMvnyX71828txie5Bra/ft+o3qZjBuHy+AbnXi9lMpLlx96
U6wESCLDmSzfE2V9K09qjowPysPOvTYE0hSdB+PaQKgw3iE4lunS88IoghT+PTnz
X3fJybkDlQ2hkLS5PRv01iLdXXDohOtZUEv/OXruKQBbJsjoFiQAcoNEPkOetFsa
IvprS4s+nyZVwCLnokhYXiz/KrFiTG01ucXNEIA+G0dDkOmHuXSMO3xD80yWHvl+
tWbepu/nrxgBvi/F9O7I+VXG9lxPnHeWvSYEonE6zj4ngZ1Y+KcvCLL5sb9IhVFu
6znJJzFtQA7SfUqG2Y28tEJSgq9Yv4TgU4KyIvL7pMLqOr+GddLFcA1GSLe3lyYU
hy3iQANoYoDtQheqRCoNI697sVdCv5KNu/iMdGU2W7vOq3enKqFkGokqdebGYjV2
TPpOrWfy8idTHCMcwYtDcgkPefeelmQUns1/Imsgao253naq/NpwCazKhuPfDW80
eisL/w87WtCcgiW/JqqAhrFhzkrgs6girsSvMMhPPATzQK9WNzdJHJ5pNSfw9gTy
bbsFvJePugVilBhLcVxMd3pUIFgylnaR7Jrg09aNegaQGSHdRYrHQ82/n82dpYTC
TWL2DNmNnUILCIObKqc9xyh6p1s8j+JBOm3DJKT38xvI3BEUVxMYFq9dsrk0wYRs
bQ+kgZ/DeCbiUsU6IJ1GykBH+JveUfa0ECwp1OH7ZHtRbVtiSJwti1iSOdswYCne
Rb5zmkX07Ca1x5XJyJnpNhqClfTlLMDCAB0tHMpSgP73RQ+HmTRn68PnzvGJPlp6
`protect END_PROTECTED
