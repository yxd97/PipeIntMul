`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2PqhpUyLYC2CQxL678c8w41Lk/MQe6cKu8ss/U7aO/c6CPXNd80+o1Uhj/gYp9w4
g8RtIdis/ebq5VwDOMmaQm73r+xBQLyjxCKefs8P/tc8ux1H0TZJS85dX4LgSiVJ
qq2QgVOVqQgAOSruy5oy11cJtBvacjPuiA1dC0+6LRHvoW70r0Xn+JK76j8+A502
dhUEsF7Ta9i+7l5jUeahvDczMLM0XbU4q35QtNKl5sQMGIbSy7lwutQ+zSvVSJaz
IXapR/yU+M3+gK73Cei6D5OAdi4lhs9YbrdFZDmw2Tq3b0J3eMaF4WygyiS+v5oj
UldujXxRzbqGD81UkNqJVmSADKCW51wp8piyziNgBrYp4VNXrVlbED20+bkNJY7t
Ln1aJfyzwf9TARkwIPeIvTUyrcQeQbIsRaEVi0hFfnmnCdNasEIsmoJVjyEchM+9
AIVxJxxJHewTtmtKvlnz/whXjV9n5aptGQXLfIKQXrAsekX+pLhbdj7nQtN/YhGe
`protect END_PROTECTED
