`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8OuJamQ76aMnjchReK3VSI2og2+Y0w0W2dl1oSsYbPnecr926NCtqcPeYr2RfcLy
a4WcYsS2xDDebjQCjWW7X/DEC3a2JcY9OXGfeuf15LrGv7oYSbcU7AM+wsuXH6Pb
orZ+arBqetWWCCEicHCKUTc3g6cdwfez6JxIeMEasc9/B82vzA0rueAYhgBfgZPZ
bn0S1XbvUZ/2KZrujVgYGNa8Bh6VOxa1x2pZtoABdTKx1eVsF4kTME1BRnMSpG7a
rZJWTa7FUWuFwAAB3IOhwoR+xK8q98IMPZVbHe9g1K7rh70UfoPqRQ8YivWuarGO
eWf1ghN9NIoXqeHgJEB8+GMQ77ZhOIIFZ0PMmrETqrqCGl1aKW0NDKc1VgjZFSU3
ZIEEdTlPsbaBd2YxTAC8yfoYQvta+mbmL/eSOkoOzCumE333rVOnc0sQv48EsNF+
4x+N4hdsBm0Ir9hAVJM9NXydV34UoCQysL4zk99leLD+1K/GUDSHMlzBXoaB9ypB
1jGl1JnxUuwFkRSjJ61TSADV7c2J7vCT8Yw4O6cTG3c=
`protect END_PROTECTED
