`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uca2Xb9XICxzJe5LXwao4XnOxIQeI6501hFx/0Z5dZEkWSqV4g/hrCxp2TtUfwx4
dRhgbjV6yQ9suCSwYwRZr4V48ZUq1RAOGJCsoRQg6nfOpWFb9mpRECnOWeUR/17Q
ezLQ5V1grtAU/RtWcsZl0tRXB5y35Tq5OyFcOjPmT8rgyUpDzcwui4jDyRRuMNoV
SUYR/t3HPIy2yVv9Ux6PTqrYQwnKO3hhRNN8hEf0M/Ij8cJx11vS6OOFgitNxoRQ
HVcfBhxA633BYTTrUF4lM1VnPqjRZS6ZF9Y/wwhkgXZKfJwEn+Zpq8HpFaicqyh4
L173AtHGVc4jsxZIqTpkiMU4rEpui4LTfR9jtI4aCABl7ruppk2YtdN/PKmCwtkj
2NRnZ1lcA/cRmelXuiWrEtYmw7OtYy3quyeJxveYQQa6cO6goSpD06sGhavDROua
sa+K0efPt6WoLtNwO+1TLGJ5t/xPg5qOflKHvGUSXb6jVoeQidJ/nNEFo35MapNN
tJ5gw2PdsoFwHRUx/6x9fLHL1aNZ6sLc/yAh0NHTYgki51fLmkM4GnGDp9C6qzdd
iPs8fRz1b+yIIxVMn+qpy4ZdVY+fo04M6mjoVPR6sibvZxlsF2OprHyFCv0yBwNs
OcnJVNgEwQR6VzLIaKd51oMKrULLnvYbZeQMcEGnvob/KmFnkvMd0W19z5ZmeTP6
WI0yFW+2ME2eOxk5T6fe8w==
`protect END_PROTECTED
