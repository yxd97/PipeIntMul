`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dhkJLObqmDwHPQjBnalkVIPr4Hn4GojGxsxTFhIkaQEzfgoA1MRiWARMfiwisC6N
p7iKl4HqlSTIlfOHW3EjX9EeRSeLaBx7LmVIWLXS0KFQyIBbEcYw9XgZhL9owbfH
VIUx94zlMp4bMEgRCuDwD+aUgMEqxREwQzLOXnB/7W6m3guyYXumrYtQN0LCy1IJ
34uy6fJjxSZ5v/Nr8qyrL0fc78ed4zBcJz04yhnQygrpy3FB14KWqD9ufM7ogNaX
tHBDyG4mDk+yUWLu33DIhd3esbRbhI1kHcl62EjAzVEXo6X+uo+xRRxhQChxqe4m
lq18iQcz8tJDBwtmtjckCocgWP6uXnE9aVkXnyDVhf81De0H03JrgP5erq7mohLL
8Ox/pOzm9FyMrPIHjgh70a4pGUbQPzBPT7htUrEBEFZcQ8SxqYKDMaOnR8Gafkmd
seiSkn0cSkHp6ErQNyDJRR3pmys8nwPJpaJD9mT3JpFcgB9XV4cC23GDtECNWyEN
WhO3cgu0XiRwRPhBkTTkXfhNUSXwuQzHRN4F1SiUTeYE4doo/O3coTcU7BZsIgzn
bC5AQ4PM6JeomIbEga+4xRzEU5PsZNg2ytWs5J5dJDjgv92XrY0tS9q2PGN+ZB1/
YZA2nBNxaz2Mprgzm8QmeZ1gs8KmSdIDTRR51gEVIgzKnOPYb5GZQpkoxZ25Y5ZM
tx6C1uMPO0YtsKWlVjlVKo8zgPNb+89G/BccSFksI0EWiI0qJ4VDOyMvJBeFLVHo
+X/IqxAH9LoHo2GPUoIBpoF7WrpoCh9qmWQNmcwGwxkuH+E0EfGQziW5ia14vYgG
g0UejQrOfHIX6T8WD3Qp9DI0W15UN8BqlHnmIdHatHM=
`protect END_PROTECTED
