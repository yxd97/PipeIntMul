`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JC9nm4VmGdCXRf7cy82c2rzw6AZErvqXEsWPguIN7mJOoAYD4W3tqxgAx1T1ab3d
2X85yU3uTXbisv3BjlWm9snNaoTHZlen6DTblnznUeWVvVUe0ua+/pXyCOViNxbk
gxowHoBsJhbVJnM9e3zmhfe0h0qJU0ZzS6VE34O5uNW4ShSs4N7/82Uv4tfAd3sC
RTzxkITHIPaxDkqFBdT84vvrs7yTCea4jkfaLt/HLDr9Z721ZVOkWnoq3jlAmdXp
gkV2AEAku0gBu4/qJG3L+pMTBb0Fg9hcGXbR8wEgH12wE6J/T0bBuJmAkBAPShgL
vpYE/r/kYLIi6DaOJLPe0iwq7UlR3EIu+o69ujLYWzUWM1UAW889EeSZFDUgYqWb
tx+aUQ2ArV1O7+mZviZN/IphQdUcO4r8fmkoPTNYqBTz2RnO6a5jUG9zOpRgOJ6q
3H8PUKVdPLSllbCKlRru0WLVZBuwlIWqFK/v/i7d1uw=
`protect END_PROTECTED
