`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oNXghrbyGh4bYEIPYB1aEnoeZkoXOzmQd9BDrX4B/aTwWl/GVdF3DkOHPyPvdcKu
MluB2+4lAEYLTGgkCtIxC+obvqSPfiy82JHHp0xTh8m2nimFdroW9ljQXv5JF+g3
LUFMMeHPEbK1NWVGi5GHyKVHcXk7grkG9rI662mcf6wQaz4LbKuxLZz9qn5UO/J7
xVW2n35rNNlbRMtFZJLvNe/yx8WAautKndJH30xRS4PG9rTOT8Tj84K+2aCr68Y8
Tvu8g3MHBV2OnN7hATldZg==
`protect END_PROTECTED
