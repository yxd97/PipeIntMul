`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTxGLKaY4vt6JUz/+8FXNjjesUpLDEGNh3sKRHDjlE98cD2t8D30JdW5HE5rQ9W7
b1UUZiCF63harnJn9TzA68wxUWShai2hEfnpOhGf0Dh19vJJjERsTYjh+dfVl0ry
N3fGiThdwIqyGD75wfk+HjPWES11Hs22diBykVDWs5+NkfOq4OPvYKV/u8nGChGm
xaKO8r3AEpJZ8j8A21NJUXt7qCOb8K2hI81IIjOCCCA4/nETHKyNAlGHgAVTZSL6
Z1z7RsxeyoXd6+SZGBu5Bpx5UKfv6cEOVMH3qlPck1PlYSeyVgg9Z/wCXjCjXdU4
jgidU0lb2I50CXEAMOPcWzKpC+rUfrzSAjKLOEODyXMUqckT1CcWXhAKpRvYEt/W
S8ao7B4fbUAK8oLrnCaiTuGE7DT3sLdBzTgIZKzgqUZhsYSnpNaLEg51Za5cRvTt
M0dhGriTPnbgkd7ztTD55DZ7yBUS4/OW4eo0/v902Z/CNIs7LwkjBkPRZKZh0AZB
IXzUcKYF6Xff58NTRABWQ0tycEPauUOFYkCIWos/6qXxU420X18G/LMC+y5ixfFy
y873ODQdiKSm6bqbpBIM0qTFvo+vmscWfbTvRQn2MWwj/i2MmFEKEilNrbKVH8Ni
s2I5qnyI14bK7ncU3aCuXyI/6K3ny1VKwF+Zcv3oI8D9pOEWDSo7IswRin+Kk1zo
Of8L9jW767Y+OfilR1ux2XzhcZR2bfP2p4FpC2HHUhs=
`protect END_PROTECTED
