`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3JvK4x1wql2JKTcZpqol+2n94LLACpcCxzH/7pl7uShHWo99OH3jXfix4DHjpnI
NI72Bat6o3sGXooX0gvGmg3yFojmLkeeLInHvlh0Ac4NZdydTFvTVTyY63EFKR98
zdk0Vx44Set/m85A1O4eLWl6R4loWYQHlwNYhBQq4dbglvncnXu5YOEHWQ5ltTUl
fVAJIZUPpomTGWR+tI+rd6FI364oOLo9ef+0bMwLLCoiTccIPBIixs1xPRe0txXs
DMivhEM+d/OzBlFsJ0gJR173NFe4t6CGzl6j90Tu3b3R5v8vEpCN5cFm/oxbXnaE
dHr/vGZjPKMQjQXHVsV//g==
`protect END_PROTECTED
