`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZsQn6pZM5eCfyFqxNuIqBpJMqYocazo3InjTkMnX1sIJRsygXxDTif7Jos42rCGz
jE18wmP8bjHAuBd0Oe1sqzXV3cn8Pq9sG4t4sDacm7R3trKzFJ1OQI9aIMbj9MVx
MgodnjkPI+xeE1kP5oLsYuKIv52KmEJ6+Xw3MZyNWSolhM9+V/KuIR8y7wq167er
woajxgTeACUn2FzD+9Cwy7gLjJmSv5VjIyGNjtm33hBK+kWXCrRpp+5rD0sfUUCU
E+yitULsNvKQwG4+Rt1dRbCUuRvG0fZV5amqh4Z2/wNScFk7Nz1RKbbkgKiEoJBp
VfX1h6MTV9HK7xp3nSAloZJ5e8F9/QzGELDwA2Ofc/65Mgtc1bL/Jb/yj74RY4dA
QtpgDhPowMhQMBfxZowovovyCTU7wtgdGJZaR43wNT0yRbyQWiZf8fRRee/1TJ9j
09l5rNDFZB5M/jbEAUwnkwvcw6qoMsqoKia7FqvvLtw=
`protect END_PROTECTED
