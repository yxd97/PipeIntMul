`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6t7jY4iEjJk2NtUx4Pjox2TbNzDG4xofzwM2lWRRm9oCsvoA1HEoooqV1krW3uF2
oYfQjWfmWOwYmP2FRkgmUzzTNB71fe+i2VrlYBXR8z+qqoeAc97iMJEKDQirsJ9s
30ZTjjk3JxGi2KvHObEnxWO5chA12FPpuvcPQq+uFUb6DiQw6IKZG7lVX+Xuih7Y
m9WQUfI0+NwcdGFuey8Jlr2vEF3qz9fpTcSEFHHtxBb0fSVD2q07MuRWHJb/aWzv
V86nu6AwprvSsUz7QsEKff5yq0oFhgXLZjiWjQV+kxBSooQ8u9jzGP0Qx1ThflZH
ZMqTxZCRRGj2d+3BnmOZPA==
`protect END_PROTECTED
