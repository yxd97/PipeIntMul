`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ia2TbE2mDW8d8JNpjKGvdV60j/f14cuNDClGP5N6lNzVU5IbrSQf2SkwkPwdyi8n
6GDvdvj3N2hGAoy4jMUZtfEi+1exU6uXufQZgK4UwLFSoj3xMfNLJ5nZ4LX4/Dbw
zF/5AEiJb4PfkY3fDRrn5IYhiyJ9SvvIlj8C43rDBt9xQIc5N45RssDU3JzhMrgb
9j51KMSsPvv3ozwu2udlIsWfG4hkLoboU5TlVMQKlzrFHPkTHXtF9RKvIF4ItQ+4
dArzSEHtml5S9BBOd4zIlYwSrpkhyR5ei1BJZIg+agxcCjfyJWgz6zWz0vakXR0f
TE12bIQJo4PJ9LKianZaDUlV7qinHOxxQffdZXh9nTGnq0976bMnvBNeZWI2fx/Y
PDRMmYFpQv2iljFGbRSjjx9ePfnDHqhjNABQGD/MpEuwilT5VLCLabhO0pPWrGYu
RBTVmB1/IMQ9woCFYT92q94CcFkTosTrSd+VG08N93Yzs15IJE13MxkIUk1QKma1
6JoQvTpzAgoaKaGwjmWRb0FvLOhtB7IX0ccsSYL2UTEsH1c8PckaGZ+q0G0XgdeX
1G/1NrBtIk2J5gIWAa6FL+Y5SpZwS5O3VyOZfLwzaILneQN3YEckMudlIOKgFSYz
T3xAPmxniJ42YjFIR9jnEvV0NYgzlLs3AnwhPSl3ZOjzfpYPHPMFJFSAw3FNSx6+
z1BRDV7ANBDlR8Sw5WkRv02Qmopd6tS+QwRQxidAmeK/se4nfnApb9lglNEAp7J0
UcORu4MbSHItwsuxMVD+ls36TuRPyNpz0aq01it91TZysVGJcQ/39JtQ+t9YIK0H
fIPXo/MNSGgqL0M0mLRSiFAshbfVoYFzLB6mCY09KW5ful8k3GPBbdMW0FADEWdC
PR5+T26IiYx0jwIhUl723nhNFWn3Bq+z5CZNjXy16334FmRGY4URLlKargP4r9ov
ZhLuGdZNvj3CBNajloqBJoG9Q5rudFsIEgzDpg7EBZwXrpMVXAGJ7aatVvJmgurQ
3eGafj6dfhBeqn8lnbE7p3EnBeHV6PUbUjmQB1K4xnN2PEF8YYZpwewlq1rJLGBY
2ik99Emi98duSuFEuEkCcZMnyzcTdXI2d/ORfbMXQq3eoNWisskU3YDtSewlG7r/
U2VrJNfh5FWjPSZyCgahBsCh91E3scx3wPto+dy0OL574j+koo0skC2fKoIpAss/
sBfUiN8o63LFhkcGb6uVt5Kucml632fGfPtTOoJRaYJyJQdlx/Y1QZ9JY6VjxUwK
nxHHT3IZvX6CRoukgVi0tAl+IIQg3J3zzy4n0oyGy7IRG3KJrZk7Bf/c4UEYpQup
KudDVcfwJarHZsi2NpeZYxjlRy4MU9h/dsSOSGOa0uBe6CIIxye0DGi5PK51X+Fn
txpINhojiBsCPFerWbHijzHtW22ywgWlgw33hh7I4pLOYMpHs5B+8LqbIranlzzx
LZG5nEDN3YwQ/SGg29cIqztqt354Ept5/Q+oI9FqZv7hEkuIpigeGdpeUQhL/1IK
kNZv2aC8wDcOGVdCuXsIc4TlsjZvLLNeIQ1/dp5R5xHpXegk25Ee+2GrzAylZF4Z
uqI1+rD96BlZ8+atXmvMONPOs8xepWppWJTx1YiUGcZhCMbXfbHIwxeHpQxD27ZK
kwlckiMvnrIoBlAhvI68JAr0EvunlYNAgtXVigmRZGqH3o4ygQrWnqfYywZz1Jcl
yr8NyKaojAFfatGKxoDxcw==
`protect END_PROTECTED
