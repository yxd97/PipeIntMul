`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJGiuA9kcB0St1oXsYFMyntGrzBPQUEwjDujkQVzoK7qTtmQHg3fTqoU+D+RK/BX
RXiRfDsNEvn6K189huXCyaz/CYMFKVy6GJpzQfhbEMIYbNVLVGQw4MRoFVQi9gtW
Lu2W8DN0yDG+zd5aKiJLsxyqcyOQXMudOACuszhy4vqg2ooPLJOa7pMMtQEgitVZ
+5oXGsV0ygySJxrWUhKhrMoao0Wxm2Us4dTTEcBtJYzR5Jq74YSngD04rL06jXpQ
PZ5U/edI+nAcM/3csV7ufhNDz/NSGf1xfpOeRJEp7odHPs1IDxNQq/v1I3dishLf
uDuIuGY3nxKogQNF+PbZbFaEwPOatfb8UcjlnLmterE=
`protect END_PROTECTED
