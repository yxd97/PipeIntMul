`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yXxNwbun6zIAt0NT9eeozN2Y7Max8qoBzeaL4vk6yWDN5biwl5SK1AGahOmNrjzj
AmLunsXkUJReQkyQhfZZ6KmpwAgxRwccM+nc/FC196uodCf6PlYBJ+Dd/cDxUCa+
ixhiRE977kbBJnoaQwqmfON50cJL7eAcVg0/IWVkIq3Pt53y4iYZRGPUL4RKbDTM
r1AL6nrd9cJH0qw6W+4mTmcbrIhKbJlbokb1VVSne/p04TuIDaCmRifOL5tyn4Y2
oiaJ/7pExZWjG4QN4roYwj3fVtdkQwwTNhPee2XrFw9fUz/gpU5V9+OqaVHOTYbv
glNW5nNbMgFa7aNrN+M4Ue3MXjaK3V6/CVrEgog0mO9iPkENKo4P9z33HLvMWTeo
0t1MwKBn0Xjw9oXmJwpBj+RbkZaF3Bb7Ze+2ekedKGK65tyw4g1pGQ6Y7AAqG47E
qbXd7pmxWAEVquF4KBWwYckphWGVkQirG8WyxauxxLYWwBEMx0la6GjEAfUrt7QB
Fv200dDH8+LyrBHJox1JfnY5hjFdjAFjNcKgaehMlY+7nxDw4X+27+HfBBkBX6Rj
dIrjQDs+iZQ0PhnHJKpKgLXRd4675YuHZW4jBo8/praBVIvTTySgKqtqmS2Qne//
GD5MJaPaHkpffa/Kg+Y8e0ShKvvAXQmFrhjwowAjcXU/YR2Q155ZM9Lwqh95SBJW
U22sVvgTS7zZIMb6vkcYul9nSWbN2eSbUnGdx6dxvrcxudhWvRpsfBB7nYo8r6xN
ORkal4CdJ/vsvOch0gdsMGkkTaN6Hjqc7LR6f7LRQNldL+eXGWZgqrJ3Sj92cr/q
4F/2pFPDRU972CnkBC2XgjOJ9ec/4daBsTzG0Y82/Beo5+Qc05u9o10tBNPS91Qd
TOZZFYwurNUncxOVrDDSUuocUOPrq8SFLXUzJS4zoHPw7opKY/zL0FNZyW9DdF6z
oz9vRDhyQcUCCHXGB7lyhwin6ID/P5Ox01wsIEI3msav5kDSAyqtIgzXKixvaczy
1+yE7/hxQ5q+9D4U5wQL0EANSKV860DsPy3t4N4U+yqJZ78t6I1IW6tdQguD2ad0
NGz0nT3IDDJVNackJAL8HZ9SJCVqy+pg2whTI0Q+WMlIn6MsKVSvYZ+ntUX+AkiQ
pTd2DNP1m/K4C0BfxSmlOmZdpj1okEM2JggcMjpVmKaWotfUgSBkpYJCwHRQrYwR
qELCxwrDeFxtMP2AoolRFyfuqPYLWpqJbWfnItVwo/EJznSts0a5GjJNyoXKMV90
LsK4WjyHIyyg0mYrD1t3+2XYnAAXVNPKdkS9AcwK1EKM53i99IhSeLv9+65oc8Jo
`protect END_PROTECTED
