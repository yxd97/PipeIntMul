`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lf+s8PnEze/Wsui5HJM4lQYKl07ACIHnMrXOAVOYTYG/0bHrnnxpsidjGMpoFWg8
/3wN/4HZNeA+AjIsM/KU4x6NKPQNZkk5Gfc1DnTbmYqf5PkjN2cJmerdkIDYo4Of
BsSnheHPokpknl2hagoC94bwGFhUWqRKsx3y5zCEYp+VSpQjknJvr+aEmHKUj6iK
7QswuLYGnWmUptwWG3t8VmINrF/1AnfWsoNMuNAi/v00XteK1ob1NPt9gH7Oxr35
VhSpUdP1KhaT57UaduNV6g==
`protect END_PROTECTED
