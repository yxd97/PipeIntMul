`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3W35Wg4QLhDFcuC8hjnV4AAN7x15IEju85lwy6t/5E8XYm7O8LHGnEzEzRsK7kky
44bJUMGtgJlG2GqunDcX069hVtNxD8A+cgFCHhzyr74wj+bc3d+jfPptvp66zb07
IQSlMB1zVrwUsp69+ByG/mf6rpYEIRtT6rPNXNVW6ydhRVw3nhbIzYnVxBGE5uMA
iYX6uiGSDh+AbEf2UKwYU8iNv2JxyPboL28h/8+BcSwoKpdklQW3g7tkpy9AyayV
Prc08+zgiRGc21ItYGkEUZOUlADZmZlO1Yszcgw/TNWNNklFE7pfbvc0h1F98woe
YUwH468AQWEwZOpYrmuDjiqiDqa73TE4gveDLOO9rTKqKl3T6UFqRCwsIDJ3xedt
3eCB9uL7fMwoUyj/iJK8e21fShU6zfEhxMDvVqLZfVbqfyzaCe6wF6is+unEJw/U
2v7WY/CnCV0UQCwaq9Ac1m0qrIBlpyPw7qyYHUlii2Z9QFcORdKclfyt3+qN4tva
n8RCbdm7H9Jki2aYpOSm82eDFDXnrVQMdRTK00jws0065bZNZY/7v/4eGwar8sQ3
o9jhof46cn7TZvRpVfRUSukZf6gfqtcyO9/RYlByrP98HBPlmZMwMzh9yv00EIA3
H/vRNZiEP918uhVuSgIhO6iniMuBWZgRBTgcf8/PglsFkflzz4GKE+QVVLFSCCBS
NDzz79Kb7jlFOaiZ0R4s+958w1EzQfcgKgGv6ujg4aqcvNOFtYhQebMngB1DoVz+
Od/hm+cBt2lpRNHSwbNaSPwidoC1vFvh7q4boKLHTehjByGVi/G8wuUag3aLCkUQ
KzRwMYYTYmgAohCmeL8FVB0MoU9oUB6Fzb78CeyAqhzbqcHaSS5dURJCvub0xvtk
aa10QMslxsrP4e7w8sacqr3XqxgLqJOqtKOp9aVUXdGk+lGQ7MTeT54sxWvr3vn0
1afCz/xnExEW43Cl1uhAGXiY8U9qgb6PKOfYMe9y75/J8ChO8svEoxfMEBbu6Sw0
Ehyyi3DFsAMGlHqhKdgsgDJS0beeFaaazNgLSKxm6UMyOXZTPFlC/DgxlfUQOZdf
e9oYAZ5E6hsgtJ+BJOEox7XceS1cfoYL7wc/suxV8p0Sv4XcDnkdvINAB7IPTFDE
H6xrFAe8S3SWPfpEs4sz4b0amKSYfFdFkMB8Yrea1lje0dfpM9WYyZ2IKB2CoFuS
aaOdcfhV3HlSqvbD5ySX33bf2y5CnYw5iouq/PCQs16aJys1V9Suiezaomkg/xDk
nSp3QO55/dc8l4chHcXKM18RFfSeMKUPLZo7k+2L1lTY/tffHO0bamU7QXnMoDOt
e82i4gIf8CA23AHY8X9URZ61i7jwcNeFKhT77si+HNcXZ48Kn1jc5oNZR16HW1Ol
iXRAuQsQoy6lBA8lwGYKGvIlW11tGbSotUlC+2hktqU5Wn4QQOWwrrDh31T3dgBq
OZapIwrgr2SsQjugEQ6A1VUbg5Lj1KSSG3icaDfIFvYh/8frsKNeyrOYWILhmnxY
2zgrci088bmBpMW4Zv07D+Qg7texkcjaGk3guxdkmGitKPGK8xSNWc1HEo36SxLB
MxnUAGOgXLz4CklpgyE8Bjrwl7iMhM3QXbp1PulZaYiP7aNpz30bwIDgDBIpCAhH
2+E6rYzPO6u1hszmc8CCN9FGyfz7TmUwKq4zukmJPla4mdNpF3aTFj7D11Z9iYO3
l52Rd+48H82/scI4FXdrtq1PTrv0ky9hfKNgdpDl1XtiDBuwT+YWlBEs+oOuQx/P
6OIuRo7pbEo0W2A1bIMGSxwp+4AajQ48WhWUlInAzOPV5CibO9tOWLlUY8c0tRMm
KLjde8n3XD/Pqnbb74pQyywPSCHr5mKZpL7IZcb+0kW4sEEAtjQ60ZbTB7wstCFt
bWStHLxrpjcw29ONVTOwdnTsvPUtCBzx8gJJQ/Kuu7fdaNhwTPhcUBzhwMqKgYTh
BWYOC7jIL/9l+6U2/yaOXiFS1upK3j6Rbx/nVowuDwaz/FaGC4YG428gm6YEvZnP
fnupWLzbRlTCerPLvWQwWITHPkA+YPhBSXL1t2mv9IkBhzYg94QygzxZxu6U0XAy
FamM8+kd4PnrjqC+vIT8l27GJ0y2bLCkb6TvAAP/9ze1DoFeOYRe/e7/VnsOFMHP
WvvVE+r6r9+j2pZXlEGFSA15fEQcIvEpFlp4TL4PgWVil+RFM5EO6r2Y09TiFVPK
DYhXFZCvScEgkyQTEwFd+flQ6kxPYFqMejePIrC75V1HPEqJkjynXV82lcOh9Hkb
Juhf5KXprnRAXliJiTSx1StAltPCrdtoo4SiY7BHM0qYB2s1NlFl/U9iF/pb8Lut
vTMMWiL809Q/SviwSzhlZDr+lopkpAdTdXDm6pDSHPlEnSN/jEAyif16NOO4WoKC
ZmpEYddgS64F9JWAB452QNfOLFrdAvtqTblCxzAK163UzEjQdDXNBfRYS5UE3BSr
SNUqogTxtLXXzS7ronPjTlep1sCTmU0Me9Un5c2DRGJJ55nsUSul7SafrJshj76V
/yG6EnD0O/ou1F1qcuJh6/E8Aj2lGf72Xk5Gcvsk+1WGES+9HwIuQDZaCNbdYlPz
CC6/xhJNs415ZE4baN7xzbn/jnITo+tIgxFbEAk3Vnsl8PUHBtsCDOqe6Y5zyf9D
YQ27+tRLt0XvQ7HGRMb+D9BhYZ3ury1n6mVJSQX011z5ZHYTx9uXCkbPV2gEvkOV
rQtz3D/tHMo6tWh5FqTZqB0ejnvBPQbVZpPfgkd2BHziDQA+rY2tfeVTbDf/ImZ2
7Pg1bVpCzANCHdOceLtRREpO88RScaiMjK/DzYU1ZKqWZYMBE4nK8eV4MYUQ7wuf
RzJIDZXapKs2J+BiORpDBz1/oen5HLW0MYBt9l6eStUAZsn2D+wVEQ4sZzodEGW8
O+4OvEqBjAIiVaAKysty9FPnVI6+YhotxugpMpAKCBIg2BgBq6nCbOOOm1LYjMsj
VXTGmLM3O5buXkDlWTvhqKV6XK7y34IZqtuAd8R95/NJmOAwzCEB4+wr5BFDS7qe
EbarpOB+to+GZfxmkvHawJeYMgd4zz5/U0L90DXv7ElLk+WhurqFOm3BMSUk6l3L
oljpaSjzuqfGDYFQOIRZKPg016ATmgDVMRwAyJ8IyL35O4auYdYeXPzqmsITE4EH
DX35zXvO/i3cPGosJbyCwHjPL2vAk9XZQZHITPy9TMqfWLCuXtIlBCRTLd8CVmwo
H8/UwB6izofN7umO4ZbIJG9IGYhqyefRc12njeChZlotBtszDz6Cy0p8G+ItPrlN
socK78JCMOhLrdzkL92af1um+7MW0wpzitsN/fQgePYDvb4MZZl1pPKht0RhdBdE
Wz6oee7xicn5KG/JJY7XfcwL/RFMZ2lB22eoW2QgPtFMMPzTVnsHzIUpOm9Hr1CE
WA/m3UF5nP/ferKYYzA83ToasO0X2w6MW1koGfT0tvXHYfgX5pa+7skKPbiA8woj
vkEFkZAKhc27XffuRLCZBbTtO+kohCb+lXPqAjMr4qsG/xyupuqOB2RcSLxzZBEp
jgka18b23wFsrT/pMwscT2EEPwPFM2Rwv1UNvQdFYhytA3Ss4glIEDj5nLkJaMqi
y4Y7P1S/uUk+AV/JN2G1zOE4Oy58AdWlssp3pdsD//1ohs0lsU5MUGjPEsGulgzp
gAWlhEUbSN1NHk2XExdwO5nPuaI7CfxWQXmS/AZcMt2QecfI54Z+0RYlAeOUM1Xo
SZWaiiHLv/mCmDVfUZuWy3GXBNl11blChqSTHt8Vr3trZs2SncuZWKLq1iRyJz4q
4Ww1yJ9aK7BX6DmEgjbYBPGGLeCkzA9ApVmx88MEHMTZusnTfF2LdyeWseBRF/ub
n7ABZhk/Fg6IwOC9zFtQnI+3m6rNhJurF/MkomfuFIHZYlwrS+qaOyE1+4a0Rvvg
3tqPsdcUJQdBLa4Gjt2pY/zmYfIA3L1OyUulSQsf1goC0yCPej7ReTipDWW28HXn
9j0o+MVCfsKZass/0f45rxuVUU6YNj0flemopx0ZSD9HZ3QJp9jPe+K2JIGMVqxW
FHLfkGy2ZONZB05mXqNqqNnWBENKUfF+BxbTZMyYnm5ueX4wYnF+f6fZWRgxQQts
mofn6KzX71B692e6botFH5fki5yKtirr6oLDM5gaWKeUEzIckb12gfLvtoEH+QR6
r9C7xLE9yf256cdZ0Cb+jG2r/1uXoXFVu08sSXnCKbS8HoGBnJ03Nsx2wki5ki2N
09XRHcuL597dn9a7b7ak87oFdWtLI5/onhgzopeNI11cRy1tgH+58jdEV2E3htgt
M65AFIfHYQwo3kcEglolC2s/VKkKI8xFOaqAvUKeAfiat0QJ+DlWTjka7QNaqHiK
E9L752QdH79XhFdBBGFX8bu83MgErAfcH/HjuitOjdpGIiTPgrVhQte/oKHoDAz4
2QLB97R3EVl8EBzk0Rv9sCPF1SHYPgXKdCT1QUVDKjcGjmNWi4C7wJ3p8wLHmznh
w9ERTr5WeQ1WZ5AszO02z2ph13stCoDqTF09MK+QCFyVqTRw6HmzNCxJg5U1AHkV
pTeHYZ9udxI5SQbEyhlu/vUPKWXM6PpZpk5JQ98W2NVPzzdJ0DH3tKjNPsHc3Y4m
FHBWACNpyWYRggyZwRg4Wqwh36+sNwFMOdCM+/Jk82dOJLrPH/cXaeko3llkcDiA
k8zB3+0KmTV6riF7A/kdXF+Na3/ziwISwGUzALCr1LidOZ5blJL+g0SJFGbCkG6I
842EAPK6IOHiKfXjkywwgcoJ7JSHm1dEOvLj49VW/kl8IEw+oj3KUbHgX9zSeFrX
WFVFff/P4+FVa4VmjoBW+JNcO8NqHJmLW56cQv6OvDFGuaIRAcgTMb+zzETA+4Xk
uYjh/wEhXlL8dOM214NAsrXo+/NLZ2BHPHOa6Cu1ItSuNIZK3K1/W4t6ZmSpf+s0
3hThoYyyikvC2BUXfPl1LD4NVTN9sDI/VMZKpa6fcfBAZETHTz+mEUsrqB2YOaU3
FV4KAnGvl/CXAeArsvvLi4xNqzanlxtVTEJRcGRcS1tSubkO3i77w5f+PilMV/Ne
QJwAW1Ow5eviBqljfXtYmJXB41LpZ+DOAJuu/ZuXT54lYnWvQKw3pukh9fOhenxI
Urz6HLREj70ryZLlzLc4mK1gtFe5fnj6smihXXbMiM2Jd25HZa5lfb0VapTX4fxq
njeg7dpvANjppvWS9Yn98xPMorr4yHzO4pM3RBnaZlwKE+S0aezT4UIvcrjTuDAX
`protect END_PROTECTED
