`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GHDZBTTH+Q5fDdN+siftwA/K5aalXwMmhwRRuhSrv7tA9uEp9PcTDHs1qS1LaQC
NwcNXKrKw7hpHCn9hF7/2OnRroJUnU9GtFIGdRFohwTmjQam3rRksby6BBrHylfa
ZgVrojYAWK/Q+gJ0ykUJfNIvwBSuCCAVQakn8+qdu8bfq8N0qL4dzn5ePMCMD75L
SFN1tQblvS89goCVWiGZv9R86kvdpf5aJmkp/DgUn5du3gdyShHakSVSTJU+CuKS
YYVx7QlrQHCns1ne2aVvveDh2zJGF1Qca6y5SIkG2Pdi+USegByR35V66FATIUnO
HcGEiprDQeUxuW6pi9cAoyNW9/UAVgApwFaNFSJGmPV1mkcpUMFsWzsPeTWsFyN5
wU0vqQy4YeFGEuj10SkEZzmvLZvg5g24rdKVuy/UOjuSsn9hza777PN3w7//C+4G
1E3OlHL0lPLwJBx4+W6Mnf8pTsTkzW8QZwtaXtknR3nRqdNZ3d72gVlUwe22HoKe
QH9CZAxNE3gYd5qPBLrW8rVCKWWkrtat1sD/JlTlgquMvMQVMF7GiEKdG6eSlWqV
sJBCY+lpAYWY5vLPPHWq69vsyOEXSvJlus3b+JkGdWE=
`protect END_PROTECTED
