`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oC9twXU1ctkiuCqVWvJZOYOBBLF4QGTtJKZO4Uvdk4elhK/vGzIwJYQ6rPKIMdLO
agn7r0FfVjNbquhj+yRp4I4ut+xAHfL1Gokf45Si97iYx7Vv3475a0pnFeZdr5zU
Z1FN52TqLGXY67hOYiI5nal/lbQJANDrtA40kL9AgaFYi1VEfvjbeO60+vbpOQdc
kjZme13pYv1zgs9aa+Rp5+sVNLG225vuhaeiwlqezz6nTNRkRQugNRxdVR6UgRQk
g2RT2p3OId15M/iz4fII26r49BRJcTjt2taOfkbe8iU0U50PmQobzYPtS8BOrXX+
7cYrwQR0jnWrrZphZAQqFTIn2nlWSM3Po5e7TEP0aqNY1ekKKZssUGXsP1/xRaP9
Ri4+XlL8ZB4ktrLj7tveegUw0cGDJguuQp2rDMnLUOcBeRxodPvk9zzMY0dRCd+N
mrsG0gkk9vOH2K4obS/SHjtoI+TBxu0NVCtTC/y9xhth1nKsIg87IYt0rAkao0xi
IMmIb8uCf9uxIu3z0GnEg1ceJboHOweDrKyArgTaZ2Js9cA1zBjEun2SRXGrjVS0
OsICBOUYSUqKCWA0SbvVwPrUSQvjT/h1QGB5KYcN0a8=
`protect END_PROTECTED
