`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OQPK8F0bn4NtJJn0AkOD3aeeFq/5/0pT+8CLmqJXCZXQYpNN9HHmWTFkZlRr8GBd
Fg4uKq3UCWMiI1ygHzT9mOe53SEXQqrVB3gB95pH9LWAx8REvaEnSpfphQTjmvnY
765PeffdVZn7X+SXAez+yGuj84uRaTQRe98SyET6byly0TidhJudWpCgwB4BMxl/
buaHmvkNkKiV8pFg2eEuvJBKxa6sohokOtfTnHzRZVMWqdujGhRuYoH2JVUCjPYi
7QVkbYH43XFwHG+SpGPdukGbg7Yal35HmyIwXFzdP/L7DyFt9/erYtPt8NRB1jOp
hcp4PO0maAPPmTyPdoO2PO3dmuHeTnicejQNSWlk0AKIjIwI1RL5rWzXkhIFykrS
MiVaDR+VapnEsb9AVZb7QE+NslQoMrOuI2gNVDH8diq+oWaAWOIahC/JU/OUzhUK
ErS6Vu4VADWWQaGUaZ7fEWG0sVwPmQy3+Ix04MCV3lpj0HgZFa+1G6GRuUMRot4G
Sl1b/n7sbaLfvcslOE0XICWVS2WlNoia1MgE1Ti39wVedlOCaIFJAjnbGNIGkK5I
TOPHBle0sctRfqqg0nsj2xdjynkeDP5WEWOdmmSyRi7iLwnH+VAk8fQAw8lFZT5d
WR7XtHMQY1kKe+3SyL5QB/GMj/fr81MpeBZOb7zAik74KH8GNMmcolezzFL8XiA/
`protect END_PROTECTED
