`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Apyk/TqzCPK9U/PZxuFlOX3EkmSu0uNUcxQ53uVdzCkUjhRe3hOH+J28SgFZTUdn
CNgX6nDgufJyPxCAoZWjt3DRGmNp13C8cugCylV5JBIN5A+F88BSMUHmgNCXGDow
NBUXnmigNg+3w/AiYNxebuwMTDZQCFeQ4ibQXZ3QJcSLUNxxX3CVNk/LwcV5tPw1
DYmBkDanvGUy0MgRrD6jKF0v9+vPi9+19vcQqygpKYcQRB525M0ES6klWF+J56w3
0giJmm/G9PD4BYxcRqG03BaC6fABuIIicwxiZ5VuIPeVrfeadU+6GsX2KrDssN0Z
7pMw4kmrB0VWNOLMegAO5w==
`protect END_PROTECTED
