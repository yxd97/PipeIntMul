`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OtWQp6f6iXz20W3IUPUR/0nwHuNdVosy9jlY5lg2yz4Bf0ytNytAEstdrlLOBHa1
VGjc8k1zSVfcHCRi+qC3GRQfimv65BffzkG/sjLVmb6TmnYh+a9KS9aMt5X2r8Uw
9SVPv9K6tLRTvlFJ2i7N4aWetmfbuUDHevVxJUPJwIsYYL+GSRKMtOSekXtkRyDt
5uXm1RstZnDOJ+36vghx85qKo4csn0UAf+U9RIdgIquoi89KZZMm6WJ8JrFCSpBr
wjskYdI+siHVen3QpHlIOPN0AKeskKVh18+LlvWZhiaaDCHD3YBGFmSZ4Vusr784
gHzNKOoA6zocl13YmkJN+1uq/KOVJu8gVvqQ5KsE9z2kKuX1kWN3CUlIRVL2zWfs
5HnD4b/2kL5tllHKriixpp3T722vc53GlSvnijV/veFJGEn3L2U2UFOx6LZ5ggyF
gvrpWRk5rr3n9zgvmQm9on5knr8KZxCA/pplvRbu/2I=
`protect END_PROTECTED
