`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
38CpNqHEKw/2tG9aOzEeaq5tqO8mSzapSbUhlInQ6eML8ydvp2Nzan6juyE3/Dtp
Cd0CYSJXUA/+FeAkT4bTAmRTWfTs9+UVPl2UXOwdH4DexWzpxqXe1ot4yDINdnkv
Z1H1BU9VifZ5HSb99whn7XrQNhN6OTI216xVN88U3Lqsaw/ny4jLjnlyxHqVdWQV
8ktZIImbsSYpHLSmLFTFlLKkTryj44/SmVqJz7MKp4TmqcQ2CKFUamyFXFKRrF1q
3JcUfoyq21mWaI5y2MYp2qd/15ZzwWG+eETmQAXCttP4ZIlYP5cuRKM5LnUo4Jg5
1m2C8hzIjFVy3QwfAoVWK5+84QThpEoksR1K+IABHLBS51oI9+omALz5c71vB+2Z
FOPl73CSShenzIj5TdYumpOWZT6VjA167DKeb70iaUnsk76jfMp5LxDB0EciTk7V
IjmgdyQjE+gwsIVqzvKGb0IsU0iXuwgSyxCiC2z6boAGxIbp8tXrhtKeBBrny2JA
dsoc2AfqKemxJLBxV/RyRA/wpSlhwRmQZUWtguek6oFp3NuBFDVKFdkL7uRXfcJB
2evubRgbO1sbHJEAIWQn/yzk7HmB71vwSfa73cK/gARcN+8ywQ60dy9bKbMfsf9x
SnP7Xb08aCDKRdM9+KddhZeWq25f6XwcF5QhQEEkEQHAAZr9GjVPdImuCgpFfgBU
YlFZDsinzTyjvXXPyttmBhPBP9ERazxhqPo0BEmByqkIvSyhlER6SrDI05s3iMwv
aH3tV0q6/BEfBNYX4+eajWMTZpMKydNN2DStMP5Tj+CoWHB1Zx+DzxeSKz+EB3pD
AYS76mDP4k62m2AkW2EdflH5THCPVIzNthXPFFacVnNt7zfncxb9CYs893Isrf1n
wIO7jHks3eqTatAIiAsPULvU74uDAoyMZI1MQqBIXeVC4CxOblC1TOuj2BCf8l8f
`protect END_PROTECTED
