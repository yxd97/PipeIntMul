`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxglMHcBZVfwFgSFGyfHu0CnC0ftvIq8mi+VUEjdIUXvECnzMOlUSvqh9z964e5m
+TzYJeacGZhYOkWqm8lM+Z+RpqFNAw9egcTDl+spIPzDiFSG3OSNi2MhbkIvz6Ki
w+wibWHx4txvsMAbKBfaXX1326vJaqp/Jro26e5sqygutce0QQI9tv5MLIE8jCdm
HTvviP9j2XRp9xIfu5WBZZfexqOLSLJpFjcXDAT+FEpg/L8m6b0fKleg3+qBfZyl
rM5+Zmnpn2kwQK3EOCimtpCy1Ymd3zawjm1qHzBX/6MzZFs4UZs6sXJ+UgLWh3vD
NCjqgEaJCmHLcJ6D4aSJ78hN/h0BexbWPBnMuVRagS/OZTNi6VxtVJF3gd27INSR
m+XiolBwc7N4LzF/QMgPcI92P1Mr2b3+HgUaARldwiHzU8S5AqsgEJt1gWBt/kLd
ozC+zUKgY9LN/eBFA0HuNw5fSXIGDTAiRefsXm86cGDAF8CD5bhHI4Bp8JH1oZd6
Qmp+AsmC2e+qYJ5v75Swc1/i/GhcDOg7xghL6q0c8YFPEu/1eDNClbjHnjsGKsd5
CIoZzsiR2TPtgh6UOzc1OzZxz9qE2txenr3FM3jiw3iYG2IKSSTmvOvJeFbOwmLl
Qoj2mTL+3/yUR+Z0j64tkR5OsXN7Wo5IKlMVm0U8RlM=
`protect END_PROTECTED
