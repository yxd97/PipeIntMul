`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JtdM6SfgouIMUUQ6naPxCwJq8zNdOiek/qVUnVuYf9zPuvv+ljn4HedTNEdS+kmK
Z6rNxXzIDTG2HwotdIb9PYRXCoE6KJhv1dxdVmhqD8obS10I5nyt+8zK+bl8ceb9
4tweemb0kY5kJblGOo7AHsnfahzgIk9OzkW9ZFxrj1p+786p+SjQsFWKe4AS/bbA
IIuNEXSRIh3H/o9vYV0hIpNK+LbadHJeMuwH5a3eX3jSiJVKLrEAWNm3gz92mUnI
WZy3HoZwpN1Gs2zmCvtQ946R0h+AiQZ2SCTxQhezpZSsH3l1ksXlPPHRcFbiunbZ
hFbrCx/aipFj3TUHl2GSpQL/OpzaU+viZkMO9FVAQGKjaihVbg7LP8ZuaTty8fCn
CEK7ZbP2re6jZwU7y25GRpQKl3BexgPUpjze+OqhQWsunZCfsA6ARh2uDJKAF75R
HHM+PjkgB9sqlpVyobEqvKKX7xE9o4Kc15bU0x+kUunJMGy5LSusSafoGUlrKWAt
MrdsW/ny/rwKIORnkUEYVnhV1yMy+9c8jtzEqu4remQK0zgjmpKlMRnPPK9X4jom
d/vgpLAXPCZ0Am8ITUYY5yWhTN3tqPpEGWJcamZYu1fg5Bl2Px0Yg4uBKL4nFhlI
Wp2W84YZldpM/qZ7sE5eUaXA9ZWovyeU4p7tBc+JvZNy+R28c7ffAnr27/0fWc4N
donI0wOBpTjJLeKba2lp1iPBJd4Y8UmcZemAH5aJJrDDP4xdlBFu7StM8ejxZgV0
yU/+zYmVK9mt01lqyOkTAt5JKINcv9zy+HY8XQF7lC1fGyBIaRDQLVbZIZUZ2dQW
3ucYBO21bzmXI2nMoUGZuIG3CwcHpKoHM3r7qrrfBLfmI98PAoZ5Qt96IX06/1CR
sEVTO4AgWaTsgE8gOCP0XAllk/EBkxmBFOzZgS7oNQyhF3IRnc9m6It3kuWEvQtE
njh02mmaxi/BoapLj00Qo5PuAB7jvPeGg/yI4O1mJW1of9lBaEqEEmqDAir10Pdj
1pVVMd7Vvcg/Fx6uqnsypDp38itao7FK2JsvtGQNfa5XEcfUaPXLxG0RzjI0rnOM
l4CRiq2Mho6JecnQBzwNFFmGKLlPYsdLz5crzgRGoG+F3QfZ797JX+nBY4Ef3EyX
9NU5GAXoNABr0Zn5+cyO9IBapkJi0I9DT/MYtSktPaGp6XKqdnPfFczQXpW3Su8j
iXDB8XmoFjZ1Y+u/CUKbgTuSE6/jJ+AUlty5V+GDDxH0GIrYAWY+ph01hCGeRmWv
2TU228nme2JKgYozo+inmUnNyUtL/R3xJG6AjjMiJSepzJruzorv7qC0upeHjy4g
gEvCLx/Kb+6uknrO6l7IBTwzkZK54vkt/EfNbTSsfljkmwpYODnHAe/M8jAGlFuu
7wLGbBW8C6TmMmhfg2Xu9SNUcB5APj2Z/sXd9os1jcfEKgwTXW7LRRiC68BfeG/H
5cHzHiYvgX3sq+8tCRnrPtynDERqS15FdAnt2sr74kRZIcg5ueJQzzwtzkzLdbe9
oPTHP0+y/DCD7xvXZh4k1QYqM2J6q/xuGDdAMiAZP2tW7t+l9+9O0dAzipU8cdb1
qwgbtkdhhiR11Wnz95ldjJCVrTMR8NiKTeOvwybEMClVfQf9DRuxK30KdBk9OVal
ovYtLnABkAJHmTvKXtlGy7EKe/LGeKY54hIvm1Xb9O+/YgJmNJ1ninmOw7dgk0Wg
YKl15JhitFKWUc28CjxX4JYzn/BEhc2jPd94WIKjGFnd7OE0oWB3v7o9liCaUrt7
TqoDNmbMdWLtDn0IQ2M4AHMJ17veFOlCgT/6bUwUetZQGvXrNMIADRKaYHmaxIbB
xxAV3FK/X+ubycCVAoEuTIImDjClX4IShm08YY4Mg0sj2URAtosqWXooWk1i9czO
Jiz9nkFcK2Qd5RujgGY8QUHe+b+ydxGZ/U7UKEaJLR+zTPjikPWakWFXz2OEW5qz
pUv0rFnzYkGjO1jUrXfr3i2/PibkoI16d6GVOXxsuDUCE5fnLu2k2YaWqZ7c+bp8
H7yEJ+ZXItJgH1Izuarguo7vyxOVk1hGN7WXHtDK2ut+/zv7COlHvy7iUE74JUL5
wAqGygBYQr6UrD0+om01fVbWIW13o0wztE6yhqD9S/Oi64m/Ln+lj5oLoj0dxlZE
LyRy3T6BUTb5f8UtbC49Y5e3m3UE9zRZuNTCOLtR59rFzKmAawfMsg4YGn/7O34S
FDpYFtZFxPA692yDJawlcCSZbcl4US2paUBJCHBCmoCenf/DQefE8Wai/oGbJST/
67y1er1XuHSsyEXzDuwvkgVbJKEGmQpPIkjakemqyJSST11oNShaWU25SsdoD+6l
JowDySTLsoNSFQilcpN/W1uB3RtkthXPS26MdNF3epHaL6gcFwEJZtiFEYKjt1or
z1i4cb+LANnAu9J2725Mifyh6Ty5N8xrRQDyuDcznfhQ0+DYo3hkNyWYD2tRGdSa
ibTFAMrsaTRW9n1aJpWcvv8tnucJXEqHC/6t4mIXqFyD2RRxic+/mJDjPOt+mSG6
18+wggVrKTehtvd254lx7LN6HsqcoiU7HT/+fH/BZvOnyXk9moBHM6L/9bf2XrMd
p9kEJStOlrgDrkcBAByXbrcgojKFja6Lz4pnCaAuBP+d71PR1KiBburdWjnbIjUj
bolEx3BpHoEGotBxRRGjJOWDfamBH/T2193uNyrN/TlENsrt8LX8G8pEudN3CAzb
ZCOHygqvd/u+i6/0id6JoKGQfyJ7y0QQE17ADoPki3Uf4g1n5neH9aR34Qu0Oz0k
1tpUSvaNMcFFUG5C5Hoac8IaWA0iLyIe4n2ftCzUxkWHd7HHTPk03ZH4VITStLTN
Bs7mdmkgoTa0x9fkzZaPtYc7XAEiusJmrKDfQf6nHek1cHGdlupNrKzPrB/28pC9
7tnyIkfg8xV1IUPleLxBehYGpZqy/qgl5FmrJVYrCumf6GwSw187C0HTTTyW/F7T
sChZD8PJgONq+WzSGnwyca81c75mImfOMF09fTAdGs+hvYtMF0Nth3rHQp9kDJuz
W5x2DoooEnPxbqQq76fGyg7SmKj12hZZiL9ypfwqIUKCDQyAMiGP1BQWdzM+EcBt
PYoortDC2msCEWdErPO374d+O4zb8ZzBcSE+n9Rxcf0HFW7fw9yXkYV+CQwIQDW8
pKCA9+uFvD7KyTWxNBTN4kXnR9f/TaSoCh02bf1phkK3Fu1W9+3lEpmXQg0EwVo5
QgVmUr0fXY8inNaYJy7LaxjPHPZX7neEGZcWmD9d8aw=
`protect END_PROTECTED
