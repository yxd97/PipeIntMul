`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2KaMBFovWRRdPJ1TOiOy0JZZcEdNJwwh0PVB9Gtl7yGHl+crKeLp+pQpvXO7rLfm
s42EZ7D9pRTfpu6AQYxmdt03a6ybcCKN4Z53XSt9dYlAu4F27cOSyS51HVDKQKf4
oUHx/E02TDbQVNG8PI8MGjdVnmp1OaxAnFMi+HwwultdJxUFhmyKydIIw8pcfIl7
SHO4mYtFSNhI2D7G2qIIcDwJgew4Sl7GIf/KwKOoPLifuL6GciHiYcw0w70lCwVK
uR76jQBBF4SMyH6UEPmyOLhsJbNKK51uU9slxaoM3pMJtIUkqDrSaKh17agzM9MA
VPRfzBaIUldibDwzUvOuzwBGJ5wz+KYopdovYNnyHVO3Ai3kSmkBn1F+fCgiKRxB
kwgg1uur0mfFC/Pny9bjqULQEG1RUVFXRnL1AKOnsFkxc7gN7mAd8tnGcjELfsgq
vAD4+jcBS3bhHqyiHyHeqln4EdzvjfILSNTvTjCb7L9R5+buI4qkU8pDwoM7a/wC
AWVvujqV7MZmT2NGypfvQ7T33lUGfJLXFpM41qG0mCUgMj79zjIxPGLHeKzDA8Da
eWyEgwpmzPwbsD5nbBaaAd6TJCgvbRR7sxQoPquc8m8=
`protect END_PROTECTED
