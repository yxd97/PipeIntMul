`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IcA0x6/Z+WgALZQ2jyGzEeQZpREuhSx4A5S97ayoAxB8RyXqPKrf0YgIAu126x6f
JC9CdU6ochnEBpTJD+tcr9zWW97Ok2ZnqTb6jswkha+1qM+NL47d1e587Ok3qLKh
Y1ai8/0/fQhJ/FfozQ3rb5WSYuJmpJes1SUoCnOp/I/wdmV0V+j8lT14g2vhy4BL
qw6FQmGSjvkMSQcIgR0khI4FjWUo/EeYUBhlt0alNF0qcaOxh1NL2k43hHh1iH5K
kQyeFc9PmYdg1zRW2VTVHg==
`protect END_PROTECTED
