`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B1yDVMa7iEAhBfZWv5/Ku6UlBv+DTOboRLDoXZwFav/A6FQRG/dC1pBg0bMVilnB
++uC10PheQjc6KrfZ9DQV1mw1g9ctZZcf/vdHWrJGJ9K1gp9AbcTzhLqhfvW3pSW
EFXLHmnBIyafwU289oUIRqXN1Fe4CJ6L1EOdiaO2S9gHFcM3t7zPObYcOmUNgzSM
nljaZ7XoZ0Rcu8v3Us2AUQKzXjg4rdjy2DRtwdRoMs52hkM+QWgdpR/BXgY6IOix
L8UPmidxKo7bUG+oFF/BObZKcfqbN9NJpuQwOwWDkWqvGtW2LiCheZLKcYWWGEHM
FtK65P7yp3gbozxw4kiZb0hExP2THOFKKuOyBxy9zL5bePafouRlAnVR46NSwcCF
Ov0svnz7KETCCIjsUsbAgH9jQ81tTtvqsadI85dWE7tjzv1PyYAvSObKBv3cMTN4
dPiv1+KF5/WnqlnG6ajB533WrhEj+IQA2tA7CwN1XRqvKol+x8o8a+9EzVhlaeCh
wbiEku0zAIKpb4ed9EwgdZBbQ1clYvJ4Uq7554p+tWOMRifyHSCYwSnEj7+s2qnw
`protect END_PROTECTED
