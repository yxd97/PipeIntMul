`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQpD8oiZVZfKFtG/hJ9bTcOojkEjUs5/5OrdZaBHy0K4mOUviYXm4PH5K6Wh1/x8
ZuMXuwhSh4PJudZR3D6SFX0kThTK7XuYbIN+Grv657DPpHddVzJB9TLlf5FbKJpn
D9OIMycAEY1Ap2Ivmki/fOpjjhNzCEj7wpRNupVC2zUMcPNRzVp2HL2v+O3i1W9h
VHJwNe5+LTtLfpCBrXM6xESX/2Khs5W0FQAOOMPR8k7PF3ZgTZNO50BHU43QtAWN
JJdN/gclBfTqVyFp3SKtN3QLe+lWnfRFAh3UwXJcddUFEC6ws1H/W1KycTIlCGHI
lmkRZFeNUnivhtB3Wv9HoO10rv/myDwsAk26zqSoM2RsW1Uis7dJ2XgqF+tZj7VN
HRDtoAGI/MnmUg3hxVX2yfI65cqYrRS4j2Hf45tuDBHUEWP4AsJ5KHmoMPQbevD+
ApWSk1++5kMCGkHqW14375FVQTiKI07c2bJIAPD80QASBKVqU95ItvGh1PbqMdaL
/RmzySIzTDtE1jeYm6iKVo2PJSlLOrb1NuVyb8NYsAM=
`protect END_PROTECTED
