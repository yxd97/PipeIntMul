`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ttgt8KFDs+C7pMq1Gs6YQRQ8O6YuH7d8EXNRkTU/WeVzh5/9JZD0x2n0Q4Hvho4L
x+b1osu1/0iGVn/BH3sBNsOaSpw6cq5qIijN5LmUdvnFv/6rUxtx1I6uuQwT/r24
8NfJQR+ees6nB+yTvd003SUXgp8JS3qBY7/qDj23Yi0kjyWLtrgvCdipHc5thdXH
YVWPJsC9IY1Zf7NbO+9ZZRwxXvOItO9ER1CvG3Q4524joGSAWmSVHJJNTUdSL2Xh
uNyAyWI/k7fVlKr63CsBtQ==
`protect END_PROTECTED
