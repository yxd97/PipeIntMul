`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFGhC/5BYsbyVP6+pniy4tGVCjgJwLXNG3FHykZ9JALa9MwDGHIFyNhcGS/8xHxG
7l3STYSsPU6bfCpaHFJ9YLG7FvvoKgQu7bBc+sv90v3eEU79AjYCcX8fTS2b/RX0
SFOWjfDV15rpTwdHAiRF15KmqFoFfGmLaKOg4C5Baq46lRsTWmSxXxbsKvz5iumq
62mAmYP8cLzBOx7xVagX8ZJhCNM9BeuILx2RjgpeeUTGOoV4PWS8PRws3hEyml74
3byusFWdNZ3pjdIg4B+0IXrWGb5JsFRR2B09X4Td89zUj8fAruI9qz3cUlDEjgo2
iSyjjCd2c8LHW1JYR37sK6QzH7KaqtOuwLyZ+n3/WhAw0rw9AhXlAc4ihgr9nXGa
De1sIIH/w+tLT3WCAnkOOwNu96EbzMvIgbzKA8NxbnBAsb7jTt/z8vtUL83m3wkZ
cAdYg0DcfC40VFhH+qXlN9p2Dl3fc8UohxZluE2hU0B+0cIErXwLB7zOleOojDrM
+nQEgaJnfHlFdbCL8ik3Ds2DMHgl0ObWg0qiJFZNgf5/ZoLTGukhbO9txQjkAIPo
hO8k9ojppJYzeDGvlQzd08ObXwc07lk6y3AqcJHiM/tARyx9yb7P5SEtKlo7VJtx
8OJRccURpsuG4MBBtLzV4gvHs++T109J8F4xSpTBiOLi6MswzTf8q8xv1XOCf7OU
anJPUfqKId4FYOESbrjBmLUNvnNum/rJzuV7OBO57xVkanYuuvNps3V5tASbLAMx
boJVeoltiEGVDmFJyUp6n4EAw7gdepdfP91WgMbvxIbBPzvfQdHRkw1D/w1tOkyB
7wqdmjPHvWjDUiVuX9DvO0l1ldXxfhAEEc9W/0T64JGMZty7IFph6wPLJspq+aW2
hsg89pgQEeGgWeSOcG8HxwBXfP/pDiqzLB0+yZ7jPuwSKM9dA7mPk11wSxGyOLoi
90ybmwluqMF+LI5VMXpCb9bt1jGX+Bf6cU3qpZTvRfNTQZnC7c8yP9oBWg4yHalT
zgQzFejnNB08CEk8vDGaKUc4lKFT6lkPvCplUE4WNYKfCrm/YX46417xh5nB0NnL
LvnW2j7beCmnstyVxa/0/5ds+8XKKMgp77pW5tWtPvjqJUL01/xK0Ep322PfhHLq
m4egWf7a7VrMCauSCEvzig==
`protect END_PROTECTED
