`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ObjbPNhRF7DugsZ3l36Q9058yZeNgYD278811hpTp44wq7uvT8mpX5GpnnbJt8l
5VTSkJaIbRS+8SaVmYyKYuG0YbfG4Q4SrutN9P23fdAeNjoYhGup/Duj34bDWCE9
h5KvleqeLXo93hK3KN9m0gmilHu/4zv6Yfuh4nPWwJPQfMTF5GDRwE0uwYIRq4Rw
uVpepWxfJ0wZ4z0GImmFASe9TLGavRl+G4GvkGgFafP5xIS08qdVBowhhGWHYgG/
UOF5BIW7RW5e3GbtGcKHydp4c0IJGHAAJ7Lg+i2NgfsTGC+1jTGk8IZEaV2EWGNC
LnHw0qugxjXgDKQbPMJVBSoK/4yOPK/eki3a8z7imyNvzzkfdoKl/+QIoMn8tbI6
PGAiiMpWYK1D9E92Ns13fBN06Bcj98CSSFc0bnjz0xouRVNh3r4K69ZtwzE1TSIu
koaXl6qvpZCTOTbUQd28jHo9LFBKzmjhbXJL6mL1q+wZGMIEpYlC7s3t2Euiw1c1
iG2rpWTu8nqh7K+9yS6x2duV6ZDA22PVKQn+pukmhUCyxQhE8cX9eaa64qMcdv/Y
q4qqVvjDUFX6gJivA/cgj7ANXNpF70mQMs5Cu2M7cJa1hP6zOU6U1nXkwmE0CUrM
MddF5qmFVvoZZ5Zefchz2gGwpP+tm5wPOCJVNgxKEat+10WR2LbgnWUwrJFxrfKx
b+xiNF3QShoVKrf+btXKMw==
`protect END_PROTECTED
