`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEUPyYZvFxGsBZHbeO/Enc7CGDfIdXLc3lCsPlfbnpERMWZdy5YucRkbwjGaLyG8
jwuhWzU22q+JnDrGnT86x/kKDToaznB5gFQtalNOQ6bbeH1s2AbCUMFsYpVOK5cW
3Z/14I9sxCfPpRuKKwahfBCwMbOc4L3/fHbdwrJk4a3auimLC8nEwgdqUb5dIApv
hyd6ZN2AHeqsMnwyZywwI6etXNIT/S/ivVoEQVo2+xpqR3gS+y6qdkWkYGyzEECu
KqZu/mp7AbnmB9Wf1y9Ujejoo2ei4Xmqs4Ql9keFjQG7IF7zX1bkq2L42dmCXN6B
WI+03Vzc7lCOVgP7adeEGQ4jUvMKSTMas1jpIcU69WoxHM5fBRDCrGoeQW4CHNjj
huJ+rScqhFe/6iTzfuuNF34Y0ajBargDaClk1xRPenCb89L7AZzwz8gMoU6PfetV
7S+GfGKQkk7NYQOgWoJGx3KtMvqETNj4moPo9eyfj8yHfjU4VPVovZrcBhC7YhWx
`protect END_PROTECTED
