`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7l62S1PfbmNGCzH/ijoVaEUzuV4AkKBeQIXD/l0lZU0AMihXdGKjIfQxhLVTFSK
3PNWt0H5pCsUA9lGjT3ujFzaih5CX3wOolHYAd7EZcYS08rs6az0o7eneTq5Ad+4
KrK7uctoNlNpjAp8MZ1Qen/qTMnI2DsPUyhVzbYwhSKXroPZXUM7AQv2ySimF+iA
mmWkS/KpGC1XOd1/5/FLBY0GAhrMKjCNg8otiyOVwJFJJN9RnHyOg2ccjqQUdpL0
8UdZEAxZWdHKxxXmOZ3O5Sk+C3ukq/j7Y4uOnB6RKSMsmwZ90hZ+tuv4ZX6daE4b
y0ILiHtihQAfxy3Ud2Cx8fBVfOkLB9ZQkjfkBWXtsKcmcbsDlBPnhCL3TeNKmFE6
B4Mw93pX1IVDlYp3aJnrUYQJ132+iUOtt1lU8kHb5bLbXBhxyuI8RozjBDg1Bpbr
u/a2r9gMfinXVbBfiUrqliMC3qKp3WT5wjc5OPgyYqS8UtJnO6KSuaoGBe/Snhiw
fwIWsF4wiNIWiD5G2Wjp5uVOluiO6AIcMxzXO10FICkKUF85TZFGtkzZ1QSyCQ1e
Oel4zfbcxwAkMvwl6PCbRDjG8S7AGWOfCgLROx5Yz/Du67IkvwImZIpMru100fsG
kJZtG6OAdsNxEUzxDzv8ZKk3rwr1AOtmYUY2d5crRpB/p69ViD74WToMjBty7rUi
s/o35zXXg64AIhMKIta/Ti3D1Ayx9SQxQ8kuNK4cXUhiqK1j7gRbtKXOIo9KGotk
dt0HQIr2VGZP+I/JlBmEqI+rl2hIkzbgT3syidNT4amFVfPk8MEMU2luncKYNnGN
hWoM9139+K6XB6XztNv90l/1ekV8R/GOXsiEaGfq9/d9ELRe5Q4HxoaNP516iubp
ob5LrKX+3dhbM+BEasrNkc/iJ5hCGUatX8LokaspGcJZuu3eqhyvXJ7Y60/F2wvG
4dPgFbTeLvCNekGT1nQ0LI34cgYmb64UkKWjgM43+MG1MwsumrvrkzNavyWSv8b9
C9qT2MDteRlQhb9DBUWvUNNOfHEGL9dDut5ZNJ2xgHuiPbPvg81Am35yRWRoDvtL
px12w5m7OUVkfZraZrLI0Pb1j+k/yc6wmgufzZY1ry1Ej0NSRu5n/qZQYQmki8MV
ErH1Vtfvd7sX/acx4y8d2s1ZR3mVdzirOt99GaNaxAhdEEwj/ntQcXbK+l3GMkMi
nr7eM16uRjyWeujg2EzWYM6IQZWmNFgPLLs61eKFx4tqadVlo92v7xqXURlDf0tS
DMZNGD2PlGK0thU6cr6z0mWlFshTjL0BLEr6TZJdCcALl6YN6ymte6b+Xc8qGRC4
vLJCHLKN7t3YOQQVbQ6qG1dsiuSb+o86cU4F/EHg4Xy3pxcE+g3Yxxxgfp1OaqLe
OnsZQmo1WkDITIMZBt0TlgLzXtdkp9t/LBYf1QmDPellvuNjAAbHN5RevoGxje3X
aknGnXDWyyhr3lI9g5hVxCsxfc51abJ4xQ83rRexfeSUBscALIk2Dixw3CJ78ujz
fJ22jC9Q9JOQQi31Hi4pHIfnJ7tnkAFXmJmQrGHgAdo7a9XC2vCMQuBi6UCIL7nx
tdGtQo/dIykMX1WWdHwQ/TzeXahU0VzPt1HG1dsMpMakvYmhDon68G+0b76nS9v+
rHI3P+DJ9f3dgHYY0Rvx3lTGIXsRSZC7ZzYvNrxkPETomkXhfPcF2lAgxKEB0cuw
Id2Bro7lqBOQUAGi1IYFb55j/Z9BgzgXgM0gzO2Gmp17axIG5AnzQV1hKQACcZ+F
+nxE//s+jhvJclXS7dP4MWxzV8YiQhgdfT2Gl734EFWZtAfejiXmamta9N7NLQ+9
1OskdJapCdPLm2hBTbgm1dT88EywI8W8nNMQOp1OtEZKEoiayF3pPl/kL0a9gkHx
mCJG1ykZAJ/Nc5GkLaOqLUwHQkeIfMV5R45IZf0afKcgPhZjQXedZ9ktI1sxv29s
12WVPTsuBJqecDcJVIpCkDbcONPx9cGxQLL610kl6/NhBqokjrJV1HEk/BtnhCiS
gFwKRmSoQ2onmslvop6HhukQQjiUCnvn0Fn7vLem/ahvDGnfxuSglegW/QI1uepI
LX03Use56EHOiy/iJ6BVzJvTiOIApjc83FvScVqaZkeWKbjTmCjr7u0H2oMqNbnd
5El3/Vep8wZ7DzDi1YiLXoXQaUMbDfvDXx7OIUCDucAUA1H8+YYLOou19eB3y0u8
oHePopd09xmJE3D+AjNpNXpUkiaFAdms8PQq8CIY7qYJmLNMJCUNcWloQoXpZzzB
gQuyuIG+Hj3yAY5xFzrJqoIIg5N1UzCSiUWfbyJwV9Em0azf2oDsYsqFkLFrhg7Y
pFisIs/T2Eqh2oJRackNEIuMYjmc3ho+tcX6kJebQdGImmDRGyb0Qk+r3FMlm2sF
MaNi+qzxp4zACyQiGDmzbNq5+q8sPNoAuKJdvgQcjA+0WLbp+kbJIuEtNKSioJGo
o9P2FshVKatFZbikd0tzl2bFc5fqmHZAFCtD1VomCu7VANcMkdN9PNwaAxz1i9e+
SyZgy9mqnS4Q25PLdzPEC82FtQo+C0RTaiQ2ivuylRIjw2nWC3rP6gwe9oLXKF+A
mmMKGwkodIg/dUkzPvC6WozKqemMGr8boFJGS8CksgToPFjHLTWLJWuWrhiRnSUO
yR7G+xAPRaAh6AEYISo/COAKf1rLOCysHUCp/Uk7vlYSyb96tZ4TC01SbmHh6rav
Yr7wCrzIVGf7Zm4iBBdV+K9Sn4xlsKSRNfPYwB8Yi5P/wGajXEipArPWxxXg9+70
zjfra8f+QW3QcoDGzKnvUmSv5DqY3ZRIB+XsLBMR9lnSXNnBje2MfUlyOCopNyhE
gopNR2D7ZPzzKukHDgmMRCTkYyHyG3XvSMltAcjVFgduOjTEBmDWSaU7l2BLKML8
ZryGr31Xzm0uGeTq3hYSj9OakVtpY1M0+lK9SmHJliUKUUfluxqOnI2gpiSsswcL
D1qUGZ1gpgEsduzPnrukjQcIaYOitdw5eQC4Mi1eOOMrB4XRacOeC9OOwAv+lELh
Sbi+r6mWeIc9bDiQt0yrz46ja7zz8eHqblp1jhD0snd6UESh8msVt9EEeXt6aSGc
0GaxWxpcpJuXbAWZLn6VH6TrTFyqYyKOWYoTSisA8VVFPNFv82HZlNaSFGaN3cXF
ru6oN1xv/H4lHsNgKZa2aLII96WGjWJASkb+idLk3G7WfTo6fgqaPuAMjwPhyitz
jyOWA/wkNp9TDPE/7w+h2fLxfqB3qWd/9QyJxe2nzfU4Rr7z8fN8bCzH8GOFreVk
/UCZOF/aoqqyfXMXGh/nMsPiQH8LNQpicZSMv48mGOTE7JhwI+HahjrOMsvVxdNp
BTeZ6xOnVdKSo+xs6KfG9PrwERETkRaiuYNJbh9c4jfqfTj+AU4YGN1KjCFSBmWj
Lh2cBGFeufNEElE09Q+Ro2YfS9FDpLhMeyu5B1YuXpkyyTJtGKId+mTBYQ/GhCmv
T+7O4E2+eT2ImN8EN1sM8I1acnro4Faipj/cv2DuqwhPFsi4JMrnL467gvSf5KNV
YioXBa4d+LIHaG9A7JJJWiLAxw8wyHa1saSoM8cR9E+dvZdTJd/qcFOrww8VOAhj
9yEfhMGNZbAbrrOTqDBF1/PWWCr+l6AF/SaiUWkKR5GeEuqY82tUCrpqORLwo2um
4I0ltxkCjk9kvM8aoT9DmoP3yTqj+o8niqS9ujVIbsmgRW+cDL27x84yq5vRFJZK
lXh1q9wd6B/8yPYU/y1iJ7EtNVeOGf9LsFB7/yfAx5IUQ8897KSUcImJGW8dvzGW
UfEMz7YG7V+HbZ7tYgcbRbhPYHIlEZlM46un7sLKP4pTrTQCdXfpX2Dsd358rgSo
cbauKhXIMDCcmWaDTy+xiT4Dd2n6YcFctpIbb7/hsOnWIz34U+VpQMQtSEzRc2kJ
fGJ3SRpbWhCbF8zJxwo7tbWfTHp8VnBTzmjPmuM4gLnhGq7n6RPITbp9n9FpQyHH
LS8SmwlAXuCCGQVkl6pzkdfsqZTOlM0nfWfhHhDvQ9WYOiPC5UNJXk947l8phyUa
kYIlxwC9O4BiCrSKe5INP8ov24m54YnnQaSfCfI5X5/6LqgYjkvHYG2QN4Gk8Z6M
UszPF3+lYtNj0aZfloenKQrt0tr1HpRlxUVpOpyVeMbBtsR3mOz4u89NUSJWYVpO
NQkUGlt/3Ji7VX38WdpgRyhPCznEhrWBC3ZtxsWVv+WM4Hg5/5Yj4HQP3lih03bH
M0qB/9cxJPN2xsJNjfjKSoBo4XZAzuWY239Z92fZax3R+LeRyCmZ5aGKOdfWqt0F
kl+WnKNRlybWkuwUfIBdpvLPNZbTW/Uxv6fg1Axng/2HnivKfubotMjyOSsqj9PL
gyQxlFUp5xCfDBCCmmuEh72HbHWZpAD33gTYb991GmzlMITyhARYrqGfYawWHJRH
D52dJQjaTPJKymMHXdufCp0Z1bIwQoQSGhqcDdMwuRLTNEvTRA3BIHe8Z9PPY0zY
UmX4giwr9SrbjPZO8kEsxoI3iBNMpfD0FNh27n7vjVRfkMXDNJgu3m42etIO4D9d
F4ht+XLyxWlrhdA0D7u0umQdlbOLvD64pMsde9+x6kYwKOwAEfY615Ip7+utSpwz
RgO1TpvKgG5iybtB9KJzkLwRndNzpwC6NRSgCHOA5ndjUs7oXDiVaHR1x0QaFeFe
mW5UO5+aeq8j4xCaHRcgeBH9F3Oe0IOFgDTQDfIIO+ynxvoBPfFRxBHa6TTk0Kr8
8kK4SNHgIYLUq4OLYLNk2wqW+fzNNGSolnFKbDOlCGdhX3M5/FSfDTYPeVqLe0av
PpCByHOlOlfWA9l8UZZsyZbe3IMYv9TO/RFu/I2euj3czBMjzVS4nbO8jhzJWiqu
8EC4EIiDzOEkYlEPoVpj4cRxtYo7aXkjAH4UqpAYNTpmBy2l522P0JdNsewl7HC2
Rc3NBaeQbc7vfxMVApa8cJgvGF5XzOzBp4ZnhnNPi5pxs1iBAZU6e9tJxMkzWZAd
oKdDgt7p29pNyJsKokGpX260JWopWzf3S0bKyG0vlvGbZSf+XDq4aG5BoUBivLYI
AWiGzi6AP/PxRLs8O8B9D1fOLagaOplZ6YTKL1CWrMYaZhjq1WjgN5azFkSLz64v
E5tUlF29tcRGsr3A2axs5vKZUPBP4r7jgb6j1sXSuxzCuo24sou11c4z5GeI19eP
vm75fiaUHMB5HaoqVJQUdeKy7CUKD3wyEPoDy5fkse3ViW0C9CmICSsJmD7spKeM
w67nLSFd7gzOiFRIypcPv35FgjfUtyR7+WIZ8CigBX2ZFhSmNWEUpAbu8pHnLF/c
vSby7dF5XflGlrGp4mCAcpeKPUdNn7T/+Hc/ffLgt9u6XEfe7GENEQd7dqcSwsTj
tZ4dQUP/pDg13NmBNq95erlp5lBHjZROBsJOmC7tsfUJunjNCO5u6eXRMdN17lPd
viMXmVUKxgD1N6StRJd+bJiS06cgJObgnNtSoVr52umsED/+7PYw7+n/eZiQg1Sd
qj7fpYuA0eKCrf6GwYiVey9YwuItxFJ9+s1oEz/tKR3SyoJu2hAdVzGaWCiDBJHP
85Jb2/NR74HVrK595BgDxoqHJ9h6OcjA241OKziki6dgD7Xe2kiVLms7MZkDmByk
iDqPBBOmwl1SOdgtB5AUMnikv3qxsXlL23t3mG8wTbQRMjqeV0F7H0phXudcQPKo
GeM+TJvqkweOt9BD2+GXph5GVdeU7AtwSIw7MxjkRWGazEG/5tO0EMNNgGVcdRpX
AZMe1pwtGrckMxPCxjtPe/226Td0ol40wKOIMz5WmioLUEeTfmE6MvFou5tHZGiW
oIRGIMyjLcLC9XJ9so1yTTjZFh1Z93/iTUqgMM1N7QD3FJhrmxnIZcLg8hqu2J4Z
vRsDKt9+5Q4USt+A4YaYhMGgk9C6XlOIl2Zyptt5phN1dugicoXBixdO+3E5U9TQ
PqPA45GI28HZZcwRLDJA/kgVzZE6y953GWmxGAxjqviBqDGMtRkAnwHhMAM3dPeq
/otNs70Vb50yi/NMEmX9/zc9rlOVEvbtGivHcwGhv7rGZzR1X7vcTmwXMfVODD2U
/D3QQMfdUPPWabXNtj2NndA5so97WVg1snrCh20/7M0MK2BDLrpXId6GfT6Fy6uw
wyYb/NYF3Xds65KQJ2hzW3rVTGGdOqXh/nKy1MaGo6rqL9gc39R/q2hSFBH84+s4
6D5LonTKXp8FesD7nv1eVoNRLDcEYhDg2dsIJkHhpoPEcVUtSJCxoS+5YJrFw6oT
dcwMDyOvgoURR8UGzZNvAb3cumiTkV4FE9vEpk/L7/soEBZbj6Foi27EC9IRQ35O
9EZK5jJOdMArVs8BG/d6Q83iTtmJQ3uH4YyK4GQ3wlvgiLW/1gWiTR6WLoyv0/yF
GpnJayQbPlL8g4WFW1Hke0XQxLDQHssWXhwhtDyMrdnbq9w1awSrBq0/rJ04N8wa
+r/gNPr/P/kXtboFYT5JMlLgsPxd9yn4FgB0iyNSD9upMHx/IPE5Tm2juWwT+l5f
Hu9K6WtvxVYnYH08X8KucTLCxkrwrCU846L6Hm5K5TiUG8+tqETyuI/pTwOvSezO
bNyRjDCqGzHFL+ydTh1p+r5OZmBpz/YdLENdQZdT1Ie/dsvihLl0XhlfBZ2fDthD
MBsimchfzrlyDKaCBdS4NYbmhCmUy7JyEgU9D1UtNtIR3ZJ0Q8dCPRaZrsudZcsc
CIIFU2FPVCiYTF7AIwfF34O3/OIchgn/sIh86rMHk8OhE785PZs62rpaDy8747G7
LV5aUszuTvSF/ZEB2AJ9/MsRsBmk80uyB6Qbx2lw/PIHGCGkE1FTxF0A9GfXkElC
5sxLXFRIvSqQVXdaMJQY2H6/xD00VqpYA0wlkFZG+QqpZqUqibpLp7FgFJHBv7qC
ZzrlHMbDWDyhQn43EBgXUoqef7IQB2RbkI2Oa+xG2F/W1Ys6zxZtITY0Pvngn4h3
F9ym7AreCa14VruxaR5SNCz+OvcLPOZOn0doPSf+mVP0ZQGSGM4ZNfr60OI5a8b+
ZyTyUptlLoTkYAyQurCebTO+3sQR2eCL0Eoh1Nf9C3J/SviAVey20b8fYGOm+xqh
jwDrkCPGWv9kXJk9ciXomK7zljOY/5/c4S6Jqs4CL4sP0B/OHhoecOgRVGrCtaPV
hZlG0HB8mcHWZ4JQccL9xxcaSsYbToPbWIPeetprgHT1J0EEuLz0WWxk+PSOCgWk
/fd8XkgkD7jEXKBK0NXGy6EMNysUarNKXPAd9pVi69ASGPAk7P9Zc06lkW5AapCB
plj0OhGk8Nbi+AkC6Au5V96e1ZAqVUriTpocHQMClvhfV4cQsOCeW/hOkBZFRU8j
oz2R4bLTDDgw/09g+me8woZ1e45Rl7pFMrolAElJcyYirT1eiKd8hMi+XuBZ/M7L
hmQOKbbJ1JF/GL8/9Wbsdl47sTPyv119vYpEBAohNxBM7lQ/ukilDOBBCYyEzJN1
pHPtHJsz2Tg4+MDb/tqA900CLdVgrHGdSBzgaQTzTHFBV/+SSM7LHydTY38Km7uS
Za4DBeBHQmLCinF4XflZVf+QbnD9SLyTqQG+peLNyqkY5TXFbc7Z9vw038lE4EYs
1TcknGcyvrFQRUGvtZdbPRfNpJcBXnI4a8juBKkq99pa4xBgtQDnMOvU8DpgGW4t
6BR6qWLcl+F/seXEVEXctqZJUpkXwkslGwwjR5M8TgU5aMKgJeMtxFdrtoBuenXa
y6B0gvC7NxQ7SU5c4ELF2OkqexZoMStmI5snbVmx5XvjL6WHZGHBIDDW9bqWq6jb
zZTf5v+NhWEs3/ptXXv6c1vv1ueGT8jTwR2r2w7RvQSv0F9HlLZrjXC679xm+Mlq
EvQ31HXH1z4TJlvAYuGtfGj4Bl8IBeAbsIFCu835ZRNa7YPxMr244bDbtPJN3Etk
Hoba0dXBb7waBoBxTlIYtF5Gf6D83+cmEVevnL9UtdpfKRzlHZrJ4Uhykdf5MpdL
Q1fy/auorFQ76KEP4XCVx5GdKtUOe5afLnpimYd3xqI0IQRPYJ6f3/PGyfLsWzmC
0v5Xj4huyvseUq1fi77RiZrRdzWRLVo7xqHsLPud0rNxQc5vpZgEgzvQim0pLQfC
mOl/Kr+Cry/e9htjy/ndUZPjUsJKI1yXItDNssL+QGgdVb3byxhelASNxTiHZphT
UVS8qZyFolUEPn8W/kviHqkzdCGSOt4u+HQ/ZwoHyFG0CYpmO1eq3Fr1Iz36iPva
sMNsbBiDe2ivFB38SzuypuzSaUDkypVV1EZoHOXV/lKh2ulkJYi3Mqyvpg29ethN
gaZqG5Y6vdSCR4zYz6RahL/QfSQBGhdlvUhxlZAjKggc2HNU9IYlhOpX21uYRw6y
QHarao3TxZwRcCrWalIMSxxdObFIijLyWlDA5wQOl+h7iNdHUo3u//J2RtNEylsl
NQI+0ZPeyA9Bdsy5bltChLfYlL7POb8mwU0WpwUL4lzEJLb+8wxVALYjpbKnCH2u
EAEMbF0jJhW9zJ+FIYX7IFRe0fsLpgW6SbixeqpDEi6F83mX1G20Vq9FDcWm0CRx
QzhrGT/Y2uavOI95VFxAzSl8mJ2gc0V8AVjqMbsCp3OLafBNiP8HOrk44cO2D5TV
r8/hfjT+X8cetZRgbVz+Ac3UI2oqC6WJrAwCRR7MmUccIaDy94NWBso7FeOi891j
dMGdU0akqgoDREKYCTN/T4RMmqSd5Ky44ItMABpfu/qURW9lp14sDaxLTWfJa4xz
fdtFI/jwxopk4PtX53voTxHupGqm1K4mp9xx0GlJ/Mfv8JpgSy7t0/K8Ax+QmdS2
KPDtzeQnzUQi/LVMFxIfyV6HlwOgexcL1spuiwV/gXY98flNqimbgqXeXMsihq4+
DFAokV7GO6YJEdLwlr0khuu2GRcYFNcwYzEtikpQ3eV/uPfVIZeFlRi5G6q6xST3
01oSO2iD4Yiotum3nd02mTbECj4CdoMq8MySHqYPoxW9jE9yJsG53GWLn9HbzrXK
MaSLfCTdKshEWco9Nc2lBDw9zS2kMm2qInTt6OxKo3sgYa03d/h9pn+zTLNWAejn
gsCe/BmgehfVAeI7x/M8aGjaxE3H3pW52w4Y7noJBmhq1zeIoo99sPdXtDG5sqFi
ayFrHe9xS9/yyDGsOi899unrKhJEnMPFOHkMlqbqSxQnPFBM58NL1arhRCenlMrH
VLy02Afyhz2uyhlRkqwpXstAMQ+5DtZaV3pYqMX9jOB/EctQm9pSMgAc67V8lqSo
M2divP35i90u6zRKutEngw5rR1I+w8/PdEyULOu05wAopClX+Wzq3XzAEKazRFst
hmr8D6SBVlRAyOykVsJnjnimKsxmTtuhmhNnGmPnbeL72L3oQh+Qu1xHTPDrfXCw
uprgLsGohv/uyr459D+NuC5gfZfKa/s8ZDLQubulOpdPIA0Nps4VvKWefHMBmiwH
7XrcEB0O+Usd5D9hI6qJhajRiz/DNqf2a5L0btj4kG3jrqkG3/v34KbDJW2iu0KW
ynYlBRvHB9dh4vaknKZTVwhUuDgtsr7/U6mat31nd6HM3iltdE/JBrM3YXr9y8+k
3HmuXbHLpCgo2ARP6XSTXMfPHmgMqfcMbYMCzdVyn9tsjgWe2ysmzcA6D5n9SUT2
zC0j4WSsruX3OghKeFGLyoaiKTg4U+FoNWmMm6Lro85TrOzTw6Qj//l3VcmZOqKA
CznRtKQbkaKhPrM+ACQ0LamKq9AlsTS+3k+wOlZvjkg2S2yVm8SWQ7He4KZajU+2
tvodiLO+4LeIxJE6+A0sqyEpjr5mQKG0zTSJncJ6qQaEKYBMPgq9KfeEm+SB+XI0
dRjoX+uY6cHkBMW4UK6BB0wASxook/0+IDSZ3eDJXj2V3/xgfDjBhAoHz7CUTLZg
25UJcC+w+N60GRqCn/L5QajEUtQSthzCGNNH1PHyuf8h16eZdDjfgwvN0aaTbs3s
q4cCq4dThQObkO/MxBjdZbKobDEet5ZcTJ40s+X19SLEpM8ZRxG506UW+mTT66ht
ETZMIpBIPvjy/90ybUyJPwLedFpHYKOIRCzPHrysFYlVmeNmJXaijdZFcRf2y0Gm
t0r1cYOldBteCY1H5MmgUSjqk5xFqjzCTP48lnVmVydxHQaunnjpF0qDQSzT48v2
MCyl4y2v55uxXqEWFmOzfZYPXq9JV/1n4pBOg6DUPhLaflVlxOkQ2/QUK1nLPU/e
nPzlMXv+0QMxv9lMiWV02LN5/6QUl+YuHVRGd62opq/SQIlF2CErqEelfMTCOEwu
LRRXbU1eTagDVrQmpBC8iFxMgR1INcK4CeKAEoTTguw9HeqnsDSJyYtsAyA+obph
UssxWklquv/5QWYM37iB3FTY3tSSQCY1r6rIC+VlIHNqCXDGa8Kmql6wk2uIcXug
NSaivQX+fUR1p0fbZeeTDIJIpYBWb8+7Une+EKX0WamrDu4aj+Aqe891jo5ZUKBn
8G7iPp2gELXGFYcbLqaFyT8ZnYcEQFYjD/YE91oy+IQ1/sEgzpUcKj/NxCBZ8/pf
4X7ukNhSnPWgwM4rh25k4ySFKzxFV0GxrlNKG5CLyHr9GD9k3iHOn6muq2t7FXd8
jaKaUn4ySK+gwCxpMw9L/jJK1M7h56Bmt5vz2xHGS+I=
`protect END_PROTECTED
