`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WgeXocnUMu5ddsxd6ovEyG1ZKJ5lRclxdQIKpTLNFT6v/98QqJMW7LVatfUXC5cq
d+fVptywZCW4Hfa2HkWIiqmFg3Tn/9UVfJy0Y8Zd4Y5fSCJ1+552oWI6X8BvPibL
Pv1Os/sYkxVvEXjBn/LCB5ZZTVNtNUq45OXTY2flgjpB9o3IH4sAPXOv/GtdK4Ix
jqPgpfm7++C8i0dM0gb/0DsdXKAgCxeoJmjETl78hE4mRMXyKvbRAJuQeupGSZfO
d1tPjgxYImlICM2ZvUc/lpCAkOxLcMKTW0KU1WxHJ4bseWYlEH2EFxScjsuGNV3a
J4GUFGyinWo6xO9rUWqaE0SrjDtQ6q7Hgy8DMesU+z3I6dl/r/PkAzC7vNDMsu7N
yvehLg/S7raotKHoMVaCBKfci8ITpODy/lk/GBfWd7Q3u88v+b8fj8We10hJXoKb
+NdulUtlO+DribQUvcmt0cx5tBPdIl2QyUbpsum0urfv3OwcWnLjn3NuIpy/OVBx
ESdg13HckhgdiHKhg16umHXqoRPUZmhTlV+OfbHuN2r4EOsaLhqijIBzwHzicZMA
0s9tQJJ2STwnFNIh0als7Bb2esMD8TIO00++ftv5xMcOEtf88aia+6YcN2De+bi+
CmEecLZ/mVo3FjIe2Ju7QjbFo5R12W2YJFuycUwmcYy3+R4U0IILOxHvBEnj8IwV
FiagEn0VN26AGmY7L1eRdhHjDnUDwRmIyhA7keLtbNb8sktC7enICUrqgieh0DFL
3nCezfMVhPIIo67Hq+RJna4YfHlOGB3gdECB5kJpcruuvXzrZANo5LSKr+tXiZtA
fetkdJuKg5z/NiAF2Cuqk/yokXsNanH7n3HuI4Vk2eGA2tCRshFkpWz7Jus/i4se
`protect END_PROTECTED
