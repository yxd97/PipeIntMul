`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cu6DvJY6aTptWMYF7Maj9ztliOr/CZVHAOw+dv4ZbRZExOC1lmz6YPDlF627hPC7
/49IiOJg41D8oWApTrGZewfzLukUHAEuzOssDTe1HwOqQLce0xtunueyOlcUv2jR
ORCucLSA+OzVwJYCSZ7nfNtZUTq0aX9t+e/egMrhnjkJwvQcglXaeEXTZ91SWhTt
PBvi7XDpslERFnDtTiDlqkFng5ufKpW/GJ+cPO8oRRebOEssefm0s+ZlSHYKiEUi
O9kLba8NMFU8pbuifWn7XXnMMFW8UX58fMpQC1dmlsOjv1FeWkn5NrYv9pLcdSFR
C1zA4Xlb1CC23CnENdO3srrZ/Nua58xvEN2NvC8jZVDm2zogedhTSjunRmLc8/qB
W/PktS4flkMqBs53vw6qx2LCYXnEwPE8DmqV/e8DyvNkEyzLmNh+rM2pRAzh5y7u
I92o/By7L8E/Qt/uVmz4yn8m2rLouXW5eNsayensnEZsDLz5Qy1UUPKtLz1EePln
u8FixfACTD7hcY6OqduOKDFpoAMvUAuUkoNiRmohghTmQwTFusQ2IiYwzxreGoGx
gJog9i+eIUOVwCBYOEkFs9AB+J8qfar2I/6UgeIo69NOA0e+vX6sOrTwXdIGPvcL
uSJRe3yVHDGuFPWsApHRwdB9os3kGgETurURdM9fiZU=
`protect END_PROTECTED
