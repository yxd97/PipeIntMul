`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHeEiCL2vAW/tfa0LOtf+CTVFdqJY2rqBkF5e4F3FYLcKAfoWN3HsJCRJ3qx6LUo
UrToEhSFMegE/kQNUNKq+XiWpDT0gQ1SYnnOCM0h7hS7FyngfLeMtK9vCvKcgcRc
xjTpt4o3DlHW1Cli19l2ho2pOB6R2Rr2wPM7l6HLrryS166YSJwWqd0ztGbHnY6q
usIer9Hb3BQt1D1rTAKBi0RwBXGnBApTknIySx+Inf22OmS7BlJ5eOWSYcS54PTm
rImtY6vNd+YIufWdAYVRRdwkv7nFx5u2OcuY8lKFwc7Q88fVtgj9oXK1MS9fux2r
plAx6VKGtFgwx9QiVkOFnZBG275Z4FOJz6RMv6aaQhhpJDHYxQm8JIz+ZvQWA6No
96uHD5loF28FHuptgJAGsLIyPlqHrYaUh+VTUyQzWZ80Qf92dQmMM5cnes7H6pWi
Cjq48fJEHXGUdcmPz2GpLw==
`protect END_PROTECTED
