`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zH0X9tQm/D2ULl1f6qs0F3JGDgKkANvnYY425ymN7h1AKoP4vliM/f4dvabwUr9N
CrvfXXGhM0efFK+9QjvnvU3Dgn43rPcDDatbJ5t6A4+BFDfhw9qtLho+IjRXlcQW
CPmeENNEVcF0x8n661Q94F+P6Gtpqh5xhXnSW6lnvNAgtGw8EeOL6cPGMBoDduhs
GznY+tYJOYDoLtkmoUOiMwfy9cl2iSBBiXoojARQstTxO5H3f7g4UkHBIHZp4Lr3
FrIAlTDkp8FvyePWXO1mEBA+TlpoJ0TX7BhmGpT5tuC8Z5X7qTJ9vQQvGyvGuUmK
nuOLDlHUchuzwi5KVK41u1iX18fx/4vix0UnTJ0po2IFLbprSG1RE6vDiqlrGMXu
qfdCpevVtKnzxU3YuPwFSyie5bgFuN2PnAX5lD8PjvLnABJqL/vyU9aE8tVxYVLy
ytDkR1lseeeD5v3JK0Sk4NowrUVCOxx32FBErUmi0vIO599sP/hv8dvKgtdDxJXp
`protect END_PROTECTED
