`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqYX33jP7TC5D1c6yWakx10w79Ia7ulF1u6FxHUVTUPTuIMuhbDOKlo4sOzGTKMa
Jpr6F2AvbeLLT/e4e14EMGzC0NdMqqj3ySSAHLJNghG7m2euFtWY5SsXBeQh0TFx
GhZ/USIThcyKXfSLaFuit4+V6o9Kw+ydNjkm6Aq6cfRfYIAeN+EngpmQOshlNtIY
3xUaQ8NMcSCV14H8Cylj1Ol2uNB00copGyUIjOymHpqxqE2nPIk+dq0ngO+jVHjV
I1zbf0SY+iFWslhNpqIoKCunKs7dE10N9wnEpsjDaT4=
`protect END_PROTECTED
