`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCHJvvOcxPfOl1D1oVTE4BHQFk8KHPsMO2lMRxiPvy5XFUh7NGlTWO01cNFGE4Fb
o1xZbOoHu11Q9BGpJkIldNrgrp/CDBFDlsn55KO3Q5juf7OQslKg1s7cB3nsFnYO
YtHUPjNWwn8ZNeIEBeLczVU6Pj6EwiL4tqejsWxxlL2OON7dHre2KeXSbveEXkAV
dE4qbj4NcmcklZLbDmZl0wYK9nOj2EfAtFjLIUl4PH27qu+CyhfRHJ/Wi9mQdYdN
y14/RGZi8vfzDmkOD3RDcxuSqtwzbmu8mYNwYLWVUO8NEuIx6NlWlVa2eNDGFLQ9
axe2TuiZMLzYxw66/m+d0eXSV0ORNwzKcULt1A2pwx6hyNBdW23X90saPciMUW9q
MXZLEuVkUBNG0E89Z3MDE8pyjFXBCyav8l+cSl3wN+br51mmYlF/rHhMr7FJHxOJ
`protect END_PROTECTED
