`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vwNu0oKe4Ur9h6ehHGpKKRRrpyRJbN4paWA5WL9oYPaf0/X+4/voQrFHMKXftH0+
0QlZAiNYKI+4GGD4AX2Ul4+1RbPU8XuBFJdQEPkHndeqfLtYOQhk9/NIi1ZpVHDE
JA+k0J8EoQnPKM2UCFjBoK/TVrUyBi/wWTOWxlbutlpNtbcd6Mh+BC5joFgRwu/4
JQDQFfHjWA8ngAeqzQyz4kQGfQOA/3DiDCrnylHvVi3Gw1V1ryVD4ZaY/VtA4SU9
zPCfa67L/QsoOxaY2+iErek0s85Fnj0bj1xObck+N+R+zXtYZhiGtdK24PqGrKaX
KPfdy7oNC1Df6xPp8mJy2BoAq3Ee1PB0HR/odFmfV2INVIqGaZR1C7rJ3DJwJVC2
+pxtOVCwLWSNa9vF2ToLzBMnfhPU8nAdXulHEDu1vT7Nuwn+AtxTzzHqxsEaBaMM
EyjcM6HppR7gZ8P3OA9PlE0eXT/6Wuw/qggZ6bZGJuzUevMZ+0Y1fsoqM3EdpWhE
t150IatLv2/zNSH7pizYKt4yZlQ6I61jTSsJlE99S8lQZYrjHFOMuG/U2P5hoXQs
rQY7FxIq44PaJMlLH50NMYNs4LFVXwfnuSy16n0uQCV/eappEc9XqRgypNni4FdB
90/Fc48g7kZT7OFO7uf229e5BvGa/rBBfB3flY5ze25CD7kGR3Zcg8hbzRLcuYb/
L8i1dgfs7n5s0s+kCLEY3dTDAwqnUQuTgoSS3+040pjWJFaeKevob7I8ugvEH0e+
fH/XArSVZahgNiOiNzs3I7L7IGTRH0L/JENpvT/q8iH2NoMYjZYZVqXQAVPVvJby
D5R1JHzPw7bQtynD0QHzVTOtRzhaKG+xTefBI2nP9PkMw+7jM+adGYH3WEV9nIqE
8GYpleeROepSpSMOq8PT6XcewVjCso8NEM8IMjlGKur5gPn/ZJlK6dH9tswFl+Fr
4v3iv+uGTidMkqSVR/4m1zoyVG2CaAGdhfkIvNSMXFnr1SgWV/B/mzcafGqmt0IV
+xyydCsDMbvfeR6fBFUL0I+5NfcB8HcD01KW/96xNoNX0FW0zhxspQgdE9FBPMog
+Yh/p8cbgT9OQdfl4ltWEg==
`protect END_PROTECTED
