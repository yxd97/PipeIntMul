`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v9mKUsJiwf3f3siPiZE4jIQlYhS6vRlkhQUpsDXgxLCNegsfx0Fe5zEM6oHnYiWb
zAbxlVlOVdY3VMZ4Hryo1AiuEtvTMQk/A2AhfkA0jRHRxlAkHjh2T7tmPznnt4iV
jFFm3u7NVPZLLie2EAurJxuVq3QjCvlfWCMmgSJLMAW+Xc3crML3FrlZli5/P/9Z
fjfY6MljD4NyecUNO9sqIMljvbC7s8iWLYL8zgH63EG3biHyhu7YFuaCt7bbb8c6
5kj27B3fEQIjNuHqtnOVMQCQH/NvR6zoiLv0HbQftMQOxiMCf8WQ0LOkDCa5Z6Hk
n+rLOIvpLuiDPMTorCWdg07suP0DOyFW38SiS7t9WaxufEKFie/voMrRqEz0sYMJ
u/7i3hjpDILjuWpvMlKLykrVtI7ZTKyQkOs5KTQSIUfzJAw5aYjkIZhkCuzfaOac
GzbI0j8NtXyFKTb/yeQfpDDAlMnZCYD+yHhYst+KeBg1A72/uVbfl+TXZ4jEYokY
`protect END_PROTECTED
