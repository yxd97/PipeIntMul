`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8kZUmoFKtVbHf6iFhN4H+1c6Zf7hvx4Y0DdkfXV03TsJcV7aYf/GbAJcH7SO1h70
8ayjyDm0E+OVmEOhMO3kWCOIqmNY/7wCh0L40KG2oOs4keCtCC6J2PN06b+QgjVb
IR1vvaq/kUgMQwv5kGqFNha1qRfJt8ZY9ik8Nz3eim8bKTPd4+kJ0MdvTutrcTny
aT6rdqi7E+tLKe8bwq6VA88TzIl6owzhR1IYwT5kCHujLohhGq0Wq1bKvmRWZcPN
kRqj3zW3n11U7jgVQ9O4BNOXb1oqAmRwQSFd9aOUXySPCYthwCw+kE5Hny2JyrEC
qlFAt84nktRLrdFd4mQ+EFdGibL1/cYVrZtP1AaT/7FtAqN902RApI78C7NIpAQp
H4cEI3oOdUyy3Wji+UmpJQ==
`protect END_PROTECTED
