`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxKWA+v4PtzOZ2Yg+OBQI+EYrXunraJyeobnzz7RP1lw0X7sYqIJkRohQvbhqjDp
r4zzg191dfuC7hjevqMUgw1MhF37L4yjOQt3MYkLyHxYj0/Dd5yJLpMBFdOlX1cu
lrfzr9xnrM5n0qfs6mv6EkJT/03H0lYcIV2c8HY9ANEgtOEk5UOmYCkUNIMLIHNc
FDBRbU/nPXoxFV8fjFNifEMhBhltB28GTwIMJd1hH7QI1eOKcuuSNbEKPxJiDkWB
jlA95+iBHgQSaGFgT6DMDkxSzUz31jk01tUvrtD7dwwyJX2c9DFkmzHEszF2TyS9
6+58xOoJul2T27kzAMECAb6hWxcN4b7BFh5VmODkxABQrkaO6w8+8CxcaDMPz/cV
FjqmdefG+EKsSB/WJM0Qbssgklwo1p4xAvMLwOY7yJc4NODHcLOj0a1Tp9pgcGWp
ay79wI+sRcSp/vdzcUjQWeF3ErTMFw+/VbtPHb8vEMGnwc6/95vFW1Dmeh2LTjX/
`protect END_PROTECTED
