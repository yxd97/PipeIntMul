`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ljoo/1nIRCzFcu93FFdFCq0ftokd7HDWnRTzK22d01iCZxa735jwa+NdNs9aO10j
CaNtDKrsOIIf5DRMsaXGk2mRVwbHDvwSGHgukGT5reuAxXMKRRl2+iEfEqjsvrPP
c3Ep3uSNI9qVbwziBvRYlyVvjxubor8DND84EnRKgmsFTBe5YA2IW770oY+JrLwo
2ujijpx+3GARkKYieOnKir85iVDpARlX8F2p/D2LrX/C+jfMily/AJvrqTyniqyE
+Yd3TadoRjY8XvE2wY7VKADmqxINAsax2cKdFGG4gJ2Qu5TgPDV4zn3nkVa4pvF0
0fn51uyXAmJUXUIuLVwHGR/h3Eoizd9IUCBfkLiyu5LEe/5MNLpfnmE6uwtFm/z7
3SesTamjyUN+x/7ayjZ/9AR1EdAu6nhtEQbG77IZFsITrqS3gJWqXhOO/HmfAUX2
jyaDyYoCJa2VRt8XPyLst96LxQx3RMc1yEJS9V6k+i4zNIdQVD5Zscu0Qh5dJoYe
L2ZAqAL4G8LpYmEx08z83vyoSGmyxCXIB7xOFoPevRmBrSk/bxgNCV2rLEBgeSV8
que2HPyaX3F5UThMKm4SOO/0m3awBaj3AQ5sbAPvQ1ajttPEHHPEAVcERrlyJc4i
1RIzu3Y+ez92UG7497z1jZZbmLy3qngX+0cx2z6/TwvqWeYOZmKPrnYnKt+2I//O
bSOfVOze7qQuu4KcCngHhZtyreeIa2hbBjek6tmT9E6jRn+Eb0Ejz130JpgpOYII
puSvR53J0lX9ZXUxhPuymI55V8GYCn6uaxN2e2Lh3PlGCAO//LcHAI/UlEnpIW9N
i0Vs1bWfRSM6XGC/H3ZnkGY/Bfj59bPrQT+LKlf+Z3AgQ1qteY6nHFvMXw35mUii
KuLtC+BGuSbzjZmbn3ry4/6XrrgmfnH9lybbfvwLO7A=
`protect END_PROTECTED
