`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FwcGz2hzH4MrtjPFfdFz14cisAUADDk1ZiFsBrRdRGyaoXSWkVleA26MCf2l2XRK
vRnjbPU70YcDdfcdT0d8n2YgAJALm9zjpckd4MMSYNSsnl2fvIsWlp55cwa+76JK
lSBFwj9wtcMl5hNZWLOl1ITbS3a4Vj+akK0SK8rljj5M5RgVQRd2VTjGj3GV6q2n
IcPLgfsa4nSk5soR8bhqzQIZZbOdivdgluD+B3eVYzS5b3xsi8gQ8KYrOxNLuXNB
i/TsGYLiiUrbODnaDq87rI2YFl0g6rvgiUhZ9Ytcil0CupJHgicH8rAGT5gG0XTu
5yKs04nQfFnceCNNuUSFdw==
`protect END_PROTECTED
