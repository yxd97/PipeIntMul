`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jX7YbkuQ2Gx2NPUKgM+XNsFkNIlhstUJCLQ7/L6lpMKK7mw+qCbam/1JM/gjT+HO
W636Hvb7/1ma9S/8IOS9mo6kJ72oFgg3Sr5Qj7HOi0FrLbD88q/G2+maz+GOtwkJ
KfGAjLsa+KT0N+VLY+VHNGwuuKG5f/QiWcCpQrOoYX21EaS+1Deof27YNmrrSLjt
UoYw4vfnmRYHFlU4c0PlWv6ySQhvdTRIg+z8z8/xC9T+bNRGS9FDD0scvDQK3z6M
tFbz2K5elSjaSGNLk1sg1kV+LHvjNxYuXLe17aT7u58KhRJZ0pcQCIDpCXp4o+Zu
r2Xvoh+XgCxC0d9jFzi8M6j/le2Byjg+UtcmwGPAuil66YYJHOU4f2uHgf8owuD9
Et/vklayBOh3EPTJ7TSqCPRIcPoqOEpsA9xjxKV8X662fRAQlMalgw2KEWwF+Ndg
NslIqJMQBF8U/Qy+FmwHYGKI/xDqWFRLrhZh6F2co3vMM65bwITWCAg2T1LuKLET
`protect END_PROTECTED
