`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
82PoxBQjuUHCzpNU7LRFr3WdPxM2ubOvu/00y4dSCRw6/37gTRxDcoqczH5VZPrr
m9hhZPk3YWrCfoIu8Qg9thcnsZB8NbW50ijTxjvHCvzetCWgUtO/38Oz/e6bndAp
qEVlX7e5HfGHeri8wDvlhIrJnS6W5T+rDoGyWWEh6mT17rd94n0jXjLOBHdWm/Gj
2letEdtcHRfYB2G3Yq5jMKwOSwHAHnAvztSj3OSIdg/yTDguwhuIJ5n707O5K6Hf
ou+B2HmJ3B/ovRcVjl2Hl3Wx2mXnodFSzen2DuXzHAQTGXZnyrf335nMZjPHMkvB
w2c5U2vol6232L5HPpQX4qkOjC7jdFjX5efm3OezAZ0oSsnFBbZGbWQBVAqCRVb/
XssGn7F1WSQLFEnE2p2F1aoedrUAIrRuA3yQ14VX/TQsgxJKGOg3l9ZK+fTVlOaA
qb1BMkuCFZQ39T/d8dcXGZOz4oObEXjMNxN72Oc3aR1ymMi9m1wSiuD90jiEewG9
ZAx3Ee90qIZ4k7iZ08iU+E+bw7Hvkdsh2tfkQCnVKrVYqQMX0jMhb80DDulYQaDS
+M/D4kdEcdLbATYN8mOby3IKX6pm+sik1TC5TWlDS7SC0KaQY2AHq35h9EHOFzqx
GBR1EeFMabtiWLbyzPWW1fu1ONme31X6cAmqXj7yLSw=
`protect END_PROTECTED
