`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
87o3qczWHDmJYMvkmd4eB5CP7Pm34Fnm6b+EfxLL0Im1PECTEy4ZHmRKBSF3SaWF
17cWmsBD/xCkD5oNgBhDjnQMDGeZk3IblNJJPDR9Hby6zD9eHFkQBAXFBgZ8CJkn
Lcyu2HkpSkCFJoezFtCfq7wgLncky7lry+ImSgQJ+sCV1W5E1JSUFCXtXJwfkhTR
jFJE7NHwR3f8Y7Q+u/JqcziVqST4Ml0VvFTOojaobypFhINSQdK7TKpEhRFqsQ8n
D6Nv4RpEAB1KhT+Jc13Sww==
`protect END_PROTECTED
