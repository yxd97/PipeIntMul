`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wrlkN+S2mkN/Ltx3F8Goo5QuIDlCTtp/doAhpsrkPHLvdhH2MXG7FmeSNuuPVmXw
Ehh3DOBADdwSwHgbVJaS5+fKrnH6ZCERIxaPaokRnFke4OA97IfMJ/5qZWF0L3iV
C6Ywdv9PQleLEtGytV0URpX8za4nQqbSJRdt1uWLde5P6YrcMw7sx34qJLDg0BUk
TAf1SKF/L44KPwPbrOq+3f4CGJMWtt2EVV95QQlaKb98yxCV8iehqo9vHMKSUhaO
uM50dEyYxxsCv14alIsHC/p5PzTCA2KKOOgg+Cl33s04uW7qZ7DErD35z46srDiG
ZeG/R6iutEsuhmobPqeOFg1mG7wf0ImM6DA9S+Vs+M0jzjdu7R12+GbeEboM9jzH
0/zc/Ob2F7fWit+n463ceUp/noYTsg8aHjnHTC90e8k9D/JNBOJaYdcwSuLbUlov
k4Z/XXUwlA3sRxtv++hBPqEAjXodvX5uMHUhw0JBKc0=
`protect END_PROTECTED
