`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SPabBQg9+8fVvZMAlSNRmdp8sI92fg+FDh0LEjyNHf9RC06d56slvfnDIH68OveI
gGxKkyZzhLk/0js+6qHGM1ex0LvAtcoeSkI/c+G0hBJlMygJEF7z6am42hj4SkSc
Ly8k4bA3vNh7hV2ySzz6g+opoRZxDzZLtF6+lIOp3YTJOhbNfLupXbQxdl0Ify5t
L9AATKlwNm+D1lE4JumnAu4kT21QcVW7lm85YqK/XzUvYjlG1MsyjiDU6lnqs6n2
QSJRfkcDPmC/QOzEIWisej3/x2wLB8QGH2xmF+m0V0hkL7iTx5sW3voK9jfRsMxz
GfLsMxXiJOJlUrGYb5d0JN8/SshPo8YSvRhnJFYrwRLUHTHcD2aEiUYyk7eOyqNf
`protect END_PROTECTED
