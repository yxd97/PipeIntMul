`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beuvQX8AV7LSZv47vwootwUahYs+tlKVw1t3ha95YNbk329GokMcdYPGVLcvc+5F
ZLYdITHyA6thoXiR0HMSjc7bT9ng5q9hQqAF4+VyobvrCOArBtO2G61PwAi46C3B
5wVOG7tXBxHG4NSjyCgwc3HorRAPlkW1Ot8oGZbEOIh+ybYFXvfZAb6EXfSPgLEW
X6mqkaP1utCH+9mIlzaMYH947V9giScLwG7dbPHTPJ6i+jRQH4FbKvnqZFqre18u
so0ojWaQMOYyYF02AmMMeNc2Xddt1a1+bZEF+sMGcIMn6VTYaxZitCEcW4X9sA22
p43jKPY1H/CZWmyfmDhsQA==
`protect END_PROTECTED
