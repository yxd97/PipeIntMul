`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SH/ZByoJe+izaEp58H6vNVLscy3OcmUVHsl/d4U9sU1ucO5LUI1nJEcRMj910PjJ
ma1eRUx9oDGHJiKYWTL06UGoeTRjm+WqAt/CfCUAC9jPlWgYcdEXhF/7Pb255ODv
fjATPJ/4MUxAz9XaaEkL3W+gMnmDJ5eRKQtWI2878/wP9Prn3U3b5G1VvgzMfjz1
57G9rC6veBvM12ob+sYblmQ7dt2MzSggZmvztyBIgPDDHqRVHLzwp/NwomhAHS6g
3kTWvbWm9yJxM8lS/tUKEssyTUGCiu4ccM20L2CNekEyFtmPyN3P4RWFbav8333L
y84f2hIiLX0UNrfrEa18GyNZHp2ErSm5BKQ9k3pIYSp2PUkRZclTiSzCHwL3jxw/
YGEyj6ej1bJbDLKay0DBOGOaxV9qtj7T8ue6uijdQ90D6ciHpzMHp4jA7k9Hy++j
DQr/Svx/YfEpwKe+U1QnErdzaPH+GXkGIyxiN1Vxcf+urwPpWjiJ0Onaj5nMgKl4
JYmLgbZj4LUA2ntfFRCQWc8GGZK48Rokrw3JI30ZVWe8iCyT1we/p04rgCPDG40g
AIhknAPKtvRFXqak7F3r5bF0QM0RyT/XwaD6zjEO4sFXiTho0GWNvE6gtP0l3zvn
pl/I9mr9kwvddobwhf8OwLTE/IaJYybqdW5c8nDFk+azEC2gO/HHFh/s1ACV6Aiq
e4yJNla5hG1c9AeolBynDWM/t3E98DqcGOWXvXONrsPn9WQ/c7YJuBG6sw3GCYs3
OJa3+rTBMo987kNbgnUGI1YaHh0Njz05LS+eYbgq6f5fuHdptAzqvGx3GJuNB4a5
2sgeUv8Ty449jZ/+Oza1NZ7wKbDucIRB+NpVMtdQmk9+WWyaPm5wFCLXZEG7w8hV
sBkV9Fb6j/MTOyAG2hLMKXCzOAA3F1+MASj22fghqE30IYtII9MQ38ZK9up6H6FS
Rj0Y8PbpnYD0tDeWtiXxpJfIoT3mEncN6z45b19dUM7ssP3iQ+I2PcAYlXTXvBKZ
QZCyaa24yJFU9cekNjz7fNGvgttzOiPyHhsHV1Op+R+geI9KNclyqWf8ZdqHrjrl
LSec9EzBVbNKTrz0eWtGLVFyFyktyLrUtFMiivp/F2xhCRSH40qG0NQnbxQFsHGV
sF0GOVoO/bU7X/JRxNkjBHsqKI1LrFlMJ1QBOC4eza1fxvcpv5pPD4ulvrH9R3X+
LTuOVkfFmQT4/zaW/avJykxK66dTpLwGOFxtuw5Ef2Zq2Wpg8nwMl/VdJ/dU/YU1
+DZ4efCf/PknVZNkNDKZkIv6P3s5EgLMH/vjAAatwu6HnEx31teIRcuvLTtefgm3
zhEzos4vo25bckCNWQnu4fsVMBf1k5Wn9rBtFm+N7ee1noKzSdGoyvQEK3EYtFko
rFBEt/+LM9CQHwX+/bJ3JtulD1/jwUpsDyy+EYZzZpWeGO/IvqciKUOGjWYDsg8g
XkhoetNNQSnXISBSSXaea8LjtyFtE7IhnaBjylr6BVq9xrRy0D5I9RNKy55M9CsY
NPctO0HESJH1qoOikZRfQ682aZEuNziN8+4R/9yI40UGLMDcwLRMQ8hvrV3SSB6b
r5dYfo90nrAsEHpRQ75EpOJSayn6N2D6CSFYLRwgDMaR3bAvsiEGG+lUOyRCUNpA
KFbL7K+D/HE6MhH7wvb5siwpW1uf36N6kjfU6QuW3p8cS53kn3qO5yra8mPH/si1
pdzBCK+AobxuGMlErcoJ0ZEFM7ow54PD5bl9rMoEZ79WV3G0qLE3nP5ZqNlzt2bk
Ai0QjkcMuKKPJno1GbJH8eXVM/u0kgUA7D2q/eI3jT/A3mIiAWjUlbfq79gOwR30
/yKOKQ0ckICDCMF8L+T6UeEZPH1HwvRgFmuhlcF5bPkCn0USBcc8sFub8kKfxyJl
kh6IIgAzZbGBOXKrSDgJ32mGyvBA/nUKBHJkACDWiyaMv8Rlk0ivw9qxCKNifLNk
7c1zeyoKFOvS7/PxD4J4GXEOig2dgO3b7886xzjN1Xud2fHn3nvpKOl+fJu19Cw8
IQ1gsElqby+DvSudB1YBiT1fcVQLLzWgXCIYX+SJs+5osz1qikmLOOZQfpTCFa5H
NoCNlOQG9nS/t5IqOGd6sTKz4sK6E074RAqcMryAzAQ=
`protect END_PROTECTED
