library verilog;
use verilog.vl_types.all;
entity X_PCIE_2_0 is
    generic(
        LOC             : string  := "UNPLACED";
        AER_BASE_PTR    : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        AER_CAP_ECRC_CHECK_CAPABLE: string  := "FALSE";
        AER_CAP_ECRC_GEN_CAPABLE: string  := "FALSE";
        AER_CAP_ID      : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        AER_CAP_INT_MSG_NUM_MSI: vl_logic_vector(4 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0);
        AER_CAP_INT_MSG_NUM_MSIX: vl_logic_vector(4 downto 0) := (Hi1, Hi0, Hi1, Hi0, Hi1);
        AER_CAP_NEXTPTR : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        AER_CAP_ON      : string  := "FALSE";
        AER_CAP_PERMIT_ROOTERR_UPDATE: string  := "TRUE";
        AER_CAP_VERSION : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        ALLOW_X8_GEN2   : string  := "FALSE";
        BAR0            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR1            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR2            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        BAR3            : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        BAR4            : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        BAR5            : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CAPABILITIES_PTR: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CARDBUS_CIS_POINTER: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLASS_CODE      : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CMD_INTX_IMPLEMENTED: string  := "TRUE";
        CPL_TIMEOUT_DISABLE_SUPPORTED: string  := "FALSE";
        CPL_TIMEOUT_RANGES_SUPPORTED: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        CRM_MODULE_RSTS : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DEVICE_ID       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE: string  := "TRUE";
        DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE: string  := "TRUE";
        DEV_CAP_ENDPOINT_L0S_LATENCY: integer := 0;
        DEV_CAP_ENDPOINT_L1_LATENCY: integer := 0;
        DEV_CAP_EXT_TAG_SUPPORTED: string  := "TRUE";
        DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE: string  := "FALSE";
        DEV_CAP_MAX_PAYLOAD_SUPPORTED: integer := 2;
        DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT: integer := 0;
        DEV_CAP_ROLE_BASED_ERROR: string  := "TRUE";
        DEV_CAP_RSVD_14_12: integer := 0;
        DEV_CAP_RSVD_17_16: integer := 0;
        DEV_CAP_RSVD_31_29: integer := 0;
        DEV_CONTROL_AUX_POWER_SUPPORTED: string  := "FALSE";
        DISABLE_ASPM_L1_TIMER: string  := "FALSE";
        DISABLE_BAR_FILTERING: string  := "FALSE";
        DISABLE_ID_CHECK: string  := "FALSE";
        DISABLE_LANE_REVERSAL: string  := "FALSE";
        DISABLE_RX_TC_FILTER: string  := "FALSE";
        DISABLE_SCRAMBLING: string  := "FALSE";
        DNSTREAM_LINK_NUM: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DSN_BASE_PTR    : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DSN_CAP_ID      : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        DSN_CAP_NEXTPTR : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        DSN_CAP_ON      : string  := "TRUE";
        DSN_CAP_VERSION : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        ENABLE_MSG_ROUTE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ENABLE_RX_TD_ECRC_TRIM: string  := "FALSE";
        ENTER_RVRY_EI_L0: string  := "TRUE";
        EXIT_LOOPBACK_ON_EI: string  := "TRUE";
        EXPANSION_ROM   : vl_logic_vector(31 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        EXT_CFG_CAP_PTR : vl_logic_vector(5 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        EXT_CFG_XP_CAP_PTR: vl_logic_vector(9 downto 0) := (Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        HEADER_TYPE     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        INFER_EI        : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        INTERRUPT_PIN   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        IS_SWITCH       : string  := "FALSE";
        LAST_CONFIG_DWORD: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        LINK_CAP_ASPM_SUPPORT: integer := 1;
        LINK_CAP_CLOCK_POWER_MANAGEMENT: string  := "FALSE";
        LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP: string  := "FALSE";
        LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1: integer := 7;
        LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2: integer := 7;
        LINK_CAP_L0S_EXIT_LATENCY_GEN1: integer := 7;
        LINK_CAP_L0S_EXIT_LATENCY_GEN2: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_GEN1: integer := 7;
        LINK_CAP_L1_EXIT_LATENCY_GEN2: integer := 7;
        LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP: string  := "FALSE";
        LINK_CAP_MAX_LINK_SPEED: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        LINK_CAP_MAX_LINK_WIDTH: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        LINK_CAP_RSVD_23_22: integer := 0;
        LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE: string  := "FALSE";
        LINK_CONTROL_RCB: integer := 0;
        LINK_CTRL2_DEEMPHASIS: string  := "FALSE";
        LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE: string  := "FALSE";
        LINK_CTRL2_TARGET_LINK_SPEED: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        LINK_STATUS_SLOT_CLOCK_CONFIG: string  := "TRUE";
        LL_ACK_TIMEOUT  : vl_logic_vector(14 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_ACK_TIMEOUT_EN: string  := "FALSE";
        LL_ACK_TIMEOUT_FUNC: integer := 0;
        LL_REPLAY_TIMEOUT: vl_logic_vector(14 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_REPLAY_TIMEOUT_EN: string  := "FALSE";
        LL_REPLAY_TIMEOUT_FUNC: integer := 0;
        LTSSM_MAX_LINK_WIDTH: vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        MSIX_BASE_PTR   : vl_logic_vector(7 downto 0) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        MSIX_CAP_ID     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1);
        MSIX_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MSIX_CAP_ON     : string  := "FALSE";
        MSIX_CAP_PBA_BIR: integer := 0;
        MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        MSIX_CAP_TABLE_BIR: integer := 0;
        MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        MSI_BASE_PTR    : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        MSI_CAP_64_BIT_ADDR_CAPABLE: string  := "TRUE";
        MSI_CAP_ID      : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        MSI_CAP_MULTIMSGCAP: integer := 0;
        MSI_CAP_MULTIMSG_EXTENSION: integer := 0;
        MSI_CAP_NEXTPTR : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        MSI_CAP_ON      : string  := "FALSE";
        MSI_CAP_PER_VECTOR_MASKING_CAPABLE: string  := "TRUE";
        N_FTS_COMCLK_GEN1: integer := 255;
        N_FTS_COMCLK_GEN2: integer := 255;
        N_FTS_GEN1      : integer := 255;
        N_FTS_GEN2      : integer := 255;
        PCIE_BASE_PTR   : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        PCIE_CAP_CAPABILITY_ID: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        PCIE_CAP_CAPABILITY_VERSION: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        PCIE_CAP_DEVICE_PORT_TYPE: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        PCIE_CAP_INT_MSG_NUM: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PCIE_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PCIE_CAP_ON     : string  := "TRUE";
        PCIE_CAP_RSVD_15_14: integer := 0;
        PCIE_CAP_SLOT_IMPLEMENTED: string  := "FALSE";
        PCIE_REVISION   : integer := 2;
        PGL0_LANE       : integer := 0;
        PGL1_LANE       : integer := 1;
        PGL2_LANE       : integer := 2;
        PGL3_LANE       : integer := 3;
        PGL4_LANE       : integer := 4;
        PGL5_LANE       : integer := 5;
        PGL6_LANE       : integer := 6;
        PGL7_LANE       : integer := 7;
        PL_AUTO_CONFIG  : integer := 0;
        PL_FAST_TRAIN   : string  := "FALSE";
        PM_BASE_PTR     : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PM_CAP_AUXCURRENT: integer := 0;
        PM_CAP_D1SUPPORT: string  := "TRUE";
        PM_CAP_D2SUPPORT: string  := "TRUE";
        PM_CAP_DSI      : string  := "FALSE";
        PM_CAP_ID       : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_CAP_NEXTPTR  : vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        PM_CAP_ON       : string  := "TRUE";
        PM_CAP_PMESUPPORT: vl_logic_vector(4 downto 0) := (Hi0, Hi1, Hi1, Hi1, Hi1);
        PM_CAP_PME_CLOCK: string  := "FALSE";
        PM_CAP_RSVD_04  : integer := 0;
        PM_CAP_VERSION  : integer := 3;
        PM_CSR_B2B3     : string  := "FALSE";
        PM_CSR_BPCCEN   : string  := "FALSE";
        PM_CSR_NOSOFTRST: string  := "TRUE";
        PM_DATA0        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA1        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA2        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA3        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA4        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA5        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA6        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA7        : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PM_DATA_SCALE0  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE1  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE2  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE3  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE4  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE5  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE6  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PM_DATA_SCALE7  : vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        RECRC_CHK       : integer := 0;
        RECRC_CHK_TRIM  : string  := "FALSE";
        REVISION_ID     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ROOT_CAP_CRS_SW_VISIBILITY: string  := "FALSE";
        SELECT_DLL_IF   : string  := "FALSE";
        SIM_VERSION     : string  := "1.0";
        SLOT_CAP_ATT_BUTTON_PRESENT: string  := "FALSE";
        SLOT_CAP_ATT_INDICATOR_PRESENT: string  := "FALSE";
        SLOT_CAP_ELEC_INTERLOCK_PRESENT: string  := "FALSE";
        SLOT_CAP_HOTPLUG_CAPABLE: string  := "FALSE";
        SLOT_CAP_HOTPLUG_SURPRISE: string  := "FALSE";
        SLOT_CAP_MRL_SENSOR_PRESENT: string  := "FALSE";
        SLOT_CAP_NO_CMD_COMPLETED_SUPPORT: string  := "FALSE";
        SLOT_CAP_PHYSICAL_SLOT_NUM: vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SLOT_CAP_POWER_CONTROLLER_PRESENT: string  := "FALSE";
        SLOT_CAP_POWER_INDICATOR_PRESENT: string  := "FALSE";
        SLOT_CAP_SLOT_POWER_LIMIT_SCALE: integer := 0;
        SLOT_CAP_SLOT_POWER_LIMIT_VALUE: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BIT0      : integer := 0;
        SPARE_BIT1      : integer := 0;
        SPARE_BIT2      : integer := 0;
        SPARE_BIT3      : integer := 0;
        SPARE_BIT4      : integer := 0;
        SPARE_BIT5      : integer := 0;
        SPARE_BIT6      : integer := 0;
        SPARE_BIT7      : integer := 0;
        SPARE_BIT8      : integer := 0;
        SPARE_BYTE0     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BYTE1     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BYTE2     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BYTE3     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD0     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD1     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD2     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD3     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SUBSYSTEM_ID    : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1);
        SUBSYSTEM_VENDOR_ID: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        TL_RBYPASS      : string  := "FALSE";
        TL_RX_RAM_RADDR_LATENCY: integer := 0;
        TL_RX_RAM_RDATA_LATENCY: integer := 2;
        TL_RX_RAM_WRITE_LATENCY: integer := 0;
        TL_TFC_DISABLE  : string  := "FALSE";
        TL_TX_CHECKS_DISABLE: string  := "FALSE";
        TL_TX_RAM_RADDR_LATENCY: integer := 0;
        TL_TX_RAM_RDATA_LATENCY: integer := 2;
        TL_TX_RAM_WRITE_LATENCY: integer := 0;
        UPCONFIG_CAPABLE: string  := "TRUE";
        UPSTREAM_FACING : string  := "TRUE";
        UR_INV_REQ      : string  := "TRUE";
        USER_CLK_FREQ   : integer := 3;
        VC0_CPL_INFINITE: string  := "TRUE";
        VC0_RX_RAM_LIMIT: vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        VC0_TOTAL_CREDITS_CD: integer := 127;
        VC0_TOTAL_CREDITS_CH: integer := 31;
        VC0_TOTAL_CREDITS_NPH: integer := 12;
        VC0_TOTAL_CREDITS_PD: integer := 288;
        VC0_TOTAL_CREDITS_PH: integer := 32;
        VC0_TX_LASTPACKET: integer := 31;
        VC_BASE_PTR     : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        VC_CAP_ID       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        VC_CAP_NEXTPTR  : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VC_CAP_ON       : string  := "FALSE";
        VC_CAP_REJECT_SNOOP_TRANSACTIONS: string  := "FALSE";
        VC_CAP_VERSION  : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VENDOR_ID       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0);
        VSEC_BASE_PTR   : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        VSEC_CAP_HDR_ID : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0);
        VSEC_CAP_HDR_LENGTH: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        VSEC_CAP_HDR_REVISION: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VSEC_CAP_ID     : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1);
        VSEC_CAP_IS_LINK_VISIBLE: string  := "TRUE";
        VSEC_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VSEC_CAP_ON     : string  := "FALSE";
        VSEC_CAP_VERSION: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1)
    );
    port(
        CFGAERECRCCHECKEN: out    vl_logic;
        CFGAERECRCGENEN : out    vl_logic;
        CFGCOMMANDBUSMASTERENABLE: out    vl_logic;
        CFGCOMMANDINTERRUPTDISABLE: out    vl_logic;
        CFGCOMMANDIOENABLE: out    vl_logic;
        CFGCOMMANDMEMENABLE: out    vl_logic;
        CFGCOMMANDSERREN: out    vl_logic;
        CFGDEVCONTROL2CPLTIMEOUTDIS: out    vl_logic;
        CFGDEVCONTROL2CPLTIMEOUTVAL: out    vl_logic_vector(3 downto 0);
        CFGDEVCONTROLAUXPOWEREN: out    vl_logic;
        CFGDEVCONTROLCORRERRREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLENABLERO: out    vl_logic;
        CFGDEVCONTROLEXTTAGEN: out    vl_logic;
        CFGDEVCONTROLFATALERRREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLMAXPAYLOAD: out    vl_logic_vector(2 downto 0);
        CFGDEVCONTROLMAXREADREQ: out    vl_logic_vector(2 downto 0);
        CFGDEVCONTROLNONFATALREPORTINGEN: out    vl_logic;
        CFGDEVCONTROLNOSNOOPEN: out    vl_logic;
        CFGDEVCONTROLPHANTOMEN: out    vl_logic;
        CFGDEVCONTROLURERRREPORTINGEN: out    vl_logic;
        CFGDEVSTATUSCORRERRDETECTED: out    vl_logic;
        CFGDEVSTATUSFATALERRDETECTED: out    vl_logic;
        CFGDEVSTATUSNONFATALERRDETECTED: out    vl_logic;
        CFGDEVSTATUSURDETECTED: out    vl_logic;
        CFGDO           : out    vl_logic_vector(31 downto 0);
        CFGERRAERHEADERLOGSETN: out    vl_logic;
        CFGERRCPLRDYN   : out    vl_logic;
        CFGINTERRUPTDO  : out    vl_logic_vector(7 downto 0);
        CFGINTERRUPTMMENABLE: out    vl_logic_vector(2 downto 0);
        CFGINTERRUPTMSIENABLE: out    vl_logic;
        CFGINTERRUPTMSIXENABLE: out    vl_logic;
        CFGINTERRUPTMSIXFM: out    vl_logic;
        CFGINTERRUPTRDYN: out    vl_logic;
        CFGLINKCONTROLASPMCONTROL: out    vl_logic_vector(1 downto 0);
        CFGLINKCONTROLAUTOBANDWIDTHINTEN: out    vl_logic;
        CFGLINKCONTROLBANDWIDTHINTEN: out    vl_logic;
        CFGLINKCONTROLCLOCKPMEN: out    vl_logic;
        CFGLINKCONTROLCOMMONCLOCK: out    vl_logic;
        CFGLINKCONTROLEXTENDEDSYNC: out    vl_logic;
        CFGLINKCONTROLHWAUTOWIDTHDIS: out    vl_logic;
        CFGLINKCONTROLLINKDISABLE: out    vl_logic;
        CFGLINKCONTROLRCB: out    vl_logic;
        CFGLINKCONTROLRETRAINLINK: out    vl_logic;
        CFGLINKSTATUSAUTOBANDWIDTHSTATUS: out    vl_logic;
        CFGLINKSTATUSBANDWITHSTATUS: out    vl_logic;
        CFGLINKSTATUSCURRENTSPEED: out    vl_logic_vector(1 downto 0);
        CFGLINKSTATUSDLLACTIVE: out    vl_logic;
        CFGLINKSTATUSLINKTRAINING: out    vl_logic;
        CFGLINKSTATUSNEGOTIATEDWIDTH: out    vl_logic_vector(3 downto 0);
        CFGMSGDATA      : out    vl_logic_vector(15 downto 0);
        CFGMSGRECEIVED  : out    vl_logic;
        CFGMSGRECEIVEDASSERTINTA: out    vl_logic;
        CFGMSGRECEIVEDASSERTINTB: out    vl_logic;
        CFGMSGRECEIVEDASSERTINTC: out    vl_logic;
        CFGMSGRECEIVEDASSERTINTD: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTA: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTB: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTC: out    vl_logic;
        CFGMSGRECEIVEDDEASSERTINTD: out    vl_logic;
        CFGMSGRECEIVEDERRCOR: out    vl_logic;
        CFGMSGRECEIVEDERRFATAL: out    vl_logic;
        CFGMSGRECEIVEDERRNONFATAL: out    vl_logic;
        CFGMSGRECEIVEDPMASNAK: out    vl_logic;
        CFGMSGRECEIVEDPMETO: out    vl_logic;
        CFGMSGRECEIVEDPMETOACK: out    vl_logic;
        CFGMSGRECEIVEDPMPME: out    vl_logic;
        CFGMSGRECEIVEDSETSLOTPOWERLIMIT: out    vl_logic;
        CFGMSGRECEIVEDUNLOCK: out    vl_logic;
        CFGPCIELINKSTATE: out    vl_logic_vector(2 downto 0);
        CFGPMCSRPMEEN   : out    vl_logic;
        CFGPMCSRPMESTATUS: out    vl_logic;
        CFGPMCSRPOWERSTATE: out    vl_logic_vector(1 downto 0);
        CFGPMRCVASREQL1N: out    vl_logic;
        CFGPMRCVENTERL1N: out    vl_logic;
        CFGPMRCVENTERL23N: out    vl_logic;
        CFGPMRCVREQACKN : out    vl_logic;
        CFGRDWRDONEN    : out    vl_logic;
        CFGSLOTCONTROLELECTROMECHILCTLPULSE: out    vl_logic;
        CFGTRANSACTION  : out    vl_logic;
        CFGTRANSACTIONADDR: out    vl_logic_vector(6 downto 0);
        CFGTRANSACTIONTYPE: out    vl_logic;
        CFGVCTCVCMAP    : out    vl_logic_vector(6 downto 0);
        DBGSCLRA        : out    vl_logic;
        DBGSCLRB        : out    vl_logic;
        DBGSCLRC        : out    vl_logic;
        DBGSCLRD        : out    vl_logic;
        DBGSCLRE        : out    vl_logic;
        DBGSCLRF        : out    vl_logic;
        DBGSCLRG        : out    vl_logic;
        DBGSCLRH        : out    vl_logic;
        DBGSCLRI        : out    vl_logic;
        DBGSCLRJ        : out    vl_logic;
        DBGSCLRK        : out    vl_logic;
        DBGVECA         : out    vl_logic_vector(63 downto 0);
        DBGVECB         : out    vl_logic_vector(63 downto 0);
        DBGVECC         : out    vl_logic_vector(11 downto 0);
        DRPDO           : out    vl_logic_vector(15 downto 0);
        DRPDRDY         : out    vl_logic;
        LL2BADDLLPERRN  : out    vl_logic;
        LL2BADTLPERRN   : out    vl_logic;
        LL2PROTOCOLERRN : out    vl_logic;
        LL2REPLAYROERRN : out    vl_logic;
        LL2REPLAYTOERRN : out    vl_logic;
        LL2SUSPENDOKN   : out    vl_logic;
        LL2TFCINIT1SEQN : out    vl_logic;
        LL2TFCINIT2SEQN : out    vl_logic;
        LNKCLKEN        : out    vl_logic;
        MIMRXRADDR      : out    vl_logic_vector(12 downto 0);
        MIMRXRCE        : out    vl_logic;
        MIMRXREN        : out    vl_logic;
        MIMRXWADDR      : out    vl_logic_vector(12 downto 0);
        MIMRXWDATA      : out    vl_logic_vector(67 downto 0);
        MIMRXWEN        : out    vl_logic;
        MIMTXRADDR      : out    vl_logic_vector(12 downto 0);
        MIMTXRCE        : out    vl_logic;
        MIMTXREN        : out    vl_logic;
        MIMTXWADDR      : out    vl_logic_vector(12 downto 0);
        MIMTXWDATA      : out    vl_logic_vector(68 downto 0);
        MIMTXWEN        : out    vl_logic;
        PIPERX0POLARITY : out    vl_logic;
        PIPERX1POLARITY : out    vl_logic;
        PIPERX2POLARITY : out    vl_logic;
        PIPERX3POLARITY : out    vl_logic;
        PIPERX4POLARITY : out    vl_logic;
        PIPERX5POLARITY : out    vl_logic;
        PIPERX6POLARITY : out    vl_logic;
        PIPERX7POLARITY : out    vl_logic;
        PIPETX0CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX0COMPLIANCE: out    vl_logic;
        PIPETX0DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX0ELECIDLE : out    vl_logic;
        PIPETX0POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX1CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX1COMPLIANCE: out    vl_logic;
        PIPETX1DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX1ELECIDLE : out    vl_logic;
        PIPETX1POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX2CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX2COMPLIANCE: out    vl_logic;
        PIPETX2DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX2ELECIDLE : out    vl_logic;
        PIPETX2POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX3CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX3COMPLIANCE: out    vl_logic;
        PIPETX3DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX3ELECIDLE : out    vl_logic;
        PIPETX3POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX4CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX4COMPLIANCE: out    vl_logic;
        PIPETX4DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX4ELECIDLE : out    vl_logic;
        PIPETX4POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX5CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX5COMPLIANCE: out    vl_logic;
        PIPETX5DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX5ELECIDLE : out    vl_logic;
        PIPETX5POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX6CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX6COMPLIANCE: out    vl_logic;
        PIPETX6DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX6ELECIDLE : out    vl_logic;
        PIPETX6POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX7CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX7COMPLIANCE: out    vl_logic;
        PIPETX7DATA     : out    vl_logic_vector(15 downto 0);
        PIPETX7ELECIDLE : out    vl_logic;
        PIPETX7POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETXDEEMPH    : out    vl_logic;
        PIPETXMARGIN    : out    vl_logic_vector(2 downto 0);
        PIPETXRATE      : out    vl_logic;
        PIPETXRCVRDET   : out    vl_logic;
        PIPETXRESET     : out    vl_logic;
        PL2LINKUPN      : out    vl_logic;
        PL2RECEIVERERRN : out    vl_logic;
        PL2RECOVERYN    : out    vl_logic;
        PL2RXELECIDLE   : out    vl_logic;
        PL2SUSPENDOK    : out    vl_logic;
        PLDBGVEC        : out    vl_logic_vector(11 downto 0);
        PLINITIALLINKWIDTH: out    vl_logic_vector(2 downto 0);
        PLLANEREVERSALMODE: out    vl_logic_vector(1 downto 0);
        PLLINKGEN2CAP   : out    vl_logic;
        PLLINKPARTNERGEN2SUPPORTED: out    vl_logic;
        PLLINKUPCFGCAP  : out    vl_logic;
        PLLTSSMSTATE    : out    vl_logic_vector(5 downto 0);
        PLPHYLNKUPN     : out    vl_logic;
        PLRECEIVEDHOTRST: out    vl_logic;
        PLRXPMSTATE     : out    vl_logic_vector(1 downto 0);
        PLSELLNKRATE    : out    vl_logic;
        PLSELLNKWIDTH   : out    vl_logic_vector(1 downto 0);
        PLTXPMSTATE     : out    vl_logic_vector(2 downto 0);
        RECEIVEDFUNCLVLRSTN: out    vl_logic;
        TL2ASPMSUSPENDCREDITCHECKOKN: out    vl_logic;
        TL2ASPMSUSPENDREQN: out    vl_logic;
        TL2PPMSUSPENDOKN: out    vl_logic;
        TRNFCCPLD       : out    vl_logic_vector(11 downto 0);
        TRNFCCPLH       : out    vl_logic_vector(7 downto 0);
        TRNFCNPD        : out    vl_logic_vector(11 downto 0);
        TRNFCNPH        : out    vl_logic_vector(7 downto 0);
        TRNFCPD         : out    vl_logic_vector(11 downto 0);
        TRNFCPH         : out    vl_logic_vector(7 downto 0);
        TRNLNKUPN       : out    vl_logic;
        TRNRBARHITN     : out    vl_logic_vector(6 downto 0);
        TRNRD           : out    vl_logic_vector(63 downto 0);
        TRNRDLLPDATA    : out    vl_logic_vector(31 downto 0);
        TRNRDLLPSRCRDYN : out    vl_logic;
        TRNRECRCERRN    : out    vl_logic;
        TRNREOFN        : out    vl_logic;
        TRNRERRFWDN     : out    vl_logic;
        TRNRREMN        : out    vl_logic;
        TRNRSOFN        : out    vl_logic;
        TRNRSRCDSCN     : out    vl_logic;
        TRNRSRCRDYN     : out    vl_logic;
        TRNTBUFAV       : out    vl_logic_vector(5 downto 0);
        TRNTCFGREQN     : out    vl_logic;
        TRNTDLLPDSTRDYN : out    vl_logic;
        TRNTDSTRDYN     : out    vl_logic;
        TRNTERRDROPN    : out    vl_logic;
        USERRSTN        : out    vl_logic;
        CFGBYTEENN      : in     vl_logic_vector(3 downto 0);
        CFGDI           : in     vl_logic_vector(31 downto 0);
        CFGDSBUSNUMBER  : in     vl_logic_vector(7 downto 0);
        CFGDSDEVICENUMBER: in     vl_logic_vector(4 downto 0);
        CFGDSFUNCTIONNUMBER: in     vl_logic_vector(2 downto 0);
        CFGDSN          : in     vl_logic_vector(63 downto 0);
        CFGDWADDR       : in     vl_logic_vector(9 downto 0);
        CFGERRACSN      : in     vl_logic;
        CFGERRAERHEADERLOG: in     vl_logic_vector(127 downto 0);
        CFGERRCORN      : in     vl_logic;
        CFGERRCPLABORTN : in     vl_logic;
        CFGERRCPLTIMEOUTN: in     vl_logic;
        CFGERRCPLUNEXPECTN: in     vl_logic;
        CFGERRECRCN     : in     vl_logic;
        CFGERRLOCKEDN   : in     vl_logic;
        CFGERRPOSTEDN   : in     vl_logic;
        CFGERRTLPCPLHEADER: in     vl_logic_vector(47 downto 0);
        CFGERRURN       : in     vl_logic;
        CFGINTERRUPTASSERTN: in     vl_logic;
        CFGINTERRUPTDI  : in     vl_logic_vector(7 downto 0);
        CFGINTERRUPTN   : in     vl_logic;
        CFGPMDIRECTASPML1N: in     vl_logic;
        CFGPMSENDPMACKN : in     vl_logic;
        CFGPMSENDPMETON : in     vl_logic;
        CFGPMSENDPMNAKN : in     vl_logic;
        CFGPMTURNOFFOKN : in     vl_logic;
        CFGPMWAKEN      : in     vl_logic;
        CFGPORTNUMBER   : in     vl_logic_vector(7 downto 0);
        CFGRDENN        : in     vl_logic;
        CFGTRNPENDINGN  : in     vl_logic;
        CFGWRENN        : in     vl_logic;
        CFGWRREADONLYN  : in     vl_logic;
        CFGWRRW1CASRWN  : in     vl_logic;
        CMRSTN          : in     vl_logic;
        CMSTICKYRSTN    : in     vl_logic;
        DBGMODE         : in     vl_logic_vector(1 downto 0);
        DBGSUBMODE      : in     vl_logic;
        DLRSTN          : in     vl_logic;
        DRPCLK          : in     vl_logic;
        DRPDADDR        : in     vl_logic_vector(8 downto 0);
        DRPDEN          : in     vl_logic;
        DRPDI           : in     vl_logic_vector(15 downto 0);
        DRPDWE          : in     vl_logic;
        FUNCLVLRSTN     : in     vl_logic;
        LL2SENDASREQL1N : in     vl_logic;
        LL2SENDENTERL1N : in     vl_logic;
        LL2SENDENTERL23N: in     vl_logic;
        LL2SUSPENDNOWN  : in     vl_logic;
        LL2TLPRCVN      : in     vl_logic;
        MIMRXRDATA      : in     vl_logic_vector(67 downto 0);
        MIMTXRDATA      : in     vl_logic_vector(68 downto 0);
        PIPECLK         : in     vl_logic;
        PIPERX0CHANISALIGNED: in     vl_logic;
        PIPERX0CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX0DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX0ELECIDLE : in     vl_logic;
        PIPERX0PHYSTATUS: in     vl_logic;
        PIPERX0STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX0VALID    : in     vl_logic;
        PIPERX1CHANISALIGNED: in     vl_logic;
        PIPERX1CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX1DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX1ELECIDLE : in     vl_logic;
        PIPERX1PHYSTATUS: in     vl_logic;
        PIPERX1STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX1VALID    : in     vl_logic;
        PIPERX2CHANISALIGNED: in     vl_logic;
        PIPERX2CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX2DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX2ELECIDLE : in     vl_logic;
        PIPERX2PHYSTATUS: in     vl_logic;
        PIPERX2STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX2VALID    : in     vl_logic;
        PIPERX3CHANISALIGNED: in     vl_logic;
        PIPERX3CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX3DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX3ELECIDLE : in     vl_logic;
        PIPERX3PHYSTATUS: in     vl_logic;
        PIPERX3STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX3VALID    : in     vl_logic;
        PIPERX4CHANISALIGNED: in     vl_logic;
        PIPERX4CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX4DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX4ELECIDLE : in     vl_logic;
        PIPERX4PHYSTATUS: in     vl_logic;
        PIPERX4STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX4VALID    : in     vl_logic;
        PIPERX5CHANISALIGNED: in     vl_logic;
        PIPERX5CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX5DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX5ELECIDLE : in     vl_logic;
        PIPERX5PHYSTATUS: in     vl_logic;
        PIPERX5STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX5VALID    : in     vl_logic;
        PIPERX6CHANISALIGNED: in     vl_logic;
        PIPERX6CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX6DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX6ELECIDLE : in     vl_logic;
        PIPERX6PHYSTATUS: in     vl_logic;
        PIPERX6STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX6VALID    : in     vl_logic;
        PIPERX7CHANISALIGNED: in     vl_logic;
        PIPERX7CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX7DATA     : in     vl_logic_vector(15 downto 0);
        PIPERX7ELECIDLE : in     vl_logic;
        PIPERX7PHYSTATUS: in     vl_logic;
        PIPERX7STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX7VALID    : in     vl_logic;
        PL2DIRECTEDLSTATE: in     vl_logic_vector(4 downto 0);
        PLDBGMODE       : in     vl_logic_vector(2 downto 0);
        PLDIRECTEDLINKAUTON: in     vl_logic;
        PLDIRECTEDLINKCHANGE: in     vl_logic_vector(1 downto 0);
        PLDIRECTEDLINKSPEED: in     vl_logic;
        PLDIRECTEDLINKWIDTH: in     vl_logic_vector(1 downto 0);
        PLDOWNSTREAMDEEMPHSOURCE: in     vl_logic;
        PLRSTN          : in     vl_logic;
        PLTRANSMITHOTRST: in     vl_logic;
        PLUPSTREAMPREFERDEEMPH: in     vl_logic;
        SYSRSTN         : in     vl_logic;
        TL2ASPMSUSPENDCREDITCHECKN: in     vl_logic;
        TL2PPMSUSPENDREQN: in     vl_logic;
        TLRSTN          : in     vl_logic;
        TRNFCSEL        : in     vl_logic_vector(2 downto 0);
        TRNRDSTRDYN     : in     vl_logic;
        TRNRNPOKN       : in     vl_logic;
        TRNTCFGGNTN     : in     vl_logic;
        TRNTD           : in     vl_logic_vector(63 downto 0);
        TRNTDLLPDATA    : in     vl_logic_vector(31 downto 0);
        TRNTDLLPSRCRDYN : in     vl_logic;
        TRNTECRCGENN    : in     vl_logic;
        TRNTEOFN        : in     vl_logic;
        TRNTERRFWDN     : in     vl_logic;
        TRNTREMN        : in     vl_logic;
        TRNTSOFN        : in     vl_logic;
        TRNTSRCDSCN     : in     vl_logic;
        TRNTSRCRDYN     : in     vl_logic;
        TRNTSTRN        : in     vl_logic;
        USERCLK         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of AER_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of AER_CAP_ECRC_CHECK_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_ECRC_GEN_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of AER_CAP_INT_MSG_NUM_MSI : constant is 2;
    attribute mti_svvh_generic_type of AER_CAP_INT_MSG_NUM_MSIX : constant is 2;
    attribute mti_svvh_generic_type of AER_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of AER_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_PERMIT_ROOTERR_UPDATE : constant is 1;
    attribute mti_svvh_generic_type of AER_CAP_VERSION : constant is 2;
    attribute mti_svvh_generic_type of ALLOW_X8_GEN2 : constant is 1;
    attribute mti_svvh_generic_type of BAR0 : constant is 2;
    attribute mti_svvh_generic_type of BAR1 : constant is 2;
    attribute mti_svvh_generic_type of BAR2 : constant is 2;
    attribute mti_svvh_generic_type of BAR3 : constant is 2;
    attribute mti_svvh_generic_type of BAR4 : constant is 2;
    attribute mti_svvh_generic_type of BAR5 : constant is 2;
    attribute mti_svvh_generic_type of CAPABILITIES_PTR : constant is 2;
    attribute mti_svvh_generic_type of CARDBUS_CIS_POINTER : constant is 2;
    attribute mti_svvh_generic_type of CLASS_CODE : constant is 2;
    attribute mti_svvh_generic_type of CMD_INTX_IMPLEMENTED : constant is 1;
    attribute mti_svvh_generic_type of CPL_TIMEOUT_DISABLE_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of CPL_TIMEOUT_RANGES_SUPPORTED : constant is 2;
    attribute mti_svvh_generic_type of CRM_MODULE_RSTS : constant is 2;
    attribute mti_svvh_generic_type of DEVICE_ID : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_ENABLE_SLOT_PWR_LIMIT_SCALE : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_ENABLE_SLOT_PWR_LIMIT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_ENDPOINT_L0S_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_ENDPOINT_L1_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_EXT_TAG_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_MAX_PAYLOAD_SUPPORTED : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_PHANTOM_FUNCTIONS_SUPPORT : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_ROLE_BASED_ERROR : constant is 1;
    attribute mti_svvh_generic_type of DEV_CAP_RSVD_14_12 : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_RSVD_17_16 : constant is 2;
    attribute mti_svvh_generic_type of DEV_CAP_RSVD_31_29 : constant is 2;
    attribute mti_svvh_generic_type of DEV_CONTROL_AUX_POWER_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_ASPM_L1_TIMER : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_BAR_FILTERING : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_ID_CHECK : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_LANE_REVERSAL : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_RX_TC_FILTER : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_SCRAMBLING : constant is 1;
    attribute mti_svvh_generic_type of DNSTREAM_LINK_NUM : constant is 2;
    attribute mti_svvh_generic_type of DSN_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of DSN_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of DSN_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of DSN_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of DSN_CAP_VERSION : constant is 2;
    attribute mti_svvh_generic_type of ENABLE_MSG_ROUTE : constant is 2;
    attribute mti_svvh_generic_type of ENABLE_RX_TD_ECRC_TRIM : constant is 1;
    attribute mti_svvh_generic_type of ENTER_RVRY_EI_L0 : constant is 1;
    attribute mti_svvh_generic_type of EXIT_LOOPBACK_ON_EI : constant is 1;
    attribute mti_svvh_generic_type of EXPANSION_ROM : constant is 2;
    attribute mti_svvh_generic_type of EXT_CFG_CAP_PTR : constant is 2;
    attribute mti_svvh_generic_type of EXT_CFG_XP_CAP_PTR : constant is 2;
    attribute mti_svvh_generic_type of HEADER_TYPE : constant is 2;
    attribute mti_svvh_generic_type of INFER_EI : constant is 2;
    attribute mti_svvh_generic_type of INTERRUPT_PIN : constant is 2;
    attribute mti_svvh_generic_type of IS_SWITCH : constant is 1;
    attribute mti_svvh_generic_type of LAST_CONFIG_DWORD : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_ASPM_SUPPORT : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_CLOCK_POWER_MANAGEMENT : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_DLL_LINK_ACTIVE_REPORTING_CAP : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L0S_EXIT_LATENCY_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_L1_EXIT_LATENCY_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_LINK_BANDWIDTH_NOTIFICATION_CAP : constant is 1;
    attribute mti_svvh_generic_type of LINK_CAP_MAX_LINK_SPEED : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_MAX_LINK_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_RSVD_23_22 : constant is 2;
    attribute mti_svvh_generic_type of LINK_CAP_SURPRISE_DOWN_ERROR_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of LINK_CONTROL_RCB : constant is 2;
    attribute mti_svvh_generic_type of LINK_CTRL2_DEEMPHASIS : constant is 1;
    attribute mti_svvh_generic_type of LINK_CTRL2_HW_AUTONOMOUS_SPEED_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of LINK_CTRL2_TARGET_LINK_SPEED : constant is 2;
    attribute mti_svvh_generic_type of LINK_STATUS_SLOT_CLOCK_CONFIG : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT : constant is 2;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT : constant is 2;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of LTSSM_MAX_LINK_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of MSIX_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of MSI_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_64_BIT_ADDR_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_MULTIMSG_EXTENSION : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of MSI_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of MSI_CAP_PER_VECTOR_MASKING_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of N_FTS_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of N_FTS_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of N_FTS_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of N_FTS_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PCIE_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_CAPABILITY_ID : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_CAPABILITY_VERSION : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_DEVICE_PORT_TYPE : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_INT_MSG_NUM : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of PCIE_CAP_RSVD_15_14 : constant is 2;
    attribute mti_svvh_generic_type of PCIE_CAP_SLOT_IMPLEMENTED : constant is 1;
    attribute mti_svvh_generic_type of PCIE_REVISION : constant is 2;
    attribute mti_svvh_generic_type of PGL0_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL1_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL2_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL3_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL4_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL5_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL6_LANE : constant is 2;
    attribute mti_svvh_generic_type of PGL7_LANE : constant is 2;
    attribute mti_svvh_generic_type of PL_AUTO_CONFIG : constant is 2;
    attribute mti_svvh_generic_type of PL_FAST_TRAIN : constant is 1;
    attribute mti_svvh_generic_type of PM_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_AUXCURRENT : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_D1SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_D2SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_DSI : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_PMESUPPORT : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_PME_CLOCK : constant is 1;
    attribute mti_svvh_generic_type of PM_CAP_RSVD_04 : constant is 2;
    attribute mti_svvh_generic_type of PM_CAP_VERSION : constant is 2;
    attribute mti_svvh_generic_type of PM_CSR_B2B3 : constant is 1;
    attribute mti_svvh_generic_type of PM_CSR_BPCCEN : constant is 1;
    attribute mti_svvh_generic_type of PM_CSR_NOSOFTRST : constant is 1;
    attribute mti_svvh_generic_type of PM_DATA0 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA1 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA2 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA3 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA4 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA5 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA6 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA7 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE0 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE1 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE2 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE3 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE4 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE5 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE6 : constant is 2;
    attribute mti_svvh_generic_type of PM_DATA_SCALE7 : constant is 2;
    attribute mti_svvh_generic_type of RECRC_CHK : constant is 2;
    attribute mti_svvh_generic_type of RECRC_CHK_TRIM : constant is 1;
    attribute mti_svvh_generic_type of REVISION_ID : constant is 2;
    attribute mti_svvh_generic_type of ROOT_CAP_CRS_SW_VISIBILITY : constant is 1;
    attribute mti_svvh_generic_type of SELECT_DLL_IF : constant is 1;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_ATT_BUTTON_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_ATT_INDICATOR_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_ELEC_INTERLOCK_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_HOTPLUG_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_HOTPLUG_SURPRISE : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_MRL_SENSOR_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_NO_CMD_COMPLETED_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_PHYSICAL_SLOT_NUM : constant is 2;
    attribute mti_svvh_generic_type of SLOT_CAP_POWER_CONTROLLER_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_POWER_INDICATOR_PRESENT : constant is 1;
    attribute mti_svvh_generic_type of SLOT_CAP_SLOT_POWER_LIMIT_SCALE : constant is 2;
    attribute mti_svvh_generic_type of SLOT_CAP_SLOT_POWER_LIMIT_VALUE : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT3 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT4 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT5 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT6 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT7 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT8 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE3 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD3 : constant is 2;
    attribute mti_svvh_generic_type of SUBSYSTEM_ID : constant is 2;
    attribute mti_svvh_generic_type of SUBSYSTEM_VENDOR_ID : constant is 2;
    attribute mti_svvh_generic_type of TL_RBYPASS : constant is 1;
    attribute mti_svvh_generic_type of TL_RX_RAM_RADDR_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_RX_RAM_RDATA_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_RX_RAM_WRITE_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_TFC_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_TX_CHECKS_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_TX_RAM_RADDR_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_TX_RAM_RDATA_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of TL_TX_RAM_WRITE_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of UPCONFIG_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of UPSTREAM_FACING : constant is 1;
    attribute mti_svvh_generic_type of UR_INV_REQ : constant is 1;
    attribute mti_svvh_generic_type of USER_CLK_FREQ : constant is 2;
    attribute mti_svvh_generic_type of VC0_CPL_INFINITE : constant is 1;
    attribute mti_svvh_generic_type of VC0_RX_RAM_LIMIT : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_CD : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_CH : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_NPH : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_PD : constant is 2;
    attribute mti_svvh_generic_type of VC0_TOTAL_CREDITS_PH : constant is 2;
    attribute mti_svvh_generic_type of VC0_TX_LASTPACKET : constant is 2;
    attribute mti_svvh_generic_type of VC_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of VC_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VC_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VC_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_REJECT_SNOOP_TRANSACTIONS : constant is 1;
    attribute mti_svvh_generic_type of VC_CAP_VERSION : constant is 2;
    attribute mti_svvh_generic_type of VENDOR_ID : constant is 2;
    attribute mti_svvh_generic_type of VSEC_BASE_PTR : constant is 2;
    attribute mti_svvh_generic_type of VSEC_CAP_HDR_ID : constant is 2;
    attribute mti_svvh_generic_type of VSEC_CAP_HDR_LENGTH : constant is 2;
    attribute mti_svvh_generic_type of VSEC_CAP_HDR_REVISION : constant is 2;
    attribute mti_svvh_generic_type of VSEC_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VSEC_CAP_IS_LINK_VISIBLE : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VSEC_CAP_ON : constant is 1;
    attribute mti_svvh_generic_type of VSEC_CAP_VERSION : constant is 2;
end X_PCIE_2_0;
