`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvR00/XInH4CequbT5uzqG0ReZ7mBJzeaZMdOyeaNdhH0Q+bD/UAEyAXqjztIL/0
2RTRkq+kLHObz17bWVr55jGGZ/lD2mx24J1B3WXE11niKWenwvtS4q/ZGGZ84JqS
8gB63ejrRs+ONn3BPBwWcI8t43+geCYNupY1eoMnTuzeS2xIhCvH7wgcQhrNxklp
RXhODwgirL3leKhrEElpu53TOQ420rT005YIELWuRnyZZls37LUwYP9u4Z6dzt8h
g8lKPbNNKvga1pHzzylcqw8sOOjqBOEK56qAAm/RgcKgSHg0F2kkL5r7LZmdGEK5
odMc8opVK716mzoUygxvNuXzKGqKbUKF2ifPzLq9N7QXavsBs6UAFhpMl8ngSML6
gfAP3JCPmpITX8SHqTMTt0SpakFV1prgAubOjn5IDJ72tpRklVb7O7ZyOSe3FjJf
`protect END_PROTECTED
