`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYkAiQP7FROTgPSB9W7OjL//Yn+0DdudrbT9Ce1oTkYdIRBI60UmiKKsfjjEXSgx
i8pjR3XZDOPfBwoiL/pnVEoNH3vyhYq/9qi7fLlOypM8Nh62WViXi84ozI6IzlwK
cfTQvbfoGQePn2VzCoAz5HphqrEf3wwMhcLhJ3OFPO6YB60+v3qOq6zOBC+4qr9S
snwzYdse52QFlDPm79jLREJYd226Yu4n+F8MJht6pzXQQgRsL2OUcVKnEGpJFJfx
O9VBovk6cOehs41tEZHrJgRaf8EOa0U9ExLdoncyd9KtErLcpLDIBm+2Dehzch1o
CX7OGq9dl34/jsPWLGtmJy0KZR10M/GR85iBeB+6WjF4Aq6v8xKMR453nu8Uux12
wO9NrHCLwPuGBwBQEZjhPa6EA+H/R2p1FQ5myqAM250MWHDu21U+nJW/LM9opG/4
sz180moR3wCupCqWj62pv0BGZWIQDNuJydPZfWFLqFmyCLRGZWafF9U4cAZaFMVn
`protect END_PROTECTED
