`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yotAa1BR+tro7G7hWX+c+7oKQiPjsQE6Ff24b+ELnoMLHr4uvjvxWzv1XJp2W0iI
9Vi4yn135D2qEi007NoeA9mjerzx9TV1Ym2bmd5CbBNEV1W8zE2X8efSjPI6KmRL
k5nqklJEJz/hViNWZe0Hxyg+bqyKBkN0IEaw6QRKrEculwEfEnJPU8UvyogcfMBf
WnLvDIRjQjfjNyaKMrTmAheSVyTyTiy5+W/NcNF+aGlw5nSx7pjbyuddQij1yyo3
DkgVp4czEx171vP5Fg6pk9bOg1WYXckQEsalE0nzC6g+se5n5GSqu2cHh7d1auyD
pCnk842Ku07SKPkdaqC890bPQ1YSXw1ex6l9PIlUntourQrTkD0+Utg0hflhtgIv
ZXA6i0xGtoZwcVbGMImN6Ud4h8mjk2NAtZ3fNbA3RS7qmWzjdXHWqR4saldK/20e
gzgmTscsBoF3CCpDXLpBEihwWqtS2jlRvy6+Nf5MTLIwY/ELXGJYKdRrrDaTI92w
Gk2U2olPYYEdPvst9IOH85pNJctOgtoKQIsZzkt3tl3GxXmymfCR1DxIJSgIZ+D2
mgBhlTbei4sRMrssN30KgQ==
`protect END_PROTECTED
