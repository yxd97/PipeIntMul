`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vl8LogAaASnOvUVLcASWQoacOl0tHJZpbtW4z68Z2WEgnqNhRHeJeLLUsqslH+3M
Rx7X8LTcKB0haYPAAtV8FC0ZZWzJGfVWvbqwKDUqVg+7i2oncWpj6bBFrlxXoV0K
z7DNI47cN3EDxW3uJTbu4mQgJ9NEuTtYaWHFLVvhslGSOf0xu2jc/hPfxWdhJOd7
1qnoxpCqVHoEZdGdRvVDKWatBLvadM0NjLH60Iz/KHEC9hk6J5AXnOfl1lgu5FvT
A9xYXa8q18K+bVN5J8F4wQe5+fY7KSle/8h33EJXAsS/q3Qn7l2alefQgSxq2Qw1
lzFFf0b2W6O0tpX/fwJ0gQdbDzNRnU5PaVoVYmg+xkYXFs8eahckKZQsvpDBtxjI
gfX6rgxbSeJmkB4w2SzYlM/qSbGQXb0wqJAwtIapb9jyaCyH4R/BJwrQ8HzJ7Kta
HYvMfegp434cv02Wdah8LURFieAp/4QQWWyhWECDDtlHrJY7OZHqxYKS5xZ8luAS
dBNA0pD+0J1nnIYFPhkr43/tYopATyjWzPudmRJO9qxSJbwLBoX47YMmGQnRvYxU
LjxX8iK7wbfDERRcD0WvYQ==
`protect END_PROTECTED
