`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Smdo1IHoFLwvsoyhuTn6D7ZUeMwb5swuUmR+oHGHTsZmuEydlrThXXJ4wt+a2xWN
i1ToJYzk8EuwRB9q/S0gOCRQOxg7ACXtc94nHtKO1M+ubitr/KESGQyGeCCD8712
Gab2j76qhz039qvFwe/+kdpxVHLQfUQCGQtGkSQ+57mmyN6vgoR1AM1T36pGAoy6
6snzgEaurZXlY4pA7IjM+PDwrFjKUZYvvYRDbgqAtkLVziW9WSi1VlI6fjtu8i5U
kQykFgkFEbO5qdvhlh8HRGkok5ZChmTaEKqoBgDFvQfwje2AlUnH5Lds4CrT/GS3
ZrYOdij+vGkbn1IckYrqz2j8w+AZcN4WNZ1E/5gdwxM2GbBsDY4TTiVL0nNXfPl/
alI58tAG1J/bWrqqQghc3RxHHGNg7c2vez/tbDq1nI/oCoP1MbWHzKKyhN1tVoWv
JYfHHaJhEwyvD0TAtsnU4FR1UendbEGHt58YVtaLWVUDuM2vjuN4+eW8WMiwEOra
6mwj+rnfE2iojiuciB/7xiqYlyWJgGHh+V0AJEtKpGE7w41Bvn6BclbKiOpLc5v0
lLkyC59d4TzdwfzE4yX7R/Z5MrPbZQ0fhCPIbbi4fNFV5AH05+NboEyQdheCMIv7
b3B5Zzl02LcaR0yjZQW9CwypfL+SfxghVzYLCqlHwSWdu51trGN+n/3PNDI7xaIQ
p6kLALqIu/QSiJuiXjtYd3PozlHZRTeKq6nDrGFCymTUcQk7Rx2hg1dw3xXtjBwb
zWdwm1YGCNsihLEcqzUll+x4bUPfUdKGS1i1rM2QKVfFt73HNy/8L/9O8BWhPru5
UoQqBK6CKkEqLa/jjiNqxrCnUEcGCDjab+WwM2MkO67vvvaPC97SHPLIVAtpZS/S
uRNNAeMo1ID3H3sNHjTR8P0oZG+hXl/5frrMqCYBnTUnF+FrpZdu/dpMYg7PyA5/
jjGYT+liwg0hhBUJWAN3rjw5tBYcgPBz0Dh2X62oIxqA0CoqniKalpvnEMD2Sv2e
vEB1WGCOajlFVqVM5miuAFxUaFLB4Y/diT8PwYS4XEmDIOWrVrBj4sU+IBYLRZWK
q99STzuaGAnjEAGBm7F9uNOD6jx/bNd4V+oNTzkYrfj6LVptuc3h8RblJl8B3KzC
Cn6xbx99t9XlEmrqPf2vyB+7kwUUi1McLfHDulzTbqCoobbx5oO0XLJIhOUbT69g
RqszLiGXV/AErEkEwygobcFLvQ8oCjUtUlUqVCsFT5VkusnSU+M5qQO84NEHO7VV
m9f/2FXOsbbQj96OPlJRfBuNG4wFnLjlhm1dqDGViLCO7EVIx7HeEawUZvHbBAml
9scz4kSWqbp15+O2urGzeDNXQs0x+U76j/4cbEx9bRz27tCbJ8cWeybaCWgpiGTz
/lxmzW11fUzqVGPASgs5BI3mnutiQow1SP6Zd0s2gEEtJaJq7zI+j8xc2ax95/O1
YaiW6vGFqQyTeXU0l+iABZZw+3AqCS6PzA9m58A26Cvts9ZFoo3LMi6GGgba1BV4
5uFM0Zf6o3cazye7VwaFzw3OnbDZH0MUcw9oRanklmnoZGIz6A8r6s0t7IOK4Rmy
mbvloE+j33ZUWFobkGEW+jvrOldIlkvi/MNMRgjS7gZHnN5Z4/ZU3I3MTUwB97I+
jbcM0qj75WpbBVhjtBxN4q2dgr7XQcwgnvj9FFBqMtylmwSK5RarXUWkD/TgGUO+
i1j/VHc383nbnvFUvX40MyE7liFvNgSVXk3dyAfL8nogwHgXni8fE5QuX7GnDgTC
nNOcbTcf8BiXwUEQtF09NVpx6uMs15KxQ7OKtk12xarHmnyz0Kk0fQRJQsCsIato
w/M4QKRCpPwXFTzVlNgvqbsALbh+Fc+F/YGyolHeyrQjExlyOTTQnqu/JJ48Umco
cz/EJ0YNRhPGWzj22zkKdI9UwPr+cC6bcoCK1o/1TzPv+zCoV5CebMQSbcg1+WyF
`protect END_PROTECTED
