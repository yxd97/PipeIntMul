`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oTkqeZBXyzZAEB1tBKN7M9+Qc1VFd6wEtMCg/hUIsAvq2cumUJ3COj2C5LJRlqgV
RH4ktdy2P/32/YzV0iUcIrIaBVfgnBE0TZDrcpH4OKFAZcAQfixw/U9/auM8gT9v
6jv/dV75IYEbqMNIsrVbZMv0kAF0kjr7foOHhk3m7slXXp84kAw7jlFJzKl17JWY
Vnfcy6ZKFLEUh3uDiK/CbqiV78iFpwxQW2nPvzVeSgDnv0NjkFCJOvRNZDFHsQv5
egU+CnTOPUkc3qQYwLIf5Jq0u2gF+O08FI85ClsY/iAeQqw+wLf9QICnWQI2N7Vk
nnqtcX9RHuwmJiFK3ArlFA==
`protect END_PROTECTED
