`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
alOoSGEKFFkfSzUEQCP+Upnk5mbhgCzPZpFy32jJhadUEXY+aQWFXPM2LJPnZz/0
XcugdMSdnoi+J896/D3f6DXIAhrAX3GkEpkiEX73SWHctN7nKOpsrLYcGcGj5peA
w8C1YzlrRG1mNPubL33t7hNaO5oz85/KgKRekAokaL0+yYy7vCcwExXcjlZyJS1J
YJx6z6zCm9GAGqYHJI4osYTt7+bD2j4q3NyZq/VkRRxCmTiDlxAq2b72pNAo19ij
RdbftleCgyuRFf9EYWYQIcWt30aGMilYRFKp0k2o7Y6WYcSOEiOz1O5YJTrw8lif
2YoEYIv7tdGANTfGDtnycG6iQK6M76pdwrdluQc6oXPxoB06AoFB+ry9vHhohblK
s2CSixMzMj8Ac2jgN1Rg5khKgOAuPExNTNGqgErleqQa1jQoNODAMO9mYuVZVZz8
`protect END_PROTECTED
