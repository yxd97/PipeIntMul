`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q067+k7CQ9mtuuRirlfyPjW4Qk3jiNYA5nKj0MfX6LtdoUQAq+85TFGm8ogVp9B1
Zl/MZBJW1KmsMzesGLDdaP/30udmSFLeK5jL95a1F96GeaXhfYAD3UpK1DTwn01x
hO9heKCRPEyEgBf6QemL+R8FqFOxfFr35b4zNjCkRii40W7AvIv4wl2SR38b+Rzr
7gjfI2NjGtJGnQigSrOnXcuBXJZhBVrAIJad1PgWRE6k7gvVstkg7LR5eASfssht
7sIuc/nLpkZmHv00hFvjErjCVsO/Jn8BcQtYeoAYx+BVY3kgCLaZtaqZaLmd2HoT
PPsfuIs5k94Rq9EzI38hDzEO9jxDti0RwbrpftU6+OlKbJF/PISMah7YCiww0tNc
bMumd9pxclBxUr9i/GbAam5AAKiGkJcIyQV0rW7C3Mw=
`protect END_PROTECTED
