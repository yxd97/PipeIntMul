`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zaFY0CvhxrlvHpJZkwEHVm9hOLF/P6T4zLehhU/345S6w6ND4gQ4fHPG6d9jCIdI
VDxtAxq8DfVgSwYbf+G0s8pwjp9dl5Fag3YceK9FYt5LvhpElZJ/kBlJ6IuQZhxi
MQbxfxoQA8FOFI1hyBTUMVPX2nfOWok5rY+3bPcrTZCZkhp++FeyOZVwPkNL8425
BN/HB/m6c9AFaHnOVPLgjR2nOXKfeIdZlPnV8lW1C/AaFtvDsF7BisRVLIpES2fI
AUASan9CWlz8M3l4cosRJepmTmRqA77duF2RrT6GBmJcdWhZzMSSKYQY+barpcmm
AxeXrmR1FloYv6FKeQZFoP5ze0uV6kGj6KD7wIzR/JjyOIAjC2mchod7RHLO+34b
NjUgcCXK5cRvle4ZSQFCaPIuflCmd7PDv83F+AGii0XLR4rymOAwo5CK/62k0VnN
iejfRq4PiHDKGBQr+r4iFzA8EkHkv1vsvcWw950aIYOI9cAAT6iyqbHO/tZy/k7I
HpYmew8thOgKD8PRIixj0z1tRZtU414cZNee52mio7lsSB3s5SI2W0baYU5gITBH
eMaBfiF3Q8gznfHijvs0Y/XXaVtoNBbkZrV9XmfOCJJyv2yTf+s61zsKWNYXtgRx
oj5o/pOmaJq4nT9wWHX79krxgeLiLB/7i/dsydZcnibNpGTCGBRQHRlWrv8xWGHE
flSYglcBNbQm67WfD+ESmGbLLbSMNcCxbLF1ggtcJzqb7KKupP4vlrLZvlEeO/Lg
mFE+8w2SsmtO+0IyxCShfWcvMsnYUVKYzto/jS2TaopEldLGuFe1SmzrxUgXHpyb
aZNa5hHBbfz8dsENoMknBZAJrl9Oj05wDFGO0rPuuTvk/Tsp6wklHADHZ4KZl6pF
+H7ncZ2324ND2waSPe7vI0toyOtg0WEtE7G+sT4Ehsd7JuIKbluXcWjcYSP4Yzuv
53MDg1QskMPMAJzRYpg+5ZOuxmzGOeYaTluunf0Zox8R7RGZncXcuocrEAZgpWnR
mRaQ0c7EvMs8SY3iqSXgvKfWHak5+oLjVASfjut8L1/M+Phs7j2Qw7QNhHptD25w
03UDfcjz/cFj+xfMwAylvQLwHe/Hv9B155uF6sMEDoYS/jxOJGDv69Kl9wp6EkKq
s/Tm9x08wvW1WsliPjlXjCuEPiwUO5lao0CjULNnMWgm9/FMTeN1AePKW3R1uZpr
L/Cux5MKwgY/UuOj9DUiNBE4QPHEUNvGeqFF6KVQ4BD5TpqdM8EXV4MAxVDnMzaY
f1cf2W/2BtXvIqeZJl1e2Q9tFSpylUIEgQhMxt2hMJvczp16LVKq7UfMv+yhqik3
Z/CJqHmIiNYsCCPigxWr07jJWuVGBKu9O+tdD/V4BOwFfxmCKI1EEpVeDTyaWOtG
Vt8CeHsqpjQARj2d7gXn3yf2xylRUEMv6AIIKAhAOPayaPmTiPv/WvS6mGCWlEji
imHRnJZTZ1fjogsacz8sg1TeCqhfG0U41KK6YCMZy5o=
`protect END_PROTECTED
