`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZMX3VcfvHFa5P8NEfI4dGSPLj6Mxfztp1hht2ZFmcZyB8XKEbhPesVVLXxdOofgA
9oXQTUpREVPq2DZEXt+vVHL3d14RnnZCM2dl3cMXB07DLn8s0TMaxZkVrGbHwbj8
3yoPoz2X2hav0guaNfGVHpaK5UJhYBhWl4xiD0y07iyDBTIU9sl0l73qbx8JNOYS
tS1En4Tu7jpPQx66/dGQ8epeVk4jzMc0pJw3tXqo3NRGx6H+F3wiUGvzt9BeWr6a
wmzA7jU6UvcJZZBbea2kuPN3s93+E6RciDQ81ZgbTBqapkBjE1dX6WqJimA1JF3F
/m7z9MLVSzspeB2UUgUYQ5Y4Uwl7AFZgcDSItav0TGhRU2KlmUyS6TG+p0tXQgmp
ebSpqbctYFfi2+qG+BH1AyDejJ69JPLY3FbsgRLqrzNmawP8MqgbV72se5d2oth/
/a+utVRAQG7qdpt7ttrwVUBn0OONgNSj8vrKCtl2DxNoAQhdcgMpEND7f/Y+ftri
qwmf5c1uMCaFfi1DhjtJGGKDLRg6cGTW1lQYWnEKxnc=
`protect END_PROTECTED
