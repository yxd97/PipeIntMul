`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gTPUWfa8CHBjyrCUWQDhbV7AwFuD4PbTGehtPRkn5Xk5FIMtgfgcRuetmobZOXO
1d/BoH2MwuknlXhyN9RwZy7EK05E9w1747dbIcusphRQTDG8h/yhj6qCJOLT/ft9
9VM/vpb7+Y+TwCkFexBGIjDJsfurOmusY1llvyXwPDth7hzHZ3H1o5u+/HVpU+Pt
bCSPeuCBXPwIOiY5qQS9ng==
`protect END_PROTECTED
