`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tprq4uzddf8V6R6/se5UQtbU6pibPq7dc2RqaStxnsqWTzwW6X+PZOu88RUZDvkH
HxRrpylNLCoNOGC+CyNGvv48kIXnjTja+avssNvWGe8KNquB8IZSF6JxhZSBp8eX
AGS8zG+XeymSYRdM0X5H8QMfIhSNWEReRAVvkHfK8aya/bQ0j0L1jBt+586rWQBa
s+fJ0bNtJX2dCSJfG9yRFIjgD64FyZ37VAOAdWNuVW8J/Ye69XtH8O7lxYA+MbOr
VSqoGVDji0OJolTNQf/rYOiHd4/etcXarFk/HwPojBdBXxdZCAzrEm7biSvNGpgz
ZQ31q5ObAbTK2NH9mffVG5ZqF4zZSVW7YdVS/cpIMva10sbtMwN4Gbvt6fyHGfbH
h0ksR3HCuVoikbkKnX1LDdHiba5arGfUf/NxgQaLwY+ZIak7j/3E7xRuf10vvIKt
ZdAsRaNB5cG4LMp/Zc8mt27/F5R4zHiOstml5ndOzL2Y09dSOpTqqIcM0fVpqbt+
c76tvN7R2L5UOTOUTSIMW2VmBtYPAIwQoM1j0Q7YErLnPj8qUwANbYFeZELwfdPw
W7LRduSKRmNqT+rKzUxP4lS9GD+RpmCCYABsznIBlYSbeoEcrR/Uxk9XR9u4ZUPi
ufLwjvvC6A4IjZMFN6c7/qh5bDHtUT/RGpipZZZy6Z8=
`protect END_PROTECTED
