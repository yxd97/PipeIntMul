`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLul8fDG+2U3ODlvzm15SWlaBXG4Mef/knjxnyGoYC23/pCuGbdCpwDi2+nAymuV
A5wU6ZKGtBwa8OIjmdIYJ+ph0OODCuKHtHPlxlAGFP9ZtoCodzis0KwhOek/tWLl
ECXSwtypu6pX2+bZmnzJs3azL1OvDiCz5fDLpKT4zoenJR6bQVnkw/370jdnY0yO
tf1G2w+5kSg5nLcuEBKPMCBfiuq145V1v4Mq80U9RA1W38Qi+znEE7+ZicMi0S0q
U0jvbeMyGRXW+TW45+fnxw==
`protect END_PROTECTED
