`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XFM2Rxz7F/vAGdn8iR2dhmEPJ2Nii4oIHZKb+58nPq3TAzO7L4cu1NqKGpHKm+WN
no+2wK5kWE+CgqXB7D59tYwus976Hpn1AMKqINYtk6OjUS07KSWHd/gl5PWZozMl
OS/CqXa1wQjxalGatdXFYxhvT1NgI+H3c04X6Odefduao8WF1pEef7UwibqvNcQk
7iOXe9H1OevCEOJxMQC1th/FRct6wUj70UdzXDfuS1Oz8uVAWtEmWod5+Yi10H0j
dujtndbPPO/UprDk7fvW64Ovu/OZTA/1Dlh9flfKz8ajXgCfvL8NWjjqr4Bp9lQc
RkIM2J7hIFZpdKfLD8QTwOtdHU/puHm51N5ZVTrhGnXlU+JMdSogu923PTE+Kh0n
t6qGAxVjV2Uw65sImaAJXz4XTWcVVD8jVJTt9+8GjwnO8V5+wq1sDXMm9/on/G26
4AAGgK/a3CIksm2xMitJ1BUHqCzE1yhYPpicgsMokFiyfn13/vWUBDIWaIreYAI7
Qztr0FI9YeNTmI0yvRzGbgiDtMASdE1KI8f3gexxB0R3lqiQzXN4Lppo+nFPltx/
4fa9qZOd6TqVlfbfxmJleusxQf3LXg5gqH8W9TGjsDxIuUDzExeQQtygvk428ahC
euU6jtVakp3al0SJdSeT7AjnF3hUSGJTB/ULBgGEq/VSgHRC2cz9aKfduS2xm6UD
4YTj1XBMw0h+JFAn9Oeg4HX4K4Nfd9GMws6B1yxP8othDlXdaIvqZcGD2qiYl+hM
h+NMV2iKl7DL7gjXAslZtK3f4CRp3OnJaYBPk7/EBL5QLxYo723NpkxExwcoTvzh
wJ7aDltm1SPcKxeKa5+QQpbTEWmW5J6fC8mDwfdXzlpnchrWK1yPOS4M5gwxX8SU
mVIptV/bDQnbivhI2G1Wepv+OVns2KqVysUe8Lb8Fmo3S5gwNcUihh1wUL+MWFj+
CgCWsEBUfgBRf+jOxx6kdr5jKAi/4qXfr6fzkTXCioRxNldj0j59kJRXgHwk31pB
MIFZ59Tqu54oLXsplMs6WEbRgd7EagJlwvDhgVkNMEmVGth9skrbOyXIbYI0H4fi
karsyB2Imcz7DCNCjQCJNLJ3FZZTeCo/Y/B1r5ngUZ60fC6n9EYl7X8sEYYQvHTy
+iaVMChyCqgCpFnzIj27ZwEwzgBeIHIBwFLOgWfBWroNpEyNydIv7+P3HeZW7rqg
/Y5IN2KJ2QIP3/V4lSFBwXt28d3D6U/0M4fBiP9LXuMftNGVhrwn9fG2uRob889m
D+7Z65CW+LdzgPb5g0g9h10GHll/I8NoISIAz8zBL8CkjeogK2EnOfSfEOOfTIbO
iQSQLZL8W44ThrswwkueDyTRYBI1f110jMg2+CbWUQd+tSzIxOi7CP7jvVSFB9mC
mqQSqbNqeeQ8XdthkLzG/OIF9lEDqQsTz0aAEsWnOKihADC6Ufi/LcO16qGcwer8
i7sg8rNrB/KCP5RF4Q5OqFMdCdHS3HPM2HelDPexVI9sdQiBhYLXLfUinbJ5HbIb
TclOI7WQsIfBLOeEaZPwKKRcEL24wRbxLXt8EF6m9rmUpc7+j7WB6HCdqn60aJaS
iFF7xAz/cKdSXgxXWqClwGIV2PxUGrGcT/e0j/Astb8RyG80NLBstD+t63VZRnru
QqyNYRrdFNDsRxtGlkRO9AigQvbEe6cPkJlCdD5DVfIximngujc+bRm8P+ZBzyMV
2bi99/3Hvva6UBuK7GN6CVSN8jtFdeYQ9dyEdzVxK90Z/81Cg/U9uaQWpevTf0qk
`protect END_PROTECTED
