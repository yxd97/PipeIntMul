`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d11fLMe6TQ5YsWKOstOWlcV53cjd+PP/rDQLfaIr2cJ56GJIz2LlsC0bZqORgH00
kTw3khh4D5FCza+E024wRV1cPeMdbZ9nqxDv03zxf9EnWrlnKASV1QsZwA/wrIFb
uku6vHvpHDXLJC6kEBPwdG9RLZtFObRBFuhP5bDj8eHdFYcu2XY6DB96wZxQn4n4
SSZlGVWgbc8JofRrTcllD3yAWHFSxxIDN3SI+6LxPNuCMfAwOhVXCk88bCJcM/oD
DhN6ENFjmtYXxcqi9FTN5Tk2zVLd/jjpfHgOhh6xZXJTx8y3LGt8+1QMxaUF97NF
21en8mkvBzAd9EJAAqJBPzD8JQoJTRiGcKM0+whNqyD+5M0TS5/RRJPYFf1pB8Wy
RL7gkvymj4QuFY1o3UtGYN3+AVxD61jJtbm0H3MvWsY4BOfikF9Ydl1kRXVqdnxF
RC/lgAyCPgG+OuugHBT19J1+hy1h1HvnXLLBPIL/3amhbiWsWeIuggKEgxegHzAk
yWzC6jud96GuFqapOmXKmg==
`protect END_PROTECTED
