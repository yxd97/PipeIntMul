`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+KuRVy1aI/FQRTBDcTiPPxJ8Obcx7kpZbBPrY6f7Gq0TB0kVigiqxYa0DfZyphtW
W4Xn+3XNB4vwMeRPPk0/liyvmA0M1Ig2T/GI4KG1rtfxwpcsPApfhE3Z7irY0msh
sbotMutsJoBISJsIZR3tB3Fk8t0lRkPEp7Zalln5jBrSOWx/YptzidSk9joyLT0/
pwmm8vVxzOyh5kEgKlfr6I8aE7Y9AFB4vZ34dlavGgdjD2ktoZFo0trs2H2U9zyg
CqIs+KZvEMAllXriYSGwhL6QFDrnRvTQnCrPQOuUlzL8CGNFFL9E0cKljEmbrhAw
QDIiMJIimu/zu3x7RU7Mx0/JjPO1uAGp2EOstevk7Boey6p4iQjxTiImQlRDNc3b
ho06BD/0DmBxv2Gzw6IpHGp2Jm4PzMy5B0SyQQBTuDkd0fiFMc3YtihSuoQ2MvA4
tE2HgaA/DKyi2r8PKaPZCZ17MUTK7NFPC2Zky5NzMKs=
`protect END_PROTECTED
