`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
51YRNFcIrLu0wXg4LTq6+Kjiy8MS74eRBYT8Ejkp5T2HNXadSS0ZyhofvWHwdlub
P1w9Ry0aiC0C1rZBPU3KWjct+S/q67W0F2mtl/5VIZIArLK6IZ5y0woQXuwnbqUd
Cwu8/1xj16RVoqZ856jLN9YjEu8fGUj8whSwluFhZWs/cQ7bPu9GuvApz8Wp6b1l
FJPa1+FA3q/LtscS++hMzqMjvEHbKmfwROWNL9aqwH8pCf1Y/VQ+j9DlsMf0/2RU
YBJVY76sXYknMOiD3Y30Hd4NRewSqfWRDTd7B7YzQVUy45VhqNdI/9tKnBf0DQqj
is2S+NHhXwYAZMD/qhlHsijw7UbNK1AOaYLVJUreGAcKYH+FO9keyQVgMCK8O9sD
o/vuRonlBO0IArHurUYVgyhhqy/F7Ho2/OuDCU9/HwGd3/4oGw4PFm7uWWsyjlXP
`protect END_PROTECTED
