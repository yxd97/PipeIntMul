`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kjf2xrB2hsdE1d3xJon5r0ntAt+qGxoH7rkyytoZAZ04r8KYpZ4xhmcjgAhCX2GE
JJhWFKdVTDi3HVWzfUzvQq12IqiEOSglxA6+Xk3FG+dmkRUMkFA7p1c3CatRkDtF
gPyzZhDwFgFvcDzSt7WbouVkcC7TbczcEP8ptE0ZXQEeKXgT45fz9gUyfAD5gyjb
j3JFUCYVaViaTLm6eNAx+lXy5gzm2na0TICdy5X0R9Ghzie2KR/z+ZZ29CWYrIGl
OBoS8FF5ek/Elsh1RS4XNg==
`protect END_PROTECTED
