`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0bQOlmFeK7ZxFMEphGjdTx4p/5pIssdm7VTnn/m1oqKkKVj8b1+HcAgOSnwn+OOA
ojbvnU518ZyS218f8LeGWZgGmpADTLdh3LnuH1wH4bBOlgJ7kgvuaGBjNk3yE22h
+SFZRX3E8n6A/1b4wuZMWQeWZebL4xOCRTN0SEf3qC5HEzzmUzq9cJQIPdj5/7ys
ePbO0nrKUo1tBUbzT3P3z4qECpfJmAMmvdtR9Mpr7v+pRPkYqY1yqGgpWGBHO5NS
vb245wOwZbaR3qhhfPHR5Kn2HQjfA0c78DpyBQxjpqTuDPpN/k1PraRHm4MxXh2S
7gfid3gQsKzhBaD79gwHpPx3HOvMukH/yyqENQR5/3HjLZubXoTmYVoV+9fiV4Am
egY18rZCrN0cUg/UKCnT87p+6YCGStIxxpjONE7w85dD8tBntq9Xq8xZzXoyNiEk
0tqrtjSQ8NSJY2spTyxzoxrrcTB71ENqvxSWK0QtkTXyZ6ClI1FYEhWFts1oic6z
c6O7uDiEm/xYmU0uWJUvgSbhUYmz8H18ncpS15M8Q0j1adCLCmECMExBF+rbZ2ib
uYu4c7HgPUJyHMqO3R/IkYv1KHg4pKrsrHkp5S8+x6g=
`protect END_PROTECTED
