`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TdcDnPdZnTOstivEtBnPIsnCMaqRbdpooIneZRF2BIxjBI6461EOfG517xP9b8Mx
5rCyZglS4qmOqALIiSsAzk975Fr5NuCXaxsvJdME3qVnXUv54uVfKkMOQUOceA0Y
rZbhm5b5Hao07VqDW7XflFYmH4mI70LL4L8z1INmcBsQfZ/UqHrBpYtxFB/6Zh+h
8suXxFqh4fG2YU9vKlhcc4Yu01R14CkIjPocjFwLtdgJrbvtFttxSxfBmzTbm8Lu
T+po/TddweVMKp1j9rAJSUzfbHXtsX8UqIOrbzJh1zth+vQ5z+47xEv8QG22ORyF
ofRRZUTCjNLYKfCfaefHLbfd7kqU+eEQNtby4/T5YXQVGKa1jlm9LAVy3uRX2Uk2
p9Y8U5pblDeY21Asqt/VbI6iZqEu4/d0+Pr8KdruusNOCkjpZ4anhaQWGIU2iboj
eMHYAwrq9U4wQywxVeLq04O/Yoxwez2To5BLgqp7CykZR9xTzOsGzvkpYbKVf1Dw
wQLj7AqXvvSjNGawHOxvDH4UaSEqr/TSNqeUxCIjbDBKouovj0qh5xvtB0PgXgC0
dYCU9trjMkcKBQGHIueKxsJTIYGEQgA2HCbyB8uo2n5fL1keQ88aJBh8O20jdPNe
var+Ui0GhwXqUX0vUz3FePxDvz0F9AdMOS9HeNDxetBGPDr4lvhHS+RIEUKDLf2t
JdjvXCHyO7xYTwc85PUmM1/bJiPyEE0TQBRJ31+mwLp59mNu+WWAQKZoI/3nmin+
WOPzRoDtAQLbCNW2y/HRgCQpdRVvUHhoyeQT2O7fxl/ibxm8FOXJVHT29eVF49dn
+zeRBxi0TNLBJ0CxDmhtKYigq2X2nhOwDmmtvvd2a3iqfiOkTPcI9dkHmEPJ1t+u
2GpJW94H9PBSL9PvWqPA0/y1V5QzRMgjBNKNl/uNLWl4+mbi22LN9iZ/FugCRAce
`protect END_PROTECTED
