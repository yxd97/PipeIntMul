`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVOA5DS0xFGnUmK/t8THQBXPsHHr+sPEhPqtm2jLnbb8VKMnp0P156GT08lfrqnq
PY8BD+EKQrra3DMZuHLpiWoiDHeKQTaKW5VpLCcGuxtHE3xepsFNhguYUzKPoa05
+WudqcxJIbBTprlg1AV5HXLc3bzjSQI135CKa8ENCDBH3OW5TtNA4qSLrbH82Yyp
WdRbwoGKyneEpD/rp3+nb3dh4VYRf6qguCzMVBqRfr/gqFp3nDVjn1tD/cLVD7iI
uo9D9IoMFNzIl8HmcJu44mHhE2/VnaRtyonoN/OZfVDWlGKuxlbPZr4bTOavBa9K
QlRmE28GoFIkjibfnHFkT7cweJcArQPD7mnAMZ1pi+DASFcoW2Hm5m/90Q8E/Wiw
`protect END_PROTECTED
