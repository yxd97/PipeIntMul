`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bERtHvvdYkCL9MxUSwjmO3qG/IeobLY0jYYrvzNy61Ga0U8E5UQDECespYVqPM6
20+MUrThRKOEn0D5Y8MZSsXGEVHyqVDvN26YN0OyTu8HNd6JRVSLVrvz3sUkAa6v
AEsn7+DkokoRNuSKRITM8G3prXRzTr7sALXAeQSErqjHXCmv1kp7QuJT8T+2Ee/h
GB2jDWxAqqAoE58gv36qGF7+wyNWx8rWTw7iquCleJv/0fpncVna4kIKTF7AZeRp
BpGOZxYA8rW1wkzEXtZx7QmvG5fQdUAZMwPtp6YQmXK+EzBd1lyxESSos+1L5QKD
99eHfUSVmEPjdqwV7DgZvARY+1yMYMW/Nwodjo2PMWcI0GlQXlB7u+8Zk35FoAXL
gPLLtZZt/ERTvelQJ3y4odU8aXVPV5cRaAA1Tmi7tQYv+/CLzxxBD3Ly9pgpp8yp
GOTguFrivKYLd9XoRA+PyKJS8wdUeR3wqZIo/I0GcoaTNGcVyHvdV+4MYDY4EdzT
9vS4Ia6Iv8voUK44Krwkcobm9uGFdiXgdwMugXvQllbIM+ZSesY/omSvcUZtJZ9S
CYIIur7oZXrwQkPtrn2zR/nIp7bJtVrQ+yqkteo+rUGL1Q1vk7aJg7cfdtkfVKuc
tifk0FJ2SPAhdavtiM34Ldr6r5oDgkm12vaE19MRZtL2ygx+zbxQ4XAAiGDmwNaS
4N/CcBEkbEN0BaCVpfDEQTjzE2hw3Pag/DxHUlxcIK4IfuRNRuL5Spqf+NU/zImn
PCTMq31vU8bTH0eOChaTG50QsNXYcfRncO1gasF3SZxnJL/YbCqshGMM62XP6dRG
7DDsCdGocnI68FYlb1GEwjfy7PMCleFbpJh8wcYk6ro2ZYnxBu44d3zIjR2l9DL4
+UgSLPJBP/c7yaiojm04CoYlXFwLAoQvloIbPtwmNcFn7dZYVHV4eRUHjUgNXUdb
VjTqQZW60zAVYkf3itmTKA==
`protect END_PROTECTED
