`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+g+6V3sqKljMDiyGRYTuLYfqHnCjuuffuHhjT0whwmMzT8CRidVZ5Xu9Eq2eXzkR
nmJ6uiHHrw+1x4FLgX8SoGmlo8B035DiJ7cNSYimBiWm4OPWGqSfxc3texM04YXt
Vs2e7fJIyEFfLVcwi5fonpbvPLkSWNdvT1zugPqleYdEbxWQTpIrPu/eahR5J0QM
4xVYYyQPjU6psg/uhy957JK1WKk+J70blmZuQpPp2T49blUd10ub/LPyIZLjwITX
x+lG3xdvWTrsk3hVdGsTowcLK0HFLTMc+hoe++OFz9z580Lrcm1MlEL9JWjzrE6p
FFLCjRBgCP85zyq+srg3Kl/MCl23L7zlZfFN6g9ntrAgDvFsjTuVwViyNdvJbm36
HugNea9I4rX5CPb3xcVylb+RYTZyf+12lEKPOSmGG+IBEGFwZYq4uhsHnQeqjFzK
BImti1wfvflfm/aMuErpSdLqyrPAn7oJu7agUrvFWmw=
`protect END_PROTECTED
