`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pttDIvCh8BRH+MiWzwYpfmrjRxPuMCQe4vfFhlVJm9fpkx1jw7+F/qXFw9suUUtq
vUT56v8rZBeO7Q1gFVzJP+ZZn5TRpQUEAE5DWvoiJsnsz+0OZtoI3eDR7Y0GgAgL
Gc7DsVP27tCkQejsPY5svHQNtZWEwybI0NxgeBWXoRHJHaRj7H+yu3ltlbErOQmg
6fnW6pgEDTdPVIL6KhyjNtIDsU3YitwQycKp6jUATuMUfI3Fzo4Q3buPgzX19gTt
zl4adM1hEyU5SgUiAhPcfivMDv5PlskNrLX5zk58er9Jz+bbP2C4PtGCy3RLXR6c
zJ1SGymsRd4bjYRy2KkjcMVfp4FXYcLmijorCS99ry9GgdjbpiqjqEOqsuil3oBG
gfWe0EjLahtAYpMJ0W5Pi8xgT8jxw6o/0cdEaT/rgIMPfs/abTebZaVbS3pMEEWw
lWhuQWGtLgRGyf6VxTo1Rf6eXu9ZOkzag2MBZ/BTDOC7WqkUUfsZQ98RJiKhdmiB
pdj2m6TBUhQITtlt90Rf5hnzBNgPXepQQSsKySBQioZjx3jAe7wWcWfFYLnZ+1sO
Y1eyyBE1Bj/elT1vfXwCcS4zIDQth953d7EYG+n+laqY2zTqCsHGZ1VyEUI6uaZB
wE9UUMDoYrgi1mFfaoVEd9p0Kr1pyq9/HpGCrWOYgdI=
`protect END_PROTECTED
