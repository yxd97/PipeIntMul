`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mhQ6BTMs7VSp9lvO8Fio9/ntNdWkXjxaTlsqtv1n97ZQHGf4dqdSgkmN/sk6B1IV
XQU7YjhD+g5vskz84h804qcL0nZcK+1KcosUxB2mkH5VfzegpLFnKAq7pkaCFgUD
/4qZqpIdvOLyFg7wNQzeJRG/8Pk1G0Yuq+ZFfHQL/EFw+0JELMXMfDXtbtDBf3q8
4W/ksJvZIwV4kCnBv5LUt5zH8QN/KiasbaYp8HVAg5AwXKAWZuQdlWUD6L4SEsjh
4xfmWMn8P9u9PT8RTKMvmQn0N9BI532yHYyg2bPEta4Fp5p+gj3/LgR66YawdAc1
0IRVSGhbbT+5PfrSZSW/4GFZ5319UaWOd+Apd7XqhbQdbMePH8HJCC+dTMcwifFi
xvGmLdEGMNwAy1JfriSztiQLV6YaHhZT/bOyqNJ6Y0q+4Q0XjU4laMVm/YwTS6F3
reQhM7xki6xfyk57pMiNxe2pdGBGyojWIp8Wy/1P7Uzilb4RYQ+eCVTHV7Jk3yPV
T/byUBcPKs8/Z1tkBC5ky6MkqjQDFSZGbTSKA7nCcekTsORa9aTRfYi16T9GVq5G
g5qp5K9ZC+pJPJ/ENV/pFNojUMIJ1TQQW8AoybXnOooiJZRm7lYT8nFy8nZiDdUI
odalwIEfgq0gTe5CpssHOknKtU2Xd9ca5mEdg8uKAms=
`protect END_PROTECTED
