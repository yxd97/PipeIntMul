`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJqVhZXABwFdlcopMgAQCJIvDS/Cgy9l2OStD1tJ+nJPlQ4shymgq3LXwVkcX/aw
PkMC0oeVXlvRN+LQ50OPmL+3iJ7lH3QNZkukPpwAAWWsSuHFJstKNwKM7HH3cLAj
fuje5RiwYHUz32ZOLawg+5b7Vpa91tE7LXLL7EcqPz/c1new/pIN3FzWWCrl/ScP
tIs2Zv/G+M8aT83rsXRzyE9JUbbvJTVWnvOwfdWEuhFSWvwvS0/sNlFcUP0KLpZJ
QkRQM9tafjELNqSts9qBxfqRehkebMZRhQxlcJXI2VivajQIHhNp69pYrw0G3m2T
NSkX3f5U0PUoE0ep01k1rlj22vqXvQpUH/pEqp+MZjNn3aO+8CjA5ligsCWRz1aY
gumnXRr4DKLSUT/5GEXQR2jP9ka4hNCSpPkH3hYyG+y+alcO5OWHKrpcO4ohJx9Y
0JqKiwdHRpZ+Aj+mmt/xeLKEm0JIMIrL546FW/rlFIvDxszgtv66bSJUkCAbzi/H
beDDKsVxKFD2+H9fuygHHYUFT364aPmYgM/mQ2xYB4KEusOqw8I3kOEwGdeqU52P
Mvj6KqAnPmo/NgpYEXRaZsBGPd0Q443w0ryZn/ACf9Z4IAQKkKu7DSmI0c8VYsy5
+h/Lc3imBYupoC5uuFoRi/mWQTrJDhBVhGiQfvgfmPfF7dD1XKn04V0rp4PnMrkJ
LaXHEElq5rw7uBx/JMi/vjH81Lf3FZDoZIJlWzvy6mwhuSMimNvlFE2SjSxzfgP/
v9ISkfUW7XtsRGnRw5BbKrK7QkgxlC4y5C1A9QS40PsJ3KI0nrAQnoJH5pOv7us/
mxM6rSXppLajSZchEm+uWf1uQFy8GUwPLHqDFGTiB1N/4xHJrEwZ4J+lVfsRIw8v
kx1LUbV55fJQfjlY4uCyKbV5JqeuQhLlwcEF1pjTLx367SHks65Yh5kch7v5ZB5X
DF+9BRlHv+tFRrwFy38HZ8EqEEu4BByyx6mAUGigeb4g7/0AXCr2F0cdUabUXKG2
Cn+uGGtMyfT3XGZExFOoW073b01J1BzwbDR/k3286vRG45dQ3MGwam94yK3mo3bw
CzfaRdsVIQD3yLsYopS0CLA++cR7BMahlEdpFmH3vaY+chmn9YLLWTyj+kLuoT5n
`protect END_PROTECTED
