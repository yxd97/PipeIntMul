`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vIczTl+JZHpHqiBzrhF7904ZngUX9zWoV2NxLqVwMiz8NBuf1MuEqL17sgvJTz1k
D3i/TSA5uT837DUF35A3FEvdDoQixKNBPzvKUTQSxWbQpTbJ1NazGboYdO8KoqRB
IH1wodNIEPCSiiDDOl+bEiC/uakwPoWdnJUkWt7yF2g0Eiy7IAs8ubKs66E1ktry
yM5kgNbwpxVVvDpkp+sK9Noj/cqh+7qt7TUA9azJmKSJIARrca287OJ3sxE46f2g
Ol5y6nNRFrM93p83ro7g71xJz7LSfMGmxBlPV0+OgVIO3QAWBEX1+5jum+P2xzDg
Nwj8g9sXGb30ec/MfS6xS2iDLtkC0LOgM3wazL3NT30bf+TVTvJODzynmozG269K
3tNc7VZbTZWsyFoF63cG5fgfKTvx0XD1zzwi/K4iE3E=
`protect END_PROTECTED
