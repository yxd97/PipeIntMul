`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/fmX7+oskmQybjjvqqTTyyck9iJDQ417c5kUgALKUostWqt6HV7lKkybcXWZUM8
Lb2rNVEgVYLnJRFk841gV+V6au4OQ0lAXOOLKyc7irxn2xlwSo8YQod+AO41bYrM
Lj65YSMCBemD8knrhc7afXAw1JOTVIQKUxOpyeIHaV7OxwJD/TlyquFnlZ3IR96Z
8RWgfaTJN7F5bHLhNjBTcvaSL6T58Zu5anltNbDDDJ5zfOuGMRDXpacUICLi+lGl
n6h7iqvKQ8Vl91/ViNXxhmd+xBiYgWiTkTjiZUXCpFGGYbW2T04IFTABwyu+tk/g
mtTalQ/mcWDPxH10quenLRWr8vf2oPlFp6kg0eeD6vQpIYSRxIOmM+gptR0whFIU
iWNGdbAHB7FgL8ZfldfXjnEZmeXM3DR2I0bvrb1F8UWhfOZqTl7KlepVkxGE/R2+
xoGTvtxEdmgUfcCC8qQQX+P0WvUcKuOhRrnMNKErfJqkoVWNzckCO8mjyhrkCMHH
VdBNhv1mbVRJjKnSK+9+DB8ZQPegYQuRFhpHY7DqjdGLoKUtg+l+TFGJBdG4y/Kv
nSIITMaEjv9iL3Elm+bZwi9Y7bgnEJINzeIHywZ2h008JjcU2JMjFQlOEWUQQuML
o7CEz8i0tyiOqa4Xp3SAWaud3bylwGKbq5o+pjeg0/w=
`protect END_PROTECTED
