`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WNkG1k0h8IsymLIybECZSFSmg4BI4clZ5zMJr5J3/m1pCAkwjffVq4nqoxQLCdz6
ysgRYqNPCoOU8x4tDCFZqaU8Xp9yqYUBC80RPk3vtzpvIb3huLp9xM0zqm47Rcls
bRMRWJ3+5vBc1/ha1QaUhNZTfEqckinDr0qwENwxVTuhcdp6Wpq90pZ7ho0Z382x
Edz+4UOKgWqCQLkRJHgQEojyXhqdH19qt5EHe+SgeJW4/lBNTd9iigTSLu2JSYnQ
Q0C25qDzZoV68UrW48fbkOkCC08ssf5NS528uMNyg97FWTrD7gaYmoNY5FINSJVK
o5aFQtHSCRq/k8702ir7Lg==
`protect END_PROTECTED
