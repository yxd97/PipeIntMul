`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrljOyLpOyjNlFGDvXFqv98XRJ6GMkOuhv7ynLdV2DGmKSeKQk11vkI2AG3oQ3so
HPCFkWBLy+Zx/pHwp6wb/Ddv1FM8zxYr/Kq5Edx6/zgKJQC2vbCdZVn8MCuJnMLG
naUdK3gbbw7/3hAQu7ZoK35tOKCVn6WhHcfMgCUM39d5IZYuHqe32CC4xI5n2EXp
foWyLjezhEUUODY+cVbbo1/ohW2XBdlSqCAhVy4IHowpOYWgJY/+hXgYZkxsZ8ab
0WBbTKPhD6eesE19rCrNxO1r/c0oVA6Qenp2Mv2Ub7p3OdcTOocEbMTxD3GhdNWs
4VAItwd0hz21K/gHA5MdhrYb3ysCBpjznTrvuCEYYVfZKpPJKobzJF4et03DyVTT
wEcnBpYgyPc/sWqYTjqe8ZfAWXHFbe1BdK75VQukDS1cxdaU0CHw2wnlUVXL6Jwj
D3AGUtemfiSyJBEjHQRnHvQdzwV/wLVqAkgRh1iJM3pN8g4nFWhY9ehh96mqrLJn
FiOfJXgJVi1I55Ba0McHUkktHbk26DLmy7/86WE+aJBqDv9IbN/d4qEhhSqDuxED
URclySQ/6wOqv+qn4dlN+wMejvIFHBhvZg0+zLnR4gSi593uGV3VJoAT9/j0wtHt
qF02Yge9iDhukQeXrLGHItjBcwr3+VxScc/g7fltZhYFxYij6HRje1iKHYDiSays
gME2pU2wjKHgT67yRXI9WA==
`protect END_PROTECTED
