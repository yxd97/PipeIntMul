`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ius5L+MZmNxQzz185W3cr6sNWnjf8f7abPTWBL9XDZXNMU/+0tlw/PRkdJwseu1M
FNFuv7FTmNRBc6RHUIcyMdlSB5t4OsnZOMuY2IAP7q6zhQMitiARR4qVV4e0W/zb
0WxK6pCjmCIZyZ10Y5vX3d5OjJDbKKbjJELaZmpeutc/RrorxUuO4bYS46tqQWwh
QQZEF38sGf5DPvgDLpoQne+Fa3u3TAcCNA7WnBTNJjKuEuUhsKFAjv/YT0KlSYW6
145gLgJoMQZMMTqyJCfCH9f/AKBMWWQQqbwqufnTNsU6000UADBcIq7j9YqIq1bZ
pB/5Fmi2uUbJp+OQTKVY/FPw6zDpSf2eiLgDcTyqANuFWqP0brZGpQHd6XtQz7GO
LUvrLa3cmVtGAnvTiChVQ1TVJDD3zjG2a3AXjFxVv49ESqijCa3+fjiFm0HZg62v
/oFBIASJtjqF/I1dR2jKTzqSSvT+sct+cx+ZXieiG0IsPMLFXuc0Sm9JV8/Mw3j/
uvSzZEWZp4SLg6qyj2GmmMblB7xzPV8nOfgkbUdNPJEPeo2erXLDXuxxfiaMQCNt
phWZxfQCAmT9Mm8Twlgg43i5IV/D5nBzWGPPb4aP6KfPEXxmC3oUHBpdMc8RPEH/
EU5qUPras56AeKTjPrkUwhz1KD6i6YTmB1kkEidDy30FizzAt1hgQP6QgQ8oXSLr
fSscolGHxRW1TCObmM6c09Rq1KiDMSmyeBmIcrEiIySrd9DIlOTELyJXKInjq7qm
xKSsu8pO5auKpPB/GNVjjyjKR4gcNwd1OQgq4GBLdFruZidn4hgHc95G/VFkdT8l
sfFrAMg0a3Ua+odoE2e+DOJJ8DcEydVZkiHDpXmEOn338uDSzhOXyjfr+Mwjf23y
aW0Nu7HFU9jHtqkyr44t8fRyo47kKNTyAzG6baHiCxA0S62ZW4rnC8DCz+z2SXEJ
6tV0W5H/fpc5fFJaw/zqkpmkb2W5wcBHRmJlD7pDqoyjdRvxmGWcsEhZCYOjDWVC
3drzzP/pEDh2oSJMij0bwKHMVbYBcP8nuCBwJJv4qU222Ydwz0YsimTGUeajHdcP
uLv/dlLEEKptfwYa+To9gUWBgqgjPSHeovMT+x4Lyc/bZsMB7pt/CFKqLxP5WxCH
uwiekbTV+B4EtGsmu8GTE+22V1wLbxR25yMAj/8tzXvO5z0Egy8Fre9JWF7CN6rF
da0vA/uzVpwywNZIMvcaxT/F9GrDO9N4NRPFmNQS48Qr4X2ZFB/6pf9qUnYApMb+
LUPVu+zbyR/fV7T/Z8AzpaO5F1HhV/aNRZXd5iTD+DeRcxDfhk/yEmnuZMIpTAiS
mkVSnfWGw3heRt1/sloGnBOkspsFYuL44t5QABp1c04BEAAj+EknpJvklCXOnezS
Gy5KSiZ7uOpka/s0ng1zqbVuTDqaSIN3LfTShzyz1PadhLTFlnSP2F5cp6+nV0pY
5AIclefm63jrYWX6mWo7n/Hr+BBirgLRvu7Gjx92V9MYEFYo1SnbR2OZqT06jKj3
GfUe7+iO73TLfClGTc2naKkKe8GHWag3yeYUt1wqppRC7TuqwQZRJHSNOxm4BAIJ
3+/59XL/3hUtH7gxqiIZ+zfAlEkdBLJG3GMHd9jd0kwWm4JpHWQ9/A/gFsfCUPWq
x9Ydp/rh9EGgGlRSrMWGU7hnfuGpKj1deP0YzYOs18SUrJ4201fVBRfspSIYkHA9
CEhKCGeUpX/+fCNBimNCw7inWbqAZA5uFjud8o+fwQuDvMPogkiBo0eigELDXpCz
QxQ/t2IOOvksPszRikUUcgfv7o/UTNQ1wgWjLqQW+3lz4M3mYsUY6UJ7mDcAo4r+
bBvSoWTdumMpWo6ldfHN+63SYJrT5ngxIjo1ahO8K2dOHIUJ1bpZ22cQIxOIEAhf
OuXJk4k7oT9ji+MOehdATQ==
`protect END_PROTECTED
