`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ri6L2uuUnHVD2aoJACjRCc013SUQeQQJbugBljM1WF6E4PSfAiyow4nbtz/gdWbe
g9j1/A2DtMnriQyUmhMDLaUOdx4wBTUIhgkGwRuqK+dyN+jSxdnyYyvrPnZfPC1w
U5/l6UQff4CYKebn5PuNcLor9xKb6VIRs9i7ZL5oLZA407bB461Uj56YtoqA1Gvl
Vys+wa5WhQwvf34Il9KSPhcuHbgDnnrU9FQno/TgqQO8et2+EPoGIllA1zdf/Gul
QRJzPKmx0Q9EnIyAdmXmSLv5ri8Mxmka/CRCsE7zBjuY+GBSgY9bSluqMO0wLlys
E2FndjBCHCr/FwzGEB5/qgD+fbXCWmUj0JqT1Xp6REOv6fvcT4TG6wJ6W+pWiuvm
xMSgQPWt4NhAmajJZR7dZDXDzc7PvWVnUp5fBJylo/uP12sQzNRYFkPquOxmsrAy
NEdwEMUNziGA5/btDWe4bg6Zk/R1kDrRcr+i9HXS652F7I7kgHtB1Yk2HXjvd2oB
ZdjOj2VHjN8xjkQ3Qm1i4qeA/Y3+UPifQP3AMXJYYz4tbnxxrkB73hFRfcvCt8rP
JjLQ5M7U+R8JDVXzkfrK5o4s3msNkfkGXwkbeKbsMPQq33jigpzVRYZ+EAE9saXZ
ubVVotqEhq9oFtsmu42/IgQp5IdNoqSjPmJuxyjBrD4=
`protect END_PROTECTED
