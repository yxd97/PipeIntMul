`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGeslSGN94vzqPw1nVe1M+NQsu8rsUYIKHzh77V+L3oHEO0PBZQgA35Utb0z89NO
G6SQOLPXARmEGj7OOU21IrEKwwz3quqT6jhFk9U8Y3aqgEUszSfSQ0Qd5nHqOEKn
AB3LHgMrFGVbqwoe6JHYMwueRqz6a1uTHfLdgCQj6cIaepzhswT9pmb7T/P7jNEo
MLYq1IuMLpFgenGU1PNnBPeosgthlIAwvmeVOVg6Pl+IlVbbhdS9fKtwE7CJdhwx
AaisXrIEnbN+PuIE4J/3yYlCngZY51QVCvWBrO0xC/59M5urkBNDM7koSQlJed+l
mVIGWyGdt4+ZKgnz9RseQQ8Hsc8o4k1FK/4pNAr+fADKXrXtMFZLm2LJkVp6YrDR
NQqYWrg8sAWgL994dOwhVgUT+lHMeMWVUOOsDEj7dbHxhlG6DPzxjUZfjJcwPHzx
Wr+Gu0RRlPoDIhYKewBAsqhRLxUhmNbZhqdHkBAbM7aDH4D/shzwWaSgA+1sDozS
fZmGjggczXHG3W484CUMRxF5btHbGGK17jtOSxt5bekdLiKhaI9bwSKGKzzcbf+f
fzHCOPv+Ql598u5eLo5uOgJuKVF/CgW3R+uFwxlRL9dGdcFjLvlIhSdOtEaudeT6
VUD+jo/NvhiEBJnTOgLW5GHJdSO/gyEb5HasAKg6CoStOu3jEoEmXggWWmxWdyU1
5OuNK0068Z1F+1TTyNP2zQ8EPlRm5yul2oM/kBks7UlYOeMJNhDA/GVgkvPsKDfc
hxzamd3sUGJ35tipLnQdvNhmpWU1gslCAgkRgXqAZKvfwXY5TnkttzQMEH4b+wnU
8hj9QQnGwF9eSTM2xYRHAZNTY6NjrPog+DnCM3jRSgzF+Ba57aSc9EMmk1azDqnE
3Q8JBaetpR75pFLdh3dKDRoJsSch7/6YbsnBe7d2nluECgJsR26lvFgd8Fbi/G5i
zu806sT9HVMoys4knbDZlT0P8LThZvjjbqLWLcKTcW5nlj6kl5MqH0tLT46951Bb
ngVP+iY7oRFWfIV1GG8ya7y7CS80mibGWz5zvhSL4aux4uBDpL5xEqiYiUpXgmFn
dDPxzMavxaSotZO3xCQzTdC1d2DKIhN0yBYHjfMtDSVTJxquqvNMEONpGSorThfg
BPoUBgQfv81R1UQhYI2fy42aMraB69S3YKD4Udug6D8QoFvW+nSxHJJMG5Zwyjdv
Y+UOelhfEAcyksOHEDSplK5kB7RRWKEGgI5qYAFwmyH5/iP6O8D2G3BWX626TD6g
kFr87qhXFyvyXypTiYU/fjJhjb+p8aOjphJAhsiGQnN6X0PY5DvficENqY5ln9SI
7bPFCk9wYLu/jokthi1eb0vQdQuHmdGcM9D7kkYaUrB8jL8uON7rLxbrfMw0wM/F
C4UOwKgA8Tb16YD85IzuHhA9bDXZVbmemhhsyN9dYp/zTQ3vHGns1axfs37BhFEb
9D4MSMc4Y42ramBROtZ8NMPb1l1RFwcz3SnRXmpkdwA=
`protect END_PROTECTED
