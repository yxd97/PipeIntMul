`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N2FGKO9lihtLviCJ2dInLOden44JyxP5ePS6EE2LKwTziCYZPSVFhGc38G0K8wEc
FPWaaeFtTXQ38hvLD2J0RQVCFf5QBvf55l3IgAxl/av1gCFWgf4wHe7dm/R8lWYF
PujQfkoAjiIbB081ay507jnEvaWjcjZo2Vqqp65kVt2at7h+uQBcQ7N0yTLl1I00
HCit8rR3S+8kyn04CHAWKEfphHfUbO1ZS/SQamnx8BF5okN7KTE/Sj8+dNTRuAy3
cTgnjjTVX9c5S3Z6/e5+iZ7Uy49C/tQsGOEhOHmPfFEzWrwi6+bPSOxKJVjIU86c
qiU5J2rw6UDK/adeXqTBEC/uDuWo4ydsEM2hrxRftYrLmvXh7z8Q2SDI2kD9cTkU
Ykw/Ixp6QfNq5WHCdvJN2/za18AT+XNTmyS3A2x6vciTZLD3Lbwq0nrfCzkmimxd
ikcFtJkgQc8Udf+jUKzeoimwCGp2VwUemSqAvFZNijR2vimjuYYulNTZ1TjX/+8X
4fLLJIEVQZb+SceRk4jNbh5iNd/Tw2iqKJ0RezDuAsod+xhYo33FxX2alKJ6eX+i
UD1imtpn1t82H3l/oSeRgPgr2lLiSy2KBbZH3WXz/jaROpn7VyJ7YEEBTrTeYt1D
DI+M/7RsqrHW+hoYA/G3QMXOGIjzgU7W0HzVRGyBmSYeHD1SNGe6vejZPzF77WjD
elG0UtQknfqgLBJ6I5VJPKDtgEfuS2kIUbDxfdUEyTGmXWYV0F6DbCSRTZut4Oox
VQQ68TTIlm8vISjgN7UGTzu+P8HJw3V9VsK8s1FEl7f/lc6c4cWmKyu6qOwFo18W
gLAKnpWJBi6z+T/5oeNLpH7mcMkP7kbXTkqbqNaHG2kYFWscxwu2pWjLaNoSbgQ3
fv1oGhp8m27FWRdr3JDUY0SEzAw5ROsajk/dpPfwhOCDzWBvCwiaW6GQEiOFDGN5
AuFDprZg+1hVz2/Wx2xpb2LLWEYyNiAUUczTRgxBACwNQQEN5+NuB0oHwbltgUrY
mjIwrqLVAswLWolN47SR6CHCwuR9u+9vtLx874VTp48YksTapcjKlerfgebwmXi7
OLfeuvnBfK8NB6VmZhUSpyS6zjirNRdOt8Ye76iV4m2ItgOkDhoFFN2NuoZfNFA4
XzMs8kAPFXgvPkhsPlz62JlrzG4Borc/XQGLMH9KMH/seNFEgWBQ2jWvAkLWeBy/
p2wKI/b4ZdJWcX3bMl+G1GtiXTAKvy3QcplaJS8DezfeuqVFxPdTFT5m8XlzXN7A
ajfX4mJ778K87xc8hROoi009i3Pti2frs7qAgyAllAoG7qfg4UgX+nfDp/CdXB7U
wBI/bIXXOkjYDyRItUqIpybeYf/njCWQGkJnM4dnecfypeVXQvBC3oOt9P9T+JCW
SVkjFqeRYnPp+wFB8lqWdZDqtDFjDcaK37VV/JI2kBFRlp0nU4ob590tJUwWT1MZ
Z1sLG2rs12kbmQbyIZrU0w2OZ+teFd2Smxo6hvmPJhOEjMuDmErWr/LQRzsTdbNg
0cy/eS3jV6XwenWk+BwIwsz8UUDFbj1r5ZvIqXf4OIB98KXKRGxTEcAOxR9RYzPF
2d9P1GwI8MXu9tWq168iAZTkMOpRGfmrFR738ehBT2YCTnb7MHz9nOt9KqtajR+q
1VG8YfUKAMu1jOQOcJ0BN/zHmVAD+XKFoLHXnTk3BtvZ8UI7VsVSAx+cOJaZ5TqX
gZFxKz8Xes9EbQZDHMf6JP1P2VBasW0jXQaGesJ92tAoX+6VF4aZwn0WlmV+Cerx
bq8zlLZKL9xZiFsyQC2Ks+js6dSx4A6A7Y68SRby5svx0JdMS/HZ4sMugqi3TTTp
oKGevqKO8YhKelx6h1aFvn4tOSgtrqvKcLjMOjE6jtmwvJc9Cvt9vPSQC4yUBMm/
YWi+nTTBMTNHQFNQkD/me69ZQIUYcQ+zGi/lNJR35hdDacUdg/JBajwDVr5Rj/q5
dU/UpCi4NS7wBiYWMQKjJUN/Wg73QJ4z5HjYJbNUMO7YneMiP4yEJLHF140g0ljD
WXHZPO4wuEWN4UhC27Ls22e5CwkH06Ye7RCzaEe4P5QpN/6Gqk3cixylz7iBIk3H
d2p6XfDHZ2Cs6+ZoksyXnkbOxSfWrZfk1xKhCqGSRrZhfd2oTtYMyjunuJtNOCaF
q5uZJ67kmsC1uCj+pNX9KxZpAKtkeMtU7cw8LXsTP1P3fO7My9fCG7iVAhDe0S67
o1rn1doIvI8jDlyBU7FCdfA+aJACRSOk8E8FRjueguIPk17rjpLIWhY1Pj6he4Pb
cmMPxfc//d/jJhvRlWRKswsXGkq8F5YRLZJh3ATEJAYC1deX3dWpQ1msK5+K6GKU
IYztrRQ2s+LbrVOpt1xjclMq9Z23XmZ8pWw3tkx2u0oZmSmFMyJ5o2Ph1sxZ4g0y
Qn7HK7gOYty7yNumt2r6YZwK1P0BvutdQGE0L2fWBLDnWWPtY44Z7kndw4EiBdDM
Ee5j86EkNZtZeg0MwIc/302CmwxeeSt1W/U/2Rpr8UH6RjAIE9mmxmoiIyXHgHXN
7h+Mk1jYJ9u39TQkRseOIEoV+5Zrf/WF8r5/ob5HkXu0JME0hfIhHIcWp8qbjiOl
KSsiJICXEhCTf1RJf45NMdO3uNimKsC3HsC2mteFHJFihgQj6Y5q8NuyNymNH7z8
eii8uqyCFeFXAmSz178ZJjX0Vn98RfhM17/RN5LxY8FMyEf4XXoqvmwXkrJ5AfVy
A1WiKcq6hTmj4NwTuwwbYpEXOWXrRHcOP972YtHIFkopqEsuMd7RGRGq22yHl7l8
WLAfYsa3J/hET7n+0+ubR3z7oKj7DlUtEAnAadjJlXFjCIDVLvee6x4Et0SUFSgB
tg6d2Z4rYa3w1a6X6l/MyoyMSamAauOXA6Nnav7zYfTSKFXfuKwjN8n1fyjfcmB0
9EFzCbtCsenBmpW0XD7+NPlJRPqZrG57htVS14DfEB3v/rM6n+F99/CpWJ+qQWOb
d04Qf+FmeeRSsGppisV5cjj1xz6Kglp4aBMEjzi2w4UTrnJ0wLcFW+PvgTIcQqIi
Dy3hHe6XOykiMwHIiKATl8evnj35UKUKoFSATjevZDofo9+aX31vI7NU490PBMnr
7mw6KBqn3ziNCiFZwOQCxGcJGTRu4divhvZDDiAo6haWqG3TUZXWyVIoNzckvXpl
K3tDJIyJPkSZ13syCuEU7s2blR0Htqu+LSLT7eCZ42XRfYvr6I2+GkKaShFTtV/r
8Q2lQnIF2V4HNTuO0eoSIzKfTJtChCmD31qJBXbrd8ib7jgtB4px5jZf+V1zZjBA
qvzJtYGB8QO/8oOwXkJijSpTujo7aLbGK7FPEp/X/aZUl3XIny37zL4egLm25PFb
OH0dNDI49Fybc8jDgKh1FKt4XXKkACa3Nyxqr9Qq7LlQN0B3boVvz1EaB8BipB5A
5oIoUv2j+UEsbotq76y1Bmn5RCFzdp7eoyQcq84mZQH/h4BVOklrOgiOEAbmzcaS
xIsbP/KLvFAZg/KMY6QRg8Qvbj9TvlegEM6I7a1BcuYgLaaUN3P66EgBwx5tZ5Oy
b+xtFrG8xUgtjwHUhuOSsDEnTxGJMtT+EjXgyuQN0zjzqA3fwGx3hL42RyXtq+zl
4aOrZZQIWn6TvgpACMpHsQFoBFLxjomDFgTL0uH7+nFvzaHYQ3GNWWjwwk+O8ASq
tyiQTI71SrKPBj8NAl9qqkllyMRcQAcj15ywotMR6v8uhaanEcy3x+LbcG5sRlKJ
/4FfDf7upbed+wFFlgiiQQABSQprmCGleCuUv40nUjpf36acbTv+CFTKqwtNxW1g
QV5tfU2it6YHVL+AtlWR7Eh0SKO1p3KoJ3eg4684sqwk3VTkXOuZeL3Y9grM2dnC
NzYVxH9NqRCCQymZ7u2FBWesSOaMSxuNoxpyj/tokdxUBHhdpYNO9vY3aTEkzhDf
aaaNxjOcRec7VBGgKmVPq7OjW3Zy1482ZvaaVPGzu0CFCGS/l/su72o3V4vJL9jQ
rMZ8BcozLHNj4zL3yUx85DyAmrffp6+NcRJWwezLEIGjozIpq7cxcE9R3bEvZf4H
xKyMckZvVa2OSuWehjImSwbjrgvalapj7ygopiQn61u9FhABm6esAqXbrz5/KKqz
a6iraWK7Nslmtookaa9wWuFLUc02PiYHmxwgYHDPnhvI8+qvsjp//DQ0bz3wIcz2
yA4N9qNRZi3jlLw5c0p6Z/MKTAfX+HJ87LSWjaedPOroTH8vgM0nRpjCd6zLD1ic
asXkBwP7kGf6stoQDVRofRH/D4CraM3q/hmxH1mZacMnAmI1u4HpS+8zQJJjKGCB
sOTuwujErtaou1BAJddTJRGB1QewpxlqH4QuBtIcAEqabqMfVqKl5pLtHKCCzF7K
WehwgesGVC7YHJUMzyPkvHfv7EhuNp/qE9XI/thy/p29ByvjNFvDkaaVOxg41Y0m
wc7hF4zzQl5GKsq+xP+neaN/TsTmnFeaWf6hClXGxWONfh8XzaId4awWAxB8PICa
q2AiokeqxhdQkGFsK9KcRfU2XIui7trZ0EJGEm3wMog+fTpOcccKTIOXNhe5RNHX
PkQ94/KFj5LhOjeakdTPdcjPcrZddTGnXgIxMvvduOtLBKG57+OBY2qR9iPxsO1r
sF6cBcz05SrcxZS3/3KcH8Jw4y6ehn5OpfdxIZnM2xC5MIU6kYPABfdcPYZJ6swi
v50J32VKVQMN8g0GRR5Iip+nrNbNCI9RwCFDcDEhsxJFW1nfxsgjeqlWuK3/AXYG
UOmO3bSO+g7o94nmYSIqVpDZxl4KSr6p26SlcoWthvjDa60o8k4HG2wv6hs5FZdQ
+z6JkHsNRm5t/vdi+NS1UlMqJkuxeg3aNYU6PLPck+eCapwM6sRjdMFKoGLwFFgU
0pNSOMvCDKLLsV6246r8V7t+EHEIKwg4+p5YPb764bsHRHa4ohK/kzyZd59ABjPW
s1bbTuOeGWkqutsUZMxotBA5J/Wlvrcc7zQXUVeR3ydb2w4I9FkY2ljJ31maUMEt
0q0ZZXG8yuRMBLQbftjkv6pCDhO6yrFqIQFJsKdrkW/cM9OPne+aITBga2eZPUSU
7priatdavJejP9Bx5jwf+6q7hC4C6trAZjGjkitj3t6EFbXfK3ibwEgsyYhEv12x
6xoBlc0OAr78XA3gPScaZmnIrqPHMV4i/Y5O4lidn5PQmkqlj5wpVNXPuqFxg3cY
359VAWq2qSZ3zxmM7qmuq3qlVMwWjUquRueWwOnqgz7yZi/LG4aag5sHyb9egU9X
w1ZHsHKK8jqOpmFUExdvSXI54GEdXNy6q61ZOuuquXLz7uAMfhmpDE46z9Z9ZL+h
2Bl3u/R229VpPp0UGBVPwsBeFvSkjnMdxvji88RcT2SljoRvKi7MtLBc9sv2Fv1D
AGR3y6Cpv+gnBrP+L1FLUXZf/avpMfngUFo7K0LPJbWaRPTfnRLRALFwYcpX+Crb
eJu27gn2cn6E7yrCnqLCPg8SJXCF8/cSxha5u2Vk7momHK/dCc0kCEZyxkVWbo3D
S74mmrvcqjBLDIuveO0UUneadyvcnHjC/nmE8l7Sq+zW+P5ZiRGRdp6nXlsNwXb6
q/xothg1e3FJrd0KzvCGHlLSktYyA3r0s04QdDf7b9+Pi0CWwio8g1PJUvHMdFDX
ST9bjHT7nrBpslQLadkrDZWx6Maq5wRLXbgpWmyTa5SGa1Ti7dZB1D1MapKMrXox
o6G/Wj4d4XOqGofILgCHGu966kc3yLChvd6Jsqlx8Izvh+wRzh+rnxRHDtN8Vz0E
+U1LgMrY2bow/0YfAfYoVoD+TCJvqAjgsRajl/varWwQbutpTyD/p4BqOzTO7MTC
kw27KYT06UWHXIG46yy6Puo9OYq5ZS1kM1nFjuIrmvxLxknShDviV85JD3rWy0cK
8gZEhcgok94LpF3f0ch43sOuLaV4NsTRQkwCjB8anu4BjFzlFbNDxAipaENd247m
zsjbr+QxjsqcnHRilhRleIBKl+JEDg9oJ9I4Syu959/DGtxn0fd9uFs1PUECMeGo
na2+dl+dJbsd6etbgBH/OmPugvpCT1xo8UKDp0nYDMznIe7LON2ZM6XjSxpJxn7T
ZyK9tnMseSBBG+itPJt6MGAj1ycPhMJVPnEy1XRQa6WEyhg/0PsGORaLlmmkTQDU
dCb5PXZufw8VhGyaADmeRNLXRs1smtZaT7Unyzzjts52bm3XF8uIOXempw0wigqW
Vd3sQNbPvP2WhSKY8dNn9jQtfUIQDcfVJ7UZom8J5t3f9ELHcHA13WITsRH2dj/B
pBiUh+SrHGOS37TQ8Tei4J2hK8ccIU7r6b3o/PEWWfDKwsQn+kCAYCJW4n81ACOA
xxrFMCi3NoKL6T4PH3BZ1Yw2f0JBpe5H1h3U/uPfKWl8nhgwT9x2KHflq2ymCo0e
ExRVwpK1hYRXc4l3SKMPYDlOs6A+mRujbz5bLtM04iCLK5abMMToCkQWOUojXVdh
xgnHacVbQoIywDEjDt413L0uVcN1iSYFwTLcBe7eQZ44kySYk7xdhhEkt8rGzO+m
5QRIl2flwcBlgyZk+2PXLKW682fg35vWgd0EoRqPrj7cwrDDXMD5YPUItOCkFLvo
e92gAN3vInhVUSs5bawfiYgdFJUua1HVGZNMv81hBVmEAYoNLzg9AQiEmFCGI5Ut
lVKp3Mr+GvWtwRqlt98GCPfI9kBLx4tGzIVrkWMUS6UKpiUrtQiw7c8WUJpDfMZb
XNzuZqv9d1RruZhhRKh8VvrIvNxpG83wgoaIMr2gfNrk91/xT+l3uOqEAsWHTG/B
NswX3PXb6gfc0SuH0fxqU7EVgEAnRgeoZI19a/3qnJqQ4mgg+cICU+g6aKURx8AS
HZ43x0E6LF0bpy75BuWjZqVJ923EdA3ya2ma8IXxuw52IN7FY5eZbz8yRtmMdPD+
M6ARd/hafjUG/dKTu2DfF5yV+dy6tORcS0JS58RRBrhIXktvqrvRTruLMGI5PjNY
cdUZdqgqQteaqxx88sUrm7Q5T+ecjA6upLZW7NMG2/RvybSXhCJ5b9fnUsh6Be1O
HNUuaY1WOeamLMAzheygDRsASejauM4kwjlcdAIv7WMvAQryZ8/LGHcmZZMYEPBR
waI4v20eh62wCphvEda50+ZaPr/UklI36wXAi3a4asELQHdVsFfpfRtlahjrspSE
PyorpXx96HkKJy3e/6Qj3YIPxHifc+OMLzAi0h/X7pQmi+QMoPQNNxG+bPXofpDT
/ujwvV668jnheFGiEp6GbEsGN6xpOTUj6S9iSHRy6IXV5WhS+QWUKlQa1i69Qcg/
HEOJ/UFnDYz3CqdpxeLLFW/fuarJ4+qLoJc8+219WBgW3TpZAb9NpC8cGqiOuIrn
OMrDSO59GLe/ZJtinN6V/X5g85RBrw1oIjGZYbQAd9khxqls/0nRYjrIcgbbGz8i
T7NsgyJJ0CXbvkHaW2bkCx1wpcNM+ood0cbpkEPEwUViDUk1bGyBwf3spgIy6JkT
xmtmr9mD097uy1a2+mVgVuxXpeQEBfWhtK0HMUIhe3PHw2pO8mpvxDmOc9Ez8PkW
+OzTxujk8KXpX27PkszCCoS71d25mPzGKv7CJ75nf/Le00zgCHPjo+y16ulq+man
xVgSNlDIRLkgSPx6uakSncq987/iMClifj9eY0wKJaifAGDuYIBicTFK23vaUCH4
cqxY5SFfy/dICCy+WAsljQTPZHzSIMoLHbjQZB2znfXedFfbnDUmrn5XA/bV7pji
1c258+nmnxxpQ88QKjojp1JqMT+pUwXnpdRQjjulgoN/y98Ch2iJDSGpUqUwHZ80
DTY2YXnbBdOneTDiEr7M0dQ8lwgYdUppPA28o5ErfFxcDeBwzEcTR79nj4MbtRyv
Ri+IGiwJBOx4vjPtx3V0wdWGdRs5PswUHCjohwKlLNyM5LYZDrZ/imcTYcnWnt0i
JfV/iWGMXuDjwtYbIHGFSF6qQHI34tBTl0pZrK82hZIwb29mZmxK6Ep28IV9Yk4t
sKrUvRjsKlgERcTR8py458BE5D9CvvcREElM8gId+AVDU88cYUTpsfn9Jl9CfdEI
UO7JC+oEneEcP2hKoLqs+DzUAzYVVFdBued8oS0Uj2vWkd6w0TK6gacKwoP8hyU0
clLxDE7Bk7RqLICn5FbyCPE2DrI08sfLjYKWpqFFq4PtmFtFJ9wmjVSB8O1KiY5n
/4gnO6uzHtbXLk6I++FiXkLYvljAqqTnftsNKpiHr1tFFQtRKYmN1xXbgpk3ThKB
XzAckXUWIzscrDjyDxfcq/f5OohJs/llk8cQzgtQyMTMkLXTFWBVY6K146Vx0pxC
MatTyxe6S19/pUJL5AAstQ08oi0o7TOngg2ZYBUEXSQ4j3+aj/amR1osDXuGVNkV
B7S4NGJ+f/kIMWgPVCt73yQyWAM6x1nNLcCyUmdaajfm9p1UDjRdUD0dtFcRagyu
LiXhWNQgDFolI37PQ/7T4KVu+BdW5aWmqR82QB6XfXS/epl3Dt91YWC0SJYroOnk
XbIBIMGYjcfk1BXwWiN7hmvUvnMPxA+BASMlKlgE/850dP84BagyKF36rCYgAQZU
wTCCkPWF4go0RH/FUh5kCZv05bUB+WDTOQrhep9Bep/tSYKvrdmkSNM4VtDtSKIK
CboR7znpqz8rOksjZg/j4JnSjAl4L3uWfvAMxbvDXnia1pVkA3pfySeqbMRi8ULe
cPMydLwwYHLpceMrKG++bEXAMQxXwsKPocCkV1yL+m+qL3im3TPXarefViYu/g+7
1cw6Va90ZytjtF3K2YyS/lm50yk8WhtSErSMvs022fvSm9P+tW3slGufu7zYBiMk
dp6Oc3GoiD17J6YhElrdEDGQ/T0hz7WuEFFp29eI2t1Wd7De8tPx/hdsij2BJDk5
bOPvz+AUwDO3+Gw2Qz1yf6Bq1GaOzdBLS2flIrUY47LynvERRID1loW/UVUCdUlD
H8KMU8VpKI8Us03D4nX5qgt3Sh3UhR1RA27njZ1mWLyQNeyD/K2Mx07QCbMGxQUv
ItbbSFkm2MY+NoIp82eeqs5+vanjMaE+o5frevtNhH7lXp2WYOk+DhHMewdV/P3G
r83HZNUbqaDgfi2VonN8XLa0A7jQQMe0Mz+CnydxyEBzeNfpDZiMuRsnNLj1Nt0s
u9HtsjHZsINAVE1jy+Q+Pn24nvOSl25OVLumQH0i3vcw77dYrrNQsJqqvHBE67Hj
MJNfHIMpMNDjDNJGbev4Fa/wVVNahAs8wftbpp8GuhTxomdFnoSd+1w4JmlntMNm
5vazWUKz+9eJabN2EB2gJH9Oe2JW2vDVn7wx8A2WBhDUkwrN+k/m+SZLDNP9jXJE
9kVG6pE45UoA6ZW+zrWLW882RHOf3TSa5O4/tFFOaa3gahZi8KnrSfXfy9f/vphm
uudDqyttVCPUNrWRNDqTULW8uoi1OxqGGuf5d2LPTjMyqg8FE5IBHMl20rzOtcSZ
P1/stHA8kW+hklEBB05kHLjFD5ZHu2Stj/zCwGEZmTLgtWUgWdxYR9DJpvFqbAlU
zaXA56qGKutLFdFsTIDqE1khbQ497vhtKDGFl0bKM1SVt+U0mZiXmngAxSxLilGN
TDDoNq6m4Wk5jom7ujOxr6uhHX2fmtbEyjPMVV8p4Cu1E6OyV3PRP/TxD3zSQwT/
L0rpePEatU8mLGaHI6udt1lRIJoQMq09rDvw0wXxxTilcoZiONZKy6hkcNLK+bCG
cvzottdlE6RcdBFRQ1KPEQYoDJ5zEiJWd/ELy+ovb3u7YJB53aFVpQqpzTi41rs4
phZOu0lxoxA575OoAR9NbvW+luL3Ng4uhghRohy42fSFRRgcO3VoseNWdHiFgr/F
YaMWcZW6+X0xCtM8ATYX4CyUOK268IlGorwvLID4JCO6aE5vYfUS/k1cEgUHYgFJ
KP9SMRCXzEsGxyLvKBdkz/rXpVf9aFTaFblS8wjHJvfA20srH2Pl769gsx0WmzTg
iYfz8yxazrzTwuWCnzquXfA2qGe4aLRNBZgczn858T2lcliSEp/R9x7v2pJsLRUo
XL3iWMMxMb2rcbHz5GQDkd5Q2kzwFLOya3nkSZr0oIkqlZZsNTPpS6/GeUpwSivS
xbsNnqKlgTrWM/gFLpxJBg2JC5xeQi7dv6AbabJbxUZ+u90WetP7e5NobvugEykU
WEvPW14Zzm6SpoZrUgzbN3HI9P4+QFJsaMIOUYBjn0YT47tegcWljvbtohAUN8TC
PyiMtqkVX9/+aPwJjIn6/NhGtf6sVV342T/VG5zco7UItYv5NBXvA5Uac3JpzeFK
QNIVCNM6D/OmzJd3ZfTbYfTCA6dIUJk0CsHu4nAPpXWB7/Tn0MoQYlTdqrJCnIEG
Pf2VyRZhgW2BnulRPSIoIHgsR/+qt+7vR+KQhDS1JgQvZLOpO2OU/0+6ZsbKEsUr
hML5DdSPfm3nT5YxnUg56JcvhNXKaQ3PcnirxgLXARtq+Dq1WR84YvKhKWklryaL
ZuXtaMB3foSL2cw8gsO5nTxsGzQ2MvB+dEmpBbWbuaxWkbiC8lIBxI/DXtK9kXQd
0RSBE+8afoSAEXozZXuJIBjkXVqlGMafjC+Q7GWHEWsilBzCi3LkWRFmmdqDHp5W
ZeIBwNw5ev4E54Kj2FGiWgk30KieiiCe9tYgNutZ1JzQdRqR5CV9AeV68rnSpneJ
6EqsAtxPjuC75SP0aaoS5T8KBFfjiX9QmHDLygfrFws6kcGBMmJNvBivUvQibuD5
lmyNPoVIjgI7vIyxxkpNEjR1G2DHfzNXr9Q+JbbjQd65DpVb++NMAoeam0tsf5Ih
t8Sx0q9kwNRAHMMstF0wOmX9ZLayhl385no7BnOJIQ2UJfjvhQaw8CRAe9dLRNxd
ZTtIsGfaiicw4uWDbhp6VxJoorvoVJDd1aeefJ09b8kY4vNGESmofYVZt1YpH352
PMWGaullQ851YYNKUwft4p/YsEyxvM6VBOxkZV61CKYhHNvSmqoxJzVAPvD2ZLeZ
JDL6KIRe8+l3in/UNQLVdXYYa4ojJG5rd2sw2WFUDTD00WckBctp6MqTSXptqV85
dle986+sPM8wTyP89TYJKcd5QbnFRYOmuRSlKvRcqUzjBENgxeVd3WLyykWtL4Gs
nd9z8FBaNHA1gvDtLY1k11/5uyhqGlllzpS/BW4SOhdo2MaTavxy4yEi6nc5qElH
GTUv+ft5ntPohX3HeNazb09OB0/M1kSSIV58gzqPuQjuJ1Jhc4w6QbUk4IQW98ac
2JTj+teOHz7DayQm9Jf+5lbi8mp5v7nZK1tIVNwfRI7WiZAfGe75hz9T171RbvA3
RvjbqH+b7WsBzHtV65+ZvrUAKQdaVVBpq8q++AZs7HPbnxIL8aJ7Tep1RL/veXDq
tZ0p69yKcP6X6XgAtYNqbopA6GkfwNSr+8et//+Lu3bCqvWNtB/qZ1V/Ddt47x2d
6Wt67a1c0Nkj4wPg4BtuWO+JxV2Jb8XLnKEfqS0PZqoEky64QgNU7t7dYK9XCtl6
b9gi+ZmhlqszhD7aFlydz8K7dxSai5QgnyGPG6qzGSxmR5rtl/56LN2NM/ApZLkm
Z12CRMntNEJHWH8P/VMDxOYW8W5Kp2eeJoTBspxDzSyoyu9Wn0pfZuJiobUEWad3
29ypDTnz80oOEQ2u3SbiY2H0voHajWy2yd1BRLO53uDAyljPmbt2Li6sPiBgfQo4
o08jJaX1P4zPhKs4izyvNnrWM+IsgFKKUkbu9qHJKqhmXzolIzKeU2an+y7h5Ymv
I2kKD1dFj8wLU2RWe2onhFg6naNsFTSpqS+YuDeZi+ngKidO5/A5a/sUFkWULm3i
LgyIjmZsm/07CpPhduXKHOy+RzhujYfztWc2GbLrgxyTEDg/7VS4iEJmc4qK103M
Gj/8aeF4V41fxFC+OzXVzWy2jVLR4R7WsbrEXbKNKPqmtu5MbayMCWv+aQB9X0K+
Cbx9MWcFx5ya7WPdzssQ44Bvs6wFEpz3YWD38GgSa/eSnpnFETbirVna5kQrWy1P
J0200HlwSxCz3SUTZqTtVaza2sE83aAeNPUTXPMsC4Lctp3UmrsdQUAo7AYRCdXL
97596P66AOC1lSnlHYGfi+LiBaEHm7b1V7b7s/zgjvw99W3AlC0qW+9q1V3f7Mze
JbKaQC+HnN7yUhRTPTcw3K0wnjXHSBEWJkrJOVoaR+RfP9mkO0FI4EmclOvp2JNf
7Jx/eD0OG8NrQF4+12Z2GL/AUCXi72SR9cUVEIVef9fDVuL4mA0GP1NIAJ0qE2EA
VYyGJL+cPBCagNXTNcmJDoBNDlrjKQWEwX6/3uK4SUapp013ihbMgBTyZbpHMh2p
CjVEOf3+mQgW+X5khrLEhdlPK4gEWx3G6pXNTvpVg8gHE6RzjMppZZsFaq7vgt2Y
y033/EIERXucGZvBBEuh6e+FoNO/KGyZnCXhQh140IJ9AcYubyRJPDrqe7Ncv5ZL
grANgpfpgSl1iHHEGa6Styhub+sO0vyhH5KfNnKviurobGESIRk14kqQKOyx4cWW
1eoRoPv27t6gQZrQM/ojG0InsQSdERs0JahyDWhLxVj4qM3v6gRpFlxCkzsQKzeb
MMaIuCSmE3JqtVh9qmE7F5ZzHW2DWyOaUZGf2yQMKlqna+UPVo35NYAemDTrKF9x
2idBFgb9+qmI6kjQ8NvWihZZBmh6x4dlce17274OT/1IpBaOzrmTPDa2cvXDkiXl
o9PDCYF4QCXlSXCsyEQwp9VDM39NSCVVytLW/HfxlBIyO2hx0AtTMzHwYDJBcLc3
DHKuNyYGIINsQFwEbmij7R7dOUzUV0JRodQsgxoJSqXaP3dXB7LK6E8dNqNqkE5N
/KKjUjFfCwXV0J946iBmEojS4TQb3iLqeY7h0pT9C1u2Jx2OTpYxVQYp793kCLCV
r/2qdXbIt+xy5IRIWhoRmqGqOkMUgBKdg3qCRo3fntVP3rE2PfsrVFCaTx1szBWA
4ibzdS/AEsPubMhnu6BKiDRmTtcGcsqCuRydiV6/Xu4pQHB6MACSB904R+dU0iBr
jabWtLrq2b37ShfIeLzI2E/xNUstBTojDN1SrwpylOuVrMG17UG6jMSxTt0nS2xD
XY8tp7oRudpmgMlnCN5CeVN98MHD2Y+ARGTZ4V1JpLrQ4cg2FG4Q8GLMHqCzZTJg
lwK+rxpKrWG4DtR5AwUTSfcpNfjxjAQifzDktYy7/jqu1JdNMn3tEe7kP/x1W23Z
Y7FNdPhgLAi5vq9h4uhU/nHNyoopkgZHG7N7btXsKMJGsfTw6pi2eSnlGVP04tXw
j3T8nzePP8lmqllsfleOyF+l0leJGf5pmy/yQCW5wJTk7RYU48Fuz6/Yzi8ytp9r
bjriwbxdclIy8BMOKpSTnkcDLy4dCMXsVKZh2ZnK3KeAQdh/MbEVSXXveiew7F01
B20q+p+YEfo1GC1Vk17g6nHGFBXXqEG+qH/wZDZmxouJcMLDzvX37FObbLFlwIQ5
RscyTr1SKbyGxSpxyx6E9Ln9+4QwOKd7cQSsjC92Ewadc8XQ3qHs0A2EP7eYVvE4
G99x+OfJReYNP4tFc+G5qpQOLfKhBjC3gFUhp4L84i/kYK4C/HjyJctB81u82722
yhIjuYFP1zxXNWe+dl6rlXQDiS6RA7HNattJiYKQb80WCNjgj2YSnNuazDuFmjV6
ToAahWi+Ku/wBy0zPZ5A+9X3OtmBIoV+CIzufpNU+AHIwgJKz4uv6VzqtS/r7Gih
ZJNHXlCOj0HGhA/6iCAvCspjihxkZFoa1h6HqDesBiZ3jOWa7r4vEul9JxLOy2gl
hU4a8RaKZ6AUzwdy3prN0HMXavEPLowzWKHvsBdeb5Jnhaliu0ymmWqawZqFlxEs
fPYADNkspeQv8H+CUNdO8/M7/T6C5q2cBYZ7752zplsSECspgVtorSLyPXDzBrwA
YC0F3bMMpZVX9U1msSYKLZmcsvi1NnYqJUkyEOWdRj6raFRAWjmYOH7fnPS/lnlE
oY7IX6Ddac7XpLlGS9TpE+a7JdxyEs6ZtyGJdqjNZAZ0t+ldRHxNA/1OkcFUOzCb
xHMSYhXhP7xhPiXb55ecd1yQZZioHT30BhQkvje+etbjig1hCCNvJJTKDdSLwNSC
8UgHUAtgxZIn/ZybAm9ruGcCN8XsLdO9RNy7M6zi5S2ZzaI9CDSDhBuksS0gl4AW
SWZEBXui5ca1ZmsmaXtZz46NUdxwHDwY78HLzXmOi4VsCNZxy1e+h4+AazznPNKo
LVO6rvrAZyrec9BfA2yIIoxlcBeHBoobs1kSbiqU5eo/5ObQk5HqbxEK5sL7Cukm
XgFbgEOza+RzRi24peOs3WRgVqb7zASPEvoOQjXrIXVJMFgFnTK0f1R9fElDD2B3
2BhxkchlfhxvhC66pDaAB3TOhrsWbGjQzQAYte/5+XO16uuakB4o/klMTQQNoBf7
MCp834TptKCjfj4fqt0lgyXCEfVsngM8v9WWjP6ZXSteDYD3yyGeRC+yCcHGWk+9
+sDW4vVcFKpbkKatSrtYOYoKpdthA3LoNoxs2MHYLuspC6GhNoMTgv0KU0qfDjSU
31bLbS6hNRquzWA/+Wd61HppN5pIViasguzV5LmkE3j9N/PstoiHBmUgFSldWegz
/M0fW1Rx0moy4PwIbNmh57eaNasVa/l0I3F+qY+GqRyGzsIMHUMvYKXgphouF2Dh
ltS0htxAdRoSh00RvCXjq4TBhYtUC5DmxINcvig70grunUAsZYpAPn+LG6+yZ7Yo
IWrt0UikywTlB2Cs84drEZ8hHZjYZWzCurF17Ss/l+sUhGcWOp9HyM1MgLGASe22
50iBc7DlCvHtgv/A3lW2hA2WJf+laj/lGop8VZq7foOILIqG9dJe7NgTCrQjDofL
mL+sel7/LH4OLSvi698qerJmNYRYCV9k+RxlCKW5EU6kmNR2e3af9gI5zTaTxBIL
fnQTXLOEPxgO8b2qAeHyLpR12uxN/eb7UIN+zpQb9AWQbuhFW/J+EkXr7nhOg48M
sYPok27IqoapVL3OHK9g89iqmcN8ElOWJdVSmN+siLkQ4GlNvLU0vNySah8xNMQs
pP5hZ1y0d1KS2dm+lcdy3hWewtBX4CdymO1pCNnxRnFmCOOixoAS6PXGVLyAvZx/
CP1HQKhozPORcjgG9cQri+nIczf5hV4oTfk4Voq6R7mVZL7cDuNrT0DCkjwHURhw
uI0pelScZpcC7aiCdiuyDOx/S3BMl7IpWs/gUSyqRIM17PTPUT3QsUJmx1JD9s3T
lBfVni53Ve+KvFeDCNO3c/z8LINGYcdRvdvAL101FUJeEwV+w8q9VPFqc4dIWWU2
svT1LQhA3HszM2Yb2FIkrO9OjvKnaZd4OuQL556IUiSxOveWUqeQGjA0hVj+SRUQ
5ioZi+C8QwbbE6u9l+jX64Grtdxa70pLYsrIFmjOQP0zBu7KUTHNfro1LWdKv5RK
QC3EKEBh8GiZM04rArgWXIh9Flp6YuO9HVkuyGN2ofo0OxNQoaM6WDmi/TZgVElC
jVgCaqClvT65uI9DNxFAVnog3aA1CCo8IfE7qssuOkUzaNE+KsjgSRX3QwLuDyKf
Uz0GHh65zz3uHBb2oP7NAPsneyZv9HDJ/wXS9gI5VMEJpCJFKTMTEC52nvwwOvKL
N7ZTCC55P1SxZ8ccnXGeq2LH4PwtamUZw4h6EETluXTnZ8vevGkkQ/WPjL74JAwY
90xsMNaFa6Jf3LgtmeIfAjwbXkTCVlARacobVmINcnYg2pehBjoR7y65Yvr1BvcR
YqXNo/A0utmo8R2THpyZj3gHWMwR09gP19baHxcchfHwinenXan66YiKety803PX
1NTnrx1MmMJRQZigZfYgOYUZbrwGaTlwgtEjnNsHfd/4PF2K1mIgOTUCoJL1cwaT
UIWczJQMw7OFZIyijD7mDSH7PRPPxl3eSSrmvt08H4JSsmOOfsvyrC7kdk1zWNNn
3jj/fCg2Jfdj56jexJqOBvewVCUYb56vJm4m4xNFYlmph6IFJu03HjlIfo27+L5p
M9I1A1KlXPzk4uEe4qQia4ICL1lBOhHmQkngc0s/Zt5g/GLBirFaLWk8d2+AvuGC
kmrd5H2uERx/6mvrpuvQydXc+sbD13lmaz0CveeuhXSLfuFI7NPJgXt1x84GYvff
/NkkawHFL9yRVeEDmZMXNow3fFBRVsAjBH15d47fpvWydilVFRGbSMGRIs2VvjLb
Tpaq7ML+XVgW87eR074B72ErJdl2IO+53iuKE148YDuWKIVypHg2bJ80ArVmJSXc
6fcSONmfIrkgxQcdNGrl6UnAzP31bs8uviAV47GhJA4wXNK+PQgLHcoLb+m8m4B2
LUuBsmSttIu3xg3jIGb7fhebNY6RpeQ4uNEQkK8UOwvIRy1GhuoTO+BIW3YTLwy9
2UwUcK1061yIjfKOaBdAqg9pBKUl9lfVucCSxXUMJYQx+u+YEoJe6KvzQKA2MLHq
SoyyK5/73VGp+JnYVC32GU11rawomz7ZfWtNecsqeiUj7sRoOtRUDLk40YlT3jZq
gXamb059tma/NCza4wzaK2M46b1vq30W4V2JD9qMQvxhpocluVjw7zFF2+igRPUU
cduvQUJKvOwA4cCYw4OzO7xiwTzZ+xHQ573f5eVtlsbkgROQM0bV66YCmUq7pgQf
Zb3T/WjLVu1FMXBjKBF9+1FvHUZd5KV+VAASnEZL5YgLz8wWn7xD5G0SDAHCPQNG
EIV7sKhT1ZFax0WNxXZBvdWIW9bfwY7Z34fF/HjXfWBCLtNKfyELsSN5qwduZXBj
izZQ9t3wJDLV4spH0sOaw5vyxHo5UFScA1MAZ5QLc+IE//ZMi5pLGhn2kIi79tRe
8P/mbvN70q0OGZ2cXRsqC/Mqvv6c+4SEGFC8v47/XaA3Np0BKKqAYjB5Ly0IKV/o
5gP3nr07ji2T5wPWSypBtp+0dND9D0TKc+aiXtbWNqQbGqrXzwlO7k+G6qnmUtVx
bYe9O6CRZHCh6T2YQ/89Ckpazz16tCxMYhLPxnDG93j3AET/+UviFJETlNsznYEQ
gbSFVoMYmFjbVo3Igqm5UIQlSaG1VhxEifGdhjhGU9F1P3PfcO575q4/T+4xLP/v
gXi+qKOfkmEav1dlmcRXKwn1tt17F6rRUjtVAAbEWBLf9GkC+s1qYuzHfZSTTUgE
JUJ/hNgt6wHPrm9MX8QZp1Wgmg29H++jE+S6drtvRtVfyqvuHKX+Hanxnb7hzTMB
2YYHlpNfNZ1UwDafcc0opIFFL5mxK+pHkLKQkklNkoPCI6QfTcsVWzOiAZh4eAH2
IwzRqyy1+WHKQnrYMkn/uZZNTh1NCiIoM88TwD4dmPPuLal/toT5sReGARR3XVBu
fY9xlgrgpuxPWVbyoMEatIDYAEewZW5GUdQHbHBrxrO7Wn1FXXFGan7EVcufKDac
6KxleYbX5Mk8hnmPodE9jIVZrU4vU0XyW8UVP1QCAPa6uyjunK6PYYtSUOqzy9MC
4kB146Fmbc47zhc/OSCVyLMEjmZGg/CYkYO8bCD/xlVVN0uXOa5n8VdWdkpEH07m
KWR5Hv94x6TcWoXly0XEkp+4j37av3+lvJWmPXvIV3IzY/P1ZfWm/jCK7oXrGu7N
ElKQXMjSHGeSMMgS+erv0wXYjBepz6RO4vWFE50WQ1AmSVdcwHX0YW4OPoXvoB/d
3U8B62wKr9kUElB1MA1i6rBVI5LCJRHqBCMFkuFkGJznVc9sO3yd22LUMMZyTohH
HMktOoH/dmOtwx8gkxOCZGL36XdSTTKzHniefOH919Ou0aocvaS+acALrfKZL9od
yTuah2YeLmCN3sYKBaf8uGMG3VI2oWPSmXAmPsfJqDWZkS+IMeA3O+0NaYnY+5ej
zsxGMKiDXTSZjVo/XkwpzyY+uqv9Quynixwh4mBSEohvf/wBuFceK+E2mrbWEZ/J
yoxkQWGQQjUdB+ISTj2IivGpgPEhOnyyFDEgHzt2H9r5JLRwYRVOBG9Q+mljzhma
/XOM8aA/s1VyHOKZJtiEyo5fVBoEj366+jZKJQ0azf+nuv5ClSc1/6La7CSfGoUO
WPrNj90IX/BBMVT48QBmciNiVw8nYQMExHZvO9oBIo0Hpg3J5staf3m73zoiS8mu
qmUi+9volZqdRTXrOo1RAfMmSrQsf2xf49ALWZNx68fEarBntP3qP1Bcpx+/zxXB
`protect END_PROTECTED
