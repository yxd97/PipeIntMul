`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
diCpdb1nLXyRBazBbY+JlkaU+Xp5D6lP8W7pYCBTIGORuh8sYp/83/QcovESzySd
8e0Jrhr4ePW5Ur5uEFHPuP40ylwggv6NMUzWgSNZxCA0n5yLLVXXMUMl/IV4HGCK
vSm7kkZYJ0s6RnRn6JdPjV9yBEKzyiUKEQaXIoRxfJBy4ye4+qvozMh+KZZgRqmM
OjzU76zwpKGBEYqzrX5IhuwVmsaGyCISY8xBBjS2odAIdpqpuDU2CkbuX53BDKEm
EnzuDOuRyspM9SvKqUVKnp6tP6quw6LFfvnXa+CuF+bKQ8XbctMDRkdJlySDDG4T
7Ul8/TNLwvh34ASHHWC67ZiFlbv5riPyChNTTEyGlyBtoSLT4dTR6mzh9TirhmkZ
ifBGuqM2W6D6RJnPc8K+BXhLBOjNrnWyd+QiN/7rhBZpxIAEO4WJODaURmuirmsZ
Jpx9Uhk0Ml2D67+wN9+1LH3zrC61uQoMF63l89SM/gugKZupDLBn60Gfl2riZCGN
z+wJgLgE337/s3/cEppHiPUZCTg33mlo2ddeF63EvyxLDd/ZkmVTHgoHtcAYREgk
TefGcfVCTwV7XbBUMJzX+HzTIT32qXquaBZnMNLxzAo=
`protect END_PROTECTED
