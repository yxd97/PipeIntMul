`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RTsXNLykPNj5IsElOPfpa9vKfGEsaW/rBSOA6FuftGt3x19nPUifCVyJwFnxwqDO
ZY1rqYEPnKUdYSPQ0QNDxEL0x5Olw6g1obJ/RE6TBTjHvSVKZww/UiRqqg42X02w
JJ4jSJE4fmfIg90IbrH+5lHk4Nx7JoRUo2YXRMZtMyjzez/zNVh6smytJx8ejI0g
ZHTDIY2RFC6LIRxc+P4qJT05DAJ8EZjJoByK65o+k8fMi0AVVTsdbVcwwYdLGdkP
Iw/fHiXCWb1nZiei51+sRdNSTqGbNmI/IIYalFvhlDA7oKyYLagutPxIkV0O+yXJ
CiCHsNtm3MJk/9iwMF9um0KSDlB6v5UFb3POGekFbv3XTMXBlpCNfnfwGlD0hpAb
YeEU+EtFFq/kXuslm48qJep06raGuvfGnAMoy2dEbq0Ic0BTWWwbMXwzoZN/1vpo
4eUzbhwiVN0f8tXNV9DkkcUqZp7gTxlAs32rnIlNDUEkaxrjW5Wm4VtEUCbBc+nZ
5ppusmzvErDpmDjcrs2QuIRsS/Pj25ODfCv3SDmKMw7k8tFqFgj/60U8zc3kb7tv
Nv+Yk/AgBbDR1eUY/YhNm1S+fptjzf9Rivy4PxpwY581WR/xqFJRuFWmLlBP7C6r
A7l6xvhnPBasuY8Rog+WOFPAhVC0HSKt/IZjI+V3IigE9Mb8RbRInNl/DpBhZtpO
MI6W/d0N5iyaQGV+lP/MMB2GwHdMM6mXwr4OASZFt0Jqw4xAafo3laRgR9KWI6l6
n2Ex8HguL4XCn7by6BB+XQyfWGL7sF/aXRnesd8C9Xz1CJsxb/ry7KDjHGO9bWB8
qcsJ6P4rsIMH29GC2nYehB9uMtRsSCjUITzcKXMWHDWR5rtXdIZkquZCO1tFFFsP
l3cGckvbOsdZSgCWwASrtQNDhfh+aTap3BJyZVOj0et80YWGW2ew/1w0JZNIp8ir
wT8hinTucYY0/EraGJEhcxXgF2rUTj4SmI7qAL9JYQDv52cM/xacG58W29A3ZdHv
a+Hj7yOmB8woEHYtyup1rfiAxq1/3t0VKqubMnWMlO1bjtme38kgPUBjs4olkw3y
dFBd/IynDQk1m4pzwNszyrPGwKZ7hgA2mGkj7scEq+W7T1N5rMup9TqJFrSiu2S8
C67zvgRfyFnvEYe1n0BAXu1+K3JQorDOFbYMSdybV0HtwJPX0NrD5/VfKz6XtoIe
91cXn9WTOujl3pKeWklRkrcMS5ChrKGX4t23VYHp7PgzPHK3zXuIsSAXjckl2tLR
xU8jCjEe24qtTmK45DmVlzNgYrkW8a8jJoxOjgBZR6r9iuquh78W0N/fj8Lj/M/K
sesD6zOwJPuujXWoSsT7h0tC95UwDKAwFMFS2feuCT7cIME0pGL61VDZX3Y6ChVt
DI8K8irEp1hDl55wi4KReqC0RdnoS3qWIkS3EazGl/raRyWA60YweJ01ZWVbF+IN
ZDBKVRVKTymtPdOrvuWnNYHuDl5ynhtSUL+snB6NBmeml3luq1hRl1SG1f6XcG0X
Z2EodmCoSDvhwFwN2knc+uLemHMeP6GwKe/hVlwTQTZTQbcTIuZ9RKh7oCfHcQLg
ExWRr9No8pg6H4+9r89w0gzo7GWuXdt/L6TZ0jq19Qz2my11a8m2TUfr+hSsajNC
ufEGGkvoiUazRY5BVVej2munJa8XSjn8FuxaXjMo7VgSQgny9sM6oqO0RUKbGynL
Is1Our0CPYkEUiEXuC8lBzgxMm60eVy79HKm1UbuiQQZkotY89auB/QiiW4RA+6s
GuyQjIOwIWcErevpDXeuvGNCEZc1J9dAMxST9eenXQ6/rrx26uOd65T9pnVMbkdK
dpMfob274eblLXA8ZzCVFsPoR+MfvAgate+BzSY67oVS2lpnDlvsASzUKjDP7gQF
VPgbUBDgsrXq8zgMH/BXmzuMeykgQA41qe6P3H1stHhf/f+qV06bBaMs25AyY6li
u664U+Dfqm2mWbmR7DWEv+ZSAnulklJgq/pHtrhvrNZJoJLE2LLh37Zo7k1pRSWk
fixuT73Lvq1QUW3dWFSloZ/M23nVbsQpIbHW6MKkJeFkHuoWxe/TRJkb+kNmgIQx
BG/vTpXQkDvO2eGzjHdDBEzMjAtZGKJYvPn8iMuRQPsdkU3YNA67PvuzjVN9OhwS
w0xp1TK1f+m9sG2sEr/rEkb3zDmXco+tVed9Pg6XRmM11pnpBtylP/oXNIFBfyC/
e7fhh802bIWE1hEFEZe6m4X+gTswBSSreiL3DZqxVPBCMrN2iLfKk0Kz1XSz2v/5
QJd6HKh1YdhvpOciHr5eDcXQ+FLk9DzP+LEB9HrU2iACrU9Wj7maJpWJcfzN40de
Q/Odt8wXjjvHkJjsJJnIxF+dkaXuk/CTU7CsaGrh5DSmD2XJ7PmOA64F8KgwHOgj
yocbBq6IILUH5FIUgDzIyx1ZrHVDdL4hEsjQkHshhgQDsuRKRkgDz2hQ6cUoLp2s
vgeGf2JUBJTbGfRQAaGz/LvhNd/C2s1lad/dp9Fs0qzFpHIpPPjiWZH7Tq8WFfet
EKH+5linJ5AUBmnnAEfYK/ucUlYNAfEkGi9fe84ueW1ysfQGGt4Amlsq8tCLiSDi
OpQ7QBcb/MzIvcUnpRVwrzrao3hGULs0hlvBXA4J21WFwoBtD535enijRJVx30ms
ReN21whhjYDj9BI8i1Km07mzT5ixHNQcdMW4Sk+v+Wd9PTT5JoM28tF9z5zO81ax
yt7jyuODVXfiZLyQu38+e+Zm6eCyBfkR3ERuU68H6UevVnQWZ47JjgoSAbCLmyFm
c90lvLCbFZlEisYbJ7xP4OPuTOS6gv7nYIeuNfb7+MT/ZIxe9DVKv7HbmGFj6EiT
d/aJGPJVvREIwH/ZjK7rGDr4Q21jUXywy6FMG2Dk5EZFmKWGUb/R8/r+UKdQZspH
WIbpXofzaXzdceZrpiz4qHZT1lJ70tFDYRV3QvaN9Ov9TdiQVdq1181zwiBRvwAy
k4uSlGizeFxUYoG1a7BwPUP7pY99tJfntOxIrNLKFqO2KKMPFC5XPmjZ0Mht1Jbb
9bJCzdOh60yIUBKv668eORTR42Nb3h0zbqFY3lJ3J8nGaT2ndrn1ryY7Z1rcDtk1
Izp6V9BIg2BYJyrlVja6yXF/2u6kyHQw0Dy+Sy5DWzz4klTWgEF4lgPI/kWaGaSF
4ANk28s4mkDWj3Tk5LBObJd+mvaS9G7LbZpqbKDvrDBH34udHk0lhUJFCG7Dam6Y
kV2gc+SHCo853yuBjbtNyDF473Y4lc4cYCLXemY+tUJ9eJArQFuH1nTa4Lc3fsXN
5frvtH/2FEiVYJEdGdgSl/wn3PzI1Hle0TCm9ObnnUJ+zUvlquFcdyXsNec1ojWh
NQSOW67HoISGnexcEeeDfJdLCPJfAkaz5rRpJ3z5HAmSYrkxnu7cCsoXzQFda+Mt
rQ4RwhH+3N9k9rYac++B9Zzjc+hzhCU7sz1hLIZzJeVHrKvDGHez9FKvaDXA6BRj
9dWv1RvP8CcXgfmPEHj8KjAcpCl/Ajx1aiiqzVCkbTyLadFU1z10dqK8MpDVQ1GV
DPLx4PpCabgGhDU1DCRQcA3a4Xg/GiGmmhKi2pcz2KwYjcaTuoAEAel2E+6F0dI7
6sMxIjAHEXG951iyBw8Y7tWa9rVtBTFntL0nP5Bdbee/tpkNihpe2Q+fJi1IXitc
GTkG0rq1uc16XhOjPnQ0lTh3Mnz6S3SYBRaQYuZ0HM27V3ZhMCQ8rgNSya9w5DKS
camQPGO7jSvQ7fPFHhZ3T5/B1e3QX0XIy2P0b3EEyl9nVQbuMVwzmF7aW4bCoEm7
ciO84B8qNAvHLKNlRbrb7iIt09svPAcWOL5THeZ9JsGDb6KhJtRrXVy7yugJLjte
eU69A5b71l+qNKc1VH4reJzMdV2vmtqYLfqC1o6ibGbXXxvOHj+PS5gFj3shf9fL
wNHGVnM8iGF1/dXI1Ma5QGyX3RPZdkg0ukX5etC2izd2h3AbA1wO7RPiVSUzJ7PK
BNGtdF7mzc/jVrMkvsrEsJDp4TXDv7bght6wqpTdgSWuWoqZvhapNxCQcHP5Cvlj
1E53nABFP5/vy8JkUzXpE7j7i9146ScbLJfzhc3m33QPhNsRpvW5VzG5v/kgcdVy
Gn/gwGdF+nzi2JRH3Ya+o4mW3ObniJnskBkSGQWqPmnkkbbjrhZhPsxigA6bYJk/
cCuzSVmd7H1ZN6xjYjg3MyXuGm+DRoXD6JhDY1Y4flA=
`protect END_PROTECTED
