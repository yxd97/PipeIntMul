`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9NsNZu7An3y1NVMYWeU7sTvryQ+hUQ01rqFTAM7tbjl8UPpESKPp/6nsQmdbQy7o
0tiLSxwWElOkjlC8jGrJ+SNIJc0+6p7SIGYz8BCDcKN2Eb/xxaW3xCbE+8wYQdja
z/PpRe8DSi9lzUBXnnXYOI6XWvPwKaW0eZo9NwMqEOQ1kZzXke2X4ANxWHUdMlaX
WJ5KIycQdHCk7omdko0QWahzVxbqo9VEZ7dW/bW6wDJ1O74L/tYDv3pfYyOlNi5U
CvD65632K+DHuA38eqmmEgXck71hMjCIGvcNMeUbv6RlsDKMyzuqjQEiRTXYu7Ae
zXYvs+g8p2BsmpNb0b4fQG/DuBBQGWwog/KwnPXGO9YFVwdJEmzk6jysSXiM6bcm
tWPHxAmWiAs+GxSCU1YnedIu9/PauZ7QTDIRB72cfUflfUXR94Xvb4xLIdcWfaBq
`protect END_PROTECTED
