`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUObMtOcW8Tx7TzBxfgkjzFiuF4QK1MPva/9yYkPsHX0W046nu1LfcoiiGBbtxD4
A2nYr4vODMWV9/QpjVpbIfFjeu1xn+4IN5dC1kjxN6QABzz/MzkdJqbAXmDt/WQV
RVkKj4GkLBDR7F7OIpa6gZwv7wwqq7OX7Y4xQejhOe4nN8nKdwr9zC2oC80a9/PL
8KAMIsPLo1AQlOMasz7ids076vZHRD5DzJAhzssHXAOPkE4URSB5sKKmLFG3xXsY
1aVqba+WR1qUY+8PBOIDJc0dn79D5xkJE5Jz68SUcj4mDa3AENI49HbhpLGU6hU6
RjBKfnnmIr3xdhU5NasOsS+Cu+suznN9dx6diIMCUrA832axqLUGl2KSPtN4iFlm
cdKOnN3cT+6Lg6faE2x7DrR2j6Vq4Edd2NEZx4WoZWDEhTeMi4jjjLC8yq6DiKHl
fjnK2M6lDdt9qSL1U6op0z8xCfsUl+hSLMmGi2DNIhKBuTE6c11odAuKCmtaXsyz
quDc4Jzu+hFpPt8R8HIbAl0oFzyH9uqkvCfMyG7aVaG+aVIMeFVspVE6PtYyZeZU
vtS41sqCuJMctjI+Q9ja8/6cFPicD8wytTKLjh0vzVyxKw2leC+4ycd+QhhwSFHZ
Dc5RUk0pJSc8UjbhgSlqRiWrUClFmR2d1LimRb0cfyjnaXFGRfBpmHidNQBw9aL6
KnYrTEIidWb0ZN1w4p6Ky0V1yQ/4MRdo7yNpQoGi7rdP6v0A8Zsrvd2xTWizh/oW
2x0qrNixflUXgEDtAO/7oMHczS6+vFgS8E6DGg3XR4oKRA6lRLmK0oYQOp5lkELw
8MWlPYxjqR44gcigjPcZ3uhZKfnnsX0HG2ep1TClf2tPpDFC8+iD7JtfPM2Htebw
ybkEDecVoHyD/81B1AdNYP5puzmUKMkVCbjlA6DA8il7ZiT+jBSbXuBcLzjZhNkI
feruxay2QtqkThtxGrtIkLcxqMI9wYrLVYEPVpGFp6NjTAeOPXeNqZ1ECKVRwlT3
vqmErUzaromFAUk+VlRIm0ZN2elSS36jIYooXwsjml9tMDC648vatLHZrfz60OPQ
tLljiS5iZFxbV1v1M+ZnheohxhSVjOlfnTg44ZPav9IQ3hXqOLnetNY9fnIL4vDm
tpUfVpW+qapfSK2fqdSscGcmq2rstkw9wyb1icLlNsQmgZed0A2/EmtY0XEcyI9M
lobYY4GTHx7SNbwmy7xxLHm+QsWAF/UadHsIw5ITV6HOLkUf23XRIvVXNiZhzYAc
9sS07syRh+j1tQuUrndm5Qz0oS4jQXJMQ0W9z3Sl8/x6hhxo9Mit8l8UNVGH0vIL
7Mo/zZHbQM4ZAe1YNk7TY7T0TSmlsFHBRyORPB9N3FZOHp56DS/2qFTBOgYLsDXB
ds6TMqvdbs/mA8Qv1XBb+b3wXVh4DpAxqAMpouXa/yZAZtodLVeiuP6VvW7cTCTz
qHaPCPltLwJUquId/Hn9nDYi1rJRU4z+Em43T6vJN6VraiE6deOmXLaeQb1KOhNA
zXc5aL/DZwSM4mQ5Oe+LxIM+YCdYmjtd2SNy6qlPbUrzMQ/GOEnBK/Y9ffSp3BfF
Osba0QlWToKAPhOK7qf0WGk8pKQNO7NhJuByPg4RggVFQHsnkHEJhX6+NsAT4ygL
oh+1QjZ0vscH32YYsFidSLSRtACR5SgiUxAm7gjD+xxquWPfcTn81kecpEEauVLN
uYz/ZXquyj8tPasKSDNRc9np0PXJo0O1CrBch5n6vtecNONJBaLUhSBpZu9KzDLM
5nJmEhyNIzcj8y+AllHV0UKEO+auiPzypXIXFT1tk7jM4YMAoMjReyCICghyp6SM
HQOKnDOfwB3ypitIq+OCIUdVSkx1hoivPt43XXwUV1C2i0+XsMoQqvxRiqvmixUQ
feuv6E6Cyft4KcmLgtzlC82wiFU3ypcpKbGI06wpd1HHe7E8/3y/VsancD/4Vde3
NzuTZzulYNFG8RG7ficSfYz9H56Fobj79pepEjVhynZfYaZjc6li0r4ZpXrE90IF
ndXgMCz5LrAxibAPh0mdcO1UvEBFgLKO9+BsYdbAiq3cT945IFdvwczFgNtuKphK
KgSEYRbQAp61IR/nL6/rydeykNsNvktZ2kB7Vp2bsGGxM9n6kOEfrhskA8dhaDvv
9AkQIjKzSiHguAU2sOTxHXC/CMV3GSSe3Yd9Y8yPfi88PH8rd12BB5P62cigONZj
XAlVxX4NnZj7ySzHkYZqpwZIrxpXdNoiqtvYCmk0ot1Ciopfr2Nqh5fFCnKM9IjM
gQParDZ/uwtFIFuG7npLqn/6/OHnNprLUfsisw0XNdluCRPMv3P72bpV2xIkrVL1
eGBTNrVGOkTz6etR9n5SDk0AOwhaVzSxrulO/ALIlKvIJAzi0rw7ofWsZUZpdXA+
jYst2ivz2IcCQ+JkTkFYg1JHHRZj5Zz8kIBCQp7EQzFs/lMNtmL7FPx5uRs9Otjg
U6aG3oLQUzZIbLgF64KcU2CXhfEapapHNjftSPQ7ghacP/pgbGvt9OqU0bghZAFE
tCBcMr4UP4arRO4ew4UIvrFnSGkNC6y7xK4qZh7We2IM6CuFQCwII7AZOtR3lNud
ZEUqFb4QIw7iafZObYfcdA==
`protect END_PROTECTED
