`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dda7PnkViduDMLUfQPhWuorBZ3Rl+1HqNPlLdfg1/t3scGIcZt0PGuN7Tb28y9VG
onBlN3AFZHwsFmGzd+kw+x7G5ganvqkNuX91uYNbKkH8EvdFVrUUuKHuKDxzeWZp
oZBZFQzB1MIBMLULUbkxRD2FH+2P0tzn4rzYGtofioKkxQH9Xx3ejU/21GNc/whm
kffZ3/DVdDcaNUsKNCnlln1iGFn0kfHuIKF55Fzzuhg1af9jejzDxcyqwVsg7Gve
x0QLEEAzNe+SeD17HATBPfndXNxf6rLJTEEuzsbeiFpDEYUHiIJkGbdpTFKQPAgc
DSP5uwnkDTlBfgUZTgST4lLGEyXixsmUS2EUiGA1G0/uZLpwcxqySYNDXVu3Yy2l
Vun8lrr8hJ4kQD6Qj3LN7aAskabDKRDPFZ1JWtSEVzSO3gxmd4JTqmjDkqPnCzmW
1g4IY/9iJlDl1JCyzdqZ2pkjttKHmbg/cVwLBjFrrcXbv50VUdycmzjv3vfZIFGt
BEaIDsnyTra0QgJuUtCXgmRGpUta6bwc3W0sJJuLFAOoXY/D6qNwNEmS1ThvHMgh
Mi9Qk9R2Zk7AHvOBqBcVWt28gqJp+Ktcg1/gqrPVHmuMuA7L4E3m7xCe45G/XtJv
pcdqQJikre6gDeAmVN9gAWks/r7qsBTFLRTZHpf4GUSnMFCpLN+rb5Z4014MidgR
zl+Ue0hqgL4JgDaU5wcBWvaZNIVTNWJgQUgCP+9hoGMQdUV6si83v/2qpj4Tpw5w
BzuJeObBvdouRXkLJf8zOTu6OGAXiCIw20nnISgtGia5MGXXqfsF24X0DZ5PqJmr
pe9ePai2g/b39XtPtQExwOEcDFBp8goAf092WeywwHNiqrZKtkNPyTXRUaYQHGNc
95JH6m6RJL3XHn476V4ecg==
`protect END_PROTECTED
