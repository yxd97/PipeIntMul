`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WluF+Qc0O5AMa8vE3Xh+85gg9bh0EcaYxKDQC+LXmG63bxIq64lUgos8UVWpXpaV
uB0ego9s1QslmHHdal2o59RSEUGQ+pFXqL8v/xuB5O/jTWbitoP54mDS5wwmJQZq
EGRKdj86oGQbIfOhf53g4rYKTwScaJCuQljUx3Vl94JrVY0woKClIJqYjp+XxQlY
W97ZkoB3cqZw/jH1nlqmg21y6hyXmeaCNL1NUUKeqh1X7v49NrrZ97PjunW0p6z9
KatUKEIwLO5kOeEYYeVB4mpzvR+BO8TYPqBr/ANpAvTbn57f0jaIwfXCpvj42MNK
s8Qs0ANHaPK6Puf2kdJF1zj/mHeVG/n3yzaHdQWFfs18V5lwRvQxsz8T2BAD4HJr
AXJd7Vis87pJHgFLgHYUm5r9GJsQnSIUssHUieYE2PxdWNtVlJDWeXJNLUENuZFl
38NgJqH7ARTThhOSHR9JCfVAP2ViD0Sc8QF7PV16WzRRkXfi/SS/+1dZv9pxfodp
yDynfOuyilHrZCrrNK/y/ts8JgVFb992c+7vH07gDwdR+G9LVSDwIpRDe/mGQAm8
vDQp22oA0ULPFbaf5ZpCidd21Uc1ivyl6x/MpdJhiLQ7XZQ0ILnRnEO7HO5C+3A5
KYxDHXPIKKFeTrHtTMI9W/GJBJuEkZLQcXU/13uBKaBlw1Cs1Y7rLUn5y3Tck2dW
Rlxu1BBO8HfNgdBBmTI0QWdahQC4q16VZO3T1Paj0IM=
`protect END_PROTECTED
