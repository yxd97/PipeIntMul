`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
igbP9NIRI+GruE+ymwe4dPMXYhUzq4EEKZ1If1/m+phuOoGwmrUFt+ulmcgz1dz/
3tZvIK85JpyzzgYTJAEM5uF38Ibfb5KJ60sOHGXixDomt/XGs76u65iU4G2NuXO7
HYf38r5SBBvOyM6rKSJ/WoodVeK3ICtymp0ucPFr1iu9UtM5j4d0UP0J0VK3j2y0
t5J7Ba1mRWBo/Hmga+LzoM1ysL3GiJBnwua96fHCQq9XDfMhVyQeNGL9s5g2wf7Q
nzVLISk3y18Dk8Ru/lW4evYlU+M7JBEuVe2hzjVygoAkcDuwmDMmr0Gx2cvaJzwR
iRndhOOgOI1jmhCrAOVttrAeu9yUUU7AmtehqEhj8zGRt45SNUFBIstqklV1HXa4
3vf4i9j5kH38OiM7vxQBVaEVvlVGGfSSAAEfMiF/ecbVreABt5FsdgP0ZlzX3xme
j/4aLgf0aBBatFMcuL3x7NNvFnN16iBJXAmSCyjI3DuTBxftv7+eO1HZnckO9PTN
hboKY3ft3C82nyBZWLSeRf6EInNM0kKRiOp8APDVSfFFctJ4RkORFrwKxGTGeuX9
mmacJ8EV6PKJ2B90wbXEXKtJhTaGoB31ZipZ+AKhRcDcK7m9Rfq6hK0j2Ztic8GB
s0cpdLIXT2iDVyAuB5YFbI5pQ411ItOyGw+Cs3a4aRNl/5CkMpLUh0yiVcV28N4G
8080yBw8QhtYANEXFU3fTqj7cq/7gIRVbS0v0+XhGwXQoXATb0704mUTgN4jwt+o
`protect END_PROTECTED
