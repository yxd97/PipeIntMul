`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkIn+t5/TKTmFgpLmn+54T6wWNz3S7N6NaHAIkA6T7rpAod2JApIQI7QrLafbk9+
EN+aG74aP0DzunYos2lCnH151Tls6EHxDY1LG+evwwNVTNcFUfoCsDEwqrHsymbj
h7k7a6976GMPb8IFzPm7ZYrlFbnWU/9Xsx835j0wXFW8acdIb1tUFHJwwtN0pMsJ
QgIqOAEQcpFkSwu4/CI4xXpdQFWjELXrGd91lHe5yu154ptSvZZKYXJreqFowTvF
V0hd6L2KP30+R/ywBjuBVF45dIJ1oLt8FmqzmZSvc+cpzL69tIFcU0y5X2n3usR1
piVdHpa2ZsOOE6/G8ewZDpPhzF3oXAXlDh5wcyOggR3VJBmvQ+rBxHvP96uImbOM
wRXVgyn9D87TVfKagF5k0aYdB3+TVvlGpbu8ArjcOmRdD7gm//FSnEjKpM+xWe1I
WbAYmImdonjTXcItAYkPuNnIIpCAtiAFnBqTjP/mSMApqpe5WkzIojhTmtoy82bM
W1hnPz235x1cpmBUAHK36lNrjUC4z6/9taW83NyI1/w3cRwF8Rv0OivRvVZKLvFT
lcvovaptFS+VHEmA9OR70Ax1Lwu4rzGSLThdZH76eJAc67pE3k9+XhgDLiqtP9GN
NZJzAP26T6FybIPhIZzaxLqTmFpwikJa6Pi3V5PnJAzOH0c91n9WRThwYmSSOQsL
aM7ZZbQKwWK+ce8Uf0Xwcw9zz3QSbjDt/EgrajiNVdPmtSELOzoX4V2qkJDSNx1F
rvRaY30on3oOYBTJ7Cgn+Py3Ra8z00L15x23kUoNlrw=
`protect END_PROTECTED
