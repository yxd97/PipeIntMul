`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwphQ67SfbgJranz2jj84FsTuPXycCyyFtLrKR0GY1TFo6+12piVxn8zMJG49tuh
dGvuADGFGlvYKCVE3jsM1Fc90hx30KcmYj8/ErsJyOIiyZ6022lQ1D5sKmjejfhS
oUpzMn5i1X6KRuJQI3yvrIXYAcqldJZ0fL/wQB2U+V2MWFhjXqxZmTwU/iwjQTiz
d17+ZEUsFMlKvH+Umvu27u0xY+IGBklmCwM6X/VWuj/pwPbVe/Pff4b3Aor/8JbJ
h2Uxg9gOdbvb4entSf2/at9bV/CI+6gAW759NKtQLDYkGkpRqtpSV8H1ysPxF8Z+
6Fl46W95/nZKm6OxtgSVuVomkJVLSLY75EKxNlxlODyVmPy+bm4EekTEA9znTVnQ
W18+A1P8T/23/XFBWDMoU7o5J9iBxnCUkIgVmTWBA+db3yLZcTNWUAYXVOK6o/Dr
XzY6E4pGyLW3S/6kYLVkLOFCZwagw2RDBOxAlR/N/sdNnu//5LDsHjZka2Mp9DfF
fbykufjdk9hY2IVOFcoH2iUHPQd+jLMJpxa3cAA3d8M1/HYqbM6V7zMg14T4vbu9
wgVSBHzu2yh9SizDX39muhuVsWkR5k77ZCbfplQ/vIYXPqYAvOzRk/g/ZXg+cSMQ
83ocyk5cSLhv3FNo++66WwGHYIQlUfX7F8KceREHnGj4E/MD9qzxPrXK0VOxG9E/
IDN0pavA9BMjoX6oRp5Wt10sWytTRno9duA0Ohq71KEWHDzA9jIF5qklci+zj5Y7
UXIT0a7RUth1GxhYCABrT7fOwtUziz1o/2+oLnqUZ6RaAr+FmfSJm/iRVi/Oowkc
6URaVJzOk4EM7o7LuHftxQFKmGCopVLuRbUXnGauvXCcxNc7YPhYofVrwYJhUeGr
PRl/qRLK6ZnbkhAxZPNGiiygQP/UDnrJftSs4bwvktUnCxldD5uJxa0wHPbCRytb
n49bsBkatrR/iiPZzLc0RHegEtEp9OJ/8IM0xUIoBA6jVauLjS97536bY8wBLc5x
73Obq8Arph9ztdJiYKG6R4i3iCa/fW0KZiUhm7YDHZphX90sSYCy8J7sVxhbaBrW
YSIruZKNXHfKx1bdXCB9OsiY9up2neZ6wMELjnljXQj4CdXaSOz8vd+7Qds8+3L+
BOkQn751jxBnB4dJlvf8ThhdTON6g0uoKfLTEUvDhHMg4vnzItM3PnIrkVofcR2y
rjXRxI5hSt/R4OzL9dMyLPK3lUP/WFw332YdAPM/J+qLG9xkNSnYwsDcGU1Hme6E
ehMSkl9vDAkXtzYkHBD2G5OxmuG2zPq0VMMg7N1z2tPTXDnh6oHw4cYDDanKOfzP
a54VFxtleRBT8DJ0wJDq3lQtho7p6VyDUoE3/+fgSDIDcnff2DHDkIPJ9jmY5lQw
mSAf1vFa+WnLD3PiAhn+uEl5c/JPbAe/tAW7yqQWVTHqGP4b41C9JHZpm/CZESv1
fclQz697rkySxsLDLPVRGMDRpTdWpgfpAhT/zjC9yuL8zQ5Erz0Te0bf1MvkdIGp
Z3szdnxATMPj5EoNArgKfoqs5Vp4E6cjcOdw/tHuZ8WnG864YyhEnPO5YJx0Eo6x
RGdggB0E+jYzhNDnkVQqvjHVLqo7Hre21H+VTko5Gkmog855EmXVfr1j7id/zt5o
knp9VhjX8jm0reStLP+HA4mBP8j8/g/N3WPuKbPLuvzbHzntfF3JaO7f93yeutvI
r/Yo4HTjH5qs5JYXNlyg28ZgxYzBpnz70MDkWPLtb9hJefI4WBW321RKZDP9u8OY
s7VOyMplj4RoP/9gjc0hVQ0GLKf1yh7Tj789EbbDxosVdIfppHJYIIESyaXPkHVp
5iJjCjzBX0ATjxP0EXe+/vU5QS7bHsmyH1tuz5Nst9ROe82wAVbAyNVYjgqp8ES0
+lypVST1dBQWujV9zXHfxHQRraKNH/2LFI3Y+vdgKov2cb9iXB3OZ3mfmivaZcDJ
l4WTHtjozm7QD4DW+xWabQ+Fp3VHWgWinzSU4F2nrhxNDmYSYeWD8QCMCRTOMREV
NCuVPHmw2uXKcsZbZTNOMgkYoe6D2y8QlH/BAHpRVIdM/i14GvHpyewm0wf98YdI
CPVzlgG6Xz6DpSQV2tAwWpy91IQ/lgpOMB3BKtXitabrxkHi6py42H2PlbG5kHet
JTv4GzzluThfZ7mMN1CYw7dTQXPn9Aet0VoDiSm33oOkX9WhV/CuwXPb3dULIyn4
9KWUzXwoRBMOhkctbG3UKK4v42UDE1rjyobvlYRi9irNIH8G4D6/Y3gCdVSgRfvB
BHlD2ztYAcXq8Loj0f1Ns9xwnAdNnP8eEzcmlKZ6yxrV86iewgcffHwHGUqislnu
ui89MwdWO0IcOIyi5fiNCfOG1kY2MhF2iF2b/myG61Q=
`protect END_PROTECTED
