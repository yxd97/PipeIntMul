`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/k9Y751BouqNQ3g74N7w4trcxQF2eHtDE2dXcqGg5dIfzLRCvpU4VYoH5gz5J59o
gg6Hxau81HzzSZLozS0ZpjpW8FBQ1TXVmR6oTHUiiQoYLnDbhFgHYqSI8K/EDxkD
VGeVcyWrRm7ZlsvtpZ2ZnB+DQ6qMOK5oJkEMaWGnVZThTOmCF/6+u6JTcXtJBvCW
6BgMc3DpJSAQpwgD0zxx1vxdm0C/DkBLgRI+qnRSwe1eeIha5+5eW52g9IBLw4gZ
/++OXS/8tX8usKpqq6lrQGNsZQXTqkrve0F8qKGjw6YZJ65adzug+2KEYbqBcsso
MCuBy1zn2s0G8Y8i1C63ydY0Nan0L4kSnvtPS/fVpIxgIMdpKKbSbgd9Q38ONqyi
SsgqZakxQeNzmb+8AwBKZkw/S+0uZ/uNBB6G0Wy2fC9EyrrhBsbgLZpKb4tgxZNL
7uJkKvGhAVTI5kk3ehwigg60JlYgo741iWZyOgTSOKnLyFFdkklCmlV0CDf7Y3xu
aXRz8PBHA0QNl6KIzC65PUhV0f9mqkN21wrlkhnpFPPG18ZweGXzyGQdGowtkFn/
9+UAJZoB5uPk2cyoTq/M/F292nSmPkCCdluuYVmACn8=
`protect END_PROTECTED
