`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGpa80a1q6rXjMZhwCI/1W4+JMG1bY7mkEHvafsmucX73qOQ4ZUgUqntQ0ZZ8poO
9oM1TUWM1v4K8T2whV6yRmy7WS120OI7/baQx4mVAmSqz3H32XdkSuj2IfBQxAcr
BKIj2udvdmojSMsHGxBL3dxgcNTBCGgfVd8LXieH4inQ50R98hi+mzg1AgxHd2y4
uapudh9oHxqI2s5PPmXfJzSDSdrbpCnO65yE7YHv3AvhvZmuN3pnLz1Ykzb35CeZ
8GT8HILSdjpYtE2wBQ7o/jY05ofi/IDKt5C5FCAeK0J7OnCIKz2EhOrS/YNNBopN
hNrO4ntyZPe6ivFeSrWgdaXlocbWzniU/Nvf++bZEuOeabHS343PZtuZjiOgxI3c
Wdmvgm0YhoGMFHaG2hMIATKKHPpIiRrhD0N9XcVmdlkkklgSGwygy+oe8CNAvras
T/d+MAKaqXVSwVidSDcp+q/0hNrify0iR9mxx0bbFuRLSNKiy1oCoSjPaP7ypdOO
qcQfbkKUUJrs2xh2R1amv9oimGY3RV5f1nTEcQ6q6BMJf68TNjeVzo7eHHZcMwPy
9d/NSuCJDvE2FNXZ8mMGl1nQBeOhlIFvSemTgPoVx5EQILpSBsREG36ujra0s9jg
6De89TD8CdSmuxZuTwTxsPl1Tf/tP4G+i1O564L3yrdpk2VdfoEMmBHI7sNFl83t
PfoJGK8HrwISpu6MAxQi6RwLuWJDxnXEWtYj07P0C6W1AmRiMFjehfuVGh2Jlnq1
jS1ml6KATULSng1pmPRu3hYE44X+RWRlcF/hrtozLuZ3A27K9J4j6WVUrwwF50cg
wiIoLwg3WzfUmgdYY6+U55Uz3BrNKHV753VeO02Nuns=
`protect END_PROTECTED
