`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cmbp3oDPCZjcBlY32BsIH5SYLcj/ZJ4cjT9WBfF9qx90BfeDcuoQVHuz+SHCjX6L
Q+awIVx3B3oWg5jhNJxw4y6XUUcXYxTUMopqg5s/O+Nd+yVIcJeBa19B0+yiPPQ4
gxQk5wAqIEK/EexCooBO4YXxxQ8HWURrMRmHEu7MDnX2BNfHb7iUnmdyf3YBm4MR
OhEE55YoO92Z8sV8I4zxFgZgvKAcNH6/I+4vUf+3pvyuNHal5LGgQHtj8tEVFp2o
8EyFBTJ4I607fP2xbK5xoMHAeHgAXauRygOOkpqcAffuyX2yCeTKZneqOcbzi4vk
8R3mx6h2BPDU7d8iRE2aV3FNxI1MDocirvIFbQR7HDLc1+S0AR6QElI2bQP7P7jV
`protect END_PROTECTED
