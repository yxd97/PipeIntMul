`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZoF6LTokrH506t2N8XX0jJzCMcWp2QM+vgUhZ2PfKQBv4H9tJkh3ymF/KLvYLbc
AKIe+Y8iArF7tDY51lfwziByipS4k28d7lV4IubRe/YDH/giPCNOKrYA0UamTrcf
Cmr10Sk1vvw9VqW55r72XLLn9YAbs9jW7B6FPnNchTL9eXtEr/LjSvCvZQr4qiro
MsTqeMokLTLKAsg5Z7HJGYxVTeQqIjL6/sXFh9InDMOCXJIjyHjj+LGOWpzWoh+y
9jDLHmSGQPW4Ez+43PcAsxIOhc91cYtttjoditD0BFDeSzp9IQDnRorIWC9EnHbt
JVp4l1LR+ceal+Gn3vRB2+NMRMdEQPMIa6vbmOHiL+rOuHPWcG8NYqBLU4DZ9U1+
GyOqhd6n3Aca/0RW/aD7tZUsJ275ZdBLwZyLXP9jK7C8dpDRM33HisljmwhiAq0v
09PWPGJ7zoFxsbAMQRG6QrAMYIjyy5FwRFKDhwmjoGbarVprKWoT9iuRby15wF0A
hm3ydLcBrxP3cN4L1hfMbj2mJJPUGyDnHfd1qMx16c8TbrUkdgcDDQIR4myyQoqD
0Ib5MehiP7uCUmDUait1o0Q41lIEa2ApxcrEFXKcx3HizKDi/77Oy/IiE9G0jfi8
McLqk3nAdNn6L244A1PrMG3e7dwAd9hU52dnTOf0UMvOXi2kfexaN6Fgac3NPpKO
bd7mL1zZkCwnMNiXT6q2FiXqBugjAuH4l1AKwlTowrFKKNxpWygn2iLzw2ujWQv8
uQT2GWoFrcsV3+aFHqrAzaMAE8OH/KrOTPhAUMvyWE86RnJ4g7HiXepJO+juxBpb
0x6+/ZSqKxIMv6zifSReAASEZWQjS64zkRLMfdZkUQwL7wD5kXJZkN6yXquQ73V+
jEQ0a3m6M4YWltyzFILqKEA2PEcUaRyyfzp6CWPJs4UvdoBJD6/U6C+nfdWpHqCe
LDu3FeZhNP1sF3L2U1jcm76UdrOCMAgTba4idF48Vfo+UOK+zllajoW5K5PLLR48
J5/I0bew2oLq642aGFKjy1Omtx1wFrF6g18FKb4PU5xLB6jy2NuGs+ef+5tGy6BU
Kd0CxVr5zl5wNLlzjgEkfLtmZFN0OxcIJ0Vq/iO/Dybq532DN0x1+Xo11LYz6S3K
`protect END_PROTECTED
