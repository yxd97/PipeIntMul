`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gcOkVNIOVECRCcdDAt91oicKW9mAFkKKvsPODzZWpbXYv89e7kaMh9mF6KFf5vvt
6Z5kGjD6ko6pf8/HRHKchLc5KlAeymuxH869mGYu9ydqJLCLi+AekEbREyBI+70l
YSq/Y147wDMNiQM/tFaQUdT4GpFcYbYcErfOu/9vacejkWNTh4P24UQU5J/9qQoE
rWfsJDugoD2TBjrgp9NXb5F/zJdiO4MksZ9ucZODM4Dl7ePFzR9kt2RFcdfYo3Qr
gUgZlrDHL8bAXyB0LawZYkilny2fcdWi+W/F5N0rI2tNnu/q6kG4uLo6CrD789DZ
5VwW5uA8FHeTlmY7pxfYn8rMHBHvWGnG29o6M5oYe+mdzY8c//nLvA85wq8SJRV6
006nMoehPzQQuIG2Cn84lhh4Mpr1hvx9K16ddmV2BAT6YDTIypZobsaQS/LXu1i9
WKjLUKYQv1Bh2ZaF9CL8bXD6jO860UeZ3CY+fWpRQGyxC1E/WPLlxsq4D73C/E4H
60OVBr4uzzEscXHUnq/zhb7ygzaTvY/OH8EnXcDwztXq79NUNa7NVQpxv0HCF/W2
Oev4wNZJ9+h+LJIwLYU6rIx1Y2ueauNsATJOP31nlcGvUnlm2c+HrrpBrdZ5syq5
JUAx8ixDQoGdFyxtK5ayCUUvOxLkLCjcsDXkt+BUPZn6aMlKJ5jspTSXIFF8UQ/J
xp66tTexrGKvxMv18DPHuUrNlbsI6qtSyAZ/Ogwpfh1/8QI58TvPSemJHAqml1V9
HWHiPOHBT9sS+4q8zy4vOhUwSnHuaNiluJdr4rwW6ZZ9n9/TeGFjaGBvKAYE2D0M
Ru4YznL/zAIUvWdLQq7gP8gH0FFJu1E37OAQcqeBHRiDQbsIOdI8F3zM0xyL9KB8
COKSydCOiC+qq/rlGaHKQkDZDz+wiPdN96hVElxa0Nw6PVyaYnFvtxurOQ1bp+wU
`protect END_PROTECTED
