`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BsehiUwjWJRQQCB3QdBe0cYcBUswxnWgYIJC3Uazo2wzBuJ78AlPdB71z1PPehDt
X6N8mZkeMCI6WgTieWVvf1MpPhmTZw0nHNPttEXbMeQWaBvB+DurEH9jojIrFjEZ
FD9PszAdoSzG0woyZwaZEuut8aansZHpX1NosCAfPwIchSP3F8ySHZ2ey7GVA7OK
XT3Uamy/qgh9wDFlMuZsxsznyGKe9A5nk0beQMWWn5tDxSD3b1VNyQ0eOXrboRpf
aZpXA3jf8Sk/tyU2vJCK3PuGjmOTQWl7JGSpEnUI3+OBsj4XZG56lUlinAz1Lxku
JioUv7DFdWRG8gElJAWtA9ik8B3X74qnc2xN7/vTZfQuP8SsbqcbUgkJuzEdfVGd
JSli/MlfpbUh28mr4Em3Cv4SMqxFpkOG9XIrbFbQbsadBzph8ZLMecJeugYmMNIz
e8Pwx6FWdRna2252CgLePg0X+V584Zm2i6A8SCrQkqwDs3dEZTy2t2KEsKtN8q2w
s5lPU+fDEzPXhGIjvUSfH0y+PPYrbDd62yAXjRPyOY15vBzFDWaCZBHUBd37/GlE
zay17Dm8JqbryKJrNmTd96NaJWxLHI303RgUG7GaRkQCPv7caZZHoTyCVYxCi4ec
jebI2ipDebvs5/Zpnjr2pDzydFOn+pDFGT5r/sxGkRPiKYscoP6Rq2vOshRIrzXp
U6pB7/ymQCWHunfOpkIHHU8SC7Y7im0xKMYZugNS3LaFSh5xei0Wl9Z0J0zgcgZI
JecvFTQHTRr6Ko0XEHn9alvdxuDvDZSeiTS5+9xnkeT1BxVIW2SGIGWOYD+FluZF
DwbzD5UKPsmIO3KzbboKJLRNFUBy3l/8ScalO+AC42C8iEiGv8Cwd28fONXSgYsl
AJn68U5rTo8WaaSMk8Hfd0SLjidRr0rA/Pgetwci3RDQQVce7IDgaw4jOZM3p+8k
o0ozzCPbdMU2KKsnW/tUPz/ZkLSH51oecvNOxoC57u8h0kWlszCKnGnKX5Ha3Dpc
IS2LobGSAjkdLyAves3t3FCuPHDDlp860ksc2XRXE/pQmk7MyTF40eOhzLWDHO9z
sP5Fr273uL4gfswjVw65zwJjs9WjCThUJI/F1w2p57AMB5JqVIdcNvTu5HmHwgTQ
Fu9fP/Mpb1BSrBQQM8sMiSeQTKTOy1fGODrq3wA3oDVh5wNDmMZ09atNj53vq3Ct
1f9pW+ZypW32T1fj9gGbKirLjDsAiEsDieVbsry7X5Xdd98mdA3bIfriJ+Ek/7Kg
nQbGvllx9RrW0tcu9hBvhQfdcML6xcEHwWeEe5M2dW3P4Ak9l7CuuIpQExugb8GU
L6f/FysYVY0ACC9ZWsb3y+hTeAeq8LFgRE0XLdehvtUMx87ZX0jMIOl3V+mxIGj6
gO8lwrDCEGPVv0Um8wzn5EVcfP88ugw0uD73OqOvdfAYq/YNghN9ZQ9Z6tVIeonV
ljPdemqU1ayrEuVURkhaqBjLEYuirjm+sgPvmAVNSQjny2xAVDQtK0f1w5plVfD6
mM0TwdE+YwSWdf3XJLldIert+7yk6j3m5eWeePWKJ58r+AYv20K1JDzXu73tYTRG
iQh4S0jStXueaAYvrZOeiO9IQIjXExGHAEwoD5gfl4ER+gabFKXQe5R++hKjydkq
ljwQzMJMv6+0Zi9x9dz0izpoHhu/Uk7nYsHuyXfjQQLMvLpBzxhpGZerwUaC6uSc
XTDFDmNavtK3Mn0OkwVyUnqElphJUvxxetKYWqkEG6nJU5xQUpAvZsEC3HucO8t5
+C4uIery9/V+XVYfMdDTl2h0KhzPyqlqIwLbpPvbvLqCzMkGwi5IJWMrkJ3+G+zm
z6pYGSwUtt2pUhnhISN4OSBuPVnra00uV/vFFSo2RlMqr4LJ0593wobj0mKSPbk4
mrjc7SCAz6CQO7UM0EbqPx6wzpKI0BgZ1TDKtJh4rQeMdx3nEz+3GFMHeVwAWS4p
QMpUt9uJdEz9e7vqcJZEG8xOoihe7nocz+W4ttCbeMY6TtL534IldCgsdb5QbjTv
PUv3rv7MtQZKG/0hqL2WRMzwbReIkdREsEfkBx7LNOXK2YAIERVVtBSSuvUEJ01M
p02HLgLBegqR7AdPXwdBNIJ6IVr2TY/k1QPNv27MazCzso97HrZ3eaqh68QhZflb
AcYpb+3mXUEA3w0J3fZjW12ZJ/HJZXqUq2pnbEQWcCk36r33odkLrS9ij3VX92P2
4OEQ/y5YnrFlEv9N9oI2jugOtpLH9Mn2Vc/t1K9TAh7XWcoOd5/F009Qf/OLaDhE
Ne+R9LvB95QGCy3WA3NNBkUpTRqB0dDmWivsskz9vcuiVoU5P2GKvppsx3if3/1X
bNLUkIjawQHiWxBYH8dCMSIRWjdLLLntqukOXLTqE6oWI0uxAmt9uyyx/UagvXpl
65P2XC0sRpH/ZBLZq5D6ksk6GfpdY9exJenDi3KsMkdoQK1ug/7gsCImy7UrwLEZ
leub1U8C/FMsIzOJ8Sr5vgK+OIw3r3PrcJgKtLX5VOGeFym4bAJNALzhl1vT6E5o
7wRB3YozFGXUerARzsU9V0z+P7x/+IXLSTput/Ta5H/Z3w8/ayxF9/9nAsjGwpl8
SaRz2G18rizz+JEPtpvEFubsA3JRtEBddeYypZq8lJholrh2LdD2axfHuct7EBqp
VN5T3BHAGQt606dnGjKLj9QPpgoZFs+84Ut5CGIzHxTZA5+bxGWfmjIx4AYhMhsx
KRK9M7EmLKzLBEsJ0iNoRGbcCb2SqbxrrAegX9UsiUOfNnTS8Rs5iLUQ+fOoPifl
7oYWElQevQd7o5ytNcDlPjfI/gcYgOsxLIT5Nc+94buTCSm7f+4KmC9tP7jT2MKS
mJ0OvwPdQjJMP+eq3MT3KBBV4H4qWWsAgfKG71sESl1oNlCRQKFVisswBdYVQMt5
UB65XrRpdNDGBh2EYK7wr+Gogmhg00qXweihUIv5BjRqZ9QZVAjTzhDcz83uzIiy
Ehclmk1MmPMjeo5PvELnxhxHDMr86qxXVMdiaH/DXSIefcokVxbp2IrLdgmEsJQk
dLcfYTXCYnSh2el61OhrVziJFMGUBNhgIplp77pnYCb/jqlQavHHMETGcgNlgpyu
vLdaR5NdEdTMbVTMdcVbUFU1ryJg8Ziv6lzY/stzW+ihp6bdNzjiZJ4xH4K1JQJP
EHb8e+6xQfTZk5i+PDUpZDrOTry54bOmgRW8W9I7AaeADvCwG/sTFWpvRkytmWu0
FZ86OQPXoVzk7tYbow/kK84LWghAtOrO3SaSSVcDpB5oKOZRQo9jDCwhLDMlQXrd
VJW9O7P90hB2VEH5qHFT0/OKA6kuN2woMWhz+mZYupHJGdejO+pVB5WXcvC2GPrk
ltprl2JL4MfpzigK6TYny+H0GTHXJ9pN0G/GbYOBzRr9Jn61iOZc9QCp8NEIOxSw
xuqW2WPBUg0xVn12hmxpL7JKaNOVufYlSgf5zLQwj/XCVAMNtJM9EimkDQmRx45w
Qq8sEVjQfFPgQvGTuylCWxcwWUT94HgmZETw522p+DSFuxAQLPjfsUOc4OJ9TK4z
hokqAoJq7PjAD0L93DBFIE5qQNRpLaLUVTNR15XZ2RxOXU8BK7Gj9m7rf003gter
H+zC33S4bCyUTQLK0DmxIqavEg0vgTkj2OwtvKiKLmtsh0/exulDzvWdGxrJ61Gn
2qEyB9AbWYYQbU1ByCFGGImmWR/FjFJrWCeS/hpBnbUcmxA4htK0VsJrrZlQ9/og
8GW29Kxi0vzYDMsYZxeeRQS2uvDZ1bnEhx6Bn7NHcXShFANgpkQaBO40ITXtNulF
p5keR2GQHGSAgTn4ou32yPjvWue+Va3WgnIY78pie0YetU2sPCnnkz2g78zmsyZ3
rzdSMDCqGGyfKWb+66pg1GVKUrQ0dXBSIj/EeRrNNuGi1rCsxjCpicJS4dXbvLzS
66eVjHiDXB1qpqX9M3AkJr48AeF85CXhRv7NgyOIES3cqEMqmxyCDocXzs666hER
GW+Ke39dsmbW8JOPUox1WU8lCtIO41WXLdX3DJSFfn98YI/BREfWdrPTeCN0j/D1
gNngmgn/69aRJX5aRdxAbzkdm18hTEWHp9twH2qqc7mfl27+2RzxGQm4v8drsuX2
8K0HTh3hN83n4ZCjC/G7xKx8ATOF5g31SShyTdK452n4WaZS8ZMoABhUBz5SDTqF
znD6u2d47Z9YsF6ETMbJrNv9LuKWkAqJ2RTT6MyXN/qG8j7yWzgkyp51/3JSYbkG
Lno0yCV5VkEdGhIDVZRWL1E9wEQCo4XJxTXUYePnW4YIfpK2/iHnp0thGjwMHyih
nZl+eK/kqizuEm6QZAYFEhTt/Y9TwDBxv2UFTJ+p15Le844q7nc6BrZ8zA/JDiw3
+LY4U3BE4ea98KCkJcW+5VVA4iEJudY80DWoShZ0RAj/+HXKQiKzl/fHamq8YKcK
AA4NoYBMofzIiT9t4e3Hg4vTDlyybOntEZFGorvbjXwL+t8tnCn2qeOGAGdk5WZw
gGJb6eUy6qCn2p+teo5BVFhU6EmMj9KRWkeczkLw+AyqYp0OQxm9MAuP+Zv090Nz
1+7nFg7dpBm6lKXEGG8Et0B2hagVpGbEU4kqUfS/hJ6S14oBdZd8lJTiiTmQgC51
9j0/ZgUr8ZAj1OkTCpLhZ6ftJllwOQAtheHW8JKM8GXN1nrH8C5v7Vfo1bdJ2LGv
nDA/22WA1pokuowlK04Dk2KZcjYaJEq7qeUKrJv+21jgvfiYuFwYkHPQiwKsP7Z0
4sYk8BK8eM+rWV0MAaW6eVBivrjwC74NYwReGU2+QpQNSC1A9kwx7Jvo4d/c2n14
hvJNAeq67ax7y3geQCTMWraDMTGwXjV7bFc0E7O6n9omaOSgBV74NgyrexBdfF1x
CaovBqaO2jls1+lGLeow1Yyg51lY3axun7/+tcE+3xcOm11rJ1y1P1QVEffYLkCB
UP8a44NdjqzSaYNLXK+pDKBD6zTS1JMM24w3MDqdiW1InbmSL/D65Ow1WFvLWg4Z
QT70kXrVYCYArLnTAj2wSqiYzbojjGkMC8EewCZF3CiicChyVd+onSPYHDrA42Y7
fx/wegX5Fw7gkuPG5Vt83Vi2tKykkpyQiAN/cLeldIchwGy7fsRrF+7UBwUqf0P0
kaguZBg03Q5/2Q8z1grhgAh53+nZ14KWMtCUNtl//74+wGowSW+BZ8Q6a7nLK/ct
6y/L/QlZ+EKOslTqo5cOS85kSgrauAaFAeVdY6K3dJs5cguc1MsBd/w/ccO+cHbC
gQ9P43kzjD9QO4oYvv9MlIzbuodXFVyaVvb7xioMSo1muPAlJHzqAV4j9cOimMtr
Dcaq43afyrDoHJDHZwPaSR+wIFQ9lW3bcYP7TKruGNtUDP2qiNUj2PbaATpviUMz
TBKsw9vgccuaAHCVwz3JvhKLoOOZOdFfjC/qBeADWmC5I3DXX6YEShhLs3CkoC02
zH103jYPE9IMCpyz/aJ8o6LVkZWaNZdDU5t0tWppgbkhATHMH2R2o3Bial+IQwKO
OtCX4vNbxzxqZYRxJHWDftjWP4NDe0r1k6QIZOygcPa9wjzztmK63iFKiSP7VTZj
9PgFbIfGNmJqECes/7r01q1WnSu/GfeDlzztdMAUynzQyVIC4lu37FFA1ixo1GBO
tXhEAacghXOMYW4I2seaR3M+XX6zk+g+8g6DjvBTQmlsBEASUPEohhVaSUnyz1SY
zDxbyN8G8aVpWvbFNlcHLpbF+abeFnR+6PtXLqpcG+VAd/OpmEbsF63yv9qQC4Ah
PiaYbjPzHmFp8TfiwKMnkoXIEFeBGK2D4MbyrE3kde6A+tdEJj0RtGjNXFcH0RBB
mWrmWXIDahSelBfUxqDfLHmqS/TC1c7tfWRU8SgnSIQjk5dxpIQqbDX032BjWpUa
`protect END_PROTECTED
