`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4bUW2bS/hO7HWhYFaLT6PFiUyAyMpIw8zgSAhseueoHjHIPT6laEQAgdYw1RdpGd
zf12xf1ZyCviXpsfXPh2Kh70n7eXGFB8QAMqjWFFTo2xcZKwxiWVoRD5kETVuLeS
pxc7bYJBs04T8Pu47yuzR0CTZRsxTXTkjtbyfExtcZKDsKyUEtnKmiwETEakd4Tb
de/u3nF46T81mCCC1ArkMIGsdJk9pPaUp2VavBNg8X0GSHZWbDVohTiLFQxHerZt
e6yvWVpuKpaqKuQIRh2EVbrkDt6buKw7+9I4XBs3NNTlvwmYIu93cgTU5J8rBHZN
C9PcFurfj0MOVupnBZ9l8q92IOIMrZZVpmttBDI/6txnf2VfLX6OT9L0C01axf90
+IMxk3EE/RdPPAOCxukgiHjEQpQxs0qVfzZQz7aT0FTioue5lCbNPNDHZNQKqKz+
OHT/H1uVYaZbLH0MWWjtYpmPjfqLdUmpDt/fAoASXvn303AUGd4/SL7uGvKhKiSI
KztrGHUu+MKzTAoddGTQ7xZacXtb4diNPAFBuIOiTvIJjw7OJkeD7xOyqrF4Q6nY
xuJ9SUP9VuojIlAdsXD7uhgXTH62S8CaZVann25EGz0W5DHAFZatRegsImDeajqH
Ow0Jra/2lqDm0udnS90IUJ/4HGkYdfVs+Y2WVQXsHFQO2bTeAUfMDTm7pOc64cEB
k9Xaj502JQ8ij2B2j7A0ZOxLFjREktDRkI1SWAMoSNOOLFWNUeTbfb2D/0YJiSmD
ok8BfKB1wpY+KyeHegMBpg==
`protect END_PROTECTED
