`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9ybftcd1e0/C0vuc/iL4g5OgywhXCLXtSfqMwGxioKId625uUHtllS9vTzJBJ3a
PoNiIka4AEl/M29TLF/9tbWgrkfFIlLEf/Zaa3FGc5gUyEpVNrk/xhrkMsOeQijS
XjXQ25SZEZ3LlSe0dWkPkFgOfbcd4NdUSgmWpUJ/mRHjYnahRvItFK3Mb8qjBL/d
jTvh7mMksPq8Rk/cS7wMJF0NReZ6yDSVYIeadu7WBWfad/FLWq8cMNzDr7p8kpA6
/rcz9NtyL7ITgTfKOI9kFAbVSPZPUfMiPEFE0/uh+p3rQbo888KrfrF2ml2+8BX1
3EX2DRoWb/ESvPPqIlRywK4+GwHvPd8Jx3wNsLb1hSW/CapfzfuiSSyz4rX/BkZT
sJrz0Ty9YQRGwJ0hhZ63zhs8W8S9ZkGOOz+uR1iHmmm7eGYx9W5nGkwh48r04Mpp
Djtuh1mmLZbu4pKbIyA2zwcFIHsY8mmJM8US4+L18Lr2DSaWB5lTVMUrQRPm0DFf
41ClqiSWaBabExM5MtmgKqC9bZ8P98J8KLx2UpR4o8cyEb4KffNVKQjf/VgtQkie
2IT5YT2FMTHLb4MJnHhCH07YNJ8bAwToN166TIwe/C+SIdZoByx4Rt7f4L4tE5DK
FR7zWp9cycPP0YBtytcgkXL5FTwbCB5AC1orKAxZc+tqJqLhQbBOFOePey/DOm/h
AnzAPtCj6Kogf/cDzUJx2w==
`protect END_PROTECTED
