`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMsjZlEt8XIm7DdqJgB3uj/pASB3ITtaEyqpNJ6XefawvTChlEJitvPjN2s8BrpR
AwKHbNtufrBxD1ITtAVxPrGfnuXoddAVHstYWpEdFe/Nf3INI+dTmMdAnQXAJOgk
3boBe+bjEaTu3Du9W1mjsNXhv7I4EE9KJOPM0eGK3zWRdRl8LWUhea/Pidf6QBZm
Ub4eJThIwKGTgUxr2eZMIFrQuBdA78Ipi/PZqVbOW0UrJ/0UW7+tjWV18qz1tIXy
y/EDePhDgzvvz7x/IFnv7AKhMAr1sel3FcjoNqR//x/S9E6brXC36cK3JEGbjT0t
83DI8lxBXjP2VQ5a1kS4oiEPQkOWhDhVda7o1gLpAEGXr/0Pn96dp7x72dFc742/
NIfDh/on1VFWG5K0oQzJG16tPB4mwYQjpb5mn5zlX/Xthx6YnCIPJL7RqtUFyWv+
VTn1ATm6a28tUqKM+eob8SIsVbTG9a8fGQIb9THTLN1O427ay1VgOCsv3aoa7QXh
`protect END_PROTECTED
