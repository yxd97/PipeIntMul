`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3uE5NHU1khPpiScv7rXJFeMxl7OIdOgKJOxMTIDqOfeqzMXz23z3cbGmk2iS4d0o
4o4UVtdFpPcM4FpqYUs/OpbyO/A8Npt0Hc8o92RH76jJp1LVoAKQRmX0MWD31Kqi
3zoTJfScAJGRYcAVcDdHI2Ddr4Q9uwQDjmM0UMLJym5ZpBROkCKdSn0ReAmEYISh
lgL2quOtwRpY6XoCe3YsSNKvAmYr0rhHRo3NVmNbhm3ihWQS/uVazYqyEP7tPoLy
w53HaAhnjFpck4LYN7IW0BjQVH6CbOI99rMYWw5NGwqIjlEViujDcvkv27xGc6sZ
h+nSpmlj8s4sV0SNKA9y/Rb1xr9lbJ4jXaSiWS0n67CBu1aKONXDzJUXq55W6swm
KwizKgWcVjTNNHJahznYRw==
`protect END_PROTECTED
