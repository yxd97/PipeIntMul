`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSRaD2BytlftnQUCvHOfPk5pz1+YoYP7PMG+rJoesszrSGeaxus4TuReuR6msth2
/AhIUYDDH1WBTxoaEjhm7Tz2Eph3YZa2Kp2PiXwsFyIRfvOx8EOWWHDXBPzKfhHi
Xk1CcvkuEJ85t9sKxjylieDWoqqgyOarsbU5zrGibkRifapcQzoEhCgECxQp0hGp
YHDvzvf8Xf6o3HHxshzX5tFoK/E2XHDBejihxGAoCPdwSdy7XOJ667zdPWuNfXE9
qJkkZnXdEtMAgY/gyK0Xil7xynjOcqqUvD+MAuTL7OpZusvq1M4/m200kfLp1d84
A3itlU7aRe0EZLXWjYHNG+saOnQSHkkemBw1Qizg6ilxMVut8Tb0VTYR8fo1sZ/V
Rwa08TPYFq+9tNsoXHw3eB4rrTRvawh58nMfspRi+MNOevGPAlnwDG9GAMw0qsZY
l6laT1OTeIiSkwLhhNDa/eKNhZMUEf8rtrxgCViYUtla+PbQJotcsOMGl3Scot68
ZqfgYmcBIT62xX8V6UaRBG/njSpqbrt+2qQ39fyKaLY=
`protect END_PROTECTED
