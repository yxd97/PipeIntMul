`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fc8t1tDkAelUYSj/Uq9w+r3Nl80wM0LenToCAchRQPsU3bz+BfWBa6iipBKtAgI
KSxStS+T5s/9i9I209z5pNU/zC3BpCsHG0QeclFKKwODhkRwVwzmblNeEXSyN1D1
HI0Z2sUpVfbKnZeG+asSsANKgk/uSABdI2gB0QJLzC/hKrAPARp6VCEcyJFpMxrS
4+vQvdK7W9zifE7UO5PfGf1cBCW+1axP5PffXMdm8JGLf8NVIvGuXV1pT9BA+scD
vBK7aokvoT5vKV4/I+Q7D84Bp46VtwALCZi2HAfIQIIwrExzO0/CL26Ph5KouMub
VuLMMDVXmyqmNo/n3KB/uQbwIVwhNppjRlzGlPVNvAKJCnPGzai2DOhucNxZjSIH
81Fm2OVzCurdA7/k2S/Qv4e52odoV2c8e+ReQUzzsUYvbawRc4iJ1yobDVIDyV8D
LZqlObflnLFnWbdVMf8FRG4DmgcuTp3ehsH9jzM2SLZ1nKXRjB5PH9VZM/c2cDg6
Anoq7FvgKS2gvwHhFsNhGg==
`protect END_PROTECTED
