`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1KRBy/IoI6H0tHoA+uAGOx/qYQf5wcADff6KSer78Gb5Op7EzChLDgbF7wmYv7G
MtqLj0EvghPcJXdcY4spkfcPdo9gWnJmRXJPuXg/0f1VgqAM7w82GRaulUJyZkhN
CK2v6hOXl5OAno8UN4Qn9vxy9GCd8KPryIzNwwywU9e8LdZ+aqMW4QYkMJwkXlVA
FRWbkl+24nF81BaR2WySxfaem+4EHys9QWuSdrPe5yl5+awDtLtQF+4TA3EMzWHN
si8c7rJ6v2BigRnOysrfL9NUeyW03b2Jxw7tj9CBNoToJvk2nNgJpwwNy/9s1Dnc
VKUGwRe2f5yvi4BFtKZ5udATXdqlClhOeu4iRR/PnDHeW9dUAQk+rpQXVhVG/bK3
1xozfHSosdW0ck9aCIp4GWknzicLxpfWZ3TTvyOTjKLrL2LdH3Yr3xQdgj8abrLd
ibPlV4v95sOE622b95B2tP+AjB+D6lbJGX4p8Se+9TTsP+xCJvAyUz1aqJgDxaFA
35qLAjmb/Ra4jOJvs1922zIdE4vY7ZJwmWlxv7i/S2dSWCRpIeWyJ/m51PUcAmCw
kamqStZAFUwnWB9JeUGB559Wdy2huFHQv6IrHBkFlBlGHj4W3rHXxxR3QvloOOTo
3CP6T2RrKTV/cqRhc5eGz64Gx5VKLn2xRPHyuAuiDlPXAH9X7ThoEPU1YyBYgR3C
TclGh89wK+CSaKsLs/Ynk6jhgc2IxkHjm8P5JLNi3dl/LqCJOzZ9qY7/x2tnYfMZ
cFCY/Rd2rRAbvtMdAHZcrtmkqlk9SHOZkD2+3AF7vGugYIrtDGlETlhVEYv5hVrS
WQEv22Wma7pv2VFrIZMOcw==
`protect END_PROTECTED
