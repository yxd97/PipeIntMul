`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xtMIpqXqnYrSBxGeX4wDtDmRFTH8dtJjel4Dx8HYuUtcqqA+rC/ez3Et9t7LN5F
yhg5+aCrZBEwQxrghHgoBxQgUSGrVwV8jEGlwnCPi1g+gxEPN2paobqFVD//Qh7x
oDwXHrbNV83nhR1kghcZlkKMZo6fAR8ACU4DObCQqirCDlFXJzif15uUA0flI6qb
a2DzDxlDnrXEDQWBZLfLRs62KqW/Mkw5oLRpqLBfYmFs9HUkRDJBQDbfdW+tDmmI
052I6I4JQyHWX9K0wwlWPM3oDgrMceX7eUHrI7ViqLFZAr0JBDNMkTsFvezdhp4b
FAiXwAo0HojV+t3eMgvfmn8KPWVRAE3g09tf6JGuQmzZSIFHV2qnt+xeGarFI/WK
fCws0GsNxrRHweHMnUZ9b+GFCyE0Eetf0pSe8Cj22Lg9o8LOgdZmjU94KSummZ5t
hRPqXgKajnp1e4sButoiXA==
`protect END_PROTECTED
