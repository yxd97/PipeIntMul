`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OlEQOGUk1HcmgOixLGTfR27nuo0sqfwDtGQBXP+8ktFIiTL45XZ4UN+vp/1Q789f
oPcuRWHuujejr6n01271z8HIwvR9EX+mByk2g8FFOfm4Kh7IsgLj/DIBdtiTLO+I
24q6ZutNBUJEzG8d5+XHrTZ/XZ6OVX8Wvkl68/Z0L57E6QYgHvUIR8N+0dy7w5Cz
EjPEqj+YJWwUyLHasIW06ukKuk2RDjWOrgH+x4EAYjVsYGutsZXYADKzjtjepx1E
XxZf2eLVau4UXGTSp3oUweYdF3ftEGYkAIrpepd8RVpk4IFCu8h9mI9qD1ZjAFYl
vmQhwfA+QCPFlNd/0harQRmzTpJe7OWdW9oFZ5quSS1revFDL6i4AeYWApfU+Kw8
W12TrBif3n+cU6RVZ586nJSGDnfT/h9SN0yu2uxABvqLuQnCoegc/UaQGpKpzcLE
lhf3fyL6sjPNOW/B8Q84kiPk0FIP0y+SUFbVIZLjtkgjQVN30LQldGWI0ili7yFj
WIHpLgta05PqRlJtfmwm+inst3/SAhiQvVVvRdxMYVxJ1CmUdhrZ1H90tjQA9i6V
Ii+1oZcH/DPP22EoG0H1hLO+GXPoQXw3IjGbNuzHD4PmLAa/4WLRgQn/BaLYnVt5
BeLO1CgX/H0nLDMNS8ACn+OqSTiQuOGrJpfooO+fMke5wwS7DF+dr1pE5kpEUEHH
`protect END_PROTECTED
