`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CjD2bmUj58A0LNeD94JmLn6fx5XBBp/6dx8/jfsLooCrJpdR08gbAm7pESApk5a6
aKecye5oaslo5OyLCjRB7erEGScWmrNZIhxFRGaj61QvSbziMrPZl+klem5VlHTN
zyePbKOYdgY39KYW2NaZ3s1cdPi3LroVKmHOrsurfpF2O70jgSPtfeb5efMwktWG
zOEHsh+fXkn2QbTlNjubaYiQNtiXChFVIzH33A3ROWzBmg569C9wQZ6PBz32ccVJ
DxXi97mM7BnNfh89DXbk9gPv4LEx4+6EDDNm6txOBDxsdWtQ1E34TZnXiPgs6f3E
bXPLWNKq0me4Cd1TdyvxIA4jN+ftuPYAyo+cdWLTlmOABLUSXbdhWcwgtoy2lbM3
5lZUAxqHb30r5TVF1apE/Utgd0BDgVLUn9FQNwHGpN+Hiubt4UxJycZnmHAzkrdT
dpYytWXu5/VZF77/JYT6/LqgNKonPgaNhkKhQoGzoWxt8QPG5AW7fy6QDX5ZMhWE
TDAfmErGp2vpYUznCD3tWXNUf0H8Qfm+0WiYOcHyG0N/KxqAFkBgcRPr8orjWtcM
g0HgF9CDzCbMmteYD2s0YQ==
`protect END_PROTECTED
