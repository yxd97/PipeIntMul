`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5aX7lHn3ds9AeIWOhIR5gSozxHPp95q/RwtapLlvwK9gPOcRQD++az4oaTpB7cR7
sD5zdNeQLUpIiatMFU2ZM30zJMA4/l3UwPCzqqA/2W1tv2ZvwIYapgDGTJzBJiYT
ivcFQxqPXFlXJEIKYCWc3CFCUrooR/28JLtkQ8ojr0GQh1JB5YDnokJ2YS9aFIVt
Eabfl7wv4/OU7iWj+IRp8h0HmFPtP73Y4R2GTOxujGFfDvxc5Au+Io02KNN7KLWx
u5Oil+5DUedJ4p+kMTo2E+eJIQKFYuyd6Em+ZXv4bCUgTVH7NKll4hjjssYiD5I2
LAn0Vcg0G8iTsu6HEZr0WzqT4P5UEeo0AZDX0OK+4XZMpr3aQlYHWGFnUCD5EXPj
xxK8HgApjDSsgrBggRF6YDDB3ZtHj+yMNe+27siOkO+uAFB02drtSvBNNA3KMtdX
Uh0PLglaPmCz3iCHZ5D/s3ljbefuSjp300s0RodSGqfktz8bb7Zu/cxY4Bu9mLV9
G1UWgVdA2UWSB4SSR/Jsn/owmpR4Fduj82D1bShdSizdmFJhHYc/efHltkhb6BWe
lp/ymQtQGqldH7VyaF/WPQ7sjDZLJI6kqxjQpeaEGvpUY0AqNpLzLesC9Yb7jwzh
4atSQX87TQwQFBxT8ocwKsu2um20lNFdcDgbLnk/TLkRUBmR4qsB+Ty5RNLtzfya
/bGkbIrcQYgLgrJLXlwOedIb7zK5kkWdX9RoL3IpCdyWzzxdqufOIk57hCBeQLWN
QOeSZnDB6IZiPvsS5U3dMqgZfmDUMHzw+UhmFmzXkMn8PdX2YPA2XvCS8dk9gSbT
TjlAyulDG9DPsbfWXbScD55AzYZavJQ9IXFTFczj2Wh1pSTtZW2nZVptJHQbjN2g
1wibaYns1wgwafYOT7bmxtkwM+ynLU+N0/Wjk9J0mqmoHge3VxHrY1Tp1ywfovbd
oJFrmVR8o1OcKlte4meRTslLn/Kx7SpsbPFKRYOZKA7H/JFm8lG/ixA4L+6tVu3U
Gla7XYDUg2Wl7WvJINgczqxESEmysj9lQDXNluZUIZ5fEn14merN6C2Xt00l9KQb
rVweSGEEXT771jMmvVSbfOHLE9a5QPFGGuBEQ5fxHyEuPn+AnRhonZqXqLl+coaU
ofweBxN798tc1ii6EVHVmSoJIwnpbJ8Qjlv38iGvZgNeBAw3xLFer89r7j+b8fJ6
1QjN3up85JxL5yPGN0PGDldd1L2lOgseJ/5GfAYdxRakevNj8ga3E9nmj418Orkd
9421XTZVr4DiAOCcOnuzt5xO62XOWLtO6kr2cDUQ55iaATxQWIArb10u1zQ6w5XW
u5VZd+WCvqSsSOWiYNyXKGd4L0vTIQTTUcd63SFg3M66NOBK2kHx6b3RamIdufNd
nR0h0BrQmKZ/JtCdYBK6gaQhkoOTHc2SO4CR+w9Lp7C+na7Aa2AqXatPG16WvqXY
w2hGVru58BUi1hbNcfzHrwv5H9QKCK0fJZe2bGfq6IkrREoELR2lA3zUAaJmRRXL
nbTxvcv0u09PZvRwwKYaGBeMjlsOWa1Cp75Sm2tAIuPPLh6noZpLhxQoJrwOK26f
54ap3t84Y9P0xb/SPL0CfZIxMO/EMYWSOvJunVTic/fyiOSoVNr7Wur0YyTDPt69
GtYzry9tKWxCpLUb9UHXs0oXmaFURy4O19xM09kdMBDUGd6mwgK4QUR8x4MP9hmG
S3tCHQ2fKxULOhUGS2veORgOyd0zQ6/emLzofxqjOqwE+mnDmwCY0qH5uiV5d+M/
xP1wQAsT148rTyRnpKot8dk3pRn/u7KLVqIH9oDAWBOS8lcszQvaJuT4OMdKEijs
tPF9O0BRoGdFWDFBADbMjvUnrGQ59K+N2MBo7hbGO50l8cSxA2HrCiVaVUTso8pH
LGh+asodh8QOSQp2yXX0lrD/vUnTgscDRXe0Tl3jQnf1/yESVhJuwkgSJ1KSHRVd
DDGEueobnkmMI+2K/G4WQLH1llsHAepIRVPCckwtxIZimr4VULpXCCZJMUJXSRI9
zolwdV+zEfIiBauzhKx3a/OEDfJVhqtdFdRVasCjE5VUNnSzF5PMUeWCKUdZjQ8Y
Gxp2rDRbsxKmRPwKFC7H5i0YrT6RvGN8X/PEXywo68pacc0IieFAj/IiiVUzRx1x
aRpitH78osRlvTiECRf87MIek0pptuu9kP3BpWXPTF04ejJg93wqiBvK8dt9iPUs
gEZZF/GlUcDpXlJbkZ4d3ptvuigErpr4NvgGVt7emOL2r7wLTXUkHLHloyu06wNT
1moqUXTlJYe1E0/ngvNK/a95V6BiV0wKYsI9njRN6WcW3iVpqGZW+81JiLxyWiXG
uiZEk1r9C7GB+6T7xCh6jlLMm7q+VG9NPH9BS/S1bYfUH61Du5Gsoe1Rvdm+BKat
bGGDBv1lLdLI4pBpWku4rt9TZLpV8xAZFvVH33YrA71XAHIcRhv6Phy7uZtsBUZ3
JBg+/O1l0htZ0+PDXp+qCf1LHu5486DlaOwPAU2P196AiTK4udgTZZQe+2KGbkZM
7S0A43Tf6tNGyLGKSdnx20nBz3crRq4W1ULuRCdQu8r6xUKU1+SLwyPweHnZ7tSP
ZrvYCyOuc0RasBsg0tDbd1yyl1nNKqvLRhUImgCMRlZoeMy+AVhHkgTArs5mysj2
xNiQYW/sZnKFzf6FBAu8/YSQY/Sa4Wy8/a9AyQTkl9wr1qhu+m/4y1YRuYPn9A3i
XeoKgpR/boB6tKKeP9HEceDY4YUZYTlG/nSbio+pscgM5BFxOWLv6SPNSXzDS5dw
A67LGMclit3t6QItOeaqVlYNIlwD62QsCohsUaXwgXrwDdgFi9rRfHf58z3j9Er3
BQZCVZhMNRLschxBQxikA8bXOjiNHbeN6lNeQsHzRFlMO/5vpBRNKCbhWK9feCDM
MDq3zMGYLJA6azWPbHkI4oXjzGGM+r0WPqwzaetXJED1VzCzbw0KBFhV2S+rO+eD
mPe1N+6cKi1qONW/G5iFSdfyI50ayIdyD90QPvEaaLg524JJGp1vsGEt+IA86FVi
hNyMt8UPeL1Co3K2pwsfmF9aag8lys0yOi6GtlEZYQLQ6Kw+6YWPPQB9YxqnaOoG
YFfR4IP2gU8IP85z+gld8vCm17fPhkJETG0IRsaWwuERwMB+eliHZU0BFoCPpPJ3
vXZfdrk/GjWpzpVCzq/RTFZ4agZ4xzQ5pM29OjfK5wbZcb7Qi61dbGS/APjMvGWE
YS+ffd7Q9+hrhehN+0aTWDGU+0Lx+krRvG+GGyGqaq1BcIJlyHbFXn+xW0d8Gyaz
ws9RWqZVujavZDbgeRin3x2c5m0V9rllND6zFBFBscCtOPklz6mT53ny+w6J5nvf
M46IbzlLCE9a0+z0iEYzmciPZcsl02DhDXaTgS36YApM7QCO/Lkx/LF9zH0tKq3S
KymylVMqvpyREH5GYIgWcoer1HR+djfdGXTWbhduWRVYuNopNfeXwO4uYuedGrnF
k/+oPZPv0iFGAnrTT5onNqF3Hjt81KEcBWcwNYhaROBlcb0njLkJPY8T0cgB3ztq
zKR26dLlbpzJQxC6jbqWt4+t82oSiCtNb6JvFKL7W2FbNav3OjfuSiSF/0lrUkbD
ado4QAaVgZTycOA6yfMFRRHh8vhtN1GtBI3U09x9iXf1eGZR1ocx2RAuLEoY5s6d
bZO33fA4hqvHXiJnzJfzK/tpUjlZPOO6YORSn2bmVX3J4q7ZwVxqwo204ubZSPpy
fmcrqFukx92UdElanSP6S9ETDJTIedQv8l9bmi1oACVT7Y0x5T17TjZZsaQFpcu3
iedpxUnI5Hv5zEIm0rG6FSF0LQYliay/0PH8o+3UM0dpkxpAjxT2bqcWxzBo9sq0
R6VApKjTk+gqUMa6zB/jxCFl/My8R8Nmomz/1QG6h2gx+3SJ6QzJX4l0YqJ6xKZZ
bT3oUy2vG9/eTeVUvnVCg4xKIxXKBqKGTGtR0EPo717N6PqHKtC3YIBYB+1p5sUV
bOMAH10G7xduOAUQPRNqSl6qNIGwR0I3codhZYc2M6xPncu6uVtNBm+7W99DjGpS
P1N7UVo4lXPQLwoIPUOQa9hrcUJ7gVJoYOErsFqhc4t21hrjGqQTM0zQ+uK3tJEp
IPJFVIB/PaFhZnix5xkcVeWzHUm24+0FooRG99suKm98GqMaZP3+eOJ1q1khyP1F
SCvZW/Gkq1XDMgHhnq1nUosh5ocq8Owd8QRM7uzW5leEhepjJ36phmqryq29FSbJ
q0SEou6C6zpvjAsFyglhF9pywj9vdGPEhSxV4PCtJMMKaqQOU1G5wzLu+ORHA4Jp
scNXs/768U4V9cf+KxcvpJhb6GgfdDdMuMSTqXj5NmDV+QSXrvYoZRIwmDHt91jZ
zmjArBhc8fpLw66nElPFBdHT5aKi+NYmGuUzqauXuJronKLDhvCtKBGSkMciarkD
r9hBn2tcrUd94uQad9uEA4er8tZoR9fEowPcCWpIXCDuEZ83MHf2DaGfb2I9xiku
hiMsduhgNMxAVo/Keleu+hQ67YAtWRJwFjECWUYcr0BHLlfSNF6eoLGHejGoj5Zc
TV7pmJxdug8uYuqFb98Ti/NKzBFSpHff6sjNEelwzBeRnzl5uBBb3Kd2tg9TpFdD
Lg/msnNniLoFZo1xQjFHWp5Nd0nScg7Spam4khrilZdC+rbdweTA91K9toxMCCRZ
SKnxf4fWGkYLF1K/BpPtJjhzRfeB30+0fQPwqMPgWUBDJRT2PJ2JXX394pTEe4x6
BKwAAi6mkKpOzCqn4F56QqMdnXnKkfo0N8a9UpJNX1WSR7wCtednGbrGaXvBxB8n
I1q+5lvaSE9tYbb2S9DAh3b8BMyy0/vUVMc5vnnbXfwOJ+MM9naP5BeXE4WXpeCj
IiZ3WYt1kKrG1slWjmIoVmL31dxVxvsT9zNfTep3+7gXRumED+0bUiD1I9tZ8ZSI
r92JHqmnI+dq6WEumIFBAux+bLHS+5NsDCb+uVjBNKtcHI0lNG2HylIpl6d9vEND
z/CKYhB8PCBJoEcfltkQTA==
`protect END_PROTECTED
