`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ORUA8u9giYxNVOuzBPWmYU66o24NsT79J54MK5KmmipY8u9EHMPG+1Cr4efc2hAf
WR5uNhyc8GlsmaMAudQM5PQJ1ItuZOOQCmTWF9Oml/1r75p4prV9+0Df7wX9M5u8
ouQWgZo9Dh/DsUoRLKW5J+SkNHwxconSHGKwDrAJNGaKcFS7IHwF56d7Dde+aCf1
zgRUptZNG2N+CdxJipA6CAunYGS5v3a2i1pbdRepZoVbf8bSIGcMFiOJWUeksW0d
96F5VGHGS+Bqf/MqxbVSDi0febfELv/xcxZ0mUhRvyrIatnjmK1/wrNY02jfE5/8
FPVef/CZhVuyPnqaX0NH0Wzc9904l2r40Sqj9t8vWlpWTDAgpjeWzJbIvNX8SJmC
mI6130el0Yn4yryzaz3cPSU49wSzkg/yJkXBx2osOFzIvCTBjWzHlxbk3BCpHSe4
HKbDvhMM6HMsHCh/EXYQHdsa02fH3IFn7KYc988A2+6IiEbGaedHStC5HbUF0lIj
doHlDYBcPiisZOGi5PZUnL7LpcrepXNojXSRHFXqAyr5/vUFDTaolIiIbm7O9UY6
HlZGWGfaywSbJsF0BrMpbmNKEb2jKISVGVkmLWli/UCjXNtQ8VZWAZ4yeSAeBf41
nchz/9+MCcVUNlddWHx8/JKl8Dubb5Tl8txDXrt9o4oAdWely7qeNKWF1dUzSQP9
1Tt5D7B/BG3UfBkOn0K5bk8sgSfH4hNncOXZTzyj83mGAM2kNxkPPl412273aSJv
KmENmiqB6mpIQXJYDY+fU6HV68AMxXvr2m1pFJLZrHobtb4FUx5Itzh7F6Umx3Lu
DctN7DbuibNii7bCLCdHSJHDaNNuZgYyDpUDm5LxKc6ynxSJ7VU0I3PS9D+sEHu9
DutpEN3wc8lnUfLkJBNUwpsWlgZ+doS50UIa63K6jPYPz/fBlEy7rTZI+6Zf+6uJ
ajRih9Kr40dJYvJD35iwFvy9tm/9r491x5I2gDkgg5qGMdFPFVeSBtuafFSrV4Zp
vqwFUDaLY9Gf2l669CQC1yT2jS0dVn0yThnjY6rsU4ck+yHoDZ3VPjUHDNIzWbNc
85JFnHYpBcV5j0yDKCz9u9EtkyPLXpxClgRyRwxn/VxkQduzQj6WEiRhdJ+tm6qA
6OwyrILNvHu/iDMlE6lRE1t9FHh4UUKLHyxClQ8kxBPG7sAUtYHUsKhvVdviYi4y
HBe1Eoj/1xf1hLc1O9d9woI+N1TJ8gloDFskjLJLairj3yhYGsNdQAcPyBVuL1jz
pUPdZ/tZ7cpU3975Folt2hoOI1hxhrBV1l/R2SDLdBvrxLoEo4GXeh9FxA6+oC4a
I/TFl9I8cX+HQ3uIC23d/Z1cXz+RjmgOcwXZykV1rc8Vi4pyMUmUDCMog8cTCPUI
rrlsHR270tM1YobYSsCJVZUVldiMZuC00p62jmAOgoKa7E2SAxc6RbkpjmmtVHaZ
weAet5F9GC7qeyKKcCp2qQh4fLoMVV0fwvTT610Ce98OKo9Foa3fQPnLXm1Tc5Re
xRI1BqB/FEvH0+Cgu+9X51NoDZqYutL49AZKJWbGyuzBZmPC53zrpZieXXgrnGLi
YXvnvhFBFEnXE/kCW1hACrnG+KkeXRor3JBEaD5wmJSvvnnIiEKjx/n3y0L/ABCL
4h4RV1bVclBTFqzZ+DuJrMSqWOLFYEMVzU7f1zxf4L1NHoE+DDYOpD8/09LTeXF0
uZkYFCut7AQhI+nRBXRgWU5AGo553WEG1H372nktJk/HxNTASevNzn0BVS8trW9Q
eSyd0pJyzm8F8Kecn25+7dyTlUa5kHQMdjlVNkydxfqGInczGB4gTRm6gNigyWqZ
2MlbLf7fr7LEfWqFSlwsYmudrya3X/t3r4mFk6JcoPLhIwrY6mD7e+Q3A8BY9DP6
J2aTJrT9JNBE3rgk5wu0B8TLzlK3Yr1wzCXOUYpmtOiLSHaUnNHmmqzO15kT6cJC
/Vq/KJTUcDHlJbBYKlmmsx0dM+nIaTLE3+uw/57wbeeewtc8MDgJHgVTdqVpxuHL
h9KPeXNyN5RV4VpIMgW9ngPTL3dWW2hEWV/UkgJXQt2ChQbgnieA0l5+J9ffROEz
QEuSrLbPMk/6P2OWt/luZBhJO22/VMxWYbA5q4Hf2lid8nc4qBZXb9z9XP8A8ZIF
L4QBAYWvv4DYUE6GsCLCzbzG02UjiBfMZUZsEVFJt2xL98EDrQv8hBjVDSSDef6z
rviKQsxC0H5nc1IPPPViHWCjlD7Ey7aebi1QCElSMBniE2m3P93g7yqo4mjcUKrA
iPfRMFX15zZYDcRD0JRDmQZJ2E4NQeqqhiLNJ0HBk5wd4wvVJBosjp42yEfsY8JW
lY+TtRy97dN9FO/VdT7nHuq63M63v0BqOTAIMR8KYeUo4WS7vONpHCa3lCOyX9nU
V/4NqKeCsIqIjVB1aDt0N0CE5zE2LHlXNqDZcT8WbYau/AZY8a8n5OQpzzpix6ii
HsQ9tg3LKiyuWdMu1UPxy4v6aHao4mGf71GmcZRFi262OaSmimXBejiScwHBP5ZJ
jK4bisoHUdWmfu5+VglRByWsu2Gc4s8FMa8Ljm7+/0AqoMOgujEN3aRI7/rIkMBL
QqW8S0cLfqKo9zlV85hf0hgkYrjPMoLcRFs+qowkFxOBB2YllnmWqZECIN1O3/qV
31b7gGMxEzgzYpFzidyAWu4yZLebMZSEvgDj+2JJQEDJOxYSH6oXdG3g1g8ztLVp
utMTckuc9QRyd4g7S3zp5R/JfMManLhY9b/FdaMMhWotgnoXMNBanpzge6tjtj7s
4J8qYgJ9TeHxoFQOR61VRsIOwZVwyl9je9oMWjoDWNPCe19tVrkYGZ/R19e0EcUt
O1wZz27DJAv1tPVXTS6g43YlegASHa6R+m5/KUYOQRDUHEJTGjtkNiL+1p7oTX1b
1EF+uo9zRla07FU4HjumBSTUfzquMEMRmrJge1yR0syL2PvCpllqXdxIXbbyRt9d
5rfdjxS0p7i+W1cu64jZQ73g5cPm3wvROSVAB4SJzeZC7KQDGK72NCEScjarOV+r
a31JFA1rNq97Rd+pX7T6v8X2A2hD4duVN4T3rqMyLRxuwGgqVBQR4756Lz5Vkqeb
S1p0XJaOOwtdAIqiaRHhkIY1MlndZ/LXf9sp9pQyr/BvNFd0t+VRQAu9nSnAgFyr
114tv9l4vJfam8oHj/3u77Vy+3FaaoeudCoruIN6mUpjYLatpgcwwakrkumZqD0Z
bfe3e6F2Nl7uyokNi5D72dU0rE0IOOYvL2kazE7ek4HFDevZFtBbf9Md8KDSZ0BH
+gZDegUe04+NasVfr8860TyHQCrIiLvmLX/g5WL9Cso=
`protect END_PROTECTED
