`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6WsKSJ9M7RbanQj850s8i1ZNigJy9CJall1jovRW6J1KAA2loTak4oP30UsXfWjE
eu72SvAmTddG/Hv0FFUJ9lSw8x9++5cX9B+5eGIVVq4tkdbwzLgEbCx9qvxZ3utq
jXCngJ6aFIO7rUPZyrbOJuH0aHNLq2PDXCnkRkqKhMEHIfI1tZHzbD9lDPjG2Tve
t8f2RWGOEHyXz4BEFymd4y9MM2yimEcyo0AgUephDIyajb3vxFBLWkyI0paUa3gx
ToBL8AqvYV+uNXd5c8NmVUTFjU6yscDOTg3JU5UHf+o=
`protect END_PROTECTED
