`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VBU2DM0YxV09BC+Ai7t4WRx9VIcwUI4TpW1yx6x1GsQ5YLdFi9G0M8fIF31EIZYM
Jrm+iyPr2DsWajMEaXkVYLDpGty1aNnunT+iktol3KLwDMSVZAc6XXUFHK7z4Qll
OuLvu21cixDRnM9mD4w13usPpyNEB3XPe2kUbX7/HoKM1b6/+Hgof1PKFRuqlL4n
+PPM0Mzngn9PCfMm6hp+/V850nQCzHuNOhIXwnqin3+pAVMvOjeuUilL16Rcp6/m
K7p7onYWxtO//jlJX+ZWkaEbbKrPSuvuTy6E0ivyvYzoQzrGCeRCmJS4PzCN6gRV
U6Xq4KquORYNKyJStJTlwM3q8J/6sCDzglMYxywWeQ8cRHccS9iC/7A/nvT4IW7L
+LERymAnlYUvRSXuM01XTQ==
`protect END_PROTECTED
