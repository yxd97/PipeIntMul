`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c1XH4Sarp1wpMt/8YxypyD/DJHAzfrABYKIl2GXzMkywRsHcvIIL4MdfMeuwVlr/
oo4m6zNqMUH8cGZ70SwmigFaL0M7lo6D9AKhQDLCjGu9QeATM12sIaI8q+rgP+9z
rSt6H+E+6NFVek181jBTN6jPrjlEe5UawUfN376zc+lHBjvlkI350yK1X9hEsJ5z
MvkVmMTWPwsMW1h+FBfX2gm14WjDsPeP97pWKN6rkVz6wEg687qZEmC1VeAp2c7b
6IvV+3QVtxQKFVTDpVWi/+WK4xXy4nz9LkKZJCnZgCAb/t70YZgwlDNaNgEH+hsl
sfuPC986BnrMx8Jb9Jkf6xDlceg7Jha+Dk2wdx4W/TXQbxQAJq+6N+sIPzE7cvwq
Bpt2LpSUiyf8YwSHD+gUrA==
`protect END_PROTECTED
