`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XTLDmcjqhCv2erjqVZGMw1rxqK3iUgVizngxmLPPO9KoFHlYbuR9NUvhRIHOS1h
oILKctlN9vJG7sR3VAA1O28wZvbStCQHLrnn0KRpneb3sofZQo0hH8cy+vWsVnF0
gVf4D4uNNix4WqAkBlO8mCPJeas2XwLhNV3+E9RcSC1YZu/0tgg6br45zHseTp0k
MPY3Uhuv/ZvbywiZQriZE0Xyee+4xBxOM5UidSUrvB03eCmDiQ3KUPqt0Gr2Jvw7
iGB91zevJOk8f1DamusXQsM+L6uGHOt952wMoiwURscPjZutHUEBBYKdZR14pZkW
`protect END_PROTECTED
