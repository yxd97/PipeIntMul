`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8eiSgS1XqLrBfgJZUTshPWtSAlEHe+fn989+EJTsciEj0KgcrYwgIJDyrdx7bmIy
BbK7cQNEk7ESEuxXbu7WlmkaRGI35bq+f2DKXNGx7U+uuSwEki/6PvuneEdqfFeL
cDmKAYOpbO91fGCSvZ2pYppxNdmlhUQ7PKZnlOdnsiuKMVQSAZmJ/UKaA2zpviPL
1NhitNxcbM7GkfCTQ8yJ8R9pVhe/vaxsas26omFTi4PPWeUM4JQJoywCDKLbWKDY
J7dFVv4ni0n9pt5h1vd7nkJSx4rmAkHue4DGv6JodDmA5lyTykXmmP121eKkNL1h
t8a5lIjti8AUBxiJcK0HiNfbSCfuhU6TK+V/2ozphvQ5dV7aYUCrEsT79q4xvBLv
qHzuEsqXv7Toa1fCzC5X+QwaDlzhekv3Uca0dKtchSm7wUfY2ftONx0otJpJpMbh
v0zWjVeMCjVYzD/zJFncWmcYYgNs6Xx+kCykQMxFs/Pc6XRw9E6w152K1JYlJ4bc
0633TndWaDuO9hw0J+6Gyckjy7weEBGJFGXOostVfxVFm0J6SToC8cvPjhpLLCXo
ybHgxVvlQ8jaDfYtseEXWCOhFaBq6k+IGlctyaf3fRVKftaRsVttIAxULY5s4u0n
zBETvxoX64Fmbwrj5+kj5j0IJ78B6gEdFEtv6KQ3kec=
`protect END_PROTECTED
