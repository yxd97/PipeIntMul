`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKXa/49emdNOV3+vOg4DWUGvS21rpb+K5FRxB06q7+YHUx0RqxhmHFMhpOW4dA1d
8inFVxC2GuoLb3+1n6kwTUEPlmn2MmQRQDUOhVeFm8v6eULWkz9rN0/VvaWF3fsH
KcK9mICYqkLso5m61qdW/jOMghX/shfkn4HXfVt48T6MaB2BA09vtkMI43FRgrlS
Hb5hVS9q+iljysNjDI5MY6VCQx0EPIz/yXfxS25IQqEr3YbUb0jE0TRRcwuj3cgT
KPrh2e4SfVUroOCL2JkwQFJc1Xmnzouw9AZBhb8JXRdk71ZQYHbZuPWufx/CihsQ
Z0gYBELtCwC7PFi+bquPzHPwrxCf+eUSHNlnxUIenJok9fYcyjO1Nyc6FD3863yO
STJzIx41STWF03oji1SHpgAVf5V6MzCK3A4/ZZit0nZy0wclVAbVEmZlP3udMjwO
KnByAjdMU+akWQq/GYnQ4ErZgs/GCfsUjr/eF8YL6QP3jXMmPhsc99cLdj15mdRH
Vw5XrqqGiy7j66SIWjNrx00U8LZfFGs5u6GQOxmIhVcRdnCUONTfhLa1MD/SkaSV
JhINnV9l7PxPUGG3wFI0dTBZT2FdQg1y+p4p2RmVc5KFlrGQgYPABcYudIaWbh0W
VXS+mHvdmp5hVP0sfpX2mIOQsWw/JlRrWqAC8hDTwNTQu4aMXVKnXiud4f/UcTTP
`protect END_PROTECTED
