`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mH0RWEKzUyOBAuU1/0ph4VtQij5aJHefTKCw2ayl/nIHexhxMWBjPCvmO9mtBBWn
P4iAeOhYi+SyVUXo+DRjYBywzjE1g70FGZTO0rcQsaPJGND2OdzV4uSskEzc98Qy
7JgZBjNDaDAWYWfZguUs9qScH+wCuHoYmvQyB5UaL7THlpB7AEkc+dbbNe41jIoa
81eUP1zQvYhWig84NJfrS/1o051c2b1683pYOeAgJfCoy0blHALXDHa4Q9u+EFKO
m+ab/9eqzbkSCkc3jZACSV85mAdrWzQjE9rw0PCDEa9USFX6UHDNZSE5Vn1yrkQF
UwcyXAAeqvG8uh/5GoZhiQriPPc1vRSj1copiQMoAJzckdH5oG21K9ppTVyh7tJA
x3w/wcx/Up2Kv+rW2p4OjYVYnPdQICi9Q5WNKRKs7/+rY9vyWD9z9HlPgON3iE8k
IIpRgeLRXyQiLsenpDTOqq7mQKPqkZXRSgIXejYepjTcHrhbxP2oESmysgdvOxht
KgUjLZBCBA3Wy1Pb6i14CN4t4o4BniDkCbRu4dVd7BKIJd4JsPXSyPWsZBq29him
VuPwtVbIRNBXqT2DwCx/U50jKAyo2VvFgRKE/O4x6hK43UKZSl50m/fKWEYAN70a
tQvxIWNkYsKozHRSV3PLRNnd1mHzdyO9Ny9DtvXeASt243ZRk8NREKYIeoHnMIPq
Tl1opIc6JQE5mV+2P0wzTK0C/77xnibzynLiTHqVpJEjLlWI+tUaTasdkCsJRkz3
AyAyes+vnY7Rb2e5OkeAImUB0N4CvGJWbdoXmpk8jxhc2UR7rNKVwUtiZ2S93K/t
EGLLH8jiX+CHienAiuTafph5WUtzQo3q97hiN72YBc92tfr5yP3FUtl+5d0I80o+
bYCMOU3KxxbWVIN+Xv+5WTwIMW8lq5W0T60bWkxstEJtqU7rJ3jeqaXoDytm60UV
rgDEAr6p6EF771b3cox34D6BSmbRThTxxvTQTn1IvmLnQJH64wccnY1pD0AP5x01
Lw1vki8o5cO+eXA8DdGF0A==
`protect END_PROTECTED
