`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/knBGIP1/MqS1DmcfLqYfZD1YS9w0ImSikUPSEtdO3BEsIqjgrs6jVx0BkDEuus
ad/FF4yKu9IXbvLpwghRBtQmOsmP4oUWuqbE2NQgNuWL9qfgUSan2RAxtEA7IQnS
rcqb0zlB+AK4NceY8Qf6zrkZ0QckeVSNDJpSSfbSBFW8w84pBiTufDbvhKUu54G6
A3C5g9sFTDDGhXhdtRI0Yt437Oo3mXuVcTjjwiaDmVMrus5Xbz4na3w2UDEgUGYs
WEK8lUUBDVEAkALdkAbN1u2C8OjRLyI8Ir8wX10CFOsH1gkDRc/OnuQEkOvDWn+7
g42Bycx4iYGduG/B0gyQiYL2QvB7j8fPCvkSQJojJygkSg8gKjnU72yC3sQYgieT
3aZeNHnhyPGZw9QkP53vUQ==
`protect END_PROTECTED
