`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DuPdVFX87TjN9YemHRMEAHWUhbYm6gyA/RevbD1SyHd60guOjmfDe1f7Pud997Zk
xeiEJKmmsjyAw8W15PpDCdieb1YTH4wikoIWORdP70xhYcEIHAIk3IIUyYt5PXbK
VR2SmSat1VnXhVmnKfF+n1hByXWtJCsjh6RDoz9UbfczvsfF+ZpdVMbFWXR3+Fbp
et9bk0kUbvfM0QX2SvvQfuDUlZzxfJ5bf6+BwXfPuelyQtKE7ACAyCykdznY6SCl
fN3GYRE/B8z14yPvq+OaSscnhNw+3HV/hLcCto3VVLzDBBfvq/vrlPMiPGVE5Tfd
YVT12yk2SyNneUGDUamN/7EH1VHp7Ysw71TfcGkdmTW2sepvL/vgmd+EdoBEf5iq
Nwipu8aQu2SdWREM+yTEqA==
`protect END_PROTECTED
