`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KbgPyJLmYWX0ik/lvyTm5cAWF4Rvhp3ouyZ7wUMWIwWwVc9MQQAndszPIimRHxB3
fHUEK/h00a4fnr1VzH2RsgFGXhQvEjHpjk1UfYhnwc2cV04bjYRN6DaRrbwonDih
cS6qBsGPvlQUDQxPftDU+NSkf3qC3hsM0OajmBgXAsFqTUkT2pytI3308KaDRJ8p
W8Xs8LIsVvLKuu2PjeHar0SE45tMpyC3pgzxoTm882XhfuYQD+TOmsRPo7W+SKjm
XpBFvRruY35tXkUTcbipxQEM+6e4GjOrp1QmtjgBCQU80VAc4zRlyciToLvPzliI
4HQxSFynmxxeQ627p3yU9NS54srEPh59ixrQ4+xRREZU1WeM/aZ3Jky/Ai4Ro3YY
M2fme65cl7Dms2AUUTctlg==
`protect END_PROTECTED
