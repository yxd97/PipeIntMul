`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXBDP1LH8EnRTwIu8e9tl/HvN8UF4mjA3f2tMn3jHcB0o0y1sOJPAYX66kZJ+H9p
/J0NRJkqC/6ZL/oDDf9/OvEXRJmMZ1W8frA+GtVs6lGAyJv5aKITCzjCWqrfEb/M
hazieaWfBC+vKFrC1uOhyv8e9VvKk1HcMaPX+ZGZe8jqj8bgMmjBFxJ/LxVjHuBQ
TnnPmuywc/OTCN6xZxcmZE/nEAKk8gmMSINhKxXLqFtPZ50PDpR02CqVnH6nAp1A
u8DNaLxSPxT1OFZq3RitYYCDpfB/8/851Wwpb5OkOZiXe45Keu2dKV86Vvj+acmH
6/B3L+ndWwssziO43m25kVQDvts+PC99ov1x8rdApHSKz0nytjlysB4aHUmWbaoW
s6KmOxaQ0GYr00c+ySq6ypd2g8YqXlG/9dxBwCvgx4mCnHfChLyFKLZ/cJOdhz1a
Ex2fYhFxLwVle1XCfTCKhmLdgB7INtv9vpGrKSSVDhJyS5EHs/Zgbyuyj7nACNg9
v8bzm9ahiqd7WMLm47mlwm5RKBK2GEFTNfm1lX4sAbA16fCP92GlvlJ1UogRn+HB
oQlm5Z+9xjSUUEPXKpVMcr9N8f+VqX3oZZkBR8xWyQsVJ/mPxmlBKjxLzMNCnbDk
xV0ZYPuRP9juRdCU9h0GDeIDKpVf0tSWK8pzMiygGwJI6wTf/x741u8vf/2EpMJw
O5zdNOeohBNcWiHwiyJUKNwv++VNASsruNBbQP1nDL/Xnsly2P9ELs3prQcuM8q1
6ESqqICk+L6QRIh9xzCikTKLVGuMO07QQj2MYi0ZwYxe+kdOSZnUB73eYusRVqT9
finVdcFGeoDlhUX58ijFK0hxrf7BFb3BV3YkqPT7NuLDzw/NxKi+Ak7kX1LohIdR
+7Njjy153ixG8egc4N55msWs149+gZuu9s98um1Qibn5BmmofEVQusjEdmfa0p4N
WaP10o2D8AqS6FJ5zYvfq8aCs4QeTh7mJ42e8LXBZr7qbrEear6VRMapRes5Lo2E
CBONatN0eKF4+GM05YCCBgTOvxGRwvz81FA9Q7T8KdrytczAcRWuF6CsV6N3K0Am
DKFUnV716+QG2+lJmCkQmshKhUhqf8/R+M6H+qRfHbOrCwAnbhKF3seP4+BPekAu
E6SpiZs9Jfoz9+CwTXG/BuRy2s+hwUOGGyw1vVspz/Nrl0tIdeiGvQL7Ul5QE/oJ
55Qs9uDmhtFleVqWUuGJOZonxIyMtGPlAsMscflhFdWdzqiXLwmq9XJqwbdL4Vvp
W8gw+W2CwhmsSBunxKS/+h//0n7oxqdYll9KFeIKvMN+19GrbvMVY1IU6npQsUm3
zzR++Yr9032fV7Tgu5yhnlVQtj6qGnI7BasSPY3SIw3SnjnX/ietmSvPBY89FcY9
R6n5ULKUE8+f17H1VCS4oTwa3TtQc84Q6cfE7XeWLMOwsF1MBhshVGoKh87kEQIY
anlHkquWsjkmUCZ7gZ2KG0ZdDhGcBDz3Qxs/ZOSJmLBwlzuJ1U61wMn7OchYy89Y
FuYWE3Ju2GPb+GA8K02se0MoHn4o+cBkMjlOUJ/ByCpygf8abp6OjWPZ1C5k3+Xn
NBNqMFKkfv08/rZDZaCmvn8VEHGi6+Ge5FLHNAS8WfgDvU7PflYDH2LOYKGxmsSW
BJe2shdRChCtUUQ3emlDApiBEIcoO13JuggzPs9it4bk3+Yks25JyIRoflQHKHGJ
JpugbeJh9CR7qhq4nnI5b0P/F9bmP/yywA1ov5VR02ITG7Zfd+GpeRMMtTRs9Jpv
1K6l70wln1wnf5OGwrqvY1qARec1R6iigfhvwXXSS+vwYupbSYBzoSQ+2/NLARJy
Ar+GBDffSFV8Kt7nAo9I86T3saUDqZVmazKZ+Hzk5W2dBdQe++lYCbK1rmDvkDS4
/PzEo48Wbiq8ynAx3b/bWNMwBaOHGkLgeRH4hk6bDWxVl7FvRCypsS/eF0qFE91o
MMVBkq0nlsYotdw3Cz0i+0R/KIhPp6yQJZylTniI5pJuYA4RJYxZJY3dBkgYgQh+
j6Xm9M3qNsmMvK7Ib8fDExs/yUWnRI6smcy1THhWr5ei4mwHUIkK5nsXfpVgsnRe
wzwzGghfz4JGhpDQX3SxlhzvghAM8fpJekCU6oOpPTNldtfd6Jc0VaPC9Sna41io
iEDeBo6vY1QR60UHSuaIfoWFY5ezkIoJsuWvdqo370RDpchZousSweueEO9NbMrH
FH2Wz7WbFWoR2x7x7C+bP42hDdJ6L94orUJt3Cx233jq3fVVh1l0IRW19xI3Pltj
pl1DNsbMvyP1jZt2YdErQ1SkJJdSTq8/yIdye2ZKVUawH/nJ27JhZT4AXyWtFp4Q
khsmBEhMwDFgO8oM/9Lzw8TWSoc5WBWeefrY0t2jCUtaOPCvOx/EQNHN5SbhRlA2
EgEqkAlKlHQTn83hj+1Wc/9d6hedj2+VX/e0ELbRyzKyZzhKANrKK2FtkEoGD88w
BRXWcZY21sLUzgiODk/5khCrR19g8UWZoUEQOPdJ68BXVBZSWgkxaNgoCOoIAh++
mVECQPa2u87b+cT0ESExj0mmfhTzbWekuye3nbXxuld1j1gQiOgZVzhOMMw/d8er
Rttme5upxxUj9cI6SOp7uXElXqFETY/jAKQ6sOukI57deSX8/sHNvcl8qFqwgsZo
6zse5P7BI1kglTpBvh2jt6IH5gCZxER86F/vUQWc0lps9ph8lPOIvsqKZpXLwDGu
bhe5a89JkAXl2YgtSAgKUwDS2z0lhbPXv0B3eiqinxoY+jj1dibk4OOygJpcigBc
JCOtnIJsKaQvLEVwvfyg9XkMOIvyIJ55pJjCPAqOQLI=
`protect END_PROTECTED
