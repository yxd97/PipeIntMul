`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FnnQ4orcyZbxUpgP3m3ZJpLNs6c2CUleZDjkuvIIt0U33eEOGJyp6dgrksVR+7cm
/Y1JKPFGH0ax6BRkVe+OYYs9mas8caH9TjHRdwBxg84V7oLPNGvXQzd13/yHwwh3
m3uFHB+AmlJpcToXMxAjq3Tc6cCOg7eO8SzPp9iC/NXXao/UmCllqk74h/b1QThZ
p6Zw9xlY3D76U1U23MruN4y066hO2hwFZr9mzDnX1wnpVJMW/rXiei2q+CI/L+e4
y8Bly4TsWoYTpGqMqqZJ87HE7DQYCZDhkjHFwTAGUPV2l4IhNkmj/idRwjeiSRkw
6CdYUBh2c3aZ8c7aWeSolAT0Z+z3k32nPMkF3a00EmfKtGTJIkl+sYHoQazGEgcf
o7PacUfgH37QONyhnxrlOsreHLVCVAgGWFH/Blw87shgOd4lR/6OFWyrv5AsUPVg
nOyMqVIUB6pnlzyBguv6e6UdYH/i2fxNcAseoPfCfEvSiTZZoTltqFCA4QwEgocN
r/OeGDc8UGTs0eVI2tXjgGFKscEXQpxshEGqU/tSH2fEYE7BWPHsWPnr9+yl/svt
5W4hS1lv0K9pVZWU3tn21A==
`protect END_PROTECTED
