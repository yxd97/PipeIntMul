`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V8RXLdXX8CxTk24wrzmdJJ/6eZsg6blO8Drzwf8IRUk9y65z1prbAwjF83wHZAuz
CxTKoYzuq0u6xRPwDjtNshh2FnKtgQbmicb2nAbvPU/H01i8vrGYcWYUkefOAkSS
nCOzR+2+JvQFlbBUIE8E3usrMsGq+nhrHv2JYa11zSsfgl3nvxK9bOx7dRxdh68C
DvrIBlOMnRKBOyGFOvAxihOXV0ISB/mfUTDzxjPXf/Hl1sfepQX6OQDPLzaSKjEZ
6V3rQEjnUbTntxwBHuTReWfjTJ4DZkvD8EbUUTi0CC8q6SiGuywi+olMmW7rN5RH
CwoRrJ6IzEhQ23IpyNiYRxu5C5vCDXhCoEydAS9B7IKjaKr6onzoZSRUaKXE5WOR
ce4RdBeOZQ/PzuIVZsvE4yiHfx3N+1/Grmb2z942/ShylOODYV9h6bXZI7apHfBm
2DnFQGJ5CUP16oc3h0U8AySEqPijuKM6UZaJoTmYwK4Miy4FnhLcFfuQUu57MhkT
Guxz4sHkNtiG646Y44z52Q==
`protect END_PROTECTED
