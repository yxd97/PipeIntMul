`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIfyjrmjqJ7OJQAS5zn/fzqxOZVlG023Pg9bFJuSex2Aq0aCgvUDQjBySJfhJnqg
xjeBCiGVZamFj4th1sf8ZSNlVe2RI7kBEzagw1yDSSv0Uk0zNDWpYbJs9Q8v3lJ4
KKhIX31oXGtVHuP9dBn8dDeUNcUWBpnWKfX+fbebaYLA+VMIoyzPt3jUxtlOBOry
ZSuZ34VwZZCo8xhMOEGYVmU/ozvFxZTbOCppBjpnyPOmu5q3AmgrjfuZs+vn6CKV
oLIhpcCyIxS2IV2aF1jg4g==
`protect END_PROTECTED
