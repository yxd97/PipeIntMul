`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yofuvbCUHE/nrA7z55sSa2Z0Vte9Xfo4gDgPMCWqNBowfneqPpffsuowNfz1/W4o
58gnS42NCtMLT5SSwqbIEGSM9i8RdzJfBXu3W3qoaq98IswpLjTwrgHgrZMcUelv
J+byTwN8iirr9eSBr7wSj00StQkA3gYhakj3tMBc3yP2VxjqqNoU7u8n0uWbhJhz
fcCUWIeNGGCfH5oDRIkshFCOPyC3CtwaDmpbUPWaYeCXeA8K4eJzplebQxbIYFLe
G1R2HKl+odih2qDVyE13VcFduQvitchk2YfMGHJhOaxG3JMn2R7SBfEyRMNMWPFw
l48SLv0sCj/WY3kM+mpeCvIFZ9Q8YnkIZilZIZOecpv+G9nS1ITyCeuqZXMCNYSg
`protect END_PROTECTED
