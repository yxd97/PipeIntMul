`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fCYuH+F6Mv06nbcm7pk6CyCnRq0I+gK9ryT70niuHeefnQPgYV5gwxn1ZETC8r/T
2DIy2H4pcxcNprL4DESky0MaXqaw+xCQBxa86L6ojs8Ry4YROeI0d54xZhOprAgO
2Hpopk3mEj8/XA2vPKzhxN8ST4GGlx1cEn57UENFIc1k9lMymoWY2ta1N3B/ry1a
Qtx01QD5/3qvs1lnV10487A4l5xHM3NoMibgwP9oSnXGBD9LWzkMbhD4ZAuaIK7u
FTctJFLa6E7c1aOiCFLEMJP75671oBtQRT/cBBisbvwOv9wzrDKVKOJaijAQZRPp
eolKIZsriRj4U5b5kBjr4nvMqAieMPJowOn0o7cohiI509EbdbUkX+V8NXB9+VGX
/Ex9Ot2VzmfVnLUTSgSNUm5lhGIlHIBt86dyQtDF2PklF4C5Czh65eSL75WGGuiP
d+P3uas8nB/VUcS40oD9MQc52CMcMvgUnqiQBb/DcaYMgqZhV8ZbWZkWh4362qFm
cJKrlpTAv4ccSb04wLWBheoqllfFKAoiXWKk0X9FiDmPf6e/puj8THOe7BgqMn7i
6IsKTM9jM4i5bSAqtAbCl0KD7FRpWkT2GElUklSV4nLY9I0jF+Vt1Y2HmABXrAyK
t6gBAM3+XabbaYg0nbb7NCZqqZvrsZ3o1VQF527m8AA8HbN2bG3jOEUCjuHn7tEQ
2hOvih19uNEwS8vdAC2Ft/SxedyrPeh9FhnppOwBedavviABpUqgWf35o5Rwa+D8
H9CXCkgmIelAk46aJtDsEY/T5fb2O80nyl7CGCcjFjD1DdcIQEZpgZFD9Az0L+dY
kWznm4rIUr1vsCWd38eZ8eYT8Lebn+MNObYLD2C2NhY=
`protect END_PROTECTED
