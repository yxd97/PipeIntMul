`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1MxsoBlDm5LNdeigy5MHB8Fb/55sTIvPALmaQVTS2wrN6FHM2W/+wGJpql975/0M
GywcoEOjNMKHhVAIfsnXgEBy/sfC1ewBDLEHu9RtDkMwa2YinMwfG3j01Kq3lLCp
t9dE/T/C/O6q5siWhE2/oMa0NIJkKG8PvmQoBB8xrBcHb0rUJDPMjYEGyD/z5EBd
Vo5gZBA0ZICJvGAclrh0BVOBuuT8LxZtOeZnlf5Tu/l7UlpMRFaBitdDFcUbfWNt
M2RQFK4zXIs3qb2+gs2p4WccAFA4TYYnjkOhsIrJxcI0cBHJuLlWzkJZZ080p4U4
QpNrohd2vpdFLsPeuE4guWMa5xobTsjRM5kP7puxmyPJEk0xJUwMrow+rQYVPZRL
T/MqIxFxLszriTbf2gqMVUsc86kwGDndrupmEQebglkvqIiSraIkh+Ngi38wk+jQ
rt9N4xbFy/3sBwgxdhBVFD2Vi/jaET/E4tAC/mSuC48atqe0vONPP/IbVkKf6oTe
`protect END_PROTECTED
