`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1fiNBBk1GspiY6roMKTP69H1rBsRA/7eSx6pkjO37kelQQ2KnFNPSjf6xJzk3LkT
wPWIvOG6zHNLp7TkO2Sb/ZgvxUNLZc0KOC+2XXohBLnDltWWsEzrSQsEyHgGbYH0
f51rcUe2EPxZ/Qz9bMAhD4b1+xTTKCNRZycjgz1EaFIskwGEP+FPjPqybdn3fO+6
bfltolzUkmq8IVjiS6hMKjzDomyQ3ifpiNhZi+BTnxbzn6ZvurJdpc2KNsSnI9YB
ez+swmm9ilgqZk/eKXd1xjloPUm0x0V/2etP1ivFFedaYkNPR2OAx01yN13Ba8Ea
EfGvd0GPDVn3jhtj+47vD4HCFhnz5gQB0ebHN3bAcktQ4VP7UYdGswUWdn0ogH4f
zR38it91+L257GDglCg79/ok9adSEuThPK0knxhGvqiu2QNa6/0sW3hGP5tESyq9
cXLRR8KL7dIjus93I1aFuUMPs+KCRZtj5SMLFhHvD96a+5D/91arApsGiEu743Xx
b+sTvAGGP4qwuq8cjgQbEEIh5w0Uo1iqO9FAQxjfubSprLt/nfH6aF/jHyRQJlNw
2JtPIA/3/Pakb6IY/BEOa5WP/clVFeDQsUHsSgEyXcntiOW3epDOKHqXXxqgUc3f
lM9da7MqiZRuXi3iIJgwTDpIq9fPGp5VBnxCivxeXeZuPEARk1B/ZCbbsqNpxqWJ
n+17CVx8dEQbRAvBO/NOlWgIwsZ9W/o/8ROCxMTUVDFTYdZG0AU0O2lGfzDLjpIp
ycbWHKo1Z/C5YycvkeNR7ejIztF6L7dohgEDoEXMrddw0JW/AeGVhN5b3hiYYca1
O5qMMOdzIkfh9YEowRC60O/YYXcAWSKuptky5o6LLaNdG6F3fELWp+aCEH3EEiLL
VynW2RtxqvHtjAOziBWq8AaH+F5kuJZtpDmvg3QRFEQc+MW64z3NNZGPhFT7pzOu
wDpGrW+E/kQIvO4X72XNPK1LvNUO84H5YnflVZNnhs/8gl8vUpd74bZUzMdE+tYd
mvMRgbW4SgY26N0/Sd0V/CZ5HpOHbcsEoQxtguQsNccmaAa7+oRvyOep0OWoVzKS
51BO1kp366MhROuJrTckpl62V9kqLpKCJhs6OrywPPaRC7bEDgtz/rL/v9X9QYf+
mIAmEjybDMeHfik2qVAtahi3pOWmgf8WnpqTf9mU17WymMdtD7C8voWyDAc2qBQB
LskY5BMUvSNb4XQAy8vPnTtqytOV08MhMFUZu5yfDWQrVAvhReRgUDMSb11Vpn5p
bX3NnlL+s+PiKCvQY5kQ5AGbAk59hsB9/CUUhcPXVsSKmnwVL74IEwgwp/FJvWhO
WiFWhPPAqpJiCTfhPTB5HYl4OZvxEzUezMPd2HODOWSprUqoTMkR1bEfBv646jXG
aoGF111nADAfd0di2/bJ9AcCrBYRLMqrbyrJBX8ksdrJpK3HKh7RyWqMq3mUOi4w
W5Te1uJwMGQM60GRentmVehMzYFBAEDJe1lm602DA0oDWcLxPtVTHs2Id/ypAud3
PlPmElnfQMvKJVlqpvARE/1xtKjDdK4byK3OUUGS08hktVimZOOgfEw5A6z8VQpD
9saJVd0EYhpnbmiDusNkmb5QJLNIEx5xRon4fUCfB1fXEhLCPBqUyMWxlazXclqb
womxXXWanp23NDKvJnX+AXdHbqNB7FqM8ASLB5U0FCLT23/1x0ShyoVRnaeZa0ph
82xYQxWJFGjWclKMy3NVSYGliK59yltEQBb1R7E3XKyKSurK5gxFJx2T8/Ys58un
lGkjilqjnAYfoHytHDyRsEOC7e2kRJmWQ/xEWwkA9Q86KuGG/zDgtrfd1cQYSe6n
Ui20Jb9ZIDyLbr5aLkGTFp+Nvc3rjz1ckS7pYpB9m2lzKo2NQ+BMUDp583czCFyq
ZbjOhHTC+705FvFO+kfc/TWYvtp9YWTFfcA83J9IMQ2/ihauYi0BoIZvv6s55sGs
mpOu8U6wFYwxILsHypw7t0VY6tiMyboXhgE2PwYmuEz25EqG2524F8zG9oYpjPXb
Jfja5dihZ4JpHFHf54VaV0rhfc2ZkXmJiDdu8W8+CW4SWobEvYVP229ap5CF1pH5
j3kvAnE6yeYhHDKcP2mNpZ9L2X0ukdtM/v5d7Si6Arf6tuWZExSnU3qWpQd46J9w
qOydnMQAqu1gvrImIiZsBaDmukASaEx+GtfnojjvsgNU/gM0UcpRgR19duEe2rLD
x7ABxm5Up8xabvRdoncLwUNXlzn68ItPqh4IMSKhJ3WksZ/VUW76KN6WttpL1jZ8
uaTrCmnXPZsiUka9cLf7rQ4nkt3PrjL0S4qXYBJB4pHlnrKgkSdkH5939PeS54yc
vmuckwQew5QoXA1pVd6gZElP8f/yKk6E0TPeKj5Foqx18hmnpiGGVyICyPRv/uHL
odkmUr+T1Pb0LT7VVGXfbF9hskunQXDbpmdgeTm5y6MtgbV+hkaIkEUx1s1WXsPS
CtjzwHm/VDOyEe/eMzfxMcOIBViUzGIDLs3pDkf8AwCoUkuVywxm9/fPnJ8cnezG
fPGQzeQcvM281K0HPwXb8WByKciBvTqU1S9DnGUc1cnzUZ0v0AN/rfrlHP8aBKdr
ZEOA7SxzovvJD0dZEmATCm8+efpo3dwAYoYx6GeRz9l0UacRq1XmWyrsIUU52orE
dRv98tgTLfMaFaTwg11518xVsxRpnPqIiUxZRHm5+6fFMvYW80Zo3o/jGe034Mvo
K90KqzoipZJBRbo2nsc3XXot7RFKglBYsQnSc83XotTTHxZRzbzEizM59FWNZtTO
9x3amFOKiczh4dsuYjLVS1xJ/6ka1LwANlvMAkaN2N0i0HwWUJvi58rBhs541OYd
ewOZtlVG17009kEHLO3xmBS6XBtXAzWZZozb8BK1oPy4nsh3YDHBoPxfh1zMdFVC
VNlzzIS2WYW6xlIPxUkDprt75fNb2ZLcjuK35FBNIqPPT8F/QYqydZZIQTFkKmec
36yH62xCdXGWK7+G22EvmkmRVn2i9AQIAWDPizYYSnQxOm5zc5YePITHu5AUAzTE
6H5lRkzmWJ22/bwPTeCkl1SVUUibsbKYLcQ5eGrLn931vFqYjSG8s5DXsFEpBoB4
q9/Xe9JHWKj93NOedNvgeQ==
`protect END_PROTECTED
