`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LR5SBFqwUyoPLGS0CwjjSNXb5kiWxNoRzS1DrlXKC6fv8G2juC17W080XMOEJifT
CYxInPI2XzJbu0C9CXn6sJ4tCZy2hCfu0f59jApA8Lm4soswRRLmDkS7mSAChlhr
vUXX5Uk6I+sb4NicqXLolXWxGsSJiN+UtWAvQFFEUBJPgOgkd4hAVfoBQHnDjiCj
GKDqOF7c+P6OF6/NZbK0BBWVaoPncu8emCst9NVHBclE4g51wfu+8yNcyJjiXqUg
vRh3o6d4Bq4YdjIt6oPStasgHK23FY9BJ2B/YqtcvpgK5xR6SPwhbPRD2OnBC2sy
fsxQ/QoHFYTTCo/BsW0uWAg03alIqcVXPnfruqXIHpi+gYhfU6kJVBZFhsubBIAn
ZEkL8CX6B3IhCaARbLIGSnPIxlutLtfhQ6AByLgRVq0j7bm7uk+IgSF2Uwj46pJr
`protect END_PROTECTED
