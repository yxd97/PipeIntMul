`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5K4zwO89Hqqu78hSG+iHk8KSlRQ7DMyhSN9VGl3W2KHfZeDCa9GLFeQggzW0e7n
8eV80Zb5hxF3LAFHPJdYgCJfFeRNePM+xGHOeFnz/QUSqnARKaFI9MRGyuou9hQN
kULi59dRvcxvoq15RPHofztyA64CmFhDmBNQFdsbNpiBNLXv8gbowyOOw7X7mxVs
FjJWsDv6dkIr9+JDbEtRyPH0yJFHkJ4QeBJTMkqhov3YQdn8fQsUFMYcrJaMGL7Y
rx/b5mYMt5W08/yqdrkm4yHkuJkjG7/1WDLSAK5UI6mvHByclow4iubG/7l+k/wE
2499hA8bDxPsJlV2Ee8vmwlN4gS+tsBf1r8eBB/yLvUcnjUehCs7PEVqB1BLMyRz
jb5ebTX7UdxAN1Da1elLv5pLmrracwxUfZ8j3MN88+q9pVZkN03VXZloQ2x0RFUN
C+lJ4nVJ0sGHHHb648fWfDY3+DTj4g9HiE1hud704jxT/DhTcUJcWZs/gtdMbyJL
bLUEY4vfZQaVEtLNkDeL+YQ6/iv6YNNEv3cFrZx0bm+RtIT3Crl0ssoP2gMxeAXR
6LGrQVVs7dUW6V5zwJ79GZJHWn07A6Hi/5I57GvvrCY=
`protect END_PROTECTED
