`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c3reQqO+yLAO9xhBUhueu3jG+yiHXREAWB2Qy8AUlLZLGrR0qCIMe0176X0kb4y8
WuB6jAOcDUviFt0eneooZ/UkNjd3Lgs64Wjj8pX9uFZJs+GSP6T9iacG+jVjeoF2
iEZ8tWi1fFqe8wkNGw7jpqUPuZms2sGSfkIeKe9zg7wyZXkU92C/ZXegum22m9pV
ryP30+ctdkP6y0mR1u7F4XcS2pOxCnyigbI1CiHZJxGn8ziF14+yhUpR835yX1Rr
CxbpTYMAtjyXxKXCLyPbbK6Jpwh/VAx0E8MRaGL3E4NDhs/YvdNfjTFYxMWv5lfl
OdtuEHSzcwODOS2JUeifZ8PzBD1pLyI9IcB69h7alVIbl4Ly92w4zbxfr7lyd4yc
r9pQKC62YKuM7u5/UlRD5JNAQPAFKdn/ng6I6AArVwyRczUnBhpNzAlvxhF9NQyT
GD4uXCnaXgk7MSprNYN73yj0Z8OVpa3uzxNKCpMaUZy3EtFc1re/aKoNQERDWV24
GkYyS2O7klqSrl4pvDAwZ3rihT6EXi5ZRKtMc3KdbSnA1eDTRUNOjbWO2ot/DsW9
YT78QMiuh8hScUor0yeM6DTSLIY0PqtEsy4RRpOUxqogyb2Z0k71sb5ZRV3ZHqrV
acy1MRJntEDtXGngEPbJps0wjd6oiT/ZzU+UefxCkPwrfvfip7QPChvcumBSCW85
sQYdfEmAsFfbNDjwTrNLFreIURKqFY0FWQa8tRyg1ycsMuA1oVOzhaSMB4zsVWm+
XBEXBWdUe9mjq8LlZ668TIUs9rehQcbETzaUwv8+POJ8/YGpXzYYX11UF2um5+i+
gtOtMjSFVZ2udH7WMDZdWw==
`protect END_PROTECTED
