`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XW5ibIoV8xuNxi3XSbbO2j0j6LLuGvYAvvO3DZvZkh8han6gL/Q5ci5+cdlk8pkk
4850ljdpRqyscrBkYD5IyIpwrSMrY0O5vUhBXs2KJqCwYPTtEMMoT5XQhpv3hPa8
o55XljDB5CAVihyLkFaUu3Fzu0Nwr4dG65tlucL7RaeefN/P8w7mWMGGVx4Ati27
deTka529doehaeLj67DJcxpU1tC+Yf8fOH9Q252Wm+8dmyEaoqbtrG2Pmm0RywnB
f5ENgr9eSHFhm15+xA47h7p3BUeUieBAnXeeDhjT/Z9+4IGTw8FYet2Lk+87XSSu
rrLSobHD9QQ7Js5lzSBo+hoB3Ik4kaM2TlODfGTE5A10sThNleNILb9xfVxuyLuj
7vQ6s+F7BM5e8MvJVXIDxuPKfQqMUkw/ZHtkIpRcyr/S+Vt8eIV+a219XZvNIV5U
Tmi/oXSIWx7VgIev0/M3I1aT6F7cWG4xa5AuRdwZrvfGBKEiS6VRAtN3jnpztnRL
W/nNa3Fb82OPrZPQhA5ENVIQ57OAXH4aftK7zHOoK/dltKDedh6EEV42LUrwHqvM
ZUxlVQ6O3lZUPETXRK6gSYfOMkLg5iq0gk06PadjuepdjlZmnLOCWveElJSPIOIh
vFdKGvgzXd1UoZ98u/J0UWc0tI8GunMxgqJKIavPa2EbPk0TgWCJzUBHBpYUzO+/
ZyoU5ryw+WqKJ/OUAMvg7qnQqWEQVd6sR3dSJgvN9YO9I1M8ijh2UCIALUuauiG6
`protect END_PROTECTED
