`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cvMphVtfMTnbGnNVQZrK9mMOokTRRi4ASdhAXqodWOvzItje9F74DZfxhKTHjbQe
LMI2Q/RxnrrRHOrEOxhA2CWe3xv1z4ompIoXpg2GNnzfhDMbJIAoPuuzvIYQFP72
UxVsIottmJtNSEvM0XI/icBE9wjKRYq311Dx90y/lMqJ3jmqwIA9RngkZHq5zHr+
p1M63usLntSRCDe58feFdqb6deU5iGHLTHPCTX/+HzHwJzE43k7EIguQoP3Q6tzH
t4VAgdFyD5hfHVnQUAEZGfmgUu3odnkAqFvzUpFDqpcjr8a5Sec1R/tx/lGO64wz
OS2JOYA94X61zGwpC5FcP/TmHLBiIUahNM6NmzGgWws0+A+sQyFLl3J/Fw+kzMe7
pO/nqEFbhRL5kVg6wJlXFatE5SkqYQ03jKrTHBdoBWrm18UvLJ/tpNFkIwnQDpNJ
8Cr3+GaEHP/DorqNM37rF6RCKArjUJCA1wvr02nHHzNcdWlgt+fzMyjBS2HUIUG+
`protect END_PROTECTED
