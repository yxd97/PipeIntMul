`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVpoQ2Q5Vvo+6qVMWdjrTpi7bAnEdnjbOTpV6TVCfncSvZGwrzkixP350VjBpdnQ
RHGXLrUV+Azq/VxxUUMEJZLrU9+l4/y6LLZ7YG7DxwVf1l9AI9Xtnah7C/kAJ1KJ
Xia2p2UTztr98IdEh68JNyjHYjmouHBOxMu3MycW8GnwLdG7c6NwH9tPxPzpTLFa
lfaYmGVetIIpkwQB7RplftruT8DJuKVnGwZMJmMT4l6b6qb9NJJ2Y7l10lFGhmUp
jEw5dzSO3hfEFq4TIVPS7g==
`protect END_PROTECTED
