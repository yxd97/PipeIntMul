`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s83ZoReEs6RCVe+/5Px341nI67yYSqOmkc99qolto/uQxLadD2zzSkr0zyDRvIaK
R+uryv3wVDkwnVx58U04sYrd+symdTuiDHYyvLoUbXouRyl6BnAuIYhJWzbj5Lhq
dbvGL/XTEXMpJHDrClHHX2a26UJGzOlCI8CLHdJ7Wro0lc2Dio80kp8pgHzVu9LS
mRAHPkSyEe8ZmagOlepbw/I+ExFN4ZyjV5jJ/xzBIjYCzwkwQoO4y5UcBIscUs6v
F4uiSu9ygBmNCUdhSjSGVW5V1/x0EbSOVGqsCrdsc0qaoWNowNb6ukAzl3EnfD3X
b2SEVJkbCy1SRWKk4hJe0XVJoknZwtUG9y8t4Sd+0bM0LSgq8Kj14khG7P8RPKbT
PXCs/3ArxFcOASFgK00oXUrlcu7+nsWt2iB8Brzv1dA=
`protect END_PROTECTED
