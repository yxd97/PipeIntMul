`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tEUaMmdXf3mwg3PaL0S/MC22fmHJ+i9G+Tp7YEiCi45VCH9CIUUTOlu5o9reu9b2
BMTt6R3ZC8tRYXXE8UNo05uOMaqIcWA4htxTGfVxakdVJgossu0bzLT4gkt7zB/P
ZoSpcc/8NsRBI7l8EWDK9BHzBBFuqoWYDjnIaHzZ6iCC1We9dUfsygJKFmbRJyB/
NzEFGBpeYSvQ6NGQ7CQ3GS0qgOxBbRHguMW6CvRHu7H4PoctMRt0yMrF3wU7jlR8
SZC1cTCFVXJfBUlQEpm7VA==
`protect END_PROTECTED
