`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j2ooWVeka1VNHvvJkq0lBKDioIUFDzue5SzaGjZhwNTL00h2m1iOKicqTDD3J5sS
J7gKlyRCYpwhfcIhfxHnR06XoRoIgTxIq8fCboCGe3ANAMaNtWIMfpT3coF4Wqk6
nYyCaMf6MCH3oWcz53RgBTfJ587sKMgFtZ4DHCHllKpfsERPlKLzfXgMfTc6wMbw
gR5ksFMsvoOBm+QgYos/H6GxaDQKqOCaYvAe3FkGrtlvn+nPP8ctMrq8Y8EVv7jy
BeL2g2NDHx9KcMtk9l2LORbSnwXHrUoKqFYpiU9ltrep+oNttWpHUbVMq3Wv5oMB
wR83FzLtv+Pm5jnhezIZFwK8kCJbYQ2eQDzUCMsdQHTmbFwAXvuHD5KsegqGUpfG
g0reAxdpAjMYWVKBJs7rj4VCgMJ4nEfzTpreCTOm7s+7aJKhG8sL/oQ6LFOfDRxZ
FYBgz7onewffezXiRq8c69cmrWA+2f0RTMFJiBxxdWCdsGE0UlGXUf5iOufaRS7d
+BOIM2+darOul/aQbgIE3F7AdrIPlPX2MCmxBQgvMM3KYghahUZlu96QwcHFkXGI
VkUrif7en7UTBkzSmnZs/NI+NjtdhedHNTZRaI/QUbNmZcJUInqDCiuXrG8wcXu0
24W2B8JSJIp1CCVMnv0G450WPbD/WeIwWalydgOcB7bn+bsdmxzysngSJgsys9SV
3tviz0b14wnPm3J3xFi/FbpIqK8pX17yY67N2Yy9nhyAbOEBmt3lO9DoRbxVHyG8
PUFcP28cfjoaWcUgAz3WtAnueaJDzKSgi3JbTEmsc+ZQxXj8wRoHz8pGqPiBJ7Id
exbpxXEEQew4E9qrf5o+4m5Ni+b/PJ2v5MJtXuMa81vEuBsgFBlHh6JK7DVdcp4M
gCZhXOBqsXRK0OrSRTFV/6Y7TfLH1ATuiTN1DlGXR9sJSlLyQiPdPeeAHD5Vd79X
D0qI7FaQTZQAduH7FAa/6mGBBpsZemZwMscSmPOon7vuUKJuEFldzEgPeshq3BmA
/XG1AphTLl38yYSEOEX6uk3FvBiTkYcEGvP1wmedW6iwOycQrs7ZCnOnw1moEs6w
`protect END_PROTECTED
