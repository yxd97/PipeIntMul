`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lLGjjqh90+JPaJnUupbYIq1uhgvWjHF0cy4KA5e9ATtlEuXEeO43tcxeledxkHWL
wUpVAB7xds/T/QaLXUe7cSDbQP3ADQBJPGPXb54my0syAyYSVS3xGCUkqqBFAGkP
nI7f/l/rTJLJrlapXDIld9B8D8v5MZFYBFESyPXQzmiGMziqjnJoOk5HlTWzf3wx
m8sXqK1SRpPDqdzoEVHPTodmo4okVElXq8COYthUk0+ShzL0zWPyzN8b2UjRTAoA
+fRg5Qixl+5OlUOdE6J/eKDUYTuwE+2HJfrV10IVURxMiI337QmpwVKWJTqjOLfs
9eNmvBpZnJMN+AHs+gLjkJL75/cpMG3fWBsQ6ftgwub63DO8gEwqlTzcMQcJtstm
pB5FyHafrYz+0lhw+haiyruCFyu34FjopKwtAXOkncqJZApZUrjogp9kv3jm5nNN
sPLq/v311eh7itNJsy+fuPNRorE8ByVR6OziAHmDjwI=
`protect END_PROTECTED
