`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XynSDgmTrpD1Io5TIRVkSscBK7hQ/a8W7CxmCsJ1aVXkH1KjmQo5eUlD50QQefZO
rEZhwXaODhP/HoN5gr1T+xj0kp2CqQvxlSCTyuQMTXGyd+YX6pD1eMmKbbWrMxcO
DlkLhMv2Yts9Q+bVSKtaBsjYzcYXgla3XA0+37Z1rq3n5AIyJ8HaQ0wdO1lZGkgh
hrZ9OwQwEdzNRnX4mSxWH/BKC59Bo8Yf4SJdvDs7GHyHgk3A1e6S85PRROdnHrIw
FKfPfRdc51p/f9egm76Pjvy/G4OywQean9MZQZ8qdtJhilfWQlGM7XjVGq5cv+rT
33Vxbv069/wEAjdz9Y1zRY6jozblZxc2ofsFZrZ3xIJMbT7nv8/how1ItLKxgjnV
y+tnVAWRlfdgpWJFMO95cJdHHMWUWeYTq8WG2nG9Y7s=
`protect END_PROTECTED
