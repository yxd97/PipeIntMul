`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gdFwS7V/nqRPhmuhPKL1TeqgSu88eZfnB2x/wLg+QCpjAv2HL0HIr28Uu+aFhEv
oXpWWSVUFQ2e9f3SsvTeUVtiAZF4118GovI+mqJZGsMrHfTULhvboVQaYrD0C0YZ
WGUXLgVuRoLxwg4KriERitxvMPOcZaSWWegEB+ytPCrM6EaafbNza2on6cjNSl+b
McAsfLjMFx+HQvx6LEvIgs2kmA7Fxai01xVgqzY5e48H3vFq/bSNNkvxvA8hCGHQ
`protect END_PROTECTED
