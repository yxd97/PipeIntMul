`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Joa8WbDzA49JrOBJNmZAhZb7XmLmCNbDH8b5ekU73XfglpNEI9nNzLyCVZ00vvp
3kxJNBY8JqLUbxKDun9YF/VYZQ+osN5xMW8lEj9OxK+NlXi3+eiDqwkLyl79D0UM
lG6ZtR0UGxRRp5+1jtx86y9XDJO1gUedRrvjlNgjg5k0yNTQYxg2I9uRNf/cUngw
weKmUUEBrc9jjt2PxHC2jtDFZwVj3BjbmWSlEADluFPojjn1v8siPuQOfIRk8Ut8
KHs3xgweCHDM/FfnLKVRCjM4qNBW7aTWFGWIpCk4SslbLb/AQPlmgendE/8LKFB2
U2roZ0YmNLCFmc8GxhJgvploiMyq6jG7V46ziE6gHnLZojFDOfg6wMrPylsMmeDM
FCsFSQNam2yYg/bGM6hAY5NMll7SrMEC37Q+FpRHgyVoxkBGgxD88OXIpnVFfSyw
3YP4Z8HnbODkMJk0uIuBMgjzRdEKNMXWMTY8nyb+tKf4mA2efH7K4nVVm6dJt+Us
v/2ZChsxH52A+n6kKnxTKvD5n5xoTO4gDgHBfFZ57O7Ih9InGXU1s8Gm2NuS36T/
5goj10H49XIQyx5XNlkw1ht0+51QnqTRXS/YHG0Ceh7LqkXbO0dsKeAAQ19wSXkK
fa/V8wTFzxMHGR128wGWLlIUXPLXGu4GRBjn5LWMwMdzlDdZ6XZIRO/DtWcraKA/
Akr1SXwk0OMU+FnQVzok4bAcTXkIvbCFybzZhP6ynHWjNhxCsZXARznmkhfeH0Sn
py+vKkRenFsQCSMaKOXZfA==
`protect END_PROTECTED
