`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sN4t/yhE3ySXvXV4YVKEzEbgthaI8AbluFZkd8q7zcvYFw5EwQGFJLL8AuibS+Tf
66WEoKuzitZlHtThZvGSM1D0dk/iwGAnWvGH9X2CmVYWlSZV1gaAGsVC5O4rD21N
YrdI53aclg1F11gS3U+RxQqr71vVR0aVPM0NKNfm+ulSWrsOKzj7vJZtiPWgPaka
MpL7Qg31NcOM6K0knUDtPAnTTbAsvRxkyB/REBShQKtydrP1Al9fdZVH9DfMqP1w
TMRoBGbubsnuHJF+pwk9gE2f9smwSMHekSSwE5ZfT1jP1rMi9Qg8UNPDoJTKGqeb
TKWNTy4YIXyTCcKsq0GeqVRiSNuvelColjkBE7yIi5+P8aPGATBqC+/dD5uSpTNr
rAMrsOaa9DsoIoakvvWyrtOk+Q/nsp5nwwJWnIKpAn5lo41Vj7ouryFj9rV0D86H
Nk7uEM2rR8nK1T9EJSs+hv48FbZhWQE+52d6DoWa/gqgSj31To/6cuD6/6bsV9Kw
M1GX5T5Y2gb0xfv6L8tsqU4eRG6aO3LFciY9Txlx32Yy+HpzJi94QNuhfHZJVTIT
fqIud02fbuhIsHIOBZ9zb7b2MqBvkSsYtv1igZ1IKqTAiIsQwmz0EIsKgX8NjP5H
PZGi5D3Yuk8009XNqoHPoQ==
`protect END_PROTECTED
