`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XwH6o1irJ4JgjnITWTmwbfxtXH4BGxCtWU8fSVJAOs3McBLHpWlfkhguSoThkx2b
/Nbs9JVGmYxKXVE2v79fPd16EAsu+oLWsy7Q+SUplefcC+DRLSAN93iB5HsTiiM4
rO2Qg6kj4WswyC7okwNpAR+eBlY01uFB8wqxkr9eLNU5WF66dhd1fbHTcOEEsGmh
ykNSZ9tsTfFuvSaAkLjHPjdJuH8UV89dE6IHBLMFvH9HsO7bSsahoymfDEoFmZGy
TFkuPkPckAZCpC/bH3kmCUFHpzqZK4o2Vf2oEp7T3CCXsLhMDSCxchuyOSXLyMZD
M73MIF+cejZQgQqql+efx9hYHflTK7uLfSY2Cja7/OC6v2W9U68X+1GWvIpwfsbD
hqfqVhkJiKkl2SeGrwZlbaBtNV6LEMHSfoUjk6tgwVO7RCUbPLHsH46t4G93vx7b
SPiU8gRKl9xIC0QwC4G/fuD76vaJGNkMGm+mZM83fqQ5OLBuehV+PfM2Ea57ds44
rARt/7RRBYnxZJF6eMJpX8X7B6YFrWAOd3p93oGWvRDz033lgt2q1lWtLzNDlcY/
OUmCesID0/V41aQyoZI3dhSeHRgrkhOkoIr+Ml3xyHdQLqRMUJnSLDxsoE6Y8a+y
xAT5MucPNPR3OSZW+aXzW2hDNVogApguNXY3rkaxtbOewNBu6UrUTjGwaFZXaZ6c
ASZCuIwG8oVwJUPc6c+ye7iUj8WKhPvAx/h9caldKmN+O1J40m4brEuR0c/uI+GH
VgJWyD9ooYqnHPxDNEpeu8IkQHFa9CWtl4e/65LOUZv2sn6j9tltcbAJUmzHauJc
cFh77ksI1i7/fqrxFpKJFiFuoYRGkdxcW2otJircnJhnDqjvbtpBRpVIODOOLUnv
jDmu+MQVc8gKzEgh7bi/WEWidrNjbnP+A7zZDUXl+50Koe84WlLDSl7kkm6WFpxR
xbGHD4oblcrdzJJE7TGL5zdbszik9/vhs60Nml7SXSOuGN8w7Kq+WFHsuQT/G+a4
0yGkHD/I61V408mZCXRuOLEr9UTfIFXTreuVYcx6bG7xb9+1HQS4upg4tn6f86qi
HwtVW8ChZR6iVJnxbJXAGPjc+PURuuLOpx2YwhmCu7dJu4WppM9icyUUGEpuksz6
4ceLtwK88KD7ju4wlMkSIksm/EDLwx40qC8UimHGDOqGrU3DYPyZ12QlhHwiVTU7
CVmFeKXuqEb1WPVv1IArynZbxUrkmYNnGS/08Y76Zl1q30fVsVP9aL/d0ayFOaKJ
OZ5rrhkhXnNy92IJ3rUDccCJR/h5O5ZrTpQzag1QzeeMTc/BRHHzwhZWLSMUAwP1
uWpvRFWvJtMS1orv1/kINixbUQV44G8gMeTiZCO3SFMiEGAfiNU4g0BshRztjRJi
ihO+4vNdPk/NWbemqsCUjeEFJZC5/Au5Jy80QItGSmvmoiF61cxGdXXsXSojY/04
paWFm68EV911oyX+zPWqMI3IKeAh+mBBEREsvYWO1GOBhkd2mrygJpHtOLsK7U1j
kI6GvpUenulMMG3X7dXOK+wMYpo8NiRuXly3nYXgL6DRFwKfX/6tMWIjihhqSjQA
9rGIl5u32uQ7LAbswA3N3TtuvWtXAThkfYOZ0vRKuh9RBevc9yJBUjOV3gnkWEE+
fbHYdqpqaJtOvrPqzA4tFze4Tbwb1GTWjQxHSo86z38bvQEbcPDQzLb4pF67yxAV
fUhXR4PeokHYOgz0k0d7ChPAF6I0HyJVaClZIFYh1L72QY5JHUsWqqZNxIRbqnUr
PawldaNiUrIyIPZ2hcYUuDHpvIcHycUc85JbfRmwFnh9NtdecV7EHsD6icDRmU1I
sI2S52QJUq+S2hVcIUaB7VbDm5EGN8NzyjH7QdwS3KQxkbfUUIJOPLo/dLOI+9/R
jQWbS/BXw697onuZ0E8elVCriT6F5AXHxTcMMe9aUQSqkC/utvmdJvKwq5hWDdoj
unHiDdDx99sx1sUpx7KYlOf7Op7mzDGWOjdDOlDLVGEpdZFYbKOulxDBc0mViqjS
dBNS6oVRB6mF1cOEFuduNNQpFawwk709/fYMcWhjS7zRqXvdk7twRu9u7HWqUvfC
NW3mrZHu9FbpuNuiGg/3SVbeuRjSIiY2Sy4htB+KCg89M20N5khbdjQidDPsSGHg
xDbzlflS/F0jtam1/wDkqzFOGv/W9F6/UuKaL1wtFRrm75aJlQMnrNjg3x7BN0G1
yFWJGKuxNnOSYa38O6jAALc8HE6836SmGIY29oy0Mb9ZJQREtebQJn/xqnJYVe87
xDWCIeb5WZmgkqhDewmAdERG6eiiG/OW/cg3VcnOjdCVa71QwMXvIuk6ToDOq6ut
G42Xe4vap28S4Rng/UMyj3+wYgotpuR86utZMrT3BGDkWtEZ261mgRCm2FNGz8Ww
zWGrjHylaqlAlf2JUabpThK+dZvkl5jG3jLWSUN3detlMQ/U4bjDGHPbJweU3ZLM
bdKn0wLlfQNs48+qtXvqi/2Lf+YrGZmPaRPjHAtpT6YS/rMBJDNbZThQB9/w3BDh
uw4s23j2ivM1cLpaw/o5wIik9V6dJc7vnj3t25jV1SKVccgqbhsz7U9JrZRKEMJ8
NL86SO32LS3/Lq5pIMK9ggvd2jB/zOBh29Xur52HO5B9M4EBhH4SSwyag/nYPM7M
GrHjU2LuTuVcq8nxFXBIzoaLc0cL0P+2e4AL1/ch0HyeDkdOOL9SR5ez2md3fjh6
u183u/Ch48OI4mkaQPbEWFo9mGH2l2e3Vvz/RJC5Tcv80mKvtuBdRXpoA8pMCgeX
fzkkzb+qb7ZhzXkNVg0UcPfETsURtFvOoTa3KmzMSZ97UucciwHkH4rBLe2P8N0I
wFXECuaNDq/NH2JgTiEbDaLPZtqfKys1QbxDUZ04u4Px337dL6dqrpZBl2zJcdF2
mk2S4il3KIDrZx3x3VKboyL+27rPIGOhQh6SB4NHsbJsRBf2dTQ0vLdpYtLVHOfW
SD83KVrKuTxfVSHrzZ+Bb6G3124b50m1i/yyBMrkEO2Wv6QLS8w1YEPzuVbRvYvG
LuQqK4gEGxxEFrvMK3O7pbBVFUrQfNMi655hVYqEh3Py+HkhXYDkVGSKzLvhQ2PL
X1pIresQBtwyQImk7s9I3mr0cKx7c0rj9m26pmBWROOY6cOQ8AtVXXNWodwruRPH
DgP8lJX6K4xFYT35BW6JzJL8mBNjUzntBlTXjE8lvUr02oOkCWz0jNw0b52DhLLG
iR6qXxlX0xEyk9RCb2YqJ9R1lY1tL6ziWFsppuD2Bqv8mfbKYjoQ8b3+MDmTXLXI
zNJmWwcjTPas5jm/Y0gg4kLQkMEjrbrloMj+KPld268YumH+RSoHZX1rKhFmjrQI
NPjDq1LvPya7ui37IRGfygQDFU0bGJ+cpIcUor/Bc8kH7gb+n8/GoPKx1HTz51Bk
KHhlFvaEI6j/c80JiuPee26p4idMVEXlrD3LDP3QrtWdJ1+a1k9BK+a7xZsF4Otb
jeHUjG/hkKz2Jv/g/8I4cbdasBv3OHGhHFcRfRjcuTgSdCdNjIc9CnBehE+bx8UK
6ngYG7igoctiyI8/EbNrZVKdpg+VXPWm4LjZ/3w+VT5VCvXz4C1d9dabfnbO8Cao
yZpbUXoV/iXjaOAWVIGhJTHZlTzc8hcQS1rKeYU60NQRjgJa8CjBdJ58ipt1JC0a
Z02PLEpt4z/fUA+kxMytL66eovJVEF1jOZhfG8yrXK06TK0wT4lwBozlJewteFpd
5PHh3vebcglfhysWPZdRuvzjDyXJdaaIvI28w3vksD4Fski8FNV00Lh71Y0v8L/4
1+c7Q1tXK4DLwnrkNsbHdPAAdoRksDCLmI/xVg58tC5wH1ODjweciukyxVBZAZsZ
n8IY9wMQm9ACU9IeaflNPd0/Sx+mpM27ezySYmZOsmvonLgGwBNiZX42Aillkg+K
JhYYbOjpKUttrqn01pYBrj3hh+JzJ+Nuy64mjkHoYIGdwHV6lbN9xoCVXLqlNSUc
Gtk+zSf9I5WdMmBhPXC5FrnBqK/osqogd/KXQf/1Ulwo8cSNxCY+eUYJCJ5eAbky
CRCPraVUjdhBt3YBVkICl+zb36ERt4upDrvExmnHXgoJ9j2b/RhNekNL9FwktU6w
IdsuuGbVEMUreoS8UnygMAEgFluybf+TymK0uDGjT/kpNrzFezh8ZDZFrCjrZ1r9
nSb/OG3a6JmS8K0HUV2s8eK0tJW/AUJ6CUppaQ4x5HMKWwWVSt1CgkkeftLPKTr4
Fszfp2g+YNUAtZf6Zhoxh1/oOpDJVki7pXVxZT6/ENCoy/8D1lvLfi4pGqUDSe8I
CjDme+24YebD2ECGu5l1rQYTaIsDYq0QB6Xz4pO9Z/4RiMC1w0r9FanxIkdS/jxA
mGSG5+0Taf3+bU0k7vgzbpzIxtfdBJslMNVe2L/CAlCMLnyKp2usvmfUzuvQiC4q
M4fhsEx689lcpAwJh3dcsQnnhOogyPFfjj4mjJbgdBTUHgzfv1Zq4eno9Aa6VvXC
26P4btDs5Y8j+WAHP05pwM1NOrmpnk0e33XBHhoFkdTNJNBcduF6TTFOr3mRkzJl
x03UTdhSwsgL3dBR/rFMZGM+ioE2jcTHIgbYU6bWo76XrzkTG24NzBuha4+AQ/2v
S/FeJWi9bwQIF7y/gizVMunJgC5WeY1VDmJteNPUp2UkXHv+IK7zNnKbI1sw/Cpg
G7jcbIFVrGGGV16qyCpZPeaQyWJjsnMT7kHU/C8aR+N2pdsMHZQoGtOUU/mefnsi
rwgMp+5hdhASY0Qgg1jPMcsU1aypPpnHXzDgtmyGpuZ/dfERqBhReaaUAk7aF1kt
8h8t1nMTsRvQHx7ZQcEDFyN9AuJWjwuph0wdlYnxHZm0XsMX0gxZQz6AGytKx31y
zwtuyg8sZc8qcRXtbXuzPsW/kElDZRpejFyOxfKWLptibNvRJoL0P73s5/uzKi7G
baJwkQVDeICranJqB+8B4Zq+/FoT0MlxkmBIt342qstWIyyhH+B+JYe+DOHRhlpl
rOAVjA5Wm87l9N5u4Z+0hf1tru4UMGZwtjypbthCW3sWquQ+BsKq0jDu8jwOHSlf
XtpFcApfZzm71zYHP3p3Dw==
`protect END_PROTECTED
