`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDeQfY0tjQk8gZ9aKdifa3SLX02icjCHxAG1EKnKxdZALwb2MMrnUaZ8tpW8qKvW
zo9geNSgMWjLO0Qzzk4PZE+TujJbFtqlw1KDSI47ls47B8PmBDeXaRkjpu1AR0MY
kSGnXFlT/UofVbDO43ghLXQ96HF0AV/TxOUVn3+AnodYPJ3Y4Ve9MwjFnXE6oonv
fsDsAS5ujn3Ghkkr9ZU4GTJwJc3/Mljo2ri5zIcvGyxT1Y5mMJzZeKJtW1rpaBIC
CoDC1ly8trrrbwTuNXUXxAPZGvC0pEL4VlhApuz4ips=
`protect END_PROTECTED
