`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmjLoWXT+3Z5Q5LEaL91YVHgkqUQdxdsP8E0iZ2kMcSUYKeuv4s2tgjH3eqHAL/e
HW8g8e7O4qF9syKtqDBYu2P8bk8eB7efRmu2bwjqcPbVhzR+FJ+TQiAkkxamdbmU
+TYG7lkaRQMikmxjly4KarPgiCBcNmAC/97dg9TRvLId8OEt9TdTkPjOMQtiwdmh
/vLq7TehtVO5KiEChOGI9CmQDaUQiI3ESnbbP78B7w3t2R6TGOv+utfIPYmrUU4+
qCc92WbSgKm7MK/8P2uKbQYhYUz23NPaHJldvijQ0QY=
`protect END_PROTECTED
