`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2UQrXyoF2f+jJbyxufPwytPcFvVjavsRBVC29A9eCXSbYCpdRhUuASnSsjMGjPuC
hhiX2fKgU6/+IRBNx17UxJn9oflNOpeOboA75z5+hbSSGQcRZB52aLmDh/hqUo3z
MzG6Wh3bL1VsYKcGRdYNaT+0XQAfXoRuM1NB59RhlAU4c8CdgXvT7XF4gKk5goRf
MKinCkNt90jl9cZ6taw0qXVkE9vHXxVuJViv/Uegfflf2YTNbErt3eOAWDImZtU5
POZ5bF2qQD6kHZIoavLVSbon1fNBWvIyl0WAKp/zA9ygCN6jO4i9tX9PWBXocxku
0K7RnN9NhfLf7/PqxIUlhGiOtLPBS5qbLR/UKjyyX0R4obNPBGkEcCPNQ3Y2RGKx
`protect END_PROTECTED
