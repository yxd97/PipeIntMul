`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ISypZrE1tr/2HvNL6T3ylyLwhJD+A51cJOpUWUZD20gaewJBQjBIMSCrdU42LsnH
2MnwR8rqPVBzeiJuTYwILHBQyCbpZJRx4XOfRc+vl7x0JZ1guw+SyBql3CDUioa7
Ma0Jkfg44kLHFecUAHs5FEWkI977vpsVT7DjgGgUfjUyT4R9JvRlX0ozOmD1qAcZ
2kJTwWOfduGMNeJshdlCeffB5ytJEIve4CyNk9H98dFBNwBijWUAbeo7Hmnx2jpH
zK9n7LhzZZZaxPVAXn4qbZLIaRw6Q8stoAj3rUPk/9CBddd9fzj4ElXFV7kQGKst
yoQkfShuJjxroOIBCCPcyUfiq7fINwqUaA8yeNYw4A5LyBojFm40xyYZAFUjN4TZ
PyYZeCQ81aP/oS/6skjK7J6cGZTNFbvb4Cnn9PawlcyXl64mZDcRinqhCnJNgOge
X0u/uo66vvS4EqeaOqSQkaGYa0ljlK0RctUuB1H30lU=
`protect END_PROTECTED
