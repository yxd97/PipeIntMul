`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RdvNhxv6q2Bto1VBo1cOR7JCdDFng+23E3Y9s1IDlVCpyBWIAnhmMxQh3nHdwZJx
HnoTC0exw5D20udTpMGXEt1uNBeAMc7E6lQD1RGdKA97SZwj9Ii1yH9QucK6sr6C
yz1AhQ7AyMrfEGegZowWGSuNRv1s1g81KievKh0Y+OlgDeMZnmMYneaKqA/7BLAG
BkntOueoRiGwH/BOGJcL9Q1Z3CFJyGL8IAQCtvY3xJnXW2zFbKn7Z0OpNWl5B7mo
/TRuA5JuHnPQVnUW+Ug8Rv74Vmfo85SZwhox5dq5YMo=
`protect END_PROTECTED
