`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyFFCNJnzobFCNKLUyQlRlTjY26TsJqL2fB3ysTKB1vE6Lp1U3tgMO8hE0s0CjBn
C+mtSHWgiNtUn1PigHzPbwkX9woXtze56QSdG1825BJ3Up/I6K93/821PlOv0ogd
kyV7Za2Fn0Jz0aLxVMTDgNduo2wKVSNHXJN4bdF13WLigI7K+ShDRBz0eEuz+dhL
1fQd8ubIpxyExqRCRxOWl0icjSeGcvle7rx+ZXKqNAsKHWLZsC29DvxF07c7O5It
JUmtR16JH2NHG118cWSZONcIsu3uRE7cnudmPJwex3fxEH3yxGSV5CGe2WpDheRf
2NGBvtTk8r3fWFqoWlEnBU97nCS6boVqOL9KdAf7xSG4PCuwIVUe4JKHBhnZb/ZO
KWGz5bIl3bo+h1oNmC2LjgWKMiaiyRA/6C8M/nkkOZMiQ2nxLhaC048r329TWRTU
vH3Eg/prwgVXR09X0tDNgC0sDlQFXEbJh5NKRc8QIgl+Gr2XNCgGjTOzKtlwP+4G
6+i7TLm7ifoce2ElhSSqy1OXpniqUZpUJLb1AxkWJd+HjU0ta8F/u3kl7GsgGyqY
qDhq5OvwbpOE+io0APktO8xBlLMG2lVwr7WepW1vpwMg+su/fw3jb37BHGENYV+y
BN3ydgvYx6Zofn/QkF23RuVPo2Ac74CdLpIHglFjjdLA4tgWQxNIrPN3XtA64cZL
1B6SrBarlDzdLhVenVCEVXMZnIPo1hVFbkKFxhQ1S9hj6XB9qalRbAGHji4CbbII
7ejzcbfasBmPR7nivAb7O7//WxfW1eQN1n9OvaRMOB59MNVE/tz+BTaPEnS/c0bR
DK7RsN3J6prubv9JBloEj65aRMYeeA/XYGGSifP3MG8=
`protect END_PROTECTED
