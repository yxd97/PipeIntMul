`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8nMg4TTDTMz1zxckpwQCKcviRJ62F55NYtIVB5Qa3d6O9GntO2IMzHwse3NFQDt
6B69spuXiq20Rd1n0CJ5Bav3XqyJges2JsF3Eko07CZ7YS6PPf4rwyCyHgyT8j6e
mEpYAE1dLERjI3PDpnueAAoG3/MoX2rUGMbobcg1kF5Ug0CCyVuti2IsUTNk2CH6
UP4yANi3FZkB1QJahmOODRLk42o4FepnhOJShCXNLNo7CsQJ7S3H/A2FML5za3uH
8toZSGPVAJC1vS992/HxYRbRWkRX95FwA/NzFGJWofY1Q+9RTaM5Dk5kPJLqSIbh
5CZ9Sz/XuGxS/5WQO20kYoqQin1O1H/JAeEttY70t+3z/YRcy2d79M/cfSzvgjrW
nN3ha4mcD+vxs+eN22xf1GxoxG0ImOYKmsLpwE87ByL53/G0pxZNm9qJZENmBapR
gMhC54jdp0tYzWoKz1fAlHJf8uZnL22ePdb81tg9hBrNBD10wFvr2ZJxaUaQPK/o
KRYWxvZmIukX04eVg3jEBDhi7IW/Poz1nMJgVKU/wYW+5pTRp6weEQeMSKGqKvaG
owG3/rjKbTf/EwwVFJalgdWnCZsnL/eS5QjeJRn2Wbh0mtydhnBxQPMZgMdAVAB/
s9YYGMJZO9AvzAjDu2MWtPyWj+Rxbrh7hrXvr2Ztkv1pZV75nIrOtPW7Jf6GO/EC
QuMoyk8E7zeowBxC54bKgXKMee4g8hxDyVJFAxjkDUgJKqJzTkZbhnWwdIsgXgWw
3aNZeKz9oK+yNrcEKHbKSkXt62QrRLbjRIfpmWg85V4U6YJHx3N6FC/fI6TGQMXA
YGVoo0rQfHheQCjmMtwRPfsehvu9u3VbviEXVFjAy3wv4mpj9AcwhPArdOpmYP3b
xLirTH6UV6pZ4ahh7tk0NwVBz4KdtMfcOhWBe1Rhc7jv5/NTlbjFOUY/wirTqZU3
v7J9MZs9ytfsbYVYCo9wL3lnAmi9l9wg2OJ+QoAdNuaPGazNupiyh0kNNQLpXvd6
N/KA0j+C7Rdookm6TalBDh0V78rpjGrNSK08xSkf+62FRLfIpvfrtgMpKzCMd2eA
GnW7ziqVBSY8lfNT9gKa/k683dMZ5tTfPGwFQCFicbUsa3q0C8jK0abJqBQ1Zn/q
ZclmxOf+rKXAK5dnFWLHZBLuwk86jfsyMiBtZI+A/X4I9RZ8W0CyMW68aI3cZHyA
duKzZDj8xIlhJ+Qa+3aVK5NpCMC5ssD87/s16Iwqq/Sg1yDLhpWjrZ4gwflcqDSX
8T2kIwQJGGRlOAh/rRNkO5EJF4hqlDI8bdETgevH8KhEMRvo3k+LiAUrBFXq8LaX
`protect END_PROTECTED
