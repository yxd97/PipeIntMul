`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qEMrzJpv+nYxwrq0EKMdOgOQEzkopF1AaqqEgMGyxG2zk1UAXQizY/DZBo9q+BOl
KCUB0ldTxE/Sy5W5Ftx5GDGEand/2SmQ/yuqjuwhTrdhB3zJ4LhqPT2K7wn2iO3b
pUy/ue00Jj8lbrgvYwpmgoKhzAc7t/n50M/Z7juhLqkum5y3WSaQ4wjzH4vFuecN
Dn9zS2IvOOwT6irhuXQx+bHJQffMzMdEG7dW7lY/0MOaer/41u10ijyWVBbumzfk
wUnepmVDKMB6I88uzteFyiKFlJ/l6QgrWAr57MAF3kUSBMcS7RnKm5WIsS5ucygS
Q6d8OjY3QieubIE/7ihaTQ==
`protect END_PROTECTED
