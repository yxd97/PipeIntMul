`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gL6Ors/pYJ9NlOebXFH5KEf/LvG+yOpeXC4WrXcdGNck5jJjDupPnBaociG3SMzu
yM08CVDyEFNztQ3UmOMX6zWcv0eUD8y5dlAh4JO+5reAEQrvEvnlFz8kjqPkpGgI
duvM/rWukK0SY9n2tdzTfjNLHWmaK+bI1VjfglBbaUf2/dy9KpSvslo9i4sIe6aq
X5mxQ3lSR4v8hHmSgnvOOS2Wq9XL+93qKZHu+CWjZIpEIB7Zf0LUy6Ury1r1751l
jsaXzFT3TC9oDKONKNUCy/khxnKYKKoQ4l4JqOtD/W/24LBQJpoZpL354uVdDZ4x
zkbSJ7YrGpT/ob/nCsPbluWmjbESmxlnakJZGdBVMOtTXLArLAOe73CX2SwTJr/Y
kprvnORob1XM3qYpw63ICBwI3NJ5DFw67OPrgwTb9T3FMsC+aPi1iIlESEtoJa0F
gOEhIeHWpD1tJQpeL+lvqRAAlvkQoVsOzIJamjQilfG39blhEDE8xBPxD6D9nzG5
8fwMvZXKZQSFlQnI9vs+HNZON2zil72JeXX7duLCBVKvo0Nip0erFDSFa0cs0Ppx
anG2/X9x0SJuFaA64Sisz1GNXQNpsurfMCSCiWfofycEYC+j0cv/LwjgdU6/Vaug
Eo0B+9eBS6TmC9FXNVUesQ==
`protect END_PROTECTED
