`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsuXyqnwn4WOy9+gTtl6MuX9EtVY/wts172ZirXPWCbgdqIc6/d4qng2cJYWuqki
HFoQUA8tCvkJdjk++GIPGaX+eh9VAIR31z4WmqjPJo5ZZzrQO5h1FGo8iCB/MTwL
4sCtja4yaLZXBB6yqp20k6CDMH4jwP+nnDbvl+/Bxjh/Mvq/EXLqmLXt3P9t9Trt
kDDR4WsoC+GoLexBCXIFyE6UPeVJbcBR41mKC1wqnD1d94FDKrL5ZNjO3t80og9Q
19FjHNG4aZGXYNdkzBIujUeQFUJgC2kJiGTS1W1/9UuSa1tYwOpEJovbBz3jjvBy
NwVY+mNzXTbcE/DMtOPc+AG7qUaFwvXTu9aF0nW6lyW4HBpZEi+VVO8qArzeSazW
f+Hi8S29fHEa9sgYt/qkB8smsmmU5R1R4MgucPbW7uFfKUFUVQoTGr8qzuukZW2a
cycM0O0x1EVl3ThJZjccaho36n0LRrDFsVqyKD0BwpLPWRMGrsJnYiC6T2XSQ8qg
YkHDL/sbfeyfcLYxKJaY5FaFSqxUiWJFcoAY0IeW00NbHSHbQbOSJhDVYW/xjx71
w/KrN/j2wlOMu3UEyrZc9225Fi9cO5laF8vhmO70azrF0zuPEMMSREDtL7ffZbwA
YAvLjfZZ6bPuxmgid9IcJMT6dbIr23H6SIKHBtwgIJWIqiURn4o9Qz8NKwJ1aC0/
45nJEp8e89wIHZJMVszuVKPpp6G1uZ7tYntS1TVrswPVWE/RpZkxudxKFb7SaHW9
WeTUZxTseqV8xjysJTaPymrfxT+4m6FlQ3wn89DG+CE=
`protect END_PROTECTED
