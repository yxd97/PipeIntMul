`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tr4KxiYuMUQm10LkOC5xgPuUxYkSK/pq5t4SI769dMBNjVq06BJ6rdc1TC98UQM2
GiEygGJjRePvt0c1Cau+mzfX1VMySH9wC9qL9+cgGoNso5mBhCrCNgemi8onWTX+
LGjg4ul1v1VrGpKjsHXE4J2vrxSetm8R+sPJtRudMzTKnfYTKzTvVotZOwv7pQIG
EaeKt0qfPQYFKX4ENBYYqM/sANKM/9nAkFaZkh8+qTAmVgUijl2fTFVhgVsgihqT
LBpDavAKndwB7+Ixba5SGSbgGrxSkXOmmEFMlqUJ7KEOflJNpL3HGD39vtVcLAAS
NAbaRS6RRPuxmyLf2Bq2XCQEt7WlwqLF0tOr85PZg5bwUPuZEjSxHwQ8sJCoW1Dh
3iknls8qHDfLCFbaFNpJsrEfC1T7IAA8pGi4z/pay7A=
`protect END_PROTECTED
