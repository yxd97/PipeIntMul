`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGXL7u1GUNFkeWtxugpWYpLdQ/zyA1FjfRlF2h5ANF6jpnqUhUWW5JA2HTdZrb3N
MT4k49BK7M44rS4+187AzNSnSA6Ux3QBikfQ4IrJyhU74tgtWpiSMVgH2wFiZLLM
UmZLa1ACLT2inxWZAr/wjGGuXnAMDyQu2OawbWwsd3jG/jiGS0vozOE/nPr2Q/0c
y7p5IkWZ98xWJwybaRtONNKmFOQUSUEmfZszDHkrMXXon1WT4qPYoPQzofnX7do5
2BWPLB8RbvuiVB4gJw+h8613IuB9oxYii+2O2sB0w1ed+wb0O9Q+3OwFPQBySvfg
GX08RYoF+m1MlAWMl4EJCg==
`protect END_PROTECTED
