`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cK2vY1xgYCu7jUiFeP7UNi+voutT1Bn50vNBhUmw/Kpu58O3pMk0JjWtJoDkDDKL
s2h623RXoT7BmGnABAAlbV6piTR3ypv28UQxSYxDiaVjiwnP1zawFvNCtpT2uVvj
FbylMfjzNaLmHeoJJ6kSjFtIs/XqBPdKWfP95YIitQLbQzu7kex1nDPLwjs1q+B5
K2WHzYC481wU770Tsrhp+DbWUs0WzujRwOtrY9jXBYOrJr75cWVKiIXq9Sf6crHt
F+r0cBEUFICChAlX/42CXadA368wy0q7hrBepvoYGIVOzyq+OIChkavCXLyIKWtu
d/dfpbiQadN9kwQQjMAtpf/GE3/YNJCohniBWh/kZEJhmWNWTIoaGtZyN8cFjmXr
TF7ySNU5kSbPR3XcpDifx6HfZ58AWHJ76ceC+EkQwVd9YGm5yrgTZpkyxPbQ5e09
0LrYpfTBnUI0JoMcqECddk8l0/lDwrtTbQJCteTOPCAcfBzeFdaOARmumvIU6m/P
N1ukq9iYlBjn0+DVayWBojMKHkUNJhAJrx+KpbN9828uq9M/Rxt9XGyK+cbS5iO8
vQVSPw3fruf+ltJEinSPMuiRZIbKesTTqiQMo1Ohpd8HoizXzphIWjuLE8Vif1Yj
aRGIKARm6OU5dJ7CX8mt6Cjk9J/TPgrIC+FGet+qsX7VzTzcIBMS3rUkwjk6fVE0
o8PhzTR+YehdUkR2OKqRYLmBuxtfldC+xR6rKJT6TdLYEXm5/IbaWQckrBunXYnX
9/5TbGJq0rjfCP3Qqt6CY+IBdsNQw/xmaMpiE54crCk9skxWq+C9yLlQ14NWUwa9
No66udlD4E9V8cRA0O8Z60II4kvVcEt0um5mfZU2NhHjU44cpcpbcdtqcrxZLPug
wU+fabwcr35KCEJuvjHOvMBOKbSHg+rQYAX1OE8g8PNuAjHN4erIOaBFAMOjebYO
G6khMOI/D8T7Nc3aGAObG8AU+ujme4YuC8ocOnTWjownsCcreyUtsFcE0AnUX3Sp
uT5mjy3drDSXuNAc9PAHdiYi5Lu0HcUAbwBTe7pB1+V0+gD0LrP6fv10NhGMmNg1
kOpwf2fbv2EaCwhD1TcRIEHX4E9nvCWfowujRw1hLlqn/HipWA6Wudrh5nPMViNo
IqP5/HmLlZYZh0RNxzoqVl1ysfJlnSOYZYcfrJSz7jOYHlSmzT+MuocHFd7r+WIp
nO//DEd67SWbg/w8fmwzT2ThDqUtnIL+1YkO6vkY8moQDruM/1f7Y0vH5HpAFUVE
jQG1RUBlgXfHtb2+HBM1Y+3MWpPEF03J/Gm6Es35tlynxtZo9uahi9xTeyp4xdhi
nEyKSoR7/jhdXg6yT/pafk/O2M2/H9Uzwct5KIF0udval00n8rMGWUlys+7BNEQc
1e7HlmaYT1OhdrLf6XzlzJfD/jnV4YvWjP5Hf/smft0z90iFiCaq81KcRHmiOLo5
KNZPixH+oxUERI2O2ERwjJsIzUmrmDnST+d0kU8FsTcIKIwVUKZ15SfoU/2PBmDB
XPR66V5JlOUO0N6oZj3wNTMNvv6Vi4CcELN1ujF39UnK31NB4uEDHyVn+LgDrDyq
Az6jIHSYhBYOtUuJM7+9T5vqLwp0j0V4/hzHdOi1RUxB/+O3TRI3RYhWdfIGBmQW
wvwXR37KW5Xv4c0NekrbTQNKMazFAvPGCAUTaEJzxkcrcd4M3PG6DkzD/1VqBDQf
lescE3RQ1m+Mn/UGn364+HgCHkBoxbDggPAoH27jhxPsw+4fSweOPT/Q9t1Tj/I7
55ERzml3ysxdA+uTJsaf9t+cj5fgzGgIZz4uw26RhMNd00wLEHjZDzy1IN7Qvn0N
6nmQXmYnA3AxRTmP+mLoP8yh5M8CbcRsR4oChXyBGW8makx2kwTsNY/AoqNN0m12
00WFApvjDVZG5P6YnpX3t9b2iVJTdk2Y/vkI796kRQmmiq0WHl2wad/vYCMVGrje
bBiHB1T2g9VXppBfvs2ZN0l1YK3rHpIjSksTfX/xlRjeUcbTJ+MSk8p/q6HWRd8p
MmECP9fWLkdrsHboEUFb+autg8Sbb/YNhrI1Cj2ri15Ejt7ZziQxCGQys+lWq+OB
0wwUy0xH38Wuq//9TsgXNHBtSRUhFsPcGUeGqeVX+ucysrij8SoOxVRGUpcFDHtr
T2IBvYHtHJXZ+xE1uGmIu8f3UL4RK21UebmLS2PsUDFrohafvWCu3Xvfl6Bg6f7W
Qqsq/WorWepXoPB00bYiPzZ0aPHSMcgNVwos0vCqxjXS6zi0OmuT9vDmWIzcukA5
WusvqUxqNM7jBiMHwjHiBtlmZ4E5fRtSmQscRYM4nvrvuTruH7e0P/SNXrtKrhFx
fLfSeqfh7yJ/SX2fgU568K/STNefB4McO6hO3G3N8CZHklYu4YOR0gV/k4SMnF3g
alHt21rDVcPS2VSuylhcrnSM9tzLmP6WAFDtGbojPvuiGJq5cDycX7RADX2vNdnW
0qz2IO2XpslI5TXFNCg0Hu4EDX5OpadgVhzc7tY2e8gP/F2spm8dYuDQTfWAlEJy
NclRJCocWAjYH/zO2VLFpM5A7cQ026oAnct0DqQMlyPzbTAwC2KEYtlaUqFXnhTX
CFmwj4FMeKmms51tTEKax3twBE36/e6w9lOmGtjUt7Brq7jt+xdvFfdTjXEpsCqP
0bQbViZzeansZidY4NsnEx92RWRkwMyqioWKTYMLDmJ3lKiD2qOi/7pQhSxzrtAf
HVCraOWZPbX0sFOJCOlFKt0mFa8U4SgcyrgcN3gfO1DrposHoL0jC21Np7kqMJ2Q
KoY7LKho8u7artut9FP0j0dEi3izvsB6BnUF8KUymDzJAFtzn4MD86EHMkBkHfeT
KS83hSbOyZs41UlzxInXQHsQKslvlbtETFEuWyzB33Nw00Jxm2TlbYEqnT/P3o3c
0A8uo1iAbHAq8t1KrHHep0lBas4+SnFXaj3YPI9XHJoO0WdBmF1p0I0b3zTHgNE0
eU+f+mG+gMg9TWo5pD9k45eC1xNXjJbucHE6MCXauojmRbGuaD4uY07uZYgEHBeO
jTPVeNpSx3eo0sPVTda6OgBk67Y5q67cy1i4Alns9WI7Zk2OwOJi6OCkK3rsJVmr
qRek5MbqcLTw1v7ItPj8QDszSzbOF8RcCsMZRpkiYryjPTZQ2gUuTnoMXDdcCTOy
zqHvalXgLehMGBdTrx5PXCrh68a5xG9v67nGJnt1uo/yJlaLBxETUX5rYGvXDPpI
s3rI/CLHRf8Mn19jDp08DXBAzoxQnwDUeXkciRTV4abNqYdRkzQwBOjH9sruxTi+
OtZ24gDq7CmjJPga3WHhndw5A25Gvl7UQK7wiAyYlBpXnw0mOvJzyu96E1CKOFgZ
wbPjltYW4o1XD7nco3tN4vSC0Q2d75ok2eBMhMUHWOp3tSN90izQpDkIzIpOdGJW
skb7lOalYKl1bjhhjY+2E/stoaqeKAKhp5gtrp0F7ZgSeNlH7nDba0Qhpg2OgDZc
u64w5j7jkWBu6CJgMm179yx4Vo0M5hPIzs4vOVqA+DYWBvaOs4UgWWQcKI0T+HoW
VNkvDdmiQ6vZygCcpURckNlro1j+kL3mwx4Bb1e8NWBHSfbsHdrtULZlmy/RckSP
EjKdyImQP7BciBae79F7IW4YxAJB1bG9ESnYEbO4/S+4Hh0qV7cFwIAV2udqPmmh
zJft6F/NWTOLRdEOZrwjLdOkjoYPfgs8Pht2FQSO049cqYJ3tYQBHlSQKcEMxGOL
d08P5u67QHQsLxyxrDXWVTQ1RK5tvBw+RMT+qH+LDzH/j1yaBH9BE4mPENRBGBIE
toQmPO+Q2tp+oyKoKfMD5mVJw87DPFal+mDsvyPZWYrMRCcaw06+r6xvbVpFB3Sr
Bv9KF7KvNN1n2GNgBgOImfUbFcA51WTWj9yzkRaYinFOm+jW1hCMcm8k4hq7vbbV
uJS8Gy1FiLf5ePga54+j5WvVdU0FdJ6df8/cUpPAK7LsclOf6gN82OH8wlgGxDOt
Yhcvsq5y+up1j6sudlqbtzV3KhS1hRhcH2hNpRsRFGYJ41gIHFSkbjHAqCBsDoa6
Oc98u9/CaBjhBNM9Ee/fmMJgtSukaIQfKMQdDBnSRFbIC1gwVOyNnC4mOK+QvQN3
O++HgOUWyrCmiceKATAj45JqzKatqhH7AsiLlGoAJt4ipoHvcTnpdAH+fYMB8NOI
7diS2+9dhqAi2txk48c/wuJARuBO7g4/eeXnmzBMLZHzsC29i8Li8F0TTxiKYtwy
WHS2Hbm307H5hwsKCCMAxFSQFGKCRpocwTD/IOvvbYguEbGmGNjqdwfZoNsQamTp
OcNtvuVbxIo1jYkkc+wJBBiGumtu0ECJ4yGSCyx8HQ9Fv90G8iUCnejnVL4GvjgM
ulyh83Um5g3YKShk74WN3gxJcKCk+9NvbuYaE27ShC7UCw7oOrzr4x/FQ0GZVOMe
kQKOSktZyq0RKOZdiwpsTswb9meuesQiJkUzYO/u2cv5aZn1KaKQJdGxCGU5z5Iv
CvffDDdvquAJVe2lhUW6pFs7zBD/7LE60bzg385W4xjbIO080F0YTQ3ZptnyxAx4
S77SQw4wBHleUs1aCrkc+FfXLZF1D2RrUjFDzOWhRXFGjtsjblh2zhY4Tya0ylAV
qsT3Z+xqMFkMfKiEfmODNJ5l18MXQQXdCPd6iIPfJaDbo5g9vgJFE08SaQt8mzeT
OiYz4Wz+NzS1RMg5rBxGBKW1PtrwecyT1DTVTOUXeQqA1wX4O2UkcmUTsy5xKctm
pedwWUiHRfdRmZ6pN0lEaBh3JAT1MJacImQpgMHBQGkVFyoJUzRM7Leng+tfrd9H
u9MYvw16WqmErz7591D8siaupN8gyba55hWmL1Fl6m0BF+5Wo7KHh5PcJD/PESGq
Atzdul518hZSg1KvGXhx1sW/rLdKSgJ1MuSO9ax2YsmO80WY43vKY07nzgNy5qud
XaNts22c9J0p+1umO25fEKeYijGXrhMMTCk9kuVtsa/x+PI1xf9d5stJvMLcYv2e
29CYGKoPTRJjK/pMHXkliRqA6VwiRo8eQx2TWdlNLbNgpCQ1sbk6TVnhPRBfjpor
i4NFiOlWpSSVERC6wnHy7QySnwXezGeaJCL9jY5z6IZQT8zBHTYyizmfe6hI7wrm
s9ARxX6jnamhGsWfCBeigPKYSknUfL3cnhlq2XH4mGkPgRn6OKGrSa+rXc5Tbmpo
0ZWMubPTvdpzbLIlzUG0edygZSI3307mA/cI/z/NuM7TD5wLQbVEcb6jsbDT9cVB
skTLZWS/PJUwJ/idUHeOWQGIKxda4SmejJrdKnvxRBh3Usz/hHv8qOtlmchiyzyT
nbYYFmrpQsgbCrlQOEdoPSF0o1zY+seTmbLPDss5RCgOIIFMkt89SG0aJqOFSQeu
UukEUBG5pHI3bC3MaQm+9OZdUagK9EHN26atuGUj4BCG4+K8ml+WBUsyTsmc8HZb
qtpOFCfkK1M8hMIz0zqPdWtkJlai6W3MSVQ5lMsxDX6DusImPUdnjlNZeZRdXWUz
VEVF9nm7T2U4xfdHhNLqOc13M5SlytPhZz9SDkf2uFrBgbUXIeeVanUwnTQlFNZW
1laJ4IoKVSpw7gEVWGSObJSvu81aWor0UVZvxiNl70Gu8jYNGzpYVTox0W7HYTr7
yI5TBt2KPTqrDxqfL/BYTb7qUtyuFExei1L0Wcqi1A6BfPrLyKWVQcklot7e1Aky
B0JsW81oFs8EQhbnHOOiJK5lBUqTICD2/IiF342ZyNtmW+yug7IoSsemvQEFw9kv
VRq08QaQOJ9/yhcaEpgjOIUUxTD9yVQxskhXaNEG29dxR596akZQlUw9hXDF4lP7
NkctFa6+VM0TJ/GNiKYx4xoHdn3zEWAT5Nu1ygWKzTL2JyUelGK/wZ5ivhOoVSi0
y6kSe+JmQ0xjz4Jw+mpXkhhIrc6b3iGFG9uzBObeWVcmoYQO7XVt5JIwdQisqOrk
Js4a93NTBygqcwv2DYxo+seRFCMCbZ+X25DAqRIhRZjUXU9HbRb7plRfJ3x7ESuU
1UCgpX/kwmAgLOi57mNZaBsUAgQXzdImuwDKIPMTNxDAXD5RZRk6KRIsiMP4Q2mz
SY4zqNosd5Dpe7Kxfwp4B8ZIPpm8VSjFCBYnxni6oSM73vwMGbHhm+39m678Za0S
64ePmu8qXSTuk6nZvO5lQ6Jnt6pq+1UzjBAalue+qbqMRyFJ/ojCTdZWbNbW60ZH
CddgnZHup7Jwn3PUFnetpvvx1yC2j6iZHRTrG7KXHPV6g9DD/sDvg4JmF7eG4oSM
qnRX/m01V2mRXnMgC5pdJaXF7vzxNz3zaIcaOgKpA4PU1QdMijxSC6N/WbuA3CWu
pFhwuTdRD5Lh/WpjeKNIaEbvnHmLpovu0huYtxcpKN2GxzJ06ksXWTVaoeJoczKt
H1rmF74GUCMBh7NAucqFPamawTQub0sy5y0kwZHO4DbZemKuURLNQpZjzfgcnwM6
Mia5FDzjuTpxU4pNEHKjw9XCOVub3GhsrxNlyLmqoiq0zU3JowdDlzMhKlUN/fEn
6/MvYmoFBS5EGEzLkaG8AnljQ3ryARfX+olPF2MBQ0bH1D4jAcZyhQGpCt6PBD38
2NZAsJS6k7n67LSTX4iC97dQoU+AYWNaY5HtEyJMMCOqTQTs0xxpl3su11DijoFz
jWH1tC6G5QaFlMcA3PNCtxV8oKFop6e29M1dH3JW8EpWQu5G90yNCWLFm0jmHBye
nSKogsz1Wg26zV3HbZeH70cm8GREZe12eYJvZcxcvsP2QqRu/fY4EsjM/7gFc/Kc
qOEAxPrgxWx7zKr+WFW+Milx/z2aG6qo3HkHdHj3rWXrVDOVaKpUxPv1tsgvvXIi
7x60MLxJgaCAM0Ue6tIT+XkD/oFrUbAcne8mdP02cLvS9XzJBjgQqO861iRIDfzg
6KAE0b0q2D6auSqToehJnlLgp4cqeowU4J60TKQDuZw9urc33sLIoEM5Bw7ZFGOa
DswzDc7/yvgrqb4rbw6OO1ULfdx5D+RsgfJCALf5kSSy0wZFtSiGjZKHvfwoPknH
IlV7UHZx6wFFmnTNgjZoYPI4xQawfRfOn5w77fcKC9O/UnytbJb/PKdBJUE75ioy
Rm59v2XvwE3ojCpW5zlezh5IVK0Dr6+c2VgesSTQyk9zDUeIsPqL5dcbEcznjGKv
52EhxN6R0Wm+H1D1l/JqWl5WxxCAirfgKCE2tVzdZYSZChjKTiAJ7My5YKnavApt
fv8nAXwoXK1OXlSHIVCKldtnC4pQRgrUWxHft5UQSl+bi9pVCNtC1S8rnJ14YOKk
/7qNpVhbkC9zviw+byhizL1aIY/hgl5/1pZ0krkr3JfYEZoOwGzrdZgpxZfJiNyI
mR3YcLJqUmQtkxqbIZr/oBCDKbsu6Ym1BCPYqGgYGp4IrOw9xlZstTspp+MVicAm
cua9uiGfsXMCMxi1iAiPqHkwXbE0DJ7EKyXM3MaQafazud0XsrIfHdtRLBYvoFAO
bIfSAQk98UcEjcxQAhND9q6OxQho5EjIzamWmjPFIQGSTLkMEEltlXGBY+hfx3Vs
O8hOKhaKoVHTwREDlm9tynszBy4oGd9SriNBVtnCq9um/5XPKVXNo40Qu4FgGjpE
xvF7biPf6klSSGY0XkbsgIAH4ZzBQqJBoj+1fPmk/F2aJQAr1KWiY2l/mPC/gYdB
YX+jT5NfOrOGBtqRjDTYiN68fgwafHSq0G7eVpIfKHrK8Ld4xvBh8GWH5HlFTymu
o+tOpmFmpHlFFVedPjwVaLXW5U8jVc3W5Ovz7C/vbpbp9glcY/tNGx64TVAzU2Zb
Vo44ZQxZ0BR+SLFYy7fZtuxZyiUNvgL//47O8y0tV6A6UJ24Fm5sF2doGY5NttGB
wJVd2C9sLE48ylkAiU9tIu+pY+mna3DbSy8bKmgRxiESI0pjefsTxIZQsfB4ICnD
0iQAmQMjGAI60crfA3MEAgfVQCw+ke1x485m9v1LmeuiehzZL79tEGsQ+VZrUY2S
FV2cm24l9bf2eT7V/vR/VA==
`protect END_PROTECTED
