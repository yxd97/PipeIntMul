`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRcMuI3zT741neCPej1rr5qzi5Cf+C3cZUkvxt77E5UsH1zYN4UhM8TTM1wvybK9
0tsUmjQIUMlpEe6L6nhuLCGG0oC6BxWiHwjSMDAElfSmeqBSf1NweoPSziHahG4y
ZMJnUJB1VsG4ra+7wJEVrksXE86QcYUnNKb67+SiLF488fkgLLDzer0IXQ0xbXrf
xc1HroRszKE7e1VFE9+PA6VYYtvkU3xnIwHpFvIoruwOb9ESVGIZGkY52MI1C5/B
g30I47Tl8cK9Bok5GA6k1hnI+dVg9qn7Eq2pqnWBIdT6UIGSCGNEH23/QoWIWg7Q
beAJPw50r8hSRyVcXnqGxkBGZ8f6Hrjs3yHOJhvkNQgsS/Eu5WKdfUKNXrdCg3PV
oePx/0eXkxfJV1cTxqMDiB2aHu56XdbVIyGms0HcxXvAKbW/tTPZqj8iLT/gAOiN
XX89KjUaCIP+SmRCbhgVF6OvA5AFhcL0CQjV2k5IgLb53rC6S3q5QnA7bl+XuShx
+WWkOzfxHRXIVKQhEANiag5xCTgB+87NE0zX1dZgRghcRQTb+Xq4cXgzrQfIghf+
AWyhwkuVKnWeV8ruivbMp4WUrRd4nWYeJ6WBQGG6G6ct/eGrU0DitG7uRf3I/YIT
xlqTusaXOKcHbWzyynjpmYZt5v0q510aISiyf8bHMArd5DrY06+iLdAQVp0QXr4C
MrrIEZJuyyvEOBk5Awc3Z0njndBohsfF+PiVFJbt9p7H1RqgQ6//DyHNNlZvjTPG
g9b5J7plTp2LfCQm6JG3ELHCAW4e//mAWukLWS1FTHfvdx0upzlZG7Gf/MuxHmaS
KiY+XKbQYH24kELQQap3vSkURflSIFc503uQ3Uil8FHA5EZh6llTa58Q4T5BFQh0
J+ufRK301vZKJ8OJJ5xe8AF2ZqLF8jMcYqKry0cTJQrjLw0grRyptAVT4fgHC8bt
`protect END_PROTECTED
