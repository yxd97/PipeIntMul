`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWI75e836ISUvTVeGitBtm1zuagdRPkPzXa4ihHiDZz3HUswmEM/GTrz7x1P2cxN
1sCYdZHNW+wfF7W0UUtER4IyCe2oFb/8ZG5ykExi0M98GJcB9yGjljCjTxRXKgPV
t2zEwDXY2XhO/oLsfNVrJA21BHTu87yZ2plU5AbVME7XcgmiqwsODTJNXslSqP0G
Xo2yuoxOTWjbufIqUKwWRIsSKzlv3AC+tQdyVSU7akKZpqyTFI807QlXwwrdGe/m
aMj51eqOd4sdA6rY6gVZkVRYcqyxN6+fLCxQPCsL6x9I0bx7mBA5MPxh5q0j6DOH
p/kTl3I79lRZwXHULgPwrstKRqBMvZGrVms/S6I4FYL1p4OjrhG3H1wKMq1Y23p0
WRv3I9nn1rZMB1CL9SEi07iS353Wffz253B7KSCMj6t+fH8ai6XiVKi9BfsrxU2/
p4TUE4OL96aBbXJLU0QXvhMnTJQHLt2ooJqu3XqMEZ3CXdSbogxKgYh6bzDHYvFt
ch+Lf46qpPq77HZm+xxInoNmy8y9ABuzq13BkZW9L/OPH88hCh4i6qaR1sAJ4gu7
uAzYUwikDKkByWNFYY4qS2b4yg6jOxhmKGyCW7pquM4fPMSlmxzJqWDjLu07XEDM
Sgod/BRynT3qPwgXaK325UNWF6nSeht4VgKYix4NRTDksFOQ1fxw8nkPQE0MZY1j
DvsIewhopLFQIbKebsMMzikmVqYueUw0v9AfCyuXsGfIyPDIVIXeybcHRbnM7kl3
YsZnZirmYvfMQr8zTbtLFg==
`protect END_PROTECTED
