`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
go/Rtcls/jp0GWb8MYlcY9heBlDkuPnvVBozaD63TdpfTZQ7HDsxtcn51BaqPnb9
Ht+WxBpsAdmup65M1FRx4PW820+J2Dr1SoMH4q9QhhfvMJ55gNXuiLwM+5iy6t0q
jitp/6gHxoPpoVuJPHuTUTaYJZk6ZwSPG6LRj/cDIv4fbij2cIH8DooC2bHMxs4P
3Zo8Le62+YVa1dpyrksP7q73sOcqGSCTuyBw1in5bq1EFqCu0TdHAEZ4i/rhEJ/6
JQnfWG2mzmhKF1gz/PdWVe/myWtEZCEw9FIkKRs4hoepjprOkV6cNzF0884obOHN
dHIveL4ekxE9pYlmzHduIVLZrsvH60Ibtb4HP7vbpRFr6eGeLyFPtAB4rCCanJ+q
RnILB3YsgCNNuHaiXmvJCx29ULQaMd2MZjMrfqLF27bQ6L1LMxHDGQ2cKCp2B3MX
9IG1/UOuoQrd466IUv4yw6wTEXW5XqfdwnQNMSAw74KJb+ZP4tocXLdgYKcjJNL0
kooWKal/NCiC846rqAzvC5jgXsSzy8S/RZ2sWYhDjUwJmFawurucNKMogKwxGzH7
BdFhmRKwhItuPS2DdZdDhu982gELk/TLBPu0fJVBG3YUIix1CW7lamGytvXErlEH
`protect END_PROTECTED
