`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZXMCLL6JRYijzYtjtXHkS6gX/j7QeIIMXxrkupp1E3VoR0lEfaBlKDxbWJZs+fnz
wi6oMj4MagoDF9V2LC3VDcvLLSKenmk8CI25NqKmmUYDxKyamkWczb5BQWIDkwn6
2NnraDpnWeNabGQrRs9hWvvfmO50XVnb+GnAlUJNzMHqT/OXWLlgzjHWlUhUY/6C
ex0JRMSdhRbYAAPWOtBNUpV946CS9GB0fR8eYwg5hJZIJU89jzzPGCTdcnHoVNwR
HRhyp048YJ75SVP6J8lp41rWZNA85+W1bEPWRbCl4MKRWLDrlBkGwXoKZRU9G/37
tTJRqXl+uowAd8ToN+8sklxhH/soQD9KkTlgGCKJHNcLxYNsY15qPUn3UBqKKwi4
WlFWlqwL1+mP2aELuunk/y5DH9nCXqdbGDwSRVgMqsEGCCpfwOQojV7gp2/VpDbl
DQ0yARACQh6s3SWbtW4plL7nNB3jmLxcOro8FKcSxqDXv/R2qn8vpejj21tEuo7g
lnOCs6ZpQtahbEUos+PimlW9bRXXdtxRhQ0rzL4cT9iTpGpXerowIXcT2GGl3bQ4
07vn0653X6EgG0m1IPsl29anUMpRyVT9QchpeAX8i4fC6t8M4UM2+WEZinV38a7c
QEjF0Xyn+/1JCrzxqn/GOXrgJyG4dq/J1hOKLfIfgQ2JM8oZUgz8lDEtY/2eymHM
+i3TgDNsSUQiHtJM3PGPSQqhkS8j7VSkTq7/f5y+xDSNdp5XPRsDlYNQuZUdTSkJ
OSebxAwliNL9TLuCgre4kAL+7ru1VsGqQ85GHoiSChHAflXRH6a286thkiR3Zm9R
oM3qOHloSVMHd+jtiYII4rhiZgBjtbZs+PUNrJ8Zt955P9+Jfzr3Qfm89OlTLdh1
0ceFhOgxQZJcfEfGn3SvECQ/AS/k3lARMOes4Yfgpoj2+CNQqhWxiMUrsVF8JMKN
RGNX3xGvVVJg4zNmqQyMv83S22TD4m7vkgIaDwUodSuveVBcdaae64pIxIjk7OY5
NV5ecBqrvWjpgDi347YcRM87cY/wvT9rr0G5B3D7uJc+PfMpY50L/nhpXw5F1MOo
qW72AEqlJxvDV3gH7uUSkNso44WCAnr4gr6PuVk2TdBeAYcXK1zYUV02bwpBhBXh
`protect END_PROTECTED
