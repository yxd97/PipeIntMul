`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TtVklfviCYEwVhxJ5myKhOECRubGsZiFZZA2FnPDaszs4OwOUvbHOe4hbJp0fxBN
JMMV+/uYp8/NnMvmyr48so8xzf5DTHHkLSJZbo550Kl+Acrc6CZv9TcR2l9T/2E+
nKiUxcf9cLhBebAzGDRR8b7XUjVVvspN2CtUwotzkS6iYnL6aw3B2nagDrs2Sq1S
IJGFwU6i06Oh0B4Fq/SpDtXmEDY2ZB7MNZWWASn31lL+8h9OUmovlsh8lQhAmZfU
Ta38C8OqBop/QzrPKcKXK8trrNtRjeTs8/gDqqnnF6oavC/6V7pHGyFzs2042DYw
QZt6J9NGLeYR6kj2Cd9+C3iHISCONABqH+bwfGFXFzlS59z4/KSjv0vCI6f0G76D
LlkIhZH2mtTrrGPOO6n8v3yYmnqE7iqywMLplA9W6/auK7bGrln8Q9cBRJSI851U
Eque/uj8NIPGltqWg+lQAuoKBU6O4IkykbY0+2l1Qu1TN7wnt6FesmF03riuMZny
Po8RlheRzkV8YOToXVWlg1V7QhHXKw3aJz8HTmhikImmli0Hc9Wi8JtGhgO/+4YY
JiU6EXnyYUm8vhlScB9D5vGHBusc4N04v9pZ/3K1UZCG9KaDOrH/5SnuaTMLRkbD
D5gF6ES/P9SzOiLP5pkhjGdoxljC6808k0rRv46Yfx/XTn0HntGH6aietKZNoSC2
LX5eWU2GBQ0qHB9dFzsybA0SDjycI5hrit+o2n+iCrdz8kv8oDzAfW2oPTZxfBTO
fXrKE8+kwJvBQHuQ6gm3d6Ak3DmkW7LjImN5/dEzp9BTZkCYInYMb9bKRNy5Lq6d
KbH7eOyT189hNnz/qmDZGPn1rFb6mL4KX1m8zWFFSB5azAj2GsGniznaubJBZc79
wCGnz21SFRdUaE6edAjILkVbPFH5dCOJIsaonNpD2aHncVrg5DVBsvZ+HFL/Vcte
`protect END_PROTECTED
