`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cpj4TZksu7EAUXTFlzDgrA7Ly1gYjEPj1s8p+OtahmELAkwmH8h49M2EgBU6eGBK
MNpukbQSPIrsRhYaHfYJDXitaGxBq1+s756i4K8pqus7cKU/fA3vcdN0WWqowB/c
wk67BracvE7vjAWC35jxtcJvuRzyN7OSuTtT1vkZJqnujAxMzl8doMKVShb/FNo2
U8DKZKXQwMX23pnY8C/597n67pv89z161abkQRL186I3hwpyNY04D8pqabQiqGSe
Z0s4m2C3KlTGeaES5pJvRHwtxB4DvEDpPxHFPL+3qk0eMUtUw6MZK1O5bB2PXNYt
9j/TEg2/5gxiY7XzIJRUwuAV4Cq6Q+S6x7u/XPg9TVCr8Qio/khWsKtGWXMPmB6f
3Uz5epkN02KAcL1yx1j1aZ20+3vbCGpwwP7u00F4IFuUuMXK8lJujeOC6WXXhF4B
4csXMlmJTlHjXZ+sx1QPVA/RKR6SDMR9L2uwSQroHVhy/hZLZGIyzQ+kkfQK280b
YzU0SAd5RmAQX401rDEm9HwNaypVCAmD8ZPwH0HDzjf52k3LMMjX/n/3YzzdRXyy
Um47kq3Xvi5Ie3v7rMbTCA2Xui9SMjRLOU1OIXBSAG6K+nS2GWKhjRY9VVDB4y7R
29Sm4j6uA0k2nijk4tBfXytG2merw456B65GNZZrH84R0GU/QhHlp9UzhEBL3PXe
CF4twLBKAy+BlMTiizLwndsSLEK1r4zYeFeX55VJvto=
`protect END_PROTECTED
