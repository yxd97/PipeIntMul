`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w81Dy3i6Ce0vhH/k4PKgeScH2qBDGl7+yLaHw3DU2APg9TmyeTkDWOEVH+t/eihm
OVnukXW6dpIi7AADzbZKy1NcRtTh79AUDG1OUS6GadFo6G8gRjFcbZy75gtk64q2
FqKxAhOQcT8vkKnwYNqBgV+txpCWH5InNqSiH/0wRld/nzByELFGm2stsF3LN4p2
Dg55dzOsvoKA7WJWnQ6lSgDA9BvEJ8yBnDd7NMd6cIlRuSOHl6scd4uyOoDeZLcd
IKBenadwuDWGBRpwTDAw8xU8MyP1zJlRxeZnG+KzyWBpTmqir8yGAFG4xVxQlfuo
Pl937GnPMcdQuvDJYgFteMWMt9ECODkTBteLzQH3DDXpbWuu2/74nj95QWa8fYl0
Z7VplcMHzRrNzVwReruJ2ooSu05heIvJ7QyXA+3iJl85OJIMK4ukFXYlFHGypdXp
5HSy0H9q85H0ytYbdq0/UnqsL9lQRj1ERCz4l0oJ9nBSOsBKE2Oi789ecWIg56SE
SLPvF5yVru9Y+qgHLhiWhHS/KoGjYlACk1V5LcW86ksDoy97cg0LH6ZAdI0gStQR
QKVpsngbiR7yNJ4ubmaMQ2RAGs0DOUQmskQi/glYdLiAf+ABZNMQpq3ZZor0KUH/
v8mA2NFAEjyIb97hqi88HE23xPRi6KEQs8mNpHcAnoXISQdQCDtrRjwb8t9Cu6nt
3i+4aKJX6N6NV6sA8eHd/7A4K7cizD2dgaaearByrhM82RmzSh0jm7qWQS8DDopz
aHfv9zWrZuRuOHnj0/yfAS89Wz/fOjsRPyB3KQH8uRZ8EgGAy2hc68g7XW2RXSIO
H4gynNEwq+Lyy6FCZ1tyES+zxtngkPYIXATvMWSq00R9m1Nvt0l5TnGhHEEp9Vb8
gxqszlhMjFonYh/ovT6BJg==
`protect END_PROTECTED
