`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INXPfUa1nfdRbBlXIsDwz7vB357SKRAFhkC8A7YeDU7kqeiWGAmxI8LPFPvkdOiO
fOZ8ZOjpP/7JYgwHxS8KEhgcg2OYUVxF88YEW66vsJtVxtMp+OBK5Fj0w0TUErqm
z3L/47AbNtkaTPc/w2GB7g+X1ZcTGszoTevXNuylj605BnfIrge7Ejoe3R1DM0P3
WJGk7PuDv5XzT10CaXALZOW4dYno/ruoYBAbHmBOLPkJb+Y/0TCsWHmlqblJ78/j
FzDyX9gv9D9QhYYWyJaIeBCuuOhmwzeaM5OqjWRXJJf94/MGvxeErMGZNK0ekLU9
YjOTEAWc3EYHezX7g9uOjFDoikFENoLKI8U3rW1c7ZePoBD+/cAOuA1l1QWyQF1L
hLnaOYyrDbaMvtWJcE+G1c3BATLzgfBmH4Wkz7OlKzvWjo8HWdZYt+pfLBXb7AMd
oaKaYaOhgz3SREMH7WbSOJQS2paMeTaFpZx4We47sG53d03NuDZeUCl3KhBMnfhD
WjH0/bHZsmYw7jtZ68+oyDnBr3EkvK7wakoBmpO6bc9mNdxV0g8EoLhmIW+NTE1M
7uAJ0RCx2ArpRxNk1e4qRJDLcI8kM6uZJ9fvS5hZKLIvqtUKk69JgDIZeE9mSd2w
N+qUrIqfnoCDLrCXjhGn/5RjwxmK+R7EXhs0OoO80QXl3q0eOVNb4O76id0gloyg
y+gbkEh12yIMOBhU3v17RbQ8vXb+BuekgpByV7C27ZI=
`protect END_PROTECTED
