`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsvjqhKnNDKQ+MfasYk6rIv4qra2H3VfCYg0/89H751I4IkXGUcdmCLzHUVxR2TO
6AjjG+sAJxPa/sIU6rCZbaMMJcg90t34HzL6HeiJ/pMr89WLFiyrrIOhtJBitefm
HgeYnxtCe1+AfNbJF3aA7rTJ/9IvvQJxlkSmzaAH0QvS+U3JvW7YG+ejkQN0gMzR
0uvmtBO3yndI3Zl18aXPe5NLGwSklWT+G64s5eR0ceWwReupdGNe8DOYeEryXwiC
`protect END_PROTECTED
