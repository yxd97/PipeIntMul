`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNsJbT3v4r9jF6T+k0mAtwDNrAZNEJ2BSAKMJ0kS0P3bPhS3wkXdrgCCuyHtdthk
/gNaX1BZV1cdr2lhRbm1gPCStSwASj4caCiFxWxDuaeXmOI2fES+etfYK/kghjHO
uI7EmeLryvERWaDy01A7eyjnhPu79Q/mMvZVRfP+Hb9IihvAJSyuAZ6p5G+6RpOf
QKKUhb+zQGuZ6y4E2iqfdRMh29EFgie8hN8yl02LOBD4+aYENMzxf1R4hd4bfd5V
w3bv5BrSWPdJo+cXwI32OpMSZxWxaZe+AOwnXQsZEL8BIbQT7Y4zfYrhSj7HSYLG
gVxB2mqNHvaFxpeszRHwdcvk7VP1Q28t58Wb6/7Bpv4sOVhlM3qSquHJyRvy20vx
mflFKjhax5v6vHGDdGFH8mAuhV+I0c4bg9B6MXuRytY=
`protect END_PROTECTED
