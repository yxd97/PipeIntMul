`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jmBoSznEYFJRSB+L/+QuevCBo6Sj/ap7V1d242RfwX+BM+BZK9Fjj9E+5yUBsEUc
kMyTE9vRXIVEsYVg0Qsk9Xm/oDU8W6OeA78aLzbnzP+yuLtoJ/ryJpFXkpJIU2Th
d0eKaKm7VukYlmaJuJf55T39Gy+lbojk99LqSA+JFpVB6QGxXQm+fbkFM/+LpzVx
N24+ckbzo7K+gSEQc2ivxrS2oIRnweOxu90PsVqCEIsGcJvuEp5eIoeJ0YfnAYml
hS0R91DOMY6IACaPrD27Egp+SGrUFfVH0K9VxqxDo1EMMt2ipXwycwmGRpKNyJ+H
tp6UQUwn7OOJr9AP44Ab6d7yDupyq1v2hb6AeepDABJ5BKdXdx34g5XIoiuJ+DcN
HTuIKifXEgvK4jx/cBumRYHsivcxjinbVTosZsaMJAvzUUXhPZxTz8ayxXgNYcQ3
5fXt6BZzaTh4dAw/aNsvSVh0UuaRcvmr5izAP8+FpTERktTZjxhQZpGlLSpTbO/h
bvBiw8bZlLblQiRaygBv3xl/pP7UUwV4HzclMWx7+71G/CYYwo9nprk0dNfmiLlV
hPFUpET9w0/NEBu/ir1XUfbg2HHzsn8wKguYlrWKxPXAHOxHMvvSYy+vi8keIreM
0UNMargU/OXVR7F7JjCytRAkqeSDbmm+4b7BpefbFid4/Lhy+eCH8W3FYxBPQtmL
u8/hGJigg3Gcl3HoxYVYdX2k//ToiSv1pofTIxDIcgJ9lFtnlzh7lWuCLlfkeL79
fu79H5erqQbscwOd3DaaI1QDE1n/E09T9QUUlG0I/q3HZOCvmWfnhTGTxQzBHxxG
e/OuHcjOthYrWXVy2XtioIz3eQnhgDnd2/UWL+TYbz++JyqrtXF8BHNzSjHUY5lh
SCzFDRj1yEyJHBE0bjbeg5iA8DMNFALvEGxxI7sbxKT3I/w1KpLikbKyWDVEyCZw
kmty+MRcjTn+nebuwTpCVYhJKayhkGf4gzE5TMmZhePnt51ES9amE0fwJ9yW5Tmz
gJ6GXP4Sxifp9x4Ot1n6RmDVt74rAul+P8jdJRlfvp5+Kt6nB8pl34/dbFbP2fDQ
1yjyab4xDN/NKdxEgdKk6Q==
`protect END_PROTECTED
