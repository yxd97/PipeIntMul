`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8RtedDjohk1rpl83GiYcL8RFqGtco3N77B16Y+2IRV+ktXxc9R95J58UAriRUpzX
ZQdba32+fdeDMVUHxLuSQI8yWtGZJmS+JolOZsirAVhImOJjdaAOssNv0fLxQeXL
tj0ttw/qGO5IsmCqXojt+emdzxAed9nhAKLXPsROsw/8iwoI+H6aWYzjEnet6jbQ
4iuxyUMHUxqQKwYQ0bFEcuXeZuegdgRl67vwMAl1mU1cE8eSUqa4/9eTYkqbHiuM
KTsZLTSc5QohokeQGs1w3HHymUmVNFj0AfMg+ID8InAUEnW/vDaakFNocBlAqPMn
fnyf2xh7OkUI/7m1wKTW4J5/kPjje4G90wcxTzR7igo2molo2B06UsPYKpxufpD9
RWqCE67AewpL29Y0QUCK1A==
`protect END_PROTECTED
