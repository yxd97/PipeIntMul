`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/fe6cdwq31RyCi38f7jai6rWKIFWbtHZSH6dGvu1pCxPaFzzrMLhUILfUaEqze0
TbXO4Q+opfWSb1b5qZw6aB4W1SwGrCDsmtvZLS0h6ujinJk+xsJYkfUnrwWoF8dJ
p9lOKR4XOqA143kFgI50QAkLu+ozcjj2RM6UF9gNlaP7p0KT8GWaUxu4ZeC/Krvh
jV+O0ZC4bjVxOyTHmbdHONpDKszWDQ2Gbxg8BGkgDRBWodTSWkm9nYXbwub9QdfA
4cRWsxi7EeLIOGNf1p+PBJLak3VARk9hbew+UV8bDT217O4RLkFusESD7z2Kk9Uf
tyKQJ5cGXJhr58oMMYPw0oV/HtRPGpL6NrZ+NhtY8M7xqIvUfHGWFQ77LPQWATwa
L5IoKWBLBACA2RD3Iw+FBtisDFJ2PjWSn7g0gBbW5qrWCKe/6r90Dkw3LNt0w+c1
`protect END_PROTECTED
