`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pilkHagLzU4hxdo1gmgdtHR1okmTs1dbMotNljyyvcFjeFe3j0b7ayb7ZB8LG6SA
fpnfqV6//fdJhvefxBvbkf6vshihB42Evs9m00UeYHaiLjodhRhMfEf+xOfwP//a
HY52OC5cgAO5DjyxjfcEd0HJNWIwNr8Grdq6pqD5t6mbP13vFKq7BkjNKOymBirJ
N/g4LVU5L/CohAAb+5Y+q14GGktoJrjLJrAPXwuMd/rX3odqXHO3PmPkiAKRSRlU
tDTzyi8w7B8hlQ20pZSTC1hh1bczXQcWsuIfosWdVo28h766JxxYxQbLlUlj58Ei
dj4KgY1btq5wVa+KUumBVA==
`protect END_PROTECTED
