`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CgwzcLzcPMjQBdtdHscT6zfjPtHgr7FpQhUl9eUATkRE3kDVlYbljT2dh92+KxP
Ds4fKzc2oD/C3puY0ZEXW7tnWtQFQbtG+6Qmv3FVZVAShVv4esVX8BfBwOJ9DNCT
bKWOwiyZS2uTjzylsOA6AzAcNj1e4ohYRaYbk+03f6xCLUav47Jxm/nYMruQM6lp
PRmYim+7q0Gj7x9ydNiLHwjU5UfLvu8A7AmJ8wiG1SpUTD7HWB3z6BBmYdVRwnp9
KFhegJRjAVEElmiU1XPe7F0PCoOxF6ym00plGgFhbLQrmthCjYRProCQ7TezgBXR
omuGqM1cJJRlvM3psOamQRRYCcOWodd42GBEUcymjLhH4u2j7DgKjWLkEUb8AxKp
GOxEMw0fQH3PaK/VkxGOsUBH8zd7bF935tHJBq3iQmhkjek9ud53va5MEmLvPGHM
/2acHzGIrTJhL7HjSaSF0vBIpsmGyg9ECTY9tLf4GSc=
`protect END_PROTECTED
