`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtqHf4xbhCiqkrrYLUYD/5RtuYM4XK+UgYfOM37eyUe3DJvf9iElNrlYsV1JHZQE
owgCJw2jTb6wxBUywUvdfbXTSaHwttCVE+LpW0dVTL1AbpbU2mb9nvsOmTDhBiyY
FfycIO39G+/Q6qMo2n7q7CAYueHcMVinaATYqSq9R0imBj1TMlkODgpO2ik8a/7H
GXgzWJihcaYdHQ8LbAXvtxr985vq+wnDzsQv5QvvaczMkTiCXe+zQdcm+A8+5mvu
NKVZp8meGsE76pXMyCwi44Yu+PdOMaLL1DKSGbQT2N+1DsplhjAS2x23rzjXlxbw
v3DbnKeRyJOEZITQamg53qgluqo5AcYG7aXrcJSTjezg8xt8bZSMzZidDbq1ZWZh
50RXZrOh+rUJ3PVnBqmNC0u04ceajEpnU4bmprbT71faWhBYip9hmAUa/fiShpjW
dHBh9hXQL1+NCIWICBlw4nonJ4Jxxl1yFWkP4dGxXdxuS9lkVl35fOwAskYRG4Vp
lHyI0Zk6TRsTMw15T2IQzftY5uBIZ/BXZ99vVJRLGdDj1IKdJUzpvSTKHxQtkqf9
8uI552uYBCj15JQWVzvOu6TtUfhubOzOl5q8HgBGK7HnGP0deMAh1OPkljoRlWhF
Ul3uluSIwz7C3b7+kcOWx6faGu2TL4sAtcp/Xw4XaDhYEO5PJMOWh+kdSpr6JuZn
KM3ch4XTPmFqPXTV3JKvZNqsvJSxbtMBMVJcuZuoDaPgbjLCtxuLuL+eu3raNPfT
i+lZ/jHb6PMF2fd+nwrNTz5CmgtZ8l7qwSGQyxnVO5WkW0sTtzm3A2gKNu7ItJGx
dWqxqsa2m4qUtAh44qDlCrdxWTauRwwSUU+qgwLeU7ZiGZqNFC9hAi07Dq0jV/dv
sMgkAOeHIOPw9BNi2cbJbCACjT2RJYPWSfFIshQqCJ2NFdmId8uwNuUL/1bMlsVz
wZw/yqv52P2pb5ylAFX+1xXFadhHSpxmf8Zsby7Wpq7JymVxfgxoe2G8bVrH9bV7
UCuDAoHJII0TM30rcR8IipmBbG20MujlaP4rnMkWIH9F36DOyKCxh3zikBaA5F4h
CWGqntesYXJFdMIB/Td6+4pyILKdhy28QD6yi7PjMQF6/hkLXvqtACMh7jJTx9V7
1JKdFDzIFerh9IFBoOSM/Dh+Z5VoQ5xsxsJ3SCuoFeK4agDFQa2JZzSLemPkA0Lr
ujE8Rao6VtZB5x0pbq28LVmxSrc54AEU7YDavRdvP3mNyvVpz8Kf01MhnTm0TIwU
5fTRAaS+AKPlA96ZHZW0D87qll5436tkXcSEETJ1MAo24YiG8ZpXi3JG55UIor8z
8XC2Cgwn08BNSHmnUNHGBa9u9QFiQ+FlWCd4CpdCTcwibZno+9Bvu+/jYSbFkRuA
5dLJ0qMkUHRJ0xmdgj4bDwq6dQlZeoXweipmQq91Wck7gKtoCqqphvBWJLiKkevH
uR7pmz32hfCqv++Earl5p+IC9XlsuKfKxkffia+hFJy6jMNYRa9bpitC8SDsUhhS
sIihBW5+Q7/8Kq1FzW+qtRuzplW9+AuoSctnkhDAiqqag0S/epLSZnuvouarnQ3p
M6knXoKBgNIGFCOGMj54T5v+sAYMwa1j8Epa7RH1NIV0eERF82VO0GYjFcClfaT0
Y5e0Hrt3EG2TXt/owXZ+9eznXHeZ5GFmdThgmvkQwL74hdIwGO0Zc9kVkX/BBaCI
kXP1navDArplI/nAow/IciEcQrwtZurGGVc4cyd01mu8PoDch9Itb9qSHImF0/iJ
raPZVFoqaQvO6/uxaxBwVzZv+SRIj4VGQRGDbrC1oT3CRoAerv8F12ygNyivdOR/
YAG3UOVg9XrRfPVJISpzWtcsksTomebNzQWhr995tvLmvQV9fvwdvcMRsYfVm6en
qJ3noMGqHQcyjfNzzJeX42aKdw8stW/74Te8c4/WsmSNEG+ImmP1FyWRjoeg/Nvt
mnD/40Bqf2cyXYiqmeJRYXKqyrxJ4L3K0vcIglUWEjPDOSyPq9eUqOnvrrVBdAaP
QgvunMghwX5i0ynhlD57R77mKF4eXUYET+STSqTOujO0Xn5GcsyZ/hoqIonLSzUS
RMBZWDjEfoehVG97ynQaZLAJehSX9IfkWnHPEwuKKuoiiC8kGAdHEbKqL+JRRQhJ
QTCmmHrDYJTiXAP6rLtaGjsX5RVkg7T+gDrYqftM7/qs9CDXt72gB8pUs8vOxa3g
KAzC5tnH17C2vo0O4XkNw5w5a5Pu7SJwqVux+8F1weS73INRSO9bAcj+ST2lLHsK
F1hSrFrkOap8U9dvmEA1HS/vD5ydrKL/CT2UzHGYDytAGLowZk9h1axKLvmlWex3
6HB0nao8e9d2iq9SwA3fza0Pwhea60j6tEea8kEA5+u0e5YhZqcc7v8EsH0qGlCP
PtJ0U2VCfYWIcjZfG6yydhsC5Cl4yb2zi8MqM3A4f7G6gqy0DZ5sq/UP12p/xO5g
b9umtfzuJL9PcakGmoVV76WGrUtoF98m4OKWVSG25tKh38s5+QtxwFhqfkqwoBdx
t57noPDUY4qf+Jh0tQGOPaTg/lNGa3SSP7ZlmXWpaLkavmvPL/qR1o5QSvZtqQ1w
LEyoHPJdwjVsDOGAPMNumMViiQiNs6RW7VP1ocBFQF9e+iT2W9nAVXwbrz1kfQWh
fLFcGR4NxokkfCv0N6epLIGEvBnV4H88uvoQoyCCFfGQiiQkaSLU8ZA5q5M4WACw
V83WOEeedErM101CigRwgYhgzUPN/77t+M0IfBK8gHCLt6Qa3ankh9BidyPvthun
X+jUpCF2ZLPl5HQItl3LLM9GzLWA3/Y6Ax3o/JpUD86jDMuwiAzFDDB+ac4F0k8i
1S54oBWkY0AMJTkzLJSNb6cMLpnzgKn+7A8hx3Y19akZABC6G9gRGfgFJaQRW2lp
tjbIujINNCeYa0/9inx9OBiwrZWKQFJfHLrKFcQ34QfJ4dg6NpJCVVLLWmpxlV6U
tWK0NuRlQXdGXRwMsrSh7GtI05cCRRgH4MfEAvuqbxija+VQXiCkNfD2bP+8QKrl
gfBYO6bCg6aubSt35GB/hy9aG0O1AFcUCSUb1Osaiadq7Q7h+Vg9mIj1/O9gytxd
swcqaouKfFKdAOxtHaWA8nEWj+PhnwOhxsn77rNUHFs6pRblrp9bHlEKFFjJtOkw
ZV/FgCbRYhdMouCkC2PGrQSpgtG7Psye1qQgB8LAAA0fuXVI9eLmO0xwFUen5kQh
yA1mW6uD2GO/EXSOPhs7kVAJ2WEWWzhtdGCA3yKc2BqaftwReOPOQ/8RAXupFqKv
lRwvTODNiYEUSJOIPK8D2ZlOmhB4tjym1WNnSUeX9qNAanOw7E3sNtUPQihnZpaQ
C+Xcw/aYESQteYPKQA1jRMx9bQmewB4lx9y5MxUnKTDUt3jbOziQhOcSj4zQMcbt
nICOtKpY3z68taaQl7/D/9Q0nsJ4zqiA9G2HoqudT0c7oVnto5BkpPgSzdb1UEAa
ZNsDM6lq4ByDWO8tv4PrRtwTSMdMgogvXG8ugJfJ5fjZYPWE7psytfmPiTXsabDg
d7pt8xOGc5w2Rf2eThTRCUZhDp2PY+ztVgJr8mbq9V/qKPFmyZYsit7o510e23x4
uq6GZKXOS2G4zm4hUvTtmWZ63voYtbRX6uBhkWPfraLuS4Y0Fmw9tCtU53xvMqtJ
tU6Z3P3CZJTwqyCg6mF240WIsONL4oebNHgi7S/zdkokxezlTEYOUwbZt4hbRC8m
skLjFCx3T+n9jOJX02nBWYT4/d74qmS593W8ZanWsJ3buFBzQfLrmbO3IT6Roqyc
lXy9XlxSsSNSUb5TrLI6WlCGRrFMPd2qrjLbr5BThsQmM3eLgH4hN/YKZYqKBXfP
bZRgv5hIF2MFZEdowoFvEnEazl+hdPomGPNpeFev9KNmY4PgvpZhkipvS+O+HrZi
GZOmHcyjfwDzBuhkkHpMJznu1qxDguXHJQbCPEe7NPwzL301y/vsCtrrVi2oeEEM
zu88YBl90OYnX9TyVS/xAm9jKwXRhEXggGHP9XT9JPah6nMkJ8ftEx1BpBBFHidx
jWM6KfHLzOnNjYPNq7b4aXZsh0fpR2CQUHiUJbUxxy46S9nOdLVw6t1vINJCumTR
eq5XV0ag6VRqG43YaQWV/6sjSlzLXT+FiToPXpHasw5U+mOn9MzKLNTU9WhvbziQ
qpzblE3wyz8XaFzzxNykLaeoDaeacw777M9yEAKTVUi1cEh8Zt7ZzI0MQbaCIfaK
6a8xoiooDYg1l//naaFtMBwaFa9NtZwo4APMXUZC+Tjag5biy7ZbmvQjR9+6HTq5
/ZlGs9pn8lMxcM7ArQiTR8KmGMOl0lSDnPYZQz6UkeEniNL1gx0nFe6sDHif4l7v
AH2CtuHVS1QdSM5J1KScKGqkRfYglwiUnPyoJN63p9oTAzKlLHporJ8KGrWr3RCP
Ik0JIggwOoppesXDUClVX7X4khtvgJQmmV/ZvrAgw1I=
`protect END_PROTECTED
