`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LCI9Zo+fk2mHbGZ5iiPAiM0UaObCTBWkMJ62yuwyZe5oHeX0V7i3DFfxcFpBfZxh
wmaH2QvZJlj7D5a7g+98nXdqHw9E3gkb5nkjeXTKUiiVn4QJ9XBF9okRpLM4ejlM
IfvpR68Y8ffI/TZbOGjV2s0z3yUHfNknRPSjCSvynJv0AfmN4/smm2sbA+l61F54
nQey3aO652WDj3HeMMEasA4UYFAxkdJbuT6ZfyZJ5/C2GU/9hsiR7DUVs9QSg87U
iiipXKGw0RGmSSlU4qFLm0ZXgbCH3J+JHEXdA+HDYJzvhnfDXgvwDby7jYZNmxjW
9wDWK3gThjJYpdqFPXmZ4w==
`protect END_PROTECTED
