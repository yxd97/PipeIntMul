`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgFrP+q1WHoliYAwQGPZoeaiDMgns4faN+pkTLebVuJ5opuUvseYZPZeUGHzQrtL
+D/HiZd9jGf8+uVLA5ZXychaB7EA/V0PcfWYlqYPN/TRJIXdaXhas5zbDglOBLUl
X1EC+Yg4EI9DTWennqk3hTx61SMKuHACgzeTrs46kPV+w5w0nh7E3RJ1tT/CzjtN
mlD9juqWmtt5s7mdQ51jx+vaOfVb/5YSEJcYlm5FvT1VamXnAZQR6JROE5DMQE3q
yphq1GIYenuwoQeUlXVY67BMxIrBLNHko+tojXIPLEFTI67T0kqbVSjuWXbv2BQf
bG6ygVZoUd3K1ITeFbe/dZVxFxnHJHfWABY64wvfxxxj91Q2d9fC7JJUzhEmVy54
`protect END_PROTECTED
