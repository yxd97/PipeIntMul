`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8oAhM0cBz6NsWolD6fhm3pP80+oyF3qDps6jXtZwC5wOirb0UL9OLLro9su4LUi3
NiR/0OJVx/p7IRiHQo9xYnZawP4FHkvZCdscyKx/IhcKfOHY0/oPA9L4aq8qZzJi
KH1tBGNnDH4FnMRWEILuxnHAFU9hB/h9hlXeOlpqEVAsCxuJx/9U2GQLHpjMzI26
F08KEHZtaaaKmDtSaFYqA2qOvgf7xnqTv5bUl9GEXf/7frfQ8h9dXreJI50GjDtW
GHqgGWjXYcHY08nNSUmW0qNrrJkvfjdfpxPUxmDDZ+95SsAAqlNvLFeTMK4PmOFX
qPvgTK0kjaGPluNt3/TCgD0eTs2G+xv5SkieyQap0XMj1nFKsoqhGt9DP0pQd2UH
jkS6XNOdwzr4YgBiRBHH8F0l4kouqgtesI6xssRvDXusm+2HRVSq/QsrKI+7FZRy
`protect END_PROTECTED
