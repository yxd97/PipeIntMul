`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9olQI1FObH29acWS6J7wB/rsuIRPz760EFxUKq2qTr4JsnIvcpYBwpexQQqEWxue
qFd/j7ZNeZoZ3IXynopqv+Q9Aa5qLKO2L0uNfenZwEEh63BT5ecKrGRf0C/WZxYF
NCKdstvJUZa8ay6Wnkw4IQHPzbWluiNeIZMmrFyKHqex+gUoaKDLoxdKrk/GLAnR
0J/922P9DFO1wlTZYSreNEIHCXLpTYAoRqGcQtTuOkdLZ+NfPahpz7X0Ui2qpjJF
9jpmhkogrKdPIbcDrwsn+Zqgag0tnrTcieFKikxz9IZ+HhPicyMtMgV8d+aNr81j
L6BjUINKNT76PfQ6oAUhBTd3E69VSPSvPZW10Jc5An0rBaG/RDgH1pBSDQQhvAE7
RBaNJFK8x5/ASxgVEUqfzIs0WrvGDUDQbS+q4stF5EaukIc1EfPp1bt1TMGgEGw9
aOOJ32yteS+VCk6qRjezwjF9CDUmt+bsxVEGNHy2vod1rm4NdDysz9bpwjhYBcP9
wkPVU7NuKGEy4peIwPYS8VScKk9rRgkTpv34gmM5FoXfRyvT4T/g0Gi6hxjkKp50
00GEeMeq8YcGBPeQ2v7IjaKpP0MLMMM3gVI4wD6Kmt2k0NKjsi0GzlLp7zanBiw0
xO7Cs7jPtv9/unoH/DeDnRx3eAPkgVOzpAKVEWUuGhHOIo5OCqdvzzkvZY38+bfD
t1t96T6XpfETd/S0CMKewgLrHLu3nkBNYnZNsjrdBsmNExE6drnv/fE3/zm8LnNi
rIrquLia+yMXCmeApBzBMz//zuTcils5q6w9vs3gAjbqA+3VDNBVaxuXwNOTSk7A
m++CAlsf2Mc4g4tKjXnfrzUWNB3AQU6oszEPpEqaD4KPhNKw8c4FwnwqHyqklPzF
SkFa1ZN43qPF8taY/P4l6zxcIMM53B8xAGsTEx9tqLvuj+MDf+Y+r7pRF/k/Kz+M
N1ul9gDWgdYqtUN0+wXK5rrT4v/ALldRxv5NLT0+FVfdPGxX+19Kbk4gmRbZ/FFd
iwNpsezPsepGhEy5WTikbX3V+T92dRNkIiNu26lmYatta7H3/cWctUFqJmwZHYK2
ahDIqAP4KANjFFkI1RkWZQoV4xlUvGCyf40yJkSYxRtJDFVJhv7HxK32LAmEeP0I
2WkoLdeOvpKrOBl8gC4OxnEq6mWVGAGl0TDYx6A2zVFmbmwo72Nh/fMdPPyyI/JD
M8HxyBwM6PxQtDSsuBkeII8HJWad8ai7uXVUztSUw1GUfcmtoWUqVdIMV9ajnQPQ
rVwLj3ZXbn65HvBuCN2nOX7sq6sKsFcCWxuH2M+0NQjbBrHUgouOEMu6SbrKnWbH
anNFyUUZwaXaDCrIdCpJpQTE4yilYu5D7LHI6UyGoykrksXEaMh0Npdnt6LhrTY8
05Gco1qjy23fg480DODR4Sw5b1E22C4Kf6r1Dvp7FcZ1G1QEIKWm0DWoseqxlSA4
2d6e+5s4LD6UP0VQCG0ISzvsT2eimOCN/KMLqex64u+4gxMeeQIu3R1wo/4byuyY
cVZ9Bet4zQWOkSrvp/pcGh+yQCfNTIPgCiQBN3Z3b9nYfmFT40+HTikbCvoSNUsS
rlMNXZBSpWQQ7YrA1neWczXrtx0pv+B25JmcA8wBfSTMgaoE8wxcNGkO+koaJm64
1WJ20vxvBbLq2NvyL2HM8dUXBhzz5gItInBlfXHUwcZWIM1KhfdmrYfShOGTf7dL
supTOL7mByTAEA/CdNs+SgbODRr2ZsJ6fBrSbsYHNabHTdz7LhUSje0s2JuEgIVn
j4vyLGIOV7jziPJkLVHJfbVssbtQ53EK45aX4NVRlBrLlwvBVOHFuz7I2LeHqjeX
5w6CNvPCD8AzVHEwJADHdaUB3MSR+StgSvrqDpew+ycO1Rm59gwEWdaSvevgUiTG
i96Lt18D20XCo+/YXOKYmEBFQmAvIEFx6HXdJE6Wn5WOPY9LVpaTc3zQjJ1INAv4
rn9AALz25b/j8T80Y4SMLfMXPrltX3ogrVVXLQCzD6J/yRJV9b4z3kma0pQQOETu
rUJeR5RRRKN1vKpA0wpc6q5yD02Ez8AZTrS0zVuicMpVvD5s6oemEs8rHgfcdhgm
8m/8Zp25vv19DnloYR/awBAnzd+2l/Hkm4BXKiV2Zc4kJo9qkq8Sv/u6jnQ1E0IG
k0I15GtVI3j9qVq/0gs/qW8dLiioQA3jSTetfLVUbYpexsFOn2esZqKMUibce3o8
nzzexxBnXT4vAUisjelpUSFY6JwH76ZYPSxhey2CtLmJ3siTWm3pepNVmsDboKeL
EekuBV67q8Emwd8FUJf+4tUKCTZSYCXI6Dl9twyPFudByUxTTaOz+waYkb1mTjq0
CLf+OacdlYiSI7Sq4Pu8Wbm1F1zqlebM0x7hXNXEkxzIiGQrMzc7CvrGGbrMqyWB
1gI+yKvYwxBqf1dA0iyuPdPyvHApI8YwH0UjcV3SeaRXzI7oe4PJX7r3ma3Sw01M
8MVXGAIfwWPb1s9oZAzsmjbsoKdIAuP700PI3sUMiQfsvxbbIYbqSlMbF3kQVUzx
/8oYogaKudBj70NH7O+ir7zwSvOxaS5Adrfb2BXpCDTOFxZn+I1wO3CKXUYRe1zC
2/ewY7m3siFXC/IygalXPI1K+2JRpS9qTyUu5p8a6wv7OX6Li9u0BOtUV96+EpuC
TmfhDsFbIexyIP9RSow+eJMEuCKHkN3vwhavv8NpBHmDdJURit9gyJbwQSJ3dPXM
+/kmQyMMEg1UzOlU1bnI1rV0nswylE9rKkGGA5bPgoQ7rg4rUJ7eJNnBQgUaBlu+
yC22gsVD2hQ0lgRxCd16EwJiiyOOkyjo29XiSnAXIF90EF/LDSu7I9wfN4fiiXoa
u6uEfQIDEEjVvtx52153zXegWTXiJuZGX5YZWpB9iwNnfAkeuPtPpmt3iyNSSXXA
IDBx7QjQw+XdIaoFQBrjuNFF76ICN9OewtxK0IHJvPqvkarMfXA632lu1teVxCzR
mc0k0qdWQlunDH9UtuGw3WwbjqdEFxNHAdgwXZ8Xm1CD174hzmAZeORFxPxGlrUz
9waMCmJe+k6EWz62h9I8Obyo/kmP5xf2eQZ85JCbQRxPCx0fXFH2LvS7mdMWdD0N
aCaN2hScMtnNUixcbSNz3JHXUCI7cB5N8LljZmdEA0RWAA9v/jM4C84e9d8wjhtY
9VT/gIbsaxdLYeQgtW65Tdc0AsOvMWD4c+/1Z2NbBqMCF0FX8lGdoUdHp+QbdmQf
bPkh81SzdU6DnWsbacZSsmRHojhDNXzn6KFrlewJUOSMPL09UsIDmtOss/xtPp2N
mS4mW5UmHBTEdMYgx0KOQklYsFOIcW+sV+H/BF/I1C7HBv3ocVQxSpQfGgQHcMn9
4l9yO9bVpmrJS+CqojumXSOVOroFAtEPxKMe9tqpbLV8+zpjS78RgwShViJjdx7W
BWse3devbAyV7pe3G0vXEn3boD7tv9NqZHp4ueIAo5eUU4f9LGRSa/PR511a09Ay
alwV1WjhtuVtlNLtxxakS+uI78kh7Vb9/iw5ZdmmZyh80CEnkOUmwsOap7tlTaOG
dc9zvVJxBrhH+5c5ctKOHJdsajliEUWZ7/P2vZf7tX6kkoG+wg/v5l6J0S2sX6TA
Elu0zqGJgMzDUBk2oSv2X8hN2MS1Tbwkvak/VM8P3xJHF4E1n2nbMcH8qeGXqVAr
BEOrDj/kNdhuFFxGuzTyLUGnmywX7ByQGwqNCFPmG0DWkUf0WhJCC7m5mIQQUzvb
5zxCu4c3WU3K/Pjp6nlxrljNtKmU+opDM/wxova6i+Bgg6HmPHqMM6RkpjmbJUSw
hctKWqBqOlsiiy5D8Q0amc4tuIbLkz7f3Sj6AfxQkg4F3MDdbYPOjhjIcKPfFiLm
cQB6dmFo5CuEmLJ/uf609kU4Q37NzedK4AZpoCbA1gTy7Cd1OfuN1RF5MbpmuxRB
e45MI8Y3zRAlOtetGGChWafYnE3TA5lpekkGWy1d7bfji8j+xWpUtpeBcpMoYdg1
dRyvf9bcXfq7KE8u+OLTXQZoEq9TbAyZQK/MOaeuNug4NfNMuIwoYycTfhxtk/+b
A7Tsqji+/Oouaw88eahE5u7IEGmk1ULjMo70we5xWNKEBW5kQELa6MWvrpSk9YOm
TzkvYOwc2y8BB1OLt1L89hz5EC+dJBDX3ORIK/P1wgdwqRYmQilL36wI3Xypwyk/
Fd1Zxq9WW6uKAfj/x4cVLAv4tVzWxvOKVnT+JO9BNYEOW6zCSWmd4splwkgDcMbJ
GKjGcWDVMj8p834kIDI29KA0+nS22kuR30V0wq1JRjOtCCEyPCe4ngCknENu/vIM
T3VpcO1XcR3LSAtbCmGkY+bIT/zZWrVzOa7bQJH6VUyJ3sf6AkAoEkyPZkOsLeWO
MSxgHIkXiQhm1dzLO2v9P+GvZuiiDgDRwEbrWkGGG1fGSZ2CDQnMaLqhHhCm4X0+
+QXbgczjtN94OlffvznyBYoiTYB+Q5W+grZjOds16dztKqQofjv+emehPI2ON8RR
ipsZ/FrTUtiEWFqztFFP/6MLIsS1gSsuL6M/MiuMJOlzfXQGW0XGlqN1pR+AjpkT
5gvXmebU6N1f8mhQznm9n+X5AzLXSi6TbLL2PBnagYd3Hg4Izaa9wPG4cqxvm/Fv
drRM+A3Ud+WFnlNxsCKcFCtdo1RVq8fxqtrJrOQr/6jKD3AxBVTqbel4Trcv8Hdp
11y/L05yrqwDu+ZtGbKI4o7wwTjreE6S6F61lDZZz2z5+1Hhrb/M+QTTiEOw6bHD
zFg1E4nLyp1LmWkXulvHOlRQKJ7CjYdZt+Y0igIm2TwoqODut/Q82BnI5sZgGVCH
nol/VlKjI3PfGUcFqPwtwrJdMFDhjTDaEtUozcLB6eoK/5KDmGco92uiX6Ku96Ic
qxemVTqf4p1ZiIVSH+2PhGjUt5a97jz+m2gr2ybJH2XymTC8DJh7McUo8zfsi0ys
OkMKXS7ifsm3t61QDBNU3ItYV0fbrP6ef/Gp+jpr0dezdesnQQUNL3MHuLh5Gc8d
O9OPQm6deLQfTOZtB8rrtvFMVEd/5A0o75DeXs12xa3FJgy8SbQ9gNG36msUgymz
45tvGjlrKOXi4XXHnUNdHeJ7fzC1T1AMRPl4ugxMIkR1wh6ED5rYU4wXeAvf3s41
IiY6C71bpSK/FcoB+e1gn8zMDSrHG8lnyBjmchRrDebFy9To01Yg9je3AZkLInYZ
MbgZ187nbrALYRXtXluPITHVMPImO9+FmABxkWPe2MziPX/o5935n/6cXqHM52Gj
xZuSLcFTgvBbloP5Eiukwwby/KV06dq6tcDnbAE9fGmNtOn4nzFiL0qNlOrWomsR
7PoFh1Dc6aLSiyoxoKgnkNN9oJuST+419xwCAygpmVr0o6bZkwuSQRKp/BJtOsSc
OjRncB8QVcp3j+ZnlDkCyojbEW0JvQhFuN0Qx1xPKDtnGKGxpTeqBPRY7mG3m2lv
0hLN8bqivVrUR0d1JYTIvjptzpKYrsmoGlP89571pXgcrNS1jg1a7/eceo8YdcBG
sAQZB7KT0iTmGnC7MC1YocCgFNlKOt7oSVVIPB/wJJmhNd/2jdUP+xnFYJ7pinAz
W5C9AATnnhl+Z1c2B4j+0LRN8/l5IyZ1UaCPuW+bgM7WxTmsMAhE/hHLosiLu118
AMJ7eaKWRO9m/9Cz8yRINpS3YvOpmeJVeEdtW1/hlYzT7gdXaa/31iNQR8ppBAlo
+a3wYFIPRZc308AcQ8j4aGkWS9sk0ROxR8xNhi3NTs5cchX0djibfUOS1co3fbUQ
sl4e0tTdtwdc/9UZpzQmEzhTu6bOACE3Ca6Mb/mfYueRb8od5AekI3CWe+XiKoy6
KhrmeVYgIIinCM/TEcwv5LVCrWK+xZgqheTFG2I48rhGIDdUP6uUSuJL/+QIWmtB
Ynh32rQUbLkgwWpx3h/TmE/K6v0PY4axx2NCCUpys5qMY4D7vB+JE3KYpQ9eqK2S
Q7/xwK5Juq/Njm37L/TCXSx6/6DbYhufNY++er3CKIkWjBTl3tapzaGUIvuz/t1y
9qqpwCLOFzFFki8jKJkxdEW47RmUXbKJZeakaSOetz3wE+jSXXF+Nc+CbAmvwLjF
joelKd962cAhrn9v014M33aInLeyUsDIKEgN4gVfFRi4exBYL1dj0LYOwFRubaoK
DFgT8oi41yoitJfCs7WzpVAHNDp4uHTeospJEwji4834nui1Wg0J1XcYBg1U3yzg
ZLg3AqhbivoUUwQBTIuICIfAYK0vzt8KTQ2AfwOiXkTlL3RT9rcl+ZcxofCB6SqP
/xtSOH6C99X1fIWDMMpazVmGDoiOxfsgO2mel9Li1senajhBLv1FEvMwQColqYc1
gWX+S9lvQ431gFon10j5DvPU4YbSgWDIRcHr2/EeD3V3a55Q+kN6qYIONsHiPTu3
tZ9A5v1/HFh/EzsFrhghc+QqMx39c5U3UgyWPpVu1Lqe2Sn5k8WgjElutBi1HFRi
HtzxxsaSMsSfWPJ2uFt0285B3tgUD+XgzbYK0FanAMxi+P5dcVl8MyU2e1Aau71u
2+SAc8UvtclQpPL6uHNqt80gUcGOwsDirwW1Xm/x8yoBrUodhMi6aKko/vTMufqo
JrpNY1LJpsOwph7yyLcBd3v2H/c2m/3zLuaUx16kGtFpN8asq7cjMgQfv27wSCfO
SfNhuQy3+qleMOnvJEIbB2fzggA4XhxXFMoVBFquZCCus57pm1AZYdfFdAoXnn0f
OLvrunjS0qsrD4Oiw7nmaYT/Ft5v4wPO3+HN3kIZjRSNVuJoStjpGVP59Sm28puO
VmJlSGlScO2zGO7tw0I7EMPP7pOzTq37W50WIBrVk+qzS8A3/yB3D/J09OSX8+Yp
5y0UT5jw+6IxONf/HD0fUzxTHFHTjN1dIu2ZeKC6u3oFPuM68vbljDeEPvFqkZt3
eqwnNwvgZBRTyvGhuVLvRhPjUM+Dl0XVVdNf3pwJGyB3jR7zUDHM6z0FDNkgDIAP
Bs2In2VcNffG/4AGIFwcQQRVDkoqZDVgDygmG+rfn2QFzCgoEXu54vXHbEYVM17x
KeMLOcH+Zk7YcJEipcGClTSWr4UceaItOBZZnZqMgDansUKk/Cl3Qsf9nz7AWD7D
mkyxLZlaC4ZUj1CilH0esYhUOXCfYpSQLqz/BKl1Q/hgbrNqMgPTkvScUcj0vDMh
yJfAocvMqLC6+1pCFI1nI8KFnZuOBWbkToN26E7HTe7klOiIIZdOvJ7rXDxEnDWq
zMbJnSdkKM56NXo8zNHn6iWg5auEi9FBVlatC7NxW4C5OCaS1Qypg4ltWI/f6pSA
pqrBnKu8p6HfBCiymKtMUXECOYR4gX7RkZYv2O249ycMo9r7IM47x7yf3PQmec9g
DWrH9JAXLknzeqLhujcoaZ5oXqvXjJlEuiyXFY7QKtHKxzTJWqb6hwzktwfprczH
PSMWJ/GTP3hJtOr18Jes1WzaNd4snjjn+FAmaPQF94Nljwgtg4xjXaVteSQe6P9a
uci2VrFhv1zHBj53v9gLs7kJcOjDyA+MGtvuUxYl6PetJMmCQoFYptvZ6sJ34eSV
NimoyBKsAagvsjDQ33ZmBJ9ECPnaasnc4hz2JuYke3cCqrhBBV9IvSuKA2ISUEbc
+x/joRjGaGhyzcSDj98AqCHuG+mqdwurgK3p4VQvUkZINU6NwRy7Hu5f1S4Csu6V
Wx1+urM9S3Y67FAT7mvHrU16BKuG1XDc0HoAkNJqXN4CwpLdMZxKfUeV0Quw1aWx
7ZoOLqcjTd7dJpJ/L38lC0rWSBuw9t++99TxAzTPS0c=
`protect END_PROTECTED
