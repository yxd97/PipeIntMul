`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/UxYTe8vT9dJ5zzdleCSk/pXGGbcXbvLN6rzlatx/CUlazkbqSyjRNDohaYl0Gn
C1a3ezE8w37dyHsVnnOixfbtDBhb/4jgZTRz1ba75a4on74XVAc35WNd9W7+Bmne
qug0wQeI3YR3SylDanene6Kxcgh0CkPcxrYCFqcN8GWfximR/YvotPdGUGh+KbWI
x+3kv3h2HWiPJKHhEYyD7FFbjU8p/9Xa5WabzEAIRobXZ1NPDL0M0XWJvA9wlMai
0yIKa1Uf0UFVdK9P36myanxZT2t3Q49PsZj/0vlVj1hofe4Bf5sm8j3+1ymuae2A
eUVfZjiFjMzyGj21WmgyeOVq3YtBe0vI2C/k4kHTnNVFHsu6t2elaEmccCxHTw0s
e/K2bzAA9WymGNgzyUXId/++ilSyUrk2YpcCbDtmy9wEyqd14pSb9p3aPY2LLLvP
Tk8zky92kcuqAAca1BoVvLjuX8mmKCMDKOJdGq33mboS1nL46z2Li1jqEiMKf1Ek
SLBBeXNd6/fVeWnSA2oDJNrNYF5/dK3L25oUrr95mAeQ/KmOQH9RjAw0m+OxWKJ9
DGUc6DXxyWwyYuozYxLyxZ5xqtATK/r5pEFHcIgl00MyYgQmjjYWAT7QeouiLu5p
gBHNaBqFbzXpEtsPrvcFQDLdo2IStDiswsV5YqSENusXKxJTWad339QXyxlvMSpv
A21YF6LwJugu0l64dWqtA0OzovSAJjrj21RBJsujU1Xl6SvIi5JQeMrxTDR8XjLi
Y3tLNIBNaMuDx94g2DUFXO32zgcFCI4FoQXwSetMbYMPSREPEQ46BggoA13EpDLc
p9L4hn7urK+qQWOOG8Rs5g==
`protect END_PROTECTED
