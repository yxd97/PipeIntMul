`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AMI/cXjrhHwszaq7wbHzizjdc09kIX1dZmof5kr6/MPqTdh18y+lrvEHo01Xa8tZ
WHpQt79AYRCrlILdqWmsldCCvY91co+2ueaJmd3LS126riCpF392oZsfas5Jzr9D
AcY7TmP0L1JEfoqM26J21eENmlYh96mm7iDjk6EPdCFcq+7uDj/B67OtXTqw8Wp4
h582PrT6mp16YDyj9w4iuOOV6ywzQPMZHSXvyi6vcwZuJCPITJNr3XPCFb92EVCJ
a8qUtctm/vW0kP5yoqjC4tf9LqW8Du4MMeyvWIuxOsj0dtVA16VMkJ7cjq8KUAYn
oZbTUB2qCJnYHJEvCVPIWXdUoKV6BS7NJQQVQZ1dER38fChbDky2VkmGJMer1C8z
i/nWYkSzxn7T536u/ZkrdSRyeaJpFFCLI58+b15b6qabR/PBT9fcSYhHZCPoC7eB
p6RLvoOcg78t6LxmqDESOMRPHP0JS+Cr7WqFS/jkDuh8KjwZ5kFef7UtD9pUcW7z
ap9nT0bsG3BlTzC0VfdwVMVuXUauhn9iTW1qwfsLRAvldphCTNns2VhbeHZuejZk
J2RAB6gLB1vAvR2YwqwMZDR7mocEtC8Jmf1MOTltvtuG4JxF9yJAF4joZU1dCn5S
U6CMqhisGVa17vSWrYQBUba44xGHmOlmZTxWCeMdcv12yYdS+dApxLx7k5GvNMpu
Hd0K9tSaGWzfbfTKaiVTaXyGQNXCiJhYJ+kc1M5IOCGPRfm3eTESrz9+q9rNxibG
OFbVgXp0L1I5pO9xzTptQuYZno9ZtBAgcoMR29b0LjTmKZwlKqJDCwtphoCcpnty
Gkvn8B+fSwsr0/5IhO4UcZyu9y3NI8rQCMHWkn90Wu1ZCm8tAyss0+Mq5DKV/smT
Hp9ZtsUbAtxDbFxWcfEsq5yMAAP0w9D/WHWbIhqi0ds=
`protect END_PROTECTED
