`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63ZFLG7Gj4/lWJfX9P8DuJeWbGXDHKKdt7DCJLXUAM/CgoWZE0dG6t0Lsg+QVELE
jEteHpwuJwk2OGMAtcSJH+phWiOcaFm1gQse6FdzEVv4MhpQBxAq//N0CSQ1+cOa
4TgSOKRYn+4klplDX8PJG+zjK4V44T6tQcCAYHX1auToJ+4jE+NHq7/RR7K442c+
Ge7x95xOwaedqmoMHLpm+k/smPcnoXirndyuJ/DDjOfDlly5sSCfdsZLn56QmSbv
vweMb8vC0BgUzYJQmhIohpeNE9A5/CfbSGcnR3NOLHH4cAi1aaX/2b3LXbjKvgny
hZPeLTw53o7jv6lr00JRyPnWrzLBM7DdDKCFpLxcs2K5E6C4zepu1eSfG3pgl+ss
rlBc0i8NDPu6RafnvHPyyA9cLYAc8Ed4ZK1hj7rCaztsV+byj5MjpclNx/5D2mwp
EIMmuyprtRzqMQWBOMBx2PEXCL5VaVwrSR5VnozHBzmKG/DfpVRE+yaodhmqaZgl
FjXpXZll+8dmqDxK7YAdnEPWRlzo4YrYq2TAsGyip7ijWDchsHKTdNuWnNb5xIRU
ylfOgYecgQBxaj/I6W3nDzDbUiSxgetUw/16BbE+KYuBbprgb1oQLFdRyQxm2O5w
s8twXNd/hCaySg5fIncQWnoF9l7TrDsKjjxlHWbghIyvN4L+b42wDoEUxxTDi3M/
2m5sE+gH+f31vzCgoiQyaoi+MdjkJghh81rlYELEBc2JS91SqeaEOzxOrQdGOoeJ
8pA7RXovyeLLb8PI8R1gi/WEKfq/XR29rog8XeuYYthHb+sVOGcwTrQG2/WSoyGj
tXnC7nSYNC0APFEI2L8ivr2M4pxgY57+ryY7rOFkJjHwi4QjJDwCD0u1YjQM7jZt
YGn7g7pjaDWQ+7qvroEMhvVydM8CLX5jvEJaAx8z9OXYkSSyeKpAe727QR4fGx3U
ycqxMLFmdN5fcSvPVhf9PnL/u5kYe2ER+9Cn+gmun0Q7p1mmO3oMHwWn8kn8Tfhz
NE1U5BL5iK2dx12f4DUBgAjXmPFAI0zJ5OBLIg9yxM7JZD6rvDLjoOPATM3doSkQ
44BbcTW8WC5ftMyjrz+3VGWsmxgbJeFcB2SYr+RoSVbSREwQkA50DvQ60z+ZzUlw
VNzXZYIi7YPlGDDluevHjEASsqgMdehP9IjJj7upYA0AnJyABEFbTqUAJgTIMA4a
7fcbCqV4vA2bb5a/vEkuzDy9Ern4aJjkm5rcP7ixArwLB5/bkBbdpM95mR0ZVK9Y
9za1bh2rCgKIFAHJJPJYnmhaexFhftv/60RskLXXBQSUJn79c7WTVSMhZ4usUfgg
QZEeBtvW0BswjtXyu4nHwnzSwirVYY7SzcWLLtChe6e7T0kMtXLMSFDt8Gbllyro
Iy0CMNyn2SM2MiN5zeQaBkrLc5t67Ns0SZWCddoZq4qG+e1egIFarxWvY90G9wqW
yZBJa9p9ba/xLbqunikys361/tMZMUysYFrDCxzmcebO6Q7Gn8sxLWY541wP1vJo
PiijRr+8fbcwWI7qA3vTfy+1SASaaPrEOFCO9JQGmVk7RVz9iFXWJvtK1SyqozZO
C0UCfEczS40lsLpbyqgGUXxX4gIV8kxF7aJ4vLiHZisjXZ3u+MwLcvCqz4+uK+DJ
YmYef0VKVRHL0LBi8pK8pyzHtki7r24YloZu4SoS9VJWZoYkBsKxH3l85O0+BlF8
xr42BIma0Xnal3Cp8PR3uHaufgSOP8mv4vsMKmBtgILkt+c2B0G4Y+fVssfivWUS
oif/mh6b3b0zYbPIuNE5zZETW2252hCvWfD0VqsobfOLdEd9hzT888KZwkIIliKp
7hAugdtclIC76rNxf9CBWJoVpFh7HHMnm/AaSWSExQa9PYgDPyAxgUkpwXX2sFPb
oyh6o+uBHNWsJReqZ+OwxPLl/u8W9zEkkyF60zblBJ8AcySbAZ40RNrJyY6WEjnL
HcUjabPVZ0LDQBQ/axl8dAmIce8TTdfGxlBvEyBmFk+l4RiXaPfH8RNE3Z4OgBsM
FxgHeyxDfm8LB4viWG6vGgVo0Wi6uJnI7skvYga/UjUXN7Deor3bm91/dZxmxJUm
qBSqFMM5QZg5utpqNxmgyDmobO5/PAL0pv4ZOcscFG/jnhR/xjLGpyU5wHi4ytlv
n1rOR1CgTeqRAOE+GJOfZL/Py4ifIIia/D5ILPCjD7X6YQK9JI+OTmQ5NieMBfn8
KPAw0iu93GM5Z148qdC0S419MWGQ8TfMpqIxp4Yb6Gd7wHr/OunRobbEcCvm8kMP
r3rj8L7GJej5ZIeGLTB9rz2oPMmeZwYp5ruZuzB7yZbmDO4+d06FfSl30y6em8gr
gL+Zxxzl8bFKoWBGpw9Hzl4KOPJwyn3KZHn9pKhdf53qJmGC5eLZocfTOebTa8z9
37riqn+FKdtxsDuvp7G4PdUeZOCtutlE/SGNrAAeSFSI6dQdtNeGhfUqbGjYfvKs
OR//fNu1vsspW/saR/bIlU+y+oz4uS298qlqHU6TYWXWWdPYxP3zChfPwTDK1LUX
2BDYgU1gaO77WFQLwHc4kDGa7UCwNLWHdoOq2+2+ZOeqbpai43DENjSc5Tp7BG94
q1fBcLFYPLaL/iAf+SG/y77KxVHucIuo7UvtL0Axb/wMbfmjXv7a4ayfSIlcX2Vc
/8tv+pheXfMDfssyBqC6rloAL7ibE1zPWdoOfvyYbVRKiQxQhJSJ/9qp9aKiMo1T
8lFi7feOJJr+3eTR1WKlNyccZIJqYkA9MVawSXXQ3MLwmikD0NeifmPZlCaukzJU
mUq25g63bCgLr/YMBZLJpQ6E6BwD3PvFLAkkYruip5EDDCJjHlJ82wlERlwz9gXf
uTFvjZpfNn3q8bx1ygmZbfweok/9yeMoYi5oGl7S6GBHTh7KVx4s1Kv1Mw2vHF/y
/lzcOGZFuPcSCf29xRQO+i3kERxv+djxPaMXitDrT9Ug+V2c5qtZnf8YOpqQ4TKw
+gXgd43CJaponxQyQuwudshcPXNiHxtCg0uacq/EwZsuqD+Xi/2Jtmy8COzFPgCx
QhI83e9hKshr5TWi7v9s4jSWErkE6l4erVV3RtysNUSv5Z6xRUEXjc8UAOiOOZIq
Sb9+xsFn7tEVET9f0frtWkCICD2Cw3jD/L1cnGGc7oJXkRpV0y5Mubo8IXF1g8Uf
dd4Rb2MosbcjHupagIKGaMoIQo0Ctc0nGrlP1w4VgMumV+Vb39e3aQnR31oP15wt
EFmPeIc9DC7I5dJaWQyM/krAdtomBpdZBNbbh1S1kmY=
`protect END_PROTECTED
