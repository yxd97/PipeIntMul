`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhjCAf+7jGKR45wnRBy+oUdC4cA5zGQ7/pm8hIYaIFLC2e4KqL23FO/W107OUfX3
8cXRNPL5L9dZAcDeESWQjF7+kiqyz1pCpmEPmgJVCH3wY6KMxMsc6RBle4U9dt1e
UUBrTVn3TWHToiDcvIrzhVUiDb9sRVRe0Kd9aAPWQdMj3cLQdALMqORHkFbpyk0c
/MnZrzGgZj7csU/uexsI5r/l3a0H1AZMwC26M3b0ZLGmOwteWh02DO1PBoK6X5jk
DNmnAcT5YklI2hdWASR8tGQRA0zY8rd0lwkO1W+9BEM=
`protect END_PROTECTED
