`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7s3V8NnW41HgUy7kqEFjNmfzGMorNum1MnnNJHrGb+pePB2BmowBwAKt6w21bWsI
FQHvGAYl/rUK6V1NNeJ4LKXOFa9v9VJRgXXqZILD3gPD+2QY14rnSTr0xdWq3Mf0
z1fAY+yKWvta+qkDuk49uTILmrdiEOiV0ioW2jGTfOL9c4E6mspboMYFGoCt1aZg
RF2T9mQ3pEmAw5NhMOejStU8hqeSsXnw5GRG0di+LgylCQLZwpMt7sxuqQy5GQJV
0hOvk0CHs0QesSDYqw/37thPGicf10ert5QOvpbyMhFZzKfPVXFiwDG134cBl+iz
rJbBpY6fRDaOVuHHxa2IQM2N+W9AU43QWdYDf19JUMDcRmvleKf/+T6iXMXXTFA6
i9+8GXmQ0NdXp2lvjRitZA==
`protect END_PROTECTED
