`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Cp2MIN4tGcTlWZ5tj/UW++0u17xbxc/ShBNOXNtwfhsSkmtKGm7hMZv8HAk22+l
oG3SjCuIRmlzmO/xfb9Q/J+aEGz+40gQy0BpYJxgawV6n6E/oiAhU7DERbOT9Zhc
y6+0G6AVmbZKAZhx6Cd4LFjryvUdGK3ZUpcUKhR6DlvXNiWPSbHXeCsVrjvcbFMQ
u8sZ4ljZq8/5f652CgA6cB2p6EwOC6tdENCuCzvBOGNrmI/yxZZ1b4ckb2hgLSJ+
kMPQ1b/VX4jTgyHNSa9zErATUH8KDtr7XS8ZqLWVbenPhiWSqNCjKwrA7iOToDoT
gdLGLg9eMNEQd4F8AHMUpg==
`protect END_PROTECTED
