`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4G0oaxrevvmEKLMVKt/Co02/j/FqFabKLiQ8KrKv1cS3IWuzkX15qiRigtXJV6YL
aEepgCjjsmQX7pg/2cADc36EY4rSJ0NgI23FVRwlhk3c0+5ghraJBe7tfYqzRFcA
GoumlaNYnkypdJMrHoEwM7jfXJBFK4pN9V4YE0HD7wmixQPbAN89xlAU22xDJb4/
pWsB6Xg9sMG7hLuUNwAUbpPsI+ekQHHLMgaqccikJ4f1yC/rbFUOTHol+1K8GQGP
tBLHC/vOTbribmZrTmkh7sDLGGAhT/mw6JEuv/WJdWsP0wZqn5p0oFXnJ2N3hIqL
KpusBjdOparaQWGPedpLYq/VyHerJqi7joqH4ImLBTK3qgQnXEh4eUhC6c/RrLd9
KDnwccbAhl/FmwvRP7bb+5zzD7Gq/VF3dpbkQBU9Kv3+003QT0KVucEdWfgUwBsu
azm2w4tL7SBiKAXD4m820sZgIcIOYoxNU8ja2/nUfEAhrfOSEZ3RCDUyKoMedGjx
pElCK1xPCj+od50HlDLLFvnSxsHAJqTZDnyLerwZ1u0JCYyCwHi+hVkRSKj/3oY5
t703lZlFHO79YfgLj01ywHo6VKN5+x4w94DbHJmROdGFswXwyysaHFfmkXYSCbzU
3F9XZPLHveOyNEuRCiyRkhIN2RWKfp/NuHRUlzsTJQRkJa73iyxH6i0Iem6/Jebv
QuGTJRfLCvDY1+Ok4tOmYP6jHq9z3dA0bJ4R1pBNCYRgdtrKCT58RksfCg3EFL8U
CmlDBaU8JONSPFxvtFJLRx1/oeAuHSfH8KS5DNBuXLCxDqzNmTscqQcEV4auPYQ1
DOQAfTXkL4YboElEjy2Pmtu6rNFzIgOrZu+2ZTWEnaORxHApGiAvxduZU4eIIdJp
ByzkfTNOcYZD89h2EH4uAi3RLStocQqzsdP5Hq5oa0obw7UH0b87MWLTDsdpsRJv
DQw7xyIwTdR327RGNdEttLl7Sp/5DD4E+R/veVz/KjDZSW9kHXBV7EVfvMt9Oi3P
640vy/du74H+9cRNNPxsg1ZFbHMesxjrt/5wVSi+AcWzvu2wydt24qWMzHWETFu2
oXhhJTH0cNp7g1kB0ckOJ5cKQR6GImiRkpLMUqe9rCfEaVAGgemB2OOv1Kn/gM/J
yR+zHQGYedL97opNnYVwTR/6BOCQl4O4ii3k2YcxPh/HYQvJHuE2KvYxXhi8uIPt
3BJZE0uXKhNbuVDrFS6cWx5Mfz2YuFctKtEQP88LJcHDgMm9zWQKbBQ+Yl4qWGnt
e0PqlaLaLxFMH2hf+DRVXrwHh8/zk0hmwOVKv2FUoPyxWc39WOBMJyiGUU/B+Hxq
xCDY7I+Hrs0/W/7oCYyn93QzuJ5oZpzcqy0eEmSh/6FbeD1LCSfj31JKcp58aN32
EG/ZOa6wUJPcTC41/41udytxyRAvhZd5HYQsx0QEuwXZZ8aqmDaoSoBVBdYDijkJ
uzOGa7w5h67i0hmIHPRCO1FociKeh5qP8IGdjrWLb3h8quolQR2llWSXj6go7l3U
8zBmcHkBvidE7jL/alw2DfrrGRmvQUoL1326nn5Ydxo=
`protect END_PROTECTED
