`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3RD/Cb6UIvczNmWXr/GeBsWHBiuVtfUZYZJMagrHAm7AqqYs7NU45WuZqODp9H1K
R1iUJVe5pp8weKGppPklqVIixHaplQwfZZ8rjSdEX25yld8mS3ROaf4FOVsFk8v+
WCFkPM9nxN5ahzEjdSrCQ+mg7T0PI4GcUpzqgSPZW4OtEp6aJRVd6xpWZ4UC/irO
BKDpmcTBznfDxP3RqEh1/3R4nSU4RFGi50ytSjylnjq0Blui3Eu5uhX/7Pe2Mhuc
GEdU+uPMOF4cNqyO2UK0zA==
`protect END_PROTECTED
