`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yWvYGPv6YeBxRQd+UwPe1ZiCha07hL8FrJAXm0vT/9pV8lTmJbMMs5EXUkJX1e5G
XjPYNaS2S9SneC0ZFZoXBD+ES8nCiVXN2dDYZZcP5EjCABYcYYrOGWtBzfUJ1yf6
r4k61zhSLR5p5KOYth0GLXtmCU7OSSSYRBXZKuVE38TFKgCgl392p9X0OgeKBz3o
xArZSCqLlGackJw7zAbvF5fXkAkjSZXqraF5uCOq7/1KbawKELdKMYrzC1xS3M6T
wIkM3GZo00SuS91tz3UGhtEn9jcC562KuZnrMQZZ9OU3wwyzRcoqWM4O4MWl3OTX
yWlpTrExCQpEU1RrHv+7sGTvkwI07ioECBCMmT7nedQ=
`protect END_PROTECTED
