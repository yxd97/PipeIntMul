`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLrKh53eDNHkdgQX6vRXyno55ugb/VkKexn4ytH4WDclfJ/uuwV9ZtprGwx5wTZ4
A1jcUGYj6rlXNQ6hp1fPIfn4tdr8OoxticvGSXc+PAmT352QA2qSOKGuLPaPndav
BlKYgr6/s0+UVJT+AJpM83obBcozcwW/O7Ej8w4vnegbwEG8QPMCjAuVxdsv8hzw
qMglwzsAR0LMxRedKxZE85gUSplJAmfUkn9nCEixHTvKfkLJil29MTNlESgEmaJ1
swt0HwmcZUyQajbOBnS6P7CyRAVjSEN+KiwU17VGLcPFAGMBTD1hDpze+n5L0uV1
WPCc32PI22U8Opu1hVKhY7aLDeSh1+Xd0JLAIXqqUohAgIKfZFmN4lx3hqpETkHW
Xackp8URCuOcQWYkMMUBbw==
`protect END_PROTECTED
