`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yvR6DTlTvk4G6pyUXduSYNfdaC5aT80xZ9/+vsJDaDkgKtYBz1iLbKWhCOea28wv
DNKBoOhhtXgk/aY8rJICAadGjJlna1IOypRUiVEcjU+c+UY/Ucbfw7SM2qyQfOGe
k2UWfgkLHHoXZMYU10MuJyX2I2cMMJX2W7qoiszPwikUX+IHOhDm1f3EN+eCsprC
wuyuqwWnpJyM4/9jchcE4Xurxa/NLoWLqqXqHjxRrEYm3Q77kScBCSnFmsnHLz+5
q2fXgRAeJiHUvCEgHNEBXCQ0zbcoSWnFSc6DHFatnGSN3DSyF/tCYCG1dEm0CMo3
lxRzRpttbELH72FqOJckGLBn6WHQcSG6SACCgsTAtbuxrCchkazW+T/KLOlGRM9I
mQziCQn7udxSHUh04F7aC/G9JbIYkT/Nkaiuw8vfb+m8wOdoITWKuNLZjnUBC0Gf
uZSGYkCLkURdZY50RDRcD+cm3Uq28AG16Bni598iHtuU1B2dBzJtK/osTkT2w2eY
/7DPXywTjRhVcKJHVEb0HQJDmH9njV3KWXENMboedp7x5HLypNCHQfowEOX9lM9W
4Mpnwe5DpOAWWJwocPtgMQQBUFKjmNFAuSxq4nX14SccAz9akKdBFHYSElC45cVo
8wADlh4LmokKcS8QwUD+IY8EDw4suB2jMrtfNRYequKLOLkrPI+QXgjpVaLB0GOr
ek8XLLCod96J4GrLowA3yORGQEa/oAw7OykW4+tonvv5h/LoWcw/1LHS47OUuHhF
YIGjVD48citoP+ER0fN9FB6uKG+4Hirfe2WeGTljwzM=
`protect END_PROTECTED
