`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/mw0WZ9U+hk/nInRp4qc5KNPBTcIigoDTVQPlixtqm07odzKSX2kY2ff01Is0QZ
+9+duKgf9vILg4Voc82WxQY75S0VpX1WNjLg7nXOQdJtr1iJQJkUgBkgaJbQyiYj
tlm7lEU1BvY6pFoWghpozQuA7bC6NRsuy+adNBORrul7uZI+8drihhKqalHeGjgp
gm2iHOipZPLx+JkN49ETtLKDFvlGmggOT8FSY1yzQFXwCvn6LjvbB8qilHU3Mnr6
845936q19/k04LpbHEwv0JF1tpaC3V5Y7BCITYi7vugzx1FrGq2vAqYoBBngfqm0
GOeanze48ajRYQReEuJU9/XnP7AxlTJ9j/+MmUxYI/GRVyHNRkPoH3/a3S9zEi3L
iJHj/LSXZhL1zTjP6+BS+E6wIw/KYMRvfkEIaqAjywdmN1kr5mapFjTeqnUeNrA/
fn+KcrV1lxTCH+AMqb0eSZj8PlFUu+tfSpD0U66sf0tBXAU++6chumDIx16/qWbT
/2sWJZq7K63IfEOrqwJskUukEPilpUIFHDN/j8cvcuiOHCf9RvsRjDudyB2DFad0
FHRXzY8l/WnMF9AaNBF+ABT4Y3KlUzf8yi9Hroqf/Z/qZ/Csw0tNt6+8R44Y72uK
U/pt2u0zmJXi1ld5TgO5m/CprbDz/MDgherR260klNCeqAPfyDuy1xigmTf3Asi8
e8+OnrqmenJq7DXfeFEmKLtUYwl+nhB5FJoh6R/2kJN5zZ5FktL9rA8WOeFgI2sV
1ZKZtqi8d9hTNGzAXKfnRYhs3k7+fI8hq0Bw+Fj9hArqYRsYQ+ardXpHQd7f7IwR
V0UGqCiFfIYMD5rfhMTQ98io/UrwLKM3L+NW44dNWU2+4Waytralj7imgx0j/XhF
d5hd3KfMN4lxJIe54KBhUQ==
`protect END_PROTECTED
