`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYXH+74NRdNiDC1C/wtN+iwbYObipyppDljdbuyLTRrhgXQU1nu4iZ40gRenyQT7
I12pzMgtILHBFL55P0LUWwNIZi0t8EqGrRiNYxPRXCQ2ePHUEmgU6TxsrQyqWsMP
4rOLFawRyz8C9kXrLceKZZWOCujMIvfmqcQsMOv6NloBvokexXNLvF2nuWMgAAtF
YjVZ5qJf+GzUXn80hZePRzM1Zjr7rJeTELRv5ffqck8UZBL53oGV+5oS1sakYI0F
xFLRonoqRCFHyiccynEkSLRmojwp6620gzb4qn5fKOoyBlhyNVDbAGiS5VZy7C+z
Jk2WgdtfBFlBHX7rQ1/lEHfUMvUO/eBFIJ7kW9XW08PPEpvGuJx8zYWfR4q9Nxos
HeRv5UhBypt3nc/CFKSzmrY5yP/uE0UxohRPJuEE6c5EfVr+Ia9P6bSsnZWt9ljP
1zdJo4guKVzg+0nC4ZyMNFOnBrYAuxx1IJiB3N/QszHWnHFMJ6RsSC+qtyNTHF99
40mbbXWoUL5cIrsTbeJNlwgcuxy/zCIxy1DqzE8/yfcy743ZASiL+k0Qghhj/CBn
fIsO57Ix9n7DFLuSGtUnUXjCMli1408nzbIJY4OX6Mep4lhCz0Rn+Gk0hnuuJVmP
pWDCZy/4nifdcxJ2KcgsQe9wj6BneICqZlB8i3ufBBm3WkpPIkFGJzwQ1y+DAEOO
`protect END_PROTECTED
