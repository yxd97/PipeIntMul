`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/kaKJzYN9ap0FY9e3vErC2UR1aFrVmM/GktMo3aC4p7S47/fNSHWnD31tf2gDskn
QyX+0c33k06nFyn9UNsN39I5Uy+/O4RTJraNM7MsiFs40lKCwS2gLwZCWe0PfDmr
BajzYFqBlZIcsPCTS5efS59Mm1W9v3ivsyAAB14bFxYp4IIQ/yZ7XeHPyS9SW/kd
Se4CPFdJOYzL9IN3JPdZAFxirTIgsRlvKGrkLo9jdPKTIUnirnbQeSVNIJMiwvEd
RQepubAx1RzWAISGDct1HhVawPKwSK+VzqXKQJtzIecs+72wIRNFvFI9QdFeRKuA
uSQ4LRpMjByqDALLGZugGMAxeLMGXx3MAHFLXKnMXrpuwxTPw7O9I4oKVt7LTTwu
`protect END_PROTECTED
