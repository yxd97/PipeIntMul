`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlcRsAV3yrafNYzh8N94jAqMNjxCMQhMewvnd5eEXdD+jlNqyscE7OafEwydzTAF
JMQP8HFvA3q+Q7Wf5N0vYHbqGnUeD/RTrn+dIyZbEI0w9mr+ny1Nx/AXxISKlWox
qSLhIk88jZXdV1oImLbO+Dsh4rngyhuZxuM1MGhP6hnxkTTNQgGV1ibi503dBRsk
l8zyOpQndn85cGKfaoylD5eSuAzxevqH8RaAYGnxehjq7Y7j0J11mCZ1RkP9Y64A
yZ6sgLS7lW7pizjp3lEmJJqwW1nWD0oWPuXeU9y58j2CgbNkOq+k1Q4/se43qjTv
X1GmF1F5iJdYV8Zxu6FxQkgUK83g2q7S6PkQd9a3hB7XoStzXCVX1BEiuaQGohgu
mZuszQaWLDZWTuXfKPXgqTXZOKnT+LF2FxJbRPongDkAeU/q8fxl0h75LECUOzhz
Fg1UEW4h5UqaVjaY8Z6YnsS3i2+RunOjNp4ggGFqnYUcmegW3g+Z9MB95kGqnLNj
guE/dDH+9GIJO7SQhab/zC5I//Tsv63P+4aziigJmq192qz7VGeHG7s2Ygl6M03X
BeYkjywyVXz2khmg532yiZx93jch3HUi/hIgee2bmwK8TRuMITFCmPPLmyFSX3/4
OIQbgsWs498CxQWSYQ0sM7fzupOqK9JzIMz/VVdTl5loKFu/+10n/CC4azDvuwAU
iEvjgy8TKYC2pEEGXRRr4dFvv9W63ccvNkdYkYwcQ7d1e7msQnhcim2IWCPR6nHe
KoOPl7f5YZRcMm8E/GcXV72bDea+GFpHV0j/asLFx/RcjqhzDYu1pVAgZ5vaFnjP
LbSX9BKpCwSuLF/x/Lk6ZsiryP3Gu6nIY0urvmZPkGB9ib7v+wXuO3Q598HGWOXt
Cvwin+hkTjgexhcfebSVYIysKA9ffVGQMHQHUd20N0vqRVK5z+MWQrOUrM5dGT57
uaAVKu34k5cnpUILfyEE2TVEWXYem+qVkLHEiBbGJxM0CXY+WXZED11AkjFV8Mmu
PybhjFL6fgZt60n356D6A+ovZAvDX7dW8KIez0CmvelwdivesOMP61xPfDJNaTCY
gCpad5Gy2Vp6Y0LJsY00QEaXyCFOrvbwBOeFCkmn1yvz2ZE7MJKTn+LpIRnQ+lo3
PutnWMwCPkOmukkBn4x2gfMKMVUQU+gNmwVcK5XeC58CczWlYv6jUb+hV5Lnz1ia
q4fnnvUxlnzYzKfUF13fJTP8j/H58EPE3YdZCBiyTcwZwUUb7x0rq/j2CxVWpTo9
gb+5f/55oITdG9nVfwSbs+6pNXDSqEsUkzbJGuS8VW8=
`protect END_PROTECTED
