`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGJn7fwgTHFLqB1adjsXEjYWeURptUbeq5yD5GNlMMy3X8GurbbbJN+S0zqGMiU4
P3hV0RRlXaDW0FyNo+hrbC/BgXXrI3mkqYJBDz5S1tBIQyjGpu6KeLH/bXQibdLK
xlfIDSvjJ9qmNdbsxbgt+3wj0mROGXmNK7iMOOrSX5tnBGwKKgZJNeevqHj0k0l2
/m5JQLQM5tKcUA/6LZzh7BQeoNGZGTldABU4ATUrY5696mQBtCx+Vi+iBgtLuvzk
KrCPA2kuNRgdF+v06pgDDSQTvuQJDbCpnbP3n+9evaUrj8vI9KYHDlZpfVuyHuoM
IxrCsB53rmxisyKh0wWX5UK3Siv9fJHMKakImtxYz0tay8XOr+aNUV3R7I+7VgYh
76evwV/n1Emn/uVSts6XL8S7+4k8U/ey+BRoYwddOzCpMzSbQCdvkRPX9b2T5x8R
B9NYzeYU+uF4jnb1Y5beW7OLB4G3FCfnyuejqkIikmbFpSkl0z7CY2u1FQAUHrIP
rezvwpEgvaLRDya7Y16uFQ==
`protect END_PROTECTED
