`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XE2TYgdbr27H4oSWTnGON16p+rltIrFq0lQT3vrEcC7PKjwkG2OlVkOf5ozz0J8X
0GfrsgNLSc+yQS8xydpmvdatEzNf+GkU6IOqvzvl+LUZTK3y7FnzqV/qMYqYfDEw
W20bFKCZ1CVtKUp98MBPCxpg/XerUtklzgqB0brswx7Tx+VEodgt5aGd7lo/BP0W
FM19ZLV6/wyJtRsJi8mEzYUiMeBY/ZOjyR2ipFrnswqJNSvQI3F7Hcm7ZqyTIvZl
411prql24pLCyFJfQ88banU7jKPieCh6DvnADWwDeBtgawQGDEol4XNEsjRKza2J
jcnfDJrfoMimj2UfjBVGADni+llyTqVUIKSAsc+tfnDpNdC7cSfXweJDy0AHOn/q
LGs+SYKfuTFxIAmuoaxc29YIIydhQ2uEKzEAbRHZdGTqcmxBa/ZdcveypjcPt87d
Q8CXrmP8w12620FrlpiVtLqp1v3wNt+ifENQGUjdweSDtNWs6naihbti6dqhkCS/
Xe14HQGdsPrS4oLFA9WHIjQBGGUqH4nElq0A7SpIXkm9GpblcIpGehUykKj6sSSQ
8L2P+GgxoLBNDgMQIzO0oRxNJbfg2mGW8317QuHjxVwnfY0DmiF3+M1brr0qShnf
VSB0cEm8v81TKl+m3eJFqK5i/dH1zUqJV0EZfE8zhOJ8ocr++F3liuvhpzU4TYxB
9y5XQ3JGGxa/CTiOYZnmCu89rgNIgEgGcdxZSD4goGUGMW1uZzxSMIQow4CN+UJ4
DxdEd4o4m/rkKgUv3Jqxfo9aMB150yPB5MyK2FQ9obXqXYEWb0TfFa1IwjvFRJ2n
IqoIwlM5H942XK+J0hbiClKN81ZeU4iQI2CtEQZVH4Psr+A9S7d4m8dPTJoddgiC
DS8uw5qoRT0wdRFQLrOeqh0MI8H+QIYwpwRi3M2fJ89ckmYToePuaw+u668h+zSQ
if4JlIqnhJqvE1d4FxfZ+hlfA2tVnRLx1RH/hOAfc5PVrKWD2CVzyosznUnkzpY0
0OFv2C9eh0tD1jyGbWIFf+20u03AXZBwy+h6DqvIawZgXZ5LExwEQDcua0YZtrAv
iiVwXz1jo8ejXbnhM3AfshhUfbKjiHDJ2pHBcnjM0lRgUyOeH5ttNDEOplGg1Wzb
/x5WsTTHbqC6QJU+7hyvlr502Rx3XtBiuFn4Isu0OrRvqex43Ps9Y4/kbdmpQ5eD
4hbVuknXx7BiWul5Tz+HyCD3fIxxvbbiRDPUy1AHA0ttZjQoRPvT6uRLbZIEt/ZQ
SfsZejZDXrkQcYSRx/8fz1fIAeQ7qlJY5t0LQliELqWE5hN3Wmgbxfaxy79pIGed
6+4Kb62Kpz/YRTU49kkx077WOucOxm60ZKgyPQRdPe+V9sjCUi3lVfhR0xzNjr+i
lNO5e3evah6xI6GGs3YeiAl7OIiDyllbB97RSV6tb6Xbr/gOgtEspfnqjJnLwDy4
R0KVKQjnkyjrXtSul9tT0O2wVKCl2unU6fnC0xFHA1iZckKyoalLCGcyc4TtfqTZ
BvAGJF03escHJHBCIsKlWIQv/4/j5dQDY9JFaGDtDSpKUCwbvOc4+mXskt5MAltc
la59K0nI/bvq95dERXRPzWnSpdndcMlkQviqiLFP/av1DyQ24Y1NGHRiAYS6b46f
Yqqi8mx5DqaKR7lMSYut55qfXC3fPlPKmor6PvRFI6xG8MSH1ymiyhNCRiPx0xzK
AQYTkOhwU7hjDJVk6xTWKvzxo17t4BS79Jcp6Hg9ywGPSpEdthEzUjt0HbKkdCdj
lX60+0dHfOmLJPWJ53cC7LxS35h1DrrA0pkX64oQ1eFEwau+H4/7GElvweM/+gKJ
g8lXJ9bsT+AltbkdDJcnREj4Twjy3ZlSgMXjIBCjP95VCM49nhKk3G77/aMMR3MT
XtFncRlKkjazp7KTGLCJbCdH0zYtt9RiZoUhLHdlf5rdNYO7ogSBgyCpv7lHb87t
6tmcSZypjooL3o65p9rS2P6toLOzBAQJAggVyhgyq94FxREYHfF4ql0I1mBVrdH+
UI8meanssEgMNKVwlICt/0+naQMtxa2RH8dql+R5hvveGJiL7dELaok+WBFvoKkR
dOjM6Iy5SfYHQFRSNI+bBJy/s0iVRfeTCzXN2h+N5a+umsqL8tT7vgRjrEGnZJnJ
YCHh4ZHZ0BqGMf694PEJZR2VMAhGY8wtS2KJxmqBfPJXuNGqOr24MCxl52CadCL7
v+BXbUKcHKbNbSWmFOiaMEff+hMT//ZgtUyr7RksnsVHiELEaslIvfFlfLNBvSmX
GlkEtRsqrXChXmDsDM2ESjBlncvI8/ieS63CnQemp90TKf6tCQ4jRaPEntuFNLbf
rvIzEYv5MRt0WzxG5IADH9KcfDoPFbLkcz77dp96n84/OTxsIuk8nNJ/XbugQUJe
iUPUX/2/CGuVsKhzhOt9gbebbaHl9ky1iVctS2R/hL8ZimEJ64jBxZvMWuOcgx/A
EKL4C1upDed/Aje0LWDg37KFQZSYCJPpXD0bY7TLIxMxbNxZPrJxAHc6vLjk5flF
lPAgo7NbF+Xq2UAuxzTu2MUgg1hNgxeJG9loq4WWUcrt43Ur5T0IBMp/zDoMIQ6P
wqHKrKEV9q9FZrub/B5OP50eUac1Ii3Dh/im2RlmZjgqT3j/qLjrMfL40aISz97H
D1D8/E4mq/kzgjf3ZLOf6iyWhnjpN/gJVXvbQ89tFY/mIF269jkTE/MsUxLmFgf/
hBUpTUs+mAZjAEmmUuS3EX8c2rzog/TGDXmrcatjnGdd2X4I2J7jOR7tRGQ3wodR
Ey0bn61j82sSamYSPnpfAqfY/i+60LDetmw1WpjE2zrIz6TzM7S3DgLzya5jkRtX
Wk3kFgfjVUDdKo5ur93GbdGOXYUSeXBJbJwIjy+1+BYxK7NQJIm5NIjCeYhOhMFU
/EvkEqUKe2qyp8d55ZyFSt/zndFHp6amZPYLBd6b/TcBGCw69wEPD1NiQ3gwWhjT
4LT3/3IFLcu6Eg4m+VXyZfTazincs+YZ8D0h1St9vfjJvO00rWwyYKgLUgw7sR7u
pU7skZbbiV8Mof4xviboUIu39wF+RwC/mGCktanpBZWbUsU9b6HQB17IZQvIP5nM
YWKG+Q8zq6Q/fI+qYOj1nxWkxxMz/btOQ5Mmbl0vMuplwxHQN1yr3XXM6zFsrHJD
89K/U+pAfJLRE1OyTeurhWKxf/fCHMiDaFpyH5FhIURrjGGxvwybTIzEuWMW51JB
AR373vMbEPAm8XIeP3vAKkjKcGU3Cpu4PPoCHs82i06ow/fDvLvB4qhwB48MQ1/Y
Ph28R4/s6nxJBIyMqSYtkuYha9VBJ3Rh/Nn+21eHLGS3S84Ot6Ete/7nBC6k8xGd
wOFu9es8A92E76LTOOI7TclPoimKtmLf/rKKmwfL3oDVXx+soGfYqjFrRqytwIwQ
EjsveSSqCzLiuob6nv2hIpq5BLC3GQ/yztQqgbFziFyMOtBwBx1L71xDJlNciBeq
2LoXp+oDEYPr/UZt8gA4n1B1ObDDTXMuziTNjKLeLXRxM5LYYS2+QiHPRKJn4f9/
DzLFT02IIeeLAElXOtICe/GSQDpo9QbNKhFrmRPUxRtDacBsvHTDpz1rFMzfpO6N
DMoX6cBQwAGGXaJyhLkjHnNardSDlLjdVRCi6LAR/Dg0YuitGZxSdzvj49uePoU4
AdRvrNfdMxc5SMzfsqTmfOrWRMtieHeVRHcHsWs1XUU+6fRaj3ucbkdZwLPm4+xI
TPDfIhqVdPkOQryqGOO9yHAvU6dDg3PE0JkuZoIMZx8yflIqfzwJGvnIN9fyAtSk
VsIH1kzGY3UkP+3uQA43k3/MaF66rAcUnyTh4p3c8rK230InWp4RyDqMUbILihqq
NfOCuilRMflUKmJjMTN7qQi7EYIP039bhGu6vAiYp/LRyPYXplkRUm3tZdR+aqlR
R7Y9i5rIrkBgZIm3AUJE7KIzYCGvzWpfmUY1w0oSMSlRL7LDo14RdLOk9TfoDP23
G//J+Zp+NQxRg/XiLZWl+pfx0+IOTssOk2WNzp8Wt69uw5EKKEBuHtUvwV0gkNzm
Gi2wNTnzucJ6CpMsuIYYVKs3Rsdrg99+KCApEe3r05lA3VnHBfcw5dP8oCpOHnUK
fLHm4+36oUpPM08td869Z+GMYIYKva+IyPrWTUv4UEzu/Hvke4InzwleGGWekUUa
4j33ts22p2Bf0HTweW+Y6ERlbRpSYnQzh0wHeowXYMHoNaulCb0sjqoCwDBBsLi0
BnSJm2Feq0xGbMyTo769KvqkjaQG8O794jOqr0t8rC0cs0UkvXOytMn+Bgk/QTYh
C0N/HMiNBrM5yVGonyNhrPqMVP56N+M4cLSTVNjcxPtlYFc1CE9NuAgkAQaMzqig
G4wHXJMcSbmmIK5sKra3lsqg7BM63iUSCXXYDzHJhgGJpzY+M5+i3h1SsAAUMhWT
eJhZTjDiiOYsbDaEo9Bwpr1YRl+9rn/5wBDijP9ASuKXIBARAiE0qH/wrdWlW+wy
Jpvj7lLUwP45wICNwOxdIhBlIGKyzOxf2xJAqsWTl2PDruUUDDTXdFgJJwAP5429
UOYUGqX0Q+ZpLwqwnM4LrzjCkWouSOG+oh0ToBkOf3ljPsfqTiRSgBqVO/dQpDbz
jJN8vb9UMk3gxcgBPQhk/Sd4ROoZTgNzkgA2oRGibGLQlZx+y5NGQxxqGC2bsEM6
tdMlGvwDjT43AxUXW0rC/u/Qcosbyd7UUbBpUO0OENAtrT8ClwuE63XY6yIbdoCb
ks3TEoqwsTVJj+DJS8whdt5/rDuli1ey08mY51ZywjkvP+1I5Kr5TvoCcLYLPswE
cK87AmPY2NeOZqd35b0oWJpCOxLKkJB2+JdpmQcjNb9afcIAgFw7vO36w+LwUQyl
ntUiYPtlPYx8KlFFi9hKvI2c/7XtGQKWp0O1PCqerOrgwLq0oCvBMzZZhuY8Yo7M
1TZifnq2zh0zO4+V6ZMgOkReoNx/smpgqHieQECD54aCvhK3FlrAl2WEgHjgCRGi
56Xp/Fwwdb2StkCXZNqbO1AsTFV5CbW9m6B3x+c+i1CNd1FdUhc2qRg0OdvEnnIG
U5BpV6riJzDkWLOIYyLvGP8WhlNe1LVn+jzGs+VP3tIkti6NJTBzwEJxwLI4yX7h
FhyZ3VRl0pJ+4a9UxRS1i1Y8RSuH/ls752YukF2KPfjmQcNkOxUaYrSxaF6nLB0Y
qxnENK1nNfnoabZbeqvrgVt6qU/kZn8M1nt11W34hcRw1f3fSfap3srj9obK3/pp
CyfC2OGUwKUBJUmanbTI6tK3lKrGk3AG92oYC7RDb8NOTZU2YFn/n6MocVYcAtOK
HhbALMRLqD1NPQKqUgKnxMuCMmspPCxpRk727+r5uXe5xPaBl+Ok0NDZFAWofdyY
t7I/NwBiS80QBqOgrbmDqwRghYRCEvy74Y3rx1sLrFJYmr2MY3Hz2x5TsO/ftczi
zU+0+QwagTG7jT2Sezwx6IrCnDLFUnuuiqZ4OBpr+IEZRsRlZd8aD5YGYKE57a5d
Otfb6PlpCRp1ZkCwvtyfHxF+ceoLmh4WxZSnUd2os8MyOCQ1sBmsKlsCDgwqcMn9
1qQHOU0xjmk3l1yiVvEEOeVq+q4yoHfN/jrQ7q26dztlq7BdtpKEkUpxkLUe+zzf
63UUabYmXx9mC/63+Je5XRFmj5kWScjez7bYb9R8M9XsLa1pLuH1zX3m8VSNCLvb
heRXO1ZXLdXhpSyMDVkhg7TwY3O9hAyy/kEr7sV9Rk7avHEJe6CzREC0mHbQXnRZ
oiihEXXvISH+XBPtWMdBh72+oQqGqTtRvukFlI6wwtveVkRJY4JkDyQS5SwibRoz
o1rGp1LGPKclbMYM+zSXfiGfTi1pZH+OneAYlkzZTQASvZmu92mGZQhGh5UGKHOJ
+gl4HhsmyMFmOLEZ1/ns1Mup47vXFx3iA/vgM/q3lwTsJlbWCu8IPQ86PWw3A7Si
e9ntCkI1oo2hAS5waRQZpPmfO1kOtY8zXJqcZIPYjJHBATj9aIvWZBFXxzDsblN6
nbyZWqZLLW3g7H9I7VlkY0vO2c/JVTdbFC9QcLieIMiH9y2DkTbfCd5wRUNN5z5X
MlHrsAlnd491hK6mmplRn35CngofpJ/AKyn8RaczkLY+YexSphWez324mSPC8DlW
XhXdhfYzlCCvrDKcbVvKMvoROMgUWFdemT6aK2PDVVk8ZIUO8ovM6uXrK7znFR5B
cb2gFq64rutAN3JPRnQGjXGE8DmaC8iGc6M3CCI/kyrI4zRN299gXp0EdnjhkClR
owB04ej+EqbTjMFWZgqBkLhIxld7ZHfLfucZb2jG7U+Kkg/+3SwWGzvPABXwLN0i
KcsRLC6X7tXf+hQwL9bE/2w63eiXPzj+kpEcA54c7diJghCK+gdFzUaW+Hx9OTgf
e8aD+HAGZq+8uGhGNEq/sEUnXWfUM4bwotJGJ6qnCfAqR5jWfUaI8eMuIduHOTuk
I/9aNRo50mNThozL5CD2jrinSPUmLVnkm1k0www8ijWwsVRlPyLbC4vIeTqPsNaS
k8k43Y64M7OmuGAOCdLsHkbtuQAfXwVN+uWaPpzbucbqQbAWeFDYUCUpLzMnHZYi
Mxyez2y+q6sPbIwXV4Q3Pj6A3vvM7mhnswWI63YL6LUXIGT8wHaoHLs9OSvIdRhW
Cn7kXVCc4fNG30dB/L8GOnVjP4hGpI5foyVtrQVwJ90gOZEaDKLesoSkqQPUM5wn
bYYk9AN13rB112mTH6Kbkkf812774/BhcyBJx5X2C9/pc7eRYGjc2McFmxjPlr47
u3Swmiu2YAuO11GlUkVcf/4dpbJ6/Ya8dxfp+XhKkHN06bI5r/KyR5ruFbhhcmwS
qS9spDTZu7mUjpc/o9EwONp+qGog3JXoiVKGSyTaaasGjdMKrSXvMcAQZHYrrtOK
lI3cW6bWM5rZrWnQ9VwU6laJV7BFkWQyXBps7Pl9RQJFmA48g1WwJ1mOjS2B3OcF
TpVusZW2FaP0DWzzoEu5Q+brBgRCLR7wpRgqRX0IAalBwPyagUjQGx2Ef70GKoy1
1DKUvbFniwd/baiOFfgsnPPFI5mru95k1Ou/8IU8/NrYi61KosJxw4SegbBnbJtI
PVlThe3DORgXriaMovSCd0TsUuTSYsCmDK+xfF0arNCrf+HvcpkDq6Yd6GqbH1j5
NMEmhgSKKEpOpIh5uFHAL3v+/61/XAnrJ2hqRRkO5bp/GX9hsUvEDc+C+YLhHUWH
tGVoG+3hOh61v7NQfuST4iTS+OevORTJfgJnlPlkCaSsu0m9i1mYl0hl0qzVq2ml
2RZSsiJswU6+rxsdGwFlylrCSnVMhoBuYkEQF0OCZL+LHBVJhiog5MirRULrW0zS
svr/efrJP5Efl9CSoofgt1PP7fZtLsNaywhPoPrAVWxRrJYABIgDq2dubx/fIMEV
DHJYfJ3xbkKv32OZg4UgWlhT3cxx1cRqQp2GYGCnf6F7zotAb3ppGna5WgR3l2IB
QaAqIeyw2il/7UP3ClEudSU1ES7rzt3KUP8uUUy6w3GzXdmZRbaU2k9kmbxIJpua
scKCPM+F1x4c3jRE6+ZGNEGtCb8qFFsySQw7pxWHdVyJoJcfVUPB449XNROKF1Es
lL8lKGiGEcv8A/9tRDLZfuyd9S3/IIV8WB1fgSDhG5U1lqJWgtA5h/ilUo11b6W3
D02bATQcNNsYudWEoLKbPY3uGr7v4zsmFqnEenRUjGRig7J3LYHfDUbPpswTVGex
dyu6ubw3EjHkiZJ1OmwQD0sJtd5pQ1LMK5qI/BBmEDBPbNIms8QesL2egdvCbSXX
Y2+OSDEaQpaJQmel52U1qIQWpswTUoZ02Pc/cop7HkWEO2lfKyupz1RX8kbw+cij
w7EuMBUZ1I34mUAln8HTBq6h3RMRw3NzWiFGJ0zZgDbWoNyWLaZRoiSv16+wibdH
XWPERKuL09H8k4RoWdGyZHFSFHqxm/5lbSuLms/IBu6lh+upMsI0/0Fz9zX293Ye
u6qZ8vaaKNlt3BUPf+V0dSP8rFlQA9Bgnyyly5Ui64E686AaeZVxdcgNI3sffTd6
haDeCtOKZqgzfYhY3sW5LeG7tcdR5RDlBH/pk9UVR5ng3bPq6N/w9YiQiusU8JLy
e/mkmgTx13ABzr973uJ32CcNhihDTkQvrAs7k62TRHnpZFINBbotdCn/R87i/Qo3
ADRshRtOopvVo3p0BU4AlUnEIQTT7zGYcJnj/KA16UXgV4eAUTj5JcCvjJu4/FBZ
IOF7s05hrpNp2pryCPPBwr7yO2uNgSfm/egXZzp49KAkiPzpUj4XDYZLCbylZaG8
`protect END_PROTECTED
