`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XGjIWBu/L1B4znSxpH+aVynod4n9kf2h6mydXDCPAixnUz+iRcgsV8dRRODYiBEg
dNRyobWUlh+cWgu971GJ+JOMmU2HVkvFR5k4E9ScYMB0j4OoS2hIGmQ89O9lkfyL
PzxyEWuiFEwb31Lm5QOICudDrYI1JeWGEzQnoQb3a+QjA0C1BE/U5wh/XM1bSnC6
nhD+xiRJmd474nSSd8PkCKt2lVAR8SyHLauHIUWhiZ1w1Kxm1fViIELtMfHXgWvL
qqNCSoA3uB38XwrT+E2kj6w0wJOzDoAbOv/BRc4dV4PxgnPITzh2DTnampShblOF
/fJNLCf3JvrfEkKNolBGNjgJIGaQe9DGRpB76abzay+jvtHoRwS3eciefpNtkPHP
ap5nLuLjI7CN4piGEmnfHdsg9RDCo6fkiZyXn10crONrmquzx5pHRdgM2lVsiLe0
6pYucpPhPzzfvCRqnv2ieIQK4WzNzmpFJA4fCz3KwZU=
`protect END_PROTECTED
