`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uyhyIkjO40ZDW6s2Dd8XCRrH6lxPRPmC3+GgXHcEG6rWtdhh0QJfuYXdSG2qqOe8
+H24IoA5ktkcMrSPsMo9rLlrkvXotXkrhVLuQGGCejBSPmTReoGfmpmxodIwNvGG
up4qkYX+OqD/X/JvqUGEYG7LLP0OFeRVI9qa3JrFzPM7i5xq+m0zrE97ngXWwODj
8C3+6EAWe1QIJ7/hU52weM6E7aY4ElbwdCp1Ry8RuFS/hbQ9ZiAImrek9p8xcSMF
cEisC1VpQ1qv010uR0gPv2PpY8f3LvE6rWHLY+AhXo29Myx1p0db45fkVYD1UF5q
o79k53UyMe3+Fibka5QNxCR64bD60wjYjKwx9PMtWZybQS22ADqZSC2uq1ZuBBqR
APf0BgRW/eAeAIp2Cq93Pwf2HfldMplxL189wj6h4I0=
`protect END_PROTECTED
