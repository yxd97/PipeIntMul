`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWq4v9x8csTxU0PIqIEQFn1jSRVOy0EP9nhDrF3OawhvlIALwdvFBx/Eg9fnhYpo
4KuTVL4VsBIrQBNDt+csTMgu3e/gRSOaIGeAqP4uHeylCAUhyvKAr4KySGzGOq8O
hfNA6x3i/JrMP7+lPkGxTkJ6RZdrPXUbviSYZ13UY9IS8D/Bi8NCFKYpDTJ3Vmol
c3ZGOAdznI4SUUvi0Yx3oN9PI1Dr5DcOE7hT1jzYgqN0k6bKPaoFshMvaY0FfY2H
TMCCy9Mb12D6wf0GVH5nAW4YJHCyPGwn4SqYqoqnL8oirnEwX2iyxuBMBc/DjY1k
OtkRghm1DE2HT5IqyZUnMxylKs52uZx+sIvhRmNa1nG+tX3gp59/3w06ZOQvIrXg
6AMnwUY/SAak7r9JP4tcimZZl+qm1ehqOfrS/w8Uzgw8d2SnfGW2BnGk2N7KRAVt
wX/92sxmaMl7peQSpYQqxXlmftmnq6yFfNPmOHqJPtAk9nsdg3d19z8K+WWvwitx
WidaLmHDHG7c72ostHEkFIWoZ7kwRB5lYxxHOhycUB+oXH/WF0s3J8mF+AGhhqfK
`protect END_PROTECTED
