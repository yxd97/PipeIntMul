`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4sx9MQOR2dB7S8WVCMls5ySL2kH+aJefmjRBE+/Ic0DNIkVTM39LcRNl4pIDXl+G
YPCu7Q1pvHLsXUslIqEbpq44F6ucRb0ZaoKATQlsbIZzHdCSA3ly2I20yVaeuhw2
x0gyZQwR5VpECfSb2fFLrDXaGpJbLcJhT2VaV5z9gpkeeAYIp2g3V2ap19WhxXvV
DBog5obfKatn7K3iZk/lyaWhHYOiu9RnSx2TYl2qowpALzHK14fV8wSSy1C11cCj
zQAz22zltfw9dd+9/zUpXMq67dTrewHhylwvEznkgJ7Cm6EppVN0w4oZwnk4Yt02
Jg9ByXolYD+H+50UZt01RhlIYqb0Q/YFQ+He+Jam18N74qf7SR+I851VqXmMLlJF
Y6ghAvETjJpJU5iMjtTLZTHcAw36nUEhO538iIy47dJuBiKMlaCMhzhBze9ubOhK
sXjEOk8p8oYgUSl84N8/sOkqnUriWqMjTkSRNX6e6bRDXLR08rOTYC0NwTa60t7c
6aPiSWYzjR7Ftqbb3dpBl05R0++mJU9cX/Ii9UnNJyHyGCQGCRRSEQfszmb8LtYy
DLJqgT5vwdW3uzfa+4aZThiNU347U/9/0pQ9DYcRwlSC63Bz9U5WUxl4rnsz418m
MYJ3tCHsg+q/knEriBGpMJQgc5Q4qKZR5HerupYieZFpt3UFFehkdDrUSuCQj8WT
xL/40cAhah9RVNM+4yLiqRqBy75jFQM/EKt7AjU+JMvRpZMVyhhKuzQXtawrxYuc
VjbuHj+j73NZY2Pzsf/Rlte6ZB5fTqWJVmnp+TPrtXAqY1nKjAm/YTdNiQRwDmn3
`protect END_PROTECTED
