`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qH/1jWezlW3refXU2zQfnP9n6nmZQOytgU3SDoGd9sm/qs3QAHVx4lrBUNiCEyPu
hxRNJqMi8jzWtBV5WKRGnnGpr6PhpELf4FM7ulFruNvoN1IqvOswwynQo0HWL+Ah
9SRHTiQj430JPpTita476alGyrk9mQFC/X2HwX8H0b7/LcWEPj8Er1NxupXmeL5s
LTJrgEnWfwWtG5p60G15e6+YB8J6NLlegy4mn2Aq2deORxBBhlC7qdllRQLxHwPC
L+mDg5q/QFfOJEdpI0ljxsyUQYuSPj86zaRHePobPHM=
`protect END_PROTECTED
