`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fqwZoNvEaFo4zZBdbMlCfEdz5HQmGMbbk/a+4sGcWCa6ibg0rg8D15CgzJpyCKtV
kRLYF5L+richuQ57pXfMQCMmoVWpPwc6ZsmC6T5kGoA6k9LL8Z0228zAJGs8HuDU
BzdfByz4H0vlkZYcaoe6oW2e9KVEk73RZhq+pOTcLXCgWwz6dWBOwrjcdMNeL5zy
AKOIOZaF5IutmQk0rliAxYedFI/RcMYXRKhjImLO0TwMtsXeSbI1Ykvjxz5b31dw
ydnsZybTWPfG5Wp2hrGizBKkcKCD7Lq1oGQLspt9NL67+jq1KXG5Wp9dQfbGuman
0xNGysnYwkOEyY2/BfcgH666aZDww2yLMA95uJVEbT4=
`protect END_PROTECTED
