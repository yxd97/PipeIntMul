`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJuuDbFxA9jC+VwCWF+o3KpMalPhCMjcPuJ3jvtqGGeRLWI8ymOq6kSD0LM7nVN8
jJDdfy5T46lu/pvLyPFOx0rj/fY8Vk8M39QzYIMy8DbrBUV/vTw3QMwLwgBt95UG
JhLih5XQShGJIWg3vyuSC09cwwbTQmoN8RFQDeK7qulJEpP3kFIzBN7YkZQmPbFy
kwebLvCr7DqyUm7YNThDhWo58t3BTMmsOjl6YIgmEoXygZ3XRbgRjn4MFrUJll3q
gxL0SEcNyctibaMVX2HvKOPenvSuhhgETdssJZVvQedIbbnlufGjwcXpOjsDGVeQ
CVooUd+1hKvBaqRWYePNn8Ur2qWrG9F1BuvJ0ksF7ZfaxMu4qaMt2jBVZ17bDkyY
wqUaAhPtp/rQTcL0lU15LAzbm3bW2ivtyyTBDuhRMTym7xsKp23BGVIIP+KiUZBk
rJVwyRVfPNBBde3sTbrYEKzLt8bK26ELMamAO3GoGC/jG+aS2f7KAy0SjkxV4+jG
`protect END_PROTECTED
