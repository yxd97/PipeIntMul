`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2NSDziLP/ARPSWqZsAH154xN9Iswrv4m5YFCApC7GQx9NajIvHhcQn6XCDRLqsW
6ZzT1NdaqsoFZijT3hxWUbGgsIE+bCJyNdtsOxJzYyveyRyXMVzQ/dEOElf8/06/
DOr2oyFc2qaI7nmp1SEt+DGcA9GFSc1fp7WZaYyyoyPUskiMyf7lAup288iD84qV
PofhNyg4yhN0FEVQTho89KMMbg9QjRLRV8LDWxHDZ8ozcqChf8XY5PoRKnG1/Iqu
JT0GtEq4owokohMNKRwOkS++BTR2ei08kaMAhUYjePFA59kHcARIW9UYzHvQnxL0
Y5TWOs2kKKkQIDI35HvctKfCWHaJLoYh/ePtKeWbixF6b2FvYF2pGQd7XwgXnIQf
Mm1b5kqu7jL/fUK6APikg4ALhOrYo5GqjKDMt+DO/6CVluLIVLMLB1LFX0w6kaOn
12WpwMePPJJR4LWr01mMicsIh7gvzHhYRp9OfJdZgksICW6bxa6lm/GZLUctU9ju
HThgl4lIHjoqIUGlwd/gyUOwvnx5II0hpjOyJ2QoCy+hRLoM079uQUmGoBhduAKY
bnApqrvwuuqHMZqpwndVCqtvoodfjuUU9L8aNv33e5RNAGzSdNq5bbDxdlAAmPCE
+UwbhxuwzNTAyaLJO4yH+DIVrFSctIerWhxFsGZPIjZ656hSxDtg/PsRgCdPxom0
2NsMO0R5BisIcEoZe4t9PA+nY4d/p8+D8n/nFEzuesyvNEdeOJyM/AAY1CeD4okS
saczSEOtfWfl0LtYJOYEWw==
`protect END_PROTECTED
