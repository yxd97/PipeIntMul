`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cu9Dmj2of0nnP/rPwL49LOHuflZGLGt1u4SXfk19zizFdsd8/u6yF8nyXz7XyCj+
FLTlzS5fI1JFtD+LIsURJbUtDXvrWNE+W5LxK7qS4wKzyEnd6k8+9Vdi70Jst2FC
/FUNskaIxC4DwL8jv4hfuxa3PePe6f+FKreihlJoKkJd89E+nbWfoi66BPc3rtnJ
pOnUssp2jqmVLf3vBn6SOLzGsnq+88VOlqM1sq6V3Tj1X8xUvBhsyxHKpdrT/top
/QuyUNQa2x+KDjm+PTcyI2QkPhrujBQyNYjqJPKfMqJz/WhM+Nbvigwk76NjA7b/
HiAAYMpinqjahaIJqe9KgA==
`protect END_PROTECTED
