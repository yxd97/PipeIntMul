`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5c3rlrn+6Zt/8mQ4yJXJNei7Q6wiBnWrpUhd12BTHpSE5r6vKQgcK1uX757ssJWE
1CqWdPe27StpokMULsC5ipdrC0lTKoXeEk9vYZbxC31lw9MlZvylAYy/p5p6HhA/
7mqTmXTXm3ObiUXWgeZG8Dlfhw6ZbWAnzT3lm0jxtn+DVZ5+3AFThhW9fIKmp961
KISi5fHmW01sw7UC/iKcgqA9d1MIDgZMGwammMts0Yd6PJYIGELFww8Y3DTcRsOi
DTtCkT4uMS+DNdgDqNQZrWtm4t75PuCJUwHf3XMUqHM1qH8+17dXrd7drh1eCS6J
Twdj0MDssfZTgT7I/nfjqMnQkA2KMjqY3Z7tjlBIDKmpcyy+mj+V3ILU9qT1RmfB
e+z9KxYFM6xrcYfRmj+j21Gr7mzmz9AVm8Rsl2Whg8DoHXqLhPzrFLFFMkzCQjr/
B9yF32KRL4jx6u0cZlj5sFQlLnx81ZLsbQ6zxAwpw2w=
`protect END_PROTECTED
