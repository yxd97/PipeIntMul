`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FibdL2qYnU1Nt+rvPnEQG6tyrSadAWuq0Tz4l6oi4e0gRvMQ+i2V0eMnHQPolBCU
gykd0lUPlQZ7la547P8z8B+Yo4tMayFIcW5fEZ+ViRyatGZ9RKTE2DzGZbSK6tT6
JKfZUctAIrKz54qJc27sLsfbhVB4pVirvThdKj9sVzwAlPji+Q/cezOVCVI8zldf
KMigX9Zab2SUzLk6a0Xxw1dTW6iJclfOW19rL81XGfrZ9bTxDjZAIsaP3FkWeEh3
nZJlwL6DXo950PVFVM8XvJ1/biYJWrKZrYbpEuCM/qxBqHJL/lXC73X2dYNIYenM
GcGGcb3EHSNMnlxiYQqmo1a4AIDVycod/ynzLqeL1FfNyocNOHTffE1xtyc+AxiA
0B9pWmbKe/4/edm+dFg4GVIcMvuIOqW5Y06NPPRCmo3tNzf83vgzJq+nsLGarp54
Ss3uYXMtQUU3dMR4bQcVYnDeuTWzh3aDw8mkb9Nh/cV1sBcKpLlIm/S8j3Om1te5
A23WFj3FqIK7aUzZjHz2gve3x4SkqrCO4tuaW/21MnDpX8pWzrwPhtn0ZGpp3fNq
3FSOLsV4n7JidOQq5RzhZBJv+vjTkjM8JGzNro1mkHjWgtmGLE7WFL0xLEF9Tn+N
HtZlme/6pOf/lVpm/MvkrH4LkEY7luMywzkHJtw9X1cV6L3Y1QNG4+k08sj0Fclr
KApQZE3KVCCMkAEd7XAtybwJFeeiqEFcLOjoHbqdhurmnhFLrM/c/CTv8IXob8DI
7flTJ0O/OZdl7QYkI19NtuQDCT4SwMdlzF4zBJR8uMZJDfk0twYCLCu6eUi2BUdn
8Pb26AH5aOZEzIeejUYUEIaJLzjMuO1CxTc+78Oj+KS1rSI7jJ2QmE0VDUIthuGl
G9ODrvvgsfl/5JBAkjkCz8b/t/1L0VThs/wEnHcmd9ln9VWRGYjd3BqXUWDbZlQa
JZWlSugriSXAFceKKwTe4PZ/HpvVDwvrqcDExtmVNGq9jb3CkmoQxE5XO8/653GJ
7AaT+NwnoYkuw8dPYJ2u1C+JBXZCDxLW64mcN6C56gXp8hfMzmwzpaaLkIfyTbs7
EN99Dshh/GOLa6nehVOCiZztWrUlQHRZeiaZNzLjhCHntv48ZiY/BD7OPG1CIIRd
8oqr3qxDooxJ1eBQumC3HEjnEKGzGHzf7bvrZMMT8UP9gizFzx7+phKVw+41KS4k
AR+iKaC6+7VnxLzZjYO23iFaDKrC0KnRPg1Y2q/p6mIKe5jhuaXMGMgTUmV4RIer
bpYo93nfJrLr47ej21jjt3XOL1xuhjZ3Umd9//Vd1jDv+k1jArYVg3am2GmgUstu
Of4KX5JdOd6Bjrjxo2ELTeF5uGRpGTQpEYakVcuQ01cMMXecKDE8gPVW3VDSJHyP
ciIbrG/YbXnXL0j4Tk3nLgLs6gKgPLc0TgaOnl3EBC5Tyct3B+uM0oH0L3U4sJB+
`protect END_PROTECTED
