`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ioaAim3I6pmTfTNNiU5EBkEJOzqYEMMpL51N2xDwYRxMI2av/6rIpAyem5xMIkLW
zGu+1/3RnUUOi+qHhH0D/idMhDJkr3ae/vuZLBzVcfJ7R1iyQxOQFury5Hr4sRUS
f+o++pfKtcmhOj3Jg5ptOd71YS9gHB4xwubxLbdWR9ckl6JdcpLBCzGzWOWFh5gr
ww5NgveOCR6IKyCznLCMaG6+KRwvKT8WJpbHIaWzVK9jEVTRwgxzzkFneDMkPKb9
K2YlZ448SnSFYOeXXIEXQd3j+hIFpXBhP7l2z7Ltp4sVWh/TW3mlEuupGOBs6PLK
5EYkdsQ4m7LNXG5lwzJZv/V/FyEAdE0vIQkSK687A1a80YLDWS4u4v6fklczZxCK
j+zs995GR74sWnjd1BbDVqs0zmputI9Abw0WDQgoxEddLZ9NyLeOky3XaCRSB2wq
79rFXatzrP1aeR78ZtXRBodX8oQkwCbtD+tghUw9Rtbw0PQxOiaDxSmawebGqNqu
wvhQzacwGp7BFhsXfOJBKQ==
`protect END_PROTECTED
