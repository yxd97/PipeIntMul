`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pudv/akuWQtT3SkYlM1J89Xc/rkhq6R5OimO5RlJwbbJCWiAZnOY55hmCnxQsiy4
pyzBcHMxh8eYEzSPsgs2I48nDv9Sj9tgZRtTz/ypKRC5daKKtw9K2r/6Por4MaP5
LJQV2twCuqT4z3KTCQzA44hZd4aGhUjWnD+bqrKbUhlisa8FcNghfyTlvfxn/WEs
XWUK5hDjPYIxPCk25DQKfHMEOb6vMC3q3Jk6EsgHTfHVvTDH1rGHZqT98+ifSTzG
OYxLAuWsrto1htElz+DFwRi/CozNmlwpyE3RuVq8nipkK6SUT77P19NKuRJC+n0P
3kYBMl0Rim03A29Xy3Od7iP19y0rynK6bpASD+Zbfy4YsfBsPI52bcgII/YnhYw1
mpZi5/uLIm6yz2fJLnYvJeI2glGsXRO+9LAKakxFLowwi1jE1eNpzWYakvV/t6oN
GD4v4jfz3vMtMMTYckFzqRiL9zo3IIasWo1uqLHYICNPd+rnf1K62bBkjxyiOheh
ZR5BvYHTtwrzucY7wN0yikCrDh8Z4FtwAXzoBO+zTnhrKBDKlaeGPqDqId+ltK7V
OyCawd8k7pwj0u3ecuU++OjCERJaFI8OA5f7YA26xBvCUJ/zyeUq0uqzNeS2OIi4
XCsBuWh9ySSq72CiJSMNQw==
`protect END_PROTECTED
