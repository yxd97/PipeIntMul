`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WkRhoRGALIQNXvKeux7cf3u1jufdIX+gXd6mFKOzvF41KoujpB/2nQhPZZD2r4w/
X0LEI9hoi9jB9syu/BaFk8SW+bB+JcwzcNi3zPHPKyivq4/2eA90AoDJS9LbAuN+
XirxdME1LcMuc8kvRMy6jOH5BF5PfwvUHlBCU3F8c6ebkAR/3KipY1GIKZZm458h
5gSVdIX3PL8W1Y6mnYikj+4byfb3bCpE+HSi4o/diTH1mdzyay4OW6Gfor4LDRiX
xOS+GWFt5GkrKDrk75pBLcShG2WPh6iUvIAZFFuYRcMU/3JdMvt8eQ02EFr92VYi
SHJnhxMb9jgBg0pH1lgYo8QkTqal5/xX9MhpLT41/ROyB3e0KpFJflsfUzx/37Fe
ctI1rqjlQbPumD8FihB5uw==
`protect END_PROTECTED
