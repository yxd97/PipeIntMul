`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jX3vnHgAp4dlKeyNsUtWVd1JR7DyZ6MSGKn5wv9weqrQmqwuycLujsJHm1xSS0cp
YGOUYEMvESHDtT9H4xwcVo07e5IJWGFvWCO+xYDtSVRNRr/yav9y3UE1TprN88dJ
NqhScv51Mkecn227mKS29g6CLkZ1vAdVAZdEEKFVSJ8vcWkqA+4a2qMjtq/2OZ17
3e+4CiAXL1dfzTBgnvXhYiRnKeu/N5bHzibHIzFmgnsR3kBqx292Cv7v0JbppIiu
+gcg8p480K5e28prxEmozts3vxiyQGDCT359kxe9qa+9PIPWp4OM/MFL0dsdlwbj
uJXUfl/ZzVavlLZf2dYScTlzC3Lzua+2btJqaJYD94nWxd3CGR0K77IezoLbz2n1
VnVS09TuMrR+rRbJkvkgoOYAwBMJHKSvnEnXkVOfE7A8yjgreU4tDbYtk/CHpUTs
IiDfT2GdOB42nXxcTFGR1DmabsSj+P1LUSrVsbhfNYPzXAb151/q0XwjkK6/9JBo
izR8UN4ZPI3qHqCMLAsKBc4+d2itiRzE0f2ll4/WCdv25b4frYdKJKn3gDBrKVvK
yT+n6tyfrAj+0+b2we8ShAuhtivzqsR8O4WELq99txM=
`protect END_PROTECTED
