`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0KBXKUf5PPshIGNGVVI9L9mrd6QW2PzATs/VXIe9MHhp+z/+NhjuFPXtY5vVKoj
rRbsyWL8eMGqMh4k6dO80wK3FevA4tkN8YUYBcbe1sfjLa7BkmaoBMUYDVN7J0oz
Ozy+dH9QjsGoHxhjB6X2e9/8jC59MkzaOvFT/kwvq1Dfmd8rrG7ni4RLk2VK4tSJ
DVQKUP6LVJzhQODLuuZcvrp0Dafdw+c+TZm1p3nEmleCT/uovwdqpPpAlHYAiV+e
uFjBUJit87vXFdWYS6e7owzvIGBod86kxx17DV34hlG6vjs0aq4O1Fw/MSszCvMI
P75QdDcVw/+YkaYU8tGtvQ==
`protect END_PROTECTED
