`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AFDKFUf8Wm18C9Cu8W8OiKk8X0kgtFJTl2n8NcCns+aRBhxOMiTEtlDeztVE9VQ
C+Y3GL8l75MGerVwCHPoiRPW4xVPzsdJeqeoORypMWVyv/uz8NTNTAzsMov+v9Py
RgcK4RoP0wKivtaEHYtbPonVBYReSFSY0Go9zHqFpsrf9k3SCP3dT/QjKfLkB5dF
g1VrSsGJsfal8xz0Bvq9D0FvdTKB24s9Zt+8p9gTkObJw+/bhBcJeLg0A6cBai5R
12sS9XfWGsYDzp6bd4mVYxik1SmLpakFE62dNJ8gYkuWWCcja8uTyuA86Z+yKXlt
hZ6xhJMbHYC+YgBOI6BLrxZLwPzRVMDt/3hmvgopvqBMYuEi6nnWZaKUYkuGsKV+
`protect END_PROTECTED
