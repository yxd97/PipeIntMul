`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLYLNpDtEEEkb4bdzJUv8ob6JnkBRq5M0UTpeTbRulgnJQadQRRgmJEYwvN8orxY
jMaO5DykiiFajeoaBpQ+oCLXnvzu7T3LdPY3p5TWuhElQj0hiamJ8S49KJwnix9p
EFTQTAs2UtUyXs1F6uszP90ov6NEn2CuAxrTe4ab7zwQY2eTrl7yonyBBZqTosid
U1/tHbApckln+F0TRTM2FVa43piDINawON0usmhQz1w+OLER2mYIib1LZAJ7PCGU
bsHkNk9jLJkGEZ6SGTfQmQGshc8XSBrxU06Jj7+MtmQ2AG2i2QDYi2cbG009cDsi
acdi2Te2qiqFSGDL41bushdGTyt71ZKTvc561iCYNqjxiEu6ddyenITVfI9yJc7E
WNk0/KDT8+LIxQhPGThmnKXxL6czX0xS4mWqpTwz7PXkvfuxSq+YIsuLb+xhqMOZ
/ipP3BRonOWYArch2Aug8zeHIkWjizGE40fTo4lqiSxyi+ELvCKsbPc3jaViaC9D
u9MZTtwnsT6LKO2IDJpKk2mSyGTQeDWQXHnfco4wELs/p9GkOjCU8VzX8MLXFC8E
Bf7iNo4j04IfRiv+iZkBFA3Oa2wmXkwkm1mliMQoB/8=
`protect END_PROTECTED
