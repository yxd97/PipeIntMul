`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kw7tWk+uggjPAaoblnJlmfNL3INJrGJR6RmhjSz2y2anOlTcUiMLL3UPSp5EqWh1
v0y5k0qsW2a90j2TcVai771oeIXcRvw7MfVY4zrwS1jL35wVTDKYDlppuLff6e+R
r61WHcXj+5KmDi5WXuFU+9GyBLCQ8Z8WaxEU2WGMfj1ifgVjP3C82BbZdnvyM8v5
o8F+c5oxXfQsiZyXK6I+N4c/mXVU7V2HvcHa18DFQ6quR0qxSFdOOdo289YbDocF
umFwePcLO22v2K0Ay1cfE/5b5UuETkr7F5eD1275CYU3PYZTRMk+VQKUJqsphJPW
7NZMGUGgcWUSU2PLJYJRXeO8UsEQoWpnO93LIckB2DNxDcaV1jh3yMH7BLQWBuSl
VbfJyybrI7hpHPFwD+L1AR9QMXb53mauEaH/87SxqpbRdxZkNAyCRhKU3Z+vPML4
DdStTKJR4SEIHlsPdefgp0tg6bLYFjzofHuskucwkrIX0HbDwz1Qve6exbX6lrsK
3PkrtnwRdwF7i4w/yruiPxnKYlYmUN+nnndXF5mnIunHnifoTmtd78Jm3XIu4QY7
SysPjdJPdxuLrm7e39RYPZh0d15l2kvRD3iRA1t5zvmWCZjK7FCe2AZgjxeQUZrA
cOvaIndfNBBpaNoM7Gj1nXJVO5QhdGT3L/Vbck3VLH2Vsl214dfRjSyOZd8Ntm50
OnQtpmQk5z5Kj3JuEKwJ/WTjY3tNTZg08SgskLmuu3T+4i53HCwNvf5HR5GbO+Yp
WsFYkDEt5Ni22xujL3tZsaQjmbsUP/9v7dyDaaw3QaWsHadjl6bvRjA9PZIFV1Dx
WJubUlpPA5aqRDc1nEQhefTsfrNepLgjW5PHwaP8/CBejLPZYdajHehih6zibT5b
YX1s/EY8yX5a1zhnCPDMLJtgiqmGxZP/qBE5gyGT5xe/T/fk10srUu8x2HIUEcdZ
7BTGyhr/4/a2O0HVWMyzWHaRTVSAsSHR0pwLtVP7MHg2wIwcbGyes2T0q7KJKem6
bnEe/Hti0lB4epBRb2EHATv04wA2qLrvBRfL+j6AnmCl0t39L1Lreo+zhOJvXSdH
mv+Bi7Iuc2YYUEeRBVXGYGHQrBunKHSDwpa1ogyXtemE6MlLXOYIAptIsFQNSd4l
bv0eN4YIrhvBtUQ4h32rBC6tPM0q6LTD6zy+aMOB6i9qDTRfo0ZxVlnyHNmsNpi7
7ZmXmKkb+294onRhA2SshJWEofeSIRQa4ShBCNDYmAqoRRZoJh9MtRqeNvg3SR3e
X5nfpy2vzpOz+kB2CQFhg4ZqgbHjG7+UZaK0XXk0Vjtu2OoikSjAvc9x0o4H6Nr2
2y96jDzfKEpIx37poUN8OtyDzhREaB0UcHelABLPiqGXbsGqpiYWG1T+sU9lODh9
HGGzWrUvYVwsMBEBUlXX+6QqTDBGoSfl4Xa2GomZaGBnGd66cc2mYMU6geAcb+0h
FT+bxigPGWsxsUjJgmQlNBcY2F6RXUn8NAPcdF/16ekg0/8phdgNMdUIxVGbmfaC
FKU53uoIZme78/UUkISN3n+ey4yqql4iM+4bp3OmPJxxGymFRPpNhAYLTasbKZee
E6K2EYm87msxFdFGCCQzbMCEPrZyYFUGx8GdTmJZejBiD+zs9FtmVChxNmO4LPeT
bQyWIUZ3HHhylpHiYp5gDt3csmfXiDdOTBwgZNDXWYV4yLrt2+Fjz7v3AxTcY9N0
J73Z90fyxD78uWOMvD/KBSsmk/Yi84OUSjmGEg4R4cMT/E+FpgCK/bBMsDZhudeP
6FoKbx+vC56CWaJxCE45EliCDyox3L4IvWUEAGm6DUTvUnmD/kbhsUtxMkJI5cjD
cQWCleiD08hvWzsI/ZJ60VnDChpzIlreom2vQOWmr/7oZ+NuxPScJfEMyRKpN3V7
S1jL8bfn8QruD6nv0ZnAqby92dEqXF5PTXXe00fxkn0l3Py2toGIUplX6k2b38as
CnZDQQoTV7lpcgyFy3RnQio2DRILCdjpJ8DS5n8piyRRutKLDNE3z+/cFKJG7N+r
Z0W0N2XWx29onh684ilcL7cK2hKuiKc61XOrweqVc9RRtU899MEad5sXK8GR2b7u
asJ/S+6oPW70j5LTc1NvMtZoVBkvbJTTTVcKr1Yh3TtQHBkemiUR0vDaznEcr3BD
wgtTRQth0msEYN7bAflQ+zE468ENmCHj+43QhVnZUXj6dmA+OkYlzsOhejb0BUKr
/wNiMN1a39Jhv9uJYHojCmVrumEihOxHJFPH6yg4tE2bAIQNqOXvQkrZNp3rY99T
hFGHi+9z6ygt3E0aOsDJ23rt6NujNZYfZ+I2IKq3Xv3NpVxUYI2kBzXLnyK2InTk
MQeqogukeVoDd7yIclN3rb3HbOGsYKC3vRbD3kiS1DA=
`protect END_PROTECTED
