`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hhMpE+UrcK+HCTv26ip4WMqm5rmsxC7ic58f4MQgJaxIlkxECcUtNmBTjc8liTlu
etotTyZ8fcnVISvIjwQnWS2sFKHV3QVAdLWOinxMm5I+5ze8gubVkiVT00i/tX1a
7ONbZFN3F9oQo95vm7ELa81VNTzOAMLEjjiHbcTHXNhTyG6GTVIAtuMqO1SdyXD4
c3K/OmxNk7FCWbezy4THujKXwAUePPdXE+/T1luNVs6hXN4Y1U/nz0O/rXHs8tAQ
R6s3K3BPZp6A1YtBVh9IvB3PReQyZJ7fCPn2Gmiwk+PuqEFe4p0BupsgZmubmH6L
wnoH0jYbecyNrAQz+00A/8JFRC8KNj1VALa3dBLrw+Z2tgqNZrXQvX2uaPhM3atd
Hg44A7jIWrPgh56mvLEMzHZ2dTm4zJTM9UUGz4zXLTqDE3WRieW/IuNJAtC+tpvY
97kXSPgynKILqzhXikFNLsojogcrD/bH4/8qNHKHj1KlfGLG8zc/+JdfhOGl6+4k
6WWgWK6ErLqRrjzAMsJD0CMm7zP6O4nJPc+8lkEUuQBni2ELbAExfbXosmQ2R5in
/GaGd4lkoukMikx+j9mA9/vIpdUNUYn66rwyOe0VNU/YrQNBhHwe4F8ozQ3uYUq4
v4Vi9BHG6UXm7VSXj+eSZthVYFdubhG1IWi445e7icezmq/Q4ypwTFmz1CUpmK/I
9dkSFAfjQlRC01rVl/Xv9Y5s0v6ToTvXdcHZZAr5DN0XiPBbPdHlCqyOrl7/Usqq
ATNcUgagzQxUbwPdj7YW9zEJou96JeVCv7hWdaIK1ElwiHnyVBu8IbmrOT3bx4B4
s0FrgG4LJ6twzMTFtETqPLh7pC2zeUSjqMVHrdug3M1jvvOr4k5zd23vIS8Zm0fM
hfRHHpeyQuwGJfwILkwy583rVzlOtopghqTUVWM0W1r+P1rHPYRHUUrjN/zkjFsz
eG12+HerqY29Mm0d6EPjRQ3omTsNsCFd6CbGaBRrGbVkX0QcfHM9tOLv7nhWxZ+n
YS9A2wq2VkgbXN9UwPkvrHOHg8Gn6op1b5LxLJKEW7g3F3YzmqOmPZlxUPtf3jNw
sRz9b/QmkOCI4Zn6EP+M+Oq8htSgGMzck5tz2rK+KDZULXWJo0xvzS66K4fQWpvZ
rZpArS2aQUMagWnG0g4GbhEy9R26iy6EXu9dheNQkdMUuUHbb9VsV9PyeFaQmIXl
T6zA9AQwyqpQJ4J0bAQod6V8IjmLGw29wD6AKsp5rnbMR2KZChPFvbdUAMPuV3/3
IWT1Affzd+OZR6geTtkGKHC0Db4sRsDXCi494/b9qbej6Kl0EDfVFR2WDmAgU8aS
e+xb+NWJ/Y4Bd2bVwQgc/xg0/0SdOVXerKvvm8yk43koUROoTUsprggSADFg+8bF
zb/D/zBgp+DkKUN9oDQB51JdezdVKcOjHb/J3meLf51J8kAdGE7F5kedbiWJnjZS
Zf8lNM60x8voiT1QBU7/so8x0wzCmoWfUGuHEzteY9pGk1BjEBgkKjrzd+knJ3kY
gTLJT3z1NxzG9MUT/Kep3ubjucQZFSXrHcyRTrTZNvNDsEU/ycCzR6ebEKFNDjNJ
0zkPqfHP8XQomVLfDis2sE4qaB+yUnwda0/EAAoBjP0iVO5NY2Bgxh5Aa7z7nsaN
8grrOgxRPUgRzB8Wo1NuaFyEIoj7hnMCNDdgOu/u4nN3KBsYcgEc45hX4GTR88PZ
1qt7WI2tjKsf72uMUn/fWjgAl98wy02HVbPVoSup99r4Cjta9xpexqAjxUkVKXrZ
B8BrjqWlmolTQMI+bKV6n+AyQ0ctJk4w1iWeMM1phPu+Cz3apwgg9ZWZVqfgtKx6
Bg2bDtnvXDQNFnw1PZ22DpzhTeoyJpGGXDDmk0/O2s0gtr5rv9I8ZN7ucNYhvQTR
vrhwCYUfp0JI9MEOpuwj/GYXmyWj1ecoyUKYtt2zf5a+36NZijyQ8sEl+yn6FPpi
aBweVg4bYK+P4Q+N7rCHv/SXWnhJTN30FFDkRxhuP6la4u33v+dAXzS2eYEZoVO8
XGNj42xREUrz3NiP4mw/4L27OzZV/nwCXkDh/3pH+XCJTm9ycD3mrPgGuGoVQCNS
QagpsAV5nqONwAJeTRsx2tESc11TmNd18nU5fJ/MjUaReDR5kxplF9+gvw+eHchU
lYvjEViJ4wyx+ccWJ3cjBfEOuFe7lqaiM9Ht0mkgkkpNi4dvwMm89/SfjeTq0uv6
ypEuCs0eXZIFshLcJ+uSevfey/tsFgFx/FG/aUpQXBwKWbzx90SYRq8Gg6LqW3A+
8EuGFYD+m5nbCpbRehm/gFWPRMz3ep2QIqTRWc7grLgk2B8ljTywfJaucmcd4kMz
1jNu63d254hBkzhpBMkPf/DHZ4d9bS29T/9s1sDIhmyIRuqkYiBzNiB9Z4ic4xws
B/2WQZ7RXBR4yY4hF0PR0VUU4ZsQyxptIHuf7CuaVVgFnTD95JWjZNsgvmBKxCFK
TMm8u2owO5Beg7jvhMFedasc6j5g1UJ4AXHHoyBajJ0kczSoxKnxoi1vDPgk63WX
0fjpE9oJi3+THAQNrPiPx5vy/H2GkNtPU5+kJs/1OJlC965mrMIqjKbyFTmw/met
G/IBs21d/eJBUG0dCD/88WOWcinBRhApYhMoUZJSX0LCppFCk4P9lappAVvb9uyC
HDYSEnSQz7zUkIgOnDVVt5v6MdsScVskySPZxZGs9C3YZmcfPp3hZiQ+PP+/x8Hq
uctckuE9Xi5FFxTRJW6ufRB5VFX+wR3ORkNyxu9w8J+RdqxMvTs5F2yn6rrlzqdb
eg8noO0AZUhrXdma9l859d/IWH3uVjOAwIfC027gwe80rUgI6G8CGMr5qUdUlJ5C
m4IwBNP62Nw+b11k9Af8s6iSPVdp9PQunc/JAYv78lTvd5zkhjjJo2K3zoWhTbNR
B8dqOMaYKugskrLE1OMSacEi8RJBjqpWoM7b5qe2puaHX+BS3S5lix6SfyfN8ZCt
np13oq1Chk9iO2p5l5FROgK8XmbNSRPJCD01Mgpegrbh41HNK4qkCthY4xiA6eIX
xjkeyIKFaCPwoERqqg4EYGomC4TxypAnFs/ACSYEKVX/sStpduo43AdLppRKMHlJ
r8Z+LYlzhYXddEGMcT9yYOET3b/fIRDHV6kPrACjMj6it9Y3Y/n674h042tSGVGt
HYaLwfYhQnlcULx1ecMnL0btufNLn4AetZoWtjbK5ITqsJig3rXO92lVRP7ZXI8a
NmqXmzCnX3V7eOztTQjomOXAs0RLUuPndXPwZtRCd6cKH7vFTbELGBf58PRXzbSp
pw6CnkswLO8G7bWtXUrLgH/rtQTdLnV87UBsHAmoSq09kOs8kkDWVrdpYXlRQcuZ
/hD6fXwcf5bUFvn1YGi/158a+ibK13wSGPrMgzTx6yHeMjL+zX82+jvhojkeCmqr
+4ulIA3zKiulaUGpHOtnBxV/ER1/uwI0P70bJd6JMRNTeEBBFQb+SBYjianEVLDW
TqXeSkNgeabdroSaptEkQJ+/rbjozTS7Ai3ZyMc44VimycP0twMshi+XaJk9TSsQ
SnlzwoXCx1IPjAykftFKjjHqluDI1eUsrWcFgSCwNmqntuhR/zy+Y+Nbn/G9EcZF
4qKYv/htUy3EXG5lac3WMDMShjhHp3ULFpn13Lhxz/3HL86gAqakDOv2t+rAX90o
loHYV3rgzkwxpcGEkaM0W7lVji+WbPoOctz9Cc4wWzeGlVd3HUQZytShh9+JqiB7
oxH/Ch6KMwCnfEK+CPc5Rfp56GVHbCGOfoL2uZL8PZQ=
`protect END_PROTECTED
