`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BVppmeL+IJ1IOJsxd9R92jZZxeekDE6rAgnYfkeALz6L6kqZRRvfrwoDV6Il3+CA
jW8mjypiEBMsRF01Ez1XJWxTinA+7gbZoxOdMMjmZew3ZHjc1RyeszfRJRqC1Qvl
Fiv+yG5n9J2xNRKRu3tH4coG8QJ8kfXnpRy9mZCXnJZt9ppY3VFbKUCiyUfoWzud
OrUOnwLMucMEqSd4JPIHLAa1jmfkySsnLduGem04puXmoV0vxYRtjorjxGPu2RUF
VzGqKiTK4joy9ss2FjuzV7MwuAz8I/5/kLvzZCCAP6CnFJj+VU3j3l7B+0DxM73J
`protect END_PROTECTED
