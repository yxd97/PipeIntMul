`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLtxRZ+g0P5E12yI/jV4BFtwQX+DdxtKzNQVKZQmy6odsymDNBYN4zvKg878dix5
FdUuC7eZMdZvFm2AFgyMKkFmMUjSMp89LgWFVU/FMGgbSFXLzfZA5u4mmWcO4LvJ
Qt3EWoQbrlRFb22TS6st5nsVA92xLy4Xuu28N9FeTt97oc7oT6DRDd0ueESUnER3
1Xd4HdBUKe6gYJPUQgJHk6ynCDI4ByJfh5+LZZr9v2HMo65eR70TLa69lSl4vPzU
6kcj2w1tMYwamfJEVl5a0AU9INxgwVBpKNIUCbr+PAhSh6qd0nlDYK04Hg/ytPgv
+6I5/M63G8OGza2pNprG/zJPPkw1XjlWHC/NQCw3oYoC5xMZVw3nHD++TFfQO/pY
vK5ej7v0RDZ64KYkevh9gw==
`protect END_PROTECTED
