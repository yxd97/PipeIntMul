`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3NibH45rCFWzYJhN7EojyJwqv734+cXbrieaijbZ69/7o/AFwZxZNXPJDWBXMWLu
/3iDq2V1SkVMTjwfz4JGhN1qNjNTVnlKraay8p8xbj1qjQpFl4O9LBuF/KTbHd4B
yQ2T6j/Q43YBgKo9wT92VLCBnP/l86YtYcne2hAEbTID4pwjhgZUZG+cXjys3Hsc
9inlhYZ6o+/jt7/xK0N+GmX6IcSShhBYiiBRAfHicoHhB3EizV94eg26RK4jIcCu
zdubZ/uHWqq57+HN++w1zJFPbtwFoGKga35a1BDkDzHTlfxXSiKMN74ZVVmsHciR
mpmLZpQunPeEx2x6ej9vj9kZNzK/dNgsh0m+iEDDh/eTJmYfDJvDsDwW8L2AcT/g
h4GtTzHJDwdTK7u544uP+5+koJO1GNINvQgZndUkSrt7KqXaatM39+FYWczKhL6y
QsX8X/FO74ZVrchrNqAFwXcd1iX/Z2r1hzB9CZy/WWDX2ntgPZY1J907y1xN5BDr
f6ubIpp20oJDk7OqGWpQZBOD00GYlDXQrmWy6yFdyOYJvYd7GKWvH73kr2XIJW7O
dsaiuZe37jiS0EtdMjib4OFFSV/f+NRcf+c8jEUDTaOvrZcxxQiWlhD9Xy9T8let
jyL0k3VVy2x1vO1dk7D8UR0Th+f5NDiT36kNUDovfm8FAoOOpWxMvvLMxDKrplsK
jeWHdn9py8hGvY8F/+uCSZ8LhzuxS8orl3/dzL3zcE04dlpnpZuZT++qNdbhNbeI
jWpXT0Cvkr0mkcJH5sH+VMwz+rPXS9UH4HcjIYIpTGhK2ANVUsufLfPIA4O4uVFa
W0HVQx40HBD2Oy4YY7vRFM8w/gKi7zsJFaszlubPjEPdiaIKOmA0shF/zyxrllWh
FlNUnv7ugZ9vqVUQKeZ09mQWXseeZZIQnie1iRRVywX2z3EE/L+kQ7DS7sWK6852
isB4gKfe8/aiiJv144RK4xUblactM96zLSefDCMKPaG224YWwnG0PYtjIesOYanX
qZMyluOL5YE2+Oct3AjE/34DHlCN2fSOf+yBVSi05GrZOrFW/CqVKxa3igSeuKZV
WmQtCjFUE+zbR/y9fgEidKt4cyglsKzhX+FOUSUcra2JUIq7671x0vXL2jx169Ss
MlmYYubQqFM0Z2a0hVGkq7nSyMIbLNkhpSSpOymGJ99A8CwaWkm3kbjcpm1XwY7P
6RJWZQa/EBUFHGwQxFp6VZGwpFRShHrYXR0RAR25vOt4AXaR8d2iWnRNgq9/h1Dl
7F668IRn3AkE+7tSiDmOWUWrMkXrdzb1teTaiSG0zRpgLepgCU80TeTxhsL4WqBo
kicoAsjPIpwniJ5yF/LTnJ5TR3DWrAWDjDTVR/iqHqbL8msf+z7YuoFkMaC69c9x
dRyRh+5zY+R6TnJ33gG7EydGvvIvb94jJSYRtQN2uid+QN/qhi2dxKXy+dRBCYQW
/8mvbFhM8e8OUl+mGml4fU6QGXQ39w/XD+zFdq39QNWW32rOqxX7q/dTwmxLE6h7
PjHmGapqbIdkFU/Jbm56fOjQawsT6Iovzq3J/5o0ATuJDAA6i08tQl7Ph/oP1k0T
BrAmIhDMZk4l5n3I2Q0mLZ+77CxuADZcsnPIkPRuJJi2FKxn2CS3sinlcbci7HxD
vf979E55hqAc6rZsZFewFVjk0oo6lNWdCgwM6RNs2Nb28jO/yva+lWJ1R3vu+RBe
DVCNJkr/ey5JqR4RqbEJ82XQVOe6YhIN70PRPY7HVOkPxmSkIeSH5Lw63ULSREuF
K/7VMrGLv84rRJD+HbyVWVGbK8vJsV2T7AfzowdsZG6KYaJ7DdLqdVdjxYNIsVo3
ZgJabTTo6PtI9aYg1YT2mDr8mmavhQCpPfhzEb5zAz+6CIFoajkUEhg3Dpg3K6yA
7y454ckT8VazXrqtUcdKZOqT7wFm7FLugPl6ifnq9hK8aY4Cr/XOccHUnDTjBaPb
Be+s9x0yM+hRdRnyfEjMVHrFS45Xh8m5X6mIPdE4WHHbYzjEnEJ2NQcGNXOWi4qR
7NUfVUabRd2qV5jV44IS5hF47ezV0KfHRO2+NcxK/JE5LHjrAcvkA/TjGKPGrhEi
Ylznbe1aEwRi4MnM9VdEJ+TmXa2EH42A/VtVG95Mv3ypmCk4mTjLhcIIgBKsJNKJ
Rman+fbHftws620+vsnwQce3qrSMj/3fRaWC6UHNfeuGoh2uj2uZyBnNSVPwP92Q
GMEldlr3EVjxV9crtNu9aksQqW6vxLvmXrH0xVM/huyYdCfBM5E55Ywd287rWQd8
jl7al6jlzPUO8jbHsiS6/eDuWSnJ2Iah1zV0ZwxxuMJr7XVIl3TiGN95HrtYwXKd
Z0Xro1KDSfTkzy6Q+jiAeR62cqIC2dobyyO6wmuz3+bgcZRK77kUzQ2Q31G5E8oU
sgibTLZedN7p6QMpQC0400PG2Cl7tsfkotrKcm8j/HMhpqlGrnMbbWjF2r47qYWM
+UPFYq3rNahMZ6S97ME4uod2BAvyyqxXmgU+0Hh9E/KyqTU8Sm9jYrrGE0XV4683
arsJQ3Zyv52YO3U4f/4PwS1VejlK27C4KEsQfN7F+n6jjHIXP83/UQLjUMVbP8lc
4lHbLlWyFUhpN3XshwgtbgYdmK6wJyBVuBFPPrvAQ6r3cMPqFcuz2DLT+Rle2m2O
cfyVQ2xFHkSAjOPy72/bAiRDK6MiTenkqOg8e9iXNqfNBH+ot8dtwjwoqC5sYoth
NQXnKTfbjUdRIc2p1rfoQhCpdArb11/KUV2LuyPwevcTr1hGtC4CeFgR49iH6D1J
VWJOSvhjOc4ZggY80It3ikDmJohdIPPD81doTkO9RTl58lCiP2OA/GKHaZoYcgSi
zuBF3khswRyqmhHS4pLDI7d2wGrfm9fAH5eO9My7gYN8kx5zWAD4ocMfgY8pnp+3
rmnTdbYr2avnMTdgQbCxOyzsXM7kCIjnyK1lAOuN3/krv7a1pdetr+xLJqCuDnMa
xnv9bpspYFMG21GhEbv0oQulxVbJCXAqCLHgIj1enMcQbgUPtLsuHvJHZ7afd3ai
dZlkd/fyNLE5PHBP9df9Reh7tzb9jiUNnmX5MkJTC4WzgKkYkYdCqGW/OYJEAJN9
lcFH6fBw/IvYFq/QTOdl7ZPqkAkWnaXs8gi1coCfJDbtspOtRlMLXGjnY4+LmvCE
jtl6vQOhbGQIRoYsXXYi2EOUYWhdWbPVhIRKN4sUmoWMgyhor6T4+5zEAPKhlKJH
`protect END_PROTECTED
