`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9nH5vvsBY93o9jJzBgBqCzl6epFPGcp/buYmbPEXIUaJ1sDSdW6ylChvYGSCs0P
2Wu/aZ7cHb6TRkcvCIPiJHrhO37itXZb4tT7YWEwUtpppR6mIf0K1OJqircTMeew
S5+5ans/3SDzBOe0rEgBNJ5BrAcx8wUPfYXbe5PVBwHo38ILNLuSlUx+/IVaz4/z
HEH/IsZJHXTqkwpb8S3UBsxg4EHiqr7ah+G1H7OXbo1GHdsAXLzQvDX2M81NLXYv
ed5xD/wStLKuJMi6yqIV0+TJX3Fg9uc9+8udujo96XC30Ki0mP1T0YzQB77GVQ+z
6FtFOWO/4maJYrlN1HM9CDvmsML96Ttzpgb16MHcnkjxtag30GdLFzPNuqzBi6UD
97sOZMOnIEpVW9byL08nsm0Xy9Cr66KRQBSRhsnzz/a4dBVnlBO9N/iP7+iPZZX1
h1MAV3FYgn+b62jTzjwN7mNCJwlm8hwQwPVB8kofLmkimNUcQc9th3w4IPTjvLQE
`protect END_PROTECTED
