`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7V9ClN/lGIRm6ocTRAZgN1pT3H0dN5joADQknyh0Oe8LHnHvjavWovs9Ls63wCOm
k8E/vIPV4WsjGDfHRCXEPyOyGQoBA68rtw+UCvK9Vuec7KsH8hoxYqIRpf6993b1
TzHXgtyCzweB2fJRHSJ+Jm3RlXhayj0pW5sEOP7AcKVqdDeLXMaH7ECH79cWvQBh
cBlGh29UY8y4ydu8VglkJTgetnSXthSgGefcVWI7HAl2cCFkWFjf8jvDdw9y+m8l
Nk/zn1GlJeVDPwmC6mulJPM/en3vmJxKGtd6wswZRFyBPvGjo4bzyTPrGDFCfee9
LMg0CR4i+fBCMXi5jp4foRrXGWK5MXqgmXGkRcjKnBZ4cSV4sR9gNQYeQt4htouT
wbOaoXwtR1R+Y2bEf9+MkyETmHDhZ/GZ0iAhxTeOMVkH9Niadk6wefnN+q7Trt85
3qlGv8Yp14CeSsaOhbivqI3hWA+erneUcacgg3LPL0Qq6zO+F3zD8pECWfca2Ao6
fZi/gjXW0YQDBT9bVwDnjZIIO5cfq3OIeGlQ1vz5pV+ldFSSZQcBqqPvNwr7W/C2
CKntt0Pk7NbLpXWGsx7f/eaCbr2VSbGelPFJlUJpatSPyw661N6+tAuo/NOmomjM
5C7tEfMOOWQ4KnvTbuA2N7h7jqp5Q+jpU5+cTBn59nVOhnlgflJq6eZhTadquIAe
hb1m/NaeUOSYLkKJ73SEwQN3pvTj3ucPP8A8PT8Z06kHiQrA++VKlZ7FIUyKsTnV
uF5y0XVYp+N62KdwXizgqOqIJVN73XSVGb68nTp1kBFVjwkJA7TPvp+M0AsC5DYj
Bo9ptT5L+Ke1nigiiy19XCkGNnQy0fHm2tePhlQrQ84GHVHv98ET1dFiGv5kdWKw
`protect END_PROTECTED
