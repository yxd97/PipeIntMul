`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b3dI0K15VH4L8tf1vPp1OSdT8fAJy5okYjIGwPPSX8En8VUdMYy3MsnB7A0d4WRT
SKAFrVOZdXQlTmr0+ZHEm7uD6pOcVa90cbK+avu18c7It6w/H8WKJ7Q5o//GlcE6
S2MFDa+BKxVEydL4cXOiyfHk3A6g8spUZ2Iv9z0Tg/uV79LCJd3I38R/3134dEas
twu58N7GI4TjeeCHs09x/0WNd1rkvyQhPtZDRjHjGJEIinAoa4lAXalw0yIuyv2T
hdsD/HCia5PCQm9sHTGMYfxaHblpn3YHghZBqCkAgBvtDMXaF7qDXq8IEj6vqFJM
yNPIzhseECy/YFk2Zt17LQwRnFxZSSMiCEYV+1cJfv1KmB+IAnm6EYXD2IXF+8Yh
OSA31vyWJSvztK3SIKf3BEaRTU+kINM6a5HXyA26naAHXNchHqAOU9zGHlhemm5c
`protect END_PROTECTED
