`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNdBYkEQS5QNAvNJhS3vCPdNJ5s0WF3bMfJGN7AsYcVMidkMeIpj/LKmUKsgzR/8
VnDvbTBms+3i4W5+LWUDndgCZvoHD4sziYrcrdNpZjFK4kpMuNJYbOKK1eHOpHeB
MqfEp7dlTzv0T6KfjZpsLWXKxuBiYfDKbqmL1hmqRs7cyddeuT7Dbk74KAYw6uIk
5CIDD04L/47eGoALjYDoq/0tV5DKzxJLNUPxgM1NqJUU+7BPQa3ktBzYQ9xmnsT6
gdXMBs4ITn3OE1ubdogfFjB/srZpYYy6OKcUkEZkxBOHvRx+y17MZLPLU5YE+Sv+
qGnlBkM5g5Rv47VMksjtHpLcfP4HZ8V+Y37i9GO7haoU45Y+C5QNxnXCKtVhtBZn
zk12D0OZ8ZWYbVnk8hRuXYakihhW0CCDBcRYssyaZvVoTxjHLc58iBlkkir42dF/
pzxNkkH3ZHEDS6xhvVuiBlx48Kdnoi9LEK2of5ZfobEFC/A0QHmjxxmjqKYHRAjH
BhRRuevKacuR+4ZcuXoutqcp/wtbQM2Eub+J/7Z6tnWNZYqiFhuuGMOVwDAuVZCa
jnVimLkLeFHfvb5JW8nJ6kj6Q+hmQUlIjCfSvtrAXfHWT708mI15Rs2v2/WTsecQ
uATg29lk/vhj+Zjp9+LNWc/RJSfBtojbGB34DJEoXC0=
`protect END_PROTECTED
