`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
auVNGlZuHGcFUboOe7ZqajoEQ33BbJUpEWpureCg4TZvBGiqUJ9hr4sr6SPYk0Hu
dmCPf/DleCsUvMtRZSNs8sryBroPswaPpYvM7mCiuBhfeiDle0OvGTFkOE5q0XYP
3vHsGPZqbmg56Aj4qUNFQt96L6OFr2Q1YNa4Vcd/tWvULzjW31JlN/2c2Z+VUOWq
crUHNUsEoCqFZYnmXyG5ar480xxfHuRqxjyOLffqVcrNPThYi60hVezWuWOkEN0y
8chqr8g2XA8NXyV3W+OIXaB3EpSr6wm0jt6zChsx5OqW/uvhFQ3pEjhKvwgUgdTe
GMazID/b6LK1lpyOjFJzzzbKfzGgjeN1QcbPeYzZEduzVxttWwPTuJSj4JCAGNY4
l4l5wn/Lv1zZ2cfSlLB7FPi0aU3ERm3OlMHetZJGpt+At+lbgjMR90SvHzOHbzBv
Bzbc2mUdyK8zEVRPsMvbIzTM9wikDkXoUdCOxF4wHZ7mpAJ0OCpnEgCeQv12ZR4i
0fBZCRL5E/8M3Huypfpt49W3F1c26r9X8sxmD5Am2VpIgz5oqrs6opyX9kkcdLcg
bXFcNEW+mLoTQHZ79RU5Vp/xv9L0459h8QpX8N3aRTa8ZlZX9U6j+HHhZ2qlPvOI
39+esVfxwzNXwu3oGVaEFg==
`protect END_PROTECTED
