`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2HClAnfqcuIi4rqsSB/g9uL22dvxz0fzlLKSD01ncQLeHy6LonhWTvMPAM4gxU3Q
0v7UlWWVPfGD7fQPHLBkYP/HjZuMxU7EmsEpMiWKxhDLDXEozC2milhqghUf5730
mUjykDK5pzc5EOQpAoG//3O7Gp6oMGkWPR4nH4oOe62ZicbvP/oshY93P0ge8Edt
wJUbsbsqK/ny3oCaZT0ZORSrWWqw4qVZwfu5zOw5+cr6mEKxu8zbXrL+O91psnAD
mhx3H4wUQiIXZpLRcpBNI745OGerUDNqqHWx5m7aNfpewd7+uFZVVNhGpz/wETbj
UUJBDWpPJtyZjA5S2BdQALmugaye1A4xXymlqgw/Y5E1cytKjocOeZ9/jzrQCyMW
j2yNR+25I+NqJwlFOKGb2Y22qqqBVK0PBQcnLzzPebY=
`protect END_PROTECTED
