`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O+HJgEMtSqsxmk/i0fQDUv4kKHjmjt7qBZ8ZzhzJWg0otMQ5kJzQyVKKKnd1Ru3E
Gt1Z2Axd2XZJEVsD4QOPS/3dIeTSIHSlAV2heYNjEyd+w9iu0wsIdTxBYP2+OSxB
huRwxmDLhyKxbsjyIfOwDgT0RSPt4yxi7BiB3LIj740DNpxFeyloIhH5mr1OTxTr
jw4XDcuRPKNvMruusUb7dma4QKvGSL2j9Qa8b24zWNVF6nOMVEMK/f+ijeGbCvob
ENqeESOSGbFE9ta3Xns2IE8f8MhSjokeARasNBQuHLcFqAGCNV2eV/OVfPceZe/A
IfxVmLLE/B0MJCQul2RZlNl2n0XP7+sWyiOE3/pE+1DtB4J/kS+XbR4lCI0AzxUJ
WXaPLNObhOgp7nrkhcAA/wFfk+pFJ9RZlLWPCCanjquAlD3YWsvGStIpCV2t5KVa
yYQ1bU3fVGWc9by+YgkLfXIK4YQG8p9nP+4jyYwFi8FqZjtTXvdsbxQxnxCoO8wx
qG0bDD1ebWuv576sKFSWNabWTQa+EF6SCjVGTmWns4SNYs3F+5oDBP8HRrbAqpeF
`protect END_PROTECTED
