`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ko/EjhRhHbSXju0yeexzF6OfwD70CpaWMS3vmWCUmB4UU6MAOPIwgJ5Y9KiZD9sO
VEql4Ev6qamw22o6hSbTR0aYJsSPKs0B4xO7bJIzid7h+7FWZw+Nx//Z7bTV9qi3
EW0IWuaeMOmd5k/l5ikiheqAPo7SDJW2fISbzCldrUqzj9f2OChZK56KmESWEJIe
gSAYNf5DvoDuDGGzGtayuLnlGgODOLeo4ZERQOvpyM0IO0ZFXgCyi9LkDc0EcJXw
gaXSQJzDDJWa9nuXvy7e2PO3DmnTvPoYje2Cqlg708fnlE7CmbBlKCwxb/ha1PHB
RWuOCTLo+t+GXoZwEcnHotPYZkVnNhe5Teu+AG/OO9HYgEb9jqsFI42xjixk5eGy
MeV9NzSIujEcFIkfsCu1OQ==
`protect END_PROTECTED
