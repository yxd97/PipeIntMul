`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kI3bKmAUqUqqfNW6XsrwrP3W+OCsgtoIlI42nkoqwbyPu9G2tPNHKeUJHgbhHGC7
S0KoB68jjaTRSyAR0/BzE+1IN98HFP/cDDXflhJJ0T/oHsO09qMU3McIlDGmqRra
9Td1hB1Cvhm7qC/l5bdflY6YNM5KZB1VqMV731p72zE6Lnw7LUHo1bONYFBAGY32
Cg02CfRCFw/A99AptOW3rP1t4A9cj0rFzYmrhy63Oq56aahblqsQCqYhkG1HpcBd
k+mVdqL1S7zPlpGTFGOXXz3iNmtvVOdOPQjoWI/gMEpuPzLM8nOBJZeht+PUR9UZ
wM5gW5+sW2eA+x9X1rLGOvD18MXXIGzehCtfPll27v7rE+vKHLeW45V+3zBF9qCn
MLphiBCixEu2MxRCAl3PsWq7dsh4cYAnm7n10CRUM0M=
`protect END_PROTECTED
