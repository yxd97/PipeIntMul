`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tua/UHM/exq2OKbabQuyUvJW2uI6r2Ll2XDTjPgjya91wrADnS+rDNNiaxPzdmEU
GfmwSYXjC17ZP9uS+NG2bFyJaEeiy+r/nGCc2hoQHdtMaunRqe4pN9KjXMtnkUUp
R65UAGYrc33L3eZOQaiKh74dWkD2+ShR7Vu81MiOLJNnY0In9+xF6l5dnoCwSCZj
OBrWEZuBu4zdjea+jbLCPrHev9o2e7x3rBsr96X9zX/vf82MaJ9arJZblbNRJjRT
r6yp0M1EvKKS1DZsnUZp4zrm54yV1iOTZCjq67cSwNOH2SflJUVWVQGcoCkwhAAx
Vgufz6+gj7cciCY/ZiwB0q1n/md3HNrH2ibi+RMcSOrRYEg/jIn2wi1te3AwGFHK
C7yA8EwrmUduFClA1cIUl+nNgx40FZhpIEPHCIr6kVIKs4IP5fkaJ8ZHDHNn/7Ux
YjUoXHosXXo1JOZv+QPLHf4Id+fYpkYk3hEeF+QIuhWUjT3OseRLkPTvDhLT4JlH
si8IEjoo6VghjoBwiF/1OCqM5Mw6+tgUITgA7/okX9JsBZzsc0eidJ+qw/uWvPk2
Z03PjuuTtrmQ8kmEW7wMcA==
`protect END_PROTECTED
