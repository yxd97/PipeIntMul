`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3yD1fYhMMLsCyHII827kZBvEMOQAbtE/S5bI/FVU3iDAJfPIZl/TAtDhOYcmeKUp
COmtPv7R8tF/B9enPKya16k8ypmBLi4RWreGRZuD0/SIz0o+XM9F63x2x+5txCHK
lxVyqagjzS5MetpoMLmh8MQFhdUz4kigUZXoBU16HiLMfd8znLcRXqIeTOTFTYS6
QAhzzSC6YD7qxVZHChXDBvTfyXiO4YKtqNsva9npQlCFimqk/uwPoQM8MI4d6AK4
WQmvqmKY8wi+Cv9ZzQLx6xsXg7lXdu4ORLOdjdWTK/e1FkOeBH3qmc4iDk2rJ4gz
vhvS5eT9PpSIDF7OYIvHjSBcWpILT+4hB34uvF4zy/Ohd5IrmTVZgfjTNgCCChOG
zSf0lAf5hsz8wh67Xtp7CTe5Eo/UaFk4PgFs74wIaaYerj2/D/30WfY9Azbzg4Dx
35MUUTDG4MOViyj/9ZSl5DDLHZUJYlaP3NSxAicI4mgYtpMXseFYgFBXC0nNIR7A
P0f8G1xpuTz0Q6fI23fSTv43TLE8m3r+EcrqKK+6AiUqnLyhfq+CdxYWyOm+UJfX
ikNgiZdH7OvYH4icOPD3k0p5ppd9xamFcxUKw/wIxtx1dNhN/GlyeDkmKNlNI+II
JehR7d+r648je13RnP32WMZhjJAQCQY74/eg9+MxPeTNXrnupM33Qs+wB+bNTGPJ
qczIebz1bE0lPp79uV/Tys460c6pSE29Ypt5J6nbthWDrQHJRqj5+R+sxJC70ycx
xOcYenw6606anaEJnObhACa02vImiP7OwKn8+WSZD9RSnvG4Y/ppFLEsvenbZfGN
STkuvA6cMIX+aWabPk//64RSPqc9gjfCKlFiZTv8+HXZaHlUeoBEvZzxb9EUpfEN
c8MsqUEW6oyqshB3vlii2Q==
`protect END_PROTECTED
