`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dDWuHK3f8RI3U4juvWN3qcBOa8G2gR06KKnBMgmPqTZdmYZLV8IZOZYkxug2CofV
SftDob/0zz3k4vYCMUtrQe1tdRYbUGwMXISGVMnm+y4hXcB3QJ1B3D/sS4OSTlcx
FChZvTvlJZnuhucG3VTiGDID+0S05GgqVSoxnvwexERZs/ZGG9t58esh2Xn0RsR0
D/ls2WdnHzj8TFRXBnXxfcg8nMlwLTjJ/lnJr+2PrcZVTsRjXvZJdBvJ++EgyxRt
UdgEkqU/lfGKg3JzogWTA7jHKu5s8+IsoHqMRRsjyJVYMdYGQnOUu0PFcdjVvzAa
68PwzRpDDM9HA7A7jv249W3TWpEF4VuiUaQ5sOodANKnODdd2Js87JIPFnL99fmn
fzJe14ZAZ8WQOh9jvb68dZws1rRfBWG+0qi/Sn2kLS0=
`protect END_PROTECTED
