`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P4u+0pd4w8s19kqkDeW5Qph3J/dt/T7/iFN5ScpBkZqTyMGLXPPJiDxLwXgBfuR3
65qZtqmbmBdBSYKlcgelOUMfnRGcfxwcDUKKyhvRR1tAtzJEZX4c5b31HwFYDn7N
6zmqm8FrgvbcjyGHMGR6bqaVaNzGXwSOPV1vsanoEwE8ecamTiSV3cPcYAclc+FN
+zrYn25aQ8oNwF/7bPNjm0S/Ro6yy5I+9xOMXGEYJN7D/RmT899ycgUKL42y8qRx
osCTbZY2IQqI8QLMdAKzHZrkFUwT1u88ciBeCIwTtqk=
`protect END_PROTECTED
