`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfl/0Jbeyq2gJW4eHflO3Wxc+3KSqoSca+xAWC3ZGocxcJfId38UKats9KMOBYPn
StojdSZa8W3LrgdVibh+okxRHAW4+69hxOHMxElas2kbiFLkDiPpdj0QR+aMNHr5
oMqcRUbKiJ8xhdh9WVGeaaSXc3iu3uxK0kdZy+qs/CYToGQtcfZ66YOcktwy2UAl
hkl67MwaCWM623QENBp+aejiEAuukbKmXNaNSqRe/dHdkjR5b3AqrIpQwqqa1cju
EWVX8BjABCLWR3XlMcDFK2Icx1YXXK47g2AKoLHtBgKvGpyDpxyTI6e1ZsmlESaq
+7NloVDxarlBQsNPBpv+0sIkfTjwobHFmZ38nVsmgXOBg7IIRQWTD9xwalIvDHoA
AXpCQIf7XUy6ncFLFWPE2A==
`protect END_PROTECTED
