`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmaWsDgNJINw5ULyneDQkre7M7TqXQ2MLIAa0SIapskUEnnU5dUoBMgGanRQt6Cl
g2oe/dvl2xwy52hSDzHgeEQlkRmFxjK/0ta9aJUteOfVa06y1sxJW4PW+6loLgXR
kXHGmyenU5EsYOVu7zBOxzVq9f87jo7YbrL8/wTXmS8FVmzqrhr1GcVHkL6KjQFv
X4cv1DK9Lsj7Hjpfko9PhRHHR6E3DDlLQyCkMW+9jIyDsLKQP99ePu3HYPTzm60j
Ee8bntuVNPpzz5U49pROLNON4sMGpD0vwyiEMm02d0YF84h6VCmD3tmMKj5PHGNR
39ONhJQzXvC8ry3opBr5KVHyxoVEhsY7yn7opD77oo86Q67Y+Xw492g3Y0mXmTae
6/ZiD2dcl7Uy4qCWUwJelWckvRHD05jGZ69y2yjf3jLhfDhxmO3n3KXj3PIJiKad
8LZqo9dUW8GodWtLyeiXKpAP+EtwDIQETaxBf2H84ajjvAZ0EhvgZVIup5tYrhR3
VWU240uXF8neIfkdYA5WA4K32G0u5htPknE3LJeSKd/EBGHttDyVNHnkA6Q3N/0m
n4CimgfY8tbU3kOTYvKzmwIdaQTRLg0fcIybPIGul25lAQ2pHT8wxlsNnFtx2bJL
W1YJ5s44W802RAq2LUzBU30tq5qfug9BXfTILPF86zDLVUsKyrTEtMGDdeSn6os9
ZXYYkjYjg1CXlUtWxyVBJwwDvHPL4iprMB5J/ttCtgw=
`protect END_PROTECTED
