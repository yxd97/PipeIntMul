`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BtOUx8I5JSuq048oINyjMa52rRB1B+sTWP32GD6UAhyqlM3QIMhkfbqPq17ZO4HK
Objl2JRpLKiP8bq5gYTV3zXjojd+8/Rj9teWTl7hmvzOxn2TUOeZmV4raM2L0TL7
UMI6uW4xbDSx0kSSpuTnP3VVilyYysXyxeqJOwFOuG/h1gsAGIS9+ZDukURyqzP3
nrbvmmCmUVYB/qMwz8UaSaRAaPqZ3MwRCH8UT0oXAg9xFaWK7T6zEckRFWPkvlQT
oB12FPZTG9dt4yotHanb2aImyOKd4YnWFqZiQydWPHVIgl2H+WtWeNj9+Nv4Xl/z
1ayv2oQIoq+TQUiUmlWbRRhfTzzrcCJMt39HqnfaXJFWpVwDwG36Yj4YHfYV7Ye3
wrVdauAdtu3gGvxXbiuJRNE6aWGKl8DN/s7sU+wAGWfsI/mO2Na2k8TClPpPr+EN
uM5U80+qxwUYYcZPsiDA31FTPzJz8MB9eYAeaoDKNa9nXVeFyQ8DY5c931NE1/aF
KVl9Nes7vetzv+Iq0xZkLFWktd1oPwFv/bmI/rbrev3NvaBxpmVJ8Y+t2KT6n+/s
NYjCqDpicXWblNV+6kh7Q3JA5tOftk3vnELRLqJ7SYk=
`protect END_PROTECTED
