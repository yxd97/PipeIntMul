`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZSZPVDT1MZxrwwCe5OTqh6wxynO+wwmKxB1w6dZoIvrxKDZqmnBSiKwWzkRM6Zj
6VbPdb+q/LPBc1DBytvUf/tGNDseywu9iexDNxG0ZNiApVKygPiPiGVtgnAdOr0b
1kOn/+P+iaB/Lwy8rMUChpONHVWqIeFO4OG5z84OIubAReo60G6z70UqE4E05jLi
qlR9T/EBoKEWrRkrdzIzKllZnafS54xI8AhEhfzs3bc9QYMpMNUjijAns7cKwDjF
xUWjZmn4Cts9BfuIsLKJKaCHJprhbf2YV82P+L+FzImWS07fCBwygI0CvyGZgtPV
ieixOJYB85YimoHE7+sXNS1IaY5p4kKRvZfRJj3FBd4Kuib9UMRcEf+FOABgtRd7
AULldeQleFXetPuL5DWwxBWyea6svr9lsHYliz99ytObjmmhZL38ASbHhS7FrQ+E
Tv0dnhlUBRJt1Rg5V9MtAh0z1vDO8yDXH5ZXaljxn/s+Ahdkrsj3NkrzT9n+XZ7j
4hneeCYPty3uHR+6NLi8A8ub3cmdz9K8tAZJ1ituLvG754blY9ZEFJTM53K4Hh41
RReGVwRzuQCKNsXjiNz7JnhbrvFpEgWh0B0KxzHCCOU=
`protect END_PROTECTED
