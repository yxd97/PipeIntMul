`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cu6Ytnh5bFJF7G4+hjIuI7wJLZk2rwEF2EAK+tEzk4+mp2xSOphaqq2ruCHAH3Xl
lyjiNnu3lbEuSmzSsxKNG1UTgUA6et+F3me+y57Jt13K7N24iRbgYw8qy7sfqjFL
iH6CiTJzT96SHqngZBy0smut2QVd56Eq/UjROa3sHxXBYWVkFZYZn77QMMQMTsPT
bBnOJGRmPUm0qT/xtZh+RYnRJNdWuYOXmSdOaVdQL5IpXiUYOwHI6mVK8PYVvzeq
yDszS+fbHftqBhDt3KTRl4qEZtm8NlIs6ASK5UxP0wqf624vnj5ZOvDpnQeEL+Cx
zI/SIwUPq679G9DGkSZjSrsLV5Ci4MkBtVeFkPt1QpS1xTWfsdAsubv5NG9WAqnt
hAEUY49wZ5MR3DB+dBMqduE24C99V9xVTADMRDKP0UqTa1b5fOxfrXplGKB9+lrb
`protect END_PROTECTED
