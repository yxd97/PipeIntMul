`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCt9AwTXqn5vLJdDxe1YewsDgBB84ZVbcpXohvO4kGKHljfl++xoUsIxT10DN6uD
VprJBRxIC0nYvnBJ70pW0TN28BLW2iMO28aNwOptM1qBi9wgk/aadgAPIncs4ONq
ILoQmP01S+hUmWAIwTj3BLZTttx5FiZVmYRgS1zjq4bMo4fd7y2A47HH1fHxKVQs
ReTvoFOrdtzrBJ6TjuXfjm15tQ97SalF2cXjbrVjsjOCDNlhQtPxlxvkFqfwEm0i
lZGS2mAF/mJrT7FhRpehXw==
`protect END_PROTECTED
