`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpZxBgs/l+tZO2l13aeSGehnJ6XAuVaCwlFreGacit3yRAOqt6Gl2SEQlI8Ml64i
7AEuhqHf5Pk8zg+/GEvaA+fn7HZnFU3huURcXGjVfPfBoiZRP2+DkJNKDJnbX1Y6
IQm1/AIMVuOxx+ijv8ee5Z3vJGCSjSkEMZ82cOoXurkOH535TfMeZRerXjSdU1jq
qQvh88ekvNkdACCkfEwAYuZOUryf9j1ZjZihHXIWM7qy/HLyPnLottyemuAs6o+R
btfnPKCE+4ZDLWhezfzyCzci3qII5dz8xobA8vikILxbZ98UlGDkwQ91fe3fp1+Q
m8fDZ3Hb3rmUU8/ER4N/diH90kNJPqFhEWBcDGFzgu9AwPh3lnAz+FwjX6pPgYx8
mksobGYUgZ5vT0clU+z78ppRpaMdthldGNSNCFe9I2OD2MWALbKKFbFq09VMI79A
NVGEWzV3OsBCDWrxe3T7thkKt4O0AzrG4orvtHeGFTqEKRV6wSo1ExuIGYWKrZ2q
9kF66sikDAv7L3wZZJyiiIOaOdb2NyULp0aXUSrYVdjkXqksEzQsE+fm2w+3kpR6
YF3sv9jV8oQB58FvjNn6aKWfHtQpEgfY5iki90ilN0bHW1Cm5KL+Uf895ZF2rmpe
il0so5r+xa1g53T2HPKuEYJtIKDJ1VuAqR3JhSnuUnVqA+2aBSBgZYAAxMvXYug9
AG44CAQul2pNMc+hdWKNam63iW11xq61rTFgkPRb1758DIQTEW6cYOMQj0fDQrmX
5RcWwvJU6ofQXysDuovAQC8uDvVUCcIdSnx4WtxqUNxPSkCVn76rlb0VebU057Jc
7zfUEm7sdg+YDKZkJpzG0ITD2R8OYFK8bEutcyKPy5jH1UNedDC7+zD7Sit3fyL2
yPVe11Uqx1qDFEuJINHYCIEwv4asQ0c5oqdNQVu+PAPDLrvk1Egg5fL68kNKV7va
oxxAYuoAZOZjWF7OPUVe4QCkC+lAIpkLPFVYvXkSn8c8HK432mJzN4URuXfIit6c
xuFL9bUpiOvxNA7Xun5MC7M5J1mzo+4fDR3YSQzSl4G0CtetP0vsfgBxaIkNNTX4
HOTiGm2XwvzuVy9RAZOwG+E73v9GKtFzZTi6h+4gwmw4ePmfocx6RdZ/4pi5slRN
snncxj9CejQx4NtM24EaS1JoJmHESxzQF+YqF3HcOTg6qzQkUfh9MLrxRivKo3dz
vFwp2t4B7SPEkjKXrobpV6RWZ7U/N3zxgHosgU7KaMZ9QVpJqROSApX/9QiCfuTx
8Kz01vV0vvPM7HGmla6pJkvHEsl7XkCbyIZnZ2eSLya80rex78ez4UOU699hjdHW
6F7xH39X0vbSuMFwTNcFspPK7Id+MExH5rQbKohkkTxREJ43zf7+fGtQMzNDXFnd
FzSc5L00imaobh89HYpIRA==
`protect END_PROTECTED
