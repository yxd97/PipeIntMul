`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wcLSrnHF943VOfkhSmyd/arnPyKbEpJN7j9HRcWjX5eoYqAwn3i7ndEWR3QeXbR/
sjMXnSB9XbHDR7zYN//xvsknI9ndxvC5HT9CoetaZghNBFsp9hT+8fauIdS2QL67
SeS3oO+/2L1I8dqsuE/2O/FPJn4gt9cp9DBdg93HKh7oCXD+Yx+W6sRKzaHZS2MH
AOqNZHZu+TYLpsMev6nvOW2y2GqDWBs2CsgILmCxwKJpT0MgTtB+iU/MLDlthC1s
bPhQ2vtYD+FZwPifWbrTEQ==
`protect END_PROTECTED
