`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eINOno2dfPcrW6IXMtqhETRA34DdPhvAM4tJrytnf2cyfHZl/Ah8WOYkUpEbo17r
KX+hKOeJIqdE/H+Ptrr/2RuZF1nfpokenXWMuut77Wrk1M43yaUDmp/R1VfK11Dn
wO88AVLqWMceMPZARfVWB7bnJWN79DY/k/FyBRCCYQhlCj+w82UUZMl7CG+JiIoh
wLjZv77NGqjltx5xWO0SJpru5/m/w7+Em1gNorcD4jZx62Tjp+wa9XpjepPvpWNJ
AH0FzRnoswEZoVAOOin9YlXns6Req6rA3mo0BJI3I7+bv3405qHAcN4ISUjRWOap
bQzoyaaVASHiQYItX3F6PMU87oxwEGO3ixPeZDWkP62Zy0rSTHAeLjqHVbm85XH/
2k/JfkvILQTYxlCsPgZWvIPPq8HERI+tqJO6/I3KqyE0Dyd/oDxNaNwz5L3eUQPs
vpVhk2tKLKPo7DEuCgmg8yP8bXyXUM7kyAd8XspeyAOfIbP8fjD3mFMzNUg/UgS8
V3B9JuP8r28r9NmenfxTm7ek2fIce9k92H44caKdtq/+QfGtlGrw5YHXeXze+6tB
aiXTrPfSWitG4/7t0dsTlk8Z7aGCxCx3M+A20eaBJiYIjXqPJKuuFHqwJ78bM/G0
MMq3KkI6BraOiL/LIxzv3HgNg28D3wib3pnKc6/+c17MIwmCFLpu+5KLlOVRKI0O
dHzcuClas7AQys0swy4N1pMztDfNIQezg8PwqVBJK1NEsfuYPHwnSr9hyhpmz/8V
KtwaVlAJBbD/VTy3MyMbPEgzqu2YotRjHu7mE9B5P2eEMSVX+/kFCaP9hbv4xhcB
a+BY8Si0+nPUlnqiHyEvc88q0AJxmDTU7YJf+V1h1R8BbnilsQv1ZxJ0SlUcJwOR
ExhBA7YRva7+UBTdymbHBRg7WrGiHP+xI/AFFJbwlsqy14M8FxmXN7IqdH4Y8qRC
vVmUqch6umJlxQdbUIfQDBFf5+bqA6jIdNVOnjAu71KrjLADhSpqdEPWRhhGvyMn
xQU/X2TByk9GBglGb8EMkIb0URF+oSWpB+ouwsOaNZ5S2no2cKyJVMyj52Rsb871
hH4fvt3aD8R0nypdshM3TnvWm3XuPpuHGguKiKWf/irbr5BM592Ditrn+nUtkQPR
aPClkKjQWqUE/4fHOs496vfw3JR2KFqICjyhQT1AT7YJdCrYsfpABiONCWQPHons
I3sCDcQvTTRA5fRw6NqeW+Lw3Y2eShG/YoZ/Nx+eTXI=
`protect END_PROTECTED
