`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
au+/3wdtD+GPhFs345HgDOw65neSQTEj7sOqiiNqQTa01VGECkbAb6uqDOs61A3e
01R83uh6CmPKH6ANRaoTgFVwdqk//HXeTf6teCUTJiDSF7DeAgoc23fTTq+c3KCn
nntTv0EPi2n/H6Rxpz0UaITLs8Xdo5TwCaNu/o913lg+npfRzweMg3H8DvWvxXUc
L9EYaHsyLLPX8stzkzDmZ/1XlxhQyRXrLIMZzTH5g3g5yHdxm1g02R/SkH1Ddy+t
xoDD0NldKE+LAVQoc1BlQ5nhIWnTbK2AXwzjnCxWQghVovwcAI+Z2RcSP0t8N4Qw
tQaudQnMHvChueZqeoYFMNCBIpHihmQ5ZOGp2Sj/TmuLFoVhYvmq5RoZhm8Mm+sj
p0zUkztF9w835WiwINJZ4joXHwlddqcDLnhVqQYNbHCXOH6OcjnKIpRpQJhlgkvW
f4mm0/bcDtLetgodh/ywcLu70nq0WJ/Ojv0H6RJCzzQTHhh0Ok+LBu2vEeKHntH4
qj8083ZwMkhaQEooDNEU5FhX1pMEfUJfamgX8SHAECPpw2J7V6NOc2+UKlvfU5fb
n8nUvlUJECbHeFq9CrrNcm45Kmjg8LA3RjLzO9RfbEPnBcSeqNSfTrN2oQ9sS5PK
sGj48hA+T+YOXjevyo27Yt6xlVTMIkB8bFK9xUMM3tE37q0cb4XfXSC2pLmRNO0x
QkmfwwkIIQ6xHpBMKI1it7MDfCU0jFAQ0ciRtjThMnZNhHgw6Q409kIFBo6Nbeny
g7tZxYjyL/vbFWAxdk7BVKonbvjKrgsKsBz3rX9Nwf/NSggUnXkcjHjFb+WMy/iN
B7JVmcsld1Vn4jDLZNAWWl1IxMbG3xIbCJfCg8471MP5gdUcBVWYeX2ghwBHp1V/
LliPfUDBVy5WoMEKAlVgH/uwuYZQZ/V3ZL/aV55MN1A3YeCQADj6dcmn0z4T33tM
qCT3Momn7jgfX5yGoh2OZwTEe+7G1nxyx1b8AT9JYhxk1S6g0TnzjJP7hsd/vvpm
jpm1BL+nbg3dA3/+OLW7w3HLMPc6KtmkITG/q8DCxh5f25H4i95Rvfml5MMOwFtV
0+VINqgqgdUpvqM/uvD+j+qgl5n8z36HKJb2PAr7GkPSpZrrlQqtOgPCwg/AkdyW
D0LwXuUuw5zFfza8Jxbr9TIlVSD7AWAXwZMlVguik52vDXXvwdcwhH58yvL0Wb14
phOfmEjiHCTxFr7OKufE9hCsLQ7UpTdU/t3jP7gMGNMPMaJ41QV8hHnmKaUrN2p2
QrQkTtHhMbQ6AkjbsybxcZIrmtCcz/hoeIylN0MMuSZmCfA+GzYqyGLwAkU0snPM
VEvHISs3cg3mF2W665kQaXRRaiNjN4ZezbtJ/8YsMJp+V834MQH0EsHU18BKGq4w
Rf2l8dFiZX7LPyyvp75Pd5C5jgByvR4AtyoHKmOx+RgKDYqVEuptlBX+4bPh/tvx
yPTmguJ9omJmXir8LHE4arBZg7cSXKsQvp+irrEB7tk03PeH9IhPa+68+d6C4N3z
`protect END_PROTECTED
