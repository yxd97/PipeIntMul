`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qeRtBnoVDPWw+LSg0EXonXPmO8j3/iHvCDadH/gY7wKyBxPb6rLwnfB5yXKgdCin
ApweDHgZ07OIBySXF4e40FmH+E5CPxACIkxP7k7ux+cvaGLmTCHH0eVebU2YKQmI
RwjZHlTQHAPzdrSCem6y9wyPcBw2AT0TUaIzg0XBbMhI5mFbR9DwMlE2L9xCKMRx
55EIWTk50/im82tXfMso94dZMicsYVz6Vyg8NaF/4dbOc7IIi+E/NbJVLZZkZ7da
`protect END_PROTECTED
