`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRiPObkjRzu5tEDfnWwG8TT+9b+r4edTMvnV5i71Ipg9BW23VKIuWniHuF8QikeH
HEssnsTkgGc/HsciN87EKyUCmdXraNmfsJBP9f+LLvjmMl1Jue9qN9+XS1QflfVt
HJCQy6NI0YbyRCHutDAu3Wqwiy18uF6a1NSUCUN/zqnvRfMiVgv959AMuSnPnMio
gRT3tJENWh1BFcjSSwOUsbAJBJV7p0Azbr/JkH842bL69jmQivulwJsfDIY8k9ir
EynqUqFU3RlaCBmgnbMOa4iuDrestFSfMCrmXTjOIP9QeeXEGYZYZpb6L9Kuk8nY
x5YvmYnbdhQXmTUfZKHnWrXszSbII54niJeTeH9SZd2JMe7IA3hv6Ur8NwFiCHo6
jdysxtVQPySfwmslCh4IGSibJTF2J7HxaQRMYXxgivjr138L9pZuDowcI4+DT4ss
9VQrHPb2Rlhz7HuWHu3U9R5W0C7NGFBAUeWDRFOk/La0FmGD3EmxluDAPIITAfBb
gzWkVlWzcsjLRt/4u17j84lBvF5HQ6ioCAaP/Hus+cv1PmfYk4h+ztvhQwtzrj2A
kNrqcWdUOFFBHJrYXSHaIFdnzjtWAHEf/iFJUxq/FZ+XX84lzRnbQlCXehuvyomg
sBIfQrVTIBQQQSDAIZf9nAM5Q7cGfa4uHJjedfCrRaWNJyJ6yXGgWuXwqGzLeH4F
8NeUUqa6pSKpkwaBYOwDDEXlYmU0kn+2C/olZyZJ2I49UfgIVW6K56MOYH2KuU07
6hMgPZIgbxqiCoVwZTYb3t7TKS/D6rjL/7qkCQmv7S2Db7zgWTA4TrAhl5qHhBbS
srjLs9GqXuu5Gb5/jy4O3gZuiTIPp1KRFiJAdjBzu8kgghwlynWLGvRfHDWYYVGg
VhfEv0Go7vRXqb1GkpwzQEp4I8jKSjeEzVq67TRBDYiTCLKJnF4Jl+gzswIAGXD5
RiXcYamns6rkpdHV+VLTnlrThm8W/F3g5zrX3q4PV0ZqnYXUxFDFJfJLkfcMqaSI
KitJ0/Nu/u53CL+VURUSHP/I1wvGSl/+Wo5Bot1XzJ+QMqTothk/YZxIXILoxvuR
pdWsXeJI4Xjs1ZzT37zpxbiKUdpyl56XduqavswpZ9ULiAlmfeZkCmAmUqX81Y9y
z3/ng+RBUKC8g/kYmbG2w3wNXV1lCSx/s4OQKyy69El9ylMjGj8dx5NaaD2Ta5MZ
+f3nvnJTv8IzGFxNPig4bQ==
`protect END_PROTECTED
