`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ViJGj0zVdVdVg1C4tCFhqqJ9FtocAr+67XYMGlRe2P2P5WxJzR7iGZMsfyFLd5b8
6aJoVgBZFfGhC9HdJkA19T9cFvd2oEKoWkLHGKpDykohh4mBDb9sMjBiOPrLcea2
P+iviWVt77fY2eONqbsTKk2Jwlu5rAK8oeX94khAd7/oxECUIEtk4ANRInLpIMv6
tXJnVfb1KLyKaPvUDBEH3TxeCF8p/QzJpZ9HN3e6lIsMy7nXy8OIFlNvyShHnsva
4+0arluJS96pY3oNqsIJBdFgkKBRB5gD7iC+V5hxv3E0ssZgCtoILARSjMuZVdCS
5PKykE7fOB/zBSwAQypf37JpbhXWDQTaBsZCRU1PW8f6egEXKj593SIkrGvqXIlg
dnli/J+u9rbbND3MSUZwYSH+mddf7IZ3HLJwyJxbRp0XS2RmSDm7mukh2i/FYpzJ
4g5xWJGxrhRkWzkCaUUrog==
`protect END_PROTECTED
