`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dr5ljnsC7damCuYgDEfooH2eI2lwAE1dChkke1hv9TftSKBY+aJpp/tNELMmQxMZ
2nC/M/EP6dzwyHRjHxkwk+H6rPgRYQljDfdoBrLbthLVN+ZoHbV1FQ/q1oXwLm/V
Ufz6czpchTTIhhEPBs241dF3/XtPc2rtZLvZbKl2RBftCvjnX4HZif9MPrXuuzUQ
/+EgQmiv5UOtVOSTaeatkMMHjuMd1V+aI2fkQW3xaQuKCs2cJB9Pra78JGEyzcDx
67xS/RpUoHwCYDgyRUEd+YK8CFfscB74uHV1jFDXnthpsIHx5oEc1NuUvGMXCUg/
4eTCN55wqlh5214PmFZlx3pmLO7gIwIBEw4ltceOJBXTZHwwGa1lMelJNNWEdUY8
aCld1MP2VMfkqAkXKU5IRmnewKCO6zvGcCRIBQZPCOfTbdI8Dj/H1AE8ANMK9mHo
M745zcCHmvx/6fX4W3I16ez2rqr/4xktFTdM5sygwuAfyRjKY5+3KoYs47/+iJTU
cRMlfoZLqiR+EnPh3Y6vEMjTzISz6xrQglwRawuepqSn3E/vzsJ6v0RIY+roTfW1
OuM0TrByM7MbONuSGEypCaTrZKdQm0LKU0XWWSFTfbbFJIizzwmxCtnRhm2vIDLl
EYZH7xH+Aq2DZRIMpDOv5rTXGECoNoNVjohHLqmTO/qDwFbfi8tCkmarhAioS3a3
mB0GYyliMTmUbzCgSieYXLD/VQPoSUb8tbjeGC2ASqDREhiqgzUR/bi6IlDUPh5U
t4Q2G5h/VHNsqtWX/zi60+zc7hF9/q4AB56skrCnk+eBQVMGfGnoYRtz2UVvMFSp
NEJMdl41+fbRG/DYN7K/+ZDtJsdIaeT50ooBxocvK9nXFGCm1x+kuf4s2tpGmxhc
m11/mCDNQXc9qootZ0OOlQ==
`protect END_PROTECTED
