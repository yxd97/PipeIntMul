`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KOvwwoLyFYPb9W8E0Qp8jnwc+5XZTCO7tFIsO1O38DDOhSz1+9qJw2/YGNO2mywi
kgDOPBAHaOCV/DRmBd20Tftqw5Yc4idJYht3eoVI06JYB9EYiwGFW6JN9GDSyU51
4Aza1VlkMBjyu+5+4MAweHWJc2l/x8erAuwuAJN3UcCActAQc2XGVigY09kAE7eF
1cnDsWs6P6XWG53sKAsya58TP2wAGCaylyGlsuy2vYK01YJx5wlHNQS2qwLj9Am7
DSC0xGO0sJWFznpByi5FT4cRuCCc7TbCZi1PqJhdyVEoC3My09nJD+ECmIfZePAk
abRklIhI1lr8I3ctwXNL7japKDZ1zW0774Q+DMgLtmXRWpW7IaOQ2sMZAzNrFYh9
zQYwrc1cAIafpeYwQu7lNgqql2fZk8Im7aZ/FothLiZtSaRhsX3RNalhwLbj6pr2
zDqCOg6UyoNcX5nFmBzrvBJsh9Ok7Cvo0J9ZXJ5g7lv+ZPjj2YM5U5ga/5BeHk11
EQU9DtWnjtqn9NMvb0Gw/+Z/HAWXcCjRCXVqos78jow1AXIJlofooYZ5uGqC3Bu0
zlYQFLEZRgGp/1MLWgVjfyIlt7OY76MErCJpe1KUIjEKGrW267Cd4KhJdOfh0N2N
D1M9hi9Sep+FXbS8UjFdz2GtI9HHFBnLiXNqhTjPo/LpqTr/vQZVmdCqO7Nb6SFW
AKOxwCSTqSWY+mj+N5796FLJxGb2htccHVBKYfLZPS4/NUP+XupcuhL8zkGOok9+
AJM60JStr9C1OcGytx879PaHAMCwcUYrszeTJUldOIQ06LmBU9NGuneX+I777P/t
T8NaxcvoRQ8dGXvKMMV/6pRI8ZQ4J8TcLNudk7fU/cqJ9vyUCcuJ4dRVBBeJozJI
aCtzDr5TnVftyg/ZDr9HTKQeaW8Eosp6VVQv0ccXt2v7HYuYaw5WPS59UgTFcvC9
39WQoHk/j92bxn0zMThxYgjrois+zZX/4cTnC2Jt5+ho9ubaVwzyCij7TC12q5Ml
eKxFQ89YYmZvEY+QK2e+Mr3K2Zhcty7xTC2wQK+ALNhzV5AywYI2xQatRjmc0lpP
zJir6hvEh6g2rz6ks/KOmywekhdkG5adOuIhM2vcFj4z8NPfPqyRQx6BsUeLznWG
aJLDATYnsMvsqSdYsfUOYjuREl3pvZcEY77I5ZJFVz1upgcNPRXVpIeF5S8g5wE1
9QAT5LjIjvcS7xqbQQP4C5Sjxi6bkB8wfPfDqdEzXbodyexlBJdTMgo/pJcKVtkq
J6yYtC6R6X1Fl/vx76kwNStPJSz7g/G+owcFrz7OHDRe1pLAAbrkvPXBN/gWwZb+
DDoD+x9ABjOBOoCpKlBRP4uY6I+rPWM/htKiFtH956XTzmj4zkbPRyHMtKAMfFLZ
oBXHzqGK7EiBb4iHWmFIyvQfANmAposlDat95+T6Q9NM8cal+DKh3u9f17NUeBzz
Me9O+PKUJYQk7ausnaFZMAXwsX+9EFJRGpzpFOP+Ge8jRVYTuVLDx96OZyaiH9p7
vPjArwbfH6xFYjC3/Ze1GWBraHjxmIn+RPigOEL5abixW9INp15h5C9Nl/tYBfUa
758zqHnDdZX5tll4EHOy9BxiGvZPhvB4P12UszGgyCnVdrIpuo86JviW5b5tCYSO
4wPvAuOzlSxMO+5eS9bO7NZ7P7hbPH254GNeTLgqd91SJrdieOHn30QFdNGG/N7+
GfE7MpXvyuxyiy+dAWOsJgnnb6L9ARZoC+KuAj0aRWoOp6tr1IPwHyny6BrfwZYT
aswLLRNfEhq0jsmzrpYUqcu3j7ToKsY7XGsl/zANwbbWQW5+WD6f702qIHt0jDHG
ffw4MG073k0v7zeQ3yL9nFUqL5uNVvwZayEnUfzvz1g4OzfEv1Z9/m5YZ7CT6Rpg
LrS8pnwUOaNu7bJeuOpCbWh9yP7xrjN+gMvn3U9eLXOeoBnhqZcVOXZrH9Ao7ubZ
KxTx2y4eFrJVEDSsypCzDoeWRIEvfX6OcKiCHVhuykvyQIXf0F0sk2uVGyIEeLaI
hxdnWtCkivhjH+G4Zqrfpto97zHRV5z35quCjoY9bHF6MR/AUM+gFttudqdHiE05
dDEbILflHfHSw2/v/Zyj4IyTN27VL9lzmCPBTu8kFy7D7p95sTfMBnh1W/iBKBjA
yXIWpya9wLDGPOTsTpHZzg8XCTyE33A1y7AIyebm4+SGn5bkeoICputONjizWD86
ndxQeZomIabDBl+MGWHXkOZgxTXSMRin804GW7B/1DesVd70bWdlUW9vOTr9rtN4
ita2LrEdZ7AMuk0s+UYlTcKUIAL8louD67KDQyz0iJiLvUjgY7v1ygb2GVylHwgH
W3ClpnPXykuZUCfl1rkvhvSVCaFm/PWyv62BWR9zbkBT2ugm93JJ8SV1943/ZZr4
/lva1QRaJ3gjtNWfCON8UOKS1Cql7unTCWvQJYMVujUQu3+ldM3lEw+KIXgV0ujS
YUqhHFVZ/f7e9akvsPuUbjb/tNtf+LIvV0JUI9LkxjJZWNrDJ1GeDo6IGLjm0eYV
GjDxPE8D/W34hRChXgjGGntkFim7WeoN1+DDE5KdjwzlBu4nvAmq1Nj8x/eAleQR
3OdhahExPYIBYHYZSv7TIylPqSX8y3NIeUJRdJ/BcqMM671itPqpsYZRKJzj3uRW
e4FasuopnpMBs4US1ocSuIRjVJKCJL6D2sjxCnApvlhfO3j7drDPbGZAZYRDuQip
bU8oCWWqV7m/wPZoEIfTMsfI9awwzz5Y3zBem6KCSCQdvNuwJlf+K9/RYqr7Nxv6
EQkLy2PDpX+6NC8yMvLbFmj8w4hPzUXk6/ie0r/7ZZeNUgtnVP/c1w8JBojIugC4
gYf8WbWtmbsNPpsDffdnaT2XKWvzeK4ZCC1lIhNLvYaEHvnGgbHTEdXOOQkL9JXq
L9pkxwOZfpeaFTP9p3DUQ/G/tccdhwxjFd8HpcoBuPvJcbhOREoKRjErWlbIamf8
WfHL/niqRg38LmYptPwsRgrlkqQxTgaYve1yWy6q0UXXFLgvifDBO9H11ilrUrIJ
sTZ4J7f4cERRqhnioWANNxbGfyt5TqjCyGVS1c/cqmT7FMSvciKD07JFRYBTQ8+1
IQLvdrdPfwWaAxocAlML/rbZNjIqDNOwyzwh5vXrNahhLcZmnlxQYWa8sWdtfijw
W5WcbaQ/Q106fi8kBwr8u7LYAlLESTFCcwI/rwPDTxRLCJDjtigAvrGZbGy17xiz
F67o5egCivxxnLqx1vG4TqguBBVgkUJq1toa0tFT4XvmxVWhgX8IKh0e5+m2al7K
zoWpuoNnBYONGzDgss4N/OAJRu0CLIuUgXxJcmAdtvtvo8MSi6K4I9eacfnhofjQ
IZrfc6iIyPMT6G7HvV7BVj1IkrcwVAMrvGYMQKtfBdNI+2wpvam96Qw1mOAkj5k1
9QZUMP1h9Mp3EX+bl6PLshQ0+/D1jTpDaZJSkOuzGP/7k1JDscUY/+mAWqoitKYQ
Ippg/hua9JAqJle85sx4zQch/nVLMcVlsag5yRh0keRbX9SajoXIQbOCvAI5k+ts
J3+iRAwNAMO8uTODIJ68ZxVEmW0vzCVe9G4yEFQtA8e/vZCsfMdEfdpXWB5SpKgY
4i/1W6jZ8O8gPm9b28HdDh3VQpvqHr+z8fLnDDthgXbdbAhsNanyE2Wo8zN83vSb
61jxyXplgtWhZ0vOwmcRoxbgSNKXuOA6YrKBE830nyHkyWt9Iecmfw5NNQns6yn/
SlpgrrABp4CkRyLzWVA6MhaC38lVcrYSsMj5bUE6e7/5oaKCv698HYPNQu9Ruojz
9n5xddV/mqOH90QpSwXM0RSnTe37+8D02F/litZ1gyje9nxjCM/xRZinfd9fnEBQ
1wMkDW3KjQr2xRN/bygqLlksof3WC89jbx1bBjwhfzPuvI/9J2pRMaONC36WWjYh
B1/p8Gv4kacRLEcas1x2Nd0Bo++M3pOBQK/YdDmjsJfZwLhOXrBNoKExtljjrgtm
1377SM4y+iQHj6e7BEPqy2jPXGtqtSUFTdOBrKe7L1afypBvnXh0E6mLQ35eDOEr
i2w+B5gA/xfaGDGxbiHDDRn6fUnPSslRw7oGrFrBrfPcqoXeo004vX4yEXnydgj7
mRTMWKhMYMUBPXaONcBz3yaAw/fSMYJFWB+7hp+E66L/8rnhGTcKBeYfH+11HtBY
KtlENoXLK2Xf+c5JOVfwrK/u1Np0TKrlrjnkhFQiXPggTLhumqP6LWxsvLI9U05r
TLrvBP4kBLZh0Yf6bvbiDAcVv/mwoy5ocuIqS7Ndgh9W9LY0G4JQDeWMO3ouuZW5
U2PrWNcyqA60nyt91vTfO0QnX3p6Rx5unWAc7bLmaXzhntqJL/7+G/j7+WwU/ml1
VEPstfypldZ3WoRbpIYhFOKpwYg3B7TqM3mGW4OPpyyA/3jEaUV6nvSyvLUFgqUC
BkbGR0stILInnIcTlc0ZQkDcce8f1W4zcNMrVIruN3COZYcjoS0Y00UeIqapeR4F
cyEFsTY0kPMTq1KVOm+b9ZkL+LiC6O6rZss96d9hdlP27tgi1xTv77DE8RiTmldn
hH9W0gcUcVDEhqQzpD8MGBF53TEYNL5p61XJxKguZWxEZ7tsD973hmXg/utLI/Qr
Me+LitV7iLp5R0lyzVCI+zDgs1IyLPdq73xqnZFv5sO8coSQWOLveg2wf0GDG/EO
QEK5Fol73Szm9vefquhPymwPQvWi8Xc9m02MiuMyQEfnYdZslSZN0RcfYr5MRX3X
wf59lhiA3BcrGKVioojvqPmy/nV//b6KLE6niG5nEmuKL+SDgCc6h37QO3766ssV
jCGXMestBQj01aoxtr/LnifHdiPZ3yj6nZRTrwFXYvh2DpC4RQTNHvaxJEQhdKW4
6mNL+OgFESCceaZsxjy8AHrb+gpbCHF5XjK05dwnDLGpTqAqgzPxqsEM8CkdN2l0
qWEHvIrnwBkBCQeTfXskkalnHmx2PakvsKMo08F6NPvdjgdGLgoGSAbYxJ+ZkHDk
DWUCj3++maGItPwEgDdHNN7hivScQbcOE6Y+E2tdgIDvhU/LRT42lBGxOUl0ihVT
+y3E/UyjQkPyVBvFQMj+0wjlMPBVIcZvJ1B1imwukCFbfPJnwLsGwtthU1UJbTmf
c11J16MsrWg9REqPZWE1scZjB5YLOkYYIOopFhB4e9gYyQCJbv4VpBVJH493KWYh
QF7neGfPxXCgk0eK08ovxGe7IetjX4EeqHJMiehxjtE2+jTFyqEbMhnd4LOVXTat
jc4wxikb2CoGYBChV3pHwN6WyEH6+x8WXEHulyZfTxp20zbdkH02g8CyvPS8T71N
mDdGwIiEttFEnc+0ilQXyY2p+no8lTlIqT9QQQyG3Qh42gM5IFjs+MqpbMZH0gxH
aG/2LKfVhejYp8NIJk4+U68lyFVqfnNNtJy64S4gfw1Wekjlq4pDPQL7eLcX6RAV
1mDnXL3IzdATy0P7va5ttBH//1EOGBdk/TKvBLYzjs/T7bHb2+7wkFNF2hN8UoHl
4WMnhxhfNmX+GLC7+OvQlw==
`protect END_PROTECTED
