`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CW/a39nv62h5PvZEicUfEWLnHEec0AMJ0BnZq3uZGs15FkbB/i45Ydf+jAVPGG05
oEukV1V8hi+O4PgyG6haPs6oCi2tALEqJPI4G0TqIB5ZBpPE5a41/lIJF027NYeB
u7px34m6ZgYvuKPXAFO0L7/HHm5p86sXBAfJ1zOSXj/LLUUp+XzOZjdNb20A8CnJ
HjpSqIkZwoShz6SmcfG6rZuUVL04p6MZltTXGM979e8HTI1cyFhRAGmYDxFIO8Zt
W5FNuCoFctIc1+mw16q9XsZS6Bd5i5Q/tRPVpiYTig/f33z51/uopB5+B0W2sH/y
2SOumXKX6Z2BLaAzD+TsTA4z3YxawTCLpFTlQL0KHWcxseMq6gRL3RHFOKO8WNtZ
38ZgGtEMRl+JENruPJXcAuTfRRt4TuqPXPxW5ElsAYdo3lqTWzyIb0Xt6aQ1kJif
cKAMtqOLJUyLdrAtWvfNj2PnzURh1iC2KZ/dvG+et+ZPPJvV+KH9yG/oiSAvQRx8
v2kn6H2etjf/kwR3SAtXTcS08xypZWiGAv9mzF0ab8OvV/yU31GBoqwN2UiVo/Zk
plvT1FhYcICGCxDVekIODw3HKbgbz5ayDEE+72JdMWUrCIaWFdCv3bcFSl5/F9vr
`protect END_PROTECTED
