`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f2YcQLRQYa1f5huZANUDHd3yo0Hf4hjFQI1PqwQtNWoss5GUzDGWiPTHp/GfmaAv
NP6nqi4ku9eOMfi87b56ezsOmGnLNpwNukt9GclFyk1R7QN8LkSZGSyxv+07LcnQ
opTKixD1UHlYmxf33SLL1Ec49o+2N0Qmuk7PsnM5P1JsEsyiHLTWPpS6LJOIeJ6y
Cp/C0SRc5bjye1t6FPBCFfwGruTUoWFIQg+6mImXhjXESiVzFwJ4xidnJ4TY8unT
`protect END_PROTECTED
