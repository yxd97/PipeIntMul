`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76OBpRa7Zl9u+doy3N+GZfsCNK2wHFP75zr8P28k9GNZ532q8Zta0E2IiZaA688u
TEzJ4tJel62aVVilsqz/9vms4kJBGhB5/k+rnRKaIXO30vELK/DEh7YQFbmTecQz
HceJ7y35dncVIKMPo846PY6HE1/9zNEvzQ7Nzke1ll12pcep8t0BOZDe1uZWvJG3
2p/CyR/jLDlwJ+GEdW0yTpUmTuk3Wean03Bfa6k72EIFy8oz3HwGaZd/zW1WqL5P
sbKe0mc/eVAMEg6zicMxWfF5qO/ukW2d9WgAkBKgOBUCrXT391dxx+cO0pZAnns2
S9NAZf9BvhN8ahqGCWM8fZ56bDWAM1Qn7b0nCfSYUnWTIDDQJNkrmyxDowcK7ZYd
vf6yQT+0LZolrPPYXbR8MiyVr4SBr7Hl+GVjBUqFGSU=
`protect END_PROTECTED
