`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tb+ZLW3J3ovrFG9goEslZRXQtW3FG8vZR7sysj+h7k+3jFG50xismH/OY7hvIhoV
lMb34ehKtjASIA5UQHhQec5M384HUNn5vFhhx6Yk+28By1+oOLTTEHhvhtn2sWqa
DnaDnvqO5SU6wW+ppBCOsQoDCqkkAwUcqvH8i+5WVDEksqrkyaexfHly99JskGdB
ef63AvPRJt7GRGWuYIVIcZmRyEaD1wy73BDzlf8fhcQSSGLrNStv+k8oslyFEB0m
gp6YnYgbC6a1mw3B80/MPAoqaBLQqjEv6mX1gru8KumPDQP+wdlPCLeRRPS82pdo
WeAhxMEev8/qy2AdO125GueaY9UC30bxUvmhMxweBbwewx/9u11TgTvwf7QQDFuJ
Z7llrfCoqLOrOSIxG9pFIZTqhZcLnziv2r0PvYld7PA4s6CEhVpIeDJ6KYt95PI4
vaYeVNjZQ3NAqOHdfpHqzioWEQe/yFOtvNaC/ty6L1KMU+NLi1ajlt2u+0djBR0D
Nv+dO8+3lWdTow+lrtYoo994tCi+VYUJ/Cm54Xo5OJih0+/vniIBITce4sI3AaPc
Gyz9f7jlDswdTA80G7tI8FtnQMTzw5sD5Gbk9UhdcydXSDgx9HYNzBOgIXtS8NAt
kT12gnzgkpau5uh2HFwM16Evrq65+KrtqAlcpsD1jII6GhSB2PORxMue1lCO3h2W
9YNfaIvsqwIXM5SjhCwYQ0iwi+Jak9BBq51JITGUfqI=
`protect END_PROTECTED
