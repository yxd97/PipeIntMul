`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yzv2Lr26fN8pOuJDM6OKQBf/NkOldK9oNuP4/YsPZfGCx4WcMTdM9v/aNV2LRJZu
LWhI8OM7MveO87hBqIsB1s0z8ZWOQvCSEa6cgObId3fCpXkGHfGXnCmPiAOwaPB8
veVl4IchQ5/lf6E16obALLtrg2iwIrCbRhbjxvEqNucLjJ4Xiyhualfvos49fd5q
A/QferJDc4X47LcSk2PCiKINYCSTIp5ffWLU4LzDwPQ4eYaYjEHIvPNA33ICLmRd
nHsp5FkMMwU7/yaBQhzw6RLio1n+oxpd4MH0BfcBTWV9ZxtIJt+2eWs1gTA8ouwh
XxgxJoBvN+wrHBkmdcVE05g/1QAd+gZyJWE2JwgdS0el7UTBRCO1Y4nTIUwqax+Q
RolIfX6FSlBvcH5agt/IodPIBiS3zB+hJp+pd5Sbz74zL00OjKmtXOJM7jie6Jjd
zet3Ow3e0gJs5jaM1UhGMF1McW7iJKpNPrvQJJmJJvSVtN3CGvBQ8DwFf8ETwp3g
YeuoIO4re2Pp1I7KFMCkjXzw/PuJT+qwR+KrAKPGaDyr0z+snGQGqm4eUXS1fkf2
ajLVLQwtHqPY0cz7mnmoskLVL10+MXZrYA7elouOWCcVBQSSMFivmGRCMNpx5uUp
1P4pORpJNbib+fg66Fj7RVIGBRO085dH/A1kVvhvXoI+eFgXbcSNzTOtTx9LiHxa
/y+lLYZNObwlpS2R25O4t5zzH+gqQFaO5TQCtDvC5MA=
`protect END_PROTECTED
