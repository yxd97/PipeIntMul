`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1APqJcJ37R9LmJfssPys5qY6ckdUe+5rsymOn3vwF6qTh/BsR26yqxWO6lIn8FbZ
AumtH0xXdvl7Z9CU0VFUR+u6+KD0BQr17RJE8h5VXphBj/25mv87swAwVnLDXKu5
cr823f9tcIItir2nh4a7/lp4UHcJDhSviua/QC62EXcyI0YaMGiRZdnDOFN7rjDK
O3auFCE8EGKsStb48RPkEwGM06xHDNcaueAuTgLwzNcLPQ44JWqVPtdE/6l4A1po
Pxmy7yCYXMrnAUmWzvJunzGj0Bj+AYK44zL0caUACN52lcjlEIbmr+HTXrk8HGWY
YyQl9Sc6jWexnJrQG1anPoqbka+HNvxoz2Rn2Q4VDKLubBDvfpi3QNsgNy7qBWuH
SLiOdfDvbQhI0jj3AkD1aEKcr+fkJl8jOFOHc89n0JzALiJidGbr74xq0wZiR+3X
R0+tXTDJ0xX3rZQnfYJzWSEz/QJSh6wUoUvsVex2Bx39wfPGMv+gWrJo6UvklRaS
bYEPYNbNjGCMSQT2PZd59v5OMl54mxejd676x3MjvrrkLV8AlmkLxIW1tyzbum3T
cynNaE6WKgZCpKCWgqLldG+rTDNYkOWvWvaksl4CyRSAwz6YENGRpLuCa3wn7c/j
60hxyPfN+sFy1YGgn4c6FRBcVKO0ymPoPZnkJ0EANXgAS34De2YmPyQBUGF/aYtc
VHgHKAlZLW911BS8qas/UZDHHPi3S8UiJ/Kmxf/dawfsO4AbNG5TQTrN3MEMHWJ4
yI1nP19KTnFx1ZW4fi9fMJaSkw6nUC9+SszHmolT9u6fatRWVRo/xNvqW9DVpSKC
chUVpDOtwGQ7rjhOuVMPyekz9pxqEBdZNEQT21VgbJBX43p+CrpuAMSOA/ay+YTm
SePvLJ7PynzyDLa+Z2hhJUHmcyPLssN38itFfZy8NpIZYaPaUrddr43PKJI9y28a
/K9AucSBkxZemHCCfx7McRf2htTADt4JBGFl2YSMiYtbD4QuQGrPHLk9yFcqyIfb
lc4ZZkRAKpuDMVspTQgkMSiBOGsOqv2l+y3we+Wnd1taC8xSuQ0Kk16H95Th4ENE
ZChNt6NK7KcoO0b7GdUuo257jZIf3RYduO6Y6uLO820mouhsmDfYcHfIED/WTwg+
t85SxkxmEBRCE86UZXZ743SY5pqToOCSwmgzi9S2A9/l+LgF7jqqXYb/iS16+ga8
/FgbM8VFryLvIUj2xQOoFkuWutHi14xV3sZTHN/DZqgXAdWiGVJlkU/TWgqaxci2
oit93a5twx0w9Lg72pMzYnzeCQNNX4pj3OWqFYwCQPX1vqt8ItlUSLno5kL3Ly2C
jtFUNS49m+H9gs1fgkh8ZQBMB+XVZIQPoKjqcFIqbW2J3XxPN+thSLzursFKivz9
KnFs+kA5VAQBVp8frwxOZ8BwIC1uYpziHytOp1pishU/0YLrK/PvYqV9epRNrEqN
bDtIkmVnP5t0l5jZgOcIxFuVOC25bfCecN5wMMrJUQLX8KVrHDXekSqOnjIvYboH
M5V3Poc4WsaT4xWpZVdkE3AAtvjcljCD/3T36fibAOzCDWF11595ePKLz/aZGyl4
qssTZTemmDzcAoaW8fdD3WQEaujEkdD/Wylln0NKltTlIhbqyKE7qQZLoQRc/Hbx
lvraFj4+e+f7hugfhoT4zg==
`protect END_PROTECTED
