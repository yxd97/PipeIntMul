`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWX/3eo8B3foAxTNJ2eKJrzumCAIWVbMmzw4g0lBh5q8116/8Shg86ou6ikponGY
0WeAVqDp5TU4dmgQfytoYkgZeOsTaK31Om/iv5Vk6reXNl2XqSrstpdZpCAvKJdk
7ew5Z0eN/PSCa47j+gzlu5tWAwbhS+2nRMrHYJ4DEK5av3R2udyhJ/vmAKBvR0AW
fDXVSejUPa6aoAXBnyb6E8jCTqMcTmPUvtQhrOwu3ealt7LZG449ai3qiQCXDkDC
4SWCZ8L56uNVvBmmSO46M1Jg/6CALpT0b37bjbCxXn6koiOa3M6qF1NI/sRcBYZr
0Nz3zx33AmgQH4UgGMabBtxbjC49kbGDhUigIscBF10sn3Z8pSjLxvnzeqc81ApH
3ccumdclRfT1aSbxaAto2gZS5BxuhQ6eKEx2Qb5DXWgDjkQ+lCEfsR3QLR5QduRz
gdrHrX6FEB9FX4I/3Kv+3sZ18h05GipaQ87UZF++sAC6X+KvVm2hjD/+SP0GXX0X
QEuLIP1ZipsErmBd12lkmrwsC1c490C6KhBF5QgGDeoQ9Fq9NjjXfaQ9TkszwLsM
pEU+F1wOSVFqPaDWFM5/amD9QvdWiewmgGXCQuwQ4HZpnCk9EqUnG/1IXb6LWAM1
FOMQtx0uiBqvCs/vglMkbS2h1zwEox9EMUe/E/jrn1OySdI+MbT08ovis8nvqhMD
JjrvzEQF20XMCRO0W+ufO7u1mi3KqRFhCTsTMMSEaAxWDH9v6DAGwzrTsyVq4Buz
aPzhdjisrVpZ6ZcIpmlMZYZFF6gvaJmupPSW+/apGgq+JaT5yQEpdMWbPugnFrK5
rDbztDrFp4B9yOofoAYRE3cWVsz5cYkoocTI5fwZUzvSuRTDfiWM+QTkqvK2wTXY
AlLRL02fA0fIi9sz0vu2AOBfauo5uV2IqiSvnXjbFcyQPecxwcINvpB8pqPDEPyf
WhsbhB00vSZHsB2DsGw0BA==
`protect END_PROTECTED
