`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wijIiFhYCWy9v+BgIq7f0JnCTVYiCcHLzNYm3RKoOG1L/ckt9eHeSD7IqVonZWzP
CX89qub3CqZWCp+eD3vKGO/d19B6/9u2N45H2cmnLbXwUWOXkKQkhOoAdWwn/ZZY
jqibmwdn/A/texrG8I5DytC2QcUZNVa0KkQLh2rlb2JYjC9P/ojY3/BRTYDTU8LU
Kxv5v3hHRP0Vy/HgBNUKz+h9CrUwCWdAI98BLDiFVzFD6VIUbXMJTplNHCDuRAOc
ighifPS27jpc6xvMmBVtsYPd8YgSbMVZLfDqnhoh545DF8sRWdC0dHSy0ehg2Dj5
VEw9eAKj6wRiWlc+02Ul0bRgfSC6jQR2whpc4hz7Gsjhh/fgrdKTYJ8wNGgJhFd4
+xPgaMA0DhggZkb2cspCm39m8JnUqOXx8L4EhgCh7lwp8GRk1qJckv/4iZPrfg0r
bmm6rYH+se0SMQtCv9OhBuXhtr5QlB0lWYfNDPGcySY2ILntTYAGoSiqQYzm/yWb
NbbKUEDkK2N8OLBjgHoBIsgf5bnVAnZliK5IIubkCNvz4SU0d9o2IAkIzffcSoVh
MuFxdqSYclz6JdiEb5G0lKnOgVA3SORqqpM3Ov/FeUX3CkhmUD0iYTG+i+uYX53t
m8wH7exNn3B4++Rh95/HE92AYDwI/qul8hXOzu25/Yv/7Ht9O8QLuWPGYpMVnjK/
zSHKJCYntAIgV72mKcVUcTxLyt4xmk765uupve2cS/1YgC3ByWcVexzKQjXSBVdR
v9MLDZvYQhsNThHeKnfDK7cUr0xDW3L8mRn6NKYdn7tqF84kqY+s/LtBFIEJRMnH
2hn7YSKK2Yxq7rMnVmpFl5Z5QhEsWkDQpyA/uDIEpjj0qnW+/0c77WtxfdLS6UJA
e9sP0m1NVfhK92HRdJ/4fiRE4/OVip79bmYBiBu2g/2GkJ4QTSBoU8MBqtFQxc4y
AN38gfClQPO6OFP/vNqM7l0pGZvcBc4oI3HTp+KDxxzSZL2zrMpZ+olqMt5zG/1y
Lhhu+EenWA90MqEuezxRYd7WSdrub7Qrtc9BOI7uoCQwyKnhPgp1ftKTStMiXbXA
nawpTfEFc6NxNP/VsWBLehr/NISoIPZ70o4YdNXZSmTs4JSKRAiplUKSh9K/1xkO
igVBjoQZuD0B33U6GQtSZfNnSGY9pLmAJ2quaSGKiCVJ0tC3uXT0/I4d5chylD83
88qiCix4jre+Spg7/7/oiDg8jD90O5QLNw9RzDLstCTcuBKebT+Ur1IDjKExwIuy
cZwR+bAP75qmeZF5/iLvpCUzOwFTYdbqO0Gf7yuBFJBY3jPXTWWblWqnSu7uhUF8
2Kf9klQfmDW9+JbdGOG9LL/dSoDau6KUuW9uthGg3xDGDhUcpq9eowmhqzAlYxuy
tb81YrE/P5yHFAsQqlikMRZ4X0IhNQQk0dvvJz0U63wMfLD9QV/Hbg+SHjO2UbeI
ItetyNeYETwIl4rXae1QvLweQFmesJWjKew7P6xPmaEVgfjx72/oQ9O+JrA+e00K
cNwbwt9+GnQJafMyCoqrCd3Prcdzr/2Mey4pOuuEN5g1W/WPoiVOgh42k3MRI02L
ZdGGnb69CqfPwzsmOiegKqFOHlI/8v7IdeK6NEwvm5RqOEiuf/y/h1Iyk5XQ+e7j
t1iHT25bmPYaQhytKtRnIi9wQp4cZJA+lGLGD5QPhXy6cN6iSuEimxA3cYS+pqPr
ePXPzaRmx5RkJWN4sRMWsLXJlYBhXzflUarCziHJ5W6vPvS7Kt61StnvkIzrGxVe
bZoCd8ad0/qieuxWxmZ2nkRU5rd61tWAtpKzwYjOMNbnemykxD6eVx3NA1ss08JT
3FcSOMhoU+4RngVqq1c0X5AFHnY+WW41/rVjG7Bf9XUdN9t3hclkiTH5RROhxUg9
sj3SBfSZzLW9YExMW0o/FfVfF/jfzobvngRlEk6ZUVRdgUNyNFC4kNDhpxRDYseM
uCc8pzR57Ss6dCHWm2bf8T1ZTlzippN85LRcZ+zwVv6Z5Q3Q6O4Yfk23u7FN8hnR
toXG9Ggmj2uk/hjsW3oV0qs0X+J89huAw2gnVe7F8kbYp9Wut6hilElj2izRrkrx
iJO04dLSmnvFccBjzUDqqPI3YLO862NxykVSHAd6UZE+h+bZCB3IGsoZ22ljRs2N
b+wmJhxkwEQxAf/Iric7G9v65zvudQh5oTM3RCGH3RIFZY5u6RNRW2WgQ+vK9P84
O31ZPrgcpwG+FbM7sC3cbSxJOLdlr9JfcKi+m9Zwp7hXkjPkyHb4UvYoIjGa2Kkt
bWSNefC6SshY1ZqEuuMZFahGlTSBOJFC/yBcFchA4H6DmIGonl7J1enNz57yjPjw
eyMUh6uxX4vPDIe73Ej0cAt+zMJuypfb8bYhNn9T8N0jVcEs1QwE6rjQjR1LVJ5I
gbAFIqyIzDQQb1VwTnxcjeiav7R/UuOjxTY7oaKRORsBd3hmoSvPcisPwG87nhXd
txfSqBK400U31Nirc1waTlbyWVWaddXRwwTjKSRgmz5X4vDi8fg27K4ELnZTixbp
eq7kHGyPgsJst6fk4NqhzyTkzBW4Tm9Mb0wjoXom9GGx0m2MlIL3E7ZEtobCmbC3
gENOM3lNiQtYNczCMaCteNwB9ilXCfs4FMTxBcZghZt6oYg+PObMFdCH7EMU0C6W
FkTigH+8nUaZ2f07pBGBYi3iLKj98ycxfwme+FGR53Wcoh3jumPQ1iaXHQ7gPMBQ
GKM1UJEl69FG4rOcqPhPPKR9fTWylHnxK5yGfxh0XAKhJId7opP+oyxBp85ps4+p
zHl4zw457dhbFDLf6pB9yv5DSGOdW5MOrIVBLuroKLdnmmBqJ8FX0H1hyE+d+RFW
dcZzgsX10cc/I0bsiHMs9bHcqRBfSrA1Vr3orzGqwGOtJFEqX2zIHmyfhnirvDWH
zjvnYA2ts0PHJY7TqPOsv+rJebZlz+qzuceRpEZ/T6UomUflVAMozZrjCHaTEk7w
zDSzNJbiTtQU7gdlpIDoS/TEe3TfgLdP9iqSOBrpS0aI40vTXPdoPI8aIFY7zODW
bva51iNY9Ct47raWN6PyZeEJuZa1he4FJ+xH7hV0VQRpG1/FR51PS4Yhj+6/1Dpb
TycT5V2wFcMsLeSBEU6eFDWog4RrDErkGXQ8u8jZr2w7NpPDvr0nW3MH3nezVvtr
tCKCA55QWzkLxr2dinvRUZfn2UA7lTLtW13ml2++KQPLFJ3irfxKhGgMys4J6JZN
K60360e2bNa8wY6n8MQ1Dpvt2i4rYbwmqvGSyUQ5OCCEA3gHj4XOZjFHAkT+TuzJ
lBZRkKkcuoSny6m10RJ172tXKQXNlIld70P1EINnxjaqrFa4q1yz6k9Em6vIeG7R
lRvx4dQuGfY7a2dptm0TDSAm0Ukkak6KvaSi4E8wwWR33VEg2DKqrHRC7AmpymGC
sUJYGUsYmd+13UDkWz5Fxv9xt/BW2aLYkEbdaZgpQlkk7pHFPwJHb6PUtifMq19W
+u2kbLGehbYYHsFnczFHUQJ0ZeZfaMq9vc/smM+MGssF9dlrGs381hfugbYmB40T
+YBL7oRTonojMhdaJiHXk0lRtz6dcjGB4sCgHWHG/DskIL3edBbjVSC8uG4mrhYL
4iiQPOel5kYcd5iPeWJqr9J49NMple8gR02Gg5GfmnlQ26JJ6oZI3sc20Fmfjjyz
+F2VDKpVEPM5PSAKdLa3pkUF8VqkzVOtJDdQ3qhglFgIAhMagfyRmRKtodmSGfme
kEhN2985BLdXefnDqxTQfBOHfB9meUfZKkzJYozns+5QEX4mrnMEuemgFiPNPwU1
Hv30M0r/NUNK0ghIaFczWvq/zu303TGdpWp48FU9JBh5x0D3bZ4KXfp3FvY7BDWc
xZZzoJCPfXlPtYBNjqbiMgO6/omAhQtEitxLwjD+KGvWJMvOvm2nk4ZZQMqfO5uF
VHo/l2341zLoME1jZQvurkZ15UhDyjAe0kWg/gj55pjzW26D5JpPKCh/9HAzeXLm
96sRPxqcVDkHrWxFd3JC+nUBC71VdZCLMRxyLS7OAdyHhVTqDML6xiLZi6BnACFI
3DGNAOdfAn8iSSvk/zzrVOB9mzTY3Ky/CceTUGaGMtl4OXWp/EpvSXAESqbg3rWL
ckPC2CZowgn1PwoPkje+dGNHjDactGLDU3biY17rIfyEv9+yXIk2gT9D0y3jQpwJ
+BBEC1b5LZMtge/FBHRcLrUr7oGKdrCvrwryU/wweuYQLwKh7NvVT921qB+vIZt3
23J4nBteW/cUewRyCJM1rYYHbr5wCUsZRVsyqGnXv++PXPUTb/PZRHqkz6YWx3gt
nQphz6ls9W/58OMigHuICDxFSnUyq57AjGcTCxjDBRyU5mA0m5AETmb3YNEgpbC1
91KzjLplUADAzA+xaRGAy0q2HWyBxDPSmDT0Ym2qSieVPXnFgWArJVLQWj0F4DBw
HFxqP6R64IQR2wjz1HcACTGPw78PRK92Pg0pX/mZ5L3PSlk6Q6u9FovbkHz5W9dH
6o1M1q4cK65Xrs7w0APqlFPsFbsGra5toxqFz21XSKwHv9tFI3vdfsE7PefilxkE
1U3vtVMcqH+I0Pb1D96FhbYcB8SytIIp/+r3AoVzA1DjHXM50LMQvsGbf1eRJ2wH
BOHC7eusW1YWUzSaSK+5qoaERppn5iMmx4aUX/bMfrSnlPxIO+BzVvjUfRYP64AZ
tIDdcVkacElbKH3eAgDjBTX2uJxIQD2XqgM5httZsSMv+p+mBTLmKxjKWc6VobP5
eT0v+5vQRq683Z1EVmgs+rxF7bFtO4H7ED4vdQyYF5Od63qNyN9yva8feHSSowpg
zh/ujg4RweHM224xyazbl4mGCGJw+nAl8YKmxpYkmtpGnLDWtUcyfETsxPqPmi4L
Wrn9vC/moQExsyIeAVvIbAV2Lq3xiY8b3eJdM4Q3bcHOoXh3Wg76HxCz1l1v3lDH
taSNObQezs1+Dn132nNIuWd+BGm/Xc0Ije7JmvMRtbsVvrkfvolI2OwtEFslozSQ
S1Bj9eMpNE+n+w73AIHaBE83r17ReTsX1fEixU6mmtGlmooiqGylu3yHkcf6wGKf
NVWx/HONzl6rckeZ9fMQx2h051krO6VWg1Ycl+elRX739xCZD2ph2cLWf1W+x9GF
0He1k4XnduSDPWX0XbJyj6yZg1FEcx7rAZlLa/gwbtbbjERhNyPg648Gl1tBgfSj
OHT0+6Ikx+JfH+uQUtoMv8BeW0V7CQsrfHIfM1JrAuD6wv12Ebx69QQX6zd410/8
Pu9FAlwXHm+pAT5+DNvLXYIDeTO70tW4/lgpLrbBdYBsqGZ4frvvRwkKPYfFKPmd
X38JG7wutN96IPrYFHu2AkpueScNX8hQR9Wh4MZbYt8C8sBydfkRjwyvexrQuiGf
dMwj+rZkA6eTAH9zIYd3tjxjOLu3SmLPASJk7JEb+K9N/D1qIzPgH814bHxJ8JJn
9wSTabSRyzd+/+oHmSNVNgAvFjrEsTFMxVH/g06SJEDE12Ey5LYHD3rrRHwSznKs
8XC8EKl4HtgSiTff9uDmAdHhdH1WHo2CWZJFbDS2i31OvEHkZMVB8mmnK3O4Isp+
k0rpDem3EYOghcgoZcbAZeFliv5Vmc7U+4nNhzDKJt8wm/JwCnvm3NFm30VmvOR4
k+c/tCW7cIL03jHrrg+RE6kq+xyRYe2s8q6L94lSSyZA6bXUs2WMd/F0jIR0cZRk
tl141idRjvgCm40rFL8YMivdqfLBtsIbkqo3lr4/6M5uqX5caDSfM0NYaw/GPu2l
33l0+ScoxtiMTbrWAxacjoM/3K0dDn/0QvfD23yFYIa/T8alAmaX+shLoYCf3TKz
gdoKkAiOwvspWJGVFY4bUFPYMJNF8LfJEwfCnYSevgatrfmUGng8MhcJKK6SPZxV
OKA76rFeGJetMxVnW5tNRxoQ1HwgzPdH8m6Hh/8xBnkNgU4h/U2aKbXttcqkhJQt
y7zQk060ch1eMu0E+Yeiw2SpF0AivabVuKGSNV2ucXE/5itWdrOPPV9HUaE4Den7
QKgBR/FbujGLqyBybxy512gtsual7fmmdDfdw/8fyudLJT51CkiljzcTCWLGmFUn
kHN2ivPmNoLi1m0cTS6LhxbNU9p0FE4qceHWgdYRh+hGTTH6NNn26DCEcEBtnSae
JLv9htwnKK2NvRT1nTWidskuyHLyumKYcKAzr915f8JcbwCPi/5pzG6l2mX3hbex
F92o7WVNaoLFQixQJD7OofisEgtNNekxLMU6BtOgZsqdWlNzJQqhKEhshRnwv4G4
RK02jALiHc5Di0HNvOZLubf8TlO/jAmAGm4h7176D07q6yIDucrmdRQsAHankRrz
VdjwgbGMbI7hL0dPgcVGUcDbs6kk8nBxKE8fXhffJgIKdothIWd5tdl0LmWqjMFK
KG03a+K1cmI8xtNZBMUXheiaJ/wc0hyHHfHFaVvjutCLNDjisppPqBz3JWVxI40q
heE0tYDvMwCopxGhfISA4SB58oFMN0t1WPBDl+8niz2zmDaBXUESGiSXZGRNO+yS
+i5yv24l4tvDzBk2Jjh/z871tVpHUxeozyh33wa+f/QRUZ2+xZdorBdh2UbN9UrA
RGAHC9ofsT3jM0MUSqA2IGaMf7JDh1szByurHjNbrA9oMJGox7U7rMQ9lMFkeJS0
HmcWJxHIETVOb7uMUFPUwad8g8c/iqOmsZyclve8x15ZMlaDRwHu6gHzRFDjCYjb
xnijnbiWxJPHYP/QwHWD2Kd4GnGc3u4fzhHgxXr5HjpVtkyl1VHVQuLPzJztpm/j
zT751sKpfdDUBziknTWR2ydE+me8wU5SF3iMjXEtsg39jOhsqVG8mcq1Mj+blhSQ
kM2FBruDvZM6+dUmg0PZTtIJ4yadlZCin+hkyOmaJ12pIf45CVEPaopBuJWYoBp8
5QKweLXzJzO0a76wT5oCLpjqjR0R0p9MlGa+KlV6Jp8eTnNODGb88bXdpL9tDP89
pBFJyPffw3n7yFE0/FB+2RJ6b75m1gzPDUk9iD9U9IeKcKITaGHpwJTcIP1Swf4C
umcaKpLu3g9v+JBXjq5KrIoi4YMkn4K7k0SbwO/Lzv08r+mZeiPWxYS2secfy8Ts
ux3gUxV9dv8FHGbEstbzQVBx8B6sj5pTzuU7APHkeFqTsAm+rTMRzSJesit/4XiZ
0dzrZgY3k34Yg7oxu1L4f3zNAo7Ops0UOAIQotKvX3zaGbEcLkusGAR9N3vh6X/c
Py9duXetiYTvXecWtN2lnvu1bxQVf84Wkb6SIdSEU4PyA0c9qqMTp1u5zGic9TIX
qzIif9ASUOLxjkQcClfNtUcL4EHtp/hZq0ZRXlYwHIaXAa8EvHlV0ClSmnYjelLw
mTre1iuED7J6NM424idw2hQA64ebwJY46lr2RjMRaxF6cOLNp3AADmtsg4AgFMR9
Aq/pr7sHo9D0rHEryIWCV9iu8o7Oo8wJnuuANT2JAw+U2hVjAyeFmg1I7TZEyqZm
em44GD3invZ5+EjhJm++Zau39B1RK/kPx0W+WZHbMK4d9lavfaGmle6EC8hvYreR
iEXrx7+Wtq0+77pTq53Hu0bCNHV18y5XOo9IrUAX1cml2Annuh7HX3EZ/PJCQYRo
uWt84ahsa7kNIriFxZw0mn8yn3n1j9gV3bJXP5Q5HJOvveeHCuYWHbOEqhU70+yA
/Ob2sLrSX1hoypzsUGskzl2mqfvV3ocKBcA23whXXcV+E64WkM5NCAcpA1AN14j+
XBq5BHaS0J293e/JrNKt8qojwLkkSfK6KS9bj62AsOnx7rP+0kLe75q/xhjIVh6l
wUEpQEAYsKxsQl088sQ5lq5q0y/2G89k17Cldoqpfp45VKxouZrs/0LSWFFYwpkJ
+BrzFfuG8Isaiui16Fuvb85FYomGE6uGcJdQh+B3cW0ImfL0SFtBDXVuYXrZffsj
45TIMBgMoEMJnD6PnoMztdAYfCQCDLvMk8RM4z/KzxJnW1ScBR+mwxn1Xco9dIFV
+Bf7/dDM/tXOmOSvyohL1NQU1qqLjeXwL61O69IZvsHducnwBsoavNvD3r6v9y0S
1xvD06t4GKe4wUxZiJd6Fu2Y3beXqjUNb+KxJWP9ccRcoeuRuCzTsCjKSNXjsoCZ
TQU7sGIxIJEJkKbWZ0lArbZNWMY0LZAZebDJ39SSRZHRerTOLZ0kCwZfOcX25VFu
2V8v6d2JOYwXfdwFw/grR1VprHEvtatwH2nRmIfXYA78AOony6vyelEC9aiwZMLT
Coj+wr6t6/+51DYe9FVeZWntLWY7zZe6QwWV4qNciJHqYKWxF8cpLMuJcJ55/XTO
aq84LFZ10tfy7/qWXAR/+x7ICiNQ8E5zGsuj7jfZIk4vOIBtFhD4WRNlilRqq/f/
sSW9bGz0Emt0ZrPKMVMjyEww31+PjeLEZLmyO4gYSl1nfDJL5sqhnKidBoAcvKxP
So+0YNReVgsC4bnGux+owk5K9iPyhUSmYGgeAsce3NS0QpEdNvrr60DCxK2283yP
GX9Ylp0/XC5BBlAeC/wWJ0q0kgcOqbcR+srvNOFnvay+qrd1YrYNVKXtqN52ZcMX
cNauN1BSoVntxIPYabn8RpfGiSILdJv2LMPOobbrN9xp5wT7Nt/q+LtTvRS8kGo1
0LG2t8PAcA6A3Joetyq98kNiZAZt160DQ+Roud4haUliaUYPe5/JQ8cyQHTRioSL
7jLVelfP4j51WL/zSvqYoWd+ZGSfxEkMBQIhI8cuj55pYGRThLM2b7JqXtcUFApA
jp1nZwrp7/Srm89WlJhokDfpuqDuMx3oT/tSjCCOQdA3W/1K1LRP/ExcQNAiEZyv
zpn3f7joiCFZ6AdXACoYoVb6QEMqhlPcKLIRNuPv4X3AtRQxw085buJR1+ek+Kt9
SDZljuKR/i/VCEDaGSIFxwKtxT5fVIfvtK2sj9xI8Fay0q97qTYavMcpgzOpKh5K
jitxrJJm+UEXGwegH74GPW3HfqyQD2mB/TB2GqONG2Q2Uzf45LegkGhlgeisz+tv
uQaLiVdm/i+1ehIkXP8HDKgANgtdMFwS0gT6uw5VVlHZzSA9uBWikqlZGQ1Qg141
JKVewehSmAObx/cx8/nPvA5cQ+8fYpEpu9H+mvkvrSjQNqDN6hktyo61RZuYPQSg
irvO4eN8tvkdbJGwDCOvsEBKcGC0YkbXVNSpZgPLr0Jbto2OAkc/gzwNby0DMGF4
dJ/1HoewZxzSeM7+DRB4rmKjHHm9gEKvqvtUBFCJKnd4vrsup6n4TAwyWxeUDYrJ
5gtAeR/VEPy3J+p1uY4gEcKHNGM41k1NG5ZNvSzKi0sdiAaI4VWkEqFGnLeNMwbw
fMvECLagmzG35juZMruDhN44hiBWZiwyUyvpypPvOFsHhuHrofc5id152nrD4aEm
P0kaTgWEf1njKBSABh/V7PO9F1bBUI5lt4G1qqR3EY6bf53wI+rHjUKxf+2dBXex
OcaYoKdAiefe+Yvoi5WgBYcOG2Tltl41nnl0ErRRrZUWHuf7TgXe0RzEIWUO0iCL
n3Z17wfGXgCPyspMQWd1xRSrU2RJUcdgvPn2LkEOHzwVSI8zmj9f/BRUVEgRlYLg
RTOuPOUXdQvv9PRlOVI4Dg3YzdlnofKviX2BFTjG/wtszLG6YMr1DBiSCX5Sv6K7
2rxdNuvTa+J6gjHwwB27lO4ynPOUJdTmjwf5+Fp8UR5aUID3katZ3FlPXENe0Htb
vJWHEgP7UCif78x7NIW9rgWggvJ7uGqeBkcGasLMdYj9VSp7o1TUBLoQeLUpEdfl
JC5Y1KwBZyi/vRnidmm5st8Ou8jZ6OKbnrOv2dH3Cjjo75immRU4yHH+6xdWhGpM
dFcokht8HPTwI38nFreO2h9aaY74+txxrKn860BqirFIpB+d3lfO80VknMXo83iN
adC5l+j3FRkXqU5Bhf4RxNLG4dmYgZu2Hbb/KMLPfsfXW7dcYyBwhhSn+RkmFjtJ
wjG0mubO74JyS3kJTiyDLdZFKoqRZ4XpEs8Nafmzucqe4rhsEOUj7/66g88X/2xC
XrpXbsPzStT1fDclK1pdU1rEgfyPcDiCYNgaIVsAE57SBgNMGXTXFPw3pdRADGeL
MbaZOx/7lWolfOknKtWKH4rbt6rhk0+Swel9EnxNRAXQxftmndRRYq2zdcFNrUzV
f+fvtPaCBu+iqL+gC8FPridmmFGjjVG7l7mBnpFskxSdOzaP41xt7cYfCv0+AvHK
ZMCfFtGHjLJ4W0a0CNFZSJl647AEwTkumu7iC7akPBCJKOPCVYjeeGJK6I0yuPtM
F23tQ/Y6n/q6B4MI9jwVq3PrsWP+0q6rQztiXC2x3nmNXZhNSVdZtWQacaIqH7iI
Q/PSL6lj+JqKn2klhcnjPzSNhABFV1QX82k6jO/+lXXDrE3Fqgojpj0/5lZv6PFb
f/nQSIaDH1MfEqt7e/nrM/3bsmwTRbAlm71rJ3//S2JKZ2G+A9eFt1bX4xbVKpzb
nf1GLJ77qzA5WfJ6ZezcG6XQXDqWlwhAwzFTeQUmsrfK8tjyx8ROns3Pkr3R7piJ
WHzfliz39b1oN1HXsrcv0o/5KUZAIirKX4DwG65WgoYyy5IMGY2CuwOee/wJ7JyW
NNyv0g8cmgvnPIeqdsEjQlzPPaMMOEqb4Jsnxi1RmPGMH1m6jhAi47nWghcfW5Qh
VBmNQyHRIvMq+heZEYSFo6lqoFKZwAKHVCxdhUEgwyodUDKL0FXV5O7KW7lbLaJp
uAN4gRRjmyVGPFqhgsUk9ZiQp4zXZcar9ZQKn+UI+eKe2t/GIuRieTt+jwF2YUSd
qTyLLt10/CoSuV+RReZGFnuEZud1zE7/W6i+UpK9KksdbxZ8V/lnbyWQLlGwCKON
D6PbBZCyAfpEZYdYOKvqTE+AwMDJEGeGC/GQUqCXitXomlI7EdmxdjK6xD2RAV27
JKlqs1G/NZbmG3Ql5L9+NoR/s5NlpOhAeH1syyumRnaEJLpFqCfyttBZNbOCe+qz
H9oznTYYbKgxbJejqmghcj/w7kAWHMu5nYeuFF9/NdrqA0EePX9PuwkBMvddEd3N
8jxdxIJqWOS23ngY5hRdjBSzcSIt8s7Ad9b5wLMg1peRQy2dPlG7hNTgnSrQNxnn
u5DiKnwme76pE/B3e9UHRxB07T8p5oUEuhWOk5oOF/766L3HLiGBi76yOb+JkhhP
01UoUhEP6RdNOlXTNARV0RapkJqAYnmVtyf7xZNE9SR8Tm0ciYEYgkJ0+hOoxwyD
4935mA/JJTWYd+i6s8uNJ//G8+lCe5kBrmI9cP92Vcuokut5Xtc2xSoYZw5Vg0VF
OtlNgywn18YKealGgY5BDp+G2LD+r2htElmeXXUY2MruclPyt3vtbYDjunyc0PEn
5DNqiQkmTDNp2+Dl8GHzZ3NUTMv6m/MzqkOnB0vbMYkj3nwHuznDbnfcWFKGKCyI
f8CKHj9JfZ+TcU4hKOVn442sZPDnlyy/61boqZrpSTsxxgAOTTh9ZJZo/jwnHnjV
e3n58qcaesS7U4okY6gaZOZlfigvyRa3pzzWnbkPZ2Dlmw1RBDfjtr4bmK9Rldsc
OVwysi0bBi3MyVuIbxuMDt+XQpH+J3dJSrRfpifcAO3ugTLEjsQAsB5gYb9SSLnD
W1wFZu+RzvCamqqEbREa5meJQiDK7KSLZ8cn3ZU+gsczZY8UQJTx7qxcwhRAtvnh
g9bvMNl7iL2SkYeCY9BO90UzN1OK5kAV40NEs8yyS436bt832TMrVTmpowWZgI73
dFcBPWJ6TgZmqUt75r7mDeQ57Y8QX2XYuKzxdZNxmA7WRk+KEzQrkYEZSSArL+EQ
s5/PuB5MCnS/l6dYlcNI9S79gkHhZcI3MIbOu3Sih9Tc+0TDNHh9SXPDOr2BIXwD
poklX9z5JXsHrLF9af4XAaFp/F9fDcHdXsk0yCndG8MnDl6mzuWrJkL6ohlRE9US
5axmvAidb9nmWB3js6LDvGkQnrfaLdOICo85pY0cuIHkBbIJyaRa8UIYvbSAWvLN
Lc2TwMTqOG7rssEhT1G+V2eqCitAtM4SpaxVDzx08w+PcbLDZdxafnO+zux+U8Vg
59MPqmQVqf0MbpnOeRaAIzZ+iGLlA0hOAlNBBY98hbXtR4OeI8HVQqd7uNx8iClM
E0UcOqJYKVLa7FltIDXshQc9CyGEajVH963JAZw1IHoco4Pya6EUyh8hVSkRcns0
ys/PEv53jvlYXtNxu7LhSQxXae9KC2CehIdiAYUxIrROjqfU54KlaFpXaqEht1pF
kvUwqoUC9/cwVtLfpltEL6c8WQXyG8Hw9XHAdZtGDHmZF3eciY+bQScbKcZVwr6T
KtdjCC+d5wtaoMM+BTlVbRrcK2j2KsnuIGuksXf3lKBCP2YMLDin6mUcSeznaxmZ
XjJMKUr8ewGUPSMNkRadH6WsqON92UN2DBF6MDd3qyvWxMaxShidCxz0xA0HWzlO
I60PYp7Ys1lWnFJ9dFD9Bcw3n8Oy7eAFR/DQTAywH2yu15Eo8w3LXBUF6x76J08f
YidWQGHud2wEjgef8u3DUjQGcvqYWNcWCQbdsYxFdmODbfJQ/wCEHT6dqawdOrJk
RsCU52dGPsm25nSRSsWi9ALFKcDu9xVrr2OeCexfACzkufV29R9ggWoGNK/qfr+q
wCZx70UVOD1nzRUpIAM5Lma+Hl41lgxsEpGX9rMNBaRux6GK4Njg+lG4M/plxmXQ
7D03gWKi19OFMAyFyfU5u/aCZCay0OZTbsc9WlIiiQBWgeWeovLrlS7J21Jpbf1f
RTDSmZhmsw68OqHEwIX2BsnV54PmbUluktetYBYGoZkNmF0R/qVRKPBLPxwuq27R
ra9mc2lAfFGwYT2/5B0HIs/f2ovfetiDa2zZOR7VYgOyAVmVEQ2114Vbf5r0EnqV
0TjwRLtiRnxIoDvZpILcsOosKweNZkZqRDU/Z/5yjXDF5rhcIJtO+8gRm/8Th5ya
uBzDV3Zyxia7Qmam9OZT/VqvXsj0OjzZChfOBsnkFb4rQMiWBav79MM9ptCW1Kp7
R9zp7Aateg5k/VgkBKAHAaPNJVL0IN7+WmRqIPWL6OKXrbtZs+GJgrHon/1+IF27
xY5tqMM6zb8Go2a3AhMiPBCp66HEUVSTX2no1R7RqvzzRWruAmS1Z1lF6xdoQ4al
2TXT+Ur8noeMUz7nY6hY9UjjrH2BQ5T0zQEtkZ2bVDNB8PD3n+ad9FwrgPi0qXWz
YPOBLhUzhzgRIF39qLQK5b1IGpDJh4cBaoI3vIHetOLQvcIZhtjhVNyPPAlPdbsj
FPdvNNGZrR84CyEP+BDbbSbz9jTUoP2emEpRfHG/SqgqtlOWiqhFJYDiRYXdaT7J
2VyFZlW7VNiiZjGvYF0vzrozg4yHbv3XBltCsJADk3cBDLE7s4GNYXud+FV5GfFG
yVFNGfV3V5SVTBhLsPgR55PjVrrWJsigLvx4MSpQ+mP6L9g5yQJ0KRuSCW8WU/eW
DUNGZQrqWgdG2KHo8kV2cMEFpRHPz7eLNVVWgaNtgOnOYlU8uJrFub6BHIqMBHDX
jLPuJURrBNGvJQSrdFH5YYASjasyKpERIErCbhCd9LlOY1KERKrntWtxSu4gsYYA
keU2IqFeBiWnc65U5GxanXKxq4oHDIY+EeMS7yRVOb0mG5V96WwB4RsADDjjqj2H
mg9JGCjCLk862PuGP74CursSyJBhJ1WrT1F9RG1dCgYmWAod8qFQ3zR6SWdLw+zx
BYsHtdwud8h9R5M6JRWXzTidkNShvL3d8vz5TAxjRuaapViraq7tArI10ONFHdpF
Xv6JGoLCiS49XRHTBHqDOe/RwjReGzNoCj3lw8zvtCerfR/MSbb88XGHjghFauj/
lxFh9CRzDpbpycsLgZOzyZ/+pZF0q7CJckQQqJ5HdVVYo4JU2QC9dxgHplxrqZLR
AVSHcp/wFCZqBx67I5IEUanHTkVuwZW1P0Twa+dLBy7ZDFUKl8chRMXHCfsittuV
NHjhQge23BQ0W7QElGn4dOkV2ZUZ4nh/g/7aHma116bg8QsRx0ym2ZeEVGVQQioE
QHd8emaHJ7LisJEetXlDyK+QiAlAqQ+BMowTUfZZL7Hp6ehwZ7/uHwFAUfQ+tua9
YiePqIoiutJLoo0nNkUGtWqK7yVOeEzlTOUXWfEEQZh1Eu/B/uHoUR6QPFmB/2uh
gaecQZCqcqkLGtlWUSbaTM9GuRmsQXQVIiODPQJ0RwMYwjqDaDNCGxxwQ65aJ+vQ
FsFXWCJChP1f6nKaQSJb4iS6ogGgW3hVmvH1sAdkEvKDLy0Rb2Z6ZrFpyZLvZBcU
pK4KuvY5rxed+exw+RCrG9f/1Th+g+puLrAGWC7YEmv+N61xy8FMyErEqgPcfeeP
gp+S6qzyPwyZ7pJ0cyGPdPEhMqKCfJgyL7iMirbQU+WvOLHTsqmhUBOaTrKj+yef
TFsOLel7cxMMGAWU6vb2+GoAPTd/zQJnQz0u9lOAFgDR26E2CuD5VijMEIGJTVH7
JTUNcStGRlPr7GkGQ7WiMT7USqpWRHYec7QBVgrB3EPC445ghwLc6ztgbr8hkP9z
x5jvKVplVcy/LGmkl8eAc+QGe4U7GKfATYI4jprzvER21rDc+Nx2cjh1YR52Ufoc
C+no3tZVmtrESh7rCx2zWvVArLIV8wBKgeW/Glc8VY3uONZV4akVoR41B4gNY+5P
DPqXdXgdoi9+KikmTFnz0AlpJypTw0pxRLGMZ5knYSbQhV5kVc05DHqyGAs3ZPiv
ln2kF8d6OhXQi2nXC80yXQeBMfXr4tQOviG+lrfQQI1OppJ+3ZRDh/Zo6j7M7IVU
lGr+QkgNnvi1Nz/S+TaCrunfkQ1qQGBoA0DT8WFze4iTFMTrnreHRiSuE9KWC4LP
ZjCW50EiJ6SYey7OLL+OScGsCatS0ClTZYe5UP5CXdaxY1yfHaQv54FC81xuN3bS
eFgQ4+hAuQRMop4wCgMviAVBoJ1IlSzwIAV7dOOnF9RjTnYKQM3IxD+Km/vUSMDh
YczKejkrTBpriD3pOJJGi1YkO8F//QqcC67vHxPIOS5rCi0X2e1knu8E6clnRnHD
W+oLv3Ufzmpww2RpuO1otcsTrAU+3R/R/kPBKDKaLUl1cjLJuTHqPck/dO8i+Br+
ip3S83TWwUdzp8rb/oTD+GywElA5AoCe+ePSC8Zp1qWBs1psQ/Jia82G5zOD3MwR
SxPkw1CzCxNblTfO68CG2yYG2Yx25LSQ34XYKl5B9o90hXaT3z5m3AUDHGn5bADq
/Pei0Ri4qD8N3otIx/hrva6m75uCJjziWQy1sAG7kQlpA7/XcUxW8ln/UM754t9k
ZJqlaLXLlSZN4uT44ZvJb6CY1+Cka9lRlnZQreLPczyI7TebdNxufMzOEFX2sTI5
FC57IZcjJF2sQOAFXty6nvTxti+y4PL1bEBtCqaPgrChd5+Jlvkdf0gRltCReguI
qNIedNMpM9hwEmr5hAcRu8Q6gjvUx/jX7oApRdDDRDtmHQksGUQem9tPfuuo+Jib
xfNFVyJW6YUwV0RRcNg/DFlY2jjKu4TFSw0v0l1a1QzNbxSXg6MEdFmfWHd+fHyT
OAgFFv3+G8OptHrrqDxvPvwXvSqC/B7DtX+A014ISeJ3HZj1O0PXOtwqdx7LcHUi
WvDAcoiGis451uDkN4pUTWlsKkgXetLMoBz5jYPVunJOKb3wg36Grjaob36MFmd6
CfPBqX5E2xXCCNSKVZMzmXgwjPhPEFMWUsA61m++H7FWVLRl1PDEqPAGbgw83DpQ
IICI65hn+M5NTT7hSeMy/x1LHDAXZ02FWhh/zCpYK46ULva+Fouq5MzNaRaw9OlU
DJs5djeNkpWFlFHXRbUh5XuBarvL5Khh4SoJygZNs2Se7JlKFQcbFfy1UNV+ytzr
lwW9DT2b5cjqn7bhE6+bH6KBq3X6ynQVTDuRUhMX4qSt50Ox9x5ISq/nF4VLhBLR
1ULY0tjAMyYPx3+qSCxIjPneORvSg92NDCvjU+cnrklX/SvpwbL+68LURRI1alM9
vXXMqv1qftJIQobfGexCAfgO6w75Vzx3tRAMAKdxy8pGdlNK6QRXbkFQ1IiZll5/
hAdMW995g5hXbh9gBZRPBBstuk7XkTGW9P4CGkOROHZ8kKNcBvvcy0R2eyzUI7zc
+lMBt2QrPBZyXbhGineCSsoj4KGV5Fmls7yKMmY6oP+S10+05djO+0DJKoUU3/JU
+YUFERWinQdYK6jG4cxze74he4qyXKAxHTswVvLjgp69WRjPK9Ec5k1WOiLr8QOY
wvOttHveqifYaaVgA/NtdruxuKkbfH0RN0SwrajewUXwO6yLXdhGzNlaaxrz7BA0
9BNZVt+elIzUxg5JG1QJy1BwsV+0wl9KysXNalt0ubsfGKTXyG4zVN7Jsb17hpqA
hBfw++qcziXoo7DqHlY894CmjP08WTtcPeqmUXmzbgWw0CwGLovkXCmhUIYOQsn+
5l/ba0a3oWqdIvkHIE1n7fwmtUCRgcW9pgAblxCMRo/n0hFpmu3hGi2XUvIsAvpx
jajzeco7yPNLA89hueDRiWVLMNOhK6Y1rsjuhap6ETRjJSuSTxFsVXJDhpXVIRSb
vRoHodUfbLNvyqh3VGcSXeJYC5x4LP+gUnlYaaplG86YGXlxRtctbNmUqAti3MS5
9sQX2erB35389VL3EA3s+oM8ZJndmif2uVKX79kns2POC49oAyOZ79YJQSH2tEgS
/7h367YBDzS+R08qi4NaAG3E5V/iOfTRD3/cGFzjEzCC4yxY9+K9uwf0FBzRn4ch
JHXz7yR/CqAeHJ1IVcDKTaFOMQgpPl5fSqObuucKVTlAwBj8CVcJIJaRR7nNoCJy
wHerlCTpyFJgAIuMOzHmg0QPc0ica3BLMrDVAqZ6/LY=
`protect END_PROTECTED
