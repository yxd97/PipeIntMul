`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66S1ByenIXVTtGPLYlItqepMIc6vpgp0GfQoAVKTMG8fOamDxXbB3GkTxB8eLRd3
rZTFOyajfRD7wRX53j1Z9XFXr5thjMQHPpAIDJLm2Iax1x8cR/kPkYpGHRVtAEzO
9p8HtMfwcDLTEWBmqHmH/l+M3eMh2hgARWEOHsDJUpnHzLUbtNhy7+Vu/F0fjFTF
rA1VV+g53/2lqvLp8zlkGwPNtKKt/FWwDRnUcixAVDvRRIpJnlHoXs+Szi3pjGVV
9/L/mbEncKn7qaoPewhIrZdbVIkateP/HRuWZzpKCuBC9+3ysqTFr9nYMUS8wa5t
YhH/grlB7DXwVJ9g1AFKE4gMd5TDvDNNE8YO4XppnKz76fWv2ujfG3CnhJwV96YM
hSqip9aqUUyVui9/E5Osh9URyo4Zop3cUs94btQb5OVdzeiy1dOtf5J7uDqt32jL
0qrVveSnbRRjfEhgBXobmwby838NmZry4hr1Dv9G7OUR677JEzUsqLqd+PlaOkQZ
e9WNWjFZ+cXwlIqu43MYzvGyogrtGTybH5WOv7gE+j7aaxKBQIIS7VdusjQvKwEX
QDxb/RlpBBu0VcBw8MUD5VXFE32t+3fBRv2x/w4JpkKFTnpiBIiWeFwMsUtkgkMA
N6z4dI7kK+5xM3rv42ALO6HNhhLYLq8r65emJDBfG8X2GGdpELN6kqAIScRzNPca
Jt7M3L3NwVrKK2zlpem98Q==
`protect END_PROTECTED
