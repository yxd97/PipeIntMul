`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F1JgiuitlfqWwVd9lSZHjfkj+YKE4wUUvpOBQQrZl0wuuQMQMKcRb+KJgUJS7oiy
l026PTptKTEM6rMoTZHCEq4FIFSsBGjcOYlBad+aOLj+ejm36X14Ob1ctuGI52xK
Ly8sWabPQfAydSITklzQCB1nP4SYj9xKGhjgmLbgpSQGL0NlCO9afSSeKuxq1JF0
D/jVSuchwJ7KzQQEulhkXmsbNQB1LbdA62c2GIaUhgIkXcGn65otpHL0wfkCAfaj
RPvZZ0veljo3eZvC95jJk+iqFdG5bh698UmbZ1ThmSR5AzVqJ100Q1WTHLBClku8
y+NzNkmk9++SNlb/WR9ZC+qYg5huUwGFr0wm5fYuMPh5n3K5AN/hDNI41p5CLIKB
KNVNO397xAbQ9N9QIjthkAsNhvIUO/au3xA/EahDZD2AhhVx4/q0VVUXSzsQlIhf
sbvSv7q5BlKFHDWRtzGbdX2QYHqAWVQfu+2AgOMAPhlBmsWFx9W/UBiV5dHsFwTP
xJvAPzbxhz1aDjcwdYpkthezuVA2A8xVJjVgdGsgX+aSWIjFLt1bq22kUugQr4Nx
Gkd+loaFTaVL3xNNzEnzBhfLSS6tJVzU0DY/iZEloR6oIVbwrHEbPy/FKQn/tFBh
+D6xZX/ryQX2k1W67A4vW6N9VFmt2NlZvzsKLU8VOPQ=
`protect END_PROTECTED
