`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LuOfZnze9Kfb5cqJ1cCLAS1Vm/b5C6rozcCHLydtRxiUqxIRXNmiqowU2ZN8gcUd
b+QRV6iVH705St6t26QPu8i3glwinloXe5CUILR2vEHCPiEpmBTTW8CIy3QmDFoY
vyJD+IhsBJnZ0Kw8UJimL/kitqW5MCtJX/OS0x+hWuwCrTlZan/ci4QBUddSH8hW
17fNmLBJ3Px2Bw3EXUHdG/ISkR6ZdwRIj9jzd2Fbyb/TpX9UXx98NKRGtRmR93BY
I3X37un8qrAqcFdOjcbEm9AkMJKJ2sdsTPp/3m4KHmdZD0nGpr+siEypgKt4CVl7
hvl7hqGTtLHoudngDlXn7kk3Rhu8Ure+zfWgl5MLZDfd5M1yESpvOD2XvLR/dAVh
oupysxkHN7Y516aKevpD+d6hUNIm1LU3J7F2xydRhWITjl89JykLSGlrskQNF8Ul
ucxT4KfIbHQ+LEQ0Ig9W/if2MpALEWCZKRErxpz86jdOFXJKK5Hw1/D2Ide2Nslv
MICqzDo78AwFEpSWiJ5EZqbHN8CX3ckpsPEdFR4SwgYw4j2QqjydScw9xFczD/gk
C9ehc/0id+s7vB2A/mCfBYZPvaB8T6mdXkGFhB8icW3enrwpwu4lGx631qVzDUNL
u+NOXXiPvTATgJ7GQUxWPA==
`protect END_PROTECTED
