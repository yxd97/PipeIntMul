`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGChb4Q+hzSblge7CpeBfqywZS9KgYWScrc99EL9h5BbZqg7TlxPdECN53lCfjJc
6VjM2+lleuXHZf4LgZtu18c3YG3CE5F1BVFYM1Fe9DTC3EL678hZQRF90OgYnD0f
8n6aL3Vf7I2hwZJKA8NSMlubF0lvVhYdmCt+2PCVlsYZ+mYxrjpn65pnmv/bIZ3i
jn9oZHwqrroDL1hQtC3FdGtHJZr6dr+00VDa3ommEDcZ9WhvTC4qS1r+ETbrGorY
wpYeOcMmswnYQsgbOGJ1Fw==
`protect END_PROTECTED
