`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6Kwjknduv0ZB2UbDFR0FFvJckn5zn2zglD7From/V/PL9m+EfAiV/BXeLwOfXOQ
4ofZp7/zIt3PQ2sjPCgR/079FiGDbzx3sslXQn6GViL04G4B/IiBqQMC4Jlq1HSQ
sz+oPjisBjmGObJe4O1rhzmySINQyUmWmq17HbEL83BeeOd7krMSI55cYuW0mxVT
lkRTkjfYTAOvutP3H5BYj8WvW3TyF3LnF0jcCuTvnR/dSqaHmSEj2c8+yvhp4+Ny
8w/SXXXzyW7Ig0H3/FzTdE5NeYHITqWugvcpLPGPNw9rrcOjMYA45J3nQnq4nbsB
vbS5U93w4PFWWQjG1T/N7HMQgXvmk+JLBZKzr1eLnylYM9AUP8ivneABhZntucWr
Nbuxoy/ZJJ1DjF2DqsNWlZA9OETu+DlEoTSkQpBFqPCmdW0AwwSLT6phJp7rGqvB
Jbjviy/imioijA8D6qHRFOyCP2vtCbGEzjd2TaRPhlCiCtndneOcOLmP4l3Xjby8
x8+KS8AojcT6mlNEeTlnwVk6Pf2rCQLRCX9xfTLJSkTGNdm7WbmpBHbIt1ixr/7i
RC3tGrch05lFOweGS0ufuaypL29GAM/xBNOirM+FNEi0ndKb5pQCpkWnW2iE/kvN
3Hc6slFitKcl0yxg7JcfNrDQXDiyrRbwwTs4rd0AaQHNecZLjU5ixKFX/c8lxzEZ
NiZFpg7HnM5scoyG3qaNoDS8j5wBOhyHjFE3Xcg7nE2AlhmJ31vkPCaF2vZK6hU1
TYOzJqj+gKsAaFWMWjO9yFJ1mC+sXNGp9J62Ico7/rve242HoDn7q5ZwnEUgc83b
v4o00gW66wQkF25PIVkod+PbDc2LkWJZee0iggAlc/G6bQojs7jmXiTQsdb3iR5h
W5wwk9ZXMdM5oEgx9cg9L8UPNGt0hqlT2hoomZJflOoLn7hXwf6B1y8GOg7K1dG9
HQZSLKOWLmGa7urEm3u0Br4y37dYcCxngj/NEEItCcV9NNUV0Dg4KP7HHjZQdWuh
Uw5xkNcel69gVBD4Uq4Ojpv/dFCw7Nq2C5lEBnyaycMH6AkZwC0Qh/LNYhvg68FY
uW1zv0H/GTKinyCuFATlbUAw9XDe4qq9OjZuwYe5Tde7WzO8uoxCAv9olJ+hQ1/e
1AIMbHW0F3r3VNcaKe6wp9z0MQSMD8qKxvlADhMr8T+ULKoCaQwJbG7oV8wGk83W
rc5cH5hoHjNg3cJ+3ARLCn5TD7OVPUISvCR/aOmVJoIhw/MxZ0Jt6A1Bp2YaH5eu
N2J1YeRqJnjenvc1l9nDRYFV5s9Rjv3TFkqp3h2MUsd/ouNiWuRdXTE/YgREpnEp
2IyOZ8FddHYQbCc5C7d6unsvh7r4TXYPIgzgQ7QBfgeYhR5khdcU2CGJ9piuzgqe
3Y2KEU5TTGswEMrbB2XgQkQWHh3LFnv6u+KGGrBdMhTSGYnwg22HViL1Y1gv2T+v
KIbTpwVn86OCZ1G7p7I+0CxQR9aN8c+v7Z7MVyDGCp8tQGzfNmLgmyIN7sQDH2ji
JZrL25irTfhuKQDKhn+xRFLx/+J05dY3fgKpMFeDIxFrF/2WcAgScrCja/Qzo/9E
S7F853QXIksPJ4y9i+0rW3RypUttprQyLLzG4Q17AIVU0d6OJWIqzzDxZYdOICDE
PnQCD7eVwVgcJ/OlP9lMoVNuvPSzpNEWeqs9z1i4Gi4BmtCGSlc5YwGO0PibrdQx
V4OkR8mScel7749bw2yhAxhcUqXJ/0UEx7gGTtnveyoeXdjBDaeETNGm5cJIic7/
+jY3PIvVzz6h5sOoi6awFJWzvWQntnKdHbu2n/Yf18LaHxiGlw1EGTEuwZl+Z7/s
uHPgrfbS8E4AVeQxmMb27XWbGIEwx48IM9QhT0H7NYBO/U4QZR5DkKGuCHedilN8
R3bjIP0mHBy5QBgApUGhVwjzbBbWmtLnTTK3eIg5ccG9ZqsLQCBXWyvJu9KVuk9+
gMWiA2BGP04EgPkq8muryTeGYQ9XyON6iAthsUuAdSpzZ6Dlxgb8NlcJJ0HcwyZy
+Yz5gz58YR8mUZWAySD1tmDUnKQEwGmCkqUHQMfCU6XmOfipDIynBkugEnL5VoVx
BMmnLtfe887WdEUd0iY3A/0524py3L17Fc/Rc0VyZE2ISDcjWubJVKQPinvCoQ2i
`protect END_PROTECTED
