`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvwIXCesXRcEhlJz4p0pCpPYFhakPAiW4QBjGSV82N4nEz+kUMRJkwpv5GwE3YQh
v6r2C6Ks2zivjsIC1UpV2Z1meIfpuC3KW1N1MiBfecyNj6V5Lj3l2vtda+gpz2wA
AKnWF9siPYjoVj4hcB33Fh6ceN2MhhaoACA6UD/fgAbbUVwVbgzob/cOMyuKyKH7
5/laLw+puEuZjK4jjOv6BdRaRZVrYX9qSLLv5BBn7jJqmMsm2wERdDhavt/g1UQt
nKzBXEK81t5Tguz+j5oYx8a64PvLRy141ddPEB2shQBkj7Zs6H6NKK0YmQ0QcDNo
CAee2KFjOKwKxVn46Y+PXF0zlnLeCxFSgZhoSn3qOT/nKUjUM6BSc+ANvaZ28TxC
My6RrbbjBr+ZvrMIR5Qt0lQ95GudXegMbhz/ERtDe3M=
`protect END_PROTECTED
