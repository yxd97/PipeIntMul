`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWQYdtLt5v5QW3EJ+sK9C0QGBAF3D+FtIiiVC9hDlTqlQj2J/MW2Urc7apSXWyrJ
yD7ePVK569NW67goNSW4fBN7C5f193ePTIpsA5+rquTgg/URNODWtphHQ0T0WLkd
4YqGdlMFOhqvh45hlDsHsHhSPXVL6HxZ0OmTWZ7tB8GeUHJMUfWgxrXbnuK7mwIH
dCkdGN0noDDAzXVocrItrDd2MJdfdPREOWiotcMKkrXUqSNTZNfKausFLX+iIXLx
pNdZ2r+9aifQBeBh9OM/+kLUYWagzuX1sJfmkjhie/K3v8ZU/9tlKPNpceW2wLUc
tmVYkw/YJI4EgNNEEObRMCDdVjBZOaaIZAQbN1CpQt31PzycGqchVF+R5KeGsIb0
Xeu5X3ijEDSeeXDFOvEH3Q==
`protect END_PROTECTED
