`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ldnKTj69N8mWqsec2cDux9on98Ytf9YrNmrb4qTu4jPJLPtbI8uG0DX2DOybZx0u
fK+d/5GmPpfCU33mQk2b8I/b1Miyf2zZm428gDn4zRBNfX4IKPHSjwBJvG3hzh96
hb7UZxG+3DP11wt1L6+XIX0WAI0hM0bMI8cPXLw8BjEoTqVhCvMqG6BPeXiCL723
DBk8HtLGnB+ZQVRWu/2BjmdD34ZLAWoDSju+7a21jTyeqHN0d6FPzUddIrRGBg9+
2hLWh/vShtoltMuaBa7fHGXP1U+1ywLJo/G9f+iVJHHiULiNP30c0Bqekage4Pux
Y/OxyxEmnLf+OrlgEHPn+PUbx4IYZL6BOEtANiP+rwAmnmtJPxPrpCiAnCWw4TdA
hWVBRgKgPqbXxB7kWk1xmvb7pzRexE/O2ngVYLkHckBRIh6larMJc5Pz0bHX9yXr
rpaA/ZFnfVylcIavcjHDaYQjz2B10NvdXhlSRaZTb/NUd/ijl8chSpRnuECF2Gam
tn0JVhC4TMXKaBUMwnwY5a5tZHRsXI9E+gyNoPoZqHp5gvX9yan6oBD+1kqUoLEu
F//b83zoY1JjZP/3u9BkppI1pXli/YKzglZNWmCsnuLcp+iEhk3L7zZmd4Okc3xY
jLsHqWoRIcSCQUj6MQj/UeSZHV9JonKB+z2lFHLe8VyQdCJpunrYO0PV9MIU3u61
eoCljRZA9s+O2jH4zBeq/+SG2UKGVHHL5rTfCq/+eDpjqJXsy3Vz83BuOTPDSp53
B+3u/iK/BzwVL7USD4if59f8wlVF6q5iw8Y9St/YSFyzNpZkBVmnYtDMIkwEqQTB
iw3wx6ptwdfB4QM15UX2SxyWy2HqHmhSth1J+X6qNQTxbpZ1yr+m5ycRnpx6xBh3
007C6XMGR4xIu09of7uSEOBvyC2mp2Z6HtE3rtzivIkJwi6tTUKFDdMFQE0gUCh+
V6szkbMtX6dReEVne5EJ70Q/pqGZBGU2HXsoxRWy3UKYuL+rcBQCLW7HuHnK+KPG
hNiY95Fg5pYsmsgI0OWPfmEbM5tZYtIKH9U7YE5A1apbog+3IxeYsy3R/bzr59MS
CITmSiaDjZoTm7Fk/jLd+o1tvoKfIXv25bUGoNl1tAG7nEkxs4G4ekSRw1IISysQ
CBtK76zH0IE/QWdTV2khCof3Z6J2ktb6k4o4e6GOpu7WqN+EBLaI+FX9K6Q5l92v
iGqqeMcwY5itYrizJM88uLYGOWsBTwfT+FcpPjd/yA/+utHuZCUeMAi/HLL2IXFa
pSLANHaHUi7HLo06TTz9EwdzRL/MUPfaxpsw4z5GOo9WtiISTwGVL9vGJynAoSY4
MTKOrVgTUWkYqu6/MyuJYMdD4HMdyQtJxrqZIno/welNIGIsi/FRWGg7jUylL57U
OaqomxvO+TMpGUX2kgcrYkYHhDr8fI+1f7MrMWFZvbpEuGEqBUWT8IkYdNpnt/VX
m+t5+8PyAdHxZbgLPBB/Pm5U5JngH3j/XcrsJ9X+rfvP95ddznU2wP6OPkndsfyX
jwwbuOklgcfNVOpuF6rhBJGhYpopTkfFf/r87THF6+doYxQHRlnFUcoRvofVbyzl
ylxE9STjk9hOqMgL86Aghns6MI0DPith1qGPWU4pM1gqEqoy5Bv1M+Gi5zYvNuJ+
vYQA1HhJoKGrG6XXvWXe8mGV3PFrOd9N1WjWottPjllJtsv252+6H6GLiDEFoxSf
tDcWyfzz+pIzCpJKjgHtskbBduv3pglImIKfoJQm+Ig0fVkkmygDSM0VuSD4+wFY
Ng0OoqPSLvieQZbyqWmxbt1WftLV0meyB7OkDlnXdyc8M2YaPhdEdKQgXFS6raAx
1+HcOpW8+ZNe+WLKSQLi8MdF96DBYTaMFgWc1q0Ug8lBxIYmEq7osZK8/hLPm6ZF
V+iaZVlN0DBY5dEn94skFUE9Z69uKyej2+/v+WyZu5yRnSzymXvzfcAzmtZUi/3r
NRNFNQmVpGNpXAibirwTk5Z3UuMAfVQTZQRro43fA3ULX/CTknmU8bi/TA0xR0nE
ZWDRiav4UrFaQhs7mJvRo7wzxeVMyxNDc5U13SizfJT/iEbjtsxi0uch6dR1g2QY
A3Kehf3/AeM+35fuEbejz6u7dtKaPEocTQYItYmU/fFiIWQjpRVza3moq2+/zYfA
7XaTvqH7B8C5+FbKK8K7ZQdgHozx+Sc4JpN3YyBNJ/+u5AFg3XvpBK0FEDTlLb0F
zmXA/rR7GwP2X8RBuoc0WZgeFNRV4MSoIGsSSWuaf1ExPROD719nAJwscrMIvp8C
PMPwqPG/hWfiyBe/+gUY0LkBQ0F1u+eV5eY6fmM5dO8J81CkuW2Ko+dwiudrZW77
FaQf/Ru1kazfiEB234umOmiuIX4WsaeMxpuiCj9PPlBqZGwzjU5uI+MHwtZITd6o
G4srrZGmJscLcG+MTN4s+lBFDI2wkoWgE/IiRmrXzSaR35beYreh1VmH2VjycbXe
+K2qUqwL73+uJg7IiHQKCEg/S5T6naKZnsfX5/gm83SlijKHctiZaivs4PX4iUZX
+vgfFIDcBQPkiO1Lh7Xm9TYHXqJcF6TLqh+/lapGns4tlzo/3qxbpZF7diNoOnKa
IuDbzQaZQkjIBqtBGWuGRiBfsR5SRSAQ0XuYcvFxbrssMaHYxbpHuTkaatttgKni
TaVHWRWQ4//9LYPYVH1cVKb4k/+JdeDYvFmA7I9f92a/ZxutN6s9SlSqAlde61ch
PCuOJ2T83ZoJ501kVZFtQ++5knn+EsgPwe3bv4empJup5HfI7OKjd9N64Hy2hbUW
ualsd22RVaxTgt8MinNW0lAsK/Ea8gn91Mie44md69LTVgWOH3LWvqbB6Hxn8gvP
x0vgQr2ZdtNGLgyyzRM+TXYqDfwihPQA8vAvThS23v2zx8tvr8mzvbc2Pg9wMTeL
F8g6jpadjAuMq3PevNoxJcxmz9k9BmRGlgEoD0tlXzQmPnAd3e6F2J+eD7oNaB4h
TbCwAT9jNf737/1ua3MembHKG7U49ZEvzPwxyEb8aTTgmY5KtkYr+x2sI/ZXsIMf
xHE7AQ8tY6tEcHwa/ugM1QI1wVow3UtUKRq93c+n/OXlkpT6HRKXMhuCaZbux+HS
0HztWpZZulCJQ13ZI+PAYUDAwACTmveW3X8AzitUOLSmRl0rJrX/8w2b/XV2p2Fu
h6N0oP8JAslGXJLuosmf2Q3yP+Qfzu+Y1gpD1YQL8HC915VJkNEgTi+KJlvDtqoS
A+ZjfPio3DRs84D8Zu3YDwoYQHSy1QkGF5+VY1AOXLFCOFr+kbLQuip7Z3vrMYfb
7cBnTuSEtVQOFEkUunRtVgYwQrzwoH/Q9uIr5NEnSAuDz9R/V6jtx31NtWtrv4hV
ry/4pJKmB32uWypcphQhKaO02VZrj1/nXVA52n42KulvFuIZuP5NP9fw+5k1CLcG
uQfa/jEgAzzCBYAF2hOwRme9wCAdWkFQoz3ZqEsWAULayG4tjKj5/R049+TQcilo
4zmXySmCC/IKDGE+tGjieHa0lu4xAfLEycNNT3XXqxtvZtALw6zub7fK2pnqMAfT
qRAFpjPpxvtoP0+x+pScB+n3RGQBNK4l1W7JOaJ69YwrNYz640KNFalDr5ruaH+L
PZPumwqaVbeKY8rE+VraD3tsLgg+k2CRPYS0p7ia2/sZHr/KiDlDzsdz/SsX6R5m
pmDHD/O3kbvyVOTypvomhcaEDER1p8HMGAYEVhgDZyJesfEmyGYw3j4ds0ONa1NJ
W/AwVGbjXeIT76eR8WI/DqHqulAt83M7SKReSapuhHtdrlPghn7e3+arQnJa3B1E
/uCpww5Ixa72zu1KM1m7Po03bxFQZWdS+CWelpIDa5x4uj4SH0mVBqGMBPS5Oyuw
I6iqcihea18TcbYnvehiIfjNXBlGvO+ws0nK7oXad4uKP5/7zygoh+zSJX+Au8+C
bRdMyUAfEXV0Mxwhh7mnm3eR6ZjdTQRzOW1xDnialBZB+fWRmPXy4lTqtbKE+1NM
OOIG8/JCkwoXGi+gT9p2Y6uzVQVyH9HuwL6/Brb13Dj5lDYBTRQDN/SmFijYt8G2
ImhkNyMBih4uGtevWB87E91rPOKsMKbOUQ7FhYGY+shexWBfPTA6aHLzq3XwIcFi
nfOC4GufZum4riRUi2j559eTu1H/3cra4K3N/umiBp8X0+JLrQaLeP8qGu9krW7E
8ATcqXWjzUQJ4MofiGMhWkR0NbcqIn55dqj/5S1KeyWateGkipQ1RjylNMWltmXX
q8T9qiO494K6bk+a4GV0q0rwBbg0tq2yzmtAdicwDgHMvZA/y6hvU74ZyoYlT+M9
MYydG/pGZVRQHl1R9UnokbL5jbfRVm5lnoTXt/rTVJLf/ssRI46ZsMHLZHWU/AMM
Wgu0UF2mrJxkjQp7OgGcaXjtKm7L9j6FFJ3bIlw/4kHVm97/xRM3265xZigcBIdP
7mu+HjKwGBk1GG7wg7bBl7xhC58E74y/ka99wnEk7EWS3awEp/8ddWpH1Ll76geE
46IxsKRfMLyOgAkuJmeM9YV/J6JcKHROoDVN6Ezvo9DT511f8yrZaHTtFA9dskZy
HMhcPmTYjp+XMyQwkcZdnBK4nHT4EUfylI5cD2rQIEB1O7f5mDPX5rhizNEwOUGy
Sd7r+U0mITCLq+d4VoziAFhvO//GtrY9drAN1r3V/WDhKU4VaQqXaagHgscvqH6/
TQX/H3RxS2st9TaQtuhAIafIDeJKmDGpazvqcNxMklNxLcJ44k/nbip2sFjqkIc3
1Tod5MoB30NoEBxMZAlg1QCpgnYIWaBY+SF1yygPsXQG+Fky0ayJQwj1eSzj15Rm
kI7GyxRoLoDNIQj3mg1c/AN3RB3hGhek1ypvR3AczeAQnHCsOfzcipgSqTr5CXph
Zhx//CDiTEPwwpphDCqu3e7xI77wQY5VQFSPiUxcUDLyyB0E5U6/JeQPCkp8PYog
80RDYpfNU1yrTmESFTzPy5K09Wu6SooAYEcDEWOjmaVlb90KGXKmeURGh/tlFarZ
iIdF/YmwFwF3+6+nAc6N6qX+bJ2DAMGw8bLgSa+iEjNZ8toJpIOYiI/igqT81fIy
n6s57vE1x949lRB1eJEawr14VrekazW6hihK8dRahgqXxf37omM8QgQACjiUFHAv
Cyqui1lt4JhA0eS/P0SwJcltEhojhsE4qRvAaZRLsF9V5DGWaDvU7764tuyKEAk9
o9cGE6fWlLsOnWcsFC75AgtJuAin9/lzxbCxqmvL3StvrKmX9DnGWfgXXbfKAzl1
MoA6YA67EuewuLJwk8JEok2q4SHdMqgg1ETTrC8yLSeCb7GevrulmA58GIX2oy3+
NrfavUS/0u6fEcwI2ACwqov3H0yOg077iXJNjzf+CKMWUAhqhdlnDug01MPq5en2
/+ddzlCLgXwq7pFm5XT+i6hoxcEwFBBycIShq+BqPI/0iuvo6j2FDC2kZReWx4vS
Te5PGRuC+4RcPLemunPCc3qVMN6rNwaCjdOJ7rs8pLXFxjF6qHE+3qLwa4svWQ6X
QXhfs2dyUh9qv3bI0yH+ZFbY6cYT0EMTfm1l9luv7NfHdsO40BBukeaHRyT1dY5o
Mw9AfrRA8tytSdYyhrpeW/8gm0Ijag17Dr/JF9Fb1vCGASPZg2E5zM8r0It7jqri
X/ky+5n54Xfr+xVFzzVSNC9DbaJW+wuLOsWhCqW1PrgWmV7QCcpWpZM5ecn6vOCG
q+2OWyidMbWmoYdD3KCYWh10mejrsiYKUDMD2DwHW9rwrnSvJGL/4Xlg2ohUtWt3
8lJiTX9cIIDAhHz5noYqVf0/5dw3z2gZYWcIMamMVlaqtoGKFJxx8cBi0Jf6La6h
U1X4pSCT9clWmwQ19AEu/YBdv9w5lPaxCBZp/Zg+gFdO/rRMT15TrWWjSfP6S/Xw
0TttZw7tx1aSsFqwfB1YMHbrrDGjrlnCrJyC2n0uyzMAH7k1kUs3Ww1hO2GOpdRz
fXDAIxmhyMtSMXO9xfE3J6g923849io2T6Z3Q1cBc9iihp5E/6ZrDxW+/6H77L/h
KEJO0ziWyzdsNEJYhdHmqkuRA42Vty+b0Da5U+vNAEw16ga0qTppusesv98dOsib
WcUfm25Xh2+6HHo/Nr0/ejyPatRYDPKQsGMa3vnEVasCBxJMjodHJG6s2vDXiPIb
wC3eQUcKjOM64Hr3cDZNH0ATbzqjUpWO/rTjm3f6Ak7Zhof+kJHQFTP1JYF2VBKQ
Ovj5H6NBH4N/CI3WyPScJoBsBqlpDkvIMv38U36aPhJsdFJvyDwpfkX5YzbRNH1f
vNSBxsMzxO3dbl8KosT4/9T7GlqqRZCfUSALB1FgctcLDkwif0aIMY1FAQQ4Sd5h
aqqh+GbxxjV7RX1uUw7T9m4WvJj3vD5OotFN2PKykO841KRk4Z2ciQT0mCAFBsin
hd6pt10+1ain9qE3Y4SZCEJq24BrwhIMBUDLK2yCyj6rC7hiqbCu8yPMPcqmeWrR
V0ak5/iZW23Ol4vKeRpO24KqyNSlbWcLrLOB3r6MwXgKY6evUYP8+qUynOw6XNQY
Y8fKt5FmIpaogUtxI4Fqp7nOqOGgPawQ/CUfk3sA+mdxfvGFTq6RugIvJ+4Tt1ZI
S0Z8+fEYDQ23Doovxft2bXCgE/+KHEQO/auKcKmBeyk3v7ELLG9POfSwmiAcM0C+
Pb9gY0c9wMRNixlRu+rYD1/43M/s5JyJfmwzQsdMu1d0PsdwF9ZY6mi8nhZzwPDQ
kGCmUquZY0L3Yrf6iU8WUbDgPRfoaEMQj63qV8J1JDMxsRt04FWXwsUNUuGvDjew
h2wThoXHeeCGWKfIx0DlLEPl0IgEj3Y68i3fZeG2vvFvbkV1Nj1a1D1AO+6HbksU
26KgOHsIB+bKiBcF70DVep4uRkb27owejQZI9iYNRDBEVuutn+cryiOtYkBeTICx
b8Esp3VehPA1BI75ckOrAmIjuWSKAS9VrxZz5O3PiY5AS6ma20hb14Udjd8aetVy
bW2MpfmPMQaUL4SLi+yIv97LDktU8sSDph9dgZ+a5NC93XjU6H0qf34ROHehAjpv
JvH+iodOFlZfinQE5T61myKdDauZqs+h5K2SgJKzwHipso75sClQ8rQWeFd281r7
Fqc3NvUyn5/X/KyIGnSRXRhBC8qVH14mPf2EGnldReNCqF+HS5Hhv+xzTK/zeV8a
oKfna+F6+/oYBlL8zDQuyOw8mrA418OGihwy4kJLPSSwBqVOGu7aN+APT08CJkRq
Sh40/on9mKzHZ+o1CkYr3rL+1Sk+lvAQbKqUgJLo9Opvg8DiZSM3AUu8nc0Ku9zm
OQ+Obmunhup3fSFY+x5nvBmYpTWBIUgaRSJQ9C7B2VYmFGdCEKRghlfx3yMQRCsT
tCvOAgawfJAozFeujG71pTnersr42bvUWpriHq0+Fyvk+LeuS9JP9wOMgm0ASw0J
3QKp8s/OzbS8J8uAKiFQT8mBxiIBDNWcSDwl7EDJ6o0v8vx2azX7Pdq1VqOmAg+z
g5RPiZKbw8pR4VilcDirQ++uM1G9qThVXKmuqJGTlPe3dyfzjxVpTcAwWW5/1xxW
JJOTqzcpn7FtK2akwZo6OVP2eLC4zG2wozJIVqOURN/EjF3aWOO86DbvM1rmpvN6
i0S1Xy2tj5nkbC4g3bYYF2NTjYqf47L6lzkD/Lq8IFr7dB1V8393HplqDOKnnEwa
5rvBSNvsRGTt/X+yDDt9U1U5Z5fx7d6xT1fjm/0Tjzcotul3I5acbEotAlC0N5z4
GO2CPn+u4zYLDn/0HVuczV6m7QTCA58JMRt0UZR1/cyJ/QqddC5oRNZg1/qhng2U
bSIhpH4oWjeYnVG0s0vUbbrMo/CxIWwrr2vJSXsBuYqwYrO9xd1Sh4KlyuaA7jm7
KXs6F46AuUuOAo08GvGE6ihWHcFbHGnjY7PJhDg35m91x4EIYEoB4GF8KqopPwlz
HONHtLptXqBQXh57prpAN2iE51bz0irzIYjgZm0SPvfs5PafsO1IYS6motdGl7Z+
z9lYuWM0OSWcckROfj4UMESu2lY+38KNwTCVtZWFhR0=
`protect END_PROTECTED
