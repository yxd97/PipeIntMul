`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JKAepVbFy5BYHRhdT90BfMaZGBqc6TA1nI1ydLIZH3W6VGitddeb/GzaGlLVtpAy
tJ1SZmk+WnMFkL0Esu+Hf8Gjcb1gl4mSJXl0WhDNbt3++J87UK+XwM5PS6wOkQH1
xAGRodLWOBlO3kwZu+nTl6k/5/9bQbm0FB5xuctHjd81ALofZU5/M7O3TjlUX8Jl
mSTOadf3gDyda6kEaXUB937HEerv7t5nnXZFkVVfHeOSReVDd0WiFryPjI+zVq8f
JbV7njA23pzyxhn6Gl3qWPVSTTZnPbfI+EgEa0DjPyYEQKRBH22CKziMwQy+OCyw
yrxrCIonIOokKVMLHl/E2uAuBuo0nFzfo5m90FFfNtTWmrLFQ9B5nPchTEYnBB/d
FQSRAz74auYCIw+b6RVLiwersGQdUZ9bES2M1LS5l5xGzr8QQOCU8fVt/zDKq1tS
47w7M9SO5KLgYmqaW6wCMBEwHc5MyY7HVtkM23buIWAU4T8MobZl6Qob3Th9J1NX
Qjsfv1GqjuDZzH5RTXgqXKwK4Fs6RSKGeqprU4Tm66GSd9bilK32YNvE1M/VUAvR
5CqAO3Fi/aOINorcZKy2fQ==
`protect END_PROTECTED
