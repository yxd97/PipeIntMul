`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ctXvSymd61qirL4B/6isaxszoiH/vD1i49qmCRgDcsZQTNNHpF4s0WtQsUyVCbak
7mLrCN2ilgOkyEZzNOXTWVHgGCX2YOeS7BYUQEgMOgpGL7RSCeBpgR8Lo9luJl7B
ATQA9Nl8pVJ61v6mrpnmF6TxlywcXGhh6V8V9p5WBJ4I0zNfPdk/chUgv6KKo2Um
vMELBUpZ6qxc3QdIsGwD5oIjKwEh39bsWhiTMVNQkotSAMktXrU76gbm6twcdh0X
m021NiSNPzs6Kmg7QZUdk+zk611qovGpqfBJ55gKQnHiO4SUr2joUUx/Eu1zO8KO
530D7W4SFHstz/o63KobRw==
`protect END_PROTECTED
