`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZSf2payBS5kb7bMiffDqu64q02uQfx40nyHlpmGaaW55kYDIJeK0WoLpqBxAvee1
Rtd3bAmzK0o9QcnpEkLdr3ITDq767oUQ73C8ksgVqGW+zEPc2Y+4JGRorVEfsANV
Yh7oKRofL0QNwfu6hiyh0epKA9VpLd0BGcdvoj2QTY9YZTNu0HV6GGmvLkBpt3/A
gB2VqciRvjWcqFnelFOzj3S6MCqX1cSg1CgYgQu35BEuDd8xCOr1umF/7sm9w+oE
ucE2EmSlxbpxPSyscYsXNTAEVBsuNpJ5eJFSlm+J7SlPYgr4VYl5j5nYqeNdlfag
Ztk2iWNeH9tF0uIKK4ijDuIHvf9ndY0VSV8l6vtt+j0RCSLx3y1KJ4/neW7p1WFC
XpT96k9Hd303m/GorKjd+pG7TLJlbl8GE1m9gPMV6MysJo2ji7BVSeLOYh3qChCI
Rg4cQkk1dqTfTwxSv4aKpSrkwGG8E/jhPPHT2+w1YWCxiXvpXu6G9DseFG5vCmuh
y4i1nY6sj0+q8dmSn2XqgLBB0iRbzvaqA37D9zhISEvtDq1jHLBUo9Tm0fOaEamc
08ybQCjVcN7t+69ajWDASFHhDZMQwCbXyif4iQ81y9TkjuqZmJOFIaYDNlbLn4rn
eYHnmKfR0owEb/AkmmlaH5p20Spvj+tlscraFTPcLM2YdjyZEnq4xa9OlweyEjDe
bklRQxdUvH0IEiPKcLuaCqXvKY2OGmnoQABCANhVl+sdxRFVhUQfkRG+P/i2nqvb
iyrkMBlwFu8Qe/6jPdeBobJgcYDI5yCJvWKS4l8puWp5k7ZY7AuqLKLilVWmvBbD
DmgKWpzjA4YcfYkmL6k2+jgi5BrETEbBjx++434/becGHUJri3eEj3u+DL3C8LYy
JQ8d2mxXWCOXjshwj7Fb5HKq1rOXWXYo42GnDjVl0kiovLjvXzR68ZRNgzCqPue7
z1PgplHNApx1GiR2V21C/mYRyzFgJIw4UxjrGeqAh9wBwqVCb0NzdGLfrZWZ7qK7
pLz4TQ2qMTCrxqMchmmNShqmMmVtvZ4ys+8vQHmn9gAdJl4JIJiS17zU7SuMRcJL
rxPpIx7tqytd4/dqlvqkAgx+mDh4MYyngSxAG31L5aE/ZjmUS+ZF7+R9KMm88p7L
1F3dMV2jHMdHeHGMwTYIDME1lbLd7i4tFjwkAOR6cdWeO8YuT0kUfaGgRMQfWeiF
O8UhLkFPFDDuOKQ8Z3sn/YpbzagnkzEHzmlQaqcEggyGhp3K/Kaevr93CPvuXkFG
KhoGBHD74C2qNFUgpk11jEaMR7sL/2HGOCA691717fozaPEjzEGUAJjDFPYXmMIv
xoFJsnyFl9UZkc15q0inD7NAoRbKDpwgd2FNcatqtobOyNQiskCgGmyZAqH1ZBek
8UW5+WSSd4+ql58R5AEhNq4UfHQZmcL9t736SR9PhJrOn+mhbMnntT5vIJZZrdNe
lBgdbsQYw1NUZdp7sA46Ag+LSXmcgi/QUu0p3ZuRxTKAkY2VEc6lI1J0XB5o+zu1
NoZ/ZWCXh4F82hjH0NNphwBCuJ2XsbFmHnv660L46q707om8sFwKNXXkGBhDqXo0
n2ADTUXKQisWEcusMR+9VH/9G82KA17hdeh+ncSvHaakFaMGC0eGdjGiQv1v+jY8
H6BURrqbsI+eQfJRIqRYRfSNbc2Ol8T6z5qA+LKISHQPEZqbosLzTXkkqQQvqhod
uiHzfCVmVqLTCez7mXcvObXBEAtSpyet1LgXEXRxY3KoBdUCoO9kwnjXZjpZS/1v
3iUXs2yEw5Jko1o1h5+QVIwjpU7a1iSZTtGz8y/kF26NLlBY7+CXcl0UZk97VBRb
hwtGM9/lO9ARZG+fEZwISPt7xyY4xCJz1v8L9ME9G8xmaYEcx/oYs/683bu/9CIG
OI8SNp6Wx0/VQLSSJcP0kyR2rIZ9JKFTDs5Tibvtb7UEFmAa+PYiU7z52FWzsN+w
uYOHbGqb5ZIcQ+WlBKWjhEv8SyRj6YSzBHWVkk53XbLNEXB6CfIf67uWxXAZ0wP9
O4V5YaD9R3FNPyuvyS5Jd9u6GyPIbEUxpy9agjInaNFRRsW84hj2i5snzui1/HFr
U5UNIO30jl47tL9wbYiKMbVCUor/XE7FUZ0VKS1CRDrcdNKBrOJWJXN94BxG0mMC
C9b8eU0DabnV6Ew5O8+sD4Zk3GRPHcoV8owXfJYKjUB0aW6ZiycR1Vdhq9tPguir
GofAhu2ChaUC0gBkahWPFkI9dvdZIFsnsqtjFwXBD9fzQNOrsU3yDoNAHwcZMsD8
fNxUCyJDc7PfGK8x184iWTM8RFElHasdl1Qe1gXAG81o3FGFqJsBVKNHa89LIOAO
xv48KGpSEvhHWg6VPWE2XGfzWesWVJIkUipZUaeL3CU8YlCYZZJ5zZF/fqFU43aw
7C5RiXE3CD7zPkFVOylq1Mrw67wIq+wsfhZtVeMI3Io/1XySxpmsEZsk8M7TJVnV
eQskZ/BpcmkWCC43Gi5Es0XH5CKgOj+jW+YVPjMavwul28fB10MqriUGArNfFUiP
gKwkCdivU9z0+X1c4BEPanJn8xlny+wwoTN1CmPjzqI30KuPlf0pmhmCd5mGR54P
iZ6m5PQ79z/CSxr5BxGwsXrrVIf5lNcEMznqQohlsr7cbpEvASBMpBfatA7iCMWG
26KeK7EWuH9qeh+7ofGjZYLzttHY3kStCZ4PK40cLa3aFrqoGQFkcURgBqXmCygM
rTg/6ETHHxmqVrcm7L6x0oF74OXQW26zSRvJBO2y7DrmsdqVzjzGqLcHk7N1cSpT
K2xdZudNW4yrgW9ft9hWMulGOHLp3F1xPaIWCO5TO3hHC2D6HK+yEwPoZeqkdM9P
Lwo22tt4OtN9ii7cv0Wkb+AQ3blBe2/HQqgB0PntoO4JfAwAEpNAPYo3l1nSCWfk
giL7uoMotluSuYUPfuKB85yNVzmOF4OQzIlRRMnlbgStytMGc9ArhhXih68rT2fr
m4zMYspPAPaUHzZKaEjsMY+/+o+xUjQI1w+786HT/FGY4/XukWqKT/skx8IG94kY
7qE2GkKjIqs2J3A69OqfQX80Bk1qV0RtMloR4Ba0Cl+8uWcAQVxCls6shILg+gJb
eO9A7ibNdudhV2aYqYyEnP3M7MCpOJytg40/c+PSWLPcvJ7fq/lncD1BlsYYuZ4Z
Vo9lS4ma0vNe8MPoojYDuSOoc6vlWCLDEBbN/GYBVrz0ZrCc87fi0WwJoRH0x13y
px02ADpOEsZLYeeHGoYhpy9Vum/5+3VtIY+yCle96nPrSwMMIZbTMyyjtzUiqDTD
25aIjx+sWDZlX1NOAVbcGiJqGafIYG6JFvYMFrCzpUrdBWFshbPoiP4y5pGRPLpw
QTnE49SNcfwTBGVZrlkPQOQFDuGvBfSzAd8pempB8hB0wKPFfMmbyxhvWMhkV103
d2q89K/plPsG87Yfhai9qX1EqvLGPeD/3wi9VWr4zh9pEsAP1nqQBGNgrtyG6HUz
qOAwFG06y8URLoLYNuptLFaAMAeBWLgjg3FwUh0CTAY2M7jeOashYXe49trUdcTL
MCIsNX0/ME51lCUXdybjHpeQe+iE25XgeTuDoMwGHqU9FFK3qxjvj5BNmEagbQPc
LUVPMb+VLZZXEvTf0ZAMGHEPDFwsq/zWoSxaAHtUobRucWBRnd9BLbP0tploR9J7
Z7UKi36sis6nqGPbdMh+IAE9K/QjnC/+P+VInjAK7e3nXloHTdCPhOKVmO7hLQjZ
Rpsta+nTOr8y44dBk57Bvide6Itkn5iD3t6fNAkq65m/VCArtGApPI1MMaqDGHN9
XKPkhIXGbN3O7QKQF7N86MxYiM2CaI2REeW5Za1gPKTDo9wDXGzdIkGKisWBhlKT
IEEAct/IgVvxucOWfbPLSqDEm1DtqAIwi33MapjWr3lY003VyjcSeQ50gWYncM6P
ujrK1K+qLWU0GlExCz40PhaeEOTTNzJVYu2Nyv4hUPDfHv5AhqWM1NHoWhtFazSo
Xum/4yrd+/OaTu7onjCx9ot4Qz7h9cmkTUMhCUqhEW3SMPIOdfDx4DWAiBQOsGYb
rq9D5MDkIJDbvknldR36yq63Z1pgSwYBRg0ZiI9rJ0VB5EeHuBUs6lUaN4AFgGP6
Y7nuj7g7ys34I4wSyjqB9nHnVCGj8GBpdFST50rkeHs0SmlyKutdZWza/fJsTJog
mfDK23GT66blCnrqs2xxjQSOQwXVJgH/z+hllTqfg9bcPT9T6VvIYShveF6X6iI8
LBUx6ZAOVj4D6DtNRWjj3J+EM0Ktr/Kj6FHiZtU9LvRRA4+1SQGeWRyBpsFZNgz9
TtEupIRcV/KMrNXcF+Sx3kaEhwzGqN7XOLZWw4u4ZljsNN//Xzd5TKSNTkFGBByD
HVWVdj3sGYNUofTxiuv5CqP4xQWODd0MrUaeJG4CdKnRR3dqxr76HmyoHSJmx6Bf
bgXlGup/tLTDbMFENsgW7YJp3zAzkxyxFiSYkiuvJyoH4IljEHxBr2tXdWCnk59W
h4H6Zoc1Wv1GjozR+6NL3gvi2bUYLjevEfuN3MChCQGy8tGJ1/46nzC/3R1InsDx
irQPacJauF7tWUptfkUADFxOirx+K3xJP6kIFpTBueksY3PR5Vz9CvoD+Ax3hLwO
bzHBRlXKdhgIaI6T4La50fcYAENqpwA+9FnbNzpm7UphrUnWrZx0PYBYL/lCF9fG
s6o7Ti3q0M2Klpie/o2HKh6RK9clnWHISC5csQxRT3wtws+6QfCqHSBHsuYsxPg9
UV8lmk0pccTomaYZxlMzKejMuMycHdNqD5+rCzInbv3ji6LORvEz8TLRsN6o6FCe
2YunAM5749A12WtQ7j0tbh9XZd2fRaGcd0DRorKA58BfucSyRdqV1Ul8MCcInMZn
qjF9YD7u/zwcYm4Fda4vsWHBYIxpU4ddq9tcdNpQL4xgtJzFeY9WzOlQbdrB67kv
hNHGroFdKjWWaarz9XDGseCccOjoIyx5GZln3m/0pvNOmS7GI8n1aicKW85kJVmT
wb66L5NKIzRh7jLKlXLL+AoPDI8NfwObiH8nqjboQ1yHniCDpEeKpmxt/2OMB/Ck
siY+c7In3KnJ7lpqSVwKvzI72+94LtATjriPxaFQIcP5JS8q8IG1o70jOsRbxk2G
Ej/+zOaEyVxSUb4WswuAngrNSBUXhuYjVr0/dzuRGWiALxZiw+l05AfTWyMHBaFi
MGW1d1EaZb7mwkzY3sTPrYzrXdiwJfFZpy8YL1g3aY8oAoMoq+X1B4eAK1FAGMOA
m3Vts3x+JreBimS7b/qg/DEYrI/bi99O1qRqSlOkoMYMM+lLlGzpbNVszxSTml/3
YN8YueMQfukM93FBaVha4Y69oN/bPvThD3NWrP+7Ec8qE/sxMyVIem4yMX1enBHX
FCpgkU5LyHmNKtlYZ+M7I3UMtegTfsY73/Rv4XlJngMxUVAg7YZmNZsv0qIH6EoG
j3+asLycroxTvhW6xIjg32Rm6W++2pdXw3ZDk3Vnbdtds9vo9/SpdFv3G/PH57qg
kEmKcYJsFIOUSeB0xA9LT8gHW/j6SpzQ3Nbo0lcqXxZaowUJD10L5HIl0FVihsra
d6bct6yyV3+XknWBDn8nbNIwOUFYMJoAJJexFaudAkmmsvD0Rg7gJtprV5hqIv5H
GBUqcjbHd/yTQd/ZXjJuJ5TbbIUQIv8ka686QGPd4lwngZpPVGKK/LBLHwTyTkmI
SnUd5R/RzsYsYXamX8IG+3JbdpDtZ0Uu57CUUmbVLUZqGyhpqwBG1O8CrtUBaDeo
EB9CJBUrtHGH7zU7JpEFE3HgbmvWYTHlBZ/5Wollx16PTn3h+GPbgodklUq11mN6
BFAmKbuxIuy2QlYPCdRYTcU93ZLh2C7C+WXDbusA+7w2BEt6HPfOLp4uC+0pMa1p
HJ7ZOa7CnrkIZ+8v9vvudwFjODSnhv2mzr1id/VnMfynNn8sLrV9PHsflH5O7E8j
QEZEwPSyYGvsrCcxN1Js4zD35E3XFbhUZ1F9+ztQoU28LDI2GbhU2xwzFRCqmKPa
USTUH0FRlG8aBbvSoEg+htik/CoRJbp3UASaenHEqWkMobamgF0+iPvb4FVyJU3I
z3HQiPLA7F+6ArQMAsIFQL8ewPsvh8Fu5OAOYvxZQVNwKxL8KAZlvJOeZlZvp01W
LJ7MyWlmSwBbunfSPhwKT+D8Z5n121x+UeRbmlpPUZTWQXluEUSLlU5IWoe7UxfN
zSQUvwjtdONCCpuvFgGRGHP2s4jcytEIbB+eJG0htpfAwCJBlUJLY/zRoWaUatGL
nF4TF+DS0DdXfmfmnNWmcSeTwczk9ZSsR7E2PPpHepN54zp2z3scLpbWTQ5rZj2Q
oegOneOtQRLLbFJse+Wrqkr+GMO/ImvvqR5FI0TbF6ewzpAJknB7yChO9j1tyl2A
WjoonSNDFUFw7QzD20PvPwW3VTrJ6fh+mUm1fUvn29QDyKXCzLLDzOk87GBEAA+p
c248h/5PXiJpEDZYyf+QmQREojTViMEgM7kHreePQ0eNprSkUjhZlqD2Cl2KmRw6
cenEogmpXsaXEMN+qz82oM5MPJQX2yVoP7f6TIzR7hFPmHBhgsfZqDCcUuIdlv2B
ZTESJsFnqpyeye0cxlq5+LbuT/PNZ72VVrk+iSlboahqjfKhUsJ4WSxyDzB7vmSl
rhlYOnM5fJ4tdOWWzrm0qtm92VBcDnYz+xTPdemnDjaVUNOUZRw4zbeGCNq3fbfS
Lj0XMmu3bUwrnD749MZ7iwU+gu+zHVk7NQjHRMWpIwWpCG8Sd4/5y02fb93D+fUm
UVwQvp8s6Lv1Lde+fiaS37avK0H8KmMUBY693SiXuDAhGgsmY59oyhPV8XDhC1cJ
o33lPqflSDYHx8jUzoEqg+o2/++fO+IglfKBYTs1b4NZyJ9N/VqQR3Ujz5XeHDo0
tHVDx6+vJ6F3xQolXsKqt+K6WuHRpywLsH9ghw6Biw0o2eXpDn+ECQlP/Ao6fQ69
73NFRLseTZFVhVCqVysGM2HI7Vbz0ORSdb2bBjJ1yjDmrpbUdwBA51/MPmrozUvk
7cmb2DX7/S3eJajUMUUEz59bHT0J8Df6IKIapGYkO6yQp2suW5kO8V/Y1IDzPGQr
jSrN6hmuvS7s/Xovl+FSOhqZpWzn22oAGjID4Pix0e+M+55qqI9fQZmRtQn3LHM5
e+6lnw2kNsiXu90LXrt7ZqgavS8uM5Fgc0/M/tga7AKFSDO6Np26mA7D+5BGeacU
YZkftG848K+27vRAwSnRg5Cmll6GyA+xQilnheoaQjYULHf4vQLpH6qDS7u0b1Z9
TzmXLApYivR77NqMuL9Kbda6PXKkqS9jHHLcBEnCVJ0OVnUeVBocC3dSY6CiUX2l
PSxclWv5gVqAKRPKVLAPc+hoePGict3w7t3KYxYQbMM/k5SL9TLK3rJQ6pUl1kqu
uTgkwlGiydX4vrOZOYCKgEyIsdvVIm4OhdorIBDUEAaJNJd/Et6lK29OdJYp48Fd
ys+nc0OAQeC0iv9e+yY9qWPXNTDcNcXmDJEn5BTqvtgBEi7b3nxko01k9frePY/e
TXiaNm16S2zKmQoVcVVmYSj94noi797wN/DTKh756Cwzv8q7QnpAO7QVfMPgY2xJ
D3hVYvzDL+Pnc7HIcQPGkhA0pbfWMSAddBfI/CrWDBvj1nKpAFWi3RjIp1hqM61P
daKZH0c3B1aRVKdNN4eDuLd6WpoCM4mMe3mIp6St+YSyvAL0D2alNNUciucXVkHi
48LetBzNh06AQmw904xRH4cohvJbGKM1za+wMOnnPFhxsPCM8WaLBSxwhhP+EhWs
EErI8f+i/4Tm32jkmI/YhINUfey3rsPTRMiW8YlODeRt31mZNML0A42n6gzW4t31
0yiCXAPQhKnbk91AJLAJmaiMZgm+apPpBIrWTVbnjhhZyLsYVxU1HzcxHaSiNhFJ
9UuP5LBiusN7kKBnXj0fwdKm6wBS/n/X5tcXa/eDS0Z4Dq+VoUrOfMC4OT65Yb86
BTeBBPYBEkFtovP85KMwersS/msLmM0/kIxYL8WS6nc763nLADc7sMxXm3DHH14/
yh8leAJYjmAUiQM5MtV9jOu3PI8t2o8ia2u9pIdlKC6xA/VdY8nYVahIJ2LgHe6l
UlJP+/1s2EtlqxwAnLUmn7A+ft5BTc/L7cVo+AAxxiIgws6SuP2sgEZb0qdojsdK
TDH1uhJnq2nBifw90mRrbZ5L55S1af/CR0n+4LjbP4VeVPxpTKLD9Pgh9d8xSOe/
1SgvcjSuQhVQsUAoStp0Ri/pV/KiYQcXz8ecZ+6HRizA9q1OGQ+XPZzPmlLcr6wW
KDNlbBfXlenN9cxLBrqJn2rjTz7DRLMKXs8JRHHQqhURof/iE9wupDH6qWGNqEdy
zjtvXTKr2rOteJ8cCbWrSUijgL7O0BnJY5g0XbIAdovhObEFB914M0vhhQ20qP0b
Ls0jcljB6M2KmU9H+qgrQX1pWOb4PkUF+MZ/TVXWrZBZrs87JD91blnP6/fwDccV
j+80ZEbLfNwXEftxOMCk5B1mfOCKAzzLxElxu1PytN0gni8sddttIJXKwMoYNnsn
RBIa97z2OowuKUWPoSYyW6lqEVYdtZdCYe9ntRFHEPHp7fgN1uThBlQo/0CVTjxS
I4PhF1Y5pHYt4mitsH8kYAjFvaHwVv9h68PoTQe/zW2l05MZ5NUtnbYDSxF7vJ8b
f07Hmi0UFwpOnHi92JeH6Ebs9ovHRa8qjRDCCUMF7F5yiEXK0Fxu7xXuHOMwE2BH
F3i/Hvfn0PldiiyjiQM+7jR6EFKFonmTr3dWluycEUhtVt3u+DpXENOB9L0OvNHm
N8dwobIRXZK8XWSzD6XeZ8IYP956Bhe+rhJPKNV6gKSclGCqGOLOwgneadUVM8tU
A/3Zm/IHsX5nyqbwAPckWtSiGq8tUAWo1hKHNdsqfJNBSKmwgrFVCrdPNhTqIztQ
+VmS+M/W5Y4B1MRA9PJ5dL9+BsWESxavPY6zszJ3l4HffJ5+KLQ6CEbMH+/0ntd+
C+QAJuZEtdOpWlG+wzQE4Jfsd/lOkhjq1P7ixS9VTLzu6F2TE5Ob28Qd8ar9ekPA
zj5SnIGJQzuIpnpE3WyMVXrG5VeaZ5Fb/0WILtvQ5qjOTXk5SQlEeKwhW5O+zv7B
Z7BQQ2f8ss/X8LD6zB6NXW0k7OjJBjevnF5jcxpmPAf/dui/ueTKypT550v5f2as
tiEhXJPpXNnXCJxVcpz/FgVU5yeQGLQTL+BjlxOdsjuXqfO3VWLMKP8cQL0WRJ2i
P2J1bjX7m7CDVivUDHxgHpNK3EXBwZHcz780A4Ifs/SkWhXEMJtjeZm/LfhnK/VT
mDgcabAxTOr42g1ujreJA/tPYvB5l/7dAHQ8dgZoEiHEJuGoLsMAhl8YoAApSuUp
/yLCoV7kKGpVLqnMl3tlG6dsn6dnQp46oMJLV0SyIKznjoqSKTAzIKxWLE3Od5n0
VL/MoCVqBZzpP8RR+mG97hZe+u5tAbnO/nlBZ4KO192ss86RyVjN8Xvx/zhwZTi3
kcO16DzuYenmJVGD82ehJKo3vIrCDKDLZrosHcJaqKLZ5GMFFgxmcSPejUjyQrup
+I4GRvQssUtlbi+VAaXXc0BhBibW7ACszmOeNI2s47Zqn3g5ggeck67OcLFUIruw
Pa6nrsNSK0QKnZgRzZNhslEBhr45OIHQfjqf5OGGIOcAfolWXkNOFvEWQi10jk+z
BXG4uGP78j/qpUqzJ4PAE+6MVFwGbklx2MNgf9B3y24JTe+Psm1Df+AhDWmstFc5
2TzryrK8YwUpP94nerrMH3+M710XJcQVLTnLx/TL5O7ToIn1Cu6ob4pVYJBYTxsR
NeG+4Z31pe7wSNUGM5W9KDvquHAOqDXQ/LoCfqhPoAU/uWKgXSRT8FCNeWDeMCmm
7AXHT5DJk8E/3YQMTKs0+iWmVIbQpXW4WDHXmO7W7kr2FoZdAJn0PAFrMNH6YB7W
u1wMAAWvfgvk+bahnFGsa9EiZ3AD/wv2U9MAWUwzmkd9Ip0LbEiybGtFay1w39dY
tsTVSZbqqIPuZctj6lVBpZdPFyFVpwbnqyxocDiGAJqjsS8w1xRFL7DSbg06qq5m
yqKxYUKzY9rsriBI+yXHY3lyfEpOi3BHTWD+vjAjEu/PjdZomtnb7LbZCVtZdreg
QCOe7Ckg7FmTCnmL2zr958Rfezg2tajFeE/1Tbnbr3cavCW5dvAaNx0+ISxTw+3P
oonA2wEDnBMD4UWuGdahEOP/TpZTIFEFmLBbADdziz4xF94QmXQIfy3GsMLoQ8Gj
HlGRwU71yGX1Zr+bnY0inxxzkV2GTiiWJmeeiRDpRvq5Xrp6u7q/Dh0lYlCD6S7w
PWMTY5oqay8el1tIjy2FWtxRTOjisFQZ5xSaUcL7wwbOgE+CJiRwV9uTeEu5W0Ab
/oXio0ZDF6raRNt5UWcjlFu/ds/sOL6fUPvDlCc+92au6lsiClbL5+0QL7KMVmEY
tiuZ/YZRYFjhFRlYF24UDzlkXKNocP8VIXiRgQXjsYz31XrxySrU7jQWPPXqdDPp
O3C+y1wg5AvZe8eG/XFSIckQatcr0NhIusztJ/EdOeEE4VRn37aS/xcXG4ezSqn1
2+7l8OuFaGNwBqsseY2hA1CQ1Rh8Z9LhqZYu6mkbk6MXu9tirIkfBjuUiQ91AMWY
sPwKJQ0YIsRksopDHhUGVOGrzm6ONzx/DFR5AcIlQF/J1iuAyZ251jMNDBnYstzt
0UERvGslQGKljNOqECKhdqgOPO4elpUPfnla3tjjxHMtJ1zJAIqRBeAy3HTIzzrG
fFPccSmAyNkTnjUu7cpIED8mwNcGITsY6Rx4Ra1Dsqq3Dw/41PlOwBvrfYzteFWU
Z2FSSOFKsHza5dLSW6veEydtjtgP3e6YjXBLldLfsXHc5NY+VlbxQ+NvqEwLkl/H
xjBB8oGztjLP1SpJv+v/VrqXmGVaS6CkjTV5sUIzSQ9LLTb3/7xMmTAtaaWk9dWq
2jnO/V8gJOMTuWYG+h2LPU7u4BnMtdhcJSZOQvpr4z49WQOiMnEpkQsPAoxrlsOf
acpRGKp5FR2Xae1pdALJj3tVpIoiboRmgWl0TVEABBTuiF0NhSZOSgcQCD7QDeEO
ZZK++6str4+aaKyNqhS4GQdFMGRi7pkHuS3xdEjN7AmIIAhkZAYOf36k55JNbktU
nbG3TP+6/rlSYA2zGkH7K9HJ+EOlR2kSG1ljGUWTAjfWK76eSvrjz3Ku7TOqRoma
fiI9aoPCENOKZRdXNJPbTOAtqF7tcNRas43GDsaf5Eu3S4LNvHP63Q/jN7KsgJ8O
Xqo25uCI3Kir3QsUa/BfJ3OyInx9k2vtKcaI1x1ly5OhBYQU85YqfXL9Kn7lT+lz
wO/WYheyWrQLhxql5bVlgcqK4x+NwJn1eeQkkgDhGXX5B0RFrXjqLdkVylZJfoqy
VPfoSZPZMCbT5Tue8LPFLeagQ/R+j6cUvHWULtie+yHhoSVroowalXxxQpNywMyC
r3WrYtLWf5bD3FGNqKnNUeKKmGKOR5yxgPh/1/N8+gGAakAKDx1E0Jt3CuixQyOI
ZdBjRj9iD9fjp9VFAtsvYT+gIzW4VVKI92rLmFKUemgnk7RfCRofb28C7yny+y02
mUEa0R/a6pncWs+QK3Jh0hLbPqAnFB3r64ej+0og+sRd5JnMh99T5P6HRkXA8Djq
bbfUx+n0mDwXGiAJGWRVu7GzY0i7+Xu3VBBXNtLoFZSO3zU+/ejh+p8kQedTsUxt
FCm6hhqxIDlSpKPd6z5Sxi8cOLA9F65S+mpI82A/lqkbm8es8K8zDbLj10dRqiUj
l+UDiQwm+eKl8DncVCr4rWDQYSkk0OSiRHQ7+S0AFLYNbIQ1OXCbo04AfopomtlY
Zospglk6a5VCGHjzCF9wS3xT1Go85/FExWQ9Q9Ywjkt3zKbIV6F9X/IR00BTalLZ
dTwWft8Ra44j9pv0t+f4tJa00dMeZl470NcA5LkJLVPeS73QKgKn3CKkOwfnW5iB
x3HIz1AwEc2lfDADEAUSjyYqfBDvT34ylqSNwsGXYAP2kIIs34iwKkqMHDobVggo
XFQGXZNM+ofO7nOjNBsIg8NUMYUHmhNbTnLF9WU0wn/2mcev8U4eqQoosDbXDnGx
t1ugBePXTY9hhGFyUank3zH7U/QQcieVCCyl6pZGtdagnR6D1YSDO8gt6h9++YRX
QI+36wmy5UPcx+VsHCHwnHA54ir/OrCFnn79A3bZRtpwkfqPg8ow4zgaNodqVQ4J
j5fz1Ns59OweGQJwq0BN1kHD9d3+YiTEuK2hLgzGg8OAXad94RDYESg5+gDQbg+o
Jaa/kvdFJ4AYUGRgHkwCfjREtTBtfZsTHl4N+Bkf2pYM9uQL3HA8kBMwTnwXtE01
YSW4wCYInbWOrbsAg3zwLBqBlN9oIGRyWndZdVkxq8n+anv3EkVNjabea4Dh1JXr
Klduoy/y0XPdgm8VwwKcaMkBKtfxsU7WWLyDt9BIqN6i+xAGOaCZ1JkxKcQsea7E
/8sI0b30RGz70wV3ogwRA2mCXY7o7KNTphYe3tOE0rFZqAw2phr0xL2yjIOoLPsi
56SD4eETZOXc2PLovuijbNi9vxWqkDxXHyfyTZQrGap+n8dc+qj0psWrZG5rRyJV
/VHNDq83H62324bFDmBkxcN00DX1nGg4sLCXpCDTMDhRa03PNjuHCUdMboq1wnLJ
5AYxe6byvIt66nkhsoalDSi8svklOvI2X2rihNdWGj4yoQxxZCTRndgRffO4ITVB
WFlFiej3+72hXTWPB1NDes3NAij3ihLjpSN7hdvl8NqSidzvdc52L5IM8bFRA08y
W0danZgjMKJEJYyqwJh9aqxVLkXDaJ1+i/gD2mVYqM4E2tfYAyZwJbM1ycPl1+6o
fMMgpZH+v6iiyycFuGQ3bZ1UlGhzjvydCSXJUvhsrpTo42KpRpzuuyuG7BJ0QHGD
m7YKoRbvrolxPW/I3C4kWTuCadiGezWWSMnHLCPtClLN9ZvJqOp9M/NPNlgpSqsL
IantF7Hfmw8HMmvqhZ1gDSkqy36jyw2rkaUc8lStEwMjaw8JYOHOMBft7YcIVELs
RsmcTE4Y7ljvN80wdCEDvKmHTQ4CM+6sWyutK+j7m7ljhngf9PhH2Rn74bPHrzd3
kr6zX9DM1P2sv4ZUtdT0avs9o9aeq17omTXxd6HEh+uSy0qc+aRfeHMlJZ/2x/Ih
yY6r81ZN9K7sT2BVzawLrzy1Z+LAmhuMlv89PHTXIFC9NxM0MbYkd4eUUXOrFdn3
MtgtfahASd0Fia+GlSPQe0q5GqvOZSwpbDHXgmYmiM//Ol4NJex7zlJgqIV73QEO
cxugJYQsyi79dKyl44eL1lEE21ODc9MaYyV/vjMVIjXmpsHo+JvcL6J1Ni+GiEaR
ORBKz2RXH6muhfTbqSoCqeGU5UrgYX7G0ZzU9skrwdjimFEndHJdHNGFR9e8a4iQ
U/9+b17ux7PxipHcqD+BmEW6RaiNtacbjREc+V4QQSVJ69Hg1q2R/Op/Dvyb0qN5
s8oy+I/qRjwk4g3GIF530NqwSVlfRytyJ6O8zOEcSmiiwwqrlYJEEYorkge267He
P55/Rjt5PTsiEjFBR9Sk+D2LHojFa0OqwhCWnyf3eaUvTpeKFfXhfAg+5O36XJkT
VGtKWQjZK7czX6vLeSoDltSGvYyZEhwQPt/tB7ThJJwvMpmZFM8fnUKIqffwK60m
6GGaQDC+rSUKAKML5IkulhLA/iPevm3+RFyRMy6eyGBZmWftXWQs5Ayjlb/OnNMj
lbc78GJ1YukzbUphngpquq4ckBiXjgBrm7BFGO1sZ7PoebW+hQhWKerd31WLx4wy
PPlmpO3TT03rp+31vz9sddzNkrO1VyYXH2Ts3o6TeXAeJ2aeaqgXK0OHom3IIbVs
4zRmeNCXW4rSxQ9WgjjIOi+J8WbZheefJui6O8Y9oS/EasEojdDyGbwCVof6S8UG
J9+2Vo72qGMKH1quBI5mBDlrZsfjxkozDUlImqqv6BO65MYBC80aAFKBC59J0Zyn
+onlhk2vwtBnroU1eukkzgPnIcGoBvykYN2IE3hyA0kCUwAm9702ccbaV6Qje5HQ
ENB5k58f3MWMSUFw8tQtZAbo6J5IcG0ipMmE68KI61NAkx2sG+y6YkMBMw2QN/Ea
Oo8CsJUrqENL5nSk0aKLU0f/R0/Ct5yoIeNIrpQraw+kaDeqP1shQU1c60fEju4P
Wxa4/k2AAF4CZuX/oGwAm6hVdjtsuIRXS860O9Rze1rb9vo/gt5lXpSODmwGNp1j
iMXNPshn2iL/SCUT+rS88sr1zYobv8xXixBoV9q7Yr0m7DZ9m82fh1RE8UD/+ywH
ej4sonEplLVWyqHnRofE26Aqrkp5IWaXjBiLW4xudXW2FK3IVA+oqDt3Zm7lKqNq
73XfcTd/ZaefTt9MMZlx1KbbS75KKJtB3dJ3lRkb5JPBEC2/64gpiASYmGNtAoNk
t+mBOdFYgGyr0VTzMbpYuMpPv/HCQF4OG16RWJyEQzmJCXz5vUBYUFlvfc9xW9YY
RLtViG2fhwq+4STCIAS9UPI6hPy7dRB4S5bnuED+ZlY1oVummUDuqMoU9uSIS1UP
P/dvr2ILL9kMx1v2ukuJNEwdjf934jBbPkircAjPOVdwvsMCVj1yoxVNNE4+TN9T
cvYBGTsksMK+0faBpBbkW/YMgMjYPmVpK1HlwR+bnO2tgqdhhmCaPVGj2Q+OQqf2
gY9kB9hM8asOm37pV60FHAHqwkzjB2a0DSiF9v0r6Js6nsRDd72Zdb8qCbAl45p+
XDwQBMMOZMxG17JmTB8NA5jNj6L//LtWnuwNt4WpzZg1/FTAtN4ha2rTrU8BPPEE
vaDOjDG7YlyMbVcabtlJI9UdA3eYAbAzlO+mRs9CUbCDUOl7qhluoqcyc3IoVQsS
+fRmnZNOMCT2fEDOxV7N2OMLZktTvD8h0i4h0Vcq9piW1FyHt8e5kxJp8G8B4Mpd
p2UCiaCGRNVvJEJrvo2tM+w7wZz/ENk4eeZvvHi2swx+W0vLXdzVFqH13OQK0u4d
jKx42RQVNjqN3M0YjRXhxkNNegr0BAxaaeyr1pQ5PrNCH5JRhXlY60iJQ4Irk7ui
VeAH083c6KRi/L8GYFw4mu45oFLtLTT/0Uf1oTRmfFr9znwewOOc4MOiwvRzZdIl
9t+2f3exL/dOSMT9tR3LmxPR9tklK3/sgcsT8s4M0PeoM4HYnyeD85BRW7KRa7Kb
sNiiR1Mpd5C5cNBTrtT5Idk66liLwekERI7NmlIv/3e2LkWEM/gj5SbcsRFRZKNL
/7i0WNuPsKZZCGs7rJtd4CuEDAJTWjpi3RjxQ69lgWKO/dXNqeSaUx+a03pAiCIg
ZV8i3hYD344sIEX/GFRynuAc1hF2duv5kMmmngW5UKx+GTDtuaPPFWi6TmeC4jqA
iBVMs9FqJWBuxXCps5UaGmwGb9/hrOZm7/1D7XD+gaZ8vhL5FrY1HvYDIj8XhV2k
cZuf/4j7YgLyJHZGCX7aBceQrs6M5Kl3aQL8UTeb3nIU0ixd7/RNlJ1riFdpT3jH
pYIml9DX2NtLTe2VMddUYJ1+gS0Vq3hqVwHe/pHOWeI1opE5iOycLUt/ujGoOLoF
6lEvpQYIaFTyRxaDRjFoZoCAxhkAmcUgffvSJvQkwnfvjHfaXkBe1fpC+HcycKeq
vRvMd70bw9qXak+uULwZ0wgy69rssxs19bYFV6J65x62Xp5DjWFuf11gvZZMmfd7
EtPxY6dbRcUrkbn3Rq11elqwchk5rvvjxcemPnUr2fQEQ3zGeNQwKyWS+FDpT/1e
OSiQFFevW7DVx4RtdpX/0f75Gh2aiJIAmAv5q7uHccMy18hZho2GwHiBOc7Boi4b
t4P4xz1999vYYunkwFZhN4264W33Eqhl8KooG369ou5PrTyU9p68HL8e6uCwuL0A
5TSYdEp4OSflhusjupMIN6xE5GMiyINb8DFn/2GSYXieLMTSBVmD3ny1FJoHqxEC
JKudGWvwoa+d/a7GkkBbXVvpiJ5U65KDBqhcDyFriYgkJ4uKXWXAop3t0M8E7t6P
AuZrcIhi2YUE40w2O1ODj3INdVl/QlALIUQS9i1PO/m7pECWS3Ng3Z5qU0agZawj
2rAPaD+CTop3XIfeCYdRflgfXun9STDePb5Y0SIpO/2ebzjM1refipoqP5vhl8ym
QHdfDMC1vjF2FwaJKLv1b0b01Kg9t4SULc97mhT3oph7YakU+nurmjocDzZHdzVg
nxctZtecYCcshNxl7LVMTrUKj3m5YrJeFjk9VtGwynCIywAR1Daq1MU1E/PDmS5f
e2ir+k5f0MAVo4ArIe/GFgSx8iXKpcY92IWBn+oYI7Q9sX1XU1YbvneLx6nYpmKt
HSSYXWUiWJe2gAXkah+5jr9oJ7+InZrMDU12m7gG7Jtns5Hf+xDi3rlFElzteBC9
zy0TuxJaiIgVVO2qx0thqclSO7qLilOQ+MneRYCptqrALGlzaNIQh4Ob3MrYIM5y
Vr0aaNGP2CHKZ8oJ4nLdoRkCFa5LvpRO8tggO/ii6fJwgLKQ3tkhcKpcKfbFTCCy
GxrBuJaF4KV27xI080DNn87LgEjTicXb6jUKh6CliXQYml8PeHXYCJHBMRvpPxL1
cMt5BWw4cjRuJWAiXqJFTzR9hN/SOIlX4JFNNto6duBrSmn1YW7Eo+G4xnXHMY5K
f4mDFaMgpQQPSxf8BjijDSpzIJSlmRYxLRkExMKDt+fbPJck8TTksv0eiby2UEkG
02ztZH1AHoVFe1HBCY6U+4ascOZF836+aU8E4ne5p3gYKxy1MoRkYEB4fz+J7Qy8
ss5mF0PBI8D8dco4sH/ZPbyzF1ealOfCRg60ORGtbhwvqkOitUcqPTD6dauHkllp
Z8TGP5h0d4M0pfADiVewpEWJV2hd6quy5cXZhVomkfZ8ar9n6IneJxkt/2dcDkm8
RfjB4a9GoxFOVasmiq4/ttKAQu942gEfvnicrJ0BjFkUQJgOViTiZk6o+04Q51ro
SNppeZha7VJC6ugVS7SEYEW8yUvHjTd4Au6BLdoAV3JYtM2rXcpyZYzZhQ7aZyju
M2mE57Y5N+mEVNas9/ZZz2R9m5dE0B4+gzDliBicuO9jvBTXvJ1MdVglSHC6TSOj
ylwk1L8UxIUpIeYYaGcAkt3TwD8DHQ11Y0gZljtSHeHL39yhpXbn8ixldSDN9heJ
aEGDql9rnLU3pQieWrnTb+rQONyJJ8fErxwpu3HA6emPw9lQAf5FPl7Xw05G7d2t
pSzvgYFKJvGdmGjK4zliEBEwjq10rpU4IwW61MwM/a+lBsjGR4DTGFuRSIgAgbGG
3J3Dx/KAAdquWn+Ql17oWrsCBEmb6BUX1BQh5Nl3m0/YuBoGaSQuqRD9Z0GqQnDy
xoWzEtCq3f+SewyaF5u605mTIfIWQnySAQQOAOlqUODKTpQomVM3DLFROpwJmjUd
SikbLf1gFnjmh6zAZnKVK/sqwRoBE/4fug520TA/EQlhUcQ0CyH5un/UahO2UJZ1
V5nSoM2H0l3JNA+o7LlFQFuTEnhArtdjOaFJ2Gbns3oFYPPw+0coQsQ8TOtOy0Gp
nIffhHXAJS5xYPT3mv+PhZO/pdUAp3+MouSWF1n4xnBqDrbbPzcCb1ggLVClOZs9
VnhnWn7IXR67TosFBPMMwyhX9GGyHEzgH8rOy+n8EjijvXpWFvUyUSGZTJ3vTr4J
m1x0hG0s2gxtJSMQgq4TT7s6AvZA5iL5sxjzUkjz49VeJ0x1hk7pF3/WJpRCRnK3
zletjilXWANHEAZLKa/E7do9FH6SEBVH6WCHPdQLk1hQ0LEmTOXbNXYwBKLVOI++
wmit1EI+Ns78G2rDPAaRaj3/0do8YA/ZApMXQ4tqwXQVi8CHUzvopGRduB8CzkT0
Jjnyxnm8tMmfjkjePeXmrpNUU4wv+JqW4dJ9FXuTMFPtcI3dczInXo3vCjSraDsI
g9LyyVaGn7NqDJMi1exmkCTv70c3/31DsWUcFWjfyefrKt71bnHPoYlA164la0pS
+6S9ApMsVPapIl862qZf14TqtB3Wfg++IZnMiHd9pNs3foiICPh3BxQLnJEAmPA6
+IrfVz5Sf4ZmYmSHwRNgSGbvflGfwoJaZ4LFRxVZvfmZ3Di4dXyBEXStVi26tjgz
UOPzWHz/j6wcJ4ODeVEnrNrHkMu9RsC2Q/k2qf2XvorxyAMsRCJEwgMnMo9Q6MWH
Vx8dANqCDN7o3pn1sahFeTC5nWGYbKjHvk2mqK6tsRFlpXvMkM98NADblZezB7AC
nQOcTp6JyZarplNsFqooXK//QqZyYU/ZV+KEYYQ2+G+Dc0Nni6qJ2cnAC5rHO65R
T64L5w1GTgIQwebotoNAwCsC8PjcjB7wbbLvUppQuiVbg18/B4SJC9saWb645dzU
QKQexz2ibTK+rwVguB9uKMnOjQO3JSWLOUmfuzST5sUOit1BAxoIenqYlMQIzXN4
PDgIlh4qAKwK3yhCIjnCJcYkSShHOAckYLzv/7ZOsKb0M463hXhpW/TNhSUuRlpW
b4A96eXwCSzmBRiobkkVJrv+6TAnYIQMOS2SqvDK2XoNsjl/ejfZ/zGdJe/XoG/q
ezuRm5bjcQKg52iM6vShQVvqV6xRNzt93fS416m24Nrsxg4Z+rnZlG4o/k8dQB6y
PMmvjALmdR6EAtY3s0qmUd+Zv9EDmSoAa4Vxec0XwhYnN3+s+fAD4hbE1JU6La+b
7MLNpzW3CkWauy4sEAa7rsXcw54EcoGSeMnN6KxEuwhcLeEVqqde7mBgPQVbWUES
6fqaVBlFDltuP9AyI7vFidMCz+n/zis97RNvPK6umE0bGatqn9aVBiSNKjUzjo92
XE2g8HeG4Qb1qmWeXxKVHaTkCXHDfU6HHcdDfOs6etbSys418SiwxVn4Dg6EvWdZ
SLvGN160KQM8tv6pOPMAxVh+dEy9DUAlbej66Lau+FsYmE0BqGG6EgW1cAtcs35/
LcTk/IJZEdqRi4akkfO7pW8RSo9rYRmCOvES4Svq3Drb6wVPjaxzWpM8TTz94iv6
CAMUdCdIXIqPf0QyKNF+jTGFOEjD6lqZfIUUTqbiPQUFYsXAZP7p/Uk6DMbPa6pF
PUv3PvA+cq2+l2AORsNOUQLDx+JsYiMt4K98XaPNFZfdwoQm9Hqo0oukOqeoiC79
rmElPmfqiPQE5Qtgaxvxb9lEAvHE6kXw/TC7H2/bO6Yi22gBM1cal9g5Y1d7qlud
Kt1CMjd7f2eXnniQHJXBnNtdZwHr0NolV1zRQkgDBNWfXL26C3Ez7zaK/IcxhRTv
bUR5X1bCJxe1/wtYO7NWplnPwjl7zrt4H5B1mY6ZdR5lcLD+1vxs/aPCiofd8OF8
ZIpcIW4f1Ad4kbIczSNTHy5SpBiYslQoMgKKDSjUHLfayix1Lr6TLl9deYHqN//n
VnWj9TfOqTPqMne6piaH29VEExl0SY64ZkfPGYFwBkCV68XM8EKkgPmvxkEp20Zv
7sHHHfZh6AzFmz5vvUBt6nQevLLxP0KyQ11ERSZ5JC8mwaearFZ61TtsMfmcFADu
cA1JdO011dDB1967a51xzcFnahKTVuZkyw0gLym/ykvPbzKHL4ejEFgySLSJCn9d
cGygpKv7i+d3/zphq7RlvUQNQeZ+iAgLUTmVXACg6iuwOV6B4mLaKmW5Cwo6LcLx
1qetSYAOtJPk707zAAleG/hWmB+3vYh10u8RNpZ+pmxwh+UhFAqTchC7JDH/jyWw
CsixaqNnlq/aHXudAtOz/OzxYYjcI/fdSkTh3YG4/WBRuwE1MPrXftXLgfj/2Nsu
UsVFSCfgA3IIDiHDD3UsaGCr715Reiwrgftq8B8bAj+apGSVssA4TihFrPJoe0Tx
LPbvwxOxRbu5npIdQ61q16qmnth0ofDYqLNJV8o1GBP/9GGA0tWBJR35BXZ7RaDP
lhaSCy3gb/G2qSPl1eTekKWdO49KEFgo/DW5xTE4mKtgn4wt7pEN0s7S8FU1nmnt
zoLuEs1EayO4vs6dGADPDnxtmSgZlfqzgIk3ZmqJJQkTlm5dwjSLhnXnLuMq0Hc3
PJrYRwn3IGoi6qfqjz+TWalcTlSVT6nDViqZdrqO2LRidwPIhTw3q3cJDlJUoi/N
TcHBzNrasa3z6P1iIMc2JywH3uyVJtkFn8zUbLH7wb+YoeYv4qzlpLacaE76uxNA
dRuw6Cc7Azj1GUqdk0htFTE0CO9MzkEHSwZANmVFohp8uvLrc5PbMXNGqDCd0AsB
00qROusRcms7Hp6nN09VvtiWSkiye7qM2tg5SOb1eJHhmRmnegPezRpGUSrHQaPe
Jz7mU0fBH2Rn/imzb41TRkGHEXbMhvzDy/Xe0XNExDaMucpua4NUz6zLh3c+iwtI
gxGgfijdFZmnNIwJT1K5Ts1ikaG9SnYjG9TjNaAfHn9o2NBdaNajaTedIEIFVD1a
qgGLvYO4gpHcjqWpE0KHXklcvATOfzSBhVTerV0pua00ekb05tle7BUhVRts0gQO
j5aq/8GTNVYswfN2fir3psAf0gxAmtkC4GX8KF3Eljv5EwQWCDUs6FsCkP04rOqD
G30G+Zu3bM5pkAsQ4hQVExaB8sZpbAn6ZqlqqmeLBFH8EgYK3FEsbpRDEfCCreSq
NBznNu8xgLHuSE0CcnJdwWnC2q0uoZZJKy5QcbHe5Am/ZhzL9I2kGxLJhEHm/54k
IG+hJpnIewuVfkfxJ9eZhJFEFU8woQeD7pBLZpM9EjYeJO9xvr7CUe2cQ7kLOQC8
ETS/mLmJyQottfTl0yojzhFzFcjQNxsZC2h4NI/coWoUxon60bnXXnYeJMMwgB45
Ygy4pMIR5zfxYmLNVmaghf8lMMBC3HQVwdQ5jiapC5C1nIBG2oD1ZzuWPbLQpRMi
pu9WJ+/WSaD2RVymE5hchg5wykqxxrZaiVbmgeZ4omW6mMEq7x61sjZmmVLOrWzs
VihpUuPNI9SZjcLAy3W2bXRDVQqFJynRmhUoP1lI/nRhF9Yw69vzN7DhfpZG2AV2
0ngE0EeA9KH3+5xNVjeiiWyiTIYuC31YQu5y9fyKyy8zyPFUJucvoNVTwn3A9RVS
k1y8hg4DW4tKej/GEAA8Ff+F0RNt1W6Fs1VdzMv+VcwW/xGggtN5E5Xs6BZ47QsR
IjvqrK/Gcw4qrAc4jssp2vkpQLOEzGdIaed/X0T9PDwnUpBi4WsZQRBhdqZvf/NL
/kgHVIw1ju1GtZP5MeTNnFYhCX9s1ePXZ00BRM82K+L4V7CXn9QgbZjY6fTl2480
qirx8yTg/bWu68ASzCqkHXPbpotBsFmWwHObhH7a8lWvK9gjfrCgL8HVjxOfoFyn
sRZeeu6Kisol6YRlg0tWtdz43mNsKXsKkDsb80Wg2jhOwNqOBGtVJlWD4FPSnFmE
3irG5LTmKpqATwQKstBCucLG5qnl5Z5JuYQAuDEBR5CkL1VgsQKwCvOZ33KkjPZu
ybL2djeVsgpyjFizuln+RQ==
`protect END_PROTECTED
