`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJPs6ATLi0n2nIS1QGmbM62wTVzyTCyRzkPe5f8jUBOJPS7xEVm65ZFRJeNQFiRd
ZcBeLLVtKpsgqoKxwZnQ9xgKIsDtVdCnS2dP8sA8CJM6AnGIl+vp5iLP8RBIPZqD
dry+2QGZF80EUziE8+8KOFS/rXUIXDkC53Lz0K1h7BX1eXrhRRwPFbpNJkXulADm
5v41Cr1DJmiaElB//4+cvCCIhuqKUvJx0QvGxtKNRWiOpGX/9fCqKw5RPXML2aTp
GP+5pCDIisWz/Xk7vQl2mpLYKxkl8OziX/JSnT0SqrXSOXrul+UyssxBxNlZF63g
cqGxThHcnyzEO8BsVMopSfHf3X2KU0PYvpTaY1muPMwPOXz47or5lGbXPyqkNuuI
cj3cxZXL/ZNiko0PTKMX+AqJCwRlaSC4OnOSQF3ntva+9b4Ua/cK3W2n9d+VAECa
/kXMVuhHtXTCkectDYOJBDS4Yn+7ULf4t27Jx7f864A2+f+yDE/TF0x9H7xgf3KW
XerE/n7h8xP69OT25FB/h8pbXvlQBGXdf50L+nyFbAvcMDoP3APBhbWXmdIRFDHn
E8Yk3DFiiFZjs4Ey5hoh/8urMkIgd/vJCocOIWxtxlhTNEwNcXrqkIUBrXV5/3yP
tmuGDBUSqhkBn/CX6pcie7j70GPS5mj6e4L1j2Kd9Eso7c8viyJ+DJXiSnEjrQAl
A4tAxWZ5LMLyOmwq81iK3Bo/uV5O94xcfa4zuw9c1EPeAl0nfxMq2xMTHMsGIN4c
Ufqko+Y9VH1eG+N8mSNBO8y6TlUNjn3FfGjhvgs8w523qbup/R8t+sKqhO7SbevE
FvheeislcUx4Wy/gmTCGyA==
`protect END_PROTECTED
