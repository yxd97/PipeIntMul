`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HEWH1UlVs22ex7CBnKUEd+fCHTvJTBMlKckj1+Lr9wqWf+iGwu2d9fZbNJQ5Xz4D
G6zWidG9/eW5PldkYmddakpWHLmAw6Oof51IwxQtTiP2gKrGiU6dtKnPRGuU52Pg
eoYgn2Mw4z+uidpxz8SvF/LdBTZm3WP6kChdjd9Huc9rdJY0e+UnNlEGF0ZWD25d
RDv9mOCpjMb2Qilq+lTSvTW822GXGHQCgIBR6XoNbZ1YkwLhUkgaIG48WgHTwCao
QpK4gFlQxkCSvHd3gth/ebdwR6UMCDXCZnZZHWjJK6b644pjASsnWhVgWRNz6wHu
k3KIihPak+1DJZ5IErXJ8KoDl1Q31pPFk1+GtKszTo8Tml6xpttx2SEny0Ek0hcY
/VWKFKDegC0ZXkU+8SMsrA==
`protect END_PROTECTED
