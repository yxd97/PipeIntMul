`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZBXUQOUPEbNqX6uq4pgAfWtV4EuajnpzQlZ21Ro67VSrAy4Qgc0SXdG1lDgoJwp
s2Pf/hAjdHR+0d78XJEPLMox92VqgL2NA8wjIebg9VVuBTpDpvCR9RRLCLMOjaSO
oHDuyrbtadOrZISp4rvhtpCXcc9OmEW7dp+2/4D3l1L6GO/2F7wsHiXMVu0QPP4n
Md2wy3rwPaI2uft0WXOUZ+Nbw8FxcSivSNAFsWIalFldzcdMwcmy7AY6iMlGs5YS
W6bhggJVFg8Osbj7MT61s9LRF8p6I2R/bfkl/3muTs7edFINIgntA/UuM3w8mFxH
mdCYOK1/MVNytzSHCibJ1+9uhjIHI2/0z9hbsrA3SnzSd41prz5v4Z5878zR5idi
VCzxKmKT/MfZsgwUkjlDhEvSDhTtwvfLh70tNq1JfY2jtsfUnD2h+AKdlp17wUUB
jsBW+5N3qUt+NV9zVPUOszhnfgPIiLk/mlOMCn3cOxISkzk0btgZ22mkIjz5rjmG
jhfvDveGzcoo93+rHTUOL1vTqPmIE7wM2D9tFTjpN/6qPaa09mGU0BhBYY/P5QXA
mGR/PtY9LUNInPk9pMJLn19COI65/I75MBXbOQ9C+qLoSVkC4u8CtBEl5UmR3aht
Bo3MdBwSuk2cQdZlMLYLA7OZYx9D9LQfpmGinwwM1gEnPMz2rj6A+xeqrBq7FM0n
mppHdkA2q2q8lH/X7OXmIh19L3vsOuhYbt+AlFkb98tZAy3Vp98SEjTedbFp52Mq
TCnYbn9YJ1EnO8k5kqnwZy29/Krgzc9iQJVw95QI2ArgdPuehDJU08R0+gA9vTZ5
Ph0jA45GBnxk0l5GmZpJSEQ91PucKPyM5LntyP3XqsS0vJTrWlcvRR/f3raYo97Y
j1PTSN2G4Ms0zYqcA/4occowbpELr4cA7DTccUOvE5fBd5vOk6Zdf8SiC9cclYkH
TAGpGPUYW2yiePthVvxzZ9x3+xRHkGrFRajHusLKKmbA2SObAZxSuGf7erUMZH+i
iDpaGEoWNiLJhYF2zCAe8Mdh5XntzzbK4q6SqijvNUmPDGo5tr90cl2rUQRaHM0h
oydJ8T7RBio03pRmW/KtW99LIFkltrb1Ng69v03Me0CjxiVcA8+XBko4O4kr1Qji
oIVPuusiqnKRSIbTWgPY4HQzm1yg3MUdfvV3MdiaVLs28GVaJd3nnYFRwSegsfQ8
rbd1S+frg5DWW58V4eOYT1NhGWukGwiDexWlRUOyeiat9ctEE/vKvlcr4Y8oXs0d
`protect END_PROTECTED
