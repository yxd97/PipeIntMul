`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6BSTbSs6T06A97YOMEfRVyJ2kkLkFGWxcSndSSvtzcJMs7Ra0CTCcGE/nE8v6Ov
AeZtL4kuq+DpERDvZqvilzN6e6cUzRCGUmg9wgfKhwAB4oAYbmEkqBjQCb6cffMr
hV/hz5xUdc3kRoSbvXeQjRDrtGEque9h+mSdZ6gz046rpY3IBQK23J5zqksFiQrh
D+sGH0vV9JsX+OMx6fHLIfBrFLMf33X+KVV0/bMbJQBFzRdZZ4/glOVWwMkNM/vf
k1Ifv25CYk+aojMvpL8BYJ4nArN/PjGESSCCluR7aHsTbeh9gOCxoTFRhflP1PIj
tF6pwukjPCdeJug0kuftQNZ56YYsykLJiuPiBDYKrYL8RJnGI7dS6tfZb7cShP56
X+pHQ+v63fRRI7z4uRblaG0omDfaiwZ9l8HNaAA2e6qnJOb3rYbEf298/PMBr3jq
D0h9t0BZsXdY/eu9xA65h2HXUwo1WJQ7tq6TI3PNbs8dY1EFXtO1sI4FJjGRDN+c
CIgyQP7zvwp4LWIl7+7JcgHM2PyJnGNhNQQq24AFmT9B3wbpJiMpB1KuxSFJJzKe
M2nTTx4NBwE53Yo7VHYh334qBujSzK87IUi69hdATSWEqac7h/rK+xlTIPPTSN0w
AxqO/XYot9HnlCqyAtUzOxTrOVOkQe1aBYmQ/kjGqV2rdmXqHW5wGKdU41B2X9xZ
perGGsnn3kbeS97ZSJN4MBmd7K6YItYBz1K+xw08ED44aTUnN4mTI/t+K52TQxsv
c6hriy3f8O8VbrSyyC9Hmn/flE0Oa7SEic8Gp0CHqBYUKNvUQkYwaOu8ttTtTtvz
H8L48aWnXeNU/S+3JEqhGCZNDCJhubhK5N0sD2nuoxNgyBfT7imNNupu978TCGNm
QMzPUyBdJVAwI3mr1wyDrv2ZyO5oy3sXbY0VGuoIph/YCzXiaCCqVghuRTw5di/s
BQ5+irtZF/uz7iZjIsomXt/BGcLxh1iFDib25pAZGr9sTMVfq1l2NAgoyDuafOyn
cfgj32L6XaAjjnc9NYX5lwWMCnlEhQcsPfckdlsExY9wfPT88LJdkazVGQesq8hY
4+1gq9PpfRPU+wyuDy/dVptFpCrYIk2TSH/+UoR2DWshhV5ynfe9wNDd4F5LM52n
CHSba51QZiWiqIrWzpXXHWI2HF2f/yuWTO6W6OFCXm+rBQpMUUHimAna7OTwZtng
U5jebntRz8vf2b7J0Py1hVW28gPhUOiDNkVO+rppsQbOg3TFtO02LMK/GuEI3vj+
6otOAOAmfAmGGqKB7S0GmjkDneTuO7LkhDyzvH5sE41Sn8Pnn4WSI742Tjti7X70
Jf3uCZ6VMewFGTxhratoDObqAusarduWedCMw58QlQUFVF7usJdk7H971mRn5j8W
E9+d0bXjnn7ToGTMLlDz5cxoNjQzVEApvTKB+rMH00xQshZxkDdFAMpBAYhMPs9A
aSy3GvmZ/YOLNrbWHACioQdSzIYDjqMweV6z/zmE8MWFoZbyz3Qg2UUjW+5yJOCH
lo4Eh6lpw9nPT/eFJI00OZpn7LIOWDpM10Sq5u9rX0iWQx/QnqWzv75oRjkzJb56
yLi1RrsrCFtHUyngnd3drZwiZO24dNsmAqxLPDyu5ycDxQQn83+5Fn/qYk1BFQ1L
vlVog4ZW7dZarwVgKFlj5bLDYKgARqnJhwbtMKRLi11ObClqzbgu16DUjABuglEP
P6GKu/IeWg6ChxZYnyEnETCt4ZBEYHiIenNKHg3GWJiF1wAWrl2eJ6e/F5dQI04J
j0nzSJ8fq+uVmwwcpxLH4EYgjH6Xp/uFUMcFrSWaGW5RHa4qfPbjqtbsjSf7M4Nq
gokxLvyWX1/JD+u0z9vHLVxveQpyL78gEtAzVfUpFcUIzu6eNGZCmLlCSWE/8vJt
cAkZw+KdEB+R4xZEuvoErb0NwJTrUm9+VuzSCpzf4dtswgR/402pD6CByqWF/UTv
im0GqhI9SuNS/PDwNG1W9aRh5U1K+iFnN1VxC38myPqADMiuLrTz1o5h4MOCowA4
69/vD8XvzQnIhQuxqoeQqcZ8y12bWpOzK/x8Eh7TaorgqfcBH7tQQ/EjhI6nhtrU
Li1qfP7zRFAODwtaY1MCKNQwj1GKtKpmsglWugyfMBYmmoCAwba+92R+uqmx7kvL
PpZIZZyMoIiNYenYldLC/FYsRJSFNjm0j1zcwKY2ddG1g1/+4+nrAR8WXiO0XmTj
/Amy+TJQ3XvFELTHBnLDu9pWKGBQa7unKyFZbxXir2wi0kMk/LEbGDjgouSUaqhK
f/QKcg3QDGnRc8NoNApZX9MHE1R+itfKd6LnKPm5+PNccsAmjQGpExalM6lazjYa
5UNGyxILWu9xksnCpDy5RwH5v9JTkXA3GQfs2X7u+n24MPQnwxGUp6j7/11Vh6Wi
IMbNtbHKDcniyzmA1XLVrSQlC0HrpTMq6rf9Y4VAy81jyKk24oKixisBc8LYF2ot
vRR2jsmtwnHVN1XqJvfEk2eKGFEn4vvJaEj3OGEHna51tf3WNtuZFD6W4T0PBrJy
3w3Ef7+r3/0XC0SEhY8YSkcpUCpt4dYNY8EKoKjkuahcz/0v6I2i3/OCE+6EM2DY
9akSDM1T+40PKv9+ahDchg4D+iayeh8cAuIHU6h841I06bd73caAkaAVxqaALsoD
yK8xFcPxyMyzuInPDy+3YSL21rrXgHkzuLvljYGK30y9VxGsRyppEN5K2p2E4wcZ
mgbHRv8o6Ri04fAgjG0E0OvgmfzHufnwNKKmuByEil6/+W+AWnIlva7d1PPa1F+9
HBwAOXtlohmpXYsmx8WQg8+nSUO7CPeoJGH4bwKhDHttPhhem1202y/cSs3mnEMW
Cub1RS/VXdra71sYZgSj777DjakmJ7B92EvLH5ws8R2nisPptGTdv0EOhBGapZbP
zcYP41SKvH26R61fhrznCFXfpxYsXnDZpy7Gxpx2J91mqMHCOOru6gpWAsqeVqw5
agJqJQPGn/pZ5INBcHvlNydsOKuR7dtiIAM8qH1rG9zdxvlwbASM8aWjVVHRouzY
NQxxLYYT7D8/2O9/25bKvfFKOP4d+a5/FOQ6bSiC0nuw1sQll8c8w+1X4d/I2xAm
nBayxCdFjUCuuAl1T6HehR2QMOa2eqsySULHH7yuX1jgljv1uricYtlfur2U2/+R
9D6CfGVbKiDqsHi6kWnX9IL2uU8+YHRwMILxAyi7fSND6eRKfzcQmy2TNnZyEmD2
1Mp5cPx9c7+rFC52nN2cVWLcQuiK7Ohsiqcp69E1oBmyO7yDchG3/wEMM1tK3Iug
rqH6uDKmd7iVVvCNxN8wmo42zUA5LpHa5Jb/CCCFfnkeyPkllfl5j4EvTvUar+pb
+ZF5xNjtm9/WhkHyIgW+F4D89gOdz2DmYdALuuZAf2Zzt5yIagu0LJHpHle0e6C9
7/90mvW/seovbi82HYUPBODtOYQX51++Lh5ci6xu0DyAVXdiSWRUIvwaXXb3ZW15
Sqbv2WslRj3p/rAGaubK/pkIRd55DD6Ltvyz+kjsLrxCZhLS+bpgllIAyZEuCARO
EIxaYfDV6k9n5+BOL3G70RPc7R0FKmwOzVNtQOD9UstL6vsebeWlh7b6Fl1ZGGCK
0hOnqM3OsOfKxgEIYawRUhKgNiupKhBr4CAWcxSxpk9IezttNU2TrLC72j2Iezlq
jBMHFpHwt16u3mQkLigVbWiWsy2UvDGlualCaRTFBwiPtv2N1ST8w1VkHUFdw+FL
p1MGWZEnUGkqd4tPAY+OXAbGsGKDQEvAcqrmKQF7ZYf9WynHVLEDJHaj2Lf9QeCG
NKSxTUovsu8jzc1DM2CnHgCU+ERJbkFAaHqM3ECc96WAVQAtxgC+lwM8uc+O1Ntd
L7ewK8mCTulD7LmKbrbkpVdv5Ozxy+vPGB3TunmPHujXY4JzD85EoUGTlN93jDl5
7sHUN1VxJbiLBI83tiUmVQjRvXtdA5avfClzwqrogSWQ/xgRFv7e8Fotxlz+Wncd
a860/QjgEjDoyXsxHhB4IEWwpWf4WceeM4+w8ac2/kI6sNsM6wrZQb9kbc0kGEMO
nkmNKilTzvR7WYMKrXCQe0UX96AGLd2DxeQLUSTvtP7k9wWLWQgpLJPiP1EzL639
`protect END_PROTECTED
