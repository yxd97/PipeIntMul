`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OKwEtBqQYGKB+A6CBzeALzW+IPVjkH5F9paRyXYI4HrPsWg5fIKCiCzF0aW/rSgG
APfNWbmhZKYdDX6VLnsNHEAyZzCnRgdAQvCwBwV5pgB8xB4zJz3wFdqsIm9DgTC/
STE6Y/7RZczfKojnx9Zm4phcIiN+VD529SJTa+snQ0mEXme801okwRe6CCaqw1Ia
GUSkX6QwHBJkQ/WvjIU8CKMyq5CSt0Kq9TL9oOCe0Yvqcm5vT+rEIWrwyX+VP+Zj
h2DeponmhCRBWq8DVTsuPv3PgmLapb2JXBKlXAstILb85QlSpYRLPk/IucYwEcan
+i1F7q4yPRJSKYqu/G09x9ObaMDeVzeafXPt74Ok5GqEKITn04BZ9J2bKscDAaD/
LtUMBEexotki+EEzqaZAUmmksvM0wuN/P9lKoZqPsFmq2bFFFPTuoWEqoLnF/oSJ
fv39D7ki3zVdaXuArt/AMnDRsrLlj1brT50G6CcauAYDmf0Lfp81fVXRbGUob0nT
aQ6vbxEg5enHtLtDd9y+K7IY+U4gRKeAKEmTdmY/g7L8GNKMH5ixjoJSCX7K6AGF
DpUnjY3gk0OID5LAQxX+pftQ55USau31CmJVwqtnjABwXOjmSxhk4HsnL8BgJrsI
FMBUWqEGkfm12MKybcvlV1MPhd76xNlGPSqoLKd31ByQcFGKlp9yACKhrCxNmgLn
pYb5bw6FNx5eseJ0N4UuaMqa2a7/jMGqUbR21DkS0UrV4BRQDBj9r59aLEwP/CcA
YXLli+j6qrwW4dGZXHmm4BhHQFpvFYAyKdqunOLxavXvSY89mRZbSLPI6HZrGuP0
vOTNRwepYMzMjVz8q9g8/cXTiRo45AbP5Q6elTrgBw6PZhhLmPG0Dxj/25Gc1Mcy
HUp2yofD/eiVkojg9QGSm9IpVT+3eZChpy4jZCcJOqbNiRl1qgaZQtd9xHLbANVr
JFFQl79Qf3v4Eg3f53T2DPMFJfxcHqXOFLT3SRu9uz7LLw6w69WWtbQVxESAAHKO
/3afdOX3O8czWGH39tGBwFyL5/iJyD7aLoUjvu3ja7ba27pGJrukXn/WI7cXwMiP
f0UDp265fhvtM+hePbS0QGWZ1voVOo98SeKGoG7QvSp76Wup70IbxfoQKynD+NTJ
jbfc7/CPA3F1s3H01ozxw7g1G8ixbGrCdpnIJ82Rx5RVDynl9Mg0wYIC1BHmA6Ro
E5+QcrNoWuNSW5Pkt77ifcHLGphsmG4+S2zvKXDk2a4zHsPwuW+0djMUKJqX0qfE
AFZdOxSx3JEZkvcPlYwZBpy/ycBK9KHkzctpnmopcpPxDt0DXgDxMkL/jFOhc3Ps
AtOF9A/MCJjMaLIw01quY6zH6Fu4buJiWiDW1jyuRuclMGfbeEUegHd0RaBVejvL
`protect END_PROTECTED
