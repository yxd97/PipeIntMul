`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5FNEPM1meDklw9vZIQYccQ/mGzdPxitZMgS97PUYDTvOlFWAZCqXEo4FlbGiZrxS
3giuFzwral+K7rLQei6Hx58iQb4I4VbOTdAfhi8WXx1Qdg5mHCK5EztkQ6VDfsjK
3eOUd5r5MJ2lyFM9mCPTzLbFyNocrXmWZPdsnLrbfIg/HRafdmY4vvaiFdOYOAEw
z5e5OnpOralUlxxpxZ9Bvnut67gNdUDDO29PNRJKt9FSxu0Q88VwsUQ9BTPuYNyH
xbj7AlijkWyhZyLW1KsT70JOIKO+2bEbqRdztkx+IRoHDsz/IJ4L00Qtk2epVxq7
ZkrVCp/9ST1QCsOxkozF5VLkz8+RxUa4vVeSi1ry3gqVth10R/iJw4nHqPB44s3w
+G6VT9t5qSCn6xFkabiXkaIm8bzQ7Mndf9Chtwrm7NPYc00PGP0fIuO7MNzx3+SA
+5rLiTfXElfbzYbrv9Yj1RV/duDjavZzFl344T8m/XanvlHGKUXyZnwm+JQKiow/
QAP5LSJ5MxG/b/4E2UZQsLFsaM7aOv4D1HZyWcpb4dBn6nV4VqPKsziU4LkJQXHh
P4iC/wB1BF24RFRbVAojmkpIyhae1B+xxhBDO7kOBVzOMCvBvu+YMomcc1ZiensZ
uHZ8bDQUDWrPDiGc9DYU3t2iE0GI0Qw+lUNriUpw3wk=
`protect END_PROTECTED
