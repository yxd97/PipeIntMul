`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6dsciyLLqwz4ZEdW6uZnBUpGPC6mRfNZ3Tg4sTE7Aa+PaPkxV3ZhDSK1Yv6oQ24
SyJZuUk/DAaok7iVP0F6ekymOD910kNrdd6RNEJeug5vBatmF9u5pchpYiMVbFgS
tW5TssVY5l6I0ou0U0OSZ5WOUsSZT3R5UE2l3gBkh/2pXxHdxJ3iYZRH98H628d1
8uv1YUwh5t2YuDYByENVUinLizix0APGYULBt0uNxkTjz9U85DMVryRpulETQpXz
r8jBJddGpMEmTDM7P119Y3XN9im9iSjwRExcetskJQy/0dbop9emWziZDo8Gv0mH
qBytc0n1+J9YoK9ixqfd3NmcbollV18XB53887mSqA0cssBniSTSQCWj9fsv6zek
Mk+CbZ+ic+XgG/82XRMO670hz8NolpP0lzGaWt3TVUg2nJDJvpUT5NuY4tgvBcMQ
j19k8X/2cX0JtO2E8Jec1m85gBA7Cchz6IZH+Z3xviiZyTRIpxZlh5tZkoyunTVO
/U1/RW5Tgs6WjBxj40CUCxmxGhziHN2e0t6v/6XVRhN9eOdCe5y67aou0fsYRH65
Jsz0alUC/zG+K8ivo4pRahSMy+SlSASNGguum588Zvzw5OUUbXvFVXuFmB3m+BYA
XnEFhorIc0zYKyo3WQQef+YrymT5TKAlb2LmndDr+9vj+wTDTy1JONeym3nBWcTm
Lmofl+WDzlmvipUmxD/OBQ==
`protect END_PROTECTED
