`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uEzpetQ9IMCJL/af1N/icdhSJKmikueAxuIzzYOgfJ4JAzfNTUmPQ3BHVXWqzv77
DcHUeWRiCzwUPuanyhDdBx13Mswgn0ElwYTRf+muo24rbKKj+HARVC3dzUxKfp3d
qyVWvvlItE5kHOXqgtRX6LXljVPQ+8BI+MAsZoAf5BwynY1LT2D2XlqsE9COI5rm
FGXZ7sGYt7x1bSbjkXoQk1GReqI7Tl0XKpu0twAXC6f9H6JG/LsnYlKD21uYmMd4
wKS7nR8cXYZ3eDAOmahtx5nxITjgDVHDMYENmaFDFSXBsQTuA48NlqDDSGgYE1cT
gV/Vd31loAXLG7VJwzW8ieLnh3sWfsb8RMy/QjLo5jwYG/2aMJEzC8hGB6Ld0I7z
rM7IXuI1PHRIOo2tkEbURG4wCeMEfPUIHTRHdjn+daTxcSap48rzYPGVSV2CJp+w
FEF1/adqmSRELdOce14chK5cLGNw1S2rFWtN8JJCrZZQxuRVDHv+LYUPAE6AlQr1
CM2wusjylsojwue6B0L4OB1QOKreYLcKPBPTu5QtFz4c4mdoMlZIiqq/cj2X4hyv
/M+3Q+dEOJet8OG2GNHxZ1eCBiSlFl9elNYU8vD4qhE4soRB96ozzwxXPf1/wdXz
MrWMrgt78jDnzqw/klvH0JhU9CkmvhzGSaGs6ftTuV8Xb4Ur30lhh8TaJbKDhguX
Vmb8Zf7bmrE2A/aj9RHq2wUvYX7r6D8IRtVqwQyBT3NtggjQ8WtsD3ApGO1qCG0c
mQpSNplAA46FChvPitqz9R7GI0v/R1Fn3vdYhHsLKfCCZwP8p2IWfrB178s1zLnF
TndZHFJWpBGUbjAIvd68RmmslanlkMw44hEYqbUx8LZRg/0Y9L6sG3pi5Bt9z8Vk
R3fDUXkYBKo0oXOgadFMZ5w4J6eF1U6lim1VSTzm98PhuLq9V4aTs94GPKk+hWmR
`protect END_PROTECTED
