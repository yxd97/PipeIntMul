`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7cAMDXLHyT7z22P708GrblphUPYUSXBoEmzIuiGQzUCXQaWAozCPPJV32jfnS7iX
1ksZZ0nfbG1MNngNXIaI4Ab3V4lOHUocjnAteGinx7xnGq2MNh6gZm5MNXLB5Fo7
w68ll23SJ41Jp9pLjZThmvnaaBypiwVEXTrtCR36YgjNbPOI8LSJtoKBYGPl3FHj
dWYO2YWZNz6XskcWGSM9NeS4C4vvERBTlncIWFvBoq6rDNgwuAuD4jJU2Azc3rIM
q3jsX5+v2RG4xO+Mv1r6GIhaoNVHzH8vkS6uflvk24iUPrrSRdeeSep1zwgnWpUj
iiUXbQB2WpH70pKIDMXDs2WoyJsrC8ksWTrgS2Lmrq2Jin2+9uDuBH10z9e5E6W4
MuIZFEXZdNkb0m0s37WAeO8E7NiojxfTvhjb9YFGbvM=
`protect END_PROTECTED
