`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IO//7Q/qJ/D1sFJGpKPgwoTs4GC5sDl6zGcH9MAwnHFSvQteWZsqi93ldQzml/iG
RA9RYtTOQbdsZ15QnnVXYHunT1N3QsbjZVLFqGwoz0OWmI+J7hLTcdWTih4VFw1Q
ujaTDvUTxFAdzSpcrMDCGM5rRslZBszt+dLOL2KNI8OVhfi7N5SaxFl2dg2Us70Q
3EwQdA/PP8chOiaIojd5DNiRqJPif+d45MVHhZvbq57FyjEIyHbpJ89tF0ujdrHo
O8BdSm9G8LU+bSwu3yFskZGTpQ/UwzoAOgXI6P/fhfLukh7qFTEBMzioel8q3yPa
VxT7U0SfrGD+jUSSji/wi4S1/iqN51cQTht8TrpGrjr8Tf+Xw6IZp0lOHCXmQMtp
kdLaTZCIwegGYH8ibaXaDpKi3nH1z5RH/xTp/C9ebMpx9tSEetP6bqJ6ksExtFfg
yyVddu77XlNP0rTokL6CntT1yOAzKnU0Ik4jvfTzo4rVv1dovM0pPbJyPLjIN+x7
9hirGi26lRWRm03veBjREvFjycKfnJBWFVaZ4ghgpdOmNo9eZ0wt2t+hyq2CAaWt
8ABLdHqEwEcEawfQI9azcv4PaBQX8WEl0OxqcJjT677yZfrqBZ8nsDDb5SO1rFhT
qK0QLs9CgEaoAZjfWoXV7g==
`protect END_PROTECTED
