`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MDNLo2IiSvsh8ulH3WXmDBBIgZGVIJ/d4ic4AIJ+Q6bKyE+F1sBjirTjobs1vhpb
f4SkCMLcHyJgrtwEvhaC+W82ma7SsQrg+R9yZFQVEqnqI76ksmNHEjaz0TUhz+ks
Q1xYnRP/7VMF9/2oKGYcQ1Kk/KA95rurAvoqFRcHLmqBX7Jd1f1xD6aW+Su9C1Dn
IjBXDfVfvt1T6IZGVRYA8+jwFyEWmFLx0s9C9D5WPNkNwqyX9rIVZg5mcSxzkLv5
aFb7sJn3IwKXxgFkeGBtZPxgnYFhF2xCeAZlhE4nZMv4gDCmxBVEsE57P+Tv4a1l
tN33X/M7pWyq7vUeoGGEJ5yCql6x4Ig22XBozMjQHtnZmTRbRmeHkuA4blW4PFkq
ue38D1yt96ZqXnbhd3Aaz5c9FPIAk7E0Ia03AbrMUF6V//CTJuEwFJ4NceHK8Tm0
1T+evr6n9Pd2G5cuoNRY8HuwAyuIHQxj42rSutfweSbBC4xJMtdoYw4+EFUqzesA
`protect END_PROTECTED
