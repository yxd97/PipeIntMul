`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1i+vD0f0E4Qxhq0n/F3Q1b9OMe/SBA1qInwjHp0UPCZ9EM/J2+EY3jBaEzC5wNPH
AuG/S3DPrF4/5xanYaZ2WFgi5bSkHlqPqa7ThgOPruLV8h//yEsaXSGFjfrhuByO
wnvNHUWBdSIvzAxZq1uDT9umTsCdC8s9E4qxEiw2PG0pVLQSQrGjKKxNp8fuhRAP
7Ya2zlB68wW9eSrhUnzGs1c6Ei6Ii+Y6QMHIa2mYFDeSAGoiC6wTfid92alolYPi
Rkksbahe3XLG8qFzMDdileuc8HSdJQQQa2ADSNWa7dVlFTGtwbTz/4RwfNZ7vHBz
Z3eKDoYRacEFqe2vJW2k+s0DwknBcXOSpp2sO23GHVCTg7tN6+/0AXnEgI+fy7Rr
/LZ2lKRA1YXaZ7r6oiIN5c8nS7CKPBNXebWjoZ4BWq4JbFSUM98K5Dcd+ufhdLkm
064dGRgXSWaMGNNCzdEhIDP1KDALmS8WiUmjhMerDgWHX9Gna6tkyoxlKSRQ7afi
FFXccA5fiMlUNTqi8ixi94B4MxFB2zl7Uq2iDmer5WUoQ1W1rDj2Wnl5R8e93bfj
4mtJpZCX1cbJCvqiz5/QwdIze2B50gAbaAP+JL4vg905V2kWZd6sjcmqHKPQ4KpW
pCAtYXBG53j63oJ6ekxOeMg2JM7xbyJzqhPEMh59ZvQjIchap5cN/yWvUqdwzMSj
3loYFntJS1DFIkMfAcZAqkv5P4NsyZAgAQ646YF6MMAJpouEqH4FoGG5IYRVwkVv
e5ll72W4i02n0mBn2yxCierCcvFB/DHmmWqtmetX35ohk/vkkWCv0sTI0SzJSpnc
KgamcJwyZ/zJ/qtb5xGvDpJM7+z5GMZ3NTvKewez5hMGTIGs0tIMU+XITsjdaaa4
zYWp4EzAjs4RhknjFZuXKjMObXmiMYl9S0WenCCySJDAVeAIboKkwYIaHVYbbYv0
nuPK9eADxtfAVl0nb50l8qcJh5qN2L5xPF9f7vi0GCE1GU+YUHkspZo6W+9ESv/2
n9P0z6I7J8X9mBxUuOeQbMGLRmKLUMpgjTpxSinNmZxIC0Yd7xaDKIWcRsf6WLxk
8yigD6B3Vn8EpI0RQx4BHicPMGn70uYQyhJbCoPP0C5HvKhqW6zpU9xyp+dPAkY9
Yk4VxnIeBLyLvXaSHvnYz3ex2PbhNsrZbjLYAwCGefuu7Nl4Yniy1n0EZHxjexhV
omHcLfIxE90J79HhMsR2Wk9RIvHNF85H+9nnMqW22fgfmya9A6M456UR63CjTJJP
AHKhvSRkFv8dZGJ/BOwQUVuYjR1lqAPIeNM03TOZIkp/oZZbmYkENF1dVEmz2u+6
peTpioYC4mJO70i6Qm8UH3oVKNifKJk/eeNM+ovW9WtiRPsu1yn9PsREyY4fb9Ca
PSJtK22W9fS459c9I6ZwdBsuRAU68a0qZjGrUBpQiFtW/jHVGleyi/4HMg9XWeMu
tRhC/Fo4SbrmOUZGprEFiakFfnVQ+EeEpM0+n3H2UzaeisyfWbyQHPBsk9Watb+H
mFjUuUP7smwd/bo1uMgH0CLNs2xJ6S6eKPrUI4tZ8VuN2HFUCDv/hGj+3jZxFEcU
oIPNnFOf5HKU2rP9DpPosBkHGalntXU0qa0tcZvJ/SD0yiypfpyKB+I/eIIj+5ey
8hIEN9kQMSu2ubKzog1EbzRzLminYDUB3Mxv92x8YymFifhEiv3A7abz/4YjARpN
EDcWrXmLKqG4cTk1g6ssJ5QoMY+PAzjsli7v2AjBy41IaQHT88ny6KPNwzwmNk9f
v2ZmEGWK+hQSXQFFrwwbRh8yGquRytMKwZBCYMpT+drtBijPtVoAllDgyBXxPU6g
+PXj3n6DVcCYuiDo7DSouso/9QnU766BmxP4MHckaion2H+gI4dHPrYODT80tLjL
C6oeNgohUk2Dw/fJ/ZEzhNo4pXdSVLXr3Qso6h9qKwJ6JsIQeEi0tIgRoXwMgYPn
SNmy3kw4b54r988neIiyrFH7p0wuftDJBl/Ua2PQx6gsyOoMu2G+WhdZU7rMtFgp
39HhqKSdrx921bj/+dp9qdbwimK9x2I/4fZFItmFEhwSXwdua/TGETtWGFU7nzrc
1JpUmJydHHwkFEmGO0bP3UWT6FFT5sD1uJ9eaZsGhu79WeOQF1b5U2TfBtW7n7xi
btECUjFD1yWFp7w9mWQlckBBVFmw86klfDjGJKpSK7cLlo6ooqS7FwUTTZw+Lpae
gBzCoKfZWNPU9MFgOfkPEjQpBO7a7XdVESOKq1uB5yW7r1XJqK3GNsA4lfkCds1E
LaLfTU8Kf/tcOApFOC/t9dD48qGbO2kip8FebgEgqG+/Q3ZQ5Jk64TNNrG/8TWrd
MJI0HoKSgL2bOgHY3FeQ5GVc8hAZAAho3CV+FxxIV/b385pmEk00ECGYdDunQSja
m0AWuJ7SsTZSsKgJMJ0KKoGQTFP0SG0JW0156SV6NKd9oRIPgUnOPNCVAIpB/VCy
X4acswHoMlrXHso83xyOFBZ7kdY9om0/3RTC0phgxOWO9S+L/KEAHc774WvT6voX
NgEwZTwYggG/+cI3qXLUNL5LZjDpXUMgIiL0eqFZXNo8N/shaok/oE7lgKOAL3i3
ISPb26GXN2WEj6ZGIBhRzyOLEZvd8NsTAw/OHRKASOdQe7W3Gssu2oN57n+H5CiL
dwqIb4HVBxkWy6xsm7mpR0CO8rs29gbj1dITb6B14pY/8VkOCm51ymARDUUMHfby
y/uPQWUTw6mKKasWJ7ME4pKew0i5LliAZbLUwY3X6NCqk5rSdyJUmKL4O5tNLa6h
nHi8py2a98Uz4qGDpfVHIXBENVeYy4VUrFO8rtpv8Y891/4SgrUiiyTZFMANHe3l
tz8FTJ425IwY0XVT0J2Um1DIKKvn9a3VZQJLzICniuFetbHi9IjzAB30ZQ/iskLf
fzEnrTjMuOMzRBAOenXv+5iFFRAhdGQE2poPhF3Gn7UMb5C6qVrZmyP0AKDE5ZHp
hNoyAJjFIn0A7mzVl4fBcfcCq3gX32X8skmZIu+QFon6CiVqXn7w3LATcwDFALg1
NjwCPF4YjLV94fv1KZM+/oOWXgRIS/Nvg/em1mgRzXpywLwd17/vx+YS2fz6h9cC
XtPd79h67ynQ+Fbjx2f/8u5SPyskxln8sYfxhfXBqJUPtJzZCDq3ueOoIWND16Rt
tRrlJqlZ581at6jQOo3AlaA2D47ql5O9N8MfgK5/hA697SZ8GJzbrGgjvDGM+vaM
/fA6dnjGhiKV6vAcXq3NvXX32Mv25ArpLh0EL6mXjHxeo1+E6tUUUZp8MYH0rygP
lQQTL5UwaV5FktOildkWJC/JRHqoX3h++HJM1ztNFeSBpFN/S5+1ykw3iUe0mx/F
IAH7JiCq77ONCkPadjt4cLJt0psI7lmNfTUg8nGML3LA99EVX0S5S6AtaE7CpyZX
AaoZGo0EzDGHTl9FDE9lj4Z89EXTj+w4fNiS1xtJmS017LoBkX7v8KvXaP5hplHX
bYgHyKVoylwdYKPlUM8dXKNtmy86GIJJaOB4NpMtlV1vbq38iVI7oLtaKO/mwpJP
UmbuPAe62SGWo/qX5CfBw3x8XLtV9cpJkpvxauThhPChVvUSItpQT0FVFpEO5Tqx
waBA4MesU7P6MdIr7+KCRtQ/ULybVcWHDTICkvZI14waRi2/J/rxfnXFub7CVltg
pn44aIzWhy3PZkyY6TiWvEjaVOsBZsZcmAwW6ADev09NoHbtjbiIbP3I3VobcQNC
kBjzm2yuOh89u4l+GO8hrWNUlVbfzfzVpcXIrn4ihBB6ezecFrXSSPX0UrPj22Vq
J1b+D1mXWOqzGuBBV13vD3sO6vzmyYWyzEfyvUBnxs1wdbBW0gbaXmldHJKkpJDo
HoOMlj3X6iR9ofFEkmDKiHghiNlDhnl/w4vrmPRDI8I=
`protect END_PROTECTED
