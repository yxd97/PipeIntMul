`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m0SUfJQZbbRMRlOOoQpy2EPbaz0d3xF3Ihi3/SIBPzF8abCVTWrW9ntRKJRHImJm
oxZOuoIxO4XN3wtCrMFfmM9qs887/PemB+oDk++fgmd+RUZEbIr53dz54PCnjnBu
TPo4Ps6FgKWh5Qaw6zwu7PEHgPKUja6qOcsKheRWP61gl3/LDs0AVaxiPjSxIcpT
yqbUCyypqiuaFUXTdLJUz7pojhrlGaOOjp6LpSGDIi1BAfJec6Y1f4opcGjXiIKr
u/s6ngdy1VeBjdy9R6sTHI3ZZ2H7N7MrtLHHvUOSviD5hVNLuACXdKPKNpALcmRT
erBV2xdxElf8QGnT2BVIR1VW4B94kT8hQj+7ZhtceGoJwR9l+xtVylJdn0nRvRK1
4+RMHL8eYYTaNf6C3MjWNupebfs5GYlab0Qp25SqEtL4k0Ldi3rosJIYEMUujrff
SulH12MCsjbJwKruLnNYLA==
`protect END_PROTECTED
