`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvvE3sqL2ebtTuWmKS4t7GJV/Bblf8FLt7s0BAxavwFmlSlbt1zxSThn1vQfo3nA
cERLNULxpArKgAoeBdo6oCger9mF+OuLDpum/m36yUIX00xfKFyGxkwjr1uZotHS
kuE41l0LkixDVoM6FWJ/hvOQYJH+pDbRr60rvNGg7zxRYkvLdCWQYwfAUXjIOeaN
D3UrIaiw69TVlan2ykJljLRDijsDciZqWYzbyxgzUJOylFLxcSifekBtcVYeky7d
1LhG6QI4szqec7Y8yitZHctlMjdTE2QKNZ/U4tOEprD46hXFdoJ6wzuIagNt2bQk
`protect END_PROTECTED
