`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRnWxuDRaZ56cctmiqf0s2f+eoONp3dhOXxqfjpikDwOAwJu+A6y3yS6LBQ34QDx
N57t2tK/aLyqYhv5Y837emXt1Xy6V2IX6VAFD6UaOehb7Dt5B7RNmSHr/P3XQt0u
ddCFEOm5qQy7htb639AwafjNZlG3/X6mb6iUQgG99Sa4w8RAmvJg94l26VC/7+XT
RP8pF9pE/cVFIGlWcigayYQaC6jV3xjURgoK96zHuWT9I7XzRDUWwN6ZfX7UHe4l
LDs2bri7zJ1hmlsKExSgaRt36lLvvd8HCvcZFCPznPJTOBjly97rIx2CZCyeCauD
vRxbfEstdkekaNqNsWc5qqRYf5XRaVV0ThDozzdwLyUgWBylFBYN/HxDo/MUxiLz
jr0yE3G+EgO6P7ICJB7YEkM19I/zOyrQReDvXwxd5NKQ4QZajvxaRR4zrp4iJbqc
`protect END_PROTECTED
