`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsCD2ktK5P0Ts3YMqXlEsV72QS0NzJOq7+S1+OhR4TzwpbjlbAzvI9J6C+wjwx/7
nAOcXVd4mVT56L5DhtfI/BKPKgqiE0nDbprxFZ9HyldcuVLvqiQBaiY8zURQlabr
G3ojPxJnHef+XXsf3U0z+X5l/wQs0PBI5izVig9G7b1moDOVfq+TDdr79Wa6kms1
uyPPDGyk/cisBeoV4Ml+NE0V2Gd5B080MLIsPQkQKVY3Gs7uc69cgXfnTQNpf+0U
Zn5qNqRkQe5UKT+a0v8/+LmQFQYenYFiPRl5IfCtFnKzYCSW63ipdfbQdbrs9SCD
srstDb1/fwNktO4ToU1M2UdJ8itj1ddVc+QDstXuoi7YS47Jpe1EM7BgFUHpVYec
`protect END_PROTECTED
