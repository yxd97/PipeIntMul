`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yMlXU9beAoLXwju8RSSe2CLHeSdKC+7OoY79gDqc7Svk/p4DmIahIL4LB80e8eMM
cOuV8gALhbv85D/t5R/0SPyXicnxsZTILuJbVBBgC3QmNrTyZxTlwP6hTWKiuGk+
G5Ib7o7puU+hWYfkS38Mf/OxMLnqNbbchorWa7foq/7SiuWwEkWx1jdg5TmDF38z
fuYMGaJnUs2olwvZCzvpmOX1hJWJh814poLi6hlAwh3QqOCpbh/J+dAJU1dva0rL
cqsGv9adhbuPlUCyaX8Jxk7TIFfVzIGBPuMjNjU25BzolEkBz0wnQokPokriWSRu
tzfmArXKl4d2kF0X/M3McG8WCtnvWD7b+MYFpUOHpM/X5sQeU1S10PvATgxAZvbk
M/i6K/UNbDSq8APKX0k7u+FbpjCaVfpGmwgCyBIpeii37n757Q41htKFEaBSr+9o
hpXvFmusuCEAlANQq7rQYWEZNvQUBMlXOtJcfUMtcZbt6XYpdHM2/CRI1VptGuNJ
UszJMHGqmJ89naOGByQcFcg1xg+k0O81+U3F1MrX7SvDEdlP6fsA2mTJNSf+g5D7
L34OAj7qVBtMlA+a3s/Suv9P5VajVsW48+6eLATfNItRlSbGeU6Fk3TBB/yvIZSm
sTn0PEyUnrr9KGzJAdaYy766taFmEgU0WvJLCtmP+M3evDpToAth/1cg4erl/C/I
VJDDEimBZLdDGIHcy9ZMSgl7bNc3NyYIQOkk38zV6yVxcJSN1evA0FyPRMKCLl90
nqSrpBNcWWWPlGrChq7rVTdnYyusBX4yWol3lAzaGtKZxMvRRwY68ZM/Qkk8m5HY
7FmLwL2WgAgEBbmqouk0jHQtSAOC0ANYKac11VaC8YmgY7Sp63ixAjHDrr4ykFo4
43qz5ozg9xfIg7yH8FEtTZp6mYuU7dm0EnxUVlA36ms0875mXIX0XnvZgPl5pcAI
GSJi9qpfd8CEXbD/n71VNSMpG8Es4gilhf7iLNVC5CpIfFEmtuXn6wJ7iI2zVJXq
soh6866c5FNN+152LNgiOM+3PuTIQI2z3/d5zKSKbtgw/bOYTl0rEEGNFRYUWmy0
zJmc162wwOT5AFTQ3RHReGvuNtO5uQHGsac1toh/nIn/wtTu8i4Qpn+PlMVbzTAy
ZKnxKMAULkxaKK6oKTF5SuGUHUwqXZkNLyaCZFwpVBoJ5nhDoObsAtS6Db3GuN8Z
iCpmzmpstRGcgxNKke0FAZbkg08j/IbP+9cgwD4MEicX6LHxdla4FO1lxN7+sSNV
QEbqzBxyaSwn0Wf+JelAwRJ6ilCg+7k+6LHeh/tK/RxPazjkR065F8+DnDa/Cu+i
tfdYlxO3BhzCYj/cfxQCOVo2sBKAGSk8se8WvDJIPnFWaWGV/0WO2jQD+Eg9HiVY
X7R0wvIhmRiFwp+GAYdlIQQ6OK9FD6lpqlGZdAxAEY3gFGk/4Wm8pJGldvdNSRWl
UvlIxXY0TCEVYvzNtvdeCcRzhCURAJHbiGT3Rwrx2vyEffInugZ/hhzkrJMTYRW9
GFpM5FpHYgD4T1agsf3f+uWvNUSrMbXgUqiaWZexMrSc2DJ/U1FTmCpt+b1wsJoC
XhRU4H7V6GZa1nBmulRtavEQFMpWTKuwzGeru2fZikuk0UCfQZ5tRCVEb+QSvrs6
dZZ5NQ8mZlfTugUbCtMjlm1GdSjk62bsI2SvBF0yJk2n4oi5UyvtthW6/bjpTX6R
OtI1S/2VQcZ/wuTK65f7IIyJlvnNnKO4EVnlSrVdqMW2p6WxctX6wO3RWO1GfqNW
q+jxuaAG+EQ2RucxbyR+kn1s9uqBJlwcUMEjkB5i5+4Dh06efo3V9KnivI5lNXNY
24LjQyfkwWnEDyk70Ml7EOsYxT/4Ik04dIlhf6QMg25aijHBHpWi60Cu/sRKzD2W
ONxyeHzMU+1NbmcBektrLswr7UxddPOoWdkSq1j+aFqocK1IF1nwd9KMiWjNCcXB
BajTHKi3oy38B0N2iFISMYwVz1mhaeReQpU3B5FdIGWfWA6MoiL/dA1m29ZJf3E9
QVmdx3um4RIXQ7n+1Pt5gbEhXy0S63QYJ5v/5bYlRog+gLe5X5frajybur5tTOdP
VtRkZK7OxPDuJ8LUK518XaNgVRuYMWL+uqN51LASq+MsDONeG4xe5wUFykU+RYEt
P8CcGKLhya1rmEvRGbuG1076BzHVe45wQ1MqmwGyQ08rcwsPHOtu5/yBF+JTqMyE
LfHitdX0mS5KZJnvg7urGcz7graMASijJ2fQaQcYJPp1j9WtLaYC9QHmOrvFxOrW
CF9ksNlc/Z1F0D3/35/UE2JwpNPZO+voPfp2azo8iPM9/SwUQ9MWcwMOBGnYp1Bh
nmA0gRPIuX/LSTx67GsDJy9GFOvpSgFMbodK/ZbDcmiLL7uzA6fDKG7dQD/rUNsr
ILSIf3qIlocDMvFuGRbCrV4RG+QMk0tKTkqbyVZ/dysNjwWzUUL19L2EfWENtOgE
66nJ1Ytvykfzu5xzGxn2cyapN+SadP7PrxK8ibVKc0qs/Pt08aLMJmLxI3MDBR73
YfnbTroxB82ydOmWCm/xH+6SZNSy3CJBjPrvFcDWPCIGWuZFNxiycOYeTrNfBolQ
WCokG9smP23ziuqtmcnwEl2RXtM5pGFpEjB8yd0mYrakCNDBVF6UjNy/+SBM4Ms/
LXw3Ea5Z94xruvnI81nPjoNjZ18bSiE9pY7xP6egI/80ZSjqgsxrXzVIuNpQ/V5J
vyyCAMK6T0NBiUIQ4jLvVhIW3ZJbnOrpErtIIhCVQcHA0gTyWLfRLsoVdcezx6bp
Wh0JqHTunZvSkAWmUZziaMKcPf3oFjVYVo1jkl90aFolCq7JmPi4qjOgSBNPtm+8
Dxitk0/QCepeXjP91odqUC9P5gYuhvFnZfP6smpcWIGLAbdyMQSmgSWHxoN4hD+E
makbsD1ekfDxJ1BYRaeuQv3FKD5BGt5T/l8v7LykW+ILAvQH0tDT0Nu7sxdnK0Dt
ev6pjpdNN6mNqrbskkbW6tS2LU4m9bYGjFbGiyMF8gKM2XsWGtxm9HKvY5cM5fYC
W41k+akOT/3rP3L8virz6cmnqdoq4j/v5vOCvtrYsOS7PcjHXRV0Mk2WCORrTbyG
lYztuIskmx8H6xPku71886B20SgBJFnrVUBo6+AizIVxoE+YRUMIV59RUQ3/bqtR
60Lj8Ga41OLPmZUJcnf0rxghCpXp8z67AtLfHU/mH8g7ynr8r0QbRlOVXGIsE6VF
XQuf54ZYdI5GMRR/aTC/GPAgNHqJOhRfPd7qg2OcQL1izfh4Yo3SYAAp4WOKUfz3
5Gr6wnSAOLsIxBHoXU5plcVnpjJsT1JsxSEcC4HBBCOHE+BfAsFeNkWURwcayj5M
6lGLwZnakCNHqz3xIf3SuXWhRYBBe6dxLzojkUEL8u+rVxS9PKMTwG++jBUGazhK
CsHVUGvfSRh4KgD9vTVPQqR9DGTQWxcAf5Aj0TdYB4ZxbXhpvvFWkPtDY8sN76fE
ThhSDOr26rl/jayU4o4c1vFqcwQW4MUwUkkiVpjfMbaygeOevzk1X/iQuCne1P0s
zPLiS5gF9W4oEW+QHr0ViMs5hAwDknGlzkIO5OEyxmPGW/A/ajEiPns35dzFCF4o
jOOT/OmxW9AlsBjA9gA1uhCCF5BZERhtdWLaBRzJFD+ihEyBTQ2bdu1IzErVdxA3
OEY3KfA09KCAL/mWaJxFg/+xCZN/dzIzQZGK4YTc36tS6RFO1O2vLma9Vy3C58+6
uh9fGIEiWU0Hgix1iRdXLDI7lOkhBh8yb8B+ATeJpLYlzjZ/ZUt3XiigkdsnNGQd
pG5B8Z8UiVm+uvIQNWJxq4ZUV1Nx/TRluYlF2Ou4pnHyic/UBiHNUWak3KpM5rro
ZNzCamd8Qw1c2fozk2ibn5TgZBx/ebuayJKi1PNakdfF7LI1t8J/lLzaa2rR83b3
UdhUIYoZbYi0y6rTHUCciuPqIYD2qmc+SOvKiryRbr738k7N67DgU/I3FR+LShdq
yIvAOjJZTmwgxIB12Mk5EI7pLRC95doB9Pdbu8NMXdvsL976IDP2ESKonQVWO1d1
CXGOvZ8IG66rDc9Q0U2RWTajikALsC9tXl+KAM4mRaMP8ssHkdZRJbr6vBMXByfL
3xXx5NEKjg3tuU3xYQa3gC/mffRdrzY1h1q16lEbjBQllKuP+7JOMx6oJiBsEAgt
UM1Sgx3cCB1wwVdZJyxq4mUBKEDlKqKukvGZO6sLqVl1F+IkaSLlsegsKMHjevid
rokI5GYFN92mM59+jgQxaHLnqT9qwkOG6texEXHk768Uhubf59bFYw9M4uIxqb0m
JJNDIObTLw/fVQM2tYf2vbxRfXt0Gu38Voie1PRjnj3HY69SUOMVOie4J/R9Lp/V
nbl26cVAqefASpgJT26wl8aANovOJwjBlBrmOA2rDn4EvpTrYPSAE6cBF65/Rmsp
8ycjW0A48OCT0hDst9ryBB21MRRvnIcA85/slWyU/Kjoc+3VOH2iIKGz38DwEVgJ
7AsLFPuokoI16Qn7+HyO65tKoB2VCxvQKGSQstdpJ7Vut/l0YkcY9XFwBGA2G32I
CQ8Qg5YXjKDIWvwmVp26p0dlXmwoRjdLw/lniNwLMMK1zy3f769MbOAr9AJj2yk8
Go20hF5SUweTWpgW0JSX5Fmnbd2gT4DSxHIf+aRzTLWEs9A3u0Vqr4AmjGhTljSu
VB12IX5EPZfY6Rle120M3wJ9P/2PaqQ67bBsL9EDG7+vYJqhMY76LXmdPzHCJH25
zJbIst5gggCwCpc87YRrd2dm+rD3LXjONyw7ieynPcZlFl8pW0w4U3wwMUvwBEjs
8VNkQlzmIf+EM9RK60lo1I1cfQxrVcKjGP80COjjcN1JC9DeVQiLB5IOatnPnjFm
SvaGhg6iFkGZS+TLxq8DkL/LMUToyeHLqFAz59piUKA/+otnUXTF5xUGkcTF8qXC
uIb1/3uTb/RZ2mK0AjsnvTpTCw43qJxMsQKVRTj+2WxihPKoWuy782DZ1xN/VmRH
Rg0USu/QcpRrAS1h86PWHGoL1Msm3bBAUwfNt7Ey3BELCx0Q9tunnsQee3y3IBKZ
CDugQHktixq13R5y3WMxlc2T6umy63mkeAa11g0CnE110mHtzmDuBz14Z66t7VR/
CZmLPqaITzDxRcu77viubAM54WtnvsW3Y4uDvvxJXlBxuvNvYv3gQbwLbAEU5Hvp
y3QzF68jkGOADgOQJjpQ6aGuQtJekklVPtRT7218pcUWd0rqhjUdNrmUc7f5efju
Ub/EHlXFRVRR8JOB94otKWuaCntaw3ABFksWg0OlW1eu5YRImoDAw+XCHrN2wlUH
ebvtsBHHL3jNMIZ7SSD+62TXFqg4O1TICqJDg3h38LA/M51f5E+4/2rOmavnL352
S8IKgcAbf60JNqMxfFuqa/Q1kl7jHACLEWuSIyNdadmTlHVmpXWrfSW3PxM7S3gx
1P4hpiFsRxBD1sTMobBHg8ueECOHI6ijShFQi1pyn6pIfJW0gV78A4Y2QogPXnkD
5hjmSHn5wttuDoVIFBvN/FFsSUHdrlpHesAEqw7/J4SYEjnNFgjAGKp7gx2Jn4XO
WyEEDzw+rbNXTYva/e8cyl7WqYV8ZIBUR78HtdFRtWOHlCO9ULcXSHR2+uMckjqt
AF6TFUAoBzZJDazb9jqkCcDiCZ37Mx2HsLhqaOVOliYhWhg0Ygcg8KrM+f7Q6wWO
olm10HzGkd8B+L5KMDl/ejh6lxxP61oBj4OnRe0X1Ozo1EAw/tH2flZCyNbKWA3X
Ami9b+mvjIl/RzRlrQWnlLww6b1pOub0PGQN9vZnaOH3XZfmwLsROH+7ygv1xt6j
QKjEm0Xw7yeHSyWas37EeJIdF4D5+TqAJaq76qoxuzh/uxJrmKZtel0/7Kitp91B
IWXHc2SE6z90anmmpojDfJmCKRNLmiPjrJ6T1r2wdypoBq4mKEq7p3UWA/V9VXK/
3w/jnRDHDHm8U3BeSlKXeVuG4whu15Pb2Xx9BZgPiioN4dNiQ58yAoxdcjBiez6e
y5LpEaP44DZ9cmxC60xMKjxoVYL8mwTODzn+nc4+ZB+KuYtZhdVUwsS/HKBUdgr0
ivMaOSTKjuW6NojAl9vHKvr/tJaHnsR9AFJ/yFHUq936cSek/PBNYgCkpLGiRf+J
E0+irQWtfge2JNduZ9XmR/dHIjSVWB4eDIZZQ7ui7VRCLAPDENaoSpfyK9284uIP
MSRxsnHbPGPuVAcE8p/VZRRglbQbPpmNTISA1GfHSJGKyJguEFG5bmkOsKGrf623
txHMThak9WYsyEhx//o8Qft8n2RLYeyg+WcgCkLwzu9fNwBNm3rpmxUp43Hyi4sQ
4j8LxAm9jEn1bUNwApeVssKcf1UGpzf2m0Qh9fc7pyeVzpETJji6+N3KTzT5tY4E
c9sfzpM6RfkBNYXUE3696jrLbtwf6BLfH5npKoY1KvITuAaKZQ9otrSsgQ2FwX6p
diZpvyNpFiILnY3crvXfYV1T4BYlhYs9ehoFtauhu1FaGzYUB96HcPOBQfsZgPYf
uPUA1vfJiAC9w/mQeZCaIjEomUi3nzzNtTBWKOrsMaXNopXC76S804G0gzEDdr2u
L2SRSo6BVYVamex3WrZv4ngbue5qOKdWmgMkMgNUpTlE3WhWFLAOfHw4sboEU1th
WDFv8CEPk2cgvFDg8h6hJQaYoBJLg7mW7t1ZdKy92wtQI/4CHu2bJVYvFObuqgnD
OIp7yYw4NrkrkI0Eqvh+jcriBA5T4N5T3KtO0JOEQ3W1mBveccFf9uVYlzOAWAmb
v+SK3mVVleXmY9jsV7ueN8N6ZcosHB7PtWo6pI1gOM8M2zagHQwAdzCJMlnxmNid
AfzurliE61ppVmm8nUCOEY5mtLFJB0caP3vBWPe1v6ipczG9jMWRegP1ypgNnLdC
eNMiXQbwCsC/OM0Pi95yaFLlEPMZdoJQjVV90Qd80Hncz5ge0Tzs3Fo1dhSfLZOd
lKzXK4Q4yHSxHsMxdMMp5TCA+uoYWPj2KSiN5O7PyD7nFxv61dd4ufe0L3BCT1m5
MkAHr41iDE3cnhIeVHsE6ko8XLw4ql+qeP6iXdOs2v1XZhW9Wrzu+t8DIoIZvHuT
aKc4X2fU09e0elVf/OB+mwkVpruIDKqdV5D+eBwxDDvNbE2+iFuGTCeosNnZCgL5
vCfkBfd2yqBhKqkSQUDWkLL+cF9lMLTxOL+nf/ML3GgDzDVlRaN5jIjSjbpJUaBZ
ylMKdU9BP27HNySvf/lIxfLcX6tzLOeh5uXENi3KnPw6FS7lX7PZ9+9EFak5AuLC
SWJbkLd58J8Ry3WZ/e3K2JNzT7XQeCodDLXbLh348RYt+K4PTiVY+BYSoPuUAnQe
KdZ1OE8uG070DaRkcvY+IBZzYy1E1XoyDjCOFa5T0fzFNJN1AZmjkMu3NRCyD3U5
aXB/GeSq8PAdgPWxWzyjfrGa81tPVlYzVcDClW3m9GL4QzVwkdVPpdKwZlkList0
2Ng2cNtHSQuc6PllNILsH+kLb0jh3K3Bi7/R69WSTNcpSX2MCeuZDLH3xLmtc34a
pm5B9ph1KRkJlaB2uVNNdhVtezeTuGmAnMhIUIF5ot+RH9D29UONZ/u9nPovlIg5
MfIemMQkOr6soKwBF0h0zwQGjNiXFZR27OKuIzxVEeqOBeLl9KaxQIBz33UoLTtV
UFAbsjD175a2GBWdm5V/zLCsydOF4bh1kD5sK76Z6CnWZ+hNgx1XaHDtWE7aRBxx
oxQEWCAqu8Swrb76JXqrC7EoINI3P+337uby6mNZ7DYMPGmfKizvAftq10aezFLx
3ROmnEDMusMEJ60M2KoAf/gww5OAYeNQHml1uTEnvBT4SEDXRyrwLV9IXsSiydTW
X7mSqGxajHtTax7V5+WQ7HrEa1F9E7J8p/h1hGLply6pj8mpNMDNiIMp7KxYtkgM
1SuKHzZVq88uIsjaPAGk0wvTMf0SXPUzYzBWwq8X9Rum23w5DmUWa4czscAB/0GO
KHmkIV2waGcK8LpxRaM4Suad+5ort5B8v3MVKNWilfovLGrUFaPJe3hKSHpTlMYy
7zDae/wLyYdBYHj9qfPEE4VTcs4RfnOhcqvWUiZjbwo+DHYAQjFPH9KORIhB8Ri/
3cdyM147dtsim0NltUt6l2lPwaqll/1jAinXu7cVZkdBCCux/9FoxEm4HZ1dMbdj
1jcY/wC8FD7Z2wcKlfLUfOPbug9Dbq84QP7YRY2iNTKsyGgFBpc0bbPsINl4ZF+R
0NMXDF9i+h3Eh6fUINddBdSxr5YPiixYvDMNNzoO99Gw8TzYRRRGJTsUFWpszUDX
IJuShjOF8Toy8Olqxnrb2pLgrWtyuoie5ePByfScfXcR4ByRLIpddLGxiPk4WjYx
x20adRWi1A9WqhPqc0smw+zpAyJZF7zkXH2TwnWIPbw0jWpsrEvxQmcuePLwt++2
7gJ6wnRB0Xq46JUXbR7LPpnFcQuhRkLDwSfNuSNaSFa/ELnZD+lOtusM+M9+MKdT
ylM9F5uJLcB9WM9Ydn5/DtXf1Vt133d3YqwrGBDJyh0Vd43qo8jF3e/LVDFvCiH4
uaYoYIoQDIFNB6Z/nDqfzlPGUOBvjtl+knar5sVH7TWr32GFO69mYkrTUh3mkmFf
vlvKL8Nuqs5MgLfvmZKkHOSEHsySUDLFhLV90HL2aToHPVf3vi/54DVm3oYfUSgU
or8+8nKdy9LU9efuz6XAxHLzBWmdPwPB9tw5FcMFuKtyzihXVJdrLtosFiIf1Ps3
a7ZzwQHi8FdsNSg1jZX7lHFGOTjLnufPqW+KEpxC9y0XodHjFLCFtQdcy+RehNIV
Mq3w0ZsvKkGrVVbD3Kb2NssA3Ykh4rlkYcgzlm6ag+rbzZAHe7m9rlG2k8RGHPIo
vCN72NVRVWEDpqzEk1Fd83fr+v+rrhDg/sWLbmBLw3v0EqFfzlEVVeWmNJqwvQXB
UbjTQDEkWLTw4LmuPg6mV2Ouw5YXlvynLhEoR2/ZV6KyQm6UEp8NNAn7R/8rsJWv
KpnOc709RLYuk0i2eRd4Cr8nWDb9OwhCh5SYEcSGFcldTGsjCpisn29K3AO4vaB3
KpoeflxSmC7xtvCA1gNLlpPD26YXotAz36PkdDgHNOZIaJvYUCpOLqVcSFYv5yxy
gDNOhHFb9Ln5OYOL1IUOjjVGu8+6YuNHFajHY8maxHBF3m5miWnxIfY83iR38sYz
nPNEw1Ig1Qo8hmjFHw0YKjBO0nLRBEXMQOzTHIm141Z1Gvz0aHvPkr2VfPcZhhth
vFuyjAUPtfSwRd6Y1HmdETEAeJnKhmNeK6/kF3DozRP9ovm91oQ2Wnaba60ZRixR
cVxJRnUWSey/hpBAqnY+OB5rF5p5Ckrx5aA15JXFI55Ie4XRAkog3YA9bHRsWRl5
rYCvThdduBsFaB3M69FWhYKikjQXH0DGMzPkhuL6IwpGISa1Y+1o6gs9clzHENmv
j61qDjpwm/tfJYnOusmIlna+4AiCCqiMVhUfkm7pzSnGWyXkrYGqIQ3pozmWm6U7
w6OyX6guM5C+H0KzjOwVpEpSFcRgVO1NqHqUD0TTDYXOeBAPfxa4L7TViTLziHBN
D/im93Jw3qSmmlB6q5n2mOyC0LtzwwqOrekKk8xzcEN+edNbBia/sK1BxUmBq35Y
AoZRLkXL84qTiU8Z8Jww5XMwy2HQswsBhHZRB7m6QaDZD9nzKRQM5Rz4x3qqKSEC
HNJW697UWVfP0cPDSd7/9LYFIZZbFLF0YJJ6vi18Hw9U15TmWs3hgQZbWY7wTmVO
4PofJeUHXYLnXFp6zVCaP6a59NAqBQY7u9DyrBxoJDwfLjsIyoGyzkRc9mYSGqdN
SBVe8+5fm/9RaaKul9Ey0zg2iSapGmLJh/RomDd839PagTI/bA+JaumRVjeorlzI
Imc+WNduRR4/liHBOTunLb8vA0w09oi9tH5GYcP96InEbwNwbB+vLWHWB3UBN+x9
MHQV9jHUXE0W4WYVVSl6g2/cI2bBezOcKTvXTS3Y2n0hO7KAeT6x+BKVTdIriHxQ
MSfDPa4Q8Zv9WaBdqtZKjiqv4nhfq6stbCgNZPOTu1RKlsgpizZjG0d6/VvVuOXI
fz2A7I4P1XPntyM/hI4gt12VoNJa0O5oQAs52wmoU3Bd89zNq3G+ohVMjOdRxGWx
YHl9yIKQ3ceOlyWrHF/7045g5b4Bg+muhDEuRnrBinz6SRzndASXYdgElZv8eakn
/rUagWWFMMKg4nJbRlMFfJmOYeazl/vrWRrFNper2X2tZ+Iz9hjP6FEbll0lZHoE
Rwuh2jEXFZ9l8spXouz5u9QMBRpagt3VDc3F3H7S26hQisIroOCbqJddHvOYxuYo
xNVdmxljVvIp4BiTXhsQnblvm9ZrvNV6MaDUQfVjVKALchhCtxVKjX17LGwYVE33
E57/5jdrh5KW38wLq/ozKIk8scJPsTrJ5VvWeqHwjYU+dNvfnUT51Wmuu/vpq4Ws
JroYCTNNceBuncoS1iCqVH4LzOwiCJPJ9s24f4lsvo2bf6BwALA71w21qOvlFPcZ
TmSUIEUFB114x3fpkIs3vi8YCDcBowDR86TLLBYUSKVej9e4bjVxcM5zIlqUQvP3
rp9vi0cxiQiBeQWXR8WpIl/kxbCRJYc99+jwzFb3DwbdgUBWxWXn1LVlOGF7enFQ
lpoxiox1XpyeLR8y0B10+eJb0+jEKImNJflSTta2GegCbcowdO3q1hywxmAcLNo2
gB0QAA0DMScZfZ2NHtWl2SCMAp7L9uC4tO8C7HcqE+JEZEQTTl3E64d+/ezD1dqY
fZJFg0dqrfLAWHv3idcJLyTSo8MBaLIWonYGWwzViqEdsq54HDiFM/eDiTU1XkQn
NNhMRb9cte2uudhxbsTOWY1fi7TUKqHdFPjYc6BOdy/Aix8s0n1FZr7/cYDYZW9d
cKB6hZWYY/dzMw6p1BO7Oa4SsS6pvOV7bjYMtuB1abbuRLEa5eKkajWKz3GrPB7Q
2sfup+hVDm+9w0bRA8pHzj/EPRhxplnmb/flyXswFypbNTcwWN/pFHkhrdlI6mia
fcFjioU6TXAb47IULyMg96tDLnWfCsiHrNGyWVI6vuRsr7hzWanJU5zSxRuUqg5Z
ZWKJJYs7rt4UDAwdIf/DhcrSAmx/Qz2wXu+0re47t2v1MdqCGOLEti4T1QuM1og8
fR1ad6svWDlSSC8RoTK1XuxLPdIjNwLKpve1YwAnDoM3AOPqor0lecgN4Y51+JqZ
WlzNwrtTBhye9qy+9SvozV9nOs7PSxitki4azARcoihzFBCrd9sDTkis3RsfNUHU
MMJ1iwVWrD2pzjOOOxX5rltS9voopPPgPlwW1Si26cpAGlKpMK3kF/lxUtlW1Gco
YSi8gcy/I6Aa3dM6yezvEqdAv+Id0NCOgf3atPf1+JPO7O/uvltFhLcSeQpWmlUr
P/y6o/rNb5qIiVBZR2oCb8uFD5I/QQcU531VBrEtVA2T4zXa284bH/Yjfd33flNx
5bF6UryngqZsF4NPv0b76QiyrJ0YXEt9dykHzZAY9bfNu+rOYJs39W4OZs8/FmoW
zW0LkD1Tf5C33tDKOzEr+pzUUhLnm/CaDx40F2LxoISvDorRgn5tx/+PyNQasQCS
sg4m8QSo1l5EAShIObydwybM4xzoR3WEekeP6U7zmtT0qa1CdCB6IYMumybsmxY0
rydctI0swrseGoX3XQRDElRHM6ca8Kw5ghE3HIflRDCK0zrjsJWPC/MRZNoGKi1J
DYA9GhqS5ThEKcfjbU0HsorhkMUn5tRo8Nzox9C1GOYRj5vsqmJk5CAQILmV7K2A
NI9IZHJ+PxjQJyr53hw8k583+pq1KwCZRV7du5T1tp8m4hB3uyvUBfJSYYk/5fnO
yiHuIA5Nu1Vq33S+WG7fZ9eGQceo0ouUYP0Y3mKr3DShsuxDZiRzwYMXi0JIIZaf
piP9RIBHRsnrAb+9y1Hl2Oah/isqjLvhbmXuR/o09kQAsZwiglPPTJ8t+PqoIQGp
2PELAIrWPFvhzDglXU1NY8YzqQ6GG5kkZDoy6sG83zuGw16lZkOzxLlL0+tX+SeE
4GDJLLGKWL5MjPCLsLlDv9jHlpCODG7JKVL2OQFVmLUJpM7dQTIDJLeVcEGjJ97E
dQKOtr+JFsAhBJKB5I35Y3hnySOAJzPJD1CZ+2Y+Btww4bjdhb3sQLA0dwF/Z/ym
lD/lml5F5YYlzeHGfAPgVlGf/wHoCWXHI+IH1gJL0PZXvX4NathKasKys2WemzS7
PPqXf0JKYCRm7O/SYAXIla/Zd2+j4CyiLbjvqAlcpTU4F7EV9/gX+0Ee/Qv0emgQ
Q4iaDINOPToj+vQ4R3UMwJ7bVjyot2KRSU8KuTQXN6419whXtEM4lDTKIl2+PCvx
P/ocm2QBeTlhSz4bk3wqH+FY4ede1pJGDnwmMAotCCC2d/6NSAjCsOk+UUEwH6g6
je/3If+694oJEjAKtLSjXoaAar1acvUegpxGLTvm4DsBDPbMYAaZMDlSx+W0bwq4
o4bOMVoeZiSL1fUeeUFDNc5F9fLpyDRWjhtUH4puis/eenSIGGzl2QdWwKJ4Btyd
+gbyDh6mTARXdpxnxqaTnIILaDMlXetJFO3kz9rz8n+OfmUULAT595mlGUckt9My
sq3ew1g4An48IrLk2p3XkNFbkIptRjUQJT274W7ovBlwjpHAX5nyvv327mD+aPko
3KkJoa884zgG9p31HjF9fXDUITruiVyH0ZH4un2zw9MshA/M9/cYavUUfysg8LhQ
xEVkYuZvW8z/s4FRbzscQfa24YwY5WhGhH2GwotZCn0bBs902zAKUlAeH1PvCxTg
ZXngHgZfdGXHvdXpnpwwpR97/Bl/nut9e3bEmct6ZpPvgoh319ynFf75EXGoQSqr
8Av6ev5UlnIq97Qo3xU7nX+5NN9NBxFyJQKW89IuET0LTleSbUxhtzToUFhshkqT
51h1NALxpuIYNGCFs1EVcI1ePxG0P5Id2pU1qbMK1Qwrbyqs5okxQ8MY8LfZ4Tw0
E7fyDp6/au01LBD4SALjSaDjIg+9AQFO33jy/0hXisipr7W78A+YYsILkyskrj7g
rVSY/8x2d0m1JBr9LjI5jjIVDiY4d4LndbOfVYOUXKbd6iEWM9AlXNt1ctYRsS5y
ss6W6N/gwfO4xORp5zoXhjQxnYNt78Hm9NtraGwD2ICi9TXY2RpJ+soPIWN7v3IP
S59I9PlSSBnLC6z9yBAlfh1jpj2VwaTOLk6bGmrcK6+Uknye6R56RZH3IO6AD8VE
6HjaRN5+GjUKnWENp0PmC4bqZuG77xkxTaFsg+R6u1zDZnwc3VOLBQD1On5/3X/S
bC3UynEg+BP2mHxt4yzSvOV3vYxeKcFsCAQqE259sOUPLNswNaifGkezTv5W0Qe2
nCYBHd7u+FWPPN8FyP2jQspjkOWR1CyLILJr8joxhsLGVwmluLcPy1iooJSSaT6+
1l6sJteM2QnvMjD+MY2NuniidvM8HOUPY/pVu1sWbOhvJ5Ke4TVG4ddRsmMptpTw
QiD5SX+/q463R/OOWJqAYCLE3QzAljsQ8ifoelTjrcxGgWYKq6MbsSu3946Nfb06
pcHPye36fp2ZoivcE+WY8WFsRTBEfY6RcwQUkadKwHCJ3uZvj7CQhsZm05fEHCaw
wOgUtWqQssXaBPPTa8jDBB6094CRvBTq6SHO3NokEur9ExKtrxDIxkk67wJGC0vl
FDRTO79stHNahHYFiMxpMRZl++GbGmh3csXp8fqcgh0B0BG5A/4z3z/+xs/ZZzvI
+ALan4WTNHc8fktUYNh/K+3r6K92FqTA56MTrhgwxWfn4Dt6xfnwHbYn2yU3Hb6W
l3+NMLyyoNVpExvU6LmYwesoKLwMIb63WMp1rYMsz9ZsTYy4c7zTG85qqi2Lvpxn
eFQyFi3cNPJYz2Acalk+U484hLaPzKN1qp1L/CklaWbziqpK1+Bzc4i21mwF5j0F
r873GxAh983E4E4G1/p9Fr6KtaPPWSMkkUH0lO0Uv/J6Ai8ZVSjHrfLMx9S6hEAq
CuSerBZQDGkdrQhsG9Do+FPCX61Gxh075qyb4skI50Y=
`protect END_PROTECTED
