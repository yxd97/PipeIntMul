`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZYnL8ooOqW8BW+brGcpi5oEL2ZnLl/t+vb82kDXwWuzyh8CxVHKqiWV/Nhw4ETr
v5pxGadgRtDOty7ORPidkaMhW+VCZTJxOygIunueO+ceo9IFMbX2K64Glhmzcwbz
Rgq28IM3LiCoR/mi68vfScEqPbn6B5EWi+WzuyMlWWShjxzBOmqsDv5x5UdTx5T4
t2xw7i40tSJblVcqd3Gtr014lCxQSaDxF5cn696dnjHegFzZKspdyO4n2+b9PseD
9EJkQtiT+q930fIrInCNMZkDlIWU/+WsBx2LpalUa2az7NKbr0/ogUaY43hfnVoH
GsB82W7N+oyp0+oIxGst4LDT19w/vFqprzp6PYm8x+sLvrRgxd1tJBcZzqlhGYdk
6v+viUN/hkXvP+QhckRMQQ==
`protect END_PROTECTED
