`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PVZT2Vcju/DWSyeT3pNHPLVvhoF/fD7WKdVt9QPHVvkEQAreX400gq0dUrnNlo4X
yJCd+59TiZjkzWwjZrvRFP6h8p4ulXsSY1Go15+Ly3usCwtN24cJ6cMSnhae0LHK
+zeL909wj5L5PrSjdeqiwJclyF7VWYUvlKkatgDXOJGiTJ/y06e151MoRcgIbwX6
gdam0gW6kCRr3xPB/tVfqLJZAo5HtyJEfTee+KMkH9Lzvdy1+g6VP9sLzQy9p97e
N/eSQ/1epYNDSZS7TvcuwhEVuF5aN+l9HV6g4Ec4fyz8D9RLW7DQoNuz4sisTfIt
`protect END_PROTECTED
