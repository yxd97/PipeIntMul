`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnINnDOm6NVHKyh2OVUTUhrUvq0Qr/OoddiViJi8N1e33SfoWO73bMqmxc+FrnMA
UqZDKnhXFMc3zqODo2CFezbkXlALck3W4I2+IUSuyzFMhnn8TWTnvKDJDvSYYL7V
tPsnK/FMEnRnTAPXj0NyGRa7vKwt6H7/2CSTy3S5JnvRoZIVXMwgNkjFtl/rjhM8
H+ojGQ1GDDUqkJCfmFEii9o+8pq0OqtnRZ8vqFJe6znd+gNdduKnmEb612pkjT5f
xL+bOtZ3GfOX6KIR6KqIGrBdu+I4L7dFKslixID+NZowBdiCCyCqhbwioysNhBip
ymhCxvkAl+ZCb59SmMWc+GOpq0Mp6fl22FHA7q2KltVUB60rVByhLatPBgwJ4642
sEbud0VB5ufYFfQM8vdUuwXH9CBiW0HIlOzWVF32I/tEBtWNOPJxWKGKy9LAzyZB
8Jw2pCmR4FoQ32xbwURXkYQts8gI6lcPIyXL1eXcPAcknaVCKmVL37/ohankqL3L
vfVp2OKPtlJKm6YAEkGb4R0b/xS5UEzi08HJotRe8W0y2OWK8iZCoYnEtryhLhe2
GTqGcRO796nE+11oy6nTaXeV+qdvG/WK99WrdnHxCCjzX9vqJWL2wQgaAuwsbvhI
1/m5C5I+2GMkqzv5uhEFjg==
`protect END_PROTECTED
