`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NslNEmrM/a1cbqR4W+B4W66IcPrAyeKBsOqM3gqr7XcjLEuakRcvaoRfrbxUr1ZG
YEAkjhQu8o1e0nNrb+iGFnZF73f5PF1qHelnzmb8byZYJHWhkVVeHiRFA56nPXTK
wgh0hyjbNOE1mZDamuhdyjJjSuSWna2Ffc84WpgLyt5Qpymm1O/+vevInKRYkXJf
lnoz+QdmLEjIO+0eu7Nlcms8J/Ek3h59dEZXzCp/btH2iYCeHvN3/ecgNGcF0fqN
CkzlXAfAiz5YHIG90l64z6CI+1mu6chFUCYWMBpSqpGTpM1uZ/OBYdOtNXu84bU8
Lk4QAE1cWHgUQoDiASt4YrUqepz6gzEkXPaBkAa9t2rfiD0y3iuKKHMpFUn0b/wv
qJHhMBqwN6GP/fJlWAXmj0rKEvYv+C5UEAejK28JqeKqOqdfMYI7ZcNXRe76JJwp
PSIsHfs9qmxBn9CUiOiNbvN7GnwaYWs4gy3k+FvifKvZyfxDh1jQU6/Cwvsu+ImX
UaPEQt1Gu2xihHL61s4VQ/Xw9n0YblZrnAMflqwTV6BVavytRx1QiLLpw62rvpJ/
YREJB+06Zzyn1CrfAZTvyG+jVCp+HYXPDEyxs935O/L35omvbxRYYihllC4J3PkG
`protect END_PROTECTED
