`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydnGPBVLtpHQxY9tosNvHbEsgc9eIVK5kF9WjWFhoT/zw11E/gcBGR8UllmfZhyL
zBMEJG35dBLmkiQpF6pTB4f1Cwq2rMjDr/vmSdUlrL0ilLrmTp7nabugAR05MuRp
/hCERIadVTyFVw7LezKIy3ZMSVcMdoD8rjzGt9HrqNpNdA2WG3/1w9tJwUfK/E1d
zwoIXFrUNIEf5SfHhzxLu3/qd7p1YdG3j+NTE8COSiXFO7CCXsIp1f7cVohdEWwu
arxp6uRZWwdcpqbIOeUT00czFCshuaCt7jsD34Emo3qJXAGciUYdMO+qU4sLqaPh
4nVZNTVIbvzGCgFyV+rqQ8rsPsx5QcuF1Sn4LzSpFl83YRbW8rpL79USzvRn2i9r
zBl2DGHpLRx4vqsO1HKfs9suvHlGiNI2lsMTkr34mmuQk9ZgmGmt95kcRZi85XIj
dWP8fAMOMxTXcmLJUgYq5RsvsZxlmomZMhdvxxUgdWlqLskplNyHPXF1Q4GJsB1A
BXYZjsZ7eIBnQ5ph0rCSvKhle3/yP3Rsganksdf/QmL/9zYQDX+kz6e7+ej4E+jD
p1yEpKsEXM0Jbz72E2AujNBoVDfH/hZzjBuu7pUz/KEEodhSeH+WZIGr8s1a9otU
ZUy86j7veRJAZBrt8Rw1xQ==
`protect END_PROTECTED
