`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xJC2EbQ5x7pGF/+UIjavvJwiBk5o9Tdo1X3tR5ffqOg9YaBRcBXG/TicjFHdO9HO
eoKJ5wLEU74UDoQrCYnohcsUrJiw5wBzSZVXIhlByYI3S+U2FLsOJ1dOGOfHZHl4
PvSyoPtMmMNWhRIwndX+XV44REs2OeuLt9ovds2T72R6F2JtY/T8Qvak+6npfygJ
Dr5PDf7MoD2iVDxsSLSRhAugb7FrB9p+fUvbd+vtAaF9LD4F4Ymsn2n3gsmSN7/h
6OCZD3InZW6absFFa5tQ9qgOam+32VlRdWNX4zQom1fSnVMTbXxWjsZ0ASQnK0rQ
dfR+y0k89/bZ5jbkCoQdUF8otsKRqkIEy8D3lQHzl1Kxs/Iqu4NhbqiEcQUqDDm+
GU2lf9C9QLHrYneLgr2x2e+AKtau5Ybg1Ojr338SucuuB4ViZUfJ7eUSNlDPDiuv
Aca4Nufp0eqevwsn65wJsiCA+fKft5WkqCx7aQmkbz/OpB+lr4PdnWqxLy0CugUK
UrgctAeO97/1iF0yGska5Fe3j12z6IfVfFtWraKgyWxwktMi++5SF3v9k7T7i5CL
A5j+1XibXxtmn49BJDOvyQnLO3mIBGeaCHR5G/qypavWU/72l5yoVRO4m7jMs4lU
qKqnaUjvnfYwrR6hIPNp+H6ZjYT/m3WKqfe4lZJkSj8KN44o8KkH2urZSI8tNpsq
Th5+HCAwOjRyr++ehhOfc8E1P7yeAdMP3Xqduv+nIaBWXSNLQzGbhTk7wyd8eytW
60whVoHiqm8kuiLGBwFHPk9Vm7ETZ5lhleZJngtxL2SaGvQimwbqYqwwEJ8gbkXs
XtPClYbWLq4qjJ57cIaKZ/DNAgtrFxbrLbtm5Y04q2MDkkIn9DjMITaXdI7Iz9Ev
h4T/p+ZVEntfK7EFIhq/8oS0wyUY/D0WKFBYat94lVLj5dz3dLHjcek/c52knxLs
+97iqijmOb5wibDkAQuLS72jnAuYgQsnzGbg4+8KX1OiQdRhtH2d74QTPXW6AftN
S1Am9EDCU/B0RARv+fPzvfuICqsG944PqfVGtPtV97M173Tb7n81NTgN5VidA/bJ
wnMALGdNOCy4aTX9vvhsdjTfX8+2diafHxEvCyw0PI157MQB6PolM79kJjB2SB59
ViqcpJj1gbtsj0EomSNr0n5U13Z6blUTKeqhHd/KBW1IGV2dZmpZeXfAOv9kfM5D
QN8OuDOv5QSbdBnD+8cRxRAjrde2hElMexEbXFKYWLinJnzvIhYaHhKPkU3gW82h
`protect END_PROTECTED
