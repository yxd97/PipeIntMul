`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmLnXZKVCkeZBhHH2h5a6nN/dm+JkeNHno1f+3Rd0+woCCByRpv3/74DpZP/CWYI
fLxKw8VpEEAAD8gqsSFLKZqYQTKXJ+mLEd7eeqOhQcxIgIGP56rIlnPMs9gWEx1w
8UPoe+u8EnpnQW1ZfvpL72EtEkazjfMhQ19/S8I6ROp01RRhCMnNe52S8m2EJM7g
ejAIizyC8BpB6ASbjeegLKlupm/wp8xXSSCkhl7/q/VxBDDeXgILAN8qYen1Tt97
d6xPCVkJbx2LyPB0Y9DrjoGXZ+Dz3jjeBsetGYHFQDJDKZJQKLBT1hWnDP/ixNLp
VZMSILuvzYhhRL6QgyZCog==
`protect END_PROTECTED
