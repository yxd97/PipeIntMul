`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cc5hC35cW5LYTrrLuPCDZQsw/g07F8sMxd4Qs5WyFkdEgJ69oFzR3BdnnKP2p2p7
Tc2xT5sNQyrqI0FxguNUmfapqhPiHekk3lEcxwAVC6gFCgB5dJu+FsSmYoKOqhrJ
m8EOhBZtt6dZgV8/ip5filvT+Km8AxgvBHReXqfiYt1sOfzujC6RY6NBrQKFz202
YBQ0fFKQHijG3C0X1Yp4S8H5P/qSZaQsihXHxgu/2RTDMOk8moFT1iTXTsH81PYY
BL6Yudp0FuO0DtNeOuOgPNe9iRg59ZDxDQ30yRhsJO0yFez7g+/rZ5irUHTKfqDc
6fYdr21FzilqlSR8EXhsAE97sVSsNqJZdegSupk10oOcySDR543XULfkMl307sUa
uDBGbGKSmXkUsoz9K1SbMeZoM4Wiavro74a5xABBJqZvGOT5T8n6KxCHhA9zj82x
+BFFPrQ6ax0gHAxMxugV1E2sF6ityvxpqwW2J52YXoTpSzsCw8i6p7lPZDFmlP4P
pHZiWTVOTKhK9miMoOy17spgSbi16ehrDU3BNdIiEMqbMeGGVmBvlo6Xidt1nN7l
/xtQKq9dT7xyCL/GJqCGYnM9Xd3Yd0wYrqz8n+8YTB2Y+U2IY5Ygandx6DmEZpnB
ndp8/9UJ4ccGIDjtmH/RSy1aX0X7+8DgHhJHjDGq/DTpNTYCYM/dWSwZBSxQ89x+
tyB6Ma6rSbF8RG8UhBwGNUJZr2EFl+4WZohlve+VrgYLpZ8ONXxVURJtuT+s9kZY
QFqsPUPmmHxcnR3zfzG4SGwu4bIXvGguSbYbnV2AgWpX0UQ5gAjP6Us89kBO8qMV
BHSdJmSBkN/sOGE9cvIWtO7H3sot+ToLyi+vHvBUDcHLoheH1hd3vJYovEpWKgHH
NopRXEJdPGd+Dg3mppZILaXXHWy5Ml5BiXFgSqJsj/OLwL8rMlZu8ZZ6R8EXYmKo
mQA3DTkbHE79L0v8UFEN/odx+VHOZGTgATrMN7xrGYa8qGQA3KH7jb/WkbAOMNPE
5r8QwgwJKnpCoJ9vA8dw+C2/nyHMb+HqHPOH73OvPURgv5nDHx90mcxLGJMGXHoY
NuxrZj0mXjl30VnocUtAIeUUtxOrOuat0HBWvRY/8YFjkLMEWRnbX40E2kvjPX4x
1PQNLTBlVJYMy7fA1l/VJd7PmOnObG6MtJWSu4wlmoWqPylkuwvR3qwbxfUPyViU
kf3k5gixRrs9g1wz42ezpikssToHckwQwhpyJrcQQQlNAYci/Jwr517MxVFWtlUy
Ziw0BjHALTKE+Rua7KAmMEn3Jymo4xJ0l7doFAiSTrAP8IUvHGboJKsAutzlA3ee
8Nbw0b0Wgyh6ErelisfXHmUxZfShk0MjSDATxjY4umBmPMRxw+O0lwE9rEHK52Pn
GLzWXp7yzaOd/c88pZ3QagHWkqnCMsQZ0sj8tOdSeh3HGnK4WppUN86PhSsGqwTc
aMoWEDUEIZPgboiiBBxSPTFbxTWS1lc6OsS6n/4U+TWRv7s0wEMLfHPyVwnp4LPK
6d7n4P7rHdG0e+vnTTizbveosKB78GEqz51IR/gKoopxjUCpsaOX9EwQShaOR5aa
XW0njSZeaaKfpC5kDHB0v9PQapd6qwvCQBAWLoUGlhWdTAxZecSSDl07EFVUV4UJ
27ldBmJoSbN0Uob0VAmBa2Tw5qw6MqcEI3YE9LsVXNm+3aly8VY2BtB2kqYIeASI
7Dj0lc8XLO0EAmG7MvUQno5TmksLXMJN17N3iep0TxdvNxzUFVcVL9yyoD0nFA+4
FPOQ/wcQUMeL6nx0CgO4scAmJ/7F6IOzwU1o33s6Oz6Jw4qdy84kkX961pRsS0tS
N3oNQNkdLqrxhhbzO89elL7nNdSG+15X+KE8rGGVoJ+UGYPhDU3jyoIYb7xYYoxX
Ce8uPKI8m1D9ZUTeqDBrMZHsepuFiVsvhv6esC08LNU2iYsBfhwaNtHXa5ZHFN+Z
BdrPay/zlUoOC8IXi1qWrtIXlwoKg0q2IOqbL+tmQbeFLU3Uvt4ob536fRPrMbOZ
/3k2mAlHYC6T0nIhDH08xEpp+zaSMPBsHJVc6QVCcbN5ZRmaAyM+p9/g42AOoV6r
VwljfzIreCejTVAk31ozuZHdCymRr/Yk+4wAGDo9MDsH6m7O4bYROfOYrzcCVRyb
nz7SHVSNLkZ2LoSLHJOeSO1TlE6BmhQJYXp4ume3UGtnzOxZhzUPd9vdvQZ560UE
ymU+PCKevj8axfm5k9FXwkLLPLpcYb6UolwtJubsK7m4z83g6BcOR0BCKLv3dYsH
L6oqh0ooNkfmDfHwRVQN0P0nY63iLyz+EqLb11dI1mHfrxSymu3WsSwpv8M3bfc5
xPNLzKMaZKIJGZ8jSkagCKBg9G2+EmJgPLX3S+X8Iw7Hqb7Ch78W41cv2/stincJ
FErBVY2qXBrwO5oVWc0Ml6frudjd141sJ59ycVgOI+vidN4DJl3Tk8TkSSufA9yG
BXExna3x7e1O4VrYkf3xYqIRN5M2dtSe7oUPf6q8W9LRXBfr1ZLjdNJvUal+DGHb
bbq3c8vbPDJzS7ZdGBVdQhidWemIULgEhwlI7YOMK8kkgtPstRWTmYUx1XVjC3Ap
aHAwfK+kAtLGMujAThTI5V2/Fs/nfpW/WXgAUmy65E9O2zJccacHaxcwvKhQwATH
bKm2KPo8trtHDhmDFjljMIz9owVyyUrsZpivSgywiNPe0o9lXgXWW0KTENA2pIxV
RtKW4XgOw58DPf4Fk3zWr7zemqCFnclcW2vNEsJ1rtUOHbUyvukobzkgcz5kwLhv
mAF+1sCvKg/YOtyh6z0CEnzQYW+goQeRfr9WrM3y/6Wd+dOb4iKf78rhLSqEj3vW
HLsv6qHnvqauWcX6krXZK+7QETCOj1RzLCl3XLrqA1d9Kqw+0devzMbnV+DFfFDm
a7I2NAdZg6Qxhk1I5xEpV69Sdhpgw2eNZ1BN0b3sTAPxpB+Fl0wryvus8PXQJMuJ
W5seUbQC1h/wFbIdSr/JmYRhqQ2Q6+9uc/YqbaRBi0rl6V9rZ3HSodnuCbqHMBRe
upUzXj29EYYR6q+WELy9UX2FR4Jd6EvYVQUsmP2dk+V/M1Gp15y6sHvk7UouDeRP
ZUqb6BedHJVnSLiX6DtIrghPTajvOfjY027OqjOCorUECOqNadq1fgl5HwhgUdSp
bZzGnp7l8KVY42NGYC8utC9sCB8J3T9Butvzr9O88gLaP8oO1milJNpO3zNYkild
ukODym1WOmjlwTiZQRBmxB11sBLAk2uqcXUMsxSZB0cdksXDhi05be9AWVakBN8+
P5R9LCeJ33BxQTx9vUfxTYTnG5QV8SxUp+PX2rwGNuVaUc6jGC2uwsGiRgtZQRuA
3i+5ztc6Ts9Le6oFzCN6kUoXjMpGjJOhHcN5KnxNFbNqPBlM06+dUvKXdVXKWIGO
XRx+RD0e1iMssMmM2RLyrCLvAP8Tdne7QPZsiuJ+ghFux8BCC/nI7KuCMYkFg4ok
ljbzjNNvpcXUNuwecm60qTQdSV7oJrLkLbtZVT1Y2A/W0YzvhMgFpI2+6gFB1YP2
7dK47Cz43YC3JDjmR3b+qmtiA0ACObtM4YjS26WtsWkTBAaPsIaoXDEaqWiOrPKk
KSEnFIuUFXwoQD5xzyKPjTlqTLuMveYeLhHmfi5r/KmUf9fqs/Ptf9BMVh7XA4ZJ
FOZ0H0sY1H7aglAKIGb+4uO4spjgHr6uE/l7sDKfFA+c68HLS7d5sijMEceXFG1A
ZEOcLySIJuQyM8Xjfmd86BwF2AN5HuBKNznRX9hzmQXruC5nWDU9UKMQVYfN12YH
LlOABEPDNaef1ENRri0VCRRb6s05kciWgRMLba81KdzatKzfxczsUP3ZiV4fhDD0
bdLm+Kbnd4jm7ytDczZSHRo+Rrqs4oMw15lr/h9U7wx94L/bxGmqu4U6keodjJUb
hcTXff9fV+R06ObkVy6iC9/fxtz/l1TRJRd99ZoRIDm9iLdB+QJy7rPS7sWbS+hV
2tpXi42EZpEOHbOX6Et+/krBYVStCCeiu9ilek9msojFaacv8ReX5hBcSdtUYyFn
0h3XwC/pirICPmq9L9q0I2e8ujoFnJ8dVYRSOuC9wrde/ME2jWC7Ysmn3t1NahKr
GF1qd531lZo9/8lDQ9QpQE/sF8Ydpi9mWSt0NtZ2iIgV0gA7+7R4e3A5IprZUHdZ
T9wfFE0y9oL8SWXWcNaNG/gDis/OIA9afQPpEte33EmkxJf4o4VU3OtRy89luncA
HBqLtMuazswemoB6Uqe9zmIz58diZZUZ2OUPen/G9ORYsMyH7VohuvJojQZvd+3P
Y/JwMnoSvVQEFKIDax84I9xi00DM1GrlbEd9GddIggV74ZXbKg7AQBLG7sKZYucL
j8a/zW3DhvRWSpGN5Q8+4Ek+5ySVpGvcRzYMgqwWyvlBtQqqiDqrbg2Zl3Z2NdKg
zcKoiqlYtF0Sr+L25D5WgqVI1EEznohet1SprCtnsh0inhqpJTAw/yDdzNzE7C90
8MLODkkcbS89iPFMfgTxO0/9eMaidck8sA7Inn19umOpG3RWb8r7Cq/ZTJNlT6ic
FJg6kWlQX4Y87YaYURePPSqtM7JYP6LfN89QQGpZiPlOFPgm5Ipkcg52EPPqJcQC
qa53GG7PjqiboPwAnSO3di/EZ2u/S/fHvjnuNMAF+pz11oKaJlHyz+fVMF6Kkb1b
DB+EGJVyGr2K1QcX3gQEzjdbzTggkRU82+OGrTwW5RBR0mNBqwMw2uSKox5n52wt
0cgpQLyy4zNuMyqZuHcnQdZD49atzp2y2HVoWC1YPlo16S//O1u08MbEh2ou3WkK
eFwyntiHWJb1aFe1LdXyWZU9vTi4Ju0Nh3qj44f7XmVkiObYmHvq+Sw/pBowGa3O
yPrgY+VLBmxUYW1247fkHMF8d0sEznaygmYe78K1pl70YonWV1T870HrJn2aHlc3
ea+CyAJI6UIqt+CVoY772rc1rWtNBxvofyOogmhrfPeTOKvgRKxwcAslJH0YRV/p
3WLqT48vulcDLzhx34A4pJrnhIpNMR1DmzjLCCZpcg7JU8sOHYFtwvxakB24jFpv
cnqCk8que2ZcXCFop12tdc9EQoPYPVe4wnH7m7OU53O50cQSXieRbqPhTHETgFsp
V3gDIJDu9Qxnutufgj2RBr7t+5uJDyguM6l1fho0O0VxFoMZCBAZPEnHrg6klqcE
15bcbzGojkOhqhQQ8jJRcZbj5Fu49BIFyPL9aZVXeJMMk+xJznvtaJ+2bAp8u7jW
3+JDF2+0mH2TureBvF4+zmDbefRg4NuoTgAgrvCA3ZhmYAsMjqlGpRdfWZtwdghg
4wNwaK/BbuuMul3VxxUVnnIPPYutMq1tAeqZuNl6nM2hR1i50Un1futtznwCm4Ak
Ty9D9nQOU3bQMC4lzATiwftUvRGRkIF5/43vYpGoxR4ZjnQm1xoa+cVX8Reo5iNg
xrY4YjbT2FewhG/ij0bn1YYxT5dOzLX3rS7U9HoRJ4fcr7xjZO4nqJIARdXz4TQE
hvglNfnFwVpoOu8rc96xMUMO8SeUvbEiXyCj0+J77Nmr5xTG4n7lJJsDe7oLoJcE
xQNaoLhlVBwhreQGZ5YsKcOitVwG+qz5SsM83TBn/gzC6em4szhwa042iBk6UCtd
owWH+HTFjThx5KFbu2LKny2HhDtKjWSuq8zv/RUXTjB8fQrXsMLV6pMzr6vlkj0e
AWL242BdWTp0C4NtbJ9SrGcOp84am7QIg/7TLU+KbL/ervx4sLTLINOaIbisLQd8
OZ9V2kDibBNHIibc84tzQQDwdhlfy7zw3Ci+Hbw4AnN9ZZP3W3cDOzyxZvH/0bNQ
0NK40QFtoOQkKFwK9Ui9JYxH9yziTpl++hMg6lilEhBLPD97hoGilCA/+dvSRP6e
mYDml59KQ74O5GRqGkU9HSAR1Amw6g+bHqg8HJP9Z6wJfoRj8DqCeuZjShdND52s
/tUw8+4rmcp3/814yeKTtBqQlp0D5gMS7X/XksIlXQdyC6dPfF9dC9pLcg++7E+V
ghyQ4olTnKuUg7HVrL0Ie4DHeF966bf2R8hDz23qOM5XZcNYPVJFPxda18mo+Ez6
cIanoWwCRZ2fie+9PLv4pAcfWSiszo0DtLvD3P2EZ7RPhQF9J4qHN7YYgBaX5Ifz
YaZ9fUf0vqXHuBLJSI2IcsRJ7uCV4ORlGJ3aQ3JCum5AlteK/zYsrIf14q5xfw7P
TkR2HTzgeCdOogCPig+X8UcSglSJSwt/cEIz9a2Vyej07ABPMzAdg26ljjsp77Kp
du4RNBnmp0FoJRsdk308o/1d5/kvWOA2/r1PP6sTvhNWXUnsDy6Yf1czRag8SNA1
rPkAJgyNYdAMszt2acvqo8d03YhaK3DfqdZrmaqzTzc9zGEqNsOnOXzxFhtAWCrC
KHHIVNMvVXYy/oelvMlJv6nLE8RTHbxSCaK/CDDVAsh3531ZLupkeh5z5c/lnQqh
QV3TFlNzvr/ivuF2oZP4RGpMAcvJ6Hpv+34BDkJkJ/899JK7bLJoExm+jBJZrwib
l6KY2yzOo6ON9JElwW5xUkcgGCW3YICrKRub217yQ5DNBMIYAZ8H/zBZwp78AdWx
JP17PI3AgIIh1DohCj4Fo1/8qmNWWdHLuAYP62t2hpwU2ybc2t7biSu4na/vLUSe
iHhY9215wqQJUA9c9Ty09qe2TGiTuv3IGz4Lvhlep+kqkXU/E9iz/Ar7IfCuV7bF
IY1jh2+AdVk204BO5qQQOEQnpPncyGKbffNgiSRiw/pdE9aMhrGdys/WJ7Sig0lO
bYOJtm0oNt8nVpdSCMDLGIO3fyqfUOCizFKTzrP81gq8yMdG6bMNrN6RH1tvAsUu
ytkKUnIOT7eDd+1DEv8g0mOhVJPp9qdQ94XUTYkDiMgStYX2FG9RbT0GB4hzLmMM
rC9GOF+k+iIAVn58TW76AcSThzwg4kdoreFwh4jpVM8iMwvOK98Vw4CYL746DERa
zWNAVvsr1RTo537Buy395HpwRJ/ob5KFwtCTtYSv0LfWhMOzojfzv5Da5rcJYPRz
EJ5cBWbe/vbVaC3hpIZWMfsNKaizUe2sRTRLwt2JsoiJaNL0SldQh+qZMwrIWYsH
k0YhJhns6bJA/odQvTQC/u/j5xTXlr8VEdmcC/WmuD4gkiF6w9iOxQQcYyjJ1lUm
vSyn2jZvya1RQv/wlIgsCeB5Df+wYVg7rTbGMHDMqYyp8yHD2iSRRaF7LuwbxkJl
X7TLbgG1rwAIJoMQNQL79XDNHYddDo2WbiLzskZi3BgsZLiOig4aTVkwuWmm0ePv
6+7SvCnuZpzL/9dtD9x+8V/W/ys92KSwROTrMYV6jqE44qqgjBjkhIBwF6hrLS97
P6golMCR2ehaYoI1ssAWJTdyyuh+v8GygNhUqXLEX48yWv8ISo19Ht/3JUeDk2ZN
OMAGrDC8dX+nH9cIW7hCTSZ+wnEU/h2j0syCmbGjX6EW1CtVooE1B53auu7vIECV
jnek7NRqk/DQYaHn6xX3Fib61hipfRDEvjLh9N24Hq41v6tOsleFmufrYTRm3pc4
QEVN8ut0KH5sVMhVk4n2ReuXi90k2vNY3AJJtmASwYDq7+AcrbmLfwCRUOTriBnB
opQIs1RTeSbFIkBwPW8N+03CiEBPSXKc8uZ0DHvLd414euHFqe7nHSAywp1Ry3XG
ApJ+Aks/CkKkCSrv/3TDPqtLerwfX8T+uJySCngUv5dVfuPCT3j8Vc3w4qARlQfE
lQ4bwJiFyple1AZ48WE2L+L7miqiDrGNUS0kPJPPJ40tXHwXe+8hecNlhkQ+uwSM
E/LhxGj6T8zmujIMRYKjkjAncQGRM5uYo+UN+zH/mIVzzp9KJ8ckfYEq2kBT3HBe
sCwkRfVKjpc37A08owL42A79gGtDobVkNQUle2O2+D1HqUsIqsNbayImA2RtOfia
mHfx62BtNQoUMhDQ5LJiy8wd3xZf55ZoYXKlByGeVLN7ReHfbHvYgxmt/kQCbLs1
uqWY2IZkXJTCPbKnI2R4aeCZroy5qjBSd/3G/3Wq96Ttdeyrlw5JifCl0Br+XCLx
fZshZMdiS7Ke0Uythmb04M1J8ksIaTyb5n27zZdjjUjwzfcrWYJkXTQmpirKhdPm
Sd/UmT4kvVCkv9jmcDlZmzFq5C8J5KazaelS0hSOT5XlI10Da+yeGO5hi6rwH/no
T7TmHzTyO+Gz6OiLXAwVGc799EYrOTlDyMIbQJO+eu6KfcRadoazgWYCEOMmzFVW
erDX/4wpliORlmOaLKior2/Z9gnpbyquG9tGW0d2gEF8foa3wnqYZbjw3WOfgg0w
uwjHp+a/ac+lFP+1QuHq0bjxBb1Ey7z4we+zErC/gfo3pFq8gXQsrGdX7GWS7Vdh
VzOzrn9xuFdc2YxuHWdGfQbD8t+XgqVNgaeGArC2SPMHqqsDY+8PNnO29h0HcIFB
QT3ZGGAcK3v76hAVge3Ihrk8OAFFbqvhYWsMB1FarIj5fDkHgGb5oTMYhtlBSIbL
DcvKdGXaiW3dIDchTVvAF22gW2U1HxMMhw0ihY7EzTEJAT3qotPoHe/HvY26SMDo
6qVgzPlkhJeDZH7TMd9JEJqYBl/T3dS18KO/hcLw2OadrGuIWS0JV50SGlRzRY7o
AOGQ1gWsjrWkOEu5LxAHQevMfV6BloDx0dqWhsu+cxnzc9821pSNm6ihhCmeFTsJ
2NT25ZN4PS/g6pSgU4TkTmG4IeY/7nRQQOG+9A1fBLx9hNTdTquXmpcJhK0FUXoE
yhzeNlc47bflgtCvXVFUw53MNTmYIZSyYBditdjsn6ui3cn5bw71ze19S+99xtFo
/Lwym/8kb1h5t5cEjYTNdWyK3JwO5p4foCVqN/IlfDRreOcmyiDedgnmxsbW4adT
njmrYOY6Gq6T8L15JjDZW0vJRy0QO7F08HqrkSbva9yyktg2ft4R7VxXxanlGnSR
b/7+cGDDIySmuHoGn65/p7aN1dAhDtmkpW3yjc6qL00ef7y5ClqYkF18xJzcYvDq
LJX70wQ3a+yBmdKA5zLcc3cwqNt8nWcB3ApgHwBeDAMFuYcZk+6MBJmqAi4r1Kva
pqhv5xrQNCJU06F6Qeme8+9O0l6uL43uaKJ+Lm6CRxII1tz6sNZD2mGqDTvCUquk
C3Z8E45A89H4bTlMYfmiIal/9jeUsGwttISnVjLrkm6ST+bLVIhUL+VI4HBOx6Rn
PQQ+DaxNf2s4gORgIIFrzs1MNhgly1l+tWHfAI7/7E8wpAVrfkRPbirRCh/Yze4z
RLawiLeQO5i2VXnN3GWAIHYhE70e5ZCF7uHNbDS96Kh3Ee+aUoj2LavB47tSD8J3
cCBtKm74UiAfZ6oLyxUqgYJWtdnHjdc50fNTJ5uIl/ovrAamPec0/MQ85AK/HHgk
4kcTlZIar5p1ZM3hYSKsO63RiLDRNGEsQrWWDZ+9WcJNvcG1/NVIfYT8PFrCoESQ
REhhuyIXg8bvZiEc9DihgXYtq9FhgySdwyc5F+zSPP/xB/2N2/MypTwkFLC2vNRs
xQ/FfO320AW8+MUY4P8Uak/1bBmxjie1sid2Rx5Gg1MDJAhR8QDWEQXDoL6nBSz+
lBF3I+hpLh/iKzla6x2cx7xYV77fF75XSiKxzsaDNdTxhWBq2lg6XCG37R4zUuwy
NUGG7NDqnyEQxJvomgoJWuTiQUpbuhjBaFRz8CYU5oQgidCylZ2Rl2fIFWpXbc3F
PTD536gJAqD97uY5/LRGNzpKrJu+5ASdCIkQkJY+HiG968RhEhVOqYId/S9frH7V
ukQsEwT2afbgcCGpPehUnacGHUmzL0TeMPKlVqGfe/HDHDd17QxBw2w+icz8q15l
1kUJetgc9KkSL+OpCj61Vmjir/TD07T2z8wuecv/1wD3duz5J+nkOTrCeDXJnEDQ
KMWHe2J8TLPCgZ8Gz/FDLnNKR8mI+S3tzFZ/1EdjFGl+OUPQHtrijIFN7rgYJy1v
Tp9SCuZDww00IGjCUBNp8FVyCg6D/862d7NUbGwv6sy66VlKz/Vp5K8t4j8n9ZBh
5F+SU3mW2qst7y6ZD9KxhqozGUVIR3guD5UBiQPQRcCNf+4n1U/ifHjkLVzrDroA
gAeeI4wgLSV1ZE4CqKhYLr+59QWS0uJBxVHjS+7lH0MmuCgxmQ607RtllfCvCvQm
Xm1w0gGY+g8EaLyNUyWO5fkLDEirFIAnHi02XCJzbjj8xmrPyscbiHJrhMChk9kt
VAXF17VVMme0Nr67z35898GLzWykfRVLjOzLVWfiZTcSQ+385OcYppCWarRzGRAj
C/aB7h2bDFHOGPmqDfI5sup8JwRyd4rU9lRXnQCxipzLIjEc9DjzJIaj1wHd3gjg
so5HcZnG0LUYYBBPB5p2JPJjo6fQ1iAYktPFN+A7rWzdCamydQa4RBK07eOvk7NR
Ee1j/BKPS1XufFuyie6ukSPOp2rwQIjadMqhN5MYpMaOazAk9BhdnWSzRhC//kyV
rvygejlG5+cFqB+cyt0dRyxIHSt522XMew/ySl97RIRPuuevq+MprCY79bMhkQrf
Ke1/TM62tbfwOPBRpTl1L4PawynaYZertaokzbbp3lhBL7Wh64/nZYYZYDuPveZ7
nLxZTCOtv0nNy6b2FSyN2eu/i/sjCfGQ4h88Y+RC08NQJgfH6OWngXNqVtkH7BYA
BstXmzrGlWf6XLnG1AxUEBxh4c4FE71PR/KI0ZzFD/pBfP133hyws3uvZzWovkfN
bmIvEzlI71UMOlmCwI1SazQqFXptNtFp9+V15+NgtKJcwkqxR8tFCnVIxHpz9M3v
5kEgDlX+zpTafMyRThr2oqH9+hl04SrN/fq2b4pdQSxrx+f+H+5x4Xc5E2/tTS5I
x+Bj7gZe9FYfWmkJxXeBD+eiYS9MJ9FaD6oTnt9Y/QEpDAi8cH7Ch5Dg/LH0oZz7
5oFBI3DLb8A/SEy/0g7okdtIizTWgbuMG53yaTpVqgER4F2ZNC8mNE/jiz0gtdCq
p1gYWx6pF+D47Rp49WF/BlOG+rw76u7sfu2hzw6JiW7U11QGo9j9nYy583dIlYn2
JQuyuT9K17wIeINMyvQDRXrRgwi4TbeP3E9lwSTJoT4+ANpqQHcgOX+fERxsawlT
Wwn1wmd7McUG800t9s5li62ToOExJS2Kk1vAQGPZeg8bo4IwB7eMfWzUrJYsLimP
Nd1SOehsq7G8y0K6xk+WWqvGBv34B77+3ZT4uYu1TjWaKE4RbfJgicfTrzo8FVtp
/m3qivnNh1itFZYtHeQ7hbNYh+Lnp49WVqBk63Gv6VM8s9Bjsd9KQfdZ6ExNFsyF
MWa1iXeI4K9h07qBs+lqxHb4pMQM+gpdhCxlsG4654pWv/2qGRzvm/pFOFQagEYp
tcM6eLC5xWb0/bWYJ1AD4DmQpXTbds4Wq/8WSaK5YuqaAUbavcJe/QjMV6T8YCef
t8+2MmtY6yvV5Sy+kjHSXxjgSmxAaKemsUREtHUWjz0qWYhgzmXSbsI5O/ywqcl+
o67HbgMcT4InDT22JeDpUOw7iWLAwWom9qR95c7l6ihyZfRKJZNwj/1v2oG64CbS
DKbO74j6UyRY93bztXU1fsqS0UJpcZIrAI+Q5BQxo668AFS3VYF60ME7GaIlTLAB
Pba5MkNJ7Be+3PGH3NewDH8OF649l0QDrZoAwuhHJOsWfYxPUYz6TT4tAxRpqp0F
mEQvgMaks1A0MdFMEUajlH2OTAVgppqxyP328ytFxeRE9NG5EHf5J0l4EH/KgSW5
SBrllFJF+APp8rLuVrfFx4Fi/zFuWMjKg1awdHO1Ox8mmKFRrDYT7ExA1v043sah
wJp7m4G+a+ziO1Eov0CJbilRMF3ljMdSrSMLiPUwNqsAMj0DWzOFEYSBy818FZ0O
xBkqckoFHgnZNL8CkWso64NcVTIfc1wwV3eUJjLhAx+OxbdjylBbpAa6TdmcvZAc
dJEbCStSoOdAJ3T/ekN0bBkTBAqn0wcuMHXoJCWTWOT5zDPG6agHlzHHdKHtojv5
NMFig8/9sqkRoUSEAsTFgR67xafggl5ALaqyNo+CjekRmbXvFu15PIzMEpXMhCbh
l8+WmptpSEqkd6k48rSz7sCUZctO41aw7lW474nDoJ3ir/LuL+KQuG5t7rKEJvP4
Z3HEkjt91t0mPr/bsweSt7c/UHPBWtHXkcNe3qCikwQUtNdya25BZdxQnNXhhUEQ
71jo+DZND5NUjSEhJd1FRewJtNN0sbKeKY7Sb0Fu1/kNJ4F/WRQ20ZnlhQawU5DB
wFOoHVSVS7iOz+EYdlqhD/4S7msku1vCRMXkONCwkEQPV76ALs0YNuVS4S8o7P7a
IAWnDxdqGhFxnqkQnKWv958ahU8gH0Y5ZQeKdYu4v/4oQtVkl77/E6M82SUVd3zM
p85qwDIJwXlWSXisCuF3gW8XIeIMsgSCCwH+2rlhcsomvJuuyhw4j6HzR9jP8Wx+
Vx5T47RQAlYc/BN/gJlhWllU/a0EOH8Nu21jCvTyLcN32D3s00WW10ZB/Wy0NZbF
sUvSh+oi1WlxP+3oJzWAcpwnW3PETbzmJBs097V7VulbUxvkmeQrNqh5NOAOlLbi
SUg8sEhoDpb0UIq5nuCGVnVul3k0kfwQq5wFMha94ma9t0ila6QfCghYSpHMzSb1
l7uM3VwJolMXCaJauQKWG4cPY+RqEu0jNmYgAq9gEefEIclkWvH9N03hgzWme3th
D1R0meYvKyDATBTkY7hrg8lXQVMXNCq2vShm7Cf7Gg5sju5Xe0Jclgs8zl2bb0fw
xWF/Lb/++eecJVtxZcxnlTtv8Xzkqqesw/5/Ax0SRmbj5T/Mevtuhm+Mu9hJDoZA
koCx83rCDiYGupwPiJ9FW0s4RQVQjcNbCbC0M7ErlCYskzFNERQwJtcHWAuWTyoz
QyCAvwO7WzvJssofBXtem4qr5bRBdtY80xPdTSizEhiCqqGvVjNzVJSlE11wmf2B
0DCQFmYm7V3rlaJ+n33ULnpoFnlngRXIetU8RgWOAHv9wv2+hU7JUc4fZ1852HgE
0gkM91PjNelNgQy/bVsSBE5HiU8WIp7dJCuehY2M2tx5ZQhZeCVKkshv6it8aU5h
TEv0mykJW/ezmjMO8xVaYpkXAJThEt3OhckFp1J7snuBIWLfCJPKUiPoeC96uLdY
krTPKQ+1YMYzIXNHXxKMjQD2tdfsqBH6dtRBC+GkOSOCNpUzbz8TTlwCDHspuATi
OHoDBaiVRWAtUC2NKfByL4pk9RspGkNc+3Q9QjxR9P7GqAaRGHEUwtXnfpVJekx/
0te6opgq10tviKvUrCwbhcwVhIUjpKdyn9iMM769XcBVLoI7Vogy1Okhp4UKyr1o
PZ9Je3SRT1Nwnsh5jCp0zDVn5e81KOZe8Oi99rD5aaAbiJF8OV0eTIM5VFS10f2L
fTOCgeg7S2YPEM1hpDSM493D175VIQ0FT3Mb8Abz68Kb/iZ8baVtGKWf7h4JayXo
DAIdwddDJaKBBXIFUq5ZE6NzY6jAxf29G5BfKAhTlPISBXMm5lS4ctZGxlLJg937
RO5mn1a82cE0VIf7dQuLuDq3GKNw9m2OxAKdX0H/tsCCOkOnWRepYKY3UkPjcJ9v
xPf/e5COU5NzI+rYpcGa4ir4547b8gzmCjnyqURtye6ChKdA0sEy5QUGTih0j47A
WXdJPCPKQwRJUE6Jc5XMdcXlmGJzjghJUGl29D0Iy3+PDyztAOm4mqiDExgTnmEJ
It/ulcatfsJIQXXX5byYVGKJ4z4+Qvi81epkjT7QtCvu37oC0iQQt0gbIOjiijXJ
ctpS0xF6GIvJFIjDvqoEgjgSCtzS9IPP8DACbOkn8TTqOIBDZyAq5BI+tCiI9ye+
HZ0hZsxD4aVOS1+sM5wJtd/AnXu3c4uDcjYW4A/w1hSX3/eCxIzJzFcXft7UEPhP
Y9Vp+KaelKUFf12lc6NvgT/6eam5MFhIcGNsr8Vpd2rvtboVCu5/DnpKQUSUTeIJ
dbuqpDmFGMubkZD6lDO6YdPnA5ZIh5ViQAmdX5CJfQi/zOyDIXNNCEEnmAJYjn84
myIZHSyiNRkoiRtOGektnBAp22btSXmQrMCQa2KOEv5LHNNcM9+nVSFIw0AolXtE
EnB+vctaEWPIfuIDfq/LVjHw4XZdpgOnTOu7104NUufJPE6ldVy6xaQC3pLdCtI3
KYHo1IrUbv/4tz92MTA25BpiyLWmwgKSr6EiJjYcXEzazJnzOjnRTgq79eo356zw
0zllRYgxgcfH0DcuMZ4z4HBhcqrumINr5lG3bVBSr7thQw2h4qJ2QeN3eHCnqRm8
fr77NUvOqQVI2GNxhUwCgc7zw1zjdf8/dywZXwesQ8JqGJuW08IjfthxJY91ESA8
0u70dUVMUjcM4GTrxaUPRxwwbMBsG509Gdf4UYyQiqBSSQC5894YMHe+aLmoDvi3
egLMqg+erKNevcenXXP+b+MHTbYctrok7zTKgqjwUBOGTgaonN7XNiyQAMYAbULU
LQoZ2Am/nQW2lbCfPQH4sgIJpcOc/Pec9+EAIC/RM55zoJ+myajY7I2K70+o5mS/
ov+oTlLxvxlApzYfb/7Q3/HPFq/yZAz4TRZPWhF+1uetxZOLI1HVEJ83bl8UNrDD
JnpDK5hV9pVq5ljaMtxeecZUgssSZZuGhM9uR3cpiVM4HEHFNWtGSYeaGc4ah8oI
CnrxcpJjw+24amRxxtysz6IPexiVVmy00JRvsUZDQM4dpKoYEnNlH58gL1mIiG3f
RQhTkWGwpnkqvcmhWt6RZoXw33ZeYfCkXqav/YT5UYLSGAbb7QLMDTIzIRtjAwLY
Dmis8bmz5qqXv2ZuVSsZQrOvO+nmaLfcIHYtG/TEhgcSjuGp48RU4YWRDetXDlhz
6XaDXKlK+NkpwskL5sWVlHDDHtWleEk4hZKt1RewjmcgR6eb1uwKZF29AfkOf3UE
zupBUjb7FOWYWN5YismMPwMhp0Qe6rTBum20h2zXlOiggQylMZSc1fW/h/OLucyv
EFHIoHw2gyTCOB9SexsTQzFNGk0NdwbVIeCmbbxiTbUnxTMDtO46U49RHdtCjAZE
zSA24nVkRNCqpMYNKRxmqRtQWRzlwa3XN2t+wc9VJLW52wzXcpcB4cYIBFU6aIXs
4kZVJhUwUizwiHAAsR3ZSFnpCnU0SI3u97eWgKf0BfO8pxOna9ZamgTihlW46scD
KKJK5eWUkHme7NuweltgUhz+CftgDlr+7+8TobQAhWnuhYNlubTAbWS1qALmxny0
l7r3B2nYabxAlx3XEhz1joDs2YtCfGqhBPTLlbG4ZAIV9WZLzOINMH3kNp7XKL9k
rYcaT4wRJegbL18B4zRptuifkrY3be9kizABXR9SRxFMko3bpvRw0PcVwcgyM210
mA1KdP+8lVY6uHvsbgAGI5dWK180g1CBBPSarOOImmA+1pB4CX8Q8cRsr/wJ51eN
aw+Rl8zGTJS20xWAR0sRM7/qUCPYal2+lzKwS5kProjci4x5hl6w5GUPyEBhNeJo
Z2sv8GXX3yuzH9d24iLXYM9XZBkXYXoLyKvhNJgdqXCke8M2KoMu0IdwLTtCDssL
xfinXmig3UWK0TQnBGx7Wt1FUhLhTPfYpfDcxIgE65454desyOn7jXVIwwGw9gPr
eVEoyJkzf43h4e4GnOQxC53PuschhWT3W0feMjK/Wk86QfpxJMTb3FNURG/pyqx3
sjOJincs0+7WJoRFg5ohzCMf4VClDNHNu8Re67Hn4qSTQMNxYAjBOdQsYSkr0d9x
ijs4qAXS+on2dNRDLGWKw1Z6j6PeSXulrj9Mnr/N7m27RzmTGJTNZ5UVhu59OzK3
uQUc0Xt35C3OxD9LP61mXke71zwGNYX6UMzfQAu4xcvXDXQ7GH5A8MM8OgIIdHOo
OZMxqfnsLYII0ocakWyjuWR5D3srHS8GR3+By7DJWN3QDCL4JsqMyJYvVI4FZAZO
T6kc4OBAwU29O0MlyvliV6z5PEt4pah9gsJcpAMz/yZYkhTMzCz29hTQrKkynrbI
VHytIT5WwEtJY2OlXDb4ambrxiDuq+dhT/One3KO2V9y97mRcxSLAuPyHVmEeCwB
v4VqR7cYG4j/CVC+omZshFB3lFgiUkyuC3uDDGGJ7IqzosJstPAGyjjr4O9ctJ/r
+wLekDRR3+jRCt8W4o6RHhRJnfQSbA+Km9FTC2LgVQYG/1NPjCoG/5kFJnIv9BGu
THPJmsU9f8JBUdFtuZOtkhvh+oeJ0WzolXK682TO0UOObHts5xQ1hKTHEIx+AWAs
xgekHcn6XVUPyEZFt9aAsC4FxUVUMqZjxQuE1DEwhG5KoOFyceBWlu6P+sXpRB1H
HoXkBOpslly3mLpq74vZy1wTK6nVvA3Gug79C1p/UaEK4nz9JC2q7Wj3Bhwkga0Q
i1PpymaAuUHIX4kBzfZZeTZbZGIragKkeGysjwmgFfSwwX2EEk6FA0hSfVhYI5Lo
d6//EM1J/GsbBy4ihhcLfX7l2DEDXcxC5yPJq5cW/d7l0NPdgyVKrTvOrvCh9p3Q
j7oCyTRskNnDpD16bwZ3Cwgs99lBS0WlQK6lvFlte8yiUZucp+GDhgF7KSLJqDzM
ZjQ9In03Xa3oPPbidm5uBk2UkJSmPAOY2A4NcJcbX6MdJjnDCOjRpv7q08uggDpV
xFEEA6G50h5uDHGqmMOXGngeN4RE+Bs7baPofwUR6VspiROCFveD0i2IM1NClC3o
KyGxl8j/naZ8JwLwMby9gBYKp2btileYEPQBOrlGXsnNIs/qY9XMKs3xholgowM7
g45sKUVg75uSH9NrOo/kIbDaim2zgFxb2PxYKavpN+47Yczo1ETEfAc8vkoKfTUF
iuTSvuZmqH1LEip0dv3ptAA0CKjM9FAl6Vr4xiBVL9eaASmjthjJc6sSvuCKd/gZ
ELk5F3a9298RaFQaosVX9BdY4HGdSTRLH+fNsEOXCHd0WSO/+CWSXpcL8Pp4cD9t
FLguAqIrlSffHMUOhqI3u+pty02IIvJ7i5mLonkuAeJ/ZHpEAuPOzTIgIamqQjMp
j7bkYh6kU3RM7THqG3ITlU81NP+LqSxPGxQ/XPY3FcTqANguudRqpZHi347ZLEHv
hZOggWnF9S3BSE0uJmX7pLduvnOVUY3OQLFJxI4263Bi/p4gGWJ/tA3R3hXzmXBx
kOmI6V/5LNcO4Yua5d4GzG8mw83X5Z9HvNZgH4LSpaVjWTyIUxu8FUxy4NDCqE9U
MfwNcjjW8Tmnx7WtN1jSWf6Bn5nl43NsMC893kxE3aqZknFP4zGbAiiTXLlYY/yk
uhYk/dcf5nv/h3/TsbqHomfgZ2T1NDSJRtEN2LZF/7fX9nsyau76rDgAgtwIqVP5
JB8MIUi4enOLVi73nM5QpkBYSI94WkhQn/l7Y3tv3dRHs8c+X16Q+FysM2MZp3T+
iEykVf7Mp4gXnM8QLgYO4oXuSQNrhSBkN5HM9YXFU4GftsTvkLgP9U/h1f/0YgGF
pPT4Hg2AU0isFB4IPYsUXfmE4CP0EwVHq/oETZJqXisHH/MPE1Tk3xeqWdHAwcO1
YwDSZ+IbR8GLmNkjYawyDPxyV5ICIN1R6PG0vrH4hkoHiPV4J9syj4kWQGeu0dOr
if6qthZZ1XiMIT5xrfB3V+dhGFVdQ7XCDMTke/m8zZZrK0gsNlh6D7++YtcxA8ZI
40tzD7ltcna/xRZR010X4syj3rhcGzf/beHqT2mEMe5BYUaFuMhgl8Ip90REOd3y
oTyjW4OivU7iwAaAbs1vOuxDQ0zS7WustbT6xzlLQ4KjQuy33/q7HAydaPBAJZYz
Uca25ndJkV04gbsyYTFId85BedOCLVN4wrqzfq41NSOBmii0v3DMLs4TYzjxNAVI
axzo5YcyUMUylXQnnHhcVinvORXoWhEr0MZPsObCPIL0rmO5s5S6uSr+PxJELlpZ
Gw4FCggTVRZJFSZYYSKHb5XKlDTzeDFh0dl9tIru1qp7uLweEc6uDAZr2A35wCN8
sPIV4f756N3fSLHdh0RuniqjlacDldCjg2MuYTfwuj9yD7aS0qR6RBxeoZMC/d3h
yt6OSZ+/Bk9FWYc6gOLD/kMmlMs/l8LFHH+FUQoj6TMd8MXfkRTIhmtmfEYOBCGb
s/i/bTXSklflyHRuvX3hIkPW5wFUsgJG3aWCeJDpSHU9LT8Svn/MAtu55/LGbHLG
6y56ilFWeQZp9qnY3bf3tfs4Gk8/9ItQu6cGSmxYrAYFVBoj3jHUgMUdb5mMyFew
C82o4JXd3OXOFfU47lyQw1lXc58HzgA7KsU1nmeFqxn5rqODMLVHeCOyfG/Rvv5t
31Wqzg6AVsrpo3Hpzn0MLRMKuZP8S9iWoFAOZNQJKlktfm6BcwwRykphGh3OpKgX
BjwFkkQqMGyKq/SdbMkCBlZ7ZF7HtLY71MjY+xKusaXDTiO+WyRhx3jpQ2wyn1F/
D43V6ygYTctv156ja6TNm+thLD6ZX8bX2RHWhXQr4o5q1Rd4f7E9ssIY4APQc6FA
iBkEyqj3nOkyN+S8Avj5EsRV4u5k33Kk8+J41eNkfZRyYfy5sxcMaNVAE4Va5yAZ
jU8sgU7U/un5NWjOT2/cSGzy1bspJFhkVyD/BHpqjguHsdOUw0o9Jjnb41gdw+Rd
Q+Ri6i+VKSItsItrUObspfNOkGzVgjQMA9yl+aU3Ejrm5qZj6sSykn4itGLnNp8f
6MM2jqcIKvkeP5tg5JVEDiIYnFor3qINaD7eaLw8M679529QCw2ToIJnnBgQwMq2
O/vV9c3ut9P0emtpPLkQNruhdeFjs81IK8WLk2WbM3fzB7/fZF3H8LAYbfsXjfg9
xuYFSlo0IQQModv22KBPeM7YYTbKwkmlLiaZe3LpZUKaTPaED3WPVZCTSDRkK5vt
qq8hxCiBG/gqpT9iMnM+ACWwNQ5unHPdqXrKJWz/ASwg64tvZxAaPhZoRl6GS/+2
SarLnJDppnckrz8C0AxtP0QUnyuuuNiuaa+31sw18gDlvvYe7IhaE7mtnhVwE9Vt
7SfUkPwsDKfFkTj5y5eXU6us5cH0hSuc4ASPdDqqelhJXcVDyWKjSBBA0nW4WEM6
e9w6RF1bjCQzNSOSTe8Lji+YocdLVE3XQZso7xMMPfpx2wPAsBgTBJ8Wfvzc4+Lu
Bb5mSLgDRumk75VNymQFGnkXqNfsT9qrIdpOsa0Nw5QDqjfoJiFUlI6fQzFqFY1Z
Rn4e1uY+tEkZ2oUJHePJoGUuNsbqrqk1mQPpHsxLq8AGkt769qOapblNcwnv/yce
zWEnqLO3NImVdgM4fUidmr0oheFk7IsSXN3IkXqTfTcmO7MInGPrpb2NDtYWM74C
qx336DNSx6TiI0qmyW4SRqOvFczMp4KvN2vGgoaa0IwEHvLxXlAr1Cm1SpxBr1Lg
tFHFol7eRMr1BneJTCkj3cWYo075ke6VBk/0ZpHvU3jZ50JUh3Tx1h6UNeLlbbJI
omOn81w1EdkEECTlH7C6xKSZyz4hY1Y2by9oPib/D9zXhaHU+riYjU9vyXlyehoO
nkFFiaNRlJVcwA/EU4Nm5rXBCsSHsjfFpMbg9DAYOHqijInQdlfKD4alB0sEaFMc
sr8Vc6L+q8bqxXKwkRpTpW9Mk49AhUDGHjYj3vXt9Cp54lfGiHvRMVvRpkSoIdEc
1d24T9g5cgyguf4SEmTE3MzUKAbktsYgwkXpeA0JC5iauYP2uHFR0Y2hjof2WaB9
E4yJCJVKwA4XR2Lup8of8Z3P63diJlyw3X+S9Jf7NJqarm/6gEgoHdikE9szQFtu
rpH1pDO3uYSziCUOKtG1R2uZMrcGNkw5JxRQlV02rjh7Ge03AbEaG2d5Wiq1UFhg
cKwkZ9qM6MHVaWnunOX0Ke5aFxhWu6kFxQ9SpV44nHaXAZ/v74KILNU8x0feqjpo
qnRTek4wIEtVENxwbNHuChAEJ4Il5Lt7VveuHbYgYgMiaHXivD5wu1vnHtghSaPS
qjvojYut7jWSQcwLG8yIaW+T9WUJErv7nWDZedvbS+lcjIyAQXu/mhUe27byDzpw
Ak0S6URRCHe//LpIkvjmLTaIoWWeajXZPat2VmQfPtWQEGxNgkinwFPmBNF9m34e
H7a/pulovpbgH2p50I5XbSsL1rlw/UW+JJv7SC4/neqBN5/iUlsH0mSF1TzlrKlb
+qkxG4qdMo8Jnfcak+3G3wN0Fr9ZO0sTxG2klHNcIgr0kY67J2E95/9E8yHSPNs6
llGnaX4hVKSPrHbWjamjIHXZAsTivOYUEFQmhQkYb6IUWWgljPqoSHxWnkji+YB6
MI80w35mqxKZG76nLhU3pzTe6T5wpjZefB1BJT7Ap6Eglgpu7AFTNUWdsz/x0PYR
Tqcd5ohciitDRA1HUYMl+eaF/BKBmNH6IeIyGU4Ky0OIi/zMLzQhGKBGxgfF3ZlB
ucGP8JKpeIrBQcPjmekYr+8VUkhz6D0BIk6DU79gOdx7NIOeyP/5mS+2CcVd7Rlr
CUgA3YfAoPQ2jSFQs9ZBbT9xdZWSXw/W9EmUsIdXJWOF1Id8C6MRozmTxKXCKahP
wMUkzrti3zpEwWzGFzP6mhgLCHuvDAURa/BYFBD7Ac7j2J4cLTP7akBwBO9u//9v
Jz6zh/IHmgS4Fifg6ojKxHP9rP58K5Gub4rG2kmFSlhVQx139pvGLIyeRsmWNUxm
8JT/hRXVBro12rxq8U6AumjSZaBFuFXsV4EyXp1MrCr1DMsxpGE0omr9qo+ohPBq
WnvMNJvBFN+vH+08XVVzGEChXnAQZO5njDSOyf5Zw5hHYq75ZcV25bMuC4pG1kve
zh9XnQ5/y1nyNIL1C51p1pF/LqXlJoFyVQ5qAf8/0FLW+Amqb++DINtxsHFWNg8Z
cs1SaE517MA0e0PrQTiyMAgqXKjkFnVfxk54+kZCILr4+fSGZKUmFcdLkwUKWDxG
ATlwtmSgjAn1+rf2IRygx7uRKTT2P4LIXn1Z10ekDzhSGoUtJjMN2GU9UFDchE2L
nPwwAOBM7Wy0hL9QtYz/LZlBNNwtmira88esJWmQ6UqYNEi5R1gX735L6wFUDrBj
GFht1/O2LTZ+ZXJN5wRQAeoAwd91z81bwB4/gTT3hI7qA3QIxv+HZZ71n3qbe9ID
wyUTfXsfH8PsrdI22o8fFmw7gnKEIdLFHX22hnOU59XifXZGVEHsIVmc73l8t1zB
cz09p0vBuk1qhCd7hR09021yhoZLdcMcjDpXLCI282gGk3U2xEaSxl08ZJG0+WAP
iZrKsj0LDXc8gVBZ5fv42SvJOHP8zvJy8Ey4EN3gQ0RokUunkHW3IqCRX2w/8xH4
ho5qn/sg2rIyklq5FMT1IxRo7WAuDO1uqhw8x89HxBeRc2ewF9jr5WjFP1UwKHDo
yS/ysA5yUX9yTKY+LeSvhES+ikd4yDxTAMdGEiqZG5MvrbXH2s2ejLeFzDoQsUoV
+Bw3bo6kdJHUHBpmP9LNMENPqCGBdT1o5yS5BWBNVnLaVTg/76vKk6k1onSE+bfA
J5/raNjmFg8iYmi204Nz62GSHDiuLCtGzmCIbQ4cvT88fZ8trFMuJMJEw+PiJCNg
h1bWM8AoGAOE/aWi5nONZQR1oDbfUarb/dhmoTQWksT0suYWRBvjEPoZyXpOqsVr
/LUVPTIXQ5HgPD+uUdgnApJIxApF8Olwppg1G/LsZ3O5eHzipMHcOS9pNyq5t1Xz
F7xiriU2Q8Rct37ioPmwskGoEazwXx8mOlun8oRBwQapaay8yd1gF10ofNL1m8lX
LBJ7ANK6D/7gJZCjvGz6IMEAnxpmje5hiX7SqLIPIYEEm3kB3TyfHu2KEnhyrfcu
GPdgJZN5eka/nX6KpoaoO/GqRDAs+nZoppMxmy/pDiPlqAurjiG6qiWlB8UK0kNn
0td4ytKdkMwzuzlJAuhej6aH2mlX/Xx98NgO5YHJ3o77Y/VoSj4nFEEVM2vwrXz2
ne6gn922D7/ueffUfWzDLB/STIe3x1P2lI3Z5zGeCBIFjYHSSMdF94CxrB7UDh1t
R7kpXIor8jg4wKH2n1cfE+KdL/tvT2iIIw0rVClkRth7wwDqNl+sJgmn4PNgbIo8
sk1RGJFj1ikltZs3HUcepK1vUNLAxYTUnrqZx1pGEqrlZAaN+RpuRnEaqt3w3FGa
37Q/7ZDjfZaQwVNTHMOEhUF0yjVDu/JUl6qSFCMMpIYkIBu/R7tw4caeghhvn6T4
iRAzQ6xS9If0TCcCPCqG7fMNcN0wlpjdG6iY3VWKAunw68rEjh0mRoliAaIKr+AI
bgsrix/9sJqW+IY6gukOyXHviZ0J2e80XKRq/rpK9S5BYrCSRSattkHqR5eSC1BF
Po76av+HlzSf4q2NB9aNvXW74febqlr7CkKIrQ7IInLae8mfob1Ge1w/oyxbWAxW
c/6XCs2uWuD2rMD+UXpD+lVvxTqNhL+h47j0X8H417FVALFMcrekPHz04leyBbCq
XwbVFFEvzlYABDPdW/1ftjyYk77BbYuuIAvzxob7lII91WDypDy+jD1ZeDEOg9d6
jOWk2i2dpUfhha/E0O9fQ4mp70q3iDRd2JN39W8hx8ZBWnujHqCt4YdIiFRSZGy8
/jvl+j0estE/nXREgFd/Y1Q9Kg+4tPNjFopF18nME8FHTYfd6gQ3Yv78v/sGh+cI
N+cS4MqBjg/iX97U6T6GU+6NAJTctI97n41hAfJ7d12KjujFgkz+tKU3NDerjhZx
EU3XmmQwgb4/Nu1Z4t+GbFyv+lGUiWfuehkKbeoRybzTaH2IUiAeJJNT6UPqOKmB
580/L5Hb8PNmikjl52F6X2OSEN3ycB3a6ca0bMdI9t2hrcoeVcihaYNa7ta6GLmq
7dRMjOQjLaZA/WJyCObCxKhK3BLUzZNukfBnRuZ0taLF/Z1kA+q5Jr0T0ShK9e9c
ho+SgVdFP4pmpoCVLg59wO56jBSa368acgTjPmTqAuKvKPVh4oFY3L9ymZUNTt5g
XxXh4tOKQM3Lp/CnWV9PLDDm6kBXUskN4hIqHBSKyxQsNpzxV1bPgzOzXuV6aymg
TwPw7riEZmE4SenVPiuLuIBs3MF4s9uNpJNmKWQ2qmVou1jtGd3k1dmChhpIyckL
E5k1+8eOeCkTnKzN7tjXNbL1B41UrAV5OKy/tCIcg7OvMTJKx3tXKJq1ucy3mrPK
ADrnpGHMhZaKIdEOB0PRqqBfMtw/u2IdF/wrhgut/FzEL6yaPIHGcY+mPCVKRi59
VW+rhS1Unw0YTYThWEC5lqrccey3Clle9iFiQOYRLMXGv0CRaqNdaGkY1yHbB2IV
vbt+aHY+irz8iV7P/hnfX6UIvZ6g51n5E4DDlfwk7GgGlrywk5elLckU5hn8FYZt
cV8c+/HJaZQp0l5iigfWr6CgAeumKcbpEIG4aQWlzR3wrM+OgKkBIprSEiR37eBu
l0rFGSetZ53D4A7S65hWa9FRIGLjIRwdDV4Tz0QNlmospjdm81s8EQ1Oo+51KDFh
kD+YyNP6baK0HlGoHwU04pUiA1RKj3sylaZrWK1NUm0W4Gcs3iWTSDpAOSHBpdO7
riHBt+ge9SVLWCMrsVWOJ+CjbnosltEGhVcoYjLuTdu3rAYmnaSCGVcs8VBFOZID
QHoQ9VJO/AIhFkiWTY6Oz4WALgXJDa/BCLMMFoCB0XhqOSyg4Qg5IwsghB8ltCGh
VadeJJnBLKgR53AuqrvMHrW5Q2hR2CjSe2hTNFNDPXas6z9ka3O7dwzPjQ8wOefr
GG0RY0OQw/QdsLo9ThHMidfY7sT29Lljd8ObsapBVL2WoXm5n4huw/dOUpdu6N58
bt7E7R+OeOkvTMLlbS4JXpfcYvVonKOJA7QI0F1ru3ytjwk/+TjF2no8ttDvrJSl
uxCHkG/ZCLjX/LfSnR86TJNJaxf8I3LzhK5tAyJ2NDQA/EyHs/t/YQw6vbacXDyv
UIdW7/q7ErXuTs/uPmblglw8bmrvrIquapBENMMbGbl4Ciulq1C2g315dnZVFiw2
Vw0nlw0I6ldVO7sdv2MqPUNVFdDaQP5OWWOnNiCP7RQYkwZK9Uqb4PokN0y9TxIj
IbNYRbGgw+mKNFWB5251SeaorqSW5iPAmj7xCYqgFLiVurCcvrP4N73ns9rkFiQR
/ZnCuQ/sMdtttwepLQzjW452de9z6NvZ1FEbfLT48mOjRIXAtlQ8zuEUJ1kL9Ga0
q4M1D06B2o4j06EnFgC1SOjtru8Lyzy6NbJIQ6tOvUcoLJbhgl/UPZdzboYYP8LA
vOX9fX/WCkE1WGRClJqpEPYdNX/Sd6hr41FqQltrEMlppbtOjRWF64hkdhONGJHv
XBiBacM40M2ASR9ZS9ZkcDFcoXr5dGefwY7jsdNAKZf3gTr1Rbl1syak+RxXYusg
CMHrz+pq/sn/B4l5j7rKFJGa+c60lhtSB6+PIULZm3mx1XWPCo+jb8EGtJ5+suCH
daaT9g2GNwtfuxZinWF3QHdYrBKJhchKmQAZ3DZYUFoDPiMwI7ecT1L+QWAlDI44
rh7SME41kn2S86WtmfI0m1kQ9V8mhbKrQQBCuhfSLjUH/i/qqh7a5X//x9CFlbAi
+6fkzrz/fW41S/FkvBE29uv6pfDCnKuxyx0E4gr6k+v49hF5fiORWQC6YNqFgDUa
pcTxmwMLM8pFobvS4VhJI84siyYCxyj0/7IqmjQKQMLmz+AU0we4Wu3twjRohj2g
fffq7VrapGXMl4uO7DC5Mz8vI6fUnIQUpRXiH2jIWXiAtR4G4ntGKKBOvoABKWLP
Yd83AOtaIsT26d6+DhPO/5cao4uimEtDLs0f5WAZj+8lu48FICEnW1VRTN5U8r8v
aVHGzSnNQtTfdwDcdt1HRBEy/k7LaXR+sX5XBHH7WrgmRLQRpqf3jf5lLnNDEs1O
YQewicN2tyqKH91qESv+HEai2ankzEdj2N8IB5wLcqcbbGiFLKJFxmDGX0bjsT9F
T0ICRcG8a4B3arCOwAv4SQ7UQOj98wBfpdev8m6e/8jMv1SmQ0c42tRaIiweqhQ7
9G2Goly7F0jbKAqTp92twH4SVctAB4oqp3EnCwkfjk/Y4ZvM9E+flfk4RTOt1SgX
6II7pRncULbQUpYJFagrQPfSgpeDCftsyYeG6y7HCQo1Jbvhe7QGkS172f2tFi3T
umKVwHlLDsaV5e0X+E3pvfTvUffYkLwdaqhGj9PwIzxBwdsSma7IWhdFpH3U0+cg
nLgi4QL8yVEcpHP9mwsq/pn2UhkVuVj0ycXkt8eaXRVwnHm9BtVheuO6sxhvuHEZ
JgZRFxGIsgowcDVtGM63kxDUbRtdcM+zpsi8r80iCxkWLHhXqjzfIMRAmp5Ts98y
oM+zWF4HnCNZWDY3X9b0t9bjd4i+TDYUiB4bx1jVhfNEIpXF404q1kPklJUp0d7a
0pcxD8jwMbREGcu4AVgTPLjSXSGL9N73qrqEgU0B7+h3Hv4BCA0pnKGwiFuMOlUk
voCDKRCSIpc3DP478ySPJiyz9XRG/mb3pFN4gQ22JNe70c1Ed/aiBslfoQXyqzdA
Kt81fsLz4J0ByPRzqATQd+2dz77Z409F1JBQ6D+bG22s5U/5XJOeMVtBRFM9U/tX
FL0b2UGyxaktC8jYravmJxNijN9TYmejI0IDw+TRdSqXHeeaUkqaCg0Gl98QLamR
nEatAYOAVFAkD3Qnr5hOXxYMF54/N9UYOepKf8sOhdBoK/uolF8sGBss8vAKqQlF
8Hq2gHNBiU89zqvezqSCtd2WeB8rJrCP/heYf8gApTyxZWQvpq44qmXY4FZR17aR
TT4z7Fzxsm1IXJTdqBptmpPuGmLVVgUbMimvwcoHko3h+Q6WLL+AjsMv5W9WnXCe
nnc91zcEdqf9lRj3TMXjdAL2RJPhamQMOHZbT+uc3fW3k0pj9rL9y10fesOhA2ie
aVeEjKnsa8bS4BMVVPjTL22pemureRQRvVwmc3XkVt99wyOUDYlCZjEdnPHNscU/
TSrgKaK24PBFkaVEWbIkVA+sNcaFQILcRXThPbAq60GqJXS84Eop+HBJos0MWT+F
OaeBjQhjca9s+UpcLWOYzb95gdc6ddw5SGerFeAcmziU1f9t/qGubkPLNc2ZTV1h
8Le/M3Hs9NQObUKN8hnU+BXeQVLMEsXXqxevomcBj28xP9BAWTPO2Bva2xxC0+tW
9fIdfz/cc8LVqREGlfR/Jeh7oJk19R/OPps/nd0yVtCNwU0AfLKhbdSfYmkYD6WY
UfQBtu6XGygeBzNpCrOrcCINe2gEzGzKOHljY31JvTgKDyAre4po3Pshk0zGaiWc
T9i0Bgo8sENSoNFpNAO9YVW1fbpmyB04I2flgwMSl4sWkYdGNEJhC/EsPHL4X4FF
MQhr6A/UNyn8qcNhS4tPuFqmlCptKpYF1Bq92onuZeHHREKYhtX7G0pYdSYrCVdQ
aPetbxVwWdQe99g/uOaIdcjQ5ASAy+9DFIngVRskcR8wSA8VGsd3dwIFxheQ6aG5
FvwyOuEgy7DXIU1tZ2r3e7OjxsOb/H5B+7me5MRZdXCF7LuE5TXAIbaCUnveSe5i
kxGEi5fFZaZhJjtU2VBHKxqIL1djbuCP2CkNkzbbys88Nm8olpa/qceE+7E3MH66
NGDmaS8niXRCU58GfyTR+aJz6A6Hd/jb99Fjf+9PhXSVYECKxi32KKgyCVIi/ZDz
E6HFmVArZiO+O0U2empdvVwzXoQl7MIPc6oe/Rytqo4Op+CFqVebhhWQj1D3YJKP
WrBV3k6G5bHF2waIGlk+PJNkKU8JCxGRWRWMB2FHettMyPxPd1h6QpDMU6vSrjCa
u9O0IX+UzYiVP0ADe2EkzJn0jMR2HSEZCMamr+9xHICfrl7ZI2BqD0644+pgBEBS
bRwkJQOEvvJY4jmzZQlj6Ae1WGmdCqIb4M9m7bf+TnyTlkOL+/8ejpEf27kpgyNe
FNnTJqPhr/6Yj/JvSdg1tgzKcSIiW9BNpLYhkxP6O+n6GVgHv3CR8nj0vXIUOVb3
amr4OWayyuoQkEUdi2c6Ug==
`protect END_PROTECTED
