`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6KcO7J6Bnu+pn+EzF5hD0b8jIlsFipLW4Zkc6aN6jJlIHlpV7O6O5taLzw7bUcBy
xJnxK42jaTDFFAxfwhZit8Vch/k3A2KXtQxq6TJWxmdWsETxhfSlqyBjQWTNY37/
3NNEajQACP5lwD2rs7G52kciJFQJb0K3fJ9E3FsqvPQJdpwYvfZFmPB7D2HXGqrj
BF3f1T74lGN+rZWrzlcLXybSwcp/iELEiCpUQ57xKvadQYFYYuPabmWJ/7Rcawd1
cQ3T2rqUS4B6/ZHmQE5gufA7ZMHOqs2RJDdlQGmiTzzXHryWcNcMyyEoSePjyeM6
TE965lRsQW+lAhfjP8EGIw==
`protect END_PROTECTED
