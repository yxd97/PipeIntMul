`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iqrq15LNx4yuhS9N8s2GHx2XFW2w3qYR5FZpRhboYlwV/fqz2HjEAWzktKdoj16a
hrYQfOjk++PvNPbch9OIMPWOeKfrtZBomA74rCqjV379xbj3ymimwdaDja2OJcYV
bnCqci1tKi7DFKrIa+pkKS/csr9St3iUYFJU1FkNT+ZbKaxBpD7VhP0dP/G55fYe
TUHGB2Ri4OJUlxHFr/Yw1skBtkJtofonSpBdw3hDtmXUDDvuVJDQhaAU2unxfQyk
+VjIjwMD8nlDYpfqI7x1pak4njUJhxVkSxzacvN1fMGpC4DuBjq9kkYR2qMMr4kA
XDjRlDIztKxm3LcpocC3nhw5l7RwxfadOlXO5l6RQBXF9EdD8sAx0WyC5Jlt9kcv
JBpf7NR1Q387tgdzD4+M/tdYRoc53mZCWsODOjvhDxGZLTvTd8yk8PTngB4UQ3AI
PEy1kqWT+c0nFd2xowLuRYGEP4Zeky8cFaasMN2Q++g=
`protect END_PROTECTED
