`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HjI/5M2kCMNFByzKqGt2JRmZmlAL8eqMhDKFom1Zn/fbLOvWajJzpvKniHMw4Mra
gi7iWMbsbbQ2nXt8I7GAuzk53IUNi5u2oXZucP+7ojJyb212u6XRrevQn6WLDHAS
uOnwG09v2mlDeUAEMisb0MiO00HpM4B3yDCfVcjRsxo8v3ehUlRMfq/Ih2ZY58f9
JThHy8Gq4ynIaDXDmF6gbNdXAZTxVNwaCwJ3SbPwxBIhKklJL3dlzSC1FlLZB1zu
a+Dc2A6gS6Ej0NCtwZEqtMLYBKBisWklHZlluUJyVb/4XYvjZM95kWxJV1v1nvms
EsDYZDPLVVsxKG0nMQ5gN97nNpPW2QVVxjewL3rLGQPyg6bHfprQUpQERY57mJCi
ErRzTihCtirOeH10CW7bykd6dRIR8nYrmcyy+g0MO5QudETqGAVmyi3pgU++bADk
TUHdSfTmJTTgq90lU55Tm/7FRrBD1AhZBiCdjUg8eoJNR5Es0qgSJ8PcemTAyxCG
TNqjD0GRa+jw4nnLl4iDldHCopQQL6nfQorRpjm5N7KgLhHBK3iGMQ+7i9snI9bu
9UcGJIkoLMTMvKsFWap5WRJL0M41RM5mniG2OBSUpgr8n+82nEPZLVpW2bJsnXYd
59qSCqOK/Xv/Oaex2PByeg==
`protect END_PROTECTED
