`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vWZciHz5cMfznOQ8w3KVNwdVDyuUHRJrtB9SVTNCRPxzQWRybAFW7Bfvc9ChliWR
0SRozNFNC3wM2PrbKCO4fXLffj+TPjdXsWuVNe4XYwfyJ07qG3BUaxFnUjTjJWbd
W09XrhT/29tE9cj3uVMaNznkABwp+VtoyfQedLOBeAfPjwhu8wIJYnr4O3u8B57P
+m00VrrDPM/6lLac8Og94lybR51vONI0ihh0KpkH7Ap2L7eM3qoWqviiJ6SdUrTR
caq0EptPLCY5nQ9pHn89kfM1G7YXJC3k/RqxKEMv8DPPQxXo+r1IcLugMb8gC0B6
5BFOYb+5Fljt0ePliFir0IjbSZbMMP/ZV99SzsUcbgHZbOgszkaFrvyT/GdLaoQO
4izK7NTgPAortXVdo4Js6t7VV37W3bCQwgJBDUsSRYdBUnBz93Y2FpDCpoyE5xpW
SKYVWDbcuNEfnFQ0pifwB3+UYcjdSFsZU6gpMR497hW6Q7w8xMTKv3WmFvznVSsH
hS/PQTKHuomdHVEWxXtpO0OKeANpXft0qm5DZ10gkSLojlNdCyN33vssAogirwqJ
tx9zYnIKuXuvGTq0QeuwS8T+LVbKTCjqGFG0buLAoTY52FzUUlApGwM+pm3jeElq
SlyRrM1i+mwHE8pNNgLkYrYT5Q3xgEz9munPc0PB/E36PKd7eIeWyqto7Qvk+08n
LyZ3+J6MgsNzKDDsmHNwz/ya7HX69nEr9a/b/RiyEsgajxz+sfvHdqneSKxAYB3a
1/Kuc5QEQrKCjm0vzGVstoN1BxBDr+dM6cvhilZRzOopR17kbh5sKd5aXhES7hq2
lMWkUgv8Bje5ZgbD6Hj2u5sQUne70Ms++S4vJ9HSBuWku4nPenfIkGSu0F6asf2u
EETjMGy5jb7FpfIpqh7hDWpMdgzNBpOQHKXYUfG3lfS0Z5Z1ekukvn7dHI9GUa2i
25rLiCxx/qadBh7pARbWsffMtL6/A0yAtWuXIkf0gmK7YOo7fdHhSza1enfzOuBB
9eidA7WS5iC+rGpxC/NavRLHsFyobTkIkDH19CgSgd25B4FAQEJuSbe3StpGJ5Ak
FKwMi92KmddszrzebkosbkJuxHpK2sfIAVS56R7x8D7n0uEpVNsNs/iSVcGJVeCd
SkEeAc4YKEPS6OROA/H+BaHZM5PYBbQMeWabz87wzB6Jf9DmMiRRDa5w1JSi6w1v
Ep7179Uv8QTrci8TDmxkjGRnv3kkl3kn6Q8uR+nkNOWtR18+gO3/w/942qzPE3lN
HGWFUkNxIbUuD9DTlEWA11t9D1KPtD8C/1Vwrds9bKS0j9+eDTi8ZDdaYE77hMQQ
udY/8JRalk423n6/tD58jA/ItnW/13JoiQ08DrHzCU/NgJkdygkG7KvW7dWRCxXq
cvC3i63ltbbfWnn8hXeNMpJVYsWso0avOgUHnVy1FN07NDbDaC/lsCooFxd4c8GS
5+MSBmAPOzI5gZuV4Cdhj9RzXsUmblpvOSD0q5b9bYTPyhDs9e4jFDXra/JY32N1
xjUAyoPNLSZj1ip692ilx2qPbZoHjzD0F887jiam7Nzq+qnK7g1hdRIiGERd5X5C
eE7SFZKmh7pNwgHEtT+Mzo85pju7fJqeVMGW4elLzjYLBTa9LlY8syAcbC5mqGCP
TvnID338F+i0OjfEPS9OoVs4MxP0uRYQM6kbf7by7vif1wPrpY8t0i2t4kG2OjV4
5sX+89mr2o+DKKEVQvMzUsPr7f43xqILfTKjIPgAlFWSiSpg7OgRT8cvUPZgEew0
9LFe+CCTp70pfrHVrqDbBz8EuOR4kIHdsiJehWxffxnGkRO1acgWz6JPDl4JU2LH
NDb7WJkjLLdzq/FJOqi060unqPZEqQ1ugKe2kw+88dkg9Dj6SQpdZr2vw7RFs6xg
GcMRrihOm8f5gCOwkhMYWedsjaGWgPjpq7OeVyWlNZ1/LftKQJ5A/AvUSLPjU2TO
jfcL4pI9ec+LNPWv/wiK5qqnY6ru/ntL1HFHKe07NgUTVsTzXEL3lwJkOY7Hndps
kLFZRseXLdoeHZXwvZsWGG/GJFF1+uf/jaZEAeYIcBaOlcv+NIPax3BeBEDBSJpb
w5gf4bT6Tr933Ar6FCVkPciBeBSD4UUodISAqIAnCnS414PE+1Z+eM/viGLPMKFM
RckBntPoYgzJj4UUgtzJTiOBGBZJyiJrwHmvW6SYvtcfUqvrmeF2Mq2XBEIVZp8h
+l2dGY/uvtRJNrT/YTIGmWwfUeztp4VCQhC33Hjoqri6d1qD55Wbf/724W9+xbT8
iVMsGbvq4ZsUqscyxAW251g26dvZUzhH3p6FI/y2+dI/rXxtntoHUFd4irhOPXgT
WOFVGYMUkaCOb0qZ+NIo3cS5+LWYnU1LeIDjEViBLFnKcnfHEsVC1UYBwNwrhBCm
AmP6jd2xZF9UJFBCn2WatBY6rr09o2r915gdkFxFiOy+vcHIKnE2kBLg7W06IhYD
a5jizlusDfK/AxTy99B+PLR+pqSR2xisN3TdYYKj4/686+ulErkvu8E9vQBTKgRo
WfqwyRQMPeJA4RJ9+zQxnhJvDvJfOkTVt2ociu9BJ9KOIr4WTTDhNifZHGCEKgGr
iONgGVjivCPm1ngIEiVsM4FuVnEwER4VJe1ZNq9/ZmPSRwqtROZsGwDIN0uhSNQD
ErrOfiBxlEu3QOoXbH2sNsmYzvuKZfH+UifO0uQqf2T9EL5gl+37HNdsUkZHjO4p
ce6qhiORBW1A90pRuG9pWQ==
`protect END_PROTECTED
