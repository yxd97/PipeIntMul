`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e45K7hniyT/I5pNZnqX2OXJbiitVuqbN0kLDw242/BpE9tQkrNwSHMZOHhA8gunN
Cvcm7drWLNG0F82hem90lUONmAS03ykSJ1zQwXuRvOXFFWgv3LaZrI2Jv9PVp88q
svcpjalzgXtorMak+WU2G57pU8gvjcUmPzfvOjVQ/S1If2FV6DgODfOvifwYS95v
1eY8ZjFwdK4eYXpNWGMosQ==
`protect END_PROTECTED
