`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RBWvoJkLtpZKVz1/6rnZHVK6DZocV0dldNbG6tN3cjtJP6ihQW25VLiqSdvNNklj
uVe3ZwuEqyLnvTvLG5KO+UY6U8pTf7F1lRuBeIMN4wFs5AfHGInwNXZS2NbQ8Zr/
oLFM4FkixHoL2p2odbjvQEjKfHoWVpQsCGPCdS8Wi44GFc7ttaY1Wy3VAfLFDFiY
E5X4QUEyAWAbGuk7ijZwZd0nMZYmfc6mg5qdM8J3kGj53lPF/3ZBo8HF53H81KHn
iC4u+bls1Ib/yeOvISDhc3C4+GMzm5T7ZqeoSh2B5MnRNTkKpewwVVaYfVSIBsQQ
J94dJt7psX6wbmeWqakwwfAZGMdKOGvAIE8eOB7wEdYZrsTEAn8X256dRSjQ+6K/
k2WcR7cLK+U7g8imaYESVLnQ2X+JLolvY4DmjQguNOg=
`protect END_PROTECTED
