`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fe6sR7hvJYWy9ZyfXNK04miz3gjgoJhZBMF0Cfk89nF3V7PHUZGahuWFt218g9+D
f6MxHMrQHnOA9SN1ltf/9d1aO/H5X23WuILkQYUxq5AcG/gTlIyr1VNAII+da82T
kwVIJsyOCdYOq7Z6RCebtU/+Xcaj2bMUFvgR/EsG2jTWOnALVwF0mA3ybMryJyoA
0u1IJhVMy/8kch3uqZjMp//S5cwu0UX9/53OGFXdKnqG/UKx6BYiJ44da4xmOqov
E1JDbWn/atLcc6XrOd9VbKYdEPxYAIehXEdS7A31ZMahJYQMx8Yb1+hpAyH6PTgG
fRklPJeg2ZMfac6u0GJTlBA2RD1ORG7YDxy8BXMK967+3qxIdbsgoqyhmr680jtS
+fe0irteup7CAD3fwaWhB0lATuRjKHdxE4MtYTn4hhlR6Adp2AQ+EOfN8r4ETE2K
LPvNL5zvMfxCTKnKevS6ILsW84hukaibc3cRoLCv+fEAknv8rNddI9DJqs1zoLNq
sgJdaGNz1VtQNy9muLf2PPio8AGmht64L56BRDeM62SKf/d1k2hplCkV61WRMZd7
FThw8rM/N40tSlvDdkaLnx71y7J1olpkqLJEQ+kor6PrLk5E/SdmdkUaMfcyfaTB
rhkG1TskXmdUMZB/Hrkzqp9gVdUi8x3VIrkP+SKOkcI7sVZ1m+wW4yzrUX0/c3gA
6wr7ZYi51wUfy8vrDtn5BmNEIsOlhv6qlwDuZU8YOJztgsulrOB1n7R0R7qKnBq8
WdVAiS7GtFWRK+K2OvgdmTBwTR4diwTT2t3q1V1ehFMxq7bh6nifcYiWi42Mr/nL
+7ugiq+LPx09yrJNy1nxANCqONeQRQNHAfkWVOvIq/pyG66NXaQ56UfK6DsLwL6v
ol6FHWmzjO9P9ccCSsnK4OVHvdCuquj1C4kqK1XwXLlqZiScIYZFHWpGCyrmN/d7
eAhHYhOe1KKFBLwWoAKkdMshnOwhxgbiLaziIAkV5fxLxF4+rcdkc2bhear7kLqg
WWZYaxBch4VOWQHa9DIq/Jq9Gdmyki7WVAeYEpZzJAwZO3vG+gvDH1bKS1VBMN89
oKqEJWQlub5J7vNmRlakhMBfZ0guiILCZm7zQUuyIkugAcEhhXeAf5ZMrJTypcmL
OIShW3tmwx7PtpBKAjWl5/XCPnHg4s+vXt+TlHokSy4s+bS4y/SQK9t8b6NaFfGw
Blp95ak8KqnGpIw9yWvkXwnfyReahVrn7rUK2tHemtCzRzqnnh24A/1AQIo/kChn
NpFqMEiNFr0QDua4OT48ZPIFS1X2eqgxFUCnqTLDD4l+DRJOVF64LREMqWLXrp1u
ficlUDrMK3TOC9J3Iw49WAJoSLerxUmkTdD44mwh+dt68sqbb6j3spt+EQ0sSC8I
kpgiQ26q0Oh3VibVNanLfYgnNIqbRMSCt9kCZBPt+RKz1ORzdBZrxwievRENq2mo
B8u6gT3G1c5rMO2a8+58FAG+j0uIU2kZf6jcZWMEBjPL0WpWr70vYri9TKqPb40K
nW8+H72/zgbSV6u7pIX0ELZb2d3FhWFqhoj8ln6Fb6o=
`protect END_PROTECTED
