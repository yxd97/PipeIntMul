`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fUyPoEhB7ykdmAILRqcbamfARXCVVHGPWudsZ2y78drEdkbMaYOC5+ccnQ81quZ4
ROY+3CD7nlPhL+4R4ibGZlWDiyy0vFuegeeMyIbAyYJ6zUz5MEw3GzPndsHJdSog
W18k3Bp3KPhM7olQRiimXEzpEeOLBqESI83pJxq6b4plHKgOA4Ta/d0Z86orFwwr
q/QxrDWYHlDOzHcHeWOFq9wl5g4emwgTriaGT/3EAuUvDbLkbjLaUh2tUFQGpkOx
DedgRuJKADKcBmwZZUO3mS1ggDpq+6QVzwZvg0d1ynTd66TE/7VWU6paugW+YXk+
2aI+/hliNg7e+dBwQ6d5rSRZ/Vba5gLMJIRIadiToj4CBGk9xQBr8uYQOajQiiSI
F1KZHSh7lj/QlagugCCMEPpctUwRIJJvc4cLVmLY+Ok/rpjgIo6I/epcQp+sD84S
uVFJetmPO8VzNYadj7t9ZJYovU2gYtSy77RhUDp6qwfKK9VOmc46B1CgmA2HUB/I
3pf5wcriX5VoD+NgRO3+Yy2DjWKfs6oqvq4XO0fyN4o=
`protect END_PROTECTED
