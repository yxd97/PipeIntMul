`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6BLPR3FHQfaiTAnYYaoj0GplmLEpUMh18nDIbKiX1i0cjbbymQrPIK8w59E3zL5y
/7xCNKEeP32bUW1xf30DWoUjAKWZa7byug0FMGaVxehvb/zXS43eb5zZjhM4ZNYf
cnC0ZlVmhz3GHc2ij105uzEYMTzhk9zxuXsOOEBdjDwtEDLdV7G/4you1P9abDHM
4odUGlvFzhMCbU9wGg4jFdWEKPHvZh5pq6sBicwsYXLNvDAHkcgGhBKF0m/fKdJr
66TkdjY41/HMBjthIYVaz/MUy63sHnSJoybL9Yx84Pr3M8/CCyN9oBOiOXRgenkt
WE3TTVADEZOZ8Ob0jvuyKbxzPlnVub6zd6bP93h7DYI3kXzXpiWmHX7uXeaRjEL0
`protect END_PROTECTED
