`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FVclKGulQwczoSHUp8SX5ddNKJqyKtbY3T6XG+L/NOTUJpm5Xw0+/UaEVzOyfEWU
ErccANbjoE62WnaQTVOHZSlXMRhJGyIl2eFJW5SrfvKEYvc0Py7DYVbAdJQRRf+2
fdWXGnywLpEAA9GFASI1fGuQgMQWz+A8seYIj5jkPLRJn+hYqK6t4gx4xVFCn2YY
2dIKC61/RA8/xBVN1MaOSSTaV/zpPAW7pbRBvCM6CURJXKEUVeS1M5ZYxnGlfSxo
GZXVY6OmHkW5Ur3V8QAk+P1/RX6PIAFRhTKICK7+lYToV3qJFhHftd8cNeuN1RWz
lxaJ8yxNloeCjwWYb8DHOA==
`protect END_PROTECTED
