`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W85PYtPqmTKS5jOXp+JRSfccW6LS9XOEl33kL1NVXOYDXHTeB+iNHYpuhwDOn9bz
oashinUARTGFL3g+8KuRf2ON5Dtt6gYXmpUEWbx2uZG0cGPyoyIMZvMP2ZCilhuA
oLrkcm4MMVriL0AvURe2dy+h7rOKOifHO+iIIh+M9sB1OLHbGJX/9IB8mViY/LD1
cThetJIvW5LnLZnl6i+OzCtaIePhr7/PvblA+x5F7bAg/6NbaT+uiDbf0TB6NhPF
LR+SwDtNI9Uyr/LGRQzCf+ZQfhEQvzWNuDsliC+T6Z4PBRN937fuWV/jC5L30dWt
+qKc4hPYllYn0u2QLJrwjIopWXjeWbiwXfFQjZRqOxehGiOR7qy84q/qv9hFLOLf
khh7O+95OFWXG8qUm8DSPaZ6g2FCcLRH4fRiWlQcd9w0C8oVi8NsdB5kD9R0Mryg
uJC8NmbKrOhntfn5yGLZgm0ZMBSm+mv27wg/DZofmqWUHH1Ly2jIeEfrcRNix1zI
NT0C4o6ulbTon8+X1HrWGWOriag3OM1hvE/uqLZN4hVwkm/orTFjbdZWyQ21d35U
0zOMTfnLeC7M8Ncq79R5RPo33xB98j4W//A3VEyo2qmkVbpXjbwyq4c7YJAmpc2a
6TIwZcP/LcFoA2W5tTG8tQdTtKoNfizBGDJ/M/XYSFpF/5oWLmHRL65fHQpngzT8
sye4W+MUtJH2636N8S9Lx4CcvXVm3JR9lbG6g1sYEUB9Oa3XntFGRFuZAkgtqvHf
aPmzLNH/yld13s6SrpMPTdOudY+L7wTrE8DH/1gy7UfeHMgQ5a0+u6+TgDU6GQ+B
ptxOSLjLYuvVRDBmGEO/JtmCqpFmCA+EJEQsNsLdD+GNj53MLLFiJAZawGK9Nsr/
Z0rkH/SqrggAvap6HRpmnLBi4bAOfvzvitZfB+7DMvbycofIAELAtxd6DEZHnrgU
PdDnbUeJxmS0l6Dh1vIJfg1C4UI7oP+30/QxwUanjsrTHzPWVZCs3hR8P5Hl2lhP
499+7cquQoL1DvidZ4+DG59ubK6epR6IbqHrL72hd3xc/nCWNWppKndfE+1ihArU
Zak7iKURQutDt8jR8zwqgzL8+LT93+Rhxukx12eI4R4zA0HLbJkv0jYgWMRxnCIU
VxONLpnNqP1ROS47crT4w+FSxiJXB/c35yJUGYnykzvWbne1DUSY0HApaMjULKGG
EWgJN28z/433xQ1aIwA5OBBUhuUVyAMI5KJAlY/L3c0S8VXkHKdwK9cMoxKqYO3h
Ip+Ai+osNcIwUkyxKLi5QMnyMXGu/OInEeDNqeS6KpKZVcj4yEuMG1SxgQhj+WbC
whegDzOJFaiddTx9uKQsVuD327mxcv+skTH4oj/rSXp4NsTW5iavCXwhg1GhzOFf
92BGtILgVO0ImDmRZgudONDfaERpDTtphRq9DWjlwEMq/LS43NyqgmnBzWWiWYQ5
qpFWYE2+RnkJYXuXBSvJVpRavdZqC/88QpSec0IPI2YVhVCBnVkpoFie0T+0422S
dgjWqNKbr4Y+8mCM/e2/z5Bx8pO3gPTYTb2KTNN/vGHQTLVV7LeyuW+uXGlBQ8ZB
q6FEk6LDnKaEAZ4LTxiq7SkKGwDu9isf12Wod6Bkwc6xwvqYLz0qkQWNpzYndANR
DcBfUGez366W7gqRtRwcxo8vAR1wddHSj8pvKw8rWxyeqXdrqjB9vDXJJcbPajEL
SsEluSZVrdk1HG9cx5jo8CQiokUdGl/HyOVtwfGt9ajHYvP8rW0236VHdkjDqG+y
VLdOQEb16+QnwBCvMYOYU2pz+tiCpXXhl+u9KerdR8HrDkg9sf6Zp+MiLU323GOa
zJQnjkmy3ZSXuX7WSCy7M7BmtcnlaOjJds/rMpo1ygw1o9SL9XpEAm6CDySWRaUi
c8Bm1E6NZXU7kVLYnqaKYmflnNx7jXMb8jh4d1jbhkPlNbzqtT5i6lGqwwjZdwPI
tGTcp7QdFKV7WdNElqybvItvgyMrqqWMEd2aoPKBjFYn2FWKJfyvoArR2m/frnX5
oTWKfb1Y2g12m6Dt10G8GVMzSlMT2SGNOcQXUI/sJTTp5H6pvKbmj7gdWMKNlxvA
9eTu1UwA+rPS06dNxIKmVK+fI87a3TTAbZC8bgxQ/M90MkdEehLuFrDWTVNgqYgo
AFQ1dMhCKOfwva9r0+TneT55nMSQ5kxI7L5On/PxoVeQTbMhhu+7BH0aR5r/KBOS
8xsZBWYKFKmYhJFCaKXCkSNtDr4MrXbRCDkom/EJ11FP2LOqik0dveEwTdJQnms+
KNjTfkVpjpGVSUVlh38/G/r72aQS0o9Ucw14ps/EJQSW3mn+ZdIxf1Avls8WeSzH
LCdfkarLoVyOEaa+Ors0+VSQKI7Fxz/46m/s2gHiVAmCESiIkgKgeURKXO6+qT3J
45feyBcnvF6AkNA3MZFykY9gXxo2BSUaQ5Ky8Kbb5PD8y6nnJx6bSV5W8M3Rnr8W
7bfTsihi6p/exVYtwQvvU3lYV45gzuOHtEheazslHtvoOvxoYbVa2Nt0CkBFWLNr
1rcLEV0o7T+7MucyJqGPvd28V++EIVqeuA6AbrUkQSpwHmVDmmXqORPAbwtMmszI
lIL/GKVt52ubS6VURpUQx02QIfYHmlw5S1nSwg9AmOhPLLEw+pcLwxCL1WOxA1bH
0CpbYPCUbZZFAMJlvU0o/LOaRatw+wj5ercJ0XiYVhp/C5gwurs+lSRKWDWaKFak
+1Yvf1W9T6xlWArHiAcQoqmyh9jW/6foSuwnlfaaayJ6UZkUS3jNchxmg9Hyv3CI
AfXA9DFWddSSuOZI6uiHnMSoQC9EehW9OdR73nJfzsa2I9czL3xvqLDKaTiDeSHR
SMOrSmeHlVO6sNATGt5BdZLgqn8zdFSluHe9dJvEMcloo+QzPvjxueZR3im+UzfA
f1jqSTr2aLov3n3lhi2IuoUFth+daqk4pw8hBLWlajXAZYzv6ROP3efDhYEsacPy
mNtdYwNiFXceUaDOmmlsIb58Xu0e2NHFm9n6F53SGzjFnuorg7MfbK/LsXk1A2Gr
5wmIOj0nxJrGrlPUrVqC+M9PTVMbL2+Nt/RGj+TQOUsJa68mvkH08fP2SrH+s/9s
1DZQlOlLBj0/l+NAiVBH2RISWgvwaOZEgTpMPFG8DrH1eRB8orIeJBOkCr28uGui
J3uMv3+EFR4wvjHKAJlqmj/EZULVO4uj4o3fp+d078QiZozo4WNvlzlobUWPTwnK
1P5GpYcts83lGt7AcVWMTAd/amdcaI/dxhvyYKxxiXrFt4+fA1pJ24UlsF+KkZSR
I4npJCNcG/uxav0nTiyiqssynQgOxkrpwTCx879Z21b8UX+tP/tdX/fikd33AV3h
krYmPnnkFBRuW4si+sGPnpK02gNzGhoaH1hApArB4CyIcVIeBxvCezWlF2m2vOXi
CEGJ+0yaj3C7w5vSmyPy0wD5H2WVEMIimNijoCrr3valOjButu1WceNRRF6VPWHU
q8cnArVLYckOKAQxDiyfpw6INM8odIAeAmLzTEkZ/xt8kuC7BRm8hdK4LUFbIcJY
5vcXpEDQkOJ80Mw3MXAt3GQ252VSM11uxMt+MvbT/uUeWhkpy+ApGOf3NS3hUM10
mA3gijYAVvhUlVKpnrkGtYKSZ/DnEr3oAgmdQVYDj+gA735RhPm8emDdyFDrYmjt
xdGiq3h+TIAod9DID+bbDgVHi8nKjIpZqD8N7AFzbaV7yj/CQEurH1oIW74z6QrO
jNJz0g+P8QdJze9+bYJxqV43qr2lpgVu0dj1jKFYfcIlvhGYwNKiaEj2u/4Puf6f
UA5XooGlbtezdjLQKaT7T9k8tzqTk6nxLPhqMPN0KqrA/0xSb2OSazRT4PycrcGV
gnh0mwhw+1DDBYeyuUGWiSeVP75eCyeNss1QZZk5LerY6TTZQD4wdH9GfK1+z3T0
h+waHCUzTAvojnFjOnN6aYDkYdCjba+VHDM1Qa2D193uVXvjSN6yW1Auwya/HJ5s
IQ3lspoYwvOgaf8CF+Q8HXoCeiojSiS9W02y+4LzoBar87HRIbxBJPNc59ezP6OJ
2gJfPi/lr8jB7+WqMJbIuM1pUdx7Ac/EBNX+Y1CEoKAfh39OifqCLBDoxO+amt4O
kJYU0PNoKIGr4ywQ+kwmC0hPyKrZeHtmKzo6zZK+E2G+08RPZN4giR4y5KNAUzVE
B45C1xOZfILXhwKQ7YB7Q/RqBlG3VQClwOYFmOmCb+ll5UkJdKkl0E8RFMxW2i9C
h5HR+eTolJCqYF1XNX4s+FEWwUxPNQUop87aVhzb68dhe5dIygRaqxLCJyg5iDgl
sxAlRh3IbBMTb6Szx5QGAjjKs72TJqNy+W1ZbLjITtBk6cn96Rc9y/eqrRen5OLw
bXRHE6A9uj7c0lvvlJqVeH6bc+ERQP38c+5qfFnnoxxyiYW0/vt/3OHPgt0UdOU9
fpcQDycLWKbVB8+4Tq0ASrc+klwM4Sgc6Ia+tRg17JXTlynRqOvpiDBYACyxNqBT
VowDN1/k9NAe5liz8h9mm5h0kpGheWX2+UCFpx0aI3bVlc2ooff0H1MRlkqn+KPF
QIur3h57F7zSi49dLMIo/ZE56KTzgXnnxxSaaPgOB/o27EV9enTv//ZpebwEUnp3
gr+TrbwfBGaNNIMgyGzksMc6OWu6oUVap3p98hR/FyWXeKTlbJpuI2jiJ9oxSLdT
RqojKlJqv8GjYHPxEPXncDjG+vHeCuD7ejF7QJ9AOjWswcToVsAJWsIXvtbjGsu/
wyHbwhJi3oc5Qif/aJkXX/DCXvs4U/CfF7U6VQe2b1LSTMuaI/fs1MWJl1qXvFvo
xLwiTVhVANl3Xo1CCIzblF+9l9YyF+uUJMFFE33pJsB+qhFvsp5Lgf/X86NeP/+R
Ve153fWD07DKwU5iG7kSNHwAw7rFvz/wuInyuWxkb+6JJjYTqyDwk3Oxei6BQO2+
UK2ft8jIGmFR6XlW2EguGomy0VmO82Hh5QgMvS85jmPcTbOD02aBxoIkMSQ1Hqyg
74JjgM0NzoWx5HxFUz0jo14ttyBuLWU0D4EOAU64maCr8y7LOJrR/dsBJDm9//sO
lTI2W08dkROPhubpjp6GU9Sn13teiaQVV1ECV4r4YyfLWjoOY88ul/ivnQtOKxDf
Bp+3bec0VTr/yk5us9SLQMoM+mNWbkgppbPDCAmTsn+iDiG9XsxWh8ee9tOa8Qaa
dAvWm+6hMAMjp2KsH99aOJZLAyw2c2G6XBJsF2OId7LaNleRxQEZOb5Hj/kQD7sD
MYhMcpXVgiUz/NakBN3tc075cdcSBqSA/bH8CNCvLBG2pmgCdW46AqUPw7iZRgye
DpDKAxNrqjAqFc2O4ViaLKAINNQ0oOZ9amBJ9wS1HkkfTOAlXwtfucqPHT8IcLjW
eAZassBNjmWwhcrODHjKlmFKT+YMuMLlYq2UYiYrdCyFUWuPKzQIJchZNbCCMVuo
DCxHnEqwW+Cj040Y8cc2qagvtUg1hCBaYNxzLtmuoH03Mq3dDKYCzF0UNEmK5GgK
KxrMCp972BRUe4zIdNFs0WtNOMbpwP2k4u1K5vRUKrnYNfCJ17UGup4A9Eur0w4x
VKPLETl5nl6VkroTXZ2H1QbRmD6jEnnmL/qAqfnfuXoNKiAzmbTlDRzvKxuOFXVi
FqgMW1f4Q25Ge+n27Q8p3QRJEwTZaHgpInyU1CjWP5YzcgWFsaDkrvO6PNMf43le
DoFnfL3MdPLH8Ls8kN2z9cJU17mVAijAz5TjTPURG0s4KDxWeKzxh3xUN7WKbWp5
2mV7akiqCKl2XY9qcaat/gOak0rSHY487EWmO8uexkKwIXcMfhGSTEaa0IQdY6/P
oQ20yd68k/zGLA/besuUflUa9I3E4CfuDNl51ZeloNdCZO+9t4D3x8s72r4Gw3My
S+hm4vpQBvFfST2LZGHYpydYZXvdRjA5TUS/NvtAkyZBt6a5A9UJYBIyxZEm5k48
Mv2ZeUWaHOfijg/ZYB+1J3Heno7+VwjJmPkH94Lm94+bMrZ5qivYrRD7Q4kUALYR
yVM5g8TV1mTqFQLyWcAqPP2KTbWDZ+4uZo3+R2xEB3HG+vqplpMes8ascO7QXzLJ
YlWRU8VeUsrw4g86ngsmjFX+SappTGICYfY3OR6DxwLjpG5eyqmgOJhhaxXhFAuE
pETHOjldqweVNzsv6Z/AxwgQH3PfmPxUP0xIINGtfMCpD3oRqO7kMLi75gMdkWiS
0n6D/+fDJbPb7+s3gAlsCahi9sbk8uT0zLk9SsbB4czx4l8GqG08bQXUM73lEMsL
5SA7h3J/rmSpZPbidSLi5UDOCmkW86/BojaM29VyPiAQ5glIDAIX2LdkGr6yw5SJ
wW4lyqBpxFh6EYpmQHKIrx17eRGSpbohQEB+uqpJVFSyU72IzW5lGY/jHYn/U83J
U+bi4DY7oPF2g7MG4WFuFuTUq2pl/Aa9XhHW276mdn13LVIDSurFwguD13ujlke/
4PIDBtU6lS4AN8Y6xwJxR8MFZSzElnSu1lIbwNhwxXNUna2fZsHMGLkj1hNxIbVd
HMdq39VbgloCexbQ+/N+7zsE2aIACDJ6olYXsqSJZWa5D3AmWWYQlJJNPMVHWKyg
rqMKGyyAe7ta2dBGADg5i2rRrePmu2uyg0Q3YkqP3lsW2FD4cEosT32HZ1jujA+J
01IZzIfMi6h1we+es2lPOchUYGSyMJanPPjU0dUXwaM/aONlhlZMQMP8ZvOOGJFJ
zjO4Pt1MmH7IJSL/SGwFhoTyFLu0FCnL2uh3JCbFoARFgAuEnTtJDED6RPXxhpJi
qk/mWY03KeHzhUUmn74HBegQ4mFz4PppALziq779xJsDNIfMomxZzb6qJ4gM54Sy
QOUwMYuR6rcVEU5oyr05ro5iXxQWbjaDzsKNjqJD0cz/M+fzvvJek3sPXN+ufHj8
Px8e1ZkZyghon4HZTXWS9fTEwJZFJA6xqihK6fJP3aRGJMvPXxSNWAHg6btlUPTl
3M0rGhsOF8lI7xr0pDOZFzrW+Z9PdwalVnxr/BIUanylvnREOXexC+DZpbqMeTm4
FaH6KZZTLpUMyShvynlQR3wEcY2SUVC0TSf/xrwPqSrHMAfrrWLQkazABloKBIR4
Hf8urb45Ofjw1lcxcRHNI9JWhjnmx3Jd9HFkfefCMROgZpANi6lVPlo389dacHLc
32/fVyNBAt3UgUQWHUcgBy/3t8c0B8cqk/o3zvA4ANcBJgK+IkSG1V6R2SYERUUD
gQ8oSbbezO6j6Bn+ROGloZ7uvlpVKnf4TfUlrkOi4D2HDXBSw27Iflb+hh+Q/tE+
+ECpwhb5Tt7+aHqDs/t9lcXscQaIK/hGDbRcd1eirYbjTfwKJBu7xdpqi1mc3gnW
Zbbk++v2nHLTOma04ueds5yZxvhy7azjQ05sIuv8uWOYdJ3atzieh8LVTKYHLlVd
aw8EgirkqC4NnpxSXfG2UkioJRtQYNIz9yzLqi5fktgs5qT18+4peifCdgKeanqQ
HTM7gVB+Cfq1mpgSB5Smn5mZ5skUrr4fWk2bwbWCU6bVJdhKb8bh6mO2prjHWvuJ
TlbH7aIlS/5yIldVrNcBT9DTxD5kRukmdqU6Tg6HDGU4pO3QW4SGtSRfK+IpOdl8
Qj8JoIzPSt9ItKn3wwtqJ45nl4wVGuSh3/3PsI3uXl9C7W0rnWX7Nm9IdEIuSKLL
AgT5bbnjVkfYjNWFCFmZX5yJ3u/qiR0P2ic2HKf6hctXr5Ueb5/8Uun0psDT4/1E
xoWdMm26x6GRu4K/4SCHsNMDPR6IxfrIx+wvIEEYpBrNeWyFm8QNAtogVW6qnF4U
dnTRW5mnyAy1Ytf5Y94RDLPtorWBcsPsngL/bzHyX2sRlP4x+skkABo5LpL/8jwK
+GsLeLBWxCl9Yas9eo/QE7peQfXzR4lzdd6bazSgvaoheTq4qEYC/xmxZHA87KE1
8V+/+4z8Evuw/15aKnOdcSVLvNhQUtXOBDXlgURYDRLJwzWDF1AdchfFcQWboNMT
NWrvYVjhbd9FAiVWwYeEluTHBec79gVpPtqEdi7UtQKJfZKGK49D0S3NrxOwPDlq
WL/wNgILE+/Mxf/YsOo7YJ18dQyXGKMmLeJjQkoBVq0FCq+MM8IFFzo4VE6wYafI
2xKYI3E8f4XD6bmopRwh9WVmq6zl0aD+YP+K9Qt2PmwIIdRLWQe+/CWSzjyHx3CR
`protect END_PROTECTED
