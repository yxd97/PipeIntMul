`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MXsOkp3AEL8bSlUo8B+SEFYY2L5tE5tehotNyS1jVHXWSp7K8c4YUXz4bS4duF8I
KXOLkCPOpUww2BOUe/B08a7RerBgcs+270YCfmZRfu9gg19Id+GTdFXz3S1yrGfF
/C2UiXsoY6nN/czeev1i0MhHO+ugXRj4AzPddNVYQEqNtmfgDdIXT7iLDHpx0x6o
wln4O4cBIYPRTuFxsF15kAFTm51FJObw3jBOW73tL2bbZ9izcP04+T+dyob3WbD8
gJi872hGzDTci4/oDuT+KUdehm/TTnGoSgyqs2QIMTElFRGwwoVtpg2y9D0xqNUy
5+Qa6T4qrmNfdqZlHPyzI33XUa5I2kdwJHqOoH5wzttmnOtD7EZu7lgi3nAOqxZB
cvsGgAo678D+TWyarzrYSsRwpb7v8v/km5X4E6a3Y4TpjP8ZFmMHcpX9MQqv9DUG
13vLrAYF6RDzNDQpgzVHpvXKBfJGOiq6/P3XEskhGIOrcBKbHqYH26w36XNym/gh
uXIWE9Ka+pr993A/823GH1kPmzqMIrgqr8aqLgd0dy0BXfoxcR+ZCytXs4zwyH4t
aTe6GsUcpUvkdQ1Kn6xV6QFGGJkl55UPrrYx/X2ClZ/rMurN7U560xM09+SauS6w
qDtW2VyYNH0AajKQWEsYb33tYnHfSjlyYpYSPNSNimdE35JuH8YD4VxOMeiooQVH
nztH9CqgatJpGQGEYgxr2ni31QA7F26V8vc/EBIIbxNteNduBJmuwbxuXBSh5djd
GSg2cNp00B1oFA6jaKC8bJj89Dgtmc70j6G2hPEbP5M=
`protect END_PROTECTED
