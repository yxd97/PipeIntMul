`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ULNz28HZB4bB+klrlGl9yV82fhA5U60zazY6fPYaDoz2tH0O0I1jyn+CecQvHiWW
KPXAUqJXfx3y0NgOVOjrDmjF/DdV+9R8Pq+3E8ztbgAhJXzkbg7r/+190V7UXrDz
sLthEjUoKPVXNtPgn3+G9fbcYsYRa4jP2VmdDuidI0HhvZZY6SpSKzxoPTxrSjjN
wUSqjxGtbgYkZsp7hoR0bZuqC64NLWhiLJ2UbUNKzJv2DwNsHQB1VYvEPn+Htsez
26aOADNE7TitdVSmW0VvnVkO+B4/UibVqI8kgzTcb27XmYmG4OTL8E6lSJ5IYt3d
d8cVFvRa2Q/bV3YV3vblwlnDWy8wzy5OZhF1WMQRKXPGXxS2NFj4FwbR0lX/mbH8
n4zI9F148XTEokjYOHH7ht4VriQgVJtdC0q7b86jUm+UBLk7XL8nyO2K8DWoAER6
sGuLMTt20BvVXf/YgQtauxBrCcHWNxvJ2ja2md3nN0CR+31/2QbFHs1RxL7UjYw6
/ZR4iF/mOUTsk/HCynwEFfMVZxnEcSoDTWIHj/jQUby4VSmW/mYoF7JSdFlzemxd
l43XgIRKp3L/f0WIJjJ7y2IsR0HuKQLfCL+8PvE8JqYheK8vFByMccVGdzsdKqD6
g+STVoL3G4ngClq0KoPK50KoflpKXV4qrnKqZSCwrMoUMDrbmr8xW8dCTH754BWu
rq2+tIdiiYdGLqgdpFkRPmYvQldgM+2AbIeFj7PCpfDIP+KxiJDDwJIeH//wAEpq
HKa8VSVsWIOWlCouCdTUI+ACdlkYoofl1cnarvOz7KVAX0iZfalqM5wHBlNn7frr
3Vuhs0ndGYnZuzP1Un+Nl8cifx0JCmb6kmXEhOVYeOE=
`protect END_PROTECTED
