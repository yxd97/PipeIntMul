`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zmrcjw/zl8a0hYz/ujVgVRxOHcrLwnAHVqNGBvaOGmq+Ip8N+li9zz5CTty32AVR
t3VW8x3infhNIVo0+/DOh5mFG7tC8Xg3C7gZKnIFjPvIgFGETTIMwZsBP6X7PKmU
fuxtXjt3wluoGMl0mlzCParzQoExIRsg9ttBfiWfj0ffceWaMvxL8JXrCkBYa07S
InlVxcV2j05UegXsPgpPkKF6hbtFg6f9AybMUX2gjXacIDk3LJvLKsuyWueTxWUh
5aJyCxxZ59Xk7o9fJRgJbyJHFSB3KFI60+KVoBtzkW1KA4USy9QBajGNLRgAKsEn
8f0svZ98Tn0dQGcII/v00yJykfBVIAKr7cf+A48BiAqBw6NIDa5N4X06vXoz37y6
4mq1vjZIyCAF5k5ffwRG1Dy4+q5A9MLDmacTUSupJF8K4IU8EJ3yICOQoafFYmma
6Gwczzs0aB5A286Wlo8YH9lY9v1IFwg9ros2agJaVGe//FiCymAIKBIB6Ejx/ZYX
lcBcrXCml5owOcQQsNkWgoQlKUAYGO17LtiAEEusfzOuX71NgEX6y1/p0DehZBSE
NNSgi9oE8fgT2+zT5ZuqGjmjpg5+G7rdDvdyqmacHvDGVK8iwsflt+hUJWQ39n6S
iaJo576HHUBV2RHnjgIP1bGvOlKdd2QbuVzPzcwupkuvLtc9mQzpzXqefZqzUk4X
4cvKUssRPx2DACeSRzzM+Do6pZK5P7YhFW+ag34lpDHuhPXCtcFjcskPM2Sm9sVA
U1afyNA5R6tTZwT1onoNsWtDkW6BHQDk6VKjDm2AUZmZ97XTlFE5HGUktYwVtyPF
0E2nAkEXHruGtiilFDRjo3cKOBSifI7hV8TBSf58bzV9dVrFZRXkyVKE8QFmTRRR
OCmUG6JMybD0rS6Hk44vzGooUG2Pzd5fbbJzUZM49bXf1/gLlFJBXJBn/4dVblvP
Q6kkCUKDNbWRPLiBuXscOVNuZmwAnG+W1uCBl9TxSaZJgDRh6gFUIfsN+b0iy7Av
H1tRv++GpyUa5YlcwWuSP0/zwlGLHVfCX3+Dx5d0l8VKCwKnAkcvS77187kdQuZq
Sv8qSGk2Xx5gi9EIBbOzfYwhEucIf4JMNdt7OROmCBw=
`protect END_PROTECTED
