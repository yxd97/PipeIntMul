`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkzVf3905EE7b2btH7KWcx3GXYUPzXTeQ2ltr4hmY7Pjk+/BTiHxT3Viy7qhMGJX
r4Ow6DrBicqFHBzVmL+Qjgtv8bccpGK7GFIIP/py+pDU+e5/LJf8V7WeT6Wc/zFu
PhycalmRijHlzBkKAIrfzfqkE0R8DmzDdcZZ3+61WSHKQCbt2QOwwYdymjHGGivV
Eai0RR2VHlW0PW8nH7j0IBC44IQ8Q5nMlzNcBASIVhdl33atCTTfMlFmlf6qzozt
ScWv6tgF3R45PGCel8Na5IvlR9g8F+lTH3ZMIQ6MxCnxcrcPPCJz7R/4UxOjrmcY
hi/8XDiog6uw6sNInVTGm5aPymU7kmo6lB4fIbQb9zgKqA2BSY6+0LDsxm0W9vjJ
oEMboRjh4ZnkNAOXk03Nh33FK7HO2RX+PZcuuV0aL/NeKqpFf136qoGNRvrWbIh4
PtK9oD5xbcbRkZrCbyiLT1pUgNIbM5u8m2ziw1b//WBtaX6vlxVbxfG0ZROFGSPj
spl4QMrC5Hkq5Zfo3RvUvzYwAfjqbMj24BeXzDvLnKSeukssViJlawDBPNbKfROm
dtiPxb4niIpg3xrE6MAcThH196qfu8qJARuilkOG4H2Xl54kDkskl2z7e9Q42KyS
spgDno0Lbpu/3GUg0kqTxVrrmOxiO3jvNZI+MlwjwGp/9dNgBXnN02x/21z7uO/s
eSjjqNOYKwQubiCeVsHV5E9tleprYkZxvTZLKpu+DInR4MmVWSc+9KEla0uT0ceS
epbvDgAywMNiSoYvb+Lm9G/hIYcm6+JWoFinRqGWvkWCLYEkdkW1Ro7wZgUKp+G/
7C/nwJHO/GcTkyh8dEjmF1htzVmYT5YVkjaHTXzCianhnyJ6EBv9p0YpxIjHfQvj
aLXtD/clY3+77i+XRgEsLEJIrgeJSLm6WOEcGBbBiRqetYSJr2pDZTZRa3nRtrBR
YULAO8OGVL81xtej3d+hi2FbRxhXURterxjlWmm0zBQ7hrwUje0ayRm30OpJOEFf
Bx/drZgrine++a4tzBNTrg==
`protect END_PROTECTED
