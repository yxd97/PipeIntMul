`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
keJKCt1YVOMtZSfqTjaCoZoD5XWsdQuDYUjGIcVDTpJsF8Hi21xH5rTMfsWPEFuf
jkr3nkjs85tWDy/tPnWPCd20TM+oa6Rw5S01YmNWX7VCnl6MAFs/SnBKEtdhOFC7
KwqM+h3v3qKbqnaMKi+VZPcZiWQYOw39bL7n8p2mTA88Flge6+WA1mQTkcEhExjU
mOQVeQ2gRUl6Vrj3nVEXzp/iGZ+Hia7eA1T03aPCii0h5NYq6v8QVrEkHe4HjVwL
mdRFHvHpUwpy29VmpJZlxg/ehgVuyFRTWBmFRpS/7wgIEWdsTKcFNXaFxNLn7+3s
wE4AGobPne2zv619/P/dEBosRP7o7mkvdO0waUqiUg4Zn/offYtGPXjH6rUIWxz3
ZWFXmUUPeyPgOthvjNFpwks4S7KJMWWcUp4jwm/6G12EsXUNTLA4UNhSV2B9n7dR
gtPhfY+cJvJZxjeVLlt5y3Eea3T2WSGTFrQ4Pvm4ZYw/ZXGo4estdB5ZxFSZEvO4
Yq6nsLOs7tOTp3ej+KO3Kti3Z3yhHsczGFUYL4RO5EzRApYh+5NTAyrFnh2q6udp
`protect END_PROTECTED
