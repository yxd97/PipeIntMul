`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BgXX1/gETaf0Fer087lMvn7r1N9P5LVIfgt++7ypxfDu8D5EsRd2c+0Ephbv0a2
wUZanLHyLXaDf0agwfogl/yggwR9K5v+3qnA7IcK6K+JkB/1noFxaHr4Iuy3vqcd
q+Syc2gp6ebUoE0nFbia0A385fOw++9xJslArh3bBxlPIWSmPcEBKhuIIfQREI7g
nKVD9p6HE76nXS8ykS+oJDZVgqGaN5fxC30RZhYxUk0UYgzthZckQ8fahWpqJ9xh
MmjFpmvpU4TLP3IC2XY1UmKSDE29sTtEjtP/t006xKwuzolT5VUWRGPSpy8x7nf8
AUIXJYx93ox3ViO2ZAB9xDseqFJAefo/HSQdmToxHbDOmZzx8PhxZEouxImh5REz
Dj8vqmNjeplyyOEZjIdMHcATIKv7l0PahFhI/vHq2K3hzxqcOBNEtsb046/nbeQv
3d1B3YkxZO6LGaOY/Pjn10Hn87Nhb5pC9zBK46+Ofc8e13/iptk1QrNut02xLyni
drAp7IGSxyabkP2Oz6ogMA6dycLGxBMR22OCC1bNZQYnoId+4PSh7UU7veIvOAK2
6LbF998neFuYvWVdMIPeBZAFub0GzgwwubVaZe1YfngQGmPSJnqSTfN2CN+g3AKF
e5N3XZhGSq5rLI2WIasxmDIwZmK6/56tb06AzkQYIq+9+aMmp9Q72fyuSBYrBA83
Uui6epyIT4Pbzkvp+zK74FNF8TtJFpEzVvq+SjhrTuQnzdLz+/jeLnv1ikQ6QHNM
NPkrPFv3Y1Of04kFwv2z+mCNU/I3Wj7xIUT9A6rByewYfVyQpl+UPCweK0D3IpyX
WDZLpTHDqecJF/IYcoDjo10HhtKuSra/3rKmBoHiwASuiBJ/XpqMP8BvrBt9trCv
fh0GQ/3BPxZAKnqZPjIkJ2SYJMjVyfwKbaW6qRJ9VitQRivpmMQqYS8T3wXjpQYm
ZENto31x+lbT/qVKKBI+agXU9lAfHph9kJm2z0Cc6cu4l1/VhEq/47wZZFEteaZ6
vCbQdO/nHrmm8zgHvnBDhvtHsaoYIH/HwNGnTbOa5zRXjqB9VyKLrLZbTgGzu9NN
eGoqh5Qm+jjbAUe7w/hG0o1BJKolTPY8Cmlz06NGV1XlLIdR3YNS7ytunuiD8+o8
cKdi7tRWApIbzO6sJr3LS16eRT2BRzSIfw5SrSerUE3z32UPyyRDz5zCWcq/klej
D7A51zZwpa2ic2E7IzmaNm3qUZOMQUNhj6iVcXw6VDfqhfxFXXf8ywJVg4gdfzem
Pfk9/fnAlIJ5o6xf53sCWldPaI5lURTTtZlwKwMpMQmNxywrvYKlg8QYr0lMutJZ
zVteE+pQJoFDuF/LZbV73ytgG9XRECQi5sp44ggjapUZ+lzHPA0fMutdvyUsNy+k
BpBRKxV/db6Te4x2LP03ylI/K7fG/+ITWK1mF8S1Tc2SPmxhcgPED8PxonX5RClf
qgxS9jv7ElKxsvb9R7KlSiZuJhSnfFaUsmahPUJP0GPGpnaiMPXMMn34zxJRt1Sa
Ir7t79OcEIy30kRUhpmfzOvXkVtCMY9KOOD+FvvVmd7Y7XC6/B7SaZ+TA2TYsLjr
ZmgamTnKVzNBETWTSr3mpblwzeyTSi7xmz8Jo85fYoZjoM4esFRomI5ZfbgDLh17
paA+QleP2IEumJ6Z8hzRqMRQ80Sb3IT9KqjYIuhnBbs7ZOaFqF5bqtgk09J9esKs
RpfoH5VXPPP5Q/pY9RWodMrOSMlwtwp3TbTkKGgPA9E4Ye6KO7WSm5yR/byVdiX4
Ovze6twXaLvgS4GlCIAwT9BKzO1838/tF/UvmLu6LnfIumiJLI8tqSWr5+kiihSn
n9ys9n1zSrlLRLrr3agw7jx90IDM04WfH6OKRc8RMI7x7akGsx8cmlJnMRHGsQsg
znK6bu1EucQfIYFpBR9UPRKFPtgsF7tnkyzZJrUqdhCbyBekTGTXp5ztGDhgYr7b
WwhfVaXAmt0cQk1NKQkeGmsUg6B7tusmgumNESGIX8JS1oGVgVdhwC3X06+qdOUq
vQrJXc3Ub8PZtnrOyD6D5pDDlw+G+bjtzuCuPR/d5NPB+nCLHETnlm0YBl6+M44t
S8iypwWvR3zSd/8OjtPgl7FZaS2Cry7zQ2LxhhqpBlDz+KESlkAYdWfIXNnS3OgQ
W6GjtV+Qw2+fvnheE5iTmJwMBtUd0m/Jxj3YC6JFqPS+TWwOpYIxis9HmiMUIzXa
iChr1o7HUx0PLYNjKtDkKMIVpqfWkM6inf6ximvQxYWnaSmLl1+Mb0bTc0Xp3fvl
obpzXlezDTdlbEgAtJr58XG+V5CM2JDmCaxVrZ/AZYNoa+MWh8MmN2tuKmRbQESH
ub1TduazYBqkj6MBBrAbLjR7u5tAoZsKKiYxKzHUlPNwd/V3m1Qn12cea+f4lF8+
ExFD8gP6kEDNypMIee+oDhmUtgl+BIpQmfdcLNPOfOpdA4ZhB/ySMZvjRX8Aj+07
jCRbk7HgMxcCl3p6+zk6BK+3zxvUAoJSRWPgnNAhkfqc0NNYi0p7qQFL2alewbUB
evrqft49gRMFgkP8L/EG0ImzQ8wUmCeZ9cIoYhgYZqGvkkBXw78Gtr0Lvnol98e5
bkGcg4ts7yQ/MRRQIRhBabSuaL3Q4TUqWEaEeXRUMADCgPJkvtXIDTk+yFDUySw3
vmJ8bVrDvoWgES9D23G3yRqHAtJr1sgYP1/R9Xy7sAkIjuDarRXUYTBl1/r0uyB1
2SA5cBnVeESmbEvHlBZWiys8cNYQTuGLclh8GY0dawR2fuinr4/FZlznNTDPaT0Q
ysf2XUHMjHW4Nf121p/pD517HIEwHr91t1J06Atm9aS3gmErScju6pTQv6UKf5E7
X8tSS7qKm7J0Uz/Do2SN6lGWr+NnLA0nQvEEq1uWCkEU9OGtmFnl/JQ4/3zwbdEN
/X7gQo4IDq2Zr0U7p0QjMkMd3Iry3096Rh7XO4XOmfxPfrrbcNb+PzSEbixGuX7N
PZWIpPCusnscL2b6lingi87+7zYWnjuDqK2UBpVxrLpiz7A3O3X3h4F8IQFLaAU2
QSs5mPUjPf29gsUdppVHcb88VIKvUDjsMn3snhoYgV6qGMQCN/1tSQeRifZ5S2Pv
snCZ1hLFB8U7Jx3qtm2cBWIkmNOhccPsQ/lKeIsoxG8mfW2JtTfwriC2vQXdMzCV
OtPsAXAhXdxDboPQ8qtD60PMmsHwfQOkMkkiJqzwN/BhTuTtwISnKxhGJ0iJlG+j
p9i/cIvHPuC6BQx/491GTW29A9t9ztOgIWbAFpJMjSXvOLk6IjkiqlbtmmHyv/W0
BYkIW+IKV7GGpZ4ql43aqVgWZoTiJf/o3Kbql3usF7aobGHxQY7JmPqjI0LK36h3
NdZmOStuYhTb5NLOavVT+JPFx88r9Knxl2qZrqPxr2t6LnleXsse+Fz7yT50UEYX
9GoUj+igefuB5HvE0aDQZ12dodLjGszJApERe+KE20C2UNOOqy6Xjlx+InKb73WX
BsVAnw0e8E4kL8anMb46waHmHUfK2JzHFMmDD95TkhRCBTh/RMogRuXCqO8NXJOV
8TzVUXwG2v/P0vSFoIf7NTglMV6UeVm7CaAZqiqHxOowT7IUqGUXsplEP2QNuNxz
9CZzQLa8f9+yXcRklf25kXBBE57Q3GjIgQTc609tkfHTnJTKeuzav+zqWLJIYn0g
G+f1+incq0ksK+KLJsorzWRWkpkzITDJ3PgDcV4b8O3uh2ms0NpSDHoKQqRiY6OI
HZGQo+ilBkSGc67BEgS0P2zGhUJadfZeUq68fpIdsG9OS9y2h5YT40tBKmHD8HOM
k4PBbakLIVjLu1WXWkZQp87pDx78/XWHpgBfpiJGhzCEebaSelTmLNgByIjSfLdI
MqiYK0bm0ssG14f+n5+rKHi9s66RwTqNE+n+dHdeLUpemt6weZRAlEss5dmbuaZG
r1rDeedvI0aT2Nj7UtfQ/Uijiyc0H7vUMoYjXNo9FFpObKVqxEE2H9TEh2hx65W5
wV4SYMQmFKq8yDT8Lk4XPykv/h206lskwRWr1sfGgKn491h+pNk/MRYEK/Rr8a3U
Xr+4mw/MB+heUB4c8uVS7PCO5Panwq89dvctdhXYwEfQQl3KPTkzS1eKj8Yzfz+3
ocKnlY7p4i9isaRKkcU0l6i6bf3OROSUJ/KC2w0JCpgPpP6BXmRKZMOa2mjGSo3/
X2Vzg+HRdQBjllG2C8CuzGlu8wIe5/zrEQq+DvVz52DYxl8HUCGuI+YgAfNHHUHs
A1/jgmjYGWCKnXLJIoOB2mBfZKw8J++KfNWacZ6CWkV20GkEtZ0OB3sWW5NAA1jx
OouPbYWD1yuN3M5IChFK5pvy6o/JJAkHdtEuR/e59tpcy8omIZKeoMg47prNosq9
+AF9tp4mEmMubgnkCYBTdCZjNzehE3mkNthQRtLjq3OGTXCTRVoNQ+CSQ6fuTIzp
6mpCk8zQ3SfCYACgZPbEwdVBpZpidRCreQIQZm+dflxlmADEN6I94D6xfavdP1ul
ZTlT9f0EwlmputWj8FBfC/XAtfDOKGg6fBd4OX7X8EioDG4SwHteGqc0g20OZagr
hRQxEgz57wIWPjMDfyeLpZ56UHo4Ofm/+CY65Hz0j0C8YaI8ISzKTwYMME4Yv0Lt
rDcUOqu9udZkDSlGuFQcpJNUlqvUDxsfyGRxVHQvPY2tue9sFtCC79NFC3e14/ju
ig2V2+1XKohXHCzWYoIxlcyL7Z3nxGD5Yq80SPqmdF2Ll8DbI5zagQVE3itDzxGS
UPQGnxAA5Ycxc7CD/0RsiYV+T/p2m2yZLlEMeWDUedvd3BEdPmek4ePlNYztFA2C
8B3GPhEdUiefdIZCIZHWbf22gSMD8zDyK0WB5tvXmkxvejMC0DgZXrczSDX3vA43
7L5fi/eUca+CWkeUDjmck7MSWke5prG4lBMp5Xkf1i24RaS12kVSxHWJDMSkP1dl
UWwjWS9GuXWzEDBsBX9Ev+YdGBBMee0yob/J7IuPSWWI9pDS5iPUwa11MJmUiWY/
AP3u5Di8atluH1j9Ix3J0vIrF++61io8ZW51ylXM+FZHb8KKbtcziT9o1fGG733w
Y2hd5IAbCGmqW/l5SnPXrQDsm/zBzEtCJnGAdmBEmNWjHii7hcs9x0zAIjknQOZH
9HDsJbLJJMYUpEJ3NaMUrbV6yZ85QKhJWPd3WUQIL7pLI9cjZ6fj8oDhSfXVDSPz
daxqWoL4CvgsIfbBELnEsu5glo0U9xBo9QJKTN0h5m7GCWXLJjmv/P8rbXtZAiIe
29UjNFqXprceSWXjGxvV23gvv1nARdIdi66G2w2gDA+00TgyQOV0KaQFLA21IBqk
35ih5CC19E3JqQCcbjIk+sIFqEEq/EwsTHOhnYl8J75NFRJAcGy28UrUNTJywTYk
9IbXfSZK6x1ualEBtg+PcyaqIDkDSJOPl+ScOSqMQOQY4zrPtFyL89SrkLk9SxBo
yDIfjd19wT7ImEAPy+SOJvCwWXIsL3nKR3KJrIJHECOeznI1XLyWcE63soMZ2LRl
zssKLF938YnqWyTwrdTogfX+BUKNfYqWvdkPoOU8Rqaaxv+66Ko5I9qGjL0rwO0h
O82R80hIclUVcZrUldsa14IZ268Kk0QHZtC006PczEhUXal+6XtLSXScKXSYtl5p
aSvgCBhc38c+DiktXiAYV/CqKZIqNAmQz5U58IZ/1q6p0mpqT2pqooC0TP+7lLFd
/1LmUODk/d7+30f9lsM7eaFMHWyP8BTVIbKgE2yYwRVUZkNzpp9ILRa6A791sojS
cvP7Du9xd9u1Q2paBF5tyXnwY7/lirZDfNGDSfCg4XhuA896s/uVFzCFHik7L3E0
/ILtKK24FFNY4FOVdd58q4/uhe5ntsm3DHqhXg6QomkQTgDePKQV4DtNCV8aIBLa
y7+ajlS10AXiOtBCcs6gDO+QBbhUIgVvc9QF4cLMEJqift9nAMgQHxhBGNxX5qc1
ZRieMfR8Q1IhS9BSiTu+wjhRhA3B1QV3kwBQ/pyqUT2ptz+9yCqd6sk6uCuMuJuF
lD5e1psFOI0lcLlOCnVFPDe33eWyFrrJ/6oj/r6+tR/WM5KVQ+VIOq8EyrNhPjjT
bxAKHAgfN2DhCqpeAQzTjOKyEE2tOc+5+QFm2bczzuaD8/haEjN1/n7cZWqpK2Xj
C9AthSOv5ylVooL3IfQmtFOnR83vLvseT1SHmFgjaTh8VsU4bg0kvMk/FJ97+ad/
VhShNceqs4W00wLbBdGwRldIIC6hlnKhI1opxw7gRFRD8cujeUjm7otAmaFXScu3
thJVX/R5W55qLkzVUGGC44joR/QfeVNvby32wUhEMA9AThvpeIFLJzjRU/93junH
Z9UFSz4/ZqcdvEGFRBMQTwXaMq1ZvbuOWLO57d7IeMTBU29pxhaSm5cuUk2q678b
trqqYqPx49047syAX5APCDTQQH4+qWLd9CJTtsUz+VR0I2xnWNjqw58mhiXwPMg2
b1GnEqJ4PvszgCM+recjecj539dxf1SlTKi2vxnCLIE56etq5am2woRzFUjauELl
OlI3VVuBo4fikizhk1yROXvlBLVC7VRX3+EAdAFXGY6SKrAhBnRPO66cWns9VZo4
VNUPLivL3Xl6vWhWlwhaHxFT/bQR+WGDYzRvkV0CvpH+5xRS2Ixp+XjusGVQ0hVi
m9JGUSP4oUOhwjMiH0bo3PszvDHoPuFezUlLUO3R/uFzQ9WMttV4rM54zA5YydER
zvZIHL7UeT3tG/gtWNUwWmYBt/z8oKODpge0sEpUOkbv9FAnIf0EvfeAP8ivgdSI
6svtTcLXWnE20nWyCyVDLoq9adcRIrMC0kYMTli0LsJExYBS1AIgpPonOLljm2Kf
kYlRch+HBW1bIpXZmUSla03k8BRBHObl+3r/qc/IDxjuX8LhG9KKIvDK2EClSpzg
G0nkJ604Z+yvi2+ci0yUFZM5bLNof2DiE3oDRkrYV01Gn/h8tLmwzM7U/hxZNcJP
0gRhOwQhgOaG+aCCPcevJirNp7KIaAQBiEJnOFrHgzSRQr4k/e2g9buks8tHZo4N
guO9v91pbsn55KD/xKDX1UawidltFetPgZc7h3oRJeeLoAD/22FkL88CRJ2y4XMq
lIj/I/poZZZSOQ0Y2PWNmr5d1fxPjy9slNxhwwIb2Nyd/NJjz1WdTedKAeZYD3w+
a7HNRVvEM43QY9+3gqa2QA==
`protect END_PROTECTED
