`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCjJZOrNTegSw9ZT0G98ziwSso5tLwyIClHfDMUERwiJYR0WvJdAKxi1ZHGsm6+i
DXUp8NentVay/aYIWKEKEIBlZ7Vq9MNDTOO24ImK4yTwUfvtjmpcJEDdN2PEiVKw
ovCmpN1xa04SDlq98dTEOr7daJMNGFBelkFGrR0pjt7kduhJCzG8V6TvR49FQjor
GFEKMahb+cti+jAZ2agb+aFY5XmzTvj1NGeDXM6ZA/VzT+uKlAG8xyxEd+YYq1/h
IF8ZBiiLps5FnQEdDtpRsD68bLz0fftGB/bFQW3STQp6dMhLkj9ITpqAY7IAQzUQ
lAi8MTAZUvr808eTTiD0UqGUXes6Q2kqRfQq2w44mIhv6gCLKhdJJNZck1k/Ah2K
eNHLR4xKeVT2E+fh+MbzbUaj+jlTl2THq7NVXNGKqp2lbz8Qa8berI7u/9z9SCC9
+Zbq4QIp482bHj71D9m/MDtHE0F6PeFXK2x3d43Aaq5nC+1CPL6cajqHOjrqs5/F
nBb2pPj7vVDM9hPBgoDnZjpYWX91JQakwoyQzUsA5324cb/G8ySpb93YnE3Nqk/t
+Y5djiAIreFBlXMqmAVd+x5SSXaMZ4bW7UrumqBUxtxwu6erNuIw9UPn8YCMXOrD
eWgt6c2fB79s2+B+Sj66dw==
`protect END_PROTECTED
