`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ztC4eHHfqu4Nq/sGhygweqi7Us2u7w56jP0yxCj5Irn39u5ify7k8+0Q48/hUa25
IB5BH3OL9AdPLcle76DOpTiaqd7Dtp4r7n0ydzqVvkM9nzgUjsErP5O/GSwS0mi0
CjIhDaxpMmtZvZ7BItdgVDvSHK7qroCRlxiftxhVjsA1QzzxWtucdkt8SlqQ8rcR
EjtST9QmjJn1rYwnt1w1u93YuWJYSJE9mpbGMBM06Uznf/qb1Tl+cX0SYGZhb9+i
R9zbkTg7Fi4RwN89iVGeMij9U41vrE5v0PfoVcU3w56SD7nSKKBaoBlJ/opGaaxH
+a0uPkD/19KjJj4ahng1UmHjuQ/Q8xAb0HVWYvaQUhmVSDg1ONJvRi/a7FLxfmBy
AdXWxOt+80L8tnp8bNvo0EftQfYKpY7kLQub293gxVIW56fbk7Ui0y+/KadDPKIw
Cqe7DK1YN1r8FU1vQv064wh9kCK4+CIazlIF/GmO90wY49jh1hlj67RvLPAuZZSS
`protect END_PROTECTED
