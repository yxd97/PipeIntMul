`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uFvtsTgLO5HISyX6Hc+rP5D6p/WOyMpFWI/7l38tgQbVFcRnW+HNyCaNyR9hqP+x
0gm1DdWuhjnWHzui8lpYVmtsZnx/BPGSd6MVEDII1UdAhW+4sJT9Z4w9vIhN5bqT
z54ZofoykFQp6V7Lr2bqD7NZc5P5BhLw6EKb2PJfxFhgJGI9PzUKrKnYgxbpX1Vc
kK7qrB0Rakuw7dRTuWdIVlmus0mOgR4iFyQguicjpYR/cmwrtXTXyYU5pbl+N1Mq
+s494j03RSdqhf9FP/On6Qk4oWF66Ulmu5ewO48de1e0QNuIbNIV63sqGryVlUQo
uAuhZK1pekKNXjlZxTDq6jw4YXqwXc3Lz5Sp4JnEDxWRFpZWAVwdKISanHnZE12f
WGQ3gJElhajrefFWB1OApoMc4CrS+c42x9sBYg33aWBryXbH6QErbNJfoLzx9HNZ
sg1XS/85OUlVQ+nFaiPp9RiyolwTHOnQofmheUsea7m1LnWoLwzSY+pPqBIZKX9I
oc2mfmtqNjUFvMQIPcyE2p1D21Ma22H32g1nLvmAJ5w6fi+XgevuxB4RwctnlUl1
mdcH4Ha1oRAgvdDvPP2h+igyzavD18pxujCVkgaLOBsimtl7/S1jgW6QD/bgFug/
c7D/AThtsCBVqZW8umk1B5vvX0HnnO8VJ/pHTZcyuE2iVKeMK/L7f4ZdXEswHH0e
DXjKi0/ZDAkX2yaDQScCaC4NuaIgRMCRgKBs1bFGvECufMjSU0u8YgUy0LeKD3Pc
9jU+7N6cFvt2Bds4myWvbB6KWvt4eN+ILvJdwTsi0Vwt4Zc3xbDVvKz7gRdfyc6v
nT8dcxOmSBsChLwJzSIyAExh38oXWKPsAc+hQXO2YAqZGnttX+KD+ILEAHB4AfSX
gBpvzHD1C4uF6TqRPaURm5h7V5zrQSNgv+Ma2Uqgu7fHpGHsaIUFtDeBjfOUyl+S
bl9uv5QgqdteGDzgK2z3L6vVW5JFa+fWmToAOIMzdIYdrT0ZCHkxnEMTY6n3/eTb
J3rbMueFZ1V1vykoPnUp+zi23Ay8QqIdoWz/VyetxmI2ULGo1tQuOPU7GpDhvAL4
nIFq5/zB1y6dZL72Zdce4JAZ7Oaovbo4Hhdy+R/YGGfTW0h2RYal4PeFKtfcPGMW
1x5GcDBTwi0xs4r9Ddr8awhY1Gjiz3JdintA9PZb2/gYnl1uw+ImToTS8JvNls7o
OaKUVuUv5UlrSi1qKQZX0V2tSFz3AE8JhF7cGtpqAWRqGPtnXpT/REGcqzVwyHfE
js/Fv4VyUvvDon52bDAoEPsHjwQv660bKfQfOR81R96ySiFh3oVNb7LF3RZg2upa
+N5PInTJPYrwPDonmvALLw==
`protect END_PROTECTED
