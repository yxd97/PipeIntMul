`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6o+XbngWBbP7neEkBKkYdQp5A1kAyoQbp7R0ZIkSA0fZjibXlp5R3asIV1MvFNOO
y2FFzFxeBPMM9qtm94dH7OxQDlhPAGc6Re3eA/1FjPE95/fDmb8bXfZG75KI2j66
arGnMPO8nU57x2RfmRcM2leUMapuy4u+rdj/CZmP5Lmie3LUV5kpUIx6l3kyq6SN
ortkmXR5rPweqhVZ2v8cwFZwIPkfo67Q5rZ1crPCfXk12y9wU8fVFU4i19Z9tRSX
sA63tYCXu4wPdhp5uEvtFgklbGUe/qWz+fKXtZ4NXxiN7gTJySKHon7H4UINKbEn
3UcYz0m1p9pE5iiX7LqTNDamn0AtjUFxfuy+fbDkBhpECsyqOdtvUODWEzj7Im8C
81qhnmyPY3V0aMUpBlDrn61UJiaQGvXJyiiy7vUU/GIvb1MSvZcrO+tH8zi8nU09
P6MgyNjMbs0YscO+KErGhcXyY0a/g3lSo70Wlg85wKe3QS3aCQjvD7Xh0+tbthSh
NbgwXuntIYPPflF6HMwEL6kmhXMzjYWGaA3+h6xGoYZuadutzbjh9G8N2K1gMAHR
rdCxifkl/mdzfNUXk6WCTzOzaMAnh5bH6f6lgcGtmObBL3CWNqOoYwigFFoIaDq3
dW6yDrXQ8OarnN1bNQAtmyNBOThinCMPjnhyVCjnVQsPGInuMKsQMXS8zwAYT/aN
mMDy0AH6ICJ2l0ORN8d9GPqQGAUxiKHlMwnbH5In66W/Ggjkw3clxcH4sEqgsKa5
RbLpN+5UDDs/C8JiMIJJtw0h8xw/dWGtPb+cprWiUuLA0UMJt5T8JQqbpa4G6c9W
FFlxHCW4eXw1wpNyh7D2XHlzMg7+67EFu1zh47wc5X0VZ13L79UBJvlXNbq+zFik
3cVtm2H7YRlNt3YFQLk8XAQUzG3DNyBYmOHxDc0/WM+koIlyZd5cZYjYhGv0nxhu
nF3J7wrxO76cQw7GcCbiz+NPObjyryTEiCTTblZF8fuJPEMRKla8npxwH2Gw6K0D
ORd2NEDOPf5m7mN+mpGogdRXQKS+Y/rO8SOb5zuIOoB+ok8TBZE9Aybd42FYlUb5
76Wy3QGLIPNNrnejtSG+MXc/RqNj+lxlJM8sbKmEy0bLD430B5uhu7x65+uy6QQ1
bhX1Ezayn7YWNCAylR//si2FhzdBzTAE6TL8KweIMmamA8wVQhZllu4YYCBrsYLu
o7K2sYR7grZSNpabKdWZje4jAhD7RWn7OF38bxjwuQlSzNphG2rVcuvXG44RhuLx
DwEixX7Ikp9ovb2jYxLpiQTSPIRFAhw/PvjloPYSu5KU45haTjMOWsoKxyfv+wSv
1Vhsj+1gvARaPti6uky6pXsv1/3IAF3w6Hz4bRNPVrUwPZ6jmhKfkNBFrYfgtAq1
wtTBHZh3bNOUgJqisHPMxnkjb9Bzb8fzEUKZB/iV5hr1aapien3zzjWZn93eDSlW
ON40O2MBPomml/RPd9pXYRxYVYyjnvcm2WBNEtac7SKf5f0GOwfsOxZe7t7LFCUO
eWy5PPGuH9TBcmLWalgoAw8TVcCN4rOH34BSP0OmEI9g/MGaVoqOPB29aiScIUWM
vsyojHPpzacgmjItxj67TVIuoJtDbcCr3PXR2CNOF0M0fEQ+89JXJ+0GdnC5wKAp
oVIT7vcWaskFkTkQig8ILj/ITVf0RUXpnVO4/4wUxWp5inCjRqiFWu4ibwt7Y6pv
y3gxRNbBcfz+4aTKTr4jp76yj7At/DzU75Zinohv1L2QpDkF8lmc1kjnoDDspzED
cl2WROSnBHVze4rvSJRdI+zaD+PJ8kLR59VP2eCiaajIk6Idi11p8SwEYFMNfIgz
EN8vlnOvCJWl07iVBh5Qf2eNdAm7Gbe125vbtuQSOOcJrr/+ik+SoAjwcQOimbQe
+ePF4nVofoQxUOgbE0qbHKYN85d5V8ACP76kcfaEmPzNwvrjuQnYAzfzDOl7yjoV
rMCmyrvn19wjWbp47mb4Zw==
`protect END_PROTECTED
