`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcNBIv2dLHKgK+sed8vqWhMCCazXh2eJbPJkngORbGDk9+VKyR7eO6xxB7WDdbSY
i4qaxP7u9IEZNxzI+NpdIgUzYiHtX7jrDWN0BujxChBuzh+XIOhJ4QBpUOmd7gl/
MQl647DGclYygWmH64xAlPV2zKpkx495c+7gCcPQ68dRInSH/qOWMNG98o4g8Kmx
yS2yPjJtPI+dPG60+ULTCf25eHuaX6TbV1NDXJidSx83Kjt8THfGvjPcJYlF/kl0
tpBmZ05mhXaaFLpZ4jQJPwwq2OtmhsWiVJR4CsmgQFnyxaOU+fB1MQ37H3TldD8h
xUWZ0B+FLboN6fbd4t3gQSxInCdgov+VKME7NrAquG4=
`protect END_PROTECTED
