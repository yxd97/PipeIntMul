`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61HlysydwtSjxduZVSvW4TIXYv3KKyD/LPODWdmz79bdagahma3AZPRtqnmDp2hq
GaSQMubyNkD1EmnLpPj0vhkYs/LqdyGKHqFwzveDnMt16c89KQQjiQ/vFycg4Zzd
mMpRgXWo1GvXXEc19FX1H9YCP86t/IVFP2kkDHduc8RJyin1NBM6jye07b+BQ92I
meiPyZY0Gg6rwfByqqH6qgDvUlKaceJeIC211hSQ6Rs6atxQPDhsuAQdoWXIl/q2
o7TGOc/P9D6wI+4CuuPfGRKgP6lP7lexLsSu/q5YT34m/Uets4d4rEYp7T5WiOQQ
0el36W4nlmIeAPkRToisX0/pw5lj9U8JHXdN5G96SnE=
`protect END_PROTECTED
