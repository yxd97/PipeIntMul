`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eXiVe0cpTz4MQ0rWcD3HE9UZntZ5plVWBC7M5vp8ypKZwtgGHZ63G2MQ9mYyOA/c
h9lebzEgLJgwi+GlzI2YV3W1EKK3Ph6er2tNzg6uxwqMskdahxlKHiwyNcEIbuWd
i/Yk7iHzsf5vtBEGoDObClh33Z9po6qqbQptId0hKwlp0CHfCe4cyJGpjfnyvbtr
lbVUS+6GeoS7EWQGaIMQGJJF7znJPgM6t/LYArgwqGvncsuH/8AHOTWCUaB+VQt6
H3yBNHelkF4OWbhwah+dv3VZFXOl0TBLYqSE194do5b5LJiVR7yK4seDlv1QsDLJ
k0bWlsgLui8HXgXMyCXMPTsApGYH6GrL0EfzGY86H94qQTW1K0gwctQYk4Y2H2N6
4JuRwqUhUDWu/BFv6j0qr6wi12tIFOUHnW7/07NUzJXB0BAQNRBGVK6qA8xDb1E1
qv/Y2A3PvxB+KtJXwavwfjowgcPFxvZeQd0uc6+D9BYcfnRf16kOQgIgI5C0L7Cj
lTp7HhuNDgp4tRt+kCMVLAI7RA3ecsW9/lmkpDG1YrYgD9TbOLk1W0fJaR/wa/gG
vTkROdcNPGQT6YHEUqvrF0+BFc2Iw9WttzaOXTppJ4MCv8xhL2l9g9TXWtvEn/ZJ
8MkjIPE8cVaK90aCVuf2ho/95MYssFO9CwJNAckyObiwZnwByo8/79tS0Fn/om7m
A/+bFUq00VIrWHHUoEyn95v2FYFHEqK63kaCbr+3CaDpSKa5+ahdDtCab9s1Zy1Q
65UqVXQ9O0MPwNkJlhgk5d8kx/CfYTqktPyTI9kA3XP749h+yhyc1PBfCMMzAVOj
2loQXqt5OEoYMfq/22Pg8ScK2PvSVGPDMDjG3dKiZZI4FPoxc+g+K2sLDYLKoCpd
gpQ2ZbcC46dtfGhvn9RzPTCUCzfUELnLiH9Sg7WOJbkwjoK3jtbjDRhHzMu2QJfL
ShX9FFLKgHa4pxeWFQUlKx05oJsKVruX71rGp62u4C77IhC/3T6cSV28Nur3XVP4
uPUCA6ggkge3pTVE71/7Np7s44rEV35awlVugBh5PQe180hLE8Nk1Og/EJ1UHPG9
6z6YA9znEMluU99zW94oYbObrNQENVjy8RhFS8F6SRx4qH55FEcMJBWl4n2poUhl
//2Gl+hqtyXyVE1MFjAP8aYAB9rpjE0CICF/crJIA/X5aKLzHn2n+ijen9uVHvQD
Qddny2zcc7K6V8PPI6wnPkyFR6fLgCkeOh3Ad/lVUuu7v3S+J6FFnYj9d/JqjV+K
9HrHdiKxMRNnbvhVqwghZX5wsEGv424yJ+mcFj32qYzTXQtDNCFdEJZ+m6yho+uo
OHCl50YR51t5oHZ0DZj4gqu9ql/0F2wGzCAoE1tTj71xTRtIG94GvfbmGUBk0VeL
reZzhhqFlqV1TEOPq24fIbTaRwfxDnESjXAvuqx4CMp2ex9cfP//qb9h5N/LcUjl
8wwOSlHSBpAYh6UQ0CnwxisHebcav8nSy/ISuw/ktt1wtTdCuBaJmsu2+yErIXHa
Zz4z5wtg1U48Aj7eDoK0Tegdn4IknmKFeEjSWu4flD5kFOmEC7u1gGZTfWbPRCNX
d5ipm2a0gZyRD4FTYmlJmYaNg+k9OmD0SU6LMu9/s4x+Xeg3sneUPuroadDW/03Q
h8hrexKR+TUY+hiM210RJbeOKwAOKJbNg8l8RH9bZCzQBP6EO/gwWRd3ce4mIdoG
bFjuBPvgEB1q8D0S93PDjeGuVtAAGUqAHhQcOHg8fE7odgHpA+339FFa0Bdzc2KF
I/GmP1o+OKM1XC+roErQDW9R17be1M6pg2Kq4b0C4ifXgHOoiq9hdJ5i11g1qUjp
zJkBLVANm0ahwN7OgVd2saLcnCisK5Bhw5BZWCDheZ3mtUxQOa4XUPPZpN7tCjUo
MVbdzSMdqd1+oAXwoQChPEe0PTDd54EL0zjfPP8LnAxNP3kQWFrTrUUJaXupLfAI
iCLf/frYhSXRKyi1PSe0GyTeQ3kUo4tbmKltZ4uJY4a8NQUxTEG+znLlikNQRLtV
QXJLAip7LTfU4uxgudZWsS6KVnrhZpFqSZ3qvHWEiSpTrtvvIt5buZ48ZnFV/ESj
dnQ16xy2PJsnvQj+lUcRMCE7ACDcF2P8UtO8iqcAw+3KvnxYtDRYfeEJzeXorWTO
PPy79cU3Clz29Q+3NCZ9Mr2RZSTrfz/mZ8qhZiZ58VSPcZfgcBoKRtg7XM/w/pYh
758dcGQCdONzsws31Evh95LNXw8mmC7YqRDjPq9MTivHS42SZnY3nZod7wsbdqa8
ZQ944AvFwPBMd5ofI5uVrx4G9CA8N8nnWn/dM1lVwb41NbNon1vDIRxSPceriPgM
VG9HQddu/su6atklPwW0KNZFpErBQuBort161wa+5aQQdoaRwVY1LSb50yaAlVIu
KRRKVfY+qxE8H52PrsnAXlKPfoezlITI1qxo+iv0+werwQofv0AbSE+3vNVJpTCz
UDS3igPNKHXef8Kd75yXGbcQPjti6L1REFbFQgsihAV52s4TRjXWiElnnzf01W2N
DnNQI8Eb6MVM17qtB7ncTktI1iKfNt4sAva0HOmB7suU7p60PKJmyOlTGaeK+mTi
Es/jMtAjhfvafRex1cbE02Ng3fnash9jVkH8Sbk3TPqudsPb1rQo9c3sFo1mkooo
Wk829NIk9kyJ5Zko6tUgAFh3AwDSlXt1eexip8kpG5P/kJlvASqK/Ym+OoST4OZK
okUtm5tUsuBG0Q4Nhj2CZAELdgVd3MEpqg+qU6CeP/VvElixqvgJ1Qyu8sFvlEFz
sE2pU9cgevvqb1vgTVaa3sehDLp9TMICUvVI+8J5+QhIxdji5Gz4kio8FbhT90dY
RzKwKLGNirFOtxVrGCkxwRz95YcAyD0Ev+hSCYygdZdvT2Sx4myRFF/hKRrewGLP
5rvj3qewKbI6ziqLD9x1zsrmlp6/AvZhWR1cqAjsw1wlKkg5+6afoqiI+J6YW8Gs
fnwkPkv1W4lqSM+VEJo24bDRMFIv/JiR6j0PkudpDB3tjc7qYLgt7squuhJg18Qm
QYXKM+w3YHI5b5nIp/G/V8Xsavx2CvD3e8FAI1hIRIwAxOMAo3APrTL359Q2YIdc
+BZMdVDJBSHM0oifhk+J8ArXEpeQUz87tmLBeydJFb54YoAKVs8eDF4rZxX0fvha
1hH9JIusF5YglIzqN5h+PmmdHmDbAKkpvJ5VfI8AZKcx6+zkv9Fx+O9+qcB9omXi
4LfK680aQm5NL/gtk5v5ntdiLHRKiSKAe3AKenMAPirc9kAGnFSzzwSzfuVmK15k
0uGAfnWNesUTqn4I9wHOSHDHQhtnM/wrYyEPW37seRGPPJits9yUmwJbswkOjn8B
TlSwupcOydj0pN6/PXz84DsZjNmEaqIq/sRMZm0hv1UFv5WbbHSHQ4exB1r5+He1
OtGyiKh0nyjfgzDqYq9VPB/VDuLHhEQAL+i6JM9gVtdN/PHT9i7gr/kDV8uDjc/h
aNYGXZMjBRgmyFZyIfAZrJtQZUke5soLsyblTdX4mdLjEC7dyiTc2vIBUHVbZ3sk
qo+dStSLt4Dw8OCjq1SvUq6pkRBxDq28HKMHNEwCVdlOvcClzD7SOGG7/vNlk8NY
QsMq/bt5NKAej3AL2aJQj2ERxenPIYxEHkw4IQzOacAGo2sV2AkH6xX4VL4GSUJ6
lLvtTUu8/GBIPpj8mh+kgWtkGR2uDATsqeOEFKiVBPxDGSv9NBoz/eIp+Hz8KuHN
/oWp0ggoosKwT4bQCm3E2THIkHkJajo5rWCv2vSoRmdM4J1h77AhgxqjJynsr8mR
NnuuMZZ5MB+sKme88ewxl2S1Jzd59Jrk9flBaLu1tQuCNW5TVZMvQK0XYdPXKQHH
VTlvGdLMUAI7r5fSkhSdZnYlqtRINdzb9f/tmk2+sOrL2m4E/dD3a+xut+wHMASt
HstdM9JTmCQ/80D9soBwVGH0h3I6neDktsbFr+dnpG25UwaT7s1Yfhco3rkA4n3T
ab8escsaGszP6qf04Ug3V8pV8SJABo0YAZDoQfekfzSRTkslqFdpjM+I4ptZKjp0
ad26iZG8nxD/OsWrYmxw7PSlPFaL4G1nWBxrue6v81yMLph1+bXDlB5Idi6srRQZ
PK7ItjMfBoB4Wax9YL25OWK/dz4ONiVpdCuWdBIMMtU8h2ZFAyDMSh7V66f1jm6b
HAhdFu1qUp9Hsk2lZna2IB6VdU7Nc8e4wO6zVauOSqhTavwrgIx3B7bLsyP9cKtF
ykevsv6uhUT7Xi8hjZr6PfvHvCHyCcj8b8ELQggKV9z6/yoYZAs+eP2LGA9ipck+
SXyCbylVGosrh1SxFcwfmDrK0qRr9Y9UBOqSWhz53kE/rdwZKnpUIFRRR1QTpmSf
wHVnn1vvbWvy2Wptyt9qh+hp5tc2FAwpuKYga4hlSMaQJSZOK0D+dUAZJT8wTJwo
dmreMG7851PG4QHvQVXc8i34jGNc+cGNOj1DHJApvkcFyh/ww3CcjL9j9XTUNeDn
aZuPFhAKlNvPTFSvYa8dKj6l26zfRcr0eKFlj0VrX4YCU1HdQnL38LYOSA2ZGDo6
GAYq1h/OodIQrhm4k6Izz0zT+Fb771eoqqSjd7XOdogfBB5RcQe6P6OkOnbkMBff
6Anmoi7s+wRT3iyQWMyK7DJ42lJE5SVIrUYBUqMxvie08iEaaecfOhQDVOZdWRaH
w2zGK5VSOzT1YpX/yrpmskKMpUAx2TjUZ6puy6B1gmyoGQzHSlf8CFzkf1COxmtv
Dm2JifALtXNivpfpvugxyESNHJM8SH6KLC440IscM69mUQQ94xuCCCZBeuo0uEaU
500itazacVmlTE1ZAng224D/rm45UN0FlIl7fF9S+XUQe4uMioyUgA+eD6z6HQG7
xb4CGYF1vPzH4JNnyHcxK51zntVBdbyT4OTysZYgrUeiu6LXIZwQTiJrGCQDoJJy
6/1bPZCnaqXlSNENbrTHIu7aFFJxd8MJ86wV0xPG7efxtUhcvCMbYLxxg6IK4rNS
ncsn0ntjaISP+MeyqZyrJ0CCiwzcXV9rY+ThFg8qugEOwcsNcKDMCm4TgZbjAEBU
2468dntaupNV7L6OiILH68FvFps6hlLdI63jANJLrLMVGNRTnkVUro9bkVlsQkfB
kZ9AsH0fPdgXKiRNC+GPWkY3JKaXRyiryS7iQjNPEdivtwBvAd9NbvAfPf+JdRf0
+cMcmQlwwFsuHSBsY84DvBZXGIxz6ps8JKo6S8uw61JqU8a3axvkgAYQI8Uxfh94
L6JvZvbZSIt9nHytL4hMbLwMEo5IfS0Pg7e88HAJEIXK1iaRl5hAMxe1lg9CJc0n
TBDTJ8q7G45PHFpGiMmCfYNU6dIU6IKnbdxlfEo78MCGyVwOE4WJ7Gh1SFibgB8e
Agpi5NWXDKW5dC9YEfHgi78TnQTgqMsY5MYmTOIPQP/B3rjGbS3qQCyt5jOwrg5n
i6iDmFxqLCSL4rYl50+cGLG4m7wSZGNNoBVlntqvXCOfNbp+ViOjiJx9LuqHg6JR
b2pGPxw8X1A6N5XxUHr2/s4TJkfnYuBOxL5M5Bme66wZAA6XxmbTDsx343MSWS1b
tTvHOZwZJ75MYMrpeA3xHF54xMYOhALeBC3TJaUGxZ54txYJ5RJrCUvVR1dA1xVZ
RQsrTdfAAO+005UBb2s2Jvx8GgxxuUzpHQnTgwKSGp4GFTNYk83sTV/Z/7DZCjKA
meOs88iPbsRScNJnPL2TyzLW79xCZ/lzYXzg2gd7iLyG56XtkGuMBd0pesj70Qxg
zGgpfze9VMFqh6fkl4PuT6tAJPPgQWvgHubhFwIbqD7ft7UmJGH4SkrnAdA6oKzj
pZQxPqeTGEQ33uZ1LzO4nFRR5MObbw61030tcixifRX8eaSlfn+GGHzm8lHXqXY6
dCqZ4rM4x2Tygyf1JhiQ95iHvuGyr6p+rtdgDKcUmWVVN1+T3n7SL/uVvv6dV8r0
SFRAysL+6lNVsWJuhcQ5QcunmJLyK/hBOEjnc2krC4PBktpxT/BkHnEBWW70OT4T
kJfOcVQporqXfCRBVK5pkLwvKG1L23yoQkayrZBtGgOwoDNQHUKJpx0S9OZGlLjN
VpQUBCfeh5A9Xg+GkxMC3HKw0RTWbhUDFzZ5jqiDRznSGMK84HQH3fWDJg3uXvv3
LA1WBjPr6nDlnqvicHhv8EsF4uZGptOusrLOeyhBhxUoK7E5vyuo0gMJFt9QCuas
SeVC6vIxeiioI8LlPLk0lUmcg43HawIL97+CQ9dFPY1263Lc8G5aMTZYpLoz/WsB
HhxIwoNqX9elGmLvxBXcNXVhzVn8tFezJukyl8A/NX5EWExTcxS+I/l2eoWpVMX6
3rzG7SPYhYtjsGFCHXuu6jXqE5UVe+YfMmgQ5CpbQBfEYTNZqC4L/UWMOMdU+11T
/qbUG7XR/dcFRTFtYNn4+qYGh+6rfIT7DUa0GlnYI0QiCFGrc5/OXCGAuRaNaKao
f23kL3Q6YyNm0kRZQvCvzThYH7PYI1uP2TThpbU5bWB1R+Sn9TjBmuFBNCHnFEay
P6b9A+1aDVfcyepT7TqAPGsyViX6KW/TqcrxIy560Otb/xCkHXTsPF2YrY3676Ve
UVr8t8CBIwHOsLf7PVJ3zDCMybopa+Wgxl8BvU1fzAMBlc9ivymJhIdVxuLRQ9jH
LOLT+mqpiCIgSqPZ7gPD59cshCurPseN6Ji6VvGBBZ9HtNqFDr3hEfa5PzuH5r+T
99igSYr4KeJhepQv9VLmxXQ9UNyNJuPeSiamI55pIc7htKB+cK08XkgC9Bna52oS
NXg/ZZqY8739650rtHTqDpjK/a1mCnoOJAgTBt9HiFzqWWlJ0PT1S+F8Tb69t0vX
hCTPsFo4MrIhlD74C2lrsN3Ofj4w5MpAqeuAJefevj5yDu9E+PUIAaJxi4NZsQxn
5WW9t0vuHYXNUc3ZuF3F4V1SIIZJPQ0/2gi8LisiKY9f8qV4Xw8HHg5/KiKQvn9b
b+5HvDiVWU68iNEN5/2kiWFiUYGxmVzzFhTIxXJSYGxjMzstsoBmsUVy+SYgQBzn
o56iGNqxUgyFUOOyC50I2RxnPKXJSyKQcxvMZSEBVGdMoDQSV4/2tpqxD67pGouH
KJ0pnXi8RhdMWO7OQbaSynQUKNkh8vYsHbrQlewM9LUGTC1fCcw+idf9ipFeR3Vd
vExq2xQkK0i7nbUjKiFwNRP3c4Vi8j4nZQOM6qWzERXPz0ghj4WOUwEw1iou5Bcg
94/ny1x93MqAYZWoYy2iOvlqj7N+U8gUjFjHmGW7C0rtNtwFVGXiJVk5f2+bEau+
AROewQtx3vjPDJQM9KMlHl3NrKXCuudmIGOdihb7v2XsTMs3OhfHMDwRoktOS8RH
vH2WVppCaebWfp3MVHHcCPgoIx/4+ceXNniLfSe1TGkjysFotXKftSWWF1S7BiuT
WGBdDyeW7J/kT65lSz2rDLyOloTzyBijMZH3WHkIa8QBkHPTAx4ZRxwXxcTWXN9F
9YdvLbvqThWbcpDPF+bVf/H4oFB3lfZArvSMKRCm87tRg7KIafr0wphigx57gbei
bN8CcxYyBi9OtMpiiRs0ca2iha/31XyCU1ycDmMrj+kRpMQyjiETiY2d4MnvehAN
Ka4xb6z9g+oDLoma0nlim7vMfeBENT1s70SPe2Q5wgK0+rRE+quDx6AkytyUS1bb
YiDNdADfLuO5vB7vsM9IB+f/4AHJLoE9StuJC5N5DDfoVbdw8YYJpkBWkwz4ZYzL
LSX3XE653P3x5fgkCtdOsOo5i8b1N7DWkKrrOf7uJclqDmJO9MIJUrQvosIEpOae
Bu2jPJrTOBHJ6hnShLIIuHXV5IQSUHbO7dsQ1yC694kAIuvLOurxA989mlADV+xv
QbRtvZ61EUffhzAnzpdxb968YqjL4KsLysYSKI0jXtP12YreTQkczDxBPZz054GU
XGEMy9nfpeF7CaAodJgUhCyx+LLd7rzFeV9bn/R3GSBhUuaTPPHG/1kB4TH2R9Kn
gOghXGkBzbvsA9VbItsoCqD7a/kU6VKIxuSxXgywYsyTL17cTWD3ML9rJCiv3kdY
CnQp+o2OUpcP/0I4tQXSdIrGwpbQLn8WWZt28mR8KrA7Gg9IlmbO7L8j0ibbc8v6
fCon4v2xA51Th5M42PLOqsoza7IYQb7vva+Bj1OFv3KZ1vDBUfKx4/PkTOrW+2vn
uP2WA3+770mRwcwL6stpirpgnvxMDKAK+6kVq32a1bqRifOss1oOeOWYE9Kw5zTJ
YJkcRQq4WjRfb6IBDIOdNZw2A2/P4mYUT8Q8hlPWDvF9ecGjncyhNgiAzH6CU6DW
DoWyecVUawke69VytvDm47ddKRD08FjYwu88hdTxsVovvN3BgqbgCze3bWuoXoXt
d3+YlLC36Fy+qeGxvkjBgg1xwkg+GnLrnTsj6sNbOkAxek3I4f8qvSaCSKjeymvd
+FmKlL/0O6MbMH4G9f8PY+H82+qAIGCwCzfg0GR5bbOhXVEgqVnMUxnfNJkUSl7Q
uhsEaUJF/yMf3nlE4Uvxq2PloT9DO/Ng/kZwYorh02HNWKeAI2yGi38H6+7G3fWj
e3muT9gd8t3dWvkmjvwvNx6+F9HLF8SizvvpKSPYzywHapwtNWVC83Z+x6BrhPD5
yAvp+npjUDjb5GUeVXjMi4UKJ15UmGzoHqwj8niyPsJP4k50M6UA1yicPdyaLqaO
zA1dxPTT1r/IjO+hZP+eGJN7GaB9hol91PKzXJdn7jYVm5I36bYR8bAqZij/65Bi
G63r9aMebCsKJ4qF695RbTm8ifgFAqZiNJS3HpfBLZir1zYpiNKISJFl/zi/6Z5r
p2Qht+OsSoW8xr/CsgPakR+r4Mh9WTHJuZrIETVLXK1Kequ3z9NK6s9tQVQE+787
JewReQ4U+5R9KSuc/Chjm+++oRao76hAkZtQ/RyMZUq2EUSq72mW8A2Akt3HCUfw
ZscdTWF3iLbZtgaJ9mUBuBcEfhuT0RzfD/4xS4jiMhUnUQD//l4noI2GkMLO5+zF
XOzOYmrUenDKBWagS9IgrEATy2CaZk/XHhVo4kHTM7/8jr04OAk3valP5rwQE4ae
cmCKpq3OFeEZ1WuMQZGzzyZFW3SjjAMtyYed/EHZMxMyQ4/BFR3qXeLzT8KsTvmY
V/6ppo4pxK9/R+SyefPzd4b0oYcPPezgarvF1yrvemvBk8uLPU8i5dNnoVxm37mh
1nZhAE6LxIEHu+Dq7KRiLA0008OEfs6AyZPHSyFgCFiL4aI0d93Ycqs7Qqx9yHwU
55JtjWu0EX3NbNTnjLbs+1Pyrg+lUSyTn/N03bZFtVKykb7cbeoWcjeJcODEUKo9
QaBkYw80x/niOIhMx6jSYD6MYc3hwzqp2m2pwRWsDu7Jucks2hMi9VzIpAw3zSit
+wTmx4I4NV/GOW2aJ8zhTzbdC7RBmy06kQ7FfwJkBaJXUPldGpFbE0RnwFABpGh6
ksmPOBdd58aONtGoWDWatX9hCoUtQX2gWQl0vy0leXDnZx7mzj0HEVUXPjZ/Y7vk
zW8eRLg5fkj0KPLw6T4R4zvyYYqJ87oLUx/dBQqMSXd2J5g8DOHQ0NPg0zwdmUeW
2GJLzVi/zgNX4WNPQle5dlWwZDE/KS8Ex/F6MbYuLUxDZNHNH5vQeYDB0Gw72u/+
NyOHk91/js6CbSZAv/5jRA7BnvXD9P9SP1Y4iEDT6d/cRgxKFvuYcx3G6ndB9TO4
LFXy+oaBLmddh5r1o/MxQMiCzKzBosKfIOEhvxhDAfe3wbcPlfmRau9ZnlkG1NKZ
OV9FzUuv35k+LBokbenls0iuFeuzO2KqnP/El3NUF+k=
`protect END_PROTECTED
