`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tMMx7X6LoeLEjrmw0RNnfTXUgyDB2qu5t/zi7AgedOIwMMJkObMdq8yYtKChUevD
4xQuVgdzS2Y6wWmXuxpkmdBlNguzkdCXzt/xouZ1Z7KewYorXxMKVlDUT2pzw03r
gLWgu9HpeH12usVxAnHPlVwP6LNxi3wQZxSNzjPxW7xBX5A11HkXTw8ob5L8dSOW
q3oIZJFWXlctT74LpMmllJ2nmzxNj2SZffxiS6vSksQ8U3Udj5idebY33ZNavT+r
KGDHFl1Dvm926sgXz5f5ZnBeWkp8ozac7nrCKoRmFaVNag0C6lQ64rKzKHrdH82u
UJeaue6p9Bna/JZhqS6cBa53blMC5mEXIXAhMe0E3Rn/NpkoAEeqhW5x5+MWajEf
nRdTuhUS8WYyoHAJtcu12eHYTXnFQTXHxIlmp3d6fcaHkwAhMKk10EzUW62F5m7z
7045GjbcA/Q69C5ZBreBbAiug6OanrrUs2rFZd+yQu/rAaDzY0VnpEcg1izTVtAo
1OeIwY/FltV/JPiIY96BoEUxhKQKdG5CkotaNmmgt2OMFiDExC3SiM8rj9WZtlyo
16816ANOPCxk4INLUym3Tspuw/ZoJ8rSrXnA9p0FeD4GprD0magR8DqCDBdYqjwj
tXc+JNdKAQNMVesrxBDa9W5CJZhy060MEUo3dfYR0VQPo0EfhShRTukrMMwHgXj8
MiNTwMzoGJJBDyxF6wXJfMxqUT5NJHouuEnl3DWxRK1CCYciJ7YkuJrhK8dF6OJW
YVVnpxjZ96Hbj1VzkBF3rjEUiRW/MKohWcyHDV9kN/oR5bigUiT7jXWFNdgb6AE2
cEXorpOQ0R4+GFhlimIQSdyLvQymgvw6Cgwt2dls7ynyA83Srzg53ZVkoGUGuHA8
rktpseq5PCzmv9aNAL2Vp5JY98oU9xAZ6JxUu6+jot5LMLHZbodZaH6PV1ULNwbR
S0vIBLS4LUI9TNSR4f41arutfKXieLIZevXLkRQ83OvxeOLdU88sCPv7UNpPTfw2
DtxZ64zxuJSXsfqP1k/DfFnstEgLcq+HHVjFjk0OoEcPNS/WZzcQ/ycjbbMoRMNF
EsxC+0ZGBH1EgxNoPHrhwWINCEy3d1ePMrANZ3VYJbao34NMr2uNTxQoxI9qCy4W
qiVkstc2wODJnbLbL4DpYOSE//1sCciRRuLmDLbfS29u3G92lSFKv+LZcoKwp6+n
Dp9kJ7fxsTI/unQZQM6/bfWOM+Te1TfqAJeR2wBTuDCWL5zN2PGnOqV3+AixFawT
4KfC2O7w5NtcbMDZrw1CwxS6KS0mJitFcD3mvlt6+2sCvl5bUIbgqyWfUfHGgJR2
PGopsYymBQUUlEy1GVf6+B39b9IJUQlnYl7FLI8mLEp1eAEGp6TutaPysXF+lIkI
Sgczg+k3JW1zEIx28i+qPW2VRdV4v9zmmm2jpOJIN/tnCSR/k8FFlIrfuRBF5m41
ZzERZIeU7GCsIiWHjyPDzxqfW7SwPIEwn63B7e0gwnJ0a0fbj8qOle1uR1QazQab
L+wRlXQCDsa+Mj6hZo2WPRteEMV0KDlfiQZi/GxZTrSJnJ8/j+in5lEbdLOxRbjH
/93ekJhJKweyZD56xM6UdB6A0HLEYPp2Qp071Hb4Wj85pESED4aVdl93mKlKCHOo
6NP39vYGBCLc5u4bsZCuUUTDQ4k0UQruPEFpkyu2B0rebecA8OBrOEvU5OvCHore
lm1vHX09tbxVM41FW5LQZ0N5HcB4RC2wjmIj7P7Qi2v6PoOgePgzWLmRkQMNMS4U
yWDMtbwt++uFzLLHLny1Q0DTRiW/ve9E7HRqdp2iTwZ3zffG59RAKpO3jEah21eK
wxjtocCc+0tQDrSIRA7pS7Gq1hZd5F6g3qfvIge5pkao0KDN02otZX0tLho0pHG+
XZHXkUk5/27tPDbrKQQ+bSDRZTldOx0+113rr8y/BYs+V38wSZyNRSFgLSmYUVQv
PkrfdcWQvJjLzRGAdBiomRcmtKYWj5tZGiBD/itTF1ReSSewdGt6890tIEwKCITB
Ov8HHYRr0GUAwaLeMXRf/m8MW3ooOIIeB91lUWoH5kYBmLiEuP7epDFyhg/asHrM
jEyC2t1lyMf0r/qQR91TvH1A7GYbRUW5YpaeDvGpH1eClvbaaxbRnDN+WlUaQOM2
OS9tDrIwaOnZMf3VZKl/fjCCerhp5OlQ5Wq+r9S6qd+Lmr7Lnf8h1q0Qp3bRCGj8
Z+X/g9w2Um3UeKgIwu9mrpLFs5m0/HRqvmj4xo4bweqsxDuc/ujXYklyqqJy7Kew
+OZ12HMBoBr8LaG3BVTcoF7jpXs7kBkLuAGtpQ/QkbRId9UP8HbE12ePsx4xmy85
TYNK8KG3Cms0VtyhMHhgenGf7+SZiVOdV6zUP1tlNd6f48n/WQeTcJaQVJTs1DVY
JvO5jWdPu9tj534ADceHc29pYimk0EdY6yhiXAg24XG5hClMjn8abShHMNl4ZTkc
ue5wyWu56uYHCdpRRvAzu+QcpeVNGx440225k8Abmvb8a+hlpUPKWw8Zx9feCi9K
4hyKCT97L43fcboqrE8booqlHPJ490QGc3kyznLHjQv9nAXwcyAwMelvAdZoJSx3
mESZEnTU8fVH4oQ+mJ5U4eSFjbdcecCUsuwEbU4HOG9veSgfKuc1+stxszNPazwn
8A4No5/j8wKjhwtS+Xx0d30lDeHzYgt6dzvZDHUq8J36vpGHIBREpMRgQkI19MAI
/5uuIlzGeqPyCmGYfkUVAa4mPY2vZqqKSHsyXGIrHrRHAOBCyr73wkNKC30JOQpN
KQugMYSLxztRTbYYHe6Fh60Zi4K8mqfjN+0RV8JehbDaFSNl5hMxXurj7Hkh7Qgz
lu+3OHvEVIGkF7FsTLwC/x/DO2o3a5/nthAT7qw2HT4HtpwMkP+m4+TdRC9GpZwa
Md+/mFb+aZ6FiDkumqRNKXk9xgLpG3IIXzBxu6ACiPLu00DgcLUkKVjHNP+PZMKC
`protect END_PROTECTED
