`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DHb33QWOsWgt2b6Aop6m+EjTH2LcRKdFVxCxqw5RIu+u1HrGs5wTwkO9ybxgJTe8
tlZEe+ZhBdximqPu9bch74zBgaQqnvE7Z59bgGjgWwDYcOs40XG5F/mG+oVgau8k
ceD5sxxpSGDjoq0UB8+ZIrcJmVxvUQ7Hrvvx9Q1xBuJTvkjiN0uE714+5tr0OX21
jKI+FkhcjdtQZ6AuBtlcxl2KD+nsoa4mGuyWNOmlsGvAltms7JBwXOdeFcFGGG0y
`protect END_PROTECTED
