`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EBXNHwBDr21BWDPo2GWV25YYAJ17qgjoeZn85GpykktDXxpqbBnZTLMRfOgWJ+8O
7PZA84VcfDHFCqFzOxlH4OebbvKl5A/bnawLoD+AZ2KQAMsjWxrYM8Q8aGySwGy+
parBsZbuTolsZNJ4vNqhXMZvTcVyRfol5oEwF1LjfK8koQNqYOX8C74D/taUbO4b
uDxqXi4duMNSQWTbr+mjY/3QzchTPZofVdP1gUQKkk3y6a1r3um4Cepzr5T7OCw6
0gjbdZfffOo0RY6lJeBdVHYqect7enIgIaY9zonxS76p0RptfS0zSuyfl+MzXCyZ
c3FqZEv8dXHKV2Xd7kxRz5gNbhXtdBX5SCYZykHsbLy5/K21HkGw4FyggpQEuG8G
ONatzH8nrDN1JLVt853JRRcEAWaSbD53CkyR7WS33E9mo6pm9uLp9q0brJ7aWxMl
`protect END_PROTECTED
