`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vsvr4hLP+2CziwiTMY7JSS4aCvgp+CE3YZ8JPCOS1lzUno4kMunuYKnOMkHJIk5U
rRX/DeEytOda2W0UDD6cgUZFeaOvDaN3j2wAC+JGp27E+jZBiTNfWbwecC5aBO09
Yx77outcdtsQ3k9fGbL89te6k6oJBohmA36/9fomuxLKZA0Jho8XG1nv1MULlaOs
FS+u1Z4XsIpJTxqS/5WDCr0paOW0L5QwueBYYj+6tnrSDEeH5qTRzG36PwlfGTE9
JvEA7ObB6lqoWZ+Ss+CjzA==
`protect END_PROTECTED
