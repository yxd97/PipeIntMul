`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q5mpy5h8ueLFC71Np7HsF6mXYiOOAaP5lGczP7qR1pXiq22kxmSARrQFe1vEPxMR
IKhPTn6AHf10TqUof+4PcZ+RX3XbtIy2WaRSa6YVxpDOCdrG//lYR9W7nrnggeja
MeuDGhW9NZm46YQJagtbnIWQqXFsOIRlbCjQwA82WiLylxuSciXgy4My033EcFmF
fy9RWWQIjRCj34lbUXsC1+LmooOYk1Vp7k1wl9QlLCEvN0F5BRQlYh5nzLv/LkiE
BFo9gAG4OEtTtpw09WXrpLC8+QrBDlFbRu8lsNbQgk8dt8a62FzdK3MmTRN2t3ha
aEuoVfqeIRAEWM/UNXNNIR+biAi0FsbZ2/CqOsvDztviXtBYPVokIq9/y8MGznBg
bich7b+DImk2F1jJ99rLBgwbFwAdQ8+bXF3Ge7s+rs5AiPCwqVceWxOQRRhMQSiz
v5KrvZWKxyAaXC9sxBgZw6Kld9bQCZzAYXz/so7gWvSbo6FXBB+cfPSYkvEfeVPh
YBNDT9lSIXECFmq5d3QTMyfUxpUABzWF6V6lK+WaVpQvMYPTqYUcdRYzkRrMmuwT
zD3MUaV8jUn85FDbWiTKq7F6jiaadQBpfvFn/cqOtKsLRKkgezbuLYiCxP8eASdg
Oq3qJcbjeUKDk0urYcgO1C4SrvXMvDxCmybcU5EqXyNRJ2Soksq9lj3gwwESy8MT
w5Gl62s89SZ0Ai8EFrv7IExt4z2LvfHA5FVt32H+8D75zb0uZOkyuteI6W8nZq11
1MJL1fZ6aP+LpYPCSezEVzpWBwi8OUi/p811mEa/y+r/3yfDNHxU3W/2p5ncYF/u
241RQXvFW5nzgmBhUc+jnAUxEtDCJM6K0Ct235jWpfstmTfdHz0XOm/ZrXNSkms8
yuUhp+DisqKNkc8X+Updmu8QZrOrwcarAIEJymMaGaQ3eRm+w+Q4qpOekIgEQ9UM
n39sGUVRgc0XlCVkduoRZA==
`protect END_PROTECTED
