`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0qusBS7BE3zmLmyPDnE4w4vWQDOthSEoLCCEQGGapFZnqvLbQGheLHGYbL7sYQye
trl4r8JEDkvncA8owO0Q+IqZ1lcNdgKbIysHQb9cN6LFjq98o1IaNUeEWBLKRNsa
a1KBfIVRQ4GrGnMEtbq5AyH6o+OEkXD+r547pChC1ak/gl42IVIV4XzCYPTFU3ux
5Otzf6VFm2A5iBwbJwEBahhxjYk7w/IA6pE/BzvaT4S2H3PYNmCR6oAIPUNbFvB/
sLo6/Wf80OIn24TsPQP3LlvDzwZvcm+eGLg5WLOO3q2UOhqmbpDHcsrV/CYL1akU
7sZimZ3uOcmDVvR/7/gswQ==
`protect END_PROTECTED
