`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGP2SqZuBZJ8h3U8O7E6+0lJHfARb2627xygAm80oeE3zbo+1PNBcb/Y/J9I/GIp
wXqsPGk2ukbkeE8UXbQwR3FU79p3uPxi0OKixgQWwLT9QEFYu+d6qwnXAgFXymor
lCeCOkLrD89vgE6WTeP7nu4ZWZvEOXLYNjM87GY98XChZXpulZjvFfv2Sy5mR74t
ySsH8XpRRO18gLzaOdeP689Je1lko7l56cXOJCLl0rrMxYG5AwAKEsChPavoZkIi
hmx5qMnySZBxWSzXdsIxt/Q1soHIhWyuTfPfhSrm8+xLYks39FJnPwvU8WswkznP
IfDLWhN6ddaHdVBJSEtOhRrc3eew0mF0rtoXShZ1sE1vFYDd8JSVGbuXiY9tCRmM
4qVpDlIeFok65M1Y/A712WarnKCy0LUmfrHXMBDpCeeGpEU+kex79ZhB9lKKO3wN
3LatuAPzApRW3WQ6dzxWoj7ziDUM7RTWrafgFiqxA/5cPNebXtdgZh3Or7kuCN8m
FUdIaoo1a1LPyykKWu2GLXXidwuDUDhR0KYeE+RGWz8Uv8AtxPZ8BRvAoJAs7Ayr
sU3jhIiu375hE/407Onlh9SFfOtVFmuMdrTDkJQ2SmvtmKIaW27WYru2ybnCi0iU
ovJtA/3N4aZWCQr8M+GvRnBEjQlEb078eB8tbR04OUtpu/d20bHatYUnxDW+Vh9y
IpHECiDp3OinQhZwvQCzB976Yqh6JGY8j8gdzuWMk2U1slJjnBGidQrLrkJ82sfM
HI//m42eZz9ksjEOjoVFRZ4og+3mugPOO/6AnvDYvV2kK+qKBFEI7ocI+MBR0kzu
9DFTtTd42I27aT++RDCHpDhCwZ+g/M8NfbGLCxp15zRC+QQ0oekH+3G26ETEYmf7
xXjT8c5GiA8QMe0dQMGaWnGekR/Ldq/G8U9t9u66VMHzluKfNbNU7far0tIsabKc
tXILfFBn7pfDnWfHuwtpELWP1+KC85u/8lhUny6VXKc+HMDHXIE+wrt4kVmWEokY
MY+vgvx3qwUnIdXEh9QnihXnQ4lH6XeqBpqNqFT3j7fctxzMEVC4WMthjWYW+I+n
d6yZ8/fJgLHI3lfTFVKakfNiSZJSew0iSLCdegrgi9nfAWkeV9ka6JJR/AtVptBp
cDBpxCL4BalovP4bnBAtoZ5gNXxX2jPYi1hJwp9VACqO9aJOsvAi/pSOYiCZIJ91
f9Kh7VuRrrRLtnZ/ktaXcs1De6BR4qz7lZD4+AzpebZSXPpEy4r7AWpouvXbFg0+
ssp/H9IY42NQlaLu/cY5xNiM3FNm/v7Ja4df/jbYKnEDw/0KyeGNNIwNR5dQeMD+
t4L6M7hvAkP4wRna9ErDF5wwhEnJXAyVuyJNQPrXrly0rz9TGEWVpU5Gcu2n9g5Y
PLbbCA9TReFjLg3agNF5JcZTh4LFZvhsNvufMJtLf/vtg3miOVepxgnBrQ8VrW3b
St/fIUMbTu9M2LO7PO2zClZ+7LjZrTd3qvH6e7QRKCX7C7AjNrMpGVYcF5YyPQ6i
ZFGgTRE2kg0wM9eNRosPPXlWTWP8Kbk4oBJN7oJPdHGcaSIIK0awHGP+e6w/erda
2Y1Ve5/87H3Lkw1uFaVOAn67h30j74Lkc1xJtwWt0xyYSRXh3vBSjVBtPxbQw4Sh
kitVM90vGIwzdcMRWa0UuYhGtAHgm/O+TLg1P/UQmvb8QIX28zSIHiZubF2Pdd1k
bl0Wd6dymueI3xj6BDXxxKubA7dFvzP0uE1V8Hwg1FQSRZxQEUZ37cKTXsbe9lkJ
eJ/e+Uf2tlJlLxmv7lcf8D3Dh7QOCZ4PUAIIN4MpSS5zVL9G0KBPUMLGfrN07SKg
QiqawNex2LtYdjuK2tnaXmVcWauGbr8RjVbQEOlZ1NlfnvQ6dkmr7PTmcaPrxfuN
jy9fucvxHYSZBk3d9Sgw7rOZ22cJ5d8EqtG72cvwHx9gxcMghj8QzfTCpgx3HWvB
dbSGET8H+g5QpwAeyLqHu6d/CfH/04vDJ1r/XPWdmgs3lltZPhUJAcWgu5CW4M6b
qjMpMBGv5BELmeRS37TCcL8WnMhk4RUS4l9zTLW2I6MlLruOWtvsXCuPwD9f+yLX
44ffw33UAxryerYDVwEiKIiMIFHaQZscVg402vMYdSnV4F8OpP/O5BdSzIc9+COK
rHP/cs0xJlcW1SKI0rDijjBqSpy6tAaL6WPPxF1l2h6Z2+nF3V0zBs0+JVUbfWqM
d+J5YQOiNdfl9udBM14XkNN1F7murfOryRFgoz9KXPRD5a2/Gy3xg9dAFIr4NNYd
kqZjwWqA7XqcxDkn6xDDzmkD5FyPsfu8pk5zLQcOPPEW1RdGHSJxwfxCUNwMlZEi
Cmnhr8dTKq7tG13Qx3l54QYLHTD2bz9hvRcVV/Td7pHWfyNy0ni5iR5Q1p7stf6g
/DG9P2J4Sr+aHKOeO2V1lJSOU6XQ3o0EcQ8JmBTHUKc0dgGCjrX36mAsuO1dmMNO
kWgbSTeC7dQZ3zYsK1k1+Tzv1OgKXAQk7nrhkboRtuW3zSCWRKDN3QwsO8hDy7bu
Z+tkeGUgCizYZgmaOhboPyD/UY8LKPPSGANxJaQj4Hf+xmI14hvRJRgErDL2w7UF
X6UDZWNy4mSWBUYI1Jsq1KAewxW9c6V16mRO0HzHhy2PXlTCgMwTQ8S4dSGy8Sir
DdofVU6RwuFFJIsZUMGts+nYitXNNaURd9Ps9GoYEJXTwwrZW9qUS+8YMdUiSOH8
gUfXUWl/7eW0PhT9cJsf8DNlw6C+6ooqVWDJ+pa6KGptcbJXQgPVgIv1OE5ZO4nn
0FSHYqRUdFi2B9DFLnycXhPJO/B+79bKeg2ykNxjIIaSv14LW8BHh3nFeoplW0vg
44aSBiIxt6vWRlEHDQFWMuOkZlgeIFaQCmPBShqozGXS4jqsSfN8fopsQeK+b+kZ
yJrEk4NJCHq1S1W6yGib0HHYXN4ig7zLifCMA4/ZexmkgcymElDbmn+cKmwXXmgr
UuzwtBblV3pgnYFDt0sgIDyIs2D+BbKRVAjnv+NTqe3MJqbB3IxcFlnnVNZ+Pit/
z3pUEk/4YevZ2E4ngVUgqLLlB7TK8Z0saPl800H4KmmHDfwohGwAyiKIGm6a6wIC
/OERGjyuOeSowX994vF30MAqI3682gaolRKPFj94oL6fCjMwf2I88phIzjsHzJPR
RJg6Ke8V64063tZF38aPNIOjOhpF4xvqtsCKXLK5YAIf6hXxMO1kSclW0lQU2JMm
H6o7SThJqqrYAuOAYn5s6lzXEK4n8sjFM33Ts2Uj2DbF1go09Mtox8OvUuI9iXha
rHtqbCBK8D+e/hrk1CM7TbuMvhoDNH7U5FSiKmYeqDVYCEYb/kyTQOqrXvKFJCAT
4dTBzBU4T3W9yuw/5oLK5Jjt9tngTFTLdc4+spKWF8BNm53DhaooEhrL3ZobJlHP
ZlkY1kkWNWsiE4BuUJPyGfKOGNqrGMMgwLJtGpbLsHNwz8NMgfMnGXQXJ4SAvvvr
pEfRFJXoAAfTiprOou7+rwzJ8DeoklYVSFkQoq+K1Eal14ZQV5YJTnwE+YfYYzDH
6BWC015QL5witdf9TAwA1RbV5EKrOLSdQAii25YUSVj6j7Ax0DeURdBq2V/yYg+T
FCLX6sEYjeF+q8yaA5PkPNuxwVQKPUOgWqK16bxDvq7NkSIO9avLZeh/TF7NU8v2
+bJJzND5e/e8OPoEiseQ+/NwFQPoD1hgCynjcphHZY4wIwZxJnJ/Iydux9P3MZt9
Is92b+fSc2mM9uc25t7dLnrQFxR7NShAVFtcot8ZVrlivN6mr18sH67SXmEYaJxo
hpPQ3uh09rb8v0E2garc3rBEoMIm1S4MJzyGsOW+vzgwWVrtP0yY2O1MUiT/79rR
Ww2nJJdioSbG0KLXmaX2/wTovRCw/JLm1mKVVt44SuWbUGsz/vW/02knUJRwEEPV
6N8UGoG37TlCi3fZG9EVAJWPneoKYuoa5AuqYhPyIsSQ37pgwKaYhB/ZZBmJX7j1
dta3jcVvv35sGkiyrOvbtIMTLD7YOsNACcaA6j8owngDJnsRNwwqmX0+EXPszIlx
TGa0VLaUgeCwlKAbtsYNM3XRnHQWvGERoJNCZpwCTfpOSaLEad4/v8isCsj7Chh6
wrfwAabzdOJPKrEaF2th3cNbfS1fJYvpULNEqu0k0HnEGhgOhLV6M5CVcSzsHUW9
iR1t27LLhr5y2Hbtv378Gspcm1fXBB4GH6zcTbi77pLQcIzqbpUx4YyIObUu8Zg5
9WlMcOWy3USFIUVsRK7c28zmwpcNusM6lPMtx/LVGPX80X6T8UqDW1V+xPWs3sMr
AQtAH/mIbdAiLqI5asPlaKisfD+qgSsrQBB14yjzcWfB71VC95oJW4AnhfdowD6A
bY+CD4bbmUv1Q9NMm1rxnXIcE/ggf8op5MAVBNSVjxQtRlwcfjIDEqiwUnWWOB6c
btvjdCR259OhFUQ2X2D3BXFMTvH0BRPRXz8SDI9fZaK04VlqID8mf+hvRo7SPSQB
JwLTAUgwx0kxXbzdqtcdXvlkZxPdfN9Mui9RxP0jDm7lHMWG0YM9Hc0t1XNxVdw4
AxVQ07Ww625REgU5tI9ScVBHWy+MKhpHYQDzzmjAHP2UI+Uyw9K+E9yIVStTGzCr
LD2UsI5ZKjo3+iceezQZdF5+/0g3zizP1IjRw5VY1ZM+D8HttNn5wZINNPqHyGq+
Ji3Rn3no2Gr4IACMaV9ipE+5ik3M48KkeJB+0IwEx4CELh737RFCuBtdqjsvxE7f
xChada18D+jxd0fKp016/lbGMWR9pRYbN90pNvjJi0caZitk31Yf5d9USHY0USsp
7StIAHAg5TG9QN5FeHoVeSN19zu98JSMLdJlAt6XBENAw/JT9oY0K0AyJponZAwf
qbT6Bgym1rGTd0oNaXDgUeBv8rTwRN7RlaOZ8i0RB12kOwiyXQz5EQs2zi0On/ep
brU1b+jtnNAT7MtJQcZMl5Nt1C99QHNTcCJtVNQQe7tef2sUezTAok2RHzLdHgFj
IpZ/+He3WFanXJ5VfWqfq8Mj3QuTrJIemXRYviBgALtDlfQSPu/XSeW57FjANayz
BRw+KumsW2BOZH4zAVa6+ysrjFZDxShtX7dZr8Eb3vTnwFuFo04Moso2ONvxau8p
UNNa9QcV+86aWG3THi5j/fqUkB74CZa6cNT8Bs8vjVpiJfMQeUA9yizsXdWY2+bI
GMb1QFsp3hdlXZBmoI6AZAnqpE9ZBOanj5Uz2uID9EdultXv82fdABuUudVPtRQL
uKC/N/AgR+9IBN4lbWRhTs0qho7Pp2x6oeSOLOshS8a1I4g6iLvrnt5Ly1EijqFb
eVncyUtpdz2eLeql8dhFyZ35QQ7AHOqMr3MPf881Cz1mGoN5fjvsx99DwJcUIMtu
CvXLD+E6WYGJyDYRogf9tye/nX5D35fBiqGcWhBUow51ftm7yKjMJkDrw2KOe99F
GqngQMvnT5gX33UNY6Mk3L4Ypbzr60kXMchZPvSJDmY2UNz7J03Y9WstrM7rogKM
sCXxSqLeLuopA5XMGuvL1Gb1ZFgqWXFrAtStIkeyfvgmW1+G+12Ti5zgJzOpQuTO
gbxSv6j8iimXmBoV7KrFpasquKPOgII1/gDNBN+K1Npw9SchRhgBFKaNpLbBJz2u
MNEwmDrlG32DKVuze8euVAS2Gxz9sIRnntuxDCJyrlOQyoHkwOcq8GvWaiAzzeDf
WA5WTOFj3vqheEPp0R8oKCUWdbOs0OYeVSvjAQUi0h2YUMCQsRvkrIVbMLM2eUav
ed4s/oN+Y+IDvP750zFRD/hWD4qUHhbync82uFIOmKYdqeuoQpk2WLaDL5ssy7rT
OrCDAjG7/UIXjOZkE6q3ZFFuBltDs5hPQwbMc6I5CUlP9RqR9Yg9zPeyohWQ8sEK
brZld853YGwBx901BYyhVWambazZu3He3Rp9pyjRbL5/A0qGUw0+ZoXAE9BkAmuf
HZ3wwwdIh1wLWb7Ueib5aSYpgyHNFx7EAuHdN6HY66qN1UwD4O1UDTwt8cxKuMf0
WsrDNe5tvpLxtJxcqf27E9JCUZ7rIP1Vn196c58SiwuD+fhmghJhGhT6isIJ2ofj
UAGw9Q6dlAIFWfXECm11I6KLvewc8rXf7UDZcj8wIpUA4LVRiGvBWoyJoil8KW/5
VNSoZHJ0cX/ImsGCXLFsJbmdJIqqQNVZAKhxN4M0RHafH8VolrQbJZfGsklVRJWw
bc7PeVcKdamey7QV5SiT3VyaF+Io6IcL6/nP9QyiolHFb69+o9fRWPkjH8lSU/4E
vOC91gk61xW7c6nzh1NlDKTzrCvHWyMrgox3WpEr1K8Tb4DBo76AP0Nkpp3QWGeS
DtxXj69pLaehbv4J26R3DB38Bt4z0yjEO3Tu+Mdqiuq7TgfX8xpvQWOV57Tb/asS
DtK//Glp+paT2E5IflYVGyH+stWCbXYAlqO/mHM/q4RLqDHouX7FieNAkvzfrGh7
A3eVdVIRYC23JAapY5ktEQLvvfOQdTiAIPaA4q9jvt+xcEKg3vwmmEKDA1sZCnqd
PEp/6Mh3lRMiNifEVEyCq6/Hd0rbC/Sig9Fs40pRNnKoD3BJDA/SDFVM//pg1JME
KIiEhBKY4JSArTrx457sTcfK2ghS/tbs6ey6QSg5vXEWONcTWlKwBl5P4X0rvkQi
4mFn2MB9zo3pNnjV3Sit9wGk/8qLSoFpD+6nS9lv2frUs+HWQRbFSt5Swd8DEmS7
AioL1VMubEFunQ3DrOJmYu+M64YJZAhNhBs40SwApOAFqRdQBaoAFBn2JxjyOwfY
Ndxxnv5KgVtk5QFPkj88/4nuaMDHCPvtVTDqKORekJjuZDodp+8V2r6FgSPHzI/h
SBAwqedipr59DE4wD76HxqhAaYDUIWOdn+RACTvYbvkaUXGWIYbKDIjxMngemWjQ
GRek4YoPDCsPAki7ua8bMastPfV1gPfIgwerlOtLIsFfxwRIg6GgyBFSy8oMSrMH
323IQ46lNQUJzI81xtu//FYr7mC0lFPj8gAq6DPFy7XX1rQuGD/freArIe62aMt7
TKb2sqNNsuYXXnJYIXNql6+BnC9xLD01XAHX1SYar/wqblfaYFYBNIYAAc7mMepi
5V1eukLOrHuHiWrvRvMGXn4v8lZ/3YhihiF6I31gAeqrIw09Hlml3Z8D9NisH8XP
1z1/apmH5+dG0Jwb1v4yzYdojH9P9voJepJCQ8iIye73fTaqwMXr/MxHj5VpWN4E
OEnYcvd6Y5olE2qrMeyeA2bzd4GQlXc2d+WFmo30pXOaN+XPBLlUhLB31KG2nINr
aNzPwQEyNw6hd5RIM2ez6IMyhs95XsjCClQjmUK8m22Td3ZoMXpgxfZiOZ1luGHq
8GR8CY2aek6eQWfhhp5kyc2SpFeOAq50BVD8EVliWWdJY0pTOYwfLRn5ajRMNsb9
dEEJx3ZjKZDZlYTehIK6bHmBf23ZSfBI5Q9t52Z2YwD9FTbL9+xUvHZwGOEQwiah
Sxo0sfNC4XKghiuiUVugZs4lzsc75nzeFJycOAYQV97Ied+9JGDvPpRg/Nr36/Hs
TFyOa1tjq2qvxh4tYr8bi/coVHNfaHJT0IQFau6Y8x/Ebwuu3NORnNoTOcF/40H4
CQ7bBPcBrjfMdEqoiFSLc29eBJzLzPT5Gx0jW8/T8Tc8agGfAv2S4gzQmpuRABjD
uq52/Gc5zd4+0K8Q0qXpPqceEBe83wUY1WWCpBqs1sBFjjKeNN0tGx+S1GDZ6bdg
7eTupyyDftoYID0sKZ27kXQUu6kHSbov+srgxj8VRBALWyrwsdjcLQUXNlo29EKh
q1oDC+N+EQxuZKgtaraoLXhr4Wx+WIeCC2zuX2gKp7xLHhHFEaiF67WsXlg4Cr+M
v24SlxiROJPsM5Xe2AY7aUpkWO0bZAe2t+RFvDbnSMa5fv0HQceM6xr3GURgRzxC
scCaToqVJefPZOLCs5T1cF9Y++2xDCkh0D1/73IJXf/HEpvVgSDWaWvXeBTbK35L
hGqpNsszUZTnhWB0eGVAybavyXEx6TPQnrDhedSVOm9Wi+7MIgVkrobIzU7+0VxN
wTfjDvrH6YYPujm1UZvsg0bzD6ctTbCT67IlJYI4VRiMdqZRHn6VjMkEd/UpqHNa
+1lb3oDuXl5Ish1ikmuJz3kkFmXUbOwWZHraCymdFFxVUbVjFoGyzc6n549Y7p8u
w0W0RN6uYnyYpKv3Wl5TP2QMG4VaAID3WHWBFC3+NlPrtWkX18Tq2HGaiNR5JHl1
hU5UqSYImRDjCyz/o7j2ZkcW3Pr0LJoXNNXS8cS6hJf2e8h90zsIw42B6bz80253
WWn51l8fWrfhLQ7FD7EXIBkeHCYp1pyPdjHXG0IrBbQnfArCOvd5GNwlssR/hZzi
0N/IIIed+cuy8YHWg7rNGYRArXn96Pn4Z7nkXWFfj8k=
`protect END_PROTECTED
