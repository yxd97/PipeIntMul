`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJFbHcz3B7O+PaJNEUxBSI7uGGryJVPceJQ7W8TrQ83SFZXFWPA7MuLDpJjrTdQn
Sbm6PS2DUWCdjy05fCshEC370dL9tx8Dr022gppS+0Wz6cNq1PC2mFFgK1n8+4GQ
MEOsShslItUeCzkH9xgVW2pjWmTyD4bktP0ycognIu27Rzsg+N7bVAGKihJ9DN5Z
TRo8x9GfW9PepFs4C+AWaER1+kUD+/uazygCoYvZPhSEp4ccOZb7qdbdxSsB1KDa
6f5MAPuKAfPKG3hshkfH03d5Kjhs4CsgiqLaKjNSjwLeAvBVEWrl8tOw/wA9wO0Z
1pW0ah7wwT5li3iU3sMQSAeYOTwB9fhREkR1rNVpSkjILtX7s6qZv3TKE5PGRW8S
eW7Z7hXw1IyPSzQlhJpgFT/Md1xuK8qiypYgkYVFLvkAGxIjQIRh20VulwffncH0
ahVg+HmnlHAb2fCt23cSffhQEb5VjvR9SyIVQlvPqDEBjZ+JFVZKYC5/HkX1Xmn8
FMfo6NkU/ATunxo36p0pdq85brxnSf/PqlVGKsRhbfm5P4JiA3qTD4I1EGU0qbq/
ZVAZ8CEeVq6h7uzFjx93+Myoy/WyrqKmK6IvguChYu3Tfya0TQEM5OkaQwQ8CIXt
5OBsSuEsNTItXrwLsfNNKZPcnYpJKTjTrJBbITbvWiEXPVSXodAJtW/au/NyO2Ng
mqYGjQYH52ZcJ+MZc7KVdqtxXViWKr2Jh2mqlQ9eDDRcXGAocoqubg71pKKAPyu8
iyppOppK3UDyDG/d7+dJUDNdyGEED9MveR4kq5DXg2DkJxRRZiz9hB4N2Sm81uY2
LMb3fh23mWVJ5rOV4wgwefilVG0lJ+zf/Jlpfnc2P79EI3sGTLNeVNFwHncinLw3
Z/jEkCuVOuXGc50/GDQITH+r7YbcIeAwiUJ3frea06oa5EqROKP7eiXWNBNoPUaA
wAamlz6COGKZo9it38kSKX8jus10INZPFiIW/qJeFcadtrC201bNYBONeXrMUwk1
EYoPEf50sc3guf7/lg3xfq1HI2fFekOvSrhat4qBXCyOs6X7xrZ8o9SK0u+SRJJx
JX7bvquEiu7EsSt5rHCO9pZaNTaWrI1e1qXa3XFjduUQ2xdUX++AMsJUpvu9nWcV
2+TJL6J9AkGRdhwN/rh2pZlRBqoCAjBQ0IH5RRqSsuE7yB7FbGICIzhNh0ZDg/3d
WtHnHUwq4gl/bsA3PzY0CVKfPus+uM76xKXvSn0vVBDMJlQKDPq9Uu1sJRprTkXu
Mxk4PrhliTG8nRfIFNDdkaaDPAgepOOrW2nmyA5xhBx5mHhAFPE/T3ai1MxVpnp3
oMF9MbvqQB0qpArqowuiwdmUiWKbVthCNiKfrEwfKn0r4b1uyEgEh2xn9zqYR7Js
6u5KIGvrvaby0j6gQod+W9NbmLpYhsBH/7Rq9qtOWmrYSRhk86X20ZUHpDykzKKR
SHF9VBDN3AfmWCU6nMCAQHTq+w/Tje/7MtZOl/PlJU9deRHsEdBSC2SdjUyAhXP4
11Frm/od/KRUraKpm1FgO5MQcZ2HY3Ud6U0mHWWqqniS66oWo1cCSi97BqqTmCO9
fEJocuQCx+i0yg95s4EpbKmX0lFjenJuu/NA6o4xbfzrAS/PfN3kJnaG+z0gDLDL
z92ag/PLmIicsKFA3qWJjTR19QI0OvBI42ZUj2bubY6eqD+MvzP71D19MeA2squA
jjJ8V8ch/MYYK7KgZVQScLIsBf9HYefDkIkYgAtzrLtIHRr8KfagcDBqmnXs7Zdj
9zZxM6+9ffEk0mP6lOXpz2IRw8OdHiYmGlrW3fM2nXZ/3wrhmHgYxCipaqaLdksF
tph473dkDtzMULImGI4PhTjRi0gkAj5HCXEQDSUfzIGQ3w8/HIFmTO1yjn/elMKe
uWZkYD4kLF7Gfged3houCbZa+U/7ZGfZ88npnUvG4ymwfE7HceZtKZKREQABnp9Q
DcEp7+B3Pje4nhI9crxwFL8S4Cp83uDjP8/e3AzyyyMWPtOaiRr0uSbxpDisQRz5
5r8QD1dR1w9NirqQAqW6FQ2wlx4pktoXyXwB+88gcPkIJ7IuM4wcGKV3L/eEKyWf
gggWtVWFhSWg8XBo2/HM+uDGRBlahFiDRFPZh/Ce7b9gogG3wXy5hZP3C+fQtWve
8D1IsfEYXUm7IffUgVQy9Wh9joVIASQzWeJryNa2YzeS2xXv/n2xcK6mhHzRSmml
wod7OFBjlCReIxJWT8sMz21WSdM+OIr5FrEz4mXVqsgF6rhV1OMXvH3TykNaPyTf
l0JPFBgMYdGrZ66gas2HeCKdKxDG3LvecmKUEaFX7mtWW6z4RhYagWiFiHQpFGnS
1XN2B7+yXXAlLYEMs81GKX69oWoI6PJO5/zrahYBwQPo1mhY+eES/V88DLSuGsR8
XJ56FsCd0b1ZAE7bpzHOx/Q3tdJQcUrgtPcRYR4rJ+xSZ8fqbt1ar8XqI691YPgn
IqvukLNw7ZDP0JBvsCwoBtU5cUW2yubNn5sGOBtao4Vg/05d4P5J7FEb/sr+rGcx
bd1hUz3r41gbJvBT0W9loqGtYHAdGtylGoveGRAljnNpPhCUMjZydTWUKwtasUV/
2p/oqmXUeCqVsbTjOpVrSp1qmIXjwWygFREpm+pc6y8kQ2YcVrbANr/AxLeu2jxO
fOhpbNciZkQqnbsjbqF+AQXStv4gUGzrdvdm1avgqRJLhEOroFsQCaW8yPmvt5E/
q0Ry/qsHEyA25zsWJ8D8dWEhYHDvX3YSQETtoQ7Yt7rfsyASRhast7eDySa1GpCp
mdxm+FrI2EWOljlFSHrleP+kTdKKyGw/KtoUHKey+e+x0FbKVRo4To4KBWDjv897
zFvo3JiiMhO6NMkq6ZSb7Hl4yWnEiyLs1nferypVEtfFrTLdtREAE6CPD6U9ewi9
GVVpSaemXCrOAUEDS4vhsDMs9dDGTPqSrYw7/0JYro38rmZ4MYI28zQEesv86WVG
Tv1EQPylDN8Ji1jyF4ofV9550Mwj/Dkj63ktVNBCUq9Z21dYYUKFFQ33dJ1PrA6D
yxaUMmq23V4YSnXUriLUES55MPdzwUQfSYZjJia8EXufUQK7afYZQAmo5gV+N5v9
TSIzQDX1EO+31JuiuV+84cffDq2s0BGtEjgZUNhWBKgWGy2te/hk7rxfo+Z8L/M/
BZuRgyX6qEfQnXlRryC5PBpu+2pbcneC6CQCY5MQWjGRjOQVqPBhEwsQru6Q9reB
yNqRXJNG/hSEEy00NPT4xe0VGEFVEs+GfJ40n9OW+Daglfbo5/MP5THqfYbzlOyc
TB0aTrW0iSqJR+3W+mdpDSeyRzbDdLbUDVGtadmmetiORrqvfcG/gHQCl+27KwbU
y+lekNzBL9Xap8diM0oqscnNA2jxFGSs8fXTdNptOJbS+iZ7tvzEeTffrlKXfCy1
dvMnJr5EoC3CG2Vb9lC+clGhpnN++pfK9vY/e3nIXfYZXs2yEoeqUNC0aIMn7+g8
txsJ1IU8xtfkaBbHCQoEbpC/Cga8TZXpl+8+kd8PjvFDYEFfNTFkiG5dEmzA0QbL
lSaZ54MjKYPP0S81pfRXesjah2YUeW07Q90Yooj7BPl81RKq+xUb5/RMsPO8srTx
D9/FJVH8iOMHNGtQTobEWg5LxA3P2Z+6ECv8oazaiATIAmAKYgAJk6e6ntxPPNuh
fsbToVoxFNGZ9CSLyc0uMIcdf4a7ezRa+m0J5NUXfRhsTZtnoO+aaSznHTFHGjfb
G0czy2mBegY0c5Q2v+BW5oF9d1cP+illQ97YPySHM+A5yjIbGT38TPeKYxain+mV
A41z94eMOKQZEoSo30dniVLzuQPUu9BDDp0sIZKEIKo2w6rRsoe8DrQrEsxIZ3iK
LNIb2wH8+wJj6OXnN4dUo690Q/exjMc1o57ksEEguohiWZvY9/3fPnY1urDFtmKz
xH2XIHsdSfU1XKl7x3Lbffw77ioLaNSRKxIsBzpb1A9GG5IpP3/Sxs7tqQ5tGWZq
pb7B3PVXe7Wu6lel8bwKIeGUHW/XEzpxoepRe0vmIHCd4PRvibGW2kzjuYLYhSC4
7XRJA5tzLE0jTc50hBstjuELogmMikmSFAox2S5v1IR5G0yLWV1fpyhPSn9f5K0k
GtkwryRtJebUDgcgA/eFpeaCm8CV9FGQtxmC2IEHKFYzYMP9c0faad20iWoDR6DI
7Fhb6nHU8AcSHeBaY7RvnkAGpqBmgbMZ5W5B8tt7sCZ6RfU9ycRxOsDO7EMVK17B
JQNHbIKcQTX4Sl4LseCwTghAx8l9xYbsYRiL3di9HAYSRvo2Rip1IElXsfz4/2Wq
oxxO0cThFuQ2PUI1bzlSV4BgVL0gBBcYLDE9ZXyHkpijVtC4jAHXrj/kSIWXfo1N
n2jMveGG3h4KXIaVkcC7PsPreMr2eQmOvQ5Jtq+6pQf6XshbFAMZ+id23czuv72V
otujDswfe0Ye7BDoeh4FwNSRluuqn3TUKfI438VUpPr1tAXGl4VLB+Ca6wrCmUh1
trB+2H03vspuKwkb6ekyyfdjlVXrXnP7t7U8xD8W252u2JUXc/XWhmz6NWgKvmE3
vkve8AapBrpnirmV4wREqwGCJ0r6dpy9l6G5UWVaTtPcLSxkRT3O7Apv5pKH/naa
cUT4LWt88PXqPY9W46aXkeUyX+KHKaBJ5BjdAWgazFr7VK7al0Q0SR/Y5xApiJ0P
ay1DZHEydsdVuqM1Uw+bofaSQzrqgIDAa9blZ7HLRH8krTW5uPnPiz7N+BqvJfN6
R0nPYZTNON9nYuOZqeOntZavPml+qqfkG/fq/gPWXiCP6/wPW5riALUCJF3oGnUH
BMfa9N48f+omXA+5ZcYJT2I+x2mkYTcFwDG5eKznleqvSsP9RGQmdIDytRHKImE9
+OtKjIuBuLJxWfa4FPHVCHkVqqUUP1okL2qb31frTTMDEVAUtSboS3NRVR5ERIDG
btmQclDDYurEHCs8VA7AZ7DZEROSM127E41qAEp2uDUdd9558JlCsKJmnYJ++wVP
C7pEY6NCYjiUuq+AtO2tFEjGuckWKuAD4F+e7BjF8Klh1LUtFrDWwddr+4yKh0/9
yZ05eEqKbdINXWOqwFGZyNNOWudN43+mS1fE9Vt2MkLy0AIRH1BgEyzZo8IZUnB+
RPQSJyOOU86ZR6RAqCVa785JuAxNXKLQswTjulvbxuy6e+jZu/hN+DdN86fAe6BR
7g9vb1vlX4FBo1Syu5eNO0tE6QO4rvVyB8fV/IF2UxPqLQVdDfRnBlbWHjsunegN
MxAyOMRPGyT2XBFRVt38FROMptwJJYK36CSm42hGYWmYa9GDiQXMIEFeaKcifMvP
QVDbPy6DgCdUy4Gd/cfwKObUxRD4mukt57XSzOcxx3tsinfnokWQws1L+DnSG9mw
S5tmrFI7xJu2bsZjHmzzCIqFMftraHbC+xQBRXwWPjqe2HH/GbrZCybLmeg0niCi
SZ3d3xW0A/fGMtCNVMogvvGCLGgw2sPHWid49mFhCqihaLDspJ5gxO2GsO4whd5J
IxMX8HcWEJ4WbXy3I2hgbezto4eaUXoq0Ib7d7DA4s1mC6zjyhe6CpNBxaBGN6LN
gQU5z+IkvLOa6wZxdo3597FtTW3evlW7uwnbIbKB99cEvCTDMQ8qauRdnYXzjvrt
v6Wcc5DT0WsyjqCU39ci5y9JN7ph5BKZd0F/GePygAAKMO4JqK7vO6zaw60UPWWM
/x5mM7+5UkqWPuwmzfq+421g2xL01E5HkZeX1uppd5ooO+5VlLHqWp/BGuyMt5El
TrPQFSdDZnpzQ1f81zAIHUG9zuiB3ibymKHODa/yR7yOD2Np4k5pbCnA9r2wNXor
zgq8S4vCaI7l1CzjzI0vMwFnHGE3rr7AL/8MHk8PBSmmFDwuUeXOtaceffoi+l7V
P7rQaNZaDG77wPdN/2jqAIv3aLHR7VV8ROUR6AH9xjB6DC1AO6wpkgWAcZZt5RfO
e4+VfZiJdeG81nf0jBchgANV/ckra05UyjF1RvYhjKmU9V12s2EAB6398fzkS+bl
lEsrNhINfKSBCH8beRuVprxzNmAAspy7RBwRAktZlSwDv9lD/P+864Gp1IAon/8r
pWSWrwIWpNTtwXSYvncUgfnmC/SrMoXlzAGBtkPO8jugorPEFU57MWM3rMTccEDR
bXik6L/DE8/69XcNHOqxO5LIPmjEmgV+sU26omoZYNHJAcEprAP1A3bnG4rfzcBo
AppW3QUB7U9sXUO7AHhzb6Jh3XU/3z+mnEuLLGgB7/DKvX6q+TDend0+y4/1+yEl
zXKErZ4VrPwrecmaE/gJPkaE92af55w3MNUE65lZ9kF++faINf/ZwZncpVDltgSW
MluaLGvsQpaSDgEzFVfGTEeO+tGa1foDWhXggWVc1kLoOb+SZbDiNAj4FYp7lxwl
+8s3UgrDtMI0mOe0SEezVeVPnGUWEa9N23j2Vw1KyWeB+zylORqVW8vhg8t65U9C
3mnaRuMUBcH56h+FeFaJMLbcZdcG4E3efYctagAFpGuW3NGdtqT7g4Y99j298F9/
oOEdRzQNht9RhhHwBxliQyycFflXfncHJYVx9WsSfsbvLCXMjfgpBdB+aeTYbNPr
GFpDB0MNB8IsGSXxke56jOlk+RW761dMnHZixDiHtSRdVmftVYvQbv24VL2QUt5l
kWB51kS7Mdwnf69bKdJQor6Neea1zaUhLoNwa4x7Fr/ZZr4+MXwUbFHlX3rvtnxQ
hvUb5dkDEvQl7tllHX15zR2ZJiK8bXL5+4hRa0hBDOpnMCaS9ifE5WUJFw28Vw2e
eVZOmINRF15MwD/FP9totDB//hjZXsfZ72rTd7j6Bv/J+jdAOQME9lzT9vzCmQXO
Li53KEgHLF6Xkl+OPizxwgbkNPFXn9CUJINLChRvnaCGKeuK2lkwKi0hezs/kOp4
uoA254nt1LgIcZmnXdxr1n03HlcltprSxsM2qCNcq5srWRAR4qK5o6/zeWtWRO7d
smDPcwy71VseLDtb+fgZJvghZR4ro5uUC6gZHUezyi+Y3Ge4rHzTdAr/zO8BXv2Z
s32lrRonFcNebNk9tRAX+w17tFyFSo0KvIZ0fMIlGYeAVEBK/+TgCxfm5c9ABF17
zMecM2SaO7coCS23wFxtfUe9C0tBZFNSrck7XsSA0P0wQCeoCDf/e6W59mrZyrUl
XAraGD/ufR7nSBpRvHeGGB+zJHkUBHWku8IcgPKCHU7Pr5krYRY/V9gFtJF/qMum
JRb/dPDQSP2D/9D/LYpr3AgHeGQ5TFa9+zo7K50eEot8SjbTGa/5hJanl+e+9756
Br/wr+I6yQhiCO84DF7KrNOilm/M64YNo0zRluewtcILqtTwvRg9FEz09z3QKFzL
ZANV+mhpB3zfOaWvFLDKMrqtlAeai/5FtjnBC+oA7OIORqGDfbfxhjk9a7EuEnYV
XiHwElP1TGQxV7NBrhZEA9l5RlwL+ZmenPGDTBT59B+ufuuKL2BhUGRNzBoAm3h8
UOTms2MbK9rqGlBzKBzuRgPkHGdCeJ2HAIpX8ipBwFkqsGemiuRlnQb6uzDlhc9C
51i07vi+X0yjrg9tPqKY8PJQmaJmAlH8Iz+b6ZUyFSUFrSWX2EF8fAVry3bVFPc7
KI/7u1NF2OIjR1LqXbe6iiZW+zvaobEL5PsflFDQKmQ1yWhMJ154VgRm+RH44Tyd
+duzjemlU0Akw9N+3aNSoQB1QE8VIRsnFNGlt4jccWB0Dgk0GNJ3W/PybnDps5Ot
rAgKF+nEXA5K2j4ILanLzJlhH8NjNyg3vepxr3xGsQiLIOJOB2f9TwAeNRGXd+ML
lxtbt6QnuGx0vmspHcZP+dBoS9LMMb1I5ZF0GbcPLk3iy2PACq/mlTCxyeTByqIw
RWUTS/y3hf1SnjAUH8Xuom2VqjIUEKy2Vz6qE2HXBBmMY0Dgs/JX3ZXStre/n5LF
UQCwlLSD5jXe8uZEoxxoEkf7BxN/WJyNaskT6U+oWOozvvRA1Z/fPMYR1lALHGD9
vlOQvlZ3BZHeIsUXr8mYn8jvOC/WHzfeVpuAZjtin5K1AhIAqXo9KtxF2jXYGxCs
sO3+4319lPRbmMz0Tp49hpOqFX1lUE/ydzSHq6v+G4Qt1WPh+BKHb7XGSbiDWXk/
BMdRGciWgvhOhuVihEnoq+AlfZ88uhWBlniqpGULQHWHrldnYBkR9GBf3wCS6fnm
xKZBt3OJGlAxaNMC8KRcIQMAeOkGFxNQe+WrUBiAkj5Ru4eaZtWTGtxbZeYrIzrp
yVaA0Zc35a0SOBcdBmvpA2C0jk6c/CPiUQMKrH2uo47WW/Na+jxuAQ7w+PpstRqf
S8MV+FpTwhxWvF7qR6Gr7H3NKPkwMa3wRBfAVMPYB6cY/UbnLJ1Gy+wCPTPcBdLK
5U95i97HXr4rfjbJQON2PzNQb2/N8VdtjtElNW8vljlXQ+9Fe/AmnUGOq1kD1rQJ
xQFcguI6wnxNHWUXz0sHvPs/Fx1OrpmvXeTyGVPyCAlUcvSzQP+WuAsZJeuPHJko
6E6t9stQA0yx9GtPUDrihQ==
`protect END_PROTECTED
