`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vS5OnUTZ+kkHyaBcmVEGMAPGRwiepgP+7Rncy2XUiC1a0vs8RY+fskpcvh7LGMTt
At0bGHj/eXutRIODrvqEwy6xZ0YfIPD+8jWZ0UEeM/tZ6/fQkfYS6avpS/u5u+4b
75J4BiuQ8hun5f3t0RWFhorwqSV98DIe8U0J6gMMnt44SzHO4zymat+xZbD9gfF1
QXQ4WXEdnwcmnuYY1d/H0wFaBapdKRZ3TbHvH+Um3+cF/huA6aEEXPhMTkDpPx6W
m5RSQng62if+tnc0Ngx04yUcXhlg4kRU9u1/XDxmFRFfRCVFRANp3fZGOvzHw5iP
YDzCTSIqnfJgDIHAMJYyFDfk26xOx1Ct7VUCA++frgaHOanctlGkqEc+gxRdrwmd
LnrIHsaaci/ik77UyxiSdC7p8X0iAz9keRJ7tx1Rv55v8CIz7Rifbm4WLHkkYiFX
daKrG54jxkHi7udhCqpwH5DDK3cHXk1rldiBW5OKxhRU0ta1JzEA/SdlibbMuTXV
mERFRKGlgGK/YLVCUbMBigHbaL6ldXoFzM9C4Hqu1nXWGl8aFyZX7f9q5sukzXpG
XhaenyIGFFgy04jDs5csbhdoy1hNCasBrHfLsHCYJciH1L8xvZWR3rGxpG+rey5M
VlZCjgWO2KAwxzF13Gpx1ZwkPJFv8SD+bXb8uMWApdUR/tqamswWqdGJReZ/ScUF
`protect END_PROTECTED
