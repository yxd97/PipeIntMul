`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7UqpaWB2Vd61kyJ9JFYu7MK1iT27N68anlMOfpk6re5bzGb3iGWeK7jix4cmlety
ZOihGhfXJEvFRMSNB9GgWB6If/zKyqwS0w+nmHSg+Q2kMWVG7uO34QJeU0RmMoi6
Nv53uDfXrz8W+WmibkpXECLobPV+0s2q5BJK2P+CTrQPoKx/3iFBa3CHsdMh2Ji+
FavCvp65qM14RBMewtOj63lHiO/khnrnUJubadIta/6rKTKzlDZNbQTKf2f4x+j3
jKQHHUv5jMhQSI4Uqu7L6LMKQcq/5NdyKJwsZveWcbQtLM3z7wDURM1118645Tzt
M7sCbD+e2ycgJFptYAxDsrF1UdQqNHzSIFkj66MDcYpgoCswrsfbwVz+znqTe1Ye
ugU2KskVzf7tDHVSJTEHHw==
`protect END_PROTECTED
