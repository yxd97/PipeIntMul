`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
szs+G+VplM340yQhb/Q7O0cKBDv143H2RQ2vWVYuRQYwtCxH4lHHrzd+dt3HV5mO
1zsYlwhwgUkDO/2l4m1aVQ3fVrR+kytDdIYhvjmXecFtx53C0Sn2UNSZw8peskSs
wP9zVWGpdcpzUfFzRlGTuGjATi48vLSV8RKtDuzLQIoGbyCDg4HmadoIAM4oCLuW
8xSxfPRYXco0IxyUsnIXqzVFicJ5TXmz6LzEzMlhyFU8D7nD841k1LFVUgwWy1Lb
SNuq9dbViQFE2DQv3HqVTM10A1+iFI9brJoasheF5cY8VCUsH/X8gDKNz0DMV9ey
gX/mVDSMzrerF/KthFipahkx/4yr5VI40fmQziTWEXTRSrtf2I8+IpmJAAfe7dMk
vK24zVRX5R4Su5QDhKZq1Y8S4kNZ35vEGes10y6f2gH0PFDbUeWyBojTUyl2I1Vc
CPui8vFSm08tpICU3/3Hea6kdaKQOTeOSsXahscf8u8=
`protect END_PROTECTED
