`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0joPFevXqTYI3reShvQAoHMWf/yuZbAxQ9KPRj3kZ9qQtrSsSFawT2HzshdzrlBD
+ZRSJSMHqUSOIKW3zYE4ZIX3KdWUdgkjXW6fqv+mXQnJCKmk5osTenI/BK5Jkusy
VrQItDgGNRGkCtM/TJ2BtFoiGm8QDil5g1cqQ5rwECy6nK2DatT9kmlUfoN6Tkrk
LLlIWfEEqm7tZNIJbGmYD16SToa2Oz/DToVs8+zMtwaBvpzqIbtKxD0RrNbZ5Vd8
MTD83XTAo1FTNLIPfCpeIJWA6fZuz72OSGZ0Fih3LNo=
`protect END_PROTECTED
