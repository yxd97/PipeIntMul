`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lV6MB0dLF4iHg7eWdghvCJ1H9UPlZ7uH0ci1XUtxUQaLYFifVWMqyNdRAztcka4q
2QAgqS6SpLaRRq5SRbYPA5vzM/fbRu98UQINABViNK2u30JnwfMs0TQfuOZLHhNQ
1UGTq5VaD+nmGAhCUSdCsqqhPyLd7/tG7f89mhDVeJH5MqAAdwCBbhjFKVgP03kD
uHCgW+3isGoHSTFTxrRto3U93S73mSr1EU6rEFTtoq8XP2lVVqH+8s/3xU0TVg5y
w4ViWIECK/DFS7oDHsRTV4Qqt/nsJnwkn89sbTMSHsUhBuZLxUSSWaxBjk+/+Hva
jvtOw5SJ2zSGw6TuBiqgQcMVuD+2tMxreKws3zCSfa8sGda2wgvzYhd2OvtRFGlC
gZBZCQTOKfVvEgsiEShTx6J5NJKPPUgGySXXpYHeaKoOua63hptYtLg9h+R0qUGd
kNv9WfkS9+vdnmTugJUHCNRv5JzxYHkxlOqetvIkn8mdqb9nAm48utskWTtyz3uW
miFrDOWvBBTohJQ+5FoncYmEiFybXRGUnlsXdPwBKZKfugqz17NNr8ejuSrIMsc7
HfNQNLHiurZuj6AEDrco3VvbQEhKysBsT4VmNNGYFTVvX8cCSV24ok8vxSZngYVz
BTbd/tn9jYlpkW+aRpc5EQ6gr55mI4Sv86iE0UqoHYyrzDqmvUy5brcsetgyLfnZ
eLA6ABc/w6dm6LQTRWX0v+AWV+6wN550afLd5fFyKyRvAbxnRnquwpcTVkvpPIGH
K5XxUhwxxwgFlkifuq8vqHjKsE+p/f1SDxg70s7upgx3Dr9goTGfp7oULGfDCOyL
d43iQnHQodAxIoqRJYWZxwfbT9jYbhyxsyUzAjo4IGX4dH7svgPtQy2xckzkEDjN
cRtxWYnfuGPvGTEgEpTEm7z/ktC1xAEJiy203q/GQGLrF2cBLsv4kU/t2/pD7juU
hivb0xhwsdapYnEJss9Jz+SwftCr94QaaSwif1UJ2yUuZWXf0TcpzudlgCOglMQi
VjICvGlLrFoQdNju1CxKLae+pU+ef9IGgIdHTwWz0Jv5BMoH2sIJthCdaS7MNxhS
BZbcp+MCqG7WCHlJ4QAmA26DB8eRdYlWRFGAawSIRGzaEXM94A+r0RWZUfh6yBy+
`protect END_PROTECTED
