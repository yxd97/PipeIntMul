`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIsfo/xpPtNnf85AFc+GJa0VXZ7U8F4+zeUOUpd0L6OSywt4XmqsJdEaQYXrVcsw
Splv085k3YfGiWC/yQEC5Mp7QLN2Br39Gu2J17Fd/acxMCRn8+vzYmfGiYtY6isQ
ugyDBpbqJ2fOI9uNBvd/QCYd1dIhRicp2vTY13Bh5Mwx54O39KZJSldJlyFlVzqn
/MIh7dmIAIIumSDLiS/9WO96Q4+2f8W4kMPodd8j0NDyv20tU3wrCS2J+6N9jGv2
6a++tCYkgL2iq6SGlBOtOUFmG2nWGCBRpWVkAASKV8Qiogp9ug5s3qqz4Gh4Jxip
f03g7g22QjBB+Y24eoY/xTtvA30JWDePLAh4fegdYzHvY0mKtYT3J0CV+I/Fuk44
jLQ1keK7ZxoIhQRV2A+Uj9xXJL0sNvFT+Ar9Nfm4oAeCuVVyqD088osu8zn3yhR4
Dj1w/9Wr3slKpRxdj+nLswZ26QC6LnYtHk+6Iz3P475qCgINkJxWPNUDWFA4PE5v
`protect END_PROTECTED
