`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kCq874ISn+MK8Sdtcmhycv5HhSUUnrYNcluXuSWhQOg1Hb27gzsThe935Q2P3Rv/
vUQbI9GaclvyRdj9w90QXXBTjL7TVzC7kK+Gl4r7lRHTJyWCyquv3kQeMGkIkE2G
vGEmAzUPUbi3zfknlAske/J7yQgHLgOdmGEOfK1m+Za5v7AsBpHgFW54uWLEpY8K
ItogNyorxynJdkOCnF0rA4yn7TMUCrDREapBUMVxvZOq2FPfxBFYj7/AoLaWT/5J
AZiWVwUSz2n2XevZgbwjBgxxw6OJqkzqxI6RgSJ5Pkvp6Wr560jNib5jvK9RdnA1
zDfp8c8lXQ+D0GvEGGKYz82LMM69JmKD8q64h7rSoHHsJZT22iHf+7kKW+EPTrro
`protect END_PROTECTED
