`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEvtkRm4uvBF+TjHJRCQbQW7QIrmKNcLhcaJU41DeVXmlrWLGS57gXITPVzvRwxQ
BYE+uE4tyR9riQyBCAnsx5q6q3JrxH50h0ANoPX5PG4w8FBMRnEWlxBwNBfccUaR
CxuOyNa0Z4Q1NccvaePOzymKobdTk0zSVb3KIx0lZ3r62g8wKfYcVeud0uCfLMhe
spn7vKzKG/XjrLuaedVfeFCDccH4p0P0D1YrfeFIuXIR1q2t3dxto1/RlFV9s9Vp
NBW+dTu0psmhtEw1R+lvznFhSU2dmrbnohVQJ4mUsELq2h1VsSEMxCKCNL+xgULR
fh8AY9hPUjI8uggutaU21VUnoxXZeNDrY4buKFVlZOYyXVI6kHKIm9SkbvFvhMS/
SfKalG7UmxtRBdiXyFD3F4jCJlMJjbWm7fBl3+9i+Dri+4a41vYOckugDtZmUxAq
`protect END_PROTECTED
