`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oMIXNEV/d5cBHftOhdpDq0omXTW9IAnorjcSYq55ae0Zy7kiR8EvfX+q/+lSC/vf
w4wFLCgzKISxZ6sYpCT/fUMzQQDEsI1t+EhIZqevpbptWSdPNIZfQXqPWSJyHXgL
WYSvpg0qM4952FyOZ6SE4ZLUGvKPxfLmdVH1zemiCNCnLFIfe5KL4Pi9oKQnseN7
1gFptJTUny6NgFwOn+L+AKAP5qoVlIWP4z33n9OYroNpX4SRjOtZI/TysLVxtCYc
D8lrnVDsjsraV1B8IOW8uYP7tHyOIzzUL1QmuXtfU8UnwwN8OMIs4sAJYdeyKLf7
5eyi2zYZC9YMSHq3LuLumCfoaN42aziauSYiev+UqsmrfJ+49EP2RsF6cXigbMUr
m+GgsIObjSBhYLzw6ScYvw==
`protect END_PROTECTED
