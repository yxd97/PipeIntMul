`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGBGpsGiYQiEPUXGjIqI4vliqOtbYPfTDvsev4eLTCPy25cjb57mdtY/rvT9NfEW
Xrf9HyNscRTGfU2EPPU1MF2147Rc3lwMsZaeyte0re8wnsB1O+KHR75XX1lQ1FIW
bLyXIkqq+vudKIrluq7s9uW8NNOO21uD33ud6ueINcMuP8DHXWIYFfWfyXCGCWXq
OJ/ba75xWforgbWLsgOhos22l7Z5ci40+czDmgLokDxrNi9DVJeYQrLIv9RJbqsn
c/3GwzQRKpfTmWLnWtMkgL4mppoGfuaTxBJMw6UiQtF5hS7++Vxd+XfM8uDBAAYM
6S1Fhb+U5ukm/uQtdAJ5uST7hkvrpsOjEPJkZ6dRjBV5SIMs/zOkbUAAaAOJf4Zp
lI6OIsPvjUdVjcnrqTwol+0u3tKWvrlPcxcY0/SWsANpnsdRhoSXgo9Fba2Ck2GI
ybkeK0VOtoACOyFWk92kKH2EWnazH8dKEOQufAvHRjWXr90cMNtmpw7iD2iqUK1l
WFI18T/68D6DLrcWtaKWvRQtjxuFGewvjIc1f8LK9EME3E72UrL0N5BkdzEL12jj
C5B0txgV5x5EOLQ8I+Xe5hkeJeVMpVJPHgT+vkBYfg/AWYlhRz65GVcc4v/PJCUp
0M+//YZcz2ODLlsjo6upkA2At1lrVhkEPEtNeQ/Fhe6fmgzpdDh7zybAoCoLqaEI
jAhHgCdMfshUvaNdZZEVYvxOb9sGt1XLAT/ozDPq2BuWMSbfYIhy4IpU8mffuNCk
AKeKwOCVQr8je1hr4IdyxHAtnN12cVqZxHilkSSjYQkhfKoBOTshmaq2Mv04Mj2j
4ybHAacjdgvHluyK1CkNGYmOlGotAm9fyBvPGhRzM8pF2gNiGjfMdyh8lU3lEQBf
RouG2EprufbAz3hjbj4BrRNVLmqlwe4ZI4sDo/rVjOHo7mn6q7AGAGMIrhdb0ybC
eBMbvv+vobo/Gj/ncENYT3zJOu7fWZ8RGy065eV6zcQGrkJN9W3zeV9Rr4y9uhcp
QCJtHFRgzXOP1IgTEZOp9tj/4EzKpn7QqF+ElRC9najdYXVPqONIK49JlOMGur+F
1FjYKHzoKvt0ZUpt2LOxtTPod3+XT1s1zbz5yNQsHTTWxtpKph2BSN0izZOIuavP
zRPCMLiJZ9QuieM5PfJpLjW7lQHg21ApTDwrt0RCJaArvULuoSDPwaV+5jA9ne56
+1SaLtg7E0U0j4bnIAJzTYvo8B8RVwmANElkwUWJnxC38KyNFSXAmZ3l6rWWILm2
wtLDbO3KNK08c5q+HQlznSo9TCOUiIgv3hdCGR30kP0+nssuQUDTiS7e0CDfl01x
6TqHOlTnKvylef0QHT0aUjivAE7mQtf9GuMBqTyYYoKF4Nutefg0LRIVkTNhTWlY
4swnqJeLqKe80+5dHJgvSuQ5qFBsTbxSO+GCS9XBL+4yN8vjjsJlP2Z77itV94An
FdanT40VjGvFADvMs5vyYr/xaLV8VBKvD56GMBZwLVgmAMGTI+TayrwYTEv6IzVQ
1Rgnf6p0o5EIdwdJ76HBl2yTSP0hbYfMS5Fb+ec01JoCOFfCx0VW+yZ+rH7iDw8M
1uf4AEdvqUaXlv3DJifHLSTkf85FhGs6TAcZ0WnT0sdILxKMRjNQ1+k7gGuIG7BM
KD2V8LQ4Mk8Jaieg2UxtvurNueX3bMRfBtZ5lwVEfywORPRFT7dvPqibkDnMcCyp
lFEfOt+FuTdAm54SrzfykOrXzSkkm/k1QFQ22f4RG+1dPUtK7VSctJyIpeUIYkET
21XUlpmildTB2hhIVB9swLVRmrzlMwHH2ZLSmAEH5ScWq5P7fpwTp7uhhqbxmdfd
xBjxyWjGaojF6aHCkYd+QhXZdrhkUs78NFNKojH7YYaPLlZ1EAloAFq/OckYjPAz
ek0PCPRpRZl1P48HVcZrIVF/kegWkynxGktslJ3AXZxHMQDWsfzjZyW0OzQfRK/g
k5hvsDq6yr+ZwVjZSwphwLLH/2V2+RzhLhc1zc5J2930/AZ9YMKvSZ6HEo+YixX+
VxyFMbx3fOk3hWunSCff8VVfimAxxmOwi2Z68xXP4xgzbG5LPbyU/nf+4HUMMmce
hI1VnKbZ4+h3khPRAfnXHtfncIqsjdofuqolep1X+t0y3v51pIbPxbj4I0x/QkHh
8LW6I40fTOZmGD41Poyy+ktK6u2x2zxMICnX9vQ1yprSGXy/dRw8UFAn1z9PqBkB
Khqo5soCJbLrQ1HB+KPa+Bv9d6ovJo3kqC+gu7UOcrAWkZ5Pi00ejxjF0KwKTEC9
zzNuQ8/5PQK5NFL6eyfXAq6nVX5Mff80FPyZSDVygjp+zqz0RYqOxvCsi7/c9ttN
ur0B+/jhvTQJzNHGnCeVE5avQTk67Mq13CNQCs9asG6Z0t+1pHJFSeQu+xBnvmYu
T8XjnVjGdMaxVuHgqthBjOdW0Y0wBMxoGogrKBxNO1Pu62cKgT4Kyfsfb/171+ov
jzZxkqMKj6Rf6IQnFrC6tjCazqpXJUqJlUmPVFND/bBaR3TQ5mf9j5+dU9E5yg75
HEt25avyVFZdfDSDwPdH1OEm/iIBrlKMWWYRL0KabMKxqY4YYMss6JW/f2V/zgt4
yim4znl9SKtCp96x5RsGufajMxhNsGr0hFyJFIwWdGWj9B5lBRswhgJriRRmL024
J7KOY6qNg6Ceg3xhELzMBcuWe//60TuvkheF3FzROQLw8GOezKR7chti51g3dV+q
ZdXEIdSAgogbuMpPQ3RCkXVSbfVXQwZFuL4HrC1VKUakarDVsYYlzaE0grh6ae+g
5p16l3DpWitH7KKHUDPr9HshMkny0j4KxDeFwB8A1rKkTUfI7o7YfqGc/acXPbsO
FBrvsuXaaibvRAb7uKP+78jasLyTabf60vAbgQNBKZX3gebECAMKVrDCWJaC7cNI
`protect END_PROTECTED
