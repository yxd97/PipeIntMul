`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30R2Ktm9jFYho/6N+iPoa1drTn0f/k85cTBeKaNjZriXNsiis3OFye9rIeGR6p42
63wccy4ob9jL69fItv+7rOjJoHGUwqw+R97HrRmrk8Voz36nl5VkbQ/kyeJ7COl0
WFSPcvzRr6pQ8tFnbWQoho0X+tmVz1HUUPYSAcG9TQO/859lorpqdRfLW5UPojja
yXcRlKdnAW111rTdbRg3pIYYLs2Ew2NxOivG8D+oBRpwEn/LZrIjRQdiWFWKjkuG
YzhrmBXVYU+WS6KcPp+cag3ulB6dBGPRxVPXDicza9UrYJHFMifso22W8re9nDUf
Lo+0qUWKtpN80k74ixYnJBjZS2OzhVQJy26e/ZWClqQMfQpDl96t5Nh2po44qD4q
VLNxJ5jIdJwJ45J+TOtEVQHhmUGEHyfw2/3NtuU09jCOi3rqAv6/qaVgg9BPT1aK
`protect END_PROTECTED
