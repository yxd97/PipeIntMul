`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QiLSvZDTDrATdfkhMUPzQ4ZQVvcl0RQ8d3PEoXRJ9OAa7Kj76irD7MPYXmn//Yyt
3L4sgz9EynbDCkz0pObL0g4L0hwecMeZxhuzqlgcGRGItrWTkS9kKOAD2ySU7EUE
o2uNQed6Z39jCroqgheo/VsTTZEuApDNSZmmUfVtfjMAw3/bhDzYnXPfD/Bs+HmC
unXw7tOK9j4ltfWctYxrisASbIfuZA53e7rLj+cQW9OLT4rWuO9ig1e2/+1vcnZr
fggr+TxL53ohj2ruCUU0O2WXhI8OKZD2apgtT6h3NMCxorHZcVv/jyilmCIIq5vm
rOW4pVCB0aZDt7o7cJesBVBZpsagxRWpKht4+KqIsSLQ78Nb0mVqh/g4tXUaKMMj
FLp5H7ZafjdNTIP8LQvq3w==
`protect END_PROTECTED
