`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zFc3Q6sWsum+IoxypIX/CHrJVd0N86z78QAYCN7CWFNnWDkVhzTEjnrZVITKhOvK
RehTia5w8vcpfOtAudGmg3dezmkUuMuq/Tlle688eXKjH2rGW+YaIahnnRBfdhhS
+13WrtlX2fpcqZ+djiitXc4JxkW9uw4JDSyIgpgVAKzq796Pa1XOp1akZ0bwL6Oh
wiE36IhxwOZAhdumM6X3IU6DYQFaDkYuUF+Y7T0iR8aDj6NqDyk3mPrcuVyfge6H
rns9WysyH7s80jqiK0GjPTNUyoy4BYrWZ9jL+wki94Rqzze4XiLsLeo5ix+M4V9u
ES3/AtwqREkHyMQ6r2xGtPhZufahfKMH34g8R4w7ze7xf+xkP8j7p5RabJavOV0w
nvogKGkQ4weialZ+nejEvRSSBDFPYLyT6WZhgXHodn0=
`protect END_PROTECTED
