`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cT3p4tRHe90P6+Fwur76UYGITvfGlwUZwxDAasaxwJGEZN3mq9LtxAoNQq0nJu2n
ciTOmN4478BReNkVyXoJ6VsRfcHe9Rdak2sBQofcoNWN7UYSwcwGPoP6pM7r+SZ3
eQZOX/pEKzAEGac+RXxkuahVXWE9brsGFlh9225xSi/QgJr8E0ASA59t75D235w3
fUOBDY7RuWHiTyFdPI3Ocy4HluEvZKwcbws2kd39tm56EGuYUhUhbOR77kqOU48s
U0nR4+hJi7492/KLSN6JmpP55wzJw8Nst+shmcwhTk+6mohNuKHnStDhrcku2NSz
pVGon512HEc5hBSfDmWb5NcdBepaW0rxcqPdpMUG51RqO0jspUGoPppNQd85vOEH
38CeLmC25AZe8YUWAYLsP7ZdNNbiO+grsQ9aciK7ZHbFnT1bTg4DEXDWiTKJpY+D
NkLGGlz2gaoeOB8axpOP62PdRO9ClGnIthS/D5CN7Pq2zKRS4NpSstDy35arTF76
rcsw9K9csBx49ItoVCJwwE9MDAEK/gQP0DQOwVCNafLreUMIvG1q5l64d75cxQvT
/T4o7v761M4ZX/IF7R/zlVbNMsQg10Mf8TuawkWDAj1eOpoehpzicj20d6zxB3Hq
9qgvDNlR/z0VeNjQhpH2F7WmumjXHycO7kpLidcecxhst+SDLn2KdJD18QcrnFAc
oT6y6nue/NR/b9lRRXh8Q/z/y8WNaSB+CqfYaLPhOYsVXTV7xAyi0Q9pXkFYmqRA
nFMKX9NWzdvzLdan9hLAtjzhO5sEhNACBI7jpxl6kSZIvGJ+YnTpRaxWS18sMbwi
d/wXa/SA/luP0EZY4CLUpOnqyMmRI8ILF4i2zc8mRwGIvHKdwCpMqUnWI1vKXOZm
SS9INNlxKNxZRb1tg2RzdFcFgvc58TwhBYfUnjvPOr36BftELUkqk/aWCgqrFm8N
NIvH8hmb+ZlxmVzKrI9vuzAsFIBrfoLWMxJ8iRMHsMnJYivrPc9XAr9AOjn0Yyfd
jLZoq8yCnSCbhMsN9gjWH7SqRvS7ocHNYbzVI1RWdxvix2lzvti6RzQPwX5FcfVg
ADKIUne/SfMGUJ3YVkGboyz0npPO3TT9lAM0IDluXr/2K/7kWK2cnWegf6Jq759i
xKLK6T9Y/KNYgQO0wybnbk3MWYqIfSftV3fbTsRG04GUpbVWCRp+TI1WiZEoX5zK
Ys8+mJpITtLMM8a61LOpBuXhXGYN7IsYJzktYpZF8K5ikCpgi8AF2Z2HJZ7PTKGH
+C4clNvvuBIBEbxwjvqhcH4hGrSrfXBuT6Z9Pe54Ays1KNOS0v1T0IvEATN/naG7
9ImW3hV+HcITIUF724f6pyuzv31cPHnLdRd3japl2TMVYuatZAusul7Y6dJzu/YZ
WS6c+XPe3oE6dMUiQoO+OhVOJ8iCs9nOsh/M5swFVCE6qh+pjiO76qXBxqDK7yB0
D8tZqiGtkHgARdSiSSC2if2gi8MiTqEjg5wmjgWWm+pz0Je/tqneDBrw2i9mQ6ME
7IeHrHhq9jpMeTgtjNXkZ1CfMahmKRTXrk4KStdVYQV+OjVo3JhKoiy8WHurccla
zi7Vw1/LMXuc88b2cYmwO8mNHxrkNltenEtmbLmn1asRJJaaLQIEcl55Md9t2V4q
xe/fbxIKg5BOR998x2GonrdAPBp+8SjXTOz74lfxrMbYkBO/kTYe81RpY+PfimRh
xDp4Vd0U/xFwL3khj+f7NiJ0wU/iC7pl4kwoJceCntPIxuZPVVrIhNlkHhQuYiuH
v274hja9Cxx4eETSBkpaIGBaeVZHwjPpUvEoyzTSKHtgU7RvWy9CV6RTmhRC08in
6Y59cwTXeWwhFfoWdFakUb5R7rIbzXpkdouCyPgtVZXBpzWFPdsa0rGGOFVd3Wj4
qN1i623mbp/L7jpDN2k7EcW8dYu8kkzPMbgJT5hyAXNigDDLb8rpCd8PZ+/o0E+C
I8P0kyXcEVwgKvZMEMwoDgv1snaB4q/dLQ7CvUTrd+qB6LuWrNooV+ntUjno9ral
0X5UacckBj0pYX7BpKfYvE4330/hxTbBhy4hmgnc2daGLwvkTzGyO8IYj2eRXUji
Yct8QCu0UkJ4mF13J90vDI66gO1oqPkE/Uiou7U1iWnDpe12iwmya7Pa3kVj9vCx
PZ5cvVo/02zIGBqUKr8s9gQ1bcrlYFTz0oFKw83KivRkkym3rXK117Pf11b3MohM
cRBoiRhqk0DE8pJfiewWghE9khfJNejQZRGhEEpnQA7SYe6CdtwS8iAs/DwE7Et8
yOpjxkDXeN1XGY+2L+LP3CijCAGYI2OCgm8pJctAlxqlyBN2HGXeYbHEYkXnxphA
i5DloAlCaH1yuqKOzdlbmJWdNL6JYQl7CYN3J1og06r+TWNTKY+SDN3DBvGYFmok
K2J5F1ylEmI2Mh6sXOs+I2wSbYS+PTX9tnwomDAerQecX9oXAN/AmnK3WhFRNcnA
khobGJDSdo9V1W1ozsVJPgbaltaqTMwP+Vt9KvyKlcLEjiLvET83luW/Gv+mkmTw
gvjxbHzC0Hy5cR8t0Fydd2QUZfxDleFkCFa/NCNdWPjJOa/1At2pWwH5nJSp/xML
ZAr9YAs7yDQHDskgGaTNl8ZUkva5uB4Dw2iZaFuKCKKRjKVtPz4onCAPYGobMDQ9
THz9s0lEkD9j+5IgqqN5WeDvqOYFptrxthL/xX/37F2rRTtKM4I3Sacb+xfpjVli
Z6uehsyASoKtotVk/ikJi7i7Vxt3PyukCVdc+B52DK/0Xsqu21yg171WQGavv9OS
SicW28KqsnfEJOFY61bkpP/5prLgNS/mGRrR15n+oP+D/q+JOI8VneAXNT1jXPkv
joDi6GMLjgMVr48X2k+f+HVgZIAsYYu+UCFm2pJfllFFj70tcj0M4SD7GxzZBDVC
VzXbQ+Ha3dVftzUt3SI3R/KFDBSbycgSCV3fXTMwuZkTpLk2hw5FQG4KFIGnlnTv
XpO2W77QD+82fvg2ybN0QstL9fyv4nZO/dA3ppocIiA4AmMjtVBoR3upQC8rPdY3
CtGG4KDlt55IyIGY16sVc0I299lf0/U/GZdxxiVDkaryeeJukjmxfFkCw4OCMZaC
lX0XLvnj46sVDdxXqPzsGi3V5XGoO8mYeFMFhVQYZ26f/za6M779CdWqzYMUpzSO
HrW65Pjd0j4NBojp+BxTrW1kBSqignDC0NXIQ4rm6PPv0/8ZbHjeEDleiaLibMAs
iiyhvdbb2VbrlEM2my2UYDimmLX71Nwg1KLQ4qkrKJ9nen57WHgddn5jiGFHEzU5
BJ1vzdx4gt48JsaztEw9G9rfElKiBBA2Lwvy7s6XwkHeROAdvs5sMIyJO1WzJrsO
XEvQ56yP9IOexklv1pd7bZdsDa3GZhvrqDhutluuaI2ufyRB287H1ktzQcVyf/1J
tATbD977jRyf+B+fegYdZiwYzzIlZb8scwoYImSgucAEaSWJci/7z9E/v97lm9l/
hsEutJ00xxZ0YZw77A9xn2P/3Ef5VjJ3nCllAIh8uT19mQ61K9D/uer32QnwKl2e
0GFarwkG7BJO8KrqJjvvhRvZ+9TdhktN50y1qKi/113N/mFI3K5dNL96zwekZ90/
e2vTmxT2uoKU0io+o2AakHB4DNvesNwdaBowdg6mJ2dTiC5lWQ1p0aDhTSXTKjq7
rpw3fG5N5GKqmSwCHMb4DvO0jqEHuBMCnjKWWZBNdYrUudpCYVndBk+JG5eoer5Z
fwXlRzx0X9UfpejIIc1aBgG1g46DWX0hYG2+fROmlYWFaaa5hinHW9n2nBJgLU7e
CG6T2U5+pSOn0SS+7VGz2iAA8v6pC6LCx2529fd8rdqZc8Avfx0eJHRV4RyiScgo
T6XyFvrFpzbyc995vObDLBgi+omCX1Q/2DENpwPaGT+D34ExIAPa4nGnoqfvi4Jd
fjIsMRkmlO4BS4UVRTu4isqf9TzyFGErJntlEqse86oYQl2FjRUFC5kWhgC+Yj43
JHjKE+2bQSWmSEhjIDAH4MDI04XaSEMIP6Ofc+zTxRGnd6foNdOi36QY0lfMEHLA
NJM7/Xl3MCvlf0dDK+9m5KH0XTtuLTROckOznUqycuqF5MlNucRrfEMV8yNaH/uU
PSoZtx1oERHTrEtPqPCj8gBy7T+h3K7+SLJlHceVbz9vkKQcjgNsemYqJA5mY5XF
H2ujkCSQNLfUL0RlCmwGOK/43EEJ6HBCwsFPFLwHCWYY+t6JIGNCAssgDBGneD/f
dGZYd0KvFajKX4uJG6QuebQK2VKpL+NKn0FwtCuyULgid9AXf6H0IjnQu3fWN2dP
kxpXucHpGJyfjv9/iputDYsabtAoR6dAbrhOZ9SxveTL8/UZRzFlTy1iFM87829H
5/6UQtDIPYgAngPujkl3PIAAN99++mBsMg60W1LM3AIsOCzOyOQvNgvMukJXaxrw
bEZNahUOoeR+uFURbQeG6ok8inizvZlyh+YQwzmF6Ew/mCniWV8h523nR8P8ig9o
Oi3y1JJPutQSLm2R/q4w0RDcWeBFOWMgDcXTsvPg6OReea1P00xOUIl40r8jmJNh
FnuwASiJoX8dzJhuNAcA5cKdzEo35pn6PHI7lslZn/0XH8k8GcxxdRXRqJqLgIwn
sl4XfvjrGgeh0OSj1lN0+vbB2zzTPX3qwdxDs/yaF31tx4mCrGPAg4aOY2ySPrmY
cuxXA7rMSCjDXhjxlXzZ4InVqZfblye8U4iVGAHRMLJ/0BUrdzjkBb3E6ltPzag1
EBTgDVpmC0h1YP1JKW/A7vvCS7ctXTxhZCKyCvxO3zmzbUkSgDhKqilN439y16Pu
0nAU5EBbMtb7emXl9TmDPaPzH5O6xyEduqQ+24Acd5Npp2Qdb7Z4C9P6W9jaApN5
bt5yG+PBJp5DTo3e5FvUtJLCCYcYxwmh1eh2pRMvnp3iXnIEcTl0Cy17SpVloF9p
y3KMEqPszq1lotQzac5yOcY78QKevyu10geby4iy9hX2ATRn1jsupp4DhiuaNXBC
TkGKKdQkfdlNmtl2JOVK7GUTQ0OjSm4lWz01Y/hXRjpP5VN1mEnOlK3mo3RLGeSp
1ezjgsl2oJ7u5WWwEy98TVaAIO576VltZJNps1kQxHxGNksCJ30eokv19GNwVRLX
d3U/RqYNMMyVZEj/XlDeIfXeQqmu1Q8kI4MOe76/SXHsoxe7JMJLt9W/75msOw0e
j20PqTAn6mZPcV+S8Itn7JpDsHMudgc0Bx5OIDTetarKXPOx+JTN04nTuMsKx3xv
pHgVEi/s3aMESvF+OnE0p9aaiCs6KrBgmiusciEB9w4BjIfmncoYOrtWmT8vaZqO
eHfj0qxQPdEYp6zhubJlPX0B4p0ki4wavFU85YMQ49lJ1O63qBSuZfWfmeD0LvPd
jzvBoU4QCtTVAqGFlWi30y8p1YHHxWxJSUqU/ZFRvB8uhdoYd1iaeVOyGl+RClQo
itQ1DX1MV8xW1W74EOdwwt1l8hLEKfeydsRFXz6ZvlMjpw2cNHemFuno72KpCtgy
qqahJ/JsfCL5WdklyW5gBdxwJd0SEGS+/RcNcQBt1IVsKod/OTPTqzLndSlKFSVb
nxl7kuMeybkmAugU+uLltAIAqWKtlym2ox2KbWS/S7K/HQmx9XpA3UpSJFvNNIyR
2WQOdvmEPibs4aDg1V0trbqliwaLnSjzCpjBK1S50I1E0HludRw4VXKKRfjn9OCG
R+XIqiDSgwfGR9xsbJKKBgTrZoKw5quMv7JGC2jevRN8kitmIXoEwvBOpAKE6WGW
8W8Q3PNV8IhEvCrl4FDtZpK5ei6rA/Og020pKz1E2+zJhUJDCiPwpG5bsI5xpbQR
2uYdGILS+YREpX+dFI1NxnC3MiUtLevrrlv/KppTgXpA67eKYOsYeVJ/OkH9SCgj
TqdbVtSPL3OCsxRsdqJ3Bc+2AOoY+Lc8CW+4QNBtB4LOsnyFmQBwh85otyu122ka
PUvlu/Qt7BLEkihmMQGbRGMOxEgFCUOLd7fbTWeZQMI+M0NjgVzoyh+PfBzLUcmN
6lmgs0/K4ldq8WER14N+VIDFYR0R9iGHVSO9awobBsnvVZ4jJRoINdZsX/rFTODB
xrzfbAfwO1M9Ho1QLc1tQJu7U0AwvRzEoCrW/sihn33izXiMG1XhsOwaNe9HKvwR
m3h/rYluaWfS7pO8UvUvhD0+HYf7GbTwziFIt/xZigoAxtPtXxF3rB5kEXS6Aht0
PadmRapa38xcmDuQ720Ikxqx1RSkkjrMCO5723RLt0zgrZvbl1sfcDz9kXr2yWSm
0/AJEWjLmBYClkTtczr9Wv6xk9dRCv+G8e4bqlPMDT0Zt43xqwZSa55vJta+TAr3
ippvOILL7h81C22V6RAGAGXBtgt96b7GOlYjKoXytaqCmZIef6tFhvcmVLdMjZW7
Q6DM/QfOPiotxSAQtBIUt3WsZElH4vTMt7PE2vYdJHj2NpkwMO+1Wzi9u05CuY+o
D9R6lEA2TPveQJSFJLtXN8lym1Wj0jXiKuLczEh2UZcz8fYGynevkk+LRhFcsMEk
vAG43k5gQUUBK4PGW0yhDXCp45BJ+EhH7DtT2beKsAPQ3isO5hcuHI1kBIFdOWet
PKEaYXJ4reeX5C9xCB2C3BPPSpYZGrX+wML8gblxms6bBY4eQVad1RDu3Tbal0AN
aAbpvs2yC6G9MWiMtJ+zW+dGqun/S3SMOIr0a4s7s3yYNCRr8hRzqXHRNStsA3TN
Yey4HL0+LrKrL1Iu0oFPxLWWNUWPlA18gEiSbLnn6sSa+H3jJ5m28ABWJjr6vYxB
vO3IB1L7fghVe6kWHed+ciH173fRirrpABquN9BvmUACC6WxYPaDRfg1NuDZb1ET
p3+bBzvetzlHbV/EoNtRBbUKekSYwrg64bzhFDIJGSmt27dwDbTbMaZ+UVoRPdwy
9OPySx2AoVlE6UULQR4yl17iqb90TuyRtbe17TOAhCbG7EGcMXfpgbnpU0h9o+4X
fLMeFFLXgjGGPAWc4kO6O1g8JQ5VyOUVV+Pri9foM3szGiKLyXRNYXw561rqnP48
DYRiV/neDNheCHfHVTT9pq/EbHIpK19zxknQTt7QjpyAFhnuWWf6gYfVB7rVW+2J
dksZT6EnnjjLBMhw4eej+5sxj1bH8b/2m+yDp/KU68dSUEigpFPbltaivvser8Qf
b5AOG8Mct8+iijfixlsFleks86BfgoCmRGCll6huGLlC58n2v5DkRk4VOiW9lrYw
AzDDFSunPOE3F2DhaifGag31RC+rxxX0D1xCPCEjEFA9m99da5PrtKAhAQsPQYrG
SiSF4TFM6tIJb79pGwoLiVVRLM4ZEqZhq5rp5BDT1VGMXAimQjiDCmx3EhGpzsie
/jQAgDuvZF1rW9HEk79EihId5mVcaCwRH/G4aGJjQaIqpdNB6aKfV9qD0nrejbO4
`protect END_PROTECTED
