`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixRxjf907gPSuVl93HDJaw6yqMrA44qUaXI2Hzx3NmHDhCdtk77Dl5zx+spf6JFC
AurByt/CQmZbpCT3EMX/KmMk/a+KI+qcfRcFr3miMbOFYkHbI9ntvFCYpAZTeM1B
hLJu/KCixBf2EFUKvu0Hvt2f3nvM8I4wdBkmJTERzybjKAnFLc9D6ONLolFTgymO
GxSXeKiv4FmjGmXiNRCV3TmwTQB4tD7uV0FiLxxh9ARhUpjuEy9ClchWGykS+VQk
MzCQaNmu+VNkKAccixhqTGWPAv90oHZA29mYm9ocogUVDquWknFxpH3K59HnSnob
U6LtKnuKR66CclAicjoVeiF/UBzgauMjZumQZuhQ+uOh5PKJ+uyVovKdTAy0QT/N
yxcR/bfDqqWxKTTyFx0i6gAbwRqP34EBb1czosjHGR1voNmVOrPzUR0Sino4P6/a
`protect END_PROTECTED
