`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiW3yzYN7gMr1dD3sgJfVfW/MuC/n4iHbtLcVtTfht9eEBxJ2wZa9r879PD7uKpE
44tTG0uCPnslbqg8AU/Wf3Nfa9jlrY0uZKP6w9noRZXs079+ZiV8l5YFVgZSmp0m
qGj1J+H+BAbtjB1Q/s5FbYwFhiM8Me6bW1CvIN0jrL3QXMcFGLmfXF7c0YHfZLoz
GOMRC9UFJ+9YuzebFcSjiQd+uF53rKQib3eXTyMnQlsclNLWTUNnID8NxAS0AraI
wN8yMmRa2BCnnXmltzaaMVwMqyKRw67n0isi8F5vV/w5/WVm0zP130wqiyHbyjlt
pYdsplpULXB9Iz9y59bfG7PPxKVJQPGFB4PTSp8PUgq/PjsVJUOnYx5vu6RBGHhl
FZxZF2b5Il0Luz4TCXtP/p/tEqF5kPcdWkTEMaq/mOot3OE839Oh5gkp8mypxP94
7DqmDYCh9H3hnyAps+3BumL2ZK3DIVvTHJm4oD2bIihB1I8M7Bospu3frqyQno/X
WklenmE846CH3tHdUkNOn+oT3jWeUWHjGdMbfRDqQRvPeh/QunjTHBLRGXQSicK+
qQbvPEx9jUUJKWlin31BWQbRmO95zNvdcjgpb2jP+WC8kV8G32itBTJs8wAugFfB
eIUuBoZ5cfJ311Avw1V0N27rpnCWf8FT23+pNYSS6oZ43CSF4dhB5bi17xiblpRj
f1YCHO2EHWrsBNH+a5arO9Um3+nwXXgKV8pvUqRZJP0XAxKGjMN1o2YyZ+X7QV9O
7tGm+WYwEP6JR9VuaSfehRPh4kp4CaHaf3sNrSUgx3DeoRoO8WMAd68HrFmQnWn6
VdGb3j2eht8Ai9MsPVlDkVVvR7mcb2lAbX4fsj3sQvqkz5J2o6l7QWFphjA4P43m
3+owbc5EQBccrh69AS3/Cw==
`protect END_PROTECTED
