`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hFOXqq/D4fy5BOTKsa2KU+2K/oLlueaDBJcWiajXhmxyvyd5JKgdh27YzeAcvvY0
FiHc3kvkzkjsGuF7zppeod35/H/4N13nPDD9a0j04BTi4GY4nwnzinAkuJC7cqPq
/njptRMR7HqcjcUxWjGvCNLAIG3N5uZt/Ilwp2APdZ2E1SxWBG1SqC+Y5h9yDiFj
gUIq8JzfUCnjPtU98SAsKo7oCKYsOUDSB/Z5zcaA4Sf/kj1H5HfyfrqS3CwBDdYq
JWoRW7ouJQocTz1mWIKoKlt0Dy3Ke1St33h81cVlktxFHUkYT+amFPAQKM2USJHV
3YLv3vZXU04uqiT8NOtwspIZ/5QBsMYmTZjUAZv6/2kNlv06IQtTGChx39QSWoVQ
B1h0J8GV8kcTD+jiwgWIF7Msz8r1sdDhKOjRBSoEGcVZJCAH9+DWOz1PbKzLB2P6
rbdgfzt8PL9yJnNO35cd0Jp9YC+0iepbgOOEnHsqHXXtyAqQ1qTv90SZCzxhB+KT
8fS8VG4NMjeureaIa2Ue3Rd2CJKJXHcp7BHmMaoO1lMLlAWhfg4trizBbK//pA4W
ntgV7WWoto0iJpZi5wG5T6s4oXzT0jxnftmyCjugCmXZ2HqRACAJJo8cDwe46Mvb
4EiCwEGvy94Y6Y23nPm5xR590hlwLKpYfivtG03TNq25EkJRQLEmIvMbkpk9x7bo
`protect END_PROTECTED
