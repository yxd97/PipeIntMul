`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmPionqapp4Mbwoq7+GUmHDZH3B3WCyYXKQYrlOrSKo1Bg5ChnUSpOJMQmnANQ0K
jW9JG+lMBnC8zoEvZ0MLwFYp5ztaCsiDCqJbkg1GjBvqp1OvpGycfCziNhzGDkL8
6RkUi3fCUzvPfADKnZ9veJ4fq1C9Hk22t1/9mwjIEHlLp9CxtyxfL4/uUZrzJ8Vb
i6E//YxR56nERmQlG4hUDdFOYqalVpTdpqj95WNRO8peo0DImievDeZJPEuZ+yfa
9cpQicH8Y6MR1rdBydoylqafXg0IkE2sqYPCN89UMrTNtJE63hE6YoUv49CFGlOc
+Y1itE2JKPdU6dwSarlUsDdVwvYJDa9sZ0m58/Rf5Ua5IzXk5NNSoAwq9a5BjH4N
wuSz2dgbi5BLw+bjg4IcWmZ/AzrjSAFitMsm5HXnzAKfhsECtT7KmWfiyYa8BcTt
QKunvPwNWkQyiGXFq2r7CSgveU66BLJOcg5Zq6IQ9H05L5Ym4yYXzCJfUDh+0szh
`protect END_PROTECTED
