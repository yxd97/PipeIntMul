`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWcxDdKzSSyG4WPz0Uzr9kJf4bxE7v7JYTWI0GP8gC4i7Q1deZPjUprZhSrRjQ9n
myq3TDeTX63vG+AQKd7h6Ks3hU4PQFo6y13C0+L5CJWTlGV4Fxs2QWYdFPJnu3yn
hBvbGZycn1vQZk8K7Dz1fNwUBbHIVXYWgpJPW2NvADmgKehUUEMPYC86/1rMt5ol
NvU8hf4eBpAvhdbCMhLUAYzRChmo4Gr69ZcQTjLwQFNQ+pKd3pWGyFuh85b4GFp1
fDmnq7skELA+JiniIeleHEN+ppwF3e5uW5Ncdi+dwdLWuwLv7Ko3l1IA7Nkb1Iwd
fYdmgl72AH7SH/92uYrye2EI1OAlk1xc0iTikbzmg96zmx4ZSvh1Ad3ZeL5DK2Uk
wig842ZiaDH59pTvNkKMcBxeJ5PyF3+6VMtQxNKJqBrcJZJteLa4QxiVM8AGjbjn
H9RebJxBh9awIZVLgDNaFVCSK/1HBFHnNoaVsbvSWzVSgKJz1UKDhXAnOEfhqfdl
`protect END_PROTECTED
