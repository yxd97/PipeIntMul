`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f16TFZifQGk9+i78zZXlbfBJncBN/q4IwDSOSlhi7IQcfw2oW182yrLZrTV2yxf0
eAaMdD63CUWRoxT/XyYcD7JuxoV2/IS9lvzDPIlC6YflBymQB4fyNH6OWTTWKiax
BAFSMFmwDpNhqwnvf9SgogZvnHaXTjz2rqy4PPUxADZQnadqs7iN6yRNGDyKcUEl
EzL/BMCYCc2SA/znuQM28t4CCinVZLTqOIE71ormyhedd3UaCmBejPBB34u2vYa3
jSHNztUpjeUpe80TFNl47ymFRsxkD7vl78+i8xsxVuiMwAg+DhDr3pUgZGr+hiEB
KvMNCuXQmEfc7B53DNo65GpUxVRGpqYDFynj6pUEGNlCNH13cEfwMAgYNCipygMi
KAL/jkytZsCoj7ZA/jg/c0EA1QwynHfG9QeQF8DW/gH8M7TG2G8mzPUpAmy/xz4k
4WFAyeynhjIeqCPbESL0lmK/gvO36rfIkKpBWdJwHqLWqAWJ7ihPVLaIbXpin1kQ
HOfUYZubVOX+IOSztDbEzwYWR38YWGEYedmEfrOOUypjgdRxYucPe6dFP67EkGGU
B33brB+iGbF18YKS3jE2sXesQlosOSvdBzvarvdQpYeGclEbFF45UhrresJLvQom
+dC9pJ8VqfGaqxZwRLPVSxsFJGKBakEOmj5gsmAsuLSRoBre33rPzaNHsUq+1oyD
AayvowGzkcIS6mVbWv1Xpw3rmMKv72HMNnthAwMOILpp0ZG/E5w6JqPlqU/mqmnh
0I5gDtzXrFi/7ZJxrO979khNI9xe8Uea1lgSz6UOl5D36PMDjksEFqC64C4hoSBq
qOFTskMqmRb342jxzFGweEN0mPkXLCc2fdJFbHDplmIiYSpkQCPp3ui4VPtw1PyS
KQIuvdofUh3ev0a1ESAnnwtqgwvrzS9Fe1ZmqmGdVLXpMDPk8csentUhbd6SQuli
/GG3B5GUdzgISjeJCNP402jesSU3p1TAhIYQw0Koej8I+i+2SaOwgOBwdMq3CNm3
WV7pO1YnkiCIQA695A3vcs8ib9vR77ZRrdQ62OpojGNmHtJA4vZajjXSLMAHqjVa
JqoC1dYQa/ZhgvIXKrJj/DuLtxhDl+Z5o9S/a9puiTbneZ/oa+kbKlvGQxNnlDwL
MW18/unyETjKnuGcOlNPGY2DaaDzZfhSY6r39LY6uK2RpqXJvm3z/PqLwYp2rl21
52FKQdNzYnJFd9SnhUz5SJ+Je7LFvaHEF+M1fGeuY9wN9JuDJviU1IN0OHEAOJKi
JztOOB3IHGCNvNvpR7qdNYIURlUWv6GSCuwRSVt0PYNiUXPg9uj2sJubW1bBkWMR
ipQEyhbf2XY6zMwsojx3npGBFKxQjnhO3xK/CfGdJR5TOSu8F0i8RRU7YlmajoUX
QIfXKgfMK20w/KXTVovXKE3+DZ6DNh6bqD5Gn0ubDcbTwvbF31tY7hhPnRXV/9zB
GMkWpkEixuMbPz6Lauaftf1QyWr6uQGx1Z2BgO3nCbWj4jfY+kpdDO9C1/lqbR9b
qzzz/s1AdTafQdKlYkWpXAd6ELeiMpHj6C3e+QaAyCXSrKnsokzwvzT/AQ+CvyCy
SxOGueZHNtfxtlkjlNw2uEY/eIZzoqBK4pVmSv2/KIx6hI+PHNCl6G8W3EFVDbnf
mg7XzsiTVd6/kX09JazhAKk2SkIwuMl0wsmV/dfg1zfO+kn5ENXVW7wgcB4oynw7
/Ol4NtAzcg1s/Woj0RwLLFLAU65dAaLhsbkaGal/zCpOFpkmq98JC+h+TskEc1tW
gIUzBrHVfJ3+Mbs/dpdgcuePN051nl/qbfYoZq4tz4nci4pEUInkwjDLmphFxj6V
NkVmf7vrGrpaGdwW17OI+fkoCZ8mNa4FjIFOetZCuX70ZeXmc2kHvAUiGiUcNXIl
qH0/wT2B+1wKb26jO7kopeWfa6A97ZlHXZQnSmpi4Nb6A21RSqEzDsooUirV1MN6
kVnTcmQ3nBpvSRpj/+x6t80sKGq5tISceS5QpwOKHjALdmmgVvLjMPzvTCWotmHT
hMLHw4ohNazBkOVNbtTp4BHh3ax8stdWmiChjYKKLqGf680Dug1MtWE7YAf6eExH
woEZB2vuDGon6awZYkWBzWJYQztQQuGSmPyYFmVjfbzqyRzIvMQf5Pp8fSWAAMeJ
`protect END_PROTECTED
