`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9SQ70YhG1CY56BIATrC746drwtwDAML1MzI49B5fObvAqSNAND6kyh6HkDe4rSJ
9qhkgms95A7YZwplAas9UF8/XqCDrglxbOookLox6dZgsd60fRA+/4eyhq3oWJo2
xqRn4Z6arK1L+4awyeF86k9wwxqkz0QJT8mEGN27fqH1kwloMJ6o7B8Wop6fY2yx
fI6L2AwzSuCgoV7Mtw82af9gehCVITnNp9kb9LgsKNSxBe8hhWuxiQSBMbexBIuy
7FphYgoCKWOngBeGPYm/xBcDnXUt9kHxLhVesbWEMnKsUhCQmOb3eucbRhp1UDit
oggic+TewuFxLYdMHiM3CL0Y5m8rJSOeCsm6welrhNFk+MhpQ+V4dK0zJreWGCHg
VzVoUl73VApOPaidQ3NuB56julTASmgpcZPQIm0LRxQ=
`protect END_PROTECTED
