`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y56arZzreg7XlueKg/bUKuBvk6w3Gzet9BPUnhNj29BPfANEPO7nFq1Eqet9e0Fe
NB5TKVpuPdsOUcse/2Vw+wwzipz8grJbZoB2cjskYKNyTpwbIG1/r0j2BeQCP+rF
Zi3tD0dTkMzTUBTMtLGeO7e88li/Ah+t2UMyYk3a+IvXFgkD+BW5vliXfoh5oU+z
uZiL+atL/pJYAvI46wCBfOeb40IbMXCjEJ4ttZXVC4aF9mNbEQ/z2IvKOTCh8pHA
MXRlUspLnDFyTEpdEYIOE9u3wRin5h1Bvy1uRZtGlMLo+qvGkGR1tU67eO6scJwL
RdqW1eEIT3NGrzWM8bUwUy2Wq6DoliIohPEJmZhsmR31ZSIBW8LzOFrdhdximbHM
bXS2bi3RjewB7ZkcGbCk/5SzPGR2y4eU7CSgvHuSLT3fYuLBZ42nm1ZPndgRFKkS
5Mo5ZVp/L3nViHr5sIw4l+wHp9O9xPsibQniI9ovczxwjo5sSOvSHvqNz2KFAb1B
oFQxG3ZfzBLPgF3VmP64vaFXqBi99Wb3cFfgfTsRSdqq5HAc76et90A+/xzqsSus
0kETxdM0QhLy5PgkotXge7WWgCzT7gYplKD1vXSerGuJ+A5cBAj4FFsVbifueLbA
/ymHFfkHsNLy/0kG4vaFUZkeX+zceu0VO8ClVH35xSRZfmuwlTEC5pzAdVJw3jt4
1Qkkp6dwXRwNELTm7egaSj1PtSO69b80iXl/3pkim2TXdvOBMEoqpA2TaYbd4VQC
2xbGh5vScuYk8qAn6bTLCc0cmUQ8+LOmqlhcDP/i/8KCltvFsqiin3R/GnFGi552
ZiT1ix5DF9Aqm8SwEu7nD/LhlMVuPHk5mo17lg63po2orDci1JkVaJD5ANSsjTlN
5WzSpz3t4913L/9Phout8zHMmtf80z3hkhDZss1mjZBN3mRImUqv/HZ5O4HDsV5f
O5ROpAdjCS77n/+Y3PB8rWN4AAToxem7SoWX3JBX8S49sPnPbvcLYCPpnsgl6pJN
MwUD07pmH4ccEHFVh8FzROYxCpWcbYnTsnOdZef7/J0LwXnkGiW/rs53LqVYILKd
vX2N57ULZAHj6sOuxOisAsL7XwB8JuQ1vJRZprMT5QawJkNEUKmraSL2fRfagGIV
6tB5a1ZkMnsLrxDmo8qWmgAiSrLullBiWHEiAcZNpifD1nHjXwT7D61tAusmjerH
CTivyJLafN3q/8dpHtra03ciZkgVpqZ0bJxpVncgivYJ+4hYt+jczariwiiStlWq
1PxpTjecDRONVtZZBh53IbokP/n8VQ6RWFzqVjCgqdCTJja2dcomDaGYZgFCkJtl
e6b+mxHNoSFtasW4NtG58MRZblWi3jcZMvl9zYqOzxqsu4vJsFieTvQUOOLNiLKh
JeLcQa2HrcP1NGuBcOnZslEvzUe1jkoEzIimeWHoBPz2fRqc3rRZak1aJ+cYkdyt
oHuog2JJcrQYaRAdactVcqRCaC4sbE0eS2SA6PAzJPs6dkHQo5efFJqJBgjlKCa4
CknR0fkhHGrNQEQJZLaZFWKy+ApGsk7vXZDeaF8kZE12K7cDCEwvm5rWVsmuQ/Wm
VRGlk0OyG32txS/4sR6S6fJT9ztmK+U0LRkXF+Gq8Ebts2tBmPTNlqOoQcJ+tsQr
dq3YKIZm6gcWK0VWlqRD2/XO6mNSK9Pk8JyZX4cBav7EJbVka3PqSh28Roh/fK/g
3mPsbF1JRkSLOxZSM/wqBumKkhksr0HnZVGLA2dKgFGzDkEflaYCxRKU1floBPKy
kJ5u9Kjbk1TH/+qaX46KCs1DihcTlzln7BGcr81/FM8U5DKPB1LM9rFD+dTXQ5pT
d1oZVFmFHrF1VddmLWFzz95zDIuuVPjThF5oUtW7BrKC6Pa624UHzlGDJ3pZ5vGk
z+TrBuK6sFsNatPCMiKKMYo+LQExJtEFswULLJpup1ftcRUHwskExA72wUpYog4m
Gh8ApO5zNErEaC8p3d7F8yKFdYP73+mrsk4zVxz/bc8=
`protect END_PROTECTED
