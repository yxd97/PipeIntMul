`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xUO9zw5KNPLzntLjwP9+RAzboEbv2Ku0lw2JW2AB64KV1Ed/aHDQnKitg6Fitv7p
DrtdNaTkiJogYM14N1M0NC45dDGeAr3+H+hO8LpH6OhGb5lGSNO4RTG3lKT+UqjD
xh70pj0oIwfzL7tz90F0wLjLm0B/aey+q0TufG2WnBtddDaVPe+isJFBYqvoNmEH
10rYTXNsLKbztGsEa281o8nvw6y5LXJz4UWUz8jfP0yDrqzsGcofXrycdOMM48Sp
s+XeUf3vEUbft6dz1ukUa6mi5+XWAtMxKx1FOhRBk+xSqkCccHyffMKXSyB8KfbM
nZ0Y2HVmqgScdhBO+k2bVxBeVHjf5pHaTVvA4bt9qMg=
`protect END_PROTECTED
