`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qT/fu5TJuh6uOuH55wIqytci0NZJiAlRJ7Wbz0ut9JXkag+P9/ZbB1LUufGz69Pu
dzEHlE1cGrYkxFtYpswi0dz0F/rSsk/LOBSV65tf9qfNXtCQrTT9SSycuwHaXkhx
tZFcW0+Qi5MjJ5GeUslCrx51xalZ9GO9F+69VluiK6GGXBPnSbce0x5K5/T4b6nU
o9R7kUetGlLVv7itF+0VlstRTcUZQVNc03SYSBt3IH83MoNqL0rgys1ZoFludvDN
7vm2r99oVxIMYLEGmBaJm9XVXOoYzq0CIa8Y1zanoZ71JRz2/neSnmm97sbg/sCK
FQ8/RBwcnH0gpC8PRZl/lafZtotecpLii0/ww5hCamiF13x393M0rUTVyR2y7gKx
DoOuptLPTm6Ot0ekZNm7ur5O6uYAXq8EdSNumZcLli8goWDDF8iwTrD99EXps3yd
gmN1K9+K80gFHAeBgZb+9Mh8BhMfJihQAfNW71mvNSUtYND/+EgfHQ3AbeZgsGh4
i26XsDTU9TVzXHwJWOdx9jXa2w76IVb8gsAe7IRzqkzDyz4rNVostQArYj5jyHoL
qfflUg9dr7U5j6X6OeeLTQuhDkCZytEv3xvZK09phEIMB72Ou9JLfp3W3LPbSRpr
ZuVo4YUI1mcdZ1h62PTLSayruI71Fsbw4s+gTj8b7ec=
`protect END_PROTECTED
