`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CgkwXKBKCqB0cp00Jcn03qsti3BGwosa5lacDfhfhxLmJYz3DZ2XdAWQhNgXMk9o
lKCWsK85IRAgioyDRpz+anrylMgifyVQSKqnQawFGD/+/CP31OLuo0K4OIwZQoJD
2DmRNR/yyJWFP+KqN4p+cvbgBXKktxE2h/7czsqldsY9OBQPOkX5mf+Vpv+LGLD4
LL96jFiKOcFCSf6E0/75ejO/fRBX7m/8bKLZwHQCDM8ZdS8TocFslkrhV7hvfFgJ
OXdXHbZ4G7knSsNgyIvnSlmxn28aNne0q8MWb9bad4OT5sC/RJKJQov3vVKnzRC8
kdHClI/Y3XZvUQ+tR9ClxFNZqfIW2wOwwETUMnlFtKHS7hQ90oFxHv16KsThQ32Z
FJgkz9A8FMbMz0c/bTSo9N1Wf26fsA6qDWlDAd2HsQDBL26RqSe9RybKpiHuot88
`protect END_PROTECTED
