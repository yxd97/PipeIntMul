`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xO+MC8LrMPC1gfeTlXZyiBbrtAt50/Z4eXsihYogQ8TrN1n/k0sb9KugOf3kqbF
duugxuOtIIL5mT+Zpshj//7fEwdvddA9IelUyf0Aq5FXc1W8cnq7Gc5USEeUAzo2
khitG8+aSAZ8msStXfIGaPL+RLEHbO+DDFGGT14xkDzvH1JsjsmhdR3YwgoU174p
Y5kywqEZkAqgT+3NWKhB5Fh3qdT73L7i2sFU8Tg1u7dYXTXXdhhtcCEM4ShCw5go
vTqcyTUHfpineBkZQRQUZ8B0x+KLpJkhtQRb/dIz0ZXMAN1Oz09A9HxeajpuZnId
ABzFdeUxQ6I33Qe+DhH9MRyJkBy7wJWOAil+kruxKjPAMuFz8Y1JjMw5/okwesmL
U6kykOQs8sR0sua8NQxo4Z54NJ/qTDjcGqLyoQ/9WLsrr0nSA1LX2mz4bXM0vo5E
igLkh1/RHZBSV79GPCy/6c5dCDYwlH27c3pNYmD32ZdAd8HilerhQ0+XK0QOAggM
OREB6X+RwwUdEPImDM79FTRdF6Z6e4Xh/dqwB3rvmM9CQv5wfQ42nfhS5RfTy13q
Ae+A3GCeuZOk6ObS/EwtB2L5kj5KRdDOZM7sIXQk6d8rk2t8U3dH0eCZctWGF8Js
ORzJ5SiIBl2yWC+8viTS/ORvj73fArCY9PVQ42ThEkGZR5zUkFxvsEBtYixhgX6W
NLteo4dQsYCbm1YPV7sRdohEWsgjxKegS2sGgmXHq/Q04pW8WRE12z/Vyyxn0fvO
4wvDl9lohHboG+1gM0irWeBX0vxG6EsI2l2rgWg2l/pyR3ESVNjrwYFvHWdtLNld
QbYMClwN2K4XYC4X3K4D65n3BQf0KNRRDcSXgRgqkpKRlmKpHrUoNKCVT59RyIIk
1Xpwqj38xu7CZtU6TcWaETehqG55xz3TSwWlMksVHI+P4wKfPFvAW5CbN6SUQE6q
2eFw5B+yNTca+jcXZFQZmV/A5KI4zMu4Q65Fd6EX/U8hGrxmsaT8sqwP/OpIPJNO
GU/rlMe0yFT+TLyQQnW19PS4vgnVbVyXUPdQBUYe/Pl0QDn4UfS29yrU9ri2JFJN
dd+0SEDRL9WnEj13/liEm1CKeTzDDz888ssHolaAzqDqZqH/AA2ew0p17y3q2Aqi
E6WxbsEy5eXLIyI9zbTX07qTxTNXa1/we6Us9C4Cuk71KCq4iMwHwQNG3K7mluSh
Osl/XXmB2b27z35G0nrJadR3tACFoY42ojGGJmagNvziQRyWywYZwEPVAY5KWlqK
En6icX9P5NKgwxLI8fQVs2Pf/C3E6iA0l9pwKQRFGhl6U8rjcxR89cYsaHjffjp8
lW2owYjDzBwev0BfAPl9KzginKQJhOp4nM39Gdx+Ucgb+T5sjeNOoXJL9GG2rSd/
T6aC8FCQQImgmW1xt9m/vpOC3bfYAXwPmbwC2+7yO71fdnWQyWHJPz7q72OruvNi
fvSXtqcZyCK9LwHSF+dFHpQ6hNNmeDLcutVvF89IZoejvFdFq3xCN7vbv4WAyiyt
WJjF5XRHpQxHEQchxdq2fVQVxHlMzVydJIRPU5qdcIb7f5hvZQx3f7O/tmUjGc/d
QlCSvtYYaTK6PLW4kWwYyQBDHk3L2QruTx0ihVFuo/F3u34yxXEaemlbqAWeR9yp
BMtYgne4wNnKPGplut7Nub0alBmlRnnRGOgMEYezN16SuftOVj2mwHa3ZLaQv0sA
nyikPKdCuASxBsMHhhn0NVodfXCeU0JdLOOXQIHzfML11U4bM6bVeZpeWtiBpkF6
99LZ9sBz1cFMk7VLd98dgDu6IIyE4QXz7I2skEEV03tLbtKxayi7e6e02IBWnKho
XiwnvqOpSBT+qiT7d5RwFSeRWQAyI+uWP4U47gBp9sIQadWuiARAoNY42WnRyOgP
Hju4UMZ37m49/PMZRRItJaeMNAflEkVTnUbAERGfO6M=
`protect END_PROTECTED
