`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3bXXg/vAedyUTKNlkmub3iMtiXQ9a7DGLNFSFQzFv8gQfdMoMkl2waoA4UYZ3+n7
LbyfI+vsUAdqNOFRJ7c70I3qCcj7NhHy6kYU26ZG0YNIE0EBS6mYbDqjvyCL1num
39h5UpcVBao6y6uD/K/bsHcsRr7QcXtebgT0tpuOcR5IUHqcEVYQK69tbgTVflcS
PFakhD88Posdb4coMIhgus2ryUhSNEywS2FUay+mA9wjaVj35U5jxxfHFoLcyJIE
7175ChrdVindqyQMZhS8v9ViuqCqwbRgrLIKlrhI9yMGVMt2T+Umd3tAxFPsAWzT
h9m1WSQPAA6qzBq9nW3mQc2/iRDNMvv7WIDkN66SmEW2r2mwDHFWXNLZb5N7B3kW
QP9WSwlSU9MhPmcijLveADuOvdMifP6WdOnTMBRIj2HBjB3n5ExMbkoWPuuUGpek
GVZpvkxGSR5JhgpQbErTql49C5M0kionVqK3uGp8ROTGCAAahn2Je3YCmSPObTcD
`protect END_PROTECTED
