`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0CcNSkn+LhYL3Xl5fE0rTPmQjkOscvDunPp70GY9TDQaRClrVCY55CtIleeBFF8
jDfKPfmq6YGZkVzLBx6Refys6TKk7sr1cgAug/XvjGuO2sZZ4iLYylH/f2H1U+WW
LZiEqlOgleT5487AeJV8YrlyThgFuRAI0Pu5MuK/tAm3XSd81VeyQRPaKoONjhAD
1lc906QPH9IuVpdC3JhuDtIBHgvrKfJ0a0uZInbFJpOQ0qwWWmOB9m9Yac+2G5xe
1DQokSZe2fJBHTPFKc/4l7fIhNqxChCtfGvAo6+bMyXt2pO0ng+EpzGHsrJnyf2j
S4Wwy7H1CCXLU0SQ7NWCzQ==
`protect END_PROTECTED
