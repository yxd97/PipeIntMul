`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0mTcFtJER3njUvDqRtGmB2QHkY2eT4XoIEgOP30uj3g/CPxtLuNsO5WGlzpU6zno
rNizT0BqNqFJm6p0tBNOdFvmhZ5e8KAPHV0D+V4JUbh4HjaEVn2POAFs8buVl2lz
GK4tySZK2NiWgXFaI71VOwlyFlW/LJRDH6pYcVU5GNL5fwd6IVAAZACZaAAmpOHH
/NxQ5iOFFwbwkS6p9tffvjV+J/M52J+vrHL9MOxxfmQRsatj934rAqgfcUD0kqr5
OZQrldjS/Qwfg+ct52BppawdTJUai4ffm0VBvOAfsu3eUw4/3UplOD5ScOT5437p
moNy3GgTfgcZi3CrdpjZ8jSfgXLSWU5uVCcRXVkpuCKS5rwSj4JDZ4WO3xcqq5eW
/Iuhh6k5PXzrEfOpCjRhEisGHoqJR3Zo0iksH9qF4VDvC/WD4Ypzi1Vq9/GCtofk
DcYSt/1+sXovJJZeRwPQ3UZFnDQBQdHsex0Yayn+dFqch9Mab5zjcsgWSpxeRe0Y
Zx1eIqcozYnJ+vnw5YkWL5SbTkAFk/IfkInrj6m+hrHo06ZU/iv7WcMmHATXYGC9
5LJesFw4k6Pm5D3RsEv5pvSFQcER7XvXkjshXZH7C9ueb7JDjFNJQD/vp7GWjbbH
aqFZCOjOSGFcGk/yNtmeBQ1FqppUUJlxTYeyQERhM1osSfCmTXSQ5JFKhocstDAi
RARXOaVzWYhaQueWZmNToM1MEOKwjJOwVdD+ubXGtP5aGuxYeCKPXl+OA9DyKUT5
FVejLOh/5OG05FKwTetLaAV1ffZtFq7D23t5r4g/AaE4LzuZdE2Zok/mNh8eAscR
dpzts6vzCM49GzC5CPy3H5vdWWoXfCxW8ZgbLKXUq2UTOnfAb09zqi3GZ5+yhi9K
EZaal++3v0XS0goiKQJvweuM0Xf16akbgS1QHrN/VXlOZdC6mYG+fTUA/DIJDvyu
HAMLf/WvK40VtmStQ2UNUyOejvWGgly9DR6/KpkhQLw5r7onJ/hpCV1EpWlw4A29
rOLFBKfbAOH6gjzBYMWD/vJ1pW9HCSsyO4EFo/Ca35txZ0caMawPd0dnHoA95b3p
0m5XmOgjVfZQOqrY4jE0tsPtFl7/NWPPoaxMPF55GE6MEGN3UziQmfyxXaqlgunp
sl/Ng8OrK0ugOXPS0Yh164G8DfnJlo5GYNCB9R6Oe209R21tdFmK65U3XWdrLrW9
uSxLO+lxPTqpj+2BK1RSIeaFyVNpPJw149o3CKuZGT2yektqyOnOei6VCp8MYcx8
ggBdu4kk0hUKDsTfMwwfshUsmUaTEJKy3jgcKi96RFrhHsn8Lq2wWa/+ORpEzTLj
4WvTO+m/zKz4f2M3azDvjJDEl85lA1bmQXAlRl22+rDigJU4fBUJ0uRa34dg2obC
toEStQQo2oF+ZgQKakxrBCy+qzBaYQmGaX/XyzHLvt+ANT2At0gP3jAkDmmnrQYI
UI+zdJdQid9EbD3pcjG6Hf6dnWjWH/9oAzGtVyDO9pmR5jCEO8NtZZkUjK6MkYZ9
rusQvZNh4MSOx+LoLLrnVHvFAPCRfxgsxyvqQ4+3YglFiQ2y+148bhgBeWq7Jfoy
hYjo4A/PdoDmW+uc/IzQ8auJm/MB09tG2F+xlZa36jmC94lv6d0qb6OsLwOwrCAE
euMX5og0lNATRt+2trEU/uuw/Q+obuZWp6v6x9rIw/wqkE7bsWS5bADeiRgO8KXf
gV/Q6OEz0ZLOjatPFr5YQRB8eF2scT6NDq/y3bHcwvBn2UsWpC+JBV3JFze6tCyY
IMLGlEUj3Zetpzw8qYwcnsm87+XcXt9js2RU7JpLvmD9IZToHjtGXulmWUhBiTni
hV1SBPP3gcGV6LcHY7yzQxKSILlB1kMUMoZfxrUR5Yun0UDhWsGCZE5Gl+3Qio8k
xT3h36oTxbBL9+AbuVzpV5kgsg60pNQYAP7v13f9Dz3wQaJrummRyv89Xs4umo8O
PMQxQsqHakf9J5r82zpwlnR6QoM9casZZMNWwid/PF8kpNUjPZeH0oveQhyQKj04
nJx13qcYwEEFKzQJYLqkQ1EmKP6dZV4P1qe1KhRkl9AZrqvS4FWf8e3ZI/z/rnQR
AxM+utGl0xwFPID3MyHClWZjmRVcSJwmNJzPPah0sTffCgHon3U6koxSMbl+ilGq
0lc5HtTu49/ekeEs/yJgGJ/7svBisFyzKHO+MbHDY/3PxDUwVsGRa+BNRbb8qr23
FBH6QV1z/eXtRjoZ50t1olyekz7/8wGPNMIqgfdHDAOCDlmpJStNaNLs/WAt3gCi
cvwCaKEjZWZOieHZcs7OjnSNL7/zcUwQdZSF1tLJ4W29ifOhFgYVxSEbWxpsQrtF
aTv+aGxMbz4uAROBfGgJsgesyYSiFzv9kGjTsSNydDZZ9W3zkigseVOQjE9jXty1
nrib0jvj1ppw3Kjn1BU64KqCwO4JQynafzoVjyFwCOa+lP+B1ACm4axKj4Ba+6Xi
v4ge0GZiUo5P3Rj7mZGyT0aoLwO/tHx9zXRvjYUrGhZRgJGKS2dOZNHcOZSIwVBq
d0zkI6HfRiXoIydlYgM3QcFzD2RY43EnV9eJ7ibIEyfZXeRYMcpX2tK4TW9++q40
CrGri9uEa8J49wkHzdYNdEuFcze23yEcUUHb801fvsrbX7FeklfTduNyxRlvatEs
JWGDZRMioly8tRoQERIeW6dfDMVJSCXspRUJCP7mWp/XGkwCTT3zxNnEmJxcf9hf
97wDf1tQFoxI6/NWBjEodUC+NBb85X0gyfVh7hVK3hf5bxMt/rc22KzRN0SjQ+FW
LD6lZNMSLE00Bk56wZjVgFHocw/+cPgbJ645wGPWKM+r4aDYqzpCveEPFWNM7DlI
vBLTG9QddZhn7DqVoopXDLYghO33SLr/232BHU0qNOxm8mGLkJ5AfbqDHNDFAkUr
lNZOVsAe33voGUDPqCnwnRFHbtXx4kaeBpgsMTIhSbOwHXIpPE4YDqs5O/HuCbAB
Vt8Ef22S+pe0rp7sQjXz/g/ba+V8tn19VhtYDzEBCeMU7IsQEutrd/PkLYCbgGc/
LqMpewdbttPmjgYIOXXYRf2ePmx+zOQhaaVNtJKxlSm+kc+m3wYtBSNk9BZrHeKx
T/oRCXdrXkXMZiYBPSmfMdj/zQEvWzvjB79KLfHIE7SFdCLefdk9b9R8BOOO/voV
dvB+FJ+rwV7DhVw7/ErL96/JCOd0QnqkY8tBdGPDzheqjKQL4TdMqzYSBwhfR89Z
Cn3SlcV5mwAsHkwm6ase7Ymc99+c9vHO6KIdmUEGtdEvzRALHj2jVJchozW1pP7N
UwDuqoZQ/4ngf0S+F7EYJQlA5FWMDjoPOuwFT/ufefdK+MIoRy4Aoz7V5QMa2a16
acOKlEnIqyo+mPlByF02JD2tyIjKVqJVubgKfHVdpULfyNkkFVzKaHBM8fA0fdPz
INRLYYlfYbFIUVY34hIv6KIDwo3EOm6xXfJTBL/cN3WQMdI7AOUZ4bHru/7w9eYr
3WNvqcYa9XoEOFPOLuqPxiwh6mReTIo9qCo7d0ogaQI3G/GO1vc0QGN7XX3UpCJ3
TnzxJTBBxcaTCUOSOaIXqLhtMQxpTcvDSY27osg3IBY/wk/CyD4YMp0SFpP/Hq9R
hLAZFaVeA/mHnEgjaxVoVWAjxV+oEtCOVTwTH5AG1ZBCPtQVXJYxSqRKFZDKWdL/
sC4YqX5mvd5gkhwmR6MzZvg1bQOTz+1zefvoxiJR9vvg1Yb1VZaNVksmPJTPAr5p
PsQpvH34Gi6fZCW/gbhQPIpOuxwkQC0GE8FW88BMyQNUKuXLM7RFISuux4kywnQh
Ml47rBlcrwiRwxnEj4YVw+SI/YZfY7O4XyNJiD3WBKUmugONslsyMV+HaQ6CnEI6
77ZdP+dLbpvNYVB8UJQXxPcUJri9X4jnkArb9PhXjkXdMCx4UAiLDp/2UsRjv9fA
zw9AG12Q6TscYo6w8t7zdVk8Ets7fvfL4c4/7HgouSCvD19nTNILqrxjP3ZKaGqf
Kz8rcS75fRrQTd9RLE71rc+2rAyt34zBPzVHB0J4de6AyF5kY4R6oxalX9tF5IJx
5FrO/sIh/MHWzFftCvvXnG4Jmya9mKd8Cl/dyXbkpnh4OpcZ2whCTGYznQxUU5IN
dD1T9EEH1o8RnIN9TsxaqZPRF3rXvPlJ9PvxZmA28V59IZ80yOWpppp/QJafCQce
0NBTnktvm9ZLOwsf1l61bco/BFortdim6MH1HNnnvKboxPC8+7dfj3sYmUH6fAeZ
YxKBOaiEgO5KmKb+/xHNgp40D/9hIzrcuXxIGC2UynF2Ln9pjC9LMP8/HNlk7gi5
e0L+1B/9Io/+KBHHWbOMEbXy1VrmiWVWTZR1zE6Pm8zRzMNcYgVjkS1daSoMlMIk
JJPkdfbNPtZjSe8PFM3n6Af9PYfZWKhJ2NNA/VF4T3XxCIBR8rQPTEmdgh47sBpC
BFr09gYRne2X3q4zYf4Q4EIGAK3X/vaiDbMAaXK/AJv4Tx2cXEM9DFkIopx0a8eC
tp6cYkyY9Pl5k1Ukc6FLedojbXXa3l6tnVEHYj8S9sNAJ7iGUKmKWzvtUpEu4d16
k7UXPDr+V76AUqagiLit47YRAPbrPTF8XQcurKMdIbCopY1eXEu/SeEkK4Wmy4qz
Z1IBKvY0Ch3+gDec3X9H8pMfORYNsm7VBymPpK1oNQY=
`protect END_PROTECTED
