`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a761vjVnc3Zo8p0c/0Efe2ZPEGDcMVt20jxAVLWTYV5TLmIxljUqjWrvNSldG7Zt
Zsz4ITOHi6Zk0ty9G0pYCTWU4ltHYxuh1YXb40Vi8OVzJrOMG6TgwgovQ6rlB+gD
R7fnjEiJqygpckNjKRuJyv2xXTDBGefwXkXTl+iPvlwkSE4qufNgNVYQaCRgxjYL
zJIfsdrGHyij0F07FnTKutBiX59bfV6uhGSIGxJBt5nvUGqPuvWxZb+Ufvb5jo2N
CqllYt31xTtqXJm5czRJyTAkX3/NVImXnnnwG4rLoTh/ksPsRTIauUWGR707kmFV
W71dO+5Oc24LHSGKYCwpWEeQdlosD3lp+cmTGdtTYlxzUG6GyOhLcsO3QSJ00Tex
vMnZy7yTH5K2MwBbj1Pk25X3y9sJbAfp4YDADFViWbo2VKDhzfHhrka0rqlSQXgb
LQlF5YqSywFVOCYendsK2C94dFpp+fqsUpHve0R5OSDFi1Kxm5Np/uW0YfqT8gcW
aBbsn3oCLcZ2DbljeDhSM4ax8C2O/i0MJDTmElB8JgLfCaHK/YKUuZRC8oUhxLaZ
D7RNC8DX4kxtC5pauo1JsaZpUrY6fnu6zCCShF2sB7fl308sF1KvrLdtWqSOCMq7
hy8SvS5M6RjEPU1Skesv55WW5SID8IXIJ2I/kDdDfwT3E427FUbTn2V6hA2l7wJj
3F6Krn3cIgTK1YNbgQjJrKDXqZwWWMQSYBqAmq1UawKnqlKb6kPifXu5ZQdanHHT
VBWqAbGKfAXnROfLgGc+Tcpr2zCobW408tX+UiqBmzu24/ENuBaxOvHWPeXlyNZ8
VdHYNpf1k/+AtwNNr6GTAdjQ7vFj7rrovWlA0ffmVpcwy0lPuf2DzjQ5ZcnLVWm8
L4hE5jgqDrWriLmIlArwMJHTgaRhLfIBdUA/My3A/Q7zPLNTze3NvTjkmufFM34T
ajEp5Zwg/SeK9tVeMmPgS+emiNEjtLWechon7O8u9C0XjZFTCEjYPwZFaV7xf1RI
qJTSH9pG+eCFTCKHHFMfGrkP7lEKCt1P6Be0Hkb0rn07R2gi+CuRRDPaEs77+y1B
eQsPKDgAfGyId14xfYQuYs5tRX3V106rxFtCiWoW6yiz0I+MjYyf5RZ66uQkisZ8
IwvfvUxaDOaIoKI1XDlL3i8UKbAsQlDOkWhqcW9y6IF/35uUkDyFU4weIH9sFyHF
hD1GqAIUgJ92UgMdpjs1hT3gQFUGR1okPjT7HEN+p3B9/FCNbBzA/4SblF7H/xMh
spsgPKfLUxheMYUM8Sa3SfrEK7QnCIIDArZnt24kFpGmZBxd07H3UXY0/VpOkvjd
0uVyWWUs41MZOhqvHTduP54aWM5YNPRbyCTAatSB6Oej3sQMoN6jekJ4PXxYQ2uv
fY4/Zv+iw5q9j2Cs6VbzY/L5C7woyC9qkG5g3DHRXcVE2KH0ipMyfgpLFTt0bhsO
DLOA4f6gNUcz5dvgZoq6JRrq/Mt5iWJAdVeAcZSSQHJUtM9Bzz3AxZeQAcZHn2AX
RDoOCP208Px34//o6mkSiECszutb2wBDncoVoE+PihyeqbVF9JQyuiWT+g+W1u9i
8y6upSiYGEJLznSEXc9y8OwMqckkaThbePo3sCxWNASuZPmLDEizoQ877q1xX4FT
AgB6BDRS5iiV+vqhFf+vHocGxlVCBaGuwjYwK2JV3UV2AVKZYVWZXY5pUdVI0Qhp
nIglk4jvKjnfMi3Q49YjOmG+49htw45vVcaSVwGWlpo6AhwPx1yjQlS60isBzkSm
aIe2dy6nOIbwV2GkErichWCltQAXSBKOoMBlyrVhj1wa7HH0sTjUGZ5DM/eSUVSw
pdY+AmtQj5FA8wgQetWOhGLQtinSFRVar9fmJulMcd6HO98iqUwwWR5JpGLpqFCq
MvAhV2Dua9ga/4Oo9aMTBVK5glz0dTyF1IhW9JQSYYoYtIbLTxJQ2lXcjKq8L0bG
F60sAs9LhGprRntZK7Vd/NJYnrPmOCeQJ8igQQWCSiQ++RIEolMyQO4vIwKLPq+l
AILf4T/7IsuPn8h//aXqIiyaJ3gg5OrpVB2jJdu+lV1BRJWCEYZ2Qstg0xDbB6kP
`protect END_PROTECTED
