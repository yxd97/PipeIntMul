`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxCDga4uIAn6+AiZFtvco0HRIHnfd54xatwRFJomxKdK0ki6xitCIRCCeWIYKrPn
W2jP44DQ4KmYnHXeh7oNqzSqn7wiwu0Dhxu7usar2Lf3+Wen3HF9/1I0VB/rZdwS
npP/4IYZTT4XgusZOVCiyz7IAdkciXBlAHjaYgNlQ7Yd2NW6+/ySAjX38FNjHcuU
tO3yii6wUKRvrPLi0jOC1BYq/SCx1VuuBd1jCAF6WPvxxhyAvYm/7eH2QXuFc2xM
LWiWcY7gB96bL3rctqz/MARNRTDpblsNOB4CiARqbdY/Yx88WQdJj1NOcjyopy8F
O2DHQYoJilpF1IOUOMVVug8hus2n2nnL52ORsXDoxolTWJ1OsGjnmsL+0dS6uz6P
EUbax+Mdd7fMMKIImOQeEWz1QVi4J/J9ZS3F45v7cGuCX1a9GaK7zOkK5tqul6jd
ojCpFbwNUz/55adwUMuFsj2VdSBQrfh+YeEApYhAuqdV3znkRCAeh9rYDHbvxb2S
Ni2WXSUyX31lW9JqJ6ISKAr8woSUf18FkdKECyznR7hYqTOG96ZArwgGh5EHzV2I
25kBKQdyH3OkGck2i0PeXa6ZtpRW4YoVX1GuwHo5zdLmc9ICPm8by4sOkJxRXLXc
W/ETWqSJHCFYbE3A72TOnaKy0nvDco6GltQON8eUvYRmoid5tIFomnDu54L6ACB9
0afaU0qJxzlzesHN/eGipzaEAW5qHXvsUFX4o0nwcuZkXvuxyeZh5fsribMFRaD9
uaPED/OnLRZgKw0otWye2yr5Bd2BQehxtxM924Ck2zlw2nZvu8A7MalPNUENhZKc
gt+1RdzBafoWQcXXNnTGBNfHbAO46Vf254u1zyvx0katROIw4O/dn0cKeH0e8on4
Y61OPX/Es1S8WMm/xAnNyqAWnz0n/TLgx2DgBexySOI+J/kMLXpWu6i3mg/sQof0
0GNAzrvtPQeN+OHE18wr2F8vyXR3fXKV/YEF/k90lLT6I61sgS9P30IpJDeqTPVl
JZNLpoRx04LDrzD0vZttv7Uxhr3ig7w3RW1Yk1mHg+b51axuyuIHvXdoEA2ee1Qy
xiPfIC4IwIizHG+oMEiwDOsD6ZG73vkW6ktcO50j/Ghgf4xyQG+UeajGxyNBN/fG
oCppNrlJ0kfLjguUjwESZxtnXVIxE02xe9oLGoEae4q/0fpbA3sbiznvo/QkCd9l
Sl2lNJWqNGIFEgMBQ24knQQyOfDbzhKsjGCOitMz9Q0aGsqYCIV4DTNjDD3wnVIy
UbuBuaiepFntPoeOhtYqcRyXhVI6jyltetQoMDhFP2n6uhKDAL7muQEULbRObVTq
DDJneI0LLS/bPYj21vJAuIMl3awiKywbm4pc479A6rwYLoiKM5dsSe0hMvvIhWCW
qyNkK7RzF5ckEl5iYJJVDf3FicWLmT8ljJSAJahm5MDYcfDTwBKN8up2AEzvpiY0
XIrl7gab/1UjwUjuFKce2x7j8dDkMHpgijKkPr640IiQ3nry0rUSnpK6DxPbz3VG
7Qvo/CpjQd6zlvmgojpFz73KvAPJHkPeT7k1kCihVQmuwkKGhdcHCMXMVijXAolE
jtbn0gsjv2tcWo6i8VqU39+Ok7xB3LTS+31PJw1zs88RmHaN4DqTcuD2dDao5lCs
T+0oSclE5Ov93oQhYucL9NBKb/eSxkusDgH4/iCSirJzk+uBgPvxHcjLveqg6kdu
gDG3f7T7cmEQqwWnTw1AaqRjRXxl7GBOVn3jfCGGsw2d5h8Udv95HW0hx0ojeX8M
R75dx5ZOQBUdEp4jgvc2iQxMtUcYOTFVha9DN++dEhg2fvIwwFwzCn75KMHT9si8
UWgXWyqq7iXE2ywQ1AQvhQz7W8gTPGhBdVw57Bs/m/XrH5I4Ku82TAOCCOdIQLvz
DBkaxKizq+A4E2+MTD2+3QX85UYZYUhYPODOex2BMXDUMRQdSi6jKhsDy7lLBcTn
pxLgecvL64j3qYXQMIfNLZWqlT3HEv5VR19QBfmDVdoYLGUOXxw8nnuZ0oDiM8wd
PIp6egbJpK2C/ggLI99crqdjxsjLHdWCeucnVnHHtLiF+EPCtMAgQQtSxVUaYMJh
iVLfiCUnqXjBil+IvyKs8HLdqF5Y3gd2FfdBez3IOcqll+kS+KZJ9ZLk8h461y8O
GNs7ge1Vl+0+5OWnYQkTJJMu9lf87iJVncv9RL47BpVvt574oUarDQRKQrou7lT2
z/qngq/ZyhGC1TLlR2uDDa4x8DBxgQ5ul/A4HVE1pVQW+aBPTAKgs2cQmwEuvHZ4
oGbJu5FpNgtRiBblqJ68XeEhS8rKbSw5KQBAN6yF9n5ZBjiGdcY5aeolL+JI3RhQ
ZIB+IvJI/oEIZ1rU+GnrjKbEnlMpl/0Jga5m8xUPL2ETCudYGOlCWRb6qwc9q5Sl
iR1Ub5BhR2fdJ69ptKx1k2CekFpq2lb4lQcDssisVMbaBWYVugwwxk5H77/oyN6V
qJT92Cv5PF0qo6pAQGo3dy2UYpBsrjEoA9HjEhYfPxttbRwFaZLZdt9LG3bTH5A9
AJ791L4Qiig0h6HlJVVp7zQGMAA6ZAS/XMQwfFy5IAf4/xJu9a73BzrIay3Qrd4N
NpMJlXYuOaD1Iq5YQqIqmvM0G26ze9ZMgyiIxc5MaDhJ7nzOMoiBkMaAKpXFXof4
7VUYqIgSJyKDCzQLF88mB1aFySJE8O5yuejuaXoEtX5XfOc6wKb2jumx8UFy6QZr
Sa9W67Do0oG5ltDO9f6mwgKZm+128yfLONTLq43mzZi2+L4ZvZqoaptZ7dBCAoQR
51KtcnE1KKIPXggmqywofBTkRWgZZnRZes6v1W22h6wnRUURyzSYudVDHidKKYMx
roLTJff/eHEFHrN1MLPOmdwnd8pmzcAlDA8vYtbgF+BCbqvhhN4FRbgHq1eTDzGZ
y4CmKyHE+gXf1MzbpyM2oVi0geh1FOUDPQYWHS6Zq3LV7kxL1gx8CCs9G2x1oGpp
aPDkYlOtfb2h7l4VPK75Z4E3awEjtjlZIqq1rJMvSNuVLZYiTXW2+yp67eLiMZPm
21TWGabw9p9M8NOuKUgP06SOIwhBzwMcoQ6XF3zSCcPwfzZAuJxbVaSjuUeUVAyp
MMQGgHUGv41bgvQQrnGRrdXwGbMsj5fqwRh89L6QuvoLXmU7kzSdzJubxtoRW+nM
xREmBQUtuvafoq3flWYhQzCZEwVV64xlvSkzBl+GkR+HuLlfAuN4mCG2uLJnr3z6
s5qGux7FPGu90yTBavVvTzSPXT5NvN0AZlB0ITfT6flwq25HX69ISz3obE8klo1q
bpauQyA9hDWP7MFtQVC3eW0i4ACQ3KRRZw6MJWKOG16ihHILWtsoYA0Ov8bweWf5
+tqk9Uw9IglPJvNjcgnSiuKcPLzVoejXD/ou/1S67gcc2A7BUeSb7bP5+DYlaSmW
dDaCwVfE3ViS0UtJHApMjHEMbcecVrPZBbQ2ix/pb1UJL1VDZmFIwshrqq1DuvEL
ZNC3BR5JWhZA3Qke+aMd83pEhAPcti+EKXPlRYrPtTRGoh4Hfx33sR/ipm772bFg
YYK6Ilinf3mBgu//Uh1yPLvyCSkRS/9NRQ7m6F4MkfC8nGnHQ8mTffK/iwcWdDkT
9pOWNzyq3JH9t2eUQuHerJnFSbojOaQKPGUWuoiXXCPu9MJy+JVDBNctoqkvtAqH
khfAZxvPB2l0Sna7Za3sH9DV1uinSNc0WNulQrl/PFIcs9ndeVbM6qeSpydVOI4r
N3VO8A2f5KIJSTUbXULALACit5TXHu5mB8G5tQ2qVJMRzYouvspmrJXOEWoc33QE
nPJ9O1NSpS9xVRu3kYT6XWMHaFbDZg24/1Y3A5ZfgIjUSMmg9z6UbKMREGHuZhjS
x6wzlL0riI0xh6y/MpcQI4Wbv4shZxZjfa9V+s2iTJdTKiF3TaYKVhgxUSLSez1G
4+PVNns6AtWGhpiYCarfoM/L72fjWQvMF2emn4tokXNJcwp6+JTztcBXnPY08IEE
olumaMR95+DOTr24Q8hTSRx5fVmZR6UKKBKdkw5pnVIcSAeN9206NWUSngXPmFkO
F3K4sikqh9kRyB9xAFLfr/TgpT2xuciN/VrwPqyNMX7suTficpSEyBHJ3kbVxHRu
0W2qqJKwk4/TdCN/275eUkXqbyoKXCRtoRZa6N/Pu7brShSTF7vSm4Pk3rRtpPK4
gPW/a34ADryedXWfN/pZ6WpWuS9KCKxR2DdzzOk78RtDfG81vRCfBFcM8mL01nrs
K6sute/Bv51x+Vp8s2UyMnR4DKWpo3QBqeQRFLfmZCtLzf7MrTywuUa8GawOLmm9
RlJzZfgDHoUrQHCHO6+/Rl+7HEiMg8BVT7hpUvH56es7+4KkZHqcFr4kxzz2sAr1
c/UhSObTnFG2xkz/9VgMCT3qgOeuJo4mdjVMfdbTqw5BS2wVDib0kJyjocKYE+vo
WzAGoQkbpvP/2S6JaQRIHY8pNx88uh4l1Ds+Tz3ZuFOp0A0toGC6gqnpiy8I1DuH
6mN6NQ3vzwpzimcfLzNl7HdSkmDo+VmwTnTRg9SPiiJh08ZWkSZnxI7nwYBpEZkq
BUb3fILfmZMRyshfwroiLoNPwg2NzJcSkvlHK7h749tJgbqwBwnjfKlH9Gc8Bf4j
VsWsBpiZHGQINWrNRZeuem9vo8seVkeaOFW9Kxtq7SqX7bIlhnIW/K7pebvnF7Pg
jl14AjK4O+XWD05IP07Lt0CFMREyBl+CcQ8PTqZMasHJfs7bZPANS9BbtXsZ+Sa+
/VNDpAEpt64YSCJ/p6TixO5R+tzU3lqEdRSca+1F3DvoJleZANP0+bUMh0fCfxUZ
qoLmOnPGHsnEEhfeTXuk6XS3gxUTYL29zf/RoRsBnPYatBZ914W5A3DbbD9BaANo
xXp7m0fBqzZjIDBMSmXXvxo8G3EOL6ag9VRg72CVfGDYsml1v5iDyAZVh1EC9bMF
EjSdZbyPyNttuUhSpTZC12l1wdhD087/xQZbL/ixX38ai0ARVxOmbym9DWhzIoTZ
dtH88a7h7ECC00lDH7tpu/ivRQQubU6ZxqgYeQlucWXy0FtfTnPjdoG18cKeEmQY
YxfTI5VElYdlUmEusCh3Em9J3O++Nza0r/UYbMbz8vmcAVqDT51FgZVxX4pg9Sby
1RMBcYpUDR81KfqqA8NXovBItsU2ZJ9ibFjwm9iwsfD6ejRsDg+Bz8rcso9X9fuy
oYUy5CtlKIHYWTuwd0q1ghnD8cqGtQkiyquLGUzw41LTJgxEalekqHeTAvG8iaHH
BCFxYQzGgUhGjsgaW//Obi7kIYDNR5dtCSkAR4nJ5dndjkBTOAGFkzx/XBYLy3U7
hEOYX0h4GWWZLjoz1w9IBa2SJKKjU1mO7YmeDnZ7B+UugXdgdagcCQhrgfnI356T
6ly6QxmybHLip3agL8IeGg/xLUOsnWkBjmUYlnrZtEsu12rVgjEHzY6zpJLPUwk8
Glwww70zDEtat6w8Wq7V7oPSqdHu3lXQGTx6JezRIsSYk/BiczTujAXQF28/ZgzL
zyrwH6ofsSPWmmfwOsBLawOzHuJXlt+kojc4f6rDwF0EBkBjfzvq7jxbQqNmUPmR
ualBph1/5fzXyWqjC3CN89icbCdTPg3+HFN3zfGZ5wc7ahy6gTEhCazt19ri3E/x
bxZ1jG/gbV+awX2cH2jgVKgg+hQ9BL/WIEaMRFbSK2Ei9S8HiaYGniDXSrMVWYfu
ACfMeJ/fzaEnt65NSFgYFLkrZNNIyYLgyPFthhKPVoV+ackgTw3KWundOR7DpaJP
QbieZQ2hpto6sNZON1OgErHpxD1jxsUJC3LFGBYfqV8VIb4IVeozO8STm/ZyNwxA
/otvLceAWjQ5EWh3oxGW5yM6oGvAz0QfUbC55KTaGu7HZKGNTcf/TFb3F48/NF/E
OSxpOQI9Kh0/+MY4wLE6lFzDaG0x/5kU83rG1z54lYOTwmoD2mKiZpjG0fNOReq8
DyqAz0grmhmORD1qQrHHe+Bk99dlmP27rrmCM2NzTQ+MUs+wJfyKvlWaNKsSFjYd
6yhr3m5FDRCMXdIcJgchNm7YgZnCSP9SHOc5FHhR6pQBfbKBp3UMtOQq/Lz5LnY9
mdw/PtcVHAwJEYH0dhaMTJEUhEukiksXtK36spPZUAwJDosEuAS+//9Vk4U12wbc
O6n4RbZZBIOZKnJ18+c4D5tmcJOJaoGwPAgHj5gMygiNy/habyLdn/s4+x+x1Gza
favGf8HOx21PZ6/neSV6fwNzRtRPgcJSPjrwAsYV8SA7qoJzfUepsqxRdwAsdWK2
TvFZnEyFgVSjXqtq7hfpPgiu4c/qhiFGtI+P92pJ8U1njMJYiwHA1uGBSHp3s6tV
g1qTfViTPFHz13xJl6qO6/LlGsfTOIx8dai0ccouwJ2BHcVcng9yF760sa5lhFB9
m2WdJpzytjFhVIE2VDxg5uVbz+dTDjfjB7DCf6uw01ALGPvoNsmMUVz8c1Av49J2
87gjy6JdBrzhJMVQWk4ZRqNexJXV6/3B/KLpFqUX5GdznMOFP+wV+rjfKUoUN1xb
jgC1+BmSMwDhLfopISQqHrCPTJlE04NPTbiwzCsweSEP0JcGV74DLazySp8Cg2Mt
nRQXE87kuVOC3XGsjVwrN0AGIpovyHynI4qc1abnsTuoF8wTA3U0qBugAkKd99EO
5xFOw/tHtOewy15U/GEBq4IDgnGAgiIENyAcaaGlSP5h5VEYjuWC8Vqy+6sJ1Fkp
7PNokKjT7zCZ52kh7qKUkkwwoI6N5UlF53DPDe2oupCJPoelrpHjXWR8TRvFcQPf
yKPfyRmxcmw/7NPJ+Vk8mGFOYPNkwkfIqxsq3C5gONHhk1lHC6Ec/EatRgNRZBwW
dAlt5AEx0dhWv2Osc+sLB4GeWOs9fL9Ci4irXzuIawzJdnKB2I4wKUr2uzSVGJON
Oq4P5kd2R/VVe3RkJKgwbD6Qp+Up4PFxxcsuf5QntZ8YbeIKJqRrPfrObTBntZct
e4156rSkgPGH2VQ8YF/7hWOgqUHkvpaFEIoPDgc4fiMaJOH5BTM3G9txL/1VxW3I
Qiw4hSxGiLANWgh2pwqBsf9SzB1Gg9Q32w664EuYBpqQzk6i+VEyks94M+lH3wgA
1T3efgcEyIp9j1tUrHUfTQReywPDQquihpaNsjRuXZmW56dXlqlzEwU8uGhkLQ2Z
vCqgbMYmT2tZc1yvsDxFKTO+sh7AokvkLv3eKrZFHu4WUwesXIxlGLbUmL/+66KX
0DOF9QRdYKKMOBDuDUU2/61KZ+HMUFO/zHTbPsIqIt/bExD+37H4Ah54MWZYJTIH
pxeyJOFyxF2L6vu6Z+Qaxpb7oSG6z2K1yVkYuW85F5Fpwb6mT5FRaIFoSmcSbhPH
r1NCy42MVnoqFh1e7jGnkzC5j+EEyVr1k9QrF5T1E7ctdIJL/8vfa0ER2TIjrPxL
oeB7pLMkBgQkRqZGiX2spbM6E4Jt8dlLlSvX8kH09tqnj+4v7tPcArvL2zQBAouE
1nAHF98QYyX1cL0LB3/4j1I8jTCRIwANleyBUCRyx05broe3bHnemEAhhouKiIYg
sue79ZQlRUEWijqMTVr8gsPdiqaGFwJ9TbkWT18X6al3HyIbCIiiGwOT3rGUyIIi
7Xx+4qFjVIpFx+YWHKsFV6cThB1bWZrISQLjfkLhU2JyDtcekhzgWh3e3FxyMFHa
PctdFeHVDJc8mtGTBb/OGsl3N8HymDfxBoqWf2hyDwM7DIUgxlhg/CGLG2HLkAf6
4xjZcCSldWIxJw5jYoD8mK1EYzV8Bnm9pMpZj8X0+9OBeQIRqT5jg3qrT2l4c6Vu
v+/uuQrelfL67pVSVaEyvcO1p8sMIdAt7ULrr/s7pth2scWHdPygoph99ckaqLXI
6LZlZtxmfFez0siJzGRXFNIZBL338fFgAexYC9u8YYUkmIHh/alX7CTPo8F8UwlM
rdJxZ/75iI+cTJOFfFYdNS62ohWuwF42iM7tuiNPaz2z9GcvdS8VY9hDdqtIHzvT
p2GlkoFKEUMm6x/mB2s5ZwJo97s4Yn01sWmTztb/oC1tWCFmLnf6NDdXLgytxH3B
7FwgAMkOfK8+1wIZCv1n+jfYZA/VOMIsslYuhsTgOr6zbgNMGFELccw7cJY/CaIv
HrtPuQ54Wm3RYicmrjtjS+Jxr5/zgjRKmxuk2CH42VL0c4CxSS+YTxVg2xOqjtSC
oc5xL86VaNDdcZ4MX8GzePeaO4gV92oXlP2LZiA9G53HpaDNZQLm3X03PWn20UqP
NriHgqHq9kHN9fcrHHCneIy4FmM4sHCPRgSfnuTTeZIOXmiVAekkwlsD2lVZMI2l
IEwoTbLh97UinNeNruunT5dZUDovHFnbogghcu66BJYxZ5HPTMWIbEuVLp/Simnb
kdyTJpso/gNhgxO65mJaJByNJhufR6oMAyy/tdG0ijWxi+dQ3iQzkFC8hROjMhFz
BfTqzs86qm5qIZl6CfuzTcpMVnYY04KPyszHajGUAkh+a2lRJow8SACi6BRQKBvM
D0QZesDDSx5+dEjmV1g6/dRxrCwYw/ER6Sowl44IuAJoc5W07z44fCV+TlQ37oFg
TiRM9CFSMzI9NAA1PRsBN863SbxL/S0PakxQLBcVm4PfEfQxmFIAVHftbPxhJ3Q4
cv6BRtdpV3Hkifjn0937nhctXcLZHaEyATzYk21fTrKhEVU9CtmlmDewcHuLMMKs
M2v33ElVGyjT/LRUCy5BYklq+zbTk1DEhEct+pP2QsD6K+eOPLFeyWoMQXYAW8Pg
cfMWei64a6yZtTpl0l5W3BedW5/WNkPGRx900CMIp+pNpvcqsp9O+hVwxKhJgNzJ
Mylbot48rn562nx4V6yQYugzg3GCwv+UJiur+dmqhYAmRAvBh93mDy5xzCZjN69B
pFKXIdiJlx2W5UC9jJG4pP3G6rCPco7lejbFQBJRdt9D2pOCwkIZsgb22442dOLS
iJAj4Nt1LdCNJiLdR7TKsrE19qeeaB81FC4bjthcpMI+chhipFAJzbg106qNmAao
E3Z/Q3fSIiCVEHuyeBTVhETxDVjkbekZWZCHn+FNsRtCowkKQ5TElwVxwfvtLR/w
9ALNHxhXtxrGBShvFj86wlCzDIwDx6HanY73l/E3kPNuJG892E97zpUgucSiA3Im
Fm1UGIo5XSbv5XRpFP+0s51y0QwwAHIP/4pTUYIUCJ23HTZvcVPEeaPoTHfYzBte
f1HdltPqrgGeyQc8kFWpSAD5nmYkRQ/uPEYXSmatUWmYoi4BNNE9Wixp5PCYtD7s
DWb2Ml+4o8Dubv39A6F5bYB6v336FL8B95ARlgDoJbhRqI/2a4QsniSn2k0f2xvt
DWr1jQukFG9EKPSgRHeOdoWLokTAWfDQAxMy1S3HOJg3M8YpPRSDZrM8Jj3d1o/4
KKdveb0HWU1+ZvqtdDQ3nPx9UGDSgzwsKjGSeTJzh3cZdBqY2zIlR8NrnRhisxEe
nYujs4vbwmYPIrrs0Jrf9UaRstpFLVFKWhpnGhjxgrwPU2796b9g3tRs2OhMSAK9
SMRAGbf7XxLVl8SduJ7uL0NtI6vGjk4iCQrp1MIpYYETTdjyP5rTwVx0FHjLBs06
AC6bcVdYpg2s9TAPx7K5hveFqqfVUouOcfnqOppFzfGx4DXb24TPsGm5NyR9sRUe
U1JNRs/vTpXxIiQY61q5hGQak1XMCsH13yKICC4jFaOrMyRxxKp/soD1iEvjxWKA
rE46DKO6vP1o0hts6cvEHbuQFauQtd7ap3xlAnx2NYlSU6p0bQDkp/ZoxUSladFW
Pc5a0WvuulIX4KriQplO0c4HyC3OHq9/NpL8x0hCbonv//9I3YsXzcE19WfnjUd4
ewrWfJGPBl5gb+2DN5DmAay+xOJ3lLGobJE0tNtlRIUIQnV3dYRSsFpKLo/C6dMn
g+XjTec7UfbGjRKj2+4cLgKtwfSxTLxLXan4GCM6Q8iOCx83mIRPIkRUO8Ac6FVX
1HKh8AMxqHrvRelmHl6IYb7J7Dd2i683X33QCL8m1gdWcIAwrkpmaCEQqnVwxvi5
luJMS77EmcS9VIAonxR+mXB7i7MF7LbpxSyfMpJJb3EWbB95Aigujb4stbH8MM6K
/POwmXHtKdR1qwR/F7x28X6T/yjm6FRfNh/84ulN7MtxATW2xVaDJ2b6FOy2OG0c
Vv39Ug3Fy+xVcbSrsaQQL9qwBe//iYyLJ9HrPRWLSCK6yX1+TCAUIxnIQrjntorj
unyEmksj292czE2n1pA+B8o0yfatxs7GDnDNfNpO8aSr9XWvT3oR+se8d4XtUfzE
NF+6GXM2DUN8tK8KyIpmqslw7flEjKPdeYDaoHp3lbkhlgCnhLtKzuI0XmK07rof
0BaxxG0ooKMgoaeTXnGfu1WmQUDtI0mlzNa2CPobpzZyc5/T+LYip7BierKBwXBS
yWkob0qQCuISiFIl8ChdqD89j+eK6Gk/bWOJqbpYenhYj1tE9Hfd2UjLLbZYpLED
mDLMY6kLRQCJqhqBwIJFOkf2oUjupWEkdP0A+cZ24ZlJ7AwXKWwqb2CZxrzI5yqm
gSVyyIhX2OTySYdQ2sGhMZOEzYNhQXwgx6zt1WoltKm6UQSr59EYRCb6ixdFmLU1
r0fE2ncMeCAQ0PVWvVZ/uCAn7znoF37CBlBUR7kYPIA6QDM8B1j8enZXhqeCkjwP
KY19ttHJR7Ll7qlHPRkQH3haubaeyzrtw2lddmWU2IMfFcCLGbMxV4ChKYJWYd6l
ffXlveK5N0du2MMLlov5rGRCPw9WCaDKSUHCZVWCcNi52/7akWi0az/YmcZsBQOz
/mOIUmFWNkkFLac1mX31441pxwsVNpnHfctJD+79dUCTSuXajS7hvrD9jXnKUH24
YxDkD0n7UdKaprvFLhD16cAvDK3az5NWkXn9sMVm86b0hshuW2KgNxwX2sa+0vV8
1N5xbVQwO/xQC6MFRM4FtpVXGkUbiKNDgIVdn+WCuCtZZCpWMj3E3TbcPziJbcsF
RNJtr12u2EPrNBo3aWCAL35jX+eW0FyHdhYYas3IDHWxDXarbHaNYrDybaK7ePik
OH2eOq3HxysBQcAVgJ39szLvV3HbvqnXvd5p69n4uwHexSfOb/f0z4+A1MLgveLL
d/5cC21WcbfVuM91H7fpskrVb3NLOacTSKvsRJ6Mtdzt7M/XvK/D2eO32etHSzWS
CRaTN3BDl5uxnLbkh9L+pjp6gQstLS1daRF8gjoOEFmoZKTl2B2whlh40Zba3qy9
rYk4bFgQZgyAUD8a7l14VlaVVVI0X27zL3iwneUyA8Kv6XSLLhRm0IqQDg621XXd
rOwRoQIMJWhSo76u+809ZygzrWS/+Qk8y74oZTq11di50Ey1Witw7GfDbwko6s43
ooWfQwBQoC0Pxzu43NVhUpr3yuoFj//j9gJZ+c94VrJIV4whhjtOwiFfw/xDHTAW
MheKTlKv5vjK/gNz3S1UIQ/UQj+VZf+8rMAPZLZjff7O+EoU4BPchMNOI095Cmao
pg3wCtqxlJ7BI0bkgCVAO1rXENdoFrPo4Wlc2ZPoKkl3piJsI9OCMbR6Xb5bA38r
n7EcFJ2tw771LFPr9TzYgokCeGhvDCtJ1moHCqVhy36U5cPm+tSULfqdxkuzqYFw
xYQhJv2WMG8bxLshfNtfRzCuynodkFWaBKwZNmhM5w65zinSMAjTgbg0g83hYrNL
DZ/fx+cX1vyuRJ3BKvQmLRXoLY+seW6QhiVp6s89r/loLebmv/PJJ48NIYy4bCp5
C0fTMJnz/FG+EFTgqWuq3+j3mbQQdMzZ6YCIvqZJySmt9keoVDJfn2Rx85FNXZS7
Mal7UY7sZbTOJDeHSu0ftI/dCoc0l8KGW5rc23f5JyKxaGl2iM9dPz49ZS3IJ5Tz
9fBw0ZsMGbsndyR9dx74qKi5hpjwQiswd8vLQZLq8hFk0Vi0R9WhG46As4RgpmOp
uzn3qZgx1nooR3qdZA5kEThYXmtEwv57JtSjj1l4mYgv3q99Tk0lHmpBAL99N0vG
Z4J9NtbT2Xi530OfiTY+cP+je6ufQrvdKcURo7KflIlONCki875/kf/j5CIh13dp
tDERP0BOS5G0Vu+4u/7bB1PDRF01IP3lQdo9poDWAw2htZmNs/hR8Spv0wXfcXxN
zUs+bMYCKgXwwmHPChmqyabFN6bLP0rKsZqkoMS0LWjyr41cOKVnKISg/+cJi8V3
R4X4AaXXK+0KrV71qKhgRPQcWQik/gzZNlpVuu23qtso8dxSWQpJpPg6c+wrwNO0
ZyzCeDdakod82dNeWHSdBw4NmcxLs+oJNNihjWlZ+WDl1jMJND6cWMnHSc8XvFJh
p3fhvZP98TPzbgv2FRFtxUNc8q3aU7DJsFeOKHpGOzd6lP4sLNCvtdP1VxDRFQQI
bVS67FaeaZg7GIvtt0C+AgwuOvgrCTGwYg8QzNN7G2B0JQ3gTHc2j3QwxXxbi8t8
y1O15TPFok1+uenrFYUsVxzgDSV0rTD9iz+CKTC2IgJ4nOli+Ohyn9YLIZ9a5ofx
d0QaSGFpYUe0LPodPoW7gDyD1OQp9WBbdf1xDGmrDS0DBw3Ra479lbBcpIuZw5Xh
hg37mDILVhMkHbcQ2KuCYx5DnCiLkcF8VDUwNVcAkgukZCsDcerSaqs/sxtqmntV
fFMK+5ddPUJ+orl6Zpz8qPS3NggacVpJ9xoacv+IMS8C/Zy/CrKlzwiDPbFgsQvn
1ZYnarTAZlbchcEGeu5lxkd8GOCwl+tV8HU1lA8Hc2ZHrQSZv6QmfvMB4AMW2+Tt
PB5WXlCxrlqcF1xOshNDQP8xU4i55Rk5Vf5O49fVNxeFVOUO1//MFrOwXMlXPMW6
4OjSYRXpcjRsorKbvTVRCvqNag0hPZsxibpn/70TMmRZCE15jTtdWRJ06oFR9D3k
0HpetYj4Q1z18jXn34D7QntsXBVG02RkTn2FQINV7kzzpGE+Mzx5EL7DrVNPKkQh
Bd85DwBYZIglvNTnXkAYQWYxSn3MjXr+YS8/SSRnMA6AeeznM1zxKXOOYvedFFpO
X5hEHjHpUwJ06FE3xbJbhNGFSnHjRpvK5lFy1UhCSUg=
`protect END_PROTECTED
