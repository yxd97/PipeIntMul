`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YDy50+lGEUNhsT9UE0s9y0oo1Z4ACPlLxwFtya9hYtZp937LDEJT4igJ2reqfUK
KGdVts0m/HdIvwrIfb56+ST/Z2yDlBIb2bi/03F07sTA1bq5Z7wxTOb2Em65E0bY
EABXlqUdPfOfwvTdBLuGFlZ6rP0tM/FFrOS8Igh6LoLzlnUteQVWJOqKOwwDN16A
W8/ozw71SIIfu4Ef+Jo/H6veHPNRam31jbYG/uToSPxEay1GU/Z1CanxgC9oL983
8Fgqs1a+8j4I6jQmyqwuEpdCoF6yUJKsYhrelOwtkkqYqRhizXmxApTA1elAJhCd
Tqd/Myylu5KyU4twJ3HCPEhYTckcSVWtUKXivoYyotl0upR6bbVHH4yLRz9PsJS5
kncZiBBSQ/cmeE5ITjDWkZ0S+QwL6TkZcb0vA0HJrhnmJ8KeFtPfdFOPUyVUQh44
`protect END_PROTECTED
