`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mal5OtxKs3RuvllqRj1KtQvHqbHO7BoEU0swb/ptknaTFqWqq9oTDmVpLLqV3Unn
+9N+P1Ep3zx2yLfETKdbnWmEjCr6cnMJn44JuPRQZFH30OhQTFWVf2Lh73afNCwE
XryA7R8gvu80+dxWTZC8e2ISP+5yIc+/yoMYzg1wh0ZPOd8mUrPyyhiMC0avvxHo
g0yM0edsKvDQI+AXO0IGYPOUUL3NT03G2ieJ9yoYNoAH83+Qa+iZqjF9te6LPxbU
f2xRnjp6ibgxV8VOUt96htiPLPLLrZk5oPGRW77E3Jqy5DcQpa/EWjBLuWXlk2Rp
ovM+Q7P8VmzBWiF1AG+MIP4YHllrSKR5kNjsqEHfA1goWXATTKHsqX5zJSmn/X7y
QjxHZBdbKmaQASX2K2QEBGydtgHjqz8S2caNN9T2ff8P3mDY+Wp46scqVgs3qy/E
OyS3DjFLE/+ehO93JbhPEFH7xND/MvkuAp/lW1DS2kQJdMxkMZX5g1XHLOjlyCwZ
+YK640mxDybqI/8i3IxqcCf95ediF2GnQiY6XUfhYHfE5NY5LncH34/Mlwp5bofE
oHq70qrXCNI2qq7IVHR1OJPLLmc1FIkoslZdMl08ULgWhZ34gkU4A3hbU/sMEMFu
VxIbQI2LUU3KUF9gox1X+pDsho6GThNq8kA7j4TEp770jGBzGEMVQqBppi2yVfiY
wDFRuqDuTqg5gA+7XkUlpo3wkHaJ46tkM1h60H93VbHR5EP6dp8353bclWSMroFJ
`protect END_PROTECTED
