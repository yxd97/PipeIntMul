`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOiWBE9+xym7YIvejPKha1il8E3uS1T2hElyoLBUJxRHSTlxR/8D7xO8wkc/HuwD
bwWmbAu7yz3QtrnGWFhzaElg2CL6TE48MlrclJ7k9k0jeAvsraZVMIuw6oiFhp+R
l0+cGnziYjVSYSNUGYHU7EW11FM6aTLrXTrKVOhjbQ2AYBduDJdGi/2xEnI5h8QJ
MCH9/ftYL5GOy9DBAnuk3wUa4MalTATgE5Eu3k4no4ZsuIiIAQAMD3OUdeh5tYwP
t78XaEsOKOP0J27qZQWBCPIaI1WcmJNq0SLg10tk6WhD11qXHqfxVYWHGibhjqq6
Lw1vel5xijfZgunGhHtuQQ==
`protect END_PROTECTED
