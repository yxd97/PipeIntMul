`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jAVRZBrMyBOuAjLHDdZ6diPUrw3qSMNpbsWjvJvfvMb8qFuSzUsO6hDgM7MadusU
5GnnR3gD26eCOkmE1eT/38JMaBMU0FU5dCRNfR3p8HTWPRa3KMJljAaKnTPu+yjQ
zJGDtA+PnU13zfJXoSH+pTdJZOzg4qyDqtFQsWVAXgE3hA2nbjbM5g8g7xMV2yvo
pmDOyML7mWUv3fVXu0+WOAqshvNEbFJ8hIbD3JsoZX7oTSIKIRI1fbqNqzhxQ2y3
S9+VVrSy5H+XA291ZG6Xag==
`protect END_PROTECTED
