`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LRssDDFa10X0YDjCyl8rLKJHXiaAfkOnHttXoaQIiekEoh/IZ2oyPCe9uLZIbaO
1M9q538hGZ/9kLbuB0IilJeUVB7k/8X0gSrvggpb8c6W5vvlfUGSNwCCV4Eikhjk
6kHG7x9H9QZaAb6/fgqnMUvnHPf7kwpqwV1oQEM6bVBB6l5JCOAxIPgQfQUGwXw1
7ZB4Pq2ZPLw385F589xgLefkp9H4nj5hvn1gSF6lDm/Oo5peH/roq8KdzQhYI5jh
r0Fi4cpjPRCSXxQgfdeYq8FJPh+g4zkstIMGi+vmNt9iA/lqUurjZP9Jt40M9YB5
wUwudLuFuToc4WTOI0vICw==
`protect END_PROTECTED
