`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2iPOlUNBKRJi/q4H7pZLJRBQEBcQixRVe83/jZuSlhO+9O6+x7DAvsR6PeSHoNBV
zPLfHaU//6RHFCvx247J0384zg05a4VLsqSYfyNw3PNs8+VyMoIu++gPHlTmXScE
ptKGNs9/eGuoma512IpyykATUOIk69Iq7+wDQBcL3QdYkgwsOAfs5WX+NHBzMaUc
H+20CtGhix+Hw0SltRTTcRR/8l2B2OgI29zxlCa8ChQ3Ijh9VpZdRjXMsxpKcIpV
dzKTtc4gc9djCPNXzTyJzH2hSKOUcQChlDIi0gj378byD6xhKCKWjvkH0TkuIFie
gVzCBHdw10IY3kDboKArxmPspLdrinaAl7DbymfAug/7peRdUc3p/Q8jfM3yaWXo
dSJc8ViDnK0ZsoHP7YTkvw==
`protect END_PROTECTED
