`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QqOADP1D/O/164+4T0ZMMmi3u0KOGBw6sEYF9/ldHQOSOiOSyrohMUv37ysQK/dc
qgWasA3R+Jjf8RF+L2C3xOJaUhzz3e4owun3Uy93cFa0T9ASs5q+xiEVp0R9FAIz
6TsEgikx06ynt8wlIrIVzz2+0Edq2UbhEu4bDDRYntMeM6uu7KF1axEDX06A66XF
21/MRbNML9omjoM473qUN0ccklNa1QQqYtWe0gIwHGdHmv38a2TiH+dvMVcHOOqC
PR4XfCwFZ3D7mqjURzUKnSZGB8pHl5ovLd5YhmD2S1UXIsYVhidCX6qWokqyqFlN
l4PKp480zBe3NpTk/5vPHPZm8No9YvBEDkcBow+V47Mjp4upK5XZJhoiX5aq/SOn
Y2FqbRgtKfWE0pIyfGzmlA2BX993SbiXabGg9hVd4MDyLu2c6dOp8S6gVgP3ziNW
rZOTN77S7sWja13EU62/iEicb82eHHH84sZyNMFo+hJpHTxF/kd/dJdEKD78QETZ
BBhSxJzw56qy6MP/rMHtES87Zuxo1Nh/TPp7Sg1jp8r+jGqgRP9QwGRV1pB8kRsz
lYsqkS5qw7y9b/T7kTL3z9NOIohN4DWyrgAMr2dmff7RFL4EGbeTrhoJhobWRfxJ
uuG3jNiHbnZsC8d2fM7lopp419WWpgv3jZkQ3MKTDILjUHVQvM6UGomE0T8Ueu91
XW3NaFeXu/MmIHAi8pV2FGUoGlAtrwfr/3huhMj9tzTuh4NOrt4Iy3kcu6j/Kymm
fcqIi6d19+BcRJHFhT56S3nTr11iGN4y0okDdcU4Np8KNs+g7ijDAygsLHEZsBc1
sL3Z7ZeiRPnUQbmzNMvHvoGHNIB/ZZZvpRSiUsBU2Yr6SfKPMU7jNHCfnHyVnuHe
DJbTgXHPSEFER8LkZFkRhA+Lx8viGpYO3/xSQbnctaye/irmIcyZYFjaz/jqs+yT
no146HuCiGJsJcztit0oEJGKgEa4ACUyPka4Y/KxE0DnBV1Y6p4NzqnzFW/GjEEo
k1Gx5IykcNGZrF1PhGKjKZX5C8xNQQ1PUdOf1FQWcVshhoN7mkEae5dZADgMaD2q
aib+FsWJ8bw20F2JSHCr8wWrVrN5mxAE1JyoQJ3r9wjm/w+2oyjP+tVmTtpzwIcE
LYZGDUnHhlbcrrBQukN3/aSo+JydE6iMZgc4wphwmOdsKkIgMXZLerNl1V/cLP9H
gCqE0+V7f+LDP4n1t3UFzCdWMbYGHZUXQkOqHTG8Idf5kV/fa059OmFzShho3b7W
N/z+IHvfW0iiey3iURASJl5FVExGZ7erB6ayKQKIv8Gn7RtObJqoQA3QKNUZVHAw
8jIcNWpWW5A5o+2kMeKuBnYhc2AFo8V0xaVXU6sehvE0Jn1Xn9dKnAgWqnkk5LqL
972gYneE9JuX8/WKCxJqbxxCh28evwdwAr5mEiLFYZtm1+mnQbAZAcIO2zBlsFpn
tvbDOqAGEkvFm4xuF5Phr4uZG761ezbqlZfobrse9n4MgwaoLckD9bKC1/csBEXY
YyNlpdmLn5zJ/ZTSShI8n06qTxJVx/30f6UT2icUwEVqcur0LJ+W9oa+cg0+tjZf
kYyOJd2VMC/sGSvgFWjccB/UyemuMVTUbOpHL1TbZLXV1MUFzdkRGwhbUBspEuFx
LJ/3xRlZeDLYpQc5snWSxq1VZjvS2A3JOqXmeEmKn5Jl7BlI6dYfFKih3CEomq2/
Q9BMyxaK+TRJlIlWJ9jGvC6tXJQzbPM/aosD1nw7KWQQw7m8cgum772ceDYUb24e
tyZJIdrWs5P9KK7QbdV3UwX4PlF3LH14cCkCk100NnsDTw3c0u57SQ/1/C2XC6yw
vaGZLr4CcCWR//UKTt3E7+ZOjYD0NqTfhbVJxQcA4GdSLuB9ZAPIvCJLuw/PdjnZ
b481yEQyQCV5gRPdJ1FkvGK7Ky8o2ruiXhVqxfsls1C+ZcdwmZuyndJEiiQQ53/V
//Q2aqNk6M8GCaVQaTtjAiQHXeLvP5iVbuPLxqx9OPVV0JXH6XPz4LJUece3C2H0
l4kfYB8MgGOOaMLB01Y+m8AYqkxc+dxetkoUo9DEualpSmvLi9yJYRQk/xLgCu/N
bASSAaL5us7BlXTR+4fzYH175o7RoNT8OuYoXOH5iI72wkkw4b+vQCChU1rX1EhG
mQ4K6v6gdbqpD+81jOYNRlJn715d6pkZ3nPkesVAteD6oTcyEkoHXRfrqr8klB6u
slb3+p1suClih/Il3S5mV4uiKv+FlHAscKpKi/8drHYhiSAENDgLeRVJZmNldGeo
Hl0mQAJDDxtlMuqmiK4AOSUb3bu8uuFTEkSJOwTg+68oOLEZZmPX9GLKpBLo4rC7
4vB8bhmXVz2FQhsxuQhf995VXN4COUW9uVXRzIj9LP0J6zCzto2xw6KYNlGcCOWA
DN0r+kW1KJIjy6E3EUGHQDQTtIhoAGrpx95DOi7r4qFU5Ee+m6zBKwJW0JdMWgFZ
o/wL8KDDjXQ0LVtx1Kh5VgiYtu5ppTysiAwxK98i5P4TOirZDwU5nt4OpDqcXz2g
RAZjDao1mVXQUxWo2M9lCXL1RiBZ+fCoBV2PHzguoLVVbErS36/ycxWUVF6qtAs8
zCYDekWo2LtnD2mXPOc1qaPbdtHsWJgrYA7gLaTrHNfAW4u4ZQQvwSMI2J/a5s8S
zyLf5NcWgx296ra/Fe0YJUXdATOtPjvbYEUxQK+RUlUCvWbUz/9eJWcm0BYgYQK6
uyFJVdHomVtaKY5JFsWWeRTPTYeFvmxZWCu+B+aTfUm2Uglu3WlAR98YKGt2CStR
dgKdpkkOOHsqaurUEqwqXwD/xvAGMv3PcuofFrR4nOdXkbfHzuWSkUfYHFDDbDvL
TYmoBT0ZK5C9SgmWPu2LJ6EBQ0Cm4QnqjBEslmydRN3bhkGzmgLvxKGGwubtBcZN
bPUukPBAv4oeVinGxk+1OPU4XQ7iyakc/CH2mVfWI4p9vnJbHgdGK/H2L3+P4yOc
8oAl7GEK6tEbDAsfFc4Bw07ErHmscklwCZUL5K87BB45fbftT1nqqyFpFASn5BkV
6vegQwexuhiIBi/lJQNViBxRjX0FtrvNCFTqZQP+rLR4i7w4zKRZQMiiZqfjpnJe
jo7a9J3nGhlsYTCMhX2MzVAQADzLG349p9uyG7TB7T7JeDnOSGzl0JrkpJkfCilD
8tB63SqXYUnCF68XAQh+sFLapSg00HxhS5LXh/rP5g69PVtEy4tIRJk/1MKHvtfs
P03Fr8vJRG9Yzy9rjkwN4HOmoX7Q4cFatCK/1dSW2Nt57XQaIoJsaE16lyfFQQvp
Fp3mf5Ab3Ozeaw+jVx1Xk/Zi4OQ3ej2trck7YMKnlFjrUvILjlN60K603+NZFs8U
8gJd3fovwHqonwAel1hu4IlB0LvvQE2NZg2WSwA0I3ec8ldQIb/FRhqqa/ltgdRD
qep05ES5GCBJL67fs9XWNQs1ViXYpZDEq1I/wWhNQZdqs33yJO75vNDTFsHDHqvk
q0oo4R0o+HR2SAHe0sglez7H8wCdkhjFhf9NVaFxUa4KUTxUEstk+Ai0tN9+FQF7
gWcJY/kB2W+CtXpyyHUW/5OnaxxjjPu8fEp4Y5LG+6oi9ejzC9fgke56EfdqpBXL
iXvk89libHjBxS4VZpFjFaWKUdCQmE1m5nNB6Ct+Vz3fDyM5jH9/fSliDsZfzfPp
v1y58UKk9IYdHI/CnDsba4yR/j2PrgoX3tsAoja1S8p4x77b79CApdDuPlkROFi1
PzfTcMTcFxYMddNmW3fR5NA3z1CdR0ICiJjU6lgXEj7UKkdn9IBLa2C/Bh539rZf
zpBkZEi6FJppoTIm8//3ox16ZFCJ4qRoNoLWoMYWuMwMeVTKfqLBJ4k55mp83LBz
DwS0729/7vN2gkaSjO2HotUqsr4DLLHYQXo/OoNRkpmNRnuVVcyas3smE/c1FLvH
LYe1U45KnPaeEIbxWdroEYJnPwXbUHg2092BNSpXG/fPzCknggcBcW1bkTERnbi8
QeAh4bB3INhVVxHYEvpcYNt1dfmTtv9R9mHnKX5IAZ5iMWA3JhfoE0FJqgwjNPk5
Prwp8BjuY5NcGyFiSu5LzlC1unWw2r2Sf0D1CuRxIuyDpAXPo+mvf//KTbfoVE/Z
c7zaj+gsKSji1J0reiFtnWDUrnP2tE73O21f98eHtzVr5fr3fdN/KOdrvCitJAGn
zl6XJxOqt2cTH8nlsBdGjo9CHJcMLOYQOg3BwUbKVhNgZYUp3ShIf+cS5Qkg+HkI
/okIb9Y5tFJPB4wgnkLOr7kTUqTS0jNbEJNQIoX8qmgbWaCfYkGWFt+4i8LwqpGY
acSq1iAlE6Fi82YHl+RfzS2NexOL6K4dE4oHZpiOqwJclBW+0GM84F9//TcgJ+/T
nrNgrcwtMv0QobLxTEseqRetDTa3ln8MEx2Jsffi99st9mihinbdvTYnD8cLbBgu
K0yqtuXjnfJoDi52LNW/geBU4rN3zFinnxmXdG4dhiGn785Gs8E/noOtTzlMhGCO
Ln7/mu4hnUf7heo7JR5+sOaRvF5F5pnC/gjjQAJMaTSUUrWMADmEdeDusp5FP/A2
/ujoSQOPaJ231uNcTJQjVNFTiVOyKgswFbeX5iPR5u+5mb3SYSOUo9k7ztUt103K
/82mIqLWSqrsFdeZyXbTQ7C5B/ZINxMCsmuYQVFgd4AjQjWMI7Lz96W+rV99sZ1u
NMTQM694gl5rt/nBe6Mvld2a37Bui93bN7j/R+Veizl+lFgOAz0SRPdNSi0Hl5Gg
WRvYbU80ibUC2UOmCA3kLYJAMmGCcRF3s4EBblWPGeohwrCxi/msofkTK78UwQVs
1T4UMVBUTpv/BSPK3QLdoYEQLmbWYAf2kr+ONp/Vba4287zlFfNxEY9DZ669YskG
95moy/2CtUCVhuzLmVnm8zaXNr6y45zzW4XCE1As4pls9y9ZsfUrVJMDIxXThJMb
AIncvhUH/uz9aLZws2leaRFrZznO+88JMvcxnW85MvsL1JurG9WNU+RQyqQJR3d5
5iew/ou/W8CkFkMhko02NjQzoq6eVpM/h+ITpBmXAGnqdd6FJvN6Q+/l0/hSPGR8
Q7Na3Dzkl7U5hoPpwk7SF6+5A3sXBWlmdnx0NaR23//ZJeNgDsTpcW/5zF1iDcpK
jFlRr6NjY92kRD0S9hDCgCqQLadxkmxOAQ9PyPODwUyMUL1I+A3N4cktDV4ZqGeZ
quoKr9aM2pPAzA8pImfX+JnGGWrsOiS/VlHqufJrImjYwBE3d/vbuJfK7hSnZaXf
fXGgv9J81fgelGKSCinBRm6rSNzhqfL0X4paADxJjWZ8Slab30BeZY9FbSQuXLCu
SRO5zwkbqcf5QkpAdAJ2mECjTVHA9HHOOftLuKtyGkMqdCPaRTJ2GSsdaQ779lXQ
3kbv8r4uMw2iHuaO0APOVQ0pkgrM0QXDMOqCTnFzBNNWHbA7AJsEAP0d9bg2LhjC
9Z+7hnZzr6Gt+wpGh8YTJRMIlwGTSuvRaRcbLnMdmIXyIGk45C9JhkTfLRNLIKa7
kO4gXi2O9DPq6uv+yGNeKFnc8HDN3ndxzwsDQjBuxlJPA2XhW5KmElWfPkFxqjtj
Fi+JRhQS/QR0KL8G2TmR+Fiz8XSkb1aUx7YNJ32+nCjYkToZWt2vSLSwnHgnPzq7
0nHazK4VHwTD0vnlvf1amGO9p3Q6uLrMn/FG5viwVp9HOdeCRQ5BYqsQvP1UK7Ko
DEFh/ZAb80fF7F/VKtfT8MCXFw6+wB/yq4WJDDZWorX65dsN9C5bvrVCvKgM+z1Y
P5DF1pgxa4Y0Kw+kyZ27ZDnYsEQjQ8ZG3BXp/KJJzYoyKFRkP3qZPC5u41K1FXV8
sguO25ph2IuthwguOoAvPxrJ4U5oGtVOHjHMsVhuQiwC6KKVvi/AUuy+GTev/hfv
QEjk8eS4bP1qLNlFmir4i/oQnTzMnhNYKTiW2PVl+LHlIN1THD2c2UZ5F3PClDPo
cbYvgUvtdVD5iNiN1ZhIW4N+SXrAC/eJr0cUBvdHoaTx+TUJytUjxm16yKkJR0a2
jI022eYyPzN/LIfZhIBlXBpFKctNdsqePoiwR1+b3vndFphOcA2hN13j792xDg08
Lw4sj1ejq/6w1Zoyi+Ep8pVQ2KLpC43OhGYsCCbuSqw4y0ITvqCr3YsJXZwecfVC
JsJ6yDd8bK9ajRy28DRUPp1Cv9Z1TdvPB/BJ6LrmgsbhPrhJlD27Qfpn1bVNJjv+
IFj0aS/bvIF7tIhRJ67IDA==
`protect END_PROTECTED
