`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvpB9jzBYtbFvSCmokbVa4VbMOv7aoryrujPQsxLpsjvUn2x7nGwOHUDWaS71plF
RcFXTgHmJ6TLuCTlM4BwWxnppNBj2S5vnEUB3oQ1TWOF8Cgd0dIkudXuUJZ//OYv
qpVkroU7BPpWO+71f4M5DA==
`protect END_PROTECTED
