`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfTjlkAMEPMgHtMd+9v344hjhAdlrKakFmFgsytS5OeD90PDQ2l0wxPfUX08cQ8L
91/SLmOGmeXLBm8JiGZg8I/h0VqxeKVJ7qW/HIDUQKKTzt4pledHGYZSIEs6CG6N
ECeKa/d5+iV6T78HRJvLJoeVZ3lB5rKVLDp9tIxeARLNxmoQBgN5Gwa54gHHkd1g
7rjMnxsU5KWSvaITxdzhT3ijFvPZXoPZU1+o0PSSjpd68x9MSTYWI36f0v/roiSL
Xc3UrSGiYcjhPP02Bj6ZovbJDg7YTRLN329/VXul2q46l/CuBGMsovE4jN8H5f1c
wv7cgVThVMU/AI6GvnEvR86mH4nZqzu4vog9SuQbrnyEteneb1pviGqq8a1J20VR
CVddlyKRZunEYaexVLG1uzpsEPIMnpWZSDvWksxlJk0=
`protect END_PROTECTED
