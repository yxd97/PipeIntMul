`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yAh3yRgfjicNhZ6F1ob7tLnXoO5w6dNKqvYAfNtFH1S37w4B1MwNATjAr24xWTPL
jPyQaSiQzNeCzxY1i4deJtJ1NJABLySaZFEryaL7P8Y09SaQ2WEuNJC1FX3ubGZL
K77E0zdpDn7hp+1jgWGQZJi18Ml34oIsyElOMwY3m9kSeoUVPxaZw+Gt8TRTQJVZ
dkvOOB03OMtMZlNgP+otzIaE9G6vWLw9gLG96kz2TKM35CfE/MgqxZ6RlYFJvmet
FzvPUFkp0H2YiIcobbub/fvmFc5mZDaDlreCiyN3mhRdUFLvKHU/CMykn6LVXNcR
uUqIwjs0CidmbMfN8qr5MICcZU5FHjvlx6eUnVBD8DC9AxQfrt05QNykMw/+pUUL
AxTQESNUfZg53w4J+iWSDqmEy39KMp3f6UVuJjO+D/27rTx8OVkBy6h8bIktLqnK
+m9OuLWJeVNI6xkOJaFqY0p9ohjJflNuIZTngABmFmdMtmKGbILOFZNj2h8I2Otl
25BQTs+5jrGNmMJg29J2C2dGDnVeQW1Ox/JvAgVlKoJxZhW6livc23DHBDz52pkp
8x+PAnHLrbhbAIrl499ehsnDWcl6w91vFaQutX4NOECu+6V/Lzy+NyWAQ8oeDSam
ydWFCA9MtPirF00xjW6lOPY9CmdDmeHLpZ0p5ePWkNgyVwCimD3od7uEp9DOzXpI
BTGhoqAcEvXABtQyHcDnI3OQ5B6I+h5w2CdgRnAkznSpB2ZAkG8NC/tNZL3EyiLd
cUW4yTPTbyp1w3AGRSy22O1fIwFW6B2ra+qtGXRoyp+45uReNTvPQTnBCGnk5WKo
Suv4GfwVP2ilvQwF4mGTXHe5C0CcDM9vs+nq7f0QOnOs7gjLoYvXXXLVP/WIC+wR
+g9y7ck7Heu8fD2VtjU3D/YKVfYlrbrbW8QkUWGu64cuSIxOPYltD3Z0wCuAxH1+
s/DYzUpV4ro4JOtTi2pij8IAjbpBorscoBSUsIXgCoD2HnuGt8WzmOjmUhl0pCzO
G3tnw0ggLiJlguA5eFwfB2NjEwKjtQIoVOSM88dqNwZsy53+9lugV3r8wgjSxN61
cTGXaq+sNYO2/JRMteFF+jkVn2b6G7hloR+UIpkRmHSQ1yeRwjtv+oSx5DkfdHiq
Omivsfuw8VHB6s0jmqE5YTu2lIVjlcYdy//byzilig/5SdoAd8Ak0RPXETQB44SC
jnpFcgmOjYbxbGQBWSAe8Txp/EP6lXWo/VQo162MW0YT4ViEOCM/9yYOZiSOjJiA
5fWu/ucCv42b/UE2LoElvdP5fba/UbPKyw9bzMyJ/OO4rJp8wsfn/PXz+EOeL0ni
Cr4iqh0cPFZpP6L4n6x10hgKvJMPVVS92qTt6WGbHz3mheuvtUGn9SKmk1FWQbY9
7M5pKLtN31t2unUV+5jL58xoUenRifWHrJGMPchgFAfUkfRU4UEIpGBSqy3GVOgL
S01BHrlvLo9ZLG8C381Xl8AkHLtTzieGyq6fQ8SKlSaqo0qZ5iqbbnrxB83vdapt
puf/ps21MneJNf2SwRSaZZ3rfnhu3eGF8QYqnesNrv9LjABffd5uQssuSIgPbJ7y
bOYhaa5GTkfiDFmF9YFcL/tzas0pc4rKjpLLXsHpfH3f0/eGJjoo6My6/T5AIYkb
IPnFFCn+LQiTCvoCAoLRhdhGKBv4a3WeoFiel5HhXrdYg0c11MLEpg3kQlPmhDxW
kSQ+AiL2CjC5cu4xRnAOVubW9x4GIUC5tJ+4U2vhiwcwuTFChztzRM/SZmJJoGt0
zrDTZZTltuMeR4KTzBTfzNbA9OzGyOARIfGBg0cJ6KdALPPkJRiQg5Z3jCJu9GNR
zkUwINPnEsOfJQePWeBYCoS9wyoN7tJdvqLuPb2vfwXsWmeP3WKkdz9khrhcZxwt
FGBASkQoDQF6SG07rmnw4Q==
`protect END_PROTECTED
