`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1gC78fmtfkIzWzgVUwBb4vURwhlFEL2Zw+rQrmXIGQrJG5kCDnr1dIfcPGqNl50l
uqmy7FBPx7306z42PFos76AYqYjXESCv+QNmiv0W4/D4JtwWkrJMsSU51zxM9FF9
oa/hA3RJlM5NSLoDdPttMVJ8F3jJb7iiLVVsDFk/Bi4LwmgY6cV3Oq1xPPHfJHU6
kphKPOg+ltsIu1VNGt0WLzaHRmDIULvu1wQeWomMEF4eYe22D6GBXaPMF9FoiSjs
1OQnXAhPXzAELwh3QBGN3MATbF+Z12xCrXxZ+7ve/4IMCN7CKqkFHgS4I8lab6Yx
mhmy6wVZU0liS3mO7CKNiS7yWSiiXtEZbzKpSESOkJhZCXu/V4k/OjLKvRANSa10
Zybr1RwRBVgHpGvp8G5zmoCqKplRLHtFP4ns9HmYV/27hnpjhMVHWrwZDwWAeQBL
byzLVkBHWi7QfeTScTd5QRQNthrcOQ0KAcPcoNj2GePVWwaJ2s1RqhuyIXG0Or6v
S3rvRRw7iVqGxzDkQgj+rVvG58EBE9fNZ/zYGE5oFhqASp4p4VAUZvbsDhRhg48a
aP4CDQ8DkPSdJD8yoDHfARhqGY9Zt0TcfAp47z8BMXzFQmg5HPTKJvIXdhECKj2r
g/MdxcnUXWHHodrk4gC8jyaLwftOEKDP2UE4Ofx14rW89i77f0kbl/ACzUokYGZI
PuME5VplJlszOMfIKCbSbVbAOSXkg9/TojP8rj+RGz3t9lOt3R7Coq7DTq0/cLf8
`protect END_PROTECTED
