`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4RBCSbN0iNOEJ/SEGRQqmwpmqlfe2trojKkmqu5DDhmQnGYGlAzg+P2HUNEJoWWK
xhUFoWPVOD71iNf8siHLtyppCt/pRZl31guJi9md2cCWzfRT1Famuw/cV9m2HjIa
nAHxOenzFPhPNNW7ZF3zrLPfVaDrwYuZD55iT6gDFMvYPDmtfIUAWnHjrIX3Kbae
InEGTJLwfXpE44jg4IM5MkE226/6tPSousLJlys1uuLo0PoxnUEC+FwVTZcB0elX
Dyf4aTLW8Uaj+o4/QRW1TS6RKQWWzHYq13/7QFqbU1fPmU5F9atPZPGdPEqMQX56
xeO82gq6WnPdBLYuGA3aIw3L9Tw3ZkSgOuj4VFFhD1aArH4kqP4Cu87Pk3m3+jIY
Rowej7wZeWi5vo0SA3GoSReMcrQB2Zx7LPKbqkZ3QLjhVs13BeKKcSS8BjDPOEGv
VuA7VCY/sVfYx7FCpvSMQ8I2GQzNLn7Gzg7tUaCb0CKdFqDeI7iSu7vp/lvm8xj7
UpQTXBJ6oz7KfQiWrjZyPhCeFaTLySYsZJfht1amqLhzgH8sJ4qoqzF1wY9E7XW4
ToAOF0uFd3y77UwYm3p2iVCLY64g/ui8Ngh5IHsQmm0252yJxmb1oW8VLsVt0b/L
cSdIjiQnHNPTc65t+hGc5in3fLQO6+ZFI6Yj+BUl60N1NNuRwhGZcgPCVkAftMCE
LPoRlxaeUSEg9ajEvU3Cp4L6YG1PnguVYE1cjqrUovXQxKOOliLmFUwKybPe5aap
taHT2wxVKnXmQ89uxx26OmPTT1oRG3aUdA3NIEH9jJnV1HAYY52eMgJBu+7QPfAM
Nfw7eTTjHiYGtyFxZRSSLjUMO8znGTRireMRNpxRhlRLCDA/CtYaq01yQdc9N+5M
QDPH7M6fhoJscfQ8sf+rRzQNBNz9sUR2DyDk0cfZd/tlR7iVRksEeAdxL2Z5u27N
STIedN3QyXVgNmqseorIugYvGJcQlTAhinKX/hn2mBe0leSRMGpiXpYviAOzdLXA
57xyUfpzyNll9PBtKHgR7qIkDNNBZZ/AwZUstIlRNGuUcaWTr7l5H+iXzvYZ1+r1
G1gSFJeIshGV6oZ2IYBU91+3/eOZmjYRNOPywENxoDT7MP+cmy9MXEZHjDHTeE82
lAEmpidaSqWbOtxCfkdN7DRPDlwq3lg1cv66FequDRWv2nC+piT2itxjRIB0pKae
WrT0DXYz18+SzCVsU6uI04sO8yjLnEIXTtbh+lReHVzKd7qcsGb+GxuUjR7TmWvu
GGFgx1bcXmrAs+qjZB6PnqmnVV/rQIT6AxkehGS/Ol920rVxjmi0hfGSGhwdfPcH
LSsFgc4Hl2Y0CbMmhCLPyjBryqnqmfa4rpbH1z/qmkDKSEb/d27fdtS2AOHqVXaA
wEEZYUH9rHeNWI55Qxb46Gnj9xm+vGXgYB2JnZSm3BzgAwzX4v5djy8NrujjDv9Z
p4zEAAbsEIxzCGazwko8J8YYK8cxJ5x6lexpUvTQiHCXKQLgD1nzWwavT5OxhHQ9
VWMeA1UfvKC718pStBlUM1nW8/yQdfQnKvHYLPIJQi4xcCMWOZqQ4eVzQL4I9C/5
dOFHL6mr93U8m0dY4IRYzeNkz/QYJPhSW+DMQxpgADHXz4VioGYBIyg47BmvGfE1
pcQKqdGae/oTESt1wp7fkXnti5PQX/9ipvTnBwrgU0oozD2oTXOjcwI1wW2D1yFI
4Y03TtS4EcVUyUmAYPIpbTr/VDHLAS9lKvgFwK1Aa5PEdNC363iPQol4GN2ZD03d
iGCkESzbkM/QiY37MAMGSBT/eF9ULCEQza7kbxDnmsEMflz9prdOj+W4Bx5l/rMy
OvNhLWnknB6QtHzik4ozGtYk7EjcmrE3TrpLGjPvpPOjWTT+2J3EIDZjk9wkVwYa
F2BRcAwDcH0NNxtoYqrORDJoZCBp3uOgT0s0EV/00WCat3lJm+8yxEcTM66FSI1q
Kkxr7MJEMuTYwBlCIDkVY9SKmoVjVVcFf92zdgcP8K0NTnoXK/gk1xD7iyT2Ga3S
dOFX2FvuBcE/QVxGqBAUZam4SIzF29oSc1XV3k5Eh9vOaZM2pKZSK8Ibncupy8yW
4q008Wwrt9bGAgDDfDThR7MDtRlyn+9b3sc9NYVEppsbnFj2XUulDj+qL4WInQb+
7aW/u6RVaq3PEm2PDFZMTouchKbS4A1IKUH+Tf91yhTC0vRkRZFQQSFX/asG+vje
+Jm3PdQBnQxlpZD8S/eFFSf5yOccLBdJSH+VNsUmFcUog5bvicLHgSC7pRa1QQFK
cGwEmw47hJrvRB46F8LEpn0hilcSivjSNzC2dDyDO8sT/6BFKRViirSwbcz9t/mi
2LCvQdtI8P2vzvjGXrp1QS1+xaK+zNjnny2DJYMIA53Hkpw0gzr66oWnZQb5qw7O
b4BsjQkwY9CCLxWIxjhNkmbeagpwhuz28NMMXRErsaSvYiHZPnSNgQKzmW6lnQe9
qLTsyC5pOwbqoPSu8leS3CnyWMFuic0L40o37xe2osTz8dm5r4PMOlhYbxSzC20p
egpbBKCbTrICxgfxzU4xoLRTkSI1Nxmcg3pMJDTzBsbzbD4rnYUSyT79/HSogzU7
6y7Rh7sQkpUCZs83/U6HGeIHp4mEuoERisiTDPct2rRy4h/on8fuxM64tJfu+inO
PluKSLamXm/BKsWik+7KExYodbzmH4LLHFITIlZzzV/8VJJtOUPUc9ULJbu6BYfz
RaudNAZs1XhAgVENPFPtJeZ6ejkgYzYIXnVYrniSVDjYvt/FAoeM/eqojzKCzhYB
bbtr1VEEqgPqSMC+dJtkt90x9Y6FacrB79+a7xSTjp0rRWtMQGafMfGnAQVFuLGS
Xmeo0JEqyF59gKwlbVXi3v9Kb7AJanLdMqTcONRGu+EU1+i/tDuatvHytO4zxnbE
JIQTCl1OjFvyathVfO/o1+qZP2ARHKIsKiSH/NAKxY+V8ZY5L5wek/1agpkBE3QG
CYsHF7yPYDwTc66WgqCj/S0jRkrRqcfhyXOfx+Vsmppz4khSO7Fya3RJWvBk0yV5
`protect END_PROTECTED
