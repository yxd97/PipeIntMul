`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4oNoIfiKtlUv/ZcfGqnkV+CNrFL8s3AzNemg4BOiBkv3NDxKgKKAPXUJgbFTR08t
/aIRks7ma30U4bmc1dQAbJqUp9+AhiqGOjTZGY7o2CdXCfGjkKjRD1MDpUI7dHeM
UuzNJuMyBpVf1EHb5DvsvNg3azvbxme6tuXiGbTMqECzTYMPMDb2gCujrIOvKOn9
aDo5nddjBE7iNC735FWbDG82AhfYIlRmniTdLgsl5rxz4oTqiFcUwmd03xNNo4UU
GCH1P+6N6NP0x5tMvY4KpVTcAC47bIEENrpYgM7a99B7ghVDWKFF8SuDXoQAPoQe
UNr5HSm7BTqiqj+AqIdIy3sYsbylxNTZV7LFRIimPlXO9aLjXxbvZWTE24gdr01p
vnKfEW0GJ2ChzHYUk6Z+BdT74ij5pfgEadPvTvNI2kkkcGbErHimmA8LYZqFvSdE
E1hkg+vGxDYcappbMVuWuCEkeos1hJjv0CP6F2FHIt7WZbKwaYQdx/0mvEHElzJ0
KLezJXaDF23P2x334nzCBeyELTvccbM/F7YC3mmRax1J3+Anwe5w8pJBUBn0do9W
S+qFXzrH4fIWsAiIuGID9Q==
`protect END_PROTECTED
