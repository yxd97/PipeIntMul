`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TwR6Cfyz6iYqvWfa/GWttrHHSwyuev4RlyIiZZdwUkuaAHLxV+CtMgW1bRL6g9+v
Br5q77AEquedeLB6uIGroXuiOCgI/BqDqbmvu9zn1u9+BbduY2r6ceWxCF0vX5Xf
VAWLxYPXHSezqGKTnv3u+jNSvaJuWohh+mSwxRWhGlWDBVtIhPq4me3nQ21Ayzpq
D78yjvqO8enJm2mUDtsnKVFx9xPFZujh4MJrneJmTzHPJdrlYXR4rGKKMt+/GOJ+
BBSJryuDU/9Fx6W02vVXq0JFvr3oIcZrN+rXMd/KC27api37QZoL9h+y/YlyxZFR
Qogdu2VgCMMXJcaj5qqpK4tRN1//aCBXr7jaa+9t9du4xqBtVDm0jvFUNJZI5MFS
Ozm5x+o0V8wxIyxQIWOQIgcollBN6m1lmVi3Co78/gdOaudsay9bHc2riDAgBGqE
QMcfhMNUD2+ZrjFTyQ3G5Q==
`protect END_PROTECTED
