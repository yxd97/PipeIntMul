`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qDxvx1wcxwt3aQw2dnR0Hb3cKd/iTuvcoKkPXlCmtYb7fdNjsDkIKSh/5UVKrzQW
rYVtnQovFG0gDEBgEj1UoC6L+SRv+T0Z/lD1l8NXiEJ/sTJoRM3JqMRqna2085oS
80zpvl79bV+aEPY6g3S1zCEhjyjksn56IL43ZuGfI81SzhVrXZefVCD7/s9S61A8
tnFtE3djBjxq1Aun9woSMeMTJFNsWfbEQLQQ+EWMFS2Tgd9vsWPhAanIR+Q+uvpq
j1dX9FKeCQ9VhLxJAnJ5Ss52lrP4owexDzi8RtKusio=
`protect END_PROTECTED
