`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B2mHSIY3KklrlH9sIQ7avPPfue9BTSgZs7ll1Kjs3192as6IPRrH7c5K4c3Ncn8X
B7TXhTzpMmOu4SuACkxf79KgGolulwWMc7jj3IONJyGjZk0cG95rjGAAxQHgpXsY
p36/2xj/GUkaYklHlm7qbGXogPGC/MrFYVL14Bu3IBpJTYx2WXWvMt6QCQPnW8TS
pW588uTR9B3oi0USSj0/IUgaqDjfmIlg5la+Ou49K5WSK45ugvsar0VYK7dmcFkN
Q2vQN675IQfVPiwagFEVfYCaaw+BZWzhym/m4DshQGUsJEzotIWJPCdA6TEh42Bu
1gARzTKt4naoGCHsJAl2QkJi7peZSgTNZ4+9Ji9/vLXygQ8UdZLba6q0cwCWztWe
2Ym+zEjAQkcu6yH285o8FN8pwNNlW0AywEYpiMxtpMNbXa2LJsjodB0DZTp4FE0D
NiaCiyzmRKrROmzemHI2Ze6EUx7kmHasSs86G+Ouzojnkzzu3HTYczpe+9DLkBX0
`protect END_PROTECTED
