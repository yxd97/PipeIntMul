`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oVD+wAJLbdGM/t8GFUuAckf4VhJn+oV37DzPBmyk/TvVfqqiG4pIdhF6GMTan8pJ
WaT3XSpVIhHuWeSjt2jIu0LfUyVQ+Q9mrAIl+0r2yvtdvqm9xl4Inl4niyhGe2to
I1PjGqLoimynPvkJ/mm5ruI4HeS5VdI5n9MQC4Rm2s7KDKa7jTLSMm8pfPp232+S
ECyDIc4stOMrcdtalN5IBn1UPStHWHUpATrOaDQZ5WZtaNPv2ZuYpADDizTT2biz
OefXiQHdw+6CEmq4NwxbcjHtURMTfq5Uv43N6CXN/NcoHBWsSdar2AVPI05DT1YJ
fYfDW5GHBwKDTJaKepw8/A0FIOnedvtTufTOL3+bUGHQRWCgn3CIGOozMoVyH+JB
/bEZpP0i3j8EejC8ri8rXUjl/brpltZkimqZgBNmmbIRCv4IEuDERqXzI+boSesq
kpSRpyRdanFY5r6Fb9AcRpkUR31P8HHz21XE3kK0KJ5+yHwr0ihk+kKrAXwUoj5g
taZTzJ0DqCVTLgAJRRSGjLJ8XxzncF3DToGzOkzxaAFF99RGemufhbq2j/geV47A
6SPyPapGv47AbrP0ibIH9gErXPasOzX6H8Xy3rHtkDqV/sehF6WvubQYvLp6qcjL
pJTd3XNpa+fZEm/7Lhu7fZkS4FWlKhtAowlh/KCrIr7/jW7H2aYBYX5+xEVWOqNl
5+sgFLXGoOf8R0dj9IorWEW2haT83DGD+Dc7rP9KIBtE7iVTxUtvitTwQgMWE2Ly
fXV/OzKzmBdDVLORMRnPQh+E09yvhBrMyl9bqb5qBL4oiMwyx9PieNncLaLiuKNL
WsBLs2qxzEm/p0stRgKnGrvwXZ+kB+QDW0UaH+fbEsZRXfZ/mpqIgu9XlhI7y/GE
QWIKdtMPtn2nKK4KErdBN3FoN7YpZpyjIDynFt1BBBepO2iEkKGEvCZSPDB7umfz
u3IfrM1knW63oDJyosegLqLyb0Rr+QctgaKhfiQ2V94pmSmSgpHLB3fHPNb9Lgcq
lXUybCXjNdA1KUPNswUqEob7CILx6w2wkTf7jtZ4rbMg/goLtXY7S1gte9PkdQTS
5S0ZZFEi1DWwPDNs7Rfk92wrE/DIv75tpAPH+glZKnVEuErzQfqcaylbR4kA+UrI
78wGqP2nB4OjzyfdTOnD5PmCWgznppQf8g2mzKq/oOd7Lz5hRSmYtr8bdd47viTV
vi2F6CkHydoM8TFC73tnoGH1wZ5q2nAAY1Jk8hXSPMD6paIeazniLq3vybYYD0qo
`protect END_PROTECTED
