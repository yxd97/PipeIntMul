`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/lkgDRQxi06pAgRk4WwOwQ7btnTX0xjtqG8gNQ09aEY6+Wi+ic3MspdSMNUnbGKn
bfnjPziUVKJqJjZETc0dodeY1pkMnRCsWsXbJyVsscHt70yxsW9uGZuqqNE9Rs0i
KTJUoMwO8nB44RpmbKEk2Se+hxT5VlC2rm2xCuUgz/hgdTlwebMx5nV+sMODRefd
O13n7MrLpOxc3y8PH1Vovu/4wedFuymp9Mk8akVrgeIcvROkjX2W0EKcw4iR1cxB
TKRw15+8ss+SVngEGteVpW7Hs2AigkzrqQlesm53GbAL0BFtVz3ljJlKaMtWriyt
qesXVC151JMIAaENSnz7L+Vb9Y5LDjFOPZJTBXy5tO/897vnjWkNQTNGqf1AQX41
h2+vl+phZ4zI7ut7qtj8yGFbrRXEwAIjCsHEAu+V0Wc=
`protect END_PROTECTED
