`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fAS89UiTcSt5zHBNnBeg2WPby7xW6SNhOxaAdfxI1DX6tWf74py8NT7Bo5/AE5mJ
FuMImvqbf47eER3/jXAWHvnkaDwKvtjxE8IFUtiUlITvoSojDDzOC2VBtC5GyR2m
5C7p7W3KmZ0IQ8IjhUEuEy+tL5gN9zawJ3of3u1Nl1P42vCVxCrVTv23xgrovyiQ
8crP+q7lkru9mY41PhXbkl0ngtf8bZqxtV37nKVudKaDvAqNGC+ZtgeFa3QK4nBf
gIDf9MZeXiOzjhn54BSlDeLHi8BlFKfLsqPkDQFHK/XI4IInjl8CNKNejV32rkMK
Q9WsvTkfdt800wWKZIsGLs3rbLlc1rsz6E/sDlwyjmE0c8tIGgQIfg7rQ9RzeOS7
15KAmFKfO++bPeRVz7FavY09VkgQZvjkZXBS2reGSnwnHyLICFwQgOoTINz5EqhR
x5l29hE2AsLJiZfZ5VVtXWJ9mCcRVE9hm/ey+MwW19ha+UHg5lG5cukXEwRINmt2
JRe1WegYoneaVKnkkvlMZ8yNWW8JrqTRFoXdydnnSuNrqo8I6C0yVC9Hf6f8zAxo
W06LLnHqLhecUp+d4HwjuIYhJmCftMkvtnfQpz84FvNGQdR1h8oJRz574d6uLJ5Q
Amzsczofq12igjiVKwKIsOvdxT0HKBVW/VQit6Ghvu2xN5BE+KLjLPwz5GC7KLR4
GbVJWoaCN/Sa2MCUnMcphvWeBGI+LznMZHg93GNA9lpiLD5/DUjqr8RMIroLBtDh
56rUmAsOpzEGBxj73aklGdRwxSv4wipXkiRGv1V+/k2eN4/SU+uBeZMIrO5iS7R4
yJE5+Y1JVHd8rOgKLFlWiKHk9mhX5LCXAC7KInDYYMY63tSNgb0N2f3bwkvHVa5H
iWaUWN9no9aXj/wfEtC3Vc5DB9XeKGLEuSXSDSeN6n01A/po58f4LcXKM5uTBBD7
sMe162KhWpjhiKvd6pKMHjSpXbKuxXpTxtI+G2s0pmy9+Zl8zitul3Pd8WM8Nrl+
Ywn3FSS1f0+hYpaX570NYas945DXNZpEqwTEj4MO7yuBdUp2wSqKX09LvwmE2oDE
KyPClK3OoJLoFqCRHr/lUvExCAMSS29cdybkV6h4nhXoi85gvia2TWKyJ/8LnbxY
h7B2SCsex0pzD0tK/kpcRdRWhXCPyf8+Xmip6IYUWVbUg1u2eTyyGOelcN5UrDDv
xBHcH6grNwvZcQEPSsr39g==
`protect END_PROTECTED
