`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EEJOef9LazeUstlC8nHpFKp3Qc8jr97H+26kfnTtq7jtIkOGvgkzHBQwiWhpE4Jo
jmB0PVKtfxQEfW/3dQVPDI7c2PyD1epphaVNWR/P8sbUPonSrUXFgNBsr8tEg7Qi
kWw+wWI+vMlEs6oB+HygdVIhRqH2qfxKaZdFN690CINM+2vsUemcK05/4Hvb20ko
ytAJSwjsDHyQE1CqEj6kbOzMNT85tf7dau8ze+RkgxJz5pu8hONxoH36LKzkPyRb
mNrvthSOQe4XJxwN6yXTIXLU+4EBK2Rj6ozP2s8+33gd0O6TB5koqAEHE+tfMA0O
lDxN2KIWDAiGTLknGW4ug5ykqWjKgg7LmzSJn4ShM6jVlLFvK6O5JGiNLetNa9YY
AwWVyHg5Bpl8ZM9l+DYj8tzgHCz3Y98H6yv4ntbvrhL2I6xTg1wjZvu2YDCwLxvN
LYNxTciQ9Fsgk4NqH9ULGfBRD0aqZPRb0OEpHv+HTalRBRb677CZpjc9blnT+zay
BrpGKzRTZVqKmF4SSr9qlFTISzZ3H83z1YrIgf+OG3Kzq4s0DJpGo4/2IgYEP9FZ
GqNLfni42+DJ7XUpA5cF9yPDNtRPT4eKp4VR4Q3EUF28GbUFypXr6AA/E8rLW0sU
COFKO+6UUfKsGUNCYAdLcfjsbka2K/+zah2f308QmZuwkEiXbxpGYw9+Gpc8CSj5
Epg7AQOE0dQiba/+5CA92SAVO4kv/4A21ktmTyM5kHm72SLKzUWifwx91QJgApDG
nwNCu1ofTNQ7QDe5QFGRPFlfBJwvap5fZpN+ixrRe42uq68VNf6rU2kVUb/uNF1B
sbgY9tz+2sll+B2I22AxPX36kPouE95rUxDuhPVbi90UmAk7Zrw+YVPx/8nxgKz6
+Cr76DB7/ncSwtyCl0lBOugXY+it+sbx0yjcp1V07jkxvmVQFh2+k96y7pti8uQT
QMw8tCbJhmqi6gmeD0lxsbdC/Gn3jMyzOJlZun375aKACgl52ytEtQBGongUcNSG
O/WK52ovLVevH+YLcXbYKO4LIIWEV4dnVSBPs+dvF8gdrmLcyouEjecSPmwLvwOb
LCXNfzsJQx+WzJu8v39ZlR3ulb6JFOti9+xzXLTNOGPpatwGjOT688G3ZNPMV8c9
UA73U9iWMzM0XS+m6RVO6+0axwRMSaf4/56UyCAeohDWGKUyrTFTuuU6DtPks7Wh
55QY2BfGhZ5O1Qwi2GzbMV4GYYsThHL6D04mdu+Pn7kMdalV5Bz1wDC8kTj/wLLs
v8npKo6GCs0cJ698Xlb/0Sun4IElGJnCyXDjO8k6fXs0vROrCI4/m/pqJHEJK8lc
Wk+BsR4cssIxkfOQm7iZzEtT47vDpBrFnuWW5sLyKnZW1mMZtNxSi8CCKsUDFT7r
6PsR1Hlj4L1uWtYvJ8CvbmaiUODogI8vAH58rZznB9b+y2atuFOFtPIfsjyvW358
PTIpZ/oMbKMsd80L5mMtYDGdrk/PscdZdRhZsY0kRY/ufMcoKLlWYZwT3KX9Ti4g
RpHj0YFkQ358gXDJCVureoYlnjMXMDleibQ+JHOuGYEA5TuH9uXz53iMW4SmqmMB
IBERRk1Ci31B23qTFMCY8TskIZ4ObJ9iKdr+X1J0pxqwbtvww+Ws9PdCOiLfCDKi
uraCWW85PmGVWeKXg9oedA==
`protect END_PROTECTED
