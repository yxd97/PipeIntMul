`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2RCYmjyT2o1KGVV2W3enS7coJmWb++6rHKdRxDQDzhAd/gTKtvrv6gB0zbh3aZ3i
gQVGcdga5Yw20AGdB09jB4o9BW8tXDbkcg07V191A1mVLUCQGg7MZwyQ78rBXoa7
abDiz8fhn79zevkq9/AKCjcTDFkhCQoS5QN+0rX9UC2b1s6ZYUfmQe22dv/xyedP
bnv71Ef6+8ZVpNVKbn5CaKiKoVOzrVNLV+mi8wl8XlogIRdAIggYn/bkM61jj7LL
dI4JZrtkDSHzWG3ZRmsqVmF/ke9SIc/BMOj74vsSpKRWWO48aRWOC/OYKevIRXcm
Fj2O1QQfSMOi0KVHqLUELjjKh+rxBNTVW6AGao03UXZh3yFv3qQJPbeKEWUfJB8x
oJyZZ1GDoEIqlZ8fZruJf7nIZXak+2Ep2JdWMTkGVBq7haPylxYlefZxSK7iSEUv
/nmewCtaofX2k952ZZYsXsj1VHQTM7c4lzYAKe/bh0SAE7MqFKpOAN+aUI9r/qEo
`protect END_PROTECTED
