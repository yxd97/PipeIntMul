`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3DLDvqiwgsaC0PHb1bzLZjwvBCeSv0Ht4XjE9R7rYFx9FhMATzVmwFkx/zOliCWc
AqI73mL+s921UJBYImABDRGoW7Cq/pc7kwoBog53W42AN0WeOmJX6fJIqmcq+m+0
Wku8IQOjH3fKRtNHvpUXpmoOHQvrMZGXuUcWfxeOoPA4jqBdYrngr/kJqrVV3WWo
WJa+BXZgxHLtxIPwaQecrEQALPyHaWfKm/nkqIhvPVFO9McxzBhkcjS0f9kinqL9
+3e8pot2x++sA74vRWbwgvsNEED7kU1rIX0tJ9Lax5cHmWthnCaN9b0SKNpx0wDc
6QDQfc6WUsoEhPi5tRh8NkeLGCO5NCPMGpLaXD49oRM4/SDp05FRawJpvvP99/1+
UW4t0Br/qkWmhw4wm3l4BBOMVs1tB9Dbsj+4QlQeGbiO/mNp+NSyR/Z+zgQ5kUu7
5lKeOjWBk0NAyKB+q43ojN79EQ4zpSkdB1qG93Wnhzn+I/kQhFXtYNOSFKcU2M6W
8ESdl2vluYP9L7ZHn3m70ME4Yvu0oOv1FMknRNGdLXS1M9sL1CoGvWDB0BFiX9Sy
DMd12bDXpxRUO5Od1qAfkA==
`protect END_PROTECTED
