`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SHQsutz8nUViodwlPMqVC6cyhsXz1RfTdtj3uYgwmbjcUTsRwe3hXmOdxvxGHQr
v5SylSDzq/j4iPAeaboRbwnzMI5fWtpm9C1423cG/uRkQ3KnnkZl6Mh4N7Fxoqf0
lwXsSL0+Vzku9XPHYVNTYbuADZrAgyCs24h2m6rGXhjtkJz3yZmhHv+UL4Sn3hmB
NUEeuTqa7T+ZMPpRyRwjLsn2YOK9FhoSllgUi9Do8vm9kA27cNIHJrU+E+k38N/1
BtAIpDGQFXM6+iNz1HTLmGJZ89Soe658l2d/sfKOiU3Rl9nkmc6N5wTmnqmyypsp
QtFesMp2GXiAjsS7S0FEpXlqxbqNgTojBzemPNzmXphO3FCmgJaECkw+eBYJdq9a
wIB0rvJPuUOm2NjSIBPHKZqjJrahj6omNCr3ATnQwY9hRciUSkjhYV27TjCVkTzw
u4t2a0FQ0+bTiQX/Rhj8E/Nlkn+eWfj4pr2oaG0XG48duY1NP8lXZYxgza7gicP2
CZxxyD3ZNvyycDRwBr13sHVyqamjvnRZNE26dj303wrrjq2fDQfrr/WytRdwLMlS
wvIBzf7Ry/PbGkOOycK09OdV3NXO1Ipnh6279rmsUxw5WwMCNZhQDAh+7XGnVRhz
eAUEJ/u5T0bDxfSzjJATFm3psrF60HP6rHoqW7X3SG6F26q/kEDuTVAL5sseXrsM
ifLcvt2TQg3C3/yPYMvRvj1RlBsV1El9sdLH3yRkKh2J629DLjN0vMVRzzO1WCmg
D4FuzrxWtxnAyb8gkfFC3g4yK9YKFc968nVelEILkRtasOl52B2ee479HOAzU2jX
phtyQWAMdMFvJKIIfzOD6h2j4gwvL0QgJFUdW/XR8w+bN5H6NjqCFD9pakITqBWY
D2sLU5SPZu9vpGtMxSxgItHkY5edYxU/X+lXOLuHGN/ngwhPctkWTdcSYpuW1y5b
iEhsuZTcb7V/jre9ycnoI+XHhh36fsZVUi0zwMZaPfwgyYgK1VP/G1kXTcM1sxSj
Ndgc1xIiBzega+3MqBsqMgtuxRBh3yc2ZziqY/aQhBVpADmUosiNXA8QDcWMxvvb
sCY3HeRYTr7WrCiULKGJlgHXSVpp4mk3MvwqDc2IRy3ETQ9GZ4NQ07KXD0KinfII
7aVwgLgsHcJf0c5omIF5fXKcOkdHLwYcwiBRXWxDNvuMaYqGLfYnDJW+7axb91Vq
Pg+ZcAtRRCR5f8avlv5m4u2ua1SbQoy/8Rs575fJtF/9tMmNk7LUqZ4MkABJcohs
`protect END_PROTECTED
