`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GWxJtvgSpfziROUWrP0WvJNpvnaiMqx25coB/TxlKZFKAcau2q8OKW6oYDkZM+hG
6UQsrLSRgHQnhLWJIsFGZ6oc9xXY00Go/s3TFXUDt07s9Ghk9sHE3sWUtYOWAH72
0cM+o3Il32G6oqHthSO4iMa862vJw7oVbnPdLyGZGi25aRY6jvyuE1313m8ULDVL
3xAOujk1Pou+GvD4Hhq6zlY1CHPmm4kJHnAyqGs5sJ5Vr5YMx9t6OUWlOdlqFZeF
iVRav+tbMKVUu2gs+9zM1mrDvuerLSq2RGjAJahwaxtI/I1kD1/ltizelodVp+UI
QsWxQx0F4sJAuD0tR1hlkQHByE5Ca+RjkVrR2Y5p5ye/LAhaGjn6Emss5ZfjVyF+
yWNx1pkvtgY734M6CTA1JOtBnBIkw3tdVlUlVAnEe+Du1gLrc4k3ckas03mRBHiF
`protect END_PROTECTED
