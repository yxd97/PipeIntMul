`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/eLdBWfIpiHiUJjkMU0GGYx+Xd6Kz76AsqNeumRCCCF8nVemtuipklC95r6ZSEd
buxjUFzeznxgXszF/Z5S8nDyEdsOuhY0UfYAjGiADa7QsyyJDhT+E+Kb/z1NArF4
MCV9u0ZYqOQx71WYanhpu5AhJr2/EOJcJxOxJfxbUZhWXqEND6XSP2ET1uNUPM5x
Z1X+1p1uaU0t9mjlOLOC6MtSayElZxutyePTIK58Be6ZiswCEmAUSZspArXhAlkj
MH8ydjs2jsCYWAOMi5l7h3SqU/h4P57hNwZMSuld7mzZz7xndxzvFA/nqYgpnJm+
njuPG2j03UeUI15gAjrC/sf3Rja+lBYh/o9nnSNp9B3zDQH0en7QMd/Agbiop97j
ROTiDN3i4m0intOik74z5248b7m39iCPomqr1J4Doyb4akPUxvyhsxrv1zP0/OFi
o02jYq11uH/FvIdfP50oO9ggKofzZt037Twtj5Fbl2iF+5GYWorwhsNXYt4v6VOv
m33lfHqDUY6jS3vv5dWUNtfyq/nMzcRHd/uXfVqZtbLXbQ1k3RyBzGhBM8O/hTlE
dNUpS1veKXkb4uXTtsDFqbyF9TMKUKeXIiuF5+DSDc674OIVIWHGnhdKbuHGl5nC
93FROgxRZ6Xbwi8QQ4mIxWKCxvzneyDaEGGuLdD5juFIXrPMOJCEhGaRT3GGxy7n
nrGiCb4H+B8c9mfEFpzmKrIks+nwhNvBXCmvdzaQRcxN5uQ1ZvbJ3FiRb3jDfVM8
YsVAfKRafH1CnmHu8hYWmEtaU1aMAc577tJ154GbbJGisBa068PUFGVJOO0UBQGC
n8HIvVKm8VsEYdCo2OoStQ==
`protect END_PROTECTED
