`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NcX+fezLYKVS1afUvVJWexa++gy3ejAmZ9gAaVFU61ALiXStX21/2TAoOY8gMXd6
mlkMuHIIEFzEaxZLbOoe3i0Hh7I43t/IkW8mE+S5g8Hh2hfG5VP4b5lbubQNBMO3
hR3vsZwcsH5C3Cqm0Gd5Xur6CiIU7tumRItCpP1M9F4eYeZulOmIlUX9KXtz+/BC
Jy5Tssnzo31xo+QW+uGzfJBmpOEp5of00YBmDx2WXDIA6qHE1cgJBEBuJ2TT9BIX
Iy/pkx3Jg5jRZyPLPKtcRkCkYX78SMwKda3wvxamnTgSEgLhj8U5JcuhazyffZol
rIpg0PV86F4QTgqluCeo9Qn+oBsXCjCJauBQmiOQ+H5qUhtCuN6SqTiJADZyD7rW
IsW3DyO4QwYm7mUIp1htP14hrWlXb6GNmZ4YCBgC9hH6RZ80Mhc4KxQ+CWJMnalh
VRp0kWe47iYvJmKXKEDWJBJNn7RvWzP70OHhvANH7nSYeCv4hwFeRS6syWze4FBm
mMtDBbvXLjUTPHWXL14HqvBMI6OsjDreoiG7zHoKwSPGsJan+Q+P2S+8u3Y8k1r1
mzgVt5SGI7nJ2AJQ4GK2ZiKQenW4ySI7GJUQ3vqujBfA/OrkeJz4A8ZL6aeKSKY3
oqtFoBPGoawZATR3JGyyIeg8Eb9puNX5CBqnnSGSLQTl0Q4SMhaIUUFLiAZVzjB8
G40lnV7EYZkuBMLoSxz/5a6BZj6DrP3A6AvA+XGXawB8fWK03nAPs7Fi4A5KC0V8
WjFCGc7gDDoBfeTg6VuE11hCfsy4zpuxpIRxR6UPGZmgLqAIvSu23a9+NF/uT7+J
pNGpEZ49YjOy+5+ZV+vvZ5ZCHdeFKP+HTq6WSxyKu/aINmIfZk6RdMaQiLu03+Na
yWzGrtuVe70+NX8Q33yzPFfaafZbEujvcHgKR+Z0ZUNtyxTom5amgGDdYXP+6uxA
W3oNtK5DCBnCZMQ8gKF6tQHbQ/CO5PaBmYvcAe/HEX1siZHaAdPzPBqOQ+0gu7vA
eSRuFyzLzXFvf9JHnpNWn1UiIePwJFUbjujlKviLyIRcH1l2PurUbKkDYYBfKGKx
qEVLejPnczCnxsozulKtvPH27C5o51hCDK0z+1CTcFO12Z7pAYM7GIttngWRCOV6
KfA7So1ZkxLWarfCcVANjw==
`protect END_PROTECTED
