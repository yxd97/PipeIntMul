`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3JX1TUtKrekN/Z67TG5Z6xoCc9tDcY1cftyA2OhIW4NWoZJmFh7MmY/Zl7qk4Ols
zD+xo3TYtDxhAg43yQsaL4qMWjCQUFJo2LwVP1Yom5JYfpFAI+PRBDzv8hkWiSf3
Q09nLcIFNl48cQn+xgGWmjD4saQDaXIY4DoY5Cay/NWd7ZuexsMSb0oGkRJ3Vu5w
sIp4tvQ6/+dfw9DucGV8ISSZoDasZ6wdhaz82GU9WBS7U33rselI3thiQqIEA/pF
rqJJITWxoBqFwaAuKEHfNU0y+b63fxcWH//yzJV9Y7yP+dlAbPnoQ5z4efb1rIBR
CXAWWlJKbNRe025di7kfAcmgr/0ygSTuWFiRnBs5gSFBl6cY5AeTiFC3JhC1ysU4
0YrO+8kqqI/rcrjeQC1kLur6otEdFhxDZK6Do3ji38W6NEPylmHlmoMxU1HW//7/
zxJqSaVZIh1JhLqLhdFN+zAlv0wewE70Vq002uWGfV+Rq42BFLH74UjzqnTG9hmA
cZ5FQeGcY8yhs1A38EXuiwvtplfa1/HOf9SpZYKir9/FgjNY3/RQRi7baMaFqlqO
RXNff5us5NorVftEtU3FaPMdmweaNy8SzyAz6Y3AJgRwqi7ebeYSSTi+04qFCij4
zCHH5PoYtSIYkyPuZMBRXU2RvBoPuWXxxNT3jDkNeZI5BPkmFs1ehD47tYfXOAuf
TRPQ3nFE6j5hkPmWkARIGAZnmro4z/MW1YOTdJJsO5RNR/gQrDs8q0n0e3tBrvvG
pkaCXy6zuqQeIeW7JvPfCLu0NFQZevya2AC+EibMldG8rqijSj7/QD7RRWLqaBnf
`protect END_PROTECTED
