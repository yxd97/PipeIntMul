`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dL0gRCKyg6gDDEfO+vqywh7n8iG2hw9gdZ1a8SucUVFNpzk/5FlN4Oz7UL0oSLME
tLzJEXIB6wUntOSu4GL3irZK585dVc5wzX4JLfjsQFEr+4bz5scwVb4XvebzzN53
Vp9rWtXYSKkKwJp9uPrmK743zoOFdJ+5hbgyhqR/w3PO0wHn/uMcUk3iYn+8t/mq
AaNsX8IhxBGmWXjj1Va9Z6WC9e/cdNe2u+TUXu2NFEczaMHVifi949sDY7aB36kV
nabHHZbNVWBFhELMOsbdR5qgQ92HVF2hUFDYxiY9/30zPKVPHRF7nKJ/GmyYmSK/
vzs3Vt1RXs1Bh9dap0tDvhgUjZl/HnA8DyzA5cxPba/4JZ5WwkKrg6oFdKr83Vkv
f5rZYeQqNi3+c9b34Kssu8zz21tb783jmQHn3QiU1tU=
`protect END_PROTECTED
