`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03xDIPM6mHkgUcC+JqIMnthoyLCXhoCMKasA9Pfp0b4PcPmMIyb6cC8ZXDLqT/jj
pMLLQFVsP/E5m9B2RQpC+9oNPF2Hx5YC3xAmhR0IRe6b7CwnlmOnKYro/zi5WDBC
34Ud39+UDWujGk3sFZRq+EASN5MIRwnLW2VOKeGxWE/lVTkSthZI7RflkgmqCuAN
inln3tO9sh2fX6wdy4x5wrNof9h7maRY1Xb22x4zFikGzS0LiF2ze6GUeULgEMKU
812KHdRRScGrLnu4Odo+EsZHJ6RxkWOGYAVo2qx1gpIooBQ7trpn79E9OF2p7OuY
spke4/hAwQbHYwnPQQwBnM4CkR65T6C4Xl7VHWTiOMPre8gf37SovHDNYr9yhtP1
nFRe1Gys596AiVSOPv8QZw==
`protect END_PROTECTED
