`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hk5qf8qzpMWeQzapU1UFh8pgoaPwRiJkmm8ohuZGiS9P6wrUJwDxgDCGSDNauyj6
EGWvto3mIKnkgkaFywLV6wlcbuUA1JBBxeBYQJUG8DgDh20iUNOzY9U545s5kNWe
Kan5egTxNS5KcxernHo/1yqPNyimthczjhin34okI4mV93mDPdD51UHqsW8i7773
c5+1K2sw7HGXQOT1qvhg17/8H98gcbdt3g/u1G8/vBgjurIx2HezE5empeH3Ckyn
0GUCDtRk6StmKK0GUydtWHSItltnbbiPEJwUjcu8X70RggtlYXwxdxz0nyBa0+uS
zS/NpbzJTKnGNWJOhcLOvDFHTv19Ds5r5uplz5SiITFfXM1CddqxqPs7eQTeuUWt
WOVXx+LTnvhBtODWW/LOqILW6l7Lr2KsqbdcBXlloE78wOtbEipbaUkXXH4TC4Yo
zPaGmQc9J3bl621v/dk545zTnKrEYpbygAcW823SwU8=
`protect END_PROTECTED
