`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wME6fs3TEvGGck5VYfGjBYtjQvFHmDgvNtNUUjZsEHa36wcdH+gKEBcDIqryoyw4
wv3Cxvh9H2+3lIzBgApZZl1XwbXZfLW+3mJwJJ02Gh3nanIbxLd3tfMjqRoVmO4D
/EpiFnEp0AXRRvE/oUlh0JkLGhOD8lweQuwxm+XJ9HdggRUYUoxbdu5bDjPRs/HY
3Aey/K0mhJlfecunZaisSh1TSrA9fPn3BEfqxLa0L3KZ28NYk274SErZ3Onwn8UI
nleVzZrof3sg4O4kE9/yMQi4DqcnwjHoMT2IEMY0lav1qXPek3f7dVA6wG4Cat1T
n5BUrvEzFV9fWejQHMFuGk4jR1g25IdyNZw9u/0+4tJUsZ67Ad5qOkDvd52nkxjj
588vAKHrpj/FcKc2j/ik5wW10lOFgE18pI6Ws1BEdIh5lLOLFEp4BggUOXUoRSgC
Prf6xLWq5w8nIctx4dSJFw==
`protect END_PROTECTED
