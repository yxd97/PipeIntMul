`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BnGtj7PRfWSei9+6XXr2lxAi5HwYqixqODOho8v9ZOLfEyEPvAqp8F/kY4OYbqe2
CfUzlhsHGZ7iEMu7K/vLc7mA7pbqcXIIP8dF7tf5Z0VyDfuzbOfzy7zokRmiW3Db
Z3htMlc7lpwr4F6i5rtfRN9fmOakkTzV1eGMQ/HYW7KUdCU1J9/rfXIl7droPqtj
gTbewoAuhiNnZrd1FxK1Ou1HnpSOfMmBrNMTFvNNarKFbXhRi66KWHjBA6+iSeos
XWtO2M0gnmY7QqDcdC1NG2MoXCkrr5E6KIrQ3f+16Cq6dYBOtKhYjcfeaHoexhh4
Z5Nv7srAAErMiQzb9aTN6tRI/Bdl4kBJQIeEhyCn7pmtfpCqgbGsWHJRI9orilq2
UetD+NP+l6rJ+iKds5m4eAB2IJTmdhUv+j94wCua0Jw76LZkq7dIKHZtC7vS2TBb
hvJMLn3mW5Rixr2qmq/4+/4Cemhm9PvSthlCXRSE2S/GuPYaUj+e67RG8ivIqHHA
gxeBEu80hkisS9k7ufK8r8LfuUgyr1PKEawssfyuIJ6/3OGMufAqGR77lw6obJlL
M2ZE8y2Hd+ICu4j2jvQCtJ07/8Upv8SIajUm7jiqYoql7PWWPqAOsl/16Y0OAXnW
j/ayFU4yMbWGwxyN0MBCzLSzfoEQR3CXvBuWHoIbdEKYDgGbxajV3BWyIFDA8dT0
SujTy8NRcxV/3R2BRTOSpIqSbH07MQ3ereT8Ec0Nyn4=
`protect END_PROTECTED
