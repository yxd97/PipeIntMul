`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOFn+DybewV01YAjHAIQ5jxv0XpoLzrkaJyxSNqhe4yWFUi8fpnGkHZwVOSRPHTz
Xy4in/QmIJRQEWRRLyjm0IWI4T5JVwd87Pm1OhyHcL9OdRdtkiKqGJKbwQzN4xgj
7wndAoZSfhWCkjYNq+qepatjk5tNz42WsiAdH1pMywADU5DmNGHocgYBndrItyd9
85XgFX1W4uvdNaGOr8548VWcaI/8DjdceF9hQ+cA55VeB3ePB/63xXQ12qjkM4RN
t7btei2qO9nzuWq1Q+jsviBC3X1okY0DB2Ysl0u5uy58BznudltnzN/NApok3NiD
eMJxh3fkgeMxbQ+yGWW0qMv5EsrggAJ3FgmM82xg3DKZJoBcZmUJQELWArUN5Rp+
+q3ASJkPBrVmyyOAFiCALFJBmgPqrcyde0fZenHbkPw4e3B7Oo2xvIrPulej1I62
`protect END_PROTECTED
