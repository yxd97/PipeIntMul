`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/yGoQBQPvaCcQfLp2NACoJLl1LqitMQYLpXR18B7l/y178bFVDukMEjB33j0G94
+LogK+KOMKedogD7wbBURIZGtwJONluRqLRCnWvRxyvBT3/QnvNDf2Truv6sWJhM
6j953c0llGBkw74oX3OX1zAwdH7eIkN+YSsmV8GN9uctZuGjA8TVH2BQKRpbYyXi
bGK6RQZwLOfy6jKZhGul2Vc6CJxw7pULeLWwzSxWrBfl3Mx+9hqsBS66gcAgqfAs
ilABpheua1h3tAnnyVDzHg==
`protect END_PROTECTED
