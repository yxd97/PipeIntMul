`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W/Vo3KeiUjPE8o/doLDXHf2yNooq4Mp4e9EMWNuscSuw3+tVfHhhIxAvPxoGHrXA
PcPNeWwecharcwpOqwKCsMuX64DWhnE5El/lTQO0+roN86vUs9HoFfiZ6Zmi2eRz
Q/Ediva7h5znJfF+p8tJKjtBLJXM3yzzwJ0kGcakKZIA3ergt0Mr2kwM19tEvuRQ
wk1L2xGS/ZCne1Xnv+9cRco0FfLv3fOQ9B0K3jErySO3b/7daW3dw225RjGGzFdM
JQRnHEJNL7NOR5NWO4uTcOihJcosAvG5awgiCHjq7GG8Ihdb9blSMGjTaL+iIcYQ
/W+01ADhwSi1OoQQGHC047cfidvTqQX8FtpIypoKqJiM/blm4PZB1citivGn4xi+
v/awV0vCi38kABR3cWRmrbSlfmDnESA2kHigPdQ+syXJWlBGdRYavz1UT+4iZTj6
guLOQ419gkMtysXY7QQJReSkTENtYe64LI5Ei3PjZxJX8vRrXRx2/lFAZIRNGIvS
G5IbvhDLBqYW2Uh1H9GXF7L2XZG/L4AfxDxiktF+lZTRYRvPmSAmxTnBZwtTCDmi
q7tkfthjkhRgMenZRWPouoRp0hZRAb3foqk6dB8ZcquLbvfAEWpv4/KhgCwP0USz
Eogz/gUIyBX8iynRxvkNkg==
`protect END_PROTECTED
