`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryKqCyOq6p/3AuJcveibEjkxEp65IBpSF/W9F58+M0/OGTO4O/baPxoJYJ1g2IX2
dsVgIWByP004kwq5hZRWf7Fcu+gYMMJ4VXbAzUXg/MnGlFpAL7vjUW8gIBvOU3+Z
s2QxX/GQ1GJ+Qj+alXGvt/yoeY4E/vMIAjujk77mzz8OjGJ271wOCS3czo7sZW82
bwzGwfoL0XzBWFgC4XtB5iXbYgn3ERSongQd2ELR0ei5hjHCOk2AS2NdCiHYtb2f
tRqdTpelfUrJ4zjorLsMFRn8kc4jpt09nb8VuLbNUtNXIdsFjAmD5eXZWguJbrOS
Yn5/XcvNdZVxXcLMGlD+Jg==
`protect END_PROTECTED
