`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejVCbCRzKn8/Zi1MsUn5IzY7UFHGUeWyI6XVPm+gWVxDRcs3zNEnSbauy3c7dnoz
abX91kj+f1MtCC2CW7lqfnLfSOgOb3dp6buNslnYCrd/bFO56qwdL4UpbRE5mOY9
g2Mavnpkrdk+1rLX0u+dNRJURTxmGuWmEl9C9754eiPMinygKh4WHR8FNoqxqo2Q
90E2FnxneJdc8RokIRy/6i63eq7B+TeBtA+bP/oj5BqeULaZTwneZc6dCQm6L+2G
gyMctLLgIgh/QlcGk25lo9s/5alG5WhkEY1rrvEFsyNshh1upKrxyI2ymW3kYvvC
ZWbtELvuS6LrQAwvuOkUN1H/0+EGtup7UvfoY0FPsckxixR7wV8SpHf9fF1a4lyq
dCyOwvCRAnBiMNYgcrzDaikdnauKGxwrz5KMxkvvziLC1iBiClOfpl+hJrQ9rjPh
2DrWqP2LjZhFauxdx7g/3lPqLzpTvC5gFnO9WAH2eaSs13rA0alP2g8sFMso53Zv
JSCc0cYIvRs/1U9mUplVWOhXYkW/txBK/8Wq4N59r/A8rDflg4O2mz/wmnBu8WIO
vb0UosMhphn9SNo3W0oG7QFic04pgK+hkBjjO9o34/RV264bAupOIofZSCvVIEBo
4rQgl5ZuYPzD47POfpn+GM8yLZGXNbb1VMxCafUj1GOcYQmYPQwDTE+UyWNIY7ld
tu6LCfz2cdoz9E92CxYwVQMDwNtPCuWiiHCdM1ZGpE+WqQZsRhLOdjCzMcRW2her
X1FPKTKkaBcOmImcc0GxrsvGggN2bhdYcjcFTZ+OfaYG8DD1bPkVd41BjDwybMwZ
/GHc6lqBVSeNubrlZEpSq8Ihd8+o77u3wu5w0BaSPo3DCiJMcbAaQGE9JdTy2XdD
9d3rQgH7uj64xQ6SpV9q4mo4vE0EAmht8PYdWIVJCBbsuaIjVovkfQTM9opP3iEr
9dIvHfEFGA/rKcZ2oTRPYXqTvtcFKXBYhpqzs0FWACUS0rU/JNqMoy/j9DB5EFqR
HTtARb/grWJRq0iOEP6RE6VXINZNw4bDmctMvMSw2Xwuumj/zpO5f0jwbHXRebje
IuLNo+TKGJGiqztgrJ8cpdLKOdde/guNly4FQtHYnSVM7lIK+iKDP07yTckbKp2x
FXFgrmGyXYjpjVzr/LPBLUyBKwtA5/3FzpVH5QEWZG3hamOaTsXCdSSt6l9bGLjx
xV9ASSrqcoHN14fvLfduqDWqSMgwwE6jyAOu3RakO375VxFbzDGhD4+wKj0Pobj/
h9nGUEueHwM3NX+msXInNncUldFMbGdXkCpGmYUsclXd4DBv2tvkm1HgiCXHADS3
DL3Q4blwHdx94EUNEIG0hi3X4o74IDHWfDtE0t1Pwmqf1symIhWMrOD7fOmVXT6o
koBhaaIvrwPzRpncVGnybN4Q9ydY5P0uSHT2dYIOabMcP5DgUhT9RmWmG42TO06K
0NhJSlWop6KSeHefuVsoCkdLJI0rEWeRCVSFMPhOQLwMbk66IBAWAuTrVDeobp/e
yWARkt7JLWcSRdWa6iyf1A7WowuHGoPrNUsgM9Vp1lqzbem4awBmj3eEmcIwzO9p
BzQPUla1sud/wqfjQTvGkPihTPyiVKrC9Q2boyYEaHW0zXYwU3dTCA0gOkAlHtTw
60dfaLDFrQRiCZPsKTTuxUDTRg6WswRdppqnAy+XRi7U5g5fUeNK2EltD9Xb12dI
f0SHVwODf53yfD2lRx2xhrxptzkvQd669tAlIqj30Iwe8ut8AMH1xPtp7Cq7nNp4
7y7Mg0CuO7Tf4tr68osddprnQEcVL5KEz7maamy/fFz3aODRW8v7ZHX0lfWI6CP4
5Qrz6SJtgdFL7PeUSCeKNlwyHa7T+f4lTRA9uFwqFz0xCphWB7JyysSNVk6eKhdQ
nENiOZ8PASEeClW6nox3phxIBVZyi5ZHIoTmt2BE3AEi7ircLVJYBBuJufD04gBY
2cNMics4kJ396ZUH0qZEs1lwl+/zFvGytZYTm/ieWgIYUpSL7DhL+EPhIKM45iB8
v+wbKKOFIq+nN+luQwg7jdfFxbfO4YChyMwd4GrHZkCSCw6IYVN7/aGHHOm+yQ/9
7VmR5N1F2BZgnM5xhm82qagzhQ8uTIQuXzzzIlYnRM2jVrfBMh2PhULtE7ucec0J
MfQzSOgYErhOVtyzi/qTg58JoWGGYM16Fg5bjDVC04TT3H/nyuMRCP8meCAyPTMd
Ecp532tX3zqmzvuieFUiSSDfLhYFuNG++yXGQNyWhjaB2qvkyaTCuoZb58EjkbnS
IUi+7jZ9zJfJZqxvvNhsGaZRx7OR7ceVDRQjZyyZN/5qllGh1rv6Vpx3xH1bl9CD
R5KBglBo+8NBXDWQxi+NDqHLsyI7mR3iSTaYbDaClp9ZDbRJtwPWhheBRYtIePLn
IUlQdV2uGTBRtP6tmSEe6r0JsE739WfhIsZ1CDhW+FK5J+CLwumFZekgJJhWiiYV
XMMM4XaWQ2MdJmp3jIm0x6WCmqflm6kBwq+RNKBXrxAkSQQ9k8Ugu/qxVno34p7a
XfcIjQB2DsS2IznIFFGfSjtduqJb/ptwmWNDSqcdeLsvf+Th1ubz0VoOMeZ9ykcZ
Z6bW9LX4GPE5M87AKo/rbKQ5Ht1GbSPF0/vtoFR/7CBoG5+YZODDppHyB3aaZKMJ
QNdW6SkRXUzxWuBF0/p59Un46j2NbVCLl8QqKouUBfaRwJfMqa+uhMmBtrPc+R+9
ZOef2r4U2hkQexJ3jseH4eUmLFAwGz7b5K9VxqiAXAxqOdkt2bItYM/vDOGBUIz4
lgRn9KMsVp4MMK1VxWGQj0N0rLTwCIfX9Ova4404VIy/8JBQ+wC53umMNETmIgYn
XsZn5vePTPom70RgeLrMlfRDM9hV2cys9a5omwjrLZKEKreBhwVTvCEhANAP8QJk
781K6C2QMD3eU31kxbVrEy+YgZhYbG6YR9GlnSmMBYV4zpdtkWfW8C6kJfd0vZYw
wE/j+XNscd/4PHUgH1LeHZpduCipztcbR45FPwX3zXoVAvPnV2tisyP2V6YAKQYw
HCzj7sD1OgnrgVNCqacvb2Vm2qF8w161nk2KsE0Z1VmJqxmqz5sMtLIBxDILk2mx
a/iKNzkAgAYGN3EKy/WknLlivXuOWHVOWPQCZ15N/k1ieuLRRXcsCMSInS5wNKo3
dKjsCao4d5N+/uqWPLb2BcrMAvGfvMvYs+TpGyFXzxalP3XTJ32h1X9JSJXbe6Nt
XvnbXf6fwV+JUrZtBdizGtV1RNyz3xknvUjgFOkMZ4sWm6zVgR1swI1VPZs5iEuD
dHzs430eDZ2JQp2XRgNcXEGArMk+wBrlum3s6lVZ4W3324md4U/Wwg4XCe19yHCc
26xd4YGy3MvYuunZ8TMyok2E8IAIf1czHOoBDqh6U5WGHQxas11o7Nno5Civ+zDp
noEzcb/zQF4JsTnuEaIpVFzzWNnJsBShK9cZJHfVcpHrF/dL6xPCHVO/1HRwSERd
K2Ewtq8JR8OC7HWi6rYktExb/NqGHEH8QZGwuizvGR5HPUMSJIkBKixmfdEChJzT
aVW23JPwKdxZT2XBNAjCcEErj6EN1eKCVFVU31eYbKB8HXllMVDgYqsDIy+HY1xc
7Uuk61DYouxd3bVIgYv7YcL9SGTMJstdkObEdyUdklc8yd2MZekS/aCpJtNDpzTw
rZ5GcfLnQv20jLd/TVRRvfKeIctDFAqUWpUkdkZ9BX4iBfc4xuhkiFSKEbrLTVwQ
rN734YzjP+u7tCt1UQZe1jJTFRlVtB2fujVHTnoR376qSDeTEAu78KB+F36CubPo
ZeGWTTNu4Nc2IHgRJgm+/EuGLcrl44x18W2gdz11jX2rRBvL4OtUnTNUGsHTI2a0
mgStmY0Wj2sylH6U7owC317WkocoZGBLzpuT3e2WK66/u7pKYQbhBUfH5zo2K781
5dv8VN4WuNnzBwBdkARrzgO+tHhE/j7VVlOYJjqL6ZZtg42o89vm91vNddy0CKml
OKT7aX1wjIKaNH/WPh6jgDIuzweR1BuDiro0mVHU1t5z1gRzb4Qyl7gWZ+jGRJQU
NwbVt05n8BTH6MQSl3WFg1ol7tRQdn3PcjfaZSBjP0XbRPsXJkbqXW8fwbt45eUS
67n/VUoqid+Rq+lp5SvCIAsx2xL1O8x6mDSmbgNrbaIjsPUaZw/0d+b8FLi9PV5E
DkWQjUP50h0hNOeUJJWrfjdhQRXWeI7UftrrGTehWlrnvDtJQYemVnAaQPe/sqh5
XpTMnJDkKZtwuuVkY9WmFt3J/ct/9TiO1HlFIDmoc2IPt7POWxSihr2VOh57F/I3
6Vcq8QiQVy8eAchtZuCTlEpwcuNQfe5Ao/EHDCODhI35lpCF+fBpO79RhO00uwcE
ITc7JzhKUzLcZa93yCsdW6LP6S6iqE5xdGya/f/EIX0FMIKEltJ2n6UpXbP8GpXK
yFKegCAph14g/yCo+zj3oSRN1IM8+EVf5LH2NP3w8WhXEbY3n9pMhDgKnkLUm0+K
xHz6t0ASjsMx8BM1u9L+XIbzQDgKBjGBUw5QELM+1nU+d0l3s6QNzjtwHXU+f8nU
nTY34T16S/r0T57tn4ubG5uYCPQLXMajA46NV1PxK5vgFtAm3cczzx4nEQShZm2L
c/AazweGw7zFOablNTLVR+bxQ0NYIYU+jGf/fiXqSUgOSo4hc+tmUcT17xpGu4Vl
ylc5PuOWrW2BahbDsmyII7599ICg3/f7U/mx1/h8cJT9a2owzcnKZl4jGxu5MALP
zpnmFD/Bs/JOHn4YLMgORqSC6LptKb+V55EwOkEi+Blk9+ECtaG1ornJ2QVxEHxW
MYyUP8SLNO6LkwSaXwKcaI60iRH7aw+N7JwJhNGqv2ZtQEsgaZgjL7EnaVocl/4d
k2LwttSxIpbRmd0TRdhW76YZYiHI3yBbdm7D8Bp2bc7KZRyaNGyCs9GhON6aXOya
0xtxLM7pQo5UnJGRJGxPS+zDJij0Vr0rSJ4wNkfmqx1sHZnkOLysy+tmLKhFrnhY
3ImELlUJ0gOxrupIIE9ShO/VnGkgBUseRRQTPo3G+tgfNpXlWV6HRCwuEHFhYait
jXPT8e3nUW+VXdnhonHJ5awv1ror40IrgI8lfJho1olJbfYEqrR+jKbYsAB/PM7M
FD/PKdJXaRcUF1vqtEw80xTv2Ygc4QAOXloSOVvWmp/C0rlHefgIZwJ+IJR0jAee
lsTYZs+FRFKdcEZEffXLaq5lxQFryj58gdXEIg6e3MabBtC++J4fiNHSQI+hOl5j
`protect END_PROTECTED
