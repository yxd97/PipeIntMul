`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ew1dPyxbD4vKtgz4/+Nz1muGP48vIX5WLZmibFEJbzForVZ8oROMd6rU6qL3Mm+U
bmSVrhidcYef9GxygREv6/AjBo1j05eUIY7uwhXX6JSlXgpKeJSrMe0B1YAG5YI5
vItXsLmARI4rnQgR89mYFX5nw7LnWn+I1KonahYTIMrwujSVmr1OQzfvkDAfLv/R
WxPFJZlBJIY4ZBrc4fx5Yb0VrJWz4Ts+BnREyv7I5KDigI5CFnMZPoCIKP6G4jaY
k2YRC2+GsQoBOEA0gI+1/2WMLDuZiVSSgQsrSYHz6JowXCKGVMddenLmCsCe3g2K
Wz0SqvNw9LBQrmGKtu/f392sj3r8ScTUv7gS7oUfgtgt9DLDJ4GI5ibzNK+bREX6
kEhyfE1kus1SMD3UQDxAGJj3KLejzWeAYBnG356GB3JDXLLWAOmfYz9z0eQhJxPG
k0rD2XrbiRKWoNiQDoA3Jxz/pQmiCaOum00gVT3bouUGo/KyopiRsgzpxq7mepQ3
`protect END_PROTECTED
