`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fnia6rwn0HYO6uuoEdiWqdpckm+4stUAleyptSlEibvXrpSkk42pfmteeGpo+2qb
NCtQCVXQ3BLKkSbvlWXHbmBg4GvpFN9vn2l2kVkjOF9YYngtRuLdBKIfuS31YyY0
GEfJ8jXzvSTeNzSUn6zvnAkgLPOH8ugOMje1Kcu7PbBf3cn9FhSi7MeCI61D5vhj
GWIcU1LAZDgyvTYJgYMDmG+oK+htepjRL4f6KdE7HyFDkiRZyTJIRi1ITC80rdUy
DtAdYDaB/TJIJLwSB+qfREXF3U8P5NCFmfrhaCvOb6BoLbf1PAeqrdxR4KxNRgbE
46v2z9XSdlYQ04M75HOzYVaBFVhvI1iOcfZmsqrVlA1s/vfq7d2JOM/RtTugX1za
0bgnn+w3Xz0DEzFUlTUZWcPPPstkZGE/CTvGz+xAJ9RGKwH8M4BJY7VE0yoCR4SB
`protect END_PROTECTED
