`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
14XF3JAkzsX4xiVabYrkDv5xD+vi50IdvQ8fP02WvCgTH2moJkBbtXAXzSGjzMgo
VjlNJ3+QtW+HxZNgEQrjVcvAGRchktjSjzKsUVBgGMFXoJke/J2pd/zydZGoVDwq
VIMPU4NeCITdIz7TSIpypG0JKkhl0GHSmJpQ/sN//UwwFZBXcGM7FULzd29VUYJ7
pqDio7lqnTQMNpnYCS2KWqGMx8Rt6UnbKkCJSdvYAwcNUJN4Ff9SfD6cJKCE56bA
ylFOTqFl9x6SCA/J1m4xYkV/sdWVFRjBLUNDiFRjgaIHFKUXFBrktcbWaXI/v88w
+ZW2Ymp9ReaKw6CkZeZN+1hrGWlEBJQzgj8hkXRTqtN4Z5fJZoljDydCg992qlwF
3iLB0OeOF2+r4F7uvWDfs+AwioFEgi01OhawsgxA+kMcpjK3h+a9HmHKKQLocBRJ
VCo00wyGyrix+Qx07bQWYbwRskgI+08dXRXm7m6io3WiXR4jvolR4KyM/NLckhLV
`protect END_PROTECTED
