`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5ZTUE2RkWuVROg6JAohw7F3uWOkazdfel1K1qVHuytPumv9eHXgUT4vbENNEm5G
oB6rIFjjm0Z9y2gYDl2KkYgxdBNr7Zq6hSNIOOf23HPtWIU7w6+c4KNCWt4eu9hm
39FFiDVmyMVhouQKrd2kkxI/Pc57jXqN8/zpSPmWu+du7G+JM+vkEkYmAFr7LlLJ
/yF3hpM12jP3lcQ9vkAkyigBdOxK7U3NgsdM7CxKxqSNuxL3DCfYFG34K3gvd3pm
CvJFg8VIOI53KQoCRKAszTZZVpUzaL0dtE5JZbIDfqTaFv9mj19ETZyRv0PlMrm5
6+aEsmw3g4jaIgyPNy09MEY9yw4pC16zzgt5wgGZlBEjTECpI50/Cp97mFA+OhBb
mFYzEIuCpVzRZjhEyjsQLkLeEusWp7BrrKcJVnob5PR9G8CrcYURIvzoMzv588uV
zS4JKBmpiR+YaECZil188pPkZ4Y9r8nsnelF1T+PP6sgw9Zmglpm9/cELCnD5gIx
ca0U1IFqSBBtSawNgJ+wC75Zq6xR+BwvvG/OSyG/qBa65g6zqkfEmhmzQWda2URH
YFfId9z8gOCBMd1NwtobLruw3Cjv3iYLXG1ab2Mu8efBh4x2MwseMeYVAZWqDECD
C47c1ZdkU0zkCG3aRmZS+DXzCFTF855h5aYZJ/uriil1rB7X8HEryEZijoLiNLw4
ShBiiqOZ3f3JqspJGsmW5gjgicrDbiovDnzEB1WM9POVUd3Iol4xWImxxvRcD24G
bAIVXHqoqaSX/AFTErdWJw==
`protect END_PROTECTED
