`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
grAsqkvPS2VmEiuvjDwqMO5++u7/bMiJBGoQSw62Yg4Y+tu68uf3GQmHyrwzvrIU
aVdovZCTL6wFdm3tyuTBi5NQDF1TpBoCzQ01q+Yywzu/PL94cox47hjbqoNCmEPw
k7y6/Pz2q0WeLXN/6PtrlkeqYjR8PEr7UcQHb2OpM8a74R2UD9BXOq2ZDo79C5+j
djYyP+1gV0vLHb7h56tVUNoaWTw3D/xlYYmzln5f+FqaillNKXBHT8Fp0MyhesXk
EpFxqPbJYC3qdf+vilHlmfjDZdjYEXHphymCSh7JZNSu1t/XxZcJaGPa5gtQ+bx+
PeEk1HoQ8tTrWUjBSbmL+iyNFnwnBw/rKk7jg3bgz/U9bt1bViY3u7FFfJQdLkFv
XbVG6leeAX4K8aqOweBmQnSCCaymeKFueS42zkT5ZvEL6AunYtVBEscR0EDbS/ML
+H6UK8m6nOa8zDfNQavX61aDeZl9b2g4+7bsX8RmhaQjWZecT5ejvfX1syv+0mBa
8ToXKEMp8SBK2Wzj+CWcfxpldesJ+tb9/mBIGZDT7j27Nw78oeq3ek5co82Zet2N
2YSBcORIE47O6b/1Ebiiisb+9T9S7DKqAmi/NxmX968v1OdRxdc6RfAqR1nyte+e
nf1QNU3j6bXlgiFOUFjqaw==
`protect END_PROTECTED
