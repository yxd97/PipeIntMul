`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwDaOUwFlgpf8+Lfj/Oyzl6UbX/xqsavS4mqel7ds86dQ+0G6rhTYvrwXAz/4FeI
jNFHXk6xkj6idRXMPVL/STY8JqXzkxPi2UMoyt25MxIxkUgV2LRRJ3P9QQfQMeFx
wVltp/QnbJKCsJlNdtAORiHqQYaNHxR91uoHMprHtHyNymc4EZwTBT3Txk+maAXn
0d/n87zPfP4CQ7CI32RLXI0D1sg3wzKRzIizGhqEe1w8PHSt0cpxZV4titYfvGFi
4tiy+FzClkgazmoCuh6yFZxxi871Kh+aGOUCy7sN38CrrcyATUjupdUCvLjKuVVW
LYFDKSt00ZuTdbljiuqCo+XlHBtKIC5SBZR2GqBipJlpQrj9dT1fHCzuw4Fq7d3t
`protect END_PROTECTED
