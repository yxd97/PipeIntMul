`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a6ClHM9WGnpz04/R4TG5pPDXBDsUmVmh8Ogrrtrfc5OsXuY5Y2R0VccDi48yVGra
QBaJHhX7plRYsecQkR6iEkm8PY61foSNsMQzt0zO/rQ20JupxAqrqWP5TALX6Z7c
K8DtfnhOjOSWTbQrduKMIf+vROZjPoKMgcswtYbrQqX6daFwynK5Dk5gyU/KyzYl
QmaHrin/ob8iTgHriPHy1zy1RWmu0UtdFM/asU8s2cBgid3PUJCs+EWTt6Xs1zdI
Wb30wlLZWU3tJFM/2pRWLjS8Jpy4JIS9z0CPWQcTG7yevCVQtHoJ8tk3xqC3jrnG
ml10NxdCpHlNJuf38oSMtbnLn3MSJ/Nup5f5YY6GH/yHNcfkzHl0rFXacW4nit5H
3gqb47r7iEfkQ8OLH5YR/tv5HyObegxyrTf9coT9Zd+0Jp8mHg2DKAT9zcw/EF2K
sFFICG/bXBywaCDVHRvu245hmZPtwh30UQwUvuuCD+rFe4PeTeYCxLU3QfCCp9Tw
ntZx0de2Ok3582zW+hylWRPVzywW0jqwuq5X+3G8UXf/21b6piXsCBEsQsv6Ut7y
wNXO2JYgDZ8tc/PynGTLPYmnck5xRTyjikyFA86FChA=
`protect END_PROTECTED
