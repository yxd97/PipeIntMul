`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zun9DNHexCK3QmvKXc5SIlTvRxOcyy+3Ld8zzup8yLNFhjgwJJ1O6CaF48CmINNz
vCPqAEqKzhBFgvrUJcLXvEoMsAIfdkTV2yRbmCF0KAkwLPr5kX35x2Wdtqen6i//
4k0+/bJ+nHtVFvRxBfSPrgRZJXsscIRUocyPlTsh+h+Z6BiMkO2gqCIcSqBbRLdX
phu0r8fWuCGwFjnanD+M0u4IZh3/A3f99WfobAHkOYj8W/fgn8WkfrWkTNIWoqUN
lKexmTXpRUzVqHoBT42qd3PA+l8rPOOWRkuuLUrnnEeOlDtEd05ns65hHtQA7zEk
2y2swPXOee6DWZtclVnllkvIc6/fR9L3At5Fd/lJoJkf81SxbOvvutgdUidAE7A2
czeQ9cmBjllk9tiu8n7KKqhgQ9mGofTevQiYR7kGxsmSbmZI57yrLTFr61cPSOgd
H5mYrSw1mD4y+mUjRPPpIy5eamT8w8wJxXUsTWb0NqWtCt9Nm5vanXvbk8of5xTb
xolTfWQ/B3qmIFHAKk5o41w5Req9GmY5QLGrPIbZBjo/MpXwPNp5MJgnFpGLI3sq
+qlMyyJRzEgkDr5mFgt5IvMX4nygr4hIkscq9SUhYNeeCzoXhXadKr+xwLTU7u1e
urXeOpThARQ/vvfAqPPpsEf+O2nOi5WP6km/MCViEuHeCfQW8EIbsplNa+6zJJs+
89CIyc6FA0aSS5oG+Qd8xPkOM/2pxd74m3bpB2qGZvY4Y082AX13iuKtu9q9F/8H
Adn4+uS8RZW5PhyAeUm/k3QkZD1f5kyA0RhAqhljvg4Z/XKxKXWbEzmDiPwUcudO
ng/LL1EtwpmCMgpKhBzMu4Qhqo2nPkyzStUMObpTKuHLhkDC4u59BOnusXF22jr1
SPuohKJQFe0CDfmICMyWtWJvBnXhSKsoN7Dus9l7V7PEYHtnNljHrg1uoLLYw1Cf
o74IUlF++Wdsj0WfNNxklyLZfJW737WpjYOB5vL49+gER1fUIXnDgYia5ZY3YLOR
eiv794LewG4GWXUy5j61J3JLTa4xx0lyQkYSvY3lYvrB9MgKJLs1Ek6XP4movoeZ
nip7lrXxgc1JOEcZWbz3ElI1hwBYmrzRsjyYpbuNsN7O2ArqgY1HNXV6MJL9ZZlB
FCGA8/ur44X/RxVjqPFPQq5OQa1zGocxpuDO1Uotn/ZEQ7eGEzFIUJpqwJ/DmxKO
94+3HdSl4lkx6YsztCncUg==
`protect END_PROTECTED
