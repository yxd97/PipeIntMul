`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwdPk9lhEf7QSP/BzRqPnsu8VzFlwuoojN1dh/UEsf/RDJ2XzVS/1w8+WqKUnkL8
fa6VJGpQuZu06fjMpXsr/Z1TEyaqWYiGUiGb1D8ctF17AbP4jivTWoYDCEZqX99v
XK/BMWj2xHVIV6SkYLLv7oCH7Lrcx8nD1BxbfDTeX4XMT3PDH09VFaeMMFj7z4tL
zi/ZEWkfG2KKj2pRex6iNhTnJzSnLTJW18CqfjdWneZzxl+bEVJRMTfuyB3GRRzM
//ozyRQ2oPvmXnE42vnbMkdf1Tr5E8S+mLFPqPlrn+W0n4mKVHWzzLiyv9pSTmpl
6cUgWeEC0Q96DrwPk0R9AB+bWXYxVGLpR+r20Eul/hCPncBdt81hbPZP3LPKS43e
yPIvnjrncK/2SuJ8DUmNZpOVz0lGjRVpnzU3aUId35n7Kh2HLBwcC9ntTYdB8z+w
4D1DbrYvN/h/iyiy7lUzSw==
`protect END_PROTECTED
