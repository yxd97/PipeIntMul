`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6gMxwfIJgfKI9JGlSGv356hG0ZOLEaeO+p7XsbCY8PnUTdGItuR6HYlRaYUgj+KP
5p4jkuNS9HbCGkxSCXF5eq6m3zG1yNY+aQ4sYGvYj/mRmjpvJjFPMHmFCqQR2MjP
4wYUy/SdxxSYTWdnchSQBWZqBMoqbDESrDAxP4pLMUdZtVZvucKUilwlizbSg1lR
gKxhtUK0iA7qwFwVs5pyR21sYogiM+Ry/nfkIrD8IYmMIvdpy3FMO544XT7PC7qL
3N17gCdKYWk05H47rvhPQzmBu0bp/lhAZB6AVo+chVHkDHCDhJx5ie1GF2fLij/3
P6Pqj+87ugsZMXB0+kvMJzuJpf4kUEaI28cXjEpjcLUfvSZbGCep2+pjnmqzklN2
EU72hG3AT0BVV9ohYCa1NAUo+n/Tl7oYOwudEEQyGs8=
`protect END_PROTECTED
