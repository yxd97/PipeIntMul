`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwXCMfXf825zU+vennSVvM7W8dAjVFAKK/9aiIC2jPIcdh/dd22EHBOL17hxzYne
VUW+ZBlx7jui6RAyQuK+iF6zzqASfiuQeOYgN9lMa/bH4ZD0pNOufV1s56PDxafk
fPFNJj99fcyn9fyKYZcGhLIkklfFnDjnCu4P7P2Br+WeCSZpBi+Y/k98rjLps0E9
8sYz3SEaGMpQVhsgXjLUxCXVAAOZe5HiQ7b8e42cape44n9XSRurGvkAlGo/wlDA
sQpxRjpk6mZJwaqJmZp7k5I23nS4OXSIIVHvKDIkXiS+f6yN0dCrmtsUTxAlbAxM
fPk6gqkpQPWK0KIT/UjZYtYkTbRd4cViRxuQaiiyUv737ndHdqxbI9Chj+4pF3vB
P9JyKN7XlOZ9+n1zAL5AzUNmANF4DcvK0EUMgIb+sJs=
`protect END_PROTECTED
