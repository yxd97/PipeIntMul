`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0PksE+nz8QgFIuOfvNWtHs5U4RuF4kChrX81V3ycmLOYucP5YJyG4+QRhWuI5sZ
h0Zl6sEenzx6sVHNwe/t9fAQNsZM0MnT01XjnhRVG7HUq+jw9adM9nkvAVpnyvkG
0z32OWzDba+bdNqku3gIu72LfdeeK9l6D3H9kgmXq7AYxF/jo8m+u5JlbaWNb9PM
9Jzm8usUO/CgHhQyJZyi0o3tK70LtBs64Gd5TxPRDkDD22LCPqRgOfjPory527wc
`protect END_PROTECTED
