`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JT/1FZ4zS+Z7Sz10PAvXOHMWDuER5uYxM0d17ZOyzaz9V+wMjSPOXQfkLCZFUa5o
2n6dzwn/jhCCBXN6HWw375fKMzOVZ/KAmFRkp9nlet1TtOCOzmBOkEgDU5ePWLtN
5dVbnWigoS/cnSBV8VQIa9s63JvjfDgTsfJvZvP0xW3WoL6NOwPQeHa0GOvruOb4
kH+2yUCkoWD9neU5rlzEDVTu/VkJE9SkGIj/pqQbu6dk2A6oQJlY/ZI63eAL7ryK
Sw1Rwpj0bgkK0VBs7TcnzPZs9PDLTo3zos1DjBkVKM8gCDI9u2dCEnl+3Phr9RJq
3WaGvi1QeiOGFi0XIuRautBLbPetzfPOVFEA7RNjGSjKI2Ias6RVjOPv4FsVQHCs
9D+G+6i9GS89Y0O2npTrShS2krz6f0DMZ3VfOQkfizI61za5Vm01R03h5aS7QDjX
`protect END_PROTECTED
