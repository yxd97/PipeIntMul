`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Whbl84cikwVsqvv7nm+TEBwHamKg8yB1PO6SVN/srI3dJ1AKayL/JczxFhWd9yRu
OCVKkjY9gMyGiO9nh61Sp3XC/C6z+zCYCA00N4gfB6nkhbotB4esvvQV9zAUUrax
kbqDf761f3EUjCKIuL/8TSzpvRyN9PqG7D9s4g6YCEjRKIv9ageKLXJsBp3n1DtP
QqLtq6MBIVcyG2a22uZg+Sk+SVGP8os53H9PXIaH/IIyHxrUD9gAuBHzCzOO2zXZ
/hTYKFlIiHN25p61HHZT9I7pzGRn2wlUDVceliJIHhEvpJKpsBhOk0TsrQZsZ982
X3h1RIo3K/l79OykQ20+ou4MTHv11b0PicPnaDVYN6HHDdhj4XHP14dgHynHOItN
3F5irPMHGoRbdn46QfEddHnmFw67DzN+54g3At9NfaH4bC3rbLgFxPGwp7WbUch6
`protect END_PROTECTED
