`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdKCwyUnYItdp0bMgRsC6BJxiD9TmwX76+dcezYGXCLN4IYRyFQ5/y4MUvCFHxCE
7OIkd69v33YkaqwGNZkDCNYQK2F6l2AL5OOeRBG+tRrfYjeil6NP7QnDaiDfbnER
CLflMGG7j0svHGCcK1TNmULPGr2EwDMuy5zgcaPqwNpB3bpKUAGrTmFVbrKKX49w
mvvk8yz2aY40hWk7rh5AhpGJWxLSjw9IV2DWe+g7elXgb9KWeKbRExUP2OE+gcDm
Y8hPTP4aQxO4UNcYY0NSLZMX78z98jxiuHDYItsGXeabwCpznTrAn8ulM9Y8bVke
Eu44I5r1cuZrZVwyqJ4CNgkZmMT099InKzZWIAZqUTOyxM7qTffN+Kjqb9PS7Kmz
`protect END_PROTECTED
