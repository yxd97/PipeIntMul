`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CWIRtuGF6XidvHbeUo38wmiZ/Tq24XD+/jXQN18AGYcmENaNf2+wl0Oj5VvoOnKz
wAJjEwgtuYcuOdf9Q3XxobwpIU3ETblrsenRw3HQSvJY50U84ED1/9eUDQ91YTD2
+2XYpDISmJn3NpxvX19PhsoVQDKadcHF51U6ggAaDjpP5cDipxnwsSm2E6VjE12x
isP8OeDQ+TwsAAHhZ7pqeKEQgRfgGmbGd3NwRaWMYhHvZkzy9tSNMth/3lfUSERH
kRncMiQWNdLtJkyBmvFQ0lVT3pTbOsD4dMaRQAmF/5SNAgmUdb2xZfdZmMveYF/T
MCJSSYbSJmn5sPvlcaYgrG9Uox6mAtAXz8NV4q6jOn0wkAC7iBKaD9GmuQPXMFDt
FhlnICQPOC9AQHu59PsR3kvdFajuty3K/Zu9J6cEPmPRjVjp+zjZWZABvMTK/SBg
vfV+jbfBME9JmZ2OmiDBAQL5i/XBrlW+UrwR0tiQ4DBh9Q5CbjgCv44Y2wd6Jx2t
Pn3J0iE/3VdxdbfjvG/bhPvPqVAQcv8uD8QXfyF/uxK1hR7G8CPFTqz/cQV0igob
ic/5IKFaSh7Iu8aD81MGaBi4td7gTC/Ij/LN+WNdA91RDmoyxdpOz2HIiV5i9iEO
kqC2yVNZTOMG53RqNa8ma86pgeRNRdjHNjLRjNrSBBH1ck5rcndOCB9w6qxyuZip
ykcf2DhfJl5EaCue/3LQhqEE5qc7CNGd59S9ylKrZ+g8aKRZ9sS4mWbLPUhThbUC
AHjUxlxpIqMNj76yhPkyodkMPUrXsREz8VUpO68zKeNqczPFIRJO5sPu+q3hjofv
f7E1+YrzS16gegOtjgqWzA/JGSOwL9HkMvYqYKIDeS0tcmItxsxhpWvtMg/QIDL2
eYFEgWz6dhpNSLD4bi3L+SEKeEqDbHDMYkHX/iuN+uTohPsEgF+Dyk3dDfvCjkQC
PskBQR8A2QjbbUejhzs5NO8eux6TXzlt6zMW3vS9jgzT/yJlrP3dYR/4+9BgXE8f
T5KUMfnt7E8La3pUBmKPZfd53Rm/ab4qlpdrdyd7vJDY3xqz7WqO7zBIMvg/z/LW
iG4Jyea/4rCzANHSt4QbWSaPrxj0mozhLCDo/tLLuq3Aq2nAN6ZpN5a6o4f98ouF
/8euNGTB2rkqEbgNat0e9I3a/OuZp5GrO9T4XIs9QWedYDqYgGZFO+kffAEJJIfY
X1MvWPzUJiI+JPZ8bHzysnzV2F07ANPDgF/3jBOPp6givzpgZFzR+WVI3rz1Dw2P
m8N+W6hyT2JwKov6lQpPZ26ZdeZWbAdmbiKB57MVWabMoYXAc+q+d7s84m7qkdBe
EVaUcxTjw4JHUQ9/Tsk+tFZCXnrBpZJqz6Vio94XVMemvZIXaCz7+Vvq1lwJi9dT
OKEK5UW3js6WUXcJJkyA3jc9RDoEBSo9cqydIQpc3wT3d9BIWCeXjczqiAzSOtC4
wJt0o8+ytCHxUltyoQxZwmo1L5RrF2fDXWxvCLZ0D76AMO4NkWtv5G01FDg0lYeJ
LSP45qnJKLzapQ+iia/bMsnHbw4zyApEK/WK4pnvvsfTYtmBps6470/IfEmzZvv5
UPIkTUqy+8acq+W8c1/jdN2Ks1lenUEqmGzmSO1LO3LoCqD4tG3wWITOaISbWrEv
pR44dnpzCiLvOm7xR7yoCoeujBWu0kPJaz8P4Yl7nqGB5QDVHwkf9PnXgthP4PV7
RLJtVF9Fj6aLnuoVVALq4JTmNnC2G69iWGZgO5HpYep74/TYx/nnBMRNe/xk8RV4
gswF9vVtGqVaqsKri57wSMqVLLM/UswI19P8XRNXg7MAHknqMDSqBf0EWNiOp4UR
ucJpaw1dGJyBUYo/ReTxi0ITrahTxJ2GyIgFVNb15RphCaYTvkgPc6oWCnNSLZDT
cUZ+g7Qk1Vj6oKlZSFLVOl4kf1WVPrMDgPf7v2s/GrvyNbmY7Hq+sVADOspMG95W
f4lJQfkTQfaOi4qZd5atsdwEpCYbCFI/ZyHDv6jLH3rDxR1LFtE7R0Kef1CvnY22
I3TSavaXlq/a2kjVRuWWMj3Fq7Y/FNB8HahAwnpHWWFATKxuNwswbZLp1hPeYKdI
JLKfvEouqwZ7PS8fGNk0DUtnVIdEIiTnmqHRXGl+M3Snqb/ZNqOhMfeN1IkUInyR
EvwpuN3WuYwdv3o5GUXUT7J3vfxxbEETkjcT6nTLdDmAES81tErI0EPMbd+TCMzs
ZKfI+2cLAZRS8ad5PU3S7KqhlrIpCoKyqV0/DypWmjNSMHz95Z4PBzSgEe/awbal
k0I47ZC/AlvgD9Dagy6xOcoaoS6/wkLegPKpUeZ+P+q/tG+VsflXE5+tN/yvGMU6
h7eJOKZmkEzU9dYvGhkMMZmOEQ33/IVYx99u8VHDY4ZHuHavWQFqX9OrQK2pDeU1
vhjnPgt5Q542Iu7CZ5toRkFKTbf8exgPJqsrMkF29lXuNX0m1tAuMI/S/Z7vBYYb
eChJWIzB3DKv+ZhfpFMHseOEBmc3OtHe34bpJn70p7p+3RBVlKwgQ6EuWHQn45NI
n8+e5btVoUcc4HX4pKu6u3VktgVYlbuIs9CVbwd6oOGbslxi3tTe43VDSOoihReX
OuRRQ6zHyXZAEfB4gTpiH3PdelZ6Gu0pNzVFlnQbtqLSP++RQQXQcFf1U9BVBZR0
MJqx3HK7YbqQqafPASI7uAI1piZI4W4ZtKj7YlCQ74E9zwZBvtuyEXHn8z3TaSzf
U9K5kXuqom6unZRaGqir6pNx8RTfYHcMbAT+/PVvKZsHf1ur2+/mW0oucm7F/WEk
CBsWS0Y0D6KIVZL6uUT/hcZGuG+UNyvpgNNAzfYnO3pSgIcPFpyqJzTmKa0TIRc3
p2ZZ5HbwU8EsydOyL5i4F8Vyj5Ts/4o6FYxgeTLZbavNLi/+gS7HxvqTOnDPKoSa
5THFDdO0PFCY6JMVe1zxminvNGzQ6PZMUioMTp6srYdRmx3EWcQwh/xPafsjJWoU
tlRh14AOt71cNmRPVVGKJ1Hx/+Q3ZI4JZIvpzMkvwo4dWnzomSxc65uyUGboe1do
VuVCdIz/b+RyJnB9eYe0QIjCSDa0rh3DmVwzNZo9Um+sImQrtjrpDsnvmzfXHVaO
LOEfyajOmbYQsPWdnEDtG3MP8+fshB+EJvoJk2UB6Bc6I4e9pbUwvBM/MPGM7vEk
EBJ4xUCVF2vP56yxTH89Nxnz5g0o4ajVQY/gUKQ7liLemn5Oq1ucZ7iM3ojUp+UE
BlHsTxOWmOn9DY7oDomKRvyXGgF/Ftoo1Ga20u5GTZo+RQCvl/uiX8tBb2pr0xJJ
4Flu9Ka2LmxKAx3+MrLcW25Z/I13yBWjJ4K2Kfj3ubkDxYk0vQn5ngGN5dOUVu8Z
SFukcDKxletojLQLGInG/mEpuFuvtlSx/1DaFaH/ZIcm8JjxxKnFTCH2nUsZt09P
Es/uJ5HQACPJvGHoOIX4JggAAeCmmFCpvaIIc2PVLbJspFLoAaMs6vgZumQ7P4zP
CzLg+6GcHNXMK6OPeqPJNyXgFrNUsxpodSVZePKdS3sXhdrb7pK9XaBEJof6Vr6Z
mqFaetBj/SALh3qJOrbjk4Q0t6wnSOIhwfJ3vit2b5so4scaklKitBDVbQKkj9JO
ei9kDAorwTc2I8vxmbGkjIb1d8wmHmUpkMDK799pFZtznMrITm8NymkzV/sBJpLi
xJhsGTdRl6WcRTEdGIpSxty/eDg95ixOQhFYx1EBpZRBTufC85IGwuuJjiF6/wjr
Sde3ZLlyI9sH8BGSzldnS1+868kzuCovwZzgr0zI1IFhg+Q/opVdBz7MmWiff7tH
T7IsvIfcdBSJfJgY0JefOzQBuJnMUlthNDEH1eby9If4bdoedbjN1CiF34XVOjrE
cnzinpUi6qlONjSfo8Vzy+1DGzzO7ZbpwPxLbj4zq8NweuZUJA69ewc1MSxVYTET
M+6O02YtqUwlxgCu+ycIlCSj+Oqxo4uaFFqcLy3m1wH4wVOEvmtDTtPpO/LCCYIQ
J4q54etT96r/u4/eGvIeWgNS2ZUbTPtGX9u8ax2eaZdj1tMnNHLgKO5mJxEfm+IQ
+Mx1q0gMBeXw/OR8ecvjdQZVgZhGvnP46iblCh++O9WIMFm28Sysw7JgSpxJ2SBV
IrIb9fRtvPwxzc3Ryaph1crZEFmAWQu4zAMYKIPgcSgGF+/ekcccwxk/mJD1e2Nm
`protect END_PROTECTED
