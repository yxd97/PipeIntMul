`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FS/9vZmulfo6SxgPSSBgcqJWsYvKMKxQxW+edfIn6Te+/w4l4+lHiy1bU7PjIoa6
KaDdX01DSNC5kgf57U68VWcLQw2E4GMwIONyO+N2dOj7nXsE/p0KkM4KxlKy54+u
tfMkP5DxaDmsooGJo1OqVJ+OgzXWuQe1/LBaQxYV0lihVBveuktl0jxtjKi8Rhn+
Qs99RfHANuH8nKA3sOIaYnWuQ/SoGwjuy2R/XrbPCffCz6SbsRYxTvWO1xu5eiXr
AGHyz4qGqYaqlWMJdmQcmypkejIcS/kXBpaKjbEMwNXs3d9van1HLZ4xxjMcfi8G
dEu7bTAZ+Ja+El596m+5s1iyzt9sjsP23cMWIKNzwdETdlsKRt//KQ5WuEOvh+Cz
p7GPUgGS0s2GznAzgeWjZwFdGjjNAmAidUJ/mx/W2uyWP9EgIiSr1CnXffOlfRfN
OnStrGxw4xGlEk332GXSawiE86YiLuooAJInGhBJtf2hJs6u5CtW1BCqdeQLG0QQ
zw+V0ohbLiv/hB3xNboqb4Uk3/vDAlFlpP9+h7DH8zj7Qv7GhrRJXl0x9NOJ+yE6
yvQiCYfDAjEwfy3T5VOeyvWCuUJ2+1fcZ2zOeLwQERKLJnjwXkWZmcXMX60Cbwju
XT83VRG9uAdIH0o+UFdGO+R84BvyKFZrW91Kj8+VDAONHh900PKU7SqKTyzMCAiS
9cFEIKVnzXCQLsR1sgFwXz/6av0/vkdTCkhjS7r+g+CQ+NEbv2Zjty3MWjAs5Q6D
Q/tYAKKsdjillUOFU1Qo37ltzYin9WHF4aajBGrlvJyOcCwcW54uJsyzKhRYA2eq
6CP0d2P5ARez6eQ7K0HYGt3TKc+Ss+D7/rPoviQJLkHhX85e4CrNvJgouI9J8j9v
zszeHjwGV4Ag1t42hJ4g/68O48uM0iCoGL48kY/fjt+GpraE6rAgJL/ghMuu7oOM
`protect END_PROTECTED
