`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FicNfeeOkuOG0BeERSqrn6YRCE1bOF5qdlQn/YUcfIXatc8t7lKcDAoZrqTK0la1
9OFv6XoLrhu6UqA57y4rUmE/jBQDdDLBN4JSib8Mjfr00NzwJJ6jFCeoY3st7ko3
KBqsFM387fbB/zfKbZ+eO8SmdIfBakqF4vfONEwfwLP384a841Mad4O/k2QY1XJG
wOW8TpeZpsEAZmnRZo59rWDt5gVbnIT+oHGim/7YVP7TzdVGlPIyfgLG1MaLw8B4
jVs4is6o73uEdQgjODEzgtk4HQJdWRzbfkXcJSckJAo=
`protect END_PROTECTED
