`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cCiEvTZNzbu/aFfXAs762kBV9a0vM8v58GHV8gqmnT0WbSEDkS8/scfN9ETQnbFD
wzYLmNq4z3nzzhYJD1tn6/0pYRdbZxZpzfOgdgHLayKqLqNLgPgmJ7peeNT6llKt
WuiroWcN+Z5cZvADrSayvni1OIyKzxADmK54HVc28TuoUk3chvtAn2FYP7B72QID
ii9lK4Xt66TuKLtowlW7OBCYPYvU397cKTezDIU8NgJ9iKC9ZfYpMmOS4tJGkobu
j/l4sNtJyWHTJDHZaF6bEiYrwdfoAL8xfHP4M3fcDGd6SgWHVaF01q8IeRgnT6L1
UEbLT5UR9wiPZqKxppxUYmqiSIrz8jansljfOjpGc3xl5+EGbNFtyF/M/4Pvn5pq
Io8mt/ZnN9kLxfZUVZOJatMufq/jinatP+43b8mp/ADUI8OchUeqbufI1ty5lz1/
jYVtyHORddPbYp4GUyT2iUtkycz5zbIcayCaJdPY/gmoSSS8ev7DfwWyUq2+TKCC
fLSY2u/i38poKLpNvqiPsUigfHIvhjVDXjheswpoJdourcen2/s59N9N0JTDRnN7
5agQpB/A68Rt7ZDLn0iTmaRsWJFws7YCInPSrRZJ9mqffngT8tsgu32ic4kHQ0DY
GyWGk0IQRkpKCowdm+8LLbnJTMac7T3GVNCuzgl45/Q=
`protect END_PROTECTED
