`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrQ4mPengGteak9EgeLQEYQTEVNES4z869Dgz8O4qu5WM8uPMflU0Xh5dRVlE0v8
o8nwsBqVyDWydQCWoUn7dZ1xC+e6JiHeEAvjDzMT6wm4Zjsy40/o/A8BLer0gOoz
LBLro0+ThHB+MbHPqBQdf2WqoFBF1DjU8cKd7SBhgldA71y4n765NyL9FyJenMmE
eJh6CaKaIEuBEvzVS5s1SaONpQA82ngfl0AKwvC5BbYl5Rlz5Ry0TiLkTjS33ueq
mvZCk55NQve2XB51SpZhy4HTZTicTPiIyxiVVPGCIn7KOMcrYiFu+3ZwfXzwR2gG
0oJF3bFU4CtTRjRGF3f8VlCAOlQw2Whi5YxvxDqme1PAEw3XaFQZI95dYxKJlGXs
JIV1rbNXrMCxBQ90PuGH3/AgKQekNJM4Xy+UZ3RXjKDPblLPCGVj48jCG1PWtyTh
5APGblhUp1HPgBpGt8UCap5FeLkThVSELHZiBJ7DirCTDdM/LgZJUvB/dKbVLTJ7
rzjYkhgLs2M4XQ8Xdzu0rPIrl4vzSjII/SG6bkezzApvtgfP2XgPgCMAsuq4ympv
UQZbcjRYTOPxjqM5KOQaNJd5GrgXWgs0S8kCCJaZ36mg3SYdACuqbFp2Jq7uoeNY
EyXRlHMOmWON3gNy3eE/6BGDgqU+Ejmg+ydYebz4NCfUsz+hN7Ir3yREfwxB0IUh
ddbNwugVLep75fUd3A4djYG6JbEr5gCzjJIg/MWUna0vhKJ6DefNNEXD/+Xpwzh8
RWLIuKtuIK3xjg1hqVPdjQS5gOXvlNcBa/VDaOof/gqVjLXAbrC2N6shzfDcscYW
kMmTMcIbTrR7nN5Gf1YipwW5SdDv3DYFz9DwmNpnX7Eyt4nAUHxmqsDpw5gUHjJi
IChqglatDkTxmiZx4LXowMqyqHGz7Ra+Qqq3lkN710u8NXWaZa2uhPMzMMLz5Lf2
en5+JyUvcNwxVfwnLFIR5LunDCjJLZ4dRI+RPt11MReVxFQWnF2+63R+YqCx4bqs
tjNxGhapRw+sf6xm3CZplPw2x+ZOAnB4Xn37/sph4EgScmW//4Ee0hiTcZd324Fk
SE5JNh4+JOJRgbpYTNVVqle9ocmMwlL9FlkueZsSvw4VCIPyF/3nR7AnCOXDzP8+
HMR/k4fONIGpbzjDXV1cbBi5bI/P9vQMhtiPf2Vg2q3+xTevxapvmxRRvYsPceco
Uqv8JClsO8DsyLnJ42pO01DzjJH7q05sAOJJFAHeBv3K0ArwwmNxxy0Aj1vSm1IA
1U4AMU6BNWPC+zt2BN/Al/3Go4Lf4Z5WSOSoTxPmCA/kqDtB3NW6tfa0nTRAwwR1
vdOkw4zZA//gIBPe94sD9nVcSEuRvGBwBr02cXq+N1Qazdg3b/i0RBDX4H5xeyJX
Azk6mv3qWTAe6iAtEx7n0xJ32b1Ee+WPExo6qN3vESzTMHnXumI4kaphy4ZJAFoR
8idcj3B4Q5y6TPAzZgeYqwtXL2UqtA6CzxOFdaHF7bCyjD0c7UIFY84KYs/EdThT
594OIpgDRVN3UNKg284VsmXdu7P0aVZd6cDfNqlQ4WdkXybQhkj6XHVPUn9fkz/d
6WyZEonJ4xLRCruEk2IzugyVLpo4+fdD6aFuONaLTNqrxMSfcyYpCC8suarl8Jh0
sNOtCDWjYS6jwOJP76E5peCfo/nZuQUrD/aBTUXKhOEELMlFCscqe6DvRcB8yS2H
S+7vBLYIlfu7X4+RCssRXsqkqdIrAzDhAjDNGiduKErVgqtkdJQAdC+P9g8EiKg+
x3TBpSl77xJvnv5sBsycQfzzxjdb8dnbzXkWNt5V33dD05fnuk94pjRWJELo5Q1R
iCCVmL+gwt8WDTdVpED7N+j//NBINY2HQI88ApK5qaVO70HbM8i6bD1IbrzZ6x0R
b+4kVg4WtTQKtuDYUXW33+DUsfiIBjsr9X5+gSbQtDGYHRlbRBok7XkB2wYIXXD+
Bv5Lw2KbbVB/WnUxhbN9z0RffllQIp9b57z/z+U41s4CBjTFUAlCRMnZIS/zuKuS
3vheQCkxHVMMHqZuWEX8Z2vM2arOD7cnM2uhFSOHoYorUwTxEWCEPtcTVedj7gKo
Bk05gd5+scTkqy20hmzNOJC6KJt4Vc94ljyek/5JSV2Xyp3DYsCu8WfVEvbQ9xqn
CEsLNFLkS8a+z2PMnyOu1hEV6qVYCKTMUw/MqjAkBedxhRA64GSCyPP9/Kn1XBZW
cHXOKEoAGLjqikqfSIRC7RIPFFE09AlfKu1iboAvFC5qvp0Ywp7RQAVKb5i5XZJk
QA5fARDLqaEZssn0nIu22mew3YKhW3EmaXxhDQhzLBhhQbZu27vvaM+t3jmT2n4U
oK4q1bEYQ8inKGwitw/JzmsVOSGo3C8uV+1/lkGr9i1Pga4P/NAbEF2yAbqM4vk6
UJU+EZgc9WqQbU1id1Ye6hwaNXA/78KWIS9nQbONwNrBZjo+YB5l4iSLY2i8VeES
gGjiQDGyYe9HpWpvc6WuWB02vAeivjIUAV8xCFID9b76GrAzQzkZlP+EYQHti9TR
WnIkrXgFU4OFnIl7H6anl2psP6Azkos3kivzj7MZYDITEsvFsIIrzH4FC25NcxVk
qNKv07bQicIkyAS09qjbk5obXhXpxamzmO67FAO++oCvLKtuyq3aykisg+FmsDV0
CfUH7Dj3phHS+cpiiypd7WWrlCK5hX73CAoA44GxISByeE8vSmE79KguuyAJwi4M
`protect END_PROTECTED
