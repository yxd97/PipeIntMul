`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MN/96ONa2cIoew5rCT26BdxxFY4a6jfmeadRGtWlDqksE7aZ8UYCI4gi2kG0keb4
Nu9Q1YlkoBvHFK+Z6RrpxMIjQSJbjwVxW1Qce6xW6rEAZPjyuY/VsEBEZ9KgPtna
DqiFWbrmKfCZ0jdFlg8aGIM9Y0hB++fm5f59wEL6+jwmicF00Dn6Sl1LQmCYyvSM
/OmLmvy7x9I3dSg4igex19ELp3wTv77/28GzN9pET2ClblscbWDGt8wZZNlYwdsv
jK2mJ/5XiQKvKoVmqzHNfUqzmgzBxnLBtZCMyynhlwE+u8NVnnFd44Wx7x/2ZUIP
H9FYkcZB4yPrpb36ZAspRlfVUkElmDryVO53dNGBjRTRME1yT+2THoRHlNhwgPkJ
IHdzcTDqSWI3zGlnKf6sq++bkQTYr1GDVJKhm35iHOlLCu3TBauzReTIUvB48blZ
NQ3iT9+EsV707GMC+TWhkVare7e1/OTZRXrZHab6pviZBB4D08aOutsExHL8Rv9U
F6+kzAf55SHYys4rk1kEmUpnP+rTNplqpf15G4K7bHdJEy0a/I7Us33dpjU3B3Bm
pzimqKD+qRgzPf3dJ6nFyzaiED+d9oCJ+aNroDrjEFYJaI4HqIiP/C9mD84lRAnx
eRvDXSQlqmibHW0AQ6LYipxaBmgLxMEtV9OgRBnpYxAYVLTj5W+ieuoQfNYzpe41
xp1+wl0RyZVep15qCuSGsEnlhwYhasiF+CFo9MyM83B4SJP6CQob1tbJiMafYqF/
8oyLq956x0wZH0fAPUmHaHI6lOKTXIAmowju9tYuMWRIszEG6vk4sHrXrc5Z9Pbe
grzXlS/o3QtV4I0Sk36IKP0r666qUFcqmGirImjD4WPNMV03uSKpiaYswM2oMFRi
vAb+wnSe7pgSkF6GTNyfYCTv6ezwRveDo9AJSuX0ZGZfT4v2ECKsfj/5Q5k6FhSr
JPXvyTTzR5nel5eaQjMATlcW9lhiAKGimGgvImDYtOqlGjGBRDn62Gn45oaocaA9
za478EJ9Asxs4cJzbcWVv6XvycWgV4gV4pQzAkC1+tushb7adz7C8ttjqLhwLwtY
cvjMzEdRmC9hLjn2JR6k6k6IVni3KcwKiqF6doBSEQkG4K/8F3lACt5XK70kgIJY
pYn/6CORDvwn4bddwjIMwwxVm8LaAzDS8JmjYWWlRm7OnvH8yG3R43KcRCoTnPL9
WCEWbmXyMh5C1OBvJwBYMWb+DwKnbyreoFKD6UX4TTVxcTJ2gK5H8YHfw9arRng/
ROUPG5NJ/sU4/2HMTtwHHP1PqETmXug3D6rBXaPY6dt76+dI+I1LeWM6WVbvTgr3
yopqWZi6rx2NUNh6b8rhi1zdlFxVikBKZDfe0yUsCYRjDQ9X39tQWPMH4S+GSKRE
pRXK3OqlyO0IgtcZUp+coGc+1dUqjcPSyZrXFmc9fBo=
`protect END_PROTECTED
