`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EVoIO1GBPqwPi+223NcBtsJQUHb6xqHM1IagxLAHBIdZwmIEMXBCG9dyTrzJQHF
OvqLgXT4cUYWkU3YyYk7bmxUkRNgv1M6+cr3Az8fHVX30V1tCqsq8S+MYFSZRQey
V3fICvof1iQz42mrxiWoy4lzCGD3Srm9pU2xKgOm7DdVUp5jeHUbDrcMSx20Y3/T
op0PgmlIv4btCmMZiy52F4Ugz6N6+kkPYGwOU++2cjLw9/dnax2T9/vIWlAU1Zig
r2CM6QYMeEkzamo8ZRvPjQ6n88k5R8EQjWRJNGoLIDFE1W9J03JdDT2cDe1EYZdq
4Wy1le/AUI+XKpZlYKERL9dZlM5jPKofUBT3nuiMvoFDj6e5L937CLg5L89fOl14
v7gs/AygBJw3kgHOtfc700EJn1dUNtnycuBD+HvEncwfAq4qkL5v/3N59OaGTF1N
/xA6nO50IqY4KU2kKehGEHrJMY/SY38h8zc9RlfRm3/z7uWauXYNrsLRwGBnyqqv
AwjUIXvvCz6hCdwl/yAdQlKqqwI4S5oj00jdzyUVG/+oEMudgyWU7f/k7o3/A0om
4MWblJ8TgIA1guPKgdutH+bDUeBRTW5CcQfQUqXfn2YKLZ+re5LK7vDMUIk4f+pz
gjqECF1zTj2TMI9NIVHmeNQaS6yZT2j/2lSDhjpxSrN6al0fLHJKa8py5kpms1zS
bXCtFAJR6ujUyobFeuequbBN0pHQ37cjYrdIStwjnFyRKfts7LJK2salOJwsTy2M
DQ0o0+20SYgjFaTI3nrF1tq8rgdo6P79JifcQpEUUfM7nsAyedlRruNFFcxb7Qe3
qxZK/zjx2WpGPa93qF4/wEMZxq2T5/gW9UDMOm99+v0Et72I+8IRVv5Wlu+kZ89U
Xe3YfpyhlRLKmPPHfDSO28blgSkB9bm6mtdkoH1nWL1FZpME002VQhgdB/G2FWj5
pm19yMjHLM7FLssAUlxi/EgH2govzxSNYKlCs18F0RgeqNdbQqu/wPF+p2nH9f6a
0aaXm8w8e7VdCFZoAkjoKQNHPhzAc7AHrUhH8WoiVJIslXdcNLRAIl6wRYAHXc87
2GuYGeQ+rXl8QgY+PJvIolNNm5134sP4VZfWzDcBqir6Yk2D1J3ldXV2ZlmAacie
GRuz/AGLv2/T1wTjPurxHZyNrLaHiSzlWomYGmwpEsydgS/ry6YMBcpB56eH7055
C6MpwT0luP0OHATAdFSj/oP3co+17Fgn6sZQ040ggvwsiKduoFihS1GPvGPQ0uz+
V8tzxwG35q8t2T4mgvgb1V0MqtSGdfUUKx/vI16d2Q6oIGaracm7GeTYgg0EG2xM
rx+O6430jluispxh8MF9x169OwwvyX87qUsC+sukD7Wavs/oVgd5UKjCVS6fuTjT
R1zwoAmc625E2jNtUOqJdI9loKNuYenfG4VqL5+lqae4ggwPIiKms6P+WfH2mGWA
c1IC205nkDjpHE4k/RBCQqSnVu1lyLHeLvOSC6ghuaPsjkzc5HVHrxHWVT8dC7wO
TalCAA6zz1gi6GFs8WO+jecsFHr1R69bhVZ/2Grg4jATa1L5dwfB70j3b2HqMLwe
G9cPBW3Fht3iMtLbq6JuQht4g0gpF+PK6DbSKADv7hw5poszE7dNKC4kK8geNVpF
yI6OLGnjl7k7fDzyyTONY/kGmTNrF+QdJH1FqR989ya3WPkgt7OG0r4d/wzBJ0/o
9Io96ub9zzKaDff4Jhes9rp+EVgQKwT70+GzR9gbLXxmY2ng14mvQ5TYlHE/cjwu
XuHjphxLYjunjYdvytyMUSN6AvR2Uwxq8SxSWVs/yyOVaH2dUQeB0nVlmnbrH5//
bv9vRbdake1WkdNmlJyzqH0XtgRYsTb/Twmg63LzX4oaA/Ej/32A2RyjPFOmtGHl
E8OSbWoNKOSerp3xjL9vlYHMKPi6xWg0Vg5+7/ZzZE6oAeQCTZaiV6Txl3Eqy60k
6tCnvFFZXb681+MXXARqqj19Jdpossq0+ohB88KPTlpOE9QBGnTBRgyUNTazu7+Q
oaFRNS63etN9F75/YZXDrkGA1t13syqa76TqHfrdQjn1lnLqllZihQDQlhGxGIWE
dy6H+s+4PELK5y1+TGdG8o/nZFVvgAyKBU7OBSeZ/RI=
`protect END_PROTECTED
