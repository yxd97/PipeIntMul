`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AlTeAkz9vu/DZ1GyV+v6JAkqaHMLaoa9JVndCyugdwCNf4AnXk+IddNLlNwgGQsS
k7Z3HDzvNJap5wHSxcbaf7PYsOM1nUTth/WVjQw1XHDFtTaZoPl+8FPdABpci250
6y5wulDrJvw9PChbeZuTbATkA8a4TRyAQa0p+1nfBRi/+bFLyOf6w68Z146FpjMO
c5Do9K1bivibrvJea/LTZ1OZC5yB4seCxP+heKb1M7O4i/2DfS+1MznrNkHchPJm
n0p2IzICwKpZy55oc6/jq4vomjSQWCCiVD7tSmplLixQvEpBMWsCOyHFk1083ZyR
9pLY0hvlASLtw1wPsGySkmYvKaFS9PkPx5/aRnMh34JDmNkVyLfI56HEET2LanC+
YAHZgXsW6mg6T9+faxi3WIFcfUw0xBHl7u6v9+TmCcg=
`protect END_PROTECTED
