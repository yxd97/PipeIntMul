`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gt4RayRCUyJjI/u+NUwOvX6nJkSREm45UFlBRV1pSUWVuUO0jJZUt88LxzrDqhIb
6FdYQ66FXW28ZcEuXOsXggq2wxx32fZ2+Zu5Q8rLkNG0j8JeYmVSObOYPnSzJSfH
FJPFgQDfQP6FVPXUDgLM6ZXjRGZpxjw+uY6ogV/UAC2BnZoRkXavyPFRsebrzBvj
pJ8JuTGnS+IkYibv03q+PTGSkd5ltAKuUpMvuIGKzvmKBmD8II+py3o9wzoWYGuT
jxkJ2KkOflknYinSo+hw/ewmJKPJLIF8KtCeNyS7vAk=
`protect END_PROTECTED
