`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9iGFI0zrI2hmpm/mdrOTaeHYrS8kUt/v1+92I4DRd6g1xferIJFvYZB40cRJs8i
6m+a7/6hjDi7yvwo16KvdlhU0iNVR7eSJbpjuUVPTn0nYIkKGwxKTzBL/T99h+59
3t7HssWEqBwNXAIGoiyCc2JADZAs1lWq3QWNKFfbFaGuVpyD2DcWLjNlt8/D4AS1
ku2XASv6Eiq/6ortEny9YJfgmAK3W1tIvWLHI47+4T8aUQ86Yil0hjZMRK7s/cuE
7raEiJMpfOC5486cIZ7MupkwFdQp+DRqQsK+rhi/DZlqZoM7gu7MgcmYW+Fcmp4f
8adSGFno2KRmD7jKg9ASA917fJTy9lxSvlYpbnsyup+XXi8H/qwjy24eJrLh+by7
/EbEkkWaM09aJxiktCaVgqa6NLXba5OXvdLR5REuWxyaaxI50cp87TUSlmuvMOnP
`protect END_PROTECTED
