`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9oFj1/RVmgrDA2kuhwkYCuOXFiqbnI1cBJ3+kszxty+p/XmiLbiRmUZmZq/Gal0F
V01TZ1ESCGAdzK6U5zlyBYkNi8YXoV61piC/orb310lGsVhlI1xetEodkPba6BKu
2tRAJ5ZQlWgcexa7kaoifStreKqPIHFJ4Ceq0vpwl6EvTLx1tlFvb7Eg8lrsG1YR
VElv2StxH4LaVXB//vsdN1OlxfJPq+j5MBGuhJrY6ZE8ZX9q5/n4eRKevlF0oD9N
Yu5f4s1+s98xBseeIyv5QcdIktAJj3T5HnyhLZnKvPz8NOX5YBNe429R+Lo5Jo6x
zekRmvcHzGoCGrGgUrq4w8BkvpZL+5iuV7CsCw6+4gVhw+C4G7kE3X+66Xv71iL7
ORoMGGEbD44cIU+t4ajCQg01+WTOAM0uQRtL2w7oSBPLhk6ojtIHZFhAlnchgQzs
e5EZI+OEBUp/+8K/Sbu6ArgQMnPAJ07bzqzimCDOrpLk57LSo1ETWvY3qAAMU32Y
xYx8dGsBqpVjsuxO/E7Hna4aTlJczOE1XmIJsAYF+3OGqdltTqYPDKXfAI//WhwA
N8SAfP4FaPk2e/ZHEbGh23oNFKlQWrmBu9DvzXbGiblbX2APx8JSK2bOvmlg5oKL
pqRq+MDd4yASkHDiLDF7/TwQMhLJzueiuAk2lmmfGKxdVj5WDB0aqThM5+0fpT48
lrDToOPkrt5dQuABR1aNOGTjcsf93hU8DIv5KxeVbSI/WtleR+7U5MmuE8R6+ONA
7XThsDVZyprx1FtXoQrgPPohue9f0esthq9TcDGdun8622skyUYJznjtf6IS4H3h
6znnj18crey0VnhuuZsJD6tksWR4wcVX9UidhKUdmLJuGT0WsljS3xRImGjzQ+Z+
lGMa691Du2yrucCjtcSNbOFaVZbfutc0OOB/o0kFXYFX73BlWF6byAh7RcFJwdOX
nCu8UBXPESMiQdv+lDsN+8B6gZLWWvydyTSFIPgi+qWCoKVurnB1bdAeIg6giaw7
cg8R2FSkDTZxXJZGiobP+qGH90f0ZSbGZ+Rx91wRmgMLnEO7E8t31/OoDDVB1/av
PYnwwMVeBec3wGFeZIeXJ5ud5IwjQ89ptKI7DjFj23yPyYfb78aqjbN2vFtYAkGX
pH+eZEWWgZ4yRaIXpo2Tajl5d7UsKFygV9GVkTGuSgzGwJhX4qNm9ukx7nijyzsJ
/m7YxPqCEEXO7L/Lxvw9maSK3pGVrDryZE9gnb5AmST5Lj04fmjVfMz8CZt1MnxA
SYyK2ra1RoRRsUlMV6thuNKEwjf6/rVEmfot/2pBvcqoTGrwJCa3Y8F2W9zuplfl
JP87sBSbh607Cd38XorTXG98m67Uw5/VBSfW9iNny7WZUhSkfkuNZc5cAeJc8E7Q
wjaLp+LVmabD2Tw/+gARX4efK/rNsaW8mDFERWDXczWqk9VhYTaBZLQ3hpQeWPCe
ldhedbrWvprdKcSZw0f2lIHRHAXpzN7CxeCOmUvCM4t6l15DMa3FrD4HItoK1w0r
SfERjqQjI9lw2inXzl9yAv9XNqNDJfxCB5A0dExDJSc5v0VTkAoTGxNevBvSUshh
V0Y3eRWbvnkMVYGhdZQWW6d9EYsqDeE2PdzhL3VpmQVk03Dyaxu4lDMWfNk4ZD9c
UJvofIit7YsEPT1qSxSRHzTSnFotpYPdziUEiKsrUMt7aAk6W6b1SritgLC69AGo
TACLpqj8Hb1WxnAP3IkJcJGNSbPACG0quo7u9HebOv/DNdN4z++B0mmUny79Uinz
jXBQQxFvcqZXYmfeZqzqqCHwB1exSx3OlwU6bsYGzlmTClQ2f1jfltFUlKKVCP2E
oFL5eEm0aGjkYR9rYsnNxnUPAWkq27hlU7hcEJV5CcgXVTPyyrNnWdYSblZmOIvb
6+OfZrYszlO0FSobQ/PV3v9ffIVdC7Woe/BI69D71nJ4KIT5ctEJkgO9A90QqYCE
1TEHNBJnOI9SrU8hEsZ177lOHdhIkIt85xWdcsrh5kJhlLZohg24cOhA6QrivmP9
ht2/zxqXPx5Li0AiIzWnFIcbrcNR2FfpdV5BcJACFD7ciujES3S6jbu9BBzoRxrh
ugPO/JG4NBeDI8l0L1z2bMc/2dOgn2E2NTCCRczxuYbzTgcjVE2LsZZSBWxK0sse
XTcTyTQ2mw4GuF1ercsvWBfKwyPPpz7SSGp8+0W/mvsbFrOY5RiELuUZRS95naml
cbGT8SC0M0XvHQmsPG6p3fZdi3RrLoraBge0ODZGYdriB1y+mstkW2vbmjsnEAZT
QPG2sR9QbRqK8UiLfOxLrvru8neKcaIkYAnGU09zagywwPNuyCTRkY+GnU0SD6cL
`protect END_PROTECTED
