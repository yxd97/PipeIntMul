`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OgP0jHDG4Y3VojsXAn0NniSC6FIyMZS83sr26yD+mHiYjwzK18+WrjV9HCpXwcQE
09uyViYKN3uEy6bwFMmh0LEuGkwVtnuLDewOFKaVvpR76sn3XTrDg9Yt47ohYKoQ
uHZZxoAFsVMDIKqV2iMXQnWAhEIGHpoju1+ouKO1EnDW/5fudLYju7tMYLoioW2Z
6zT0GHqcnfxwJI+fpeQC/yf8tdyZES1Q/dRT1kNa6h1zWG8zu7dMFLGOLRM1F765
qV/rj3CknOfhFwDc5h9oMWKOTgEJqAgWcNOmz5YVha8w+u+Gc+LC4ug/1RrMf1jf
mudPcWCe89ICiEFgW4pfptYC88KxE2TxgLwYnxoGrtAvw29l89xrh7k8+D/2Nzrh
RVrCf7xCacNmKsY1qXHgUxqJF30w02gfpCPdGiKWoyNpS8LAsljtdLGcWRhGoQVF
`protect END_PROTECTED
