`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Atmnh0Tz0bdrnw6lhrkB0xQvEg13psrWDlLaSb3uSKA/X65zTvue2OV8X7r6tLx8
SNB3efPXjDoUzoPKgGfYUffj2aGV4phur6RCAjL6F6j0avE4eNznjumjJh87m2SV
aVfCJp7s/ZfBwr+gy1+X+30N21bobV1TOy71/dQYIGgX+YarE/fcsXvbSYUVBxpe
yxY1RVhCVd6D99Friu8LHyJBb+f3g0wAAQr/aZBjMWCuTmKryBUfDEvXl5IMJoBu
a/Rpc0YJr5sRhz8MjvbaRsurFgCSv8RgOF4qY2agXa08kt6sfVS+ohkWl/M8BmoU
6POBVCF3y1RI94Z3IYDWQX+5sa33XdB/JVRXj7TQCumTByPAfYg4HhgG7iTJNe/v
LL4r9O0GJ79X1/Y3tLf0dWAhB5g6Bty7IRqQG+Mv7XuwPgZFh1zLz2JWdFaxMK/k
HcMZneU+Mwmb9rl394eby1Yq+LK65CbpDdaSUTZcchKjwbkqZMNdtdqv/qTFSETd
y+miIekV3LmThz4s2kVwubDZ3dW88HiDiuI15ssGpBB4Ngzmz2SuiPZz+jjKZnpu
OYfaHbr8a0dey056U6jH6ADBwklTctDtZrLx0TAdAZl3PTfYr97aWcFn0QQqz488
`protect END_PROTECTED
