`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BIbs8sjoHdTwHkmM3iggMDJLaM1xABJlIrSkywsBe17xsa+GEJwcH/2e0YLWYp1z
93oizoyjAQEDUOWUfN8wXHo4PGAdb3ICAnY12YUApSdt4U8x2oC1kdjJHU6gIEJF
AsKJS/5P3813sE40UE2lvH7B7D/66G0WrKJxoKmyf13+6Ge6hNyG0tf4tN0nlV5h
H49inJCor0tX6MXyycdN4t+rcCYjp+85Bjn/EOnB8pHckbYJE8JptYAdZ6l6lTqD
mBM/uzQJqht8/2Yi6XHVtpMsfWQVdVoScvVlNIfRaYqcPXuhYLJBYDDYlD4erJCY
EfziaMaAT1CTchgDqNQlfNmfbf6eHQmF5MTCiFuf0oD+bEGLuGlovsIGuHmNF+xo
NF1uT/kMQ92dpxhAE5b48+sxSdjX5Yrtg6rVuj69OVqWGh/jTz+vL93TaG9hVBXG
8ZXporiQZwYxl5yu/ysOPXsYjEzHMyXs3LiteuTPacsRB8hjfNHwGCCErpEqRbKv
ydHWb/T+mmE0q9eIiSmuyFnja03uFYhPtJqiqzqKpoS005Y7XmI0cilxx0pTXd1B
T6cktycw0c7Xc3ZimQFbC2F3NzWoaRNlMXP04hEeTdhpY5ugiIfrIflBkNMWFoCD
h2Lpa+y222U9hukjrHE9ao5IaiQmSqmHXBla/lypEigqW2JP5uU9O0bm0EdvIpU2
sBeKylyDTMLmjlcLQMExBC65QsyAsa3BFDGSoJ7rvU0dPI90BVHLAu/nS/SsV7c9
zNe3sfHdE4WJUgMdbKXr4mMEWLb9IVOx8q59c8WzFwc=
`protect END_PROTECTED
