`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJLDPFh25H6gk9j6zjRRmjO0evbfpT8R4+c4GD/WzdY2rDVipxxV2HMpRuGfK2i4
sQaBapvrYsVZz60t5RlHhQCpuZ3rcf9LPUl69XFy4GsT4ykg77aI087sgRxjXvI/
TTbJHz2DWLxPU1nglpBboOiXvU4WNXH/Ug0Xna3MTr2vA0pP8VUHBKcUMGiOoB1T
Jo5p/VB7yve9K2XcS3mB40nuW9jr9GkOgo0m7lT0Vv7yMcB4VQOdQ0PVgadXezxc
M0ZdNprYJlDhUp1kB7yLoA==
`protect END_PROTECTED
