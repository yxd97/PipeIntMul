`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NhAHyTMH00gUNDboNpikam8hUtKoBZV/vFzuOCkmIeb6rz5mTc15IC+j6Z9eM2kW
Vxq2mLnDrd9c/qHUUGMbaJ3dabgBkdPdsRrAoT6ngiVsZ2dGzK018nKQBJb+alXM
3l1sQHmAAgPe0uQE6o1udOfZGYnulwPCTIzg2Xwjb2UeiD3lJppqM32g4V5coyTq
zaRy7bEHbrx9IwkuyKNXp+ZwKQqh9RTY9B4YDFdA8WZbkHubsao2NomoMpVFjlQs
L5dtyHNQ/Y7rVm3AJEVoPQ==
`protect END_PROTECTED
