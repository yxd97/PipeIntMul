`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fTv5c/rHaur0msb1yxQurfOcuCrrEkfzSYg2jEl2ehxLhdJASWEvw/yeuxilw06P
ngNKR+DiZW+toCAH9QO0ksDMigkc7QdV21zesPFj7nwWGfKjwj/8fPCDqq4f8w48
ngwjr+yv791dhIUpIO/ksvtqJrq+WVNppzDlj+xgs0sMZAkr+t0VkE7LjAdVb+vy
1uVlBBnIipBnsYfY4+NpVj7vxuAObKI8riDL8Llh9bCeiviWHmublXVk5SzFQQog
Y8orNNQa6kJDA0mat8w9Wrxh0aRZXMDd02/OWnDUs7DII6pvteHofvEPhXq2ulY8
/gY34ag56c8wxHErnpjWzANYF3xq+STneOdwc2Oqc9ilhnnkqxa4YxeJAdsGSOog
EzB30dY10lwA3aklDWrs0cpAljKugelVCJ8ga0Z26oJWcV7DgagmdSv0yi+QT8BB
sC61G6z/6dOt9R6YJwKSIbbKBl/AxvgtMtWSRKEyNmZTdYcdTjFtnfqJM2DSOVI8
592l2Os656Eba+Dz8aS43bbg7a/TIXGIS+tV7kEtdQvgNrJFnnVJ92RIcB0Jip0Z
keK26wjIfLWv0KiuCtHvCmpmQG0iw4JUE8vym1Lt5xQcX9IXLC0hSYHkU+pHHtLr
dFr9AzPvSgjdxIDnuqqvkzuwDAAffGWGOU6aVAEiblB8DAX9ylhI811S7JX9yf9g
vef/hvtXrM6de0rTUUthmMHNJT6OtNol2cUlvEOG+jUP7aCODeKdZq51e3diECwP
NadsSckofaTGNEbfYu1yO0lkKJLz2CH7WDoNwt6NH++EdU2gqsPNmr/kt5/XZhyF
PBryjr4u8Mxx+MGc1wAm5VVJGcIULHehLVX+pfBv0+p9ZXQAuK0Dfk04gZk1KdxN
wzRDxwVystmZTuo3YetUb+9d4FFT2rT+TirukX9cn6UAEmpKNYYiFm6F95c/RS5f
7t9NPgksmwigDtvc8uHfhjfJlTQ2XCejTfpHD3jHnRFHxRVIzNBpDuzwJnmKkJAM
aZ/Yv4of3R8EPgsvytw+TA5sYYsxkckMvOW4YW3dNt/pLdTbdEHnK1/07zjhQX5D
TsZ6PNPR1aDHcXgeqICy+ANWy/Ds8ixXVNJKt0MRkoUiDohWUbd6fH+6GTdO5WFL
uWA5wJa4Z1PXCLodurmffl4yrFBER6PgBNCgxHfpgjBZuwep3lcKqVnL2KD5vLPR
AvxoeIFUsyE3DFBdM0ibGc/gEguOaab05kQx8V2W/wJr2sAe++kAMxy/xmZ5PuwW
J3sTiA5wig0iGqdmbsd7SqZZKp0xM8Eq31wNYaMMSpicpaE8fd6liOm5rVWfU/Ev
p98C9YeZSjLuGL5Ts0AKJ5NG5Arl2scLmJO5LGjCHmDcFR4QuycF4Uj+pYswjlKh
dXzAvXZAdmVdCHxAKN0/Wa0thR3hsS8CoTWF7k7ZXa2ADzBdHOPv2WdMStu2Vo10
fFz91ddFzI5qnfq/qqeVrccmZ3fITTEG6GR0V1tB8zMBtHB5vT//PfkbUSy1y9Ur
DM9qHWzxcatj5GH/eish+JaHkff02QrgL6YdwxDXS1pTH+7HXTmD19HFGGcnIiOl
YJF8gMnqEjt8AVjHqRLX2zN/rMlomcoGFG4vAc7NcczWP3NgeJYvysiOHCfk+9bJ
6U9O/Lyx4T3fd1yHgWEELrASHN756ungXCDs2ulLtP+1Dr9zpN9gbQzGfH8quZuT
YuPrqZisxWoimZks6Wvs5o9XffGVTbbeyKfM5nrbI63zbnF7xwgaUAQNUt6u3rlv
4kknEBaPlN0keWzuq33OZgLFKQkF/w0pPc/ivrjKwximqwKyI5aZuXWIlSiwamlT
dblL9eELWrfvX+hkdsbt5t/aV6kXX4ag0CBYlqsfmyfl2Ua6n8s7i/acRgVE9PD9
tgoxluougr2aBCln0H1HyAuRVUUoomd0Gka/lCgj3LbWR92rBSSBDtrRK/2IRRVK
1vpfWzMBccwg8xNwflfr7+GzGX5nQ8reJ2PR3s3C1mjwNiHw+7iMz8cNUtEGj1In
PvSHteW6Xtlj52sX34weiQedaFyoSkaHzO7WqmSM1MOJ8tlA7l0XhdS5dCX5kSNn
vsinIRsozPKHwBq6jgz7m6IiZ6vU7QjqE8HHO+DHwpo6lHt/2UJWlFd+hFECYkGP
uT5TnddPhlph1a/rkRz/gcEC6TwMtDgfc1X0DWJ3R7mVdroZnuthOCgNYk0/J2uq
b8ArirBUwHcYuwBGW+Y14uvQ2Y0xRkiOJJfq99S8XhBTXzylq6R0zSDdbCr/pS/L
h/G/5QeVw7iN1Wjxmu1aj+Oy/pboi9vgU3+PbE57lXhsWOcfUBStPwlOGfKPUZG+
uFg9X+AKWi8dpsbqhWNK5lTg1zgsMnHn+gWFVnLWWXJHVhbbrLcTf1/qvlf36tJe
K4IjT5pC8nYEZpiEfG+jiYfhez21nimdMuoCg34h3I68o4gZdSGIyTgd/KiK312/
diq70aGTA0tdTTbsvH7bqMgb15WHr8Z3hZXKxQ+7UrnMl9i8fbyXJCJKKLUNWd6t
dwTcy0KhOyNsXmXFo+XeglPhBpZ61jwTeOrk3I7XXfR+hk+LBjVx6anYjFfn9tVh
`protect END_PROTECTED
