`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q4Rcl31WQIKo3VxiSF0MfmAcGCgh3NkhItdaniQdmSP8VOsrcJlxcVfwasNKTshf
tiQ52Di9c6EuVwjIOAmsHXveJcThGhYRlCuJEIfL2dOplqLot+F6NNDJ55hOrvpJ
DNp3vQjyD2tJ3CDYgfo8EJ9YOqpWqdz1uMtaMWmmqevHqW+Q3fd5/pTVya/CsM8K
8wG/YCsxweLPXNCtnC5Heo3/JpjesKu8WEiQwxV5AUQgL6W2T6Tndyxjx5cR2c3I
ObsOoeLKNtsfaYl/zpFh3OowdR+wORK0yKPavnQpsEadzbywrTsMer00I3RXCx8M
Sb+/LkuGkDINHjfAo/8kXxxmAqFV0De3YZhMhf7NSG7pj9lw4I67qPyEUbJnAqh9
yTU0Gb2PgUqPW3mgUu6so5/okswcabyzcXI9q1HS+hHmK3Nloce/kZ1rYW7MDctd
`protect END_PROTECTED
