`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wyZINQz7c4rvIiD/Dazfv7oA7wkbmPJgNJN5zMOgyPFQpO0ao3U8EKW97tz9y33P
x1331fAR4Cgcu00slVzKuylkSUkFvJMcFz7GutH+zlwtlOqy/YfbkxrppMRq15+/
4uDzPCkf7RXIMhNXOP5pxd8IyoQv9JjNIteeZbUBzoKHvtzS76jUgwlSUCPxFdFT
x9FCREDIBBNQkICworRYpf0sTBq1fARBbKLX7m6Y+UtZ2J5mpJaKeG2Wk61ENNka
DFwY5M2GZhX2m6qP60unuE3Nm4k791qdWfPZugQWUZmza+S8lI0/u4jWVQly0Q/+
BePebAC8nV/YgGy8ZFKiro+wcKeU0pDwmAoESolhBny4TgK5M9TojPSUwn//1xtZ
3qzVHzNwq5UG/Cc2ip38lUIhfTV2STX5JN+KjMyUUBIy28BrQ/3ql5i9fbIZYyQM
Zt3DmLCdu1K1pcdAnLUajQXViVgU/hHE0UAPLkDs6Lw=
`protect END_PROTECTED
