`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5ZxFvQO3Bv7fDmoFWrpGs8k8U0iYZY3PS5fx6IwrpMsa8vO5+u8Xs1uMeRmc7++
Ay3jeTzQ0rxkRwI2upjyPhSdCtqCTSwNs4Q+lvAq4VI25Qxq28m6Dmp1kHtiT3zc
ex7m1kKnfWdLDP0KKZPSQ8zen5ySzCMaXq1/TItEPfl6QRXQVmJACfliJdhpQYx/
k5x/mxGGYYDFrU4NjjmPaLRz031dKMujtctpP7Vt8u5K/FM2Lx5+aWQgjWIaxqWh
DK+fnE0vV/zAgtaEt2njgF7bu7Cvs9ch7KKpkEbz64DzgXc7YKU+L8GzVt1oxpcp
84iA7YRZepxLuJ4wulxSNH9Z2+tx3hZkmx7SWANI/bWgNQhLQrdzDYKcmJsPvlJi
t4sk1ab9WY/c5QlRYciP1a9FtMDm6EFkrOqtqd7rZmnMCux2s1QJcQbW/gP0qczW
XgybcSHeWk5D78SsDzc0/kEy/DYQO2Tiq6tW2K8f7dGEUplgSphrgCvTvda4n7JT
dBRBUMH67e0utBOc/fDV1yxZaqovFtJQBGm634e6Dy2GRpwgTulV890/fu0/7ZOx
yijMTwsJspcxff0NmJcqY/5839ULSrr6//Ja3sIfiT0=
`protect END_PROTECTED
