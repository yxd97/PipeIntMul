`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfueCJUWpmqhMTUVjGwqbWiyI+htGb+smZAEIP5Pb3d7BolRHtqLHJgOmUnGUQ4F
dTxO/s9/jl06FExJ++ztamkHA8vTSxr5L6hguVzdzpj8QyhXc4j1HKSi5xXS2nlO
a69LSnWONLGor3Yh+h0Z8v9x5aOeNmJYdZeUU+QmosSk8KcxWHeM5hMQ/kJI/S+z
kSSY2H8H0Zxv/iG3u21BHUKe1LMAQLbWFfX/K/vB/HaQoTDc2I8XaB/dE4vJBPbE
uawfgVKLV/N1RVuSVEfAhNP/f1CQwpQaI9PdzUo9NdYT1hXyBwpJJbQ9BdwAVkbF
TUV+JNunKIHpk8Al03FKOh7CHkVSFTE2pgkYD7XTaNCJP3VqMmaRuEuCiesVETWs
VLnd/CCtaHwM2pFBe+qpZw2I1y7jDhP66Hw1KGEOFtqCQxS5Rev6abNevWmLHrTW
YLV0OS42uuvgmXvDxLqWgMK5vYj859roLIl6KrDaXMoFYDJqAQwngHcit1BNKfVy
5hpxMfT3S3gryjyfdcbhqA==
`protect END_PROTECTED
