`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u/6yFet2eCmwxRtnES73asZrkLgDMK3JtQnJpcowrFuHWcU5tq6Fd9eLCSj7CebQ
ezasufFXo6q7Kd2kh36KhvM+CAMeA/xu4upqoXzaZIWkoLIqbYo/wfHfpSoZ5xPs
/aQ19HAPAjal0rNZPJubsrnd7oJF0J0hiBP5ENSOlH+pazoGo1mLHYhx90NQqub/
i168998ETzI6Uyc8lCrFTnv0oWNNj6websnaGRR1BA66br0n8Rnx6NWJIgVMDxpJ
uhWHLaUVqMtmV7D499vzem+MQqkIKmzAqWCweoyLCELXY35cJuQABquthfMi/kpK
OMvaa5r5OJPZLP9AYk3vR+jhToRybVv0ONQBrKDu08o7FRy7Hs1F50c/ErQxqivW
rc0uLN+O3KbSv92vePGxq5USTEhwGcFb4kepXr1j3st5KLuqGJHLOXnm/Bf61KxJ
pPy7LfC1vk6gUvRX+b/Pt8zUpczdEBpa+1JuaTY9b5M=
`protect END_PROTECTED
