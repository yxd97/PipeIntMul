`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJ6kd7wqa/eE39W6WRg42LpOje8aWCDyJS6mRV1MdQ1m+C05xqtFo2ONvQRHguK5
sZuaak2mk0etApxDZcLwg2ZxO4pT+m3aouel7rS0P/2jDOBj/NL+gIrDffIARiG7
AzkLYmuqHgHT0pCFhYN6Fm8BrwfdS6M6VQE+49FurRuUgq+WKRv0DW5o8vhcAPjs
BEYuG90eiuJ7qXXzODwv5wq9R+DLh8/BhxTvop2AavLa2Fz7NFV4ppcJlyvH1w8t
i9XCt0N6HXquW60rM/AXDLIfuhyWYbkgsxPZ99UcedaBo6WQxPsUafYmbGaQw41K
4YXbnJAKO2bLCXaZY6nBVSE2OJ3hMfwcKtRdFJAyAePxBK1T1inzYrcGy+ci4vEM
jbganPrh+Ue2jgDGfTBEPqGlAJgMEUEYHhDI69m8Fms8hTBhDx6De7qrqY6n+GOz
zckIL5gamkXqrg0hhFzurN0TWmIlqwjMkJ0wEzph7z449n54z3kxLl/tntGpk2S7
rxHl84OCwIF4eLPUBEgfmsA0uyLco9VPVTgxUAT67mzM5qPx3NAekNRybiS3gj02
fQCVFBspOCdV6Bqh8foPwRYYnFI+5xxiQ6B6vc+4Yncu8ZfiqUYKBZtHw4Z3ijwc
omtWPG1qsXNQ9DXoZTU9p+2+tS4wO8Bwkq8+sOOaU2qiCMLfQ4TaV+MKdDW/XFJ2
eZqKCoUCqFgVwU15OlAAauOUMdwtVlQemfV7zCXNhhrgj0wd1fdf1/FsG1mAmrVr
YL7FsrwJsFOcgMu3NwlChsNACQkzz62668ZOfB8A2wyZ3r3TzDbXdAjb3QwGL4wZ
mA/j02dARdLONV6lnog67jNMhR0Ghu3loSRpTuScXJrOCkgoz3baciPLkWmVJMtC
zW5qss4inL4REA3PoLv0eLwMhGDyw3/A7dpIN84JqV9YYmwA39uKyUmzbvvtiw5g
BUaKXUvs28qEwa7Mc4xxl7Ah0ERKN2doMx3QTpCwWBsHff39tCY7K093xPbDJGSl
0aYh5y0PHNTr5DpkEpRHMrmsChWTfek6Z2APUd2cSdHGeRH0b7N2+jj/SJrnSCNg
Z8EFymdd/Sgma27FLIwO6wt1ADHLT6pDKJdkzb+zBDgJhTgdK1D+Tb945d3rJy2K
`protect END_PROTECTED
