`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lDUwic08aSNAHy2r8NzaGUWiiu0gVihQrBre92PepbiCkOO8fbOtkSjQELVAVSTx
yiTelESzwXg5LhU+rmedo35AjZaBF0vHnHj2+OVFQuYAGdBTuKPnmCgLJaO6inA1
nlUoSa6p8QY7Ec3f7v4cblDG06I8yer2sdYnjzPCJR+2KtyvwPO74CdbhkY58e6k
49mJ5ybKljA18+f5G6q44W4oH4RoGhffeewI1ASDo7N3sbLKnfGM+RjfZP4auypr
517GZqEYXrxJbxPfrVs1dw==
`protect END_PROTECTED
