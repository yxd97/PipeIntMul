`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wncyMjzvQJrGrD5PhI4DryFnxmoluXMA6g0wGcO+hnv68xIXmcfbvLrJklb32tjP
/Mdp5bzz/BhWc1lU0yRHkurM+ppS/UIvtPm3TCiwbHVZ2XeDCou0UQSdZ4yDQ78p
rX4w0gb1YkFrBU3TiOBK4WDU+j5EA49N2/6X9TM7PHdYRWcfnDVM2ZEmFJxyAvPT
cDmqLeyoqaJhkmjbat1ss7bNPlQMSC90XvbioLh1ivPRy9urka7bCqtdB5wTV18x
QRo5Y+b7LetAoVPgvqw6oCZP9h50/cCt6O7xAH7VF/lGoleKrDIAilawq6hdidy1
Hfd8ZuhSOgTxTeMNlPIUelYFes2VlO7biRfeZ6WWSm2uKSnJGbwVJDpecpLQ2fYi
x2g5oJx5lSUTrTb9X7bp7NI0U6z9fyBC5c1DyydLZf2MtjJPsMgQM7CE5hLvW3av
pk+ah9ozwe+WzUcLii99tXBT21kTEHkUyxxZA4R83CJzBVRRvsjg/DsFv6m1pK82
e2b+6KQhb4ljMfa+oMxu9jGbHgNPgkN91QhHy7lSoZw=
`protect END_PROTECTED
