`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HlcjPZvBXPLqvF20c8SAit1cf66bynwR30P30+Wo70O3EVBv3pUgmlnyyycuBYwK
XiRiILFDfeSK6S+sKjsVRa+CEWzvA/Lnrkf0bpK+ZhiqlgnBiNpjAoFka7fj5m0Q
J1CN5XxZbFKGoXwyIYJASRUmfJpL2GH49WwWnh2pU4/EMONIEiP7K8e0q+YPuLa8
mIXS2IVEBo6P3ycXnaWNpCxd5uSo77TtKXfeCd5c4HWtCDewwoy8PwnLOLPd6/BG
tVdG4TlUR8D/BguSn8pg+DJgbZl8L7jrzZ8xx1yrAoD8HjneJhXLcEE8u61C5l6/
`protect END_PROTECTED
