`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXFmlNb7i4DX2W5+jYJoeU4MBp/jsiYA0roJr9sMoe2oMLNZJqgMxaF/ROqYSBC/
ms7699rvf35DGGSfyIZLX1RhRXnZo1V/3T2A1q1yVbXYSIdLflFbWplR0NpwfktP
oTwdcmayn0DA5uEGt3VM/E4/RtXrSX5pUohaNHdG7hVDVwmqRysT60XmYlUAfdY4
ccTN/tG/pdeqvclswR2u6Im5th3LhRnRnpNZQHm9C78nw3Lu6Kgij3B7EUI7Weg1
wMN8y09yiJnMbf4RI/1u8Q==
`protect END_PROTECTED
