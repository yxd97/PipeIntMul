`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBm2nFL9ZKrjihmbP12JQx0hPH5K8IV1XKAbIPOGTGjoaaqn5ep8qcT90Y0wxGlh
qQmux/Yq/+gWiTRjgY5XsAeqzwM2QB0fyVRbcMJtZUtS4lbRUe7iSV4dYngUlj1f
8AD9PhDeO/sNvsPMHGWWul06y5tb2A6XmeFrx+DSjmIhMYic8vpHJ1fEjyqzQqvM
kzSQ/fsYbm697meGtJUnj6mCDANwAPOol4ALJiCTLvpoOlLF0l5oqCgovrCYii/4
KWnzu8G5lGc+4Kn+lOnIIZ2cgUDWZYSOPIESZ8mWu/PtUMswTyRBxhvmn011yoGm
r5cr80cJEBXX2E84vcjlxRv5fHZ5ZYVFf0eaZNg+UHnhnvmKX1OACQhkbnsFiYXq
vZ4wV9MYG+STOMiUPJnFi3YUVi60aY5qb/BH+09PROanf/ZzSwK9FMcBTaRGT110
hi7/htAMKgl3H35c1/spKlYoqdsh0q3lLWggyGbYKRmPKk19AHZA0WQN6ozNGhW0
LyWKpcthXMX6MEjP3be9kcoa35ko4SSgy90eyowHfyrLGNAhxHaDhLnaiUihXreq
7wfG09BSa+SaVNkbCwyNilkiQw62zWex2roqDGx7DP8RzT8q6nB98nnkS0fRS9Xo
n/b/+j6vhWhpo8SJBMoMau620U+fz0kBEP1hxyJoCNhl3sB14hltqlNmf/yloyQ2
`protect END_PROTECTED
