`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a2djdyqNGOeYYUGNaM8Jg4aSdM2lKTVCZpXFuGGogshUWspWe9mnrq5iF5ajXKw4
yUQ78HZ1N11ivdjBy3YmVkuPxTW31eniGPrppC9E460kfMHT6SXtby7yXO+uiyhW
umDxPmLmimBoeV4eaKkaFjhhFuD7gVc5WYVIeGITmmutk/4MxVsa7S2HY9EdAF3n
pDJQbcF7ENxEkG51l1Fe7MfEehDg2puqP1dosgnELe3Fx7DTr5NfuCup8SotuXfk
y4VHlBgr2TfybmvJTl7MsRR3yWCFXwgHuWIh6otMOI+rESSC8ihK1ysjlY8R7fxl
FPfzlCraw7lWXzUET5drIQSF6Pvwb6Fr3b3lCleT3lKVixPO0Unz/S+I96LwD4e+
jhTiyvib2X5fLijre2obdImFZNaq2xD4Gimk1Uv0oSOsRVdv6wLz0CnvRbZfs7Ro
1oUJifRb/1ibIcFLnLy6GbxIHwLjNA2gfMtpZI3hZKjxK5b5JQMw8bksHrDyrvyW
/J+V8ip8n8VnW5aL/74hsuhBoglVG8gXM4OK+QI/5HBfafKLhx5D5HJihiMm2G7A
ZHZHEjLpNM5rJFxdM05zuXFucluJ91eHF3us2DWyMtGK9ujI3Wv//eH6KuS8ah5T
s/eL+pXkVLBJhJc3I78Fh0Yz71FvjXTD6a4yNvxFzqoPnHi+PFSiURYr8dIV2boE
wakjc8TLotqEkFcB2F5bUA==
`protect END_PROTECTED
