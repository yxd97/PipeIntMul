`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVljaoBdvDdqQRXONNS7nqe2K9Os0UIPRKu6WMHyP7JHnE+NIuDEWh06RBgteQ8A
9sZ4Kqh5wqGsEyH+N5KSt+zMMjJC+zz+LeytiIjj9Cn7ZE/LKDjndURvzXIEsI0B
D/F+azswm65KuavP+/ZLSIORGYqcUD5a2H7zKtZoDh1O2FDHzB1iDCgbSNqZVl5a
xGNaogfnjo0anjXZhm7yLGe1Cv5aUDMBMiQnw8ehwWTI5xVXcM5MmpuWvIAjS92X
KhABlhQymiiutCq4tqdc6jhbUssoSbErlmUyFzKByrnDlg0S4z82ZIosDIo0B+JL
DXnj78cS6qf3R6iKVfaJWm3+OeSqz8LAT1Jw+POeMdv+OelV51oCcuhh7oFEcbv4
ryWv8FLWP95w1KD/WhtvJQyOd1Y77BCraj+oB+dZQu6qe6fZ64BhDvAniJK8Mdg8
`protect END_PROTECTED
