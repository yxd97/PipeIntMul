`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J/Oi5KZ1sWFmxNIg4M5iUDVZw4wLcwHQm7FMtJksGYlMOi+G8GFvQBJokD1aG2kb
RdWohoAIS58YunnW8hWaL0SINHxE2vDaatM88orJMLMmukvXDvKmUBN+uO9aMABw
hsnH2m6T6xR7TwL/EDcl0XdwRNAFQTXgCPBqcWxx5NNcsKeCMIhK/gS3js2frev3
GZFsMT/2qD7VtnqneSKbabSJEdjkSdpOd3qZAWcEXtu95hT+7ZMdV7tX9nZwOCKw
5cr1CnSERf/dthJ1AhEl1edwkZYviOQo64zmajzQU2HZt3EdHHnE+CIg4l8dPxMQ
7WGkg2C98yLnrQ5JT4cd83uXWEAd0xPRDxfp50BW1rJstFJHmAOojJ/MHH5Qz5H6
EJwL1NovsPOygIoQawS1YS5BQLBS3BRc1yVHegDnDqk/86B1zP86yB1aNAYE9kil
K7RmITWTdpRduJuwNVPkhVyIjTc2LaOdryE2hEtNvV3fjNBdZzhJau2DJSKFyHGO
`protect END_PROTECTED
