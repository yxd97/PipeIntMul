`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rSd3t5GS3Y4m+kEY7Cg2Q3hV5YEC37mIcrmriWc4AiDIzxqvF9toVVG2XzQNBOCD
t2VA6NMNpxbMkoAR7r/b1lmpL6loZn40WMIDa9PccTGRFOM03rNgmh6TDCndSsMl
6z90Kdj7zzeV8l3ZFZrAJdSUEvglmUo/v8AslVbWi4SBmu+AOUvLm4C1osNbC2Z/
h2Tg72Zf/lku/jEKbPXIyv70UMtof0zk/irwXQucYMTWGRkhg97poyErsFVyss8R
vify6188pNSNrIDZmB+i+QkgQhYH8kDRh1KA14ZkUA9j7G705NzCx3Uj4ZPth04c
76aHdAs9YPok2h+nEGVgV0iDrKrMdsCiuU7SVDF1dzpqmr7jw8dtYAg/GTk2KGdQ
O0f2SJuwX7Ui4dZZxZ5hLhyQPkzNx4U4B7JWw++xMI88sTQyliHBcnC20JX3ITw+
xKnn1iMpNOVBTloPXYIwWzeEtRDzlVW4/YayLX565otvojX1BFzMnAbzPoAdlBkj
Rud12auNGucxVai0kTv/IzXgswevTfspTjZg9bHPqKoRdN/wCGcEKyeGKKgqkqkb
Ohr5KUro/dubXf0CZw78dCzPDZvCnlpt5WejQVPkF6vnt20ELhjzMD7gfTYmJcOc
QhcVrJ428eCelz3K42V7kQ==
`protect END_PROTECTED
