`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1FrocFFeGNEr84P531cpDNGKZQgYZ61o8yt6c7KMuSFseBf/FepIgQIL+5wPWPvD
S43HctFB/OnmOjJZ7tZ2LoEJ/MCJ5Tjo3Cph9Yjn56tnzdMOxPhiVtbHhMf8GZOX
XmtSEgjcCgW6KNYt3j+rT/K/w4lS3RtCODFH4GXER5Ki+rjRtzNkJDBcyOp5NXyD
4+zTsY8Jzr8RhKbrl4HPArIpJ+6HJUeorLGMZp9yDua479rceQoXJXqy6B7Wbvvz
nXIHQPslzc6lzBffkeDXPJfk8bUk8OEY5sXmFeCvdz7yyDRIf3W11WSTbmN92fUC
N5mO63B13fto8GlTp+al0A==
`protect END_PROTECTED
