`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uJibwHTh32mDsbSczNsZphQhaFJELh5mYvpT8DwHHd4zQ8N9GRAkkRzliRbb7eHJ
Gzt2tRyW0o3DvnjAI2PWYl0zzUv3ulGN10UacGTCp9g4lLzl2eUA9BUBy7J4pwgb
QNL81EzI/04SmxGCL14A4E9CHSkLazE6dLOxamU33igfuhl+jT33oKg7MP27YenS
yweO9ODf2lo6bCTRnrF5WStFOPOG9q5dJVzgc/uWiQdG1o1AvBPkIJxAYzKTij0n
sUlXcAJnpjHxmTNSfTKhwBouwlZSkLvV4ljvLIpvrEC58Z/yswf+//hX0SUUJl7S
pEtIdaJikGx6t8OfcmvjzOUv8EmeUGV6LhRcMKUKSuBLZQdg5xOIb9OG/Hm/nRVK
0Tr79Y7fwuK6KdDFIBvcUVsB5oGDSM8tqwh2JuIYLq+nXVZLYLWLKJAWifeM5Ixo
`protect END_PROTECTED
