`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9ZoFnMYTC+2pBoCwUToo+L34e9EHoFTNpfjqrKG1kRdPwIufFa4kzFLrNzNGMHj
J+ql2V4RQ0wd0Qu/WoDAzNUJ8HuWPPhNBsfqIFHETnmA9CGZ6IzRZd5A2HSbL/UR
4cOk5esUeQkZVMkfsmb+/grI6l/ytImrcvKyf5crPQyfS8SotW57xNgbLY6mKGxX
hHPTL1wM4yqqHqXFYBk+yusE/cciRteXrByqU68tm13Dhdstjggshu0LnVYGG7lJ
mxDTTfXkTKdJWmF+FuDPAeFS3kd92zVLskRWBTdwQHSOgphse+pTMJ7J1ynf7xfF
B3RuRwAqWKdIuxBUzuBMOPq/V4gN+xpo0CQVxAT706s8znQ7UAyZ2xIIgIXJj1ms
JwhnCTKU/GnS3+B8+XD4ho5WlfN34z38IyxIl6C7VXYfKaEi30RiLFZfTKp9DAnP
Xwt82aKU4rSSUTh6zP9XXw==
`protect END_PROTECTED
