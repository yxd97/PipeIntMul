`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jfec0lbK+XdnPrk49MMhmjLUuuzXVm38CcfRTTGiwiA4dksJyYqnyn5/v5gFUcr+
AY7KSgsO/hzvyR/56DhrtbMT4Fcs/0JmK/R5zTm9G7ysOvfwAFbK3KPTuvNhQpyS
XZ4+ODTrb+Cjla94C+8fa72DrMAiH+fWN1LGYlDWSL/wV+K56kp5LjUDe5FEbzlT
gSwB7lzQwE3qA00IiiWOb8GiBZQYAT3lD7kiWjo13MgPev6mrL/fv8/frSacjgtx
LsOWoOjLQKN9Kqk2erImKlCg+mdcUS/FjpQV9C4ak0Rb8pasUfyQ3Q5Qwi/IZdZ8
rr7a3aZlN/6M2aLj5FD8Q0P8e6AQYGQ31PP6GwjXrXIt4XXjolXly+ZT/G2xRImW
lgSw3kyPLdQqZ29IL4GvIxNd1oNb3WQGVhFbFrOfB9D8ZlCwL+xmPn6nuUZAGglo
fesOXJQnZEg6+nbiJYWHruvunTbmVOBaUyLEz42yiyaEFwx7vAgscMIDZutir5VY
IRA+GK3/v/vd19n2K3EJlQ6eI1lWQuMYcswBOKAnYzwhq+dNsCRhUJFrhpiSQSt+
XKfxuazjt0xgwSVoFzC6UickZAo28LLXRnB/4781YQGzGTDoPClYBzbEFrA4pr+d
I4IGcnXFQn288x0QqNfokUua6648K+/sKAbHWHVw1qXqW75mqQixaILVt4Gb0roh
2A1dVcjGM1FxgUOdOirX+AkEe+3n4jRcMw+Ot+Ygr9cyWI+Kda9b38JtQ8uZmfPQ
5yA9mPALrHJZabZAWaaq0c0mcXvPEIpYjcK+qc0+xVLwNRa/s7mY6HZACmiZF1uD
BuUyejro5sYy2xCEzNForNI9qrcjKzjh5iV/MMeQNoTEyvL71lbghdaTaroynBd/
VfJpOBbXfJgiEQaAh2Fo2n1zpKdTNYtxFijJzWs4qBzCMNt2HMznP96Po8ujYwMh
UfM5RCGyGEbFFr+AmDBLRpwTQPsSo8A6AilCRRGHnwHb6LqKHKUkbb5ux9T7Xe5a
fzt6OE1/ls5dcZVJIm2MohytkAS63RfCK/sSF1urYikBX3ukEsnhvBD3MrRL8vFk
aM+2YUZFXfo12dP+VZJ//yHnEnR+I6xOLFbbNZJJftfLV+yrCQr8NCyahGc6xyqj
90NK65+5SphwCp5Z2mIazc2kUhHu5UKCSOnowHJxJpwNI0BWFfjK+WXvgzFANsvi
myaGHd3S8IpoiieB4fuxrBcV0XTe7DzZDGRwe6CYHBSfNrFUD9OQQ1glxgwK1gW0
HqMnId3iIbZ4axyGrfgxh/0+qj3ZpqedTKhwDOF53r3TYbcG3gEB4a/5ccxB2EoL
JiympGNxGx7CS2Qdd3h7y9Iy3E7n5EZZ7wqYyYKkxsghK1CMlE2VRcP+deZ7MEgI
vqd4OBWUi97eAX3GnXQopClXPiqhr+gh7WVi6NDZv6unh+knTBgjDW56OX7jV+oG
zkck3NPjTwXiugtuE4GLkzNiuCk3m73G1JLlKiqfApv0kIR38wR6ol3eV17+pzVV
YGHkJXDVjPE017Wg0EQ1WOgdeOxACnizpuWzsP9Ip/jx7Ym8vV8xMJ7Il3yWQYea
j7qlkSnfWzWpxCt0JGNRiCMuzPn0KTsxFtiOeWgTVfU2c6evFqPUIhetybw4dUEF
EDoCCYRa40DgBXQGFrgDVJ1vUPwzJwdTIe9J+3+rOcG1NTnN4gS1TK0wVbcYDMuO
HMmUDBEdo5ikF39qgXebWnXOqCMUehI8K3Fa6vBgqTx2XRn2jDRwr+a+EjYvQQHH
XgV3ZMyP5QAgY+YeKF6Ezyyptv/1pHVTehtNeLY3FXxIeoWbZpG12puIswBJV9V2
`protect END_PROTECTED
