`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HWIG+5owL2zwS81xWtf0GP187PBR2wDGIFMQa6rWUPdZH30BjS0n27ZQae1N2T/
qCfet0XCoGl/S45/fpJ+xSHUwSil6Wapef1WqA8E0TG5Z8ffKy6mfxLzcqdJZHWN
O1IWIgcgfVe7/qLL5O8nZZlkbUFrSzZDEkLWEMh8xp4BONsXOSguQLkuyZXxz+zZ
EIwEGhSMoS2KRCHQ+Ao0fVi2fxsCsXIa+A334xoLqBYxMD+6j6VXY/C8aeOa+cl1
PSwXI9smbtVnJS3L/AZZnO4OviPZ9fc1d/HczuPYtaTOZXPS9WoxK0bEj+8nVdcO
OIdA73t8VFIeAYfJu5OWR5YaxDsCox4lAP7WaRvoF8AHq97JQITPPSJtICHAhqBi
vnczWmDeP2zGmXaL4EVcedSpcf4pshltcxeaV5k9LUGO6T4ySLXUxp/Gnpi8hhDf
k1FV3d2wOiT2CROgWOVji71I7jpr6anTfwK4DzCLUaY=
`protect END_PROTECTED
