`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z3TyagGcgMgMtcuOM7fl5HPywmIpfiSdxGwsABJmvNcpKS00vSTdzFegKUriaeD9
Ic3TrLKyEWQCRWzZXG7FCW1pZB/pG2H9JmQF9ur6csrOpLl4IPqzzH94qo+uZkvq
vToNOZC1Ve34tf10ksNLOXZUUi0ZNt9WfEGZThCNN+yAxJy125XAWjFcY5zRTayH
S/ZY1NpCW1Q1zzsvgzZb0tFy7F0i6dmeoWqbjkh4Y9RJQ57f/f2gBvIONK13FNkU
FOEMWEoSL2hlqauEIPHG8auTv2MpxCHMcCSM106aaQthsPxtCwG9Kn1J3hkhob4X
GCOVEoiXCUqrhDha78tJYG2lhEELSHg/yOMKAVztExQ37q8r/oAnBXahElDpIQEc
U3YF1oocFaEdfNZOnKLrR+ztqd7ztT+fv4pM/Iv1gaBCIQglMgyHFJLwzzzbBhc5
AbZ2BrhoevRQx1zw5X9RA2bNYUnZS/jfsbkPcaCog/rLJYnXmk110fa+tMmbem02
nmAt1+KgGEzC92YggA0U8iIF4Ri7vzWJqTCqIPjgOVFHVvRH5Bo6ArIhTeCM8bl1
YRL5aXerADeUcdx0dD7Sd5N30Iz2MSTzs/ynSv9i3gdcJ1pQTirH/8n835ebSxib
zDXAJwigfwT8yeD4ma9iR8IrsIM/7rhkII5bBV9DH1A=
`protect END_PROTECTED
