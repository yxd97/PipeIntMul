`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hc/3F+OYPPG/e89QGkvXuNY/aXWvInf28wqC+33NEgXX6WdVQoRWc1OdiWCbAAH0
RJbuvK0fsGoVSSoOzjjUdqa27AZqkNw9Nt5gxejdn6E/Ast/caJ8XL02gQjZHQeH
aZXfxFeDAvGNtY3OmFW9RsiAGbDUeY+PeeDLAPfdH0rwyc+qp0BXFS9wX/W5nZfu
BBA5g9s9lMo3UEiG6cnqCDHULV79aVw+Sd5LV5Rrm6lc3ezuKg6snFsCf1SEYUa2
+rbPtlSvmGmjX8okwxSLTQGaIi7MHja+r5kDFw4Va/KdvuQl4aNP+x8gdbLcL9Ib
Ol9ew6Yq9wc3HNHYGaH9+HqaBEsAJYXQOZFuu8gShMi7ZvKC91nI3yEYcLbgNDHD
EZoeYgyu+/TA+BUoRKdf6w==
`protect END_PROTECTED
