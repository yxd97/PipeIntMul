`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sghUmOdupXJ0mCLHP7xY5d+DNy/8jB4N1l+gQbqvKYKtVzngALrDn7QlfX3QbXfB
m4s0VIqcFM8DtkxyU3JreJ+qxPlJ/TX98kORopAgbpnFeaqaGiQ/27D6uCLdgnv4
Zm2PUCscH92iHuBGaIKFIzfVlLkfpm5qLSIMGEmca7FKEkc5yik1jVF3ZiPlEeR1
gVbFgo/nupj5A9Z2du6Mjz3i1kLEy0Kju8HnOL5CH80gnAcMX91qOFkLKJQtP0ca
vMjwCmZOhQgexFI1VvN+89+6ya/I6OyxKKzVhEF8ipXNadql/dRKANuQTck8dsmJ
5aTGheINC4Qn63wrB++wJmaPtEPgkPr3MHpVqk27MPdugWoBDXDaBfKmiiKPjXOP
M6o9Yrk4mU2Q7MKVZX6X1SyvhRKdtiYifYujLQcdb3HuajWWyeUT1hmg8sI4pvs6
jjrPx3YQC7pVpQAHFLLjHcNWkefMUdNwe+T550YyNjVAbduD+8Zv0hausoz3BnIf
g2sJXkMsFtXEENXbh2Jt2Q0cEPeHutOwaRY+xdhcTIc1JkSxyH9WWYrJSBwK+E7V
XSE9Y5q9K8EwMLFHMrUEfg==
`protect END_PROTECTED
