`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cv6jZKZFO2kCWatLz90jg/U2DZxZNR/bFD0XPyMBd+W+GUlftX+qMDJVNdGUJjIn
r4wpPQ1Udrj8FHOwgxEcAPxYxVfy+nD/HMK4eQQB6SxS10igJV2AWbwuo9wXD2KL
/PA29UEKy1W57cLHYAvjib+H3gNV9Jw8xE5tJQIqV2HL4WBea3AOlFglioUzkFqn
6PsQN7JODo1L8ZRVfwn0ifnHga05505qCVdKykA9Chbo3/xzo8udS7u36jwS4SPF
B7NPagO7jpVOXCfV/7wsvXLR9Gl9mM2Xzg0D8+0IXP2Z586v1DP1ZLvlegr8j4/w
kh5scGtji/M5TVX2e7+45APaCj5s7ONgtzvL+xDqdbgvfKr1FftsUqZcAyrK7/5z
`protect END_PROTECTED
