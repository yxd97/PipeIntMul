`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FNDhlDLpLQVEx2KD+sGKnUPXEZ7gPrKtC/R3CtyiGNdViBxr9hGubyL8yXL1IC44
wcawUhLllBs7iNp8VxI0Bfu6HxJqv+exVtIFdoc8D4AroManGFg1lmvuYHe7LJ4T
JNYTRGTGEXv3SmQCWmpD2utkg7r+WCkMl+duOnxzAS4VirR4TQgE3mYOyaX9Kq7J
tVdjOT1Z9EAty4SK4giWdmaiQjTwgW4LmSPTgdzYRZ+/G8Gsr/FxS8v2aNIn0Nwi
QfGNKVIus7KyKXhW9RwyNxtq5tQSVLz1KB13se3myhRp53YiAKxlrk1ib9k1sDOI
`protect END_PROTECTED
