`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FP3SEAUaeoYOOQMlNKH1sNrEEL5Xsh6iFVvyd3Ts9jj1OgQyenHVsUpGuHUEL4yF
H7zZj8FiQZ0yRWW7ez8LeIc3x3LKoRQkDlpgdkMJpiI+17iR2a096e4ZRpUqCxO6
0qkQhWOE7LtQ722ErScuP4EGItE4xcc2ztgxsxEgtpHV6BTpmQzNg6AL5vaQVXi4
s9+cOMjfRpfpyUMmAwiQmOHnrGdWVpImvVZnVR2SlMtmkqmItliVntQuJVFVmCYH
IhTTNwNClTfbWyQ5RMIcaall5pQeJCHJm9gvHq+Hn3w8059iKgxlgRVXceu9VNjT
i1TQ7ceELBTKmQRExlEEBgMCBDOaHsQeRTrgxpKBgIl6VMjBBUSphdWyXNEu0kvg
NDfWuw0cXzOT616EQaXX+3LVOTg7mSxc8w7ZuHkM9Fu2BhrJJQYTM+kjHXrsaLPr
pv61S+Kd3KBQyHM/CuGf8+g7eX2IXHgT5bxpZ7xyi81mpfybYbrRCidFzlBw4PVY
IjgBYzPxaPDZRco41vaUWTB0hWQgAsiu/5jmqxsUjVdlSlTb5nlpyc1aU6DqeE1J
8ZtKcgh8mfS/kUwxIHOd9g1/HUKW14oedmhdza5dZEy4YpHiJiMyw34N1mch5AQk
RBdN6TScSZ6MI+eMeUqh4HAA4URy7VqZvvMguduwyLY9toyF5Ml+4qJSgxtVXv2e
xM/xhLprLoXot+7CpOdFUg==
`protect END_PROTECTED
