`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3b6iIh73zQ0cuB/CYJcZvFVQJ1FuST2BXOrzTc4PDagHv9/4cclCdPcc3WUfPSw
XLa7uTJhC64KWeABIGopTpSO2TSwPBSfnXA+YrIGkCmbnKcltyQ78jfjnyXtwm6n
wqNCXilgSJSXsixAC1ZYN76HAwnSpDgROJLQj/LrWzjje5vWN3Jsj8mTvpLb+YUy
grKtEqi5R93hgeCA6ZnkH3Xd7ljDzGTdPl+j1989IZzW1oMkA7viscRqXBcWVt+X
ecBAKA6h9n7CQnok0ZAzGOvha8CtFXsAm5HnGWcV+t69Qo9cSxU+pZKJwxi4eVN3
quDenFbGfC13vxbZ4tBQ5Qa1pbpocdyZqaV2OQCfgQxNR7iq80K/w8Sa9k7CSFqs
bXUc8j+3/nIk2f2ZBWksBGUtzcS3cQOlVuraGbl/J8yxELr2pV0+CYIdbLDYR/Fl
bXmvO+mYWsM0vdfF/RIEahRpzPSR74erdpuHrQKReN0KOKRXw/NoZGy9aP7AXizT
ppxFVQIF41Ngqz/eg/NN/n5XCZGz5lkRhwsVtwfvyjohoSVqF7imsX21Zp7OXPPx
kBBx65qZE5zgypdBROul71WPiCU2RLnfByiEdjqgTTcuHPABMZQg+jv8ZoRdacJD
TvKg8WDgaUT2QpmTuUuEZ3IJ9yYcc6OD85picg4yOnUI+yA+GNn6z5RgpFDZlg5W
FCSnc+0OhS/W1H85xWUaMAfOZ6QsYpyf2rUWowD2d0TlD99T/Jc0ffKjKVCJL05C
FXiyhK7cQGSmyWbl1RlNARWth09wSPs8lGx7RF1xJCGLmAm3e6DUGy1UBIBaAHWe
WH2X4o7TSzGYR+GrUFf7G3STd3RFTAvyS3n7NcRPPKQuLtAPO2EpqQtznTqle91C
PR+GArj0UAiWP7zzHUaXVUeYMlkUX8i7+I43DexRDgIwh9d3oGLzKotiwKpF7Yrn
FOhLW0cyxkkOEQ2cwvFCAM4rIk+fSsRc4Aht4GoXCANj5CG+g4yYvb8YuvMQsLXu
5bygwRF4HDf5+77HmEyfsKNkosh7qyjKNbgMYlJu8rEQHy+Vy/0N8iItjJ5SV2gi
mE/aLt54p74AscCDgttZHg==
`protect END_PROTECTED
