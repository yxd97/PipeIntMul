`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gyyjOPBxEbvkWeiEJzORWEWT4tHV12amUjd0m1ZUo/SYfsi94GDNg9+FXOWiRtWP
W3DxXsFCVSmbUKVGrD6JBPemcW1HL1wI7+1s9o/hy5/Jtm92MzZnqkeTWQ/vbf7I
PsOXsAcKAWG4+cPsylgfo2CJ/p0THPXwbU8TmVHG+qK+wTc4eKib2EstfffebsM4
RkuYTBSptaiik4yOh0TJHxR3a0Mfgw/XgdjqxuvGH//HURLPdSbUoqelF1Fh3fO1
DjeSXzKE27S0CiojwsHeOpAlZjEJviKbr8nHJEGo5R+jj6CVpMIkNl9ElBxWeF5T
730Mtj9awAnThuGkNOL23/FjKS53DqgU4QvJ2bcYyZShy8E0dZu3qBmX1FqLncH7
bcJuCZl1r1nNA3tv/EI8Rcm7NODTOMBVa9YNcLmd72LUPBIM3UpbOSc5px3hgmbo
4ULm2p25/7td6r7vMAR9iYhLS3Npj0uBn2WkglN93i9cewwIBQU47GTeL+20iZKr
j1AEFDtujSrm+Rg33AeauYmutHUYVPNDUnT1N95Pd8pzVIui65u+3yYpm78LH9Cm
WCwDQkyM3RnxXwhwTSaR2yGUIp1rDnZEsALiBapCeShegNsyYHDpW0K3ReQMi/ke
G7GNv9fG6Tby9sUi1h8zjCiKW7WS/qWkmJ4473BO5wZeM9ujDoiMezCAYV1MpcTD
sSVusdyyldBHMrgTLO1qNZ+Xyvglp5Elqc9ET+run1c=
`protect END_PROTECTED
