`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mQdwHu9Krynews9n5OaTnjY0ynX63xM9jCBv15dnkE5c9y/ikcwE6jAwCqABgjki
roNASqfEYs0nci/Mh1GGtly+1EvWKdSg5Ld8x7ACDaAmsewHv0wET/LQe1SD8ias
/4lsnUiRMQCbszMN+pWY0pcxFX383V92wF/f3J00+F528Qs2Ae0K3XxWA7Y7zlD6
OsYcymDbz3rrsFBWPrWGMIlZ/pt7gvJUQK8S9sbNGd3tvYbEjnhLUr3fg1lor3BU
y8/loB6KnkMqpci1H5WVf3oW5SBYhqgHZKv5BALPtaH31+GXq/qSeVYfQSjX+sVQ
IFCanTtsMzEz14VpAZ8R6Ooioad5cCBMlpiW6vBYqkWnemr96Mk9QjZ0mn4gQ93M
KdO8rPCKOsQwO4GCJiy2dm5B/Y+s+d5HMNO07l25TUejZq/GTrOX2m6e2KvMNMvF
G7/IH4sZ+ypN4obPNef9gRaywkj8xVVYRIUUci6yQa+BXKqQBVddhjBaz0ImX3kL
LJlg/uQE0PODOMmG29PjE5SiYM3oepFvF0/lFVCp4ZrsL7eR7zbtcvEFtrq+oVID
UTQvyDz038/8ccq6+huUpqRhk5TrwcEQP93liDXU/x15NG9FuhJWsAXAYUY0RkhL
bQhGZ7M0PdMnftY1W9p1W2Wrsno2KC+CSZxzGRSZOsNyjt5aPPsjmw8bwySIjYzq
/Qqoz7jQV7PCGnDTVURKVmGdHO8iR+ppPIkkZo6J7PEqufHCSguVFYnn9bqv0j4f
jtzQGv0xX5Byr/O0UwxSenJPw/i7SyxVCIzHfUEX4G4hiwn4xWzyv6u1txdrdc89
zSfs0T8828YaFz6r6GlwGN5vUpDHyUNc36GCZlW3MWXuLZb5rCYvAB2orUCkHNUy
Q5xDoGxn3qZ7RNBz2NBWHubnhGqrHN7D1kRJ8cG7KBb7pqO3lMGV77PYehoUbOm8
5EZfBVmpIJdhcragONkBfjBPkUQOQqPGzwljHZMOXR+EryDGI9/XY77UjoV7ToIk
wILRBGlmzTq5k41Gj1x18LnzJOIC0vh11veyYmk1IGSpNYWMPJfPtIXq/AY68CYE
sbyct3Nw/of7hQ6NJ9ZjXnYZDpLMTDsmH3qRkMbBlHeMbdx+Uyw7zybUzuKTP+3s
kPzsrNMqtQ3U4TFrPHo/pbrueZdD9XQHlRbhf5+wWGQMkVldI59R0Vxzh9InE45G
m25/LGhmpqb3CRwAi0gcmiSKhd9s0duGt8r4Y7FU8N1QJMA9P+Ivst8DnegbXeI2
OilqPYoLG2vygbd1vppFAYU/qCLrnWRUJjsHzYsyP5zy5yXo5avuNqqKU4nBPHGU
EK8rr8wj5ABZOWmObFYAGhFiMoapoSmHIu/oeQvT2/+RK48kfh479I0tpSyMRL7h
1qyNMp1FeeAQgDeHmtDSB3m5lAj+ki+OJiPB/yFoZ+4Pv+HXWbWRY9SRGKijqnUu
2oCDy5e7tDATgxg893L7dgOW1NUpfpWrbFsyRn9esx6DBREW1x6gEIp9AFjz5pY8
GpOpc050PrkJ+Wqaso4q6xYMTgN9VNv62zEcV3khnX/RLh0YhsqzsZgmWapa0Ral
a0yZAbJKP0TQ4w0iPldk0caBVi3R7W0qXub6klmmi4tLrAlvZB0F1U7tC1f47kw7
LGGBWBgRN6/n3HBu8XCCsBxmj2ZQfaFkG3OJGxUK+7D51Br8FOftQcBBekh2vPw4
QlCu4mXG4Yu5lfHVAvW9xw3Bwm2Azumsbmg+igqreZWX1Mh02bq0m8W7fvOx7JvS
nKcHxfoX47UKpuhVeTjJhDa/RnJmSB5Z/WJGKS6O7Jv4h73tOY7D237C2Ed9Bop6
DsO2p25do1+kSbKTk7/J2mrFgv/czrnA++URqtiy1Btp3v05TTOBQloJZeJIeBl8
jabOoA5kci/hf96ju/dGWamyjVHe3JObPNPVyGxyOnzk0pTZ5xpAt1wjIyHZrhK0
IblqH0+YzeVYYh1kRjgO7Z1hiSoaaitOgevVRss49uvT88zi1NIHiBTRQxxjGBtX
QHXnNHo8FrkjlvATuTR0BI+hUuTQ4KcakU8YuLIEp1sGYw5Yt9YBaxFUwIT9Fs46
3ypIFuxSi3sevVbB7yNUhIw3kB3VelridR5EgSZzirE=
`protect END_PROTECTED
