`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+ZeIiC8Lci8bDPR69ddE/arpghzn5VnWaY8ih4CVtWJdIgoaCwLLLxEhFMyjFhg
Ec6UHIgmzYDiT0h4mRjSgUeEkko4pfLMCPu4tDRQPTFpfLRzXbBTetr7qLiEMXWm
rCpKkscUHD9dkt3QVXG/bxDEscX9JslJClkks/VFTmLH0FjvLVD090B6AshuIhxz
2nogWA1FY9CPI1sC9DIf5mQnMiApzF3wfgP9mChNu0kyOJmeblhaQ3B6G3rlaxQn
obhG0K3F3+4oQMBQ58EueKnaHOp64xXeMQd+OMsCbogI509pVCW1zFPdtLT6sPl8
ZVc3JurTpy/uRmeWVjRspogpq/GuGhviUGhnI6AqXd6yKDJUmqOShAD3Dnz79fdM
CLd/CZWSBul3KRKECciaJcCQfdzR9SkQnSGkB6S784kFlnWc0L3qMU/nUCJMUDxg
U8Ba7+mniD+5Z12FTx9k/Gygujh+wRP6DorR9hFTNDra8/ODH2ymdWmwdF5WmHC4
/yL5wp9Gqn85mhfLGi0HdrP/fC+UDt91Cd2KlxGVVkpb0fU+eFQln15yRNN0iJmz
Aq+v5rOtR4+IMRBGwvAqTbaw0i8HM+ZxQ114BRP5mn91yBfpAh01czmdD6Rk+l5r
t4uYxWZBKao6PDh9oMKdie21W0Nu7gcrRWTxOrhGXblLTX6QzHyg9gAUVdjvdg7l
219a/74iuhhe3DrL/zQ4AIznoD97p8Wyboyh1CMmTlbINNoIs08+KXHSLsz0BRFg
D4g8N+vjhic4TRNL7fofyKNRkYOgG+icgXoonp07OHeis4G1m7S3yzoZqhnsEywI
Ll0N6/ThR/s9xRfhsP7bRVaBNseyUNks/azzJLrY++R+ewOSLS9FklomxA0SE4CU
hKHqLH4xE37jpV0zHXv8TIo9JhQ9g+a3TYFTxxGPT5oOjM7oJglqq6Zb7sDpR+Cy
sj/GHtWghN9DJRZCcGJrNlfxDoptuxEI7x3PDhVkwPv4pqYlJY5LZEBat0egMA4t
`protect END_PROTECTED
