`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+rKgjwTDxN8PqvKiLHVR15R1SaLVZVA9uApmaBIbJXLXC25e1SXEAXURo0qC5FE
8VBsUed5iL/zTqKoQre68aRxNlZO+BQ0rMw/oF3W80PL5MhaWPL/zeF6pX8g2Mg2
2PUioN+qFPdd8/nyv55tpdOCy9d0GNpLe5r6EvNe0rhn7gDU1BhTbSQLfAZ8JdGZ
MrFluRwIOTWtsdMBgIDQUuPDRA1ky8+3wE5JVGuP+dZdghngtGKMFyH8EI7WX/HK
QcN2snZjyhNhXK5RZFo9KATxKSJypkTAlefDkcgKJM5ixxESuU5FUmN1nqN+zoxj
0cAWC3MmwMvMluPTQntitg1xWq5UfPeq67AzwC0HGBYmjIuBk5l14C1GXyMplDid
OYcpdrkKf+pMvbElHs+q9cxfVcuXzmMIVbTiGSy+mNikHWO+o6KmbMbiTJYGyIop
dGg9cMlBVe78r0XeAIznLKgIhov/NFavqaJd54Dh5FA2KWDFspTF0lt0ndxjP0wy
CuA8Vovj76bnrSIVr37A545y7GoTI3N1MLcR16t3djBj90ZRQBMVUvg5jx/UJwip
WV86uzzDXVNX6rSgdT/g5KvSLdPvK81xVkb6bUivSlYSmRGl/JZEo2uMX3RvB94w
Ax5gMMRLLxdnFDjwcaC29/lVuNiVYPMPcSfgw8y63Kc7ZZGcwt8nZ7RRXX0kyyIQ
a6HGy4pSzERr3Wu1UFn0xha2+y97SrGfDthGbuDX9eYd0031P2BgT5QDBu22YkLY
bT8nXI33mISZXaexB1imzaYmioAOUxSVLp8rCmcwEPsETeIre+UjtRZegrmxOhdA
smHusbesK0Ls5zObk5uGxx7cXiJFPE5O0NnDDqVtNV6+fcw6O8HEBuP00aWJSTmi
UelpDsGNQe6Npe5iMFTjEboccKTceNag/FeS0x/AT8EPD1fI7nL7+m80b5qQt1Ga
2Tf7H60wcAEXeZ8FLsagodJKcIpIY2I+ce7CHC966eno5ypWWy78CLDj9G6PZMe5
ot2sh7GAE0BCZJDhxDz3C9NNpSGTt0nW0XcP0NvB00wZZ5SUANNNv9DW0Mk9di4v
ud55McW39BTHjZUANyFwxJq7E89HqDj3EQXhmRgUuyEJE5a1YhEYqfN8aBogDE7G
fQYnG0Hw6pAGJdjyL1frj9RvEuMikap7XyKhaHnfaUOdZz82ba//Ics5fWS9cwKh
nGTG8uyj8u2Ovy0ZYjdeobLo5PE2LCOqG3cKMwFA7KPwXDYVOKD287HAYhIHdjtG
9/XXDZdFGhmYN/PBMxL0dSKwGxD1QEU6ADJoX4DknsnwgSGi/nQUePuvISqLlWPt
ax3bxOBsUZcN7WSayTZp39YSncZbJ6vgjVTMAijvyXydPIhY/IomtvSy9BDq8ZZe
+Gou93ARvfMDN+dj0R7S+w1+jDrzn01VmUU0GsbfVbI4H1/XLI9Kl8Wv2qUaFNtl
ern547/g/8UEl8Az4qNJvomvfA59ItCyMjb1JhOSsX0MyMOZmcTEDGpw5SjMZfD6
4RHhbRXeLJzP8dpN+i1RwwunJ6crSIPUeVY45CwBW9hj4V/+h9V+CawXLEpCRxAd
ctD+wj6dQ8dAg50oh6Aw1fgDHlh68ZFRc2q8bpu9uZDhdINmDrFVTob3SZKOIqiI
thWMTBU7N1Pmb1OFtaeOqKCu3QaZ1o1aaugP4oyKcmUSCvU6KOTRX9hZqz5p1vyn
OMNYYfaqOfpEC+KwmE7MEiGkZ/i+A0orqnKN6O1gCVliudLiNTIcjychcLKJXY/P
t7535XNV1EJGTE5vr0HrCxDKCSsi8JcbbHWdv+KglxP7kdiCNgB2ibStj804CW2P
ApFXgADEoItBg2QlNmQwpHmfdOrMVyOHfC+w+idd5RAd30HB8AIZnFAAtYSN7UZj
oo/21smm/nTHjxO3BHvvhXcom7wetdTgSzcUOjx6YZwe9Yal9d2tmBt8ESZOQL/h
qlJbOT31roDuIIPJ7RbAvo1HRlJqTYV7TEJum6Sv+YzdKGSA4D/E1fU7o5JaLQg6
S8qVSjF63Itr+dH4kTk086aeRvh90c5vVaWDK2LY1hwYA4TlP7BxQdqrSum4mMVp
zC9Hx5gEB0LaqDl5ZVqUfYn5hJ9Ia4Oedq/klF7Z77VfvuBsh4Z2ygZQROatk27x
J4ehQ5dsObeHAk8ztsvVv5UMVS1Hv1oXZCUftdVr10j4GYWHaN7bkFTVrF0nznFc
LO+J+iXKaEDtBTVB1I955jvmYgCzgQ9v9o8OUzFqdsbaAeR4nbzSzGfAxZ9RpiBS
olVRiPqun6s2udk8Mfhl7z0WzGuvJJjJpQa8v1b2LU7yjnil3wnFKQUpsrzkSVSZ
mlFs2YGrPOWFJoQDoVBjpnZuTsaubvEFFhvwkBAWT7TXwcogGThbQh4u9T+iYeOA
pCrt0X2PlgpTuJkaGv+qLIHjqgdIG7jBBDPOGaYYmzBoifY2adkHbdFdT8AW1vnE
ISETRelSx7dnl0VjR7QQCwELDJ9jpbVgYzseXT3Z5VlKqi3tF2G8GG4IPAnWUhxH
LW4wk9Ia2v0FG7o62fJP/YazMOz/GNyh8tCYaEcqtON861k05TyjF7rBz8K9J0Qu
dJ7akVgycPK7wD6en8PSC2WwMyHaKpKRBBL5OMnEBPJii9vekJDYtW3WnyQDcRcd
jLx+FlY9drJ9mxgB5v+kTBWxprQ1Y84FqIf7hHO6GcI2JxORkENbqZisH8CZb0+Q
DelG7Rqr+0spMs+yz6mAzVzo4Z8AXmB8P5hy7fTzRgepkbAJzAt4ktSawpH6Cq7Q
D8lNowoepfLHU9sCwQ5yv8roy1vpl6DT/hYsmwV4XtfR/ev27CsewVqvAhYeyZWB
6AYJb912R9EqA3pRM4hC7IO3oc3mhiDRb9XUz1y/iVBOa81urJBYCPOtyM5Jv4GZ
axglMV3sF0qOgpmy75lhzYo+uSRjDalZUhugcfA7M2891qDu9tl5ZPBOAwsUdY/P
FgmZGGK8MvwIHUMs0IwhsMH3HXx5VS1Sti1sLOG1jR7ThvQmzbEQk+52etLN/gSi
mRoHIrFfkmMi0dh8g03U2vnFUHwx6OP3n4exFH+kbKUegPxC7laBS9erGk7ytrEV
JLqGpU7idq2i2kPrCxotPNggPZeHM6/VkviwZAUWUO3rgJP2DWxZy024CLhIDbgS
2/nXWApFK43TB2HPTewtfdD3FL9sryoEOwGFpOezJd8CmWWS5BC4XnR9/GSz8Dv0
D0wmfZgJtFaaUpPJpW6dqaNzx+j0J6tDt9atl00syzknr9rjo4oNQxSDtWf8m5hY
MS22b1PwJERlEuywWbYPbL1NLFynMQLHAlDp3B1e4uWFCwxlCATNHYAUGvO59epA
W8IuQTSc6FCN5ZjdN11DIJvrT8ps+m884RXWagd08OiKiRxppqN66HYUPLKD1qUY
vHLt2OcWr5idh3InRL9AUJGS8RHabLxYNVkJToB7NwkwKwGHzoRIfVY2uOLxtVxl
IK8qAvgMeFMQ442q/kt3w2cHqDmBSwnBR/vjRFTvbL0WKrrO4FxO8ZQL7Nzzpfcc
WWOiGK3zvrAYTR8b9nGeAuxdmEL4LHuPZ4svsZsVUjBHJMUB8z5IJgW98jqOlamq
`protect END_PROTECTED
