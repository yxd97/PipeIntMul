`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0hkHKsMLK6OeqNplBz8eAn82TSBVJyk6BkUISy43cpzeiVcKRADfi+THU7Oa5PEU
+X/HfJuapgY8+vkydu5EEdQPWEhIYBFvt6CcAiOYRKXheOH6G+yZCzoSnWgpQhgp
ANUauNo1c63i3BaAio6eA4Hl1LJuHyA5BOSkJ+g/xx926ecC+P0MLAS2FYU+9f3r
KFyTkpM2xCIa0nYaTD8PA8kkes5aLZNr8lc/LCcCxrkMsXVLn331otAbLw4Q6MIo
xRAz4xRtAYGLDlARuRiAMWCZ8yis06eqtexvp8fHxsaeIUUAXaecDBFjKHihxg+V
lS1e4qgZsfPfZETBWBC6rQIQlosYcefr+0P9MFGYlBF79Kmqoi+He+JGRU//nJ7Q
wKL+hJAa4IHjJXcF6G58xx6kwEpAYP6sbCgD2P3DjYJ8yO9cBilCxn3M/eEogywU
7hJBPt63JUx7+Q1WeIQeahbzoaapU80EtsFEwqnpwBLiVR7FXbXDlP7P9IyAcLtF
YphvGvonbvRSyi4Qmn6eWM6nXrOj/X8JFfcwFnQtc17slyQGsax//8sZC8QiaHTP
liDjMKXmdlKI0xEYS/Y3RzKw3TW6crEg190CAznY2AeRy+pTtK/eLaQ/H8IRGlfy
t8eKw3hp4TAwZkF3MGMXsipA3THvvO39/1f00KKBujDHBTPAYZKYocTyG5QYNv2e
BjcBzvjXsqqW5Y0LAlVrpUzFryRrnnkgrBHY0ierqLW5qCwmDUN0tXvoVOm0ROYQ
teK1sEQfPUw++4b3RL+1tq2jIQk1oTpHu6I8XFjUkw6v4F9ajoOHUFa7kA/weNsT
ROM7gvP+9MiCmnccWoodup5k387lhu5Ik5sHfJF8z85waEGllqqQ1X7i7u4q1FAN
aT6AaMtrbiPK4+X0SqGHEvE1umBVAAdeaMLAdrX2cUDAXqHb2mbJ2haKdaKHTqfE
W0dg10vQvescG6T4GDAwONFZmtXJtuyopkdXlPZYH0NQDMPDWys/vUe4A7FfiNDq
seHvMdOfg3nYn0YuuPbAXPcIs7Y3LzQo1Izg7w8G1fj6Xpzi3RuV6iPx0Tpfy4GL
PcErSLGLQPzhVLw9FIX2yew1nlpPOHSOagMZI8r8HX8R78Ism171eBlveGor8Ypn
FG95I6hyT9QgTyMJ1UUUTcmK+HoBBw1aCAwvptsAXUCyZK9zbup3xCX/IKzem9pX
r6t6z2bE+C0oJtjvneaIsuX6KrmbsCr3yi7rTeFh5p+C5f5Qgz3FWxfUSMuR4D31
VZu55zAa7ND/DY6oDoCklfyy52xMvym0oavO/nQ1BpdGZeBgt2mnCCQGhhNfiLxH
s/CfDIMK4JvNI2RtYgWApktaMriVOrA1a5G94QmIdF2TZjHFDNqZaoHGJqEeF6pu
Y3IcijcFYcfv/KQjLnHGmEVmScJcTJiXBWcEon0rM+PZ955E7jQFr/LgPdtR769B
qUzJ8L+KG1Ic1fgB1bBwQR8ZzV4HOlsBBCw2HUul7ra3df6ZYdPNIBxphIBwk7vw
rRp2HPXNrTCKYe5AQ5Xx/Ze3CyfgtGqBAAwuscjW+BDRI3oZQs6fitgRGyv0nz9F
xTcT43O+tW7nkU1HXVI6cadFVCI1Ski9MMIGShNfcLVt5EwVzpeX2DXkUbuJrzbF
LyAY0Dox1trIdE85mO4HkYrKtLXhBgNMqO9F2WQq53Vdx5SCwdD1/oImXdYyUpvG
SXv2l76/ib8+T6W+fmSVvrSno14K6IducpBErZ69qzCMB3VsrKfAut/SlMTZc/E+
cEeqkxB5LJLI2m4JVftciVDjqfYvl0eq1qCHoC6t05gJVIJ9FGf8ygZd14+BNelm
k750AJSRAZRJEyOCVJ9A2q7MHm21Zr8tkhK+PI1SlgcF51VeQOHSlgrpQKG3U3Vm
KpvHmQ1C/7p+qDmL3xv0bA35IdJHYiiRtIvZuzjcaX5DJqnNiT16uYd7OIRHAq2V
2kgIl8gB2k/4w6+ePL82waVw/pZjbmPinHOQo2rUul3hlPf2INLCZd7Ei94bHB2+
GSonP5qqxxsZKQF9bVYvTxnvKdpY5paX01OhN5iI5dHZFPWazAb/hDJ48EICAVAl
oF4SKEKaSmZbaGEMMgIH80z8bD4iOhvlnK1rs5kpCPzzcRexdbqyM8nR9ta8O+j6
AfU/7L8cOuAXtlrJqVY81mpnZ65kJllP7/2Zs7AKc1JIYi3sAn6sAf1KnmSl3WT3
YZniFpDN58Kg6CpW6RFsPr3ty1XFKG84brvrD+sZzgS5ujLY/chgdZu5mkqdUQYS
UURK7U/rABXtXZk4rDKuJ6Dxv3wiZOiDBaFSuo4XQ66Hrb5T1NM02N01F7wFL4NV
JqJMDHVXu++b6tJAFi59lx8aS73EmLQvPHuyDEdtYLhJuu6diuVHN3me1hkM6LER
2uIVnIOfgEdL5Po0NHqJKSafMDMSOVhwbw7Jum1NK4rw/W4XRfnPxR3swzhsMvPu
uQv7IdaKdlqfBgK+iR65dEjo6ItQU4QGt/Y1H5Dov++GnuL3lIGE8wnYD3h5pYB6
2sf+PRf+CJXExTZKU/zCR/FNxmVaWsC6f/QhWcQ8hxJH2/C4onoputWPxUyMaW8K
QXvCamyChmryYkc+QpDPsQJUwzZ4H69fUl4lw3abAM+TIdwMU4eX0wACfVaafpH6
vj+paPuHbDhHVEjqafomuDszVLhXhLWyoheM1tVnak2L9Ql3k7XVeowv+Fy0gGPE
+/ptU98LPwXTdsx64R82W3O60lvou4j7yxhT2h4DsU9c1PH9avxfDpSP8cAqsHXy
FHRqKuu8+64RIgNxhleqszXDB8AnR9fYY7FqC/AaEFZZv1UxXM8h2JBSt73VW8RZ
ptseAW+33Z4Q+4Z5UpzOsQNQaO+P5TGRCz78WAgfL8UAMRBwaACD7ZqSOVuUEwOn
vlplb9OtLiaddHeJLX3f4v/v/HZ6NLcLIrBFF8gN0z3slWAfWJXFTQ5E6YDOMPcl
Yx0/rT3FvwyW5HS6WIT9hgWg9lrZpn5eVycRoVSvz1Nb3pwTDzezqMnAyWe2pKzC
I0XoxjeVVqzUjtaJGLXakYYg21HTyPv2kQABbDuAKZC40EdlTskUHNKRfYrr9k4W
fZjqRApXrrfw5aytaL35KguyLsI6dr+j4sWE9tza8pmY88F5Yc9BOxPE+eJY1cUw
KUcG6Oaq2js7Txl6XxH573TGm8u+hCGOpPvnHKvAwxr6QXSfy7x6iirNai2InMOF
slfr6+K5lEQyTRVpfWihB/9yqDgTQ60aywSg3g+HhUbmHv6o8o4ni7KGhGhQVE+o
9wV2g+MHUGKud9XKYmz8t56vC6byyXF8zU9hdqqkbsLwEO/3l0A1Y1cdpcj/ElHe
6u/Qjjcm67EUi/1EhxyRYq5L++MyNHV4HM8J4/kQFZs4rFfcU7cmxmjNXG4WLgfg
zY/beaDyQ0I+bhV1jxbAnslDsSv42LFyW6J/V+ggk6psKP66DTfRnXALMAiSmRkv
w/buDMvqlf387f9zY70i298QxBNZ/H48q4Cl1RLqFaqx1zOl41WKmeIU9lDvHRRf
lm/Ck3ySOPTFk9xmOrcTKHlBXj+Guzx26FoCdbsadqiSb5ogrr+SjJZs/xUhNEsP
5wK4vyk+tYEPnQ7/6azIplkJCrqKsSvtqLtcHoHA+T+/eZYp7RBc9P3MEJlwax2I
ml6fKHABvD1eDrz2L1Sv43qCvDmphRh36TCEkX2fMWYjaULxJVHHdy0oCnlK/c7t
qLYUvgUBIPeZMj6eD90WuNzc1wIwb3CMhopasCEjQ8wDbuhHUTzqNAfYsDOvFLd7
CtxV2/XrrMAbvJcMypS7NC3JCkdARNKtEig0QQ/MzauA0jlI+zD+bgRbXL9inI4h
ty7aG2sN5vwE855Dh+INCTKsx3dOqaGAU0MN/wQPMmQlLDnaWcx89PelpLZ3DaIG
NivHgvPkDzSBStwGhmivBmLmrodV1dKmolU+3FlnGQiNvl6IWmRJq7q+8ZWdavxY
uYteiYuzJ85n+mzBWVF9lo3Ydh+ffQAGyJGoxiO9q0eXYf7ey6E9GqULRqZcJVW3
r6mUAtz2C8JFiuqtMDjvBmYHhG27hroiyky3/GppoYqz2PXFg0+LiLbZ9V3f/FCt
ZH1ZByVuStN99WmFGutOO74+4R0R/iHGkLxYEOtAJWbkEFHNvugyxnl2JWRYIasS
1PIKvG3chJMeD3VDD6PuhJgcaNTMHNpq+laKAStb3U0LfDsirVjT3/PCAJq4lBKJ
v4Q68J1YTEXCzeNYAzHQFf3QxVojXjh3JgaJZbjLLtKXynu1RtZR4CF/C+c0aeZX
RTUpxniBBPie6Oxzn4xfdJ4EQJ+NO6SVgVJlWTzNXmpETfQCfq57sjSsNWlNtcsV
9KWyCZu7945vYA1IDaBARMgrquz+SQvI2XgPxRhnY3U6rCuttY7vp00Y6g3zmEc4
5KQCqh9TlhmVV3yHE18HeUoEGm47bH4LsGA1E/f+Y+Uh9/E0uMsYDZiVPKhtUBJx
6MyxG3O2s8s8V4Sffs5gYjL+iBji1uwpQDJh37SdNE7wrwQOjPtLSrJoRkEhQTSI
16EcLGp+biZc1NwTpKLxhFGfm2v8cGTPyRfNU2G1fu6EyUIq2ik6xJDBEIwfO+PB
x6F/0LI4UyIc3oquPbrjSU5Vtykc8A3taSQVKmPtkhw5AxaE7WrQ3Euec+K+r5Zg
IUYf5dba1DNHhJlRY+JkuqSSMvwUI3hbSp1qkep9uakFRlhJxXGdJzSMNpvAvyKm
dWT33uSoVl2IopMTD3kPCsgB8+lt9SN0mta1easxoziIoI7f0JrdpWFbbyK5yTzu
DJfvVR+/UnKwf+CfTHZGBnbfuD2ADE/QYVrc6ILpje1ZJWMg8H3Pa8xPSKvXvC8U
gite91u0DaPJe7jaOjA+OS6zQq19bRM1O4bw5gDzURO53a5lD64EFlxYPt8pylef
u+vHxT/UMQUsKDaWRvK2swSD1TfabO3kNBYYxyhV8O7+nVhm+pa+qvxr2vTr5pL3
+e91jkQIy/4ZVGCvglqRoI+yJ4eYWm9eyesqHHXtFuC/pIFxLg4cT69uy/2mio8l
rrG4+HMxxYgkhtdyGm6k6vYU8ht9h26ceQw8jI9YY8rYDGA5r8p8dQiwKLp1bpD7
4mgPDl0vElJtxCg1EFL0huSduS57NjrZZeteji3hdThlJRP5N4T63Uqj7enL/mjq
fqLGOovlVPrpFSp2JJkwOfbWUDVQJj2fWarrfwi+53Lis5HH5YVqYEoAxeTTU/NY
N+QyqiDDuAiMPngFMB4qKmNoMcZyp/iLvozi9eyvjxgbZeORiNQ2uT/hQPaflDQS
Srjf4PDN00Sb7B+NJoXLMNuaXP9hXO2ayNgquWMoea26w4XvsrcoLJAP1q4/rTk5
wL62kfqd9fHLD6sht83VNdjbxJVlRiqwakqN+eZxSQXwUBlm9Ld3FRTJ0s/wBzFa
+Xv127kcPJpDHzq3OSh4sbXKYwxJkKxIPQ+aSaKC2hsJxxXJi7ffczBm2WeG1EWl
X27HaPC7rmOZS8NwAwTWWklSY/KYyXknynEG78RmTfPmjVZybxZCE9i8mr0YSHdj
xlbAcGVVD+sxtdkPq93RkrY7FYv53kLSx3TvjGPXJOWiIW1/dAyT58rrmnrfdulc
c3sutA5ZMCX+XCAGNJU9tAtsRhsOO/9NsQP7gTfMnLrehazrjk2O9SRSVwmH+a+O
+Fe8L5ZMc9aDTnWTLcEU9+lfKlpv7RgIXJBV/iSUXUEUk2JXx+kAEIFjUKSoB9/k
misWVI3S6m9q58wVGKXQRt/nD16PH3GGSHSgRbzXjbsk2+2uhKIRVklO4MBrXJXM
/FNYPdt3xbVm0DDeYXWkQef45u7dJSeQIEfDXW3RmQE7FGXc8V4icnX4co2WT/76
wgtIkkwzJSHLmxvO2QzPNHHhHiMH65INL7eOkfysyAVtRNF9LIx6xxKZ9HE0fo3q
Z2/NAIfHE4gDm0TtScvpQp6Ntq7EDEi7bq3Aki4T8D4ic+q7J8ILn4g3FrTzga87
IHhJbsO/F4XYoeomsbGjgl2yZOox6+/xwHYuxZVVN2+WYdeWR6QOavSdvLPu3xWf
gBsS3pLBMrcKV/Cth+IDY57MRya7I59GU8K/kHD7p05bhdH2NP7rS38Sev7ix0nO
Ak0fM+hpb9xOujR5JhOL1C7j5l5GPs4D6DxxS2aEDEXVI9wP2qu5Fz0ZIKi3EKfb
Hdem1rfStO+YoSy1+7fmz67igUC6/fqYAxZQ+EV278SFSVL1teofgEUEkD4prwcn
lLgy3f68+zZ8lcaTb4r8cjDNtyTl3VqBQnMC+fjfoscI0QKO/ETahDDBCY0HASMP
jMVMrmCAW/zpel3GjV02IMGfadpLkpoEcrYvwy0HaZDYzVXQ1bDOqF78DKP2504j
5TTRJwbfmpR6qZyMuwICJbnIEfoeC/etANZWa8wiCg/iGrsyNHmE6/jKakYJ3mZl
qFTa83tPVGzaSDqBd5eRYyyGvCSaw4HU4IiPG08C2IjExTrSDptPRjuEYuks7eFH
ydvgw0T01EpDWS/Uh1Y4TYDkkzbhtpSdMo5YWOsz+5MRKB4cw1AhLzWtUPhk3Kas
vy/2RvzwCB6HaUJhft5+3s8CNUyMJYXjYfi64uOfcrJ3RbX1f2jfo9g+Dk7dUBCD
u4k4iMBVtnQrrbIYD2H9KV/Aiyr7+ad2uFmX2LeGv+QZ6cJvXrzmQ7mc9gpBi42A
brOnLEFYQoOMDRWISIKX1Gt6kkSrJomWXydnqnKT1Xgnj5NxkgOmfcuK0xpddHig
F53TjOGLGdwGgY2hzMqI8NP4HUwKuQvIvh0DfX5dL8nDoq4o5lZFsKoFpnMg0TCF
dWfqX8o5N6i83TYImFi5nx045lY8V2GZFvuGqRfPofsF/JISp73tL6eVzgRcP1aH
mSx3BwnsQVht45cwtWWj42Yb7ir+CfQiMgdxeth3VVdgbOqdqS5x2vcGG0KSjMux
xbaoZxvij+Juq0qrvaHafdk+CYj63uXnetJ0eTq9RPtfhSguehtOkhSSwM3iQtX6
EuyFw9OCMqcQJV0M0hEUwYerqLQh9Ei0j/k1Hh6cHkl4e2YVEX6hxsPleLRcwOLr
kuEo29x2UX4CfxhLXuu0qeUfALUepAV8smpjZ7csKSBMZuWDUCfZ75Xprk6AKF2x
F1lkcDoPNEfHbzko7WfAD3TeeoCCan6xyuriDaBpVSl36+xIiEkwEXLofh5w93L9
CTcUNYNM14nqtb4zHt9UcCd406xKQw43rC+0WnVctbgRKeb2SEdXRP0TcnckkX6R
q4gKI3KtGNEGpTk1JSt1BZQS4N5Dw+VrXixVEcf0tUNslSZkumi01RQWlVQrcowg
3cd8xE92g9dS7JXAWKN3deAKeyTWNnlt1YtzLeuin9o78n0xBgXP6NRnuJwI28bP
mHHFtpzqqpGfODOAGN8fPpMf0QbWw8Ls1Vo5rBufTxECLludZLShjzFe/BVlA7wX
46kCeC61B77EOn9caXM02zgsuwjJVmnOPvFp/zBxKuNfV9viLMYWe18ZZNFG+EuB
w2ScMFbGDZbm3ojtkjFkNmYSjMgU5/BzIwvp+2kDTYgiEOUD7IvDmum1rwy6EnJ3
OkR2ZHHZvJjxhkQKQNtcUzEH52pjZjQcMuTzwPliS6+i/ap/mFra8ifcK/ssmcpN
qr/9fpBG8pYtsVMwtBhubsFFSZbI5/YRcltXl/tuow0aFq6yrpxIGzRjhZNo3WyJ
PQ6Oqg8MAuH+LLrFDSOEF8d/YFg2wR+NZxhapnu9bTGknbqOef1gB1kdzs/hDIKE
eZgTldyzk4wGpHl1+LMFsLReto3DjCherm39etlIZtLHZ+5POzfous0tf1NG2bZk
TSMZ/OFqcNoj+/hfXlu1bNsBYu5Svb074BvboxIVu4q9wCkQiiIn2/ZcUf1Gt2Zd
zM+h9jUJzwHJzSJbNejUB6epK3xEARfFb1zpBI1OvRC9g9/9fzAcpel/9Rs+71du
LNsTHra22bXvrh21Ll/aiG9Mid0kPqv+lYNU7OP30BO6jfEhydmrmjJXuU7pZRQN
IUoojjIebhmeBgAWMA5aKoS6dBNC+MAQybR/lUi0MCcBTj5y+7+WWYchuBdZ+47z
EmPCTvxTLWXKf8w5VxDzFWf7t4OLUEHLCUcODx1RQdgx2XBmgguw/uNZMtiy5+oL
BGLXuaQRJQPYt4tkTjKVeVy8LHBuA/1JotPUImOmRrM3m1Id0Wlc7RoxI04FrPmO
jpC5PtGM9M8o8AAL8OZP78NFUEePCJ72fUmBR38D8MctUDUYyLcF0jhSj4Gtu/ke
gfe6r1wHGksYU7lJW1JFC/O6nGoNAbZlM8docD5VOMavkeMGdpde6J4OHhWPJECW
YID8Z2cqFgXSw0H6+OosRwlWA9gP7C29WvuWMu84RDmOpZ3Zjj8xW9PGszXeCxQi
TQr6wSt8kgC7cN39ooOOlpx4g/T9upImd490w1IxRCPkdd0Dy697Uw9+NcRbZvlI
GgFNXpok6URBefng/fFna+Pe3eZbFJ6eQ+KvLZrq9flcJ9ffu9lmdhbwSUkn6xl0
I6biPP5g4dcvXt9/D4ddnOPIzNhtXtzo0oxHRGiG7r5zHBZuhYxgiZ71VSN7yLJ+
RJRlBPrJ/Ab7wLl8a1Rh+J03MeiCqT3DAw8OtEUqxPLDyOO44lbwkOim3BW54wgC
Y/c01dsfh8O2551GP0T9FL2UcKJ38wlmsf0kPyanAodc14+7dM76XxR4RH6uB0FV
pidnF7P8KCVACAZIRiZGiBHsBGOtTiWJmbKxrURcD6lU8Pkq+9ErMlbWt9/gjN2o
uI30u/XfqYkKTCPnBynrY1/xFWw4Hnj/BG0mnWjXVOHaq3yqCOAEtiIMV+CSAj2p
LI9l5w57LfWgdf/vKoZ44eWqg2+y4ndIisWagKfEkfFYEGPHuzuT78/S94pqKesL
RIKb2zyltwkAWD+KsTiaDsDscywmGlLT9frr9SYZQiG+3e9tcuqdHQxiljai/tXr
NTP9j/Vejc0sds0t7QcnfYAxmpEbsSCu36vhVKc1jHFTNPXPfaFFUkWAKoYijURF
mislvaUIH5TfQ3qWWTNXDmAcjA0meDwikF3InEUBH7l9cJrX06i3FQM+Wb0/qke9
+FPgaUvyEgYXSask3waMuCLWfnoGBwv7lDTd+MOCW9CDQ6IC1S5LexSsDYxsQwtw
C0bZxsB1Xamra5CoEAA5PqJ36RP+nLuUaxN0KcdTOKFm+hriRmV9MIv7omK3wGat
M2Rm1nofwq9U/r9sJdL5q8ocfZoI/trUkqb17TP42hk9HMAJdOy8YtalPgiKWVnf
RTPp1/QNvnpYQC+uUZQeCRxgPvvfgUgGD6M03xQpOzZWEMtFMOMng6gz6kZF6I6r
4UzVEUW7Bqnapq1ngTqHm0dy/Y3OORBaFG+A4XePFIPNd/VyNSUoa4q9QPaptqaA
Cx38WIilmvR6UQisbiE5z9fqIdXfCRokCymvTIf1Hmtv5a18UhIt6FxuaZQTWWAv
0QYtnJeizdjdR2p0CTxUX1eZDC2jWuzDUe0mtYBzoqXhwSd0cbhgmKOQykU2ypOP
hcmxDQdaUEsuUFu5b+EYXFb6YagzHVY3BFspfkmvJnIFRUQ3Qt8e2J56rbhdP9wP
c+D2PwZjcCLV/p/sHBWHOKxE0sUJxRlxb6VvaRVJss5+tdBxKdMYwVRhQnT91w8r
WYGbU5Vt1DHx+V+wB9l5+Pfvzadmfc/2Wc4Niv5OfjrvM6J1JaZqScgDDVyAlLyi
sfyVH3YEVt40mp7XROq/OhZYWKiWbHHQylz90gwqvWSdAd6NYrJBlIRhCtKD2Ffe
iMTS/yEW0Dhf8TzDiu+khFomysZXb20DP9Wkj+/CRJBepOCJacRFk4sH2fCs9Y2+
IFuJR4fGttPdT09IkHtq8dKokRRoN1S7VKXFvVJKpXvmCeyE2TQtDoEmqhCYkLF0
bV2d6KkE0eACAqOOY4KOr3fLu5IVZcOD/Ybx1qKoISOjIAFkSakFiNcwfgKD4glV
ErzW05NRBLKIrV1YUNbNKUoMsKY5cF1yA7hXSS8oaPL+s5EY8u+i0LkOjb3xsnG9
7gZn/AtWod/bRSw6K70R8ZpMJuaZUQYz15oWBHYqtafrr9SVqQQJB79CKOZUhIkq
70EBQqHFisH39YdFb20ZwBcKg7AUzP3Z7m6kv8PzVsbrzs8uF3zzbKVqgIZkct7k
DLu2zeoZ8vOV8vvcAbzuRK5YTN7Vg/fJKbb83hbCdZijNj+/DxnAK+FGvsmY6q4R
g0YN9KTJRmKAWYF9UXA3Qc9CKGw7Ds6+YChispAeJ6XJcMhBqrai8h9gbr32KUz8
+iOjxLgsVQSdefZ8u9or1RlDxBqK3fes2oTCot7bJnDsZ/o5Nly9vxBgovwou2xB
EaE+3w1PIy9mVGZN4r3DWGidJDDRji2eKDqlct85BtuOpxehzZGh+wj0vMjkuHup
SHdc1QdAIv/I+7RSP8wKYiJmlwJLU+cN528TPhnAuDTGBX3oQzsP0TXzPShzBU+t
4Ti3gRoYRK05xpo8pQjzBNXKj2O/OX/dIOrSDBxsfPuLzdRptH+ytW7jiffifejG
+Tyzd2j0Ldy0BWNW86nUxZOo6YUxRUzQW5SHY3WNKQzWU/TkSw/HUJQldxPI1m+Y
lUjQXIMeZ6gFRSQDjU14OFfI3Gy35n0K6tFBDQHmnlw0QIxAaKXZwz8rZeAEm4a4
+H3P6ZGS3smoSATm7vjL+UsTdP7r4DqWvUs8rb9vC+dfTDKGvzXCxAPt5nTWOwHN
usbSDckv9qLFEXKV+NV4QDwlw5yFPBG0gFy3H+fZTXv9hlQ6hIQVIcF35GNIhJUv
Fvq0oMWiMXpc+9CmxRsRh9JOhjGt+UDZh23QfuRVrB+anPx3HQswmZbVb/5KOV0W
p/ELxZ0As2bdi0HQ9mHWbPJQB3vTe87+t8Uedl2j4O0gpk9hiS+AQ/FW4X7ASAiC
CUSsbW7Q+bZDxM3n0E4uIGFBKEdr1H1xnDOkuJ17PJWUNLruO6WiosFv70G2Afcx
t2YsofeP+7LAJVbXi915Cp9cL37JB63fKuasPmuGaBdZ1waTuDVXvfuiKAMLATF5
WB1gCjmPkOw09GVw0YKlBGMmo6MJL+Pg/AGla1dv454Cb3ycrq1GYxnBJY5msdnu
916ETdHrjjxBpPyGhOlGdgaom9jGmtrN7AlmuFQhFfnIaQHKHkKjIi8/1Imnp+aK
b64cFP6Chcu4v52DvYa3gtmiHm6P66SlHuVuDKl1g/MmvvJwxdzyzFfrU/cRqfGA
O2T2OrM0w+w9FwBS9wOcn9nEEePeH1/RgXctzgX8d5QOjwA30bfExGTzcIoWd3qK
3+GExMyPO0jzaZvsiDwR0t+m5IiPfWvL4utG6j914UjziC4Bwm0ddZmi4l44UJoH
NPKlsLYKvJb1afZOSAakbUFXtF8bDWqEX8hf8Z7mQ0Q0MII+YdHbJKiEnkmZAn7E
DZ9OWf+YSB4xl7qYh5TVFFfkF+jTqrZluDTcBWUHUAxJiwqAOdlKWLxOql8PJeld
mclHOAdofVaBsAW9KgX+ocDZlazmvDR8RmfUiGxnWhsyoH8969x9v8pT4Uso+Szu
VItKWiR4K8GeTEYTnTYO7KPpiIvFdHFqmw0qRUq3N14ZqHy3brSZotci8Pq5rzgz
R7njZp7AJlhiPV78Y13cdrX3HJ4ueCnO/8mp5WDYyTJTGN3EK63Y8Dqaxi3kkazo
z19Td7zYYjmYiM1al95blYFtzR4RhO4HcZCQRyCaR8WZx0SwkusiysmLpqW/OSYw
Imq+oxe7ut1yP/sHjVbjZO53qgmgxgTiTcEjA95ARCzyvyn8CV7JB+O647q40KQe
ahiBOYtxqrYkYJXVNxzfYsoZyZyxoDkb4upcRDDL0Iy1NSGMEg7cfuDGTKcgPjVV
I75knIVkmAHp3U9lXtIuAxgxrKsyZFrSHbQNuB9/co9YqnxaBNuUP3G/10oV9kM/
rWTBCp3G9FeQUI3T3a2u2kFAvikt4K9ot0evucidlOhUYsEpESuDT4hLFMuLhg55
nEZ3mRAbg9yqbspktQPhCa8FjV8jilytMVelwt9IH3UszuqFi1aRu/K951CIgdNa
eYKZJYfuKFU5v7oqp03PqiqHroxdEMZDG8sjiCC8UmC06vNdnrcWzHG6ixDJBljs
wPr2RFG0EqHiQgwoG+IgkfGiFyic4UOTnAdyCDOLtHChjfJhlca2Ful73jV5Lt+0
vt3c0I+SO4h9b24OUMyJhkT43H68jCCdTPXen6/nKWRky9CHRzWEOcbdui8bCOOK
GrYbepwQ2kyU32HfU6bLMBSDOvDDsw47TaohSTK2mwkm2GHNOebKyCXkhKXMK11J
iNBf5c7nPz6xV1jzIHusBLM8wTnsoTK5iz8CRkajfGktTNPcNPd1ZtIQyzXjng67
HSKhd8Hk4Pa1dJK60w3H+XvRu/BO5mqZNReus5hxAFSPqGC4J+QKh7nXKPgskfJm
tzRnHhAE9V/qx0XxMrocnBmh2CxxVuxgmMbmmEfpnMJWQN4OgdhemRj9R99mv224
Hc4lPStlJrN863gpLw3Gy/Ub0fop40eSGacDdXcTKNWJg2KHgBiWbT/FQe0Y5nW+
EgGowIjJiGOlvxxZawlx7jlfR2x1XGN0oJYjrGlboXTrkn3FM8e0lmPZY2Gc9mxY
aiBLPBAv+mQeZ758G0k5RYTIdfMxDc7NGyctMjKAxeLGcIYgn4rGLoZlC/21szGt
JqIWL9PZUQJY86pQa6nkq5/izT3TxT5atOgWPkzZYD1DhMu88xisxLdM1zzRufjz
M7SK0KHqW88rNRJt0vgn9zQeOmVTvjoP0GZSgwQO+ERrE6+78g3+66Gnz2L25sdP
fpN9rYv59ylBVOHsScpI5ROb7yg/cFJI84QCmJAlPUKbJfLmOFy9q3HQbWntmDz8
0LJA3WWDvCOiDe9M/j2Wu0W7m5chSQMfc2QiHQ83Xdpbh8haM5WnYkETvlkh4ISR
sFZcevv60679tQFUvFKI/GRaNIaOyTaUTAn9GMjHXtc=
`protect END_PROTECTED
