`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JRnpTA26+nUAKtD3sgomKtIDO65+1/CJjs+JkB70laGZJLqFhfysNTLmRrriz54q
UlGaVpi4QMf/UCvGz9Fi0mOUzDa5EmeQ44O+fGL7n1k1VgRLDgAry3/DMgsCZjh7
XAc+hWv3JiFnB1M/3tsTCwWhINBLMNa5zjqYTLBEPxVVFIZxZYNsm2zchWi9vC/l
bq6d9K3zLuOF4J64N6k+rZrYZhKWE78aJ/XC9nP7jG8yKTpl32FJhxzJw3qzaOE8
QqQFqj5UZ2XR3hiUhqkk+ZL5YDsqa+8CXsXhy/Prr89u0wwBmgm0R5Hz0FsBn3tD
3WqYgR5l9bM4qd9wchFOuA7uWJZZ9L5DXMHL7WFhf6dXBXzJrKh3Qyq+9GRj9sxr
4xHE/0FKCaKH8Ccml1Zoinf9z5VkpyjddfgIJuZvPjW+Tr9qaqMXF438/6dChG4K
Ipptw4CxzuMpl0JezQhpDYsJ9D+wTyUGZAONJFUAj3l6AUNZBhnzaXdmIt4T9ckc
fzeh95nbJLPNELMZko0xgR5HhBg+oP6QdCINJ2IyKUiWjbLqrmsV0l7ByUbE4vlY
833kekpAWI9cUAbKLy9NF6q5ID/3o+leeAnf1hpj0Sm4b0YocHXwJKJHOrlms9wW
SVeQAJYnkH/Pund0pYJnZ3hdCf/SRz+pGxRIgvwLS3SSEsBnJfgpnSRWYcILF9mq
5DnYl6uSKIYekYX0sDjkjGtA1N4zsbYdjmosl1GUDgAlNJ9WDLgRdt9+gJLG2e0m
mafeQ1ZnkQluosR7ZObWo2nG7jd1tUQpG5RnUciwYnK5xaW7HPUDPs+zd1xCQ4Rq
eQ+gUvfNrre1NSazMs5TucpJlNhQ/2HpKYOeZVL4dC/OGQnOrVDV5xJBJnAGZwKl
Lsky5sLlLSyMCPybrocZkLM1R/9hTzU8aSGGNfSg9Qs/2jC3jWZsIhr7ZauvdAoV
F4GKgOsbGDZfLp2N51vOFm3r0HRHt8pzoNz1+Ka2leBXndQ7MnHFKbo5PD59YTHI
G7KM+NyxWJsSZYuipUqiyX4W7G/VLvrgAOmUhFe68Y1rzIlRFsXuyS/ZPt3ei0o1
D+h03lHl7n09kJBhbcyQeb8gJiP6wIk+Fojp1wU6gd6xXUP0S9G9pP3ofOAKt442
QFBeCJX1G6D2vahLYgUiUEseA1n44nwTLmMeFJPdHLgNlLoUJkoU1cROgtHrv17w
TKQKnjfPlt/hH4N1WSCBDDToG6os3c2x/krPQ16PFhmDFm2agWl/RM3Ox0VMozec
nDZIdszKNetREWjl8kJ2qDiyODuusgOwfErqCaHhIPcMXOSzmolkeViH25o5Wvun
UzJ9TLtqtN9Cnu1n6UKPGL1VchLvXpsVSkDITPwaWd/xIUP8XLmoLiXzLIAg2iBT
aT7xgcVZiMWQRYIfTMjf/uaGHPZq2iMkovp1AwBoRng/JwZwDpF7/imx2hDMG0e2
7YyMCmJIM/KorHEI4eAhxVTchtwTkeXqdqqO+CGyofSbZcfgH29ITgymx4c1Xwgq
AhF6UvLKLzChrgcfG7I0llqRjYkDzk+8lWO3lBPH+n3kOMdmrxv13wZVTbXZd3GQ
dZOC4otePAjLd9F+8Jdxn8C7hfsv5d7CQsVCmJLVvVtrVV49ukTcWRAGnI+05dAs
+WW2cWwjplzBdbNeUvPM3jJm8s/zgvZGnAIjZ/XYAUfWg78xUkZE9/8E8UdRwx+/
m1XqWxbm1mJqHd6mv/W+vqptIL5EgY73mLMFE7/wd+63RVqKQ3rE4Xt8+FENjMqv
lhB78FC88UgUHolY0zQahd8++JNE1j+P3hDAEDTmTjH409+hoPzZ7EX7d9p4SIqo
vY5vKp1Yls1jBmhAQOY7oxUIpBoV338ocVxb8pxtrwwrQXtr1BLAjmE4xiH7P7jN
W8Iz2pvi4WEpTR3iiyHiNFQr6X7unGZFxSjwUUCx+tcQxWeGaAHuCa3jAv/RNYse
8fi+dH/ud9VArq7/YLoqyHmKJkPfmJC4egldHhMmg92qPwO/U/AK/nVcMnSskS/X
67SdfCWeR95zCvKnjMJahA8wTCs3UoWnY48VqzOecQQaMlgTDejWkEd51OETUu7Z
U0Gm+RPU1uX2ZtH8QRdLkZFyrnCUo7wx3z6fR1Koh2bqTyOoKwVy9NqYm1rNNMg5
6MsMXzVsryAVIjC6VdYGKAzMMK2x9d9ElzcHGptC3MqbCintnjFq0lmTkObJSNKR
gi4S50neeN3ti9RjVKIJKLxXSTSWV8aSNHZEPw3IzSM7oT3MahyXpF4/xck3gDAp
xbdNoF2zmn2g5ZPSUu11+aonBF641n141ksYWo1gnI9XZwVBFKpI6AM3tZ+CKPQ4
Im9rTZCcEFKr/6D/D6/KyWRIDpXcervQM9wD0gYDJB7kFwAQupxndGChexMSLtjH
DEBTe2VhVes/PqpmZdLsidpkZWKVGtapAsCW/vlC6r0oDR9WZWKs4eK/KxVwfvR8
2eTY9saAweEFF4SHpyCC1+IdcNz/9jhmd3hzdz0oFbZtBog0RJPoNZge41ANPETQ
`protect END_PROTECTED
