`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMBl2nB41PyYH3UaYuoQ4c0YY7WRaSz5M5WMpjdX+771MbRmB04v1OOImKe9Tce3
Q8lU3l34s2LqvnvqE8yUGlO58URCw+xRV3LyWq9OSdsGSjHe+z8FOhtt3ILOuEp0
OxqNvlY2V+B8Xpc9oAp9TMK/k+e2sh84hGyXoyxHVA3Adpf//kSnn8UGkbCnKdA1
d/p4FY6Dkg9JN68b8xA8OFoh5uQSzizAa+7oPz8Zf5lPOgmB+KhzuRA1086aHq34
lAzUskps1KTrtkxt9HmxFRPbxMaxrWFINQl6bFziPxPmyi+RPqc0cGzky0+RiaB5
ttMqspxHbUHp/Ra8jycJH6JzbUWAiwmGe0kCY26qpJQQZQkbonCRezHFmxPfjE3L
8fj6Q57tecda3h3fbRs/NFgueOtWIq4esSeLqdRmLyshmxUozvoPMublSlnZ9D+1
QsYHSIxa3nRoNvd/r7AJfldggHvFwrswBpqfLzS51Mqhej7F3HiUNArZ9TAirOE8
mBcv3YWLhYpNq1jSzQRohyu2VmwsI2TLyfM1zi0mZzbFVtotBfJGVhdtB3tsQ9Y6
1PKWGSAv5e08UV9oL1W9IA==
`protect END_PROTECTED
