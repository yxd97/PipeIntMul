`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ni6qUq1lOQrPeoTAl9I4UZ3uSTtbfJHh9wdPQ3mknbcDZw6ZItqM/NfNnVpQWSsX
ihzP8US4gdrFzElWvsp66DOvp1xtAmeOdpPyozF5EcdsDbVSpt4RRf+RQAr0Q106
7jTBqcuajbkwFrf80dIxwhI4al6z8nldFc0UBmGl9MaAhY+ZdgGGdi0s+DwZAgpZ
aW27fLtKQbQQeCZnirz6XZqD/CYLx5EdVopbdqywCHbDdK5WT11gGJRep9n52D5n
beT3TXfSr63uw/q+k1y4GQXmNucpbjNr1DeKhzFXqUy5PFEQuwaYOKB5YZbltUyR
tmdwewqK5Zc1ydggrSN73XNd+YMxyffKHp+plKV4EaBL3Crb6YlpOGe8K6dnQdM8
O0PjgIzsV8pBAsVoXXx9hccJaiDgKyhl5prgaFO6GBPBNEKwNGq2l8EuKVEZ683e
+BjoVJVahQjJWRBJLdLePUH48CAyqJ4LlqSG4e/g+kQyBK6GhsS8C8EhZXK5I5gZ
sMXPOOGfzQFozuW+jfaxVXylc6CV2EJqM/NJlHuSfw8BvbC83659cgJusaCjkbVx
1eg4V1Aw/T7t//2Zy4/3mT71KSryokZvoNKKSr2EohLKyOepkC0YWu2h0g0p6iGu
8T5Ow32q37JKxF2CaUfZJaGd7OLjHZKmLRk3cYiocrdSOVSNJZ691NDODm7xePrL
CUO+VChVLdlmZizcgqZ5rkvgwdNZi4UbWzF6Fmfp5LAYHC0x5N7DSOeiD9I2oRO9
CAHayH3/ryZ/mkQ2iAo+hg==
`protect END_PROTECTED
