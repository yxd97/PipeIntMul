`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpmqGUBBeR7w78ZsBz0nmP0pScSjJ4FjpGnpwaXP9EN++hraAf15DzgOIRV35k6Q
oX3B2ComJFVdwFqXopKyB+6h/BI3QgITljp97Yp+DSIQtNfzD3wW8ooBxEego0Iz
yzW2NzmJ2ffmSOpY4mAzwpQU9Sh54MqRfVaoHXrHlHatNFXECUdwWM1qeC7B2bdt
pNboz9AOXkMxWSHOFCqYxaDiGxy9nwNQUdKNup/tWKopZKburzlIhxRBFq9HuS4s
azwtHIOJkq/RsBdWUP17iUgpD0n1B47W/ETWSR97w6sC3O3jvYE+W562zdROb5uA
YieouRSD5p4U9t26QMS1mm/vVxBVHbWsqwYem8zTpWE=
`protect END_PROTECTED
