`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fApgvgZrK8KmmnqMriERtrDwzAIS4xV+dsvswnFjMKrCBwNNrCTAuf62dmla6I8e
xBivc0Orp4kX/V4Y7XgF1WePUQCEkyBTHLJ630NoRfjwhpQLa+1DVyYAWqIPCtmu
x2ghj5Nj3Wp/Etjjc6dg16gclYsw3tC1Gaa0iHPu6+f081xAprpR7K3+MA64geGc
UMpeR+rzqaZd4fbYlt21VsbImWwCcds665PODYP9K4aD334sXp7kMWt8nXjMJGp4
wgTeAgCGalEnyvLZF3ItQYknnJz7uc+aIirxA+i+bGJC3mo2MRMVP1UOGVmqZv6f
VS7YfUxXicKVKMLAGSqSD6JuHpn2Ntdwj4KDbvlvx5Wx6/5lJLseFQroN9F6v5By
jSrHwsKF3W4ny9aTVshFyA==
`protect END_PROTECTED
