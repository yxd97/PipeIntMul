`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbBQ5crziEtt0FwSDpUpRs8nAVS6VC71IvST7z9zjyWA/s9aYQltUWcrcsk8axZe
hFzhXgA+tgS1Iqf5V/bqSNTBHoI2KDI6K2RXPSEtiTCCWU086Ko8BoGJGmOOfx5/
ZqPHmGpG6/vZQAODRvo+WcfgETpTTk8HrwTvwObxY/2U/2WnlyiFbCDI1n96An0a
RJ5ZXLJyU93oBoxq5c7/n4NfQLKDDNvKppDJQWb8z12rTLWDMCoyn2xAIY1hHdDy
i2mBKhbL1xBqe97tICnBMFwPhQ8VxehhwtWQ+VzbBD6+PUHbpV3a41B+kKpih/WO
ojYPS4NZRzYXJknEWDjnqecqtzikk9GrLFYrVJyMnLGqV1J0iI+ol1LyjkfATjFO
yHFdjWZSn6Q83nyT6S0J5b5f+9KJZsF2oA0VMXiF/W9jRrejnZtklu/0oBkeBQVU
Sm9Oa2ZXQ1ixiaX6M7fMsplYEWdco15EorEmPz9ls8A2A1YSDQFqXysCV8n7/xBV
`protect END_PROTECTED
