`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eyHRYBqUbkk8DPnF4W+BsslbK+Y81aJy+6LIn547/dJ2TXrL7k3OcRamMM+Fvgh
DZOtGY7kYEjx/gFNzEnqGirHbf4E9IXEyDFYgLzPIVScy8oqy677UkYT/UEQbNNa
jFUD+NxqjpXR2Cp5TNTXNSfILQnCt/tlfXMKggzZlXUBErSjjp6QqMHzcR0nBICq
DUZ13rawYae9daIi7oPyX+iD7R4HthWaU9AYWLO8+aUAY+JaNVi7f6xRSAran08g
eGbidd4cAukHX2nJLJwLr6gy2zb7M/zpnvySvIR0kIJFx5+VIH3YnnuyoOYHoP9E
0PzJhZnRnP08fFVI8V/krx1bgbLSmdHGfudWkNqD8UY6N5BMq1wEBDmcd/8FiUrq
HIHd7YyzA2V1qwHtwMIosy5OjS4M9mZYRnMS87ZcoM72OBR9peux1pa6YbhZtQYj
vOfqPJSoOXjwyRI8dGqcsbysfrFUotFam6J/pZR7Sh6nzELvbo2eYQ8nr9D3ipt4
/tzxlbMhKMoVlS7oQDYa1R0nj3LEn+iIBv6NY1OhxNMT7QsPHPa4GdXWtoBOaEsd
KARVgV33k14GjfsdeCWDvkQanY6zy+KfNFEDn6DlILATJdbdsUkNmaXAXUJ6RlMR
4fuZ8Q1xFhwnKdZvY2kBIt0djLlFLH8JoJ2IZ/7UgugIV1Z9fFw75hQmKwlvtMTh
xtqWDcSurmGWl8IkeW2FejgrFaPcE8uvvI+DXytJt9IRdB5JpaIuzCcE1HVGhZQk
uiJ0VvZ2+hYyYcly0oc9/NFYmrViREtsOEHekIObMnvRx0y4ycAiHYGxsF986nV7
svQ9zHGXoqIY0qmDDPRM2Nzs2m6syksDh+9LHAQHJ+wZ4GAy0tPTlRhrczJs5vLG
/WydFXNR/DFT7DP/ubF36T47lltCb7Ep+O0ryMXi6gR2GUsanm64vxlSyumytXQM
Ujcplz4Fw6XfhNz4fAcCW9XcCuBVB5OFWYIxdT6va/31BsxCm0QnW1HBbn4CjGWk
Af2rHX1mQ+1gIS4WwKBj6rimhG2My6Uav6J7Hev1JB/28OhddGhrxUqGt+91DFu8
M94176rKuPOSRxsq9N4ohPgW2QWEWz7s8yo6PPq/KLvaCuPSI1paPojYtYLlsah1
yvpRF+ziNbIeauDSG7FMT+/Ybvz4TTeIaAtjdB9eabmflci/eF3M8RQdlBTAHUWM
XFtxlsWbkr31kJCTYNTltOOappKqcELv77IOxg9nJBEg6OppuyoaAga1YOjh3GTT
cdX41cAfsuPtrwiWJPpocGIFnlvNx1tNF0vQbhO7AItmZA48QcdcQZ8TWyYxDXU3
Hb7Ydm1qN4/c5iHRxSC+xt4x9M8tOiHtQEOLssBVzLVmxf51hcLESTCuVwH/tO0w
9TSn7/r9DCBMNhlCErrcHg/9iikwg5xpsOmXL67qJ/+OajKLlC1yDBUz1aZJjIoG
2JM4ADzQXwjQkpnkLR+9ZiDMCh04n3vnuiMoysZQHvSvQHdtxOacXt4cV3LXMMc/
jE50yyYTL++VwITvZ/FQxAJxIxj7KRmigm9a6McGm/Gk9N/tyLxvL+w5uU+SUZpg
UDDF+x+vOL8xbPht0eDqWVsUdDDSWjrd4rLPaA8wGJ3P2bTCIlUq0DrtVBQ1e2JV
+0g72YaXT2CFBCdFt8u6VSpFRLBeAVs+KS6d6jCEZRtx6UqYywtFb5FvVTT+hFdi
FLB6I5uMos+9z7e21+Abd7xg04A07cSIy/eAcMMQFQrWI/CWRPTVXfsla8OAnTe2
KMlpuX6CuzHv9vJr2aNr/Zlu9o+H798hBm9w3/lq3kpYi2ygi5w60I7UmIM6MisA
bsomYTAWYWYUco3dZemjiYlDmIyo7kZGmEfWVGdpPmfPmcFhWdSt0Sem0hpfWqbD
YyRyvMs9ajjbmIMS4l5fufE4ucposg/m271s85KHl+OqBidtcQIT21yGdd7yv5xi
`protect END_PROTECTED
