`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fTtQr99Gx5CcHRqxkETnw4vlHIqZPs8ex3Bqloe8fReVIcU+cUm62J4V4SL5l0d
J6ZDBkJvsPMnlj+nh+A7DRhqP04u4LNTtcTCMd+r/bTy8H89Z4BrJA01MrUlK54h
eCMrghFmj5tu24CJ0iy1PqRF11IkTyCTZX3OEytQJkD3hhxu6Eu+Qr2qeLM+ITnc
dj2BXsoDsEjiBHL5BwT5048/cZnZ2KBcYCT3PDjloVuNRlAcfH0xlD4Qr2Xz7Zx2
nd4W6YW79J5a6f2KiiDX9iOcIUrWWS2cD3b2we6WhNbDcgLgHicWrgPY8v3T7i7A
37ixcWFZL5XW4H0WqxeLW4+6ckR/gVe9dl181M5kt/NKY26r0vnBDkPG9xpXLyPA
E8aBl/Tf8Q5m4BhI2YWSKYR7R0GWI/V81wQIh3pmKXFfl4q4nlIjUej4ZBHVNI6S
cz+tb3/dNY6nr8QK8G8gJov0nOllAjEFgbBzCSAScWO1PcT0fuXw+UYDUKqpGU3T
blh4Ri6GNIw3mGcFE9QLQfUJ+Nw1FNA/yz701Y664LCJx4yXXdx7T6Ey0rK2WVAy
5QlTBwLn1OjND+t2lyK+4oKFqGhjlZ2Ix8n0p5qyUWpHffVHIbnZw1kxZdwLtL/h
rsPQNreT3GqAo31MY7XkR4QuihkkdQ/ccChsOQNsIKtEMo4Un5+ui9dVkz4RgV0k
wGIND0IIHOWWSv2XnRFZvr/5p3bw3Mk7zKR0FKEo254ofFe2t1JWB3xzmoI0n1Mt
wzI/CEB522TYyAX8SZV27HyV8Da2+chcZsJR6JRnLM8qsFJTHtrCmcW+BXjzDvZh
dSaY9tSHbybxrTEmX77TyS2gjw7Wz5A6zJux7FCSztlkrfjN3dXyVjxEmFaaguje
CC+h58JHwktUU8LPwG+R6nce8cETPbbA2m8fcr9XneBPKB1vyXAeRrWle6DDXHt1
RvsSPkdzCzWJOdRzsq6lycj6Q80aPZdRFuG7NlkEDJQYuTsnx9n23z/VpYxAsaCM
AAYuAsZiaNrlpsCgHHVx1hyNah5F5nlUJPdWkYfNI2+VUPvHS3j03ESMHbXvq+B3
eg8ACS4ssOm4E0uVsMUFVTkw2w5lRHpxlxP1IVSdjQa5Ax3ArkNn+1FoOxsuHVQ+
uYKFg9GGxLiV+6W3R7XWLO5SKf0CakoJgLtONyVh2DAUHdH4OQ5GMyjEAJdPG6GQ
MG5Yb2oKr8djZ9a/kQ/v9ay6A+nInlL1Q3oRUeTbQDf1oa+dSeB5BzIbmm/zlQTw
3z9RBZHoZWVZELDSYyYXk4HkISz5tHcOYVYcGyBYOxThQdZ92S9JCYrOAW+3MIcR
loQVeGw3u9klT4kd0dtn/kIGZoPYzBmbv9QekG7KlTak/Chy6hW+xqKZkYE0w2JY
UcZu07UxqbYgEIadHny1cA==
`protect END_PROTECTED
