`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
THX/hwFjhU2d460umTovD0hxB6d5ImOTbstNNn79PWWxlPMrfVx+mRkOwruQgdYF
KtYcG8EcrcyuzqsR6t+s3j77nWRatbM2Tr27IhEcscUkhB7utd3fXG6ECbKCvr+A
sHkP5OOyoOpreUzyjlsDCdUkFQEA4nh8ac9areTtrt7ar5BEsT4qUMbjhNp5wTMm
Wsj2UZcHc5U/Huwep/SluLgtsIP4zPoaAnxZpeEuDtc6oxn3Q7C0A0B9BPu9gXP1
IcoT4AepEIu7hALxMVsNQycgGyI80Qrnky+MPcFNOud0XO6fdqyBYJuVt+BBtC3K
YFjAf1SKCjFH2EOCC9wNNK1fl4FMdpIDohyNMV1dwR6ALDA0RWbi0E7wsU9+MD2Z
Nuws2zDb71InBOhGrG+98kGqB63Epxy/oL1HjJaNA8W5kBGfqlUUo8N3ppLb2lOJ
PZF4gToqcky9gWbyRYFlPZnJInbIg0lqzaHiCi2+U/y2E36YR44DSpgjkF0vt8c4
`protect END_PROTECTED
