`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkSVLKOcetY1wAUm8SXSZShujQgqnNMw5ZJOg0AUtpUiSxw4FQtm2rudxqJPpxuX
rv65Y04V8Pj5pf/ipLfFR1yH0JHHwM8NCrXrCW/ug0PUb+MqWJ3XVXlubaM6xXWD
B74LzD3LZL4mjdbRCj39WDbGYvm/dlQx45FbgPvy6qFnfzMmbjEfdoVZ2BZM5iv4
72NGJPVCgH32yJXr06qyPX0qINeDiQeHqkgxvHZBhN0d6g2riODRoGqpX5GStfCB
B+qong7dT3X50X2iAf94c6XWExmzb4QchUzeKQV5K2Cqx6xQ37Q32yvhfm5ZMvxn
ySg6dOnOvfIjOlSDma0aA0qrQ8uptiOyCAnmt3x8z3ZsrIFiKZLLK5HpYeQ/O5HB
fwsuN1D1Q8ec9+AmPAAVUodarX/KP34jXgYUF8q+wS8=
`protect END_PROTECTED
