`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m8BqvbeDi0vfmmZhXfEXgvl0uXnYFLCZND9KS1PLl6zkJB73Q0tvYBXNPewDaR6a
hr5ENpEkyYAm+f/czKbD5Q7oDC/nSeIrNfDOWQcZLt9KXIqVJYDYIs8WfddTFLVA
rJuws468lQBRzAkr5PZRoYXAVL1xS/iJTgYHmFIHrj6+yOzu8C2HGYELNs5voPip
ANkNcV5lHq2v6+K21QRt9fZZokCxofyl/TLqvyanj2qs+BDEKm9lvUQJR8LxEp+Q
PCQSe7+Eh5teuGnOKrAM5oAP+zU68ixYckmh+CykfN7iSXwNo6BAA8I1d9hH7BdS
2gDucbszsFJx86rvC7tk8xgc7PENnsq9uIB/nxlU7oyZhlHgMcEIbFg+543x0P4F
4pNYyGSJrgg5n4KV83zaFL/rMWQQvUchYLy0wIUN8uvrEEfRcDMoedAUmWzzGdIG
pKgWGWmxLnWm31Gjgm5anO/ccMCJ3xCNlgRYM8b4b4oZmWHTTiZCq1Uttf7/hAyf
`protect END_PROTECTED
