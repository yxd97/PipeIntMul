`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8WFOLihLewSsh69j+FpKROhwF6epTxdNCG3Lj+bx7lXY2qycu/V9XGyMYljbNWF/
N9nbXLdu44mGsGNugqgMvPeWVl4gBDMaT56LpJvpB4en41kfQo49aHa0pJWYoc8V
kebMjHk72y1wgAxLmf9V6Ha3T9urmoyNUJykgbG6FDY=
`protect END_PROTECTED
