`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KxWOS6QB2j7ekd1Gen1p4dHYG2z2kkWJTUmoTgIVpRX9OHdv2MyyN7Sr0AXRgs25
DvMdY5DxFRP61YCfUtZT5AdLd8cmr4LQaeEN5d433KapHuOt98/mR3b7uFbRfH6g
J7hoGsKuKGOU/EA8vnMmLcpqRgrUVb7ioBtihF/kwKAwg6mjI9d9GOQUfzrkELVB
Cfaw2DFoytTm9dlK2TVmclmlLuYXGtXkvsyN8AUFa21nRKrzcr1HF4mVMFXIoQEl
ZB2HU+fQjGm/KUuXIBnK4f+C6ljrTQdGaC+mOXXp3adsM8SZlUf46LiNYi6KNy10
9zeMk2mAplOCILwebGQag0k0kswGtB+kVYZJIy/Ua0r32rtdUhs71cCV16PxSkNv
4SCqXdSgBxBPWWaRU5wfhIp4J6TtiqmDAF5z9eYtASAIzghAGbNzZeZRLm8jRUab
kvxhaHihTtTFRy2RrDM55XYZmXly5yuFWloRqY6D8A4r4sOFctnZDBTfUpf880jL
pSC2vqBFigWxlNDkAH7wb1GescoCc3ObUL6hmJnF5SfCh4oJfvk/4ctuZEK3zN5M
iljPNoACgIbJvfVJU82NidiRO6+pFjsI9dq7Xe3khDnOfGY3cYMMUSaO7p3iSNFU
TtJNjz6UKWenJhilk27kG7zOaTETtdU4LW/kS8S/xmZKuUWD3YfMLyFR3gBPCOD6
Lrof4FYsR1u64+S9DJpvdVbsCMMmI5/7DaN17o5+9/elZobvxO+nOnz6Tqs/CG+z
XNc3RNTsdWrKSC+qAUiUJm0rxRjq5Vv9cXMI8PHr/OiVfT6BM7PDrUi+R9Hc71Mp
eRpTNBuT+qj/IKTVo/YOqA==
`protect END_PROTECTED
