`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k28PZKdEwoRnSoeyzo6VqViSGMlbiQjdwYTU0m20qXFafLS6XavpSk398dfL7/Z3
+wCsdsDNa7NxeWe3FzJ/WRrP595CLh+0HM4NwrgM6N4JzevaBAeF+4RAd54ayYEH
5SBBV0iLFB3ulP071hJvOg8sJQJtrocccrzgh4l0M9XN1wdgkk3WlIaezt/SLY59
XuV3w0Zp/QaQroigUq32tJ8xWishdcy2zs2m2Sdyj3eZLEaNzk4oMsMKX8qvo/wP
UVwNQMteGHyTXRYhWvAVog+NjInw66ld7sGNXLo8HAx0KKGefU5yv071byotZFht
VyQ+n2/eXhHwdRCH/cYPr+CAsmVtgILQ4Ut5Oj0+z405b/lLaS79SJYuhST8l6Op
FWq87X4uH54d4+9/l+il/AlFXy7JlROUcvEjHDQHeUvU7ide+w05Ldl8ZgagAH3r
`protect END_PROTECTED
