`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hh+SPA9dup8YhQzetAQ90lPbDwVMD17cSiw4/HR3/FRWp4mOjl2rpcDrX+gvwoII
ffPsz6T8iuuibjo9lRUSo5eBCEFCkPt8tfTOvka93FTmQaczZzMYQ1UZChq+qewV
fbsNtS3x4c9QDROAud+eHKMTAq8dYT1kyZKwADqO9Iuqjl9ahIGt+Ghh/77zsaP0
/rEwPV9j7MxBp5PtKtsTOyEgNf0BeExIwO6BCakiFkjB22Wc3mvIFJvqKRSEkihT
FXDi3b1PBI1sM7prM82flvOOA+4HkED2BdO37G0WewNd64HH2nkr4/kM1xBF+huK
45B+nICkAWozDjLgCJlRGPoM99UWgxKaX5O0EQp0hYuYwSiu/hN9baJfxY7xXzpE
jsu3Ma7AtTZ+DD2Kvcf8xnWdOfOPfHP6DplNLZObnfzU0Q7TFg4JHdxT3Kcm1NAQ
9LDmy2V+qCqMztYoDL5bvO103U1/5i39PG0oazAeyuOpJ1IMLZddUiP41ycZlhIk
WMa7cyjaMdyX0N25FGG6g7K1BzWpbLA7zadMiIuK0IQ=
`protect END_PROTECTED
