`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8quStoC2YN336GXxx5ab0kZYlBgdGL7ZWgWvCN7g/82/Go2atHJLd8GoMfoSrs6b
bxYWppzYBtdXVsIoF/KdQOmpXwg9lrmmzcfnWC1doOB2WWqh4w/XLwECxuPdqBti
+mFgZ0YhU7bl5akuz1Df2tGrYWwKck9CIJP0kh1/hCWAKJv1jpY0Yk0/F7Kjr7PQ
7Oiznt41AcLZrjf3kwFBdFQtsMryGncsP3sfDrV3txujpCdV3QKztaHODRdE0q45
UEZXRic8zro9BglOwDxGQSoP5YKR1Ra24UuVO8UqvjJVgfOAxFk0E3GZ9IouCjuY
ZB+J2d1oFrGtAmCZzSBSe9yVKPmk/PVIWti7pXlwBo4=
`protect END_PROTECTED
