`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Gb99nggrVo9ixvTA2W9bBtAJLhQiCyZau/+5/KvjezvZgp5+Zm5w6cdpng9LgUS
K3er39Rhn15j7/QWRmjSanIocRxzJR7DN6n9PWq1BOBE5CA7iit11aWCuT9Db/vO
sQIPIOnlE01Jf/1Zee5z4laEYTBvKFjVvtNLR3LcWy3YGZX6cH/OuwWWnCz6MeO/
nC3+LqgE2ffZOcBrGCyYDtQCzj8VZTQIefKYf3oaIMn6nQkd2tCTaVD6o9fDRmiU
N2sn/y/wfIajESpn87pzJkBA7McyMMTbnQ0sYQMCy6Ngui5ysoNibQaEoVNiKjnM
2BGKP6Umy7VCaAuNcNTQWFVMoEn0unE0V1FjjquufbwUGfOocgN91hP5RjwcGsca
r2RRAaDCgucjcXUwOEThCymZvv7kxB5geB0aiNERDO8bT0rmb0bwz7auYTT36J+n
hgEg6tTnrM+DW+46XVoeK1TbJmEEGC/T/ZWjILlNUTUpNPY0jqqfmbxJcFRhTmVR
6L80b+iM3jyzwlYxt7IkOFjv/pyFX8qUvDk9jXSIMcpWaYFPzEi7H44k8zaNuera
5xgWl6+d+3Ad7kSWy7Kyn42pKsjGQCiWDvMWSnlz6PgZaWFn3nZXqbnErcz8FgIz
6LQ94xYmC3pFf00q6ypaOuzm3ayBWDJM7R09C5C0gJnlS1RNVThM563nI/RYivnU
1HVUE0Cl1zkHbohN6luxPZ5eUuNp9zQFp58cjf8d3VZHVH6iAyUMWMeqkC7P7nEx
Ziu0UQ0wtzAksJH/YxLqViNqF3Qd1k21qSxlseVESJDv+NB0/jAHM972DVmtrkZ4
76yJwiGbwu9Wd1+mgSY3Aq3XRGmeiRQaC55+/YoUzIYBEvoPsY7AqTcpX4ZZJCks
t8q+uTWV89ZpTo3QGxyUY9imkxw+H/c39fEiCmOf8oR1dPIqf/tODUMvwaMdMi5t
BW0YUzf2VO6ONdbnEabW4/ajglpZ9BtVXVROlCqKxqgNE/kIi0nEpxAGB2Q2BKrT
uM8OBbTarpaSGHVFAGg/TDOgcnycEs9N3K5jxvhujc+6kQSmtl/Edl0GJQikoInk
pm/6KFcOLu5pIOrlFPQduLraDCAiIasVDaxa5osnE0boOYHDjRBSJRHGB0JOBGG1
m6WGumHvSI5XTjKOQ9Bj5HAUdZJUWJpLtvbpleHajH+FyYARZolaiYeg3GftYDZE
J7ZKiU3TMgRipjOR+DyW0+3PPceaW5dMZkAtwU9b0QESXFrmzEyL56uFxKEVv4/E
k6ygQVk/+4w9Wadsh3xcpjdEUzqF+Mi5+2/+cS2SO0XQkLV3DfINMVjE3tbSfMxg
/IQ9crcxEcJKuZVdDHDGng==
`protect END_PROTECTED
