`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6AxC4GxP3oYygqRP9NkfXaIEbTI4sB/EHU/NYXGjWFuPhnWCFLyMy/X+kWbNYdOk
qkM+Q458DaH2gHRvdNbFP+Ny1HhMOGQFvqOTjiGeuWuaVJFnqMWyqo7Ita1VixDT
UY1457jHJYv7ippdapGwhlSIEX5KdpG9D53VFBFZPd9zF2QZUyTBorabuCL429cq
DfiYfWy0xtJ659gk+c6S3z+tHcdMZ3kHv+LE9AS9YZLs5fycpJYC3uJA1r2Oq83g
Qz/anVTi5xTt2byQ/muBHBeRqp6bVzM2KfTd+rcQGrslh88ZUb1HWFJnHpPn7eQQ
OnRhofW4zx61k84Bkc3J0Jxx/vqWaEIUC80xtjDj/sKKVk9o88m5dp4UnJoXghCL
7QRmSFtKY4aLw7aG3GP6GqoqBBMVTp4PnBtyi3dmLuHZ0+PXVj30ZyLaVKmylKvS
EoQmVHndYIoth3TTMJPapRkDg8edqydV8653t+x29VJvsHVrrUS5GIBKb7XKQu7W
tg0OkHuGxex2727HsSPtzWBo47IoFn/HN9/bs5DC4P2vaoW/Th+93ebp0UbXmD1D
ht3f6ZG9tJ1g/rCrbwoGuQ==
`protect END_PROTECTED
