`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63/IhaiLszWM9jCrnJ6FHUCkTHKdbYwVeixyRWe4JBLxYBafXzVtWF9gwBKbzlfQ
2vqYdpELsz9oGtMdyYIFtkJeBaRSs1YVzk6I+IAzUdpAHb8WTkg+zbhs28qQCODi
/9BzJCSnxEd+q+ga15dwTUw/gaYrQfteAGEXUFoQqgUD0A6DdrGFZI4AHP6tc6w2
a/7u525EAAGUE0XnoqRMMfpC7S0+ZzYx7aVNc9cEz8zRcpundv/aO6FnOstWmmtF
YkCMbzWlBBQ9FnaDiP5kbolHNY3JV1640qqOsD1zjEr7Z5PpSQnjsD1QbaAYknOW
0TQ1JKyKu5rthXUqdxxGL+r8QqOuaRIBD+wyDCXdFaHa/iMW+7jBV7ZI8kOKI1Js
IsFBraIIw+xc/FkmnXL7JQlZ9BC2gdXy53dx6Zz1LzfZMgiaSAYWn9BwUDgq3axk
rIcrMJ7tJ2BqtpRX9aWL1z0Zafyb08J3qHJLQhJlfx9o1Nh4Pq3FSVFCWjld+O2I
xJKQsHM/IIpOqsftYu+PTxvbUUnzeNF9mBE8LUfrOfOK/WH2wppsJ5CRjS1DUBK9
p/qzg8ShhV5Tld7O6KY4jM66TRHA72blRDJtIxWCPb8zUVdkG/bRz0TED7mfHcRM
5yPWcwgM2OnoXOGfKb+sxAR6nDH9/aYctSoP0Rll5QCgIdJYsAzl8iuHFEn/MExk
i8+sfEsGCCatRf+MyKYN1jY6EYcVuys2at2PBHSso80R7xZ6//onCJevkpPqETZ9
gHi7MaFw4ch5KkVYPkRxie20OCW8GLDkvXvpyiA8eDiHKssxUVGUCtWhWfPlcrfS
r4xfXH9d/bqkAEq5T+giMOE2E6N8VtczwmrJ4lKsKa4ZAbRFevlG6Wb8ap4PJewr
xgSKXURETnJv6AZg/nFlZqbpgMl07ZCjr5oLxMTn+jSUnhSB+SA0UMCVYBy2krNB
`protect END_PROTECTED
