`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jrcTYeD/4wgcjv1aJ6R7ZoQhXD89D3he+fkxqXhqZKuMdV3H90E/4eSMDt/4PWwt
15Zi6JAPDgHXg9ljwyM+t0l6rImkibfiLMaSSQO9IVvHXjkx5k1EsSB+IzxBAYYr
Ix9PJnoSdkuZvAEWuIQCBLC7XA1h+oNd4n8ZpaF+S/wvCHjk0i+k7WTp4KOpSD2X
8GF5NPFDt2uHy7X5CPjF7FVhMiFrh8/DFjw6r1EIp8NJJdDYdOne85i7TqX6ahFz
8U+QYF0hBzYb7G2uRxn817V+X/zeRsz3SppRr+s8Tk1hcjbPPk1B/t3vN9n20mus
AXlZvliQlrmGnn5c01OVGCA1ciKd1fApu7LS8HMjLlF3iBI5T5Ggr/VQ58El6fhM
eVxgjEhJPGnMUxBG7Of/kZyf9jkYtrBpLpyWrzgG9Rk=
`protect END_PROTECTED
