`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMvSIRlZsYjszkKnewFTeR1UCBthM8hvrLDAhcVzvxReuc0f7Eb9hGs3fahtZeOp
6sk4ta2GmpkYzvqSdUOrDp145TVmuT+AMo4R8YNHShWQEXWR4y5l7fbrpxrXeyy+
UZbyULEeRqXMO9g5JhljulfX6Qfnq+2SATBL/2f7twULoUu8RMVUp84928/s1Xwk
guigF2ZethdT6PLN9td1cNPobDFOrh0KX0Y7wlXFVoovT5szkBFEYISCAEaWV93A
I9NSchyi2dc4bFS0X0XbtReYxc+61sFoId4MvL/18+cByZCHiZdhlU3jtVcRULrt
MdL/6PW72ZvNVbJdVBYq68Xx2EuTYkd3pQnL1ERfA1OuF+0jPSkdb//W5RMYu8Dh
CvmCZ2UvPESnObJlZUagxcZAnVVEnaA3DBy24446mHcymBXpXRldz0HrhHEnM3uB
cIXWymHbB8TMXEFwm6OZ/qWZDFIl0lFNqa+IiLoYvQlkWRM0CBwJshmqv1oTAceS
Nl1p37wTD1HPsvbA6r5SNaNMUlqpv2eNPcUNHRZUihE23PgHYX00Ej9WbnGxi95K
vgSZ9Ccjnltn1mqKAOxfTlLflrToNRoSyajzB6LcoI4t2UYRugsC9bMQxzA23brW
kX7AZtrnE5ghyNBn3bBDIcpnuWWZExZEM7DS+3PC+BPzdy59ELkC+/RfDb5NOie1
vc8k3nvzSAaY9x2pNrp4O6IsOoGEgJsISiT9M0oX6HbXyyyX61oV54A6TuFLg3pZ
x4ycqBf2VdXRdznynDXd8YUDKFi7a7Tdf82yCF7QJE5vt8N6cfzQeU/F+avKals3
XJ/foTSHdGJDJkmQ/vqZM6h4KNrecL8kFJgs2vUL6Onutesg4LXGwI2FcyujWQ3u
pmDUgPc6g2hd9e1F9mA0GQ==
`protect END_PROTECTED
