`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jzhPj7jdLhxHFq/5urpPWbft6apcmq1BYIRvq9OnalDEzTjdQz4jbydFzWoIji3+
5a3hkF3bbTvxy2NyYi25I1s+mRK0kJVGVC76nNXNNAV0NZP9W60AW5jk/xFjboTq
7jmyuLJEA6rbMUCFGiCFDsFJaEqtDYVUfqZ6dE9hIu6PuK6XG9e4Kv4iI3hbAuNU
1CMxuRKFhHwgkZ255QHJd9751k5mm2pG9AuXI5cq71o6w633oWagT0uss6xYgzi/
AVEXA5aldzYjJ/MeAbM5ndWSPL2fdA3YZMmI4isvwpMTzkowd4wGxbeuvKIBSIu6
cmZPwpKRazM/XzS90OUc1SU3WCdNAKcac1ifTgJmRzh6+SgZCfVwej0SuCQEItRj
FBvO2JhDx2vMAtQxEvBOo2vaoj7iyeqyGFcSGvvFNV4=
`protect END_PROTECTED
