`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTatRATC2cwDQHBXYK+4NuxBktVJePPjdU4YtXViJLl9SsRnA6rQHGefqBethBRn
B7w0Z1xW7aZvPUej1mVLlW57551iFnlVjBnjkZAxBdeKazA3JdUYLSlWobdQx0c/
kDewuqGnPEj9oYq6eyAk23JXcNNe0jfrwBY8jkNPQukfjV2o/VbJdEfozNZBhTYb
KGteeI74INvE6TdigE66AZBsP+tHekO0Onqo+TJ1sf16UMCuwACQLg/9f0cEOFZu
MhkwL3TDckkG533C4u2beRuCkB47AgRT3AofYWcCo5RxOhobksZVYkFjz8tDQP6W
5lnxcIGY0JdXmHxdbWiP6Q==
`protect END_PROTECTED
