`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52BytDjDRiFFVMVx4SeseeeXY71t9KNKdJ+riXUuB38aHrMTKrTPZakZyOH6ejyJ
8TC3qJrq+435+L2A8g76j+Jqdm5lBnYmFgcRdkYsUTnoSsWcvVxyQxUkTR24pxbW
qJgmGo/wZdvstxhV/m8dHXo9AoZ9xKNoakd3T9xgXV1UBu5EtHEuFYa/Di/3QfJh
vh+18U2ZpjAfhFgh9+uCjeR/nAIm38TrQBWUuu6vaiLd2oEgeGjDB3sgy5lz0Aka
lISsCfJcdZ+iB+PDZtaJF7IUg8TWPqn1g8ksXBW9DRdLsANq5hPCrsRwKVhTiBBx
wp+KyIhcT/m0XYQQ/Lp06w==
`protect END_PROTECTED
