`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MP7UFeC44d9SivspWnwsNKtR1Jdbc/gjmNlPhWJBVvOTpKEKlFx02pTo0PHIPacZ
xSx5qEkC6k7g3exVk8Zg4IqM65roqSJ6YIKju2hGaDCYCuoQGeHYUoKQeu4VVPRb
rNNMEHa3baWqnt9ncPKDIK6b4WZjn0aB9BtN3J8Ou22GoREi3NHraBzHrZYs27a9
iSdKctV1GE/tKdUXnquNXRgqeJUC8s5PM3v8h620j3iEYY47NLdaNg/KQa+Lannn
BWqhLksRv+eH6H+wt/OXDsYfsUw2KcYns7M4zknHDdhg+zbhvFodPEMNJHlL3yqt
RGUuvzjm44MU/NQ4nICGBoPcRn3Oi+CWHkMI7Nlb92Ju38dqGbPkGSz/C4pAYKVT
uomRf4Abwtys4+K7w9szKD6yxlKOvAFjYbhTltDdYlI/OJV+tQ587dIX8QcgJzCJ
zNQagv1mZpJOXNViMCEfV+VhRaaH1I196cHqqRsB7v4wcMMqsQLvu9DUsnXvGaWK
vbbRJWcLuIBqqtYSPypNOA==
`protect END_PROTECTED
