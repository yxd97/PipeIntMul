`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGGm+gNoeVbiZMuOlHuHM4H6iayalwTtEt2qMU+Pcmk8jrW5+oZ4OTwPDaZueyNr
DUQtipWbf/Xtj9yHUZw/NRDk/ZMyl4ySF9f8/JO2ycg02mPmpda3k/48OyVDJu5D
TCkLRC3YTUN35A8INWgf9PvslBN7ev0W6KTJkxwJL83KZSNgeG8ECqOmEC03EYyz
R4DlMazJVvgLc/54aUC/4okhZGAP1fssydJSAk5PIy/Ieiu6CLYOChV1CX8JtRrY
vSQXjkoKpv1Mu84X2JuC5k3OVAAJcC3bG6I20kYoJxjUmLF29XG2rl+Q0jX50IFZ
tkY7GZuFeDq1A6uwbAeepsytTYWFODxiIwpcuYlKeW5L0lcDdpeGVIy26f65zP6P
7AGOLXOR/B0PehpmT37lG+Et+NlZDtojakAq+Qo6OVipaqk6lEYLnYlGbgx1W0hL
GQXce1plvQku6gW7qcIATA9SYEBlC6brfq7j3dspXIx2zhC24dvO/8HoHDUmr9Zx
+/+b8CAb9yJuZFJmp28dnweNy6JiPMWfn7Ss86Sf09Epq1G962qND3D+Bx7+hav0
gdquIIGTbktpV/t4/1QZx9r/oYCVFQlyM5uKXbPmX2Czu1ECyL7PhWk7sV9FEX/S
UeBWylEeqWFc+/o2wVD33mNMg16C9vDYfGj6FOl3e4BlevpNczJ9PZRAy4iNjJPE
+Wyu18k9JNE91S/VwMZOPFv5Fe6/0kq/Csuri0cmk0x6bZgEVPYfso2f4UytQYgG
OIPu/AO1zfOB2oDZ5xyoFUdofQtY4uO/JgKAtikiud2qLLjmluLF6PospXd4YtZF
mG7Ymw9Fw1qSj9NrptHPnH9Jd3kKoc5Xld8wP2JYcqXDZWzeWSQCK0dbDxvl/U9j
0eAvWPrkkAou0dTknVCKbvcxn389XaKJKQFkphOknq8w5BgyEDu62DR+jjbCfzi4
giFGNa0sUIHY3GhWhpjgAP5S4S2PPbcTWaPXcwtiuv/voDWpXAwKNv4tCMpkuVIG
HuWrg5FIf68SfqG+xROmMJF0erGkZPl4nkgl4Y6cUoa4WubN5jc0DhGzgeyoJB1I
YBCG9Gw0yNv2NgD3kWmHs+MOMXHEcjF9ycht2dlBF0s0bqNqk8+SK8ohhk3xCAn8
YJweyu/0f/CnbWNdIJjT2CBDaKepbn7FSwTwCK0MwEfEkhvsdRtaYbt9gb3C4Nxr
gvGT31AQKAUR8jXQXTTvqWubsY9y2GTbQkF2toV4DeHhz4RJ2amqmbBhomGFEQWC
q/Fmq2t5NU/2p6YEPEyRkYgA44GkFpBPMARluhnjWh+IvllT5IxUMCao7yrYdRBH
OHfybUQCzuuvINK67/lVGvOBmjsMlUEhYm59D8KvQgalCX8PsnRIzSgMJ+YqA7Ei
MQbSTXl0PnyKzjrqvmkOUxUNZu7lJmQ6ZH3ZN3izyXJmoeCkUvZRDgxfeM2LQco2
lr70vJ27cmBolfyuKOfeNs+1I1JyV8w8UanZ4MhAIrp7rw2YGG53v4YejPtyV+ak
YCd88IF0xG3GJwPrl88B6fGtqgNtA7vN7Aex9MhZqDf5Sy5vzlE38FgLZs+c4Qgm
MA6b194yI3cxtnFLDXINepkrwuHrsXO+oV9RVVOlWxA4EsXKsPFwpNPcdXNsV70u
P8Cyn904eeA4qoLsvih/NLvgiaU23DwxOqxeP7WeIvCSTGPCpVJjCY56gulJu2uY
6mL60Ao1fUTWwc16Eb8TgekI/sGZNU94ekGdXxo/8VaKAN3m1nJQ6JC2iZDmRHGd
RkNzXAyrZr9vOn+XelaWUhPkLWy5iRYEfI30DtncMKccJiRbHVN8V5KwpozZbPYU
3mb6cvx8jVktYG6voPhAE6JlsDsY75IO5lYICRqD43sYitKj+BXnvW5bc9vgRZQf
PaU2ObZY3C67XW5OGYhVhALoUrXLm+3b/UmIspqchBr9qsksLy0TlgfbFH5Dyk2w
sZUvbb8xIBaYKkP+Yk+GBj6NtQ5JH+Y6h7k9VxMgbMAwyZn/6nRMP131yxC1wAGr
bZyOfkCWyMqfiBfVeP8LeUYKcnckUF5d0Fui4CmusCci3t+yxuEd/eATTy/EdACi
O3mIG/DvowkTeeli4h9Rfw==
`protect END_PROTECTED
