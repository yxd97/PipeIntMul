`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fu7H9VlyLJL9l6reHk7iHc3ge8ke8SOIw6Dn1uaJstltOLSTBiL3DwHu0BrtsiZj
i8K2RRzZHrdvselNE8eKATxMxnWj3VssC2BCUD3z7sqZeym/fpehg/bNlJn+GUkl
vAyHuoWDT5dOXR84Vf+UBJXJBJ7dlfMZwiG8nlyytjGeRpJPXWbxwyzfRln6xLx9
9Fp9FOedabcc6sBJTnUXSEswtWpjaofQstD5jBNr/nB5mFcZzp8IzByGuXGjzk3W
sNGpHGCizS22zcroHmI6W+K8xMHgnC/BXVVBzU7l4lwTvPgJySnXdmqrz2Yy18r3
4cALlvqGYI2/M3NEQkysztqwdP5d/G2xFvGHBTLeIHiomiTzmXDBIKZCTgCgLXl+
af9KNdmJ19acrwQExSLd4r84y6cYk/yWoeXdCjdDaggFbXh3tJsu8kEeyRsIXx22
K2s6qbkBTBt9GlDQzLYse07PrR7fqETdB/dNMg4rrkDnMz3JRiuuYbUs44xFyK5D
sZgcMYlz5iyRnCYFtPIb1RwZf4nI2EsR49l2xy4IcjMzzqg7YbSUt7Xrsl4pXYWQ
dKlaUd/zsgmasmuc0BmQSg==
`protect END_PROTECTED
