`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
62sSidaJqx59FFcYboDi4lQ/PlrYbg8iCe7bCgL8oqLzuGRbzTge9w2ga311PnZJ
Nr7xXiT3stG+os5Ol9rtAhnZqkWXrfcsCf1DbLPiP90DhZ7eniBXhKH47TnBF1RH
aGRF+cANhWVQY2o2L4fmxrfLUdYPHIYtyivIcqxvr9+NTEgDlBSkbQY45FPQq68J
qgrbF48Y+eGp89IXnGuae1ZNlDAyuabcc0ABgs8Oz9QXSrhQx1gNaRlw1cPbQafV
X6wNv5qwjZC6F024NDNAWyyRg7eFNNk/qQuyZhrzS+oSkLgJ2aGnzZhtnAVe7+8g
IMydm5Yu7AnHCjKzmdeVQqlToBrTV3uQoIfvaxtKqh4ccO8j37zTx4VFrX/eXAYv
FEWTpGANGpDFpYpdhby5zw==
`protect END_PROTECTED
