`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AhP/IETmzP5Bs7gWYlbcYvEzu79w+KjTfnXS29ZZRYNDQRYucibVKJCGBlfOzGHW
8JWc2fZbrIcGv6achrxb2SwQJcl/rXcAjuwBIRil2tTv9smaXNTeqlCJ5ByP1fi+
WwjDhpAtl/FL33dq4sQ2smIF0PJm5eLsuE12ivKfSWQ1t/RM8AxmQl/Tmw8XGPkU
5LgQYh1M4kvitSahHO+gzs21RqSzTwXyRilHPqxKPTTX5W5BeHh73Ovv1WxZOCz3
ADphH60TlOkviUHE8tNa+/yCQytrCOTWN3Kw/Q0lC6QH/KOQBvU5P+XozVhZB7ni
Un/LR3lEjOFdlXwAnC9nSKEpeJ/MsrGTibkuScsW1Hd8RCUNxMzEIwlBd2emmQLa
ItUAfWluwakE7qjvfFw7jnM+wstuWqw8mMiFLAvhHVUj2fVwDwWsRYlJ6Ztl0tKv
JQGI7EACGujvNfoYvGv2HnPs4WHeI+acFzazN+GtaaMXNbMRUsmmi67khvkWTFbp
8T1TF2EY5j+Rk4fqFZ73sVCcruJn5FFVAcIDKnt8AWkoV/ZxrNC+XFMwszW/ZoQt
/fLTyf4AS6jIoZz1vwGx/w==
`protect END_PROTECTED
