`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fnKaeENUJkhtHMT2EVrSAAQyp/OHWgpcW3Y+E5DQ3JOG9n8HrkgeFusW0qFP09jV
gMzpTCkfAr4Jf59Qx18YlAWgWzRHAScXKW33fNu/NywDfZYr8xt3/3LwB0BmgeGe
RNh9sxEcfTugfmp8bFYzEr0Umw6nMLvxv8fKWOG4mxAvsbHxQWkYI+jHfOn2pcpR
DztSWgRwDv7YqT5jQ0MttHKb4/DlifumkfvX6wWAeghNvxRdlkedFXN3YmLVxQmF
BED8lFCFHuOBuBmnjW0CwUOrxXlh3hgfbHKmz8IbKZuVtA6KQNZHu61UbQXpaCk8
C1b57i0IVAhQyFUyb6Kl76j5D1kzBxGpZsOq8ruZkRj9es6WeparPxzzzikIUll3
LZuMPQqmUovxr3UNPxYH5iwmXl+B+eSHFJAQhuSSCwI/5W+PKn8I3XijAcC5FN5k
VLi4hd2Wt5GOTveRXYGXLTTr4v519OEoRMjGj43upLwNEODX7se3wVVsDwdIWuA7
0eW0r3nT0dZorhUjN4Cqj6uUNI3QKkxJiVM4UbchASrPJ6IrdqvpiKVO6izwjs5/
DVZgrhxe/aUoyjGdMpuDekQU3kyq0l3b4q8Kp7H4Gls=
`protect END_PROTECTED
