`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HXDBwv7LutoQdk53+Z6ETaA+1EI1UOg9GuOsCPzNLPcWJuVrUWyIMnAKsi0u2noo
KFv5Hr2MYbPzR4kehwUb3itpHZrVn4VwDyjhnt2A5a9VXoGIEfKeeqrpa+TE7S6/
dpQxNcag8vzj2+wj7nbSiGC7MgfSPaOzRD7wkomVrcvnNyoesDfvW5D/RiVZerdw
dtWnTJZmvbHEU551vOeYYfl/mteUdgtXi+CzoB2pW9sAzsU6BX8vPB7XfCxj+dLn
CcD9hweXUxGSpVkOH0OrYPz3VktuoVDsifritwvXh6Kn7oXNMydSx6yYJuZJRWO5
siWxpJEAVFp3pHXS/tskIX95KSkOAoiOsj1yXVRBVns7GDsfNfv3kdZf/7NJyyNv
pCNNMfs3EM/Keu8uLU6Z/ahtdZer14lTuDoHRa2cnlWcGHEyKyjmEJ2qblL60Alw
lyZppAx2CgzZYP/Bj3ieKurpusTtrQid4Pvw1Z5lDkURsSw6vb1dIsNqKlLKfVTR
kizDmlzWSULQz66Auluhq4BWoURB5YDyCbhJSTHrt/y+KovwZfjTIE5qivro7dNZ
mVCEHyk23M/2KQXRe2VoltCZX+QXMlNm3yxXvCZ8Ps7hP7zDlXyUjOa823YhYpdR
QZ35wM5eiK5/zLEZqri+IPmX6TWqWa4piJA1jPEaqrKbK7CWnZVKTqI8JtmlPi+C
`protect END_PROTECTED
