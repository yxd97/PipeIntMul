`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Zq8C89YHvl1dj+m+lJq81rwveDL1L1FILndTheOnjrRDTS2Xd9NLFMVcehjojNu
ZtJAaDxodGKxZJRHNU3F1n1+TwLrlQFTTnBvzMyuZjeu9s6wIFJzjBoYMZVaAkZm
lUpcWtTBSB8E+xugiqgxsdhPyA7m3yPRCWUN//EvhOMMUB3OGfhSbiYAvrguUYvs
6lE+wXC3bbnMQRjR9UFdVed24TUSZjHy6oL6TtO2ViiYD27CnXeDKdBsk4flPuvF
n0gAzMWdtBOxweMy2gR+atAzlNXuu0Up85Au6ywC/DQq83WwvU9Xmo4sHml3WeKi
QhzbcNLVQNhx+RgK0RpchxNAfXmiYU0bpDt4O7jxtVa6mmnsjoCTEczR6XioqHcB
7sdp+vmdv1R9FTg2PK3Y7zeFANFhq2/AiFBnjU9/eigBIEqNRaPSjsnHKGFC5sR+
XtRhtePtlJ/+I4ZgzjEL7tAL7rdk11ks4F0VV4jAIaG4cNeVoYVdOb1ot3q2pbpu
CNX1OniCNLMKT51DmvLa0wUQOjo2UmWA7tNNqd7npu7gZlfG3KatXQkeDXn4rY3Z
NqwJaxT7dgEl/ond2lY6R7T5qyAbjIWYGzJN5WgH1/AetA3FdeluN47O0KKEFDeT
N6ZIrkToNbrWQaehH9m5kXP4WGYBtFbaQl/amq383hjN1CufCGEUL7NvKC2xbQCq
vvxc20+pJFY73srsaWrl5VCit8KebTWUGyA7uT6h74mjo37RrTf+7FbLMODDeia6
fWuNLtuFLVEVFerEd0agwPcv1jZjHiYZ0n8QbLP74EJx9CSUf2EhzqlwlyKlHHlM
xnbMou1K/AzoHtY29ZJaw7NAOyFcG/PcjyUVmTiu1zIe5dvFzCT6swhc8KRQ1XjG
r6EeUJ3p8cKfxFXwqZwhAaO4yJmMR4nSZTOCyVpqTLqd7i2glcW1nZWcl5nPbVFS
p906Dfw32R8kQqAF2LvCwlhKaoYO3Gy5RqEvH0DpyqBhuR8vtU3PAFW1zdONqu4K
HNUbEjKBvnsMZFGptRiShjtERw1m21CSNcwUkJe0rhnMG2fH5PTzzxMhtgXDICRz
M4zuRjhdRduouCqzyvhrIYrlmVlokVOjREtqfAJKI4tkp15QJFgSUmq5lFqEAKIU
zXrjZnKrPigwKscr6068yUgxPGl2o9k2GwJgR6v5QfjQWuZcwKjpFzgk3emcMbLF
4yttfS+FpN1nn+1xk2eaYvwxQLB7Di6Z6qX6s7Ee7WcX7uznaSP4H4QqcnP7MY0K
WCnn1YY2Z5q0e1DT99NswwZwr6zShyTUnZYu3wnCWfN7+rpUtZAHw4CUP3UOK4eS
XlPiTfhmZDRUFl+/XiMVw5rrU83yQSbffw8yOzvJb4n4aDYO/mBYcRKjPkAmZS0M
iLYsnzTDaq5Wf1IM+O8Pwk+duty0ml2oRdKWPbPDAUAgmxKBbLJ/F7b8OzonZBlj
39G0A0T0z/LUgU++xOIEvBp+EPvmYV23PvM2oMg97nNkkFjY0GtOnXHv1rA555RS
MpvADw+2MFJtTLM/YCHQ+rvcUGNzdJogyqttMxUUCGCaMfqsDWCpKoFN334Qrwz1
usEY3735Ys7lO4MsDcIjai86XITVgUIJ3PgqzsV3F3BuHdDM2HNZZKH1aUq9a1co
eaCrryFJob6MHvyIrRhCK6PcxJlHzSNwpxdS0DkUIk/peVd7DDIvEeCAIVeQa+Et
B34j85bLtyMbFFPPOmGTj9Yp4UQ/KC6pix490h9Z+IBb6W8ImrRARFbPL5rVxkP0
yDyrI07GM+5hiFUrHkb3tJ3nhOIalofgAl5SGZ4Mv40upmeHAWvyWfwYXmwhY9OX
wkYtTkfTk2wDRM7sOKae7l5Vr35QLqlWpDweui2/Xn/dSq+d5y1eYg7WU5e6wMTC
dYzssXyuEt1ULJtQRz0Xzfk5zz6GrPX4m9qWgKNaM8WxMuV7caKSnXSl9GzWYgEk
+NbfvQ8t3FTrydZAH2+GRQe4w5CNkFpO8MaLZTPwzgXC/Obm9XYPEnsy/wcxHXyn
TQ1wdjTDTv54+4t6GHHbwsWLuqSklD2UJq9zF/Q4X3z2ru7jNndu3k9waALP2MOK
HETKxoTxP1dGpOXt8pbKUFW7+AkFlRAsVT9y7gDNXqA3vhkx2JoymwjuQDLG9pn7
NkjtfnSkS61mtMTAscWpSayA1r3etGW1O/82puOhw+Gsop60PZfakVfRgHw202+I
dlUPKLY4NT+YpfzynUN84QHKt2xe5ZtKgXKnRn4R7hJrSGKnQPFA8NxuOU11owU0
lo/1vcdyfis4rcru7hilRmoUAyjfM20J7IzxVTRCjtLz/ZtMRWqHUkdXBIaaN4dy
vSXhegEIj6hkHXKC/ytW9GPcoAdKUXWrbf8N5Xp0WvmJIq0FfG8BFjR00FTZVO3+
bYZyyq/9frXCPHQkqASXmMhuju3ICx1PygnlDXRNtoqnc9N0R/yhA3V85M8q8g6r
VQDg9bZtpfMepnRl1r9je08kV/NcO9e2GbnIf1L1jnvVrJfWVHzEY/GljQNoL77b
J/FgSWj+z3TTYAZZoZTFc7jYunL5RMtFP2pyYbfOaOCLVzjFwsCMryWU9c2PkW2a
Sfjc6OOX0gIrrMfxppliVyEg7Gmy9oemS0LQryBAqct2MFWlKBCR6sYebVbD7hhv
WTUuWctvI4TlOoJ1Nz0cYXL/INWH7HmJ0HasnzJPGu1wmjZlj2nupOy9PXy6DCSN
rSobJIH+0CBMTbMc+0hmhdL4OsbZ+DW7X4hhov3B5gHZjqMaZYpX2TNugYt93krr
ac0SqroUC08W1U6LSQlJxdcjvrtj/xvC2+3lTZquaVZ31LgW4oE5O54q+zbedrtH
/ijvkOBah6RFlydXjCN5NtI5ehyfzmLMO8Ivh8ddJM9wvJ3Yhbts6myUiJ0mMSIC
fOtrwgTI7dhHspMjp/Klf0P3+EqYCnJisL3Wfla2dAZSkMpyTM1lzjzyrzM0gfzV
RA2tdHt/MUdru21DrC5p5JtwZHCe7gcySADbBpGK5UDkcUEBmlFolEeEW/UKxxow
7fD9SUxt4y92yZCDl+aeyNSNbpdkmWn7b6wVtXHzHA/Fy/Diu5Ft9NuDg524b7cZ
oc/SXeZwdU7MPbtqI4VxWXDL+y+ZNEOGf9450I1n5ZJAX801S77P1X8p5nzEoC8P
IiwT6tg3hPeSlwLwnr097PjWJ7kYTjBUXNErcNvNpx4Z6qse5+hCO6Wj3T68eGjM
2K0y3gjzLdJTltir7hlX80Rli6b2rSgVpuBEOV1CHsR5okc4LMLzDTG5L+Z4E88P
RbhW1mVtvu6meVhuxRRSi4R23Fa6TsJXzuOAqO4hvJrjN044a94/2YFvA9B1NMbr
kHNSVhi9Juu0rAZ2KPXWD+EJCQsZt9O9Sp8U+tKYGRthpkSor8JgSp8o4BejJwjH
y0fqRhfT9oxnX1p0/LIzWkfBdSKUlv7NdOVbQSh4VuSHYpkwhLf01WDg9Dfjs/0e
N8AjeuSR/cCisX9qGmV5zRdYa7JzcGp63xOtIAQh4pHERrEnZLWoBGhTUmRWuOPL
K9vMASjftiEqD7ZoGLbSEHX1Q0r1Zwl77L6GmDylJnbJnlP5KbRQagfzg7VL61BK
dtLflNWhbzZEQozx9sPehQ2QucF7PnDuNP+j/drNTJLygTkR5Rh8IpE1N4S3Pwzp
1t/C6lukaOKkIcA0NazfhM9/Bou+0/D3FGBHd4ZneRAzNThczhYD80ufreQ4ga4b
tu/1Pc2EOi/lMu4bEH9TRnfce2Roe8eUcJbBoivrhkCLAcn28V1qIHbOm2RUA65q
2WPw4h7giTqmxYYkM1WKezk6wIEtHEJR9plI3yNTbDSPzff8gOjsRXuK1Tlmyief
ujcB3iEoOm1ORrU+OmMoqMJ52k+8ZEAZhvnUPmdsO1BQFSfSj0SzH/imYaVvSVvb
nBvunwv+vtZZNBMT6HDhMRleTajoEUtccFWoeXoHPKbz0psdCvdN2NR3qpgID0Gr
2+OFd6XPn5rPMyElwhq+IBj8mzJXaLth/QkWBG41pVWdkh25cRJBBv1VyQmDalwt
20fuCinoo7uoR0dVwmHIwiXUpc7x3fTaEC/+Nen9jI/q5QKANIfYA5iT2vcQFxNh
xdOyJBolc3fm18dJwweyHaaecFD34D/l3YPz4K6a0hbP1OmvfJCwOaeS99avNOUd
K+EY9rvRE8oKSigjfgUSnaVaD727Kx542UNNN3bWaW7V2Yihl1nFyeQWOFfATihq
JpycT9EUka2U4r+JYv9MaPgh6trQ5QMwaKQ8+fn74X28D0R0O9BbIjlQOOB9AsHO
36kTtiWWndKYGJlSLh9o7yitO8Flx8Zk5uAvd0ldt1U3kYAXzWkz2131Fm0vQpaF
tQ/mBP7jfJDniZDm5tC32nm3tvPrEIhAjaamHMqzdRB9K5aoYSWW0Om/R9JeVczz
SUENuhn4OH+dMawMmIU+2JiPP75FRIO5ocuGr4O1zRuoQOFNyPIhYMV+tXckLFo4
gNVR8HfPJq1EYyG3Df/GEdespv9ZG+3NM3eBBHuZGfHBlG6EXbzu/U4sg26Yy5Ms
3+peunG33IxV2e5IW+Xx7lvY/pjr7tc/pyijmYVtl2gBSumsgdh7Gxg0Y/mYW+LO
aqgH8QQ6LOHWDYfwhTYi4rdauu82B/KUtC6OwbnBrOYAbnYEu8dY7czOq4nIVNEJ
c8cXNFAMK3Ezgx4mBY+7vk/+9Ac0bBZ6lpS6C5otYJ1ZIlVBBK/jYqEdxk5YqYS8
tD4WvQoi8/NjH+4WA1XPPPOA35lkheliwK6zw4w9GR/aBcAuBrEoQEY02iStagp4
r5opcLkB+OgpTlEBxwmypjZJIgZm4Dv1ay6+0i5zOPoujNPhReR1TGfpqdVkHlWc
LTUs9B9zyAVmZTqTCboWFNJ0Iwx30AdamjlLtuPX7cifrafhmX4HCP43Apx8GD2v
/RUysUQDn452qV/ctfk9X8/EWtT1HSG20EOJer/N+GcFruaImYN5pD21JkBwXOGk
ghskXnoPff6BuMpxr6rkgkGQDwehxBB2vGMoXzg1VpQH2Ou9GtQigfgFt8NW4IY/
+j5+UiPZAQ0zwY/KPEkKslAMoV1rmoh/Z/y5W4hkKuO5bk/MJo8jxBrFOPVyh7K8
F7GcN/MlXy51QRv7K+goA9YbceTlsqiqpugbG3ZQXybXYEdWm6aMXvLeGIvp1aea
IcehiJkFPeSpFENfYXvhULARrJvg38aku/Y7iQFdP98=
`protect END_PROTECTED
