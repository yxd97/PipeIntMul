`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ysj+BbTOCywKcRgYTZahTA99G6HPuaUKuYKHNkOd/pu3bVBHM34zCiDQxQt45mPw
dvu2VPEO4rSYjzGR7FAj0BaLLBmU2WGb6yIGtjIbQHkQxcuvB4rqGF5pchIFPcne
xXNhwx6iI9sJprNlwMeHWKdi1r4YvlMzCcqtpz856tcwSoosUc/YSzC5yqXhNVnC
w4RTDg+/VF2Uleju9gISXidLeftHBwx2GeVScaYrO2VI2QNKEmCp7rEhYRumqFPU
GR3D65j3nXCUJLsoFkIJHRv5dcKO/IK1QfiRp1zDpeg0fuhbArL5SYu57Ady7RHT
T//P1uLoq2bISUS2HEg5GIpWNzMz381h57l6pJbQN4G1wajp26JlpZ0UT9F0VvVE
+X29n8c4wEeJkSLbvyhDPQylGPWIFyV6BydkkOgpXJgbk5lWqqM9ouFNmDUMLSh5
otG8EQEYoQmT5V31pzBAsLI27hfpf8gKfyS97JdG2poCVDzEwCAE+Aw34U+zVSKO
`protect END_PROTECTED
