`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/keDQ0R/lUI1dRabfUp/roRoZEjUUSP5IRBn8fW17EMbrbzgGF88st4N0CB6i8Z
KnX3+mLL6oMHqxiUVf/Ru/DL14N3EB9V19HenG7BXvlyy5o/sKkk84w4eL+Dq3+Z
txQlDtjlXHUFO3XfFtYtYbTy8komCgRQ3jNy9FVfLmAd7H/qyO7qNazA+nQw4U5D
s4Tdi+Zo6Ugv+0rKQGI+wYMTF45eN/EYCZLtXwfoQj38mAZ/mSYm4ImjCM+dwmhQ
9EM0sIzADPVp/CJALTHAIX4fCaHf3o3nDuAx0fvnTzM=
`protect END_PROTECTED
