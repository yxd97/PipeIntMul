`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
anbcUI0V/bylyV6NCDvpIMjOpSmCipDRCTPMI6DUj3+ApQvypBSfGAI54vWhSEVT
lRuIQub+58E8fIFjEXktDN736WRulQccm+GK8f4YVGOD7jv2ZsxFahG8S6dkko78
MstOOMzpc6qXjEMAahCLOVolVCUkbatSzdjfhyqDwDMd3MaqRiyzfFPgOIBJSHTd
J+OltieLI11kGfX6I1moruvZpXGSmZtavrTu+U5qH8PNTx4bc7crlOnQ3SzIdv/r
Dx6REGmq9cDZc0BB5zK3Y2r4d+xfy0JOvIKmNb4BE+1uvPvExXJS09pNTjF9Kyo0
HAGu5Wnk6QK/Fwgzfsr/Ekc9/D3T7YKn8ecqKU6ov9N9gzsAr2zAGDCdckNs2IB+
OF1IsfrNuz837Uap4n9gCkS45AfVVEwjbd8NBxs3tFLi9qpcp9nYFmPLJswstXzu
HOpkAVEIpzbX4BgL8EGx8hBYXcfwUzVr0g/7dmJx9ggKzwzLneFCzmJ7aWHzSsbc
YOOH6y2qzCP0MigN2UGkimcswDiwLk3gzLau3xBAkqNKXy6yFMzOisYpmg8UsQjr
ER1ZIexqvhQhUdPi7SxqbcdJGeDgokO0r538ufLqqBgElTd8qNn+1gLbRZdfAcUo
yoieQlQDN6hdokDwSYWBtCjzo9xzutG8IXaKMP5nWaMyBrcDCeaeCFo+HW7CbU+3
pxhylyajvkSbIoC/27RNa8efikOeTZWgWLzyjIySk8lt3uoDcAZDXU3HpqWAfyfV
wfqZKAyXwlmfRT7+JmHIB5o34bN91uClN4a0i8kyxYZuozswDH0UGS2yLWQx7eHc
tqJHzDNV9mtWUa03H8lKeq0FqPI62qKYUER3mkt9ONfXkul5WcqAaVC734IRwc00
G6F5dHf/ifTSynnlhhmimLQTkP415EK2Yf3gQNkz53MS56UhVSR3Hy+GyPz8qCAN
toIXuPzCXgs6TV0p/LtscykeaqEjgbzV03CuZpETXWVaBo6xtGdJqNhkRSz320u9
J647ZwWI8Cf9cPo4q+VRAgJ6A6qiRX8QbcouqxvNt6ZLkdmNrxzcH2Rzm51+VmhM
WqZaFR8BJd9rRhQLB9kir+I6DuTKNwNhiC0zxxVZfzE9x+waCSbVBqyGhOf6O4Uw
ACXAcpbWcmdfrZTqzNcQVewwE6wzZB8YtgMHubitLJIdVar4ZbrkIeUKTNRE9pBd
8Oknp2s5QhSGioD55CVY2bTid970CBr1sA4+fOJmGejpW/dyxIFTAymXmnFRSSFp
mOUyJLpo4P+565NVmCIh9wpzFFKlZPhWcMr3FbXWTAipdmYd8A5l4GQBGCTCNcj3
Q7aWsSFAYx8dx1vFrLStQJkgPqTg2YYb0MdYnC6/M+SrSpl4J9cSkko52vbR401l
2bgvpMNqBydkNqJTprFthUFgf8UpgolP9dUN4hdkQCPIKioAgJ/JVU68T1MCYycK
6A/PWB4c7uNC2tSj7hX/X6U58pIVsLZVPROR0BqFGmyHC3saFDNEcn5LkOYW1Rp7
iS22Pxw3BpeUP6MkUi/Xkluzy+/LPTVPOv+CLgOWQ03/A5JZlm+nBKHiaO/RrKuk
lRlYjVUYfFpp6jbpE535Enjiyu623CTvEcM6sYOS7jg0P19MWdhhbi/BW51o3cG6
BY03RL/EILS0cx6xdAsxANXc/ZqbNYWCOpDVP9zftWbtUEwn3hsV4ET1b/NHgELH
OxHZaeiLmnpIaRKLkWQxZ5/VKkWuyst1HGqwy0zrmje45xjxIyTBlxOcOiYY3Mnm
Dk4N0dVzRpSuXjpUE0tbUaZZjVzSGq1LjU/tcW6VLNN35104RyRB5bE2LUsATFHz
50LplbGcBrOgC17w2XujxQkYL41KQTdFSWFAyvmwWksyXY3EPYlkeJql86lZ1Gh3
GfyKvRu0rd5O3TqXzkdv8Zv9jfgcEoPchro46GEenk3FoDbkNzf3lMsNpEIJh0Fg
bfSxsdIviCG/VooEtVKjEQ6ShNK68uo3I4wB9PdNLsmbCFS7Nc1G/jNWFm+s7yvl
gC095RvOK0EagdApLUTXMl9++tKItNw3USRXFlHNTeZi/k6czT6ebaXcyyZ4E/2O
`protect END_PROTECTED
