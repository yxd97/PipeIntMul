`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9aF1hWOfPBiUHdzrkARnCXNKAsd2w4F8EwG/ubS0QtjQTmOJq0IUkxBMzsSlHIq
TT+ZFV9UpdR6H3wr6QUWp55b588TNXJ7r9tbyLRMv4Utq15nTRGcMJr6QCpZChj7
mY4jKC4Wp6hgrH/giZ74bp+LrXR1eX126vWMULGn/nKM1CNwzlG6d6xY/MYIH9aG
/61qZyRn7DUg4/BqfBi+aJBs7P2BihOvw2iep/jymRnlAhsZMhZtWOKIhqOPKBV6
0UmFgSqKOMnrJdqctcHiodMdyTlWh5/a8kltDW3U6Wpr2MM92lS68e60Myfy5YVj
sBEmEVJ0CnpRr8fU60V1d6Kul7XMhZ0dIV06Rsw2xObgblfV0dl++lB+SRVNdgbt
j7/ZuoSex1sC1KyuTlqbWjHPpJGUyB2TaNzOu1BRZBfO6067zBGEGVspnEZYod6k
Db0grLqa+AWoq90X8dZy1IYsYKUX4Q9jk48KK4D4wrX0sRSK5UpWFRNfy8ukbn9F
hHPyyC6/lh5isDV9c7wFQgHn82L2MKVD+rjDDOnSc17SSGLZ5S0nS5YGmcltJ07Q
C5v9Ga78yynFSVypTFxgQJ9pjaP6ynoFw6WvRBQ+nOQ=
`protect END_PROTECTED
