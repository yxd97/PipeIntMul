`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P1lIRoFErQ42b5lEf7d+TT4Yf+sI9wW+tiB6KKTAp/jkzpgCCkLpOZPoxyg1waJi
U+p4xnDAGX76kiucrRj8Ijtfhl/3l1/3IRG4YAVIBV0cAh3TFP5vWQ8S7btvI8Ah
uBrzs/2qeoj++xcAzPw82UByRhUvW3mcp8x6ZgAfeizGyWpVmD3RPkAy48YPUNIX
knM96W9pbvbuWOkm7Xsihs+pQENbTd4HslIRrvTrWh2vgGMpdwgPCMUj6l71YyRX
shtkYwO860pIGA92HWok6w==
`protect END_PROTECTED
