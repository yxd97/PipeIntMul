`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cB7Yz+B6rKpnXHXjN846QRlGzCdTTjkaMF7cEaWHqFga1QA2FHMlJkKPdqGNooVa
8Xc490uzszWtuoGwuXSXTGcL64n8W4dDzTkzYHPzsOaJ1zbrezRO8oXRncsRhKce
gWZuiOQQzUX9RZ/1IJqscnlh5Uqlssg5yo6ewKxnnB2sOQTXjHNmuJ4bj2hRZRJn
rOSF9itdAaYbowk4GyDcf+RVpqVl1whLnMsPHc6+9vuhNu8guicBJapCkgwChNnP
CT8tlKAiEbrZdUxbwmOseJq4IB30H2xoErND8HT/WcHyF0hjJN/tm2xvViQ9lor2
2Lg/uQf2gsw/RodZXoWMe5j/z10DaGxCL6R6FB8TdwxutYWnhzRls3FHbZ+T7Q3J
azIEJoI4VBurEyXk7+NbmFlN+a3Muh2LhEVPXLnfjCLI1pierYzNugsfzGKLzsss
TaRVjRGZvetYu6hMO1Y4385nKvotd1IB+vOlLuyVeuIvV0uH6zsVGp9HSNhxEqUS
BNVm9rxccaBSQbluSKUeIIbSTiecuLrfJqWQQqvUw6WMSfslzn6lW1WY5MLJrjc0
`protect END_PROTECTED
