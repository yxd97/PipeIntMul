`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i5WalxJZGxxtJ93w3F5PRolYrBSNJZdUCdxHq6YbqE62xTPY2i8dTCYJQ1y7L96z
mpDWcdP3hNvz/ahpGg2PQGDRC8W6XFbRw1pSbId9WNWXdeYru3jS25+eG5VU+jNM
jSKJZcpEmwV7IBawzhHryzvUjLScnJEmaU9sJ5VtK1eYi6aWWq1bJ6QQ9xvBzUcW
npVn2Wac81+Cx5eXi0xw0tmjqFKe3dgFeZIQBf9SuU4LPttHOmgUgtO7UQjmVDTi
d636Ok9z2MLCYOghVGwMs4evDtRXYue0Br5IqNycR4mjsAYdE6rCSZNLVQ9he7cx
Qm7QNyqa8vsZZkW7Vq4EToanAdI5Uu7yElF7Fw5Mpd8HjbVMwk+qaEOa7mmhfyWP
GkofIaPGtWobW5q7YulWjZNgXu77yi3JAdmvdEBOZzqzFQukE8nGwJhDfGDZLP4q
tTtFbFcoGXwQ7w1esItiT9+SRx63Pld8+GSiv2FHIjS+AqBjg9oEk2B07qat+3qM
wpNWiwnAbZeG52sxsK3tWUgahCsxx1XaM/9EToLqI6WPXGbB2g6CwBmxO6HicQuo
nKpejOiYBMlXvIN/WFKBOw==
`protect END_PROTECTED
