`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qPrWGxVysE4GwX7Fu57wSyC9bLiQLYKc4JR4VK7Q6xRFmOZ4rQEwu2I4zInkQKj
TW78E4+mStoUu/caJl5Si4Ov/a7kHNd3ZElnA+ggFak5RgEPSnu3xHV+DtMW2B4u
Vqtfykm/DkWjuwVaP9HDdo6Z4reO2bsNjdwKRSguvfL5jbNxptXHPGpCDXEFySym
ELmYJsP212jnC2fFddf3Ll56qId9Ge1Mur2hTm/XNV1cT3Tjw5Kkvih+DAYv8fe6
JniP3W5OQR3I1OCrbW/3IQ==
`protect END_PROTECTED
