`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HFfQdeb7As7U+szkajNiwC40ozoc4HXuHupi+7rlLtDVTQ8k97u8CeFhVN5guSkD
LszdA+Iw5KQXeBnu3PmpjTnx+HAPlnv5+fNemqrstTLXdT4HMbcwARczQWgaufsE
5hH2jDR8IqCYyzdOQFHiWwcqfyw2wH3FESDnf+5Lgrk08pMxmhqSnoT//6igvqo/
VlpwpM5/gVc4LtBfJOgwDqcg2XsA9BeqzLh4jvH27JaPP+yDsAUQNqECLKtxlPNJ
hBGt+OS0lCs64QtOzFrn/2l/5nL7EZ3SAw5SSZa/FyY5yloPemYq/jmMYvyTLwrN
+1Eb8qgwnDDmSiIrsa9Ff3Ch/u0OOKiY68deAPUSSeaW7gnozEvuFmGemUZLIpI5
sSkwR7PUWhOqGviUkpRoYXtqBv3/vvzvrWeFcvXlb7Y=
`protect END_PROTECTED
