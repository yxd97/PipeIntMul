`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2P3CHt/P5IfoEBJ7LLsyhREaNSxQnwoNpsnVAdcMOF5RBXWn0IRyyvBUubfD8aNT
WH+r48/HcemheD7R8ZzqxI3KzRRUY6ailIqfzqf61qR9ZG57ZA5vEFz2PnMCEAGc
WmBVpiuOJIV9wypDkfRcoxDtbP/gZjHBjQXo/U9Ml2apWVBkJ3igVZHCcLt6zYtc
T5QkR+JmHJ2n0eUR6rQBrZNuXthU7p/aAXMYlAlteJ1thm9lpQq1W2Sy6IUxruSr
AZUvRbYmMcBHQ1rTepLAckCeak7RBa0fTnnlo+qVKkqEGerEENZzzgD7SyfZLGWD
eFdUJCXEhzzTlOWTvQ1lGMFwhpdt2MlEmjWe7Md/JykjP1SQPMZJ20vCOpfVflH+
D8nRDOf3w/iDerI64Je4HgsCyjd202LVuD/lT4gO+KzBAGPGL0FkF7rT7bnSWOU/
+T3YNI4iPpiK6WjYkklDIHZVPQrU/HCkPjwQ8fWwqs+hhZulJKHKHUHvEZDAZWaW
feFSAL/jBxBjd0ff2IJ+k4FcJw8AO5PoREwg3FNuvzOHxFMQkhXroduVreqqEQ8z
ipC92xpsZDxAkmINM8xpWAWguEicx+u3ChNtRAt2YMYSlW2QQ7paehWju7jHo9QK
d454MeElw0FATZN5Wb8QQ5i5sLXvo1qXriDOVO3+PfN4pXkcizC4yTdoEwvCo8t5
24vRs8SYE4uRzV5D3lTpeSM/+P2QU5hXfMReU/YmMiZrZoGakeLzGSccGoGcAd5E
tcWIp2cwRxWCEPduoWMbXMeqEWtRmVMW7rKgYI6/LCDJMsRa9SsRvMFBS0fv/hIu
+6+DFxJjsjWfRlz53+wYAguQPJQQ72YxBPPsSSrOpRG02Q8i2qiPe2MUyanJx7XL
5n+uSZ7jUnFZT2U/4RvkQaVThFShA4hKZZusMgZ8phRnECl6KDpJMg68hXZvq6ux
f2dSyDLDCBCWxuilMMcf5/n8QlorWbS1e9T4p+AM9lIXKoZBXZxjv6wHgFZqrRMo
wgedIc6T/EeTV7DXBQS9Jut5i6mSwd5piOIVC55JUTrYu+/1AVyf6zsP8enpgJaG
RpTNfhhKLNdCa9Z0DFucAV4dWulEMd/tyx5+Ei/q0JkgpC6XBvjWbB4aa+q2rbaz
Ge2JI+ePvyJhtaICqiTl9Bvc/WahoVSVIiPWmFM0WH0OSkn94Zm63Cw3D5OUB4s/
Kaiu9C2IXRCqtx7Ip3kOn7BP9cgzt2PieRriUg7DoUDmdVY5q4wTGNqGeS/9dAe8
bb+L9AGEsB3H/onee8VKTmoWuB0NthW6TX9fXfbEkRLfIt4GLifYSy/Ao0VrGIu6
uyj0u7t09+LmB0mgpuz+0B+on3ZpQ1vl+UQRjdJqFMDj8VimzdBJXUTPULO+Ppfv
hrV1uALohUE0phBDA2CEhj6GvxhclVs7cM7kRrjcAfDlLil8Ibwn5BfNJG+2DVtI
tTZ+iXtS1EhBmbrHqWZ0y3pFX8zrlNeFuwlLGDSBRlmqNybuujDjWwX7tKyUTqRL
lnBk1rwC03S7/FkuX4Lv528kSuwaaUYIeRDH6R20QY5oKV9c7Oor5Vvr5+y26pwA
DXZ59yYUN3kGElHhpNBBH9B9U1YvHEdLD1b1ubXZYLIOm6G27jEpWBw1Iny5i/xu
Zyryg8OJqbDYDOKWIZAS4G2mYPf3aVF4PZ2HOF5O/BFKyPqUOqItQnj9jni2aDmZ
kInXvX5wLX+xpGLTXxhmo+YNZT7ExLZ1H5t6jJBGSiD4FP6w8rfpRhtv7zSUA7Bp
LZtx3/qNRlhLFkI5giUfdOMhGNI+1ayb8I/GzNYGIgPNdZWxSDvDDiAuKbfAiuIw
rPeALB/lZeljF8vWtFtz1K3oV3I8hWaZnJcs8qewMiSU5YaXfAzjHPbZGQcTZHjy
X8vIsIsefxdMLM6OQOH+dKWnzGE+FiKoLbVOLLCCQMIMqBKW3kycEB41HOcwdfKe
Qg8giQ9HCNqgio6NexmIqNX/ArtrAfzDAetjT7Cxgy4K24XxpTWrm+kNsCoQY2D0
8CLXaIAHUZNzxYX43JnSjqPWkeJ3wpGw5SxaP/jWJ3Nufs4ye14Ea60vHhSqvrrs
KuqKafB/2HgtWnl3+Pg6ITt3+k468jdHd7R5HtBNTj87uuR0B9vSnPhCan+Squ36
enBz3iUrLJSqOnaREKo+GWzMVqhdmz56dwdFln6mw07zTYvCs67w//IlmbZ1aOd+
fOU5YF3q+6nAzw/YfP+RShAw7BtNxHfalF8u+MR4Uqnj+PWdQ6WWWamB8bCCC/P6
Zv6YxvG0Ump2TGn++jGkJIbUK0zEKfS4EVy1glqwztQK1ovWQI0Og6re5h6Rvx1O
ISRb/vEjcZnVgbglNWZd5IULwWnW1CrBKC7U/BdQsOgYtI3F2v9czl3qxbww8oYb
7FZhcJJ7hkO8clRqYSg2Hw==
`protect END_PROTECTED
