`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWTjl2zV0xf6bwMU+lCs2G3grX6exjLiDB10DFc9LURq4STsA5vF16hov0lwreOc
eP0PLdHw/zmGM5HwTtLngqYo46FKgNl9CGot1HBA3fIrQta3zUs8FrW2FCm2DFqT
SuV5WKHbiWS1q+CzWk5Y+20pxSraaOns4OtyaBT22vuUNWfOukx/HnQ3mybSm3ij
b0dXGxQiGOCn9ashoib/lZrkHvXzNbFMrCAunUwcNpkb5DnwsXXApEkUSEC9H1CH
sCQ+gtWbcpLzvZ17Apv6NB5GJzyasj5HtepGtr5Q0WgDAvuqbzeys1gK73knCIDT
Bc3+vt6XytekB1wOZwsyIlq00Cnf8bKoxVBBFTS5dql0pplNs4gJAEwSeGfkg7O/
Gw/vQUdjcoO4ZPmjP0CTmkYeP2ifXTgB7U1s8CXbccb6wjiU7FS1afYwd1vnhnTF
XK0iVaMLXUGrCLYnpJ3gBxeHRANSdqebnFyO0LhZB6SuclQkpru54A3zV6+h4b4r
L5vDVVqCcCltCAcaVwctEJcTLO77U5eAAiQDV/IrpjxxQxuMBRJB9grfMIbF5TPA
brOg+jC/U4SqBqG+JSxyxnn/Dsc8IljrmqJnLgXhoKI=
`protect END_PROTECTED
