`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KsI6d6bFlUjOOwmoiajVupktTb6Go5h10RKtwE+pSvH8S703hss4qYsPa4zAD7ip
Th1D/tz260CDxrVpyHRn78pIA8BJAhyximCYcwyL4xAg0R79QIzdPYyFE7lB+C9n
FfLQ+nWMgDkQDiGXyXiKMTKOjsvLQUv9nr28u5LVNFmk8tPCia6uOa6RLf9vNGuC
Xrm0LpYtc3/CcDfOBLqpAmR0Bw26/gmU+vbfxo5+FhQcVuLqJTLHQCRoaZ/IJeEN
`protect END_PROTECTED
