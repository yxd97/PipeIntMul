`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cYgH/qT40X9MvLgHRSFt49AIRdMbUHcgs4niPPR/wXv5wEf403Sp9YS0QT/hyJCb
/1NqaPzCnrOaOULKXq7waEloFWf74/Z/VHBIAJPtdLK5Tbo0vE8htMd8LQraMtsM
CtDe0I/k464pkHct8+vRN0wrWOJXUEorAqyyGE+zYiGmbb6JYEptjdkaFUNlT96O
i3kj1B36eZV731ESa8nVOYJVEmZdiOvI6JscV6pOWnd9KUTotcQo8r16hHKtBP3n
CxsPP13rqBsnnFZ+pxOXUctFpSh8nVHwPphk9AlPsw93GJWMsBV+rLyoTvHFqs4q
lQWG+tYzq78IiQ0OHeKylyDX0yRVgSpIqJGlgTBh4JLBVbJa0Qcti6jszX4Yv/BA
94+5HgxtVCFicY8mhUHGoTeqb3uvydhJEQ1+ZbVV7ZWpbtFZfi1xnxA8Dd7q0oY3
bFhm5Zz4oRzhzg/Z+c3nZTKLDPaF2ROkk8kOuMPrHt/8K9tNA8oMY5ueLM3jePGg
5FdOSNBzZCj4lhm9mhA/IjEQRaRGTaubnixg4XV4wpKR3PrZKAoH35HoUgnw5+Pg
WJOBD+uZEHbNFLZEdPz4Z82NiOVE7aPai00f5mQXgb1It4k7k2Kdb5TWMZBgzj3r
LI9YaK2kmj2dMz1Hjhx89mut1YsupgajPSUoN79s8P1EDiBhoX4TmEZOs7mRCdBH
DN0yPoq0CIOnS+MF7ugM00KWX4t9JzlekqcVOdD3jdJKvXVjeVj/+eo01RoBlVyv
9ILWlYhGrHQ1EUsMNOoVPPfVoWTh4ZoVAiWOlH+UL9n9Qgd3ef8jJSXqalFM9l0n
YdA/tRDDQXeqPLLsguwjK8DmDhiePdn7Hhc+zq4L6TX9IWqSISVgZ8JvBDykE5Vi
lBT7gyuom8DmNqy/ychQdky7TavuH3VlUldBHZPcdHfKYQtBIGQLttRh6X1yb+73
0xTPKF33K2pFWQb9mbctfjiG80zWvTooQjTpAMKgaAwK+Rj9wKVzVntKqWa8/nan
22Jg/2ttpy2FXeN3awTfMycoG0AA/8JNZeHWAmACAmcU2+Ucz+mkbNxgjy7wflcB
SLmgfWQvqcTrvniRx8fC9E1YdPsZ3llQ25Gx1HRtu9tlKGeN5nJnHcTbhhXWu+nF
E3nm/jq7jlc+qaRQlgNqyCZkXOaLSi+xeSul/ywnaOjRbhsXId8OUshNx3TPbrBG
6W/NpxqQd8QyrajBgiBPCCrWme5ZXTJ6MUu1yNZHXIK7LA8cjIDraO4hfahdGtoZ
Jn3uQt24SmkbN6Bg5RAbMRtPnvptkz3oP1EezKGnFo/cofMU9JD3K/1lRe9hubkg
jIR9JARJWYKOeA5Dk+OO0Q==
`protect END_PROTECTED
