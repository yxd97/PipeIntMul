`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cFjnG1O8Exjcn+zh7SqzBXTbTpi7mVw/9JNws6huvAIwm6VNzzztRAYkYEAIazdM
3zUpzGAEB01CGEIYegpgpdYWzthcd0htHPjfL2IOb6fASXetgwtiv4oX7HIzh5Fq
hQQQOhkxmMM/jjojEayNOqbTM4x+brDUbmv+FsEm3xG93VksVZPXLPkwZFYmkWzg
T2sBJoIZNTwklhqiyI0l53ab2Sk2IbnbpT+PJsPDOaa5DRgNZr7BgW4ziJsmFZuW
EGreo2fzGLtJfqV9ZHSNlhrXeD8GUgrBoQ6IpVipntyo6HERZtUSkOUlEmRxAXjB
dqR613Qn8dhv6zDPhVECOuIXCmaHKomKLR1zxCLwBEskPQabAQ6EOVNKPrkzzCsZ
lQANQ2Jj/GmbeitBF+WVW0CZZ/jfEC6rTs4srBXcl+AClhvTooBlJ3QvgRGi0Adt
`protect END_PROTECTED
