`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BxaEFHDJQj5J+XZXf+XeX4XpYGX/WcrlHRFVvx6gTIhMIQpGj4XF3/CBG6cPY8sJ
/j7RRskdtcfk/GV1ac24hbTXJZm/SOQqhmeEfiLaqLuUDiNcpPTQMh8zkIVQGEAJ
nilsuqeOiPBFx2aQNTtQRqRPMCnA9ISW4VLixs8aZnAT1VvAu8uRp7JqtQXxgqk4
tiolFlIEXeHSwuDtsupLLMIBnVTcWLdakzE1I3m42uXmlGghAbTQPTsaWYrfo3x1
uK6vgXBC4IWhp2ebiEAgk2gqMkDSs+pkWH+nhKX7TWI0y25YMN5Zd60/DHeddrNT
pNontvBjtGRTLjqWRSsnZzHpfCDu4FLz83Z3LbmhegFzWdn4rowraECVy3Zzl+yi
gaW6YP2wH2cFgRZkkRzkS+GIvX2QoFPKKy1PBRwmDA/UJSnqDbDdiRAsn4OpDrIr
2ZmdgtFg1GVTqKsWQjj7ji7hCAuH0ZQmI5vPTWcyZqo5iQ3vFJ1r76jCEYPeAInL
GSKf1tyDV0m5oYCiJLKla6R68MUTtbLE2wSu6EcaE+5OiWv/4WYPdqn+lefGRH19
rbiLH04KFUkqXmY6s6oXyrw4qc6upt/IZG3CQJK8z5OmOixcHxi0xSKKo8fVzh4o
LBOt1ibqgRr2u4e/Z6KeOA==
`protect END_PROTECTED
