`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSR8iUKL4o5zrUXU5cZPslALVLyImCUsQwkz5sbuV/N2RlA+z8Yxw6SGq3YaG5jQ
I3BcA38G1n32PnEFvC9QOmjHVERxW53omTxWFeJovefSk/ZyJ5eCLtfNX/XDRB3t
KUrswTcEaxA8bq2ItJwhCYMpitUUSJ09V4NhH+GZr30+AnJUkcnn9O9r7gzJrLjB
werUcu5pAS6OT58lEmBDIcFdzDLBbv0Br5jr8gvgMVNQ8U7WAScQaqW33/8/wHyT
KKzS8ms9W3B3CY0U7ImAE0PI4heEzWFpgwpZsQVetNL8QgN1VFNVkrlkxkeKfGs2
IhxHc8FcRoQPukB/EImstqLref2/cft8NRYrwZX0HyX0SCbsAxx3VZDKFUWLsv9z
e03Wi7nrkkhJVskxLzz5LeZXenxEZwHsa/jbbEBpquoRrzSf+k7rL0Pxt7CHT9/D
Fe6jSKjyZDLf7dlWz04yxtjg4pV8njfMUndETCYGRen5v1QNFh/GuZzyvl60NRda
7x5n04ai2P+aQ3k4WvngZhKkYHEQrhV2gYgF2ELeMLvihE1PVTmRrD1RB4PSoKmO
HOlDUOaKKg/4Wzh/f1d3cvrH1GbeE8K86ouSuSl4U5igNGT4DvVJ8r+0/n3lCq1Q
tIeMv/PKgM05l1Mw1NDSEyJupwqdzQQMEprE3QzDrJwdcyRlJZElNNo5eQ2FOHJK
DgHzNPJBc1F5nxgE4p5bNjWK0JiXqiich9Q0wNHO5bp4L9loEp8fooCloZTgAREZ
xWJzaLgd9jI+4lMbaXKkptZTFvsSsxMAVHM6CUPW9UwTjQYSRnS9GVwP+yw9lwTz
DnTj9hmftyP4hvKHcYP+u46akrVPbm9KT7PjkOnAf+Ut/I8XWShCXx9LCL90rkfG
mA3tgTYowguKJbOTJ208EfB60CucX9N9kJG/9jtrf5kVIBd+XzH/qpaP8eHxXc69
ynN0ueisUT42smmHQyBMR5vmXLW7Ykt3sIj/754r3vLZ2HK1NWbZ2ubRO64LuL07
oe1bPlnRiiRAyo5ItPOV+jzkxrJoKXCZU/6FeeJYfAZqFdnCYy9ErG0AIJBsYRLp
iUBfn0kGIeKAbcIGI3Vt8+67k0heMPOeqZgP9SQ8F1GPTCAjg6byKIz4/SojRTCa
i6LSs1yuA8PIemoPjqHgypNn+xJTPQlVYHQtNJKIZvUI4H2f/h8ElxbvZ92xbIiY
`protect END_PROTECTED
