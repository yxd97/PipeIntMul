`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QOZh0tEhU3cg98Smu1dnMNjez0gQbL+TpeN1etLZgYVucrlyejl1Nqwz9hKJyrgX
j+KI4rFmh5FY9GXPw6F1HSJkhFKKkSJrgI7NvvP/woX2r+BoegvxJofRAEu1giHw
s3oKZ0iBAMGxn9MWDnOAFCvB+lJS612GOw/8V943VU+GmC9ukF1WipPgZuUWcwAP
I3SR6MuDXW/6JyHTBPY+V7C36aXIyO1Sd9hKT6flJRHNEHYoWdhk45tRQxJBcF/o
Fp9ZnxG5AaxZTaxARwX+pB0nF4lATJqyzvxZCezm20GGRJQ21fo+chiu4NB1XKjv
Wydt342vziN12LqM+culz3BCca6P35GH52MWIuKedZgfS7isde+dt1FpyH1Mt5ct
uoqfS4phZziMtYUrpYDa5SlOt9M29li8lUMJjefHPOu1CGI97hWS3HFHV/58dbH2
OqrAk22zz+Hpywpp4+jBcKpXkfS8GTmECUavpjlyYO/1V88ZVCoc6UJqWIgwgyLy
XQjnVgwg9rNg5fAKi3iKaUm2UycjyyV4HN0p1icK7nPaihLhVEHpW0a1EVR1XJIi
0ZBaN6/YBqKkas1J4fkPgu9ao7K93xVVtV/l141eP7xefL2lLK6GSsKoaZHj+fA5
oWJLbdskmgdZdXv5z7r67jDZnGxXNN7iD7fUZMLrXnVVbRIm0+BPuIBmF33NQ7To
KbkysIh++mgDfZXGpwIfqY4WLXTvn639Z61Dt00qBzJUWJAzNo7ASQ125wzqUC7z
g65tiWgRaW4AQxRdwotM03wk0HXR7cUZNr2G/XKDCPlfjhVMP/5q9mD1Hd+fm6+f
oFIlDXNXxM6ZuTF+1nsOvc8IId9YRxh9zHOHYeYEowk8jd8DFBYECl5isof3J7Zt
FYAnNXhgQlOr2RUvMrAXMO5PNvnECnOKEcsgaGDhYMI=
`protect END_PROTECTED
