`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7V78AbYfv5xyMzwpOg1Y9ZT2bBBlnB7gzDQwSlPNmaKN0btDB23F2/DUniyltsl
jCPgVGl0bJH6UBQrn2RWHaXQEc3c34qzbBHAc2encXg/u05NGW7EI1XmmEa+WPPa
FesKwvE0grxVsxw2Hj49AXl6TVq5FNcoPaubunFXMFgNdCgfiYCK+NfBehht5dgC
fiBhgPTiViUfswU1JFqph7MTppdvMkneHLIpzwSKCXDiwWALEyZJ7HHvXI+QsvgN
vjH8TIJZYFMXNFe6cJ9rgEDhlJJk9FHfye3DVIq+tjhiIuPzLZ5D+mS/VUUguXZw
om2rMCFXqti5FolnABbSp12tZXM1nQb2YsnuYCfeH9xCieutRtaYw6CZO9FFT+WJ
tcqNNmgLSKWq/azlnsMkY2degIz6FinACi4n+1PFhzQttXbLFtaE85NY04lwP4SB
Hm2Lcbo1uBWXIbHIykZWfAgltlLiWuquAlUzfAttdlj5jKtRZXCIdxbzFfNnMR7x
T0Fdi9OZyWv1L+shNinE2myxD65DEFlpcvs8p0guz82r6dlPO2t9J3izbgICm5js
cWskn+vUabl7iENb3rqXJ26oztrOZPFj0D9dmwSaljarkzZxP8i7gWW1h0evvYqf
jD9sAuIcbJdEjJ7jiJbOfRN5yx2VGvpAgZHiL0jk4Fh+dtOAPhcQuu9wOGJYSZRo
CPlrtLoaCIoupU9+zEZZcw==
`protect END_PROTECTED
