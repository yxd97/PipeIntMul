`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lPF/Y2H76Zrgvn0geQdyoM0lKQNrsKO5MVvu4xORqvmvXTFaV1erZf7By+K/jiPr
hwINIiWwrY7VGzjk5PXPB1tKSPlDkSWffZZey3kTDmBaYH7DXnqWUazrNBM+DEhf
0CIjSDizfe9swAo2UzESX/Tszi9lxdax3QssWmE5/rjJcWImwdP9RDH7ZCvkzGOx
zsy1eRj5oBwE1NaAJRaLc72ekbLXGNW8540pvHL65DsWwmPSvYjL8v3ZDkjEiX7J
GZ4Fm5EeX7dTNJCS+DIGl8D3qiQ1Tf7hiMW0L8B5TLhViSGfi5R8YOYYXh6a1zKk
n12mHjHqIQot7STKYDG9JFUb2p4Tc1g5lCtesPn21LBXnheiVP/ynhUgRRxqFzo8
Aai2aDGGtgDJZvbGmYVtWv1qhc2Gezhf3BjMYS/igUdi6cz8FZmkXJAag1jSZWgH
kh88IWcq4uxX1R8KXBDEuQILGMhvnwI8v8nIp75w4FB8oZiYdwWqvHwY/GCd2Ess
phRC0bKvrQqAyIemOP7nU6URLUIoCDAPLXUq0x+5ZPW2l5UMKTjqteKLNOlbt1no
NwxLPhEjodvo7plpvvcuXJ+LCgMHPJV6NwBDFuADNgdRVHmBw58E5PfS8KZsapgu
Lttj5yIT9NlbjcuagfniJKCcEh5zEHw+yK2ZHaALk7bpCrDB3Bx4hFEP+TXaU3mU
BZ+eyOh5bXP6TyXykCh7S4GyvHkRq/yqqyahKh03jYk4YGRTBwqM7QKQhWJnB0S0
s3Xyn3dwxYfHTJ9Q6v2z1RhBPh0gcQfBVpPc4hk7l8ZPUqvxJEQiTsrlT/82AOTB
7fbI0qf+QPSaXRDdCOKUcRDl1JapSJbFPirlGZhv4YoGXSyeW+zo+ljZlHHeLZIh
vvklDZ4ngbJAA4mjDM8RjD7GlWmqIyZ1R+R/P/wIVaBQyq7oK4GF1vyjXO/PVGQh
FXPzG4/fEV4sUQetmZI86n2oofp2zBTvKvw0pFJR1KT96KTwdrP5OTfvqJLnKILz
h4EJdiSFbCrk7Mq5RyOCsoSPBR5QBUxPnbzJTh7rih2UNuWT6SAGV13/Oq7PiJkp
VM4VPhCIIBphkLW8MbR7kouvj2Q0Jk8G7XsCBgbXunD5GHVhrMXAyZhOT6DdgVjB
un9xwitUKIFkauXlllg0FlTfOJULNBLVOg/IseutPlaC1X5NbkTIwpBScDWeF9SH
z7ZYH4xGh/f2/xAjBfj8us5oK3L2x12Hxv6gYAC0OX9P+fQ2+WdIl2FLfqoRlec2
fm5VJFgh+fEy/as3ip1QY+5SDmVz9dq6ghhpIyzUcR7JYbDmGZ0MXxjphOgT/O6M
qBvJz4DWipLOeOscwxdMWvnNixwXJeSSEbTU+A9UmJGV723Awc29JqXihVfQLpbZ
uPCUd7c763E7XJ1rNzp/dpwBZjX99VgwiViTBdRMObQtUBqaUE/k/vWxILbWbyN0
iNvnfYz0/X9/Dh+Xz2CMn8PEP2SFD8u6rJeKjMcmHl1SY7KemMHFNuk9RepyZ5Dm
4VuPP6A43/Um7Cnshd98/EtPGDOU12dZWx/Lb3GQPBGPzN5InzHbLywTaJy4iMEz
nz1Od4wQ+VC452/2sCSKjkuSi1SVtWH4COwHVun4GdZdPO+i8bPbozDBJA+6BVMB
iy6LjZ0TxdbgWWcNUY6aq6Yv4S5hhfPwzA31GOQDv8wr19czju4A4Rzu2MX+DIUD
SqXIN+8e8MWABhjM/YRLKB7qKelIAHeFftJyTcgUdU1JeL+sIYRoovkNoIysGhQN
EOxWqj717g9/tk7DYwocFrUPP6orzdjlRu+jsiEHfyIcz12uQwbntNKXHRXyPBBS
l5i1stofzoFrubojmAyp/8226hqJjlNRxFSFw2aHs65H+kEUV4niR2FBKo+YP3QU
HrYqK3SOsi2evw7YZNnUtUu9c30quylSYYsjeyJgFMeFAaPeERwNtcBijtJgSQpq
h1pEDSMuEq1ByUpvB9QrWCAY7rxbBqI78dpRwm1AUfqoLJXUxlYlnn7TulSPUpCk
rGa4KDr1Gl6zkiAkN/CxosOfs99QYhdyLmXXkOud1B916E1KqrDNz4ainr6qpCUv
xLKT23DTPlO4/8kUNv0vd0Q6zYb8/aFEDYN7QyzvVXkb5Wi0qjDY0V1lgMRItkWW
1xoTayAo//EbJ221fpwofE5vSOP16FRYig8gcUwNOuu8w4cF7tBz+RYlpDQeYmg7
0pgFIFD8URS6g9eRariKtMOhznbsY5b/9vWShpeHESJNaoNvRaBxLJ1hTuM/F6D1
nPbyun5z0ZONQpUf4xevS1tMGsoRhPRE0Ga+3ampoJakauah8u6t8BK8zH0ACttb
WYn11cEAKESIRi9pMm7YxtiSpdfE1gV5st4qHYMFc56CC/9PIvfmTofKGXwLYh6y
Vhn1Lsnq21QEvrT2k5S5oqN3RB1Actuy+fXLT3ZYQ5bz8CLZnKVrXo44Jq5vf03D
0jjP7ewmgRPHniLO8/sAmoULG5vs9kUVSr7lWvt8WPYmlxEaYD7mB+cXTVcHxv/j
ZaWOcFTonZ2vUjwbyrcLr5QShnnfd/LtVHkTqzQVHjJGxucY1O+ffnTTzPkG27IA
05V7hHWuiEzc9HGOFE1fsS8aggoUxvk4ORwNaUlyevLYszywzA526DRCjGSnV3zc
rT2dsMDH3C9wTLySq5BRav8Gx6KUgHta6OuQAYdroiQfhD+drl2nYIBti3EzZkF2
yoTgpiHtXZpJbkWCuOOlnCoRey9dkFxXZhF92DxVXtLTIlZxYGDhYePcCU74qMHQ
ih9qSSAvhRWarq8WuzQ+5ZUJQlcMza+CQlw/47d5b7VORj9vS+6k6U0xbE6OO/4V
/TFAI/h1BuX0TL+NT2+kbvegt7pDy494dpEbcIwUrMR/1E0p4dw1py/phaKC3unq
MdyzxpdOOOItfBoMUjywrLoeSzvQaglK1hqwvV5SHGbRAjtfggHyexT2FLpbxEIe
eNYNoKk0D8oFk18E/pHxqlNiPyI+ycPpRl65iqfSZl8H9wxNRUfZ6OrRuReNTtUp
Dbw5+M1t6uhiNdQ+2WBPzeaWz69oN0XE1LJS65meMZ9Z+nrcJmajJmU77BPcdHJX
ECZUDF2RmD/sshnBdSz4LGDL/cnWj9q/FMkKDjbD8MyasJyT7sU0zJeKeoH7NI0V
XlQr3ZitYkWnJ841WLzB8eYmzS1iETt3v3JSvRF+qrKJ/Uj3AwsrtMyHvhtai82r
EVh6Iw9segGBfP0S9LXKGKah6OfMJtg/pr6s287HRlocOowy2eugbN5uhtR2eRvg
Dvm7QvvHtWZ+IvmlGr/jck7bhAgj9c/MKamseqvKcU6z2NsEplcioEbtBT3CyuCY
jmh7ZrOuwgudnpXism1gRHoBd9X2jiRdWZNhsSJMp9cV+MJ7iTLJy2WwUgvyU0hb
JDry7NN+tmnohN7Nprr0vcgAMN4HAqG3QqVX6SSiGkN5tmFWxyvQ0n2AvTFBD6bJ
EtAk1S8myucdd0M7hyXoPq+gRYwFoAdaoPKmpcurJXXwtL1lp+5T+pHcGpZbYU5k
3xlt2QrIULN9WxtnARItk8fbFd5Ix1de5q+ds+vEchU0oJItbXNNH393Kr2OFf8d
096iQosfOd8aRRqqxlxGEbTZPMFKe6Ds8Jt732Jz5jwIApHR4BoueLdQzmOvGvnx
goNw7HX0/hYSMcmi0x6c/qlyHczu+Ul5vjcTa3gNCx3mpJfTIkx3ecWFGr0c+fhI
guYZwcIcPy1ADD4xb/x2ZrjaFlYdgyrkPCBU9NjRlWJqsS/PKQyGeWz6XCYR5rHR
Caau5Ml2YHWafdez9TRLN5n8KfS30yy7CRzWetY3haBrUn/fPh1vjM5TFWsjOPgZ
ZG3q8Z81uMyM/+ehnCe12GEZiCF1Qe0+vYQLQzZQHtDaLRAPwFzvqZIFGJGxmm2t
WkaXyFSfisj6qRyDuHbzwSz9MPXKyBk+SjBmlZCr0ZvIs4QVW31LAfb5DQF9mMMX
X2ZcEGvM0PWzvKf7bLW9TZ/sxSUgQO9XTOhveQPDJi0eVaxI1x9byFvWUh2LTNRf
fxfy/9WvTwTypwGHS3zsMipdpzZ1Hc5eN8m/Uj3/0f7k+5ljMby0Tc61X647QaWc
PuSXVgWTsr5rwgTyPf0CmcuOmK5y/hessaUyzvPIXXS8uLjm8SelPm9K3mEaWxL/
yBdyhQ/ekf8cmej+Rjrv0QlJOb/ZfXlemA6HpQUQpBtE98nJ9QgK3AP4wXi/p9UC
1ON3Dv66Bb5QlcRwk6WGw2mGKB/Bg00SmqxdkxsdLzHWB53go6ZhsyUWKC1hIL2y
fRUaiOkHcY0kfyMbZAzLWwlJFpWOUZqWVAYx21BauxIFEKW0SYCygwJNmkN1Wjfk
AZ5p+i/xR3njestL/VwNm7O63z9GJQhAL9vy6Xj0Jj/Yoz8gfSIauxqCrC8ROaDK
gZneRmz93ol2hSvcHwyHFmfSg0J7qNQmqbkqafE/zFKardtZAoTZRuVSc4wm6Itf
PDyt/wjqOywmTSPTwm/25DPd1dJyPLyNtCd1XzViV+nA6k+UVp9vIh8nO8HdIK3M
mlCwHaeahQF6tnO1qVuBZJaKDwOuwXdVodPmJepgBSloyiJAuMz7Hk1GSYKb1zV+
ZyQJoja3sny4Pn73RlA3pQPufmGsd2MFzFkXQ+imcYZNDIkpottqJW4INBGcTFZg
V0WPilAaSjGhGHC5WRC3Tvf9PQ/u2WI1e6xcfQ3zlmeWxCl/xj7FxV4JmeUS8Xk5
RlfXt1nbAyPHnPXx69hmVd5OF9sF9mXFi/4qbAclmjkp89dC3H9i094Lc9mAMHHB
cqZm6wRdVS6Mq9SAT4ZxrBC9JzZ9pVvCntlIl7cLOT5NDCVn/lSQM8V2kwb0jXcD
dKZW8TWhVLOsF9UQgGbL/kOHvLa+5tv7DdNo3VV0bTAmZj6oYR7kcZFDmP3UsE2U
gI9OFhSISAllK2LjE7s27uD7U+VwEuAuEs/u4y2+LRmCiGXiFv1cSJ6I2oh+W0le
+Do4zeitJQVhd4CykYjMXYtj17dDYCAqk+7AebN8Ux19nIxrA1aXjpdptY+qGcfI
fLcM2/cIwAI1nZo/7h1tsxuwltn80jtZvaSx3Sj6CmwR55V6vwoFM3vgW04ImRjQ
A7KGvTFMPgYb4pjN4tUXfnr25KT7mPZHBkC5faLhkPs1pPSgBo9uW16hwZQJkpeU
TjcA0vZvBHDQgh0BbDMxVg5QHC+s1r6mOEaeYDWpQDsyPI9vobjS3jXZILYrkufi
q3mMG4/s58iJ2KTp4dFSNozQVrkLQIP7XySufDjXtovMk65sc0705GhF1Ko05MCV
GNrDoCekdP2HYXeN/1dWBTf4r4obM3adEFwZ/oAQmweVZP036PhBxluB0Qaq+ei8
ELjZfQOIkk2xdxzSWUoqsfTLUPkAB3VUDY7S65/qmQKSGu80WGKe1WRJ9bX1AH5O
GE92Ru6kOJ7Mjx2HymmafLyA1QmF+tf0lC1vXVOxgThQUlBlDdbOM/JlMG00dJKd
z3Xwwxd51nsx8yQEr6Xs1WujphEzxF9ES9cYD7tMwCGdysXrUmVuXFonE+wBz98o
18fq0vQR4w+hDs1sAcGZ2mqT4cnjUs+vefXPrECOT/m4SgUT9L8B94kG6ywZNQuo
OKrspF0lLFx8gIIr8GBd7FGGEI0rf2QJwdX+E3iRIKNDK85+7ICAmDAxTTlNROXI
tK09UkGkoWfQYOBDjVRyOvx5W39xXl5Xc7UJ3+LYVLSqH6owf1VJld5fu3PewUAf
l03QPuTlOlZ3jRhWAI8bM8ID1OqUd/GoLebI2moqtmh9zMJO3iWxgI8UVfAuNCMW
S0upGeJFEdQVVEBnH9nOy6TJGd7pBtC+lIupy37ELxCbTYx45STgEAISRyy/G8IT
CbjiNs1BiC1GKtoRWLMPOG9hQov32dyO8GR111dt5fjYuKZR/zn7X5gXyLCPxoXp
F4ETCykDhemieNekxTR0IXoSFWEZUK3WV4B5RCZ206Uzsl9WAoBvt67tcK2PqZhH
tGwmys+x2sy5A+GkLKt18MWg3RcXms9k5am+OEAzNdF8nfiubHR13YgA4PxiG5lC
j858dQW2gXMQM3D5iEYpap8lpZU3U4HnpSqsAHEKPXG1duNXGZMe97Zfd7nUrbF0
zxUWvV1Xla0wp6hT4GpE+VxCOOHz9QIZINzgXBBXg5MhaKTN5iCiuW3jlPx3wwWg
1Pa3OFGSRSH/3taOrnD+Jh7hCOCiOEITJcBkWqxCNtNQJuPie8un4RUKjhFc+QtL
QBWqre8tvxTjiBmz+0d1ITNRAl0cuAdi+/oUN4X9CfYIgDShgTKLrXhJWaQetU3S
9zfUM4RLNaGtx6y6ck41hYXbuF5ZGliY3DGRFJeUihE1kbum2RBic5wpRTJk5Ycq
7t9nnL7syIap5rizDOP3GA5tPtMzpjrcnwYL012S8iYpGmQTpg3C9HrfoVkJpzwt
eFpOXa9d8UmG5EsEQhscViSjTDmVfjJ1QE0GAQeAfE9DHvhPvDUsyD1Y+RXbN/pb
2sabZCOP0G2aMQJRwXojQMcLwcOzFmScA6HihY6c8x839rVXcTgQjlXJLy+TdfwU
r35a0iKIDsmz5ZLC6pn6qEgOUH7nYd4Wg4UcmYBa0WiqTum7/SdAdTnWTDxDHfow
1hwDCPqHQeFHz/2DLFxz9DsCZyka98LNfg7nHWEIUYb2BWcEQ8mhalYypkqKBJRK
n9VDlUIMlPp9rBCGxsyXRwuh7iqTok0oez5ByoywFmy44ACbT0+pyY3oftlekBfP
tEy09g/vzpvWnc3hIifC182nkhb3XTVVQtsL/0owC3Urs8dWA2ooFZrpHhklxGb1
vUuSfDO/sfeZkoUmAhkj3pplL8OPj8D4i3fYnCTcwVSuG28rPHfbuiImaeoShi9b
wkmCe52a+ZibpWIGHxaWcFJHDXimMNz+jA0wEeAeGVFW1TAACgSv0fOFbgXg/VYk
SkGKsDojpxW/YYeAiW7lQD+m2zKdDJg7q7lvaMk2Rledu/NfNlzY0w0PN/vOZRUJ
nzsFxHPjXd4wefm9Hel9kR2W/QW7hqQMmJATTqhTkUggS8n/1/ZbtUj5ni73o8LB
YbAf0HFx+x9nQqnsM3MkjX01woTqreucsxr8uJHo1U17QvRyHhMXz6w4GaVJ2My4
z3GPLnVemLWcQofkRUfjWqMN3x59vDVIu+JS5ogdXd1MEf8KZN8qj9O4BqF8IFTc
uXpcnqNAlVwI98bCIaGLzaSJ5ve7wyhIzoJP+YF45kAuJP4ule8NejorKld2xJaS
iqrR4rEbFPCcKjKTElWWsP2wwjfZJFLlAHM5DQNSV3zrQLtjta8poMVpQGlPCSk9
aZ2AoU0XI4DrVjLsF3upvBQP3l/lWm9y75z/yoReHT9Bort1OvJFhX21WolDmN92
KijT3dlYbmEEgerQh81esHhmok8tbnbW8AkYHquct8QSYAYP9JLx6awtbxk3adNh
YX1WB4gu5lXSs88kTNQlqeG9pPxmMLqYBCDjUl8wy0Ee0J4+DDSzdO/mlnQ9/cFW
Nq1V5l3ObbLkUcrvJ3q4FpMbghlva7jmxTBiujnNfpVaATOUTe8IPYoELWMfdwR9
zjJ9zRlBbx6GyYurzRQP30a/ajXGO/Ewxzpk2VqZMRvdo2xfSZQy/A4F+pH2agWT
SXX1uhgA9pcXAElJescBLGXJ8ZIJi8l2OvKhepQ2GvZrCDdDQAZcaELOa3X6j/Lg
vR7nzoy9DPbo5rivAndEKyuzKuuLSkZio/+/qQ3RLWtNYAxsolShJcEzvAfL+fO4
QimtPd9O1lezeIQGewk+LE7tv7pxjih8QabMkfSb6D9b4N2ZCTEXaJ7PZV6PEO1Q
IR1CodxCb09WYy6BjDfhnnkhJudUvbbAfB66DamzUHGQ6fCGlvu1mlIHwlrYmMhl
S9hN079ovaSMRL/U5S0e18/npymXmqDPkGgIaLzO108ndVxadqn8ujuKhtTJsP7B
G+gL0LbRQnsJa4XLCoD2+4HFxCrjYxl4FIwkClyu2dd9ee6WX8WuiyrM9uEk5gnN
7+qygjOOF6WVp7HWefLcMMR+rKo/yIgJHLxMmFG25Iveh3yFfOC7r5RSkckLvd69
uOtph3ZBn9zfXdfz+y7OeBxyoDeqVuUip9pXEaAgG/QagSPVfIgzHtiC6QNLnuhF
CfKSh6djsTWQeyvOFJkB4qExHPO73bedOcEv4hSJxzZTp/fV3Nckc+aQYPD6A6uu
AiyxZfX9KSurR9BybWFilGB8x1E8fbdDn0pTjirtp+n9ijYM9RadMM427kFHXzF2
ITyvY6+Mg09yQbESeXG94pBwo8JSvXRlfJXFgo74moQia6F1VpmspQL5m0XejQ2d
BH5+iRbu2UOm2G7vJSoCIbsk57psL8UsF06IJfVkm+xgdYjj3T6yC6posWnaq2Jg
uYquzcr2UCFcbquMdWR8ygj8RyRCB4nusI+EXcBBotpfo1vMAQJ8NN8XOZOR5o/3
8HuVvZYippTKEj8XrB+DKOCkm7jocVzqszeGNLP3GOuf4n+ynSSpZkiX2aDg4fYc
iKYvIOJqnt3Ba4DsJxJFTWPc0ks+zO5rjyLTmEv7vK8uVyGTZ+ciALRJKcTxp8br
LzKCxmUJJaUrKcPvfxKrjgThkkBjnhdyCP81Pe7+xKybqvuGOx2/Wk08BZauLxoY
r/d+MiPH+CjYET2doxvE+W5q4XTD9tfgO9ikgpTvEkJ2aOUsfQrDfTi2Vn2vMc46
ImXT6QUB+pVakB9iLKM4oXhWsy7jbjZCDzGwpAXiOteQ3hDzmQeSs3u0pcRv/J/D
W3fpM3PBplRP/wowxRuWlj/D9KcpjodJ1ql/vwNKyeLha+DEjd3NyyTPmURB2Dlq
pOLcaMfHIHN+OPp7mzqCmO6zwup8oBdd7sy2nldkOtTXSNu+aJxbg9RZA/1Y1BZl
yr6SIPgvl4UDpYd8oq0fudZG9+HRmOlGVlFrckZ6nOBBc3oF0Z/UV9eLsrJ6oVu/
Wweu3tTPtZKNhGJb2EB+CZmbqJvU4fa1WbF9ZRw4mACFQQZuh04r2Xs6t2SZ5xul
oW0OYc3UUdwB9bjOJJWup6qfDIN5xKG/1Hh4AFjziAWspjFKVAjJrXHHPEJEumdn
Is7wUEKVtEkJ68t/F44S/kTfQYvynRVgQkoVRScpmvQRilJg3oluL2f9xUMh4QaB
KFW0bnSUvoxoyjwuiSt/Oatui0OsuaatolRn7c3ADHlQwjNQoVC9XztvEm7QIoql
WIhOmMgT5+m5ZPgJE4eZybDydyDxKLhV/SK6WvgT1dZQSdHzU+sulrjoWQqR/6X1
6/r1rPaXjzHH06uixncFL95yq6ZNeEL7H2fBn8FTPAEy6qOdKxJHtYwIeiufYYmf
oDGRf21GyMSXT3tjzOpRxrET8vAA9TTgv5BfVGronejj9M326FrTtpbBEfXb8PGW
ZLikY1bJoK4/abkCDoBQXTPoAiQJGQyryaT6LWaeBd1nx/MCjObBKDxq2p7+Ds3g
atfXuuJgAeSeINpdRzZJMShuKB162QBsoUCRWJ/MFjDDu+a4C7p0NjROX76t81DT
rzOFYRk3fh5PK3kGgHmSefoGR9UcdjCrIMki++LjBcTBpN2t2lk8Q70zLzlRKS1B
/mjCX0QXycoloT/WZ6ZfbYjBV/PuOQE7yzfnMurYJIfRAcH1zCGurkY+b0ljTFIk
vkV46USmbQ9II/lOmr6TAdT5eJvbhKGKqkIv717G3eyXxLpQYXE2v2TCJe5ZdSKy
u51ysJegf6VdTC6Ru5kBwVA20sfR3bzygUU2G4i/n0XOi7gwZs3XmcMAmn+Q6g9/
uRuVcUu1SRZcDHZz2A4HHwS2XbxcMAfjjBiaZ7QO61wOnE+L2wQomd7cy34Sq7Ki
tfHDwY1T86bLD+gnn6id6y0VX4CUTCEV/mSJIgBgnhscqhotk6ziE4A1XQYTVrCS
f4OWK6C1ZJhyQSMKvPZ3mbAP7qzt38vYU0pgIiMowQG9Ljaoj6iag8SehvQLA/1b
/7fJQ4twCqlHOa2hyxPtyOcvourLiJSzilck9BrsucZDpcnzr3FXI2tGncNDmcoo
th4py5c5rjIDVrlYeCI5fKxnTrZmEVKhELnfN77b3ietMzew7Jt8QnQjkqy6mSSH
R5cxZWHb1AEak5mLSZAiDv1hnvu79SccXmc/VzIfHXiClkvZDcTS17RZufkYpL0p
+8B/8uIT0UFjPqy5IYoXQO9j33ey0ybhs9Gxd2ezC3Q+sPSekKAITlAiU0qn3E0u
Ono5mE/pBJtHBV/wtxYWO6yw16LFvfC3MW6GPU2sdzrF4/RUhDvGdIBPJZTKnJYz
n+j1p3LdIESZ6UZKXqICuskBSydbPkYe0MBSCyo4deZYmnGYXJvCZ5f7z5Xpczxd
3FPRa4rbpGTIUNjd6UCh80KyAFl4P52uc/oWU61W85KF7ryG1krXr5Ej1kAQagjp
yQACpmxucYIdfShAB7VT9LWohEl2pABDaUHs7kkmo3h9OKSXutXapqcLiWCO30AU
JiqJWoQLF/IXMRbsf5VE7gPkKj4fo8Bl4jzFQeJgmD2LynjMavApa6umq1X3hbOQ
U79F34UTDcUwrdnSJNDl2UKz5PejNSvHv/tFCYgz/8cTlStKO0Q9ZHHczh0ZA/Jl
PL7lT9dOP5QteXRaZDz9WVnlsnbEEw0Ue5EFdJvw/FdOTdfLUrL2fQ+DRUg6XSoN
8Uo0651EzuR6jCCMT+Ao7Rfou9R8ewhQ8NeTnc7xi9G05yU5pE/bAz/eN5kXjF06
MmsT79mpONS8+u0Bye/BpJx5yphZv4TtRx/0VCSQTmYGUZuPTZhZJeDWUbbbxeTl
DTVvKepQ/z08EhUARFnf0Fdaolu/OLLLy1XOzZch31D3rateFq2O+VB5sfBuQ2th
/np2wqEgGswGC5U2xkRCpv7nRBzQD/xMJrfhLWeFoLTSlOrdxfj4nhwUtuUF+Tj2
Jv2Lb78w9ooNhry5/LkeZggbC4aawNZqztg3PfR5FUzah7scSvWCATpo6eT4H4AW
HYQxNBHMfmH83+MNUmtdEJKTy7ePF0t3tYU1D2lwoIp4bW4J8zhsc/T5cvIuiWmn
kaQMNEr1OdZy+D55xw8e2jqo6/clw/BIs703MK2UcFxFMEku1BZX/ffgLH8fj665
SSc6lSBbB0XvSjDo3+UbdNPlmq0iyN8grj/SeuK85i4A8JhikLVTWt7/LRbPtejF
71iyZQigSjP2YmoNeod5cajT331uhXw9DiyDAcOuzgebCS1ww6pFsBDRyrpgMHop
Vb4yzn8+HdF4/fDLcDLBRveKlvE8wxZ9ISwVw0UZVNJObhe0x9T930+ncmeVXXJs
6AlQTsZygN0ER/TsUwAiUgfMyud7wMf3rHiOAUIP1+lxR9fJ/eM8dXq3IpqAy2vt
4FQV4Y6WgLn+8KgKlya5a+nq0O5Z4Z5CwPfkBTdLloovAA5Ikd6M81xlVKOBM0Eu
maWHpWykIe1moeHexcbZw25YvlcRkavHBpF9WkFRVWF5mhojQfc1G6W2VvTIUJmW
oxPp4kalL2h97Zj4iysPU+l/+GrmWxTP2JlzuTa6Fz7bMywMg3DKeDkmGAdoxe4L
y6wpSVKNQ7pE/WqHMGJBinORoVKP96ev/tICDkANLzFbuQwXhZy3aUL4GV7WpeCZ
0KJjEEu986SZC67OFHClv2kgSe6uZVqKmYMDOOhM2k9qDpRtZ46N5owYAswSJoGI
H3f+f8p3SelVQ+Dk1zVLWI/DdOlYXpFhl1fkKuFXSvKz+kvNH8AW9xtZ1tRtsuJq
iHnOxu4jj6w8CBnWlKA2fN0eF3zRS3oZRy+iS2/rAVHAlbjOQ3r+zdUn9TsW40gL
qt6qePRMY8hbmz7PVxmuvRKhH1gQX5IQSvo78VWPc87Xk82ZN3aXg59B16iFot0L
GhEib3EIsG7H1VQthkXiQpja3hQNJXbw4R5F9+5WUk0U8oVmtDR24P213xKUhgYl
EypnlYeuy8tnrJeWB/WJptMBJxgyTBwMvXbmm6SW6YYV5RjsyazUDIMlWPbF0Zx+
qOl32qYX1thfY+ZgTUbH1FerraMEnwIsAyqmEGpfe9clnIxYfgn3m2KRS8Mrauhu
kcokCNzNzgy5U5A8a9292y1SOQIjKe0lpyRMXm8HVlJoKexDR2I5zc5Xa4XGzFFL
0rZya+Z71QTh87nBbwE6WrI0cisn9bfL5V8tKOufP0znRc/Jv10jfKYC8WbxvXll
w4njRKyWNCB8uzCBhJ7fpiZqRxpeIBO5KeH08IJTS25vqDIQeNCTUepqosa9q4jP
SJarMDigGq8ISCVOGy8e/SlwlDXSS1/8n6L03aVZDXZK8pdNPBD+ulvw9xNk9ubH
4f7P/lnuT9l3NJ0j+h2gHKgc+nf8DDdiZXj2E8dD4B5saoYwbhCM+Oh9Jwg3XrOj
w4EA20ugOZFnjtemc7MR/uQhFloXsO1SRbsGcJumkHDa2X7Fl2A45MLrnhgjaMA0
36w6YNLIr6Fh+jEkG9/2YIjS9axeQ3WU3ByEVOW3f+nNmZAIP6F5ovZKV6SeZg83
euY8ao/8t9Uh/em0WuSqRY2GY91ESdsy1UwnTW9Fi/N9yePrlYXUAqZpKN88MHEZ
WujjxNYsmJ9wqN9VGfHapqGNH2ml8CxOrT3Ck9XpUz/HNt/EOjAIC+7EnLSX/RKf
wY6XJ7t6+eNr+QjzeWN9yz6DcbUonQ7HVWE47QOQKWged79EG8xuO3K7yPedMRie
zZRRtYNI9RDxSRNpGq6x5sNUR6R+DxFeuSS4/I4QXYOi8q4ABm2AwZl8rCOsuKca
e4z+6bnTB7gwL+MsBA5HD1sqXiNSWrYhhfJDc6EuAW9JaNXFsPmWSY6s+/shTdXw
zNKRbHU24hKjygkDxF+OYqGD7AdQQG2unRFMSH81khSxG/dTmn/jZfhhZcM49Y1Q
1+bi9R5/bgklYA3GaB9J1EAHs87rlS3eNbELW5BCwV/sjar/vq4sNDh0yX8d2kba
lopxP2Z8tAPhSvFksmccV4VXV0bt3TR4+w66exBX2buFODCnFmdQzkV1psHNvu3T
yjkwTtJeB/tDtNwt+2WcOZrHB/syndg+qEOHDGA9K3ZWIhZ1E8XDFh074BE+OfZV
0kPJu1ztH44lTDNr3X7x0q2UliCGNwnIKHBpsBGlB7db8kkQBXgeOayLCgxI7hrb
g9kWs9QYOhvBaPMP2ODoP7WCRVyCmwI1sCmT1YVhfcGhplTeUxadXxIHMR/uvAH1
IFIEUbKEFKw5CQn/TCCqeBJQ+tnxqwwCiKyWu+QCePK3VAOxWEPIKYrYjCef95vL
cZajM47l/H27DODsLSPwAT1S9oSI0eHhJ7ES/69fx5wbuKPv4AEaNWVVD7MruWVy
d2mpUwNcJ/BuS0fQI2k5tqIQmcglRBa30zrVuVwj03Cs7ZiD3veXLlNAU9s9Xygk
xB32Kyad48oV5QIK5axblUxaxt1tQhI0Opir/3PR1SZmVS+/IufzuAxfKfVGE/aW
AY/kaYxr863oUCD+UvDk0qOxLl1sv9tKgmTN0Om1BOSC2W24hoJDcvMDZKiWgZ9W
PdtDIIE48+i6G7u/60NpAp891zQiAcJKlP7NR2W0u2gtCHzqtaOhwQF5Fh1B48zW
SNx0y1a5Q8H/2YusWGMDJ1KtS4l0xA1mDQiF01iV7BgKB98nU9QIxKkrlJMXyCkx
roumuQcfaiN4x/o00tRHnPWiNA6cbxghs4CB7Lb28oV86pRGXl9gzdvfGGDLq2QD
5t5wf5CjOBq4OCFKFlgkVLqHRxAdz7Ym9klDKDMwtP0f104GkJjSbosOE4I3iQfX
jv7jApsCpE0irqJzT+KoBjgoHcKZI94Y+/qY+1++3qQ=
`protect END_PROTECTED
