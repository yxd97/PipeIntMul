`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B74KBiXP2Cj0hCik3DSDMaZxOe7030Xj9hyCKM3SXnkOOge1EVg8DCbhW/6HbW/d
RP+6iFPJPBI5qMbQgouJN0WbPAKWljAk37CBRv5PaiGCR5GOuI2dG6tDwSYl7AM/
BkoNcZkCObDQMSQO+b2BhPGJHR7O9wc3AjhEOyyTo1A6eCEz0z6yuF9/JdRcVXHX
tvM5te16vgam57o6q42m6xb/BP7HkT0+i8btcxvtbeRykSI7nG6CnrIKuWdWg5vG
3m/JTST57xwWTN8pDXcCuq7uEyRmVcKOKeyPdqjLt65kmVT5CZQg5BI7e92hqmeE
bfZJHb6+J8aVxB2vvFHz2SSNCr598FsZBIzn2xNWlIU9axYVlM16joN7rO2MOktF
DZNJtosHUhQVvh15KPzMtHZNz5Dk3p4/IAWxh7WqomdNJ4c9Ir3xsb3H5NU1psln
LXKkzt24dcMq8TgIvKNUfSTSa5zAT1VtMGhRr4MPCE6HDCUEO2Bq+i1pjdFi0VrA
75cuL7yt/TxeZ3pWqmQB1MCT1ahfTrxHQWrkIWiq9bQ9+sAuturxnHXS8HwscYAB
oTvBckimgbg1wMIwCMiXDqGDP7athVRAmQLGpXLy69P6ckWILIynSpKDmb4zztML
TAbR0QbATt/BD2GZeJJNaAqlPz25pwHIBa+QGtwCwxqG7UwT0zjo5YK3pthqPnaT
RP50wExsAANOnmf3JzEjwAUSuwFPrui1nYPTw+vedssMSm18aJ53oYlYz5tivflj
lxLDlmFCLncOzYIWYLVQ+w==
`protect END_PROTECTED
