`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QkzDODzSwNVg2T8JwIDoaeWUnJkdb9xBsWvMoKyR323wQQfZpHetrn/sZJZryDKG
gY9dkwlXA41dt4/Wckzg54LY75aubx1VUsUxmU2iKJtWHy0UiItzSkaQjVvo85V7
nDFV0S+mDytDjEMcJ9OnQV/gLpQmDfLLjhAo7jktKH5Ox++oVEsvMyanrEXvhdC3
Ti5atwXqI/qC72EcnjLrV1cR3P0JYy859VGtOGbYEr3inrpfXZhN4BbLd0+5g2Se
0vBn5sdC0JtfuxWSfsPIMHtHBNYdA3am42PC6AKrmap/Gri7VwyrfWhDvWYr2asC
Wt0welePpeABf1FJklMHFE6jtPTRpevOtc/0lWVWFLeJt2oFsnZXOOWX9yr8ISKO
0/o2w1L+BB57EjEplERPXeMvxsKqaj7MGZbPxmKsXRAAi3HKhd2kCFJgSPypRqgz
mmTOYH4EzO43xCfYicAUSqbCy+e8BzySICGYQXUgVLq6/oOunLXC2SHrv7Eas2v/
sCvfju0fnml54IN3WaynGRA4zwblMsa7PVqv+Ee75pEI43Z80Y421Xf9pJkv0v2T
bb9mn+LxP3DZ+lt4S1s3Vd+IF5fM23aJm1Hp5TUx+Pk/k6Ybj/j/0AD0mbmLJlEt
1OioNEDab9wh4KaUbb4AwEtUIyjyfZP8gVOq7iZVaeEB5xIRyAJtygTulZgNiEFB
ek0F9fScbF44CPP3FTeuh97Ss8wbjBeSbZUIXGZ5CZQnt//1EeKJlizBvpKRQqmn
Vj+LfAFCpYEKj8YhszlauVUqEJVu1AmrzCx5kPx7fKm1JKryhjQydbrPZppSBWa5
U+2FL1RckD6CI2M0iRE8VLJ+pr/mNaY4bsQEr9NblAaIxPApqCkbD2S3SHWZvO0v
AbuhIYTA6azRUj2niK/J4s6xhEr/Jr0GzlNP0rJBRpWkSEEB5VxoT8Oa9jkW0Dti
2Md8Pg+faWAh+Hr2MwvvtKYqrAN0GYr0krUGg/lXspJvccDcHGa+5Da49vJ9DTaO
LvQEn/GGheaaLhknwjPrDohERFtVuqr2esiuZeNvbIbzVLEy/AE9VxCUGNBCfid3
YOH4nr+8K5qU3WUw8erMcvQ4EWPra+q1KpyGjosKELCrdRY51HhTLsmhGF1wBtnc
kc6st8p0f129Dj+jqAw5icH2q47DRNvFFNlOQY79dmLMFfk9gIHmdTCwVShcVLCq
4gaQlylUbYl6wZO4ee+J/rzj19gU7Xl1MCcRLNGaVhG4sSXDZLpklw8CaZfAVI8e
`protect END_PROTECTED
