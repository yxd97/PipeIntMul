`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5AvVLsvytMKW6g84AzDvQtBIPy0EGZzEjJLYF2SF6aT5ii3qCcjr+TPEdy9YsV5b
XkABBz4dKTUYUz40nxKhsCQlEkdMbPodoNvaB8WHXrmgV6Vv7GjYDU1tos+u7gsP
G5AFXP6GywfdadvdAuA1fHDfIH7fm0dVwUSHfa809MXndZSAWuq6bOLcDIbodyDC
kRjBtJTQNyA3oynCsW+5JxLiL5p2XJCvAFKRax1jpRDAJogYIga8mseKQcIHQcBW
az0PBN4fzn7SQdcAKJtgZyqHaGlKVRDvjF0saH0RwfkcAx61J8pKQ18Yaah3+9LZ
IHMVkmOKrzFDbE4vYLq1yFwR3PS4SLvh/pps7wY4OIxohamrYnXhEgK9XEcmh5Fm
7j9meqRWUtTeil5s5/MMKWUYLbWu3eGQst/AItctwej56AThAr/5GMEC4HTtl6nN
5FPY7ya6Tdh1pEDbulzdq0/01kAtaaiysR04gmZX0P2ByAVgpbhtJbcEiCtKJI1m
zGLT9BE5KkdCYaHmznf4LxYIfyZKLNPGiiLe0fn4KKDo+mpfy/0Tf2CYk9AIXf2Y
72phhJsWlOyULPyGCkn+J+bt+8h90a7u00Kk7E8CGVug6zZgj/P+k5GCvFq0KXtt
v+PpCVUxX1KVsJRbFlNwDXqBPi6LQyF9/Rwh+qF7ih63ICsphiUQlBj6wN0q0FPZ
MLH8TF5ZkVeViXsvjmUTqGa/2DBrgXyHiOO00L1NEYguimEXzXDuVmZcFhvZRB3c
ND7mArRXCiAXhV/3yZWQsUYsZXCguqz6rvozB20wUQpvCoyXyKoPVQsjaHroIi5f
vbXnC1WWqFqmHARkh+9IaMwPjnzOXpFoZQgRABjEtZ0yqQgORW4+tWSAW/yzgetA
yab81xjten0zkB/T9lrr1JoRbnTlMB24ymSOsdkuFYy184ybCVLlvQJjv51fwwIJ
lYAyga5w33rQE/3X36Tti92m6v5ULEKgdcTpbL9kKOWNiNjSk2cpp+55D9H1sCtm
Wfk/qInG2eur2Ra0msy0Iyrf1otuMeyQ7D6BYb56VUMZYSGLMXcrGXKucSR4AfJ9
DNf0sJ82lpdte2/97mv1sBow1HWLAcQG4uNN8EWu2fil19Uy0Lfk3WxdmHpOJvSV
oR1txY73ZxcjXsrIEtvyqJncnvMXAmCYbJAIjJpscwfHzYOmDAjArgN/zaUQnEkU
eIpo0ODqntbHgpX1zxfDi1ZN4sz8883wTMGGlxqZldyMGyKmd0PzrDAr/4ELuAj/
vnna5opfcxWpo+SY069LIPAGvECPlT57XspzJI6pjwGluajI2zTzIq1FXSZ6IkjQ
KQbTYFUDoH5By7j9x67DLfQ2onBCtOija/3ogvT/pQRtkcwxog2Bx5fzuhnKugVc
O+RNNHN9xObrMSsYmYRuf2L7s2wW4E44ROvDCKm8WegjKvONZDnZyx5gOXGi7XMM
rExWQlrMfTwQMqnh++P+BZhTLw4Pn52/H/cu2FV3SKjLA7ekF0+CpVA5J9bmQvSj
O3STCOuyMk6vB1y/h126yOVR6I7G7bXsPsLrXWLg9fSwQvqWpKJOLnC+UQunMtkr
ZgPJvrqdFa3sSLjYe7PFCWCPnyFi2PobTj58pAqjR5JMaDRXq1OOMhbYVRmpHsQQ
SaAxAsrpRLmyO//jX2sIOIiRUiJYc3D9j1Q485c4a2ZX+94bMB9Gng8e+kYoJPcn
uog+IK8yoiT38xZ1xokj2rBaoCdqtIhVo+gVZ6TlbCErr0uF/pARQSIwi1Q02+/m
mTz6NfBUks9h0D9tgWUNS6LpZZvG9TeyZLGZw8WhPHQXix71s1mW6rlP3doLwSV0
C+fSvB9lacsqihEIGO20w95GH0gkDDSvxp4NCPsSD3KNeURHFnT+MyXwGRpPmACP
QkAUk0H4AWGjvPsmrK2AZrz6Ggk2Q4xCvf40AqcDSlFF5J5iCiJ4hEnEbw5Z91M2
F7/0HiOciuI3NTAc05UO+kmwUL0HuEdvq2xNxg4TsrsY1xBgCsH0/BzVDq97Ip2G
JaZYkamNNNbmUJMM/VRhVX2Q67tvQhcymAYxYfhNZIEmkJ8bvs5AHwHiO9pUSxyw
t3HeSJP2+YJcYgP2Fdw8iQV/oGAvjC5IBhJ8uSLdhl9l0ZkRUW5x47hbE8r4eW47
m252gfj69sfeC0f1Hyeoh/kXsr6c3RYVKxxFmplwIpXvJVjgWiFCTWu751m1NSZ3
v7fggYxEMtEhInZfHUSAVWGxIaaxLyHiWwtuAwgS7Ch4mWptki9K3gUWhaW/wd+e
af8dj41EAuba6jHPcRKP9lW9CTW2KytVOKAAGRUHNV/tHLe0qpKoErw3ZNgKuHGS
1mHA5jP0CWt/6okl2DRCdatYEYFQ8SfNBw1dhLbt2/k+QD3QgdAYz3sWSU6Gv4rc
lbJfJedfXOjtSvzr+cXtvZIIOa0sB0pUp/TrwpOMTIYXTv+aW0xAd2hSrLQTrTgx
fI0sEsLpE/t+kn9qoTgvOiNXNYxCDWL06pARcKIlLmWkNnrL7NHr7HXTtEEbkRCT
2JOX7fqKSPkIfjM6vYZk9FwYDHM+pYDmmMY8Rz+RS23nhugL0yThvggNELdvTUMS
cB9CuhGWiVnau5IzY45/DdtkGHU9JSo9VTvbQ9tb8TVbVmk66uQ5+dIfxOBLsI4F
CNA80ETlSrEfdf6xxJRiYKXXJ2pzNcyBfFPnRPkAHIU7mcMDQ1JBIlYXlw3GN7Vz
dVcPyIM9SP5GCgh2AohLbyvN4+ciHwpcNwIMPfzBVrIniiQhuzmUyv9JDEZyvKMU
fFsTR8l294BMypWIaqLQCZLHlxhLjFz+RNZ1OL03B706ut9n/fd0iVLO/bGY1hA/
kxmmIbE21LHfi/efoR7Vyp+O3yoZb+6IoTnfPlakUOGbMmPwRg9PxTMraHvK4hVb
kT+68cpxGYsg5hSzEYNzUmKl//RjKeqKZFvd6I6t7pkCRNEnBpMjAR5BCVL8xFLD
pG+leAs4iDxeCkQXptb1XgQC18glPSL+yVn8VxqVWPrdHCZ/7QevVa6IYcjRQUvp
QKc6jwJ2AGp/JtjtXfMOCJlvqKIMazVyEOqCLyfkIOKhtt8X4z5F9rZOTNl9c7x0
zigBhZ0avN9+n2yrYKtrt/hw8lmhP6M0ki/V4RH+SFPsnwQRmLhPbv9AhFyL6K7q
LxqUlK51Njqm98j2RqJW/BoMHg25q6KbgE+FzFJYT4FnVAef8nqs0/KLPI4jkWYn
YXm/uh9psOEt4mF3+R+cgONCIAPCeDiDr3/tNP6ZQ+ohHAcTvFtAaB7BEmT8ZfIN
arwIRzKe1ZaQOs/yQdmsemz6C4M1VZnmbVYfHebvw0Ch7nypAY2pErAd+OAJ+oQM
ZJoIBS6D5T+E7/WGN5dhs0WtJ56+FMIsVva+DbNmlPDPM11/toa1TAyEHZRQtdHq
97+0PPvobXIokINxedyi2bvQfwEvyJ9Tj8UHvgv8FwZjzN7oE89dcOeXWfeE4Ebr
PIp4qgTQGKwyYCVUQWDgVk0AVwHrEsL5z5eYXUDueJAyH9Al5+Ifmzv1A1orPBUN
0NCHaTaxX1FJHbAJh9LNjWdeacfIhAq/Zw3cnPc2t7Bh/2xihJTrw/4paNwqfZS3
X4hmqFFa9coifXaECPrpJ0+39OrK0ilfbCm15uXZQsruC9WqtFaxuNCgwb/fiUVp
x0G7fbnuAfzNFPSF2m4IcpfwiMp8HWEFuRgYzRWC7eBWIrhdZsOUw+pv80CRecBu
iORRNHNCWJFsLibUzsFvcs5Yiw6pXV5P2jggeCR97A+9OVdGXTtPsqHYqb+gqDqb
Ot7FnQ3lxXPHnf7fG/J1KojpqqK3i3DnwRRajgYLHo2XZ3GTrMa3Jv4+VZb4B+xF
r71NoqDtalLxgAFROGS972rjsS15vy6ptyHqTtl1MeFI3UMUn9219TY9zfzSnQvR
a2EREKCIdLT6eeE2JCwBG+1L1AvGxjWobDUEDrPPhUIplgHNvFis649iiYtNsArx
i0NPoaBNVUlh/+Vn0Br96MDND9zsbggWONC5h4cSt5VgcOoQ+aK+GUw/UIPKvKui
yHDbyNSRtQsG1pNQlhAJfWozm3P/CmtDEpLPZ9JkiWGsyZjUDuFRZl3zycf1f7kI
3LIFLu6edycsmPS3lrBHFvLlbUEuDrE3kSBLzhEEROe4SpS6tEX5jty6CO8JBG6q
UW2aCCoU6eejrLSGVZBkPoqE4yU/hE2u1UBSEAag0PqrQzrbp1XsPZc7+2iUUiL4
d0pBN8wJDXQv79XT+m9TMFOYhmYSVW3AbDmtLHsaHAytF/kHaNpGjn+tWv+oumpW
nm7+jvWDQXkZcPmzlBZsq2TsjRNsFJgKmQjpUBedeSwM6AlmqX6E2hCxrWl4ig9F
V6Wjsbn9FL5JjkEvpuiUj6/+dNaidUgxFqN6dMxbWKf7HhNniz/8BDE7WVFn7H3V
vkr+kQ7LRleKHgpT38Cry+YC263aFEivf4PFMf32+dhGLf+7qB4qT2dOt2gvuRwP
iqihZMDV2YP05oWUuRGch9r8P7gseTIy0vgMgGN6jHJUzy2mNE3Zomq5AAUkLw+L
YBOUwMtCo1v9jfnDmpDEjCLrimUm6t3dK/jkRnazH7t0tK3tLfGA4LxpFnVkMFSW
QLZt5JqUPwxdeCFZdKSq0SduAN19ecAeMmVTUKpmGvKb14Otcv+oxA8Z+7+FL+45
WL6S3oTyXB2IJ3yfuPRgh0hZsvVMAFP0nQhdk8Cfow4J+tmRFlRy2PCMes4X65+i
ypSlkOZWiCs02yP5zct4VEpmrZxQAFlAPu23aBFE4+vJ0QM8rPIOWDtg5I1wIDtC
p2PQb+VlPnEVB+5BX/ot5c7HGINZ3Z//vi7NO/x+YwsWmRXNQNWWvLwRRy80EvDb
9lj2FCXDTIXbMgQ76nUM2u8mgWaMy6Jm3HWqd4FVnykbL1CtNr+oNWkf5Cr/JB2R
/O15EK4jks2LNTkcmGqzijA4Hs+OXp1guLuLLUUfe7xlwpNi7Ys50s0V8fV6thdR
m1iB53+mGpbT8fannoKp6wTKux4rEl3dqDlbUFwITp0N0RFwGfKyNWG/bYjKfCg1
LtFos0CtnKXj45YgK9fV8Q5ylKAEJbFaCXHAN5GDa4aiJIprpjsJzqzdQhqXC5CA
uuiiYL9qXYntU/bqgOVkZhRvQ9jcO6OmPC1UAZsoJcj2WHgX2meyiG+W8xOoShVD
XSo371igZ6L5AamlIKL0Y9B0OmOl1Rw40zqYX66M6pEgXHcoZB/4/MQu4XqsbVrG
GzGHebPD49yvU7gSWHiWKBu7MfHeEMaJfRy6rywIM20d3CcijNrQ7xoc8bHESJT5
u41ssPISkehRXrvoOoQsfRXSp39QckaAU1h0LHBm7J9mBoP6R4Wny45LiTfT4VH7
xMLfigfw8iqX0+aGwERAku1+xLiAq3Dq200HdemQB9e8Sc5fPmNHGNixtE1nsA9u
V8QqYCi1tWtw/4SxqvhZQ6XJCQFNZUL4oOT3pfvaamaoT06BipnNZ0GNLQD4D+2t
7OW7dh8O62oQg2LCZgno1OGe+60sf1aaAKhUha4RcrgQ+pnSlkIe4SKn0XdbJjux
i327UPxzmsXeu/lYdNXbNlYd6/IJFVbk8WiSGlEt6hCurHzpMLGVBwaZnTjgaahV
6uKROAAdoGG/c+xRUrVKia/G87NEkuTaYJ4j23zN7EFC1n3f2c7S0P33h4FkgRTN
4cosQXKmKeCD73RkI9nDXsz382Ff3yauOg7NkHPTImHvZEtlh+LTcwh691kLCh8Q
tDsPI0mGU2kctE2xPsI5Am1+aqShEkwoZKMEloZTgFv8p8ScoQEh8b2tMOmlmOGW
Rnla5f7jgBwb3EtKpyRgaQqRPaE5CreRNEoLKMUL7VELLs9RRyrdMKUvBBT4hiX7
BuarFMZP0nlBFUqkxK/8bSRgA4f+g79NmX036/hReBJTaX947Bhr7dl9nPxrtPZf
eJauMs3KJBN9r05SROfXdt6SGVOSUr9LOKmPTNOQeAQ0Fe7K4YvoaMQwwhPMRRV5
xinoBuXHz1l4cTmoNs+LlCu9gCKX7dlzAX4snmToB0eSIYM5W9VavgxOUbwK0gTR
RZP+S/a9nxIVEX9tavTdX6dBuJY38qAZbE+dAXWc09fV0B0JP3yFr/KarxZJbfFj
N0scNjMGh9mftr7gCD+ZpmjnqBPcXwUg/6pPPPQbRJzpYJTCko9mNcIv3WZVdKXf
+uqS18T7X3CgZIMG6qb4U/zVfsrhSjy8Ne/O/ia1eCmP2kNaHMrzaU6o/ifdAlZz
zr1lsIIESSOcW53YyBGzgS9h5ejgzdT6TiVTKHLpkkFePZSqcLmefRBy0D+BHbHs
NrUJMj0uQLzHI6xAimk2bcXDYnhtm09WUaZWNUeOtwBr7SS67GOvOI+jrGZ+7MPk
BAZqzF/hmBdvm5G0fHMtoNWBTnyMt4R1lvgHXRoViiollJIRnvA5LIW35sBfpUHb
Tkj3YixvaEo0wakgzkktWGApX+5J9zVbd/KWY5f7JxKSNhwA625K8uZtGTOHHs4G
IOXagVHBskGDMMvRWwbw9S3IugQQ9jyUJJwYbZPUEsBQYxFcDzg40KyY/S8Y2/iG
ao/h8X/U34QvnlqutFrc/kkrE3S63oHzn6j76KxjYeWXx7yp+wPDMq5mFmlFWz+F
t54e5PrwIgqHQYLr0FEh/Ha+9brNWmSgfkDOG+br8CpT6S8sd4KG2JLVX2gFuHsJ
61pFY60dJ8enHtRyusb5uv0l7nBeSHLgQyd7ltom9ULp7G2gVR/OXaKKZDWpSFO6
m5VdXhA5xMf+G5VvcRXOQ+rj1WgGE3pxQOEBRC4SyAgR8MZuacqf5kRH3RiAMMGY
cLdyWbEEff7ISNR3HaXRT53OmdPXYZ/5Vw8tK5s8d2RRvP6vIUDO7qQxlVwfXour
YtkDwx/89w3FURewS5QQr8B6e2ffNGy7vfNP+nzD7Gdya1PM+gFAgvOC+Sk7fAZj
FMkIcuXbhDLmPqOwKePFzemfBAViO0zObF8GY0u+myBwR3feGuaq47BHO5QxLVKE
OLt9PrrrweXjdBaonPsg8PzmEyLoX2Pqytal92BlqGvAzEJ8VZlvcOCbuagmu451
csy+KadcZQQl75UfAIAzW2Iy1EGRjV2j6fbdtXDJjcmnjV9UJ/BkFMV/C2syPGGZ
HVs6BBYEbHKe0hm8f2h4X9jQHquWwCCodSe8nLhE4+/rmaSbUtyY+9r40QyJoong
8VgngCvdhawKJlcYQOXay28ZQhckx31AZHIfSIXExlnmXYQVb250vfFBpBlOhc5+
1P13wpqawENH42YAIV91YEPgsXlpnH5mofCGQIgeYhNEoTFI7a35LyBaPsArCinx
nQmHF4rzT3jfU5fHKI31XL39EHWAPSMNmeFyn4Yl3IgsrIdZcZRC8yV61KvrT3co
ZXukYdQdB4J0PJ4fLMCKZAg+67xKx+NTzTQ3wwaRqwpS60UdAKwtTvGetgt3rIAX
m457r5KDe2cNrUb7SeXGSDK2pFfYZ0MpxB6AJfm2afHroAyWo/iqdzfmf/WZIQti
djm945ErnBBNalfSXzso9G9DCv39bKMhO8mVmzUU1TBwH3IsmgeoY9WOeqLCiGWj
tmY/22OMhAw9phEnKkRnJcV5NMPO9NFxEhHmbwnBx6FOYBf8m94UpzWZcWaajaRE
KSEMkcWu4WOKnr8tm7RnLREuJ1Ie/aYm1CNwBREKbq/e7uUqXTBdHkS+fzk+72AL
5SA2quXR1hirKvKWQhihnyq1jhhKUylwN9B896Hn/CYV4fyaPKXCFwPMFHKwwhC+
4HIo9CcTY+22jjzYvBlR85N/DN7XWpVK0ANKy0dx5yPYeWSPdPrYD/Rahcd0qtRc
VCVTOICTo4a5TBRd+bXzsyLglehxrw3lRdp6JnXufoM6BqtCHZ1iOthUfVxROHRj
lSqG3/Ju2WovhTLuIboeJcyjpI1zi/iB3gAOyzhjsxnMSo1jwB2tNvwHP2DT3dro
YBsRXMrnetzG5h6Kv8Oz+4t2v59GSBilRPkWJRMgi/QgqdgJgOaSDJbXuF5Z45oh
voscWDBX6bFvzcMfS6OLiRPIHDm6KZn4KFe+CaBFT8stmrJbpk0+fd7CvgCUEhPK
bi8qEbk1owijQKzXxJFqQcOV3NsVlILtsafhHNplpDO/L9OauudHi32lUxmymNQN
ORubw+y5JNkMXE97salcZ9aYxNc6H74oL/1Vd4ewLUoO7AT6kyO3vJwCjJ19owtP
3KXqN+RrxCSs0pYz3LWGbvF5tFZgP8J3K9CXC2dKY9DF2NgFXhXq9SLW+r0f9mXZ
9lrde7swpay7KZ4pSiGPHScGyWEj0KE8FBdCJpuRP01AvNJRJFAJ7axzdeMXIzM+
6fax5p+/p9uPpwYOMdi+mVnoOXSNgXYoiNgsa5PPflsgNJYZib5Nedc3pvUDFez7
a3navvnCe0BwXX4OZSJKAl0KVRH7DFUxklQE5zxrpxEmR111d7wc2Sf2np9Qr2AQ
TZfxehkphBb4LMG0sAMOuRjwUjw9t2A00h7LSlJtEgHh2fJeiHgJYwdgYbOE5wLU
sSVt4jFRW7WkMZpkud1uT6DnV8a8bqppVRDMVeAtWGVWxNc73MLgLyJ0HtEL7j+8
qJV9QbpN2jAPL3Ir0pIYKuu7If2t18prujLEKpffFlVc6v3g2JUo5crvw5xQReTE
rA86sE/p+EaMSs0ApuYcagNCy7pZlP+UL5Qm+l8kKQZtoT6F4Pes0LOq/bHcmfCx
ApMzteYwr8lstkOKWm8aiSumOa8Sj+F9eFucX8p6L9rs1Tio6skoaVUSifyYFAZt
BbLxsrsopHnkREu6Vwo4a0aNguso84j9mPT6d9Yh94ksuhWOq7SPN4XD/KsMQ/Lq
XS9vJvANVZznhJQb+eEy8QxeEYYZXmxYDEDWtVp758H2+XNoUpw2hYoryExpIFSP
erLjR40rtmpluGWyWHyivWUMqKWxGIph41m+gmV8B1eY0gt7WH6aGcgQOgRdVex8
KGCwiUziHaxhKRbbzvjxi/Q4iDjJx51Ndm1O2TdU5uQfCsmezd7AAxx6kDScdQOW
MVrGN42ux+Ekhi8t595XRwV7bUp9vSCtVCglyxDHE8KRrpQHoPFYFgl7mbdrZ8Ai
mqx4Xsd4xXJPGBcN+Td/s2au3u6x+DeEEqNzoHoq3nJa8pZA0n1HN10tqMnXaRzw
EVWtRWFLlHPSsRT+h2T85ctxrRpyrR2OQlkLxF/ZdT3lr4WgGknzct4sr9evcBkZ
U3axP6cMIep34S43Kr291exeSieIoXAWTokDLZQqIpIJv1Sa6e1cTVo7nRwlQCxG
rbKZL7GhJ4MRK3NPxJltrU0swG1wtDhKQx84qGtzfHqSluHZ6cPW3ldIEoqB2Cj4
Oihc3IxweipVN8/vLkzux8YnnajdG+0het78lbOSW6pXM0OJMUofGEVp4dWgANDU
+SNYGRRw2te+hbWNq/y822ogayV88DXlgNeilxov5u/IUGK9FgQu7W8K3aGWZXKb
TwVqMjq86Tp2EcNFL4iExQ4RkS95n54XXBkHFVSnbXafQB6UaLR1bYlueC2Z/hfN
Afyqufeh40s1K/UBl8TAuzvz1ZM1n3v4Dkl/+27646DeN8bOoM2Pn4Cbl4DKbZAD
HYGS9YUnC0Q5p922+w3P2SYXp9Vxk/m+gO3zFc7xC+UanOmNt39jHXseaBxsCOHs
OL1SUNzTMWlMPeeUd8Qb1vwFB0iQuuGZaKLjwn7KNw4BJsLRmsgwmDToZdLX1Jb7
JOAa2VcH6dRAA8bcOUpnqfwruvNekOrxW8/XYOmkQTCmNAsAJ3rPYfW6f0xpAl7o
tFDcN6CMUzknmlNUCPvVSwSGfjmTEV63HaIab75Zr8fs6mb3kk0dCXVh41YfdZLD
zAZ2BQxg+Pe9mnoljS+GacsI8kmtXGBLPKY/gLek1DqhIZcBO2S7FsswKen/cKLT
mcnoZSXsjz/h91eGm/k+UZxb3reCpP9pCtTEEBHCzKtUEuMguAYoGV4c3zzoG0z2
4DRuAQWs4L0+Xuzb0rZ8gRT6UD35EcPDH5vBjthN1cUaDqqUTWmBiBH7GBgwaJtW
EXYEucc3QuFLj/65gxRP6+ImJghwHRilB6w146GBvZkImOMIoQpxXDeb1IDyTv2a
KiYcSUk88j77JE68L2Jgss4kZ7qsnLBmV5Vr/lFjT5ZGzJG4poJT2a7T5K9KpDyG
cNEnRz/bhMAVln4FJWDKD6RIMsAo9rDVtfA2YIwQNERi2EpPIMhjFqRfUO/KwPtO
QGVoyFP2UW9bTImiLkKAnAl4Krr+T68hi/PQ6l3A4s4zj37jOv+7Lmnu+nykJPKF
Kr34iDO9VkHH1Vx10i+K8x1+BRECPmNiFxt0QMpLMXFwxT4DUCA6B/FCMFfajNB9
8LDzCYZR7q2B7Rdcs4vGOf4abzDDuwPzqVfGXSD/uL6uGsXxvOECzMrjVX1ofDw5
dNBdDrXZHYaatD38fY9SpZkQI+4AusoS6P6u5/zvz1RK9WdFWSj43fl6Y8k9sX+3
1jSNES7f2ML/sE7+HnLPHz0jI8gOiMblhVMY1WEIPLJDe6VZOKOCta/UPgE1Rmwk
WLgn0lUA4RGM2gLp7qd84AwA4G7rLIMWicpcE4lmywPX9u7BfrIa/JyOEy94aOb1
pAG0lKugaoHR+QzrEpzGv9aSpvx/RvjQb+hs/S/Z5Bfgrg+LI27HkXgFylZc3E3m
DxiHwUZSYgSi73Azzb0mZqEdThJkJMlpaoinYKJ9F+f/iBJRKgbcTNUanVgEp7UR
o1kdeUOhY9GoOxPDY1M0wZSgdnqCpSZBeZA9C65fKsmISc1GS0LhtqQwQ9tMOSMf
4dRYrR8S+J4mgwqO5zWrUp8z4z3OgTM5uzn7ubvUUl2rEV+4Om/3cn6wc2NQ1QgG
L5B3B4k2aLfex6ypRHSGc44DmGbrPNSJtliRZWgD3JooS+MPg3Y3ud5cWQf+eMjv
Dd4RS7jpvMQj3vlMmMkbjG3SFUmltZP0B5qoeDf2rEpDBXeWM8I/qLLTU6jV1vGd
3jl8CoKO92QTp5sjIfepbz0MvSbGlcs8cnZJrMHDRqpSenA8GsFICzxLr0Vlofbw
+qwjqjeqfOHeZStlnMbkJIo10s8+P4UiVIhegbWFuWBb1BAecXb/NFvdUmK79gni
bd7mZhJEu0ff72vDfR+9I5dY1mzlcpm/S6tFMMTA0JaF5yIRgRWCd3CHi/Dk1e5f
qM5lnZi03513a8VuY9gbDdTt98EGBvwQhLxB9d8MGMqM6ZhjPG/K5s1s+5tQKqtk
7CzYkNu9+2hTeLt2bIpkx03l3l8zUQNGFJRbPwqNTNhYpnGJ74jH6sd3C+Yrgt8w
H/ZWFO5gl8Zd1JsOhUUFpQORZcma3rNnDpXfltldpwgtxhgrPwSAn6MYJhHO8K1+
QnVwYxHwYgC1VRAa3FWtUA3NWN9tJ8lpCV3ZNnQM01j58RzsntI04IdPn9nWYT7Z
CAsLi83C4jDgqZK1a6Mfi7Yx3xb5aSU4kDzFvcq9pp2rw5DOI7zrS1HXr+t2H8vJ
Ms1Swq91Rk5knNTkH0gWCAHIJlCLp6DeFPPLiXe9lRmRtVM5ieiaNA71fHX0cBx3
H/ianlWjd+wMPlCJQCaMk4sb8YzW+nhYlzc6/UBkVIMBubyaF63RcmE8FF6CMY2t
swguyb1yL4zyTG0CXCBafLJCxqHLzpiHDO38DryP30sh3a04fQVnSI1CApR7Y4Kv
e1uuGV5P4yqIIHX2IRso75nH+rCJah1CQnR8RKLe3SEQmr39uq3C5P+DUCw3iFro
vbEKfm5I3R+Y8nVjERqzicyvpU97QrW6GRtzXeBXnv2QkBOuhZV/KyuG7jSWHPpP
2T/ge5OeNoMu5kkFqepLVQEW6m4RsV+PyoE/GoitFII5+JJRXmbNNC453kWIp5B0
ypbeB2/HWEuOwAotvGq4J/KT2WZhTuOqV8tmDtAu1vBE37VH5Jfg/Awvb222HVI9
Mk7wk6irN/pHlakO4tAF1pgPwXSYwaAmLGFmmvS1aIXqTk+2fZpz8fdFkue+Xbmn
eNUIjp3HeEiZFZ79xe4B2fTfS5drEkyKjXB6C9FZ4cLoiUNjgKuuuSKEhJxLMpoW
p4+QACbqOZM+gfDOOhhOtUsoni3jJmgQN690cMutRbkwc8a7ID8in5vVgXh44/uH
zQxCuOhTwW9Ob1zgQq9VN14mu3fGzoCaVXU4KRtVZDrdrHZ4tp7ojHmzMxj2KsMk
zFkARYwSw+lkQVisNmR4GjoM3Z7UthGBSM8hIjkCle50P1d0CRScqSQ/a3Aba6Ea
J2vk0o/NlyhCyhtYitHpVnWk10LlhDwmsQwRIUc+v5net0Jn3p50fVqdqozEZl8J
PEzFGXlT1+ML/ty9KH9QUCz4QITUR9eaVpz+IwBamo99yoRIsVMq83SaP9XVU9Pu
2UwPsoVyPq3Kw40Gmw1mOAqc8drZaBF1kywZ2k+QzeID5zwVoTZGHr3zH0lmSxix
g9ycmqO4R3fmB0govbpNkUTh5srlj9RQ0VqRoPrPTpR88LidRD9PRTWg3ym+1ZA4
S/yRic7SX+1wDZca/V4nHTVD/JgEOoAzCVkQqNI9F2pHN8bs5X4Y/s5WtipS7x16
O9bnuOGF1IX+/XHS+WNNN02g/j/jFSGJA9TvuLPqFI6EM7CsZ4MfFbrGYtapdjht
gXKERi9hQeU7aAQsUXs1Nq1Fw9J43TePSIi9R1gn6b78YsWcakjfVy54DfftuQ+s
XcUwwQN0UzJGXG1MSZVXbyG7AUq8P86msMeVB8RgYI7mtBOApD3QZsvaQWa9w0Pu
JOiPKR13dO6uHc7+x0Cp4EjCmL8KTOTjrZwGfTnw/gNenI+yz1e1DPh8F9WIrxrz
UQOzwTTLXjSi2ykSIH/MKeizQ0qCouwGXETDV4NEVTt8zXSDRO6OcbHicHVYyNGY
Yjw6NjhfCBxfgRs3YY+0743XpTqANU1KeoibXU2Cyx9dnAglsOeF7b3fkM/DqQpV
JF0LCEGlhy+trJ3O5EHc9U+UnEfpEVeGM1/n8krLe9Kt6K2y4LHGnVnS96/p3pIp
WZ+XnYf7j0GXp3cEYpg5RSAGn3It0jb5RjdFlxTa9FE6JmHBTuqWhz8TD6t57Cex
PDCxr00vIvsDhVvf+uSkQWg503T966mOrMPrhxvcQU27k9syOdH2pAA/j/2/3g54
YGYWwj3HOUqZCxR/AXxJ2an8rdiulzKYRDHpzEN9PKTWDb0+8xQdyWe5Xbf8/8Wq
LqwICcEL1YcZmeZFPObvMvke8fAbpYsegBYeggIyDKW80vGVfJkRIgiu6zR0xu+d
tMVJ9qGOYGQV91+MpCDv1Qdqkm+6Mr2X6i4vEhgzEtc3MzDDPiwU6CzQ2popaFjZ
NUBCiT6xQvm1LJbgVqJeEeV56IMd+jUoWf8nE7idADpHRZ+V0igc8a6eD7W4Bwbv
HoyrOV2SdvCZr1XWq9E0uxiiCb8CBWmOGkFvbIliS/3xT2ngnrW77GSayDXn0ekw
Fmx0PLKhGehFjkTeYCCK7mX9jVw7eS/xWaL5Gfv1JQJXeRGRfcCXkTBMkNrSan/M
MT4pL6KJKXfqJTHxHgVUvGbOkk2kM/J8FHcyenND/mZxP/4FEjZoqn8JOQPubere
ZLg3NeXdOaWyLdQtD6k14aOYulDDoxHbNIMSXEdmDJbUUcaN5Pu8nHOPIhayo97W
5XrBhze9KOvEiLlIxlvqVJEAvOjQO1sGFD9MwGIVFKk9WwRDF7YrNDxHFGlWuMRo
Uv+sxfNLs4AkXD12g6ape9noJGrTXbNBa4ECob0UZNLMQ6H0X/hjtWcEq/YAo5st
/LTIuH2Iu65YzUTFDdbqsBMkel/lzI4GJ52rfgUzysND/IEkSxiXEhLuYDLEId+3
oBTv5VNc8+8w7vL62334EjDcpUkVFbtoveQQElmQw7LbitlnhUDwJCHuaDUiAiHF
beTlwEBJrSk5Nw1HkFm1peGD5doj2QawNbBdDXPDlUbyqFXDPwzL0wW32pqW7ERG
QD6p5sMwn71tlWOHSTOWmiyN5pN2iA2A0q1FYI9ufaiw8QDPmlHDV72ZgZ0mrHz+
QJ2Rvyqn9ZGLyzhzbYKMIvo7vYcI7iJSCVxthzSSWryBpfouvC6d5Qg+78NhXvsk
g0yK/r0sUpM2dtOmU6StrtMLe3bLBBDnTIGqwOvNy0gLaOE9xViZw3uXeAvHZ6om
ZdmCk2DAgTQbZNkIIPim/Lxy3bWAYT5MCyzEkFoPYcl9ylLDAXleEQlxRftL8ksl
dgVeGR8lQ/Wk4F75F/vBlaaDT5Y+HMS5bA+x4werXX1qnp3cYAd9a0TVUlXR8Yoj
72NzCwhJx66eBTJutdLO7YCfxEZc2qEtYoIbzLEQ/l6lhQ3wdss1M34P+6D1MjxW
ucz5EoYWqtbD9jt+CWn/+x2mfj0ApRDCubcm4Ro7b0FI9xngDNriqxMgsckRquT5
paS43mK2m4LuaihsIY9A7f3OkNa1+/DlJkNT/1Qo+Z7qpTcKnJBj3bO14k9SeOe9
GxZMb+qRVOsBVNQlL7Z3nwxr41ZpVwOeuoGhCuFoSlbIg7EWPK+pZfNW6z0zM4Uz
Yeh6DBwyL0YJnQgcMK5wSdPQEoAC6Gykfn3HnWj1N0zRwzAACfEK9RE5G+6KvdOT
a1Fud8d5kiEJu1AabUTrumtWvJtdcRqcYtKkiwiAKDp3EFFOQowwbcz5UfjL90wu
e+h4LQ9xyh//dtwaJDl5Ha56p4PJabuW0AyDx9F2p35PNFA7qpae3sTdPqHKBm3A
M3TA3JrPb8mgDnQQLyPdIm082Ue8Fk2xDhEhb1mDQYGrjjOJuK1SpHMLLvPn/CSk
Oq5MEzX+LlMeXlRsmCOMaBSj3zxd0oeWxVtlGTl3ctAeDTDMQC/ay4lBvZViB28g
35pWOUJ8brFwyd2cJm+VJ+SmmBBF34LIBdN56iMS65EI43XNzoBJ29Nz3Iiavq3d
D4mq2UNFbIssnx0pDeAn+5m+InehjcAH/gEeaeufgh//av2om0a9yEB7oPX+iE35
RbSMcdsgY7pRHCIvctTUFaoSZhHaznqKYN3N/zK+xrWpGewfUsqtfEv82J8R8QJm
se/yAXljf9dszWLbrX0OPbPJ+k2lNqaJclNijcr0K32OIrYZWLDldVzNHT3+ep1D
fB9qzqbLjMdWEUjXzUM3X9B+I5IS/wj0Z+0JRiFjVG42502h1/oHkVezj9pyxFBM
Gw3SSBnJM6p4pXJs8HkQNsjvu6jifk3s8uVDAveN4shi1iyCZA37An2ManTBvEhP
9vOhcNa90HkHXtU4dV3/5A0XBln2oOb09ToKohgC8mxSj6K+6u/PCB5DLMlhb2JN
j3jEOzuAyBm3dkm0LbCjLnlcZjNkBvWkIBzwNcFBS0Z3PbAcsEkyzLp3tk1qen8a
8vF4KmUSwPjZTnsxbE0X2XNywlDtFdgaupRXUfoiMzZ8cQ8bLJEh8ChgohTQcZUp
14EeHxbbfay8bcCkUxECZRkgrHzmedaNW8lTle9x+kEEK/IB79j7MJlqDKHAGVnW
mrCOeMylGvkv/XhdBlrtoXsz3+Q+LQWtRzYD1rQ1p3UWNxIjm6uhH+Y+l8t+3kOh
Sn3Q+6Tf4R5eC44nDRDiquWsVgbUkdsP32d2V7boKOkBy0KA/z+eSN9lDapQfauB
bho1DlYl0y86KjAGnFel+XQHfaXof5WrnPStuHxn6N72508xkeLipefBaE7fea2z
coIxbOLkJ+wS9ViI3/MSX6QjnfQGK3Pbl9sQ09Y7VyTdhdlgKKUl1uHxYKdkps66
3GVA0/9ORhKEtz/lJErNfCKO57dGgLbq+ApY7EvMyDTRTrjRCN2VPaj29UELRSCC
g+jeIMEXIjW7gACPybbduoSXfEBt1kKpwD+ZNqd+PyQyA+VNs/PBI5HLEb1ddTe/
WZcQPq1tFJkmg/daIwMnY+SWho4RAFnsooqgSn9SG3MluhzY5ZLb+B4aaDebwdqX
58ukvVI4AmZmudS8oiuoaX+Qsp11pT5x7YAo1WKkulxE02cztwdoYgGGZMTNDZku
wVo8Y8ejkFxoYttomve8eZu28/xODg9c3z+yqFvpblQHPAMiw/+QxIiPK2agwcku
Gyn5dpCJqIky3XbgBhISJGX0LCJ888OGvbxPHZuQaY4c+9dzBBhaKO1QLDu+FcDh
uLHWmcFEqazzflRx2dWOJ0edoNP8DsLsDqBUbmFQzmIAVMlzIM6lE06tAZFEJq4j
Wtsr6gcXVWqY6ALlQvlunE2u0SnmFQUuAOgIRLdYJFVygHLA+yulfXPdYFrd0LEu
OGyKeBUVK143HiF5JaedUbb5Le6MbJYWyPXa4GnGLD9yiMe2KpFnv7LKUzoSt35/
vs3QgLkJ87DKqRmn1Y3mCnEtxBGjfJIBvWWDkeRugUQGGMUUJdM7+dg3xn0QWvtU
+4doeILGeXgdg5y3axCV3aH+FL3RRxex3Upa4yXJU9kiEeh4HoJlJjwVtDRcIg0M
2TJIuWZy1mmNGc3vzdbtVArwQqMutxtGl3uDghOh9hproyYZYox9e/QFCJGLEptJ
4xYZCqWZF8rSU+xllcJqabXReqU+pYt98RLnjuNLyAoGPjCUkpK5CoTU24j5Qak/
ThfsJuBCYf1V/oaXj27H472gUjrvigrz88QFRssDWJ2LsTMddQ7hdAoQ7FnRLa1O
kDXU9Ke+B924T0WhrZQzIFQ/qafHKhP25nIKLAy+Hxk3WldFL38nYWljgeONbPJZ
OsXeKewQpM1q3z883Q6/mBeJYWi3Q9+CowwqhVDMEqX/+2zf9keUylGfyJITUXKW
fLo8YsNnMlJbs7MUbejav6H/q4m3zxquudAEfWlK2IKLH+mEl1/UeQsHN46n26wQ
/h0KPLQ4c0TqViGrev0xcr8k9wNaBRxg1suuRDhH0zI7kT10OdTaihCQ1ZTdpqTy
GBMjSUDEjjnVNL6nc02GZdUPbePJL6cGkQWO7LLbQobpa8ApWkkXMlkYT1El7mJF
WtA6mwQPCQx7ZC0dhbh/4iNxHql3nXOGxRAvKmPi/ZTJZmhgETv2nAi3C++JZkMo
y7qPYu1LsgmM8DGoPSNuYDlRQmeoujCiVjG4yL7uV4ZLIsulRsUHLWywaxe5qR2J
AjUvx9TOuVdlC2lPHNeaSNvmvIU/DAhQoogbnNsnOwS5UiwiGcYjheEz0ERKO9aj
cpGHZ8skx/iUx6jOCRk6wNxEfOxIWGk/k/jsbInetT9C7BuKXrTh+y5UuZOuwBSf
SfWkxP0YM4S5UjAsRsoYcuEhQ/QgPqm8KIrr4joSRf6fpOzZmMoDeQEx1nZCrubG
DAD6+l7IKSPrCeLLuDv+r7FYCeOfe3HneKyqZ8o7k333Avgx/57P5Q51S+QOAU3L
8k+QgBohC+m471w5xGf3pNNa6/uprQNEVWq+W8T1upgA1RSwj7+MFKXBMIvkAE7L
E4CV3B8hz+wi+X3bIg9WHvyAMyj3DG6fuz5lbf5u4f44VUTTtTyBDGPv5uN5HwJ2
CAolLzFoccCqHl2/xjEY1jO0PE9aczDgK+/MDSCnJs9Pam1cO07CoUCfOcQXCXd1
Spw5DOatqPr41rUQwtHQBQt1pWtCcNjcWAQjZfh9FPfPHt+dxegCAyVVKpwKLN/O
zC4MJ/JEhq1FS6mcyfDxK/Bzx1CZEapHbcQUrEmSKNpocNw61PoT2s9V8Lo4GdyE
8ERuOmsbBpF5U4rsfNkCRXN9/IoD7//Av0cjJ9ZvM2chbCKXvSjmDKCwjyAQgK8d
xU+MKz2oPqFNXio2DXmuQ7oAtv5YXFDXG5qNx2TG7nCrtI03wrpCJskokzmRorHL
uBJ+gBwkpEXNv+XaFzl15Uivi/5Yj55j/zyHrPT6kzi9rT/G9nzZzBuEHblX6IqK
5Dijb2sXkDNruSjEU4CotvKIoLsuoQ/OVT7XLcKZ7UlFb6n2hvwlhWuZhx01yOKY
EmCP5jhfqCh2L9LJ5gDmmaCXIAZsKKxro9fvIUytG+QgoQz118OH2Kq2CP7+RFxv
GDIbSLBRDRFVxvhSMfgnvaHa5sx6yndRoPU93YFI8AU32JS9SrV4W71PVvki4u81
umns/hN6gjWuuTKwVUgpq3T/ywKSm+DDJfqewLZc81RSY8a4mR9Vb8A8cfFEjav7
emDdXDhLJnLllc4WbfRob0QcX2IzCZ44Mjmu8qf1xrgivtbniR29B4rnDjGM4weX
JUeJlFB50bszV1olbhpJbjSvdhthPFtLc0ikteaguLNVFe+XGyDZm1ULDLh0VXSl
9Fi1z+DnA6etlfBx/6N9H3A5tiwzwgLsEpTSHDD+vW2lfFzGDNEYhqZIa8iXQU2Y
3wLo9yNCXF30892gtjS6ovzLCN5B8uiT8qHPeQBMnaXNgo3KSqPqQuNI/7PIoxG2
88fNHRyYhe5Vb6zFjRFOg3k3e/ZwXnSH0gsueqxLlXcKKD+0mqb2I/vmBsXsgoEI
L1GChzOEw1qlDG1RMnySr/cOx3nU0qkKlhqIoQdsh7XGxqGyw6Kyj+QlvBU9dOay
AreUz7jfsfW37ytDHlCGxpXvI74j87ItNecKdNXPn+xtWIoSv+jw2T9FfipNJ/Oz
hjEQzKBMdoB7riiQquaL+l73WEO7us41Ey2VvLA9DBvz1ffRAgMCCkU6NFl6U/vC
0s4EgrPfQeu1kAIrGMM4WCTEMqIp/YscjECMFI90Se6XdHpViMpJAm2NdVCsYckx
sBezD62XUYo3FGsd77dCB8qSBTrKqDtFvUuPiio0wY7V54p7T9fLUSO21k65qW7C
COsFSdfoqXRIPwVOMhFZkQtrB8JMcmk/4D11ubfWDtFohIzLVE4Kjap6LaudJz1A
+ABo+d9YfwfB7Zy2si1Wo+gNBnOgQchXY6E9y3oTG/w/CriEiMCBXdCRXla9am8k
TYKsD3OWDbrTlGGDIgkukkIuW92rmnE60pCDiQqCKXcMA49Q7D6Wtdt6gBmmzT0X
UwFnJQmdl9aP1pPiKrqlD9x4Ou0QdrxieSi65hunkKL6qASwGDvGRXlVZckZ7YNY
bAmcQ96DrRoPlwcsKK7aWKUneZwAHbqvRqnmrJPG7mCXB9ssloGFy3rrlD+B8B3/
8QE/7AA8ersnO//WxG1XHFrmDqp7Joh7MWDkw6pNec3IgorXedmSc+aT/blYMQRz
J0pOL5pM03ulnB4VaxrYqy8jo5DfKCoAnOd+GKilatcM96Xt71isX/DjOLmvkT9q
EI3/QXXwoRswOKwWyNVRXUiSqXx2NOH0BxHSmTi1LCzgO8ivc5VXHm6oVM57o6Zw
FIpMxKW5FQwtSEVESsvUm+VFLslX55rReasj4ODEsA2hHUPnuoUBy1ZBZI1McXuo
MidOg/tqS5hslj858PBW3yARdsv9IjhERxQ2qm8RebtTNoCxsu385+PAoEJbfgvR
SrwOQyXr8bT8ETHxvR5eQNsWSpq/Zbrp3fHMejLuLW0D66AxU9VJGaffa74n/8ps
xOUr/HEc2NsbY4aXJA+OzlFrjT9xzSpkrjidVt2f181kiFlSoY8UwISEKp0VzV6M
kdj77h99lcPKz4+Laa+c6gMW0KL7ZXOpvI+B6FPH8zUzASC3sKYTw55STSKWa3Kh
dl2r9ZdmTZmZdLOd+rvOWFI8SxeqPNWK8pUZz/nPe8YP65VppCBXL8ezZwY0LzNW
bQUWumAveL4ONLdGZfc5p8pOazSBPs12jeOYuiN8V/3LEUhX/+dcLczuAhLMC+IE
fdPRO3mNAyj8t3z4Pt6FCucGpqWWlTjVt689h8AN6gSoHpuR61TV22lybUa6kr8r
v+OGDKwZIEJ3AOCL8H9DpSJ6PT/1Dvh7djR7doIPNNWssULvkOgFBrAzfaUgKUPT
y/KhN5DYZg9a1jbjK/MHfrD35+SoffZO6srziKHzIFxiZ4Y14CCOuYsv48yBwfuU
iXx7U2NNAcrnY/SgaVxFWKp17CaGdtWKB2qY4nua/fQnW8ROWPSVl3d4Nqtw6mpZ
szJV3bufABp+GnY1ci6PaWVaBoU/IOJ3XGxP68347UxmkIF6pa11RteeoouI3XRg
xwkF29cEL22J6sROBvkrjYs+39gpyNEAlnMhyV5SH2Y4hIKQ8StLf2dHXuGUhaFn
CDoJsUjS60vrMPfJk3/H8v6ZgENi2ifUya/BKT9x6FIfFilOwtDohXqEZYtYPPAT
+7yBGaWaDKIcN8hE5cJsLa17cjAeiA+l4EBvcJavnkf12BS86Pf7Z+2AH14clzG4
xWMrVEoXI7FrOiCN1lK6BKNKvTdouAlYYJObPj/lpV9FDymipswXtA7hf4AIcHmt
jjzIwXLFRjqHAyYQk3Lbg1qcmACVIwD+5LCirUU1mk2U9jPUnovPqSppS0caS8mf
a1KGehTH6ObD3dBGDTPkZfsYV44UefrOgZ+33iR/EiE5ovzj8mMjDwde+uBAdjxq
/HBlRSV5aabrk5hNdY2pdHEyZ9sVfmlSvpCqnNheLXIsIyAo/ATfRoD46yjFvfns
BFEcoPQROfahQTxugFy040asmuzDI1Bq22IWoHSHyPVd8dQK7cCkBx8L9HR9VTzQ
8/dq4JQBLpG6ZyxOAw7qAALnjyW/XwFOBY7BC9EzKu63FeUdG6M+OyJA1ReT1b1B
y1g7FFktfPpqd8G5MZVOU702IbRZFUixFB1uwFaLyB+QJjaqQPegQqTKWIs0Bwlf
nUI8E+wRVvBc5l8Qbxkwd/Uqa6KgU+kSs8rlddww/wTJkACHrLB8EedI1qefM73r
RQyxE8AplpKh1TYkiz+95wwO0kwNTHAVwMX8WKsQAeZ+eutc5MIAiFKr7gZW7YQp
rpR8HbniojA688QIA0m76p1BG1W38pdv72yKPN24inTHrSZtNPpeww9zIxq1IkQB
wU18pWKxLNOWNMt9UDQpSG5uBEvdS8zaMxRvQz3qqhqoSEQlW9jDAqkW0TstzDQZ
sZcBLf/FjIkQ9Uuds90Hebv5aVNS8YjmRqSODMAt9NCDJB6a2muNeEy4E/J9ByG9
3XsKXnlOq6VOXrdMXaeDHbMpEwdGWkwL4qGdnZzuoEsOejUXCzAlvRfSO+ewWZC9
fX1D4mGZieVcmET2YjHv4MGdwB0EgkwZ3e8kv8eBE+6VdfU8BUBhrOQ+tU9LX6P+
5wTexQAK2Sw2no7isMNQrxmSFA1nfAFWgFXazoInGw05JtBJHl9Ot7KKXIHu3Ilq
YQPOLlEJdI6Hd1G7aX8m8c9yoGuzqJih9rXD2Ck3/rmXmFgzco5TaOzZPLtCgcw0
SjxAlo6xbhXztM6OOVUCBncqZ63OTdHF2CZRmGvBXOTuTecHGj8i53ComIrP9XPV
WJ20g601MVnfMGE9J2s81cAqLwnch0mrhRHHat1CS3GqyobNthsDhcH2NHWYt4Xn
TsZgZ2YydyNgwqgQNEH2I/C1Caf5sTo2p5oo3dWe4yqftSznYuCaJvQ36bAieSc4
Vw6qd3gbWFhQ83SS/IRzq6USeMLJ0XHhBlpkdkWnhpX6knyeSWuhU0qK9U8mVNG+
UVxeSPNGjlQYVvbN/y32r6cqFoNtrloFvOdbndummnPZ0ncEpbrUS1vpBtqFUzlJ
imnYOTMLnNBnZP5w2WOPp6eugIh7ReO8XGauWA6iIPdoHiHhhsMIFA4pHyx3rF03
uiOtmFBKJFQxpU+PDVroMLiDM2hZ0L1xtIsODLhsGZ8aphc78slCaGe7qIENHU2D
FC1Bj8IbAtC0TAaBtT5RohtTort7+/essAql9bb/rZAsHTfRGkOGxZni+KLyI+F7
walk+3O/hEev0O2D2kyR8vmvzUPZ2LPFF8IwKKvyTLadUt7S+vWjmn/XPrChDa2n
YP0SaCyspdA8K8he7ry3tvBvtbHutIoUKrDRBh8Uw/b4BDe26e5646PFK+/qZqXB
vq5m1RiYNN8NE28cJNDdjFQxtNZ99/5aW+hh/gfgm6cYKCH/r92hO0AGzxbGBdHN
krwfCTG4XgCT9hGa0ZM0lSbp5hRrIGGlJ6bzLmprtVYgQKCQ/jhiTiXuv2FWhyQE
0DJYhB6BInbVAuKFhpIKe1ejUYolcnwFVSxmgMz/1Uik89uDSE6VrJQn05/Bxy4D
/o+zfulk9Or83aMR3oGNtfuDWej7dACLtpw0mogxtqYuI57kC4iK+MuGIogVvxCK
4iF6nK+caWyGJeKaKGbh0eJUuAk08TIEX9EqYbW/paBTcI9Le3RV+9H+jsZLRfdd
zMh6PWUphoNi/V9kTcBsNkLaGpGN9nMdXgLquKA3PjqiVtxaPNcadWETDbIr05bH
Q1PLQ5dCUPj1y7GzxrwI6XWGEeqWx8TZhrmsXNEf/132DJiAvRN2G1DRQc1JahrJ
0hprHGCb4kawqS5WfrMZOcSxyn6aRrZZOZodPkssN3Hr70isGVqobPDkB+O7sSs+
TfsOFthUxGk591+axdv3+sfksFi4l+BNsnmfczVxcja9XD+c4XLWIgtk0gMfl5RC
CQoihPDTj9MTaWmohxAmSXHaF5iV0FwILRz3edoPNXHzkvt3KXCB9RO3KKyyKxU2
XTxweVNIUMUEqW/ghnrGNI07cXQ79mBC1CxOpczyvAnmLm8KonANEvohflR+vaY5
f+0cYCt1sxuECuCwY0m9YWwfGuXLQWZ4g/pw1dW1YsA/TeWG81mOSOQUS0I9sNcu
YpCYkNjTeA2dfAllEl2V925iz9tQ43JoINy5rWw2E+y4LNJQbi+rlGMCAu6jTkev
c6hGNvsYNHALDavWfhH2YRmchPylKfP4juc+uvcsXycQIxV2c/YoeI34tsyT9LkV
oifwb6lHRen/jAl5g92pf6Js2wEkzA7IMBVJNoWE7UHthmAvbFyzels2nwTywBCR
XDFcV0yMnSTY+FeLhY5V94ajqD/JivuH7dfBOZwjl2+sbV5l7wpgtlJF/lOqKmzJ
q1NT5zec4+N4l+2FL2jh6HdefTko4S0gx+4hBbEzoSeYh5JIX5/xI2+htW7urgHL
XDHgeWaDIu5y1ybiudcYhDV4FIsA6iegdoKV28HW1vCU6XkWMd/Wmx70p4EU+jrx
/5s3RwyWM8p9ivkecyACwCXNPezrkRzvNBcLromti/yy6hFZ+c4v4ljrG1Q86Bt3
Q+1mRcWBzHkk126sthp2xdcd/4yiAGLDmnrxgELcWEfqgfgKVWYdGufV6PzU2/+H
fKgbO6d6m6m4VOZjpNTtobd8rKKW/imvnT+PlQKcjhErCseNzxeRQJvgkzaDtBLY
yoVVv2FQGHKk/HCjAxCkZkAtnzGKqJa8g+sGdFxltZ4bN1yA5IcP1IOTsPxCiO+/
TwH7Zq/Y/t/X6Az5EBsIHEReRT2SyXr4Gx6wH/Fn5i3twDD8q6h23HOrg6lajBTH
w2biASx209NzpriPuyDwZ48k0UoM4TYAkQBLfGisfTVSDFIE0cvrBmaFPMg8mJdF
FGaBvM+LVNhkxeIuUitYO89Ja8TC4wThIe5Ii8Nq5oqjiJFRh+A8YpDtufpla+Q7
cgwE5gAy1+B8wexo0lbG3edJ/AF4ObD2+23yfkGPCPXmHE4+gilMyAC4NmYgzv9i
uX/M3rjwSS2uedp03P9fEW3w7FvnPD+SZcugOx2jpD4mSSZ0Z39+6jVwICWiMAOd
3g+b6doTLnUZyg/MiP/rJIIsLygnA+yHmG4udXcG1AcQpq7kJQcy1+cIIn7+0YGK
IAMuZS1hjoZtdcqUM1WehwOV5DkguStzMOcxNEuzyaQjHcbGEf6IQuamCW8q/ruS
+hpK0OemL4SfbvvMtWBNLWRg7BLGJlsbZuRYtGCxuk03bhuFuxM6C6+daXSvVhzG
kEs/WKkkDoAfa3GPu1yyN6Waij2hynYNR6envnSKpIZFVhTNOJBPGqeeqUeQ9YKy
5yOc4Sfx5F8qmWcZX2i5gKwJ43SD6TqRdKDomUQID4h3QyODX0wjwv/z0hTaPx/x
+G+oifd6pHZ2WJBBAKzFHFq49w4tiJDGOhmZHjGJUkSXZYkytjKkw3U0gt643egr
JH7PPO0cpJ34BEaOB4Nnt6aJv9AItatOjn/OsbyCg2xBlxCTw+jKGycNdvzz5Fp+
oi9voXqb8G/HFAdlFvtQcaX81P9zaG5nYa/w4GaxO5wfR6SsSvVAqiljPNTLMcrV
of527Pmapwmkh17S+RVRytJmjyeeXSWv+S6hU4goA2PIZt86OBShc/wxLXCzW0EE
kU8M96sV+C12iMyAldJYO3ailslg/puWMsdymnFQqUSe00V1qQQr3rHrDe1M/9hq
t3sYeuVDX7g6X4MUnL8QrRy1r/FFm3Y+VCkpqV8gbII7rnBFIVxEJ2kBD2pxtWXf
6Ub9a+Lfnd6d05wGRZNKxZyc99iAtVxMd1f4lN0UilYX94huoOH6NezGLT6lvd9i
SC+7Ju16i0/FCU9QYYVsZXxAgJMZ1UYAMOPDM3HH034aW0uAzbHdsChVcQqoFPXP
nVnzM9NpP2RWx0aEcEmlnURBthnOWJJsVU87dCL3EwKbf/HL2d2oabAWfaUW+vmz
m5B2QKBWrkUgQchD5FiiltUvvyubanGRI9Sv/DjXvWdpbCONSfGhHVjHXHQN0Qmw
nv2cu8O/cBSMKA7GLXhh0Mf2imvBB+aT31jiq7l+Kx/3d86YhWKoiecijWZJWzkr
pmLWPivIjRYxOWn1lQoCOEjyl4A8zGBINUIBwcnaIyRMRSaFMog8dwMpOtqnacis
wx2KheSYOOBEeyBVrJF5EaaHpl1iEEY0TBv+lwUwHjpQYKU/1biaW60aQrjCpnEp
1eancjWytO1NB1Ixrl8mSLl4PDxvr4dY1Z2FgefSrrU2ZllAZLION1vxSUeubVIC
dl4EQ/rKDHrJcvG26M+U1/hZ68zEGOu7kQNQu2D+vaVpBBEhc0o4xc1r3MCDGfvr
wGm/37nx7EFVREniZYNhO/qxY/KbI3uHI+m+Eewws6jS5Xjlj5ocBG87+rOIXzXK
u8RdYIYZOyW5uptxajgEslzqBI9pMZGoQWAjhvS3RayreZVvhUwA7y0hdPCVG9BR
hoQZeH4zjrt8BTTwGDh+QnIHN6jFs7XPGlzALKdqF8tolgOLtp+smlVP498euw/q
2XQppjUKl0tYePIg6zrikOFYQ1EjXCQmeQNZ++dI0tHiVgE/dHxGg/wPL/H5xqNQ
RadNyjdazbz0ISFUI4FX7Qi0eWrG7ue5O9BZl2uvqsZ7fJKewHWFTLmAzKx0U6xG
VP7iuszVc/kwiXozNpnbncH/PAqtFoa6YtnytOPZcdSlzWRtzI7FOhZvMpFxN/3W
ONuHpjMsgIrF7ykNJfDN5mITABYrJur0H4E+nNw8cpJzTG5LWa6xdD7kWs+6eX0j
gCNcZQ56IbQElTg76czL+hyrzaLw2fXWrPR9ng8h3iVfmoYxIznO6j+t72LPmrWo
4Th/VCPul4kdVp7kydmj4j5IQenpSVsCuGVaxI5fnWs/OlJnpSUU4Z26100qa3vy
9Mz53py8+GX6sMNkxYwqN9lOMjiBzwMrB7nsjyaEnw8eqqb49Gzccpv91Fyxjf40
5Tgtq2jAS2QPyFcdT8y0WsvIQjc6IyUAoUTEmb5UKS0EdztctIp/Tuv3zhLM2ul3
U0Ah9zT2ndhLvMoSahBkKUdFBd93nqsuRwhVUbWngqrUQB/HsXEVxDFNpeVXPsRZ
n4pUXyjh6pU/GTM8vbXQo26nxrZuTuwSR89XyknOxiwO82oL5CQmFrR+XVHz0di7
lblH5l/3XGQyl2iCxxzvYPiImeyvQQ1KCtKnwpi1y60fqZlNowPiXtM9m2Pg6Tlx
KWcSqQFLkfvn1qmN28oOpSWwupWVxMaufwR0UlFCb669LotnhhcFqIx1esYI/AP/
H/8yZxxYlCiAA33efGrzC9iFeJ0jUrn4rpnJceMZB4jwOOYkMQh0rcGtRn3V1H00
kcM8q21ebFR7rl274s/fem1aUVKo2SZ1ijsJOd53QgZpBwn612pYL1fX/Uuze49x
wxRLWIhhrdE9+gU2ym4KYTDaHdcjP903wewMG+hSQQSc/sEeTHJ9NBlyz59/nDgZ
SBLx8mCPY4w41IYvskaHM/QeLl5IpvGZKdWybcOb98jNs0AQT54zBWa9hSzFkc/q
ZZnXa30lUfy3MGtpPw2NajJ2PMY31wnCrEYZpj02wtcmPCxnJ5YIaLLIapL8MOBm
AeVPWRPWOVD2MYinlUne5PFEsmcHSaXl6t6J+TvCcmMieBYuG6SXJENmUJ1Pbf1y
mUEalUraI5bERxBzGeFTGwvHovE/caUJgVsqu4/IRJh+GF752kV1PXNBJHiYw9JO
zl93K0kbUSgnswagkKwiDKffUVyCWS30eotiwfeSIuMAKSIDenr9NIGlTAYIkhP3
hLJr3kXQdLMDiiX+49QCl3KSh6KPjXM8k1gh4F+ZUwHCnU8qRlEgB0mKGY19t4Aj
vDfusqQYY3liukW5723+kkG+6EywlyJKA+PEAQQx1BIrSJXoPSZs+/RJMLKia891
jKKZNz3HJrgVwqFL1GMSAyhtFAt0ZdbwaR5H29uLFTEX/PNxx89+QiCeKB1xgMyk
nogM09c0t/hBOOkGxHnmgEuSdBZLTbQGgdDf3Y7yx6SszwutKlpmXx/ctHc5wT0S
6EdXu+ytWE4rjZYCfO1GaLyMSQVoS3+uvlDCvnIvCoayNPWeDPySmc2lYGH8pIW0
ZIkhY48LPyFeKc0QIiV3eaPxV0Vxtv37I1GVg0VOL9J1KLWZ7nVJlonP12ZhdrzZ
pux5nW+etnlhJaMvLlfU3ubAko+SFwV9X7djAi7t7XL5zBSeQda3OlGs5vCK5tAH
LuUIoGHYv2Qb2FtXFJQqEvt49oxaneq3CwgCOCRhAc+2MwCO/NUJ9pOQ0mvlO79K
CYe9c4BhE45BeQJNaa3/pESTjkx+QBHJL1V9mG439Tu5z+Dlcf/WbcCQZ9ZmEOoj
1CvLnxsRjhH0ZASLFxUD3EcfjzyHrr6Q7hlnP9LOmlq4IWwU6OWsBoSX/K1E+E9P
K0oa6HtmXDJ+oDMHRTQ7N4OeUOQJwaXSKRQ2c7CDfIjQTC83zhYnE9TFXMKZNAjK
cW6q52buruV5Xf/XLxcwVoIWRAfLT/VpJQ13cDLxiFD+4Uz6hy49j3mPGn8RInXp
gJCeabswzHZTjhlpYp6EjfZh01hMOYyz/tzHCwNf+UnXeuBJu/sRzWv74GRCPSum
xNK+GEG4QK5HXPedDxwRQkWCYf90HmQ6/DkCAx+Oz1m+zpQMfov1FTVq0PIAy9+7
vwn+FH+H7w9I1GBWjkUBt0M6p8hROPjg6nfi2utGAgtbcAZrltje3Njl9+8Twq5d
72lD/5Ru8mORYlhyGVDQZ1OA3GhNlpgxeZySFZ9eDebigQNqgOyHZaNC0yzd8spC
tgQfczf/U2WcT+yR1/e3Ghirk2Ub/A79TGPHttikXdKENq35RdXfIZuiXr31zpRG
C3W5ICwsqWGzSYUajGFnTuYKCO+1M4APKB0YbA6ijNTStiYJMscgOuLd9HSKDAd5
Ka5WjW8FlZQmav2JtEruTMev6nl2s6Mg/OBwk9EhLicZKfyvF78PZ3litJGVEdKC
70mMQxzBqxs8iwv/fGRxv+VrZ3OZf6GAulWepJyc3VTDlAWSyKeEgB1AW/vLhjnn
AKGgpR1TSn5D21ucrJEdVoQbw4AAOVirJ8aAtAtL6Hbwa24fM/0om7sqWQfGSoNV
OVPtYb3bbe5skOOZVhGPw6++RXtwjzCEL2ZpMipm+t+0ijG0tQ0n87W/4eLufaIh
Zk4j2YX7/UQVUsWBqpi/QhNIs8rX5i5y/EQu9Oo7W1TJ9jegsLXq/U9o+AlQu5lN
PBGq4Mpg7+qN/Og0/Ace/G65uJpf5uzjTeaeAcWSrtP9Q3r3bywdSd5L5DcqLe13
mJLr54XHxhMpvbFMMYREAvJAnmBDHYdKw/LN8vZftEP5TWc8Acsle7A1l3mWnr/i
9P1PkYJRxWgyziZR+5dhsa7B1XtmO8UD2zOEuj7QOoLbElyWJEXD2uShh14BlQUb
tQmmj/cJLu+iojefSFwQ4CFSsTzG1+AlyliuP0WktJBRucfbDqlXBkzesmjITO2G
wkzRZR+HVVpNkXtQ/p8trMyyrKZES1jkdjH+AkbBWyDSmRXCX61znNUg1NpszwSz
CFY8xaL3oHx6JiHbDnR6G62PN42mWs8dUK6tFTVI1hdqbfHoVDvZSszC5UckAGw2
Ny4pdDRzN/Ubg8G4Ir0U24X5u+Rp94tl9Ren1w4gmizrcY3O4/FKA3fOtXgusEQC
zxcfP3uO2E4Tehmvn3Rhg3kO8E1A9YUB5NgssmSfgaTD2LzetgFhx1blKxNPIAZg
kZxQDq/vb9zXm5BIrdvV7iSiSxjvoPKT6RO7tAuUKa5bLayb68sfewN5AO1tp04j
gEH9WAo/uG4EA8st2MCUgap5dK8x6p9PvVCM7tsMS4RT7U5SVHnLOB6eSlmTNTkH
jbDuX+snhnal9OiPh9f2TjaeJHi3pqLKbvpW9dN2xI1wDXZkaRcwuWOFF5Sucpb+
fWulufpIxW5DBYLWWhv0ItymYxyUq95SdkVSAw59pSQfn9phXtpjmUH2/0u0kQmn
iOF8GRsGwNKjhb9LuPgY1UJjUHgRuusmrtyxr+gDXCs2BGnVzaEDLMDar0+MdSOj
sgZ6MtwwzWIo/noQusRqL4ylfV4P7a/teNiy0UjwAq8JnYgE5I1Mk3vL6GuZikNQ
/H0OIgKMUI1abV+5eZxCWy2+5NhzrOlMGUE3iOmElpEeTsPwwFjyYIIrgROJn/k2
GY9M1Oy3f71r7KhR80T+cgLZsCGwTrIAHDl6+L9TutDiDETSSqYLWJLng81pdTXx
4ntsCViPMZsdQuhNAZ6LC5o02jhp7twBXoJoNdnds5djEitmtu0yp+zVNSCuBoPb
955HTwEzLE3uFmIsbdBCxu17EiEpPR03gIKV9XVm4WGXA+ObNgqr5vvq25s2y+S+
vnEBDoW5Hog/FZo66Z0+WXw7HHsAMu8T4EQftgwN7XZZHkEaRirxy0UvA9+8D1dP
AJPPz33YeVlKOuH5F9G5MPS7foCaq0rlD9V3XUmXMTZ3q/RLajh1eDvya78dlyGd
zg3Onfd1Fp8ksB4VknbtN/3H8hanofYByVldHXPFXusxwDvu1/N5oXRPPBS67tMJ
UNKsWp2sKC9xXG908mnqAN75wbFGmhMOSCLf5Fi7lMUzZ285Tb3pW5Ew5D3wsVK/
Ypeo95taJJCLYgeRhoLCEs4XTmLA9S026td6tzny51s/4afE5o8RQYL/7Pj/jr0s
CRL58Gn1bwusaSrOZLxpfmVv9Xb25EIPQOoViPsj+j+cgM2kGvgeRCxmqoaETjyW
o+r7aq4bMfD8yLciFly4bMAAVZODOYPHcePOCjxs5X2RFbYnvdr+RnL8TknuRZ6J
SxvAJru1ndbmE865dvHkXilFVJ9TkXeezsdbxH1m7M4qFRi4ruzzahn8sOM+CHfO
cy2hN3nxsHQier7JixwHapQOcziFX78jfNnphdDhqmzs0SDnO+/utSS+lTcSi+2a
f7x94bxcVfP52Jz/l5jY3D33/BYpqlj4HSaGQVObsaOL8uuX/ShAeJMP17YHLqtW
IHlkUlDVMyq0D7LHLtrqrcbbmMXb4wKP78Z2EZrv8GpoDwWVc5/a2McduU+8CYUr
aHaav3GEld+dysy99n9dBss3DEnWkzUhRWaYmmIM8UQZgAbW6SQNgBY5OXjtM3nw
SgdyoDDm2WT99QDEEg3FmXFVTx5+KAVIkqLEFp6K6uDwiy9no186+T1os+vSNOdN
PVJH8L29eqckP9//Y51vgJXHYIci5UzropFgoIVi3boi6sKsEojxrcbnBHsFml3s
tg5kXqQZwe+q6FozhW26YqlyUeOEcoURlzeWvbFOziv02p+UOom2L3XbOXbTVfW8
E2WlsnVTk0PE6qhxmfG69m6b7konKRwBigG5YNWyxYhZkmVdehivXVWdbMY0Ed9f
7B1nW43DpFrLq08d77jhWlUZy7T0H0Yw8NgUofF5Tykpi4na5Iqc6zM18yu61nPq
5fgZMpJqY44LMMkR6SO8pMxtdzjwh1nZUGqsFJZssbgvI/z5nIonEkMW6x6NfLXx
AX6RiVZKELmlylzK+W/5q4bMX8R8ssTSYrprsDOObqWye3YXvDeZX7DC8n9QjUtB
q4YiBQn009PG4FTQMZ7ul81YhKsRflPN7qX7WE8QI7GimJoHzfoEErEsSm7/a9W5
J72Uw/m6AzV8PZstJF9TFHpQtKmx/ZJJvlz1rzVTrSh21fgmZ002eKluvmNQuoSK
Awm1yD2lvWfdJU2BFpuoPs0EZzh+GHExBriPldoFlLMsKzRrBLp/tSlUBJtW/83J
DZCBRZ1K6xhCsNkabU4QcG3RjtXfqI1M6IkkUxM89s6jvbD4cwNryXlY6SZmrZ0g
7tokpuQ1EEv2v0/LjrJyCeBb30FkcCqhPs9kD5lOjvMLMAK9Dh0unVAFyIutzW/4
aLU8177IxZ/5coUdg86KoXxhlus2bX5qT3rOXu9CJS143nXe+Mdi3S+uPwb4Z/zy
1JNmSESEW8ORP6ESeFk96SRA3EO+OzORDZeVWfIRnGis2+gpJI7Nw/ouPMwzHK1X
vIhjcn8qstTq/w4ZRlBs0QBg6qJzvXvYAUi26fp4MLzgCphM+yYMEtW7Hcf9++lI
aizEueiZSwJpMCeSqzW3qvgcHfqVGKfSt2F30eORSqzwB6wZoV0EG0dPOMzAF/cM
5SSOzqpdWqVCJGCsmERpl1aJjLgng7rkG6W6IoPeOEbXNzQrQ3srjbnu93yyZI/w
MVyPiTyOPny6uj57Oawh+nIMXvG1vHi9+3pv6kLaPEzn4dw+Q1LchPMOWSWa9Eci
KRQ5kYmeiHZHocxXgwFZLSny4hFvNbE/ytIVfslcTZo2i0+URWoeL1JA9eG+yLHg
EWEulOUr31mgCAUDv9ItnlyqBXOyHDkHbQ/uGaZaKdCyVnsLFIiBnVIfgtm8sXdo
ZSqnLbBNV3L9G5Wes5TbHIT+JY5xxOOFal0slnvfnXxWUJWXNRZJ+0gTTe2TkeuJ
tfqB+tPSr5r8DGHgjfbVH3fBYde3OmlyogMRj/jdlXjHQLlWozIKZR2PdLkV+qmY
5I+xnDVYMe7jEjlU275VhnapVnp5muZ/Jtz3PefTYwA6iCniWWpzMLajVpy23Nm+
Ly8ZyhFth3sxsYOLH796osVbQGL2cPZNxe5VzJJqwN9jn8sWVly1V88d2L+HbWvV
busPeOyEY/8RJglDsK+y0vXhvQdo8ZEZ7qEWxNEc4zhxfx0YvAWUFVKI08Pf4YdO
EE+IxwbpjhWgwWyE/19Y56H2VRVMnysr1SitsvfqZpj4AWOQJ3kQ09Ux46/m4axS
LcI4SWZxS0sbtD5e4feWMPwGwp3qfRrUoELdykXbjNeco2bDOEEWpgVyU/Ulc5ou
0zodVl+DH6HD6Cgq5jr1+hS5XUihWPrwTrDimR3AJcvtTkhdUux/vLeqwDWD4P8d
yc27a7fxns9YaGNcJrX1tbUf5KwUwdIZa9rJusdqz6wzCbL0+1Pmd1AdkbQfM1Bl
VJvA3sE7kOXSl2ZFvJ3QmRC/rIjfEkZfOmyUGDGp6kQ7F5DVoArsig66M6qsCS9N
haZvtj4NCMDOQ2zK0ynfjT8NGFdTTnCbqXxIg4AsJ+XCVLDCjgESi3KEmqYPjcmt
sR+4eG7itUfSXqawqtLcoK0PrJ7N0ePGd4CYLdv7gV0XhSULb3dwvsbAS580Tii6
Bs0dVm/oHpdexgBMn3KYVRZ8Q+YZYXibWwQltnusLoOW9Gzo1tbXE4heFg1wApiI
KTZi7iweHJkfKRQu81cykEXERi6sSqgZp33xMGUBdq06dY60SSUD2aUjjl97wuoH
YW9vpjYM4XMQ5pOdQU/vw4y0GanftFQmdxaqiKFwkjc3Sa+BLYisYZuw7uaPfodO
280hSAdVyinGIbbfOSqOLdEC1q/xgFT2HdV6kT5OZuwLBrLHIDp0zcv1cAwwLDlM
I1fLjrbdIpNx32+zBidB1QLmPvxsKf3CTkkTaOHnGF7CTtm3p3gmQ6Rag3SwRDNk
NrjOI64OFvT1fhnxtUB8VUnnae+u5MGDJSSg8USbTRYmE04Wr+mu90zO4Bf3drkh
wCIUOS6jEURlZeu0cwUhBhSTjNM0TmZh17cd3nRZfnh7/jRgt23WmlBpmT9AFCXx
EIItz7YL7dZpOTg2/EVGhE0TuWjoIaDYjlw2XrjdbDhfCLC2VuARwsG68GMsxdgq
KHYBCIplN8c6H+wmvwRM7h1ebzKwTvFcnkVeMVigi5Mxd5cLK5F/fWBPAdZN77II
F4AL+4rU67Q5oDcLEPgNyv57sofhGWDr3hWAbv7PLOAw8MUOyJ3xjoYf2lmgERmr
SOkJjNYDDkximX0W7NRM06wwqD/CKhuv1sIYfbXd1800tqzcJesaXfxzYY9e6xyV
sCyxcX5J7E980ZFzcl65ERI+WHPa3lTobpWBay/J1L3Pp6UxLJnCIgXfMKV1+8qr
x+Mwvzz74a49rUS1lvUGolBMuT0z9taXbqTgVutl5vMM0Sg5gNWwMnHb8Ei2oyiN
cc0HLJwsRLkYnhIw4OwDaYg3yGIu5qNnNohft+V/CDEGuwJ9ai4UqM3AllMX7Nyp
NQeGB4TzQP/DueKNJMKXwJLHfhZVjCMaW6uA04mZjnIaNsXzUS2kyXw7r59wmNn5
/4GLjNXevJ2mQAbk0uhUKrS++Nc1dlspQRsKde8nY7ANfrHaw/Cq8DRfmBlh9OMX
AL36Vuzg1V5zfwBGXw+IsJ1vZBAFGEkYML+8QyNTf3XL7Uv8vZeo0sakpag7V3e0
CzNOIjF+9d1TF05atzZAIRrHB7KoQosAqpiazylUsGOJP9y4+xmmU6xPPZer3HtB
wM6ts1VFvSXaCZh1Q2/z5eMXZrvABk6kgqOL7b0FVOAknmCL4UcQ/A4f72cOouj7
nKODNlRDH6Mjov25SrVDP5a+YZwaU07hCV+fy7C5MYCX+4Xd9oEj1NwAIGZ//W5k
393UoI3G5ppdL1JGaUq7OLQXzAg+7DwrP3EEQwXWFUuKqIYKHHjoeRcXaBpxpNPJ
OWBfGOh2AJ2TBn3iac5fERmqZEnOeKw8HzKmIK8RG46c3JC70j6+sx0P0GCkdGsF
zw62E15fWACAX/hKdhxPvkvZ9ye508GJrVzAnDOxDqLuAGGsy4k0zOtkQIO6XLms
sCKEBgnU3opgM3jypDecRDif7oLKb6AIMszTQIXnWsYZ9w7NGcd/qA8F/7JYoXwQ
BG53KjzEnxrdOZGMF2UkENzZcPf5BeCmRMWb0U8BFvWhIelPGM0BXOm+6l2hgn80
llSumYw151B+5aLTnAdpZHc2FaCHVkKGca/qtI2R0fqagnMpgFUPyyNr4pzWSsID
83mN4MP0hEFlf/zkDIWJVcu+G0p0dSvZYuIIJDUArOEBmp6NanozY5iOyMN9zmTa
okpg2nXf6qFiI/25usH65qWmlhDzXCJTGemnEuMDKLOh/gm2EUpqsrSsmjKP+PNM
w0T46xCi5gJziTEgyqOl/ihEk/6H/3YmqnFy0cMZKXK5KW/Adfih/ZKOIYETeJWA
Mt/UESpGp8nWLskg//pVuMPF9vPTUWoalV+B51zqyMgx9Msc06wBNRoCXaygZ1kz
E25e9LEz9V3pGTz1SIC28DuFNAwe1Rt+pQCfuh89eO9fRGK6cdGBQRyTc5GMOgKf
ixyVkxrO4CPvPqLHSyg31qFIE3VXVUPMATdyAH66xjhku2oNoDLZO1BPSqSyOr8E
pZPNeRsKBT7R4/pIh8HaL4uUjwWH07SB6i+mkE+8mk2d4b6Zn9dwoOn4IIQAwiLp
/pbq6RbYwQQlHgVH9/Pw8TXWkY9oXLKoLQhYIQX6QQOn/2AesOHT0O2BnZxtxSCU
X4shOCqkIxB+eALk6cwLzfD8mmhjthENPXk9tJD6Nd5GXruqRZYFYABkyQr0Jylt
N1ZPyVJLHxn2odxxeb7Ox2molq1UR+WgdChAAnE7ANjo7z5hIdIGDp92SVP/xGxB
pOACvAIfqD+hhS71i9DtkLsG988F86WK0f9IMIb106fz/SzJgKuxv8C1YKtwyRLI
9HrbPyvxAmdQ1250Ne2iJspa+lEF/xLhmPoh6GcURvG8kQO3rffcMixCmnlF8tFN
mIFY7mJZgG+E4I3jERdGgBZoR2qeHiALKKrbMDLp1MdAAHa3eAb2f2bwXb6bvKKH
NPJpDkw1lPYQmGwWPEQFNSDvSgl4BzRxbCeTzOb/N6GYLu1XMf3eBdGBEZShSdV1
Uv38bduNwkCjEdUFSbi81MmTJTAvIfQrY2mmEUkAf84H49xkLHjs7eEhdpxY5pXt
zoPjpsVuEEYOoUJhKRgcbNexnANCwP3uZ5ExoC7e8VJvs4ojC1VR01taZmojIPBI
/0IKEdqECJr8dXal5jyZdvUMim561H1O5dOrtDOQKakIEkqwwQ+r4WbUkWRuzVvp
c1hKx+0OnnaMMEnNlF9TspWvVvbgQ5in7k+NY40SNtCv8ey62AUyQG59GpeIBcA7
DIonImI8/x1SgEu3yl0fglJ4E2jTGA3A7ccnRfESi/w4D7mMa/M0Tf5HKDS9/j1w
I9ZTJwsSyg8XpfXYYMwzHoSN3ZhKeyOXnYmE4Ydf5h483Jcq/9SjCCZLCHI4psp4
FtiWXTB/Zb00J6C5vWCCuklBEf1VOlctp7Q7t8kZpoO3kB8WOXrfJAu4dxR0Ceb0
sBeiAL1GMYVEcReC6JwLDpVFrkbnK7AoIP1bdHjmX1dd0QMgNBdqB2MqyHyH18m2
vSNVmqdH/ZhyJwZrojybTWS512IuVro0tz6jdJwb8tiaLHS8cz6490252i8Q6WUj
ZJtBUjzBDFSgxqPBhAE8e1UbOXw0OO9h873rQEfcfeT1ISDVYY9uUVaZGO1X9P/O
aJDmIbx5FLdYiuTfLGfoJH0SrZxEPxS2/R91rRKfAZziKUf6XQdQWLImBBOGzV+R
J22f5NPkh5CupNceiW0JLogcicZt/jeueXk/3u8jK2Gnt8zR7nrP3hkHElUTpVGH
mPI01M6ElyFRhUJIEGJ76RXd1cPWnFIp46BOcm9DpRiJJXPoqZ2bNps3GYvniMoI
37soRKgkmgA0bp6Fq4TKFm4O3PvYlN8LwwevLHgJ9ZvMU+Mh6zbdOVfHtdNiyhGG
Zh9EpIi8MZg6RaOStxdgD4R4QUF//w55YqmPdXX3S0t6OVH+hQf+VSu3Anv4FU6V
DRXZDb90eLfX+a8IRU2gWAJ1xeKNLie5gYhpkIwSvvuJI7HtPNYfeqf1CV/Injkk
il+rY+ANkkCd5Y7IbfFMzLYeFeMBBWEJVUbm1UgXAljCk7i8/2q2tpe9rnrY/PEo
hVDlnsE4sEaQS+1FH3UdSPmMrNuFyBekrAuKmPB8i1UebG/nystz7ZDj4RZg/wik
Xu51yIMg2QwfKQGMyGA6+A/x/sw5l/nT25FtZvN6PEXzqYDWUUESDdQB6IEZSfQR
XOizeSnTSkYEMeEvyhSGCJrFDbvP/7cJJMx7XBh5SiFwjXsmlTm5/tL5iARzkD0g
5pJ57zntU54DHnYPEXv2y033OjwG8eE2xZ0+H/keS9KyPZmJJ1b781xs2duoROHi
xRtIuznHNPGZh/ZR2QE2HV6Wygykc7ai4WuqAsUvW0Ks7XlNOpHgKdUFln2t4U8q
B01qurepg9Bsjq1/VJVJ6WLsqE5iDAecsobzpObL1QNFt/lE4oXZvsndU8fg2Hg+
z9Os5vUsgErEfEM51fZgYNAZs8x9gT8YD5hcNv8IvlCe2UhHyCpdxd2YSuOsRb5R
kX5+HahB6ouLQgZgSvA8nXgcOCv6TJrwC187M48eG8tv+S3hU/mWjSi2ltRubkNt
wZiY9qOHeHNtgX/mtadAUWN1QwPH49yCrFhHkRt52KkJD8yRhR3WwNG3PR3zFmB8
fuKHZyl4ybX0Tu1F4lOpqYz2ENGYIbwa3HpvFjc3JnlZ3tYGWWlHfD110yytUyag
WMN9wlO8o69eR45fSEj+RP6gM3zJcBZ5iPY0K8D+zhX5HHhNhJN6hMjJhMbncdYQ
mIGC503jWQ8bZ/0kd4/ct5QNXyNvvEdqU6SKhL0kItDO8Ao+OEs5BpW8izySIWAr
h7Txxqh6DSEQpDXsUo4Scx4tC2QiRk4ozrewhVFjm71C2o9pS87FIeV9Yg2OHKnQ
BFOziFXaLEk34rrFJTm438c+HRYSiZolO3u2ZMZPF6tVyE6mAZmNbFTSTn95BzFR
tfe1ycBcoMYs3COp1+bt9VerHbiZ/g8BBRruvckR0jCwlpkmb1wv1ygh3gmIwDu7
cNcZnfDlSJTn8s9VVRS8hXKyWqjbepinsDITJBwv1nQ+gMxwcyimgOtKm3ZyNSDq
TBIFRkU6dU+QI7SsSYexRapT4LegQg79A3OwAFMXXqBX12ggqefjUcz1mmU3aeNI
67DlJ1ZtbEaJCaffvLdeBE/9CgRO2Radyv7gOpBKq+G0KEVQt+XLuMYqqFBU5gRU
zLP7ID93MoLbuDImjX/f8BmYW+JZJrVymW9Q8J24mxC9DsIS5KtTBzyTt3Exf2ts
44iNx9ttu/1+aXGjeC/YohS8p/mFO4flBcKAzabM6TDMEEUAtZVg/iVmAJwk7iXh
oUBEZ9MFSyEoftOa8EyqCTiiaDVhbIf1027rpiuzBpINDLyioZcjh0KjC6m3DoKU
E1mxDROLW6JhyDaHj3a11pstiXMb7dbqDBrtbAgzKc9FBdld02WXOkK7lQuuyUFA
GbMM1eTmb0KljLyyP6g6lhqucdm7V1lsjo8k3MDemCerGU271/xP7WVNTt39MYoy
aTw6HW/FJp5nrDQsqmT8KH+zZxwcDSDBnfoSTKYWhzL1wu2n8Sbgt5imovB0AJhQ
Lrp5Jjslvrkkb2xrmSDHNP5Cj6kooAx1MmOctMgrYkPmUesk0pERy7L7Sjyd2FB+
aqlk1/NgNLmQBAoQ4fzc6YtmafnHHNB59V5tDMfqe8Q6ZhDNjAhe3eke6oV914wt
gkUmh3RCrdz7eqMfKdrbP51GBsafgcjP03novuhLwZmM9ZkZL2HsRof7jlxBrmF3
sGDemEdnktx00x2IOEFWonxn2KzEQBVDqLGNKiJvicx24eISCsJLn9vM545e/J43
UUvMyhn4vAMRz1cmBgqi+OCJhfCcGYlwPavUh5kWqMf83/3nw1MZKXzcV1Ovlg2F
UX7vmJ66eSTkKdfxjVHTTyrvME3QA55qmiKNQJpazm+gkJcJQp1wq/pxuOVCCpvk
dZcZbd6bpTcYX4ANtR9cW17Z7+zcNhyAsXfVZH+1IJelyHGe4xwsFNbPqbMhuBPN
/ifdtaGjvZ/KggQchFO63vhD7gCC4ugVEF6mvyNquLndh2xHPDio8H8wE31NEyl7
6ijOBtdd6RV9YWkiu3MmNhP/LVj0j2LIx2g32foBlgTRMobvXZukba5rOY0dWFFd
az0eQEgGr7tSK/4CaFcTX4LHW0pMaRDK2q3Uzq2yY9gkBD9RMqwgCT8HlEz1xkfE
EM1qwVUIt5cXqmZMQvZAE+N4imbri1+mZAzUfvF9flh+bri54xbEodMlnVHPQrdC
CR6htRjuay14EIjzHrs8hyKL5CBhSGzMDfdAhl+/AiZ5DZCSCakhNMxQPAK55IQV
458RZlB2pd5REYv3tvAJhJQaj+zaiBRD+GyudochV1GMv43mI/2AfBO/suOWrWto
En3GBr1bm9AGCeFHGLE354Hypvdy3D+oZSe8uTcaDUovwJ0NiR5pfDhY6NOF2Z2A
mnlq7AWBhSduVE8X0luwTFcThnnwJo/uA35civbS3YoC4JgZdAgycXuNOflLitWm
fu/ujaaK3QsCu4EUSSbjqMJXhcPcK07J4kq0AoI6d5REMIGXFFtXmPvL6a2x2TLW
uZbZ9RFUAmDH977mFy0qhyHshIJikb8l97i+Pg6Cd4hKJF1f8yeZY3we80pIxBHt
/+EjiMZ0MZMSBpJUb98LE2Qg9WlGXyaZ4YrTL/Pi9Mand9aOj4jceiwpYY+lTCFJ
/UUzrqLeTonL+nMGRIydXgv7t4LF0nHWBZ9Cac9sVhmF1fQP5wz9NMX6w/0JfNqE
6sO81qklmuam/0juuU6T4R63Mf7x4N7XWzavmRHuaiF8N3BBZS9UoAdDvCoOl2O9
GeMBRKr0fRsNwkt5YsAjOj04lpbtUE8tzFnocAi6F7jHIB3JqIM695X6UmGSSK3E
WIYkWv9DdOzg49qdQ+7IeUUctLjYwZ+u0gMp66CsQieRn9yq7Rzdca7178Bqq4ON
J1SPb6MTu0lhUkyrUr4vbmy5Tqpohj1C8iMrV9TDPWE05wE1VPuW7cv659nJRJPf
iJG6NCR9Rf9CJWoCrtpSsoDc5HGXzXqVcSCGNJEgJHOzYb3Y+x9UGKvjGu9I32wa
YTvPHfJXK3H4xMgSh8cmsniPkERoIQpJV7FAvuL5SzQrMp/Djf/LVhDCiAIKjqSX
bg19OP2+G+vrFomVxPlyn6RB/NYJgTmuGm+j7VAj8cc+lNEqRFwjsBwx/d7gXu4W
fVVxz+0lFOJszk969kku/qMg/b4Drw/h4GWpxDJcpcYCLeyn8y+eZK1UApU3/mOs
pTwsGB7qgiAvhdOFT2qSGX0Kmln0GYf2OuleYwDScJ9c8mDNCPfOT/IuBJgfY5dB
+MgneuhRMkjyt1GRXHV235czsWaaUWhbHNdfFGVJoEQ30n/XtDFknNkOnbNN4FcP
B1QiJeZlMeQKuLFOLaAhkgFZ+KnHPHjcJzdvlQJbK5dLQrSGR2Y/c7hOjRKZ4TVZ
W6iGKzKCr2txdGVmjjrVLChZsO9Cob+TMh8M4PE98CO2gv+q9CdS4u1tyvAoMB+s
E5VyLJ9igaJYDaTnrDM0dTjp2lxpBnr6p3JlnyzRkfkJddxujeUyZDyu0Wf7Ro8M
lwWLtZbT13PzpNV7c7MlJnK3WDUPW5KLiyeZK+3unlM2ZnX1leoFFB/EW7NB2kd9
ormLefiQoC9XWB7qnY2x03AhPXLeoowvWPiKOUtfAZ2RdxyfjK1szlJRFrCGgFN/
GAQpB7OVAVbjjVQW98m62c+mWbikgQzvEGtfHk2j8CGPx4c3b1q5eNBy2Fo2DWBf
bgt1W8rqbfyoHsLrCwBj+bU3ZrTI+DBkIyQaBR/Y4O/lIwmgze9zXUoVwj3gWApD
XIOC1UNF73af3YRA22YLRfvX35y55DliEPtI4lbXrYgvUKJ+PEActtkZ+65Ok5co
8VZUvXpSnOftBELYCV5k6erZd6zi7D3alEzRwVIr4IihYV2sGwC0RNQHb2UD7ZKp
Mu8gWvfF8XuMxFfUWVGJlB/fnh90DqxLpcFjjjptKy5DfnlJ+ytnWuCcCZq2+Jfk
jIZbvAcAVKDCEFUUn6fzxkeMGHiLMtYhFw5E4urmYY4pAtvi5H3cwN1hcYVTpn68
KbZ9pZqT/V4CeU+bPRfD6VRNjz0Ej3KX5aM+/OdYBftJ1DCpER689dyq4tWZoEuz
LROkr2vTMKQbdpTSuIHtlKXkb9uJ9kLVFCgbJWsx2CAtLqt6IjeObz+ZOhvq1PYX
UsAyrsAVNk70i+nL5Q8n6S3+6eoU4Ogh9dZH++fciHzP/hg2aoV+OcErvyJq6L2x
O6pQjqrPw+yrbux4bmsm8naMK4SaameZyIrDckc8dttJ/4F4JfkmjmbxDCfa4h7U
02SDafwGyAwIW3wqyaEjRKoyydDCGrXlY3QWb5iBb/lHEkGwQRIf5JUhrHZlKBI/
xSCMoI8deYokKirzukrVx+9nMCYMpP6YGWTEIIKULlF7Jd7uJlZEVJpMmox7C3DG
BJCTq/E/2lfgVCt+peT4fKLhFExZHYae+Rj6lYexGxXjkMHuYGeKr77wHRJ87rFt
AUeQSbGEobWJ8By1XX1aQsgv4Pn8V1VmA7tGYtIvLtNfXkPWvRm5ShMwDHHxrUhY
UdULG5zAm89qugPu5Q00Zoi4zqyCyGFU3eqh0IxO1Br21OfVJovTH2wYlr9izDlq
qvu9umsZsnybemEs/Dyxy4uL1/64oWkTTef0317KcLawEKP1hhc0LxQn5m9Tdgo9
WEmBDxog8+JGl4ZjvK1J9b79RdwGLKlfpMwijz7uH3b/+ToY8tKo9AdxIBUBeATE
iGA7bn29OuZ1rMqhedfFJNnsznDNhQ5imPlkyonyomkYEVzQQKrXLN7zAlJB9vjb
6PiSpX46+dOOz7GoR2vreh6dw/nE06Wm+yMIqYhM/C/u3XMUKoi92wzTzhkmigHW
U8J05J1M56DxDXQdaQTC3UWt/XtW6v7mOJH3RNVSke81A/OnhOmCQ4Sd9aA6xIVt
HnglKNI8JNTRjAghJ5mbH6Qjg5eRgNAdL640tCEPFUKIYbAhlpazvhuI8HO0BWWN
G/ZKVbneGDfaBbPcBXcAQ5EbEy++GADIomfpPldtPWDmgnECP0NFc1wNWnMdscEO
y9eiSCRMS4Ks/XiwqElrGpOlaUBV1L+8tSBFInTXlnY3/qsEHfILr9Ha9uuFZpws
z9xsz9ea2O5Qyo1Z+8bKZ5Pk1OJbRRD9IkRQzk/YM7dD09S6hLaJXXkJ6SeDTkHd
HrfrRmQWszR3XdcXvgvSgkvC7LYpnaU5APr7HY2JJZP3o7cAdPkXgD1JGJWI0W6f
leS4J2upLN+X/3U5QMv9Hho1shI1L845HQ5l/uHKUXsrtPQpasQxnDucj8aK9eC5
ww1QCssvYBHVH6vzSJDA8/S0Mzj6UB54Em83+Nup8jVuOoreKEYyJcX+ggdrBKNs
1nTnQxcQJaQATPgDYhD326WStTxeAy/u6oejPVICs7doTn/wXWmcfGp5zbjREIZG
VN2kfgqmk5sKapGnEZWSnPnbGEAcWMC3XqMqyFX8tpdiUAwji0ZR7bXks58nlp75
S7Uf8wSJ6+kmqQo3W6oKrg2JYKH8XliFY0ItnSs1PWMYo1UFl+Bl02dPNkb2BKUZ
XEbRNZvrAuNXcDU/fqtwWe/3zIwspQZe/9/NjJEesnW62MVz6Af74azujugnjhMH
oGCyxI1tZovJTUlRAdAwtYXQEJhOFvcHh1tNtELLIMA33bohBdN9GWOmUtViLdBa
foIdVG4J05JS8YhpGkGTyDcQV+GvtULe2GeB2SB5Q85OIYq7FRIC7eHyNO/bR4l4
75WScqOfZHm8x5JzzpbsQ9F6y3Y+6j1DZKB3sDlDgvnSulm01kUj7KsD4rPFLRTK
UvyPIWogKyyVyeqVna9NOAH/Lf/1A96wQFeMTEiec+7GqO+7HAGHoRXAIMzwY0sQ
IcwBTpPWx3ltdWIocAloVvYD67UinDKMhi74g+ABBWKm3l9ovd/BaNjxVoKL0vCp
Jm+f0AaJFjO8sxivxMnZhUds9WI3LIZcVaBHEB4JA8Dh3lp7cNRI90AsrfbOEc0B
/fu0FXtClYAAWckRnl87XGN5F65ZJCwguJpICR+FftLrprqB22ZQzFAVU8Cj9Kry
y3ybcevji15t+OGFFchMtO4kM24mJtFrwgkTvMOsrdWQw/q7jTc9IgtxERGC7IQr
N+pNVmKWhyHBSTkkzsxxzU5ix6r0T8sFB2xzPGqvn+O35sN1eAeAqvsZEciSJG1l
lZmBjmupnWRH5rYmisfhnJiHiRl7vJ526xW6pNYWOu1kf1UXUGMLMnlQY03AVFK7
Mb3CjZFBTwaFuaCfyV3bZC7CqRog/iJJiRyG6epub1Xl4Jdn4q6RJyiyTCwOVoeD
RmAgSmXYNWRrRtTAYYV9pfWlop1wOBPApTg+Nl3uKzrNF6ILxcrh6axGcP6Zucth
5U0uQsp0A2ef9mufgKgSoKnCp0+Pr/3JxS1JvyqYV2ene20ujMTebDgJRGZURv04
TPb/hzGanyKOOwxl+9LxVmEIcddoojseb9WwJUhzqxk98jVg7F9GiGegEA4L619y
i5WFDgCakN+mw7+iPwLbZ5WdQx1OmCg3mJoPQfLf9oZ/zXFbLjcngNgi2kh+PU0w
DWD6QHNXFiIEPJXvmpkXWJofFcqEQcHie1s2mKJTvRLmU2lT3BA83IGMKyPt6cvj
jw0+oLOXzj/ni+gqC0bEArBUkVyXPvmfJbc3WkGK0qccxIewnpwIp2ggAl0B85Xs
Mzc9//DgQBxG56ARszUL66tPAadEVFIvXk6AUPfGBOAV1SaEN945HRht99272ieB
GLjIJrrCanvGB4271oA8CTyg1LgC5WCQjfWK1GP2EqdIaSfW6IUN+KUVu1HZvJUj
yGQQZqBJZ4TI8Moq3Gb6xXdqKI2wjZYimmryp/gcQrGb/hS0LKsDqrE+tgWq35dq
SBxijKIZtr+9lBvlSVbguLC+oz8Z94jaY6l/hEUIAFy7PV51PFND+ehSeD5weQgg
/DTR3Tdnp21d8ib+GDnhLeE8eiVLH7gX+DxAYAIXaKhF8FEzk9OdU5DrwWwXTAfq
GCC41liKfYGLXk9mv9uLfCEToimxwlJ4EDUSm3o0Cy+dHjVzHGAOOls/j/TikTvH
VRf26S57vWOHxjmW2HnVxG3BNKjO+S7tFIJgx6FC2Snbbk4z7Am7kecVkKX9qqWS
liJlIFiD13WeQhQpLS5Adh/JXMVg62VH2YJgr+aZ7T+5wX3X3ese2vF+6FD6ALu1
5EUDDhaWrpxMQzccdzLlr+EsuxvFHt19IQAS9UE8kFamGnyzJfa/RHukeFP/LqjJ
6z6e3FO/3U5U7lppLP1wvALra8qceNAXT1XAc20BPES+ui2u6kwtOX4ptx9noieO
JFJoHOC2bg/eD+r9xJ78vSaip2pLqvZTmoYNsOHKRe7ZiZSD3x4AwkLAh5Q4husW
WoTDo/b8mGaePJn3qal/ncsHWgZEzjofE3ddM2jVOhlYnKOpBJvXy2+XOXzgA7hv
JH+EB+I3XmodO+lSatTjM1nxY4k+qOGSmtL6E8YZ2CZk1pzlDNS/rJUcQEe4j7Bm
DF/4mmnxd/RWdDOz8Kd1YFz0x3mg6TWYqnRyVK0JZIrE1KU1L4B4c2123f3gwy8M
n8Dz3neRZk7XN2yh4FV3RdRD83VMtlttNIsxHOcmxmr84GQmEGq3vmct0eLqhb1G
rd/zlURui3zCtHl/XL+A3hWnMt0LLj4FhCqFAENHy3TXhxsZoxU2UOYnYWp4dOt/
yXNQI65HJisyFisupKs2zICiNbfAAqyCcVenHkZQfIWhWr9iMl7hgNDYcqBsbCa5
8XKGlc0SLLarBPqzQOkDdQ0ifcxeYl4yp/O2L0yGdSQlHjTk4CILzXv4OdDTaU92
kbgLHXqvZHvEppjBopjx6BaN3AfitmuViQeJ71dcZoatNjL0mD49iqbyaicMIc77
VU+DA0SancP8J1nFO7QkZzft7KIAbw/eiSdP+pCF686624S80uHHlXAgtrP3aMz+
SDIF0MUsUBIC9AWEB46Wk60m0IRZeSippHcIUKLpzDeGFtw64Ok9a56YFb5NsnTz
m+p07ed41Eb07QZMgX8gox34HYMP+Esqewco0X+B6RUQcXhYbvXD9ha8wFy0dzP1
4jEjEMXAEGr8+vcS1mxIVW//Ye4PowtcBY/XNlMNrk1OuEOd8jPGMThYB/T2ACks
T0rPpJrpNUgCIDNrWCj+XCBW9Svc/QXrO4e+sFdV5ph0jYymQj50y+6Jc6fZvtn3
eaXV2ja+wEh6L2AuJWMALhqlEvXyx/6wvU0jjqDeJuJBvyguIpS3GQNExOuT8Unz
IzLOGHjDCC+2t9gjkWK4ncXcdw1KILpu1QHXfLNlWr2qGF+HkkualtXJqp8irE34
VVHzxsHS4D+CBSCeSYrbz7X0/Iig81MkojPZovIj9EXLLYGtTr4594P7hcKrQQGf
ULDx6cPjED9suxw8IfobFSDdLyj0Xfsk89Sd4JnuoUgtluRFhELC1wWmxDs0qVC0
0HBOza7rpzWPHhvq5yCxOdFgzOb2NlJjuQq35noLh5wYiV78QjZ+85fmpO285FMd
11RBWBAfSIhgzNFru6Rz1Tzk9YveooHW5ofImaZ/UW4Z8+2/tCgF7B/mGAAm/NYj
RA3i6Tgn920Kms1uIQ+GdnQpCac1GDhItT8KwBtf3NH2P14RvLxiT/+zFvY3Jno2
DYZYiBorTF4o7wx1qt/7P00D/R6y3ZEtQTs2vYjPROp2xwyuo9r5+qEGfGdH2R/U
C2MEdaR6tvGprWNnO3h958lmm8nYwPMxCSGNF9Ol6rSGlqR5deODP9GXRLyBi0Z2
60vLSiPLp/wpPgZ4FlTAVbfp0Yu4NmU/RB+OqciQD7idJy1gyAfal3/EzgM0rDLo
U1MkKzvDijFIY2eTwGZ7hEcbS/tvCE45TUTEVoLSMrgpRkMAqFNOzzCO/YvDIZyZ
4nWqpETPz/TaYiCfL620PKAiD7RlnLQ5g4/zXhaZv1SRwGsQGjtgBYWpKfJbKYJ9
9FkOO/oPWeoYCluSzbNXHVCmCem8jAEeJuFZ7+jDS9I6xKtBjoLq+aFLijRrhkEk
SLmtW+qZ06vp02bSc/vO4dO+GS12eDmdYpMIlwiAWh4bS+Ld0JYgYOVIOsY7z0RZ
5bmw/0jE/CtMKpEH3JBDNgnbDHviYvyG0BSgUGCtQkeKnh0nWNYa6M8QxKsrev/p
cmNBMmcbpmP3Fz6AMoUSFTJ2E5/dz1fT71iSfxpUWHEWquqeYTZllbfAkeCqjvyQ
vkRJSk0lQDPTRY5kcKS+P8OmNU39qYsdq2gnYQ/RqqJtRv1+Ph70bYA6IgtiJJSn
ZMuWbtmqkHQCMWG3p7i70jWUQU9CKW8f6sGEi/pAABzvFRvP6DVEkYeUsATIAP8U
mjRnH5VBh5tW7bpNrljvjIljIn31HcPu05sCIXoS25Rv2e9AE+BOrtE8Cjo64Fp5
6kNFOxvkT9MF77myzJQ6FbIhgUfER6Me498l6jdHth5sLj1kB0FGg61nC4H33sOz
bgdftZ5NTR03Pn83wdg7fX0a8hclmC6PDLaqhnzCm0YVHktDCyA0RzzF0pRQ89CS
oqw5YSM3vpnAedyw/WjlSjNA3GVvycMnN3Q7YmFyd992jj++kIZtMOJm8OugTpZ8
3VUDOxfiMUXcOqYqQX2dziEeUMuPFSXnwzCc8ovY6Aqkh/ktX0CN1BesrHAY4uOC
l78BudZUBV0RV5fUvoLzyJe1hfYkYBMoSPuaQW5ZlE62o94CrgUhN0zKahO2wVJV
441tCbN5gYMMrKrmSXj7FzCtd0pPcbO/mweLveo8MhXi64ZNAyO4VlzO5X6LIsvf
nBBxElZKsrTiA7AsChj+OkcuKRoe8gcnft93R/gJVJMrThbxeFNGKNsToK9cqaFC
TQxbXaRVITxtnU8gx1ErtVFN/gtlLDYC46Zpw3+03FnOO3n0wCGNoP4nIHpG/f0K
SQlqOecceHyvh20ZVHr2jjiC8HcoeQK47O2RHjY5Tv5qm6ELz3MQ/Mk40oabXZ1a
/8TFx51bZggo9PjLWVo/bgsVNrKgN9BTOdLaf7Lm9kx7EpF2d7RixElYl03ra5BF
oh2YR8MntmM5e43XNnR7d6NLSbvybqBl4d5XllSzXdORuiDk5qGkGxGEqDoJn6li
DgBDO7DOQVbGKwtfLbaCW2PQKkl8Rbih8zDUVbS/DofTkD9/N5AhtORupLTRmkhH
KEyHPuTMfvxMC7ZJ4LFJinu7i1q0GjXilwM+LR5oY8rz9S9eCXLynYahvKOANZQc
jEpB40EdKpoLcg6jPbp90+iILow+ZLBe/nElefSuA7/gdwGCxj/TNn3fZ6ijnEZd
fgvcpIHiWI/e9iyX8A+RvKmfQ0HoLazJb2oV6fF/2Jflv03GyuKJQuBS5vKT04m8
Hzj5amNpeg1fK+Mje1sWDhyiEXaTwvnJj7gJEu8QK+bTp2Gh/2eiZ1d/bH7b+bCF
8A0f4+nk6gJJIdtp8vzSJT9S+OXJDZd+pcEKAt/aeQQq9M7aaU8SGXLxOzk98HzJ
CmCv5LT21Vx1WpLqV5tlqFlJShxK4VKYWBS/gzfcZMFFfihnNubLMUN48E1T7Zec
to2qUlrsInZQvX/2P4uTXGyjmDGJM5moV6NhC+N8mp0XUHY3Yj7QoecOA4y4qSRc
+s0Qe+yiSZcewgjECwKVcL00ggATGKDrqq3x1e5Cbt6skfN8cGukGO66mclMJTBC
DfA0oiuIdGFDCTrL60YQoRDgrJFBTQA8zcqQ5ThxGoSfNE6YEVkVPsYOmVT7k5yW
DIPBK6a6mBIx540Y8/U8p85zDWf+61Xoq667rORsX71DwUl/TBOOmal5l7KuJHT3
NsrEWKzmLQxTe1S1Oj44LHE7F06r3WYwE0VKJf5/h/r8xABWimAa8VFbvoWPj8r3
3AePiqd4ZPJB+v1P5A5ruZsskTJBWYjIHczBsR9Ile9NlAzbdokK/2PnhP5JTBey
l+X/JdXpnL9Hai9IxR5pKMfUKmnnqrcsopglaXWRHCm23Tm1DBabWLVdjEaZXWBX
I1+6iv8OONhI/P7Pxu6Erod6qRXLOwB+jpCY7VII7let53aMXWXeOKGP44j2XA8k
Cq6rSPQ49uAZBHShE2Q0UqdQcPQiHwWxbOEor5FdCNNh4GFFwilMTp3IPmWwp6le
/2VwL/rw6M4BhG51VVT82z1Et9hZgmVyVJ8PrAtHpeJoJFSSyxaZWVZcsW/AxiMP
gsbSgHZpStLGV+DZo0S+4jB1NCCyBh9jHxF+NDIHj+Bi0bqLhxrKTT+A/jecxwqC
RvKrqq6rPqLan2s6arR17nou9UEu2mYzg4QVWyHz5FfvUHBODnG4lt4594x99edS
y1NsZXKvdREXY8D2/7Pra35HbwCSag1aVpuJJh2BEsrdMDZhIRgvRBQexALabuM2
xSy4LUqCmtD2RDJsMJfGCoGv07cKdnkFzeSzBcjl2lWg0/307QUJm5XPwPhP5Ue7
sO5LcR8Jt/ZmnMt4su4DORVO5dFktSmNaFFYTmY74s78eOiWVjy1w7YlBjfqUvle
WkNC5z6CWgyRJCmgUiWHXLgA9dYVgMvFM13JauYE2F2ESTxji6DPeTSeFguiKKu/
7ZmQNSNs/+Gc84Tpa6ZbB9hFjJBOXZgmsGHgEJESakLjmSIJKLnyM5PC9Y+gV/At
lBiJq1dn8COfkecXUTrPhjqy6Y5BDzPZxkwo3hM4fx869DuyNty4zEakxrAJIX38
i7MQuKLBe1nS3wvZAIird8pP9zE8CCiV/txNwgI4A3gnc2cdcDXon1eFnXPMXmCI
F2lSMrMFWv3vwZTg2zTbhY3XWRqqYWazFG8fGUlxt96rFp5rvPtxyJE1LYgRnaaN
f2mA9TgtuEHXwiG2itSOCSzfbxnS52WRZACLEPqzn5OTypEq83NWbEQGFFVbXosa
V17IEtPO7h3OgkHWp4wA4+1cObSsELehxZpdMDbXsN0vd/aF77r5TOsKZrm9rwl8
4KmPBXa7akV4xqHlX0s1uJhwYsAnOF/EMQfJ26qUEANTNVoGF7MF2F2BiPKcplVD
kYHHAQl9vaw0sPZK/+GRu7kVye0g3Qk6kpEsRxIBEDmvCFigmV57OC1sAEeTUr50
xwBboRHG2n2yqn5pI9wejRBp9G0DlFHLbX3Pfwx12pwiWI3787Vmb1JMXgoC90Pz
PmqG++LcqIJ1+Qv0iD6FfHV0rA0xkix52ReGel4QCWvj9QRL4+Du9CNzOndNwIbb
SYaUkWd+0eWJA5+5KcHKkow+wcznxJb5iRULVAoRUtKx21qCW5okhNqkRRBYppkp
oF2IqNdcrKtBKlgJOfBz/w6xvmfuzqWsX4fcaFM6jiblGbjlbyey8yoFrG+39317
pI9y0OGnivcRQmklSnASRCROWnR2hFRdsW4evhTrryMvACLnsS4Yvh5diWAdShFf
UwursxGf1DpvyWp7j0FN2XcouMXbsNgKtOky4mlGfio3BFqvMuaEEFea/Hg8g2gf
9Bpn2U6jXoj5TxBPTYGsu3hsOG0Knrp0up06MTkafFci8yoP6Evd9yu5nxHCj8Cp
k7Ax7nxKDn8531LfvgZa/aB+EVuu9FmIKX13P1VytwZxv1kc4wprfVgEZAY1b/YQ
tOE1iids0UU6WdhYKUT6s5lzKFE5Xb8Ix0aC35aJ7Jh/CdPLD0Z+cXPUsMqiMSlO
JoVABE4rBm6pRXqSZEg9S6DBt4AOX3I4y0fphuB+HpYwCrUBMORVLv3Oyi/WeMpg
JtZySz1ylpL24+oPDDlFZQfzzmN+d0FJPLSH3R632uczfxFZzzj8C/XCSDnR3LCc
SXEgEazcslDHEmUJlYCYwvViwOzdKDeU3WidLg0O2OMaXJN8AnA4wjDbnpx+wGFX
TvDCRMjwN7xEB5QikvGWV7Ga3P+Ako0hVzdUNFXN/E/GEZ9RUHSKUy6MtEmte8e4
s0BMehpgafdAgif9UHlwEPHuAEF6xyF8Q7o1Dp+fHpsNVhbt1TYQKECjhEFR0p78
3UubFd6MQBtdhbeAosEAF5LfKz0YaesjhBvlfE47Ck442VPJMTiJGgItFd8BgqCq
A9D6rPVpTCZ5YSidqi1Jr6Dti1p9sMBovGBnM4M34ucdOh3UQAWk8oZQ483Vh+Z0
ddPGA+cZ2ZNq8PFWuWOqGNXfMD3b7oQ7AS29UfuWgN9mMe/Ons0Frv28Zm9ZoeXW
TuICAexHPJotZAu0dFvF8ofbzAk+t4NGJc2yNHkWq+COAZBvqiqVysZ5VkIcXOOW
vCTsboLN7HEQmh4X5wVBODYM1UcWJUtOGv64Jr8UWd1Vw4hrIHvwwBAtBQ+5lXiJ
FZE9yYG4/F9rVO9fTdn9dXwVUigHPd9kGYZjQXktZZA1Cxr6ot1iBh8WvgRLFKi2
GcamPkqpfYHPe9pJM2ay/i26zCCa3wC9qRqA4+H5Uuosav6wXyqWLkbNjkk3BOcl
AkzOjcUFxfsJZYawK7bxXkOOFhpqSCKzKvS+wihskDXO1I29jXDQCg716G5vRPpR
kPOhuhEwtuZ7HTZKD4Pa/FrnYxKRw7XGKK1xtykc5ugFn0BEVbDa73dCdLUbpn2h
VgWJY70/GhLBdgNdpAl0Vtdfwko9GEhwINZiwEUrZlRXWxnlGJN9e50dLLXcDjMB
hcIKdRTL/PFNPxjNktUVSalny09H4pPO8yIwqOGPv9lIZVIlYUqbn5Y6Ej9BTq+6
QROvf2jLp4RW51RbyKZ+nUzKRHFl0PmiOH9t/YVRkEbf0Kf/SqkcPQUfBhGMZ19J
e4f4/bIXPUslQSiMLwbWzSKFK5JqvPRysC20raUvxzjpxhyOIGEz5thwBNDsTEBb
wEFSigfmujKKK4qJ/zsTzWRCyX3U2DpibX5kJ5KsdR8VMduEgOIhKCwJR3veuYmZ
gPvU7oA+wIor3an6nOdYRmTRTwQCaFs3wRdrV5s4mMm/uSeOs5mXhX+PzG43BQw+
2LHVwCw6rftHDuE/GFsIwchBk6+uRoBhJn1wSbOqRUfMhmxykcLV9S4R9CETD1DA
qz+NxituhIO1fWVO+Bc3zKm/+7QWXRVHHLTIdoywSx9X7yDMjWyHGDWii5wU7Tas
m5K3DEN5q053aiM+itO17rVADorqJ7B356dpd42pqlPffHDO82Yba8rIODdudErt
a0Tx41bdpuKLDPzqtQ8FIth4E469UswXEFahtUaa1nmqh4o2Iq2pb0VSlOZDvJp2
7kgUeyk/6gI5iaYOIayZlNIGwR0AB8VJUgfjjC62P6SCWaDn2MiOppufN73QuIuL
yEz27Uj4XctZe+xO/e+wJDy/C/XOQojhRwcprsodoBlXPhnCIW/SVm8dRR0FcFgS
7y4O1Miuljx2Aa3OUc4oPeWvu9smfP1afRr4Fg1SieQAdWAn1wSPA1XA/p7LLPP9
oTrbP5WJQ7RTOs11aCGXTfD1+5cFwODgRuJMSLQNTjD6sCixINYMKLTHbKOLYMEE
c/u59opLgiHd+2iTIZ6UiRnc8aewRKPgjgzCc3EJI+DO2GgKrhX/29GnQMfp2yvK
1xasZR8hycTk6IelmgFdvpJnHEvWM8l1+22zkhCHb/mexM5BnGcSeRhfCpl1+ry3
sEKoiwTeSAI5LhUTbAwhhAJNwMmVB+NiOnLaxhAK+FLlc9yqHDciGBFA1UUZLBAx
4XrISgFIlt89vDI51RY/NOUJK8+RvdPwII6jvCx7Y2unb+fT93CoqXdBE/D5chdq
YU2iGdbspLwjvCtVId3Zmg6ivEgG1LzAX5etD/a0uDX118Tiy+eQhtJm3ichdr+2
qBy8O+3rZepP+gjiGmJi0JEtBsTQPEpbEo3f0g6cDbk7sYnk8ehYPFQfK3gCFlsn
SBVYDwfB7SEZu3sBqGSQop6RAgAaKVduSkmLYNcEzjxg1Da7pun9n3M8QdJ0/Bwx
xdf+wOiKZYI+LOVTgMBw5SU45tmnQ7CnJ2B7yX0woPPgLz2JyPAxKPLm2MIEbwzR
Ja3xfFZp6s+PeI/SKQdl9fdqa92risHUqSdzycF3JGW/k43AVwRfABnJhSxKlB3C
7wX0SNZRmdzI+c0gj/5gXOpOzoS0fKeg/qFbIOTVD3QBze7VvR301QRRu115NDkL
BcPeKH0Vm2tOU7uifChdkvmelqp1LjFObtYTRQ/g2VIncpBda/Cb9DCaBaNdMvpB
IJK1ja2iKxVdThsCYpQdxQioloO0VZbvnzAfHMvAi+jEcktu1kOF09FwTUheqsv+
jZyz0n6V7zPDiWPiYQZD7KbCtF6t8+EhA9JPgGpJOIpvvcXQ2cMzK1xQtbDt2asx
MJ7gtAepWG56tvs9cjDfE1fzDIXS5pf+tQpvFknqZJ4Po9wwc3mFYbEP9wmzVBU5
rPsXw78ULrmUjzM7Oeh6CK+597wFNcuQuJwcHeKrAS0oXJOVvrashZy4N882SAeF
XJ4Lj73VwEXF1DY9GCOrIQ5jSzO3H03Zve9dak8xhSapNWhl3CoeR22pCNW+nyXn
55UelAKvGBmXJ4sl7SCtL9AKELhzN+WA/mZLir4DODRLougTiEApp31UJdE8j+eF
f6BzfTFimnB4CFQHTCh5PLsIGgxHEjpn6sBZhJX0ZbmJkHat53cwpd4uWtVMgKfG
YPVttVO6aPVqCNYHu4LWyUkrENu/WTFuea9t1zVtFzy/YmexB+0qlxujDjJdxwaP
z82tMU+UIIRwRZs3zBz57BKiMbeYY2my3A8MN8Nci4xpJnQnD+XlR3YnAdWnzitk
lVLL1DV/HQ/Q+09FuobMG2exm8p8SZUe4SE189QMB4GsAP4GynyYIJshkosjmN78
N6wibI4JTvZAwkTGMZD/Oc9canmI/7OY/mV3ouDOIvT6mFIw6DYbVaXE7bxPJXV9
8Z1Fvu9v+TkB36ZPqJ3192fkRe92Tu5j2CAZH9BuWQx5K3tuhemoK2dc+xoQC5yA
3/3OoD6QA037mkTgTBLgNpSmhal/Pl/+bB99NdQhzZPc/4Hn97jsbedakDzHXUq8
6eLHP+YkPDcoJUILiMq3GGX4gmMHLtR9rHySxVTFr9ltU405B50heogpvckMD1Jq
rTCAIjHwILB3FSdjmZJgiuDIDebkD7EA8tTMMeuPwD9Pszm46uw+Aip1g150qYxb
vyfAaX97IgC4FaEEzTpfeUlX1S5Xp/9kE7sckBHZW2SFr1WJE6vLUcFnLHVm3prM
F5l6fot4UnUBDdRx2pefu2+wTe+9xXVrpVlTM1H6QiCbJapqSEsy6NKu1J/NHaiE
I75y6Fz3gtfFFO4syoAXJGkBCCg4r7OMNEEdBs6O5h5owin0ScDbQ5N37/zh510B
wxG2SSZP3IGn7vjOjmgAYSldZTLhvniTsWSNTFCiCsGErHIqorYi8QNbx22W922/
HL/iWmlQciyMDIQqaNl79cYMYnVi5JxzhPqaGGbKclHPCkMw7imQYkngq9zFvCUc
dK4JroWeq5p3Il1di0BvKRtQ2YcwmLen0IjKXSGRTWFU3I/rsQSkJiSjcb5+zcLP
3xzjVoBdMxtqj/r3EvJR2Q4H5c1AT0iOiSnGMgzkR/yzvL57U+eqGHcKY/4/6Yow
J10goKGPApccC0O73paAweG0vPyEhJapRxECQ1Gb4/xWnpJZZm2h3RCFGtTb78aV
ZvuMwLmUXjCtS5v0VLTpxIKtpCmPc3nGV2UtxQ+6HfGa8uHRDKc5IBeV66jdwx+/
862obzmK5oqoFe/etOz8lcz2B6/b2yEVesvx08KiHvJ133gfxEMrgSZCMr6J+R8S
DVwDN077nDOFgI2O16lsaWeqrl6eJ2HNJF8rJPgwsrzT9iy8w1by6r2tHu+NeBWn
uOzLm7yDUWaJhmxvtXfs5fDo8uRyKnGSWaHLlTl21If1qRDmE9hr1c06y6lT7/ZV
hkDE1ADsu7FScpExwwKWdYmUajlnH9IY8k3SMa1AP7sqPnFaJO4xt6Y+U4uo4Nzc
4llcvazMAhqv79idwB3lXyhDixvOiSzh9bMNu1nq113i5jCg1BeDfAdXS8i998QH
xMvykX/nGH/RelVTAt4qGVVlL61va69EQCs8SETnbYAQoFwmhYYQq31OgUwBge8t
f8Irf+dh/rZHoTDY9sMRq6wAIqxCvYj9VDs/Zs2NcVtoJwdmnc6RJHw2rmpRROik
QKn/rlSOwncHS2ZZEGIQcNtp5mAYmvUgke3h2+1hnFn0X1uHnkV5A8K3xkcjnEhO
x7RTCwKK+Pu0VeuuZMN6MkGRk02MKj2uxG64ixuZnYuCyzVVTsTJrpvQlf8NbidO
RRg0jiCLiACmaoTnP7KJqSep2XeHkFS+QBq9wleIwlHAHKnMWDlif3S9pyx4fapG
8rZGykBp01PYBhn500wvdFJfzZQT3qhBFVicb48T9VLdAkhJJVY+wVpZKZza3biz
1Z7sLqoZwz/q+QMaV30WP5sol6ao3G8K07P2+cQoQ+RVxP1l9dXbxCPdELMu/J5K
DxNqKy2n64a2CIK0Bpce+e3hR9MSQ52VbeyUb9uj7sfFAZeu8xk/9f5e0p/BX/dD
wQmqQtmhZMHB5suZnQgi9UfjUfB8GXH3wI6v/R86vTwX5DFwCZ+xwkqNHsiCoEE/
9PBDDK2ani6V8Dqlh3ZY4EhEfOFNkI5Mn7y0eT2QgxRGvZny/QszBjJBNLjxyQ28
tMIg0zVz6rTIbVjEi3oAbouH7aE/qhabl2wvrzMrWR9180a8UTBkQ1++EfqwqO4k
V+Jn1/BYpsVNv1uaQ+Hn198qj2ssZGsiAmNXKKW+XXoWyINDvpdTH0NDPG4CLwVO
I2VXnt8xvS5hTkqOy8KTuNyAWwvQ95boD0UJpwRIDdBfkh5y/DHbvmuCvy0JHKRb
kq9is2gGvFUz+miqc6KrtyTYezynx4/tcGLBJNg5b4QPbt1ITsrkFGYv9jywFh1l
nsX8qAtkVemGLJPiSIf5aDM+v4MZNGyBgBO2/11DDZOr8SWKThWwahVv+QmyxJua
WQpWG9tM1QOON6VCRRtqSVscJjrRHvZ2cvdAsGDa/jSz0dEUyjuxKPzDH6wy27Gq
5LzSKqoqg6fB59rawAA3DZ15MJbFQd83R9sPIE6t6DkJoGn33tYow+L0Nhw2UJVW
R6AdyUVISF7ZJPLFhYHwjDkIK0yY5UbNiksfw8Ga0rfx2PNuM4undtstq2c8/LKd
xUeyyu6tazTXoIiuECHtliuLvWMBt4X6cwPQUj83+Sgn4p1ymcpWNPJxXxEAKNF5
rlFW0bpy9F+8Nim+ueqNXwW2Cj2aTGeROFlCITBuBP2VahgL1TOlYDVSEGlmWs1f
RmODGZzNGzOggNTS2yMGemJv9ONAwD25hu9bOipjfwdNzQOI74M+oyZRZjDfC9GZ
/T5kbiVeJ2gOlDD7RUHvzupYmCJzCIzPR7+oC5WyDBavWHXxZM3ExDHb5TvMi4Ef
3mtvWeO7ilxpTG8D6y5C0gO1s8DzV2NR12YsV5/tukqM6o2l48R93g+9vfklzLrx
IhKqeB3WDcSYpd6A9K3xNwCZrx5IUAiU6lecuHPxcu1ozMm6AOUEIcHiZxpvP0zG
evqdlkFZJnIP/abPLLTJ5hjsiuumTsKQW885ei9FiwstwUhCdB9vAyEQ+8GXTbKw
HwjaglTWbpCmR9ijNR7IN6CLu+7BgkpxSA2y6Ehtoe/BdXw2/XtcqrpZhawn5w2E
gWYbhl3ld0MiGs96OhDmVhqiXSew6HXbuZHWMl/eXqELjGH7xJU7QsCrAAYpupsO
jDwiPPltJo0p3DxHd4LDUjKWDK1jbfcADlr8+IutKi7Zwu4tgOn/F0YmeXS3/q7j
lVIWRfx6DUaSUAsJYD5z2QDKWeDYRRcqvKvcsNuTEpJN7NT4rtX2lhbsfuZCrQ/K
cYi+nVR75B0NBus2Oj9wt3Tdhw6wlIG71THBYUITwflyIH8eowT60DtMzGgCFhg/
qDjjepTQDCDiiPrcGZ8ehna+naCYTECZ6rkUfqp5Ogj5uygFxHTIaaL7eLVwhQsQ
nVPzcRfo333lXjanvSuUOuxL9ntOzktAXvEr7sI/CmNUQKM1kctpcTenVfjp+xz8
5QWUv1Ndk3NVgdkrT7uo1TlVL+cu9+/gI5x+XeXXvEA5WK9O/Y4SkBZTfFbTOl0P
f4pQJ5rUPG242tvdAoRpJ0dLER1sBvo+CxWG9Bmu8q2qUvhiiRTxysVT0/URAr/6
PH4Nh4S4mcMjCGyVWhpuPBRg7ZKLwqjx7n7YeCQFTXeSaJd5eCWZEFkWwjWACJ+d
uS3nHeIbhGUVomzoggGHgTIxpLV2ZT+grwRQbcZnAMUqe28umMg4/cTAUKccCcEY
9iC0OUOl7wy8sTx1cDajwVVRxy7zsUwhZEriLm0LsGps9tHgbUFfCjgB3P61XWCE
ghfW5F6yLGy1zA84pLjlmc57XUMs5xyY/sG/kU8yWLGlubsgDS7AnqqhtYpNi2dg
/OfC8Yz5PvahTOdKnDtBPUjCwLJX0MfxS1h8pjOZuL1TcoeTzjK0iZzSbua0thxY
54keCiCC7+YdPWoGtqsXt4x0B0m7SPq6kIHRJX03NCGVGC2uQfzDygkIq9ZiU/Dc
Jch/2R1dUZ9Y2rM0BBadmnJU1GsGMdOTaGGAVsYvzn1whAIcRw38J6XdOwWVXb4a
Pwz5Se5vTEQHiWTIeFeSTE8TYk4hbFMc0F/qtobSZE9JPsSyIt2/IiEGx24kPEnq
/nkxyYen2xhTcUDxEvWC50R9WVjB2hdBBDzkHciJlbcJdcAYh8qd9HZpAeW36PTL
fW8IUb88/DYX8dpSgtTEJC1H5M04JAYQiHttD/g9JXlrGJrgDIAF/PnSQzET1Vbo
WvX4fl5NvFkmNgBWNuOKixjRPn3+Q9QOJiOmeMeUiTNpQJv6O90Nyz+RsNNs8ra2
Rlq+0Dr3HzoHQcWyZlVYCRbLfDY4Bvr0FLRA06/lJuwKQpf2WRrQTpFSE2TSuNyr
kdkmxseOsWGRbnBN5+H28TKjaQP/OpAtkxtgAjgOLcXkz4TjLMuo1CrQdzGMSn28
MjtqccXJwCEu3JY3DFiv895B6FYtKBnUZEvXy5k0puseYLp5SLMxbU+03Zq26Pg4
y0K7K7c6/5IUBsv1ykYu2MTr4vy+w3aomDf8HF6JgUFPWwBbcXARDzzHDGeMA0dv
MxLaOWae+Hc7mhjtv568Uz4+TEY0D+zprASPVbpU47T2sKcH0j2++9+wmwVLz26o
YALWcR9+ZB5w7Y2gQsp8nrfLrLmcSXl2X67hvhqLBo2z/XEiJ0fu/1SuvVq3MrZP
CAwYM71D0ANcYP9b6ejbNKFmf3tHWLbMmf3kvLvhtdzhTtuoD7/cGlmtHJcmKWPs
hrsA4OcG8cl2Bxz5hlB9mf2HbK2Gh9gWiA9OAFizRVA3N4Ks+4aFrhpbQh0X6SGE
RdzDYZkYZkhoTzuiwNuScvNnLYwxJcuckGyfKmqelurItQuF5R/tJQxfQenu7uHp
ecAIoXq0Yed6FSx3ZmKkzVvOjDfBLRafuwINtrpQK0VDMUESLBMfdxF1rQNDzux5
70nA1voxRLml/Qn+8KNGPu1g+gzAEYutVmxvXYhsOJPiaaB5eNGx52K3wrEoYfiV
zYDhP6L3Sa5Rw+4Q1cPPPt2l+e+VrexFX/CkvFgtA1aP8E08rpmGh1++Ev0pVzBy
2ETE3yqbr+TdIp+9DEmGBqi+Em/k66lhud/dTyPJG1rNuMPmi/p2fKfHEefJZkzK
xe7CNfw+n64KIV/RUBKjRKa6YOKssHRRVpHnA9mAh1Q/GhDYHkSp0Gm37hUv7T93
W9n+6FO8IUs5kNa4NWO//hw9motidk9EAmNmr5Al4BoZWPxEMSEE1th10m1whKyy
fKmyYZR5zcc9Elo8XCdmLJHcXBrRwUbPJGOEUKYUHWgvtfdYWpFuZD9bp8nJcaPs
R1y7YF3//UvBMWxR4V9o1lEsffrwW+spPOMgu+djrYfoDz+TM/tI7dcV7EmnLEi0
9s0jFkxzBPTXUJ6iZybfQEXRmK0yvIJiShPfjp6hWL7EXGpPaeSSv9j1WvU8WUPZ
mcQMa0RgFsimgKLFboR7+Udu1gJub03/d/lSmEsJmsVMFc6CNGSOnRG4QixLg1GH
DkqY0hbm3sbS6ZpOCLf0wfkzRg4Vh9hNq13uPGZcqQvpF79UTKP4mOEIz4DFM6B4
TxjysyANUj2udvc1e/iZw9hzPE9TtC7FlbTpx2zgI9cShFVsR9jS+RVie6DFL8Zx
Mt9joRv0axsRa2/uyzxPa4xYGBeM1faraqeyHrrWi5ob+L4cX7Vf0+VfBSm+BKWR
BcYSGtCqrXcsui7rWbOtRLbbTLWGKRdx8B2RFp4eguyGKkKbyeBr1nc2dFOYTkK5
0k2BejfFcFqMtndC6u2Lyp5x9E32PERR18vcR+WfZd8B+l06OzOfE2IdyXjnsnvG
xI+lr7U2otEapXxm9RIPaEEkOFKlwOIbdVhX/YQwcEFXl0UD4Qok/lgSS9i0bymV
2TdwqkOWpxLrNcNDeLqrfcJ+T3XnImiy1M4PHGfuVvJZxgAafUPk4EnlsIxbDJ4e
fINT+fjsCfwFq2fTBkhK1IE9XIZtPT87DcyfC4S4zmLOccCfQf4VFU9guv0If9Js
OWyr/IPqxdhldSA0fxFC6epTc5wmn3ZAgz9ZRyr64XuB+AwCgkg9ADe9/KBPa3aS
aLHfcEc8ECEkVuPrgwY2mxw1KrcFfvGx0Y3/yYU4E6SvBEQX2m5J1jkokxRCPKsk
QA5nPAOiPHwHeBZHitmNI/eWAopXiIpNWeujAf3sQgD415ni6hH3khX8Cjr/iS/3
5gf+Vy3GpswKZhfZDlqiruH9Xbrhgqs/mb+8Z3hBxu/gJqeNc06vkPi40LglfJd3
dTbkwvggA3enm50GIajyMt5C4NKwFnE0Ladmdmfqi1G/MwSXWuvDYU6zitP77yxY
Rbq3GP0bXA0FDCBafQJuOhOsHr4nbS4zsuGJXbTu5UALoR1FX0JgVy5W7fRX8G2m
tHPOLGIqKJxvRSyGpAtjZlsHi5S9xZxijLewca4Kw5YTyF7syUAB+atxMz2trkWd
NsmhdtaTEdgti3G7na851yd1mpdBqgOCh3si11QHtdx+Y5xu26T3F3ACZ8hZmHok
DyvvuvnkOHao32FRNyjfCxiLlmmbndGl/yDnSEf6citSdo4mcK8V9gDZuIZRVvkT
aCyfLCPy4MPKv1OBrbsyBw55GtySuLxEfA4TeGVoRLmWwfvkw4H2iVsFqLmmAR0R
3TlJ4foOGyi9PSmKTNBJGSw3kSsIruMTJHiAiELdGbB5v4KJL/hJP8iNcM0WLOx9
EDNAG8a06gguyMnRGq8WTC0EPYAhh6NV5HjEMvaONTq5qaXdfF5/nOMv2TtyGjVz
qmkBXfwN8halmRmOCHTvlk6a8OpcKkc/1NKruByKf2cA10yBqMkRWB/BMFcmIt7u
e0etu6LnpIEeQBGdo0j1ttiQRzZFdyfzUoHjp6qrZLNRcGO+23EM+gY/axwD+V9b
720+sM1HvwEUeQMgGGWh5fEuvo1HPkXY7z1DRKgpxG6WFmSAR97udGdjcfgm7dlt
jhcYEGj7TsvDReVVum732fzYTORErR5aGPN2xHnoiM3ITp0pvmb9FnvCuHW3ckDr
zP7/9r5RNomFJcJtc0lAYQyAxQRyZIS6m7j7r6ku9j5sWfOiyhhtltMzcUOtiQso
zphrtRaJB5rhFLd6wJ9I4pyCMIvPSC8u7iJyrbsedO4ZLGBCSjF8puaHb/oAMIL7
bgV0XdgCwNbNuybzKmNZd24+2AhlFP47Nxw9DQ0ecrRue8hRgcCpaNsZxA5h8z9y
xSIl2fppkqa0Ayskrfl45yp0cPnJeonmnDN65iX+L0Xur+OSOxky/aRC5eQne89a
jFfNnaWL5Mj6GdVKHV6h/wnZw1qu70FFrs5Gwsm7gI468afLKlwldIosVTXpSlH3
an0SCcs1J9t3mTTiyZF8u8izRY1+zL8eGwZnxd7O/nLIshN7WrPYiqiFGxNCsbnN
dVLwem130QWO+zhtEBwLijuKoGYSdUqU0Ncw3iIwWWImxGqJX706SBBiZusWLGnH
t1Wam09BhMXT7c+PbGfp5yACqbuNdz2ssnoGaiYk4qzeDfCkkrjZl9d5IDItEDiW
N6B6AS2/XrZJk4dMp641gMKHKiW5AbXn2ajuMa7LHJdAlxc5q837EoEvJwjsXy26
OD3msVeLnFZrEyDJpjOS1mGAIFKmYQNzCTfzPW05diGAi063RnJTzeBBTg7FvJjc
XT1OQpdgVJWNtFi2wVuc353XLCX+uomeJmzxUwMZ9r9AJ+5oxAOFPzvP3LvxO2uj
9eOPcNL/iE7pkRoXvaFNvXB9v+sZSjaJ3t1HPpVFlk/vGE19tLOGqG3kUhUKGu/e
cDOhFWiiMxCWu/Y/m/d3tUhqTbKc9uToC2Jo6kBUO2dxgUm3PDUwoIzR9+OUaEQF
FRIAkXGLPDxrVWWuJRtEfpPNGV4PMwmX9iCYiGFbIyh2R7xCu9XXKaYFjUt5cV3E
hGu7BQDGV/5S7z0VHAEhIX+REGizY3nXXsF+fqjbbq9a8pT5bkDx6nhDm7BMIB+l
gDmNMOMy5sKlktoyVNOnojyanuuezL7ybFpaun4cqOqjfpnhd/hXDEyP/pYXAIzO
njbBNRM5MTlfy86Wx72iU3e2MbOWHD7vhrANGtoQPGxRaTepxxK7ishnBnMnBm/i
ONGNzmoMlXzXzta/gB4Cto8J2z6J7SWVuIdtY/DtBJhkLeU23KGQR9Yw90+dsWjN
7IGuewKysw35C1+5tmGzXddZYFQyRhCxB3w3pFIXS4B5IGg79pcBsHDZKtPMlKxJ
AFelyyZwwl6IkE2l4P5wPjUN9RIP5qhsstvU1b6inxxPqs4Q6TIs7O8mtf2PjzTD
I5cdaehTCAn/jskUr9dYUCg1MzpJqk+9YV2Cnur7SiXv9DjVQGiYfO9IcTME+4x6
Tf5s8U3fA1ozYMR0wAga3k8QAXrlnmWGimHdlPYYWsxTG1rojQEptfHFyoVNrpQv
eChjzxtMGf0odYXdHn4NEkQuAE23fR/trhDnLdPXzCMUFyqZrTA7eY+8U5V5RGf1
hDdnczR8SA5gNhzKNki1HxUmu8omi9I3X16zhRF67bKOP0zMQHSrFc8IDG0cJibW
8cZxPS4PsXXI6BdkymjjeU8Em2zuikZrHK7ksusloXnFb6T8lJR+90Lc17PB9iKh
iMGLUWByGTcAXmq7R79ryNWFkAVgf/stfcJIhLXn06NRQMz/qOZpHOn/n8yAB93W
sISQeIgHz3ukqD4T06IlrWX4E3PAFuGLJRpGpVFqKcxsZbPS3FVgzj+zqh5inviK
calyjWqG0s4+LjQSR4Rm+FSvwV4A9QXAoztkgU4v4nTWQ/IoUvaANH4kxyXliOpX
C+iLNanfG4uIgcrrbyhl4H6CDx7uWM8kDQfaes9NaYkq54lNV+KdhQ9emzY3oS8p
VcV0osLUlbT5eQwfb6AlHcRGKp4N2z8E0F4ca5KIoI3QhpYjQy8/XPdvXCVPFyC+
sfSLIXBevISwsXPFQ9agceC+HUtYD3/lxYuiGjHDMY3XXOeJKL/HCX/tHllgWtDr
Bm2gMGnm5ZdVOml2TTZrrY2/RpVYE5nE5Gticz7hueyceJzFhiJXh+22hckYZtCB
zw//Sq3DK6X2OPu4oDuiahhkjy/VzC+XmISHxNgx6P7XHJxbAl5UMkfzut6PrH0N
qDR+CeUviB91vt9zQi6q5szdinR8efi5R/oxV3z9X+pOtP1FBXEl2PcV/9wQIHss
bNtMOIFGS50sl6ATD53atrPpStu6lGwlCr/skVMYpXytfAUfNPO46JzVELYrGvAd
K3MCOw19yWgnOIDRLaN3Ezr1HrP62aePeM3oWq4p1LA34nu1RNllN9g7XoaloRgt
QZ0oECRmQz/ymSbMRf1n0HLmrmpNqUpr/2EJfe0WVr6qCa2YbFk2/pSvfknLWRn8
ZmXF+gVpPT2HmOQSP1qfgmB5DIjAUDu6YrV88oDX8N3nuEQ2zSgBABvZqu2RwnXG
2LWQpCzfiyA/Q5zz9ZLTZy1ZV65VcemjZDoZ4nQ0+t9ApQOAwJdslMwxDkBk4tOz
LORcdZdrqHUQoZ8+WLGZHjpjxwe7WQdMJ5sWdbc65HOcVVAyZOziSVP6FPZnvfum
Aaej7RTwV2HlGLWI1Wv1r5QNUhs1/2X/ioLUIOWSRiEDlcQz7/fc3/K+hGKMrSi5
N7RKSDIPQnbUf8Xn1sE1n6iZixtjVXz3m8uQshu/IQ8L12ZqCnVG4RKykblMyQEw
ejQ7z+0DW02mS2WbjcS7XMOgJ5V5qCW66YlW2cru5s+uYVJZY65VDIJ2vc7KbzTd
gTaBrJtieaxX+F8Rb7ClNv2U4vLSDgczN/Ryz7GRiLDu8AsKQcEq4IDb75R4rac6
cdTf8Jq785neRPCU30fLxerswD14TX4vK4FMC39equ/21JIcKPceZQ0f9iwbI/bh
eWr0IHn41fTBS0lzIzkJl9qjkPtChLZnxARk/c0ZPYEkvEgutYuy7j1xfI7KqvYo
N8GTdGuUCzf/XQ+D6842cIPMAiOBPGnBlgwvdaspNmeqOwdYkhBQitMBqmdxefR2
IaWAQM8dldUQ5kygME9nUQ==
`protect END_PROTECTED
