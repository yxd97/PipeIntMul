`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+YlozEobzR6wgQIxhjwwyb5MyuAGtMCdpVXvAFdzEXPToK2RQGHYt9ezQBQ468iO
a73AC+UMooV3JyTd8x60ieQ7fCXaV6nKD5oE+hI9xDGCZUXei+I5Q3L5mFrTiIDC
8fJ1MRSl57iAR7q6iW6RDYo4yTx+ub0VI0DgKCqCzMdWM00fgjrHkHTwytPkmPlF
ocDga2XwvrVin4kcCFeLxQ7InSvqz7EeOLkxVU890gs/pP4wqa6DJtju9rshKZ9t
PfcfRTCqVMMq2U+vb/aZIf5iIMKTbopaldjGxbNBicnUjCZQ2DxX7ac8/SkPRB84
bNuDCrntXRDsKjWD1ZA5ARpgHLRWpYsBsTkFln31H3G+autjugLEkValVi+R46LT
JQQkmlgxkudcNQUxGroQ8vSE/HEbluGqgifm+y17NMUbJh97BHXTGPDHtow/TK1m
5TULpUP8qMIMcrhFMIllv58JJ2Sj9GukALAx8qHkFlB3f8oPJSm7Nyjmf3oMNWbp
r1o93M/mYh8sMpvE4VQqzWW9/4mZDmRovFyHKNf521aHMrt7vBelBsf8iSBvXoKa
MCDNXmILRA48VVOEOKDAFxjsc3iOV1/5rNUTYhkKpNn3CGYt1ZRRjX0vLnsk1je9
M4GTkXFrlxK4RmmQPifqOCna2+Eb+g615yJNAce5DVi54k22quIegrM0OsQ5bU1v
wDq5W+/w6XpbdTHLr+Mto7yn/Vp9q7n5WIa54o/oWyJ0l/N5Kl5bNHPa7wangXmM
6Zby+YVNvP54E7/r72c/7yiCv2MFxmQG9nqnb+lbKK6np73EiKuDWZ2XMMz6O0UT
VsHWsv8NA2boobQLWtcGErpwaQBFOShktfsZDNsfTYRVKUif57KPRDb4TuTlvTCH
HL2OsEkE7OQUdYjym4ig4vLOjpRguSj5ycuKFwbSOMAjD/WlvHPJ1qthjUTcDzsZ
/5VJrISgK36qI7kQ7uLO55JzglsEMhvDsJwoDimoeL5JulkXbMCMBmBrlfabFKgf
xmaPMHtGF7QaSlTRLfZi6PHtISLVPYNZ2YtjVQrOmjaruBCqx9mMGjoDhxuVurCE
KN02ZFZ8chLST3Xv6uKMsDcVYv1QcijSPnr8HtgIKTfNlXrxsmZYwH5ZH0qrmOKw
d3NOMPegJ3k79zzQZca/hD/AIG+7caklrdVghmid3Bds0S4tYCll5LjrjA2u5bJ1
2R/yOuPG1lb+g6vpzSrJ7RyrxCb9ymBI9P8eSIvxlRrU4E73YlgoINl+Mk2BaSv3
KPvwaZLvo/QPLTIYwr/2sowzbkUcNjT75ydoKxN7vZVPJIBdqaMdT+AOvuY062O4
efJm0CQogfL8wsdPW1pXEJp7ckT9H3ca/XgGugKvXkwQWs/wdw+tNfDza2SKXV7P
`protect END_PROTECTED
