`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElQ2qRqEP14s9NmLEPcFWSgHHe7JnnubFcu+DpbqmVrcdP3JqKe5mPEZnHdN6Syi
Xz8kjTiOOUwR19uoQbEKjeO/KKFumdy4u6qPmDtZoODMP6yxsYE0dCNL1oLeixks
iaCoFd/QdQm2Idk22kWDOW0H99Ae8kV47n4W9+nPTMzVzPpOHVyp9F0kI/g3W628
T+eblBO8islyllW7Cl9AmMDZJCj7o08IB1a0LXnrq1VBuJo3JdMzUra3DyvQQDZ9
hLs4qAkjHQbNocXf4XAYvEzA6vGXC1D5aw1GIfSSK34QRX/RpPFSqtG4yOkQPWxd
MQHuXmb/ErmvmKdtWZjInK6XF2U29wb8nRY8vk5CjqnS3yYCOOUfZRjGAdSGu3jC
7RQOvjaqTdwUZyxjzRT8Y8dticF7Bde1VHGzhI5aP1vyB/fjUABqnuU/eG/gV47W
xGEFxliqQv8h1Dl7JExc6jzH/5QenfurS3XQ0EGXsKvRftKXZp0mwCHaZjeY7J2G
CRsIRAqDyFz6JjhcryYFLc4glZnE5aVGcYucH26uDhXwnQtpszdBiE4WuOZogD5i
2KcS+OmcrFEXxwXeIuAOfYdT/CW0jT0cgaEGejGI8Jz0NxIBllDmKGhtEEjeiqaT
Z3EpyoEQTyztVJB4e7BttzqtZgL28L8ivt2YwuC0QW+bhB/ddrxh1rxG1M5ifIOc
xJGs1jcdQDNgW3LqPfE4OsRT1+dySf646k/8N4gyI6aXUOVg5bgGT74rwEYmZ1aT
/zMZ/RdlqOmlVjfN83zWnI10EAhO5GiOaabAjZmLL3Y=
`protect END_PROTECTED
