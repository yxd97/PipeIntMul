`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gTD+66XeraNI3e7Ns7DBO5XoTUA3rfji5JyL2IbT5xyxTYToYoNoGNvC8YlU8Qoc
XPsi8hMOf4iKtdCkDRGovkAR1bGHDY67+rKNESgo+KjCImt9FAwcvzdlAAx//lNe
04lnw8bUU0+99n9SzRy5HVQfVhkPGAw0ThaISObSqK2G8nM4tO6FK4GAEkQRyg+O
iYvWrTFpzfo4M4ImtS4UoXD/hzgeqcjpDYXk8ScQLdIjdPLr7onh9fyg858IZNt0
MuLbWKHH0bY9D4fAqyvVx1ri3V6NZa4hKhCI612ST7JnvZiscvzcV8b37Y12IWo+
VaOlLqQ7itEHUzbDdBDf3ex4A1XOqP6yjXUvjriFIuKPpogxZZPW9xEwN0t2a3Xu
`protect END_PROTECTED
