`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o3Jsy/g/QK0+x5IdRIdZ7txE4eElBvJZqvaJhU5o+EqhYv+Duzj9kX9mF24RWIRX
rb8g6DSYX8Q23AgaAdoHc34y+WatiiaF3gotZATMOA8JILEa5Jyjrdlw+lurjMbs
oB9gtV2sY49cF8wltc5JtMwzzQYc3rYc3+U2+5EzyEnzeImAYGr/aqgDmocaAbjn
lKq7aFXHyrdO7qzPbctgxEOJ4jYao5GFrC8h4a5rQBBBRZcEdiedP0C++6M9wwnG
64enZXJHb9VnoZ9j483IdOLT7sYbfT01XTO6pCC1sw6vNNHlqhQTyUZeh2ggM8Nr
stwvuXDBc2QlTuc/lQU8y2RWXYvftrVr6V2kMJ/5hXZWGSuKdGSCBT0vwuYeCdsZ
P56xbgjEbE6VFML4Iz1H6RF99c1K3Dr5Zz5anWuwdeQTwKBrkvOU8jq+Uos/XLuS
K5S5LVt67VHnBIcJZBEnmXIhUGiBEh1ksC07vY4/VMhyk373bRx2mAcjPpv1Gjl2
`protect END_PROTECTED
