`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwVBGUkPVPQoiYLF+ihsfMgIcHjcj2KL2O7GsuSA7RgYvyjL2XWuOzySyAEDhQY9
QLsG5Tw2+NW41XTNN9cuCXH+RJEChbfICepeWfsUkoynGSkZtG1iirsppl8usTOU
XVv4UD+EOpbDnEYYlqwxS/NrxaJp7uhhRNbYuMNkf2hjAWcPhyuKsnnqGR3ATVTR
wzc1TggY5Ye28yGA15sN8wkwf1hAJmV96txB0atmfJUCisOtLClF4XCPxLteoKsy
+VKtTBYkiNCT96+BytF/hEtTLgS37ufmFQZVmDgR+xbAylh8ggbhe02c/fegVT1P
a7PdQmesV+OHJKoieJ9awomHvdwQBwSAbHiMk1m0IELodnPoG6mesUD4Pr3UKxz8
7PL+ZHMml5R26mPL82z5z354QEZWn5OmS9q2KVkG2dMriLJJZweA9pl+6C7/Bq06
etznvS3/UzuKOXaDLANasR5TcFgqIEYsDuz0LJINZ6YU1fmEQMn77Q1nfzu+BhF5
XWwGsEc4yO6bCpn0Hwa0qjcRzP5lcCXE5cQPP4X9doZE2VPeSRCRIe2cG42ol/AV
zs+92APD7gzZ6stIrSi1C2TOP9VyfoYVcB9xZb2bcTaLZvqRskuxYRECk424FFaa
9He4jJz9f2C58aqM4Lz77Tzfp1QpD8TsHcUQ+1aRYXEZGUzBmM1lZuKlMb0eKbe2
7l5bX1ZSSh99h8MKX1wteCuGXsWpphQe1C7J61kzhYAXlScMxGGrlwh3DNCvan1G
jKFHOByaeavMfichqM1jTb2QTPj0D5hMJ/0Eowabp6uoW3pm7KnByEqBUa5RZDPQ
/fb91g7oP+EgJWfpyik/QvuKG7bSaWdcWPm8XoLMoVtfPqkZ+x7iCc3xSnyNq0Py
ALGW4I2QCUJ0z72gWAsLg/CoCsPCl8QeWRouLSS32Gf4LQKLQVLozB6RtIvc0kGz
`protect END_PROTECTED
