`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMZPOmv7/RaWfB52ECiwHCsM17sbYJBYS5nga/jhe1EtGrl67hvt4/o/aHkE38om
8d3+D1l4obr085/UaaQyCB8AvblktG7BAEhCV3oO9x4ixq+nxMTXhHjPED7j5JZP
0MDL02dzwqwnBcn8LJe0RMQgaL4BoQIFMNfNj5rGkM/K2E8Bb7kqTRo6rugr953v
F3Mw/jCmVF4Rovb8Lid5Jw61v/0wJoTM8F5V6c7AVT9i8DVziCwro362/mddHc2f
41q9HdYZQANNLp0Iq50RaMbodNnIroF3MVASIT2PNIksRM14CcHuNm3HjH9V/XQY
rodOuafd1bryg9yyVrmxwluIcbzD8IvZPLTIr0Goi3LTEGeFj/SlbfRgCHTbx0Y1
PD7Jgr8l4B8DAGkR3XrTk5zwpFsFLPikPCMFmzAPM7JffQtHI6iuIjZGFAYWr3DT
C4Lu3dXFpqnB5bA8tOvFz0d3BiC6RCyr/o9lGr9Kz2RoRxk6BodV+MrLOe4cTw0B
bBuvnXlpvKCvLuQOPnDBrP7pyofIh9rsL+F/3EAvx4ZxzMtuG561swB6jd6/dg0h
OCYx5EnnZIlxNYsuIlKCNOYc2soKTAGx0bvWMvZl/fHiCaCf5uoRXI0uvE7innPN
cuWFVR1UD9zeK/C8HP5URRBe9ah4QuvtCCLbsIWubWNJ5EKBSVMIfF4FPisDZ9G+
wND5s/kPNtuHjJSVVR2NxR//7Lj2dO45I97aPJt3iH1zZ4HCFtH2IhAxSyQnZnF4
Zb1CpnYtONK+15DGlnYuGfEVNcZcNKczRb5oAPVXcz+Ks/nSEZAWST2B/CQxaFi/
NflFl5Fvloa+Q2ou/Mv0ONQeCp9Qpvgltpb7gQKssDyKbqUr17iPBUvH3Ukl5wK0
stmHsnK1vzxnGOtg4alrHBJyHW1Iax4P9MMQhMIg5VP/PkxPPsOzfuA/xi8JTxH9
f9ku7i1Nu1Y3KzMrRMmXtS2PEea/e3ppbGWh/FStuazqKYAh/wz4cF3MuNFL8nps
LxdT2GgDXrg1m2sumkdIdA==
`protect END_PROTECTED
