`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gQ2vBvx3MDwQun1/4khyu5KD25+t4wCBQpJyNVz2ti5oCqmUnVY7gmV2LsQ5ngiR
tzH77FFFfSgu5oQtO3mweyu0lG8KFjhEWICileovlNUQdtW+nvQsgJOH/ZuyJhtw
HifnQr77uVLW5YeQEjhy+6ZX2cfLNJFkCoMBMwdM0/9UdXSvXHH6YdKkmMtE6nDz
CaGynkRzcX9ap05WqWr80Zs3jOuULem1KLmDX2S6CjKDNp4jhwp3NtiGMdds74cx
8AvSEjI11vEYEmsLY4bgQuwIhxb59GJXSG7aqk/StHJcGf/5pSB/hYT0RA1yqwgD
OEomtC46bhdurspRs+rhgQ==
`protect END_PROTECTED
