`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFp5M3Clpip7sT2JmgESOzQCqSfiRSb7GFnruagBeqrv78AZCXgJoCHanRk/V2vY
8eRirF4W08P29I2/rDUyWYCJfR/l3WDT5jzpNyaeonPM1E9gWM+WVj7LV9Ujv9Ek
bPG+AZ25nPE0ohN+UPDx0kfMAFwzFqIg1kXupUL+onrTeoP5s/XXzUweewyfmMg9
sfDfyWIM9Gvxb5tUlCNNQIExJjLF/EXShCGFjorkQ3UezsKVWHQ3RCZSuesXdwrD
ezJW0ASvicnexACPbSB4baNW83BmUheWSsv/sQDbkV6bTsl2QqM1nkux6qjOsmll
ukIZ/Y95WBU3ATALW2M90i8SQyE+xlKkkUoiUSKSSeCtVRGP4bR0qVZzyxiOd+9o
q1Q5zeaggB5XTadv/ur8H3LVUSUbzDJ350gTLzdS8ZAglHsyXDGogRIoV5Sb2h1X
t34UjvtYgdoOclg8Z9LwxVuuyiHxlCxIHXum02EbUs8fj4bf7E3Rgiqkdx2txQI9
QeZvTepcCDj7qP2zllv1JNHoimCnrlOOQ0KUKR4Wte9jHoHnXNzUA2tfcl+01p/i
3CjmIpqBGOY6iLkR3o3yCWzkgoKQhB0LYlCsTz7za+KYNyXQ5CTXKnifqNs5z8IS
U46Lo1J2biKauiZmEgINWfJumYUR1Xp5XaU3OINK/J8mKPIPLkLuAJ4TVDSKydOj
Zqz0xczS4zystgzCXU+Qg0AQLA1WcHj+mp9e0VQstIk5uHYOwOBnCKdj1H5/A5Ir
`protect END_PROTECTED
