`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lZQwiqY0xpudHNKVXnnQK62am73NHgPohZTA6oQNS4LQxPG9TuFgK7Hrlx0L4J8t
k48o0C7nNk30aVSc67EJrX/rW0LPfsnODlxZHJFMCQoN9PEDBLlir0ClObW4gE2p
5Mpgo+bjDUwPO3uEmSVD1/W97O+owX27MjVrbQXdAa/fGU3cOuCJ9uJ101SfGsBu
+EGV8twE3eJte+Nen4ycUyaRBa5dq/avFxa7oK5v8n85YqepgjVlj0l3AxCuRk7R
5BuNA3XqooOBkWqMut8eU24isS/zY5g/LKffpmflk/858xmWLy4F/zfKiMJzYGVV
`protect END_PROTECTED
