`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0wbIYYEH9ARohVicN9vdnblsgj6llRt4DsNzgqLcyqeet1uPqwg6fT0R9efaMPuT
y2n8eCQh8/2ZMHixL6r6Flxy8rX2oSF8cj7vRLbONNaS3m91ilRl4d5o4qfyVv15
Vs2Px/58XizYPecjESZq5rLGctVdZHfryzhK2vGiGKBjugbvctld2yAUvkpwivGK
0e7ZWWbEbQBNFKsHqj0Q+VJuaGm2XiJpnG+LVA1nDwUtcgwWY5BOWw1n68WrzET3
wFio1yC/yFfhb87zBVz624c+WKCSbBlvvlgJYDPO5F9ctIxD1W5FBGxGNc57Jt0Q
9/+GJGUo2ozoBmwu9gqaCBHIX17RSW/ZKd7WexxwvYUUBi3mTr82WLPPWtGV0mZo
6hSjrinA6isadOaVdjhFUhNs4JYhKKqu/h3Def4gVBxW4SLGnHvTdcLis01puop0
qvZySXA6DARwrIxAUFFDO0bCSdVVVh1io+JChHugH/InRJjlC88w1Um1Zm215mBJ
KIzEYlmwCELsmVBigaptk2Vmc3MHGke7zk6ZpUYGskRALRKUDynH5EYUSC5eTjUL
pYksKBQ9vUyIv+HiyuUs5RJYNzBEaCITsjNMt6hfDVShPrnw2O/4/fZQbzhnHttb
SMafl+KxWKIYj6KWCCio+nRl99hZL5GZz0CHHXwA1yf2vdo9dT0Z2zr780Ty6d0R
7WSs6t6TPQBdb6i5sylYdM6BJOMS+iP0UJd8GLUCY2cH0jNXGfqR5MgXjFSLYMaN
kfGsBUiibbZ4bxHrGLT7mqdoFXylDm1tDhI4uNqKcLEQRR1vHVobysu8xNCyJVqc
OJ/6owu8TdovmIP+YIqfkKY03+XJSiSRWMLYtP3rwLpZRc+D7TeAxb7tjmkJbIJA
BTCdYgpvV80Q9RqFzUmzbKPNRJ8PV01uLxeHoXT4ils=
`protect END_PROTECTED
