`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pW9eZQtorba+RXkZ99LWr+QNF9NABYcNyQSbjz242VtlGzxojBp6hinyeZQZhnmh
WgZu+9OhwJ9YJov0oWd4Weaua+3FMVgqk8C7l89por9qz35K/qA/UN50wnyNDXby
CJ64tKLAJZwxfyWrXGzvoJLiXe/LeqtBSGHU2j5znV/NtqIear+P0tUhFsXDtie+
gdvo7bW5Jr5bWgt+Vnsbr8/u1guE3udVjyJYeIJV1JRAgXIZr2c21w2O5URIj0dh
kxbh9/L9peRXx5MyuclkCPVcMf6U+55f9KRGR3cn7DCpS9S1DfqEFaaYtT1yQWEw
va6vhmLys6zJGRfwqPEGWFFRENWzph2pPOAe6jrTVbh6TJqtV9Vhljmci3xq8zNg
05qvCgLTcTX0zLsU7790Zf570vPyEwTUR+WTOxOif9k=
`protect END_PROTECTED
