`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Rpy+PxQYTbLScCiBE/wr7gC9RB2yoHg/kFe4xiXToXuFQEoeSDTU6adl1Emniut
/wjyqf7Om1C28A5s6vuPYrFmEqqAahu141moJ45F8OqM0upJ4hw7iwiYKurtIhbt
wFnnf71eGqMpYfjfheH9s6TfQFt+4adnix8/skmBfk3/wiThMeY74iNDHs7e0sQf
BRmbuvyibPfT8sojcjltqKEYy8fHwkQ8UuRA/Md1SbKui4vN4xkMEfncosnY0LC0
qQnqzv2KUCgtvjcnfNJ5LC/j1j/yjOUnbIVufjnC7MxxoZ3OWD75xlF+M7wCTvDS
CtaxN8ckYv9GgKOmBFUJ6xP2++OVRNO2p8gifPP/Ap3WhJI5Z9JZACoVnUFFD8y9
TpwY7TpO5k0UUFXJ/Gg5kDCS6mGvRn/dMhMaQVbwgFWEKK1LnVFZgEf+XSjxKQnn
HhpHvusmzMVl5zNYrESiuzIwfwaAHGbKLQEjjR4OWP+OrGfqUFuLN3LfZFpx39MN
ywlrssZiICtsG8lOUx9/NKSChaFbD/9cON2Agy6QxcJhSii/1SFapePzL+jnyTVV
qSmjaSLkgdM6Jr7mYpQanWF3PQIqzrO6f613kjKiItT3BMkrzby8hpJyGu1GBgme
nuQIZf0b5dR08MsGXxhgIapcHN5QZonLT74bhiXkUqIxOXthyh0fhF8KBd92P/Lz
lJB/ZSZ099tRet+VpcMZIZBgCXYlfB+iCZf9BRqa0pVaHEt81i5IyY8e9zmLx837
r9kgEvjeC78NL272BmuubF5VDmhI0FktblEMalFO6cWFIoPRshvaj/kRmILnYBhl
VXenM/GqZwIx0uiVtbrFJGrwKyjpXh7vM77A9VvImg1+mEboRswJe3WXj0+PHp12
ln3JRTOZWCUCDyfXPlhgfBiYON99t1hWwGiCR3M7z9uy71LXuitTfJnsCWhicBxT
Q1k9dV923jWZEw2q2sTVGfTVoRMokvy8o20eWrOow9eyrkiIGycHcH4yXzWaQvj7
PODn59ldf50hKacb03OwfYTKX2TKzNa6taTCYCLV0Qt/5fVcB+1FdM32WjnBfzmL
sD+0kb8qsdU7A/G08HuDXxYdc5JqHkxtwLLt2w7TIgQ6XVPPhlJi+zqyfrSI4EDf
mDevRjT8gcDsfpEPYXzqWtniviz3Hx45iJly5zDLjI6jgMMqk2X1HhkkUOtkVzZ0
D/A7nTBu5vRe7GAbll1CYQ1f4v9qy8UxIrLB6prZVUUUsHIW9ePxoC9ggTjwUV8e
`protect END_PROTECTED
