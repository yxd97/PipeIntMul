`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pu5tXMGyY6/S8ALpoO+n334ESr3MO4C22BFL7A2Zdw/a25dTKMKYvvoZuEdBcHX5
qNp8Cw0V+9B5ucUM3JXW28VD5XO8hSA4MBVBEY9fIlhtM2s3pdmGyULUVKtBEchr
On5ZB8h0KpMVJtYEAv+aJXweMWbGyzmROHas5Z2e6lQ8TnaBH1T1yeDFrFvk3r6H
vSzNXqjAShRacaVmD1XmMmjnaF8phNzEhx6CfyyxxZOSQuvTGjJ6gmUhKn8pM/AZ
DyVX9HAl7RrRmapLGDGqxW/nfKHmVJJ5QwBQQ1bh6XrsLVUMFztHvG0OFkr6AOSf
9jwHKi6SJKG/oUtFEiiBrbIGftngbKhkLksxe2/uzhFTd1ttPtrKHquhmtXvmXBC
7Y0WcQMxhx7EB8SY58xY30XH8/1DIUEEl4fIRqFlhO6pnMMC8BdTEmZqJKrckcEa
Krr5lFwrVCKHz0a9JIP2HXFZ/l6pMBt/m8xAl4N19iE48mgDVXUTeqahz8n4UTmd
`protect END_PROTECTED
