`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UahsGaXwcrxg5wFEdUvnkbnS+2B3SNXZ2j7h4q3Wf3hSF5cQk18SysA7ZVN3VHTn
KKyac7jE+gTwv0hjsi5W1lnyb+vYmfDI8NQynH/DJm5n715XuhxA/S66Lpu7mylI
J5P8U43rbWTv2qgxyQpEfdgrse1+mQCro9HhB+YvjVIhevYSoxr5ymLzu9GUU6xs
h/rtsV7hHwLwoWe9CK5UogvmSIH0WG51GlvDOug14ttVQX6mTkLY07oRQoAZJsbT
N9t0uYogPeTQlgjYNpBfUbQj6DIL/Q0zOSa/wEhcROdSnfDKTLNFN7799vplE7Dc
OUyvMCHkiZm5OGm6jL6J2pptNpnzIWj8iYG193EOuU8aRsB2PPrfj7e+UiyFBo+X
lY5qaAOulmxzAFFRJBsBmb95lGoP3e+9qlLWjLv494NmsuUzjSh0gGhkMz2GBtfc
MIGjxf4iD1eaHkOXO7SkrxQ6z5aR5sxSSFsDW2u8hAa6AN6/B60sMC+KKiUsY0pU
ZfvQ+Y9o+4bBNlxMBvWMWWUwMEy2Yg74tj4cWSKh8r/ybapVePHlYb3k8VIJgp5J
RooC6fhCV3KXHG1aJC3pMCUV0DPKPRbdJIpNOymr1pmCuCFlj8jOOb+6TCNPFj/v
LyFWwt1MXE6go8V7aC1vZclzy9COsE4xwavAWvwuru0=
`protect END_PROTECTED
