`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EmcxmdeSshWPKaL+quvMuU6WoDLTO7BKJRMPY39Gzyklao12diGWNn+M5PvIUaJg
iBEtccAZJku4dtWmHte5lX1Kk9nKp77dpszxgcjcbz3+NS5V4VyEeVQ7nZ1ghNVE
+J4AbpM6xnuqFhifAolOEsBdqOAxr9D5eoMoBArjFvSvbXYK1bkSuLvZh0+iJqoq
MxkPNfs2oDUGEpwA3/xDimbFjYuQV0gjPJdgCM172ZctQpTB/3Osnu/ln+OrS/kR
TbMS+fMRNeaCqWgaQrPc4fS3WamM2W9Jd0EI5eT7HTVVAFYzd+TAGMncSDu7ctoP
sZqSORfPxut9PoOdUrKw7A==
`protect END_PROTECTED
