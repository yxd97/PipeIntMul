`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rOA5+jGfRmgGSXJFQQsAX0KW6KZrbdL3Gz7TqopoYEDklT+y+TOdGJCeVWcN8DqX
V0fgOeZ/HhHAlAqHpC6cKvbcjRX8TT0FniKj9QZMayfOEZ5HASEPEO929k7BJKuj
81OMIUyNtFR3aqMjgpVPHqFIcWTXMt9tCjUWr2rZbFkum4PRct1/BdmapSrTV+M2
cv/FN9pHlNlL8NZgUqqmH/LOYtDLV78m52k7YoBEo+G1dQPcWKZ/U5Fpu3hi30Mt
ay051bNlQySyRNdVmjEio6ZpGmLva5gjGdEPpU2YrPAnt90wLrUp4BxgsLCgLXAl
nnYqIlhyxNFXGzeqHLllMcnGp0FJ8vppTKT1/tI4Y6V4alWN30QONe9mrODmDebF
a1/GDs1hpUZ6SR0JC94EHbl3iSZvYYGp4kidg3Gf6HOXy5nOVZguyYeT6LXU6/yh
sswy3u541G1yWUDz3XR3maiARmOjh50AbooQ/EIZR/w1zFQIjdGkbsqJh31g/hIl
oY7uHYrzmqDNUSs3l7M2DsnAfM7gbNVIgtPGzoEmwBqEtGAwaDOnyzyc+r6mabLi
0SZFZihqlJiHbLnSmhH+9859ZnpnN4eahzZKGlYTACzrEzhQvw4yd85gi4Xq01Pt
B7mri0FVdxtGctLM+AfnmqTpN9xypkQ4/6nAt5kOI5GKvZx4EFcO5gtYxj18wyU4
jkai2aP7Zp8ZLxN2ZaT+VxZ5DAkC3YJd8+TWzoyvfgvzUqNMRuKljUz+91lFo95D
LvPXpQ0VTxHW45BlSKSkRcMEqIzMYhNCV2Y/uqCS2nE=
`protect END_PROTECTED
