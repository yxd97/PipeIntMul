`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEgo/nx84DRBLyFpoT6mKbHe5CZyJOMfg85o/d9zacHtEaDvfthRkmHz20lZydhJ
jI/qGwbfEDPfzPeP8MSEHyWBHaKRHREWcONyGT1S4PCDyEEkUknnZj3CQB7MSMzt
D/o1ZOzCCzyMJLaGA2YfnqoJVmTMp5/932N+RfFCCcHQxfWO8+siHfgUGaaJCxOv
K/QDYCVSXaf60QRpiaWQA7yFimr+NKqDmTTXFmvx9jJBwrlxstcIS2lkl8gjIhwc
27LaKnPcE4e0H46i1Gt4zpR25WMl3AzXQX6pIaSSglSS2dEt55LR60yLGvgFuSOt
94LRUXL+GamVhknY5DU7KqlXpA9Of83FNVAQI4e4wYkpvryN7VDOq1w3mhzPgIsK
Gyfdy/y+ND/eity0fBS6m/4hqpgKkCZIaZN09VF/nUsZRk0JmoS38ADj7oA3haS7
qWJBqdFLot8J69lx7qQiq2mg8iET1nN5TQn7lAfd+OlW1WyMJolL2+6DMKwSj/xa
EMZqxNHymlEANkeSgFdJapYSrp6pngd19CPUug4/Gp8=
`protect END_PROTECTED
