`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xGzKkELofQLnZ27TgTtmNQy7T+8W8l/HbeOLTP5CXpu4dJrxg2Dm7TecZ1bgk++8
tAVrZLvjtLxzwBS/n7XpM4qX72Rg5YcyEcB8ICP4SBUzKVUnV3/o4m2fr6DyE26C
zZivwM++QvCcsQbB2+UXVoSjsM257Np1vLMr5ehgIGszqnLyfFfpkqIiVI8gsiaJ
xvekKg9o9g1cAUbsudihMOXF7aB6I8fBPRwk3Hti4JmBBpHWqANk3JC0A5v1pnfN
NWFmvpULELrJ1FPbZKEKiaN9DfkpIdal34AMtDImZquqY7KAvRgyzQqMGLE/YHEA
FHU17fR3Nxp+wrlD36YS8fe4VC+s7dHqpSJo4hd9gnM9JzzM//aide50Gj7w6y0Z
q/P5YSx8OTGML5NTDxfmh1ijDbX7TKQTlkWRuZBMGEp+qCcW6YBuG1oihTxV/H0b
RnmnF7gr94Kmn9mLb/HxN3CkJMPtIm7NBWQCfGMRLrPiPaXJQt1lUVMyv7PW5BD5
EbdKZDRKbwfoH7A4MQGkSY5StyA5L1LVORWibUMUbe+hyTaw4X3xkUupjyc7ggF8
cvTpYXt0hNq3GD7c9M1cVZg+SkE8eFJH7x0PLF+O6C1+Sgh9nJytkijfD7MC6Kv7
6lkJkK/wjqPyXe9qlT7zIa5bDYWZ8cBHWCVgCnMd+Lq3vzox+1pIY1ngmn/0hKpV
UZb8Qi/4uxRPQUMuCL7Dkwg1I5NjvkfICgrxD5YSuF5WO685mYkq2keFsA7cDaaU
r/9UmtzZZ0ctB3bCOFX1d3DobbtJywpluO+SbbI+oYTzNzKgdAh4hZxDLiEAMQfy
Swp9Y5MRFWRCTOXzptjEFugCxIl4fB7eHKMKfWASPMCtbmfFdataYZvxc5DVlHC1
JkvT99tfsRnARAI7RUqjoJHwxU6pFnDUvJYHiYxUK+R4hhqGwTBjutPmVCOwv2O5
`protect END_PROTECTED
