`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qexbRf0V2zysptMnaemu/+biINJhyJ0fXsLd1Kh48fExIiQb9my7EuYpxPNgmvLK
ICZOtYrEg5ybvU8FYPr6+mzqDHQMj4gTMCRm/FJ7a/bBQkECAkaKw8iWrvSQRp3N
0QU7ajjxsM2c3Z5mB+wcaeCylKbZSkHLCDpzb8iKZZNE3N6rPCNdAhVORgltt9au
sCzW/ymWCqqpNul/KfxejP6AEv78PodSYbWWnjt9mAU69of/R5CrTEtd8AX8XO+F
wYbnpIXV7Zfvd+8Ho0NLEhmHAfVXKjA+6GUP5WKJlGwYuCHuMrKvD+W6V+FsNoGV
pNBvWA3DFkRhYJTrJY/BhKYSbkOQswTSg5vVvOhk7HBcL2f842ZXgzpgwDC5s9Br
ldv/B/rIT54Pg2bYEJy8rM8YqCPQ53vx6hVvxL/6AB72jkYyn+6cw1/ugVgZimHX
d/ZMJqkO5/5ecjXnkCV7Tvl0Yu0aVefQ95wDemaIDbGYVa6YhqL51E9pZ48okaNI
iXMaPKhVg/d3DgsQ0sx/CO+rOrMMyhjXhVeJh1nry56fAGQefTQUVBibcuKf28jm
jNNMQ50+ACx1pYdFvqDotQBDveRI6gSytWyeQd0AsqUXXpWpuwaq7jGzBKiDL1VH
hDaJV+FqtvE562xDjLuHWfPEVZuH1JSZgOSTVbU49R2r4H29Bn40aq4ybnCNBj0o
+g8W1KjV/yKJLihw5z9ducCw4535T0ltiqzOjnYZyzcjCCZkd+F0tC5ZHnN1UVC8
2gVNlZUy+seyMBtzOp2IKQfL1+kCyP5tcV05cyqA7rhQgJ/W6XF9VZgNtu84ac44
F5sZ18hP/CoQtlg0m+n1E/T0D7kSIKr5bZKJTcBJpr4ep0iyKflM7TP1DhNiRVtg
tOEzIyRDQHSpflmEpm6yd+FhEtqxUqi9TNu/G4zDk5pjldjkue4hRsc5y/XrB+x1
B9Jf78q7QX9lAC/E70k2W+ySPYafVY+sIj0xcS5VyfuJUaZc4n1FCQ928ZtBgQc3
rz4xHNdadg9pXc8/OOzjwZTJBkMwRV9OTxa74qU8IJGAq2Ttv4nftE9BG3si/d7Q
JXSQWqBlIBlKzp7uYd3IsmP+yQvHnnpIoc/S500NYG5NjF/RdeG/r2G0eLojBhZL
+8hs1KHcw76nWOybwNHXrI48D0aObZhh3Xw/tuFOHy/oXI2P5aToLJB0WxVKWBOm
3Epi7ZQjTZywm2RTKWv8ihJl405q1zZjj/rmAlMxRB7j0SHYiu60X9EXKsNTvchj
CD2He+0avvv+E+ZsA2sm7ZHC6M51uInkFdF3F5vKVyfky/LK/fpOOx7dx6snZm6N
YTUqH2AHWrb462IzhNwTVEH82FVnSx9bXad+Ob1m6Zvh+lOCIFF7PmtxiGkIMeR/
tvUNvFcycrakRV7YT1TqvVlj1jSTyDd14V40xbUlafB9iNeSsb7TaOKV8EhwwoY8
9Ev9zZyV5/yYhjG5r/4r+MUpxPQ28peWlJYZgTsga8BPjAm4bGmoowY3q/2qIsnn
LOtpeOB3KWsxT3Sb9XBUciUdbyzbMt4aONl+f+XIv81m97bgvq6xoIQpUjwtYTYG
aAp7Lm3/TrMj+YchR+JT214lxGmg1LlO/OPINQ4zNGu/BM0KXkXPsu/xLvDUB/SV
XUneqEKNvHwCW9+vPlgJqmpBA2ZPps8SyChB3OBvrAN+OVUqSk1+iebXuvmMX+Et
PntaIiXteUmLweXAm+uYIjV7yIZWLCSsCWvr9G87MyiDIlTYut8qD4Zfm6PSTPsV
Dl3DgxfZgZyc0kiOqfnuKVQWv0NcPl02r5N25kf9UqfJ1ckuhSIuPY2MPyIa0Akt
nKu7YBRPtbCWbRrRuBrH8Ya6wiuYVvY/GI4iqm7mH8cSo8NOJqEtn736orQ54z4o
ZH+th3FhbJInEIb6BejF1Rdjg6/mDsTUwKYt9Ljt5vekexueveMX1ZIeY9r0EckJ
HopYLsRSIVnk5VrbxrKU08UmHS9AMdioieyIL6yqAZy+afcNroiVurxMAZPa1gcL
6tj52HAPr/ly9WtRrr+GifZCm8ALQ/RrM04ZGE6XFWXO76C2yt5suYwpLcqJt0fE
BuPtND9DTIazv5iHVe3RWyQ7So7f2dH1U0eEavsTeP+o4nQ1uPsSullDfb1BAjy5
71OEk2/kWqB+3QvbWk8oTMBpIVoahuq0qhMxGwlFtM5qVBo7zFHMqhmrsoOUmyUE
8/Cg73O+OyLiby9ghjDz07NFxoxhTbPuLu62mesQf0gbZ+cwDIqUuOa6gs80O/Fc
adaH08hdvECEmjpM98j4juLSh208EYBm1dqCRoF46WnUkMkyFzqba6eMo7isGGEp
CzcTH/Cp3yTC9aP7sBz3kezPKNh6ltImpf/mTNNiFZ7POsoiQNAsbQSHGQACHO7R
UKTnP+7BDMQOzjawddnxjxyrnMPpPfBCXsvwtabVOTqRmpFiSsrITX1+LtVOJSfs
6IQ9tQGug5Ga/+IffRJcZCJd9Ux1cLF442EC6fvve+6l3BGPUu8Qbsh7PyfqzR2r
A0PYRuekE/e8CnIBR18Emn61txNCbvYoxWRRmFBL3V1B+afzj08pDquudKnPqDPR
daBJweICxSBgsQxMS4dyuOB+hQeqfKfMC2rqhjiboP337zKJp5MazI2KpVJwWIGv
AuLlyKxGrhtRtYG/wg3TBsH9edfED23/P2yoeR5sUSZ00GSQz+eOXGuYDIYhNM+h
Ng0mBl464siDjHCyRQlXUovfECFMFQzh9v/6XkSlETWvl83C1jFD0/U9sNHOdqsm
N2BZRPFhJfqd8NtEibLCxR6eWii1ypSh95HQHI8vh7Y35CQTb4nuulg2SamgjQ5k
8Gr1LHTgrKXaprLSbHHguUhWxmdSHiJStflfLm9A+FAgp0/ANtTtFBtwDnEvz962
gfTpXoZLfCztpcxB1Z25l0JPocfW1WGwMEG3dduSjXo2zJictwx0M0mC0JidyV6h
PIiWicGspY3yGFuniTlafNnxazjnXQgGT4BPNtqpO1G5UjabaprHwB7aBKeZeC1f
lf1zzNByb3/a6r3WP7Nf5Mb/e2NwH2tjjN6+JuG+zdue042DuS5AY64UQlT7S2Va
B41xSLDGARIXWfRP6guJGNyWPIr3UBTY580tErQPNv1DkwJqAf9H+1sMkDoPZ44h
uONzKj9YIWaqG9dqAUz+3c6ibldnJz6yQuVj+l909VwzOpiBk/946LpQOJNczGIe
UldSYG836UXuSM2+ZXsgi/7JziNzs64Yvn4eSXzRKrCTHY9qxp1pPcnekOhSP4Wh
T3tUQYEentch/tTjg3g2/f5fDRaOK6Tr9dMcm26MOq/nLyJNzsDQnFrACiqeI4en
WFwQ+60cHZ2UkEuteSRqB+ig0wkuCm1rkmBvPHZBdRV9Q+aYWb5EHKpRQzDAwQ8B
sHwOIT3A5BfoXtyidhByq9vYX9VBk0IMLhXFLwQ27mX8M+wX1rLiuwpDXjWqAJAA
i4kcqTerRH7r4QJud4c6ReSOyA7Fv6lOrb5EYL3GVZqLGJqRzpYWvuoinXapsybC
dDq9kHTtvtuE2kp5nxS5vOFDP+4jiXxW5kxaajWhEx33tSqSXySWOGxb+/UEaL8/
LW2Aj98zvAUTCl14ZYF3jdSw2cnzs5Wn+fpDetyLYZ3JUdIUN3IovemGn7PRxact
mufEPB7Xm76FtiW/tR+d9vfpE/5IeZ4gI3e0OpZdj4ot34P1g1HsEOK6hfxxYKcr
XEfgHEm9FjPde7YwVC4FIOt0fVIcL/JkmHNquzz9n7qe4zrPRov/lupf+ziJRnSY
BhvxncAeGk5e6VdCpwrcAvw5XHYOLsUIIJttn5c7wUY=
`protect END_PROTECTED
