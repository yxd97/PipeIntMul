`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eD9uXX8/VXeLTn6AUZI3pPPrpjT/zb+6p551xs8eSTDvA7Ozrcqv2xjDP7ofTnc4
UCTIwTRZeAPUNULSOFm63qgV7q3HVxWsJek9vniQUkMSLqq31peS0mT41lwNAvEV
3pcRk17k9IfY5TYkKJCboP1LOuQj11jBTkL+RT0yWrXC7/2Scql10dwlMbRtd0Tp
StufGA/8ghtSVjLK4xtw5IiycFCcUFKmPzBR8fAm4yY7CltG3J5LbzobkZvu2llr
N19uTLVzubU1zZvPnNwqH4ti1AIuAhanpCpOo7+TfK4TRvrUODfFlVsXwJMnlANo
2eA5KNcJ1BJgbPPpzjGfrwSmt+5D1edrvDZGZ5rbfufQhE67RtuqYhMaQb+9zaEq
MDRvgu1RC1cE5+4jCBhkkx9HhzpCQhpmGftoOeXpbYk/3LGLLSas6t4PcO6QgRvf
3gNGQ/6xCmYV2evj6bM7sAsQp9EScAoNMRYYpmUsBTsLdOr52kSZrfOMxKpj2aJ3
K49ks25L+oCwH9UlEAE14a4HV3pXJelF0SlVWxCt/PXwMuv4oQUUTnORy7BYkBWY
oyciqzgMdX11+enPrl9TPPPNywIuOdnXpUbHNgXQwRdtobdwR05DN2Fe9zYupUDn
pwEXopn2jTB5SMwy3nq4vCu5vHvEHdsCeSKc+8lWayRI5msQHsg/sWCglCtBiIdS
GKzFBFUjtjnN/+LODSp8iBwl11j8c+9GHl1/jG/poWZm7frIW5+l/6QBN4AWZFme
QZOSg1eGq2JIvny8tHQv/rCgmU0h3MXHYrYM0x5TrqZgrPVvUHEvSDzNFDlR21RH
JGdhup86Rxv8IsiCW5S+ojpdPZQCA2/woviCZls8S/qrlQCDKBSt7Lv75wBwBzfk
HJIu8Kz8u6xeyfyYC/6xFTNnn9EFVluzxbMYY7BlHflUFUW3gGTXs4xWbwPZZcB+
AUkVQ9R9/9y1QReCOF61uTmNY3x2o732kbkmj0314tGSJE1b7J+RVYWQh2ryn36S
wzyRuSsllzNUtzxANbPkoXo6FOWUNs6X/eoQc2feLWum6+ENjvO/FJmH8nxIq/dq
Rz4OGzoxxjvhDIKHpgFlYHabqGlZMIguBgw67qccScweCY5lwUhJxV+5iXtz1nbg
0b2Od+2/YJFz36tiRz2iiWys7jA1H2AeZb5bstDIE2zdffdLH2cM1qSH2rAczsSL
ExL4Il3EB7SZ+qPbP3kRbLC5NBdCvxCDJwJ6Sll+GyTOwV5j2BKZfQOvvXvA5B7O
3FyNjueyy3ToHX4SY02BLMXTZs8QyH/XjA+GR2PBe++lrHCKohjwHv1hfRl51hve
PqGqUwIo9U68Dflt48JpAEAs90dy+EgSuBcQyD1udnTCzvaNX1bMbcbDdIz4I19i
tKeB9EvqUaIIHt61ISZUQ9K7nE9RU+i/NOji0PoUUymkh0/ct6sAnQ7NqR4xjfJj
Q8Zp2+ZVWQ8cNqtgwMFpooexTTNTuomlLwJlobaUDa75BxDgjSHc+WujTLvbZQW9
UZWtxtJdfxvSsN23CAx7Z2LzsYn4iqG4Ycw0R4oiovrW/gyZOZh4sn1/HDVRTPPf
6Cm1beuyt19DJZB/38Fqscc5HAarA5XH9g8g7JVuayYhbd5K7JzfWV1RgM0ID2VN
x7OmIaBgrcEJtuajEjwnL/4KcgzmaamVNiDEXl55blxxlEfhA/8xrNgEROwEOe52
BB4InTvXQbhN11YexATHDXwYEG1bxFrB9/QpCVX15HGJnoFFwq7kmiL+y9cq0kQP
u38hSEUoJtFifzS9uZKRSybRv2ypZOFn4j4f7ucM0jloI0oUsV7fbn1rONumJ4M2
VywbDYYkGPNv2kvtK5+VzTCyrW7LXBDe70PRReUy4eo=
`protect END_PROTECTED
