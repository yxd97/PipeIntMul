`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KOXhFeQuOyaim8aJ+DgwRWQTmznAdJiUAITmqHuEdK829FOcyC7Nr8CO0cDvBFk1
CK0t5UFvCWHMopf3ipXjG81ipQFNxGMLp7KG9eSUDWrrLqJgBCVTojdWvaGnPsXZ
eZXbo3a3qFIr1h+4oyvdeVLJhBE29Ar5lIU52C//kmIQ3K4C5GWlkXTxr3iNV8EK
DwunYUuqZ6YvfYz5uiFIpj80PhCdyiYitpNnGEm6CBGUO+f/+7+z7c2Gnymi2ymo
+c5017Px6saxqUDulROyO6c2SYhJ6OvaCUYa1njp+MNk+o11baJKQSj5yU/pemH7
rQDuIEuuZyLPXw3ahevO2vcZK0jpHJ8uZZzg17FmQahk9VYcowarY4wI3NTEDH0z
UQ7+8YGwzF0DCc1RHyW9rVDmPa8CCOo5HvY8X8ATtOnAP7xvuJEiQYwfJO4RhVq7
VLqVgd6YQHnHd4KAezErnGyBVpBw4q2tm89udluMrD/vd/kmeZPG+32qxRyqWK7C
4O3usDG64q5xRZcaBNLckWrpQyL6m1lFVUeyQnEIMp7M+FjTj37ekQG4qcjdk2mN
DRrRIyrHza9OYiCgG8gVa9fLnr1AJRX65GCimAsGqfU5JQ4uS8/bY4DDxYt2ay2Y
4lSe6s8vNSbO+qmSnkOkcZfRMIfWx5jHhVrga4i3ciuT34mYyiw5X/O05sf8NNMm
wVLLYY95iadqz99+l1n/uG+ltUQM6tWLyHJX4EPijtqfVEXabFEDcoVvQM1BrEBz
N0sXgsFKgQs9yeiV7Msn8aIr+7ha5VzOIJCKm9+fMOvm8NMR0j++n3EZHAX4sQdP
3xCQLmzhbKhWoouXNObK16BoYTXwutTNvbhUkevcy/9DlnzbUkWS3KThgI3z7u8J
agU/m+qQfIZCYjlO8gcOAujWqfXT4ZilopxyIhdSxtjRo2qXxxVy9AdKz/e2z0Yj
`protect END_PROTECTED
