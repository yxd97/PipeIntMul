`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lbt+5fHO8DtFk4X+td08R60KKN9lOBViZgkSn9tUEX6dZZEr7rSSWhrw3xfap13g
pnoyt0iOPu1xd/avkvicKibsH13iwn0QcYl7rpfXOJF96zlWRt70qa4bIQh3axfl
0Zm1aCNo+zsrdU8YaUjU7bEduRAexbVQ+tgGRYDFbQkq1G1OdtPbWiMNOJzenrwy
/6fbEq2D1iI4djdllomLDiGvmcHYt1xRDoZtgvKNxfWNNaBY6Tq1OAiktvnXLdB3
xQTTqum8k8Nhftv0zbhGExYF9psEqbTlYHSZuTY0rdiu135Lfw6tSEmKGM6MKTJF
Z47+Y1GdFkWkpUht5O//9pH7HntjR3Ipo7l/ctcHU5YlXHtGTUNkSsZ8oUbm1KW/
Az7sBX3CCjbSeMRiIwX073phARrywz7PYADH1uxslwESdhPJ86KZzCwn2xAWMXmQ
smmIMhFMlCsYlg5zyTTRXjsRW/XSm83xk+JBgeHzW7bgMaT/NDCMJ6f2eubUw9Np
adV34xWkLdIyv5oaLjJelm1AU88DvUpCu7pptv9oTfgBxLdzBL9S50GBK4RzPBKO
63/DIcsWmMhwuW1lIAnarNK5n7/++O42i45LzA1CuSIXZETTrMn/GxlSSjgDWgj6
qu8jsHmv7HQzyV71Tx8WJmuPXVH1QB/6Qj3YR7Ln1nZx6PcamJqgBA+svGSZPNZ7
s5u8vgbibpjQHTqiOH3ajA==
`protect END_PROTECTED
