`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3nUc070T+M9N9hMZiXn7tmTuc0cGYG8jmtJKFcSvlRDFi8dgQArgxbb8RHIYCVXR
MtVpqxfLVhTfaJzz3E+VrDe8Y86f5TCkchbkSGIqiJbXma8PiGxtMbM2hjAxnNe6
aXEYfd02qU5uRtyZrc+rWagyIzH+Lgzlt2NMO3YNftmHQGlfrcYPu7Me7HE0brXY
tyQq5dScElm4hKdhlQ854thd1EXYGWtIjcMTF4uy87ij9AOPAi+2V1KB2n1CetO1
vfP0tG4N526Wu9pV2vg50w89ivO1TeEpEgO9HnBevVg/U04to/Mc3txrCBE4gAUu
/vr+0v64qTHSwrtzvSf/70Lif9/RZFxo8wXp23KRNyaNCUGn+QRRcbvDZYLtLD6b
Ra6p7PM0rt9EllVGN7YO3nOUumt+JeBRNGVUD1EIB6k=
`protect END_PROTECTED
