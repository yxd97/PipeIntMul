`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTFeX5DWI0ZiAbl6rZ0IAIJh/EKPHztEwAq99st18G7dBJQ6ofMClvuzN5g3AP8J
zRyBBOJJdJASd0ThiNudwSKxaOF3O16NVVzB3uGxN2dtWzky71g7SWyZBNOKjd1k
jAqoMvsVxdpB/rDiBAd2jvBYazU9muI+uLPy18+Q1rTmXcflA8u4t+0QTg1P5xyk
yaGTJwO3e+02NHNmB0PLPqNKZgfnqseuW0GHK4KAKF2m9KgdFhVn/7FkYfE6AsNl
Q/j188PbKXYt08i7Y4hrN7VCPAEhdHtQsF5jF8Z2hpY40r36qL+MuIgvYpxB0XVe
BvPb6sAz1+kmZO4D97yQRFgyNWkLQw4sLoIKZ7dAPiwdlffMdIg4RuxOA588s22b
yKU0zjQl7s7ReX3I0xxjchtfdFEEWHzakdnqLbtdyiNmlOLIPY5Z2R1PL+iKtpyY
/DZZq2m/eXZ8X7LB1xgJ8O/Yt307bs78irBvjC19MeEzhN0BHAUSAy41JcoiZJax
tiipAaq4NPDDGpMRyhKCRbbl39rs8Yri5ufEY/cxup8=
`protect END_PROTECTED
