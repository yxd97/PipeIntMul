`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pApfNVxTp1XB5zDcU14GhH05kAh06yiWez2MIOIULs0EslL2xgCG3cb+JcmnEOHa
nr5AzYEFDt+Nu+oL+PLQ9d3VPZgmLVTaKYFfJglomRuc2YRKPMmU2bDqR9WXiAcj
mdgjRp9SRVo0V1wLmB0eTNkNZQ2et42hTfkk8xe6hBgO87G2djyMVswQFU5a5e3l
Fwa0XX+qyFtqWp0kJJm3pr35EU2ntw52aTmbuYuzGzPxQPlnq8xlsnXHa4NNGZwJ
iX4Io+X+/5krUlzzUUqXhNacjZnEBL1o4YK/WjQ9hl1dZPSXn+EyPKeJtwTnV+rS
WJboEQIpAtNjVjIT81NoHbeZQcZ6yWFKy6oxah7x2uDOh4EyqObTStQXrsJP2CKU
hA3v4SkattzTV3nvUx7/XiUAjyU1sotyDCtmKL5sWz2/jYxmkhSzboLqV5uBZcdE
s/+oLw4KnZMX2t3NSUwIjw==
`protect END_PROTECTED
