`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pPolfvqkKzESGQNTvQYkUx5xjD1MeuyZ5Se77iRMZhaCRCQ6GvqNGLNnKlZR8Y9m
VeJzr/j/0CQNioMW87OlUoW9pNBNqiQ8sexJEqV4N7uGarGY7cf5+XZFHOh/yzva
xN2aBNciLwuRw1InnnEVUw0qkGlr8deR8z4xKBqzVohFnGiBWmvEvMe1bn0r8kAx
mUeni2PPu9rgOnDr+uKgE3nmBPwcvj7KPBQrer81cVpKR1RZuD0uI+t3AIOiq8mP
t7/z5M1CaNTxr0aeCt6ZyaDilG91Hlz9AMzbmh2Zdv9yaj1T1jPAV4F2iDq2m+//
5A8z345bl5KNAZsyEY4xdnkaiOhUuAFLLz18lLxH0uKJKNGHkzvIO7OCcgcFSlx7
`protect END_PROTECTED
