`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hafJGBYIOJk86tdmatBeJxQ87vYaRyGO3SEUKEL76UyTQLdGHnmpc+B/dG2qW4U
zlUM4dy8Xh9OSaAogSXiprwAHsbcUHVwne7bO0UFbBGIWDotLcZGvTXJ3zYBJMe9
uzp4LNnnxbeDCS6v99+gZJmvs05WAWPbmgN7H6igYvbCUNJ9yLOtOIF8VlFVvlwA
3VL4YSAHjCib8msVCjq7Mke7/rw4a55WWXSkzQdhxKNnk99o1vcLDgMPBr9cmrlA
h/FokHMOUqNf1ZRsklvWSiJLWtavab4C5fXHdXGz/gTacc7oFbL2OcOoq6vVRLt0
CZvUHXIefF6w/mBvrPxbyzSb7clmfx3KnbxRYUJrfgbNRO4sc0tb+u81kHn/GCCh
JW3ThrM3uJsusRbvZqsLefRpv6Abnty17ZR4sa6jGN4XFq2qevgv2a5zkMaWjF7O
pURKQeA7cr66deA8N6U1UUJnkHKSoJKZYLoff1krOPkcJmAnMzLcFSK3ONwJ/Ey8
1D6v3RYnCeriewiTMnECSI4blzT7cK6B5gQs4ic5knk=
`protect END_PROTECTED
