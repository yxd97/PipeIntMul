`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tniX5p7OOHmWhusiUWOx3hBlxzue7CN3GFWm2BcZlPBQRtdBugMCIIl4RqPA9jE/
vpj+XZAnYqEVghL8ZpQFRgIAe3L1XL+v6PsRkueSCIjdYY5fWCml75LpnqQuoCnz
LpSeXI0UkQBu3QW+g2+qkmp8ufqkwz/XtD8SvUQI2yzuf0N5diVg7e/AVUZmAbj3
Dqsuvn3480O/szV/OzSIO4qy7uj7hGQOIH7lCdH+IG9yyUaz+aXgljqvK+Siqv9R
xOm5zkFjqviVwss97pHXcztZW7XJZ2fmmVrivo70gRjWkMbhS7p3jEX/PfWHxU/r
ZZ21gcF6jJTWH/5vbNLBdjT2VF8HhNMn+Oe0LYx6TJUlgmvobuQmo84O58ri2LcL
`protect END_PROTECTED
