`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UISF9M/9adgWHHucqUGGqHQ36Tr2vjmWLQu+PxbdB1Ol4W2m7YdJlkYNEYPrOgxm
oT8c3+WmOsLLP7n+8DGxDE+q4Cf3n8aiZXQtJpx3rzgZnZ8+mz1I9y/d5b4Zw6gF
cCuZuBkYSEEr7fWvVfvyUTeuEDVaB+xUeu3urGljE7VNFUmkbJ0MAVbwKAVMCcdJ
rAPYFTcJjxrsvf0h5pF79huy5+opdFDcS65y7wZYO4jQ3g2dxTg1PFw+nbTjGsNh
uF2qrQB8JrkeIZPJi9WcOY365jgyx71lgPGAG6fTQdT95HnZqzHOZXS3qOiblBew
Qj+Q7ahm/VsFuHuAs/mkVt/qIRjzU5/mVXjR5MfrqyhlZ+hUgEiyj9U+8B895nK+
at1aglbpCjg+pgE6VjHYIYGajZutt6ysGvJ8+RDUzSg=
`protect END_PROTECTED
