`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kaSuGObbYfLD7zyo82r6/mbJ+UC38xqgiM/xBj10Y24ZweLXRKC7c6kCks72LBlA
YSnkT6hYWOHv3gtmx74h1mYhPVrhKoACkAY5YBOvni7U0uX8pJXv33EjdVgJCZLU
4Fmn+QNiyXbRODFHPqlQ82GTJpBV6KEj300ILVi+l9h6UICCHjl5TxpyGwY/2FHW
qvaGdqrxPxi2G3aDrSzEycizb7tIRY3wP7Tc/UqEYSgnZs1Y0Ob58s8CwK6H/fBQ
aclg4IpkOb6IHltxluWg6gWyWosJo+8nTqsIUZQDs/eGvuUOQxtOqXW7HsjHvPEe
ZcLlAnp2G1cj9n6x+nXRCBc/zGUrP1JxpEHMWqX/Ak+pxfthEPpG4Bo16eTdTGmq
ZSOPKXs76jD9DSVd29/oYfaDD6Afx4c0efwIgN/EJsxh0SPcVgI4uHbl9hnP9x/C
9PqdtB0t4yoPmH3T90Iyj3c1QphgXiokLlqeLoVe/m6P5NHYHaKiV1Is/bjU6mzm
wvgMPu1TW8tyAk913roAVn5Z/ExL/j23fOYV9HLTJZwTahJSODL+1jdYUDFTKyar
D4mxbmIfDJMPhzYUL6H/qBRMneTMburRlmxHJfP3zZ6l+gxaMdQzB5gCus/56Yob
pBET+RTx1QEo9WmxxSeLvA==
`protect END_PROTECTED
