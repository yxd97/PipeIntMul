`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9+RorbpqAxQCSpVxX3JgHT/j7eU4oLzlT6cnwCd2dQtU2Y/LvMHh7FThXzh2puEJ
AezeG8tLZ/tK9kLfNVYxUjwXVi8r4LMsTwj7T42FklsrH/TSkRHjyvPbqIPuo2iL
G0bOKtUlCbyoxd07Or122eihdJxYe5dT6g/YhJrap2qq6SUohWQi2hW9gVc/KIsZ
wyNSh912qCrLX2fQTueh24+cBt2rEJ45q01vHcKbJf69WweMZChHKgmZiY5UxOV1
6l7CSA4t6g5FB4HlQneFRourpYQ4Si7ivURphKqvecLP9W8YdT6udbtwDI6n24WW
Vjm2QcndjrzJDdXWB9YgYRphLvNpOK58UHAWbbqnxnSJZaZaPIX+zsjRFBjPKvCp
80YMc3GWDILkujRG8MI7AmDI7Qt6hu/yCVsa+70WbuHrhhmWbs1d4FCgvKdPbB1K
aDfRZmnKRQHNbQ2n+MEgLyK+XMlsZlUTrZdsSEpJod6fM6wigw6bLviVV741JW4B
N51LbhuQpKgZhoU7DlUPQvKMpUj4qvsD6IWIc+5vAQtMvzjVVejnYhXTkWEciz+H
EXPr1+/S4aqITkK1hb6KDw71aXFSrS1HpiKzEUHPsm4mzwk2ZGw+QvhKHrZXL+yx
VJLgFCcUbQ+xe6hOP5wvwuSMSxw5T+WMTfMJNQHdjVSFZlLtZ1pb2hjzM8cL1s4m
3F9Frg8KIDZYC0qGBrI9xuABANFeDtYl2qM/0/ReeYrXrP+ffCycLweCSNtXjm/m
a+QkzWy2BxzI7vnWDTu60itbMimw+x2t7Vq+PNes3TsJmuzMWA7dUIAIUzb0gNdj
tn7Mso4vqSK1WlPNakGd5tJrOcnmsA+QuKj4MzbPf4fI59VoIIWLIKM0Esyn9YZa
5aH1R5ul1L0M4tlYo0JvKotIofv8BG88a9JwBc+d3oops7hNRFILAc72oFtQt5Da
mNOxjfTGslP07Iee1Pue7BGQH9ZTOjVaAxTDDULu917hTKliipKHECxhd9a8oQpZ
5TcspUtRiKuVKLE+AAQai0YbGlfMRuhnlEC4Cq17eGrdZ8dxP7Qwf4djSLA4PIm/
S9FmXjCJwOPbds4K3TofMrBw+q85kXDlZzmRQ8wWEqr8vxqK4/caBYBD6IuAGpqL
qfR7IbSsNp0/Rd7aLxNnmCjY9VHWEZz3a1j6VoCVHNp0ddnPkBfZRYs1wEfL6uGd
727IBfRc5HriMsulgT4nDXR4KxJ134RFDO63dJWc2cbWCalQWg+8dtVm1cGaCmUM
zhPX4syKen66FxPvw66GQk/dWZ7vUneSE7CpHMi9kg2LFv7FFEfA4zAKiv+NFPPE
j7cnk2AabuNBRO6bHyjG2Dc5qqQgyTun08RjEbH1ZFkvnMqbDppmfq8QAYdR2wFy
zUmmQwqr+6pvTdG7FR7UmJGn9okMXNXDwpDP8HcmHsknWv+Sc/rwync4y+KJsG/G
Rus/9afEP7Sd3l2FsG5cMg==
`protect END_PROTECTED
