`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7pBg3S569eLPO1sU7oeTAWpesoC4rCRN52hYGF6F6AXHoG/pgNMVbCvzoMZsjpa
xvUzNg26SDCOxYNSnOxRmihz9/qnbXJzklbNCJwPt8krfqOf2n6NhcTnWJPocYva
EvSznfR1lZEmAU8izkYbFsBFYud8Z9iGgEZ3ceLKpmoTeackdqnMqc1Rgawr2ZNI
doo7lxgUGKkbBfO/slsqrwpnENuqX25BgRsoiNLWEQmndxAEl9Fm2AQKhMuamtRM
MJtyABW+g99anrf39KCT2I9d2HKKlQ2O38vjeK6YGWZ7xH0SysHSEcqVu5En7fBz
eh/u7f+34ZZB80k3aRddFUm3hblVQCqBzvABWUt7w06ljVB6evzb9tNGmfiC5r6L
qOQ12vA6P+KQOWLcvJKNkEjmJpcGgZJY6T+bnmnUSIEk7cV8B6vTyPSd7Pp6WpPo
cQhyr2bXR+I8HaOF7n1wLoxVO2V8ZpVuFVfJ3rJ7fjUWHo240UHdLTS9lMp8MbNy
`protect END_PROTECTED
