`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLIC0KlfpoykAAQuhbrCBckoAYhJ21KmJdpnKrbwBS6aCwFNqeAfyZJAtXY6ldkN
T7MRiZtHa+MdctB3n0nrjW86wkXPCw07a5omaSst+cqo5N+tliEl77gxclkaLj+O
FHXKJrtKY3pGcSryfpbcly78SmZiNOP8JiEqIfOeFLob5wDadWJrMgPrH7FoXA+h
B8Xkkfi1bJvPQOkCW1G+7zV2IbUor2w5kvJb6SCmvTH0ZzhxH2/uKFC4xH0DVSAW
A6iyvXOIpe+S40DqxOgkoMt4Nm4F3zb17S2wbG4GtQLOgDJFBFoXaYyvJ244ggcW
J2J7rGYUPOJVOPOCT5C/uf9lr0f5RPO62BT8ll+1JacjAO8e/wPpaftiwGuKkHHm
4+1ihbmFJ4dQLK181+GP2bqpfMRTMWwYwHuwoRMKLuHQ9CX+K5F48WyW26Zwv/Hd
Dourr87xLBlogCCgScJg6Mu44wU/HPYeggNtQX5oPsfuUipYjop//6l+1K3CH/2f
m2ssvlQ9WVBsUJsCtkFacdjd9fE92KZP//1/kI/g8zzAIGwJJO+mZk6UeIQLPncp
x422ztOyfFwX+GPCGEdhFvFS8Z9zqPhJ3QhC+oL33C3wgUc5+4RX8yXbMOSrCVQj
KNYUzyh52VsU8KamHM8L8JDqG4vt8ANCTnL7mgkORqbxDuXq/brKNBWISQ58yLKG
MmdL7TYzCyhsbzDtlUW/LWpEjYUOzsk3z4J7WbHoX3FH2L9KzYtIMHv3jwzRAOkR
lMUTG8POHEGjEHjTjKnB4id45Ig98l6fmDR4WuQ6ZK61KQdV8dR1DR7o96FLt8hx
o5O6NJrh11VbTVI+JAPNYwR8PhHZC71IOEW3igiSuyjK63ivpgyqBQCcGsErUqTL
TNmhUwJtk9rx6TcDMcgucigl626E59tltg1PLtqlzrA+TAyT68sOxnMiciDFRX01
s5o8gYTScFvvmrRuUMiV/4I3X8vcx9Ga4g/6cQ1/Xp+x3YjnVI5bxLSW7rgdLGWE
VVkPzAw+7qKdA2Fp5jQxspLBQ6uRs7HSE3MwZKJ0Abr4jm+pc7wpq/KaH5+35zib
P/NJfIFZlGuEgc3JZZZbQ0e9Oj3Z64kYbjCrEg2NU6lkNh8fWA35E4bX8sIjs+6w
tftcWjJMDU0IiRwhrtN9CqTAAxTG0OBbDp3GQcWkEBWZltvK3zjgGrfD6y5OEsjB
u4o2S32eAwRdf7k1/azdKsG6rADKslGYLK/U9LNhQ18UB+q8HpnBRSxyyOopjF5K
Yd9KLaa9h8l/oL7XULC7PdOAUrQyzwccA6mnpmyQ98xlWLlWKqiXwLLtI4aSDWWf
KAgcTFNJUhDk6BV9IdICuEKTHqnPkRUXZgb8lgsjxr4IXUds/V10N41T+n5rQU5w
n6BsRhXhfgBUAl5mBIVSpMR7eciTQ6UMKACq/H3YlNw=
`protect END_PROTECTED
