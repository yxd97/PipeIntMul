`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XoAO3cddxdVUuIZXaxczq0NHGmeMhWr4QB9NUX+i1BXj9m2DtAy0y2UDARUOzJX2
HZp9MyHtxDIe3sggjy2CsR4OlH6XEpVyTd1gS7yPHR69N65chbiBRZcw2M1aAciJ
v4iKumsd+yMd8WC6rfWn/YeeRb+AVJiwGb6IUa1pHVgB4V3xvgIRFdXjL+dL2yWa
H25+4uYD7cqR1OLOdxqLReqOC8rdENBk1Vsv8YAHpX7IIG6KcLVL/9BzfL61lqHv
qUnHE0GxdjWwvYYn7klGmLlKXaGU1immww68cHf5MQeSOynvDGsT29KZI4o9VWY2
CF7Gdl6Vc+jcDVyoHHGYv8zzG3FaKO+ogBKbqFd4uCTwndc3G7sMHhmcQyGmv/pH
y9+5u+MmzbtPaOfZW9v5xtccTdhGHAHLV90H1YaAx7HtbT9EO3PE7+jWuyh89AoL
/8boFhq+4gqQryShAlPL5jS64qQUySk7hPjv3fIw1S00HBp2PrCI2i0Yn32xmIW2
dfSDNFQ9x7ebOZQ0IP4WrPPqR0GV5eNbg4SHsCnomn9YAsErE0y0R6c+hWsc9mJQ
0bj2+A694af+JUhJ/HY0642c+lxDcBfoypD3HQn0XtLVkMy1EHE0BafTmBAHmomh
YCUDtYSkIJ8y4eXePgAgWbO9MBS0bz9QySTZQEgnwmyu+b+ncL2R1/1XquymNX84
ySrt5wv8Hy67xPSSM60dgQVCohduPlRptrKH9tKnOcp3zoVN1Jblbz4mYtCaEUrO
4lqaF63jecEP0qKPXaIk/jo/9YZ57u0CwzwMNwtO0FVjH9cHDjFGrFUfYQxR7y1U
nequ/W57WEygljgBsm5YSN2NNBxjKo1ATrLUrDFZ/H3W2V3DBIICGz2HTcmj7oBS
Z/EahiVdoFq4dCzTU7zCRxQBJTjdTK6Olzl3fq0E2mFbZX6Gp7EDx1mcPNo/4sXR
nCJ276AzNukmr0G1hO4fyYRblWpbcaOFg9PMPZ3a8QNHS+70+hH0s9IJqRxNP98t
9G2r4k+a6xO6hOv5Ij2laBNbGspGQ9kA+AFqvNAunl2+2X6UAHSXG6CMnE4eSYhz
VzNa9cEifh7wmTxfsDjZeB0zJIuXiuwsEsbw/mpmqyzXEqCW700pK/q5HXuA+cCD
m9CwkACH5y5ofLaUVuY8AWbwUmAWRte3j85xPk0pzDiLflF40/BsB1If/smzz2WG
1PoJ9BViUyhrqTemxJk5aQJ+u8LuFjVHOMcWDxT6qqEa+/dFVeASQop35T9uBCgi
ZZJZ6krLrwZZAVG6CQ2dIqoF6zn2uSTL1YWVTtNTswUZUjoJIZ2efmtTNL58X06v
ai3mwKIkSpC27pwlCd2nNZ0iYHbCBVKnVqMvRly3ti+wl/SsK9WHqi3BPn3/OBAF
V+1s1gG8AQbwf7bGKuL9O7t/9a+wglE8r6BDRSvp0IIvNk3h18BOC2ZPr+dtWH/J
ecGz890CFSRt/4R0updYJv1s1yf/HojpOmZcZDSkFu4rHNUgwc1QpCvZlaymBAby
sz0+7ZTL+mXaFwq61I4EXuNsyyox3ooLlh1ACQVXvi98uLBWhiGfKvKIF+NmPltS
/gSOSlYHnx8SbgzUXf9q6IGrTVLiJpLfbhzcmTiPyefvKsCA3tOKybd0Kjz4AJLZ
aJ9VZsM1RLwfbvwprd44NkKDzDFTKfxga0K1k3N3CRjvXQwt8jH3jwnvOQn1Bbyz
OXqxDf4ermumOujcLADVjsMeLMcmoGKdy4C4ya7lM3D/WhuOW8NPGv5nhmGX1Erh
ul1zTDC9VdGZf3tLZp0UwQ==
`protect END_PROTECTED
