`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hwMgBuT4F45RPq9QMZnlRdkG30YDVCykpL/IkdnDjGkaGT6dH3c8o7wuP6kRy9U4
d0HqafxZ1VVSHI2gGSAivtY6E8uN1xF+JJOm4dwC3TgpzJVQHBOjfkL4YPPnU6kz
Ixi4C5yG8KVGrfTbaCRvWfGKtQo5xGffzKVfm2O/ruiCAdEk4sigh0+COd1fQBZO
tZrosUKixZTTA3unnIrx4mRZ6bAmHpR2+n7HY723+epFDuTYKla8IinoPTdGOO2l
AiDm7QGMmoCB99vgo0OnhhT8t1HqwGDfCLU87w+TT/VXL0ZccL77iS2F3mJxgLCV
ix3+S13rc4E3ZNBHtp2AOg==
`protect END_PROTECTED
