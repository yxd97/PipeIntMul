`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gyv4gkdiwXcda6pzpqYrIv+hlOZOSEFIBOEJiWzzjSARwllgCv5UYQ7Z4OqKo/As
jOVLspY0TKk0jdWNjCbd65gJ+9TBwGoEP2UEguziAY70q+FwmRlQPhmIAJLiwYwd
pOveuKIQiDLFZO4WkNXKKBKr8RJ5xcZEirHK/u/GZ4pvLDNw1Er8sPRyT5U3xc9w
2kKKoLUgCu+FT6gjc7VP9AGRIG9sEwDg1GpwQS5WjcPzTcn5+CXjuVX473s+BTDX
hJC0NRPADwUIJVLVgBDulEvIrVJYbRekE687ZdHehWd2GppZncf8eDJX2BIjofWB
8c7Swj5DEFuHiIEWEbFfhkEKNXcIkn/UIswPNpXjHnOa6JAbibII9lNM6L6pS2UN
8nyoDfrc+uxZVXcYzHd0K5dCQc5gW1c4icMcEjs/xtAiUtY8nDRn8K+eP9UegaZI
2SDBrfJi5UcZXM682Z6aswWeKEphwjS9hNmAh6Mj8sQF8SzLBTh9aOVE/zA25LdH
AU7/mUVj/0YFt7E8kiqWFQpf4GxfpeoYxkTq6EIvXW8b7KUm0OlVO6y6iwW00RzR
K8QFvrzic3zgHsDrJsHATaVoDi7JSVSdlAsNInMK9GFy6bC0uwg+7ZQL0HrIGPM+
L5VBu4KDvUdRAyD6SHsx8qz1Yl/HkjNTwOJWYfeADnZC5TmmiiMUDWudhEFCvDtw
fMx8lGhZoY4Ziwtqsc3e+ehaIPP+1EoJMEjggGA9SVBg7bQ+ZHkp1J/qKh90s5Gy
dE4Y/juwteghoTiyLcFggwmCkUZyvZ9ga0LMd0LFkzSXoKjXgSZxAdda/vO4QGu+
CX2LbrZj4T/v4RBaKSRAONHyy3hyuCXIfSP3YClhht/ar67+zRcpxVg5V4qND9dJ
rTE1tc0I4W2glze9fQwnAMwzZzeaipTenfkBhGPVgO5iAPOB3J/QmxMGGg80V0tM
kIpBpOJtNMDuQPOQolZfywV5VG5ZWMmPjFp3jZrFP23AeziFOcKUcxemRnvysixZ
NHzEQ7MB0mbb6Ni1IiMSe8N8GKObOP3+M6vyhT8Ebl8Y+L2+KUW0mLqcfTCLTf4p
fpzXX+pRQSxcZHzcr41XxraGG+F0TAr+WBmIQkjdb9iXQz3X0KrxHXFu65Mjqo7i
mhREq1AvB6taZYCsBemeJIbpFnqw7WRgIB7AiEOYcEt+xCW4WtE3eRCnwSodasP7
Ow/LkjO/ONr7BXx0Vo3nsmCjKCDZ7MWtIdM9DQy3r7VxKwEvrBtduSj4dSTm/1MX
i6hGGG/a4h5MRbJoZMBk0xNbbTCjkHXLcQhN3Il53z5QLssn/3qbbPpKx8bJvmpb
2zj3P45cSIAGs2ZdfovmfZV/CBCPWPh+MgF8mi7/p3l3EYSYaunTL0v6SB1OrgXz
EWwDAB4jGFAKkTElrHQosxadeI084hqRUl7t2ssJEzjxQYY/6Rsz3zAVblRuSPT7
I/as47Z5wN3eQzJG1nVIhvQheN8OQP2QcZAR0Fip9thdPaNZduERxn1GOH2FjzLA
yHrGBXgZDwkb8veV4Jq72k+H6idi2elHJVyfywROknxprGgqKOXQH1KvfLyUpx5/
LCu7z3q3nkZEABTgW0uC4rEAZoqUzyAyIeVQWo0nG3xxbhNHa29NKyMSERcUdm3P
/uMWO0W0gFdnw3VQHotNpqSHAyXWxLtwhVGRaLJm4TFH5vaADiCtJEIaaRMRgSA0
Z2bNnLMTsTQUb9VPWJn2ou6Hux44legOhq8fxqWWFbeekgWxgK11E61nNUBhbam7
ioYVn6oWUuxNw5dm+1iW9VOnjfb6LJ2Qk5ZKS4GY7fRkhwiUxj2zM30YJkdr5Yju
DD/vJHWUz1FvgNLz273WH/TJtTeW+b0TfIHlMkgTawyCRj3LTkp2n/6t7kUmH2Y0
vvL194aWSbsBfS2NZuXve0Icqu7cQrsHbeQD2q9JHaZbKqe2N73pS8Z647PhnON7
JCPFZSjRDlgr0rDN5ZUNnfwEY5m4w0V6OQf8PkakCWFSAXvPiufD5pQ1nZ0oZLFq
Cz3ujXfA/shsjpmiK5s+MqFBgwCcWxacB9RxAR89n7wpVICL7ID0yo/hXOElsfpU
LFroUF8Pu3pM0MnW0W1tZSUW8rin5awntk+QboPCc/XspSpKBw5Se6fNCFxY1jBs
bJa9O5PzSLZXI3fnfozXuW3mfdzhMQXTo3MsaanEFUzFFMd2t/Z5aF+FAZd6P6ea
C+S1LVQNcbHjJytckD0LI/vFJ2kuNOE6JVdN36WoOwLK1kMPzKZHrv6oYrvoawy2
0l2Pdu8XGRXzbiJpd+tSi+LdELe5ResyPIUU//lnaS36mALQbksnxavpNMZH/Eew
UkDadDZsN9Hqcmy57o6gAw==
`protect END_PROTECTED
