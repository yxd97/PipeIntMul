`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z6o4cGClhsFJoP9QyojbiZqW134AW/mQ4Zff0RiCvbrl4v+abjtp9GkDulq3xzq0
zaBwVFeLIzFBmxdWeCJSk8Pf5rpE5sbkRFkzDat7SZGCZuOauUpTMNuB0Dg9taSu
Fl6mHbjZCW+imH565TMdjGynVTxYxbJigl6bWfXM8AWsbKq6yFnZ/Lqy7TR0GFbB
BX+Fsuc01I6VGLuA2tF15gvcVwENXvJbQCaRGCk6LIWhxgkBFdH0cLyg07m9qi2A
H5uNa1xgUGKX3zvS98kRN1VKCLjUagvQe5EvzwPHGK+AoWpDDkgPKK6cKJk4p/3+
NBVwnB+xMOSi6Ikze5otpyY8uoU+GawjsCSwYaghvDCWJmzr9NXFN5UrvAl+N65L
f799zkAA21g1qgajbkvz/5Rh9swhgP4m2clVhuFlE9E=
`protect END_PROTECTED
