`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2hriqnSWx0CXUTQI0bVgX5/2AE/4zXfV7YMd0saxqLYzgMjlEqbw1+UA4dz0FDXO
0FYXfYcZeIY+5nLCycBO3fbLRGpieLg8y76JT24kDC0WW652JtpjdMWCnp8+3IBK
2m3lW5NIsM/GxvbBl13B8cLjJ+5QeoDcAvHbevRbxDxcBGpNiWqigo3FyCRLBe9t
FIn1aHpoiVVDsr5ENQHFMFXruHzOKmZeG7ebEQcO6dI=
`protect END_PROTECTED
