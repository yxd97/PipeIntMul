`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XX8qWsIEAAGDSv5oMvDJ+9Ah6sgsxeDA3YFwixtJi3lAdonmifMi48U5vI6TpPsp
JmvznEAWti0AypIDsBF2bR2a0sDMpfERImZplIF2YOWRVUKDKw8KhWUZluczzIjd
cyw6wb60khr3nQP8M/3ZNHylCS/MDNfeduD4Qfy10PtKhYxpctcJMA9o3XDlB1FE
ffrfhgyUcYGEia0Hdb9RwmVFw7WcPeE62ZukPHz8D6umpA5UOHmSboGu+oYS22GP
nFqqg9kL2w7rCbhbxJtgmvkya4UsfZU/6ysOVHMSsMnGCAzXWxEUsqY98gqZFBsH
cuDrl4gkJViLcfJrfoYtyyJeOyojLJ9RiRGsEKvQ/xnVSpQ37Ird5Z4ZC1NGtpJ6
ctbCIpJSpPjkv33JPkz5AxInRyi1lGxXjPfotBAzBpV1S/MwzMqwxuw+WRVBjtNi
WxeuV8hk2gFM07Dvk0ANCXnKBnM3IIM5hnJ+w4fa3Q2v/YW0Q2s4YPWB1mZWdsKD
lMiDUvbXHOPSncNvTda/YdsvYwAxZlEH/cqircJzqNgoC6X72PVJBWiIFdieOJMg
5fA1NE8Nb4gOBkCDOXDI2frrftsO7IrmdirAZEt64z/q3HqD42kJLyGno9Pe9OJ3
Uv3lmwARvDVyQMLZh3imAN22U5Jy2GSgnZkCDZ3aQnw4yQWD+8zaY4GhFM2+1M4q
5Z/33OuzzX0XTyCqIFSt5RJNRc1gmN2TALwq7Ca8yTQue4nGizI0bSU5IJiFI9a6
9URpK3sP9Ege+8QB9t3Z/ILThcos4FfOh+WluhL+Q1mI6wiAyqxKe2LKoRYUaiyY
5KM75iqLJV9UyPjJoXK1JVwVpgkyfJ58je8iWHn5/f0PusO/IMdyxVyo1TEA+JFq
zZKvuGncbby9lTX/SR+Oju+XjPkiBxadPbOiLY4wgjJogauWgycYgBQx2qYH2yjn
ra6z+jVz1kgvXuKwKKu0Vwqxj19v3/hRUVjqokJENGkHGylpIb7GFcMoePFlWDmq
mkhTTkUKrk7SX5AaKz6t7OQLVHqfSpzwwDr7nuFe2+7ScPgiohYa6JbOLJZrYlLK
VAGWdCqbYsee47Od+s68S24S/GcIZ3dUYdomRSnjtwWQviSf3nqt1GrvDzc09KBw
`protect END_PROTECTED
