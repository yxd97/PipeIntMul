`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SyAcH21AW6AHiTuQA08GIXqSF3/Iewgf2gafocZtKIqzKGBzPTdNc8xlZpF771iI
Fb+tBN8PAYt2u2tiXayrY2ZLfi+91ATetxTFrbFJvJzhNLu11P5Mdva9l62K/Pod
N5ctwJ2TY2XsJ2rw/9PGovSDfkU6a/Pj895UikXHgwfxgboKnbQswJvRz/Sp6jSy
ylODZP6bXtJywZ5lJ9rL40dR43oALrm9fPf3KCabEOmOGynCSQEKhS+5CfbPO66r
hK2YaCsKL55Jm2b86sCK5rm7Sot+9pVrq4mbqPF+oQMgz8FQZertqdOM83yP4xrp
JTc/WeSwbYTQvaDzdOS2//JTuQY55Te/P6JDGDD2KNOEcS0RzdrBa49G1rlvAYVX
U+dff/VWZA4xn8SOeUqgx6KAY4hvPUyj5d/s7Mw1Gx5maKAyjZmcYscwWrdrTAs/
LZw7I2EUcdkMTEM6VgvQgmYv/DwWLA/iCfKbjR491ARyikBfLkXPEHfv02Cpr0fI
8BuGM21mU0QckR9ls+oHGkUaWlQI8eF3A/m7a/Tv3IjtZCJ4Lq0Gs3PzDNJ9hcNI
ly/fQHWa7qgTPBfRUogaZQbl6BYESVKXDOJqKSx70/V4A2+P77BDNZPMQTbP8E08
bd20DTTEONM8HdNPE2hLg/A7BZxniBSaXiEtHFH6sHV3S+OSf5TcqPKfmEN+zswz
MtqTIVimv8WogIcA2AmPoVB8JcgOVluAw/p+sY0yCXsdLWzlSUXNT6a7fYCYYDZr
2xp51vC0yTivxWSKygWqJKLPE8qGTzYfM6WW2neM+XZbX8QsySROfCOq8m1xP6MF
LZ8OfE6Y6Iro+YVeDViH72x8gQHg0OAw/2iuW3kML+TdmEEXL83iCMAVBShc5gee
STdzATdhsZQiohEGLDIlcpsAx7a9vtjRoYOXqRjbDDBnGWf26xqJRl+VEiIMwtei
k1rkTvWhMcMSjlq+fm8aj17wGNasyxjsqIHfdZk7fQvY3UwH0oi9WuASqGYqBp9O
UNMIGRLNN4rfB0QGSEZHNwarCuzk+oYNp0LUyjuYUomfQ7+3WHvxue1pmRS8t1W/
+yUHIp5/v8gXcBpvXbURZQ71SU/JniBXZWAdDg6R9YEumm2zR9MW7F52M2HOO3Yn
cBCzjXwNHnAg2NGAlcQSGpagujxc2V5LJboOTzVzdoE4fhyFIjTmQIvHk4e7U9iP
j9FoTuXCuQdS9WLQiafx7osU8anNREYKa7mx9bISORlxCGjLx2yUX/B0D/OWyBdr
`protect END_PROTECTED
