`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZwwhPkV0RCXj6Lw5gKX0t+vCKV6ITkBZVxI3nxsnAX4ZJeC5a2zZ8SeioVn/fX+R
NJv8t+lb2s0BNPHNzNMkUWgeJURRX/YFGcTUEyEWECGnWBSR0Q8T87wb6r8bYbEc
ldED/hDf4SWUFS/7Ex23zNv4ZvVx8fTfv59jqaMUewJ7KiVgrQGax50gmPeUrLj5
Y37WGGLQA0ljrJBKw+54wIx5YiKeNXjAvTkXpugNd242CYT9P25lEwqAy/5ECWXP
6APbwclqtoOmmzeR7+nJKyemUh+4cfzon/N9hK1Xvw9kFhxIgKbFdG7Xy8lsnhBs
xPBC7pnPkaSZazWzK4EfyXLYvdnDIoPM0vJcOxbXzOyswV8ahqMu5CqcfRCyPvqi
0hnKvNf/ASH5Yq4bScvdSZSmIQEAw4A4fzng5WA6icUqhRLZ5qPzvM5q2jd4vFls
Qm56FGpbVnwyZBWUQFCRrA32lFc2jJFuic/gSY71ICVHIEUjweRs1wBhsmviY3in
dnP4sGz+aZkoJB7RcmB72/XrpTn+Gn6MZOPCrH1Y1LA=
`protect END_PROTECTED
