`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ft2bYXfg3udVyYIRSXg+sluuRv2r3Z/HWvu4El9NHGLF/TzT2NAJEh60pcdNQOly
m8n6t9lu+use2V0N+cLkR35htr49RP6BQFvaZh/qdhBFW1H1Oy7h6XVl++Yo/wCS
cTPfboC9kIcw5GOMzLQRWMfq/5xUOwGORUlLK7W8QkrcaAffg9WSp4Dhr95W2k+R
YKcRLLKAnre4QXrX+QocNARoBfX9x7JGmoRpgvlrInkN0x2CXRvclhZYrIWkJ4KS
eacl+OyBbbs4e34APmlOdrqmRQbBPnFRNnlcgQVG2dYuPzfPX1IOu4N3z6C58Mv+
x2UD2mpJfp+ISEFr0M0CWDG5hc16EVpcvHsqZAn54/MFw7J9fpaoXkSgCM+QC6zn
mY9h2vHLDIcdBvHepKBH54SnkH1GjXsQNaGId2ibzQg=
`protect END_PROTECTED
