`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ss6O5Ok8YdOJEX6cri4O2Wre7AGeN5/H4U6VjUeScOkBr7xuEIF3dwmabV3s7x7i
BcafT9h4mQDMZQncZNzlYw/vmfioDsxK/1vITvqAYxnbIX4hIpp2Tr8yrpJs4doK
lR8yvCi+DxrQI+gV5I0oC2igvXlPxVwSWoA3hsUjb7l2/k6MViS4N2fdjfFJ29/I
02khGop7RnenXhxBYrSO0TAquXRNfR4G6vusadMG4X0qzcQC2n2rH7cOAjpiOfPy
v7x45ZzKPoS1nBp4VDrL7hQDcQY3Yxxj2HA0zbZocrcg6IxuOQAMcaePX6b5HviN
LmRotoWNMAOpvOmYuZSctLXs9Hf6Sn3fy9VqojsxTMgL/1QGW++7U+hOexteSSeV
6Rhb2YdvO+lz5JCdwlnqgw5JiWzgTjtqtieNE56m1AjRjXKGLKGIvQioVQDfiobp
tg1mWk2ansv6c/TOxCAHFANl1z3RG9wmC0CHzia9q4KLt90Y5dKrO8rxRBg0bBCx
ZL/poU9DrBGnGDt4/uNW2ZiVkBIx0x11UzfbefWA43MeSoWotXrUduoREhpOtsxd
arbt0zSoKGWPnmSMRniHyo6u2LvgWYbeiUMBMn1w0hKroFnXm2onpVnaFZi0/g5p
lcniz4k8zkm3em2mHpOItGpPUhltB3F7Uif3WNsZyXXR74fFy5PaKKQ9stj6JGyU
t+w5iKHt/Dna0nNGyXcsWGj3jBk7skuNL1YoKthLD0UhE/HJ67cfvoS3MwqTtfFD
RPglV/opeJdSJ1uxK/vTFZWRKODcPBlDIqiKwlRR2rdGphFQgEniM5ZdyFS52pUq
0IIiwYEDX1qQD/7rczUB7QGNP7lUboaoxuDgAB9aF+ryssqg3B0qLZ1+r2ThD5FN
b5lmDUbF+ND67u/h3b+p7jGx6q9KLprbjJ3sYuzDPSZIkbuor9bf2tG3oZ8vG5w4
`protect END_PROTECTED
