`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0PKvLUiiQDQN9N9bb06ETonSFpIELw0jvwmwDbmc4ee2lne+3CxaHt1dAGnRekA6
RTrEsBxO1+PfPwJSWaChQqbuTnJzNkxhvAX2QDIpTVkRXq47ex1qXOyeQ85yMDU1
0yK/Qv/2UFBcVu/yJfEWuweFdTE0a0pypKp29/f7vRLRQASG9jY/NaNAj2vroG7V
e9LrxbgNZghbs0bo5I4I1Ou/KJdAnHw48mUqHqnF71SygGtBw72F9S3KqtkXwmJC
G/1YBoyvlksi6EszEb4gHMiiUDB1dHyT/xM9K79s+LhxIsZNyaal/BUBmP4mtWPS
REiBj5OXVZ+6OPughExtcb48pXe7N9gloSAeWo8blTIPSEcQv61KPx+Qo8eg9eih
/r1tXGqzXClt/aCgfQzQ5fNb0MHC8YwGKhTo26M+afMIiwsZlxOhCzOutPqZqnR/
C+uuTzQVGhd39tfKnZVU/ANLzeVDliI5GAe2EPFzKmc4cDqiDN5BaAYImqWAIhCj
CmAA+lDmmSm3mu4UWh+njUJTxXiTjSB+HOp3e+9NyYqGtRwy+PYgMKW5zwh4iy1N
M/fZp/T5dh6eIpA9ca8mbtCfYR/Af/Z8gwe733R18FQQc4qqT6ZA7cvXpHtfn9a0
JkXd8vYs+oU6ddcLIQHDyFWjVpyT6TW4kkY7Cx9UfYQBLFXSL1bcml6EuYGP9LDH
vvL5dUOa4HlUmDB+rY3SFQFTLkL1ScLhB5diE2+FC1LqOg1RFEQ1PXEkUWczavEW
GuKe9B4qDGvgvvDh5oZQ+VHZ35VKHlrZ4MLv2+1moXBFG2GiizpNaN/XjVvUyKn6
rjvqRwVcKizcG6Agnuu0eFmY5iEu+BIkjihVCPoqaymeszVpn+wYrqtXLPy+VtGK
AlRMS8bYUGQkxyLTDZaezyI1qzIGDKI/W6Cj15hjKHMg00TbstDtxsBeUlMR2L6x
TANLVLNQr7pfew1OEWcM2eyAP7VVlw5SmOmfU5hfWFl7IvkaRn+Jcur4vfVQDHMq
eSlb0dQQHT57lYES0dBRDSwZbQoCyIx1fgX3IyVoLDhzz9gRRM3CSx0dVfzObo+J
WTkwe9pm8S6ihkqSKTLUf/4KdFRsMxOM094+ang2wiM0ci+65igQ6R7VksfPNvLU
3eIT6DQV5k7okA6PKcjrE5StmxIYzhIkGBkmb5yj2y71UPSnA/mFjSDZpfahLUQ6
rNoquMpJv1Ht2Q5tVNf7n2LIEVP/AeZq75TrxtZyj7db+4Hiyw95WljWnaTNGYiR
ARYhM8eXcAFr3ITz8SXFWsEzzZMlpm7PRpXq3t0i+Bd6YQ2WZgh92N0ycQB/KdM4
WZACC1peeNSbYn5zpwbB0OBWMB184WfzGx4DI9I7DMExuYe+i6gvSX8lEItImQel
mI/ToUG/k4oZ3R5Upj7UjMJRGEm/rQlUiNKPQLOa6lCY0/Hbu6g+8E9MI09LcCfJ
WaMaaMTSGRnzAh/iXIvp3v9KXqxLJdz7xzdwgYU/fR+aum+605fSQ8TEPRNh0OId
vNoGYyIjOc41IoTDE36gsFxLuqEr5fJBgS7+QB6K9BsYD/ldhHtLjSOicDWCGxue
7oJK2+iFi8P6SJ0cZgNbmfrC9evxulOMdtMsxxK80px06U1ghKhedzg0zcIl6zUC
yp7/RKqTKCcpgPG3vP17PgfD5zcu6xPI+m77gtkJ1pSSQPF+yudL/o/269O7LVMx
4+ubY67XdJTUBpjZuRAQQJuXxeiQJDAhyJAw0XOtqr8K1dxxoCjHP5+K5HL1cWYO
mpUyzwhqSWGAZwWjm4gbrhhQry64zCMrl2FRb6yFQTyp0ZqNuq9Z9SCgETyrCxt0
0SpBYqdctK6i0+mzErg3EcMKYDEdX737eiZSjA600RJFfcQ2pWoXHeaI2TcSL1ha
IrdAcffk2OYpPxQmmw9GkESOQw2rNlV4QOtAZ8HSZdJJ2L0bQX1wU+bOEUtDCAko
2ZBbV5RKeeDQ1dVH/nerZtlWYUwiVT1WHxy9oQoCey2P14z25nCjZ96hYhpzzr+O
+O5Lx/oh1grzhDuhMweuMVOuf9MughDE5gJgeXFLVOy6WGCKevKDGrJRtOvJkcSq
89QMW/q7LRvPjAtAF/r1O895+yS3yXlYVgWE2+zbjLQmJ3fifjckotIsPFBD6rsG
nq2ph69eZpkbFcQVq9PpGBcWbSJnL/itd3LHBfwE7bgxBho95C2nhKQgnGLp6iWU
qMm/Ed8h9x4Rq//r0ar6XCm/MMUkWvD/xc9H5jTjhlN2sQbV7zSR0PoHrwcVfUhp
hsgQQPKjyfQfxrG10VsiFIuLZmEBMD/uH1354iQm7dIdKs0jwuF9/LzU+7momHnP
AfWOvq8Z2bTVE9xUnqt80mkWg6KTCoERpnvFuuYive0j7zQP/n9XdYXUD7oTaaH9
0zigML5TMlsIyyZYuQQif0r5K/BFQAuLW/X2IOZTXJS/aeOiOFdJyYGjjOHs5JGM
aC0kPnTdHnwXNYccHjXRzCObI/Y5XcE/uLxlsHw2StOisphmSWwliicQ/iELbf6O
EjfedO+IxMP/rZbZKbCY11hdfiUVM+qdYy9k0yZ/Ks4gRclKP34janvF7HwpdQdC
0Z86HSmkbVnob8n3JSOAwrOP4lQ+h3QcXPTCiJ6EkMsixyBNzgtgedi1ZKXvdaIZ
f32l+XwsMdUH/tGuxw/bNkZMiMfrckTqR+BgLWIfyDxJcjQQ3GoCugzIWWFM70mF
rikGEkSaNqBt4Hu5AcU4Xs2CwyT7flIFSozRZjxt9P6n0a4VQZDliY87Kxow1MGK
Jjv2+EPZyrUei9E/dWDNxXPLYnJAXyn6iTaItshq3rO29NW7TtOlU4tHSFXxymdw
MA40RfOuwWANqcIEu5sgj13r9f/u0MDDFt2ikQDhIor8IM+aPd19KYI4CUcCfADJ
/hzRWzGM/ou5Ofka8cSQRJG+0c/n8JIhaPH/38jABrvKaeaNHsiD1jZyHXcweewu
USykagCtX3ntpwTqJGUche8OgOBLlSup74kwtt1x0r5at0K92zEVPwaRPug/BFWd
UMDFO1LKIoMk8kMeuWBqA3RzumfpPPP6qbV/sDPcxBm4WqtxSa2OzoqX9yvhYJlO
BGYL4Dwv7n2WB4b7+v3UL4pqGArFVby2gvhSVgMT9wuCp8/rAjfWatfMFoEp701d
+uSOXLU2NV3+1gsgGxv2u2TcUS0aWzDyvofUDQtzFe5c6Wxi9XUyte746YV++fZO
f4Dmp/8ibeUgEw6mz8AFW5MPNxpIyrmpTXENHo/Q49WKLq4gXD7qr7cVLM1CpOfG
NNu4elTavAH/f04Ja6O7Zy+qNLXRTKjO1iMsqETTa3+xiXDXtLCyEqXJrYslBKVK
bmwKliqtHykad2tfHQnGS26JhqVmHHSOlu+JQlhxvYYDmqjN1Nod8nr3/RYkpIqy
Xu9idpo9m1iMzaoqCtpA2sWBxSUtqkUUia+kCGYaC9dPkVskPHVgNklQZDmwzsaN
0q+puQKyqDlq7pPl0xG6F5h3ySkQ4tBoBulNOWWzI2Doqdw8YHBYThIenAtlGM/y
3etiAtLIhm85KNC+J2taQFia59wQAG+nRv5NFAVE8gOQtWEOZqH2wC5NOMHHjEu7
eUzPwXB8zZPL762L1xSeUXmf3le9uejIhy1RE36mEeYdlKwNTqE3ZNdTrykewns2
nNAWalPioW6oOVwQ2Wu6eTdVP8Y2yzlo5iOho+NUcSeUH9nxgAaLf5zOLg4XRl49
RSRxPvyi5JX5UzI9JJgMOeWmVbaWb812VKA0yk+uXIVYHLmXPOwKJP1cu1GfhVZp
uF5n5P0U4hxXM+rMezlEduZHXIoWcrReaTBp8s/TIIL8GukqkgkKG2bT9jI78dOR
ztYIiX3wW+vfQiUSsPdyD/r9Y8XZgFYK+fOKScAnjVcVN2SYpYZHe/K9ZPkaWV8U
0Fvyx5wllC8pOOFDnHdm1sBSztCIVtHU2C4SGbqauIu+05pD8zc1cPI+MT7fvz4L
+iqC3kG70Tg6R1WeoNgtG9SOT0Fy2ui9+Tl6Yyca+oVCyOCWg1AIs02yZAxPoQXB
yDd7oo1cippAoIFiwwvebW71mJAwcMu6m8bo40mOZpz8oB7hcdjZAmNSUhWgfak+
mlEldVS01moijpjhVY0L4lPNTinT46nw1St3OZoQn/+Br0bLimyY/rqwr344scqD
GJM85VhB7vO+eZda0Ycp2mGvW2EkXW9ZgQVPlHQUB5oIeiuOGZxyxqcVsi5H/5Fo
NFBDacHHy92QnOFqE1z/qNfJoNoCilVam0ZTDIqp+IbREO0K8hB3OvJRWKr1ercR
BJh37VBa3CYZkxUDpf96Tsj+ibdBMvrrBUwLy2fooYTqNBZdH59fq4KgKt0HEoaj
2Qq+VrvSJiV7Z3Bzr9Ol1b9sg4o3hLr6PVa+hODaQN1Ib8Lx0jb7i/0IUJ0UNu1v
OOWgUzVExGKnPX8u4AtL96Vjv/uFU1kQ5InYVloexp1Zu2a/9nikUtK2HG4t+OqJ
Ah8j3Z8t5F5NBqxpbyqf0h9EvusciycLKZo6DgM5DW5VAvKQEh55QNSEkGuU+8a1
S2BcuQEFNDuEuvPDYw6fAz44bBjRoL0bXlQz+JKK0uKtpgpHgE3LDOC+hfO29mCr
5RA8GhGMI58iT1cDmUXmU/0uyhk921lN76aUBtK1vKjbVBt2c7TdtjCsLwyJGYAA
wLz1mZd4c2ZoO0Fvv+d0u9Wi7ZN/4Yiclzuarbu7i2DO+lHiWzvL5iiuf4lZg57G
FNqHDrxrHTrxcyDu44D2TP5WPECs62tD0ftQ6bTC0OfyvY5aW7CID1Ss8OcGuH3d
ziYHHTzM3cN6PSZWSZpyYPGn5bdnU0Gl4HYQFJMRvg46AXsNBbf36uH2Xh3FFyQy
YWdz/w5E0AuHilSzQjphdsaJWHeooPIwirmBaJ4hRT+8aBLk/6VqLGnUfb8iqlpU
eJAygyT/vQwb8G4ledIVfbRmc72n4Mps9sAYGqm7apAm/QJtAJdESC2ZHPmV7VAu
mDji2qrfBycEHsbPPIKkjcRzYxavjZI3PnqEorSwoCWbzaBY6eGiX2BCM/c71Tor
rZ9oT0uhOJRdf7Lqu6UqeHc25HEgxYe7pDatj8zT7kgZVHVGLrgOhvnDfX5448fw
7nKWz4WvKy/7MUJ0Yr65rEGQeRFK3rPEYs98bTzwoVdqY0L21hTC/tkuopgA/2eb
D2yNj6jY/RcMYnLBWk44rUd8zVXFsTxV6v6BioJYzulXPzLdg9EBBxx53SPRAsjE
7IGtmgFYLho0qkulgE4n1mu5lbQ1TZUd5y966vH8spU/cg9JcFJ94FefGqKnHj1h
J5tgzfeu5AAy/hELSiCAhfFdaQBs/WbDi9d0rt9y7KnabCs+Yup/tyWZ513jMN0e
s5B9ee5ohw5i6ekwXkGumoZawR7wYcaYFSmHq2LQ7yvZva6DSKS4baUbyq6Yc5fA
4lpYs22Ds5+q2nPhvi9LOqu8ys1Xzggn+tJ0//9lAL1573jRcwH+6KdN46KXlZin
G3y33ZI3JwgB+kaDXrsgZd35YR0hlx7vSrp3/I34uBsqwGLMKNJ7MFBIYNcuF8gJ
Lz1b7uARyhAM8foj9OLnDWvbPZm2Ecp3OHF08qoeFKyY1OaXQS47GMoH73CZV8UE
Cdqts0onstMIeWl+SvB33CrQ570fDNSbKiFuiCvXwA6jP+ymy1vQZ+vfeeFwBY9d
vhoRJVOuvRHK+dyDQlHLZtHwyzpwmsVus0jXL1OHH7r+1RkmTKaDAfiyIAIfrrHY
I5dGAKB5wnTThYWAaYy8x0UPwz1HzbUkISAvMDBA5xYxUYB901cV4nGSk4kitv23
JWPkMsnw7U2wOFUex5GXc6t++5Tm/WoATnaeZvZRrcp5pz2x5QkVUsNE5AaWR3ns
p0eAUNc3V8HUqz94By58gK9Q/nf6kBi8aEIaYGlE6C6ptSjWvRjdr3FJcOckUip3
Cq/kxub5aYUyW+ZIVvqeZxhKkF3lAM+mcifXIsQfCnrQDPX5gF1UxPlyagodgk/X
Hg9DNTct0/ZXF6fqtKcjKeRwuG9zvk+O9zUaqLqRFxJhDv+rVb8SaDWtkMgiz59t
OwZT8ni9nkIR4mthgw/O+dy+g2xpKMKq0WyVekswCb4cKyaJsJhh5/WmWeTMK7Uz
Q4FogBjDSZXwnmsggNou+OeOQlNnLsHzZrZO+alO1kyooyWDb1eyzhE1TzAcblGa
0cbONs2BQBIW8ERCZdSCS4A3sB3RikRS4c+Muq9YKOIVGTuNRZolF7RO89/ozX3x
PZbxjQwS4MkNGJsrR57KinVr2wJc5lMxsxn6VbvxPIH/RAKBEs8IFxjyILRXlatW
zNpSWEZtIZzhekNNklXqD2TyjWavg8UvKquu+mX0t84+Rst6qfYJNIaF1AMF/ztQ
e4dISTFiljC9MHvWRfeuaDdKSRMG41PhcHWLKI+l6XAOCmAw7SO9lkNMi19NR+ea
iOD29LNrPul5V+imG6qqC318gig6GKvKT0MweEwbTsYxLGobtyFSbj//uTKdEhuS
uGC+ujieDWaq4TuKmfhAch00QERjgblSIYs2O8oV9D6QY7uh+ACxOLHLK1xnZ6Jn
SaYSbbjAEuCanqKmugloA/8/5Kj0FYMK/z0YrlwLz1c1uzCpXj7Hoi2nbs2MRZEP
vZlW6VqYGGZsOu0h4vH67emo45oNN64ySTpGGgA2XXoGBYj8EMaQWRieUPRC02JT
NAsAat9SQDdSHLHqkLXfQA7YA4t2ny4io2O3LysSl9PgGaYSn8HY+vBmRT0nMS0H
N4/6UMeWpnn++r6W/WGwp+DizFc7pFaygt1EABsHyu7N1TZdEnyY1dFosKIDZdtc
O7iVKdDv9AugS6oZksCjfaDM52OQb3PLHPll3kL4kHk+eJiSyPifD4nKdFrlHEa3
GL8XjVSqslXE+UdJwHXGqFov7i1ZAnUWzYb23zUPPtFR7McBF+a717IQSxgO5m8d
Yk5HagdXqBKHwCgQE0Ooz8aPMMrfoiYO6PKEw3aCjJL+HA+6xNtG3r65+yW9NF3F
u9WiXp/Qb7qj1YmIdonuUvHThA0uXBEX2dZEzhfTQ7vHPIqKtBJ+5qQjh/TY4g81
K8moq+Tn+NS7QuIi+vn595FR9t1lKdSi4UxuxCIRKW0VNPhaZJZsg9X84lHHTRNk
gvIZL0lA6vtnCJL8fIdTaSuY9fjwyGDpL3ldjDhJfp0qK93MCQL9rhUEProIBJtC
688LLCHxeNw+z7YqtP5XwBRAvS0daBKrzfzGgiKEe5MnwJjw6klFJRQlSOdJ5A0I
7d7nXtk95dchL8UBTBu4m/lkDF7vYPApqt+F1So7muQWAH2C2C3ahRDnjojFu87Q
TXRb0rAod+T0HtyxpQX8n4rxCsadgWDRqoGWNgW55xgCOqEWgHNqb3Mdeghg3914
94oKyrMAf12qKB90oy5IVTnry1FSAyeIqCZJfMzF/18NzKxmW7kpqzfI2eAeGM5b
ty6G3znIgp3kM6fU4lJMchVZHpesrbBSuRL2q0XV1pMM/eissivZ9f8bAsyFZEj0
YEIOn5seNPGI0fl2iA8KSBkepijoO+p700eNcUk3mWqKsbIbrxqh+3RC8nYosuwj
pXwGIy6Ck2RxiVKclDdUFHtzhB8TWC/sCc2VcyD6+4FsR0acip5h9rqbEVHzGNnv
maSHV3oItpecXQxqVr/hI+nK+QQni9HNI+VNV7RWz/P8TgTOtJ1aUzEgdgQMQmDA
66RZiobZSgBja4IVetibdXydxwQ09FUEw6b4wjNCC0maI9/8E/0yzpsK42mRDxKW
fFqax3Xe5rSKEnu6zgOFeUlK9ezNsWUa34Da/vcE8ZiXN7t/GSC9Rl/FUq8qamHe
opHVgEwB4K1OTXd9zH1BlqmzkDevDpMNJAx2K0W3SCzUeiT9xY873FmB6iR21xHe
qousmC408LlZteUNT9Y1BeMrQzWrjouYPjWxzEHEuqPqq00W9qQFGTuB/5iunHJs
1tu98Ba39IKsEGWVEkLv5jNAQq+kUdzbIbUhqAVzkCkNFLwagnY2A7BlwHgFVG4+
Pj3t9lovcrPsCch1TlhhLMA7nA0PZ9jQESHpovsYyokVwUHkcSefgNJ2pBHWOzS3
cWD8ab5VMfKniIbY07iqT7rpMh54EINTeyEs8hJ3/crlZzXRm9Vl00VPwr+SCDXU
bJ80OZECn1FF5SqnVqIlXHGJpwyD5+rqXnxnDAakdmhsJZqwIfnVoDKJOO+eRY5e
VvU2QnFg4e3dzkaAuU7SH7PbGahvFW47yZEPygLFr7SBsOul11J8sORsOhr/zWOz
zra4/j1o1QEaNIPHBuGkAWECLNidzwoeEhZuBg02iZ1sPok18HA0OnpGD+AxUVUB
nJHz/aZEgpdmMpG9WjS5dp9rNsMaonlblHfdP+1In6AQLyt5fJTzvVOvjEOxS2wY
iABkEwbwVvsd/DDKL3qI1VEBH2ZaYUsxh7zjtWb0BlUkdxMD0VEKBJ7iXgQN2hYG
Kr9YdV5gQVnRXgzG+xSTUVbqEha4/8aw5jOntd8kVmB4k/kxOtR0R6PdBn+Z6QIW
r606FF9Dwcf8KUGo++wXeq11KOMpYNEtuc1M7YJL02yvAH8twqBtiuGJvN/J9kHu
sgpz1SSKzee/z0dTqyXOw80ntZKE678aH46NVZHyfzQjNwhU3OOCmK68/1FzfEjN
hkNtDsw5SuXJ18Fve/uvL5RswNox9UbG4si/vFhOj5gb1WS9FwbtopMiMWzNWD1N
NdMzh7TExsqQaULQXCvAP0mkEiXM/Xu4y7HaPrySivfsjuEeF+WLvj23+f2/umQN
COXh31Ecwt6sovZXn0pbVcbcs0b9HHN76cr1Rj5f1cINxyLfxBShx6WXtz0OcW3U
ispfANTCFMMS6DXqo2/OWMWI20LDiMTGAqShzn1N2X50LrbikX/2EI5jm4DvquZg
V87L7Vb2FYsqP33PSO5uI+uBrAGLKB7ieEZuGm7Plij0DIxZxFPOQ0W+VtlcIBl4
VVVVR4s8q8XL9+y3C0zPexYrjAAyby0h108aJq7Gyllv8hb4KIoHmi50OMlLqWSZ
prvFO75RB4uZTeDdQ8XbJu+NGvW+7mpL69areg7uYOZCMeASEZR6V/y53u5wJEfi
99Pzn5wxk8lNKVNniK0Ece+hWffMv33+xF3ExNoN46NJGtV0/6VWq0vijJKJltFj
nNLhKX3VrFXWwIPayNcE/HEZkqC+UFaRZ7TL1WOXedJ9B94PVCr9KyVn/IBV6XF4
av56kvi/YcFEDDxFg3BmgmRebmXnX4qS9b9z7ug934WAHXJXvOCGPpjPMExIt2s3
5nE9nt/MKN2kdSF55Szg8vA6nTck+rGJ3IWbKKDrUdPorQVM/9OjW56t2B+5Cmnr
dEoWEEVD1j6lrjmIYHqChpvYoM4os0ZNWyu33CRjnaeG69TOC0dCa/C+nhqed/Sq
R4zDuLTTmMo3TvE3UlpcJF3FAlFOQk/4e+KYYG4C51LrMuwfXzIf8O5wOk3IQeRI
hmAPaFsWhiBX/fxCSMIeITOexEbZKWvIcc8geJaHN3JCMcd2wP+8j6R2Rw9S56no
iz8SLWZ08xGk5jdufV0X7JOUBevV6bHPFzwSLonVyBgTwjAWbPM5a4cmOLe+hYnK
cltk2noB51g0B+1ZeVcJ4alO4Q7X9t5ju9/gNXoFK4hlI+zfrFQxn3S7PqDSlwP3
Sxcf6rbHNCasWxB1AFdycAL66nPvS01hG5LoiQbwqnOX9V1B/184I/1hqAGyYVo3
DItLHaQ8K2+yPgulqxF2iYfGk52giVmXe47YCchL0XESjLYigPvVuE5/R10Zf+5+
GzyVbDBV0yknHr+m7WinEtIbje9vhESki2bsB/fsQem/kFmxU7Jt4VdOmeeYHuHx
ixnVVCuC12sIisnL3hXjzDOxs6lMTJ5xKNzMjBvGg3zwxfvP8r6RAF00P/OkAgcw
WUJub5Jrqv0SuXMFQ1f4+He0nPdc0hiDSTFQa9h1K1V3F2YLPegODhXFlrDHV9eF
vigimAGieAAKUdUrvfTmgfvvVU7RtvcwFvEdVNqDaBnz6zMw2AmWj5j5mIuKwaxU
gPxI7lEh8dpMUppTqiBrGpnmH6kuPM2rrwz5KHI/1Vutznybd+tBB0adQ3OmK76X
ZQ9UvKXPLe5+OzFsIC2X/mW2y4AxazHrzEYW+DU1/0DZrHVF0wjy9D9ZyM66K32K
Pw54C4jDUQANxvxGChLiaN8aR3E/19DSpMN9HbzJVohKfOGPQ/D7mrWo5pVgYgF6
Oe8zTFSgVcp2i0j0FL/8nPhX6pdUlljzyxTQ57kOLUIbvg24aBJ0VS4TOSS8fShO
vifXlCC4IIhnKe2ttLm8brQGyEfXm1GjZaPcE3Cl9As5tPJ1aIQbOk9k/hOEyYmI
vbNrEQE8JD8+IaIfQtGfcpAxxFxOhJIzbWMJy/TZe5pXCs8y2qyom1zlsMHeEzng
irUs3CAmMlm7zfaTpgIM/nFxXgElNHCsvZvek5dFrZZ2mPJI+hcFyEHGeMdt0Fgy
j62gnfXm60AWeUaB3AMu75PvPS6wdcLVhp+dGj68LO7ZZQymXW4sT7H0H6ceokKR
q4JnIUhw/DAkej7KVQmuyy1+xmmt0lblxJzuGKFlEMxJtuDjtais1ZleuH1VAEji
JxnWMsnmOPlVTNxUXaxV8Kk1aBIZAipbpqIZ2WRYO5zqfSTD/KJUjPnYLgNwtWFg
EJXXoXuTaavuekE4pAmyzz3MdBgqWZWKxK8yjh2ViffuA3LE0i3M3bZY1jLiKFlj
UKm93WpI8tk4MggzSVnHS39QS1iwEH3lY8WxAi/Q0TExyQbrVg4nvgMgy+iq6Ewj
kCpWWXASAyiGfZT08mt8AscRdkn1AFIJpgAk86H4aJM2sLim7mJSnzKrCmRL6mby
D9giRJhCr7RCzaOoU/HFnDxpSKpawuycgsXbZV2gfqnAQTwKtVOxMfj6CrQXjo46
iBN1/6DHtIio5eqQmjczV5XM+Qk3pGOEjD/zPT0lanC1r1XaN+wplOH01zGeCXVk
JNQSbN1ls2c76FVM5e6lvIPF5UnafEfeeuCgPt3+q4S3jhSRENrPw500LyK22iY0
/wx24ine15jBYN2Gslvvcbfr1mZAaBAFjhI3U4AzqUHwZbOio/OzSONgmhVJWqWy
Gx0sM9nAlj/xjAZzu9RPH1ZJXLzmKqeHLM8NAC9DWeNYGDB1wT6hhcyM4kJmkBXB
/5/c34OhOIzNA3FJmg0L4/0/kY4H5yAidCrrr2n4tQnqaTtd6k/iIdK5FguuLXpp
ntcOyD2C7/Fw0SbnsnHnj0z3oz3gqG1oXQyFs1W0YkCD3hfEkLab6a03j3QizjeW
XZHH0cLcdT4V0nLo5+qgRX+qpEBshzDhkcIKXSMZ0kflM1RBMyW5Tz0mWoICRhTC
QbZfi8Zx4bLK8ri80Kc3tCrDqSz8LhYacaXBSK44Uf+pR55eY2hwC1nywCRoZXHK
/6e8C8mT3yQOrVssn8wZCilPj8vHjpIq/9R6LlTP8af/H+eBnA+i/xnAeCrmThW+
s9bUZp3dm60/veZuQRJeKZapmP2hbrjx1geftkYk3tds2yw8oSL0hvt6hTXXqJsa
H3vSNvKXPaS/VSwBKBw5VIYFA3grmXkfdR1JFKjdCXPEHFOh+MYOTDsWRu5v5A9F
n9d8SDFZw7PbCa84PNb6GK4Kag5ym1BFq2apiQ9YDwW9V0lWd22t8ud7fpuz4DQ/
cN3C8ByHXZVHk5IfkvR1QIrLtwsfDDABYAl/nKKq7k4JDn3t5Pk7herZB0k/uD5J
FQpg5OlEHcuHDNuUX2YeeU2OduYuLdvClo0iOSOstaH8nhe6yDDO3buRQqEa/TRf
Un/fp6AB/7lPMOE3ybR3alP7FxGcWQ3jRi7yh5nx9yK0/Br/dKlq7O5ToWMHCplp
TDObNHgqUK1n8LV1H0qekODnXr6Jzo2nlTlJsPsppeoJXohiN/AlGs4ykWDfRGRZ
Fm0qDPcnt7J1c2W1MbbpTllXFzDWoeh8enkC3VQ5VZcF5bDFgjXMGSl851PMY3GD
quwjuoAdD+YbRmePYhhrxdDvo9i4t/WNigV4738ZKWZSiaGbaGDIA2pcy2wV7yDj
nVL05q81EwrezdCDAI8uMDpKqynI5LoHTy2krBF8ZilYoNIVF0UkTdtg1xS1yH25
H2PvpZA2coQzcsOEZSy3JtESAqNIKgOf+5+c3fVLkaNQOkt/Wh7f/8CHiNidvqmz
avSl3IVmuXTjgjK6iFD2X+wLcB9v2WM+HUqbgnKseVAT46nQ2dP3uyhhNektx1BC
PA6DfRkhTePJEdnXWqi1KOkV0NTFuI8EEBrqqvHF1FqyigogRifc0xUUdkzx+ToX
AiXU2xTfBSDM8QgaYJAAP3gCFAHsAuxSaPe1D+pV7b/EJSQVcU0D0uRfsjiQG7er
RxPGqo+fRgPCZanz2LtYXzvai7W9qyl4ypaCsTyULFqHglzGYHyifS/4913sgneM
cGXUPj3lS3mKBNg3JUkZzl5EQPUXY+PiVLcxomKMkUjfuzfzAFF4wKhQBu/HDv4Z
4+WIlEKMR3m/35MRvmMxscmb9kJKw/3F0aACsaagtBc+CmZskO7S/beIOsy+BmsF
an5zk8nhrksKqmGRcA88G6i5JrhCtDMWkgwdRD7Y4rDlVXJsAWZ2isGHdSO8jJWu
JPIR1dSeM9aPxcAy0Dm3KAo6eh67iYPifSmvc8fXRqnX0shOozrXXHTaM28OYAPZ
T9aRGRQQnO8B24uleRZMepUN2IDaq1cqJsCYrpIv8D9M5ieSFIFMU/AIYQt/Z3+D
83RxVEj8LSxc9PgvWMVs2PxLFgIiGn5d1jrUW9xtHlX9+KlrjWFNjXD7NBuSHqtr
iJ34RZmfLInxX90YlYfVCjjDKPpkGMKc4DzqrGCK9OoDJB/IR1pX5p5ka0KVKJXn
GwciqahAnWCPoNldprNv7QFrV/1vUv+LcnfYwGdooKQ46PkbIr4oiGOnMD/wP2YD
BmPAj1wCtu7VtBtaDPpPPXFzyt5833V2s69+5YKP2q551/1cT/hFbFDnXP88sFVu
WMZeU0U3+Oh6v2oCnRY/QcsTsU7D08iILTE/wB5k2RDu2jL87whCChqobMIGr0DR
S/yxiYIfmECxmkgbSMAd5F4Sgl7jIxVenfo9qydBDuuiOQHqk4rg13QirX4EqoSx
mcCSkcUfnT4ynp0Ehj9ScjpkLJdwxGNjyKEHgEx/go3x9YvBtGLc17yK178vJlDQ
fI0J1L5yEY6mKqVM4S2TCiXZDjA1gGZhfJAvhj3lMHGm5ecGL1jqshhF7e8w59AQ
xdSDmQs3Gvi7BMGGwcf+RTUVFmUNnXAxdlyBKFImHpmjjKFdIMeVgyU6r983KTAv
RNbSsSlr0EadXaWT4LtHkn1AyDfgF1qiBKFDwUiLgH9PKTMjrqp3gpgqXmOnzXaF
M/Rfxtbi4OJT2RQUD5ZDItZKMEhSdN0IibM5AdzVCjAjnHPhcyhZmCSA4xx0LIrP
Rnb278/7S7GMTbjTG1LOWfDiJi2VX9lsqpToQVM2oTI0WrtQLzH9VyPqUWelQNgn
fxpaIWWaSmCmpnbVLTypiPA4SBcKx0Ad/EeKAFI9X+M3/5ZeHmSqOVpPCS/5Bzbs
zhJ1f4kHyI9sP1l/lWLjmisM7996NMXZ3F9FOGh6FqTg+FA8pB58Wz60AboTzM3G
AOk7aOX+O0Lt3Oqkmkt3DEBBInSWwMjZmvvFqIvg/AHgbmGl6ahjpM7bG3o+H4+p
s2U9se2m0y/P3vbkaJFMX2arYFVHeVqkk4nJfmphR/axra4/3onPT9CRCdYLO1Vk
bLkT7TGPBfbdAbTZ7PvS5Zn4pv4UDO11kUipUrHkZfODSG3VGjtl768jHWLNNdzW
DyPVkTDDBdpLRsSlIM/ZBWBwp/x+iJVN+d9mCwCN+kb6ZQFDAmAcZZVUwCzEJIfS
QEceGATwoYcubMU5G/ZNdwwNfXZD00X0bjnDB/yF3FRGLvUkKrh6U4LyJHOyv91J
lb5AS/81WxtKcEp6hkHZ5c1ww6WEhQTdElZqonjcSaY7o/WONkvKQyAfcnSVBwn5
o6vWYxhsLPvspxk+/MZulysBx/04t7Uxpi0B0bFHJHKSD/Nxow9d8oyRZqaYm6yZ
fKfozi+2gLpxnJj74gQ/8X1wXQ8ArC4u+viM/Nhjd1HAfpWQNwcfJU9Vm8LxHFI9
36FcaOJOJ2pfl0u7D4v2wD88wtiXU4HeUCHQFUY5NRtPgbidkWzS1D451sXpwPqF
udAeSLWDUfHCj80AEjF0ycKOxq0bYbt/RaOp0jwLaV3JWt7ZuWx3pCBTratUmTmB
gR7Ugphv0xK8nx/9rGtfZlp5+58QT7IBZE5Optq4UX9phc9h9gEwU9/+2C4/KfNK
S/ZP9ze8eFQr77vy5R1b36DFYMxtxNERFus0SYeswJrlc2HM/neKWtZzIq0XYFiA
Vf4xvgJjH4/f7PWjS6jt6uHOEWUJ+3cbRiGVLgltJTS53mZEDtXTV0PZUwaPzdMn
Frvfl9lDRT1TxkBS8iHHdU9bhEMWANMhZISdjYJTFEWBZlhdo/FMim9kWv15y3bD
lxFDpfklgCtu8J9W4qm9nbEWLrXcmo14eEUXzJpUgIa7M/yGcZNt0f/RuXB05v55
O2B4keaiS+kN0ljZbwdke/iEQ5/9/Y6GgEHlLHP5Zx0DssI9QclkQVqJfvMEqOOR
HW51REQ6eDoekxk+7XnatebpXwR8dIhuIM0IjA/pyQM4NrLjdqZoEEhBF3PhOCb6
Xa0GY7OIU1OaVsIAJZQDdg9cX/1y4QIeOXB6tHwvEgttuckxCZ5SDMIOOPf8LPl/
DIlMcJPXZYrHWlw/HQ4oR8vzLHetPCY91FGFCmMuLS0LeWIEo9woL3hLyxlCiz0i
AbMP/wrViWw3rPfjRw1zU8vVaxBLcVFU+HLeheEY8i3QLy9FREnpCr48VknZlAkY
cUh6Q50rLAlY1khpWyJmQ6vdjsWCxeaK4Z3FZrqBJqFGnCQLf+UjdoTYrmuY9/gx
uUMrKKr82suZc7nI6sZEOqTbXg3IH9Bhz05qZGI63qV2nCb+O5ilQ+zWJOfW7188
EoNQ7mCqrgdoGaQP0Rt74kZo9jlVCD19ZJGIRa0UN8nOJ1ORRiK47Bjv43EhdKyl
XciuozH/4ERLVDgbE7bCxSFy3SU/0MyPpKajLXhG3qJVVOQU9IvBwoPGa6JDm+0C
LoAMTAkHWZGS6SuQFaNAZzl+sHvYNX0xZT5jh7ZS3jqETMTqLx/GhH3pDKxoXDht
6sGAh4FWD/APWTk43/raMDRrhOOVTx6R4SPrr6qbTd1SmvCvg9eqJVSQbYXvnQTD
MyMnrrigog06MDlXmtM4/6xuqFmEDTI9L69OIL1qqdi9EJ8TVs9FrdJrAjOOgXjA
G5Kxb1gL/owAOnlg3vKxH2jSUgmZ9NycGL1sfF4s6dbtm2hLNBe4XOkGUlkklKQE
rII6tFnz8rh0r7F1CzHq5MfxjJkxrN0qy8o97NruHjq2m85yTKBv6ZYjhq0eCoRd
tHGWR5kKXG8SpsC7VwAc1PSGgknQkwUc0kMhV2kYZbo6BHE08xAA2w2mHdRQr4RO
Jycvupphr+OMF4dij/ZZxjQtWosgSd+kyDYxgXqtgtHII1cCh+6T2wH4MBwldMe2
dqWNyfJvtkunW5/wKHAQTHNxBInFpPE7+vb/2cTZurxWGGl+sXFD5fPMaUpeDtnQ
9y/L5sjbL2VVCWppZsX5x7toJ9yJJlNcVuYB6LagtM6HXXfCAHqByuwjdOVsHWzN
+iXFo4cYPX6Rw2Wb7camhZWutoZ3a9muHrQrlAZUKMoXgYWMapBHzITmYT+S9F73
/vVy7BXd3xHSScB9MPErQ8UK0mo/4LTdZp1iFBmjiskYUTo2Khsnpobj/y/GwjAg
JDDRyYUZYYDhobxLdf0Hog7dNRLmZDJiHJIeV7k+uq8pjYY4ME/NptzMMKJWNgnu
Bvi+4c/LlCuouqUBiOrxiihwcwpQSrdv2ffzoq/W4IYblZcI0GP9kDR5y+XjY99t
CfkRR+zautAXwWVDyjeh2rw5ziwGp0S/ZGQUYCoZLNJ6Jv8AzcBiokLgTDK8V8Jf
uL5E5f9+9KTjTWWffVhYvwQAG+EIUdEV5KmUBadq8AXW4ldsmlfK00qURShfEMQk
YUUX41pBejSZ5XcDUujAETFJB+R6ZHh8F4TuKGAcP6JRXXG/aox6GL0zg4wamhJy
rnMh0eoe+jeVlLCzisI8MGxjVt8l5x+3T/HTf9uz0H+VIqjKW5JqG9MTqVaNS/sN
9SmJHXabd4EF6KItFX7CiWXd0OkY8IKDAEqYDzuu3SgcK0btAB18lYvgn6Hd3FGI
Qcn84UzTldj0jrcJSqmpAOdU9XCmh6k1QRRNlUy8ZL51ShrIQs52ZxaC9iNChKdE
pZThV0BlaGJId2UexUFejVLlz6yBwa78vmofzZILXrcgqltBfuqA9VEzCkxEywex
VvQboCX0pgPnprVmQsT6TA==
`protect END_PROTECTED
