`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qu88Jezklf20JBYbb/jZNK8W8tvrjRMytmI3RqGEyc72qIrjyn9uncgCUYvoOkt
qw5WqLCziHX5dXYtQZAzd6z9g+JuMj7D+Qcybucl2FuuekAQnBOkLKB4QD4D36kY
+e3yQUbXtRsBii+SQE0Xxa3cUKBSRCq+M6Pk1Fqa1DdhFw4YE3Q6wjvBhm6/8Vpc
dYF01gBe01f3sIr6M3bnGSX7j5sIp73FnXmNR+lAoTu4y6qeXMnsAaEpSHMPdEwP
2vd74ybUjLp2qYq6R+P/5NULe+5UTCOSRMwAcnL77quYeBAufoZqx30BWeio72Sk
5DLHUw2QCW1IeyH8rP/qE0Fmfdb6vVznQK1j8jg9LU09W3pGJHm9MotqZTSn94TF
yMSyolQzknLfJPJGnUh03iXpgY4jkV6N2ZW+Y7EVYmOJwsdtXWY+CDb7AbocAtgo
FXMA0wx1YvzR9DFbL6I8a3DhzkMAq0fOf/cQ1dzs1/18F0h/MF9b+mnhyxB1Ch/j
ueqg/tKumaEUjQRKtSks80mH1vJTqfohOMW6UPCTRomfND7lCO/c3S7rXHyltPb9
W/Tm6a2FKDTDN2Ru9RVqfCtXPw3TyPO7j17hxY1tobdn7t1kaxlAxxutc51nnm3W
iUqMafWREWS5pl4wLc50eHt81G3lZ/AlFJDkGZm/SR2GiWflGZOQnoQXakIVdmZh
7IyxQW5oY+nQPjMtnihjB2ya4kJ1QqBs0UntrOPbZarXzhRizc8cVlWdY3vi/L/Z
X25AYXKsNjumYAetBCc0ecBAHDtvW5s8nuoSXUfZi7atljFFtR+1nXIpK27hdORI
HiSY+GxBglREgrLyNe7XeiETRywYHIg9CQi8uuyRfjGDCP15Vm2+QyZsnyIgIoKS
RdnRoUcPO8p78Wn41buiUYw17YHpZ8C9WWmxvjjbOnlYU2IBCVM7kFThof0pJpy+
oi3r3Z9ubQ4Wd77fJXuLBb8Afkq/kfhJShXa2bKXfIU+48VCq8++zVJhYPdjc5c5
puFLo1S4kaBxzIe3PSFLg8nQo3EMEo6hye+MAyCo4/s50VAgXUkqppMEyhQX4pD4
+ZDnM5Nz/tKSeU/onl5/F0GiyY5Pt0TVnm3gSVNpAFaqR6ScR5HkFATMz16+u6dN
ucgEXg6gm44G2WA/GR47iTpE/g/lSdLMcIunw/PK2qrbyeWbJlsLPq5S8cgpA5AL
KICYh+KgbMfV8/QdK76B4A/VKXZPPtMjmy36RmJ/wL1yGZ0MIQvfS/TCZVOHMvsF
5fXNBdhAph3aRF/gateSDAdguL2tsA9jdPj5EA4BW01blhhL9j3SRo0Z22o0SSk8
GqLxRIEZWahFfOIUQAJD9XPVhVf+C3InUWa8Y+gB9gaTu2OuBenxtAZv0wwHX4yo
tkD9gdql0/ed5KRbbg2dcJWL2L9E4dGQJLRyClcWz6WYact7yiEqf62bnbzXuq6z
ry1pdkzqUh1a7+wcobRRAS5/zATl9kFOmj5D+rnk8rBuXa5wVRTbnUYs8cTUDSHM
XPycJCvC/HT4/mXErgwcFKKwaugMr2Ap4gGTJ/nDNZ6LzXcJwr6LdFCi/iMrdSNc
UUUyFlwJaL2kGsJQO3JjxIGqWKkg3eItzZFtiFN3C7og52CC3xKT9v+EAanJYzK0
fDM9e9GCONye5Oed85yyylnHhl8oqWcsxUjA1vc+sKDzkR8tHJ1X/UVjrGNQaoUh
/MJ3VQPg3lEWBtNdgg544wXtPHwqaDskxkCknMTR9gd3qPQMkO+8gXTIhgnt+3Kl
u3wCjlRaNw32bCOKyEOrk/9rG231vUndI8nA2diRfuDY0Qrvmgbu5mvC8/R3LV11
NAI/NnglPyhmnDwDRSZqvVBJrGvfg23IwkvNYh0W5f90z+ZAHoq62TIqOQGeU+Qe
BQAJF5jZCj4R3cvs53TCoMo7YmX3O8G/8NbJdioSukGvzzYYapR5nmptqpWHkXhZ
irVQ6q8yx2NkMJioJUOJUJDjRhdxF++WVW2DzV0l14bmxTUTiWqbiOYCO5bxVZdN
HNOFuAhULnGo0yvo5iu/oWw9tUwiC6PriAsYZ9XkIZyvCAbDZgB1tXCXBG/IAcJM
Zh3/+8sJnRfmPmn6HMHkrUM+epWzG+jf2Mxu3BPH5iCmLCS0kFxDI3ohY5KW0Nnv
wHeI7N7B4S0HuLkzqlooR3LDoun9NhCMIHCWf7QzPjLdZfnH8mGuUSlaR32825Tl
BviLmHlGgeontVSxHw+8iBDW54ss6kFt+Oypkn9C/kjjUK2IIJ73766FiZDE+58p
WXRlm2ZTF/t0bbtKlmc4ppVaeqyz55Il1Ppo/Lm6/1Zxs6gIZZQtLsfr9Ekr6ayf
re97BNn1rJ8GQfTQJBezS6PH3+S9x2qKJ3VlFoc/GS8hqK8STccvdDd7HNmXgLPg
TEgZ0r9Imp51eCjGqo3Rdr90Ss7ZReTtPmMrBImy9V4tb8R7QqInWHV/g56H/In4
n+6gMb184BPM3sKZMLPbkjgRP4S2hxYUAzMdZIe6+xCG9X3SjPShU22vn+UIm68J
H4K+z1x4AdPgz4BH/pgLQZk1ezV3KBuz1h0IC5hi077M0tEK9BX4T+2h1QV2XuTz
VOO7HXYsri+1Hbe58/Zto55M74sJjH1oGQTbp1hl9xQ=
`protect END_PROTECTED
