`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H3c+TBIiJJM0Ma+J+HP5Dmx6YFK3889FZBQPSceLvIJf2joue+5R5YFtW4VcbHvS
2VCy9YFZIOiDc678wnRhJaaFYeL4BeSwNSoAqhjJ1eP20EInzGgc2G/JIrBR1xuu
FtYvnuTVJWOOaLwtrSFOGCkQgoxhGdzw7vtvxGV87NwvDaECsQe8cDKNiymWivXV
XU/AbZKVvleo4kyDG8JVkFZOWe6+fyf07Kv2XfGFhlRonl0e3NJURGYKqM+jtNDn
2bhYQwJKzsPjOIRJ4McbonKXbuD2lEsjWKmQO3BFO4A40mByzSXzJRHxQx4axSNx
tPBH+OwKMOihyZFdeQah/UqdKBmi+u43S4Bpy9MljEK9vQHUuOA21ptdMRJzQsMh
YfCCPOyOfvTetUugYY+XhbtNRXKbyevfC01MGV5yfb61ZEYt/MmalMcO4+e1wumH
DC0ir4tmTDb/H+H0MQX7yjqKOULl2DHSKSO22/jDM1fTxnNMhtLpGF5kZW7IdeaL
6Sar1DtMBtpBGXqEr1gnWq/CHrAYLZy+HknpEO3YjMMPexj3TP9jdnoBr07MzJh1
Y2yoNqS0xFcn9Fe9pzruynGrHOvF97+LmdsO0F0W6eXvK2wMZudBv3wwBs6SG36a
+vqsW1glFpE3Q8Oy1SRppMl1eo0B0sxtNQPn2M3h7u3uFi4FgIeURIND4qdfejWX
WB3O0d9K/1l/t4HusYE6E4HtZUg5Nl/8+twCQMB5+udh/26IWFzPiKbpVs+UdBjh
Dwk8toLYieeBW1HXTUhXxwsL7VWl9l9F5B24ebZJ4rZ3nzPrMIXJcZj0IIDqDu+p
3q7X4gsXmgeccQp+/Y+YAeIP9BY1E9UAamXDFAUxNfDcg8xtMxqKZqPD3SebsX0W
q2GizzEjPYlkXx4H9XlqhyFLII65OclQjtK3uSfJG7D7hYcrZZLIOv6H2Q8wvOuo
ljNcltRnk/5ZrYo+MzorDS9+m0fH6C+ujhiIh1JackzefqXDuD/YpyQj4RzqdtH9
/AwW5o6++bWV05SanLkFL1+bFhVpZShVTDWbAb1W5GQz+LgOxGTDowPPPw4/4aTM
is8au/6uyu8GKtzJdwUP1XGzHeVEte6l4EvQAFuwn/kr+dElbTmScHX7qcCZ4PcZ
HJYYsryQ3mTa5KdlEBE/eck/WPqXWP2vcoqZDjosbyGb19ufOJOcxgtsVglLRxii
WUJM3gYJNnope9xs+Cc5z7T/AlTsjxk2ggY5YwSGSOIsbsb2mhJFPkLjjPM7l6u4
xUjM0+u+ivtabHJBdU5Zr9xOlZNlzD54feZm49GYE/NzgW48KabbzG5b2X3S/xhv
/eYTlIMrLrRMu30Ro6d5sEjAxrFk96xfjyMo6sZ//NYV2RlGSUpA1PEWaw/yfzuQ
HeB7QSVmwYOP4NC+e/gYFu75pm9rgxeO2BfR8+E71k+HxajdvxPp50o7i5WCI6Mg
xlREtfgoDNRkuEqCxLg+tOuaL8W90dIDI06pfCcTyEMJwC0d5V2uh8O+vmZWXTUX
`protect END_PROTECTED
