`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnAjU2nGpS6VozFXRgEHfQeWiUoCOFZMbz8+L1SdqGw1rmnAkm1FwbUgDzxGVVBA
IAOR+He2srV69LGU6ISLRELU6UbIE2lrgb08uIiO0gucUUnre7Ksic0CmqTVTAR8
ROgRcLhQ1CtvyVMiM9iAxmkf4GvSDLuTdQLBtZ+DhzWibUckVEzVTnBiE7K/Gxdk
g1EHPudo6JtILZUADsP+mBFO0NX/mdWSr5B5CVcKiP9xBfe0pUSzCB8bgZ93HuTy
EnFeG2UEw4+rF6xGTRLXERfU4UGxsQaqvMGsnOkZ9d/67+RrW38zb7l4yRTiFb6N
EHbj7tQDHwcuIrHg3tllyAeDmElvQ1YEXeTtwjkhwZp3dgi0mnR5A55zzu0P+Vjl
GehwL+PZ5BJxFqiA8PdXX+e9WNQMG7kCMMYrc0BdXYiOFhSiOXarYQyGfnPTG2nM
78om/l6+0uLwkWHKAye9VpzbsDXizVKYx2NF3utETO0axy3VgGh4yBwyEb/o7bnG
g+1Q4OmkBzef4e0yMEkYkom9cVGyu/240/buvwYR1lI=
`protect END_PROTECTED
