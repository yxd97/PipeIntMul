`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TewXgXWu5wn2EVIXkwYjc729pwkSRCrwklEOyoNEOWmsg0ZCkZqTHUCi7UoIeG5
PqFM98I0xB9cVuk+CinDAQNIBu6LtS9s36bLM5iaK1dbtc/a+JU7KZY68KGOgIOc
Z8cDHWLy0zmOIRyXvQLaGaixkyE33eMZqJD91PSSqy238Zh9aOy5Hxqk1yqNrVwB
FQYYS4zd1w6Ow5cndbZDLJrfbK4mOxxebwVz5Xfhx9694lvbfNDfNLUzMW41u2L0
rl+P2dLZe7Nf86BsN62x1Ah0/+5axTzWpBao8V1aDqA9ANoAdI3NAeYM+oN7/HkT
kVwQqTpzmWH7LvxPtk0+mV2DFGZVlIPnxT9j7tz23pQNvUc0vd6CKocwh+ZmKhEV
`protect END_PROTECTED
