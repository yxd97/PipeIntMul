`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Fe+GSrMQzgJXSnG8FIRQLYg94EFZfP8IW+vH2J/iefTtgsskPXibnN4hgo+kzQZ
tiRM8UQf9CE4+9rCUEy4U3d5NDKpa9l/V1w1UANT8eHWbscEj4Oznc+PtnKXL0lG
wE5aPcgQ3bn7d2LCVD7JhQEtZBVaLM64mldzQOCx2G13ScG6aqbcyeSgpaYDoLW1
CdsvT8VOAbpCY5uvIDzS7RAURpiSdTsUJV1Zu58x18mJkdR7/6Gd5xiNdgZd0mJP
5k6OnFwLceD8zvAPgf26yg==
`protect END_PROTECTED
