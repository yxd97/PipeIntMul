`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aQ0OJErq7v1nlJD7rPL0Uix9akbIahBhtXyi5gudt1TUDCLiLoozFpO3qCLkVUvz
gcbK/3t2yeqTS95LkyT1t8YAW0R87BpxIzGY9CWszU3igW8lqfXjrgDl1lFmqIgK
Ps1uJ1CBNDCsmbSznKR8v1bvsWTz0jw3KluBQkJZ3NyfMw7cOtcZPTByIKF6jjU3
wlOIWFuTHzIl/slkrB7WcPO6ZUarwbRLEgJJ63XnfCi+AYdn3ouu5ZgOwffMMHNv
k9B9WWPRy4D5LVEyBAzbtZL0mYGwZ52UqMWHaWjQJQcmksI7TkM3lFgjOGpka+gG
DoeviyPmn6I3SXCDkImPAPA0YPwGUIdNu14JbBZ9c8VLFYu9ZnEQOTNJBhasy+Mx
HU8tpl8QOHuypYGzElKacO2QqFGOJvJudqUh0T9uwUG7I6vKq4wf2Wf2DPWMvJQC
CSl8qT4FnGk68y3PgBDdDavhAIQEVg3G5tkPjZcaYxgkMTlE1plJtssfWCu75KZn
P9U57Bh00mYQNak85DeYIsEZDlBuDkiaRrWOp0+N1pJKPeWDEp2+CimXJ/F1G4jb
SP5+POePGqYVNy5j7OOSKbEx1p+9iEPpXaZoMh3Oad+/CUihK0qqBj4Je9irpdEt
pPg/1PZG8oX3l8/mo/SO4REX910vyufX0I6sPhYfxIMmo/FFi44Ftnd/hfOgFMRV
NdiRB8oViFzcIkZKlG+/vg==
`protect END_PROTECTED
