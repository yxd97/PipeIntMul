`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JtUFxaXYPjxDixL47YgSXVMSJ3jfsIqsyi0rcT5bz5rd0JTAHWs3VDKNgQEJTzAH
4acoYsOXFTX9kGsccZNTjh8rQQec90WSTG1AiL1hbqPsmlbeQ9TSSGm3pBxIYFhP
liVx7Z4zwLHjUx5UZ6enn4uAxRn+M166r5a/9uhkDoGu1CAJSy4ZrkVoDolBtK1J
jn0Qx5iAcdpVDrLfBKmjfcd5FX3uIXZVEbj6iFjpsCXjv4mqMxUmukNNRfXkqvoC
/mZG4GLcrQbLIi+Pr9kPe6a79cF/VHHrxg/2jA9P5oUZyHHPwEuXyJ5heGMtNqIb
bKPzQ/fiWVOpQLSDsH2b5qpcLKEVTMhrO2Wp6G7opA6m1+xHqOdMzP+i0EmTaFYH
xMCulQaMI6ctRCFHxPiEH67AqwZgyR1DVOzVdl5avy5lekkTBelJPjtH5ASCl68z
YgK2pWDEOzlUG1wyiw6xEus9mUTQZj6T2UL7zaFj28wxBeJa94HLy2+lnO6yZRN6
4QK6y8ah7iMLj6/3EaRD4JwaVfkNMQ5WzJVEdcPSewu6NcWNDv6Iw7URscCFaO64
In/LBDkAt0Vhgk9VVIFaNcAHTilsq+fbhig9FR07OCVLLp59zejr5G04VF3Fptbn
X+WtOHWne5tRD+0Q/SzMEsA+GDBQj4VZe48G2WxqivRn9ZQ57VNIiP2a0VxL2aiQ
B79prfiU9wfbJlic+zv2Vg==
`protect END_PROTECTED
