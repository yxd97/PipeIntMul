`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RieD5vgKcwNnWG1FvLGqVNidlzWVjFVboWxFOiXlcxO4Wy8BBBvig3UnyahBzqvn
+bAJrACkKWJChCy8UAUbvmdroGdbKLoSVAag7a4meQmzktUh52iHzar44ho2TJFS
9sY+gkiAYmAvk8K9c9rZ0IBzV4uqUxDm4XO1UoMLhuSKZxN/NC3QUPOHMOaZJ7cM
qD8N/zSXhOUwVbX3ONROIdTTDrTcv4hHkK4Gyd5pRh4mM4qqxSOu6kfoJZqsj5YZ
YPM8epHtQx0GtbQSqezEGwXsZAD2Oxo3y5ACbNAgcVxO0IAKDLMM6WK6jbOC6peL
TwUhiRP6xD8lflYtUARX4opEIMRutYbVvFdevOm0napmzouWy1yq5mLVBSOKC9oG
zmdpSAVfJmPVRHlDM4dIBpGcSnxmiRJGE4rUx6tfD3Il5HjXBX7G7ZR1nvylqq5j
2XPC9XFBcwGQwYo2My1iB0rRgA/YHba/W+ALQ5QHcIAye653fgsbzThLqD1vIDNv
JbGndHnyf++P/0YCM/cfN6tIVmfXBGhMNTcZd7StYo6jGsgmn+TM2DLHCk4mSBwJ
D97FiwhKcio+j7adormcshxSLjwq9qdvCqYILJwutfKLrfTRlDLVw4CcVkCx70ZL
mPNG8C5BAH8LHKSKW7AGu8FD6CdbJZvcDiYzoJkHGZDRIUHIXtFsrEEMPT9VtP/r
B45Gt4fEP4C4WPvwoqYx6ZJiAX8CtqSLuYK5+WEn4B0XaJOyg8Jyrv2T+VkJLzcx
I0lF3JMw31+9EY8BxLLJvfqU/wPctQk9Q9dUjKeFFTzdWtKqk/+FHxegKCkm5/D3
WohOt6i48MJMs9BQryR5FjMfR9OZM0tG7JK/Md/ACD3D89hSurhaC6ZK8FGMkjnq
NGjdjEx3u+G+4pTYKtqttYmmEO5kKywKFIuwLYY5JUeLG0AtLzYGRwQdz83SSF2O
wzQ5fah4Q8XNR1hIcPV8UpcA+wWkqF0KrO3J+nomFiBujI03m+TCLqrhbKVf4MpE
HRad/uAJ9l6de+TGVuOmWqmZpZDDKAljzwVvXEVFbN9Zrb5MjiBehWb/C530b1/Y
FsPtFrjEzf/yg/0tGUp5r2f+fwf41xL7+j8IBrTjqpwRF2OVmzc+xowQfNS34wW9
SfiqYQA5rHNHdLOyat+OhdvqNlDJV1Pz5L6zO9j48kZ9d9+AeEsZiNVyGLjMrg9X
ifZpKvsyyiEotOkd4Je9YKliC64ItVBaS9zjUSLBlosC3BFHrK6bjMN0E9TNU0Ce
elR5exCycYJIDQjEG2LDbpB/GLCBsX4LcbzIF4ovcQJ0zvvRpJ9MKLZVR/sG6RgU
J7eJ5K+YZ2aUvqr0DwT+gcQj5ZF0D4h90BEXyLdH0QbVsY45kt8p3yIyn7TRYiiJ
UNutVMzdoZeLaM2exvhpO18skzRcX9IBTZKMyQ/dj3Kehzbe+oPb1OuhyCE3ZrDx
Q80WvLkNQ+D3NobtyEaqL4EEJW5qeli4lATXyZi2wZGqSiVphKyJrx8nPJaFmLvV
abit8GNMvdGr1w/98H8X91vZjWflFYipEJIcg1G6WFKOlp0VBapaMOwSyLFJspOT
P1F1ja7R9NiBV64zuA+kh3/AqwyocRPQCdRhS+mGVomwDsXOO7oR3YB6qNMWb4Qd
AWnVQrVUMyQ66xYM4k/+pRYe//n0DfgJI4Z61nwAmXCj1cCrLaA59i0pTPXQpzKF
zF4/VVRAe/iHJnjq//waZojHTOXoKuiIMTNHJ/328lJUqRmQ6BdA6L4O8jgjUlp5
ta0ftOKUjmAOGLx4burFdcvXmHRDSQgX4nHTYsnUMKWZenpw+/Z3pYPT1v+NvXYv
KrZQV+Pdm/OZS79wUu18k8OaDWSWdfUzSSKwoFDi8VIreA6e2WJNttLPA7HPTyOi
woN3Ktm9kdaqSbMFgLhM5FRfSHy7Q4RWHZ2z61iz9WBQY8LJ2Hav0FA9gz5qeEOc
acgjMWZwiZZC9E+sqR4FPWLNLhbKpSRvlmsbYViNnwBBbrsJXGHVZ6Cn83ICMsoJ
cMovBvfX3e0UhF/RrCoUe+e5Kj6EqjQ6dyjEe1k8/KWgI6o9GrKxNlwnLFwYYRKf
gODRKVags2BkPrR312E3OkDWz9vxaMHsXaQDx1CbxlbOENXYKWQn+0L9Fb8IwOVS
3Q246O3Qc/7zGv5QEdeHbIAORHB52sEf7tuJOGth68hcaPpq7BEYJYzjeP+H+qTG
fdk9ZVpq15eqcVkt6yJBfUCLCtyw5fSsFvgPyLUDbzBSfdFldSfeG0SlzsihfZo9
vrE6AyWEG2wna1KeBAe2WEQVK66s5l7rOIupY/rXButHrLS6gn7yf0D8ccFTRadl
veE+rkZ+Eqxf8JVlsuOPg7xa8GiDDWP/vJZYld7J3QBvLHO8AgvCMoacyIFFMhEJ
19GVqItT2luajqWAHbmHBLhYJIdqpTrLvMad8eW2dA+F29LzBS8ZZeLFUogHYEXr
NQ16B3ouZgU09h7bCNoXgVB1rtS3CeD7rkUDgZ263uPvleGIIuHf+3E/lIXueYy4
VPwIFIebRQ4MpwZneyhAGDgQ2XqG4MTeHgZ3Kk9eNyhhIcGaNXkvNyJH8/BIgduH
rLK3GtmO0vI0HMbYXrav1epN7P8Ni/93Dc9a3ijmGFr2E0yokWvfjCDlDG0Gv5gm
jvRUylIPYlow23ExXrnyuHb7rZ68ZLouYuLEFICuppBsJZzugbprAQIV2Tnt2Pvw
Sz0LnKtZjPvU3ZX5BSWgAVRWUQLVvf89gT6V6F5I6VDcp+I8ISTJMiv2u4SyXEJf
7DEYCWpVvSAHGCpd/4fT8iC1cHwx8wdbIUlkHRkjWajfEMxQGTbxWZYObbNIxRj4
B8QoSqChexapV9mchvAkChePCDFeIpFKbCrJAW4zP9Wq3HlFSSj5+ARkJ6HyZxRF
aPvLx5pHgW3oyU5VLSbIwJDDTKSmDXnr2qnRivcMOkdYLe2cy+aLlZ0RNFImPoIJ
m0cEGk9m1cCPH0j7Iq0d4z4Itu6+vh/k6ByefXGoYhzHxSFlY2Vjy0PjOPkfNS7/
VtqZF5/IyBVyf0LJAcO2l6781gNbk6tPhhxZFgYdZKEF77H79OkeXPn++5XVy2LY
Yne3b93xPeCwwnQFWb1AngcRHRrlddmcfCu5M1Zu5i0r7bKqRUWCTmaovQmZNdCT
6g6EsVmkQzMMheHl0FwFpK1ViCRycw33sq6sHA1ritmRp9ZP6jAi82lGGlryBI5T
mzaUujr9gSBsFucSVVaJIM2vkURk/ZKLfdvkMfY6zRxx77qFu6nVF60y4UIIYIgB
cREYzwaWeBdNFdw4buOeqJivAals7KNiVYP2v+DRVIAp2L6QwM/ArfallRQcQJfU
QBWy+WrpgJQ8YuuGTM/g3pR6d7gmRAsMgEIayb6+pnkdx40fiShO8zcNlPGafyMH
yphYc5jFFjnnEm8lVqYqddAx6GNvStQneOMBUiuPH2iK2LWsClPtKu6Y0CGhIHHn
eFi8XTKHHFBmVOo7C4Ps7IVXCRIh5bzXyCFFeLkQdaxpSbNGAJ0UwXMgri7Qc+Lr
ZrfNDPP8a177DA0bucZMJdqXcHhYUwuk/Y8p94J2XI+jZUcZaz6ZcPQEra52IWsM
CK0f11cahDznRQBEpXFY+FSZ0/avk9p/6hfV7IJRTxbIGPNeJvCCcqY3hHtzJ9DU
7SDEBAafHdMwIot3BdO/n7W++FSojxtvxm+ShmuQnAeGoE2irqwsaJzBbrsWAzZg
xylsHX+y6EI5Y3D6v35Qa3mRX/otZ2DeS9mnDFTPYCzi9LTcKV97aW/3A6SG7oBG
UtV+Pp/Zr+qKd/aqb9ENQnLA/dbjXyjQrEEaAAwKusDVfYP6LF6bWbNzK57kGETa
tcTsKHak5PgdIoi59Lv4iXtJxXmJahgGKcFqer+hhvSGhJoZ/cB19exCtMXCsT+d
A3TJp7h9E3n/Z28knTP7iyE46XgW2JKb33K6T89GAPh66Zn6JbpfcYFEvT1QmVnQ
Nu7AXTbaT7tBkA7PDbtiXPYjREqX5xKtOjQR0TSgT+4ZB3PtwG6Mhb37FASLJdpP
mjwF0bi6pjcaH5aCb+wGaU5pu9Oqy/gk0zfrLOxgIwXcCqaOs3H66/11EypDY5DD
sSAjtYllm45My6lGbq85Jq0wocNGkQvLC/0d/M0eGtbgELJwB0wflrg3GMMEHiG5
KFCOVAwjNAKAFn/M9yZyaSxoSTrX9t1zTbiYmzhpaf+++LI0qi4vLznPGZi++kmx
RGOdQK1bn464m9LQ5vnARRHLM2q6xHSUiidBf57Y5T3Pad7MVo+c8723avhx6gUs
W3ZO7k8/1GoRnS8n6sAfFwOUFhUC3o7idItMKZ0y6teyhKmCC6nJ3TxnRI2CqcOw
EfFX17h/okC7X6zjpkeoUgY2r+kH1Wvj8mViATLVVUIGuUu0+uT3aKyuXfDoZKOR
aHHaPW2GjNwNIekvB5QWpnkP1+ORMD9XK/632NDLrUnXSjcy6eM6SW0O8H7kbDXj
t7TxP5DXOI4YTx3OnK0SywaPLoYdT/aW1AqzRcqdlZ7qul7kMHfno5gydWyUGqfI
t705QYF9zVriGEAPP9aPmkGSpKyvzg/uhAuKsDBT0XGrzinEp7WrFn5j5PBC/MMa
a6YynrIkrIDmIB5hcmMqjP7hpVYvKMXS0FRtuApIrpqT5d1bWMYTbYRSrTRo2o/v
L1EHY88gh4b8mqaoAIZRb9j5clnZptQJxSi95KxdzmNgRYFFKWP0e2/GTdr3a3JU
pfhKeXLJppJTjpSjoHThksmkemZYEhZWs8YiJ/lJfWkwW7Puj7uRg5JXlLSXgIUj
xbpD0Eakizgf/ngWRuE1FrTpaz/G/FW/LF1463AVLsc46VV7ow5dmAG1WNksG4OD
j75140IXk553nVulRDuA97iY0hmEHxXBLPrPNVIJkcmi2nNXvkMKpIXs04SX/DRU
NQnPjlq9g3eRY6FEdAcBVO8R5Gmz2+WbK9Uj/Zr9Y3Kk2ELpFmQBqn/e33x4GfPh
Xyfi+5NWD4vSMaMPvXPjy3HRaDx6KmAz0GEcW9wdTYbXHxZ+PLNiLoEyx05w4gHj
Bmx+roj4VhJpV+0pO36uWcFZNSzlrEGHWDNJIkUQMmORN8eIc9lxz4Ru8DJrcEN+
j1+/zE1ITo2HWi+8WVqW2Ox02kvdrsvVk10NRaEFKdi1M9BXA7V29lu9KieEmxgQ
4bdBhIe+7+N0CfCcHTDRpdm3Y6Y94053bXUgAB7mWTvQv9mcNhp12Q3WpCF+vEPn
1E15U+nUtlrrIf0pnDVh1foH4w+MALi6MYf4qVwJ2xwQyw5bUqsTkU8Y3+FY51rA
FDcIQj3eMrOOFOjw5qcOqMYydSti+Igxsp4GHivtMzUz3ZYLZ7ARxuAXgRZuKzPq
ht4PxDjWzQPowbZy1QLs+UKqurpw3OhUszO17+hTleyKnShqgpEE+/kPsZYgKatY
CLzcKL6u6IdEmgIuCdWHGxIMVKrscttFVHOjG7isBYPJNmZDyqymZbPsljh26Fe5
0a6GdkDmFZzu8vhbT7dZJ9Jx+lhRDm91+sZNk9kFEkia17z1q1pvWQZi9ut7pBND
2GF6GeXPsdmstLFgE48VBHQ5B0IgbGUEkPnJVbRIrulK/2gUbCo1HBRRBqgYc/jc
omHbyCoHtYo0izm7dkHy6SAGpe98xG26GjeHzfE6LogYdlAle7Ct9kathVQwdrTd
z7afVJMMd8zGGgJmIsKtESRzmUsBvEZfiyKU3QYlEU45f/mDjMcm98vy1Lw4gyrV
ig98opb7X9x/7hwMI7y2hu0XHHVK2di7r2nDhwOPS8evlJXk6mzXNihnMk9w5Ak1
TeY/rxIZ1FfJ/POv5ag4xB5Y4zCphv23/fYl8IXIlLQkapewg/POy2r3PMH4AfZg
pc1g2Y2NuttyoRrA4JygMr66jrppFFWQW1uPuTEhhoYQJcaXpT9+rxn6JO0HC7tO
P/gx4LOUM/OLTCxq/PHwJRzpCYGiENyS9mJ5kwd20g9faBeaavyRjjnm0RNOIRw+
FSh0vg4tT9PVIotaQgRzodoHiSS5V1NzaTKHNiQsKPoFOAgL2t9KSO5tCCxkdiW5
EoGriwp4LDSWCPqZEwVLjUw7StLdbD7zpmrdFzDtH5LSWPOyjrre44tRxo+RSng5
xVYb/6Lf5eRsMbeP6dzfEWqALQpe42bWRL7CRQD/xeq7mZqcj3V8faCBfFmTtsJg
bVPms3tbRpDMG01G71cHgq+6nhMmi1iD4bSBNU7zsYhW8HLAbc8pAboecNKsOJJa
5rsRMZBnYqFowjdC6sPtn5u2pmr8MOjRzuz0Fmi7NDAKPNippwK8x2JMsgqZFO1M
j1eNDaS8WAvnn+Y1GA7++ibMwYE6X1r8YdcyJ07qRgp725TxEI5H6GgJbTo+QGLL
5zg8ajdjsuww/OzRCUUZn6HRjf/UlUd2dV8i93O9Q2NHG9xliaYS/a98IN7Sk59J
cETkmmY9buukxF3jpIN8E7BFxsizk7hoANsIwXIbOjG8oz1PKV1PwFHpEv6BLQyA
G/tPU0hX2N4jq7jGHwGrW/W1s7zuR6lXTLyrEgQXMHRrrAgmkGPrJZL8YlpnxWuV
r2uESE1hX+aRfX6jC5JDbOFatYA3r+ol2Uqs3RtHYpfstInlcnxBRqyMMj/sIeGL
6IreqH2sxhAGuSqIraDgaiZedms7t4isTLUFIxB8zh7xklhV9KooK0SzMGw2wgLR
Nd8nqFbh5/Gbt8GTd2ZqB5tlcVzE0VQ+A+5tVYKvYjg1twD6Xj9gJwEx+ZH3+acC
DHqK8sPNNJ0tbNhdfgBKcG3WfLGLJv18hDimWf/ruU7xcqhVoZHbsz7piJV+SAzG
SCrlwB6lXpcpWJaL6AqAMyaoygi7H5V4mM6VP7yqG1xA+yh7bBYvhWHAhwUZHTgT
Td5dH+FqX+hlvdlz9FZjyiDmDTJtWVFcKxiKS9MO/umhTSkDzkZbD+4yhQlRJKg8
pSfxY+8gRrvRuZBXg1zDsZYTR8WUC/LmTcb0SbNw65soQFewIrPLRYIWcsSt6Zqa
nJ5WAZ5PUIThG5IvthYUgUx7Ouqq+alQRMrt3/p/nFsY9GARQRvRexADO++mvSNO
4sHD2GiLCsDgRAZvWLIh18fNrdKDCpelbDbVfhxwv6qTt+9WkcPD5kkdEoLhZurt
sCUP0GwRl7kIDfA7tj7I9e/ZyNeKwnX4uB0lpS1Llw/VDlLp9lnt2HWr5UynDMUv
0tsvqNfG7g6U7RUOHZxX4+tTK7RKmsxFXIqRTIWp5tTisXF2murnoK8TpGNmMcoD
0GFBgxasx7st/9c6W+BsBlNWO+3vU3IIbxn5sSuwUGlu6f3YukVy6Jv/cbqujFL4
7UVAlt2AYv6itV28a18Z6DS48tVVWDObhh153lrIrrnFR7Jj9+8CquJEvJmrwa2z
fWcJLCwxpYsof0p8UtNcAAtjO+NXQSkPg03bN+R+ptDRzWjpc2NuTpxguPlgWi8Z
ZyTSXs0iAdR7RVWd958Wqq/V86MQdX6RFGFRzYYE0355Vr77CBWUUpAY/gYAo/CV
vtCnd6MSjXZ8gf2zNBgDPL194wa02yMzbgZGKNtkffhbSet00a+afDmfZF70SEON
SAeTtw4VBC0CatozirlRr8VpEUluU9R8hV64D0J7KmYefpdO2h65gZvULbEW+DkV
ZUonHZhzDS2h2JwwVSuRdGruB3Paf9y3aMPZtjIPL9HgUnClt5hKFulPIuwxMD8Q
z7+UrIguuFqIiMv6YrDNWLQfgQLYEprSpxqWnGDdVwufglmWSWfmpPkgORsAbx4a
P2t16iwZg4bXrjf7+iDOdYepNjHA2nKYQVXMMdKieC0=
`protect END_PROTECTED
