`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8oyneUV8keHePpM3XfIPnv3kNiY4oRdDv0W4wY7oXrRi+zUkrT+d+Wl1PedZj4zl
ELPog3NyUQw8CD94Moc2Ao+QWuqdBOnat6NFNO46hyGiQZdcGHfj3qhZymarGUMH
kxikvbhSqSZx6OqsHuGciDrwthzklK5+0uLhpQbNx/t82HePM9kJeoX5V+tbL1kF
1Rl+zxtU2K761YA2TovLNmEKq9sUBhjtHxSS2dTCCOfZv6FOoGQ0pyC3RWiujFEc
uc8maSt1eyebXXIhrVWj+yifigQCumZ/hfBMfImwdk0vuvwchPcNz8FN8+GMbmFE
aMFJ6KIPQcDIXdB3ANE5iP55sBo3XBHHUvE0db4w1tS8Co4hbvZGLsPvp/BqSHnc
XTmMIbel1qIvfnfCNMoR3FzAMj8RzVzcQ1uzh8weT/wbgkw26dgJXZldXfN/odsy
8rTz5x+3anEbBUPm7uDZULxpGAoCp9+AhibaoFanWQA/gcNg5EdzAbximR0UxMuP
hR/pgEDkN2eHBsKYDgyL41GXVEgbcmOcTT0xQUmeHHd34wjd/TNoJW0PMmpSos+r
WT9tJsfRKQTpKROPp+sh3S+McFNbbS1VAQ3Bx/JvmBXgsEPG+llbw7UC5A84GNYt
GyW8WUauMOy9PckrmW7rjcPZ/i8pib1J1yql5GAIEdVsXdTsd3gTWK+HYUL8KnAu
I0oZYRZ52wsYJU//j/WihTiTp3e/+lvfuqmdDDo+n5fCW7Db+CTCc3RpWEOSFATC
+rHss7aJ2Gv50LFT6e5T2ncnuieikm/tPSg8YwFAgeQZ/rCuGyNjfT5SX+uIUy8f
H3BhsexqqUgGWwruv9k2Rdqn9FSx3Q4kcEWHuqx7Hbpf2jGXd3Aabdye3UVNJOuZ
XHqno4Q0Tj580mon9RDvc/JwQc7yRrsmlDRQrWlkOD/HUtBmn5HnnNE87zedf9pS
8VNiKMsclLg7EyznjkCXO2WrHgfp33xk7CWt7+UpdCgLQwxMD/VI0h4q9ewUdNSw
4HsCB994BI/HQXxRT44NF0Q9ylTQ3a2DS1qEBoNJAqLm9UxVYLC66izlMXEMfYp5
kFhcGHpj2LsLkbUBt8+f33lsoW2eh3biimdn4HS6k70BB3quFExZCwxq5o8ZD85z
8+eIJi7jkv/Xjr7W7PeolHEFyIxQwUL5PtaHBkKuetTbI+BBEfLZDrUK96N1sg4v
bM1uMG5IO/YKWbQfKKLpziPyU7jtNQ5SXbvC/eNgEGkFFbkZMie/Kbfgi93Mc3og
GbxPUFcj0lBX972fzG2BA/vaQxXToVlvbuEn8KrNub54MrBSbXniyx9t4iknvzdR
eif3x6rvQ7Diz2zKtbfhT3MhZId/S6srU5wPVHW+eN8wvVzbXz+Nq69LwZt/oTfx
OhPUIhMBpatBs7sDxNGyK3M1n7pO/Jj8GUOKeHDTqzD5wF/wE1UAGwwQLH5JdBga
SL8UbXz/WUH0euyXYGaHw19R4KzAwIpQNsF8IvC8Bxvy/haqW+QauS6i2Q3477pL
NZagAVsNQJiL2Ujzw2HKW4AkHbpDGZWwFiwoVnk/CcvKfTlUEJi+3yLO/uS50iSP
zNmw1lH/EM0Pntw2DgVyYRSuvzgwKVG4tbLax7bMaiIes0AnrSL8SHXdaUdXm8Pa
x2Ux+HrugJnbLbBev0mHNXU1BVXwbIEGGegZI27WgY1rUHaumdEWeVNmN32Wza0n
cw4w0S0gouY+Pp74vkGVzNPl1WODAnGkglNCEq4y7XWvBnjHRxqOjCTfyT7++0+y
DDX4scwaqDlrmxxse7CMluzFUK4Af4aK/oUyDd10lmqknHSfcJjR2+mIEUdU8xLX
mJx4p8gltAn4rL9+XL/LfGPotXIyQB8poI00+rK9y/XvqrdbGDIofdIyodPqp3dk
UedTAwzKKjD8MsbostMtK56OhLwDQyCj2AbGmSmL46H+EqGemJPcvOqOqmgyh5fU
f2JkpHg0mVgNWNPNmiTVVOBMIGFJh00zP2cWNmkQplRcEWcf0aptPGH/k5izX/Hz
FURNfRnT88nRpjJUHgEPdnJ10oOSKF7b3Drr6sEM7kNl4r0qrNi/0vECdNMhLl6D
5V0+rJehNCThYvH4ydmhIjDt1I5QHvCD6jnsstq637uu9bsR2Ig2b9mAztK747R+
7m/tLML6CGuJB3x6LFawh4O3T3mrjNU1+JyrQGdR8X3p7FUUhEs2/BwYuGMkk2wk
9k1XO5Aap7zM9Zw6LqcMIYFn75GYyE4l5cfjPacJpFMpmSRVm2gY8Y8IbMBXwsJz
rP/8BM//4+GOk45x0StZFI4P6t3CLA1GIUE3oqfTPKNQF18KUdt1IRBs3AX/2IUS
g2eh2bLVluEAwxe/zqkRhzfHouwd3YNHLspq60O9sv5SHeyXRKjXdP2Z1hYxOwQt
TYjUYGdzg2fdM1PDp1pxT9MPJObjbMnKtL62Evm4ZeyB7nszItj3B3j3NRdcUIMt
tVyjkgcqLsf505RZ+YCc1MC+8ZJc2iqv6ycBbnY30kDk84s3y7//DyPd5jzRsNEt
yyIr571F18yvNzTdvl0sZAkODh+Fi2WVUj3CSZaW8VJLl+LHRfWzni/m/Yonq1fR
PItGuzXX0u79RcrfFooAodQSkg017U4bVZCslg3Lni20istEv7HVfm33bHhoodhS
UMBd2GYqIbjfuv+4SeIk83RH0xiIBN9paGk09bxHmuQW+vZtYHgN4hmtOimJ2dqb
H+c/9lSzDfrJL8mRF9GIFjqMje7wDefP82ylCU4BZYHgWMRGMG/zf9djVMu/QtAl
61PMoPMbsZ8GD4U8n9Z5djiYBw3EbOdNDVuierI7gLgAgR8V1iLXI2gdebqXzGtP
2SLnIMWW0nwlAhcj/N+e7hdgJ5T60mp/PnWe8UWDXx89452XcG8k5YbXaxl7Az6w
+tU1jHd1Hyxs6W4hxRiE9Kz+92DCkiI3Knl5x6E8uijO19gF1hGNxYgU/MwZo0cz
rIUWf8+88m8J8hPifiNn/Ow5b97qysrjhkAGyIVj16c7po1kXycpX7z0nzGo4h+2
6edD2pcWJoeK0Qt37s5OOFOJZcnGXndAo5adkMqWeC6iX5sP9P+Lp752ny6zopTZ
4Fpj36Ga5TydILRetaXH8clKbjygsDl56uGNINzdX5yNGgw6ZZfSmQJaHOM8bys6
3DoBz24HbnhORiVVxVfY8jZ5VqsoBa5im5wozOXymDJEWSNFUsE4yA3EzqEekJaR
oTb3HLileHUH4v5xw2h2dEBcPq71hu2uzIP2cGYYDtohZHrFmFesBPe3eEomBx19
ZgkrQsi9C2BgSSpIo+YQae9/V6wfu/PDdM/CoPairJ84EOsPeKv3+svP1Pn171Wg
wa0MUhQXfsQiV37XJvcALpcCawZZ1W9XSk/qVJ4ABAp0nUkvjqqlCAXxp62Xfnf5
MOMvw8SWeqm5BoDgK6GQeNF9jw0BVldyk/5034uo06XKf0UV3iueRlqMoLk2RjTe
PGDjVfruusiQSNxcVcs8UbiWm2Rf0sNXb44Rk0MD6yT3iBrZPsd9MS2nGMFO+gn1
5tONIM3FamXU2+PkEqNVS1IKfT5hnLVTK/7Q7pDybujhp0xULkU9EUub/xhu0hE2
L4Kf6szhY2k2hpKNRemLjn8wwGThRn0MT+ZMHrtFCIw1qHhp62c26t0b1/Z7j/9y
7tP+O4PMfFsnLKsXTMYt01arai+ispGaTh+ZpRF7s562t7tzptT09D7AH1CUrZIA
Bp+wqVyJ2gEax/S92yvOkM4Hd2W6hnzFh79XMcMD6vAp4u25SPDVI+hHwExUrh+m
hL6JObHQVN/0UHpmJkwY8AjxepwsduYp0jIStiRUHTAaTi6XNx3fkzCVzCvYw0eg
v7ezesGC0/lYXRhFYx+f+XB3TFToBox7RaBc0uZTimEJ1MOzZeQKIMQtZhACoGYW
xS+MaDEam4a0KIiYZvi1X32P/7vCCn/EX/VeDHwSbn77PJHM9+kb90vC0Pq00T/E
rJCsIgOvmwZ2s6DpZL6nNg8WUJiWOD5sFFbdWRaGVPNvYVecGhMgQI7mEw93FnpF
VpMT4Gk1Uj7pKWqUAHOZ2twvg8X0vCdPDwtml1vI6yl0WXNT/3iq+gwby2JluFlJ
1ilkCCSOQzw+chSWDfntFAKcZm77c43lyHk2oXDWhstab4FXBq016gbud9nfv5/N
hDE0x1LgYzrISSFLHeAVQdpcML9r3xygzmPEzOU4gVqkh3kzIu/yJ/wrY8Q39VDX
VXLROoZe6gxnWl43ZS0wzkpAEn24l0SD82up3xo2CJLeAEK6YRlBQaS89Ha7x1zt
4ORiXqxjWM3thPjLArmRwaI5CpahsoH2opJh4a11oGKkOnoHp5tzVD1nwiJhHyDk
MWwHDj31CVs+DZm3iCTfYJ3pkrzqn9xNfVeddhF/4xjCjSgQFgMyK+XK5i2cbcVy
SQp1Nq+UVx+9J8zi4KQNuJsmY6Kjjf2maiEdKAS1LXWdtMbQrdbGysxoIlbgSYQ1
Sb/WXa84bL0F8qOnpNN6O8ot5JfOuISaiinAJo0gFp98a8MtVlvZ0i/wxwNfzrfJ
0pivseAowTBes1KtAY8GFRSdooJqzu4fxo95NV3oIQpSZu/1CoQshNOSxsX79ti8
Mg7JF33dRdoBop92+E7GV0Kdde7uIPy99f3FGI/26nt1JNwQHp9BlamnD7eobVBG
u4k40r9oSRJWP4Yo6EctR0YPZk+9fzRmAFIZQ2HK4tiIX2lvYEAHceqyLdeIwamA
eQzoWnbuBmMUg+hzWZi001Ge4HJZXBRgpmq6W0dABICkRqnfsP2LYDm4N2TWhyzn
f07Z+sf/z35zljAfLrwi8bGPHRraTZ6/jqVA6oA1DjA21zDwjbo5q4iYqLTnv+x7
KafR56RmEXg8+MCKyDtokkwFxR8d4ryIpHLa3bYCHMIg9NijEd1d9/Wb2ixKpM57
v2ettNVK1PUXq3+lZMzpquyVOhUwbSuuX0D1ZOsi9KEtPsRGNn/TttRF5BR2kFdl
hWV9LUS94ydLorxmE8FxvMsDVe1ofSFq2AREjPSiRoWP8VoxfvSoAC8AkgOwAVdE
atxBR9D2O5FMf2ZEFF0qjJ89cXOQUtkwf4NalphDlsyQaYWtRlaa4zZJKywPi9yG
7zoP+FwltN/h14psubfLfzwIpDsxJC7uF7NsXIAIBfyDf75xXDfdfMZU4UwhPnbS
K9PkrGB6vr5zgqYFuRYZzYf1UhswCVRFxihoR4GEUbCBgBTVyDpJhhmwzqAkcqaj
UQh7NUk9GDEsLH6+PROlxSfCd8KLK1T40EfEMUG4VJXaSvk4rqpS5qOtm0Z8BnyI
1EK8/xGg7YJHaPm+S4y7talMd0XLdiGZEef39IqK6M5QZgufd2yPhx7l5H2Z4HfM
bGPt9EnrB6L7PTW0niLd63FPbRRXO8T4NcMcGTMHztyp4Q8OAA1inaAsEKVFLgJB
zbhlZzCqaIZteY9EkwPRbbWngfeGmx/LKQEH0TCbKxIq6P3HS1RUHr4vD2f1RtvF
M34ktQfHZMFgukT7ZIHNZMSbsxIDT3AjNS60uieQQoyURcV7+XuzydTcVIOH1PJK
8M7QqD88WqKBDy1/Y93QzfAVkHrPMGqU24TFQHyqlO+4pmqj5g4cD6zabhXL3PD9
t9z4b7/6hSFPi+4bZLGTpiO5cqL9dF6Yirpr94oTy3HWEXCMPay7e3z4BxfsGCyt
U4/Izvwe1sjz1ABotOO7BCy80irIfTmRrUqKaEboakplpQtAGs6rDDLGipjbvqOv
I1Tr/hMIdFaY3ssBEJDYKft/vRdndrBHTwLblWm48RtB1HWb0HZXdfUTeoefcqXr
hVCsc7t/3vrFAHyAjsRgL8YreYIfe6y4bUvg+fo93PlzcIjYABqHKPi2DGKYn0lp
PQCL0FdihOsgBWLbSTJHct4M9ZmG87/w9HgOE3meV3FvwLAstohy/xVJNPCAwI8b
2CP6OyphbaUUbExLrrgRuh8TIRk8FP4p35h+zXWXWrFnJgJ+B5PEYHETZebx6iy5
/yIhKV1GyLC5psKpRbm0BPTwAlAYRRkCpflUKN2qlmNFkmzHkdpHNrXiKQCNjp3g
dflgSm8QQ1rvhb3B92B0gprh0lJlgBR6APEDfDTlHvC0dG3LW3YEenX5Uk0CLGIx
h9vTp90duSrSQbPNV0iZ73fG6IkCR/Yfoi5mPL9mrD0TLB9rPgkCYj4a02l8RcUR
jwZHzt0QdqrMP3Z3X6qrkwWaYm1oXdbufwjQv5l7xJrKZQD/p8FQMug33Uqe3NHn
jvb6Ggpr3NZmdPwx45oTgnNn0it8UFvhgU29DEt2VbzbjV93r7SMe6k/adiE2hkM
wCdfME5jESiVcHW09Jjwfa60aviMsdow70ru9p2+3ficz8Oi71yYSQVP1SQ+kbNA
Jxcpsga9ZpAOfZhtsFKYeuBl/Ir92FazD1vGLm9Ca5txXzK5TepnWxRVx1/sVMxw
aB0ma2oY/90MNl5rgnWxJwh7CWJtut2uUuTT3b4LNqIUEF7x1OqyD1srg/mjL/+M
WlC9o6yg/g7jo/eoUFqutv24ZVagptmiUSejCLPRL4ZZyqeS3zx5oGg6pmIS0oBj
fSZL4PbONan58XqtSeOWSsDRwElGniQOxeWzEOPd8Qni1nUtUI8YzBcJoJegIH+d
O+61n7tIUQDgggAbCzmn0/F/JYzbuOO1SYmT5WhH05C/rbjkaPdQcStKpeRXY0Ky
d3agWr6NUJPSzdEEOyLYc6g/n3eiMR678wRBAwacRMlGF9nJn1ajSf9JFi2F3y/Z
MsGg7dBCx94CsxwW+T2lh2rMppog/sa2vhMa3dowGHW705sMoXeON1diC70TaBkw
irA4+mnPi44qifCKwvQWE4p2cs5w6eG2GEiTZ9oPZHNee3FOyW9pz1ZMwrQDThXR
UjoU0cfOxD9KLuEj1BYx64sdXkNRgVJYrACuj4VrG1N+SX0Qt9anMN3X49Mlo4p/
Q8yoBt5DK+QF7vcHhuEFp86pxQREjs8SAn1GU3CStBcf/d4jlTK2XSGqCkt8e7LX
bSK+Ugsb6pHXd+9TzndsiChDDGave+YIc54VC944MHWVKORnuphBFaMakqlq6mKe
k9/s9zra2eazvp7pkcyVG8rfCYxoIhLlQu5fi+A7iZw2ZxPZnWg6ABcjiNm9N4BU
uFWGGNe/hw8CWWR80p9iPvl/m9TpsROI/6ojTQYp2c+SOGw+GNz8VS3ecNny3qSV
81VvZpmhrCw72Rjam1408zbR4uD8nsq5dBqqdFnNMog1QXzhDT+t0bUjwl/935N7
CKygUsuAKh9qIvQwcAdFX4WA5Yv3s5JGE1i0Y5LW/Jvq5y4O8CjGezbZhVUf9ANV
HScLvi/7V08ptrjaFE96COTWtEgNdkDIqL/XQvgARG+qVmyAy9rgZs1BS7/dJtqo
Q47tglNyf0cWKZ7vAWurn4Uy8hw3Qcwfp3IwjIRgh6ER1E3USbZZha0hWK2OuxCz
zxJCBh9eKXkLaWOqnXmWM8BJ5KC75TZrAoOIyVuiMhlLEUZ3Rg0ZO9DJWY69BrIR
tjScENE/rFrhWaumrg4kmTqOcWk4g90cVn3EJolJ9GrnAWf2rIZO5QjONyvydvlb
HVZ0W1WvdRMceoQFwhdkoec6iqwH2f4naMNFPZRDifSc0jEVVYN2TyaqAdU/Ibzo
+EBT6xWxZawKtHX0IIvCGS1O/WuhzvILVkJ9nrLXdqm8X4WSpydw/VsRu4mx0kCi
hDWJiztP52DO8uI3qWEPSAzICqycDUuhP8E0FOyiWI1j2v4nPtb7HirIoMeFsgbi
eMUiDGBDpjFYueS0uE6Po64p6YIGBwoEqUY/0cMo7ZAueJ2GGFFJVw8DrJ+QzcZa
pYvAIk8utExzb+eWwNaL9+glzybg1i1vxShCCVHgxMp6gqtKogbdUnut2HBGHNR8
qeEdCMw3df3hFUhV4r0ovmiefA+FpOH2o2+k+2Qm+WlJ2CvCXTcUmUkAKYbXYOZU
+cFV38PUzIJsVG04p+nLDqK2npBiJjnrRx/MY4Y2yV38AhtXkrrbJh2UaWpUMt9S
AjramyUy4MAAa845jS834oH4gfUWJ7YqCWKkvUXVuusDIC0WcmRoM0bE2FFoiUeY
WMkD7vef1QWJpf8EmgsWm99bFyRXt+lVijUruQFlgAHRCwi3KK6Letmq/tB9KF6d
cc6UdstvrujZFpaasucu0tZu3bUZZpN4c5jnsLMFrAKq2Nm9AHowqllEShJetfCx
KWWZo+0HB4EQwSd9xt8VEIgd+zsWkNby75UWTNi5eEXVP5jLXrRPyx02TgK6m1OG
8Whz5DWF4vmBqk7SpIng6eieOm2FqRef7qiwY3omrTn4z7qQGpDGUwaEtU9uA/lI
rZentvxws9jAm+FaT3W1rPszR8qVne9f9NPwH5a5L0nNnQbVDSTfA/ZtR4U0/ZPk
Uh6EHRsAAq4FabeBRWoMS3jr31iOQEnWYTTYOdEcL1OO/D6F37gBpmwTUw45J0ZJ
6L9TuELwBZt48Rek/6TTnHD4E+A9EDgu+ZCN+9l1hHY4XqmzXcf1RdKjjicS5cqh
Ga5s4VmYr85so2npqUv/cOvLlcxzbgNG+D+lR/Uu279yph3QhMkmR4IsueNzeQ7J
bRR0+HuxtlrBqlTaNqgSaxvnyS+OTZv3BXb6+DyxPgRSJSkdhDLfXA8vVUdoPdOp
pv2ulSk9oRYSen/LVaNblKNGxWn75DzhF0tL4uNZpCHhoo1fJiygRG/Ym7Mh09iM
kzBuVmPuV1UcMRQRzfzCk8I0GPyieepkYQNOtjooPpeyCxMnIfaLMuvWXMolL1ZO
oSfF9JLONOUWIcgIhdnJsHpX6uVIjoBkc0ehxvpUmqTN+EZsznq7jvpLmFs7WGK2
4MYymBNN4Gm6dy/g+EdhRvZmUkPHVD5lHj7FqDjWZbceDKG54qY/YOJJ/M8sI3YC
EpBRnhrTET4yu1oqZJLvhHUQGdgBBtJuh//0pNHEkgbyNjjVzdWOaI0BktOMgGm5
m8evuH+v0aUwlxd/5zkntX2NI2OUY5ZzdpcJu81ORDDYpdw+pGHwbZk5toK95oTc
EuyiJbNgFfcEgYieNStwtTqr9tJQeim5yRRW0N5SQhz2K2PBfWpYjoYV2P/+Eolv
5j26b/C1AM1Tic3s2EV0AlaBAw7dZO+ZPFKS90sikNVSjoBetc0H+U/xws5kn9ZS
LeqnwnIq0xSat1Tlk6bn4AS3tVari7RlSuFZBuO5ABBB7mQhVrQxwatsE7AuxmvY
FruL9tdjy3kuN4uw+nu60bix3nOtEufWcPMnMRpOShhhaXnwn0SZ5c8Mf/2FJhWt
IFFdHdQnF9ddrXB0EAYLnhGJKgzvycoIdXv+RB7MzSK4glwHTawCwpV16OdXdRnz
RZtiziGcjEVhnk/3c/0hrNSO3dO9u7eruvfOtUJNccuAKl3wQhwbhhmotPq4vtF+
um+n8rq65GERBemiTT2iqH8XzFa0HxcedYsT/VNcUquCYPGX6+519WgBy9WGcXhz
3CmXzapR5lR8b3h54LtgGMRbOMpi0H+jaZ0PhcomgHDYGtEfujQpkwXcr0ppk+7Y
HjDiU4PUOBOe3DV2UGPnTCpzDJsiGB3fX6zLv/q1beHf1/U9LYJjTaCLF67HZwqm
fRl1sd1OOVeVqDMGSYdCBB2FCDEhorOo9JCm4E2I2UT6djTI/q+2c443OdgWFvjM
`protect END_PROTECTED
