`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ugPqYHDD8czmxxeXFY92zohSYBffJyNmm2lxYjIRZS/TKGI4eIofOjB6yl0As4wP
XlEuCFIdpNj/5Yu/MtHGAzJgGhC9F25w76vebty1JOTs+FCeSOjvmupcbwHCsYxn
0UKo2elMHShCUiOr3m0CBvS9D5I5f2wHIfncQJxZWrmRjVxqGnL+9wecdE92N0cP
u37Z3WDvnIhOJiRfBnAGK7C0TymRzcWc/vaADH60DParANZiM/+P9a3YLh+JD9ib
p5RQthb2w2ix50PmOTSST7ryR5mK133gi2hSPK1ILc79bwYU86bAnp38SPj/HZdm
HCy3E5juclpJiSUulDk9tfTJhVxF6oBnkGe4sw/dGoALsii4iEOrzeXoZCBa+jQs
s2BRJL/umpubthKIExPFNryYYRNPbc5929MiiyskjbHroco4Rl1z3uracNJTSbus
VsAj/RETKa2OOxNEm1WV7ZAonttxA7RViIKzv+n4pUI5OwBNiLdlTWjOHkvA8nWq
`protect END_PROTECTED
