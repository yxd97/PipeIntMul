`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XSmzS/0Nwvg8cPlBfFmERgq8LSiRykGxW+BO/xVGeRQUk9rXRZ0o1VeopwiFK6wH
Qkaj3u0T2oXbBlumksTkyDXQxCZZGBOMvlVykOXHgAiaO4zGOyVMyToA9dLbGw8Z
kVeKplG3zv//dZkOplOgyZkaXsiAmA6tVZcj/I/45B548RhwSwALAFAORCHd13/E
Y52Amlv4zQbXjICTClsIstJg8gl9/LaCQY5HqUZXlVjasnxNgy5RJtlCJcbPX/Dt
rlnNwnBJRmbcrEK5ZT0CQA==
`protect END_PROTECTED
