`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/3Zf8DlaiXRK4cS/Mk+7SgOhVRp+h35//gMMCO2kc4RfU2HoFzKHcuxdPaj4K1qt
W9b5mI95VGkaUgYyiv8PcTKXR7uVIgW8xHgUnnQjsW+fWt9Y29iLCLglLHJOcAmd
Bwgp4g6I4h9m8B+2EH90Whasb5EeRhBo9lwLsj0MwSsOlxUxXeZQj7QpKRtm9rwA
VQXE9KLldtuKgeeFV8QLd8RsJPd6pBwOQJZ14wY+Gqb0i1iDEbtBCrMQ9pPmNM5n
GQ5c7otKCoozZXOusWNqXO+dcwQ9IcrxoWH6g5GzPR5Eiy9erZq3YMl8qvB9+Vjl
tba+FCTONHPiZPi8xPK5vMEA90d2b+FxfeWb+4hniR3rBatMdd5F029BzYozTS7d
sycEi1j4TE7ct0wOtooU8biSXk8N+EgdtDeRQZcKKLg=
`protect END_PROTECTED
