`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gKTEstiJjEqlj0Tcsn7CgSh/RfUp/IqJYRz98jsY5FOXljOJ1q0+bcT3tGBZLAnh
MphHHyKb8f3AZ1i461a12aeUjL8niii4uZXAzEEcCZzcfyesHiVZnJugD8WxUWZ/
eH/pTQR6cc+0ZsGzcBeWK8n54TTomllvuckBMGI8VAfHn//tl3zVEVQ7Eq+sF9VU
9QLr4s2wtwdeuVJ9X3eTUOxGE7r+5hVGmU3XNh6bS5c7uhrk+MZGMzhD2VRb5nRF
jIqHRXx0nRjOqyHTbqHXkaOPfNVEvWL+nYpcpzP78u0UK5+sSIfGiegAFM10hR6L
9zH2K5SVhVhoyqQfH3AHNOUhZ9Tzlg71lTOSZCSMy56oAI+cVrE0MhiUcRv+okEa
n/P+xuKrbBTStELpBgKn8Q==
`protect END_PROTECTED
