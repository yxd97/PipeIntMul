`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f04YRt+nVOZ0p3SMhefrd9Bl3GhH9KjCVEml56ZQSHkVwaJ+KVK/GjIR3Ii+1hkE
p3pny/kiQaGJENjrAAv1RpnIMV8LdyEWczXtZbjuG4O3CFzhzofGuAuAqFVtC9B6
VLWodsWt8ublSQ3hlEbI8xHWDQzPNROwnNwIDpAN0bJZRlGKqAa9bO7fMEDU1Kdr
CRW+reYoKubPsAD8FhkErtrAzbk6SCXWyjULfaq6FDKx/SWL5h3lj1neaCczqAqn
PAhp2eEaKsDy0NCOyCAdkprWyPeWxdOhSms11g/GajVYVs6Zlql4yVwTHQ4/ADoO
C/jQt+a7P0BFbrQ4g74QR1soSk2hcQN/IoTSsvt4mZR9m8XizYefdtNPLLwOdGmW
L/XDSXdr0f2KfDsFZ7GtvQ==
`protect END_PROTECTED
