`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/S5KflMVylhSa4b4aPB9ZCVFxbKtr0TGQP5Zo54Mv5x5cuKWRZenS5/g3JFGDg9
QgNVxqrXPD3BlJKIjtCcU2FR7Aftzs2JEqNJs1va1jnZ0Jn8uqwHgoXs2iRwvOjp
u1mj7BOn1+mI5tuw8QR5OcSMcFB7+kTFFFj0nbWxTs5eivlaiwBBCVb7mmuEkQVP
2sy8Nk9ydy5+kKEh0LGEaU5TsLO0BuaiGQCOgSppZMQMQTBv7kFADT7IR36RcQ6V
VFunMQLnHwwz6Qyqq1ECg/OaMAnWeJO7Zp6Qsqp+WQC/gyiUS1QtuLF1AbPAyu/W
GEPCRu5B6znh+Dqr6HPyXA/57C+1K+l68fEHbCYHVOq2ISk4n64TZfoYecEpSGHE
mQJXSiOzt4v8sSg3j3BHkDvVc2LIpR8w17MESk3Tu3Z5MV3DUzmD2jmT4fZyQKH6
t1Lj4YVVdKBhPGjfls71vMWWkYdXpFzhBex6QAt5aSSoqBEgiPqO+hY+WQC8DNn4
fYV80mGL2qBJ1IwK5SXScDgc9DwmITGQNdB3tnB/lfEQLZwYuYD6FjsV7YGcaCOP
TYc37tCKNbpth5T4uNd1F+7e8mMEygpJpcMQJTNqu/BRf1xyZkcvSuCUiAj7wlp9
YqjUuD42YaC1/vUrZsdmHE4Uo17TqMcPWHu/t8N70tb4nwlHVgRVOTw3YtxFsXhz
m0+FG1dk6docxHkgyoTKfQ==
`protect END_PROTECTED
