`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDTLxG0gnVPlZJZtJJzC1YUTd7qlHN7PF9SwJSeb7pYkRTGxoTbiETqMTbVL9fZS
9/SIMeNUWh6DFlE76mP09BU4QgwKmmoOqbdFnGviSXafMNQcV3vLlWizhUMJPux1
1K0UdMOLhukKxVvHilsa3RM4Zdj2XRic182+h8+/Zot+uQbLiQBD6u0dhGSrBDuE
ZQjbJUpxZ+R/licqCkp0S/I3xTHBpWElilNX6cNQdQ728VvNgJrC/m7nP5y9gOij
e1aajmBkIfg5pVSfLUjhj8dBKMBJicw3z2cE7oft014=
`protect END_PROTECTED
