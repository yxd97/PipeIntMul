`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xKNss2ZSfokw67W/g9rYd84ZYTmxMs6uhrxUkxuXC6La07QXeElf+NHm+W3jmpyV
F15gBqcwZPMeRsl8qKu5FeiR+EImH5ldt4WU/Wnr0CzKmFB93gUfv05q/173YCMV
auVoGC8yERgdmIRQJlQqvNE8fDKM0NoUWx7+Io8Wfs6KlwvYedyJ/bXAKJdL6qD8
6P+55F0xKYxNHw16160d8+gl48UBpG7/GXC8BCcmHu6JzRJ04uiYr81mycTFG4F+
qeJnuRLUBZtJa4jVnCE8UTia+AgRSAc2TxoUqes35ABsHu+oyWlVplfhg2knx4NX
EtJud7nLDSQIaQLa7H/Aztj6bqeKyIu30hccLdAGIH4HEqikaMEYF3OZt4lETtTW
IeOaE8JBvcKbRW5cLVQGng==
`protect END_PROTECTED
