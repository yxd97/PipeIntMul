`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2zcR500FPu03pQdmhW7Uy79yXQyS2xqA7ncqGGtonHq+h0UqDIVj7CgGA5PU28b
FHYeYrIvezyk9Puly+WBlNen7mnJwHP3dbCSVazC1zRTnvGfHY7yFqb7G4z6g3Pw
ixf9RRkH0luwZawNBSyyTX0w+5+3Euwfo0Z8gLiV6+tQO3O1ct41yRQE3AjSAyYs
zu0ecyGuBFPPONwLcnMf8TWM1UA6uMKPLmr3jsUyobPjWUNUIPYjtprcVB+OEoC0
th28CiQOdilkhoGoEgysKU64xyzoKb6CyZ+ZCQby3rkqqWjne66pmbVjXxUO6OGt
LZA+tg74CDjq1yohXEex6JqI7bQhghaXlvMJdcDN29e6lefC2oJqtaaFTLttdsdJ
XSqG/UDVnG3B0mycdo35JQB6WYs/uKD2q3Gdti6g+zfSwSOiBOrQgGUkZiMQBZvW
i7V+ESXiqquC9Qe68zZ7glIccpftDRbrsIIr0NfaGxH4coqKkin64t7raLtO7jJo
WkFoK942hVnSgxXHSgo0AwEOkCrMgSRQWTG5ZKXhdoeZd2O5RwONvtIjgI1CTY24
k941wkzlw25Rbm5mypQsEcuSuUTdVPQVzWJHwFlGERde1NzuxZfCv1OaVMeHOTQw
ZzckcZcrAsS03LB5KvxGz14Qt5NKEk8m/U37pD//4Kvd3Fj/kTOMHp+I2hTO6xaz
x7ImNWiF4YWsV0Sc53GnHuWiHnOFCUTJRqnGrV6gOdBI9/YK//c2a6Dt13WjikRi
NVph2Good/3yEuncg6vjl3Hhr+3SUL5hTpWTObYEdPOUkaqew87vMXKNcqWOlO2B
4Q9Z1xmEho9+BoV7PWmNv1wim1PxmVUwD0RqDykLtuLrU2gxO3mwM8DTdFcnMzUP
8WH9kT81N3PumKFsKJn1kMY9g9MmcZh06QGQEJxaZqbNNL9pV1T7Eji3SDMdHdS2
+3xWWGSvTv4CeBdfgVDwHJX1OSMrsH+N0fSZLpI4sNy/f0OpV//ZSB+iVsuzqVdc
nXKemsxu3VuklvMC5atE0iYx2gdFWjWf/MaxfVdo76/auJd06x+Cm1+B10rQbHC9
Mr3n8PcimvgZizmiS20bAPG3YEXMBsiCQNCskdWyJDoQG2m8qEe7Qc1/ihgnX34q
p4kHGc+sGNx+jB3zUIY4dYz4So1HQWbb2nyOPAcCbJ96O/fRJLDIstJ13j4CPLsG
RIhbaxjak1uhkqi7QwM+5vYUDeNziT8b1xp3smemAoKvMbiUuMI9ZqcEHmcwI1rq
S9bRZCMcNeDZcCfE8BbgdHvZUpSFXZM0jmIl0RbwEeDVsPJ/1euW0zs/TsNKj599
xFOztK1+CAE5lj5tjpegz03rxA7n8K+0uASYDeWj/JoG7ILUncgiqjWoPADyc6X4
RqmiHd1rpHt/rtOQGquQHYYemAUp7YBhzBwKucFMEEN28iEpjYmNPzF+b41e/FuX
H8/oZkKv4oNBkdSDoTY6kc3Dw0RX/LZeFL2BcwYt7OfyPJu/qvf3m0HElJR6wyjN
HVFvdQqNozdsUpMPQOuKZVc+ohOLpFlrn8zzwDiJGNPb8knyKTJtwEoOiTY+Sqpc
hejAe+D/O2VobcIRFaagTMv17T+fVrtmmuU796i8edg3rTei9Iqb1xheFj2Uz48h
Z4fR6DZv3ZsjU7d8u7mYf81qUPbgZevcCDqaHtYjo9z7+WuTuhLntAtrNv6LczCv
ve6pnscj7SnnCYZqQydhiHnw5OwH0ymxEzBKgD6+zh+w8Mz0OB92QEYMuhSATI5D
bpjrlX6g/5liiNYHFAEocKIiX/MqzE+3lmwTtqQTuWv6oIdWTZii2D36vLTTEmoe
d1jCtXqEt00hug1Um/FT4qa669jAmaWtFAc3TLrWTnFG3nttBtav1rPRmSJZPrp6
6t1SlqZWmfT3lFr7A/QBnHUzH9GmCShONVRc0OWCFB2Zb05HE9bvjet3kC8MTRCO
WQKDonVF6K+qTBsqFWPyqMBU9Im22BvEFLDuqdmsWpwGB79xX4B9GDUmE9G8k3ma
vuPjdVpET1e0FDgluhTOrG5N62u2+xnnjaHm5JFd/JRLZg5o/HiyE4FGf4Ito5wW
0c1wwPqgZ/BxIIMrT2jPKEvHV+eukzLewyNNYoVSgHEsu0B8IMRsKsc/qMa8Zn3h
Sdc2fZhcmlIRD0YBqPVfjBxnlACzoZg8vHDrz0iEsgTICyHJCc0l/MItOeTyV7RS
Z5i5+JfTglFSi4J9V/tOvBo38TlCLQVPd2vqZfQlR19L/Jq03fzmaTmhZ42/qQpm
MTe4wDI5c7C+GMqEpwsU1wXTWzpi0IwpYjdejBFvVkn5oI1ADzN6r7Ee1gkitn9m
w3lOLnS2523dBeewxy0Y13OE0JN5GGYZ+2u1QjFZxkzRu4aBp1FKbQ8BBkbeRAav
CAyIljGDCtojg+xkixFon07FK0NZfwygOfIlK2sB6XOcKEUiF7L3pV4L+KPyiGGk
unTwsEzjGWw2duh9ed5dr5v21zoiQPr/hnoQ6t2IwWI=
`protect END_PROTECTED
