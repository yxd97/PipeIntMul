`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HntqQ2Lb4qoxHse/lJFswo6JkjKp14M2COcXgXb38AjgBzeZ0STUrA9mteSdA3vE
GMJRw7GaYGwfhTeQryCauFoGQoeC+HjzR9Hn1ik77BvOt1IURmoxqo8CLn4zLxXT
ctequCD8b0Zp0BB6wA0Xtz4osVjJn/Xj3z4nLaDM9wfaTYexqvVjYxRn7/rq+ELo
BQSH/DMRVW9fo2NhNK9XnzZqpdlBNw4tsEvtltqncQNs36YjKwcMdKNuPVK5FT5T
btbOMrrXSXHwSjr51rDqOqYKD0InAO0P8pp7/Tof2XX15rCB4Xt1cp0RVklKgxkV
+82qWR0hA8qIxmtFByRVihInaXepKQF068FPIVuHPR6l6IRImI4cfo+Kc7sgEaVz
VpA6/I8AMocTO2DUVZM2WpVuR+aytOmvxhUR5eysZMqvsbE3Spd8oK/HbOBIo+zM
`protect END_PROTECTED
