`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8WuQ6NyZ+HxJjZYkNQycFcGZXPyushVWR6HL7M8/nh3bLja7iGZ8n08gn1+F6L+2
KZFLZUAdZ586HrgIqebZqwjQ8ff34PpprYmMrgckGBaAimSQInKftkQ5DwfxtQ9Y
zZvMoqqESDj/WqaKr2R/n52AtzziDCQNMXNPV+mSZJskreLBddUZ67ymGioGOVTx
OIvQTo5D9EEt/p9RFn/HIYNFC0mu8I5KFnJLbCuhfP5FAdr2IW5TPiyds1KpZgod
GywURPck7KHBzJnwxRTnsOwkboI9Uf2sr2VX6+VRi9vrQuNK3eShmUOhJoCxudOk
2U8wrTdqaJL53WbLZN5z+w6K1jlkeO8QsS8VTp5FTV7RNlsWai7B1+Wmrlk4LA5g
30UPwzeNftNxnVi3Ah32Oq00OWy7IYuFsU9ZZnSaiUOYJ6/W/gV3JtPhbRfMQq4/
fTaii5aU8OOK+CvlicZ2RDGcmGfqQiJXghA9qKp/eVBvWilZtsv3R7sL5cygajnx
AgpHwOMycdLoRj9OHe/BUen16YFbswDMrocUCXa9DoPauYWM+QK/TVBCEhSMdvBy
LUcHYI9v6pBDnE5yC1UwPo0nI+zWL7D5xIU4SGU4/hcn/FCZmEjfdOcJ5+07kSy9
iHAtrR5K+V0ZRG8y1RTh3w+t33WzSUD+X7mP8fgIbViDen1B00Nmf/3JshLKKgpp
CtrTknPgseNn5JCnlYq+0rBjsOB/N6AXJOmbLHDRmOlVm6m6VtdeRfdjZKDbNkZY
heagf/joRa/a0DwNoXA4JKftyvolH0Uni9QiaDwPVRZyrVMPJSElWd6v7drIVJuq
Zg/Xmkjg3yY/TvFDcjIQYLEZ0g7TJPSiHG6XFJ5Dc1lzYkKps5QbTz7H6wdK8PmA
GwkfX0Z/ClouYvWJOQ9EzH4YF6ANIJgrt6Vqg2DAT4OZ+Snouosc266pY7c6J2dK
fVkXeilL4ZJPnsg2mdkmAUMvr6rPbVBMAktM2WCORRz3YA9cOEyDyGZtAfukZWcP
Zzz6z6OlQQ2EQmpXhGYlQXhO3OeLhcG74/QbU9Sv8PE7oyZZJlvtc3+5E0NbyZ5L
8mhcgaYYV0LN6x0pVC3nCEaFtnOlxzYnWGkfPxndhr7LJSAdXZWHb4zkBVObr/i8
cHnt9+FTIi+dO9W46ViPAK+g829L+VfS9kEIJIRsR3rzWzQMQjsrWkkRY3pE/LYz
WZIWnqsNSCJyzLyxD+X6KtMJ3lT5Dzrh/B1CcJfmg7kz557MG8abHoEppHdfgqu/
APtPFScjsID1BGVAvHJ8B7EZMpVVlSD77O2vmpGCNU86nL7N6hfWzie0rYgKjPI0
alMvxqYxDsRYqY8xsC5HO8ZS4Yd3B7RmVEIiJ2ifq1ocNa/kdhi/1mC3im8La/vD
EOrQkv5YnLpAwBeYvHCxcMbd8N7SRldulNAKpyin/89DZGkKy9iGcy3ceSNzxH/y
307fiEOqrQ4vFH+Zv31DHB9haLmld8DQW+P9I4uEfrD3F0tFSjPulkfOoiv5QVca
Uli00xbgRlBlzQm4kh+DqfKo+m5XJadq7qVWCrRI2PToov2hpnYh0l3/cqAsRgQe
5c/ZpVL1toEahsJPLx5XyvgszSbMzfZitIhRdF1ABURmSkVMuwY7Xp5aKRwZKT4X
ZhwG9nwKtOSjcMWgPqjZVkLa5ZdiD98R+cojJ9DGkcZSUIh2F8iVl3Nzl9JUfJmm
P7pi3pqXAxKIRzrvivQZtemmEdu1a/gJlhtDuGUMz46appLbptmr8edwyPtQyJaH
a0OJb8pyRXvQfxqGd163koColsHOU/t2kPjPDeGeSFioUGO5g6pDH+K9A5LrcktI
oEWN+fkrzpTF8j5YIyWVe03vXL5dP0AOkPQY4UFGIeCZeRJyzJ5mTc2aP2X1gNpa
7+wdapMNUTC5/V+cEX3F1IOq/rJElsSpm3ymIkwUldFdt/QR6L37ggfdfER01K0C
zWkBWltALUwP/NbBJlbL0XV56RUFLcrM6qk3vkRbqNQWZB/6HHzymcxz5MTm8uvZ
H1O41PnJV5Upzr0UxGOdf9ndysKOTXvAA9Ybybi+pT+rSCFeiv76KHgmb8CD+2aL
fbI7McMl5yEPzt09pMFOGCXGAsY1YZlnUi+bpgnOG131KPHXqF3iK+zSy3Yh8lV+
ICwpoFKcdDcGzVqorgSfYbpUX1BiS1fX3VTBoLyeo2eoyGOEq93P1Hiu4T6Emy52
WroxeM7bhbygYaNFwayfPlfS60UXZifJxy1RZdM+RbnZoycmGdJDp4a5r5aaCCKE
6xZbh86e1W8NCj6vAI6h5r2KrE1ng7tPZ5aUSDNupuI=
`protect END_PROTECTED
