`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jrp5JBqoqbU14oO/zOaXN8fcOhuvCyJPWTUIXJ2U0F01m665KLgFN9fa4eMlu4ci
nrfwUELsn+IIVHYX789Nbs4UOYUzlpcVJ5tbm73IBVj1AxBc7NQapy6Xb1gGEk/P
6ynh37FPxeT+l6icAOfJz0VInwb56Hc4o+YZIsCIfJdEI2T0VKm5Ch+pOMhgb9Xt
6Vp/OIICVvaJSr8tNnAo0XK6rQjvpFxt1MZtSok/2+vcLh+ZSJK6Kx8PyZRFTFsw
zQu3mlZ4JBTUNa8/IGHahG9wGWB+m3B4baf8yTxP0zitcUqjaMt6nLD7Gz76/Zug
Sedm/dOjZP4WKsBYrxmj5w==
`protect END_PROTECTED
