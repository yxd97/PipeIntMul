`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x9vVZym+7flbHBLGSzxSEPH50/AiUSZrjBecu6cVv2+/yhM+1fQ/zhZMJsFPEoc9
mW4SbT8LaLTsJD5vj4VgTEwWbhWpvgvR/O7GaDwaLzPmJ/AROV9FSWVwr2iXosA1
5s5mH8KGGEEFcfsEqS8A9U3S352m0ANtEfFjrLcDLrt2JP2vlL646GuLPTF1N4ML
pWysQE3QbGmB/el83QyUkL5PpofPkSrZndYG6qtIRmiX2AWNmVslcsDwJp+LykP0
43oeFkoRD4SUXE7gfVXATtW6sSsy7PjyfZhDG61BuOqOARF+X8YooIIJfvLciYSP
pTwsb+yTht9NulHIH2ba3Q==
`protect END_PROTECTED
