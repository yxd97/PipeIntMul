`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5XDDhc4PaEZLWRy2V4ytYPSJHQVbNs2ceyFoENO4SFcgQr1dTP7f69EOfeokzI0
Pw19L8fXUvRltAkc7jYtep4IVT1hik8qetxh+Xchy9sF9YqU61xw2WbfOqKH/LQy
mBqZ2J8+aKXWOjRLMpsPa4eYESUf1knJVIUdzxSJSroKatVJdApsmFdyDWW7fV8K
IhH6W1MwIEb++OVxyLr+lZ9s92RFxuCstPlIFGCoV0t8jHGhjV8LuSGh4FBb/sfT
REpV29mJ4FP3dzp8Js4MSsv+tkmABRprNQ7SLVkdcjhTDpPaTPpowGH9vKMYl4/k
9YeJ0DnvN13vmufompEISqEQTprYblHGU23iaCIskYrPC1cWc3lOMWjKNBVa3DsP
UhvyH12dPg7wwL9F89FAXN3wZPtzjy+q+DH1qszmJ2TDn71vjDhQXwJA5b4ZESQq
vDae29JtwnRqIRH2CEbpNRkdwMW9vJuc6MAn7V5e26lM2upNNl1B0fy1h/zKe6UK
`protect END_PROTECTED
