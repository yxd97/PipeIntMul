`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kedfELPV4MlaFYL4N0lBfYa0raPQxzf8V0Zh/+uSB1Gd9XLOdK3vrINiD3EKqSXX
Ba3aa8KfMF6d0SO1K3SW01VaHouqPaPF8ksB0TNmPB1U6mYm7tv4kCjAjWvhqC0L
xeGybuKX7IW4iHM17sua7gamd1RrTS6nLC4VUIxuFQx68DmMpohpYBz+G1GxbzFo
/3WRKnItjI2L7/b4Imq1FmPYVG48FDdFVUhKCP7sTKyw6YP+X3p8WFiq2Zypz7I5
AP4K8rwY5+Sy/beZwUE8CXSoOpxwk93EFS1yk6cL5HvTEeVjyB0/pDMhPX7jyg8E
udmFVKygqBG9MwPNvjuBHwM6UdLwjbhnrHQoOmoT4tlSVfO8IR/HP1WVLzNu+LkW
A3DTmYuR+f/rCFKEahHediU/jsZgKAw9MFFgIl7Pg2PMgwf69gwesXQ3Ayxo0qtZ
NqZiqX+LxjbqtXdA4ElifOnPTXCqvz8GJIvNh70NzFFfs9d3L5yiZDSHNQhYNET5
`protect END_PROTECTED
