`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXqDq6zbWkDMt3gmmoG029zRHdFeIXFg0vPb6yy5KJgmtRa6efRz75OV/0++bE3S
dZncQjuJFaBpbBpaDogmtQc72Yg5t58js1Cm+M46x+PpQ5wysKfNrKhGopmpNYer
LAzgzjziyeQNdpQjFk3tuxRP2j4LhjVsbE0/VZE90VcxgXTqjteRv2gji8ZzEQQg
naBIDotCHEqyz2di1+xz6uZa641JrUDu9V3cghwNeRu9VC5hlcPKmKxz99F/80+g
8Cbx53rl9mrRdvjWA48U+0OJ2K6hLYmyNiEJL6zTpW1gqlAQ6mEsvUQwM1xcmf4k
/FW5f3JWJNeVeSzcDlE+kqbZrnLsz/fsBJw/RAzQmID3OFjdAzBBTzrB7iTOyH61
KcJTp6N0jgQszuL3odiTJlipHFjxdmDHCMmYFroZcfziGVWh6pnJoGbHukncPRoA
r0+FoZxWMtBx/qToTdzpYbTR3VjNmqg1/SgBIgNMEE3pHPA1hDD6AU0BYbaWqj55
1UP8sk0rBa6N2zZtqgUKwgyMezk6YTB2Yq/KiGGRcXqgCwTBxs2UOwafrSD/4XR9
v+I2lb6f1pMvUT/dD607LB3uGwj5zkuCg2uNBxwFAQYrgPjGuwtXkioFa6OYB7kO
m/Xa9YJpKnxfIxssXWT1C2lX1hujTzyjDnvOzbaP488mi71TR54yzZw2D0iVzxVw
jhYSUw/U/cn9tX3HccMUX/RnqEnaakn98YwX5MEfr030BTiGLfnz+eW/wq6yP2Nh
VC8dXnmoiXbLSk/yA2DPxxbRvoz2d7UzR7NkMRUx3yVDjoMdmZU5jfwA/P/lLIEb
W/G14R8Qy/7wXoesU+MI2SaO9O/iiQyaPLjS4atb8t0TI6STxIGiVHo5ayuEUx7j
fQmwq0iofmUzveHdo6H9f4Y4kzpjCLhaXK/XjVYgdPTLDIFo9GVKPu1E+wZojVzI
EZliO25CBhwLc/GLChXy2qFqHTd8VGliN8yCeJC9CMnxUzDKS3Ry/IyzgmwAy8Dg
FtstdsBrq9XP31rx5aytOR4U/QGo5Ymav3f+jzSd/bziej1jOQiUKhUY0cK5ufC5
+biYDb1T4JRBlbjPLdfJowEhGtlxokTaDPHydaLzyrvpxZYz6hSCVEMsub4MMuKu
5qMwDuim540Rpayrx1BRwqohETP8L9epNlHKQ6xbxPE5A9UpLdsH6qX1+PA3dl0J
OCPF8altvqJTqGyROM9hiE3IIxfK5Hj+/B+ec1w5MXNboZiQT/utmQ11pQoCdU5e
249tt3jsa4pav1TfqAHdAXdFCxYEPQ0wBdXE6Y+KHEo8v8s3uT6nsBPnIwRCNk8o
cBg3hXQFE28YiI72OHs2F8YYWttHz/jPIoAA3pRqEwni4P8RkeR+QRA1HuGxACqJ
Q9j1NfjqEEPtVpz7M5719D8iQOMsySJ3OW6z4F15VZ7dwFkCzvQQssPRVlKszZyi
chadazansgVbGEJX3oPdFhoManu0ZBjvXBNm9FjEQUMfr06KJwCw1dITXac0Vx/a
/8QaNKXZVMHJCgM9E/who8H13CtB0Kf5uWPn5ozRXFaI4Wp7zfo2FE8tNbxwIYkE
lxsCLo7pRUjG4gn6r3txEe3E18NMXqgqYo4QrUhX8i9QmKjC0IoJdn6J3BvLme2J
yVW3t3+alSG4vAYGWe1bMfkbCKNg3hEMMuMkWKWTOuC+jWvHrGV3KU3TD/iDH9S5
KZWN4igabXSlDSogWuawfCffjNetDZN8qjs/YgpFANAgMqmiD4F1pbeY2k3QTWtF
KTvZDD+kgu2TRi8o98R4AzVv2M8AJpOuJ0RRaDc9JH4GC/bNyaklWlPKx2rl1b0l
ugc9aazj8XRT1rz5+VCO3sNR3YRZ1f8eT6zs3+6vkNS8hUtcmcsjuu6P7YDSJJhI
Yu9uEypbTO0GaQxEHsC/CxlbfHdLUOcIJwWuC2ri3UHXI80t/GNfHzZsZybiBn7Z
avVs3QbknL5x70Y9lI6sTEByMQbRyq9VpV0KKyE2mhp4LkVnwlBE1kASfUTiCcug
TSbhXltgc/3ryuqZyqYXFkIMW20hjtDxIkTZIhr1BFbxaJXej5FrlvsWJD7oH/bG
aeWFfp1OSyibGYIiMHWE4XVR4xab1B9sFc6cmVtXE93lYgXL5k0ZnB1ypf6/WakY
m2g6NzpT61sH1XTpTGE30eo1jxoYayVf6Mf0mCYh7I63X8BGtQ8uJaMgymGLP9vS
tRACXPdEf92lo4Rb9zpx/GcT0Z/gbTY5dmBmcAdMMUcInzCI80p5X5HTlkeZaP+e
O2WxzcGBNdArQcfWVXNQ8mt73vt/+ZnHoV5vQnnJGxVgZ924JZe58s0yStXZuZP7
hoCE7kJNZP3Fqa9GzbyCe8S2yevSPg2U/D/sqDOLLYyt0BLkE6CRH+sg8SqjWebb
3VREgieIe8L16I5vE7LM0EwZKBrQvHuDe8qpRbeeZrWAhsgYWa+YDEZ+oF29wNoV
tJ5glfxMIEAPQGc3Y9PcIrFb4rqQeC0Z1AJBQCyDteQApUAlFOPcK4wCvqjFh9Yh
2eP+AxRI3Ru96JE/6aAxE8AzkO+9DX/mg87cw+mHHwp0WimVeE6nsdaqlNFA44Wc
jKIx2bHMmMRSmeOdS2TeiNHW/qPuwPz+TkokrAk8B7/VmGi9ECwkpzcw3ZwpGpZE
Is8eoRxtJb0DNwwYk6jSSCo9ykou9q8mqivWak+M0Cz1jPA8TiyiYdTQrkI5wNJJ
SYkD0aOmWzpJYkC2/iPYQ0hBGZ+T86fXr/j1NVQNnYqdgxmNF8Qd74U7hH00Yjv2
Vr/nBkaku5o75vw1Cr1X5mN1Cg1sAePoKpVrtO3Xk/vHbP1EYWjK1elAyiMxld/N
i0koohB4VJHncHcWOTXTmHcBOGTfm1wTkHytD5eslJdM9+zB+kv+rcabFm+k+154
9yeBdFzuu5pKBLl7cdF5Iu0+NwcuqzyqFrs5C03hUqfVNClsGdYv4uq+tnMeFTYZ
34ItNzOWMAFlh6HskxzjY53XoWyeq8TMZgzBnRX4lz8gKM9nUATs8tHV8UVOT7n+
S54qmoMxg10H0BBczdguHio2Btv97mo+deWFvVZbN6nNetdejp/6WCT2lE7uTZyJ
Ztc5FrftRNzK2pFxvDlnCkmFBWMxqtnHyHwBVWMzSeDUu7isjJjWoE135GVGjgJi
Df6FBFq6DNVVColmcoDdzVJggk1llEcgjPOHU4SEeG2fCqQNHsF+A300eJbvI7HU
MrpXc3s7r+FWakdFwIjGB2sIVnVVWcrnzXIbDvtv6abeyairpfrWUnTCgXB0TbSb
Yw3u5YvEczo5P6vkMYz4ncImGjtwzqfdp8dr5u3eVAKVjquQzfAce0/RUtDyHDUa
7eS2q94bXOwvwhklB1UWskebyrdzWNE/j2hHJBwHWj3Hy7YrEh+kOXRBzi8ccOek
N3ObGC7R9q7yIUnU8c1tPmSdPGMqbIwxVTyxzVD0KwS9j16SJHzshKmFc33Cig0l
B1pZq4VWuPVQBElaVKNVqXdObrsT5WIu+Mc1dvLuZ349BCWftMgExS/c7PZzAwFf
Hrj8JHoELhLETP0ydJ05pNsj8xZILT+FVvOuAevhZU+omjIVGrSNgGHoOt0lPoK+
a4Q5QNWVmP4KquCImAHICEL2SEUe5+7ZcmS0mDhEXtB/Dxtg5NAT/dsZ4WcbkY/2
RLFrJ07uSDw1RHQBewgaMjYaMx/v3H6QBvRz0zgUDWmkeGNgGlWZuFCd88WTmymO
FzZpMFrNtUp7lFQmgEMVWhiGGd6KwoMJOc+5vCQPHO6boYCFwHFeJ7mlK8JJeHyD
HWSUPBrdt1X6NDGW/uwCRJ8nARmuaJmD5bbLWIhfI7Xu6sm1FpqYfK5Y55+lMLSd
KUGcEVHMBUeKA8E/OLCIPdk9AP0QRaA29g9J1Ht59od54a+6KWqKYkCQpraBWLo4
RdhmWcc00rbZ+CnL50035IxyYEajKOlkDUoIVA1vhAB7brewWwqPlp86g0W5q8ky
J6crGIuPg7QrZCOffpyl3svqbU8vOYH6NSQ0UG/Ik8HxyhglMcvt6UP0dfVzn7rA
BaOrhg/Bp9Gi2na6hGiDA3A0T9DfXuTkgDDdvTYONwZ00lWNQP+63pEieFdfOMng
LRpHB9jwwCIDPtu0egxkrJg1QJnvQqOpcnDVNERBOHTbrQEuLMnxojlK0L0eYdJi
Zgr5bxF/BK02c/bt1RUsgNFjMuxC5OTXJLd74lokPJ7L7Wnyrrb7UKuYNIYTyM18
Tl4cBRPNZFZFuf+2j0LtA/uUABlyOnHBXUF4By+SIytwSyhxOno+So24xkLqV4Ll
apNGzSwtlES6aGoyoJGVUV4r25UwcpnMh3eZTw48W4Ldz6okjzslnG8NL3xUvUMq
qb2MZ3FXO8CsABReOZML8ORLLO6klSbeBFVGIbvw1zM/o5hv8RfSxU6SOJ4XGTFF
b6HjVEiEp7q5taiSNkWY5p00jNH1deiKcal5W+WIeQZXBNQudkxx+KHYQqUoGyeJ
dR22yYgWM+9o158aQXHa1NX4SdZo3NcHHhmGZ+FYZyvICHrwNL+zpmOgzXwfZuhh
mX8xOkm+4r3ZoMTU8jOXaQWb8HU2lEW+wQ/YFLZtfK47zQ5nPaGY6HArxMbfV2XX
jmg6Q9dlRHLi2H+blVUR8otWK/GiaGtxge8zBOqwJvaMXU+AuPz7a28cg3m7JdF7
7MDaz+3lMYTbSllUGlpu8kvUM6oUkRDDsEUC2Q1mYfiBBix7bkaGFDJXou2V777h
QncDN08IVyalOMz/w48x+tR6tUmgGVfkgw7ZL28FghW+CpBbXvRJilMLQ0rA0Y1h
rPgIRxQVncKAczxWkZoMUS46M1Ycs9vIYooRTfGr8V1FwwF2f9JB1dRv49P/LFqU
mTVLTw9DPnCz6CO0tSeZLt0Y4WgRXoxkxXSUxCj1AWgaLIYQIAt4quDbwxo4O6Bf
GhvBae0hTqiQR5FMXL2ue1qno/tMFQVACf8xLyxvaEj+8UQdyhvRebsIOj1geaqK
W1dDnS6f4gQdSR8G3nQFaaC3WG6ybgj2OXzP/njeLngrkiCGGk0ARZ/2onytidCd
uzqJbRUiaj5vXBVdR3lpW3TJdLZSz0rot8STHMIDADHdsq54jZrP6F9wH7LDYjNo
BjAeb4UG8/6VX5f7lj/j231LEeJPgIF8WedyWr6wUeoGZt2uwZ9ZRFOBrr2Gb9v4
AXZyqKd7dK9QmYZUm/FA8oYNlDvnjZVznBP8SbppWtGjKhperc7TveU5VMMe7bte
6gr/tmUI/AdZO/1m5ua+4OU0P6r/Ng+LpN3XJ+Q6V4gPZXTFSGEzjrmLu7/j0av7
RrhuoMVwgiyLwytQiZqfbm4qaQEhiFomTbSfhBAPRN0PA7PwtWwjxPc3/HE68IZc
tGxXvZe7MohYrLLT1L3pVDf09G5UvBosAXSpeNo2+Y+qglFbs9ZDNrjxUBMWr/RW
Wi3aBulcDoHeim306ZAsLDszWbuKTwpVvYe9ZsBL7MvbJWKqqiErsaNtWYtwMDov
oClhUlEan8mOGoeEuSIMvviW1EFM+MRqrcUd0/HaZIQUr/hS5MAyxPw53/zJo/oT
qO8uFFARZfuSrsQn7IOKOtcIBBcPyER4gEwkKVNimHZsdxA909YP3EyuhmtxPiEb
S19cnJ8HXeHhalDV+CcN0B1GBfcFLZI+0HEzAiy7S9qGl0Ly3Mi3KOnZ8MlUuRMr
e99/sToYbzvrcAt9y8whwn99TkaF0r5gbRZBio95nXVTuWczNgXTCe84fG4Jj4rY
+IJqC/cpL+OrGjciWb1i1/SWTwi+Cj5RqoHZQzFcVlth0o6xord1m3mQaSgWz6R1
eV981Gr+yjUrkrW9rajtKuoAB4ZgF0+d06prcYOi+oh5CkeGzTTp0iLzQwxhyGdi
rIi0I2+aGtSJSDe/K+1ZJa4MiIWxLGQIUWvq31IiQKBX7X97pVGQm8YFHxzfgJD2
LBMpeV6UfUStGPEBc36M9uQybnWSa/ABSfQ+Y18X+n4tYlzOLjfHclTiiD+V3ioA
ttvnSV79J0UjHNU8vwWLoeYlN8I6kmyoABOiHF7HoOweGBOK+qqC3UMPfapUPRN8
ifzvljrHTekAsO0bB4ZfI/uj2RLZ+DvWgBsab+o6p4gEJlDXVq68eEgwKlGx130w
Auec3tW0X5Omb6Vhjo/w23fyq0boO8rjL5I/m+S3Ji40z/0uMc477xjMJU3bHHbl
0peU99OQ4iFtHHcmDcE2q8OZsnjURpOcVriuVYn94x5dYYaetkvjN6pRcclrOK5V
qmeSugTT6Ln71LCVtbqnOxjZNljpJP44OHijKVsboQWshKZ0Mi6XFx864cxRsapT
O3A0ogDjEmscIeO6BQqGecHxQxi8Atzq9bi9bHdsaToH+daAGiPopjCXG3BFNHDG
PC8dLaJIIvhBcRp8WpDt0J/HbxQIsFNraq0nQu8wnQIHJeLVSZEXUQPk5WEHKwU+
A3ygCwR52V1IbOKMFo2Yk3ZmvUFDVgbYw6vJIWJ5H3ROALy+kbbdW5YNE4E7Zudb
xlC/RjemLNiQKZ5RejfLg0tbPVK+Xk3ube0ha9e7CdtMkzQoV6LHsihyjhVyH/H8
Ss7FuK0lJt6qYMDKq+pkqsd9VTAIlL1lElxMMWompXVzFuUWn/iVD7uR7KsIPaiR
5YSxsMS9nR8c5shr88xo74aaO+gqjxIyOQtfXWpMvWPYyy0pnUe4xNKr4ACM5NTe
ejzV2ClxBDjgZCAgW0DJPfa+Udf9rUyJ2GJpf5mYUH2wrR7GD+uPky0k1kB8bKD9
gwUzbMDCGVChaQhCS6jbUT+cgAsEZgluvDxUZomWrKNdwcIrlRaCLyraUbeQUakc
+6W44zfqr4KkaXAVbgVUuYuNrM3f2OlVt2VPLwvXY07ewOIBKyIhCS680GqzL78C
hO2YLGI8Ddnox10LMV6wbIhZX2+xsVqDJLt68gFevVlYwJI3zU+9s8ejL4Y20pCn
u4V5QVHhHAtGZm4bq9KPphWkR2IZl9Wr84CmT6iq+g325809gXjyL1gjOoYk3b9z
oUZj/j2p2JpkwMW0xQMa9h/Dr/zq8a+qY4MXXyyFVuNFuK2O885Z9MykxW0n2iBu
ZFD46ousNbKoLfqQd0n6DI9qT7AysGMMWweGGdYg036oLsd+5EfnSYGtR4c96i0X
dsX1qA3YuD4TDUkf5KA0gAVlbT8HMcG/tLVoOlEdH17qzX3fh0az/5bYbtdY6BDJ
LTiuEbqsF6kvXroKGOm6FuCrvmg2lNV/s5P2cGCcKWqmkT2AOvdfFDtqj0B/tTJ7
jMSf2eYSo5PpqQf+h9yf7cePhr5mSYqmuh5l2U8YEn8Pj65yPwHZVKhzfsABciPc
rfsYHru9rAemK2ogoaTrCEBZBWtPXYLrrRBQ0oaXZjXHsQ4BKV5bXAvNWXg5JixN
6k7+7QhsMdv+6g0wiJdOda0tazNlHevOvh86Jd8KG/+0ZudpARAKKQtudwJGVBbS
BSXLjzSlcDgt7XqpEw4xDo70gBES9sp3NzVMzcOlFLg20l7AQMJhsmMIT4qLFMoP
6bjuSKmhB72CiwmpittdCUAYEc+SqkI6xPZBTHVcpQPXS8q4jfKqldISVJc7HtZv
Cm7eBJmY5LFg2fKwCNS6Xq8gF3Uo8hJjSYCoHoxWOudBsLwMxkWfHWFO7kgHKfd4
V0kyFpt2Hd4c2vaeAkHUBC2rsT0X9VqBn9RcGevqsncpBPXKFezrWK8K42xVXtfN
By6D7dxb/2WTl/zcqxbkofeegomeyfaukXA186rRcjkSWSGpSt3gLL9LYyUr48A5
YXPvhXel4hhhzaThHPVDJSpDkj261il4V9DHAVmb2A+ieThBiaXqxgbUZqaYCzKn
yy14WIyBYRYUvu3DTic2Plnwcs0xJ04T41gS1jkxrqz6U4+A4fWBcMwM8xs/PLd3
OT4RvSjElWxZxyDRMNthNcvnwT2wL2dLTQacK54xszCnSejvcaQITlCiEEXmqlOW
xOuSYE8XNM62FozcwYFStR2OzD6P4FgxNEoLWMRPq3jL/mIRvMUT2uLysrtxpuCy
NNNd7IxhUJS9eW56U975Rma4bIV6RKoxpFxLhhku/n8Cy7Jta5/bGZSTo41hgfoF
7oAQ4pkGheWHdYYo8LUa/mVIY8bDL1qR10HSrm1r2nPRsGAJjsd6byP3NS+fPGkH
F7sbXFIu0kNgFWIiDX3RmA4t3d+M3fFDNi5B7DyrpDcQEIETw8hHtm1KGJw++jjU
ruP1bMIxVQ69vl6CUWVPfXSGdgalcYVDABqrMLlvbxM8Dv82JXiMVxhxPzXpNJaF
KWlxJZ9BwNT/FeJwJBzhY5epHGyUkcSGIiaFVxiA5TOSuc951mU0+EGWLUluXqtl
tG7uTohVKSFR86CynhiWPD51y2DMBDFf5LLbQaGQMyf0Ahq0rxAVH9hg8Uo/CFTW
/USo47Bes3II9klnSFEx363XPBUPxa+Egxc2vPS0HK0IBbo8i5Z96TZDy6M4sdoS
OTsAV1dV2wb+I/0hutTbt6hD/nHGP16Mq/mQRaOSd6+Np4fvocoWIoZRyJHl+weu
auOh3qaOoohSAu0bo1d8jDkxMB+FIm2qzVMz89wzHQjEzDZkO0yIDoiTDr/r6hIY
dN9HaRtb7y8gRTuT7tIKx3jWsNyI80fxvFa9ihyAIbsF/VE1rJHwfrn3Q8h8p1p6
bcLCTDUnHfnLQUVQHRxkfivSrDjJbD3SvJjOIdo2eiszogdiJDz0ynblJyTD7u39
tXHhQnFtvKZIjifmKF9yOnj/VYTSPM5sZKq4O9q6x84hukG2aPahxot5diWaMf+u
ARokWCjiONk9Xf65YkTkxhqSeb2I32BY3n2WZ73tleCYS4zxBryekYNVv9335ERS
PcmRXnM5r+kZ+dvmmKIZ5bzjPnbaGeLCskJmHvJUfjtf0Q/1njRneEnQNk7APRzm
1N8zZ9pUNC46xmOrt1go7z/Nwpt7VHiBGdC2nN3mVZApMel9I2Rs9Jk2kjlag6zD
RiMb0lshU0YL/XHKMDpetZsjdM53ExwrC6hVVH/AC2h+Z8MlGY38qpoHNLoU8O9E
JtiQ+RyPEho2JRBih/zaLf73ltBda/Ja2gf6q9f1UNRb1sveAhM0LTdwh9Of9rbI
nAfbrjE3p06floudGDtzkscbR2bLDHbPP9wfKCmILrAvZuevCs4Go/9FkiIEsR1M
OhXmLdN0zWncBWzuhEzjKIIKcxqBGxG0knrrm8CZEjkhWBz+hCJC8aedscIdXAvk
Ke/XwG4tEa7aFWvY531trV+7I8N/IB83101ZsoE31O5fSfyyYjte871vmz4KoX+x
TZPoUAEf9YfQAEXK6L7Vs5Yq5krbnzHq3Uw8Rak/2s67E5Xp4m3XkfycE36o74Xx
pINJJ2Z5bw/RW6NOCVPmoe92tfBJS1B2BRlUfcc4viesRkLyMgl7wN+yfLG2GUNY
pePrRYClmHtx6NbRslr8v1/xoxnmlGVr3MvZAL7oi5y8dnui0sIiYjhw4SZJGQXo
gFPId9IS5aGK8G1HKuA+nLFVyzSvzFTSU6KvAuT7YgoYELj2kPCZDGj7HX6yTHOk
RRrEO42X3X+ECpWUO38jdOp3n1p4ce5pW7x8rz3he2oxZYThAbG5UA1NGOYLzPMR
rO8Qzc/COAwwT3D3mpxKrNQ2njPPJlXT9+yHoH4tGImWCmZtmNH+QEW7UjL22VuU
DSaDK2v2/Z8FZlg8mrJ+D+Z0WpqEhDeYtX6Y47LzXCysa6IPhCQWhD3MAfK1c2d9
LFTpAYhtIrRahSRwX90WCtic+mr7ITDJ6cnqZLtssjiesTSLWtfyn7s/9isoHuhx
TQ8N/aDg1bPd4KjuvKKSWPS22+lsUA8cqmgOq3+ztbHHgFWWZggV8cWI6BOLsQoG
EV5kVNp7insgY8vTucnUoZQdoHhVfsF5m7uT+2xK6l9Ew5Ov61T1zz3pgoXy/KhR
+CU/h+zfOjJ8TqvEzr3454PYtPXLVb4aO+U6sZ3K4xxb7E+lKVF/4LwZOqMmMcXl
QUnDBJVHjMzo4dwDms7mN8i0OOq1AAssM3RmuyWPxK4QtFI3qG/4ewi9jN980tJL
ll7zs5O08ESG+a7Ft/vo1eLlmNO5hQCE6i9yWs5ERzTw3SoLeJPqp6w059a/Nw5F
+6CFftGsNTCxi9R6jl22Oh22Tw/y0EXkUNN8nSlUOKLAToeZuEkYCpy0zH0jOZVn
f9F5uKr5fDo5N/2cpFXhiuwUtGiiA2zmWJOlaCe9no7mGMk0Rl40jyovRnXgBlEl
ZgKb+LiCViwUIJJY0Gv++AtSxCJYUplrQNi/0qQ1psBN50N9RF+piL7Dgby9y+Wr
8hqIMdvFs1bpXhtkHpOCA0GwINzmOk6tcGDlja6i2d0+yK6mFau1VatCUGb0Niz8
ICrQHjQywud8u8XquO118i6uoa7yS/mBAuthk/5n2WpYAnCgaes7bFGUP1qXTEKW
J0ZtAzOnUo730EcMkj+I8tNjLA4Q0DJ9PBHO22SHlpvJ/9mrv4UUdVLWGb0fnPzv
qU4jA8HXJHkb7qlgVdl87zLEjprKmPfn4lqvlax1gK3jCAJSNyCkKUy/jbgpVNO0
f/Tze1JbcGioyePh60eGps/fLE6Mn4eKg27ujdVWl+cwL/pzARDU2qrZvqWpHC6g
Jl/zhK5a63yVdXTa2AUzn8+stwN/S1AQEZCN2a+xoWHLt3fXy0wjAgYt3X/bqNSq
LrYzOL2hBvmGroMYAo40Bh1mE0ONib4+5yuRluNKJDNKek9CEHZBLHu5QWuwaVqo
/nqTz5BoHWL8qG3cAj2Ofcwp29dTiBIwQJp8Ddk7tkiyQWsJwQZf4bRk8gnRFKon
tAOUvorpfr26eWForxQcpCwGym5iuYtGJAHpiuEJMvmvgwD51ZZNykdUPmMmwlbh
MfLaWCYGscKxC89SJt6dFS1JsIZIT5ew6Z0v6E++lhDaEiV99iB54OVhgzlthWtd
m7E5LglVJq1T5YH/JzJRbkmLMfk/iU5Vl4gQff1Km8zon4XOUyH+MCMtwXfRDxGj
HXKyHXyKG+S9CkMksRAMbie8w75TH1hsMwkVS262/gxzrog2zO0t9otl3osJmxDY
wzYPRBiNUV42eBpinQxkhUxlaD1Z0bUdsPJ2xwhEi9DysRZovltvzdkLQ8js8na5
EODYSOVIzy4mBEn758v9cLyfosN1dfNt1AeEgnjF5fwrvGUZR0Gb16KbrKH7DyG4
WHrCo6yZePsih9XxUfjOZ+EN6sZ1dbDRaXMP8BRKOs+Od7gqRL7kKEAdnVoI2Jhk
QF96MkUHt03I/QcANAtaz9L190pUG9mzifc549xZw256iQz8U7ti4AsVqb74pQss
XRwxSi5uKKH0gwe6YK0xLOZvon9Wu44i5i3WTPa3/cNVNJBc1EUizYb171bracNb
sdBLiQoormns95oIIoBP8oRSIILHIemOH7X29L4s8qa5Td/AuKN5S4dB7cZps2Bn
9Y5SgOOLcqPNAww+/8akBbISrg+x58Gm7mm1+8XRDmmsT+bN1an73OtF2ai5VLXk
J5dAm3ppc1W5sbsydJWbrIB0ubZ7kVR22WvMD8/lGLOGJBfA6SwiwDxpcjBh+OLj
mYsgZa0SjAb+O4j0cLg+xyKi6BEMikS3yDDtJb243G7TZ4W94iizJVdnaDllWIHw
aSxb66P1rnucuParCDANj7XjIgyrw/dF5UrySTCZMbJ5+jkDurvN1XS0a9+zRA/5
hXZRxD+Uvb6+7agR60cGkc5F4unGg1uML0UzajqHfK5Dz+T2fcLdW6VcAoReSZLU
oo4rSKkdv7FDCSmAJTanBH4qjsTKvi+SMEwdcLfNqYGMlt57bwbdsa1JFKEd/Wj5
yRzj5N5VB229y+IIQttcX6n9nL8GiyX98PGXjV7QvnFbH3/sYRQ4ak+dAmsHfZiz
7hIAZ2sNADP43dV6+X88cqgZGL16byX8XQZLhAM73bFYilV3HPbZOmjYB0PVekM1
P24h9Pmh7HDhJU5iJPmNvSzsPhB3FNxS89y1pnzb4PmM7kAJ3LNXJZsX4YHYeQwE
hhNCwxFJuZT8JGBiZYQthijbSX/l6f7bTgLuolXRF3JVGVeyb5NSc2LYEbv2NxhS
hHAB1z79XFeVwSGhBJdPiVYlMxYUp9yuUYgF3FppR3NSq0P0F631+6/YA8kh+7mN
7QwodpQhJTFf5bKAexHJwNcAobnJ/uMoE+Wbt6fhaSFAoA6A43HlIrk9bcT0/g2j
7YmoX5cxfLTQbU9HUWPmIELxuQSB0ekTuebCOlCB8L23NX6mDel4FmPREnh4TSfG
1tAUyBUztdDuTZsZBZ0kydOoo/74glP5zxGnp2yyZ+2q6K/8tNkETmIpxOFfKQR3
1JOY3d/n15GJXHxn9j+a1BOZJFlJLJ21Wp8cwA/FQBoqt0U1t5EgWqmEJUV/wdWf
5FP3TVF69dRav4oHpxwAJWXb583V7og43Ka3h0NmU/N7PhyvOjRlERproJyrxEBb
ooGKvSd2M4yQjgvlSrumjYRW/IrgaZO8HNGRVZ2ijEteNyBli1w7wmNaBkur0oGC
Lb8MGbbUQ5NpVh9GfdkAhPVpkiTtk9PQ6aTrxG68cBIspygino4bSKAC3o7erv93
yJGa6Aaj0CD0eAXRqAtmbCmTMRm5z5Y5Ot4i/STqEwlraOp3c/bQRBYw0HwMyI/3
tG3AykLrULpr63LxUUh7D0N9mnnpNgQEoy8Bu3Xp15cp59SdDIZjeFAtVwaje4RV
fyy1ZF5CLsSR+LyoNo/2yjZFEkIkJO/f1DaXlkgId3Bxy+/zafRs2eEd5gJIPbdZ
1WRGwDQZGqsIB/rJIaUiic4i6UhnVeHbdbqWuXRQFDvLOhFVzrOqFtML8QxsGWhD
YeAVb2TmbeO+41l9gW/yUSefhVRhY1HZCkP9hh6MWby5auqzBn+YddisnnqT2gPm
XYMN2P7ZuYlQLzTolZtoFsH9EA7Yt2bGfSVJmAIbCQDwmVGi4IL1sa5CkCQl0fqy
cDlAHTPc6iWEISYAo2hzYnEOZZpuY3JNjGZuzFYWKO9vk8q4jlG4ybZpS9rbxG5Q
cZhyqzS4kzh9LY0zN1C36gugT4a6s3CtVIUM/IE/ldlxCHsGKwahgpz3r07U9RhV
2RdAvWEPrBFsY38AAhqr8O6X3msrp/ZY2G5XzZIuqcOeTUQ+JH4vffW/Jl0Z3Cjg
yjohdgHLhPsev0C7QlxGcDGbvSC3hn7ISxSwSFy80V5Jb4sSKV2z6GbC844eNt0W
Ll7AfMHquaf/ve7wBK8zM7IZk5fQwA93/5nekzwIpzt/n7IannhsN63YYOHy61zq
oWIDlIQMMY1twBX6gDBPOqE70vOx5DpoN+OjRtdRK4ITxEIACNCzuva0i+uOUNlK
+qp32fe6DhTCbxgngkFw1fltUGOgyceblt6N/iT3bfU0KIOAyov+Z/Sh9FdKh2/M
dxKcl1O8SrvQuPpFUpV0rgPvVQl3GzEXtOOdjeFWWGsKqTD58b/Ox/FRmqIN/a8v
ijHDDk2fO+ZJA8J5W/5A+y6deN6fv9aCmkoWraXHKcb6Kerma56+6jMUreFxxCZd
UJJ6PVto5ABtpi8hCZXYazIfK06A3Ug19yBq+hn4STTvSoIcvDcxwLDykgoTFQu/
NuHz1ougthpLr2kPMhhAC7tOzvsjNIgcAzmdyG77lkNu2ocIVLpKHn1ikjM27kCO
RDxqlwyOPt8I64R3TlCQQLEMyYETy0sZJqDtnotmTbq6l/nSqVFwNcyfm4tNwMC3
DFXXogQbMOZmv6ZQOSmKLatPm2G4DTf++tZmK1c/iXrAntDCETmaks8r3wr+pyUM
Ro4hbVaiLI1DYKd5JiBrDxhvFYPR8XvlVr17rp+SlYnL8Po3Y76Z3VHu7Y9yE5B/
nNFMXBgiZiGsna3+DQ6O5XSzO6blow1jkdPqK+PdhkD3/q080STJfNnOIIPEBFHZ
X3/NstBmxs3piGB+bJNkUpcmssn5t9w7sQ/U5M98mC/9OjvzfPtssB0UGv931y7j
00wWMdXaeQk9rsBIHlFnLtoJ6KZy6cvOVEDCfuwMm69e8Qyd6Jr2IKzRPeqLd1NZ
XTvYkzyQMae9kKMkbHGhsIzOllm6EDcyTOpPzO/ZiPd7+XLTQsDhxQEZGEBQDBG3
XVuqR3r8bD6PaNsqoOSWa3FehEWGplWs2AhCiu4/WyP8TLpwEcg3t2ESpf9/tDgg
tElPhVZWrikJRV36O942aWiuDQLlzi8jUSGDD/9yxTKppV2HozYxDwZNTPD+dAuc
S6WZbLOvSz3ez+gKtalc+zLWvbzbx9olSvrHLfnbX74OnlLxre4EulSVuvOsNbbn
ZSAOER6FkpiQLj+rGNhyJL8n18MJxn84vhNJsl9xvKmdrG7H+BZ7qrI4tAELq6AM
k35u2Ow7ijDJQTxS87Lxa0snoAZf+w+JnI9DEYZFN+eySwfKTUVxEMA5iUXevNA9
Z6soknRzjCshl+8QJM7jgdBvudPTLUklxHfABqhrtjHD6PxFu8UH2XlQqT1gtGBD
OnHpBIdqL5cxMbMENJvqQq//X0gjM4+hD/2r+I4AMOaWuxrioEMmdWFyNIqN6ggb
Nu9FdFVpdnUDArkuv33YeRU34bymmq+prZB9nl3TGYe4VkJFB84FmIef2qA6qlcs
VZxI4ecPmqant0xUF9IXf+CcleQy9yvQIcfWr/3FnXD292DEolFGbyDy7K1ydkcC
ksEd8xgq/wgu8y5R+2fb32GnEKCT4FcPGRMHHYhbiiF2gmyCPxZYlyXu9HseWsKl
LMniSqVXVXP00703qbCHf+eoJ8JTat2pwKVYo6r0Y9H8+B6WpvIj7b7nBvgTCGnJ
NgvrsftEcVdNdrbtqCC5dVPJLtrcg09zzX3RCGKBiSKKP+z4/7VlJCh+G6Se6kbi
D8DI/LmX1S/vRXgAejE4wAupVwCXZRdQ+spqNrharixZ8DAufT1tdRqDjOFKzDXQ
mpAnzXoiEDpvcKnFjDdtwTt0mhnmgf8S1xhsrZtCH+WGLId6agAq/sLvQantQXrb
J8gMH19GcsLfC7iBvsAhoPNF0iipoNrQYmJWj6YyKLAIieJBW9xSXn8i9+1OljDY
Zsxbxlc/sSZ98177v7A2t/iFpxdDtHgMzWTwBuxY6fHquRc5RBor2UHqpmpAS6GT
HnuxJN1P/lQYV3P1FZhTacO/2P0lpQ8Thrvc1hA5DpEV51Qq006Cus4B4/EzcvIt
6tqGvc1IM9NqsfHH4uybVQ2uvkkWCr1mHebwFkJzRXFkEG2RsuNqeUIMp1J9g0tq
1MgLu83N8+QTzXJZYVdk4ivGc7dJHmDgn8d3cdAqxnpjar2q3oQaPlNS778jFUVS
VU3IT9QKUT3stMPSjXeCwOFOvTsjF44wVAY2cVNiSNschuHguntgFZykUI+QZj8f
egAUqpwDAD1NSzh2heuPPQex4s4OtBJ2eCpsGk5XZCtjXTFCT5M/L2xDOiJOTiR8
uZXh6MJTO/N+c3CkgBmGr9zyPfeglhaQZUXmPYq/fnvZvnlkYUvY8QoxI55IxjEO
h2ULeno6U7g6iwGpi4ibA8DvDdDybtkxV96iZKNTHGyvU9bvzOu1lE45NGC1dXcY
vpVONW4USREYgJOgGg2Rz/nagRvT7OS+jjspJ2NrTPkukWC9l89WN1KaAOvuFrkK
4OrjFMi/k+b8MKFlrpo4dFPT8ijF79C0a1tz4MYdvH4+JpZeZI1P2DXr0a5miUwN
nw9WhhhbqkWehBUMru5AwgZfWWp4/B8lU91BA3e1yU9AJlZJWoqCMWon6mFBpHUo
i1v4eBubmLuUkOR+JRtmtBLArdpAQKeQAlIPkohHEx2/GPXjMTjL0f/VUwvhZ5Ni
j+HsYTsP0f11gp/fFujj0nGhawzSGyQYvQADk482acn0A/OO1qt8OJWSslUvoYGY
AMAm7yi+9x8u3KbmCNwU9gVgzKhW7GnZTYITgj+15vYB9rercnIAy87s8B84dK2e
MtXer7BCrtvtouB22fensPRRWgipZMA922+mOgPTThAVuZG/Z1p0N6vBgLwFnB/n
L75KoWzk/7dLd2BjNWPwVYsZ1iXXGoteKJ7h96qISHFtm8RujWSxrVKjDhkAdBDj
7+3UB9hlV8kOkzAP3ncuIRLJ+SMi82BOzLpu6gu/ShKAlBhsXPkk8ENpGIGZ3TDg
Ax1dVGaw8zRSq1RzPLRx/VF0LujHYCIA4cxqD7zsa1PE9HYJSRW2vEqwjf3W2Yat
mLLvZPgj9tuazEehXRq4fR8u//I1+FHkRQ6dPrspKx8qtaPywsFV9ObUR1Ap926Q
DD4EhPlEntvhZh5KXUHZmgqd9dEWe1Se1hQHL1ZagCVqrAWzOyp5swBtfsU8/AUM
uEADoNAkuXgognqfs/I9pt1OlhQPep9F+gS2MI+cbt5INLqOKfqagaWANg5vFSmi
IFqw06iTybz6fch8snNTzaZPyVj3eSm48ZQr61V74ETklamI61kU7MbIXQu9TW7B
cQcG4aQq/HAYMivQayrw3d59e+29o2A2BHQeB6aPSxUXr8xvPYTifVjC7YyClW4m
7M5FVRoQ0u68diSC/VJFOMIycHFLd19z6B+o1oPgzvg6n7AyVZ9eG0YeGfX7nM31
mMN7hKXPBgdy3uH0eTfgbabW1hU2kGlbQi0VqtC1tDTBvcUjpo8SdAQtu4aWCErn
asN52wqpmgj0izxRnm2VSvllLhxhrY83HU5KjMmkiVKakOcLFAeNkMR6ZlZtS/J3
MeJX6JGqRjVj+mxDRWzYUkwKbzUUAFIRgc5bvIGD+UdzSY87lfWkhaMd6hdmhtqH
vIKcsUBcVSanM92ktuvnH42kHTD1RtZELhsCddupx1Qsp3Ac7iE/KAu6HH1b8Vzk
MhJVrXxVuZI8Bx/id+iypismjZ1sjBMvkNv5DhvmtAb8dVFiUn05QKF6sCr8dDnG
oi3Q+0Oj73tIfSNLaXzqLvyrIKsYkpJjHdtseTeWmr17VaBNHewkAt7f+7Dyu3fF
bTVsCWC/+a7s7IXARDyIZFRVP+/nlYgYouSwokKKknAf+3wprBW0V5U/V+d5qBq8
Y4Yhj5FwJkjV+hBSI0aKoz9/Gdy/gGIzfWSAyIpIDZ4BP0j+Ao/pQKZKermYY5z1
2xYPpcBWfOTWX8fbe4rEWMWJUmpAIJU4Kg01A01Dy5zCo7RzUd/ko0mtLOuyPrNz
S01+KB0mElfZo84bd0hA2jW48wyqK58eBOmiFjXTL0gLXiWOa5D40kVVe7FIbc0C
NX5nqLwkjH0tQJ5hwMck7fEPxmUYdkYo21UkLqzz658mLF9GKKGmXMa/Yb9V5wQL
coyjuT7IsM8U3Nkndx3hdZW0uvlNzstIXSVSSeJL0HDMF7SZQR7zxNqyLaFrOmq4
WVArOqJc/h8CY5FAQi53gj2J4nEgYlr2d8Z8xatr3/pcNj2ScIE6YcGpnmlaLhI6
LY11kyUwSN8v68polOb5RDEHD4yVB7aI0fVlfFFLDBSOsf3kBJXWLe6k9zmx5VPQ
jtj+XXKo92YzToGVoyvqYztjFxp5v0OyOiFMMPqq+m5oQKeUstCpww38MqQTW4Tz
T4m3EjxmLFgHrH0THF+SbwRMFLKWP+w6H8FHznH6BYJe5gGcIU2fSN0Kybh2QhGK
qtnyGhyLAcmM7mura3VAPOD0hhzmIKyVLUDSOYa+A9rOIoMSwim4fxoxov+9Rzwe
AqiWfpIA9pPNFb/S1w6XXdz8bpkV0OFK0KTKfsSQ9kp/z7ToRJfZvNjN0Pb5lrJQ
65nqYqcv4qzr3PORmh2CaWoLOdXHR/SAXACyX6Mcro3NO/486i8GZ1rao7uBKRJn
9XKlisodkLiLVjbLQTeJ+UPBu0Q8Ky27PzZ9KYqQGzHFuuov4fY+VPU+tHMpcRpl
2ggplzmoMPYYgBtGpA6GrEh2aJRuvq8Lba+pvapEnMp2uhfZDE8v8K2SKhpFAm42
coLxtR9hUEosfofwcHqr4vfN8m5ZtsLu8aMNI7Je4UROQS9JO7ok09uZ+roJX10Y
FPZaJBjwqMXtN4NiATrBZv+f1X5lDkvv0fmWz+J6eOlcZiPtj+2ig1y6Ahk/lZh3
fQGhhr72Na/HggSX94rlclE/jGXRQTNW1yrJJgKbp9eFrLM2JFGDJ49mU2i0jseG
KRO424kywzehrF676vho2gmxe2leXpiZUndxl8L+MSsRM+QfEDgaUSoxvsIZnZD6
aFyvTq2ljtDKCUZns8PWkGajlvxi1Tu5icOlhkSxBrfQ2ls5QhwZTvb6g2z4Jm1O
duvhL6dWFLmW+NE2LqEAzbEV53nt7jJyhHdwcivmwjI7OoWPZ5mMRJx6w/YCG54C
6ZNmxKkRVeWQZvb+X3F+m9l+9/zHrkPQh0V6Kh5SQQhwnhv8qgPHKxoiKY+63yc7
igiyo5JsdgP6X+8GXYtRtVO4uOWEiD0QDG8s+Tvjw3EX1C9SWISK54jBynKVLYVJ
qZpPgRkdmv7p1H3X6WZfVVEUhcvOUpHo2RBCBLekXrCLW/YeogPfTo11bnKFfxnD
LJEFr6Asq6w2+9+vivoNKIup7Y/s3ebraJCl19vLV4LqJ1Tpj/5S8zklgBiyLgc6
JuoOaK1qbhQEI0r26zzSlbI6mgDCnwecwYzIaLglvNA83VgnI75VcHuXJJGIm74w
1bcE3Opm5a+AWYVg+P3HAxChWETOekYIYUq0YB1Pv2PjhLG594/crwY6bXj0wnrQ
XP3PVxxf9O44N3Hb2x0E0KuS3xfycH3KhknFFVWDz6qP9e6+1WNVSZy3WMQCmqYd
2s60lmCoEnJ7wuRdJJbDa3JrH6ZArB8W3VKGyg8Yvs5PCYdILNIXiz3Rv1H+FqvT
nb02gKSyJzPZI5oNLxLOf1riQQ1y/yQamb7bGaw7aL4PpEEiQivYmq0i73Jc8ZqI
/5k9dVJYcMyXNJi1D4c+v71+y/KEgHeqG8kWjnCJJCF5p3JtNrfFNA+0ns5UFPyX
aYaRvetdWwq+Ys0m+3UytKW4XE0TZesJAhSfb/YEq4KirK7nbuH15DhuiVCTa6Iq
gJoGYJZsMEiOxdezC3XMkD0Th1hsJ+BAf7PvlYsZsdQGcZ+j7qIeMHltPmLNHGfp
6lwPvLGTeGcBAZ5sSRsSz9bAbffVEKQjWRsdKmaWVXSxItWYumd0PcDQtDYGfLL4
t+iW4wY/RC38fnajBNMSmOHo22t+CgFb/vyBJAI1YTqz7PfG4qf1u1znB5+kZlqC
TMy8wJgFzMrOs6HV1ugHhVl7/Gy9LASyZIgH0MyhAbHodEplidKxsZPNNFv1fjmS
+WdseV0t+2B4ETPyoWpxDv3Idm/uwrOSn1td40hjX3Xv1CFqXgjY2DhKX/mTTwst
JHyysbbOGSl23su7eZAio4rSKDlGu5d3zhi8dK+yJP87IZqIWgxAYYM4ucTN9q7T
Un56vqbI1Yy3u6kFMi0jm0Ju7pGaNjz4XJCZdfT+cYQ7vo7Jbs9YUQ77RKkJwxSV
Kqh8Sb0JQMkT9cubEoYaMtPzfjh6oQXEE/205YgInfqF045SvK1qZUIQxjspZEWq
EhjLrSdhH7BwRFk6GQ7ppTMIj2MCbukng+c/AcyfK9+94nXSGK6r8XZMCLzq7w0j
4IRMEOgIGx9dqJKAQWVU31UZLk8M85biEMvGjRp2dzzvIlY8CxgTEDdluMP14gC2
Ht9zfT18EkpDmlJ9mTf+HCWI0W1Scx60p+dY/CqmQatPbe2RFcF6OAltXfQJySQU
31rqpunEf42UIeIgqGt5tNtkUtNv863GkuPstQFLYazFHXLa11BXoDGOKa8Hp9j9
NHSAomMX6t53jNyVk9GZg5cpQYDFHTWsekavJCaA10ywE4aqQFJmGPOv7dsmfwSp
RilnYdN/3nKsk3qNsAI7a9M6OdbpfjWhg+cREeTgvD+WtxJ2hT+hOzjKR4HIN01g
8p3pvh0WBStiisjaR1BGyeSTLsBBuV8vQNz/CyQdMbNEE9cPXrCECOW6189HBuNu
ZfM91yR1rMJ8rmLfnA8YDRWJv9oPldEsMGnLM4e0BvjnGr21bczbp13kT+WJ47zk
wv2wCUlt62ISfv8jzANxe2RodxC4cGNEPNQ2rImQLFsP0qVUKIW63mWefiHeHTQA
+xhIxIxmNcRdTx3VCgCVRNxiwamUL1gNG9ewCs0oujUP+CVcLEA40P9dWPNyGkTe
5InIcC56JESpIED+5HYPomwOk23GQQw53sETbhh4vv/vWdJJAsJe/IbdHaHH9rvO
cf6lEIfGEleLcE96z6Tg/cojJSTbFoSWF1sbIDLvDkfq+ZNgnZ6sZPrlIZnaxmNQ
KorrX3lsHcdD2dfBSE7Br+UpTvuLa+27SpNl5Zs8A0mt6m3USeDE27d/X0i2eWu0
bF1chnMgvDsOKEzP6XRDiRBXW/NSOj6/ei6uxNST60nZhCAkbfSGivL18JFryUzB
duWyHn2o5aJjDtFLo6wwntIxpYm9GqLzkFEbys0bS80Gndwhm2EGPz+hLD+pvygk
m53Bc6T00XuKl8s3rFjlJbLcLgVAXw9AAhFJg06PPNFWZjXXGQ0rTx11/VmIfl3a
z8Sz6qru17y9atJ4tKq1GeTibpFtxq2fFcILlovKkeIBtqtGrY0vBrxvmCDNUeMJ
72D6UHpnN4DQM9gmcjtf8QzXumtE+5LEUULf4CM7s74nO1y8SjOAmKORDTU5pnke
NjaKlA2oOvflEQ+qIHf0jzIRpk/NNw9L0H6OIb0ikTwUCHfQQKmNlN0S7K+mUc04
y4lUmWKaBxr7hgPiEuB16OEu0FyHLW2IsMSJ/dSazeGGZagfs3vIbyKz5PMCJo3g
QdF8hGIsV6RFgqHizYYKeyA8/dHMcsOqpW1hfYZ7pDX3xnfmrkAn33GGD7PTIS3u
iGusKO42mKCyM3/AYrzI1WaQycEOVHKGkbChJRLUShF/SHyoE6O4gDgkxL4c/Syb
sch3pt5Bk+4J2MVTCkkoubULy9+wgmLSP2WwONRnIpJzFlLpt7b82XrZBpLjFawV
r+/EzYljyoCJMat7caVy+gFQ7dC4RTonRkFEIoRu+zKtotT/7v8EJMtXw5a1mhL1
NI+55TxQCNeVum6TvZQSNQUM16ScYYpL/DIm3TOQdnPwtANmq5Q+maLbH84OYqsW
oiiTv9tOdlbfBGtk6LBUDrirMpzn4HSp2H2bTSydtY14yRN2ehXXWPTQ7FWuASrY
CuxpvvV+/7ksve9kgCoARrvMdAFppNKnXGsAVZac3QCIpUA30ApcHjHOmeO54IpR
1qnWFzNA9JIYdFf52Ej1HBacDGT4zUPRPAXWKiGIJ/VdLizpfoUz8QrlQJbT8kPw
qp5379zZf45h7W/JNGqwMLb3UFzfNmucOwfu2ecBEcQXiIfWmVXPjLzP/hAyov+p
QExBQmh23YqBKMGpj+/OmLGoF3ubWgkCtvi2Zcof8Gss2Oxus10AQX+eAFv8968t
yp2dGlLxyRsC/Nr0Er4Q0+G89X4YBLXYCKXr6hJJqAY14I/XfQF8uIoSehVABZhr
DyVm3oubOgBu0WVncMfTbQHXecXTaQK8hfeXvLghZ0klZClHInLz9+MpQQyG0R1f
aIrOUNtM7lQxImq+NnEeDbEjE/IOQDZFQ3M4PqL3D1TcRuBeE5G8uzVfjwYxljBL
BugY71/Y/ElI2iVHO2HKt5oJA7NXk5DfYn25klaw01ruZxCfh+6fVQXRhXujCDk1
yGL0Yk/H08KpgVp+O04Ww+jLhSHrxxLzDnwXFfymHkiuY8Gs+xEa068SQC60Vequ
jJNVmrN/+KQyA5SHuNLis8RlA45bf4gkZt7Ivq8lSP4sjTMPGSWx3xQh1632xt+c
fsTMeJj7dJh6Gbqbz09d+9u9AIbd+T/APiR27NlY+OVG08cZj/gbZWtf4k0cOFqy
InSB7QyIWv5n1DXeCxlkhdRcFVE3bFDg2INL8KGtNdZ+ptlafWznqQRHGaSOqqUQ
n1K8WdMBvrhQCKRc80ll/HQ5sueEIK+/3MhkJLF0SWJpqG50t1kRJXLmTrWh51pl
+3byNGfLnaEcaMxNOsTucOYi4aAYq7dKXLg/TQmFwL+lGYRlj7aRrm+0LfO5r9Hr
mzX1gmM6UvMOQoIjzUPsRU2NPyQzzjCsadcsVkDC3BK/UasVZ9egmhiyTN3riAmZ
bAyCXCQpm8/xoj37YTlpOP+c3ix7O5F+QsyXmqUIWpbnWvZazhgLQNzAcgeJp9f8
0aIDEP1dwgUT83ZYciIOvXcSDjb5eeCHylzUiL0GsDbMya4U2wyke54k4wBORhYB
IS51/IHDtw/7JiI7+3G0qTw1WEd2TTwpMLFaRW2aKFm++5TWwFgTxnzR62GSJE6A
XqE3p9S28lPWktUK5V2T1JGuLXDfiDdRHjiGClam0ypKTkLcXvPySdX40CexHVge
9rpRh+FczAk64DnR8BcPjP+hzMm7EB4xcWDsZzNdIQsf8ATSCimhU6xXFT/SZHYe
SRKGcSL2HBQUikfe2A/XC2kPumAcYm5A6Y9Q2sW1BJm02x7fXwF14yCt2hckGxnV
mibnALnbjY7Xe0zbNJQtUIsoajfGXOPuXEsYszL9cwG0dR6MoCZ8FgBR4cuXw8XB
z43kCRQ7T0kVgs5KKnC7+hxs4nW4Y6FszZWeFy9Tuq/JA+v4HFO0nltk4YkkYxxs
6vHRpdtYkqHhCubHjjP/+gsF/cNBAHNjTnLu96KtavbNPlhuHVjPHspvlH7Br4TG
MPpGPqU9rzKuIDplvOsHX6W0pfgKe/ghv1zsdeVw6+PYMsbKUS88mzEBz/BjRmGv
a2VJ3mJNkR1qeXo3wsNA81lHuG4a9cq5KfzlglfqeBYuXNoG/BWXN23kSpVDcg71
XOfbzB2M49O5sCXRc0Ttyr65ch07ipQekt/LRNdOsHIeLgVcG//3QD3B2dg3SR2+
iOolObWUx+JOj+fqh2OHi4gyemw76fgYcW801Ol2cRqvzdOUdJtLXv1hNF8Nfrqo
xpCzDwjLJYX1YQJRHvJfZsL7EaTXdzI5mVAEPF93nx5PAM3mU2MLjpIb5mV1OgGa
iBbSK+k/tjkawpHEvjpzSmVXQqA5UMOV34QiRYC+opXaaOyKzEf2D7Vat4KuNhLQ
IAF+JRcPe5FI7qqZs90pb8PST2AXaQQdsl8qZthPNyitYlnzXr9DkLTkqNsFDCFl
ezV3EvoU2T9K2FUXvtao/QXuOitZ1D3e8kkhwUt2jATzmCsDXo0rA1QltrYHYoHD
WuRfiaXwr/6cddyF2nvO6/kso8t8LK2QVq4DH2TZIhZf52MSqtjBMxBGv3hlTU1k
T3htaTBhC5RxYzrJ/QJiE5LyXNhdqJgfxl57ebwPEJvC4s0jybwtfvprAZfPER0n
qn/gvp7OHvocK5W3FbK5we+XuHY62Ud8GvcViJqeT7XS2Gh3a2FhmPuM5ud8QrW9
UbKGjzQaVyLyi9vEZ9fNtKYfS70rTRQaAMJQHgfCAD5LWce6I/UBZRp6u22yii53
Au4xyxip3o3NjNf83JfKKIZ/+1nA4FI8YHuhTmb0N444G/I/t2iwspYuri0Q25Im
JV/WP/mv9xb5eRqxEb4xaHjF0UmE6VW79ceURQYA4xcPEHl2oPALeJ7M4uPtf1MB
LNdFALuWcK9kzhD80wvjuNisRhcIuMmEtc8sqLqSKnCr5nTZZYBHS+5CT6J+tavN
Wn12y62nlQZpM6u6Y+qj/Raxk9T7C6dGqktDnSgU8uD2LRi3/bGi+WUM6qKSJUos
NSq7QSDoeE46gqGcqQfUfPZxHFv5PimPWUJzcZ2NceySq2V3f3OtN87VFP/kmkAV
k45SpQnXENJ2OgXkfBy7IrFLXaTb4CczINcA12iMDhyF93UJ4xM5hQS/79FfngEP
B0YmdskWxfNMPc7snYrY5W7MJE6R/LMh+2yprAIRdRHvqfcf6e6+He0Jj9CDtMOV
Klc6n7a+8VjnX3b7GTZbKyTjuVF1TwCROz8/iiZyEacm72nnXH8vKstB9H3S+AB0
JNw95d/OxaZcAnJdKQ0FTbzXmKDRVKI48k98OGh1cQaI9gZVdGXDkzW8a0gDBFS2
czs73XAZIxeWHUgGILZD1PsaO9meh1moTkEd72Y3SkM3enlINUA3EDhYHySu2y5T
Hcz6yelhbqQQnHIf5+ayfob1rbAx9K/UwguGEOBWyDgPBkFQU8HSr7tMezOuX9N0
GvxlK8iQNHAK79fuw1RnBoVGetOrTgg1YfnSOHmzLSIXugckt1vsjkLn6gWrlUBd
bBmetDsUwn0Se13dqHdaO4Wjy5LMWHbQXPxVy6DZ3VCSes5n5a24soof5ZTzVNGK
gQCcrLdedVg1Xz4CEiXyFiX8L3YZoBXsU9FdIDhdlEJcvvDGQFUlqwId0oF2Ztp2
7lNwxuVY9NY1XyVaO+C58I1zfGSbho0zhJC2F1Zu76OrH3X4yIOyAcou1GJw+0ga
wbE0UHULrBnSCQW5qm0r5GgNhNbtGE8rMp1eishS6FKqQdQF3z4YDiDITMLf5TbR
EUFs3W2Ht98ZfXO0wl0BemK5DyfPZoXZdmAOwJI71Jpemgmih93wDVLfALYQ8hmj
7cMEkjXB6b5qZ+af5Y318O/Xf8CxgW8yLayuC9yTq+qIzBhSzrVWvxPw+gyFGiNM
x/E25ElJdSJ5Cbr+8k5h35kONy2xV6MazdqmCmLRLPMZXA1NCv2uG9zYlxx/NEDg
IN3HMGAqR/2tuqBUbJveJuc4Ii3IEUQQL7hB2Vd8xaknrP0jVqLqNlZwL2v51UDW
WKh2LcU+29OGj2qWXjNuDneeaQwxJR0dSazmicAy5fnZap/WupFukrj6l4vUoJ7t
VuGWeAZsXLGqtq4LvlcWJS6umDPelHOWC46l1UbCvPOen4gPmMjELCFNTCxRmEur
nRJLL+ha16C+cOl7XkEZg/s1DFiUPXvHtve86P/TqPs5nOaz5L1DUxu15Vl2xyss
zgUTs3wx6tn5KMiwNteMH86k3vnSGBWSeq/oywko5+uBrqpGx3MRpqL4QXFN+182
O5/aX6tkc+Hs+TEXDn258HOnELXYZQgKXYlIsZoN8doIE1tIw7t82ngFzQfjJoHU
78kN4s/Jv+XHRhMh4lXBiVkWqek/JOCv7b+qopqcq4/8IMIFHDV1jNI80+pVOxF2
MSGIJjqG+fFCAvZiv7+8CFKFUaXMVlltJUHc9mLJmkyYYUnXLEcZzenrotoA0stM
F1eR/w/V3yEqfUQbh1Yz6msYxQ/b0mrDu0FwvfkauAFJlQaIbK2AEQNMnUr5F92Z
I67k6aMnqeWJ1MJkAwcfjhLK9sQfJOh+mxiiaWr6qoG9XMCBjOwWC5ZIMIqf1m9I
7tVWyoC4hVBcVE+E27aWdjt9N7YLYsrXSfzV0M0cmUCqFnlxmreyC+Jq/90JrkDL
H8nj9W5cvOIMSKQjWM5lkEKJgkqcaWedAAxg63CEAhZLJ+hDbPGxZrJNGaEB3cvG
DJSpoU6ZFl8a+eqFCb+xWczLPRr1szbuBCRtz/Aa8Z16yBaY6aEXmh5UbdC8jvjx
lUViV1eDjaLxiSpHPIP+ABVSRnxmXEtRDUe2j9olp95HSbD5SNGZBMOh77g+eCKC
8kpQ/s2UYI8x4YC07VOOuScxTXl2bKfEG0G8e2oemwsRz6rR0zLLSxK5dRsY11vs
u8V2zlro72z3ZEhxftGy9QHuw43KXaYC4g7yq3qyblCJix4jXOTMAEggI/79nNVs
KRf4kM1o0/n4zixboMNakctSoLjoj0xLUzpkXiYBL2w+LXii8TNhTR8KUbLNx0rt
PnZJd5yJ7+zdzuEvXoGfHw72SPxtkqACqnpTFDjzIacdYIi54/84yP7XV0CTe7tt
e3rOHne9Zodjmd2jbbOt1P6C5rZ/tRfGU/llPiXCMnkC92THkC1DVzRTEoCpem7z
uiuh9Ngg9bYD8xQvQhxQJisBpJK3jXF/JOxyO+eItdVASYDpGh9mR7dZwYGk4IYr
qP2llrLJ8Pk6dyr5DyKxCQWj82bEU9Hjau7HXL+F62KJWWWsioELgHvrGS/EV2sN
M7XEtcIszzVHKe/vuiGp0kTHm8Sj6VTLnX5F0WNegqLfn8CMu0yRwK4Z4kJO4G2o
U47uen5H0OO00M2IbpM5JmmH1asACMGY11CCl4qumvtowumJ7OdVBDZOICKs68IQ
bj+Df+H8egnKpmyRIIxTAMtmDcHTZFWSpKUoukLWiHukmhfkYpOosJJkNWIQRxSD
2v3ayjv8reZ/eNaavZw+z0D3zdEruAfNNRvsJQ16oYCzHiLkhhWaJYsrQ/dvFgHh
Ey4JKmoIQp5syMALDcFygpMji7KRFMiWSCvjX7rekWq7Y/p78FbmKSYAekMfFCW7
DUD6lCZ7mVL5XCSinr9wsWIjUaO8QysQirHu6LDds6dDUQx8OmTLeNHh7Fn445T6
z0ypuvra5eBCNfT/iqIphP7jewFJDzyAe0u9OsPadkG5WL80YUwMCnoed2HDJJ62
X3BFPIYFjjGptbR6f+Q9yhylpy6jTA5Gdgh7TbLp1Kr+RJDsjAKnyfUMKJOXzTgS
3zge9VRTbiXCk6vgBD/L1PGe3ihTomv13awoscgock4MNQ0UcZmk3g7vWBuPjIiv
RtrqZ5cnDvBrd22YvXWXC55xahXn2sjklYfoKa5j4Gh+1Fovxq3N5ti1n1W+DM92
QcN7zTkA18jwiATSxoqEuGrcWJU4nbAaKzM3UnNih2Roalm+wsGIBWX+KbF/vlJy
80qMfD/kCdo4U8+eRGD9LdLk4Mlba530QoHW8ceclRH4zWPIbUitM2K7iwuy+Bi/
z003VzMIYyNEhSckLj3mKkID+ZSc5T8nRnd6XfiforHZQAW2E1+ed6DNqMhiNkul
vnrO292mVz5NTvejYXZ9fquMiU3MclrJ+6NhR0S7RqMnPu/qM5pKOELr6Cqn299P
P7mUci28q4tK1KbwbCaOjemrMMSwlZ1EgirpYkBPbzIuBJATRAyCY66lFpaqTqOG
LEtws/U07p2hJJaj7dCz9vLVm1mtDz/MHFc6dSOAEgDc2KBzhjO6e75KeZUPavAM
lYkDnC8WSczud7M6TqUktVMf7eSg0VnkcU7EgDsFHpstCqxQhFnwu5DK5cq3CKFq
G/OTrQEi5a3bwPzwcGanBQP4qIF8GY+OGINeDllfMfjOGR+sFaw0UPEoWT2+bZLh
5fuUuqkjOrZyp8uU2sSAlmcvZz+58ohdXowv4JoTVKnvn7zSteBzn8x5pfgoICzd
FbHRF1T5ZyEZzXKfw/y0uWbknAKCmqCu8NpR5HScURBS/aE95gEhnTJMTQECu5/v
Zw2LHFDd0oHyT03EpV2H+9kNf9WNv6nRnpVTZF/9rpFciaQO/OxIH/afDEOfbTau
s+Gu/WkiJCFUuRyYaTJSdstdN8HCr8YK8BX8Jt7xN//lmJZ+2fCNgmrworrELQM6
cpeFjl4mYqmtKqRSe2AD1S6TH5nIwgXO80PS/XbxMb7sr09rXErxWeJxoejeNIsn
UBDgDVvJJnRQ0soLattASQNEpUg8HLZcdSjVO4F5T8e0ZZ0thdNECXVy8aohqpqH
Egw5DsNsDWD+0/S/glpYpsWwZEMBer3wbrTxlzKV/OQvhpr90qGmroGd1mQepQHx
R8u2aZU63F+PC9q7VrhCr8lTcJe9hJgCEoyZpPmKpqZggpAJLQS5bxiMQVpbaoQu
qfFg5h9lF1w2tPNSnqto6nF4NgrTPp9rFggr6KqaaoIQiMu5WKxXwNnvcF8KMeU5
yKlYf1rKQCi9CSi8hN16cmyMnnfYndbR4Q58QXcHiL6YMPBIQyduDDXEK5f8UGOb
UWWY/Xyz6GXUqeHBZkG2xFRyh6pXh7Ztx5TfwY0Mvq9MQwj9HMwBngOvZI/CKser
4vhEERl51GFEeLtMxC4obdQt/sal+sZ+Y8EeDrlqN0LXaY+PVI6HWK2io70wE7Ad
I2CAjSq7DsGWyyZNHoe0iIJ4AwcPjiT+XBVVNzsOMaq2ZWeudcb6TjVZr5YviKvW
FzuTouzZykWwFPhSk58A/h8iqBOCBbI1OU9mNS7K4foLq3OorCGLOHc2hupeCbCo
f7UugOWlN5w9MvE+Ia5L1olrhqY8Po0TXk/6CWBayMdZ2tDFwP/2JKb3Kypyx0L6
lpkMeijH65n3ELqb7PSirKWZuaCGgYD0ShERSHB+zfJFNjHBJIhqymQID+ViL4ZB
g1m3VVIf5jmnSFBqYg9ULkyPfk/AHPQd0iXY0+J4y5H4ESfGWbvGwFo6dHlANP/Y
6F67alypw2kRqS2EUCpIR/HQnMT+r3sWlMe+x3s3htm22pIHpYVlM59jvyH0srH6
htys0NiwrSlXGBs1XarfltiOoxMmLY77Uqdav01JIh2Cs0zyWz7ls58nK5PZReJI
ab/3i+4NdbGz2kJXuwaXVugEcFNIWbx9fi/8d0SuhoXEDpX4znoC6jCN+0qwuC/F
bPCATbIjaebX6Jm7z+hB6ZmcwACsVV8fukF8reHjruJXZfR9wEIQmiGRK6NrD4Jb
d6wRQekfb/2Tw40Gl5B9MNu0zTxDe5sKi7G9DHHMmSG3/IyvbZNjM0DJt6qJ+Cj3
0AcyMGMrj8EKLjnvlZgg7mWuJk5gHuwvM7/UC9waJ3DYf4HXu7/5UOgFesmQ9dHm
2vVdmiJnoyv2SP2eUmOC3fejJL57fb3uac6MGEjF0FSTK3dteGijfPW+1JU6zScO
1jjodbpXZ3paRjpIVbq7fn+cBbvIXrayGgY2iQY4448k4EKcd+a2Il5F59oTzSA2
1R7dlscanue14y8E4SHmRU3iVZMNPgcKKGvlfai7ukJBUmqe1HN86WqUuhTTl2rC
MmJ9SOgqlKUcUo2aqNb3AQV9VKJUXAIT/SXJLvrcIJwUWGJZ3YFqIOiiMyad4/ny
HrlD5g56EaMFwJGHLKEJutHuFAULDeQqnIg1xrnIJR49W0Jo4Kg1THqVl+IgVqw6
Cmy6aeCCn2P/5EaIqiEzWoA6tbtFSjCBvI8jXuarv3FR+ycoYLaRicUP48HHso+A
dDWANRxgJGwq5FYRrz+5CQa+4wa0zRk7FxVAhxDtIgNFwpjudCjWym0iCczlwfyA
+D7ABny+MCYDxotUlNDB9fVvILu4NZ0pCwXYUw0sJk6DkeG8IumIajpwvAm+kzRu
LRr8WfQtrY8AzPxpMiMYXXXcNfm3/DP9V7EWxQug52c/FRyEHQfHM1jGzUJZZEev
fzpCIxuAS33sVr8q//6e57XeiBVgkNGRYV4vb/yZb/GFPcEloxLQ/e7mZEWW4oWK
6x2aGlWyH6fuItfiHsyZpIYQjYIWbkLxGn/kSS4TRoqQLkiTLOrWWsud9licsg6X
1OwMnKp2aO2862OFgSVZTh343X6XM9cBBLNdnMph68dDRGSRB6vMtgrIhnUry7E0
oa6KbhW6pYxVPHM1klwBQy/lPny09Is85IUWQ22DwJah3lhWS7x5KuFK5wz4ngWl
iLKx6WZnIjZcGxHHvHSXvVUfxcBbDvxBmiYtHMAVUti0DctQT2q82bf39nAiej1p
724cI8K8KUylYzJbS/aFBMQ1GKuFBb/ORdbUlHBz0uWL2eVLE3Ty1ZSLy/BecIIF
YIez8GKjDjpcQLuJdp8PmRnToQ/RoNzKsbuDnJK3SeKL8NdwpshnNaCqUehjQ+YV
QVoqRV1pHVLeVFXBfKc1gsGIVe0pjeEOR33Y5yHD1nS913H92bDxMCr2jpN50/hQ
bK5Jw6B8CJ/iNhAxX9i0kOzbhOeVfnP4hgPUDNVfrkVQvq25kEmKFB6fs4pPF41m
GsXD+HetA1zic3WuZzkdxDdLU/ENOagyA560nZsxRtvqGVIh9PjcyX1V6DlaYthj
2CIuBCb1zNo/1YgvzVj/EG28u+ZmrkprHcLov2rH3AO5GfgQq/1NiokuCGmRfGX5
d3TbjDwLAtFloC5OqhuKrbktHOu6p5AnzroFX/vrxMntkhWSOkLmCn6ooSOrSWyZ
rf975UVSz4xnmhnityyXBaZLSXZN8Rw9Dc04O8MLfNt4nMyp0MgOE5ensT5tcyxb
7CSiH5zeD1qW1UKNTh9akRT0lWcaEv9P7I/eBuz4ka3JK+DXal0lGDeSyO8YAPTz
nimCFoaA5zP+Yy33YLnqgcS26CNk8sjsKc8jPr7ZidtXcn0fvz1k6VxJ6jmjkTMZ
rCP2jGsqKWux1P3io04AsJKZ3WLxkELEjmfAiekM9uV+K5a02RCCWSZyF6gVtHVh
vLbPdWy/khJrm9vdK8qQ/FeSj4xJeIRny9yQG3uT0T0kCTotmjJnNbGqPswKP0PQ
ANC+aku+rVtuAcg9JjJQGAfy2MkCBi9ybf0Sc5t24WE4PxkYvQ4uKzQaEs2j/tpd
iqBwlbWs6bXct9dFe+hCkpTtWDp2npFykTJu0ALd6CqYvd3P+cO3DtIUsnFSNhZw
VTlp9LQUiZ1toQB/eNtKYwPwD9rxGFR4YlxXsyvfjkh92ERZq1lVGnG9PAE1DxI4
ukv0RGTKgsU3zbUGbhik8zQ/RlUBuqNQEXlE7ODNNAargufyHIb5xEd0OWhOeqQs
o45tZI2igfj6z3/5FutxREOHzJ0bUniOQo+zq2FdtGhozKMRmrV7ghWrh4B8DeYW
LUYzRK4Hv+ivQqBs+WtaBk0DiCAgodLNfj0pWlm7lKxksHIfK2Y6kt1pg/qtiICu
yA7eM00OnE8bWBQB40k6C8M3Z+fsrWnTVutaQJZ6HgNd3oBJrBKwHOpyE6SR7XeS
CAWNRG9EycR63Rul+6S+SkcL7bivm2CkORpfOYeMAqGPl86toZITejxnVJHB6r9W
hyMs3JzsfOpkVzvJAgy/qG68j0zNlxK968X5krkgqwEzjDHrJLS1WGuoN4E3k8YU
F0IeJVxprEyXu+yOnyy6kRksIM8kMUReDxsxtuOSFKoAGhLUphzVqk6ZUoKh53Eh
7NoixHbhUmfF6+TR911KKIMi8PJ5TgUtrVCnvVOv4NKwCE7e1gsjX9jT8vyCz/MP
jktftH66PGhz7QpsVojQf8IoggTWUBrirhULVF2QPi7AfSzGVnDhFwmdd636Llan
w7tI6z1fsrfLi2C65s4l1zY1rcwU+WIbnTmTikNHN7JvbBa2bKwixKUwJNh3ZPSJ
0m/FH/O0fPQI4jOnvD7Kow+FBSozj6UdMJiQP4BxpDkNuwpVWV96FASU1SbzgvNv
iTvn5vTvxtsFYVoJjK8TXWU6G85rREGMy7Iff0w9JCjfR78uzWFJ1RebsOI+X0MM
S2D4VaVCx9fZrc3vYTDn3YpAM6OKT1fDKjgZoFBQJR4dgTb3HV+uTLf29z+d4OUG
1pYs3Hfg8PQL6kQU4yAQKux86pWuzFuS5cRQWPYgHPAUQMbjBIlcj3+DAtKhduAW
wtEx2cIGQAjToOmwzhmc0Jowq2ZJ/TVXs2Lt7SahG7Xrdja5fMUdL/uxirjisjti
XZa3s4PtHDgD2ITPcKPk1w7j9JALZEo8v8KpxL0EHUxEL8D953UkWT4rx5C/+M1A
wdoTndcycN8GnKCz3yEwU9hNctuVsDb+RXrdEnvp2tEymidRRHDTcvl2IDZfuFE8
x5TltulOXwKdxB8cWwlkesd3otoLHLNDeDKAQzyjwsPBaZdG6+dpMlyKTrOxfmd2
anKdxhz4XF21tFAjmgjNjezkHXhU5kQQZ997jQFXqjfUth2aqcrTsiPeKnGDk7/G
Z3ilvEKrKqhEHxUgly3CE8DoSZOQ8xUGqgslF+FwGxPK+t1J1fpYQ8ena+oL0IkI
9nGs9yLBUiwweNOYRYxq1TQ0oVRlb7CsKrUlJ5AaQTI7He4ryBYUQTEo/DBpHHwt
MBjKRLuqZGgJKGq1F4A4BiTjA9Wn2HLwkVoN1xCaCroQ0VK+k+YRMnA6BSeG/WVx
J1a9poPJomA5a9VlYFwqh7uGh/dY8/vRAdwb05cpEHXBoKNWmUUMt9pXbWmwC4uL
MPrFeQQd0DVHPdYpJLS79jnx5e8l31aErgfJJVvGjKHW4v72Qqfj0EdVkqaMjc+T
E8173v+cn9QDWmsOlNw326KdfnTmDlgPpd4Zc/9qpuYmxI7AW33nLRzAoAshmel+
psQtLNSKQqZZZkmI+0KvPFerND6iE2gLJa3GFye5/f7JUYJcCgZwg/0UJzdXVT/K
DIltTg13N6X3pSSIwr4SFAqpDXRc8NesDCDmmK6mkPMzYCVE8BLmFlv0OILVYXs4
LZYUkQeyDthvZixKVH5eCnrw9HfW2dT64wkHjGKkwKwUoOy04BM4bpnpeagTa8r2
WxLZAHK7gyg0/5ELYex1+OXO6nVW+WEJxuvrq0l5NYKNz/hPFC4oh2AfHBmKSQZi
dSmt63z2SFthCz3r3r9wgbD+triGy7S0A4qCIfej/WtvsvkXefWAiM8BxcMyWv66
fByy8IkTQySYl89WEE6rzpfKcpX089h4oy9d49/cayXWTACiZ0rAg3/VMr22Ss+e
YQmYov7B7C6wZSPdOBJ5ZkgHxZWS/qeBE7Q3h74hVNItEWo7R883XkW//W31VBMt
iHPqyOOHhvx2u0g+Gx0gtMax8Bfww0hv2prv7qGHF07cx9tzlV/UaKd6R8i1GQUj
SSWtQJoVJVc92BEl2AN+MQ3vRW1c7ugBN1QRf2I8wk/6IcZ/oGpiHZyBSMfi56hY
nJlgur/Q6k8Cw6gJ0PPz9ECUUF1LVlcQIyZFaIEJV2TpFqkCzkyOfcZSsyDUbaxP
MZ2/PttJe0XIzSMyC5dxKaWr+8+qRUGaVcrmTg4SS6gOYElDxhTLA7Jx+8viPUGn
rQNpmyABUrcZzdxEp29ZfYVnc42xN90aKBteBRpx41GDsRu4Bz9n9v+hP6sdcU0s
aKKQg2ynf9BpvIqibAy6NdMt4cVO7Rv5MJiuphll3KlLK3CHRoVjfmdJ14Lur+J/
MUERbXjI8flCyMGAzOZV4N9OHFLz83NyDPKdpVUQ3zyQrAc3ML+Kk5PrraoLq25t
b0HYximW4Up9eqPzWb/jMCuvsU3EqoRySKvXf5UrZzkTyOTYI0YerKpPQEVYllIM
o7iTllqf8YVMA6Gu/BOIcyY1vRxPaKoTn38oPItWbXAHbt/qYqPKzII5J3daKeyL
un8C6v50YHLB/DlBAbJS2szS+bti5gwquTmvXsAyk02ORRylHENK+seMfBXIpdmO
e99NJR793RaMcPsihYIszoaOUWMW82t104Xed3LqbNtBdeie/BhzOr2S2a0M/NnQ
xBfLubLWQAD/6ZjMPiF6+ZTijOo+I3Y/GnlDe3VsBIUoHT4iNmPOfDqAzw8qkpK/
6k3Ar2kYo6BzPqpg4fFDgDBLmURQiHIA50IMu86wAJlZUA7mCDAPMlIRA0ULmGZf
cI+4mW53eoVqtz0Wk5zfEF82VTvfAuw9UmnZDMW+7KjtdwhlmHuJHUD0pz3u0NNh
fdcarvL7h4XIQiEKsztK2tFKENe7AI7D3ZNwVYG9xU6s7sZt2TCss38FRP2nyRRX
zNfMVq657MZdaRHCrVdrQ1Up2ESHu+WlSZ+j7r2pxfzXi7S1NxbQ2CDFBk2qex7y
B3Bp5M09l3zuzymRaFcC1r/Dwp8C+MPtdI/zcx7kqig6q4u3jtmGgaAsvow8kKMY
w0z7+4cLoFlGakFKsExG4EFYrSa7N0a2WNC3Dj++rQFbcUlrO07WjDNaDiMiq0hN
K+nZwLgI+WsQ3UCXKyTuOq9GcNAKTV3LxDqK987iA82IZZOZlX+H8NSJa5NNLOOC
/gUn2i+31Bg4NtX3y4o9jwUvGejDlqlxDKH8O5ABxousn/HRVc7jRXNPAqSy4nV1
kJwpwZ9OGKihSK7pDZJwMvqRsIBoWJ4xiIBfPsgMtbUxi/YTn7VXZuYoc1QF5/6Q
+27isZNfaUhdxFxhp/EkO/85RkWGkicDGCsFIYGfvTRmRH/2mgsa9ctunqWUwPzL
rPqYhoyWN4hMrpusH6zdaxK9PtVokvIB+SEFTnYayRhDXO5KasPyEBmbUQc2OZpF
tPWSRodMYtVZMKqsijxrslTcXHb+TkyVvdbnZRO0OUkYzSMDbmSXlfvRwP772GFy
J6cd8XqospU7LjniHjJv7zCXOEJHYrkEQ33752F8lKiaSRifDOpv/3rlrucI8wSu
p+Yp9P8v4S3/8pVV7VSyFdNfrjEHd4MbLu36e60e1tzlIqLhJFfA/5mTe79bHzNK
JIRQa9lDDOah6glGvC0C7uPbjQHLDGLagUANvLC3TU+oK+eoOV6y9bIpbaYIBe98
ffa9MC+5txsVvgEJNeapR5rvQtPOQA/+o1syvq0oQkXdbrkVCwhZRHcdGCDnPs7p
sLcvKRdHbRlB5TRdz6fSC33R436HkTYOjgzfcFoBPN6lJscJY2yp/MrA9sLiSzPT
R6fWUwpVkl7pHLr9VSyxqjClbCf5WDHzkg2ewEktUhjhajDu5BbfjXgLnE+S0mpE
SUisQwTQGVl4O8Tiv/idRKQXgsGGOPw2Q20Nc/vRNdR/v9nJnSdBNEOMLiMHES7v
40e9mRIQTR1egXcYEnAU5OxOziOwrEv1vsuv4V4a7DpaOc2hy+52kyQPROfRmOik
LLcXCiDSdSvn4+zRRnIxJDfschC1Bnl5d74h5Aa4/f1BiLOOUEJUmZ8JxwBmGpPf
EdtBYlrv7p3acHvIJP4oiUppZwXWYZncok3r35twdK2DSJ4DuGhpHt1alKso2Itz
cXLzODTYzkV7wJJipQ9+gdwp05Hp0usmLDsX/cRcBvy4mSmpeVdiFo949mE4BxCu
uZOuPyvCvqiJ9DeNRZC9MhqcT9Z/dU47mWIHocSgyDbWjf7DPA7MclLZO8Csa5tU
kf7q9KcduMT/KxRwvYpiLRKCdqJFZtkhQrYA6eweuqeJb3UCwi1HXPZSdjDtOncW
WJxkaiDfz+AcPwDNy7AzUHjgEpajl0Kd51HBAdU4CpkuUwHnCP9v59p0GdXkKgzS
OvtgbrSc3ATKMnytFoTQedyT3wgBgP7o18QnKf5yEFDCejPj2AUnNN6dAmAaV64c
rK/aiBAmUjyka0okoyP5MUzgdnnImFdpqW866lSkGGKACRisVMTQ59L9bCnTxfho
Cd1Y4fhCegHhOYMTXTRPbqi/hQn0bkq9lifeFGYw1sV0k1DtP5j5NgaVlPTl9eM2
9mOUO0J5kWGa2mg3dJ3HbflEa89Gmf25YuHrlg258vsFu5IskHrejgjXEmvFKzA/
cT5Mg6db5ooi1fg1XUbuiEQoh+VoxE0DB9rkSy8tNcmQBJE3hj5FAyDVHpHaFEky
aGrNSFIDvKiNwY6MMJ734m5KpvDu/UQdcBFjFc76bLBgrdxPnCQp0r946MV5Gt+I
cAoGezWVEMAwon3U4Ei/S6tlDd9QqaaKQ/jtv2FFShjq0ln9KaQXfh5Wb3HuLdTZ
uWBT2REge6dlV5dI6HEob1qSVFhA07abuDnDjCFNt55bnCuzlxg3YC8HP4hKU6Hd
vOH9eao0tRDBR7wkbFMlQ5cstXHYNkOUj1KL+tUbqrzj8HdIcL0klZNV9c11afQP
6gscPK/p4JN6Rhjcd0sbMmxfGGtuDHQyvFq7OzfRsvYJrtRBsdg7qiCGS4gKrxHo
1+3r/cOyc8abZtQTTicEVMwyK0bHlc046uyYPVurFjTVljQejTQtZxjnTV9wvT9X
LlXmH3dLmYpn4fvgBk4pP6lw59FNhRGW6kqD3qQ7XAkSfi+ZYim/Gtgmz9mguw3T
bBEvS0mE3GtlXTOpU/Y6KagN6K1bMx+1EdYz1UZUHXxEkPHZWhdBd3sZ1eWqMkwF
AyBNKsDUgltVMYrLtfYexq/amvtrRvTvgPqwAPHAm4k40H5WgKNKNQ1utgbUd3fR
q/ojATvRZ0I6e0ofB2sQm1BUK1C81zYzsgHwT58kvYZK8vfqNfMFUOqfqrK0ZMb9
/3mBKIkFOJnLWwmBeB8YyirnwLtfHFwdmr+DCsAJNSxgORVYgcxvIoNb5BE2xyyA
AUnz7J7PBbghRvGLRtSZbsRQRd0SOiz+6uoqAVfJqkQPPKL1Zkdd8mM00ozsORKD
G3VCLDLvqmqBX3GIzXLdFFcE2+0tHE1GdIlkYiXNxO9mFb+eLkcHzDkgoNWXGEsm
07+59d/dgtcZRJrzC+AIEYHJoXBoc1grI+P+ipKxZFau88tkCJXxTN4t5sse58Md
lj7ROs9VXwU+2anWPvptfmmzTfoH1EXBQZwtaPmi6XE9qXy3svSS0dke22dQoBEJ
AqvF0iG9FIb14sw5wkPYaj0LkzfcWL9KENkEz0KaNTwhFS92tUEonZHcF/9gsAXc
HJHVazgGRSBMm+Gvq45uPjKjB0iwPGc6dQhlPlqVFEC0V1dEauA9sFpfqWDXzvid
y8dkYhLiPvh065efYXZuZ17asR8Z/r0WXpJwEg+cIupSN7SboCOhkFz4kwwM440G
/ogjItMzhJ3B+d6OTbz1das3fpvnMdomBootTSt3FolZuERRtAaqH9xmUq5tBmNI
eiEfuiyF+VIUPk4obuB3RxGo759u7J3p0QUn8aCt2+x0y9Up6tCphmfYhekX1K7B
nqgUUeVLMw6nmioXmU4gYFhKE7VrgbRCap8syyYit08BM74xiXcNDWJ1ztXXIeHV
j/rgUH2xz5OkRezDLrqG+DvR1hhFWGQNplB+K07bdI04OoUpRMl5CGEvQdHfmhg0
3EA9F9LR9Vs1o/89Rwh6GCDHmBwOYYv8reHl4LUZa1v3EggbM49UaomnMsPnDasd
cGWiRNqyBfZGkdQJdQf3SfFlOOLjPOhfuNeEluSBUVs3sOvOHKcey1nvFAG59NUR
aJ88OuvOlob900bKYEueCQFR21FoBgWR63nAcHX/aB3WT35mK//dLUrdi4XzS70q
iOv2VkZFBSiWmaGYF4OUTAyqD9qw2HGDNn/GREITqn8v26xBdAclHF3GHRl+GcQj
AUGA+4q5VAf2uV4j3BBnA9cp0XieURIUM9SzmZKlIyOUX2MmUkThMsfLBhA5nyhc
A0PPQBS+YTEwVwKA8P5lo8Qk/+kkBW/7GfsbXwdt1P28HzLVBtJpxrziQUH8duBe
ElCHiWI5BR+8M7FttZ0q6yoCpussgiUXViSYdzu3ro2UrF/kT4Le2n/LBn9/OIWe
62Q7Ho/B3lTSJeVmhU8DAmJAIdHTaAgC2/2eDTeS8hOD3WuLtzO9rBjQgNrCuaGI
aS/4DAUtcCdeu7SIrXhXclyexEgzv8y9a9KxCtotjol5ku+WY4v0ulu8t30yTgHJ
6gQ/lgeTGylhmp489tuxN0657wTZuzdAyTc5sQqwgTFonB9IwBF5QlFNwwhIxNiu
BNM3o0kxI193AdoX5Y4q5j4us0l62AZmM6avvhhmi5YRjw4yRF7oZKGLJt4ih3qD
opKWNDWyiJ7vmpH4zlw20RQ1wPKLBazdC5qa7ybSZo9DWtt0c5Z6BOaWSfbfwHN+
c6ZptvU+Rkc+Sz58QZaZaw+M/4QBUAkfnGhCkdganiZzdAx4aeSoOAQIiF6foo5X
i60+gBpeaz03ht086YWjCdmW0rGKMZi5r2/PWFNXM+QyTgEyPuL+ddEii3IVohyh
P/9erqIKFEpKNNwud+K9PV2dJlT02JltbXOQYXpgImxm6My3uMnU/ZNMRxeq5/gu
w7jekkC2XUNPJcvUCnx5z7ESkNIra8Dmee3jqERCDj5/6wd6Z9wkoZ1+czBevkHx
EFBS6vAnh8DgrHbxijB3ANWjgnLgUnXFnkYpieXlp0az7rwfOAv9j2VBfOCVrbyo
V9OCYq18hHhm/ezd4G9Mu0eVTRz8Dj+8aasmSMnu//m5USmWTzgfjh7YK+rbzj/s
c5jELrAeSnP+oh+7fg64J/Aj//2oiWXkgg/nDXsnLsMyFFDR8hcwGwxW/Pdl0+ND
rUQAosoEWXFX/4BmBbVmAXAuTENORqLu8+lgkwWL55Hn+mlJviIJHPCzxk80cVet
WJziQwamNR1oijVByk3LlZQ+l0JTMucB3cKkXK6aaFriXU8106vU0tPIqHCcRoEv
7zuB4xw5Hpd9aF1Lundj+GU9wxQ84a4HoSvW1u6jVtNSsNjSlEYgp5CVM8067Z3i
V/sFYJDgeCfl/GoOCooKLDdH6YSVp4r8mvQON1qgmlv+4mBuskHT1VGScNy3zoYL
9QKaZLHnTVNPVYvet1wPflxCryDQTWHl3EhvKdum3Tr+elZGgetyo/VPCr2qUMTw
uo1hreFwUahkW3ys1ZRyZV6cMQj47kriTuzd6ABxEZzfOXMfGstLz0PUVET40t3W
tGVP743B1fZvBXgo26JicQnq9PWvSzl3g9O9a5V3jDh+9/fYhaxjTXUsaAS8j9j8
xAcHSJRTOMFnaSocyz1h/nPcjwvqR5pqTTr+D4iWqRLtZ2/Q4De48ymE3hUaaPfP
PtMi3cqbUsjN1ZhZAxK7a43yaXYt56y+s3ypoYb08xFv2aB1jAxYmIdiyAbizRfl
paaUxgsiuQri7TskRzuuoW566I0WbtR3JgS2ay4J5E02Gsi62cv2uZARB72FfEwM
fTpCxneeNtDsFz9Hr/qG5oJ5X8cAk1UXT9HzrvOScWTz8EtUQ53Iaeh1T3ewxHEx
EA4WGjCt6ZYxC/Bb2/6JV9U2mdvG12V99bW0kVD+siUu3TSqaHZn8ZlO+cHjferC
3X3A+/p/gdUPGAyKnIIeFFE067orkhzHGvK5eqkuLaRMWt9B4JvTcxZ9YminnPC5
BtSoV+5ybceLeE4tEfh9Zd9WQbq+Ponvnl4ubyiFlUOhAifMI3H3fry03pRVMDTo
1W9pHrm4Z2YJ9EJyI5Px8IrMcjzXWK0AcMFSpSfo5ksNNAFbqsFiB1RJTAk3Wv/c
Pv+ZKKpSHxytjXKWus19pFHfMVZd4vuGTXQWiECpgyci8jB9SZ1V97h2iN0JOgJY
/mOTEyRQQ5Po9Fan7SbN+WBxg2S0M3pq+UkVvcNRGMkhwxreKRSsfaO9PoSuDSNL
ascFFbuberdbTTnC0Vhx/woafbZwrg4RqQL4g1Z2kM26hfBzVoYg4odqUqaS28yq
epLVs4nUTz/CTRA4xdiGwOsp0CXCaPyy28d7SyHviW/ad0nQ0z1LgJ9OpEuff8Qx
d5G/stYsyQ25ZC+0BQOtiTRas/OD3JYu83ZPsZRe/wPHvm8+AuLbg5OsK36tzFHA
LCb6M8YCiZ4sw3nntDT/uTjQXQSVhetnwwy0uDauO0uh902RzVdbEnR9O0RJUJe8
/EWOxHbVp+tbZZmqGpWvvWp5FhFuWksGa8LJ6xcB+askNYKo0zMIHKKP45UmWM5B
ZaLO4HejmzRPaExNXrU3VeAtXT17tu1v0Tvc7Igv6o6aig+mX/fN6bBt5bSWOV9Y
XgDsXKRqTDqqR2RQ7OiH7oOSBdfd8Iyq4HL+88VeOnr4bJXxuJJOOi0wuFhqMZGz
2hGkNSu4+Ilmqjd8EfXd8m3zYycauvCh6bpIFdavmIXi8kkAe0Rsj43VboxV4o6M
fSzbTd9/Aa2vYDFtEwiGrZoPkkS6M8qMrqRQstURCqwH3Su3DkNd1oExerjH0jq+
bH5rKm51rqD151Qx9u9cllwSRWgKevicyj526yPuobpS/lNp+eQgFVOFHJ6F2H+r
xJuHltdYmlIKs+wd45Wf1N5eJFgWCpxRJLtg8Jd41rz6eSPIDWyt0vKXniKKuDyn
JOzX8K7z86ubl62hEmTdymhoDaR9SpXIbKDevZ21+5zaUNqKLTWekRFkFB++E4/c
MxT75dvCnanUdBmTxPx1W3bfrsXwbBczh7SSfrR5LxswpSF6+Lza6SE+NJl/doVi
5yQ3rRL6UqfEHkKRgulAFRDc8ks5PoW6NQ6ZQVUqB76e0l3jgIt0DQanRtKXomW2
5BsFXJ7smV6b5gAcyyTO85M78j/WOMan0Qs+Q4tK0LkU9uJUEZhbsGK213Lhcoql
ukdxP0SQ1wSVhPTiJ+Mqc+o7v+L8C309YCY40F6I+e4WW/YPZPAwrYYmuYD9dXOf
hs4Db26/PWrE8eL5tdhDmNECn5+srcWHC3YAFELb3DtYgxQUsVTdRVSTimZGVw5k
wIXb2P0ELZky97PCszt6ZU2qp7C+oa4oEw2ZJtViEGdk2VykylZEaiHRdReWKfdj
qnCx0VwZYkvmQ20qno8oDDEaPoQI1CkmQWqNdvzotFSdoW2OaZpRIuS1Frif81jh
Z7tU1I/Dn7ZkV5gQLtlWam7rtAFTMBp/mBOoleoJpzvV/7UKRrLrLUDhSMvZS8l+
tnt+KjZvl4khw47zisD/YzDbETyAffY36APoq4+gyYmdcxm8AtYOmcknESZhzsjW
UCnJnUH4/ayWJ6sy4BdlC399BYPt6bLiT1klM4Xy1Oc6073IUiA0xYYP4zDi1CYE
Acs52wQAqpjsLHUSHYQ1gNqeQEu0OGFgDinkpesKfJzAaTvXKGVQM/PlFBvBJp5f
eHp/mXEmtCmDBox7HqcXZ13mqj6jILTD43pLS8veB+3EHy5zwnCjoqr94jdv7+ro
NivvNPdkjJtjRwKbNEZN9txAuLBwrxmxHr4a74wB9p5kYh89kbZ+AIUY7oDJzp1x
8mmKCiTh2SG8K8uqAV6TZJYv28NqEZw2pX3p+N0wBxjmKsFaK5XjeYSZCD/c0ofv
f/QhayOgyeomnl8JsQcAxBt5yGLFNWJCuWMbYs24ASvadOs2/WaO09wWX4g1F3wL
z4Rsfnu/ptXgY+6OVpeD1Vyt2y+ywkSrsB+1IKMqB3tbQObKJDq4wacnExbyAk7B
N/0HIazeEUQSnxTEDSx4Zm7giWe4dwWLkfJHh8HvxBabOEEk55PM1fnpN5dnB572
zueCZ59oh9pmXGX0yU/PMWUxcl5mj24fYhpbyO9fMV3H6dGVvPxouTIdyy6t6qbh
d3W6yz1Zg8Vou3utstmoXmMcvdg1lCIyx9JXu6R5eHetNNJHb9RkjGJd6JP9lty6
k9B0zU8LElid251i9u9KQFn0SvEMrTGK1MqMtJYC69BuzKFGZOwt6KMG2uy64P76
TwURM9ztXnPwK8366H8SB+X+gAWwUZ3JbofJk+KeJnUvhCiTXUZBbbgvND/WpYoK
sugNHaGjdW+8U/F+ZxRPH6aFJMa0UDbzJrnvUYkcvz1TnlXA9jNbdc7wCVsaZ14h
K1cOY29eC9our5nBg0ZXJFXXy327IMtLqyxVf4NrmvRDe2jUFnYQwtUPX0e2ELMR
B10jo8+MpurqWD/ao1Ena0SZ0yC5j9wMugFfco/iSDhjy1gz/a0kdO/gQwYXAjU6
bYxb4I14f1PrD3kxzUSUAU5W5+MIEo4YG7P3ABwJ8wd7wmrFllmUVUNDLhtLCU2h
8zE9lxVocwrMFVH9MScaQxtV1AhAL1ygN3+JE4rbdJQZDKoGOKmmExlRWFDjmYo+
SyoZrOYK0PBx7MhEZuTLIMD5W8t05qgUwcgALS/P2uViLAsEnKM5/SZev6FkgVoi
QgXMPfSFZSPe2Cxs9YOe8hKnkgSa+q9Qo9V17Ji4X4VnLpLb20zct0vDxEiR3HBN
pHpFRv2yi0TSc4bd89Y5ilOPH7Suki8E3ojulkoC83hzVMJvEe0uCELUPssiOYeI
ihg3jLfHjANYDouweS+IzALKQZ2fQpsEtzPQIZZRFhXVhtQXxb857EXwd9Utr2Li
L2H1NuF23AcUy0trDrDuqJZNbxGIt/sciHwBVPpdG3wUsWLjDT9YoQ+I0AXWrB3/
dTGCetGxeMH4AJX2BmwKDErUrNUghQZBE0z42ga6TMyYhmnmzxKHSqBRF6DYuN5r
01xmfmCR8qj62D1JoatGFbP4COM3ocl6XGYMlhiG8Lm2haEvvHD10PaHT+4sXf8K
2H2/gc35iJI1mTQei73ZtshxbFtFLS4k3az2Lhwlf/pQc8leP/Ja6t/+DKs+AiVD
cf4l91iF8C1miYPE6wulTgOzALQJWhYZ3pGJ7DV6j8JF2UM01iYEGhg1EdaFt15J
LoSTvVHCfdWqPsStm37cYAv2cqXeWuqMHdzPl2/dnxl38rSrNG9xlErzIK/c9kbw
8rBKa8eYkqNLGQ0dElryrth5sdCFgwBV+kJCnBt+a3UoWX+rs4cUWPI1fFwTTEHM
w/oGoIAHraX+MSlZpOAXcdj5m7KFRTreVp+zpgPUnHvW/gtZAN37WxlB1MZQaNUN
KMfFfefyhww88sjN3w4tck5TONKEwHlNny89I74MlOeW9FAxdVyjoSwmNFg01XW3
Jhy3bW93Rl5Cd2i5QiN52ueJSgdXFW3BxPEdy+bpsmZDRIehZVLtIdbbCPbeCbcX
1nSrqe0VL23ZBs7jDW6wOEm5pPfPCou+ygFeHr3BNBgDVmEudYE5+LelcOEWaLgd
Rwmbbr4De3qbpHV+CESKU3vgnPUOHceVFuqokko32qIJQe5YJO0nAIqG44+T/xvK
lFLl174hHFJ/QCd2fgMMofaiESoNeyE62DBfPzsoKjwTnlbfFgju3QAFujzzTJoC
ylhXzCwumOjYJa4I71aXuXoXPZqCba9sbmhwDXGMHegHiGOzI7PVcvK2k2t777IU
UjICVM1rOuplcMuI2HLndIPoeDCyd4yGf5qDjft1ivfjOIGRcFxtaPNVFb3rP75m
HGDj62L9nogBIKKyMxB8uQVqdIkc5s9P4vzwfstWW51XnNLaC/n7dI9DhD5a2DkP
xZJWhJxSTk3VZuyAEMluCDpVoDCN5gPJ13lr/4RyHGhx3YzyjfHJ9U+qmoOIpC02
1VEkfmUjrN1X5AutHAbeoPXr/hFeOkVPoLCdCTnFGAWpXggcWCmpsM+6ahr4WFLL
SgfNpsLjXKKNDHprssOdkPtTmaxNtUwdfLU6p55Bx4S/vi5Q5uFmbpmbNoiGfGjp
Gi8qwtjR7uh7l5w5BrrZQKUK6d3+uz7cceOMnm4KM5YcFx79cy3Rxb0T5Bh/C6dR
IG6sYdT4SdBU5s5JNdaz3H/tXVaay6lXdOrCuU3K41dylluPzHGaoMqz9ZKdK7mh
bBQJbm9lV/dTfB3i1nglb/ftcnNnf6h2idWiuncxWFThQihNjtQbgEOCbRMtZm/q
8D8S5FpYyjOhWIfmSdYcvl09AMEuDQwQmjyRNJ4XHm27YwkHTLp8HYCALCLxFrvJ
bI5QIr22v56Pb7euRwaoBZcsFt7TEqXclHeMqbb6S04YsTNCf/y0rDMf2pcdvsM8
PV6bdR0i6TTYFAXo4jyLHsReXhGEZuEHM0RZoy6MbRkSAmx8NFRopiGHEafCL7iW
sTCqaDEBpa08UMVETAQEbv4cl4P9SAX1humpHUvOFsrfcVv0stslumisaqy3ADIG
aHe1Jo/5kN3iMzEygGxpphrZ+MSa18eS8NSEwQ/9hCEA7UckswP8X4hx8Cgp+eKg
tI+qMgxkQddpcJ2gD2UeL024E0NQXl6ycD7XgqEdzsos7iX9ZL1aOHCnPWAB3CLm
5s67p6hFxn2ZDsOrJzCODKavPucwI1L8XmJIx9+tiC0DSK/Tr/CdaixgJL4Mc4Jg
Osgg/HA6ELaUGkpoiu5qAD4oMi/RV70tou+eevkek006kOJPXhX2aT6SmPQtzXbF
RQrQAHKQ4FtB7PU0K7EwwDxFCiyq7OviRTAHlPKhTiJ6/3lZGHfojXogbriRypG4
DEI4t/Sapbz3OD2y3XvKv5R9SlFP5xGME+ErQ23+ooASdEIPmBNnCCVAbihblPx+
qvgn8xXUsSUxELM4G6eWrfxJGATn1IQrxxIUi7c22z7BdvVYn/Q7v5/sqBCjo6lq
y7fOewv0KPQykfXkKUgL+xtQvbWkqZaO3PDFN3yhbXKYXHjKYfqgiXNVVhzxB/5m
CvBOjxjBIv1AiwErm/wX/34M6LJzJWeQ1OSOltwTZoFv+LYyNHY1wKQ8b/+G6nZ2
t3BoTE4TbDrZ6or8PB7pxq4zipS7lj93YZfTmBBgzFKgbkQlPQbMterVT41oPQ6a
r/1nDLWzw6dCgGqQgddnFdJQloKA1ke83XAbPeSOJnmIuAWdYziR6EYPzjyyCizR
exMVVeEkhJ8Em5OhpoWVKuiwVGl0CzPe7oNyOPEEl+vSiBYLyhzrwrybl6at3d/F
Ncd/0D1uxHW2dUNvzO0TErOnigL7b/ClWpgSUbV5N8Ts87yVz4dpJ+COmgn6uLo/
ZzSvfAURfsj822+HU7HdHMKi/m+dh8lxWnrvxREZmL2UmDuX6w3rX1ZWWzKizwoF
F0P/JiMLyGJ1KLoNxmt9e13pYdpMM/Vc6tYAfqxnFbDCKrl/z0o70eI0mOzJljb3
KNvflwEG/bWwzDX9yGJqUdqHmrHN/aAZaruPzjEyHVZ8Dt6e9KVTpE9KZB7bYWuM
8srvtAzjRMQiovuL0P72nAa8cp7i5IQWfjP/RUxjY4kJRg3p1jBM7F7uofYpV2Fd
UrSmLo6kUiOyw+RYZ1qv626Rofu2JvE08DBFea35b/dOKchSTY0Rj4fx4iYXnFE2
XW+B7eqe2fnlG+jYwaK5WNd21SzCewFCT+bJKna/nNGjoJQm0QLMyK82NcTFmY4N
jpMt9MZZSa1Isps1Tjns3AuCtqlYfRMa+AfWSoOP8Mjs522/xkk3hq5MQzxUFpI4
m3aXzrhshm0Kv1K2ej/m6fBl8atPR7FMINmPcDCa7JdeXI7yrBld9M6WLczQWMEe
JVVSny2uW85XwkdRuSodruyIs05DTopn2PcS8FL9oDNEZvoZS0H3a/tdHAnS1LfN
NaG4KflaIWrQ6OUnvhRQ/txmK8kWpNZEuXeURIpWdrM8OosIIjuW611j/O1cUfpz
0s8dDW1Rz60wgcbWb48FyKk+cIrLEMx8d4aM2u9Bt8DjcQ91jrlspuy5Ez8ck7Um
eKOupEMGw+MvJrxmt119KEOhBSgWm1h/k2mLCizUYAJNw6SCIMFKsFRBpKXcZYB9
Z2/a8bsjsuNXuEY4IKSxytg3VM++PCTyTmxn9GGGAdrNz22JfCQLsiY3SKjlIukJ
sWMuTB8tJMgalwIexOJlpvDPIf70XwEYZe4aPMJRiYX3YCqj5p5n9JKKrHj2vi1g
OQ9y+LrL255Il7HpzDRvGZaSjl1epe+ZE3+cGOJbu2szkpZKK23ACUdgHz7vqtcE
Q7LSHJ56Y44Juf2jPIu+S810RF7Rqe937eh5OSfjlbUWp1ISkqmbZy5d3VvmDXzI
m/ZYgiSZ9sMklegFW2Jy/1vuqN8wBDog2TAw5v0wC60tj1F3AL9Ju4/xkKD5DuUH
CV3QT1794cIyQM8EobctCHuBYhaRUByThHF18PkHmU7cPq+sn9M3IB4Yt+K2xBvz
sy79G+bGmj+n9oOii7FOc1gjfuL/SSQk6DMtowwwQ5oHJ/U1KN9tAOWZL0NSZXpV
tg+lPgLcgz6g/JcGtREFYIlgk37G0qA378QCkaodvQhwD1FWBg0+6yMYAotGwGgs
DD2hSqDsGUUswnHbCjiCAYHw/hzxy+ELzQJs79yRrPOrHHJYyeNQ8K/UfE0av9+h
mhI6LElbLLAq9C1ZO8o7GcKvTKOk9tP+tO54aLw9oTC00vBcEJ9xlr4ETXrPxxef
3n2urjbz9riCstYyASbYQjNjjMJZvKcQSS1u8NYNKD/mYAf2bnfrxjEW/iUbu0rc
FPqRApIX1QBKAVhxAtdZJKvKQ3xRyP9RH5Ezp5pHflR4XfClcbv6zsT1ZvN/0epn
09zQmM+oBWacasZ/SMicxepdpIkCQjDKe9sQBeaVl8LsRLNkR9lPZn9Be/6dg0/r
374+QW7Uxo0T9bnnCgh5kd35WtgU6cih45bl7V5daI3XugFeoPdQXXs5HosSakTV
UNnTj5/iiIBWoRUtcGrLgQ0WLE2vsK/UVrTbM3e0xFkfpBc3hB2ee1JSoKjXJ1W4
prfyAC4dWBwzDdX9yZlRx9F2WUMbxUirdGQvxDRxaYxeGqIa4be3MHrLMeKunqVB
xjtsj5yZy94UZGWMm3h16TVeQyUikZuGVbdMFgVKvK+QpeRfxYMWdV71AbC/4p5d
Nrx8IfkwGGMkzaxAKb7T59vjOtp4tVKAfU6u7zxkZr9kPi08oAVBPQ/uLpNETdA6
1IMLlIvO2Fs9WxK/V8mdUgsfaNTULsv5Y+tsXlWAFQQZBJeA+9rokzgP9OCf/y/s
TKjyQpHwB4iJocUHHzSHc6zIPaUTAaAZccK29rC9Ri/1jMXUQVmFXqrpUMxujAzg
AoIulgRBo4zkw/dUA7llCkYNyS+DmCz4sS+BUVT7Hitq03lOCTr98oN+j5Wg56rK
SMyWbtBugWPtlxd/8tuBn+Et2o0YYshK0YRBmdaRYfcHpBmaYbksnUvWrMyFWKaB
FABPIHVCZUkJIPmEzKb9Mb2suXJL6gChp06M4MWkFmfytFQZ2MN9svyvo5ita5OK
TzTWAXbXJYQlBLCr0E3qIXHq4+kSth8Rttw2umAiSFPrWepjEpHTInRH6luGQbJ7
lgafW61mRqtrYWxWT2GeZRq0w6yOqHMMrND27eihefGoY3dY/CzWeh459WxG0b1K
zGhacuCDvGMA5Tg3uD4zjjW3X/VWwE9AAd2av3XRloMD+bllikOeTTxi1M8CSUDO
ydTI9UruwPUX0ZA1bU9Lsko45vxUGExZtxBPru4QpJSXXcmkeuh/fu+bnWm2u4nA
7VquWTgiR1VrV96eMUDfWpLeEVPezMq/6jSMP+O4cB58xRUwcwvc14T2l3507Koz
xDTiWVS3bkAvwDIIdlQ4yr4a67WEJwjcf1OALLssvbjlGVhwkXgb9PsyOqGTz43H
A70wxNY23rvJgO//SIXtcCNUYWON0uLfNGnfz3jRvS1tVbBB8GVvu8+2GYqWjzmf
lRGojK+eA98Q3gAMG6Jnfn3WlYpd1K+2xTZTXENSkZuP0H79bwJK9sL9jary2VQX
+HSZibxCD7E6V1WuwN/KCdArID+ALoCnwIwC1IVhw6WIVWYbAGx2aItoHPS/0BKS
u92LUvPAwMNevI5xk4DJWGoiylBO4NuV965OT+Xg1XvaCeDImu/cxo13VCDKRPPk
XWBdu2VA3gj3Cfu1HsW0zokvMKqWnVhuwYu379eLCaxY6+ZzLwTtCI5CBm2jJRLX
5xXL5HowxdfThb+zzUNSJhtbH8oqF3qL9AIgYSbMyWr4jKsESqkAM5nOnG5E97in
Pb/GiHyqgWo4d7v1XSYpyBuD9avHG5rOJYcC973hdGFx/U1p35SUq3ov12DwGNyA
iQf1SnhhTA9hnbM4rY975cbbt8iC5VNEUuq4WqM7Kou/hsa5mUsZnUdrw19BpNIf
LgaB8EWBTmlzX352ai9XA6ZxSWsS8KFxoZo6bkQDbpAjJSJ2gGufOLDBY6H5Ejyw
1mzhw4ro0iBf+knmZ92HU4G8YAaoQHAGQDyUlhCku31cJlKsTAaLJVNkEy49U7Ld
xsgnSMNNaGMJe0eK0GBar64Tk8mZOfGMxnkvAyRDsHbwtPY3/ykw2e5U5WkESYuK
cHVmbZyELE7E3UnTn0iHQO5LO2HFOarx/ZUrfa9hAWLOV+glw18yrXm7/CULTG1S
1txSYIUEF1eL42ZJlMWN5uuvPUq+sdMy0DLkrDxDHA36vQ/8sGmGhxOu5okWFjGt
wJozjlZqIsz3D0yTXZgJIOTfM31xLDVOjyOA/gUEvOST2RHwINxbdieB8/m3xMkE
oXvzGYyMjXRmtMtY4gP1Jdvhn72eHGnWUigI6UZiYAT33yaqMCSqE/r/OHf/G8iF
wBcma+ig0/Hg/peJ9HUSkiWz4Vkm+eHKfpxCC5wfbxXe0CgohWU66CqgE/x7I0Wu
NTZmzrzp21D8AxdpV7prS7fXoiEB7Q+VNSXAxoF8FtPbMw5e0jnKujfiqbhXGuDA
eg+fjj7riXaNTcizdIkgJVo/dBQ2W9+6q5Wir8kGE8BFLA+AfyqMfULXUerFOTq2
gOC1IJhIHJYk5D3kt+913W54XhtxAd4DorsUEWFTp3CQH5Bf3Jl3krWWykaLHM7C
Z9afqERhpm6YmQUsKabw4bTK3G0dcSpMVMXB0Q1pLPq5mtxiLu7LKLcHjpVBZWWP
W2NeljnCf70iOlGQKPSh9psNL14SLRkInuMYwsIAPxy7a2Ulpu+8vBCu08DvxXmR
bt/DwcdwID3gQJ5Dwh0eK1I+NQnqqaqyoiMqlNO0UMOIPttM4YTRm0PlN4ZYiI70
5nw2WiwgF6FS3kQJ8hqKZblevCfRsxCb51RWR/MqvbsmJyXNM09TjeCBjaINxkUj
Qbr3KBKf8rElJOo6LJOGn98pwf+C4IxLF8zJjioPDgeuXn5aEKipZ8WMke2ph3iY
ppDmaVlS1EGVsF+/j1r8V7PtwdedqstFiGN42CDH47SkxO6/Y7yhsYk1KEK0ulAy
tpZ3avkkoUlMzd7TKQhNm5LmHLgKzNI/b5DSsOvdoxZnbYjLHP1e7rkjxWaxmbv8
LXd+6HVsFOsIuY0b/KxtoHOhy3hzN+ab78+SMwetUlcpOfzRNWbN5EBGJm5AamTW
oov/wwpNBC7X5HhdyLtV2WjHHmPFgtIxZUrAWAPZf1JqEYWNjstxLMNel0RJ8xsO
cgRjq0rTqvuyf2IYn6lJZ538Xmpu1O+rqQxEqMtFZfexsYqLg35q24jrn6oxcnmR
dxTpBOrPqH8NaJkuCLYgevtiVqE7K6E7MKw68vzJiqcn01V+jN9k9O6V1/Cgflao
BX4x78cYrPF6jrbL4m/6Zy4UOJOu8lveNHX1mIOtplXXBATmDQ1pjF34FPDGdHul
UPhujyBgFP275cj33NsTs4XOTb2O9SZ2/aqjblpjczCPpbimwvkP02q1/GbFIwlT
0oi8NmRCFAnz+VU4dTLKWYGedJELkxh6S4ls6R8furytF428qSYdizNNcbA1dpeA
VtCfujPXCXaRNpj3zVJGyrh12Vr7IFcnLMvqyvAgitapn0aS8sxKGBRnNuUVJa7h
kBjdoLhZdXwTmMYOBSU7vNgP7yCEW9djGIb3UiIHv89oOOTxXhJCpwu2KaSrle0u
DC2Qf45ttybypK1TyZ8gz9IbLZr68sUeJ2A7H6QQCws0urzDp2075dK+AKb0opTI
x22SKXA+xrC8e59xHp9/8Wr4Xf+JIeH92ZvHQuZpEAqFUX5l43RUNKwv5cBMa1JB
1w4qt6cqAAXzWabQrJ0bBP16kNOnGx611sPAsaDyt6YUt2P/hG10S2JrKJO4/LHT
WnvBlfxtbWalgIMXaJpt6Z6XM29uwJ1rX01N0/nsWppSRM7dMX/uMfVRWqQrBjTs
OV6KaRNgx+e23GynB0Jtah/itgLRa406djF9sFAV3fFaUZdi+1PzuvxFzJpbVVfx
HcgPtLXK2zkBaw1eIGC2x/cDqJDKUjja8bacOfipFCoRtL1VrRjWj4HvxbK8FWW6
V5kdI9Tx8BFVUDfcFa/hPCS/9PeTaX8hcM41TJDFwnVpvtWXW1luUsBf942sKzxV
HxcGhflOkspYyYsnImWGE5Vds7GgmWN25e7o8avXw8NVnKyD19OvcgDBKSirCC7P
663GherVKC6jNbO2zf3+WwcJfhlR048H57EtVOG8AoZY/zrt5UkyMKxQb14UMzlw
bECVgOSaqnoBx3IVkFDgssG0LatElsp6hp399Bj0U4Xj/tcJ/NRdEw8LdaGCDGLq
W5pP17DCksC/C0w2l4WD68R38aPUsehyVibPOLAznMYQq32VmzPn53whrJry4REg
daPYDbLy1P09dNmvH89dH/iu0PX5p/Mggx2BojrcvfMfidNkcQnYq7NGG/ajLhaa
MVpgg8oLxHNtVdZfXuk7K6S8WIvf10La8M6S5ViqyCmooxJeWCoSkXbDJPVEAcrI
Mt3ycUL10dVX5wMIvds66ZfHULrmAzyCby4294n7U+l8uViVpDiJ00ASMg8Xvkl6
vADZrSE+8O1IiM1YIshmM6Xk/scQdFdOz3lnrgBbWyjicx7WswOfaOHWr82CiFfw
5BTRGpiYIDfITfefyG8UYk4xdeT32AR+EeFyt0xDN81O/av5Eu502eLUG/t05loY
87uaAXfv7OFncw467KdUu8jm8B27Gz3n0quAF/1wbAe/lpKgTB/XqAggUf+5WDj4
N96z/pSUoj6tFDp0W8XJcA+82SUDR6yFxSR9N9PIZK8cQ8yeToeRSHH3KPQ0OvwX
awq5GqDdEKTMp41BMbSq7bEcLZKRN/P7qxi5xuEmTXBZkozdT9CytumnOO0ANdoS
1qPRQK50Kccr6f0dVAOWtD97JXxuEIm/ZdWWjmhtMgCe8D+/I9togaLdI60KbDJQ
57/3KQ+1PRgsup9wRuwm7OscJ021BNM5AIjPh4o0tSm4W04ClfeNGzDhGSFEjCv5
CIhaDbvs8e9elIb3uIgGzeTBHNhuCF6o1PZvD0cnxZpD79JHyly3lOaRBEG1WniU
atrnvL+hBxxrGL2XBPvGoNtQ1/XewQNLWDZIzZJ63jAu4JSFMWHIF5hU4LrWTNA9
hhYRR55GY9XPA1Dj1Xd7g5kiZlaDlpBJCvYQspDPDKGNBTzG3A5ShNLb042gXO2O
YouWLL6g+aypHkudQ9U0S0lmyy/OVxYKeIM3r7lB8N0jdwv5xIV/rU5RRAvE60cF
Qff5ePxCDZEnRjMAjL37H2KNPm6f2EJVqH9YpLVXzLLexDyrxyvcKRhD405KGuco
G20nioamKh/Cf0jiMscH9K7mz4f3HC62U8208+A0U93xWCTj2PO0QR0Gi4kVnVcW
Gnm5rWUDBh5QEZagJyggu1zOsXE0D9eEGmVFX17LWQuBYJmrL3C6OoThcL1bs+Ml
bQG0pWba3mSwPMVHLDoTiaIN39wPthj79sWr1mBSFEJZCHNyvgxn/48KsewtJdSW
mhOjG2x47lE2xvAste547yEZxHYdnlF79DidBg9G0w7Aev8wbS5vBU3Eg4D6pyUm
ViwR7Rs157OR8bEKfvqbtKEquPLufpnlCAZABs0WZieOKcXR/NIbHuR6tY2F6QxZ
zV3Hn3m7pVastXXmMBzeGJ6PYlBPV2jxVl8KbGSxBVTtiiWwfov25TUOPxQQVdhK
gVTztasdePj7WO1RBJWsoMNL3PgJXWQV+rewhqOkxpJZiyfkDqG2Clj7Prjy3Gz5
D0u6q2I/GaqxDJnAmBphvBiIpFhbo6U+KY03fAvwiZpxCD7l1rCBYpX/80lpR1Vi
fAobFl5c3sGjOL5iACpeUti5i/PvE6ySCnPvUN6a3JMrex9i3vtPA2XHJDPVt70i
TfGPQ7SCj+CuDUWgdhLLPYdzQtOyNpH2irHZLqrUSIf6tFQM/WsFEfXLnCpPjF0k
nNmBVTe5hFWmPwYicO2CQLjEo/1KlLnUN1Fz21zVS8r0458f49N7MQRqmLN2dz1k
edo2yYypVVe8GRCXdBG06EXMSqjMFfVYDfs5R7yL1urJxSS6Belvq0hYAIsbrSIR
kMu5ToRoQsddD4Iq5I4M474vB7np/aLnjJpZSlRxbKGJNX6vl+LGPJLABggkI08R
3IZrvq/OCrFvwNF/WK1EOdbRh9WyUYnHpOEWCELQnqAgalI5XXldmFuji2rv81xD
RhlN5GABYBzLjnHajkTOhNWxwFSgPiw+O0CELjEQRLMXzSA3drQ/17ay0PmQdq1x
T2lv1nRIUIgmr6BuQGfPKuSTXVEEppotzYmBKe5xR7Rw6mzrjkSdAtmbv7b+PvdX
NyrgE4J6nx/p6hAAQUSWGNMzdtq5C99GjubDRgoRcQhzE3VVtSTwcIbg2V+5Lb2I
cxlol8rGRm1c25EwEA7HEo5QmUYKzYo5lJ/H1pCoBBqGbS3iNlefSyRNXSy6wexu
43oHfHHKe2WNqBmg4siNpOJ4NaCJE+KajAkSkBaOBEwSH0w/j/FZ459G5nSiryS/
+HV/XStAFXMyRW9rkBHqb88NAg4K1B/HL2v7OIdvnzL25C2TnIpeAe/60hkqyG+6
ZC+o4zCQA+P7rnXbHyI4tN6tfrwQoG5KcpBlOcrHLmrCbwc9U5jUI2JLCBzXsMoS
FcdRBP85BuDUPRjEdJvP7ovIy66vF8D3uOQtpn44hm/GzyLG0yNW+x+P+yVNjeCr
muMkoG5PEGDM8dmv7hVP3KoLTEJw0LXnEQfjpbd54dOlni6fmUWF9CDyvgFAzWSN
5bWm+KScnjZXJYN5l1XT8krr6tWisDynnPvTY4+DHHul/Rw8b7+y/aux+Wb63Zp2
4k2gJTBuCEqezFTF15vKGwVPgYHaU/4Phiq6dsbAPZdjNf2xrc76xMG4H48vGNaj
MBhGTLYfgpobcNjknXhN+PeNvJu8N/r0GtmBnSkLUEHIo86epro5pXT/nCUfmdpt
7AeJkVOHfqn7ssl21icSJTg14eGVOHYIZGNL3/QaPnaLhExtQpv2ljDsQZGhBQFf
sWX12AqnDjfk6jhju/mQ9y/zXEWiP/rSOqnrFuWH1fNeslQb1/mqLWGrOJYXV7Lh
PReCBme72oa7CZHszpBRLY5qylCbZuLAgWnN3xjYUUl+Qs+ySGub5Y0fdLGl22JM
IgVs0FOrc8thxt0sWNH1pSgckS7UlnKBqC0ejyxhNHmoYrp8tvoAnjJoqT5Q4mvy
yjcyZXxQbiWUyOz5CjtZ76hcNTB+i3jnU0+StFcNXR7fZtE30Sl+4ALvwaNpdAAi
uorM094o3xpHBcWBERc5Mb41OnVux9BpayNoPthFua6I32A8zuw7KH7Xv92hccvT
a6pv6INL1Y1iXmqCKwjVykClEe8X5RBv1JyQ8ISisDWp2zHtxvbNLHHbTLfdICWJ
J/tTiv6KNACB7Q/zufhVTGAkckez4kHeFlprbwSGdOxHIm2Iocu7g6f8Ck34eV9V
V/mWdoBtvfmQqXqTGJHqKmcoWSz1UiipSZ79smr6rWxl53BkK4jwU1xu2JBJdq6l
VDUPrG3JYDFJg8SDLSjhWwy1YcOQLBEOxlv7VMUygrsTVtLS8yY1vpAsf0g2+HaZ
Ym6yQ9vS7UIaZxyEzSRzxWtr462tpt00MeHmemY70PZJBztjeTjNKEtfN3+OEdAE
jH9WrGS9PqGAeoMFYWP1xUPXYuxhR4gK57BnIYtx4REF9iWS5VMB7HRAM/uNJqeu
o5EfDuoEzf9Wcu55hQ39/aS6xRw6SJ1yibf3Dk5l6G0VSm3uXEdWMm4ndjVzMWFh
0yjR5qrjefQegazsxFQjLQG8NTW4piBvozmq//qbGv2ZTF9u+7m1KUh6derQ9O/U
LNXnFAh0RE317fHrCMoULgZpewrt3i7NQ40lMIXF/FsJyRZhUKODjwxyeyGEFbmm
QCv1XVV2Ty/eemAvYI/2ULkcguMxBqmH5rt8lGJyqJU/rNgl5PtdCE/Ab3eiLbsQ
Lqk4Ehf2LBaEs7HAU7Sip7uL1neA8qRaOklgwuIxj9JdV69LTU3Vqlc7iX4s2yxt
t7amLC63Y8VDIJxbBUQQv0u7aoGBnlgO9QaH5K3iojKkGwE7n/CBjsgIY5aDKPIq
eTwdDHN5dKdPSdyDOGRVsx4NyZ4tiemd4ZFsFuJVRTl29pHsH4EvoUjhJ3BvdW5Z
R9aNSYunAWoqmlealZQqiHrzhre8SzxKBUoolAMKpB0mLEIPngFgYX6UCznc8W+e
/ZX9Y3iOZaVs42K6Mulr6u6bYjl6rSsnkg45jsIlfaUmrPVK0b/mI1i2jYxJpAW9
DMGk3/R+OPd0yyRp7sCZYXN5E+21axKwFtL/in8QthWWi8bVmqbdU9sNU3+Z/IG1
kbD6Hg6v9qB74xj0Rej0OhWbIYak2j6zLDpUMibWMaH2MWVHRwNWV8udSmI5zcCU
cfDp/jsMXKI5FbaUoxYRPHUFr0RLGP56R0/uORC07ll3QfAbRBDiDljxZenHTmmI
aHdbGW9RIyJwVz3dTRmEGUmTIq2BXeFw16JbbTvFg14yyObhUeTm/8HRJDWsw/TT
LQ9UN1vYWBwHvY5KXoZ93yjzLv+k8M7RdhoqAIiNgbusc0HXMXGrG68C/CBl4kMV
AtMbdiccWnWwfLvCZX5CgOaXfJVtYmOiD+k/L4Hr+Dsl6tTsCzU+0C4TxvTIV/pk
lmMfkV/A2Pfcf5bttM/Ym07NzQQ+XdGDfYrLJ1uPKDZvx8gClvvobnwXmiqqoUgr
OQG/cZ/4ZLRXNZ7Dge7vTEiRTHw8AQmznM3jBJIaRmeb2YFOt7k3Uf0xCPh+czrc
1iVI7Sx60J72pdEelmql0IFsLHvErlPWyBKrUn7MSjB4vWpSQ4oWwD1xgKenwrdO
mArrrny6HgvnLKRSokA0idqNW7Ib55noqxtYamE/SF++xyvady+T1axDhQ+ysxZV
CozsfXbIkA/8PqjkydZN8FPaVxUKIal6ddEn7m1+Ampw24HQ8wM5RUuORIHtq8HJ
Or0jukSSobynH2gCIhxZ12vOrcKafMadTY7uN0+WDWSEYEJN2dylK4XiHIhobbYW
h9o7YH4n5Uu3IDVAJEJ/dIZ54/O0ebTocBSyaPaYp4owhB/Yfdn/+1mBQ8/NIHU0
rlqXyB9viEIloq711jZWInImFT68pYw8RuoM6h5IqAMRp4AXoFRD2OfyLLn/w8zl
+UveOgmDFAi2Y6GE+RfPngOjD0jv5pKIb8h4/sBeeVjntfhnws8O37IYS99i8BzF
NNHREk4kB9wQ0rtbMRmH+d86Y0V8bsPU6PmDYwpBAOKoMgaaeib7ShQDmlYVQQa1
vprVVUGfLmQGkfKLKwXPPsgvjsZ09oiR7dzErWHPqMjR/Nuj7iMR0OJ6nZVm/QJa
SP3cQRnRfe+gX7ItTJXxcEZX6j4QnNlu3MiVpfi9ysxPeVFdRDO3p1+96EwOpxDV
WjF8m20lFUC8aD1+qkoIqfxzx4ckkvszNaxAWNI9msb7kqAtxPGspk9jULhqAk4X
9Vp9XZWgTTYmrIqcu9EF2guLp6UnP0g/t7/ULMknLQpLDaQW9Gr/Nquz7YsayQP4
1i6/BgnfEYeUgHou29ry4vRufuFsLOfqtdqotUAvZjaLTyVFZrCGpObalmK0LLXn
4dVrYQM6cxrmtx5ETIhUIRj8DwBPQPuKe+NEcT/AKJ64+fTRcBLOTXP3AEhFsoDA
5PDOwaYN614XTRgy3e2vePRIeXbgYB6fOA5+d7+1ByCJfsp/aH/NuzMYVlLEttJn
iOKOpCN+S94eJl4NrPs9kAu3M+fSnmKz12+qeuG4hKIJQMm1uVnv4JRKnVyG368P
Ln5LA9i/sTQRy94OP/+vA1kNlcXro+j9ugQGzU+utHSvKaSHXJaTdP9AkpfI/L78
SKkeSSVUGkhJ4m+WOF59OpuRB2S95nzwvoHNp4LvRJy2bsCiMb2wQUg1MnT+qHc3
plmGg+2V82Q7MnmPsS7Nd9eh1eXBT4dmlHHJqLMIYvxfX28giSqU3LLh2By/yCWi
VVTN9wL7K8KQ4XQB89UmfzXFtVojfD/gJH/LftXYMpNKSBhXeq7PVSZZlBPjVDBu
1ckNl4VYkHyTH+wD/eq0uiegZZbncPmNVhaoLV8y5+WmO0gEfaC2APkaFX+4ECbI
pGKZpueRzhBENMg33/VRkwg07Ytk3T9Tk0FQ3nZZ93Ik45EXueGHN6lYb3SYFXBj
Ihe2IZK8cCg0n8oPXrizeVIZt3UyiSccXLNE5FS6U5CdafB82U9evtOpW4RUMvde
RQAS9Rx8ttArmKYaBkEYAp6CrRxQQNJefQn5SGbbKWYjC5Qa0W90UWeQ8/FjsvBj
V0yeC4vhuDNnkOa79diURsY9GozIwyrqc4ynTFCMoQtU83tdx/ElkEzk/8wOXwwA
FL0E53XWRPj62mPm0AdPsTyRxdK9YJ/qJidSwdMd8tn09qBOGJMDtgVg+QnRezpY
WwcBhGtrAvmqdM7XE+3ig8ElFy4SzkV+8GFzTxBJ6sZr4WeNs7ir8CCMvcmxNYut
stRPeBH82M/sXvHm3BHZwDvukNzFREsfbYc1PAsTHy8hmOWZ56AslPJfJVo+dqLC
t1sLWATlnOIaP953fS8K3kJT4LcDBnlorcjCtHoqgIe1yUOu95wdQ4pyRcd2IGb4
QXFKlPJmnjrI6Ml318gtFHU7I1Wj8gMi//jS2aHfoOCSqi5Y3S7ITUcuuoBIz2Th
gU6TqhzCNZmnVEtDOxUTCJCZt+l//ZLZ7A8sbCexye+K06QZg/+Gc8f5cSTaLKjL
ziG5+BvqK4oR/xLHn+BEtfiiemcFNdZE2wWhzOgA0Bby2z5nwRIh7QWVh6n17tee
chKkLLJt1EFPN5ICFrDKvkca2b6NH+09b1I119kk1ziB7iR4dY0ZyJrfBmWmXjV8
M/48mSfsrmNa0XTL5ocznnIOlfuTM/4j+t1udUZ77cI/alguW9njMyzEVpZrriTf
gp7vBEBGtYs3nDVfO7S1eEiQLzSO/lRVZPCbhmmdzfYYttIC5MQsLVKM/HE6wOQX
8SUpfWPUdY7ng4pr6rrM55XOvQvSIRwmviwDbFgzkeDCEU9irVNPqxVqheaQfofx
AwMirICrMAyiCFUypqMfnEOQiFYEJVQd9IDd+rZtgBake76LSc5Wx18WUIuvftPI
nGVpEO3oMvmh9/mg3rXPz0ZWh47loF74NraV4CewCEfPbOvwZm8AGSaqGz6Dn6DM
Gs68kCysb0LD/VL5TcNCzR1bGLHA9cNFYCXZ2RlZbaOGjPoL1X0Cn7m/LHXDYveP
8EgbuFgZcP+vLMw2WcabunCxbegFYUPofesHrmQgcD1orWGEZQr0MTPI6rSAG/u2
b4B2cDHFnO6QlUu4Gx4zQqB10vJsXiMrkvqipzP5YXcd2v/+GFLcv8V0RtyUHU4o
UpFwyqlVfwyD8bSDzgzZAZLm20fN6fwwJqmb4HSdxaWlAvpfzep36dHn73ARn0Vu
QNwzqEx/hYJy9dWQDMzxy/Y4Dh34iAqDxM50CAhT1tKNSV/AwKWrINDLlw2/xSwE
VJ/TYOKyqJiUC04kLkdOa/90fAHDihpGOtaWRBYlTrhQY5qxGMihtvr51kvc1B6R
NW55LM8gkyxIBEjfCUVMhtsYV9bmnC1akiqxjSYMZL/CvirqEnZQ59okrQBCPgpH
jJYFoiyxsfQoJxZHqwZjCzY7ffny9WI3y72EfgNZrbkp6s2wjUsB2UapIJ31X67G
Gynu6wqlA8zb6lXCslsdvVF0gXHdEbJ+3LDC+nuv1OPIdi4aSJ2MvUkUk1l/FFkz
AEmz4CEKcz1Lzb6fqnNtaGXgLv4gqtkRZD4QGNv5NlD3kZDKau4rgwOfOj5087Wg
3D7waAz50aRX3zuUdktCNJwrMDEd5L713YDcBQbqn+G716njE4EmtyqUX0DTd/wG
3xjByMg5qzUmSTsaAUfCmFilZfU1XlSAlcnMAnpnVAq8giJPT2URhsRo01KSDbaA
VvDiUC3xvR50Epd82Iw0RJxhTnqNHekK74yshLfZucAR00hq1+3wgXdMVBS6ySST
xu/AfgRYU870Sp2igmJtysuyRh6WkCPRaarZQPZx0RDcXqRwatZUFl/0KDtVUKDQ
CCsUK/3iyZn3eTlKSTSxGaBpaXkimzz+lEprFFTqmpNtYMcPJIdeGXOJbHfW9EGs
OOi08DTnFTCb9eMwvX19qxdRTYSx3fNzu4RtNUjJuE5LAfOGgex+g3OB+JarSz6t
1vI8IjUspRwqJmElFXbxwDN3buDTzhD56ADnYJKvwtjDk2yu/pOKOcLaJAzfvAhW
VXC5GFkXQEYh7lMlIJlpi4ngzEqME74SgSgFuvP9fIerWmTUyl2XGf2E75jZWJyn
uqO6sss01smkB4V+nu9oFUJ3KxN3qSttMf6BVwlvgjlghkZXUo4Y0be6m48sjmUT
rW+NenE4vjVyE8IYbfNlmFe/47d95Z7uKeMR5vBhZE0pGU9mZWS3O5p6+jZoL9z7
KH25KgHAXnmW2KieS3VvZ/jZ4GOb0FOPkVKyPyOXmlmV5TI7veE7JlbZ3indxR4q
FLYevKJ4lTeMnRTdFaJK4FWPMrkQX8wq01et30DhNd7iPMmPS+cx0CxK8PU2RqAP
HgpEy2KYTWRdD/4bqMqVXJVHcLpLEtOjun8SSVrnx+n0FDN4cwUrXz9IpeOnu0ie
xyEwOlYJRKRZfYWBnExykUXsUJy8gpMwMaFC7/u8WdeimgC/OZCUOKG5Ijwk4Rpl
ME9Gs29XZTucpACP6MgSIurUWtSvq9PcP3ci+fK8q1AQtH8qlPUFfK2vXeNHqbCP
FXQtOYjqjCwZUOgWioYCKggn+0VfSbvmBMNI0uZno3vPq+FQV0mZ1q/a6HJqIOQb
W5BqxCMbRl8chkruuYhJmtngHmjbVwW49MMxIv1FZUUD/2KT9l90pSl+JSqmoAlK
H97fZ+apkwYBdk5GxkbVXtjynorw/XKcVWZvf9qjm1MAgfFnM835adZFYxjT8uxe
KcIe90eJfpKPgg5AGET6aDgnyN1foyRijjoveYc6uT2b/RLYzdOYcFytJ9f8S4+h
mmslSGKuVB8iJHb2q4Wd6X4ju/mAGA/Ke9e8yzkq9IuAjOx7Y/AqPC+MbK47osLl
shlpG8O01KuI/AcUrXWkSgPRSI+1wRyEuetTFpMsWMxMgf4BYpqiKncrJOSXd7T2
zg5ncuIRDpY/JO1dTNfMBqQoMeAmm43/gpvRsiabVEvdmGTLSK0uwk53yHoJ5TlF
WQRCRd8uCu47ozaluDAMznq+PXYh2proKrCsFrAS4TPILWQpu6JWgsZ/pajflWE/
2rtjPjs42gxhMCz/FpwNRGqExtQsOG/HwqBhjBuMdjgvSqn61KIVSehlWelGYgHb
mXP2QzG2TsUxDLaO7TdAn29kwYaQBCGeyPeaJu0WeBca7YWfgQ9V58o2wDBAem+A
EOa+NVkdm9qmADaR6n+HzC5IJLXBlhl/apmS2u1uvLmeS+cMmfcaGG94/urN+LiP
NXO5gJb47jae5JMRSyyNYOC9R1Xnwd/5jX5kcbMzW8yyktvXqBZN9qVa/yj4uodL
ufWv5f9al3St9eqz+V7OGSmkPtaP7N5jr6UtuS5Q+FbdUiSkspK97V8c2UAjBN/g
zqm5nTaNuV8LmeyyPCcdf3e2QhUs8pnnhwJeElf0SNlEB+/aAOQBYCpQ7tsdeL99
QgeFh4NAZhkRY7xVCc4H3TIZ5Tgpaos8agUwyceWEiPjb0b1QaTF+TAyoQqRHIzs
p1gqKBbNdNJhP9Avl+NWZ83+izx9v9x/M6/fnhn81CIGvyikIHluYq+5ImUBGFX3
Nnc6hfruX6AgNZcv8TqvZwZiWDQgjICFl+3UUgxf1qH/A1W5V/91lEGigX/WDamZ
R4UgiKGn0YV5TimzW5ErL+5qj5vrOZvYobKlzUIrbHzVy4EfBQdE4BUm7T62X69K
Ub7u5dMamURkkDIFf4efyMNa6jjEu/HgSyQNxklw4N6IVjm3JOtMBSal8+G+hq4J
u7e/21byLs00Bt91A60oebSvcX0uCBmgsiql58FWUmToL75meZA8iNcnbNY+K372
kNmT/DavxtFIAcxfFiJe0SPWm3WXqdRjXAkB4tlL8s2ubRPKRF52gYSxlM/Fr26C
JcNGuse533WUEBxWJOedr+0O+G0uYi3WuPEYV3UZ+H6ViZeqOLWWrX4QeQ3IFX1B
wU1Q7hA1bsV7cET/HezCVCBckysJ1UKkqy4/0y33pu90yb579+HScH2kikpC9t4t
lFu0+jcndrwJBzsTYl0Er6adPI4hwVSCuvEJeyk5iVrurZ2k3j1wSM03Xz5lFz/d
msvrrxm4x6b8rK7WBX3jm//HI3OhJdw92Q0G5n1B3k81tjpsOl7lT+PyTJw/9vG/
RJhj/YR/K4kHwfziIyN+uhu9GJe0lJkuZd62YkaDoZWc0tu+bqKBP0wtdRXJCWKE
g9qTAN5H2a4lsYk7Enyf4+vuD4Szf7eX2KVcmg6C5N33knDpV9g5+sFXQDeRt4++
PRp/U8//K6NPy8bzukKl3qgdISsYUX70Emv6tNOZOYy7Nal89FIvCJMsaFrDNh+y
o+8TnWCn0V4+crJJV5k0kSnrFPgz7IJ1O8lxT36tzpBJ9fJsarefGrkME+K2YzsS
X6Bi5Hutypt225zzZlDpvgtd14hITNl6uhqeyHL03SdubcR7bx0Xq6CqOzFshJ6a
XqAHFA0bYKnhHcGEdkq6i9nRAw8gn3OmPnBovlilE7fOcy8nq606kSAcF+6SPM7K
VBHruCWBr3loLx9DH66VfFkLzH+gcbP0J4mSeWE1kU2TLPaDfk/0n737JIgbfGz9
XFFoSXUVRu/raBR9icSzJ0/u6SJP3Tbt8lqGdYg+lyUk63Bvi6aTTQQwSs1IKwgY
pxjeaz5slA76Df0KwjEYFFo3pSglFHhYfrniER63gBvXUHaJq1jrMVjywxLGw4BJ
CBE83XVeJjeAPncDJ/kWpyklfr7qdquaMsCQFkz9PlMJmKdfQSXIoKRbdFm/CuKz
GnmyxrKkkfwhyW0vdrY1zjxhdBqxMD+MDd+nVJa0x6CKXR6shGPzLpdPY+RTXSyP
cE9hSj5QQE6sELe/gVcKflJO/QbuAQCzfIibIKOzWHZTskhN+yHHcR9zrBC1NxyX
94GfvBbb7vRkW/7LQgUd0kUUYXmnQJNJ6fTNk6eu3WEOckXnvqE45hh5Hw+xqVpA
k4+E90Q5qkzWNyWLYTqKJqq9b7DhKrL7Dp/4nDjZlUqE4urOqJejiXvTxNU7ctn6
2mD2idfUnoP9oHiRZIZuvKg/yD6xJxZRokedD9EwMMT1u0XnDchXXnKRdzMOXwO3
K/RSm290M9NCcA7fi8B4W9Tyy/uNCnEKPvI41ReS9o6J9DOOwWGty52ErDQT2kcY
uwwqyd68QZz7pzWrWlfgU/CGe0IYIgXOa5TmWvt0A0GTcFpN4CBw9MhcHyrKghA2
yyMr6p4J1tesosOfEeTjqVZyXjhcq0f/cYBD+NRc0cq1AYIFOBXtW7TTg53pcti1
g9u79vXYthvTfMmFLe3w1l7BZ380WOfNGU4ffSPYZvDLqKWNpmRxcXxE8+D7+n5g
iklJxOJ7/Pc6eXmZciBnFTVvKwqKUarPV7QuHBmTi4BVmzuX8iCBwxDtImsfLYTk
nwVWxq9eo9gyVJsKJ8ru4Uwk+y4cQf6RsBFDpzWEfJKYmaTpt6WpYp9fLdhHj2N4
jfvOSrPvvYSaJy8AjHhYf35/sTIUcC74nouELwtz7T9bitKJfy3WtnZ1fHeOjRDa
UkhmCUYy9qGr/n7QT+tcG0Tn5u7qwGhG6M2DQefdhdRRCkCj2yRyeldM0nkO+HA4
xOOUiSPLEtKVfC5aKNcLMgVrWPezi61SWn4v7lykekt+nROTG1vnm00zuXmfaCQL
BdARF6304y0zja1hvc2fXZhVdCyl3aRu5zris9UU58jFhoaRGG0CNlPcDfTGrwNA
qL4mGPcrvUXAPprYy2Tz+AZqt8AoENi7r1wpBrNIMO8izEr7NNIGY6Ocwj6OKzQb
ciexF/RuzS7ev0ESRWXvm4dSZBnQFE4XcjPU2fguNlRi43rOx/XhavIgxF8/FWf4
/qmLpFJ2I7KhwXU8RI8X45jjJqJ9U2kf17Qo9sdz0Px/6BXHA4IRo7oerRLmuOdL
SpFeZI1zaOfPw4MCo6zDbzPFGVPjBW3cbPz67vJRno1XxyqT6aTvAFBnXvoN0ius
L0BZxHeSmUmJj1PVp+eGDlU1Qpyi3K10v98pw+KmX/nhmCcU8rWqGJ4CG3VbTckT
yGEyViXkife4d6EVJdts+FBGq0/WMS2ah4humYjYGfahmqPI696LaXSMDqV0xlOa
pfq4KuFyfXM8l77aHNuE/FT8muX8e10xHSMdBM5IA1S/gL7FWZ/yylV4xx3+U3f2
wDs6SbPLjAYMuVZa+f5R9ITUqwbwTlbaPfgHNLxv/7oz5uDjWX44pvDxn7PJtN6B
vtrl2srn9JiVyCtRIzp8QNiUNTHTIWVfYT1EUD0Nf8xqhZKmTInoldhgoE0uhoRU
hHcZq55iAAD+2BASvTMKvnVOLSHi+m4IAW+AwT7M0vorlkp6X23yAobQ9Uy+MbgB
ARkxj6yLzXkag5OR2/bYIOYYiRpTAaDlw4DBq3otHWDhITkRd53b3f5G+PYkJB22
wqRjSw+Yzxd3WKuwKY8kauRN+aktt30alneZaxtaOB3lLlbsjSN0Rx9aeNo7LcWb
hDoKLSDZjjmwPGhQIlAaYa+/Jg8YmTmg4DXk2PjE6Idoo2zcT2xYtm6rFscDGzy/
NFm/1963YdVqfv1mIahzxHRkQqSv2zIyNbNEdadoYF1JfHkzeCdIIhVyf+9QR/XD
G8iiWjQeG5njKzcoPQxvcNmB4KsGfGNyJDV1ImimvkRoru/xac7zC/hz0+JfoX62
lNrDnjCj4H+WXzHAobj9ZEJkFI30OQ8RusTSS7BgOF79kxdngkmI4nhkQhV46tPx
4S033QUaS7+bN/emWgDC9mfV9YS8pmeGrT5U5TbnAIJuZP4TykhgjiQWQTrvEwq4
C2w96/cicaC0NqLc46xZkynWs805X4CfhjLyNx/QLWHnTAqvp1LyipW2k1Qo1HQy
D7Z0DOOo2GBaNrJr9fF0ZYsMFpXaCJH9q567bKLNeORbx0gqkH8O7UagW3Th7vaN
B+L3A9Jc4/TP/rbpMppkYu7HE1xALqWVJ7CN/qZLvHWvAMWgsoKe/3bpK2MY9iqg
0rpg6xsm4gn9DGpIq7ySpMW33z9FS2Cwk0MO3DUNgOQG9ohOwEqtnKdSY5uaoABi
XCpqe/4mFBusKqN7iZn9U4LR2USMY0uijMUEYg9+GdY2OTWLn3GJllEbQgASYG2Y
K9X4olcg9gQWSIXdLu+R2pzTrgPZ3G6//8xL9F/dK5nRU/jxInxrqEE7KbHhYYNE
bnrPFBKxDCyWdVy9aVZFCcLgKNwnvClbjZvnffiAgrBORvcT6E5nk/Vh4k4V9Wh7
RV/oBiqBZj0X+iySSpqyJmvqBhYnACLwTV1iQF6HcEYxAZrG/eHkcEYbJVkgaHtX
kvcExZSdfYRYrlpspYB2vE/Zs2Nl++wLStEr0Y5cZHzyRV6g4nvpSA8fX84tAETB
SMN1O64MZg1GBviQF2Pcez5WFTg+meHWYRqU6H6aoT6SZsedISsmaeMMd2U9Ptzr
ev1VgkheEXd3uWr0enbvlRt5uL1LUKYhg/7PWj+OK7ljAnGAWgwzfAuWJr7xsyfC
+OvkwBjKPLfmz/pjq9IXtrXadoUgP/8Bs3IV1SRHqRh2ikJCFC5YlZdZawNsL6I6
4+3Kjv5ZMFnS25M64eHnzjVOzjssP6vCBSMCArAZYACaBu4Vq3NTVdjPwQCVGrZT
UZmU7OTxB9HZllgAS4K5qU34dSpw9b4VPOQVztYB6fOrHjp27rGYJ36qfdRXxs99
LwQChK6fPHsNmJEQi8b2pt3FQ3ogo1hokN2iLBMr6nga8eRiXvao3ZPLS9axIB/r
rUS+7GVhVDYtwXvuYpbphE+qJxagZoTlvqaoq/Ae2cC4/+rTbEFPcat/13EwpgFs
qmm5NQcjCxVR7QDXt+ZbwJCD3N9+rWfUhWoDowXTn2l8Ub9Zer7VWrnYjdK+jCc6
3jQNiFQ1JN+838F/VtuSRbqBxPEPEPTURp8/TsQav2YGfXjaCIPDRvCEhURJyWkD
JsbcEFSeXaoCWjEcJM/6NeztgZDK7v4hl5HJIHSgJAs2aV88fkKAM+/QtKK+mAV/
MXCfG+Pf5/K4Hqct8zN+KQR7oLDeThDEwuSHCrh1hTeL86IAJx8Zxc/2Kinty34l
VRrFyjnOX1CQI5n3e0A0dbYqRji7bJl2tyB11eJLVXuDqOmDlw1l6puHqKpOUWmA
/Uk/C0rsIdHjUTebR6M4UcRCg5DzuvAMcrQlpdbl5tA2gBPNdjCOStfJi5J08evS
qx4HD2rzbaYtOvQvDiKSYNqd8gnhhdqozqDXYMrY1+IcOdvAqnGFv7U0cGxkuf/8
t/LOYf+ap8zw02iKgrBEjCnkn2WlVk7DQa6rI5c17+VIV5h52IB8os/BPyAxaDeX
4cWeB9NcyFbRQiJ7UcN2kMljpAz8c+0oqOoyH0FMmgCoa3hkJpS3sdvuORf3LlyV
ANz7SWQDFdPqDxawN+JFRYJiqfVSip9gY2kKCLG04T6NQeSLxNkc4jQfqG73wwkU
Vky7VtaCBOnJ2alqYTivouaHZLWIaeemjAu9TiX7amqBUrzkITbfRc1wvcq6lhtn
oabVP0nA6E3NkZuRxy7wbnePeRQRF5on2bNnQhfiOvkuc4dh3160ypvlj8gX6/UT
32Dchs+gNOqlrzD/dpnAFURvXTxSUK1WpsBr9683NiFRUM1sozjNb8GSz19dL37Z
a+gMcep5g+mxs85VNJm+VuKK3lkElhsN7kLwnq5jsfSVi8s65A09eajxyOHmWc00
vP2dB6IssJPWth+5uKO5KbZdBee7C6CmLKyotwsJDaIBn45y5JSvVMxIoUcP1kmV
WqugnGGyo01/PVfZN5wHIHZKrwhFgdI0DW5XzrrzebCEoUNE5K2esG+fcxPiPE6o
gUoqa8cvJjkcP3Tx9fb/6im5IXhMeP5JNL3YZZFB0X6g5s4BCATssPWNKJx95qfv
IdF2BryNwmo98eLnDnmcVnBRSW5dMVcvw4Zazvrrtl7hECVL87oM92yFbD0qRVGm
+c0COTr4XcBclEa7fRblteCgJzs7+ch93zxdjr2YYjT81dVQXZ0w3YFtwSMLZjjO
rOU7J2XwaIGOAjz9lyQ0vHMvFYiHRupQDzav2fz58m/zO8wbkM7Qh1o0yFnIasUu
I6P3ugsU/78IPCCFgLQQciMH/ocSAoGpFkQDHS62kFtZdu7HdYhGcRZ1a6VO1FXJ
5x1FhH0pJf68cIG10vD76cDe/GIkmp5eY8tYKXS2aQmAsTOfLKdVIx6xWYmzM24+
Sd7rgmhaAqCdcM5m2pYxMFpKNA9O/GPnwSKqm4k9UNbcm4zzRFcpt5O1rUF+1hjV
Cl9xzTIBX5bGB/DpHHXfkBjW018zC8cFmOHyTyKtnTh+CKk5tJZrNRvir8upLpBa
2KunTIqrpKpgPxSMkmh1SEvS0UyEZFiSFZRAbfETripAIzOG6E6SwfMwvz5SjqMC
R6CS9DGSp3gROlXO7MRjPZS+sNDDXXvnRWmIipg54Lo0FEZZhBjmzsH8NemcElLk
eKPT8jI7QKMYTCUqH8/6xpa0Un769eT0Pdct/NSDg2ZwkcMtSw4KgggwNKKqg2l9
TJbE0cGOVR6jc6MMKZ/Y9+qtrYTGFXIS1Kkow7rtKbA1AxnDTQuwLBNla+SnVSrE
aPk1q6CA3d8uZjvCqb4IBc1NP8k4wP4U/wHvu/dsC9XCkqxIkqjylqzlU0+eL8/Y
TAK7pV+DVXJI20Jg8YsTu4OgywNj2ziueKT67478CHzAJS+q+1G9tu371R/CvU/x
+BfbfXOQKkFxoFRC48f1kusGK3S5MtxzrPRU5FlxnvWyTiwDbiapTDHiuVuL5+1C
lF3f9qK2VbK2Kb2Rv9IpW/zLDi+JsNlwxof9DTml0xqPY2YHqMMx3w3+oO2OdRap
GkKW0hN9bQ9pJ4HxWT0CgVtZe32i9Bq8kONu2y8StEu11nVydhUDCMOB0gWzWwZA
3ocEvCeFZhxNhRwHxZ3F2y9QIyehcpckOW/cTQsNPv01oma5ghJP9tsv7OtQmq4e
k+kKMGTeOmB2tWwZPpjpR7DYtX6s4I3Y0ENxpmfyW4j59cDlWvN4qnaj5PYNqw1E
Dgcoh2Cvfhf0dad/Q9TFQhlSUdCIKRjE4IeolGltuKgnPoCq+M0rGRLzdG6pnEA6
y0TBM3hpv3mNugwnuD+ZoMs6zsfyd0V5weUHMXEYGJPKNrJ3bPohpvcwbv+zoJGq
0LIYf6yjgwMzpF9g9NdA6eUEAVO6/5k8NWxf548KUvT/FO6UV51X04BNEJ8LmP7G
f6Y968ZagwyrGEIokCW54A5KBYkwM16R04hkQMveJtl2nYYLppwgfalR/0ewS7fo
3Q9Mg5AdRnhd7GeAxxwNMwn8ahx67WJL9FKSkIGiWA1lp8WMQ4JVJ55W/VLf4dnH
QQ8tDBUDXRPM+owHGPe7nT7nSduZOVR9BkvkfxoLx9YQaNu6+gmbk14v4LsJ77kB
5nvQEjdRz8GbAV5OU3IQD3ficfKOid8P8pWQXKKteoG1z4/ZAvQ6ce4zN+HDkHON
4xXUdvzRYw1yJAAWXa86L6tm6i9vjTOQoxLSvFoPFMZAkbA1XbY4M308QuIWFGqu
ZnMzlFp7+V/CQYG2f5PqmiF9SEkqkRJ5eDvVkkkhLQaN2sNsYGUNP+yQYSCGhOjC
YEK4sWNqHBt6MYDPV0bJ4T///5vsPgWdPnrLITkm6nLS/r3O9PEVowlGD67DK+/b
NgKz+aj5+ecUDkFwVdjVIoEJ0c+THjjr1a2kXAnrSy5h/JztXnDDVp6UobAOUs0W
J22ldaMp2jv7LB8DCBWwyb4+qkc4ns5J5rYkbBYgTc0CM1IrNTEcIwnIDx+pTJh8
O7Qrj0xgtdilPaR6KrC93vRUdko3itXkwls4PBJuiWTGfxDUX4hTg+I4hXWu683D
8Cn4aIG85I3CrjQNzXK/T4s20I7Eb4Uvxy26vjqnrvbdsPJKOSu8tVBt6mEDkGz3
tncbuDRIM5dyZKY+R+8uTvHM8qawfifKvJ/2OzRzKn/QupLbw9uSD3HOP0wECiek
ArBnDVXU0fNKee6/Oqg4NDvrb9d5PyadMwbKHCiD+SUpxFHASRStb3ycncx6yA/w
aGMCBBhygqClGxJvDHoZvpCjK0aU92kdgDpVSgDFF51jgwxLz4ByO53ueOP78ZL+
2bZlJfgmjV4BerUb7SlmDz/M9Hrrzg4BggeNGYIPQpTBItF87EncJ8JI24siflt1
Cq1nGaWeSN4IQ6kEqEajTqSWOoOxJUjyGRB0786FV+BKzOVbii2FI8UinH75EQRF
bybZV0ThZwN/tw2ryN9yojVUAk65i12xCX9aaJ4jgA+370ubFdQC9EkNpmGpPbbx
O0xJqarAzznQu0vS2/+tgYI8g96geyY3879cpVJP3JUkKX00PQRs5w4PmGTIhJTP
g4ctcBF96LKFn6JzcqEvTk/8ejzAiCMDqt9UzAh8Mh2/i8B68VixTCNLgY0i2csv
ON744H7XVhuk9I2yPNIzNYp7s7E1bPMXhB5aMR9Tqjw8p8KkxadAuA2f9L8tFo+A
B/W8PenQ/p0E1kVN8BTbdASrg00mSpMwYZcMJ4+GtwwMHXti5gHHRFbCvP3HQYA6
/VyX9xe8YYObsihOTYo2eCKt72V83gKzixdBC+XyAsAVT4SK3/PT7VKToQrj4u9O
7IqYGhBEV9AljG2w0YueLvfc61rvbE0VYQzaPlWzCefuZ4ysWE2N9S42KJd9H8Lw
qdBAFtPh7O/CHkppLiTf6GKxafAIfeMzJXmBMxAKuccutkkrER8LZ4izuRPKhlKk
P+oioSkbrwk6xMomFg/+sNftkm/bA2fEG4PepdQWDQ1boQ86V7U2nBKwnMzu93ze
8FweRrtnMvHyIE2iXCF40bxCRCf7CiNrdROjV2jATQS1QTz5s3OBIznR6jf0M3gM
Q9toMKX/bKToYy7bEiBXHywV0fCcgMP/Ry3UAGpaAW3HRPMyY3K5+LnJv1uvCIoJ
SmXrN1hyE80BII3A6fG5JUSOeVxkuFRSWXffLdtKbRNnRwSfWNILF5aIBYUdZG4q
OlxXQlW0uXSevWAHL3mNxjKvnjm7GgYunyHgzQgax+uuH4TIWVL3BAitusiFCRpQ
bZXRlKa7HwncvbZCOIa4SqTb5JHf7uwS2JNPPxE9gmIGLjBBUqiuMG3TDSxJDrGJ
Ugsxoe7j+tZXJy3jBzITtnBo63g9PbNAFKC6OA15nHtWVwDWbH7kWBCLI7+8HxYb
U+1xuZxsR9SejVpmALBCP5UF4rqIbO1uSZi7HIt8jWrbuoV0vYFs+uDLeKpa5Yd/
2MAZUPT1v1akoapX1HgPbVjwaLF5GNaMnDcLUA7hsK6BnG3VpTKlAwCqT1M82O1b
moFy5DWMmML3wIM3GkxSW0LJnjMJHfU3BW/MaUfRARerKV/R3ExtlepSLQeX9qG5
fYPFPmaH7aP5CPb6aPj8zSpzbiyNC+QAhDGJ5D6DS+UWMzQ2RfmLb3wYEI3peXJX
JrW1BY4RjRmW7rWnJMt8jDaq7xBEFufdSXW3jePu63EHq0gqbs3wbaGy6cITWGwd
mIZ7H2hugRdHGfFuEAj1Y72i1499OabD0CJm3YCluwmeVFgJKTm1TRdiHlQmUNRH
/jCr7zsuvEb9SLM0zqQ76twaK3KL5NC+QN87WPwHn5xOh47hvnK2MNqS3NVCZ7HV
3GlNpCt9Rx28bnY97XKKdqvqZP5dTpD6QXJ0HjVMKw8CbmVffhC7Vd6YJ/SeePDq
L0q9k81SlgGLNvLj4aMBCRbu4ALenQJ5hnNfxNWx1hgRrHQS+Uc4ciny9oMKKphq
VDEmUpfUMJcGJrXAIW84EPkuPziqewyUAxNBMTQSpRp4cB7IZrhiNCSTCNsbQHHK
kZCAj3Nct5/jQCtWF1UU72dU+0rA/T7wIgt4G3y7lUHCXfFe1GbPl9O5VC7faf84
O54X2zppq9prhDLQamiHWiyCCdBA48LA6c+/YiPzx1WcvVUQJpcdutt+EESWxDf1
7uPRPAk8XkWkO6u90rODyTA6sg+CmI3R/7bMeUfqs8v1cjfX3pJThr7h8KrgdERh
60K/aCUctLe1fFMF3AbqIrXjulkeUMo4Ny2P63+F0OFjPPH99DGxc5VMkccM3s5B
LfFXl+DyrTpcc9kCUONqP3baSL3gC+y/OOQpHwjNO3kt8VOnv9pXejiBXLeW+KOS
GcYVVyT/JXWQYWE6zlVz08HRFh0IHT2MHlK2Zdroj0NuQnREvl6cgifMwODZWA5l
kP1VoE0U/mDgDaCf6nfeIeOZ1ubV5/IuEccHlM8EduEftdZSsGMfxIQJ+rUJhHIk
hovhUoZGILubNly7UGX2YSFTaNov0xy+1OBucUqx32MqdM6fwNdNVyRPFCpO5MsR
FdvRU0fQOePLO7rAenI3HAESxam3QuXUIKhYq58WFuTWEykPfpXr22C7jvZb9LmW
zMc1Ofvbhf4HuLaAY74fR6GztwdlrohanvnjdTWIe4kdKXvL0S9ikexWyuyiG9td
yhMIEk2nnTLRJAcHoXzDbyj7Iaae/BWkEVQnwcrIvo2E6b61cGkZYIxWaC96GNk/
pxk14s6DWx6pW4icaeG7+dlZX5qU4qsMq5Vvt6obiqCT+WyNQnyfqTFliAmUmAaC
8iZmjAby+lZvh99HQLNd5ionlxI2sj7XzAVbB20XO8ghUMzU/3a4Xd40CvGlsIvX
nGemDsBTpJMKieFyvwYDHzSCLCfwCeQfznLcqA/XhHkxaQsUUTbLGQLCMhBmdvC4
5zsRJgfCMpMZO7zouDug6+x9IB6ddFZP3Rv2jwLg/dqw2D4FB6pERAWvUHyWKvry
GhUXZgtOXEZ6fujRXvw2Mzo7djvh80jy7pYZAgy5OawvO4+/BLr1+gzZhl412U6/
3wQ2VrPH3FqrLBJoXGRKjNAUpYl4JgSaCrQof5E1h+dLb3W29bhje1wKe+fFOvag
B5cmVZ5xSlFta1r1hFHUxV6HD5F/uxeWq6vQm3Ja3cG1gkj3qn6RIDAYw1LwXQEP
3H6YIlRgLiAVsjIsg2TtxHNFMwa7jykjvmecJzPf0ZnBXkS7j7IQAXBzkPtaJMEs
brhWT5MlM/TnRJYnk3saJPlVCk1DvdWN2+GJvpS4hJhJQ9sxaGf+Zyc46QzspkVY
ddq1SV28M92qi6TXs1LNbIcBknINGEli024gr7RkR5rp7wujOaQ28ovRshBjGx/v
gqu/nA06x/HIt09qTTuE15v/JVTowVHa8TWyio0ItPsLHL+wNoqMSWTKOXOYwDiB
/93n0q+0plg9Mmbx6P9/aWG/P7UCUPtGjrelyrrT4WiDsL27Yah50wjfvOB7UBpY
rQILfQZqcIL3hzlzqiwwi8ofhL6MRqnTfUTj6HdtjtjcH2q0vk+XemJN+MFlnlfo
fFciLk41JBkkBwHjZ6pNHH3pnMVOu3oNDRhM8rSb5sWJghcaRC4kezSkkL7HPRuj
vTw3yEddD1G8yQA+P9qKCGfWpCVCT9ys9nsfatTpjITbk/UmeeqGBMYjtQtLOqEk
CDfsCdhZEBodH7DDq8yg3UKSo6Ums/Bfcq0zHcvqD5ykWXFCveSCzemmXmg4fYJc
MsO+k4ZIO5ui/99zuQ7gnogTaywabwjuwSIZx0qKf0EXEhxajZIokW+mEzoJj7ba
J6hqghmuhKiUzhfJQfjtgryca086Ixm4y5ExFIIUBW4iGenrXSlkVdcalKEEb2Q+
rwalBNVHuuS00INVK4QZ6VzdUTzvIF3gAhUG6PS8EEfApn5Ir8wNWgWLfCVEPOeg
hLnyInvtND0+o0osyCeSV3qDYaTmYYf5u/g1XO0gj5zxZa2U3cF/7NC4/xNCYRX9
HuUwTYKhfvh/xD1KhKOr3UGssfmq7S90p1cV2xwBXAFkbNsohSFnk4vDsPIuVomN
GoBnEAY4dP8bumr1LnSj+Lp75cDRlQQZlsbPrj5opQraohEpXahom54VdfqXxK8W
xVq8zvVJippWpitNgVuBJd34Kkft44zHUA4UjnnrAhB4ZEumKFaZvoYXVo9XktUA
li8RkMuwoMEpzC6UIysyxs29847UoZ6Piyvheiu7rfja5lDrT4eFHjigkSXfDgBm
JQiPkCIPq++KovxfyWH9uL37ab7mKiS2zGrFKcZl2L3yYnFJUQYYpdZJ8nWq44nl
RoQA0kz417EMpAnImHb2RiMkxlpbxK3aplV84Hrvpa3gA+g1SJmQFt/GimDAIPMw
cgPX8Os3MQ2on1WLU5rPWGSYH136iLm4xz9W4JmxpnGZ3vDyVKNxgTpRQ0u0eg3b
kQ+bpd+6qI+6rLp86V1T+rnrWERGSCgMEAM/ggYuyZFR4eWwJJx1gjuEyDSQf/Os
i2R9NlsiJTbU2o2VnvzmTzr6yuyhWDL+zh1s8FfJHsi2OC3SvhRrgZS+DbJfsapZ
C7cky3Fqubkfq3gt/HBQHwVwM2ZxRmcPU+nOqt4LhW+sKA+P4ZFZgW/ONh7sQyQE
Boiof4ENe/F2Ma6dTIL8Zv0Lys34QQ2er88NS8PbqFV5nMh6dZRbXCRSWJFCLFGF
xrwyzvvA3NAVXKM3Hv06fJi6ZxQEBnpG0/KbgKr3lOUIh2mLxdtSeiRDgvDZTLLv
/4c7pc5BxcOtNKDPOkgvchDj3p0+iTIXp5vCuPPlnZ6VWt/Op2Z5uHWTFOgpMfQv
Rr+2gnsyZQpN4FTAkfDNekzPTqd/avdf5h9TNluKmBjwLyFcgBD+b+/BVB9h6Vkg
0VGf9293THZJq7q1CPyOq5lwfi382SXoK/0EhYRgBNLSRUPq1XMvBmAQjUgjj/1v
eSWiUEPy3aT057xzCK2mFm3+TqlwrVcb6yLqp66/nsYl3ANRKcViXUPE8GqrE9WE
rWQ/fyHVryQUAiMs6C/bhsFL/IOrtOdV8sovH1hQ0ZHL4B7SslJdeKKY9McrBmZQ
1vSPLHE+ONidZ+S8BFZZITmOHIKYMmOT0t1rhcCXK5uW5kGa0Ot1/pMjpD0aN5Pd
nqjpZt3mmj5w2q4o81kbY48qyqlwHIlDSX/BsVQraOaackuj2I3h6OmZX7NVzao3
UGGiJ+UNHBsNEYYnpTYUnooCO/Ol4vbAFMHYpWwgdQxwSX5wJuUbSeVFcJ6KF2Ng
G7J1KekMwyqSuZV2qrNRFZSMJDVJkHmoQju/+d3BzuTvQ1mU23aOVFH+rB7qAnnj
jRUvdnQny3TETsf4c7dEsBD2Z+yS1HTGrpRSosMjAkoBL/1XybvVsmIuInaSEMuG
4NePwBbx3KIYgthyjIsPkAnjpZ423WRYBo/B4uvlJPbJzbDRNz5yyxzhOVMAiHmr
9LjHptfJb3diL39m8Vk+LVbwy3oJ2I/ZZCYvthgXIZPitMQMWIJne0JnhavVttMp
do402ejiFgX/Kq3QaSaBSKwX2fKRxJ6txZCYnDHnBlBhAPgAGuoKKGgKrvPWCQp6
xI3nN50em3n78qoEHu70TEjVaieLGM8BOwyLtURkbubQSRiMpxHSg+7hnO2UPD7u
VM0rCGtcHxaCZCJzDWdMPjwgkzV4AfLgWnJzQ1DoVL7zt8cdPxxwWzKNwOIGxrLG
SBpSzxVk/zkUK9lMxYXmg3KB1RNnQuo71CrcDBXxrUcJLnnhUQWkKOwKUCd4j3Xg
PQXgHdF952TJNaE9qQ8keLWCBh+4H3uCxNkGj2M2A9dXWqvCf1fps9HM8hc4MODF
iXnnnhT88srIxL4moiHLUVQBxhHvexPnk3SKQDitYm4iKdT4gIrPMJkm6s0Wdn6l
D3MPe2JFVaMeqpONMFq5MRRrD7q71x2BwCGDLhiEp9zTaEM12DNNyPT31SzXUSKu
DbEr6iK4nqIaIJZk530ccRCBf4XHOM5uNiMFkfC7RCKT+2LHkE+Fy7uB4YpwxgOe
109nwF/wmwoSDSKiIVmP5zMHIt5WqdigE6Ck+DFrhDvRM+U7xMJys0nCOG80FsBK
RjkRViTMrP55tcJd5MhLNxpXPjLuQv769+lsr8iXVhBf7G4e2rBLzSuCrh52EZv8
G8PK/pJBocu+384hRlwFxP1MEmLnlnQadSuIOHTCJGI9PCWlwDv5JMOUOwhGd8Xq
cCp5U8wvAxsx4IExpgiCPS0+IxcEGxmy0JUeM56semlnIjHLHZMjlyr2M4AA8Uug
B27rJexPC6Zm0ppPxto0AC30zfQJkiLGR7uu6y+DtmVY35PNUJ35XOSz9V6nuwgL
YNewcY+qpmMexhLhgvAYdLzkPGYQHULziAXFDCvDRVXg/4dG+TDoe2pBqTNwGVXW
iwj7UAUmz5YjyUMmuzvRoph5ZN0AUmwsbHjpMdBF0TRU22X3cHgLEtBpFBy9tXo1
mKMxx2tq6H0n4q0tGhGjQW8f/6PHsg3QeWvnjUWUhmu8TMmCTg+IneqIBkzukacH
cHs867z97OOGDqEa1KpsSGvn0sjzJF/xpUGbomVXnzLxtAk8JzgLCU8oYstscAw/
glAGXbCf4NO2j/qofgNOeVK6RDVgRjnomHfenSp7ME44suHwz8HdAo3YGwpgGoIv
yJhY5gRVYR/BiK8IWX9M6BGlFnLMcpC/ABfYok9imIONv6qSx8g6jM7yceJmiF79
vZOUFrpWq/FAHqH7mPI0Q1q8ho270TZZiiH70cuejr/rgWYO7xXZpzP4B4t74+GZ
fIpVOG814SNdUVaHZi695Hw9Ypn6mFvorgGlGndP3Slb7ExcQ+UnCUz9vMkNXkLY
TXcKDjysy90fjXwN9/ALMUzpPknFdg+JmYmYXinml/qA8w+zalIlN1Kj76bwGccj
KQmTCl+77HCt4A+NAF+5vs5LOprIx6mF3GZ2qzjWzAyU6FxSEb/3vmJCrwU7z+Qy
bDLgMnhAOc7CIngBJEJrTzt7b8et8XvETKqnL11EaaJBxFzs0h7Vf8dhfb12iKw1
pW9tgu4kCQZH9QvCZLYKRscPVVncf7LtG2L9zRwXz5HF7UgsyUOQvd8cDb0Ovm1w
VCvsNxahTW2mr9gZOElNZeaQima7WhxmxTWSGK17WfoHCQuPGQhyqy2yLzAw5Yae
fBnUum+OSVcdv5EtScVEqbpHrxe0hiQwRE6oTHaxSshhzpK/CwJ/SAfGMLF8NvBN
ueawp5IsFyWRjjVV/Z9GAUTSJnpPp5n1esQXXVcN20cjH9H4ICeUiMI7Hp2i0Orn
rM6DEWah4YXx2d6k4c6Ep1hQ6TtiSQfDpGBnTvpmZlKsRsNa+hnYM8kxUwolhMbB
6nMgIELAWZuRhoPPB3OeTS41VsbiJ844nDy3hoPOQsXI8qSN140Zhdp8vP66B90G
kjTJ2R7aAl6FtbopQreKxPMZbrTcLGb9uJceG9S8xLahZNBqI7fganFLzznEA850
c97gZDnbhicVPf4v1/fHSSnddgPEoIYXQhnhZrA9SjlXLrIj3C0BcvwIZlKmU7XS
kSmuWdsxPngwOROWT4/3bDYwsiUdFrMg7YuV1ML7gt0Yk9fsJblJkvvUYA5w8feG
I2dKh5lHHypAPAuGHIig+3Msl0cPZVuCAB2cSZpjO99l1/AOeJDLER1JaBn99pwN
QLTTvRxY+tndsbMP8h6iMjFbiv2v6hQbttbePXqnNuQ9eWEbpfqHCtF0DIjcB6lX
s6vLOfiCSeSLwZVSFqSMumE3DYcsbvyZFRpK0rbtF+qAS1Al/UJtcCRMPyoEAzGU
rRT5ZaPOAeK0vQn+bkWYyGWKCNf4dflFiS+fCw6pfdXkE2TbLWTGyzna2gfYYEQ6
qr4GbiYz0tKLkbArJvUd0fnBvMzi4b2+jMnuhPu7jhAXE+gvzWg3N02u4fgZlOB2
Gw1fBZtx4HIyCuILzQG2Tzq3/UfWobH52GOw4BUW3T6dV4ZXb6TDToXRdAqH1J+0
YApD3FOwmwSugrCw0Es3ZtXWMp6DcChArg7OqEuBIIoTlmibhTzoUMZhVwdvh9wf
cvaAxWcFiKvQNGU/NwLL1hhJSIf3PhlFBYbxylvT/k7pBinzxafExatgBIEdeoIC
5yd6NCnrI4Q5KLchpSYZmU3BsAWu8kjdRnrykDaqne2pWgQ7XU4klpY7wdSi66Hl
+5mUD/P7az7WaTThJOQIZiifUuUYt0NT/DfRLXL53ppnBHpldggSzBdP15P0yCC/
43ytZN/AI7kH3Ty5Ovc2QSrTOIUf8A7EGMUlSssM1bqH4ELXIhPXtuQq0oTIiBCu
1lBRUvIB2YVR4yKrLzYh2rc48ilrvIZcWJxf0N19Xy8FC5cDfq1q+bFQTIASG6GF
ktlLZM6KeGNivOzKqKtvkXkzrTGl4Hq7X2FQsTb3NWvNS0zbLoekibyT04zqXACy
cNA/JUr7JB8Q9GpcyFOp5uT48HORS2/JzyGWlgBfx6z+rDAi9RL9bi6x9UyKNMR8
3/8uyKBsIldB5N+8AC3tfL/nb2BXfOCiZiGRil9QGkGDhf0BFdPytmrlOMDqxNre
3qchiLiOiYjHoqrIFHsgRUyIiZiTqSoEspJVvggmf2q0f09uyy4zLyCo15hmPuk9
anoRitnHpIGjt9U2gLKZTpHjPXHD2T4jDDKy/X8myVb8/1phCva/YaY0sRLwLP8N
VvGWbztlWdzsWK/w25Xf55By9zDu4GypPIPJk/wTy6rbUvMJHYIowrsBfoAWbh0l
fauqMKAjlS/DtCT8j4W7fBtQZl0dzcXWmvLCbfTAVsmJp1rlVcSoVPa1fz4Unu5k
uQAVQx6yvJYcpKv+wek88iSv2R9Nz4JKTDtQTL7D1TD+79I038PqeVAWa7dBkrQh
cGJcU3w9wqsy/uo52SaOwB+o3wYPmURg6qyAYHgTjQOZhGNRUJ5kYSupSucl34rK
QOXE4tpCzufMivLyhmPsA1NI4fwD5xEMsuAqSjdoT6aVTsbYB0/FFNfmqARaUVWg
HyK3IyV4bc3yorUXHzLYoC2bibIKu2RrBNwS341LdN8Ay/dhjiwzg0bq1kpTFl7z
AkHZmxHS4ywEm16LHKv+cs6or6exyjqo43KL2K1lfgHmwliEN/i54e5IaDxL1vTt
faA1JOkDN3bYh85gtdju8UuF+vrNRpvtVpFz0fvZG+UYaiSCbdwo6d6CxpwyFnIX
j/+dY88DBzkvKxdu7xj/sI/OipGgJwBHbZeav7vw0NWizaS35y0dkv9ynIHiebWc
OpioDe+s9ByAFptpq7HjHPV0xLat6/lf4uXzdbQoLnnqsNjg5YdbAoV3sDF2T5jk
DulBrKvQAU+Lc0GrlPtUC7Qr9ebGWhd+nJFl9lw88tg8wjGNPgu/BEUH96uxoJrq
6qi/90BAWR0R7kzycmxMysrx0B0p7oT4J4BLUlKXEPP0xGyzI6nIGSRW1L2lOdaD
1JNTWLMu2emDJU4Zh2aQGkFpIEhJlQZvoMb3LOIjL+B11/mduxcbI/KkfSIom7Jn
QVhGJ9ovi8MSxz2nYn/S8RaOd8y8UOtyiZk+y0KRh+Xcxz/H1Hs9c4PR9sduvHsm
0KcatG25/T6PxLM1vfzh2dDTvzlsZx7VkqkkoV4Gz1m6uhXTQDKW49Gl/52vNfJ7
tyUkSlY53FYHDCus1I2TO3pqwAznw+CtWgvXzkH57QjLVHjz0U76fU2fqn/dR1WK
58j4puT7TbkjHM/1IlTBfAZs9BJ/kENFWUka+UD8Qh5AIl43yMQb78txjKFJL3Fz
shY+ErS1H+jLDWcvdQSUHYDp8SvZfxYzhXaP3Cm0p/zbrUBrdDgb+NlhVeDgXLa9
Wgl4I2NeXekC42g3lknQrQY7vfjVJES1od3+6g128tAGAk6J+IOYoHv+ftlCyPlp
XfhzolXfk5QxCjI2hPtkTYzbE7i3YSh1n1s2JqfMIWb8I1RsAT1hY0QEXrQaqCpi
kzg00MPUEeS+l9YJ1KB842PY/GbyENC6VPjoHSKOG3QzIq5a9Um3OKJN20oGob3V
A1z9xf96UMTWHEoB4l/VObxU+9BjkbsyquBHf1TPMmwzFk07f8seuJieXbdn+UQE
UEQ6j2IFIzNCfSXr1v9ZaVmef54tkySVcTPLILeDWXBNAJqe9uyq7JbgJiyWj1v0
n1S4C6aXPG+mA3kc58RSKX3jL9tldhw5bIRbFN39ZyFoVxWGkCmRfAHR1G8poVrr
h2sVAQ3dNr/0OUWrpIIScyc95kLIPm5sLjw6hBfM6SaQNecdOcdsYShLwdSjdzjg
+5orNqZxg1mO11d/fQek1cnat8sCpP8kA5AXMOlpTWrde1HCxU49C+WMvNtik3o7
RN6zkzkzz5sUA9XbIdTfx5KV76egI0RYEgZM+V84ox3Y4jYCrHo1mGbPXNDv6SrX
71VhSN4OJ9ohvgyS4Gdf/wg2tfnF7jaA9hZkfGku961pYaKd9y9ZLGhUzrJjKrai
hpTHy3dGz3SHFcNOsZTm5I3ReVMuwKFnUpGkbDOZKc0Imfk/aQj6Qc4WlBGRNZnf
eePy0zl6QENH6Wc1coKzPvgWMRdJlF7PgMRfHhLvCmCaemhoM1bibOqr1pnBqd23
GzeLcldSOt6VXnfJgJygUEvFq5NzWQlLKQp8Rwnnk4v2VeiULCIHnS6zmb95ZgIT
PS28RqFnO9mUtSZfF6Oq8VfJ7+RhGMVLsXnzAKvONZGByhQ9FGiqufg8HULdND1Z
p995rK22M4bBJaLLgFnfTYQGO9wEFZsQNhdHOddJB2m1CXWl66r4OImqBuX18c4Y
6NdYUF4NgrrOtmRjoyujweOTfEe76nqrlzqCPpSjoN6jayf8LV+QKwc1xd9geBRZ
QhZuTKP4cx9WKXq4DxgaHyzUCepNxve5qR5d2Y7y7eJ274fQYwfhJAquWPOWypOy
Gd36JBd84CkNY/nrb39aLoO7IdaD0m7z/5Zrez/CVHaLm8mgf5fi+ImySA+YuIE3
nc7/tidhSQeZ6BHX3gPRnk1aMXO+hckeFnrgCmQ28jC/CwtYX5CP7eC+DdjaCYGJ
kUbvqidQBbYrl1ELbwDTFnG5pO4x5rJzlkQ8brXEIlcnzJWZxDMJCmpp/jz+L4BK
wKYeu58G2OkSrf70c0mtVqePqgM8hkl0oCfaZInHnhZ8DBCkrwiN3jhlDdasur6M
dasCSxTcvNixfNUrUgEaX3EERTJob9rxP95qXGOKmjXsyceHY2dbDCuzOJ3/5NvJ
lrxkYUn1IB5Gho/iAwAIP0pm2V0k3Ck7Jh+E/bQS3MQVdYbXhga6ig7Uw3/oXy30
b0ONYlL0SmIa+uMQWlB+ZVrskE7N36bf3BciGCPLW6NzYJpTl4insvJ3RDXjC2yp
5bsrBPmgA1mxIX8o6EXTVa7bJO423Ftlf1FbQbXbXMoN29JTvH221sJ63B9fEGlj
awZL7XEDnGQ5kVXpgflc2pWgOA86vrR2FNZzZw5qLMqwWNuyO1PgkxCsH9MJR9DD
SyL00KIT5GYelp7rnuk4gOCJwuuo8X61yHL05i3YI8i7dqsrsca9Yi3eTxCKUkds
qD2eIvBBvOypx04dxDCVffJX+YNu0noeRRYc8eK/XCB37MJnFmOtoA+6Gugvi1Oj
l3WKtl6yFfnc2Is6k+sKTZJ3PRPgK4Ffv5+dUKqthXvlucHvdqmd+IoT1L1fdxST
R3PptcXaLAnlo35FQoYLiJyvISA8oFulXXgLehUHeqb+5DXGE2zgwukEZbSu0rOy
s1DmU4KeClJNoqdGSJWuYORN2Z65WUlg4B5FdvusLRcxlMFZiIgInXu61Numi5Pe
Qf/fl7eFCaxzMM8gnAegewCxrAq/XXfoCH0OfBV9Ibr/Y1uTtR0dS5lC6xDmtYiz
ldxn4DsvATwXu3T/EbAj0iAnllFa4hZST5WNnx1xEzn/XozTcki33YLIFO5yt4q7
NTAB+A43AzYwbNptG1R45tSCbYLBO0rYv0TMR2+3KpNissH9hBza3r3OpvpcLW4J
kcV2tmh2uhJKrZx3/zC+wmXB3MYhxF3JDpVIuhN1kdnW8BA8yx3U92GmceMUZ7UG
r/LIcvR5e3MSMgRQsA6RbwOSQ/i3qbbFdq/zjLjEwF25RLk0MjrBBiEmukqcYh+c
sVQjfaXpC+a1rN2mx1z+0sGXEMTkbW3UIp6M3gSRivPW3zSKvD2Q+NTL9Od0gYiR
j4n8wTulPhRCeqcDmNjlWIaSZ6B1jfwKf/jf6lpI5AvuNdS2XnhFQcKSVvGrRrXH
va7yTKLz8lQR8eY7ZBWAfm8cJSQlA38ceXPVjvDi8gxdtL5KU5Hs9aNceXXuoYqS
w8zkjdkLhsTzJPcqt1bWCbozsYqIyr/8DVH+NQU/v7Ys/o+QMQupaLTbKZcx71hC
Y01UqmookUUiEDRQOS4nhuMIRzRYLLHKs9DRaDlq6f/T+dsSdo3Pr3AW9y4C/djn
lsAHRM+lhQwk26D+G98OTBGm9dzd9sx++MnHtb0TpcOImiSVYa2v/Q0NAvarWmDg
4bZdrAGJjYlO8WY0WEoQO8T7wZxSF1NugBMrqv8VZeLp8+YG1PG3qq65evK4NF29
lJCT7ef8vXmPDwhNxAZScaFC3V+vEvNfNZPJS95Jsu6vLZFU3O3pMaaThdnH+H2V
nqPtUDttw97Ht7mMc4yXRy/PvB3NurWuNh0aZ5rTZshU6jTKpaN9GvPRlpgjpYzh
2ZlUqmPuW9/lQZzCAIKztWbYxc9kJNvnw3w3NCeloG7D6SOJ9DXztn9919NRgFjQ
EQd3xPdFhmNHi94zRnLQAxQegTK3ZBr2Dg62r094mZ4PG58ACa/MjzuiiYR6S0wC
cfD+VfXh9t3xs8rwtwoJWvKkyE9n7mK/BAAM1MKpMw95Mi1Tbb9VGW0tByDhvQvX
Gj1gBfepdbQELdJzMJkcvxV6+WtGU0Zopi7dLLvzKvRFclClemeB9YncnUZqtAx4
nYiEIdP6lJye4q9hzf7p8RDbv6uZARpJ4XwcX3BqTh8nJE9zRXWZNqWhLK8YTqZ/
VEmGwCEirf21ApDAampZw1bWYB/J8C9puXoBh1xI3R8clUAN1m+O+CQ3QM7sQrpH
d6YoK+T11J5tv+Gv2L3jSiwHJ9sZ8xoV37V2RIDdt8YVp2JpZ7LCTFvpkVfJ7QNK
HmJ+25Mg0KBHEldhoVy3/lqqRgObFjdyt3Onr8jjeNRhy6CNJU/lZfEgKf2qG7ds
xtiB2SFuQQVBSdzbylKMSt0r8hvsoSIDIaxJJGqKeTjd5FRi6D8KtiMJSvS9/hMD
L2c2bgJogY1AoPjlA0YVHoPf3KoMIkoz64iMMGl19z9MkvnjRIUof8/YnNpomKpw
kNaS/E43nJ5BKwYPtrQTn/lq1FOMGFIkeUPpOlU8gmRARCgReVukCwwa2BfruDqf
eBzPLUrqhklfrD5kQPQtZ3w0nCflU9j32sEs0iBDbyb9jYW70/RtuZQVqFuFYABT
p6MXQ/DMUTBdyI42rl5Q7fGNaadKAJchVzaE7R5DsBV5R7XSldBL2o6rpzCUco4N
NNxm1XzjD8AIM2S2yWwSV/ZqEDmRsjLxfIpJ2/8DcJsXjmieDsMAOom4WIGqAeXG
ZeLvI7c63ldGRaMOiNgq1js+xPpZSVnxE+V/lIW+KL5gTxn0ty2rJpWkCTzgpSJv
gsuRHidCHyNrdbiWq02bxXHocuOUnT5tFt2sMDZq/E5NlPwqIR9ml19r188uJ0Tz
MCVnYQOVsyaZBj9odVxDY9erVbT1VMbIr8upeYdC2HGIxCpMLMUaVXs/RdltUU6D
5EUz6Ax8f3RYE5kOhBTdewPZK0uWc0VX5WF8D70L4TyunYsLvNVt9vgJ5C1oDCvy
cI84gNEi0YCuu0xeyPx8o5QYtABl22dR0rFNSTyjUvMbbgMF74j9ZO600e0i5Quh
+441XmG6xdvrILXC21mhurG/Dx97o5kKH1qV7v4k3aavG9vv2C3i8O9mYc7+5MSS
IF7690AnYYmnDanGu6eeA8675gZeHe2rb+WTk2H0mIwYWFmsC+S8Eyod8UyU0EP4
yeRnXsgpNzoxdQL67y+nM8ScNYMZbeTQvqosL1JPVnDXRgVlcqXSRDK4iB6L7lRJ
rOeyoxjRh6I1VdQdzi0D3hGEIku1snlicRCS3I/6pIQrZORNqdJfz/LaCUTLypNU
0irkOdlj8Zr2mxjIx86Nmqeih36EaXE9EkgLCGG3BGShdOP/4N88P7ibg3CT9CJe
i8tOX1abHPSDOLXMNNVrAK6aHui4pGbEuXH5drsnna2GLVIQaVqAU6spofUTRT80
kK+TNwt1fk2jNgNYk741pmj+Hh1YpTALZOwiI3//D7O/E4FmcXbwTrryXrLhgT+g
wIR5fZBI2tgokU++FkWqUGlgJ3fbicuY6frPQoAXsiaYRhBz9LHtZCL2nMQQbBXD
n76sxFZ9iYnMQx1gBRZDF15+Ajrc9j/Ff+yOCAeCzKohZIh+1SKN3R0VojHHOEnA
/AcdybyUVP6RWbJB2Wrh1eZ3E7y5AcIWjAKsFyl/BE5AvMiKskaVBvKoyMOX7BSo
jwRqkmD2LHsoaVr8nJBANMCBgu4tMf8+pOsKMkm3WD+3EjprBq3tSz+sECRhTDyA
4A/RhCy7lbCaCS+lp8pdhBhd4oEUL9g5+WpugAoJdg4kOFo9Kgvz1f588uetrz7f
/UCLyuAqFQMrNJWoBStcxvjM5HRl6MsX4ZOD4W36atN82yDFEPgVDF8Hs1BvsD9C
XHZir3ZFyKl96/hxtvUzTopaW693hGcAyyj2fi8XE83qvoZ6nuKxSEST478guhtS
W4EDYcvoCIlEx/Ff75Uq1c20ZnW5pq8eQPs9wK9PVamc/Kye7vCGpQCKD9OwpFoC
37iC92JGZQ24QkxSmO9iCTwsAcK2Fo2+2sKFLiQGADDvbkwyv/G1IKfXhOQGMhPu
vV2vluzqhZcrBtdMTWMy2VKYNx718EvDR+mhzs3KDvOi/mFM33QIrKHuHpBErzcg
XA+xaMtY0HXR4lYptG3mjXQIenVaZBJH188PTj488P6mfOBd9B11guDZ8SEJWxtk
ODIZAB5br5DNBY6w1Ikj3D8pgSv0z8PrRBlqwvk2ouXzEnAFIVw0vnCYx4tYlyp/
cWbo0xYlpj2UFki5lCcZZcvI53gZBqeEXCi5jWC4KnR4/bcUha6kQkorcR7uiPUk
KrT64SYF6sxCWPJgkPaaLp0OPQGBW9JSGQ5HUwGkG7uC5ISCrBo/+yGl69iyU59W
l3LFn/QWAUfjCIIQ4cYzxY7KvKIrKxknkxhqW45wK7wwTjWQk5oRG83qiMPBwmjo
bJRuIRFsZy3zaCpuWvmmh3osRvp8fZ/BP/TbH/hY5BL1MYLHvSc16vZjBGuYttI7
xGhdOymrb5283XgtpvslIOHwV+CY+yH/0hjANAly/LY3CYUUZH3m0xC+7lnQef54
XGb17c/gs4SPxbovuY6UTM+F38R9KfYFJ+zau07ATc43hLVGyB9mfi+63vDbMVIH
eDmTKIX/acAM8b1JMxdxkVhKK5CTyIU7LFewRU1ggtX/rXKu6KQo04VpZn95Nk9U
9Buh7LCRZK2gWEXm6AuGwuIV4GFoOdDQIP1V0M3UZ6cBs+CevRXGjXhsbiK0BRFM
Gp545WGw8nWcXqJ1rB0HdutmVLky9+4X+Rip1n9kfxvo+srWisKyM2GZSFqt35YN
RCmpstIEo1dnQfLJRmSjsISJoKCwYLUaIFlD0iVSPindHqDa00o0Ea2/9wc/SOOk
7FvQHFTYvyQM9l1bRSEX47gATMJ17KDrF8AAL1vVqAt9Oq8YEc9RfPsrs9C9Orjo
lNSsUWar7SeY99k2DvE7iBJ6KxbHO2X3L5tvQ8HRztrscSQMkTNQuL3bht//0N06
ZbT73bClzbGJONYVBqWshnJm35k3V/Hm2IWKHgDlUg/x3ISYC4KSvzfHF4qVhnvE
EVocWQyxUMaWT4olod3h8hrn51ThN9EFH6pEBPfxb/2u/LWnDgk8cMfHdE+vKb/g
a/VeyM61RJJVjouaU36Bm6lMDPbsC6fdvbkFROJ0+JOgLOuiTe80Ki7brIwv0Dzu
XZ5L3YLt8jJMA1qI9IEvmcqXYlY4cndLl9EFdaVvcIMT5TjofLpb4vhBR/6/yCtX
Qmx5b1NJ5bjFysXOEGKKIt/65z+Dqw0cVkhxiqmIC5MIiq5woY+sM6Oy9pjoZEMC
uovrUB5ksjgBZZO8SFTELp9rpILfyzGKnOiikvuzDaGpXvZTZkaRbOvx03xDXEtO
7TEI9F99h9tL78P04V+2tge5bIpkvFbRNy1xuOoY/LtYs+lyNLyclonwaerP0iYe
2H/M/Q3q/rQm3f9e2/cSIG0jqDhQEx9Y6FEWCaINoiNYaR1V8VNMFVy7XNAFhI42
gpfL/EAwsrsFoAuk592fzHHd0E4v7Gz/wZ4HYAV2BntozFkTZBmz9RQ27UFRsnju
N/0fg3mht+P4fqPvB1YXll/lkOJg2au1lj6x//4MCf7WmRfJnWoxwim7DhO3NotY
93Wx2+fr2Z+UQI4+3q6AE1asg5z0x4QbE7W6AulwDzA3WTmGfiEnuzvjhRGCsIRG
b/be4IVw1QjPxkbBg792Fa+l2r4PY7G/iTmKBjkZR3SORfNRCcYEiCoHX4avAgEl
hhQ2QQ6scs1QJlrzqT/Bj48NivB6iPvT1dkc/9YB8bB7G+WHLFImPjkUxC0p/sAo
2Np9u4ilGA6B7dqgxEknPdzL8timSjjg9E2ZgskMvEEUvPPuooRBs/OEaSoveJ+R
sgzhMoZm211iVL0m7j0e5g95b+6piS/Gv7EgfMAe8aqW1tUp43M4rR+qI/yII2+/
oGtSkDPAT4p7qcfERXVtS1O9iMlI8hmhBiw6ktEjDNo8wJP3zXzdzQIjNe4MBJUH
AzLayfgnGCHT4I97vQf/qlI/g6l8SX7PRjSCldB1lB/h8fJeH2m+eLCbKUgpsPVo
lQ0ZKyr4In0IHAjdz3T+1S9ixfsZYpSvVk9byWlkkCC6xxTcvjpGF6nticNBSF7l
xmn1EHDHr0h4mfIKMXxoayeXPW5cUXevlmIRQb3Yu+VkcPpRksdbbkZLjh3eJp75
I9Awc/OszXtPW6VsKxouKFFysRmx2pOag7GbpDkVLTMwShnk5YHaAh8l6TbtChgs
XyuwmPWwjATkvuBGtgGhUtP7r5JuCybEh9Vv6k+CYjtNiEZZ6sNRb5EoqwDzTDCH
LAcyeVkAudI+8cM5slVT2v9nnfdY1kLaeJlhXPdzrcVbVobZEM0aWCUZjtJJR8nD
vpfPR/MaiNkE1gx1sdejBWvhBOPfBJX40zU/xptXrvQ/ss0e5YGsH3oWOSJmdKQA
QFgWpf4WTH4z7cZ3buqG/g7wvx6F2rgew52KoIrP6Gze9Dd/Ny9BI8BcAt2IwFP7
lohJ6uLeBjWDg04XWR/ousMVwDvRHZhoP9FnZ8KhXFx+pvcCm/5ytrwJc1oU/KyX
DGqKigi1IspFNqqas90zMdFtbfbSOzkDbtES5GFd78+hSJ5+h3Vx4pOEf0rXkXr5
i+fzjxI2Sk8JL3RYsueNXfY7RLjeIp3Brhs5fP0S8MRL4Jqbm+3bypoKrgXVy967
T4s9gBbVTirFiMA03dOqakJgnu/uveKpEtv52OmCAvl7FnaiQiOm+FuasmjHVG5M
aTRnmWypmU02gdlKm5Od0y2KPZ6T0bxoC5p78oG3rBU=
`protect END_PROTECTED
