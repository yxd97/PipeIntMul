`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WyInp5biVGaR1patSOFcmUwBp4qNJHkA3N7Coi0Cg5l91UAQxTqvtgOS9JjmLEKg
LZnttnfnC2hh3D4VjTeHOTLcZzMLsaCl+kijAE/c7knNjt1b8d/NtXGb08jXUbvr
qqe1ow4RQrP/7WWVGyxgZoUDDl15n2dfRgRSru3/G31V7DhLY4Xwi3bzIIEwdt/7
fNIv2UKt3smyohWid9hSCi4Zm4xf6oZDhpO4MaV5Z9xl1YR8Vtq/U50Qz30d2mBc
x6mJrZKsd7NwzlxysW/vkN4dI15t3X8QgBhqm41LkRUGVI3dUbnOAlht3L7lqnfo
yKsJ+jTsqzey893aGuDIA9NtcopVDVQGmtf+VEkzd4kn0f26W5OaM6kCdiJ3pdx2
`protect END_PROTECTED
