`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bd5t07wVji8Je4M/GepUta/+Dk0NAoBoUd+Jbv7l93Mmfb3wd9BaYa4ryGx0q00+
1a6D+6x0hhgMM1vKhCmKzKTNWguql0elmbDFYcdsTd0gQyFw0v/BHJlHCC4kxCBC
lL0IfKJYl8hHno2ImI7Umg3r2MVC0vMb+I5Eno82x1pDGMh4akY4qq+1M/jm9b3Q
rNFsqczjjkSvYzKGOmkoyzIiLMr+Cz/K0BOk6v2itRcCfRL0C0aspDTsqALp8sHK
YmI7F73uTjOa97B9+Kq9jTRTFVAV/nMlAyCrSn+5cAw=
`protect END_PROTECTED
