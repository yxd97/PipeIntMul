`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BMkZJV9kMbVzwZbr5EPsLyBNJpSpbASMqRqGLEf3irVI2z9fkGGmnKUnh7q2wMQi
hFkxkFg0MdCmqZjggw89xZUX1duRdZVyLsmJuTNkIWR9ql70IR/4zydu/9pEttNS
A3YH1VF0cdKP84uhao200PfDuPOBtWGPTRmJVWHwxHQP0XYpweA/IUC4c0sdTI9S
PJIz4wbxPQ/ODVkyB2lwgQBjlO+jsbBTF+YLvRB3IiI4Gk+1bpQAI6r1DSww5L3k
w2v5H8f55/a2BLk1lu0eSiwxdgKn4jKQ+YfM/zO1SDJtM3+z9AXLdPFu1MKJch3i
sabi6OZAL2p1/H4zL2IDd6SL/3P58Q2RBQ1XCVfKyopG9hsv0jS7P3Mh6xcLLYkh
9B+Vvu9P34pCQjFSkki5kmx7xsYMS/xOSXLU54Ng+9bFcx9idg5QHR2Y9qtZOs/D
VmjVgW5pNmET8vvUbTracYk/RA2bMDvzVVc0k/bIsV9ecD7vdJPL5xE+fuh5H/l4
wA+IIQ3ucx/x+fWDuCibVrlZbm5nTZDFOZ3wibO766nc5u1jNxq92eGEYQgbQO1c
MqWl1e0p1c7P3qJT33rk/osE0ICZqyk1aVOr8Gm83YAGh9byFaPJCTrx7uFoDK/R
Uzzy19moj+EyhThOCTlr9th+UYbb3iy6HmyF7I3x/I+Q2ao1jPRnTxMLMcTqOfGB
tvMs9C+QUDer39yufPUcf5TQcum1yqM0da7R/FGrWW0//SutOOJUDaORpJUlLiKT
GXQsfHCmomKUKeU00hMpiaxYCopZcXTbP1+ckKGq82wc7zT+1LyXF+PQDyUCCmYj
Bk+XHuj01nYZFIJySeYVgiBy7pOcbEIIqbUw8J1nKLmFZGwYDSgJEJIvgbCZdmEY
dh389PYV82lACjjVdxOmLPCAGpmBFknRVo+sa6bAH+Tc3Ede4X2tPPK1K7c64sAf
sVdMJmF4zHspvFj85dTbr4sOWa47G6oQuaaaiegWgWTOUDF3qtFzLUVqa/LfY4X7
2Z3V829eAexC2Za+/Oy0bryhH45fSV7VAvE/HkwADABgRcVWfQcs2BTRfiF1M3pS
rJ/Wcy6W5+xq56OJz/puzE8QObT/pjWQUrPql+EyjpsHVNRkFx40L2Q3D+gYRuqm
07aOme1Z93wx1dTjaN/SboqhyCo0De4QUYMhi2ThYRF1G5dKJGYbeyyO1aFJgzX1
kebrLDKZBOMgnvPIXnRK8vCRiRH9bsjHndWi7wQQkYjGZJ22oH8HeeZDFbnAIrar
WpHCO4yG4LWPOG/odBCPjJ2F4MYZ6QBnk9V/9jCNAnHH5RlMF4EomUBR+zWgksei
Nm/V1XKW+HrACGzT1ZblZcoqJaD2GLj033nFc1e46tdOd3+zO16L4OhdsMbzkGw2
dpr3Tb/Y6IbHE/Qz6Fk0YsMAmDBkA4UxF/tjqywQ4HsOdHqQJNHlnsBvIArxBC84
HswY4W40Y5GNOXS0j3OfhcpmXRipIJz4HRes8iKeybarPMPukdejrI2QR3jMEqFZ
ypziQYAUPmtmZ3o7CheJn5IRHn4FLoEMbqitW/EQt6souKEcCHv65xJZxgk4xSl8
UqfPF8MHZtS1F3QuzUtJ6kFtci6vsPBfw2CGMS+zlJpEbAiu5+vxQOgb9zNMsjGs
0cs7hHAl6wmDsN/2wMYWsukjKG/OceufwkmOflSqPjK+o/FxfcnSiwlqjfx65o3Q
88vYlTj486VTtdj9E+pCjnRUZnD3B9cGBv/jqAIopQhYN234Too4jqXGGdFkjjzM
T+HO4LRz4TrTMSzkh0budpeo42cEzYqKb9PC3uZy7YjvTBsewOzAVY/PQc3WI4Lr
+Nhq0/7+RYxKxq4DrXndLwV+cUSLzSoUZ1klEwN6b6nYHqMxRj6ZBYF0NoEyZV06
2oFUcvgai3F6y2R+zelblRrXuglQvLjMeEPhNNbjwNXPeBElkoHVZQ/sG8uOMelZ
UjPw0kbEfuC9Fxd+M62vJ2eQhUmM23rp2nnC65pvkXvG4nrbbs5Sa2CJAogZjsxH
zF8bpDd6ELo/TuK6AdZAwSn3oS99ucuBYWYokF73pJljaSeEpyQcoxyBHdhG+ZOl
EQPr5mY1WX6fC0qxX1h+cExR2BV8ak+rWcIKNSBP/jlzt+ymms/j24x0c3X5AwSj
BhhDb+MJq0de3KXthYqL6dYcFFmAqD0Kfn9i556djONeqU9CGVWh9yNvU5LUzqdJ
80UIojWx+36b/J7smxcSCWTopn6SkT1Z+tArT/ELNQ4wKx8GBKFHyjMGSvNJkvfq
5g3+zKsUMRxLSztDfiWyw9oLNoL54JrWZKPzRE2XxESj8zS8W8pHawa8bf7EOfPi
OV0+5laGx+UP+GzhdTOph5BNiH+3SzkSUgYsudvgY9HatWYUopp8uJCl2wfHdyLD
VeCCWche8vqOQ2crmlCeQaraGiFVMQZuNiqS0D0ydYByYgWaWHcMv/7WBBcBHXFa
vBmSPny4jsMQlJ0nw45RvWv9zCvVsJGNkj/RK+OFoG3TcYhjAFRJiWb4u4nYiIO3
FECDlWaGVnZOyxtHJpVhl0tGIhEL8b7RuIZ7QjoiPrPofrk5XR0G8miZEQNjjDdS
g/kl9R28Od6LERLTOAkuyRpSoEcfdI39WQUOYcTBfLbHly/XS4LGaOaPTKVttuAk
qOT+r+AoRx0wONMp394CuyshwqkRQ7vEH6IyngaZiWLtf7cqtsgUG51mDnfGQ9W1
+4mLntvp5+BxaiMeLP+xJn3BWC2USognJp+3Cw6IJW9vGCzhnDVAqt3QBG+6KrZ8
/txiCaJXnXexHO6eiV1EzHdqUpyal+CmACR8uuLwCGxFZ5Xu0S6oVEv8BYiVpIGZ
MBRnS+dJy4LC67UkPj0ZKDthmzgVUrP3ELep0hmwzFeI/TPuNt8dmDhX0F29nHDO
4w1jz8YUlbDCY/cQ+WjJiJ/1lySC9a7Ygjr9SxIqxXGi4QL0lXMp/5uYyDvrKWwZ
dT9dNmT0ZdxxW0vUoZBOlvRJry6yBBmfI2Ydzfibs5fkrSxIe4P3HRzPIBpgUF5Q
xkK/aT6aSOY4SltqV9jg/yPPasjd1RutHf61/msK5RI7pe7Sq8mJ8Wyrwl9k0Gih
Gn91yicgCKNE30Z5xwiltESHu22QSaH6qQs62BV1+RvfiziONmdGFaY9EKKj1ti4
hJRUH+vkObu7HXZ7CuN/1VwNZ2Bz3kUW7aaMFjBJX397E3Nc/Qy5SNrHo4yHi42c
HqqD/ibwoXmIyP7xhKdw6D3lg1hupILMNJr6ACwRBenyUf/yCG2iEVWPMZApQHsI
JS+rVEKk0zmsNdbJmIUDUNmnZQCZPWSN4rT053/sraIXoO9obuojW1kiSHrWVmcr
vJfJADKPfqOzk501tDV4t8opirAUW1w/9PLI4OqphA3M96aat+4VJYdxfeQSiE7l
RhtasEgHyziWmW5fQef82BTopYhDAJldhVK6fdqBBPi2l3TH19fltKcgaLHhYTdX
MkiZLoYFJUK9cqOVe+Zvp1hTmqMG50wH5iJUNx/X428p5WmReyxRQDr//w3Ka3sL
DO0DlXmEkk+voj9xMnDoqzfjmxqe3Xg7O/pGVjqa2qMsCKR1Pud5wdwq4EqnRZ2U
`protect END_PROTECTED
