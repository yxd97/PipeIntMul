`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WRPMbi75vo1yFaF9yeOadGU0C0O8uZ2Dflwf0vVibCE7G8aC8HiMmw5FjOaQ3XQV
oHZO9jZTAS047Ip4UAE2xAv2zd5nBlbtQLZbbZ3eMvYymWF0PRf+RzDRMBWGSVU0
GUMPwPxNnCNL3oemPjd0pgMRfH+YerZmDpbURsGSNbYja4bhYCn4LjB/jiRcTix/
dfhNsrBEJzJa0T66hW/9cUUbLTuPCjBDnnILdFqhNQByfpGaNvVGBWUA/4EW5SII
a51j5ZnYG4SLSvG5rRWebA==
`protect END_PROTECTED
