`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1s72olnJj8iiXUNX0L4HR6YdX75MFPdD/q9DHSnheoeBlNintKUM2j8YTgfffiX
UvmdjTnDElPCr919bY7BndikdFe0a1otKn+LupAFDCW4g5JvI1MbS2fImgyt8gAa
zXMBcZrvNhvGsZr9u6sYFKVEViskhMQBYeSAuQlr/GOc9jp0axSVhXnh2LF4Lv75
E1tYNt9GvuoihoaZe7zHpj5IlAVISCkov8CBoCnsYru9QWfCKGYqyGC2SfDaqNhC
p7D3RzESxtNjf0sUJNAQt2WY7T2lMOZ+satyQ/GKPbxJLgk9rEdgHCohRYE+pKKS
1v5QPTO7XvKHzD181BOwFFUz5xjRwM6oWrgKLGsDIfqsr6lz8w4DVHvdkhaEpAm9
k+/O9aMVQ2xMl/yYYmTPMcDmlXY3ZpZ5c2Dm63SosgEjQOmjQzpCCSED4Y1gRVan
4QXfibI6RsngigMEN7wAWPEZCKbdFcLYill/Z/Yhp2+6b8O53NR6WOLphfHmXeIm
f1Vp2WuuvqUiLoADHdO+/xlEH3hBnnxux+vHGQgD4AwW1gEVzi6LnKl+zGZAYd9p
pw+7mXAaT9kVWskRxfN9Y5Bl7gPWfJ0CcZJTjarhHjU=
`protect END_PROTECTED
