`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dZnWzPt426tpYu/BLQLwYAe1gKjMV1O6Ycy49HEpSjzqt10FiAE5sMpdMFaEQ7Y
pbMcY6lSKblHi8Gp6/lsUpgj9S28D47xw/tASEjd9bZWkMFtn9BPeAIuTVi5NQ99
R3U+STJzZk0P25/+DAvjENk55Mu94WPYSdm0tl5pgKxfgqqbKNIbEcqq4SZTh0It
5ZRkqmWlMwzohuhI9xwJF/1H1mcZFsHfJfH0E9m0DoRbJ+LsKoPWQACOhQg+omU9
9LWX57rThQIwTPSAApIvMr61BSXQ8kVNYk1XNgRSDrs21M6/0f3CU8UGOlQZhwZR
Tm7k6067TGczSYZ8QI1E/TtXpFrnDS8ClA5wVx7HIa0kbRgv0cTVCRp8fSjjYf5Z
1lTELB5OnqwLey5Holj4fCchkhIfSoACwhzXljXGmcmhBLB5bTluUCheBCYE6DxN
CMMQgfWPSjHyoc9/9Rqu2RAJXpZE+cttm0SuTw6bz2U=
`protect END_PROTECTED
