`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6aaYU2AluL6rvA8U3OIGo3nM1pH4LAnTmpw1Z5vCaX/Nzg4BD7aoPeQa0ENmEo8/
zwoQQE9wyownAZINKkgCjqdj7PV6/jm+2Io2X/ZSSEzPPjBzbFJMZYo8OHNUBPlA
2LglBZPcp8VSlDDPYVArFCQwWJA+Nn6rcbs+VW44sgMrgZcO8TVtaXLH3l7TFUdC
yUotIEVeIB2uM0YcH/iiMFXdcnuSWvTTqcRi9cgoB21r536IE9vW77UnldGp5nIe
OZJBqAnQDO8lglS/WNBsbGnM5b52CMUTNCdl+oMiv1G4ojULU9QQjXPecc4rSSCk
Xb6gKQz27x3TUmdmxAscEGBgP+umTnlTr8NBiUqanA3qdCVBxUZR0cRSvXlruC2j
rB9yGZe3Z2LCKs48wk4KDuSzpdHh02DC30VPNg+m7aeUsc/7TaicLWrxZ7625xni
YHrYIwzGrPxvASFFZoGJZSUClmrXLSdDk0VSsujex3M=
`protect END_PROTECTED
