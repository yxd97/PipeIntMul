`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvwzoZLlDrcXEzaCUO4dUijJrNTuvhJai0J+2A623cGvAS5MKrJrewcND8Dm2IM1
ASWk7a3fzkm4m+rjzRvAJzOJ/XSKRH5jKRi9MjiqKQJ+qEoAq2Ij6WzD/1++47vw
/VexFLpBdpNPcmb7Is6cCIwAKE8JDMAV/LT1XDsuUMtE+0JCHtgpwksTf47Xwm7L
3qptN7pVu9VAW/KKkspQgAS1PeZrBPF+8mZVxP5pps11GC6sG6T5Fvhg5EVY7VpV
XBiA+MmfR7Y0z3T99Xe3QHuzjYzyP2SRrsfOGZ+mM78=
`protect END_PROTECTED
