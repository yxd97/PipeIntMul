`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3pbMeyx4zWxD9JyRRTKH/3zYYkrJoJyyuPwVMXfrAngVH+boJH8V9CwvVglyqxp
s0gfXiHgMeB7SjtgWFN1kKSEs8OTxbFy2uJ2DsPJip9od4SOkxO91KSn64FMnYkf
npR7jkavBkjen0el4b+tSRo79oGAIaWUaMMVU4Uea35e0tc+l2HIbw3DOHO6N38Q
pae7XBrDfe4FbqFasgJwktxrwLz2DvCPUB0neVbZdUXADThGSkfcpfZCHh4WiOuu
COa8uAK9L49yuVabYT/h4Kvql3kMDj7H/+Okm1gAxeI/scgJQMGgNd/NzjMl6XAx
+rrKqBRkQTkovweEB4U8tg/jNGFHcdDxdJffbsCCQrsnmTlKg6wIliSVNul/xzJG
vvueMT2soQwYPjpNY6nm+YYJUzLEzcO/oo+gf6u+ebnL2Ff7601ft78CfhL5ZYq1
sjoYRtGblRr3iRekIBH3fWFtbFZzcskZd4zrA0EQZ/Mx/Aejuy/YBLNU9br/Em32
JKgFoW1q6lMpovH+QUZ7TbXbzFv0BpHjv9KHOuX+6n+4j1x8V4J4dC7kMJm9j73V
kaViScOVPOgXZJQzWOQBfXIJCnBlqTG07J7KgoGb/wIS4w1vCoSyuAS7M1Kw3BYV
TafPdUwladvJDV4bG8t4Eva+mOWU+0907kWOKTFk2RTAKTLxJLFWo2H2C1uLfFoY
n2hBribi4V8bjBIo0CbiwHb3iKDj1d4CULbf8mMqokPBXUlkWIv74Md8xQiznUGE
ffeOjdb6bB6RHouqLVn3NBkKNqffdzXUGE22uNMGBcaHrPImo3K7cWLX+WDsu/7n
hnTn9U2/kVNtTCWOK87N1mgyw5DN1suyZh0tkUu5Vae0opToY8rtRkKZUDmBvxwp
4S/OYsQoUCynmm/1gUGcxFMo99j5MTJqozeAUUE2UeXjc20m1fOWOsm/FrCk6pOW
bs8+vEKypEfAhxxW7T0QivhENmA9/+Yrzp6zrXxCb+QL0YzdmzX4eotfuDYiphGZ
/1q6EcGQ9SAtk36CrzOkc1xBizxzCv4wkjzI8E6jXR8qNPXDWZSFjLRxQblqaJ4J
lZY9LYa2TJPQaljQ92j4ld/JNv+Cp/uNmy/kVfYnZT/S5xqtOdFjo+0Rd10HUGyi
r0uVooK7UXyr1SzfPLNeEg==
`protect END_PROTECTED
