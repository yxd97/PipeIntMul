`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LfsVxyAqZ9F+hPblZGXXzJfjYKcbYm23tCbPxpjzhUcX9oVQsTlMX1a0U5oQl9Zh
+6X0Na501YQAAarrsep0t2wfqwI92kSnnRGqgWthvf/qqDgp6ZWOy3OBA/Yd5FBF
Oyuv+IILHrI4RKK5UPk6MaAebrd/BN5q6xv83v2sh9+LZkB/ZGL0ReOuWIF8YdE1
mA7fK1+IzRSgbZFKN4DHOwoFECjhbaqqBW2zmlil6zcJUfyRxoKPPs8yZ9WJB00I
FsRzCKRlwIJL5pH8E66vgW50E+GCE5Td2ckHmyhtYyE=
`protect END_PROTECTED
