`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SMf2ijef05BwdbZQPYJYxKkgzL8r7qi7KQXMHg5k+FnTIc1gKz6jTlZdGCko3uUd
2VbT0jgs4IFSm2Yx1ziZ+jP0rlA0Nl4nxdO04HnwahPIUz0i+g8sjBRvYew9uEyk
FhNg7dEsFnnqBjpYWqMNi1TdnnGeXPCrj5nxLu2mM6XMH6cTkSe2cu5uy9yUHEPf
zm25iaw3ksApkikeUF1pLQDbdBaXVkpQGl+KsqZ7VZIBOoCUs+WN8WuAjizsuwoQ
442pCPuk5B6QtyigVpVmb+llKmZ0rP/nv3ZfD0aMvj1gaUzm5c07MdrOWjbf41Rb
OH5JnLoEHwyxPCETt2aT1AuilTOLyRdgku5yde4HtQTiTJyoPsfSuJ1zgmIH0m3b
C/yKlQBYSRDv/yCP9OdgqYGsOY8KWcAgWXZ/U3M6J7ad2wIBJ1V2eLUYFLE8LbXu
mOqL8Rbky+kKoUgCUtawQWbqKlnSOXiXE1GOKl+Dk1LqP/l5IYgtMLhdJR7abKOE
JEwyhsCxYqkvYKMzHMOPaKjjyRDEJuypH8h6IMJld67Rk0/csJfxIXJgZsXvvoUq
qkon5oeSM7QVvKHmP6wCQXfmcHfSpenkFqL4krK3GzsHuXBtx0/JdpF2aeaFl3e6
O913OJO6H2xYPbVNNDD0Knjh4C10jRbVInpzzkrYRXGTv/dj6DsDXEkKUG5l+7H/
J1/9Rys3+ooyyhl012XB/hosHkCwMlxc23PyFR3qMC3F0WKydZr0wSKsv2k+y4ZB
Aewu2iw7zvFC0DxL6ErRhGnYsaiDMi1qiK0h6fKryjJ0zsczc4rLsmWBnIyTMXHy
w3BtWFmoBQydWj7az+Bfk8R3mlm0m2F+cJ2nx1FS2xF5mB89bHBV+KXPRra5in5f
IrBQTBwxW71cUifztKKgClLJj4h1N48CaPMySsEALbr9HAa0O9ajAGEwE8BcxfZk
S4FKpzdqHKOYuLEtvpicZpUOFMAobaAm9ItFv037AYWh68sbSU7WhMrO1AVc3nsQ
+5+/cFGACuADsn7DO7EQYIABynr/xy2SMwiDIQk//ZJPYKvPldmUtabq4rgLCA67
AvP8LBvOz0NUZ/TdXD6nasDLSda1oojyVNDBTxfJZM/rJmGlpfwzCIrk21vJ5Mw4
5rxBvm4y8k1amWgpxLZABzgvqmtnvDXWWuKT9mMboA0ZVoB/nnqbqWN2eHe51SbI
8ubQ7PH/i0wbhiNzhIaLp4uEjrdAvz7dvqm+Sqbk7t7HyZSgbGtq3fPauYx1b5P0
1OQYfUuwuoKkORGzmMNl4TfgCuPZ+q7rdAvpzh0L2pxSV4CBQJyavT3Lit2RHxb4
P4G6Qscxh3TWJwKNXgwXs8OPAe/sc1Qn6hze233/LeXLPdVG//FtuBLEsSt8cKuk
smt7ycJ0I+Ac/90A1E+Zc4/nvtudAii34jOqTypW6Nnic4wrDrx6wBeDuP0UEbFv
VtebdcrA8owlmvL2f/2+Pt1nfNRpVitIYbq21sQgHcTGVP/Qh612l2laSz5GEAdr
2gn1woadikgX5NSqyldj24YaUYirlROBvjvTrg1SYtlQNOAdgAQiXF6hzFBZMmC7
JJYtrKQRldb2Y308IRdgJF/9WrG0bk9xRhZ431gU7M3ghSSh+b2M9Ea8POHsmliz
DjAsuyrPTEGcWrnREQt7FG2cuvV2maghYKXQ15+fqeqzzFhmW9R7+51mcNAF9Tl8
I3M7Kg8xBzrTxO5MqQrPtTEg6W+vUgWG3UaW+QVFxG/Oj/ynNb7C/SbiRIhnzXcQ
VHxEGWI1GAssrJPFvg/AbvNO5f1oY0m7toNC8RmN9UJO9BR6OeZZ2r83pY1NWPxL
boE3MviH2t+q+XI92/ldELmdChGAQuDHcA0gnA4hvFcaNuJkGAxo+4jS83r7Pp32
slUj2ufgBh+MZ80tSB5Y1MLcd7Ls8//P6Q7rFWD3Wgay7GgpP8WHaHijW41TYHEm
WiWGABTZrBFrDVxSzGZmZXdJQJnmLGgbKU19J0y6I14ND51/0kZpZS2gPUW6KTD1
htW2pAvZ+Efa+dDL6YPE89l3NPhFzPPt8mzJHUaMJYAKMiICeB50b1ux5V1B/0Eu
pjM5ryzUMqWWaUYa/jlm+8nyKDDmafYNCGGqCnZYZjNQrSy15MXf9o2sIt6R+NTh
1V1zGsPNcfa1EzRsd5LRRwp0HdECvyYVQKcLZ/p8n9K8I/pXMYvudojlCTdC3Qd/
m+VllVMH3nSYKLt/Q5M4fdHqnrtXWzUC/vi4I8R1a77TEjWf41p76IGYNMczGf0t
EnRd69pIZ4tDcJkdQPDsyR4/BqDJbWpWGJYDXtGEKHPVUvQAdYSOr83aaMl+C/+C
cpUWQzviGlc0n/3ELYVrQJfGBcJxvA8en+T03hdwS8onhnLHjTRrHzycDGySPIjB
JtD96Q5ZkkKREpfD+LSfFZ3xAzk9GJQ2IPrqx0iL6dTRDexVDk/nz/VGyUfO6xIJ
j8/cgaTaI/kQCC2pKiXayE1dm1G5yq4wS8gEU8Fcs7iOwyuhWIuvrq3GAcRv358J
HVsSxTZDMtUanMxEUG3sNtH8CR6cVcPxRd0nkakMnijge//pk7ffGW8yAJEezCFJ
dE5AX5oee1yIEosKf3gWStnWMk9HKgROPyj1Pnpt2ueScNJ+tOo9pKPGWYHzFZNH
5JgJVslhmfNoUZjFTim+8NlDaF75ujaY10bSvZR4KhAz3Q4BYYt3jDuA9oJSV1fH
HSTNan0HfJyKQnfN6eeZW1ULI6mQ34MvnarzM0boOe3mRFqNlXDxrnXejp/BgO4y
mwsrTk+EAiWW8/aXwsMsnjMDP2kH2LTfPSVZFePUUUDRRQ6zb+xN883T1jVc1d5o
oNziX2a6Lyb6r3ZNvQDmPgOjEKAoJVKneqc/9bWdqvciB2XawZpBS4OtRUwgqDs4
vziH3Qd+ZuH0NUZSYVZOfimONea4pn/iNjekfMIRLF+hiMEf+0U7QQ/9d0aYd4Ja
UvfEcKz/4B62a+ViIIK+xcf8IC+XRxEO5DusCxK9KH//Hrr8mHeoWjcihEe3/WE0
2pzdniU3QBXq8ffgY8RGMspf0/CTHV3hMb5IwojeRXTGf6FALvf7AZhERzVpDlok
pEDdGo1zng4WfV2/neQu4GOFQRMeblKVGMjqEGKgmPNP8Obs5ixY9dOKh/gJJMAz
6WH+c1QWq4Lz0jz6jZR0Hnp7o+KylDHrG3iTqEifHYemfjD+Sw77lT/xkLZyXX3h
I2WOprDwJo5eOiSDx7id64HgE85qQ62aDBPghk+jsN4Y2a4QjBIcDF6DW/8DvA8l
gqDdCyJRmovE14jAF4w/QDab7o8NwMq1C3yqeIuj436biqLiG1cw6VvZa/4PtNhP
zZeWNRgJN8VWrUvkpugGFUYBdEGK+RNH1/eFbYklAL8QSVIv6SO1TSgexU8FuStm
Ho/ZHOHnDANZ8IP2p8Qa4RBe1/qYFj4SEVMpQwaqY1Ks7KCzb+q4pvu4yE+fGaxT
e/Xi+PAjQZk4ADTPFxfbTawdsZbJ/GlIamgsb+CUjF8apioc8FhIMdrL5ddw2uD9
oFbMM9cLoHraU7hFx7OthR14f1mk12ncvd+meB/gEkKfMZYwEcCFGCZmbYOe/67/
YHzGF10sM3kmrX/7X7r4L13pHSc+w2PC7Cqm5RLTVP0=
`protect END_PROTECTED
