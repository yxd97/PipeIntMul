`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JBa8LULV56879dWuzvYSG9deZ9ZTEYKB3VhoEww1rrus6p3GZcsyYTKnyoMRl+51
NbnsMlBB6fVAKjQqwTcapYfm7IooqfGuvdEVDS5zxPiLJj5RJfIyIwYMa2/KzAEJ
IFyjBddq6mIcN2dEVoyVUphypkfDEPkz2xOQMuw/WuKAksOH1HRaAjKgz87L1lsg
8E8oN5to9LTnmHL9IZIOB4Yt0MxqjDOywGffAOcTeVbVaV4xbSeCVq/XhK/qA4Kh
diiIzgEbsyY0N4v+pdueKvWAyu6+YFJeIqxXoSYoeoTnAol0H5/OHLEjhv6GRrLP
g8HeIZO18oGdb0uvm9yj24Z4Pu3wj6waFiPlGWCmIeTmM5wu9rjYyhK6AvtvKYcu
Z4IqrL0eonIUxivUctBRGqdqNPoZpxKb/Dv69PIpV9Ao3+5GGQYfa0uJTn3B5877
pxwFNI8H2h0HZNk+nmd/7k9AaCPeLoaQhx/1djGzcjPkPP9dmqqcLRpd76bUNyxK
buC1ZRCKjcWl5cFjd2B4nU1HY2r7vvg6GfTNmoZW26j4IIzXaDxBhckhqohb2/Q7
yUxV+Fhx1PXHVMmSvuqgeBlaU/yrBBiUjeTV+ovCUJbqpqIyPUQu6vqcJPGAafnc
I2rw4vYR2ZgfTHNV27yYk9BWQPXr/JPiMo854QaQD42Xyp1JqEr5ZC8eZdgBovZX
Xj8mqCXFnz2QTHSeh1v/isRnDhp1HLtj01HS/0rpwQCNT8nv9Il0HPLsu5VIlHoI
oZENq4XNskTvgEtnIvgEqEcY0MhwLYQULthOp1uKVJ3SNVFkfrcQksPFWhYNkoHI
79CYndP0dW5+jQ7p9X74FjPNS7eNTj7fQgq7CDqFLjJpNrBJdbyMOtWMk5FdKpjI
OiJKxjJKzFDn1SVuw37yCxSAYwCO4DEHbelpYE4qborOZy4R+NoV4BXOlg7Y0BUU
Y62KEiNdby5fUpRMm9+rlkcgU0I/kXGAU6cs3mG+v4miEElxJAKU6hFP3T3DHKSL
xgYais6d8/C/hcouhCfceA==
`protect END_PROTECTED
