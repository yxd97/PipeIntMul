`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
09t1WjvibdPo27elqX1MpDmMmHCXnxBaXRvC9meTrt8hVaqdTiYI25/n5AO2FMcJ
8AgHLOCnfdyn6MV+gS1DFlzbR1+zUk3/OEhP3rKiHeQYZ4y3mYx7JD5lm/IC2aMF
SmAiBEd6TgJoVuIuxXGcdPsbEfiAQ51D/3wPzGhbS7JXloYhi/PUq1zFJE2UgLeo
bEYaxH7yY9hR7NHzgcIR/LHuLopYZPISTnIosl0BfV7y2q6KWRGHoyd+rHlq9GPW
CWU4sl9aGBBRsz6asBnqRUfeEqswChnG8k+LgCJJqXRmwXjBrtphR75IzFT/5uA4
UHCFgjfx4BgNUvNUUkMbH8gXHEOUI42Y+JkOnxS07oZPoVP+Y5lA/8nSbpD/90Db
sOTpb9K5ruqID+Rs7Xqd1K6iS5bTiu0enYAmf/Y7VKaSK6wS3ofHvI/dZt9nrKMq
jt19z4zAjPdh7FpeVKF5JDUNw5Z0pKJZlaCVEPG94dFxys4+8r+mRQzYtNhgViy6
BVxDsczU0ryFncNZpn3l/5XbElLwoGq6nmOTToUh02fpRDGKvyUZ6AOndbYrplKU
GmF/lTLM+jVMG4CorcApoKxPQ0y2VzNIUW6F+YSy6IE=
`protect END_PROTECTED
