`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jKLbpRN3tAP/Mgu+kCDAEblobscQq17BA7F26qggBx5frzbwaXqaWA0okw7tk5ML
Lgp04M7lrD9S5dk2tzxEGkmoS6pi5O3nB886vFYDqLhnB/bfUWJ9Adwa9UTOuTMO
MfgVNZKbaJOXTfah6qhl6sNLC0HpJaHGbXz8vWMparcGYPuUgtFGf2S0nCj69V84
B9sz/bGX9WJdx4O2ez3a4oD35f1vuClW1Y9tmudGfWrDQZZ2jVEJaRoY1WscxBi/
z8ouapc9f0qzvVTAOX8zi/Yy1fmLFAgYAVB1tXwVisHc1ornFDxODC9CbIWmBWgE
xZfhaaiml6UoLvA3yv6jKsTARBHprYMFC1Of0tDq69SfQeFsP/vmaDrUSXaqNGO0
iSXIgTStJUgwTDXf4eOCdHYSrxDttyGQIx87H8LP+CtTeJRe4xuu2jtUum5qr05k
srxSbskOi74Djmq19g7yJA==
`protect END_PROTECTED
