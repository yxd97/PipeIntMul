`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mL97qR0LPO/9XrbmyOz1q/KHTfIhLP0LBdKbShmFDs/oRpwynQe9A8ZHMESedzn3
1w0dueiJECTXtij/LEDu5gQX5pvLjQPacWXzWEh3BOirMEMWrpWLCfoM0q8nquW+
xPGNh6QWpztmc/Rh2yeJQu+vO+KOiYXykhRQvBuFC47qa0LYVBJXMW3rxmnIR7fo
a4gusuvL5A/toy0FkZAtI17yEzEqCfKJnbrvJOFETe0bLsCo7XTtftVS3JgO2+/K
PIaWYzOdBpk1Gt3pP2oCbgnjpIbs4zLhZeKdjrBOXu4=
`protect END_PROTECTED
