`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AP3BnTPuHyAZ650aVv88EWK2HP0m7qHhlF5e1BUZifkh6ORR1z3+T4+Cv5y/+W1a
5E+KIPHFQuOBaTF+lGmF5O8AO9rRi6nOn5s8RauFFPgl5P8lA7rgdGseLouPhuSS
uDRHio1LHDo18/bjmSPxKvDlGhnT8svT4/bm9LWul0BzMyWKvvzJrhrOY+qq3b6I
A/iPRUJ9plPida2yJ2duaZvJmuPWzTVhG89lv/s4X3VgXxr9AvEwVfOS2f1AGUTx
`protect END_PROTECTED
