`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eu1b0CpS839ks/0hxe+nHvZ84kJrNWcEKjL77YolW7RO6hJZHEtVtTww0/clwyWP
/S1KsK7X7YgO0tLl61RtKzZi8uGgCRuN916qKepRgze0OLLSnlhgXCc8z6eXS4F7
9//z5sD6R67nvJK4PGdS3MIe+pjyybL5CiLOZL6myq1W1ucykpNicz1Eq8WYjAvM
B8F14AnTWEhVUGKCCsDZlyJ+t0Gr+IWs78JoXyJF9dDj8hHHuFF3xNYUnPv3re9s
9/df6hqcTAJ46zd6hmcAOBQJ/V2lZAu9SxqMnIMdhHVoH6/7K6R4jjDyEB9dJr2Q
vF8ooQdHxFWsHvNv53TQdiw5KyrQsgqjEpxdVViS76ofG7xGn2aZ3FwOiut6gnHl
3Jfo0njK4sFIJWLtmEO2ZlkB7KyCa2Ph3Of39Fuud3tXbChoxs0BCH4wBMDdfiss
kipQOphBDUGgmIRsaJIiKXWqVzpscwOgXQTDEkOFplva7r8fPDUqTb9fUszOJuA4
tQUs8Pbh/FWCaqEG6UBRzwmcrCzpHghde1IlNhxQK1bbit0YYoIZdSVlpLQx1Pre
gVpg9YMBy0FJmEP1tOZsCrJ2fDdFG8OUiDsHGc5pQdFtT4igswHyI8h3ckR9qLQs
Nm7RHmE0lRouXZyJbA6OgoHAKZ6SvcA5SWh83rDQTUvvkPil+nIT7/5xIiGkHw+u
etAOAkFRTguFOh+/D54mrOpHDfOSe8eDTSuJmB2jbq87Ee+pQNuIDq/870eesm3i
lntR5PV6VIAi0s0zyuhfyZvOWFBw05Va0bZ972eAtREpkYrrVzxzz7RHVRqWKJ6D
IG8WCKqWpIfxXR7lYL6QGDn/LKm5lcykvpxECTrYUbMnadG1ZpivZ0WCH6/HNjks
lkogFb4mB1cauNEevCnz2ZKkRD3qLtIn8M/kzZND/M3XCFruQugbzk0lB01Tzeon
A5K8UJSnWN5z61xsEp5oyIx5SlGAZSDpmW9wQYU5ejsMjLFSQ/RfSszD87g5s5yb
SpONu8Bq4aVzZ08KiVI3aerYv4rgmMH0Xj0c0MiWoI46Qj+ADRaV8WkYgAo2Ie3Y
vDRZw1BlNtW1W2rV50QeFAaHEBbXc0H1EVHDmj+/SK7lZ2lhZQUjIqO4qJ75RnGY
8KcIr0KT0FesBJLWqxx9wKv63DkKVDz1PiGjxCLqaw5vkuNiiSBkUJNuEBfSvlid
wbJ1wd4rN6uiGFoX9d3v+4mglCAGpEtn2MIiOiP4PEXQW4fXuLlIECV78Utwig23
rAaudrTnPmHig5nI37Y3cKd74CD51LE2+Z3JsU6qGfcChE2Z99S6hmF8uBHEk4Ry
SVRQ2IehTXtGPmvR4cC/ePTuhvQp3zys8vFFIsrMyGQdLhVZsXeuoFD/dnmBz5Od
x+Sp+M1xcwbp7WfBzqLTsMUDLotdakEMLkfvxyHslF4TCzrKT5YqkMU66zPywh7g
DuNjzK5cOQI9G1GqGE/jXJV7GkRDgGO1ZyhDobdPOZWJVqisGchxT2otinlX+Cgz
hLHIPGk45X5XJ1rkYXSL5EDlVA000NaOl8Nk7bqKRqHIMhDFTJmjmh5yuUslsCnY
uU609T2vnafhLM813g/ztltUoj4DYI48JwXrY/wA5aIhAYzMrEGTSqKXftFHh64f
zbYUpA72AU5D+H5livgwf3qZtBv2pBAxESC8RlSlonOTpPV3QT69BcH9c7Un8jhT
5rjHdggLTyfh+Tkuqk/NR16Y2wWOgw4YHqhpBh9Gpi/L3zFTpsXWjQh4Ht7Epef/
yT+Wv8wMvYOilI866b8Vli5HcNfPYCn3OcS/zHSm/HxgSaatkTReBPqkNzYHnQ8e
1KyiR3lFmMDT/IIB5xondEtnfWG9/cPlCb1gPBgmwl8MSMwWPBVcmp+RYOVOLDlz
H6bIvfqpiwrHrOKbFT+eMyK9z4rWL8snkOSNGkLjIJsKY0OSkodV9e1oDeCAtQhP
ccMNcQK2VCG1xQX7Do/ZvW7TTggDY33c4xHw62KhVWl8313mdgUUq+diyiTpNkiG
18D4F20o6TRg4cBDFzNYWbpnjMzbkCeTtTJfUAx+Ns2umKJ+KKd0h3J9pDjm/jRI
GbMAJXnZLSmZ0o61EDIev80tGSQ6nKwX46Jo5BIYJ88UBAUYuI5zNQsTvDoahq8d
hZYuhLrQ0qOxhXdwZw/S/HNajZDaDgW83zsglcBrI3o1NnN2WuFAQASlBG6rnwWE
GrFvDYmNpSzd+V+4a9Ai55mkLWPWa+iutysw6REm/IH8U9zmGR1ZdoRI8g2tTdi7
q6+keKGi9nhrpAsyHuQjm1pwn5rJFxkjzdtyajkpwsZAOjeSTvStnx6uvE+IL8BR
8YWvtUWyo18ACBJ/E4z8Ea6XswtmEHkvBRHpgMsJUkgzme9w6B5QYsXE2Fa87MDX
No/jYT831KAUV4ReX6xoIaegF1oWptYqHR0zWJM1TEFIa754eqxgJDtaRVKPBvIj
X5nG5GqA0wSmiNuqIcbixLKq8l5sbnrLDDOx7WB75T74pH73E1UGmrVN5990p3XT
MmDe7ceVTSbrg/C0OFV9fBmZonM18HWHwmPdOW3amCqobbXlYWoA72IgfdCVOvI6
noqoGq/iUzsVC0kct88/puSoyUbJB5205BmLajqZMwlOoWVw8xSGLwjS4JsmnM7H
EeLLQD/vwWAVegxwtp4xw+w4KlwgpuB/uJteKb71iD61R9zKi4XcJIJRznnYbkDt
LNGcBKlb+K9TDRONzaIlCOhz2Clzk9sQaZLONdT9C0/cS0Lg5l92UC2JPCxEIgNC
/EziPV2AuXHNth9bqa4igimAJPuWdP9EiOdrlmWVDBkfcd/8pbpOblU2rl2WxH4S
WBJY4qft6k4hiOoY/MMyMTdvWzGA0duR6Fs/0S+NTMEXpfi6Hhf1VTR1oW1/y3RF
g0grAQw2rnNQa7rA9RqCetBXKq7PDy3rQWGVCY4PcldPVO4zWj3esxg/Le3UkKZF
gkemrgIqr7LD8TVwc96KPunZ435jDFCwevvXPbJJgEzEuOuI1W5J6PXKYWOsrdX8
YTW1drzP34D6HPccPSFeCO/EpRuIj6vNQohZzxhgMEJZdpFSy+mmyXzHxMmfZhlV
k3YlrTnEOGYTxBD9KaTnZKgFfyvgwwF/Q2fBGhPYOjVTJOzKBSI374W/x5bUK3Ug
ehLTdAvK5R3LOIZ9bPU0cFdVef/74LFt0uOEwmr+I8H7slRzpnK+lktF9mnLDo9Q
QN3JSRGochqVqno84395h75t+EoZH6CHqnQL5pUooVLVTkflPuIl+3FQj/uRGyXl
Wxx7SGLS7zNvneFiXGUFsoLPiLOwLDXMr0/A5ExMbRBVEIC1YgUpT9wh9MfHLs1F
v3fJ+flGDQpXANqPHnkcNzx1g0Qt63/qnP7L3mmVZXKGY9TQJZ/YgZE3ip/cmy6D
2KOLJlFdU6IfUqbvLg2jsV2hnDK761KZw6s0HnluVDB85Td+ZZ0unh21MtPxDcdd
U9yr2jhCkFIZG1Xj/A4IxPrvFmLuDdQLrpHNhlIn1QBgultd0iUpS6EeyLmPlJBg
MKl8k78HXS014rlwmCFUQ1VywMpT4Z68DVGXUPIsEtGJlbb9+dYVnDniZxByj1UI
+pJb3gnIol3daqQ+z2rhKERAxjSRRZIMqrItZOHSooA1vx0mtPnXHeOiHfCGJ+0c
suucRHzX6l9WnBW+FOmPyyVrofkG/c8V3fn8oXA7dHx8qZMcxjCnPhEGC/5zNnrh
tgFAveZYXaexByeVEIevo09TgP+78DKxXk6GtyJVqTd+1rkMTCuqQZt11YZFWE8Q
ky8AdC0p36Gcf56691hK6XAu4QJrnqLXT3+OcN0jTrNQdY1F430iehlDqSj0NMXV
+NF6zRdeynOHgP1UuyzC2QVx3CWtPbGgdm/2EJ9L3HrcMJDdRlDtTqkBDj34UhMT
3w2DnuvB941LwJoTZMZoPnkLkmG6azAbortl3RpBpB71vTU1ndAQSn8xKT3Gto64
jQCLBRb9SWgSELxU9hnsv9ndtl2WtpKYpjVBvm476KcPG+vMkfochRASyJ2BMfaB
+3Dnlb9vE9msOnuvXxX6AZEa0q+SGOyWBR5ONciBTjAZabFYk/sIDdy3hHLrN956
jeqjbAi9GrlhnpOzuobnJWYuS1hx0sAhVZcM9L4moLG81E57K9AWSr8lY0iDDdlx
R5lfsqxr4/JxMwBEJ9iFIEkUhlYu1mSD1zj5vbmosAIxneKXFHqAcxdbfEqONPh5
9tkfQxs7Qm2I+eqntHUabggrG8zfGGt90QDSx+V5BUfrhyjzytGns6LuFpe3B0P9
1j05uOnsI9JdXDdroHmhRZDFcBS8BmXFKRNGftgFrJD/9LRxuJCLgJjZTC40Fd1Y
JO9bUoEnNdfa9A2cpjxfyj1NiWRVSaqCsmBRbFE5tobkAjrLvXopTnHjyifzLy2z
9m8rCuvzXysWEqBe/vDSWTVU3eqr0ms3Qp1OydmbDvk3sIwtwlLlOleqVXx2pf3X
9N1ZWgbcfhvK6YPV9GlwRcYEbXZ7Ix/Dke7M3LZOgoPTtvKVWOH0WQwO0Mm4Tl6V
+9mn/ucIy9XTTBh0s1mb6a+cfWPQR4K3my+DFdFzhYG0ET4bHynBS6jXZgT5s7jM
vQTJfPEtSTGEPefGQQ/FhknNusMV5tcvbhiOev9c6C58LZbyIIi4dPiU+nngeC/e
bue5VkR3UGdn2bjRGCcYBmNCObKpefY2Lmizu1mqYbxsGReiTC1TKi0QeGhCYUSa
QLWM86v56TWB7WAhYf+imuuk8i64AX0HOJSBVNP2elpZWmYSili/HiBE9M5lUSoG
ljg56hfAu0VoBhz+qkeMWpp57X/REsc2caSas8B4ZN6CJ3HM0LDfGRzrV735aLzQ
0VSEtRSC5bhfRuPsGSeXT/2EceK/3qB/icuStQ/BesUCNyn39uBQGiNNSGexMmXN
VAsH46UDgOT1XsojVIlfXLvWY/CbHhPgC0NPvvTGiqtyYn3+x3ahVtcD1RU5d4Y1
Nyh5s8DXvPRdHH6o5HVL+r4UTFhoxyCf9z3pkyFjs129mjZLEYFqLHiSx5hfhNnY
6Ng6fnMa0OtWDLZGAwnGElif1gyCl7UEY/A8OjSHITgL9+9Utowq2QLTvzoYNgjU
p66fewXBHj/fefF9l+gk/cz4h9MGPUA1GnFE6A8DtXvdXJ+bAInLmiJFO/PhcRKP
w3UUjSjYsPinnUnUslqFlRBw2ffRWgCajtgVSykCOqq6hwGrCYTiM9xoUSdgmebA
rgcZmjFLDoRr71DN76UaayanWWrbBoxex6A54ilOfL/5lpvBaVoPwCG6PZXY0kLC
fufiEJFSCKvJQg4tBa0ct+K/zqhzf9bCYP8hgyj1i1qRUuwDQn/Cdj4v//TKc1dv
G3SHOc0LvzKq4xQE4IL2fFH6by7Ub7sOY2lK5LUw/knH8VuNeXbo64FPnRYY/s21
ZoCyiTxzaCkMwnGahg7yCrDtKql+thRQIRo4/MGEeT3Ibd3+E5gaH1zoLvK4wXWj
jiLFxQXU6u1F1oASz/8vcDX090gBd5pI7qyM320+Dk6J10h+2wpbJZedL5JZKOCz
McN1j5dKLbfxkuz2bnHvOQPBIuT3VyWL4rNgogFvxVpMNx+fACgwcMNTCXnu/y53
i5vuCLfEvwt6kT6DDtmF8RrdWu95aKYvhsVtGcjm/n6D/jilTpa/zBsb0a1OiW3H
Npa79vzodIv/jtnl8mjXnnQ1ZId/qsUFCE1p2vXi8cmHaXhd8JuROKY/CYOulzOc
rq2I4PHoP3drynb0u6FNOqHup0K5aa96NYAQc+sS1+ZJS21CxG7bJrXAGLUuX3Wf
c8NgeRNl2OwSVvc2tJTZumsPoyp0gLwbKbfUO8B2AIA3NcyKULegvs692c134T4E
69vLA2+7mlrT675+ZX2BtXbPcbwchMwRt+p3oSSFAOOAgzYLVE1LiZ5BH/hDRBcX
VrUwnFHINVUYw6IB8zkiKfdNmxsCfS7TY5lGztCOE+gEQRzIi2oROk2Sd/WDeAQF
N7RyDRRIqTwe4kJ4ZW9NIsWSER0I1lwdaYAQilKdRdW3QcMnL2kh2tKPTuWCqt9N
Tagim5Z9ANa5qJ03eRIZ2aUiiZq7HRdKasgO1LCBrsIOI4rPK9WIEyC6EJ4S+GMJ
EDpo9MDwxWTg8uEX1+VKh6hV19Aqpu5P9GWxO4KGGMKAk7KQMDtAF6PelhRIGqjQ
iW22tRqVtHw5XBeP2F2u6To/SBQYvv+Oh9WB3IRAT0zinxrxw9xgQhoczW59q58P
MVOb8n72lmhOsg6rmwfDJ3fyShFPmVJM3q3GF7pXz1zTHTAWib7q/52j3E+naOgk
fFf10YH6DXA6CxKPao2HeqapdP/7ljEpmMDg7DechvvVUWZdreUOvJz4UINIv72G
lKutPWXCFk2K/J33VhC36kaTXA8eAw6cYHAZZMAh2w5NpEBKoWXSGT+EcE5Q0BAF
EMsEYbfi79i4dl98Xt+GGsCU+wNbsh/JjhjzI2w/a9SK37nLH/FR09pELv9tjbLm
tmQ4wIId4BhCoQDdH/M/43vL8Fj2KbcOsv9tSevqZIDQuTyi7aoMCWhiw+JWZijr
HJt18QoUh3pV26qlyhSJGA1JQAql6HgDDBTYkhSGg/LH0aZJI+7PZYfHovH8WFJI
Oh+65kKAd20D5+Cj+Nv6jTatBqdJsjlDXK1mL8a3n3TLM+9dxFVHEsK/ap1beqks
DF+qLKa5ForalKgje6UwQF5kAK0Il6DmgfRUdFdCHsfPzcXGiYPF3tD2WK1BARbP
6nh9hZ0lIWVFG/zIAOuDGzp2IJckYmx7TCduUzW7/YNP5JLnGkY9hGBeEhwg4pHu
OHrpNYszbEO1ytggIg3/AuKwMRCzDfxu4uFqwMX5/yWcrdS4H4+Bq9dfydjqwBdQ
C0tZ8w3DV4h1leAMKbzGkw/s6IKoDmFbiiv3B45PdFaFQB+/vMLylAEAplqL+u4S
z1ya+0N0DRatHs+f8VKsEMObpKx4ebtLj+s3i86l4/Q6JLzWWuSRuhZRe20LXXmR
/HldWzrURLbnitMtuHwBnqYNplO8t/HWMEdIssmfAH7JyJg2hvZaeLoOhgqhvzTE
L8ZHXG8HYceALa03MD224gSavwOytmY4zIkWQksbFTCm+fP4XIao9O5tEEu1XAgE
ED0UZITvarfSBr7P89h6zRHmH9y+Kba6e88p/JkxIXPWE4eSSIZlIFIXBfzx7fxs
7y+3owmXEc4JbdBQ8h2BCyyDDRV5zcaz+VolFzk0QLi5uz/4YLFwpV+B03Af7dTU
kmll4oPhvqUJQgwWYOYMHMtje5PiOfyHdv836lrmjP4MIZDQLdl+DHFMtjPNS1y0
n7Uk+bzwMyNbl/KhThfJqAj6xdPFZ7NEYADA+tJOGE5AmODKfwEgwsLnKQVbFw8B
UOI20TEPhc9IDHRmJCgtIL/owbADbD3rnp196CfGLhEdCmEmx6u8yA071yBZ95jz
uZ26ZDvt380pT82ZG/UCd4tKabNKFScM2QmGY0jGEwTe4j2QQTnqD3JOlJrp6Xck
w0T+paxWnaD5cpk/gNtpcS8j8DEcunuZix9oN+s2GbN6jGMWRfgLXBQJN1YZJbjT
t3KubSofGG935CCq0lQ7LeVE21uy5pV28lqnpCHkoXcyzRFPXO6nhRZLVPqPLcjW
LGGDCIOFdNkKDi2SpjSoa1Tf8I5rjGHpPnxuybduvgmfy6HFg4durJP3CRhzdbIE
L2sq6Md6By5YrhL1B3/INrOjZNk1toVfu+adDuM2Lgm5X01lMbL+SpO5uER45Qg+
3giF/pylU5ifjI3P1Lcw/QjxNBjx6BU34MttwdctF/GhNTIt2kRJXqbU/qzJOIxf
ZaD7KH49XsmQJ5pMdtJUNvqW693YP2gowElPu2j/pQBs1TOChMCcxu4djSxv70ag
hQeROLVuiZYDCQIJj73KzuqXYVLG0x6rSdtpg4UieydpzL6h6I2AnmiJvZM4cwi3
JuV26dDPQ24Gz/b+1Y+KMzwmzOho/VHE3FsazyrJB/5DOb6q1Uq25eso3DGlSpnY
VaB41o9lmFpNCx8Hfg3hwI0Ks8hvEKTZcmVq+rukhqC2EaD3IJSQZPTzHFPbkibC
cF6dx6D5TRGacNO3nMbHBQsvDJSbO5t9pF+vvAeRx8Ifiw+NPXHbC/oPqIMSi9UM
EbokpIVK2/GwslTZWy7IV/Mr2Hlqvz/2y79AXElpQQACvRYyH7gsgLkByNim60QM
c6gQHyuUMeBbfaehsq8kmwgkUX8bTXqDkafAX93nv+zcfSXgbm2/Ris0mzJfzOWa
ymECChn93ZkfRwd7z2Qb9AbyS/lPxLgAsEBCEfBZr3SbdW8t7x2rbd7FsOtQDhIz
EALqo0uX5SotJ+rI3IVE7FjOHScOlBhvaKncycCDprwR2ce+TFUJI2OUy7gM05yb
qGV9+qrp67PezzTjbW5ETTFbOz4cQB5s2T424lwd7VS6F5Gp17oLDnqPhkk3lpSa
ccmfZNAfNtZv7BkIv7509Hl8y0U4/hRYT/Q/i8RoB7Axmt+0s1hfTzabENN50H4H
34b7xPcl6sIEQJ1X7URfYQDM5YJg+U0WV7YvkKKav40=
`protect END_PROTECTED
