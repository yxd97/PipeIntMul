`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwS8dKtmIymrCb5g3Q41Ps1y90v1Pb3gAuGnB1vGuH068k3Xxp8K/jB6uzcWNpm0
FCfdzG0tqqF64R4GVTbMvLDg9k8NrG6k4JA1NjQimKRNFAd3BYjn8zL5XS1g2R9t
f00aW4MrgL3TV+pMg2wDv8mfloL3mflj4egZ51SH7t/3HugzMExjOcJ4RzmjSKZZ
rr41R5Mk960c2BZf6ee6pp3w+tA+hjWMYYtEnG3ELY0aPmLH2RXhLQ0UZVw4dxHN
VoYCD1ScO6D7MfCxr1151vMkDrKlLFFnQUootdJZcwrEBad/KiNqyCDIFoPPeMDD
Lwytq7lsJ6ez4huWjeiwz6Ezq7759ebpVsgPltgeRAAlxBhP+mueakMjGQhU1PDb
xTG+PrKJwaiMDs7ZN9IFQv26Dmb3RWZw5PfuHb2yLQI=
`protect END_PROTECTED
