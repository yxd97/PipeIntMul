`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H/niwKfQ3GB5DVNVeqt65Qbxctr+iwjbvmApm39W3Ri4RYI1ZUIzJ2zQaFdt1pm2
lXMeqPAtWwSqdOjnHw71U1HQDMCbuzUD2BPGZMg+SvWd87SIIhjHQPToD66s7/Fu
wg39CLKCeFKDnRgHxBcMQZtQUcFnQcmcLQIKjLKm6lIYoRjnfjXd1BAEXfU9jBms
mkzrROGV/RuZMa2h8Z2yOzueU54WHzwunuFV4Cf9UyHy0irPoGV53/aLJW1NfgQw
JnOLLyE4DcF4x0ScCcI0OkbOWnn0wL9c1Y7hxYfHBRZ/q0j3BGceaDlsLqHLBg8N
sCpkpyWA522qLdzwx7iNrQSBNj6vXSBV8yEkB6bk+UtHODBcdd2h5pcu8delrK2n
qZiwORkG9If56xTYUHaEluSAUu6moZSW4fSI5nJ1JUbTOwmgh9N4sKOyrq0Dr47O
g8h4DmB5BL7RgPqEKN+Dtmgxq69aLx7MQFKdIvwgAV8qEHqzgY/RhQvxUG9D1+v6
6FT4PLh98/1Plr+UEj1KOuvbZhkUPXcDZnZSAEaHd9zseNi5+ZsRYgzHM99zliBA
Q3Xg8d/z221OP4F6sjeiQHNl+WwvPj42IaDVrwRXbDBXLDjDY6/9DmXvv5b9tSmf
nZPLzsdwnhOH5muDyArtGq7QWhPJkHtHI0kVYkDMdt1JT/ozAu2jz4QIDgJ00lOx
gyW6J8vGO65BRobABaLDLLMfoI7ud/Fqv/myQGgzX6T5UhTMrb4+eQPN5ApCoYlJ
kNfbLKV9uFjdgKT5sQSqTDpMZEg3R/tJVV3oLhzdclnzVeRKFdm5Ul1c6QcS7JAU
GVnBjWV7ZWEhXCnBW50DHmFKKLIE0DIJR2DlBIs/hHPTrCIyl9E53ZwdVeJMpayb
YHPSjPrbsMtJigme+ftwPlpjtBJNTlLT6tLc7ZmanjrFQHt2omsHce+ULT/OMuvR
/Se6f4YET9oT5mrJkFHSr3e4eSywbP0Cr7EO91lj7LFKJkUM508HYRoc7Vk3ZCXW
C618wfq6cJlvuCX4iOWaSwRsJtgNaQhVdda2BaMam2o7K9X4VKI5PUr3nGo9ts7p
IvbiOI3xC0K+lRivG8TIiY7HJ5ZqSAXmIHzopb4XUwqsaEPRAw7p8YmPAz1dkLnt
af/S7ALhauGDVLncQoUkXyOydoLRBAD9Odt97/JkCzy/36N2QYauY6R+3MyeMXsi
JoGc+7H20vVFqe7w1adSROXHk0osOzHZxdq8IFXzT7dFRvuKQILp8Dye1p7lJmtj
`protect END_PROTECTED
