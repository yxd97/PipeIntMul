`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kqoi2/mZH81PJtNoqeokTgURMo64ZhmxIJ0vW3aryV0uwd7dozF9Ydld2bW+Ss6
QHQ936qL1xi4Dy5JSds3q02LSyEBL8FpoIizXPUAryf40pPgRh+w5QEr3MDxZjJI
YOE2alqC/HcIcnLg6ydtpGbg4xWdx5lZ/AU+e/oyH+1smKkBQpm8RecvFpnI6eyN
aI2yMPQlf9WtRq9+XE8Dric8uttLMZhL0+JT9t9f81smBR5CbeS/UBxUaZAT2NxV
/Y2yGeZ+k/CTtdGLnwTXb8XCzD4bBCYB72gVZB/c7bYRvptwdY6dPzql1Yem46wu
SV1i5LLQ7OVU1XLVp6Dr3wl1Z+1389CcCYlOtu+9OhNthCiW9pXHH1C7yFMCvX4I
ZV+xcvkFPXdhqzoA3U3RxdvHknxKVftf0vrEeKgHzfs=
`protect END_PROTECTED
