`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hbfSnK9uF1Di0J1wgFL6B6yoj8tUMXJYdBtFyVxF561tkQg9JD9JcJv+LUOTc5r
4Z14RTyi4DcYhf84gRgMIHUkPqGuwxm47Sa3lMaTZPC6z265+kx7CIneO6mCrftJ
PPwuI49LkLHmN74CoWvCHWGSW6szf02iahNIDaR+vvG2gPGj83R/tPe2h+DNwobP
0IdCs7pwtCAimCym/zBXrHh16LXtrC6qI/i36hx0O9eOZffDrw2CV7dkPSeLlJgr
Rbp9GaqEwkzEltJJB9LML/1dKtmK998VrYwqvFBlZIS2K9SmpCb+gbeLF2A/9mbJ
Pbk4Aa5bit7NBaroxiP2odKGmMi4ixxjBRGOfQ0e2dP56TiU0QqwBD/rw+/W0DI5
PR56OuPg5in+9wlmencRy6IkS5kc0mGX6cnu7/u6PNpZgXV/GE0h1t5ZCkwTKhQk
7lAwPO+eafzVQzBorBvBUx8jAszThZtClDoCHuIjBNKJSE2XF3UThKgeBuK/AhpE
yH107pacCB5rBMWCI2oQTsnxrZz3uQssUurgSIFr6ARyIrBfwrQI1tw35ZiuYlne
SzTWQNignhCnRytUuukMnQ5/8E4/SPQ3cGPystFFBhibocs9i9z646oX03gDijOe
Z5+uh7jQqYeuBhFCvf96VRrrLPbiaN1yiZjBj5dWRyFq6b4N7BsofysSlE0N8VyP
kZL5SegunZsFtQ8/rcSBg4rRRjd4LLSovUBn4tb/N7UK9qnowmWfsLjFQ+4oDfBU
JRglA6RU9x7qjjZ+1V44F9xYS3eAbreRkTUOecc3CnPEZl1ruqT3kskGKBgHXnBJ
Q+th6EhXz11eLPat/aB++bdQApQOB9WRXfX5Zjqu/OfdsYsC+1g5ownH/CnqO9HF
rbw/4gpbG6vfwgExOjYlq0GtSXx0mKt9TJvPkkq3Sz5xk1k68zMSPf+4P5S1Hs6K
VnKmcHgB3qLZlOW7GsI0WOajc3uGnuM57/TMcAVzJd8cRrbeESqkxYq3AnYfPlI6
uUSbmbxuTMnZtHwtZNq9FRbsqsVGcKckzORBWpC0mpVrApstQPBxkjhgXeFCbLgI
qy+z5TwL3yKAnMCEXflNP+v1AgIMJIiGOogLPrIpa0UZw6Unsy4jW3Cx+xqpeHOi
/VVIMclcqF1tw8lXnCbk4AqmD9hVi2y5r/s15YpKZZmejeMaZzi7k3ObV+0XR0a8
qc9PzJMyI/x4GWZq1Ab2bhBkTqg72HnS4LGBsR9cBYA6tWLHBTUkqZdsQVJs6A3P
uoWJ5eai3TYZEFfykU0mybJ/Rz47ne5f0DLIH8mYtFNYn1ZTo1lLa6tvJqo6m/tW
21CtVDvWL2EAXawWrLHJG1eLYXgBUXOe8oTFBX35dS+miduS6giOXjcavfp6LNra
7Y4xIZX9OIFX6ztrhtHpWZvoRlbAQl1EdyA0M6LmMwKPDVO9+ck0NhEaLJ/J8767
mjKCt4pfdLrZoGijkMTF177GkFlJZ3kN2HJT6jqR0UbuU6VwJN1TrXmHOxRj2gkX
UwvXKgq3rTAcL4qnIr0nlVFmoYN6cM+Nw2yHdWCgS9QbBCYYejlI9jY/DOTJgaDO
cGYXvwhXDyZnBTowR01N1ztCe44P/c0rxxRLYOHI8VXnCTURmyenMp37e9q1Yl5Z
8pRO69LdAVMq0vm3OHpYC0G9uyZyJChuvDbHdvQM6me5GgUBHdKPzR9M7kI/GncS
sCnAOCyKFv962ZBrz4Y+9xHudP0Uv9pCO3n/kvi4utT0x4ANkYBApKevAIP53q83
Iz7NEeBjEYEiyeG4LvQCRWxTcG5qaJ1BF+8IrPWqatpg7gmKuiHd/IRPg31i6qt2
EAFkP++E8FcrtTVs1vkXcas5RtkdRTU1eJdRIZJLJJvREf91dk8Ody2qSIUjEoJx
nd1f4YSpHQgKMxBA0kdb02K4a/OX3YFVT+Q1gX1Gd9dsFMYNumFOQ5HdtQisq30U
uMx5IBcTuxRPYy1SU5DjXO355cG/eMvv8Vldqxalvm59yfQRhzubPPvYmNycT/ah
s5wnbyZQns5xWvTLcp3cZuNcSftQN38KD+G9NcAc1a1bSRiuXIw+B3pw7BaJSSSd
gs6U4XC8CVENvNkx94z+JRlVlnycPahx2+4Gx0P5qCvuAdVc3FXVJBXK5k26lIA9
DlJHdf8iaOnl5H7rOGm49F0/0qTH6+cTDh2t1sp4WLOdImm40BJomMku9eQRu4Yp
GcWZv6wKMMC8p/7D7fJeR3PI5ePY7kwuqe4ho2+Jvv50PuvqidIjDYR4nP4KkWSn
e3mgCLB30EbDYzTv75UvXQsUC8+L/bVfKvTYdoaxU9OOBnu7l13AdEcsP14GY3mC
HqZNE03hxSHqMGMEtnJZuJ6HRqvFwHV7T89t8BJQLMvUyVf0kPPSGsRa+7LcVUmd
e1YS4t+GhC3p/5WmqR0RQYLfzX9FK5hEMYK81vct4IVTP2/lIZq5AB9hAK3Eaexq
1blzedzyKWoJsbVjqEMHKaqLxitd8UYVfjLQnlgaK8pgb60AtLLLUZrRFJAglrEf
wLuZR+gn+OvwQkl99cDvsc6D7x5c/2ZRm62XyYHw8vzzcxCuzOqoiC62568tnYVd
4ym6RIduvViu3BsFfOomGNI6RThqQZA7C/UxL/W5tNDA3/aZvJyagOOcKmYvSE6w
bUJHWEpmDWWA/290L0j6oTVcYLJEVw0CJeWLo/gfWq/w+hKGh4jjJygKnSZy5cwr
mV9H1cETwRvXTruKJAu+mdx8kGLRAxDICkKQYv8wEuARgX4FWlaUQrJKNy/H9MXZ
DCw+N0tMDaOkWwlkxhntEHZ+vaTHuU+rY9cGQqBMxGKgADnqiMJVHJdlu/G2XhK6
NIbkTk9nqVPuBydJuGKIBtSY1sophgoyCNehO7MaNn7PzhLMneoR3uF7uhZ5U6q0
IbQUys3PlH/POOmPWyru03vUdKHo9/20znvmQbwiCdD8t/l53DhQV6/jtXwGW6kR
GqSUb/8uidVwJ/lIQU6iAUxNS1wNk9wb5j7ueWGb0iPb+j5gdLFMZ89BC9Ump0/9
6ILMoaYYw9Pig3VXrMSkbsSUHZxdfuxc37WCUo1kZi7Zn+tCw+9COypYm1KKJcP9
5EWA3r0+tP2X7oCjwYVQVZEv9k5j7qv9QOEiY/jkUp79ZxHu6e4+f+9Bft+brfWE
2WipUTZaA0Mc9PJ8HdpOZ//WDH2LkGeJLqpqOayXj7obpsT6exQxw8juALndUBIp
PQdplec5p8S3/dS36MjVsb4IX8P+3kiQ9AJUHGL1RrCUa0P3sNG9qyQ9NcVe1pl4
r3M491J+UmWXKBlJiYqqw4ts5Z2mRYCF+Qgz0aU/CxUghk10hSd6oS18/lShdzHf
J4HimVxLwaIZmBd+Icpe7erZiseD9mi80cGQMMUU/hIkcCdOLeWO+dYH7p+FWDuc
5KdoPlCCmVs06J5aaxLOTnendGJmOQKRNGKzuPxiExGTpBP4FnTvU8e960fWr5t+
yCaNP18o7rbFAlk4VV91XcBI4cVoQdOEtxxlYXPAb+MrzspSDWMcKT12MWIlxDN6
jAwh5eEotV/rYeip8g07n9daNzUXjhkBqt1Jamk75jG9YXywGX8EZF8vEtI84frI
WU8PPazqnqbkZJ7+OwYH7dj3tpyUF27OZ7xp1RE9sZHOzvhDOTL0ZMkg1ziATd6q
GhnBo4uo5T/0oZM8DYFTeqi1wDZFrAnAExDS/kIWhe1+hlwbkXM/oI2/2nIiiRy1
UHWKHlpzVA7xa4qs592ZnNUC3L4c+Cdxi8Nz8KyNHqMySDTmiuC28J2Ha1tTQIFg
vtWSSomm9ZPNlac3HN6+Un0HIa+d0crQrUKg+kCD65mKV0gW+JttuEkEaDmlw2m5
KTb8EK6m4QvkopUHikA9GZwPZqZY9ImGprM+98lkSN4+raVnbB7AilHUQwc28o+o
rs1a8znTgKucb+4d4F3SxdEI953ojB1gizGVIxZDOIlvLhNaWON9BhxXdhkiUc2T
Dd5sWbUfaR9BRFjEetGU04St7+j4gvAsIrl3nEScsctP0o8S7FL9P8KQFiPPTOCi
PqA+Meizx4NhvfcWbLddzhuVtC8WuyYsDOWS8xzAN9J0w+bmlsNq7XJF0HSpGR62
yuZZftBKBy0VH/FJZlxXRrHBIJBbXrfSGxLm/Ekf5db002jGb/1HRYy64HLYsONz
oskE8z38zoPuO7Rp0Edz8Vr8SAgbBpY9OH0VA3QcH1Vw1DVjJmq+tajh0S2Id8FR
Jcs+rcqeedTq8PySS+0nWGhL8QH9chtBnjgVFjFWxy62/ruNQlEm44MruVr1gl/c
TJh3IXxXuhrnSkO9ouXpWFuFeoRiUUGecEtO5ZgvSv/QY9D9JT/f7YI0cEUeT3HP
d1VH7t7u6Vx0tyQInG2jMXvl4jb+hBESp7UCZTPJABXNpktJ4yMvTdhWsRNT/685
ygwYiuRYJWauGJhZ+AFh1uYo0k94TmsOGrVLl6CCCEzjgObE2giGrkri+Y4wW1eP
9nJry/641nL3KXhX6kGtzTj7NUorcI3GkWcw2nnFFR7nZELyxysSPHVwgJVgFa2k
lHLMjkgKIs1POiRY0ho4yVOAm4tcmmYPj1S3RCFGdbHhs0oI+PQTy7bH9S0Y+6+O
U3iRFa4QWx1U10ucP4gnK64zi0PZUzGKwsESQgXlxSqEM2gE+qjElKpRxnwAFgaG
jtdMhmK3IQ6Vx8jdNzGfKxznrE95ISGfObWxx+jE3ahV47fVaZpmmLqfV7pULfIT
DE6rCIbuGICPnCn23EqbJMUH4pJZ4l/yyIxpKAxV8wppiTa58pL2sezTGpl49Jc3
hlwET9akmRHygnLc3zJpYjbgdhu1fdyHT/sCUOWdnARfT8deKZat/deDoiv0yXx0
P4FQ2zt4fPXsoqTwEKEYqcQfY+4S+SpRZHTWo0dVpj4T2D7jM7lP3V1hqDc2WgBV
0UNAQA/HoJUOPlAIFGmLmWaH+xUAVW+0oD+LnmaCw+1AFCHydrOBP10qGwULprvz
AEzZpgoRGkemrx0SgKCiCe1vmO4JKpbtWckADnZ5pU9jPvY9oj3x9EAUix+YJDs3
Ze0KF98Dx1cU3+YibHn2BFasX7WUXlY3hcM6f00cfP4phiD6Kjd3PfFGle8qrFQT
Qqf8fkEiIbAwN1X6aOWUsCu6sTN/uuhzuj+B2iwJo3sRimikdQ7i4wl4pa2+Kzeh
O3da0QHtbZmIS/1vqRifc/xPuUGcxuLp0bp7kEt2peWW8pDDCKgOqP5LYdId517u
LaUuSqGrsg4ahSwR+TyO+0so0zYICkaj2VAHwVIXaQ5Y4MJ1oFkb3aoVEolJi16g
K6Ad/EwaysMkbwGPbI+Wxjtuy36KM+Bjxlv1xmzyAdBh7lsF0xqzD771jjxGkQdz
S6xuH5MGgJXAS0AuD+TVPjhpeTnlgNtCQIp9Jr0WAdDYIaCiTxFJcium9FtfzYeP
qcw6F7U9Tc7VOYQM1IE1RzIV3WEbD2+ghjZRsso8Tzr7es1VAowD1SABI5ayH2xM
PaiIkRufgsZm0+B2QvMp2X5Dv/083a8d5nnfKDPTP0mEjy8VnVF70J7C4479wKJa
MMhi70QEgckGyABlTQUJ2A7cGqNQQe9rI3ukd6ToUM57vzD8v6Z4shnkMRjJM2ms
CmP9l/J+B26b48c7/ZsK/fO/XhR6t2Dw2ruiDriMQpVM2kqQsfF2HpsxDQGU22L2
XtFQQ8lhzD/Gpqo2Y/l34WXI/KccITzYErTm6fkkgYvWvqrc/QQVKsMV6uT22nNP
KBO/MAeCJdXOP3cy3CC576JxDzj7UIPUe02w6CE10WBj4YgnJA2T4f9da7KUPy5U
KUON/nmFUyST6747OWMR2rwpwQS3kX2KU7mc8OPQb6znT3N/ObuY8Utd3nxjrCUq
Rh8wBdr39AcTfTnAUnkTiWbPWJnTBiYD/oOafLVAtfRQxG0IzGs+Na3EDdhBceN+
8NZMEh8ft2gew6TDasAXM0IUOC2ODzE57mJzzuUT7AbiaVFkuZ/DCOPIDRNlFdpq
0YOeAeXg40qaxI5IrHLyEARrCux9jtn1/Ng2RRnfWYnPEaZfmGwHp0OV7A9IJSKG
JjzvLbzoipVM6x7B0OkVUdH0MtnTxkaBc0xYLo87HpY60o4Ab/+PbFJBSyjW5Uk0
EgqfcXcbuyDUuJCMMaJnK51JTXve4er6FvL3ZPgWMkyIi6ZeOAIdC2NEXD8hVCvV
qfvAs2GTDoxnPEq8pHL5+hNCONCCyMa2KsHlVnbvhcAg7FMvNKIWFBe8oln/yl0O
jWBWgo77VXAxCPaL/zJ9gfuAtcTQ5NC1rRyl9ip2xSkQu3HvFnNWI/H9yqHMQ9fg
hZK+D7S9+PjWl5j8EC3GtS4J3hwlDJeljGxSuDMnDG4JWuBBB26s1OXzezclXTOa
xmbTlyUv1yKsYXvYUpU8QZ9OTuMDDB7qVeZhHMLT7MSXl4L+elDzJUcC76qHMmB3
JgmujjoOjOF6TPfqoAhnGKCNE0odBlTETAMSGrbhCUYKXcXR9G2GT0DRrIJ9LybD
fKwrZBpTdFJb/cVOjKxeFy5hU/8FRzRsIRCc9y93T68T5SJRVMvOBFJEluyU5R6S
ikNtSRDF6x5tbcuxR1PWhf40duoys5uDS88WQ81/Jn2rGTXzThAY8PWPqQ11TexN
xlJf001v7tShAVSLkFZ1A5NCdEulaNa1LS6yDvDd1NDOMeAPPZgAgoYpZ1s3Amgx
wtAPLj2gEDDx+RrnUY0hcIKmG2kOmKLT6Jfqn0zRrORu8MWKrFM1GIPpYvH3je0q
8/1bO/rDrLfz2CzRkSKyIGnXdzWhshrYSJJVAMHl1uaRBsSYak48IGYJGrFTMNUy
Wo6feVN5IYDLK4k1KGB/cGEQeRvHZPjyLZd7eD1nCcx5jAl2W6LbUBgD/AZWvVzS
dqoBsA808LwLVp8CcK9RU6rwWHv+CSN1xJ8ZfN+1Si9qtMuVEc/+5wqdgmU1ENvz
sZ+OHzfgxseFf5NhYUma+MgS1hDDZbM+vSiFck/UVPDopO2cS0Uz67aeGPiOPrtz
aVPTwq3MAd13zCS7+rxxzjvMsPqmhpTW5divDXrWOm/rulO1X0iQS5PmemYW8173
nrxJ44FLwNvZ+DHPmRg3rwMD9zM1UOaDocYrb8MSgmMcehIxZmhxxZzZeIvyP534
ePOeVANgGHaX63HmsneJ/253qO2ErL3pYtRyR0iwCZlR1rWZ1Dx8ARHf5EJX3gF1
+F5N+8tA4xmwIWbLMjQlwuxPoO02EBq1kNjtqXw+HVaYAMbV76Igs9K7KzFvfLfm
qpu5azl3a8lepFMjZRy4zDTptzWKnf474M3y3IHyBzTc2yURCG1f3gTy2KYM1u6C
cVwItoiyfgEet4DM7gHytpTU1zHl7Kp0Bcvn3fOsixDjO0ycxKx0xO5oV5z0HPrV
TAgSs1HYYqTKZ78/bkUpr3LmJxqMn7/hTLRWkv/qKtnZxASYKjnMKEGYsNUtB60W
M8Nw9VCQEUIUkqzbtSa6gIKRoGzR0DvJU3C1J94sQn+rN8W62zrxzCmz9cbFfbm+
FmyPkOf2Paon/b5hThdk/vSqiQFZJKvbu/DWCLY1h9iv6K79UpKsKtqNO+16R4VN
8N0BHcNQ7CMhLucJxcCuTUPZ081QDPJRVZfA/7ahIIfySHBR0J6iw/5bV/Us/D2Q
ce8a1m+jbOPisZP2UKVqu0VAHD60IcvNm4Ze18ytOKFZZyEZiUFLvdKrGwXvn2mB
zCdL/pP0SHW09Ds6cMU0vHrZfjjQEBHxwxlVeB2zGSqBkGVUK4ZjAIRZBmor/dGd
HilYBtggYL63PGsQr7KtBjYa2p38xBsJq6j0shWdSzoILvtJEyjbl4IxiQH6QBoL
7QO76om3N2+8MuzqvuTG6htlClAjXWJVDEBBqeMN645YPbjjOIoiEufTyr923RQe
xVimMujs20pj4XZBVDmTcmWbzubmRBh11ETD5pR77nWlZAZjuJIQIj8BG+z/0cdr
mtT8jkMrqYIC7XsAf20mlwr/DbSvf/z7zomou/TZIRlLR7tBblmVBIfqFIYe35O3
Q2rVR7EmwFapijfb3AL6Qlovu6SK+knsAbLMEgvjua8O/9xp9cdMcwWIWEiHTTgm
oF3+EPpCuM+kgE4d/CQbmsBJ10uUjUMDWG137ngRmd7OM7U/uXUZ3vbv2Uk9ubsI
2qj6iUby7cLPKyf/Gf88eqiRkiKyT/dPe+fzZObYRA42JgBLDAnxNd0y//96dtMx
R/2e1/YaxKrmJ0S4Ao+fLJeJ+y+xVbmgt6F9smbjoFFPpuGuv510gjHj6x0VmnO0
bl8F3AFNe7bEh+LYPEOi4j+7j4QYpwOXkASMjo9L+z6JprkhDhUiwM/2iEvK9zFU
qyNrh5JsAksiyX9xmDq58lGOq2PC2SQIf31IpC1uWJwG6RrDXCGkw5FSNKZyDm47
BUMXhOXH/OE4ywqNjqwP9i7DlUsvCsF6jP41VXk+psI52DcMimuXwQjq6w0oniyC
YdRq3dZsCuz09y2Zk4U+wJ548KLYO90Nmp407BBB+2iuD6UwZk7xdMPw28UD4nI9
KjdLLziGwQ7rpc/yvoVNFcQKPMk7khuDbKBZz8Zo2prBqUdYDEgyeGfCBtndXpEl
BGtUTDE8+oZMKz9XB6WgkCGKJtMvZi+DW9wbTmRuzM/yiCh0bb8H0q3g6USmKhZv
Tb2FQvUoEedT2TwkyGyFxGh2V5fccRDTGg+L8EH7bleqigbxoc5BcNAv8LA2VNch
M3RDusBhGMDKgcNbPhsbsz5DzbVc3CcGV/IMr1SvO898H+KC3Y1BaCihWFYQlaQC
KXoXSqysS4fiFQkTbslhaT/b3O46Bl+qr3J2aCMXwTycozmhNued0GwP07I2zua5
6zp4P2/IetNchuQ8CNCCIiKqoFEaBHXuENTC7YFCPudRWakiL+qHvmzB9kvCo2Se
HWH7KMhdKY0G8sFTPbcVfosdcX2BBi+cIiJA7G5s9Yr/B/5CrmqgP0bnSpD3UTCd
8ChUFhUb1q0K9OR5xA24eNC+cKpB9gkwGvBfQ2pWWH4TGwVGeOjNNtdG+KkTqgpi
RAHPkEftRDGmh2Qdawoq5G3VJ0/ByMyGJPqdcB+MpADfYW47v+2x+XW50NoAABAZ
RtSIiPaMPlFNTLkOwbI/1pltdSl3UOQgbAH3cWR+I8FTfBOkHMdqytGrrdx7FO+F
SIddIOmgjCHpDTjT98Ck0fIG9z+7fANtibEixeFhcADeok2/KSu7FIwF/UwbZKu3
hCm0GdyhDUlWtgZJiRcYiZ9xAianBYS8x2UWd83vWbTvRcwSvHBiCQl6t1/FdWR2
hm/dNvCkV41SX0lwM0PIKECNPJS/H8QIlHs3Lq+iP8EKnj8B7Et7+o/u4tpRTITq
2Jz4sPWQDjD3hNzIZdenUJ42E+1BDisv2AvV7WO9fIEJgT72Jmo2XKKkt1+kJKBc
7EvPs0JY5ZlDr0q/N9YsPnCkjQyOrQJl31tX4gJa2T3JDyOF/d2uZuYn7pN79K76
qU3JkYlxNu7dFlYkLBg0e3Pou/UpCx47DQvJYleEwUdFaBanqxmCzJzXy62/E3m3
FK3PK5XJw/1rz7xd8kdsMpMe5zAQ3BOS5/Jxvl9hvSRD/Voo9gn3cuN5QzX4n7ec
YRGACNuChGo0NZlOeqbYmo88tvmTdVPVaLFnDciMyZSvHwF9gWNUlLeY1Witi6Cz
1H+Oa0DSGhOLN+xm/ayLn3HeRD3iC9DHgOX5TjCAnBe/XgbMD3fCmxDjPC9GkQty
t0Q0lYW6Tgqjic2APTe2zU5VFriNMt7ZFz0rynpDa75MKmWZQeeGoNLQyGjf49cB
9YUy5Xbq/LPpjZuwCDTiTj0/64d1d83ACxkBd4kJ8WAfZ3XdHX45iZvxHK/Mh/Kr
ZFKs8u9EHZxfMWJZhR25ctlc6GjXuZ28ap9aZAVxDSU5UIU6pcdLIdP3xS1F4S2I
YZ700G1TdotH0QBU49lkepkGjBsjGJaNofV+Y0DkI/bcZ00jS8unWGnDYOTvS46O
HRuiJev6ORqorK/JGBeTWRwTWog0G7jXM5+dftR5FQaudAATSQ0gRZnjQt9kvgF2
W4loVcvZwAFZNdgQDoA2ymLePVt2Up9dViHICahbvUDM//DF8ekCsmnF2qNTKrKF
Ft7iz3n0JLxBOBeivtjt/yKAfuYzSnHPbrkNvltID4J7/AKo5BEYg/FLmG+i8nW8
x4zQWNh5urYC5rjK80o68NnQBUTW/qUOEUtVURs36n5ZUdm2OwH9JywYIqUAhByi
C/x4V7QrcF2UO5yyOa+nQwRl8bW9ThaCucbovnbtO0DVOUFm2q/HRmC3G2mttaS9
vGnMUKBtAYz4kTECNwI4d5tgXy5yVSkLbij4iXZOKYNKck4pj9s0reSCwRIO7MzV
FRnCPH3gu5c3kelStaaAwT8HLlU+lIW5wMrfnJ0666FeMrmWFLPmGxvVgp52pIfx
kTBdhXWHPUjtK3BWlmqpNqU1lKFv/opQ7RzAIEllC5XStrJdLqN3bLGgHVsKx5Pr
oaPL4EMGfnqOVnAsqc1s4GUF9avGAqwYP1Xew6oq6HrhFK7+yMgm13sQNgT7CIBP
cn/FyMsPln0OpN/PDNlNPbmFJNh0QnvBZHG3ziTXJ8i2njOpbcBMxhO9cdG3OJYH
1xDDWVpFEc9knq7UiVx0npMMhDpvJ/CLv1HLrx0KPX/i2G1VfKz6Vo/NZpsNmeSA
CnTQwU0QFoftqvAzdpPAzSRFFXIxSlSrkmlz/rKP3QEAguJPw97DYBeqDs2SvnnD
2UVLxdRXSSofVRWsasNn4PmeOvyTzaV+3GnUdMbn4CyiQLvOhM/j6n+Evk8FMnwO
UQ+l7LFLfu2TGPVJP4hrPvckMbMsl/xsE0g6nKfzC4q2kqqQi2vp7nWyS7T1bSx2
HXomHFvDig3QXVgFDCovLH0fsBnlsasUISxwFEjxEOGG03Wke/VzN+O1FjzEB5WC
0btM5cWcxvwerFzgsQdMMXqkZJ1ib8E0HwtDf3KDyVJZBuxNbR4KvCu/lXLX+LGg
4K1THOAMszSqeCozwJT9zhwF63EtVnwUo3rjCqUHKRyGHH6nFxIHudzl84dkNHn+
IFkGwFLfyYEP1Y5RXbquZggxPgLb8UAEvE4m+fHxl58Knep6hN6zptd+Mbbj92Fn
tUE/inTmPQODSTa6RE/8tLGAh/8kgmc5GvT3GM5GnKU9hFu8R4EFg7bPb+tJ1eag
FCILj+DjmcGeI2pOO5CP7RwHTqwct/25hq/e6EzTV90eekq7lP/OF7EqgrvRi8jL
6/zuT811Lu4pgarb+nQ/Xz/4G+/ndLOifEhX8BkipwuJmpaE3Ws5soBwcTC97Oga
Lpijcoy70UuyWG5Unh3K/fDS6Dt9uoNSpzl4y7uuzMmjaxipFLo6XDUIX8W/U1UR
wEHC88/EaX//+uojhwKhetB3wF7ehy5wbY5MsRAVj7ED2mEcjXkN5YF1dJEmhP2J
ITt0DMvN69vme4m09g51DNRF0vx1lmkJXPCsj2Wr4cQobJiLns7wchAJtaYiqqvP
o61if7jlOBux/O3SP68SIC6JO2OArahJtUs52u+Fo4ezStYW8joOgiZ4ye5S7PvM
YfyRshY5AbmUXMA0+U/dowabxeAd82f665lzcH4JtaO63XR+f0D08CTt6yUVMtSD
SE75pI/UWdiDeaUqYUYqT9/vz0hH77tr3gKtQaZJHVQ9JPfFIqbW2RtIPHdxGNMn
cgtX1NRUJryOUax/s8Ypp4Z+22BHbZVpAWtPo6uejBl5IjnqtAeQ3dhAyEg4Hy3E
BqcLqcZs0rdYqSX63AsxMEi2l+LRnzwHOKZmdWysR5sgMX18svtJWXdmrlyygzkP
Pk0VWkMgVrCDIPXk0tWA33sXYvnwhlGkZUg1yEdCNC92/6W8jn6DGywqpfyZgp4c
S3dD4w9IkqNG+locmhlLOPl0C8JnztXfhMWlMqs/BI31dOwpQTTafUuZwX7cIt9z
O29AhL2Er32g3dyI59QnO1sQUUfnhwg3qMGmywn25cp3Yww/FpWAScPkU23by8ww
7hZ03wo+fGXwFWdEeo04H5ye33skZO/Ldvtki6iKlhl5MjTzSuhAWe8ikYoAgqea
0VlZXk2JyPzhjqq2QHsBxWcLklNJ+Ez1AU0oRwfpsJy3W6Lbme5qod1QOLI5d9Fc
j+/bUsq/jMFWTrKkjSfyB/BG++mop+YAyIwULv3GtqZiY7skWWWFbCV2qikf5Fzz
/g9tfEW/mQh09QKrcm3GfUO30zMTOmzyxGeOhZzTyeSzvM+/ca/KMy7cQY7TMAwI
x5qu0ZPw1a/K/N5KBYmI65scJgcDAUKrJL3GC73s1varf5z2hgqVsdTSRCf9cyXT
wbt4AZMiaHkn/1UM5MA28y0B3ZNzyo+xGe4wR0xXx4jBIGFaJMKfjwkNLLYb2lfq
+wcRBwSPRH6RKE+9ez7AMcHkebgHruSUZGLsjSfjrDbWI7tcBGli+qbyHNgAv1QJ
5gC35vXMWEYKIsoZN8ekT3prwqysCKnEq+J9yJgpW+G7n5NtfZQZn9mng8KXdUgI
2KuUzubYwg9xPlvcc6AbPXIo3ovlC+NvE1VmlnJvtjN/d1ZQGCHpH4cI4w6lBZEv
bHB/c79n0ScXNhEMbbl6Q5MR/5/G4gwcPN1l0i9YkUuE7L+U9kc7ClxIDks4s+sb
Z30FzNS3f6lyO65CmS5NId4JE8kP4KPLl0ia8Kj/ygiIxMu3PlXivaStFqb0G+N2
DCrQZRgU5ZifIMtDpfUMVlLPUJCP8zPhnfRWz9mFyEmh9fx56+yoB1SB4o844rvK
S2hx/V1AglZ6+KSRQIXmjse878ij37SaLe4uv04as1ptcAlwB/fKAjyJDQO8fbt+
ZtDrn5tOub0OQImVchjIJn//I6t30bKU2WylwirEI8SlyMtsQ7DXVAyauLjASiYd
q01k8Hcna/Ih4LQB/RNTS+gBdBqnf6SEigRprvrTRbIyOOpcI3XXC+r5qDJr77Bk
/NSYLKC/PotlK9jtEfdtchFCvNA14cZpwF+MfB+0wfJ52xsKiZikFOuvcgSVh8gD
h74fGqFVFZ/NyDEZLT6sBl3diDrBwLMSmQMWoLYyyu2rYCfJxpEh5vboXVT8MCXb
n6tArkXnb0tU5HMVb9Ndz9gAg7Kk/iFv/PY4oUg/ukk/I983AL31LPRscjwDLuFK
d4cz0g3+S4cllnPNamd3Cwc+NMQqqVuLzJsK76kXw3iCH9BmOkNk2ier1pR9MzGo
g5TANJu41Fm0gt9MUWg03meVKan8W5Y9mZKV9xWQrmXou7d9VHXTtCq60V5eM0DY
REpqQqj4T9205c0Drye897BQQ91PKQ38kc0OJXSQZN5uFhRXcx5KvMae2Qg6xQaz
i4ESubefVgbtY5wPmizjgVYLdxiGhCVx/nUaO5BOpvQ3e7gUD1sMq6/kvUh2Q7QW
qBB0bfYCbJqGu/32eG/3a/PpL4DkvP6g9YUd4+eGfZDw987Hd1WbAikhc3zHqzIC
bzoLnuooriSDOxfJkgLTjqZBZxQt41pthX8IF1XGHsyz5g46bEk4d2spQCAGhXAA
29uHVRZkBsTnW/env4TRxJjTlUdun7lZ4/HJFL9HsGcQOyxVO6K8hBydjvtRAhSd
OWgbqVmNMYl1ds4cC9l9ZfwfNDX4HOtdG0EAmqiviCDMkLCmp6d8KK6ZpVvrz0xe
8kfHs8qEROEIEl9ZGoAUqVBoB9pC//ct9qnM/PFVxXRwaN/SsUEP9zP2G37GEX5g
wYwKQ5obKAYn/SHS+rusF8MIpYQmscAI+mEAP76KkjKkUvfDO5yLt/x5CKavcT3F
ZgaW7PWwRRNJDNOaFxLK+mCH5oKoV8aWnM78KDmYE6fUnjlC+SMlYBpGFHJUfjd9
2B9oa6L5R0TlWEydO3QkBumaFuQPx9Y+BSe1ZdZaHx1FzJeAS5la84Gl9RPX8ZMV
D4rfJT0fa+/iO8hZqoD5JIpe6fgn289Sy+oae50wxVRNz9rlmmNFFoU4LJdGjj/o
cUenPrB27m8sfU9N7bIC0J84oMb81HcOaBUzwz7o+DqE9ziGRuZ9/B/XDj6UP0C7
BXxIGAFlgrB9WY9ZPjHJfGin99BIuiqwDPFpdJqp2CQIuL1d7XeTiEV5WBqAAvku
xPeUsOPLugqu9YDEJTQKxtEv8CwxLmOChNYBq5cCdioQ8J8EqntmqlpntcC0m7Ec
f62+tnJ+Hvr9TzeBUKVVwBzlH24osDulI0LUWpWcgdNNKEkzlUuS6a02P6gW5C6E
JROQKYSoBwv1CbPghyJeQ2Wu5mqmkYRB0mW9TjCrZsPTWTtjtQka7qyc0uopM9RG
AGcnu6HM8o9JGK7PuKfzNIOqag5Aj/P7F/65PLYYDhRRfFEZIqYu92UA8Q2AxJqo
g2nAhlumHvDtj+yBj/n6szIC0kkqcMs5oizV0kvW+dYfESL3L8eZoQQFdgK4nA8L
zhQWJLQsbne6GOcUis1Ef6g1Fq20NbRCvccFrdwn0JOfp5BT0bY9UeRAqCnu7kBo
p898BEq4J6wIUq5xW7BhJSxCcokJhWEumWWF8sjq3oeCpfjHLFfyG6Bx615XXTUr
QWv991x5VJzWQgjL0hgw1HBTskrG5qWwc8wh8cs23tsdjXNzIuQIKUqScxYLFJOo
jSTZJDYv8Wv1NSNG/RF7HyetJqzp3+qQZ/MLgR1IBsnOcrw2MntxwP9bf0xRWwY2
Oc+RTutzTkQF1Y4Kx7Mrq4kg/nhheRm8KjwXy0CM0KeogEOFGhCJsNnRlAefY/nu
hhM6pt6jXZFaKXT1p2rh1eCiSc04KVXSkHEt8hElXHgZhk7kejMWUezAI2iOGlN8
HPlvHUd0rNyb9kYTD+siuTHE847p15HwUkkB8e53jBgsoK0IXDF2Qfsv2JT03Q8f
FVt6qp4ufOrKRbnsnR7uuygb5JOEtG7q6p6EtvyTWaRMdVvxfwLOmy3Sp6Wqu1DC
KHYsj57Sscc1pZ65/uuLgX9VwDavAp7c91K9Nmju+CIKp6TFu/r+Ua1Ee+wpX1GN
YY6nAAAUcX9U9vzFnx01HCSjKFSzJGjX/0Hr+6UZkVENEn66Lv5o2811Lzd2c413
w6XnZXNTZ5//peOOnCmOlM7RM4wjf+lEf41qEQoxeX1Plfxeujn6R0kz71t0UaBY
xbcYE3RwuVrwz1ozuGkR+iVScT/gWyU6zqA3N7shl5m6g3wHm6ltjXtjIfc50w8m
Wpx9V5m6eJVr7/sK3VeDC2k0ec1eLLdfMr3wmvKeOsb/rQq14OBWAYnClFR2b0UE
AegkcVxtn1zNW09Q2dyUlP/SNY29iWVa1piaDlVOl4oVGqOlA6WVir9Il5tRdD1w
XaVdPSm8CRBSFEB4OTEhu5w+MSZUaRnkJ+3XEHns53nEVXPRlADkjrf9YTTWuGlC
SNC5YzqAyVGLJlNgLXiPexEA6Lu+YjNo0hcNm557fNiDnLkzBJYMw8cJkusH1BTk
TjEL1paymn0fLkOsSkTMONXw94kXy1qsAIQ+/qYZZWs=
`protect END_PROTECTED
