`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0B7UNQuy5Et9pBkS4b0eMr2nKa3yoT5Apsx6vTTr2jmNsnXB0XqLS3fs+2RHhB45
qkA8lEX7VfYzP1ymjWjya1Z0Kf9TieWJ1ll8bHs/6GZqleoLYLUmfNXD/eS9Lr/m
aHlMgylh3wcxN84GxN5OXN1FJnggtU/UJGK1BpTovT5bWNdNO8+oSuccDx6OmK1L
RPv+VY/ROL2SY8F+0mdForO1ezQlOtpI1JKZCSP76fLEbO42e5CISOwmov11EJjJ
cdIikriyORLu8N5pKOHTrQHVUqGPgxfS05ivq+GNxp0V6L+MBT1m3PjXe/Z9WZPz
eCnrr8T2Pn114DayjqLVcWZTTaTNTFf+/znDjzIo0z4LgXEf0YYdXPzCHr8/3Qpe
ymNKhl28Az9rN4wpx2E5On+ZEwPQmHt4C50wKhnvijFmU+pNO3w2lT9LC2kef3dT
/mPy3JswIr10p3JTyWviTpCD2P2QBISObmvtCYQH0vGJcPgSdOEWIh2jZDSqZlmP
FsORWYgkG/dMPNQw9ahFtMb4IYxSPWONoi7DZ8yrNSXzqLj57yJA2BzGj2S2heUe
yq5fJHA6x3uKroirI4CgZw==
`protect END_PROTECTED
