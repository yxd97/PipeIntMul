`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6auca8iD8CywViy2Ny95MDDm1M/YFKu06OmOf+syJHX47KY4pgUrbu2rn529UHA
ao1XkohVbuZSWPAMJVtmXaoOVDMmqBtDXKLH94VnjoCnuNnXFezDnG9+GwDGZdm/
vRm6QRhhWBEd85U2yPhGkjWbxy1ODeWeCOIvE/VdFH1/hJ7e/4wRpsCeL4fBKoYu
JOzK0Lpf5JiSSJe5GYA2YsPiGGePClLiC1netUObOUWRqPmdMlFxDJpitMEBu0oh
fo9yGGPmMzy1zmLyfGcIIGzTAbgbRi5Wh9Bz290/4rY98Mf+wBnCXWKBDlZxtpve
7NUVkL0wFp186TEwH47v7uZpaXpGE0bCC2YH7BxA72zMcO23XsQ9cxgaM6F0pE/+
e9yxhURqmXE1WB9mZsORk6Vue16KTcxy6GA/EEWYjPJ8slfYiAWnRWGFb9ysNMbZ
ERt2d210aDKdCa3kouVcdCb5aCWLohFQEVzHCH5XFw5tfx1TL61CH30pjkBfBzRE
7vpQN4quCjrzRr7OQ7ht9+57zLHkciFySTJDD9Jx+TJoxAgFl18q21uFO6c/9Swt
nXMPP5XPIWvOzPnJ+NQtFXiP/AeT1jufAf6kEXPA7fzuTiWuSqfvf/w8+i8EfUF0
JTS6SCmhQhn6u1pfGizofV4q8Azpweclhd2CF/imDOb/ns43pzxBUAreGlJCFFmo
AkPymrfyukYtv5t5EaEHLaw1/sYvyB5nQKidQglaPWquWfugT3/qMRBaX/1IJO2F
FdScps5Y7o1F9jXsNZLvIg84MCWCWw7/aZA71LWU5A13R6YCRm5Ngb2KCuxe5dWb
vmyaB1XXY4sn90ErHYE80JzyXmDbkJY3e3PyO4wCJAaS+4IvD2uIKJWqcFMPh3Fp
xtIaZgUizN0wXvJWQsYJfwmd6jLJgEU81/pzJ0aXW8A=
`protect END_PROTECTED
