`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CBii38vmuP1xu+mSQtd13qtPLo6z3lfvc2t6/U67jv8NyJsKi1dI4q1wCAs4oKA
jX81Vi1/977leZXM4EDeTMJMEibu8Pdfle6zSfvlL02L3zOWRejNbvBhOFk7PkAt
Gnb3xeNTxX0e6b94pflvWv4tIsoHOvwPc66u4ieZdvsm42JKFVUbY3YSGEdhoRGf
DmVgu/vQhy0qdUSM39BnE2vdAdFoyOaKFs5NH3lbWci1XnNVl1sJqlhJjJVdkzgy
V4LvqiSCIz4yuJOsXJfchSjVE+2V+SnMLPyK1Sa7qfwTZihyYbsh54OXEcHC7CFl
O0R8tV1xBYftjJdc6azfGIqRuCArlB5hbCpzR8yAQ8rt15Eh7kSjVTP4pCE6k8Sn
a6fOVAUoDk8G2ZPBebOjf0CEeDIhTpzHGeJg92/k20VqDE5AJBLSR7V+jeEfw7Ve
B+BcsQ/EyhNNgUXkf9cbzTAWl4cFyD4BFdKbdfryyRy9D8Ywzb1ypsJ4vKw6r9J6
R8dqxyO4XbjdhzlcV1BviNl+iFTUpIqzhiWcy397pKwOnQGezKbwi2+sjw9OnpYS
P7efICpjjO/hlXiCHLInqXWgb6ddbvsedW78TZq9aOpcOrsZhPTZXWLDg5GxoNJG
VPcYEKLP1xKjq86d6ND0DyVzro+DhNoxnEymfK3Py/PzflBXNvVL9CAn4TsXZhKr
DbHAUxrJUsPMTrqiXIgYFNSZu76un9l1WLrju/zIacqgXCjCMTSH7L0nHl8NUJ70
9+IDoVXi3ysjt8pgOJqtNzQPWZ+J/wWf5a8pj8slxRGpOKmPALOHMaTSwg+egx09
lra8H1UshQJP/RDtHc4d+7k1rzVWHS1H5+PYwGG65XSr66n9562871nBgKFq5+8s
CFWHyC5vIwgmNTU/ViADDyqYUXgRLqlRhjuFRxC1kdPUgptuntVC3tv/DxbPO8IE
hsq7UbfQSkX6j5qGXDk2jTFajEEKONo39YdJb17XRQFk9JQ1rLkyjcF8p9EuTaOu
sazk1gmwqcRUAU6qHbGEhAtw8R8nFyAoBTQnfYVKOXWqQfwzyX6f6MU4G6YOCLaR
6k0vfhu5hiKQoQwM0YsZaIb+aDHMcP0q4rOXRsvdlkbJ72W+J8DtPFsA1FrEjqrm
vXnJXck9Mlh+kDyUxLtvyUAiW+aCP2ULClMiqOK1+n+dUjoPQZJmHaDJq20hdhDV
bsKG8JE2BEPqPPML9//sTeceWSR2/+YYX2+YiK7NGet3ouYXosW3m5x28vYAKCIa
y3tUv0tC/MNeLPlChV3OshqMLLoOEr5i3OS3unlXQkx6JBrxn5BK28pbK1PUrSuM
0r5O7TxlYABKeVqkItjAnv7+qBE4AqBhnWjECEThWFJ/jdf0faeAoYqZkiCsIrop
LEOorVmHSq+ikqrpG8XqJZGeuczI5cLpiyyAOYsu0+kGS5eW2NKLSxwI1nCnF2Xm
KW54Fdo86ZddwzxTdRgXq5IDnB5w3lihiFxQ1YS3J/h4ywfsAUDob9BoJlKh8bsY
`protect END_PROTECTED
