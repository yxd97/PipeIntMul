`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NBzUJtDMEWZMKlYBSo2KFADM3ebAWNTtg20wC7XYIWZX12hjlLlcu+wml7Jyz38k
+JTshBmYt5EEtgQlVDRKf37taLEL7Ahg56W5vVuf6Prrxba0EAovUdZqQPbsO50F
r/gMoHQdzR0oXqkMfByqsVdrvFscOCSCalZzMMLnrSLzDXfIlpqEPcEpZqtGwkyT
qoWxXnGdMvmcum56xxVuOkpRu/NBtn7IsKydSas1p6qcaq/Ug5lLZb0WJCRnYOom
vzP9xKaUrUD//ERH+xKiw8DekY2xT07x8kFmlI+oIejE2tMHaBXkS+kr+fgIGPS2
+a7Gsa5X0+F/x4iJOdQEDV2XAw6y2dkV/n58KkRxE7/zRshboBdDg7/g4YOlTkiu
w1MYb9VorHIhBaFdcTsA+aB0Z8XmuZIHawWsGj+D/Ko=
`protect END_PROTECTED
