`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JQHjDQmf46SZNVPuHor/0CAq0Aa6N112CZkf9RxhXu01UDhRU6E3mQd5N6+9d7yF
9VicbiiHeqLs+GuvP0Ycrjx4dDdmx2SbQ22RoRMOPmVjE5IfcoE3lM6+wHiZ/EXO
UC7WB1tiil+Kre6MCkwygL4rupxLhUMjiYkQOZ1lARJJxLWmvTDaOJ0twr/X2ilT
hJPfvg4S0nhuGTGApxP2oljA8FRU8nAOtWn8K8XRTUCWhlDdlo9PKDEMpB5EBmJ4
`protect END_PROTECTED
