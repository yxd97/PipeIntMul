`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zete2COuzvLsXSRz5LCMRXsVPkWIB7Z35SU/DNL/H6IEbYy+G2i7Bzfg7I+4RSFl
KmnauWTnnmw7W5/tNFb40D9+9r5eLOl9iI5YzqAeqC3Mwsth1lvKTm3EUeBqSTCA
7XuQqHObuxd70cipOLpGgH9md4hUbG9swaH4hmHniIGub2IsiQvWSA6SOwjiio0R
AKQEZnwR8JdWl6smZ0o5M7+yN4kJMMCQnObpdVEry41mkpnZySjv9cn/fc3zbJoa
jN1LBM3xZJmkd9WNPfYYWORWDiOO3/sYooOLRz/tqt9m8e7di9OPACBcwmyd5s3o
WwMyG5/0JQP8jevqh9UM8CPhXEV9wrtiAr3TdolCgDJCKuB7tpEqSv4NbZ89X/bu
1yuUZogkK1fdSiRi4IZC2lzeHb+Oov30J2ftRAxdyCA=
`protect END_PROTECTED
