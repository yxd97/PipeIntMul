`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iP9tD7JcZda5TxQzTcOHGOohgEI2kxd9xi06M34uR9Ct53Tdbc8oyvDQUfyPg3yB
JNiA78NW6TeIfrFUECg0vBy8pk9MXFwNDa2iNw3YdwTdwEVguQ2lOTUop4yz3pzt
xApQdbzzEK7NwY0K76Vosvy+xw7bhgNPGUm6HgbjWC5PIq3pJJ55ztJinbO7MIc4
055WhNqTFBqV2Dfc99U3XwWdDONwjMbVtmSHYhYCCIarzNBIyIO8osfvQdjFRYSn
QkCIma2Kggg7IJWnkNADi/UHVUmsvSD8TzwRRreyNy52ybjpKHIRgdqPdgxGdd8a
Ue3+IdCPy7ua/UaEmW0ae1CrruXBOdNxDv1bDcxFCqYaO/LIHwIZ0EU+obZD5sas
UEBcjiGxpb6h9tkF94Bco2sJ64pdDeq8xIj6KeZ5UZj688BPRBTXJlcDOPng/YDB
`protect END_PROTECTED
