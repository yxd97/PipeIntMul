`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yx9IAjxJ4jLzdIcEsVO6XoFGaozOkkE5AqfxVfevlRjy48wAizgCTg6Hg2EOX+l1
D3RHY1J49o8MaSfGaODa3EbAn7b5jLJ49hJIVmINu2TUQoh71etK+GG70XVi1oSW
2iGXWrX7HPdPNmUkwIZqGx9r855p//tO0VVzebBldzlo+HGSpJZddc0gxE+k2vlq
LD0BUpYrjtZSG/pH+qLOETt/qM1JM/oRQjaEX9UU7O0a6U8OLlyN+8lwW+4EC3Yh
Gt5SUjPYJ9U5k74+irt5NzRfeKCxgtyKr86Oqs/tR5QsqzgUaeBS1o14HCM+HU7y
hzrGHz72YJPL87mdy3gM62jaQwALuxxvBFRWpFpxcKyTSkBLtAdEoq7psUZNRzEl
1fSgkF1eOGXPBVfae53iJlnFmX5yl3CkPJ4fv/YfnO0=
`protect END_PROTECTED
