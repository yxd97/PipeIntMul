`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/wZhV305wNkETBpbsGbKm624i9PmcBmm+NwOyNeYuuhvoGjUBYnVnerCtyN/FEnl
3sAZGJq/1qAY6LHCDnpPP9PKf+Xw5IODNVqzqiR75eHOgMdos66yOSuhsbZR98W1
Rzkbk1JJe2HzxGWhiOsQAMS5ADqY31jzgNMG5pQTRNKAEjKyBdWFmhBO4VdDiZii
ZJwmqsewVbxugLPy8UxVgQ94XKCsbzC9NWYj+oAhB3UoH8FZUl93ELWX7shE7UWX
W1RU1rBZNLqFrNm4Fyqor3Jtw+dcJUZnY8CfKKknLUvGlHXLACppF2NptWqcpi8U
ZxtWSuLBBKX+BFEX421pdeCiQmRbDFdu/FG18OlhNAWX7rUiTCqMv3UnKpOlNVim
ZSvSr4FTExiOOqvLe3dxre4nm73doFCpIj9aW8A+CHck8lzAp2PzReYB9Z4a2+aS
aOigKNjTiyECPlb2AtqOS4Wp1jRfZXWZDq0RfrkLSf0kiLVHzz/GMrbI7XiMpbCw
e9LmjiT6/xsmziGtQ/ukgA==
`protect END_PROTECTED
