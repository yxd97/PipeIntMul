`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPg8IPmbKSXLUXSYyVVD17giInOvOiKNl2MuiYmXlCBrOwlhfzm3bFejuJWOWtp0
v0kk7TQZ5L8a9LHpb3EOG9X1iUKbtQ4Wf6NvhHVnxwzxuD0EvX9JAFgO+PPm7tjY
T4LzwVnOLbGa06gb792QnOh1FaUYsiEa6gTxOauzGDaHZ6/5ZEDpPX50kzjevjYp
iilFJMWMjibzNtM15S+cQf5WzMXo30PGH/kWd6TIoYZudTvPgwVgcIW9Dr4+MlMZ
03Kl1U1a1sEmLm0vAshEEfLJpDETEeY309w7igje+rjHNp6YAeb96HkezSAw+Z8b
tFtGY96ZU0FKW0CYsbyg83WdkyIwgvhMQ81YcuzJef0VVIZ2Q6CRWBSNqeeBO6Xi
t+TGkMYFHy1C87w9vuI7zFLLYW/dgHM+neA2l02XBjyobYY76dVW6PkrUdhc5QKF
`protect END_PROTECTED
