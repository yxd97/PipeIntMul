`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ERqpbD5f47pil6EEncR3R6w6hnTm3CGJ+2yR37Oc2Si2U4Nrl5lLg4Ab05vaGN1v
RpsXX0+FqNa26v+EhukW6/8i2ezC4CbwqZU65Kzx8QWoHuBckLIktcffuyop6RGA
keOUkuEfVRPu4Z3m3W40wr0QnW2HpJbT07+r/XVjKUL/acmP109sLnfMvpaiAu7e
15YMd8UvX5ifXUS9uvWk0tCmnGPxH3pIKcs/1HlRj6v71FgZZmEoWTrHp6RwSA1R
m+MtvXc3Rbb2Nbb/Ndev674QtUy/b9H3xRUsrCH32MhHQQ42lfJOzRF+b4KvKayR
GGAzqtIFiO9qEYWqX1AvKQxTIamCEJa2BVivP9VmXzmt1u8T7l4YYA+fgy+2cd5y
DM4+4l5jazVeEDoNcgatQajkJR9jjeveshrnJIhoqAOSFnbZCyX7cqut7WCURGzc
O6PoZ49tefRPAiWBNLLfL+Mf25lj+UFmqt6HbvOOGnVUfyK2oHiVNQt8EMiE+lE7
SomdEby+ZA1IZ/tO3ssSfYwWLj/JWxWi9xQ/D/H5AF6U+WAp7L/rkK6Q5sRgc0bv
kR8xCmPxX803FIMfe9+zLIU3dTMKyNSaZq4wvTi1XTuPyBAXcpkj58G3Auoj+0hP
eYwlD2+aeegWYjf6wdCVvXZ72owFyGVS1VgEUBZ6G5OFOSW1DQIvCGQau47NrZmB
260luYUOdtmxOP4vb2qZudxbI9fw8QCNbWL1klL4w+IzUjDA6U37cteRiGO3eZMZ
G21wKpjWnEqaIsYbqmHY+hrvSZcJLymQBcUi8CqtRrDruXLHcZwrt5Oczc3w4sDw
67bIhxKXfysVLyyIJeUYY/i4groOa3Vfpe4IWR6vKQcjGroirRfB46roO1+3HBdv
7d4RphX3RvcIKxc8JYMi9lfsWHF69XBI0jv0DjFvN13h+3Ith5f15+pOQZaQIrIZ
4v8nZDOSvmtjXya2WJQsLIqsxi0xPLbDSxE2R3NEwVgdxtmCloRJfwfwDAk2OKab
kJ//82fwrSa0W22APbsrbZqSY0NA4WvQO8e4+/Ig7DENkzI3O5xO/epKQFD38K9w
sbgUrXpqIMU43aST8vxt5A==
`protect END_PROTECTED
