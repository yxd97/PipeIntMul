`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CIv/D8MRD7eMAAKXhi6Szq+X9dQKI0ec5WVjGfgyauxJeQ8y/pfZ5O7IYI48JbEp
tjvGrSGs3kVsmaCZx94fkjHpVURrx7qaFgsSmO0jdmXNYoYpM92PMQI3qwilyuOl
CZnURhktIxfdIbNeDwynyC//MpBN9bt2iWizh6Baxco3LbJuc07RGLjseO2I0TD3
8Et/B+X+l/5PwHnhSD+A6OYPBBcstqEqA8KoJcl7xTv4/Ak6bFbfZT+5AFwuBLxb
NzdkyKQx2JTwyh99S/MYlhDXMG8/WoAfN3D0TKqPzRZqq9rhFmrBvelCzBTijTkc
8LhnzMml0nIWK7Led8Nw5NPRkWQwu+RqnDT4ylnzK6/NhXNJrmIDE5TwVTCR59Ux
sUnIdJlH3F8pU0KjARWbFjpQmJEc8ltw8vhhYps/yQMoKngzXzIyUIyGu9sbQcYT
TIMxUeB9GciP1ZC05RiqyZ3KHta/8EZKuQ5xprTdwMXIm3f8nPufrtHPX9VXeZ/Y
YLWq/9jezW2zlTCVcUpGpIxtwG+E0wjLWbHKbwHQAcSy+AfIpmU4+unqe/xgEBGQ
X2pXufuA3XOBtHYlTnL4Zf2KqDhRczI5M/NdJRa022HOVbHCm5mcnOBRTKDKhIb6
JrR3eS9M2ZSMmckK+SXfNtId6oxb5C/L/St1g+LKll/ropQUEIW4tl+xVyQcLkML
J3k96SWEojZPz7W4UDsW0XiIzLkJJzvM56JOzh5RVt45robDelGSIOXcpqUqTLXx
Ne2duGonsHZBiKTQPjPTIg==
`protect END_PROTECTED
