`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxJN/bwtfIaVA9bUdfTtnHRlC6VH6PS1+/rWiz1jAHrt4j9yr5Hcfid2y/CzOPK0
cip+SJejNzPi7uKBJ7uHL45DYHMejBVYt9woEqiRKdaVUKZ45KeTLVj05TxynnB4
8SRZMb1nfPc0S+EOm2mGdhGTzZvFvag4vZXiV9lidcwuCBcEYUlFV2BU7qGkFjfM
fQ9zzIZcX71LbjGmj1GE9Mu+CdWEeFeTZcFiYfuJ154r20Qz02aZdXzAknFMvyI1
ySailBZfdiLptINam9J5GOtflpmR0rkaGdPMy7i2LQ8jJ3IW1b1vxpdyyh4rXelW
eUSi4a9udBU+ibtRgEuTvWiv3OQKtcP3ghYtLUtPXmiuZxOkurEOPRHxDAaVqnAE
iJ6EM6dGNaC19FGeNQFi+jpfnkFEUEk60UwXQxJV3DcpfEtJVwfqBM1ozHQ1InSZ
8dpxUJzuHgfIbIZTMq2BhxqFSaMDe5ZcK221UCensM7lw+YZEi79nE0m/yV7bgRk
fZme3YsDsbrAhu1siiWiB2T7PMK24xfAzbPJWDdqYO5Xqe11ro/BtawlS77KIoUz
k4M9vPAq23oEiegToxBiRbtlo/+eWY0EpTjIA0EWVJSAnR0rMAeqcOWDBoakiTiX
ObXMiek8BbS550Mc8c29RhAWbowJgmPhnoTGHeMtM5GuFg1Ycp7hjEtAvV/pgDRe
b+UAfeGnixu11C/q0SmLRRrZIpSut/fQDhvP4vDa8LNWwZSS3/DKhhndYGVb4RkE
wiklAxfyVQCpJ2rP6RcWllM/qB84wxZt4gHuLLziqeDbrfamtaiHUcgkcn+GN5JG
4/N2OK/vr1h2NJVG1q5jZ5XK9j1RRfvT/PfcAzHz30LBxcN7e1Vez92pkD4EB8ui
xWpbce9JVUeHZvpeF3zh0AuGWgIDTic9q4QIEoVaSjcFYxPE7UgR5WawD6XXinLf
pkDcpR3IxSSIDPp8LurjaT8wheGMW1KWO/k3Amys1sL/IBZgDsKrBD3Qj8jjecnm
wgPPfUYNqr2ZbAlisFeRP/lyzh9yJMQJtiKMFrJmfgUKoPP/YuhKmp/ytUxGzFps
z8nYtMcOCdhDDkUIQZsZBbY9XKaJ0DxfvOWCTNi2NWw/MGMSMR3idk+Mljc+x4De
Pyq/LkMR6rP5/zNH/+IqY2+mEtFNTu1UoZEkDdIIC63qO2oLbxT6fGqrkGRL+0wH
g1ppnCJ6Yn8kay6wznIRC8ch2CdNh53lb478XIRAVH1i3AR5yJVcp5ofEaq5BwI/
EpCiVHY7PsJkik92W2QJaiP3DIrzlyiaPRTFzs3UuznNHw+2B2SbW745ZAS2ZlRD
yFsz6j2E0mEVHoJZWUA+nm+bNUTx2Eifo1CMzbu1l1qW2bopsux3z4G4CCPigxbJ
rgmqiA9AwsZ57dWyd7XqirjSiw/lLmIEqomLa8BzGL1CUBdqX0mhefQunbrM/1KC
gV2Ms7cdyCrI/zqz6r/F7PjyyexBAHao+5jKlk9M1TAk43/h2rmpBp8APPJn0Lsm
X6iQDMPJiFmrzQSSEl21OE3oxLMLXZvhBOngt18EV7ILpifIMao2+GfttjuOvw35
viPTj99E7Un6OMItJmi+6A9O49GP/rJEkSYr46XIAH9f8wtzug5gCtdsIKA5b/Xx
8WmE1WiJBQcptYdFO9eSODX+794DnvHvr1gT5ZpxxSvN/5b161sxJgZ+48rOUz+2
HLjgUHa9vgVHMpxEDgaTIs1vexXGXvCZkoHGwhnzzkt87M8QkjcNFxfi9vC9pxON
Rt2LBeVEaeX5+5MLdKp9KmTomSvifbtBZhL/Af3uqdeyd/dapda4yrJK5XU9ZiJz
SVXanG5ZE7iMm8Aqa7RVBl2v/LpKnchhDzHcbBJESIM7jJ0Z2HCcgbzXdnVADGfB
nDbI4zgS/wtGMkj2QWSNNGf4XEkik3qEyB6VzBzyUe2iXETqSlu3AUdf225QlAfI
STSLWNGsF3PNUU4UgnRy5e5xD0BPSP8WSc7pyEI/p4o935SZJZonuq505xG5+ART
6XkmLs+ReWN9F78V65V9AyZvUYQHCJyIGxvzerCfiQkXz5hDG7ST5dl3Krhy+F3S
nHVksQdP3W8N449GOVLrgTN5MAx1RbkdqOuTBh8fEcW6EPAGCtf3XhnVh2xIJnRB
/8K2cvG4DK+Fx0lELRcajBgEJA54mWyTdg7kaNqdcM2z/5fhAl4XHQ4v2zRH3FKs
Llp/ITst5NXoNx0V1Hd81JxyG+0guw9v8uhVQ92ZRmUVxnGONZ429ShZr90KDkO8
NqS2GaJUBhe0/JZxtne6Dg==
`protect END_PROTECTED
