`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bNu762suQap/OG9p+Q9o1yxj0b9obZx3HkROx09qvjJUQW1Re2czk2aDPZZ7+yaB
vqRY2JauRgdaTPsbkRqiwexJMjSkEga3NiwProRsG4lcEgllee4VRvGRNpmYdunN
jXspK8u2ftSdCi+zFiHKk8HWH2yBjn9CxyWuaX8R3uW0Q9pv1yR/L8SjoZ89ysyT
YCYgEb6sJZf+wkmxO/u6uJ9ysQFVHHh3sICt0wbh4qzdQWLr2gG5VpU333pDdo91
SKsMRCpASqiAxQ7LmwF8/semBF48RXpkVAdKhXP77IbJRXt7E299KVGszZtyjJyv
wfJHieQwF54c8f8zo91g/rhLHMrBLoYDzxP79cnbj1s3DTQAaTxMYW+seN0q95ml
cP4rRbVQLB6Laidx0FsiATgqeapACEInAzb7FN0TXxBW2O/vo0ABIA6uLCNJjfFK
gPF3KcGhGa7MLmDHHIZArdT1zhsczQdTc0htUspFPNjDvY7CNwHwe89Oc/xKB9AO
/x/yHMrKopPCrZiCfloZ6bsVoT9ajSc5BD2kSlLsTVPMm/XreQkacQYcAfhoyJv5
DpjmoluzcZcjEI56pubwA9WYUuNWi7PzwcMm86aYTvlwW+gGQ7IZZNDjfI48Uo7d
amCxV8li5oi5Mt2fHnyr+lIqcMhQkO3nJAMSoJLPDZei0gJYdSr70tDHSYiNQUGs
ZEB81cYkUtWuqgPINuEVdAJmtV3hp+INITtVwQnxl/swMULN7BRVx6c6R3yIj6IB
3d63yh4a4s8f5H9iogYZdPgSt93uIBbMUiqZSp+1IB10niGrJv3qlvefo0iwWDNI
gUnhbmZH8WZhg2PcLThAfyopM4W9GpcxymC9ko71dL1GWzhOsJNx6tAn9NddxkmC
zF1W07NxxNwwr1lLNypws1PEbfhSCl67wHwwRCnrTt6ByeTt1MYMegZm1iog0DQq
/oX+PypzABGWotNsQ3zTEldZmtk2IUwYDPV/2sA1MsSmBM4N06xlpdB0CSWB8RHk
36XHVqY8GTmzNzHLknQU+By/tHyy3cHWZ3il8Guu1/OZyNOgdluE8NAmnTBaEPkB
8LgkelvCcXsoESou9nvDPRlFLB3FeIfKdDw6squTiQdG+pA0WdmF36hwO2ZH6yMj
U3YGlx/LiE6JyMZl8xsO7A3l54c0TTSEz3N1E0EeSzdPKw69MfrKwKcK2UY+8Hc9
Ss47cND80t5V1v+vVZ3lH7enXxFxwNk7RinNs5uMqceKt+xrtkF/qn0dKBSn6MtD
4QVhY7XrCEN1Y97KeIb1YmSaIUkyq9HZxnqeSlkBKojBWUzd1KH4rNT3wEaApjuu
C+8NSbJMVcOF7BwlHGPqUjTxJFqNKPIH2WWNHoN5N9zz12FAWVabXotMes/5qO+M
i9AYZvVLTUEpd9aGktuO7O4DdtxIwSiIqNLuC2H+JhqaSt07pvhDp9qHWjJQCF45
jJGyqKXEBvOiimsoiSGtmxT07hAqdl6Vh9LKoKQeJ6aJlNViuiYossy4AIqqtD3i
APYfBL8U9D/6b/SNmx/DZH+6aUEi1TjWpJFC/zuLqLDysrgKpzgHPEau3X1hqJ9k
ZCCaNf6I6lcRmSeCYhY+l7791vQCmQ+/wqs4iWPoLrey2MG06Gjcb8f76EhJ6C6O
EikZ2QakJvj/+9uF5OH0/kJInwUUJqm4Uz0D5olndSFSdxYPzkuz/+5OjNq7gzCa
HAmNw/1Hx+B9qbjqfJo6GvKar3O4spKwieS3yAWYH/YYIien8z5A32PAZKO/IrDj
j7ZyGRImzrM+kpvGiQa07lxtxHssFSnJWj9yLjBpWIvaZUa7XZ+dTJTMyM4XEkcH
6ImCmb6Y3vVrZHzwDOfP5HqX6ix+7DIRCPHrQ06hE4a8d/LhX6CbmRJ7G1AnPu4j
`protect END_PROTECTED
