`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKCgyyQI4Tj/hobK8iHCcgsQfoW5Vze/gawxGgttWSyRRVBqOZVnuHPy0/Ogs5VA
uaTnpWypBBRuUtnIJFuAmAPspZcsccwwaKX+1TIBuBSAnM5Pv5AMDVqWEaFkE5Zi
KLSAGl8i0hMgKy/+/2hlJKK7HfUgwhw6+hlUcl2FjUiYbzVqNcTuQpgAZO+oq5Nk
iLJhdi/Ssf6tqmEvAlL5ImV/ZLrb1BsIWZ4Q1Nq3IRo2Qyq/RGCG/LCA7kkIg4Tf
mFTImCTwCYYNmlAYdioz+MhNtTUkzCWJXL8LEAQEiZo7E4lrBj5Va6atWG/ZQm1a
ShZ/tkYcmiI91q0rtbbg5+N9H2uYXrQY1UVKo2AGflubeAgSjAB2mR4PkxfaFi+q
e697+MFQmNRcUOxM0D4s/rt3Yjrb/uMi6Au4wu+ZZFKLaDQHXI8XrA9he6SnJmiS
pGn6oPvSSkiyNkEL7+sBdqE1tr+6UQ+sWYPjJ7ivoAkJRF/iJW4JIYOtoV0L/Pgu
`protect END_PROTECTED
