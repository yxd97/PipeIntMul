`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9pqBhhRc59SDZqHXI1TEd3tKwz9J3/4YcauM+Ww5Cw5wZEMJMQp852qVsYnmjmL
SO2fZ9KVWO7evEDSul7omUc7HFGwTMW6j2Jcajrke8uyZjyqUize9rzjgRATyKxl
eGSGqHVXw5du4R/IV/VQEI1MDw+tfX8OeZssbWBygGvkTzMhd16y15peDcEQvc8k
56a+n1ttC+CS/LjM2zGhvhklu9s3y+Kl9/qMMIm2fjgzMLZu/sxdf1LHLhJpBS66
1XDZnnBO13X+GsfMWsbngEoZ6x2y6B3/U41twSbQBEpTGx8ui2l70S0NOY0FxOqw
J98JzJWIyOvvoAoX5WNl90Fm36GGxUuGnOA0rkM6ZjUK8qORWfgc9OcVjkgUBXH+
M7O7LTpo1GPbn3eNgC+/0CrXcNTD5M5NSiGsOPUAdfcYroKI0nkT684q0U8dPf5I
9X4MG8JYp0TKpxH3MId/pP3BQpdufpIcoA8nofuxqnwA7pVOXONNnBGKX/dTODup
9vJ6Hj7KtFqz8afsUzi6xssnur+4TeBqWsdNqTwFVj7Hb39wgatD5Fpz7JD3DhcH
9D9qMK6bErdCyyToKljQZxovmGZsY4Tw99ygsAxn5epLP8dgJoORNSbkL2oOLCO2
Xw03VZtV+BPjSOTGO2CADPHBLKL8jrLa3BOaz+evkKPcAs0GwA0GdYZ2HFuWt6wB
Dl73pv/JjwVXDdLr2G8wyxAPPCSF2JK9VLDclaEaDgP9AjOe69tKdPknXp3ejli5
Zd4kqZ6tZvSAKpLgu9NvGQ==
`protect END_PROTECTED
