`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSC4boSBmuVudjOjbQ6d3HbuHY9jhextlaxAOUgMs2B3VkEyhVzNJg8QJW/2m78q
n6QpWa3NLTWsqdGC/3XdVME0Yb38mC4Nnvn/G9FO5et1VSO5x+wsLdJm1LiVCzjF
bR+kpr27ohPFADpOyG2XXMS7j+Y1Pbk7i5PhV2gEs3BtYpYVn+i9fRUXrGzfVu2/
GpWkY4Jph9sdhz01Kd5PjbQg1zaPnAGvJVBBDpD8+fyIeoN0NtRDher6nc1VFfac
XXajqq1IlXBJIMaIuaJL/jbR5vDRYBokj6uKyfR/JyBM2J6PURRJ1zThvgTJ0lHD
4p/zF9V4hJsLRMO8ZXQkz0PlntPYRYExKjhUw+Ca8I9/ooHTPFskTh1Zub1FuSTi
`protect END_PROTECTED
