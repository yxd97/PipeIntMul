`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vwb92BhR10fr+3xm3TsUNfk8B+lR8w25YGtZO9zmDmS9T+gfjPT9xv5NlJ1rETUY
WVsdWYmqyRrTkump6HVLsglO1AiMt2XZm1qDv5nhSrDp8LiuJMdOBYTz27Wc3MKN
/Hw8RplL+5766v0g0WgASFj8EUIhvDstQQF7qk6feBWBXYXP5999tYFK3OOJZ/Pv
QJ+M09ldspTNP3B72/nkZ7cA2HVlwxY3JsE1rFcJ4OiqUnVQIfRvtXOZ82PBYmpT
oZGmOs2T0tGa73jOTO3vPQ==
`protect END_PROTECTED
