`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3gM3ODHEYxYcq0vN3J9B5sX6Fctwc52gFArV60OjB+QXvl5EkCDo4KXRuriqJoY7
qyuenzsbymwWcU/sfIaLCDTXLXA59sOpDNQA5lF9a3fUSMLI7yQO5V7U+lLXtyth
FTTkiCtY1DLa0yjxj3HQdHgTzuvFWuFYHqzmhr/FhSlkg9I0YgKzrSZMXwxivxBH
ByWVWRghatvnO1u13LUAMzDTvz+sBliH8ehXZ3yu1+wmf9ptB2fjSH9GlXjTWwUv
0rmoVpm88pOCyP82msiWN4HDebWJwycD534rE9lYcKKHMlkh6pX+9AvjLHEeOeIg
J32awCchSAM11kHGvl2cAjxSJJLNwunfpW/MTD+SgAQ/AEh7idTcvoI37PkDLJ/Y
V3LMbPYCtjqE2QDgLYnIt4I0dvYLYT5zGy3NiCdR/y+D+8hcWS35vF5vhGjda8YG
6yWzvkT7EW/qdLan7Oy+bmCrfQyg0qI6YSBIoybbeH8Qgq9kqguZrAXu3Uy+ZaVm
+pZsrde9BGu/9T0jJQdeRD0gFfSQy9gF5Cwi1ouNZWUoYNjm0Btkm5uxtmbFEhPF
eDYaWUunR9rohpnKPN8FFQ==
`protect END_PROTECTED
