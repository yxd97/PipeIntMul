`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G2Qn4oWWFvCXyZPaHjFTfJJ8xX2d8VzqpeVOIpCql6GGxIyz4TmYmgDdPy9Cat7/
lnI7Ps1JM2XELoNUNrL/2/MAphd20cs6hMXuftLZ6v18m+dKFZiB3nWl/7I+T5MT
RX0N5Q4G03Z+8GrZtLGED4Xt1/H9QdQ/riCbT8G/Y0zB2HMkmtmkG4Kbvh/PyQDr
QuvftfAE+Dt7gpVAs7ZGDAAFC3nhYXGhD84f4v9KA7i+QJF++BSutcn9CJSCzG5g
GCb0f5Y0wQHtpYjpKyXuCIXXozwyuv28lzcCIabVoOnb8mE19bknXiOZddBSzBVH
YdgAmpL4DXOVUulcyVrB9FPehJNlMD8f0+p8o3eHCduoGodvS1WUGgtUfGQJee/5
7wCLzU/cyxKfHVPzzzi4PAQ7wXip63I/KNzVGO+fYd+T15h2HzY5o5y+HvE2raXx
moBq4YB8x/7l1mmCFt59TmpTKZpVSzrH6oqH5NLCH5ElW24kW7LAYDgZbrZ8B3fX
0Xzc7H5BK+JhWp/nUf9BtOSy4SXsa8mGb+baSoe/zmU=
`protect END_PROTECTED
