`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bUMg4G0d3OV5zeWjiZZ9qY0NDGVG5dsoVW8f6ajmdE0H0LExIqkuHOraYc1mHkjX
3GoFkg/SkOp9bSYxeR63XtMfMKSrqbEOpcn+b655LlTfilR2WEyXB8UIS6UTJbSq
/PScdA4cP5vhzNmbJ0P7R3suwxpZIKw76YwFh+6WtKXVJzY1AifzkSzyHio/kiuO
1r0lwhBRyvf+D3RcqbPM9Zpskt7OfaNCl0+3oUiKWNzsYusjiD9PIHRfAtXt+JoM
cRyavC0h9nrZMhzcUjb5V1hTJNQnrEZq16XziY6MnND0aI5yOIQj63lkw9DOMniq
iox1v/Fw8+RZVLnGX45xrxuq25wKmAzFsu2GGhVLa/vIdzIj8n3zE4GX0Fl32gfF
UXkT8PVGEUIPXv+uzDmOKwKgOuqrVe7MMQJO1SoayQgcyZrsiChmYM6TvJHxv2mx
+en70YtTxv6tAr7IkAmqakdHV6SwS+0OMcxYYZMFwaMJUNEqOnXZYaufzkikiXg1
JrR3ZHjEA4jDKt2C/ekR8fPZ5inEkpd/UnnHfblZVhHOFxzwLyX3jk5ce5WyEI+v
aQfl/+0ybtQ/3+QkQgoHTzRCqRVrEOSOfbCtm7evitc=
`protect END_PROTECTED
