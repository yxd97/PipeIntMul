`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ziSn2zIW6peqTzrXeffHIs0otllzX1MdU2QE4o8EOGl6DZvK8T6SsAOs1AFWo9RJ
JwgHfzNxR6vOh8ZC43HH7btABb6cZG5eIDEHrs66GmzJXeCa/yAhNKDnVMfzytrT
JXHYxlBGiIoq60AvtklsewAswEGgEoYIwDPBMFt0/C1ig4/bZVnIS6ZqQohRJE/h
VKbbI4rQ9knseaOvdYbEi/isa/M+eH/GVnIpAmzbV567NIx9JFhdB2shjnokhdvK
i/iEJvVAuqoEAFFX4SWqoxj40pjEOHV73vda/zzZ36U/8a2Uf5/BdWYq50wets9z
EL93BHt3y5FfBK1aN2qZHQ==
`protect END_PROTECTED
