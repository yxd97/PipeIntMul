`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vjdODfkNZjmjbs8VCktmqLGALKXad0XgBA4SVdz/LlnjxnbDewjUuZ06CuQ0xCsT
jgMPQcSjnyBf5eIi2nlOwpRtKfqAAq/E36hLdVPQ7sbQ8uPJWSkzUgAoogRhVTXo
zaDc5XasSjBNAhOPJSS87uQNE1ByioexNWi6VUutARWUQyNYOFOvqnhiy2wVz1PE
E+5ad+BR/0qMFHPSyb2ejcS2wsEHw52zcMo7I07x8yJ0PsWmc0icMvMFI8/bRc0/
y09MF2rc0pFoGwZV5B68sg==
`protect END_PROTECTED
