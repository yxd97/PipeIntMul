`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8yuVbS7v5IenlHi3NzaYg026wanAJ4HPNE8zNUYT5ZYudMWYPRndH9GQWF/0KqB
pD61d75vQlGLQntDk+PY5RvrvczNa5+yKu79pyxl8aiyTzyltNW9NUQE14rudygd
wtslwGU95CT0MVoYQIcjbtZd05jfnnP4vT54x/Hgcv4P9DDXqIQy9g4pgFNou6OJ
Oi5yzVhyf+82kqSlWqdKlpwvWcSTg5kcAWi3PpojX3ScTQLZa1+ZAUd6BsjnVMHd
GVWGMg16IVKqzoi3fDPjLQa7GPfeFGVnrcDFNUNynwa5zKAMrs/9tR/uyeXofd0Z
j2OBnn7eLhJvMHLv9Nu7sAW80K9C33zSIEnP+bigJIy0uc/iHgiq4xPzoe++9Z4O
rVZ0erf/wYzfptFdSBJgPngFWBdFu5C3anD3jDxlkkAwhVnz8SZTe03YZ4gBoVuf
ADvacvsdCVPpeE49fSnK0aHbcHKMDPgjgyzr5h5zh07s5zw9C1ffwprbeYEZe34K
pftPGzVmwKGUMlX72LrYZo1CoBZbMZ1tpritLz+v4Su2TDae8g7aeyiFoPe79JR8
C9REqyPi3IhHlPSmEja0jxWrTi4LUtwGYxeCw96zRX3ZswXscZuQOQkWbts0K01Z
vF+ha+KANEWWbHK3EgxOUl2i+FOwuKwVzyzeInRyakXZ03y6wYYBs2Xem7Am9QHQ
BMUmqYXpxAsMx5xZQlek34NPdBnF272El5gx58SDMZEahuzLSaKH/ZB2hBttz8br
LP5VX50IKPTFLZENUMZRkmH6mAp7c0e/GhV3Kcxn90o7HEdiQ+PUWMYaep3+aGyN
VDqWaCqP4Qb0qBjg3Ogv6mTw0tPzNu5MQWSGJ7MQ3hOQdKMQ4XpohlGAWqDHj5k+
rtLMa737CW2DDCyfdmIcWHanu+52X3+YJaCRpMd9x+jffC/RbKOizBtdjBYGXg5r
aPaMIPX1vEhWWl8rFqSoPk/vA2vtxoWT2cTFD/ZN07eib6JM+3SsdAzdulqZbAve
RZnOzRvf1B/Q8HtPwq6Wvjrjay5qxDnpNU/kLFFYgf8PK4B4/kiq+WR1Haa35CTo
CYp2NTzsN53BYnNVa4wmZwRBfzRaGpxRWlQ6nmZGmRI57lJhrMZdvWqtdMJk4IgO
WnDu1O5jeMXXF/Ui4Ov6GQz930IfS/vXUEnLTzb3IcJk7Bmu1KC9IBxMrbnOZXHW
QIn9FM1ZQ/YxwU6lnFgbZ6BGKcWsqD4xjAR3NJymqqqFtCCXGhLYaOwPfha/u/e5
9zwAtvzNEI3tJAzPTHbmCUhOqRdjjThgLyfy6lIFzyxCl0rUEBlSyfFmOZIgHkK3
X3r/usmD66zu5k/3D2x/YSg1ArOzH/jVLimPmlSKBvU8Dt4frKr4xOmpvlgEjQYw
40zUEd6XyVnT4YrP3L1+B9aZml6Ga/AACPkKCoTN+J+69ObvBXiUkexN2T5nkFR/
vvmGMgezuAmhaeotLcU103QF5bz3w4KGglUh5wRXvPEDaoeV6pYB92aeaduGFHAA
O6WjwiKcyn5+W5FO99uCWdduDPZmLgoh0TKF9kh2ZVqF2LJDKWJE6m6eA1S3rqn2
ltAoOfo2zTFOgLkkijbNHo9CXe/yI8BBY/RIVwsuEvqlWLGdO11X3HmBMbhmMD4O
c3uf3pzJ7QffPromYcncK+GrmC40d6pJPwSw5yYSldtF+EGD6PVwjlJ6fok2GK0j
C5DhxraDz1e9Zz6p7obFGHsX2uw8DEKIB35ygsoh8h2ce1mJPNMRMJ5pB0LVMuL/
iKQSnUpQ9d7JcYzl9Qtnjx5GGCimNcNZGuZU4xD2L8Pnz/IhHM8F+FMamjYgg5D8
0B9jTE7GU1A8axMcFo5Jt0Eb6u0aAbhOhOjx/Dt+ZI0qi8XItfFc1uWLCqsUfhXe
TAlV7P0ZEuu+h/kypm88yXCwfi7NTyNOg/kMzI6W4bdGGtEhN4JiKG4nmVMNeIsA
Skqs9COQuorw4UwDizT239i8f3HGtwNDW/IliCJbO/G08ZEoMOB/p3w+FNJTARLO
WejthFi6UMbxPsI/0hE/aI4uEY6r9a5HhD9vi53ZiyzDW8+4x2Bpsas7wra/mk3x
2e8HilCciXHP9vqn64Jwr4Yf7kZSaQ9fFZA8/YfwLQoyu2gmTxZZviMfu/FwNj1E
GVCr2ByGocNZ0DTxLYJPOeQziIAXXbTkOv7dTy/3XA4D5qoF+tz8qG2km4EPF8Ly
h96CVq/4jdI0+/pnQLlV/FeBbS90gYMj+xjQ7fs6AALqtRQdN1DSVwl3C3IRWiZ9
4fFm0INnYhOYeskrg0nNHM1UjbD4bqM5NH+pi+EtSsXMDmtpRJCBGYPYjt8cjC46
4Ml1ZvHBkpAFWD6A7KqjExdXzU3mCnCTP9F4fASzWtYodGw6sij+e+HFkh40sW+q
QaEi9y0uQXNjhml6rkUZBoSvk67hWkBgDmwHUoQ0pxd/ODYM6XnhJLEe0yVUT0rD
CY8+nFnjjnA53YnlQ+o/x2ivyKDeBGUqXn5vP4tiAY1ThdQJPwJCAbf+S12gHvOD
MskgKeCAhXfOA3bZZfsm5lGdFq4468tMKSb3L8NVIJ0CLs/uCKfQZjTHxYoBB0H8
4zfA17WHHJZc2SYE3NmcSdonrpLNEcyGjfCGcXC4yJOBt3JvyxD8bm6goQeQftPd
3gB/DmKCM9fHdHRTLByenY1WZVM1Q1EjkGLthvyxtS2LgTX6t/mirmETOeh5ftaU
byI91EGcYCQZFdFjldnHNX+fFX85AZq//Y/w7Dvhm8VcYivEwyuzcIeQ1a+zXf65
UimSHHz+uMWQ1uQlIbcpUg==
`protect END_PROTECTED
