`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wdw0sNJqthiCsIl3M1OFhKeAMBHBjm9I/uFuxGYH2BsnKtcmXXl++fLghs/3vfAf
zgVLRm81Yf9VpNEEtlRgXPYOivgJvFhBzDHUdhgjakCa988d2HC5+QO+u+Go9gtO
TUhPURr/zgDHFa2iiVpxS4Men/l9aPSFiNLEW/lRH7RXFcWDncoE4mNA5swhhhPT
nzbQXv1gKtD0+yhNsS3+K1SDeveg0aloCcsJA5sN7ryLYUT9650GZqsJR3vkdf6t
62ME1UflO9uLUUxSi23+rbpqxFhwufdYwZm/9MA+KUFywkbgZiH9y5k8YJx1vDCO
`protect END_PROTECTED
