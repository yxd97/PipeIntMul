`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Te4W0DqVTUfFj1ZQ8dhP/0ayZchqIAc9G3rzuPg/vtMjlG7qi8RE1+EsGnat7o8B
tEZnSXSXZV31TBVbZ82DMMxcIjf/4rEkesuDVFoJGiuCBEVp3b5Qf2BKhiorDEQ6
lSd1yNxqQMADcNJqoESf6mnDmRTuiAWuEPZKPmpj4QdnDKngPNSDIRp1maWDDtQo
aHBDOWae5dXgmlCMjHDcxpTa2rTcrMtMM1sxYsFQ8mYiRT73OKYLkVfeO+QE2aaz
CnyeBP7u7+4u5lrlIZHy26gKxnUpZwX//Q71XcZ29o9XwDPNL/8SiMD9JdN4yGr3
b1EtYTPAXusmlA3dFbD+eZHyvJFDkUJq6vQnRFn7LMvmp1oSjwEN+hFDIfi/4JWq
SFKg9n8tMYEDaiq/TVqvKNGSEqHGtGQxwNOz0E+2zGOErzePVLXTKupC0+Pp2ALh
qvgPOYzu5luiFqlGKcVpBxDTXgwbz5hvEakvkwZWwP14+hdQ191V10/QvovO+piu
Kn9KJQGsn/8wa+KbHeoCFNhphohzavjcsiSrRZ7LkoJOnvmYfkDcxfmYbkIOtolP
8f8ePiK1b9kdxTXExozxdAGe/GTe6TfCPFzJ6A3Wrfn+q8vwgGJdIeICASpdjAkC
O1MLmi6TqHcBR58Kmra3xL7AIJUkH+iHe4YJCvL69Z6D5UkHwHgOCfMUcNroUVwF
LIzpba87SO9Ld8BGMXaR5LtZov4UWGyxXBJrS8W4M6WFPtzl4JFeJInkxsr36KVg
koZJzyO4NaTUuFOD9zWtLOFFOXZgcS/EnE6+m57Xcp7yHHdOe3utf1od972mt3P2
1IKQ1f8i8iyzg1MoZ9exHiox6aTyX/03L9hhALcTh2lLEYkWPaTNRuckHZ5XqaS7
/yW9S3LzqMUBrNiTXKTjV9MudjbyZEXSz3so/wjJhHAV9a5NCIAACTpx9l9roq4e
wzlPNISpCsCtuEbFxXPQAt3JWL67zTykrJs0P7FDBDZ9Cz303KUrG4Mk2heJu/ht
cmIBYDhO3HBH5vdKDshxTw7zHmF5h/Y3lWv9TKmg9Wk+5vfWUZZjaDT6JQCbB+xd
i0rLqN7gaDIZXpuRueT2YnALe75E9mkcIqodrmnUNRKhj/o/mY4VQcLw1qnSzOB3
rnuk27mLCIjAQ20I1Pl9XWM4PidaJzayzjtJsgv3K5YsyclJ3/LBKAiqPwo28fvx
XGKnGtH4oaDK5JmG35qsOx7qphcWq15i+x7IxOxq5KiWBhBTNd7suaF+tjBHKfHP
REDBHGwytD2GlpYWsHlH7PH37QRlqqre+khCZDaORDdjstbgk6B5s9JzxkdVQC/q
yEb3U7sDAtKU2Yg2rs0QrSUcj1WHhGVsZqkfRX0DZBCWmIgeaBWijZGStSezBW60
Wq/0dG0Y8qO8c9wtCX/FP39g9TxfOcA71R129nxUwbvohHdnT9sSBgd3xL1kolok
djmElXTHxL8bmTtjJG1GjPq01SBxl14Z2GTxtabbORi2xKW2LSJM8toe9fUGUevT
M3d+AVlgVMmesC0zl+RmD8IMwXXCWzWa52YBlUlMZna7mcBX0v4kmjjDNdTaDnYR
NAkYqMvbiFsOtZr+kSVWmg8ciiY2e7qdrOTOUwGIH3MGLJX4+BMS6F7z7Z36z4Jx
j+u/LunQ6zE7RKrPTUqEKAPqqd3DPPIrhVgc7WjoMSATkesmGvkISCed5Bd0sLjr
pwjLNfZf5pwDEtPQ6PaFcR2ffB5nPYM+vMgv+JUyAMPCI/suhHXWGDZrc3rByLvV
P6785VXoxul1RbVUEVt7cDp+t43jH/gaWr5xaoR96zRhVhc0UvocmJpw4JnDEWHh
28Q8zQghGaV+ge1648lkEPasLlH0mMsfZhz8MLlrRZEZnsaJXm18s0Xp8TKg+AgZ
8Lk5VKoeDDnI0Ta9w57lGkB2gXnQ3PtKgGm486t+uTBl4y3L5+/61wAl/7OTillO
4fxolvjBjltVX1q/PVw9NnrOZCViWSsLWj4IAWC3CXxUNDaAgjlJ1+XvtYoX4QAP
EnR/nxRGLTzG82QLh6FPU2uS/eilAaw8DlSrQwbLaqcfsS/egBJWyfHs/e4mPhtM
V5LDBDxQ1rCBB3E8e8ePgRg/0I5SDJnY6OInMWPsyB33s1s/97YIvaiGOjoQIxpN
PmoOabA55n9/ahiRMB0r2N79l2N8kyXw8P5195w5pFTg9PaseHsYEpSRZ76iRdQ5
W/MTYMEBWg3V4QfTqVJzh+s9HayNcJINc8pueDk5me3iPu0BukB2GZ63lTb3YKuH
C3em81vCN2Vq74Mg3gXXkvPS7kKCQVi/W7opZjH4CDoN29XbByT6skuRJV6DgqGa
c5Cemm2Eq7EmT2Kp2M5HORxUS8iRDG2U9XYoyHqigI22PMS0z4H/ZV4Q10cECIgs
Vv/oqYdY5+67KS1IrP1KqoIy/SIKRq4IakjgkibtSjXf2rOK+cqGCQO+ZWUHpuj0
TB1Pv3T1LNtYSruZWfXprmEB5nYhsXmUvki1hLjFppi68jqna3XHfHpwvaea4wbS
etfdOTMdNWoHdqRtXSbOFJ5WgDpk/+lahzDnMm2c+UJH11GmXEZ8+quYeQ280cmI
ecdFt8VU86YRO6jTEYVzfH7A3umZ0RXbRpI8R/YkeelaHLLEyqy3mLh7NvBV91Oo
dzp8PXzvqdP2thH79AFnULiaKYcYfrDO/gZNCWXn1AR/wu4xeF2MJp7RKmC4fKO3
sW0N1O0krVxCm/3Qc0TxeAUMUPM8FYTNUWQopU3sgoWjSQkNXeLgEkeOZF+d/fZj
ZTE/ebGn8+PLWBJ359VV4E4bN3Q/L8tXSOy3R6rkYcxFtay7yDonxFNCIDLB+5R7
s5xuhdfGcY3PylCgZAIFfVqBL08yZnJGnQTHoYn3cMPKSbHuaruSM8VD61joAbcA
sHQ6Owo++7wF7rP3vME5yiWZK1ojbToEZP5nLuRj+DVs3DGT+ddH9CCZ6mEMuwE8
nQ2TWvgXB3EOdGI6coVoUmnVAOP5WiTGe4c5N1o3eUjzJkSBeaAUbcvJVRCTwpBN
Nu9e2lP0MOHoMP8RT8cbXE1d4TmRIZ2jIQC2EhhGeVAfSjTSa7dDs0iVJRI2egTQ
wNpcfhMH4E1W/U8SKQ7L39T0ncBH71oVARBRK/6C6/SE2PKkPHg+1nuZex9t22be
QL9OlF32K1jEFgk+Nh5VL3Q8l3X65n8FFp92EaqKOVQy7/WbjBnbuKC3PFymMywd
PaZxxPN968UM17fFujnT18H8ejBLkQy2J6YMllu/jw3JlTFvg4Pvv+cbvurZ5+Er
eYzPH3lAiUo87VD+XNxq/Awgtj1efJlMV/bxf/8/moQhMh6HCJuacZFHQ7F2m/0W
8JK3lkuyWSVo29PHz5Nmg+0zjUl3vzbeKhBNXxhppb+FwASxjlhJTrkY3vVl3vIg
6O51e3uhaOhqzWHjpdlTEd3KVupSwSzGH3ps1dPXn95DSrqxkl7ps/Oue6UWsIh9
pocNossKxwfUnyvTS/FydCZzy4HZngdwM09rUhI29o/s5+edS+5zW23YNrfiKdr0
GY12M1Irj8cBFf/CIoLHCZB9aIHRId+Ky7rSliKBi6cSNVJO7VVi//h/G+leEB33
2xc6+aPAP1Ad3QvMX8dgziOx0kQFYJuWJPvQ8vP4kfFr0MWuvAr+czWd7o6tr6it
rA5JloHbX7wlg3yfdnDpaAZYI6DqA8uEtMboeEAH8R0yagE+43mxVw310zF+VoO/
WcXq2MjVim7b8+17p9AAfs+1S0il//CuZewrIdVlo38MR6ljvWa0P/+DP8mAA5+8
DEetM9F/WVZzuM/IDgoIciRKNVFwJpFJePJX2qoRPxU9n/M5oGNsQGmuyuU+xevC
MtjXK5b0VUqHdU0GGtMFbNb4FjDLyUPwSPkgxhSt+FS8oy3rJM3bdsfiSlDITSN7
9iPSvvj+dNSJYNAn/NykFQZd85+tKNLke0YDDbGkhfUAiaLgRVLBXYK9TYLqOAc5
W0WPX76CXhgDdsW1Ds4ZGiGn8nLWga4iFljP2gZchdgcDjM/YSg/x3x8THpPizPR
EO46nLkK0xTUnKW8aHdKasaU44Ub6Er5vpj3cZOCvwF1ZyyBt8Lkzwjsa+6S+ozg
D7sdyagt7B5MzuVGYmvqc0DztR49+dXbi5S54tPwm3JI6pJBhtfz94psbczXAVjc
xkOe9X5TIJYYw+plZ+UHYNADhvKusnPGMgq1NdJjcU05AA1B/iQFa3SePqrgv1nv
O0ZiVYHufmYeBGKQMLxvCeURKOSk9jdyYRWhjZh2I0nmPV6qoKaMUCQYr2d1Y+bC
j+/LoK0lhNmJzImwHOMv5Y8mWNooFyftUWzuzZSDVTlRZh9m5J7P6qx49D2LEqvq
3gpuoqB3nC0Thllpn/f39KQgCJ5zO9Gi12837ZchgwTcNguOh3ezUX7DLKaGy126
OBnJtanEVofjR53N66e9tkOkeceA3PdK/h1u6VpLcYLy2XyNYW2Y6GzHJMweYs44
RjmVC5F5LgWS5POwmdI9VNF/Glm543dwcF2s9y+MrCg+IZ3Fiqv7dTr7JDTf+8uX
sFkuHWUxDcjuimkFs7Ekxg+AftwbkChBuE2897/3pjCirf5KBmU0KtV27R/9q/FM
qBqr/V0KNTwrMhFCguDvHqreR85AxKVz/nU6PohOsmdFDlBnTkyS+1wBozUVPlCi
BFqaARdkbIuupFJXcfowmkHDna/oxbia+P+JtaXtD/ZwcwfmFPdhMm9FDXTA7vUz
IIH101OIYNxDlWI7ksqgJt+Fnbyo6wP0WEceVYkGxgFhARfkWnVsM3E3NwRLaJWM
LeHD5dZzgJ7UzZER6mLXmxwI85SHsdWS7LYySavrFTrF7Ue8P0ZoUvuubt9K0jjC
/FcwKkOqn04W1WRA0knNy2Z20PKxYz2XPXrr3kyxSo/zFfElRnHCd6l5c0BjtxGP
BUxEXP2M8YK2g+zBVOvF+EdDa+QcM3bRIUF2aXbpgCBUkSQxqrBWihfvSE5XxFCV
6usxVWUKMfINRiuzBDT/y6KGff+wQEFwAjtetDevNAFz26kQ5jb8iAiKfOx0a2mf
T1qwcWbIvvJZi35UlGYnwzEuHqm5xbQxwkDi0HOt2P2YzleD2s6ohcyLHMRsiaUK
uFdOOBjqdRrK/exJFFsRbEpelNgxxcIEPZzc+v37pa+BmqRedMYI7gz9AcZWCq+2
423SYV0Wmstj1b2OkpRCUJSAtTM+YG3xF8B6zUk/BjysTzWclM8oSdV7TvKZZJnK
yJVkEvMZcwWebYALrb9OJ6sp2hzLnRthPtkFZTLpZxiFSRFXwwrXYHnMHxhkvz49
Y49P5H4EcJLulldRX2+8En6Pa6g3EnFkFz+95WMsZyHdV3cTeZh7IyXMi57czmr6
iGfmZ7BOqKO8tafWUcZh8kgJedP1NH/8J70YFXwnLyMGMixZoKsVeHGlTZG6wKwl
b7noldOEoEMFIf9KNbCrZcHO71Re/uW7zrRYwjjwBfecKPKYH+M6IKn6s5QHSP7u
Ey8zFE2eebrj0/NMJmXoJU9K5Pg7QYsEDKG8QmHdz9MFCKMF0+OzO2C9q/kbiNYt
WLxuO8E4S3d3xa/PI+ggOSDfzAgi9O41ZcXrLnXQ2+2FP0idlQPNKaex8i5IRGlk
nhcAtO7/IMvNTk77B9q2MNqA2f7N79zx3xPMqWuIF6HSoL0KUiyUEiyD0PTVwDGI
AL3t5+jRmXC1jfXV+ZS+1Lvv/MasirQZrAock5WqQJ0lHjF4GvUFF9Wlgifxz2Po
56HBxEupq0KkhLSGSlIKg6uwarfKGj05lkm/syNexGFNESt6PkOIR+4l/VxB4TV2
7PkPwp1SzPpBsORxRB0vzpf18ijsMyQcS5fuiW1NKsRPC0w/ljk/TABDIvHc0fHv
ggotV+jbJ/AeRIg5NtLkzOF2QP15XmqhJCF98+b0J8lf7w7gaMyMXE+AlWlIYwag
1qx/3Jhexn0T3UNIi768xlkziWqZqddCe32eMobECo6IMXLhb4jZHlnGVgltEmJX
A0VcedNNRF36Iut+S7BLKbszp0YBLphIWVjBYT4xOUubV4mtPfWiXwAdrv4u67yo
/TdDjn1+kX+/i/7HAl2qu0LwR6OOcyXzQ+0KzTr7/QsRvmQ8BS1sHN4B/5gtMc0Q
hTgJvylXOv2OwWzs0MEwnPqtT+FzzmhGgzOeMvja3Q5+Lj3APT0ok804KeIIA1Mc
hSqcL/kUEp7qZaAXcym2SGOIBom1WLD5UQsllJiGsZn9zqj9k3pzjzsT/uVkZVTS
B666uYfVaarse4o2KHQ+ZU53wmaYNp4+brEJMwjyoqUpvSNu8Y7Vw8TXzDQ7dHZg
WFGEon6Y4GKmHEdgAXXmGxGZcI5rYINS03QudOKwlBig1Ilc3B3xEbkU3CnVX2en
epXYOWhsHepLJRZgkTsxqKqsgb7sscsObMi0n1E7rQVT4QYZuNIw8INg/c2DpJwX
rj6mWa3tDo2xOSUUE02KD4Xk2J3LMv5wuwt8EcavuDvFV44QjFoLEViBpq1OUPDP
UA2vPxa/gU1yCIIv99twG6xy7Ls5f9cHelma/C4Iq6XChuAbu08X0RgkxS5j70xy
UkncM77/GT0u7PytrPNDR0x7yMc8IZnTSTQ0eGXM1s2eSQ0iqbvktarcudE+7LkB
/N2ta709JwIBVGf79fH+BVpJnKtZbVr2hx4w2vIe/SAdee/sA6GPUZIbPrgZn1n0
IQi1+E6CPeU/SIwJUhQLm6fyuEU8gwum6NQnAEf/o48I7oqgb5tFo9r+ZTalr1wC
IkEosE4Vk3b3pYSaYuZ7uZw138LVHxh/ayzZVP6jfx6lZLp/kcWYDqX56j4t778w
QVgLtpOit96q0eSYCFxUYs1kgEEJjV1rXRc6iexJS8y99jgjqPBeV16qOgfV+zqZ
G44KfRlpSPHANY53zG+ZCl6LwHFhOKzL+n/XCnAexcX1hhMAnFjvgteJc/Ve0ADT
yQPzCrJ/Y4poEhLa9rtpDIzLBH7CrsgQmxl2ulmk0QqUydd6pTbjpJ8NIpC01qfB
rcWRGCLdRjUtns51zvbRlChngp+1QWGZzndb1Y2+kGoqAIpJW02sZSQF4X/0ZJba
Lt0/TNApaxXUMGoJNxahkt4u7uLgR0ltEwvNxhLcQhEsXbUods2KeuCgK0+o1rdF
ppOp4qppK24F53kEpe1iDtHHYBTy6kUpczoXhLt5+sGYp2Rc2kt9nF6X4HklLnQP
PN61TmUJIQCXtjWMKTZ43RTgdFgxSHya3lwJgTT9GNjJymK6VKm/LZCvpUTm6vgW
csreafHfGFffwv7E6FIHcBjmS1vKw6tCOWdVoSPbpVfceiBCUOEosoC3aPhJeMY3
SQbAGhIkb9IMGBIpJx4UWv7+7g8xNEOTA/AHFDESrqxdHSQBqHA69V5+YzyAFCO9
ePQK8b2qq8hsBPSYJuhdx0qZyKdNaBkddlcC/eJB9epbOpDQwXxQ9hHYZyD8e37E
qiyT1+HLnfslPxzwkOXbFBHOk3X6mNI8vXHeuNxcEAlbllphS2bqrduirnKdLXqX
Pc8IvXMvYsnQnDAiCnHIOhmoKocQKF20UviGcYTE/Ieja0xevoOKYuMEGeCu4zSj
XjgGHv53w6iSXOCiJP7pzMO6eZ4zvl7QWcTv50L6umBzOzXyJ0A4KCJOxY5pLXvr
MabImllZp/pTTa3IoEmRpkJWGq5G68H0J6opNN8KCqs5/OZKYj7VFZQxK7xLaYmV
PCelBP34mX4oLsBLxF6B74MBI9rq/Illm8iw+XTEX+g7M59x7T5CKqIAVGCHsThh
jEy1QDwSYyJEpSUo516xK26zEDk3RFXO3PIwjy1m8x4zsH75pMK+B2sd3aTuTMgW
qEKLzeJH0irUjG2VzWF4lan04TWEud6KKphKBgzhm+y0J5VxVYjN9mehMQhTw+rk
9InacU57fTMkJN/6RDk622tznWPQBFKfuiVxuSeAZOwXEGfQ3TuWqcvDVZlDdws+
MIhOnkvvYVOXjsYO7o05PW6OawVdDrgb7GbmcdSp4Z6JMz/yVfXtec5rQ/olAhAL
RKLLadquQk275kT5i1c/GChJAoDn6G87MKsMXvNwFGbXx91OiQODCUd86iCi53rx
NejluaMG702n/GJOTfCNbBox1U1HnDiZAtozTnM4Xk6htq/yKjNkCpPdS0PQHsp0
YwW1g3N6yZXd3K1S9CRfHGGylalj2Uh/WKNf0uPZb0MU8cFUcLuZGQ80VD2aHF1g
QRHp4rPswqxSL6Uk/yZQyjHIxyd+VHLg8kqvb40pq4ae8he3yAb6wL120bBHYnOH
qgbRPKhSEtYLYVRdOMfSLUKBcuFwhOyV8WGWJ1zAUPztnc7UlsA4iSuWvTL2Ml4T
n0xj9Cq074U1BDjlJRqrnVNf0FnbI9ceLUKa7tfbW7+96UamuK4pLw0oCGPMjzad
pWBZEC4gd/zAhzoE/JzUD3rvMpW7iAGX8YCG7gyV5HoxoMIzpQylMQAuciDpD4ga
/r/cuJYn66lbcJU3mimUVcxsTg/X4qpdcPBrhvJBLrQQo80QO1LFQkxlDkrUiS0F
j8zQzv+PAsD9iyEyhk6PlMfecwNWzwmGn3B2Fg6tohhZgc+619f5vQw6cVP+0tar
Nuyi0YB1cBbyKDklEEPEXWIrQfwcEvvGc4kODE35iBJzP/Xq4g6fEKHk4N40eSuB
H3degDcgAvz7IYBau/0ehFF/r24CGGU6uEHPfq8TzdpCBiByMQLGUAUsuMYdtvbE
wS5E7f66nUNUMRullG4Z7Q69+qXpwaNfF1OHmPXKS4uwQ1C/chY3seQb+9X2bfzG
beCITQV2kwjcpSocI+dbZuO/TAryc4MVwN578r6/mWXeBVAZ2mEiPhpuwaEiTg8f
oWVN3wYGgWEhI+2HITz3YQpRZuc/4gCklEGCY942GFTQZWUljdqorsQBOUP5MViz
EfGvrfOA4wqUEjR+LFRFLlRUMHqJxnmBgk1FCMuphcZ5YcO1dz9fEdzfPIKKt/sK
S3ZyTMFAErIv8czZvPcEURCM2HrII+vdR9nKQG8OInoFY+/iDilujH62mFNq9iPC
BuOqBUsvwBa5LjmpDzPv4ISmlQsGRKgxEN7R7y38PPpUTq+HzUaHMouFPXEkVlDf
SyHsoGrrIxn8FpP4GC5/0tAYwNXlGxiTa04UZVDanfH58YD2/EaxjDVfzoedGDda
JP34PChwn85g58lDSxNpgPWvKY4EKuvZ+gSn1vgveuXc0cGR7SQ/UCrh0BVuEt0j
mxkqKh2KJf+RjMImAtu51QzcJqpAm+EgdxdwFRbxVB/POXP8x7lf+ZCTvzKDHX3o
8zk/Xh34H5hgykaXCu9bTvbuwdhL6QcDKMQ6nLiApyuA3i4SMVHRxeA+urbPO2Ps
jr9veDYz4vtFA0QT91lp1u2xeORddTaqjQO96ItXowXKhBQnWir3u4XZ+BFPeguf
u3KljNFN9jrTW4xovKButwXHYxMdnCZCcz7F7QVH2Xa6aX7A2inRek7riVo5Rvfn
jQlKzOHTjWSCCntY947YeAi1d9xfoNKuSeIpcUrLY2cnKnMlqqIejw2nbn3TN8zh
orSQCcyfBkLXOOfAOwIa03y7uuLJs11mYkcFaOysFLpr5gmraQU3L5kr13EP8+4w
kmq8OUITrAXfSipqkizzrAjkpvGKDMyg2o3eKWBqADGkv8quTX4P3Ey1ciPHmlyO
nfcTKatunm+hAJdk1Hs2bwepjwuKbohp0nGkyToyq1QPiLsk0kWapbV+vKC/zZxK
fRXsdj1E01ysfSi871UbZoIlSJ87S30mHdB8LH6tH7NsrLIL2prCMGBniXduMK+C
eKjn0coujSKLbwKUq4Tth9041sYQNtz5pISo0OjyXNksvrCp3QmnlGwS6Z5EM4z/
AEtf/hXX+j1GKDFhGWJXHpqjUcgh1icV1mdWkKC6K/vr4E0aJLj7lafEnrq/3giB
cQaLKGTllJavdc/QKIDTxjg4ky39LKX9nPbLYwx7XltBOLjyPMMCywFcBrXlVlVY
Go2aTAKiY9+2PUlFiPOi9tMwgNU3oTfe+gVbPaBAi6B6Z2X5Blc+5L0s7wlcfkRy
2TfzfWscusuDPP4een3cVXhLfF4zEB2KBbWUzOSyDYa6G/vxkVB6c1XoFYtxKpjY
9CALlnMBx1fdEGK7ZGeN2Xhgc8EoWkWYxLhZL7Ic2Qeom4cK5E+ZEV1jRnhlwNhv
Z/K9AZUFXtI+oBKmQJg0KlFrJ/442svQwtPyAX7gWvIsSDWrv5E942jZf+ZbOFKI
Z9fB7qf8x5cCcaFueTl1Vuk7iA3hp0nEyvKYmpXfPcxxyKLBm8YZCB0nuPXcAIDu
XF4qiURTl8APbwiTYOc5qAiGQp/LrL0sjutynuRa0cP/EvbgTqLaa/deTE9jHTJ0
ksxLCVjwOUxlFEmGZJhY4BXBOLxaTdw4hy8qbnQKVL0eDdknYhMSNZlaWl4isTcX
uGu37zGgdBagZJC04+OpgUMilEivQ3wNrAYSln6mJ3x6TlOgRZCTYQbOwY6YwoKO
Mka4vlOiXDrtHxuwraALcyY3w5v/iQk4kXfC6Xgw8d5q81AA1FldrcgMJN+S5geb
91kAko84Isme0K3t2ro2pPKk05KFQG3Lt95bt0efZkyglDH4u9C11r+WfHL9evMf
EOGtsXiKDAA1Uukd+r+wkjsgMMXk901aywL+K9DaWs2PDJTQcYSHt5ffyYXJRZ5H
4WpGaP/LhCwKFLFvXrOoFJKFdeq3VicZxB3dukcOaBivsIHEjHuI1dPwwB2us5MY
0aFO1yU7NFt78jOx4nLnETz7pYdgNSdvjLpA+FkGB7Q5VagCD4BHDwEWPsd8Pp7V
zEdsedmBc01CybDmdj8meDvAAM0K+yFNQmbnxIsMgJ0bUNgGgYsYEJHng/YTv6bv
wS9kF7roQeMlJ/vjuRW+fA==
`protect END_PROTECTED
