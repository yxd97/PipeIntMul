`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZM4DaWL9+/NykZj6oCxuXMGOsTtoayAoR93CwSf3J/P0OrM/wLTj8g4MrGpz8Lxz
yv1MsZ0/LShL1mantmQLtGsVznd+cWXUFRGFC3lGIgqfvA5tkvUWWgIAp1eQ9smk
1n3X9LGVprwtiP3fz28FcaKoXcxewP9dQal/rW/y5Arm8m5gO6UrHa5zvr8Ogzvq
cAaXADTvKRLFQ06r40t8R8SLYcaBqpKEthNuU0n4sb8GpJkpcC3uX4wh3EOLdeKY
xnNwJa4/vEm469psGr3Hco9yXoY7/CwkqgBz3DOO2fQLEaUffu2QDxHVTF2LzGKB
fXVdTS5fcaY4jOo+v8EL85qkr9WaN/xVxzuufihZ3czEo2jzAzR4qz0+un+cSRVQ
O9HWJZnG0GZCGUE12rGTlWlw8SRdmgynauorvlFgaEk6mtuvF6NPSqCGk9Qnh8Ue
7UZ+PHIakSfXEQgs2dC0BTkByonK5YJuXGFgAyIQK+6H0IWtcZvK6EXFZ31MUqgB
rdsjF6FZtQk7pBWB6cxy4uYhVNuhGlfz63eX38H8+KtrdQl8JdCfUuZG8N46mLjd
qtq8QF3iaiDjOjRTxq0E6Z/cEP5u80fAgRruPhUL82I=
`protect END_PROTECTED
