`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EpGkjvkZNIxFWNmSCzxfc9zbNsBHhHJdnW4hGoPmbo+DCp88ar870FGwyFVDXX6i
ZSLPxA9Qx0lqTFWFUrpks0Qsf3at7YrePmBgkDCf/6znfa2YME4Gy0zaGcoY4JlT
WhXeQ3Z5FBOOyA/tyIJS9NTEsJDi5PxrWUzgEjoDbRfero7S0kqORH/bgKFvTsGm
jAWW0NJXBzetIRRNph0AT41f1gvLlo4OUnr30HVETpikFFmDkPjuPaE8oI/Vdt2s
tDlatxBUS8Txon4JXfR3ayPiZQHQzSNfdlQcb0ZDt4b9LvSz9YNW/cM5k34fqPY5
VKvZ0LZ3wlJXYnFd3zoC5P7FGzabXDHJrqtla7b1kglZiI/9pWNaY5jUrGf4tOhn
uyb9IkGGNeJSD8QdCIWAa+fphtSdnBIqbURa/oqGInb444rqOvdGju2TA2HTeos3
UfBqLVIleoA1PYQVFFV7tMeb8rPxZiOtvF7dzcfw2U0M5zC9vFMrkntgHVlsIgwt
5OBCZz3WaBSSMd8ENev4AOe8IK/vpkJgrh7Xm1xEqyeKRBLAZfdf7kcIUhI4taq+
9kWT52LDXC9swwBVrNGzxg==
`protect END_PROTECTED
