`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KerfVo1AKzFfkoivtAepfMYDV7dXB7BcjUaq9ZUi7g3V7Y1YCd64qNKpE/SyFWiv
je1OSAYemogOjDmWRRUWSL9wqC6Q8STFTp+2jbqvzyfJjhTLeB1aXU+IFKwYX8RT
r8jz8VKEbBdcSqqJ6+JmLwiZvlO5aW2dEmyMFHdEgnbnbYkGgzENHm90wniRQz6l
2Xf70uEHALqp5a92ybVWyIYsm6XF4wheH76jviNNRC/8zojWPMMnfNciUs2ra6YO
WrzLMtD4/sDdpOeYvxnyBir7j3zmLfQnmvDFBX7u2w7LNxUib4idmCVmK1jCNaSq
nNoBvpHXaUmJS2NpckWEVkPHqUexxdQgVx5w1eVCugJkayjuJIcEo3f4boCV4Wf4
Mo+FCiaRaqpsSlHSN3u2fF8qv2HRLh8CoPKmo+JoBYYw5RP9jNq2r1Jy/b2kFMbR
uNAEUypT4LRnsVr59dnDPZilOW82pDQVO9lzh4j2F7c7QT1p3E2k3m0PWXF1wKRM
HLUfXOsPHbZtFvc+Iz/tlsR2ix7Aj4yT7blk61UCwPT/oE1mXQZgl1lzyQGjGRmq
4XClW2cZcqYqUdNL7VV7tPI7AzBDO7u3k/1gmu7YIaNWBG9Xmd7D3dtUJTmyZwm3
zw3F74E6oV/Wm6Io+dyTuDVHZshnjB1EknFxVjgmK/fH+ffF9rmaVmNaoPjU39oQ
YAmc+7mAmsvl/cjXZyowvOZ1aIfzRSTZHPP3iiDctYPJXUmDCBXS4g2JTdyQr2QU
S2GWKY1YyB/plO9uuuSYGMzYrI9BuJmNVE3Wm5mIY6WkBW90pQpXDD9Th3Mx/ij4
DMzpaJ84+i6eNYRLIUEWuRH3yZ4gU/8gtayAOWdNr1WATlSXQ20Wu3l21PI/AdEe
rNsysrEg0swU8UuQ6MxIwhVB3HsXyQMYgMJ8E5GRtrtOnbpKREVUUZSE5VXGb3Z0
NXMn24UMIMAB8CkWZNOKT0Rlb2MO9lzO0HRNRgvoFokKbnXcybLfxksVO+8Vlk/g
M2NLcYDIpq6VpivwdFf6sTvSn4UBanlYabndiVQzNh3jj1ZOEbeH5wggRX/IwK1o
xjt4l72PJC0SeqdcBMEsaeHdRhvHKjZB/jOQMKjZRbsAaucYOOSOoR/M8KxrLKBS
HNLcLZOwplWWA1HWSJWnIpUBGiJ22nYA+s+PToAddXiHapCdKQlrT5AvB5kJDLXd
gbPy6+LTAzBCrDg8jeC7KkRlWR+tmXbBnHgUdTfzSejalvBvSHF+N5xNRt8ku0CU
20IV7hEZ8v7tB1eiz0s9Xk11jehuqEr6X/i2NmKbkHZ3H8IPdDo2/B6cOD2Ym8VY
GnF0VXJZV/1cPPkARlZmtPR5u35M7JF0TnA11l+HDbvv9TOFyziR6c8ue05eToq6
c4y1wygtqJ4/Jss8xR27YV1Sqg12eyji/TucFWI4sy08deK8QtOhZhISyJrK2rFD
pRNwP5ahe/yBVkRihaFZR6V7YP6mL6q6l4to/FU0H4yjpJ9eNDkAHtvb/gMBIgHl
D1OG+nDcwKKnZJO2+xveIgL1r7UyQSQ+VRx/0msHZES9Gvxx+nez1raAuaA6F999
hlqt2vjt9sCapiqOzxECTcBFOXWE4exOx3jj9hH/cZlfI/M/2BtUb2CBj7s7oaRW
P8ISLxH58i1JHZxd3b4BdrQzfPSk6scVd78EAcrIp+A32wIkfAsQxmdDvPnXY8Cm
oQEXmCTUv3f/rWrazcj8tOfu5Zql5vCIQLx6s8yO+DE12ZL+Prvi7ItpLeRE9W8j
kx4E+W8+HHLNZZj2h0re52fvqOrHp4bYtOXz4uumfN1f65zESTKSlhvEyaIDXvuq
Qovvqe0cY3zPUqeO2O3yngtB0Rrd/+Qpdl84ws5WNTG9xZfpOU/XBNqA7fH5/ezX
Eo5OTUQWJ+CCwqfKwDbEMn7Z4SXjGILYADLXUZxINKjfX5ipYf9sYuie4lRzBMyv
JLRpJMpvl4VyZzO6VqYsdYsvgCM8+LuhJrdKQCW4TDDpbhpB0Ch26lCcFgRnX/MZ
0gOM/o1XImrbrRhaUBpPDq3i+dw5Ux3bk7iTy+/8kMdjij5ISjXy8yBTPdjvo+sH
MOtkuAhEmUuMp0eOOkTV9G2L/PADSs/cm4UwyZ17bn63dw0HdDCui7mKbSnBV61x
TKSipoHQ+Bv4JfBGP4GyRg==
`protect END_PROTECTED
