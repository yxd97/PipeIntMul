`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ji0T+mxwpP9WvmAdNBM17VAerzHtCYaPqKXcg+BpvMMjybFk2cEyexIeiTCacE2I
uz0AP9lvRjLDOwEZPxIvv33H9tOg+UvRN7DmoJUev12ndUvt/KA9Wp6OevR1IpRd
qjsH3bTeDzL/mhc7bToWFhwLX1V+lxAWuJhpLnauEeV9mHRKHvDVJ0Bi7gGXhXx/
7f3KmQmdDwdzzXWs1iMMw0T0/+ib39tY6vmDNPJZKM0+wfjTMIBiqCJh7HV6hKKe
NYArGcqtnVQ8bM++tjwOM4sTslDDM76zP7dvv7XOdaKzp1SsVhUAeZ7FSw/sIb4V
TfytYTrm23rqbhY88WyGC6ryNNLtPel6+vrfAriWzQsmKHUldNZ/DZzCNvXueO3G
cIw1vQZFwRGbj8lgg34KvgWcSOPdzOa+hhz+Gp4N8ChvvYJ5mDuLfYIzI6WLzO0O
s/AfM8OHhD4w45HH+7jeojiEsIHiu44s5xFvUA7JvfOON0KV9UEaMbdwugwqmnGV
Y3bkcuPq/Uk8qAszM8x7+c+5rxLBpdJQFtFLklb+ySsHjCi+7lNPNRRhNemFTUJF
hFdiXPBimE3u8S7amKS4aNHnrVAXNKoLnsz8yRw9K54=
`protect END_PROTECTED
