`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KN6iHJLmS/eLuFvaaDjLCW3BGljyyLLQR1GpheyiNAe0uSjffv6MDCz+KDSCvg+e
qT8MOszxZT8tYXkpjEF7TPnsdbFcJ3TVuGQqBmsFPHK4ErxPTWOfdvBqAyQDPguV
k76uGCLcNNqb7Q8tgntvww3j3lGqn18RE2xT8dDQla73Ouz8Cu7zHDYhirHJyUm7
WVYazGhxYo8s0FhaFcyfSX5UUlSY1bDWidmvUWnDG6ZHBnCwWEt3Usctx1vRn0XX
edOqtmLlOs4j21LCybqd/sAExtsIls3L8iJK4HZXJpiO2+0Cl/q7AyWHNrKv3Rdf
gTumkfgaFgtVcjkuETrR7Tl9C2ow9K5kAR4iKVPANUXoiGHNAprtIJTLQH9GJixN
GqZRlNNKIBJ1XEAl0xla/wYEddlOf3BMZ4bOI0il2p2rekipRlYKENm+tGLRHgiC
gbxJ4UKwY1midD6JWkP75yRgZZn5j2h2KKlRKd35BVuKMCvbLp1cnI0TrKWWI+zK
zmVueZcdxHkHG451tkix4MhS/m4HjUDEpWP5yR6VFEtwg4G8qCfwm84TPX4c4Div
nN06sFpa1HC7ZLPfXhhn+w==
`protect END_PROTECTED
