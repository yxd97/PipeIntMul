`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdyxVREeO7DEbq8t72DDy/hIozPsIDgmTq87h0vWSj/b8vEhGzPR3fqd4rek7ujS
W5TVxwobzmc4FqubXrvbo2VAycswXpPzXsFKRX/3LAlZa8pggwvxXyqNF058w607
DU5ys9pZJEhUyJULy2bJLWntiuPtAafy1e774PAlkkuCgOQUAm2erBgRc3K9AF/v
absU6ESKaqG5/Cgb7twwUd/C2x+tZZHGakHdrW7ohi+21NYaI9MptaCDNdy6sNB/
MYVoQON6otBD0WeJSYd+EBVj9fFauppyf8izF9mcwBqYY04RGILgZne9zAD2yQgo
FNRpNzqZfF6dp+ERtlVPh5oECH5OSxPdBBiMjt/qvsvXC9JjEcnSlDtszYn497+E
mT95ue3pS8wLoFuXQlGVNtCZsJA0HCUsSW2d5x6jiBtADeZJldVI3jvswcjpQiT5
y+IIXve7etvQhfZtFLQCCJDfNDhsX7mO0lCfsfYh2esaFd8pjGYaizFp7o+JKNy7
Xx0QQsMaXuFnMCbcEMHrn5Q4lNgh7hT248j+RyifXK18WmvkWHsm7cdkM3EAbMzl
qORNTU5f5sCJT+zmzXz3a6I98OBeJpA70E3gyfANZhpyhRQyYg24mTY6oOLi8JBV
nCFRQD0lwRj6lelbs2VWG0XY7i/r5+te+THAuZkwb10lmFces3VLKZVhhK+RxOAa
4H8J3bLkBCXLkOwFKxfDnwiOBmTBC7rYRPwUBHRkC6IrumfYNTJVKQeOr4btxgPC
PLOfU51zKGxEQtuKttwS3l3cKI2lNsd1NzRgrrI8jFSUJBIY5KWKJpjIAcqONeXO
JX7kY4e0WuZYYRBD77QmfJccZ3U0ofNxubAKZWgBcyUrNlGPTxxvQbRiP+Ao9r+z
ipxE+0f9+R8ZpNbeiHKrAw==
`protect END_PROTECTED
