`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SXpjxLUwSTX1tAJ4yqwuGiKLbP3fsTn/xemLXyoZYI1IISsded9q29rrOZlOyktx
8g7TGH90+h4NrdyJ4fpawg5ffBzqKI5scCpQq0dZRCZD9P5RW/yxGazE6FJPsbkj
VVHrbMKtB3EczppvMBIASOO+8+R9m5c6wciUIftHRGiOIFcCCZhjbxkDAjBFiK7Z
/rcnj58ZPp17m2xBy3CoiFBMqdn1F/LZHFNB+ZXGkEB8PX4wbCDhbn9gCQVumSmp
mNBYnE86zLCGhb74HTiQKxBq8pZjCQ53/hGg/03N1ORMQpmyPTw38GvpYBV42BUN
8HLLujUrD2ZTfEn5CY/0tw==
`protect END_PROTECTED
