`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
//SneMGxqbennL6YDSwvOw7HV863vy4niDqO6z4TNdROyycswh9n5K2f8RndTl+0
orQdf1hYTKp71XE0mcmg+DRc2xpifFVdSNccN/StKPQjLh4nsrmUZhBf1YYAYHx2
Vq7Ny+5/VLxXlYL9NZeUAp3wCX6xGeV1oMfhjLFq+oyQLWSInOfJAepquMFPbebq
aEEGIsT4/aZanaBTPaUvyjOFfoVvWb0vxa1CamydUGILULL4Yq9y5Fi8t5Zn2qZH
MA6Wu75fk09F0Kbc5nTBdbUGaDEG7QcP3nsaGqkA06pvm5RGVx+Ue5vyy+wQV4tr
TAkWbWTHNyuC1rnJx9+t4SDC8Muh1rEfselP+9XbYv9oL+G8mz8k+s2DhhlbhYmW
QHWxktQxGJAj9osJf8qDTnWAMp+HaKTRk8K8W1cMcdCXj+jbD/fl2uypwrxEXd0b
4IlDMM8fU4RkFdlGwRewR2kbC8LIPCOX3NTQsGDNgIY=
`protect END_PROTECTED
