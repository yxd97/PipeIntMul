`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvQZ0rLJ95kpgPUUGS/uhDuOT1R0AMNyikzcC3T38JEtLhZezUKkW/+ftsh2nsmi
IAv2JCUqxdRvM/yKVl1bX0bqmUq0NlK5v3MamlSuraqSHPP1dOuLvxUaM+qs1drn
g2rWXSVcLk74vR+BP6ZexhgA5BMwps2mj0YntjjCxdfwbeT+rd8AzBGL0fso+HMQ
3pzr8MWErRmY6Kb3N1jDbkogN0wJsIwAB7n8t7V0o4uXN031NPhSU7cqYbNiX0UO
NfoNfubRx/oVXECXjXoPJ+wxurWzYHRu5nPtL2R4m76NtUGfSF6P2+NIEmP7CQUP
6PAzE/Aa5FqJy9904tYsJFVcFSPsllcy7NEjVvUrJsUK4t4qMRfDSrOzLBfNcYT5
w8qpP01qV8MtDeS4BQlQONgpbDCgjHAPD8C7RwpEgn5Gtt3+byIiC5ibWmmaW8vJ
DzcWt9k7lHjziB5ylWEZRl/md0NYw9PRI7sDW+uucXPHah+Za3Iu6Y5pMiEZSz+X
t131ZO50SM3I9SBjIMuaCQjhK7sYb2NFNey+0TdPi5adgr31aardZULDQd0F+rSN
RPYX8tR4AarR9Qgu7HGKiX802umvtHlNm/pgs4fKIFh8aGRwxAW74pm0dmr7DF3O
vxNKFosXG+myNMwEGtKr7VLAmnL4s8QWsUKk+KaWi97yl8BbwzexGzvfU9T4FYTq
poSQ9hTyzcxlUEUPqjQjEXvi6XmQURROZfiqGQnnCbFGbhozlDk4pT4VGhH4/bhH
RyrqFax0RGuknjrJlG9bv/JUAMb8yDbDEGiHSDYKOu/Do7ZvQHQKBbAGZtfERCnT
ts6TMDXrWoZbEAq1X/j4gFJuedKA1UCBlQmxuDLPO39PjmwNAUDVcibm3He8nKXv
FSi6p4zZLrEa7q6pbBZ/Gi9viQ0lBPg+NnTjihB8Kf8DnCR1ed8h29ng32FhLPnz
me+1lFrsrdAzW080TqU+sIq/iJ40k5IOACYThnbXcfOQkWbqOZzwLUIywnCMJ0K7
R7G+mPeGkMaOTFJE2sWUmxFNn14w+pGl6byO1yo3C+9Oz4hzXbZ8s2JL5qVCBXoW
DpI04olIhRlORmPLf85zI1ooJe7kJgeNACCZcAaDO1rpek0q6AfnTAuMw0ahAbEp
FBjUr7xxlKsvskm1AhnsbVNK1CzBrmRPSXqY4xwu6VL2uccf1icMH1Vo4jpvgXsu
EJNcYhIMrGV1K1SnupfnwVZKmJvazeTSKVqbjtA7M9UZrCBrtG+EyuYwnsvmp4DT
iZ4f2sgn1hhAApBZsUuvLKMnlDAMtnuTTjw3ptyDnZzJ4FuRc/zLnpmNF8VNeUQn
c/eU3WM7CkjURV+uArB0JAbcRNujZt/iajN315I8vHWNORsR+MYROemX6HwT4OzK
AKG5JGA6JGhbKSI2ijqqipeaX/gWDhB7q02uQaHH4C0yGxXXLpKpxAo8bdIjypfN
C8TkOptjUSmZ5ldRl+7LeCce8I5D/nr/Fv4lc1eEf3H0TK1hAqY6M3zI9JOuzCh9
y8Gz73/2btHrNRq4UZacsNiU71QmaBTQy76xrdydgRvlaTPRqmqexvNVhi1T+Zf/
95l4kmW/IPJ16Ht77MY+fip91mu4NjAYX1uUPPxDNVjbk1K2RFyXIxDVdTr32zSD
iWlz1oGjvjsHwpoWZMvvVDoBYma9euvtn1f23Q4YLceBGzQiCiA9OTb3tDj1T1VK
wEzFP9pZRMj4knPzhpUIucwdGgqAPHLqK0dBEqd2i57NsamitaR4pliHCYP4e5F8
32IY18wfyDTjZSGinVinL6nMcAthkr30FC5g+hDBw3X0ZJFAZ2ycvosqG4+Bh0f8
Q2jljJmtBMFwWNLp723N2STef24sQRmelV86MNyh28/3DZwML+iiRl4WLV0mrv6F
VVf61sYWaGkLbzBAHVeAYWfN5oCmcIyRbBbJ96VRHhTfTB9RgpzdrBF+jGsnIx9H
AvJdZPWGr2OP0QiKs0fG/gk2SS7j8yL0AOn7qhFPcN9J8tam2xAeDXuRkC4s5TvV
ltAiVGYP8Th3Euolwh8Niyv7fN9TvF5H91WE1oe97VLJogGe8hrnyId/ubf9i9lA
MzyVedw4Pq1Ejo2bQ7i8zgPVzqWxKsgknyjFZfLU7C5H7nXL/oVP5Jwnm8Rvi/c+
86FVLZwFiv1ZyShymFRkYrarhIbBMehBXCMACz7AaEnqM2FWnOGVhDMer47XAZXE
jBskvoBs2M6o4vYtuhj6vP4O54yo+3O+VKo0LvPXjmK2prwIL4zalaqJ12ta7hRR
/zrmG78Q5J2XjW8lTkoG0rMEjHMCGmf4Zo2//PRpQ6+sAU339vPtBDw/Xwzwv+m/
9OL60hMKz9tR4gWjqhb2J4jfWVgvKevajDlhqG9lF7OpM51oQf9A6z28Y5wtf5AD
3IWcfahGHtz84P8rtdfVn/De18K0Cd84vJ0yt08Iw8Tn2PRBRhnGgl61aCNotiYZ
GYorAkRGQRaVBlrgH67TdBmT18ggDmF4ExBlO0GW9Mc1FewvTnKMwHGDnfjGVuzH
dfyimBgT5d2zIoUQsDVRbyvuqAoLmPY8CeTOjZO+dGcdbITF5WpovMAXwe1NbIhh
uUmsZFBDRYNMnr5bkUIbaF5eFf3bNn6YK7fH4EEPzBYoMF/MGUfADIgm4aHVfOto
bwMIJK5WNiRL96NvwLfKcSH5R0WBimzAjYaIzW9Vg1UTkXY9WU/R77Rv/FWN2Ngx
WDcYl0TgzciKjCZYpEhqjiwIBuo54tNlJJTbTbSAX3/hYi37o/mBpS5/bs/Dla+B
eXP8S3jdGOqvsKKID4THWor57qHvX1t/8rbK69z4JG//5Ed4+8pGx683Q2L+lbdi
IumY/odk2JztobLMueGt9Zmgl1cXSUNEVbB/60KK5EA93N0XyEaWTzIqnUdBJuJ3
+yeXfGcrSJ21vHcxoeXJsE5kkbdRC5b53xwdjQsALqhE7fTrj5DUVByJ1DPLKNQZ
a5tsyw3xiCQJvDrh3M2NRQ44uRypfbYSF+kyM1UMjZaCGdDaNEl/pSHtPOfFwHFa
mOEaSoRgoRoc3xsNNqMTAZSVSpa9rjkWbLgddMrjWkNyfnnVJ80KTPFHKO/BFX8T
463qLPLTUX8YCrsQQnu5bjYxxYgn2h3XcLm7sSv0CQ5138n/g77+dEPcsIC+X/vA
lvjPKX9EA6DDFl0GAf0pRDwL3jSFfw+VRFv+Ipg0dQo1f/JgtQUbdwTWXglNlAVX
ed9lbnFZI1woDgJBBjNyZvLOEKwnsIkqjuPepLs7FLI1GioFEX0RFQsxgQtC59jV
pdc5PzdnVVW44F1KnptHngfO64cSoe01JXIaOFr+taBRmkJ6jDypoHcaEgvpc3sY
2HbOLCly7v70gDeVy5/MWj0a7aMYOyzgEE7w5f+ixcBVe0bmPGDivM6ggnFf9g3k
SDXhI1mSmT/ezEftjwcnlp4A6HlLZaDglLtyEk60BPjZiFgY/xNYv1q4KkUytjv9
ySlzDdQ4KXu6isUIv0ZRac/lDRDWiaewBxGy7golc1mav2c6sFkxmxTYTR6fAgGG
n9HoNpxKaoJxkRzGYGbVUaCtVTQWFzkLwgCnbDOa5wyHdhZ7SP2YJR9w29NhNMAV
DbxX8e72vmx3GW8q4c1nvLGp9XmAajO7AGDUwJLNDNUEHrmcyg0B67OIpQZEq54Z
29HMyknzdjXY8DEK2bcn/vPjN6TgEvtSGpQhD5ZOLRUw9+MrwPLi2QKAKZsNHjOF
8S7hoOqZkA2KcQNI+ymIdaPfFLWHHkmR4QVXcsuZd5jfLMVddqh8ZVk8iuzdoJYY
4pF8C/C3nWWeni84agbg9CnUHoY1QhOHXdKy4Js1062yi04tNZgXVFrs7++/tYwY
EchcTGB+r490ofRFcvqKIw0ICIaestbrW4jc5UuR1Rm6AprOsCTdHVNDVfJJGH2n
SVyDo1j2zFHQOX5cfHa077iP8M3kAQrEdhSPtYaAB32w8VCbrJHxjvbMRIRtxBFQ
xmdnB2fkkf2dHrlyE/HW+M8aptBs5pa2AoirkPC+Ic3a4Gxb72DuRWkZLBpnMC9L
0WjewBN/7sphSU6Mk86SfSUjCoupnQ/cGokXrWoJeZlzppi9v9Gdd4B+p8FA0kEf
TWMjd2S/0bEu+h+dEvWGhFyQoT+UGk6/wDlwje/xP1FyOQSGag0+kNIrWpBd/6v+
HyKH2IMEAZUe90WPM4jHzzgm6E6+Xfj2ySSqhAp6tUmJCLbz06enQSyCfSEEBOVE
8ScCoAFa+EXkx6J7ckGnuPxi1oL3YxZk+sEHS5dnxyzHhJbQTIo74g2Zl54YJnYz
eI5lExeDbhbzrHtrkI4Vg6NsaMVgV+f21sqOCKFGul027OoJzx44kal+Z4OGh8TY
zNnEXtCgVpCObigIBqmE69mx+7/UJCy4omtsEIvPuU/U5fZodjcO8yBnVRuXgrSa
HfDf6Xs60LCOavFh1HYMCufNTmSNHBAeWl8tyl45BuC9kA+LLqrA5Hg57jUYKKdU
pKIjlzMsTxqtv6SSNgDxr5OkkAErcC3S8GpmNNRK2IYZCB21V8IgntiGaicpjXw7
XO8sdCfbZz2kWwK4bVY9b3BpHX22J1NL1L/BnZE8KRvRmf/BKatfa/7OVn7xCZsy
91EsmvvoRcx4CkiilXm/MbUj5jN5pXFZ+cDsvK5C+CEwV0gyJBikcuiiIXQgbICW
EqEvO42/X3ZbNSrcid1aVMzT9tIhfdPN/Urf0czTueOFqtVdiK9M1YNdCBbvaRQs
0+Vqo+DWAf3lQiSSYsDlt0CCGG1EQHpDFhh9Q30aMeo8tieLeHOYt+Na+wmbDppg
0Gst3Vl4emDV14arHeO5ypJ1iPiTfZaHUd4exhBsXlQOnoWqQnHHSI7oWfFn4qbK
vuLrtSCZ7yzzvQfjv955z+0teFiPPh52VER0WuMJLWhX7lD0G9LGqKFxFqvtn5wL
uswIj5CfieMY2RjGqYYKTsP1fO121Gt8cOaLRh3ccfTdVut06D7tyOoxinh3J2QM
zUR40vE7eDhrLuVvMCV7jYKOMAHFQVelV4wNUMRwAqdE6epcpM/tgJ7LOGId23Yi
LFyQbgS5y7yNRf1K+nMg+LJQtBzGusBj9FFFDwLhw/N8B80quGVE8DBSG2H5MXsQ
pFWzNlbj09NMMlLySBb2yTtpv4gpiCeqSDiJYSOfRLYyoKaK5CrbsnkdcunjXw07
3fIl0cTmR02cKkVorhb24svT1loTKXp6ZHjZHCfIwTy6QUz/x4AS/h/cCCguolJ9
DGGbsRWJGQPNg0XtYCFWOOzb3SN4BiQqIFlXV23ar+/vOiRnHbayaaOdWYagdeDC
WRzbupP4NDh2vo5hvhNF5lUbTkpdGlD8DXZkcwubpkFN/ul5ZxHqQN+YW6wwqXlZ
1aZFsq5qrilEHErtYjv2LGSSvtf55Vl/7xMhF4fSNfi7E86UQFwWfauIHc8QOOFU
asCu2HePjoWG0xhZ3F5p5Ru4fhxCK8xSmniFKX7zwQ+IGYcBZ/E8pAbN1MTBaw9e
aMAoqIzwoalwgi+8GREA+WHH+v0XbtgvCTVgaxtLhgVPwFCdo/400ZImI5Ybxvlx
UPtp+L192esAaEOvOlbI/S/m/ZjLYSlwdwk8BusxpCjWQp/uHfgv3LZb1CPX8vCm
Vps1FCNG//sdJDjpHLEnkwhI7bbp8T/NElrybJgX5cxXfutUOZzLPcYpclV5PRGm
tB7ZH/TLP7/IGm9NS3Wh4d0i5kNMqf/95mPr32m5Zplau/ObtBm9beBa/80L+4QW
NoEqXnxB5sGsS5OYx0QZPOev5K+19SkqBqr56M7WLN35l84C16W+smqNkNYExhzP
BAVoMmXKk1dXhhczxT7nhBeOKOKlpgDbyljsGwhSMO4524PUlhmvxj+dEzr0jwoJ
JFYzQrg+akfIOWqdwKbTAPwmlVT9lnGyLMtB1VSt6ypUqcmrW4mtSFA6bjvkO4m8
yZpH3tbxSNpi5MVM28CH/iTYOsGEDWBzpjPbc0P1AEzk9eX5+fWr4rj2UtALrmPp
BCxveY+HJUu1SfZ30uAf5FoBL93iUdqJJ5bOvfrnDk4jRVt3QB+c/CATEEp9PWZl
nHNQQc7wOfUo5Shwzr/8LaHKu3EBuMtmlnhd93Y3iCIZHLZyGHFJvvvo8f5DV5xq
5vXHsIDac8kehEzhbu+WU2BPAesIL6cfr6opBNF9d8IuYSu7R01L+tS/yAcz8gdm
/9r/BO2ucCXhinJN7J31ZcODh8AZJVKf8Bkht13p8JZyRcm2Ni1SNA19T0g5oSRy
aysvBUjCDMPGV6IWKWdwt5LIldduxr1K4XaV92U2xBBV3tNhIpOZ7xVjb62qODbG
ze+RvOm4u6HkVY0blz6s4wHLTHWaETZb8CseiCHCDspZMBQaiWXXYh+eSMgN5XUk
eFZb7ur3Gl3609DYeCFo4VuWnbVA2KW2MnkLvxE6A+pVRKIc/CqPhTi4heSXeE9U
GcxQf9HIGt/zRWaqqRG5k/6kNb9hwEzfIUIgQ+YIe6HmC9mTSmvrNFLoy0jtFrlC
qslAKQDXul4HYe8vVHonNrn5BveCLQW1QkbvB+Azglio50x+f6iCGIBZqi14mS4U
Jnt4CzqwReM3qWX9b4lTMvDiiX1yF1jHQbC633MqPlaf41j2kyhfaoI5zWoAOJcN
rykP6djf7U2aA9TenUDq0LJBzM4yrSGj5LM6H46oICLRi9WJHc+IRC0+1CkYChBE
5QWaEYt07mfrqFXO/iIL5htkKkyvowVIWEeejQm6qaLO4Wx14lwWf0MDgTJooNBE
XVROSUEZcLn+2Z8T10lDtGOt5ggXapfd2JRisG5o0NW4Wi9XBapZIU3JVM/cqUEP
++hteZQqSNDF1tNWSV1oJY05a26U7Zffi+MWYchdgaWQhsLEJR6s0bYeM2JZLlcK
y78Z//EnEHCONuO3Rj7bMWZaG12ERK1Sv3LpEKR/qzBT1CutjPm3r8NEfbtPmBZ8
PiYR/VfDg7ckZ2hurYlZxSfPZHdm4Ap8ah1Rvfwpj4XRsDjXkp7yupFrFtIS4u/0
W9jbwzPjl2mbe3WBWEr39Jv0LJNycmmdqrHMhIZBUgpboyV0ymI4y1H76EC8SNdX
8H/rSWNktUE/aMe9gqjUQg==
`protect END_PROTECTED
