`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bbPns47Mu6yn/2AVCSzMi7HIN+UNERqzfwpk3wNyhYqXuN/o2HxLExdAT+oeZvCx
OhoAlbig56uBAnaLRACtNsRgOGsLOYNdXQZV1Ebd0a1HizKNz8VD0CfUmZ+OPyvQ
0yrh8mwhiRIZefFYEOsFt7ZFqMKQLqEuA3FiOhpFB7DkTRRVnR15subpTLA3eXir
Opa++9c/d+sWo7vqgW+TP6A7XPn5Nb3CczPXXEJ+hmiVOxhihck3hWwh2R0E+HwB
55cdN7N0EtlGAwo3jydJ9Hwqm6bb0iAnVmOtRSuwXpDBi+yBMk6eTl8+UN/UkZX9
I/0JjMGc+4daAC7XCamK/DEvfzh+6UMuvxSpvJWjFlJbxr66/Tmsyr7q548xShA6
VNe0AVkWnZLOUDR2nwAbNW7uKg7FYt2mWNhWGZz25++MdJwWOTwxXMrENQVHSCnF
sBJGaXbTbYkkpBbvzjtrVxhynJ6S5LivXvcEHsOXBDhz2AnHJtvIUs8BBepzjwiv
`protect END_PROTECTED
