`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qI41XAB8hlriM20wr9PZzJYv5D7x/eBWQjN7ARHzVEUW0TPcipP9h4L19rVM7Lzt
0/2FxDpIw+zZOQ5qe6+2XlZDt51qusqFYSI8tfhQXyK1X76ASSke5s3OQJGmYe63
Upr1pb2Suf+wrs2nAPb5BnSRkMQKLQf+OLHeG7PO37yS86e1mFxUWer1S5V9jwFC
kLsSD+CtCV+yjKVwIk6OMoiAYf4UFOoC0tuabooJcfENr1d0q6SIvjF2rsHErw0H
i7PbCZ+zPGWbTYI/6O6vpLHf4VYNewqwAJMhib9UDJeYXynLIy/uVtCij7WW+Ec7
gPPCLjV5M07hKvJnYeXJzlEyAU3B4yjHtYDNNNFG7A+T88emdIfJoSNn402XPpd7
xJ/G2iNFOWR3/BCvNnWm0jAAwrSbsXryGLy2opCZwopWIcv5It+QFxkGywXLjq4H
s863YilA42SftCRCK2tL7EN1reJlXGZYFTE4BoGxx3lC1Faip0hv7bM065KE/XbO
`protect END_PROTECTED
