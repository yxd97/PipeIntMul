`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQJUL0A0upas/kkLl2z97nvjxMWewMyYG+Dxxb5fWHZWMXK1X+a81GZZrRf4KF19
CrNz2iM4ysXqmNeF2LDXXufEtWGZHoN2N8bn3N6nHvEXYNGH1KG4Gttv3uUn0Xu0
YuPqvbtG6DXoBcrS02PSwMhBSzw1LJR6LbUOMCaDTSIdhjMGMhg1ynVj6OFt7GnE
wT6rez5xx+H04bSCZvwa6DBOUS6/rrIuW3/SJ6LrKQKmS6fjQiK9rE7QeeSv0gb3
W7tsQjVKLo1gdIUtpjAnIzeC8YxaIjmsAmRYWSWaqYhCCHdqiSw/p6cvte0obvSR
LZA60WiL9h1WGOJ2IA9hoggcpqcUOJ7df8Sykss+iWalAE53SrvUGrt5m6R0K5Gl
bl9stHfbCA69sQZ5M0xoytZRziciV4IgEG9aB1TnK2Sv+dwGr+BSdMY1ssvzumPO
qSwtcDky2kMJHTHCmj/kcq6AAR9wo9JkVqx0bEwLsCvCaQ41rtEzqIP8vJtEE12G
OWjOpNN05KXPn7EIN8Ce2zg/EWbQRmOss55Q2i5dCmT8haRhC1UgH/A7wuOrqf+G
jLgbicx8D4hvbkrQBxYHYQJRU2VGZDwkz++QvFfmtXpKAMx2tTxyiX1yQIeekAUW
3XBEnQNcS2W1sjpQGlquDWGovZVgqcZql2FuuVo0piBHV08c6EdX3kMvW6BMJaCX
H4fuhguVhTi43Zx6qD0+9qwdbebucOqd5J14u5NE2diyJVDIVRkoWrgV9INCMlj5
E8pe7oEGwGCTiuwra62LbSnAnIkPKTaol5W/+aZSlc4zFV+y4psfTorpb6M5mbRr
/6XGYLE8127j6Zq2CNKSSeIhQfQ4imR2wURFaKs4DoZcTEDLqROlg0S1EQtWsdHb
PYFb+6vfc75Jbl7BFj03Pl3QATs0d84I6EphKR1i8Hz4Ek2b3GzvER4MJ4plqN+q
6ywIlidXzBbI5LCb7pT+HnUcRVHFrF7ZcAEanOsEh5qzguIfG2Um8Xqo3h4VkG7F
5I1E+ifpK3RVRQtC3RAe9PVWCmk0va7qCZ7n62CqK99SB/8LnOyTOopipCbr92rt
a6l94Vz97pMjuWXBoqq59AtT0xaIX454C4A/i5wghziBE9c2yItcY1zUb6FHhcbK
Xab2Uu2+rmUpUS5rwt2GIY3DGSibKxoKUZ6kiwYi/YSQ4Zwk1JQ38eEIFkbRVYsS
kLbYeB1HKSlgYF7XMB5Ul7XHSrKKSaMxYX7nthpwb+lYBYkjuL4urmO9BAL0lhUO
KU6FM1Q6qdzNAU9Iv1gRpJ1DfZmsofR+NhO0iZUmNfoX1Fj3mRus36PWx4F3qHdb
huEkTMV8edxDGmuKkVAei7k+VMaveX7WA+4eFv1H+KeD0ttGWC16ZtyN/kRudae1
oei4Aak2jhhGSo073jl0hxCjdcM5hFSNAbsGaqZO7WO2HLD45S72VB5ZCcaUzrbz
1K1mtYfO7oHAqUwHZi/W3ZswGX72uZE9ONWpGCrk9oVCeqblWRecBqY5NDWskImj
orvt3s90fLShKYO2JG8QtSiVKOF24ZDMU7EqeQFQfVtM8483lLZyLQC7Ply+ir4b
PH6o447/+Zrbfy7nYawlNcKsUGfGZ3bh7qEwhQizxjy/v/x2QwhfjmO812JO2vLh
QtpmYg4mMUfOKOu1ofqRrZwX+W2e89mC9V8RhdVAhxDRfI+fZbVq//NmDbMQs5dK
zcmQOFGs/6fSon+NHHIygoILWlfux7QTHevn/xd4CjNQLR10OHhe1ZxTY6RSvdEg
+Yz6Nf6DtcyKg2ptblrm1/d0S1zt54axwCCcz7+nRXk6xf9FpZhxJZPSMKpNHSDx
Z3qvBoBBu/rWXu515euVwf8GEFcM+Dv9sNpNlkwONRBagC0Kgu6ANkXBY+ENor++
+wfAoaROOga59QejRWEfmE/VyqVmVD0P6s/066jKx2VU2atMuQwwXP4ANum51Q2e
YdZFf7E9pXV8BXLTQXIuewh1CS4K/8IOiHcGNu3edRK1K2uQ75gpxawOBfMvBQNo
BCXUEt7hAIOUuGQRkAsk8QgHGSCn3P+nFKcwIELgMPEarSawmQRJkrneuHaY80lS
A6/mofUFhCiQ7Oz2EXx1reECdUpVVSkeu+l1SSV7kSxuQ/xBVyVeVLV11DE+PP5i
t3iYlBBKfoWkSXCn10EA6vHSlqbj1OCZxe27AAKCnFYjl8DeXs/EF9qQQkaDcPIP
MpgCM/vN6AD3ZGx3IlfU0J3DS3aIo4bSa7FUJwN5VyNnrWg45tu4ffLraKtT8JTq
w0OgO9C+m7f5P+FXkaSr+2hEhZEPYRftZ95fUEdp2N68mY+TjXGmaiYJkpG5SeQN
9XuYPZcjkBlensidVvjK5gNt/8f2kD3+ajq7fCpciTgvw0f8QvW5DSjKmrRbtfhW
6nfG6huUGKLAmdBAzbuNC9dFBAgxm10pJk1vaXfHgvyvuJnyGUXWeYMFysbQ45j9
hLchSh3F3Kghazk6yurRkyKnkijrFIlDOgbn+q1pE5+lEREym2B+C81sufsHP56Q
7hji/SFlfBofO/pDqA8nuaGmXhbX8TcRu9SCSRNXhYDJV5A0TeMGtRFcwAFI9AJe
Wt57Z4W3tHefHwpuRdLfwDKEuOndMyl15CpndgjrRy8lZ8ezSD4TBHfo5wHVAPHs
PHLlMFlfK+sfI9AQX1XEhktEvMPXKQtCLMgOjG9HLy+baKEu1zEtOHh2AiVDoniF
PHFTRwnO3Dtys+WNEah/A6A6QrM8JcF4PQpaH+LZb0jkiIuo+44nllolUQF/c1yM
O20R+ducYAQwmXjR+TyD/esGeeQ8AO7kc186AW3marpr4HJVTqgAlSlMnGLl4DsD
uUihSnx/bLrPMdSTIunjFDwTGLC2WPbLZ+6PbX+L0xUuRsIRk+KkW5dQj+b7AFKO
nDo1oxFovX32PkJNe/epyEBiagfQyHbqnDFHfeeaBRHj+2vqJUcVypb2NADKTfuH
RkPNGtwSwK88jSc4btH5fRYr2GQKbbHoXi+4iNJza3i0YYB7OnQuebisbSi57nKt
fJtet1tVOHX8mEB0OGrhY5WqUkmUnswsJcMRGlBQvY1NOIzbwq2UHryXE8tU0Xa3
cT6WBw188hJjf7hFJj3IqF6xVuwwoJbDl3zhcgJlCK91B0Y3uqlr5xtUjEMFwFaL
P+HYeIq468qP6oOkUI0AUxSmYislBSmazj9q3Hmyrzz5THr13bGAbqyGagD5iJk+
9dSh6PbEOv/ooU1G+ZqxGPkbYbx5WLAnTQZQ+4iwqClsrDb+MRIUNkoZPZ+3fouU
Bj2eIlD4dWOiL/N0VBSqwwiW2fkShLgnJw3ItKyJ32S7AOiY7d+u8kXZKMkDHfEi
Vbjwn/OJjOyauaBSmJlsBGWlhygrowZKo+2uO7BBfFitlMKyG0uGc0AroNorqwq/
Q7xfTQkgSlOiYkSR2x8U/YJv0ZNOPZaRTFexaAGfJPFCI30baxY75HLROr20pUhr
JHAlV/c1PxukayGssOaHKwIpFnIocUzEWF9rIAEglVaZ2so8mf195GOga/AmEQSB
tN7Tzx6ORngsyD7QXMNFfHgwxuF8lxW+rBRku31sVl49h/425v1e17ngcP2wUeaU
9sebOMCY4lsx5uPThKq1UCBSneSnrI6Z2bf/OEdJGgamthC4vBOPvpolSj4d3Kit
D7qsKldkWMM649ZxzNGhl6/XLZoHJlrKGohHCQX+CjFfHHFGU4QvqY0ERq86VYtl
Hr3sXs0tOg2wA8IDJIMiLY9HaJKDXRMmv5nxh8yXsaBWPqVgtYlbdL1mRLJfI3RI
xfAqjvC0cWHaxLKyQzTfnx8oi//1d7L4Zl4Td76ABAijl/POLpQH2jfdTlrVp92X
7xVJyJ8jfAClk63vt4Qg7iBhtba7AqoxFfteyAoiKj4FOtYTBuBX4YLHy1aZcSpM
6snzta53Am/eikrBYx8OdeoEcr244bhLhE8J7oTvHCLhttDlMvFTRVcydg3XO97h
PAwdg97AhFJv4F4nDbpT8rifOMCklKu7Us1iwpm+0pwGKxQrIBV4nyJ41pO0UyEe
dPt1jhvQaW6Kjskjk9Z2uqGHIr8MZj/KIrw/2o6xvYOSoLTPBer9B6P1M/cXVWPt
nfaanLMlqBuh6B5q7HnOl4BGfG3JdV4eDqPdi6ZRDZsO2bkadBKaKeNFOUDEWGLR
ti9oRBlfQ8fJrLk1zv/Wtu2WT05mWZs0aKODFDshxSa54NldrI0JVdf9/JohXtvJ
iwRo0Nk40Skz9thLtn3oh03QZSFfh9k7YcgMl/KB3JWSxPhMmyAQslKcneTltMc0
yeA1Ftp3pcQHY8cZfA+DG+W6NSg7omUxFEzMuP9OOYfgaJl8pHPnNpC+ri5iOkV5
uJz1Z03eiXDqsXokjQZuTAnEESz/cGs0ApLd6eZ+a8JMaFqxcH0gcVB1mjPA1sm7
/OUgcMi5PZ2uhNgfoRSK6doMdWmS+GR/239s6F+rekXMS3ubhaab3LsmoeT1aI8V
ZQJnEFu7eqcecnTMK353wSVHlLvV6CjwR/7itCvmSoP0qQpA+uDSYa/E8EZY0lZe
Zx42VsvYB97sfegPv5SmKXK4qG1baHZEZpHl4R2lH+6bL/ieavXVsk96dGTZqKBE
plhVnwoxOPd5wj0HvGZUf0hsTa75DFevgCZYFobGrgTqQvUzQxZoTpooAbvJFT8U
+3o5N2YYfMctMddPr73fZY5ofw+gK23XteL1qrDZ4jCoBSuRToMoiYXO4XIlogL+
hn0gyL9KHGL9TW44JlOuMjJryWxVafjec7VfJunS6nweAGY+aDHT/qG/pvIrF31T
JWQ6OaZKkHfs4gru/z2OHqosFQql2UsWOeEPYiKPfChry+VYEmU0afKz+fP1aOoS
r02DB5OYWA/TaZ6OEns+088BZaKeNz9zG6RJV243MitommCzjQJqhKCdm9fDO4uZ
YV+MMfcJtAhwLChfPNmp/rRjPOKjvcUjmP2rpf9Q+PsG9jAv3E8xCxUNlXzA7n+k
I0uIvxHfMvzUglOWLNHMrrme48T2QnEsVc/NvM25bC2kyNHuVLOxK/NKnk24AlSJ
ZPAyiFxzcyMLm9QeTRRTxTjfEcVIHk2rYgAd6Ge43H5+MViv8h2zB+8ZyYF81nYG
JEODSUP90JyS1XpKsluJbIm2wjBUdh59iBIFIhNrfjpAoBnc8w6J2DNrqybnn+Dm
Z+1Ifh0qNwdhCsjy4WVwI1fUbV2P6Gq4QnhndhQZngz+PDXmRFpIo84VJet4OpOt
th+SbSXhboGZNfcs0rkazdP1ilm2qmgwdqLe5X0BFHJV3AQ1/wjW8flrko2LiVuw
2deu6MG6tEjTusQ7Vk353rJJiAWLLBztNbyC9F5yOjMY+F3KNYvxQWOjZtUaPVID
cn7GnRChbfyec8pqbKUGrLSpyvq1ZzVT3CA6qwce0tYs1u6CBthqO8GJAT92RFdg
pah1LdukavHyZQ7MY0/ZMsQjjHU5nrJxRuqxo4b+l01OFt+C9K8xHuH8QrGtihyr
+fX0lP7eBmIVSrtUsylyRuyJ038x/EwvOg6fSCv94PyVsr7Fj5L2enNQBqjRC0il
3S/cKy0j8DdzgJb9xveT0hlYIj/PFdkMRH/T6ZpSU4X+Qrf4/Xwgz3SZ2zaFwcJF
z6sC/RFJ9mM5E4oaXru+5evjNhnfCWbLRBaagLIooovYRzXvoYr+ufH0gxn69j4I
EEiKDsbzutaYsS06NWC0TmG96+kUyIOHZBSyZjb04h5iwG4sr9JgWTjP+OL9y9yT
hrh7LjNpgGfp4qD50sTI5yXQIqzhEuVhTalF9WOk/e7A8C/ZBZiFekyGlVPEJyM5
G6onGBPdN7gHi8nQyOakPuybyDbVHMk2m6XH1NYPSE4qyXXLAPVPG0cgkqJ1lJrQ
a5Gwgc1FbT2WZMDBhjy0neCLbanzpYem/vNPiLjVr1p7aDvBmDtTkJpFRRnhDrFe
XReEgL6Pz8WGYoiCBqSYdJv2S9MoHCDzXClFGm2tUfbM6CTw/9HPIEnKFfMzFzQM
qCo0NOA7BKNfpfveReFH2vKOksyq9XJJpNT1VJ8o33OwaS/AKckyLyL88E4d2bDY
wCMwq+/GaEUQXr6UIaJaOh4RG0qxcyqj3NmQ+6Cb+6LiBss+ps7JbaeJ8lsFUxMm
QjKzGRkvY+/lqQDtJi/RdiapWH26kDOhHo7Flj411sMcQVmjYTffgU6OF5XW7n+J
JO5pYzjohmVsxIuRN5AQRDUQI8G82N0/nhRkcmzSvqrMBQGNHuzUjDejvtO5PsZA
/M1QGFYSmYlFqzZJGA5N0ByN+kxxCHy/aalptAhUqx/6Jy8ooJxI0kTxvCZuMWhA
gTSaszIgCTkzcc8aXVrU2OWEU1l5ehg67MI0JjTbzIczuiWrblSoqltvBfiLoV8/
HVUCD6MD/vWZ9koo8LMMYOreSoulUeqLFQvnA/BFDk+WENi4B9ZyAO5s+x+X0yt6
a6O+SnSgc9tOxQ+1mxDTgWwTbZ9uWP0udJ51ZDstGYcBVJbuLuFF5fR8GJlON13X
6t0bjzWtTvzEH+SVDfEHlUctn5SPecr15Mvb29QFBBb7xngkXDVnv9x+igW7gt8P
rbpA93rA5w2bY/E4cT6aT9zqGyqsbaK3A9calBYOjvLwI+y6SH2L/kMKLcZJCAHf
QyVwy3+YIzZi9CeBDBJJg+VhnQQTtPzAOJxKVGkbq+BRVjzdYMDyYR+AP5Q7RSZd
ibzgXptxBrOQCDvMaqo2YvdY3/2ZbNLHoCd9QyaDR1pfLxmt+86wO8OhjygwLoJo
XCp9dmNNdm84v481cw3W9mqAjBZviH9qnLtO0gM6fs5oHeyzFhiNikMnr94e3Hck
ODSqyBkm6vSmzRgXDQAh4DIOBF8G4KqYkR5urPTSH5Gb6GUc4ApP3ndS8N7bRz3H
bsHr/Dp09YVrOpU+0s9FVlByF7ieWPZ5zqetEB+iVOg8UtEvsjndhvx03ciDRJKq
XxY4Ri5hjUdov5KGeyCA9+E2RgUKxjR3qMuqKSOIoRFFNsmf9BwzzcyzgLYdafA1
yMJlXY4vqckkirbvGOMQK5D+gFlFCrSWIHnBQa8lCg5EtpKQpFtQ2tPTEP/So3h0
hwYffC/SZAwVkw+2Qk61uQDDWuc8neEmP8EgW4qudq/eXV5e9zuabSThVj2gx4ie
A67FtMigKq1ms+YBsSWPeU1EEau5FpOZsH1Viye2fptroZ+X5uNwdrzmSNZ+t8Ql
bwQaDparZoIsrb538N+gYeKxRD7N5fwDacUFz/ezr6lVy0M/mVRhF1CYuYlEO1vh
CMncFF1DqEb+gg/Y51WAOIA+EgC3Ew73eL0HbKkzuqeY8bJKzMWzA/XlzC1gW8mQ
YTMNqvmv2x2rgF3HR43bKxyYV4fyLVIUAqgXG5ba2QcZzz0m+1p+wj7aeIrhssPx
7l8Z42j7np7tGGtFkrE4ee9A8NHTOLB6BwB0uFsUerNlJq2LQwX5GwLuY7Cua5wX
wunVkoasqtVJwHfypLYWsV6FK82nWTbT41WglPaugz06MrVIySKM3TQAwxYLq9OQ
yJcRlMtpl/PcatPqv9j33/hZ9m+Jk3QXigO/fj2lkVDos2F712QE3YCC1SlePy/Q
cP/cyWBXbzQVC+XRGYDAKmi3/ZmA8zPne58/zy/ixSmPtn0he9VHSUehvIKy7QMN
c5wW/8nDCBjyxMA74BCJci8kHLaOZ/0dkZyFFlTGZX0pO3O74+7txy2bQuCHDXa1
cBvieCkPMFKHL/4vNGX2e+rQEmhxA91o8DWvwQdYJgT7hhlt2pF9soeTeGIbUrpg
KGsS1D7EzW55jY02d/kQ4gJW6lKDqW1+KSfiMXU45Gd3RN1lGMNK2LRdg+AXhgoz
B+qJLDLwt6uBy/4Od5BN1AUizhU5PMEVVN6+3A+w4FIrXiynFVhiXPP4Rk+ycEnX
k/Bkuub7ncRM8hl7Oq7LjNiJKjkige4qGbuWY9uR28U8gVL4JXmaqOQ0bx7GoZzj
xMNQ6V5+W9BDqJCAmDqAm/J+U+RvRwmxiWFR0K5bTpOWKv8OhrQAkWlDI595x/DR
+5WVK9AfjveLlsCgbv/yB22weAx+TfjYYprK3B4ieLJysblhjRVXrWzHbOPmjmcW
u22jC20e+cFZiyKHb46lCzNoUTcpRYwSVkHNWpWHuFmlJRSiBJEQ/7gnPLrqFpQw
725AKRre6P00ZEPvrbLU/9AJawK3rijt0D300QPErZ6DCIUStj0HB43xxaBhyYv8
2XETtdp6t8he18zqFbN3vUukpzQ/dfcmENloPsMKVEfRCWs+BpX2j8j/4rQ2qe4s
wItUVkFlxO4Pbfy8EF+QBAwouFp+LLFfoByzr+LGaO4up2fbRXKwiRl+xTJRIrZI
Dm3mJgbwJmAPuyKux/LTANjL5Ph9dK34K6t5KKwhl3YgOD5k6VNmL5e1/MCx1vzm
C2dnIl9xPchVtFPTExcM8Crm3sGTNBaA3wvql8H6iQJOxlfal5UeiqWeUAOpQwey
x/LsjwKl7BODogtRuFUHMIO1a+/nFX7TNtmOGzbWDow+vzzSUl4K5gXS4590Nmdc
EY8DzpfZ+DdXgCiNFCBOyCvLIPSQNrboRQTUIHYvhE/CSryrerABtO3Tk5XO8P3F
Et+UM2F3b9/6k511GZdUQO7A/ojo822iYN9EWHFSd2rp5LtswcAJWoNTutAgdtxL
6y1Cwed14dfOGK89X5oIY98LwVZ4byUw/GLUG0aFBRM3QpPuRw+ZhfYYy6hqEDx6
ejH9xxAMK+F9s2hfR17Jgefy3/epm7jIRMxLlVSibWF+/MK+XUYmjwWEed59GS2d
NaBmkCS+vk8pyZER93r5B0tZY9tBLIWHVN3yjwH4wCPNd90dlT+tnzbTUKspp0bv
L2a1iLE9GqJ01usBkQkfCPgTduQzyZ0OGeWXxi7UxazEWmUAHL5j1BFMKR8/gApi
uP21fSpNapY9dMNeSM5GcMcp8Uihm7qwQ+C5ultJwVkMJmVLq+I+UB3CsTBotA2o
UBzQbZR4OFTBUerpKDyKu5BKxqXdTEEhRLJPTjVGtSxIMxrye7/eNYwXhCscAcNG
Kr8BYMABumrvtkhbeAGsuodhHL+bU8RBfjZoJftSmA2Ln2TP3Ct0ZTOwtdS3TAX1
U3LUVeX5ckDfuG+qVEycuoZfwEZ/USKnUZUyMiXRZt5GXKWdvbOQZVHz2bDDNB20
UUtrK2u24VuDccwi7KroYELXgusNAjrZ6lAI5DzY24N/H3lcyzM2MrUJt3vu4kkf
xlPsfDhBSBpnbqTuKzMqaxrQrVCspXGmCtJM4EBJWGqDSQYQWkztlI1U7orsyuu5
tMdNfKi6s58+Q/hy7Gy01+1c3exgPoHC6hOg2kB6ZtyDW4btkRwqe4g6jPcQFdIw
0kuQ8FpPfzA+CWMTcIvrXbAT3AmKSeHKZw0WVg3G+i6Yt+daLjtIAiBoKp6tPJyr
4RrBX5e8oiwRJOX5+3X9gVf9LxPxBd30wEJtCM6exX2m/WLm9BKJmEIYpsMgWeS3
+cU49NWqFhwWUCMQUjwHb232a9Lu0ueU4m1CTLJbLZ3KYvp6MYcbOwK5VHwF8gtS
+LVLjrFd2SqZEumfUr+UAP/9uw6QI8c2TaXNun6gVT8VCv5nknbZTAHRrZJfQqXm
w65xrbY4d6MycNeIGlTUfs0grxtYegDSKzRjfcRYOJXlTnFAmrQHGvfkdWKyx6sB
d2anhrTVdLqMRnkBq4h4p/estA+n81yn8d/pQyMibY24jTLAbPU67dgSL/A3h3MM
+7AOOXSwJcRxrXVQ0YDcTKRgd7a2EuQv99XyP/OD+BzHGvsFZL9NIqf7ysXPzqvp
PD+IslHTNzNQUMw4Rcxvno9gSjqpabDpjLHile/Td3MCXM0LvOh0OsRwME9zFeAQ
YGXMF2148VrtnGheMlEnj5u0vc5HRBUeJb9unGfs9uKsqm6XUk6+CWeQHOFy1GBO
wYqouwnIzE5KHtQtCe5KzLH7T1dZY2QwIx9VUgfz/tbnUsKixqrb9Bpj4PvPESXQ
N5bAF275o/S3DvdOjGkVAKYquhLcJn+c2YT7zHGfTM97YIdHaMr0pcQ6rGPEAjSj
zGQzcnxiwna795hvt1isgMKwEH/7ndphHm8aDpgP28SF18l5qSDyt1SYGnBlwlEx
hWj445tXNIiA3s9HhaYz+LA3M1rDJvgf+70FruFZHXBmREbzv57dDkYGiyUR2VyB
1JzXSMkDA4TwjfqLZZmCFGCcVczphsAvE1ykatCYV+0/yTJgZMuNaa6N9HW4Ue2u
pNCpkqRJTwwf6NlbHbCJMMA0e7oetf2sxCmmldgnCHvb8CM/sMWLHNcAH1Z1ZLod
INgy04veJ2nWw8lQ2elyc/BKLi9ZLr15BxlSZpKfy7RbXC+yVAgjRzusp1vFEFWi
nE8mp/NWLo5p7PQFiIoABDWkG+S8DesmCb9v5xcJWT9SOyzCL1P9d2cPIGY+URK9
wcu4rzC3S/ljw6Oih6kR6NTEXQ4cmTu9FKgvRzgcsjqs7s8qelf7lHwKA42X26PU
jR3sGFkjuFZ2WmJUmCbjeR4sqYXckS3GIapBKsHRv7QfqIN1Vu4wYuOI0cRiF2eR
FNJRymXQ73Wmae98TmeRaPGX/FTi/yrM/0SOGXKMU04pPruo4hIX9PGYG7XE7oYr
vF5l9/c/0owGt4fyEGIvJ+L6uMu4Te02Z1lfpDQ0E2bwJ1XkwIjxgsu7NWqqGXCK
MiS+49IYZ23wQ79oRAGEzeBScJUi/gF0gaxTssaOVocgfwfNzfA5J2ptXcUdNrYa
QVfHlGLeFCA4WQYm8IWEp7F8tJXgZvHU9xGQRb29XKHpx8ef420QLuN72H5+NpAG
QFJOYaQYt9H/jQDyo0QCQrxkKbI2aJhxa4kUy5atJa8YWl6jI0Hrx+8PeWic6xQE
c4uUJyFrMEblil6chRB+SwO2cgFYGDjHnsDPuWLopzJXpfRNgyg/EzONWp0petWV
d4004HmGJHUjb9UMveWi8FJD8SDaPMp4pRA2VejcCOvx3O6tUpfqBsY/06DRv3b7
BW/510dsUnm2Eq1eNRHYefj7QUgeJdF2CD1zV7gRYElTOlE3Zsn8Z5OxYaR6uZkT
EL2+uYlZ8NhnEpYWR/I4YfPYl8z+CgIH0ev66WcamA8p2FV1Hu8rDvNqWYpypCXU
BpuhLQ/aMna7d1n3EvTdSMAJ5whRJriA90YeJTdIdIE9CqdEsVTeb6xzwJMBVd0Y
PQsS7nNmntIjSnuy3OlDSu84LK681UarO3tRe2gGo00akN6zpr+l/KxJ1H+Z86Lz
lXnBq10ihiIArjEtPz2FAhi9rJ4n1zKtGUp4qorC8fnjApjjqOq0dWzDFNAklpcp
24RX7FUkce9CQQPOlnUrVvxZ/JfXIySLyp51GyiZbKyBE1Cdma0igXMeUMxxm++5
BbkhSowj4QJvJoiL+3ihV1ck98X7e4ipd+tUl5M0afKNABrBpmn0wDBfya9CLbyY
+/+o64w2FJQMBqFeMJTL7wkOHbTsH5q8YoYHyx+O3UbwJn1kYxwixq6L5OwTUOFx
MAQGNQuoUp2yI8nnUtGBNuOR8LJRgEvTW1lvV2DdKUDZ1DyYgH2q3RYjYoWmH8+d
t5cR2SFjMdykDwjAsqIzSKj+LXeKqguGsoTcoYlD5eH7DA21aH2iuvSfpYFEM3M1
aca3aftyuk76g3jumrTCXBjbqMC0PJ9it5FOBgKt9/gp5tYmmSxbk8ShIR841Ewc
ldg7yFYhujXPqfET52Q8TB5oHLmyx2KSj20LNZ389omkkIvuBMU17n9Nbdqb4YNZ
NtxXg8lk6Ympdgdjz/dA49vohITP+RrfUUWQG9bPCnoPm9baY9BITOFp/u4srqnq
W8fCv/IzVwAh47uApAwMuoTg5K8M8borBE/A0xZnwIPIm4m+Ge/lCMmaxI86Ifq8
PXw/vdyvMn54c84+2gCAiFNxlH9S0gk04c1Ys3jUdl7Uy6naksSEoAYw8CkWCcz+
rQKXh/MgTHSrz7SxFwIs4lxgpx/N+QVCCniupIUvin6ypNypJCKo9JbpIBD6Re0H
yjr8ar4qJ+BCLLxJ9cjVHG4ocGHBeIh/SueL7U7NBlGf9HPh9j9+pK2zgNYT9pap
yyJd7smCXX8ZTBfzl1K/NbT1enpLGRyP5GpOIJ4U0qqGKVmgCOkTV2fUUJz+3bL9
VSBYdp300nelyT4r4XJcpTPdfzDg0kOZupBRW2ck7306lMZWwbrSa3+RAF1pGw1/
3iIX4KqV1DGguFacAFFsMvVoj8TIJpBp8Cutt1UYDWaOE4SaoL9gzNyu8Y3GD/BN
UdE5+mu9ymE6J61hHsBjZ4uDx1JFqnxqPGLzZf3NmSJWm7Q07OUCyy9zWwdzamRi
OS3E19I5vRh5CrKZ+G0QH3pFv0Nlk1MiWeBAampIi6FnmpEGqLWKbEnWt+hCt2BI
Xai/HR6Z5PImH/tD4oGKH6JctzVZfjXTvHu92JZmIiaG1QY/gg0Z+FqDi1FNlRgn
wGL8k4/pYSlH6J5cdoBXreCL/EVlfNU16SFlimKt+hwQrmHcY+6DUgFNE+HfHLnV
NKwByjQJLdbmpDnCKJJxEF8Rr6JDmXrKEKEhlOAaAXvl8DabEuTRqDfK/khq7pXD
`protect END_PROTECTED
