`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8gZladg7JuZ4DfDlgGdtyzH01KkuZzHvTdapWlEZvXWL5Ofe1+/Ll73eggrOI5la
sEeXsLVE4Pd6H66aH0adpohL8tXokvH/9E91eQqsBvg2+fgZq76L5CtPSr89/auc
bHCo1tUD6xhgu70Jp41CXUVsS20TOFF4T9OxCXp6apWReCLiPBmEnsN3qlT0ERc5
Y+5bTOG4ECdAsCl74TwUH2WKYtYX5Mhm+nBWJOSQ6YKrikXPjQXZeIZE1UJJix7o
hzlvAVSNz5EoOi0fluB74nDpKp/asB1mX1c6TSi/vGmYFJP+jydQLS2N1+A6Trl9
vJ6Tcq1kxiNzZyv8NBfA84uNfEuuB5kU480pXMdu6doo0nmF3hfsO0DL4Di+5ELs
EBB5VUzDChXzqaoG05ULk8hd0Z0b01aHgeviS+rNn2O9xDVPG+BHWWrFB6JGV/yv
6cL2XT4b1UQflHjGt0csyjUH4gkJqmVlKkdFsxk5ed9uq5hU7p6rjJu0DM+PMFKK
ZskSrmb3PcggiRBz2nPXxi+8wN/uA9vegSBxgpRcqTsOutm+4/xsM+eMp9GXd85e
JUBDOKbgLV9pEqb3AYEZ28qrM76gtAGVyKJlRfmkVTtiORjsVkbfUSC7Yg3PdAod
H0yvwvKyL4rXBx9zwnIzsovpQK5zWL3z1At0VfF2cGG/gZZ/K5CwvNbW9hnYbuYZ
Ob32ydcz6ipDVoXIqEXCZ3DrUTxJFt6JdBEJJDeeeAfFtP/EAYNWGSdAWs/cSlNg
F1oUQeVdUObQfL7ewgzDgQ==
`protect END_PROTECTED
