`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5TwJ6utn0TO/5iPH2iZTCxFdyrUK3hIKM1HHeao71eegFQ51w/GhFzgNsJ68jvLS
fca1PzQ7HOPPyx6gr5oMmWjmglL7GY8Tgfck2y9w1Jog/Rxg75K6+CJW8iUM3IMB
tc7OLZZi62LQG5Qq+logROzkrvDOHq8rNrBKesJQj/JWKsZTp5s0ngICAoUTURvM
KxfQcv6rFP2iOob0ABX6FFrfzl+MIoFQGynJKRXrXHHlrWVKsAE5Q0UQI4BOHGuT
1fIvdLyaFNohdOmZTqNDUtEyWYIb53YiuOQ89DNcPq7dr+hofXsqSIi058ysoBPu
+aY3cdl34n8gMCdCidCtV0vdqRmfJOCBUk6gQBxM7S6M2snMfnguPFmugLu2eDhK
/rysVWCDW6Z9qimcak8dsg==
`protect END_PROTECTED
