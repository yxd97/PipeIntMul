`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWiQtxaDAM9naK3Lk9Jyv6Xw32NNOr66TN1QUK+Uq3AcETVDlufS8/EjMh4bJFMF
5ilbgQ3KWwpcSIj3lYvThG7mevJoNI8SPkbKWuUexXa63YgPGBQs+J6/JAOF+cqi
yUfVi1XXRb2/ExpEBSXmdGv/SSPuAvOZ/09mPKrpbHmY7tRAdXs2/0zH+Z0joClL
/FQzGSbn77ICtOnPGsPfz6U+6uLPlsgBd4OtY0K4XzeTGOmaUO2sSxaj/SXBDhXn
VMvvBxqIQ83COnfgr7eTSo8LEncJQTW5VSRvdbkzv84Br7y/YOGBvgbBeQqXihr6
NzPmFnKYj5Py1DOyxek6Nr9lGMya4HNvIbPFx2BgEeElRDKW6VIwys5HLt6Darur
VHRzJ3zJw84bNolagVgkdC6ZcX7r1jicorNGah36BkbmiSegHDbWSW6RSIW8LA4L
`protect END_PROTECTED
