`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/iM/lfXniC3D57JjBYvsT0ix1T3H3W792bX6Xo3wl3mh1jZjiGBLSTeI9hkOmp8S
6ryaR6GTd89/asycXmW/uE0iAoObdw4Gfl8gteKwdYp3gM0m9a/iVN9askF5KlHd
txoYeQoZNWb8dda+/RksF7VTVBcco4ajF73VYoUZxDfcpCjx+Tet3MfI62FR9VkZ
0gCpwscYDXZ/Um5DmkYExCEIX4o9TXP1s2qVUeUPTu+QtA2OENo5XLgbqD/UOCGj
FSZ4a1PEDrUUlON7bQ0pJTPOwceB3b7Q+SLfMxfkTMDvwtTYTepISYAM3JCs+fQl
XCBfzKQy/uLhpwZ/5ECbrkf5E6/WDPd+d/Mi7Wg9Bh6R/fEYDzgmkWchzzeyMmdT
qMUOi7ZuPCRlrs5JB/xb1cueOfAsrz+2WKgHdFyiFzlGJE2Z6/PEHuAarSQKyRMe
UQQuFnYFtnbcAqkp3KlHj9RmEOD9iT6TqNCx5neBOoQM/WsmRHL8pr3eaym9xb84
`protect END_PROTECTED
