`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryTD1c1VA87rYCexZLX6BNw2Cj8w9L7wp/sQswNNlOoL9+NSstRWJ3hc+DiM+5zg
T2FRovpPDcj1GOKEh+kyy6IinOEJYbSnVDFwCKn7t4fcEWdSFtPAW1YJNvB84rFj
rc3FU3IXttBe1nvnMuDomEIIEVNblsRNXDYlG9136VKp3zZ2FhCkPavPQGGEjzog
K8Iakd8xJtxeTEDSnC2j8OpHjKuv2sCRD1V9HORxPkE5Q3HVLEN7Zlm/oMUavrTV
Ie4/nW1iVQNGI4UXaV5y31CvwzkzfbaW4chOPF0vRS9rQlwc/n2xr7WXRLHS5BMv
1UdhtcJsaUruZzpg7KJi+IvWdWOZD3lyzYWl3NpZ5NjEoMqv00JJzeRLv2U1ruVl
WSxOl9iTFkxd59EXet4wg+dUxU5E/F5tcluys8tDcaTB/fWpXXtiX0y6027KR/ME
x5+7sctt2Dgp/VcbzVkPM5pSPBaTLB/vBXiJPzxbv8oTPGUcdoUdOXvWqGBRgNaO
ham3df+I/8kVE6L/t/Ft/HXtt01OLpCWip/3FfHmQ6GqhzQnRAVmfip1WnL1khqu
PGb3+TMO1NpMExFTadcJX3Q425Jly+hZ91DFtYYWjnx5WKHwHwn7VcY3cKYp+aZ+
tkVUHhd3RL4SkSQH1ymSHkmDZZzfd9h4ZNiAjyTGZIvn5bl0+14UxD58Sdn89H2k
O/OeRfq1zaa9YiS/d++k9athHLQZYjANK2qwH6+3wcrnjZjptLeBhpJBzOkDuCDa
`protect END_PROTECTED
