`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IaH89m5ior6oLUTVHB1XIS+7UPm/ELe75rPk7tYo21pViSFZRIFcFtv82CLBNeyu
2R62Iw4NMN0HtP3qj3ILhTABQIxDmduAufb6Nqqp6g9K5hsu8YDwJcydHyct6ItC
u8Trk5fSCwZNKGYQ2m3HANGn3Vw2nOJP7uJMAQh9Ei/KHroU8izu3ibD1R/qvhE3
pgELZShz9amyCbiwm7Bcb76VNIAzqwvyg9OOdq+jGw4aHnAdFTRiTZRivF7oknjA
DtRpNrjCz/9FTOehI0/QqzaZwCs3IehliS54WTEFtjO/VM8kc3S12LkgtrCkBSwG
T7uIMx3yu5ypsMerTpuzoUJT34kEhMDHUTtBAhNM+348ussVny2excoRGoPHBFYD
UiAvYoehdB0FBhdjMz7usA==
`protect END_PROTECTED
