`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egqDBe0XRHGQRz/dInImQZSC/lhztEVXokkxp7tHOsoY+OglP5ka7kWo2LhcIsq1
XdA+McWFylRim8uWxRBkuSEmm7PQr8JLsl2BiMK/UnUStSHcZAdTOQ8HMq5UtoTK
KOxuwIQIZrn9UZ6YaHbJU6LlX2WDxSHcizv8iZGKek3cDUbXyF+J+m57iwZoDfEt
xoQVJuWzYMmAIYlMEYH83QT9usg7FENyzrG64nnwrFmwXpVTSGzEazoWlpIaf8Ss
sNjC9WWJ7khO4q5q7sdv5xw6gogbAGI7Lr0YbEb8mPITlyMJBvpvylNR9a/cGlaf
+3K12vsmpTPVN2lFoZoZcmoP28T2KVrM73PPBgj7ukBRI2N3xo6+FT5BgsV/wGG9
g74SEL7IAlfjV2+MFH1wmsI7HxDsTDp8yrRE96RdKqFiZb0Kx0AtjR0TXH9fH8H5
DhNyV9LXRtUnYnd4JDGAomPzjwl/8eTQRK+8o5n80FuzMEl+BsvMJvliMKexZ7Bv
22m+Oj+u/eqt/jKwQN1E9nJ5W3fo5ZxOXNe5Ttv6yaPvs9yRhoG+XtL8uZsJbRmO
Sy+myj0zyrz6w7E+m0fRfPKqmnWxWwLr8mnBFsewxJEa9mDgEZOVCIro+dDZ0Ucn
/xocRWcO1pkSGV8K23H9L8/MQapDx+8TiaOBH06y4JHPHdqN1JJc852qDRFLFb5d
ynEp2gFEGjWhx7/tFMEbgwLdF4byWtXBJuwtcJD+F1xuNWq2cHI0keYFTL0k6nxW
+1gynHJRYKOLZjiT8Cy/kACD7aikI2IT18UiKxzytIsIhMQ+2yo1Pfhc40E0VaiC
43cPFe/Fq1aZ2B3o98xMwoBSIrJTh4EkK5hVgkVqixcD7sZNJ4z36clkiLpqIfPw
x55OoMGbILPC1kyJ7s8x+dQbBhdntqktoDWyxP34wn/TaKmTkqh7hQQ3q1XnfAIa
AKMHBwSPkdJM5hITPz8M3QW5468e5Ojc5bStONf1GQWx9/uoO0f7+3GkaE+fvC7x
DHmlv+PVFWvaht6BaSDMpxyfgUjIWNzcM3oh1OduLDBFtz9GcPPG8npDII6JH74T
xU0mAKSnSXnIw43SbeyRPxZfdfRAgWkKKE9YoMlUPqaqQSQ7ESr+EidMs/JMsdZW
ODFP+PL4dL35C2VLPTLY2fPJPJ9rurgqdUScdRlivGd/GSlxL4bbKi+Agdy9XYGH
muBq8AiQWDwfgIT8et7/KFYhahx+X5m+l0S4IsV1ch9fTNHc8tLYhch0c5UpYLPR
`protect END_PROTECTED
