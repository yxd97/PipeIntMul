`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3TZQ6A22p3rmO7QR+vH6RetIsprsD6i1rgGAkpUjZJxu6EvxJJeWVW6yAQrBhY+g
TEIVOM6mshY6w4+mkcfCGmrTf0YIViYQ/kaQE7FG1eD3rsU/mucsLpDZdZCByXZS
JFeJ0YHSESeWnxwE/wDzvFdIWFxe8qcp2Ekv97iq/UUgq+YaP0Sl2wxYLNW9Biw0
qSJQUmfXOrrS62q58gdpIktSfHcjNpVvip/GHw6cN9TjCORWRtF++OQYGhR8D/NQ
bF4zRmqflZQkJQEBLBUx2n41gRp0gtJ/jDVKUm0uRz0HuiOj6QnKNNMue2T1uOHf
fP6XEJYIxlJXW+/kSa+sL2+RPANljnrAtI/9o9vOIfYqwR+LB9iIl88/ZYlc/5AU
rzkDxMpYXrbR2S7o61tiMIthM3lJiGQyzE7zue5oZKY=
`protect END_PROTECTED
