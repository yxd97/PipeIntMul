`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/PbxGyLNPmN1o/zn8ssu66er8VJPlPHUBNAyobvdkShJvdJ6zMVvaz528Kww6FC
zSqzaWe6tNGBcdFPUsvLCNFRWQbUj5pG3NBCkfMVgbug5B+Ijav6sFmQC1D6Iouh
8xV6rERm5/dAHp4A5RBpGwfoAwSZjGwLsqjjCaxfyVQcrnG6VP2rMlhEZt3OWjgP
FErE2jp/nB/o5CyU/6E4duMDQL/TCfR+JSxTSC5iQBTGpDvScmwAAb96U+b4lS4E
TpjcpjYl+jf54uleRZWrRePjstFhPBUPO570CwiXM+27Rgl0BBOupq61qBwlzvjI
1dqBM10KCsJHKlCr708S1zAE3U2KDSQtiTEuJXx03xqh85Hlx0NYZIo1cnzwc2+G
hP0ythNiFly87oSCcD7nYcyQ+U90r50ZdBJZH9a9R3/+OQElGHvPMObGMHxqP1jt
KtrXm5wHK4kmlrjmYkW5M2HuODnG1gcCE4femrqiWJFCwedmIY60Yx5dKXsIm3Oi
N7sUsOg9j9r9rTg1gp3QUP6l3jf5rxVHU/mL/UkWfhXF+rI/NrpjaS4tv1yOQhtW
60Sppi1KP+KDyLjfkd7SFacbb25d63fpogLBwgMxqUuuqpptSNBkTjzVTl5YdZ1s
DYZdg6MzoSDJrXAKoNn+gQ==
`protect END_PROTECTED
