`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8cX2LhipudOJkpAghZpif5friPWh6oEb32HqnnUIDnfot2YpXKYAk3S1Qjl128o
Et31VlwrqPAZj2rios+zUJ2cTPULLIFk7KUY9LcjfhpmZZI4EKoE5wbx+G5qpx1R
uGeye9RGGBZeoT3t/HzJUMK1CL4DTTIVBHrfBrO9WI3mfkVpRcj4rdiHNmf/BRZf
yALdpFZPH+n9YQE4LchujAv5WHybC7yZgdO+6XF6Srfl0nxCn1g8GOWm53Rgi6qD
VfLDImfkQ8Uv/GjpzB930r/blZ2uZPrph4eUaqS2pGXFT9k0J8aCc/pDSnF5aRWQ
yKUMygH91fL6aVt9DP+kHIYWqgdz55K/s5QYbrnzETHDlNtXmhM9hqGIu9uzUs5F
hJS8eLNDtOfsl/4Y9OAsOm+yxybaMc0Rg+9NAXPQQWxhAdwWFdNb4cZ3VvOPxzp5
1k6ffAKSgm67D7yCuShV0rYMuHfFliPOM8RktcZCrWypq04DM3VEjr7OfjSIpHy4
2RLeFS3MQZU1xSxcPKnd8QZe2dvrlF04pwIEUG6KJcGxZeUuXF2Gh4fHSpb88U0+
CodrANQ/+D02NMPK3qXi/SnGnD9J2cpidu8gt/ugYelmdtXPlMvJRkZMfkqRIWQP
fV6FCTw/v9It3HsZVSZTcrXtSAFpWPQiWCycQ68S/jqBVy7oQZiB6sGTSoFepBuT
TukGaHCj1Vt+o86zp5FGrQaJpjNzhB4EjiA7v0EGfvyqc0hZFi72/MKPLnB0TW2c
N+MdTeo+4nw5DSzZDFWq84FEHwfTtZUQ8ZvWLjzgaDn5kG4Z8xZh+C5migNJiqi4
EqCKns/8M+DXL42mVmolK17J9F6j4PQ6WoVuUYbBaZh6ESbeBmJga+IddrxgqD6R
wu2aGgcptpSzvvDo5f3HfboK4GuFb0BYZ6Q2u5mmzEchAUNzYBsfbb3TGUy694EY
GlKabNtcXj7FFCtrHiDBIZaQBPsH2PlMfEoXvHGpR3ONiG7vqsjQa6LljlIJL/ji
3pmoLFUjcNb4oWCYMRLDk8eAWP5RROuUm4V9TyXV1tFXLm7+NDpzlOtcFFhuQxQq
oCqCU0oJLzJnaR8I5y61Dlay79igD38G6FnHgerbN1f4tKCgw0r96KmZtdml6HBi
OVcjtuOW8PkQTZ5XV72LlAFTylEJrp62wB3L/k9guXIYss+CeArHBamsEsT1Agvo
4/ETfwlyZgpeLFM7laQsBdwelasxBJG541YZhplk6HF046PV9YkMf+VKWQBAvwi8
uJiuCYDZcgIBhIoH/74Wy5VYShsaLmh7UVvJS3pzxSyn+Ng1rkLreRdn1Q0rtB7v
qF8kZ4tJW3G7HeOfjIrE0i00V+hzo5EKgLSov7s0nZBnD2Cr/3qOe7t4mLwysUuc
qW6Xms8vekFWmuk39cmul9hP8HX7Pweo5OxmfI97l+CXY/FPz684+Nbj/J9IME0h
k4D5ZxOxPD09eNPfHwJ+qbLfEOHecYMk1OdgQozruJ4y3THBh2FcANqoStFSzHUq
V79GjYsrR99hxs65p0lX7p5KPndl1w7vw/DRYSnBMqL7aulGRt+TwLmfrn6CeGzA
NAn3eTAmPX2TCB4u+VtxFmzfoQ3IX8tz0re9rlrQ7032lzOkyerUxjF1wRvMUcRG
QaLJ5HsZEajForrQlOGoFnpQgIfW9ugxBnirtsLmN4B8iBAZdogLwPUHBgBj6dWO
g2aOgcgBP5UQeAOsC/3y/fjIURKnziOtj/4nA/NFQ/3xrxRll+Ij52H+dV06bXav
P/rTueSqF/a8k4aL7Kpg5PBnKCWJAPPM3VkKkJdDt/hsUhFw204k5xQo9pPpzTm2
58Kcap82X6yjaUlkf0RWMrETc96ZYE4MXF4vPXmUTWo6Q6YUTRn1QWLaazlDyDD6
X7K1dSy8Z5Qwo7tRXSObSPKhL16RSFsPCOR1wFODNvhTKNV5wSoDMFI77DNOdfCp
Z7tSJAmWepKpkqLEMJEosMf+ySBzWGjNcW1qi+H6O/KgpSZ36geap7Hr+JW9soP/
cYPPzj8HnTxFFmNpH8+M7iPNfJ2UAAQIpEF3AXzKVxHbh7PNDTmORYPXQKhr0Ehw
VCGRi9WTVa/22aCRAcZeyf7QZ5xzmjxol2jEaGbAgAHQDS/tOsJWZvwctP667DJg
eA1wmkNA6cwlYZorrXASG9L/CiGQRvgQgWW2CN+bNotWtNj9FZKEtp98DzAPupTI
JkDrGHjxvgeXKlAX95THPf/m0QnOBKe2aDM3ao8nTLG6aK6xevOEMfEL4LbGpQDn
mthHjBxeR9Z8hMqJg09XT0PKq/ZfeIZvNE+wWKUUGs4Nnah+u7Qo4gShMGMmbVjT
`protect END_PROTECTED
