`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xa22eQYvJ9pNu8XHb4SwurZX0GMGHUnV+sNRagBRHQ9TGbVneqQDUv8WWt0fSUF6
4juIbk8tXQTEs5UaixtdnSwRFf5VvyfcXGCeWIsevln4PB7jRpeFjYSnprg0qRii
2oer3lC1WA94GaClUsxThPYOKQB0du5KqLc+38+fjXFzPlEjTY7B5j8Rh6R/UPGk
mB7jgQAY54P0yJW9AfCDeVl+5UFADBTgPaGWa7FbTgryfKqPz3iD7XogM6pDOQ2u
oKVSkxPT+2Y0PFtCbS6wChsGhxGUNu/Ka98WkmSiIgidhwgZrwiQXaXe5W8wRQVX
UINdfAjvjTZafl/Dagl5yqIgVol9VFA3tS1PMftohLVyiRqBJj+D5vAFHDogxqIt
sXMNUmfa/uHil5C2+YqM1R2jcS7vckQqufxIKac4VXf6BLvAbo36ezv0wOFNyA9S
jGn/qB22/AjsMAQwetcaxOTalXs7RZiJzgi8qs/mC5/OzLrIWAQdsasLE3qlOnX9
w1ohJv5Anvq1t/Hd0eLkexFkWoAiO29xqaAyGyx40tdu6ytA51iOwklX1AGZZx44
9JCgujbJRjX1j/RJbM0iGE/H7I6FQvAL3h9JakytU0x5YsmA/0Pg90H9wxmfQjuu
pVuYh0kTpEsn9aabuYNDmhcQjJ2UG90qI9cfJj/vJUAJIHHAX8iwj2eFLJzWAX/N
D5mszzut+JG72y4xBMBx5+5a3jEarDYy88ku02dtW3KYIILG2wWrsxBGys/qcuzg
Bqg3lPQuX3Om/sqa0uatFNKdJBoUIVk00/2El0VWWuaCMIy7SsR6lHwMFznMP38x
yqwWtFyOpCXP1xMAJ8eDPV51koqOyHG2TROFGtHuogU7UOTb4xelzP2J/C1sYgca
By1cmT7yuIFvtRF4ikFSSqJF9y/QwWk91Zlock4L7jrsBLhzZWxGqutndnFdhumm
QIg6a5Ag9QHwH2+SrUaNXT6atO9eT7mqynZKqguGuZg8E7coiLrE9Ai8u8hN1nG/
dip0G7OIKFM76nUMeII/wUl6emg7/y7olKD6vSILCXRnNrWihMWgi2EElbN8c8Y+
UTUjM9C7WqJ9gyzXqKURo494lYbxsh6OsYdC6dy0kRohgEju2Lldc65fAIcSL7Lj
eFVGAXIXG5ui1pCDkxf3tB7P/SCx+A0vBfiPLnXbb122TD8KPUQnPBo+IIbezJtD
YCzvfzIhvhiyJ+vaTb9uquoCbNMjY+KQ1Q9v6J8HRHIQdoXFr6sN+xE9cvQP3DVj
gLpCvnpGuaWhQSD7+T9fQ6Y4PL3WLOZAU4Gx4cc9yboX0282Bz0xx0Jp3r1Mi9zV
LjOONI6+oRAoXUG0+/A83i217ixKLUswhdwn/nNyQNGahFugrlGJJuNH3XKxdyIb
n/5WWhhlEMWQNnbJ3fRqwKBeQOuDIAyX69AnrMA6vwZPXKFpcr7bkqDQL5VZYXk2
qtsRsZd4CgnwC0y14Db8/saFarRPLbHCr67c8bZZw8SMCgoRawfYpXiiXxiOEEiu
bfoW35MHat4IxkrkwjuvyNGPZupeQowSxkn7Ygd3Ivo5saknE+f493CR2vDi7fTn
fUgbIVKFGh2ouwl8rJZKiK8SeEUuo1QINWCaWBZj2AAke8Pa4s/NlAArZBV8lULT
4j9O0spen9yJNuc+VPyDzyMmoS96IXoMAVuZfB9f9Xbc92pPLAhzLHUd2xN1sPxI
Z8d7YJ4djvs9xHc1O3YKAxukKVLTMXGUH0vuQ8svX+chQPdwzBuF0SwRJsDN1YTj
b2Qlxj8eNdOQlKoRqFZ4LFgl+9sMvjvxM+C45tujfr7HIaEddryME3rTnEChkIN5
Trs7mRG5b3R0Ak0Cw55eoqolYjranAWa7NuiCAOd3WbK5TYgHyEm/MJGU5HmG1y5
5S1tyXYX66Qp0ytBtEbnLrQvGZC9BaPqUH5irI/EpddxoPaIbdSygLTMp2u9gsKW
5Xbe3MGB34iAgQytbLyO7W8ptJHQDHKdhjiebkE3RuSRHoEzA7jAi0u/fC2eksb4
3+m7gbrgCYUwSroVBRbl3MS6wKhhZhOJnrqFPGmgmFooUxXt6eao933r8JlTXWB5
wqoWc5blKR7nhreNE0Ogo5hdKU3VufysGAx6qHpYpy2yka28LcKkHgCNMQ7hWy0B
jiKKmsmRm9sMQg71tdx9Cn4SMnOLo8AGr+HZp0X8UWsUzN9nccJhiGRCEDXEIkz1
RUsQ8ibkuToa/8Pj0E9aYwGWozLc0eF0OSVTrjjy0sBTB49/gs+HJTzDKiXluGuT
A8xq4moI+Alt0GnRQulTqMS0bvgaxiss4ZMdXbYsEJ2ln+1e0ivgGh+hL9lGzXZS
0DnXUSmW/gtwc7l2v7wcP+UlbX0tqIrJhPrdZOTeqDENdD1U7AHRu3C5nwMceY5v
OJAuWEABjg3YlT1w8Dlc8c6yFqu7mU13C0tSvPIVcb8=
`protect END_PROTECTED
