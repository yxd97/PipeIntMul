`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MfaQ2Nm+WsVaa7xrQ4hQzPDVMUQzo8gr6cVEfImvFHOLj46eVLnilB7jq91benzM
hbrjjKmxujedz+PxB8aUGb2nRZjuIYdAenbS3SP9eRbE4tQf+91Yh5Q7A3jJ66Pc
AH1bRhY8b1dwclkzR64KRgeA+/hXSt3eNlB4STH9JGWvyreq2zoGQsbkh28D0prG
u5jUPVwFtUc66bXIQJgr0c72jcqDRWkKkzOfH5e6hYk7qc33HIy8KEGls604sbqS
2QgkPE4kJ64evBjLCYUgC1tRpzA/0S+iELgbRAU0ykuv9Gpfnfqix5XJF1HtLcti
PAVlT2qGNRdf7s+1ZAKDdpP/LgQg721yvmHvHfmRNm/AsDeph5VrMCGsD7TIex9n
15y8e7JkZzsr7OjMZg2vDhA4JeVZneZLjMa5TxkSFDufa5eYrtguyyQb8AbyBMPl
Ac9NjbrPbQ1TrG8L6Oo88Q==
`protect END_PROTECTED
