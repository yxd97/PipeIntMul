`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fZ8cbzeVXmwVWmkH1Tom0327/Mo+roq2d6xpdQ7ulPMg9abLTLPD8W7+S896Qs8/
LuxIyju3TISr9kjsoUHyHjZCgT/NU2VRZd0BV8i+0hDXvo6kRwmp2+00HGi68pWv
j3+5c0tQEtFaw3AAJU/VWTOSBUl+1ZsOGpzfLwVIYSpkksnsOQR+38wI6jh2rVCP
nGWnj5WN3wDGuXSbc8EEPJGhGOSt1Qz4hyqJJNfLDCvS9VMtcc2zbfzOi7o0tADT
uGBOTiLjgpghKFyjhVU/i6DxxXsiXsWl8GrIvCkxpDaGFrbrJiiLTfh7qr9f/zGC
8Fus1GhB6EtI9YlGewsj4j0n2a7aI/iLRFwosL/s3Kxm2J/VqrAp1NfnR/ZLMgKH
hXPdHer0KIExT3S+QCwbVA==
`protect END_PROTECTED
