`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r49/iCA0qEPqWQ5DFaz9ercZP1EhrTAfuW5Y5GiVAM6XywsJZVtmEyB+ZW+j7h5J
qNAbtfsLsZRmp9jqAgYQI2YYMtZL5vNclwgOicX79/IhuSr9BpNgoIIYp5E7w3nQ
xeWY+Q845z8TJ1e7HAwrPij7sfcWFV5+Zf0B2MGFj56Uym+o4WF4QyI3N9DeVIVj
PpAJznbmcHU8yvgSznJ4YaqTB6vXdVUOqvv+P8N9l7YlCSNsd4BLdfXZr1+ffJpP
cN0NY8YRQ7Lsd5C1uxoMci11YGTd/T9oSjj9dQSMVaVZEdGfR27d7qe6xC/uJdxc
zCyfeF0iRuxKEBtxsTFsp8eSe+oQ3syuxdxmL3uaGvZwCRiET9OWzpbRn/IqSuMl
cvIM2JXtDTmy7eLVVnDeMsXCSYuO+j1Vk7P86vw7HZwUsmWmVBFHU0AzBNTXS97H
S0YtEiZ0EfIed2mf4bSGaAFjI34nTZAxUH+UZ34/2rBXEtWVP2AO0LUe83nOpPqu
xrwHvUst2cwqDc8ULMWjap6HVJJXV/padJrsHIEg+kDYvFRONiac3S8ZxbbT0jPW
Z9KvrKyPvZcTyfQia/Pi9iCZ+OjBlGVHlUR7GDMRMrVafkfizXwMG/K1+7ZJw1Nv
90e+X4wXpBj++zqVyJpZfqCwIsg3gM6vPXt1UszQ7O1Rw4QugpbUjiqqjzkBnEfn
9SiUvtlw0wYzNCe3nFn/4KMIqmGg4hAO9mMvgf7jZ1ddoUQMDsMNR7GovnOGUmVu
tmXshUnsq4TgWaHZHd3jwSM0+BfWRjw9bD0DxkbjnTUkNhKhr68l20lDB6rIZDEz
HCEtZNUmqPdgn8HilQdokqGcjtT7yE+FRIliNDjuYtVOM42JzeBnbChUGIa2TPGi
P92QfQ6Ui4w4l708H+GVfJ6tkaEdq2J6jHWDpjT1+vCJL4lIwBWfhQxJ5tns4ID6
ZHAVE7dXZZgD6u+v7MwTaw+dMjsOI1Jty3CRPpOYN42CaX6Mrj0leIRFws/yEols
l0CnM+117kcehPJwzbZUYnsEcNGcpGbpPUDUzBJGRMqokjw8wDg6mc1gPNSFrYWG
kXpVVH89s8uh14qRc5BBbrkn0Z+J2FQvRihJrdyszEoPjp2QFmUt+fikCBMoLJGc
Mn0AhMpiK1DyejuqdLC4G9mptsrdBxIJD6NKGwqKC5ShGfPXduarVty4t3PSRJga
kgGRufxEQcR7aCBIyreojFEdr6rhvj24Nphzu7kDTeSyPivzqCrxcTbcoccdUuBz
s/kr9KKwdmZBOgN9uYrUDsNhIzlRyFuFiHoPqHXhRRlMW7STKagxXlrlXD6T8sdc
rpc2g3mKduUXm0vTsKkoZBVA7XnMtr2ZYGd8M8foVYdfSjoXoRHc2TGamGca/kHU
sYHrw3IHBDxbFPU+3Wfs559Om8YQi+r9HK+JRQjzGK57Oxc1xjxnrzWmyuCrVO1E
RAEkaCcmxXUVj8Fuj4Eslzhxu8/oOItaK7XjaWD95E7FBetUFrIHm5l9FT/L0QBx
7rHz7twjJx/4HUC4pSFFaOA55NAIl4l7SM9X2OOsGwy0uv294hObDWAYCbciHDW0
QRrysZJf+qPVBgf0jFtDgEFnBHwOHgl/dcFcUoNuXFx9zqPJfRF28ExW5FH1gWZ5
wsbBcylU+aMSq0cCLdRFklk0k86ULHULjJYLktut12Ytp+KCUgqtVfCVABcWdq15
sCwhAn6eqBz/rJMIAHcaHfst1gfSXy/myKrJWirntgBmYjtquYau3Usi2Ug3PZAu
gaHOz2oQMWGRbNTtlAOXvnG+X5mo5Du2AVQcMH7B2Q1gQGx92GGeiFeVdLXheo6X
LP+PcWaFdUdyevzOgVaarwWbF3EF4r0Yy0FQyT+Tlj4cgomTjWhCiR8g53v/vFki
j4CqNIU/xTNUzoZplUDfn8QEozjUKkflHVg6W4LC/MjSvnUUvz4JzwaWg6QALywx
jlPgsDyTu7a3ZOv719aRahLtXpSzf8AW1SnB8H1BPc9SXe4nGcNK8BoPex3+IiaJ
solEeAjeluxuB/5EnhPKy151BOoyxXOlDrLkQCf6bNC7sOPk9SibOsMbHnGMbV+M
/EMyKd/kKKDKVPG37LtIPKF0eRgqzZsRM3KnliijCwHLiRIbvxHFACkeSynM4aMl
UNCp7FbGmXUtQtwksvZADn3PHo5cgck3VRgGc4TCv+f+TesfARLsop+9pX8NhskV
OUeW85I1LmwLerUO7H51fsCQ8Cfn3fIDySFqq9YNoEbq5xc6Owpl34o2FBsS/Ktd
f7cgbcuSBoIzII82WUGYzroGo2nYSapgJ/ewDISZeDjGej0EQgfD0nQuE8Zz4lOM
/NCNMhC+ugQ+BNk3xMAMoJ7QaqFmanttc6UhpjRlKLOJ2PitX913k2t5Cuo97CB/
xiKIkaCSqnZTQXEyK5ogDw==
`protect END_PROTECTED
