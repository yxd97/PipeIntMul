`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eAxYyLOueWHN+rtlEw2Z9FrYGdJCaHzIZYENd9M/NqL4jEOg3vfOkpo9Rjumgfk1
O7VRCyroPIrjxg96w42mYqbGT75SkI2IjhOxw88mrbOGQE1zq9+NlTOUihtAwYZ5
HqRarWdPSvUpXCjAKI+O4W6tgbONhM1H9NUa/b3jnOnNnWjo1cmNE8r1ggMubFXg
BwU2GV5X/Jfajj8HMiskbYmL/SmOW1a3oWVuxG8G0kJnentnaaFMDl3L3KzKC+uD
XsTxMUNdZLQuDlQjHyRTwoFT6aYPRNMN/fG+PCKx3b31Ksdmx0NMVhg+M4hYlWsD
QE0/EfM9uJ1Y9qOKaIefZRGBoGUE/RtPc41N+LIPqablAVBsSXEhEeg1tCxxAlxB
mVWoz1LLT+enrKGXZlXTmWdvynvRqhKtmBFgpeNpIPZUS4WSxwtKWat9ZtSS/v9k
XgRs3TOKd6IduoQgrULOeOfPSh9QMayKEC3/oHAYSbqsmi2yGS19lytbSB5IqKpV
2eivOpzF5dZgRTtfqaDkai4U8BA0+hvgLVDmIZxq3ZOHWxQ8ESJBgLhxoK0wugkN
ht6nb/fjmpMBekRYorHEQ+YvQ5Wy0gxabLvCqzu/d3myYc8yw/5tVzZrI0+gvUhg
TvJmGY5Zehmw1zPtKyfWrXVn0V8WDLpkfHRZaPtb3NWLhTxbXwTtucKyov8Qro4g
MBKm7Z5az95EW0PBN1crRJ4dczbRVsAejY4EeWwihzHlTNWkueEfC09FonnSAJFL
ZTQnAX82B1TPfgRUKb2V6zvsO3qNSac5DY5HWHskstJt4Wt8/+tC8t+y+RFAZ6NC
v2/wJFV+TkNlSApA/ZTQerevryZ8dcUoIwRIEdVBcn8CRXggwtzTW35txwTVEJT/
IZCWRspB5DXueIv9tdmvZLcfCOrXFas/6T2s4++jlbUZUCGDGTvHVoNVQoWG+arZ
MPi2I0z+paGEpv0/beumeAFK5TjoiMoW0OIV6CVL12cPQyzyfjh8NGbM4lVjS3vU
NH60TdtaaInnXsxnEbAv/PYy4YfCjPJUzWoxDIp0LVkZ1ZGFrB8EArEaY+Xw/upU
YeliJS7oannAatxMtAUG4QjxVbMbfExas88yX1se/GBRqiVwWSq15IEFgu0WhjZo
PHevm58EeMssqYyfMeoTeXVloFikvgUphXZ+QdED6obKLvHSrRhS+5pn6flpUods
QOEWKsjd/x12sbBM49U5b1wM9UKQBmE5FdMYXxBwqec7loYi0Z/OqF9Yr2i7HF4w
ft5xvlIRiw+ZetoA228ynhR9DWDDjiJjIcY5nqx+MUrKa804UYtKkYBbBjfNanfG
1t2MNLALwfazkIWq8iicW8PwcKruYXDnDn/wzDuEQ+doiENDi/546US3yjmYMASP
aCI0pnLJdLUoZCNaWL/45gjw3DBNm6hS3Nc/G0XlYFdphnTp6Az7LnEFJ5/0a+AF
emzFCTOOGyPsSACJjA3d09L4Etni2T032tYN52g/30c4IXXIVlr7DCtkaRoqWepa
NaTte6dMdYWm7+8Q0LgO5izWgZULGVRcAzMebdzUe7KzvwoUBGNfv1kP5t7gknLy
oOQmgyM7n+5rDrj98FLIwyCu5RfaRccaKsRYu9ufhqaxXrzylmg2KQItfNZ+xz/t
Ag6+KFR0RrswGz6FXLlhjM91bld3Mz990IMrs/bBaRR4vGg72KbbuzJqSnLFO5cc
veNCKUgemsWNUdFU3cMM//Fd63HM5A57517uCxt/tEstJ5BWvvaY8ACpRPG+WS80
FnHBcZNNiqk/ebC7j3uxwqDQ5e4XrkvoZevOc94iPoAeCGOgSIdwab7/7kOtikhH
56r0t/a1YK5V4DSgXkmKOcTYBso8skvVr1PyqxuSHHY8ommttl59jnniegyljkNP
ZD4bLholnmnqbwSqAhwz5UiFZIku/ytBfisLATWu06ubG6Rb38Cdj5lyXJG9eAos
WnOzghniR02GICSWoueQvPcniNyYaEevYfyfxrCr4KqjA1MSo0HJVDQgmV6a2GPw
8crixnxBoyjzxvaOI/QDAUv2+dJ9A6+rzPAqndZfEKPVxWwMrAR8eA+5pJg1ZiUj
6Xd8wcz9/GsXDG53/73GrNhY5NjldjBoMWKDKugpPDlb+zD89wL9VzpqjEgTAMBW
P4HDwhNpbeyD6opSR7wynO34Bg8eA6WLc3ztuOKnfTGQg7hM7g/HPhCZOwtA416V
d4XtLhpEJx7HMuEr8KCTQSYeqFfvTl6MbcZz9f9ATbZG/Cm+TRiba5wav4Wss9AJ
iz8GU3s3eRbfN7vKToTdMuBha5PNIVOHr3rLUyLNkwdYjNRGcpXqWDjaygVcOj9V
+J6Y3dubL/WRha5zNP2D6HBMOEf8qRTYwzL4vqAQDi+h6ocIniW5zvtvfvsryo3C
FjBUazEsK51KdjuY9eTFeBbqkrpxdT282kOvHihPtmuXqS6GCeX7jMVxhydLuokw
GkXWuif2bQO/2OX0L5acPyyC/NZiY8+3RTM3WAm1CQW314v5XmlYbTwd78L6Bstf
`protect END_PROTECTED
