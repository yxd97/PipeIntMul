`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P86YMXo+OMli7W6qI+NhIoqzFfqZfNYFgy56HdN9rAuMx9Y4TPaqMQUTQD57OL20
pKKD0gVtUDtHAQOfHPviiXUkChzE1LO4WrODV6iavZMxptbRNu7qZScpDwQM1Ua6
gsb2+AhAxYSC6KBwswITQKijKrc4Ty4p8CLYgMW3Aj7bzmVV1sW3tlWmg8HKJ5MG
YzVy4o82n5LkpGFkqlWiKQUP5RbIXktRxvuRzUgMRXQOKK7zguEKws46JmO0GK6D
pMgXL43zQnqAvO7CQGSfSzWPBr+SUwcp8nuUIbALaaKgkiW8QHiqgJOZnGM5dEdz
IrGEVzmsYPLIk7Crz9aG0dkzh+Pkpfp+dCBc2Df6noH4L9HAH4KDLV4hW+iyiwdQ
TtqnYbZPKGHABZWlVjSi8fs7FxlLJ2yh6o91uiOQJROsOBp55PXzuwb1DUgSO+vH
8ZdhNEiA/anE60SlvMcU3XBOWqEGNEIuf+/RJ9EEA8EveWm4jKoMa+ssUHRaf04X
PkznYeKP8z2qd0XK/FjKcMkujIvZxNXFCT2bNxTH4P9ZhGCD4Hw342PS8CDke+YG
IODEg0DT3Fgxcr3DxE9LHhfF08IGhwQeNEY42pZSvv/TzPwUVBUBIqlXHblcAbpl
QwRB4oXu8xT78HCBFq3lUYhZac/HYEs23TXFwfdO6QnU3Yt9DVRPmxwV8FwEQ3SD
tEReTc3W4Aj3FT7qNe5plXusWhtEKfwIINyfVByrepA=
`protect END_PROTECTED
