`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rz41UH00ZIoK7+Q+xQ9s/ny8bXasOCavSsFI+IY+naBd1YBmEWCtTHoiioRAzbjH
IUWkOJwhJPEl4mX10SB7Wnb1rih48m8/qs9ceZHil2MX5/zcAVe/GOfB+VLmB49p
IppEUdLV3IgTiRjmGj28LlI4s0Lsz9J4mgkpEDktmHKzmZv3Q9JQSdoj7wX5gxPK
S2Z65gNmEPKm754OVFmBbXfkrWWDU6niXtiRHV3WKgQFTi0obp+ORvOKMoFYJCUi
eioiZ3YiGjnmRuxbL97A79s5L4L9TMI2rFvUHRJ+KTEG58xdwANwo/d48I7gNi++
7zsxUfgxTyX2u+Vp1Y18q+S5ZnHjF0DGDO9OEB206m4=
`protect END_PROTECTED
