`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8hnpiDUvXk3a4cCiokDLa7Tfsw+iupRCLxSJUOYnf+OUrTUgQbXPdKqXLnHx/WTI
Tpe1P7bt/yNLluoIDIydsRiUQk3YBPwP4We4Tv9LbjC1tfPxM2OthIpJUP5G0iDP
YpIyWigQAhsf5EGJe+VW5huhX7xxkRCZOFKiyjh6UJWhYyB1KGBZs1pYDtFny0kQ
cqeeLtpio3jzltmSZ6WPiK3STZY3aJyIkOOBmaL/INxDLru/WCURZk+vxT6a0LCz
FxYAhQYDKEUYIf2dwXOtfkQXqPkwVZYYZhTo05awJQY79WU5CIegAxIwXduVj5yl
72venztdfCcN/qbPN7DgHCuy27kSDrxj3W1/8ecnV+5BsXa8tNmiC4b25zNneRmM
o5+s6igTEVGDUVhLrrQTcA==
`protect END_PROTECTED
