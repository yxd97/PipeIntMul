`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nJUre0yJ1d6c5y6VpzBurlMQVtv1aXr2Swuc1Lf4Y3OOhxvDjKQNFHRwhUs1cHtf
TNVlqyIaHB51kie2ZlUgs5XvZ+DPMEPlXzkBJpIKGNKXQrz/JMGZ11LvUIYOlU1A
oyePIP2vQTa5Yj7Uf+XAjjKTLq0T355RmkZvkq0b70hRAhKBwxGOXj1hEey/rdJ0
zra4v4ESHlL7dEJq8c1NocRaVl6A2Hn9UtFB/SdoasJpBzO8Qst2fDbsujeJZ5Dn
fouubI5DIrVv5tWyIwvw4udVMUlBJT4r+ZN0PjFm04v/yurS8XCA/mfNgAMQMpzM
0P8jfpbBC+vG6Vi0r6oLE6s8JAq7l4XgUudYFNQ9Bj1bCNG7Jds+YmmncZ7biIgp
giDmomjIXihl5WihbnxoB+BXoq9C2qpKt9vnTaZDHjEIZSdyZXZkqvGglWbnZlBE
BjAv/Y5OGrP8B0BxE70rUzhRLOO+gEDBNfgK+AjHSsb32+zHctfh4IbS+JX+g2UT
y7zULcg+qwtwEcSurnNhuqpDTqqb0L2WuDL/6TWGjXKXnVD5zSDgPCbBwpMlm0iz
DOwRodrmc2sNlt75A8PkYLX6hXh3SYPD3376OvzZnn3iT0gEfT7Ur0r0V+ZMAAIP
6hM80npCq7rM0QWNrPFFP1EdigJGY9FqueSz67ZSRFhcbF4lWLstxkzQ0tKnt/9H
b4ANnDKj/sINH2DxTqEJDZASb1lGAbzmEF6E6qB9fZ4yKYv5dJmc5bg4ctdiR+hC
aYQotGGDKVomS7VLXPfqifv1/soz6SoZFLfKt0lhKqnKtXFj671tLs3/JnrYRrRl
7sX9Lxi48xvzoR5GPpqHkRdCorpd3ZqmqyY6uyTsVlo3DhCfBGDVkUeMmilxkD+Q
Shv3P3QtlL8ALQwVAktLVETp04eEXnsx/DmCHSYGksToXOhEHocRxQqMsVvLOClP
GfWMfph7hzf5LpU4lkxYV+EiQO6VlewHKMxezxng4uB1K7jS7709Ce8R13DHgFvN
`protect END_PROTECTED
