`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RSS4OxOn7475NQaDccOAgWiywgBKzLBbUZHJxVKK26qKpW14HRu+nZdSGmfCkevf
EIRu+dCVek6v3wHLGbNNe6ocbsl9yJlAlNYLKUnA7EIp7nM/woC3/gw11min8ah6
UQXe7Hz7HU4zFJp3xCk7e8BVGfjG4aLLROytpNgbeBlWLVFawNXUb9F6ArxmhSdi
IgF3ZkTjyFbAPQvnca3+Wx+ObL42Ted6wTbJoveVias4B+sRuZebEaV3JmlRV3ov
DBWZ7CecZMjfBcIpSZdAjLPOh08uds7R6pK1nyZchXSSDJRGhpmyaC7OW+lGL5Ht
pK0gq9fHvPF2AjiE3yP7fdck1enRTzfOgXOykmOOrKpCZukxV+GcH0noF+uGzH4/
4MrU3n2x5JSM6CmKXW8g3bXI3ddWauI6A8/KM2ZMZZaktcnDj/DA/QuCrGi6zfye
sntn+XcE4csyJeKh53ByWXtOZhpofaAPFjuzOlplzdC4cAn7Y1e6rt1bPx6O8D2U
FXJaDfE7JZ/KOYJwnfMqrXdW5xTWpKBsjk0x41dJMwVDJ3M5TTuzw8tCh4i42PHU
A/M1fsMbO+7HOmxIDoPIcM9FxPH1env+ek+FlJMNA1DNcidFuKM/r/oHKPSB7moj
+Sz61ucQWBjROfFrekWAn8DGBLf/njlGWhDvcWE2ERB/foLm3eGC/VOSMildF4uZ
ubOZhSJx7AWp4B9Q25mBIJk6t+xhVG/O8CrU2iw3bKeFghhAVHNV06LIk121HfYJ
pz8AmGrJV7frYigzKxihUt6QuMIR6ouWApg9HlaPJbAUUMga2UT2r1b32NN8dYYX
T0K1hgn5YzPA1Eht36IKkL+5yitzvDlAra2uRbPbutmUjNxs+UdjbS6q7Tv/zFXH
cpnekuRm7G3VWauMb6+HJjKbq6sYspYnLwCGCEmkF6/0axfNOZZslE7kDogMc13b
cTXNm2HX6F1tWQ0SyL0FYM7Ec6kW3RFVS6v94GvvB8/6SSVqAOZzBkRbG4sGeQdl
Ak1iiaHP6UytsjclxKmR1b5V+hcNxtRi4JZvK+9g3UZemMJ9xEedu4O5ebjtx0ei
gfBwrsURciClC5xhdRmC69PfjixzU+xd8Z5EbSffaXUjAAMbGbiH9fpTqDVT39XE
Owmsp5BRsgNEgLDCr9OrzI538kI/Hq5C/PQPep/dv/8K4ib8nt+hGrUTMW5Bi12Y
vUCgXrx3UhNiwcwxiqtTVLcq8NDp8DzkMnnWWL4ssAk9/ZElwHJCAmb8YSYUaA0Q
3rTiURdFLaawd2eY1mzbSipIkmR6X5lrl+0EYr7m19d1dwFFwVtsoNLTgdzDgzpu
ep5m6w3eJXCXBMlu0jCQgQ==
`protect END_PROTECTED
