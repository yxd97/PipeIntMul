`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+SDTYrmVLKkFFKnyzB7stzo0Thb2IGkOSPx19SOSY/fPCYHhCpiK1/uk2Xw9GiBe
rd70e1/9GvEk7lj1IaeXIcV+4K6GAIwsBH8EhsU80omjsqLZFuQbhcptzw90Nshj
Nj9MnnRZgVXvL5LLDO21FrBTvi4qqb5+OHKfbYHXMkz1eY0sODiKJ6WJ211/snu1
0zJlGCtgl7IVmc7K26igGoR85zaj9Dk9m48Gxm3tmKsWQ11t/xcQ2bxPySEUe009
SKUuKNKV4erT38N4bLo6tHlxvFC/LDB5JGYyUgVufSLDpt0aBZmifdfmr5MCPpEL
qhGsWIo8CKWNy11XKdKKgmxB3l7lPYeq1gYzlnh8PUl0BVdMqyfiE2hZHB7Idhj4
KNpGbXtb8aUigMdJ+HRAdVpfXSx5NODmghOCBaCA5ccOnp9L/SpejRbQIGSovt8T
`protect END_PROTECTED
