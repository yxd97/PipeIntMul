`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nrhkiTHcIj/f3M/QDLvKYyl/QHTAA/5sLY/HjiktOcb61wTjyUU0ZmHvzKxlN5Nq
9uCXdkglae/8vnjPKWLuNiEoapd4gp81PcinlBP5arwCEHeEanhVultac/6z/fMU
a4ITSKTaqZ8IlCv6qXLmPmUpWPfRpj2b/7tHZmd7LDeOW5OMe0bFhzndCger7Jsd
M5D4hYYCj3YDWk304m+eSP2znldcPgpVGd3CiL/kNO96hYi7V+gYZyIRZqBO+hdm
OkGyIW4CsxaO/Gz7tZw6axgsTmmNTexfCXAueZY7qmp76tZA+WCmi/63SE3PG186
2KboYM/XT4XBR2LvqOBbkhgrk14UpfNqgGJo6Mymt9nyG75jehdCLRXgKWcuneb/
e1pat3FukajYgYe4a2tDO0e0slzjfz9NniEzi6nLv+3+C7P5VT/51i0Fbp0JePB8
rXoIAxY3hcS88eiDziY00+MMUV4OKd/Bkk1TcO0tSShhrjr0Y7L84E5QdPp/3YsN
aV02528Ico+jiS4XfjMjd6ux9Dir1dHXBShm9vYN2kcPjZa4NRq77fmV59AYwh3C
fA4D8MEHYBTYb34w+sV5wtxnYCeK2Dcqjh8S1xvfiWZI/sSua7TMeyz1hQsnnFLF
wrJXFLa76Wjps7pvGLBjEygN4VEBfOpsebgxIYj3raY5RlOPt0QuLAG3iD2W6VXA
MNJmB8SfR57nxHka3hM7xdH3BEv2AH59Yge//Hjxiu7Xvw8deCmker2uTFO0ikyE
4381bo4ET0rL3fJSopishM4Bg19FAwHj5DFtPq9vqMDPrf8lV5Iiz6M56DIfgMEO
b1nBgz0xWiSj+DhARtN8b0fBHZa0ZvQJQ+uWXbpjzKh58YEyMZg/uA7CJ+h3+wuM
0PlbGe46SMXeAYQzRrhGzFy/jQyXxHkJL6GeOuKswh5y8ydD6m4irt2kMGeLjsWo
+pAjLAHYB65FfetUwCA2CbDdEpvukHeNz1P5jokLhfHtEBm0KJH66+cwYmcx8QEt
xUE3tW1B4zOgdNXHVxpAQImmNosz4IcDuXYgXrfa4yFimcuRhEwT/kH63FPvnZZh
4ZU3xKt8Oli+tlLLhGqX7EGwHGws0WF7iEA/C+iolkuP+QIx8oxwjCMMgUjbqyY5
UJUz0zrxVpelD6WYWUpuJSAti6XftswJnlorqmg7LoHecp1vf5jJ1euAiL6O9S4U
47BcyKveQkWHCMsGIfQFmCaK/8bJrtZm+UDaBZm6QkDJybkhFScJNpFuLiw6ArEb
02r4OG9s4qPIe1V4LRwOnWKeJOyc3dUo2AjqWqeriPaClSio6EkP6+5/yYZ3VVxh
WvA8SJH+yXGP1QYCaSTvDth7wUwITMdLhcMZHjf5Qt3Lba2mgdoYCcmXypETHLuS
u0OGfFsaBg3NT7wdyzpp5oULd7THXQ0oZGAAUU19Sp0dZdbbcoYQHf679XmOfQtz
YCcTp6cSNDICuxb90F2FmxnEnBl0Rzx5LTuG08YBJ5vdxbhWoimg3pWcIVmhAkUz
rZX+HLglDRiTRH0HDq5bMGAJ7lJ4hsDosaN+rbC4INm5kdBsblxcY6RrVxmfh065
bJht2bUe8FMi6sMFZgIBIbLnLbg7RIbdkqKRt3RCPOPfYtsXkllZTP+mUR1unAhb
5zjpzJ/PbBVfsnqYo4C0hLvS3qhjGBf/aSGGj0CeCIHq7LaPq2hyTPXvzAgXA6yI
sBRq6u+NaKYgPiJHyyxKnIFpFMrDBuf7mW3bMC5qQqrLu9gjrTgv2NO0v+/3M2q/
lzluZWZNsda8LKHoP9ghp0/RhkzmlUTtJeJz6w9FC1pv1hPlSfv2JpwfnkhqX+3v
mI/911y5MCm3vRQEYjBPm1UbZ02CI4X9bzpQo3C/4zi0e8v28PwAcRllCri5Jyjo
1YVsslqdyGmpGB43aamhfmHwWO4PHcC1Gv6Pynkg6cqiK6yrS4OMsRQ2aQlxoHFq
XyN7p1e/v/iVOHIb6OZoS4cyty36V5NMXS1xtUQl7l+LvLoYHJnSs1mJe2VvW/97
RnM8vhqTG5XuW+1yHhZYwC105vxJ9mipsmvO85Lnk02l9WuXjY3uwpddvXJtK8b+
KmAXy0lu99rxjsiX0uGreajBDDRzdfi2JETr+CpnHyoo7IpAiLQpnS2BDFV8n9y/
ZyHh7NgpC+w6jewaoh18kL8uE0/kBeLOBMfTvJpBcrLgR5siGXMkeP7yXRBipzek
AWynBAqA3XVfzcPbsG2oyP1skteeoa81JdGLU615cl43bg4EpZaAahIYDieIKg2U
BpXc48tseZd5ko4enaoTCCtjQWZJebZTJaZJfgmxdAHC36G7D6aUCdUEJQF0/Stb
zbHnqdiYxGxTvDODlJA3VF3dUA77UbXKNUcek9rtd6MqN0PwDd4Jza4taoR2bUtj
FNvK0IevIfueCkL5Fcyam40537sB+t71ujq/s6z9F5Y5WQI+hz+xQUA+Pz+Ybe+R
zOTmDtDmg5Eu4HJLgbPFuLvspTyQU5oCL+JUSqMpPyiWs4XAWVc5mj89W3RyhuZ7
/Eddqg3S9HsBB0F9PjXj6YFYSTFRQnsWh3+hy9o49Cd/e9nlFITK5UWahG2upG8t
cY2/vV3/Q35xkyrDqMtvqvPnQ3M+UAwyc8n0dCxbvCBbDwhauHhNkZuUjKhNwr+7
n8ZHGBDI0tHwI5jeV0HsYHqkpLT+CwHvwlAXoMYg6E05VGHUwY1elM4/YvgXUANV
p0JPzGSiheP1Z8BaQLiKeC6VnoutwlJyd2o2r4noB7cxXlQ3wO+T2v2Xkghx7A3H
hznLuHbyd9aU89IHxYEH5rIWx56uxTkFcmVIwIMTQiVeIxe6pu4G8q+4kmAATTt8
E5jQbNolx4ht2bBvR7FGlC80xH4YzLfW3lmd1VAfv2vpyT4SAiEo31nMbbmaEr/N
8Kpny2xSHRxk/Ix/XCBJcEXGdsWPsT0AiVngRMHXmUecdA1POe6sS1Y+HsYxABRr
afk+G5UH4KPIp1rc2cLfJIOsEUSdcVzPwJXKkPx8rtfwdMeS7resj0mG6wdH5Fus
DaHNyQtApg61VzxVl/KQpxE4/wD1CySnVC12wMhwVa+cMfHmJ+BSmheiiAbfGwqn
7TYtID5UUcatCGeYFmCLEns3O5UuiewGzhoigc8Kq4BCpxO5Cm+dNhuKTbmK2MnK
X34DIEAiN9VTkgmKizMSNgKKppvGslBVJZh5PWtJBTmXeknjFMSFKP6sPKWF5hAk
FsZO8SmIvjcnGYasR2s5xSNFYm2hKQBF5QbrksLIeE4bYnbRO1js7MTbt70FU0mv
`protect END_PROTECTED
