`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iLMsRUcKRFLkXhlve9eg3ww4tNzXCHl86JqfHV26VmvtZXaMYfb6L2xAZwwJxqfS
PigbgvsEq5fxTi/K0siL9PjryqLZWRzsEqNkYkm7bZ++OMmZMDzdm1bKSEJes7yy
QlhUcnOcr4o64hg/W0k/Z4aAk/BTi55yAr0cWTwCGVGZBYoNayphY3KV83Sky1R6
CGWI85MjTNKnuhsVxEgnina0MBumlswyN3/gYK0KuRWoSR0OHu7JwxkNlVcZexzP
247N0ikl/bxFrObxjwakuMQa4PgUvgCPZtGiDzl2UXj0m1VvkSFBo0X1cWb4jkHX
9X3P8eam7VJRshzTaE9dPiQcAvJVjvl+aup3y5Qy9FQvD6sUwmeq/TW/ivLo+HRS
jgw5QsBnqXSmbO5MIg+zb7zEyPRzQ+UcHd8Qrk4vTF2AIcwMCjVF6A8D8f/CahuA
inWNxFTvbmb5alramFx5xb3dYb/c5rAryVMWzmIB1d9GsL07qyRNtc3fkOAQd5+s
Fe38zu8eUvARzOFsG0zjonbTaeoxv9FKqkrQoqpNjvrnntpzvMVeUXauLsazY5dt
g2kiuUEPjocbsfDA8cvos1WlilAtMQWVrvGv7o7Oh79BiTpRFolhQQgItOZQJ8ZW
IaMvzk9nfNiL4Lrm3jbx70u9q4XX0pNwlCBgT1Qjxnd6zxABxjhq3kzxdS4UirYF
z1VFM3G4CE+Rk5RKeCFvFygX9B4SQ7rS4Lvlr1Pqu8b0DhZe0+YwWl4Q70UuZ45O
AKZtVcKP/ogS3P2V8/fXOEJgijpo+f7igmM4uh7T3SY448Qj7OwzohcLyf0RqjzC
YgwS/vO+sg3io+rExiVZpn1nbx4M+udl0l36HWYGwtokVgtbXe+OXaKEDxz/JmCL
lioyC56oOCmTts/Rb+Hd+dC1sFMWAbtGSzMO4HMDnEu0JmPE4KBLod2HxFbIGF3W
Opp8ZIraBJUDp73qPhrLIevA6HGR54M8BfZ7TMeIVYQREaWAVhoiHn5tDQvoH7xS
fkQFSpfZJOtxdajzYqOmLzhZ0U478fnN8mX3Fbr5ImaeY7/GS9OKncGag0Zuh6sC
EtDWdV7qx3swCb7opH8jQyKWMWOQsQaxDqRoZCC6uG+elU/rIcU6kbEvz/p99Rh2
s1RNig/laUKU50kt2GOOH4aIiUx2/vY10PXkJm3Ku6jykiWaDwy+zmK/iwZ3ARlf
pZDI4T30qGoi/z3Ak7zMjVES6iO4b1SiJGO/kKWvgiU/j1HpS4H4bH0AiBEhKLfx
FALXCYOX0Zyo3mIstak+I5/QhggQlNKH5jwomXyiDG0XzDvS7yRv+s4eZAM35SF1
zCpCP+RdauhnszJ2nwbpqmKBn2SNTaiOBQqsQsC1YE37P9VZ0heV0+2YYwpuTrll
9wdsq5F4K5ayQDLqSg0h8Qz4Z5CVH+YheBtDPUnqfu6ZXVD8gtPpQ55gr81wB1ca
ao/WlYK4RRlNMy06bigqOBylpgAHat58mAUufyl65z4GiMqrov/3D6UIFjqA6374
1W8FdKbMu8N/EWmsrPj383uQPuUHjX62Gclm+B+9G6PWJvM6+S7h5NvLFMSBw//6
g7pFIvl8FmzGaIzsfuWMwRt00C1a5ADvcgw8lExXFbB35ideoweRzG5Z4vJA3c0A
L5vg+HxfGABNpX2Hb+JMeQJCc0+23gRab5T/rCrRQcL2ng3h9Za5na4Ah3q7KUnF
+dMNY8NXZBXeCOC1BFPLwXcQx2NB2TBmjAFSZ69iiyybctgHfCT0/rNL8zuL1nMh
CmfDjAeIEI2X0HoUsOxSmqTXCT9N8Z2KGKEHR1cSQGi3OLAJiYH244Vm4b+3t48l
Qq6NsHuhji5amL5/waQWaWAnvLhqd0br1AQMMnsbSy9yKGBlWPd6rF4X+ayPANBL
gvinVOtQ9a4Pw3osHIOd6mNfJDSXnGYrN4RrWnEpZe/ImORoG1upe+5xY6l/TOXZ
kBwlO8B1xqq5HQcqOTHNpo4UMWZTY0wpNCQ4x5iOr+ccMf2YTrcrJlABQ7YLm0tq
cUDRrl9s0sJ1DdKskg2NRpb1wPp8AA59Wm5TzkPgE7fbTFvM23zMgXy7r9IzW7UW
Y+99qKrL7NKwvzzHkrp5wAgV+2XFHtZleYDqQlQJdy6mqtBFuzfXafEA2y+ClxrW
Y3jm5t9VwMcLcgw1wW+1cxvcIetLIp/R9rIENR6BJlQeWiKNwYt8jh6Dquuoj1ru
1uqx1BQod+Z/yxUH8TkwOM9ZLSwJRaxMrD+IgWpxR3Hh9qrNfo1oVLqN/5X/XV0p
0DMkzpZy62fi3PQciYtvi772I6P01tJ+EAWx3Rn4scuyDrKziImKkVpLLDWfKVf4
W6TfZGE0yXDtvJFS+MZ+yHKpBUApYnHMV+ltsH57Fgwr6r7d46bCAKTd2nZwz2Aw
wO+RlQgnrvJZF+apSq/DiWU7KLBaO8LXg0n0i85Hj3JsyisK1NQiiOtc0xK8wjtd
CIKdr37NhW/Zk/5/gAV5X7ZTJ2K9t/XHhd+hEOjV1CkT21+m9DkHSoc3PoRGZBIz
CeVWMoOvRayPvdT7tR13RfWFEpZAPovFB+2VDSpcLbtdRfSdTEH1XClgdczSI7Dz
NiiAOob97R3Ou4w6jmJpYtZ6O7r7gBNM04gXIBmFAkNyGa3B4xLYAj9CDycF47pE
nh1I+VXLqZr1IPx+3aMkqkostXA0PIgZZRyW2ID6U3nDbgq2A3uHkkrZzB/isfHO
Bmkwth6KU7YkkeExSReKtIUqoQBnPV+3QU40ySp0JGwESwY0onzvNFd0hO7R6atn
0OdyUWdIpsaRu8a5q9qRHysCriPyzX2tHV+nb/c/rMfZYGX4+B/0zmUhVnSxqQPh
CCAvWXDP/Bvqg3zCuCv/uauO/Gp7uHI4xkJpTXoN42Aw6Hfo/8rqbP3n3C4x5EJX
YVV1SufPpmjIk159pa0dwS8OFoStLllsctW3NpEhyQwdUDc5dQ+xNhPjBBpSuUC7
taUkarQELALOc9gzW3vb4Gx9lhT9hHTTdizjGOYaZ+q83VV+1W3C8eJSxzu3q9Bu
+Jb05AzfVW/1p/mNm3stMOBIXYlxalxSAIwnv9qcoPhuXwsF3/ByF1Mh5Z6x+IAF
lY7oJfMWm3veqgPZbG9N2Zo8WkqUV3nhdGCRlo5NNu+NcN4GzuCZTUjHB1VGKOqv
PrarkMesaViWUO9Rzr0BIocUOxv1G4BuUh9kNpp/evrJDfS1whMyIQHpH6zXp1TY
IWMiX1+v2NlHDwz2+kfDCqfPW5kGGqOF5bsBraWw5XLiQW7NC1nr0u043dv9YrFv
+nvD0H/vpXw9kj4IVgbfQnyqa8ErtBIozxjqyzpv51JUscU23j7PMo1dqcCvV1xw
EgCMS/4YDa0M6N4vkfvvKNnkI9yyJpY4XYrvPdxZGAYCC4wz54MbE08TkWkd0mI+
YgpHU4eJntD9GtNB/Qj0b5Ln9NpO1JSRkU6i+W/T/Qq5XEPUnTL8EZJI2LHKS27M
DbI8sd1o8Na1S8WHiXGXVOmIftYVZugHrTg725evVI5IGsztcjvgkDOQ/0Zr9520
DM6rSoCxVmmAYbUfWRmjmBQZ4iBThCbZep5Gc5SJKBBXenIe6VoWFrodOrSS6hFX
iN0GG5dr0y781fr6nrTVqxyw6adebj6s1rPtUUz5OLq4LqWT8HCcSev7x7LNJMsF
qexH3rqDBbRHpI0ddixwSJdnBAxLKJSY2+vdzxWuOz6rcdJasxWJ7tE2fMGx4rlt
T9T3G8bA1o9ms2sEVO/bNkL1cRJq4ipAMjBaqO/XrIvT6usjnQdVhjE3C3S32Oq/
xq7fgfyJAsWTYB73jSIw73byydMpLxVoZDi8XjD3gESCgv7h3mMQlI6jpxAhYS/x
/ralVGt5m5870uGcUjiA5q2Ay0Ep9QxX2+IuYScoexkD/3BQVqJgpKOzR96ydaZi
J0QqXT2XZqFr1HlSpkS2GpgBsqBcFRlFu5N0Wi31wRdw5/1ANfFvoCvq+Jj5+HRw
vrnIYQ3kxrtKGiHAMWcNib+p3nhRFMuKJJo+aNVezG8Zn6lo3c/tRxgglwt52C6q
8n1qfdcAYkGAiefR79+rF3bW3dZxw7zCNKD4Ai5WgbRpC2G6tHNPGF2gpYGZmRDb
cVHlDF79HCmdMcg24M1SD5r+IcwzvLIoOenxaekSV3BhqnFnuKx3ilPT0ErQVns/
HwkGG5Dm2V16pyXOJDS+xn3DB1tB3cXGWUTv/MRCn7nklfYOjJ61+dISjh6/yeX7
ZINvzlWQLvvgyE5f/QJTFqgYqphcEJ5Ut3tpQbAUHBBACjZgUu/g7alDsIhyMJCg
TVpu9NCiVYm07Nsj4z8Ow3Dgl0vQAr36fTOsHTQFBNEX5+emc9DDLD9TdOCCzOPH
hYVSlSGhsZfPcoAM7uhybtdC3YT5ORUUOfQDNkbP3RjPJx7p1OqN8W5sDwUlyk+C
VksrozjYwlQe4DKH9+z0fPn5/jf8ZJBXP4qOmKD7RPLd2lTqy2FQEaj/h4GMdvCn
aa2XDu3wCmhQNDm9dHRX6my04ZaM7VMYUnwaJTP/Xgum7jSm/UPqEOUlJHONdxGt
NmkVXPwZ33SB3dJiFnyAts8H7a7tJA71kuXTKlJbfHSg3EZk658NwRc2ufooTyKK
qMlIvMyLVh/TAHLNlT/V1ryr43/KvfhCx2ir4rcTXDk3yMyYCN3n5L452aCvAnPZ
J1MtJtbi15fvsopg9eEDG1eooFuhMJPYpnX7kDbhN1wBQ16ndTc9xQX819VAEhV3
chAoTF5GW93+DnG9sk92Ce1mH6dG79yUc8xdp2T1REuJwYNy3tUru0+ldea0yR6F
/08JdRI/PA5VoYSh8X8bQBsKCGt89JqUudWlp6qh6pZZJlSxyn6LwYBXwx5RCVAn
1TcsK04iGdvbQGews0/btE8kk8jsfnhKocSoTakmyqcPoQlJfS1bE6B0nGH5awO4
HjMCu/7MEdBXKxj7z571oH2SiitZpZrZFBQomkMxWZxC8MZgUdNlyEaiWVnRZk7r
dxec4bpcZ92USgXNgZW8HMRMoxR2KuPIA6hY3LFd5WMWR9sOAand6mHGRLFAxURM
uMcVGquxDhZbuBk7P+AStibXHBCjQQg3uD3lupp8bQ+g3/wBKVek26DV5Bfxd9Qi
R+E2ol6XdqlJ3lU56ufDQ+N/G8OPaQSm1YxYUOHzKe+AHd8Hq5W18myuhKH7BUG+
B60UyzYJJMTa2gKQ/gPXwBN8i9Fkq9nfFixnOJ6dkyzetHmA50/kdexeVMcS26Zt
dkn1WuZOEQCcz44Je7gmqnbc3grlECChewZVa3QyakuGUvRNiLgOX8viUGx5bfuN
461Rz0m0aiablt5nN4I9kJ4ZG7BiFe1XRRwBhWxlmONSHkAAMZpCCNdD78xehGTl
uv6qMAGk3CpRVbly/d8pcAku2lAAUIKwUN4+LUHmaScwUKOoEmSB0Y2XOk261YMP
VeUCFKtaxfxI5ZTkovhSwhEBfno0rXIRfoG+CbUySubfJURRTXAY3bDRvjOQhSU5
TMEqyIEPaa54pXYPKQGSNRTaVwZ17IK6iJJ9Gdyx3Xc8W7Rr1ZchadAysu/vxVkF
kpqJ5Ixk7hNJG7+iMTZueBWOXizAUHWifx95ZljbCxKtSSp9onAX3Xo3xu3u+Vt+
0fAnxaq8NdSC0haSmItwaocXXhxsiwHBQSn/OkoK8/gm5xZ1Vgt6LohF2OuqFnWB
oU6E5ew+h4dLnCbvmzIm2Wlz3zYzVoeDa7TjyMGt7RhTrx6Zy0D97FyU9HtSjRRS
h4YUxU9YXZpNFAcp5WAoRYsUslG3dE6X+t0F7hbHZrGAc6hFE+V4Car+f/tFp2T5
z51fENRCVhah24kR6Q/BTUx+Vfhm+0gMhEdFiasUhSRR0ERlMk/uiHWhe1GJoxgP
lrzLE+clwHy+aLvCgzwxY+Ad/LOvIeRWiuARvSfZFqqIgZ8NItWmEfpnSt9U1evE
vXe3sK5Ny9+X0pT6N8NMCqIdwkp2+19fqrDkeJPKfR5TbvUt622i/G6NwpTTT7Y4
mTRJnUXLO1usm5dze7dBpqctz+iSze1flws7UTgETSapCHbVWuWO75yqqhyqyHsM
9DFOVvxG+5EmYQeZyIGMopNVDRG7NF+Ipc8wV02PpOJX1r2DGCi8ycdphOywwyzK
UGRQJ22PGpep7l5QaJ3A8oB5gXbEcgzokbnXubNvB/q+CPdTa+LtRdnU4COsA7AN
f+lLamHLxQXlfFb3x2goKq+7ZPFmjcvAOodWBdpLgDwpycFOQ/RP/dN19Ag4LaLQ
Dg3agV3UpVomd9oS4VJjG+rgB+tqhwsiF2q6FzYQc9E+fcCkglo24HrtmGqjDlmh
aHxQZDhYs53oPT8kWjQphHlPL3Yn+pyCgLMuJoLH9WX+yRzydTOjtvtMXgl1xjkF
i8oiHEUxUnyevFeIrmhXISkhpJpcCA7s5fB7UZLtzBVyyzDoYQOw9yZnXqJdpQOp
6hoG4ENSq8475gW1wG8aUDQSRteZqbvgqp5em5L6e6qTlKlJDqQp6+b9qbP1mpcM
lN/7na/PdptxUZpZRx8B3jbmqWUsBbIwhgBn5UR3DAHnCQigKQVxy+GtM99x8Zc3
8WvYvJv3TEQwq6xczbooSIVc8iOzBh94EWyJahpz2n0O+d52xBiOM/eQe4ucP63W
z9GuWc1aI4oT7tCop0gOoMpqgyROoGvVKmR33Kgv1CkCW2ffOZ5nLgpIxgwqWrGk
Aauv7Yk1CCfTjfzpfuIJS5V4WZvk/xesNILY6TgOzhmONYaDJA7NiEVaAkMuNyxR
YtikYTnbBKMfccwa4gopSQPDUi55zqiR5DsCDpvcMfahBnrgUB8k6ZghLsn4fQoP
1eTVNYY8xeeyS6tACWqsnvb4j41j9BMuyhET5TJsfa2Dc1WshHZ5z5qf/H78DoXE
PTnmFVnxXoEp7HjztnT2UV3ACgx6lC2P5JI5MtBPU/dUaRl9PQPtXo3BlhBBw1nV
Lqc90XcCfisDaQvUkOFMejqQ2+/fSZeHesDVNBw0sjbMHJEK2FojLoJTT+4nmU29
VRa9OEeN1vyzw5a4avTcLxA4OAtGGXKcZ+utKnXoW6SptiDD7GOOQjGxSAJeU9Yk
bVQmkfKHO23LiS0gjR1eg1tzAkmdeNuIbd3yNYf9p9eDtPxRaSJWCdaWXjjrQOfe
gQMcAviQejD+WyzJJXgb7YP/i0UraPiQDwAAWa/B3dLm817DFj1UkCh3hXFKwdBR
6ns0BNXb+9PKxPW1MeVfTzesHF1GZq30f1hsAlyRQnp0h8x67PInIseUcB9l5eAI
hpVoVvhz+JX5w5bjGnKlCO7cg6CfR/lLB63XaYBIMlRJ8q33ocZ+91ROFr95QPqw
luy0xvU0IAktQhsk3qumLQZrgjfT8rqYlFw25FnEvVabYCgcr8AL87KhFMRcfJVS
jRuzZEu0eW6kVySEMrYqxAJ3NsGSOSGv3c+LaI+LOvQuWdUWVfa2/5jtQSh9Ql4G
JkHdyew+HA4PLwrTpVHyWJYXtM4sBubUYLze0SqzK6P/cBXXPV7l8/SfqvNLgSTl
qhoflZ8ALpTBCugkLZqoAEPzGco8MsUmKqGSoeE5kqm04hpQw285sw0fIYAVeG0k
Gdq/vzj9TGqG1HC13WDHl8NSw2TePfzSiE7fL6URrmNk4RNgIgu14o6oTzwAGb7t
LUM+QC1bxrbeg3fvq/6C7b4pCJTCUnZYS2uO8hARNPuJJKjL8WUs2mB+AeDV2FSg
krtbjA894T91tGGOudSQ88+/OxX7FaOxgvHk25iDAgYPnGCpJj2Dq5+Gbpkp2zl3
29FiztuWlE1OYodj0n/vW+gyDOfeY+UZylzZg5+EI1NLQ06fi9Kwx9n2VkH6R0m/
WUnVjPRetjFlPQMnVf+xXJNqIL3HsBaYKhf/ilwFc1avMxqvISOVPwjeb8THZT0h
bGWdRzlqIcjxwAOfrZvwYNq0KHQw7zC3CqESK433Sni+Cy/nvoODxPBNfztSMdoV
sQBvoTHmhadiZ4bmESSkbyuVBlHHUnhVNyw5Ed6RTnf+IchGzZXlumS6j7Q5d2eF
BVRLRK9mkVAuy13LGA6HF3VGd40N4gtpCU1sqkHAtyUjOuIPXjqf1iQAht+UvsLY
DqWL0ERB3tf3e7qgHgZUVI4kQkNEYKaY3E3o3VaAVSndpKvt2eTp/96hVgOWrP6l
T9DLdsx5/ZrTFFpk0aRmnwDUfBxmzKY1zLHIDgiIBrDaw8+3NGq2Hn0b+LP3l+i6
Yq3D/B6uhSvs21nh4bjMM8AE0cNDecwOnPmO835wag5Npr1AvWFoojgs3KkbykXX
nj05ruJ1RcxfBx3MS9Yf1im9Ff3/1rbUEkgshZZUIG7RJrJzndCOU9qNrq2E6QN7
hI/55tDRyyaWRdTcSQjJcvoya0scV5x8gN3g/Cei29odWNJDL/C+na0saVysxUmi
OVbIluMo6JoTh+WDjHU3qyVRODUns4q2NhILE+SUjZhgH8sDUPI/cay2P7jBIo68
EXsL3rcMDwfaN5In1/kHMD19vUiPlPAWm6LWXX+H/8ZTjWPjpqFBDec1fzeuY8yz
LnSWs4mr/Qj8VCuNsbn11oZ7ZHikO0UmitqH081qS0f0FTejAhz6adaJzX0VdeZj
PbB7mTVoGnk1Wsa4cmYMCj5GwDi2O2PeQxQr4AZjo4Sy/INe2+jOuPqrEJemaF0M
2P1SY5ttE1txHUqmCH1nFh2P1vlEVykGxXsULem4Ko61Zx3zGbmLStUvxFmzMU9v
zmn2gTFRWdw2KSSQwfUMXb13Y8mO+aolaaT8aNkrbh6onJMbNuJ+srp6Mnw07yms
cXR7Rur1bzSxgFrhKiE4pSBiGnyHCb90WMHv+LdCJaxN/KMrD4dbATQBy/MLd+NE
AZoGwk++r8U+3WuwdGlJTuRsg9MKwurXjKi3vqP3t+icdNhIihfXX9+dDT07fZ14
nAhll+Jf2romLkLgZfujXfhVyfKLxhQnDVzSi5D/GJoMciNCAePDHJQqmKzGjzLI
x6LX7JrTFmD7iKf18rC55RBGu8EX5PvrADYZSmZVh2O+Hff+Hwnj957GghlrN5NY
+AksCftzI2AGNbI8fP9KBC2mJrg1nDa8ekxkwoIQHKcsM1rI2WXUmxgHGh/UIBUI
6NfOApShuwOb2e3jkyJeDUqFHJBlGYxPUOd3sz62h7HNpRkBKsKeC/pX3Fr0dbDM
RspxxV44ptgGnTzETNHZkP7qm1ekKfmfMJ15Qgp953ZgOKHNSh2/VNQKYfkE6R64
2KPWDPicnaaqSng+jFYo5XzVL5Adc9bDl+fN9D+OJXtAkLeAecKSG8yDB1qA3kjs
WVvNnm0XNpw2yecOAL/8cF/f9uB4UYueKJOXS2CRRVm6rPdZR/CC1dy0WQ+nNTZ/
VLH+4tLbcSmubSr84fI1xIFkIXuadTUez8dTjGswmhcuNLODZ4C0nfTMxzO5bOjj
0ZMi3istHNYjkt2MU9yU2/Hqrvx2tRWzYNMkzLO3LqoU/UDameLY50gVg6FKAPJr
tUVyBRBG/eZaZoBkySOZ2YNKJ8z2zyjlhULYU+5jUbY22lfMqL0bGETS4kPqal8t
/2qeN0QlfEG1J3XSjNHzKqourHjdobGfdCfd9WQIDU8argbLI4wylGHINSrxyW7/
9cfliJPWq8vZFle3KSlTzty/UWjBwAWEhu88P4aICi8LHqkEnvDLno8DtTW3L8k7
34NPVR1grtrp6zL+i9vRy2tadrIVT8IY4olBQVJwPs7Zh8sNo5+QL7PWShRQln0R
fVAxB+bcXjEPIpXD0fEk4DQm2Ycy+2f9Rsel17OCP+JLYBMHXK7TI8/cFInUEjE0
miXxT6epeLiaT/Rc6gZQ3fxEZkA/c5wKKLv0hViboutF5CacH3S+fIm0S9Iba/Tj
vOzo62e1aD28DtnC2fWgULw4DUCSEuGkEKUdKx0GUeQc8eZVPMWhCCb5Gtw73s0N
2NtGDzz2U2vhjz3Vh12mvwQdazQxLaT5WnvRPbi8VBKdzJB9CpqDxPZzPcUNzT6s
wL58mNsGD8ulZgHQ2neomKEihnA13nemTscJeu7QE/RxFy0/zJRskWMr7DJijYlS
qj7akZ/lQElmzhPofvqn4B2inbBkRwCwgGEnqtDuXiprig+cyiNRNvljMqL81SF9
le2fdXeauRwi1HeJXcKy/KExPE1Hky39/MWpYL2Wej3O3KVc2x9WoJKqAvTGLqoM
LcksmsdfFksxMkMvQ5bL0mWqXfDab2fhJscDtfRPMnm9E28sjysghCHqPD8CATYB
g2KwXqiceLr44shWSsbcFbGK8Q8o2Gm4v5JBK8RPxfAbrqgsf5D5+43dpr3SfKWP
PfrX6lidhP4hiK8xiKocfMSgt79I846Zapy6RdmMxzIT3VU80+6+vdaK8y1AEV+4
ADwidTjKKd0I9ccSU4W/M4t0oo2QNwpduxfuLPBgQ6mUziT52Hueh+9Y8iTZKwlv
OK6/kcub1vBlFCsJr2W6hIgZVQagKp+/Nu5dPngVJ9uT90h89h7gL0k/xPSl5R25
zl9FJFBc3WgqPFBqCwmdUTFEDCt4VHB/HHDLq/EpmyrUZMt+JyuxZoOUAGj0i417
w9ThHsT6vAwn+8WI/FfMZpmKNFNhOKxl1/ObvwtqBi7SVs4IWG/J7yGbDdK6gt5u
YgIAXnZ6A6ERmf2VrHH7JNsrpLRrAvDX4yKhZTZicCCan+xYR1j9oTV6U6L54+S4
eCpN4RcOBFi/XMKcnHpZD5wdW1v1xtaiP1+0YicguoH5wEREAw58DH+ottddp04E
+K7UQN5izI2QW01984k7Da/kY1x/PYshry0ghZmMPuVbQY239kyZhVE5xaSlY4aQ
5GQBFIL2cWNMcY4ORGtBDto4/t1fTPfFYjMYiDbsAVU49L/TtOTLZay10dtIZSrU
7JqCTe+hNQcHY6QTScXJRmgXHgYm34FKY+RttxhXN/YeK6xNhOVsOAkoQxKZEvTx
MO16F2hCDHJkUD4ZTyRcISvRxx9qfc1XiiCqFeo2csnMwNFsuau5OxfjxP0z+J/U
k2a/syTJG0qWdpqRGmzaNEczVDCNH5PKWu9HmvnslqEtF3pOeZNWAFCIwJVHBfY1
k5q4Njvnz8UdgQM/+TZE6mnZNp0WWgHdvh5I3ndCmZZRzFwIajHtk/E97aR2musy
C/CrniGzcgSsRGLY+Ep/Smj5K+rrefbDKamfQ+h9pP/eCJBF7BsANxrlABNOY/o2
7HAOihHlGMSOyYe3rKNA+1ZF9KJlRCOGO0goh37FR9cI2OxwQ7vWacLt85+O+0Ho
uF4AQ/gTgRoqSduNZlTECjHLyNpVKZ49MWliHSr4oTdzh+LPVLbkPeevgwNzqRjp
xWJgBnFGeQYy9lz8NxLxOV/Jnup4rcczfwerNzjDkbFxvq1R9xLDTJzLOkqxaiMI
zIqXkMXJZ850iYfGs2Sq2D6M7IyKiqeooIve3ISU16/oFjP4PFXIkqypfLpFQx87
HMUJAY+HD9opC8JMLvhTFzGNldvlB1auvqQlRcJnCLhHlI0mKqyI0NEkiL0WwntK
ieTKuOMiQ/FctkLS4crcygjAKzXhafN7S32wO0RDE4zFPcSfBbQYnVmpvxPAwbb8
BgYp21gXpFLj0g79cBFJp5d2sHfGGY4i5ok12s07ZFJo90w+yfDSYVR59hz9jUE9
GiZ1pzjUa7Mfsy2lt3Z/rYvFEWXytH5S9W2ENzqxOFf0M3rKdhWdt/idNVmkiKiD
UziqG7DqtZs1xdHHIDblM+z0RmvRpStZVWjM72Vf8r2lq+hlVRkH7l2zl+hIqbwS
BxdGMuBZ0kNumkjDsnOQ9gZrjPrCuvxlvYaiCDCRcfvzN29RocZwe8b9kVi+KxbY
GYuNlO33MN2eTGmlnsmBW/iIpz6WzqueoRtVRLeimAWAZ7+zZTuxSkGfvlY2qstM
J/tgiKHIfT+UNvWz5FUpPayZ7iUvBQadTZiJyIeGZsVvsCuGTn32fCvmqSKC7JBn
iAiQK4hxQLPvlnppLQcvwNiGlkrM47VuVXYGpqU1+BhtGHsDeb2+cyRaIJYaURp1
FSXo92DmF/tIy6ztqpjB06lUnklE/Mpd1quYpn/rxGaoK7OYDJpUMmyw4J8OHZCr
baQ5LWEhRbKhAcRhLU6VdR+3L2TevVTyXqWw37hcq1qj/rOFicTwoEcOqF40CEad
vIApIYmbZ3awdvwvWhGZOqnCnD9DMc24CMbZbFKYZ6BgrpYfzNXnYfA5u2QQ9nUP
3yMfuRX38B5y/eO7ZmYGt4AmamP9JL+Jt5Gp8aPA3/gV02dyirt41plCEzSCDpvK
GZSfuJuSsx9iyT+gk6Z3o06qOb/GrQsXCccBPclHq9YHEEnNkusdkcLJHStkBGY4
808ZnkZIKjuytvBllznDXOTRsk1NHrZQX6nqljkCpJHn9+BLQdNCrrMP/+TXC1n1
BFiHHNTHRbACLX0Zx2O60BqCaI+ghKD0jHcC1wEZlIcDCFIC/uYtjnwZe5/KQDJh
JFiXoGTYLzljkbxeDHPckwGrb18PvbkRIBpJMzw3rx3bgZCyFttsyNH+U7ZBogPW
ppwqlFc7speAEUQ+3Qa6uZMj0KVrLbNg7ybxAL5SY1VJh2cl8VynI4tXgcw33nww
idu37Onf5PqP9qjERfgtK8vnf1cRDLf8fKwZpXeN6tl7VI/0kBwUQsvxiPaqNWGn
JlCDfN70LT+Zx08gNEmPtbH7ml5FdaBxEtqzpgWl3TuDyHq7jGKzeb6KhCS9jCvw
welYNB9ozh7gjVQPotnIAB3EXpfCeYbrOfvX4L6WU+gIFU9h5bLzcMaGf57YnX2C
gRempbZ+LI9eeRthJ0eYPEvQRy8tUXnF19Q4R+Sj+Ts86yUeMMyQEa/hjzwkowzI
rQpGWmNOPzwmsppIlyp56QGEH+zAYJKWN7bIF2J8bUndJGx5+XDuKsWUDp13J0+m
vKnuWOtXgzSt6tMWg6vflBZT2PYjfl8hFIGHh+TkQl5qdaOHd/YB1M4Jhzgc9NCq
RArKbyxmrGj80z6HDJZmAm7twad4SXj/aMCb3S9LTYbmoXAXy4ADIJ/UYvTAih2b
5zYy9zuKoxljx738wntR+qH+g6gkoQJe++ECzH9+Oh3iO2gv7d+JXbpSPqIjPIz6
Qel6A/hi1rnQfTaLz1DLnujhiEYWzIjYP5PJ/f8Kj3jExFUI+2JNlyEz3OmLFHyU
KX0rbCWJ5r40EFKEJ7G1qTjCjBmjXzSsGFAUlWPSfK4dK1l1/ONzHzxpFNwkkobi
4LZW8IXbNjwrTpfBzIxI6ti5F+ON3qXIzSSiD0oLtZ699UDcqY1DXXnEGR+jxufK
UWoYCCDqLopqOC/QbXvOrW5nLcs1vXxUYYAF8DCDYa4KcplMPlGup4PUSP6udeaK
e3B1SWkLYEZYyIgoO8On0dqoWEqbyC9vvJhbvZPJlABjM3c8oErpU+uWqPehHGyv
FX+I1/0wOEbxr641tuGTbih8hWGP42ILh3ubu0CQMBNFDakujQCZfG1dPiKxv2AB
w3B3A9hG3PwxCcMH1FlfNq0wMXRfSzLappmUj+aE8cqKtNCiR2FS6Ql39ANGLwEn
l6cY2ACAzBf2czcf+NNVqBlLLX3TKFjqLPYbKFOZotjPN1deGD/tTyq8S7kGTSsh
2rokHYfUc0Lcaxrc2YNl2mL9MFJJbR8aPZpCaYmymXV0vL6D8oOKK0FohQZDEkaU
cy9mqwDWFL32uveQTwRFCqGca7AxzuUsHLscwO9BbbXTZLLKbAHOlYylO1+YILLF
MiFEXhsvFTMI+tqxH885SNqtMhPyWeDyKT3RqjtWM+NQ9YukwCxChgC+TCJfTh+/
W3PLHPuCaEz842wE7xIBudGKZ1eAQShALynT51MUxgiEkER9cpZN9vUIzGmRXBKD
Q0c6+wRqoV72z104sXhfX6WdfBlKlYZjPNtj0qp5O2a6C3gobBlzjZEqSJsH874b
Hmah3oOj7un7AY9FnGyBeVji8u1otrCoPTsLhs3reqEOfOEIJTtgGmvqCuYU/OgD
vt0P/bWgp+SNm14i5uF6Pz7k6rs/bnBH0zhEb00CnMMLAt6dcufUHTssHeJeneL0
X1iwspyzGOqfDa0bKfe4CBMU717fevlxV5t+Cz9vsKR67Vc2NnR6u087qPCfuiFK
G1rQotJ6gt/Wcpnq2pJ8wUSPr8xAlSPw53JRcJRF+2k5SuNyY+MJEyD65XwseIDO
xBH/39p32w04TYcTCFgAxjx1ZMZdBUeUhRHt8ckVW34pNRz+tGiU7wp9oweKkD0T
wKxorZK3Lw7fbIdVn9cfu+zd6RkUY1Kp+qkfPorIToBh0Bi8jyCJKqwtQSIdaqRZ
Qm0sDkZ1zN4fwW1wlmjZ75gmfw9COTgFzsQMPNcYvW+nMSUiEdiJ2ggOKhLVDyIj
8I5xfjkMCDAapuzF11N02yxS3/z+3KQtynTkz6oTTwoU6a2vaPDQWqf2CybeMj8D
nRVlUufuq3s77U2CKKU+GdUkSR5YIIi0mVFZ6CEExawUf6mQDtrbSTk5PIPeuJlh
M5Objo8DOwpPYTsFDnGZwljyKGAwyh1beACZR6bO19yH6PJkQcoQwtJ0zU1rsLPO
qmhj8U9KHij0a4n44E+rkZSIRcgaDXbNQEL0IN3XkXA21RVKAgStnAPS50ebUuzs
qKFGdYh/stKoJbOpvnPtiKH+q/1m+UubGjkwbUEDg/Ffprp9TopidHVeEiqx02j6
1B4vgNu0xJXYix0iQ7nWUzmwhDUk7RK2v5pHnN88euAcf21F4Vrvpw+puDWBq1/Q
12fQn91Mf7Kxf2wbYRz63FhwNFDCsCDqJTLhLTpAGYqfosqo67dgBxP1faytPe/i
wSOu1qDa++/uM7Iy1NlxedvXLJu389A6Yog700q4fRanu9DaesjsDYWY4up8k8od
DYavx4Fc3ln350BmnuTncHEUbh3Cp2xj4AzTNV1yYZlvMxv+irvN+fqm5M6//mn7
O43gXyaYOc1VK86VDhVDCgxkz8QFCk2qWWovLs8PIcWXXxBmzLYaf94Z0/eJnyJI
g94OttprpLNj+FMvvjZEB1wuoYGHseX9O7LCTdh7vzsutmxqfXlhaFIfNVnSVm10
isbYFQSIMe4GQuFTMpB+eUBWkFtluUqg2v2bKbtIoy1L0VAVHtwy1JoEaMzRUDOK
hJurcN0072ZTHmfKcnY36YBUQUfs1M0PTMx6Ti2sjQ8j6MNSMzYmKtmL9RPVUMwd
BRdD5klXl0n9RprmDgdF7JP3jkEQ51tjh+h6Yqt05ofRdJITg2dBA5U2JuN6iLyd
8kzzyAs5GCvgyt1Is6kP+KPRyEkuP2VYAcozEdX7j0KUZUekBcP0m4RJCJB+8YoO
FPRA+f5eMjLWBQVS3PZN6/RBz9RdbL6ImHlM/KBXIrPPMSm64KwFS/JKOVG7MP2G
YTk6cowmH9V0w4OaTbS+GPbp0aE/b+L7yOi7PGXgUHmJbdCy4zXFyNApVcjUisES
B9tTrJqp6MEYzkpJ26EQHcSLhi/q4zin1P38jIb+zZrIX+B84ZwlvNXUr3u5CJKK
ZsuCE6LDaSD6rQM/wb59R7RHrpDFDNkyW9rAG1v7+VqiikO0VZosUszDE7BgF+7L
FvasMLkjBu9Nzs09CMcYH8VcIWi/kpoLjweytRr9K3E1K4e2O45TzYXOghPvg4B+
poKSCBQ8lIvHsc/2JYSMsW2oRV+yviACsGkzemij5UuLBOZX01rARO64KO3+58Az
6gYXR1Z4GjhEKYEHw/ewOuVczSuJDYpY6eqPZARa3y1S//Zmh2HkCmEyr7ggBQ+b
/wUT57Kmrx2th5AHgXmPE+GcXge+cWEu7zdCRghgtJ4oHXfDIlIlYuhfzUjXhp6O
4r6gsAc6tFOj6qwY4DM/WnCuqfFSajpdKAwmzhgRKaNg2ebIPMueQlDl8M3L9k45
/xwh4Qvhivdpafw59N4cvOXv6QQbU+E+ArLus516Aq/I526/5/Bo+QRm5jwbAw6v
SAJw6XhFrbO/wOdvAXWo5KnwWNPGzmsglE0yra8dBUo0rx0DxUP5QpWh0cBskXmz
grWrdM651Hilx1x+d31yq3Ds/CToKU2a9gAE/fsrTCqB+ewXutavNcfCG1bp0ok/
tB8wpSFoI90dCU3SXkrlOzSgre3EQ67fCWkSVxvI800E4MWva3XXYZFV3SMp5U1a
sR+zUzmMi+VT4MfJJOGt6rni6JBC5O+p02UCcjIogonQ8Q7XLRtWuYnA4TAkdhfJ
rkRlavU/sye7Cf9IkcVLt12M7fXwzIXef8TwlDyUJKvVctQzvMu1wslnc4exPfaU
HMpZmRJM7jUY8e409E6xSjOL7mWwhlgAyRV+rmEY+h0sHpReNFQ8MZ0qKxF+QiC2
v9BUUXFTVfv/NdnSE/WXyZCmEDJuUB9e8CS2gFr1uWxV7aIPULjmGXGV3sqDBHjd
7L+C9ZVgNxwr4336ymwy/osW1h+T40otPWfIaal68c6Qh5+vVxks7Mq+DZraCF1t
OO52SKpOK9UFKC4xAUBQRrxfjvdVNWqUwYNSTWDCvVKKXJBZWk5wlWoZV8aomHBM
riyJi74p4qA8OK0Y0wXi8WXTCNWQ5wQP1FtHdVtboGvtN8M5q7ecvNoJvuyb/520
mpL0vZYBNoFzrlirwVf4tUomSxT4/w0Gqx+RMpl3du09eZPECZEnuNRqHhsA2gEu
41IWQ4wvsz1/Sa+6kZvj3KiuaOdEJUtS4G8lABhUSUTI3Y/2LwplY7g31cp6kBpc
jmC46M0hVkSjC0+apbeomoJZZ5ahYypchrx2R0j7OLW8K2NIDY+RXWmNM+dngC0i
32BFBT0sH1COev+3lgCRKonU3MZZUgcxeC+v+P/Mg4Ih6wLzLgZJbtJnKyFA9VUN
SRfnm4fxfaWyTgMZDRjkWMWe06Dp5/F6kuj/wW3jJ23hPyXuwpQm55kNggkKZ0ag
M+GZgKu28+kmHn7vWoo14HqefxMWLh/5Y2AQho2TrZSs3E/llIDfr9tz5GkmClCi
vQeqgLLQtTGJHX8B4fgmCnV2gwEudR0DaPt0sScxOMk31WRZIslL2JmVjx6UP0ju
WwFk59k1ONHbIKGKFXCj8bFoDMzIrih6OyT8x0pEOgzUuK8lkUqDCL1x/pcNxuDP
ttPEtG/8342t+GU7zNuUe+9iUah2P7P7DpMCKeg7PCYNCm+X8ezEFThP0ugsPg4p
IUU0udmMZ8toFEk4w/00zY9IXsJBrIsx40Ws2f13i8fgpH5PcbScZ/zEMNx0JjPB
mdHUOQhZu5e9dNoExoD5huQFU4A/hSAfk5NkaoToFRSUNlRvFY+97kGH1gcNvddQ
YG1fnaJp0NTjIxnTGHKCTCndFNY8NgdCoSiRWcjan1Yyi8xemSHkPyv7A3aV3MhL
66LlGCtD0b4rbBVG1WskHReBfQtr93oKvoBm3URXsTYv2GIx6kaxRzDnlg+H0i+b
GMLMC/VrgZQ0R28eP9ammnE5lT7LQGoP53VOzz0xBXce0n3YNa/L82xgVli85/MC
Is+GMHak1Dz0GP6NwSpsoZ255EWyXGoL2CTmloztd57ZM/ryq3fygkSPTqd6u6Us
IQAaEU9sOH1FnsPu+cBV7qP6syRluSy6XSlngw1tPQnna3H1SzEZojb7KAYUod4r
tzmYi9jy8hL3dP2D7+whyhQlGig//xs2eZaAfehBNrCpBcidiJyXyJbpZfylGcu3
6FFAZYkEaR0baqRn8AuSETHsRGMZto/Zf9jPoVotVXBt28c6OQUSAOSOAkn/vp3x
+X6N2OihwrJMNHaGCTUihWV3K+bl4HRuaoG2wwGuUeXZPSmS+kteAVX8dbKWEcVZ
UohcYkA/6BE4wxKxut6qfaC4uWrpS+InuIzBPxnyDA4KqZTZDZ4BoIXGS8Kd4q+4
mB+Clo3f/fl7s4Hk66sq+O6sZXtFHv1k7alKSjJNuB2I+rx5l2OtHlpiLxc0YuUU
46FV3A/Q1EYK1ZrgEaDtX+vdfjpolV4xPF9hABW/IRcjHmgwl/chtzJMvrpIHX9v
1pFm6CfK5gt1jRpdPFfJX227Ml1jDSxBQkW8BNaQtYMOpypM2cwEJfSdicP3UUbQ
6vEzXlaD0CGQbyfFVWQDo/bEletpQ5lkqRgRZsvXoowhuYuT3XBjWd8r4eMGHH9t
VEAk9AMmfgcZon9cdQnQe2EWp0a5uKb34Xgf8lixnEb5YT7a12krHWYEWTdF9+jS
LPr+g95zOpNlVUDP8hJRd5Q4KXq6wLVWKntC4MmoJzkixnJgtOnf8eFXtlE/kQND
yJDyvaccTH7M8CYocq0ikgq5DT9wD2T7isjF4ksjTYgPgPBzkQAyEfv56w2Rdtr+
8tyzXu3Ng0jhI4qOa76g3Ak9PvsdDaz27EAmWXc+I5baG3dVsmDa1kZdq9qzZQ+N
hkZpateO9kYQ9YXMsy/WD2zJbwfzF/l5n20UJgXUn4ned3i0dBTvUQV5DutHGotk
VS7sew5NehPLFF9bLg0/k6pPl1njNtcfIpc0IbPcpzAOE5CC0xgKD5swVY4Y0Nsk
fcfZUfqCd81HadlLyy3fqt8oTjH4zhhFjYL3JoVWIaPqRJjG9Srss32fDFmseWpn
pb/ydHQt8HKbZ9UojoIZk+GWtXLhZt3sk6+1D3tFLWkXgKA7xRAfdlgLU7YJd/Ph
sl5Orrpy//8J6z+MBBVqa20fujEH8yqbDNzHwLeL35Dxj6OYKmT2pRp14RvxEw0I
lfHW8P1F39fliB3CTtFVAWSardOleALfuXscNrnezytWqTBvqKtCtT9yT1EV+cZ/
/K9Mk2wn/AOqoiJGf2xr0nMozmTkO2AWrEEgBXbyjlWM46LpXc1mLTL7+RSTqk/K
5av6cfuwZBGuaGOkesTTfqcsOcvzzm3ozsaGrOYU6rOcBk3XpwcF7ROysObfwJlq
IDXeSwTfXqEhro8jIwJNQ4e8bDBqf13JUjuEXIlWvJsy58ncrc9TRtnmjczfEFFr
3OylrR4+JehjsUKNEB4UyYBRe09/rtX9ohje7NTRiSSzCdJnlwoVGVxZiuYO0ah9
Maxalhj8pG+eY17j3tEw1gDcQsdwFZOhc2Me89VxqNT/flDCAl2LHT3SIWz431pX
LjjJQ5vJd7q57gG0YaiuxDESK8p8e3a2tXs7aMBx0dMmnM1k7YmcDmbtqkFCqaoY
1dIJ2QYURrZvoY4thlP467NyzwvtBMUDYE2tMQzA/zFliJ/WMgO34thnON5MLLd2
f36wSJrEWlhUUvpt10bimXLlKH5UWCOPdveBlD0Qo4RbXosxhoPcp3pNw9ARujjC
aT3y/TGiBPiqPhw270CE+qcCJz6ncb/FbeLWEi/uhBstyTorKrxUrXxUIjcFEy2n
mIBBx71HpnRGYEMgGGGqv0fbud546lbmcM4wZGnCECEK87kA8FQ2IzcAg7N831xJ
UoY/QlJbqlTM5QeW1Gx6lD41NkILnmT2cPDNUawuXCrGIPNptZJayJXM1mWgKukR
xMfdfym41mIMEFkXSXcLbJ3K90LEysHtSJuu1kqOCM7+VI/MlxgEBIlYLG9xVJbm
RCUee494ZrqEJNtYBJSu+rFH7nDO2r9PY1YC567y6lOgm9iqR30gBQrCcO80xEWG
T1fIU1mUSIvNN2B8vaeg/eOQNHS7xv8kwMLTtUws065t9AjHCvW8S7MoX2tcyjbF
yeeFyo/1c2RaYf6iawKmAEHbV4sM7phjLpvPBhE9Voh27bCHbF0idauQ0EJcLXHk
WC7yU+sG0qoHy+0fjUL2yZ9LY5erXhYkCbu0qhdqtb6z7raxnMDJWL4BNOSPaM9Z
oCyg4QstBwfzenV6gihygQPD89B03Iua/P1YkYZIrZCRqWp316KSALcvfyhI34ZY
RL2lkq9k9M0SUouzqHJyK9cJNZeWCnUj4Ro3mJwxbFym/ERYf2T2gnyiHZ8Li1co
y+Yt/Sh9yjy+RmpBgEl3acFnEg7S6ccmj12DSh4P8y9IRqLe1eXwQpHi9WJvreHO
xq/FMJpbxGtRI9W4fMl3OMU8UQ2H9h3L2bmIAH/GyKawluTvrqsdgm+P3O2JMZur
ghlxqKg7KQOHL4r/0+r8vjQU/1VEVgmhnUcqRcET0S+n5cuL+LFsYdcKheP13ELX
EeVcUzVYfIPTX2P6fQwcpucSlv8Hue17Kkn6oSVFibtBFVflQIepYb4073q3d7pF
a26Jc6c62oqJJFeErJo1Wlo6MsVGCX4wSjnwHNartOUFqOKa//+J3aI1MkPKS+sd
KJCOm9HWZpRB3SHf7QitFBl3pLTDYzIxDcU8DOcniGHD0EcLJ6Wf+/a1eCPfrOfl
S+0S3AbYctZ8qRHw1tGEqqgROXJRClF+4B63gcSsOsmi0+v6ty+x9Ce/cNnmQ6fK
STuJlQAK4YAX+lzNWu2XdVUdh6mwwqyyDO8uznPUSxpLM5XAyp7xQlV3a9W9LX/h
RYKIKIaJqs3hqVygfH1P7vk8a+kwqBp6JbkJwkMGXImho25Tz80+o766LN9dspdJ
XWC4SxUojIS0S8Smz0Gfkp17qD2sr05MdYJuFmfih7s+nRGFkAZV09LCKCaSZAeC
5a1yVAUlmjVQBskMf6u4+OgspXVjX5YSV9zdFrE4sQdpPMFk2aKTFchnWXTFVY/X
D4l32INg4Q9TL/AT+WWKlurDQ5tSBqrS3MRMzxwQP0hq+AYvBuDQQgm9PHLcKRAl
lCpaY44GFh+GlCA7NOwewa2g72BCxhAzIC9gnOqZxLEO0QkrZxC2ztRUj1Hy9kh5
NeEI683nfcUa4CAXl24AZXgwnU7yHmlUkaw83aPFapYDysM3xy61NhrGhaDoEMR2
t8qVpVmKv7JnUta0UwiB/zRy5vp6fe5rQzGad5PDe8tQM1y60wWl6cfdTlBUY26E
iuC7U7uLwx/HajsHiCc3CiRQJpTy6fIPSS0gILFlN1R7msVI/8ExcqnwTYUsnS/k
kpl9/l++83ApQiVoRdjkSMmqTkjlw+Zvux2qbfx9fISoo5ybYYEweIgIYI8/grEp
VC6MeiOLqONzLdnQh6aHjp2m9wroHTrA9jOaN7rP6JuU3s7pSyWx0VUA7M7d/2WL
ME9SF1sIGXNoLAtOw875IyUF97+BEK1LbUcUwZRUWRoYjV7xWD4JTfLzeBadJg09
ixQ7teb2OaeAXZrS1ZfgpJoc6BNpjCGReG7CbuCk60slYmkO8aeNR37CrSYeJCmK
KBRQQ+dXOPnjNjMCYWYLfx4bA+VvnIXcQCcb4qA+635MUAV0f6sS9SqZ20al2ef4
AwbvpJEUASexKRKQKFfpU2h7eAYsxnvXXxnwhe/9ANJZqwbD8yoDcg5WCddGNsgs
WZiz8JoT9jS++uznlxJY76xvXGZTYXLmUfORwj6hmHnfqyOC659k/m7WpPW/8HXx
TaFdzJ10wSm5wORb43SLFJwpHbU1JCcPHeBN5TG0kuaeuoUndddW8PrBG8CLDXcR
mOXF9grs93XbX3lLkDwFYCr3nDw1djJqMYMo3M1977hunj64TZg/6KNYIBAIByi7
ZEtY9QBbnzIZOySVPsEucbk7yec0tncMrp6Bwl1ZlgoTtxrkxKcp0630CD9Xka1q
AyZTHg3kMUUHoO3/VAXmUexzgiN94tzyFuDEJbkggbwv8K6+Ey6Dt6sqvyterc4E
s/x/pQUz9jI6ZGOlmn2yGNr6Gtacweb61/EhzY7OnbNBmDh2n+TbCa0lHXGv+RoT
sqGx55GpkltRzEOaVOxFFZmjjBEhgzapZYm7PPlbE9O+ta11wlpUECzhyMepEs3F
zKS1UIi1UyAfjwz95gzqMwBt27U6akZ3sp8951H5W+ZJqvMiLJ1s+mWFxLWi2ibq
i1JP0aounuWPCLh4bCgXdHl0yFh5n6Cbh68QgmfWFXDC8aKWPdegfLhIrtlY0r2F
aUk/xrhCQERZGaypLpIJYFiCfOM/DwZUw+dqstRoHDhf+Uxo+Oo2dFuJFWPW9ovx
3v5l5bhdeSb+1jGUia1go1VZzz+ghOaB1ju35xGGAxleQO5ghVPFVURTc9pH+Z4B
WljvXwFz+guaz3+zYB1rCPouIcpTox/QBZIaJAT+DQCYxGgkn8+Q5JNWqY8ENjx8
QZQdJiE6/viNbqu4hzb55xUuJvXniGSCsnT8YJlU37DT5bddLbOzE7uD7XU7Vn5Z
lRN6GsOQOpmdypzBywniJopY9938ygUzxcI4p/lwCfnSOH8Lb027oiRNK2AyHUrA
BtMYNOdE5l3sDHUJ4eH85Xsgj+bOC4pySymKlg0Br69P82/RKK661ERek9Tt/LEn
hdh0QoP2RvDbFyhYUks0v+GTDkki/MWa5vpFFvhiXu+GaF63LjPswPRk8o3XUd3j
hEMvgE5oIFiJELsCptHbtZ96q68AqZX2XT0vWqnkZrRs35pbjFyMvKTuKwJQ5/WB
6u0GZKAwDWD9TbTkw/fKNQjgNNy80hg6Fair/5VsWsmYiJ80hxcjVgIBfmAoLxAf
6qNs0iaw7rFBnINWVHZPzIt+GNqqEgl8LvCjTLgx9ZTuiF0a3PpbWl4HnbntP7ju
RRMy2adCWpho8G+FmrZfXoZ19xCD2W4KNVueHWSUjTZlBdmUtdwRnXJld6N9T9dk
3JODrUO9lgmt6fgoZCxn4g1Md0ViZiaWUdS3RpsYCeO+h2Ay3KUia2ZeNeSt8NE6
jv1TJ07NC+HjIcaQPkVBTQjS7c75xJeEW7MqtGiqyiSMWuTzLHiE2tjsl/JMeACJ
TbGOlS8NuohiyN7HCvGZ0l3K7SjuywmBbr6DNsXqp67bY3xdz2UnPxGumQf0WQ/g
5VMDFS2iU2UqxKUfriNLprL4cJfkHchHCk59QEMTNdNhTYxhql0VW5W9MIq9c6p7
jlZhobgQ5DeJ2se5QuSV9rHJEJEi/4dWCcjgF4xl7qHcNVlt+wvExArjIzHKa/fe
E1CYX2gITxuiw+j/Q3Ztgo3qT4ozoivtslVcrit0SP6KQZiYvUUyDtjuodaMulUP
W8c9t2Ulvp47stKR4IJGZJ/ap7+bwV0j07xSeLukowxa+ZACXDtktZL217K5TKOj
2ueE2CHRpg/AbZZGLeRFN6cXzvzGlPpzWJDnoL+fff75kjn2CPKAxdKzKJcCq8n4
DIBzS/SoFS5iPXMoRaOAXWI/ZDXNmJSDffMBhcq1u0a4bSiR6hszOXb5ZDlfrQtI
p+s3dmILC9bp+JonVhv69i2Jx01WReVST7IquKmaJNBHW65EGtH5/L7vKgviLzoh
DC5UJD8gccTeZQg9gEW0FJhKP1uZ5zSJ6C3/6e4k261XBiO0HOKWXoiNKLTIqsgr
bj/I7aVIC7DyHFBIE3l9OLiVKKhWuqZ+sL3kI1APgoKGw0LWGxwUJr4mlFX+bFSG
tUsdDorVkxBdlKAWs48Od1gn/AMakau+5GjDkmrIDl6eb4nWCtFIs+xBszjI9xLW
m6v9n8n6BfeYyKWZ45tH9dpByI9rZWT3NhqX+i0zPwTK4dQtcSNQRNSmPIwdipP5
77C1jxIlfIzs14/eul5E22eNO/+lYOmHHxjW3sfrNS7HswrGuHTB8MaOWJskhTP/
B12U2F0GN7YArSN5+KoV2ggoz5U2vMZF0GregFHSWnr0+Rvsxp22BQg3g5ji8Mpj
x0p0+/1V607KK/oSd0MVzTLQArQrSvtRyyQXaiq14H88gXfL04uRuqu1HKlwhYYz
TT39FcdyoHhaRa6bGax6s/CWromTOA84w/jAbs3oUPjF5XWj2V/u8MZI3vER5Hod
ceJQ1Y1IPQCRg2yPg9Lx2P1TGgdSsLPJBWCH4PutTaAfq0YQfJqhZ35g1JBFCmrd
2TvpYYa5iPbOpBukvMdpADjB8mwb9D0MRQ14ZiDYxD9g3ynhAjZFMijhV5XU+MH5
YIMXXd9tm+bAnGiMeCGi62kVrSerl1iFYBK8tFWmkRPJf6FOnU9GujS5VK2eSYeR
v1Dd8lAq3zwazN26IKAIx6K11ysvTnITKW0wCYqi17wVghrxu3z8abHME/YEcbEY
zC9YNssqormxpk5hj9AEpr7hueDJnHnw8xeMj8dQ8kJA0f2m4HUk0ol5Z13VkTOJ
idr3WefblwRBIA4/J3D7jnf58J3tIEUAJHvORZY8N3J0ua+CFylM1sVZ9Odz6oOG
iEqET0Ba2X+AHB9eHet4uthqDQH9uywIslv1Chl0D2PyuJVFBZC6D2ebB8iw+iGr
gEvN5DgE96b76Kx+/t2CLHUrOCeEyBibZOYgSWdqmWGN3Hy8ki6k41Z4rGhuN2Tp
QMgLCezneiUZmltAs1wVi7NrqduxA0WCHd6oHKzGfPm9JzuKDC+1ZvREu+98WpDy
6crRr7zmZPU3JxTVbEdJuqVer30gyh5sf4kSxmVc3bRFHZApqktitRQo7iidX3xu
9WUAXeCTZd1tQSGmJutoXe3FquWrFWbfSa4qcUQNALveHXpj3VhUWiuileSTPffY
SI9EjeKxcGqBT6TraoItFuzPUm1QE9mEpP9tN6gkmVUA6/b8DQUGx6TodevcYdLe
Wt0UzwkQEULMCD/Z2s6bNj0qNnzPorWK1IR8Z/GPHtFzvSzHfseZQnhQBijxXMjv
axDGEDsOaJqNGsiDHmVn/bGKvNdCLW+Afu2k/jbMbJ5hFRbVw13p/xeKglyaD6/w
3pvrghzgT/o15Fe0yO3DNrWsao3yLbQhL0CwGfRGsvX137dOO7BFaVMEfOLoWIy3
KLl8n1UCan6qQLa3L4VPMfEAFnFDMIZFI3RYgS3EiXyiXcyNnMZqWiieUWD+wO8K
md7Mfpc+JDqW6xqBv+bVmyqe89DKV6G3wGXXvUmpCmUsWja759yRUwF+aS20+nYT
28XRZ5vC1FUiylQqDE/LcamKS+b6ZiMfIWMC61bGcR+KfOrgyZddncS6Q/QmP5hY
0QDT/66sDk4KSWo3+XHMeCVwoB/eX8VZ8jkOoS7rBW0Cs0wQwq9JKiQTILnh/hZy
kYndXSaoAEkQesfvSozKyPWdWvBI2RmH9ECzUGzdJOuSTrgYqVQum+ANOA69VUjC
YkEhEm4h/KmbpVuCVT74MWEpFYwHLERHBsW6SJbRAW1OzlfNP71rIKpj5ty0ARDe
rkksBxzUw9HejRkFNoZX7HczjpJSyalep36E8vvzAZSRFTZU3InaiUpApGP8ZvPY
6VF4Tt4q59t1DyhOLIzg8cmiE2y7NRZ+nY3rafd+bTpPOZSIpGFJJRzvG3O51gTA
6jH0WhdW0yxRf6lE0HySBdvVKchXSRjpDwd0EQqC0wsnBrtQDE1htL7270rivooq
v4kN00+CkZo91BRFVMmOTr03rUhHdeITPy+gODAy2Lws1wXXCq24s1q7ttCkZrSO
WfVBG1s0w1RzcsWd6wO4aB//Tivo5+KWY8YPDZEGChUP51kMVElsMR8HY8ab00PF
F4M0HaCKbCon6EGPSj2GhSe8vSAr0QhpWZdi/wtnyN6OqOB8UjbbuFvC6zJgzm+j
HgqxAvp882Z8w+2BtN4e9vjnJhBk7TwcuUt3khjWU0mQv8S6euKGjEhyXxsM+aUz
4jBhG2x5vAbP+gcYg6QPTX7Yec+JO2QZU0RpcPuudyR9JXyZfUm8rM10xRTDCHIA
IHFqhc/Z1KQs1FTd60JxFfk/q6zMPJ7DnXjgFn4XseL3qBJLQqm02jLQUVSJnR+6
jczSLFaXcxTs1OVfO6fbHnvzHFpPM3sWWciA6B06FaxzeZRE44ZTUZe060s4DL1h
1aM2OM3lOipsfvZyReRVbyS/GOD6HSJTTe1zSumKWMB3SnyEjOMzlDsmj/tu6qbm
YkCBU2JTvIy68cEVP08rA094DncJr1GuqSa5Kbx0/7wQXhHr3mmyfJOkmKgR6D+V
eyexpfTSTrgp4aYLXQYqa1pAHatzoH0KBxo1NQ+SpURR9EKnofsPvVK15MFQNOwj
TKIzV6Roexip0m9Iqq1ztXe2UepexQ6JwN0BrkNfXdxcauEGIJbEQU6evUMKxl2t
Kmyob8zK0SpYB4U+o0QP2laBvGnskkfa13SerKs4zu/6B9R11zsAacTGRnSAGhJ1
OpeiE1QeyBQ7SV/ReHmL10n2WtvbeQxxur58Nr+LrYImSCKqb2Xv11Il1dXDZ5Yn
6sg6ffD16pNr/UoQUQpDf8UCiLhm9VY8RrQqiPZ+SnDY6aeBOATNVZ4fBy4LIHYw
2qzyjicEQZT/XvyQ1QUshLHyqiSLv4CY1Mxe8BARNrheeVK++x4GsqUlLw0+46TF
dJWNRB0CS0R2fZMEzQQteYSgJopTsXNW0nGan9f2DAB0QMo89iRV4IFbolBymeCu
ckJf4DtYcqIUTNQj7o/qlSLmwPq3xBgD6ytnooglDybLh4gPevi56ziWJBmdDUWo
BiYX6qDqMKsNbsPgoMhGycHuJYX7669DUYwYMFZdhgiPDZUh2n+WF6ehYjTBs7Ll
dnZs8QGwmesTUoAB53E1o+CmCoEAKG5LgQPzu8AlpWqJM6CN9r+i3Z6UEJ5tXKQe
QY7+HRcI0z55l7fgtdqSr48dI8cQSGbzcLolqslBFqKF0g1LaDDO37haZreIJhwl
LGwxcR1ht2qj7yyRcg1TBbhIxibPbA6LGmInGWR2bLlD9r1QgbE1/KgxYBvd9WiP
yFqY9IEhEzyjdL2XYyiLIjQYv3AxO6HTMWtOZT2+zlEAizU2vg4npQOiGd8xOk+8
c4zlJakho61dLpiFEEtHsAapI5BJd3xKPEGXi4rLh+EhSlLbRRQ7ZogWNZtCJdyM
xSG+3IMPrn6KgrSAh9Mj3b5doenRqv4sjJK2p6F2g95jY/rdqX8aJXL0n42N4Bd5
VAwGm5OnUcDff4j90nwywu7+3uO+gyd5WMTSz3i7q7P9wmbvCmty9IPXEpAj0ElY
2qXQukpsJw/pppFSehHY8fF6med0+XxUs5ihl/5RXq1dGPQrLrEjUiL+H3Jl2Oku
ZzCnCG+b13AzLIJ2GGrjdeyZjsg/ULZb2fxbXklYPhfb5uK5lAg5lQh8rOvggXy5
WZ9GRuXcog8uqYsMvu9HJILxL4TiAGKh4MEbA/Yu9oGusUqmFMB7OmL+O69dcwlV
VSKoLehouW+a2WnZke4nuPaANmlyqhUlQT5SPSgFOnS0UuZU4AH0AXpRbiRqn4UI
Jq7UI6+4MRTQlk7Mq7I4iRtelQ7aPJuEPBWqVi9wAef8lZ3Pw6wYtK3zH136woj1
dUCHqVcxagO4MRGkxGxLGGuLkXCijPwnhcDbUjkFa20Te8yVUzlUjAtoXGsfAL5h
FJbxMCuiTo71V1hb3paX6MuEtq5jz80PJ/ZwYJutqB/NWdvDv4wdYSckJN2MV27k
RYvFQv2UTVSmkWC8kyfsBE2HsJ0GeBNTyH/M6SnD0uKFvAKwYtWXNOqMpgScJg1e
1c4JKME4x9LmsIEpfchiPIifkJyn55rP4SxRP0ks1JJS18Yab4xx0bocLzcTa7Rk
aY6WI91ZUFaA0LvWzkd9L4Ys1eGAc7ZnycRxyhozktOjqFQ0yytPk+/RdULV7Nf+
HTyYgevKVOuG8nyMA9cFw7vXcdseyHCqcIHNsBkG+AIXjXPXyTcxGAmyNVtg2jfl
MUyUn3XENAQ7khAXv58jGptITsKCayVQQbNZehRVY7SKtxgO7IAri0AhP0safyjO
aKPIKnHgoFdssHT2EcrG9rPilMACwJArmFkoef7cOgMfVG3Hf+ehtQu1oeEV6aUE
6sudVHbXsO2nF55bDNQCEOrR9a6eqa//LGNgkDObU5eml2ZS6WKf4QyqNPEYP8GG
EOoGqkUJ/6J5/Ylp0rzZp9m2HVY66+yzmxdFU1+oYu/oLo2fWuWwH72EA1sstQlX
PFEwL4IUR+OjRAHHYK+IYYmg/+HNiDmkB+VHAYbF4CfK84t4IedymowXuv7q8EmK
Y5SAVi4L+XIqOJ/olrLtDsezEek7swzvSuGoVwcne6b8M82gz+oeiBk1CAovWAtQ
j/iw4hqaFiHkqp5kors26a3Fs3gWKZRuIJKJdC6J1GkYW6Hke51cg8e5ElY5sFfC
pQJTDWrbFpOfnhwE+1ZGi1bTJDXCS/vl6Y1j1Iqo21ZAvFw/t87yM4GqzrPR0gP1
BtQ+OcOciBJdjM02/tNxg9Wgo0M/c1J3Hc23ktiuJ3nVE9ZgwzFGxe7UNLnkDGEX
etbmiAMcwlqX2/U8F+RwF/qiiqHT++Gb0wqrCIjEruAri4ZfYOCLfySl+7tvltpd
WA2n6AxU+X7NhkOiT2CqcH6JV4VevtEByxocP0AjidayYyepN1z2sLnly4508Zke
UUQztuwYjAjClICDZrZeiCItYoOCJPNfFdQk3hGxdJNb/BQj+1KJ6Ge6x9mmFo4s
6mzNLE3tgOECFZeKGSYEfto+wV1j5Y6d5Jsae7AfKebDzV4oIp9bhiNQGXUI297E
KkIwIWg2ThpuFlTyLUxzN68ItI2a2sJ0OzLCkzAkewA202aMAaHbIjnmE78kS6Vk
bH4sGrfsAK4/5jBgDV+hlgqkYnBB6Cql8K8LoaXIA8jTCTRHlwef+L/8t0nGmFAr
rUwQuTqM0sahV5XekBuyM3iakErq4u85OzZBQHtbKICwxU0tkoKMYECzPXnPBTJe
rlH5L86c4QRWNw41HU1Fmiak+/0rzrBxK6puW3d4tfy79I3F6HZT/uJIRzLZWdy0
C2N4S5wv0SWgFip3qIHSdDNf/19ECM2lh3EOnra7hCoe37NfSk0aBdcTAqN+Nk1k
3lYNaG7FVm3uDG+s57qC7QXb5Pt+lhJGj8dLy1DoRjm1ATVmA5ze4EGHnW+66f5n
8uM1F+I1F6XnizATJoCaEct4VR2zW2gTACkTqiyzCEhTHF46gnFYWYBWIqW3IV3e
vzf3yKIWeEWdFgTzkewrB5CeN9n06qrM/h7jz66xtYZpcISakaZMs906sXVeQDLb
UhRZSwIYmg6StRrcFu5qvPwY26piBMf/k3AQut65xzMyiUsLBl5rZxR8wwH3/HBj
BG6V1YZyG3w0tt2ZYO9ovoQ2kYvM0wbtFSLzqo15q27RsPQMELjM1o5wVV7FWtsV
ETmy7l0CqGAxgBPkc7MD9Mqa8zaDg1NczRlTFJXT56y92HewAQzOlakqsrsPyyEi
zsOM4sNa59yU9Mrq615vj8zVrRyLBhN1GeRGGaEUUDi5+4uw2KR4PqG09hj62Tf+
etGjn+tkNTIXy6IpdDNzipZL04vCN1sUpGTXmmvk31VIk9tQPS1K257q6UnJCe1k
Bzpi+5rTABwgPdY6fgInbyogR49QeQCkHFxZuE7ft+gEKcUbwA91eCjxi28G6H5a
fYsqIkOi4ySnA0hgZW+kOsyod7TSEI54RVi3kmhOxGdX/NwuHhIt7QBppKRjtnCN
vpr5DIoQSlIOiPgGLJazzCjpgtoCUrZLYYrvG9q83lqJivFyPrW/VzObiAjcOA3m
+agWmPku0zirk7+qcxOtkbiXQcXPI/jHbOmBLvpB9nN+x/W1fck0XkRZxMAa8HAY
6mtyy9BG+VZkeP0CWgjMJEXhlKz9KU4uqMyf6SyrxMM7dLCsNWCJfcHIAzKHw0uA
EgR3b9YYvX3XLdI+yYxF2ekrCXN0Zp0GwCxd+X/lfpDhbPfhermfnAghox4K+QWo
fY4awfvrOtDiGft+jTkuCzxhPpaBDL+JyVfir9PAbgUFyWE7tG9n+ML9nAxFQZDs
rsau0qLg5THkRubMKk/bbnWZRCMTqxhmIoz4U6YBgGGshXh7Cps/gszGy1IlXtlE
Ud1Pz3EDMnvcXdk8LKCFL8JQulzF51ADeBT+xD5sqNGsJ9ETrOXWrXKm/wX+ab82
YxLAJxyj8aLroggRboNHu1mEzMdkv19IihIcwZFffhQ4a9mxfuU2QNKHJzkYnVFp
5v52fJLA/vC7LDkR0xbzo4TxtVddr0Htkxho0SSdxBJUTrgUhr3jSQG662HVVDG1
38KkMOerH2G82vpxBIiEwPsslVVD6MwwBg2h/XkYMZbErqoes+e0FW32kZ6vSQ1a
lk/D1FHcznOv/xHSfQo+NWv9IXeTVLz/fp+mHisR7AI8oAGLYlOayqk/Zzrxl2O6
ujO57FpOLUVuCGT54KBFqECBUl4ThlKigwrwxOpAkYHVGUSu5rGVJt76OjgVzfLu
HvWyspiQ8AOkzajh2o3/7zx8X8UlCRvi7PjmbiZgNMCGz6Z0kv8V8CZ7FsvlSF+7
UAKyR8k8nrg2a9oaAJ7ZwSNZ9v+/5l+3LX83B0jq9TbI0I/BQsmTHYhY31kI0smV
rfwCYGrFmgPR+fIfSn0bct41qlwLV979t2odxm6lKMzp9dYVoSqPnn6sC1j1UQfA
DZbEK4tf/1wPolNKHxAUVqTXHhL8w2VLUYG0ydSh9/z42cZ9du/NtDYKWMzuFkzh
Qe24YGGrsGV9tfXGL0yD4NfPmLyBW9DOIZnZ7BVYNiT/y6Bz6u8Xo1xRVfgpeR+J
EbZb8oA2aj/MXa2itUatg0RICkv4yrTnS6qrwXIKIy+5q7MN36Cwycd9xqVc9hDP
l+/iKaL/F9m7v/JG2VfP9EpkPnNLq96h+mA1+TFrEGqTjpb43Gbh8gHU60ob4cul
gnvcaZgPoj3ZFlsrZSPDi1Oq1Xb4vsr/7/J/uXvad29t037/G/yUo5lNjkvFPEKl
WBJTSAJ/gFQ9B2QhADxYI8CLYCjOON9KHEx7ghhKQ8s8VruQz5/82HbY40LegFtg
grQpXfIBl/FLX29aiaa6YPN2mqCCLJmwyS3rW8Thsc+tfO9cke9X2itNdXc1qyTU
gTiqbqlOkrx/OSvrc18EgeGbznStvsS95urPos06mgzhg0yOEk32ajKTdwUART9E
MiYuJ3cub7ai8V8gkmVqNxU2J8f/CK+8AjTMVxIhcqepfR1Brnm62UgN4Y3YtsIs
dMuyf9pG3IdXd2rAGJKiXtdSHkxcz61Gso2meAmEQWepTWs4Gs487MEMw01IKFAW
sTKkDZn4hohoJkPBZ6vEUc+XowhETT8GQuE+HEVrmnHpqUGbOoGYMdL1nyp2ek7k
MhIUBmWgS2lsPyu2SYF919/88sIQk89CzDbBVZ8kBfQpKSDOz1Tp96cZ0FBzoaUI
5eKn0YQEPeYtALwInfaGjNmz6qsLxGSdVKVdFrdR1BxX5KI7f1EzOJv1lWHY9lmc
IXtaFSWSUp/RSsp9AZ+iQex52ukcXqNTa59GMDkzhVAoEJ9vmAv5ukWeM4EmgQgY
dxczlrkuZEwH9fBwnQQ+b6TfxThcv/kn1oM7WdLIDVlTyh+tI4jKZ1AonVnkdZw1
Alu/xxKb/aMyAw9DMe3gJzka5IH1OyD4UI6S1Lz6GOyrSx9+GECVrOX4CQgWJtUq
0ry2fMBPH8hiNBoX5rPw2y/p5GvWx7ngbdyPzYJyLAidsilE8YfbtE2mv3sykDwF
039KSB/G+Rtyr2oE+2UbEO+bi1iOfJ6P9kqozKojHwNTxiUhduexB5pW1CwuCHhn
4f3qmh6FbiIXeGK8QUTrRnZkSkgFaWi8IDA+UTY84yLt9tnznZi9qRhx/3coW29M
XO3/R0n2tA0pMd1w/K+e4WcGdKFSQWNC1rkbtoMRaSimex8/ZdXaZU/pLRGd7mFr
33rc1OLHatlbGgJrXtfEcQl4OfkEW60CUkZP306Do1iO4JqDafHmGeEvmOOwhXS5
5ncGvTv0UUkq7mRnrLA3f7qS4f1UgmgdGWgCDm9+8eAwQP2UFApFJhT/hTQjJOoi
XmRYsmeAr1oFIwbJmg+71wYliY0mSeUePwR0wXCtNZzoSDMUjsAjx/Enykri7bni
wMssMPPQaMYs7h0Rxzj6a1RBqsy9N70+v5X8HCnJza+ul8kHruXBe5yaYHsdBjk9
8Os46r2GDwjk/OVwYiu28iEKFFtPpkIezbXSvyBL6jiIfLpL7k1upfmK+yHvlYY5
3PsaoysmFE6Q2ibHoQaBiTDBvztcx1aFhNvCqHWPSUi5socEDZdl7miVMbVQ9Lqe
IWz7pPXQgtbJcZbqF7y/cULYgPrgRz8alOxomxKpF6tlC4dLGesnUI31XMDBADjD
Yi5Klaf1Wo2lTbHIruca5QPQkZv9Nzw1cTIRf7icyYOeej/4JArR39OtZ66oxX1L
Ktu11GTx1UkNIhexkdNxyV/7zyHQkJRToc5iXx91PfMJyChWbmGPE98RhDbRYWCo
MyuW0wla7uJJXt9t9yMShnWeND7Ufkt7esMJFSR6xFB1RBEJ2xxhye3pvWjXi37W
yuIEcOkP2lArDgGaVecpjM1Bl7BnFTle6ekEwrsMoAh1ELunttBwiybiNDYoCsc5
PXkpapQgc+MtP5Kg2Eogs7LsKiA+oDSZQ40/7kR8950iS8idqN22i6OfzEBS/i7H
YDPGo6dLSHDGdXM+ltD36sLstPDkCWU7XvXa0+4yg5WIpEooIMAROSOE6RlBPGLX
AvstURX5/uwykyd86zYyBBJNs/du8SHx0nyC62iB5FFwTlWgXWDdu8mHKxDrTrwi
axE2hJd+Bml9svjhv5BtgJT4/prQdGQQN9RPHzfNc46qsQuqu7S/xaO+K8Mq1gOi
1/jFrpx2zsKWICfzWvQnnEkmNR6witbgKYRIA5H+W4PF/i0pu8wFvV23vSkOmMHu
gZj/MYmsfXFIAA2HV1rrOa3FAnQkTmKgFvWWIypj8+k0FiiFjTZQbVRZ7w+j+JPb
R5nTsIAskBtUvsy5LpOEb6y0z0nOxRsrQWqSQRKPfu0AJRlxISLDmmDkvgLVquaQ
1bl7iOdMyOlSKPIm/cWYcPakKp3rVxWLR1WXkP4mkIA26JWwsCxGWqDsdVAVpHFr
BhX0ieCPviBYDUHzw+I0+BWUYNBXz9ANnqwyUDe5vQvY6czf9JhYOFyJNe4n36AR
9VaN56W3l1MIHkUqIezYOwKS1CpvninPkS4Mq4RDOi9Z3giADd7sJEhX0NdVJEaC
vLNFjAPBIcVXrQXNaoloqq34L22nI53LE/C9cFxYQG//GodYH1uSbe6vRgz+z7fC
4F972eApkEpFnCQHd9YRGhK7mhK3OVTfg99R5kCaC6ai8rTJJPNIVTuONZsVOn6I
7G5emMosrNLuoFz3cax6EhlK80Ndv8wNSqYYlKuFo+oN7RQ0WSpJ4GE4himjTGLB
7s8ecRcKI4l9JnexfBphCVnZhnlZD48ZYViAKcGQD8m6mx7ZohOykqK4ZNYkra2j
mlcqTChbov1XEG+l9mXqmfiHllCmqXh/16AhLjhxRk5v3kWtRZk3kVNI3ODfbo4A
dkr0HJLbLDPolNUbXm4e4icOCr0/QYHODHeGEBouDGSgo3lSPDniqBoCAIo25/mE
B0rv7CoX6r9vt9PJo+FpEjsmI2ZEgGQl0ytVMUougFog7P51NxofWT0a5FbNFWsp
RTo+5CBYgQ9xd1pWp4BJfyf/4nsNdhhpkpOnFAO81VRNUdK4w2d3RNhfM+cuj3fJ
P+Wd6OYtI2Q4hwMb36mcwWkRZm83UQXatHV0WyfPv7Xs38+4kzFKeoklIJNnfgyX
+x9z/pJYKYj0ESoOhbyE2OeX16EFJixGUcBrrG8I04VhnAc8so6d6jYZhQcYQX9J
dojSef1Li8Y7VYCfRBLjeMtz7Jkcq+hpYbLubTadFnm87qRKaD35WiyQ3Om4r5hA
Ibvms14iRxUGFAucKxNTb1Bk4FyZtH5+2/b9eIjgNQmzGtR4DDgmmRPTGF4KVpMQ
GtBFWfSoZhQqd+WTGlPTUtg9WKjB4gWNhImjPrYbMbuSCeH52VLsAvoWVFt/yB1H
r1HRkpBSEgDBMgPXl4QfMcIu+yxYVPaSebqpyFkAk4CyYSgxSlfrns3RQvOXbgPW
eUoQ7sRofgNMetYC2wqeBuzOk5KtvnWEMEuWvQh2qRgkWPPKdZ0X0+66Mpw5+rIQ
P3wJkEljXWhmGZZ+OqnQeBzti4+0y3kHVGD6Bofh8qdAWJJBkoK4hGj04Q4ZqkFi
L8ZpC9jlHQWjt5m95bUTVmxA+BkhsgJ0PwydL5UBG7vcMIk81an8JUTYk2yy6j8V
dNF3BuDKZLzVwbJuJRP0CNWyL4CEH8x2il0O9XNCgwM3UJwz/M26sCHTh7PLbSHR
ZerWtYwagCdSNwTsteHIE5lMXmDFGE/c6mw6SsjZyVOo5LuLxhfyA8jKN/U4tjzY
bkWca6VvqTUTLh6h5458qGTX5m2+a5nyBbHGwlmzc2m92b5U/ioFC9PeFMr5rxp0
rtkUTswOF5NmezO9fbbnPkdGrLyvWYSsfMQefA3e7mWBg4xMgn4TtTa2KMcSARtk
18ZiwXSMACXMEpNeBKlEA+1yC66hCDw5a+VNPU3MkOqhV+pAYmhDsYcCiHNBZupL
DUyJlRFspZnGNPaTmgWzK1v7DccXFMOOmSCyJRY415sN+pA3tNqrSSom37NgiHaz
JBeTLnNgggn6xBpNIk6bqEMrowiLMaD36VSaPK86R9oAEAg6c4D/B8a9lht2tRno
9+ILSFuXXICbbSPQtj1WPCpxvhprhkGe/kI/jk/Xvamb68zaF0K3Oooac0RU+Xk2
rOLfUGzejiWFv1oca0QDsRSxWp56EJ/QX/O8typLTyTCxBXLllAGtvCcWj+y7VF4
UcKX52pP1x81wLqriUM1RNUW2+dP1k9U98mk2l96OfMknMsadr08A2pzKKbWjtoC
TNpxNLefPSrqptqpyROvsPbsqXTNWMbj/J9ebqjTbuFxZykN0a0lt7UjiUJCAEkw
cOPO9Q7hS0pzy3MBSLgzC26xGMCNPxi/+7mSw/5qEPE28f1uP9Q+wtKp4hLZtk+d
p0uD3IxzZXoczAwo1or10z5woFh6tdpJiMSpU1oCp7mkxsxRSZx/79y1Acg65Hnj
zJIlq+0nitAAeBHhRfgcBLZnt9+Ztkfcrlw/gu6X9qQwg/CT6GkUVByN1/JjL6/s
EJescpqA1SOrjABzsO8GnHjkdXs9Iw4q8IZcAa4G3QGc3YNb6KO9uLTx3JH+FDQf
o24srv0BHweZ3cLq3Jh2frHhcdX3kMr3cIuOTozAW7bpEXV3F7DdjLgubka/bIU6
Xuz99KjnlJyRnIDaFmBWf6VyKmmGM2XIhK5tyj13CwrE23Dbu5lnRbI1C0+mL5ul
HR3BznBF6VoC30OSg2Ou3knOCVC26m/mKSjik8vHMiZgts0qLaetQeB6VO5RH0vy
hdSP0v0+O9WluDQxnLoLtLTXCw/JvlL2LqSt2liXAryJKSTisdVvQsSadhlciPp5
3FV25apQ8KNZnb4X88P0rJY7/5zofJnkG1nLDHC55Qa5dTx+T3lHb9Ils8nK/Lnt
HwY4ms9NxXeB3tmUe+A7uAXqLBlE0zO5kHeBuJnCsAT8GywbFXvCBU8D74yEbpuw
FBEcAfHc5yGJIsWsnhEg0VWQWf7vLtiKHwZ/vrLm4za8+db6W9cdRS9lg/1oe+X2
knKYQz0KEs6rjXBtwXIP7KyNxklMBdVNBYdD7qBmA2VC8RXQ0jpu6ikUCYQZDY0D
MZhQXBo57d7FCCb9zElpnUr86T6RXi4bOyn81yilgnlJGChgjsVgAkGgTlvhjLOb
kvBmdMhiAj0sQYzoF01oQcb8RU2CuBZPAWGX1PbuYQfw9MFZJzzoCnqG75kiVaCZ
f8WzlHGH6tmSwSJtvyRixiFEH5p+9Fpr1D2m3X+XH9c7/+iFITm0Wo1GqWgqm9UD
ysnd84mPt/z8/GLiJuaNc3J2n7IOkLFPEBQ9SewVh8rlcJ7N+gxtYbpftn3rF5nu
CmVVvga2VCGF1l5EGROOftMKaQ4e+bhlim3teRViQOTZpz3BCuIjaSigvaOCofKW
nnSTD0mqFimaAzKgne0uNEIS+3tYdOGY5oUibPNuA4Rninhc+Y8XDg85BbPJ6w9J
Sr0Zzc8XHkVLJ4eab0Zmq2B/5Kw/hKK8NkXYf1VdpEFWQqvR8SHsbtbwLnwHgf1o
KBLpW2VTlUox4p/DpJ/KfP6uaRSMaqxdlUmDOzGo9LM1SfQoS63g+grk4sRCqkFf
+737dSgPbO6O32sy01+6Tc6kRsu9LxxLuNXR7gCady+Vra3QQa9jbGBlk0PqmTZ7
9kgv6brcz1ey/vuv136TA/wRcy5sgFt9mPhblpLHgMnz9WGzvHfINM0xdm31c5uh
psZnRdnU3R/gzkq/BO5MjkdloNpAn9GU/ZZdinXb5MPRhnNBV37dMPmIwHwXPGS3
fm3rjImyJrJf49Aic8S6ffVNtcmZAQr9Qh/lSyJYJBWFY0kLX9VwGAm73rKarQBl
pHNsHFt6xo/IKuvZJg9HKIUMX69v6lmD4UvNHgBtELH6SYvokTSnjNmImBGwvhp0
GTeDtkeYGL+5/CaxKuwxzpcTlNFPmDD+ROwpEsNzZTHRttfgq0afHjCxOy6OTo5R
ADDX/p7Zp/Zmtj/l4G2RxYyio9eyx2889GLvqTPzNLc+PJi+HWmUbyFPL8VZHjle
lWu6w7kqOX2hbK4EwDbo8QeLWXjHCfMSDRfJ+Z40674dQgc6GWp4TtcUcNuUZdoh
Rz2iA1/jwfK7kxhEhKXYK+34uMls+gmww+HO2UNIPYxC9+R6Lf0YkkpmInuSKiYt
vAyOnMiVdxAYzxjXLQOzFWQKSY/hEis4Bl84i+L373GRdNgU2DkMfM6wJqtgUctA
MXcpFC1N4JfFfLFEeHXTm2f9wchm9AfGL9YwnRSx0DHAGwhHV/jNZMbDchax7S88
dWSOyx1AUbwJjhRrM9Nf42GH2HzGwSsent2xWGr81Ox6AfFjkEDetRdZSUUVKZE9
a59Ng6jvAFHOD3pYQFP19TTjw9B14Pu/ev53axspcYhylsvX3EnO632B5qklodSX
8r+wGFTbD8mSkWq5LQkClxgY/a8jqKg3xfSIht3l+tjSZFgh1vmRD9d/qurljtui
UxIPLVAQoUr1VhUHbROc+UImbjo/LBBrPzw4rf+EHegs2whRfPvPzlf/sKp3L92T
Oyp008eNTzt2+6hNrEWbQuKfQ8eR4rPu51YjGxHv0UbyKJKAuX/VrtQYs+4TgDiy
UHzBumgiOP1v94tGZjeVEIIcb7aL0bLfmi1mbt5vVsBHEwWvpyGMa0gX8CWUxf3a
XbKBc88aRzhmjPW3z3vGlR27tvGcKz078qXCHzXtk+WM5AKLOG9LdZsrtBCDs2hp
GPDQTUMLQK6IMBK29FK9YUXhusYs5l+sdvExga2jQZAXmDwR9vQyLaebd7bCe3Ga
lms5zI3jmNjPNiBvouX1au/PjAK10vbptXduufQSSPVXisZNZFNATHKonSIw0SWD
f6yZb+TRRFXHmRLIfzhd1XBKQwqCqDQXczLBwkvmqaqjyJKLbwjk8BjD5gJ7LoiH
cyJ432Sj4vHOxVaHUtuVCHZejCRegJ2tQ23ijTlxg1noNk0OcVaE5Q7C2hebib6F
lWDQNYZxwDLGJV/5rbGVw2zZe1daGy7g6n0fQ2rqkmnhfuFfKgGZWuEz4mJGFm2f
KXo7X76kv5vimrTgNiegdSWHjGK/FKW9We1DO2QLSJDEy1t6MYG4TjD17UEcOjMa
sA826LjgMrrSfhR+mBPgLqjib30NDPLlMaGW2zkB+QMBwnfhaAF0JGGqdcestw4+
86mdWORYY2ytZUqwJ2iSZXrKomqfWtXCX2olXHx1vMzhAd2wqF7QcFjoU3rqZJR4
zMKAdN+up/nx7sBhAZewEoBpaliyXjd/lBysyEtafSX0QqLzJaynA7k0VfGWT5rk
RrbIlgN84sz9oDGSsrc257Iq0ZZZlWIWCLI2YDNgjjIegJzRWmhmzcobbymcy/Xn
6oB42VKNz72GZMTNA5JISC0fZ3rnkz4MxzdiM8IAwpRG0Nv/TmO6uZ2Ir9H71K02
5kWhdqdoMfy/p2OIXC2rIGzvO+80V7HfMH6xoJfjGnGzPVU/H8gCLmjxjLOHK3Wb
R4d25aLGcfi2BwH7nEDNEWMw3fY+RRXr4U7NA8K9UMsiwx6/dgQN1E4OHjS9LVur
dyumQvEnGgL7yoDprTQNAHserLVSSJTIv+Lr1hc1XxhXm2TScPo9UmqkoCsAzEeV
OdVztf/ZuUj0bNxIez3M/VPQ5n6Vbd6Cnke8Y+a1aMIXyxcSi7J8Uw7RBB/7L1bF
8XvzgossEl+TAcmmNITg6+EuPcFapgcbFgOUisK17iPpaGIGNrJRsvJ1x+B1lvnI
NoOTi5lHhlR6p0GlzM0qD27ESX2VJSlaE+dPC9QwcLg/goZ+JFwAZbFazLE35ZVE
EjHQ8cDncmvYTiAbieT8h6pg1FpI+6G/SAuWQpN5usv4sK3L2MoMNcJVBWaLtFLl
4goskKKh/m7h99sSMzoGQFcNeloP7wHUbhVDCkkEwzFNFA9EF3hicK7+VIteiZmi
71KAh/4YJR7r+tY1lgB6NgHI3GSoftkXR0/b4JFe51nfJkG+4dvcY2HXF4j8ciQO
QBMYr9vTxJ9XSWaR5hj86sNZ7QFh4t/5EKCKou1T5up4X3ZCqmG4hjeWgLmT06fL
xzGiiTFWFYuNfz9OKXUNJYD1ZGrTAe9yy4MW4BLVsvP0oyZy0umeAgEKm0hqnpHb
lFxtLX+30wpQ/MfhdYyWcp/lFHiRQgjitXbk4ho4YNkP9vqFoGIYLtDy1bCGEaoV
Nt6azeHpc643fvGEDuAK9FgxZXddWzoM7zqK9T7OYByEHJKntxMVJeXnqF2Glrhv
dfwB3K1Lu0mqIN9X0fJa31IURUpX13yKO6kgICalwSY1nHeyc9+g5iZ5ksrmV9M1
cISYVYMxSbqWWKFujsiWuCwX/ZdlV9tNA2NwjJP7Yv+Xxk80P41QHSbrnNuxR0Op
ILGPbqOzt4s6rbQpA4TJliUbOWREoLi8p4nXOHe+edR0ffxO6VeOwNfeuVajEXvG
fFG4cl8yeCUyQOJaA9nHa0t8ytpMO5Kx8lIoM0ypYTl5dprnXO8Qf/kisrNxzo/g
t9xxBOmIi0k5mJTwVhGLFRiFznbFlAUho4EhUbhRMPYOD7e6NW9sm1h0hrk/MmU1
RDK/1oU7iC+d6G28E1HARRV082vcegPA1f5g+V0yKtAM+6HAYc6Qg0rKfujwnvMG
WUzK8eTp9DSLtqLjVzkRf6ZqedZmjmWsw6hPpLVHRKHtHxOap1ixfX4hqiLOPnz5
YEBE69OzyTddtSjigGi/lpduYr7EYRBECP/W9CY0g7jCZuxVCGaoVFRCW8OsnhgY
R+Kn4QwwpnWWxibwLNNKczZnfgRr03/nRiIWMNaRafY9B8QnhYmsGYbVwzeSON98
AIMEFFEz90MMkAhMgNmp8HfTrUueV4O9R0BsVbHQEtDbVSmJ37CLMBQ/MQRCmY7H
8ve4YQ/HOEQ9OHCoABe0spqnps6Aq2snQH4zjfuHGZRMHZaFMxYzujs2/sCbds8s
UpGeWnRgYZQZ1f4ELNLT1ffI9IBIcyZd764ZGy1qsAPsa+Qqbe+OFw/sMZxNNLt+
VSop3Ce1XNkC9n2OX49vFiyomyH2CU+LAYKaTZl2GxPrzh672YWCxx0wqEozssBn
LFPWo+BEMysdxE7THBCZBSwYuLM9nlh9/64HznD92BFKmnYX6Xfc9n9G7LykGDfy
40VPOrtEoBmVTgSIRKsDBsrQVl6NhHyi2GrN+sas3AUuhyXDp1LLAldEm74ge1NO
REWa6spC+KljJV0o2y2pc3PGqIh0noOBhmB6CRkOZGUSTugm0IaRLTQDXVKonjVa
/krz8Hoy/cLAEZ+Djeq9xlArgJtVUT+DRj60PupOKpjHN2Blx31+HMFaTBykCXJC
ONV6UGeNpxQdwjs32e2MoPe2YQcKK5eYER49dkiP8/blGgvKAa1TFT+j35mGCJel
hZnkyCljyhYL/qUudaizqOVFPfwA9Y3egAWum78C901+wbkdJ2AIVH13I63Eu4ph
c/E/4Eody1pvATEN6CFZ+exK3vA8x1j1Um/MPoNEZ5iOqbCIqvyS9a1uOhGgOAW7
E/5iJka7udtrTOBdTaoNCPqI+b/dhgbzaIr1U1l2Y5LRcCIoFQhbXIxIEX6EsIw9
uiI79Fi6E/oz9ypMeukLjHNa/G8KX7NvQCCdAPGRQ9fVwCKLAVbuljXS9OFSFeVy
y/p2uhpYHAfYl4V2zyMhlpytyQJ/Fz6ctc09krYfR0NCMs99dPNeP1tQJioa3nEn
8pewA1IEbCWC5OzcvUYkCd8X1ed8CGXmzBKmpwvtWWWBKgP+xwOEIia0JSxTxDgo
Vk4wLSafzY3q76BdvFuFkIzL81LjCq5HVZ250WBJiI6dF/QYBuK3u70kCgGGU4Li
rRlIMFgDdFl5gYFhNeeiD7bk+25gYm6eDc8lE3k4w5HRsTsihOKS6mgENT3mkdSy
KBcpndEaCCMTJ6XqpgXRDK20fQX1BRfLO3Xp6dI4PObTfIEhkySnC8pwpSMjyfLI
/XXBbHCR4ofiQx/ambARacVsFnbzYOS0bRQtN+vmPx1yelmXZv4AxXH8v6Ad52Zs
Qt7mZgL8du0BBsHyhOz9U8Xh10cVgER8iBC96vQMQJBpUnAaU+xSD4Tet8Uzd6gZ
J7vWj2lVKPDMFKIR0iZfR0s6ddlxlgHQaedx85qTlJQWW/1SfAIFKcCYLsCNgMkT
5/bNGeUP00ZRvu5BWR07t65no5hyYM+oynBDxBxt9E+y6ABzO0RaMDkLXCfTv6eq
glW2AizCyd1HORfa3rihIk7WhxaXbYHTMMJSwwftYJlSUIOV6kUwXNL1A63E/gZn
qHTxzwxaa/VVJ6Jgi6xjcaeBFbjUwCf2aUtJ60qUYtt48C8HZu5+wETGSwh1dXwt
zCAgTxTIh6hQAnHiovpbmcBKPs6EfJXq/Y5pPSthW3SRPExEGBZQeln4hcztZq9f
P64iaGAVfR3VDEwkwcJFbw88pQJN5Z1qrqKPKGlEeZ2ltaHrFDh3FusXjZoLBB1p
wBagBWvGmfozBnVHug48HrOQMryif4kQeKW5D44F74GjoaUz4+VqDlYVfScwY5Dt
CH2fnjbMTzSKivm9PHT00hMb0aLJrggbo0+yGx0yB2qdVr4QDu+2fpxDLuGtq5TM
xc19x8Zbk+w3/hpP6xExUVG0az4vgdLNSCpoPlu7ZUpPqUjkL3MSh6WtR+b3eWqH
FKIy/24N2fzKfCF8fJ0+UQDdXGIRneJ35hFazX7keSHZAgb2/MoWGNpXNbq1YS0t
b5EyHbC10bHoVJJ48bxR9WpuFNp//Ofys82YrshjzkcMw2VPV6T8E1neR+4/9U8K
tM4zn9xqxYjhKjzHlY5uooQSNEGtWF4yDazJSXoZjs5XQ2itNiSUXLRAKfjxtFuo
nrTpvZmaHXRwJUgSKeZ4zPEg5uz+RnzlZmAvx0Mseucg6VaZRDYBFqZ/0SKPUzAB
G+fVk0/hYV6eapgqUpk9wl1gkMtufoj3tBG7OYLCf3gTFigP/LB1v/wyhKwSDrAX
WxJdJ3MAqYGeTVQiWFxsDp7x2rra36OjuISETK4g/dJUF93mm/071vIuOHcjIYDp
2GeUowR7qUfiFZxZfQz1fzMOqjq11Pv99dHyYK48zwtQY6UUtiaNB5R6oThE0cHE
VtWn71bjcMrL1e00j8OFf0aAktMiql3nu8F1R5cv2ZHEN4XoejnVBFWYRgrekqoI
DCrQlbCGFQMntKk/Em5QxI638C+rAioddcqXHG9YF+RR5GC/HfYVUCEJQVlUDubk
mKnFtm1RbvB0dOZrNCYvJ9otJNYSfdubKBaNLQVFRo093bsDrDtj5AWVQcKW7Za8
1Eozn5X+myUwGw21Fv9bY+ZadquX7wsS2bD6ESAno4SdZG9AFNljY451k2i9Gndv
NxFz4fDaXwjTMPDmR9xxjW/ZUl5TwadbwyhoAUO0ebXv3QJgOZ8WC8XPixou5qPK
W0VtMaIYEuTteyjNq4eoHc5MSdFFkvnLsmu3rhCFZfTEYjzvX06krAqjo1QU0TSK
ckRdFu3xs4+GhFRdoctb+Gz2wXiUoldSdXzAvZl63YTo5aAC8kTMI3hpOf7RwpjB
rXDCp7yEqhkVKfDqcjYsBn+JMHBGGds/N5aTHjAM+ryOo4WCgMvCq+2O7sCoYl8e
Tv8+E3Poc6WYDVq+EKPTvL18VQAr0F5dghxOXdHb2Sy/MYzCVjcah8TREkLZBA4O
RoUTkpTpJSvtOvZbRpUWuRw4SrCoUWFHBoj25j/U4NYDqUvvaNZuxGbUiA/BOHLx
5swiHEwyOwNNQc543rdbx585ADD9JR038BjZu1OKNLyrWKeolZOGM4I2BZrHtIDM
njX+O3zHdC2gFNWLeadyP8wO2XipDkFsyd20+nPJmRXaNsDAASLwxXw3NFn2oDrD
cDRiMGk7xs1LFHX1suR7uCXK7jDCpADJYDmCdwdcTZwrmjfZHGEarhmF3s5qts+g
G1Fx7kYUUn/L/0kvypRNmZzLoaCIH/Y4GM6QLl4Hq2arxvswIQxB/Tcve29BZZUs
HS0anCaWeZFqS2Dsn8vHZDYXTLQoqsJVvD+tWoZEAszriUAYWhbJwOsQ01HS3AAZ
S+8qBcX3FdSidABrxB3Lt73Z2DEU1VsaX3h2DVA5qpPf9XU6mehD/xBK8BbyrAus
Vw+O6N3xLU3+LYNMAAl7DCuWMzftWvsnm4UhzskuSyBw7GrSk09dtCo3V/Rk/6Y4
kyg6ksVb8iPOzFGaKdBgXHQ+ljOHlRvBssG3FcRhvtQs9wgMLEh5VXz4XmwmY4YU
y2D+rBBIk2Cbh850d4fP7jPwyd6X6uM2gmqiJRPCRfPJ3ywrGTwjFVQmgfYMqRgq
avrVzWH0d+T13iq9myOvRAzjlxsKJub+98b7+0WSL02X42nrOHVWrz8rNH/VW1b0
PbHcR59hxwXNY8Nrd3NXuoXJwQl4LRvw1BeTBubL9/BuerTY7C62vyfaVVJyH0sJ
FMPeqWRBIU1WEUMkSSt7QGn/zxWXOFz1Jg3u2SGyPd5gqhdakCYNET8oNH3A/X2y
defFRorfLHSxpmgwVbyRcw65UuPyucMfPVBD8JBRAFxf6QRNUW+xx3NAALUUqKs8
HuoaYYqqm8FDpyKcguzZKlecrruK42WB8eWL1Ekm1/MFtBA51nZynMhhlpmMFJCT
I3fzx58fkksDOWQxuV7h0aiHHFn/3r5B2ldB4ZfI/mfasWyRueW3CW8t8pNjiXtF
qliLYDfynO48gNU8WaLRG+RjA8+gyHDwHovQJBmxgBnqE+Bdbs3EOObM4eY7LdIU
y3TF8kbLc8x50OxsV0xB4BAcglZ0wuL5WpdUp4Z5F5ZETAoN46+MHyQDo+Rh/F2Q
cZPV8p/8KXrgGkyu6pMJs/HT6BwoD3XmVCoRhP+AOgQrp/Nk6dHf8nIGr28iV2VA
ZmeFsfDpLbuHORhPFPNftxNSq5tY2EeoCuhtl6p7w5GZQ/sDAG7ZoR3nYDtDUkP9
k060cvQNusK9mFOP7Um0mH12RELHo2VuviWIGDwVFtu5/osKmaLrZNSE4xjaf7Ls
DM4LcSFyUn2Z6nIUrjZkLR2lzllS3f//lULNctIoHqg2HSRHR5RBIt6eGmpQd/CA
F3L6ODgbrYrxhgnSveYbFjxqvbdFQP2EVqOggJ9kgHR1b3y26tHIG+86yla9Jixc
JUqQRBQnYOLA8V+7xyou19+auJvf+jjMjl6wkPVhLSHSrVl7gv1m0G2DRWtj87Uk
oNlI/yy6cDXj7qgPelk+cNII+rluJjoFxeKGK4ZlNwedX2V+BPLAl2JeYcCRgXss
QMxJMqLYdE0TmvK1Ycdg+z2hhW7L+KdFUEwjTwOpyxiRmc2+G0Q0U6cDIZXCIfiG
Ty0jXFW0HHBIzjs91sdm6uuZ2GVllgA6KlIA9h5cNaopmf476ONWnBOpYXm8A9kl
RSGEGrOa9ijSXO4DLwKdhzq9u6Znb54leibf+KcyxIlNZluei+7MtrP0z0kyde3l
g6ZhFLK4M2A0HMSP522t4pehf5+xT6Vgi7YVbH1wfE8hXc++ebHNqWxbcbNRst5u
ZxrqNM6X23j9VQPMyDtjc1J1g9Mb4lpk/3hNuqFQ1/JpGcIozrl2zsdFdB87pzzj
oeKIhQDOIzaVURmqO7GpTc/KE1Y7dNxoxcMLDwsxvsrnNwqGB5a1TwiQFLJpN7AT
o/ow/P4MNIAfV7Wdr2TN/grlBoOS7WXNfSvuqhupgiL6P3Idq2JJHJJYsNN5HUII
iGNMSki72cK1VxRiJqmpJS7nWPtyKFxwZPqrEh0teZIMxWrrNcNDqqLa0t6w6Usi
x7MzCy8mxSfsxwQyCPksBSAM2+Qdt3kmjwiRcLC8OxSgsfiYQZ9D+Sebz1EqY95e
TnE1m6ASo0gLHUk783TBGFKFHiHfCPvXYemsyzEzDbw3ov50Fq6VIcQ3t8c+mv1f
C8k3m9zszn7SbtAS1A6E03p48UdYbahsfcya9NkaxjWKR7JaEUuSUzGE3pOPNv1v
VPCL5I0ZYxjjQw+amOuq8razNWrrUvdRQeh/ICUSfH9Az2MPLk0NmbdY2iqDjHf+
z4T2U8svX+16LJWL4LkoNi/HMnL0DDC8FbKcPHI21iS2sdr1dvID/e52sQfaA0Qh
QBGabxpd2xyjj7yvgouDt5c/8VHKeYuVloE7ZzarURNhJ4cZQOsCcQi92Lxd/6BQ
xRh5WQRIlY1sP87uIkdh5zLECqa6V18iTjsKR02lQ7/1WsjqBxXvH3tC+s0bQjqi
ommig+45T9ffzxcpErfpMOjzSIGWaFlVameTrXl1w4VeAzTbLKyCuQVRs+2sBwBw
/Q9vaKPzakgStO05YnmDWe6OCL8OwNfpdL0WQf9dJSFK3P2afVj+X5VSmuvB+UjC
V1Wmejl1da5lMyrk0LQ8BlFMOOrbFOPY8s7Ku8m7GJxIcmPUpPvnFMJURHEPX36e
t4Kdo1xfmg5V6j3w08D7WbctAswwVR2idXgYfb3VgZU7hRleUZOZ4SIwNpdUy1Eo
zuhuJ0g+psq56ZDPSS18G9P0lolA32i34avFee/3ffSjI1TTuaB3g8p8gZYUW0b6
B5jNvJBX2TIAdTjnA55LwbuQSQF46VV651R8AgVlKWGGfpreu0oYAfj4EYXyDlO5
y/9z4G85+/W4t583DlMoDWPhQoHpiff+8nchz5lHnHos6FLHP9LUdGane3+M3IEE
fc/D++1muEXc76puSR/Msi9PD/32HsWY6Erg5W/hU6ljAX8fSTq3LtjW9GxmzQ3J
e81bCeX9Y2GwaU5Xb4ytv1EMItKiQTtYIbtaJcFUkRwRHvjpP69mSAqG9ipg/I75
Kh/Z3kgGtGAoUVccQwP4Akh87Pp4dNHFrZufJ2Sm0hnSI0GWTEkn+WAGyv+c38gJ
bG72zQnzljrQBwaDYpQsyWayPSH2PfgbRLQ/24JMP6Q+SVKRoQpIEZYzQYtg8ANu
ECjyt0LQrn3U3K6jZOmI7+08cARi4xt7ESuMOpGB2ebj4A7w6T+I3CxVq4GJ6xeD
UZqNQsOPa5PtTocOAX3bD8qPBXi82fPZ8QL7+4c3BVI=
`protect END_PROTECTED
