`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oh6vRMCmzYeCXhkdVn2CdSD2vilc0HOY0X3JNKzEyrGJRVF1fs4Xyz4hMymgdK9T
YdndRtLXbud5AoDb2MbURoaKmhNMiuKNEi6qWsupbCv0ba1nIQkZQJ+RyWMR1Paf
w2FmJgt43Jzf9+pqI63VjxCnZ5HGrTU0yZbStlAlV9udAxxQCKrqTuXAybvI0fX2
j1JdRBJ5jVKqoTSbkheGRWOz4EyWLckIXLYcK0T92G9CFtyXcDeLQ7MbiEcYlr40
asXNFLgpEnOGxEK8v9PEPnJdZtKiXfuGcty8jul0XTxM0seStTnrUspHeVf22hNt
O4KexmmtlJ7nR8uBOlDga7J4i0LQk7O7XdZr2hGvzzRouARS9bMskuAyyO/GernV
0UWZYjSlEE7aqhnmtAHmnRxEmUkC65KXoHin+wS55rXPyi8H4sM4CKfsFYo02pzi
T55Xyc4DwQ/CJ/4igtkUv1Vo+XXx5rmYTp0jTuepPnjWGvF56MAXGcVxFc6PlcF0
T2Dg8SSyerr6FXNPib6DzynrwkAsUTgrTCJQGQO7xXYrpCXD7boHXZSFuyr3KVWK
OjGKyP90wgYs+x/9D9cC+/ykmG+0CyER/qiIm6Bl2+mhGVKgRX6qd/40eY/FEaY1
OeC4Ofcc9N1h3RqCtd4ybmT+l3nXg5rp0vwutmtFGflctVpFkgRgd1+yEPaZLXYM
6ISFOb2EOZYkZE9zA6AwLc5xSStCjo6EzsXA+Lyzu9HJLql52q2FniJxK6bA2oMf
zcEKdN3mBmvyfZN5pbGv4c7xJ8jBJbsfqiEaoDOVB6kM9O1iOW8gVFXbATvf5vX6
FGClrmihEqgR9tvHKaSL91zlsTX4DLP9LTdB3eJN9EwpNACL7FcS78+qiTgJlgNe
DQM4qYTlMXJsW4VfamkqPjg9j1AbBXiRn5kuo88iv36bZmL/+/dUrTeLmPUIWUKB
fz0ms+OPxEbn6+hsQbl6RLQRz+dSt+cYfR6hZ3naxp2v3c6rYlEAFiEsDOjaEIi2
dRyY35qMje895XNZfsoAKMbQKoHOmMCll7srCRaZnAJP43VJdK35NsXF465dqvzu
P/sn2MNlHZgznX3iCezzIezjraiwXQxAKtU/0rQHjcei26ZhZBxLR2GXJnbkmFmG
6Jo6I5B/koxdB4OzIjDJCXCHLRgwKAvqLravNS5ZT5Hg/KYqZy7slTUVd9BEj/c+
XtjUiCVhiKu802+nz1TncgO1MTYRv6AUOxw1ukJEhu2UYPI1sQAxbXbppO5xdAyx
Z8aeLJe/4jfu61+TBvpB//lYZCBmD7YQTXnaa26kBi0=
`protect END_PROTECTED
