`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ElerJhxTMh4lcNogoPK3VTQUsJ0CQHIHZwaVIwHNwjIlLxQtecNDwmbMlYYgmfrm
HD6kZYBI6VEp0d1Ce445fsW6ZIozFqtGBy5rXhbp61yQY8mwwRGhPKf+BA5UoUEr
MMfOJ5R35scVcVGLodtuR3E19DXaalEMxsA+oCTqFc43v3JTNTn7eR+G4NTSkC87
d+yFU7NzqrhEQvjQKdUD+EHyzAY2EHDP1riz3r04jduqM5E9tyyV3Aaz37Is4Wyy
zEHvprgN05cwaZDODegL8UcQ7FQiYfKRlVYuStjq2gqZGTkmaeaVXlQH3GTxFR8f
wKoIj/L/2SkmbSvZYuh7ZzjnBOf/BAX5VtysVYRvHSqdbQgFIQlFhTxJY36AYSGi
lI/OUmKqqDMQGLAlFZ+DR+F8yN+MQXHGjJT/aZsX/yFwjF/2i+hBf3h123wzFYcY
/0kUSbAosINU4P7EoWZQ2BpJ+eRLyN3mzsD+WI+pvkV85WiqSeaYyexxb2Q8vNEe
JxHPiYniydDBnQqUhqMLJAEMhRhV1S3+Niy0Pf6ydTFybzmSN3o+Djhuz9FAkji7
THPmXHT0T+N7S4HV0mf8GU11nZair+inlxRJK1BODZo0eY83sm+WuomZE4SnjME1
QoSQ7SvwyoBrRHk+VsTIshJts7w12yiJgjGjUzQATR9nTyKkfoLPvtnnNy3m7aKy
GcbGgDlvd4sQV/sUI6nfhj3aFfkdWE9/j96UA4srLo4tGkEZy5P0UuXGe3lJiOza
Fi0JoItO6ISfIQNy7IpciauYE57yTYNsejanMhOywYXNegFZLVaVrlVkK9kvFb5n
qswlfxyNA2b2tAjXpw00fToAw1CGCQkM7vy9DGHyRT2LkigN4G4tqWGZs8AQpyMe
lmoFNU54/hrpIuQodd/so1Vjq9bFZVuCGXJUfpmMMqD4YkUN56A69cax916wBsVU
NprvX3rNh7IHLG6/BdMLeCq2+sVTaSqHg6UUWKlQTxdkAY1ZsLbL3A3GsY5PV8/h
ZA9wG8FqteAP9tjYP12H8w==
`protect END_PROTECTED
