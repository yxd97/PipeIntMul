`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JTtjj8RH1PtEiICdXL3M0vKP/CQjJffnvljcAcEDHtrzss0OjJsRD+9zxLvzGy72
xdFzMg7NtUirXm9oieTz30pt1ISCPp+F43FYjJ05PnlUEQbsO3/FFwKcQD+6iebM
eAEV8ty9tMUy2DOjWuQOJ2bXeBb7LORYiA+yMHoWRFRU/Xk+WWq9QKWTO8ejI70h
PsLep84HV+Z7wSoQH7FNPHTNj9MZTD5d2zQO/qNlaRk2QZvNueMlrpFYgqNGcilC
URbYdiCGoWUNoGQz+66HkxLT8vu9x7vjbKuBuxI2CGeKrxDwdHlNs0fvZBYFAE6y
rT8VESzR0YDCsf+CCE7JUiouqrqhEdm6x00CCNhPzeFAZscHfu+Wse5VY0VB73eM
qJ0CYLmgvtLrtPF88ZWnBIJvPSBa/H8i81GTLkYGY0rg46u3kQCBqwjj2oQg56VH
Ip6Xw0eXO4IhxAG/FLKKEq/iqLw/voT1ZVe3sNQSMfMX0KSCN/ZvZ/D91wwfhF9z
DTOEuHdYebj8rBGoAP5pBfyFTMb0hIKPzYaWOtMsrU00B6Wed9nEjPRc0Jm5dMNl
GtjzkQ7aBGNEBw3nRr6MgBuQSJix3Cor8Xvc0lkdzm2JQ8bpCZgOEJtod7/oIKUu
wnowafP9TFr39sAfhFiUTPezBRTOPTVkFV7v5QNk+7oMzD6XNc6fPAk/OnYNcOQM
EzcHdbm6ZIFyX5wN7INGIEzD7V0kSE6Y3Gh8ZhB8So9zKWppUCt8jAevpzhoO0GI
1D75lxm2UIymhx9DPnPThvZ046UDpCoSb3gVol93n6oruiUtKirn1YnpsT39p2Gb
gvwx8QRkyqsoER/a6rJv/MpsiLOCCzSOaFxr9gYpOjqyAxKgPOdrWl74346PsmmT
gQMt/8YYvr4k3cZFXcoNpQTi61g6GW15bmEnfPddpI/KMNGV+TL5Mb/c2vE7761t
IFjo8Bi197nsbc11tAzGR6HEatanb4scHEh0TVPmVRMFN1Y/qNMvGZq2DU6wChcB
uSRCaFuI79H7s5RXeO1ivuubO1xyNJTC9NJsXi6OrzXGVSjM9QXK9i/vNYQjnlKn
8yiZJytYh8pPN/RPFD92ANaBZ+tymmPw1wRjkvuQg+Zbh5SCi4YZxTqS19bJh5CT
gfj99D7rRn/DTd/GvM7Yy56yLZBCYXtsBXhHevLU860FCyC6LYwjPvaEGj3JTInx
uJFTc/ag3CV1xMyDCKXJuWHYjQwutfeb5RBxZLui+ebL582Ip3Mn+5l6JJ9tzHcQ
rbpEBvXtzaV++L4cUKSFUYC8mKFcoE4fsGk/zF9WBiy9dZoSke+6/4fTd2+REinA
8c7zCmRNBnFfp8IFKwLLCNTtZGRnNyWDFMnqrJNTAELZE8i6Aa6D5gQYBWJ/qDq5
FPHFh70jSdLllDl3/X/b/VdmJ28xsa+VvcTGZ2VPGr8asLiqkWX27fgPXS4O1Gtp
LGD0KvNSDfOAKf4V76FAlxo8MgQmMJpvp3hkeHHyJGs69mSefQIctS1F3bKv8UEe
yWflzBzi44JLJ3UzO4/tA55sfCb6wnCGIDCBI9SuKL42VV21Q1yWq8CEiELUoGKj
Kwk8JwnkiuLlJXsxkY+p3nqe9tnyLKS3g0EYyRtTRW5SgbsIDkDcFq/pIKGcNibS
T1uhCGLOcsxUv8IkKDcMJwpyHRTSpHfeiW/2vMxUnMSG3ZxKGNB31s67yiNNdSW3
HQEug/C0dMHQA01YFnLZYh+xNlfCVhIiES5/bawJ2jArbpugMtxX52F4QpvOc82G
9dMTEfcSemtW/V8kGbNW9IPtcjoNtKKlFvFTo0+S+BAG9zCLtrMt2PCWexSniC4+
bq6XvnEF23VqSpB8uiftdV9VY58ysq+RYVwR7qxsP11D6hlzRVk/DBbxgUO8XvRX
x/0tfWKf0bwoSAQCmcyRTxGINn+4P9cUrwgfrcO3RE+fD665BN7Q8ovRsYeb5l2u
7hxIKlcLwLW5gwjr3lXrvnId1AoIrTGwdj0JiZ21RKvcMOeZaPOm3XnsjAVSKyKl
2rpz6DBnz+wD1qnfTU7w7bFm+XnIvAtxzAhQ3D43fC2+kqrp3MMQ74HOHxTsj9y3
i/Mdkgv/n8NebB2N9c3FMZS/uM/RehQA8UvAbMWiN1SHRPp58qO0MLOy+cMnJQaA
iKtZV+qzkRTMr5lrCN8WiTY1OaUy37NlbU+4Lhj6Ga9C6PiCQQDjhKqjggVkN4+m
ez77QI7gYAjPrOmHBNw2H6NLRMuiFgBvzmPcycY76Cc/GA12ADvdNDG/8/HkMh8a
xlup6Nr25Sl9UVhsRv6GSKtyCwmg7FMId+GeYvFqa5W7zIc5A9DaltUFpguJ45Wu
CRKZgJcQ7WMQg/6q2G0KzzfhJcVyJ5NQ0PteHsX+6NSzNogU28eUAfTazuZZUXFb
ucZwxsegoa9hqDBK7KoTXBAJv+RJ3CqQGWYtcHLDROK551y3n17cKcjXRNjrMETP
KnKzzcQj8og396MFaFTylkScmDPxpZODqvwE/+rwlds=
`protect END_PROTECTED
