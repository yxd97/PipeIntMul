`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWcGfxDwgzFr/iyIPdvIM1zKrbr53xP8qpXLbDXW6sQZhn5cyhezGmgFUTaJ4J4m
YnFNxLnySUgPjx47ACJehkzzwZnu/ZmrKB5Sung6zjxybcDXpyKVm9/JUluwfJXH
Hl5RZeSLhu93xA0aaDV0coreua43CGaVUZAmp3aGSaE9c4aRhGorlv1Ka/SRd5F3
/SFIprK/Lnq6BDQk7bfnLTTllRBGPdPH/R/JWhkA/9eMs3Kt6Zwq2OKOEByvpxh2
VFuv/WxrM6o+owUPCDvpLgjDJU1LGkP1RPlcLHglmSgl8mekQtLTBWDy6Ay79y8O
0kbCdds30zRnZ4Cxa8AnIaIRRYsU1UaLaGqm88oyOnKJjVqqP/C96/zk2luyVinF
PkKJxLg0V3G2uLnSTQKDT2kJ/5RkNqbC0XT/zb+LaL0aIJ2OnR0gz/eJl80qNwe9
uKF045oIuGPomp605vx2Y2WK3NatVUnXlGKO+TZDqtCH6QdxCqdTWwBEZQDhTszA
zX6Rvgy3XTFK7ylJGF0mnWufP/mxq+PnxbHl03lVlxLAPDjSEDmw0o7a6wsNkvwf
90TDyv7zwRbTI2imvyYMG6tk8Ad38xcsIdgNdTSgZ32KrMrvU4v9285gUgeMQrdG
Gf6qnOGf2drKjheFNbN9yXZKLT59/Ifqw/maPMhvmajftT5CAf/5iHIYRncaV1+q
gUGREOk5IPSXNKUETvGqAB/8AuQnMBYWeRPumTFim3Z6WQMKQbnK5ZMm0m1ZHng3
AfdqL6kHMpxn/PqewaaQvY5eT91HWLtqGYe/4Ar6T5Y2VcxAmuGeUpYc4+cIGKia
cbWhm7nzeqzpS6FRslHTXYBXYuGB5Xi+hJKKOKF+LYbZHneGVFXPg54zI0bU8PqU
PgksMcdJcdh0wEQxL2d0IYZlx7fLPs/1Rd6YfFxIWxBfCvyZGaDuvLjDnYNSqbqW
8lEz30W2gbPtDRFS6+8RVW/AIi09XCjK4h0ptYREDXWkHdIo1EUzh8/2NS8Y2wuG
lfPfYyeIytMgmH9/WKo74npfIyoev6sZ/nFMg65Le/1rRkaTIc1wK/ggznlVsMKh
32K+G5WgCuLH4PKEkFBTquKx804YSgz2tKG+Xj6ilPmiXNacjDmwIahB3Fy9442H
LnjYGog6G9UB4F8LHwEJQDEAsSlEXZ8HhuQPJgHRe86YAUg+OYvtAKAABPmz2ltB
bWt2OS1LGBVSfRUFyrFxue0Z1AElYchPaekCCvZxOx5Eh6Aq7KcDPYNwgMFFOCEw
oDH1DXpPq6oqWy60u8qZPpCyxnBn1DFtCMJ5UtEMEI+ZvxCF8hqvQ1+sc0PYh0vZ
nmnnmY6TY4WNBjfOuu4L02Fe9f0CMjud4jR3MYZNIKvY1faTRved9XMxViqE7Z+a
6ilS2zAzEwzDWqdh9uMXNLDHcKl6Q5hCyGdqB3uAwW0V/7wHdJVZkZHuZhAAbraP
BOPu+QXxsNZfp3/WuiNlpAggMqKEC0LNII93Ct+Dv7+A2xx1JG7rQG9Elhk3QsxL
zlbqM+w9Cex/9Bcc8hbETYVZEdoWrHS6ijLzHcc+JKFdw9LDWlL1qp8tcGwglPtQ
jJTVvx/biFqG7a2rN6U9aWq9gbzzyoQHgK+2vgacF+Str2Jh5MlWBUzWrM1PqyId
eXoOp7WdOc9SovhKnausFpztx7L4l6IyHLMwDXtqoJoJ1/IxEl/0N8FMyiMoc34I
zgtBICUhKlir49x877e13oTt0m9FMoFW2KEcfvlGfY2oR56gWP3cwZmlu30Mt7iJ
oXSeP9BJQFXGbVUw3xTiDeBi1is6EalKmX1em0I+LGLhj/YaU1AEb9JvruYzPtPk
LE8Y6J1w9ehNpBXhdvZb5uskU9nc/hJH8YkD8GrIanLMkFEEduGs1tUfG/CvWhzq
tdlooYAWIsC+hNhMt7gKHcmmnQrlp7NuNSHmnx4CjuPPgCbgb3jbrYU1ZnySpNiY
YPC3z0Vf6GpNRi6qJR1R32snN7UQfA5SOU2SQEx97QDp7EW/cxgnOKjcrf/fXG4/
oWCsxORJO6dG++5jx+g+uoLCCfl8SCy7Tu4MAiYOf92fjfTWSPbsBrs5PeNQgSi/
EbkQB/xIsIuOs/8Vr/2KwlM8KJYl2RlN1j8D8HU9ZE2Jqtn9RtnfIaGtvnLXYDkv
z4SR/RI56bc78yu2UNHRrQv8g+81jgG81jOwVjQ+chKaB2Qs1nPzBGOzv8kQFdGn
GVel2vNlxRBlORqxGFsDfiMp3Hhe8NEV0RMp7amEmAADjEOZtsPRJCR7gD3GehGd
H/Tbfd+VCdDyB1DcaLhHBRGpPkZRhpkF03ZrL3j/oBkyUAo8FIoE5YGVS5OnEJJ2
OIVmCJF95pReBb1/2W5HMWm2xLPxspLQK3YnFN6NfCyRkTm22KHEyNPC9mFAo+hG
nAXydXnU1mii7aev4CRA4Lnre7Tar0gR3NZ99tPZ3RcZ5x46zsXRI409KPUhZE3N
A+JAgixRgGsAQ+VT4YNSvdiX0r3fG7E4HI6mXyz/uWk1zP9ofeieT97ZDVMdhSL+
rxHvSfjI9jOck6tBPVsKmnZtdiekY+TNUQUdVO5Lb5x8NdCleXNw3JfU6RP6OL/3
158Vk64XNLucfG9v+47Bh6CaoovRcgJaph3hmxcTl7/aqFSmVUHJc67+lAYALQjp
it5ySfkewrVy28hlKEMUXH4xRidyNIvA2XKTjM163LU=
`protect END_PROTECTED
