`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yijgQqtigmvxVOciv/IDCPT0iMC+/Bn3sQyXbLAIBPqPibP4XmYAxQk3bD0EMwd2
HaFA2flMnfvxvOhwOBg9zG2RoF6nTlYCaxepWkiggoszVp4vLCG+p9X5I6l9neBc
6sjBI5/lnDnIPcn49D3Gclu7KivioP21pkuk2EzzdOAOhrk3gfSaPDwe2hePTOCr
3ZWJPsyv/L6WiZ88yq9eR8nOE8WL4SkD0+mpfLNHBzVXB+kMmbEmBWVrLmG39faP
QRhPRP56x08HRemOaNP1Xg==
`protect END_PROTECTED
