`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOgA1+CY8RrmDWIeS/T+RoulzAVJbEwSGw9E+twyH6P3ecAjpDWM7bQVc5FSy8pE
HzsWQjd6mHmtP+kxHsk0Mo/Nof7x4A+7ikNfzPC7L+aOU8H02OqqxnYzX3CsNeRd
FSOtuJf8L2iMcJBg308YxaaaLXzXDG7bdFKUCi/ea5bsDDNUsVxBLnuqIRuPFkqf
SHlCX+aitnowE6YrOmmnzQTlLg6BGrdHjNG22/wcHyp9PMhL0ou9D6gsNm7sBp4e
E1nvKvJ4fjlQWV0x+vnJDSKYpcGHPNmS1+UU7mpagicoAg3fOr4aUt8nsJ8IADhe
NVXflydauwak/2C6Hqz9vw==
`protect END_PROTECTED
