library verilog;
use verilog.vl_types.all;
entity IBUFG_LVCMOS2 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUFG_LVCMOS2;
