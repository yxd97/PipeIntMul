`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mveoXt1YyzdEmrLDnUJPBZRvjCPqddUeGXbtJFK2dqaLDvJc/KOs4URc4PWVFCx1
1ZmZ1utazT2XNIMQ6zNUobypcaSpU9WWxoItk10vB3wx8enPZtefQSvgRke04QBQ
Wjhnwwe2w2PLGulBBXvw0/r38nZcJDTP1N79pP0v0Q8jZkFRuDxgsApqEnINt5AV
khMPyNQRmSURYf1Vx2FzWulWknuegrQKT8YnyDvNUVEd50/hrLlo89X9XUoNGX6u
L6eVxMnK4iCmH81Qx4BLcKO1Zg1bTiizvRCIcz44PzD8XPDk9wj1nQeKnmZtqhCR
9VSVTSMlbmSsOYBYLwnuVcnwfTfctoAWWGKpR30tG1vn5xhwRS/AoiL4UhcgeM8V
`protect END_PROTECTED
