`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjFA0soOV4SkzI3RTxYQkHYDr/Ls8v4l+cHK3HbRAVu259mNFKrZTEe620A+DRjz
eR5uBlnen4eHisHN86i/XogvQWoYYNPiviEc6Mf0oKttlLQ5tKq/0gQBs2/XLTas
rPiMTcyHfEncz62LSKEt57LOvSVOXzfsbbyxCTRdnGi8ZEvFE36/RWlIo0A5+SRa
fgewbuOqT7JGvRxrPwKH8EYt0kuIEFMygOrfQa6PB4avmH1YJRHHp0rcX0tHAZs8
5mjPejM/JrVfQPcoT6g1fiRoi38Njqiz5FL0pqGmUkj5577+7GWp4FMfpj96u++J
int6jv9/PVFCrKjpQVEKxlNuZZjKwc+JmGHI97Y4YS6t/zzEQY25KSUonpQ8Houi
PJ668FFOan/mvgfgLLs9VCzHU/nzULbZNN9qqP5iWOPmXP/5k4to7dtMrPy23S34
RrjIGrEYWJjcLF1vnITMGBa3afWq4BuikAr6B70b7TvVyC9x7ixyQ4zY/u3zL4MW
8IMiwk9k4B/azZ6heIR7KRVTSCsL84aK+XBZMx+6oCc7xCEYjc772BS6mXT4YYxy
NY3k8pIwfYX086hHttCL3S3DTC6ZX5YFtmIPAYyZRDTZpB1oJfER7ttn+8rfS1Rd
sH4OWQEl31LrjMYPEvQ2HGeXDz36uLn7kva9VXW/9E/FmPnYamaSkCEv982l8bk/
T76pw2XHg1wQYa6z3aj12MhsZogFw/m94y8S0kUD5edNCuVOJKMTUXfIGgZ8MZ7L
MPG88nRhcg6tt6rnvxM3pP+an7cmGZ3ZCaiJR70yESP2/qAf/t8uhlTWGoz9oYWi
+u9qF4koZNpyHDwVR8N+chv27UNY7UnmiIOEGUXE5OlpyQZz1sAVKfzHpoMy6xnf
//x+VkYKDeiixoeEeB7zFVdY2FXCn7cZQ9plE2KMvc4=
`protect END_PROTECTED
