`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iNOybFBQODGCq3Rj1HEpL5LJx0nawrXr6L4/urFI2PC1MFZHmF5SaWrlSxO0XNl8
mf7Zp9xHUR7it+1VOSMs3zdNKmd0vQBWnsdqn2d3HQRh273HPY/jswYEc480xZZX
3DnPMosPI5BgDHH+7CCcD6JEozZfgRkhySjNjx0MayiB0+2d7/aUjpI+byXGUbGC
mNWvUrF8BjriB3+iwUVell8ieZ0NZ63iAxgnb/lY6KoJZeRuDJBV1EEn8DSOgvqY
cyOdFd+pxdPkNaBOQziVOQ==
`protect END_PROTECTED
