`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+BEC5q2pRJDYS2hB+RGwqBMLI6OHMFMBIc2YmS0y5fPEjrQ0UoIQUYSPPsnth7CL
/9SRuJ4pLCnI5PsN7BYH8d1SdFDikXHDPy4gi0VVjkpSuUUwULiG2maD22s5jAoW
egHgUUIsVXD3uoaIC55EBIWS+QeFvW6JzUz2MV8NNl2Ps0aXOuOcp8xWfFsglMAq
Q/U6nrn2eZJzh1NhcMaq6J55CGV2axuJKJHUJOtcapbkqCZn9OiAQ/1SSrUZEuXb
Ph6jhu4czuteHP55NPLCJ8vrmEl/s2/79ql91m5Feks3Lzw5htWyut9Qy19QzRqK
lHZy0D5bIraRoWihtVVwUvK2Z1lWbv5I37zrs3pDAQ/OSS91f9GuK1i9m+/yiaoE
zoLTY1xW3OItumzDx9eMIYRQZ4efAnx15DixZVVGUWGtrujbEPfpYLR2P4L6hSvF
oKOZ1Q0BBSRRtEWGMGrKyOq7Lecbg2UE+lbzF6mpu45XRnkZHkeQY8+5JOipsUTE
5cx+WYT86Owsp8txbhov8voDpue2i3xgLcc16FSMmfM=
`protect END_PROTECTED
