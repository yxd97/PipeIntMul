`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o2xBPFhIDf/RmQoWPcDusZfieZ1QFus7flPy5HNWom8TzAigCLpkL97Axsiwov7v
raZHnj2Dyse4BPc3SdlU4vgy7763EPsv+Fj5a+mxB8+eC+4K1yTokT6jlyvUVY61
mtn/UC8Ndwre76kk9h1GYcUW9BJ7HD1/VEgCSKq+/jfqbg9Y8uaLu965qI96sWP3
07CME/x1U+qaieN4tkozNZRnpay5ktRvyL5GWEarshFDtYMRHY264/Dv1eBSkRi2
aJTWMJZujuQO4W5HTD7yLUVtEmTDDYDA7GcmXalF6mTqg88EfUd682PyUxf1I/4a
8HHB/PH+GuLqu8Pnpk8SN6W4S4T/+LvVMxTrmoY9uu1MUBG6fEenxblJ8j2XTeDu
ootR9y5D3ONIxY9ZHB6uQBLzUkhqc/cmj47tJrJumNOf5rHBMNFiw8G0/ek1b9jR
vNkyGkOEXrxDMSQ+PSaHidrJDI4vsoA4BoFd6+V7tejm52Vv2ahROtfDp0ziiE9y
`protect END_PROTECTED
