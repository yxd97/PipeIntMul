`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNlGf7anp4+4Kan9+RpnUNcvvWboM/3WoegncqvXpQpSsVAMa4scorgRZVwWbDof
nMKgxz14xbjmougjEoaFwfmFF8Ng2rtowPC3v8SK1J3j3N9jEonF1Ef9aKjupVee
4sanGg3HUAmUiDuchkprCl7FhSxCeiCBfciIhfXAVtKy+hvoeACXtlzyHmV202aI
iIEw7IcHt9CUJmS5Wq9HZko5olj4MEjJRaOrrfIStVk0Z8CfG8GBimTT6YXmFtRw
lN5gf78k/LRAzog9nG+ZOj1ZwAVKvkS5Z/CGRIu7QCkKQgXjO6kz2VjP52+Z/6UG
6c0+gMSKxM42G2MVLoiyPXIeKZfpkapjbANkjOmxAbsuwfjiJf10p6tvW+LxkIJG
`protect END_PROTECTED
