`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ln86L9b12NgDJn0cM8mLP0O7+nJCRDX7i0BDA9Flb7kwpfVDm+ospUT0I6Ht9VOA
Lud4tEFHDH1zObUaIVANsmGtxpk2E+rn3sLkU8TDnSbiItYrVSdmtSBmcYr4emsq
YGhjie1hTbR2i0MH0Cy7A1bw4hi0PjtVQyTgBc8I3UTn4lKCCQWKrqVO8+hGRg47
azU/rflbKyMwEIkrC2PShFcXzhmvmrKmVeQ3anGDbFLEAdI9DSFRX08vmq+g54IO
39NnNj4TJcHZbLgGMFkKjNTKjEFGJGk8xifjsZ7j76RiuV7pGyhO93ODrTy95r/j
aO3ylH23is6n8VgYJoAHCroeHms/Rj8SMjAvHgw7gDAjRM/xR6AXbdLw2dbSu4UD
c0ib5w5MDE837Q4sgx21CSR6rUIc+iXYIu3HiJGQc7MDVPT9bPb97O0atpoi6InA
nxpcGP1igV0uHI+mLQpZy7sj7qpHiOr3USmnQFr1XB8XFGFkGMHEqOB/Jvl379k1
`protect END_PROTECTED
