`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K0OQDyWkiC2BihGM1nvh5bWizZaXMK+BJ7P67xgutrASca2ZV83BiwA0GcWSIwcO
sL8x3D6B2e0Uj9slr8/auh6wkQ+2xh+8HWodZ2T/0AZtI/VXCcj1zvNtqOtB03T4
UPwwgeh+mafcXwvYivKW8x2tzw0Nj8o+dyXV3sa3hmE4YNzG9g7DRRv7sm+ntdlT
HMEVNOjrTjt0NHJCam/OCgd9C/yxncJcukdEGBh/4spcdqumEJxncZ+THR5ZgA0n
WUTd0DWfaT54cqPdB8KGS+QCERW+zFgmpZBHc5yKATRa2CpFA8rPqmDfjWzafhga
c93gXYjyOARQ5wxNY3vAPwTNIi+wAR7mDJlKnUQGGnAUcLBGmfY4SrfsQalNmLmw
GXZTLClfcLxT9xg6+y0ysck1woHZ982Nh5OSxoDs8Wwa6TqBl0/lNYz0ufJWezRZ
`protect END_PROTECTED
