`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7Qmp0b6iPzQ9HUjtZI8n4QoccV6Cn8jUaXBcAyUZp5rV18o/Z0doLtDi2DKzNpP
k69Enn11Anwx4Zn0eChGha45Ww32cnF+FSBM1YP9MU0qsDr29I6dUQKC1bM8RtyW
Gs1bQfQ7D2bHYuGM10GCL1K5t8dchog3nuc8ppb7/xgBVEjEvLuW5QD+7upxmlEc
cddB7+LRJccE7345rDtWO/P2aeUpmP4fMn3rSP9o9aWR8L2SPhj1jN8uHkw1g1pZ
uFd/+4wPZGggRl69CY3pAYkT36sj62nhhVyJluYpJDiTsUsOIPmCfXdZT3dgJh9J
eNG8jfpNNlmNsfNqZqafK5MOa11S1mMH2iQVv2Z2iQaoxPoW2sceaIWj4svbBP9o
SQsGYJYFC8J3tV28YvyMpIQwXJyi9t74hpoUxJ7b6m48KuQm04kSNBojLcQhGCDU
YBeTlkWv3XnETzdoDmEdXAwQAwnE8yWUjZh2LoxZHVnX3jmjzb+iD/pO6Pe8QFn4
XvxbZZecEn6cKTnXaHdOWFbF2zthB0aH+2UTNHxMZZmd7t+DhJYrmHhInqqcQcc/
rckN0H+qh5D5qpi7y3TYGfWAfhGGmzcerls1dKfPr6K/qUGcl6AYm5JkTATtrXPt
lz3mYaiyTFpNpbEbraEZlU5L89yGQsB5APxEMZbAHVfTp3OmNpAc/6R4NxyAvcgr
MVyMuKiHz0zYAe3PksZWBdMWevplYK5OG64a3t15MItnFIMhixiqC1fTV2rdtV1R
sPz6I9uvtb0vLdc9W4vhtzUCHkob5rg3BYdNBMwrSLA35wiKZy07pUm5T1B5/Aad
vDNPRkjSNJwncxfxai68Sz800KGOIlSZUE5r1aGm0Tso4fW5guaA9TOVn1dlNOPn
NyeYklxQI1CJkjLwGc6xa0X6JtGmLHwdqvf9ceTbJcQMM/v3jW1DBmJaqyLo63PN
`protect END_PROTECTED
