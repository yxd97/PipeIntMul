`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cS0Qk2w5lnf36q9W0GP8hP0ybnyFHk56HxZfUjz9X/mPR0XNF+/AxowHcUw2eS4v
Wh2jBTvaSRjcJ5d/JO4w32PC9oCQ/OjsSoAHx9LtezIYxjInxmGzjvoJtlYoWCCT
jAC9QWroA5s1gjKStv1BfNEDrY1OGRoOREtVEGPRmo6yR1AIlxxD4mH7xhmvj7rn
Cml94q+80ku0xeF7SfWFvVkRz2GkOw/3x9lOlmCjKvugvcG8bBMjAY9acmsYTJS4
GggD67wLbQhiMkvPKTS+vpm4V8kGWtwhuqn/yNLSbG4dFHgkeYfBwPKNd65g2Woi
OBJTlogIftSSo13rrfkarTtmGNt7tkG7O9SFJI+yStYUBIeEAwJmTdInva3jdrw4
0ORy1KR2BWYLYr+NPnyXMGzW8J2MUSAU5t48E9sGX2+fGH9BHh2qH7liTM7gf1KU
`protect END_PROTECTED
