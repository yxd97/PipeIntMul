`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uALEgUOl3E8pOZY/1dbzXfOBA/pmF80TTzlW5f83HHN2umERD4BFjXLiemmQ2WQd
EVyvixJ5LuPzZbygNf51LrZ6i+QBz66+i8b84T0BLZToT47OTvHcP+IAZc+TB/qK
/GdmVlPD4hPT3EwrW9Zpm9zcg11Byjsw99/dWR+VdyjYwkJ5EaTDa6ZdNhPm7Tpe
i053GuBw9cJjkpeDuI23GR+9MFqIGq7khxSfsWIr0eRnlCvdM+GXgQdoIZs93Vi+
F+HB3jszXMhp4GD5W/QqG+T95H4JpQVhsC66ZWSP4Asri5Ou9rn7+Fyrzb5Rc9Jn
zEqb9RBn8Gb95laLSyqT1f9pfLapx3xjF733elJa4RDbv2xMLIIUbJN0O5zqHGbF
6wh42eFjfYFvkfOYSDvAXuU9x9oy1NaStlbjG2dvmvJv96vU3flobvpFWaPzj4T3
ltInzqwySa6Vt7P6nCx6PAkYcbM7rQVcHRdPoK7r8bcBE2ZkkHfoMH6aVg+THR8Y
KNYsTL6d6QKxEJrEm+/ztVG3tAGIJRaOsoBOyXAVjdFpoE59Xk+e8AKVLU0Gz/8A
GuMkUFiCSNWk+E90tHaiZLdgM6EadourmTFxrLomGhvMvzwL7SdWdfteFL+rkVDo
xigj5WTPEbaKpC61Y3eFTGTufLFR4NxlINRNVb2qKOOj0x4IT8jrvnm59/4DvNIV
PeZmD+fegyyARflq6rkDjzjYZIG5QN1O49LWGFbtpRnTM0xcrU4lCC3ht4srxR+8
WYlkotxsLld7iF04xdA9/pfMpormh2X4bV1PUPuwpjVLIVQe1m+A7/OWvHksmY5U
WZ+nMMPYna9e1hOCr9dcYOqld3yxvTIckktjqCL0sKOAfa3Hts8IffhmPMQ/VR1i
ytGmWt64ynZ6N070nUvbnzNA9hwmJtS1jeIC35GiExf3APtm/U1N05soelblCPjV
sNhsiG+CbwFtq5jndxQ1boTcmWg9wgOUXeeThMmCavpOO2i0VsKZb3nOfb4No+2U
lMezQX4NZbvKwuwEGsiO98t3twhY//1DapluyzNMMvl82TVUZQMu2Sf/Aw8Xyffv
toa7xquhbXB6eYp1cKuToFOM63xwDeWQYOVYfmFgFkf/DbnqGy+wTQBXpZmE5lYS
VS14QDuj/rGhfKBLH1qGfSo9tH3pR+rcNz8BRxzEPPpQvFrPcEEMbzB/stwHIe1l
WcuXZqOMWaTs31oBRrFdheU9/aRhI1Iy64ul5ir1rRH8Hq/z4xn2mushcL081kjS
/pluwRqVza3VvK7Hthf+vzuNyF/vTKikbDz3P6E7s83J1XdJFzkanBtuJf8spRie
r/mR7wL+oYxyB6qso4wgp+ENRE2HympN9tqqS8cDAxKgXjQIH+VprxGI8RF3931y
pBGAXeLCfWAGEOfkSPKKhfjJjKj4eWYMtehm30OJun8xiC+Og3BHQwKveFlPo1Fk
B8E02y/4hb1TwY9jrxtSomspqlMwupmoN8Bg0ytf43617RDb3JDqmqsWjerNnuTp
lUhxWSsHhSGCHWw/jbjNfZKiY3cUurB8rNMi7Lbv2V4p07OdYqn9sTDqf/8fUhkJ
zpDpdVYlRkWuQUgDJNL6xcmd4Ih7cZsWV+3aEqLKCkDJ9AnXYsVrbpp1IKCw2eiG
91DRXrSUC1ATmsc/in8XLVhEopVU1X4EuOiX5y8bRdqbWDcEHfrDs5jxpUYZPiKh
t1eyR0bQMA48KLX1Bz5uSPkL4CcVQzGz29D6QcS8BkUDcpI+tUJdRGh3B8CCz235
reN/6ZGMd3yn3Eg8os004xlT25EWKxw12sGqCtrjBAdso8x12ls3uFHNqFV6dtfT
317TjZLCKGlK+wGBRF8AixbHcRY0GsdVz3dJhs11Nr+oKW6PsyxnLqIkpVX9rouU
zrqfW2RBm6Pw1CGgeXsOJI6V9z4aACqfp79M+WM2GfxeuEnlvs1Qobs92vJyoXHi
VOij537aku8VxQfdGvu/RASU09rKYiyLbFsffip1kpT7lCHc3Hdna79UeKBHTVHx
NRHb0P/40x6IISVAnsUll7bQoYFr2KIZV/WWT30o07tWeuXgvENyBxM12NhtVb8V
K0+7cEGcWrIdyvl2WJAN7/JGa22eTJZXIAkSAvdzFyez81ek46x4/PU8kNPTAMOi
1vQZgcsgQ1ug7QSnCKBGwjQTGtzCnx+0DPpg7+8bEfQ9qsswkglu0Fu+8Wyf+/E+
PaHRuhUUoXMHoWwncQwdtqbBY5Sos5T2tgZ0+s19nlxY6BcO11Z86Hf9rS5Ipdu0
3wVOw26qtGfQ46hBtLcGpd0GVW3JUASgNJhMgKxtgaI80fIZEeznHypQPjhPkLU8
zuARDJoM/8HRy6wf5hB/ihNEX7u4XLrHBD1bEoLWmi8ctXsW5MVNjLI/o7y3lnvz
wmW7gb8pqLOgIzF3y2BEsPnTCczjPfL69CD1axWqhOt4kuZmpSpA8qgu9mD657jW
ttQl0B1bHQzf4B9dvxwaC02sWWbhOySbi4gYIbXhm2CE5xIn5MjSXqFat5aEiaA6
ahdh8rdslJVocQIqGyM+JHC/54PS+JCYSwI8sToTgLuxISMIg7t3KHyyOrtcWFNw
fQOD3ldvOEZsXMfRVyJ+HhZZAbYJuC2J9fwSITJACPjQ+Hf9RbP0LcjZRu/298CQ
9nwt7j3V7fyIUs78RTEGEL/Es0Jn0pAI7zfNj0OJAnc3dkf7pCiAExsrRLvzvrfk
kiKayAUEv9zLELA0CLZWp6ULkzl011IgwtMe8qxMlnVd77FEqsmMdIHrWFB41CUc
vbVhcJkOdPKZXFSC02sfR1GLqR7r5aqFnMhQ4fsL9rR9GqPoWkqcgCtxLsAPvitv
/gCmvo7d3fpY1iIbp/P2x+v6tQQ8OiugUvJriN8TL+2eL4ZVX/IQRk7OLqFgHqqt
7i+g7itl/wpYW3IZTf3p7oATvb/DEisHCy7gxeh2Y1vcZce46KH1U/YE3FzouSEu
nKWRsHwahCWc7+a5T89f/DqgzCKtds4+eSMOTXAzuvp5lbg6qFTiMDqLiJpkcxth
i8BgJCWGauUg5TO/0ktUoRlQc9Ib7l+5ruTQ87JrxWro+b7BGcP4qkUOVLQ0D/VW
pFDUw1e3eit0KgLWMYHjBg06YbcSBZgDaG1pcY5dOEZaouKT5uDRiA3h/bM6YcJq
MxUzoS+25kabma1S0fWPvl8liYKYI/AxsCe/OBAmyURLFTx03bAWQvMUx7boCwJy
fXhMyxA/ts3cTRCVOXLeUAgJJ4S8/wZ4Wwqzce5Objv2ne+R3pp5uedUd1nxSJzz
RHxROquuqGntgFxy8m0b64yy7nXWJ2IxqcvXWoGJCDiq13J18wh8+dPXy5VQzVWx
rtcdm+vuf9uqbpHhdqYkUhEgMNPml+BrnN6xpC9W+3Cd13Rf/mqAq2uiCD4lnlYq
Jx9lWQwyi9vTGvjATeg7F93/l4Xe7dHg8TcBGVxU90PFq96a/UTDXaa5/TRupNyQ
QFWBjUqK8T+hYVXGXaZ4aRlBOArzWw0k8JayEi99lix8U2FmsYMJVph2XWzJBRtK
CDv02Og5XThapqMCgiH6GLLqHaWPgysQrrDDYx0iRRMRslcL6sOSZD3zWgdyTuhB
QRAdshh+XyDOeUv6OhF8svRHc1AuQDFt+4eelAXgEuhWidk6nonz/fEyboWdQrVK
vATdwgnn7Yyl11TA4Io1rCYtpht+SNCgZ++Ao2Rf/hxiWc4TMUySsB59yHBLppxc
EkDC2PpR8A0BvBqkNHvr0MVKlnFLnQ7AocPShFSSYiRUKRiE/eP6mQZPgXkpN2a6
ys15KpA29PU8IvRBvOW5yU6Webo4LGBTEnPoKh87f/EaHhzPdZ4Lrx35+MiG2TIR
BlS0tfyKKskJv/noYX5k7GOKFELTZFZASkbtOmKaIGGs0yLKE3X3fGyz/IzxPJ/W
oYHl1wkScpjy2Qqsu8A+GDaNtbuwlL0Aossnbx3+bZSzxYi4LLoWW1caLUVUBlTb
VEg6dpuGK2N3SnVgL7IPuEad/WtuHXD/mBL3L6qx5dnrBD9RPU+kdq5Ea2nbhW2L
cDt/U0gL0ZwYapMaU29uYc4t/7bE3XqtRGWqoc4DIRRNFKkBzNw3BRo/eTuSNF8r
ygBV6hyLcEVtF69uhQ6e/7g/IEDxf8K8ro7VsGYp6Wt1BNCyJvxRIf8lqkzL+2J2
ekSu1vJQQVUJOU8LWgJZ089UFrEF0B6NHxNgYbkuKtauEpuX7qwNdpFur8aMd02t
i5v9chX8GxfUuOxU8NBbZ5fHRlZG0jtQtUKkMO7RSN02lSkpj5ht5wXg2B+Tv3i+
3d8bHKn1GXSdDLlZGKDw4FjK5Kfop4uw86TAaMjqKD/YnrTiU1jM/itlZ/VT+PDs
6rgbmE7FvX6HrQWfOWOziRZ3GMqDikfX9exZdKsS83DxhhMFBkSQ5JHuWa9LruTj
2fdLVxoAcYz1LusCG9kvqNFHYcgZAaUbeMsm8LP/jKTNMWR9EPbTYZ6pXpERxkRz
Om9As+CfKTJqzhSvQpI03s2yIBWgJFaiLa1jJEW5Qih1Mvwj/noQvLJqfDxYpY8L
vmvgiEeg1n+3zo1C46amlJmDVndGFLY7D5jg0sKSAwQsVJ+KTPuT0RY8VY8VkimR
eOs4TooVib17SRziaTvDgFTabEW1XBPyW9E5gaqivCNdi3kfGQdqMxKz+9abSmfl
uauEiI1QB/QSOh8H9ONBjjEkorZY2SwTrV3nB5LywwnnbzES9WqL5L+M+qta0ISb
yQaqXs1syU329KmvklwjVVa2aQi/muFlJMT3wKyR4/Xfj1oZx+weSdtunCKfnXU/
FwXNQ8EW7vHWPNPSdGPEmHlqTqdE2N9vxxXOpR2CiG/2aa8B7Nqa9UMeYat0LEwy
5jtHwQ7RsMtU7vs8Wr1IjIBCz+45Xxxipn7IManzNrboBgKnk8k7B1KXeOhiifY0
f5pt82f3oyxaaVU3zXhQB03ESrHRMwu6OLMeMP7Ww6k7gD1o++ZktGDk5sF92Kcb
6F7/cGPyf8xQ5k7IFjQ/TvmNtLdA/gqkoO2W86gnAIYsi9+ezUd9pK3rdkaU+Xgb
xI1zUzZ6w6//WbD3FLi62KpzVFBuIwVNvYynVhM2Ho7NOFJuU2691eq/ms2N1yre
RKZvvniNfSh3ACQA/n8S7z/R2XXCbngeEC2JSL3xBiBALlmBh3vogG4iTkCCZbOm
A/otzoOfTkWmJ848/I2jXoXl8r5tAyFnBsp69X+OzZtgB5siaxqH0eUCJUe6RsgK
tzlKm7aJcM4ubdkmlwB4QIX2T4VaqM/A8TgP8wGTf7tbZc6kgDyeO9jXNvDudbDQ
AF716/nDXnZ8ufu3/an2ElrQa96sqdgbKCs3m9uO/Rqxpqbw56YTcYO2QP0LJOXF
CelltQEFfznbmJAzRNei1WROpbh6RAcsTEzGO43umXoKUGkIaVB1zO+FcyBXmHZ5
a6vKNEdN/+J5eoIatuAqJTZcKoZvCPR0Mo3fHXNuZ9Vr+pUyrpZX4hdZ/WQWjCC+
EwYEJj4DPcuNrZz+CqpOVUHTrGo0HcDmvxTTHXOL02UyKOvPEY5RZemJUcLMSBEG
0XhvDBfgTUsSnkK040ZsdazZjaWL0H5ry731iOuB/aLk+YXt8dPC8YEqnWOocVPr
hCoAiKuAMrFnAzqCt1A/QFDWdazO3aXgaS1kqz8oKlHYdVc8+8rlIzD0U2Ih2VSt
yqJu7Boo9XlO+AZtXkqHMUeIHNeYzLJIQ911jSycktmapB3+gIIKVRdWQaTadeF+
1/bE9PmYWoTnZCV3Z+ykJTVboN+xGjs9kSRchmjfEchrzFxW/u975ybCF0fqkGgs
HwNj9/uZd/E0uX64aAVLZBLkZchHE1rfyj+71lsmku1KouTxkgSX76w+4HN9yUTR
QTlnv1eVwYvSHexFNZnmSTqwCci8Muo2m6s/Uq+E3fx4vzSaYyvuE212tgScdA7f
2Ge1eut1K5LCnqPKISDSA0aa0+qliEQhJjsDLkz9yDCwmr1dM2PE8AkKl++hCLfR
lcDPm2oT+I7HIan1QnwWZAUUhqaaz6ceyRc5nRCmk9QBTfAysCoJve+rzR3O8+Qi
9MsQ1pqgvohF6mvPHnuLtp5HA9A5LaV2Hezphc5fhcun62VHhAndktBQwHWMo3TR
NaKLaPv8bp4+5d2qHNtBEnbhG2uuZl6ya1wpyuGTk2tmEUbVa6sHD4Xje8j2l2dk
fAzU19iYVmT19+G3PjknWTPSwMNbCQpSLdrxstD9zA6hQ9yCFhwcRYtd8VbG7vCA
1EsovU1YOxYvVkWisBMA469cC5hLIhgqc0vJAu7WVVo9Hrlg59of41/vW4R9lBci
1IM8d7Q/Kcx+ZEBSdh/cLVrqT2udAJAmvho9M+DfRd75ARzfuftZc+JbVUqe4zF8
98HGBGDcGjaQrS9SQFkAjwQKjs3yMj+qswypX5oAyfEChRKRyaKU5xNGk8k1td2q
eUa9ySg/XmrDlyIhwR/tKH3Uf1w3pABRc4XSWr5MnEmRUiuq4ehHQs8h4VK4dCq9
rq3lLWb8FQ7yuN8pPzlUILoHuruimskGlLaPGWZIrEIg5H1ldd088GitZrkzKRhI
aCf4SxD5/F/qOtldVWfUf06jUagKiVy4G2yMNq4VxbVSWtnKKl9LarhN5rfiI0Fd
8pwI7qirJq2XThQ1XumVfdl3EA5kbkOmpMKvvQOxfdgdaDlmQA51a/K0tB7C5tWv
nofdUuHFnb8yFCSHFD8nzdrcms2K2nmmJlINCrRUHHaGQiUT0o3pok7noBxp0E0o
FF/njaCfxtDUT/Mkxd/KelloWWDXRrA/ikUPr1TP20e6R/JcIdRoGdy6Jgj9g1HO
r2E0XXLsBIIaWtEYwzSarX0qNAMF025E4+rUZ25E4z43J70MEbdd8J88mQlNzu/p
EqtOqLv2+oBgsF9YhKNFHtLhbD/Wg2D2KZCuTEdy5RR10aa7UagqAlou09FGaxF/
XAGpmTMLupIjeWMgaea+Ui1C0FRdles49/+MkyaGzOJrbybYAhb1GiOxBcA1dGcX
zVj5UY8law8S1EWv7zCLtoT8deisXybp81Lj4Y9Ep8qxbbvdiki3laP1TTQliD/A
aBHoFd7Q4Q8T2YUYDhe7LBvxlpl1VKfjz/nSYFpl90zong4kG12Uc/m69RjX8rs6
qIvZhkNVA6l2PtB1YAT6FVUTnLih7w94pEaCBJ8Sp3TrwDPl1/1z+2QGyY5mDTyP
9JKFrxJD2Fs8QKQrGqtseIWMhxjKCp1uJoIhNVhCLr4GttPDUmITn8sueSKluwEJ
yh5lM11qV9o8KFSgoIJ+vV21m+sJOxj91JeB67KyEX49ED4b8v9z4ZQt5rnwJoK0
js9OGruFo+HS/u1ugkL9cO2STvsR6bzfP2IDXMw2ARzd8JVakCy14CgB7ZRfv6Ca
H53B70o1dA+fQ8sXdb5MTwB/8iKHNONtBJMq/llt+isaDUDt62lQ3TIX3qcX6ZMp
4yeDvlGPH5JDVMM02X3sH56qiGoD3tneTM5JArthB9BngzUGbEj+n9sdQeorUNy7
x/7V+0D3KZolJXydUnJinhfAiOG6Fu2cCgLpLmcdDdXy2ySNO53qRBdqeW43ccHB
5kAf/FPQrz3K6XV+7fVPItSNxLmS4ReqIwCdo/d6UOQidR/qMXhL0l6Idq65jj6g
WRV16sPWwoO3G8G+a/nOUrVfI5hoo6CiO4oyiiWBoThKRbQKHvC9xCOZ/NET6Dei
kLXIqJY8sOQD4DIi+w0OzyyeWR49wpHmzW48krH4Q7Kjw1EiVBIjPhQU6O8CJhAb
7ksObHR0F/DlTTcdu2IG4V7Zba6FT+yaQytrsdfT7O73aCBjh8ILEtmJxK5pJ5rQ
3BdiNPBi2ABZGP9bvOKl9gLoF9mql+mRllF5dQAe3oZzcRTpXlm1ZZAxDq82AGjk
tIVa0iivRHLW9Gpc7dsHBlyixuAztjRr/hQLHDZ3AvZf02LfemOPU4yt7P7YrM+r
7i5jtVZxeMq4Eb3sQIl/2f7rR+jb9fFd59rQGXnLEqGneBiMfey6/awciL0QJLaB
sMdn0sCVgdSkr8CtmENGF8aZKpWDkO1cfjzKbO2p+biM4LPI84np4DS6u9h4kufx
lvKa8Tw8SbYHWAkyHWz+CI0dTR0T3hEPe7bAyUyvF/abEUyJhEglsJY9EBqA7exE
8OYTQEoe+zQUyMaJklNlY2L5h3jSU1aiqVsjrFlxt9r6Nx0CLTyN/4DWx9o4X7xw
+HpHALG7jKxBzW/e7ggDbzTae22C5n99W/PDl2uT2yu2gzhAzqMfGZRcr9LbRoL9
XCgWDeMDa4XwzlJL47nToT8ISLi2PMVEl/0M37q0zQ2SDwP/K8DnclxgdQu2Q6Ng
A9bRO6RWBYmNsVV+FmHmXlFm9qTUZ7/lJ29Nk5ngHSCCVxxX8tqPwR6cjg9K/F1N
7kQGecp0RLy4XLLHfIZYiHKnacfVBNhN4mHemEXlXGK9a3g7gNGQQaIfVThWyn28
RJgiyQIQWz163BS9w96ez0ZyaACgJF8lfbqPANkHsr0EmmGSdqxLwm4RRSxX6zGl
8i7oi3ROMK8acUbHV0sf11mCX+6gFoe0QWGWCX3N9SDBdZAGcwvKZS8eDMWVEac5
VPhjoroj6XLVs9mERPTClC2HcQnRqSK6OSp8m2ldG3FkM1665MA10Tq2XHHpT4ov
4NAdONqCMPQUX5GrdAomFPc4qZfoJUpx75Ty7XWHWtHOKwPK5UNCMQQW4u+F3NR0
MfEpg+y+vE1x1cgkYCB4+zeroTa/iBdvVIWnTPN3Sg16INZIXr8z3Z7/LiKXI33e
mkyE1dyENvmhqh7JE+RnRKtnNY3ROagtVH2hzuqNaD12snZp1wVBQ36/w6r41Ifq
Sr4swzlp6OXOakaLSSewyJKLuilCfYjYpBL7vQCcJlITDSUIVtMgHHRc+JT45k5x
mc8izuWcT8XWo20RzrtnGYDOSrFNqBDIqpYXY/VJElGwj/0i1Qf4ypxDOhzsWrrP
JAhpn/lrswM5By+lGh43QTV8YMORPLHDY7dt89E2imTMmIcC4xVXBi+ebFUr6tKy
feZBRs6gXIqsKMpzrrpH/dlDESNixrOmOiXo6dY8w2TY94Dv4drccqC4fFeUGUZo
Z4VmxIopm9A9O12mTex9zZ46ZjffaRaku7CQuYNdG3t1PhIMN95MHrwo54ZlkkQu
7Ahyod26wphA+RWYA/KnpkBvuAXS0ledvzzOXjGza8IMs2fN6BWS5mrDHMN+srPT
ZfuSCoVoGGQ9SwjvzJgIv6F7sP9v+O0jlo5hdA6T4OZDM9P5CPpGqpUKhzRAG8GC
eZKmtlUuhTvIlCrjOH/Bnia4iNObMyAIBPzS4Qvc4jCGUO87GCmmy/qdQ3Hy4nwj
Nh7jb5sDdtbe+ZIwKu64ycJAdnMT6MKCoUL806yM7nkUw1J61hQZYdN97NHuDAIL
6waVrhDTJfG0FsXpB37YbqAzYI19nAUJ1KK99jspvFNpEeucTGG+pHq+R77bm1vL
dea1iiD2tRMSLpodJGmN9TWo8WMSe92mtd2/KpzHcWLnOluPUUsSCOit6eTVmeII
PuCtKAi8ksi9BRDgXTcfQ3iuity9B0JlQhypP1hCjNqoWzWD058JV6n7I3X6jq8R
ZWBkIiBCY5t5WH1S/tuPSlqfXS1VuAL2b+66n05ua4m4nc39iq3kzt8ZpH05q4WH
mmkvizJNYV8fGbkIaIEJBwruskY8KHeUK4PWFoi8zhPezx2zBpBd7LzlSlEpaxkB
ZcxFJgdine/LQrOkPf/nYWGCuy/EzAcZ7XEw0liGNn77X4V89gxSsBWQ/P1RLxjz
l34Ru0agVsduvlRt/H42zv7Dh1XIWpPc418QJib8tVIO/SdalqnXvNjLQpzKcIIG
maUHtAjP5pDxTgRjGEFkUXj0m1h3a+rPat/C/Rbxgqye8FpmJYhxAlM4y08pjv/j
6i1nHQSEivvtOXl41iOwZNouxHFEpF67DXjWjuZSg4IatmUqG4q9MzgHTQiPMClq
yTj45j0EahWbml4FvJIORzWG7mjLFltkZvl4c2kKKTwpSVTNkOa8WB2ioPRdB+u5
UQlCBRyinptX/+mu8dDwyzzHHQ39ZbehMsOuVr4api0efSZhqhksMnstttgFsv4/
ATNaj2GpScP5FrAvoX7qb2OWS9bo8O+JvoDAVr/jQQ6SK7Wvg2RU4uxejEcXKbg1
/G/MDkFsmQc0JIX5h6ew1VO2QvAN64GNKrVSU8WEcY5bKCBsDNiPK251CXSLLtzC
TWlzXsbcJ8vA9ewZTxsDhP+fboIA2gEBsoRI3wWG0cKx7x3LZEea0GUb8rTLj9gx
xVu3RDoxJdCwBOQ5Qmwf50w/Mn+ApAbx2HBqZ1gMSRPm77cW++ePVLMuVtufUyvh
gnKefzceC8o2RU1ZQb0Czw9pnSyZb6AqPxFhilaMgbgb87mkWvxH3K3h6gQ1XwJR
6BeMSV6lu88kxJX5AaZ9gEebc7LEaKh0o1qvbYP3vA2jNQBpQscFRRWoaT2R9F3F
sKrSklaNlwGg/la8cAER1b0jxdo8xBTpLm1jIUAUqGQmvyQ82N0+RvF3flFzj1OY
QlmNB/sgMYfs9FUtpzEzHpFqIj2INal4yJR4pOj5EuRXe3IRtg9rX7AzsG/OtBGK
okBKgHS1C6UDmu9AV2lM4ZfzxXddzH61es+Zo6F9GSZSds/iEjgIrKHRL/UVFmuV
AyruxDgkKHxDftIeaRRC0wBKQKDL4M4qilnWsOxaF8FAkhJcgWNGB1tDy+xJQ0Qg
jbp7859cX50yzos/tGjNjgT0qcGOUbdlhQr3Wx/08ATlS1Alh++mcXYUrVmYA3cf
uSF06QEH5oN3BRY1L1AIs9IrdS9SxxXbHj6HlL8nfdMh1HbjY2jlmxzTHbUpk0vZ
EVqpRMNP/LnYPWFPeA2SRClnxlsgugHxCxJQjifxDYeY1W4ItehOGo9ygT0plQwk
D2oWVPDFjdM515bHeSx+FNs8UDXizkXxITMg+5yrA3h/JE4BfHq26nkpFrRYYDaK
sFG7m+auYszMcDdcyYTnhWQj2P1WFyezqZaRtAjLYgDudtDO6KoWwg2t//2il8Jy
GjSjd6JpahfciC5+IAhRJqknJsZhpmem+KYFLWyFg39uR1KG1hrrz4I6aXn5HC97
r58XIjRhFuydV234RyZ665QLIAubKYsYgSyFw9Jab9VM92gwoG5ZWJOh0o7tUkQ6
KmfYZfw5Un+vugE/R6vZHQKOh9ihHjU4X19OPt3KYbPY6JFyHh5dDT4+G80rm8CX
Ze2y/vwQ2xxvkZwskYLqKt48pslz+QBMOZWoVaXMpMjjr9zh1E9ccTkC8hO9Hsrk
tfdDENoCu8Ns1FClG8FkAvvx1yrDjQ9004pXiLfkkAplyrqI9txM8vkj1pxriqrR
ychV1qA+tfqGV+7TU6fMnG2o0vQI4keJ2KZlLp3fPRRaip6dZGHfB6AAiijLiZjw
EUI4VFPWuaN8y51WdihMbNc3zSaarRjkty00Pa9MmoaYFCw8nyCSvaBRDaR73X4u
p5ory+TyMHbU59BB85qFJ1x4FC5HeQeVsyMj2au2Iag5nhWj2an/3TvCYjA7jcL7
DuPGLdc1KSACC1R+gkyq3H8OMBUXdZsG8eoyFVUKoVMd2bVbaTHobHiRZG5m54BR
QbQoxDEV9iogK6wAOuOWHtxbskwZ/oE50aOZebGqoPMJ4uVeyLQPD4P+OQY0zA2x
Y4MW+CP/8Gy5ZCt9dAlB7IotCgXNRD3oW6IYhU0U1gdw3MAhu3KzByCqoxf0Qfsm
8q8syE2o/lfIO5VXVGXvSxb7ECSncmvaHS4H2m2xCl5rgHlXbneYoYMmebjBipBv
AM23tTqrKPwSvo3lhdFFcd1JHeMxz2B7PizwTgxmRm83i9hWWITSO/VMjQ8uYGvU
g0To8qEuaBXE//4QAb+H1DnF2Nd4Mq3WArhr5+KDHWaQCVLk3eKaLQRRtiGKE4P5
8HrXlgNZMqo76eTDUKfNgd1j3/ucgWRQgfukU1mQKjcUfgTcfh8IPD61y1jSwD5a
GOnJwG2ipsiMGGQUxf0CjrqOpOGbl0BueXkUfMIjosEMCdVUM9Upd4dQ1il18rDZ
WPrfUFtLHwCvcoFOHJsMda5GPQcyEwnQR3b8KzNFhuA0d9qnlYYQT2vWJvayUMK+
RrUtS1X2Vmc6+72gccnqie8xqdfhctAZTe83zV2C+u122y96qWO0ZVpBaicqhYCo
j6Fp+K7yt69oymBV7j8dugMydUdSIHIMgmmTKzp59Bza02jFduy1+e2gldfTNdA4
CsHnfemlVYtUgfK2NDCXPqtx7Vta5w/9QNzgbNZmiz43JfVCzohlNVk50785B5q0
3XiqoL25Q71rFwObRD+D5goFIY5h6OrkaqkB9P2QonxkN4wJou121WsbByPkx2vp
wHIsf4X5jwK3ACdKAvlv0FeKHr+a2+dGgacDnSZdM+TusIrjUlsWf/0wUjoJP6OU
L/uoZDfYswbFBSDfxnZzmLcfCfoi98CjY4SNGWXzysIeZHtC93mALuok0xGaOvMR
GmUyWLRmJCmFa+2m2AxNVtLRn3tAOmGavn6QEB3HlRlgrCIFh0W9jHCwuKNjgepT
ssEnjTmJMPf06gPcKb7vjOaegq/mNZ886WkEsnHIetUeCrwUa6FrUkMQcROkfztw
0qEUVu+6fPvI6KmThgoH28PPGtHtt0NvtgH8r+cYB1xDjrhu9waXy8OqXzw1qggi
x5QquJxBGssNWRKKE9oHpflOu4O/JxipWwYupM0WJHiF3F4QifAaw8rdlvbFB7Mr
YIR7WZPJAzq4erZTl6/WB6C/abHT3VQzL6Zr91Qwh9UTa8SRbKg8/KU7EweQWcuY
5IoTnfZ14405C/wwZ5KcmMISdAqyS5lD7WJ/J+Lnk2XKTNRglMK9fGBdcpnHKoLj
BA7F6qANrQ4FrK6cZALLvIKP95wclZra8P3HTZ9O7YAydcXS5oLGU375ClO0GjlB
k132MWIPS+MJPuYAHL/+Td/skd7ZYa2rRAkx2lbmo9ZPbARi/UEjj4eYyhNvxWOd
Rc098+alWFCNWTZpsFBx3CzUihVAHt3uVwB8EpUDd2ndke3jFcoEBqmx82QqRCl7
rl4Boy+U/LeS1sBZMOBGv6Ce90AuodZ+7Eq2jeP6FubT+oThNevisz/hJsf70WV9
zokkFWFINm4nkBDLB4bZhwTl5er5T5AKnDZhS0sOwk/mXu9YmWPiCiLMLzwoxU2c
RaVULp/zMGTA0nqMXT9nG3ttTmT0chfP5AdtjfYi+oS1wBeI3hJuZKwvmvuIScms
9Wlv8+Jm6GZjCSKd2H+Mu/b7gm2wpbpFZJlmQOzS6so/6Nh62iUAyaBN0Va5WyTH
c5AjXk+Kxbdsz8fSwV1NxSzldbixz2ecVuwLLrq37a3ALbSuTyCFYbA60fAJlmgJ
Ws+rWH4Tqvn8D6aNg4MndeV83UaiSLnIcb/iJiZG40eDawBI5bLUOnrKJmnGMR1b
rNrdr1tMdfh/+K89uzWaVgW642+H7BabviE7BsqJuvbY1lnBW/zxs4xBbDbw6bNZ
p1Qy7r8/2BDnvJ16gEks9Sk2hBEj7+ph7T/Bgbt98tnvLAPWvCs1gvHvRojrt1s5
SNITmLB/O2NN6ylULSLTOztyQpze4/lSDwbTH12bXIylDejVBFT3U7CeXVDeFRFY
SDFsM2U/ftMmB7KPegdjxeCaL19uBZSnmXIXv231kyyzulQNdtWavalWiid57oJa
E6v0GOGwcQlXKyluQRYWxLRuwDqdiC7S+xyIVVMcRK5eA8/dhD+FvbS9TKZMVdpl
3P1fQsoWm9zUSQjnyzQncCm6jXoGm4t9YTqC/WOQKOCrrZOu3fktGvpVfhmWr9LQ
nUKlsaaZnbcg28VJ2RC7Jwnk6stRe+7RzwqxZJNjtn6whPAFmv6AtauDm6U7kHLF
lIqN3H6orEMEqlgwdI8OnOFVIuigjXZ468PVURFc59HUeoeBWbH/kLX09LpKv1z/
Cv9+OwY6Fv/dzOGWWS3JYAkuHtbz/YbQp12/qVrA0gQ6goAVkEOoXGVR42w6UMQC
TyA8rpM9kMr678z9vYTSUPz0/EwMV0BVjARYI6lFaYnT/dpJ/RSb+6/aP+HBuly5
r7LIk+rfzHl5CiXXJTnaLeWFTPhN1mxOG0TxOJYzxWajHeStzT/XjzQp3aZMcaY1
rE//Fvf/S8rmXtnCO7+aMY6psUS3dafyhBQ7MPOHh1a2WLUZX5Dwltre8zPLwi1O
Bp7wVgGZRFcnF5/9nDELx7lOARLlW4qAmVBRQPOc5crngNTPDmCyUJZECteMrK5L
cEuL6z6FKEvpsyNjfL3VtMOv8nzw1eB0MDKjjcgnQGeYuL0vfhdxE7clt70JWq3T
NcJqEtoU14Xbc4gq5op+KUghbdFW+l/DcbIwqPGK7it77Fe2q4SKZXzbgHjsHrGc
HFQNVRq8DEd/j2PjOKkG6dMiOBWBIM5Z208vUkFBhwpjDRDDmy/2IMamqWVk3gm/
XNbhMcfkDw76zGFk+9hp57PwEWqxeQ3Nkgjd+y5oijzy96bVCpip5xMFif8dTL7T
f1AiFalJ1iIYhKI+HC5v/etScEs2wiOL8Iig+ALTnlryL5hO+3U/zxpM8s3nYf08
0NZVjKolIPNZDYwJdA3NOS3NvEknB1icabShMUnasBGYL61Yosnicjtlq7ydZcmk
kkFduYZagOXBdDbAq8Iv8sSIoGlmu6CCaTe8gawl69tfdX7rUj9DYTxQ35l3py4S
t084/LUj/wb4TKLds+gwO3Fa6uml0nGJVCE3IRFSfn8hSnPk9sUh1gW2FwFDIT0V
Mcs+q+2bn97RVXDqqY5tYfnoFAn0+pOUrMRaaT+2Uoiza8MfrSyyXr3RwEz2sNs9
zEhWwBi0T3hnPx8K4yKLnHZDnCEiQvIrMJxUoPKbcmZINrfLbRL2eUqe9+GiKHfa
LmhPYGKeTyIo6H+Hhtk1rIm1zq68iZVWK1/Ty9hPdOcbnbezMM2cpHrGUQuoYXp8
NEeIO06GPcVytH6y/ZalSHigqHwSKjfd5ElnZ47UXAvYQyUPbQzYa9NiOveYsaYP
GUH1ekE/o9tznQZ764AMx83fbam8Mw0b3m+gPb3Vk0bEG+iuOfZWVSpdUtIGdBTq
sFdesgTYmCHGuyPsKnlgCj6vbcAVDwp0hByX9aVi/lMdJU/r8pmhMZ8NLGLhAsc4
jZVTFWd72Z30yMOzrjPR4PcfZFYDl8/m5j0TGHwkm+TdMpdU75vA6PKEKcnoWIOU
H8OJegCXlwpOz+0qlMq53IOLg5wwWm8GA9OGnwsYGgvaFI3FyfRsGDgmknxDvpKL
mW1/iosZRv6UgClUsW3mkd8v+MRYOV3WgZb4rbkK+iHy0f4qxgVG8+ZtJ2fgw46A
P6qI7IaPpONAKO4YvsfUbpDj4Gxid1U/RAqRFAX6zbsosdg5YiQOW1YoXtM5sduX
H/Dg4ZsmjsTf5oRzoskqnwjYKaKTuM2/EI4r1TG6RPOY855Pf78+Z2ftVIxwFvnY
jkSoPG9zPNW6nmLTjdN2+CRkTqWUtR6hL34yWVW/408BkKqW8GUdYZmYML7m5YwB
ivVwdcVwGLap3ctCBTESmhs90KVLUf0hK0OBN5pHLFweTsmUijA7Q3e8ll3A3GIm
nHbnCabvlCDJ1j1utkTJxCf7neFwV6C8ByT7BMnjw1LR+H0AZfwUwZPa/XN4Wktz
yRgIm2QKWjT53hjO6CDC4UGTs9ywmMt6sQxRQQfU9nFcyDqTb8uUQlAPHyWruAUI
hXHmybL+SSdnCMjlaJxRJpBJldNF86nqRz5Oc7BcWJXaOwvqn6+qXupRP5FOFaA+
WvK9HwS80GrQP4W1tZk/YUQwp3ziSTu45xihDJPSzwIyUZxFg48+5y4LshMlKih+
TKexGkU1BLlrLZ7i8pkeMEzaptisLETFbi4JZ4p0fi89R+8k2vp+3Q08sap2669K
WPUoCoqv20auwrndQvbXOvvnJne4eF100FgxFOJieY1OOFWAjpekRryxiVdXHEne
vIHNn121RDCAyHQUH4u20onVmeOT3gki7a2HQDzirxLE1cRyNMawyo5dOyL2nozE
mghaWIT/xUCsE3DWZj9RnuvNNKsb1C/M/8jF6q5y/2GOrn8FRMj2yfmrtPKoi+Tf
cXd18MYJvqO+1pCE53/KWjRGEs4kaSmhMA6NBj81WwiOsKijvj/G0nmgh0t0c/ez
ggTX3pNJJs62TrqICvaVGURKZtVE+NCb5W8ozWJ2KI2DV+3YGhlgAOEBvi8UdYTc
/2+61qjh2NDZA+u9YpA8Xl/0ogjHv1SF4ntLjR2vASTiIvjdnlOvPzEaGrB7+Iq3
Zq5hIMcYKWJsOWvdmjauZd8DPiwiG/+NOOTDHR8EcWrsTyIN09G+rCrTjYaCWE5N
DWi0COEdZEAgmznQL6VD8xbrDU99CV+HsLZbOOIw+80Cd61M28GfPxkoiKN3xNPx
hneLoOSnvpLBI3cVt2bRzhlUnWqjyMhireWIUMKLIL5AQQpbFapqnicvhC1xo+Yd
lg2hZeiuYFMtW5kjmPHtYKjJDwdlxaPqwiSngLi1aqNExJHY6W8nBnr0Kq2u2+SV
sXTYpmCkwPHuvUj+d6j3kc0O99m2GtZAF97Xplj9qWMaZUEp10C74Cwb/9WiR2sB
bLf3pNoO6UosKbA0AJ/mJzomWCglsDytkeCD20jHsQLDGHJcZNo07dYro13HrCRR
VBXcZ4/lWCemtXp1NFd/xTe3f1c2WjbZRWWX6FC8BUkOPS9UPuytKelvznvS3ut3
jfSa1++fCXm8u14jUQUNOfTCDp1/5F0xbcb5ggSDaS9W/sN0l29RQQLWAnsGbzdQ
LHsaAAvuGNgAxZXjsdVsOmLwEvkGR0v5zH9JX1669HFr5m8I6WUZeHxcCGEqtNxl
CYMQZXCahci54RusmJXCXrGigxMBjb4H+G7K0uSyJ0z3/VvYKenpHzCpOz0zpkBo
x66pDUairj5Aw8zqJEa1ZFdCJeBhEk1y30PvDsNHnsbtrAH8gx/CRYZA/FKuhKfM
QloTjZnbKaEeGSyW+L0zQNn5ZJNMRT0wRatZuzoRJaIWcfh0di2XYpvWlJ4WcBla
mauR3FIAGveJ9LwBnTsc/Thv00YAlENmzkco6uwd0SjBcy4EGO5tAh0X6ZhnWo5n
OOaI7TqGYDGOp+OWe3+jqfeH/2swcQeAUGZUYf9/RHZq7j+8lwb+8v5ZTcuQNH+K
F02gFK2G07OfDm3zT40jVm2CS7D/UgMlZ5toaLQSsdN1OUu0aCfA9+8/kelsrfVW
rJj5L7vpAfCDcv7Zkq+iPD3NzUkgxH6u98EzdBPNWIlkdE4ftEYhJgQwHDbHDKrT
U6K92+OLm9NaSDeLrYsf6yoGgu/n8JfFPYmCWQ4m6IGwa07SIG1MO2GVPVACpVmf
toNMpTL0A243mivWTYViRSQunR8j//nWhyt6j1OAtWsANYyN7+o0L/wJmjLbm/5L
enyu6FDQDApDsoSpdBHHgB/abofJx2zE08R813Ys5Eb7zmt3/duANlZP+lf2DBa3
WxY4B2vx30diR/rJ6xjzSbv72b9Cb0DCr4z3QwGTRw+3XYUh6gYzc+lG5rCSFeyv
sT5cRqlSZkr0KaC7jAdpTVrNyCbpOiOPJK0QTlgLfjdxsIqJmGlO+hvQ0gb2p8rh
aVycWZgqMdwmQk4lbB4sTCzDVdlB7up2fCHIMIFHZZWltBpUZK/hMbUW/jsM6h6K
glCXOvtDxC6Sy0IttiLYV81mhsjmUL9OYQgD3Kv+K6epk1ikZtYS4dsI1yP1uUFR
yyHnMvnX4QvWigdxdL0+eMrrAswyihLykdYhxAI/vZXJZV60jBf7i3FuPFn6kTq+
Pt45SgeFxiwE3mw9BVLrOtvxa23SutfU+lpt1pK03vhv4UR9UcXqwgoZaHiZI2UL
mJCTSK011vJG0p+DLBxPmAsqvQtlg2E8S+genkN2k3/SsTsfwOhq4Px0oNOYKtdh
0i9BMuwGyo4CBJ5v3zh0V+GfMU+iwUBZ5lSkWAw9Zq7+SSJTGTplJafaaCsfRfb5
HySftuVEGscmfK/7R3esyZRruXfJtDivvQLw2P5zM4g4VNSlnIPsrwwl7MUNMDLw
NcG3PL0nJj0MjaR2C/L2dV8baJM7KTnVTCs1gC5s/g0NnpH/QaPB8al8pbk3Ohte
XayfLuzOFoQC2diTWupafh5FDTaZMtgasbQ9CxIRZ/yKkawH1Mv+B+ZT6uDHVV5x
VDJ8q22sLGVt2sR0OCBsEVidZm35T8M4mZbFbWeSHdGd6r59RaXhWY7ybX83JPpx
445YRWJNewfyiCrE3j0kf0Jbyzlq08vreB/86laHXX4BSAm5bFHdXwBvT5acPGHz
CdetFJIxGoH1YMy2AmIKJoNnPIhjzo+/2uEXVrYCXJBFUh8C+y1CzDcF8yxDrngH
R1/pZ/O2ca5o88bmA/6U5EA5SQIw/PTrcg1Il6k1wj0dUTLmidAnKZw0Qr0y4U/w
LPdwe2AHxwFxxUjKzod2pSe1lZ4V+AjOLJCt+LGv1I7Kux68HIS6AfCEYUEzt+7M
3zhYz+haskdkqTKMJ5bUidGEbyust+nzBNXYeQSv3WZhPafG9lxG4rhR1rHTLZ2m
9TY43ZVRT0q54dPwa1Pd+jb9Zqzd8Yj9lbxMHrB7pGNq5a1r9fqCvGAqyQwGjc/F
rDL/GmR6CewTxUdfWHaCi3/GN+/XBLMuwUOnoKP0rHPMB8Wo1v6tC1VjK1d2SaB1
bCvXzOI96ol/OelT2Alg6COLWoUnYOiJ75PJIov0/QtLH7lFsVuisECGvaXMXh6d
4hKUuu2eO9/zXiT6yHACMu+wZiO/ZnP7NGnRI9tSYL+XsJsSEYgdrNI45UwFNRSL
CSRtRDVWiBuWBPaGM23HK/mxek600zVzNYm7nIbSjThO2Bn5zXXM/ngRpuIvMlFS
Jq8Tw9vLRUoK+4IJzG3I3+mypWBcXEt4OlUKKUQG3fyOLtAaXAuvSL4FEWYM+0s+
PcEGzdeIcd3NwoXYBv9voh/2zgcVdYZnsRPGEPfMeyZWt5CCE4/PVppKem+XS/bV
uVN4DHf7fwI3KdVfcmhuruuSijG2pd9fVJgpZNzz4nHjpYG0U82jBBqY+YTRnXLD
M+jJzIoaPIjGcG84o0FQHxhKu1PSQ7JHdoLyssEwsrlG20amCtrJ7Izopjva4EFz
clX6xO9A76D3bhxKd3/0P9cIQaWbTVozWyaxVQ52uC1bpjpT5JWE61eiLhAGs/t1
PB97Dqku8IF0liGIA3r3+2eFaHi5jk055xuPq8AOCoqPPoAKhDm8CeZj5LeHl5nM
UR6+rGmSdRDsExIJrhTeX2/O3OvXskDYnj+iMj8unZ6OEufUes+qEuCdhKFd7UJi
qBFCiAUwdyR3BBoNrBs2qIF+0kLkVh4UKo9tKEDzTtxvKO/SWlpbHjgYGLyyWlZ/
tdFs7ljwVLiI4kkdEb6ZA8cjDCZcnPCLH4l1BfSiyh0odT8CLcZg4AxGPQIxuRr1
O3Axi7COs4VJ6ZHZInO6cx61hdfUnp++1ken2UlRr42qWDC284LnxBuusCeSLW8v
mtlYP8vqubtCHIzLTpmfrd4TJGu1kyvXhHvrjytYsuIzJBJuQEHQqYbGEfprpqB9
BF5W8VEE49NlWTf6GjFN3805p0Oms4/vY+nFr/GZwG7aX9lNclVmD9XEk27jecEN
r8c45Ms2Zah43QkIUF5NXrchUKwAeuqvW2gBUnJr1PBOMlluDQxBiXed+KX3hOFr
zuSwdql/pndr0Hs5Fv47LTsgX8K7oTYS0Xkl1ATeKpNu7MhafERTKgu6qfJstRRC
S+T2t2eVf+NVm6tClD9ACQSsUhrE67g7Z4vIfVbn3eT3t5seyI9Xz/c92oaJf363
s3UDF0BQCbR5EBI/vL+NrHeaYlje9PqeMciFi9YuSSXJ9OupwrfqnZ08AHHd94q5
IfG1tX3YtY6clY4Kavq5B6kv4vv1BEkKX4n0b3Zf6ghxCuGCL+qJ3dosgt682OEj
PGDo4tqQZPlEyUvSRy1vKJ3AKjSDL9qBbf5ESjY+VGy2PFeVFxkRJohNt//1sYRV
on2QTuyNBReBqgmlx03JpNKMwHEa6dp448g+cg16VqWr5/dfZglMbPIFdS8NYmNc
rdzPyJuBAfn9vDKKt9XfPJzkR81xEu7Uh8px8PqV0n1QjCfKFg0TW+WLbFAHkIYo
0OU2/QvabbxpdDs33sR0lkYlSvr7038B/56DlhRHfyjNwWbhPEmSWxcI6Fn9UUfy
H8KpHPNxJcFZXpkEBXm2M3jstABbt9Vf5iAbMAWT1zk8gK17vaagufwfhd/g/9IV
NRiL3MlcULb1bfbwzQ84oZs/kU/HlZH1OV1MaMn6DLiKOicta/0XWouReMev/ld1
U+thXVoGe/pqD8SWgAUqvj8lefNtjcR4Eg3p1+l+Ti7c7yGUcQSk5zRVYtzniUGR
lhNj7lC9a7XimKeAiumEikbhTS0R1K2NwDMaoGuETx6LaMqbBfZcbA1DJzGcgbRH
ZBdWvzq3TcWyIGfMd5erFW0CiaOir9MyF7qdh5YfZ60LAcs+zcF5CI3PHsJDk01B
MJToiQVSmBYShz2obgdPwOLFc6FNH2id3x2gFUXQMJcRwhSG6j2jffQcABD1Vj5l
BI9ssTsL4HKjt171iWCukBfBmj+NVlheMAVoLYS4cTAcikekOiu0OL2WY1fXIe+n
VNdlS4cLnLrzbTgwixqzxIiYZ0MWcmI+TXPHf/0IsxXNB2cH0VAXunMqoEQC47a0
8vnkv/gr15pTrqAtOvY34QtJhh7rFQnOhDPzpU8IYWUJKRgcKfoFWdlNYgx9OQlA
mTSXPbpDkp5+koIYi5PQY7eQfl22MeW7vwbSDzqMYjKJAUQWPNQifyEmQxbKCXpr
H8DFgTYXgLbLjJ5fWMAcGJT8LNs7EMpVxQOIJhfUUR9VThS1IGh2w+F8nzosbDGf
TmqP02IQwgB3Yqa+wJNGpgdY9WsN0zRILLmIEe0v5q86UVJVvXDwnpS12rilL7+Z
IBN2i4uZfwhtYzrhHKfmdbirDTvQJyKmvm5K7x8PPfsREbu02jeSVbQYHN3fGX7u
XjRwUFjoVbv1h3GnDt80jZ3E8zY4GUe+NQK5CuHyFBE5UeZaz80meSAPO0kzf0ZJ
figJGODVEBis9PJifkGdCJKaE0MJYe6jTLQxX6+qufGMTE3lSnYG+QlzuZjSPixj
PkEgGjAJwk9tYCyKgQe7ElKDZxoPgpYqc9e838fsCNpWtgWulEyb6qUMuXDSdDnT
gkLb0IzTHjhP5K8GZRGt8/GB8HbRTZ/gNH1tMNm/jlxCACu1OywenfhC53VTEzTV
NCRDbvunTDfqVlkWC0qhIch/ggk56gIyoThITIUzb067U2V78yIVfDcMJIBZ3E/k
k+DUt9OwaVKRNVgVLUVInE+K4pp0rKFjZ/1ZOwt6sjUPqZymFBVtqPEmlr+uUoUh
TmgJ++c1AWoJhJWa+Jn7B1MbNydYlDd6fzHei+1hHcHoPb7nWO98mfi+gGLnpqC4
/3p+EgCVh77VlmAu3zzMk1rtHHJUQd2blyI1qkiLf4kcTU5jh2342KyPG22Kr5kq
88LtyKYWPtX1Gej5GqYMOX3vsBs+dZUGKloe2h5PWOcmmi/o9XQcWxAaMnVh3pAY
w1oWPd8XUD1et8aTINdu4OKXtY3H0NOgByekH/BJ2pK/VVwtnMHk/azaYuP2STn5
KCxC4/DkZIla4S5Z7eJeUJNleWG6NlIzvl/SSjYxVFnzUm41B+TW1sUGHddJGZpg
zSO41IEjEkWfwi7JMcXvefWNOs2nYW1b7Jz1T1kI4OV3M2CimQgR9AGgQBw6q7zK
wrONGbPkYMBIItjxGpum6H7/BcCps8w+XgO6j3ApgWIc4fHw/tTLotv3ia1vcEV9
Rt/HZ+BNTu2gycdXJ9VStnJN04SKEQXlIbsGw1b0J1Q36Oyh7nfayC5jcA4Ab5xq
7HQ4rrh2B979OVeaeh3gRIG3HH7ym4nZIV5YTH6yKe7Xrvr7VRgh5MfMXIoHVulz
gK5KLfwfDOWQlYjubyCWRxK1jcuQvP5Hynd8hWuYr6IRrZeLh0plPAeey6qfnNwR
xvcxAc22K/lGM2jD3bjVXyzWGTuTZlO12iZ0CyrPfRKiGSE+Qg9FjZZlJgYsEMOZ
tcAO1KGByFxrdRH51ajLmLcm6YA/0kH7/582Jeg+if1iZEmv/PhX+UVzIcb2Pxja
5JLiVLkU6qZ2tNuUxQzIyq/irmjXd8phJLaMErbvvU9E4dtJh+arsNJDAg/QJBr1
t0edgLr8bTpfAGDSRp5TBQGTjHTanFNMOrEK0qVhhdN1sfdAyol59ubsjcdcVAE5
kUnkc9VDcDp4N3iGlH/laaR0joO/mBgt/TyI8rWTBTiOBKXqlYZfC1c6Rkr1m7wq
ZVXB/8FnEDH0rriamqeu9WWrU388c2wfXy4yrnsJcTqxZZF5qoyfpuJVQWujBpsx
F/oxagfPmvDgDaEZG0ff0Nt2QI2S8EC9wIx6seo/drRrxpJ//AyUeilC05ZrvWUo
PsChvzTV1TdaGgHVKBpF1NpIoIzSJOQP6JMeuaWFM/M0XJh7qpEER5OUUMK4Ms42
XHRZrT6ZQ+p1FKWHq++Wz5f8phlgdZDNuAxQs0gabi8jrplUDwoMpNDfsEb1rJCg
TyJ0Ifd6jr5R+KqLtIqtVazBSKqFMzT5FSvzoNQnjRkWnxP1Sg/TXVbjQ3oe8m+q
0zhMASy+3kB3zxjNdy9mcmuVVXU2enPEMbxU36E/Qg/9zJWUzAPglRCVV08nanCV
zumwjJSpD7isATQFJXWL1dACW19c6VVAgurEjKICjEPAd3mJ1aXj7oU3ZNz22xZp
ssLov2jbnzbwet9v9sJ/4hW5JwfW2O6UD6g7ZT0Aw1lW36gdJF0NyLdJmiH9yIMg
Fo1b8NXbmFklPkmXPRzuSZZudZlVThEnA3qMyaaavU/48YdE4v12IIM38Mnrhj/4
4M6OXOLDF11SsYYWHzCQp8K8FJ6MPv4Va/lld/Iys0KM2vvgKPG6cXhxY7OwgivS
3MLYYSzoenBMY2ou5e/90MsmjolXLqyLvQH04tjsAwZmNUmnlPwcNwGUOq4g5P26
seaX4URl++DNnQ7p4j/jjMji7nrSipKCrvO6qhIVAUryvVxVejws0UP4ySA4BiEk
QmNUSt0P8o8WzpXS1OuG27pFlLLQgcJR/HRhPBM07v1ks1WUGIofsmIWJdKGEact
hosTH5I6aIZsxn6m2cvjoMS7OwBaw/fOH9z0gDy7riy7YrFPnUDfauXf/yr3+GEV
kyjChxd46ru++wdX2SfpxMYUtVk5e/c8Tfa5QUmu5jIr/1kopwboOKg5QMcsJ+ps
AQs1Jba7IMTxcBWKEUkgE2E1JO4dqkckB2NImrPkKdFf9wRJA8j7YHsC0jwYFAHC
EX4cKad1QHFuqSXY3+EQoD5Limt64XyyFsExGTKrIAdX3TukiQrSimqIduBT/2cr
XV/QRSZfQvfZGg8t6MP6Ov5vdTH0so4Y2MsW1DTqqUxpxaiFzTe4t8YYj13aefWz
jNp+75OD8BI4WtWzSO45c2wN57uhWb6dS5eO/n1u/I6ZwWZ93TPM6AnSrX/g1waP
OdCOlz06L1qtVb7tU/pAz+NvVzb88RsABjmkXnItQc48vBQx88QYBBU8wfHuFubE
mWu6yCVkxJX3ycLvGIE19mlNmCKe4ca8RO1jqpYg7wqyW6NhRndEzl0RXfguhAGS
w2Ro79jNEz2xN9txgcw8VVvaup46xMXknK6OTIfMySnmYb+hkbkY9woiqNbcbt3F
Ie3Y2JHhO4iY5vUpnXK0kIIWJbrdepWIomp3Ab5ZxrXD5zWoG46eNHwSbQQDU4fw
8JrFfLF/qIP8VjxWyNMAsrWw6Lfkiw8lCkhJA6AeKDsIOztxv+a1YKVV7/OytYi3
bpYpmNCZmF3sTBWhIvyQvWIz1ZJeSVfuRj8D0+eVZYCIKHRDOFmYTaesX6S7DWgx
v8IWYsW8vVLOnmbUisr5c/6b1bCUWcGCePrTxrI0vx7egempijyqWQuPey7mZ1v8
lopMwQWkzL0IUaRlZaJ/7lvitC0PTPjz/G8WmNqt0yipivKzxuy7XhbihFlr6FjB
rAgA2WgvwxcZTigKtkjWN/HxxJj2bdNXgwBOMSkTfUkwOycjoy8OEOWh6wimnoEA
sCY+7jodKQoomk6DZqTv/Slg+tPB3nGfa5ePrxR4OuQ3npZlsAgTBHh9G90XVQDx
8XLh+todkIjsMW42THUyJYBBVgx1LvA6e4ek9k6lvnz0PYkc99KJ2qNQy2qGaygW
FJwhcmuvV0dP1qd6azorvRVd4pMQF6AUrIvliOIJwGyWa1sb8vw/pASJHK8iOLbT
+gYUw/LcEawC7GFvbeEM+ZccQn4Gr8QI5fGUXRaZNPwvYU/ia2equyDAtm+pUEVw
oAmg/Wo5ypKbFJe/jwQajYSCuT+0++hA9HryOiKPTKO+rfThmKrgYj89fZu7oOOB
d8dXWVROGuJ8L25QWDJbMHyIyri1g/UGAbI2uQyO70PWpA6E8aDjJtj87xyPrck/
mJ4XBOr9F/bxXdAX1ucZMWXS4V94V501vLB2AjzG5Xoeb6yzRIqr2QKYOmWMrPUw
4i/0KShUqTobF9mgFEPP1R2k6qY/q+ymfPGWb+ZBWmDhloOOW7ehA3zuGPxQA4Kk
VL/tvdtGKOf9/m7Mr8FRBWIL6BfvjsEnXQE/DXC8hA/eOYLBLnDdXbsAIpe8Oh9i
uPUCPKklMgcFgDPQFa/AnFDeXAiFqLHIakiGThzlb7snr3aM8MeAZ4dSgFVUz/3L
+f8AMVR8OM7GZvgh9BGce6mC2GOXokXJBYcHteHQMtqIFNCbQTcNv6U9aIkIhAQQ
QA/OZsQ+byAqdUiUNzVHeyHaRrdyF+en1NkBMbkrtGGdj13jWV9QDV7bAl2nPX92
D0GqHm3zUAZAZOC/ofJao1GHbvyO/DsNrFrs+alBFmwrtrkINITPYbmRTBJJJdHS
JPoUlPJQnZvRSMbma4Xs/rF1tpkqjQ/aJsmnOGiNr5od8WEKI/lGRQ5kfVh08BT0
UZUg1t/JwLoNYr5jQPlM4j5cYpIo0V+BP59OdqZjPy30N+H2TJ7C7XWsdP825Y/J
xY8MDd48gNKLHaeHNqRRYcIcvpRlDlhCC6KdxEDLa55JnvRKvBqqeqrMlIByCxyS
COy+DsmS3gMb/xRhrgJosGUJnW3cc4K/b+XFc3rxnIF4cOo18Wk3imEvab7EV+4I
jiowD+Q24yIm3q6vIKjwB6VW2N63kkbbZkXW146gOCem9ry0+SCLrWZYel8rPQ57
UQPhL8g4v5zztWcEhRVzs8Z1fzdh5hADTLExIwM9HjoF4AlOGDLohLEK5cDC7yvR
oeuj8PfcrUdblHVgsPQJSLNHNn2IuNegk5tdcz4iP9uJPT8fWR8+ARN3/vb3rWux
9uM1oFSQjLXQd/FfqGhQvhhce5W0vymbR8GGCWkNabFcUPTEjJzZ4f//19AQml+W
ssrqCsi8/OIiAEvlQHREMuiGZNq/dsaPj3KWdesYa7oRXmDWvRZCiDa07rOLMRgO
enPHr/ry8QNl9pigHDwjSVTl/C0VjDs/QHPnKtgBExVCmq1Qf7BfXbPo42zl+AK2
VnNBqghU0dHN2eLPla8Xzj/ZkIDMC2DQRh8JMhmUcLxHex6UkX56wirfBWGbODLq
vONFtk1BrqvVTzjFtaw+vzkQSst6vpCXzJAA7xlvYLl88elEp6iNlKfuirsbN65e
KJNgNrlpkRTbhEMkeTTSBpoCHogf0PXvecY9H2AmwWDAcw4jsPh6lq4qTw6TTbTl
XpPXmxzmNPvHxBcvUx/4000VT2CBjO1+r0gPeGKMsACaXvb6V0nb2Z/oZLF2vSRA
NLSROtsrdkTCbBJOBgWFL+xW5lEDYSnibQP8OZi/F3y7rE9DQMfXOkU0/X67CrMh
nZb6EP10Fm9R7OipW0FNCGKkD8jGf6iQCE4HlwAWCAqo6Ln+IeZCjFeQG0lanp0O
g6waGiLujI9lvGFD9+Ru+rC0o4yuRcupYiuWud9O2aMaESqOqRADXINkLTCV15BL
ltyIWamBpzfutxsuQt2BFONwaTF62eguawqKcm0YzPeZS2enE0soc1f/KM+kvgvD
3T9B6pWHvKPZqZexUitSKjhpXT6KDqCOsEUmhoA++QXlCy/nN1SqzmS9D7Mdcrmi
xraUD82yG61X6vx04ooDl+mlir+pmN9Mo/TOcCb8YejPM47j2n/j71N63E6QhnOj
WizMNJgtJQkicL8SohBv0bEpsLmLLKm0JfJLsFSvcItDxNSpmzJaMsCgrdcLZm2H
77xxJnyKPnSTH44HGAZg/H9IzY1e43ZehtCz6rGCmfRjrWbF3Mh/LWQLrX4VMm+i
DpudJ3pE2u4wXMMKMB/Q6PxlAk4Wi4Qm3vNzpFy4sNpkn9lAfyZuDhlisZKJvE3H
pSt5iyKKsKZpSDfG2V+dDWxrQH5WyD9QubzmXstZsNdurhVgJKlHzdjpcQBlHMGO
Uy0IjughjTpZLyL2fli2wOwcpAs95nqKN6GSggwwokVnT+Rn6HTu19n9NuBODL8o
jc1tpNYwdpeJ5ZiKgWL5V7PAQPCCJPq0GkR3CRia6/ZHNJoI/7Ok2R2gmyS5c9dU
wxS6eRLJ+jTjCpI5SSw+hAhDE0OlXSez9qulhvgXC/H0p47CQJAjKjiDtKw2UhPE
TD+YzhPzShzl/kg7HJgWJKLoFm3YmAoINLvYfuyFBEuP80wtcS5yuYFZwoZJit+J
8YxIrw07cK7GqOu/g6wOkeieYJicf3s2HAB8+3ZRtuZXrr5kquQDMSEPPxhkPCQE
+jx9l63L700NQ1pWTbMfpfB+j8xxUvaKbiYGoAC/3mzQiGwqkZDJgH7QI3apKKJS
iGfGkxDBe7ugqB5PaBKiSpN1ljBsyM9Fc1+LcVXGjhul4nmzKC1fdv66+nwamHv1
SPbc59SpIdg528VblRG8oFM+95DSn6N8h2qVCKEaaWenBUBdOFACCS2xhorZRE/V
nZxHtVmMv5fQW59NLF99C6v6xN35mh679V+37pnysj/ndb1uK4AO5Mv1X8sSlYnh
+yqtQfA3Xols9MRyKFxynjm9ChiRE90UvoXUQlfNhgT89CGz4lQcy9/sNIGnKAVA
llZzUc9QExRFkuncXyrEFA8DLTii+bBIla1O5KngKsZ0b/KZBSc/0k8JN+HYDaml
Yk/U+oMJacVjKtAIMm0nubTZO+QXKNowVTP4tuTXIGebfuPKel9ZTL5Cl9yCtdVf
Cg0hADy3Kcs/rUbzPLn4ChpGSfcqhAoM+IPHy1pZZVeIMzrIa6d+rb7lEOR7XFew
4vjObMg05H4t9N5KY33pyxD7Fsk8EbME2qwoMuqD9uZJtBlMhT3YRk2NqYaVasCb
9lV8W4HwLyutcOiUSlFbCOIfqMxXj7/dobku2RHAFVaIPtONcPNJ5Ty6Qa92EhA5
8N2VZrYiKQzKMPg5s2P1r4vAETdXhkwAmazUupZWuovEaAjt08KG+gNHTpqcMhUa
xrh/Lf8BF0mEAHh5VpUeOqd5TyekBiiAdFgSOZiYGHlrU6sIBlxZ9eKFTpDdwmLe
QzWZXd3MnvkqqTqPGXEeNsnNkdRz01uFGs9yrI39q3X7M7hoP57iHKKTor0JXlIk
BQsCcdzf7IfrFBp/ONC0x6euJ0PAF6LmSIhusQjZvs1XXoO+F2JDZsfrzXZdY7B/
ntD3dfQw5KxTcfin+tHR4oYdtNhpNJClI7MmopgTAcBDXqRPXECbOVkZ6tbEeTyT
C2eIAuMpHIPwffy0m12ZdhCWjCzqWO2bWN/YPN3rtgx7qjb6qLaosU9WjRlxrmoC
M/+U1P00vZlQ9IqMfuvDJwOfr1aD3BXdEdULaYXHLFRiuHvMJVvsHw4ftN9j5Kiy
LT731WkvddmANpu8tRasMN4kkKtfE6kpMhmSedKKeeV3MCrHxxinNG/kz7ePF9BP
+nwKAsujsaWxxIRawS6UnMDrT8RU2MhsaikLfnXOxncXMjcOA2KcI2ZJcf5C3FtK
3vfk/IvK/+vFJcyjq0fYaw9SzzRxBpv4wXOHng1RT0uVPoQHH1HALnYCi1cSan8B
4dsxq0K0KGl07TwKeTTZkMXVf7D6bWkDTicnFXgWiK+xqJH57g+UpyYM2rX8yDPP
3gXFXMZW5butsCZsdHvpfaMlyliG3AzHbDfm2VxCDtoyMoj6job6pZoQZoSl70WF
w8lZcFJHgWrA8FFfO0FriT8gMCGeN16Tv48trrsGsCxsAsmXi2UnzSs6JAR4TYLI
UeSkSZQ3it0lR+YwlIbDKmB8HPPzH3O6Fsp4WwiZZOXp7k06I5hvTZabhiyGKEkP
OqwKBC/zkyn5iZOQ0qMNy5U8sHnNzo1Yx1B0a2VXqi2fwS4n1CjwKLUInwzSe2fp
1FONpKlsf8hJP9npCVRcTeQ4lxJTgCBAEhhYasfY/DC4WbWYL8Nlh4+0WAY7Qh24
h4PN7J0QnVwBK3ePrsYTpFZU1UlqBe5or4dMNiGrVZUGRrl/XAT5KT44iRe8PKY2
T6twBVoiO9ILkr5l+zFAmA5JRhj7T3+ZK7BtKW7mP/9RRUnf5bwIR223rUESHl8I
LaArP3/5B15/kI/aPlfxXHqnj/AP89zW3nLU34GI127yorvqVLnye38jB20N8F+e
/AVmrQytepc5xIfxa+rNR5VwL+Km5Y853G7XYdNpYGH3XpqUoaEnLJkl61w6buEs
vNJiLCyespv42z2cuWut7yyz2gco3GPXYfSTDZCAAurvh/cgzSSFpqGwh+BMrCka
ubLxf/dzk116e1JenOpPKxgnBShn4WxW5QdyO3XaIT59Ztnmj/Ut7DQDMsURLgJi
lZ/WEk5O7GE6AdVGaxwTwXFvhqnz0KsDN7yiDAOL0bFl95k4ue2nitp1UdkTA+zi
511Q+s4l5jqmnaUal9o931DcsB5veY/ukyuTtWcmKpmoXYaoL8i7zSwXKmqcU74Z
IQwbMcmJR1q/RMgseJMLWWegUfaFeLXQoiIxDVX8TwfcGUSA2i4oHEHrGJUV5HER
lGbWaBAbINI5eCCDI+Vo+ZWv8Umkx+UUQHvpjCMAD6fxIIiyA9m05/iBRHN8Wc/8
1/1F/tEqeNe07xNmC9dw7CXiNmFosjnhSspEeN6tO0YqWsFAFKjhgvgq+luJ5Mnc
q3jD9moaUkFSrucJrjom4M7RAVBp65+Hh84USNJ+Hm0OehjrPjam2XOZe4LInmir
ZdIQxUbnfpNRYkcPNuRtMtGiVPFGtwMFcBX2n9JOILDUXSnJNaE2EJ4xc0NqtLxi
/JUuAivdUeCvWF+WzYd9+R+jgtUOe1uk/22HSnP+Nc2b6HAB2HHRO2qzOsLNG6/D
Ir523PpmFhv+4xxOl2+LB11lcHR2ct0mT+aoViEfNy8KyiP6j4xjcHrytQIGaXFr
ieOKMWjoP6Yuc5f/9ngmNJ+2zfUV013cNh8W9vxWOJv4a57g5a6wydnhgT40st0e
JsNt4ZR6hBotKvYoqkCEaEVhijEEq+ZU5gt59fcp6fMyz3gawL1sscebZlv8otEX
0QDbu2B9ujr5iMcJbqnWWYDI5NYbmF+tG7XmvrTkAyfG+oTa/r++zDW7qykmHXlJ
tTuastTRBVB7PurKEleNRNLtw5ntx6Stq+HS5BMDo44Rhvnn0ar9v/aQKc5lEDkO
rBRY2BAaESWtmLxNnpgXjoGMPmHt1EB1R47ibQPRcK17gSrc5ikQme52yRkIgSds
T7h6yutT85LUklp4HdvznOlmRNSKfmvDhPlxfD9ySm/AXKE3aPSWte4lWWOqmG7B
a+QKf7TBnEoG85CAQHU5F4XNFCAxD+W9igmiiYgYTFhgi/0nRtv7MEYNnUnHJSsX
rpHdVJpD1kWaghGqNv1Xt1GrSroL4rQZzi+Wer9jsUXz63Hl/bR5+G+wdl9xII6d
9mPiNTljUuM2s+yqfCkIRANol1Vn0z9JqpkrJ39QYBJMJQp20Ss/ABSrrZIVLquS
zW9SxxmnWq3N+5eLMejPZFw++VAYO2/MwgbV/wBFBza/xGZkqQvTCnm7ktlnihzJ
9/1HVwcOOfn/HyjeJrm9sMWwmMZTwutcf3KofU/ea1+0JCfN6E8qJy95HbIg/JAL
eI5Teg+uJHnohWkqcMdSOGEDAhRKll0YzfqJF4+4GKqZP1xvU5yIWhKeqX4jEQwz
cEKMk2jsmgJGWwYFRm3ALetIfhoDhzUEnYLZPUi1xDvu966zOePtVaBkdQ05w13A
zR96ljNPDIspDMdl5et18Jz2htrPcHchEkMlBHFPw856UWw5EloU8+RGrRepczxb
VoOL9zcTlm46JgEB0X5pU6pJSIMqr0Ar90gc7v041PhLA4R4wE8J0cDS6QjCLEQs
RQg3jNOk0V2v8SWBpYt4sw9vf4NC/36oBRREsB/IroZC99hyOkr305Z1MGd7gEoF
xJFHnLBLkDVh+8WJtgZw2NXkujD62ReB43T+dPNUPzkQWbrd2KGO5W9vTltJ2ySx
kThvdN+jmSY17w4V1oncA3sE5MghQ93+1/Jet522k4k4yFIauQAUquRkYwyroT7Z
78DcFdNxJC2viVyk2iTflGfsBqKNzTObE2W7ViO/tuuPKYM2+ZqSOLlwduBZs8b9
KozoWdDKeHSpwcFnA1VAEJbcL0AgpeYJnVgznsjNcMM43MBGtWM0KdAhffMqiUEf
iHmlmXoybimnS+QMYwuDXRN5G+5DpYehuhdwHShfo5nIOR0TxU/ERJM13b9Sy1K/
Rf8lcc1AP/p0cgeo4Zf15EQim40UT2sBDoGrZto68xQLflpFAGdeeKXMggV/mR+N
YjI66+3c1KsJMA1QrRmzcSPlCcZqRQc8j5mzePrsBkpcHDvOhHItYwnyOpE524lv
7au3EG6ytxxcfbj/iGAcaGEdO4sFrujl1Ol2cfdBpYCR9G1bCARwvQ29/4byNnjI
zPPQPDGY8OW5qV1u2FsxVpyx6vsQBfo5LUgATZPqReBM7W11cxmYH7mZ74RutaKp
1VFz0NMzhUzV4XwBpRYqttz80/sYDMcE7IRH6l0kzgdmY+W6xAVufyDHiTVhAemg
Q9xmEgBd+0qVQVUw0oVgJ4aTBebnl0AO8Tc4Gq4ehABgcDHgMIqeyfmDycePjlow
iKzmBRcdFs3GmMwNw5SfVKX83vMoUqB4xYFmJzfKtNDQv0mcbt2U/JRF3n4Bj3Fi
aW5R7qeU2nunZ0ZNoCRCppiEPEA0QsPwYQz0unQ8kXld53MZaHa5HHVhkg8IbZh/
W0/l3OH7wS7QWGxFVgslyfVix79m1XfUvpWNQkzG0+1oDcoagFV0BvI5KR6RHMa1
bJa1x1xWn8XIjIW+QEtYx6vZkrMnmc23kr+/fAFYIm4sYj1WDmCeqk6iuDNsWBSB
qYAHj5j0y0sgP0uQ8XfIq1ON37AzTSABCCjScZEEe/+KSdPYIPE1ISic4hOmBAA5
FWJJau1Bqiu6LvyqlQ4Z82wbv5J2flLTI2H3VeL/CBr5wVNhyHA/t1pWm1VuRClz
biqnw00qRV9O5drv0b3xQ2eiK+faxNdR1eeRsVpD7oz+O1TxWRBuDCord8CIqeaW
ifCZvx0c4RPJtK+4TstMzBaeQ10KDAQtKg0nHa3csLyZGgM72mM17G5XdWGAlHXa
0rQ9AveXdim6Qh1R7aj4aHb4C7ugnRHVNFc4oG2Jd3o8+s6efVo6y6e0nNj5lm3b
v5qNHF/iaeufuNiS4ZNc94timOZjy5SRENTq/Di9Mn8+WDaQoWzsjVvPQBmJrVvW
nqwp5Q7DrRmt043hvw05q+X0uRLcfrQIloRpt9te730wMRoo2wCf8maHJPPBxq3w
mh8gwp19+iWc7spob7I80Glmb6YYnMRrYXSxVGGSDpATqPEnIeyQm1++h/Szo6rf
TiI/1aQVSC9DtUL7nNle6cK8ZODHw82mbObIJZr6r0+n22MZiklmeaDCOkD3nVe7
iFZtsw9rkCcW1O7yTSHfqDABkOnuOIMjssYY498IAs0zG37UtR6+k68q2qZcM2Aw
khDLY9BlFbKizF2JvhIJy9t96b1Y68dqalS+KuoOixJyz1FhPWN3Kr8GURLj9EMq
x+U+7ytJkHusH5bifVcC3cJyEYQItO8IddbULFQM0CtR5eSN7Xj6VzeiyJBrSYvV
7rLs0LWnkbOSzz0O2mc6RD9hNqh2SuSx0R3HvkHd4n6lllR6Kbbcw8KFi7dsrGsa
bhbe4XXqHLDQ7aI7leuCrp3a72ZgR6sR9na/D247nIfK6FcFGHceovv1nSPt5oC5
K9PqonLTHhLRYkpkjTJmnJDYBoXa3R4sTW+ea5Zk+z5+COmRxUFNUpXCizZrjpDF
3OEH8uECp0K4qYKspsnuPRztUUyXyvS/ssmLuoHMaRyPeSTbUUj2Sqa+46mg7skt
JU34jf4Rwn2uRb2iKdEevEjpQqh/F1fOyyxf3rV7uQ/RNelQbZu/xyKooepZ8+Mw
ZjaY1t9lF2y///CUSox0199GDafB46je3bU4lvTGVd6/AaU1ODF39GJ1mo53A8hd
wkUTZXjlqyBFTqWcvfl8R8wpYfGijb+5IUVvd6Q/dWrQ6HSIy8rBEr+7Ur6MyJ7/
wyMSvgvRAwT6YuR+27idKFtLfV7xkcwVd/kXq2Z965KgZBNXK49cZxfUih7L94y9
WinSfOldeutDI0l6X8gO5Pp2AGATd2vKQnLCkTQ5/hLbIJ9OfqYvJzcju1BJXOkm
5GX855GL3vKcZYeBEZZgeXUUuFx02AAh6A+tDrq4P0kTBTcRPyy7FYiOLjl5Vwap
wVIwTfXUhdlWq38EeNx1KpECqcjIz1+iaCyzfHA7itS1UR/aDj2mVuyk5Eck2QbL
XgiMJqLleGPD3fFGzDCKLCb4PlY6qmQMF7HOqIQZs+0yvzHbKiMBGTe3ap8o5aQ/
viDaW0qyVmFcsHpUg2eBAo4LLTQtsS4NH2rnpUnL3Kp8yunsFlWDEq/SLm7GbdHe
JvKjPhCKTuxYh1ZlYACsRS3b3pSqpdd89e+TkH61vpSElB65ljb+q9zB350xVkpY
aN+3MzG7OvR/flXgt7QeP2PB/TA45XVNCFR7KfcP7eZMly2gdEN2L28Y2Z2e369c
J+pK8fB2ioslznypxQ99rOO7uW0HdwwpJC2/AZ77RALQQ19Js284jx6W5+7/3B02
q92lK/tP6gVQoDjE/oqWG1Czf8FksSZreKsVyCZ1L/8T5XrCCytk+ftQ2UPVTg+3
KRjlv4bfAtYiCnCggPOPJmDe218ZyLEKKllE2n985dlhdXLlmPDCSKb062+z9Td3
TIhBBHlvM1YlXJ+QxTUo5HBzm/mJ1IcswtyOUOuPplq28u1WATkTnherT/U4V5QY
pxcjwo0BQdXEqa+5kfAGM38jnvKYa0NJU3I+brnfaKQ33ACpE+Gm3dQ0kC6FlEjP
xYz/cuXmolIVRl0K9NZ3RypJe6lMR+3kDYCSUduw6jeoUMRgYEA8whdnRe+dTwUZ
OjM3UwL1bSCjhvnRGPuanPy5PV9YqVIt2b7XNGpnjJemSmoaZ/t6EcVMC/7P0Hrz
BCnOYgdHKTlY1oPdUIq1OaRDXvpKSOY2eEsgFvr/tB0oXu2GNfYruqcguTE0DGT3
NdEJ0OGLWO2og4WAu5I8HxjeKYd9pVzlpWcy7cHFsqgMPctBgHzVGk0hvC0LhEyZ
tRiTVRti9UIC2iD2nK1fcmxfQ+nWGIx598aKmy+MbhHhTu94Kg5TyHY030/VzgeZ
09zTj4rA+YvSF+XhIvVQX85BAPjOGKolaU+jeCUCKv+Ti02AlZdCsklOLgSc4ILc
oScRazRCwwVg4rPijdl+GB2+V7VjNgW2y3b+HEWIz6uAKUI/fiAHOcCDWpqIkZxG
CO8Wsu9u4ZClbX7u2Adoi1/hr8DDiVBccYcmSIxJdep8Lr/tWNLO0HBg8pogLbJX
f3HWPXXFiu071rwmySu3mXi4OmOsY9nVWW2//0e0A912JCfL/Zy4CbAn3lyNBGCl
XNmZkk5JlP5plT/lKoZsp/h7RYrX9qw+k3e8mlzJsr3n4GcGtp26t2EwOL3lJWxf
XpvRSXS9LwtG2SucFyCd3UJX9bK21tL6ImjPjmRrCjeUd8/y/WFqRJuzHSxXUzNt
42dNT9FI4Fc723xWYK/ZipT0wz4GmURx532UL0AO2YzsDa1pLNeMxdk3R2zcQrQH
A+VjFwXt8dRdxkavg0qJ8tqVFO89Icny6NcxdzoAmLXYZcLH8+/xPsRFnrkcIrET
61cVj/BZ9zNVJvWtP+KVG5lDnEdYYMovqQcDZqUzJzqX5wMStLevLKHJNP5e4JuL
0h1ieQkpcqcjdBQrKLmiwWIVF8kls99crbMeazd/Dmzhu24nM9u50piMRsR1jw3e
uoIuEL1Mum2JyMHxYM19TdzD9yCa2vI2yIJ0+SUHoJTKgzgvbfmHY7VGa1rUkZz2
LXrsLpO8+TWUQ/cPYLDIaN0ljbRUbCBnfRX8jTYfmyNjKTbyNIvmV+pVznqZD3S+
QAjB3iw//LDQsuTZl97t31cME9upEJg3d6eoYCsl6hdTIJk3jNoX+J705wKN7hJp
ajTua1mpx+DYw8yozVtLYULJ+ZZy9I8i05fogPe2AUj+9ACCw5ozKnfvaYk4rR84
QEQUm2jnbWxGujCALazYx0GK3l4wrRixHG56oSnYTZTo+cEsmRcEeg5lGGMNMztW
zoHu900b1O0YngR3C+SRniLPt/AsKTOJcryE1cIHhHdRHPnJU8YCJobKl3X/xd1Y
i92o/wOMyoQunt1m5+C2DPVjEJjCfkBwS6HEZXIPoLWqfvj6Fc/Lbe6/Zg9oqpXY
BAuFl3e59axkDhUpRWx+DNB1fmi0ZNYMcSNFYi7yFwwkAF0ZWmQ+3u/yKB3abqh3
8wt/Tdb3yEOay+7BRkkoA0r2S9uKebQ1RXWhbpUK9wz1FYkTXv1jQcmqUY1MPXtI
vxcBcYCWjxBnFuJ2c5dbUngSHQOvzIlb3NFUVWCCmkLeJXLQjqtABjtHOxFWXNRK
2QIg45Vfy1CaY2eGlogdlUwhtO7Xx2mbcSEt/kCDVs0ukHHGYaKkn9hSOejQzFtB
EQX6kJhhNdNnD3rReMlib8+AC05D1P3usLMphX8eBalVhyGfTs3jyqTW47f7YA6n
9oJY/J7FOh/f9H6mziHU8b2U0Cbw6FYD5/ktGBlDsWxxFfUWsqQVOzBguGqQ/ILZ
shrz2EHDPNOtNhEQVyEXHCVWGin2gfw676VpAlZJZIAMPU+wmH7a42QxwV8T4J2c
n6eXMlf7FlkuHWVfw/LUUJYGuuLjE+G062lpWN4pi+oVlEZzvyk0H1+GTSgpz/vR
Wa6lVv4GO9ur8lmNmC7KdhLr9tQUmHvMAb3quqcd3NIVPBahTs7zmH4G2YajzWAy
KWZARIWT11XUFEzkxMYZxM7TnvNLHj6vPoPDn5ExaMh/MrPo/JvurffcpJAeVTkL
DGWx7f/SQZyOLkqLWDRuyHvp/3VfoinM63IQxCiyNvc76KnEM4wf+ucUr1Errqxr
7kP8JMafcCFb6aE4s5bD87me233Mxv0SlW6p17o0EDCDg4RyR+pewxzLQbGrCfzW
WDjuMN98eIV6Sxr7voPnob5mQ92T4XxDwkm1nWzJ43QbF/w7ukZ7AqNJuJWjYWYH
SO+E+rC8EEBpQzzdKCTnqDLJi6VboZzH6n5Cwh9hnGTJYRtPP82l/+fSl0P1GiBi
foucjGLQWPoCCxW7gvUm16Vaw9kmH4AqCPoGHGqJdinWi4HijR3DXI0sgjH6Naa7
W4NrPguAHiXKY9McQb7REH7OJXaDazbjl0pCyhDldIVnc1tpUcrGcHN2nZRGvvpe
KA9NBHD1sHKzzEwGUeJa8BOBGFWXx64DfjcC5LN5gBkrNTsj4TMyQhYBRh+ZKoVI
u/nSrfYugcxdSk6Az4VYs3J6ryz9/snX8vfA5YvCCQq5Qmw9qBLhli3zrliEEnO0
swwUsutU/+9Tq7IFifbjnAVVMknU7K0V5EeAGFhKZUU4azfHJnboYTGVnahdqgj6
0+ZfuRIcIUiNcN4CShMW2hFlFKRwTmnMNfCF5CNkMN+Q6JR75rafzYg+Tdw1OR7S
AXcBTRQ2xYjb5E9BDwtTXTgrXJDpUdZN5MVYLMQEQvbo+zYtunuPC+RK48p6X71w
`protect END_PROTECTED
