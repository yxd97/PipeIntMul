`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSeCmpKatnhQk7h2ymWU44JfHDVRqyivzKrjVdgZHQHTbQ6ucwFng9ZrUWl9MoNN
IE4tvRn6KiBcHVUGGVnFpMYGs21tDRcx4mi7MnxlSFCaB0DtqbIgg2p4q247FMdB
iI7zvHxoWwJ1FvUomTYyQN5uJrV6ShGf90kpTkXOeIoIh7imC2mzRwnzq3Isc2qy
tLsPDdp3sTbWB1qxTLaV1eou5R9KiwNIa6sFJWYdWWMgz/gFJ9FFy0wyMVS4XqN0
oyioJwPoLe1onZ76JMNTIlm1rxAXzVkvKraZAI3cV0mFEUcI7QS0firc7BNUn65f
/chLSaAc8YF/8DMLRxjxOWBSPjUB5XaCjLu93vZwjVgkats573qK8R+igLZ78MJq
E7sgWQ8OP9/gQMrgU4WkoADcO1cW5M3Pc1wJbTvn3+uYrvBfi33c6xpgC3w0KwhL
IuzNhBZvzng0c7VXWLbQYUohU70vRCAsNDdzingCuFw=
`protect END_PROTECTED
