`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ExqTRIdqoGPAxj27zIdQQei7y05J+kH/cn25P17x9zflznm0EGKeTpNVmU4FES+u
BrvcibxzN7/VKQctSfdGwXOTv57YZtK6DuHid4+5Tashe0TEQXOoNcby2LPlH9sR
H7Jmg7b6b8teKYTZx6MIrNHuyznOoR2ELpQekAxqVA4S96JqS1GgN208nCdoEgFp
DhPNufnpDvPth4Bfvq73Qtr58JrObRbJjf6bsnrDvVS8RaPcpCfhIC2/dGc0OGaO
tambqcj50Dll3dH6yx+55lOgrRg9LJdWyIqgYmDW6e3Y3918fFQh9ythDy/Iw9uC
l5iz5SKH82NV8Agq49TsEKBaTgXOTm/Lx5vq5bVQbJjjBLCbeF5cZ3WcguLGoVgq
xyTqbVRdgmpaQXSxpOEvv6vLlLPuIn5c+iY2q9V2ct2m2CCx2HTWeEbKaoMYzSYO
oGVytO9FPDk6yIS8r1KFPrC4wUpaagoqxkF4qbSlSiEdlIiYCTx1d6zD2ZNW6WA0
cBHxMaqKeWxPG+NErccl+SjPN3g7NI1a7/jUOuHMLxfqu5EBmRiwlzuV1iXMaLWO
KdXQ9TkcGfpQHcgbLHj7cXOmJSPSsPGphfULxEoHctOYjhs5W7XN1EdDaKL7tHPB
yzDJbBUjY1hCPUwO/28N7EhVhDGOxxwKC5YU1mRr/oe+sULDzlgSw3mrkxt1k0/P
LH+QHpopGkQiy32BgSAw1GCB8NtimDJb6LAaHBtJ+4OtvkArLDmvqb9Nk3gxbKvY
n2XmZu774mEAPADpFEmU9LkCqbY4GxkOgBYeW0tvJZ7glJ3NKXVfcS1kY33OqfhA
Gz625zAdyxl+mraPgVJrlmoLKvfQxAhmbY+hg3tO/V4ZWajADtec4pXR+NCUn4JD
e1XNPCNVBxa8fwFVrSPkWFsD8Yzr3JgSUK3TRg0rT6d93FegMZWxnH1omnnYZfkp
vTYUPNJ4n2ZrFH3sjvBkeUrM9Mt4IU1eptPptgDCUtfWEkUH0KMlQOWk3j2GLmvl
ObVeUl7G3Vn1Xs/piR8Z1lxnUzo0nldJVaoNoMMMq6LnaEyvfEJMtOmF+pcZrB40
QBb40peHit0emUDoSOSfdV0ntmDy8y9umxw9SgLgGUsjgQmseaqpy7csSFc2S+QU
sf4+WXalBggG1MNWwxllNgRPPrf4cftyrexi4GV3KtWZn+1dLR87hH42KGYoAucr
rreKCD2mAGEZXSeIahaYY3W82128ZQ0pM9YXBiJRiYIuwv8XUiXaWIOlFlSzh01y
/ehrIgBU2XiitPS8Tnn5XZZsdX0WITQACYXycdPxlF3Y1nLyh7HWusRRhMj959gz
AsSTBHi2DF/fvNPIYM5nKW98lfKkhNbeg7fa5Ovm+sFc1e0G93Wq28K4sMHky2ay
A9MvvVncSHOjqQwBIWQRpmrckMAaxxYYIqA5nqoiJMAkdfyAqz+pe3wYI+aGC1bi
dhaYOXPoVmY1KP76a6DVGip+cb5cz+odKyabgJVwaE1bmq301VbLG58FOWjA7OOL
2Ehd5ufJc+NeqvIaH7NXUjBRmItSfJjANkQFTuui/QyGZjMD7Bj1AX6GlVW4nLrb
d1PDMaLWSeBnnld6+HiTC63TZtjCqZAwtME2SIRIf4ycnNS0abYXwc/JE+Z8kQh/
F2jmUtJoVh+BMPTJKn16e8ejpf5NfBJJZhCFNpzxgbM9xrHOtQO6w1J4l4XyA6C1
auYCAQNKwFO/YkR4435oQbU2nr+zv1XUg6bkj9o20lE=
`protect END_PROTECTED
