`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wwh0zmQ1OUMiLC1QRTaCxzJnuYchC2aoKsavHrH3V2m6vIcZtxDnnTWqhQZzO5X
kmV9LAou7ATiwOlvMpJZQwbhe1iSzZTV4O+Js9HvwdMOSnrIFawM1zwWtJTHnmwY
7MwAWIgaVhPvBu+1aLXBGoxFQjlGVxnjp8skdnhsj0VT85WytQDvmen7SalvOB4C
5GpLG2/mDjNwwwwva6v6yiA35TQR29ky5xkcHqI/lEXInCkX799PoAbGMGCSKzrH
yE791eH0OfHxb4Pu/6GBeXIr0dJ4HF3GuRUPnbmCWBgL9Kq1LnYSqiZ9lJjxZc6l
/qPkvBJ6QF7DQ4EWsPw5VgVpm925EZHdinEdMWOKS/J1wBPFjDLRdsxFUFkCYTYC
0Lvw5Gw3bjAhc+tFBX5wyKuDkqQcJGx1zsGiKObQiIWpgdfyc5JhPDSJrtG9tSqm
`protect END_PROTECTED
