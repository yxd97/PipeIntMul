`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4wO3t3fBMsBw4iwslPiHTx3jy2hJTyaBle8OfjvZ7AF4/iFHMoCYF2Mav+YIE+dN
BCCIgaWT253q5nnRCzcrHErieeEXDcmc7oQQqHnBzJeT8WFKdltYlRN+y8KPg2WW
dR5QlqyNS1LSnaHHZh/Sy251b+EHriSKGqoiwuIztvyhQ5iCtCWk75rkq23jdE4m
CeUPJxa0DAKKwoQDZOHzdLhP3GAMuFpT7k7VEob8Xb3WW1O22OIbRCyFa3O5h8wJ
WA+JWC/5ikrpE8ErUk9fO11t3trAovl82cSzrilEskk0FzknfVzjIsAq+g8FB8l8
w05MIYY+EsPVvnuMyG3C5tdD+Vcsvci+4ifdkUlIsW5PScvVnQ5MdeVJcXodb2v2
ILk14yracjOe8oBpDWfwWsWFHbzZIoj5V7Ye8XMb+nC+PyWMqeMDrLumQGWMPpXo
SXBt0byZNb0/KA5EYCFPb0rLBmp/x4voAM7ve2d4BR8=
`protect END_PROTECTED
