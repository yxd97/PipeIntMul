`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dx8XMy3Vd6F82GZQ46WEw6/lqQf2JPeV2zpZGt3i5i2JLhgeJSmUNEdsp3giCshq
yZFKJDmZQi8vvSDWq63Oh6HuxcgoE2UhLWQm4nal5k4kIxtBA747xRbJGcQEcRSN
xBS24C5AN3dIi4uRi45uOjs27IcKrMGtOVZxLEQDI22cAinuV2U36SkTEgO+o+6d
L+rFM68977gpJ5eiNDlvGRUj+uwSZr7xTyHnYRYtcL/x/CmtKMPls+M3cGqsEzQl
SubUo12JeAgqDFAsuj0ut8wyJATlT/15E7QpBcOz814SACnRJRZs1tcuvL+eB7GG
mvAz3rcbjUgx4XTH5QdWEC/EiJ7c4zx4jGU72lTMQm80SRGZmaFsqbKxsV23Y00C
2QEc2MQDfcn282NOgy2YY/5fIZDpliTAypeu6haAPZToMrdhWmKo2biTCsG7JVXd
FtTb/rP0ISL5IZH9RxW0BA==
`protect END_PROTECTED
