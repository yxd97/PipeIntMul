`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15dvAUPB45x2A7g+1uJLNXjWndTrod6sviq7d7Qzt0a/FiZ3cgAgSl853jVtOWyO
6uswx36vqxErfzRhNjt6Gj48B7i6V3z9q2/bSAvJ7JOquwYWA1jONcq4De/0146G
joN82BwZ/wC/NxiXFz3+kQZ47jvxAuvElJrALX5NNLnm+NCXhAgl21OlwP9JS9wY
wLm1f/s1dwgrE1MsJ06JLlfwY/YYfGO+YDiBP35LTl8DRLQs8gVuR3O0p6NM3IPO
ZQYriTroMtS9nd5N/T2gfg==
`protect END_PROTECTED
