`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YjnleHhCPTFxz4CALdM/qILEe+G6XcGFZCafrgOIknaDklMRaAiEvRpuJPc6iPUh
oitI9y+RcXMzkJ/oX8u7sz7VhRhIYo7NeBDDohQbwBgEF4UfXwi+e3iNmbF0y5ch
Jq9BTz/k3nw2/A1Edof9tCFQCiPs+Lo4XwXnB1YRM8OgcTYFNlG/tIZFXpk4wWNF
SRFLeCLw/g57oWP0EobSOP1sWT+zU7RA8i0wTrxuGrXiZMFI4nt2WMFQTRFm3HOP
s6x02AaudXXCRYOU47tVzivAMV6hdaH7rPCNkR9+W8M1NONEf7aM9NBhXksleAW1
5GnpzpMXLmYERh7wba5srCZAMdJu8OBYVBL+Xv7cpiA1AX+E4qRKyWgB54/VoEzW
YOy9GD5UIt4Sz92Puj7Ap8/VAybxfLRDJh4sTaM0EI2utUspmict0SLjJZY2OrdJ
+3uPZn/i9f8Rw2NAyVig3kE8vhCCbO7fZUgO9yAbM9hJCri/DZKlAjaNFene6KCg
`protect END_PROTECTED
