`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKCVC8G7QoWZhS8oYeozxOUfRiMg/KU3snWOTVwTGKrvtyX6x4olX92cH2ok6g/7
j0O+8L1ZOYRpn0X0Ht0NaHupyhZNHvE+zKchxKLYoavb/MTPyxhuhnwLaZLxM7+m
ivp/tJqIEJUFfypnMopqA0mqqt4iVSwhK6SXR7STwB2u74gJCsv1sExdtS9bRIWQ
IZPnnClfa5LE3WQYBsMdu2zoKEFhoeCYCp+zTFo3g15HqHGPDiNb7CR56Wy3ij0a
yHZduFiyIvq/UXM+o3/ZXvHCeitjfXQMAl0aiF2kcWkA6q68xzc4C98mQIhPp8aj
LdV1FjR6x5zRaU7s3a2s1X9+Ingbrb2mpFGDWAENXKIl7vJrtWuayAiXK4h09Mlu
yIgkcp1ZkfQS7RZGwUu0J/Gl8rTIz4mSd3r/xKbnRzzkfm8obVvUojMmLy4vyhIT
tivANcfbUbQ+4sOALMcrrr43KTJjzvJl+cQ3w4l3H2y+ZujufEYQgE1sXvvZ+yUX
+srZd5NxkJzJOSqKHv3bRa1nEol2VKJc9wi98GSa9dtkfS+9O66fqMOucQeWqnhE
qS4mTqFxAudOUZH17DFIlJqJH87Z/hqqHodz1375jUY0qvucAZIlbu268xi01lxc
EYI+1t+nHHu31r/K2A0vOQ==
`protect END_PROTECTED
