`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kvk92u5H8Mz5XYnbF7+uKUuL/MBzyJHZyq9CIO/UAS3ZERVjoq4AwMFOof5ebLiA
29FxSUReG2bWZ8WDukwaCnytLjdNv8V3oMCgG1OhzKppdQcLnxI/suaB0P3IflWf
MA671VcRIOR/TyJRWtUt4hQTCnirsXIMv7u6QrG9HeZKTvl7Hz10/DSz6Ur56C5l
5i1toNWt060soRXv34JghQBlz4A4NLz60T371ro1zdRIJjCWTq19WRFVcJaXr5M2
nbVRoxpAHNm7fPXtGMz04t2Ohzw15+kt7qOFdETwsGXLDv1nSO0cW4b4f2VDg6FE
v5BZT2WyrGBGutOrZyOZTqaZkGDXyeecT4mmsfYUR35/8xMStBN/A/pwh81b0YSY
ve4VvhLhPu240TNCI/xpqWrh8IqC1TyB2VLxpIfLvhQ=
`protect END_PROTECTED
