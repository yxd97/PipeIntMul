`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7DkBBhFfYBV8JoaHDnvt3hZvWTI0tmSZNsvtCrcTD8Qk3kdUKXKDmfaVzhBtSaCy
l6+tUlPJVdNcmrWcXmCp2ko8VqgjJjEAaE0h3/oFnsO0QhxvCLn++fbOskKraeIO
cVWf68wnYSJv2yWrdp5YHRVzQnxA3x9vMhZ2yms3CypuqfgFuhW1fB6+zIrkpYN9
wVcyqCWFnIYBOQlEGYZ0HAS6Hpx1qcxqfkFPHFewNfesptLP9waaLiTHjPN9R2v4
2H5uh0dy2NhOn2ox0Cik3U+z5x7fD4UsvE1Xpw9l12HjK8RNxa2Z78xY6stSe/Nc
9Kkv9xMS6B0pbRicHPGz/OAo451lrltZ2Kc4Zl1/r7YcUP7M6YlNGxd43AYnQmha
3UzQ0YJPeAjGvNa2eIDxxSeqQ1bTBsPYoxF5wavz7ZHAXQ2r1EsjW+1mBicPhEET
k4UKg9cWHISkqwSDdfjkDIoNFd7xTfOUMGjhHcUnxBvY9m9hKd864v5QATTW18rC
LA9OE0irDv7RMxuQq+nEr+5Ek+vFuzx36bnCbBF73MRi+WgYpMSgiZty9+FOBrK8
qVJRhPVVe/8HzBPlG+cumAlpGeJZQc3xwvv9c0ff1yrWNHhO5efAeClhaS01v7iQ
70DeCZcuPAbId2JSguj7zdyy0+tl0f9EpKtz5D8KVe6V1CwXpOZla+mteMcmqStu
4BGckpl42gyZPCF146SEbDbyZbYBBPj4yV0e5LE8xJwnPvNaTznXbSA8lq5qlbQI
F8OMdzZqR6aWKQ4QxlRC9OajuXJQ+1XG+Ap1m0WRcoBaaDRIsSiw7VajjyVfdgI8
Np2Fr+gaSS/CcriQkNF4zvAjDnWzSpJhyqwwKvi6HSZyRK0ihC+vZD17esEqlN4W
HKDN1Vu5QSgAQ++vNN9r/OXvfjk1LLZepdtFYnu9KBpQ1qLruL/a+YHXBWp78EIP
4rH9fBxh5irRacWkRH44nawEzz9/957S8L47LK9PnOAEaf7ByWvBRYVSsPxvibU4
m2493CckC4nOmpQZGGmZRa+Hx6dyL+74B3JGcWtPNQJ5VeFyEIBFeh/1cJRy2Hm3
+TzuAgzyo+UnKEsXZ7emeX4PaZbcvtsGowSW0UzHFqQAM4elrmB6MqKBpeu2bFGH
oFIDuZluAX0YptVUMv936TwYdBHkOjKQchOTaLJuIic=
`protect END_PROTECTED
