`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
woQrIznRzEJofBCKTuDT3rNtguzat7yE9ep5BR/AFN7k/T+/Q0CPqfKEizXWOzbg
0AX9CqC+VqUR6iIih0x6VCVWKpuW1tebkrJ6sNxi03u3oe66HLFUnCuAmyIeBX+K
X1D1d8ZAmkyXh6tN1tGBOAnqstS4XrwdO4M05zgUT6fnC9dWgQaO5kyYI69aIJAQ
uyaLJN6LNd2DnZeEQcevyga+pDdaYVVTpC2PA84vTCI7OQDWeFUSRJKpP9mLMZAL
GwAofb9ZlI8XEMB/VyFAAqTM6reNx/8OJx+6jDFCeOO01qcta3AE/to/oEkkrbWD
6vdlwEDoVwieL5JuUnKJ2d9jhdg61gkMJ4b7tvUl5dL4xI+VXFZw06+duLurdg75
hJGhf/hdAFVp7YWAI6M7kelSVPIuUU9ptxxPuUeYiWRgGk9W7j6lzxPciMxu+tCR
6b9oQTBlXIG6Ik0c9YXUd+dBDako+wMgQt+GW954pGDczOJYITGFJj9Er8fx/gtW
sPXhnO2n7BY+EkMHI1D9OYsOy0noqReqF9llsMLWwqOKShQourBJziYkcjzfXjdd
pBx2TszEuAmXC1O4CxsrgbAuT3NCmyfz8nA4iM2SpcGHAU7eSqYINmeHp7qS0KNY
znQb1Eg3bpUWSgdtnSLXBcO1cYdVjphNTDdiYaxgqxY=
`protect END_PROTECTED
