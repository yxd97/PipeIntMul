`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PoRhxiF05xk7J4WHFBdQBghaLRUDtnrWm3YjPn/HDX1cyEjC9adDYura18wI+qk
KKtKN4hIiBGUq2eSmBPKLGfnHYVmnzgK6fCi7RfmLiNgaDnu0bynDWkLuKVarami
L79wJmWy4Qr6tzeIzaOrDE9FmRma6vwqcxrQfq7U6BSEqk1Soj4oexE1/8vTb/3R
4RhhxO3pKz9cPRiPtgvABLi3cFa1+TWBu0ayhySweaat3C7m0jB8meAf0Ci0CraM
hCWRCn9vs56h8tfEdBPHqlc5HEE1Gw1f9EXRZ4V13gjWl+2jFrPldZhQfpeLqgES
FIKzE2TbzCWClWrfE6oyXVZerxLOjyMEqsNP58JfXgsr8dypcahUlXL6tqLtQxgS
ElNMxmduRUxvt0ik15Plze2RbWF4zSX7Cx4BZOF52dN1ZLuZ5SMoFB8o047ilTQZ
JQ0QreW0eaOKU6fKCAnnYz94k6VCP33080AAW9gTT0Xh8EuUrNctv/4xrfRmqYt5
i0/2Q4anh13CynKBDpms+oJtQA41cgN1F9+pwwJz+bi7hupEgqWvQLrFrfaiAkEV
p+k0DILnOU0YdRa0mqQVLUAFK47yFZhtpHLSAJt9Wtf6d7yiyT7x3dRVY/UTToxw
btx5e4Chl5uS/AJvmKVgeHasSuKxbhKqaIy5KGZYPbnuWt7Bl6hefmvs1lJBhmso
Rrk5Da5YfxYhdm9DRcHhuDrKJ5JB10intg+ud2fqe/naabZ55RCeBc1+lxEDmDBv
WTuA+GYypFmR8hbdLzzUQYNsDicf59khTtyx2xODWKSLrQeroAwpy/Bay9BCZYYa
P3hCcJHfHYLmWNHk51AMpXIUvV2hfM24D7ojR/jGFON13XJLh56kVhd6EUezRSCi
`protect END_PROTECTED
