`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RIH8ewJrkU//N2MRxUdhlwTxjbfBp5Pfz8cudHUo/lFC6tpk3w/iqwk23cs0x0yW
pysFh1lmt2v0rXKvj2u0SM/GqGa/HpY9D5xzfpIzFhNgoaAEHeRj9+NosH13u78Y
BW/UwFvropyHSJkE4fwvowvRTc639A3l6LDW0jAMQ9pUd0HxPpOKDMyTHEcv3AzP
SmbQbLXcL6sj/KWsI8jCq5L0E5HiVNVFP0BDthAICXA7sVxpP0ia2IYgBWhq1jOa
pyxjHLFYHTLiRGYfxWEJE52I/PediqZLHwE4CJsSZktdebkOt0eBI4ghcYmamBxQ
XOQfKTkor5mL2RAKFp9aYCKWmqCX2qCE/yqRM5lM+OK5uM5JCLpRytM7+6makK8m
GUn2DPUwyQResJVYXbMI4puOSx5UPzsfpJEvW/JU8valXRNjvTbtOU8/PClI7MzA
3YdJIg7NK21bw3juFhHP/ai/0wXdz132c063550JOqIMQGt+VhaxUMQI5gv5LR1Y
viESvE2HNEGTsfVqBz5YYmZ+AUBdQrX+M1KZ8Bxo8mHiFDclfJu3cmoAHYP+y0H6
d6DpV7UXub60N9XCNj4bxpq8y8yJhI3YBUmDPzxmhslm3wqKx+4sR4Ano5o0yVfE
4CVcf+076lifLUziD9lYRw==
`protect END_PROTECTED
