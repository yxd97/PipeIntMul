`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
frlrnOzg/Cp4/R/LpLo8lLg17fauf2aAZG2pLCeKoiV5sHH0pSE+Rz08RZSY4i0K
5NmK6mQTynZRFaFIbZ1RCOX+rb/hzjOdXJORSFadT6Iw8ckgwYhZOhkgXKU12+tw
lYBjY9UEiF2wYtDs6ThoxEp+djXWdT3BCeCSMwwWMmKH2ezvIdIvhHKh22/H2gRB
018ViA3Psf/CB+UxmoaoDuqc5IBo3p0LZa/bVaG/Hxfx4bLjEmFm6w079Fx5za57
FSg6KBgzHKwS9Z4uA4k/Q8SPYZEJsrQzJBIGSkj91vWfwBP0MqrvTjlDkZoNpldQ
OidYzaGFONCShJE1BQ985fNrocSMMkNGBFGuJSMmmdSG7akRoBJBDjAG/cRnbK3N
3aiIr+HDdSldwe0Y3SyHHpfnxn+IvFZsr+xBtaldvsPFcFucTjluRpAMKqDhmPZ7
W53F/LzCKWLKRjk0BIIW5g==
`protect END_PROTECTED
