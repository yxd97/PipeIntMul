`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRPkdwJXhc8QPxT2Uvir3dkZX81VT49R7Y53qyIuWnuYpCubO42rNsQbSqqMWJ+9
KTQDT7pdppAz1B7gdWb8rOacVw6Y/juUMKoTpOnaSXbZQ3NXamAKMciYPaP6Lqz6
Qza8YfN00kcqxtTHqbCWccabT6Nc9Y/QSOFN8chOssIy3U7zqjUiOB17IUADmfhT
Pdooamhyx2Tp8cJ+HWFl5Kv+ni0vnyb9kGkABhflwZUw0ONae9BS1T3IPlCpCEqn
NcYmQAIe/tTl0nq1mcD4RJa+Jl0MAi34ck26zSVLHpxDwj7dxvP8Rmrh3m82y5iR
quJBqad0hz52NH8jtV8lHqpmIQ6TYPLHFyUj+5MnLzlih49mdZhaxHn40xqvj76Z
M6asZKtTU8N9ts34l/nr0+9J0dMmrWsQzzy5tvqhhHToBaZjUlgZrXw4TjhPg9x/
O/mkiRuJ1sGRsZNN3wo+kSocolw/QFFdfNEaqTAXJKtmRFU2uxDGx7Icuxxs4Q9p
IcUoCoDX75JS1RySV+kolYu8f2TG46SlNM2qQpo4tryjZ9OtoCwqcvHAb/bQFlw0
7yHgVraxDxk7TcsPwX49aW67wz/lK2F12hMn+yHjxKLDuj+h3C9Wo1XHZwXGZJPP
UFaWabQ05x5IpbyyLLgatclE/P5nDM/a4givcpd5VpNlYZq2ziVjarh5Xrpvi5c5
qEJT8PgnI4zh9tL5FK5+W8M04nRdKZfW0oyCv9Ixqeahw4/JUwyi34sigjUofqQb
Z46zpcGbYQhqs1t/PI5zNnSd/hxFNn24J+u211OVvBpucdkzghoJx6lyqA3GsCzX
g8Mm+4cVCJMt91R4JFfFv4DsuHCDLv5lDvPvH6Whs4Vax9JyHZyejEIb46k36DD0
r4CsxyCTniLcCVU2zT+DY3LbK1ZGpWEnGGe4mBTWr4CFwNhhffR7hEZ6kGudglZX
gBV9Gmi4QJq+DdDSNN+3Eo0PnnuYf5wlEP+GSnAwlUWkW+f8aZbV4nRmiU3HXNB1
sx0Ssb/kSLVaPg9ZbKhu8Mgn1vHC3rmgW4eY73QD9FpmJNkn8jHvDc6D2SaTOAmT
/M8isGwWAr1p8tpBOyBkSM1HWSm71rVcrwdaCtH34tl5JSMCb4EwivlRSkoPuXoA
Z+4j0oTb8TsD8b65ljpiduVhL4F3aq9ePXUGBRlBW1hIFFB7NgSEEmRR7eEPe9dU
cFRDuzHUO0wNhD3vbXcNDS5Uxf8KAK842/VwJkS0hWNpgXMsrPv4+e1Erf1xfNbu
5tytFmCHQJ4lRMVrW3i50485wbKNyCqHodlT+0aSSRUB9tYhOkPdq0Qees3BsZfq
awyMySe34roGQV2KrAdH7EOmFtsgra8pJKKfZy/xUJeStnTY5jq44sZEbloywqsM
Tq8mhRP3CFO3qoVZHWAvKLvQU2lKuyIYodgFJkYP1pEbAqFQizmce2YHiv/Xahrm
z2d2t2ifhfjA6B0HNxyK0VLaY4LfOAmBDIA17cOjDCVFJoDoll4oQHhvr5HagNLS
d+SFrY4StuaBFXep4SIT+Uo8S9xc7tlf1enpfb5l28L0HcnSIAYmevoPxLws5fI1
o2E/nCErWA0qC2I3KmVgPCs219Jj6HPb4UltW6oQJQ0WNUH7BFahhm+nvNQkXtuh
kmeP03qVSS2/6bJ1yx27V0w754UBr8/OR+IsvQimw+1i0frByqLz6ifomlJBGEGw
k4LePnnFPywjMyPukiMis/WdLQgvr7cm1pZLElIXJK8lazunHlj/kBb/Cwk+0TS9
hx+Ep2dqeACftHXOVZxqE4kGaVEL49WGoSOkpFuNwHmIiWiD5O18wRrNmoSG5QhO
ET5vCnQjvQWk3BXY85zTE9EcTu8Jrw0lB5OKOg0cRvYh7nygT9m9AUEPYQT4b/53
e/DpXCmAY4ZZIhJTcs/nrJ5bvsIdPqUmzELtdEXuh1mncrEe0a5fDRZ9vcaTNsi6
RZw643kEhxC5E8VkqLyuvYfzr115P57Ci9acQpacCWlugjQ1aY6eyrml/SelBcy3
t9pvuQPTEMLz1etnx/FtZc5DBrVEVqeS63PLAHsQIeo/YHQzmCJ0HwcKNndB21mu
D0W7PHXdqiMeVoVTQbc3p0oW3tSKnhjCJNcZ7wnxXY6/iBK50k0z93YnwVHeNb8P
6tMEy9VjCaovYaM9UeE3CqVXutquzxuH9Uv6/rgI1OUsBWio3pmAffpUeBiuuRNW
7WqtLeXlk2U5yN319qYgpw+8x1o8e21efIh3wP2SdS8Ic1PRBLMsR4C3Fe+lKqAl
TDut7Wf0wqsEL3xR20XxLzAumESrhggDP0KguBZ8AUP1hCOATEEIZ93be0wjwP2v
Yg/x/YaQ8BC0F8p5UsId5yVZufRWJNoGXANPkBs0Xox7yvjCaQSGdk60tKZDnwTR
ydQiPo5BGD2opS24s/BsTzK6+obezrvgBIo6KXv1Kg2wRvR5nNlr3grgvwIUhprM
5mm32ik247kcENYNy+ClkwugVqHIX50mDv7e57cxvxWLvdMnCiKA3AVlJNKda6X2
68EVe1Qc0jswLEpmzzjPi2Q/Nda0z6CDRAS6Y3uD+C+f5524UmTVUVkdgWEUlMqb
O7lMZFjd4D2umYNWeGavH0VU4I9HL1IwCo8N8UHC1BHu1lXxrCb4f8ESGX6E/88d
sZVbC+IgolmUlAyeBz8KELXmoSaCoIqzUiykhGyjuE5jZDDG5IhswFz1YQOhtGDh
dwB1ZuUmbJyBvoohDsWU/tjAe9XT4wggK3g/HiKKlJog53mV5WjlXBgDlVGLvfjx
Dk/9CRSijxx37bcHDwXDc8N916oZGVeh9ULavdpWjt5RkjIs4RNB3H2HYH1g+on3
eDcYDalNKIWKXwzl7uNLcMzdlgA9ugVlDd9inKHYfSRkbdvA4qlCQzUN+hkWgNf1
IUyART4mK5U8pPUp308u9rxebDXWlgWJRBEwFV6eEPO9jOJIRnEgyblU/GwOtUpi
Hf1uUlsJSvIUW0ycgGQAS57E7dyjXPLKtIf7VG4fC4JCEF3jyWPa+/7eP1vxHGxF
alP1h9jhj6yr1JMLg6qXPDcmNxHRpcdEjuuGvwFbpgMFn3KLZASy5rZUbg1bdzKK
4uk/aj95MvkxrJmNZGiQXhdRAPeJsN0dQscZCrRWh/tiQkZVJdejR5rMHMbhXHN4
gFTDrs63smrPKasuUObQM0kh9V+gGyAMkE4B7r67u3hIP2ah24PBkClPHm2jK4kQ
aCFJSMmhqZ6Kt5tVS+jzi0qwej6YRmeylVgnSkVNvVz9B8IgILJYcQjB/mqUQ4s1
boPK4L4Lr0l82sIAkIItF07Fwg5SDeZzn6nLMDGavogqwxK31QPYPFZ6uWmJz7xk
k7A58zHaMZ8Dq3X9JS9kCYeslkL9jsy3d5I03K5cF+T45xd0y9hJoTPE9OmeN78d
GJENQISNH45QNqKPrO1mGYb53cagaSRNrI4Fe45dh99jFqX/mIaC5EtyI5LG6lUP
xcs/6sqUW29chIPFNHOVN2txws7ea2kocOYkYphRVlNjyrxrVq8MtmpaapUHSPHq
x6SavGORR1fr5ZjR8zhIACiKZIbQkd4w3BHQwwN5M5kXFgZJzMAMUL+sWNp4jfdr
yypypv7Ium4OgObtXz6kKCr3fMm8Cs1+uGbLqxDQYExLioU1Hg3YpokO2sOXtx2G
Y5GqqzDL/fuEhddjWYpWBBiFqJNZgwZmuHTiDZI5qHTJ0gsUkdVgXy1QMICT72A7
LHwVjRj87+chyngeodNyVz5GXDyKTELpFpDKZYza6T4O5lUMYj8s5L0bEFMuknnN
6CrCmEVPec+cpgEMpDhMrLWsRpuTDlXjwJhUb07cSgvmYmHOnzIvVa25OdvGc2Ae
IkIMKHHwjzHNsAul0Oj2i+5r+YcOCKSk9heXRsE+WCXT8zctthTIBnNPTLtw/rMq
dpi18WBiciACONSe7ucY7f6x328otv4+BlzVLezwoRIgFouIbTTRG1rBjuq029dt
mDKJMI+vS7yFxCUmbP6KPqmYcGTJPECue7s6ywiHeLMy+usaTdYDEpDDRuUs+T7N
nnso7QWm4YsqNLHmrjFsUHEam869vywI8ZAplJwZmSA0OYHbJZKHBqFNIcs8Dv1o
6Y3beA1tirur+rtZOZvbDe1ITj+6hkB+9wbz36DfX86MfyHkcjQr7b9ioDpz0w/f
yEF1T+WFHtiULtvWKPD9ZCZpiVHng/Po0PZ07jjrcR1qR/kU6ckDigtZclQYyu+i
keGgL+pGyv3KUCzvIQohJ80cSMIB6nJKgsx7dYwZksAKLnq4Mnix87ueSsGZFQt4
1UvOP/3NRyw3ihzcuZDp6Kgqt2Dgj2SRO2nvliKuAVvViB00p9RUHaWvyKG1auZX
bYKoxfaNZYoaotp7yQoT+fT9XEHY/eNM5eTGQNulXIney+1Mh7Invan37HBE5stj
+o/M6SxmiinhMs6XSXDkLD+ncvbim9yPKfGh2gO4rp3+qrT4eysAs9mwUfFBICKk
0EZBy/5ZEWCCBa9xOL6Csz2hqCvCYAvJ2VJdEyn+4Yqg07VPyl7JS3I+oQQBnOB9
FasPrBoK1lYn4jRuyXe06ZXNA1/l8Bhv7mHnBzwj8A98USJezo1BY9cXDUGGykdp
GU7ykbNUUhAhU+f7YxZEKu3N/vvdkZ/U+2bAzcuT19EPXhvPtCTnf35RWWVMoIjm
B80BBvM3Ts5eCBFrJ8+Nx5PdOXeJYjnaaydmxIaub9Te9AgsxnuVyUfQLKpjdOcn
3oCCqK3wEO5TrpDMR10B99gYJsYnWYP+7TkeRQ2Dkw1vKC7X7GGS/mky4xUpmcRY
Ux/pOTRjiClF87ALZC+U9EnLUtuuC8T+xxeqlSXeSBP2Dt/tqEZbs29l3yRpnCQb
+PSmoOv6qkTZnkRyssMweDl58LVjf3tlx/OXqV/4efcuDNoyGZVbxWW4lh8qu/6O
dRV4opKx5SDcIh5DQ3GstjO5OoeqlgwDnMaOLIQbdXMNcV/7H+KVmPz7YOFITGA7
lsoZlLXVs2mrFAMfdzUf3XL1Dbm1IG7ILgbjYaUBMYfMC47sc8gbfuS7mlriGmr2
`protect END_PROTECTED
