`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iX6ATHLHdurjNrx+iKs6cm2JowydjVm5joQPAhFsIaAHPmv5MZjfWDiX+6QYiCJO
G4iF/yjndwzessuoawVTG0xxMbFM2ICew5McODumGZK1NIYPBxHZVcuSScbGqvea
g0HrU1PGFT/ct5xPXMXuSaaqJ/Da4LoZohrXDymLHj+7mWMGRWhYBPPzwSqbr2r6
642Tubz1SrGo9AtjNDbqHhTM6VS1ChRE6eZ7g3ULjZyRnwOkdZJkwg0abPjp5TRq
I8FarhImR8yg2atyitwfsgVRNSf7Do8MA88QTaq8/7X+gr7xpiD23B7J9urkNus9
7jy3teAwYAeBOnSph5WyAoJ9y161Zl4c2rH9y+3AwNdCkN6Yd6Tc3d0pSHupEf6b
RIFz0xtFEz3+yp6GO+7QZYlFDuXawQLc7IILzjOxGTLuAvk1xC0XkAe1nx0W2fFq
UlqzLecBaTF7eJHjqwNn7QAM9rGeNvsF9L/bR5KEADUbWlrMkjP9dtaeLrUPlmq2
gTxU+AGET5BY65RTuWhrGzhqvQEw0FbYcAiMyOEqSFfd4T6SbEMyqEohQNhcMH4g
Y/6COCfH0UcMTk/6wHhPL136LHwsKZ+VnbrBQT9ZXsyGZ7DNMpuyoNCdn2yuORgd
ABb4Q1nQ3O3WxUhUcu0LMrOfa1mKMix/z+6vUfi6IHqg5C9oUGBZ2SluL53Y2Dty
0fYrcN0GI3fm+RXumdEaOVVxD4TK6+CFnOji6UXNaMpc2BoDKXBXlNOq2pxmr4G5
1yBpgq7JLFIMfaP/uO4J5kMLE62E6FRQf5F9u4zPDUB9gwsL1jUvc8vsyBx3PR/X
wa5gHid7h5IfAuK4+c7tThqHkDwQIpLciXdBTVcMeYfVd+Fv9ISVGltOkxsQoLK6
27phtsb9NUL+VHUgJycFOM8yrnPRLeEPgtnyJLttqV2rzq2s1inxr7oRmBgpR5sr
QpdsAK7an4jv9zcgV4k3K5icK9UUbivpffW4mzEEx6qZlGnrvE2f65CMOo3y4K/u
IEuuEjOyk+UqIeo7Ll+DuLkfIkBzu2x2GZxRiqwxusQ=
`protect END_PROTECTED
