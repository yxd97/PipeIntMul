`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9To4NmOM2NfqNChjWPOtL/qp944TbSTATqNwguXT59amsmETg07LZ4tHG3+yS17
g7paKC4CTn5GwIddAM32W8LITGntjQpnklCe02VKWZxLmk3/AFm65OlqxJPp2Kcl
hdLOOn++Y1dIGVEtDYZ6AJefH+Zi7ZK+p2W0IH5ltuYnq1RImRIWg/LPBR05TSqs
8IbyRjWAwLt1ZOj2VQSPlVpoFYuxkVKix3XfS6vYX2kgZ/DT7VXRq1T1nHCQesX4
Y1QhSulPGklYrNRXCYhPTykwj6Jhgcx163b7dhSY23LLlbmzjJfiHRGKKF0E125h
iUFvcAE679cIn/PBoQL3LZdYcOoEr6Pzan9cXOYm1tmYTYrI1yvp+8BfpEi3Jz3n
FvgpEUo9X0/8j/wARIlebPcEal3bkDrXgt6xi4GO5CM=
`protect END_PROTECTED
