`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOh3C/wkSGBnV4qQFiARjLg+fhPSi0nP235gv7rEdz+12dudS9JGUtWiNznXzRNk
+dzG5pkOUo+ZY8dN5hOTnCo6Jhh/s7MaJNSiXwa2EsfScjPtVeKyC0EeNHSgo52/
WxLPqhSgiGpSprVMOtJuvYXuJHacAHMuDF6W0Bj6SUXvwsFgjKk2ATwyo5z1IQ+0
vZm+EAt8t5ug83hp54Dlk0TF0POeF1X8JSbzTC+BPncdrelCUZKommfAZyd10/w9
Pmo6CrzV1a/MN7JSRF14vQWnAKwvpt303O0WK987+WAXtOlD3EHzmqZwdQ9rEN+t
1wwi+/fr8XN0xTP3WwU78yCMrK9X9B7WqHtTnfhOsboIsolmocOTXKZxGJ6rvMjn
aTUhLUKFeNetvKvCXg8qEL3yIvCRMedirzpPqtuzAXIPbvsCWp7gbt3KQ24cpq0c
p+m2Ofd3gP/s4HvDLoq3OzdWORpRbNZndMU1sUZfF3K7+5zlAIwNY48iuyOat0cL
I3Xo51uEjQry91n1Ett6U9krzw8Y/XeqFhmOE42tyBaeHhzx7Oru0X7b+g68M3cn
jKlAqBiZ6RFJYLpF861ddpDYYaImZJctjepAMhQzDTtnUA9+ZH8T7b8cW+Wg+kZl
j/W7JAt6ablYlMXoKZHQnZ6fhSgDaUW8zrPg7QMiEAn2HQyvQGX+Gf7vamyevzq8
fsI9TwwKe+0/oXXn/pTeUCVh761t6lIBkO8oF01L4wJRsQA9sGCagBLENADnxZEI
2nrxAB6undfI9q6BA0b4CXr75/3/GfXuZ0URxgxhGsYBANLRkp0i++jqt4BgrE2Y
ZVU8OZJ6Z6eRTWipkiZob8Wmni+upv/LAyjym+PmYMn23RF3BLFV9WB1VdMjANwt
FswBAQm7G7tw0XFNNlIkbVkbUVh4XCZJRDqRTWG01EXugoRJ3PhL9vUpLjjKYU+p
DAvs6WL4QiIH38LZNtkHKHe03Z9EAIFT9UMBGPNfTISJ+MDA8+TKRTSmsdjh7YbK
rvUwBygqR1R/l7ZY8dypzSDSE+wudAZp3TyaQuLIHxkXLz8hhV7SOh3Ga9xbMZXz
N12pDkRzhHZdQeDohqjIqvJOqLvG5u6RY4yBueTAWNbjkYXB52EqNPK2ISnM1tHO
v0qS1/PQ9VmvTMQNfKqIy7UDqrdsAZ9SoeOkT/CtZ7j22NDb2XfXInGi57sTNQZj
/lITd1qXJC98gVe1raW+DzMgur11usMnNfMVd+yDE+2cSEL89jtwbum0E9U5wsDl
vUshzKvXsGa2YNuuKqBgLNKvGf3F3oEekmHnkFZdROBaZbgNHLZw63/eIEjkAM+z
BZMBuYEJUfX6iP17LuHCzKVpry+835P0OJdxQSFGrNV79C+aQxCcT13bVtdbvWTQ
IYPk+JTDvmbo/YGl7Xm6Ifuay0rseUdzclPtF1kxXTtlPb8xt/8gL5xhb38ZbzF1
WW+3+vJCx4H0UncFjJaY88od/DCwmu/ljum/2+QC63TaoEVPJpV74qdomHrhMWm7
0bFHMzCt8JCp0AWDdBpOObsR31xMFZTihbkMjxvCmRPSrztgLmdn8wNkdYyV+7+J
KuWlPQS4vWD8Fs0KagNUREzPosi6g47sKLysEGa7zAdvcU4ke5jW0hPOAFR9uqIS
K+z/3j28roRguAh0bFx1qGzhxtyQ2u8XUbgqdwnlUCKrfbISIy/3SJqJLRfxGr6k
Q0b9Yb/LyoCSLe37Wc9FBsJ8oBMzYiM6s3N7Ydt6zWkoq9jxzy07vgrkr5Fu6Qjy
2soEL+F4i1nAurmWL2pr3QNJHyEUIllNg3v8jvFEbTUUychWJtjs2s0CFVUQYPxS
16cXHyUCCTBNQ067qyW6l4SW2C46JrQhtqCc9mveTIlRZu0X+0NX9sHpSrgQf32S
FN7qCkBbgtJBawoVWMJna507k9jNT3DE9xtPMn9w7HO5t4KsO0OKXsfF31BsNyd+
nz6NxhdK1ej09tlgQ+69fFsROu41i0JQ4r2w8mm2EBAdufej7wbLAs/ujWBkR70z
11cuifZUS8ceNMLjIqqG6FFQZllvNSk43OnLqCN6upbE+UyMHAJ4JGS7CQiM+MXB
SI2++jsUUL8yaIo8TVNHD/SaqJpePOzTKhRG8e4swngryXU3EEtsWQmIO8DhaHx4
3wZXK1OaVVEg9VL5gjGQjmKD/b9cWGltcpScc90Ssz94ozD+D5rdSofEkSDNRGY0
/VCmb85m3fkstE6Y2OPiVyiAuy0kh9QkFFobjymzsr0=
`protect END_PROTECTED
