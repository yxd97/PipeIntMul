`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/P79ZteXEFE1aAG/D2aPOQopdJxLLl9fx2PcczZNRKW2wxlIrPtijLhWIE8iEX6q
MR3SsZwMazTLGYWrbdjpYkIEW9bLhvbvPC7WNrj/M+H2tXAAtXKTA60UoWnGdil2
IfeuJQ4GuMZJGtTYTM0qJ0D97IqHvSfMe4LanBf1kK9ai2fepntx/pM7jvdadIAt
+qftgu6AHJAcL4OKpqQ9eLL4DL6wVW03wXs+453L/1NQzLNDookFfgfO0upA7ptb
RMsmjS5zW5aW7bWV2rVtFmnMlDxMHuy1NU2WDfWM4S5hM9sTMXd6dUNbmTz2uQxu
aVkcoz9vl0/d8BRxCztE73MwqgLKgJDauGbs5RDMLJnHW+P/XIMshHFaZKNmbCPR
N4pWcs4TJJ+HtUSc2XaALKHWSDkhyveb60D56Sl6Z+18BauwBuXptOsa5AUjDgtg
`protect END_PROTECTED
