`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NczfKySh2fUU+rOM/MFaCosRAf792qcRQ/OVBi/ztot28rAayn2tdJB3NrJx0Z09
73hmDRzKZAqOGj/w9fa/53wNjUQbItOZelf/teOR2oL5K6350+qpZGcHlab4h1v5
FEE9v3d1pS0uF3tUs2FWauQwEVqeSvEJqweKqSeS3GzJUcal8n5ZNLHo6ZbOQW8B
4Hs7qbOb/Fm5xOdt5PLOoczBmFVWo41YCwNXTXzSpM3SU28snn8rDmVH5KeB9Y5K
ID9O7E/0gY+hHNwGGVoqjl6mPIlYaaRNf6wZf0tZFW3IWPtR0SSeS/1zpZVweibI
B4b97xg3swfd3rjyU+j2Yi0C8sP9AffhIF/o9GnR8zsQUQkzVGvTT3Wc7gVPbSXo
Ma8688Siabh/KjtE6FUCwlRpTpTzTc5FNo4fpbM3rY1uTdpBo19YjRU3Lu4JkRwd
pBwNMhfcrd1IVzNlQGfpBd3zgHBflkzotRFMISWa3+w=
`protect END_PROTECTED
