`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tROSzzxFqzUlbYk92jn2qyZXkXnOL9e6CdOAKNLECfX6D8wmVvPJahnB4k3oneGs
A4cNoLB0MhXNrRS/1SpZTMTgV1dkKnGHdXlWga5v/UcD6qJx2waZF+oDQk+jKaLU
ReiWI2nlC1ZCGjmrL0NEW8HUDzy1p3PXIiJ4/dJQa7NLY/Zft6oygOjbY8PF832v
C/vUQL0AuQpL2UqiK5Q2SrRJfRsIzQvxa5eNlXyMFm5NXtPgl6YG+wEPiVXH1yGx
bpkji2/XP+i0N1Adv9pmXl88cU6O5VGA5DPpPZGb87FUst+0lmuOhnoQLVTy6bIu
q6XW9kTdngSi+UnHJnMcWdiYI3c7AhGRdfY9Rj9bPhezwh4b1gS2riI72jeKU+hB
wJ59FlPfdBfdYzvb5/l9fA==
`protect END_PROTECTED
