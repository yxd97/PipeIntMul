`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Ze/gzAtUuJvPSuB3Qg9Iofxif0oBZiA6CYGnp0NQMpfSGjvvTfFApPJsJeMdaG0
o7csa+t+814gInVStHPUHG6+HTvHkCNLC+SKawbW9v66v/OEEM1FrFkPkbCUaMTU
ix2e8Uuv4/6DhMNzNfzPBkyvtkyoh7H1bSFRsVKKGz4Qh6E/fFOhMpY+zXC0ICuT
I3otsTikexWKfFUXzfAyzLPFOvFKU5q9p82CzCji4hm+SG6+fWwNoBpBU5MKUBXL
d+pVpHs2acZPW3i5TdYEcnXfjEskfdvMCy7Thza4yTzaBdHCor68nq3ezZW1/+xp
tPepLbPzrRd2oovc3M4nDYxoEsoI/xSpnl4AFi+u/f5IKMCWG/TOcqgTimCIcCbI
lkFftaOjyW9/SQ1ly2JgAyfD1PHKTZ+ji3hglRdclZMCnECMopZ+BWbxhJBO3ehk
yid79src1xLW4GGo/FNp9685s3mOF2oGQI4Q+JJsZddPS8l6GRmK8HYPn2HR5Of9
irO/ZQLyuVCb9j1SF4+NYdF8JIbcUP3KAVP+yItGuphvcdjp6hu1lGM1GCnOpgJY
DCwT3FKF3d9V4H9r/+UvZZKzGtxUQVE6DnUt/RSbR7NonKW6lK7BgmRUVkEDH3YT
OM+lHrUq1RTk5Arvcr6Zy56cWPmH556R3oIvmOzs0npv0sG8Q0Qztt6ZnzHdqSKP
bD8IzgSk1gTNKiCXdHmSqmGu0FCM7gtDqm8gX0hJcf7GSBOxsvqVrzSZ7xJhZvdv
80Bw5sfMZMetZKOJFh1LJYZXMmsUXOLLtvrdrdQ7qn0fDXVqVxAaAuvHvW2vpqdp
rzEwpEKsRgrguJaE7Vo6r0onpnagWPFLbU48f80jDPg=
`protect END_PROTECTED
