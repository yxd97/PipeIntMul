`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sWmm1paeaMhqMrgVFqcr1jWIb+4x+VrmvXuPXYfP9761bO4apzeTvcJMynqqvRNE
GPYA4wXmV6Gx2FniEpN35enpBiT4sgUNok/F+uvuKy4yrNKEEJzAk8giG121BdWT
itpDkFa4ZD9IFwOmlKO7qfA7Ih4OWDOfdP6GJDdk4TR9lmLjqGlq7ZWEIxC+v5ra
MDUSXyIAFupGOhEQKhobawMdhD74N1R8yCj1UYlW0y4r9h72xg5BqAbKxcSbyssM
f/DX3vA034MUYWTWU5gNy9OTaV3fBlk4bEowlv4JSn6JhbtiVV/IjG9exsQReWME
6hMp2L7m+7VM+vC3AT0EeEACEZQCIJ6yXl0Hsz4CmRh7jWIkUqBMX/3YewImOSVR
l4zZijwJvQNXMradTFidSLJMnaTtGM5bfbEg6qeU/KM=
`protect END_PROTECTED
