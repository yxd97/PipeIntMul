`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d/O7jnbQm6PSnBuyxgpcsz1gWFn14av6bp+6XkcHFeEaVcPTAFhMAfGinMJE3Y0h
V36jjOqE5i6NfIiNo9z5Z9Ski/OzsRKdEhuHS1aWKLoSiZd2SpPvEFehFi0h35B5
LwylCX0e4oOrDIYtvuRw3CZ7Hvimx+b+AuujZQr18IfUD7C5D7a2OeYg0y849VxU
n5Nmnl45NRXnVJ9f0URgX+d78tYM/xiUSXHi74XAjOmrai4V4GMDjfeR0aI+zUTO
I37x0mzYQw6660R7vS9+mw==
`protect END_PROTECTED
