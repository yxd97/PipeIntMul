`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zVtetteiYSe7Jk5qYJu7mQ78Zy2lmnKJ8c6uTjaQ5od5oFGWnAyhnqKVQdBdfwWZ
oiF82Iag3SCmFEcm7U2rfJ5TuFbCkapB2qc5YNktQtY2zBFyMMwb4X/rOLlFr4Tb
Em6hcnlXQfvR9jhX7MzxRKt5lG1Q4jwUatJqQ0MOkBu6uGEG47mOme6ZVjDJecCs
suNI8Zj7U+GQ07K3jaU5RaRK4ztWRjD7rKaja1RBwjscbhQqU2jGg1BpdkNMkT7j
4LY0VaD8JMpD+wJP/Nfo1VTCHu8FcPfmIplVtqvDq2FuSoy1XvRNfKcWJFoKAF9O
P91WBS8Jv3T6FMMfkCrYDfsG6zfRXcDxZexIUUKUqKV+jYCjOYfM7B4Vc5mzomI0
HPVHicy1qd5GEO9hi/1QYreVL91EuuWtizxK0plX9FxXNclVuy2Z2KH/F0E4/Y1o
ICPNQ2eJEncR7Qu3aAlJRt7TacXjvkRz3G0CkbmdXspM2v/Z8ol8O0pNKurr5Jn5
LpKKFpWLeKFqk4gkSH4ncOihDWpL3S6L7yoCxcyKowUGcXgOFHpbMXpWs9lBmFpl
wTz2JW0L3JFnZTqv56KjgI7F/t8hTMdKM3nulwSFEz03owB5gjwTLZ7pglRsU0bp
JL4qqcaAyOkoE0EgLA+AkylEc4Nf11az7pp1a1Pa+2yTRuAYYoNi+effF7JqJfuU
XSUrr5prEsJjFI1a8DyWL3N1ohkX4njWzsz+xLmD6MQhwjDIWCRrJdd5LLoVYrUh
4zGZYu+B32a1PeMo5wzPXXQhDzoOidApim9J5mCamCziYliiNKmlQQqZ2otGvFZK
rANkprm81nUhMu2EdlHTohOMSZrEiucHGjtQGjK8VXGkNJPDV9U1zrR0e31Z2BTm
gZ56NLM6MJoPhpIlNZy1R8vNQEC++EZLU45vrCh4JMFtu6y/kmma/C3uXRjCvezk
kotJhF32cxHW820m+y6Tv4yWRLpxr0Jh0C0Pr60mE8r/hF8JOsQcXPa4QGXQUEkL
k3qWhDfJFyhGZciVErhXYlv9tyo8o3sGHHEqkPz4J4jJFRfv2i+r92jldDWhYTch
ZjeriLDDp9vgz54xQ1RxzNMg3zJYjwccbuOd8fu4PAoJNDcNlO4T88AeGfyRS868
fSv0x3GhOXzkYEy2tfPt55khhqO2tXbu5z4T4d7EI+eOMjlf2H3G+IfLayVM/KLU
tuS4KClwM0GhukYEatXzlsHr2Ve1+M+wu6lnUkqn/4UQTukpic5dOmUn3vuVEAtg
zGgwMSfeLw1tXZvo+FqLvPb6UiTjnRILP1qIKq5l1W2H17/VbiWCpnqkE/EAhDsK
vCN6EFjlcswwL6v/wjwZ4gRzwNNXModFrmK/7FHXjSHmnWBzLTLS0NANvp5X626k
7lkDAoKbqsZc7WIgyojb68pk4ez8iLpptu/5GwPRr135+TdIuzuEgYyGS29ELFXA
5Lst7Q4PgiiH3JbQiB2yG34/oSZaaymmdpeBvtDADv9NTddNZsNs45AeBPNzBJGK
MnUbhEL0Z6VkMsnKN1OcV8mUWe63KZrC3GiSa8D5VMtHTWhjiAQKhcwIR9grkdws
fbmlFUu5e75uDn0I9Ck2Wmnb/gs62rFkEXyEK8uTf+Ywi+ktOkYOK7kId+k0573L
9dsKasaILjNc8aSci5UTjS7o8Tdo2R0j8anSJiGp4frrYFP+eiIw7rP0o9ga0gLc
k64lisK1axpaAC0xiseKl0VP2y+EUv5J4Jk3QbUUMIeLV3fnrWGKqJ+oysAvyu+r
ObFsKzO53ERPgXfOj3VlDo54e9Kb3rqSd5fnUXqGgvTUPDyxYBmCV8xUBpYLy2ex
vyWoB1Pg789ub6noqhlmI10VD+swjXGB8U66muIaRBM80Uod0hWxhkxBek1+1Hzw
umzXq+275Z8ds+U3dlrQAlRcSKEqpPHCylZrI3jaAGRgRMDhxYavKjTqiiPtCKOu
k+Du+/Vvb62ljdCz5Q+a3RRH+HLlZBw1civrszC13yr/SimN9c+fb2X2tXB8+4vg
njy5s24DT/Sv6TxmdcG6Sr2AItj5ECXAzCeWRh8g5y2sRUuquiQSa8R+v8xcKUNg
0Fw7qFSWdOOfone/wkTUS3YgZp9S3s4tGZJXPjTfRw/qjK0JQltM0lUCmV7iKukm
1qYekse7jcmj+ERnteBPfEesSje7Gizq1ogGTKfNnr+WR7uFU1j6ZunLhHch0qkY
9LCDdU9WChsjFRwZGLjNqVz+nWrHngwZfE3iONjoAOro4JDHyuqDUE5XdZW54aTY
CbycMDO1BvHiLdbyvZn7ilAPo2JDWgmh+DGisl4Uspw/QSSCnk4m4EvnhtViQIzT
aFiduOaVEbzNbT2oP47WBQ/vUzDagH9uMbgWhwq7xrcIEN/i7i5k+MRDwJog/5n9
P7hn3ujG2/1JVYgw/AsyEtX0sHw+ttpoJSa9ybLeUHO7bsYHidGhhGSQbS9BVYLh
E2k8M4LNC+DW/yZriSk5suvQ/YiB2eWP6Wu5RD79z7QcFGml6pmNERVHrN/k7Nv+
029gYPplJGYW1h3mqTDShT6tjhthJivQemM55dJAiEeq0n6bL+TkZ19NAl1dml08
UUrm2gAxks587vazKgdirz/8lHaAp44w5yxUf8ZooJiNTR3GTyN6I/tgkrEjTzMq
HqCe8Ua20eEUDqeDC4pbMrNT4Vi/DvoXkG7rgb9v3p0mKjCVuaEV5xRMtaHdCZ7F
iq7cNSa+eRS9fhMrFviv76evpHlR5tiicZUaqWOUW9twx9ombBP+5DHabbNkGjf+
IJpkU1QI9Hd/4NNunTDwv+oo6zxbcbZo4uFskZjkOGv+jfyJr9cyKCeB8oRJRg/u
GxWafqxM2QUzn6UalOiD7C5kWa5Qb4Wv2DpYooeMBiseV9FIBckzVJ4V/HZb+86Z
9jAMqWC3FgFchbaNn0h1bZNNQPdAfe9UpkLmdEI/kTIJ5flAwTPJbbUdtT0U+mQa
KUZzVTiAHXCRUeWP2CVM/6ywkX/HJCtEHzZ/+Iiv8lfcCSAYokVfOX9R0zrtcQU0
Ad9oKwA521XD/+WcPO1joZ3FAkskCwnyUL4vfuMj4PRWTNhK6BlQ7gTaIDz7z0vc
VDf/JD3XQ7OyaKL5U2lSJhUzmi0Xht8vfqvsy43ywOEgF+Y0zd6Ig5QGr+Rp0vTm
5d/+yviiF34zEykaK8X6NlcsdFjbuJYRSFK0SNzrSTbLXs2a3NMj5DL3+fC8PFYZ
5nrgk2+XRo+XpKUAm0qWbKIi3slZ7iwicxXniuEpvCOMJtiPxf/gFzWTGkVAMaN3
Vr4jjrHrvrFt9qq/itePeo5bf1HUOCfiSMymvh1Hg4+bXa/oMu1yI1EjaqjVgF1p
SCGFCD6Ca5bpLggoiWWVrQS7ka3EwDg6F41ZKtR0IdlUZE3QvKEcnwdsdw41+3yj
GdqaH/Y/q8weS3hBHWwAz3jLHt32dOdasyX0uMhSrYGCGAO+h/qTIq2KDnpW6N+D
c4h/9G/5owWbOMhSUe9G7WQgkFrkZHxsAUZxl37496wPyNAaNS7sOX5iWdkab6fu
LV3Bui3/J4VdO8TXDHGdEIhL8EikPg+Rv9jdElKc01HV1Y2chzsh+SZWYOF8Q2tr
6r2vZ3/iwGHrHcNSL5KK/VC0UqqaWr2+VRgF8fXk98UIqPgZAAXHys6ZEhQBExG5
IMaZli1b2d7QGxaRh3NSNUUCmtyXRrYPKSuPV1LbNH20a9fgVISmP1u5+fXEx7Mg
5B3OnsZEEo945Xl8uvx9u4TTrr6i1h3lvsvfCh3meha2i0KDG+ExI87hzILRydTP
toVTeDzQG6SpzjzWR/2RrVJeqIwouWZ1xddOtflfsiZdVFY4SXKOVmmidEwnxE9K
653XFXRFhzaq8ltna9t9Y7O89eE2jiR6xMalEKIIaQXJSKj24xSu6t+5kwlgVBfw
9JOz5FR6yV1GebQHngfQZxsVSPJnDZ5By80ErwL/1mjxS83CRIOeToF/sQBuEAks
2rgr67O7tsStEP2DWs1GLwir0n5zlOnk87g6AwP0d3R/BCzUi6Q9JPhjMsuOBqvd
ieUFDHOi9cmAkoOj0Fdx6LSlaa3GrOmowCoFPzXxy1Ipwexxh2kSKNPgui8n0X+/
numC/aH7+C6ya6Dm4IU7o/of79dsD35uPF6GML20+5Z9zuHX63rJ0U9yCF95koZr
Fgnin1Tdjglx6jQgd2/f/bEmv3dl1ylD0XEjUH2LBiCQ3tn/fHw+WQ7VhTYgoJyn
OR9axLvkcg6MaZ5r18w0sW8xisR8hILdrnzGW4XYZ5tLoNCbH04XdAjRMqikFV+q
J1EkxMfZpYp+y+4tdU+6vynNGZaqnUKCaVRzZeFkgHYMKRZz9hvO2RSRn7/zOoC6
hZrrvBryVGraViR9LDJFMJUh6W67e4n5cs1G39NwKWCWcY5TpEs2nIgMvN46LCrq
LLlqkqgBbY3HFD4DAOfttgo0ESVHJNmExIvPu3gAlNzpuz4yDQ2sTKu8KZ3N/QBZ
2vj0kW54vcN4Qye8lw8AcHoIC0gHWYMIk1yMvnGCDo3WLTktMzWjbYynnPEVcGvy
sfiy2rO4AsOVHyN9nMqQr8ZEuIcmKuvZRRNLgwKJOQa1kACm3HHxYRpQ96xRiIOX
wrCtTZKeCfc1ho+P9b3FrY8WmIROsO2nwzXrhCPa3o9GhQg3CV+/wREFw238k9zp
5CQnd5nF1Jut0eIxcwmRc33widkMH8o1mglERBmwpcCE7DYegEpNWwtTWkY48eHn
sIZqi1XssIXu0t/UFUHa80QJ2ooF0Rc05E+YckfC7tUcKkUmyYXUEOwx7dVMnaqY
90RmLqZcV/mJ4lRcGYX7GJatONpRqT5xeKi9x5PKIz2X2d0VMUMyqBC/smt5it54
sNm04oaDpBeDlZ58Hkv2MA81wB1z1CyyjFSi/xi1Ct/ob6a3ydqDG/82vXAzIW8I
sc7UrhsUyP6sn+FEoMKmuJXFyCVajIKIP9l1ZFdk2UJrMsYtEs48+EoGR3ssJ+ul
mTFNR7Vs87MhuCr4UcC4XOXxwbMeAF0F80+qTP6GSTTP+kIaDdoIKM5JC5ikCpME
2h2Ujfk1VBJjC/nJyRAR66MKDee+noRmdaDnFFd0jdvGE/dJxzc/+IOW6BUDz2cS
CeM97TfECqZEcQnq9CYCuISRc7miijIjrgXamyxgsQFbo23ygEhx3fnWOeun6XzE
eJw1MikCyVXxadxJVtDClpk8l761JPgVsk5zgaE9F8a/Ht/eF4kA5+y2Dd66zNsX
wTEGicW5POWgz3PS2O+ry16LgJvE+dpfi3KEcqxU8Sc8NlLzpQaMQ46zgKF6r60v
9TBDE8wQ3wO6yFPQ/fbDZOra9wLHIaCKJm1KW2fz/XauG0YoU2VZNbre8dQahn+h
s9wo+uQuZVdnVrF2dqh1zfcVGEVZ1uIMFHKB6wcRzqXlOPH0MaucLBZ43q2PC7Ey
p+jRpnJHVGvv0Z4SrlgLQR4Oa1ckxOcUp4nTvxE4B23Ixjd1vQH8YZiYwVZZ7i7C
U/6kBDBav+7KOyG3EDxzbtSY1Xj4vbW20zgUQQa1+EOC5Zp9+G692Bz4XZgrlsje
6YyuoTqOdS40tZ5DZ0Wmq9xFRJ4LRn56iXKRT4ukmFjMpEqva7zWSy7UgwHNDe3i
ujgpasAeM3PeN8e8iiqNCO0lEkQR8Z/P6Dq9r9pM4VVYA9Auj5VPD6lpBZaKVyxd
PG5N3OUlFH5UFHztZCnUYzCHYhCjD9AMwwq9PqVpyijmmG1WrzYOOMg3TVG2rYkS
qSFLQtcSOjrC3dw0VIU++clJYMbUZHn9np5smOsCNHbPVRq1tG/sStUx0RCBiMQ2
Zy6ciUHKZCS027o0HGlTNtioBgAwr9JLZnX0a3KsnBM9IWACL5RVBIbmOr0ce6ku
H8BOfiDrr1HWAi8a6hGQcQUGWrXEeNoUEk1/PZMxvIm61q977bUB/Q4HzCdG4drj
VgiXoFuRNGAQLe/L3IxBIFLSDQKdI0gtTBBzml9w8kXDE6iA0Cp0PoHPGj+FLdgT
RQe2zDxyG5ZL0OBpRfegDax6Bjem119s41tT5pqGK/JIMEtgO3btGihowm8jlHz5
4DapywvxKEjad1f0A8aImi6BxBH1CiTbaetbsK1ScFU6mmTW/WRIwZwtOb+9HeJp
/PVkuA6p6NPYZT5/v8nEaxL6PbugisZGOFo5L0vXCwUjnC6rPXdcs387niMQPGIT
8VfXUtS9T3d06ZqSbEO/ELqGNv7lRoyT2JD6f2Ev2FVYTInqIZW4G37UU/DnV0Nb
v4AYHJEimq1RzbDm3QlVtd+Vv1yZ/3yVWqY0Cd1qMGUFdXezbr4y0Ie48c45o7T8
I3Pr6bOjUdEsPF0cnG5AM78MraQLXMBpUwHjS2VARUsliiM45sUivIx805oPFCjP
bX0pNhcyNypYhmNRolmj6yE/3bNZKyVsq3Mr0x0mtB98Bb9OLRjTeh3plaRvgxeu
lPk8GvdBdK2tGHltBzHFvr33Bt5w9kWWrkaT2+7H63Yh50KjKCxIOXbX7qCZ8ZGk
OTtOXkOn7tSmFTtuyM1MTQ5GdT2pAL51DdMaURMRU//WMOrqbzJUpsbKe2bA1GAK
WSZZZfBiI9w+F+CQkQK5gRLGdlqaLnPRsPvmiQxHoBUfcWqmnBKV33MiQ+4pZEOZ
P8qqxV9tcxkk378V0pM60hv5aRDegMlvs/QoAm/xsxhdSsuPBf/Dcwj23iyJoeTw
NzbiwvYXT++MvrJxNzYSXcEIPecleNA/7jyxRJZ+awt9SfFvoTmNYLL6ZPA57lQM
mGEJolDYRtYBPyKJB75j9YlLAfCuFC3CMsW6h34QlOUeyj8vPzjtKqs+aN8cGD3G
dEQJhUSJj8NLIWJyW/pa3dHgcmd8F+gvkw8OHAfQAtwiLKmcIEaP8pMnMRvtY0R7
lGRLqUfc6Bs5z18ecQjwxe3m8rM48Z3samcXoUfXO4IeI3JFbi7zBixPeH9kYoGF
wzmGHMci/1jf1XzlDw7LO+o1E3X8nymY0UYz0BTtB3y5J16eafq6H5gQDmm05rrb
H6aV48Lf7/Qa8S45VRbjqHjBPF08c1yr1jjcbN4d6skKObMOVgUENI+d65uN73hA
U04OZq9GGmMyzD11cOf/uqcsZTqBk1bLUb2UxpKDSVfHZXNCRuDPGKUNwC2rcL6r
wKlhd0u2864Ei1etNSSi9sGa5pDkm40444W7VLdcvaCjgXbiFeTFkdn323Za/ayU
+RDMCZxMueRLYiXmcJ/Ix58j0PkPbMz+BAd0lWdhDyKkZSQUyAnrI5MZw2yoTqc3
Ds8yOXyb5OpwwM4cy0qtTdLiriiKcmf1fP/J0GCeWoNjuOYeIVnCbmYxbZZLriQ0
4BYDRHW0kQVTiGZNVWkWrgX/xEAwecNNOs8PL6WaRfQuFGNiT6zqZ3gCqHM2zjU7
4blrB7iR0oobA0qQroSI4V5CF/PWVHIgyXSAFn+zL3zNM+U7nMOHGEYbFstKWjW/
aUrIUvitKw/bW2KbRAC9wP+N88UhUqQ2K7ZQtDSAcKVNjhMFG93bpwbZsYK7UMeU
t/IBnj3Pgr+TnF1daq1QUBCs/VjMHCAqUkKNMmkAzg2+Fhxn38v062RJlvsy74LI
BO/To1zzdaxON3/0QLwN1r8dKDMATv2htXO41C1RBXIBdqzdvku2psldoycmYHmU
dGjh10wXgGGIT1fPXyEvW99poIc95wGUMML64Oe2S2mrhW39gsCxZJgjuO+OZrof
kegfHmEx4t6mejbo5VPmPuUyrLoO8CudUCWDRQfD/1QvpTsNgFX/65p9PSLGLnDM
FZCi0Dp2AjNeUK17FUxecLTJ3ozO3tDh1SsE7c1QSiz3T2r0kaGbGcADtwIkz3FE
2BFVmWx35SIId3zc4IEIfFv37uZyu8UxVgKPM/tN+fAQ8A31DmX4XcU3BaZOvACT
+OQnJL25k303UKd9vQtqyd1Z1goZwEetKjpOduMsW3UuDBoFKzFepDeM7fRkcWB8
96ykDfcCkPHOV0iF2Gi0mX5bc6F6Go/ZY8nLDlZ0q7duDsEDj8NAFcK91PC+ujZ0
b9G7wgyf4bbQdRal3WWS30eGCWHPKbII6GklKfpIUK2ldG8B7hyBRbqB3918iNi6
WLMDUi/GAI0uEvxDSudav8JarS7+wiVanIWiE9j+9anYWAuSjVCXt+WP0LWHAxOv
ySI0NfIYeb5ir11sgGntXHtDJd5hNHWi4M9+SAaCKxcmXYIbtrMIBQyUo5WQe4rV
5Ew+jcwEjRbaZJp4SEUT6ulMKJSOWQ+D56xYNbBC6dH/BloOBaK8lbVgnIt4z+64
LPzeAQT7E4Z0X6qhCYzmCd4JAU8x8T9Q6fn90dH7O3diUrSskLOSNgMLj/djQUZf
SLpQ3duAGFzdh8wOLjKTEbwDplJ7L+xN+o73hFdEM1KGxH62LFTVf9n3kXE6KLLj
`protect END_PROTECTED
