`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2/v+3Yp8WV5vFbdYAZxUNiUgd8NjIWKou0uaal2/NtdPQDUw0u+gHu9WcoXyMFT5
/sTzUq1bvfUSR1uWmIxz6gTxZVEMMZIAVJ998Q1/9RPWJViPR5IdyjjfVyMhuj8T
VZCZXhKFipN4o5SWYL8k5OS6HaTnQXQYLdsepFEJQOKZtwtTABgn8c/Msb7JgUzn
jCf7UbcA8GC2p/Nb6iiRwPXOrsPDcaYhtdwZQ07ddliUyGO/LwRU1SN/TwatFpb3
ZAGN828xF+ELsuDBmJ1UESxFY5PNoDoX2cX8eb8D8lfOlPAQjbAUokKH6NDBLTG5
JLK+93ctHFyFlcXZhyh1ssDBVsYHjDorfr5TVlB2I24AnUswMYMpViyHMtl6Sf0h
Gf41mTRenEkLvRPti3rNyd7MJUKFkAA+RkyZo2ilqzpmp+PPMGd22RaT1jpSjF38
J7Eeq8Yj261tpEeOmyiLuzArkEqukO1X6Ern5g8Jbs4Tv/RybU7tqHKRvT8rGUKj
hryPO9tEOjGGzXrX9W24HiJCwnFsqMf0YdMVUCOzYcTgAVNXUEBnWDHo6ecld3J7
xJJ2DLie5vXSQ1c2JJmOe70ydd1CryvwNaJ/LGR2eFK8MxkmoAAqIHdiIb+eE2jK
e+iL6qh6JwWV1J7pzWbdnxQV02gRL/j0YMDFjEOD4i9x1e5X7wcGCQ+Utu8I/dfg
BqAQFV8HwvYRjrqnfNaGAA9WpUYYrlcDeOwZPYWGxsy6Vdfu37k1IBaM8iSY/FmU
mo3hjWcyL/ITqIm4P3O48dpvactxCBY+DqFyNC5DTt88R/EDstgMHpKWlqiIYWIJ
k3hQbxrU0bivAG8YGkR4fWv/kguMr4mS5OcMveHfy2IZ6m9O4erPZo+M2InIZ8kJ
WwTJvulH/eKPGYtpYmOwovCqyjmPjOJo5GLC4CIcD3/BFYuZsv5UfrhzF4GFCIZQ
KGl12YVAWhTZSrYb/p8dXmV0EUiDx8U1by7jnzVsTSu0ScpLO6pPT4Ta9EkaZcis
UIuNwZt2hNwU8c8ByGlTAYzJJEdzRpB4yYcDPHPcaNmaFmyvq8O6IpC/wnpIh8Bl
FhtD31Rt4SXAvuWaOLQu/ZsLzzne18oCdNhqZDnUmffJkLrllYd2U3oTJvVtDvQs
Fo3WakRcQ3Sm5XqFAHyIu3Lj5cFde8IZ2lWhpIE9cK+k5Ih7bF4dylGokP7vstKj
2NAw5O+EMbxWROid8ygfzayyTcYDK3c+80JN0NJKClrkruwA6Q2wSqsZN1ddKrMg
DA28ZZAp7TnKWMAix0q1SqhJzfB+LH3BoEgY32nrsz49C3/A+H/Rcw9h9GdtHil8
k15AwklkJMZ2Tu0LlDDDRXJpBTchlcb0Q83xsoUE7RlfsGuNhca4Mx5mUdXLwgDJ
DeR68yxPtbskYtLwpUiDrGrDaLM9w2NImzyZoPMPUmmr0fchDrtqlzJv8Q0WggNG
es0j/42kCIfhLEG38mxeOzF8LEA9NpwiBDQqNKCmZqYDrpT5U5S3mR0iQMIJVj1G
gvBLpqjgxtnEOt+Tgkn60bzyokebKFo1+RRF8ZoFXMhr+n5t2JZ5NPIuPjJTfoiG
w7AZx2sLllvPYIWb5jd//g==
`protect END_PROTECTED
