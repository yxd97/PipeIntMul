`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHNwLUo4W0U/Q07YPqgwz3eBhRjyLOhVlP6Uw9lCfamsKTkNkMaDaIZOwyWgQ1RH
ov4oxfmwIHuI9OcTQZ4A885NY2roRFHAAmRFUh+zfKmqD4QnQ3DkJdCTf3guljy1
TLrLIDzpRoLel4Cr35BVCpsIHfnRIcCJ4XX4T4BcMKAUvhoz2ugkNwJc/hCeYpuO
rVEt/Qft/pnFbTFCY6392mKggHVOkvVlUR650fjVAqvqspErLGaeOLC0vkVp5F/N
RX3FdDT4jztncsDFS7hU97tLeC4qUAtIeoUl5z1GrIUKN++o6u4oMLaNDN/+4E2G
seu9JdV7ePpeNDieZXfekmWiov1CUDdqloULV2cHb7EbBv2GHwGMMOtQJiLSHUaX
43a6VsTkeWP/GhptSOszn+baA/QDEBzDkwf1gdzm5QSMvTX1B/qtpcXLD7vxJngk
Qm9w2ppmBhh/rodOBKKPmJxsV7UvSEsJl03UT/njo5jhcwXiPvXlPycmAjXXVgRl
X7NPbWk28uzwPgQ+nlgpvnAeaxw7AesBJXwaQ4d8XWuzJJHprzao4kn/iy9Y2mON
xqPSbd+vLsO29JMLoGFdGL9iwdu8VaoGt1r4JIeAsq986hQ06/u63P6/I6kzJt58
jH9mWSEWEJJLWPE2AgaFAA==
`protect END_PROTECTED
