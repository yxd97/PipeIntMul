`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0v3Bhowev6Pn6J7q+4SaLgR9mYicAVCECwMYq/ByARv0jRLUz+cybBX2sprMylxp
M8ucKx0ZLGW025NskoQimb0ArrDReCZ+17Tvngztf8OrreBch8+cA/zvg3VjvAmJ
ArJ/EP6XTKARzdP4aBI1p1thdsIsx+sz00nv4TrOAXZCQmZ16/HaSQesjTqnLl/q
Ki1jJlC2p2AWXfJzEtB/F3mqa0wAyTXr0/LjhGKtB9gnEC86o6VVFhcYCFtL/zBE
NA1gb3Hsl9r/uFBS6nNXyuOexa8QYcSYor2OP5sbbbNAqFXjrQ2BejcqOHelH/4A
kjeOtxGm9LfZl7O1Y+i1/orcBnwQBG5ZcJl2aSUxSxbm2OULJMmAexeS/LHDjGq5
DTpTtMMU+32KRXPvsz/KBFk9+0/370FRRVa33KpS0Izs2OGNJE0QoT9FAOp2UAGW
lkvfxMRJ1vUcOxHegbmt9C0losVVgCXZtyjyjXoEqW8gi3y6qEDzfmuI3HPKr4ii
Ia6dPGzKN2gUOm/We1CxfvWJwPPm8UiaM5xJI6ZRnzpiJPY0utTQjUzQhEyEYedq
60fmqn49JrPnClAvoaJrwTLQP4dUQW6dmVKhv/IJLLwlixINAzhmKfs+EoGL+wEC
epS1TBKM+7QGDRf4InD4d9GuzZaHjawW8GoCmtDebc4dLzUT0NELzT1KbVB4AdTi
zi0DlNcJxbuuZ5tfGj+lKk8LsbvHx4a8B335CuABS8/9khLtQTgZlQfyuYZquYJD
xyOkSNdfbrkZE1GfVsaQz7vxOR97HAesGWrtxiZBFhEJzhYWfgXufQ+EKt0pSS4l
BqfRL8Gf7WQbNSlN2B9g0FSbCOulCiqWXzBzB0CE9Sy0ELGQvbsDD0tB9R053qzj
K6zM6zko0kmJLK7BmLWzz+pjvGxmQU2mL6Iglya/H6GFVhD5vEtS6RaYCW40AVTB
NKv9VanIeBOCJf0Y6lBAuXayy440PuArEmVii1XUFWAvP5YVumazpbPILYuiIi2P
giZL502qojqfJJRP5y4zb0mza/KmXrQk9Kf4as/kEmrg4SH9WBxKOukvhHITrezV
yxSGHjTBAz4rJNLVKNY24tesWFMA9TFvPky3Hzhz6fCjxDJWpv4zuLaqUg+6UCZf
T3o85GqeNyQtWfUXzb+RL6kIVLFb+hvKa5ioxFUSatk/aVBZFUykk9pZr7cdZ3FW
XSeo6jB0xPc6nUdUaTRAxg==
`protect END_PROTECTED
