`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bx6yJ9sUpgE1a1J7RIWSLCR9EIwSSKyZRH7XBx/wPfveOflwOXtcBclWzBuP43Tl
jgWKh7imfFSnRMx9SvD9Ud3y/DlLc80gS8quUXcN8mk4M3Ro7H+jUAquqJutes9y
U/df5jVkw7R78h6+l0bHLnsd/OYjfQ+baA7ngGSb/Nvubayq79IklCq1RKbTO9g5
Olokb3EY/HgKJqWZHI6SohdOKpdYqsDmdhAYRrkPMjpAWTokXJFHfPpWVbIpr+2/
01Sn8k1Zq/nQQN8aEbYs+an98aAYLd/S6A5oN96n7LrAGwz689VLptIh11qijRNf
gHgfVHB6ws1v1nynj4RVb7ZTVH2vCOA2RLtbr0VQRoJLxG5pp4287YEbdb3mzKpl
GZqoKJHYK8LYP6tDrg3eWJHfNVPyPj28hBhBYALldiHjgWLdjCLBqDqzh+fPUaUs
`protect END_PROTECTED
