`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zvu3bmVXuXttjb0KShtaXedHSnphXQ2zlo6P4sclHB5CS1S4i6qnoF7xFITaPMTK
C29wU1LDDrf1vr/OixQR490yWWea516shQmmUx0qqjlqAsRJsY6ExtDaTa7oQkN3
cl7rrdOtVwXRW/LkTA9l4d8cOYlyqndWUKDleka0Stn1WuP0Ud4XNKXO2KvjTvwl
jHcpLaTm9LD4uIwfOFtQk3v2VvY72NLpd3wNjl+rA/1XRXa56EPHHsGbUQSlZ4YZ
gnqZPO1xzsRExdet3zqisiuI0Mj/7SfINgFwKtgTHSFn/InZIf0qjdodRox3S2Ur
RN8esXSOGozNvV08uPOf4cA4R8oge1fdUAfj6groY2ONg1iXH4TmN9QFtktj25HO
WmSTQ4VJXWtpu+sxAjbcZuEdLEovQOMwWG1kF+1MHMDI8UtZYvDXxbeWJuo7mBir
a1hYJw6R7S1c08irSybP8TpK/l+0OdCqdp1WR/h/8N8=
`protect END_PROTECTED
