`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3QTtjxuuDQfnnv654dIj/wNQx6OLUOzBtOe4EOM5Zt+8R2YgYOarziT9jz4Wv4Fw
NhYg2etmnxiO7JyVYIiWwWrWEtzNyJfL3YEhN1dmgYlBGkyL7Y/g6tFC8QNJ0VMe
d3xp9yzYroVPPIo/ngEHjXj39Ew0Al02eRuxCYAnwGL8mrRSooYzvbY8ZAcakdmk
PW1rFHH38dqIye+C4YsaLWjlFKDxw9tM0BwIWsgkuVjRnbAMoLaTzzYSlRIA7AN+
/O8TBDFFLHEPqLsYq0Dv7b8C3xysu8UjcyBFkYby9u7FYoMwmILB339zjDs8IdTq
txgOhAuFpGCEddo69JeixqqMB0ZrFNTU9/u9vMtMB+8F9mmtPP9OUsYEeuBd1cEd
1gW2UfbWWtE5caO3UKHRwpdbQAURczUSj3KsMvXcLIf2fphX6bHtbzY42WZP1Kyc
YNfaxXOx+uKQN7L/LMcmdWZi10QkGsluK/5Y+e/1Wh0=
`protect END_PROTECTED
