`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAYPSfsDhdb4b75tYLcsk0wtR4BO33GlyaqvIP7/g4aFqMfc6rFINibkPZ58ckyN
hAY4et1qPJYP8i/Q761A2S9i34K2Zm/U9W9h8zAeHQJKZ0/PVr+EInhWpFfUIZDO
LlfzVGElJAmlTC9qXaPYB0SIKpYoOpFYJCjzjMLZQ4KwhI24ZcLAfmkidhbpAPPP
v5XCBHx1HataL4haefo43f76jqFArpzYdt90ctjbQOcWIs45+3OIcq2CQlD21tB9
5imrdWSw8DoE6XT+qA0jqnYmTO8e9rTwHlxVTAayR9CrLhGQ1HRbpqs2ww3cdm8j
FKWmqMl3f0JDn8ennzu/DFN/oHpl+dfhRKa5VWx6svzxrGElKosL7UrkMyUj8mIx
c3GBRhMtMFHztxmyu2BzFDPFfT6JvzxwcDCl0h4MIlWNPjSTxuhtUWWQFxtJugbd
eOHysrgTu8wwPSdQTSEmNhb8hDTHhKiTbRp/aUw4i36NrLogg5EMNtNnalHz6eqJ
MF2OyG9Ix3qwBsOZYF2IVA==
`protect END_PROTECTED
