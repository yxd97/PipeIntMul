`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2XdVQj59EoES7PAs6990peI4Y6804Jno+FdLNv3sx0jw35SpjLIyno31qBktSc4J
TmUUMYWRGE7QUBL5Mk7N4SJpWSVfxhEngPOKGoGR/lbVBJ3Hp3eLNJ1q5PAOKMik
YcmlPzwnYjuHeCHNh121K2ZXzzQwsrTmUuIeG9NFlz+bUba4gTfi2UdYeMmcbNv6
CrwB0E3odT4opzcQsGHpsTsfbOTAYiN7N4pGEO+TD3XfqQ7GBUVKAuRTijPBmGqx
gpxoY5yFbxijD5cYJPTb0vUXx3lWpposICjdXOKtWTQuYX4hM/I9h7mN9OUKlLU0
cKsIKqa+dB3cYBDsA3ICf0bqRocM1VTtyrHNPsZwec+6malC3H1yAeUTWAsAiAhe
nMJFloOOmLwqzslTYZFOuomZhREj5hFAltNo3fup91jDXxspbJ+ugEVzRxyI52pL
qYBv+sI7aNfw3EHS3ILCQHwR9C85EFtAJf9YWlhgNMb4Q2wa94gdqOBQ8RDWD3Ts
4drYAQOnhRxbspBbCW54o8svl5vf1IM2WcPL8Wkw3tgLbEd7UN42GzYa3QuKYb9n
YoDkElI+tm8ITQDMlWl57zsM3L7GBn2J60kA86ie8iBJohzFy95M57xR3y8Dyjie
HgprRKR8U4O9ZrZn+8H+1mDH0ITe4zhn8JXEh6f/jQOxg7TMo057f2oKxA2qeY4q
8Bp06A2arRtCdPMlmXeW0xCSGsKg7t32/D65Iyr7vIIs3Ru7zGU8JEDsqPuR2qvT
krKmD/lIAJI9H7zt4EllsNuO/q12DpKlSeEmYCniRQv/Ecsrx1is4ssaZm2Dip1B
Oc7Cb2cReCj+CeomepIdxxORsaUJu2fAnhjJUEzZo8CJPYDuygPLHe6k56xs95me
yC7k1rvC9ajDINW9da2MzxMAmxCQeWMWnA7OlDfCJPMDJzNg+w3zorN5oDTZSeqc
cSmDHVY0D13a8NvG3XwI0oaxC0L1cthQqQIkZb5nUtdIRcBlsZV2WC79Rl8BYWy/
`protect END_PROTECTED
