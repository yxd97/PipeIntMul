`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+Tp/a6sw3z/sJTF2ODgXeoj9XZZVNYo9Vrw+Bd6B1UMvgcama/KdH35ZdcpXmVc
du5q0JbWIpq4yk+6QsG7gReVXbyX1pJG1DwY1VocsnSy7FjysZ7yFScJ0ktpoojz
xVoSrW5/PZ6nRrMvHK0ssWBy3C8SZecD8r6j21irwauwRDGZVI/o+NPNlHsHpISL
6/gnZmF+Oh2f93ZUb+AFEjDsAEtA1b5sXPekae2mdOWMUrMWvAyFiBUuatnsMRKb
QgUKucfgDBemezTwNxZmo+cKTcVZ7g5ALhV4h/tIeevQRlzLrwc1NHQr6Dh4MNy+
mthVXbvJRyAiuBvTqVgptFViFiznp4XrnptOOJeqLnG/hU2xEwj0ojx+GVd2lvAz
RKwlKlEOgufoEkTmLmSRf7CvWhLX5s+xaO7hhlYuoSoLrziDd8arr+/YAv2HYCL3
BH3V/x1kVBXVJLojMrMbXj++WPdltUbavfWk+hd/RyVgawXlMDn1qWloVm2Cb3oU
D0abcIVvXto3SQKoGzWRnR5SbsLBLQu7cj7gdefkM8vEgh+wrwEbjwGomaClCUyY
JtgnP8iQa5BkZ6nLeAU9IZQe/N9bHvtlG+PB/7248Et5eEhjhEzoCGm+Wc3hnquG
uHUY1F4NWppXmfsJW71eB3Z8ouvrd0xgldysQH02BOcRAYn3AFa7jcV7PFIPcmsK
tFh8jRv19dEP4L4yEfIRFWoSFvFyTMEFAYv8FwCgDa/fjDvjCAxwT/CgF6bsJtzY
AXjyx+2dScKNovHU7CbeLN56LdrQLXpXqnERneCEvBZtWiHjMCnydN6Gw+1waEdI
yqujQJFzyqkNY06czDQdsYNxoWTPR0YmQOSKoqIswbuRAhFVVfG2Usg9PEquxVjg
zxusZ6IuLOh1cU39OikELQJzi73MOiLNAUjKv/EDvvkNN3oImICv27riW/t1iBz/
sTjaZAVk1hinrr72KMBTsJK7NGVEB1Q10epF+Eny9fHKgqfTW7xOPtF09JLFAn3o
VFbeCV+aWbTkSrYzUDqd/5Jz+9yuqXct73Ls7DvBJu1cUaOYN4KQBcOzpqQDZoN2
UktvUWd3YfcyK7SfHtqz99Ol0OKwli0Ok9RHZJ5U7i+YBxWb70mY+CiR63DTnO/m
C6PTHm57O+PAUFuXAF+eBvWybBTkXm6buMSVexeFdP89Fd9492YtpukRHGN2kior
ZkYoZu++DNT/+MGJ1QtEth+/XhbZEbCqb0OF7+E2ZZ9X1eCXFs1HM8DE0D7d0RXP
rVET8pbWG0AETf1gFI+Za0qA5cKU39N3+v/AtsGjNQh10W5fylc2u6f3wFre8YS2
wqLVdlR/bl3zA7dfxiXgFw==
`protect END_PROTECTED
