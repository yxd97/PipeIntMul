`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7ScnoRXf1BqVdl1T5MYBjeX1PnMq8mLjyJMSqQl8z41itCorzfieYOFRoFqbIE1
SajYMNMUV40ev8OLt9LwVcWLUkLMSeKLqY7KoFWHZQVmhNpLriCHUnspHB/UuUuJ
FsqSwcFHJcbZVgXwf3UD+EyLV88GtZcHu7XnvxVF6HbJcM7hT+1v2diUwdLtProS
uyd6rVn1+Dyv5+yHIxHz+w9uswDRK4xE4LkcT9ktxUmuvYnOzXS2h82yRCJrlIQE
slJpLYU0YM5jriUqTY7KcEEduxkOwXhRpnQC71oLr1RdOVKqXHiz9+ghFqFusFit
PTwGXJchVa0BJmiQz0olwYxg66/QoA9tBVzW3DsOtaY=
`protect END_PROTECTED
