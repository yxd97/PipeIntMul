`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lkqaXsWV4Zbr5Qg9QV3Kmuwz4DLI6YcATFUi/I50Wz8JZiPN4SgaEhLZeTk8aBC3
H0rXBj+JTJ2CWzmis5QlfDwxoDAAP5hUfs2IvqjCcN6h1MFF1/e4/HkZJGlxPQ5F
zmgaMD90dpEYehbvqmK74LZqHkp0LNoFnHSMcIum8oJfN3AgMBLy2y7TilT5P4WW
8OR5jNOnS6vz3GD7TJeUzBlO0EElj+Oj6Rx0jNZRszq8Ejj22ECpGYyDhUocnHne
IJKBN3MRMYtGiLoq+2NOqi07GQAvvH7A7fMMUGpU0/+GEf7h/ajnsjPrq8xk/W2E
52uXC+fkQu3ahETpp2jCe1MtWI/0hNOkdhxFEpIx0e6OdZce3OqdDcBrxWk7p54D
OKOgW9DCtY+aw4JeaiTAGRwmPvICyQ8GDPiUopzXXfktJohcnjj/5yDBBrAFKfIS
BVqejV6D80PDUxFHPb2RPQiO3k0E6yt5LGz0ILmKytT+A+PqzMQN+RVlfqm4TW3J
S9TAq0II3YUPvqOYS4v8/umL4mJyohrAy3lIttPNUQd0x+0cNB9VV88hVF5cEBgc
YQddPrq7JBX86aJIRjG1oWdKa/t0TCsvUUuhWk8m8KooDdbWGj+IAJZhsthTBYFi
hNamko23BvZpO5i/22Sxd+/rNTo+4aYJQ1R/r86GQOIIZ1zbZhr1D7HCgQ60tMQ4
iCymQPRqdGBa4CpNNsX7lvAl2wivhvjAHLpj5hun9bHSCCpLodhu/p+yxrQMax0N
v9Gs9ER0xwmKihNLm0aJx0TJYkvwuGWa8GeJA4KIisXWPxz4dqM7TwOY0M2qEYiv
HDMisIT6sMSUPIUR7a3dV5CgpDfsxSg8rjzu2vhfDYESXhf1n3KePPR5NSoA+k/r
s6Za6o2m0KtpzfjNjPkbglZT5Wj+ijIqj5oVflD66HhyoGn8F+ioVACfILgVPvsT
M/xBK7AXg64qvGwrqWu8Bq2dK+SP7qlLtPvDHmQSpt5nW+3aVk3Ry3KSshm5p7st
2GqV7B9p/MxE8oPpJD2jYOhywd5mnroCYVAZd94foLjGMIrtHgcaLamG0ZNYCVm7
qwlBo7F4kK93LxI4npB+maAZjKHWwQTs1LE4n5qv1agjrzEhkmMBXQpfr0iHbJ2X
VuvzpxWcOE1giECWv578FrB9FkgoZKM4Bx8ULaLDgmABlg45lDCE94SktubuYeBZ
E/z/yvUQZYSE9pkfLkEKNWsyshk1ae6IM3CcLX8GsDc=
`protect END_PROTECTED
