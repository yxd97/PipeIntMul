`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q/AK7IwDRt4fEPxczIzshSwP02hNoAjpY/BhrJ61ubnV1CVElJH7Q+NFtCRMX2lV
Aihv3JupwNHJO7bYyxPwNLzc9ebhAUwUeDtkw2A1+eiwvRA1A1iqWPA39XVkGOrD
0mil3UCRgQc43sY65nIzOLoCvx2xPc+ra+ohIVY22NOU0+xuL4GST1yhVN3WEmnM
ggFni40Dh/0AaTIv+GokpvwwPURjmAq6rwFyOERnpDYKnA/HV1p+IFSkZwcMJXvi
Q61CwiRYhWoXl+msltBASUzG4MOau6soe+qXfwmBtLgU7yIFm1dONCbRTpKVI0mq
MEeFRLHBahmxlAZF4kqP6XHNjxN85/486UMdElFk7s4LjUt6sTY4ZjivdcnF6HgA
1ZXnf/x13T3HAOSiHXAgirEjv/qWmINAbso3+3qUJkjs2mU2LNwrWBwm0zwQxmZ7
Sy4V1A5ay7QVcCfH5qxkHrHgvV2v0/T9m0pZu8Rc/+q9uceDEAIUyCfn/+NlYeCo
O37tWM4mpz3lZfqV9FrQTT8Ohh1v/OS+vlH0sugaV/dNIeeMFeDdyhpplezb45Xz
LrRFq4ZVHfuN+Yk8/k/DzpXTKhgGyCsMlVHM54ngGqGirFjwLQ6sEG4gX9EBJtv7
MXnBE4CYVEtrhAvFZMgUGv+HBGxNzW8TRedOkWXVxF+G09FCOng+fzcBBWwAk0OH
fQYHGIM/g880F+6ZdF5lqcpDofSxhhC/SKWJx0hMIoIKdyIGMe1zTEwnORXd9g/N
U88H1H6fwt9XKYqSEs5NCLdrb3bHNkM1sxFQ5CjFTd6dh8rZQSLr+tkr/F8vsAKr
pFS+MLThOhNhPnmx7m9X6SR0hKi6JcbcD7G4C6GVKnoY3zCYQ+I1iHR0QpWqeTXX
pVeKBFmZ4utJdZr5vGSnucIM2iRyUWTD0WK3SsLrSMkQkasj7zEbwdffQnhgcmY6
xPO0xNjswV+WxFyrkzcwPe7ImV/ElzMDRcC4vbgORts=
`protect END_PROTECTED
