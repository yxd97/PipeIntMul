`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wYnINYJeYBbGAB5a8UUemj0MGdk0H0SbR9MONnf8QW+Gfi6OPtRuynBluc+i3GXK
MFdC9ABTRscRCEXtU0VXFYZrbHEVaMTpLEZ+cLf+pK7+z9QOzhfxNXrKaGJq/KNc
QBvBIhcDleJvM90ElJQUaLRdKD2xMiGcd0b9SyBga4+Z72Q8CCY5pN0FS7UvDitv
kXqjbA76nvDqnc84IJ/nlrl2UO5yeBl3nAVTFAgAc2WjE2V7dsJO/BjWf3mz9HMc
Xw1J9QxnSt2SmyhZkcW8mykSaKq+HrzpFtbpsiASdrcRMJRKUhie9qZD2jtLbIcj
15yaokPwozva0qjeUMgSyzO8RmW+SWirQZlA/fH+s+aySnfhMUulk/VjTD/6lnCt
ebojOXwLb0760VxuI5GK0gazA/n7+aDE835VakJOyiirqUK8CypwkjdVWmSZqyPs
qnAIAgilSs1Bf/o8xRyT/iVWlT2nCcF94tnGYoh6nWwFMijGeVF/Vnsqbl+h2mKQ
nWFhGBTzPJf2V8P46SmnIPAY41+rhhtLZFZ3oQaBdqpr1FitOFLKGeeuy98BcNOR
MPIu1NGzpZEY6kHr6Egkz50VKgDnqmfceINQ7MxI4bprtpzsQlSWLi0F+ci3Qaz4
0wRHzGris/VTbK1F23G9lC04HbOxhM/xIfDBT5oOOgjKs8ls8SwBptoyOhKVU//9
ke2Ua98H6x1shbqg9t/VJhrFKOOQtAcl83zzpcx72lC4hRwgd9I7UfJw+OvE2aDP
lyTFRyBMOM2WVpH9q2zIDWGd5XDrNU4uHqvQb9vXx16/oCQAI5G7fWtoVFruE4Wo
rNN7AOtpMkWuaA2bcqG3ywxv70jpB8NFLtWyy/1+F/zdfAwySN8Aym2vevH3c4Lo
520VRFFFaJaTj86DNBh8IdcuEJp40kM3iRWCyKkYHnXwBms5DUuBDmkEsv6HYXU0
T1OK9ykSXDcRKcuhOJrsCMRyPfeFhrr1LYieatEf9hounfNTgjEZaybt0FGS5cyh
boeYILR3wgBjFhEuRVo0O1Fno/wHLa4VNyhfhrtE0K0YbAe3KGsJzE6rUJ5pkf81
iK3PbUnrrgmVeNi0o36Y067rm16itclPKh1qdLPZsDfL+800UOGUZOGZyRgcDATi
roodmdtEv6nMy/tZjthw9Pi8HsUzlMttJbZdzyK7nhF0L5YalNrswc7A1nV+hasP
ZaNb6hX90cyOa+zP/CrTeAmXx1DhQFYVv5r4zuush4pOS3zysSh5RfoJCOFHXNXt
uqe+i1XBVJWio3vCr/iCCdazP6W7i5M0MRRiTHCbl5W5wdxOKLIBu+PbJOntBdw+
PYywH+hUaBzbqMGMmZNu5xhdxNUFWX5ONZzAAuRyMeyAgk58blrkF4xdouf3PxYK
2IK85fxvxp+VY2HqTpp1ZIhjgWYgzZpPxswhHxB59x1iY4BWESDS5p2HKaxL3ooS
BdTeVApP2Z+77Nya/RsmrjefWa6V45Qyga7RmC3gneYmz5tw000VuBk0FDK7RuBB
/SAUz/sIPb6liZ3CQ2teDXEnW7J+3EcAJq+g4iFtt2Kty+irLPyQNzCbZZPRhsgh
Wr0ABv2w48+QxkGbBMTdOaCtfRhbBl0FFkZ5YfkwB+D+4pBrDOudoGFliyQ8/Klz
vxkJH4OWPj6l0q9qMscwPFNEvSOquY13TmzaqSXdKQPjvrboOWWyINU0tzrnZYeV
dnKiRuWfDfvKfBZZ1pe58JeHX9mxgER6SpRBMFrCO7p8N3IipwziAn2VGSUEfhFk
AuWw33iTaJNkd/0HDL8NdRku+qmlRkZ3JRXKpmvcXvaFSgvktodygBShHfAsqHuQ
ctjbj8sfRT07q3dpjfJowVNh8n0/fEzR44cW4yJtJQmxuhLuQ8BsqDEeQLs4oxW/
/e9IaT715gTmBoH8FtwYpNioS8DjDUN86QDIvtKI7IR7giWfneCiIzs2Btm4RM/r
dCe4gdvhHvKwvqPGvxk5JmOCkcLmH7NmmVKhfyqGqHjvg0XQb8eVF7MSEXKKRqIo
tN3zUFzNmS+0Y835tkW975qmb7TbKryKTKZNopZd0kO4HR5qfc0Is+AOCxEpZGnC
cLF3AnRrasvZd/LxlUQMUqGHZowSOWKIM41/3M5SVhG2oR7Rml6CjDYStPLq9NMV
EsqLR+JObgxOEk+i0KKBjXZ6WgNCriLSPGL0rf+PMVioKlImAkcjxjrd2K/nJ3mk
EHArSR1U2hknxqWO0HZMLOASx9nUgmEnsAisL+8cWwrgWFUJ3rwXsbmkbekmAx74
zLJIaHAImyCbvWUNnbA5I/z+Zvj54/+ccLbrQz7Ve6GqGeANm2Eu1XiC+ptmmQpC
iUksX7acvRp+yqN3NxVyJI+gs6PBSU0iOZE3nmi2TWN0PdNPwxeSZXYab5m+TE8A
M+//FFS7BerYCygN7+5B6Ym4mYuSvu9SPWjXDcS6GIahM+kKz7CxM7frniAmFpRU
PwrcyHGdK7U+PUugG/O4xIxqUzVo9ikiela9kjQyGca8GgOoM+WFVoPCphys08BA
+P3xHeYv4gfqj1maX9N4QDmhz63gyV9V/TSqL7bpcuQxwbkUWhsJG8w2+GLCZpAK
g5Sd/Rrar9j4rvqsXU8LVukwPPnUgkKSEramz6uq7pr3IEKkI/aiY6HSgDS9GUDm
9wC4QGANfXugDUKTcsxTNUr4XFF0A5rolZc3ocmwtGMPXC62PKy43Crinn+XkApj
GLVnFxfs4+Dfa3iykM6F3iBRzHuz4dUZPIJbUA9t3/rwxeW4V9KvlLmqKJVbrLPV
H2Zk/qg8zQviM3uil18CYhaq4zbeHDtjmX2S+RW9JO7K/thfDkHLXo4KGE3b0X9Z
7NwpReHgBApGFEHcwCMIYF54BwtQQx2MT5Ov8TDFzUYNixXaFvLt6ByBt+/V1Q12
XrX6VzXV2lv8Na4qkltcSPDv52H8FeQ4FcCgZ0DUTXL2QBnC++3Y7ShytlWzMES/
trYAJn7Am3k9IfZ9EynGvc8XN2kuiDo9HjMVbBoX5g/CTALhRspceXB2qY6ZihD/
HLY66mriaxcyNGIfeLrh7E5zJLrA1RcRa0g7Oy0F5qdKgo2ceRweH2xxfn4mQj8E
dRTpGPmDGdfboXKzkCjq92LsYpi52vaiwcRunu9ybOL/+JudzjStFOX61svOxjUR
eKksNuU9LKmqXRKYxpcadqSVZXsGYmnqpT7LVTUEcxqNHeyFNg7SAAijF+XvbfC9
xq6Nip2n0qktM3raxZWWCw5++AlfhijCh0SpR2kxV3WMsrDVtGCt29Og9QH88v12
JglhMOp7pbLP/Wi6KYy42JSR2QOLQorWkN0eJv440xTltGPurMOpPip6U9CR25tR
02WLLrAyWOHFb4dQ6cwAcBW4d9Nw1Ot+M/7Atyc3wFfRdfssSQaiF/q3DFWrlnPT
ZgXT3y2VkLuUjgiCXJ+L4dZu1JNNBG5MIVNg8xZRdFBO2vcD4p4hVi7IjdE9NoxL
pYRND07EiLy9Yw2Waz6c6CYuAVbaHB+Pa/wvssmPCd/O3Otrlkt/aix+0JQ82Su4
ebcuJ2lCit+eEkke3mXJqNlyPamOkD3mWwWfj8g4LhE1ibKzyHuDU+xhyGvp5UOk
onH9qSPJaXg4fXFgWLv8BOOq8BfwSihHdi7G/om5fPqE5ZAV6PIyC5W/AsrktPCA
YM6YWb231lKf0PxlL+JJWQ/xeHr9E6EdSEEHjZ1IAknLwwW3a0iUX27qklj2ikkt
pHF4KDe6WjQTra0gAuQH0TGYzgesw8sTBjA1VOIXGvVcnw5ZhTu9AYDDGHfvRk1L
gr+8SK01PpN2tb2JrcBeNxvLQGxiAytfjv8k1NvGsMVNcAcAGDBiNOa2NUevx5Dr
kkPjgJrx/q1hQZeMPjIRz+vqRw4aA60XQi3aKTvetTWgpPw884CccnLjm/GD9Sct
6vetio6HnupuINorkys1k++SuVUfCDAHkBg1D2KpLRBNWUbJDtYJXqYvT9hrWbEG
87RD9aVO+30Rd068Vq/bE1TzUpDPRUjNd/devwS6DYp5Uq0WB22ZE6X+aFi/yqbv
YW/Ct/cgN0Sm7DGhmitv0h5n+NluMaThTeGEV2pI2bQ4K5cFSw+aimK7izB6YZb6
OEm704Bl0TOfOQzzDOYKpx7aL1pnkfE+oi/yTxEaAvv9NBpAtCCR6UtBhP1eW0O2
0K5EwH+50UKMTjqHUW8d+vW6MC2fpJiggsTq//T+lfZmmS85hTdFGC8rjqt97c/G
5B7D8U4isewNRXmE0CPKOa9K6YmqRizwO6Om2vocJJHHmRd9BwJYWFJD0G/JXhnw
UAHPLQJlESDpO4Fd/HG/JIs/LttQY8ZF9z4vvMUcvUve2Tm85JJok8U4aBQJkHaI
1ktNv87iVpJ/JvUgs7IMsNl4ugNQgmoPbRhQmYO8a7cmPC2GxVTiqtxjMQ1D9tI5
CyUtqHPYiHgqGK1dJVbBe6w47fzo7WhVC93cBk7ROX6kmeylY0WocIA8aP7DZW6k
SYxQ9jUPWz61tfMVXJt8PxMi0iayWqOvS3mvwMxxlno4kg2jdR4OHnOsOfTePoA8
0N5K1e5tDJRSfuhPaGdVcvmrF08aJtPU5XCo+kmSECKtJ8XHx+vrsMLE3a1wNH0W
h2L/oVCiimQo4unqWydmQ8g8WDIaMiFXn5rSX04v8jcRlWBmQWYmSsEFE39AxJP2
+WBkLjbFiuYCIW8C+eb12zysjfGoy2BeNuRJ3LX1N0lLl/NWb3Q2uUKxGEHnEAAG
EvBWVvQYgTTL6jvxewHY3golyEQ5E39UR+dCmrUv/VM2ywaDGLFvnTaz5118kRr9
TEXi6Cf0vGyiQMyplvcH7HH7RZCXOaV1+gnhCIkIT62RCCzhwCQrF7CdmiBO7K6/
tmjaMnjA3W9U8GhzUJ0hdONwryrW7DJsgzJeEFouk9HhsYQX7hxZCcmxG8ShjpnM
crBRgTCuIL5UXppW+dIDsu35SxvIJ2XMSrf4PldMYQO5m7vs7E78NNckFViVAEza
OMn9uDTMQCDol2XvYrdr6Ovvbk7rzSZ4rKwqug7R9reZ+DoBebIfRbgkxiKFVPe4
aEuNckLZ5r9iLIefxIw39JxSUmpgo8F0dtnQjjR62BTTWM1+1D9ohPGgZLQRELfZ
Ot3slHCmZuUNSsPX37FEXQ/2SsSvaQxr3GLNnz5QV1I/72ovExPwZQTjQcUI+lzl
yaIrccz28b2EGvdnH860X9QznPYPFhJ3Mx7iWvrR3dg6Qg2hQASRioQ/gMhWy+mH
tKFBnH3JPulK4ubg+97d6cmbfyWcW8SNYzCQXXkiLKq42vFVuOO7G0idU3nfoc67
ldCiiO0qmvfiLkXngoHtiGxN5gErBaJgxROmsB1DTraOxONRR5XzuIHLpEVYaLLl
4+jSNkXvaInWetp7kIxfTSL8j4YFqZLNuco/QZUicyZlbHXpXSZ5oC5M689s0hM9
kOOtKJGhznBJ+zj+qbpvGJxngj+m47H8kCxF+VfBDGMdKiraRN9cxKkNbrN+/+Q4
NUINMKjZR0odFjKop4SeIm0V+35ofJv4kPtl8FcA6ZlDncNC8fnuGX2/cGWt1Swa
JwkwQGKxIpY7djPdRJx2sNvHhc01yxd5b67vOgb910mwkIcuK2C9e+OOuL1XzX5Q
LEeX/vp4be+spZE/a6X5eFxig49kRlc576qTr/3AcLHhaJRuEnLRcuF/e+h5SbLz
mxqJW4lTfp5IRkkTdd6nzs0lA46vaNH29n1NHxqS11XBhaEN0quYK0pPIckd0f4Y
k4hLKsUYYccZc/uwWx+Zx4dMhuCcLEIGB4pGw5hMBQEqMHJgVzbfrQf32Agq/1Yl
OFqlkGZcqM4SqRQRSeHryAvKTStvTqgVMIqr+O12EfgRRZx95H7aQeXX5XdN82sa
eZjoJVEgwsxScPFoPXOAd6f1tezUp4Ht8iageI9IxIuf6Tdl8cmHHyYM+B3oKpO8
wpz0cvbFaNr/Hpb/VrvivDbpMuotJxJgbM6v1pSAarj48OUPcLTVZHjI+3Fk7ASs
wf5VYGtvfa9eCwTGUuaa0O/RPADUa5tCWyeAW1uJ7RBExbRzVHdO/kClRKpM56mI
3phk4PfB+uU+XS/YQ1/HbRy+7+r0GnNrrVfPkEmQYorSG1vMJx+t+EDNmRpzSSsW
MExovIXdJMULCiH7vmTodg+IRINIQ2meTt+3pOXrX1qNwNTO7vHjweWapaExQcS1
p2LFz7E9hKkmw5+eI5sRhYea5E31NOfZoIqqXvJjbt1nUq8x2pdmB4rMLDICFUpD
tzH16U400ucJqzd7TwRWC8F4tvIncpwDF9w7Sx9iS2iMIEqTnC5sKdio/bTYfdQ6
4XWCz9YYNJy4D92BfWMaNVjHCdHqBSSBYM9VAUEu7+MD19j/Q+MaEZ9aS9dbNpn4
56pBftgsliX7JZ5Oy9t2CVMNtmcVzAE9kDcOCxbESbuvly64jEo9Ht+C318rlVEw
bG1EOY3MX96+Svn6bzNdaSJBQPLomF4hCMw97C3WmkRolA/DOULaTwBkctwP4B4+
TBkKMn73t73FbcTiAGJ7YSHyB9Ukocj71mQ6mM/3A5RzWw8NAgv3TcKbn4jBgyEm
mvobaYwjDMnoS+LHaWLEfm5kPDhIlVrcgKhi3/6S8lbqKPjC2rvaBYsfPW22W8G+
iALPdfHbIjFpskXU16FhLudo8UafWr069qMAVsR+9tK0fjYI38r3CNQRhPbAgTem
x+8VpdoLuJbpTAAmKN12abZWDQya3vZ+spjeQF1IFeBhM9PScWhP9vfX3F9aO0xq
idt308ZVQDw0Hfi35rTA3yG0k9J3AxOEJwNjwbeqA/gQ2mAhtZTi6EyCQu6/32vk
CDAfnDQ7vP/r1MzNarXsGp96meuLbONNU9ThKnqLjUNsONos1bBJa8lUgDdQ9aMm
0mzMRFrQwcygub5bllDh0P7VIsFtkBThzMDj2r+eSTTY9T2NIg8Ok8fCzT2mlqbc
I3wh6htbAu4Nz2noLzUlWB+Zi23D1b34qwSOgiPRmMdJX6UpPCiBN7JI3XmkBhU6
4dhSHO7YqftdHaSHiZg/s9qcI6kCQ5Az4iHPrAEfUihfuJyryDTzDnsEeM2YxULU
NkoZG7nZCCxtwKuxRXzQZASfUhKjUgxfyEKaqNND1+0luAdH9LYTWaLJYXJTn7cV
8f0Q0Qx0BC+O6xhKC+qXSULC7l5ywtAG5qexlwuoEqpmnOeK4Zi81/xRxk4ccY7I
jri66TqJv5MG/p7V/2Drj8FgTEwQUCvNzjRh4HXOFV1aIV02tPQJNXt3chyG5WwP
INIR1XgP0Eg5UVSRpQUGEsN0EHXktnq5EzW01gheePiSgYDlgfMIBbSA9M6iwiYT
5JptM8sPa3zeXADFSBGba5qPQq8rtopbHru1U7xj/7aPEf6P1tg2mLkv9YafEE51
1mNLfYmI7hASpGoPBH2c4h/x3jtbyYOFIr+I67e5RADx9RXZxngcjikrkPm2kVcG
SxYTTYoT5wSWYDfTd5lSlM9hP7gsMpEHU6tIY78SRGRXOcOo2Itj+0EsQmoaYtv4
ISOd5PnS6XYXc4zOK3pYhDVPzWwqa/NDcwlhpqKT3AQVMSP01Ixu0BeIq/glH21I
MpQAPzp+WwpF4frOfkO1DbW2JZz4brC8fEkQt1zuffdhPS4SLXMUQD+uu7YFq//A
fUa+U83ZiDRyiXVxVCQKVDQip2GMr+23SFNiSwd+hGBk9oIgnPl3GtCL9VZNZzVi
fnBmzejuyBI/JlRIkw8gA1F3kxgoQ6lmF5joCjrLOh7H5K7vts6Df/8c5t+81f+9
wBTGWLlgaGWxhAOEujci6C2ZTCZRM+AO2EIEFJtf71puY+f5VQ58hmz9R2XU1Rnb
jb/A3eXfohdQJq1cY2e//ZLk0DdQgxs/x+PZudWeLt93ZbkPxPnq5C3sipMI6fBR
8+D3oP/0yasuSWBKzlMZVwXD9UTTeddme+JqSqHY9tvEuUu0OFZ5+NG6MS0iuIUp
GA4jvQ/KLCiWmKT2Q9kDkcIaGj6hwVzWWAE1+WZ0DH/a3Ra2o1Pp9YFUk2Kqacqo
Zubhst6VpXXigNGKRbzGnl2fIJNgQf0Up88806sLCorthPDpie7lNuSfTOTApzZT
IiBG3tZlPCIQX7CWRRIhc53mays10y95q2mIwMmSzPsmF1hOTB0+vr0PNELnAbdv
YPAgBTaF+cFACohQjQ+059l1g4rTFEixX1TRbzlsACfG0xnrxxqaviGNJ3bS6UcG
dHC1rQYc0+csE+UynpDR2jwcBEGF2lJY3xwMKgLoP325zjJJJeGQ/FRRQWfGyGbf
1Lc9SeCyp6o0vxzSatFav1ug+IsdluZCb6ivPbJ/vAB4DGrpHd+/j5AonynUQZeh
KWCoryDHRlqSNKypzbzP9qjVZf07gGodUbLTOKQYSHTKwoVlUSSg4/6cMYnoczBw
A2tSgfkTaujR5pX/OuJttqS+Ck6XLLAnVyEs7mDAOThChfLSnVnlguVAZ15D4jsP
M+Z9b50Bfv+lQX+T5gY480mdWvwo+vWXUQGapi8YLg/wqX0Ny9oM8tXwREo++Vu0
TmW3NyK7dy3d5PnJC66+t5NjXkythPBKPXOjnWBDEXEcYvG0zU+RZqQlQJsShYeG
SAgtFFGM/fPY84DTULQaIelUWn92lioUmu8/piGGSQ8b5qJ9t7oCe7UfKSTvR4GB
Ehe3dKzbnqIy2LNwo28q9sNhTXbUmUPhiw/CJOSWNUtXqbawpaSAtR8PLOXZPxT1
tr+Z9XjIy/g5Nmm8g3YAaHH/LvxYPUnVMsIR7MMVpLgBdqU9RVS2+OhFA+ZtHNQ2
2WZsqtw1GU+0ZodcYat+4qGI1CwuIyQcUebTZvWVgBb8buFu4LVvvlilUzAjq01/
O/bd7z2oO3RE0yDgZNG/gHCG6inVYelfy5lSD3gCmsqgXSxRzH1B2cUGHjIaBuRV
IDGYI7N5hVKUSvTFLOAkcXZWN2+Iz7EB/wybdPdWBC7nBAiIIHu+r4zD9CPyOkxC
LeA+n8dmIqCrisSOCesBtBHQkwPfJoyiub8i2vkcBGN5gvY6vx+Qryu+Hp3JXfbU
HnTdYaTfosKMMWQlUoGj29hc2LrxUZiLBFyxBijuzN2Cq37ihy6fu2Bsb6YrNlfq
9LmZe1bFoFNZx9KOV2EX20vfI14dnVtqTiJWD6UHy04=
`protect END_PROTECTED
