`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scdMKSHwmiLuRkllJBMYX2GhNAroAKFLSMzykPAgkX+xxdK54aS0KQJ2PKPgfS6Y
jlNyaMaZ8t681SPI3K3mvdpj3yLh95ZbIi9uxIs9V8WM1XaObutSS0VCmG005IC8
xsjGlxQhk+oG0+k3z+mabOCJIKme33bjuUs2haS+ozNsN24Dr0+mEHY0Gkw2Uj6m
z/zBAfmyFplDuyIP/dOMWMtNb/FdlHY4ktDO7EwxWG5J2sJamUQeAG+8AmD/5hWk
aCup4F2wfni7XWyTwkkn1xm0KMU0fqKFc6ffQPv3hEuFoqJ8D10SIqX9sNJnfvo0
hc6m/5JnY4zcCu5gQ5v83J9kFSAHKji9jJ4h79tMNb8Ij3OPH7Vj63FiQ/qY+2mG
VrBMF6+ATuszZq0jxrrseioPlKaV8I2sQvGemq2cay0xZ3ozWDadelOb+yHE+SB/
i5mdqsjJZ+uskU4vLvj/9/Lt8df+p2hVRMnrupHRq2Y2AKZLM9+pJY6B6clO4B06
f46lK+QgiUfavOem05SkKX5JWF9EIhhbi1QWm51w8+byQSodLlTZucSSOols4r64
/LY1bg8vI5gLPe3ETLXHqI2GbFjyLPhj6Kvlw5QHsOMGudt1bCMSfR1i/M65tecf
DVFg2VdvhUwRGPCzbg9AJwz51Fq/3i6rGIIrBKTktiyqc3cIj4wz+RP5TZdhE/Gd
`protect END_PROTECTED
