`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWS3ZgTu6CgB0UCnVBHximy6tAiUl5C2fEISyEpsbj2KXWBh2mUdsRYB9XrlgM1P
PhiLkkq/OCBcmYtjhnHvpGmf5wiMnLToz7sdHhwEg5vkUQxLIBFEXCpg1SiALqi2
mzLnZkr6VIshs7XnYLfgBXms0Rd5ca0EN3EKwdfwioudlv8CEMiRAtHIkJeaGGaK
E6JaI8jF1hfHZkyZ1wJiHVnSWXQwS+qQJ1XdaZk621+Y4F4greVJeh54jf1DINk6
DAsZeKp4LJuuRelfPrxgSpvKrmbNri78OI8GVGn/8ZHzUJNx3lQfbhs8iN/I8pLI
dgP2o7Nba0hKDnz6B6ZD5zgeN/kqBFL60orbfdyzIetlOWlTv2dYgBMlFerQj+Ih
KkpXuh3Fhgv0Gd/GF+Bid38OrIkYswgjpW6o1cf10Vazy+3FxAOPhXx+5/1f8Pmp
Iwzm00aXbrlHb0V7x4m/XD5spmZ8Hz3Jo8q1k6aoVO0/+kI23+j1YAXNHkBWB17Q
AQEd1/bwj58/n2L31J6ZXt4paj6prC0ma1B7/W/s8PaoloSL7xYsl0kALuW7QeT5
mEnHCuPO65ppWWA8AnLVe91hsOlBRiHzli0Z3N/iCFXw5CCLKZgcc7kXZ2jXH+Cy
WTEtMGDqq1tE4xuwaMusmyC6APBc5Ol0x0CmcPi2QyJ/xZ/STf/1o+6S/uhUMJuf
Vi12jK3fKGBPD/syCZNvVML1NC+bXz6RpjBtZx2Q5J/oE5NEX7yK+Wvn4fXdkr3K
y9wuKqy+gm5CIveSRPasPeevM0NskbDgjuIVS/8EQgjSqoZmEAIRs4QmdXYmEuHD
JNmx52fyqr7V6Oki7ABVMB88CMkzhH3tJ450/gk1eEWpidGbM5hiwhhtaeAM0MtH
QOh7A6T7v/GKkafh7rHN4gX3AXWfW09Lfnxy/nvlTbS+ewPLG7x7pdf65B6QUzbf
lMHo7UFq30MR0bFihv7pOJ84apjo+shPCuL2tnAHrnm1ptocWltWtU4fNjQjMfyB
6WB3tVwnmhYCJobMT7HR6ee1htgYT1usLePBLdIIxTBDkZujd2JdKPIOsoqTILPL
fkyyBRtgw/fAbBL5zBrcudFQddmiIiQ0yuQb7GqZJ7U=
`protect END_PROTECTED
