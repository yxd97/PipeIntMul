`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0ZHv0ob+gfMdXrIQ/qRMEO2kOZ+TD71GtZ/2eZIPGllixvK2llvaGpnWL3+FwO15
he/nVAz0phExlMn6BbQct9CDt9TjOCNHqfMpCVcs8msq8d9daBB45zyj4mSWqkIJ
8fC8TUMSmskO1hW8J0UszdkpGBH+6uXEUV8L+eKcS0/1BmU66xzXEctgDdvVTKTH
YyfAX1yhNv9ytBWv7Ykls4WmZAcslpRAftc+8El+AUwND21P/x45xwWPX6190VOr
xImYFH8GKGw48XlHqulhtEYWc5JBm3JsvouitKUCG4CFy09ZBAr4BtM8RwQAe5Rn
c0W9h9myky3Aajg8H9loUm50NjQC7wcVDKh8iHcdf1oL+B6hZSz9SsRK47KvjW0U
iv/nCPRUhcG2IsROHnHqJcnA/TLs99wR84CLgfdJjwY+TUQIr9xdftxXjZbXToeO
`protect END_PROTECTED
