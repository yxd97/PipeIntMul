`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vF0amxP3iniwl/57VZ9jJOGk/BEbOefwcIcsex6kLfN9jnVIhYtrwOTpcF/6Zcmf
LlfpwXjzrt6/yDrIxspwFRLZWe70ntHGcHqssxDForVY8ZuXiBejUUgse/AQmowm
EIPFloQEmJre93ahUreG0KUPQ2hEd5H+vQQd1DE0gw5DAw0r5h3B4dRLYxmOMQJr
hru2a9aeMKKCHOAo69xLA1JzmESIqU9xv4+yfWtKItDBa9UQJvVa33mM7i3Q5PIX
cLlc0Vyi/CWGVBkTMYy3HavqPD0E0Mg5KouJW9Es0yZprjOlypQi+PZGyv1P/VK4
Mcw4g7bBcz/0QMz1ULRK50NVNbuoCJBvo/GN4T8MBly+4M2Yg4HNky/y8noifTD6
kNRdBC2mnawmDPUUOL+MIcQYdD8vaBR1wgznzkdGBrZKM/ItH2IX6/HR987iGwB1
mL/ZRJbzQRT0bgy94y1Bdz8ThAgd7kG8Q4+Xzzr081I245+9R/l0KU5kJRkGVLer
0moISbZiP7uy9HluuDTlE7VyA4dw7KXyJkFw8e1IYSMsjocvLVv13ABaGegj+BVH
PaHS0ljUaVVd3UEBgqdxUxB6SZzbID5uKSnQktH402u1T3EjePSORKthSc3DZbIc
`protect END_PROTECTED
