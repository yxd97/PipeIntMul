`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HUoyUd/YyUtqfCUA+K1r/BmVeESPftGgmQJT3yBvQQv5qUbSSF8ELTh7KAm8Q6BM
PY4+QnvdckNEeghfdihPoNZgp1j3zoHYdgqft2nBmxdOqP6noAhwVQFpqBoxsCjQ
j5s1g9ud6PRomKGQtgTd40ZD9X6EsK0Y4eQqpQ9p3+iPMjzCa0KwizasuI2MprF2
KnAL8rJenRhDXvd8Fm97lctfDS5OEFoS5qXZ8SOJc+lpzVCXE0qn9Dive8qtd917
H9CHLc0OM1Gi5NBV1YTXaDx+wS916JLN/TNCZnqhJtBhJVQP60Ad/1PuyAD/6RLo
uPiUAvLcSjGCbXmsF6RV31VgEuvRPRH9ikyFa84cFsdHGqAiuhw+5PpbbJiufnBX
vNCYo/XoS7ylF3TFz2uoLZlJmVH/w56ZlTD4p5MZe0EOg5+xz2c1cpLPPo75HAWv
`protect END_PROTECTED
