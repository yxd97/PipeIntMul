`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R/o4+QqahSvpX9BMDQRBZXsGD0NHJeL455iY7aw6LBCEVic+0G02JBdn6+P/bOXk
rx3BUI89j8urQVnCdEtPYYOg7XvBIIFUDTHQ60nkZqv6yz7xXKpGhyQUhol4IeEi
tYDDetOhShRLznRMI389JAoJMcgpL5v/j+ryZxJBifxsqGf+PbOe7t64EggD0Gmh
QtibZo+QlsoNA0B2w8A9k+Nc5vlL5Ku6FkC7q9vuquz0R/idYQ4k3XgiGu/8ztnl
xHIv2zxGYgkvjhTN0BSXDaPq/UIhfDTHUcXayJNl2DT8L/Ojwu20eYoi0TCjbMqG
AdQScVgH267kyyTnywWVHe5mDAYjhkolnGgMUnUO8jnYRgwa/VF/L4YRsVO15uow
l4q0JVXRRf7jQTpoK7FvTtn6rjIqT5LxM8+oD37tC1PiHGkR1bkLXkLGs7eL29Uf
`protect END_PROTECTED
