`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QxFmYT3zlhPT4DjAdWasIAEJmt6nXPY1tXadvtyhMcvL9agKtviwSIWdN/ItgEja
5hZjMAHCvmBaeMI2h/1vxP52t4QXYHxIQ1uc4TENGMURtnQlR6mxBA7SZ48kmkCH
DiZ4dnwbz/PcvvxZXjhe1oRm/qnoaZcTEpgWQQw5hXEgV89i8TVVdBa9g4ln2o4i
0tILK1rTw4qEsG3chA0e7EPdiSQ8MF1a8naBufgFungh/ZwY74l33RwY+RYNQNnX
R55VfGz0fR02ID0TqmcxY6b/U5D9bM5vc5xDfKQylStf/5KXvkipxG1UqcweGVO3
`protect END_PROTECTED
