`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hxKuye4p5+nZlWry7+jy05/o4yHmtbcmCdi6b3g5gZq135ZKKfRNjl4Glu96BTvh
BlRBKaqpOCnC+j3p9mGpk2I4/KrKB+Vp+CKiMT+5/Txwrqi1dv0aalJ41OqRxioI
JBSjDSizmmVr7U1shkSt1aIjgbOaIH5tnkiypORpQAeEXDe4vVgjOp0gSyK/kkA5
LJAhA7JISOjXx6GDC34L6DmQdYUwAIwGd3Ctyi1G8l22lLTx2+xx1ZOjbPO04T6u
D5QhMrWI9Z7r0pBAPZkp5czSMSKEu96415SQzyipL5wUEEvnFs1cIugvwVKuasGE
lwh+0Ab0NPYLOMM9DEtPn9+zkjH5QviF4939was9IKQEzeIbolig9TUaB2unlibz
DcZ6/zYrVlQbEk4l/B+tBO/fg9wLtR39LyH1PVrYbIKNArXT5CcMu1C6yJyg7Kut
iDCqXk4qnC2gYW3glo+t8NfPenPz1evfmOW7Sn+XOO/C0ROp3ZBPatYQ4PmioxaO
xVmcG5TjxFeejoEomJ1PSTk3TzZy2p2nJKtwJk94CtlgZFxxkh3zR0jWG36aUrdM
lJTkMgohOr9rpRF0WbkrM0jKHIa4n4m637zTeVIWk/fGOggpT18qFbI/iGx9dxYU
/6iPm1Q03KEn8j7qz6a32DIX5vJLsvDP50SDZ8eszF1hleK3eoEPuzLURzL7wx5T
9OgLedZTB32h5Zmb2Y/6s17rNRqBxWEViWNHV3Laxgc8sYT+Vy0sQLuorqgCe4UD
cotFRW6HEd43a9yls4GZ3/Wk11A85AdSnQxYEiIkcR5uB15OqMJYQs6/Zhl6NPpW
hynldl+0st2QtTM9jC7GSI55H/ygToy2GIlxA23uJK8u6ROnycpjSqFcAlGA3E/P
HTvzjKoBjVPm0a7TTqMk9CtuMhAsKHiZYFYPGxRd6zkrR7LYWp7zP2W8wcN5ETBg
zdtIJbwLmYf5FPzKBXBi8V3Aeu/T56zak+2iYt3zEKvbQVq0iQpsS6wBTqwBVjIr
io6ylHjT0imYxl3b3BPpsF4RFImoNaSHjNDVY8uHKC4GO2uWSY8ZwTyFaJzXF0Ut
ghFTJ7toe4YpQ765x9Ec5kAs6wF1NbYIhE6MpYAaX7nvbiws1I+ajlVv825zBpNa
3gvRfHwvVqTw4jh6r6f/BHkLr9kbGIp1Lu8fLEOA1cqjWU13ZE+JQIhSS++h1Veq
tWDNWVSoEfR3QVEsnH2F1sQ94D0IFJGLAXxI+wyuZzI66ALoDYR4+47bl/19GloP
JyeM+o0w/yBuv5Gu4y9U/nSxPgqUGlHg1oPjyk3A6vpQF32OE75/kI4yPTpSRpnF
XuH0TnClDJleAnzD7V7m686DcADkEtDgSptOPSOw8+lbwbWUQ/HcaPcF5frE7MTn
XabmqchfH8uA6o5QKfIiqGrWma1AthtQpsXinlUXNmM5VKiDKTxNznW72iAPuKyY
P3/57VJ1CDzRuA7OzGmaRxCQbsWWcc2jtrLzKTdhjo/hAhWe4qBgo8/YWyTpT+v6
JwSc9JfnGPzy8X5NN2IVJlLMmvaAAhfW+uy6ofsYKWsO8MXU8VRPIc4FqGlEO7wS
0uXeR4PHD//Zzn3UwKfR7HRHXPC3J0eEli8j1B9MiGNZWFCci7d6mrN1HTb4akUF
PPwYbmPC0fUCwqfA8jF6Eg==
`protect END_PROTECTED
