`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MPzKogibeRJxslzGoA7xk+3kCpq8YTKYkU2POS3OVYuW4tlHM5MmBbN6kTe+ZtTz
VWaJjnNXnve63xFjrqNdoI7u3zown2HCnm7+SpsldIvMzj0A9t9k+rZ1to7lujpi
WDGy6gX2OFwQd1K7tCe+EMtQqc0O6MWKgAt8JBPEZMyUZNCwI3N7tiTuYJ2hQRPu
tX/53x+rimA2lydIoxEDYGNU5HjwG+8B8/2BtZBCx0PfOJDALcetT9Zi2fFWYkH/
skEkD/vIZrNouawBaZ1/ryzVqTPD7MuuOMa7RrUtxDYEPXT6ISsw2P76bwD4d+ZF
3JEF1TCS47+BZzvkR7A9920zQTZQCMQEL+LWTnyyGVjVPNfQMvW3lvnv+14lx+8C
LpcMNM8q1hQ2AG+tBetYX924hNM+kLbWi+4iglF416fvc+U+jxoX2kO3NlL7JCRw
IwdzFnVGHn0xqi8dVgxGlrvqnAYOKIiMOKfm0CRbkwg+A/BDzNmuQYJVJwPRPA6M
rig6/aCZNlCqLkzZiyhAUl1rBDRgCH959nOPXySzk9L1bQUeIbcZHPxyw7Hx2lNe
8PQigpaavgQAa+xq4tJNrf0cZtZfO2/XQZB+JF05pI4AMwpso3iDOamKEuQrO8eR
NBmuWXxWJeSxOP8Qu/w1vqXth3VgCC670WAu5ocdjqVr5peXCgfk6cUgx9OjMRAN
JOglDX2kwM/Y+zPwM3jA/5Oxn6SsgWDm6k2Uo8F5deGimqOh6fMTUxez6Hcd2rZQ
HHi/T+1MgELmdS9JnCYonF/y8YmjeItw8LjlSfcWhVo=
`protect END_PROTECTED
