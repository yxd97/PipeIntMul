`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QzEm/fYoibUqRDs/QBEvGrQgv8GLnayd6/L0m6EvSgAwogqSRncUZeYIGcuQUIrc
vFa+sHR7R+H8wC/4EhDfjGBiTJqNNo2KSoMOvhTg3iyuchyjZGs6pp+zitU2Il8x
3wGCoMHvVuJJlRjFzWDwbuegd/kRqgH59QzvTySaNySY9NSZOxJZHCE/S3EXchvp
SS4U1IQ23NokP+meX0dcAx/g4X8sGZ9b9DE+kFUhIM9gdmFGxg/fUvKsPLXM797O
WFyvJ1s0XcrlZInD4bstYPk+Vn/QCStJgTaUKkBEqel+l6nImTx4jNRNv4pJJA2q
G2KaOkjNdfHicuctPCcsef+16DblA1lGki0nCy4Tcpz5miAuMfaOTStBgFqZZlAB
Z7ruE+A4BufKcv6YXB57rkNdbvnltfc1/dsww+TVkBhaKgmYUIakVN0N+I7LJ0KM
Exqtftv+bFEWPzEHHD9bPNwgaCarRaHRfxBojZW/q5nfJoCixNObuAMAwenZcTHa
`protect END_PROTECTED
