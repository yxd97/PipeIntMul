`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UzuzHEBLqkml2yijPauRTXxK1KB9JfTzC2O0ztrvempHrTqKTfK5r9ex11iRokBU
VFKy8Hng8BNMUKO6izQcxoF/ZXSDc/+RSJLF7vtVyVfWYL1P+bnR5WHNVwArTK37
d1oNl1fkzExB3WaadZl+Guox7CP2BbiVSqhs/VjonaVqBj/9XzkphhfKEe3BTGFE
itPzXaFH7v3xwHEh+pzkrrrD7P0syN8TCdDYHwsbngNkOrdkkuezrGrNfkgpEifv
KeK6igUcr7f+DaVo2gd85PKOJhA43KEvqSzOETU6lnmu+TfAImpjv7bnKM9mZmjg
r0kqsPqPef9JOHZA9K+HpZddv37P7BxWx8txYjxQnJatQohZp0LDT2RKA8plPcd+
xNW9gYupRqnriInIIsioCKkmi4foIKYmx1srVLs4sshB/q/3ScbDUIRHWRqc5BDe
i5wzTAMuJZe+DVKLUYNVQi/cZbhxUy+q7Dr3LUisbsWzL9m0TmvqSazHrYFCsqy8
3P0ukM8by3DznF7EIYOCw5pjdZSkiY5/qsAUpYiD3vAoTkYjMU3CTWZ3QkoPOgs1
cMqCb8kcurfEnCNOmBi7JfeQqTohhwNMKE+hjwEBC9nI+H7a6wVGbSBdeEzsJIyo
oeGNvymdMpxuHmhYTtE82Q==
`protect END_PROTECTED
