`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kttKARzaQSLoJxgW70s1BLnoCmAHJSi9kP9+kLcen4vbP5abo0GJ8W1Go4b1KKs
hCr6TTQAdazkT6Qg4ZuDd8PiaomuwESiPnlU4I1oYoSFJceEuEN6c/goUxy7Kf1G
fZQM8Ud7Wjz+ADQ31Qbk31tG8ssyreJTRlJ24OwszA46bzrRSXViED0L6UWT8Ll2
yBPKD1vXheWphAYLa2jjx+H77lB3/+UtiSYHByePUzDFWL52tkrjaZNU60kBhwPd
8514hmWMZ/PfJUQBAL96J3BwRByPlTu77XJ29nA7jY5Xr6JsjU9STPDvUbK99LQA
FXl33DQiPeQ0BYKHfA98xEZUXIfCfQPzKjv4JLue0q9+81nCP/+7TXOfWsZPjyze
xWUsFdgFiPAammc/Nd0bGQ==
`protect END_PROTECTED
