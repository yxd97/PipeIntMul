`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wPHi2rm/zct5QpUPW0/8QJKKIp5sxT6GBvzhkhlkJdDmapFdHur17MEqKlgE9X51
sOt1vSPvoML+zp/PHgA6DjlCuCTwMpfqnKeOURuM1MNb1WANYRbiTvEtOJOxOjpr
YwGdSGkZzHD7RcQ+HJ4TxOC/jDyW1ajf6m+oOzgqLpP7ADIOQRc1WgWY6LY8X/VH
A8tbjVM01WqjK3vgSVyiZsf7itStgAvwkqTbQ0zfigxsKoRBZ5ke2idfTVzC6YNi
NR++VlFsu12S7u/Aeqe2i53nxQAS+C2NEjqDSU2gZ8NpSggYiNuljiiYMUKJ5JgB
dWPsqngR8qKxudrWrWGZdFrsZbGQLi+PP51vOaqoNie8Cs5ETljWdnhCBHsSpLYI
1FC5Tunjkp80OPyg+Q7Cg8ZOur+I22mpvwffvUxXoCcj8Ar2BBLwwZvCZEPt9BGz
QkzalN8WQc0jZRKwXfRktrr7P6B6BDiLgY0b6A7GARY=
`protect END_PROTECTED
