`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G06xVxAFZp+Jf86JPGpwRXu5poGPrrjrcZEA4i1bpvUgLDsYkJxPYgz7qbBEl1km
0Wvb6xSA8p1VpM5COV9d670sZU6iepMwxo6ZCT2l6r7NLq0c1zBgCQ/6XRiJUBG0
4h665Z5z1HdobmqtdIzTgku/8sJ3myj5U0vIghZz4uCXHtiuEvpAeATTlKL7PGNi
qVEkGyQugYxNELR2dsWz784mBLft/vqVoQ/2RKdD2M1JkBuHme3inCV2LMZN/HO9
cbB9gJYfKEQRGL1GWnSyeQctuNS7p9dQYi1t8k+LfuhSCDb5zZaVRsDuNg63H1TX
CwNRGnoPJ+1riZ3wMZMy/nBjfSaSVntrzHR1U21wBgib08+UcAJjPxz1ukvCb99z
C4jX1IvaTXCN5Xv5kE8KAsUCu8Pr4B7kWSTvhQtFykk3qqzlO1k+7Iyqk5n1n36E
`protect END_PROTECTED
