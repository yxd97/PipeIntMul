`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IIsoW4R/yg5hR4XCWTV7ovJNJK3XRyjwe2Rx46j66oYEiVpjOODADc5YcCb3Q+YZ
8etmZaBK1BcGb+qdmJhywVlbGAUm31ZzbVDQSv61ItQOkp93Ar4iirZCPkWFjRcl
OKMhGKSxJVxbo3K1ASIG3/cX651Emp53kCHYtVMWDKExkNRuZKlU7Zr3WqCQTfcG
z8RmOEr0W4XkC+Ysadzn4Dm3tqkuJJAYZf9GQLVF3LYhW7/h5IAMcQDvOoBq9dYS
GuHPUySIIJyjbgs01bmySCNnjSBCQAianNovFoSh3KcBfgaSRcQCgarCo1PGAgli
Zds7Ob0agsy95oydU1VDsHEvwpAktfUVywGRwJoLAtkbYzvq8AGoRX25z7niw6jw
tz6F4f0I+BLvZOWnqhIzI8aaoOg84xBve2CHkvwfq9EkHIlN18BLJ3FjpHfxbi3J
hiGd07xFMPOuAkEX07I5AF4igo6MGb7pjLDy96RZNAfK9DTS1SL9/SJVPuNfTCp+
/fclTcPXOIZHp9sUDK9+VegXeLjRO6h8/NxJFCokFuchgMey2psgRRmLEs964DPw
wTXcuzTMY5xtRYzKixzKhXRtnb8Xv9CYXuzIW8NHJqibuoziG7aE4/3d2U9SLq7X
vNWausMauZH/ke2PGDtElE0T3GYP/6hxFEPm4PEhg+YKW+7yyO/9vs/Wa7pRgXW7
wxOVOQL7QsOO2Na+5Iv6mGqoqMzS+I2eQghlr27AiYtVfzp4sKVD2s6+BX1cFeYx
a9dc8HbS70UczLXLGiY9TJZvOHOQ0tSywsSh7/WZUjvM1Ly5FFlIqPk6o3l0lQhi
uyP0vl3HqMdpEnfSP/R8srTUpzGyPiMuIgYvruoULe43JYQYFFr4Wr9cJotl2pd6
N/Ub3iTPYwDhyciBFK600Wz22RILv6xwPJ1wQNtwggU/YPa0EvuCgvpAJkdz4llP
3xlG0tRwQ/3CGlTFpNLjsJfngwz+Vm0GVSX36xhhKRcxtdYuRJ4UmkulurxtGDU7
YDWgRMHKKxYmvCU+spxvJOcnOtD0tG5ZRmPxYxGsyOxWbGJrTuuiOVgB89FWoB0b
IY9siZydjo71txVgwFcIWP8i31uj7lZyez+gpquH0g1creR+hvSMEj7rjet3tSxG
IoJe9ogxuAA18B91goecIJQ0doOD+rRMtpQQY2uzIbWpfFUb1JsOjQEeJZhl28L8
tDlmhAsAwdY/nQ8a331mzSzxgd/RbvPkjRmRszdMoV3pnJrXq6Hrlj+iC5ZKCNAZ
DuMZrS2pSFg0j2cPBuopl03m+ozJfhvjCCDU9V7y/vHjS2zfy1KSdb7keLO1hFZy
NENa4PVXJcejhkuDnwCw7HrwUiTK0P2tdKXdLz+QUz+ogCvztU0CCPKmxbIMUG+X
p1p8XGGrAR1UpwUry0ALla/aEHCZFODva6r69CJD4Lu4NHPJ7J6eAx+GiMLfs0k+
fj/jVTz7RdDyfAIxaSiHQwAfniS2hZ8yO5ofJzMpJDMUnKlQcyPIA82RsedoryFV
Bw0xOAnXYcMkvHUZ1963D6NFkzZ2bJ90DMWSrFGxF3MOyfSAA1BoQZnDbOgp0VCu
9f2C+BwB0n3Z2bDF/yN3nak7+eY6c0dZewp2bKg9kfs2BwmllJWY64p3UFHsuDgM
zro8bSuqS+YBQv1sgKy4CRby0xVhZQnMmZZRs2Wlq6PrIFki2WZyezrw80DfMzGq
QwpJ4QxBISVTj2irCK/fX/wyamn9eoyw7fjSD4Y4xilsVv9emoSfW1q+4SP71/MH
bANigUbAuo7ySkBikpqGlM+WECI8yAOx4JxT5SlwzQXu0R680ASgDkNdAvstZUCN
Vtun4IB+dG4E7M1JsugU08FwpwV6+LkznWJnUi5hqvgTXpL7bBHdez6HH2ezlEQV
uCr6C7eBEHZ3GbmVGmtyhxyVJZWc/5Gspi2vHJ6xMJpS2XpzjbtfLwYn0D0Vgzz0
THoRTlO+Xr4n7+s/JFkid62jCIHCgC2tofBF5/3FS9xytzZa2NbqZ9gOrctKmvar
g4naOR+3xTUvub8lgA8oi1L7E+tjv1PKlmFrAc0rvdsvejyPmIf+yeUKhsfkD6Sj
iXAjr/TaLaXcblZB56Yxrjte3HPK4h3hh2kP8ckvm+X27PuPhqnl1oARHauGkGsz
wTyWpnqdRW8mc22WV0+7HYeGKYa0DbkyoJhgsusO1vXwA58FDxnXXtOnt6DmDyV7
H3D1lOePaIx7XZw5KZTI8HO/LJ0FsojZ+aCi58w607Nbi8VL1zeOc/gvN59ryPp1
5Dd0LzMiagx1RAEenjQBElNKisgN9oiJefk9+6rO/U+j4CcWMmkhVaSswrp0/Kue
j3U+9Gp6DxF5qLRr439Wgni35LsfbUgGS92vt6u6BEgJDJ+w+lvzV8fSJsAnC6Ks
PF7uBr3eT5e8N6r4nBUWOtS2kRjuJnaSiVODRFRn+gT4FgD805IBZUG4D2tiosrx
prZZWarB/w24w93IBMY1uPojuccp6opcp/Rhjlw76oSSy0d3fGGoADSHRwTKEAMg
Qo9qXcZjUFuwkfmA8F0oKGvGH8Fxxi7P1QIJblhLFy5lBpGL6OmrXDF9HZrtZ/FI
HuCKmXfp2sBuxocDPabC55YyfwzicJrGiiVrdDKzDz0GymEL6yVWJXiau4VergHK
EcvxVRrogIC46XQhhIqoKShpGhL4D8cMpeD9UquK+077Z2RpjB4kHbS8clBjabTl
q7uc1jH+bnpbFe61/Ba8Zm5EzCg/+xgk3Lv4fz5VowQNLX+zynsg6guDrAwQC1Uo
SH6f0A2eIc25uFJGFI/0dWJD21CkUPQe6l06yPTMMevl4U3Y6eO/jAArLHi094D+
GlvJ+eu2FwEqy3AtLu18JVSKi9k9VTJQ8s7H5uQT1R/L2lwb83VHwUCKewDyTkF0
tTZljc/VepVKyqQyRlH0xp8caGkkJIlpkpIwa+LUzd8VRxbfVNUByl76AA5AGu/y
wrzkNVz/GltKQ3r5YgkxJAoUVM10IXTGYSiUEsLo8T8uJvEFMdLThR5AlZol1R8L
ax57c9JvbxIoiGZ5lOcwegN4bKkUBHVBJ59H1VVgT/2NrnVHnbkNQ+MX0cMBqYgm
tM+C49nFZuJR0EqgjYaMa3HhbMbzGiOHdwGdmgx6JNDCpbcwkXLoeAQFbJ5h0xdq
24pkFCzq89vgLgly7BKa+p/IRYsy27YbLsqROVNwswuQ4Tkq0SjLL9OSL49WhrtC
OP8KxbLZ47JdeRYh3wHZeW3/QUftM+OTVhgVo2CkatWf7dqjFEleorvqmum8CWZu
w5sTIqbagHznv+r/EaK5XvKVSm7AEpbPKqIyC3XE8HqA29AVtq2RHp/gxM6/xatL
t+0nA0eK87NKTMmdIewUr6bWvBxUdQF/LXPIUjYKkZsRSWTz0MDOI3cFm/5pAQVS
AQ66H9ldaMKCtbZqzYs/vB5iYx9jryKWzjsjKI8bhiAVC9D/aRLehxtvyuWAYgOi
yJMQGXGFmq5n1m8YWmB4os+fs5I7RHseJ0Aonj/FgN9NRGAVmrkkfA5yrxWhGHcQ
sZdv9UM+iE0CEeO4wnfcEx7kbeEqjJRcbb/ibbeTiXdyPN6xCK/rEBNmHft4DWJf
po6QGCYbpn6S4xcl8ua5Z1xBoRbjhu6ZjTQHrEYOaEOe1izO4v+GGPmO+crE5nMo
mZ37si6tVthh1efJVLe1J6BRpbVJSdGjmmDrJd9Ufiv+8WHNgj+fBPeHwoZxMYEG
pkOrsk5F/jeOsqNpwGs/4g==
`protect END_PROTECTED
