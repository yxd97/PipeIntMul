`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NC2HEXmyEPoaRS9IeX6pOHPngDXH0RQoWC/dyF4dttnFlBDl5Qwj4L8ZYpjMmXm1
JJUuiZvyVRiu9rAGEnSsad0n8y4Z84DO/V838rDNIf4QrKUIByMZPu+3FTzUaKH5
IsVbLjKA5JZXFmBGxfkXhBYIMuI5vz0EKFkQ6sxvpHTqcJKY+jasYW080qCbSnm2
oWZqIEWMcz99Gxn9tCLTZCr739Lv+a+T7ZH2nsm8LNCooVAa9szi4cUHIYRLNET2
KmhcR/rGV9VvHWcABUkb3w8MBpiUH/n66iXNcU6p0HuLsxVMpAIW743DhQvaZGLt
BUQl6J/bBC3CxNNwnjzAqAXgk43ZFTgjKDtobMPCAv7+FNP3AFZjeJdg1/AnbyNu
hYnXHvgigVQq1tROX6W6nQ==
`protect END_PROTECTED
