`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zowBsVo4+cr6OupizgQpfvbqQq52bRoLXTl2z1qg7F93FHbgWbttwRy+sE4bCB0O
GCzAF2NdXhAp2b3/uIGIyQ6ruxYfgsLHw7M5xnrM8JCwX57niD4vRyIe3JTijuJ/
s48Wq6EMPCLO3u6rMFr48HzAY03XVZilK+bcsYvvC5Z24CiaUtTjZhR3nJpvyKOz
/NPaG7Ue/0HyTKcYbfEaN9U5l70RJ4grzp9wqM/8NbGzESyOyXoksY32bLKBKf6h
BDy4swftBYoV7KTQgHXfaiD1ryA7ZweBIB5rMjzvUH2aA8WMtvfmUIXweXruhGsz
Dy/ew39+4n0xh2g0Opxeo4UKBEi+LxssMQCqDKcqTw0LeraNBmC8Q0kPNjWkP4yt
QxbY/h+mTUAHtluFUFuKod558r7LhEeS1lP+aCknd/G9JrjXwnNk0qe1I08reXp9
Ka9rMhw8+r8gAk33wpvBP1fXYoWXVpH/+IW8I2kB+6TIey3rmEcvhuX4v3e36g2m
MLVTRIy8buabM+AZ/GQDslfOQXiAYLihEZLvth1dfco=
`protect END_PROTECTED
