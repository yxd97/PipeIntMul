`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W7rHJeaABo0rd5iBlsjrQ/qU9+sxY+4WvZWTg94ATP+D3No5xj/yyCmY//5I4DbE
R7HqEfakhf6UFrKpRW21OR4x2NwJinmXVkcVQ4AajHBTp5janRTcAGxfHt7Im7j7
KXprXJlwS250YFDkbINn9eQaWcbQpsX8kCQbnkrxrPETnErcjtOIp+Bxa1Y3fTGa
x2qwRrBpUL1bDf0O3bbEJnKUb11cr3qgQ6B01S1vYE2P2hUlaNrQ956A4Xykoln9
HVJj61MOnk7k5vsfuY5u7W7VspTahCe/3pp6hc5hyE16aVou6AlPXggI62tO3Nx3
07bGCZE8NA6JbTp7OYKMBwBNAwtIeimVyRAjtti4KhrqXh8MmIVX/5uUr8fGPDjd
64VFjfqoLU7qLNg29vd5TuOU+FTlxhRy6nbDX4jd6rsop3wegWqFJCCog36m12Nk
0f4p0F26pTLnBN98yCAQt0T4vpj9vd2pUzW7dGbPxB1ZB7FUVA10QQZg6jcQTHea
2dxWbBwA0figxuOJSmsBXui7o4EJ3spNtVufNcPWHHCSqC7HFMw9DsnEPNu26mue
wTL/nW7eHOBhtXcxEfZkeoeQNAad9srCKA++IwLED7gG+9PZJNT3+E2D+G1Kg0da
J/rRKzl6XDabY6UzyeRyWL1y9rIHiZhE3LqOHAQUpaB2pFmN6WO6CHR1rUbRX1Zy
AvqJYvQoAGFMratTaikL9JtKQFc7CE2DMMPafXA3QSrChVaNV61lx3OueyG7RfIN
TLnY1sSlLuHX3pnobvqUqQh9+m+IG3puDp6/+p59AsOmu/4qL8X8sP2/HfDuYE1B
xiDlS499ssG/OfNytmkgVlOeT3GHI+NBvSuUeTk/ChAnjtXlqyoRBSdLiQHORm0Z
jeQZtrS0zviYakFnRsl5EymuCqYhgHuJCVMI/wMzubBE1uAWgc3XhC0IB8ET+8OC
8SdOEws+a7qYDsYl6g43X5+7aPNF5Uc5wJ84SxikHWJ33ceTii+CDIqLw0VMwNJt
flP47ewyjxgkXeQvpUq7oww3ZPYPP5fBOJiQXdRDgYGEyHaweKWCgU9827w5anP9
d88H8DwuzIaMbCqYcvnPD4eZz6puxYoeI+q95hRc39E8/BDjOFtNvo79VVxB07F/
R8IBGeAiRpB9r/CeRjQHRo27EoMTgIAjMbe90eMBpP2Zk2KD20mE6BZi8GILUDeZ
6oTdBYZt85jvBMQXbt1QfYkEoq32OmdOZmu/SMD5VwJPJvZ2Vb0A35in5K3PzhGa
/vX4q0umDUollxVoZbT2s7QawdAgbPKeU9WRGlzIFWu8brIqAgv4QfywO+YEGWdP
OC6iq/8C8ZJXMPYauf66ebHjTRmcZwNP9Q0AuR2v38tIocDAI8INaGfudnTSqJh9
/we6tKvFS4/K3jrRAPnmAtStqjNdHAc5GZCl11c35J5kUisL/ELi4Yu/5AzjRzMn
2NxY+i6rXkCxLmE5dJH8WzYLwOb17OpC4Cm/JgjSvWAr4gwApqdcaWw5p9aI2auv
cC1725WORdULqRk6UsPUWtclPjexAt32au7AL1x/yES4LwLabTjZg5CIKVt9uWSU
jMAIClGvNvmCZ4SfVMSHGpvEJdjOT7hsx1jeaUtVdMFPM1XumEW/w1oapriVxx2j
VaS45+sbMMB3JxBBPwX4DN6c8fyfxyU4N0vgefJez3100E6K7pxYdlFws5SXlzE+
NzOiApAoz/5a9ETv6nVmUUcSipAdDc8zG9qSwttBuJ++UUrOPHPpvU5SEK3/muAU
0zprabdbD1GKIhy+X3Qyr6RSJ78bAHnluGf3/gkJq/zzBdednESRMHiogkoj9pQA
Y09xr51BiBqX9QVZ47kw7z7kl0NpJqLfRqQszxrPQGxMK1Crty3bk+Uo9vAUFoW3
OHzwQrBhwjFR45nfJ3D8GAfmYn9epvMAwenPpOludrPnLHWvwaLJIJOuJEqMmDiy
QvtDDHqtMwOXIO8Dm38rvg5M4ijp/ZddCytx4iEo0jcwd+1rGDg+86HnqDdngi2s
9RIkt8es/BEgAlUTOllxIvPy4N2GjnZyNp6fGcgNcig42Q3nFc330+QiWHYvzpJb
sbaGaS0Rf6kneJRQMULpfzzIsRt4/BdeWk/NIDgyQhTRr032ghe+jgCvpUjkFh2Y
1tT9OimLz2SOG+op483lR1EwVfM4W3/3eMNfhv7enLN1nDKsriI3SNWF5HyLodSM
0k8Bpn4XZXrxkt0fbhJIH5JoUDdf3n7QnXgrVZs7ob/QzRbiJnEU1kFIZyMT8fnA
0wRs4JxAW09dCUYQHo+7pcaoJZDGHrTrCNyfvJ8gcFkkETYgHJpIKuU3sIQBhWSF
`protect END_PROTECTED
