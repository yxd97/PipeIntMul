`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDmYFVacUYh6MKrHXm19WFlY9RSG11EqhhGCN8YqKYItQU0GvxeOanp9irZD9JJk
SA5B1T/klOFpumF6VlXZ65d96PxR1m8sdlz49T4gY29WPaayZtKJiK2PNQ4S9hSU
qFv22Jfa/kebA9ZdZayUxRegXaVhvV09+w/6q9Rij2NLNfPy0oMT6rbdcOIWTJC0
MFAruUsNcVJM1JoPenfjuliifP1Cr9bGKMFOk+d+0iuKvi/A/NDCTWLBasNzEbnS
mfplg1g0YfUK/ew7urIupBqxJqDL82GhCXGjZJtz/dMmlKjMqpzAb4Iaql+IR0Hn
zw1ojqH1OUckaXX4ZO2J2SDoKhD4kORcj9Zh5FchuP1OhuPWZMEq25/XyukSve9U
+ObkAOg5wD/KzCSVw+tkPU2wVUlYhj5pzxDPOlI8k3Bp+FVyikP7vanEQ9zfPFph
9huRa0PegtlER2xmeQpXvA==
`protect END_PROTECTED
