`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2eA0ioXWOMWB3uI6xz+dE3Dq05UrrB6XWnHxJPWawCaef6uBKxVVzxeZgqAYY/aD
IXYykoArqXhx9wQLf4sde5rrotJSB++lmK+6oHcCb78uKOFGnh8McZwdzfXntZEv
J08KGZ3EsLn0TWw0kJNPRnwwZhbN+fb1MHulIk38j1M0wbzHV7Dr1xfOuaANAhxG
crTQq8MSs3imrE9VLmvzMyetDBaQ6b609yt2vDvlfvZZEesbpO/hHu3iVBSuqwUL
U5gNvAkEx7brJ69lOeA/us1gzeoCaNdvF5shwpADnm4EsbForivGKi6GV+TR+HCy
VaUoYoTyjzTPWZDe5ncb6mg4B0DV1YeLGBv193CxRaVj3Uoek45h4dw8jmuPzSun
A7B4wF4H6CmHCPHvTCp6FXSPsMysckN9G/5G6aF/IKCIuPE9xNZBNo/EaYgLaIe8
F1I10+/uavl+Nve7510n9yknVMYSygmYdnHFlo75PDKFmdtg8UIAMfAhCg7IeEg9
25iq63akGTX2d8djmBAT7ypVGEptX/4ObyZUhe+PTm4u9hJBgkpmfdbkmH/mE925
NalGW2ELKDRVLr1lRyp//g==
`protect END_PROTECTED
