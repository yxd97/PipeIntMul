`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/kmbDfqMaTSDrxZ5q/jHIUCSvq7Lt7E7sFWLefWVpKEgnL7cYl1DkdcKOE5f3lcu
XdnnXQ6f5qgrDuXammulKN5Vq5vWHJ8QAz5GzLOxO564Rm2e9T0L59ka2i6wKMo/
Gio+uJAuPzH4SS68lUcu3deP3cZtBXsbAbcGfgUGT45GEZmkCA/UaaO0naIY94ve
+HaApM0cJV2WtEx9LbQCkilTpJ7M4Y+4jNfT14GlsGcOG+IcBCQhB/4NyJqY5SRJ
HwO6XZY2tdJ5RRK4ZM+wm/lA6sogk6jdtNGjDpIsQgBOvaexAWNsitHpZD95BxRf
gQuzkjalKPtQ0RbDO/ZfL7wxiWEAlD8ZAx7jZDe/Tiv4/8TMKl8IWJiF959hlm46
D/CYPQpH4d42W3Q+P9xZEMaizkI1y8RGeNOWkJF+bdxwdo62QAmbbEoop36Uj2ry
OIksUNTgoGaHoKepktC10IbBQHTnIQlIPP0C0q2wSmyHoEFUNnLdO9bhZlQifMJt
ymmIFkPuGNyPh7iz7CgOHGwT0ff398hD5w7Jk/X6rHiG8G4SdRJkYLhIgV+C6IT6
c5YAFkj2SGGJGZK25nwKiyrfTFwM72s8yAYdTtthX97+O8Ou8k7pX+NduETPiv3N
bLKthBa5KjKkE+Lz3vImmg==
`protect END_PROTECTED
