`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+VdPHKZXxVpmeMuJUcnpFGI/RD24UWWyQct6uac4h6z436RT3bR1QMKqp+hz1lx
4A9eiAWpN3NL2QE9ukfvNjAif+qaSbbJcxoFQ9ddr8QOv/0GEgzGxlMGpjXBP5+l
fXVyX8FYhGYcfu4qPLhiRQtpcw1Dky0hadNhphNLC1Pv6aQi9POFxdxksRbu7XJM
xBAPc+WzjLPR3h8ckL5mRghu0oN2LQqklKdMpOvH4oY+irehwTrYjvSCkjToCjHi
Eq9Tg8w78wKhhaQCBL4fZrH9ZzvV8I56BWQ7EggcWiL0FwIRSnYXOSMoPezMfEOB
Jud8tdXcDKgl70LTZdl82b5d/cyinbcQpqH9C6oXzoHmFNUclTSCtCBflG0/Td0+
IApCbJfTfSbsxByKKxiH9cevUqr2XaFllWaUfcCBLnjCpjHOaB3MsbCXLA/3xFJx
ympLReKC/d/twsxcsUJs5fi/NUNUVgZ+RR5Ac6CFNcs83ICN4eGD4Dq+j1mKf4Et
58HaXoLyo5MnOOZrUTzLsSrALL0sbnPW29PUIe21pPiHisMaHBjpEfwxXH+5quUx
2J+IVIBQ8oWeDI0+s4OqD8P52JpL8dAkXWTg45/YI/jHHYuPskND7+LEoFv5A3n6
3fh3k4JZyeMeRTRGHmh3AA5rOh0XBMRDO1etf6TNEebbJWtMB9gLXIqU4/9Zn9Am
L4FOSRWB/C9xMRFXa7FUUbujnJw6tmeveV8UAyka0LMUFhYMHby+OuBFlGOHUhrj
cDu3F79o/m+7hGhwwwVM2FqAdMmk1rLbOfPgZduDZONLlDjCP0wbhbNNHGIk6fqm
7OUwzD/5MTEsPwdmmIOK9EcP4VafOu9w6S1GkveGGAxtUQLcvMxMnChSp/3pYa8y
rz+bu7LQpp6icY1oitJiEWmM1MY9BzIFxGIHWGKnB8O/VgVVdsivfvIGf+/RAcxK
tnACOCcD2wjPk5hmQxs6ieppNq3QzJoihCiaAHxbly7TaeIbrGhiPvWqTuS5tgtS
cUnDuAMgvPG7gyLsD1a8yg2PxCs4b0y2XG7zgK/VqQBKKcCvLLJSyK8B1pfMmaHH
xOJtfW49kFGb5vbiTVi56UzCpc8frMa+QiSSjG0bzuQ/77/1DZFII2BxoW9nokb5
rNl03uvrvrX8gypRBSMjzpYFBasHdEfWPqfIrbKZMZjEsS+Pp0Pj20DH0rRiJ54e
2xaQDwCorMymFk9kOtpaezwtRhtWNeeu/nAYqtp7V59nm146F0jNzmdv4y098oob
yWQa6sFomgXzWFbQ3XJc6DG8pxqCJ/A+bxGWUivQmY3Ev255/KpVabppzvnr3a9x
MDjFOoxsm/VCZCBRkY0gIbdpSKBiid4TpiF/gYrAOkIe9yqohg2rynK1HqyiD2FA
0bS34DjXGqSpppmKjJxLO+7e2r0BvU9vmOFv/LIjcimuHRXT3FmzklhTHSb/rt9l
bpK+q5XLq2eUF7RsG15h2C/Z9ZsLBTR2qACLNzWNpNszxj2KGC/XYpcYIUcAiDW6
6eY7JYYH3QlSPSTCh3OXYO0+FZQNEUvTUdbMtheYRhmOSGA5+szBdKPuIe0w3dk5
I5ImIT4tuVsb8Bg4MhAiYy0ccoBTbUxO5f4ANGtTiO1QasulP9rmj5/fO2CPSel8
/QHm3bx/avYIBMLggmWkNEPIMfAZ9QSEHGKpGuRtFBm2t5y3Th1LZklJn5A1uslp
ABV3HpbTGWq+5un/WEdt1x2QY7MHVhwPIhecye4Uu7xONOBHY1n/lxDAjKESf0pe
0ln41qCqpWWDbgXw/DCbhj2C5iv52WhBJdrtVeLRjBaQ3J9Wi3snRDsTAv7t+xs1
sjgszFWjENglMdZWnGkdJ0OHNmuS0Anwl903sq5TQ2BsuINhFTO37F5oOVmxl3Qo
y9JWhYjH4x3yqtQCQjtiyAyT7TFCrbVMFWW/TRtFQ5/toZgg/4K/4hCiezbP6RWI
Tr1npM/0FsZYWo093Pl8z1IO8tvYWL+IUDec/n+SdcDl6EYH9kjJ+iwP3Z8zxgNP
CZ6gRDpVp6N8gIUaJb0h0aPqWIqYXnqTCi9vc0lZkUDnoQkR63ZQgeqns/RmikXt
gDsHhXrNjsfrUlFK26CANWYISKup7JQfNAiRRD0XeI5yDoIuaeYRTH5vNg+JhwT5
q4k/WJ74EIB3rDKF4sRK15RNGFQ1goxjtGE1ZSqjSSLsAGIiGd7HzkIv2Kc1YKcn
If7ZPFO4vpvU/B5LX39/tJWzWw2Ij3TIRD+VIJrct6u9pPXR0xY8NwTdPaMhcGEu
LYQGhKNbQGKvGgEDeV4I3aPVfE840tGTSzbtG+dcONMMTBJQZvLwtjuP2tl2FxkP
E3fcE+kGFYchs2an3Wz45Xjse/zTBI3fHpl4KpYwcYe2Rg7uoA5e72t3jzYPRiyr
5SVDwNSbZSZcn9EKb+BmLbzdU5w/OL2RzqFwCY5yFiq8l1TITd4P9wF/4kWmT8Dm
6f8YyXANyDObbos+Ps8BQaiVFN1c1R/0KMEXMQ4JmTcgxM1pC4o+lMfIK2eueuup
7ffVN6hSob8RRTK+GeZrFix9a31rotqTNJSbVpbj6e/dDJMs4hybX5E/Sm8rA+7C
rYG4svyKL0MGpizXKGouO40PoWOxYW1c801kN+FDwtqEaWJNtFj5Lr++f6LpoNG5
wa82KVdjSb7zHfU1rTz+xo3X70mygy63GwIP72sqtrUfLFkO0yIk0PTj7UqVYPNJ
4z5p8emPlIf6wsfHRzdp1H35RiWRPvIKgQW7HHYsR988rM6qUqlm8Fyyza5pe+L7
4hRbeqtZn1Z+mrZy31Yn/e6tp8XSUdj6pmsAhvXcGqOP4Eqcrk/B4r43ZpE34kUE
J1XnkJjAg0WscV7fKGAVKm7vDHXNo6Xxz1kC9Ff3VIF3TzjKg93ede5ACdFdGgCy
5G+iE7mD1a2qaIshqia6/TX0hFDUpTS7w3Snc0EUn0Yjzzy7zCfp/lxNfXlAMfKq
3itwn/fpWaYSMnV88OuGuDDCgIDBYOSqhKUkoHnkz8A=
`protect END_PROTECTED
