`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DdkV5M7QiTLMa0oGSzMAohmH7oHztgts+7FqUo1zEAV1qTulR6JoaEQx0AyVroWj
mmrh4rPRrOlvopKRSTki2lwdHAaxFlSW5V0A55bmsCt8oGe+KFemQO5Z5+xn3NEk
VP2bc9XBjq/CQqIVBWVU8QKNoVmOGf3/uaMBS2J+cbtOcu+uyMB4K5QmhAJ9eiNF
k1xtNRKkFIp3wE/dxqcIga4w8kf4GTq/H4weq7bIsNoGkD1qU+GEJJc4JOzQWR0o
VmgDHnExK9m4CzC8u1FILw8K7mhT81O6AGYcQP/XyaPwNfPfyTKDILJhD3GBv4xQ
BAR8qPAIqqfolWoaWZ6rBpNP4Tv5jf+c6CEwgxpEA94ApjL5ZBLsKukMbu0xgn5d
1EV9UoCS88zmaniXPrZXiu0F70xU0+Vbyofz9D/YhkDity1jk9TihoHEAUoHqyMX
E6Nt/aGunZ3cZ6fPhFGVAl32LS24vtbP5r7QJbo2A5pTscglwD/5/K5WBJM4xi2r
UJhiBeGByo/ufbY8YErxIKgpKUAY8oU7tPGSuHnGt570DrLFsVL5KA2VTYwpKrIM
FcpSG7LerdUQ0TsdJSe1/+sztTtESwD69a/FtiC7MAs=
`protect END_PROTECTED
