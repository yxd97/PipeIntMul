`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vCXtS/18yOIXoXoP680BAmN9ifB0Mi6ZG5XLV1nyK9mNc8mBf7xRqNifn/WZn+9T
3pNqoA1NCZhaEO1FqvmXBdRm4inY/KxNKCB6LEFXfW5EA1w/qO2OKOQAbHEIEYjo
XJfs+HmlGCTwDzvihcpXkS0ykQ6i4eCQJ5fFNN//gbpxJNW5ztQMjNaXDCpkw5mu
OZGdqG3hCttG6xSkNjbwqP2zPY15ycPNqWkxRYYishUkUwKBLUabG84XMwWaQ1kX
GIrh2PfIHWIPhPszMC9Jx2kkMrT4ItFKyL5LVq+p7r2wwrX4JvM8AjmaS072qirE
RvgiOpn7AwEkfAIm14TpqLLe+0fKX0OLQL1akFOYkz4Vc/pDeOez9iomAEp+K7c3
yvuKTFrsefrrJTuAIeElPEqtaeC3BXGzQ6xwrO+ltoICazuoHNKFhZRrRbfVJhKX
kjOgD3OGSERtmWz2ZZeC47KbU9q1dNGkWC3Cl3jZBSI3sbzUfjap8TOlyfvvtUy2
VTIYs/6lE41Sg9D2ZXFbTwgTD4NBFLtzh8X58/9c/UZXzBCaPyxuS9dNRN3Y/3RQ
czxPf6I0C8b/rK8kRnAmpfbvVqmQXUsAxeWp1LMSaWgy34PmLRKyMaMFfeumtqdC
`protect END_PROTECTED
