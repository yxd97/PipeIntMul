`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgGqwa9hA/yTdDR2T6iXfyWJ6SDQ7fnvfsg9ds6l6mYP6Bz7NY00gar2AFC7j4yH
s8qr+5ws7tmz0nPBeXbyM2cnLivbjYmi9U5uIqEPP7yuSNOJ2jdFONosYEe1Whca
YhZdj+Pon4SvlrhBndO7/G7Ui2v/xJllHC69qpikUGtBQDo2iV3bt5+9/4Xa/3iv
GVpqllIsY8UtZUkIaDRkLPxRj+3p56UM7M916Yfzy9nHcJX2wqH4SquEf1z4O/RK
T1xgtlTOpy8VOdYVmWmi2wllecLQPJ4ymkctgPnVndP9tCTVfPAO62noVKevkBuV
QZx4GkXzFHK3lL3pB18XG0HFLtozsENJ5Gn+heGvyDat0TtJBYVc0M071Mic8bka
rxQOkspkC7UoohaKMeZ85S5ta/ej0+m+7Y/xAAuy2BKgmmVSV0CEx9MwEZlHYy7F
o3n+OHDaBDD6DyX+tgg+sQDyh8LfNe+LuT2ULdlgau1HGo2AIm8zd/aLmXKwgajW
EEnM8aaWxlHLLYwhhHJ4HEIyNBRDvd3AzrU9U6lw9FOVhIiSbN48aLAjh/T+J5kR
UcvCZTFuqupdviQCYyaCprvYdDUCv64TxMEv/tKCMWBqd/f/nDvYKf7289wtRhFY
WEUxozI4uHFJJt7CGXJXEJhxnoBv3hNCU1gG+BlvLVCWQpI/36pN8F6VBN8kXt7v
2qS1u+3oEYAhuBxUBZr1xeJoSQk/2eQ1/SYkuorDgmp8cqIENeHDtzK7+T03oI3g
X3Wu4MaIoc5Eoc+odHW9xQ==
`protect END_PROTECTED
