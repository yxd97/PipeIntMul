`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CvCwH6FiW24xjXtgPIc2AA8EgvdCj1nC8oaPsAYCHiSX7vwNFYNigZpqq4Lmo2G1
7nGRz5e5/EriEjZxW7LqD/+0YfwFpQ5ryva6mlrq3lI6K8Fl1DrOtYPVc0Gz7aX6
e7HH+tIT15IDwlGmPyveaQQ2AdCq8DIRyVTvwnpw9FLUV5RUVDW3eornlbeqoGio
9WZ+cJ3mJysoAd/Ng7lNfUcMIk7oblKKna/AK57TKl+RwwD1grMkqii/r6ZfLmbf
46e9icmh9whHTt6MbdTCKwJoiNEyR+24cQ/nObydnEOORjwuf7lNwyr6Aw6xHsSX
z6vsydb+sdYKpJnKVkGgKogsglo0PF7bVkaJv1RnRO6wy4fFp/OJscVG4MnMGebs
mo/Sf8eJIN7IydmqpXwuLGCNl2hWaAzejhzgeOcHWbMlxlvb7/2Iifin/BVB7JJO
AovlOnN4N8wirG/6D91egg==
`protect END_PROTECTED
