`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWyL9Rxm6CtOirdVI7vtcA6YicgbZjclWgdJLYrSwA6/P1fOUoPbWdd3ABquWurT
WfC0LBy4VqMkGJu2S++XKF75+JOIsoCstKRuv40OrBnpJlmdoPisWz/p8HxpTVN5
cz89TFLo1yAQqVPNVo04VMpUAKjoo7Y2skCOGGfO7csWuD4PC23cgvla0JQ/cbSx
svOlXZ7NE8exNumq8EboPT0nHDiQ07wlNaWtwoO5qATkHlObc70Oohkmc0CVLHVL
xspJCQ9G10lrqDec+pMrEwfQezEdgIKWxacJyw52R3xjrWuqep7kMFwnGWfF3mal
12GiVqYAVnr7bC+aL9Trz9HqpKmCJFT8fuVsPziHglfTV2sRtCqwjiAz5LyTS87r
IFFW23RiD2BjG59rrxsi8NXGi2XHO6fJrtB7fhUUvNpXysIf3OMCJpudOWNxOUpC
4R0+nUoCk/+zkC4upZsvR5J/V1ozcLsjOeNVV5WS7/FFLI6XUXM0eTR6FrmrKlN1
AXOQPXBgN+UY32LBGYCyceVAtJMYlnRFsg4cj/iZ0a7YIqIHyGgNHiPPQDwQPzJD
VF3dmwS5HacWHSFLjAsSY82WBSFL4C4ADdu5rIzwIHGq3g0VaCxbY8TzNuU/UT4W
wbYgFVfizDSvHqxaTddQSJt4cGVfLHmZ7AvRFXwIPTgjNC0+jDHWazpObbh/R4Zh
wmxssClbusJ7Ha3Bvct+feX2BxPk7Pau3CyRA5QUwz3ZL15Sy6uERJzJ0T7aDvio
qOO7iBhRBqJhj95z5ZhoLqbjyL/WRndYrbJS6ZXQtJQktiZ6doLxu1gwGElPovNF
11QhX7hk436IgZtV0f8z7Eb9+deLnR0apYtfkhlWLIwO8qy8oDmjINAiqiDeAfy9
nGnIWUKar4yYfBzjHiUbk1iC1Ed1DlzmAmMnKzVcH6fFcQQAu1VSq5aBbKCWFRjJ
CqWc62ou+SRkDA5w1MWu/PITRhA3dqJmXR92QQQO3J3hb0KYYW7cqN3jPKjPfNaZ
pr6y7EkGW9PN//rcFLNq107PgdBXbnQm/stUrN7q7e0=
`protect END_PROTECTED
