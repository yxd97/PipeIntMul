`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LNgdWJe/oeEQCsSH1QwTtKMlHYe6/ovrd5AIkwAfMCiXOencl+jgcN5yypoz7a5Z
098OS4EXkGmNC2ma35Jmj2n1lfrMHW+DCg0LzFcqAtOmabemND7Rxy/XmM4oB8+A
zOOBKlXGcidBbquxGMSgrC7U4sE3UIJ2MOdu13WYVTF8Z1uUS+JGyVtIK02lkerm
qG1ZDBDjiqT6MX+K7gbXbfy3fz+21e/C4b+4acKoWOfR7FQd6tEy1BLHvOqX7/wS
zwc3WQt9gmwwjnkzVwp0ut346FzUli25qYegtgivKENb+Z5GeV65+XlV2iiNv3/X
2K9YbmVyzrufPr5DstL5xlRullyE+axuPVvFgjqMgeYzRM7IWYpL6d+OI4NMsiVQ
/FYFWCOIFBMj5O+FJSZ5QNO2PrZ9Xy5mIt6CCEIr5mdIqaBQ5qPuLhbPXAtwstV0
`protect END_PROTECTED
