`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pDMXNQ/zENYfjEx86actP9tSRExbu76ifYEU+gEJ38IgZLm3yGTJa/f5Fe1qX0Un
Hq6gJ2e5V/G0gLBnlrX6fIN+S6bY+e2M3bAdXsVIFVeHMsLpgqOs02Xfap2PUlcH
LUN4bhR89Rjni1BI7rRpj/OqqrqgucsH5QimSdPjBQbm+ebdjhXjz5cqoqZJHSX2
/kmhasBaw8Q09JIWPHkyoVcSAbPumFW+LcQ8eeXjJkVKd7kgTKR3tmFh+TJt+Rw5
rAjhprPTFeqfVBxPChTYXHyAAm8PNQ97mzymNZF8zxhJFMBfLs66kW93iF8rr2oa
G8XU+jCoX333RxhW32OgGvrJu8qn0qc2mtNctEhyp0X9bd5Jy2305N9mfnXWnzuo
C7h+KuRY/AUvJMCkcZuSceB1BnqFVyGfqCMMT0nNNCkKvGv4IIup+8xtMsR4XstG
texoWh8uDlocACVpI+yqQUk9gNTRkTdEEa9nzdJ8YiJzk9y+VY+EJX0WyKBRBGji
yyh4zkuVshh+x1Mcj7E58ziGsoSf3vTCqCAEEgHtHY0WILDTnhljLxA2LpVHFHwL
ILTUC7ruxPxcZOLNq/VoFR6A53O1EEfWxuoHkqKzscD6ZeDSRwLZfklsBnNQomdP
v9yPZyYz4EVoEjNVTx6nCJTS74F6MevgjtvafXF55gBldQm5oSvYcDp3J1wxpwZk
H67plJIbx4gz+81tSoD8F1t4PXmnQihaTSGvT9hH5j0pc4Ex5C/Fx9IVg3MFk253
F1lvm5IJK7Mg5BxbKtETp+YWHOAd7sEm5tiXR3/tQYznyqWw/m0EdSteHqNfVLn4
pfboH7LW6CypIF/ycGLV63AxmEZTvkcSqo+L8xaa8QFNMDb5HgBa3GC/WD9MC16j
z05cXwaANpktiSIejPyFlpYyt8yPejsnjOTQyfMysKMNKcxORYwkeDQ8/IFEVVbc
0vbvwNSFl0pFYd3qRdjrKZ0y/cVxxwa5ufafv7dxClKFdbpcQEUH9DCWZXVDAc6N
/FTGrS7USrAstslvjFc6AgYZ+Si4UHXUGUPraLaVHIRE5/la/v6RERpN6zVPhaqw
`protect END_PROTECTED
