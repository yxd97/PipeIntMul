`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eWdd9bPHLYEb5CKhW+ItoCiHGo5+2+66bTdX9pKN+sldkHm7/tyvbxOFHW6lCjl
4WoilFyAXy8RtAy+Ussw0oBfSOozOY/pByZKHSvUTd/qzsfcwc418S7uHBe2qLy6
enFhfV/2Tests37CK08NQwmbqmTkvv8QEmF47S5utwPWCMdrcCxJ5nFr92rNgkCC
IzyxmjNhWDSJsoj13gLUdRgilLIWXFeVQ0hnRI0Bq0ioOQ01lgpc7P7htYBINDwC
UFYXjOh1X6IYuQztovWRDuFTkUSJyqwK8wbS2fXuon7kZPWvAbeV9Nps6QS+/86l
h1w+uFXDHdHU/jteXx0USu0mvga9HYBlZFN9Pyucjml7hy70IOsCxGBFRMKfD1l4
W/NyjlEnuljlT5IZ5N2kj8N4KCneu8CQFhaZBfX/vUEOCRW3eTX7MHG9uxvrqdM/
JwcnZmSBxxymd8lP3tDq6TFiVVNM5J1Vu+Wt8tYMlo0C+SPLMKsOflqWXSuBV7FO
GvVO8RD/dfS+cd1k5TobvrfuCJJifmAP9PikbuPVvUn5X9Quf5eBXvTetOXaDDXl
3xQKMMPZMTlg3cmME9srIKxt/qru1DP8uRdgu7lTWMSH1jx0WjTLi+vcYpOevmz4
T/pKDny/6D0snFqZeUqpKaQuL8m0MmJT5E40y7PP5e0PICEUw67gsqctrxEjx/PF
IIDCa0ISOR57AEKiM/kb897Z72Dmr2O5KNwtWuoWBjWVuuXNdwJuEOqH8HOYbZNQ
Wm3hlVrUz3P+0QbvF9Iza8Cn97fiSh/4Ce9hmrkab6zgBsBXYIAdJY9pNSGH4wmI
LQwghVsDOUfTHG/hDRyYVMOLucayiVJhPbgMwmmCGiykAW9uR2PLjidz07kczjO6
GW1o3eYCPLJHCf8QF8xZRJ3sRpgJHbAqrGO2bA7+TiiIbC9mmZDHRSy0KVDqKCcX
MPVef9sj5OLBhfSv/ssjdST7snRuZdUJzmzBC8TajXZNywKaBMnBGwRZ99ZWZkGA
9/C7P3DJwRiLABfcwHoKgI/7RSyvuGQe0GtlTQySwTiyaQYQQAni0vb9CcNs8byB
TvMP1xPu/AFOXLHEtvOBbdtLBEBin/at3cNzAzCr9uQgU2QnvPTYx7VxqgAFUvC+
ZSxvDyld/d/H+1Cw9dFzyvuaxf8OWIhHdPjsed+YDwVCLZPT06ldVM7co4pXQ35m
TeIuMCvz2rHI81PBiWnkxf4DkZnH9459FlveAJPYWK97CktwML+hcG7X+yViJ5ya
PGkbfouVsrPxdZ6yn+Hc4CvLHUCKp0SgDtRQ15Nva3NH/hFIFKgirP2Uy4n96nls
xx207UkjZTW7ELHzF8saBKH/RQ4nYh1VDNcvVahM14wsYVPWd495kI5C3kaxxiKn
KvmQn9ldJtV/jz6E61J1tlctsjOUxdRYW9EELr4VjCHRlYpKD6YRAADlRYC889LN
Zkd5n7xsdl9l1g9GR7gOlUNIXyMghRBL0r4xrlBqODmm8aDodGg9Ob2FAuarH9LG
qjEm/XUGIeRn9dCSZbkbOuwa6oMrNBJrm6CgxVH7f11TdMI5EH73scLQnNzqWrOV
y4dhRVL6pWSU6EKUvQROy4TpCvJ8JExseUAIBTstZNavIbYQYNmsC4aqj3NYhZI/
/uFvCm75hvfXwQpo+2K+jkS21DPBDVesVYbVinW1GxsuH7Ad8hRdMIcQO6sidoni
VH/Bk6/3fOS+yL7HSLcCOfnsJ3XAM13ZrNk8rzZFD0w8gRAUURmXHxOEiULP/ruI
rLuHY16hYBqTTa2hfhDVHjfzAzHnNHqAjnFZh2xKVI+KuuSNHfzSTmaLKgVMXKrd
OYHa7Dp34HeBTSsjisxrWaoMM3eJLjMaA2iKwAsUiOiqoJ5DBjFNU/a1/diUJbR6
NcJvUyuLfNkh/i1DTdKBX27F8k4tck0fegz2nrGhh+PTflskDx1sS2nd0knv44C8
BkgPmI/2IrHl2zpRxqB1FvWwib0nXdDix/qxxJjQ6VbEN7eGMIBrIKn7hoSUmfjO
l3HSWq4I+yn0HGPcHQRfE5ikHVURxbQ8Y/iWzzItTsVQlrZQrHwsImpRWBGKZHBv
GbG/tuUfKbLDCNHcZ+rD8Bv4ZwofP/z9acUWZQ1iG0TOlxMBKAk2bt2/T8jfkCDh
ZLH+w1+K1lHWzVWI6YnOsiIXAcRchwQAytVhMLH0Gv30SEpUaYQ0nEXaBvRF6A8S
Dk3+Onln7Ttl4w8M9ori7RWZMiLFtvQ6RH1MNyOM23LHXj7guAQlxINeVG1mokbc
nz1rssuCBshHYo69tXgUZ77fH4yNNWpSQvQJprzEteC/YTa7jtfb3akvAgbk/iHJ
ALkG68phI4d4fIAPeoJD4SWLBVJcsrKagONEoQebrHkJ2muQxiBzDPHsICf4tFdg
MmAYnqsPUtRgZi15xp+6Rk+Oj1Vi2hDGLZxTfY1aRfQTQoHjaenICGGAk32bPfkr
8wldsD3Wu+JWQchrtNHKWcFDVRC16r6YiPzyEwnnRS3ivGRslWVbSqLlJgE/Ie4y
bNyVKRw3LoOEXggdlv6HnnkWNtvPbpRMcqVrMCbhX6XOcJnst9BPjg5hxyQKU2A2
CU/nAEq2xAsGSXMQVfpcgG5OwkTbfIJq8B0ZTsWKZRjv/cYNh26/F9wTkW/1NoSI
+cu78hAYo8R/f/mz+LHJOy7jXKdsCnLjLzZ/PZvJ2QZ0bj0Jy3oYzcJzMRcmdz7f
Z0o0CWdpM7LWNIOT/+jB/EoOGrI7kHV19kiIvfGjPxe7F1XSgkwlENStL0I89DAc
9tcJfXMkC4YaTBPNyjdrcD2nRiO7Lo35kZ8LlqjYcn9LAbC02+gjSHlsZAvreuSS
MkTB2rG3iyngB8btadn9Ux1zIONmPHbTmRLpEuBw1asqxXfvMTHF3tf9rmfNdchK
4Gi3sRJWct6TqlFf6Dqso7duRL9Q/07rxlUvpgzhl5u70WkpaYf9QEdrWto/iT4A
nRcqCx45oTdQVcSHjjxd92jh9bRk4Vh6U/Siq4CCBO9I0POKJ7J+0CyXg/Tcn+ig
Rr0+jYm/C0JbaqP003ZGbiCnwo/fuzHmJaM2lXgM1x8knVNmK6myL2yzue37TnHC
PlWtVSfA5GxUBY4kb324bt2sxfwj7Gze1qho8RcPMdXoNVZz45OAvuxWGAQZmAr2
9ycs5b4QuwCs0sUwnLVGdZWUNL42tJP+3YJb1HLnD6av0YtOsRD41fFP2bEFe8Gm
C7qJLwdmngFln5JNp8VCbI0CXkL5sea4nU8xTVaAi7oXgNM4VsIxXt66c5xXX2c7
Ciwp2EiSkGSYsEtE37vqHjSLAhK1NSsNNrWGogIU5bT9rgpvtQZjcQvgBx2bZSmU
iaxJN0UtTLSs3ky2BPj/7Fhm6Fkht8hzDnwvIv3ceGHMAzWR/pHO1/aKGkthShmc
g3Zz3PtednVvcOP9Ez01fDykALxry+lTbvFZlJHQeL7lfwzdX+Pv2yye8H1APxjV
/J/UGxp20wMxbG+dvEix9Ml7kbhsBe7LfDxA6w8bpYAWWVkrIsdC/er1Upo6VAQi
E2v1MqoyhMRpC26omdZzyFb0qJAv+81gyDi8xARlwIjxhAT4RFA+XfLdCNIyd8F+
N4OA+2fcPfrme60ChMDdUkdhQcfq1yNxZSjM64Bp5DPCNCxIVszCKNleCB6eciA/
ePul0hnIzgFazpx0h4Xh6p6e9kb6Vy9UL8eIO3mY9DiOlevFqeSfEa2m6XX3S5xC
kE0h7UxBFBqfwZWTmzq0dPoUs+WLItBEJSKKjrMxg7oGK/OOuzI1z9jLXt6Jupav
VctJmH/XySW3XInwyuzAbklCTWag5LtFxkmcZSazQolf6PNDqsevNkpoc1k5klsI
r9mg7BPH66v3hCZtkP2szAtu/zRB48y1q74gk64gPHedrEsfkRQB/wTppya213On
HO/mNPAdPfXfPYauh2nWZO1t1mXH+MKUIbLGIsIPlB73JYevxqq7CFYszGIbYZGD
vb7aIZ39kf020lYm+lYNfQTGN9scRRVx9DrhLbrdcXnYqWBiSM6ooqVOedulCRtb
KpHFb8Bd3cGyudQk2W4GDl9HEAB0Kn7U0/8AlGMNNGy8i0xbJXbmwofQpkUpHYyN
NIIwYAgfyNt6IJMaeg+Z0Y5oN1Pum8twiv/dXNf5GOZp+XmPjmnqMJmKE8LkKJtx
FtRecGuTnPGREwErX35OIlw3ACzceH0p/000QX1xRB6RL16oQ3CJxnq/1p1bCKZW
t/qjmSA2lduwB0GFXfhtowXFOBadAdBQhKZnl/+eoZUhsGgfns/icFVwnqGvDsS4
BLo1VFFPXwRuE9u2VcMRlW1jX7Jbhdj2DR+y+6EOuAmsZclvHgd0MduLB2rXlrAr
EeZP50eu+nxBPvWvuPd3OQEP4M7oPLwfhIN6pHMW+FhEqsHMtffZp5oHNpe6AL85
VFEx6fCqx/jY1V4SPsCEkFyuGAoPnq0wEWMcC5J8wYL7MvoNmffukA1IAHu9Zns/
1EK9Gt8PN9I6x0VAnzqUeQsvmr236oNRrOPeInwe5pfuURp2tVjo4/OttOiHnWsv
mGtbFQ4GV4maoBdoFoGG1Cq1VPZRa8T4tHju2FjXLxCCrgWqry5QNG8ACvWdXdcH
hVTONmutU8Q1WeJdnTa0BSQHusmDSqhi0uEIS622ncobJsqBvIC+1QNHUR3TbvYp
bxJnvpuNeMyOvj7CZq6Imku8zwiyIrtpWa+8AxxcEmXnIjQqpkGpSEXMQcMWzsF5
vY+ms1yCECVJpkv06ko0QDLrgCUEFaQhBJgUrl/F94YpnFIiCs4NE8c84VSt9PLS
wsRc796TEtTloadC7Yf0yvSu+7wAQCmahgQr4ljTa8xyIUDpCMpmCrDvzlgI0e3X
FgoKlXUdiU9fNd1jX+koKrJ7II+5sPKEwHB+N9MwiGjNPTJ4VWKptZwKZKfj0jbZ
Ko7ZtUx9FnD5Ikp73OOTEOLx8kerVN9ypNo31bzhkbvWnkDUtHz9WqQeagc4ReTo
YmTCOiFi4IIfkVoFORSWLQnxOhODmtW7+17KwugYGmWp8NeAxr/mlSDF9Fk285aG
rSvvdL3RfRbWQajEME/i2X21jjSgygT2v3wn62pPNMDfw0M+RACAooJcgASJgwH6
eYhZk2vk8PTuDFgQewE89WBRM/OlljTdKRPEH5WazX9u37mnCU2ofOVHbIwCjEU7
1GOaFBn1NPABysbUcRMWXniJtdTNzMJF/2fwzL0oF4PL1Oo/RTjfDWHu7kXNwaK5
xfbkdGX+vFzrsXQQMYQKY+Lw09gKLTxMdsE0mfxLLq5DUuI19Iv7jrP8N/7K5DPy
DRgsVE9FwYVmAEo06hCSWjjpLMsHheO4FBarlHIcUMWWNoyt8KqxdT0FRbQ8/KiY
YwkklNIdG/AVedFO6s9/KsD8z2xQBj0cLuDDFz+oPzt1+EYs5+qgjrhOAR+qC8C7
FPBCxIK+4zSkycVWFajMTLNs50niU2znKTgNPF6/dM4dQrPDEBCJTo0DJ6LiSVQH
ZdfVvo8itOeQ4ePR6OF0hLwFTofqI8ek/KscCwTvUgk/tRg0aSAS5TQ065aV4KE6
MNlwWe7hCWGjBtp9uEVhhkE5i1DU0YnxSBgZo1wp+c32HKFN5reKuF4h89TJd1CV
H5vD0uEzgluDiEYUr9XhPR5+zswTtqECQr6h0FYwKKqjh54hRTXTyjYqZ5dThsi4
3soC0yixXadq/z4Eo4GV61ifo/XW+MuTb3GUAgiLpxswQByl8agOlOjZHO9nlerD
hmVOhlgLaTV+2/B3WGfC+LgD2xGO2Ku3sAxGYOeH/2vdKuPRj/jW8O6NPbY7vfR+
6O4QtREF6GPSD9CSPl/7Kek+AS3d6tR55GEG/ok5ONaPlFIJD3xXb0HUMTBxw8Lp
q120ldlyKvVgwCv/Bi2NLHnlEPPMQRCK0yd9xGGqiqYCvNyA7BhxsOAsauZeiZX3
cOsuD/+bpWk83R0pPkQ8liP6IptUsDEojIWvTzCtM/U7ibfqjG8JcLOU0Lbpy8at
P2XhepS58XX6qszZh0WChrmj+XRzhwZ57vDDInh8At56lio4pV7rveK5EqlpwvNe
CyeQd1MqxtRX+WAJYWhsHnyF/Pujp/TRia3UaAEiUUqy1WyvVrx6kVOvCG4Zuo6d
2H+Z9hoZx8/HCmJnrqGd/lIw+MCEZgJCKBewcGvyUo6YsV2ZzQ79DDJQfPxTSZpE
FQlESwFQR3wW7ZmQwbmAjPCLXlUnRGlKj7zK3s2Dxk9QOnpxPcKQahT+oVtTEQXc
m7hNnp8JALHgM/oQeFfPf1bz7/setsUZd1mVXEBiB2RkwTx0cRFbRIF1Kxm8RvRZ
S4jIj2qoWi99wrAYm0c2vkUKYevalpJT8TEF4eQMqR/oRvvlLmu3XGfUZvgh7XAu
qvCnmrY/QeYLq6VpMBD2mIbBdeo6xho4XQoTqH5WENfQOjttAmb6JAGCvfDgEZk9
Irvk0T3uV7TnkonB+9nCjnLYTtqI3loZgH6rvcWymyPXBBAc4/vqjd35jRs9jI5l
AlUwuatXd43mDfT5migJ4Xk0zXDLHCfwupTfe0D0s+jTCPvAaRXZHFh6jrYRMXF8
U7z1TWGkYoYHTnNH0q6DijcL4SRXSRT/6lS7xfJhjT9Hp5nn93Z3bSRUEjAtA7Ra
LmdbzXLO1tlJvchSu8BEh5ZdeJ/PWjuuCURW7+nBlnQB3kT5p5Wm48Zp5C0xLSZO
l9KzP1AasI3EtnZfX83w98VwW8tWruOBCWITLwTGZdHFtJRMaTWz3hEfNpZD8YNX
c3Jmq+4pRYJnOMJ/RCfWhCivCXzXvjaO0oztENjNWErwoWpIB6quu9wN8uS54vHj
hoBGgYNWyi2ms5sH4LUMbWH/5aYz416Iue7s0z6Sm932b/VNhqJMUxF4/cMU6pp+
B5QitzZ11npxepr44wwHJrapcAQSp7+a+rEMCcOzHwBW/SG+s9NAK5uzza1i7pTE
WGuU67yl+mu7TZkxx56iuacA7Uz6Z2Z+Fwwb7eItAb/ZwxJ18zDgvalk9VREqr8p
b0hrzrUiu6R9n9jxMsJOXxh18wJF9UK9vIM6q+Vt9AEIY/I8qQaYpa+z2DOAlYpx
jXLDz/YK+U47ogq2EI8EfHAPcYFG5qebsh6e1POw0N0A3Cb/YJ+eu7pxBhh7p19O
jMX+r86GbT9jQ/Ezo6p3vJWIJ0n5+AfuodbaVCwTWWMbp9k13kt6bSUfHoxVI51N
X4iIoDe2RE4tGxsMF3oHN5wzwSzEfWiHfApRCdljSW5bDFK9StAAhmQJZvc1I4dN
I35aRqyS2T6cQ115xwCcJG5ORnIM4t+zVGlRQVJZU8eAcePqVM00yfLPv8YeB49U
U5s26sH7PgYwkyaXH0z7t+f0hEWwun1nU730mrEu/1gg2KWGS64Tkx6qxvEsnVMW
+838dEwVZrsg1EZ9CfjOYJ0L/iZA86KuHPMHAInBu3z4TJqEISEyQXUjMwe3atEX
SDsDUMI2RudJRmsSdUS9KhSOKQsfGdaPJzULFPwKSDzDEAR/Niqf909iLzAPEOPx
V5q6SZDOaPergbo2Bkwtoyw6eRJCIe6PuKnvQLigUpzWDSKS6p6iDHyBrC5MT2jU
nm6TSD7QiP4kscsJzNITjw7oUdSYl4zQ9cbwZEwYYMgqCDGBiMZzDgWj2FICPYV0
AErxSnf+ZH/fBL9vlbu1kKJtxXfYwdURjGjsZwz/Nw+CAnjFXZOQN6OGFq+iP2Ve
ZCd2Jpb+QzgDNVPjQkEh52fWoWefp7t3A5W0WGyvKd/iqnN2nwjXcyQ/7aXh7V83
ujohF7jB4j9RiTVocTtRwJMjTQ8dAHmTLpzfoC5eeaDBuDWrlsYdUEHZGQ1/LlUg
XI5dmfNp+2hJAQuiHW0ctHQjcNoKFGdj40iCXH0DK0qn33yN/x6YbHq7/O8Pgw8v
UgP4KUyztxpYEStOEsxsMHzzPC/VEiBR8tEkvG1sffyAE+YJKpU0B41WnmVijoGN
IIdLP+Tfp3KPsqzG7SDg3w/Srd7deb2yAXAcewCUNyHPfrTKr2qpwiS59m11crJD
rpi5Raeu+1llitTI/H5L+1Da9l2U3Cd4Rj/03dS36l1mIO+AUvcgRNMg8GiGAQK8
A3QatapjurUFEHP7W2biK01y8xg7/lQ/F6fCvtsY5NzOtXWO3k3H1KuMbQXbhRAf
5PcOq7Kd+ffE4IzD7egR3GKkHZrq+dnYJDtFEOMMr+vQ9em0CbV8XOTSaOlGYYsi
eBPqpY0z+kdA8kYFu+SkPD0fb/lvf/HHS67yA28L/tgP712skk7EZwwPW5J1QipO
88S8OOilKJbgolIg5aFgmJd7xO23JEu2nlBBqkfGnpFcdBIuF0+u8J9CycmP/3y9
EATuuyxqLzw5ZRvgHd7N1lDgtlZSazOWwpdfretYsFOvOjq4zahRCDZdws1BYHSQ
QXpqtHzf83l2Yj0L0hq22lp6X7HNyFV0i1dMPKFVFopn6F6T/BQjsjm9+ZE9OL1u
anBtScwzGL2CUBCIbBJYL0tlLAOUNeLu3n7UGtK6zeyUjfJbKIHBX+JPSB4IbI6m
ottIXGKtRVUmK+h5ezoOEIlVFNUlAfYcdIMidtZcY7nPgkQ2Gloveunygz755v/z
SZsnwzqK4X8sKyjuL3lMF8S8kR7dpswvfNdfF3OOBw9yQhmU0RhsAAOYKXuNr66l
hk+5TegKfqmAkGvG3yKHAIoQMt/SofdxX9BVI+whKW8ktKuVbTOBpb8ogT/2Nexj
YOeUZzMRPIe848y+Q1B4+4M8xYikgXZglrZTAaqieDG/gPHPs7cSpSrP7erIwBFF
HLyX2SF64FkpPho9LuPxfMxB96FzKYJmH1UmF5G6TiHTC5iMlf/EfbWj6yFC5gnJ
4zrRL9y+EXd2IdzKlnODVB+4cVEbKgm6fwOn9x/QMjAVs27DNRvY5zjzjr8fD6Yz
ukq46G6ULE2lwceU4OR1bz+9we9Q2qx81ac8vF8giOBwIBKf1ZT3VSYFpnCeDNTZ
hhkpY4TM2Z8O9ElgtdpC33YLZjCYIl9NCihowtycGvCtSdobm01Be4UT8EPSMl/s
CWJp2YoP/QPlkvKikcGkrqJEpfy67A0yKF5sCcvUZuJONQq+R6fQRjnXe1hGveAY
SbLVpAVhux/qt5K1i4GZnA4CT2Axj6qA6U5Hzg9HABnCscdNMceSKnQClMdcwxom
PK+GE6whHcpy1VyopSk8bfnyTHOy5hOzLJJ2bfd7xA04zPlSnpyFEjuMe+SBpv/k
2YPaVD1XHvSmuMM+m4X20IQptA/VwFTkyp9dzjNJtvgheqFYMv7FYZ0N9nsx95SM
G3xMQxDXiDEBv6G3dl/84cOe2PuuLbMPjQCgIidnXexapyUX85bLk8dOCeSpYKLz
N5JX32qxAWR4nlLRXWWA9E+Cb78V2fi+lL5BZbteBNozddGQRbjRJfSkDbr1hJn0
i4uqtmQcZGaa6EX/qHRz1xzXKxlKGt6iulN9+VaD7WUtmCC5UmUHkqQuQ0dh9s2M
iQrzAy8rBZReTs+jCiSGr3o3h3RQPlgO4PtnlhlBNPME9aTeWcGz0Ry+LLDmzywS
CU+p0/dDYOmEJ8V2ASoUdo6GdgtuxhDokvkqYC08rGDMgxjWsX+ks3i6IXULUCa9
MM+TMc1AmAypMaTOYf07PIvcxD5Rwz1vSaYJmGCWELfFiHjhBOk3MGHYFYPklScT
lWeb7/a8//bvl+uCUvwsp1ry9Q1mZbDT2ISmqU7XduoIfkH1PQ9L8AzzKgLIKm8v
g3i45KdxnB60GxpkSTuo9edVKwXc8Ml9CCxPXXBLkj9NYTRsKbPGu2df/kVDV4XS
bj75xD2cwxdjfh0TOuBHsk/J+Y8MQB47lCAMiB5JfQFq7KDwU88sW2Pjm6WHUXkD
QC7HZOPgcEj8ToIKKgVHYNmoBlJkNA7bbIo2zL6vC3OJRZ+kCgoAsLyOGOYpn/en
g88RWDsZD9bTQwRtaroV1P+rhYmBiqgOhJaRRkArHjg+py/BDKvX/QqobAN4FVCh
NK+4lus5d8Aobh/xxPFt5iBXj90ILiBXABQZzrFhbAIfvvBC0qQFi61VeXSHjgB7
ZKV/TXKHYGHZGmTINbwBWATkrt5yRdQW+kTMGuJiXaYajD3l3rydLp5J2juUPlKo
CJOqxmroevpQf4G8BTYOg32lUTILJdlNhlBva+xiKzBNoUlR1o3jnnRVsL/Eup5U
9jCg0/WsgTZWxcXlW4CL909ClOJNng0obYNo2ITVD9JXo6xaDln4qA9mBPWEpQwC
mvEvz/DOfZudIEOZkb8fcqDvY8ic50ELEPpdQ/sg65EtYZaqthzwZaolU/YorW+t
pDUlvq+mD0ROGbAJsahlGcM3KQDLMUVVm7caJlvyh1Ew1ea2fRuiPOVdlEMabt1A
Hf/2z418aZp3g9E+vz2MXTsRfY6IaPHBAXlXpsz+woCxz8qjz7c1s2OEhPog+1tN
I10+80qtwldfDPPsFHQa8i6dpEBZ6s/rQz4gCUnQaa8KSop5Jk1QGzKQy13UOQcn
wOBdyTNsqfoa+3XSp5OMTBDBvbw5RcWReia81f/4Lt1NyhxfTi6wi95v1G8NLHmU
46p/lZOWkmrkadlYkH+2zLIkaIBECKbXJMOsyQI/br6MNaMLEHQ92DMQsBXfRGMt
CnzFjbmKBkLEfh9fgbQrOzOGppGcS3XdW7NeLmKuc2mp8a43mMRiv8sJ8Q7Shrs4
P46dOv9rUBAhq0kRP7hSt7v5kRlSlCwBOSMhTo+yejfxzS44I/MyP49pZARVNhCR
axDKy+3jSWy9++ujOi4wL2e8q91M7nQGVzV+ZWAl3QrWcEpqRyS5f8m5BSRTh8E6
JumYvAh7+COypE0nIGGYlymwS5IAhEEJap/X5tnZaxPLkoyVF+D+RX4axrJn2mDb
mreX7JCZtV1FztJNWXwsksAbx1mWNhJUryCPhThIFuXNvD5XOMfxKsn1lheWlPAC
BkhsWFs3QAa7xpUNoI9lqgqeaefl8y8XnG8CL6zWv6UMQi6X1Gf6VxMI/OQnUO5p
obaGOHXmB4aLSYcyoJVR/dm7yZ8+iCWqd4JtombWDkJIJwswi8pEv4c948FjQblT
9sqrbsIlS/IknXreSghhPJi7pbqvrUu41cG2oK8iHzb4eXASvPQ9MrBXqUoMizny
LGVmGV3KHS+1P+nof5DG3OMD76Fd7k10bGwIFApoeaKNjTCwKpotnt+hfQvVrol2
tEKNyCWkdgOCq5Rz3fW9QQ0CVWQN9SsebYHLQLV/0SOVKgjexdL/2J4O44KziHRk
MizIu7XgTMhmm5r3ZjBl2wSOLxjc07Jfur2IqUkNjzUPj3j7chHxU3LFeNNCQntq
Ib7fDQjtD676q6fXi2jKqG0/ohwJtJWO8aDmjHDkfIUN5+qFpV4SDT26Pu8Bz3jq
h9CY/p9DdSShjD5JkUyDBLCPgf8wgnA/CtvCvRd61/WXU4dNlNDsEZMgGrQzc4Wi
EfSNktIBt/Mj9Es9AufmeTJnESiGrF0P8LQ8YTcSO2iW5dwlVWt4Qjps+RKreumd
ZxYnO4Q/B+JGA4qpkiwZtD92Sj847b/OzTnAqnKmwb7E002V2ayIWHRCTa2GmZuh
vFZ+aKqU7IsAIXlaTJCXrOGmfDCqqpdfIc07Z93VgJn2WCBS4bDOEaKfkK5xJhsB
C23M8ThAmsTzqd8+9KE5oUyMpYKJ8NoBdUaWZ2jj25qHaa0X4BQnvCOdWgFoPLAy
CUuDMiJBBK3ao/UnVQTfEWUH4xiXEiLau60eT/pSt/S/LFQXqP2R2pPPz4hcOvrq
sm51Gcz62wo4WG6wGw1PHa9/X7JeE99+P9OGm8HvN5INnEWfUXUX4IRonwhJGnbj
dYLTma+rfKuWo33T3+kGym9DOkrC9WUkBcjNEaXuJWSnVK/GFDdEEMV8a/TmDqU4
MvnYWy6hFGr0TaN+c5RowefFOM6M5CsMkIbIY744WA82BGOvfqZBJxzapcGgPAjM
DTfAu3isu9W0ylhT2562M/sXVJZq0IUZIzmSogMqAtAM2Eca1xMCnAHCFX7ToUze
lQLp0z687vuSl2e7qmq3+ejuxuCLKcnHv+a50eNbdOW2vZa1tUtKu+K2SuPxpnyv
QUapg5zIVVwaC5INedvKdlB5Rw6Ns8ssChLd3t3YlhKrOJuCb5awb6z3seIss56Y
7UcUDXo6N5RnLYlQNbC6ofLBW/NpitGUG0OOLxIrL1H3nZQAW3qX6AFQC91TRSZT
bCE5BkOi4kTsRQojfwtnvmT8GTbqIlZshE/y6vm/GCTdpImnO6jKaMHgcr4eR+yy
LPfq1NtI+uPXSidvlyYBIw1Or3Nmj1TcQE+ynl4WSocCi0FVzJRwp8+o+BKlAWV+
+QmtCIDfClPgnhac9DgUVqd6FQz/R2rh1l346kGucbI2QNTqurS78mZFO7CTyZq1
W6xpECkGWsLIBcuGwnrYzsSQQZT6iomKlRLjexqmlz7Uoo+4or70SAeOa7ms4ttZ
SIsHkRmzZ4mbyrPzX9fRZFIBRbu5vts+4i0Lk6ZWT2+Qg/M7BAtzH5hqZYCnsiQQ
F51wbnZ5yGK19GbmSmnVGJ9FVsVqUbnJNYzzojVONDlHm6TX2D9T7MJ5/aFLBU4l
dM7UzT4jjUCRBtxZAY4cBPZ7ku7dPInSftnT90OOhqxpH32dROyOAZ7QqPnk9XUD
3O9KE6PKovTAkKZ+WyP2cJsEfGyimdKU5lGTbfLppC9yizqXFWUXDEx+IswjQaF0
yCHmxUXGk7bZNOfVTsRcu3Dka2J+af9f9arnlCFTHqG4RK1oMAOe4Pn2rzGVZVvr
+zDl3pR/DCofJm79dA+5DtBjV/I3UzJnfZDDfq85CTrMviEQ9qhHoGrR6BSlTC6E
Xl0VJHubhg1U29IyX6EDHZTMPmk7pCnaPL6sffb/CsSMdVPV8sOGwVb49Q94xpQw
wk/gTtnYvi4WV/Q02d8yf5CiAPEhkk8vkCz0+Bym0TjG5ZXp36v41FDJrnGr+iWy
dcsR9HhHBlb1sDzDYC+9+vaiGuRbTva7Ep/6pJZEQcXBUrNnvKa88f9Zaf0DcJ29
yXyfrS6EIXov7b0c43Yh+KR93zCHsDS/sTeJ24kAJPEBplA9irOU8+FNt/xpDv2F
It61PyFBoJ/2v9a9GYOdEd0OXeD7e8+aL9dUZA78zkM3VbMXaVprYNkFbV8zYcLo
ckaZRSaA+R4B56picf6KMrk8l5WjOTlBLmi4hI9H0VsqKjSgW7o/Q/GVhgIfiQlx
iIlqHUYYcHK0syM9W5HeKGUrjJSDSy8RoWvWmLxiXsB85M+q2B+bKRIUxyQKnQOW
nHpA8pRVylVcwfyDvWIM/oruaXRlDuHLQc2aR8ZYN0UPr6+mt8OQ9SINVP89s1T4
U13DxvI35NyrYWqZZ9e9eDx+M7EZRFsdJnx5oMFYbdNHw2CYZ+ogejw1ME1q8ozI
bJM2MBeFVmPH/dwiIBXsneRXhYBy9PpPyuH6KkyR1wIqcTgSfkyIVEHvS94JjCWg
p2q9FuOoozck+j6GCNg5wdj2FTfCq9DyZoJyuSJxT+3Qo9fqayMqB7f845RPcSBW
/xq7l5m4vFghtkvTSaIPzECqHUd99C8eiXxAyFPBFUBYs2DnF69TpgSEIK3vP/uy
RvgMvd9zNuvuTK7EsB7h2238xzhNacNPL4h64d087Kg7Mo4j7q8jiF09aPw3sPSx
hR2+GF9G7FYReLzm2mWm2QfinzmAmISmi+1sSVHi8YxDyLGvVrBGjNE3Q9JFuQKB
MdsXsPTSETT+iMHVdAZbaFMFu+qgPUPkErz99bTho6iNo/mMdmp4Xd37wctQFBIQ
MosfeGw5he/Eq0+OhkBGu42iqtaGy5S4gZSTezyT+dyrPC5CPpinVmDKun/g2nJ1
kFavgeXTxOPf8oOpGTiSFf3NjthAslIvgR9BP9uX3KEZRWB3cyNsrcnhc2BMXZMP
3tygqMMIJfMfa+n3oxSOkNrFwxsaz1noQXVC6/chY1vjvOYUMJKcqToy5elaDy4G
6ZZ6HJiaLdKkCi0/Ow3aeeR0zG7ZTIyXWOXNJpcPaONrJcyOC4K7UK56/KsopIWR
N/or8Ro94kOBaXZhIwNC9/bnEKlPKMIZ5QqMENXuVoJNMUypWG2gq193Ny/FKiY5
8OZIiHL8DjMaBHcQnSPM9gd4kyvooeMl7lVzBlMvkhD2YhcxDfgNAX6DFMxaKPM4
7nLJsy+Yq3ZYZNpknbCXJqJNHJJ36/mXPRBNIjquB9DS245DiINwJfdPaZ43NAPA
CdDO0/oerIkXKW92h/ap/A09GDzDV/pKLhcV/d5V1pbkZAM3sASYjgjxbqGi62Uw
FL6bRFnrKk7fWkVpOmEATic3WtofIM4rexKQC9v6OLH3ZBZ5HG0WgDg6G2pKRJcr
5UjvgnCr0ArxlSqtKzmND4BB1fy59wzD56U6fyeE8f5ZdRd+LHLrT0hZAc8Mq2FK
mr/fkNS9PC0kOz9wuIWFPhsM0ELpEK5fyYr8PfNjKj/+JJwpTW/G7ezpkA8sWatl
BXFhDTaEZ7bKXw5PG+xEdA1J8ZQbKx+I8bs46keeKLZmT+5pX4CeZS8KhA/zRTSj
5btwbyJG1JBW1mdm1jauFzpS9S9B2nP0v+59qYM1uyAzOUamNntcs1rNBlvmT333
d6piTLC7iipWXX++dQfCwlP3Vi22VZwd9tEkWQ1e/qQYRf3bgqWLTzs8NE5ZUMvW
09wLi7+9NwYIOI+m9/JvEjZRJdmJWvgj8xUf1joAKzLtjtr0HwbafMJERvrpr1yb
GyVjtyrAP+IUdlWYMl3HzcRcQSeUFDxRj/hzr8MNbmCZQgoPKgH9bPqSnHH/FHHW
FmPN2jb3Qd+F2MiOfdxXH1IXp2wiIIz5SYxgfy1MQDlcDqgpm+DKGAx7ceLA6yGv
q1LbKya9DAZ6LVhhFklW02BYR9987B3NMVLIfzmrKxrnJtdM06AYyjJnTjvy/nc2
x+SNFu/QDTHF6FHsBJoCZxRnr371t4fnNYs0StaXpRc2ufszWhsM2GnE8wwRzr6C
F9WaCzdYxahRhvM43AqpPLGmBeGz3nH61gmqoqdWF6uq3JuhvMt826KVR1b4slUr
MaLDNn5QexOEGnPbmsM4IAY0IApMfIv336ZH0JXC2Jutc2nyeF0GN+7quN1C0y3a
8NiSt3Q1MCjQqfL/WCbcYbDGuMbX5cJoDuE3HasZCIOczEuwieRixq7WLseXyJD8
pmuGoVp2nxCzaiSCRg5I+OJT+8+AxyvtMDKy+eMKJUsqtABXZDtzia7lBGZ+6Uxf
b99eSVFkJNaE05aS/AlspC5rkEHvM9mu0mtX621jrmoyBMdWdItdnHQck9ZTIIls
AysFk/PW0yBea5KCHpt9Gb9skh14BXVIp2CiSfcHT8mKja6zEyqXBeh8C2U/H0uu
zDxd4pQmM0IbPZ8i4lrkatrA3bUW5SIMdHoeXnvtHFVKNZmxh2cQ25MP+pi0hF1A
N5tUUoFJDf88VeSdn17F2SDO9e7AoeUWIZb7xQME2Jp6SDcHy93pFxCgPhdFHHxS
BwN3x74VYKovQAnJZNqn8mqn8wYMEcwFsVtC4YXTD9xXp9/vrBhB034jTdLSj8bj
iT1Tx4Qs4sAGDPFMk0oq+yG1sLollGIDB6Fs82HF3WYLjQ+8eGTx19oOsleR2ole
GXI7+8ww+dzrHK9HBk5nYNc63UB2w4ohYamgfDhnq7cpVdHZb7Jyah+wnO6W2uF9
0V3xe9JdHpWLXlADA9XhUl5U9DrcI7YHerND/5aMmgXC2Y82epsU+0Cz3eVmnd/P
StWNn80NF0GQAtOICG2kquO6AXSmXr+5Op2G5VMwJy7ZtwUmL3DV9DxKyy3ToQ/h
fXH/xqPwxTawlIbo6UsVvA5Vweo0D6zDe1eFQSGZMCUKF2N+jO8HqXfnEFtl/jgM
zqzNB9TyJeFboTdbXJT93kJ5TGvotfQy4rSbkogOvCaJSdpffge83YZbjrhgan6+
YQGmCMpu5bmPDr/XMquVsosBgqX1TxUO7AReFFlS/emK3AFKpaRDSzIB/istho38
wSX0BpLfgwjfFv9DLCjhqikC52YSpVWRSsb1cdI9azGWWJulhdY8lJfuclQ7/uHO
MhpX++5YSSMfjqCLa6I8mPUKEsRrDicgSMwyOJXLDBiWmeUTDN/SX7niFJRuKDqx
cQQxJYV1zT24d5ZmeO4RXUjdwI4KqWyMU+4xRGh6/W048jKErCH9+12iv0po5eV3
MQqHiDTluyd49qXdA614UY0tCW9itzK8+n+gEao8ZQRU1Y/JIttHWknqwcXwtS2R
xJ0sP1Ix49xTOFDLXWD6+Fe4KI4bt8hnR1XdOT64lv4j6sguTa1asVhY9ohVED8o
KKK7ID1RHvRJ2spwHehrqEDHtmPYa4zgBAthJNB0zvcd2x+9BdIrKKFgx2LKaCkG
Czheyf0J+b3SBLt9/KDgnEEii855ASJlflwRD/+lda6kVsegolWUoel2+4ec+tG8
Kw+nQKSbaYIyCLjrxDAPXVmo/+1bHr+PeRTj/kb3v5Bzw0nLQnIuzkMjR6nBLmNy
wNiNC/2KEZWimmEZalRWcRyBJ/eIHWdGspCGswELNT3+K1YtoH8ArQsOgcmqdseF
v+dTHfqmHBFTk+n6HWm2W1fn5z0ZuawzNn9TLFXv9nbqpnJb7bYxO7QGcahMa4MI
N79BXuAM30Alb4jMJvrNdVhbJC5ii/wDwPBYcckeaiT7bAP+P+MQUrhP6GRO0S/8
coOOQGPaqCxbHsEdZHLGY5VahPZweLpYeMar+qDxCETv3TZjUmADF5HgtLctZlMC
lsfoRRkhpFSRwI6C4nE6/z2Y6HPtb4YIeDwVctFENRR0OY7gqjWqu9qkV31OCGgK
v3jG0SFUcEsCnb+oC2R07gHv42OadKypByShp4dzTaynE+lYRnikZZfWQ745EP9q
qsqHbsBqBdLTj1bzfrn3+nhb/rmqNZ8XYPpraS/11a/NFEa5eGvOEWX9hews0y+M
QCIQVfsRuq9fT2xWgwM1PzVWQ8Y5TQIHWhX/KbMCJTZwB9jmiu+a5Ata+a/gg8mF
Yj8NFMN1QZj0Q/LIhaSIvwD+SmpG2v6oKwwG/MtsR9Lln2OzOTNQYDc0TbI8oznL
TpngUIvZC0NNZF4eEbhOWhUNooTsroRYneobt53zLLUSiB9/gZi3mB+dg5LO0b7b
CCd+z4QX1q6UFtv8/ccQ7x1N+3jqDUTxb9jY1xQSiUSuMqN2hJRPj0hcduRy7/TX
Ah0MtlJvog08KkDvPvH5DvmdJwCtn69xKTRx8RjjKD1V9HgCDr0ERrJF6D+EPzok
3PSCKBZONecUbVu6nD7I0xi7GEDbcbwCq2M79WR9bdpTvREodimbPaYDgq9Fci1z
2jAtUMs6o0XqEiGAif8/+6GfVL57HywVb3IjWIdLhI7RxT+8oo1nF7Xx7OLhaaRQ
wzsJ6usEh/A437zilvxb3eEqIpEUvW7bPq7i2KuhfiIi8TjD7lNMHcqCuXUQdqRh
JlYNeCMqxMavJ+D15fuYz/3Uh02efbKn5SpaFW1+Rp26FTAItIIBrTKIIHYimimE
JEdSHaWlzrRR98sEZrGAtexI2PRHqIwifeldnorqHdlEn2UuSpmMU4JAFqE9N/Dn
xRO/xSvaYjli8LRJVPsC5JnIveRE0HdNInzXy2uu0k8G0HJburu0kxlnhyz6F13t
zk5nEGaWLv7n6WgYKN4w9owbRwvrqxs5sOAwegNYKmQskmCcdIIltJ/j48p1UXgl
bITByuxlsb+lNv5MdHCBYAcb6a0awxncjJbpF66tz2olj6g3KocgJSOFKHl46Bic
8ewnWALKeQkegTW+5ELkuYoAUtHVVZtd4MXfRts2OLonDjuHXuhhsrbooeXP4Lq9
6g/paa2VclSFShlq1Fs3FKvWJ5xlXlbr++jPspyeKel05ulySKL7u1/j7AkTT4dG
2zAkGwJpCLtcZrk0Vsa4mMWl7wSvdPKGmpzNdxoLUslHt/DpWWKgTn3sRdNn6d07
M+UP3qcjYpRh54YrdR1Jn7oVdnBc0pwnQN5WMzuKw/fRaAQU575f4SOfsjgbU64o
zj+IZZzXaIno98I8QalC5X6rn2y039eq1XFl1dGcBE7VKGrOZgw9RYcODTSyTV5F
/zmemUvfwhBlRpJAdoauScpeTgP09TuvQk1dYqIy0hhH3ID1UgR6kKu1NwXBc8/A
EkdLogF/aMSG+D09/56vxsWHpj+os8a4ysR1lSwtPpFU5iG+W6fXb5nK7AkhvLgY
p9dQ1U6NfyKjQV14C32IgGaJtomULGkXxCaS6xhN1yMRuhvpwI7kLNG2i33naeA4
fW28M6vUTo36Rxeh9Bp/5xmwiCwLn/0X63CUPm+ua/Zn+5AnLYF+1zxP4tZ4LUTQ
/1RnRm+7KuFLOUUu0X8u24Fhjs16gZHIxrjR01RPVyZH0REht8XLZeOze6vYIyvJ
512kHMvZJ4ZG5DeWNc+tAz1sEeM+3Z+E/lmafgaD000An6tYYorb3LgDfjKUfMgw
B6WW76VtAu7MEVec7VaJBzwc0Z3h4bBzyjJxAz+a4+iogRJtFPVvVm8XFVCprKFr
O5SL/OI5nZfwNAFIa+oPrZnlg1gSWlCSNMciXM7MfLzDYFCfmXSEavGBQQwHaRhU
5pYnH/MY+2GKAardM76uWY59E4rCakBeI0D/54Xl5y7FOj/htgKQA+1zQto/SiZU
dwbAI770+oJ82fR2kxcA0+nFYy1COTxqCvcZfpRvv8W+8ALOx3apfjThWtCvvyTS
bt0B9ZCJp/aF6UuA1H7wtuCq3HexxYVhvsHI3VsDQvLteP38xC+A6uQSRf3t4p/a
GXfELw989kuYND+9OzKUzCyUeRiMq1IRv1r/kln4ZARJklrxkgocbAd2Uk0WyODm
AsLnueAUDH5dpdsF9/XiV7xYgX8Z5s3xHxjFnu8OpJrAcgW1By/KlFDRBM2qkNiO
6nVrjA/au0c0vt3y5zLdNKp1t7R1r0svD6O1P4XIDj67psthyWdbASqYMfEuOxMt
vwdVJUeUs68cv1L9B+CiSAK+jDJ57TF8Ukd5Y7WvLW4fu1+FD5eoGcArUTsjWrvq
sOgBGUdv1ldu1UourBza3rYYyVCvt4bgwHCYSBbLrENKCzuVcBW3SCR31/hK8zyS
4AuhM2u8lBXGDJaC1ENrgVxxXbi/kQgHIw+FJK2rPEMHwUFE6JaFlGAbLO5kgknT
pw0YynWIkJNpq2VW93Stro73zq2nmboOa3EC0i5vRYKmeR9SaPpTZnn+FOuAA2a6
qWvCrPCDjKeP5N2lHzDaYPx6CmU/lsLIoOY4DX5gcqSqFugItTYntQLZyrDl/jBD
ljjwe8Vk8Ktc35ueMLWZNkz/Hq6sLuEPICI7Oz/HeQCjAbbM9Wl3l0wjBvhvOFwW
D6SJOO/ZGXquHlhyaCUdhGWfrhAjQAMRya0cFe1cXms5bhbwc5wQBmgzh1PczarB
Lkd7lxnfsAR8WtaPJS1Jg3oi+D1tnMm6f+z1fGWY6rhE6up4KkV4FDDruGsKdHhk
ldWrUpMCelesjVOi+NSK21H4yqmlDc9Iu0kqzvR33Ok5o4sU7CT7+TdUb6KB1YeP
ZfHZm+1rHdSydfRbX/UAsXC26TQ9MhRn2JZh8ESJkbFxb9jHwOf+wp8+vzdI3RH/
sgHyxo9UYfScGG9hmZAkf/FuFYRn5Hz2Q57Kt3/d5iFmZEdMKukbrHyRQctUoQ06
Kyigsb/0qZjsNvrxqYuSsob7xTLWEPUaeXzX/XCCDJ/qMLFnW8KFKhPddH9GvhwO
9rBuhlsDVI5s+RuTMhhTKWvMqiSPI/yynz190Urvn9maA/vsxHz1OxnF4Ez9gmkb
CS5xrAPWuX5pG8Rg25wPx5vD9WEDp6g8amE4JOdwyFII8FPGkEUsmmoj3/8qhGl5
aGPukOpq/oeFg9gWUpgpvaSCyEl23YKal2Yv0dV9DOY81jWqS9sAuyITTLG4TP7b
AAJ9iiXNf9HgWwYUCQUJTEXQjqAPyCLxd2ICJfHpAmq4rfDBgMJb8Y8grpmsKyr2
HqDgTG/bB9lHptdhxc0M264O2ACuTJlMbtqGQkFVYLZ8qdE+wLS/NF7lXCPQvWIk
EY7fCjvqIubVkqxuC3UDeAiCljEOnq0ipaQNdEop3g5tjkow47u5e0h3xiSfu6M4
K3YwCjxQgppvpbPkp2BgjHddsEhE+N/AohW1GOiqoABOUHMYZiOXAoeSzMq008j6
Cw34J/+nl4Dr6goQL2ZFfYDKSririAJI4AqDsC1+Y3D2I+3cjX0iamabYgystTJM
Rg9ZDuSzFQQ5LoOyxc3rrRxrFTWtwypBaIvf4Fp7dfby89c6U0Vqu+EBofECVH6U
XwPyNL7yIi8THBANml6gfbt+ot1iHtDj50NZUXVkBhNTTYp55pHK+ufjwkjTpScl
gAhMmegsLQjoqtRtrUBCmBWLQsf8OoTz2GyG6PhjnG7+cXrtRggWQI30vf4U6+he
LfEwjgqc6sUcC5eOpKwwK+TzGyWfMsP52VdpIi6WaCy24t3v9LDR6zWlzk6u+63l
V2OvTO6GuMVcYNp2v0DUMCZ1nXgcSuzs9+pHSoLslXPqUXbqSh03B3AwcTF0DcZG
8KwvuNQfvxiW7VKapVq9rE6wUPoDG68mbLNHqtqbHqgnXcoVhPaA5ESDeANb6mep
kBpm4KCB65OF9lyRV4u6u6kxViSK10Eyhdc3Q88cRe40X1nG0kZi3pqR/XyviXFC
QJEFZcVCAzn6rmTYWrOPWmxoY5S4aXwxTC/J9VeOgYCzRDBNkgi6W8o8xa7+ErBm
bIHdO+Fru7gPCv90E34AneFOkifJqu4RlUuNV5c+x84EqUFOqiJPg6NQuy4pOLQl
RKyMl/NDhFgKwtnUEGqAaoTGWj5+wG0vfAExCyUHH/X1Wt+CeFh6Ibp4lNn5Yt14
CWm+Xde979AygzTlW8092eQ+XnFChJg0YlJcb9Vg5oMVjzLrkz61lXATNaw07nBG
QtpZo1Xv74PacKzuQ9ANPPbYSXbR2I/oaomf3m1JyYDElic7hgxnInFqK62IS2dK
LAgsBzgPoH037vtPsOgxDxMbxsdrsvQkiUo5Uv+YDEfbHX6XzkDHr42ByNLUl63x
t/G7E9eozn7s87U/eP0NvMTM5vUJFREzzLjbF8RpJjDOF0yNyUTL5ZUSiPAffpCD
AJxvDGQk78fJ79VK5Yq1rZ174cyKUiSP922O8HiMWXIaC3jEKBxMT7V8d6zp+ucp
0HuV11Kfgiu1XgIDwwhZT9rAi73rL4exyBHL9TaQhAk1xAkzOyxiwjaTKoT8JgwP
+gOEQ91rDorXDlbUP6moU+Da9VFlZW58KTlBHsuFoKDkqOph1qkEQZv94icByyIl
jxZXLxwpKMhbZLteaeBT70H7H2Bd59BCS7B+8aTdpbFyheU0m+frY6uvRd+sxuuu
UoWQu+CK25sS25g9dWLcM9CWZ2EjFA2o1x9oBqS++JhVjjgFS9BuwFL+4n7v24pb
6QTH8lIaTMk55NgumcU9+qZiN9ePvYmBhjEShfuCp9aTMhP7x0v/QSoHsRyOLQ7A
ayANyFkW2T1M/9lWRocy+nT4He8Ymoz265gQm4iAlqgIpdpx1KB0OLL6CglnAcd9
HPijuwQBrMzVbXDo4inp7gFNj7narZxqqgXejLtB6US/72PD9qruXfRvGkOpmYHh
2WlRj6lQhg/n1nLW5wS39gbVCjOapsTY3XFwR2bWJdZq6EGCgkN2SovHWwikwYA8
gbcEmOIPcD+LYO1AaJcdWBiF1TAw//N4hzL47WEUOIxXT3am+bmi6j1hRBCBa2Nt
6iFa9Jj1JdM0Y5AGGje+ZTPbuookXNXCGCIn0YJLxcPdLEH3A9E/OQnbRIeJTrI4
st08Pg3KZckaT3l4ApUasTTHPvuMVeD9svkUqfAtlwy8D6sMHzKZe/KeyW6g9w0Z
qVr5E7EGl5OrhW8iuD419HQt5yh6UN/SK7tPE5kPDETU9iENj5wZuHWNfDROVaJj
CkE0goWYRfKcVJwJc6Vw7AYudy+ST90pw/bHB7+JYrUtOom9Y1b5qcCwTEDGSBJa
Fb9tVqjIN62uywzDW92t1Wo6uNZhA+EvD997I5qj5Ci2nRUpEn2zvp3vXON/LlAx
v/tykau7ELqagvLLVY+n5mfjSKJmsXPuFHnp7+0o1F28bzSymIyhhLHWoPF9fZJF
O1yE7IAPAA0wrnlMCY7cqv0ObW90fGNvYs3CrY7xZR3xhi95VR7hv5FEan7kYZbh
zu0EBjmSLWojFa5xduU1zPOMSvhE4FW2LYpZ/OljzuVu8YT3C+T/jOc9lwexcOS6
B8e0zopk/uGwm1eeWezrPpSN3KVpJnOqf6EKz+vEcdwSKrfyDvJpdFIuH/pYBRkt
hulmaoukL11VxewuMxjBSLI5xzuSP94PApswnUNbooWjlBD8laU5wwvDv1ceLFmi
25oJ2CYg8w0eH7n1vzo4FdLSuHZqQycIGgzUFssI//ltoAkTge3wjTckk17bFjkA
eH7aW3J8srpU/fzV3ZMm2i2ibj41fEAqv95P1+pq6WspnNx4b0mdeUeCTVdXQWp9
FywemUbS+qLxRXl5NpKSROi/Ul46Ryca/+mDKSsrD6R3/PwYSLCd7VSlgCXcL+bq
riClquyafGka2CVie2HcCcbzCp0eON79S0G8KhKh/geGilSHUw4b3rN+bFV4Mww+
/KqXDfpmLtSJqvaoqQeqNFxzjura7wJdy/GTOrLNILq8nyDsgRRcOhDFtsDc9hRU
4PxoHOk29bwOUkgrUcQK4zo87k20bMKitBzklkSvjaze/boIFsmiMWXzyQFkmJ+r
w7CMTZD9iR964fpjLZy1C1YCGD2GRrMK1Avp4Tdt4xxrv4sw+Sma6G8PuIbtyhMl
g1DKov4+blzrH08KMpm2YWkTsFctzR6AK3Nn4KhB9YoRHWheq2S+wyFD0voIL5YU
FVoQGuSUulanfIz9cDapMTOSG8LFTlCz7ln19RGN38L62Jm3cXmWlzaMKcaojYlg
nDh2fueshENxhUHiDMMyKH/t2UXkxBhRmvY7sZGKEFP/P8qA7CtTTu7BDyZO9AZg
h+wJTypnesuuqmVsxgMQri3UFZJXcfopt2IMDl0RWkEAZK6dusvwDXgN7ofouMN8
rcCNg2IpsgW3Si7myhpEkmSE0h667HTBSb6Fj/rpU2lbYkUDIT73H5txpdmFAGjQ
kX9PA6Fmbvq6c7lamz5OPJuWMXp2PTFc8WUi1jTFM/74A1/UD9q64+vBt+/9FaH4
yRMAIHOhMAPEBnrGc20bItsK40vpatLG/RwoaJdtmBpG0S63FL2m7T2XQM4zpVn6
2uK6TbNNYlpB0t89e6e6tB9C6ZDjP8zvz9WZi0x/lCOiXZX3CowSlH6bxG6JkIr+
vosqm8vCDWKzkKJsxw/ZcCs7QDGVTOpsdkowUtNXTNExl9zZVE7/r98ae1i6XQaV
CXwHp2ouQ8nCN4ttXdNP5XggceXH2JM7dZxJ/T0y+3rtEHVna9yi5LivQdNOoWnw
HI4CMoOHLhuC2UQGCuA5DxN2f/BVyJVGJTbZvOIwSlbPWQt/HgGG88NfRKwzZSWn
6Ze32Eyn0MwwLd3J/klvxZQSaiFlyTa6kyPChqxcTnMqh0Q4Npzpmx3zIvFOHAl3
xaZsx6qiQqJmAGTmA5CT9W/jcewpLafvAtjt+uCQq2VxbtUyNEtALe4FyFLFPIBh
ncTX+ofnCdjIPFteLCgEiXjXgbsVrOAoFxGZ7f4XgUwqoLYGNeRq+ZbeG2/X8kz/
`protect END_PROTECTED
