`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s1RZhe/fVYmiroy1GO6HjeN+tkrTaHk0y1Vrj2vY9KllaSke284T157/GEctp/tC
uZ8IWMieFXQb4hzO/74EPBav/4VZ0wlki8J3oFhQ6Km67AnEiTa0991JperbpEGr
XsdrDsM/WRMVpCozay+3xHYAzqGF6Zio8sXtflrliLNL/9beIRN3G8urKwAbn6sB
Av9vVem8KiDjW1GzZ7UZ3F/LiN2M5dtam+JFiajMTa+JDxziYNtkEFN+uHbXy6k3
EJ8rxEGalWk7eNGhMOpvxt09F/PonqKtIU5GOUjgIQ5LVdFAyfhlvhaSTTlDEfAG
D1PMVC7spl5KxR9HQSK+xDDyLNfG8tl746hzQqDzO0uTGIkBAnH2zfBNAcbSAmUD
JhnxsEAApsAqAkf8OrSLq6L1tPar0kY40l3F+tw42RgjlncfYx554jgC+C1xBv86
0G/tLweCg9ZDdE4FOyZQDbZ1Ld+xyodXZJ4DmTwyFzyCkfZzVGyZ+9BoLsFgBV10
OThF1FmStOpgXcrXoE1RpySCjJ7a7FKKztJkk4y128BIdSp0nEv5bjqym/gpEtnw
GfOwbp/rmmnA5PQqJhcaSwBKkkNAAKAKcUY4AxhlsgvBlEX5trHZxMG7rnYM+j2k
2nJj8+uuYIe7mJFjG7VhnC9IFVDJys0ffWSh+nG0WoDM7XlauHW7twTM3BcOnLuJ
QePORDjwaiwDM9aTCfcX7PR5JDrV5lEC9QZcUXomhknYod9nZ9t/RhmUKDt42Gh0
q9bENCrN3fneWq1/XSm3VoeQ0HQEdazelXP6sno/NYJf6u/HmmXSuvXrM2lSHVYV
mN9pcrJ0KOpF0KSj5Ndn/QzOQsZCLK2XDDIIYMvXV9AkUcVLdEZ0BPKFo8ukbQDq
ksdUjhuDyTtzvKnXp4REe9RnmpKVTlIbRz7eJowGKEtvp6UIh8fK8daj0OkNB8Wz
3AkUsguDrqRoHhDemQAJppSjXY33dpreq2spyLGNEfUNzj8Z63npym52H1b1FElt
Mx5cC0qIT5DiYuy3Vgb3WTr4hsu9RLLFG7I1+tuhushqVwgupVRLDYi3RufPgXTH
rcY6OLEShoti6EcOisbAV8cw0vvQKeWiRisljXAc/EDrdnXbBnG9Upcp/DxOldav
A2NbSHiEQzk5Hk1a52bdaVb0KgLkHtZ2p3drqPltAWbJT1nVi7hz1UfHZfv9+s0C
8ZTIGWCqxC1EkHpnPgNt0o6pOFwd52C7G40sdScDdeCKXvaEL+Gw3dz46C3vgvLe
MBnsLmNfZicllVVWP2gnJMW8UZch1M38hyyYOtovjLOSTgpiE4BhLBC99S6BGjg8
fHS2veBoojN20EqMdQpuZFP0qIA8Z3rxOgbZLuqkyAYrppSKTujV9wZNKiSGsIsM
450tgFG1y9Q0PwBnoY6VvmbIrolBWl8yoWp2kcdwJdZmc6FC2suCH1WOWnfJEWpJ
RBR4abNEQ5+DXQ8hfJ+oeMqvJ4VW3K9O3YLVbqzn4gWV2rAi3R9QST3aChPGAdLS
DhxLZ0MoL2tsg54m6u+2aJMvxxyVCq63BQgcyCymk/Cq34d9FoTl7zB5WmenJBt8
LXtSECnsbltw9IhPCCD+yVelt5uXM0QlfJ0IGNysqOU2kiDnMvNTYQDvrnXJViSf
u9iif1+H0n0+sOj97zBeA5N8bU6QCuwXt8Rxfq12zwA+afixk1AW83n+CX0fJntG
JzSp8aaoMfy3EfGkMyWMkozrTaIbrYj+yMHNZyiMSAZkJF/oghSKuM8iZ06PTpDm
KcLiNy711E4r1UqBVTwmlWhAAtyYYQRojVqK0ddwgdHYydIeYrX7VC4JGZucScVk
IUJyDpnfqxC0LcWzruhOf7v+OuEORYeqZ1q8wGpiOoFdzGNrLstH+AzO4iC2rYT4
KVSqd5E5tztP196eVDTZmNNOcmHOSeRsKREa4qKJQ6AsTrt5Rxg//AQ2+iJC6R6l
hNvvYRD60TXdbhn6uaRhOG5jPQ9+1Tie9r2eg8hj3vCFvamGekzypkMfHjBlMt3V
pdQHdPCTgbYYFCnmJFsMhAI8EUy7oaBMrUoFjMqPGqqyGLQ9p9xUIslksr0W7MgJ
QKbBa3msTD+D3ex6V9y2b4TsvliWaO3iQ4wNN84/OgHGmN0e2PbE2rXbehTFu5lZ
JdrwmXBGyVszSqHnwP2I1stDxj31BL/0L+e2xCuNcFffvau8VxsPgnKsuk1w/oco
Yl7UhPk04aoL8MNBPfTwot6fBGuI4hupXjzYnZWth2a/EPTVSzXDOXF2WoJf3uNJ
44F2uVZ7/Fs/WGOE8oegGL3hstFjSyrOpbxgTZpBAyP/WHpJbGKcr6NkJgYAmhQ2
s7szFXu3VFJnUXXtmKW2S2tohalKbej+jwZhI9Hj/j/IqMiUHQafQ5NQFIKyCkAs
oGtTq9sp5qrXi7pFUPIs27VmXeWHInBlr2PWR9fw1vAtii3Yiano+od63V6d3Dj5
S/ac8e06LOAmZks/bnupXnITlKlgA6iyWp7On2Uiu5AfGlS1spEK5VXXkJmkLlHr
57WrlgfVScPrvbJ/tbKdZph5T74WZ6QLzUw+ozLqKI2rqhLuqsuF35pBHJYBP94N
N8o49+bYvC4ZCDLAjNWC2W+9rqwhJBgbuQrEsr/SsDP6x1Zs2F+bA8QFn/4x4G+s
yihZlHZI4bTU6GubLNGLhZC2PaOI8mHn5yhP7KWAE4+fcHYEjkHR2C1t2If5Myvd
Jij85kYAjk4Te6LXOrq9vTKyTyUOC463d66A2U+hqGrKS9/8bThZMTfDBbAixh1W
wa9OHiK0KnezCdSptPYL5T5BlSrUl4sf0cKK2ZAVqr2wtJQrLiC1mc4RLeUk3/5D
DuBZUzvuh2XyXo7rx72fObZ8eV5oxqndhDV2wsNpSnQ77x0P/0lfDoG2tBWPkFlN
t9ozGCVD6MHY8KesMWEw2/UlsOkyTg+O0uievMJBtXGEU47eZfi3YQIR5FgUlM9s
ivHwlKeuVluQm+7i6Mj0/shEXbNZAAYGk9NLF8iXFclTrgfjkOsO4zckIXo3eSXu
+de25D/9O9TpbUbeHOJC21etdCwu0RzJmedRm8XSrGI8cfV4r1xXxy2EsqQmP57l
EgWHsZDi/lAcU2k1GBcVYJ6oVRDH3f8ProO2RcDVVLUppt1FoDWCgi8jnFuKCqY7
5qC/MFDPhCNpdFl39imG2W1KmFvnCuTjaPryHxcC+k+d65uhZL9ggQX4kII7gIyW
v9VOf9RT7LjbN9c1dHVRAyeg6aDLL19itDRd2PAm9JcQhEaU+bGJjrl03FsYm0SK
s/EHPyx8WZcuCJGi+01CoZ9AT/xosms0ePTQxISo/j1Dd/phElH9A2SdhElFKaG7
qAca2ZiMNXPM0aw3tO2k1x01m3cnQYq7DmSC8xm535A9gHjRW8eTGFpjHgYKZMql
glhPJe7F/IB6cqEhZQEQN/2RInNZUWyhV1AmHjTc9E/bAsSZ1esWJApJkCRRgupX
iOKfOl6vWBmYcczVtKKtIpQRGwDKHkmkoy3KLI96OluKd3wmlDJ3vUuATTtMgQts
CSCbLvn/M+Wm7xKdOExhtZJ/5ItcqwgMYJk2Md4rGwRLlrKpzvcMFl9bU9RM94dx
CNCu2JwB47gZ0HMRuGFJJpfbpWeAiCwowgyslqZ8Uk+m8lq7uZt0rDQVfHGDsVSP
ycLe/S0AsMf3mJGXYmdbeaYHTrs/BO8yGQQtxJpZQktpSq+9AQZANpyLO549mn+q
KCp9z9Zhdg1pQOyk3BAuLJ4yEdROw85x4q4N9WsRSSdDVpJacnq3zOHQ7iN3CNNI
vVJU9N6PmvVz2m5xlyJmEqJB+FbYbIt4LThdVsw/cEsIhGrX6/Rx4XCG2KKD9qTm
OcNAa0M5EBlzq3DiE5p03dsBWK0Y60ev5bQQXd/hiOijr66xcYDaa8hfBMgNcZMJ
4nyB4PEVcx7kbGztf4BHJPBZr+jEADkcWtakyAO+xvAZozj4BFVIa1jkE4Kb+ABd
vFtrKCQP+pszEO9xiwn9axbJmvDFhLCnSA66IJfiysNVWEv9piYgP6siek52nOUW
/l6SNuvXYUtX5Nw9ZfIuaKXEng/kQowy5DgBpVdaIXf+feXBIu0TC9tVVdP1R0oK
hGtb22T5ZW/RD2ul6zqxfrGv8adec0m2fGnXIxRM0zAO7zA+erIb0+L5w/lj/4H5
5WAXfRVGyY1PKnXWq0mm6lQLvlOtcumhHd2+kG7/FlGufOHOsUYm1LuayrrtXZZV
fykp/63WDCz2CN+km2kEcFU64GM9uwOwaI92pL005S9Lf8e75yfzhtth9b3fTUJW
SYoYoKh/+LI5rnpD6uH3ADLaUghBe9cY+QmJ2u84bgWc/kP0uMvMJ3995jUKyGcN
SCmzHaG9AZmUtZUHYV6lsqVL0BZxc+sansMLAW360u2DcQUPlxlDKM5VR7GnmhUl
TANVYOqo8FA2XeL7AlApWmOU0TmGEekqvgsbsldKH+osVa+qyryfBQ6hQ5bQLxwI
1p0qQgQcM4bENDo2S1oqOFyow7O0klyfg05CHdRt2FzWQG/VvVZeddJ4yNbWRduH
DaNlJAXVpnMULDdswnaSMsVw9YRS5bOAeYIrHF7gxjjSYtTNrCJQGH5nfBp116pP
jbwzxqmA887mPPR8N6sH5Wb+k8sMIuC6Q2u/VRTZuZU4EWqFFculkXpKyucAGB29
w2tACdI1nkXDGvKHE5t2pSmERJ8TYDyretEhc765lUP6AKdMrRTe7UxZFXZwoXhD
dmUH6NAEpYcQqIMvLczypzr0cwOpFOr1eVbJqjLzaZ47THwoyC6LHeElX6HL/YKV
q3RQ1/jOtN9X2lEBVbIEDKXKYC/oGJN55mTPJ1e46MEfrRhSSsdi8S2fwsn3/ttl
T5bSx7HEey8Lc/a9JZC/MoPnTfyqXvS1xdw7XXs55pgrhFR9InCwzrYfa7TF/JjN
X4nXBEBn9PK5qeujOsia78VzwaT44whGRvjThPPAwSiLhilaJHe8xSaheNB7lPtI
lNTCp/bOS9H/OojBOCGI47NWjmsIT2cicBEU+PVFk8w8vUqrSsunIhkpwjL+Chij
gJER8MUQlwJ/scPrDB0PK68Sj54vV13R34L8s80XN1LO9M5aj4erD6ESpO1bcI6T
7ZjHtRQbjbnLc/ee0pv3mrsZ6KK10RLYSgDeAPqAcu8o/YscR9D4AOlrVzmIWrkU
2fU+nJNUPknpTue+OpU8Tyk9+PgjPdn+QShqkT61G7Go3Q5w8eo5cmLfZ5xw5T84
koaPDvipj9ZLoIbMJSFzo3gXeJRlatk0UnHCC0OcPyY1YKW3HwYs9LrcuzB6oWaC
AHmbwyRDepTvpKNlMA1eQ0mhaz9AtFDP9oh2vO6yWtUlJENz3w2FQhY3/SL85GgG
V2TKkPWLUX2a3wcdFBn2P3WbFWuLFNmsF0Swrq0dil0s88WKTrzI12VfPFUssA9N
Q7twTvj0XL4YcLYb+9Qs5Yub+7VGjKbPVvyQdzkr3LWC5CYv3aevurVraxFhJ9Lk
Bfngin7h4fTDSjiV8uYm6Ka4qLiJFCdF1Zb/8ie3UNsd1ayp9+QHL4XyjtVgYnOv
IHSNzYiVMjMBFo3y6RyHyNFTmkkY8sGAiBxGLWfIQDR36+xhwFdyHti4Lg2WwJWy
1S1HwXxtbmohfGJcaKboOBdXO1aE7C1kVLragU6hY8h/4hVm+SXhxnQ1FWYTRmBP
Y4YYlVadYzg5GtBFDVG1Xv9u1KTJEYsQXQBTt1DE8JXmNAiPw++PRLUjTCjhjkmY
08QUmcl2aatdcEHrXBjSXmznKDElC4CiXS4TvcEyYg1/wry9o4wAZLqT0eB2JZG2
2hgxToUs3rLzwCYxRk2iIliDK4SvIfD5IttnomGdcN69vi+MGWb1FBDk8yqQZQbL
0v1Y5gzLCZFhLaXBSqEJV5j791OqlmHCyvnXPDkkymRDEtEdqO6XrniJFyXH1U85
WO2oZqyiWuLUcIQzI6fuPm5AV2soalq81iXCO25yeUegTLgsb5f3+ew1ONHEDWMo
YZmZqNnL07KX36Y8GXmHBXgCvHb5uAm8vGfdKvRaT8HHnMVr4WeSZafENFdJXleB
XaNPDvBxK2fGk+/IAf4v3n/+fQWUfoIzdXdggldlw1bz/vtrYM0BwGewMkyBQAmW
4uG2gI6hl52Y1whB+Lg7xVZtEMbFtT2hfMEWSjAKtADDXsyRm009E4obTfik3hfa
u3prSHgs+IBfQ6LiCwarkHZSHh/PgOi/U1mtUM2DChzNiKIozeDEGtmLpCDaHTYL
wnTgTWe3teruz85U+OImhoUSVnAibS8PHRbBzQBJl38OlQzn6Z9nfXrq8F8fOUF/
FVrePsmbWM4kEgI+oHIA1S/M1gyH49dIXjX5KpO6UZEhcGnCfBbH3l3rfT+fEvh5
CIGaI/etJJNnRC2+NClpFIesYFh2Anh3B5VSUkbUKwImLHse9gW3B1+IyLW9wct6
CHyDQzx5WpFe9MacQYAAoh+cuOMylJBanzjPFBeeP3DtKqt1QUKYY47EeNksw9Go
J+PQEWKCbPvMZ+O0m2W3mYlyAPulKjJO6MPJGhXOpRY8p83O9rPWebwRscrVFhJ0
7ReSSebm5XEFSWiyzXfuKmMn+qbXkDy8WF9vopVIRxStDqxuM3vxEnb0XdTmdt+b
ObwhIIIc6KusjLf2dedmGwotjqkS0rrNML8ETVYou1XojxA4eeS2y3yTwS/G6f4Y
pOhbztjkS3IwYzufKJ+RlbEDKQAAkaQQR2qz/pm2+Mrzx0zI9NRF0gxi/QNmnzDW
GoOA+r2CmLEXliohBA3IXvrXknejw0ElUyfwVbgU36/34qS13yYyotUB3zXIR+VP
ybetJpWrJAi7f0juMGUoYkm8FQ+N/AVvKqS+mF3evsbXsojALMVAQf7MyVH54kSE
HZjP+Jve4x816E5TdqenN7tnPjbQIsyIdr6i2beelbhfW68FDBLE7/own6GjW6r6
Dqgv4/hWPjmCwmixfkesTd4rfi5+IVMh5v/qhBTAJeRB53kGVWCnkqF0KSWE+c/z
R/q1I4qFijVQgvbQ7Gz54PI7yx9vybL8UsTco16Eip6D054z/kgC0KYhBipBtz7Q
mWHkF3IRQnv9gplQXYu4pzHg285BugYHP1od08jK+miPtRmWiNEeK7jXvkYZXrxM
uEfcA9CeNcCqcIQeZFV0oQf7mEfkC6R75bUzbBpNegBthVMIvwefmIOz+TZ7JXbk
qylzDaqI0FrgEBq8H9eguj4FY/Q3pin3dXhjQHjyoaDGHzJlmrdeo5tXxC6VThb5
QiNhcfEYNOTlPrO/Wq7m3FpxOb6GwuBzr5Xc4po8gE9hJzBM9A1nVtROS8m8CQ5J
PTRqL+f3PCVajMoG+XfOpToa62xYlZ9Ea1OAQRNslKXJLY8hhxyVBfoD9Zr78pDn
rmS6PWB8qQQT/Uafsq/SioD2TOphYB3WFGxUsw71lp3O+tqE5sx9w7zfBhzSsIbJ
PbLSxThYyct+GdapSP6uaTtQBrRsOsCilKzJXyiYsZGJSs3tYQKd3TwwkQANTFGL
OqW/LI1EG/g1FmH9oYNQRpZN1u0z0ddXGv1nqg4XQjDucnumlIWsQ6uG20Xa4mIi
gChrTfP39kxXILFa5UH7F14k8nUrZmBFGhgbWfzwXNP6mmRNHW0fmyqtMdU2nOrI
yHHCO5A0DaDImJfznZcBN3C+J3qOljQd31ovVOTKG4QAz4qaD/UwraPlyfgKsdrz
D1wQNlXtWao24WTE/ajyldx6Pi/twIu2W7SNTNvjR6BOaeOR7xHuah1xZJo6Dkpg
6STtgdQLQ3VO4Nh2ijkyCEDEeooGGC4BD7FJHmHITYA3wrJuq6WuZ1gqwYD5v9qK
JqXQl4utbSzzDGumgdpd1CvYuR2tsiBa1Rdl44MW57Wv6jkV00NEgkYReMqOeJtG
C130CuGPJQvF7rUNFGMYqQRV1WfMI3wHXIB8iE4Ttg/FWNMov2SFjF+hgVK5H9q3
7r9xm9jy8zAgDrVSu2C+Yjw25+tF0SQYYiVYM9A7JYhOjfO1pyE8Hdu+sKYFZQeA
D89XxqVj8bqigh5taWitWizii8V0L/8Ff0P+9d7PyXhoqQLGfaHGvlKGKDnFfNmq
ZgqxFp/AZSmIb1TXiOrVdeuUedTMos2b7iftcdjTfBIF45aEbsm52mBcO8wJGEK2
lNSEnEXPE8KZYRCjNPTd9Pz9A1Tm048/41/+UQ9rkQOVkbiSedMJjnk9baivIgqR
6SwDelbBIObGo7EoqDujGgHjcacH/P3+TB/0XKE4Fr4GyVkJLA8GAlHPZPZexDwZ
d5YS4z/7GZl3Oi3hGZjUlHAvWmZCl7z+ZZKI0+wR8a0n3vRYZBbdT5OJ0tuKEOKO
4HAspKfUG/aXLvlpsUjPv8/Yr4q57YHAxKvjYyatJdBb4RKHyKiYseDvDuewvWfe
9j99AEdyQiPwjlIjOYmydVlQfCAn8yL5TDHNTW2BlYM+ACnaFRgeb8XEaXs9/APP
L6GQQTXaB3gJP2otosugK66+0cO4vwaOpkJ+f9nSbuq3thsx0MvG3dpyLUQsj38L
lrKVgPvotlaswBixpzMoDRBXHHPW2llD5RdnkcQ9x7PcBtJXpahLfgd/2UNqloMc
0Pdi6n+Tf2aELAH3sDQ8bo3LWSZDEnIH0SDcNQaKQPV0DjVQU3y7AA+Ufl2i4qZC
37mAUgnRZwTdiNo2jM0mMH9/WNMKYZjGNZBEbBf06ji5XwUUCGUVJ5TSEqzI2ZpU
L7I8i4cbo7gRD3SCX1LbwVjlCmv05wrk9MaUQIo4FfB7aCj8Z225x30fcKQqBAdq
5Z0wrSY1NNDiSooUwwIyXrd//6mbwEtlf9vQWeR/Y1LaRDccsvTajJsbSy1xvpWD
eu13uuqsjgcrk6R0SW/IqNRp6cou+GaZUMNYiHMtctejkmRAp3mEjqqgeGZivkkt
ibbgF8yLq3duxCjWO4DNQW1TwCb7ziiJWUnrsiJlsuA9pHVAoF5DTQGFsJ1KhXeb
PDOBqWKnGUWSNrvSfWxnlrUn4IPCWV3JCbg6rigmT4QPdTyljce4XmF8P+wTfNwN
mLYUbwPDwhgn1nV4LrhoidxHpZUiP7StgG2AAK+KVpM6PUg3skx4rwkp/Fp6SOrp
DnIWn5KhP8XUxy2rRdvQgr6tQPfyXyTcpGVpti8pG/1KrpoFHyPOz2On9s/lQZ/Q
gYkhYBKPscYjlxMP3MAis9BPN1FTCcsrqIgdIUtwQ7xPssF9H7zAM9xpvM57Bv1i
47QTYuXq1WJ016Ylo4kKvfeNRTv2UZKjBs+2zgAzrxJNXOOeX/Yth15Xpghk+rBd
7mMnda2cG+IBmSUBnLc3JFABpkvkR9v06Fod+o3+00B2aBJyq5s+QxQn+iiTvnlk
W1lizJ/0S/hcEIco5qQItYB2LZ1f5dWiG5mUFhN1OtPxP0WW1hE8cUREnsHEoHUj
p2V1I7CWGDi7KsJ9b1xVQw7Hti7Iy2S9EUzs0iW6SEn8LpFXOp8PjD4wsaNxQSND
xsWEZrqWxmHfHn4jZeho8xHkV30M93+bI5BnlK9xkH7MHCkGt09IFX7oyuzODNKB
f4bpyLGNlLrnFNa+8ewdwUZsXp4+Khe1HKV0MYD9xJYWAJEtYy1+LFxCpaVSCGQE
j/tIkSoIQpTGCiQAMtm3ibb6+R1MjNUk6XTUhx65RQN4V2oihguGw2eMsX1bnyQU
v206QZaa3tjemKTUEZI+FTFGDkK8ibVckKKkDOR6jGYSQ6f6Azy+fzkUXkuBehLh
VU7nOMUbUX5why3ZOcCODCadQna0L/ItNHGtF8ofEYSEp1Y7qVYu38h8FX9bU9tZ
57jsykqKpGOwDMahmTfYF9x6zyz/O4M4IT+IPWZOT/bZmnug3gAX2/B/o0/2Xf+c
M9jCaNcJ7d112bJAb8H2JrOIqAij4r9v+ZOhh1HgGtSntEFD7f3UrgruPUhfRSxN
DYvcUmdfNozmMYKgmDqqG/AGPQ5KuGYMz/sliRtOlWkD4B+zGASAw9QZhGh+9REi
oiCc0oJ7jQf9UbEww7UdsYlRO6EX8d632r6RsZkQTarFj0PhWI0ILQeXRI7miF7m
PgBEfZdDL3rFOXjW2Iqylu4Fy+AtmMQ+SniqreH3eInNavwLhTVi6D7rP11MsUCN
ZKf16c1mDZjWsya3G3nrycLPX8Sgt23BrwaXP4aisgcbYflnRoD434wknlfPizHI
ounEMpmgEwXYLKKIvQjEH8AGLxBb6+qQtP9zzYinpyrVutgm0hp1SC3PDBjLxYdx
IXEKuq6YC3BRqXiyeNOASmqv1WrgcC8qF8iZkSr/6X9LKIPL0PircnI+0R0bGsvc
li8CtzTxVjoR/bIRN6z+OVu+gTYX0MBqsD65ime1pOJzzHXptwLVYkYyxSEeqFx2
t6X/EXZaAUWTgJtbTgwsEmwtx4lLyYBXcKIGc+jidVj7zhdaiafjPBHEEGxRgTne
qlj9mPae450CG0sMyc5nmAIgJafHtLDeQ+zNLBDsARbxCJEIQqnZRJDA//JHS1jf
zhvw1iEMwsOSAFojkR/ScKxQedtnlVHUMYWR82d7mOZ4N36xRoEOtlAyal44p6Pk
45vJAdSsRoy4/9sEeMEDSt5KfqOK8OF5zb0bzUhpsmVxBXxbl9BDzhyngAEV+ZzF
XnLb2DDJ5FmVDrWCKCjpKf5roeAq/a4j+rVrysQcEvWanKMO82xGwR9lncEnTguE
QxjdMIjFLdY/4dirJL7m+dvVXObVWdZcPEJOhehrAWqU0qZ4rOtsQwCUoyta5oqw
t35qOD6uf4LmztxffJjehFcae9vpyjhfArASIp5DpKft1AnBAhAusnBwuBzNRpsL
zzpYhPCLuzhklFrwQVE4PxdAjZZ41mPEsszd3lR4CO2HOp9ap7gUoH+jfAMcFHM+
AS3/OeDNaLNRG6odpq0FFZZcaffdhqAexHLf9Et0VNUW7mrd+rwXwh4bcmzsu+a9
mqz5delMx57uK/RcVKPbjdAfjPKnpVDvb3wZ6b+fd6CGIxm3+9FMB3tov+dhlWkE
s2vv5cXwUWWbTBnsZawTGX70fGbK3YeY2MzmA1pXbe/BUY/m3TXOSu4Kv+Kv5W54
YWDYLbvJ4Gu6b+CiCmTJJwaPgO9TjiekVZdaT3+Oki/yUaTM34ak9hXgSrIAlIC1
I+XuNogrpqskeex64zDFxMotglbmtth1gb25mYmMklNRJIkGEXhc4eCg4S88mIB3
xOD48gcphPF7DYMngSAYSG6ZrQTDTy8wMvwLF1IpYkYzec+41fjr7PlJmqR5HpWU
xWxoFCYPKeCc0rdUC/PMmPg8txuDxRheiYDFebjb2+tskb+PZkaC3vNePRkmDW2S
2oM3cT+BfFNG7CmO7BMK1YM5Vwk/bm+hyDqDLLpBbEefW+Y1PxF/f0mIxU/e+HAm
9eyViumJ2HR9xzVSqtzYyiLTEZpaziHTAMILpeVv6sCEZmree2sDE/oN7CPl0PXQ
L4//tqDBAK8bevmZgnJdg5CaN2NWpj3pbbdyZZDhKi7AE6mKKZdeC3tabLehPKZM
1H75z2V0ipqpiioMn/gB9mWvDcAxFPcTUsCtK3LZgaYGTsn8ji8AQlL/VTKGkK/H
qYrB2NFUVLNa/eDQ+bZAmcCDTBWNuYDZ5U/4wrigqrupCXIlcl+FdzePjiZO7WcD
iU3nZmZPul7LQc0xOZf1fM7jCshqdpHcSIaCnNKdNRI9/6xPKOSE/OER3i2zZm1x
pv7pWtcVdADe8MqKhs1YNQ8HCe+9Z1lfZEISp7JxGq1dvldhh9tbmzgcp9cvL3A/
sqKw8okzmSup4lSEw741nUoLyphftwnrROtyG9FRV4vtWYPNoWKyTE5qL/QzPuGO
NjlD9L6UCm1BH0HVLvVRk1an4PoqbDzv0KzzIqXctesCsww6rWPA1rsZow6h59uC
ce6zOMclCmD4CsKYqknzS3fBSTB1h43MG+VNNUNoQEKsT+K3qHSOUJecdFfv0r8E
1BKcbL/rXvDa0F8PkNMKemwASjmnAOcgkqGMZN8kWTUYDbBYxsbyJ5Qqnxhx1QLq
GrHy/65Zo+zdQFU5CQ8TThi8VqfvkCt4A8Po2GzgLdhfi7NhqMmB066gk3d7EiKv
b+lKxWb4bOc9+5QpNhoIqE9kaWnPAKzuyOgCKt/J2hvzXdelvD9JbXvZUjczWut5
kbmDXqTbL2M30YS3XnhVgN3/MfZSJf8ZS8zHQVfdCj7jbEqZmvWZhtanSVE/PLKD
v3mm3McY0eZvFR9za/Zc0GVKOPiJcf6keJCDEY0DDjoafp1tvYkUKm6yDaqQBeV5
dd5EJcfptZUW8rDnitfyHHCPO6ieqR+zmL2ZP3dciJimF2YZPbNtd4eQByG++jek
yXLu3WdpaE4wpMRRjSdLbqTBlIMBXX/KtxSE52dp9k9a4uSai5J81AOXyiVyyfg5
5C78OfiAwRhuyM1uorsDt0wpRq9LBEGSVUArMSuR/9Tn/djQrHcHX4AF1drMvCcS
q38OT0HugbR1U0A/zvmsJiseyvA0J5A/WAipolVAMqqzUC4dNVl2Y9G97EUPKEx6
32+zfCCVmJJ1vqXxF7VqLXRxXH7cwficwNifznXz/GFkxflLfFTrUj9REFE+SwSd
qP3R72O42xqLW+3ZpDms2HfQvRcLgKpFCGsSG4jphtneMrj84uCEy/yQbnmltqMK
DDacCx8ebjnPlh9uXGRNmuywSGk90dyeDA5An+xHRoC9s+Tf9Zlv8cUgnEYc7B7Z
qzftKJzfTXE+1C9vNsvqDGMGpViLvO4tt2L5BoHV0jVpe5KzNFLcfgbnoIiBCVoZ
gQAceVGY0os5vfPHzDRXSPCkPQKd+nW6Gwf7G6CeS4RjRxesnzyEhZmvt8wsr8Hd
8yYSPLSS2wnoH/9BVWfP/+vyk7VeA4v89UtOPWeKC3mPVBPsVPbwxWSr7A3R63QL
9mNMUQG2W1OylvEiumynl3atP4heDagZr6zsHZwr/667NxZqgJ2XJ98lVHWzXO16
anotMKwTPHZfp2tnighekC10QePtxf5ISOBC9epE4S5YlwrOSk8Lvnl5ZcAPcO7U
HD8LNi3LKrWz+Dbe/Nwwz6W40XKydagHznnwXOBhNOAaOKYx/0RZMTz0+78IZBth
bF4zPDw/iQI77nRclGK/6g7PqrM5ckyi/YVtVS8TNGCt8kjc0NDGZm06nQe/nce0
q9R4sGHvMTk5H1EyrFImIdvsXLi1z3cJV0W9pfbxeXN42bnEXzGANXe9GnBxxCLk
A6zXYO1kczXrkkqEU1psCAS7TGhMtC1z7iBgz7XQnSjUOWUhUuSZ4a9GTBd4Y/de
BBJcmhBosVbxt24qT+klC/bsOYdhg/g5L5bTMy3qiOiPXnltkHr1F1Ong5pzjPbK
HUsHBezAjnY+ZaS1+esATN8dI27ALhCSNjhtVsJL748jHRm6gwQvVOoLMLuk/z+V
+xQWtQ6JUb3agWaNONIZsh4ngaTMN/ibVvjJsPu/d0y1c22PDAi0Yaa919D+kW7s
FejnyMuxWAOmr9Lb0VXK7riINl3IdzgU5ifI4FMm505PH2KwhgKQXgp3E/CJkAHZ
xKox7WROYOLoCAxFXwMNG+9FP7TXMfcq94v/w18WiWQXu9GPOWbu9c41uv5UrsGV
rY01aDiQa9EbV1UVFcSEislh/GxF5VtnNgJXGddaR2L8wVAbroVYWI+3ZUdm8KHM
0zQ1a2Yn3c3nJCirADQqTMA/CRpU/lMgXhL3OnAuyu9vCxh56dJE81gR8LL4ar2i
a0/yKhCQ/gYUgcJh7wl8JTKCcVoc2HUyAZwaDgOqRJd/QkqrKo3SLgsFhfgOpLwp
/zWnXjCp3wuE4i8Drb8n6hbJc9MKpyS7cBXwazSTleodcpNBWoX6WbehHLdHgn8k
dD36eg0TmzL9l9u2XExQOwlTKf0/PCMqUCdfU5GRR7nX8b2apNepyyDUyoR4ymt8
71Gkpz2sHeVhSkpVf44hWyj2RzK3yYvU4uUYXnW+mukJfRqJrSmfSq8dhrEUVCGs
q2RsoNr6QaBWeza9sNPlrkxoAjQ3aMZWtP+OTC0WAHcN3BPvFrpjV8BYnQchjyaw
mSvZ47NGZULyy/jvQk7E9DnZBZtpSyzalTXcsmhHqfSErovPrrZ2KXfz4YQFlDHF
OMwdsS3bFYu3iMfl9B7wYqMxTYXOBSYMHXO15xqXXk5VF0lrujHZPXjpPPfHIKOF
ZVqbbPex592GRjApKUYdf940tikvw3tPGTrTGMC4dWS0K2DCAtRdIFKzDk9cKrQD
WXldNnWqHWtF1GMp9ejpWm+VMfTpIubPizPN6KM4MaYAdKLTR9Y9MGu8MHmdjghV
+nOVOvtyDEkTIFJPMqnM9DZDLuyZigW56V/TBhJAveB7bYULg0o0O6kDPc3pUpTN
H082/OwiXRtIg5I4rCwrsVszdEHnqZbuopmEx0NhouIRs5/rltm0CVVBLM+2qhKE
NWYDUkxos3vu12NLEZycij07mX9n1vsNZbyHcCKOqxH4WB9dGfVOgerIyNEkpFTJ
qI7SW6dWEp4bqbZx/Mv9k9ek69Y9tLdsTYfzwdvzt2kBdTPpVL2Db5P+02CQ5X1d
0KtuOEthXZMjg8SQ/s6c0A65N/bEc4bjvtTzr2BS6xI+gGvf8SfuXiI9/u5/j0XT
TfjbvyTN+PNp+HmF+YtCup+QB73rkaHLSR0uYnEsKa0JIiWVZ+F0q2yQxTcfXRvb
kKhy0CHwKgpwhJA0Fc7gboeO0YzHvpSXoJMyGU58ozevL1PA0deLwY6ERT998sF6
+cipyUIvDSLkurEwkDTmHWXPRBxoUQbSgt5Qi7nddB3pPXAqIGod1qXti/bctSNa
dVAVsP/hy2quprE/xwQzyKkCmATr23bF8viXsDaJJos9TdTkKxj86yHL3rV0hlgL
vvucgFw9q6wKMtw/2bVSY3yQ4TGHY0OxRJM9QtyZhv9PEvm3TnSkHC4tX4i63zE4
lpUnueobKEcLKOkC6MTFDQcUgwP+J/sFFgO/T9KCNTGndIf1vkWof5Ji3xsNYHDS
tQ8I8s+9z7UVduZAjQMd8iqlYZ+onmFy330ew7b3BkMz+hFOYDdNomRAXZKxGrMy
I8g88xDgTaldinjoZhtt9FZ7o+btS9nbvSSgiMEjlG7OFFrB7Q9tYe7kK5Rtxfu3
4EAvgwoZstPlgwJdwzPhXTd8jGlOttKiDQx7l5xrd+PK3KQVaPuTAcAEitJvjOTk
BdVI8jlqCpzekQ24cfNykidJ5J/9gORGKdU7U9Hoo/m7uNiyOam+dp8Z2SheYibf
aBbW3E+J/iHFLssrzSTzZnqJ1C2khmHQptSeDdbu5RdwSBQmVrqJ60jwgOFUX5On
i8Ds9KL1hPooIXNmS2zIUHDvhulrruM5qCK4qlFSr64TPN1AmjljBQiKM22mwKOR
eSm7eiD0yYhFPRnY4uK1NV/x+njDrv4ps7Z1WdNbckPi+6EmyrvZByOUdnghKX7w
7J139eI5DbY1CgRGBrcA0Ek5k+D8MxHS+C5k4ejUHiFO2sPi85g1+Oynku5ixflO
onNh3YQ+9z4fZOu2Th5iX7lo5nOuiV7i1LsCy6AKbXdRUtjTaJv7JDdq1yLDWsj0
Mu/9u9/1SkznC65CL831SsYfK6juuG7ro3vwM/o6F30fDF6vqBwGcQ/NgyQ5x3zU
+3ETACTFZHOAcgilLi1O7IU0xFxqVa9F5tMhO1q5FxZ3ml6HgSeXWCT36+II/14I
gi6+rNyTK7sn00rqLaaK6ZpW7ZZQs6aY5IL09QKbfPfkmcRRaqtoNT/dW6X5yO2d
7jQstESlkHzLSkY3k4M+x0Uk/aWaKBJmuBuj8ydatgUcw2Rt4dWAJiJYr61Whq2x
E+REeuGZ6Y2VNIoJGd2QRqXu75EUmvk5MomdUIjKroKglwa1LUdQXF9nM8VHxJQp
hvFiTqPriK5LF7KWF6F+5C1GOsqjKltStr8OwzOUNH1QAONmz5a36DJ2vi2H+/Qy
lKhlINH+gB7FdxJzuPp2I4YmhCZjLRQXtA06Hcl9uttft0maRv71v/a6cojHvxP+
FBTh2AMW8KTc0LL6lPyYBENz9fXEvMpiAHzO+4oKGZXVn0p6JGeyiHnN3uyPnlyK
7q7/YKLqpE4VDW23127IdhMiljgFRIB2Uo4Ir1Mz0yB4pHb+761lp8mejcJ5yVp8
R6T9vaHjr/ZC7929OFixAvsK2UzyvjC3Im55LLtTSKykw7YsPvviW0GNWJgFNG5F
tOsq7qms7MOPkT8QvNc55lVw7dveJheo7TFB6RWLCiNr39iYEabhwE/LcLqkqTxi
rf83Oy1dQtI1eUpzmZDrzDELu6aGow+WSZwDa2XQLrqEEHeY9zEZSeyGVBIHcpPi
NpROT4tGueOm4uC/JluCWs/C7VHwcJlKfVmw/O9y8GZB+/INkrqX0LDEkJcrj1g8
WQGUP3zrGAVZA2PEf8B9F7AmX65mwk5P+8sXeqiuJ4Gr1EsMzcPDXdvmwIENqCJQ
ZjO/HddcLw58ShB2TWQ8fkp/vAADeWjwKTaxOMFffcCPiCDMDY6RaV0w+FWWBIow
7Tvmy9I/Ka3HxWP0hbfWot7KcZ4FhfVsTF86vgEifl8Qtm7Dvp8oHerEz9pWR21c
Phyn33XrXdLPaVZMxJFDPr/l0Lvah0rwVrN/PhztkUu4z46uBto+L5luCXbAHRdW
CFals2RTyIfCEzvg4lcvhBNLPp+l/Z5ur6xmMki0ThQJl71DaABRzJUX9mf2rGIV
Y9FcK1d73gtN26tCznAL6g/gVGDgUgDQLbjIHcOWs/S3OpYfmreNOOdQEY+8Ktj7
5UCUXQoL/FnUWfQQHtOQMClxvJtv8CE0dtK3rRbCkA1x2f1ZOCsIkwKBl1Tbz/cT
MtafLxWFvNeAamq1H06HHiGnKk+gE0m2eeDLXV6yF2hUKBbBtCbpa5wqfxPUtVzJ
Nbb1gn3bFOWDSodAbueP7T2RNH/iGoGRNRQhcm/Ye/1H3XccEJ96dNRHDxganTtX
u6riFNwJ5aVXWIDU8dZjJDR7i97ypEVlQqfHlc+o168wfaTI4d3P1kTZm3wRJpeU
XoDjCr51X0YuxEeZHvm2F81UdEeofVUEQ9F+aMLhe99D7hgSuHOVuFAvseADV19r
fXVnWqTGNZQg8b0LvacJL4Ksx7k3d5rTckjkbhr7wUrwggusalwi+1cWYaqqaq/s
8A0Qm5QPKAZ/MVti/QQAecLwYQ3xT2FaaYJLYV8e1gOr/hnUcAu04STIMf+7F9Iv
vuB3K843Ty7DWL2KOkePrDkULz+B13G786A7lhvefHJKjzgg0HX6ucPLCcNPB1Xh
MiA/y0HoSIVT+w1yqakPQ2AvspX2dI+GYxcAwEK/+NAdbMu5j/gFtaby1Tg2DK0H
AOKQ59v0TLf5D1nzxa5hTPrXIvziJK54CgY2JoMmNz5MhIV2ui87Cx4x/Ob7Ug+b
GGTiZ63sbmtHWimISg3rxfo86fOZwlTl/HxiFTEnLDocyrm4OEmyCJY46dSq6to7
HEIF8UfjI+XK5j5Bkrx+HIqwtjuWks8QDm82bJz2TQMEeTJyUjkrnG4M+hKm8RGC
/okEsYk8xFoKplQpYKamVLgiO4J1JEQ1Oz47EEDAODqL0JMr4UC9NXgCZHrfWlZq
hBHs9NaNUs9x1DObGHrnPtDbYLBszODA4VWQgTcCM6Qp5O/R0cdbLzbrslY8u+Oy
yDompOxVnHc2AoAjuNMoflKGOHzL/Q1v0t2ECRWl2gfOqhe7hMp/tgNYP9HX9UVD
lqJ/OAX7n0Bh5ucewLJxgB3L5452F/1D3nGmhS/rB2MoRgvFDYD5nrQICUj054Wv
JtNASCqK/3j7ENfCslEXZfUzyer3RoelJArjanvWCaP3vAnJaXY/yaQp2gFNx7Ay
u192qO1NOQnB0C4uFCIqjIUgGm8ZqOjELemNR6rn0NJD6cTtSBMDuM0nnXBhrCoW
KDwZBXVdJBDbG4E8BMUApCIwpX9J7/ZhVFYAbONp4vT4kdcC1KSBXNjj1k2PgoFe
k0zTlNnSNhANM72Hue/Ge2+sTG5Cu1OekECWl/9yi9GqZjuZzMglPyr6HYQWZw2U
quVSRmyuCcPwW+Q0HBN95xz7HLbQNYetqT2cxhB2mpRThJ6Jd4O7tkWkXNzv35Ls
jLH7iNeH1lroPFcXU6unceMCUWjs7FVjSzwdep3FoZYq/WVmGsYWl9q+BgCEAcdV
G+t4JAiu9atQZet+S+wJvel0xVyPurHXDbctAFiX2Ba5lSB1K1NpB33m4GxOB0P7
/sJKEmIsHPW3iUJeOX8uUGOvkizm9ub875eAjbYoZfbUoQGPSdsXcecOTYQA0WET
ClA7T3h4KNqGSqgb4ZMpWFsf6E/Ul87tS2Yfni13fiRv6Jr7u3ZBhMjjzF71GBxX
0CdVmvuSLUgZHNprr6O7UldkvztF5hzEfaC/d1tzh8VyojYLHR+hL02RE6m6cOOa
hBy+8FlsVQFAyjWaoYy2w2ZBBYzI3uuk1tIlNrZMosU5vjEo++XXRI9tQEUo2CJp
9SQxXUp0wE7R+n2D3kVf2OUgrwzo7gauwgs25INNmDtd8FuUaD3VoeFQ+/xv/daR
NQtO0iNmNp95KQqDgG4U9cZXC0u2I6Pplbs/wCcr0ImnglCb+bDqHpLA7Gr/rVkN
BPZKswRj4IkzUMqm1T3HiNXofDsT/4h0ULKw14YVqsdEu2byjWV0w6Dtz6vNtVzD
Nr71VQYp19rI83LR7aBPYl2QBwbGyPgJdkQtLo3xl66j0XUuP46O0PeZq+8zJu0d
Zqqg28mTtcjdCeawElvjTxGSKOd5AlWvQ5y/dmVl9p8jLRDudvlIw0kExk24dUsz
T5nAgCTyj25pNW52KI/Ig45NHwoPCKBjYYh2e0qriA2IiUqChI41OxgDVuErSfKh
WXAfch/NwPEHeJBgXXjMFHMRzs3htTEbhn714T8073DN0Lst+Zw6zV1W84wSC16n
sPLxuky6NBK2wkaUnH/RCgHM6XyQ0ilH91I9P+Y7pxCehba/LMkjUlKH5ckrfBz8
Qf2nrgmzu281S4hCofer2XeVltlFl0mULuWNM0/jZyR4KZPZRdxQ2/8/8DorTvNc
v/PFy8Fj2xW+wUm0YYNLq6MdwCWd9l+MTKlOVZ+Y7n9LZhisSRWyhaoZ+Az+Sn5f
72Zk7N7u9/wACA5q1h18ozD+KYsLbmGSO99OszHyjwcbxdqQhOZCIroA33+AHILg
/y44X0iKYWiT8Aj73/m3oaP6ZIk+Qu9sXLp8nXyW5wq00pWvXaK+tMOdr5CQBEgW
K0VTsphQCN1vE9U2AMzGma3BYxZVBh+B5qiz9trJW/2LmbThMx7a/eCX5L8qpjuz
YSAKxl9aQ+KWlrUuuqg7Jjpjk84ObFWsEUcx9xr0t3U7OTqwbn5nbJmO1ejI0G6z
0E9Gvy8FDiVYfovE80ufvL3liFJ0x5pND34xXZzjUsuLRS93bx1esJsj/FosG9DJ
NketkNAA/FkMbXXC1VxC9cBeUYXoRqKKZImV2csq1QErx/h0eLL7nntjrEFYioxu
uNOOiQK8MnN+Dxqpyt04TyaHVfET5TOvLYlJgXyzX2pT5eC/wO3jFA69vkSx3/RL
0ptoWziJWem8Pl8YgRops1fTcxCOryLUTFp/wN54559O/2Pd4IX/+xIDD8lSHL6M
0KX6poia1mptBrB9KFXZrHxDv/owSkznyE+JZDv6yf8bM+tp9uJH3YfsbHku+SH6
2rCAi6YHTG2WNWuofuc/h+W0yVRpp2cCIdHCb+81eiH41pPbv4W8mJ0D6NASCZ9e
Zz4YnCm4ivVonOCpQIz3V6NoutmW2jNH6vLoROFm+8CmajvpKN0H6qC16giGFQeO
+oRcxaZDmDzQuKaZoKpL+SAelExcqcSuvtoxtTpDtFdW+67sYikOuFQnVRYytE7n
8UX2ZKbYXTWOCLHk6BvV1ENIiIR1Ne7EHrNbMT8u+1YYE+/sORTmHSZtrOqVbJi3
Os8dySpiLT/B5J71ctpfUdiYJ335kFPdXWc5qaWZ0SGSocsgm+Gqlj4j+Bh+1u9q
T+4ZJCuQSOL8WVPhjmlvtvwwXkjTIPraxanbMIGHVKOEWfN6qPxrpCQwRKQ8w1MO
rhLAqBJeCO7hunWyxmz/gv7CRq/q99jAjFBo+0+6Fy0Yi3qmKQOQq8W2yuKWqtf7
k37uwTqa+SuIgGH/dUeA46Vj06yHpxvP4AXXahzdjPF5PFYLOpeXqFqwrrJ1nDNE
U4n3FXEKf1YpjK4v6M9V/mdcDfSBsXmBSeoZsts0vWW8Ya7tWV+UF/WEnX+8Mt0V
tFqkwDPE4WvP3NxzAJ4gJxyCB3GvgZVN6rhH2lMDTW4tkGt0u1L8wCBMtq5CnIf2
VH6a6fNDxtJhCjIXDR3eHyMPIFVG1zFJj/yiJ0u31erYta8abD4hvcTblDWXAQtO
C1zob64puDsKKzf13zkVjlc8LLQBETr3OIxYl8UZDg4IXy1x8CYL6gGRa4NRS00U
gfaUjJQ25uDPsuW7+9OgI4FjaEtzQLCNdD9ZypfoIflTw8xeVbaxWeKvzy4O9OdE
dq3ZITaSscRNfEk8q39T2YJkcHIOFWeunjMPsU8UAXGHVQ6jY6JZ9x8gEdjufEVm
AydoQcJrPwY/i+TYEfrmBqhILw/G3DB1yKUSctS723kje43XUuvc2zB/SDfZ7DzI
qBgk0RhJ3LuUz1hN2uTSjbNMVPfGVNiNAT30+i5/nkC0VjI6gJc3+8OjOgV9Ryl6
uCd3NGACoaBuD24qqnMCpD3eNm8sw/Pdru3g4qe8qrm6WHe9OuVLEnj534s/UBT+
Cd1wnaj5l5om2LedB0aIaLGJTcGPTvqmRC92qKXqL8bNZc0DF1seTQY9z6SMrIJI
h7jwURWM6toy3/Symz+ICua4ZHgPckiD6f2Hh3TU0i0uDGxYCFf/V6r6gDh0qCBa
zmlxaUvSXl7lzdvdVteqAh+yfnpyXZSdIaqnuL3cFoMmE2UCu8DzpO9WIoRsTUPo
t/EZBsfRac+I7pd+CtlvabUUk/uEhovcPCD0uJmgA12jCjKe7JiRtenHl0nGS0V9
YXOzPC+QVtDiQQQFFHkNE++4C8xiFaw1Ywm6v6dvGaE3g1xT7cJdWitiwy0FxU4p
79eeHSAqNYR7M3PX3GzSPMroKBNCZyQiSnn5waiwG2lMh+/o80zbKUK46k6bw4/M
fqJyOspD1hMoc+LZFHfaQjPgH47ZCwOFEGaYJfePexsbtVvfaPhbx1AuevUVo9yC
um0njLU+gGn57ze+raN+jPuOkuPamuPvm1Xft7NOj5F0VxlFE0WC50qB6MtTSAUQ
HD3yOg/LRSQCSH3YBxPXZ5YIEmOLZGf/dVlPCJMWm0RrFQO3XGTwA6zE+eAmppx1
LIVQZ5DXbam3pjNtP3g/CNP7B8lxJPwz7NW8Zgvv2euFyuVFRX7BP/6QY3+IpMrJ
gWFjzA9f2VzI0n1RhjjyXVQSm/x4YWIMJb4buyrPeQmLhgKxqTv0lNhT+tjvsFx6
PJNk4Gfq+ichcGgTuxtJ5hzniGnd33OdUENqRjrXFSGxSt5iEwcJROGP61efS1P4
Kx65SOrxN2ltDnlVJZLuvVjhQ/iTWzvY6qdrLDIfm9EW5CdfRQU7lK4xODSVRJQt
sc3c1Rs2xC78cQezBuyo/fHx6FPQuFd7rHzazXnSShc2q4qiVrmEMnTgGKkASMCr
YbfrsJmlXzsHAUu1F24GC2Fp4VqhKL29ILWJVivIULRupxM5Hq30U8gEMqVDPd78
y2VpCyqqj6PvXM08pN+ZHz7zB7Ese9JgoO5WTTJB7OTVPJXCa1ZfjuJ0n2Lle+oz
qqWDkVzFeJ9odiBzHOROyR/9AD8m61kblW5WsOhd1KGQblttc8WQdNyjMBW2OiDj
yClq8a+vaAbbpvsewBSc2mNKDU0Po+ixgPNt9St443NZgyHMeeJ/dQusEQ0Eq6oG
0YWrlMpcrQrQ0rOf/0+HPRp5pM28y4rgmcbjRIiEZWx7ntZfNG0cCyq9dHWEMHPb
R9+3F18oOHlQb51kaqDt1VY4epZyjobRoVnw70WRTAOsIaPaxES7ka2XKH1jr3uK
GlwgAsYNTz/BnPnES24VuifHKiwvetkrjD2HlGkLgfNL2zrv1wruK3lWDhO7Je2L
9avc79lc0x4ax/7zKvLgdUpW6t4I+f7TnmQJ1yym84yaTpECzqlWZO38y4VE9Q1k
X7zWWkn8/0Y0HgcRSNgjNYQbh5zqk02b9ao4yytfTkX/tMnKb/YCXfaUZUdh7Uh1
GLKF4sm+a39eQi3pO3Lqld/WJCn64vft46qG1bmVroXl0+9rrtgYMmjJRIW2Am4E
q8WKPfFKPI/6WBZ53517WPEwqq8QByLPu52Q4jC68ATl4toTomOqSbYtokkB3i3K
g/5iIW4hIMA9ZbNKxsJmveeYjEGQTQIZAbHdxOD5PE+G7Fj3JouepG28RG/ZrCUC
sDrAEX4X0qjhr4EnOxurqtOQt2WWMsNhey+tZXlWCpEpo2GdZwODf+ATGLKVrqkF
mPYmFyn8lvU6gonHbUWvtOeCVwPjRkT3cSs0XsPU8cpphPEoilAnL5qsR5Xlj5ym
aMg9PrLS16/GI7lbS+g1VjFCDeoEhoDeVWV8EEo4yEhdOBAlk1qyl/PDjol/pzRP
08vmnBhyO7YVmfeuxw0x2IqjaznyRnyJPT0ncpUcbYfIsMaqMc8cqnEg++p1x5WN
QB+no/d6ON9fc+o/8X+kMQGEM99d38YXdJw2FSgS3BY8PwDeCDDXng0iplBFR4/m
BTiF3fDXY5fWpTo0KNsjsiZ15L2HAemUDyv2f4r0Jc+DEh9DafYqEJvohhnTLZEE
zjjoXlPC2C300crW0vhhraGZh0gLeWp1to35/rrA+nw79b2TM+LpmqzNY4ab10Uv
B9U5bHGL3wDF9En3/lu07EhHdc2C1Izdq5BEfAz/Ov5OrFU+bXTaYWegCOeXpi60
8hp8ZJnfj88TSnJG8uouxIV+VGqSwlZU/HCfddkpHAsj/f+3DAZOHFR4Q4HEOowM
OyC0FRN4Q01gvK6escHCP0sInSiNFa8PPXVr4cX9G+NPIPgU+aMWKvkCZKyApSUX
dysZYTQCXrGGMN0fiL+Fi13KTO8U72UQk0IIuRhGOmuTFmtyBJrHBXXzDuNcRssJ
jFVhGd70zjh2DQEdwnKHFr/7YTn4oX9y+YN9liDVinroyvFGWwn43ZRvRJzDUkgw
6ocPoogKDIvXb4n6/mCB5/l/csMERcyHmzFXHpwDw732jR/n/ZQ7gCYfXk1ZuET7
ilTEUdXUrSCkjqYaEfyGauLzPmZPv/zYQAb+fbCvP4kWzib/dEM28AfjSqZctmUG
FW04VAawhFTtw7dZ6Dql6zXQZ+5HvjaZDIdSD17MappUEU8uFOw5bylc6KHds0GC
RLqbbzvbhPBCB0LgtDel8bNmf9PYpX+4l7IYkj6yax4jKwSTideinnoeqoXk3l3M
/xJMi9SmLxtquHJQFp1/zNk+pzLpS+sGppY2zIieh8fKkE232WqXmaTLXLMrzgYR
oVW4ij45VcUqLWmJeos0oDBQM+T70sE6I6fPkULgJtggLl/kQLlnlUtYGfM/jBQO
427pTnidluv+iiEENHkSdfiNoq15/K/RcNdr6yjfOil9xzNvtGhkRFFeywPSeFIr
J1RamHHJ1p+kJHDFY0IM7Jj9G9rLCyZnueW/bwJxfMC4HsitJWaivD5wCU75SSGe
teZ2jUVZlAN3JEff54+CHq0ZS3en0nqJeYK35IWWEcSuoQdGKdeNGJA7VDeNMVd9
YRnORWR5DyibHMg2x95GSZAoJcVwn3Z3AW5sOgpWCJL6zyjuiVmRme9AVTAksi5e
P5IcAnQOmFqjGObROkPpu4dAM8xrk/LLKx8yHmsIQkqEk8YKU8kMOcNxZ8XvkBU+
ELygkdKcJJvRBNzZyGvPcMETsPtDYvEMeUl1BU9bAw/NCIkXRfBqGz+L2TaxW2RJ
GCgKUj3OquBAVOpoyjnFhT8z8bfYbfHjDagE1cexaUCWJEk5DZ5+zqNcUmhGR4RU
hxvSLgpHHrt/hUlF8inYRTCUrD+GgKNUOvvHUwgyBAAf/6N+BZzMZlwleDrsrbG0
E5lnHv8IArR+MT0cUTi9dQOH+EN/IgNwo/2Odo+TWnEzHHe1EzfIr2LFPJ5N6hXa
EIswiEnfg0gBPdpl+ZwyYptS6LUnKSvzsFg5sCpvf8KTR1fi8NrkKXrvR0WrbwgH
QVYnkVYs/zuwirXYlOl4+FqakuiOIaSmFbPyfE7CsnxAozhWzLm8GkcaH9uQl/Mu
lRRGVRpYi6aDD6M1B6HKdexzcxSvtx6U2j48u8iZly5Lj88sySXyjGohhlbn2lMA
QgPMbo+H0JBwEbEol8yr4sYqAzlwtYztH3DGEBVFWHkQKcwapZpsw9F7IkuoFj14
U41kwzySi5taOj+sYirQZ+wMRWxmivA84AV+iBryGdUFJEYXX1GuNxTkp7v4KspT
VcvFJI1e7sgrH2gV5LOYzGyoqyEjhrwLemNymfWLxam/xoVPgrq8THZWZp/fh2u/
cbIfC3NAV0rb/watFYLMbIVrO94LdT/9GQtB7opS/5T8hUsTe1RH5Q09VvRtfuq8
Na40nT9TI/YEjjxSHRB0CqQ4a93G30Spy7wiBobPEZPSKmtSUte2oN11NREBy3ph
dPFvlx8RUoGefpoVsQ3n5OLDo6tmR1OaoRDsO3uQXXSRj+g3IvNWXPybPrB/slX3
7KpU5rLL0f0dhIEH73upampo/r7s4lUsYqjvGScnJY9PbzJhOwyRuJ6yOqHPSvOO
t3BjXb8ugIqCD9PSasLN2guQE5pM0pcDk/y7RlYXtIVqIFoYaEm8UgN3ioBVkLHZ
KWUX9KTcX952bhrIhKbmu52T3L63ANJ5UMqGX7LtH8VmwUlwFOeU2ZP0yE6xUFER
oUdICOKE/8cw8HaSvwC44fxfWk+kq8gdsDSLOWeNhq+RCAFbz9PVLydFqi7QW5fn
7K+otOHcsWa2DDRPM8G7OEPAH9D57Kz4B9JPWbIU2Z6KegMFeYfWn3jt76qTpZJE
5DNEkmXVS+LUuzq+sia/eSIYH5hQj/8T9CfPpvi7nzZ4wioA7aIaMuCzwuRZiX+w
xwnjd3zRHtq8x0QnWr5YFUYlQBd2mrgF4Brfx7NFIhrxn6bPrcChCnQks3lfwHhp
1eP4xoHleBAqljYEdorYca1kO4sS5hnNCmod1u4N/FZaNpyyemOzUYtgIoh/R1nW
Em9aL9K9BsjsFNhaEcuv/au6ZgEqCVtXBcOs2YFiGtY+RLzFqqx+Q6+kESXPZzEy
qfqdxTm/gwzbv8Z+2DYIEodYBS9+s1polnKYvm3EPkSI4D9NAhqSS1W31VAwLr3C
P9r10Kw67BF1PkRYgHq9Q/3q/MfJr/BTLyizgL2GFEo9jn5EjanyNUCcNIIX7s5z
EKsBX1TqhYc1iY53mFoOn5RgbmTnT7h12v7GzB/uiCLUj9TLyhThEcZGG46RrzIL
GPTavqRoVmGSUv1jXhc4m/suishRFeBDKJm3WAtkYFIwc2oUJ1vMxyuFBsQXZqrq
BlTTRVE0/vvllexmMyzJCLfsQKWn6le68FJqyDn1NYpsvBeEoPh5Gclf8wxorl2o
pCSx7L7HmaAXlwD3MeNOICLV+QlEXq5Fwesqg8IXn/ZnHw8vBwsc9OQ2T0ZBCXBN
Gb/F5upNViWKMiGHHPl9TcZplqV1rnlqq2HE5jS3mBO+01aABb5GSlnK+BvVTTaJ
rDhbmTRUupgD887DF04Tvy3R4AsayJPVtCXrqdnWUVjQnOUjTe8X2HPVhFb9ElF/
fBpJtFSrK5IZ9ZnKVLxnZEgZ391/zKFjnf+gICqDCcQpkZR/ko61SLVHMLzSCfIf
+sgGLNVyI8Pp7Es6+Iy2V8kG+LAQZnTTR/E22EJwGeKxgFOqFsnwAvPSlteMQef5
iA/qiG6ja6fzIm1dJhRsCIQTz7p79KxqoUSJCKX657JOsfanEzJfGp9gJp48OgNM
z4thCeRehFMPIGoXfK9ICacLvlRu+MPN/RACyeU0oAzaiqdOuqkBWy8ymVol6aWK
QvP9K40vHDg77q+I45VvDngZ1XsYYke5cwMNM7ZcfOFn9Ci7mc9ADdEnrUU/BzbH
wnKIB4+cm/SV4ESXr0FVMKj4ulDNSURoXiYbkblCqXwxh7BBVIkAiVgXDUma8Z0K
4keG5zSAcuaOLKoglT+czvjn2CIuexUPIuY0q3GEVByxYWhUyZ8YmYCvA+F6T+e+
Y9Agb39pys9XU6+TXhFWn0+RneZY0ATfnmFPSEETenNaiecxWgyRqO+X0aOa+Ozn
wrAD9FMJeORkzhb/4SF9EhjSeEDUXXg1Py15BLtO+zZ/yYSw39MgOyK3YgsQJamD
souubbnSIoXTrJ9GKXTtF4Cwr1FBU/X0zHJmymhGWeNhzpBMAOCUja6xtIMXyxI6
yKx1ft5EroIV/kQVYk8bwChZTrrDhxVq6Zu2tQeVZr93Wjb59pGi/5GnXgRJK0oJ
n1RvN8rWIPAhrG/xF1HaYsN0xGHxDq9zS02Lg091pGuUSy+S6r9SN9BV1sty0mjF
0EvcTzc4oton08cU/2K7wQ/FpkR+aFrVng9xMF2PI/CZ8rezeY9Sema8VwNw2nK3
UJWOsEibEGVtMT8uiE1ElxKxvnQc6I8LPctY/dmlIxs9quy8343hTTdFddL8WQxG
ASOvx6VCL9yaDPU6tthzWCcmtRtPecGuTVn4DddHyT5zm4Rx69ENjP6caw15NVlo
QOewYtVal+3xrCFZeVnBc+oWrU+3z/GRfu3lTS3PxGqXMY+UlKRof7RaTtj99gSP
pmPgXclfCf4lRww0PKPaFJzp1+FozEkhnwxza10LxjBHAz05Fwvq1E1+Zs8UubFx
Mewj7tPEyMxPI7EIwoWSMGoKbZ0YUO+5L+MxxkXpOhimUEsDHRApcVVuB4R+uM3Z
bc5m8ustJcSWyIOTA3HblMTnM2HfBv6wMFlqRBdnHdgnPga32TmOmCHsm7rAWif8
psjjO74nuENQOKe6V/K5+epLXlGLj/O9stSHfJjoaa4fPKSxOGSBErxnO/N4r5FD
ibQ33kwOGmW3KJ9Qu9O77R2fBRatdqq+DpBEUgaUBeU7rS/lEEq8VleFNR1K6j9v
hPjYQFU/vROGnlz/jhTP3FgNkYLQSycxABd76c6QAqzcP5HRP3kb8dx2YtJFM9Os
VfmJtDkW550mWMUzpg9G9pC4iW4e4f4IXuHUC0btwBILl5zyxgWiwr6gfVtjgOFO
Re1gYMhRdJz9b4twi/0DOO4pxOfAN3x7Uh9IyAW4UuCzMg62ONkXDdGVba+hkzTv
L6ey+pQFuLGDaSXgwkB9ug9d9NPm63MAzEWtfQOkr2w72N8XgD4DYjMZVFo3BUWs
ebOvIBZOJLPpNIT+deXr4uCnaL+NyonnNFRf93YmNDD01eGblEJK8a31XuCDhYjE
UW6SNJsDrdVnH2bKDhptWUrxrzLe5ICxny6MwVVraOQI0UMCrwwX1tHxgwhxMEbT
haP4fTOnBkMvq5u4lkxB4O4bbSAiDELuULIhHxuX7DFa1rFFyNtOgEFSxiHnibuv
kCM18D7oGdMfr10fp7XZ/tPz/dEzjvEjdxAm/6/kKu4f08oSFagMrcxWitETM7I8
TqMf2dK5TVLTSE9KSLJQ92gdOLCf/rC/Hn8dKRcicPWRMdk9oG2ph0Ka8hG6Wbjw
R67M7qQNWhNbuqcsVQG/WmlU/Yskcxihze6eVAPGbzlqkIKKUVrU5aLGLyy5i6Dx
mA5sx0uARHedge1HTJrZaZYOV4iD625yadaC5rY5ok3SF1QUaUbJjptBb3NF+Dpq
OtXJRwYLiU1cPqifps0QvWI87IiaW7UUQ+B5AQZT7WbE3ASsHOONuPMmKnM2zMke
gapqiUO5BaNYu/UuOyQp0BsX0rcuQz0CbJJIZgFRJ2Xbim8kBkoPtS8mc/Ozg5aE
NZpkT6FibfWkd1r4dTVwaEjeK6xGDVmtwana/UiULd4lG2llkuqq49Lj8YUP8MTE
qUckgOboFywSzFSVzZP/C4dp7cCrMefQdtny/vwMceLvSVcjOy3xsRUjo5HXXgzy
zfSuNGFCxBh2j4VMrrfAdU8L7lzhp8esGeJa1OgtrklMJunAzFO7hoTp9uqw1WCL
jlh5Z4OLXnQQrcVzljsEkMr3B/MOus6hVdK62/u8MggdJdArgERtkQJ7PtHw5DYG
9JFBBvJXiK3VBUreX3dTbYOcKvUpi7KI0figRfEP3Ake9BPIJaD6YrynDAcEJHHb
Zqfz57JV/3+Y2pU9tizGUkhA35owaWv/Dyfef+eJKDei5JATO2u47km0e42FH1qK
vjdoBokzrAhMOrzvEszWs/QM0V96VlsSNXQvaSct9uCyjg6oI0GLU+nN1BmTbKW9
ajpkZo+gAFfQ0sfx+8mut2yI9OKele1oGls0AkKuNdaaQUUwczwo41TNwS7KI243
vf2t177pqYHVUQHAaDEpBu+A+12Oj4DAoJVqoN0egUmFkw2DDNyYjqDFg5wFDwKs
c4mCjJBwF13becyWsgtw83XHUFpaI+jjE/XtMrl0iXKx1xaZ4/pC1PTZMI07xM1q
XCaOaoqw7peEoKyWbMFSdG/oe6gsQmIXqsm8vtUpAj3eFCS3tb/DKZ93U/7TLX7P
64sFJ0nYxr07jxv/4QybUZCOEkWQB/1OUAQe4oGiygawNiMFz5zAAvu+/skwvjqh
GmzrpAV2m+GoXbAM1atbMKQ4ex3+wcRSFy6uc2grYmLGMErfL9+VBzlsy+PWEhQu
3pRVHQ2HWjdkFlGbxTjzeRrXy+hxSSapn66WC/x2z2nYvqVqPAa/9rXlIhDEplB/
lQ0VjQ+wV4RNGL/dwzs+3jAue7EUUCNSslVI0Nk/Vpqg6xuYMO/eGD1N0ihd+sVs
P14uCBU9Lgt44WptCHwK7p7q21i8MtP1tgtYQC40x1VY9VAF1htkJBe15adFgMS5
kW2WEx/xQsQKUnzopQQ49MOS7siEzyzV1ks36ReUljiFtPupklh9hJCg61Iijr0v
0P1xAOSM1qyyATzkxi9Jdmgr1vubL5rpWiYhtIRbAEZ/xdR0cKc24c44L8Ke4bTJ
y4JCYkJPcV0/HTbpLtOwrajEXkwSdRBlkzYuJS2jU47vBEN9Kua7W2J70Yzp7AVk
l9R7VWqnK0M5TEOA6OJTHX8UFFUXd8Rf0y4MeGoiXPWjMQSGVE8FGGBk23U6OFDZ
Un2VPo/+TV1mDkrY6046+PS1VHPbZlmadXIK8S4AK79PBxehrX9DJJHiBcbGc6FK
XO3Wr0LKreE3JSWob3vUQT+S8VQ8amsPlK0Lyo2Tj/odRNGiH4AoAEhQZQ5/mWVe
2tt4Nj2Hr6aJqb/IdNF0/RWXRKo5KgNYVgdSjRbbXbWJXvQD78KTlFaSVl5T+iKx
OMD3jA0AnONPOeCcULYM+wuilE8lxI9bNKWGqRdIhMYRKyEvTcTBLO210zuApFje
RP2VVjshfgipi5R+/tjJcwETHMA6rbR351GgSV3xVWh4mVkHZvM3sQ8JnM0nQx/S
0mLWdMTMZa0w4ueTX12g3eVp+FWsBd8kgkIym1Ba03ppMXEBPAgxjXWbtCfYZYbF
Z6HugTV7TbMytCI1sSxIGPp3ZU7iEcdiCG/qR7951tkRLqJ52kbgqP5Tl0vEDpSn
vKUj/SgX0DiWmI99tbBnJM/LwK9AlOHGgz5fVRevlJt2fS3A/Y6DtMdsyF/X8dvd
YVnEw2/XMzzPpptgq7SxvWXcAlG9ARZ60yPN+Lt2KQDpHlAYZQDqvyZju70zCqqH
6GekLuMjCIm1FIr5LiEd6hWyGkRwRTtlOk/Ivn8uKTiYe6dM1Dp+dyOIKT/3Jqzu
c1G9OKyohLOZEBGkAiR3n8bngrjWn7L6NbymZvjMFXvxbeLW7kmHMv5TxFBFQcmE
iU52AwRMwE6eFAYxCXL7pExUkjlpN0iJicWpS1GgSBPN1jba0RURXqux04/ppr6l
jTyiExtFqzADlxmH8YD1LI6hh8dujGuUKnajwI2gzFL+FEyBniaHMMClxuzLVaZ6
zCQl1m5mvO7Z2WUdWH5eywkPzSSibAHWqIyIJeJuZe4d0Og13CQ7nVodJMQ0MMbg
LmXJk9HUE049ZPemZQLEQdtpAL1LMecwfGW0fkHKFCT5yuQc53lI5us4sCNdXgsh
yC3qeAd3kLSdS6X6stJDm5OV2f0/2Mehd7UPHcVuy6aX/ALGF0z9Il8+zpKGBXmP
F2PVnkaTVEZNM95mKhuC90pb3xuioxv6x078fU06DM0u0UT3f8243nJktXc0U4nM
oVSL9SCHJQ40qXf+OJNh5LOk2AW4AOS63UU3svLR90ekcdZGMokkNwh0Y4B9L/Qx
5WKAuUNesz6nbUEBOOaiIhXJeoNKHBd7uMohdYMhWEkfjP4sK0fZqv8SSNIbh4y0
cAS4amV9d8Nd7PRlNNrtV6k8EFQnUjcv/QrfLN3JPojgFS57WgEsAg8SDnZe+nFY
e0A9XNuKAPgGMtLx1YXibYjEJlZtVOgneexYe6bzn5Ylles0+ijuAAEEkh8QLwsU
KCDY5sU9r49GfueCPQbt1Us0lr/iPSmaW38Ks9Oxx5GD041x+yV9E5T6RXQmSOGg
lKMRL+ltmp0gsJjeKYnPdxz9QU/liTl0/8YIIFwPgNjSe1ndIw3FMBwJSQq1dj+U
43ZkfAASPMwi+JeonqCU3dlD40ByBJUN5g9/idFlYU2DipB5kYXEBuGQgeIbkN+n
JOO1GErUd7rzHPxtgav1lrOAnqxEHsyQUEKwBYr2EGSnR+FgVXJB2vUPHGkfrOJx
okKSX2Yh13A2F0goB3pWEC6Db6CyPZPs63HXI6ZD8ojfjkonkmYqg/9nU6nYc9PY
Be4XkWSFOdWoZDHw2PGz+YaSAuVwsS67EblQWiIcWfEjr1RS2UH9YEvUL+beTqXd
BnEaq1kwypl/4/ZaygK+DS7NDkK5xHKx3/SQA1xdDJteXRbqqdP1n/fGemsillaq
VqwR4E7b/EMBADRwoKGlCkDHwdBApAwSSbKEc3EijbaQgIcGo5byzXxP7JKxcDL1
BAzQg3pgnyODJXDszkxXjmEsoEdYPSiwMj1BtiN6Z/F0c0HAmqb0RWlzgevaOHUc
5tgR9BS7mxnz25W6juvH50X0nIXZSgvH4856BrdZkzuKct3Fj67SK8012/l4jkeP
2Khvdtc2gfNfgUm3atYpJekkoDPWHdHRUu65KBbZ3xY4qJAp8yM3MR0/3QFValGM
gDgxBcc5F0gG2KE5uydDfRsotnd0rtAgfuRu7Vil3NiLrt41c1DI6zelrUm7tDXv
U0+YhxI1SPJe4vaiIWEUNcV+I2ubRSmDiXnZXMx5G05xzxx+A66aFpZoq48EL7WW
f/rWH+abyrzkL7+fyQO+Rdx+HZWY4/YWIZjiZzwT54p0P7/8nV2OS5Co7aw+7NKc
WC00YJRpBG5Zb4UTZsqsi/SowKoAvR1pw15qWnOB91wP0bufVhD6zxQbXYWVFlaS
kF/nQ3wcUHNqy79/xqL3iHcBiRSxrUiaMB2V1OCChcKR2NG8wO8RbNCHV7qMcyvx
RMMX5aiATmeJLAIxnHLYVwnXtWY2/J62XKo7erUoGOZXGbRXfE+qo+zK+i0zCYdg
o2b2yTcAn7dtXW8YOHGYSqZxADRsejrG401aTOUjBXwI7QNIJfi9qwZyWUUDNIxv
Uw9l49o2NKmnzqEgAPOyJJVKboSmBf2S82KfkgSQcRsa3Ig7yaloChURYscdcij7
ZCuw8ZgBJNE1aBH5paszn95zd47j5S5+Gtj1ICPFrKgNcJRtZQtPSQY2sg8X3sOi
fcAEsIyrasRyMaj0fWCYXdC6/L8RLfofLmdht8tDBhmpbEgLkaSaxoewcvupi1y7
d4tf2XV5pu9295RlHljXK9wavysuVxAFLas5B/yDC1EN2h7/fzMOiooLD5zx4w1l
hFGVGycbChrkv1K+c+nPz/iVMiyr1YyMa/Uq9imcuzGZRoAH+p0XYpVFFlZqziQD
jZgxY3YizmqaPiq2hS2EfRLlnij+d9lnMlfuMaM4ZZWWlUOscwbwVfiZvUML+nlX
9Dh4UMVpuDnFNkcpX+qVFymZCXvMfSxhJrAUpLNcqR/yOu1BJn2t56Ls7BCJ43BP
zaST8FttMGYdVdBpx2PqV8gfhKkpJAapE3Yur83MW07Q9oJzuBmCvP8OUoUUrJPy
n500B1QdknQdJlWX6otcz/2vWwiNuedZs8Pv6jjAkX0shnZt7JJTqvJaVjMVI6Ww
r8fR7ImFqKfzF84THnx6W+9wBVhwGetiW6WiJ7EAFu4DFs9amEf9JmeSJJc8h+EE
ZMr/FGnI6Uk06Q3rBoOeXvS9PyJ1BHER1jPkcBgRMXvJul0aO+QVVdAYjcQQdfkb
deGCpAK9qnFQdqA+Uipiqojo2QUbaoQemNrabNy+rYkseO1VM07KWKX0Folx9kE8
QcV176ztG9nNyZt3poEcfASOLXHH06HG4e6hOZ5XcdQ=
`protect END_PROTECTED
