`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8a+jcBQU064Ff/mdRkcIjf+zVHzfhVT6oIsMZJ03HrWS5S0EqrnU9cc1i1rlApdB
pN41N5zPOE4NsltXvzocdiLzGGI6XkHhmNCXgix0yAa+0afwxFwdUZDOkYpkTVbk
P6EuHRrVFyhbg0jv1MvJtkUsE8C9JdQAndMkZkzJ25d1n10zSJ9dJQ8tyUums+a1
QR+GtFLRy2ShU20kX3HATVJ5qVZMfqKgt3oGXxqC/UpDM+JWKxBGK2CIBYn+tw+b
Hx2vRw/dozBxQz5NtlzMAw==
`protect END_PROTECTED
