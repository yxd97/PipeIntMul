`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBzKMrZrXq4l3h1U02giPOS80Tr/jqhQaW1Uwr6bNWy0rYp5pWFzFRNqyoWYYabO
AOjTACYp/NNhF+TLJYrY9qhHyVRvfhj00icfuKzgsWg1SjofFQg6WiER6p1eUpUf
SUNftazO+iNlYb5vinX2S2/Mr0tXhqUVMR0Wrp+MOmfDNVEVa9Sb3/BCAsKKdWkX
0qP/70Gdu4Mta+UqrUvftasWeL6PyWvTI1PwmTq3Nv7wmntyV5lRJdF0czR2Xas+
On1ZX7BsSukzLuxPSyKj/lRrpkwj6CchckW7g1/qRg9NYY9wiDqR5bLlTESRmCv4
`protect END_PROTECTED
