`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
225/0A0nui2YLuc4IT3KQN/7MmoDdF6IWhTjL4wETyYQ2L5dqMwWVtD3lkEdyyhj
O9pno5y3Y3vdVyLsnkNyzAqmRCauqPq0IAbm5BxTYnnjEajSmklvpiEl4OLKxfCD
+/JXy2O6T+4L7HrogYK9P4C5N7fUyhQstTKQB9FGOd3fWr+vHFkudLFYWCUwX16P
8WX+cvoX+O/KfOn3M5zddA5Tc9dfElku1sY7dNTafvpJg6vN77NlhNgaDPNnZgar
MemSuFI3htqoVGPu5RyN+6XEg+oAfmWWPxVKJGruhifLjSM+eJYLrmpnvgX0ubWa
Hm+uokpCm1y0QMVdAL55N7PnHjl0hXFONzvVp/2K09safnvK+v/33UgP42SbnbjX
dARt8RChn1oe/abPdx2VxWxLc3VVorR//BPeEVePyoc=
`protect END_PROTECTED
