`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j6oq/KXsfpGfJy3KS/ys+PDSZXQ+xd7iI9wfw8e/jWGXnINMKESXN4tNn4ZIvqLV
SUNKmI4IUIt+ZJP9CvkW+IZxqdNFJCtqms0F9rH+BxJSZpKDLEkUvkq5x7E9+4tT
PL4QJLv6aiF8LUsqFLUm1/lLthn3vAB/oN/Pnt109KHmw3K/RQxh2raF+quzTvaf
FybdMvnOg1G2HDpybheQanEh915e4ZEjc0vDcO8ep+45tbYAQuJGL4cPk9yJ9yoS
ZeHH1mwZg6es9w2ROnmDqh63mJgltgN27HrlveF08gzlj7KUw+BS0Z0B3NXaOcZH
yJBFSgCPgZI57RHHXk0UYDExtvif8qV+BqOAFyjsm+6c3Ev4nxfU1cnIVuHpVDX1
UG1VePIdTn2qk9IZUrV4AQ==
`protect END_PROTECTED
