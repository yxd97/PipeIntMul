`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GbpjcNmWMYsyEY2KV+UQ/6q4Qdf4aLlbOvtgdiL849wNvftTODbozie25F7jQiRV
Xi93aPC8ZXI/XY44LszyfBG9tvRUxMNXt0Z9ir1nSTKNgNgklI/CGe75cgK9S47s
utt64sNS48AuRPNxRN7Fo0yLniKxNPh55vbqgYB8meNud3Jxtc7Wb5xAeBNxz3FE
YtVJZcaL5KaTmBEurTpHDw2wJris+UGh7Kspe/hTlz2zyC1I+Rzy76H48hZ/TBRy
3RofeLODHEnmHaZGWwyM2USC2IZeS1Gzgh/UQZB+y9qaqY7jmSJvklOJHbGSVF4o
tpDQSu+mch//QajgeL1d0qgYqpvWmSYCz3vpmGIHEXLxwM404zk/F/U4ZAQS4U/o
Yy/ogS0nBzYkdx2XYKJ8NxZm3Pm5L7PvQhNAxsOh0UXiOln79YoUD+nZHkbtoGwh
LnhlAmFsXLVzwbLkAY/R3qtnT3vGJTPrtnTKMIjHG0YAG/Apjx1PLJNFp6EM+qFi
+KpJr2sU+TLM+Q0ftGpAxhvalBpoMMtOIZHkTY0/5ec720Uyzh9PJog3qx+9BF0D
ZaFuVaoRE88BCt5hB7EBHh/oCYeKv34vGaWIVNTn3LjHDnbKQSK+QXQz+Muojtae
hszwZNRqSuuyjVA++nddgRTB24LqrHpoRPUBeMrcMQOA5X0lDBZseonSYCDhEPiZ
BlFpDYEOg/PpX6qP5Ijy6D6GzB4EjGGpdNUZbnJF9JPAZ0BtCKI1faLsvr7s4cUv
aad32I6KZSaEmegjct/OS2P5krEyxHv7gtpInKbc4rlfDgAtXlVrS6WlSN0nBd6E
e5GZ25NtS1nj173jyISwCzOQtg3VdSZK2/R/7LPNHgVkLUwMGKtUpTVD2/1YhzHT
WDtdKmh7CJ9FfcWBtVcKVYsUFX51RGDBz4XGuwBPsL1BR5iXaTrj6wyvGFHhSagf
`protect END_PROTECTED
