`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ksyzk0VkzY6YizgRMvv2eCQkxq0Y4uU1Hkjltw6lfPri4jQFFo2aGNlf7cL00RXG
0hF6OiY+oy4HZFGyLu4WYUtHQF4QT9JUzCI/dFGlnRb5ZOzL7PUqMuukxSuX9D5+
tUdgse1hnavJwB8WxrPCERcAMcMUA4jrO0TxIkDZ9eYJBDVhI5p3q2gXLAlTKfKH
TRGn9G+Dwe9KkxhPm0KsUo9fKjKW4IIuzO77nz90DfOLs6/b7s8IPLSv3vzErfDa
LgMLkdR91RlxnlZFHk0o/jaybBlQ16DALfjEwkET/bGau074CxyyxjiTUQ4lde+m
zLbUwt/mzlIKqkSjzM3ktQ==
`protect END_PROTECTED
