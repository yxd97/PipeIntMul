`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FzsBDAPnsuwJ7MTBiQfmT70aIfmY1gfXn8sATtDFTp4yBfSCDWMJFo1eYzjV7RH6
PH/0qK9XWF0I+rCv+WJT7M5AaN3vXIFrgqgLVaco0oTWh70Xz0RTgN0KrbMqS64O
UBYJSA0QPJbXhdRNRsGqc9lppkF4mp9zmMb7rtHJQnW7rWZMLjtG3Gsz5aZ0wP+k
mHBlLIg0UewLjPoXcourAqNPlHyBeBvntdBW6Z938k353N/crIzz4vg2UJujBW+A
qPJ6+dVbr4pbC7seJAgZnaC76R1Sd2jDrCFYXmjOAiotT8jzCmgrUqSKRDpLsOBx
2sdFh/Lzwkj0UyqYbi+pn2n7qFupWFkOfcNZ9TCZ27P+yJk3pU2cZx7Kl4s+9CDD
3oqKwA1RMvbcecR0F11r7OihYpG0W9NPZOeqigmXyaYtr5E+pui2eXJGtUMtfHki
fHFo/Bjwqchf8GureuY9ZW8hz0Kfd6yWoYvz4cNoOM+/ZHcKUmBovCLIKvq4rt53
IUutQwok9onnO9l3GoxoNVo5T74tD5zld3mGk8lAshZmLjNXzGIwckBYuw+45uEV
uUPM3foCmC1vAgfeOIoDZTd+z1nYHXcB386+co1PN7TVtemwJ1PSOYY9A/PRTsSY
BgpH5Hu3ixBFRt/OB+Bg7vmL0OXgwN5acXk3dlCkAGanYi8zk1jqQSTRBCxzgLP2
9/Us4qZqLzSCKnE+zsFt+DHNsQKKviM+LCcVp8e0+4dKvkTfxxnZPHUyomCZazyO
9EZktUGHh+1NVIwsz6k4FrDAXrSuWri/om5xeyijr+tAXstrBuh5LwlBj2hTQFK8
pEYlZJeQg5Fo3YHpDWRxKa0bhbCmGA1IyT2OZqkC/+Da+Rabws7HMJO2DYlyTeDv
WipSrLRWxqIzREWw8yspIRmgnSYgN8toSXsLaM9+Z8eLS0f3ksMwuCDR02EYOniC
SqmCTB925xtpI85OdnEU0sq0XWmLaWsRxpfuq33Mye+wh4rz9I5OWs+8kp8lkyts
EV80Y/0GNdubVwYpifkHr9mTVzz/dG8ce8GWjasoKXlTEI6kpu0IZ4bcavmDIgrF
yHVXDZtEdiJVeJfGmGTgh4X0vH4Zk74torAz81STYfKBYLrt/gmbNIvWUrNw1hS4
5Muu7RE+mJ6sALu2z6C1na4KYAujNjyGOY+yEESH8mBiB7Yj2GQEIDYulj+aTG/+
Db4oOlPeZ324iNhzhYifY64Gtsa1+yrN5Tdkr+SD93Qwzr7SKsAXg1al6BRqlK/0
TsKnM06g1NYtmE85Sh1dsTrtlLRaWs7MIhtwTRQjfxYvzjhOWQoiaPI8aJxL6l1a
9tn3uh0P+CLh6LdptlxSlTLDWe/pvxFqy+tWseHPa6lFzLoFECuDsjDxc07WZI3U
+WemJsJF6akvsvyNBBkcjgPk3Nj3BK0SR1mBWlEFOm9uR275mUp1pk4LEel7tH8d
558ZkNVA8HMhkEKvEFPxMjNWlXoFAT4c1grFRJz1M1Usgmubg7wTmW7K1BrHyEA5
pudm6AnG89dg8aZLGDM6dsznKg4eSJuf+07AnMoEXh8TE1d6q1w6hZcmXulmiyP+
txd+NBJVEgpXToncbMHZx9b2RG2W33E3cjGiIE7M/4vHAUs/ZvhRdaBU8e8+ycnv
J5eRAQ3wMhUvbHZEfD2nMsH0z225rkM8X1qsww2EGFtm1AV08wdTt0LPBkLjyerh
/CUhQOrkwbESlHYzd3jxbMUGrDwVLU6FFO+C9Gzy03nCi1JONkld+gwkUXe5tjK4
Wr5v2gsxnHzIxV9xzI3nb+nywoJgQy6qbPXI8cm6StD+BwFJZ43V7pJaeMqCfg51
q6GYZqtM+iWLvdnhGo5RPq0d+zPn18334nESodUY9wTlv/rp0eCWH+O5LkyA1jZ+
/MzaQpTa9M7ZHstHxep1jLoEd4VUWjjmonWJxZWd7LO3306Mm1ehGSKM43ZLaqqX
IEkkGuPnubPYixqrWJX9cyE9Ibo/UreYlxy/96MCPlrp4Lcqk/JXf34+mfX2gJhb
DzuVxmXTUtU2jdhmO1p/EKt8uVS2jpXg1U9CkDJ+xPtgiHtMQHxRAbU1Ew3UGIO9
uwQg9zBwm5BGmM2ALE3FaPfTu/KPKEa/JaP6nkyEX3StfrHWhepfknMVHTQqU9EJ
KwQOuUei1O/pHRxYzqPRLwoPUR1i3UGLcnSB9Gw+lXravuCdBU6NZBlKuBEzz6Kd
TM2gzzCjlKgMnxQN/9DtgA==
`protect END_PROTECTED
