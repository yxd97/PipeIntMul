`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGJUESOJLHeKWzbeLq7OVUF85lXJ1wFdi35Qxa4X4Ba/uwum8+W9gZx97JigYaIe
SzJtaua//mfIP2O9GHygmx4TADfGpjwHZnOwaiXMwiLtwFS/6U0sVU8G7Km1BOYH
0BL5wvkZ9FHhTZvfKtpMrAbcNr6J8X8Eacrs1VDEZvAUFXBA5jViVQ2zs19ribL6
6tEW8zIU9KgcPFxweH2TgMA1nG9Tm2M/ye+UrKDm189FhDKvP9RpC1OeGKvGV1BM
oXCUdoG5iyAsuAWBXqRQp3Kp3LFukXLQNOStllFYCki++IqdkzoEYBK6MATPG2fc
+9npoJVni4dvXLFm5j32Y5DiBsJqlDiVS4i5J4lUeIWiZ2a1NvpcsZeR8o746RVJ
SrTlu6qeW1JJQcuQjmT7gbTlyZ7GtMHcw/6b79aAphCMhF1XQDm6FktBA64qr3je
lJeu63qLqLmQ0vE9QPlZAawyODUrKJPoyt0c/e3XAwk=
`protect END_PROTECTED
