`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KPUhj3dAjdWaZbSJ7EDrZeEEvkEwwQAH2RACaQgsg7syIMpvINEBPs1SlUfr3FUS
viB6AlpClHG7whFX7QV36Zn9yv6CzW7TRf0fbSA3TJkclDVk43+1C+dz7DSQ5Dv3
rdZATBHGdQNWv1Yr6H6XDO6/hKvyYscYWXcNwG/soBXK2TvMa4Q49qgLUQKh+JbD
tjkE3U6YULzf5UYJvKVKlGAKnZ79nm1GuJyhsaYKn1JAU41RPxM1BMwzxywLtm6E
UEpFA+RFcfwcJaCpkM3xH39NNaKO0Ya+15QEDv42yHEZStw4COfyFXKDUyicLlsi
dPEhnpuWVLtEud/37kADoFZcglDlwLopE0y/u1wQbYMVofWxgBRSQBSdz5JX7JGk
0BeyQ5hRMjr8Yn4Xvysz7LJYhekujKg/M/OobUN5H19et7LzYsfLY7eQlN0inJ4P
wM7C1THtnkFvSPEg5+r6W5Wz+R1cLjIHwMJx1rU+fhwx7wYB2l1HuwX6biMC7iG3
g161sm0mFQOiusyOD6yiW9/r2O40+/oqhBAknV2hdx7EgHMYYMlacmQmhkK24iO8
cEf83R/Dns+kA7Xr2vmVrfEhfzMD+LPB9gDVyT3osywhbjMLY3LiL11aeQ5EiXI3
1JT21xDTEzMLN6xSCd2o1MpJvQRntJlm5mqw7ZhJT2X9rd9jr74265pGnYm4vBqw
PZW/I6Bc9OhEUBrWAGg74g==
`protect END_PROTECTED
