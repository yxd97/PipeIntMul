`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S5a42MaZ7j7m4l+gad0LXOYBbVcBjYEvNxUufl13cfZKdMy9JWjZOqyrO4rEKbbO
m3tShptNYy2NLkoWtgj1EFajDK/tB0GhtUrKMNyWOeDjMw+KbWt0X9uIICHIaGoW
1zyDafwJKmkBr4RdewSuCBp2GNIy3nctfbDyczynLPd9Dld128yX/I3WENs+opa2
OayadGw5WuRsUpe3bduZJq+TRUkQ7ENXUSfRnUrCFC8Hen3rHWF8sDIc0WSZ8GRq
WfUBctqLv+w/P73zXPfqn1VdOTlKhFFvN2ltPDUarwv/eXIsbvnPdVttMNMPJqEY
4KWRCcNxWe/TxkxtpMfutg==
`protect END_PROTECTED
