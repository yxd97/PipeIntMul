`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJzsnfGqosi841sJ8gDzlxzGgcmxnALEo1dTfwv3+hGLWsZ4SvWz7kv0th657B/d
M6u2f7BHcRtvWmdvJD+AV79ba9mQNPqgvVTG4L2tCdqUtPYyVcC+w0JDn/Uunldi
AfP2o+tehGOrMjjgDcBiIQBYXnYODxol6lBNvJmf0LFHJir0eFiCJS8czxAz+wQf
ODaTMiskWMF/9wNHW9EFVlN6XmpWinFyRDX/VbKFY9maiuNmB8CoJoy02I4T970d
BdwDUSPA5Pn7iaTXDZaisnt5oCIG8CiXG/aqohsoDJDXK/7+BBRdzKxV7Fhpk8mp
Edqy9tx+MDSjJQUmbi/dfpNn3Yc5Q3aX/6d1X27Fo5Uoss/9DFiYK5H4yqjAv6qI
vntktXy58GGTgdv6wZA6q5lCbLf/VSnNR9rhvutEock=
`protect END_PROTECTED
