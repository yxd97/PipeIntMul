`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m3cBfahriYRmLRCtetaKMlD6n+Ge3c0kCn4r/4Dn8ExNW6EQvMv366zvqgoNDmAg
9DB5E74mhd9KXujFqZaE+czrsnrb6baw/16gt8ee7p0UACPw2mCKOD/qOjMsaX74
El2lJ7bzT+36a2A6RN1nzraj7cFGvQyoGntmLgqkVW+nQ/uLgvNf5Av8Skge4wTt
aeXZ282o/lf11ClF8iAUJrajNbTmjgjEdkuZAnu41re0CdCAHQbdOcKZBJX50kdw
ym7eNMDszx/mB8QfMpCmQaXrOsp2AjC95QlcWYWM2pF77RsRH/Cqt67hQFlgfr7o
qhuj2YeiOQ3FYkC/24vmOA114TwHedGWGO1SP0zUlinwpN/BwHC0GAL5IAqkDqqq
lZAv4cH4R/4nI7Hj3gcE2f7ayVWzQw+FdoZMGjswYg9Lx4bLWz5oL+CVJtyTknO4
hsnPAYKZAwaCmokkOfmTVanIFx5F2oulhKBmBIHr7OaubaD9UoHc2WiKwb8EOw9N
TKNesb/GiMrS2p8BTEgVZhtGjCAwgMQE4WFhlIH7H3JcJof4c93B7R5fBSP0i3Xd
HU9FG0uJYTf6z9ygzNwSpmqVgjDLsruuXjy7wEDnknubNH4a9LOK5qevtD/s+VJx
eu2GUfNJibMXyQKG0+Z0BniBk05n5ZrVUBXvYbXmw+0Hga3K9zTlyc4JRYWBCSHd
RtgdpWK4hmPJOkcPiU6nMxICOFt1kD+LR1KB8c7kDYBggxNgCxrlt/A2GAiQHxtl
w5GQlyNDIsOD3PyfTEnsXvYshErw8I3I76/jAc0+6EzQ/PjweJ5x7kx120MxIJ/n
oKWTTNZ5S9u7rW/tT4mFr3UEtLthF3nDHWx0xboGIllyi618yri1N6oW27AYwEjf
dHtZ47K4Peqj7YMhmJ+32pRs9hD6Sgo2rD5hK414um4/AdoOI0XdW5LrdIw+waZQ
PaG/epGnr1wfFnrH/qbO6LHZD8htakXS6GKBJx53NKPcxGm7tlExo7BiVdlD3aR5
ac08YmVu6EoOVpTegLeeyo0D/0KkBt10axOcDuMgBZ4iOTx0Lex8QK8pGoWj0tBe
RjgIxQP+mzvvEJfQvN/LWC6qQp9rGIZRGsoTXv8so0y2P7BjYmpGalJuRDGv6/m9
jGSuq/74/s3Xe9JM0273rskvZt7usz7KkVTH+Ns/oJRKn3tPzZZCKucBXdUpVSdo
zmt5GXN6TpPFQB0NGmyj72PItY2SQSRFZlxqPikLmi9FY7Z9z/oFBPRLOGi/RFkI
jdlASfzmt0I913EWV8LK2DiL8FgW6zTovcwClP7nETmPao7FWMAEaSgqPTacgd/K
y2yOC7BZI2sPKHAZeDovNLCPLqgxpThhA4SSD7ny0FQ1DGi+yzuxYuc7bV2DRewb
HeaWoDXtpwRAd1HZyXK5sd5DK8vWggCQQ3CE+P9Y40SBgdoo//jSDBDOgMZTQEJV
IOLwhLKnQP+FFBXkp0Vt62XGvyvb2shG6NeyzjkG2g2RFTkihZXRWgn+7h285HnD
f6c2rFSRBOx83kUI/hmG2rAoTUiaKEQcQTw1v+GErnaeOVmrtdBq2JWhwdzPvbx0
`protect END_PROTECTED
