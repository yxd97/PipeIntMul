`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GwWDAcABk1tcypenCZsX+tNBcFY2D5wU2ZMojghaxjrLse0yjOG0S5qLJkEOgB1u
iRg8p5xEuQK5OcNIfPA8s6HScw1XSpOQaPFO/I5XGfWAtCYP/ZRZHnHTXBmCgshe
7BNstcCBA/0BVNIa/B7IXQ55h9bUm5Yeg3MZe+n4w7DRuZkzufGqWeChQbFwWH4r
f9VnzZBQXD9hwS1oaMhevzfd98hcaaMGnvmZdj/eCAqQoMlabfZ7FJg4D0/c2ctt
uY/Jn755pnZxGWgB/VpvpZmgm2C3CzSaLYZUa56Q9DkzpwvxK91xbwt0Oa1MYF1F
dpq0wC9UEYiWyJCNYIFfl6YPVB/ETYme05+2t3ksKmiY98oqrOoZovlkek2So32U
dlc7k2yY8iwKVQobv3AAy10Op5ko7mzs6HjD2X8cA5M74Bo0/AfWvAmCN0qmvQSP
`protect END_PROTECTED
