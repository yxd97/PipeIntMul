`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gd1EKcNWuROqnvh008QKl20ni5C/VVdgtaf6EluWdlV/pavIr9bjSiUyqYJZLQyB
bRruV+sbacZGQWzc4URdrlH80heAhnLf7EXptmZzBKTEfNL+/1O41bkHK8ECvKm9
8O/DfQ7LosoMXFMGgv9SMHS94ajergQ8wQeFZJny0VCDHUDLMwRdjMkUjxw0UfP+
d4FvCLDgXViWps/O3b2BWGrL/+t6492j2thsI6u3byaTXBoG+Zn6WXDBxFuUgysZ
g5t6XmFcbEjlwb/RYkwAuAyQ39laaT0Q2AjhCyFhlb6N64Twl7FeGSyE0uYZuYbK
y/sESPbfKUooeyyx8G7T2QT8fAdDYMN8jyiPCLN1V/a+ayf/jkY8jkDeRtcO5j9J
ze5L3Jvvpsw+/fcZIJ05fQ==
`protect END_PROTECTED
