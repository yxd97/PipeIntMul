`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZWuFhjiRimFuhQDk6lRFnNNPrcnOxm3xo9j8sJhkSjtyb5sOZzBmsmggbZJdUww
OK4H0BxJOmTFzhaHBX00XeSonZtHTT8uRtEg1pEpu8eCDxar2V7pQYDKmpgyVXX5
TyJ03Pvz4AO8c3bdbIK+4U602kTzeX359Y1EF/gHbdKYAQLFm0UqBda/YrYgwtdM
nwU3FEgtDlyrcteDRcoUjMbRBtQltM6XZN1npSXHJLB9iEEH57NzfYLnQdKDMtCo
wZFXTMk4fxFl22vmL5OwOqecvgaIXs70i9Mixg7z006NLindsGbLYNA7Rj6FRqZ7
ogTXpWSvkfVc2+/41psCh81BFcdYeTbGbcPDNWRro0D9KCe8SSxi6lLTayCuiGl1
whw0fxKXRwqqPVOOFqpsl7T0PyyfkCJVQhq+4U5IsZBpRUuIJihRCB4WkHxE6T7r
IKoB0+X7kbjK6G/GcurXRxOVgQL26DRvtFTZuwrNDXM=
`protect END_PROTECTED
