`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1E3Evrur9UeDs1adqxN/H8qadb91TRAWj0rY/HwTM+hjdrG7YzugYcbF6A6+VX0j
cNs4gnY9QBknr2MdTVuHvIlu1N+6VxMLgepspg9xq0+H8qFfADGFhomYRECn6nZt
5SWqMxmsYUfpB/tV9nimn8xiDII8h2VQETtRHLQX6PMyZgWstuDevINIcduBwgtr
C5wAtuZHzfBS+P9cMuaklULkOX0XVPeI1hZReqBewE7xpoQr6hDMWdTXyTJl/FK2
nQnlq2rei40EBhcWXbRagBC7rKZ32TW5JqqL3rTrzuSAIGTDmayTd+si6H/hKzc4
/CWfrwWBpcUqWFj36g7/VzKMwpc45/0jv5I7wqAv4tEqV3Bie+sfsnC3ZJhQla4i
e18UevpDfAMV30LKejDVTg==
`protect END_PROTECTED
