`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zH3pk/0+Rkp7lsfIwcJqAAMJCTUcsUtzJmtt/+eWXfKFC2KSZtK0HTu4S2B6STGe
nRnZkzHjNSzZ8nR/EJwzCV7gvtBdpVuZfeDIMemgEvG2NMVup77hkf+XuNNA+t9u
G4g9r/8hqnTiosPJbdPz8NQJKfhNWCY2yuTe/nQp0yfryQQNeEYoyKRNPktOgJ7z
3oWRWuCwdacWo7htL6a4pMs7/elufqupzfJbuUWYgnLX4S3hjlhnEWDDYN34Cp0b
KkM45YSQoZFL1C9Mc5R/MBR9P3ye2b7JofQhQbiNgyd/lI/Aqvf6x9DaRTCbkm8j
bwdfufzhF/CL/0RlHynwSNyKxVX+eB8IWd4Gp07lFe/nWLdTv4RW8KciHi5LbUy0
mLvfUtA0CZt76Dj2HHzH4iXRztM6sd2KdNXOhJ/8hS1dmSYOiwqZW1Y1sjSiX2Fx
bw7bQ6GkLN2QYoi0rW1/itzj3pqbN0S/fRH48HE7h+xAvIfjgNrx43YUNiNQAFd6
PHSYPhyNALIK1402glXEU1vpEpswgFXGlCKbhvvFIlH8OUh9Gw0Izk9/2SMXEpwu
lpr5JaV5hDf9lwFIrHXljPJXK7PkNLwgkfkttPsvsTMSWG1s7zf0jpkPagrvBcvQ
t7f8ERc+3l28lE7C52HPH/EZM1a/+0T2iiww56EnsTlF6ER1fTo7X3/BZonbNAWR
AqYq3dBTj0X5636x871CmV6icO9ZSd3IurKf8ykZBaIMnhW/CynT/1k7F3kTrCvT
Dtx42M/4MOciiK1PQPCE1QeMzjTfhNformOqJlSLiwxIO5yrMLKOGiBYwVaJoYKs
FbLaMvjSKHZUnOodJYfzXPuJvRD4UIDiH3sMYhAr19gCUMxNk3EVGLjS2g4vV6EL
SDv7/U4aFfCatGUqPiIgEtpuNcwxLrL9ohy0ePogq2FTLTSKUIpvO/3T6k7KaH3L
RaEA9YO/5huc3RfaFpiSxaWJEhblh/NtVRLayUTPmM3OemxM3o4/E7ePvRKTWpoq
pgkj4G9VHti76SCW2IjRUA==
`protect END_PROTECTED
