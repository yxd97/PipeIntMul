`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p3ip6KE0SWj3NrOsNzCjV7zvNm/kbI1GGajCkn12WkHMcE1Kn9/UR5VIhvKUXGFn
uL8D0zvHjCCv2DE0kyxZ+O0Sx5U8No7P8cla95XW15xEie5Cb2lDSnEZfR1hs7K1
zXcPkfOLqwCZ9rolxlJOnJW89cVH4R+frqrx7s6j8l43Ta9o6XaK8oMDZTPoSGyj
wAB8j3LasrEzhiZaJbdm8Scn6tqw+n9LEOMGaS2ntf0qRLab0+A5di0rXebZu5ae
p37cOk7mzRbc5XZYZjjQ0d4u0/7sg7LvnxUXhsdKQC2kY2as+lcGiPioS2JLVQe+
r19EpcczF+hxXy5/whnsJlZNSUqfRLa1OejR+BK63Ijbqx4d2jho6ABltoGCWx8H
KW2MYwty4CE9XX8Wapg02O58nwpPXe2rjhY+SyqX+dI/M1DKHoIz04SDwWf4ElpZ
wwsQwQF9Ci2pfw6ds4Vj228W5Chm1xON0PWWYBv1lh5RbYjk9mmmoOmUdvliJb3v
qn1CXsn8dHdYUPTAdN68/bu7ceLGE8Mu5SY2CWxKiAUppHyiWXr8BpC87I9nTppA
oz6EN61x2LiagMbaxE77gyKhkQX0bY0K6qMKGNuynGxOrFJR1F88IbZ7WOuqA6L/
zNL2LPVWbMNlqJwgeJ8/WDKjKOXvqbw/gPvAtFlbzAz0A0HUXek07gow8horBWSC
O7XO2T2IdyYHSoG2axe3ZX6D/Ynd4GOGRCjy8hv0ClRys+hOoZMiNXzQo+vXpYyH
sx+4eEAamRMQE2E6VeX1G3AquC+TMi73IJsBnq9ML1wmWulHyU8SSRcoVdt8QWNW
mKGjuYdKI2wCWaARdfbMOTRJP3lABm3gcPJsGjHL7mcU3DoUwJtj4WiaG8vxO5fN
ND6/I8po3cmt4fCkVyfexqNrBpjG0gsPV0VEdShqzN+/00z3ouYWh1EJSS4RieUU
6T6yNlMN2eLopnPEzNJ9cCwfOh6ImtLrjlA8qvTRIP5yxXtyCR+spMnyCU8Ytg/r
5Sa/ubg8ZkkktE+ps0RMKGcoZ49lz5FTpShULrWXEB3Dx6xJTraVbVaDe6d7Mm9B
Ly3wrqr7yzU8iOxoYSauuOOq31zfQIca9N+lob+IiPA6idY/Gn7x3OXPvOai2s4r
eL9rHvnXOkiq16/gkk3/gKMiC4hy1m8PlbenIfPhRhh6brQ+EwTcaflfoFhTgviS
e2vZ8m6WEOBKyQudhfnf+dNPAoQjxHdq/IE9xvqkgCW0hHxjQf7IJyoS/QgKne0K
tav3rSNpnVi4xz5zwZ48rHBKB7YNR83IHvLcuJQ8WSQ3Gt6FJTyxzeJeMHH5H3PC
b3QZjpDN12Z3Nxa2apSDsnhTxL4AQxw7FU5//7tdu46vFpOYMs3WMdamfFXI+bzS
QcRE/wxRNzPSq8k2eKNeYNJwkN5CfHF+yhoe3+tJaXlQHeqIuSp1GlWHoQ61aq1E
Hum7SicPSe3DP1YheF8TWb1CGHBQeY9hu5cu3xeZWQXxPb6VBiFWuu2Ktu+THnC8
aIxOCU1OUpqMO9y8mzVHZCT0aJDgBAAUfyZCX2DUtnFs8BAENwPprjVMBm0kpLeH
3TEPlzhPwyZdGguNB1x1fr67xf9JsjE0RV6lIivxufgK9KUVoUipPEGzlWgUYd5i
tRG9Eb44L58JjBVJzHiGjnwI+T4SjQAJSwIAsmaZUwNWqLMdw7s199jTLYI0vgmv
xg3Sl/5t7Tvr31w4dSVEyzJwVKwv3MNie1rmYJEpbpufKg5CnQ8Eydjdjn2C8fDY
ZpycGIvOaH9ZrxlpLK2SkLq6/OgqxIHhDwXZxBqRA2ISmg1eQFK9O+j6l3sqmEe+
vggr/wmE15jC1dehZYLKXl5uHfhkwE/in6xXBCRuykot2m0APysW8ERYvdGLFFzz
dwTz9m4Hprxg/lAIbJ6UkY73qRCky/UMIr591sLpDAWQx5T0KKUboK0zBEpwoj6Y
5Q+v66DTYTJPefG74WBw+IviynzzRQYa+5CZ190fjEV/Os9b8jkuU46tyrEh8czZ
7Q0DqgGGteFR5l7UyUtQ79YsWmUgEizen/1axnoopJhzWPuDhJ8ZHhzXfwp7DKVs
jp6mSjqIeLM5TfvSxrKUrk3PvNEwQcr8JeNpgQLf53ys3FLQ0mtBD9H1hKiUhoXg
FYRE0kw7cJztRcxW2nk0t5TqiFjCCgaH29CXD3n1iGCBF/WeFqr9rVkjwG6A2mbU
gPOOemgz4DM7qA+YOvSfKADMn3yAoIy4ypU2ejQGeJ4VedeR/87Pd85qSlE69c7y
Irs/XYdB99v9H1fqhZz+G13gUlTX0Le1vcXvCX9AmV67esUGMRTkRZg4SiI7S+nF
NoR22pJdeov+OKo9mOuPs7UAxih+y4h6W9qGaUCLHK8Ne5P05hLQGWNKrWs7IAJg
evKA0dmKGaJbdLvCu3rB2+AvyDTu2BJjgm73b3irAdkXa9LfvWATzTfGUiKGpHb1
I0PjUJ/XgSpITKs9Ow2Ox+/05gDv2laohSckxe/8yttsg2EY3JSQ0+xtg5nnR49d
5v0H5Vhy9dsA9gqF9I+oo4LjdNdGEc0hqovW7kYtxqrHvIUoQr8koIVXbiTPbvnP
QJeXKlJgcPZjhVkz3fiiUV6T3K21ytJ99OAWTsRq8l9U6nbBqnwdRknIRz161MKI
7wBSXR58kSYtEGGE11NgfW4ckdet1mZ79PU5IpdOUXZUxWKeT33vDDbUrRgjIKjN
Zimc9LPqXt8zq6MG6BCMDm95u+oXEyMlsOa0yVeBeNU7mItEC9nA19K7YZq1BVg7
LLIkWSi3ovzfd0cDAU6Ri5Qb6W3nkxFC5Ad2u5M2gzdvNY2c8BFf5tNDC+IQ/Y65
Nu1w3DcKRycQHzif6egXWPg1UTZCHl3YBO3w28Kv5x4eEoSSBwiVrsG0PBUY+RLP
gWAnVf36V7b/cC8YULQe/O6rAZux6No+3gcAqYH4u/BNG/zdBz5pftwg/yb4Mbd5
x6rgJpS3e90gvp6GGyGgrMa6VGpXUNjVBXr02jCUGaecnJa5q1Rc91/6bEDj+KK4
U912ANta04+wQUNeDQtwccWFWuIW7vvO8JAQKIQX6IoqOnJ0CXs4rgLIqgP3OHDh
/QI8+q83LJZkF+1N8iNc9u0awM8DcMDpnhxoMoW8a/gGzvH+06kqsPChNXi9REA6
0MA7UJQDkX7k2T77RTURkPffmSZbhM493W0xRBAdr/N4x2ZYoLxei28mHZswbZXB
nzGkyCm2s2aIq6kUDfGYBLZa85SaSwK2qZ8AfU1X07avMlz5gGRSCwYpFXZik/eI
aY/CaUqjfCIx4QfdJ+d5y/MKRFtyHqwGXLrwmcgkeUpTJ4HCTlk/CRHjUcw5YiP2
oMD6qjGhH0FuKTKVum5J1Z4NOyT06iLVntWz8wpLSk73sbft3JHSP+RKezEge2Ou
3UcSL+18DKdSfEaEixqLHgVqILv1MeO30qz/iAmMPblmeBlY9m9QLtqk8ATrX3Re
HMUMWgH6HckOIZbCuDUJU9kHL4+RBnGC8E8d6z/YvUN+vMuqnop991E5Jr3TvM+S
N+jnsqGz9kDy9w45vvG95nWITevBVGamqXpSnXcN8bPBc/dmVo9gZbwHdIcr3fp0
8VR7mxJkSNSy7sz0Q1iwzX1Mc3FuOWQxsy7cBKnIAQUPtMkXQRgfa6rgkXQ6vQDw
tUbQAy6Hk+WS8VzUnFaGeI4mPy1auYRIlk806/gqYBYM4KclFwSECwMclVQqHhUL
refgoVWJ0ZGw4kuFwKX/YlbwMLA1VXtmWHdk6SZ6XvPDs27itdAj5j7gYbK1XCMO
sLFNoLq2yKKD7SieEZ1FyEbzpO1ENtjn/MLQsqXHu7WNmEWvWVzUeBUmhqaMCHzC
NpPm2K3kD/AphfqRwKZBP/wIx0YZIkw0bgfWDL9jG6Ov5h3m4oR4ZKLz1GJBC76L
D7PvFBpUa3j/GVyuNb0cH36OGCSFdopoUItBdYG5O9J8sb5v+X9VQRZsUpVNtmex
BYm2j78py+Xmz6Obbq815oaQyJPsDgPM3QaNg/OboarpeGP4xOt3XTArNad87TC+
mvJM7waeD30RDCBeqZRMOlStd97ZCNf6+IfWimvQYh8Hto2RL6Yuq0R0eNNInRV7
wkQnBo/FTzlZiaIfpjwdJY6XqqJ8bzTWdaVSAW62++hz2iQoV2GeWXfa7+bMZuBk
10skimi1hSL0XE3WklUoTAm65HW2Q1a7puW9b9nctYfTO8tYHkz1im/yayjFGkdh
glBSdwwagi78LXgDaJFUhUuzvazmUCb+X50Ne+TUB3XGYHkVOAMnD0qK9xNU5hJz
MyqhWY7GlX6Rg/heyVUjnWf6DzX1rIh1XV7oFlJ2heMN5qJYomwqLaMpY1VFlA04
ljSsJLF0kpBgf2nIeBbrkYAKcNr1yx0u0vH8qKyq+PZWAB+MND5BBJxHnlOoRkin
GSRHWWI8RXDlDj/yN2JNZChuwb8UvXNpXAE7gCXlDfLFVxELuX21qpGRanSJYqOn
Mh/RrLqbx9n/RXDh0J27l24ziMCuE90j6OovqbClNgVppXNaurLRtWAeOIQ8Dqmp
n2DyV0mi2YKVUY/z5XeRU8/QNc1AJaExUjK8OGMaXMX+xX/6zgKvqD9G0ddzI7hF
6anTuDz3A4Jq1ZHfAGhz2RkK77CaG70jXaUrdBLQReRFZmy/N5YfyzSaDWsntR8E
8Penc4B4swi7lMuDffzaLkTiN2ofLoPQSH4aF1IYCMRnzcujRpZuuLlmAtw/gVuy
+FldDP/emB51awqvRUigdYolagj5ndYJ/3BuvMD+rXmkR1d2pdQb9+w5I1wL/8Ny
l8kC4ULzlyJbgoqnPWVErOi27bi0aoWxqTDrViU6810msiD8kpSQWV3sdRswaFsp
TB+kiSpSqB55eEfts419ejKSMlfUlQoi3jx+QXMnQOlnLfIIgjW9cL0aNlMzhO+s
ylSXKHKu+AX/8Dwjd/8O/K+i6dpOmMFXvUuhj8MME5Sx42RtrkWLRNTi98+VJGOc
zSmenKcJ2t1yG2ChXTNWSzGtaagQA4dBWtaQp1xYb0JBuU8L42gHAY0BexDGSYpY
g2orLku1UjconOSrfFDUYpcJtK6i94FXycMStdrzvtMmtTQHI7cltQAqh81T0HQ4
CD/xzLJY7YI1ZdWnO5kjWVc2UJwMqWX+kBTuG/mVh5qlLr5Fl6yy7CPKjiL5OyUr
nQwTuibB7c5OHuprzjt8d8+W5dpDNtHaCuXl3RIgst8/qRPSaVxKj0iiO1CEU9n6
qp5RWWhgB5jrU86tuAkSml0RpVG65ilNgyTVUuUiUNkQGCgaDumvz7W08V1M8WR6
jCYKQ03MYrTbH02nVuZM3lvdqLuGjNgvJOtlPovd6L9I822d5QHZVWm350eP7Xrw
bIEuqS99f2GJL3uIdyj2NBhalZlaUgMB1SR4BnsS3E9qZfU7TgglSo7U7ZMp9EiS
tkUW/WxV8HOoQ2tVf1/DqU3BmtIHmcrp5DVEpd1nHLVaapd+3BBOncia9vCp58OB
aubcVDMhur+EmL3HBioXdZcP66Op/JdS8JissnjXNI6iUpwF+kUAkWMo66JiuAPV
A5eiXUfnpSDm8avkc+KEWTeS/fxks5juXGhSaBJgCPIvlP5i8/vCssCXdbTFwasH
0GZQf9YJlEYUa3wmc/R00k0hZbNVPTtWFUNDCXqkEU/29EpBQt6sPlFb1YLUIGuA
81Q2xKERKy07LR6HfMqJWs7OGfM3iIgjhXOyj7oiGX2Vgl/XdWlWZcWQVc+txxa+
UAdN2nP81fb+0al/a1fQGM5CpRSjhaVGTAgete/+PvlQM6gmWQOsh0QkszFhCuN0
v/iScpZRbNqkrUW8CIspgXlFEUHKYSEo5J2SyeaHk9n5C3Pd45NWvEzqDp+UzHZv
W4xPpTUup9k5hsjwILinuHp4U1Z8pwb+aoa8cEy9phu4JY7H2Favz4kws5cRxth3
f34ELpX8OgG9yj12fa1Ixo++7Ebevlxib7SaxKJUgLdPf3tqW5tdtlvk8a2omg01
S4m7xwTlPDHaRGwbd1GKhq01oVevsAMirLRwpxwJKDBp+OBYZ0Bi8Jwbvwz0s2jn
hG+QSpENBZyr+ANqcb0RkfqP5sKuZzPdqPBda6QHYbRJmwpIzcOAOQ8c0FzubSHM
IiYeME8aXD/UUl36hMSfEaju9yIwdrLjnDnzpRk+XD4b0jxa+mbBAINeWjYRxmzd
iv2s2RK3emKvGS7TkYZrYgoFAFVq4YGxyVBBIMek1senuhspjiir3iKuZKxYaZ2r
+KDZ3mzarC3uec4y0DpWenfqhFjmbjA7yQ3sTHdOasoVq1fsw1epc9FW5ZBtB4cZ
j8qSC+8ac34Dpf7/02AXyq9k3i+KvX2y554NEtdvbdPXrIhcgSAO6ITK76WJBiHj
3idIKIaz/iju0cCiFyOtHamqYLUI2agCzcTToesWZXL4dohz+UPQ9qGBeetZKw5T
s+jwUHc+uN1Q9UrNWT+s/aMtVuVzYcG6/cg+8HOscKk=
`protect END_PROTECTED
