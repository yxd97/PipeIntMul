`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V55e2Vsip0lJRC3LP1eoyNd9+ZmAlSWLW2jtNpdj1yHPpNqxqBWqbiY+3ADff6LK
fc8rvQC68nduWRFIRgQkNVTe8f8JoKVL+KJ+e057PtGdRMu2cKs72t2vKNlzywdu
txonBvbSdtIPLGKe0cUsIkwPTYWXt09FkKjE+fKn3kVkXsCrfHJt5n0ohJKufuM8
YJRJKrnFkvy9edi8iQMiaGM6XyaWQ+jKHbZ2FsISQrvl96W2l0wRQHWglJRNqGQe
Iha994V+34E6qEkEzCIVqZ927l1ipG1aM0j7SoUcrnHihwHElDHGEE2TfVhX0hRs
bMrDm6UEFDtwz33060W0JCyXc8/Q4JzGlOocc/Vhvuuhe0subCQPCuX5ev6Zefbm
frx4b5G1Y9/7FnkX9wgnFuNpxZ+hvqsAjpJa26eiKf6F7vA9tdM4H+A/gn5/9ngr
yUllRVw4tvP0Fj9K22I6VE+LMif6EX496b37H1W7ZyIl06WkbR0+JbHhWeMSyp/n
rUxDHOAi1B+bTF9CPoilqRrHnRMHuza9xpnOZP/3zxKLAzQCax1JKRAy7L7F7mJC
Yf76M9tLQ3/mgJ1ixr7qRc2BY9/+ar6TG4ZaPMR66AQY9/28BeaiZ36psTAHOI6A
+al54+8E3LRHsTdl0xTIbzhE6P+FeDGDNznw8wIfAYMaoOg0n3zkz8qjU5KEHXVN
aPeD4JxxD88L25iNFHafPK1skzP8w43d9vVcYC5SkM4zAgdj4PGyucQyva+CCv6B
yeg+Gnj7vRUrZEf5oLwL7rUiXZ6G7sGesLHO+89Br4Tu1m4NhslgusXwSwZnvjZr
gwmLnnrgzJOgf5IkSfvt3QghLba/lJlOna0orWjM5uA6HR/CGq58v2d3mOj50AGB
TKUrW1zzoJwSANBvxqQFbp3FwGHypLEzTRxPDqsMPe0Z/Em3AHUuyVeI7zMxCMhy
L0v3QN0C19Mo13GtLUt6IQn2B2SimMqvabFtepGEraYIePIOpPRYBixFH6/LbuIw
YfIm8/c/252IS+PEUGWfpmwAhjwGnY/1nQk+tQmctDcqJSDLcwZ8eA65ExMquHNr
6d2kdxY1UZfW9EMSuvLItm3qk8N6cBvqhaRo5t77hMDkEbb8TsxqDfVn8ge43VAn
xtbB/DoG9XHPvomZsr8zRdONuIRHU9K3fC+FZUGUnSivSUJ0gLRCOy84tSAZVnw4
ox6aq0ihzvCpARXHDhguHh6fZs3YxqAbOs7ZskAT+uGN/uhwMFWmIX8b//6v38t3
R2sgQWBI2hLNKIVD0LJOaTnvndt+vc0qK5eGjFJJdAacpDC8B3V6WJHfZFmMb2Lm
y93s5GjzRn+RTYdovBNKB1BEfSHDMW+uAstWYtp8xEDHxep4WIZsoTUUkvPnxR38
5z106ByJ8hJ8or+57fE8maD0fEub2M6fLApVDuNFN+AaA9wqfVdIQmiZMFKAj8d7
Tv/SOJUaliOuPHxQIxgA8JvopbdqpSfk2Y5Ccfi0vkYL0MqaoYK4DsiR84HfXaUA
YGL/+id133el4avvkNAxqmYvQJYN1pNzYn/XTwSsRygWqU/fLOdi41tndu6ONkGm
2lREa2f6xMq69dshExVR7M45R1dpv/vq5Y+27BLC0OPePPeBBqfP6U72YwgRl2bb
JRj+bADBoZB7JzpzZFVIQLB3fCe8F5F2wMZGQE3RJzXpYWJnYx/rj7bcZ96ntJlG
ga3EDQh62/H3lRtx3NkrW//tJdTQdHCCIKSXb0cW/6sJZPI+CV4/lbOeHUkK1E59
vSxEvGPov+m7K3IV2UdtfhQtqyGBfw/wUYNwz++SFQzy47kF2wypMCsT9OZy/GoA
II3HHyDcLoVpTKIUiyRLum5gbwmOJs1Ecb4UXhX9ZS0G6d9MqWD0WXCcV99+NF6+
G2uLh8pjFmcb3Jr/ZwC6VyiUFBSVT7y6bWcz6WsI9b6Mg/T9B7RxKFhwYysMcf1M
VCWkIvcaTgVLZXDA0/LoKdTnszIrcRU+4mfHDExqhrwv9ZZvQqp2bYcqi7EbNLYS
td38HeXf1FMHfjaOXe66npeKm0zVcCZAoMMVBZ8hRAsQKc2Liv4KBIG6TwVthzxo
dmwm8/5/4FIOPoA8Q9dIrU2l8/fVJxbM+4LwWVmhAEoG6FSOerEXEWtHuq4MzmvL
d38BNibZ+5j002phxu+fa/nX+8rr75wK29EGyzyv2KrmDCNn1U3VCEK3ApkHclH/
SKQaRubub/SDvGOVxzOF5t6KoPllpkzmlZlZwjt/pUtUbj8Z8BCOPplVwrSMwpb6
DYPTNXRs0M7WW6+Or5Ltof/ZYkFSP0dPc2c70K0i6IReqs9sVXM3QyFBujK1yGjG
Zl7Qe/dO+XQYo91+MkTLl7FOUHnUHhQbWjPvoiCFQtvVwGKw/KVmudLzrBylgC+p
MfLefovkAaHp9plT3wLdSKhF6dIQhEm0v8+hv6gOvz0syBq8ukeZZC0aaR45NFxi
lvmwuROfhk3fQ8zgfrWZh/jCr4k0mekF56xK9lYOIiiPMwbuYyqdOyuCAHWvVeed
ZHlSu7ecSa/KSHnANxEeZL3iEUQuiFOBrXPM+ZkvX/87poycNxvKQxzyYpz3FHhB
4a44RPsAZKEPEP7ejsVFA5Sf5Eswjfg9QkYsQwgwsTcglj1X7FE41errCJ7xP1td
L59Ty2t9g8I/ZQgQhXDuIw==
`protect END_PROTECTED
