`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/Qy8qYCc2DfjIGPEK1jFI5WE6MJIMnSbL0j6+H8ZRVBjXmfVzmV/9gYUGNzDTYi
KC3SM+mWEKsw6/bmUW7obTURrSSPBKXQ6aAdRmvAaYwkknabbJnoqpMqwOxYCfja
3hF5Se24A+TAm1fZfOv5o5jyjR8r27E77pt0BEdVa+umfSl81airlXtFW9nLlQAh
UgzrlIW7heqvlpf6OdAi0zDpbet1E/7t3Zcv5Xt7cysSDt7mkklOk7bPj/kHVdG8
6UVYVaQK98bWqKw4R0Ao2eJWYOc6x4NJzvI8bkdpTHo1UNotlPR9Q/VM3KRY4sO+
i0fpstxpVDS0WDITEI/UsSX985kHeH/YFIhlIDARidsfe91kqICJuL4RrbBdEz5a
W9FHjJ1x5ELtxN7Jnxp4228uvLb96hCQ4a6pKMEuhXmUa1NmzqL6SHSqL4rwfCEp
MME/+YRrgt6cwnarVjGcKnTteeJS9zL2HxhxD69AIpi0ngevL2oHIjGq29nRf/0C
mMeNQHxvXvtn82hFrAvPF1VAg1D/2UFqG9UsDpSu30jA0WKQlIV3MNzYiHtRFNft
8KuUmSKFzy10tBmkt1cuQ/jvcHj2AiRj1XCDMP7zXmaebIOVX3F3Gl2IuXq31ObZ
pCQFl5mc6NJSVMW4C0Al4FAQ9+LY2dfT3EYgTY4rHnKLXyrmg1bdJs5zaDdPtcTX
PND17sMeD1hQLv7J4DnB+LWdpBW3RLj8NjNMDzkWAAWWJiPsGlufIOujnGfqyFjo
QVxLPflqDqPWkbuTXcs2l1vdwDrSI4AVoZxNYQsQuI+UPG198voIb5BEvAxHBcce
1GyC+xCBy1xebFBVnRAIS527gNxn3YudoC7d/POerBmbbI0TZ6ibcbXTJZIxUGI8
zBZui216FGa7yhiF+97Uff2DOdWZkG2GvDuF7GOxYUqDkh7Lm+riYYg/ICUnkg5v
AEY7gscqx78qC223P9sAIDiG74BeKIJzhtdAhDbeA7QLc1JcLJj/i/+BkJtLgCh6
x+69xmp7nEFbwkDJT+XnpO6wLOrJcs2wEFI/QpiiMfgqAe8hgi9brXgTfJSxYB7w
5Ritw5rEdAmmSj4RMurXQXeoJtYVReWuNZWikxEvhTWNdz5Z5oXZCft4dox1zwoN
4WjflhHu5J5N1yOWaO3Q8yX3Z0se6WV/PnT4sq3tX+TP/JQ6W74Fb4EIPprgy3RL
4JPqZwnC5sRguq/S6W1JSfnt8Hbfpwxod9tdmeP3l3c8JkZ8imivaRC7OKQcqqVW
dB2IOxFs1GWd82B7WWNGI7mHVClVdu6DZxayE/YbNkBm9BrDiJBKL7pTNSQO0oJE
o25cC/Z+a3hWROod63V4rt0b1dKZH6T02wQkxXlYnEQLuYpGF+/yeAMy4F0QPDLM
h5s3n2UWRB91gLrEWSPH7GRr6rbjuxkkQO6Z7+//puacNzKyj/gzJ49stumz8nGJ
9pd9QAsv0XX9jYmibd+R7uRTox1JMhunIuGZf1+h7aSCBWAQJmPBnVXjmIPMzY66
seKOHxkpsm27uhO0kAjI7V+Ya4ZspbyO/lokyXjrsGE+xsorevtI6sACwIzeBor2
O35radOcdTkkF2oLJs7LtDhfV5pEq/T6MeciOw58e4bmSguh1zY+xXBPGDwQscMG
1I0/YryUscqk8GhcU6hgQqIxPptqbAb1QFXAMoOYiYo+R5X0KHgLz3Q9V7GgxvGS
WJD/rA6GIvLVfK/dRjGi9w0Dd7wk6K5Gna5kvz+J2ajq25czkdwbqCRracbJUfQj
yLOHlOHkbjCqOiYKWkN4DnhrYh7CGATZU0iULJ9p82/+oouVq89lw078laXwWbRJ
t/1IDID8tQNuDp386cQiE3xpVYSkk8gITQuBGn5glP5BSGf7ZrYFZaWZ5rfoZcbD
uJYTIMC9GRonFoC1ShESXS8FuOeV+zqQhLucB/6+sb/j6PtBDBn07xFDsf/sl18M
1HwCqxwS/DhVUiCMPq8AidRCR/W+OEKlhAUue4E8hP4pTz7qbEOP5hAGn042tsGz
9KqG3Vau5xb44YtOZ3OKrYrCDVX4cOAg8cLcLM9Ig0ySPJmsiL5WXn6zL1krYiMa
uGWQwG2QzBzZ9jH4w6oRcZWqz4Ori1Xy0IawZfpqaX7+KdxUvpjGwRMkSUsjSg7U
0LTLrwLupeKYBIZ9Ot8pkzjjyFYw3U3AhxaDICzYVWru2bSydSO2k3pp5x3ssIq4
YaD8WEBc86PhX0KNMtU+FqJ30aZk9Rt5sLkV9n7PGKAVYKeZxgfxTEynScafZZ4b
Oea5ThbezFg/WrbXT9OWRnplYOjOpKxhQtrhY1lCBNbYct39fTuGhABKEVXSIp8m
pJ4H3qU9JYbv2p6j3aGSU4Rf8L1kUnBrRjXCC7xh52ux61KT8v47aDhW5BWY8qxs
KpRkvkHPNQHVk7/hiSxpApdOhBiA2tgTojJ1Qbnju6iUEdCczwbIsArWGG8BepQr
UzTdZ1A2LfuC6Z7AleBDcuhUFeTGsGgvKm7z5ie6XzkjicDT2tJkStOsCEXXGlMz
VCEGu83FV7oCPvqgd56EX6hu9PTcZPkqmc/Gov2TQJQMm3OuQveMRrf6VgEfwLIU
mNBfHwc6pPKdRtYxU5rqnDJ/ilrEPSFAeyLQwqYzcP8ue6msEUc/w8W0WOIBQES9
CVy0pxOc3/9LRxhaK9HuH/POiQgUgeU33/dOaB8Ch+kGMcIAdGxtIe5pXxTj/d2a
aHNYbrsBoJTL7s2+UzTbni7wy2cVcx4v7qlS5ET1Myn5kxPNE7bYDC0GvProYF10
4WttKHNV88hhVmwtH0dZSMCfk66ztrDlwpresmfJtxBvCiUibW6Za8VGFH99972m
+NE4nQ4lbquMNH8I6F6CLZi0mute7MU9VMl053G0QNnuOD3+NrqSRzKb2zSXcU/7
eoegTIJOspgjpL/CG/USs65Wuj+JT3HcvqTJ6v8bUOe+xh/UarQza19Xk15h7P1V
1qewrIC9ZbzNMDCwDifQAj2/LlN7zB2g56/2s4wyl+3GBLPSnIjL00G3TEtleHoG
V/efAA8Hwp/pfjGOe3LCnL7RYWys5ZGfNr/LjtLVFGJLlm2DjQjL3gIaYdRlj1UP
fWcaODDmIyla1VlB8iyw9Qur9aV+yq3epIxHNkCTe8U=
`protect END_PROTECTED
