`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zPKtrLdPrGzfFTLW9r/cdObI+q4e+THKdaORe9YVNl5NxiPTzcg1+rSpIxg4EJK2
xafSfEiyIHosufcwSNvghQTeN+VzFR5p9Y/3GnEeicuHB1uaPZCM/XjoJBA2n/WI
MyEWHKhuOkJgY2MWabxjwxsx0+Bdzy2QvnqvVrFbTfiEedWsioLzLokRMpej7zV8
dHZXIVPPFqCiQIiVIgkJ03WbAUAzvZYAC6la/oOaWXSVMIj+eNelNJuZkVSvQ08K
FFPXMcxtKNJ9HCtKEectDw==
`protect END_PROTECTED
