`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFx9iWlYtHvK5W1DZPZWDugy6KULhFZ2mcFGkfsKPJf7xa7zple3JgdUsZQ4PhuB
mE+Dt/2G8wgdlnmUYzan41Gjx7ZnTY6bES+JrKfM6HmjmKmzYb88p6gPINwqZ8r2
M0TjHXM/J4GVB+qDx1BJmcbK5QjIUlYBahnUx3VeWyeLvSAStqj6EuDdzEcAI+sJ
PmMwW88FylZT4kxhzZlqZC2hurTW/jiH4SC0K6m37KOx6293N1M3rGvLru1J/n/7
smt0c7kLJOmJD9j9pgP+C7AE8sx0qIOu863iAqgOt5QXy4oaL3/5hKvQ8BtcDE+Z
Sn6pfF8pFngIXSYFdwzKUEsQQo+UmQ+0CXluIaMb/Y4rIl1EOA1AD3X4+UbYbnEf
QZBbEYAZrp9VQpxb/Pw+wbsX2cqhUYpKPh+5QtyQ7vbWdUZUxUZW7/bFf9WdHood
tjZkUQVEXzELC56mN4gG3UhzghVWecNt9LO2PgfH+o7ue6EpDlEBVjcgYG2yBi8G
VY8OS3wLNbfvqqNrntcrVa0uDDY1SqVJG2AKk2Oeil4XMorY3Su9czWQXpDXjOtE
Wc3LtN3xRG/KPsXNwMRcEb20sJgTjGWcPN6K1CLPlXd+fIoa2iQhDRUoumOUMyd6
rAyUnSrtAmBLIeaUW0TuZbw0EfIuBbGRIqoIpDF7K6gD7g41dKjr1YDY2TZYehdZ
pFp1x05dvb1ML1eJicC9XBbZiCvz/c+XQkcU4/5vU3gtND5q+0F4NlQZXcVt3XgE
/Sz6YE6e0Z1uJwTz2JCC+DkBzjjxacO2xaG3f+WfnB3vv5JfQDw8XJNGKkoOl45R
08vN8Cqz2W6Y2kuLqoKxzFX40LY7ra9J9b8ZI58sjfKosJFvoNf2B5PLBvvIfmqr
TiGZdA5zcK0RtJVKSyZ9TbWlYE2BaFAK++B+d7QwKgz5rrDuSwllPHF1nTF8YIb6
mhz7QdkYrJi7M+/5ss7bcost4H8FR9AlWe2SyxOsQIg4AWcQRfc8Oc83aeerDtmM
UAUczpVEzSQ/gDGnDRxq87Q5VJ6WRYCQxlGmS4404wQoF81oa39B6k0vCHvOj0Fk
ZnMCgyWmkNX01kK+ZVrwiRQtcZremSBZ9DaA8twPfQdfnnI4SyHaKOxVWuuawsCL
brFZasYqXpAYDiTbNZJdTEsQT3m9XjqMoxvnadk85/tXp0dicJMBSwUHEuvJQOAj
tXlzlK9q8KfbXNWyBeUDPKBfZQR40iEZSeKJNc2GwGBx5BoRjicqP7P81E/TGp8J
XMKU2j+iFGXi1R6A77le7LEE22VW/1Om5TIiklbXW5x8X1z5CBT9Hi29LdtqfZOx
2MQEg2uFpq5o3qfLSLDmMaZrenqfdKTWnMwwa0pjEARjKAbNlBVnDWXpWa2vGNFC
sZuKhydALiOpm41dSN8OTG5Lgbff1g+2zN70jiyVhCpacZ5NcDd00kiQXipXDEZO
dh1NhrYSTSyJ2LodJAUcf0iDiNVLO0bVQySRl68M4cjBm8gJrrEwvNh6nfkRnTnO
wBrRtNywtij0sCc3tBzkZshhdu9G7RIIH+urCGTjCyHqXIAAsIItgN9dseUgWcUz
PfMKFN6/L8+6RGbKwtnru4UjDwLnDFqEOKZ4bZg+Skm2zxPf7c4eYlkXeSindCle
jncWKYtDbiqvqVwcOEV7RuOo1rOAbk6Hzl2OFCpQbSFGvuL4WHUguyC2MKa196/D
v/L7jwlt2FKl7OGT+wBvjGVvM2Jg+64FhYGI9D+ukgRJ7vKPmfHV5OVPlQq+wzhl
UorJBi7vuJE1J+xHPS+DlIcoJln/eifZ+7rwXM00S+LSuYLbxCHQv5FDICxKAbxj
pX6pe0zcXMKwjubd7SOlh7J2HN7w5Qawe9RBBdzNtCScWFcPDvk3WIfPlnirFeOb
fHTGy0w6VjZEyoOSQQo9BASpDcXYj/8yN7cmyMY3ADBTVuxjhlg8XMl06nzujxyk
PWw7pZfSOoxf3JvyiT6tUk6Z5A6Z/Cmhy+QyHyfTm3bk+XODJCIEM1CaGKIAGCFU
d8Xz/hLKuSEHRO+xCOYSsG7cCMZ8eb9dAtQ3YhVvbUzyLD6u90Nk9JLxD3YnPE07
urfy1hVJ/qk5d6R7lNSJhRqkciPN7i/915zJt6IRMJa3WfyMRc8eiob1aq/qwUG4
qiP9XmLmA7VAs1KzHkseB7nyZD55kBMBx5kgRfA/LD8UtZRjPZVj4nfi/k3wu3lg
PanTLFgRggBrF1NX0BLGhkVKtm5urH2ZVl7W9+Pm00rOv8MCgvug/k3MQuxb7Rh3
AfxigmzyJjwMWPPxvlhfdpA7U+CxV/gMnZjxMQx5b30T0TAUNoS8jP+WNvAIw+f9
Oie9L2UrxAihHchYtQwVHbhB3K8fZmOuXhvVUZmfI7uzvc//Nlo8g8x2HL0AGpRu
4/itRj6hUVA9a7NC6ea09Tg/AatcvspX42F7d03FSCxJJdzxX3MevUlPGkas9rg1
EGdiBmj3rqERsvkL2Fv3WI/1XyhyRboPnykDlfxzZz1DB60bKC6CERKyosoWouoj
RK4qaCTeNgXskzN+/KbBxa27b1IMMeTB2ifV/y/87vxxLHaXUzqeBLe/6eBgynFS
brw+7O0huvjdGrLkTbNDEJa35qItxkanyCcKXpslRr9t/s2eYSFYyt1D41Iprry2
Giafa9VBr5uQwkWy5XcO6vvd+m5etBGSUiMM3ZxkRlCWJrE4R4Qp78X24oBgmlOm
RHwrbbo82SvW/dM7aJlpe0ITvlOksgEWg1qfEhLcaeFBs7XVAFE7TbtvdauQPHMi
oX9A3khIxNRchULpvszTzqoTs0/cZCGADwRrCbJkX70QfVMpTqIwOgjQ0DdZSc8x
F+ZIy58sYht7lHh/liQikXvpIiZgEBqlbqEOhJZjmiV3WGCLDigBYrOHhaHbPpce
MiK/RHi+Sji/Lq0+leXBjzX7L/ESQ3cN5HzczrN+az+COjiY2hKruWKWt5RrX0+6
iwknsCsX+PGKPOM/D04Sa9QzYCE992wHKrAaPdQuE1f5edU/QAgLP8GJ5pxwBmVN
qWqCfmFCLb8mSlJG0dLRr3THQDzcKfK60KQ0CbVb11hxMd35xTTazpvQGzDmSTNm
J1lWT2NUh0kd7maouby4A9ZgxiE2XWERLeQCkv7DJThkh39tEyHdsjdGHQd8UlWh
iOTcwmuAw10UcooGa3HDkCVLrejgE0XMa5EIWhYwxtD1UZ2SP03xNRtSnbZ9Ki07
K48Ncr+k/lMMTvli3WEWOX+ZTaESN9lSkrlOqYzp8CSYoeX3YybvZMjCbFif78ll
/Qr+RMwoN9vriIXMvfLS7WxgRMJU4IHtTpgtz3s5bLZUTcUx7aqUdthRZGREP00U
CX4YAJtn9/6QW9ajU7VTfM+rWwS71vxYMCYnO1NEjhOzCw35FFA5WR1VBKTlECW/
S9p4f1FwITYZDwODYB3KC7IYf72GQ86ATRwRzU/ukkxsLA3ymd9WfE06GN03gPFN
V8bhSIVbZHZd1wcJ9WGiCLWB/OBhJggEezVSvt4Jc8TQ3GizwhePm3jQB5afBlgZ
dnvn6EFYH2RiH0G9GkkzN2/Nr+IbW8alyA0Pp8LMcQYH9g8DAZoG6I8gjiuE/tVi
BiuxAJCa3zhYcMRlKmu7bHaCXRBO0MxKP4FkS47EPGsOZzUfmqZY1Pr+UqFIDW6D
5R6XyOd+JeitFE5N641slL929hNnIS5IOlUpikuUqu33JzqeFXJfz6SeLjtDboVn
u9x06vRtrQRcniVfQHkFlry5Y+Vx+Qz+B/1gzGGWkFuGnnMVBE7VGoIPnUb+oTX5
kTvVTGKma9iKE2m3OK9tm2+++p4Jrq3Ch9mUo1QzcGFw2MjUAP+RZKP9XGsRNcJa
KS3QmCDSWpLghcAFKSL66HpxnTxNj3BdmxGYXk85+QEdqy9AMb6gE6nN0Q8BvbIy
opzJkdHCsV9VFh9OzI9eOtB5OYwlhUI5iDHlkV2ppUo0xHmnjoUOG01clrC2sdUX
v4kvKtg/9+fB0UT/SewlnqOojFESOp2meSk0inEFxw2Z3+cyJNnn/g4fjRn3tjSw
030ESNbjlr3bWgP5/K7OGbFXIvAhKHQxvjpVknSy2ucTOlacEE5otSrPIpO0+knP
Yeldo3jfAxJKj0MvaFTI+FsHnxasuRvtnabq1YibKEmrNJQqPVdZk9GjycDBNML+
rTazj3InlgGaY56H7BsZmze1jJvULajRmj32e6jeQWyymzByoKdNgzFmfhzBFsD1
WWpOt/qZ1M/+52XLGCeqoR3CyBd99/+zAsWiQG0RbggtHvg7fHSyN8XDtt6MAFj1
zsmT0TR5oDxEQ3OGOgp7BV+o21bi6msAfbTyxhx7QbuGoS2B3TFqESZ6ggsgyAcL
/5+hCc5ey5dqSrRZ1+JTvXQSyefHIjZ1vGALHxKypcqzUN+g/QW3b5hPigCwwf6H
qLB+f9NyvVE91hFyqDUJUSUp6QpfY6as5ALE2wb/ZlaXk4XpPvlevcqLMqw//q9F
5ShXVZLQcnL0dpi5LhBH2T84ojoaIgvHMaaUe7RBfIwh0GNTWBInieLRODDlJrPN
hqWM9Yd7deP6BfIo6vGl4QyQEKfj9VD2PiQCB3Ag+McBJ0819OWnFrNmfWUOmRqT
S/BZ11EnKahWqVz2+2NJiL+WZ5MuFX5HDEGTBI0vxKGUnSC03rC+YvB51EKmX716
4l5qeh+SGPr7BGoBm3l+Dj4OOyD63N8TSapAkvZx9w1opKBc2WXicpbReZqm+IXQ
SHNZ0wefQS437cmt0/PAK7xEzIpL5Jd28dI+zt9RJAzdQAjRyeUjrbAPTS9ZWTij
m4Ml5Z9pARjWrAEGY5JBtWJzvMJ5R44mZO8+VWf6Wc0lafeHRfofbwOpwswdurz6
goHoORWgZ9p13j00YUvlPrpvOXcYuNvWe11rs7eRKDX+L4XDppoRi6+AaP9nstpB
YOH6o81zt9Qb/nOeO8cXKHUpAI3Ya3i19IFwm6aEfJ4KAwRwms4VdEP64cMGxX5g
XjAWycpRNY6RZ/U9gLLCwjIHAUINl48cJkPBk2O3G/rbJCpmz+9US4dA6pJ/4SSQ
48QyxJd4Q8Gh1bdQbzjGCOY+3ylGO1JGwUzW3Z9rKiX7qbwUrjLOZQzlbkd8kceR
E/XNbysVsNIu54aYa4BX6TRn1YnsRvH70rgv2zUcH02dCtGiKHTnjHm2S5qrz47C
Kqf07rkJSN40sd7NTAeGSVq1BufVwfK3PSiLvvdUpBVDjy5sq17vejoV+IJjRJzX
gMbE2jVM6ppZVOSsrncmY4Odqv6c7NMiN0crIcJKKWS5Nc1CyeoH1SmpwAAtbF2m
sIpvI9iTwBUPRB6CQWv7XVN+LfG/9vmmL0wCYmmafk8JyHIDlbtZOI8iGLxtLCKA
yv1JxDGqtcme8XUhBgz49ENZSGiAODVdhRduGk+LArouXjjppOsLKVKEEJtjzN7q
A4pA52w/vBI6L8lBfEgk+0W3+lcOuf86yPvcusPOxAb+Xod8Beern+e2BuFCVjgl
vxagR1em1w0Y9L/Up1QAJu7SxQ4u52zDxzFWjBHUpYHVJhpinA4g/jlAPd0T+quK
uVuhCkpDRQgU1vITGUmBRM370E7Y/8E8K1enIwsvnVSf68udpoid/O+bVNtpRuKg
4nUy8JxxX1H8k4aA5LvxfSinPCE2D7FopbV2mOHpXoS9RXC/F3CnA5NECcnvw85p
AuLj3MvCYF4kMK8Whdn1cBoE10WKihGxJoyy5emJiu/pqHRrudQYEafjJI9HONeO
V+oPrg6ZfbVlayzNyPViPv8Zb3i6PDGbM0cC4/sC5AjbBhHXO9VSe+2KFvNmYPxR
6gwe3WHLEZSdF0hNzQEzz5YIKikxzV+3KdiXFrOibFR1z+izfaS7lCejWCK8tQnf
SCuUfJ0XW44BaEgr+LLEvN3WA9Ci/J3c9TKrBnm0tLW/o1saskmwRG6hRrGk/AlB
aghqZvzYrFkUCY+L0c5bFqQh4indWP8Jcoqgaf6pgom7TeqcA13iN11bh/5Y4mSn
fqxj52QE0iIQA2dqLUa1DZcUgIsXSiKOKmD76uWddLnZRL5ZV5JpBkrVGgMD5Xs4
ZyZP+S4Q8olqd9YklaH1VNIyJNyAhVlG5xmwjFQq+h+vlnlfJrCa2Nuorgom41It
jb4klJL2bb5sV79ReLasZE7h4f2E5+wjyyygnDGAzyxu8nYcLhBgavCDyzDth/eG
dzZYRdyKJoZVGaCwdJbFcY3oR7vFA53nvl4a2LMKitU38Tis3B1IHW29QAF8bxUl
0ksgnvwo4v6+cDzF/gXJJFDA5ktniI1KD3k/mxhGDqs6sK0PTrCClIIgcfZF7ANY
6B2PHgJLgLZOjD+7LE22H2u5OgkJifEfIshKU23OGyGZ9W5w3kuCMD4YRAmU7pyZ
Dhko8OaZkZTAMlztDIb/20jziw0nZECw4QOkF0HOfG2NmbUpL12xnQNk22MWtWRY
1lojI/hezT3qIKZO6GjQgejjrmhpu9gDCXdl2ZpYAMwg2V01JtWOoRHj/2NDOArp
9bjLfBUByGurAXCOnPWez3j/EjsFq5NeYz715WZv1NmiMVviHDnNM6NnP5i4g4LZ
MfQkLU4G6GG4ltIEVOjo7O/AhqkLUdMa3JaI04nTr4LRRlpoOiPG75/Yf0w1JFKi
Nn3GyReANc2gLbUYyFp1QiKeM90SMNuPbW9lB8HLcqgVoPc6DSGrP8OJSKnBGsvL
aOuS6aM3wmCHD7yjlZUkyP+/X560YkggWrHWeXJ2UdF08mh1pEFxI49aCRZWCh9w
GMv1ugfaNnYsQBN4HUsEyhxSsmKwm8C+7eEvHbLy6uxvyo1nZrHo/3S4384s6cst
PSjnqW9NugWPsoyKCrf5FL0ymCTI4yUeiQsBWILeCMAY7YAUFn7nsEZJx7OMaWca
rXGA/nw+rX4JXKPtdVkBQ1NZfnqbu8KcyJ/QOTpyZ1nlbQ6TmmySgv48lO77+vTz
iCNCAxlL5i/D1084SOGubmolHXqrLpuf2OlEGT0xvHawch5iSzekszlLIg2M4tlk
hma9QOWEamgEjzm9XBmSQiGHlM0lmVpnlaRSeSpX3Rst8w3kQLoRCfViaBj8RQoe
8unDiJ4ZbqQDHOVxjbfNMmYNAIHtpelXjC+rvvxttlNzsLO/5cU66IUzmA1ObDMx
DDHRM2IFbWAUZFtbbspvgxTAgEsWepLCDhttjt8RsLXkxszF92GARkZyDoRb2WQR
cHLYGbN/t82su4/qXco9JfjbaSSr4gmuS6mrQojE41I1Yk9Eh7FD9dgtP6x7SWSn
iaBH5z+BODOj2jzj3ktTDH8LQhLDg8lLLnjfZgx++6ri3FhZlfEaJ/FHqhUNCPVW
9H0nfMSewDZKQQ7mHBWUbyfyqnfBMGsyo8d1x3p2UrXz/9ZuYmaaR/lBsk+I0Ugr
RL3ItKrysSQi2MZQSdavGJgEbepZ5Z3SP2Xm2k1qJ4s8uPbZzSVzxcEQHAr4HVhK
0Ispoj0T998hHEh+vOMz0oHNa1OFyiQvs1gavFbix0G2vUfGfCqiB6Z/NRFcYUpR
PZxGAg0epvTQcmljITo4sz372nWj08IHU/7deuRhv8z1iIvo82QJLfflNxcih39n
MRb3YWkWJ307cpDTet+tFa0Wtf6wGPuSObvtUEkxYrzUZhRxJNFc6aPVzLfJRBi/
20a+FIsn4HYGj2P4XSgR+0UCjxSPZsMA8/O2H/EgvPdENV5jzdeUXPpMGOAYhZVU
/xSCoORy9MrmXtAPDWu5fjFJj/1rzZgOsjeg/SJT4NkjGgy2vmjvmzK/NgmiwIQn
C7A+dl/f6KWd/Jy1QR+nAfdtT9T+9bDPgeJm+WQoZxk/CBWDBv967zav+H+eMJJ9
NYRn614dvg60PIA/JkLeeayeMcQHlOklEN5VVuZvwermd+FJsEmUeymx1mnmx7cB
+gKid/OPwhGsk9EDrXEWAoJoLwEzB6d0ZGq5QamKTk5SMkHnvHrkvsiv84WKFCvS
bwxG2t+VcG1hSRLZE0g1F/3iifecv9uiX7MvRnYEAwSKxfA0ycrx3yVt6+R6GQWM
/1HLKNnFgMZF23vAXVIxIXp+pBmFw67jVD9I3tHIByKxr5DkMJFYTN9lDiypUO0w
7B69hsAjs67MJc6FH3X1Swmo034fwJFRzQS7LK8PcVx6i3ZI8G74+E/Xr37id+0K
p43tD5/ycNdFVrIE34DPk99kGS8xO12Pq/aAbgf5KSVwRLq9J1edVTk9pM14JPna
jjnoXSlsoDmWtDihjnbsO2131sRdx/0qtRnDgs1Z0jfBrWgPTctvVtlspLAt8y72
ORzapE8jmmsw4rRyzjQn24OOZqJTUK/o8A1oSsXJ8ABYt5WA5spvotCvDrxq9VYy
pRWGycFHXk1OFo5IICHWIwFMGGzbtIpv2wu8p2JshK0SN2wz546qCnhDINqDGFCJ
987btaSfSKsSGXsqTkPAxnxIBEwP6vklnUjt2hSGP80XoemlyHPCTseHuaQCW6uR
g4nIL5fBLbs1zMcMtiR0MhSRGp+JVgo8jYBkxu3OdH8iMHxTEAoGnRO9vEISHUm1
3OQGmeChIuYR7408uhdmeXrOAlVqDzzYUqGhC0YgNrthy6auPg9gjs0WNzWJau5A
S2NGkdCaSwuAwsKPxJWAa39SKyXBrRmUa6JuH19kRTj6+NkZDe7UDTfr65pbmC5Z
bp0yBYLJVjCqLJZmz15awWrPgJZFb7b3Gw7LTwqv9/rAL6jLPBcptwFS8Dc37UZT
eqMBRp2olspfh7MTwy4e4EO1choEyjg6CR92ElOCiDyml7jQcdusT5GPp0XRnhML
pGstReuqQHQT1hcTWWAaEFYNttG8bBySJ44TOvhFxmzQrD46Bqw2WRwIeEWXaN4m
Cu6Qow8F6B8j0tovwrVS8luBfRb8YQkcC6zFnV3P9eaff1/qk6wwCqwbqmLrWj96
H4ymTT6uK7QUtFZSSNJi7xlNVqW32vfdLMp2TvsNBH6THJKIIqePLdwfctDEx5PR
83DKq5BKcIsIh5iTwldxHS6XDK7oh2eMiPV5VAet8+K4IL2PBYiXzImF+TmXQpUa
AVZF0U33X2dpZ0gqnMKBWNg3n1cAq3SGu7SfPhJZ2xpdSaR40bVTqmYBY/AnhNX0
ovKbGYKU/x6j2z3qBinUhdkZJsuU+QWf9P1p0my9/rSbeuwa04dhPqNGeoAfao4K
sQQwKd7P+L3rru1dNVqBK8vj5fIvR+/X62hcUMNv1JdL3GLEF2139R0N2ZDmurB+
KRNrrq3FBnC34cdKGExeHBw6fOwyXsRaJY+vFCw62PxUl/gFCuhgGN8nAVZdYkpH
zcAQMDd1NkwvsIuUJVFqxOf3hyPNys2bobpOE9JCrXef8O0tIqjDvIPOWVQo8zgP
ISyxrn69qSMTqeFib9atgWVy2TVX67e2ktAzUd2DKweEAYOeS4YnFOxEW1pxUWsA
JuCR9XMCHB0wY22cDR5/cVuOynIWp/QgvzMw9pNwwzlf6fTIQMHP8kqJOaSV+z7X
gkmuG4y+pdkmMDQRjJ6nEbQ/rPri0eNZ8k4+2GviaVCX6To94Pv2jt3zno8YGW7e
qNr9EufVGZt04CcJ5pFEgCtCaqak9yicDMrTom4z6Ze4h/Qxq5WWaVdvdCoVXsqk
xrkEZMNKJFZZ4AglYxt9Ep2QNR+rueBzjZRGz/rPQTk4KOKmOiSKMH6YXD37jkTV
jEoC4asgmRETt89XUETP+FSB8T8YOOd5qFfhoQOwAhPgnyowybrsQ7/mFMQG6KWu
d4MknwG2Nl5WYU6RUCClrcME54y03rVUu2tpPT3u5wqS68rQMmGkEaS8gv+E1dln
uS2e2z0rXQmdnfmYEPAWByZWnXxX080ALSBZkOGMf6bXysN4PvJSCATqSVJClnyk
cjHDlvjqaZk5GjGdKngonpV0eAPE5iQn+Sqt6iY9IwoAqeuF/wIy0kgs6PARpdyz
BKUyRArJ0cgoyfA4an9wD7L8esu7xBNexnPTWaxF9ssUTCczXT8BhpE6XaPgLBCf
1pmrQlb8y5KWfn37jAH6IOnFw7+VBoCTY/6ncjQARYHtzlUXol0VKwUi+07Amyic
aQfA/qDsD7PyIDk/MhN6syktfDjAxlxfQfjhLpYen/BbQX2j1rPUcSI5p3A6ukOi
VgPvbRzmntaSO0dumm0pe1anEhz+uhWJWcYjNmC+5UqEASXCbHA01XyokMQ7PlOS
tcrVfnaJnT76HzDJ2FUc39X5yphb7PKfRgaZ5CdkH3M+tVVVqei2RRE60mXX2xC1
k7QVHJ74EPNqCoxqUqjVF9YnAVT4S0XXfButraJPYGvQX/tDV/2NfuPPIhLfDQX1
khr2oN+aUPukO9OaYKUs4kCD3UyfQhQz4zX6VsR8pX4l+le2jQdGHTHP1wexpyGt
WIeZD68Qdux5defT/AJKLR/L+MAgoGfjCGPhtnS/MC9Y8aAgkVVYG4I4sLbIcrM4
xDaNuuyfeQRSh5/ChjhucDfSfrzHxXn4oeLNrS6GiY4BVtXQZ4C3hBvUMW46jIQ/
qxU8upm5HFwdhxaSteJa5qbJu3RY/Vo0+b/7Bm63bId/s5OIuI3Oc8MwNq9w0Oxv
L3WfoS4DUlaTXDz+ATyHkNzqlz8nQesbmNR4ARPxfQDCdMvtSWnBJNjIASyL78PI
whfmBnvjs3/ecJE6hIZpXAKsdau4uhrM2ePtEXwbRQO2JdPQvumbgqbqabuKV9Eg
I3EZh9gbi5ojmPrNji1SdNT7yrcqQBYNTTRvAn0ZMfI+8JEiNjMGDNAU3s1feEph
+JvnZoxBAL2gluluExNQ/PynqQQroe0/fZjGs7yQPtw7w+2SxChPU46cKsbuUh3h
93mOz2wrciNI0MFEuDCmXZCF5/X7FYKcKf1Wj1VCLmovIsUfhacLIE/VgruFBlK8
st/94Y5P71LmsHFrSKu9a76DyuslVVw+56uXPLU//MqcYCW/5MsujwOb1QlgAaUc
fmHKKqQsTT8ogl8x1RG9899i5I1z+GDZ9cXg7RAZ6fnXk1wpcA02AYW5q3g7ufVL
IoyLeWbjivmpc1gaS6Q9vt2nl1/xHPvEnk0NvxLSAxlNopq2vSZ3VHF8PsyGWoXC
w5s0pkK8f8R3ey4Eznvz2cQVum8w2vB367R+Xsg82zQnB8CK5eOjTXbc5LmTnMYg
3c1+SUXXRApmiMHyrcxE84872AE1deWPboHqCIh3APHpJsSUIHEUR5+xYzLvON9r
8hU+ZEyrfTPgsRZt4qOM7RSEAJ3+VXVn4NXTcrPIm9sOH7P3ATfG/WlVb46d42CW
aVWDePB9pkWeeYSZbK9YF52u1uqaVBhhsvL0IQ34QUpdCQ5pu75Q4rxsMLLPpprp
8Ws3c+HAEKRGHyrdcXa7Qi27ouEk4M++bduPIrQzPaWJM1NU7jncvnH6MtkJ70RM
OcW1pH0Os7vb8lahJ7HwvLP3SZyWK5zpT/Lc3QlK2uY/UT0LXEsDvVeNoSX+15dA
NN92oj4zhPN/qrjdJmMs0s3OzJ/FJY6LlLLnSkiES0brngl0MSLAdXr58MwXto2h
rkLiLHisq5oEuo7aWpmLw2TDZi0WLUb2GzViXiRhdsz2XFY5NDY6u7V7stsb+9md
ClnpuXQGUVV5CrYqpRoF/vDLq+vH51NsDdnHzwBn8KsM4BqPupzNopefocjc+BYz
fUba6KjL/bQ9lM+amHkqodtONjrl0ZJhCDJ2nIgKLEcrufDJFLcBK16IybYFRCXb
YhFmCHTm38NNDfICwO/Ed1l701uhG+cX1sOVMK0lWHdR65wWk8mqi2Q9EplYYBxW
8Dyq+mDij0VgguqKEgwUHskWKm43xSarCKfurcX/Yoh+9Xo9KZUEXrVy9JhU3OIn
tdh8SiirtgCNarCikjnvs9/NMgv5VA+jQswzcleVpvUQpzh/AgxAYbtBtp5XtrCo
4HidqS5nuwA8De7gq3aZjlUsfQ+gJrAsjuflBNJdCaTE2vHUOphOu5cGweSuUG4f
9SiBnpb3V1NJfbhneWC6LaAgStZyl8dtljgrwTRgKI+uLL3PqN+zUoVhcUIn+u3A
mTSXTr45lARzojBHxQzoZJwfuZTnxhNjUQfdDOND/b6Af2zhEpBPFup9KAZJWI6g
QJoGOKWuGLliUjbd9SJrUmBvPcfPHFNIAgTC8kcMJg+E502d9CjxipAVX0hfuvUm
vFcS3yx0KKjM0fue/Ydi9TVIc9J+ryPWysTVmdvLs6b3MR4cQW02JlOZ3C1V4DEm
5MEAH6OzdkjvnP8UGSH2TaUa+3wKVwJhbEN6liOdEeitcFig+6waZ9vZqmtXEp6v
i2K8XFb504xNLdUm/rHJdl9IbE1WVK9KK+ldOqII2Zwe6EqqyVheSupAdoAWa9OF
Z3jdJHA5JHZ7YiTKt2uXCrIXRHCCaz3D1gxn/5/9b3tAKwv/gSggevqZr/IA5WRP
GEGGMtRNBtAJWiFgXJRIb9jgx1c/qo9Hius7wuPhPBWkiuOgK+q/gHjDHZmRY7gQ
v7lrIsITOGoTnqWYd4umCVyFKGepMHoslLjPWgW+dig=
`protect END_PROTECTED
