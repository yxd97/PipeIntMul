`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nVYtV6sdjB09Qbdex4fcbYGVe+KhBjXDF9sBnWEHo65+jw0DH7dx7WwJui/9zzFp
sF5PB85qVxcWrS0yG8rcptweApXTdewGsED64HcqKA9l5sA26IkMPuHCGgfhO5/p
X5hKFwCacagR3sSM0fqtZg31M0j8whrdV7GqmLf9CieFIT1hq8l5gXE2iMw+2G9c
itHaVJVxEhc678IK6xdmdaEy1z7kWz83AN0P9xDE58bbedZ2I0Rfk5CbbWNPgn9D
s8AvnWe60FdK2d230sEAXc1awpRuR4ryJXx5NHw59wdX4CKzafPA2j0VMzKsuSAB
gp400+nVc6xixmkioBnE8sYSZRFi+lIV/AgFYAAQYUYhUiad8GT9dO9zIPRYshVu
CVN1rjjzu0wmh+9T1CfXDSk8tzkflejg/XUdgRqrRfeYeR4o1fRAYWjYl4U3+Nnk
`protect END_PROTECTED
