`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1yX9MRyS2AHyc9J4CBjM0aQx+I0PQsJi+XfT7pHG+fm+lcqiuuXErCKia4vT8PH9
MisygGWSQvC/TbGdCmSKBjn2zywMpyRK6lcnA6sYxH849c32Ko05lzUNzvC5U6mB
J2x8pYl/oabDA+3JCUlJuBemax4JUrk5HLmhY55rlc+rBnrSHNWKkMYcB6xNcWm9
bcJSnYU66Glzv0zkPthof8BYun3zHIXmzony7qdy4ZvklDzDUkO+QfDVLJI01WVR
K7cOozyLAF8a++fuipR4JbBLvRbHL7ELH/0ImU7BLhXBxlt5/M1BC9tA1ZPfjH0m
5n9gIz9G5/h9NThugnL2HnDb7gd+ggSkoi9twUd34DVeLUTK01+OR5YmlqDEMmys
PaWSc2xK/DJRSgQx8Kemje0CGu6opz4b0xeJbR1nxId6YRDEB6uxJehUE49COBzm
On/E9nWRSCFOrpDaU845oMVFWh4lVldnU+Dsp5PNfh6cBeZhMlWNjdffUg6Nv9n2
zd+cvmf1orCm2/7gs6KaiS2KEZbRe/5OCH2uRFTmPT9lLgfHuXOyAJbaTQZXDlL6
4EiE6zB6dZcrfPRgeLsXpWFXitBOEuL8Wqxb6/Y3ucdiZX5UoEDc72HBHxC6ENZy
vkrp8r/oK39ZC4YRUVc9DJxS/CNQrXl9sdpvnHvCqNcFhMFSJwJ3rQT/LxByYPE9
Jpzz1ptwdTIvt9KUYY+a9RxZ+RNVKdv3B7bdO5pbySzcY3Sx4cspIY6rrMSN6d4r
pISPWJrrUAZGNOS2K/q2fmFchX2hTisn71G0r8nzgzysmrw0qVeqnwbAxX7X4IlN
UB5VsmN0yGvG88i5vUZuu5rlYPj3pMEhqci/tUQjHr3fwu5ALkWmNsese9km3PVl
lJBnzyoY6X03hUcLRHHVC0U4zB3e350lEtYYeVQQPJyi41Na33W5Ba+GPqu9zXgr
DY8hGIH7ASKIZP5S8lATjCgGYAPBNc2og7ScmkHy6+qrZcxbjWIE8DTqhClbDE0+
rMKCyd0PrEnd9u+yRLO5jeV21cHZMLuGneqVt65I/z+Lrpx2LmLazDCOeem3WOUX
bA+jTwkOpQRTD144iTCZCQf+bdU0Q0TLJqVbj/rBY4gxWBut+PKVlZ0vlNBMICPq
kPhxqenlv+pwPj8OvDZj/jypTcW6FSwQdVk7ZjMPIOUfCPpBSiRzpesFNOa34UgZ
bhOd+FlPC5ef9VrqeXL00PWcNsXJdMKC2l5VJsupMaua9A7weLeTcjdHPrDl9oDw
NY4m2vXwgf6LuGS/oAhCWWvRrNVWALP+JZ7E/FLJHn7M3QZgaQqesit+eaEqEHU0
n06NcQ75DFqH1+SymN9MacEn4GXaMd/OmdlfFNvv5blka7sZn9kk2VPpbG+4IqWq
gEKIBCENzIRUFKaPeL0AbHIMtBwcK2wABwSOZHwEHQvTPlk0TOP7SAvwPtq7Lqbn
rnyuDFlKiwAk1KlfMsg7KATt7R1dRwJ0WDYlrXXZ6yd7rqtk7l6PS1yF+It32cop
CjxXs+DXz5p/OIH8k3tCSEBb8C/DTqSD5226FUvqaPiRTexlDtGb3SmkQMUvO7NU
hkgqbKeOA+nPhVfcY0q4/GlCa5dSAThxgfA7PuyZkY3/TPSzx8LQBTdHujJkOKgi
hDBHIfDdtUUfErJO+FpuElcXvoyBv5N6gcC7ZS1HvVsLmyJYaoxHrqIsElapNvIw
0dNvXwqo90psadhjV11IPIp3mgFC3WmbYPF85iGDqqLzDvHiL3ZOz4t8CnikodVv
Zc2hh5kAKhQvQf6ktRCPhNXoZ0chncr7fgfUIo6EkZTPhXV5he1HTMnvKSDgzNSE
Dw2v/oLBwiWDJb3HAG7CfGLQn62xJYRCJR11flTlsqEUsvBXcIMhXzLWMUiN68Lt
/l3zRoxyhJiLjoYRA6JW2GEvlYy9wbb/0tcxCpD18VtfebvtfoN8LS4XPCCOGKKU
i1UFI+dX/05A7/T7OB0rK3MphbWxcqJmpX7znmvTpy6VOwYpR+tt5nrn0vP+Wlbn
XELb87lgkdwfA7JuMo/K5tx9EMuk1UKVuEyUytmPqN3PiCmIzST6nxLN8TyOKHxO
`protect END_PROTECTED
