`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
147TorgRBA17bYQcoVou+JYYO2BclOA4EXAc83HEVWB1coJxVBm70R7lOoKin/8F
k7hm4g16OMgm3kGWnc4HHs87iG1yBgpbte2lkwJOz2zSnmv/xxwLaDYyv+qG421d
pGEgJMV/vfL5tKayLfuTUjLqfFA2mTvrfvxsejNoKGI2ndyvTTeMpSiwxmVgt5dX
NquBiVso3WSXPJq1MwWkiszR2P2QcXUNnqHI3yZCVzm8EcXljV7rCSbvdpGKcWpk
Dlmd4m/atEGrlIzfy3JNXro8C7FsymJ4mJ5ZevTauC529OExtfdSuMeAoTTaFGj7
r4FBx7QVFiF1FxNRaiT3driwU8OLGmEVlnMyaQc4/qTCugVQrZm0SLjacO/X+5iY
E5t8eLnASeShioCg3H2UdQh2wXujW6IFbx6vi7SjRxzADiQXnKBPwgAYAZ9/xIH2
3bJ+o37dbD1wwSQfX8W8je4IUcRlLVQdCRJkmHWOTwoTQPvZ9UcOR+qUD4R4GH9I
gc2sTvMBO2zX1p7sCrOm8wjXrmjjMmLvDB8PaAMLzgte7d5xNV5fSOHzFQLA9ooF
SsKx7dPXW3bCq+JpNeeoCA==
`protect END_PROTECTED
