`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eF3gbkxWyU/IqnF9EZGthgokfx9h6LT1N9u9CsUsFq8o7JmllzC+TUDArbArZvtI
/2EXs0pHIVZFoeW2GwbL3McaXab/sveuWMVf60fdqy9sWZidQKT7EH9hKdxuSWWy
EaV0taIRZ8Eu0Jk4dIfZinXb4HvCuHs48r8YJMhgFb6VNijHtQE7f7FWxL3nH0bc
Bo9ewRV3rcR1YTRlwo+i1rMKxcWS10MfsNAyuq5Ahr+e3sPbGVQ89XpoHNj/wDI6
HAfQC9LsJhesLkrbl2LPI/RPe6x4gQsrzUwXfGkBE4wZssdsVKuFifOJ834orID/
MD6C5Oxd8MOsbTcdAg2zt/iGtlEcXO/j7ifzP8RQmvx/NeV+jKdOBTSBfw59n2L5
1cKUWfAavn/bIeu/3Bbfa9RNJUMuoEJgHFUxqleKHvr2kmvu2879RkzbUZHoCjxr
LhrrnrfikViC1/HDiZhVKltpNaAnX+9RkuJFSCYBEi3JkenDnxvYQ6pKsRDpsOmS
yufqINx8GIhtgobuCuJJmvIWuZPgbXnB11WnT9Q6MUeKNFS73WckG32ZdmeiXXZh
OzXzq0AL1K8LOeAzrBzFFkdkiG0AdaKxZJ/KY6AmBfNNy+ALjWfbRteYeqaD5ZHt
`protect END_PROTECTED
