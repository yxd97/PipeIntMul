`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
66k8cxnMj9ohqVXURR95cI4Xcr7bO55wxgbBZyJbdJKGB/3pj1XcEKQLXkXbcZY9
iYuR3R1fbyzgAQVvGw02X0K4cu+NYU02l+kQtIavdwY9HqbDmdJXYjg06pxNRXrz
kr93Tu10D4ybytYjwyLXg8wfPonljut4G0OrWSxwudozp2OwBmK5PvSd04lF3yXn
v911sMNpTRE6kVJ+SW578SSlNGJeTFEv29sXrFRrXPB8OsrZvvx0E2wp3uFF+2nB
OG/wX+sn6kQYytZguLaCWw==
`protect END_PROTECTED
