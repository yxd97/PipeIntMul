`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/rEynbnJo/pyfMnIimaWP1ER7GOHBZvXrPycdMRUCbBGexAe+WndFy6jXaeF2UA
xqqa12oUKQhIrkqiYQbbevOMJNJ4ozazohURvfrZJGbO3i2PaLvPZ4PIE2MzoRIo
eJsn7rkOhGzzHhCBWnmDmtUEDBHRLOIJDFrvfB4Z927n3HuDMbTyyT5k0mReeqXP
aCXQyruraZFARcFgF5US0/SUHau5lkCQuJHqCDR6cE17gIBLOwkXojKSGFsfoyrX
SDGuw5RWscc8X4UbtSwMCUXrAyeoL2YunYtA/PPxH/EdJofKOIK71L0n5TKCOSXH
NQeOS4n8NDRV0lrLs/TnWPIAyu/o5t6QFFOyENt1Gzbbo3hs5ZyYNq8VX5R69tpl
qk51mR7YjyczOMJ4OfmAMGZYNLLs0etGoZSZIv1dpQC0/64KKVw0YCsc009ppcLp
`protect END_PROTECTED
