`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/keJsMzNrTn/nDo8BPqGDzA5/38x88MUVZCQSH9RG/dmDHLnVfU7aCrUZ235wucH
QD/JMpwjQ0SRd9U5yZry0CUncLBHMtSnK4aIRm0ANv2avgVR6JaZNRYREC38BjPG
JwpyYdL1ysu8cU/ZwdT8dVFNQ0XjOVSrP7PEX3c7PZNFvwph8CeTxQkk3AhV2hUu
TG9Ju9z1yvVqVNeFbKUJuoaUwTjUTqyOZtWuU/+AT0aPVJieXfKUz0UsECz63s4h
AmDMngl7ry4syfq9x/8ZJ4eDRJTWr8LPdDZrvAhWl6uZttfMjUWHF1bXhggRfLYx
CWUsTiH29z58UEdcsoRkPIUNuzXQr2qACWZEFtvlQA2S0MWF7xAGJ1W4AaRy7+qQ
EbNd87r7m03Huzlf8Z//WMuiSOKJXIun600y1pSsoR6mmDrZgPDqSb/JxDYsNtpj
`protect END_PROTECTED
