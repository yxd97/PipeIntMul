`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nzv2S69babZUwB1LiVdD99AjYafUE/jh2RFlMkymRHdfUuwUcWbrak47wICZqNcM
oYn42DLxnfjsV0CpsqtfoTCCOXgWqWPBpwzz3ODiTMGsM9j8pq3sgoXJgLKGrUPW
ODP8kMI3N8Ti3OrcFmQl+G5R/pQk9NguBcj1pzD05iGPz4SaG7DxRIhyKcQhpRDn
Yx9XbTN+FmbKakDJbXk4awZuyMVxZtJSoMBKwP1vrK0yylsT4fBPE9ar6IZAVHC0
XILuxTm9YRtWk3Jm+l2xehxRysoGJWVr0cYBEqdBjOaRw9Y4FQDVQpVSpA0sexK4
PUVsROLUXcucKinNFfNlvEt/mr9AjmmQNA/5IW5+i6b2lLGBkArtpPF+Yyeu0qba
LUEBiFGtn4YGdBjlq053+A==
`protect END_PROTECTED
