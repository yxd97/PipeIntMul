`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zMhMwy4+rnM4O549QBpQ9N6tvCHYjpIf/yDtfDHYrXaTSQQ7jAkn54vKX3tFP9bu
ByzRShiJea3+Xg+8GRbEqalPq4pADGc/YG0ZwwS/pXTFJeQtXYAqShYkItW7/939
nvAwmTy97HebgBFBzYahWHxfFeQFRtaGxwxZku7M3m4Yzn/1ozJxWejk2Ru56YFN
4YEe/7/ToGJpIBAwwwY0m5jFaeOcpFLcSugAUpyZd/0ZLTMRv13lvtFBKeSY9hRH
Xk3QDiKuzmk3POqypkP6uSHGs52O0wLMBs8nLwqItQRPUWsqYSl9dv1rDpRwJ4tN
aN8XZGyvv0a5AwEDfah6hSMbjcgqUA9wGQ4zOjYhLIw7FNpToacFz4ljqhoi7VK8
myiUrIt/PuIfs/RxkSg6bMfANZaLRB5FiaRVcrZGgEaGbc0ucLG3kLPmQwgFMIHm
NH1+xAEmvkNzGH9LE3dMRMoPt7mDV048tswm1tGknZbP6Gjya8rGZ/U/P56aZjjB
AO1C3FTv73lCLii2mWDJumxW0W/hjTPlLfMf3pt/nP96AjW03bmiwHLngNeTW1o5
t3CDOoW4m1RLLf6aS48rn3Ktb/saGeY+zwL2ueGfBA2WI3c69Dd35WU3LTIkSGzU
4Wdg0pvgtN34nlCRD+IdgmVPQUiqn6w05CD8vJItwSpeIlOGaga9SQ6k4bU3UhU1
cDw+qq7ZRCM84RDppoYXE2uQPiccSgbB4gOD/6v7D595IpAMRESC3E6gaUNuXdH0
93snwjHywWHfJHZ/NecrcLoy/ft++vQiiScqfTFl7u0JY/jzMWBOiHJXOc3Ehj8o
tfQFs2dQapZvBmlZaPKJqU/2NPWzWlYitiBMMUufeuRKWdGQx7yKh8AaIdAd7B+P
vPf2QpWRORHaQ955jxQD2mQhtcSH7LG3HkQWf0GuZWPADxk4W0NkE5xLMPRyXhyG
kdfJ5H1915CbdJNr1RyPcMPWkqlOfEPnDzLgi32GiKvJqYW6m6b4h6ZIbW3VD9nw
3sJoVijYsyID2q//bND1k8fqjn1dPeFpss5i6b9/qJ6YsVwgjfuMG3JjdLRdEkKe
bEqyQfyCwnIrPrcTSuQ6qXKwZd4I6OvbiTIn6GtkoYVc9J1+v2UIZLym6wC2hWA5
cFgaO6hIusxg3XE6k7mYKpLYl1rC/kB610jtuYoZ1LvT9NJKbCUaG7TWSTZ8d7ID
3IBBZORky7GthM9bgLvG1gdLYWgqzQr9XDF8L9lh84Gv2c+ZlePabzVZaM5k5JIx
TalNgI9N/X9qG1m4GiN3JNYx3hm4dvXZavtLJGO6MloQQo0/y4kwuG2Oi8lUwJLe
7HFKe7oRZqtAC5LoXNvWye/bebrHej/XoARL/7VoMVSyelNqv/Mt73aO95ZBYGsc
mywic2/uzo6ZlzaA8lGNAluEbXmRwhKYlMODek6oKMNhqrJtbNCMZzPlH5/T29PI
uGiAFLJbEcFVGb8HdNEaB+VHinE9nnzY59umpusg0W23NS647gsckVqG7YQNwiKV
1ohD+Dvd/RHcUQFutRqXdthL7xTRCIXPFcFFEXezWRb7j2nO9mgMxsQa9cBOh/Bw
31fNbQHuRDaj+UGMMexH/Lx61RrC+6TLU19Y2pUH6QKUhIaR8uc70nOhAUkT/PXZ
9cwceeUOKrCS0sV1d1vDHQ4N15V2h+9dCYBd6Nvd4o+WfFj8VF0XHCo6LrSDI7as
hfdMaOyRiUeS2ir1iTPuHO3Y7BSsaKBmehqHkZw5LT2u7fbd8MWrALUiGdsQoCF9
B0ltVoLX1HqttpnqYqN7NJkNG6OTFIsinCgLm99lU2rm8BYKJ4ZfT0QoGMqVjywp
0vAi8vszQYBU3bOq0X/CbMQGXuY52x8v+BWXLGwVR1OkKhM5lsV0hj8O+COOmYtM
YiiQxDOsm5wtwPnHyUdZnA6XBvE4OzaD/pOOAPDZVgAICk8K5UrEy4sr+znlKp41
+8Vy3wZIm5coiMm5i9MTM+qxPA6IRRIv7kyMSAMOb1VZR03PjGfUZy/2dWpVcyhy
xEuYWGGyoK6RkEdXw+zdh3zHMrVl16Kg6J4jcx3irLjb4Z4ExDIfKgWBAJSktGlh
5ILkk65nVLgoPzxk2kS33ksJXp/cFQkg2z+28dnd4fhqqszvioxi1lcybsxCzYS9
YffQI/081Z75AZtl2hG2YhU7hDksGD2ZMVUncR1+7rVvK/+wgFY76BTWgkHKyqAK
2KGB+Z469gOgZXqk0yHJ3FyXc62ySZQfwCh23iGdBdF9xPjxHPXezdWBru8LHjNe
DbHWNO7pnWlrMWQyr3hh6HwBnroZnbCiis761paDBlHiyx3Rctl5oitDM5IjUwVm
KAlLTGlG5axB1RT5rfmsVlvRmHPDepA/oatRSQCwnhVUiV7oNkOaZcKLCN6Bfptl
YHK0a86A64gLQJM3bSH9w+7DusHLTy5/K+/oPiGLNhc+YbV317hWma1cJSZc06Bl
et0Hkg8lYmY6ifrmix8Kel8cKi8TmnlDQGpnfhi67CxiWh7r1V40msSuucLhbPa5
lpwLz5FkSKRMCvnupUKA3zjCDY4QRPSkYRpBtxY4dKOv3UAaMSgcgKnBISJsjrVm
IMyhhlAqlExljNDOetLjRA==
`protect END_PROTECTED
