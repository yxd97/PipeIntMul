`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xYu+E645WHA6wMWvU9XOWcKhFnLHS3dcdOsRvBTV8kccH9oN3w9dRRuLbRiZe8nt
HcxsNrESpRmqB1n99f2gkKvaW+Iq/rinU8Zp/w+/eA4b7x0Lx4nJSoIid+s0wkZw
nvuUKn1CKl3ptF9ywVn/KBbK2zQFv5i9pqYepAo68OfR9dGqBWNMpMkCYqZPY4nO
CIoU3IiV0GEDCNZOHgepKCuEL2k2eOPYGNSaQI7FoKc9fxbVGbWAPWQ0d81pEaB1
j//YslnT7xJSN/kC2Tia42UX8/gG0Bz9DWdlYoVbAMROR3IWE0WhBg2gXFwp2AMJ
gIuiIFLzVU5aQqvYnaSMyMmEFk71onk7fG3SLxay8gt+9joSZvgH2ULIWATPV7ZX
Jbn5Y9xMOQFaJo73OEmhh776pmePpC1tlsVc/wXygAOsdeE81P3GtgwoXaAnuo0v
SWt6/q+bo3NOw5aPuXzdvC3Z+dV1zqxfjJQl9soUOeiZ9R2tjcQ7Uh6osa28OFeX
538YCj9nEM36nur4QuVf9+FXsepdyILCgVWEUDY1CTX5iqP0ZPKChzKo6TSDVGf3
/kajxMUclqNDru5zOqodqX+k67+KKTzxUsDEDeUWQGMkxLl8f923ZDYG9t1KBHrT
7nk4eXOh3cmfkRT+DTE7OInGMWhSefxCD7biIRVk+/EWllERySV3NPeNu0ieGCol
YUVT6qdqfF3zPlJqw1q6G5ZWxPZoA8Yb3in38HtVMRMnRvrUabAtc0XM/T+UQPG8
75ayPdWsWSa+zJCMKFlEiRqcDh+14xmZo8e6TI8k3sHm4agHxxdKr2DOz0fFxNwD
b6okhOzDhbeQZ0CsDOK6U149i0XXRnaztqj05LifSJEGmdQv0ZHppQ66WY9h26yu
rLHxk2PuFL439oWl0EAVhSiBvT5QoDOaqH4mjfncmUysLWXHujYAEkiWAscecMog
zxiYs5C8RVrrAwkj7buw7V7axnQEHpcEIR6auJG2vBtiXMaJe3AOkL8qcI9SaXIi
F3tiu9NaC0nOSrJm7oA3dsdoA3Xd0m884DtKgejDBioj05g1mQe9vTCMvBZGSxWk
P9FAGgWIg5aJjZEDkxHvq9zQ2vrfloc1HmKztu+jDLX+rGnR8rAuO7jzhig6/fQj
`protect END_PROTECTED
