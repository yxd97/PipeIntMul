`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rdZGiKcZqO90/y5kdaTB8+rDKzMzUlet+sorj5jR4Dn93zHxB4tnNnsuWwNuJvzm
5ZmBM0NT93gLvl0/cVJr//epUSv/DbbCN1DE+hBUy7DkkiHvg2OBfR1ZmsPpn0If
vrZlXGKwfvVESS0ZQ1YNvALrO1mCboLZfOzS3yM6uPE1S0yATCb6loJEt60SeXOm
w3J8ccAij+60nUJqnJHE5/+E8GlcqmPNY1cztj1wHesXO46vTJdz75W159nL7Fv8
/uTvlpw04P1b8r4oNyrrLpFZTogt/I6HJwB2C13rGJea6w6p2Mt1qisBv437dL03
UwRBxOOKghU0ZWE+YCBkPn95b26YPD//VvDC4YCB0c7Z5EyK+/AEhLU11k8Z0Ecb
wq5pDM91lnv0eHAiuCH+sgNwcUfbohuT4CuMuaxMksc=
`protect END_PROTECTED
