`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
abW9DQuTpI7rBkcL96tboBUQmJ+b5LIAV0O2UKFXfNVQHNDdgmKP0ASqjD0FEbng
MugBzWgXRSRspzuRwR6jvIu3xnaa9xAWOxAp2R87si/dPIekuLqH8wFuvKKNobc4
qCcIr8rAMTiTsX/+DD9JN18e2FtTgeXvEWQNeQ9bQk1yfTu/THfE6JyQx3NtDndb
Utih1NJMvO0zLqmKZNR1bRVtjRYA+sCD08fsska3eknQO1HWOrs0bUJtvj4kdhD2
OUI9N1OjbsBcop5AYLedGOJUy1VsICYqMQvSfKdzM8b+MSL6x0pN0JSRx13kTZFp
2cFiIccfg6vuJ9ICU4xxdBi0unFaVw+HBbVqLwGIUEHimlDtQ00jfsEvrKv1Oj3O
9vb4GMXxn7B9zt0hsQMgkTqX2GkLk4ZO0CavYIZpTEhbTEuEpbtAos3ZE+VOGSY+
wSPKh27LcveUiwfwES4TjXCxhyhquXeigDH9W9W7nDaK0HFjasYzMOs0Yn01jHC1
rg+DH5rIQj1U2xOy7kiwwhouA2xDmexWYYeJbkt4jlCumVFKxqarIh9r7FOKz3D8
CDhHv65C6GxbPL/aZ7djBQ==
`protect END_PROTECTED
