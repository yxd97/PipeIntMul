`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+sxPeoLKAoOEZBSO5gD+od5Rxw0Y1uJToy+8hsOjtRX4O1DNp2mL6jylnWWjvbCt
A2txJ/+DU59t/0dWv6oXAEmenerc99Y3bGVrl6ChLDl+06RTmRytNyHcIYv3mvkY
ESskwXBc6Qsclx2QyFHqAMPcAtDbZ9qX3lch52pDXTiHyGMKBPNyhkWRIPfrVIzq
sQZKG1sLFeVOPQrF9LN25mjUso6p6XclOG8Z8Dck72CVxn3BdVggCC/lTNydLoMp
0mue/8mTLWPAiQEUSS9FSQ61of3o1mtQ9w8cqX+MpGCb7T5aohHj/imrHyLldHcq
8G4rg0qSfZFmyOqJkeVoI7ndGerZRbb0COxD7cWVQvcIyOy0+yJt9d75sb4wqtcN
pCvR2UBnevqxd8jdrMQ0d177V2Up0UQVJAghoW7vqlMvb1Dsw2/upExGZtf31Wyq
6Y/0f86qgzHHmnMMcq/vFsOfvz7O0CLGwhlx4j8dA46JRGItfayGGpDYv4IF5TNA
cMfKmbJVU/bdr+YBLZsf1iLwmaFDeKr+HvobGH4oj1aGo/IE3WZliBSQ/4p8/D38
wH4C97UjMSX5WepaLvS7ggwG+ygZdhaVmd2svQgdOQPb6gQRHDRmG2Aeyfc7/IjT
B0WZRLd5UEmsQJrmoo4YQi2f5QAGla8OBlLSKPttKkBaokWoInWTwrR9GVzD4QdI
ZKNXy9knbseYaTr1VuR1cw35EZbHoAXkNGsN53geZ/LFUgEvc21CVgaNkkMwuvFQ
Cm9b4lbM8R1ICUSd5epyxxkkgqbjUzRMeJ+5BoB+OAO1bkHxMFjkVelM8Ym4YBk7
ShYj8I25reCveKFJ8xaeTKgkvCwh5OAS//DMO/16g01bEF40Htt9wkewKtVOACWl
9/yEo2kx0azVTnBzcAqFpPGM2X0FGiT778x/Eru1wC3aFwYzlcsMk181iQy0NLIA
ucKjD3pfGePaowhpoPYR53kSaW/poNG80i7brgqyUqWWiO1EvLclZm70cst1yTKd
ruue3JPCAJUMm26UyeRWDnIp367IllJTYDeQYGRhvhby4cQSBcrzYECtz6wHrP9S
zOHzzubTopE9tZacWdYyxzchpejjsaHY7l7fbrYsZ5pinzPuAMV7M0Fz3XvykEvF
PIW43oIkStwaQlnxFmG6LVcnrcEWaVLKPHPhm523HwxoT8YtXzDr+sXbs7T8srYV
D9Tmn7qD8wXQKCS6WrScWmaKzpk+8+OkcjQg6ebxVdIZMoZqmmtdCkMMKhXG9niO
DfNbcmHw7Fz1M+lc2HB4iU60ykgSuMqbGFM7h8l06h9mJo8UhpFWZwICecl/S/z9
Bdo1+3eTFKT+Lp45Jgk+P6huS2u5OPIWLpWOqXcjQatVS0i0SSo5Yd3avMsjN8rt
vgHxe5v7gb/EXInupALowdRXPLlxrW/0CQWNd6f3vFTZsX5hTiQ4FYfl7vRTomLy
3n3TlKgvB1T6K9PiXeFj76sTiWFlmoI31AjQkdB5QHIt2zQW7rh2CwchAL9EpsiJ
eGvysViQ//o2XPysyYjcboyjKFVLI0HxvUy/FT91HEGulneUFLkqTKxrKcFIEtgY
Xie/Gkr05seUnOWyRCjFQOWkrYuGe5TFVXb2it9kJUwjHq19RjugvzPEfPIopeG6
3X6M9B7v3CJkvoRUUjcWJLvsIi7KCeMCHHk3G77QOmtPA5zi60Q8NqgkfuEyS9p8
xBvMyDy4MGwTmvJX/e7EPLqH1mK9FIjvHbXT67DsC/WoyYJJFPBPNkZjckUh+FZ1
la8wkhrcmHRwoEcvuZMfyV9y+IdZYjRmF+kmhPPOuY7LCnOlc8Hn9o9UQBU//uWG
jiXsMS07YsVXr7AF0e59mjK/pnBUCrucCKPho7JkjpnS6tay/iYA6Ak7N4bSLMmu
JyOCJO1d3KCBjjc3QgBIeQjpRY7ms4imEa76EqqpCNg2X/rJNwyR0Rg8Y+458fPk
u12CUu5zkiZKoq1NavIrWduiRvbyr/eG2nQdGkTSPVrNLArXtxmFbgSWMmwCjHUb
1tlpcooUXJLM3YpQXZHdfkXHq294QTs7iucLVVxMrcxF/97aW5T9mopIEga2oo8p
YPRj8edouh9uQl4vloTWZ4Re1LQbqbEVAVy31RAciqjFmqKau+WNCvx3qNfaCVa3
WP7lrc5bvxZSd37oxjy/D/Y4E6khbwdznP/nIoogegcZxQsUPXxfUWs422K/88bL
GnOcGgpsVLNicMJgUm+VtUtGiliMb2NIWK2EEiymdt0WlqotWed73UTb/W+ap7N4
da6p2iUQaMR+0ChyYzchi0dLjuYfsbeAA0LI1CKLpswHoxxj1nD8Y/pnZDnKk5Rv
HTYDAc43YE6iv882pP/lKjaDJ+l+kVxN6XLzjPziUuGxjV9ylpOrT9xlECZJ69E4
Qk3PtszQgnA1GACk9P7J9ueHQtGdfNpDJ87LQMIkAEimpBuKimiTqBasuEKWl9os
BiaiiiQsFJQ7OJ2RdFHTzC5v9Uu+zHSpBtSkyBDK5ZZts9QP34WTpUaaquQTLMNh
Frktw6NPg7h+t+DbSpw4zoyw+l01/EkNJ6oQL4SKADulggi71DMhwkDeAci7eivh
uAHzyK4L/bcQI44wExf4VNUvjvR8qbWrg3c4B0Bjg0xspa/sKBMMiTJ5RCniqGok
HMWKZhkKw3N0lNV771ynUnvVH9m3rs1L2yz7Tz0F3mgfI50BlD4ZJrclYt0BA2Ct
tLDWSEprrc5BGayE5SjJuFqE3BvHpr/R5Ian8WKa/ilWjqpoPCV4OUP9aNVXhIAF
FrO+nGzd2G/sNPqGAMYh/SxFcDarmze5rTZeK2yIIb7tRGgWZMNtqUXqlKpfVgD8
saEN2tNjZsut4SKnJQlkgtITyjE/vUNAGCDOwAN4++4qqCBqumbtifp1vjN4swIf
+TV6QRj5GBDhzAOAPUBIxMhYcTupdK8AjiWYkLsQ1CXUPO9WJhkKumpOqnLBZM/y
XOeuYQVFqU9MKRE4WVvBwqli3Rwlmpyizk2DXQG+w0FoZxUYw+R434O+HUfjdkpG
pczUm8UzhS9zDkuhTG4gTtsZe6rUpJYsFV2AG+17LPPSM+0rk7trGf/l9F0CWbMb
XQBkTqXcxB6H4d28/SiMGvGfHUfg87ctHKc5ygsvp50RlwDjunTBbATEnsFFUImT
quEjLESqaasiRED7XmfOHs1kJSbW2+rIOCX8aMLVPvSWrhb4MxaMr4xJRwqK3NwQ
iLRZXq1OT6WyZjH9733QfxKlJ1EF8V2q+Xyl3FWHteRcV5CBTuSpuWHkliEiVhA6
WstBhmmj2LUDhMI8E8VuJkzUVHeC7JzUV+NpTIU4Tk9vEP/iOykbx6wcg0xxeOTA
VYQlRlnmCS/6Mwse7IkuMH99/SOzBXqyc3xAO1y7oKx6DhoKnFXIcA2ANfAr2PKI
qTVK45CaMzND9W0blpCo8pUNUPHeWlxpmTX3LY8xDptIz/Z0Ctz8rHnHxzCW74Mc
0NmnBjml5SeQ5SP1fPRfvifwd/AbYR+ylqHdxcFSs3Ew4D+feTSWb9Mq2m78pr26
IgU9JXKURjD3bpAf2XO294LjN38ewjmdh/YDq61/NNgC59vyo7mncMasXqfF47nh
WmVHn7Ubj6yu8Afghi16STfHw/iWGYJvvXpBo25lanF5SpgdYsDBJ4nJGm0E97PG
lsx90tKkEZhFVaGNnpOKLs0nEKkB3ZCtKzSUBXcQBIPBpiabh/oVe2xUGC9DIEpp
RtyF5uIV/06B59zoGJurUAkVfEs+P5k6wDNKscnkMxQkpcLvxhB9ayRqeQLbVw64
HJ0YM6Zzva+fBQsMkz5z752tQKBJQvP0PDINEEJSzCACVld9rExWgEHQH38FO4vy
ESd49TnEkAvynNqy897GBSwgZgYsY7gvIcL+6Zi0I2SCpf9PlRZZPdGZObkSiESI
+gGL6YeM/GjHGPO/wSJ/dZvAYAQJZ0BcAEdmzgZ/97FaWSmoMwv03Sq8DQQS3OXA
aqgvxeEhOs4GmAdb48G+MHMdfC83kEyuQerFzLpbRrBnE7alpntUrUkSgx7QD+BF
0+S53U6ZUYPDtZAKVN7lyX8Z9Cm+3CMFkDLXx0p6bqSg2YZYDbq0z7u0ZM77lWGV
uBLjkGjdI2hvcmwITZQhWCsybW4iFbwQgBSlMA3S9y0vMGq/jkkeSQ9xi2IdhtZ9
OY7pNAaGLxjBus0M54c5DqGGgrSnYekWkqR/qX3LkS4b/2TyLcjByFA1K2bdzwrm
A459Ze8VQokIUpCi7oWRAAHpG3GyY3zUY10Yzg0/qo85EvJrpcnjx1qUc6lgz/Go
Ecdlvs0OhU4azzv3WhedDtl6k1GiRiuhZ8vmU1rsc28aFT78Oc5QNw5p7CylJXIx
qfeCe8Q6UatSVEnMxLKZqUPjcMa4HWLnp+UG5An4cYrYLW9p93WsiqzjInT0faZu
7PKK053neDY17tEt8bkKPcrAmWfLhgEaneqWuZnYVflPEUpfAhJ8pqJDSmOYfD/y
uVU6vIe4kb26MjPComPGmWwSAzzUPyoUU+1MBojGocnaNocSjKjg+hG8cQRhdv6A
i48lzmbH5WDmWRyec/YWB1wBCuxSCxUxvRUXUBzaFdFS/dl2tsC2cKpxg2fJFgJQ
JetlIdUtQ6TFKJr5bkC4DcVAyhgVPIKhz7Zs/DICnALJONDrXD41E96pb1h1Px2X
90LZCZgza59hqmGy+7wl4N/3l2HUV+MTElYQFTb5oJyEAD0LGygsyYhsPgo9wr5r
u4eYHbzzVrxQnzAe23cTc3bChqnuMPS5VwFD73R9zdnv/recjSoljS71MYh/c6U6
JOCeIyWPEHwf8I3tJM677DAdOcMisMTBMkqBe7ErL2Dkli6zNNL37wvnexzXgEtE
yUoeHUZjD/pHEWsFQY6lTmbgtP4KdVgt0w24tsMJ0LvkJYTmOf8EbPYkflfsPR4r
cfqS9+IuwF/GFC6o/43U2uY8hxqH2SjA6eUozjFhzwIFbw3twsDbXlTDfNAFOYff
qjj1+uVVRjuMg+46gRVnUELjBeJPv0UnoDB3B1nNdlrGQA6agRPTf/Oju8dETs25
hp5iG8jT5YAo6D4Adz4hSJ8+EGO/ISjRPqFkH3dZOMKHGztttJxejhMbogbhU2pI
as/BFJVG8erbGledk5dIj+OEO7NPfU5UDDDDvkvrKReYlNndi6ZHy3780UAX/aeS
QDbglBE4b8ILLJfjY8eTATN9QQRFPoUWDkl1eYUGMUBVPAvgDNNWuzzr2OqL163o
Z6jygDlhRnBUYM3IFK93MQEntOiGYh+OI/TD3MFTBiT7AZJYWwoTJ/fc0V9DB6RI
I8zn6EIWaQ6ZpFHvGB4F0sF/wccsfktbCibjUGX5T2VVe10Z6JWnrcGeS/8v3ryR
+Jj6euWsQiSz9Zxv7K0lLifS3Cd0JhLk7JpJI0aYMiu6kpqvtidgPECagFSea7K4
o24B+MhkPs0oiICsYqmT7QIVLrnJHKVw+wK/Sua7HeaTAIX0AWZielNDGBp5H/OG
YeA/zB/J9HNzeiVyhpFPTFZiRRjs3dB55Dnv1T/SdgxDR6afGCVi+C8RMifqoD/I
Q+UvXnBm1/s6SPXNmn5VOGT717gUCNCdquFXKkcWRzB0xmr4ZGokhqNDgLD8IiKW
y7PHJW2JWnH1uVRbUP4UkpE8GeP2ZnVY6OuG2Bpg7h3ingtEY+okjz1nncZbTFs2
+EAYUNR/DsTFhwjUoT90t0HRXCjN3mY0C7j9dPf4fYLLdUUUGpiDdXPCVbctwCps
mJRrK7jiRd7gHHhAF/PDmnG/aY/fre2olXJc4DTm8Vpw66qsbhg1F7SCB3TXIvGM
ozFZLhazw1KdiXnPutFbIowqTXsV+0273MD1wCd9dpjiZZ7sXgqGZNZCh2eBz9r2
Ha7JdRdI5WgZCmZssVCUGtw6wyGLhBNG3PER03u58tEs+K4WLs25EpC6SUaO6rJI
UcSxSgBUhECAzY7Y6giw+IoO/bpW8On5qpuCV4hKah97Q7kZOUSTVkdy0T/wTlM0
JCRugJoNESMufn/jmDp0RRZW2g92emeu3/p8S5QLY2i8XRFvy5/c5+L24XOTlj7w
UL+rsazRzyxqlNM06oJzwRolMei/kV+Q7WWCQBkjSchW7Hr3ORMnf+PJa/8H7poI
/YdOAFE/w65sZ598zKU+K1RMlbWaYKi0ZoEsH00GnVbNxXLRZonpdfR2ZT7CB7wL
n2RLC2YHq3ndPSIeEIUThl7ZTYaFAHYPxP20KyhteXMNCSRQlS+pZCQlWZYGJjHi
2WSTYSolphMcFsa7ULDRn4qjhjTNVLZOUx+TVmO6krttmq5pruwU9AAKFDsexIFv
4nCwdXBYD8Wnzw/BmQOsilG+zKo58Ea+O8RqHMB8G5YQgnT5Hx68th5bW7w/g39B
MKy7hrvD0m1zlsdMjSAd9PG/0TLheFyy6QJu90+FT8ipRYEf9f+66uS0xau68fZO
kg0jRjUj023oZrhGC0MrI3XFPQLisymoTbjz3UXdK+4nZgwAm0CgsAd1Q9Eu+a3y
8g7GUoELDHC1YrfpKMbDKwAZcWws9c+EAvwAI3J75Iej6w6XR83XNt+fDIHFWt81
dI37o/3S7RgUGlUyuJKByhuH2cMHnfeQHcYJyEf3KFaGDMrvSyg/3XxMDb8Skfhx
elxXPH/cnuxoRdsfTWlMtKvZwpy38p/rfhpZuPHbNfEDAa/3Xxytm0Enhqf5WwFi
LnI+KjJgaJDWaXWKtG4SjCvBrEFwRM0MKEKzp1An6IdWQw0ROn6usMxajOHdVy2g
caGhbEdvbZVVuc2YhWbc5L/RP8OVx4XVkQzZJqDksIbBEGX82Uv4JC/nFKTvGmwN
3hguN3Y2jS285C6gQVcb/CTzy9AXqah1LBsNK6SIY7uEISJj1SpIRgnaZRWOoqHf
M7DRy61feASXJCjQGXpJtWrvDfwCLKdSdABsVHQup+kiMz8zjW//7ymW2/2GXybu
SVV3Pv065cKsd0M9HkV1XUdTW467X//FOHo5HwL9TnclIjb8UlIXcZtotnlKCHlX
rUCVpZUvB7v/U8VJvFyk1Jd8fEkE6PZeO4JpvaXbc4li8/GmauriZhXjkQ2u6kNf
+sAyPlNl+hzwHSlpZU56QaYUfbZj1uqCSGf3ykTr6fIfITP5mcqSnQAGbH6+uibC
kXf/sBbrarGuPq9HBiqizNKFJfuux29Aps0+wy2+jm0vku9EKawQ4vmoV5QaSlFz
xG60O36aBpJYf1npEFtMZO8129DReuOvJPEfUOhgi7Az84irPUtsW4rrNO2y3ng0
Kg0mHUQ9zyMCDAelE8y7dzbgTUrJ2KXRVhYrJLaaGz34lRNR5M7+OlJTPQVxke1r
bOKUbU/H8kcn8VFr1NnwFjwaBzDDm0tIkmSLYnLL6yJ/n+AYtMyHxZ2gL0FJiIZi
rATq37ohyYMO5FANlDj6DG32FAGm7IjByZ+a7QZGYDeZ7V1DCOAE7EdmoOCY5rKO
lAQtxLNi9ZySN6fvvQEHWA6PRwN9ZjXzob3TDWFKtJBat55d0ibd0FBB3usUzWFY
pI7iyz1qdJw0SQhKS1qsa5KtzEQqaSxq8rkt5kMTyuVX1rsBivXQZOISytTJWeZf
5PYekmG3hL4UqHKJJx9aQDxcA4XMgCACobQSM+cqaYcUUnzGQAJBOlLXRylSxrGh
UIHLpcHZRh/1M60isRb3BYSMX4w6c4fTw8P83RRMbpof7A9Bj/isTwaS1fPzJWj6
EyJIOCOQ1i72LN0YPQVWNYirkYS2X9a1LWtIxp4PxJKyR5witaRQfjZpLiRRMPza
VO9fur0tPaSySUsPozodrOfsA2Y7fjuZMDMa+6TBrgAUmc3mr1StyKxdN6tfqrq9
b2WzySQDD4AAK54TSxDSSQ3qVYdCrUNwWxPoVU8PCtZaABEvOJ4F5CbaNtI5zGiN
cy4YSrGXu1U2yagnD4rDQeXvQwSCadV4BWnz53SatSMmVpw4GEjhVJX97rzxHVvF
8RHhDw2KHSNgG51RNjAtQwpxvzz7AZzRMqL+OvawhdsLDoXYxWlgCmGgn5fUtYp4
/49q2Eci8vC7bz+4tNskJbGOn6h6GKTPAmckRCCrUAPZJEzIIIc06j9HOpO+CLiz
0S56/IeHexwTXGsp2Jfa2fCBts8vJs3Zh6ob00Ib93WPOfON1eOR0ixQZ+ix0ODp
XK1zdRBZDYLcQBEPu64BwsMtdZbbqDjgROI/fierou4nO8nHL0hxyvYJa+VzoD/M
IGWChm4DkktSCkV/Q93KZUP5AibmNUeIUyQNgeiyCp96nc1zRyus/0nt4oWChLQx
9axJZZPWOUWOlhMokWktmJoblY3JGFVTSKkhveJ+MMQlwoG+zxjGwhJT+GD4EDy0
9sKZgBQ2ZMUQxocySHbbhFX5cONXKmciRzlJP+rP+MtVRWxq483eCWguDeH+wh+f
Rm+qOROunfFUj1JKkj/kDeVLAhjTHf5svxnx2T3Ic8jPxbQtW8ZT47ZV/xcOQ+Hu
PT3Nj94nAFhNkV+jrpRaNKZidM+lylMMS4T17CUzc+DFNatzRoemIkNxKkc0OKl0
HJKFstOwrIk2U2NlvQZO8hP5LyiO2jRLY++t4MDkoJYL9QXTFDUSTkSoKumtbbI+
VOxQoiO79l2p3jiY4DaokZicQ5XvqjhkhcVhyhdom5GJZHULCBDuZ+ZbxxUWUH5B
0aN582w9AQP7kxkxlkg339MiIz3/0ja7M1niDTWhEqbKkbWBnwQbC6RUVGwNqZbO
3mf5sRLBdbEPez1SrIJNp3m07CYRSmdbBy24IfXz/YvTV68WkvahwTqLhivRP/cO
Gs/gtkuVH6lnZ+ScWxca8vDD36kuRpFUG0FAiPGBd8lnBXHPN0GuYp2l63vXVCrC
V+g/e42uCgH2dLdw31GRk783ki1vM588WWxyVaSEdiVugxIZfeCAphJGj7yX/Ej3
O8gWuazJGUR0aroaQ369W3VTEvEuhVdVC+kRzGRDxFxqDbnT9ZYwHlW2uKh2ebdI
KSCfuTtBf5fPFfaX6ITbeS6whdIRWQEF7xQUqahY9KUp5GZ+3+wXJ/R86KVfyYOL
/C6abOIqW1apyy3vlHybRkXPpVAXTBu22E9GN9p8n2zIvuyzsWfPcnLzXlyA1Ukm
niPNaVKuAXxJxCtWmsbH0uXyHDUNThhup7IUis0XCTOYUSle1QVbAsWu23rn7eU8
DueLrB9sOCmpb9qSs5E25uq8wRzIdRACq1R3xexCtvfPwZxxr3svhkyhfghyACG5
V5HO5GjvV+yWf9oQ3S+lUctf7+F4J8S8xAB1KgxBPGgd7jo6S5veFzEI13RGeUyb
7+5g8VBxiBjPlRFWy7R2p0nucXL1IDqnvEziSaMULTRAbg+StFpmu1P0gz+Zxgqg
+M1FtQ8lnVSxCcEXdlIrFy12VRQDjRCAS+gYIFmmGK+3/qw3wv+AAZPtM+87ek75
ogmxQXgZo4r+nb499mjoZtXR7Ofj3TvuqPV7jXewfTifWmvA1SX4mAeSqi2G/mjb
19rVFjQStUi8Z1Rj8smrQvSZ2lKR7pF22t3/JnzUY86lsJqmDEIE505jcS3JJIEx
UrgzGcgV4pSYm01QovEtMo9blczn4IAmCqoQ3vgFaKyr6voe2mFxlfxYfEMZGRkx
YEcbv1cGRJ3xhf9/hycjjDCkamPExFHLUZ7hMWrzTTBnxjGW7Srfu3NXVGjZDTlk
FZfYs9ca2vS4DjA3pLSI0U3nnOVjiBWZap+RJuqAg7wQgRJuoXtPHpbzFbZ0PEIJ
0E2h+zeSG0kUyEVDGtDZcTMtTsThzPsykb2ZXvgKJ1XYIhyJM3VzsaxRyOjyntae
13V5pgPWaypKo6ZOr/fqemvmwQpoh8B1WubvhSQuXPztbXT4OcJgXCtcmeiBU0tL
KZAG5p8hDvD/XAyTF6jv1DDEAsR4g9eEP/YHg429SzcACnrvcrxnyqnm6exp7ar9
gJPoHa1wQoaKEHlYTieA7Ga0lqHzMEwSwBI62uJJx+PQSigL5hpYB7bZeK1H3VOl
wLLVHkuftd78YkZNoVq29YfjU19oYZ+QesMWLsvi82+hkjNq2oWDElrz7hDyEEAn
Qnu/yibfQjPuu9UNG1/Z5EOw7Z7G38m6AH0l6wfmw0+3aIUyzk2sLtGW7Kx4SsaW
qIomqosGfS3C8xEkLpBwkPjP+nKmhtLGBCGHxxnpNAXQeaOP7uOTU/rAW4xTaNdA
ulO9lb83tt1C7bHp5Oxr7YQPJc5Okkn8UwUf8DhX77xYlmTV0XF6OHTFCQht0r5S
8sx/slfY8DKsvwecpSrBmj4PgmA+68qJJQTADQn6y/KmaWIJpgLWFywLqF3L8yWz
wSp1XB8nQSkeqJmhvKB/D0fu4wg9WbZY7MHbi9YShMX5pdQGSPQ9nlx1P/z/viUL
GGgoqk6QeP+37Qb/uuyHPjpcZvaMHyX5Ie4iRRbRyyvWMFtR9Xf/rxcn31oeYvq8
5dEn1da0ZtzYul9ogUMgx7ZK5TWzyyjJO9dk+qjSV9vM/Z6WxDjE4JLZv4qVIDDE
m1eG/zLnzRa7ZCPAKm9yl4O7dwxB+ZyYRoybuIYwpPw/jxfkoBUr+JArkKPOYwOJ
FeMpwMexFAxhYJjy0HoTJfTQuzZ5aJO/Xcl38yvY1rcKgervumst58N/AULkUKNB
kUTRDhCQZXPk+rioPUzb864j1yeS37EsfBskrkqpWlTnf9z8eJuBzWTv6OZqouIT
RMHq5r0NF49mQi2C1b7zBkQWByztfemq6CMXRR/QokccX42djP8pr3AL+yz8G554
3v43N4sET3HKFoB1uDgzntrwTe9nwCr2OctKjt00LrWPJ76u5yk/GnGYPgFfPvd3
VLRgOgrZJD0fPuQiPL4lf3TvhIMJCLKG4SWWTNmw7GO3YRjvQVZduU5SASfkstWd
GrJWCEotvsEE4LUUg9PpelG5vOcBmRhaE5t/Sgg2dkZaUnILrcK0U9vqedGCZd9U
rmBi8/0WjenVdqftBVyRoW4eHIfufbBBdys50Sydui/hQnXlEXr5Pzsu3zU4mvZR
RJ+rlHVYDjy6QJaOyyirKnooYOk3m706DJ0+FHqndchBbMO5+GqtZu5sBPHdAIGC
PJfVknpAxnmmHN3YrXU+PgJU+lMYydDWBx9lJdiRgDtaCHl7DosHx05RfaBXKZZF
CWdfHi1YRigmskrLhbiZ4sH7ml8fnsY+5sie2ys6T+JV5RKdHEBzj5bbn7PmeGCQ
k+b3ZNmdJFGyNkLH37Jde+qnDcDZK1xsVlRBJcNFdoe35Y3xPa3OxmkmwRczWjAO
h0CoDs3vcAsAFAIZCjiG8SaMzZHKLUvOrfDbiB/yg8PNDUn3wMSCPGi+35hG5THj
/PVjf01ikuaJ1K5otoMTxPy2QFSwYm6z+2jJGvl+3ZmtvmWg/fpE5ZLzgcIZ9qek
5JQsSC1kI9WE+drenkQZ1zVb4wixjoLLo16uiXIYZad3jniTFdJBKS7JbIgnzPxx
jkUlHWFdgAf2Z7Pl2S9IF5/Wfi3elO4AAxxRf1DyuP+b8Q/xnNbv6TdI7Xo7om9l
c3zuNPbh7VgD/w+R5AbpKEg51pOEejoQvuiEvcNBVtT3dSs1kQR6AqXo5+DKeeoQ
B348CKBF/2ZhayF8S6Nlf2Lxl4OBXwNgjHgIus26WduuTlZATm1AgvHI6Kd6UjGT
9s9ay9BzcQMnSrQpnGw7fl7MGuFPXuYys0350q2qsQSOTXhVj3GxOvaGpY0ebTSU
WQfKIXNFG7rz8+kJPLFWCQvc9TyX4tzdUhIsPg4OoIAS9GSznVtsfKaWdB7MS31l
eNqCx3Fk3v5Vg1GxjGhJnbbEKyIazZiH8E0ydrndbq/ex8uWgksIrfg5S2KarW8I
ANAo9uVUAjz3G5nMXZp4VbzpSQy3+dd4jWAXAmmEuV18jn35cqlEnD6L69Zmbz7A
yjt5HMrJoUB4ox8Vs5c/7R+QFAe/fp05/Vff6717sqLL4JX05ilEdrOCcbKhkvGp
a9AlgWOqf7Z2ajGulmC3Nk4BAzkyy9UUft2oPvdgnDyNmwddjUAHiL9EFZabMhEJ
mNmLkWJljG2ktN3S6ZqQZno9Hbff2jqc2b560F3H4xnayljiDyENKVfWunENJKps
isWzWO882ewVs16/wqmPYCObBv/BOmBdjSWz1lnncbeXyUgt+0oH7BY8ak0KFr5L
806KN1ltxqnSnt6u4zfPrveDDmffi2bYSBHLZlXHnf80JPm7tIIupWrCWxE2c/W4
9gjOZ2TO3tCf2C/V3aHmnSpHxHHrhUSu0mZ04gUFS98eV+oUYKLXRlwEuSw3QDcS
OQWJGm6ZOFvhNsPut9XM3Nzy9RqQGMFYTrPuolv8b+xY4YsUZwnOYkUAFCSnDpMY
C58MBa4paWENuT9NZTTv87cHbBiAxJYqlzFwMTkNftTMft8Mnjp5RytSS6wKl2R3
JlcRtrY7/4PFxhhhkg7Bj30NH/sNzpH6fY35FLby+dvtozRpYVf9qF//625j1uaH
ekQT78bOs1dosifszr5avVOMrw20f2+fZm7l9ReMH2TU2Jrs66np0jeRis7PUgkF
4illsC135t0gDldO5TRVPestdaXXPWXQ+gGn6rb53dlx8XAZcrviOQrs2y0EN3lt
luVqtUMnxGDHz/pE8GeoLzw9L0R/kpBKiRzlRHmuV+yB0sv5j871x88siHfdg01e
TQs0i/jJWaIi6GHU2zYBSSE5fNBMKwW/zBampLoVITaaWq6V5hdG8lc2h0MdCERM
1c7jc/549ma6a7foZeRBSaUaRy3OARPApripFYsHQhoXkJf00gft+RHD4XjKqj93
aKj3GkS9fTi+rArTCrev+RVFeeiCLnFXqCxu76QQDJUxnQXPjDS3dkFx4dsgQ7ah
8NwMwuyjzaNSgWRl9xlOfbTYfGBCAxYrdFwPRKwm1XMPHZctTf+FgD2j6JVzpgvE
osCeRpSnu355LPgOIcKWKDEevwR+RTYT7Z7+GIjhE545T2CgmAXRSLQrq7vB8RNg
RnK0uz4UXNVQr3WuFNBJvLiYkJD02Ujto6k5NFP4VVFEx2ohs/Fo1Fs7nrBcGtMm
G5NuEDjhogc1/3utC0r3R6TMXYXoxbtpzhnSNmuaj0h21A3JhX/dUaEodZ08XUqO
NtPp2b9d5qR+R0DoxXgmAglbkIn6X/khO8B64qfb9l1jmUtzDkEv2bFghi6tfWbj
S48EkdS7GoYgv+YMOKXilmmxSPkpnK2nlDnjSLUm0HYabnNcoIR/P/UWinNnz8DT
yFz7xTUqeS/QvxZtf1BwGONHKGzG8uN1nxIkOkijG8ZfaJaqUt9y59gIgK6YvErc
rWxr+IwxRrhVFil9vzkH6HkMuKyXLL5dp9B0EfhX4SmwDBSzZX20770pXFughFb0
Ttp+Dnnn9UyVg3H0VyHrhzE6Y1dG3Cx2n8VPQS1NslDLGVfLezYBn7/Ba/LSiISg
E0DhTWO3cX5vVFb+AwTOoVfbszFJ8f4uYLu+z47jjPipFON9Zd7B19cKp4GvXcfo
eE40tWdNxUTuVGZKNnGrRoxKw4f1sdF8UZQmWBz8a2aIZR1gtjFhZn9YbNBGCKiR
hMzFBLJvGhPkv9HLZ0bFSZhtQTGrHhBe9SijCS0bai5ldk1VT7Bn4Yi/Pz8/qJ7I
2QJXJQUt0W94G6GH7QtW0QR24K3nqcMGD2eoaXzMWg137tTSIC3WxPzDzBz4oGJ8
IeUiKhT5RabLPySAbCbhAWs4kwJlLDnL9WtsTMl5lC7iyTCsnu7OFF6eQIaOs0cp
WqxQ2OhKXHkh8FT906aL6jda1l+wexVR6ZD8LsZylDJ9/MrJyAte0cvuhjW9LUIv
AJ2L4p+hkha45fTEuyNOz3GqkfvH7HnEjBBqoaPEH9AH1IuM+gSmSL/Skb9260tR
RXDC7jLhibjkyo11Ds4/USk+CIsM2am21UbKnX4W6YzChc0MSNINEVWhxoXivo1R
/ohmkQy+EP/KLvQUpSPdAfMfJZF9EN8XivXuCLYP0XcLcWzAC+pRKyrYAwWEGPqt
T4puZPwbnDWsQiPTBBaovNdnsS2zcO39l3Qj63JzSGIjlDJno2ERiK6UHbA8dQ7u
5NGl9DiFIJbGOY/+TvGXUoNPXBO6QtGrcKDtHU1HlisEXfdTNI8Xe+WOKT7xxbWh
HDzrNBx8YLuWpTNLIxbGrRBNd6aoVUtyUHUAtcDZoK8nvW/tCpHMaMhlSd98hKBP
6dSOvwh+eXJ3GEh4k0ghV6nMy8qVy6uEV0I9NUKAQtl1QcuF/vFMPfIuCkEw3Vvo
niZsNqqwwckGKTr08GLP/yHrs58GSeFHM+eR6KyqKRUfms2Ai1TMgEaQxOUXKakz
VYUKK7wPoCziOhulmTzzJg==
`protect END_PROTECTED
