`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PNSJ87YoPof7omCBr88c6BE1opVufQzUIVM/VFD5TglwnQ/jf50Qnp0zkWP6gqHM
c5/MtlfznBO/0aGicXEPH2vAIafgBwKA8hwT8MT9aT1fabnjA97oY3NpDSssNRFP
wp1DSWPz37wg2CjElRJ/KmFuKnodscM9Emhnb0alpL1Sm3EcITS/WQfF9LgtOaB4
F/lpnxcQ7E5fuZBVLFpFAIpj8HRDa7qMrwLHd6MnbsoUdx+mouJM9zbL/HME6ssr
5O27sn8uU3XkCCrZGiz7ct6BGiAc5KN8hnOECkYDhlFxzcBlhnkuEKDKYO2wROSu
d8MNLikVZEzmRdxb2QXjEzJhYVVejD66k/wHPWZ72wFUwrmYB/BVFps1Q3h2iwPz
gyLxVMctljraQMeHcFR8syaMivQFyHwBlJYNGgTR3Njxsn3tySY9OGl1QblbAURO
sOgXUFjbKgqiAdGQYEOH7gF28sbnPa8nJZOdq1d5RLihXPMBmuXjSBRsnNKZcs3C
`protect END_PROTECTED
