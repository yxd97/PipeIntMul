`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g54LOkR25GkiyiAUH6WTnd8n5IOt3zyt8Zihg2/29XgYfKXdCK2cNOYdxeRd3wdU
K7W/4YNMyJu916RU2w7azhnH4RkaEe6LXqNe+eOK5qZuw4MFDXbr6Y4lGWyeyhrU
OvLsWUzRypUCyyc8finGMXKEk1ZA2Jtj7aRD9HAg5Cd/3R6YxET1v2LDXvdC0Goc
1gjdP3h42mj0YCa+B8XSx/Vn0Fkr/IMeyRpNlNLp8D3OAzJ8MMN5+DIRA2ZwsTwG
WgLHCqLxM0LDvgGpJEPwbtKWzfSUSDEl40gfTGY+zkOEKq3CSzr+TMSqPe7J8HF/
qfXBZTtJq3mWUqB3/QSBnSlikKEsjvZ5QS7AU0YDrPsnmMYc0wFyJEyR9Zrb9Po1
1Ccinp6qaEImUU6A/1Rd+mLebekhigK5wHt66fJnFc9fKA0shXBDs2PxM6wYYrjn
TXpQ9d6GeElinGDWfC8PRuTkEbReKyoDE4wfoqzr7RQvHuG2wJ1e1eFfPpLQjmyZ
DujGJYdnK/f3PI+fnH/2B3cdQujlRdOn8zW4nr63djDgGkSd34sm9GsgZv5DRk3c
EQXfdWTo1NfW9gbCoJeNqpA+B7y0gUqBytoQSKnpREqNLFw+4IiXz2LfoewTm1Hx
rprp/3Y8DjDW3l8l78pwRL2IebjIJD00IBDzGMWKNTTArN7DyeVZXXQrIR9XaII3
igfa2IrkwogzZECZ47bZ/YY0ql5688TPr6t0HwXBA/zIbxKpDogWwabv92TQQOC5
8atWZ2GeeCLLcf530rPCdMhiy26+oKHospNfbM65E3xQmgzO/hJVq2idbca0FXOw
GVxI4cFZdOHnpvpRwBQguxw9OdSzmlsjzkfnUJN9s/YRFOP9FMHWNTkNdgKHo4Ko
rwH7t91uuNdvhYc5QuHvS8U6JQJwpfn9hq9OB0tWE1xFRusdb5OiJMrjjTcQVTB7
plhda/wfxwTS9X5yrN45W7a9RTaGY66PdpiuA/k3+GqdUbEg3Or/ABpxlTAmF5sw
QK/XlFzUDDl7f7aaafdqwUIfUvB7jr9uIvj/9008+fk=
`protect END_PROTECTED
