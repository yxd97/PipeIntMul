`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oaDvta3+SFQbw6SF0ejs2ph8/QawWGEMEt4DZ9UlI3zpT7wKoIVyPWTICJNUf3T0
PZFMw5/y6PpM7Xd/yurfBBaFOQRL+g2+6jTBZA3UDgiaB6J+pS98a/Tb/cv8fgVU
nHNboYtAoPOBsEp4N69arKdlO7IvwN1S4YDYsNHl5ug/HNbSCpOXU9jmdso/r5gn
vVp8RO+Lir63QA5eCmZvzI007Rcjdwq5+KuWixy2vNvnRTA++p+XLB83Rn7bA3Ge
7CrXPdhX64yNJPF5VFzDoqqAOOBdPVE5YEaJ8s8UgmRflOld8rGKclbNe8ZVU19e
NgXwt2VZt2cnzAbuV9aoKgVh2x4DFZ2XIWuofUVPl8T0qXJfrEynE+4BeXuwkPvY
vUHBoIy2TDmug+zvLJ0Sew==
`protect END_PROTECTED
