`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUcpEPbDeeSmXNPluq0u/ZWmJDLF6+p/6QEv2DYAF9mmlOUFsumQtRusCcQLySmk
F5Va6uydCirWdR6vBFI1oT4qL5WcF91BiTQyiLrevzDWf+90W416pgCop//n4ZmD
H/60pHwPbDXZ82yG91zg42Kufw1ClpEt8DyQZRnHJch7BeVYryV4lxI4i/uDEB7H
6iH747Dl7WQrLwheu7thFkuEQI8VKacX6snf1Vc5+0QMSj66YvwhNv6maxe8rZlY
SvY5gzY14tmIiA4Bzelx4g70IbH+ac4SrLH1JLglamkkr4qHn1gSpVtPjL9EFd4k
3doZyUFobJ6RGOYoibMc9k1Toz43NGIphBN1sdi1yx0UT/roDv1UdTgtEk5yqydn
C0tZQ7YZryfs/7YGCm+o5SInaGmKEg4LcE7ZhCo0oIZfFbpVgYlTn/gfxzc/tzv6
9zN2rlAgaNEjK6mYPVR+VunvEyNv4co2Pz9GO3+zxhC5gWaJTrT/xWJrpkfCw7sX
SBsHOoK1CVja+9owJxBAZuE5zmh7hh9U9H5qITcw4PoXmRyYoQhOOE0rsLe0nw6Z
H45o9pfbIf8jF2Eju+twIKWb9PrRrjAvPRbHbOKePL0UXZkkDj9CJ42yuyiPIwVY
90a4XiV74H4U1cZg1tIjZuMR9BnwajyE4wnRAq1o9Rpu3y+TNWW185MICTK/OrsZ
+Rt4bXDOIdIvSAhd9/dauP6jmJU3zvDPjZdFY/yg/FHKpR3o5g90bUsLXBYDLCav
kG78WkXJbSZkPq8Mf4YiNHZBumqRACNxlYMiN37AnujmmiVD8Cg6DZfDE+YPA4xx
NcJCT84BS5JeS8Il/ghiXamoYnNoNsby1ylUCRDKvKBJMUfcn0iqnSvJxPiLkuOf
pja3NjmsrOwxGsXfpkuYwiqtMKdl+lOmenQMHuo86IPRl6PMz8loEduB2QiRGV40
mgb7VVP64FtJw/kHY4+oKOgHgsy8u01CyION473Ewkx+SlnXktiAlZ8hjrdM3Iv/
8CSqQGzE8I+X+d4ciDTP7wiBBFf99m7OyR1TgblFX+lX7XuoJQUjdj1PA+0j0WWw
xgDWkOzWW4kojds9/9ol7Zd6rsRjFOA+n0N6nC4hOJUtVGukvQVkN01HmW8fyRaU
2n2n5p+eifC778uZU7MI5TIBXOUvQbGREcKwYNIF6EqnVP/T65iWguZtRk8pBOcf
0lIN8nE/hc7C3jsaT0CqZFxoxSwUgnE2jv9X1+6m/Lt+PXIOhfTpZ++83fNqTCoh
9IJIdhghWEpORwEczpZCvRRkKNgtHIa4X0UF1rOcQQV4IBjKfmbRvJcR4nRwcaJk
0QG8vwT+9ETuTTDreqOPYTkrQgRC0292SyZ96bRSXtnvkDnBn5z4tLHLsXaGTfAk
4MmqeYabKPyUKWizZg7pVKw0euWpcagVoCbfm0fnb7qc6X2RI1JVEHZhyyFMkomf
FABVty4VcS9TYE96dbxfm8TKkPJIWyISgO4E6lZoDsKKA/jjJyGBtpgjTj/zIGxv
n92wdpXV9+0vRtmPuPKkI5cB/5PdMCx5PO6A9yO99w+TWVL+k/iC9p1V6Xx3WGr4
dOASBW+909ynUQ4OzNICm8JjHCUC7xqvPskJo7/Mt4qL56tqYnS3ohlv13S63Lkx
etLIT1cLwZN178mQc9TstrlvbkLdFobMm6EqA06+DxPGRKTVT7+oHRPsOyvTSATu
HBEj3Ktv266dp4kUuAVhVHjKi8ghCSKqC57gA7nOZ4DnaclpIVWdCriCJTBTby66
zY5F1mdC7+aQUev+62wuD1COOkRIcK4hjwdrmZORyxF83tyohWqjmWM4sdkeyplE
FdbE1jFONgr+aOvPbf2pOJlnZiSDqnZ1XQtPsmB0I851j04xNGHQ4sEP30f6Yf4m
h8N/E1iNf9sqt8LvkrNhWx5Pb7l1AvLdysqPkkP749NyFi/sR6SxYsKNfuTjNnUc
bgW43PDS6TrCSPoa2nko6/KWL8LvPzaRRyEVCWtqzXtdrm0NMq/JOYEfXsVc7sgr
b6ZkWgWZjG/VwUJSTEp629sAarFqTgKoD/EpoZeSXird6ulRtoFRcal8lXCe5IUx
1m6tEFdWkQPavj/O1tl999kE+RT0DaHdJaL3fMBTs6FocjPsKWV8Oeoxm0c8eS76
tAdl3VGUkEgYvxCycp1PoqpwrQEJp59+lqfaGnsGDPd9cMMI7u5VMWN5xXh3fnph
Dy2LrxiMQhElRauMHin395gN1C+XIkJ0hOxPEahFrD3H3LCn8bcuRxdcoQV5YVFe
qKco7oFNuwF8oyjMNMUAJThd+pW5FugPKHpiVZkiijyAufmUoiPo0Q+4Nsjtq0Ux
fNOhtWthqalus0ci2y9y+PILOwacBqHw1tQIj/S/AphXqKMxC0XyTNf7fnfsWXZB
LKSW2/Za96pPF9Wc9GjZvm23Tf6z/RQ4XRFZKUUfAV2hh8G1ZewLtIAH6BnI+KfF
Am/1rrpEoCNxeuKtgiwMbsaJ+dnxNUo3mQ0vTUuoCQEVukOxKBzIuO+gw9u5AsB2
39ga+khNoZncbERFJXGImeNUorxgnEP6dkcmGIgRfTBJA6M0at3CNQkaPGe1ELbL
Juj7+riW1TaE2lRMU92HOFyIE5DYlu60IW/cgRg+jN131X6KaLnuvmRBXQWKT4xg
6rN2ZZr6DwOVTlgXg7+fm/Okye+bwlKC0r7/0ZmxFrpEZi/LAAAL9DLuXempbtjd
7BwpwC+9p270Kl8XLPbmkwjDcjieqBS7dGyjRR+R+S7Q9NSSCfWm4om+kfyWz32z
80+z+OjhbJpocju/zRt4O8P3rA0XEvA76COifCz33HIzBvKjaqPaz0sKjuvWrWb5
vJVGJdD2qWLO6JxpcUCLfT2ZHJtv1L4WRT2SJFjcDYRI83zguG93xBCTJJfiAjB2
QBVwVxNwTUdGbQoTQr+/vj5VkxxNTGfJUEdlXO7zw/7kNV1sC+qMEC6vwXcAHMZF
rwWLoxH2bqO4/sjXYBno0GMo4wi2tsw/1ugbDSEFXZ+gZgO5446MHfO+SNZi0XMv
LaNAY4/AflrtcaeQUDnO5KQ98rwi2fhIzqNakTU/qFFazoR4Ri1UedpAaNxSBfam
wfmYIkzHw9/7e/LdCM+NdnnVa+HlswfPrGv1BlvdGGgwiwDaArK81cQYiyjaIdxG
ikXE33qBzFG6vbQ/nsT1MphGFb7+/nmYbKFj1bNsJKa3sL+N4CaFQaWGmJS8SdcN
HMsQ0BNbMhtVBfkpEDXbUDhH4im6fAj5COhC16hj9Ea0ZrB5z79UXpJV7vBwzSL5
JAyW9TZgn6BdMSPLHdIzJC1uUDMgwsaiRqgMSg6doT3cY/cdg2AllourfHelklht
Jj1gjOL8gNoKJts5M8wjC5PrGmxh2v7tLhYM8qds9tlxuT/wTTxwW/LI8p/hB0nZ
ZvuXgwtEkD3aP1izkTJcEeCAlJyd0454oTgwHFybPJwW4SkgJ0OlhTQohwEi0Ylq
TfhigUARQFSkpXjgOSu+v65RHuQyvU0Qcm+DpF5oJZTrhGzTpPAjVUwtAKebLSJR
StXJsfnELMhZVZqEyoCjGXc1VFbDYIpiiTAc1NjRTqa3sAcZWELk7pf2dwsi/W3z
SjAD8VW4Uat11X9dS7WCXQp54fWqGft5OrGgYoYHxHUUPpEPCt8I3SEwdgANVEyS
HtAoA/Z7rf8egaLZn6QC4Zx1X5qLAlCfAfBfs1O/XNtUrqMzsWXWbp9AvtuM7xXb
JLMBFcyuNZKM8nRSKnrvHLSQ3RMHsqJkDhP/h8in/wde0Yo8WsBCgnwFjno+fHyg
wtm8+vEeNyKKxxMwfcIuh0+VJspzrZJ8xiwFLCIClc+4nvUECEZUkL+dKwFRwYz3
kS6TAOaMFgbqHosdB8jWcHsuGR7jdF4JsdFHxmb6aiqlIliPKtz6p6WGmrf6FtPg
uXbfBONXaRzbfpZ7EZOpcSlx3zrn4qOdMVctPtQAkRjyqgkzaWjV4Qdb1l2H/Xsj
i/knPM/T47BYszEoCiyAbrkfrks11lgOeG40M/E1hnghyWv1GsB/QRARyACde+sq
s9X2X1eb1bqomcBvrgkomFfNV0A3Ojy19RQ/fzew6DmfSZvnCL4UBIGZr592jxzJ
wETuLDSM1vug3UShNwQhGO1dRYZqHd9SItGl86NyyIcf83IdsGrvoNOCg43zb2+4
ibrzBLK44eVVv5sJV0uskuVqUvhdyl2Izut1TN4nj17YSLjljSUkDzIUGhiSyfRC
EjRCJkaYJ6AD1+kBdzRpjSOio9ivUtJjxwxJdfkIhoWGHDWMZJPzrzE5SHnaMRcU
E1LvhaHhRV26KDfgNwtWJuJOJV/dA0GFXFPsb4bKIBITnpE28pDxY9/1a2Z9OKmp
tidX7bUTLntsh0UIMBaLMKIn8b9raxpx38JL+yakbYddaJ7/X+fAHlprE8iGSayU
cLXUBaX6y2BILBrJ0gkiU6/NaIdUtNO5OT2m23Nbdlki5PxviUGyLhVCjGgNx9aA
a+svWlVVJCsBg17ZXF7c6/gG1AEu0xJVcGAozZk6bpY0YbiVq3wY1wpuZDJ3aYeM
q0qEpB4UlvHr7JgblJz29O8W1op/D45Bbkfnerp3BiEG0Q0C2ygxMMM+UCt8hwLE
CghaBZXIXRZYduk5b6lesV/wiQ+X+Wzv+oO6GDSiga8Xy+DDGeP/+l8Cg3AW+Yol
S/zTcmV0HKGbxYQ8lV53A708M9Pn77rdjo5o+ysHTdDUqdNvnNKxVIFpoStmZf0G
WcCV2flcK8rUk1hN371B98znnB5kaeizt6ViKcCQeNMvwpiIgzUjfWshOwp/FtGZ
0iO/35N0HGbzQCNkKW5vtOuLaspEAJKIogAKr8We/p5lGSvRjylJsa0a+aZrcAEL
xQHUXhKSShtrkMmDiQk/xgevid0XHxbX2/EVQz4CKSFZpIyNH0jF2R7FL6dYJIN2
k2J3RcwNNYzl7nNASiHvDuvRI+Bf+h3SJNOCaou6ZkYQd5zY826UvxSLZulYBzL8
0MwkPNcs2XxNjc15E3C9XTWuYYiqitxmk0BpXoxgN5lyzxftH2vYrUHIeqTSl8lz
SejCoOa1WtzSWX07IuFHiehmlKshzQXXAcVQMP6Nlvhof2rCJj43GyQ9P42XLTzJ
O7/AKo5NJBeG+XnxEAC78fnQm68RaDstshiI2X2ZQW00MyVRTlchbnH5mQiyRCc4
dSQ8vl1yqz9ZpLjgXFc/TbynjjTzznZ0nAf9BSVLX1M9KahblnQzV6pRlL8D19bo
dT1fhmP9veeGgkCju7UmLhjLfuUdJ1mW7TrLzkZzb4hME8a1mNo9zAo1xDoIrCAT
sPVOItNVHRoOkmp0cUMLaSUMKSShV6Ouw2hQwYsLeQhmLdhiWsLkrrj/8FyxJR0e
1UYIEwi6ESoIGMIkypMcmQOBtAzozJUv+Yusa6omujPuvqPbFPVD7XCbHYEZGQU9
0eyYAmtri8bFhGBiudjjJ5eSwc/2i2xwm6AfpwQxJW8zI8oGgTeFZJ6vl/Ce+tjg
wuTHQTWyfmdkN/ZvKxcxtnAG/N02yNVMtyYpiT3gCTlrTDvXvQ9gMhBWpBtdAkMC
eDdQw9pOEWLSPM45UHQw26DzhIUMA1GImIOJ2YJuaUkE8HZ1m9KlmpRPKUHaJShO
o4QQ5hYZD+S2Hmx7TwLtZxcSxbpcUDZRbF3f7tlTtMCMVVfGiwTkidHj6dFzvCR/
Z7xkk0NJWRI7LQKDvjaXKSuYuREWaGD8Jlj5wj28JUKgGxBZkJyKXMU/RyE3hNY0
lLbFEKbjsad9iFyBZPq+sTPbhak/RZrIWFxLnVy1JqOaD/Tz5K+E58nRJNbvQbwt
U3SxQ2HOCO7z7SGxM734r9DhpRdYPqa6KGCY0/uLS+J2kVh8fLEMa0EC+KCM86Bc
CJuk/Xg9BXm4D+eDfVQLmT+D5/ADMwvjCMXpraXVKF4fumZtEl6M3DgGZs4tiHGJ
GcdHCTmUoLc1mXLRXyfsnohXPKSFvAsf29EQmdiHPzSgjmNOm5r/LLNsnEnPZN4+
P6gBmY52N71/yufQ1tun5Je9cLREzrQa2MV0vZn8bV/Xl6oFMo8snTJ1FrCERJyO
WzByOokrVc0E8YT/e8ryMnFn0cFsx/XnWKWrhlDolIX+YFMFYzQ5/IEl7v76u1hk
JJTGPNtrd+s7yEV2iE23O+DUy3ivfnDCUTxNaCYXyb3TyQ70Mlckke1szs5+USeZ
qQROFw7Z7vbVV8ZQmzyI2920qQs6itN6slYqG54EqUdePOvnKoDaChH7sjKbngiq
oXsIOQov6Qvi85VSEqNcaQA/wW2p2/Oxrx4s49QMbeiHKMwjQr6WJDWT+0o/zdeM
tCVbZ6mLo/SunBBygjeYuAmfxhQJlMvoIP9NKbp6JRQ87I9/OScwtTV9LeH+6bjY
qhywHN87/2YOj9/SEVvGcLFHI/swr4+jaQl4RufB3NUx0Uv61vsgcg8kbzPYFg9t
kmYNYGEBa3j9/v2Q34XrRrMM2/1IeXrtN5HK0H+7tFBoem5mnok+l4ghwORWhJn5
jfa8KIAvoGS+RotQBvimgVn9QbvpaDB5AIlKBLx7NIqIm12GyUvk4swgO4t/ePu9
r6z4IPguIj7K81x20pgIPGdUEM6C3E3+NTtr7C5+zcECF8seSRwEU3JJC1yetUhw
QAUx5H7GAjbjMNlGOXOOAkJ2EBCbGU3KqHGJLhNLWYbhzKpIvA9Q+KCnnVQZ/7ca
HHvO9mnKBxTx+8lnwzvjPkez7LRoaF/ojKToiZyZSxMb17hKyzzqMWZCwDx51Mul
G7i7QlluU2cLs/M5AWSN4QcnqBcddIQS2VizveG+hE+ebsgnUxJsUfhIWwSckI8P
I/4qWurVY8SZoY8ocXbTx+J4/P/diIHMcYTsLkEFFEtZbXNtTS58kXHhHmigWqih
FJOnOhxPYqP+0kGLSxUVKlO8vzRaUCJQCbkw0QKbIU/VyiRpBRQr4GahHaE8LH2X
7rYYOO6Fg+4xDvkkJcOCi6/rL1EjCp7v6HWbJcLQDC2Zh6fSxAioaMMolLPTkGJO
5Mxx+CaI71dmoRv5DEWaAuxU3XEeDn+bR51x1azeFlCKskT52J/42Ppg7VfWvBe+
QdJFrEj3e2V8C9BHqxnRSPJCP/CLKJEUbvsEwkaqj82rldMv6crQUWkb2FpSedXF
N3UxARbJsIhJLksVhxL1nDsfUjUil5VGehbVg4uqK1+x8cUzpAyLpalqOX1oh6JE
9jeCulft8D6nEDTBIYlCrGJWg34t6ia+Pki5OEGI9p8bQmY6gPPY79QlhCppvdq8
XUGDO6ZIqP4ILXcuuNYPiV9vE1c2ROyEAei+cGurfMpYN/PHaFbTVzIJyPtFX7cU
yFu1QGkuRD1ryXkgEa51QUYObgN+heR2LVLM7PXL/ZldM219iM6Msi5mmZYyatQg
NGxxVzj6nWZ9TcgQ3nhlDiqS3DIhzRc7FVs9XLjpCMkBxvljjvMnAmZpvCwacIDB
xJtHa+29HMkHJoH+Fwt/vBI/+wusl9FH9UwTX565oYsCacIhkueT7Bebm+FosA85
f/Yf6Y7sdqLASIwZ7XSsrCZxDecGXRqTxWKDRstG2t6TaDUByxN/a5iqyPIBHF3k
GTItw3f/kv7nE9CHG8uAtbPm/Ui675LC8pQEDXxBDkMKoepVCeH/CIf49PpECpZM
hkG5NuBX6ItRu9s1JYhpj1QRnYzAT6IAqyKy2eNZuDKy6rywauXLkeNm6/QLw7PE
yoZRLIhreMOFP/hK2SwVKRTxKpSma6nlaZrJO8CC/He2hDrblGxivjSuei15V5e7
djjWBTcCkzJum5CJvdcLFcY2wzC4aY9webX0nJTMr5G5mHB+XKWvIj9GKjMcIj7F
BambdFI6zYL0iQesTLLF2IIj0+bsLKwrBVWdPn/a4DYihBI8ZAT57okgqQnlAQA3
wDN5m2KfiCj310YIftKDMiGfzhsnnybf0fK4UolyM9AJhHVDQGTK35lsyeTwBXaL
0WJWgwUhCCyN76ryfWYuQnVAep4fbgAOd6ENpVXYASk9j0c6ovPRCCubY/V2XND3
zRBAEc7DX0VXwwdJ/cGvvAdbTzniMTq9wtR6SFFPuDFuKf99YUFQJ7S3a6hQ4BzV
/36vZvlCvt0ZgVRUsCTna+GxYUNSrwXgCNH2ynGhJX1L+7reS9GKfsgtQmI/TWam
/7ZwGSaClqksryQuDN6P+/Fh420tx2jVogPgY5iORI1PsO6Xpbeu9W3jUvaq3QvQ
CvcIG7eXZunV8NLuwckKe1JhyTjRLkAySjUCIHtU1CRR53Cvdui8NkLshJe40UZr
1EN8POwa3qeZ1FFGawwRSg+eblDO1c8VsqBkPaNUQy8N6paYDq1gDG8I28cY1Yeg
lGKhxDT5q8HraVqjsDbDrN8jJaak+fB1Z9EXgtDNs6hI8qp8tfEgtbQhOZRaPtni
OahESheqYYIs9JhX8dOUU1BcVNRRg6rTi06XfwXW+g26pGqVNjm2g7ZeRmQUHYSn
Ch4BMQrF27djzlStRuviUNh2dHlyld/bwBouSvLgHdj6ht5QBRo7qIfazz6dtxS8
weDwDD9On2Y0Rm5xKeyimuRAdbYLN58IGIBo/8HdIe7TkF3Cn1jugNbyHuWI4hj4
siICUGrZe9irmMP/uI4XnqJVz84DCAcZJ4sDPiwrQti020v7XOHM5yxvmMFvERzO
C6UNN6OoRqlrf6MYhYD45H0vNfUHnaFkwfwLzw/EvS2AzqihC/KC5DbRlLBhRElO
m5XVtI9Kq510/Q7wiqXP7FF21OW3mKL2hmJRzkjsmzf+9Wj7KEGpIQEQFtARDd+Q
/eB80XyyVcj4RtvgZklBLyM8me+vGLJ+0gLRiMJ/+97kcWAIagA6YAA32CunsSPI
qGQp9z85skM31HJKPjFIwHVrF1Hk6PotK61mvEYR97SqZOshxTBiAMIBe9kwhyi4
mc4PQ3hJqX5PNYROgGZPU3aERBhCWOpmZK+jwzx/vO+xxP5299JzJQS1rUjQCM1e
+Op/FXiVpBdfv7g2LuTOrzb8jg9nTJm6eqV4p5bmA1skGRdm8OZNNpIMbpjM7n/0
955DUBwt7mo8tx9gWgVcR3CGoor1/wkZG2D/XnVNnzq37QiAJZ6WkR+glD0aH2VU
2XDhuFCN1MJ827TGkOiSaWgsgExK4ur121cDObazCj1JLtxA/PW8v2EMO8TwJTfR
Fz8Nv43fAOLAIpf0Wo/WyD5R0tEvd4z5fgy3eslXra02Bct9b4oPOvD/i6b94+26
MIJ6YpvhEnA43pamwWVO5wQWTqFUhWShdNu8qsXygyMp3EtrSg5xXINzbiNpuRr1
qN9GMJtqiOrIe/YQoU3pKVemGewhViwgGc+IskUvdYQ9mw3QMrgvpQr01JcCvFBZ
sOlO+qP3xT1MuArSf9Z+J2/9G3i/mUENBQ48VJE/vbKts2SIX0OVJYXctvkxpduZ
GEOTurHOh6SGhb7IPvXRMF4Qp8vmJbnTDwYRbcSyIeHcbb61+p7zw46eVX3RHwB1
6qogeKkVO25Pl2DQJY9WA5ix5J7MMTd1LIPXX2/M+DhYopYG3e8vZ+jaUuZGKxuU
UATugzHLOVgORX0JQpueu09/l0hm6Y1q5IDaytTCzUI2eEIeE9Mgh9d+nevqatYB
zFfcO/11QrOT8Lh22rXF/EH5D8JJuMiKiRAT3AT+iH2i8FxmBaLhBDscaeaJuwoP
eBt5IVSV3Wx/xBtV7NFnGE7Es49QBKO3N2/qq8Poge5McNOKbhkwEOuQsdvKC91b
BXMpoHoAeBtZm3mM1wXeFvu6/UtoVXRYKvlUjqTG5U4thLSV2Om6RcJGUfgvldbS
WIv/OL9XbBQqjJxkfrZ1bHQ0MOLN4yyZuvtlQuPpBlfxkh0Nog5Wa2oy3Q0x0H1x
iuHg30KfvUFneNEjiL48a7s9/gHNSXZVK9X0Qc7nBCHwoB7UCcFaQ+r0MwOgkBs5
`protect END_PROTECTED
