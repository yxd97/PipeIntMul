`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iqXVl940NvEI1Sc6IU0lKMVm4rOAX9jf83sipQHtS1QD6oWwdi1aQA0w+q9HBUMV
XjivU+zbtPN6/F/XG4DD3P9YrwHKmGSkhOiz2Vmi98jDnojSR4+769SuJ95IUoqS
FATSuq75hYXb5Nu+FVKuFqQusHqV/1ZMudMV98vDLzghF5O/7fjL5C+oQAj19zWZ
5xpecyz5/qFy+d8SL7MaP59Y7eUUJyUJ9IBlhGlsXPNGG9jo/1/duy9YULj33qq9
cH3MVOM2Yk4UpDMnf17TpzAd0kRvQpO3nKR/HLX2oKUHDIf0eDSytmFaQEIcDKXx
mQ12r+kP+5W/YhWZdnfyGszzYxrpyCa7dDYGhXcpt5QC5RcHlEF7zhD+6uXZ8yck
R9rsGYcSogqxqaBJSwpZ8/BZmNihb0QWs5wsCAx/AcY6YwcF1k4YppdBeAs+EO93
yAuV0RePZSVFvn/GlbhGBg==
`protect END_PROTECTED
