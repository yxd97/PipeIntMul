`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DLTFPRIGCphyBCOiYqyM+LXPj3a+xuz4TpNClWFmGwMM1pg30raiDmf99G4EuoXZ
Lnnr6iOMkuDS2Dh5yfLwd0NhsJcaFJ8RZbZU+ktv1pisxgaEDktTv2mIS+bvFSRb
y5EPN2euX7+jv/0Hrh2jKMgB+KE28XDuRJfwOVCHHDmPXcR9Ada7PU4zH5jaSJqR
bfkBcfh7powPyYQlvpzqyBIBAgPW2MOAGyyOqNJpyb9CvA59hUSabPr3usKnvOD7
jhZo6ZDhw3Z6VreTletJSUqkNBSS59emIpSI33BZhAHunS4ZrpWqN4MoqlXKj9Df
J/mD2JV/hzYQpQ965Pvs+XGn3JfzlFYLcvWrbJyQcVi8viKxFr6BRXuYrJx+4Pip
3i3p1S1z+vs0vXPL8ehxlDcGwpuqYPhliDQVDnOfPH4uCGsyZOfK0SDQcpczd5cM
rfNP0Pn1IcpjSm6qhbaDnzdBP34mu2Uzaype8SytiLWUseOoSfcE3QqBVfytYDKq
yWCWZOME8EUS9/FRXv4TdEl1IWmKiQB1IwpCke0m3ANvdVo6YG6Ou5WzEJHNdxsd
9pziePVVDhAwNOOdx4XZfvlbij3/gfYEcuP5seNldgRUAhc2t4q8EjSgOEhCT1YC
HWFA1JYAktk7E37LZwLr5s7rhwLCle35nyhiKVgNZSVVjNgxxjeQFQRQlW5c3Gis
q/7IXd5HhIT5BDj30Pe3KHFTPjk12KPJdJipsZVQHEMCksXCphWDhoJb2ijR+pyK
Z8bsFy4skOFgoKmf6rXp1XR2BzAVHR2vDpSA34Z+tGL6Rr81AiRsYtaR3f41TUYR
AQ1OuyP0gXiHK+jPZfkPllwdhh37izxcTcNf0sNSCAjaafGbCrmNz6a25DnaOfoA
r6XpPIP10091tV8MSXpXHV1x7uD2y1Tu30eD3Xi0zvQFjDsjt9rZI5sdxrb7gQcH
Tn7l02Z26T8p89ffvBK+48OtkERR+o3k/Y0kNvnXCW0Tv7d65HGm3bjYfQUg8oTZ
ElID9i14c/BlmjZsg8P55zxzvlnWdciUJdyaOB5hPatItEEfXrefbBgkgNT3hvmo
Wv9/vcDfHakX/MDzibph2DtXsfiIUCU4VatfCJGMd3LnojXlzRUiutgHl3NrbqjE
8z1/tVREevM7Bo3DCUeH9ftBozmqEIOg5H0rrA6LMh7GYVIP+lJjCcrYMaV7frfM
fOChd596F9ZnMTx4a9ACk8/BgHfDC0aN6Kb3uEv/0FQoluCr6fFOXXVf5iYNJ04/
ks0THgUbo7u+tKgOHHX1dfu01I/BRPggMULVcqWK/3VH9gj6R2Tkmzo63O4+V7yE
4e05zUMacYvu10KpfOx3wGpV7WWFJNjneDxn3u54lNRpf1GvuOOrQNfieuMhukIE
cJEqfu55yAj8xhzuoTxHD2jRWJxAHbPlYBiYxfVhyEZdqoalcLq+5g7CzSbJyG3y
vKmT2gD+egxxxVyW4Qk/c7phbFWrmxTf0WYH83t8nYFYMbckF1DPizUAajdzifJm
Yvjw2wfiRFJmFuJZwpgWd7gwKgu1aVlIDzriP8C0utQNpp0D6c+Vg2XX5CrnT/fo
fMm2YQ6NbKDJ4O22/iVsojKHL4BSmGm5M09kW5gCJmcuhcYoAeaZUmp/h6469q8I
pZ39JUfvdbjHAt+y2Rv6Cna/fEm1cNXvAkojukaKzxVnhaD+4OwGX1kLbW0NMLZM
77YXdWK+TUBhQPiW6x2BEoKSk6YXKDf/HNGorAVCXGf7iGO/B9uLLumZAG7f1D5c
26QavPcYQYAi4IyDUZkCqj8YIwjFnRTz5de7nnQFadTgnPUfhdLH/Z15kMiQojin
mgJPGLlmxJNdjtnFex2BLBMKVbqL3+xbFDUsBNINXj2Y0me4B7yf0jDQZCXmBKEq
hAmo3SS0GTXjDUJ30/SkOtQmjWGbTxB/ha0t5dPQSCCm/K2DiVAxRDxFgJ1LYSf9
hdcaOk3wOoZaltlWHqkhyfiipbtGN8og+CXhIBmVWevn4t1SuXKOJ9YD48bjwjMd
aQKR2HqNgl7Q1t//dZulcxo2FMQcEnVcVSpg4HoB61TedcKqfaPK5XaouZepBwKF
PvFj4Sxt/D34RjiyhIbuwN/vuVjgPA4xFD2rUc9u7IN8WIRicu1XuDf7PCF/jdGi
hAxuDeTcX7eByvxotEU+3USeCqIQS+CWDUAlpySgjMPyRyzu2i5KyA1N181QdAp3
yggiqF7Z95HdKhhacEqh8WwrIQlrcsvQCHGFWNJOF19f4HpEhl9YhrTUwzRk6UJB
j1zR1gftr+j+aVTDgdfb0oyd/PD2GyoM5KFhVjECstZTo7dDTYi3m0xTIeRwVa+K
uf2hLYY4JCAw9li+df1q3ib70UZHIaztWSzBFSoRHehng71Lqy1oZaI75JGQc4FQ
O6zIVsmF+86TCaMD6Ib3DPuzaEZUavdEcpRmu3JWxrTaTKmwMBI54n1TYFWDoQtH
`protect END_PROTECTED
