`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
44qVUBEakn1aokElpedWmQFo0dQ3hxYJk79O1NuaqMr09mjDI5ZlDKaFjSeeeDlB
tabsDnVk1r9bpp+MQuftfyCS32GHfU9+Yn9zT3nnQ5EVDypvPJSsK37Xygfvz4w0
xVPKDw+wEGOejlSk/rt23UgcNRrGFUSN0FFn3oJ9X74ZlnmF1W0ltquHtPsuhpYX
LMti3HT+FPIPihexDXCaHw2MbvdzOTJlZrzS0s5KHEFbllZNb9oy6hp7CblWuGgY
WcpALJL8C3IR/n0G9tAAT3himDx5zPVHzbn5XR76juIB0KfNDN5HQHDVLXjKleEI
MNiBPo0HQNSvmxgy361dq6SzTtwnG5wB1maUsFvLqS4yq+7LG2wBj+1sk44P+V3p
So8o8CX30FjhESl+5P12UiDolzlm1XGveK27nm088qD76gGI7MkFpO3yjzliQjJC
PiGvYbSR8au/h+KRVwo1DfzDaP5OmpaNGY+cyPn+aNvexFpF+NHiT2sCktHAto+9
UxmDDt34rWCCZo2j99CYDZb5b86I3D0E16aWd791KgrcNVt4vkLi/e/EyqiYotg6
E4LZ+xPy/lzMnzxxEqdEn/PBo3U8Q1RQjAzMCqb1YyMkU7+PJKh9RfLYYcu+XZbH
Kjgdvb3uuVzVsPn/fAFMHk+2ctyLDzoCl7qWwiVDSW6Q0eB9A7tymp2p9Pp6wMp1
l3U2jpp/Pa283fy8H3qmC8YH0LVj4+edshchw1TOvY/9XOCk+JuSwRtRqUj+ERAV
`protect END_PROTECTED
