`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rvxy6/HTMlMboBqi9BUfFBJ5mML029NxxA7wn1mwUXV/CDFLbdrlR7qciHMcjabf
UYci3tZXZE3KtkSpRnXv24OuHXjGAGa40cNTDJ2osfC82Miv7GJeHUAvTqOL2Qf1
2PJw7cX6DUibJ9MrssXuksGspogzNUpRf5YKQTRMAaYBGgfycRS9ZXSQ839HgWex
e2/4Itmwos6Zz5NLDcu0ZbLE3JxwlFF5nsZcrRQiPc9Anq4Molbqqd7Iau1QYm5k
bCfPzsSBHHafCAarARtr9oLtj9/o3qRqOUEYcueuhl7yBaVXTHFo2r1qWKZDgGIZ
md1B+YQorE9ZXlVicpBepGLTb8RcPM1/xNbpWSmyZBpyDi0soj+OwcAB5L8maLI7
TEv4CaxDFo1EqEAczUlabWDLyIN/jkbXrWcBiCqp1cXTdakNaZOdX59VUV0Zbhp8
ZpGGMp5X6l5PErq8znc+r12FQATz05BGf3UetGEms2oGrKmOdie6VEddL6/KmPfJ
U7hgh+jrQ51uOtfFXqTYz7ya/lYDPocPzLishvGhtybPcuBx5BAT2/88rzMK/Dfb
ILa4i6tyIZZVjYngKsYvQKyDkjFvKc9okd1tTxo1NQtntDwGuDdc+/TzSFgdsfuz
dVleFjxv7FvBCUdCeJ4He3NELCB4RGyVWx1R3G/Fe+njGJIjwwEESVJoQtbF50Y5
WkF4EHr3ipf+YXG8zWXq/7lnIBaU8PmLveRhVcetUyw0uMMs6SUMCuo9NWRR/kyP
A9ukitm09QqUH0MtW33TRZVBX6C7lPuclEQRJYZZNt/f8mFzid5u9jm6Ne/UpKy3
F8SPpteKPI0+iP1lLRhJTjO0Ef3paNSKGUpQ5oAOOFuTt/+VWK2vXTyfIaasna5U
ZVfrVPqK9W4wrl4E2Mx3SorTrmLYr6ygx754iBaqtnwp0cRcitAM45H1ud2OR+M8
3XmJgFxEB0wlm77F9bKxauEwWUE48sWbPj+SNilGy4cnJqXawE6w6bgx0G3a3ZFE
jC8tghJ8B7U4ZTUIy8f+nFLdS3y2llOgly4O5tvRWYkw2sNdqeJRPv+t7yekH+P1
TXnePXXVn1/rKelpkWTxlO0N6ZdfqXRPjpObbiYy0PKNgxGuHMO61ivP++e5Bhdy
0tT+dwdLooZ/lX8YB40TreSaEbmc0UUP/EEBr2PLff18p22LXuf8Jc6LdGVfdtsG
`protect END_PROTECTED
