`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/FmlKw2KNAkdWeyCjXB3Q2gtIvrrXF/7jqIZyhuBval4aADiwDW7cqhbDOxPrbjq
ii0XpspowLi00lBBGFNAd5DeKhYXnPGqG4w59RwQHHT5Houvtpw7k9a5HWBNGHwV
HI/HAb0MapVBU0ZY2SkzBxFWvvkmhC7neSmDCywuNAU3cf6fYEeiR8yuKvzhVSMD
2BVbIxVtMQADqY3duRah4YSs4OfY5kXMs9K6o1tECRH14nAa8J51gNJ4dE6MNBPt
sf4eJ4VUThSQ036t0ci8qHri7XcbbHU3PQCA6x46dfByXxQvUgXdaidYqxWHFQIo
D6XG+cee1WrveF2G9MOVj9jETAXE9NufP3a4FsjO5ESJ0bLUn+2mKG2TasRWg370
I9t6HzbLXD1sYpDHixILGQ==
`protect END_PROTECTED
