`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/w7RwdLx2PxH5D4+95u6Gka8HROBDoVxgOw0zmgAUvqq5/fPXwGekHeVrzdwu31W
92wSKRpKfuwJGBtGVoXwxoVc7jPR13fWTlYkrPiXc9AG/3AEYwsDqWsfr5Ro5Jvg
rPA2QWnWytWxrY1+DzLGk4EVlsGpxH7TbPypCGanxqFBZDKZ5PzNLjVOoKYzbZ9C
hC3YtXlCqNqGt4m6DrlxgvH9vJKUak7+6JywadPbEaxVZwV8hSN2TkP8WGB15WCK
C2+/s9o3jttIQb0Cl0Sc59WEoi4msGC5/PX2gh7kp96c9km1StT/b4uN0PtfWgWA
VW1Nht1l77MnHxFM02BwlXm3Zhb0ev5upCcz4p4/7EztL8BQ0jB+c9XL7/uFBc9N
FMQCxjT1jEY75Sh0OTyiVB1leId3A8eVeGgb+7mQM9MfS4fI3NjSK+UsRht6DK6P
VEvJgAArdNU8vHupnQqWn5lPlnrdhysqLkQB4v9UKRQ=
`protect END_PROTECTED
