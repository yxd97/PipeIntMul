`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbpRQCnZz/q6t4/t8f+piONVGVSe4MVt3CNDAWEdZtio+cTGQOTVmJZkXsj1Jmrs
5iMzGZi5+ffwpc2q/fzpdVTTHxtnucNd8Cr0Sq5WlCMTt3KPXvdRwbw7NsglHS0d
pbF0csrblIGAgjGBdM9M9KkWfEheJSSF+2V49+JuAazEEBGGYqIAfSBqe7Mc8XFB
BCjTk45MIURXQ3NN009+C05qE2RjWxL8r4+ZtC9lVxnlahZs+uwHGWXBXeiw4Fgy
MKp+YK//EKj6hvHMNgK7KfEi3qYCLBvNm65sARRzUhJTS0v9ocft0oPYm4KmX3Mc
Z8jLVFeu+1pBlgCdvsFTkpngh9efNwv3/Kh2ZpF3e8Tu3aAU+xACITC7b+0CpBJ5
zAS5U0JpxSULjxHqp5I03svXoE2Ob/bEIMFjB5e0KwUH5uQTTXpwLZ3iowFkcJ2b
`protect END_PROTECTED
