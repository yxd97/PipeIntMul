`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWvXFCqU3E5v9PjGgDnYYJ94bMo3nZB9437rgvAaxllgixaZ7giG/FeuFOaJq3sU
U2cXG7xbSwxE3cG+QInGoZy0zW9649NhngTnHeaAMhN2vHf5url2J0d1IqrN9/7m
kLrd8Q2987j8vqVYDgT2imKqtyVsWu0TsGHOqW2Ct9H7AxKY2B64u9VV9uNIRJpQ
fRJ9QpEM3AztGo8rDrO6+FGegz7K/Scz5ErxAUCLDhRfXuKjxYNwn4SKDK98jHoy
S5BnDmxSuq2I3LR7XK8IB8SLePeScB7ODE3JF9vT/eTcAMpxkzWKAevMyKCfMqMf
I7m5pDcvAbh1z1PQzU0NWOCPPJvmn2VkhxZGd+00b/6qO3vSD85xFIGTr/hkeHRc
DpasgdiC/SBvdD1ON/EHfw2ZaaTjYrrLjwi+gLeoEFipO8HL6Xf6f47/gM87qivL
i/fjtfKYY7RlKNXEf6TG6TGgGcklBpM8B1962+rnCvxEJ2zpfsc3XJ2/fRoB9VMk
6ybNwtec/G09M0kHfaw0jgvoJafYPH4IUaojbVCb42WF/ned+W3MYZwfQG7Ho6gi
Zo/AtqA6b5iMiHNlj02yH3vn/wYvf/rkWdbptU/fABlcUuGWx/HTUbZ2xrpGPBCo
4JAD1mrEPAfqBSwQRdS/2D74MHzXLrwcwetZKjQsxm6ej88szr3gbCMaDHakEky9
cguFbzIqz4xvK12aMZqi+gNqmqHUCAP1UCFX/9CZeg4hRIfzmj3maZ0t0MOJlE7C
29bmDSKhbFOV1+xufle8TMVz8OYT0VbaIhu8qyOlXSYiA/qD+nl9kOIbfYzGf4aF
RnRDkeWLppvzy0BK2Bd9f4/Z7sKu7PUhPB7BuYk/6I3JhJNFrsvf+6nvyxHX9agT
3sOY80v98fpUFBOECqeSCmRZpz1lVtT05YCusrA/2re1nSGAsTelassFhKq2Va67
o5/sUjjEkUP7Xt0NvZ5YHvMZQO/hwFFXpQFVXfPiIGNMhHsdhM/sZ0TFAn6gSTLJ
wp0HqHUpuD+U2nrj7QtSS9ojCxhoouPHdANDjAhxofk=
`protect END_PROTECTED
