`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59XyOZqwoZjoWfJGiKGUYZsFVAPU9oCu89xzfLfifgdXnSwN0EV0e3IOJjno1YyO
kxUP5rmv1Oc4M9WwU33eMDzImT4wa9pWVof+q9l/afGGtyynJjVllnGqbbpQTosu
IhVAFZILwoVxKsG4m+8KcCKnHQLnvn7mvvqD1rJdMyXFu8aj2gunai8GUh90lizD
sDVmKTjyJIFrVd/30CDQnGoujlSQtIwb9Q41dGMnQxAgmRuo0p4rsgilE1s5/n8b
aXnbAblErK5vSHajmhI0g8cKFH6cGSvEsTAVoaNdIzEl7QYllrysH9YXo/+CrH7b
dawadZ3wQodNvM8fZZ0H5WAEI7IJFrQ1cTHBCg7qMofOzxwISTiYl9bA63IdbEXc
wXQxayPzNY6rR8MrlLfu5krLZTaAJFCqUzORjIqoYk869wCRE7yFm3SXUCyiWLMO
63uZOltHy0LhMGEHcx1/gGEUNbvIURo6DbMQKJnaOEsV5Bd08iFDdYEkNIdoYZTQ
Fl33IhW23KGbNzGYbnTzkgVGxOnO6D04G63Roam8RiJ0F1TFo4QUiG3P267Uq1rK
aljpbWpJ6KKRG6sOWUqKruAHMGn4/m+zfeq03uxEWCagD9qlN9Osnghn30wSKzEM
yi/d9xUTQb9QqjIsgw6qWMiSW3+xwKMPwCjb9Pa3L4Y/wncj/BdGFvc7DwRbaUxp
byNSEQfo2C0mtV3hSN+JcFddP+iVH3tDmK+C0N9V4XT1xg50/tPkASz2aJ6Jk8sW
GHoIzr+/JQhbSy7tjGIHFAVThF5qGY1VjXHIICKhUEao0eN0mIb7ZdKGXzPPuwPm
6iE3mzkMcHj4HHGTTtRrC7ifrsMhdql4lP2Sd38mfCdGuqbGBecREblTJ9B1DQhO
tvHmR0KHeBVv0o8rfkOOQbY4DkrTYms+sBwo57/pErNzLQ9wl1AC0VrtxTY1IHCo
hvjObBcizGDN70ZuSRPNye9zROYceDYZLgYYpH/3B6DNZkOG4GZ89YiKEEi1sDQt
kfCT8vc/Y7xKmEXhgE4rhg==
`protect END_PROTECTED
