`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVkJgFZ3p+oXhqXuwK4nn9fkZPJL4NqLPJ4OSmsVBKhaMCeGn5WEFkq5s4XfEeSW
iMNWV2+bQnaWE72Dec3DjPoFxgreGXQnVARg46vBqPD43O2ww3RF43k6cnYcKOly
V6WRZuh+7YZZTWCaj934Hvyj8WMMTsfnvNLjdPRlcezcwAi0PR9m117+WNtV5u22
bDs1QL0HOu4aG5qnc+pRnZ22RBvjm/hl7T4joxjF3Frne4L9SLiecUm170zfXZgS
FkyrM+0gxuFUl3XgPfJ+zuRTlW/eUyKjIuE4/3eiTmj81xJeKn0wCg7DaGk14Npi
W+nVgqgKyh7COS78Pi+4WhNXNmftfX1BF9DsooOHLONecCmdqNz8SHDd2gpUkMSE
9TPW7VbXiX1kYYdU4RvJdQ==
`protect END_PROTECTED
