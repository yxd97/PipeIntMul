`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nrxzg0Od11t4yfOKW53b7e4IIFsx4dcEJ9BzZfsT1lDoiOeoAJsneKKDvGE1Va/R
UHjj3aMcj0/Uf8kfPfbapHwip6h6TEBvtFIxfaMldiwL2q1v/eWakrGZxeJCqsR9
1K3u6gId747ZXfUovtsd4+ISe7rC7nzmLgJWY30uAYEEsRkGAm0k9RDsNWeDEtTe
MmywNY6VafWbrRtCaSYmHOnCz1a+4rSYgWes+RcGo/sL0NYamJz6wby+Y2G5wWc2
VkZRC4IPpubf1btEHKsMaupVTk8HzX2KtYCjtKssJmLpnC47IxzVtuIK/JDElNPP
WYfiOa+aFkCDzZeoJqZjcx5woRGdTugjHQEKIw0n44ZqjAL1x1A3uGMotdfpOEJ/
k218tcyMmwF/oqBixU5N1A==
`protect END_PROTECTED
