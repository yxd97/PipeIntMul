`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r06/aoFhqsOe3W+G8JVEFGik8ZZpo656rjN38dwFgeDaXyj7LAiv1Pl7adgGxXtJ
nDuK6K9ET66V+JO5b67WkjW5asBQCR1hxAGguMeBaXCwUuyTzKhHoZk0ktmpWnBr
7cOXUhKrP+Ft/de1YXcy6sCooXtu4l5prFk2MM4jEAzHdW8Y6+Cepw/V2CxN+tI1
S1EXOLLvbksq3KSkSD24kMslu2dITDbBiLSSKfZWWQWwCVv/yu/qCNfqDTiDSkQh
poeWVRdT89UkDVP/h4p0FU8am4CtqfnWw38SNbuNQDRauLtQ+uDe2Pb5TyYToGNE
ZenGEY9Ex9CSS97UpqjHZBwbY2wOk58NC1Lcht9CQWyjidweIUpM0dNhIkMAcG6k
h4worGfOdMssot2WFMXnbjuUVisIDy14TNzFX4UmqNh6J4jgkqkcKAgFho2gy+w8
u75Z+i0b9sanZp4Lo3CcdTmUNSIbqwi9dJ8YzNV3rv6LEuH0F8xzCDekwtluQc5K
3Pv+ssiDKFg7xQtEeLumtzZh2CytyZY9tW0qflmnqXg55cj9mjWGWz8v0Y3I/TkH
hWn0xZgrmr2dOo6TdxOU/5vvHTjZP2UQX5vmOMGIM2+Ky6LpCEyCThUgm21SSjzf
RS7J9rQ7GBJVg78EImAhEQ==
`protect END_PROTECTED
