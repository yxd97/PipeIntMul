`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wcvjp/2+cuoGhdu2xYRGs7wwAp6BSYisXdf3icALKWxdLLDTkMR04hAtK9NO3vtF
jjRE8Ei48yHAF7VlECXMVKMGc2k0hqKy1qQd1iSMF4gelcqBlFsCp0HpTr1itwBT
i8ddoKR6BD843iOnVKfGLa7x/Yn97qiJ4MgW304U0Mv8gRq/1wmhuBf7qmuscIix
5QS+5BN9RuUrnl0tt2cjDBMWUFlXnN+QW++00G1QGO2wdA4MxJu5JyfcExpjKYeu
qXZQXBdszASo6AHhvAgVvzAOBP3wHfcgfjIPhPqIRMG8D9yYsHBLCGBsPISoDYH4
sNH9DWKcA2R69XncqAdyABTEgDWHonFaSImmSE4TXzIa2mTXfCGcvtGUtTEvc/m5
TGzX8sC1NkaUWTlLLff66EdMcy3UfCAIT9uM9/hpMXYYX61GW7apwzjOc5QA5ABj
8VvzztIJIwr0kWNxAZEtQGdL8ZAbeCbZ2zREXXpPkwOS89dX5f59G+S1ziGNoH8x
`protect END_PROTECTED
