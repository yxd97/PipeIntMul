`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lvhmKGz4uUKlzoleydVHBGtCWneDF88oqhRnC42zDUlWRJya7e8D6f66bojsUtTz
08sE7x+CQpsN7svBEG+xZoUosQFZUeB6U9wOnoCTd35OClw/xq8QDUPCftzBx21y
TidmO9apSms7gfHDnx6hk83US4TJWdePcJcnSTOYwgZ29zmSeKBWQvhazXtgzrIA
9MxHNHvn+R9uu8FGj4w2ULbvKemffFGX20MS4/ZlQCGvy51juXuxXld5Xk124RN0
A1ndjGI5fP9TpwMCfw8jzx+wqj7ELyxU/8LdUmxT/+i1XrCpatWyU34wjePoydKD
MqQo+o0JmZZk5Q/Gb/htkrDADoo2dTTFUTjH+eHREbyiykCR4iGH/JprIFG0p5po
iCIFLxJjPyhEaD8YkwI3gFCWSsAsHVYBNAg2zHlZ9+g=
`protect END_PROTECTED
