`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rkk+upzGUFw70+oWpP7wL61084pAk3qnejeeNRQRkBGk3EZoVE/IhrDLDMIB8sPv
Db/phWYVgkgq/jTdrW0N5ycWInPwOAwm+ZcquPlFzxHfJz3eW13JIRXEtHuQf1wx
HWkDhRJvUfF9sdMdrxcUnbyMriwJxRnr0/BI62RxNdimzhoTpAP7zxoR31SD271T
Z6zThS5L0Evdmwf8G2CUrar7ckUgryg/a4YDb3/64Ukz9ai06v1yQkYYJjJJnYZB
GLEI3bv00Yi7b1/YG/5ll7LJ1y1h7pufU6f6zoSxg1tjk+OoQz1Ae8Phw3V+sOM3
/RmWV1zrO+7TUF+JkxMjQYN/XMppWjb+WwtD9YyDQJe//JA6ZzfM9Ij3DregcZmT
rt14KCp/Wl0J/whPcUj0rxzhGoYHXRhLeS1Qlw1dgvKcwpcsPiZhuvCN0gURjFrx
h24L/iTQdK6TI2Zlv3f7rh6GRQgtz2k+B0DchmKHJ5AUfWzYOlf7WoBQjnTzWfR8
0qgiGu3Z03jcKvu2SAz8pHvDxhKeFdC9RK1IFRFdkxaRGo8JVTV//TT1T2BSYcaO
RMLI3obEvo7iJ7WnIrLO/w==
`protect END_PROTECTED
