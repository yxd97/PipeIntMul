`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGo6uS3D7CNTqjGg2pOiG33XBbYjQLaV7pO2nXLGQ0ZSTHohsqBlgI9viFJS1nY1
FiLV1i/+Vgy7AUDXJf/z6VN4b6teC7azSDMOjoVOOVLUaVLre4rQVN7hv60VXaqw
qfgHE5QJLpqjWEvJ45mnDBOuWQbJomzI6s0IoSSLK3OK6zHzu1G/H7hxMa6p9Z7e
EFl3+78YnvvLC2+7hpALw8vkwZml9LaId5vH+yDjIpuAclDy1iYT16BlKorzrJrt
RvQwi/W4/hXcjr0O+K6DXs5gE06kju65gUDUwA7yvXxTJeCRwPEPXKcLPaxPyDTn
MiDgwJ4D8DSwpCVx87PvZ2v/wza6ZwDMfV2tIZBZJZ4CUSCt6gU9gC6bAD85+6xj
O6Po32NJiC86EYcYK2SJV8cJtpGhiI+WAl7CN04hiAU=
`protect END_PROTECTED
