`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eErUNIaZ+CMwl097RW7YpqCIHXBkSoW5qRj9sJ5cI7mUOJt74N1J9Df5fiOxdR/m
1PHt9Apd12rdOgvkASdYcoOGWldqtrtpzJPeQiOrHhpKLDzZyv4zdSZm2Sc8E4aY
uF4daUPlOruN/HznqLcC0G/ls1rvFUd1ScOCfg0iB3XNQREM0hz/vTfQyNdAQJhG
rD8pLlL5gcJtqPPmaBIqu8JpvsxaGShvi4xt5GmGij9RePxX4M7InRtqzrb8zZuu
N3bB1xVdVD6N13bw+RI6IcRcEVZV89rjDa0V4eU1wPSqR7pPU/6QnqCUzfeCWuL8
wDNUYOLUGY2WfAAF4Ip3RP0u3L4/rHF8zTVXYp4VIjHmwyDTMIZMjUWjIWZ+zgfQ
HhEbalvFsJGODTWEjSfb1RnLnpfmnSGDNpH2vWfJtZAuIPoTasgIGG+tlTdz+VD3
Vhh9pTCw1o4742IYDHlNF7LGdORYructA4qeYZYRIU7QLFqng/9v3f0/mDdiP9to
`protect END_PROTECTED
