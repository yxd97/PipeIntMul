`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OmYiQCRCuTZGMUmBPiAbC/k3dsu4xf4eXcY/xI+hQLfhpXzuw7Fq4rnFH7UmKCfl
eOnNu2VsIfkRpb6dNhxkuoah+Rp77cOIHK5EENO1Q39PgSicqyf0y+SOs27/ir+j
8WytgwCR9ihbWLe7mXE4rBrcUYiNJwYlk5ycTTV2B7TEPh4wONQYqdm0iqGfEurO
fLMYQfleVTOIU3YdHrKnVG7GXzBP3Px2hKjbJK3rYtaVpRsTbkEfNjSKA2wiMQ4t
blXdqzfy2j5y812Pu1+EUp6v/EFpdoG3k3cgCwYlz1OhVRey2xZw8hyZGTf10BL0
AEJ70VE6qsj9kysc9+mUNfCzIzVJwERRI5mR91NMWeoZCFbdjKwZiPDzUWgG8IMv
mTIsG7BMn6AtcOZi3brHma4l1kyOglmAZN/yFHnAn+J02HRxX1x69vA9HxXVtDtg
O+KN/2XOQGm60G/q3XZuJ+TJD7uupqP32ZqlObPcETZWs4C9unqLsXFPLW1DynYj
DEt+QHkn37ZqncUeo/jJNkDs8YYWdzfZpZUYJEF88g8iuaFDeNf953rdFjPrpmdD
bZpqJI2Pc0/g7ljTe69/FBmkVR7EgkxxMNWVRDixi3Y9Cw2cDtpGVG9knfAbRNdr
XVXhGAPdTP+dL23BXflny/25I7yOqxiPjbT6g4j8VCeZKB7rnE3BRVrzzCJzLIyj
9Nwr0i05U9XMk1usV988gXwblGB3L6j799yk3xmL9xCf7AQWaXAC0kvHAkEFa55T
vRpLCghrN8yoGkZXf1d5+VQRXLc+TLD8v7sMTtVuc9D2w9eJb6Km0k/p3rf83LGX
lE2No9SO9zJ9yUAks6S9ZZfeuAp0RwpT/NRWMdhyjwAewqADBKDKIbsmTXzMpQ0e
gJlqt2DDHvMVsX5y3xR5TbgakZwWT8flB2PLczDhzheEeyCe7HQTCzccF3/o8WOl
b5NiPBLrnc8MdA+Qz1P5KeJFj7QNONgcPBwLHR0Ie7YyM//3CEzdIFfDSfmYEO7m
2aeEnoLKysEmy4thtnltaRTxBcoAjJuNhOvWBSqKxTbKB3bDaVF4LM5ZKaLdwuT8
WhVgAEiq7f3tCBNmNHCKfDVg6ESZQYqMo9+EtN5/V2PA7YmR527kP00jf39dQUDu
AhY90Mw6TP5CJSqTXg+I5ZkcN7+/JVLukileHiF++Ppkj0q0kUmsW4KGuzmCeL8Y
aV0y842O+ZRh3VI0/zippsZZo8cwUG6/E4NlYaZ2Y8ABn1ZiDAcr528Z6r3kw3KP
vNHT59Z7SE92uqZytmWSKKTo+65akt05v7g+BU7wTnxTCfuMHmfovUz95+2Zl8ih
OXI3M5xc/d+VWEuIDxVLJE8NxDUupTsBgCpwmXY8+YB1PSvbkPxaVpeujC7PVEy4
jEnOsIbJC1qyE+C0j+vLyuk2YfgKiOzO4FqkpyNBiDtuFkj18fzDEZRkWElhIfqq
HLdRCF4G6hLup30PNi+v0cJsGDqWtnrOBOovvKS0W1HMH51B+pf2nDlAhixfLMnD
RKlg9HuQu6K3q9ZD6otKX8UxBsGsCHHLwNVJpgUzNsUSs1fKwMMdAvtWeMHBI3PI
bvUhkrVIkHIwILHqz0QEfcb1RwEL48Q8/ziQPs4ndy0GeIQuzYgG9Ww81F0ymXJU
Np5dJC7TjbzfEH+L0Dc+FJi+qObqygMQ7uK66Moc5UWHHJAvpyyCOtko79ehsk0u
4qz9DBt/Qn6eOagS9BH65R9qqupRxv8iX5K7/VHt66p7TlKxZjcIaeAMD6QVk2U3
OxbT8F9CzN93pZdzw1dblYr45WsfKkQJ+epAd9pqI0YzngiLkTDb0mrUpqRv2lZ/
7oB11/AiGHTjieqZODQAtdJcIyY4MUhZUcTxvUSRQc5hYqAKx7brB9lzYWbJSceA
ZUA+6CAN0IggDVH8jReTThdxpRJ7mHJJpK2/fhjM6Bo2BEI3mxpVgh/XMYoQM0Wu
pNKGDii/YfC+dClHIi8tJwzkOU62TE05889bXDwiPUqBE1hPKjhd1T7erBggqV+T
nEHqHaFtvBuYouIii2htruYagxu9/P5e2K4vqBTDUvbi+yTmE0sKDP3tjtsgC21d
1aKWnfDsgRiFjHpBwQ/xCfnv2RhS03ElxcBTY1vdLrCn/lQXRLyTHkLLeJn9SL2P
dBT3Xl62HpyLRk3R9golIz2E9qbM0BArcVbGwUySXm0vPzZPWan0BC1uIhSu9D9/
TIqooc5RytLnAoxpL1rp7ug9FUOCqIGnxYraARHWV8Vl1HwyaX7rF6cEhXSRCbQY
RqCIFLHFh6dadZlfdiS+Nzh3lWQMrVv+v07UYlq7e58pM4lkb1FhW4wudah+CE2d
zyi8rqGm3NxOfW/ijai3VEdcpQBDkYylDJk3U5gcmiX2lgye3P36WYI13zoFA89R
6Sp6H1htVZwhkiJpDN9AwLp6Hnvd+N0l+s2Ikj+FqnJuuVcafejZFyi95AsflxHJ
zZYmdGts7vofEge71SBsx+N57Y1VRXubF6NmACyrT22+cBWrs/nm1s0uDrT6EV0k
UGf3glSoVVp03kMr9k+/uvcx448SSZoglNOTla1f3YoVsJpmUGwc+YWgR5S5fT2g
/EbNrzqtxDMXnoZ23WjqEuJZ0MHKhgRjiF9eOQeAgAe/52oSDSykZunN2suhgAE9
6Bva9jZlPPnXcNhFUZQPqeyRlY/00lm5j5LO/Er5Iy+wO4fMgkkTVn2sPyc9VTFU
GrYX6Oy0uS/wv1LG9MAopc5Ze7xPdmblBVQAWb59OL1us07wIH8PwsDC+CrmQsQz
9jhVMcwjEQfjaSnaWc5uDCnA8a2CVHaAyveZyE+x36zBYxeX9FkEG+IHylK/DC4p
uXcNAV3Z/AXvuVm45qy6aemwFP1VMO9QAQd4b6k7UxgP+i305HWnL3YYvjkWgUJq
cn3/+CswwJCuDi3li1s7tDS1rEWRosmrbvtM/xuB9MqHVjIUKZTRwvrU5+JgHRE4
mVYwE8Jje+llX0+1kGVkVmlNEAmfOM87S1DP0UVabAKI0PL9DJD8SgCYaHQs5AzP
10qeet82U1OWcvK2gF89B9ED6VXh85jqffcmT29iyBq5GtWzto7lFV1MC2PE8hGw
6bB2Tz4am6lGM4Yz+1s6leATKMrEHOZCatvRqPyz1i0BBXLlLye5ZuzzO+LFaren
uLdosjhQ+IOPiZgGBX3RA6FZLYDUvaACROKyZbSN179NcjhEPSns9yTgnhLwsQRE
qC7arHlEFM2Qr5BfEsIrgwEVn/sj2xt81ts3A56Tdz5ufuUyRJJgjbJQ34Wnl86I
eSSQHbAFwwGCJ/OjVf/Tsw+giziGB289zB5rE6HmVc+o0HiUuh3ae/4EbbpkbfI0
MJFN5m/3wH/532kOx/JEWsh4ihGBc/VO60rQ7Gm6Aum3gasknUIBMfTkkwXqhUwA
01eiARPPKMS7/1oe4KF9pia0IOIMG8xV8OkFmVhGzwRZKIzIDvStIV6oBiFFDX6z
s7poRSn2Omj2HflAeOZBrQ5HU70k/5LKjW3ZE2VIuTPixMqGAOt6FRghykC/k0+9
GoOW4kDRRCcV8WcYUUxFmsfLzF/BhPnMMYgJEhImCK7n/RiOW7Io8HPMHQ3w53oK
nkF9hhhJaqjFFqr7XUhzw98DPzyMyf3XOhEGNWKfy4OLkWRfUMGfKKGULRfVfH/3
1CKIetn4q8/sQMKx6vL2lMpYIgYen5o1N4KewJUdOni3Bj0Bic0tGEepKhd/Fy8K
+2rtxGees/3MdTSfYWdAP/UbqOsQkEadxtxH0so4FtLcJhdYaRGw3OLBvXDeKd48
hSXK4nFRjQt0MmrFXPieGR/EX9Cl8KoCM1LxUiYJRnpwDC10QZSJjSiPRuRW4n1L
ttVaarkXGU8NT8lsZu5DMdxkpQJn4aW4SBKKvJJqyoM49MJpqPk6EF5N1+bdSnXo
TBR3sVler4k5o2AgZ3Oh9HPQh79bRq0a7JoMGJxEsxqTLj/FbBThhN3V3busDNJP
4UwHjN0DDE6ZQYYPWjy2FJ2zc8Ym/rlNWQAXrwJbXR9Rcd+XTZg9611TVTcWne6v
eq4+f5MLY4BgMTr3vkQdfII9RVKJ4a/vNGAQSeQ0Qc+NDXEUFTpzNxY2CykaMIlF
uST/n17J9nbBCIUdEUXCW9ieE2Tmxy0Q2PMnXTq/W4E7gk6ooqYaK2OlIQcDaft5
IBmL/MPCN0hc3ibXc1Q7kyvBdK+SykTrb2hlXcB+jt82/veQPMMDMyJXGu094CYp
Tr9ZgFpetFzILc/zDAW4QhzG7sJ5PMfBfMrtKBefbR0pXR3zVqD3B6pRV2hV4Uhh
mLlDsKNFslfbB3OIxf9y1VeSxukeqOsOYMHA13n2zDGGD7fV+2hPcSTZ+HfcTlm2
OGMYf2l+R50VoXmmO4gCpRTqIWh0wh1rcI40kO/4KSUY4fDUSdtM/qAlo6OihpTc
4n8GM0WIdGAXe9YCezXDVK+qbZ0GOoz/eFbry4DycMX7eegPybcQOFhTr5h8nEug
ZyTHgMkBjbO6GRQkwkrkRJQc0Ht4qz2kVVGkurzZj5tPaEylvMsdTvKdFmYfV4/H
zhwNw4TttqOG6ipp94+1AuqGyrxZZE1biVXry7/BEnBSHOnfnIDZBoYSqI8eW/Nk
1TnfCwR6D0V+6jbm00MNujn4jcE/ICr9H+3qKN5HdJWCrTj6tS3ZeC2imsw79GzQ
cgd4j1YdqIqSa/Xnyo1YDKD5hyCFXUcopwe5HSL52ODAn78c25dSW6aYOSAsR38k
A+RW39hR/ZeQaAHfyzsu9Iu7KxxzsOGuna5xbB0dfTi7GgnIncvODNkCvw0qeLcG
UWQTjWi0yE1vbqhRuogkSAUmCD945IaRQ1cf7OGjSjRbdVJ+Yii4a9tu9VopqfLa
PDuclsw6SToW2BI3mLBOcYXjJwuOekkswdAq5uryOMgbBJVXO0XpST6NVzGG5JWU
a/0zGTSuJg2BR8CXXPzW59/EGOVEEz7K2OOasvEs1gnfOBo0iq54X5U+ueFI7bP9
yGrh6k+cbHSK18yJx9kFvD3ZJVI2MLhde/xku/umTUo/XIv++Phv1CIwy6Mt2br9
pIx35IzMTMBO4u/kXnY8Q+ECIAGguzldFNQA11VP2tz8erKjjg4waGGJTJZBV/MX
ISh/AvFsdnfLa0rJuOcwxO8B669qXSpzGAAY67ZCH0Z3a0y3BfNNAsvTWAkXJYBo
2CeIGi2A6acE4aj6L3Ll3CxlTZJ6EoYqHzB70QaC7mpNf8Eqbl5SD3Nn9fDYzusq
X7K7Gm8K6x2XkazmxSIMZApRez8zm//CfVgNxxS4yIycNt9GdT45oKAf30iyMw82
dvcJX5NnJD/aQKcZ1SUJONu6RvN4m8DWwdpkvxB5yV5N5s3/pI9Kk+Z8vllbAW2c
3MV2YBh1qBNJKkytNPlzwtw3E9N63sVi/IrWAwHbji+yjgPy3a2idGBsbgog5Ces
Ks5PzpNPySZM+6By3ooM/cxgl3Q67uhERZSiDqglTuPmZPPbVvESYjUy0++WL0OO
6LcOo3ml/uVLPipgiM3lvuVTmsakKx4p9qn7QEqJlaPANDZsPpLSODAbykMSAEV/
jTsQI3ktfrdisOm9eC15fLpy6ME3GOOEN8629m+T3kCmkk+mTAfCsknkltWFnH0M
XCwkgZYueBowL1pW7EXz5veTxJWKRryXl4FXPlFDurFUl0JYo8CJGeM4feMtT9+0
S9uUo2p5s4kglgOMh9LvGw6sMp+jjo9lBkZBOuZI9PT/rVBxwxW0/FinWTnmW6Vr
IlWg8vfTnqRK71XaNX0BiPU/AltvDxOXt3TgaD8vhatHax4lXY2s7KvdQuCV+3tA
8xsE8iP2CDXtgGBm/9Jf2YY90niOh+FBzh0ImW7X2D8rax/7uB3pQ+64SXTS17hF
dZy5XHKhf1be02BfLezda+7MjKQMSGzEB5oSb8QsDm+0gBCRTYfmy6GKmIzUcX+X
pJfjRI/lKrbTU74nkm5uvi7aQcEl27LsQjZqIm0KRyV7U1qqM72RamqZ+ZdZ72Xc
5E4PbcaSG60l5A21JTn9A7ctH1wzD5O5vgDzZFsoD6ViJMkNTKjPKeRfgeD6+SUU
kNddZcmgMK2s3QAkpGXHbniyksyn6Affc4xGwnz7/PHGK+43jKuREd3xTPQbmkLB
8f/dgw8Q85l4Xsd30I2g5qmJk+Xndd2xVI/2zbwf5zJ6ZKwf6u1miBfRuYVNCIIx
Z2LVMh8wNzVoO6wpbn1P2CGcL7Ecb6pkvzVSIA6N07ElMlJ7q+WT0ohx6npxdVBf
c3ieCon3vQNkhfREdUIbnYAu2niaDnsCkcAgXmQ7L1bcmiZ/kBwwqefiVP5PMpa3
0ZKDb/POp699sTyDrgExPM5vYlmTWTXISVc8uY1CsPVy5obrJ3EnY0TcO3BwQEg+
LewPM5eSHyjahgX4sOukM4gvMJ8X8cDzUIw3m9OMW41Iqnm1TZCmeI25sz7kZHuj
RhErZF35q3uCbWLrtIm3pjB/y30+oHNuphS08xxyQChvVPf1ZdF5veTpxIN8R5KJ
pcJAxIlF9yIFr2cz3rAkEWzEP0+Tb3c+OwobbL+dyYdh20/IA9CHip+dwK/55G4x
SRiKcOmfboXaoe3S7GcgHgY/TGFJUJtLBpBCTSLM0cKRWeV9pBEKqIzZ6Sdr/b9k
reATmrEM5uCFQR7fI3s4k2CYw0/T+d5mO/Cg4a/IQUpelo6uqJS0G6OfCrAUYbYf
xbDTbEHJEPSNVhOJRir4mAyeG5s7oOINJQ6ubMKOTTijv6tzZZBznKnZ2L+B2uC3
2FbomvU6IQ/rFePymFwzAmg43qL5aGt9djydynHEQ+USJ84HbaFot9zMaIkfZ73y
vlQmcee/4GPvQo5Y3ptz3IWAccdgNLTb0k/qEmEkalrVrEZSm2+QseJcVZkZFWsw
W1reNzPTif0jLs/1GdZF7m07BZRAMDjvApbeiS2en6LnJgXKp3sXGyjtn1FTeZEq
k/wo5uiDUmpr7cNm6OtO5H/RqFY/ckYH7TvLB3Ohs7LjGJJv5b9lCoJK7feRHmLL
xqCkx0vzNw8eu70jHMe3gTSMXiPmjXQ6SkvOoaO2snTQt+46W7PK4h/LgoTSSflp
eoqhXRwX0Qkbw9j2FtNBlPVptG2s51n1XgaQyqcwk4I5J1IGf7FSvqtx+ACradAF
3PM4TZw15ndj0WYdsmHmXSucNA3mq8N36qz5PdenWaFZNmDhCOZAYtr8n4cI2uO3
oh0/UcmqFnAm5VwKxid4/CviFAUiR5PafoqSUkjNTFBNGmcuwu/qeV14uILA5Byr
OkGn8/vl5TvrNiWspNOaPSWpOnBuLsChD++8bEQLXGRsMaHtN1gVdXpMKGJx+cNY
vHgwAetxTjwWT1ofige3kwUY05Ga4ujypEEAvROtYpMfArLsPGG8xBw5reZqYKAp
XBLYlDNouNZ4s7h+itkw8ZAmGHyWJirvQ4EyXseTTnjE+xYC5F7ugtw39omM9ucj
pfkoDSAhzwsWD9S8DywRW/9nvFldT5eUdaazAG27nwN0fhdzU3BkBM5NsQa3WNeY
QoJfpLC2TiSwpIWYQjYxbO8SLcw2bNFXAl3KT2+Vp5dJPz7ShY/wvw0R/dQ/9kdB
x0tQgAeRmkod66Q2J0J4D0SW7PkalLkTH+hvnv60Tt2WSPIp784LDyAy5Z6JjfvT
O+zKtGyZ1JdIA7JVEfDMxHeuDIfQMAXWoMltC0nlRPgRDIxtFkzQiCXCNTFoaYB7
rbLGP23Pzun8DMnjv4iP6wflKsvQyCRvL1Rw5afs3vCtiumu8uqWs++kVgxlPcjl
k7Ro4xyxEUzVs3FmJnBWcW16stUSlJXOFP9GVKg9hob0QP2dniefeNJUNSX9Nefs
1kPdCC9VIID2/dO7D930Zj2I9jynVa/uvApEAGDgP1Qjm/Y5sPlCLhN3RdqVsF6K
qtlpPoxDw6+so4KEBi7JXLZ/VpL6T3rsO9Q3+rJb2HMDrqdvG+O/JYyySdyOR4LC
ZYV8q5Q8zKGXi4RzNGSVSoCwzVlScctacialy1NsjBEBYbLrNIQdPo+Xan01Kz0y
8qZa59oUNcLTU2LbqKYOjzY7R17m5WT90DiGK0W3GHhSva3W0aajMtbJzVoXlckv
Et+6GllryaHovEk+u+rJX+PotXHiSt/0uQdxL8FQWF3mTRVY5IlSgAwBkjhGBN0Y
G7LK6RXIzkuT9hYZewJtHouSJ6eCS8MpHJXbQmYOmlDfQmL65kwhNsqGwaBaiYlg
YYEGv107HJDA2ns3LfRAcMMa0OEww9fTUghgNk9+NtxsMp3TSVKP633sI0crHbdg
eSvg2bLieZGwFGuy3U0GB95BAUaxKbjSK4NUQIalhbdrELeyloohqZFj6TNnFPJb
rO9q4QSiABbPk4omEQi/4TX+jHw4nCbdQLBE7/Wot3UzBuXRLXgURl5zJ7SrnfdU
9ysiLhDOREGpTbxiNhkVWZdMLNwOsA9P2wfH8M+KbQn9uP22udqgJ31ajEw4+q3M
5bsUB5UP5jvRILxJ6eNeAFPumJmOcth/g+gZHTpaQ+c9M0EUnOCiTEgVdFxpqNI+
pHXDl6J4kVFRVFTIS2Q8B2cMIGZMzZixGX+ClplDLMv8BoKymYtrjx0OhJaQzBAH
YvaDY2a7KxGjKSKDFH7QpVJvaI8Q6B7cnKSLlnzhR0qPG5VYu76xGawzNWlh9u+Q
tV2jjKbqUCJsuthScf9tHM9FNqGVZdoHsEM8qBJjsaiHfhpF8wyB8sxQm8mtns5f
dVvsr1Q+LwON9u4sBv3lwye1QPhA+aMSpXVzYEa29hBr0m0UhC1pgkPqe0rh1Arb
WGqE8IPr0QbOANG8zRxoeghMWCfzUQbmLCrb7rWKzrkTcxwJczxxB7Xx+H8QBmcw
poMditJdRDaGbwUrfQ0DWvrUUyjW5bxNuNCAZk0vwZtO/7RHLkHrt+BFJezH4+By
VN/r5uORMfS285R3SYWnrPcW89JtAuEhII1YOarNyVWDV+DIslqWYXWZiLV//50f
+JnyAnZjbiElMQpEyNN9jfJXJ3AhqMjbZmgK1/zJtE10c4lADav0O2tDVaAlJmF+
M0gqkMN0onXQMVw/6JjDxYHubWXh5jvr3GRnZ6K5b5uVSkQ6b1x6Nxjek9FiQUdp
D8l29icLhxx+gybmCjzEXM8K+Cii6JgiPTuARzX8ZWbBqL2vPoilah1bFMy+Etqt
KQN0TfsohAxWvL69T4+hT0L4+NfP+S4dJnkmQ5ZVNxpBOUOMp67Vo2MK0be+Wu/z
Hzxb+5fHg7N6v8hRBOEDeLJvrlDEbt1TzKLJR7m4gTo2l885iAojD+mOHDO7TT3E
asJfSdLncwQBtBPawWu6b6rNfbEvsk7vC498wFDNuzCevo0vbpncEQ9zeJQV96Q3
UKS6JuWfKuvgARx01FzwZk0DedTpWw1qnWRpqCB9BbtIW0HPaUp8Kr/4C7qkbEBe
mLcM/yOVnKqxbGww6KsHpEs8kG4xoxjIIF2iffTuH5kFUCNbHSNK4TjPOp4mmbKh
j3sQxncncGf9dZJ0JD6XZO0sWMlTzhbKMxKBw6jtiTgCFqwHZyNq1VcPxeIny2/k
hr7xcWPG+ZYSlf9dZzZ7CBxGe0aO+qfE5QDrL04rwbmZ258+lmrDgfHp52f8+2jn
eHEQULlZTnhKH6dyRjya8d3Z+qwHatasVCKMQSMRcvdLVJf/o8kyq8GFYxLJ5DDi
irnuG278c4/TbneMkSEKw/3PuHbj+XDwe0+g4JwXk7uYu3kRK8Pd76w68wD17+Ho
o5xz0z2MKIuFdhnsoo6nAkAb4/LAdxWmenInN74jDd74F8zsq+QeYEUQsuTX5+ap
VqNYc9d7fyrzS0E2IWg+tl9Ps61nnlIxqFj9n853V3zLyEiTZqZ663sSGzLPuHQz
hRMRHLtPAPSoJ0kqCBl5a4hPjC7ckAMbMwspU0rdRvXDJ65fcc5hGtzh0pjQ9LKJ
doAxG//A3Khrvow7MNNoSJDKJKgFNavOGqcHzrBoqwRHD2OLkcQCdCZDG+NbGaaJ
AfTR33EiYozCGT7qD0nMmnbq50HnL+rMbv8tvIsDWDUGPSG4CaGgEYEu5cLkLJep
XJNmM2KJTuLHKsAfkCdHw//3Jt4ANkoYclj4O++U2v90Rsnw7cQ9vC+TWXG1QFo3
mblc98tIBunWrZxNlRaDWprZC3h7uxo4iqEaBwfbfFqBt2ng0sJ+APKo89pGwKMI
nSV+TjWQLCgCeTmqUr2MyRSgD+ct8wmVvtX9PnLAt5zQ1bo8WG2cQh9NcO5Z/Rwf
3FAOko0avjZgjAPugpeE7jzTEhK6/MP0n/otylzMzqrVcS2y70S8dDYREsQHmGyo
XChmmbD5pLPG/hSNCDqCaVxQMIp2bJpfuxZJ3+CPuKoIpeh9S6VPyZQkuJ7P/bUH
AYBIa3Un6y9W590GCcUxYbC3B/AVP+SdL+E6uPmBVaGJHPzvjnj0L1oRoo9DP0Ew
HzewCnClhXo//rtfgB1gn+l90yM4jrckyBq0MKtlqZlTKv1g8wbI4mecEeXYoWt/
ahmB9jXIOA1xgxSAxMmwmbqcEIFpMqdccZo2pSCXQI4qmPDfRfXrJ8HVueLuuoqI
9Bp7HbSxoCLqHvB5eHSKqUAySX9hoKfA2fCh0LE3JkcyLsTVpNXY+xWAiTOUik21
dOUP32McGbpuD+lot9avBDf5N58T5qerjIuobgh2xqFqSxd5kOMqka2ORfs/1Ojr
gJUjVtJp0RNhwof5voTjR21M7vZyY6uQewwVaAO6TDeidighqeS0dmmFwyc2cqfN
526aD6ALDBvzWTHngZ2rTyLAmZ6/W4NhsyGOYiL0w6RRBtbss4ZYT91Izx6fDjT/
Xx/ZQC8I4LMks4M2a8OYu1dgHu8/R8vgah48MyjnpjqV+dwaoxxbWipgKe/ypima
HSXcFJYLCxS+r9TJdk2+x5eUw363vSravL30MaAOdAIoXJWFk96OCEyTwlDKsvrw
/AE6cNDE6ILF4N/7/EZXVhTrt/2OaYUYYAIoQh518bOTf+xT6Xz1SwnAovvyQXDB
UPY+nwKAG7XErr1Q+LKRXqe1tfg7s7CqI68oQStf2mf5Xoh6sj99SdWJGyGRdws3
trgIZkHrXLvaOOhiIh+FlVOgJKR0Bg7fm2vnhWnk3JAjNHvYgqV/jpb6jgodvTOj
Znmu2MBb2RC1l60u3IDeodvxJ04FDcbb8zbz/Q1dEtRWxklXXUrncyc3TMSsQTpb
+LLhJ6aJ60+3zHjb7IMUQukMK/hpyE6QmgfiBcuGvP+6nvNCnAqNy50YvO1kKTIO
2QriHCQZ2l6JQ2u6ryCEy6Azf5U4Y6CKexFDJrHqoiJwvriF0/54LJf69IN4fXQn
Z0yd5wNOh7KtFx0XFC6d/qkkMAFBSmF10+FzNocC0i5dkQOS/EAYIH591zjI7i5j
gqlS9t18A3WHSH12EQV1zj+Fc7ioNawTUFLQyvmJVaPHsUR5gWd7thiAFBZ87eHb
c4PLM7i054Un8Gtax3ioJ1GREQaCwg67Bpggj4TvI6UqvEueD9BBH6jSPU03N3Sa
ZL4NOLMwer2kHX/wv8AqBsoUeSzRzsYJzidkNfHDff5l3Irj3g3Dvqa++wP1jR3K
k/jyVu4vULk8ytIYZP13CHMRAVHOJzySTIrWTQxf7/2HPTLTcLHt4+B9tZU4tvZz
gxLZRctCcRM6tE/VHLX5C20ngoWr5hCzLtjvnJpyofJrmtt85PiFi70C6rm2AE+V
wfFWWrWo7E1Q493xNGSPrx168Hqw1kclZGSFDX+9LmyIJc5HHvYnpuHwGu39Kq//
Oz8OzRvup75hMCBnHFSvZDUSfImUcl6AJco1COUy8ezCh14qdiPolQ5aMH6mSg42
mzwwDEb760yA3iuSnMDaVNddjD7KbdGrDD5aB9iknYAcqZxs5sAueRUREp1twbbL
BSDYu2rcbfCeWBnKNPPqSFgug/8PR6j8h2IN8irwG1548eYvV/ThKem2GIjkofdC
PZ+ubMbPXmJQJFwIVifhzTjNPtuOngM0bp89NzhLEcO9/RVgLrtZ3FgllWJmVkXd
Fg104z2QC87wh09m6ccfSJmISURwjUu72w6dRJQ95eAbao5D5RuJj+XhdfRPZR0k
OjYUrYk6BM2vE6BOabZAMgXe5PoeLPlxqiHIVNfHFEGsVvhqN/p3XoveJmswDxus
Fahxyru2xQDPYCCIDOpJlP7vuBQvz6GPk24P+5nBmVjRb9SlbTjHNFypQZrs0QG5
y4jBbeP19Knm8c+l/2U3eRUKuAbgIjARhN9DFjDHgm/BVvD1p6FPqnOyFAkhTv+t
nawJAxxWGp++S8VrOBnWC9bohAe+PhyTlh0jocuTHA6dgL0i05IVqi0XFFKVIJUI
QGj5mDPS7AZ1WEMjZN/FH6Kptzj3pCbks4KhGT38Pn8jMb0c66ztfmntHc6Gj1qH
aIXP//lqvksYypV672xXE5FHcdgtEcUcUivWU2SOVr/e7f9cUSO0qUNmO3Onh7NA
zAVYtDtNG4jk1BJNqgNoe07KK0MIFUYxyI1OsHfKgECv/cgKVvyw50iZIGMwFOKp
ElEZgIJftWiAuDpXYKsNNsp48OIf9ucrSit6QK4i7CamvvnO8ItPeART2NyDnLU8
/6jO9JHkOGJ+pFRlq80O/nrmZiSZGsjlw1NVCSc/jb9S4U/XewUZcLNTYxzwemnO
zjzRPihdBcBGOXUOoLWShCl+3MFsqMjeSxyiSrMZuyZQFBtrZbSUmXUBc/4vHA29
iGEZbhxvAhklGxJjr1P4YN+5WoG3f0tDqu9b/mWlK0vw99xuBFUaEojt5NeewBUm
roZnLX7odgyz6BWLHr39zA3wo+WzFMZXWFsBnDU7myyvd7c6szEzSlNBs68LdZHx
CuUX11yVSLhsnTqHoA+k2VNnVWrRvwMUB5L8NicarS74/ZnuAnFFXx/U4S0R7ymf
dpLQITL1FX3LesVd+vComWH1TO+QH77VY4TmaaBnlpFSr+JvdNlUmvRQh/ic37Ds
O/nvFKWk1Q8cad49mbJCNelD9lcuTwTrsm4PQE24LS5X5Or8yCTe91fDhNqkIxgU
vNKOawyhfkNdMIHbHUCTmjorqxTUnTD2F4Px+D6SpphJKZiQsYF1eT6w7ei5FbMS
3pDaOygg37z5DXzf/DpmbvxdOC0psWjiFOWHyHNyulvTnoxewi6v3nVkw6p1bY3G
EtLAWGHuMzbdA8kn8NgJxUnQNRqJfpapcS1j0oMgVhc9gAZ7yp+nGOObefRMMaUB
y2UqtOOScRewnqAzu/v10IdM9fb3WynwUwco59tnSJ1OCxaenRrMkVqx4LgzUf5E
N4L0Z6IUUjAx+2Ty5eEO2FeBJuyRzCmK/5TJQXn2wV8Iacov8UK0Crv1n5pE6gRd
8hIszOKvsbzJ3Yb4tLaacGsHppv4yOalXT86LwKAUgw4FdY+4iY4qY18fMWhsNa0
xEKCDJbgjeQEOmPYZxbNQbtsentnHyKVjieQK6dT7Eno6LsFBt3ZHlYB+IGqg+jG
HXCeD3VEkWm7fp83yIyPTlc6KzgajC9xMR9kn2FD5/EMRm1ML4Ipn4+6XY3bQ8MO
ROV2rRalMuy4vO7jHpok1eZgIVYsjVV07oWZrr4RPw1Nb5j8Fzmcml/V8npGJuWO
JfLPjPRhcNj/itTrEcnHHy4cnMRgYbwD/z8WOemg9bt2V9KtCKk/dEfpnC7xvevW
gAO5mylomzjHzutOYGOvwU6wNhmE1E16amO9eV54sJa6DCzN70Fp7jJTqXTbH1Lb
pX6ftqGwSS/w0gQcDw5ieQRO6uvTsN8Q4w51/riyJM/a5P0ptRrXrSB/eMeH4T2l
Ll9wo9AaTXRCqO0rGwbfpfFCE6rXbA70ecMbkoGCKuKdVZ7wzYENLGRbpr/TeZmq
F+e6w6r3Y+AUKblM9KDWQUTrCXmOcnYUj11d9XqRw/ry6kZ31PqTfPe0eVYCv1SG
e7V9quHEguUJXj+jM3LxDmNzDp9/rGrDH9B7eRtbwLQPAnmpR6PhmZ/Apyl9DyIZ
yhxqJ/bvErO3jyWIr5SHqzmBzcylAEZ0pq/tVMCioWUoxxxxWVHNCG24dBXXnqdc
UQbpd6pw8AudvpFW8sr0yhqY18kdkNLIHkMnzgFUAGD2iUpg9SvHmtXEFlNnN0kp
75BUuop5L5z9zEKv6YDwRGUjc2DkDpv8Eab3cj4E/YJTjSkBW49U86aeVlZKLAco
jeUBFKAHapv+iUpks9Bd/To7UuYt72veBWuLcha9qTFZmW9C+r7kxRCJdc0jPioK
gDovF/iL7AoxLTnn2XXC4/vFk6/s+qaiv0sKUoGcBEsRAYBkdp7mGampN/gMTcO1
IvBU/Ux1I3aSIJp2t24mKmZMvTktxkjyCg4r6iN6NUf02WGNCAbCaA3iHztZlNO/
eBoKEqCQfG57PXrfVBC2mW5/7o3bd8bZ9bYnwyY8zlgJxhx5d4A2ICnzQesKJ3jQ
cs0PN67GKKnR1dyaMt+TOruvI1891bbx9nvTNqeCgwIMIe1ECLiqyQ9oK4dI6XIF
3MbVDpYGlueoE/BBsL65ul78xqASi2t7T7aSiVVghvjEaEbDtrts6voJMZ90syNr
JM2KypWyLSzYDyi3p32oNmxzc9SCcEytcqc+BGo4jhjADmBJJFrLM3XNTXZlP4sg
egksQLN+EMsysvK3Qj1bPmVvMZO2HbsLpbEAxLBpTKZ6DYi85Q4XwhD+Lpc6F/Iw
akt4U0WWSSVtW0DUgWRrBH9UkzWdHu/jV9Jy4GSOacyOrVdaDMha37yl3uIReQn8
fJvT3JuJT3bDjO8yiojbjaCkuHdq9TaQIsuajE68nelRNfBvffo5LyUdyiUumzwV
WcoFqsdPQejUB62bFcrMnUwiebSOobFvVaDsJRHxLYntu0vlBvWG4ajr739mGSPt
JwY44hzIQEEoScJHEadXOy1oRk0/IdioXqC0+F396C/qDAOMZ7/i4J5L6I2WDCPb
BKErJfQdlC1FsPdUFgsuQkiR2OEdi0GNdf+a9n/mCfZ2Tw1eCwR+HaOJ1TnL6BVn
iZJiIOMTAfmyKecsi31j+jFh1m9pNl/S6bF4T0z66MN0B3udeaQwdsuqNhA9EhD0
qkB5dVCOoAgaTPpiPF7o/nJclbPVDR4ChVib814vQSlYBQk8ZrQppokTDZXY7GBG
MxD/rB52EA0Q1gWIT9lVPeoKcfMbqG+fKqJBVg/Ptju16TfDnH9VQ3BtAh0i/k+r
t5rFutkOOk+0gcvSXKGTpcPC0M/7vlf68FCA6nEjv5T2o8nUroetOF0iN0FWZrb0
FUzhVWX/PJOxO3xNIu8nHd99mZEwFkGYpv3wwiJVlSDwtNAf+o71Z2BlJS42leeW
TDARF/X/ROUUzFeULJH8lSu3Id9AisGQX6KcGiVcFt7efo05SMV4ND8dmL9BFzWK
2at0UznFWd5h91PgnnQiZPbRunDsVqgpIofdUsGwwbQ924kZFOw9pvrBq+E7r6rp
nGvsFHzarurA3yJFh/uR2OxtKEt6XPaajt1QIGg3lZtWFIEBYfY5Xkep6+ZwVdAU
3I4J68+M5dq4gVPHzIt3mjEMLTt0sRDwFFYQH0JAunaY054WUUzD2/ObAyOqUNVc
Cbue/kNNxxIhLKWiiJld+6wLAgOUgPcrnqi5d+s7rTKIbKeSYJ8dwJ3Yni4cy6Xv
tcXVAWkQdXUCclMrcMspIHEpXlEAdyjHhUCgzBRH5jSGlvdvKx3GF6GN6iWq99bm
/dkqS4Vxhj8WnZpB3JOlPZZte0qdnm5VP0ah/0qVXnr2obP94WoCu/OfKpB9wWhl
SEgRQ9nGO1pgcC9jG6RTHxiHfQFfMFeQfuT3eSmlLjwB7sUuaqJ1TbYd4SanLFoE
xGVdzDvE8uNfLtzo4fyw4l4/dRceuyjimXGXqA+PgXLegtUFKfKedGQmvfLu74pF
nulXzVynxl867zBmaBLSEzDHhJ5baDSfe0tg3AA2fl3h5YQnm9hDOytyAOXmg3MU
5QxnqyoWiNxHkJE2oeYe8bRxwsXJMMIrduuTf10oUmZJAe45GFXbGHRbtZqiQe1U
+O+sjp9b+2jtKzb9wTKpAgmlSta3mx94eNAGG6boqEGyErDcq0ElrzDNRpBF1QJr
JrwSrVDYPjdz+AiDiymMnsyPW1LizfN7+w4sQAHNttXHo0x8ylD7AQ7CE2/f+/I3
DEjfRH1C1zjBlLi381HGmZwWNMbNMBST/M7Po1dg9vk3CmXWToMjYsTn/RVKW5ag
4wob2cxr2Nw0i4xtJrOgKnjLjoVOpFjj8oliVtIP2fOOHg0cpkDWCh03phfna17J
KgOUdS6p39d0MQT6n5OLPrqVdD/HZGZz/cYJJKjDxFsY0hvSDT/gqsAlLdW2JvVB
lJZIfgecKRv0Yeur2FD0Sd5+q7JJ2ybyBf2aPK1tDyu2FsedcIsat/g411Dfv8c9
28gAKn1xrr90PrFY3lJLFANT7kAt4mIn5rmfPiEEzk84HceWwkZaG2q9UOd3/K2I
AnWqupgOrJcJv8SMcxWpwgcf2hkCmzT9k8MCSznXd5s6yB1pxQBgrHsvexgmU0Qo
orUYSqo2RPjzFBN89TLQJBl9f20hPDdaRO7VUqsH/6l/P/v3aoERYNsYgN2BCG+Z
3p9YQoQNZBiOpwZ7aeNhWYg08jYjl37rM2x5l3iCmvFbtUP61TSVSKmhnDdRNRgY
3++Ys1F4FX+K/v6cXjGp7F2azbuyoMfNtGw00rh28GfRc9DyI4qKUxO7c0DzEOLa
MTJ/9MaE0t33uKk7f3YFwxvBtrr/EyAshr5p+2ndNZ3t7dIJFPK1jSl+04DQC5Ga
IxjWvSg8RXPVW4lGbtp0AFv9JEO65S46XDU8OiiGsrfNrEuR7iEKxYvTQkV5sTWg
bWVVjUsUKSD7Y0G1BtllUKpZNs+0oRZaL0hUDPEqHikvCI2CXVYQbl0hC7zKlaYR
D1AYM6tYY97IA/f24BJvKHXvTLzkN4x/NeOFzL9LeJqmI3o4ZLfBXcErXKTmNoUx
uqyhzlMHyf+IqRe2xCBD9jhIrLoMfyBxbaMwOJ2A/eq2Ttfdvc/Nyxnztz0WxPQf
zWlTfCWzoJvxsHpKZ3RjMoaLPstwDjYFMhLJrzWuM3igT/KhGfwNHEczEgtlFrhc
4qm8XI7Yj1bwfUVRkXGBkmg4Uv/OcizJKZindCHvMeJsAw6Yn88T1FNxuDbfH/3F
0vxliBwwws13+yFmyNYVudG+rfWvm22X9yF9VINryuOjPFQkfnVeR+K5700e0jbD
LE4axotEFQhoPUA1wOTqiGGwsQSFewLOh6cfOufXD5UOvdEIVCdz9dVvPDpvugG9
8MYr/RqNpdDnRtfrh+xfa3CSBtlPEk4/oKmH+YrUq5H5L3j9ZOVifY2QWY8jW01E
gFTtxUKGojy2+UxS6RrCwn5vU6E9y8NxIE3oGsKr6FEu9vEWIvJprOiwliHRwWWM
Vanwww761F/roPf93F5Lndv6BOUhDuXLVn8zApu2CvZSQl3+FfmCfVTKTY9n2edT
xzqmF+q5ITdBNcIxgiD1FhvuOFB4oVQiUjbu1WyRvnxIHyAnHKsTEorTzHrRjStp
q+80ZiYCNlImyQZiSVb+mJQgq3XtgXHPkn3BYUI4j0CW+8/sXoPeWaGIkefwtxFH
WjFIZdhFnz1qYP50cKzoC4roVbkWhjT9iPGg+7qo6txuEBZ2e6/Z5mAX2CuHVfxT
kHTqfmBzmNoVH9BB2HbvwAXfDUvOEaCoIksDkoTfnW8g9wN0mF8UHWPEnagu3AOr
FhUgfEC2iMFCBOfUP65D1rnCz66fjZi3orBSOlT9oGvQBuaBfUgjZciJ59EmbAq3
akeQ+o85H3cVYoIEM5JlvyA+u3mec5GwqYpvW3bZo5Z/P0N6tVhS/pjbpQoZuZZN
MFhr3QJ4lpL4dStqtFqwOdsvVgLxwp9Li6KoZLTb81gULBzWy9QgK1hXvHDaxEc7
kAoJLPnG7IzAgR1Z6QO+q9T4QTmimFAXWC2Ick4Gnqcm0yHnd4DcoPm9/hyPpNey
CEwXY3v1TPgkNbxNDXl0Go9dnXMbecE1ka3ZY6vf3SfkWDV20LxUIiEToU6JlSCt
wrWvCNqdOcPQ/qXIT7wom7xflhsUzQgfTcaMHHfWJ83IqcBGkAyo12NiWBvN4FiE
OKDRUWc9MRnK7ynN+zGSWeszto3Um5FsU6lW2VnVtCKZvbcw6YwgYJIbZfNIh+k3
NQtPftjnudBrRgnUehT9oihuSV426Xyn9QBQEDb5Z6Jfi/DKKc9s0qyegniCu0ZG
nLafzYDzmhTimQl1xBDysoldA2fgdfa8DqnShaeZAEgdlMn/b7+vX5UZne9iM4Wb
lECiWkC2Byj5/erBNMsgKodVzLQ7EC3tBoIe8Xr+23V6hobaf2kUatqFq95OchPq
t+ZmeWhCQpXK5JcsXZ8mPkIoUyfqMS2t8l9XneXekotc7h/iX5x5tRxiXb70T9AS
lK0CJWsUoydMacPYV+gseoHawtbp/pVFsZoYP84oKfqFWYAsqNrZVo7A1ZuQrBaj
mcx1jFKX5h2OhcXk2bbtFiMtz9mS4t4iMO7Ox7pg0id6ZeolQ6kP7QHMdd6Zk0cq
FP5kKTPiGwr+ISmvbQ64vEwb9ZzS+E4fgzXJdMn69ycdArqcs3Zy6Ic/Z3FQHk/A
AoPKSyReE95F/OqpsIOe5gHuydqoebKmhxoMDdi5wvosGtDWk/79oPE+RMmmpxvD
5xmNZWEL3WgQ2k0SIibguw9Uet9+MwLo//yw/3EbeG5OFuHe1pKU0F2iIJfbpcGE
rM9i78vovFQW4d9HPQtJEytb/BT1cCA3fy/P89u9hsTver+7q5EBtL5jhCItHZ1h
OICW4slRzQi/mT8wNcI34AdCZAOTi0SRe7TEMt6FyIe2Nx7PdD+bmMZU/FNRjjGa
84kFipa+H3sEu0ShEBm/ryBKGOMKKEkysEtzYgY0zcvIFfuCYqI7i0Wk9oAXa6Dp
bYv5BYtWJnV2kLs2Q3n5Y6Co5zZ2q4I/JRP9+ap3XSx314rWp9mTR2PMd7lUkrnM
7Vpn13xYuatp9X62IoHuH0C1vAE2yg7dQ/TZbb13htvgc1OEFRLw7M+YvlW/EFPB
pemQLdvAE+s9zxQkrXCSrSb1F/gR0krJ4+iIoVQiXLLpw3vlWzHJ+9QwfF3Zcywc
Lrkk5Gff9f7XA5Yk/ypEe9fl9BLEu7X7TkrYZvc2zECVvRkQhx8c7jsu/sZbNMql
+4A0G4k6gQANRFwje0R6lu2VosNDlig21bNXVItsJ7tsHJvIa7HkjWRQx+rDKA+T
Xd8+UTsLeXlvgsvci/T8DVcjwuCsMRu3wD1aeeuFIxq3Ee2iJx7f7GYMTMakDVXP
UaXhWzdeNg2YpaTk8DTygbDWHzxQX4PdJsUEK3BjZYtT7J+gL8ohYUjH7l9sSuBK
TBZHPvpFa0YHBdZkNazRTSQyfBkweQUnBH3KX/6tQBmpud8vulmRrCY9zZ6x3xGQ
0cHP8j6umRTooVMLPVUaoXZBWU/0+w59O3Pk+j1GfWOQI1L7bzXmAkHHy62wR3S2
7v4QcndNBfMdyM+70ceHHpv5E2JuU9PMGgIWC/mrHLLaSKTMyYn3zcP21Lr0Pk1o
1nwOgV4x1Onu+ylg/MOPVE4sdupd1gOdvR1Xyprrl28zgitOGShSnC9vmtd+qgUz
7fzazqM0PMn6+ticwS2NXKXhyonf11yMUOamvRbPRgLzkg1bf6ftjq+cQQaeqEKj
9u776N6sxhkh55C4jNck3Bj+LdVrverdAxJRsFGJqX/8TqFI9i1nuknrSUSXzIfG
ljhkJFQFn0CExo7woinnA7u+XJG0SRxfoJ8xXieDjKvmGCI4xwOChBwE6vF/j1il
bzQ4S9oEZ0PgLUri2v1AneNfvYIe7pm4zggDOSyOLHPZ1Q7Ud+ezb5Y+Uctvx2um
SjBJsg29QLtZqyBOhPhXK6nCD0Gjfo7ueLufjjXN8fGJ5NHDlDYN73kmvMEJdSJ9
JTjTdlS8RYnIbs3aJpVwBA4dp1GcijgXgHDmi4Tn0yukag1udxO1wUUhC+FuakM3
NCAWhMLcmf24Q2+Z2k26IFW+oozp+YgsPsVT2fyvL6pr+Rhh3QfRqKWv4J5lbsk1
CpJK42xWkrj0knsfq4jtsQbZGIIMd9uNR5soREiQyZPN27tVIx+5LRPecjGSEy5X
H+WrCAAiV1pTD5uTZU9VtadiEmvd2XB8aItIx8n83F/qgYfx2MjMWaco6iJuiRR0
f9UR7+NzWl8dNGSyru/WcLtjEoxMJ8tTahyilKkEnlj9E62lfFUgvCiCqyotcXDk
bzVNeHsbWd/87ys8lUQUgED9crCglpKyUo100bKsd/MCqU4FhQUaCEHMIm20wmUh
uTKxPaGv6GnIHHimvbajBfCfSJn48rLALLFKQZR9ot4GKbqaLf2uA6NQEAi7mc2X
OmK/Q6gd4bgNg1bB7KHDLdNXx0coweaJVB23hWgFhv/DdbjG9fIrYLg3VVOHfDFI
C0gt5kP8PeaW2KTBL0HifIDK5+yubwkqjAr6VhfW8PNIKmQZPe9Zal7lnkT4+Ki5
40gLL6oU6tjCzlZ9sjt09hXRvWvHrztoEecULZxmzfC8LxAuj2fbcOBrGN7Qbmtz
4rlFpA57t7kLorx3t9BxMWY8qlzPdVeZyOkkqKL2XIFy2LLq8638JkQioLmMTaNy
xlnHP1rMd9d/focEQ/JKCbha2FVZbJGaSMKPYR/thBK+kBwqCV/QPspNczGqXZ8z
Pg7BkZ1H4H00jjj+VnAQ6JHrXUXWYYW6Ieg+9t3x77n+RWiR16t0zFnLYEwL6Ar4
ED/KGEd01+Hefe5FPnmJHV7dkU4SAODw2ooLNSSId+XDsTV20LMknh3+i0IzLN3G
+NL+DX48A39WZlkHh9vrwAlqcs92fqg0iGDIRNTR0hR8fx/JCJBt72TZTJLunuCj
1KX0rqbdNjsKxvMzo6Daoyg9yTjWZDzQvRW3qkA+o8aUdulcSRlpwjP2GVm6invP
H8FZuLLiqNtAOAjtI6XIJUlqO5SL6jL8FoXQqn8X8FFLX0F/sGx59p5v9wSr4/Xu
4fTOR+N268RWVnfVFWVl/A2kq/PN8Pk3B3IXzomJvLQyncTGko2iSJbaUHgqoAJt
6/ePKGu0SrJcWbI/txXuz8q39Lu3aaRUnQwCKbp4LJ4tZhqrFgIOOCwSXIrgLZ9A
RuJObI/kz1XO4wrZ6FIh7P36CA2kJ8+ZwEjcwiwoDCeQ13ia4xUDrpUXKSEFTGNZ
HCTvCgptglJrzcI9Lvgqiqs5hzvIEpkdOVNoV3WH1XRZQ+M//ukvTKfxIxeLm3AP
vD6Km4ENoMWRgoskQ8zFFoq8Qw+Fb+h+JEG+lj6vLmrEKq4tlZ3OO0NoT/dWcmnZ
O19wX9SO2mVrzeDHRraELNd8uQvmx/qN99k6boy1AgVLYLd6PrcBDoLQNFMAciMj
EgxatGJumEyHf/qLAkNWbqOE7k2BXV0FZxmJ0y0XUElLn0ZXFQrXs+/N8LtX0hYA
EApxzpA+IId/mRpEw3MW410MXZSpQGrfyVcnAEyh2mPb4GDl/Hgh0ilAvpsfgwdt
h9Pp+pxPqbDSNP597+ANCfvUbyoK81zPr66mgMHQghUQXo6S2yjKIWV9ZUqvTDxq
854YoSBVB6P2HCt5Jkt9TTnrLdeohqso8QqMxASayyfRHHguXMSkYkjpUlHJ6TOQ
13hKYj0rM2WfBI1cE50RgAPxs7W7c5WRMODGWWOUg7RbrAdsYCX9cbdA8zUvzFnm
4eRXu+s2c2zhjXHKkxTMQiz55Lj+raG2n8JdBoCXBaZ+hfmCh6EmHDl+ij/c2yLu
fcu58uAs1rl7jlWKqGdFSb5XHdhQTyJd7OkNKCwOEDbWqpxYz5gT4YWjHpTuH3Pq
6JcGXCf0rjBNJq6V5aJb1cWz7rJwz5Q7pF4dVHWRUwU2I9j9BpCC9HLQXAe+EjyT
0f0lrW9R5j8z6NUwKeNGLLIedEigYVihBZXeane4vkyqkZ6yqMZWLyHK0ox6SCZj
s9nrLGbpjh5bdfgFBCCMP6KnqhNUsPL7GiYCqR8Dqkb/5paL8NyYlpv0UaW6CerJ
c23ioI3FfW70u1qkJTOOK71F07HkAoHiBERT9DQYH4fWN7C/V38DaCvff09Th6OH
cCgoqLuKLJkwoyXtmdxbg4dcY671LyitxSEXhQ3qVwTA9yU3jwj71p9dfJksdtM8
E0kc7lgaCetWHpy6Qx/wQ43IY0VNeaszxlfXwPT0Bkbny/NsbdzrZaC5T7NZUZfz
MHzx4YWd+2RyseBnsiba1oCtFwjG2mnwP2rc0EW8FHPouP7ClsOWKWiBvs0TehZy
J1xd7ELt0UAOjdgnb2rER2rNYAMmgyaHEVAxxbgaFL4pVJmaDqwRWdNG7jBOalMn
aLfRXcWEY5Xuhyue+eM4ObFowDOF0DByg4etHg+9CrRKnGgFRHylOAFcYtgSTraU
9fxhZFdf3SCy4QT+0bGm1YT8zjrjKNsGUw7K3vUE8dNiFuF8S6dPiO92WajH3KD+
lRjMmdLjv0YnQYwzaEL6yTHU6h8gsVM6q3R/dmJO5w8fIO1oaq++o9Ss2fRvfHbI
qZTwzQDayaErBu9vGczUYvwOttaENPzU9UXlNCC3vX3w0sZ+w3oTPI5HtjTZ6Tx1
fEukO3jOrLrFPbL9pqx+mpz7CH9yQqw2x6sEUAFIngmxmO0Minx+FuCLxpwmY0iQ
b64Tv+yHVNC4/QupRCqWf5DOjx/ZRFldvbK4m4nWadJQInIcYIr0eio1Y78M/J+Y
IxVBrWrSCkLGty04vchqR289PG69Km6/Gvdg/RB2UTu8YKaJU/0Pa4Ef71L7GWfw
3w3ixJoh6bnhYtNoavYvQdPLYPXzAu3ZdY48As0320+posMZ8VdQjMtc07bJT9Et
tVuusRJp/sK1xZbIA7hzVeuMVbwG+/PEwWN7LFd8q5kWfes2l3GbDBNDeYXQztQ/
EPTAYILUL4kQd1AF6cdlHL/Ay5kyeITOmosL1nRBfIzP1U+NZ205GCPO6LjmlIRi
RRoaCNBy/41X34bVe25ODGYcjEnK0ku/OTOXpdgoTH7NYR0520OA26XtyMkOcYSv
yyyzISLcPd5t3oRo92l7tslD+J4O4ZBq8hlW2146WeOgQ1x7PsavAzqjNwFrqHEx
6zVVCVHEl8zmeaPF70Znfx0JMeoCtd3DAzwywR+nRcQEhqqSQ8ln7RllLzn5r9Ka
HQeKPJguzSTL0rDaoEHl5GJZYup2b8m4PalKlhxRy4PVVRNVou++veLMcb8S5QqO
Is+5uoBYtvU1bted6VRwhzPv594GUW6G/OsXttHIR3aVgjXV0PNm6uwOvOH11Fyy
wEeiI0Ov6b7XQiJzQyglejiHjV1AJzRpgjt8vKYhEM+SVQf2Ccye4eMbcoiEbQfw
ZPoZ0n0AcXp/SQ70JNVecYZY5OZ5llkGSx+TIKzY2CQ7f5lNJIpERK+WD13DbHjQ
eGsXq4F7V5NMP3BUzXVMXFg4WDtVNXZiO3dkwe621JHkXOSwEYwtU/oKdxDSVl80
QsTAEcnASnOswo37B7GQUpSZ68qgLiZy72Z+fqOeh2QgRY+bq7l82kVwg0lWhJAj
SWr02vRWrbH9FKnNRRdpOkX0jWENhNVRed+vvm3v6TEF5qL6GHU7agjzgEyfDwhM
ZpOB3lXj/hQFvdrkE7/mK7ejkHEYIv2svSKziccOm9LlFvWy8bfMs+fqSs1+wt4D
croP3+ejAKG06xHk0xaRXihVVf5yMPhSu7iehxj2xOoTXWyVV3fENmcMkyhrjwtd
HL6jTYRcdVBsTyOLFR37OruHFe82hmOwh2UxibsGdRB0oSYTfhuOuzJPczTCN8/t
wVfi685UcwHiHf1dui0yunz2qTZVzDTuQhvVjSZlx1Hm151O4FN5LuAEX2wbNLa7
xekkuYDLmur0iCh6UyL8eCH8kjc9MWr0foUpeQPv7ryUfa0it353yrIMo5P2zRqh
uuVmvQCZ9l0jvriVRI1vyhj9ZNB7vrIRjkBysiQyx3NdqCHKH+o8rQnvyOJVFZ4Z
Ul+SxXk9ZcXRu0ZwIv2F40rObj++7u+nDvjHM3PMv1NKKfhGvwnLR3DaVt90hY1/
7GQge3NIIXifgZHy6D177VQItXxQd+yyAbYH0D82E1wpH+WbSzaDlBDR0R3MYsAe
MoZ99zmk6ioW2zwT7FdD45yrnUgsNICyj0I8GDDO0beAlA8Ipj2U6oGZ0uKkNvrf
JNIEzp2V7xLJiUjCRZ0dhooKdj0qGLru2hXGvnGdJpZC1UbyqwxAm2fYGVVpgvZZ
L8+91mPGyenyP8GZsL6EXYR1RbGC0pXsoaJhqPxllcYFFVp9qfqmixB2+eTnjNuO
2PG00mjB88M0Z+DcGxy3rzz5Y/8sT6yJhW6WELk9aCNHYpLLxnWl+NL91SuVtATc
liF3xXrQX4Ik80h5M7GdFhoDZYprBM7jbt9RYWaTVGTEMFqrYVf71Sqa71KxK3Pf
7CJpnWKsYZ5SWIpsN9JEtmAiSdylEr1y/DT0CWco3cv9TEZoW5SX7NGdSVn85I9I
GtCVVx8PevDBmj7M4/bTmWEAACdCrXGzzQ0xnZM31PEh9zjb0+m4zzrdOy1nLN6v
qpyhzh8Eu7fKaTWM0gsOufc2mX//jo3c2XSV0hd/G+RG+FdG2oX7AfHATVMiPQiG
0kLR2psvspICDPLqwEc5ZjuCTk9geCutyC6obPtHx6iyCWgba5XuZLTef/OQ8xfW
6kbI7K1gedA5HW3eSj4FfK+s6Y3DmiO0yLdSu9fgxMjom+uz4VvOytg7p+6+1ZZd
BpOk0MdlGY4M/PpSLTn95H0z/On9m89s+cNei2BiG8qGRICG43Yv7q0/c+xzyRXb
n0Nc8A3aFkP5P1rMh1uM4LAdAR/sdw7Fqr60oX+1aDdjKVy+MlLpJC18z6dDncKY
FhI/McfZdHeUAAJzzIKmKTDEkHPu6rgRnwXwULrP0JZg/5tdUxQLSDfj7tJ8Bz6H
BiBEW64aUBiLke3D3JX3mGK1qwHFD1J/if43KIZEf/R/oQOAJcBK3aAOBUphCvEF
Cbu7n3nVF+45HyJ7DJ7bovqiO7PIZWLGuk2/y6ys2Iz0K2/lAKhvUwuHtvc84fEG
AQovhlDdAyfpq+euKOzy+gRH+oPfYcPpIswUJkbnjlWg3CNaYp9f2pL9Njbtyrna
E/W+MSFgvsbJ8idBUqLV5QtwR3GBu/82xQe8GbZu6vNgEj/WNaABrSX0lk/Mm7oJ
eg2WiD/zcetlJc50GtluY7DkcZEtoh9LoX0725t5f536ETkO54kKSbnJfmQwgeb/
46oO7LmUDQ3acV/hMe6rwcgQb4E9LBuSJZOx4CAYQVOJSymN+DkkD0+IKIAQrvC/
8yolMOuVusDwBmHtjMysgblisZQ99yqmYu78t3topBxAUZB9OSFPJsjh6vgxMxY5
qUUxxwcPnhXjsBiHUD8MJZWexteRnykYMf6T79rO1qv1wvpKI7bDiULRPdZ+p1Lp
S3K/C3cGxQMkiF9XGKPHRZk2AOEk8UKj0pTH20X0GgTBTwkiJ8bf24f4/ZYwY/td
tm2tGMQOWH7Nn4JSY6gi1gcWlakzxhSzs5bKxGFowP4FSior/7+xUGYa2y4zxhbT
qT8rt5cdE6Hc4ziPj+SkwX7xN/qSLcYdtUquTFT9L1bQmVxsat978FMgBy72P/xY
DoQyYx68oF/hS+gGCh1zbGkx+KAosB6lHci/hdZ/pXy1HIOBiQWy4aYqHJWJGdg2
ys+HbR9rY/02cI8qGFHze6fQfrF9CkCghC/M0umcCKDn1p8xfCbQB6LQvFqMJ09k
xLebi5GWw3rYiLMWALZ/medVA1Sp2ujIa2wGqkSDma+U4NR+VuHFrSinEgVvJGaY
CibSGAITeAvFeaKoW9xhATw4QhQOIR0yHE+MB29nKQvLHQEuxjMyP5C49twlSXOg
P6GwVNy82s0XhBOUAh28s6fWaVareIzMqJeIzzCfKO19r3E1fVzRGLDwG7eeewF3
Jvdvaz7TQDwcWjy9Ofh/7DUlDNKfXjNRJKdBz3oc9QXMbAurfTtsXC9jpdeT93ZP
0V/CRj7TJxjGTLw9oiqrfZqdr3X8F4ar8SyJmDiAI4XOqvQDO/Ft2ikKKbKitdin
hfy8wDWDWbzhgoLOVgRzjLjHk4/xyc1/XmHrFg28bEqkrtBdgq4hqqim0Oy9mveJ
iJhAINrMhQxoJTgMbCOUB/AHLS6nq2w/GwIJ5qDw52Be0iktH8NYhKG/F24chtQG
0CZHWhbjePPKikpHQnbevtWGs1shbT0NpcDmiRgDYndDpFzaPk+ZtSOSHWDT1xuh
RJudsQT0zSvsGHUaW/Bpq7eM0fKtESNuW5wgCi6+EWRjVMb36SReRWWyzLlQQrZt
VycTF5T3Oo5eUH2Z1FcalWaXxsh1Fkqam7uXnG6qprILX7eR4z7XPVbR/O3r+uFt
9WM9Im+RGBuoMxjD90iu67wAwROe4xkWkwiYIPHHdXowY3TWcTyKvLFWerIGmjz3
K/LLaJ3XdnLQuNxpWTI5H4tAGtMaMUjJzFiQZF4B48w803Pwifc53rVgGsHF6BD/
XfZ4j1eE/Pg0kt5m4Mvoq331OscqRnN1uNZuRAFltKykGv5QflcSeliLsjxOSryr
Xg1brtN6zfPBamdbzlWa+U5/cyRhMMC7uF3K3VcDHPZaFoX38ST5jM/otH3hMP3j
4SL0c9Gv+fwQlsep4812kzEHVmS+Zfkuurt9gcRnXuJDfWmJm5ICJwqWcw46gK9a
9B97SWKlQvodjtm+zbF3OTgEOQnvxbs7fuDIlfpwjbMiBcTdZs4osMZsv9S6NxzQ
YuOS4Kh7yeqVI5NA0C4xnesFHT9AJ7FJ+YSmTvakQCPKEqx72BxgJSwDMmQGNlLC
nqY/kgQV+AgjNGASo6pNITL485LBWstNwv2MNOxG2vbML3Tbn++VUwWsVMlL2nNO
zK/xo3hcJAsNhjitP//HIRnIF6YHnQnn1LO8AIQwR+5Ez0AVmgIkkoALICyVBj2b
m+e4lLE7HOguC8TS5ySIYLXDTnYPL6TvLYzuo1U5vDhBWr0EWkfcdK7afmHlu07m
7IUO2ccQHQBtbgM/xyEFtSxDEetVeHt5BEFFndDO2rpYDayX1vze6Q9W9WrHZgjC
P7xFrPGwny8ACqnkxPFcKNNtyeQoZxvwnpv4j2z+8pe7SyPOil2Yz18rdIQoYDN0
CZ4rnLPuAp1fXZdDuBGg2dGlZvqPknGAvQw86CWuK5WBqQj312sSVUUeXNGI3Ccq
4Vfee/BI/Jt0L8kgtXvrOEzGI9cPDUphSvSw86nBLOvUWTqK0Q9fcETErXqd1uXC
iMZI6pWlYNhicOQmL53xVyjbc62cO8q89Acjv7tnCPHvcKzUUMOFSWet7Rx6hVgN
9E6b2bzZcKx0M+SPGSd9baV80USoQlpg9IQHYmiaUV+GmuBLng+QPGRgVRA19chQ
kChBQQLHXPBsQn4eGjVVnIkJdGzb3n67HrCvA3ZDabZCnp5Y+V34u0g41gjexSh1
Ei+klXfWlfNUVODQV+icT0dSz8KxwSaOALXxinTSuNJkCT/CW5A0YubtcDUBgq5m
fUnYY7dS7/8ON8O+AtR5zxCe5xDxzgzD3Z5wed4xZJPCbALk29/l18r9Jg1kR7pe
oTf1rUEeAyYUpe/yby9BaH+GfpaNyC5OqgVEs3uDUjZxdN+Z1dQefb0yqazk/x7/
SLQdcU7XHTB8AkAsQ2uh+KEM+y39cudT1c9h0RpxaxC12nBkIyoKBu0yGcMfRL0L
F0/jPf5bZ54KycoOKRF1nnqj+0aCVzx09R+oRJtFbVFV/OUXwp3NfvGv5XO5yILZ
WK6PflCpGyIJV9MJDaMHotWxjeI1QpKfFN2SC0W1io68+UhFlWp4qDMLfrr7PZnH
IfsdvujBlRH7snT/c3drqAl112g4QYpZUcunqt+B21PB/s7ck3n+iYWzhb6elnIf
91GhldOSoIH7N40FIJAEwge26LihvAcw7XMTNAGNncRLxww0OBEQ9pzqeSo6WknI
VZeoAt442vHVXfpR78pUKfaQrEKVszbY4mXZoGrb+LO0tZLf8loDURmTi3J2mwth
PxHtQ53E9smc980RDJNhl9ZV7oKpNnbOTJdmdQDplCeDhsV8wp/i9JxzoZJkiYr/
6sye+2kiUFPNKl2Smcf4nBQcZzz/7Tpw3OZg9YidDcTM3bNHYivABoEIucHqk/y+
4/CPHrKm8QTAqhWWrKUZ1nhclEdAY8wjgCTWVx2JvJOQLm4ZZgb8UX5edmShYTzl
DmDDvrHfb0rtZQBa7OdWvpr0qgayiq62UPkmjMO6QXFYdCsxE4R3xUOFfx3tZ9j0
ZZLjVQnUs2Y3Oa7tfpTj+wgKPRgdPZb06Z/YNOCQDVz6isWpB4VXtNvF/pV2MTbD
DLkbVRxT455tjHiw/4ccL/hAAtlmS+TCaIEFKYUjTrSQA8dxYU+J6WgOs9MB+HY5
m75Ag0zmkj21MY/OQIBlQFKx6VsAHiHipCpZg0FOgnp5pr0tYeSozHfq7Six8yqz
N9K13eBex1nhuV1/KVhB9xk+DW7NYVOr/rcStLMoEWIhcUKUrdcJzjfJBIl2QWA1
r0cJWaZtlgXlmuLyUIfMH+khYsjhfmvEIO3xPFdY2d9ih9jNbBN0Orqnb5oRd7N3
Vp/f0qfw8O4y8HimNQdx8+mE6Z+ROkOh1bFSooFluPdaTN++Xxkeec5RM48Gpk6L
2v6iFGNs3NRBoSxGRh/5ZUuFVmeJzWMvMEHGBfGnyaGUqBx2p+/IubUG6b26gJsx
K6RwpO3y3m01dpXiQA3/hBAZcE/vArqAnui5cmoMCWjiUcUmdLyW3Euw2nFTFNRT
k9Vd3a1rvtuhXKfmtjkl632e9xCDEu7AsbiXq25q/02Vg2BaaFE1G0/gd4qGKf+8
xBS+IiIFnoB44eF7hg++1DmBhn/tgyVBEqrJ/mqULxbf9oy9SXt0aY50qi8ivB6B
S+ecyZB9klHqefJWS5PNdkX/7ibtlKvrY1UFq9dvn2pGtManMATX5zo+4JjDhuhf
mTN2dK+FmJbGvwrrRXqqJyIDLnLTPEyWTQqWvjRrpOIX/4fBOoNzJDlx8pybD9ys
5epFKNNsJ0ujxkaodGAybsU7infmn6Z1sdBfrwzYQ3W0ba2NZQKXxBBwCfEQZj4i
J4wE/SmW71YWO4jxkirz79xEH0sv7hnYCbe5pMzP3EapaU/6tcgC1YUuQ47WixN1
fCX9izMG20UNT8/SudtNX8+FS5g8GVhsvhBQGztTgN2pAvDrBlPYMrE5jBJzVCmT
/EFBr8N69gnHORzdaypHpfElfokD1ru4LH6jGiLrBkisDrBHbQ2Aws5ZiGQ02I3p
4N80h+WtPG014czoceuTg8HdMUpikhR6r0Syc562kQJeoO+iTQCVBnZh5oQTMOon
fjqugBNGvmGDB8R8bgPqw5EMmBmeeVusaqpFb4Yc/oZh39LU9kxqh1UdmTntX8l3
GV066yngwit9rWGdXKIBupLEMFfNUl0J7XljIs9iKV2VXk4JVgxy4QI5j9QdZoW0
r5AIT8IxcH6kPYfQjer6u5fEhZ+YR8IhIDHF73chi9AGnoZqU1IONovMhN/pLBkn
Ix3O1UfWBCTDC5p8A24QGeBPHMgsP3yGaTDKvrdJhwuizuHHP2WKK/rEFcXVhBIo
wtB3zQMcYF7SAHAV9gAI1YfcxqN6W3Wf+8cSQTtG2R5OJotsvOnlvUhmx8EBLy3w
L7EHBiVr46Zmp7QCOLKmX0eXwcihhahwP7PlUzieCSOniSOcDRYckd5MASXgfN2v
IUTKIL7DW3HT9dVY+uMQ+pm4SYXCns1eVOcZ7OwKqU0ShCJwcnft9K3vFQFZ4uup
mXkBtumnqadWou6JGzZkb8b4rH1zlp+VJ/0gC7axT8Adp7WGl7vflcHfompkjSXk
pl9kPgQMWcZkoLPXmMgksVBi6EKO+ITxKJ8OCEfFtyceWo3D025grWlcPSY1/loF
4bRIYRKwPppkiMHNEmwVAP9ekqpNfHy+r8oNwYGPBBbR79AbtFRg40ubywHSReAY
MPgqB27LgtcPjtRhlJvN8vLc3xQ9V9OiYhKLcOC5dWU1T1eCmQste5zD8BZ0SEGZ
HNo3n8VBRw4tTZSdD+QNDrZWkE5NO4b3O798eeXbdqIXbHH+iZyOoKfsbhOx2bAD
Wf3aD3AHrv74HBCd9W3XWlY37zjBNu2ul36jOBQEjlTDekmXdq8I2oKko4nptZVI
cd4eQPM0CZOzn56nnsQxUrn+KJrjDF8ueT31unSMBy+ViIjlSfXOFipy02xbs0HI
4y9SznkawVSVkRiTPkkVcg+m09qi1K3prkL0uoHpokxOpwxQNwoTHiiV7oZLjdXH
L5L7cJTiJZPeIUf8IX5ltVixENrlsZCJIILMV8hKUyysx9keQLN15y7iqu0YmgJl
4sXp5C66HNWXLeAkO1ckWW2C+GIRGvoWNd1y4t99CH9VyuqHM5jWD3KgCMQ7RrVV
3RhXW2Pg43tWHKZT+5kmQBvhrGY/YyVNmx6xtKsfNU4ae1MO0Lg5u6PaVWU/lMem
dgv7ym2hj8zw3cui0zb8NyDUnD1iSmlvIFkhHEYK0VntU1fFkh9Rkh1XNZWxjZNn
yM1irMH1ecNt/YRvQG4YD7LEJ3kJ01IT+q3y5y3gI9PFP4n71xgvwEXKKrjnif7k
/DocsLcDgKdgI8kJEvDyyMRTd7/XmdtGMPCXnxXGvr7DGOm/rUkixbZF+LnCBpU9
kS1vrXo3Ilx5HGOvNXRtuCjAhGU6LYAMdQoP5dlh2v7Hy5Xr6/kBsefwajIRIGTk
bU4Rklb9vRtlhF+IN2v5JmBohnqpaqW3/LMgs+7VNe9WDtszxF5QE6ZaVdrf5XPD
kttz/6hfjwxyY1QSbQ7PoH8gNPXyrdZ/oCrSOL/vVGuRRtK4rI8To1OnHnXaA22A
SEKK4n3X8zNOsj5O53C0t0Pa8HDoPDPLC8KdcTTaz4pKVwifPSu168HmBLMFPcov
ilaL2Bvq7PKKFdLZp2HIgOZRpRjMGcdItf8jZMwZ5nS8xKkK47Q8RaQ/EPi/0J5p
R/Qn6Jt9wOeNte3yzAewrU/lfkrdfbCcHMh+xglVo/LskVEU8FMtDzQCo3LhHu7R
RfVjobUdiDr6DTIJnTS93XaKr3dD4TauhyQ/p8jHKFlqMyMrSEIFO8LnLkiyHdmk
xaFiS0vdzAyLTitLqJQ5jnpMoctZ66cJ/J+8IhuqLswe3rBPLUfapauB/I8kktDk
LKRiCA8gJkEOT6PaobCpFe0RtyjhS3ZvkEfeJfMzUzlpiAEtSk1DjciNubHNggQV
7zWmmwNSwnu80oHumYG6fMMFvNyfsKP4j5cKM4u7Z2QQiEOUp3hN843bJGrQG3+k
LiewH2oecg2aaSAYH6wTGDe3eL69YZX3qcFex7UJfbIOhBKDx54Ftab8EfCmsSTD
qRhMLP+shuX/oa0Jv4tbn064X1H3yGICVuEZ/EVs8c3eHIqaKZiU23GGNuq1VWr2
KhtXH4NfaXgdjNrc6Eyg1QrJKlOrCokFzXDSGM5haDZdnf10kFHm6W9aWAd5zwHY
FV+H81TKGMkJHjJMBf1Viwo0VpW44ihmsw5Uty362j4scT4yJMY7Yd9AkIs61Ew6
+BnUFcF5divGkXNA4BEaU9n2CHesB1/42G7wXlzi9ESnBzl7yzjba0hxT9AMOToU
0v14GfHYsjBEpum94LuliwsZO2gGHZmqTDF/GDv2mrR6lVOPW+syXmJFhmH1rImQ
jGSTzHbTvS2S8WuCC0+kk6ZXNsYRopYTEspUrFtF5UvoJLc+K3m7JeMULkwkv1VH
poq/r3DrdJZU0oBFOWBin/z5ixGL25cH/v45IETbAYQcRWm+rbK1at9PpkqwxgeQ
zcOrvL8XziA4WHCSV6Xx9TY6qFs/ZGIZmEjAwuKoSB+QiJZqTqFbQ7xS0bqBPg85
KM1v8/zDGTV1kWlfOqHXGpOWYnBSzJjTtgh9d9CdST2AvsNI979Tr4VE8GdBup5c
VApigyPD//k3MGaMKYW9c9fYHRUz7M1yLHbRLVir6tnJobkbDcLFi1xT8H87JTx8
iRQ2zSE+7Bpv2o2F/Pq4Xsdr+Xx9qZmdQluJyGVoLrByj8fIqH+8JemDFkYN4Un7
BRtKjP8skLEbL2bClTyMnPzB0upZwbirhZScQBlUJhU+hU5P55UGI78oXEKxXFs/
WkYmWNw4An3/3Y1HqYzafXbXDl48KAMA+uUx9aQ1hsFgHqtfBpiixytSTiupI7La
+2HDZWj2We643eTS/pIuByZVpxP2bDE4qUeraj5057imafynaB6fYr4Rn3wvOIkD
vDL3wsInkbJq6SNz6QOAkqejgkb1ik2c/vM5rV9Ih6n7Vch+hIhlmIxlx/JK1I2p
k7NRO+Uly52TQABFHjNNS4gBJFB3StNMwZlwej2Mk0NGwF4EDFM6ubZ3Y5ZQAKbC
cDptgrYJD0x8hYaXw4Cta6Kg8nXfdAIxHFHllflEgBi+dFejZz+xb2IUmfvpg6J6
c+v+Y5NjA3qDh1zVwcp3Nh81i8JKilpRDdU0rAQscyV1JNa8nOO/EgmlIiW3OoFI
TicivIsKqZ1mzi9VwvTU5WsmN9PwAE0AjL0ypP37Vf5d5eE320MKOj6+yyY9/MFy
Ns/OcoiRTMI8sZsU4/oRFMuy/UFbeb6YkBN+cTzJ9ciwrAAzhvKo3wyou8VcYN0R
hLGN68E1NyFa0du3hsOicQymbBd4sfrp7iQ14DPWDtjPns2r4ANgjicbdo5SNHEW
PLvxxt7RZNoYVlZvT1SDSo7UUtZyg0qRALomJZYJOtpsmOzXXG7xSC9iHerwKZ4n
esmOspr8QGbN/beEBblM18+x+3vlQhL2hDXBqlgZfZpi1deBZXm5AYKdDwC99y5L
aZYsTyaLPxG34RqyAqifIWGhNb0IKA0PJSKVCrGwwsk10qkSJYhCIifoRzUu/be2
Tho8PGHkA48qaawquAOmd/hmiONfNSd78quCWRdcvVIyaVstX8jDYBCLDtayRgi2
eZxHFzePHfGoULjJdcdyJcucK7Cj5F45ubNfkrJVVMIlWRbBXnpe6kUAW064zgHH
KCSiCGbKoHuAfzE17qJE6dmyoyGZRKaNNEmJr2/V3gjxPe/Xu8PaEz1hDA8Rujpn
q2vAtZgDkrrnMfJoz8jLnJyT7MqB1KXw1/6cqYqbdIwau8dH5aDL7ITkC+bCe9c7
W974G+YDlVSYceq+ttpCoHgdvzzeVLCawCTFw9IDAFluDUl/E6pUMSq+mmU8Ku6A
I/0+HoXoLy0OTnouMoMbqxJeg7M3ugKkR9Gc08nJjXtbVjjOMRta7l5lJt/BcxcE
uQ+dsfRRQ7kuK6WXVZkHflP3pnXabRCeJJmg/u6L4U4za9m5Y7AScOJQFyCDqGU9
nekdTVsEbgDyAYLExsB3hqGe3z+SwzC5W3vFoOATQzZBcGcMetgJnYQMx9u4E4Hb
/+VoWv3l3zlofxngcJw2kYQhSpzA5j3hk6JhPviFtHIgD4u+8EEX/sPpQ+NtM8rp
U1o2hE+Guqznh9DaTjMOOmFcqDNK8UBtUf59y+b3B/2J9Twaul3WKzaCYdbb37js
MhzuWb8OGxd2spWvyQE/qUFFJGMLW78w1DlcYL6I6LFPwpTRGrsPH68qm2FYh6Bz
kbquRBa+JIkLPZjBx3JuUjCfSCNQ+2IPxeHIqxlE13m1DIs5peIzwE/gv4USzQw3
j70vck3BPFm0P45rV5EZOt86ENZzwuWnlhHBxaS2Vk7nlIqhJZukLYVcHllh4ANM
xQLHCaFiUwd1uelQyx67HZsVYXAm5PBHiVC87CF14G+DHz0AYG3nIrRdzOdIg84/
D0tigcIyZRTKfyBF+6BRH/Ro3+1pC/LatOcS49LHNJU1GLl5FVBzeMKZ4NLo+PN1
Fik8LxhyCOlOm7JTJpDZT64SnSaktRMKvga/0bniyFnEz5bRlhnLyUysf9HZMmSX
VhuDdSvBLGtluHBByLkO+2YJa++cD39lQGE0NdKRxddpgJYzcGrekZI6rGlvt1bf
SsFMWvD9V1lvDgjQNTZulHJqJPJ2h2FneMYCUzugUsBpdg2R7AKtMinukKm3APVL
Z/vTo3UEbJJI9JxLqgLsK1ES3+7kUJP1XS8xMwVvDKLQLT9yNq+0f27xmxJHlsRp
nitF27uVwYjWb+c1b2hsO9zrYcnVmtvCvANKnjU/PJzKzjbveq/lpZu5wpacCPlB
KIlL6LmXLSQxT1wUkzbg6MtVjXxK3vXKENZshpAbKPar1o5VkkCWFMqXHmnQd++N
NRPUK3JvoVmqinAuIEFY8E6rfOo/fMSLwfs8YGHllv6ntZ8s+mPIfvxE0Gmworp+
N+9pvkc0pqdgFD+FO4x6CxWE420q322KNGOC5FqQJCH7LjnzCjZYuXK9AqNBwQFI
gzwKwLrva5zJQEDJ9PNSLkj/IEEhRYZhROQ04BXR3SMhZNayj0WKEEAjUMFajbZ4
ujxiQt3bo2VozawQ6FDWe1VZfCmwIp21uMT3b5A7JqNxOqtsTs+EkdOkQ+fv0/3h
407wN789EkCBMIvo/TZHq1r/M775j/mxnrRGTau+GOGCxBu2U29Ij3PGak6QOPC7
WD78Ft4n9zZJVFx2MQOrf8wCY2LxRXKoLYhx6XmpM9nAwTvhVJUXM43XJYjMwjWo
OkJSYk1GL3epX3GDNGNaiGwbhfzbrONdU82HC9Y+jFwDv2gZfQCfQ6pO2piaWDpR
MCoOKtvd6lBv+Y+SMX94YIjpffrsk+2yq/wzjTIeit0yiCDjnusDs7ogf91PUKIh
cg3aSN2Ap7vLXAFtfEXQG5xYL/x5vxaszsxN6pWNv5+UpxgFJ2EVIReAxmSDh/Fr
ROoovaJ5m4L92yrFTcHesQ/ugFGPdOUEzVTuqNQsgpLfqrRKU5c3qbVrgBUFgY/1
AR3/BrxoPsGTyIfhPLz15vgKtKUnfaGbRcYkKOolUTj8ceYWs+1GnDhNKqjgW2Ki
ap5cKYbhhKbmAPLNEF6tl1xhAKLGUepE1GuIFhjMl8VqEIPOzMjOllSB/OWHNSWJ
Mo2iQJ58EhFeT1uUK9myfhdAataMIRExuooTaMKe/Fpv46ZNCqwYTeecogupKIVW
YdDXSZuiqpAeMvzhtlnCddoLV785nH4eN+C6IdmZ8yi7qTTxx9KRx/OsMpWljwOU
b2f+BHpAJdZE+rtaI2HDmtFrPj+YlZPghUephIyPKMrmF42BFyjoudbY2QMnBsCx
RsiqF/O1OOTyEdMXQhp9YeuyBPyz8Ix4Bw7xg1phrOEIfUAXiZy7DZvTUsiTu7xq
s9JvR+tLoi52opJe2IHxNpltc9roSiAd7W3JA5W8iHLth985o63vaEI6sd3CarkB
tve1Dntl0qPFBY138UuyjOO1Sb7XJttyVfHIV8m+vi1uY5nHxT/gI74RdYnLuyT6
bb9phvfrRxEXl/fqJs69RQ9ftR5aQfS736XJnDnLOMZrcWAMOMuayF7npHK7zPC3
EuBtv6UstBRXsqmvBwtTIkNvIsBkq5Sax/gg4DYOMQZzEJcXBM6V9aTjIXcHcV60
5lLVbKfzRhKs0rmG3ITgqL9j2DAYmG7c4lViATL3li42fdbP5ph0Tt9HQ9tppaYU
cW3sWcrlvPMyMMtD9qrvntO4dZG+myVhfV7ru7moIXPVbrqA8/WsLPC2OXM4s8lx
cXnJdFs6L2g5b67QOViYLGWLBOSBJVENExS6L09iOiLRR/n9IH10ERlfqkz/qKLD
kFpqH9gzfOgP3VN4v2uHpnBk/kVNyRCxxJIixs5ZhU7fsfI2biLaIBnwUmPsUfwJ
6Tr31ZA9QFuJKuZCX1KvgJNAaE0qsojK9tmKzWxse9yxsfnW/XVp5EMutPormOiq
GF/vvyXRhzxrHrSxq2VcWQOuAmi9wTDh68/yWFZIrOQoHGMSrtoFNz9UU4qj9iTm
IinVUXWZdoyn33LarIK0BN6A7p//WH8Ug1jXm2WBf5dTDZi4jLxZ8e3138WHXolc
YfTNgjYqREQ/IuwzhddoeJzFvJ+JupIu/S8TVnyCPtNp2IXdNc5PKptEo7dH5cOg
c+eBgtntghFMypQopwP0XjBL5H3n1uGtfCukT1ZNLrzTVpeAqOo8CLF+RTzJYIAx
U7c/PkU8fpJjN8BviOt4cOP+wb+v75npTk4d5qwunFLib4x4kkp/hnE1Fk7pgvEF
/ouXCdev9xzpT4qZBE3VwV3e4omnNNGIfPYYS1dbfaa+V15Bk6gPlxhsTRVWotBZ
51+xdpunl1MhQHXI3yu0qEkvhsWpAg+p4qLttLPyzW5xQALo2urmtAoZ9YMRShkk
iWnIbrPp4Oqhd9p0/8Ih4Jv5JS30zsPZYuXB+Cik0jdIrnY42aot1BR9ZoxcqjRl
ZWKGXK+97CJFGTGLfgzOFs+jnhEK53BH1yz8ixwVJqNKQ2xvd1VhQS6nnk/YOoqz
ZTu2oRmOtVcjsS5Pdhm6PClR/yGZAmSkGItTMutEu/70tqX+iqtEbniEe25ApgIK
sOMKvOEYSQrYdsc/0+dMJ7Pg5Y6X8KSOaATY2524K4c8uvXLKphcNq86W+alaENq
gGA9PjbHvW+B2bXfRZKVgBwa8qg2wx3Cn1LDBie3E2/zHSVEY64LLdbbDjfVR1dQ
HTIRQExr8C/GQgtuQCv8+NqP2T1VxhngrmgPqWpw2dYNy8yKws0V8Hy5diX737UX
eYAsJHvMB2W5bQXkwmDKvLS/Vu4cyHieMRvMnHSqykyxRU7IwrnELtGrN4rtQwCc
Vg7zNcntWiQc2pVNiKLjMY3rufsjKiMXaqvOKrl3QK8CitmEZxTIpjIldPpji+Ub
m/qq/CtuQTJaKydJVIm+LwdRIOjZp8+U2RgodV28Frwj/uAtZXzursfUEJc71Hjl
h0QiAyLox7PQ3p/4xkn1ozIeNbtXnuc1LMLKx0tsqyyxclS9nGL071Fdo0Lq1xjl
CYFnSQEP/RjPBnVHN3xo+FUAs0DCA4qRtE9AD0POFvVfCk5csiEFn2GM8EEK5Ci/
LPwqSILmF1SNwv0NIdy8ofaOc9rSgxtVAcnKM71/gCx+/CxXmeWeG31zzcJYKxiJ
31nM/WwPdz0oygyFxYlX7WyowHOv6LIyhdhF8xjgnH+6E+7BSGopV6M2ePtM8kFq
q7yEkQwms3UwL53YPI5QQbCuribmCSY9aYS79iz8ppFHrItJC4dUq0RxLPEH4TSW
GfDa5KUdID1zUWcPf/ns33TbN0Ei5CveGCRQMZVoo/8K/gK6JrbcskhZlaZfBAUw
AG6DHIkhDdTF6vYGnelHDU2pJL0KJgXBGakc0fYLf+GXYj4DWy5y8sBB/KD9daLi
FKpAZo/E3PYzQHJttZKmUc97Xhql1q2vlj+/KHEhTlds1Ly6jxNGZ+f7ChpumJ+l
5hmvYWLXg/zZghd6VmtXIwInByrgNa90Brzip8IsIv8/FX6S2ZtOkJD/Qio9w1I+
fde8j9ycvnJcBokeB6g5GWeM9y76VvUlRNY9jabK7SLiiGfQalZ3fKBd1iBvjgJj
AX7ZLCFF4edEISZpRuWSrMhJT1TITjH1Dsx/11U2jYx50UuVdrBdemKnwIrhJ5o3
NdlXXWiPxxAxRimMQLUqbJpviUj8SaTzjAJL1R6MlpH4H9rUdJ+pyoqKAUp3m+zw
uROHxCPm/zaH/0C6HZAutNEsMEu2Ym3ukU1UsvAAjliTMN6/VQG3AydeQ8mUSuQ/
s53cLwmzW7iK4+0MKH79u29cmaOQbP31hFKcACLaod0i1WV5zXJfqRHQGYCHzcRZ
5eqxFkT9QLhJsrXvyduiRLksHcviw/lUJvr0HdQk/GPh2W8Ffc5hc8jFaeQCBq3O
n45nhSqFG+SEMdscIrR98GBuHWYJJD2npMe0okTre/WZFZ+U9W9HN8zffa+Wz2lC
rrHLOEU0vQPhn/Dofs4ilraIZ5H2tfAPyazxAwueZ4jvPaSTrJvAQ/krlswuibup
I3FaDTuJcfqbPUEE8WLZpxPOli7CcsPrLNIA7wXDNbMn/nWlUgV/7E+J95LAVMyJ
5y415FDzp7VIEzQvUEyDge4+jRRkZsoN/E4GIcihMcJVSsQwmC9up7fucUiL97Wj
qeDGzlGdem7Oy3fMN1VpuvEbeyxrfXmt3gs0lEtiZQHp1GY7bQ1uAdEINF67eBrw
HB8t4Nyy9BXaTQ0uujdLzFvoBbRCgClvTM3CR7knAM0twMwzh82OXELau7aYtrvx
El53Cs/2Y3gTQ0wCP67f/DfyIrfxkGsTe+Kmdk1EudVDV9OikapRb9Oms4ejXJyJ
rL9yY9EvvfXZZ+PsI8FGYsQsRl8UCyyfbMO/fzMqN6MLLPftFuIYLuS6LcvQ7j7g
xpqbtNjcR937azKddVBy6oJ6eQfHosQ76iWo8dFr3pxU8o5mbZmll7ATen6JVhZv
lb6W1GSNrvSD5VK6658J5I7P18tHzl5FxwwsRwd8l9WQsKAw9YUO11nUmTgEhEcJ
0ghTq86HqZ7EkD417AgzxnUIpqZPBKTsM3LJJZYhESqZXmX1jNUXV+6PR7beaRhf
1p56+Hv/yzbIVwqujUJSZQC6Kcq7rtQTyGRyd8HNFR+RGh1zAv5riZFotI0bSVe9
bL2J8bVTo/D4pJ2XGJjQdDTD8pw6bzCkEMUNzCFM6LL9GF79owYrLNhA5u6iozPG
rTBEqiy6I5gAdoCb/s3dk/ASK/jVq3FpbUgTQcVdU6Tn3kfeeyf529ys4CGavRwx
8Au5GtSStALM6T0IRX2Cyi0W0BgkEFyyjldks/tKvx7wRN/25CJrq2027PfwNxK8
L4BjiSVVrSPLIoeCBn4i0v1dQwYGW/PUhux39byr/kSwYrPk7L31MI/RkE1D/y6A
HY2RomHkAa3VZZCRmdvLDSeHQO7qWXoCw5ukKmB0nW3ryudkMxiXRrO7fUaIv1o0
39LTNBLRqCQicg+zui8wtrUY91VLX8A2W/GcvXNBZsT5O0Q5fLWLVsafrQmIolxI
Jh/TZHh/H/pS9LCtYbaDGflST8CDyLD/QPK6XMoSDD/yyCtA/agUKq0ki9dmk5Qy
Fttgc3xNSoFOiaOGvN6RFYbPNKeOTM49cuk1qyqzzazabJHsMvHczqChk8bRkNI/
0Z1qR8YUQ621JD8VNxyc+hCYptwQEAhp7CzvCObgYEpJ/oYv3gOuK27940x/jDJE
0fsASVnaeLb2cf3yMaPi7ZnN2xyuHpnffEIypH/4ctRTSKu9VapywmSoG6YwBFiH
8Hl5MgG256P63mJiBMrprasSu0MtTsuLwpvmQdwD8PR3fxLz+Y8X1AkA+D609R7c
riiJ2sxg5T7BBQSsMRlWlNgiDvrXuI6412BjvMyxfHj3CtriXq1uUz3W7rhqfsQl
GW3BKCu8ue32xA4eFsr8xAHxy72AKJC/2pIK83GKvR6Q0RkT8mul7xEHXlcQ3Qat
XE2yDeQTIphwIfbDkdoXfbFHnDs6uwtLxi3qgqh+asnP+VoeCXGlnocJq5/yX/O2
bmA7SoCrOO714tm8GQ/7DpVz1OMUnXKswOjoE0dIMcOhTGZP6bvi5jwPWGaVzd0J
0L/lO/dHxp9dYL3WNzn7sadSf5EkztUvSAzJqoeJ6kWGZX+00oGwrXSopnCEXOqx
+3JkPPLgWK+vrs4SVt5y7O/R4D9Fg671L5ZiIDC6A4B0BdcaMVIor20YXYDcEDQy
Bi1JIsIP1ifSToc7q51ht0Ni0qsubTDPnfWnTEe72I6ywK2BGqEwKFf6SvGNMATs
zSlyizfk26TwV53AE+m+CHuMGfS6ybPjrOoaclndLQXbSxqyER3tg7HH6GdLW/Ft
1VrLnPwv9ZDnOolMEYB4rhE3UBmhF8HsPym//KFxAx+OIG7tJni0SWNEv/u8t5Fh
TTMzx2F2FkU7cncP+yaBaNq5BdHvPwpe8hSYiYMgUwkHBKwRWQfJrzTD3m+9KtYr
0hMBSVmpA217YaBq0ykn6sDjI4MlyOjH4C/Dvl1gZOz93FAu6lzRRnzY1DsUgT3R
ZumucKIA29w1MMD+JsbXI+cXUB/7FwCYUFr09ctdz5HsuniotTugVK1rxskQygMO
A/JsKQQEU0ZWbISSiwfiT47FXEgT+1ooXYxwk0urEdItlWSH82hO8gt2hIrgD7nl
4Xc6PiPY4uYO0Pn5FoUNeUZZR9dsAFaHQbuDIx7gm7rsonDongtBuxUngxyrEAPK
5iPx4X9jEz+f4u3VCBo/mcUvxfLJuF9Cn+oXINv/CqIfOIY2CsKEaSGOd2qTY4OE
tLrhRetE8upf0TfNnWFWqzALMw2U5YPB6IJtb2wYhcO6B/gzR0AZvLVDoUC0NOOi
XMVLyGMnAKFBvFrwkPEfkM1GjYunTbYsBELa0jQB/7fUM4mbUj2kJ7CJetR2YEv7
7pt90UjjhA9n8dfqTwkdr16J0a5hpZRyij0T/bk8XtA6x1AaHbAob7yI28wHgIvv
HCqg63vVHVARJ2hrrTVeSDYf/DhQukQPDylLCZnpCD7UUaXH4ClKyEA6SpOQM82j
9y0sNdopke/FdJ1Gmq2iYYJn5bKm8W9ZyTRcv2QK+Tq08GhGYDaAVFV4wb/JPwt2
UA017drZCXrBb8JfmfsHBeFHOIE6Gq0XhsAb59UDYCuOT1V7H2yK1T+mchkGB1rk
pPGSObLc9OjRhje8n22MPLPil248SrEfb8nL+y8fpyHUPNqaAfTMudGm+T+Kxu22
XPSdFpXOmd6PovOm4rRzfxdOCJ6D/J+qWGZw2a5lhkELEopkjgJzxVJeJvntuz0K
HFueXZnN5Bni0QJH24D7ViYDh9aP3HeuWGFGaRAJ9TlCZaAv4zsLYdH56RfwWw2n
rfkqSgXv2GA17XJfyvW6eR3X4fwqvrBlh02FqrkX3cFkAUmjm4u2s3OXapPfmi7Q
7eR5Fqgn0wkwerDQjDjpGMxHly1Oa4xboIxZqAxiFUXLFVrj3Yf0rkvi3GySyeFj
cf3KY8wGQ7lCSXN+HnYY+CgcIr/aytWvzgQuNXaGLJTQyyZV40JJ9ek2oAogOHWI
FoQJT/BcnIbijoXpvXQ/1FtYhr/SmUS/tj9ndGD9XQ9mfbmpF2A/HizdJnjKtWIA
yO3eBUM+SXhHhYyT6dN2cFrG7RGVY//L28neWzJrk0VgG9fiIeSZT+9VkNAe2rIK
SDogDCSlNh6/n/FtPHd4YihiKetumVPDt7H5heSlyxrlONxlm5CKvWsTxoCMBfK3
Hq/hANRPwIUiJUZivz4H3IMV7D04CEQtruPKgkMfWbU0//IiD/tMiQvtdErgNWAJ
lRksaGLlmvyMiSAop9q+64OKskr0cgKM8obPf2FoFtLLa5MWNVfLUFboNE1vaqDd
7aMl13bmmfB/oUbRWosahhJH8/QjKYGFIFvqVCgYP5wo33CQfx6Zvbzenx//+76I
Uhqx3YT6GTMSm7EnisCF7EutLCmykjQhyfxRAOVkkTL66HeZZG3KhaonPtLfll/m
O+9sNFpU2jgQubx3BbfM5OBARGMUYkHphZUccdd05/NCf7C/6QldXQ2tQKkZr3Z3
oEaPXkD/8HeL6TrEfwMjjtOOFqRCnDI1XTtWK4/nztV36W0ezBR7p81JjD7nq9gL
l4us4pOwzYQ8kZXZSHwIeEkuQuck/quYFTutsnax0Vi0khI+DQSjagiHbsW4qUTL
iBQtmsQc18DYiJ7+vfkTZ7Zj+9edZb/kx7SY5D9XT+7I39JqGr+2lRSqGV8Baezr
5IudAl9YY5crLuZr7RVx3wXQWWhxl+uzozdP78NvK+FhPtk5Zd5Q9Op3vOeG20QW
DDGAUZL/KMjwpBGbYhXdCpzTUc/YsnOgGk9P/hIjubbLokM9t9DNA2Plww2pUQtc
Y0p2SpuQIUVIQeWo0kq2sGzd0mVO2qU5pTna6LOv3Hq36iD+GlqsRCiT2lkBwGP3
/WmWQzLlQkgI2DP8YLdiUZBNEquoR7pKrYLiiDBizcswPltwFjGlYBjGRZ6bpch4
Thpg2kcqsJu4mKkzTK0Q3asPCK7trSEeOako/nlwrwgMN93Z7cnTmZgaK6cIk8dd
Vibt4Sf2gLA/b1wyn772f9/yKSwUkUx220sf1jmS22fcUnlWQSwq6IQgybqIasys
+k4bjnuH0c9EfoN4xbtwF5mp+nRLsBS+oU+tQWrBdr2wlN6IjsNNkkOmvQe13laQ
1YBHmCY8hdJdspU4ZBEX31yr4fuu2hbF+syGtQ2jtx+ggZ+CtZAD+YwOnF1q+ZMY
+sckO1BmvXkJrRxoYaK6veKvkGfBS+JDgiPfp5DKlBHmhBUJunbuZ0dcrq915+lH
hIwb7kGIgQKw3RWuOM9aQIxn4rdGnJVslbinHgWmhTxvGqaiWRZB5TPjRIERYI6Z
LRBdP6FoulSbgmrb1jmP46/HixR3tBJYAdA2y3jL5gphwrCxpG/AQ63qtZC9/616
biKtY3UmixgxrEgjdsIIr0hZwOfyDr/j2MPjeIbFYpbQy94pvVvkfhAQp0nEEMWf
lJZLb491TwWR8xzazWGAOUt2qJ4nI/GAEJVVKxD9FncLDYDh+YHUO9WNcmwMJ8Jg
ehzD+oSNZNJj48Uk+NZ+R7LXjF4RZQg7wISALw1u5IZpBUAfWn8yRrteOAezke5M
3WNAFuqXM+tzmDsKoBznkxl17RUV5xSIIQ9slVm82rEjHSI9b62lTmiJpRqT63Gr
ZO+KGS4szMEpu85B24XugkeOyV+nmZOm0++/Z9mTa/NAsEDvDPFuUVwb5YAhdRod
GaxjVE4CfAuWWHmRbb/13WwAcIQBgkIiWLyCk3+3gqOiCmwjf4cL4WTOzfUdtI3G
8hTpF2GqIx3k0W5JG44JzqUs9Bwwz6tVbWhgwQFXUEVl1HRH3lJwrn7AGv9BNPmT
0qSyLmduIK2TXJ+QDzFP769NGR4AGjRlcNrbyvjYeDZ9Ozx2HmVXg4YKwjJM7OeS
mqM45SecSuUUEuWU67eK+6Gigb9h04by9/yls23sAu/iLp8KohYU/cNYuIv2Ric1
AtyAYDG3xY4c28neapXeNLOpfFYKh+3IfVsu/QiwH/6JU4HE3nC4yp6NqucqT1KO
kUDAntWgccklgN7vHDUoxVE0gU/ZsxPYJz9r9hgonK/bfe4KeFymajNNKZh8ishE
Vm8q9Qf1UhdT4l4mA+qAErT0oCcUxBDm7GIie31xHtYdsSAFpLXiffMks4wbN0OQ
arAwT0YxgICf2RvEgjVZeVK3bJx5zxTlzPIzNk2NSnNpWl1XdKyD9p5g0X/0toXx
gi85JXf0oDCuR5gj3EWc0yINYFMtUBe/XOfjftRZ7YNunbCUO1epgLOT429+eGAK
kvOvLpdZS3AYRfNtWq/EWf/6T27tpfdB5IMeOBBJ44WWqNFhJOhnvlOgDDiM8FWV
1D5ZnuImA2K3itj9m902+dGeont39EcYz0180GdVbd3oC2Az7pRX2gcurqDwjNKr
qBVpEP8BAxzxUVxsRrhJP0sOTbtv72x/+4WcFO/sK+amh+wQLZhCdyogVfkw6TsZ
RcDAePkjxz3vP6QEkDgCCTqeZeQD/PaWFXNafsKfJSxCXjUgTxUshN/JjURaI59e
AfJNX4/HPbzXlOVTB3awXkqbRemv+0oOT/j19nG4BP/nq+dRcQpktq3DRun46TLe
PY1WRrZ38oHyPAsrR2MTeIJEC23njeI+j/pPCP+9MZ32NBaEiX5pj8lwVWIcUdCS
GdxMr5W23eonJxo3/itWN8qIzcUgzVwbkljPz4LOtpKbLU+DBDtEfvv4up3gjjDd
x3SY7jOSnsRoBHDlRK/grkeQ2SF8/wNNQUExxTBXpE9VKkjy8Z3AOzlFMDeHAHpH
MgqHKeH7dPDUP0YJc6lrSjvJoG1RFB2OIhvxNHq2AuBWkErhf5IUGvvKr8SiAjHg
qrC6czuepZgVMwcBgQFwjhAv9XsmcJs3Acmus/kmZM/ljAI1eIqgzHeRHLDGoeno
8liD1VWkAxa5c6+7BeRmsstw2EpnhLDGRXmoNHOaVSYTxHoWiP4xkWhWYgtnPXEr
mQDfyxYIVI3Xtg8rt0RVQoD6y8xJuUgTA3jBrTh7wlQqMMI/jXmNcuwxjmsFQ3WO
Y2Pii4sRnxKaUWoFAMQJqGxvlJptbu+PLUOcVsY5dw4HpwKU7i8xFBCAedehCZ2k
bBPl7db6E5VsN/BPqBjiY3jpaGUHj9b73tqv8qR96kC+oqvXajm0/vNebg8DYDg1
u9PV65CgCTnyQlpDGI6TeNPw9LLvt6VS9rjdTsuz8XaRH4SvGzjikCDKt6yplVUc
mTT5h8WPz7X72mQfMT5YX0it8j7lwM6X8HX8uOZ+17tAfUAvr9HLWqGvLW7LCbac
5ir0GdlDl9OaTianhVtgaEq3L6496jmMRtVbi90eJg9IoARr1pmos3iaBoHB0vcE
wKLnnpaEGEWlE4mJZGWkFrBQ26CE4cQFtnvOUw85cvFBJGBnVU/WCBjDBuDY9P86
QgM/u236Bx/cKJBTm2aA//up6bxCFJoMEZ6PAeCsfPP7sEajwUYkIfuG8Er/yZBS
9ZoW14F17LYSYYsJJ8bPGTtiVLjpNO2SL/YpYSJCN437TcW2df0L0HIO1UGOXiHE
H9gdfhhCS8TtNuydSAF1RGdY0QgWEe55Jir3/0MTOmfRwtPHXYhEnfzvI/h1Q7wC
DmfSV/9RY5GNBmQv0SZhGVhl+FSsSHKRb+VTIVTIhn24ARJexLVF0ayb/ziPkU44
CCK2XnzWEjvm1jptJq4SyYgAKFOp0l4YUJSIm9BS0gAVOdA9m/y/D0XyYfr9pZ6I
4EvN7NmbEJaJmNQ+mT2pWdsMQOJ3if3KNsD7+aM5WpK3MWtKCMFCJ65jPRWUIdtj
03E4Y6WNneoXVALoTBs5uiX3Qe9sjm+brdokRLD7lROp6Wn4btS2BHUHDgkmz0uw
P2rwyEZ8/7r8Vb5rAuU/PmZUJZcKz1yMrCHoXGYeryT9qRKZMuxw4Yor20pwXlky
BDxF3EFHHwU/QIZHGmXqShwBfQlrm+C/2+lOHHpIu0/TdQg8ImmUvKT8eDwKfwHx
cTn/L8Am8VGsOFn1Izu0CrCGyDD6rdfqXMmYnNOZKUnLDiUQL4kdw2cQwefBjn0G
NjuUcmI+fjA3H3Vj2JkBga4hIKXAIiAMzjj6Q//Ry0x2eEBm9XNG6TO9uZY+BPiZ
jodaQVcDSR3XeZYLLU0DOjunsnBpnf5zvGeQtHAn+S0CVO0vxG7/gVdLAYjbZaGx
AHGmiYX+GgoGbQk5Fnoxav/9HPv0i+38SreG0CtI4dziUKG5FaRLaHwy/5dWbKqf
OOojbrNEnfEMRPTlth576qnaARxEPHlzA3XNF2Hv8L0fcjFR1qPjmJNtQKE7COl+
x6sIPfx3/2rLIOTArROLqi9p0kwynkjTu0JVTcp0/8D1Owhs4OZEf/SGRB/ITiBe
libcAnWgCvMiGu1aRrF9nRVaFyVlnVjWzGDE1PUpGz7ajnU0m3+ex7UcLp75iXtp
Szj9RlkHY+0oxdPG5wE2LRVYzFabdXGj2SZWWrtoVnoDYX6xeZd/s/eQX6hWmmB1
Z5iQz75i+tsf7/dlM8bTurtJFDtO5LHEstw5qm2a25K9gtEf4MzvNY71EP6oifar
O8Y03GT1oY7Epxrp6ueWjJk5SntQzXUrIH/FVOvqBFRPmxMsL2tGQBDwC10h++cR
CGzY8gN9VuXfFc+QWNtRr0ZngaTg2GJx75FMqMKPQYhDV5HrV2yS3UEkS5jzIBNc
4usWzdcRrZ0YQNtHA26LQZvJvgROHus8qTZPWEabn/NE7Pb7ylvpanGl8KQy55F/
xCC8c+0QiBeKg2X0IjeWbdjGN7y2R5Dmk1idNgrq8EkGwG/JOX7mTlzuzFQAcZFX
73+mnSa/vrnW4xtKYmTJo/FTnLKTFd7pEWyyXne7rM/sBhCstsSc3dvyeG9JNOcw
N61cCqE6ZStg+Z4BH/R7h5Wf4nRw+w5AbWiHusAEcfNvgwtPLOkVVU4YD6lHaXJx
D3EKHsIBV1h5T9kYPrthIcNsuO45GeMcwraBoxZs5Lvw6dhgehvGk39Ec1So3Mpx
RQK0JrEW1bjIkFKVpu22vm9pnSLT7R038iWteSXQq8Xp/AK8cdwWbAwLTliKoDmp
qButrg66bKA5dAGYi/ycO8U02CTuEfEvPnwTLeLgzu1J1BXJOo8gnucHOM4ckjxZ
Mkw3opkHxU42DoSXTeOV33ZWkgqyasAitDyIbxzrPn8zoo0hfTM8Iw4QQZvEoj1S
jllTYBHxt0M4cprlmziVxG4cotJU+Qxq9Qe3BUYDviLs/FoyfxxDBHzg5wKelDem
3lh2SfCpl7YRiqjbdxMl3B0GW2l0Q6VFyBNUg0l+y/xlK2pgiG4/83GPfDvbLbzi
xbORa3Ftq2K2ImWIKvXZ25FDza4Dd9iKXsw7HDr3icHHAFD0Dg44AVXBOel5mF/r
1fYceixOE233w9osdgsn+2U70H+dIQGUhH53lu2I4JW6SMGp8hHwArn9BR8+zyI/
X1TgcIKEbckeiyx9Xe/rD+aTtwKnF4Cl4wp2M9KbZay8hbmouuoX7ODwvh0trIE4
Gn5Yub9imtFyJ+pMIIbVFA0/5B6QtwgrsLnfH1eL90jCHEkIRNADAlxK/zmmOjCS
vg8UqZDX4S/QDqifOS936lTacjInFh2bavK+V4NE+K28Ahb3b4o00N7NbC1nPnnf
W6J8jKaIrfXqa6Qn9YB6Ce6Q10wOwodRxB7NS0fmYG8NwqrNdDoF4771NF8bicp6
8LioQB1FbTT/T9RgIaCp3FBY+CfPICj8OLIDj7XpXQ+xZCbJ7IAXJ6t5ZZB/gIfz
DsAMiUuvNwzy8Q3P9GB0GqflwDoDxbgMG8TrJ57/akjf4Z8UWkLk9GpsQDnmylj+
3t8ee2wGJFeVfWaDLbeXM49+KgG7/DW6jXxYYGBHHqn2zhXBXJib5RpkOKyhed18
od4Ij1uDnjL2ZytgJF2MKmm68VO3rPzTP33qfMuXKj65fxmuSrv8vaai8WjDS92W
Ny3ISsC5MSYVIe2r2qXlIkaso8bPq02622blX4kBZZ5Hg/KVgFXLPJcznFzQzEVb
vEbS/gdXcqzfjM6AooxBd1bAxIeN7J0eptKB+1iHDz7E+0I1zcOjjemBkQQQR7Z2
eJnhJ4t2HTSSv/WI4umo9VPkxECszSj1o7nRTh/O5VXxfcBDmvJmJbF70CpHY9Be
NJOADewHYVwscyPuWIZ5C0S6i+laLxg+zP1ubKXnDbIzwu9V5IZA1XSL807RBHbm
/I1/wOF0i3ZQ6B74MLHaI1I8m/TVrAF84Tp3g9jTgaf6do83cFtGh2/4zSDNA5/R
7loJvlLlD1C/Hfp6HAaRBadSnDB+oUO+Cx8Ua7xjWV9KnopbmiaO0kFC8UvaFTYQ
02Vr9jL43hius0n1Lvto2cI0809Jca1boDMHjnLbIKufyJSNV41+kDW16Mn1Jo63
D0VmIrhy70QzneG+L/VeP7X4ytXkSGM0vFt7QI6xDXNP4Wk3xlokCQYfFaOwhsNc
7l5kaqLKKl27NwdBIy3gfVq0D2th0exc6hL1xLlstjCzijokDvzqPaa2JvHlrBY2
zHEvYbt0U/vqNr61hf8J70BcW72RIfTW7UtQOn8GhALqU0lvsrYjcZg57hNdNSDj
3O1pE/qrfqXiwRnwPN0Q1kiCugkymgDbh4wlf02xFmULcOdIpkBjZPwrKnT2AoDa
B4J44Ef1V7ibaMolv/Y84yc+7IBs3zUIlJVA2bi4p/Iqmpx0BTj+TU/YY6tFl28c
/jyShoboZ537qY3oNDyAl3h1P5PWKA8DFl3Lza2IioqCr9hPN2iOOkQZaXi/7plF
XqwNQWVKMxSfLKy9TQQiLvy8mkFFMbDxbmspVgivwJMH72Yv0hdiea0Yk51FneLY
JFXl0zPWfiCOo25i4WaHN4h/d2JkaBzM0HsakkNjau3qneJi5nRIKZArl9VwB3Zz
l4M0a/Ep7h6cfb6qEHOxxRTfN09iPcxHrfZE66twi3YaM3Ggz8Z/emqGHXfyhc6u
YF3iu31XyuAaBPS2vqXcsakJ+vpcrch4hxJ+oMR9q38JNEfg0S/gPj93FFQapuXH
k4Dfxcr+isfoJjAD3AKbkI+9wdWpkDxTuHfWyH2aCuEPeglyO/JdWY6zluo6Oz/W
85rdePU0qAC44mSQ5MQXK8sx5SQXkd4bE0z2iZb4V1HMI9YmZkkC43xmeclaavuD
of93Djv4azOHgfwDUyknWAP4XwIMxWcY3rZNe9hlsYQC4loIS6KJrvPmt+IqQEiR
0R17SOuJrchqoKO2xVADjjCtsdjFlCPfqNZcfq1LVhsqql9ebXnRyaW3iHts7wBu
imJ0sNuMumKK0EH4LhaqQjHPkTdRB/a3eWA4b8MI5v6YwU3/4VG/OS/nDvmUb0Lh
NBjt0YHQ4zq6rqiDN9XVtQRJTROYYgs0vnUXjbNxzd2naAej63VGvIQnXmSN0Ft5
grv9cbYuJA1xrZ98mvi6TYOTNGwChrjz1z+C0yPbUPWZ9kl3izll3tcBER4d4hjo
C4xs5Pxo/R+ewTFGSJvaNMOV7FaFAbgoE0gyxtTQCtWKGmsFohwnnm2pAXd5r+ft
zaQj4gUBPlBSYAKhCMI8wkia4+CRNsnfAUJbdqvqoS8IoWufDjlCl4zpMQ4/MKM3
NruK6QTNMSoVkRc11LyU9wJ9kVbSy4eYZsAmiHTi/9gMi67fq+hr58L9QvbteRn+
6ceYwwYUUYRq/ScuFnT1QnUuNQBKIM4VkDA7Bh6pEYX+tceS4ADT6W7vcCo0MgVa
mCMraYhZK4HAjUpWlgqf4/QMrijFX++MfH9qsRICwki/bYHKwGO7tcKDJDr/bGeA
irQkyQdm1uOwuX01kHlwE6d/mXzk9xy1RMIMpJhE4ennuqhPgEQAsJUfM+tcQ2d9
m/872gdEBqI+RZoPoUkIqDKAXosE+q5mQ+YOkJYsyg/Ds5UVFlIyi41GrvEOHf6L
ykSFH7qaJla81DUs9bsw0x0lOhuB5ct//gJ7OykpgmJD6tbTzvnt8J2FC0wWU5W9
TbRR6HqXTu/cY3uPkAyIv9C3mrTwbRe3alY3/EUf65BzuIshVMjovAqxwQdY/1mC
9bEvmgz40c5LKNwSczvEgNbU10HW7fkvGJk2ZhV3yqQ+sKXhtkJVFSV218STuhIb
0lrrC2qyP1p1nLaiSXxubrYOFk8GgGx4NesvpkYefInRA4Rqwk6nlrLO8w9+h8gm
31LxJaanpaOWDiUMDPT2qcvSjoOrsbYyRJjsWjzbAeh6SqmispcglvLt1JfGi3Lu
q4VQFTiPKDmZyyBDlHIUD4ZQt1OJUgbTQPjUV7SCbFXG0EoORizc/eGmy1in17my
tH8eWTXWTDT9CGYNVkI8jgwHLndCDBBBD3u11aR5CuDRDY0nYa1f3Qr4pqW86cgK
AyaKFNMtTJZkXWogbODONOID0hljUdjOaO+4VtAc97gGCpzM6kdBqgnyevuwHLdy
WrBNaFMfn9Z+a1R5L/kWcz9TUA7ZV83/cfhJjotEWolv84GDfdMQ+QHOiNk9Cm7O
8Boh7sV3LON9J8vacbpIqR/ev+V+BjavXJEEBgsVv1thn3U9JX5I5zuEf+UtlmXT
aeRt6jgOAys0qOWjP64785YngjQk0ZqsnX43B1cymQo2PP+1jCfoBMX/S0et3MEP
9sU9Kpl1dTz3dCAmssaSMF6IyNmzC7ue5UkPIaSpaD6c5qdKyzY/m66qAa3NsAwq
dT0/9nmC5Gou5SzWj1AOGOSnhvb/te2VRwO7EOjp1dMfpbYwHsb/lTIGMZ/miE/2
anbXEb+XOUROT+nsifOL151exd+HpRurOnmmD/yXcnMkEVHBG1ZvZmqK+M9GqQQb
3IYME/q3HeX9ycW48r4nTlOWn55082ZntGlu3dY+tD2Bng6NeiRopv4/FJYIG1D+
Ev+jjX+8kFKapdOt2huewP6L37qJQMac9XrqXLV9B8lzMPDNQxTzJy1vpmphPFqc
NpwuLsIy87ovjhtXYgmYGOkdvz2SYvgBrhqo51+YGR75K1OvIhI5nOnf40ae+a0B
tNR8bHUdoNJLFmrrzJWiP+L3qckxK7wl1irDSLVDd2onl7OzgYCPVJvZkLc0iE5J
L/YhZ4YpFC6Wiqy5dK8bKXyYi0vlBB+d0gwng1akZjNcLUc3zBXcIiVvfBlAQy3T
3YxYLArLPcYfQqIi+6oZFk81us0tueFtKw519MVzjuUkHzqnQ0kNsW9sAb/GKW7L
xSOPbo4uJ46M2rjxokTsam87zDQrP5rpyH21pR2IRqlMKSQVgJhn47WwUT6OPBwI
1LV9UZQobVNb5iV4qXRPx0QoOQ1r7h+d1iKr0QIf61X4ZBAS1DNrTB1m2v7umcl/
AXZvlJxA3t30eroNSHn+V6AAallyM0qX+db68vL+Ztl2lsvxhpdShncTGlq5TbIc
2nIMPt7JZNKfAZLqSMAnYgU002qC5cONTlcDHiDGDUeA3i8CGtQ/VY8S6dvt4vv9
B1CwbOL2CtoIpaEaEZZJs6WiuOIwgi12EbXWIrDLHJFEYdsHdOguvMgWFtErWis/
IhBbMGLIDSQDhwaPx4IVMCJCC1MD5C2kt3G3jXSxVYl6MbmUXY791Su0OrBaXqA8
24jvyqPpPT6zktzx97hs6zCLm9cjFIyh6XZesWWCwZ/ayNPOiblCxuPR7c3e2a8y
1pO1TofzhRIvJ8vB5ij+NACQ4dKxvRFFhXRx6FsJPtP0fDTMoXX16WUaIhZ1LExe
BMWbhcR7Q1GVLJTIauRejNCCLMewty6gTx0d+uy2f77bpPRBMyJGkVN7NASoQAQN
P9TnAPAPaR7ebl0u7+IwuuUdq2GjYeuKORMm1KGiI/iv+pxR3Udx3KnfWO+Mj6LD
Hsle0+sI3lK5bA5VSgBdKfopwSiK8iXZ9TdbU7N/mj0Ah8eUTxR4QFRcHvd1jRxQ
8jkSnKzayEv608rlENaN8YUl0PVIQpqZ0R3EAlp1Kb+Vp05WxG1EwcBnqhETIOji
CI70kceCuPUVuMQwSIFnAWihuB9DAShk+6pRtyKwkSH47+vEUek291wiKdl9j0yJ
iLrEDWOe06vDmaFn4m+efy/XEQXAtsTRAUdairQBepotfbRa2qziRIDIqnczEImn
oLU9Zf6FymTvvoSar/NmJBWZ4nf76XclcR2+qYjLJWUxaC6SUGmt6nhBmpXuRYze
igE6Flb54uMftjwOeZb0qr6P+dp3e9RAAGs+rOeQptL4FVW9LUiUFRpaxOqEHB8p
uhjsH8AsO7ltEotMuY3M4dUWPiBbhYbnLXTww+w5ssWeM3BJlPihRgZ3C/mo4GwT
qRQiC/2nD5fAjq46ywjkkRJspKKSY7BHG1+IogX5Hla2BqDkqM5PQHgtSUA7/L+h
YZNTW/JigaWvtBfM893HY9W8fY3cpYgcxsQ93LpfXYs6W7a4tzWoS6rBTnLlm61H
5Jy1drW4dTtsiOjscXkphl0LGTsM/ZgFZhUQkXnfYXDD3jIf9ZzBW8mlTJRRTxaF
Tl8JG7hEyg/Hl2rndpF7T6Owqnkqbf2yZohs5iKqoCI+0lCo4hqkgqIgAH8sXDv+
YeHiuun7TuD8OUUG90ckBuP9RmPPKwinJk36WFc+KdebByXu54Gg2dby6PoHuu/W
yYV6Rv4TyP1rwo+2Nl5sGCJ8IIAOn2uHIZ4GcbAsATUNMg3RoyZh/gBIy1LMUvv1
EdIX3f66sC540O/+IuOt60pdF7EbThjlZSWfsjk3ZRRWZesuZ9vHb7IK8zh1dzYd
fLEGDYy65tHKDRyn5nrf6U+eZnghpUcVhwFcLoujdGDc2KBA/KnZP8FnOJCPoI6m
qO2A2T6BzpCEULRXn3ALsKaHjPKCIoBjag/0pDQFqp3/6aQiP+ezAjlNkkh35eot
k+13AM/PAWQJJ4PBj5jebO570ucHAALkNewfzH7Guv0KZwBbP37s2STePrAsf1co
1V6P/4yFcwkzEawvzkSueBDbLxd+5cly29TevVVg8x+0sT5sEcDhy3PIsNrg9+rl
dXO6/gQ/JHY1A8Hr6mU/fGy3VhYcZA0wDVw4W61fF4sASOewKVVdCgTdFHU6YLQS
WmpZBNqQMc8GbC1ARz8u7Re7AmyKx1ekXc39oGJ5/PUchGCBTnVfqXn8Kvr8JoJl
B/qTDEgM/V3CLkxkdf+jyW+ZzyItZpFJU6RlsRvcXVYFFSXMKLR7Cagt0f9RtBlN
1o/8UEtdpXLL8S/sIODY/OBCMWL4D13erCfd1pUOsbfCy+lCvQzXno0igApMuFwZ
9ku3mKYoV7H+B2aOska2H9ZSjVIgVOXwbNjH7MTXPHpqQppnJfeD02fMCxrSVWXd
vPya1WV64Iocm1YXu+raoor7rrKlNdXE/31oZQbuRquSisIf6OFxuwVt2hWlTB8e
AzblIlJDpkcrI8G7cZHM56ufNLh7GjRm7YKPULWwjP4mE5112IkwGsG9eJHp2ast
z8w2OPg+OYYHEVpUzJ8T4uX8DMIfuhA6c0KXEnF6TK/1ARaPLQwEZ60k6rBVqgi6
fySkQ5bTwfhWNPWAOiWI6PkyjTZAYD9+ED/Kv1tx4TVwEWuW+r8W71JHCTLpwpGe
C9idKkJmtWi/4U7wPXCvzZ0uroSBj4+y4cwKTfH6xnIYwWZ9pIqmoU90nEf9cL/M
ZVggqxyY44Q1S0uW7LMRhKeoDJO0AKJYzpCLuLvR7Z1q0G0QF4jWeuzsCwG8cBxi
IZMGqD56vLgHCzqPNfnvYX0lexhgZ16ClcXb0Jhr5qkbtA9bAjnri/vANO7nxPis
qy8y7a5vb8ZGatbEeLXt8Scv/vmjM2OnL7PD4XpddFxWNvJOMh1/xiPkYkDjHiEK
Bp9NGVnBTwAqIYI2/Tk4Mh4DctmLWntRh9cBfzBPEJdE5d0Q+lNffaqN3O2Z4XLs
4iXF854qS0Fnxx49BGo8RcDKDexJvdpMuJJTU5sIpnr3LBiynERt0t73Egmc1vEN
a/cKIhEOcvVnxyfiLi6fuss4OebI8wzgMovhuFcKyUXeBXa3ReUZru/A4PO7Tbtv
pM2LBipDwIkdLDv5Lc8JZFwfbORuxRNrETzkglhZWBIzXJOAmjOEOKYxn88lzFrC
rnBLcculIc4iDkGkiUslFbmZ1Dry2qBqi81J3xRZl9ao7lDwILronzMlAnUmq0Y9
vYl5drxx13mest8LU+y3UoOjUHnInr+GbDS5wFwmuxYlAxJCglIPh9szKFzPl43u
dkE0IGXkMMQZpNsCf7chwzkTfm8VqdMAnv+55Zufd87eYEEecCLZGmjKXiN0VT9O
wrV2gIvMdJSggIXYCDFAfL0oMMaTZsci/GSamsXap3zivuIoNBmQ4sXrENJhITTT
VkeC15KvZmr650zfE3MN+UxjIw1ScxVPs9jlKoWL3EZzff/8H0JvUPLZ8EpRb4mV
Hck/66FuxnlF37QGY7D4f9FFxMN/ZO4U25efD0hVQUIzDuB0BvHbTGpFjLTMdMTO
JEaMHopRrmnE3neuDnbt0XmW5BcSkW4iIqeDLTkh3tkllwPe1pprBUjH66+0N5O/
ECyIEEHgqtL+r0jdiNck2baeocW+Et5VxD4YH+SigC4UVA8SCehslh8aD85iayLA
67kJC0qO7089coWhV92fksJPPyNcWCRCUd1t/VE24x3S4PqtwuNiFdbELrIlc5Ih
FDjQf8gxRAi0jBF9lZoS7EEGFeHl4TFGZkkWiDigoz2QJQ7TmZQdDwIomOiZpQk+
vl8Y8VVOKV7NyNqPFD9ZmNf0fnaC3luugVCfPxOrR/g42nFXC0PAAOu2KmFP7Ygw
DaGROqj4beQLrXzQ0cm4HImw5J/YxK7pwGH/p9REatAofQvml7oowqTKAB9ocYds
`protect END_PROTECTED
