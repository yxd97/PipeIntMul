`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
htK34gLuBlxF8AZplZeUaM7RZwbOA+tmckyPvjYg/XRlZgLwNWIHfWcU9wtDSGgT
bUMLm9AxL+wYXCP2KKUYm0W532MRS85t7g7XKOJy4MmD1QlsvPyQO4TwlLCa79/q
q9CpgvzmKqEHvLFd8uDRQ6VCmbCKSCgNDDNF0vnhfM4pneVM2TKM7LI/Lx/q49zk
PDpTEr0tjhuDN+7ji835jVTlnDkeU9NJOk6KkVN4diRww8FkLfjg/vuUJa3wHnER
Qmx3APaYF8uxbk9r3LxQiipW4aGRkUVgy0Lq7IQwYSsZsRTnM/8+m8tIBQNCSjHn
l9fjby9P2iqWyrxeTxq2cX3tlcaSsPAiFQ5NcWmBOxAK2QsaOYz+jwh3jB6L1CZ/
dIZjc0ySz8AFnSo8TBYdw4XmYc50UQ7zq9cWUGGEUmV2jD7Ia+jeDPmjoluHwVit
fYLqIEdewNOmAQctWT32WYI1ZHC/bVCWAWJ+pdKuAx11U+J08unHppNDWkgvq5/d
YpjdBcO8mapsWJV/AVjpGi0uGTQuGFGi01HjBoVNbJGt2QHgQB1c7t/gDdUqljL6
AwyI3OL87fNcC4OPP5psCgUy3vb2b3ijEp/CL9P9eN+tiVVYytRyhACVloan47pg
ykiQoAa1LsLATDb9gjK12QNzGaPNrPlUZDyp44OoFrzKkhYj0uemcuMvPNJhyup8
pA+ReQLVyxrTu7R2fCIGZeQhpl0zoXtovsOJPIzAfj9hCGp447Ggr1GitthDLxjg
G19zy5imGb+wqUpjV/71ZMjYVLdkWQN+U/gSoiejZGbI6prSvi26Z8wM8m7I5xRT
EpaNVz9hLL5Pvpg8XdaAiXelmD++ZqNi9/hNE8qla+HtTiyNb9HR5oW3XCSrG0Gd
jg10+fUcMUMCxxrN+eA88WCQsTOvS9YLzlWyP+iVXPid8fbOAPKzBsqbTcLMEr+J
yZaG8VYToUePN6gCMVumkkr5hwpPN1FIG0m8Dk1FQLa+C5jSwPqcY2ydnTkZ11Xw
1rQegfFffyaIM/x7LFgKzvuP+1lQL58BGa5/tkI/On9Kyf/5IPMDMqHKKvBjiC56
rpU5Qi071hGBIfd0/fkHOj3qzUIugmH8Ni4roWqE/im8oCcbRcOVJKg+sGUCMpTZ
lT0T8j42PhdL6+UwsD4gceKQUj4ml8R8ELsivW0AEuayQRIGJuLvrVFAsiK4OpRe
/esn/sfAvP4QBLCwFRcVPNSo00EdYxqbpnPE1zUjW5DZ+lPP5u93b/KmEucvCgzX
OiL9FcETG4Arqg8FnhCbNn2WSNEViMliD8SV03TPdra25m6bN10PyUFXCApJl9DH
uN3FPONWF+nwwkJRkcftQhP4dT4K6q/9k13JPMw33Eytl8nrsNHSBGwkb51WgcqW
tAojCuHKnTvwbgKo8ulJkSBQ0cmqCuXnxCP59QgGq8OWXywBkoCl2LN6wTkD9s8E
PE87MH+4xTLEmcVQd5qtl4Jve8EKfcCmZ4Wh+UQuJoZUOOZhQWoindHjBEF/t9lf
XUebjjDfnoq9NyuVyRRfJy8ibalkEK89YdRY3nmyMMjF+nMdLamxUhECb+jnBMqf
cwys5hHp59D5b52ccPtOrbBO03ob2iikSTmFTcmxvEfDVloIKMPjuYVGwbg7j0C7
8LENGDjSg+MM7u44xi2n0t+Wq1uRPXvI0FslfOsoRWaFPuiCaQ5fVlFq193BzD9X
K1Xuprofk16uEwftOTjU4XJiKC6GT3pAGjVOZ3Tw3JKrtwXI+zk4uln5Co2p3vpZ
+2vZ4bBOUswvx9MDiKqOCvCuwszRB4MihmqZ8neV/14Zr3mPYmvtDl+L08+4OSJY
Fpts8ToPZlAH4Vq5zaWer7TwV9PYMqQjed4+F3dBSk6hLVwedu7iw/AfHGSOThUg
/laT9bFxdOdLUOIAqj0krYOi/jx/aJcenqkQbUOLzXwhcP1vOz2WZ5usaNVai6gr
1U2/zqPOMVPrXD6MWG63aLO+bah5MQ4dR55kZAiaYUH7isUpwsPwu4M1AxavH6fu
AXSzfxe86YklCpLGdFw8uxYBcpJB1+UMWn7TmgJAZKjzPtykk2uk8VuiTuichz6Q
3ZsxsV5Ta7NigUYdMZ3bBPSUUqicAPalBh/5MVnjQ8JH5W26IHsW2v7oQSm3T7Pf
OKDOEaQP7n4JGCVCAyN2QroetZ/WDxOjsnJ27bepk3M=
`protect END_PROTECTED
