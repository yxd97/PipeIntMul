`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1pbOsuGiXtstUZMrWNwnhzaSTuupTjNIy5qInZtALahtvZRm1A8apaOYPg2a5vd
tXMZn0EJXoJusDyxxyI+Zui9YgKgNZ7BlYMduMrwlVjXHRBa1r/psH6ZLyGnCoX0
TZdlLZChH44BYj0X3MBxE6UdCsVNmWunFT+aR2V/kCA4B2ukz6LHceAK5j3OSigl
RLk6d/PJuEZiQ9uj8tGcdopKQHUFSAMl3Gg4QWXDONq3RZTRVzZSGuG/06TFo+9z
aVZSJ8LPRrlLYu/ZKicYwg3+caTJvAnth5T8SI8OXAY9+6z+NcNm2NBLDupzx9ce
OeOA0Ek6lNJ7ueZazmVzVqeoo1SAWW7etLHe0XgO+QfYT+gqovqvrh0SsN7pShuX
xfilcWoDnGBP8kU4iP3v06bOQmtx/1PoJ2OWwHE7GgspBj79c8srJ7TCrxfMNbOy
QGHi2Wxr20EQkITnR7L/lemFMfbROwi7S7m1v+IprxY=
`protect END_PROTECTED
