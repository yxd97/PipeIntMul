`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGuQEUabJ6bBMegzdNyuJKxDPS7lGBTbRHwqev6yYZ46upfpPfbYCGWo9l1iwWjk
t0OiVYfHHmHovLuUtZCQowydUrwz2Qe52EdhvhKZnX3k2mkAyB42OkKEWXjD6d+y
cNcG1IMOkoropxFnNGBgx0phHER/kB007VLgwE3gZOB++55aoFNBTt0J8OBcTKTX
lAoLyEV85Kzm1vbKnKZGO6P3qYhcWrpGcQBr0lOJBJPH35kehfZuh0kpoKXioLmq
uWgnZI+qI2ilDI8rTouW3EfhGaob03wx5tlAHLPJ5Q0=
`protect END_PROTECTED
