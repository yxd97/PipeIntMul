library verilog;
use verilog.vl_types.all;
entity X_PHY_CONTROL is
    generic(
        LOC             : string  := "UNPLACED";
        AO_TOGGLE       : integer := 0;
        AO_WRLVL_EN     : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        BURST_MODE      : string  := "FALSE";
        CLK_RATIO       : integer := 1;
        CMD_OFFSET      : integer := 0;
        CO_DURATION     : integer := 0;
        DATA_CTL_A_N    : string  := "FALSE";
        DATA_CTL_B_N    : string  := "FALSE";
        DATA_CTL_C_N    : string  := "FALSE";
        DATA_CTL_D_N    : string  := "FALSE";
        DISABLE_SEQ_MATCH: string  := "TRUE";
        DI_DURATION     : integer := 0;
        DO_DURATION     : integer := 0;
        EVENTS_DELAY    : integer := 63;
        FOUR_WINDOW_CLOCKS: integer := 63;
        MULTI_REGION    : string  := "FALSE";
        PHY_COUNT_ENABLE: string  := "FALSE";
        RD_CMD_OFFSET_0 : integer := 0;
        RD_CMD_OFFSET_1 : integer := 0;
        RD_CMD_OFFSET_2 : integer := 0;
        RD_CMD_OFFSET_3 : integer := 0;
        RD_DURATION_0   : integer := 0;
        RD_DURATION_1   : integer := 0;
        RD_DURATION_2   : integer := 0;
        RD_DURATION_3   : integer := 0;
        SYNC_MODE       : string  := "FALSE";
        WR_CMD_OFFSET_0 : integer := 0;
        WR_CMD_OFFSET_1 : integer := 0;
        WR_CMD_OFFSET_2 : integer := 0;
        WR_CMD_OFFSET_3 : integer := 0;
        WR_DURATION_0   : integer := 0;
        WR_DURATION_1   : integer := 0;
        WR_DURATION_2   : integer := 0;
        WR_DURATION_3   : integer := 0
    );
    port(
        AUXOUTPUT       : out    vl_logic_vector(3 downto 0);
        INBURSTPENDING  : out    vl_logic_vector(3 downto 0);
        INRANKA         : out    vl_logic_vector(1 downto 0);
        INRANKB         : out    vl_logic_vector(1 downto 0);
        INRANKC         : out    vl_logic_vector(1 downto 0);
        INRANKD         : out    vl_logic_vector(1 downto 0);
        OUTBURSTPENDING : out    vl_logic_vector(3 downto 0);
        PCENABLECALIB   : out    vl_logic_vector(1 downto 0);
        PHYCTLALMOSTFULL: out    vl_logic;
        PHYCTLEMPTY     : out    vl_logic;
        PHYCTLFULL      : out    vl_logic;
        PHYCTLREADY     : out    vl_logic;
        MEMREFCLK       : in     vl_logic;
        PHYCLK          : in     vl_logic;
        PHYCTLMSTREMPTY : in     vl_logic;
        PHYCTLWD        : in     vl_logic_vector(31 downto 0);
        PHYCTLWRENABLE  : in     vl_logic;
        PLLLOCK         : in     vl_logic;
        READCALIBENABLE : in     vl_logic;
        REFDLLLOCK      : in     vl_logic;
        RESET           : in     vl_logic;
        SYNCIN          : in     vl_logic;
        WRITECALIBENABLE: in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of AO_TOGGLE : constant is 2;
    attribute mti_svvh_generic_type of AO_WRLVL_EN : constant is 2;
    attribute mti_svvh_generic_type of BURST_MODE : constant is 1;
    attribute mti_svvh_generic_type of CLK_RATIO : constant is 2;
    attribute mti_svvh_generic_type of CMD_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of CO_DURATION : constant is 2;
    attribute mti_svvh_generic_type of DATA_CTL_A_N : constant is 1;
    attribute mti_svvh_generic_type of DATA_CTL_B_N : constant is 1;
    attribute mti_svvh_generic_type of DATA_CTL_C_N : constant is 1;
    attribute mti_svvh_generic_type of DATA_CTL_D_N : constant is 1;
    attribute mti_svvh_generic_type of DISABLE_SEQ_MATCH : constant is 1;
    attribute mti_svvh_generic_type of DI_DURATION : constant is 2;
    attribute mti_svvh_generic_type of DO_DURATION : constant is 2;
    attribute mti_svvh_generic_type of EVENTS_DELAY : constant is 2;
    attribute mti_svvh_generic_type of FOUR_WINDOW_CLOCKS : constant is 2;
    attribute mti_svvh_generic_type of MULTI_REGION : constant is 1;
    attribute mti_svvh_generic_type of PHY_COUNT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of RD_CMD_OFFSET_0 : constant is 2;
    attribute mti_svvh_generic_type of RD_CMD_OFFSET_1 : constant is 2;
    attribute mti_svvh_generic_type of RD_CMD_OFFSET_2 : constant is 2;
    attribute mti_svvh_generic_type of RD_CMD_OFFSET_3 : constant is 2;
    attribute mti_svvh_generic_type of RD_DURATION_0 : constant is 2;
    attribute mti_svvh_generic_type of RD_DURATION_1 : constant is 2;
    attribute mti_svvh_generic_type of RD_DURATION_2 : constant is 2;
    attribute mti_svvh_generic_type of RD_DURATION_3 : constant is 2;
    attribute mti_svvh_generic_type of SYNC_MODE : constant is 1;
    attribute mti_svvh_generic_type of WR_CMD_OFFSET_0 : constant is 2;
    attribute mti_svvh_generic_type of WR_CMD_OFFSET_1 : constant is 2;
    attribute mti_svvh_generic_type of WR_CMD_OFFSET_2 : constant is 2;
    attribute mti_svvh_generic_type of WR_CMD_OFFSET_3 : constant is 2;
    attribute mti_svvh_generic_type of WR_DURATION_0 : constant is 2;
    attribute mti_svvh_generic_type of WR_DURATION_1 : constant is 2;
    attribute mti_svvh_generic_type of WR_DURATION_2 : constant is 2;
    attribute mti_svvh_generic_type of WR_DURATION_3 : constant is 2;
end X_PHY_CONTROL;
