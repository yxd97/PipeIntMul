`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ierydxnd/poSsMa3jX5dhSDavJz77Antvz74rZdKzdHoGtHrI8sl1zw90GIkeDvn
ZWF2Vdzs7ZxBS/2XmmY72muc7sg+iXmNp9uOrIGKQm1m1ZL8gnuozRVbGksSEII4
eLpURbALuhIXWVoSq8RNBT34XB4Q6GB3u2foIBkZffA387e4lWprSsX6OSV8+ptX
II5IMNk1ABbpua3yg2tMbgwCpXMBzMGvw0hhopbOJaE6p0tOKw5/h6xlFjFiFa8l
ox2am2xNNRAIIqUEl+6tQzNowfHEfTU+UPAeXqriI+B/NhJi98InsLlGj9qYHuSh
/o1IEPQCU1umdCS9kgGzC2GYFM/QPWd3LT9AEOzJWse3HmHRarzyoGerOe3MLnig
JjWhATwnHPikGtnKk0JwcZnZ+9FrJh6MZs1/zFEWGJoCXTSa9SyUA5kihWekowiK
ZcH0k1GnUNQK62VSLk/kKXq+R1mgNASWGcXM61QkK/lG79+s1bv//M5nx6klaXY8
B5xq9MHVOayq80fWsEUQ7uCPUDm6hKJqJrs84On9C2Ir8OQyB5KDrTTQQLdIWLh6
Hu8JdLqYd+ASJ+S5zihSXQUp/9zdX9c/HDcMDTBPl15MNS80npt+ZoXl6O2OONRe
GOWlM9RD4i1/vJrqWcDnPStcXL5UgCBtey689E+mcGgOUjkA6bTj+QDj9tP3dNER
qm9FZf52AqS6j2ZBo48U6A9CmVFFRBEIa1apRW61DxLVNWooH4lGooOBORkpaI9A
Bo/BUWBmfdrdDtnt8HJoXFXEg4VbHbr00wnbth3UEAsGHKWl80cB5lHeJtaoN350
4vqzTlJgczEjwzqxeO2KeemPemvWsVhZxDyTCNCyfeOdzRWdjf5hOKhJE/AxOllf
/iLW7SAd2KOmAYKTlWiBfJj9ugxwwpQBJy/kRUr+iiOAm/o9gKqdbY0o5+KLxGUh
XEIhk1t9uBZZJmsTuD9rdVQoo0+k7iqNphhQNCoASAU7BYyc6UgW9pAt+WtKYaPT
iMjRdNgcWUBcog12ilFI8CIWBN1nbUF6DrF7WafY/ETVpODeLktB9Qv/4ElGRalU
kid3LFAoJjLfF/LB3iteZdSxa1WFIusTBEWOgFyYqzgP5c0JSXtvSeaqKMdYwkr0
1rY07GyIRZF2qx5NniPpY6+u1YqqnpqLiGSMVEFYIi8gb1mq2qePDG7p5O0iChbr
bJ0GFcofxkem1zLtrRXb7Cq+YXKIBQ5cdXwDCc50kgRhiMgE+/5wd6fldAurDWLi
krhuH7Mt2dVMadc2ceCQMxk6RnEXcez9W7k+7u4IJeKa0cTz7pyxwtPNf5oUxShY
me7HJA79RqkK1rtQqQwlQUTz5EjS/RO5w+ObMJkiljuuv67D7XUqPxs4vUZvei2x
x9vfPpmphKmbkFtT7WDCiGM55yBDTxzeetZR7I84rBE3So7w3qtn1hvAC7B7oEH9
t+BLCj8DNV0dFPGzlmStNKuiSiNuqcPT3Ycz9s1pqgNEmSaE5DSpch+lBke5W3WF
V+BWOxGe2qfHmtaTexsJrz5/B530eJs7YhGJCBlrZfhMsNKi5NCYIh0bx2UL8jk4
XNivwkBarEXm42msDCDF6DqfboexgzwmC4jLzdJjxxgDsQGlmr9rdMikhEc7aXqb
/5OgrYDtSX+sv8CpMb0EblcXi02q+D3aczg51FmCZDBX07pQvPt+jKfO2dwwjsRJ
qG8XAFKvrSNc3HgVA7vGCkSuDFntlERqgSuX7674rm9Qnj4MGji0RQm5agxqnUCx
LeBJBPhaQkgwych7DsiEzfilVehipQ+QB4ghZ0GvTQvP7o4c4/EmPa5EeK3VnCJ5
SjiP4KoOLThNFxKGbW0QnHHlRVvocBE0GWy+cBZWOD01TklaCgnIxb7XzJnjTKZg
oBWn6/XRlGK7JC4gx1i1QstqRIl9iyokCo00v5nwvUppFBpfQQhlFGJGT8gZ8zg1
VGExnn7lUHZsiY/wh4lczNHQ/0IJmna8VtgznBKVN8CvW/eHYO1Hq0hMJkldT1Qc
+uXPtoLIIz6TSly3D2S/jEy53VGRndFs/lrZQW3T2n/kfN7RfkyPi+LkfcEy4OTe
f7aTwcvA2itdIdV+4ncCnnCkqxVKysDwLqQEZjzWYrw6Q5uES6liv/1O4fvfuSj4
F15BJ1eCffU2BB4UKSxiYlrB2KZ8/i/hFIar/O62oOJmn9vtL0fWLFedUbNIOdkm
CSXTBi63OADPuRs3PQRfu2Rb8Hs9jEMOXlxnmnd+KzlNVuI3BcnYIljMHklvByYM
UmL0DZUFbC54eMGnXCnkrOpqV77BsqguozRHJZEFdofjQEIOBCXj+JMJuWriIWQN
C9lJPu1OcHVurDc5RdVxo45wdYjsSd+YDkfGihO0cmbFvo9GJWkWu7owKPdu0F+5
VEcxAnzQKF671DNQljajrL+jSNylfIxDWHRJf3XxfxInueKW7ErXIGubYi0burRs
dYzoavXwlbxW9a3Jl354xXGeM8SNGOgOOy4qhzvBaMjqEi/H2QcpboBXjLiNzHC1
PJB8YPKu0YcRmMJrwF9rQ872IXQasBe8CCU667KIO2bIkKQphiuXZyFd7RiIRbgS
MHNNgECZHgNaNuX4srdtEOkJqrhnNbM2Fkl95YYXCUEYl0KYO6Otp1WEoEbov4/a
zw8jadZIL8KoEJMEFrQ2CT+vgeVyZHk3yBnhprPX8tf2I1gViQDCx3EOs9u99se9
CU3zIyIYpeLo3kAeze3pszI0sREqEF+GcEMRk7HrWpnVLBJ98xhZSlcDVqlMenx0
K03VBqDK3jeEyxubrDbEWlg5CQuMIqd20IRJ596UToeLSkZMd2faC4c27W5yAK3/
Qfu76+nQseTSMWvPpiSk4w==
`protect END_PROTECTED
