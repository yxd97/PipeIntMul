`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lUduh3b16MlESbekV9cdpZDNmqBmRiV/bAMP+Z9Ev847pgxSzWcNyeHQLRCmLTMr
AxbwuXOH85WBKUKJi14TyjJ2EnxO+QvA6G24Z+K9j3vgxAeuUtAVN+o7ZCx20AGC
dKkhdbewsZR2G6jkGpn96ggymS6XH3GOe7Ah0p9WvX0HMABuhOzx5DvC7OjnbyKB
UGgZDu+oDLRUOdHwPGCdVe5Aw/5MiLA8mab49VL9CX+g3Cb2KK1uWncTt+K124g5
gGjPaiPkcXaVsRJWCVUo/4EUI2S5CrXX9E7AWHHFw4WfvOaHqkeHQya3NkOYPf3k
pMXIZm33MYPp376q/3hhWHW7injTPTtNUS1rsJPyjjF9TL5k27loq5OpTEavF3lI
exXU9BtFDuyvtRnLf9NX2LGWpAWPXQqPAg8ISXuo0ElmlBP6JMgbFV6soPU+rLOB
G7GDRUluzoUrqSvVrD850vo2LiX1ig4gdXi1xkhCIc8f9KeY7/H21eBihe5/8AsJ
QQIGe0+YxSaujrai7maTk3y7euwOQ+W/fwv5V3Dk+85EAdxgYjowlMkBpXPc9VJy
GelWqCiGWRtojxL0WYhZcvn5hVX6z/2Q3uKBrqs85SGSmzFpgwG4AOzVNDiEorZL
VTih6fBTE8jvVm6pxX1aTTwhn4DYRDKMf+nhiN/pBV4a0D1O7Gs5veWrAa6kEaGH
AAH2XxyRkF6gC2gV6/tvB6qsAj/CnwKRYMSlU4i+9R3wVTzqRUEJFV31jTDFoDwL
15Tu/ywKiDvlVicPNs65EVvPL4RSE7EZQRwvCxmN6gAZo93w48gp6MigFSwT0+Jv
7jgi47mJk8FETa+ucPuJpc19C+zEO9jY03m13TigfoLxrhKjH/txzYSEndxCHFBv
sK0iHJZRySQD6CokHVBTgDIRsirP5Kdzsl6VKiKbYmxC2A79EfL7zDe16owvLjKq
/hNmbry1o3m5iTX1lxaiibP/s0bpcM69xX5GnGC7rKX8Sdi8lIeZs7Q2rdfFVZZ8
S6aJsV5jGHt3QRo+KWbkMIbW30YiCVnWY6gTMjsD1yGp34jUmrG4Mujfq05dfB4F
7uHJlpBrtjE/3j83yGyNpTaOsAMUfvhajlqPlzW66CdrHseEaSG6tpdSt/+kcz0B
g34mLBb7j4iT6MFSZwXTdUNpMss+rtxpHS5vhIX7hj0fd1xAztwUp5xxCQeohSeA
S0EunAsIzb9iCqEkxtbkWKLCWJ4P/pvJo7gJDwaXGO74f2C9vcFnwUY3rpn4JxQy
KfZw8CciSFc0j4aFBG1SQg5OG5NbCOV9H0pRXDDySdhJDgl6qn0b+xu0Mh412ifz
`protect END_PROTECTED
