`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VVomWuba4xTAB2558PfTpUP9Ko2e5ardY5b3XpiImmO6uuNeI/1OWkv6/CSfI4fL
wEcDy2rvOCarrEPYsWL21fgD9QZstpEwLJFW2H1IPjlimLJe7P5eXYye7zTvL/+z
sqOu5m1PHpyEjx8uiXCmCIc1qian90Q/SM3FuICTydPXDBCPZAWFW0YGNgb2grHI
NtFaRZwh+JowI2MrDEbLoWCEolOIR1RC0fEc+Bhvh5AUd7SzukmxKJdsB3nF/MAA
A+caUeFh/huYCYP9l/GqjsgK15HvEx7DYzBan05JtCxHU6+FdyuWFH2TieXvgZXH
d8xfY2ToIpcor8UTkbEJtSFxtultE8O61iZ+IjLT3QIJlXOpMRYBi+2o69gb/9uV
qnasA4wwjTP6y3d+whlKlcSuIdbj7iBE+COCSE09icUvwCz0RcPR4gb0HTUmuu1z
wIAK73ywI5fNkNnF+tXAo8dWlW0kmLC38RBRtaOjQbJmM89uaKipUMjDlw4i8sgI
CyMKdYcDbAKqKlK4FhOiSrs75Ppvf1WhjzJcZjLXtCIwpK1ydI2yxqAkroXZK1Ax
z6sKP1Ssj3nCUyApDufrBuXiwwJ5fZgDU/UVR/VtKLCvlVvZUO/YUgDnf4uUYdxb
7TpwP81Lxz6FbwcUAavCNQbJO5qEUNnmVaI2cQOw7sl+RnUkoyjNwV54nTOFo3/e
hm5zLCE8ZhpZkjmmg8C64fgSCzRZxmaT++NGQtJxsviIruci+HuLT6Zb5la2jk9W
1FjnDCmHjgQircXiC37cHQPW/uft3syZ1P84Egmve+eBtDPKnr6uy2AUnIZH6x2V
OHtr5vVFtgECGEn5Rl1Fhp9mG2O1vN7Yxw6xKqv4QwyN07eu3hUn4OZeFz7MYBoG
rdomR67zjnCZ5pg0kNrx8tYSO/M1G0Qm/xV4CxJzW1fExVkzoydCcJFUP364laE8
`protect END_PROTECTED
