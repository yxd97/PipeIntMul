`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fdje/IpAwn0KDyHdppFz+sP91rBTi69VLGYzb9xzcCZ7SLj3RQ9blrr8VFAOm/R+
yh5wfk/CAJ79eO5KIBXBl8/zh7akwKzmQD7BFDFnrwzDcQu1Iu5EIWCoOiE1NU71
Tkd5t+bmKJQd5eVpU2JO3vcjzm4cN/VqqIs8RyZVkL133fKZIXz5liM794g2JKK9
4iQ14HcRThejRpM/5F0I7kdFEQtOx8Wex/Hv/c63yad7FeSAh5rYq76sC3TcYsxu
gZgE5V3z9HnkNM9BszrBpsXAY8+ILAsdfeaiie4V1wfzEeYC+uzyibnrau8tUIwz
VD7q6DNChOzaLsiVI6MY17NgPwaf3WpBpKlQaDM70yIdzLhUjYeeOHJDN9+45Pfa
`protect END_PROTECTED
