`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gDBPZabB4iAAl7Rf8dDjwZUMjx70u3nByAAQt346m3vHlo1VynGUkk26nsxE1UVx
yX5afXLi5uShjEK5CB1b0Exk8f9EPkx8DDxKjElvfA9ADkqdyH38dqLGJQa1EZ6v
E2/7ViM4FYyvkcvG0FF5G0sT9TNxgdbyE4ZJqmjQ6P0BfQ1wuXvP4o7WnFDHMBCy
6HeUlA2VXISH0bHbAwH5TbSQWUjb0AflCJ1NbtYmMvoosH1tGSOX4naG60xyjTkh
m6vCZFs/OdqBla73NsUwMWLBh5B2xYvOroNa4AxeGZY=
`protect END_PROTECTED
