`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7fkm6mDt7C2e69gEMuyTzuYg1/bVE0hhwM4q0nho1aYKqQgh+C31FfanYkSWizCb
KuL7WPkN0R18cHMaVwM6J9HEzh8FT05w/Fg1xdtWRkWFJSIJtM/PtRsiPEt4pBNd
eefuQPlcPpaS+MyuDm6kLVTbrtyWBLKe7qu/CZvlgA3CyvfmoucsRPqrh/1WIhMZ
i+a6gBl+AmI/tuR820bOClCykxjfAzI4ucinWQwDgNwQhTj3e+XKN3Xnz77B752x
dk+6aTgXOFHMMfkk1bTFNVighXm9BNZ7oTx+aXivS7vp/4AXGsa0V/CunMuU3lN+
P8YhbjGz4Z2ihKel1n7KMct4r1Lzv/IwhEFgGshiJ4DZOlV0w85FBrsdiwWM/Ryg
6Z/6Xfy6NIqc/0+iplxMj391YyaNnDotK5BADLs+GlghlfqP8dY2powYSoyvrj5v
pMv9uNYSfiAFAfyaZyfbDDdkjnaA35G7uIxNkXWgmw85MRyROEp/e7qUKFO5OXum
R0kFCM4TwG8PfCOYO+r04ox19EQw4iwK7zvxIShcdltYB0a8a1QC8LzgwAkjuFtK
1YpNqQMfDw4HzeaNK7Uzdof1iHyJ87SCQuc2AxHMqKAKGcYicuogpkkcdA04UPPG
f5GuT2xcmc8sfLUuiSad+BZXGz3E5Sd1Ang+oSHVSC6IgaUYOfgRr7SPGbaGjVKE
wR9sv94Ds0Tpuh2+U2zGjg==
`protect END_PROTECTED
