`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHofL5FZGNr9yXy4Lxk6VRnuXOAhAVRM8+SBcZXkkLBBBCuGXhQpFTcZxbDgo4sE
N7pftYjGXmp8nmLoZL7I6nnmRPV8Gf5POkaI62NixEYWAeeM7K+Oocb7h111EGfC
NUucXxOuV50R01cmYUQSeyVpiw0w/P9ZKR2sxDxtPBuyWstbVRMWCQYOfxAFcKts
GX/pFtDAjaQb3ZgPZEYNbyuCV68tMo/VUil+iCwS1kKeanDkVDVkFVnQCCBZXZFy
XKBdx7+ZRXDOWGVTs8ph9sUPAucLEmxy3IhdPaz3TbN/TYM3xiVmMWm0RMFCtLdr
jMpmP+Z/iotz+yZQ329abx5Y6SwNRMo3iJ0MOrhfGja7UJWey2+WTRn6RxK21IHq
wO8EKF1VmhQOcwZLVGv0g0CSWcaSoZVLLwoqtlha5elNJCUJC5uhFCbwe5AXi9+5
XxGENI0FKEX4LhBfFvP/OcHvOU1oH3M7KzL1JrBBdL2IOT3spMb0M1+5o3CSsf+Z
Dsb+ZSOclEB8lYYmMpRLO8EhvdvbtWyBVmcteJ5u4AydK0enzFGShq5WLoqE20gq
00gC8HAKB3iP+ZTTYY5Y3Oe6XD0evqD+pgCc6PqjlDxFb25wisGEbqmac34F2dLd
5S5dymms5WZ/nm+WokcqhBmMBDPl42GX1F9EQ0CpxdnHQtywLOsOsLgdZw1Kke6W
U2uKL7S/exSolIFAsJckq888OgGhYMYYld2k1CbWX+GLq4LN+1/DWhX/1/CJYP71
VJK2Xwew3l8d84s0M/3sXCg/gGZRTnSPj0+cdqqylLB/YL8xwAUqtydYMUGYjJ6D
berPwxqcR54tJ1XcuwtLq/Nsg/8E1gmy8L2MALlIiJNkHeIm4ryNgjI+GkKRvKo5
rX/+LQdTp4YXK3dd/9W+8Q==
`protect END_PROTECTED
