`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ne8T7bNlZvMcr+EWm3zMUZz4wnKcHuEAs1xHnW1qBwH7X3zSkRjaO/kCbmccBAJL
57jbzAkbHVFHH6X1ZNeDXah777hq6/jQE3ePQeTpXFDpVEfXzmaV2nqR49ekUKYi
YltkcCqKMbhoO1g9IxnLAxw2fMNJw18ohPo+ILO5uq1W+1b7rxRMXYJjxQZj9VN6
DM9WBeO27VRqT4TgSJnRVl7Qk3Vin/5kHCD/9h26iNgeS6GJ7ezFMc3Tp3+YiP43
nDzjSGLDk2ErZo20wJrq3gh0+iUy/Yq/ki6dKeCKZNluntPKjEZHbxLOgYPl+dJ6
sVPnQ271wwrYvY91BDQD/YqQNtM+6wZM2csNimwr+Mh7ayq/8NNAXPwq/z6W1OUJ
5jBIGsaWjDb3cedBzo4Kj3uUV25XhTahJxDR/DiZnoGoEGd14WSTzuw7xD4iOUxK
6t1KB4tmEfg0sDiT6CiuVtfEPjYXxkUqqd+L7+98RF824/xlSObxnOC0dMw6YWMX
SiaxNAjYoh+k68ix6IY4cifEWoOpJ5jbKXlNUH1QT0HA7MoFiGM3+3wLf8XqexE5
8f67cHYIPeJU38l+FLGiusrk8j2ZPvmm9jn/PuB8JTklca2L9SX1IagEgfuMcjC7
WUFgjL6b0g8qR7e57jtV69PWqJxLW1Lj1CcTrfGKl9P+pt/oBLHCpotf1fCWJeOR
8xza0SLXPicuH0gjlWT7F6ZY5lUTQOfo7p5R91UioWldKc08Pe9N9p2C/HuoKBRv
JUoGcqoM6Qm1dWQkwv7WLA/2LxydMx4TJ7wrrMdQxTLaDma4/xUwT1z/92sG6a5w
A0BzT6cM4+vtESYjRebeQKxrz/x1FBhtS7oNnHrGLf2immCjjqHHZkpFhElYSCbG
/N87JZTL249mi3CMSJD+5PJqLoUcfZ+qr5eGMQlKD5KvVsQZNpZr5MKB3Ha+d8po
2RA8ucL38e38WwDiNbBWOk+CgNSSNEYztDQ2Ge1dXLYmlPZbZnBowW2rxUuJiEL8
6XCJTawdIl/s7Z66RB/TGirwNaLAlZLRamFhc9sMZmnkjpzt60ysvB6qZncRS0xJ
/aw499pkFx4144+cj83KLGtCxSU9h8TqhxqDJrKuXCs=
`protect END_PROTECTED
