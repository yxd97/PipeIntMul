`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Buzh6i5+4pJCgU1lNLoo4nu42vpu0rV41FjtmOyQ8PXUXYt3INESZ+XjXo1yrjWu
kK2tAcBWYurcAsTT+pD3Hjn+4cjqwnY3RaSUL8FAPs1CXhq7+ERKsUo+fOq/e3sF
KvHdKIdnbD2GnqwbZCZoV64Gq/T9XQgGoLeCqQV6Y5CbDkC2T1TqAD/3RJj6kBGL
CZFKWyABgxTrvPMkE96+GbdsyahF20Wi4+2AjXDwesKW+io8Yi00YQhkC0gIDt0a
72bOc0L0T523/Pw/NQDxxp75dA44w4TN5BDnb/TU3Z//5mgKtWT2UGIdy3S5I1rE
iteKqZIF1GQHVU0CfNoyhmcf+GxqtiLOTVI+lic6D8k2aC9rxsUhAc93lMlOxMmj
mFwJcR9s6nYMrxC93G+LhvnbPkeot3dM4DB7STrC75eEFB+seKwIgEVnVKE0OF7e
76J785APAJQTlyBhdPJSB0w9OuIZ+geVUxf3YP9RCIQlHJi05+qdg+I5+NiZ9l9U
n8Cpdi7pcZyQFmY8Oa/JYKpEYN18oKPCdespR46hONwwkGcYe5b3A5v7if3EW9+Q
/7jNiYKjH9pswF/5PlzU3njhnU+YTjFluXmnXTloJ5bvubhUMkrrPamn3tjh5D4O
5vDlJs1ArtGFOxiX8SO3y6eqCZQxgzaOUCu3qNpgOVBaeO3NFbj2/AHnVxcxYbdG
fp2bpfUICeCkLnyrhqIUFGXUKfIqSyJZ7dtQ8nyBvx1EOej9AugIPXMKYPzTJVq1
SrPQIQd/XWiGAozA2mWvmJQkSoQXzKXvTfzfXckBpA7I/Ahet03FVfYcIFiEPxjQ
dLx6nEHaZizTkXf2zcoe0G0D4gCVYZUl0hD7it7ZVsXwTQS9gQ8ochOb9Mb0phnU
ZMV9cXGbhPAWSsOe+I4EydT+416GZaLsJpQu55HyUaZ8DahfHsjQFTpU94ZePy1K
pGxWGJslWTTuV7qQ3OlVNt7ZdC/aU7GJu2loduwZOKqhDGtaq26h9AqxHahu8xfk
JCaRBsD6DtCQ17zZ4DqwcCcSCrItNPMrdb5sVlWWdRLEKX8033O/7yZ3yhNDV1tI
Xqx4seIlNkp6+wbaXoY9v6PuWZkNgJh7LPfYBFqMfr8pWd3vSh0x7mKjwrc+QTe4
nyHkAs93TBWg8yn+AcmlvaCpXUoWtAQGXyempaUPIJzxUBcaPv8yu5qpwsR8HuNM
vL93fDtKPW1PMr0CF3kPyCar1kkkl6bMO6DL8N2lMNcvsfdsZ7/6C2T437QKoLEz
4FpGyzpBWkvn4orh+/9GJoee12wfvNFmARFMvtI7TjmNcNSwk5M95YUr+jKII1Cq
pY6t2wZtW1vhExor4PyQtodzil1T/GK6yz2KKDcYwQwA+lcZkUoAJ85I37Mtb461
RaGdiGTSAa8j5BjpLauPhNiyFVGYn0AOch1OgWzy7D0gquOBgCUaMxiJ2zrxlwyb
`protect END_PROTECTED
