`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bKQgZGCVSTWpN+PWUr3JHDjf5Afp9PW3ExPHzeELHpQhqHBOHhlMs+dGKNfPbmHx
moK2AXIadGpUTynBndawbklocF06+bu9QQP5KzBIG52d/DBeDphWXbS11zIm6jjT
v+Z3W58yKTNsqP3QJdUK3XCZnPib9OfSgu2DUPQ6+hKVLt1rw61j1PFCFKoU0sbX
kXoMKUjzSZSGtzbUkb6p0kK4euCcD2vDb10hJboeAzszq+xOTgNyMcZYzW/z9Qa9
lyRW0IlQWpfdE1ahaZFpSQhvRS7r6cjM4V9p69uL/qO0fvvAnzCyPQbps+leUYLH
lcdWzIJIRA3GxxLUEs8lptXrSaM6T9iR6Sy6FQiwNQ6Zx8+FnDPeqgAk6DvW4Eyv
mdp86maua+PfGxKoWqwic9guWKgIN0j8dQkAoFJOPAI=
`protect END_PROTECTED
