library verilog;
use verilog.vl_types.all;
entity family is
end family;
