`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
81BndouwOx/ZAWbyc17KzhmaqSid+o6aisp6qPVKMqUvEpl9tvSP5mHUJtA/5ZCU
q6/TDll/30FV2vdItzqNauEfO1goGIPVL1NKOkrwRpTSFMQfiSBhv+EW7O2VgUxP
Dpp2FQ4j/0R34D0Oo6b/GN6e8T/afQCIDJ7l4ihFdKXjp1KqDK5SC87WO68acDYO
OSKBy0x4aoBer7NKLnamxMMByY0YBkhGSUjWCSuPa04ZGIKanCz4BcGXhKw6ZBWh
sVMIqtzlWkloLzM2iwZSeweyK/iey0zihfLbteeumszG03SqRYWtpECQnRH3J51E
oF8m065DoA0j8K6w3F34uqGahB2w2moARznMwylQ+EKI+8FxuwgyFRb1r6zAFAZt
zhZ457DB0jkNBM7LtmZtlsBUgS/UNNpeF0YwwlwV22lOHNwUYdPB2CmbyaSDdcYI
xieWaUcg7hr9bbX7GXm1v2ezgg5zTN7zAnJa3zWz3No2wgmcXskKYfs+w87EKFJh
Ve6hdiaCLRdmsWWPthETu9ew/s6myoXJmJBCYPvVNdub3ZngRakQnDJaKoYZegYg
Pxsojv4opXktmrfq/4XragErzqXQkRlNpvzq2iUEJl/fCMvGfs2Y87S+nE4ntqTu
jjbNZ821dZSFg4XH8fvwQdd3HnxOMuxl67/ZT5twt907C97h/SULXVr/DYG9nVoM
tmtezyq3K38Hv/y8uKJOaFVVIBGa+NYcl7sAf4pBNIogce9FTihktS2P7X1jwK2X
`protect END_PROTECTED
