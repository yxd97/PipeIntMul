`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkWVcID/F+ukJ7nnGIWybcoMV1qarhAMlw55fOSd2WwZlteDlgCyNQWGm8pE18KS
DL8GyqR0PytgqPu6ca38FebW6ddUe79WxQWcatV6y3wyH9lLUbQryxHoBBtu7+zW
/ze3Xh8kVrpWTXmPMw5/GX2HXfggwTDBMzB+TcX8zt5hrhmTFBAtTculedZnUbHm
BLHEJQy+QUQas5W8vvrx7NPPzGDSZ3k7Uf7P7s1ARH9LfaoIb/ekdrAakztSJIcD
hovhx4wSgLHQIlvrRWs6nq6yy/+ABHnRw8Ll8/UW8kWnPiUdUZdJ97Q3pj6dFQlm
MTgqVKJ3tj7wdwNj+V0JMR9RbBj1zglYfKrKJNgTsGqbfAcXTmbSvr8HCJmWb7d5
/InTKLvhUkDaYSxZRH9qIb7pzM9kjyxMGxy0qSsVbQ+Lq9mDtRgeBQPaKl2xGKUf
JVNow+O4xKrUcLnX6wG0Og==
`protect END_PROTECTED
