`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzT4bA8r8uHZsH+JuD+8jwIbuUxxaHAsJUzdFcvSBVcssNBo1z5HntNnBm2p+Nlt
Z4p/U8NhiXBJgO6ZT1A+JEqxdtaIAhP1//MLbyQFrk89NQjZpzcOD98c/2UqGzHy
eoQKVcvJiWHe3m53QUBmiIufe8jh/vaiQ+N3MRTUDJaMuvfhT92TJB70PJdvG0FS
V/tlH9xMTZe55m0fYGCv1/QdxoS/InBAL0r9E4O+NzadMnKHD44nz5cOYamU3vLD
6LIevOSoyLJ/WUeZlWVetE2IsLHX3HpHyuLS+kW35rjSdyQ2o1yT6Ee8F5QuKdqB
k3SJJngy9XRUS8XbsU7zlX8SxLYALPp/bXvSj8oR/KRnvs4swvQpql8O7WwJYrkt
Qpxfe1XQJfgKzRGpP0DbiZ950G9M1/abyyrsRcfXvmW8sVE8XbjOApPZ0mA7BE+2
HKxq960Tj+GazECxonyOZalCzob2pz1NTtbxSxUTyeiDp6LkgwTPGBretgAE8i77
sMZ1BVTkh+I38rk9gd8GP5a+Ds3++houlVL8DjGkYD7sE6JX4anfs8eDEpjIOcRn
I93XnZ0K969cwW4sWrdpmKiTjk6QaATGCwl7i4eTkc8YmAot2J51rNTSoGmYWOeD
rO8A5ScTX2qzy0bnhsPI8A==
`protect END_PROTECTED
