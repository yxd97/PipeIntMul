`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N8SgJ+9Ff68zO4Vg7oFN6H4AKb5SfXUW/JBijAqunQJWMyvn0e3HiCiRUB0rTl5/
xnOINGEcEOmMI8TUtuhduPDWp4BvOZThvaxSHiI9+CUW0F1zVSQqu3WNV6bBj5ym
8MDN8dByPuoxG1fuFAy7LOG6eYXErHYYtzxsCPIJkcttsS96lQioOztocIboVE+9
GHgMYM+zCSl78MOhr6jFjB0iFpmUgS/73RAbPygmOF4ZdCxxWFA2kKjuCbJk2Wtr
x3fRx94BkkrHln2RODn8j1SXmkfrlR//NG5mIQRHwc98vkX84nHAGlGtPw4nL/tI
R447LwQrqNpJ4sF77Ip9GpF3iOL8R2eAsuRM1VipbA8k+d1bLjmAhc7yjDB+6r6D
u6w5jZdWbwWpYaQ3U6xk8GvnX0e6jXf42PT/xBkh8bdiTsIT6983uY+JtfSVcDO/
Q6yNMGzg30lyHeqh0Zw9qxlGBeqPNFModvDBL0GWf86oMeLsmHdWDVTGWkPArYFD
DR0c+j/9aIhQZjyzc0ex75SGe0kd+mmQKHreiRDPjx64HT7TbAdUSIFVsSFW7vDl
ovDfQ33ndJpci7A6K/2VQ/39tkRdzPDamYsfZr/+Dbo+kADMs9TZZxvEtQX7clw2
F64nd5QGPOkibHbF6f3gywFinbRISgIBT2LKOqqz1o3DquNVNnWvzo5mDRnq+NCi
iB0ar4+kFr73yJYVvakGGHh4kthJvXuEnQwesaxBUa1/Ipy+Y49k+0mPNwKTisqT
N576nxZfkCCEzNuNqjf9vMNaHtQ0WebBoeB0R1e8h7u7QQoCk/UbOl1iugggcbG4
TyfgkZ+tbf2Iv7itE/KYUwboWNA94x4zBzFCzvZtSjVMSYXxsNj//v54+MZYf9Ei
eYXh2PlYqo4OwrSLv5hef3p94RYxTWBb+eYaTN35uVeJN+ktLVOXnI8KsZGiRaZG
/+VW0sHp8d6T9r2Rr8suhJnWHQ24kMIau3GKpSLfLF/BV4UBfwnf2whUlLGTKRWU
XYGKQ8n17yAwKOcizGj5TVbwUAbdQJqbiiqPh9YOI1SllHEeba9vA6n/rXsQkh4l
tXP+DTkbEgemJ7r3D1/vLssNOesy1zsdDFbSLT7nuZ15eWr3xaA10R1V7R0613YL
Z0wFdeVtvA8ghky9hHYmXRE0tpQoinUbMbVMjYwwRO3ypvqrojn8HUCW3II0hEY/
mKDbwA8Q27v4W0Af3t9QSQ6BGEia9TNFrso0SKb7wHsWRs6ObBCOzObuNdDrPAWu
eZxOh6JJo4Fph2Wf4TU/E1g4m1aeJ28fN2BpN24RwcQvR+KIuiD+8qZclemC551K
4B+EUJjjLkI9t9y5cJpquhdq3zX/nmt/AocMIapmxOCWUIWBrqZUX01dHZYjL3DP
6UrvF19zQGaKScOsptMQ54qHQl6oeTb7RFON0VXMZN6x5IkOM8Eha5uEt44E6Yhh
AAkn976YD48HiTdbXCyr5a9tHPKuEfznvw89w89OPWs1/UQG6fUS+nry7eB/H5yI
MiCAN8IGq6jace62ySyMjYNCfQYqW+CCnLeaLIxsHDh8ZKoFwrbUwVr3XqoK9jvM
xGL/XtVXhJSMgbGliwjciMm/S4v2BNHPp6BINzgb1VmoDL5X4L4VXLYvNj6byEte
gBwsvGImVC+FSX759NLGgOSO24WddxqcEelRjjPEw5vTfXl7PIQqF+7fPUx2DCC3
e12Kfib7D4Ea/6T1FszNOpkRnpVKIPFVkdZLsijvd6RW62jE+ZWsTBLLGuMQeIgv
MV0jp9z/JmoDdPRfI1dfAlO4Xqhd688Nj6sf/AohntOP4SfV9GPpFS6CqbRTJ+lX
dcwZGN2bHYd9UJus6Zo6GrdKaJ5QNvEufUR1ohFPJCggyvEximsvTyxesJ+P+hBZ
8LlOKZi3LAiLNaXMH4MxA/wR/3aJ2D4SItn8GJP5FzFv3IsSGNOcJCEatcN++Rnw
G9s1yfM2/4+zwmrDiP7jm4U8c9z+9rfJBsM4hO0OvzR7yAn3iZNeXXLvLjhw+GSk
PHsYDR1TB/GynAurgBBrhFBrmz6VOcUYU0Ubd6KP9PgdVlGdZi46hbzbRDD5/g5K
gfUqu79Ym72W3Pgyv+FFTyFGPlxTydgxZe2oJxRbSmTi7FKUp6HaYKhbXbXN0Lw5
vTj118oOuxGJ6loj07qiL6qeIweXw8l6DBhD0tG3efqiyn4zaUvEJ/bv7HYyfsWe
3r56OkbnnuRudQ1+u0tjtTPWveduGLxcH2QG4EuPsDuqsIAb0jwD2eGMTSjOgaxf
1ZYnLHV3eJDe9jCAR0lyWDgxRlAkvzC35Z8sbHCL34zbLUh/jEvTYaSSqJylyhva
y+W/JLuPhKWH6zP500Wz53Vo6Qeg1JHP5KN/CoM+zxmYVWE+lsgypwdTcyIJ0MEi
QlYQlBSC/41NHHf47r9uKm1LA+z6Sq1W8xYwjmCUSn/Y6swr+6htRMCFOkiFhJ8E
lAITU4ER7dKbw2nJb2hKabjV+IUN3kT0JaYUewSGJfLpubWirZegdz+Fg6m2aMWh
VpkQid0XbUer7HuKSbgXWDdTuuA3GfXtVNkUablueK7feTQrRv/3619xy1Wnk6cL
Bj/QepOFsOi91a8lHmXGFRa3ipWleg5ln2cjQikFBG66lD5yujyt8MzjFH0CbW4x
hVCDzObg9LpBOl+fuKvrCeXvE36TJeTwTGe1eg3S3K3ETMEH25pBsEtZ1av0AWbB
E9s9y8Z1wzI86ZPaU45bMkkQO/9ra/in5uF/TacRRVik39pYP7fx5izGGx+nltz6
+1v2rZQDmd99EE/9E6Wwm4hxqU3jDvdlZ7nvKo+rYL9BVNIKH4nAet0cUuC069lA
boXt7Y56a/Gq44p/G+u0AipI5kgMbMdS34fMvBdhZGl436bmLh30WU3pwTeg8tqC
NLqX1OTDYZBnK7/lpAjaDeNBPpW6C8WcitBstxbbF4tC2FU5filXpMPGJPQ4brT9
sxmzh7xFG5hzOl9vl1a+BkgS1BHJckiXCi4ozWtVTzQvOttp16ZSA3+3FWJmOdR3
PVB9T4QVJV7Pp+JMvkceEujip/yx3zuesath1f4a1cK0dRyLAMROA5Bkpo245W/J
O4SiHli4z2A1YtN8Jro3w8MnUOQ/WWjpqvWF6E5buT5Nc/7sJ5Sc0CTnzizvpPys
Rtp1/3ymB0D2kwv1STQONckcZKEGMVUAaFet3pOYp2+4naB2vjh6pKyNlveHc0uJ
nw6nO3dOcJUD94NLXm1TI7TCvTCJ7AVmQ4CSOVF2WsY5t1gRfMhddXrOs680qV0q
VmKzcBx73s8wb8OS2VmoriwfIH35mpvCGSoIOs2e95V6djRpiqpqtyfC6FFMXiAI
vA2/Ji4ktp5ibSLSW9jio10vCbhPeaThSlLCDnd9nxL95AFkCNnsJ/jQG4ywa9X8
3jVHfkFzTJ4r4sKMZqU4LWFfOKpE1sD3+jqU3BcvoW0RqcBpIYTKUwDktYeSY5dN
XBIX5mdYgn3MZYfLnBYNOkGsty0L2bA/1CI2VFUJ4RONfPX8pIEsY9t9x3NQeuLd
W8Qv7TvxSogQToFiCRSgdNXZfX0saG7++LXamVlACZwR4x6a+V4sUn6rlsBHxxtD
Xm0/nQ1q7C1mOYEDFRrB76s296a0vx9Gpupmgk3txfj9ew7/m31mytr171lBotI4
q3vrKcywOTjL30iBPniBjCK8AbXVIEu9gb//SfiHCXrX44HrbJHaNWvDA4o26NyU
Y5p3O4h9oEAzMN1442jEwjpPpWX9H9DM2NFVQEPuFqv4udH01xV3q7wbfsb6DvIx
miZbxKteb5yBU+DbqArApatB7q3MDAJc+sKgNU33j4rog/Im2/iY6BWUwA+dlEP5
G9tmdCNaBOhvwdhDJ5Jzl7Z7wJtUQGu6Rs0pXA7Kp9tf+4NnBWluygoynIq7Hzaw
oJBuYIGKcOZLbnv7Gp01wF97TAo5syvpMb0AxmP9jYWRHj0g1iddvzUvsVmxBLrR
BLJAHNcVB0Q2ufKQXsKr5vfuUED00Xi5FfSDYQCZTkD+KBbaLs6U3mTIL1oL+fG4
ixyp3PhkEuAPebW+0+ECT6OamsR0vR3JzHrFLKucbAZuJha1//ydB77ngcvE9qN4
CIPmcHZzeGK+VsEsAkPI0pkxhKeC2bbs3jZUJZY9/GdIkOSUmMbiVM65AQsAYL1T
u8cAeJ2NAsbA0IaL5WDnyKzD6/MspkTE3eN8I10jj8OsjkFLynmBMYVxpJwHmDvj
`protect END_PROTECTED
