`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Lbk7Xts5gbjeyg6Os6qqvdxkowfFQn1an+6hMCV9OviG/UuWp97eZaeP+VWDQc6
HdiLe2e8u44AEw4N9mWN++o7PtGLcCEMTRCYmawRY2wCn3z4m6kmqejjunZQjN0C
CIzkPaP5M/uxG64mcHNydO57X1BSN4OacxpK17/UAgtW/JY//Oz2SWmerfoKZ01i
/kGz4u1QS7p692zomys9rRKbk8kJqTa7JxeuoXhmLw3GNSPfLAjgylSiEcDppy37
PFw4WorVr6AwaJhL51jGKdo8c5pHK4rnzPP2hUUuGKDz4XHPt57iEoOu/zLrP/Ye
4vv8XLoGuoD07k39jJGQtI9KjXGOwuKEfTWWR2KbYvmNxwjqj9Oe2eWxu2vMJCHD
+nDn/dldAzp8c7HZee3WqIn/9vxbpkpX6vx2hxK/fYFd8jpRyE7mrs0PrnO+pFWw
dXY5Xq5xR8kGu9jSX+9pDIYJZBIzYaaBoKP/l/BD/ohPzbZAkjVSk+PeWZneWU+8
riPPPPbzNYp44PIeSfI6yXPnMHdk/QQHue2E02pYIO1cKcHyTZ9RYUymlYQBqF2g
ve5h8i13sDaUKxy6uq8l3I0i8lQ34yF1b53CTavhqS0hABaLDbmM90KXkvTgNovL
3RJ7eWF2FyOnfJyX8zqr+Tbd/CWad5BDUwE/KQ1WxdyCNkgh4ilKKdBnjeBkwgYP
rRSo43yvgWobgj0ShNz5IljVAQldiRMrF1p8CJRbKXalkkqzgl7ZqEzMNTJiqETL
Lij2/5Hnw7M6a+00vVqq33EHKoa6TwH0IekgGVwlyhl9If7/Ps3ck8ai8W1RMkHH
R3LNu/h0AuESn5VZQ6IjfNzO7KwvRcx1lEdmVI6DirsAvgl3HOYamkV0jzp7nqzS
CuTZeEAaS8pTazLI0+LqS9FlPO2qqB2o/bOinP7xVvx1vpJK5tHdcorj05c6xqCa
`protect END_PROTECTED
