`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRmUisUvZs0X8OcOV4jcAtY9jAqILDvQRJi263KcD9KzB4BWgHY8ci0V5a2+oS1c
ydNFHnasrhNHUerOebRFj6Q2TtinZ7zYgZMeEPe/CxA9rPkQpryVD7jipYyPR83J
PqOcNk2tTTDB8wUgWFchKHOADZwgPt7JoI2RzkSX1yv+uBkjmqN/6+PWNfRrEgX+
Ap7qFnyt30nDQh8TbWcwr2zaIxe2oFB1Au/AIgwqBA+QqQMs5jspY7Zj8cB+VOFw
D4BokQJD6ttKbEIJzfF07nmLa64MqqeM9jV7fbFGspwoofLYwsu8dpItfhv7w9YO
f8jgohxZwW4XR2WmtpI65pTwg3BhB718MRgqadhpmg8zMztNN31Y1iRKaCR0eukY
sDOU4vUbFSfVT4wRZOdYNJihBHn939p/aeqZbATvFZrN4E0B9AiUGJHuwaQ31Vl7
ttpj3boaWuMj2ZIwtG3PbFPYj/RlJJvQeAbAR45fH3o9Khf3dzGFww6zK07MtcZT
ck/EIY2FBMw3ybyA7Qjw0uLKWBihrXVukcbx6+TvXl6wGIjkGZnTl0k9fXHGisDm
EzuM5y6ZfxpUonf8TT6DZogdCz3dKzXUjx6jm42gbA96Un286iGLi9f/Ctl/i9bR
gLRI6Megv9Z0K9xtaCIO+L9nTA7oSyp/p48vNc+cC11T6mAirmrYjK2e7AVGiiy5
oiVv94OCTg2XpqBUjXsSxaTo7qeI0kcgJ8RLKmJZkwEeG9q5u3QvcE24n7vil6lX
arZRGDE/ATo2Zi0J/K5TxlfjFCmPFxuF8dwHZRNNr+W824L/U1hLORPlf7+J12F8
nBF01bP1AXVXZX/R3mg4shHu4aamrstwpIlo9T1Dl5QpkLAUqRDOnh4iQNzd1dxC
ysF6ZkOPcF/NwkWTBZW7qBSZtwvpE0BOHtISBzorpk/TXsWIcfyMtBA4iqmb+7Im
n9pSzfKKH9EsEc6ehfNNrwfZz7xwCnU1JDIPPi0pNykhh+8LSXHM2zSjZNF3Saii
`protect END_PROTECTED
