`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RzNmoELFQyx40np1EfM7yoV5y55JH5GNvNgNuEHn4IfpKr/rD0Pom6UjEv5lkIm2
Z1LmObFptI1kfDSQ5+NBvwctdrtY+etvlzhhAk/6N+/ZB2IV0HCRUSvLComG1LtF
18yK79YDUj5HLDvst1LZF5qQWhrX/mtEzo1pWzEaXqPwEeL1J+MJLhnxvIzbfgR7
e39Tdu5XWDLzXOwbJ7qRokthlMXcbu6EFgFOjuKwNnX/QZocVNP2S7YdFPXMLStf
gvZf4xeYpVxDJKnveArqgPHbbDK9LTjQC6sZrzkN7sAaGx2RXWHOTwvmNJ1ycLHb
PvLCsJOmOzBHFi8F83dLm49nW5wPdsVKzCtQ0EaqGt7Pka+rz0u7pLiOKMdYTbOw
8gkkNhgW0aWZXq/CrFltQXKZg64SHnEePk2glCJzh9YAygmn7wcMhgNlkmF7ToJZ
uTWiNn81x3mApiStvsXWdBKHzskeuU493Jxu9BuXysb/jbXBeXDvmUvp0F2bkpEv
H6Id0E0pNoHD9pjacBImsURCYyh037vc9c/Yc4v5hePoIQt7B+y63KjxP3pfagtE
yjdZbzQAVochxYJOA3j03K45wxq4Q2mAHH/V6p/a5yvVc646FnTVckhpXgfx43HE
ol2LtaoDT5gSb+iakJwKJoPLvUFpLHZZxZhVC3y0i/2+RVxyM7lqTvQTQVuntb3P
NGewRTju6vO8c702+MWYzA==
`protect END_PROTECTED
