`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wsb7XlTv78AZEw8GCUxPUg7utQzOMwjZNg0HrS5MdMFB1xNtejHXWi1T1rmGjrgH
mq1Y8d7GKPP+S/5XmfeQJDRTn0OJACuVlNAqiAnrLaNMvTTUETtLM4A0NEJkawuQ
Z3Wi2ZXtmLcN37VaY6QhmxbCO9Y1QHeboVanVXafsUNkGfKwke/hAkgnSKXCaODM
WKqGPSKmVZKdeoN3hX47VnM8uTXpSIODEubuAt/+9JD5gQDur10B5m1J8zpfQyxa
0mT0HEsAt3B4uTWgqsMQVnraABM9eHDlgHSvVKL0fx6SHJDwHQtvRbGN5vbi337y
OPou7bMODjEUkVP3pzcwES4fbQQbAAvsafnxm0uNdoi2ZXliOrQk3x/GKdKP1/g1
9Hq7HtwK9k5bUS0UHwyvRytXaKrxvQCsUQcDIWMvXfk0Rl1qAy2cdpbGRcCGTK//
Fv0XCZxabARApvOY1FqDOBLa+uNR0XQWpGTrTsffM81mhtr/ozq3jIOFa6V1eSl8
Dct2ugUQTKvKYIZK3XBUZpYmcXZ6h/r5WMbKPw4YhEzl+oWf8sy0bW2LMACY0MZ+
bidv9rL5ci7CwSro0u4+i/RZ7LQ6d/puGPBbZODtLRo=
`protect END_PROTECTED
