`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MmAwF+bvUh+jXSD4MJ/DbihP5p9GKKqS3W4MJFzaRt8c7VaTZhCvODyvevc7TSkk
ds7FxScotO6USFztPm037xxGHsyCGJHg+y+T63+ZvaI3IaOZ0LFKWIR2Ff+6cZdP
In6rwPbAZ5rLCzgCWZnrS+6ARC+0qNEx/JTmuSSCATsSeA833MSH6DqcwsaYQ+y+
k7sxvzUW0LTkUyH9G9IWo/rgoybR53K1p5mqvaOo0AktFLXO9yls2w3G4FLPTux5
UL/Mig8e7SN0Xw1FUOzt+k7O/7BtaM/z+n7COhHlqoGsMQMu8dpPJvN+Z6hywFyD
0TnkxKCgFBfKdkz2yMn9EbZO+3vBwl9+U3Dt8MDRJGTs9usjulocCOUJNPKj3n4S
z1M1xl5/Y3QK9IU1Y2dodsntwpzAJXG7JopaeSCTX0lbl5LwvawMvDz77SyWKoGw
0v3YCUUSBJyjSie6p5+S9zDqsyxZRP4EIG19nreGiduonptzwjSKhWHirTywu2MV
hIzDP3mckRzZ/WLZsCAyRLRi1dQwS/cpPTOerszZ3hatQYdAeso+EMZ4B3lEmsLB
rUXIOgB8RJ+82U+Rb+AytmSBazZRwN0gTHnhtTpLCxZZmzisOPu1quPib1NYm7R1
UrFNd/Wgn4IhdHrC8M+VaQ==
`protect END_PROTECTED
