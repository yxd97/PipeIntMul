`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCcboZIAAwJncunmf7oGMaiJSsF07k8XV2tVoAQS/bEHKaXK2Izf4rjxMrMIJOJa
JuOP2fCT6O/N4NFdXn1emMIh3WcFpaPoqVh5j+L18/yuWzbcBF8GEffq3Kuo5YBd
XRnyK9lDSFDebasp7LS6JU6VhwskbWP7OtSRczfN6RidD1BeXwdkYJ8P0nnCKJi2
552TcbvCquLpJGyorAiwTxA5e1gKKRpxazVip/1amAQ1+ErfKa18W2d5hqPg1dSQ
iywwmBWcjlYQZxYb60NpSnhmha8BlqxvmWpUciR4Hk+9kOYQ3MQ3TrWmhIAK1fEN
2CNB7uAzDiLsGkq7b9JuMXd9fhmyV0eOZsxmfJUeGszHROGEX2k6VVh/nUuvOiYX
z7ESjyirxTTbG8hDtVF3NNf0eLA56ljztQTheDG9yDpR+SfCw82GX/xOfkdCCMXc
9pf54SzHZ8rlvgXGnsEmMxsi/CKAfc2olUh/0U07pmI5wofYo3id4s4WUHNbZuIY
5rPOcQBwzX3a7mLK6AsHL5BjWV0ENarCw8zqwiYO5bSrly74oNuCbyugrtO9ax63
WlRw0+tF90ij5WInUuWhCMm1jsEJr1hiLZL3HeGo/dxUvT8fnIlXmknwcloQCofv
4Hrc5jVdnYFmikAfEjhWPi1q4XPzqI0H8XdeENQcRxrRGgbZPtKDmy3z0Uzu7PfG
XfGdN5FeVMRyc9rYOGrXRdBkdbJTg3IIRucDAvkzCdc3DLZVAB9c/21lW71uE2w6
2BC3STPtWmgAHQoEAlBcw3irvvF8+xgW9hw1lnKovxIA5KLDifoWnlabER/ASIy4
84HUtgV83vEKXT0osXo7C9t2WpSR7iF3/u3oRUMa56p9osyiRCWai5f0EIZJeMlU
k3HBe7DePWmjZNmHAOeu3jxl0QtyuRxskXphNIdVKkKvCEQUvly9YG8k16hXMW1G
0QfIfGNua+/bx8+pspLlS1KnWLRF61G+T8t7S/ajk9N0JmELnXYuB6X4+LQFPjLF
H5O1LFTXKT4fcd7IDXOThSZvUE4bBPlXSRWJbk2LQOowM3v03hpGzQ6GoOjUfM+A
PNQs603GNI6lu4XSN7IIj5Fve+WOc43105Gi06oRnPzID23FzQu0pm7ntBgC2beX
WDK9DMRnOw75zyZ9tGY/kaZRKlTB+TQ3/l2yeDErJ3x1biUnQ+U0HETMtOVTPDjT
B1y2aq15/b5VhtrTAvSm9NG0KLrYJ4/DGQRi+WfU2q5kG49fSHkvdi3GyEueIDmh
eW9itFGZFMHVe1kEQGiGAvLugSMxTCCXzCyWgRpSvHH0hYUXT5GEvEwSfmmkdR/c
oqu5roTGrdje98ihpT+xRIwq8XFAmLHbWf9SlqlYZZhb99/GR6CDd0TapjQ5pek4
OJ9xl+b5UCE572b4yRPn3QDxVoWP6tHrW+BeUs20MpWQgtdML16x1+nLm5lluktB
sj2E6dGirGF4mu74V+gL+QmcjBBR0hgB7P67YQhEmZmK8rDfcum/sGOOxl/tqx1g
LW88/BBvgA6V30oQmj0jn2iSSTGCAZIG91qEWdfwPyYV7nQXUseFxFJ16y43Jdnw
Ytl7SdOszFDduBohH/VeioUD/GZb8/wy+XQAHKd7ZVXSFfibvrOEtYkfpDC+zwPs
fOa3K4xe/7S5oeZwjbwgXpubzdhmfYenzSHbInoQkR23rELMNFJWGIGi+01gmsIb
M/Pnot4pD26BbmPl7LCyboFB0Zr5bH4YJD1tgkWqArPs5a2MDi8KzXvYqhKFmmNm
fRbwBhXjb4bWLsQq6LEwofnb42rTGsatMellcjtvk9t94EB00c76vSW6cT3rcV6d
gtyoInovUPCMcaBU7LMEguVPaCrapD73uIcTvHaSifHUgEYLP55zv9jKZ5c4bkAn
l4F6xL98oMhMNqRZQ3Q7YDrYmPeiiLRRBtmJ6f+FD5Ing5ntedx/0BlEmqdP+wJc
cpemcPT8VvJaEq88AGfdm6lHK+1yIz8Qfadh8v4Vrm7IRH8cmt3aEyFH1MO8HYLr
MCt8A3gKELymjBVhKIqRTo+Xu+QvgwFWEir5Z/2ryYVSTYDV+D0vxuCCFYOdICOn
t9sy2PBnBOhFGHUf12VMhT2Rq4bBM3bU691+MCer/oubyAZ8mZx6Z8J1gosMRcEB
I1oEJ5JJUZ139lQS/xRQoHAwyyo3SwpW/HW7EkeYHBlfOVSzWkaKA9IWm/uzgWIA
LojwnyLil0g4DnqA0c4tbhUKyGNN2cKd0XBOwhvtFWYbC+pnOmV+rbIMB2Ezx65S
Bbm4aE92q9GNewzIY2T94V2Mhyv7zAZFBUbbsnd5a+n3qcTihV9i+76C21l12uFj
2VKrJS4aohpbvlDSfgqrHqXm08s+YFWMo5OVVH7R3oo+VpDqFA55+tExtsYMYQEU
oalD+1hlccohsrgqJpOroCucF0gOvzkuxYDo2bkeLt9zhJkRlE8otKWwI8pXEdIR
TE92tVHiXT11rl1Lofzlq6QA8J3gUhrRTIWINw7SKisRIKMbsci++Pc+cD6Ys3uY
i2gpG5C7iu0V4zc/NMockOr1C32d0GQeaTvCe3cUTaSBIt8+sBqL0XqNsI299oyp
rkxqQxdNsmbLK3etv/c1hkN3WLOiHEmfKUeOjS3u9FSrRrTZckKxY+6nIZ3YkDrC
5C3/otL7ISe1Qrsik3uOV1sc/1SXRw6dSrz29vasc5sRyX7qXoluUXOBn02irLLT
KhXX1uYHpaqS4n8vx4Ucj2Pm8AI4YEVQHI9wTqIiswoeyc9Oz8ot34ZYYCkn9OnV
XSAa/uitElI7IC44dIzBldHZXK6191EPXh6MdRATAIRbFYcq3J9Cew7xzrc80+NW
8LaCCFZnigaiErQAYeGtZNCfpip0gxm3ewfhggjmLFkogeYgA0RJ0hL1cI6vulUW
v9b8an3kIcwR68q3SZn7+HlZvfmW7g+K6t3w3vOgS4cfh+e8DwDiRmunfBnDprTT
cMADgfteq9Rn6ZECNhmef3x+ksX8zcc2b8vIGuPTvez+3eaDuhV3Ezi7HUrRcR/1
mgD6O/ZXUuyD7g3QCu+VBrxgHeqvULMaXg1yjb/rYYa0f0nxVpiP3747cAWrUp29
PBo7qvL2y1F8Fz7qNUY0/Akc4a52TLffEMa4WwUyZGeUkk0GruryW3q5+lZ3GAHq
Se892ukz/i1uRB+TCUUQZIRfvcNDQtlBU7RR5aCjfgzJrh57wwbwnK3bi2kbk0NQ
UaXl50L4swklOdjk1OcY3gVjaG61ZtqKPrq+kyx0sBuF7u+zLKZXYtt4bHiZXBvC
sIN/pGKyA3ZQDaDM+TVG58gDGcaMXbjX2N7r/+5Gz291QHF/OZD0Y0gEvFoS6Y2/
AxjLXTTzAE9u76xUkqNs1xBv3T4JJrM2q+Bm+Gv9BY2WjrRvoJm8Os2NlzcDStnR
syyP2HUdhdOXof2CA36ED4dRUWRM09fHbJNJxcPFjKmxHvuJv3uggc/uqO/RFkye
fWetpZbjuGDAZHaHGha6+L+FiMLwa5xHuyVPli4YeFBRIwI4XzXDbiQ9aKQylwE9
Mr8I724a8lsmDREds+c+UCNucHyXDDXuGIvNOuZtyAbCze4x4MUWf+jLlg8b74JE
RjGMrlV0w6HjyG8ZdneXWH5qY5t44KRWO0aTMmidSsgulCy1IhQ7KYaR4HBM0DDq
xYydhOJhnt1XxzQQwTmSapbHbhYFVXO2v+ij7PYX68hqd2DHMX7lcQaNka9gXlsY
eEefEoLjYsgdE//Ua1lN+yLoHxcKm/DNtMrr8SOl8yEqeMypPU1ZwLoRfedjqEPJ
Q26EQ6z9DJH3AM1DRr3gJsKlvpH+TphcKW08erfIMvu9bosnz2oBd6XNylb9HtMu
amY5WUclTqxxdro6Dchaa6VEPcsDwfYTdPRhfFe1FzbJkG7UaCKA4Y1ROnqgDLW0
eysFuY9c86tq3Md520Q1ZLehoWzGFSIbc0pSh77GrRQfsgxdvMKrrYLu2w3IVQW2
eDmgz650HUOfCmvpVh/tenodVd3CvvRGAOBkrI3JbpXvqFGVvII5Im/kdweEFPN1
c7AX8D46fNiGbqd+5jDDEwM+2nZY5eAyVcrOnJ4TjlfSfgYERZfFKTEtYddFNVyZ
PSJxouctDBZIASGcS2hiwCZhtQiUlhM+sy2RDNWhbW+PfQyCeAgzlbyfOB01jfek
gzo9psAzOYHcx/FvoQTXPOy45JbEWyW4mz8ahqp9ne7NQWN9xyAKmPNwiectz88r
dK0up/Ik3w29fQS22fpPQ5eK088ooWTc1k9D4uxpUEmEP+rTIj+ARFiEyGrHmAxa
TVUrZZ8KIV++f7+TPzgleoweLGwpUUTsR9xFNTiWZVR971zvQPRKT5hiNzmdFbiE
jmipE+Nb0I8+2aTDNZDI8/E1PkBWNvjoWJNd73cp6USJxuMy7Ul/qYTkDowJ3h3m
tchU/C8YMY1B65ZBvMsVV16tMsb46MeMemw345rzYuKiBnSV7yrOp+6fPqCvQXbq
RFqCkIX/QZTD2iYtaCBsrmZvjxg3gx6zjxIu1JYHP0FQwMtxPtWWgJ7QVopNnnrR
2yX9iziUOs/jXIDBiz73NS5H2FkaDfHd1uY37YxglHr6SmOQiZxVtRlT4ObprLrO
XUPQl1mmVSYjc0OeNrIGDBbx8oGKt2DmNPGkmerskGFxyNR7+L2wwQnmT6jFnZtE
9MLe4jdA/x02Ca383CP/mr9UFdhIfGitZo3wEVme2K3tmi1xUv+h3g/DXvn4ShB2
ZSSC1SwWP1w/t7cfZPLp12NcB18/3yCS7FEsJb8DeEA5pISLBhVUbTSj2vNP7ed0
1UMsNYh9X67dM/ErxZKmq0gHhf4TQ0whcCu7DjLWRdegVNcXuqJV1yZbwyjlapPh
hrSmqZpQkQfGdp0tK8z5+0wxMmqduR7XUIcs/RcpdJISEGOju07v4HSbLaoD/9+l
WXgOQUM1TsVNNjDIkvDBbgaDVwZ4Lfb4Y3Th8JWJZCyWphdLJL8RWsgtPBv0+XWV
8eHi0YoB84UlMzHmguA0CKkEeD2lzNrVQa3ws8v3yIMdODD6q1HRrzOsP4E3DUL/
BVpYCDkXQcV5MMaBNJsHD1cLj8xCk/8ZOstHdLTMwUViOr0YSdrYK0Cmv6g3xXGS
tC3CkVbf+N5ka3D1NqkebEQGsvxRncjYByzHPpJvl2yO6neGwir1qLT3qFZ+ZcVK
qY/pVxD0g2QgOgKzXgUuEF0q2ah9qYdA3FP41e6sxMjO6w9V7114f78CHXP6Fi5j
QVeDjSKmmZO1XJW5HVh7H6m10Tui1DOY6SJLQiXPrUaQUwHM9jkcl+NFvcQIdtT2
kgutpc8VIVr6PWhZ+E5l3PV0xInYZPEZrSF/RwQMwbITw2txdZc+Jrs9hcMl3l08
Gkp2ZBsSL2qW8UwJjJB4VtfrAnOmIFXLJ6DZ9BlG+G02Ha0omf+G4mc2fV3Z5SVh
8uCkRbio6mhC6g2Vfsz7T8lUYh2c+AJLu/+ROS4SfSWAd9XCLe58Wima70UlcNd0
bAAinXdkd7xweUXVDXy0kWnkBuQ8+uVM73eLfT0DHwL+oujpVgppk8oOm8XRrBfj
g+Wk/8SmNr84jXgotgEyfaQnaSpPMOKCxZ6yGU+fSCn7+Ovvv3ziiwinIgb6zLdu
Ducq9YWtveb2A4vmLFddMfpUo7fTBReFa0w6F6U1YAXsL6s9XLHpslUdK1+c6kJw
yB+5Y24tJtWmisXaRs4pT8b69vLaiocnDf4ALyRT95fVFtVco0A4oBlaNFNRYoe4
TsXI0TcgAcX3jiWt6TZjoVGpQ4Y5KgsAdoXtrDs2YlPjB39ZucI/50ARkj8sBP08
OZY9wJhjcrTg/yeUsgSPtnvCWbwH29xJxtU22KXPO63QA7iwTEcfTgpxbVp7H02d
Tp6lMMVbps9fli78OkFb7Jg/edmWBPQwfzbcKLEZ5bLVFLbhBGm/f2SznC9MEO55
dX7nmXf66SJRNOfyEI0OvxS5eEGfzg3SuZJosZkfUQM8vyJRODu5erqFC+uKEkq3
bFE0EKA7GC4a0mmU3vJKCPIA8IFrPh2sa4qJkXlSiSI1JgAFXI+0Jt1dUZCmHZ9D
LjMH0tu0FkVZa3Rs2nrVRcQI5s7DKhAv9M7FqTah07VW2R7ZHyRCFfBPlcsG8P9g
pac0jOuHD+cRQY4Yb8al9w7W3rlfwVghyPz75QMeH+E4a8fI53uMLc5yATlJiZ3s
PEfNNHotqkALvss2TUiXPrvDnWozsY/++jE0U3T2fke0FOdDz92psYxaYT3UvlUb
2KbeLL1HdnWuJMkU+5aJLPa5EJSRmBX1YtGMRrYI+D/HDjNtZ9zkj8xcqTZPQhLg
SkIZlkb19puVcwPm6ric7tULrPD0xn9VYdWlEVA95h7/5pGam3qhNB3ec2RL8r5r
4ex97S2gfNRavtFhC8f/z/Lu3EuxfQA2MJXK16PDeWhvlyGIDZDhqx7RufjOgr00
Cr+TlewGDBHzAPpyUMP8mvoMF26gUYov+hNn5UlSA9Nz8mDVgPVVaguM0L5q49yF
iFlETq80wlEq6qzuIhKg0xxKXDGnVcjsDs0w6T+ITGy16JXWE2tTCVCHvVOGCi/M
ze6W8elcZKHa3GOKO7i42cGmH92K5fb/+yctiStpgTEuH6KRnUopPQ+PRMOLsF8k
M1LxczTB16sj3EHW36te/VOwldgg0vuWSoAXK7gJQiv0mYih7JyrtuFYEzcaJ+8p
NCKQgG0R6W35vw4SQaCk7iqxI3FRXj5q/MjjtN+92DIdNCWDF1njrM8ya8wEsa57
I+ElqosSvfQ2XvDTRnHGXr9OYBbyAeOMORyWyBDYoR+60SFq/II5AP51bnzBcsG3
yIBGar+Hz9/I71FxjjMmGrAx0y6F7Td1YISEEHD9m1xmJXxSpmAkH8nc/qLQ8E7g
bH0hkeXlr084z3fBQPOWo0jzSGTPUZhuZ3TTf6Qm0aajSqUQPNnwll2fTkoWVBfP
KcyCsExZYX+MN9A2l+l83KHGe38cwmsSe4y+zg0WablEhha0uTx33/pBoMqqoKOX
0BGD9HrDcrpIzpLgMRbmWxSzeY7EIfH8/O+eSdHSGwS9MJa+M5CdOXxH7qjQkTV6
IRk1t0Ov4OXwCUdr0idvnEElZJqwlx9bmO2nQg1wMcW/XIqpXC+Y82E0biF3zPui
pG4ibkzFoZkSp1Hg/6cJIymLmooyVheq8yPaLR1jlohg4K9p8MgJIzQLNlqeKHEh
Y9cYx12s1aOtLgWpTGIZ67HPm/8mva2bpxXCS9kaD2J0LUtnF43NMGp4s4KW3PoH
UcRDFpk3+YS0ixnX5I/g1g8EbD7O8PzwJ81ovvaULxgFchd/y/ql+JOqyr2OvSf+
k7w1R+G8a1HKAxZUejYqp0AvQMmsoX7GXHFqwSNIHu75q1kKYqObLqCOmpjXTK4s
C3HEbnL6lOW1pkv7aeZDSJPcTc7w/UfLT5DGf378cXM=
`protect END_PROTECTED
