library verilog;
use verilog.vl_types.all;
entity X_ISERDES is
    generic(
        BITSLIP_ENABLE  : string  := "FALSE";
        DATA_RATE       : string  := "DDR";
        DATA_WIDTH      : integer := 4;
        INIT_Q1         : vl_logic := Hi0;
        INIT_Q2         : vl_logic := Hi0;
        INIT_Q3         : vl_logic := Hi0;
        INIT_Q4         : vl_logic := Hi0;
        INTERFACE_TYPE  : string  := "MEMORY";
        IOBDELAY        : string  := "NONE";
        IOBDELAY_TYPE   : string  := "DEFAULT";
        IOBDELAY_VALUE  : integer := 0;
        NUM_CE          : integer := 2;
        SERDES_MODE     : string  := "MASTER";
        SIM_DELAY_D     : integer := 0;
        SIM_SETUP_D_CLK : integer := 0;
        SIM_HOLD_D_CLK  : integer := 0;
        SRVAL_Q1        : vl_logic := Hi0;
        SRVAL_Q2        : vl_logic := Hi0;
        SRVAL_Q3        : vl_logic := Hi0;
        SRVAL_Q4        : vl_logic := Hi0;
        LOC             : string  := "UNPLACED";
        SIM_TAPDELAY_VALUE: integer := 75
    );
    port(
        O               : out    vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic;
        Q3              : out    vl_logic;
        Q4              : out    vl_logic;
        Q5              : out    vl_logic;
        Q6              : out    vl_logic;
        SHIFTOUT1       : out    vl_logic;
        SHIFTOUT2       : out    vl_logic;
        BITSLIP         : in     vl_logic;
        CE1             : in     vl_logic;
        CE2             : in     vl_logic;
        CLK             : in     vl_logic;
        CLKDIV          : in     vl_logic;
        D               : in     vl_logic;
        DLYCE           : in     vl_logic;
        DLYINC          : in     vl_logic;
        DLYRST          : in     vl_logic;
        OCLK            : in     vl_logic;
        REV             : in     vl_logic;
        SHIFTIN1        : in     vl_logic;
        SHIFTIN2        : in     vl_logic;
        SR              : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BITSLIP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of DATA_RATE : constant is 1;
    attribute mti_svvh_generic_type of DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of INIT_Q1 : constant is 1;
    attribute mti_svvh_generic_type of INIT_Q2 : constant is 1;
    attribute mti_svvh_generic_type of INIT_Q3 : constant is 1;
    attribute mti_svvh_generic_type of INIT_Q4 : constant is 1;
    attribute mti_svvh_generic_type of INTERFACE_TYPE : constant is 1;
    attribute mti_svvh_generic_type of IOBDELAY : constant is 1;
    attribute mti_svvh_generic_type of IOBDELAY_TYPE : constant is 1;
    attribute mti_svvh_generic_type of IOBDELAY_VALUE : constant is 2;
    attribute mti_svvh_generic_type of NUM_CE : constant is 2;
    attribute mti_svvh_generic_type of SERDES_MODE : constant is 1;
    attribute mti_svvh_generic_type of SIM_DELAY_D : constant is 2;
    attribute mti_svvh_generic_type of SIM_SETUP_D_CLK : constant is 2;
    attribute mti_svvh_generic_type of SIM_HOLD_D_CLK : constant is 2;
    attribute mti_svvh_generic_type of SRVAL_Q1 : constant is 1;
    attribute mti_svvh_generic_type of SRVAL_Q2 : constant is 1;
    attribute mti_svvh_generic_type of SRVAL_Q3 : constant is 1;
    attribute mti_svvh_generic_type of SRVAL_Q4 : constant is 1;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of SIM_TAPDELAY_VALUE : constant is 2;
end X_ISERDES;
