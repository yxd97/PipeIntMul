`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5pV0Jc+PmN1klFu3ztMxkK4IZrAL674G3n9Vuqrj4Zt/V0sv045Yr4LmxBrwjnYI
qj9xesHdzn4K9IdewqHDY2J3I7rmHvOYSgoQaht1k3+RC/b8OXKb2y1lbXtRI+6I
xgX2NJoHPl6WYjASxGzSlk9YO74aLm7f7SIkTDdp4NmXsJSN5eiU4Kcmuu3tQUea
jOKlhPq97AB5bb9es3fX1EQLPp4DZug1nTqJUehqViN5ViRg8Zx6c9lQ5icLpAXh
iQdwqooxemq00yCVpZLRaCnVX9p6okUfO477fcEJA5qJxVoyw54g8WRsLx9QUjKC
S1HufOTPa1Hp9V6c0u9zqwkca4TxMLboKEXaXiCO/Sk+m01ufDwC+WQV4xS4NeSq
Oo3iK9GUfhaMy8cK79fw1Dw7QwvTAQa50Wp5MFH1eVuGm84lxF9N1fX7aKBAB+wo
TE4oi3y1VBoj74OapJ1OcIxJCRZekofjRtIjyfLvVeVovloii3y4PTvlU1nLLGK0
tPeBVV5Ye2UEoy6aVffXDV9JpRPt9nvOWyvjcJSWTrhzVAB4sesoedgqmBSkPLC1
fhiimG1Ek0B6uQ8yIlH1bo2NC62MZSZBAtyXKuAGd/YetMnsq5h4tA+g+RxkgcTt
3inuFzUxASphtW9JQFTSLnnJUa2L6pRQtLrhtrcvVcZfqhKHdD32iSAnHQYDoUIy
UmskJz9K30X5KoJt52jthgcRmlkPmVM8qKtnTSSIyU7gn7mC67E5pD8pqOejCjoF
RAR8hyRIQU82M4j7PqOLipXfxudyf+GS3a8epBwSxfQtP2LuoimsUTssHfR0xXjP
2/NQQjrTf8UddG2z+jMFjWTIfUgacNSMtFgf6mJIezUFL+4EmljKZ336yG0TCiys
POSTLKguyG6rC0BtcrMwsHSo/d853eUrZh9K+/O8XNxrlw2AyEm/RhWGt4lweQWy
kUMZQt6gasSH4cxccI23Eqc/r20oteCkLBYW/1VIJdYCP9tX//QpjP0KDrRUNbUc
QrGPpLb56y7q60CCwUhWDVSIUMIQtODxukpUNnS+RnaTJ1BWud6pAaIieJCM2IOV
oLUSieURp7eYctQf6zlvIbbx+Zv5wHD73qdpTuHpMsbvYWXiaovYD/yhv+W0tF1T
+l8fPNSbgjodcqzRREJ4/ZerH00/uQybZrSivVIkj1HVWiJ5HycMUqBmXfYYc97S
eKyjdi8hkLqC40Tl0UqqBUWD0VIz10gjoqMZtW0RlDj65Nn47rGIn6SLHU+IYr5X
RDq2IYC3nehCuI8O3vJ4ErGcb5oATgdvnz9dbObA9MfgLqn8DtKSvs8jsuaQmSTm
hlIACLscqccRpEcR5pTPfuC3PzuHgKCFSYc7b/036vdbgGhrl0H9F1cHQotTHKyv
qegok6fGLJ3eEFVOXJ+TjqA9pgCIFYocyqCLaRyneFSGm0dfCryhAUAVMur33jbk
XOH//dAF08OcCDykdA2ZdC0C0anvTbVd0KvyXyqiHz8G98PynPvMPe1Q8In4SCXC
ntveSUcKkbadBCFFjWPfBLk7tslshGJZx7KNJ3jq/3bmw3h6ZfJsrG064jcQ63tL
UwTJ+iCt9tjkiAjjwTgEHX+Fjr5+0JeFhNq1WKZFb0Ts1eyclY4hs0rD/U2ElmB3
nri2/VQKmTBTSQsgg/l5qNG3P4jMSDGlbTGHB0pygeabXPO8pWfKJhSFOhP690+R
Ghi6hozD1jSO0OZzv3XvyyxZQXz3s6sFkJdBEeVIqjtuWGVrSwxTWjUXVrckEMZC
UOUb5Zz4/UhXFU8OvKTpjrqg3EBMYnLhwQ4r1slTeQCrFvkHwjXod37N58poImer
lhIioCbYWj1PCKcM80IY17DS/L0Tdklusxb+kObSo37h6yHDNMdla5EzMOPBzCyZ
35SmxnF8Ic+rA6Q3M2Z5SolHabKblDT0lBNfwYIIAMqXfYogWoXLgIUeE7irhdQr
i5c86beR0nE5MgFxe7rKzkkqZG6FrJHWa5vj4DQ15ZE+wqe9NDLeccen8L0YEm0E
0eRiu07NjMZfy6r9ho1gJJQTgYQXL1TWavE3e7ukMYHNPKnL4vyougBZgdPcWY2O
anZ9llVsTL1KDVACE8ohrv/TIk7Tz2kKQuI2jwgxhAht7ywQIY0qgbeZp9AgCnc4
UeVTmb+IVde38C6ZdAeuRxNAV3nq/BHij4/uW7Q0vZqvgp8Qc3q8tXzNYtvfwCpg
wqsl70kxq4QPiCAO0REh/tkMUkk2qXwDYxY10bXorYUYN0lzNGe60VEg6CPUqJyp
QRMegXrVPKdyH0HrfNsU5y8ZNorrSdsO8fukj6fQaKgz4fpAbyEiWZJxrh7yTfpf
VAIWuK0Hz7Ruj7j5w4lzTK7Qbp+FU8Irml26pWOMX9aZr8Yc2OcDYs7ejvV3u0UZ
dR8O/EQ6idjXkEPcR+lA/Zr3eGvpVUokmgrmfK28FK+rTNPcY2LX0zcpJ9m0QjPr
B8W2NqfAQjdsD6nj36PCLlNgWv4I9k0oVMBPE/PVJZYKa/JTmFQtaNldJc5TaDWo
2rv8MhWoqaZOKYq5OsGyogBDz1/yNIm+Us+6He4hqMvdFebXCx0xsXFjFzUWYEL1
3ibP0eNbCHceMuX6npcMkJQ3WA5kzg36e3xvdpoUdRRAWkNv+MiQR0MtQyPANFKN
e0P+33ucwDCyrgJL16OxDuR2TSxcoxweMHG3vhQJUw+bQEsFBxinbalT6TZxABoR
jbojNzRqRilMh0BNkYC3uwba/+Yis4oj4IszZDd4x0zLS3z7eKczaqlTroFyUKHD
v1kqbRphqYmMfRthp4wOp9z0u18ExkzSQQ7jhNsqsq1r6vdUj6FB4t5PP4UwHxpF
B8Cz8VmAUObf+T+wxO2BEVbfLhnJqEOvCNkPPCOO9SVyIkIlXvmdxazl8QJIlmuS
cXUOshF/rcuaXprKI390cHmjd4eCJR8kZeDNEQMOR35LwXycpxphj4KBt2cYwvlV
OWfNgmtEHstWB9EdMv+UKoDkTZgpMs7sWbXpjT9w6bw3CuUi3wmy8IV4agqIuAv0
2rgaKwgNPsowvEJdLpH/IM815EiRj9ieP5jz35FH4DPf+3+WoPkAo/gIynXbKolv
KtLi0h49r3My77/qcCWvfNogTSo9usLjvNR1eV6/UNQwR6uf0t5kLHACShwEaN/m
kvzOVt6qB89P7ZfgN01rPI53jzrT8ZQlW5Cg/2K/1Ki7zlCfpbnEyAvkXc1djz+I
7e1wVA6P6fUo4301KzSacyzt3Bw29TTLewxE6eHCBrUr7f8ZDnnrC2lWcc/Bju7h
KwuMgjTXsld+5/E0JDX3R7ipvKAmWw5mzHLXtcoD7t2h1KgQ8oE2Gg205Lf638wz
1TqDAFk022nUJB21iA5iIY6raC7ucthLr9GeDZpY2iEr8vqBV/acz7UsHwqoMWa8
Aa0tZc4pAGBkKM8jOvbDiFZSanUYsjsFahgp4/A4jKdUjd13ooJKYTDFXmZXltWs
1ka7I6ve0o2b9ALzlePfQ4nPkUbxsl44twSjIoasFU3wpIxdrpjgzms+BgvVpmNN
4NVCTdTQs+WVMGv79t+GtymOqTGuu1A6OTi3s2V0An+0VYpN0nzji3PKbm689XJy
DaXSyPdShapD/MhtAHvZm0FWNwBGdeMCJxFPhSmCGgU3A5adSUj6+vKsGynlU52e
9dd8U53R5YUjXIQWjVdw83zShsPimojk8WCD+2HN0QBPAaGHj89JtUmy+NTuLW69
ARWYJ7mpF8g3163IS7gWmYmlbKZwPqtyLDcz4y0MaOleXjrXasbzwdJNpDhZkXwg
CD8GbghXcMFS4mL1RzDn0+gImhdhC13ubLgUQt5PQq+WztHujgSVcmqQsgHXfpe/
EtczztZBLGVPdlC/JBH9X3AoKQEldCFn/qHiPif9gg/4LN5z7QCo+guljnEbkIOx
nD2oQ+lkD6unyqY2NPkGCFMUEtfiYpqNouasOW22ljglsH6/6NPZ78fWsKiTwYdo
Ulgeo5WKHYRslUVxn3hAOuPw5UNy49N/7NpPsX6/qIi12o2xBxD3+fb45MWzFVU5
1xgHKxmlv1SJM3QRb6VfFAUxjzAdbyTOPjE47nYv6mvY/4Tm6DEG9or4JC7X8W4U
6TtW+7hXg1J+Kw7qcDOu+C2zqjhVWYyM2zYnHqtw6X0B6lsXAYdUM7p1ZuRwDS27
DcE9iI+4UWfr075IAlB1wVnpe+30axNKAT9JC3yDBM6mvUBu7D1idlw2nlGFx31d
diODdU1pb4dFi/atPSTv/loNc0vsvft/Q45yOESBHQ47UO8ORjGfMe9bDnnbu5qT
YYceqfuRsxpATFC/iE/78oLddNEJdAQV9K7iUvj8+/NZj+4t3YKXqnXRaQczax/+
lnBmGpL1LVrUcBGBF16IuZwgab1Mwb24DBWJYB5UYn5wfGbqfQUQQQjaXtVStePQ
x6p75oOIBf+58l5/VR5M3vJBSJ/5MGHkrINE/IcvEAxhkeThrcJr+Ur41glyhZmX
uyUitQho+w/nVdsGji3MlH/39iASO5Nj23OI+Sw4u7VOjh4RJIB8U2BqhS9vN/Cu
EJo6hbY3q6OtxsdVuDGiy3jmvUxt/rAh2LiRW49whqvAIYRB/jC5DsR+cmhTjXne
yV7vP2zPvHw/Sjvojp2Tj6KAZqAO2uGX6AgbtqlCXE1wmoRgttjUYg/5uD5Pup6B
+woChoz8LNrOQT+0JAxi43Ofg7p2Kk3A1IrG+A8m22jWQIhrt0RzxXHUyt4w3LcI
JtFb2/OhjWzbD6/OMHV8PUHM50RrPvM+1EXgN4/cwd8DrSefANOW9skJkDfdmx/z
hj3BbKuSKhrhE9PUZDNgsWrrQqvZtEZxVTuPfBfkoTNBSfm9khPtK7OnP42CKXsC
QJgLvEiUGicKOaVOspwY+UN33nYW1JRlDdbJpOEVD+lVyavsFv+vo8laobKw4VJt
5JgYJjfVzz9VPw/pXqeV4FNuUTfs3yzpBNfxsisr2qxJoLUfBkvyYYvegm/t30IL
Kx/auh9O/Vpwpjl84GIEwK/4lRnqoPtfum2rX95HZMCbdp/PrazbNZhoeVTAverh
T1E8gYLW/fL9y4fPT/f+KRyr6SUIUBhGFQYwhnDMWFNnQ7V0nx6G4sAC+zdp179R
dmgvnx7/ZwZEvWyTWxdVtgaJu6/hfIAFbTA4d7P0pL51EETd+pnQKrcmqmn4TpSs
l/uS/C4ibr8cLYQDrhaCDyRu23sqqCTJpgY3fP30sBOjL2gX/V2iqrkP3oH8SJ4M
uvn2dwK3HpQFBjAc5EkCND6/e2WcT0oj1XJVH5/lUJ4=
`protect END_PROTECTED
