`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X84vI4ORFYiFnn4OcqQ7ICF0BpjsRMc4w9FS1nlogqPLLsBGBRWkcstTqY7m0MUq
zbAvCP/WVop8pXZTgxC1HukmOWkPyChPGvyaFFzJFgpRcB/0WT5X0JLCiTBOx9xq
ctHlFDuOyczAYoZqXt8OJvRLAXuNEM6dtnzU3wfaxvJT6DNK3OsSKD0DmYeOsvbB
RoYhtFZtdRaGqWK2uCN+2dlQuR1drI9XAGpLUKN+mGOlDyQUbthwvD7mGi2ncjCd
2CDp8K8RqL9cXO59A9i3MangmiD5eiOOtWzVmreb/USBD2TWbfKJUO0y2lJzzw4s
Kx/fPDfUucjwQOWdVWPWzwwKlqztMVHrvCpUjBwcYue2DUYVYzLlMPQWCCz2xgmy
KUkHg/ZbvkELp3bQb3zY3hPf9w22Y2himalDDy6WuAaOZOZZAvEmIYiKi8O4rkxL
2sYWz+ffEggUi7rEjMdaYj5Hou4hNY5hHJAjb3jAzxQGGUg5VwY056wdcRUKui9S
no9dZsu12vH7oWkdcKz+C92qZ46mRH7L76vAepQd7Vbrnd21DBgoxHKVTRk60S2y
`protect END_PROTECTED
