`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2VAiN7mCakC++xOF6QBmfxAkU0b3p0KKMSEzKUtZDSABbee9XekoZCRfU2/4jx2V
/B/mP+dHeSUf4bWpx7Y/gp5TbCFQOsRWJCPA9ePRgRVfqAr4e8sktQKUVk4j4SgZ
eTLgVJBKOQIH/X9BLKn30P3FX+QNgAGxTTZRZ/eCZabxDqiuLLAd1M7LVMBujIs3
3wtWCF1TgLy0lV5yfeCZddg1wgFo0zc5dTdbUcAAHqYOOEGD02Zfeo/XUDlM9ieb
1Ec+8h9WVrr8knYLsPCc9II9VdPzpDvTK6wWN+BKdq5mqYWBEY7oMF41WO7sx9vV
aBBRS6vEaBJrrYWDLLSvyx7bUbBgH5Jfi1Qb2nr9z2z6Noi8eBU0PHdIaHC6veq7
edVTOv8mFGRHVaLL0XyUnZV0MiLDc66/M7e8QQsy+x4/bQq7m9lQqpxCZcpq8TfD
BZDFW+gfrW6J8/RJMT8uWEZ3ZcQYA40AxkigZX00Wosr6VAOeqKvGs71JoSCE7Rb
Iw0YSveFfn+ZS2TMwniyAsuEUTpefaJTUVoRZ1h97IPE4E4m5BE50TylnWBP9wyL
xbgFaaIG26aUlajl/z5u8uy6dIJJLWBvRZNlFYrrskE4d4A5MpKF80ELGDIg6Hpd
qLF/2AWuZqZvWy1yPbO9+jQSj2YOgwSo64t4CWwJ+Q1XfT4+IdGc2CuIMnT5atI/
hlZS/r/5/DFs1p+qzR8cRQNJYf68ld9RjuHHYPQQ0dWMCRZbjcpNbB6/GRh1TGOl
kXM6E2+LaZAHEAAGsoS2xHoZAyROtn7y/KwdtFVfddhRCaF+c9bxcs6vbeijbw7t
UxjYfmRDyd892rF0SDRgmW7k28iSnjJEQqruiJDbjtGqXnCtGF3llvgu6WAHZzLj
3aYoZ50s+H+8z4HWe9GhiciJPkkq+8Bg8+HmySt1hYfAA/0NaqU1bTiT/b9+kM0K
jEXC8LVx1PJ1/5XNgSAxYXSIOsrSf3SXoZYz8EdFYkNLVCMGtoKX/UeOu19MJbMG
0jhX3FUheV6HKmUV8cNIl9u7BNAnFAW/hHqkViMd5m+DgQVaK2lIxEMBmcsZKt7u
zDjFGcaIe3iuvlZUn5eUgHvPI4H/kiEUCCgc7KrfKUsd0qefO+nuHS2e7xqBsslC
wSviYTgb08IItijSV7IXjuW61LYkGMzyByNq3CZmSly/cCgmmmGLlDcFaGtTOlU4
OyoHVWvgM8NZTDkJShQlCih1bOxWTunjY14cp6uVbg4=
`protect END_PROTECTED
