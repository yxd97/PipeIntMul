`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hU+DlTasmRDe7dktH3fke3p3mhc4jrJZryfBVqnaOUOeBV6SLXw9x0g3E//S/zsd
IRtWWA8ijHLr2HhSzoWkQoAbGWBG75QdvQvw/9nVkFYgaBjIbDdMa4ciPpN7MSx7
1O6H5N0bbrmS8dXQ5cTzNnz3MUmAHojup8a5sJ9Spki3SmS1gof5YqtVlkSapm8k
cFY44zdtzKGV7ocvEYkZxVwlnxvBYuvJrWgn5N9M3eMFthyXjtj8kuT5gTQKjun/
rBkOS5KoJG+X8XD+teuxoNtlcdbFZAubAfnfq2b/boOyCoWQU5lKFlhwfvBX41FT
PXVXqOAV6EgYjJDdur+iwyXH+cEvndBN+Dci0/rkumcF1PaBg/uitTFP2ythOzYd
w7iM0qJzv/uGoM6cC6bKspSCRcsVFlXDHItSSE0ezYw=
`protect END_PROTECTED
