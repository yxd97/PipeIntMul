`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XWxDL2QTutfUdiKO8iyslLxDHZDkPzie7sX+UVPDVnPOUDIpslWlPGfGXEkQwOCC
Bc75vFxz+z0Z7QNn+YNY2qv3a9P8rM+asx2Dh6zREKJaS5P2kTt9AZoneGOef1Hs
orhXGSA8duGzi5uN4WXGJ/POSwa/k7SanOpZOFN+5gtON0ORHmUYUJxaL5FB1kNT
0YOhsFQlawIZYGpzuRXq1ZRv1pE0WNEe6Qr2izf6l6/c23TCc1oxUi63H3gswKkx
hICm0UJYIDo5hSJoh/yMyofViM1ar4VjOtmxamD4vJQ=
`protect END_PROTECTED
