`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZvxwiLPrE41sG4B2PzaTYpOMtV5Z9T0dtxUcvO8zAUfk5BvjtLvLGDSL440Q165B
ibxax5BO5PPnVkVoKRncSFCXErY/Mhji/sCkZiS/C0BJvgVFuZZ6kLnaAHkB/SrO
nJ8c15Y3PcBp9MJCgiFexfBUK4mGDRQp/UPHA5CMIAvob7XLFM9VfZw3oXEinM/i
Be+iMMGa6wTnMJT6mp7tz4PmLFXJzqO6FkKichItdNsSqQiOPh1ULDXIc9yKCW3o
9VGzZKGyKbAMxEP5zSHOt4SNcJnkCo+XW47DF0mnIioRNd1pXiakQ8VDZLYBY9ou
Q6gGPPTctgjp1ZDieVMtsRnSUwvHnCZlB05+37vjB/8BQNq1YQRgbA66XWUbPGdd
bPiKmc6htdbwBtAemKUNNyUrRUZmO0I+1laWoEx4jc+vGLfWHXqCIjWV6LPdRspF
BklkKwCSTzItEMy9FB1CRkcuTyVzqqFzfGaoe1KQwnD7U1i8CVbZS//K7prpom7u
HcsZiYKm/lZNHcHtkKj19f4C9gxa4gKcbRGiX0zGMalOT4jeSFoCz1e2SuP5XZqL
d2DZ/CxLIEhGirTnihX8/P/GY38JXBrNaO614BO4fWyhBnOo//+JrylAVTj06zJy
wRg75RH4GuDTqGNX9Fq4etlBpoL6PIedKOQhPf15xux1nnJrJOnS6Pscjxbq5QQU
GoHuomsuVR3xYq/L0jMJNqUlrSkfOO9at+tjyDEiZQ+dglZ2zmAlXqrvHJvZ5oaE
bjNRdESY1eu0MSkYE0f7FZs1e3jst04yS1npOjTDm0tbu27A2RZuEfQN8+nSaJsg
xuxLwwlAJOGYu5R6+aL1aqt42JyAj0PFPsBCylHrml/jcAhBMn+JeuxqcnVhmOkU
eY/fduN8XUaBOVfN680C3y2t9dnvEJOq667DDpuCCT87ysNgaHuqnwPtPYZyYSN5
U9oGUXjzXE0tN28PNA74wAiJvUuAc2CvdIyV17XUXiLv+j/wtniQ9P8+F09Ryam9
frXGsSnHsR3dQTyUY6wm4mAQYY5sbVMAuu4Xxe/tONJqJkiinicax8d0pJsby66X
1THKfIH+UfKG1LsqP74sjMcGOjVNMLwt08dGekbFzo5LAF/SBci7JHC2k9XPH+ar
zqVJhPBSbmUeSVD12v1pqAUGLnQen5zBgiwW+3D2ESGbSeXOW+B/lQmKGe7jdzxG
`protect END_PROTECTED
