`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Er8d/V6Losv8tk4s6Suii2G5bbiZerd4O68G/8s8a2VwTChbn3wCUmn66fLvLev
WdJZCbp/u0arlNQB5zVlR9rPxq0An0EODTYSAAMwNSHB9AEwt4Zw7IV7ktt1hKV2
BmvCVDdxEpzfy/0YutqfqGLGqFrtDjGWHhDh0afAjKRDenmNZx5uNiMiTJNtlTEJ
M0FCyw6UITEk7BWYdYIVTO0j4wIjWg4D1ZVzAktfsV9XtFX6I0P45P73ZQsslvKx
BorqtSA+AScHCY+q4h/gOg==
`protect END_PROTECTED
