`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73bv5TWi9NNHII01sZGjofW51CyR4O87wa5YmHCtEEg/Fd7WcqPQVqxg4buvVbGq
JTx+WTd1BSzGN79aEIT221itNkAHt7gtBFeXNvz2XXnt35zPnGczjXUL6+KVaAKi
TDsr5NiIF023UkZ9VAMKEVZ8wPEPSLjBE/NadFfuaiVKYCGOyn28p7zbldWtVZoR
zKQNJTbUhbFEDreilRj1i22azTwZINrTJZ/i2aP84N9wxKnFlGmT5pQI5T4FKLwu
doHMg2y0qTz1OKVv+qrLcxWraE7yj7pVSDZFOOivCYJFDgAGpIZDjFACrrJ2vdJV
T80EIGPgg/UuIByusY9IX7LpwsCc09A4UEQQRMdQIx1nTj0W+Hu77u+Tv86CgkkI
VulVBfG3vP8iqF2+OqbTe8owbBW/mo0qmOkt4X3J0US1aV0yuAtI0Vjzt3awDznZ
lT8dbBiL5UIhF81mnzywKdHVG68nQ5K8MKOMEypWjMZ50Ob3kkCO5HFyk/fUk/bE
SPbVoXg8vsxCOMBycz33uC5PRTZGMTt0yYCJOMyMOZIPO3qD6S/hPts/S4wu2eos
8C+URIOzQ1z5iy7KnZ7to88hCYqXlQHalTWABdkO1sHNW5f3fmrkmfmOMEsXuqKk
pw3D1j0l53P/+6+iJI5cKdLLmFq7QH9mSfDL8CWmSmhry57gPN6Snt4gL4UfWflm
fo7MBi9rCKytZCF1fIU3+UM6+yJU+sct1Xp4x/fk0sGQfRRSrRyV3hSFT8T7LWKL
kWl7eViUwbTZpGhR4EwAa6rc6eKrXTLpff+4eRTrn7BLCuEMLOdOrHZJmCtFfMlC
v9+D5GJAU570kA2re1z3Dg+0s4rpwF7YngrxqJjN5mbe/j4nNaBAYUZmmNXJthVM
g3rk2VfC4SwACDN3b6vQCLhiBoKuOQeoN2fqd18Ox7R2lXnA6S+3yId3OuULfc4i
DauIvYtLbFK0DhUuHPzCdRtvQmcE1IuCO0XxXjVt/46lPzLE0ZFi+QciD8ghZxXy
1TH2el5rtdRxrwLWe9NWdBi1ZG4EtUN2eVTEchSKe0RMQIOkRb2ylT2a5Larg2kO
gyjjG9ZGPMcrcowcTWHFi/bVbOHglFDtSekCEO0j0Ja6T1ozDyIU0S6vhCmUGeni
L/k7g0Z3Bv+day8Fm7Uk2g2gim0HPK6ZNi0hyDWbZiitObh1/qHC1yv3Y2OkfP9W
WuCMcsojOCtWzFFUGcWvPsgcMvxCuM6Yv91BDhmYTf61t6z6JhGy+A7Gd/AajkBY
bq4NzflAiCp/8LdTpPKuJr7PX/iV+LtKSr5NY5Di4KfgyQ/JyqDbG7NORHPXk0XS
f5mnQf6UgKrLIsISSQScIc70ijH5rxvB5HhkF4638ym8xjP/S4LVQ/0xcP/DJA5I
wsf4MUA86jmbYUCGRv3BmcpNpovUCxi15brVj119XrjjyIpSDAZUiJWspXn5Febv
PtGeQOC0zKh+zMLP1X/Rl9dpUgO/ZL9wmJ5l7nvlW/vkkI/fokgy2cLY9Z0HA1bT
dcpH+sb/5MebucnWwMEZ5eukeV070BxSCU6cePcSW35iwCzlMqzAYUdjV3Q0SJdZ
ECkXBQzN1P+ayjAR3BT4OZeyJzT4TCtbIai9s8uMvx505+sCwjQRGn/GJ73+/Bzk
eZrZP3kVO2kL9XS5QZSzOnpeHOcnZLS1bzgb5RgAuqFXc7RSjRcE+x5jSfXfhpPo
YxLJVunrU2QbCP6wuRSZQtXyz3FMGd9HfgfN1SfuLJzxiyIYBhM9soHJbFk8xD8+
SvFG/TGtpZUWsjF+mfZp1/vSNk58oAwzgG9vnyc97AmUpBzC2+ABUvS8fkPX1JEN
ah6DdxP/J5tg6QD0Ha0WnAJsRWfcvX/VGo84+0BQ2taqho+VOZ7BKS20nHRe5dZf
o6nuBqs/R5U1V5c14fD9dPDcwavA2r3XhY3ghMPOuMOfETv/rjfpjPgsdcgM/9qh
E/npHoulyrS57o8O+CVkwiFryhCbnmxeWa/o0/sp2TLCkR0RVN75X7LWKOMZAvdC
uHH3zzjCbbAUb5PHXt0mI3IBl9GrQU1cKBIN0lLixikRGlv/+ZNrPeUfcJWD1JzV
dLsT8inhRzlJfmRntKwX9t5e77Go408+BxreOjrKWn3VMNBAL+CwZ70wcLPQBidW
J1IbnUtLovIOVWefuDr8TWNntVUfc+3ZgObNVF518m4tn+cQjIz+bY0X+uZwtdWi
3CDSFaZylKoo5sSXCzbWGGRLz62RH+T635MjtoBicjs=
`protect END_PROTECTED
