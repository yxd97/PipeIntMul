`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ocYqIm0C+VY3tlR3apBX6ObmoNXRmjf/x3jPScqzbF5+hjVsPmz4Ka9i0GLubUc8
DtcTbX6FvwPp3SNdpe3tUtQ6F7NnnRIXomnPOMWJZoFFwLPXmz6i8Nk8c2gDJKQa
axNXA/etbgofehGXOriw+xSlzz/C0SKI6rULyo4OnyFmP1g2O2ar8r9EQzVFvmyM
sDlcS+7PJq+2CUHgtplmcPOXTcxdvI6ihi6+fVguL41qe/MPY1AvI4guvf6Ok2du
NVqToz/co7cpGquWJs+P2ePaJAUF7YzfzgJl7+9V+JmD30oCzCKRjYGhsdXq4h31
5EAYLgGzTgRcACqNNDZu0A==
`protect END_PROTECTED
