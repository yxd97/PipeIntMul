`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hKpwx1QlqojLDSbORv8G4UYa6f0a/eC/OF5flwC27o5EsVM6yxMb394XsixhBqrj
jmcQJwqt2icwLLIyz4UVZ50t2UQPwOen5mbbg4faNrpdWVeJZ1c1jJZ6DLqIQTZc
3EMwmv6uWWM4SYIv3RDBaxpitEVeyvw1xQPaoIdRi5yVLsy39J83ReAn5/bIGoZa
adxkqGkpSRRvZ7W3ySizvV3yIWP6MEmQNcPJIRlUZzfAD82b7FFFhNtEYQEiGHAi
hLGaScPaYozPx6qh3DsayVnse0iZlbBTI43QvttAdoX+OROjqI78Rxv2wgJutywX
MfjvU+NRjVGewEeZMbOSaE4fenVHCWUQ6qlq3MmL2pdTVw7GwKCCUd7wQkhM7vW6
rCufZRdv5CeNS47HDTKBVWjhQ/JlOw2MY4KKgwTBASwgBmVQxz2k7G+7oY7wlSD8
5XdnxShz8dhChpSrPqpCEueBojdtU/OAtCuonMS8wH4OWZdRA4KJpR8zbriMEpNg
qipKgnlFVMqeyxJFl8xZPm6aMelPQ5FkP1+8UhCvHiEgUE0D57UKO647Z2TlELq3
l+eQKx3jbkvzJ1DHxcNO0RLC9Wwyxx0YqfXHRqJiyxN+hhQYi1PBaIVkFSTKU2bo
Jt+LyZKFjUcHQHBNWMvW7QscqelqlvS90a20zf3kPzHCehgchcTGIybmICLYHQSI
ZNd+MjIuFusxHZjhpGWVRpA8sRFkyS8BfOR2ETXiqPfiGmQq0MgJxK05qkcsynW/
v95nR8MkvLtGHiMVGxYrc02uW8/fJALpqgAwtvCtAN9pBk0gwyJ+VivJcQT9002v
Ll9QFZFELA4EQ4CVS5pdxADttRe+9GQuOuQCfehp2zo=
`protect END_PROTECTED
