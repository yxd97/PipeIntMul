`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PH24YwlEFNb+dJNf0MumxIyemEvhfVUwLfDQVGUZ30M1EOz/kk5rdcA+ZY+gB0LD
h9uJR0ST/0wwEnkSBVbvNxNAJ6uriTt0jDGfGv10zHeqqotzv74WZDqhdhyi00As
+Znp4J60MhO+IkvxqzqcFUunuI5nDSKzKmNxReq4nntsBi2AX4LqFPjPyGrPM5P2
ZQUwVUwRwk9dnZZ48WugGFcZi7TpATN56mSfndfTfgFVZwGSSOihocBKqcbKi7EZ
W5n1e2KLE145IF1R0ZhFAhlwIuD8ZfPflUKNbH53Sbw0MuxQDXxO80vZF30VvJlI
wn2Y8Fn4TC+0pQzKlixuVAjRM15O/NohFrHCiAvKIEPICbCEAGFKsSjA88BI4gdP
rD3XhTp0sjQhoILqea2Yv3phklziO1b3rOMmWpDCr0uOr4i4IIFqihj7hW+SITih
FHNKRu0Crws5U+H4z3BQg3oJ3LoR4g1C9XW/eeRtw7MHg/03+nII5Kz4CPNGp1hS
KPmQPlRjUJFNsN79jsaVWeqS6IzVyHvCCAxc6e9LkqJH/LV1NKT7tfGNLrwHDqDL
sTgAOzydNTgdHOOMsuxDpOyZeZfoCXaHsK2CuihIQJ+QJ+x5eVbeImF0sB0ASNQz
0jAbWFhPPzwUxrBg9mduag8TB4UkJA9kF0M7/siva2HygimUxX4kJBdVclu/DOBL
wBDr6M5f3opCqoXHPvWBA8tGWpLqKN91sj5THvmCbj2ItsvSp1EtlWW7n5tOfoBb
ELmY+Jz/O+xnvpmCyfkMVYe6DtAW4XfBzX8DskStDx6cjxV+HIzUYgqggTKw1qul
F5n0q5A+wCs9JfC8kdGbL5wkCPHH5T2e0TNscoZzSFlGfDWuFDY/WxzTvEkEh9yf
nutoYLbPaIcpMJeRw5Oav1/Cbpc0wL8/8jXYrRvv/3IFKU9878hM/Bz82y4eFR2P
1diqKCzKt9LIGN9W21gg0ukjUb9SoxXfX09twyt/nzJkxa4gOA64EQQ+3WuOjQeL
v3jDMJxx7Z0fTwmxvsXdPTtnRviVi/Mdyp9YPCQwSRHraZ/Qy/f1Ib4soIaKMMS4
J2uGgTz38rZnoeYgLZVLkUFTyZZUvN2y/7HwUu0I3k24Hb5EF5b7QXloaob/jNs/
9kZevJ2HBWLNMMQ0HyFqVOyr2TeyWUWyv6Kid1QyRz886ZoiV+kqy/o2xQR+If80
lbVPrKUz1qtpcgK7oiol5jxN4wl47gPGOfIqYzoM6pDZO/ukxJlBK+zjav1Q7n8O
yWvdWawqa/0HQ4U0yPVKL1dVqcf0dWNYGfSfkd8kirbL+sQgoS+Rk1krHGCHSP86
SH4uGXCLryHnlvxSt674mJCM39VhTPz+CPPC1TKXMLHXrf3BkYG1xR4BKEQMB1c2
tDjVkZblw8AvOoXRLh+nZ1DtQiU/rmXsfVRqxFAdaqvPdrLQDYykK4i+3Dfx4e9W
B64qtTeCbjYJQGf3IQcaRz4ls7aDvnjFrXpJVbQZGo+1gj3uJ8bzX4Vm5WvqSM3R
76YruZEPxLNJfqagqi1A0UvAcn9U6dL0XPz4XLhjC6PpkFTU6CV6hA7WDw1iCTK6
vK++ZTKz/qFyKuLC2sEdkgCAuEqoAAiq3/KALB3Q2DxZSLEgn1e9YBjZrozFJA4K
cWRPYaIohNdUA59HZVJiRibzqin5vEpc2B0lOJqgBgmPyHAn+4vTvaJU/1/WfGEk
s6UFXKvcD/fYcvcDCW6vN2Q+x1hpf++XxCkEsJYxNKbS9KhfRw+xmCMmgqXMN7L5
pPAdAFZpT+WDKDnvRHSkumhKKN+wQGGmiejFI6q9oUaHcjCGNllJVapkyBnSulE3
FJbj3IP1fi6zwBl69zNsj0H/UcK2oz3ZoO29I7+VitJG2JF6hSR4Pl7dAspmY/3b
0P21yozzBikZZqXlZtDfQHwnCU9vd/q3NZOvntBGkvnFIVLjqLFj+a6X7faxjvW/
g7AgpdwvTeM4WE8p7eQgmxSABoUvke6YQ2zpqiio9nPLVV3ACRwRbrA53ydIGVE0
Y9cmZXZlGo88CY9ayAx2wvK5H1GEu6IJw0VQc33dRIGVPSy/OJruR8OK4T7IfQ8+
+3lVZ5tp034+RQtWK55Dow5Q+0KAJ8yUPU3MhEbwsnVq3iRi8uxgt1QzvPGjPgRF
i2gWZYHhLVE4AatYS74WgZoDauCOrO7NLL5dZnAhJV4EzFwEHAKnk5zFXEZe3Vl5
Ms0XF6DV0GpEIZ21BY6iQIuBjr3ZW+dcY1VuGQhT/CKPjUCErAJlE1ThI7jekTZ1
MqzdBV/muh16tOPL0fZRj5l8BLRPDwzKIaBdsGWk8bXO6TS3DwMySnXwUcO1Op7Y
L9ieTR4hSebDQtCFj53DlfSNoPq42usM/sPzekUT4u4zYq2hOi2pzYWP1naeQE8a
ZY8pJgOv/cdug9Op1nI1aNOnHXOYbxoz9irb2HhgZGDgnIW73IZ0YSq3Tti/wRyR
7NoNgEybHpaCyfLGGbL40d2tLCZ9RgMw1oNyVX7GZga2s/4B/NwrjfgvtY/oVtoy
qxDmzOcMv/xWaPTDKo6k+KaVAkx1bxYVy1s8h1fg8jZ+o6UKczQCcKxT0Rm1nU3A
qBJAFzBLlw4I4LEHk/qFmMS2jNIwUOgvEcVG1OzqHLyr9aqxg8UBFTxahJG7IlKW
9obFj2bU7nKyADA/qcDSot6kHmdjROcKF0PlnIVBzd4BVaTw2CDQ4zy54D5xpY0T
kJR/MuseUfnL3P2a7+TDLlZ/cYqP8DkYZ6CJ3gysqCsPDgfeLjjzgKNxcgtIgX3G
aKsPNkBXpfVcy2GrXHkX341CztQVIdQMyf6zM1ZmUJ8mGS/MMEX/hq2DhzWRKcae
8L3sVHWehMAU9iFjz5iKJt6nF3vdsDyzegIciXL5Mlv6Q+V57JPAbZeErQp8lK0G
uBVS9DcZUr2oVdqPI4aUH8Vr02uUGbg/r2jpOtLzu8+F4lDmvmBe+hDWcRMiDAZi
NHY05olo+vw4EhEVAB/3FF7I9a4Xodc9RdKNmr5xK8By6dAay263N0IO8S+VDgmC
BT/qcOpZKEVCWXVVNBhvrdRLqy30KJ/U1IM/tPoND1PXNgNn3JkH6Zjinf9haBzW
K3np5tvK5PFCdqNkqV/mo+vE5Lg7yLGFx5LXJDjF4e0iI2xrHIRcDwOdIzQYhsZy
iM73vkxlyWuS11lVkiAg/BrGF86J4Zh+j+0juH/aOe9CkzbaTlnDicV+BaQKsXja
7jHTggn9VVXQflLLQEWVctbjHUcF84l5Z0E2B0K/qceyhrxVBMLIqmMGhH2A5R+P
gDFFUXhZ6B5ReR8lp5EPSxGXPBdrY4QSgrXENlBOQUIDxBCne8Gr/GKvp90ud/Ed
uq5hJuDh4EidkLXinAkZ789YW5YFjvQ0cXri46zxmejn61XmI7PvjPYliXKkptyi
YZwmj4QmFiJIkBIF6RcJxW4LQ88dCveDuIxYbEWGudqMpYPUTvx/gbJGuH2+PTAV
LtMNM/5sGRrzDRxiY6OqkurMyaHHp5mLRR0SXG+BKvlYKBa3lFq12GWX97vGfwUJ
doRWJZVs9EWhG2HtYhEsPCBSoKpRBy48pd4fP3UclQD+uJQqeSE3pXl5QqnSrIE4
X5P3N4CcOu2Pm/hjcCaLiTW4AdHM1ZrqqjNHbGrVbd17r7d0D47JGBNnvARf2ioX
93Rhou3VNNecIbjeHGCxDrH3lHa4+avcqb7wYfCO0KVfz9b0OyZwWc7m1OQsc7f7
mpFKf9RCuXdAj4wdgFRSSUZFYQRKX4rVc2sCfDW+nuP+syeCKcp3Pcgj93LglJDE
qGgtovd9cT4eMv7DKxQ3Qwu7Th/GFmBgrVMq0Cuh1T75jJcktYqnv6qSr1Ce95Zn
I/lGKWPSbbY6OjNjd0y38SpBX44RCkEUFCZM2kp/SHhRTNys+4u8NMIGzT9FuPu/
hFbK1XDRei+ehpXesZTR/8CkbVwAXuiwN82A9RsNHB5iTPR+Usii0ezOz+A4SOC6
+iWEJ+NW1OsJVpDI1snRxgCFyvX6veI9GdLFtIoJ4dDCySaYyaklyshtsp7hhSs1
i8diCjqia3EudpckH1Afa+bQwoiQJufgetjJ3N01/XbMG3faEX0VeDRFjh8fsB8g
Sauz+nPZjJotldsOx4fATv2Hq5jMLGPHOFH1GqCag/6NqRj4IwB93TQYOboBt9Py
UzkRLHYl1WsxBchLYjIiXBzIB79Sp5GgfptJMZc8WIPV5nyyJAl4KLCUQaXqfBoD
2Z4/WeU2SvLkCU2MB2tMciYYVJAbbF9vrmvdoI5xhngo65qGoSO7bZujedFBsJRY
8Yn6w3lxSyhn7F6hq242N+rn/iRy/jtVoo6MP3X/ILH3M/Kn2/OPWRKRKsOfwTnn
`protect END_PROTECTED
