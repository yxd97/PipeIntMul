`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CGcXFDOwJa/koH40295kIRtOkDJFlLyJ01zr5FQcGGEkGJrhxWGlyMPqFh9ZkFDR
oDPnqqpbtmuzSCUKR2aHQaRVhJErfX1CDUoY42Qh+pmfVmJNMSebJ7PtDy2otL99
AbMdNKRVTX0atYF1sYsov6FrKeDdCRcs3Jxq3fZLkby7WlLevI93o/CSt/C2OEUP
aNgsSLd4t9f3b3SAB89HLA3CioLMZ3iTX65KJtUuUcOpiCLcBxxLkQAPRIoqbc3b
VQAWReL+28inYiThss3rcDVnnLvGPjv37PMqK9HvzQnChFfhcyASzu4CmT/7oUZc
CL1YVGVrl09s4Y4P7Q2QRbEUJBJzOmEFL0x/GajidF3I34GCQIlf0Uzwdh3UeI8c
AMKLMaLtmnfVrn54nfJepCN9zVlbwfTbKMQlq22sZ6b1A2eZ1gnHsXplccKk71xt
teTBd7jYmmfnopYT62rS30PAwSyVOMioVQj2tBBjDjYMk87I0sH0Y6go5ndu1iFQ
74xomDyb6NkkfTtyKnbppSs0Pv57s/CfnUz/FIsV6HDa9muZqMFFHNtL3srL/62v
nT99PGY28YaznP4y4hg7BIBGIuKx+SnMdES1of6eCMA1Vyd0CvK/yaM9JmNVmQZW
tXxOjQsaenj3AP+QVuzFvbL1fJI+SMCf0iMCGqimWjE2l2J2Wqdl26xvUa6u289E
P7Ee5uyaWUaaklnPMf26CV/0vDqlUFZv22jHcwC6kdIh8Lt9hvtWQXf5OqI9sK4g
LCUQ+pW/CzHyoz2jIZUzwaPEpQa75Sq7wR1IBd5sfY9GugdAGYa3u5ODGq7Es6ti
CuVbV4mf717pA5dTJmu7PKACPdUfYydl7yQwkkDWGNmkEydznf07QnnvqNrEUprk
`protect END_PROTECTED
