`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9WV2niUcXaXElyExOg7KxFX64AFYsEktRnMsjE9zCxhoEMjcqeZ+coJv4PR/2LLi
gR/tcWG7BodY52VsL1isaq9b9TN//jwU4SnWKwIocBOc/HVxlrtdaXYO4wY2tw2H
KcMs1pvMsRG1YIr87F0352lIvT8oZlFucgRUpZysi+5QQEtMoIo9O4+cPGvQy8JL
w5bVretiW7q+cI2LgoZxj7WjiC5m1z6/e0yLBI17p76Pj7GO595ymGnXZdVNbqHY
z7bG+fbVgfUrZzfhkw+OCovqwslkUS2X58j+cgqvB+9qEtnjSpEbyOLuZc7a9h7y
`protect END_PROTECTED
