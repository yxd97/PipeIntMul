`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rmbayleg0xbE5UG5icsFyq5xFxuhDo8Ae/q29Gqq9TOtDruX7tqqxBq95I+2+4dD
fhm+cRZH3D1Bj9r4w3naroVwmKsbULdRZgHHE8BGyjeRWQPbqdAdShuTPdNUZxtA
lmINuY18No0OKotEW4bB+wfwq/A3YDZzhn0sIvZNY7NfWS49LOQMpez+dcdJ2sFy
/XJnGe3MmsHywGRFo8B83hoL15kpHb34QnH/XDPbesjUKqyrEtGBhzAwSnNnONMb
5LnSmUvPt8iv12Xq6pl4l0s+eeyTEeRfVKkdb+/O007LbIOgN69fUAttQSPzP460
RjnJS3ajHla3TpDMrcxcSTAltsGZq3nZ5n/NhYT9lXUXj8M01HxtUTziYRY+aVT3
xXnuglIookouS+SHHcGn7MK8lKmncnvXg/mBhiAGvsrwwRNRyOXY3K7LP2cLDOWF
RKZKGExQBcANULHlnInG28gyjMyBN0nCt8S+fV0UutGgP46w8PrT/ZRpb3NVCsEw
qCLtbpBBr5EMHDgjMb5PiNG5jUqb38dQT8ZAiuPpChUipe0y7yN0AbQe0Gc2dBsB
`protect END_PROTECTED
