`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YvgaLqZNdqq2tk7buDKDx5f2EGsHMIv8MGYuM5UaxI1yxNeGoz/MFOc3dUscy9rA
JUuciaRbg+q45GcduEq4H4tFywXTwLSwYxxTQZlb6VNMTvHKtda8A4c1sCT9qgRo
4imuxIVb5p+FUM/Wyiu3tnqJKJvfgJcHc+DGHqX0bpZmJin2PTTg/NGm4cqVKSs1
dg+rtsJjmIUp2vaQXG9IBOs5ZchT4BET8A5fR8i/V4E5kWXUqfZcgExG4XLYf18d
8rEEZx6a4PGi1+QQpi84ri/8bZghc3oChFJrzg+An3w=
`protect END_PROTECTED
