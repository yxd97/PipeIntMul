`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RnB1vDtoF3sTvyBeCKKsfYs5vIEXmkNFUJaKhYkXUFSwCHw2Ropf8mpb/LnQDlAk
v3AxbovRw6Mt32NMGcbgj08PDQT7CiTbmuHa8z/kl+U76nejdCnoVuB12+1d0q/F
ggXfjtwsCaszYzfzpCiSx9w5DqeNiZs8dRYDNAk4Kw1H/UKEzA1tM4MhXomcGHdF
Rx0OJ86o84tUMF4wgoHfUx1yr9oMESB8RguEPu7suqVL+sffilLSR4/RGyPFYiUw
DAM79T5mg6IJO0ISlOR8AGbWEaeMeZfWyYbTp27UwFd9ePDyjfux2xPHzOHPZkqA
BK2L1Cnu2NCGLpd0+9VodOMvXCsV0yO50siL3wcvvwSWrW3/Q+TlhqGhO7MhGq6k
ZXj4dhFdk0hyKlSlaxzO9mWRfEeG2zKmdUasolehogybMyXJQW7lepunfxCYL4aD
fcFCFFk7ZrAuv5aN8vW6xX0Qzrp4rUCSM/fdEPC6xAXSTxQYNJs1AbETU3tG6g4U
DlO7dT3qfxUPn1I/OLhIx6wQV/pvvWnHbv2YThd1/Myr+sLd7281Mo0aKGFE2Fcc
lWcA+tf4HwmbiStTSA1k4o+U5ijLzllWNKNINGw0lKwHrYaWVh3pVanoRcdZOntJ
WNVT68AvFT2bNGzjX/UCukaIjjy1yJbrGDPxDJUrUlG7D8JM0mC8kriILNlGB9mb
74wz0dV5PBP8Pp+1o4SwScOpoFsztBfTYwsUyfz7icYXgCC3aGzo2GDYeK3q//Td
G/COevjFPxB+2FKP+t+Xw1sRuN4X1HgJNZOMAGK7uHQoimIS2DDsl1DifTKeuC9Y
rk9sEFXdarJ12aBtlFyjxU8FWdeuXbYY4VHycSZw1yjoR0tnB2zl4WRo6mMNaWvJ
+QqEFJQBVyJHK2zwkmxR/2Cmez/PVuFSM9cD/VpAkcQMmiWDEOB4PpXDgltRvfKX
ACLpVxSNagKG+N+RQqaNyl4wBOVf90Gysoh1ajKzf3RRZPlaY7CN2KIdkSO1VoZZ
duzG9Df/RmxOClm6KwJftT+YSwu2uauePc7FPNPUswGEiCZni8tamDS3+XMl2P1e
lToaIV74OIxBQqN/lt/wE5Jdk1xHzVy6pH2EWkCxCbT6RwKkE3jRXVwqw7wINGbX
abgbiYFC5Y8BDZYWfoUuIlONzqR0SqDG5URjQTzqk6UsHqaUbcMyEkvmd2emy9ZL
zMbdKy1brV0wnuQzuAFKxz0kxP59dx2Qc7+DCa3ZH5iKWRlLG65f0UHpQPrDoyIq
5J8frhmS6tz99jHqDirV6nTCAc1bysl7KRLuKT+kSZkDxMcYPkdWdcBaWg9bTE5h
zFHasFbnnK1JyMhgsoPaF2JFYqa4vJSe6G1/YGxoMXAP2KMvqnvFv4nkc/Dr7eSJ
xuZacCm/7vw2R06c8Lpr2cy4W2XE3jYry+hLSKrnumNYWdR3EvnWWdmB5EVHOvpy
Ef1JwkcDqnDsxN5TLsGi+LxJ7hx/4UYdrMK12L4Mgw4zE/eMJrPHrp4MOO+aE3so
rnmERIk+fGFzabGi6erwesi6vbkxeC3OeyoK0lRNvsxInXRoerL5C3e0KmHIToer
u/gWbgMGVJEFwdf/Ru5BkraMlvveeSlcGkXOR0YwO2xq829+kySadbzPfPqBOvBn
orLb1iY+gzbRe0syiKuKKax0MV5w/hAtfskb759EVlMq3sHYVSlSwK64YTsqYDIu
wMRRCSEmm6fha3/kmxDB4KTKNwMO+qII6vb14jwCzex1u5EY7cDt1EPUv/rMt39x
mRBdrjUAcqVC0PsvN+rJrR7kjecsc23y6azKQSpCTPu35vVQfpxHZ4k6WbseovX/
WbqTZD2U46kH6RPlmj2mkSPCFmzq164frV1NTIkjqgO4DBiTIplWExNplwCnwF5q
AitF/sarLBvGMZVWfHG88TuZXVgf1Y/5bM5VikSb46fgALR7S9uJXasBqnXYwuqV
9TqwGtG0GS7uF4uthkwPJVZlWUiAS38MkP73F8OIQQ1zGQ3REOUypbcl3AcLF2Re
fAT9dg6lpRVjN1PPISkOgekRRniW7ORtitJxBUIGDNvaKOoodysdeu/4zIR9PSlr
vhgIp3VjsZ+cwQt+7TpuGknYvzk8mdcKHCABjm+d7pVB8Mwm2QaVVH8OfOVyH7VR
QIi/ODhuJ+XWG3OlMGTyh0lSLhljRgPlZMNEG6Y1t2t0MAWs7TxkcJEQsSgGaj0q
KJBSiYLrhhZBGDMhWYcarjJ1HndWLnOmccTh2UL68p5qQmkcd5snG0Lbo/FcHBYU
la/75fJfvItHufnLSOsKfhw447VAyUtaEG01ZklQtGeghpBAeOUOhJzYNwP9P4PJ
TwddRF3dEE6DawqMfn4pIyExuU0Hlg4/DGzH1KKYqPAxDl4Uflsnm/XVA+t79JdN
am5qJGMw0t32ZOj+wATTkZ1ltmV0LFOHRj+kN7JBvnUTSkKUAPMwn4g7MODG9nfV
7QWypdnlb6Xeu4XHp00Y6hjEIZ7qdjL2meKb7epmWeZvmzyB2c9i8ub18QHn90EE
X8fg/qGcAF9db1WP4wPAqpoOLU5Ftd0uPuohg8slyNwHjGhznJWli2y9eOCpDCy+
t6rWV480t82A0dScZNPa8Z6aw3oS7QjlkQdUWyjMB1wis5Ew7dl6G6KIYhdCpJlB
i3xVxyGmEx/ii0U6guDwrSKJlHqRmV3cTQKGEcZpVWeLz+CT37OCwvO5IEPPjmCX
Hh49++ovAftTbRDrrkVEf1JWL6mD1otEUeBd7djioVx7WF5Rm5HWiob/EK24KeFw
nrm95ohJrVsqy0SRDUIhvOe9//V8CJZyGd521ZKZtOI67HQ2dCSEyMHHy0AdKZ6s
KvqdzZMYc1jRXIi4FxBVKip3YQSto281KT5Y9OeE4WLh4A2bCCqkwptCe8o8qhrb
bUVhasK4Q3xemshe1krFCeB0l8RUpx9hXYtDxjvbOGy10rvdMs5qOXrlcL1xMksL
o7Xxoei73/Sgal5G64cUlbCUz26YjUGQZ5wefbieV0jJqs0KtSLOMEdHcPVoYc2u
O28h2NRxVnyO4AwnRu/K3bZMJzP2X/rQFSMAhfQj45jXJd34PDJvA66eTJt7MY6G
InzrYQfBZR15Ia+57t8wdjxc5nGpOWPZMGbdY3V2+76upomdf5bTAdF7aLdpZ4Lo
PGn0oAJSQ82FogRvl08X1p0KMfRsbdVrKBe8Aq4y6p280/iEdw8k3BZtDum3r/i5
7sBupaOn5P1a3tvni9BwQbgDaxarYStoEWFEUk00ZpSh1H65hgGZFcUlHgJ6TRXH
60qeW1oY8IuEcl0ogXz+TOdF1Fcu6Ps7oH4S0SeMs8vVT6yztoKAGs/oT/LdGsZV
+1wXQP8NSSsdX7NLp/IP5poJO32dSrf5GorotvsgkANSaBow7O4U6i6qSSIE1Yxs
MA39NPFtkbpvjoiIS2rC1tCYrEwup8K2bvMLBChVor0=
`protect END_PROTECTED
