`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4kL6eUWVPEnhh6r4VoOFgiaj/zOpfgxegTjJ8ab4iEVCp4aW3WoybtgB2ySnlekj
aiqRqqG0H+DNQphngDbhWJITmL81/7vqqpPX6PXARB5GARSgo5a8BTzlGLyjFPzS
nib9rVZ65XyJv/hq61ubWJrjrQdhCu3auDut1QzwhbkWG/GQZ2Uu/XtgpEIsyJVh
XlmvmjTA+JkGAdyuMfBEPxo+NbxtIZfsod4BzdxwbxhkSzpvPOEbfKxvCouidHCA
LkkhXWbHqsFMaMQO8HLXcnCGBj2RPIoXW8j9yys4mFOKeizrQ/jYhviXpxuPKyGn
jWQtTVrKkMFD4Zmh0lpS+A==
`protect END_PROTECTED
