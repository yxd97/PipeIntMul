`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GG/ja/IHU5ne89fsi6TQZAyxzRqLJjWQMVzTY1gGiGXJnsE35QZcrBqbBoXohFVx
uFqOa2OY2vAhlwfN8ZR9bZjlbFyuogy8BblPWskBXdS7HD4hBVj7zsYTxXx21Uc9
EBpRLpSZoSTsW/FykqdtUCExwMY+Dg8V303JG8uoiPmMyhQMB7wrqMSooh8Q/YRh
eVZudUryrC1zcZtg5gFlJ9X3I4/YT3VrEX/ResNmFkfM+5ZqzciQafQKLVT3Yu5V
EZjO7UGiBGHUdcZvdOalF1B1cUod9GbQpYxs0maxwaki4g1JnMcaW7d4/G8xkT4y
B0cBeNqz4KRXC2suYbfEzw==
`protect END_PROTECTED
