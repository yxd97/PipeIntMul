`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDpNgDGeEWxwaVeTKCPqvnrjscZdyc0hGrzpdSu4ne0L0CtHL2UQ/HXyOMzQWt2k
exEQSXJAjIpBHW8e83dXMcsUiVIbDlmHxl4+VG2PqNhv/BHBOgutNv3tnlNZpPCb
dU9MzSlt4/cBBDlo2b1uiyIk9/ttJMzwFEzO6nCjywd0Wtqctb2Gc+Yk4EDvqSzW
qeaDY05x5lqGNGE+/Rfv1im3JlQviVuXnI7M/iGWHYX/yFANq1bJ1SPQMKET1+xE
HjRyQ2C8Umztb1Ck9cVvBmynd8wEYCmR4D4iRIHGaPbEcoIr0JK3zbEqqkiDLjuQ
/DeJWGw3rXG6d362xrUCi0w2OQeEow1S6RslMYuOeBbA/CufvQxhj+XvcWnPx7zj
s7t5WKqCOFgZnlzFp4mq1U48qLhHs3uOFxwHMV6eFSz1xgI7JY9JVx4GyBH9HXs8
nygeJ0BiI5vCV4MdlkjoL5aTEVq3J2tLwBBGDau0C9EmmdNjIeeICxG1UiJaZWue
wXrd2pF059WYQ6A3UQfzuF80YGO+VtiaCEDFE/wmrClMiuBRDu28G0ObDzdMxGjt
StAyr5xqcKMHBPL0t83tccAv2lR0kKqX3TOTsaO+PlOmYSO1ocD+qKzzznEvZfUz
AnzBFwtxraiB68AbHD1DiiFUCGM/OnfvIxqgBohnJnQL8Mj4NwI9jkPC40Rpq6Bx
CAdDHiMr0Tp7a9jhnCyPHk90CrkNUsl9gxdHOUf1nvwJH7ZLy8xRyNtT1MP/rT4T
a6Qr8XecQEp6Ls7PCSd/G7wmL+12X0m+z8RqTIXY/SnMTYU+Xw04i+rbr3LfwozE
m+Za9WvP+znuH27kcBZSrEh25bz6q4yuZ4tWtzUueS0rBuHVmQEKAixtkCTUj8WB
T6S+AQwXT1EhHxcfmNUGsYWQt3Cy1RkfsCTkj5CMd3fKRQIAKEbdc03Grj0hEJy9
odYabR0PEQbVRPINPMHhzWUo2WcUl8dD2McoJGLcP1V+4kMQiFCh4wxYesofKk9Z
IQAkLyDH+UqNOtq/DQL8u8OoqL1A+wpFU6sJ4uS6hY3ms0uVdHuXISmfXEjtflxd
aOdg5JrSP2Er1698TgfNcO91swLy4l3d84tUjOYE38uBOdcMtv1x07p7K12Ekd+g
VRA2KRRROE6Qt1p850cX1kqdBFetcaPNU/5sGbhaDk8=
`protect END_PROTECTED
