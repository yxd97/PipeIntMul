`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u695XByL9iAjrOaMOczZ0b2EnU96TXNWBQp7uB2w2v0cD7AcFhuPp2NKyQ+Dkxw7
Lmph82pIDcft8O7xaCwPEQssbS/QWiyA4dS3QbxEPOXRyqARyWwq9drjTiQg/KW6
UXXdjru8Bf+WVIC/kK6HzxefM0M0+Q/YQ02rHtm7gGXYX2a0jFSvP9Wj2Qidsk8l
Tt01dE2dtXO24kkGADNZBI3Za77M3HiZbe3CJb1DU1e8j+rgiCa4nQDaMztgcKJ4
iwle8FAj/O36LRmbV1HvYHtY+JvpRxxVt5HEF2zykb5uG8cv+M/ObXQj5h/Cew86
l/yQUltmDnjd6XIsXYdh3XCbWUHDgqhfox3RFm6jWnFehU/INjDdY/gc4uDm5rmQ
VI1tfpf3yPI+auHQVIhheztm/ISf2ZEescl4bJTIeIRY62uSJTsY4LWpYK97f8Nh
+i+vDwt1N21pJ36n5/KsMeXNwgXN7RdyVU+l95do+NjANpejLqPcwP1lK4oEp9V0
p+H3VylZubqQOVKEDzoRHEjFjQ+BSsnNnToYZgJznDQvBn9s65w3+HGyDCwZ4u6c
7IjL9WMTEAfvzdixZ/mAWbaARmH1rJ8f7UAJ4bNmjtAPAT4N/erNhqwM5dAK4buX
d5PD3pfyHY5r6mZuXvkQMNH6B/J1P63qSdSy+liJARN9GtsM6eZEnmGnKfUhRMQT
0gopuubZ9esbWDEWVQuGIwA7fj3ll+3AJK3Z2bIgQkDgRklEyW+L7Spie0/SeaVJ
2INdM1PV1YwrutzQDsOzUhBzxOdEBiJTnXRGBMg5qZM9L69Es1yUoEI92DmCSf6U
N4P4Pt8Vz7ySEJIFrZodRJlqfjOeuIAhFvSNkr4PHpxJdTUjya+4nbWMWXs8BrHj
R0NVTZi66nfZqnHVB0gxlRdjGol9rzNECI++G2GAKqSVSFWxwRKlRxhbi6iuq7Ih
L5MgQidzd+arb8y2z8qVW+grHTvRmwT+8a5bcMflDAX1rxS0iV9urBtkMiFPV6HQ
4ySNWjn4D3fLv7at5TZ+EH4vRUPZVGQzdaE0ZfmF9w2/rpK7W+hYS7ANdEEiQflG
N9xttQAbfgsM6Vo3ceagbzd47oqh/Csq0HbK7v2wfbfI7Jmq+z2zqbdo9kwgIqkv
4QDpTLjzv88jLe63QzcCwbkqfl4IB4sh0FPCcQu66TLs7E4FUcEQRZBd4qsnMKh/
4uDnLF1Jmp0+vwQpItPvN0Xxzk1mQrT2sIjPJRpxYAq/Sdql8Ad68F0rZ8FCgnrB
mQpaEVASjHwCdvjWujh0+Zp1bOVvOLv+2+duwr7/Nk5M/qBg8bDOtk2B0b59Fdth
N1R8k1X31JQjTcsDmpp0saUvbL2mDYvSTxL4lNwS9StFKid/S2OyIiXHBK9qoIqs
KYz02CtSSF+yod9K2yYlum+nTtBid3L2ozWISfU1021g786D16B9fdBbqBolUkDW
JHeWD4FgxVr/NquH38CsngEqN3wUO+JNjiZrDY8QmpIVlXlLS5iiks9pSeZolmdv
6Y36vRkh2y5vm943sTWKbey5T/5SXCD8HWl8beDCDM8726iknxq+ux68DeM/lb8i
LDJyaBxZZzWE8L1dCT1hT3IJMtuXHfvEgepNNf+5NuKwb6MVo81gDHFvI5U64fRq
aROO+IF/hpuUOFdg3uYuC8MElPF3SQTUSdpsAgVdI9z6CYoljMMtzU6WHapae07M
TXVSdOxDM9pQ3HsEgvvfR4sFQWuodQ9oBsQIat1p51FKxn3BcO+cjDBV0BguhESj
fFdRJUJcyNyyRUc3IAi99d6n1R6VKVFqiH+IXLTTtcXnLgZQNh1Uf4m25eZWrnHj
owCi99ye3efaw97hH2yvhf1jPZ8Phe9Hy/L2tOMIC89MUDtdwXUXdkm7u45eIUpy
EixQgJO/yjsHG4SAlwNVenarHkaiXHL3bo/WuSwKrgjS5svICiCYPjwUZA9tqGgJ
jq2y7CcRm0ivSUVEbylBJk9H+ln22tFcOUV+Bo5SHozCZx31tFWxyp5Z8g4SE2po
jwpYAXnHngeUgAdajxsmH/C03jBAoJn9pEpo53M0yv72E7unJN1tKX2s4xgOpw/2
Kr5O7d0vQ3v0y/m9D3TRxX4fARkOoJc+80Rl2euJECrldp0jfOXL59KQbThwu0wu
DIZBy6C6KYF4To/k+Pf9zcMFVQzr81kzLmhtWRU2EnKf5D4P9LRRxEao3fTwxXeH
UPNQV4BwZzjwroYRc1+iwhPPUAH8ycV1yHCDJeEIpQoXsUMCjhpjpoZvlp9HEkH6
Od+wSTbR2pxxRIniFXx7i2jw2zGAgdWjoYII+XjzkNLWKdd8vrlCMuGpcedgpmdi
vmbAKFPLy2AUheOHpuYne/zHmoGf6J/AjP+sOYbB9WvV7WhZPW9E24SQ3Ix1/4cW
cgbXOCRRCeGhDWGBMTYwVP/tRLTLT9cz0X7AFE0s88ltCX9tA75pYIiRRKBPjy1A
CekuNKBW6ZmvZW9qPoOSw8V0K9n9x2mVTzXisFBFgRrlySHG4uCDpqobhyTr35Cn
hDZu+TC7B7czukEGaytRzOmWcu4VbVttkIbPhTGxBfIiDglqnbD7YpTeFDQ3RmPb
8OiswmwddnaZ0at3HkmKPk8oM5xcJdE35hiJWT2MMlr1FzitgpnqgKbQnZvr/bWM
3Y7082WA6F5PkAXBaYcrWbVscBLhRffRAWrljBV9eLNcQVZnNRvP6P6PTcUr9wV4
6gF/TYrBfwGYJT/tuV6dEAKBzp0GFr2IzW+k+8e/VoUKr3p4ohZvkgytgMhZWZ4v
/m90gN35mDB6lKDUxj2PFEtnFdWwf/KLBhKMyjEE8Wup7tsEWsQZbmTIvFQFbRS8
WeDHTD2MagP6fCxIdx7/+mZVWiCZ06OQZvIJ/7zYHvD9y2wJILgDLZiPERhjqji2
SDBwTrZf/vxIBKZcXT3ZVKY+Wkb1Advlwe+QsCX/zYbFJ/FsXB88MHln9NP8eNuu
iLrA+Gpn87zMFy2Inyjx993/GeiFXoKTF1P6qUoQxx4eqiuUZmHGYbhJ0AjPVM00
m7vE9PaEMRd+ZdLQB08dBJIfMogxwc8dKzK8YTbR448MgZNicSOkJBD2z+cdTwOe
o6J6lVo0JRhDkvv/DzcgGE2ZGUYTlYuXvPdFhecZ3VT0h306/NxNDxU2+o9LWCJh
MZ2V7vfjAJ6pZ7ZQ1ZWYSwy92gB5Z+qNqsV+VZhigXGEQvw+r028kYG/b2GM2+We
TYKi6MTNQb6fjDJfC4PL6gVq6ndQg9h1RG2OQmTvnAQh+nf2mkYQknL4TAa1/UAc
eCIhb+qKLMdrP4AIEo/0dsgDziNW6HfgfgyLUj9elZpsCBZj2y/wQG3/jb1NdU3I
`protect END_PROTECTED
