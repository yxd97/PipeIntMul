`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZOSOHUVr+9NG/KXZmKjtJVfQONazIhVgtrJuwQaRI8PQ8ew3yGdB2MGt9WWXSbgw
Q+sLojAyRBCINNlw/Fctr3VEJPqJVShqY03Tbijam6pqTJWjhgH5V6/9W8iqfMK0
ZP3Y1DZyGHDw5IdtA9YY+maI8y6FayyBHrfX1HEKz/h142T+jgw83eNBr0fZzmq8
ALY96LMFm76w32PTxCLYBkp361RtNcoFVdz3zyHGBolMtIKqbaNFkGGVpCM3Ub+v
XklPEGYwigQeCjaovWkRgnJ1oKJiKHvjOxRzUYJYI1Ea8KqM5oqdfzZWPG5AAlSP
Z0va62IHo4lyz1kB8OH+lsYG4xh2gyjMJlQJIQgUH/wR9yu9CGkaq/PKvVYNl6q6
taz5HVqVbl+dCXoB+/wEjwSqZtEi8AwaoBUu4Zs9NZb9hKo/amMg7J42voy3xCrs
FdHMo1v4FzYRpvvIqMbpTtaXXJ6RwMeC4bmZh5w6VAiH1Ecjj+CAbZ/pbsUAMJwC
vl5V9M9lu6u02OCmMmVRmN7n63bhrKLY2pFGu4YlH6Inj1zReIdTIweY7ZTRYdi/
cjXZnY7o0SS975SjgAd1+aRiFr91ypz7Wo7bP6B1/WtKTbs/4VB70nkhG4yiomkY
6SCCBU8U/Poo5hI4r/vRRqnXmc9P9mELX4bnNQTdgUTwuiYrJTA23KoC9jjDS4N4
0lQlLX7SBaFWiwqUkGhp4rjCbW9oVBgNLoeS0DKx4QAKO3/1/UomXa5g3VsTobUU
JoDC61b/vHRN0Z8jkqFAXvzPipL3/nM2Ohl0gDjKWL4VtXlYOPEIz5rxPICA3Ot1
3fLkLjX95xjMOy5cSqQ4t8N+HSX0jBbG7gwgPLHQwXYcvlGPtQpYuTU+K1ICjBvP
QrVL35wsMeUFm1shnSm7RuhUtcICU/PlaS6B8tO4wCT1e1It0XCw2C7Znx1uyH6P
3eN8CZ3JIb2bZkAUqbAWvw==
`protect END_PROTECTED
