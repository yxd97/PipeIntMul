`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6NI2DHZgcgJAyfajdXfOmc9z2SRhkofUmPbYDKfyrtB9/RtP5fT4asX41JgyURb2
Tda+pCBnkimifd9FQNCaPD9pMDLJ7leZcS5+EeOea8pXd0pjwoy53VORmWr/w9S5
BUeoVqKTzgcC98TiPsYLXIZrqmowfWG1zz1IdWkUgkIyGLOQfUz3DATA6+jBCm/z
7gc2Wqa7lbjyA8mzdNgG8nBU6L0mWbUESOcd/NL5XMWKykR2m4bk4IKSZLt7DUGY
3SZJG8y5Tm0/0d0C+mExn0r95sY4HOvlc3YZnd5FKVCvViX5p3kXMOWaGb5o1lNk
ESAg+/gUf7IY4JdaqpHLTZhcs/8fidcLEcOINGlZdqMrDeNwRa93K4yfM/qjhXz+
VQjEPo+sA2neVmmxPA16FkXGOFjZUKfDyZ24m+sXZkLXk2hQ/a3boVLEmCr16lT6
VaginDTQ0smJwYBzN0Tp2C9EMLs7cklkse5HNxcR4hkRdbdEqUtqLKgJti+/NaKL
SHKHzax/tk7QNH8Oib1lPXi6YfFFCmQUffbgThPujRrZufj4h+p4d8X/O1Q9NUk5
i7hoC9Sgi+QOVRfg0jfYz/yS+4fM+kdeeYTdqNwhWepC27IAte59wXlAMSJ+s1ho
eLQ57Xe1Zq9wEEwSdhoIPo3tVeM4WJWOvjNoTvUjK1hEUGgnMhINgjwaZuPJz0GI
UjOjJXe6IMy+c+hbhxk4/QcRPUg7LdIPlvPvZ44e3yM=
`protect END_PROTECTED
