`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aebwzwsywZ3g0I1JYkrnFfnUKOfiXmJKwv3uuE6WRwPIHIJgSlTFM3wL4rou5aQv
gSFOyuIC0K9HctS25WjHBiu4+a90Uids9POjM92Ior6sGhuVuPXJwpF0cRxC7vOv
di0gleSux5XBBWAHpHUT2jDuD1NiYOtomwMSua9+NOhFjFiVQLHCdrKpTomzFAXK
SWGF5WFIsNvNe7YaUpQWs5NUKRax8V9+2ocbx0Vi9I8wox2baf4FZ6l+/bga+vVX
LpTPowXNq7VRWuJO0AKQBytTQy0GUY2NnmPMl1sttwtxCKWUMCRJQ13zBCW5efmH
bQu9gIprNv9p6zgb5yQ5hXAU9v2ADsUjDSp5H9P37h8dBvwF39o8tZqhRWe+qvNI
`protect END_PROTECTED
