`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+Le24PcB1n+TLI10A3byvVaP/f6btTJAR+NwS25h5ISGErbj3RicdV8EsDqDueQ
crCk97Ee4mJLwN2RG4IRBDxdWtN4yGZJGRgZNQ4MHnJEa55ibNhMeJ6oqSgUGK0L
3sy0IEU4PTeyxscjWhj9SfntAoV7Oh2LsSlzri2ylvAZqrhdxsKJmC6graqJ/3Dr
hwlJAYm7MnChfo7apynADJPXt9Fx04kjxrrCihIlEPnFrlIy7iS43Vn85b620F1u
ugrzDHVLfLaW0sLWbHmsI2BL7MJ7KJ0tJF5HhS+UaOIexp8QMtljje5axHC9O1Zf
lbLRhUEDa1pD/RceiawCo3KaNwsoHdbOpByEQEBEBnViE0lj9A5QmujlpQ8/1Mpp
onJjN0sYkJCCX+yEHrLKINHXpUlRAOHNJNX+o5p1A1rlTJozF2QfntiAuvSIs8mn
affk91UeF+VPVTlAff3riCbqg5smHA7wcI8UZ7VspYXusvfGUYwqLeWXSny2vT1e
u8VPQqYo025H0B8whK/xRFZ0ifNpTwuRl01l8xX+PPANWpb7/qmnF1AaaaBRvvAv
/VT8ZlNRVVvaEEXXLy2GesrWi5NgdzQL8TdUCwVQoQqZWifO6W79OBP+NO27cYaW
IZ4/xni6uwcvKxXNKoJ9Ze/nHDYg/rl5VU/XH7uiyV826GaU4aIFoW+U7tOk79F2
HpgTwGcdlqn2Q3s6EM4/sg6wa4Duv8x95ds5bJDnClb0hu/Gs/cEpM2UB++QILpy
6N7JdV7K64C17cGUfy3ORB+DMU+pj8YZf9phU4ervw04+aEnn4W7cl4hJO5Z0lPh
nGmnKFO5v69l0lB9+kvFWpoBYyETLYsM4txWni2tU2e2LEVaiYllAW5o2W2cHMlj
fMxnSueTFFArBjCsedrqnP8MktokDCjDG2uRpMEU0jhj+5YHqBodm7StgU7QM0k/
YrN+kJUpSp9XoWHLum24jNfybsAQtXrp080WhHPufHDk9CFc2SfHEkqWCmT+mHz4
0Xkw6z8bj94bEUDRkuBr4GIXBUsFnW7IWDIVWtU8hZNEkN6sPgl3mANKOK2+/Ocj
NNMatg9Kec1KW6e0nGuCD2EdUfN7zEXyRaK/7+cVr5mn2Ysvq6vuUlGzviwCv7+p
kcaUX2V3Zkef1kiFP/pHvvT+skBoxLhEScvBRTcQem7NHmjvahGGKXJUFMw2/xzs
`protect END_PROTECTED
