`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SShJ/id2tumdVg2rm8ZsmLfpcqCRxZyl5nRStenYAC3RKi347E+fI2Dn5fz76EUu
X0mL9kvD1BFbNcwQ4zMXOICkaklfo58BVBgII8k9z1224Xi+eYfloES7YFeT5U5D
m5XP5HIe6a0P60tb8Zc+BUIjmh4qb1FOAjtdZDmBmUfrGNScihNaPfh5bzhsB6R0
StcvlzuWmRUCRxULjLrui9XUhVUCH0j/Buv6WItxRvQGu7P9dllniLWYJv17yHc0
TQ11lrUuI9+7FGf4Kd1DyzVYlx7Ym1JJ5oGwgtANZ+8=
`protect END_PROTECTED
