`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0n1zIRd62ZOKQwpnLT5puHLLZc1D8Ch7POorlG3B6A8iJDx/WS6LhbZFCZ0VoMiM
TvgfZ8MilDNMiONBCiT4ER9CZxtGZe66AUhAXaOkG2WgpT5Jh9QRvBNBhguY8rec
BWy/HbWvyM75m7Xy36Jc02REuJUNBxMgZMQNSr6dApLy3JC6y/JcCw79TWtTjToS
JeV6T5B/GoT2AzFcntISW0ReqFGysCOyiA5OXT0yCqP3FtFee9uLXsXAmM0c4svq
a16CMreKBBsKmQQXgNpMEHg0/K/gxDNBKlGWInZLk6Iv42kJywlcJ/E1W1HAYsrn
bBjy9Pyqx43sCoDTpSc5uAAKM1JmCTDjAm2KLsiFV3rBokhNGGNpYENiWoIh6XP8
zFkYCxjzeShhh7XBJf4TH/vQUmVAhWnnf6HhEIXZYzt1gZAkhlfr+RCoXgTNeVDl
w76zlFygPhnI3tl+GVVvNSAQvc9LZAEOMGKDtJzDERxcMq3l0yS9/ivqSxp5/Etu
LGI2M4YpOi5N1u3ybChTquI2ODiU3MQBdRwIarrSTsJd7Hlj1RQXZnFNRYecGW/l
2zJITnPFpfCxC6zrP29sFILGHP2uBWFM26PD6uSFfIKP1ptfG5wputPW4+GHnZiD
kqe77QQEbdGlg49ksMX4dTEvqTGEemRNUSSHBEFzh6oiyx5fjraNQQXQQFZhZu5r
ouxhCY+NSGhmorjBJj0WocsIAphO+Et2nwmbeOTcQDeV+fX2IjgZSepPWNaafsXX
VTaeka2h7EF4hGHsmBxDta+nElLZCOsawJQV2ysFf2USCurJiDCuBdQ60KafZOhN
PS3nwWm0Y8ypP8Uixm+Fc7/Qm+CyIMINtw7SmHA5Njz1bIZ/FFh80wQunqtHw7OG
+gwuWAmEsZlVQTFWoFnhjH2sFraeRVwxl+VWFFIghds/mOIbgpcJj3uWy8xnz8yt
aV9lGe6yOgr9i+v0yAb0ZQ==
`protect END_PROTECTED
