`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BCSvm0aeXlcU3C1dhEa/CFUD+2OjSipE5Vwj7MyrLVP1ELKOVWQkg0gH4cA8dHfL
hhSPi/OsklsuDLwNpvUgRFsGWhXeMJL/7LBvxTczSE0+swd8W6VXJbbTK/ogLlPO
eg0IiOZgPT0/PUOIR5mqz3U8zF5u9r2vBC4RQ+vPlZT6ZA8/Ez8kilzQjySNy91n
/8Nc8k2HdMkHM3DDZeOF2jDPwO+V87hY9TTw40ILeGi5go5H28HcQ2d+VEddhjkI
e3X4D0H42aqv7lOlUYJlh4Dtzblh5kmDh65u0yGm/k7u1GKT/DkZZMMbgn8v1bdZ
rL+EcnRh+gJrBCiAQDv3H/XNrUyDo/tyD7JPwYa0tqOOFQN/gYmsFOe8KyF9sztJ
tViCHZnbDczW6aAiFms/MqrPfUG9R3bdne81ntKCcfQQ8zOuWaodermzvgjc4ujl
bOYbrAiQnCspojAfydlpsV2i9WkXOfoLr1KZOBC57ok=
`protect END_PROTECTED
