`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsvkfCM+4D7YcDEVDHhXddfmj/CP2RdLrwi3UrJbUKmgKGkWBKUKFESAPGe+7dl5
Fir6burKSB9TeXHjgT0e+jysARpK5Fndqd0VxCbbgxYQj7DoN1cLlCB+fE3hH42s
yHWenzzAMI3F3ve62BR3zjA0ocX5RwCdeesvuVQTQUCsuHIXB55gKFXAuS5piJit
nx+Jde6NSVXfQeOucLI6ijQXD+5aMCWZzHuxvcyDbpXqB76ir0CQvdJ3WfHbbQEd
PoQU/ToyBjpEOMO1uSqxJGpStMJYVthpIRjOt4UY2KS7sRowUJJM4tkWjm7LcwYQ
TuTNvducg0O2a5isCc7qW562OgA3gn7ZHn03KwR3CqH8OS75792EiPqzssRB/BD/
`protect END_PROTECTED
