`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zp5pjf2p7V8/WDwUjg43H07npo06hmGYgMyQH4UxfNn/f5HZIRGTZYZgwthwDj43
s3bCqKEWIlY20HBAiUlrJb9ZSjreGwQBftGIiKc4G+3AUbOT0UbJWuHFA7IF6yEe
4X7zwTqK7zCgnUrBFfHb6eOi/IJrR2ZdrxohluWCJgYYA18w/e5npg8tMOJEGMXf
f+/PbgNS7nWKAtiE/SK9ylT9UFtnVbWFmIR+rJE+HE9FKZxJPjGRBNfgNR54Cn1Q
NvrelBE9f/sW1SvDqY2Jfy9w4FoY1HAO7ippmNLWgJal+VtqeO9fAbUrwofcXtgc
pUcxAZ8X8qEgl2GjLtfBZ7lM6b3a9ORyG+Ewd8qTarbyLkHM/XA2DMyCK+6q/k86
0+G3XkS6P2pf4BJCNQUPmP3EmUHcJhzDhVKECL4ir3DNp0h7g3S8kKxSVuSLCahM
nZwWCGzx4KgURCAwOz5NI8kAa6Z+KSndEDctodtUL1cxdqv6QdGttPOeAB+8JENF
`protect END_PROTECTED
