`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1/KGVVtbGU0jIOInSg7rYhHJ6jow0ryfTyhzJqK/akyraqbrOD8jIpa36XnQE3V3
GMWfKS/g6DtPhC8hsIbWXyyLI0Vy32U547bu+1HLYwcAM4rkU9d8d+aYG1pcWa2C
3aGSXsecbEWPVjbMHMyILS1bp2Jwvcf0bD3IYI9X7qQ6fEbnrEnxeoxxXWUWpDYe
Aj1v57xdtInaW/4cwW2D1E5oy0x34xNUtM+678Y3gXIzDmicT/sD9QchV3oJYtrp
YP5MY6QS34M22ZPYnbig7Ii6vdct4m183ammkDYIcyy+nE63x22hbOG4ngBJIRos
qX+remZBMF53f0RV1fB7yg==
`protect END_PROTECTED
