`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LqgbMRvXx52jUsHTP/aEqO+wHn8TKkuyV9sP4RB60NiLwIyH13BqSgG0l55uSsIk
Z0jJznvnsGC0DLuReJmvb0jx0QdsjM2KOzmYCDdVrFAL3YH/g2XEWbRobt3zz4Sg
WXHEr0jx3k0xwRkueJezj4QRtNjWJDcMBPmel/9QJGhLzZivW9XH/qjcfy8Ufv2k
ZpFInlxio9xEQyn8BkdlP15+vQTddABHpRmYMPoi30RwDm1AkplXbvNVGFsKFhPf
AO+PBXM0L5/3AksUYBfdFz/oVS/vFCRoqmCClB0liQosBbFHEgfPrewE3wGGsGjm
Oh/PzYtRyJX+KdokmfCx58649tQer4iOzTAwkgAtNSu3/aPXB0eRndXKObROLCsB
8WTKJ4ZfjI6xiHK5YWdbQaNPqVn81pOVjLJOEK8Lw/f4mCfuUc+hYLfIpgsTu9f+
AmPQWvvWWiChl70mMSNZAEeu6ZVUE6nPjTBx4jnIiK8=
`protect END_PROTECTED
