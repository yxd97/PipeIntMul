`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3I2pQYdlgAeC47F4N2/TX5v4DWsghajxqUf65eLEp1JHdO4UcRhaVCdSyn2HM2bP
qLM5d9bOIDwVgytGKmqUTaSz/doOlQX/rr62Ov0d+kshnMy/E/8N71fJ93cZzqVT
VEQ4MCE/ytFkYC9zKcCl0WLf8wzeUrlucudG+sb//bt1uyi9yL9SRbksK2Oc3fpH
2B8n5iubkPCs2xXtKFNaQgx+ZE2lj1Yc7QeB2HOg9Zn9Wm6tiOdbdsDvBdUIuuxJ
i1YzpRCuTaAXUUx9K2+DdhOO/QhXbD+PPwMqVJMj8UDGc8b6OT/YPzBxycNUfEaF
1qeThjfL229Y3l2y107SynRhNoAsd7nyNDa82TMj6wYrGL2YNick30rTdREFeaif
QL4E7v7BuXJp+iOCGuWLcqRItsXANew42Ndkv/cxZ3zK5b3d+7xvpTvxna+v0Emf
JMjb97XipkuHneC1hNfKWCTyDdqZwZPLowTfnwVGivA=
`protect END_PROTECTED
