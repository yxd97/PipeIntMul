`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u+aVOjDe0yXFOMuymw2VzR3Bszzl9U9UOvkydhtpQeKxqdP063ZhZJ37HB+Jas9z
zDZpgwwssh3wBr/JVOrPHhjGjytiyx32SgZSm4g9qL9SUiWLW24rt729V61DW0eQ
mUMdWXDb+ipcdMQhHiwDZyrocGmg4O4yFyb2pc50UwuOj9wOc2yTtdgPFtNIE4O7
RgDB3vls8gjNDb2sybvCUqqJxz16XioLUF1huk3UhaDik9f1KwRujbe3aZzYYiR0
SYPE/e1nDwMnPUfTNHc3GB7eJFiUjE24N4rezg9pM/BqDqGuHapvOygeXtC0s9F3
7du8VOH2d8X0ssKnnLryLsA99dt53RWgstwbx16xpjE=
`protect END_PROTECTED
