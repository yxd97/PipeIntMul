library verilog;
use verilog.vl_types.all;
entity KEY_CLEAR is
    port(
        KEYCLEARB       : in     vl_logic
    );
end KEY_CLEAR;
