`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UkyQXzhtsubf4rLqc97YwV3JBtkSo6VVw6d16zDIn1SG9JVxsj7bJ0XApj78KGVG
6X6GImIjqLGQLf25cZsVrDXrli50At28t/DAkmtHzBTVtrj+rrdowr5VpQqHQ/pI
TRVBPr/V8z16FJfnIQCqZCVxE7ngq1VAvR66cE67GPc2ly0LNBAvITABPgzmqQkX
hgEZyxuHKPF1IDqQtvx2qPZkjAWsJ9TDbB/zMsUTJ8gt+bs3gWsuWMO9XuFZagrJ
RqGbWQ8xJUcrq/UOOvgzji2lpG4so1yEGU4UcSLOqh55i8T9AAt3H41/R8HFgk6J
/0EA7gxsmArZpKhBH0ZR6jpaxxcjQFoERZSRDEJeaT/wt1/kk6PzMKZgBhZ/Edzy
c3tZW3WFo5SrbaHCPiJX8/GmxYnPJ0GCGw1jrZyhwJeCZPL5fNKOVcwa1l67q1cy
9SncUk3EvZGWszqm+C7vcP6/2l34TbH2RfD+teL1NSl9NAyMxQI+wi9kdu7WAjNC
qHUBkLzC1+RwhtAIq43uUQhlKxtt+LVmmUz/RdFTsRkNcGFZdtbXcWrOyDwlcs7y
vOCdYLzuZ869u+Uj2RARnHCGCVWPhoqo59NYkur5cbiqqUKup8OLNUN69SOMGUQM
nVIba4jfjZ7BtKgi1sCdh3/+IaJuX7ERGCyxyc/3CggvTfXUWMG0xFgBigYE97So
IgFTjG6wRmm3vQXtOUGKI/FJp3XyO+31DwKUzhp+IsXaPONlMsrj/9yeSt2IZQuo
21X664CFrX5yiWS4ScBzyvJtJASmVpDcBpXIBmiRWRrOlrzPwhw2sZvzG4i6ohyV
UhnWGey6fyZxbM2RgtOIkEGqBVXh8ZmhJhA6ijMS/HVWSv/KedAlHIDnWiYpVZpk
Rwntn6GtY+3iJyOBfL8fcZdjHjzapyu/Itv2ubvpCUXnu6vUJK5YNL3QxRHJeli1
eOWCJ/idebRTcmzFGcLkFDcPeZv8w3ROMlXCun3VaVhm+ZEhNyat0AbVoxAtRpbq
HmHa4ggqteKWnIduwnTH0/+4kGKMmx3eLFJpsNy0GurqHKme7/3ohuYUAPyxOOI8
2JiSYrzWjPBAbauIEOishTrwd/ChlD8IVyaraRqoH3Ut9KwyCgLcYt/zi9+z0+Re
aKPM18HK+pF5xVc/kvKOL5OTLxl/2ITjyaWBaXcM3PXVUfD9Y1xLkgSceJiYTT0X
P+i9YMxalWy04y0hQRDBJhx+pCNnHN6vTYEciFRPl6F4AXrBjMQ8nY6VQafkZeUg
wCLKAqb3TJ0Myy38PYCavZepnFJyyWb6icUhKv5dxa+oo6gNLM/nd6SdQgzOF4T1
kRttp8gSVhfPIjVbXlC9zzPURqbJ9NBFyXu0y1myLcsAe7s6PQprrWJAI9bd/Yko
atsjTEvZ/Ibtoy224A2/rANIkCQy4HpKxvBeBIyvsc7AcHSawsYMh1vCHCZPCB94
zqXtXiEGwce9sZkg3GTELkMoxexnpWrj4blVccwthofLx5E82F/MygqymotXzSPZ
4x78/CLtsm9NtbaB2oSatiV92u0n0npbp3lWvL994f3L3Cz7HcBzVypRN9RLKGWO
kC6FYtFmkI6VrIwJla1Aw9dPSPv8ulKnV+yv7btVvU6JszX31TOpOpJpHn7+BaJo
2/2m/O8lqBnIg0i6HZIZkXguCVlHPqltAJYY+H4VwIEHm4uJj1hfZthENkGobVBy
cHRTtMYrVwjy8XByixo/vgGnQ5Eg7lkPcaH+fUPDwAJ9lbHJldHjZeeCsI9hPEtH
dcm5/hrqYh1nRUPMYOaveS1ksSO5uiooDFAQ/cQNvkVwHzx4d46wdB2LpFQM8YSn
h9Wkkaci+jSv/uvW5GrHSmWcOGR7SfPEJEN8zYc62DoccC8f0KeaFfha/pgi+Ayc
+nEoiHDIrQDuZ7SshEu2UTs8Cz8R+HJ9QlVpD1fCzTgDcrIvVkef/yTRvjBs/usZ
fLjV4OQn+BoRlwBLXBmjMjjdEAHlIv8wI+4lKtACcYWYlXI5y4PIleXquC9CH2dK
x7pKbTVuc8M9804lrt9wD0rmtvRpq3BuatL63Y2784VdDUFNb4jMLHgYDYcx6rsj
aX1E4ofNYxV3nSnS7E+EZWBUPJqU9lNJ9/U8zkmu9GCrvM75cHil/En0U7ConJTS
Pie1liFgGjtdoghXA99cD1qTxBH0fnoYviB/sGhI3pKBRKO01ckhdID4IDUfDHR4
sMrMAWZlNidHyWxZGsMtpRxIrOMrNQeaTpC0GY6xsb8/2YHRvGs4/wxQ4L4DhR9B
s5C5ChvqawJV2EJ/6yobA7YpMqfXJsPpU3i8KBDKbAWWXo4MX4P4CF12G6sv/z6P
v+bV/mlxkQbuHjLVsyzymn6Cce4pQCfg4Kz2NEWMQPDZtaDWg70ssLA5VCq5mQgO
ypI0hP8VZ3+f34W/bEmBU4T2/dTKdgTl/RY35OhK/gFGB/2zIe6/oZazX9iUQe89
iuSD0LO3r16yeI/Qw6m1E0KzLBplMS2k/yYNTc9P6s/Iz8J5tBUsd9K/LNfOY2Yh
600L+gQPWj8LUXxl16RU7YTm+CH6crnh8+iSOqlD6dxqKU9y82JOeZHRy/gYKWjm
rYetwoTO+GqgsFynOPuujyNtxLHbN0P82/MPCo0M4/Y8jC30jsdQXRGNu4+oIkHo
5kQUju0WBBeqrAFO4bgRmFzvJRR3puHcpiaWYO3fQgajpKuSSZ69xsNCH5JsXpjU
3KgdqgoF2DuyNuJitiszQOgi49k3gvQPLjvaNOU1hbpmIxu5ln1JgSpDmCB4IMy3
H1B3NB9CDmf7cKLmt3h+LkssQseVgZg+1LApdGyrypL4Mf0N5NOPQn8T2WkJrXQs
i43zDdvGULI2s6PNJWyvuEFy037j0mphadBS4zsT8QKHQC1gCC+/Z41BHFoPwuvV
opfC3nHwDdWmp/9QjGY3qYz9Cax5i+IwqUi8j/uMmyU=
`protect END_PROTECTED
