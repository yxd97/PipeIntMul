`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAWP/wy8f2DI1R494TrFSClUdMzrGoN08QLWDp1qhlr4WwbrfTojlXaNyl0MwTmf
cn6OVRMDpvTB/BKIr/9zWvwvm6Qfj14X8Idyq7wTFwiR70nSRn4l3LUz9A/hTjYH
/3PpBVTIXCtd1YxLq6mQ4mlxK8YEZjo/pXnko3vIPiHkd1XlImZ5xQlxPDD5FZq2
cqLuiv0HFBIz5ifTCbEmbjx/gpyaHMw5WggZoJentyPok1J9cbYyS+pioMgZGL9E
ynCSRKTc/BXroz+amruv158S2sa53Lpi9Hl8QoPzmmbXcsIulfgusao05469sNYv
/O2KXrebIPLpRezsvfimRlEjBhHWfSjmw7GZ34iALodtUCHgcFsdZmQ9Z6KV9FZI
JjAT53owPBZyRcw4Q+zzRgarhTHle5Tx+BmvWBxZ4BQVTjEz2oDvzgX6QS4gFTnC
ysN2kb14kkUSJXW7dCnj41c1qFJhbnHOPWgfkzwfNRpuIxxwzSe4DNGFceUmP2WI
XVaZRo4gnwaluWfOXbj/ltiOiUk9N6uR+S48qFB/034exDUJS+gNA9iJFakkFHDQ
FZTeFeam2tK7l806I6yBR5BPa3bGELXDPquPKJxhnAQkSPztY6bugEvzMfPSJ9km
jCXhlM7zYm5nIjbFSf6X9CqTFS8B3S7cRhLLTtMpAvqVXKLQU64/qP3/qLMfgFJ2
KYR4KTac/ITTv5ISV+flHCxK8AnP/FZnqwHxNlg5leLC0UswBf4I+9Qh0DpkpkaG
Q7wum3d85qvPnVAF1Ri0qFVrKo3kVr8YysCypQpWiR7jeIz5X4aWZi41tvbfUSVz
GTu76vyr7CAGGfTJoaQ1TWZn+2Jj5+Gl387eu4lWPlGe0oYOF10j5egaghtullQI
j1dh7Df4YiPpnT3hE30x+G6QHryygOcwVkojO9WqBxxf1dvPciSoDJhoMGkfF0kX
MrvRYV1VVNfO6rd8FwKXQIJOhL29fKmxOUV2DGKx+8Ymli3mJTb0FxFHzoiMYtFJ
5HtlDb6CftGYKk31lNFWnBqwF4J2r+INDla28/SiflZdo9uqWRIaAQFSUTLqzy9p
3m9AmHbH6v/p03xapf4uS3C3DasMahVLmwzKTRbh5etzFYBgWlB/YmGWOR523G0z
T04i41uAzLUhmt0knSQ5SggShZcSq/OThHRpemsKzHRbMJSv4hBdO/NMQea3RSbe
eFRwhQ1yCATUS3F8xYVe/7U0N22zwTXWnOjJHRBA/bSEWuckIHIpVWN7FUSDUrWc
NzmTtxWfVwnQtGdACciHLwuanh3267jTiaaY9xT/gLPMrdFpgk/5TuX5evkdX6Bx
Col/KF8fQWqMmfhcHB9ukMSYfrKyiNnhRUMju0Dkeh7V1JaAJ29hczOen1lZzhWi
XT2QNyiTUKQnKSjdAhbyYd65caSdHg6ZrUtnN4Allm6DSnlFyj1AOKbEzctqtJE6
g+zplvN+DTN1Q9jiA8CeNa1iT7SL0MLhKlnDtXv5ghowb2OLB0JVO46GNSNYWFVJ
OEsAKRdX0HD/Cg9+vkTdCpuzC6GCvSa3Nm/yymQZn+CWvKYCtc71HZYA208CUzrn
6Rj8dZPJQ/K2Rav8N4GjivVfAuHN0DBZmD7V/7GmLGhZT718J4B78hPmz43N1QOX
GbJpP3TS+oYMlm8P+GgXsrQ4FcXLbOFxx1Hf7/6ge+3S6Z78L/zOeAfkaoB653b8
dXVxXMk8U40raQmOX5YJnZOt1BLywO4nN+tkXwcvI1Dd6esG6Zy7JnXoSgzPitQg
nh90OVKK1L2oeU3Ovlm8rQVvQYVEvRdUcJ3jybZYJ81mIp7Q0ADCjqNIwixvvSI1
9jw2i7d8esMyZSPVDk2rmscngTdXtRc0WZFiktMHCXdvWnIPZYyBfA4PCi702TbD
hhzCHlNTuFgs1rHlNDnzvJ5ATLRTAazJpLRVZrXaW525YT8Ue8qgM1/7ztBG5WIM
jA1BECdOWReYJAjFqFa9p54/u5hFtU5ktXXBPesdODdHUmdPLecJaUq5TKm9Y/GR
iwek5bECNcHRWmKZItclR0PzROiPgEstVMKVlGSpksCxzf0wQtLlB50IbbIzJQBO
bctwQOV60Ta/df7Il5wvPWXs9XiFP3y4iJ6muLPYfIV/Zqo1+qdR3cEGlfpfsRdZ
yfHk4WVghtdNilLNS7i85lhrtRTthGEXwaXM9YSfOtoIhKvZ1d1ok7WYuTWWSRy1
TVsdGeSDjHdvlN+iSfECnsuV3yiczkhvVKhMV12Q9JEIepm41pgy5/0svT+dyrt7
sHlqauC08Wxd0mU8IEzrduNmGIJJ35uPa5MPlkteRqsKJ4256Y19jsHYBOE/Mx8/
cEKoaiwxbqXF8jHImK2BUi1699LxcRNIdRAJLC3wKtvHe7OHIb9uXnlekW3bCTIo
PT8+4POwiux4y1LSpr9jA1+fUXCaVBLNS5c9MLgdKTFU6XtDwNwsePcjHvgEd21e
6cDoMe5JtCOpdbxqowiPnCJ3JS2nqABDoSQfwx3O+URspjze4og5o+bbH8MICF8h
HS03COoOiNMFBVTXejYMYvDTIaN5HfgA5JcMrgseuCs9+ndb7Nek2YiNIKFwJc+6
DvnktIMAD9T0b4qtZ+J/wb28SPm/f+UH5e1uanr1a+mv/TFfosNuOhMImOW6jWlM
JkUr3PYWrJKhaJU/fjxvu3fWnKdoejl8sM+u0DLdbUVibhHMMWuxrbDNLLioz+Kc
kwbikchg9uaz/Y6NBoM7PcWIjkyaK7TLuyLsCZVQtCKFyhsHmmloohH3nKRru3ah
+m9lSwA/NA2nM6r7O4U2cxOskzyHbDW4IgB2rgojj3qUnVclWHhegkF7T4uv1boB
0IUN6IHivtjkX1J+cvseQBRtjWwZLefKn+ofMI6xOPkq6lRiN9xDBoZT3gthsNOR
jg1k4+h3pRNfqPr1mV99v/uR/4b3eTG2XJ7J2Kxy+Er5OWmPVRz6u3NOc9DlADSu
q42s42ang1DJGjsfwhiNbMSFTy8Vug1yl9xuWYHjqz5gIVCUc3MKfBWOSHD8tChM
GzGaIJmIPaaHFnJB8E0ZrNTOQlRMRRIti1KBmasIdus1gQrpGgr6trjZu46DZlQf
6TnSzQXEh01ghihRLC+V8UkBwOhB/d71lYr6YcWQvswWX6ZPyJWbfa7in//Rckf3
61kVXFcWUQf/cpwbrDicZFSYfiJmRNy1ojMzI3DAS4yc4V1mragcydn2QYXZ6RZR
QmrSrimmlyQPLTXspdHhS02s/UxVQaQ0YDgKKF6K2elk+7+LmslahMmSJLJsXVPG
z+AWjaadO01A7CL9gDGd56WSCarTA7jKOuDSzZxg0/tFzrVoD25dD3zLBVewoVt4
KrH20UCL/PPSc5D23todwTnj4Wz/mwcoS9nxaOmtkFgpiCIprSrGkf8CDJ0P6L3m
m6TgzTErVc4z5/9VdmOV5PxqUGkL4525NQHv7UEJaTU0PNVeKT4xUiUUdvJcvYRK
GzofKNpnOzcownJO00FgPAD+oBhG/6blzy9J237x0gPIOSDXD6OfvOjLkpyJ7AAS
2d8Y/cPha72ELP1tTpmDoMH4JsFRRNzQ1bOHSUE17ktBSrbQdkbuW+gUDwCb6g0z
yjWO6aChquibDZ08MPlGwgHqMCz9e/CM70aDNGuwdGJyT1x1F23Bb+j3PQy4aKFW
yOZrAWnrT7VhA8WcY0Q4RQDMVmu2UujSP3/G0HZ90YbTl5ussDg3y4SO/RJsbkSY
fUJbJiEazgtXHcoWS+Y83GYnIHwFjRuF6SjvKbzRoFhSo/ppoVDbqUfZhlLvZ+v9
CaoMkW3afy/fY9eV3Zl0/uip4RsI1ZxYy/6FbRH4ZRgDueFQV5plwv//C9AULBSG
JQ/pCXE3XGUxQMqC981YpqzgPq/0xvZ1VSGXzd0H7iLo5NdYch3BnvWvB9XhI+g2
fjcghxt0n8B0qkovzr/XZMBfzn9Lmvc4j7kFwWoDmAg6stcMCHY+pV4Ty/SnSKIK
clwkH2qdU0cnLS4/g2S69YfV4YzoCp1LtumSYrjwQZK/CmEQQY17CTdQk0s7pCVV
VArZkr/ThM9q3V+PXhWrjtvMo6OK6NzKcwJB2jY2SuWXh0DImTBkDbA4AaPi/AtW
l2zDITofvNstZuOw8B+CW5oQH110tU0XD8P4n1+pZDBb/w2HcsSFe0yfP21MonDT
MZEnbNagpSfZqDqgoFj8ey4ZiZWQEZV2/4bLedlWhfhIljZu7vbCaeQpfvzXOIok
FkhiXCbJ0e1E7AJabY7URjxL2Gf0wtmPvXi0OFmwweoxmofnZgFlYY2ypPzeYDLT
KkcMKXwCx9T8QmchNuaQK9ovE0pT6mZsVcj/BTik+6VmtKRfcMTVCJxIK4b7sjCA
byB/lwdmaaPk/POMffcyJdnmhk/39Ah3GDicW2AciFOKiYp12nH6MZV86rZBDJF9
1V1gtZF6NFmlz0XQXMa5w9sJ8leCL3K1Qnv7IxDqwSqBbrccFEcQh7QvpTPVlyar
hD+EF/uLhFaKERkdKeLGgoiBvhUJxbywfq7+Y24YfZ0Aig1HWtWrsypWH9+F9xOS
yOILBMflcjsPL91m5kRNBQ==
`protect END_PROTECTED
