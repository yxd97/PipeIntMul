`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z48nLk7gUdK83x9k+AlfL1lK/YeodJTodYSH6E2er8dbUF00t/8aDM9LUtx/cj5G
nBRuvRdM2Z58H+Cp7sI4UArx9ycaoTBS5lIK/y7WSKwByvpbsd8AEvzGi+7aRTAR
MWmluTHV4rqEYkKc1Tx0XqoR9/UGZwY6pmRwwMEvqqnc62UEd0vEnPhdnTY5FDmN
9gshby0q1Fn3WANtLYJQx2b5VVNG5cxKi5dKQCbS4g8XsRsCeGGLM3dYRagG5jUK
GIQItCsJ0XsTuWC58LXQBEMVoUcds+XZE+CooGqdYHqCDZbvtMAQOGd3xkskETPD
JrKxeI2MbaV8MR4qCzl0FGkbVjA18csHI2mZGKI/qhlxRgOB++BCSMpztxDVecwG
xsupWiWcjRNIdleJQ1ZGAy3B2GUiT0CJG6WqXI9Tete4f8B1qisqzLvhgyyRMPZF
`protect END_PROTECTED
