`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iSr86IuzZsrj5CaXYOQ8bfUbwSZNMbGtBwjOXHlRAGsnjk5T/jMf4XCC4hH4bzkr
6QOvuC1WW+dYRBXH44aXcO/M9PypaIFn9uqb1NPFYVepVmmBiZ6AmNSq/dtaE3C8
nrGjdiWjwlEbk57yjmL4wAyNobolZ2CwHMZg5UjmM8iB99HCEgyS7z6k2DgJUwQU
DamZ2sgUkj7at60PyhyIjZJwBV6qRjeW0QtBW5wpiuXvtHxbRmAKvQDp61qHAzRN
7CyfRoNDYQ4+AdRiWDSSmpUwc78Meyc6PICg562UPCaY8F2ZU6el9GuJYQjU6Plf
Qkn2icYLnQckSKgaxnUamiSabMfcWogqtuAtUPs3GXbE0WPyn+GcqPTDB9puHJRF
2bj99ZVV+PR58tya01WIgY+VMDLvNqC/01j9a96eCC4=
`protect END_PROTECTED
