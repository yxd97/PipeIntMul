`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cEcPi/pZ9NwdAjZBy99xx8SLq1xRJKKU+AEsQAdMEFEIbpZ4jZpAeJk7B5KnjVc2
NgItblrsnPXOyn9MPNs9QGw+jvWl8hrhP/hsHpSe1koBNkf7/1lpQ0Tu6GaCaOQf
2PIgjtzBdIhKQPXIseUdxIc8bot9eaPvqlIr3+wHSBAjczf84zrUkjHZUZac7z58
DpgPk0UavMk6rT+xCt0Pb1+wr0IBuA3QoU3cwIj6n6DWHYtTcnPrqYeeQvAZvdTV
lC5eQttjLFxl+VyKrXqvDs8NB9hzNpKoxjgHWQIPz7CjMTNfyuw8owgbpaFVlXrs
pY2xjN5OmBShnvzEM1CC2/iYZMMeAABZMnrxbvPh3xE/k9Lp6T0LfA4DQFl6O4x4
9qpI6eVd9L39Hbw2Pfy6rtd6LtP+SlJTnGwEqRLDLlvsMeDvzxIAe9ulyWTIpwFT
jLo9+B5eNzKuUDBplCQ0oJrXfV85csRV39kJkyrh4RcDGahfmzBKEy+dR6866O06
UTmMZ/i1lu5LwwuO9VfGAOcvQFrZkj0UDMc/2VKHov15dzowENsE7nY2QsTRBdL7
NaEoX+YOYwrXxrhW7yz5wg==
`protect END_PROTECTED
