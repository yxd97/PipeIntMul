`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gtv70fHaEvw+JN1lJIzRiwgJS58XW7AyiNsfKlMNfK80lhYlYMzgRGG/i0Kb7tpm
tkco8XZCBQp2cvwxsSNcZM+nfiiDKjsq5wtLGjMaGrAcMaT6P8NFA1gy7L5cRJt0
T9400vdpHdpwZF2pCTjx42teXO+giJr8O9HFiJNK3THlZTzjh7SEkfpLuOj+oYiW
9YyNv9whrqKqo0dwKCg8SubRSaoR29ycSmC6HLccxWhIZKwTXU7IqqVqVOSi5qMH
Yp56siPGLMtEGE+0HzFoPZi7WYvN7qkbr7AttPF5zvsX/L12Jo1xZOAn2yEDnmVf
IFoAZ3L5TJMzL5rlkjxNqRves6HoS9L/CgZ2T9ifWDKHEy5RUb0ci/J1X1l8x8+L
Bd5lEck2j5BOSW0OZfIXHFLh+OVrgexXZqXV8CDV9vYVTzD41+dckicHZZ1BALPW
F+XXlM9ufKUqa+D+IU2TwzxpBhur932ZLz3qmuiyF0BKqVpih+iYlGMJIMzDskSW
VIxC8sg5v5kkyvxTmZvHHgSS2aEEm0A9nVGPAguGdgZ+9zZQv36EzkBkM1v+GMsf
NRb/rWP8PrkicuE4QVRGfw==
`protect END_PROTECTED
