`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PYHWnnWsGuhcSU/BcxsvWg5FeYd2SS5I1SJvPP77AHbl7jQ6UkvIyEMQuPWmQyFG
08qxI9Wy3LmWKoSfLIfVklL7FKYWTCRw23tBN1hqIBvV0x7uQFbhL2ge0RCeDfPE
jXFbv4WcNR9xHotLi8cfkWcJlDB4DspbFrTrl3E/YpByTpZr9SJ9VpKia4bbMiN6
45eo/qpq5MgX6A3wIYAde1bWLfHvUHPnEVKlahbZlrPS280RhwEY2cY6vvKoGEn6
jORnBvdDOD7a9dzaMBhH7YWa2Yj3X1xux0FoF99vaFuSolhgIORijlCjHWZRciAm
5axl8uxcv+1z/ibIZwRohbWeDfb2SFLpls6hyPgDJGbg65Mxobah20MTRF+WBKqR
U2X5TRSYSj6oOcEhI1W5Lg==
`protect END_PROTECTED
