`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ziiyOyuqU2kCPth3JGav9sZKDCbK/lSlqIpjOrOO9zu8RWY6yiY17lPGvX1YuFr
xtbRaewkYXZGlHFVBxbaBlk7uz7XBi5uZtD7YrDPi6jjc8HxvqVPoLa4P+/ghaCa
lmXXPnPB9m3+A4MVYYuwhQcxt1pmF/af30ao8Scl2cf3cQTRP19XpetV3NJkDhZ8
cnKRR4FqUrFq5/b28x76nQ==
`protect END_PROTECTED
