`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s4ROpRcqVfsfdCqtXLb/S/cgbMUrjSNNonE4fuA523oEwv3jkkEjmSirCH17eh3U
9KbvQkn4Ym9Um3KbHW+lBVJ4Nd0iLJfTWaRW6IBuNGfQ6oP5dVpFHmkY7pLtfaoE
lRGqTLTlTcPJPvRAAhUkiyT6+L5b+VXFB/KqGGa84I1wqcgDdPiJwWOGINHweEO3
L3PzE0E/AQTECPld0za++G25f/Bsj78rfVQtRRskOe2jbQ+4zAT5DPz1S98iybyi
orS8nBLUPQCRG9kFfn0HVqvHYedMhtCThnWL3dp55YTdq6mHX5w2mWSU1znuEEX1
bsq5yvF2nAc0w4s6IQAq/RlnVWZqTzIBPV4li25q0Dh9kmAVc11oZvLAqQCL+7Lw
kBKhxPmkg/ckYXE815pk9ibp12x84x1K2BXIvgjk7KM=
`protect END_PROTECTED
