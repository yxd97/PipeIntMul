`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wKsabxq8XUohbYYjooWX9GYQ7n65tVbt3V+qDU8hFRNTnPn8UNMEavt7jX1R51bi
mPShfkpTkxSYswz/u+C0TKRkigmzmB3NrXpjoQrkMvHf9AgFkra7eqjyGol/MRoE
rcGsluP9tj1tDihNTcvS2Ys20/l01jXPXlp8ceQtzFmJfVCzZIWQqRc0h0O5mdXJ
isuLV5wUDjW+q1EkF5sngOi4cFhChbBat81I2iL7+v1WX2Kh4oLfQYuYOp5Hr66M
j+uVpX05oOdan10cy+OKj9wXbSYQEgx6zWk5egmtXbLZtKVRSNfiAia+xSyGFB9a
Hu6tN0O920V7A16an7/G7HFzihdITGrN9OCUXqD5jo/e0LtaWgBFfo5KaopAwlK0
pbddcXFb+2uPqkmuSYGTB9SSY9EB1nyzqqm/b3HRrJDPosj1KJIQECLjA7n62ZA3
lHe/GJqrYgh6Z592PHhJxq6fl8DFxaxFwXEbhnPvm56ueDz+xudnES9zzD6Z4MLg
wkuFw5I9LaTG8p8Rb8biIaPD1so9g/EbO1HLkapfy5IU1MObSQdS2rCdpPxqqT76
glBtuliig4Ez4gh9TroYz/UTAcI3sSxilVvCuFqDMRpmET5/Mz/AYYS7fh5KOXKz
6mH6KNDJ0tTsC9UpSzVMDp4bbZZaS4OeNwvxIc2JjK5Xh+rAMjHPjx7mzURWaSj2
uXhwPgU+eVVwdgVol8qyRMysfjZNpdbYe/bt8C/0EimmpoXne/CjXVnNiYfJjLi8
HhgLvb4NGAhPk5HgphH3GcoeRqnE2cl83HtPoB3Bj048EBfqID+hk6xNgrXPQQ+t
xkMfKFt6BXTICejMDPp6m7QkWrsFzVCIByld92nOOrqEojP+l8Lt6bdIgJ4rjbbu
13ArDjKtn3VJgo79wSzn9okzvok5/fxjQcKuONcv6NJXdj4iI4ZMdWEQ8qlgK+QG
kZiLuZcWbowLCvPid0kTFouBHG0Vcbbj9KDSrQGUpV/pt+KokcTpuipzJ1nQCiQ1
9j+5pTDyRYKaoWyWUobVWxQaoPImihA3my6xbp1QewIAjYPz9Hnp2qnLxDEJuxxb
X7GR51VsobfkaoBxBRidnKKqrXaS3ZZd5D1v9jeVSkh9+lmt+yA3QeSCbtlL9P5k
OFhf9xVoI7aV2+DwFZD6NTp4afintGoebi239fCu4/miUrLzrpty+eEWQWbM584A
Sx0LT3dKwhGLNZuJ3q3DSzjeiBBy2CVIgs/GJeMql4wsh1RgmVScjeU9hWUh4YEv
irPmqq3hLjD9CUE7KUvcIc0r1k2I8xRcnpAXl2JtuaknUffFyf2jAQgz6qcsGcRJ
UbDh4g6AxFoTjPwhTUZOvqz1JIGT9y26x5eFuCt+8a/a3WzGTLKwAvppX4u48aCW
cIvaiW9Aj1nkqYqJAbhwkDPuF7pzdy3rk8PJG8NVxFoQLpi4Q7U2Mm24pU3H5B96
yw6F/18Q+cV0Vs3Xg7/ZXwmCd7edi6EQqoJ4g60JVoXjxuFkguA75wKWaT+vIzRf
9sb97y1LCnszL8Y7/GJAxakGl9JPMh6YSt3lxA/zRczT21iZDwK8ZTuBEbnP9J5H
yThOtsbOzTmx3nQBISaE7txBDJx2NH1Gg6M90BDrcb9w2RpHr7gYRwpmw6DM3xqG
1GBT+1YsvAiHlEbxq0hJP7GgMcRftH7fhqg7e9gMxpRTpFxDfbtIHfvkSaiFHh6h
fOgf3eWmbw6QPJYuZC3h4bmdyUZB5juIf7BFbAZsLM90Lzsk9QPyhR3UaT9s/MnA
xbOEj4J3oA8tEtJp7rrUMbliKNqX9vb2UyHmjewTA5aQ6OfHjWVfJvJnHjWdgHEK
7IeLcAo6ciPVr6P2A86TYjr1Z3nEvLh8l9djps0d1O1HGo1mmTb1QID3gnMBxv+E
pFgFQgC7Px2T9xyQoXLqWE57DP4Xcg8IGBnZS88dfoQeTUWM1yxt8HVVkk2mD5wV
ijxSq4lwzTURg0yvsw9Mr3F4Bfwk06359Jew4AaFEr9jcaoEvARHrb79avXIPT96
MxWVCX3+Asd9g6AE3r4Q35h/EyH5pZhmgI/OW+wsfbu/zichC2HivyCZ4oXCr0kk
F+Hfqop1mwI+Xra9ejHoG35u/piAkHSrLCkfh6ug7TyzC1E1QQR6sVcF+N9Sjb7W
2Pk16TESfsvryLAAub3KK5cMCX21Uic2FBzyJ+Da2S9WCQ7/wMu3TAS9e0t4r6Q4
bwl90Sp3hB/S5V4c4CMbrgCgL6C44Y5SzGG7ytQycqYoU6e8nkJSJwjaALT45q74
sYamsquW/oSP3Cze7lCyzAHmRERCLlnLypvtJJEJAsyMBStM4bdj3JZ1rZA4+0DY
FfFSYF46xwwm4mOSRNM9Hxpjsbnp6WNOUZjfEzVQSHi2wjPea0FcFlhJpeD5OPvX
1GAZAJFDbftq0nxdb8iaRlxyQf/C7KT0P2vcXxX5ewrz7ytbM2oK3B+/mbzTYg3r
XzgnjgzV1kQg9YsJ7PNY1RHcjl7ntpduue/IhWHWcS6u2PJG9iCXohvbYyCSQQJG
Rrthrjro36ztJLId5zXn5/fdKckkC9qgM/DQ5EgkNFQpWQY14dk6k+k4TyQDbRUJ
NNtMpgWUXu8XkI677n8TsLO+HyZXej1C66pwZETyvwnGIK4A2g/7Pjx+abYa2nwO
K4qRMqjRLWSRiawPTTmCGJ+e3xRlUosyQuGMzJkS+vKZZWF9WbuFpgbP6wc/UprQ
et9+MjcUdTaV2vkKi+LH9vHw1ZZNGa7vAGG2HFXwe2W1ZCnPQTaafQgUQcrvjKSo
e1hFOjVq1hESnsiUdVbAfBAYqd1NlkgUCW+72+UtCAqsTUupcLojCnWlKe02t6Ez
fD1nMjW3qHgY+vB3XPGyl+rik+EVp1gHEP8UgeAgARurUFbx1z3fHNnmGIzj5VnD
nseJgWEbv1sqvGIxmPEEgpCGPRdXEDk8KNQ8MfAo0trF6QSvKeJdY2Cm+oX1kqgP
fUEwaZAFYOVuLdxT32krJSkwmXUtekLCT33IGwQyFlQeRLTQ0lPmrbZLN+MpCFCK
LeFdcO7NE5jSowwHGJmWSVNF+/+cSLEoIZ4Kew2lmw0FiPeYCd3zSS7p5RLw1NV+
KcimgIz9akC75HshBek+47rEn/5Pj9AhZdzdnTscAfM/t4LJKL9qh2nwSO9O2bqI
8nd5f2m7cv7DGG/FX8LM2G26tary9MnsZwl18RMc9tiPu1zgOAJm7VvCNL0TnxVP
0yuz0En71BfaqQO9NyThNtEsyKPuGKHoNQcjPaXXB6Yy2FZ2rdxclo0gcerAOkw+
1FWiwH+GviAkgIjmokEhqMoBmaLh1/u33L924aCY8pAWCHKFCMXAxo6b0YI4t6UA
WpreH4xsYPRX1q6MPwu0ltyuEjFfN/Y7/LfFiCNIZstr/IGgg3OKlYdJ52eVQ1UC
CSXhSs1aUQwEAHWq8Yuxp1BU34Brd3cLITmCAoMi6IDM8qzRhTFkJ+pk0ZkLDUU/
ytTlUUsFPT0PMo2s+6qFpRS+Yw4vapmriwPenuYJvUEunSNhWtL1qC0LAGZuYooG
7ouA5K8Nf5318L/jvaK7mibOEqYcbjwjKa4OdPTLbOu8ulaP4kSaVW2PTOhdT2Ua
R5bVhd1TKsJiw0jgYfni5F7aTKKTjm2w8R9xOJwUprsJ2UfN3mDUp2V6bPqTfdlk
IgXlRUHPlAPG4Czdd17liGL/7sMcPVL9W6gv01yyX5F72VXZCEI/LNv8fChDmEo0
E96Q/bx9yhef/+kzkH07Y4awMGlyHkBPNQJJ3Q14mhpBtONkrDpo9FXNe3IPMeYq
Xre6x8rU0jV6kjj/2cH+56/DBx+4mme8U6V+IOY79nvHgCQodp97asLwnjloHkht
owQgiGGx+Nj0H3rAsQ0PluAYu0kS/gKYRnxCw11AjLMcNqp4nYKvFsC9DArUuYG7
CnOdwHS1J+wMJ+jqAuXp6CAD0ISooXK8VPijp7tD7n4KECswHsE5Q6Aiy+UUNUL0
oatTLyDQ6VlXJVx9daEytoP0QYIkQpf/2mxZuEFH72nDa5cc/6lGtl16CpQ9Yzqc
w6/ffeB45JUEhyGA9mwh06dNpKVvxQXg3d05GxB1tmtwDFso9d+fNHO4NkHhA1W/
zbhRSD80C7pF2vPumPOlQYRo8jBufagHrithY6gJFqvgew3TP1eLXngq0wdGIlH4
R5GS8u7FX7/flyIAefQb1qe2i2pD2GMsInS9IwX8DaZBrLrYSM85y9ypHpMRsOzW
gVF8cD+xwYfE5dd1HbvDJuSFoGh/Vxl6bKTYYlpmW+K0TUzzvVCh4n+qeWFznmwh
y00zBY21r3OArlk05VAL7hEY3fm/uC+bRDRZwy2fVoUTCNriF3PTVQp4kbUfpse2
EI7jDDMrfGEj+7AsocH1MP3uwjFgn8t7wrRWe0J6D+dLdhJWR+TBwNBjGZpeWmsx
NLQFy66HKsUZaeffJ3ULFJKHNK3A+c+NBs2y4YQI4U96vXq1al1ZYXfWRG60YfIP
Vg9lQUvqFznLRmJO20pDPmCRE57ok/xq2c9u5cj7jb3Nl98B88MwVWLgTiok3Ya9
aRILve0gfmRK78SkfP57EAIf5JA9PDAYwrPGn4ebNyfmAJce6RFCNTG7APqJYzR/
JrjghM74+06t3T1rTTsQvv7wS6/yWYTmlmk+6bGCMQrSqGQCwB3a4m18yBhV33tQ
xrv8iznLDKZ7yWbe9M/lnuUXhMw3N9ytfu6ryFgIqLAr7hkXUxlBRq/vXddwFSG3
Ik+RdFtA2q+vxmTps5qZSU+7ACkSA1TK2ENbFUYIPgiyN4j2ep6QI/YvimKTd0qL
ygn5xs/6Bv15oLLW0JdIqoHpORb46RhxlV1YMpUHX0BGLQqNzcuQDXVyKlUw29E0
vf48Z8KCGf/q2uk2MkL07fQNTzlsIe8nPk7vTZSdUPpRxdAXvXdDIQs7fWCR6SbO
CetsMBHhbIlD/JsWhnJmEXfAeMJHDjLJ2U1aoIPKGkLjSyW0Xttse5utOyuYHG6R
Iqs8uriGN4xqtD/8iko4c6mGWtlPAi2cK88d8FPjUbcrkLjnjs9PHPLzZYSzqs+2
5zMC8MJIcf8q9ZWijcGPm5YJ6rqMNaEoXgRYnNbUXZgVjWqbypCb5iFtvh8jLfET
4LYhEMXjRS+gWk2TQHNKQfETkY0w/Ghb8kprDUvZxogxF5g4Aye8GgC563Z8SMl7
1MZh2kxIwXUq7h1K2X5HemP92gOKsYXgBrRlMY6F7qIqxcTvB3M+44NttKdnqVhm
RmCK1wNJ2qCYyhW9OQXL1KuP8whxpTGrA6JXBjLzAWmBYvZs9rVGCPq+tWJ1BhZb
TrmR9yJjZBPF/Qm1YzoOpssqIIwLMaBPJTcplT9lo3ogyN1YAPg0s4nGcRRPTvbz
/GLZjgFoxVjl0ICxyYY54cjIR5l+005edS398qqiVcpDUFNmSReuHAIF9sjs4LnR
XGE3XzZ+IfO9BH7sk5iJn9wtkDMNkZPZi4pSwbQjCAmuTDHcsLpFQJW4KshjflFL
wc9ePVV4Os378eZjBag0ZX2rOsyT1n51H16JP8ZBLEa3tlOi3YKyYfdT5jd2BV6w
/s0+A37Umssa3yCPbLzMzKbUz/Fo/6+YhWr2CbLkO5Jl4CTD6DyqL/80IPwRHaeY
M7q8tn1Qwnh2yU+eHSK/t6oDXvnRrO3JgvWpHW+RpdztWpyhrWwNo6swd4+PK6oP
PQUaGKr7cJgV5GOMZgJZ9Vb4t29l3h/5jArZcZ8aiGN41lMQFe1DzqsHM8wtTsFC
KueMa2VabWBQdEWHqxUt8ic3GzDAzjUv2OfK8E+0Ju+CfWk9N5RFo8mJzYEZJLOH
BRZEfvBk703df5fQFv3lbyd3JMfOwbRhhxNEZE78jBzbyBsUtH4mXYU/p73koZaH
e+L3HvVTAQtAHgWaXBWIu6ewYvnR3qd3W+/9oKhwKuTC+NKKzbABK6n2AmUU+HU0
lYft8H3na2ciMTJM038Nj5vjasYx28Godz5/rU9MDMGEm8OJQ30c92r/T3u0KZ5W
WFV63hjp4x961s6RfacsqtRuOJ98u7w9Ue+4udFuWtSAokzx83j1FIQMX5N4QTAe
nWrcm0gMdGzA2f15ZdZq9EOlQFiw4Wb3fD6WKv9OgN50hYc25qGg22J+yCuUTMx2
GTl2QAZxESXdjjxYonUUxtSZvhZIsR/v4JHVKtHPrYJW3fADf1Lr+dMvEBHbqiI7
q5GhsM48NY3D5+jxtDogeOl2MpYL9xJ57lPFoKwstwWE0YaxxS6nEB8plZEqYaGI
EKmOBMUnpMuPEjQHS1B8mlgb4/lOxd6xSmOpSPYuU+v4W0pnwX5EFIwh07kqpaAt
kC5fUUrhRXFM94+bCWo1ttW+Lp995PBvRTfXrSQmSocg9GWVMxI0Ft9CzIyxSC4o
1YA0fPdjFRVrbRx85k9vILHFkbY4j6CwoxIOPFY97nx6S9Hg/m7T23q0JKLm8HrD
F5uDZXC/ji/66H8amSd7dSMXhWyKC0ZmaGoPFHvdFTQu9ouD57obLezSX4xQjbgc
buDfCM1Kec+9CvHIFci+a67z5yYBbSPPBN1Fde64A4+UZX+u1+7NThB8ww6upmh2
MX4X8WQwmpDu4j5gieCR1lrzPMWeOX4Kj9mT7wfgDaGBg4AN9WFnM0jjWCP04ay5
QPpKcMGr75Q4/8fUM1unKyl2hGoahGa1Ryf++nGNg04nWs/GJbiIMzjqDDr24l/R
f1Q+5Lp3NaW0hMo7n4avjRhUitqwzye3Oe/vQqYUx7LDUwCxgKKCfhVe6DM54dz2
ERuZrsLPlA5+ZBoN5dKsPN1WEvsslKsSWh8zG+m3j2bWATAJyUZ00eEAMXkvBPHb
mH1Dx8SbV+V/hUn7sKCDhNSyolNYYVxH2MK4qUro1ldgqhG/5tK7cHmAc3XX7zTQ
Qsoj7ZxJScVUEPfQbuoAavTARenS7Xm0DVyOiYPuxA0EXQbVBs0Xx17sQWe0UD6t
hSUdXrZZBahcbHBPkphCom1jqTu1weUaeT0APFeTrRYDiBxPjf/eilDqWlkAAyxq
oEqFf3CWVuGLOAqV2IIS+YNf6WpCnzR4clshlqRl0KRmL7x1m5rOIJ4uyAJod+YC
EYOi7dzd+y6LBsNT12BXMTx6F8m+80n3XptaW30CCv/jas7oZAFfyi26/8DGQisO
u/NQa7JV/VXvJAZ6akGHAW/UYAE82CuPJX+iR0aeMGs7ZII5iEyem6jlKWSEtr9x
U82wY0fAqdUE6VftGaiG3IKST9H9Pd26PYf4AOshGjP2Was5BT9TK6CDeYNvq1VX
xMC7GyI8rfhJkfe+1bk+Iok0/h9a39VqsJL3xKdqvG5FFYA6EshhSvzsy3J7hDn0
ANsLnZyQfVGer9e1zEHolLsTvi7mOuc0Qc+w4+PXMsHtZAQTLHFNWNT8wFleMple
UVJy5Xo2qnQH580vAZWoHQSaY3BkNbzRjkCyBjqbP/JoomALPjWrFOD38Qlql1aA
OtVAVpLT+Tk4WNsToBoPAGLlI2iBGLhsdzlATqnnAzeY1RC+nMwEY2NrmxZyP4Np
jw5fGzyjKet2NsJQpuD8HFtJTtbQVX4Az19vhsxW5vMqWYYUUKabtYMM81M3baiS
jwhN9nP+11ykg2qr4iP8qHtS/M1+5v0jul8igmcW1tkBE1cl/M5tVCVD5lCnAMp/
q6fDPkjBPYaBDW5aewUEWBIKV4vQoTicZiNRcUwbtUdhMvj3qgyLaDO8BsQV3KTj
zBWux5BdLY7NoBZxdjpwbG+NCf0epkpoVetuRcO5blZr61tzUHdTihk+n5DzwRyr
vWRgLevHq0+En7c1DwVHBeRfSbEJLcWAAth2BxurapMLRBb5MOT6aSRO110xqRtL
6dZbys+ERnkPUh1DBH+/yBPojMQBbgQhVqU0GYZxlC6dr0j/pqxwyMgIi2x4y9tk
N1Vh03uG7clOYOhLJjp6adu8MIco5AJCRESJ7Ei7VwlCjQlhfqo4Tiq2oOfb9/Xs
P7QgD9hgdWuWncmiUHmaWeJEqUsn5zvR6wCat3evn7ZcOIpdCNUxQklA/qfvCnxO
1fwsOteUS7YmMLE5BRT9OdStcK5Qa82DzOmuYbDDt4uhXIlIOkYGJdwdnmAtepgY
U/cm0yhlTg3NbJyrD6mESdaf05GWR7VVKznNVRTcP2+nXDhfi0CMdb7jSH569hf+
ApkzoHNlOPxXwk+3e1JnpaAV9eAJFs2j5eoPivxLBCt7bpMBhG9FTZYJ7V/jRGWt
9OrRgT55eXX5MfE5OtO/DD5oik2KNPHtaA9hOouw6SRiZB0kEsC8Fr7giVuPaVNE
w9jTYI0/pPPIvMexRnaesglTcb1diGO98Iz++P2RbuTPdQpc+bhUodFHMVVqmbpR
31qmWR+dTuc5gNJHEh/j8VdhoNvhdZ2HZce888LIIK79ke2pre411rRt0pOshxVq
IX0h4Y3s2nsE4zx9SGiLIP9BKvaoZj4xNH2vXtfiS3OelItq+QsIMyvudNy3JcR4
MlmLcsqUXZ1/Srhemz3WZQ7tmMCaaKDTI9v4RTAzBxQtGn6J8fanSUr1MGWtUyQ4
3T7vCaxacN+pewDt612UEfqfMgnLXFdTP/eg5L1wFBSGbo+YKLeg8/pGe/BEYeoa
mgU+0mI4a+IXG+Lf3wCQ9ZkjfcPj0Duj4n825Y136Ec3TfjQ6zJ7WD3QW3d9tHsy
hM/zi8bskF1qycjHlDo5/qib89U8sRrdzjhM5AlH+mErOdEpKMTmPoDnADRon0Rt
pCl8cakHyIUp+zRUZ+/moZdqXO4MmoOh6jswqHSTxvhfkkMlcasiuIQ5ugci9Rbt
5RtCizPDHwbqco715Jis8DEvX0YAwmXfZtHirH68UtVxoKyBWWdgPdkUJK5HMJXU
wybZLtcDqBn3AdCRtLuaModNFyas48Rter7FGtKsN/gz0Rtc5aZdtNEQVmE9Qbpu
boB0kWjE00C7C+A4TvrRb0rIsEUcC66JAhWtBgYLWPetPbZFlliaSzYVKWqqdO2d
aIZQV9bK8dIkTD8Ebsc30nC4qQyXHR/OZTg6/5wyYVX+34LrKAjZFNBCN2Gs9/z9
uoX0YEyERZXNTF40svWiIQeZ8itZi9WC1shxXN4tGOh8rcN7MBR+kBtKL1kNUMLx
L3QjC0voDEu/GDR0Gxj5eQZFy+9V83qaWfhbxkcvVkeoaujKZ0/6646xBREyKbJi
XDA2wpcS2GW+bNoLwRrkGqJSaIbZsdFnsAP9XsTpkDBwwfxP1SKct6qvhCPGpFHd
/O5NpTxn93X6UYOyk5l+0xKluFJ8YJlxiCqSN4dvzTysc38DbRJ3GeTRdihnyZTQ
jMIMUJ7Rl/gX5uwFAwSHrlMG6j+tpgxzHJKDASE+0KjS1+STJWrf93zB2XVAMGCb
d2EWlxyXXBR30LRYS4Diy/dfJegCRh+QKH3nso1NXjnnbUHPr7A6h26CRbLuHsSf
k/3ItOhHo2rYyYstYxc0lFxYraOM0EVayi2ziRxz/21H/U1+JcU56LZ8hDmX+U1Y
cYonnCfEb2k4E1Y/vbRjjn0LEjXWkZjlvmkOtNVzD/mRt2GtLUy55cPQ5J6k8ngE
W+42ZM5PtBz4Xoy43VPU0fMkwihUb7QtnfQ2ZxfQo/poSpsSxvqn16RZAtVWrAr2
d7c7kXJ6Xs6XG8f2K5u0gzvd9ag/GOkSCkWk1qzBOeyYsQUefloH2TTKFjiBQ4O5
Gk8FIVMVecC2uYkLlCeG8mggm25ZdRAY22VQDk2vtJhv/vKy49BPqwe+b3Go4J79
AVaS9Bl6uKK22djBf5tDKKyRXJbYwlFhP5ECCP3OaUKS/QuWewmLE63Ewktqdgo0
0BGydhLwYjW824dQhRI5jngAxouG0eekQM2LHruBnTmbfi873YuUHWwRhd5VEmJG
tuUcYrJmmjxP13W0nS9nNuKqHDhRqbFE3JKeErKEJPiW6QUW1x3iM4O2VNtHxQGr
/UXw86nvkotHUadRQ9tb+hl7CuWXcWQ9wqZoix87plkQYpv1IaJiJrMRRGOSEzPS
YXbt0yu+p5U0MJHSIDsif4mFlKcA+UvElCYFdaxdeSI7oaBciDYgOd8NIOK4/DWU
OwekAlvYNiyQiA4w28M8zm3Zz9C4KUVbtMMdG+FjfqbsS/jx+eBOCx+TEbhz7hYh
gh/59u2O0J7x2xzTbWCh64h1/JXAVqDZkhLJlMsiLUmhzxKDQGOR5WbMOt3SWEIl
oIMFxoT9HeAAAJb673WkHDHSHxsV1d6efaQaeOeVppx6vq45TUemTGsDLZHjSvXP
CMEG7vDWN706WTSy3GK65FSVs2ydQgN48STTVUvs+RLs/8KUPFFEHYksl7aHx90I
dxBlYNNsYQx/keZ5bGVU5/69QPs5l8wyBQMO4847QRWA3foDv6HEHf89bbgfTt29
rCMEwZU2ejpgWoJ4cekoguHI/P2zZY3CwrZ888jWXiJ0Xs5alJHZV68JPuQRQKHW
8qqo0Gt2KYpNRKibv8C8kgbRiHjQgpC2YaZts6kVzS2ZCMRLzpz3QpJaPXue42Hz
UXxPL/yXRir17pk13O8VBtc5mutdedNRaZwe/gW7VfA5Azpy0tGDM80nWUUlS1+j
xthdpuQfRB7gPraLgjwmVhgpTpXxYv8txiiTPQEQvstFsEF5QTOe+mvBVKsnd+bg
3hl3gTuRXIoGiEKSD8LqchywSTABUM7U+Sk91fPsKg/1c4BgLLbCop+ent7N3d5c
9zBkbhYAnnVXcWQMqSF9A9ddL5kFEoqGkWo8UZ3OiCfnOo0TDc8wNyYjbJhkr90B
yRb+TJfh6J5/Qi6m9EcH89O7prfQ6glpoq2JUQUfTdWu97pAEy3YAaK8Tx2hZDz8
lW/SdRe492HJGyKgShbOuX701JZ6DbeJLc9UdiaMGjIk4t5kC+lW7tfmnOsjB7OT
a/5vzqPDT0vO0AkOUYQfAKKj0VfqV50baoPeutYMnDHEIdUCwkRsNJNEdMYMFsGK
Jk+ug3ZXsFKDPfJxYHkCPRRHGC8lC9bIzxte/Pik1E2cPCtgoURMrxmBWUt0FDOq
19nCk8NnoXwDAWp9lTkHtWHQTScpnzg59Hfk4AVIVrBEEE/vX+AiPJ/zM/NWJg7w
gOjkkWrvLgtuGTyjRWCiW9R4U1igf5+oRE157RGVYPLWnbFz0EN16cJYTAdvzKVk
B2l6Es7f6t2pFiL405/2jqdPa/gd/2h5ywHlQHOnMtuHvYgCWH3YOFgxSc8tsNoM
3H6GkAzXawn0N2eLHOC1kLp6GxOaWJMkFkORhMObia0wMSRjXd1fLYFEfS73Ekhi
8HUggQFPSTWUeFuYrVXAD/ntYNfxVfiPrnbjjGgUYj/Zud1asS/MaxqTyaKnPgBP
BIRsL/1WcyUY8aB/kz1roPq0Ur+X+UMokMfvd3oildjvU0vu6u8xacboAPmZ9YpL
UiNzQdUyoKZs6DB+9jZ7NHT2IQ5iGcZoePbTYPaNTSn6QEYurfBfhbH5h4/Mx25D
ER/jTLaCAqNExUuRXstVYkqO4SjHeNczzPMLsu4ZO/wCXuRHlDHCzcf5PrHPLyf+
Mdk441pmS3nJVZ53VbQ7YBO5xmvMuzavmA3zX4x4yKkbGTw5KS+b7TEumkNiieQF
VmufTwOyYhhWW/WERXJfLgAJN86Ly+tzMpQNgzdfRXzWRD05RuPDs5u+9latH1nx
OlGAhjnhs0i9cXZHd5Ssw6B6pHuf7qYh21LRqA0EfMYb0YfO0hQ4tYP3/Xk5Pg11
Tsx407aE7eI8v97Pt1VWPtkLINKWOtkUvRJ4RVaK/zvoFJMyKbljpkbrqoAnyNcv
7eHP1KKp5dtqT7fUEFBhjR/E23C9jRrEUULWoryZZF2tki552i/nC97U0UNrOIJk
ZMQh/Tm9+xsQBwhM/yZU3zia0Hr6pFlB1u/YPcAD3IhijAA5aoUjn9rW/3BDWJLH
RqTFKvP65gNr8oIGJugtr99Z/TZCoLywHxgfTurNxpIjD00UfRZAkHATvFiIEnjm
kN9iIOzQG8x35np2TQSYEwbeoMm87sBfBIyOHbQu2fSAVvAlV3+wIxM+/Cx1mKCt
+tcBeC+YmdTt7PScYuTLHG9bq8nUcKxHaJ6RRQ1Ggi6ivDd32v5n9F1tsWnhtkXb
OiL426vWpMwHbMaiqtJDCCImLLgHsfRaByB1Cz5a6e2NyNUrKKotEBzr6sCIncxp
OVs6XKTAeXLzlWMT7tsmcuFRrlLqGqPJq0+3+zrI2Aq+l2TD8nXt2o4gz97AWlzO
CMBXU61QiN1it/00xmTqqEzB+Ic65ekSsfcBvHQgC/OU67Qi/2jMU2xNFHq0zclN
9p3Xs84VZVouCINcnKjH4A3/d3uhDwCSF43xVvl/kjX0VR2mWFL6DERIFswsmF7w
1S+5k1rawfqsNx4suNa1h5pRdAg7AINiboA/20K6yjgkIKN/b3PSZuJEW6uvTJ2O
4o3HqD3t/ea/hegpcSE3ry0OgX/dc/D73LcXKbwo7WahIPY8kIC/wgwlMY+GrY6t
np17ns7laVZSAD7u7FemcfWTrMaOO6tJ9vuDikF3xcPdKmWj+Y5FA0ILAR5jsASs
UuVLaQ2uDlbhKgYULm668xNLEjiK9IEOKVTAq6o4krTTncJx6B5h6dn858JvGL05
qeqj7rBJfELS5fUcYUB7DXN+xN/kLuZGT5Z2HJBXMkUOaaOu4hcEymsDcO02A9QP
E40WjUH/ev6bcTNyFSs80BBv4DBoe7oQQSPf5iUUGkUviF4Ea7QshSC1ngCNPVKI
LG02echOBuQPCq/7oqNeBsknC4j8GNF4q9FHDNa9Aa+USZLsujAnEZeNqPQuKX7w
SXFsliVRJiNmXJeiZBoquQXkzdAohX5ShFknUnCNd2RnWjYLRCQj/xs4TcO64Uuw
ZkzXOGkDgEMYi66VlqOiv4Heo7jckLaPpwlPFFkBq+iwS7+/xzQpcdtyD2zEwZ+p
WAR5IoN6RVH4iO3FX/GBP3P7mgm3P6sxpF/ck7zbMMgC3Y2zZQnt33e9MgNG4DIc
J/XrVKKwvABlmv9UKmtyyZmo6vOvBfFBMu8eni0L97I02+BenZxpAAyMQu/TPaWX
h3J4pYQUu0tVTxFkkP6jPvCqIhKgS2yLqUH3Ja7ZfGfyAUzWV5tpgg/FYdYirG45
LNTvkMFyl/8oE1csIU+acCLrbv9YsMNYF4QFT1Qx4xIVNK7QBfeRmOqcUwaImBOo
aa0mkic0+M/AakCuR+sIgfqiqZBpwziM5pr/JkypzpMuRH8oG0ibex2pGt5UsOMC
0HG8rbSVSCYlx1PCGeAn+hZzNm9gL0hkD4N1dUW0XDidN+k7sNB4587CoUW97QYh
O/RQOONGpAWG9keNPEpq72/iD+U2RairsNCJgGWo0+Sh6Yr22/E4WmhVfYuUzanm
4/a/7dQsvdnpZlSqcjOdY+3EQfcuXL5Lp9nIBK4khuNwVyFV/gVYsLXnnxGACG2Q
6BFbvg/YbwFiPL5wA90xvK4Iwh0udSp/z52lBTcbKV2zBwmdXQLIy9lmcLhsab6v
Ij2WIzLP6NRj5fvJECN78mMIGEXdAXi0sXurYhgCfqk4i9Z1nEumHkIi6O4xD5/g
DsPtue3gdpGKGQk20xgRAznLy0mtrpJm4cYhq+ypwT9uyp1OJwQkdM5hXe/P624a
oOJPyiWJc/PaLNDx5mEAnLfU4NFUFws1z1AmOFwCi1Ky7ezybZ6oVN7Jys8gWiAW
hgjf/6JIC2qmeeoE+qpF85gG7WfABr2ElY+rxyuKpF5DhEAUiJet+6RrGz9KZ29v
3KlFA8gadLt8KLE25XGFayG9cjl7AM67PKXTUxmASebA61Dbb18jfwJsyhSmMw0L
k5k6wxzfuUJ6rLSh0ViQMzq/rZvhp0+zyvPnmXkqHzM0vweU122NM/g/SUioHWGR
8WYk7uJbsm3C5i8XEJZ06ijwtQl80vfMo5mKnM8QKg5ikGfB06MqwOyhx8WUIMRZ
qdFtQQZWH+iC/Rsjp/exB80fuZ1nyN2+noIaNSw8V9JKPrcQCQnvSIpWXIJmFH4a
ceLP2/En0snbG58ifUm3md7douBTEPtRh4icUDHxRVpndGmfgYwggAtZt2FdisVV
UtSdf5UkwXd+tAJMXnGC5/TUCjrU7XsGPHdjbocCtQWrvptHI67isfhjDJZuv+ru
weZBCFxjb9bDwzvlKNvN5eYfhjCcKwrDEmkzhG/pnWX3JEUWCCNwmHjtBkR6Nflg
uu+gqDz5sxN9aJZQ/Gch31eOJL2ntNU44NobLLgQP2jv6QvgKuAcfb5GKc8eFVYz
mANPQwnclAPSf6q9mSCuWUKVUAv3vPJgcwVRzQqqrfsZ+T//ppW6qv4CR14H62L5
aopk3n9k5JZwdGvbSmKFl6cabJX1T59RO/xFteWYwit4rdGgFqLNeLIbwlybWQS/
WOaiP0ZYDOT7CeyRGMtoJlWGW6VJMNjVUcyjG6L34+wTx75hbFpY7yQo4Ip0tpMn
XR8cUgnK0kRKVunsrY/W/tmlAQhtNn3415NsqmlgXAr91hh9xoygJwMZRil0UbDD
AoxReI9QYwE1OPWhPTmlzEkswo10SJfYejr4Vy0t+GdPSRr0paOjOM2uEDj2Kj1z
FYeWOOzPu1Z/4UanpVcRV2Sj4Xmj8KTNFEu3MAY2CR/f2pxnrnUnVhexPACg/q/L
iw+MKdR+cVAizIMw/zjzwvB0vVvSnquzVSPlGl/UjnKIjVEUYFNnWm1Jomp5P5H5
DG6hoUzu6PF46mBBogjmxyKxq8A28TpasGGeU7pniSy2HprRCNGxT6R+4kJvkUsq
KZN/ZFJx1kDZBSdftGwrELXwznNeUkQVWxBkP4YiUuhlqENGXvpVJEyVwCMAfQMv
GEI/jlrcztTuR9mY0rjpgsBt0kl+wTMn99c+E77doecNucev1trtFLiWs8IPdVmL
AAch8DG6CsV+stfyLgT4hwNuiO2HYCIKsK5fRSOs1wktIy+h9JW65EbWL/QmtGHp
69c4+KiN6iHJWLW1hpAaaP+G3665D6Np7Lh+Cd/yLELYIC8QeIc0iEBQvXUQ+OJT
HQZFJnALu6tXI3NT1B5PNkJnhPGPSVogi1t7sVqetvonRPvsguBzBEDLzWvJDQda
UmRq2ZmXY/zkznTV9VpA8MR9gu4pe1cYHPCjSMzew5u7UiQMvLhspuzCRqmqIDtL
F8FrbP7eubG1UZ3xe4vf1aheG2P51jzksM9ZXFwAiI8VfoCABMCojPltL4UzgZza
I1njK+8GtM7UnvB08PRU0LfbFYtz2sasiCN0Gpsd9fD9gKA44kq8hXn5BamPc4yC
VDX9DFhCQYV6+tXYbnk5C2Iu29Ci3Gq7N+bGcoocCTAn3PSXSA4NNGnIdY+RQ38m
GiUpSH7UMmc1YyQYjajfVeqZ0znaSFJOP/MNT6wfH1QV9cnVc3MF1naYhRaOSlyg
cQXybGct15Njf8FqVrJUp7aVV1kGHemlyxfWW+Ap9RtlXEjELJ5+U4Y4DRwJ6nWG
NYQ3J2zk4vpcL4rjPoxKexD1qM7D78wsJWTbYdC2kptgEeXQndK6qJbuUjlD04xU
S1RfjSHAf4RDH3bH1H6VtOAAGShsKmqeCjB0Il/PJ2Ue0hxt8X7NX6f0dSvl56Um
OqocNdzz+GiYwmw2bY9Cqr/ulgOdXCq/Dq14Omh+4l8J9f1lCwxU7AILJxgO8Ljl
YRhYMRbscaGPCc5RVdZf/5UQgxsP1dcFyPHTVQQMckjANIRG6txiQq13c5UN2hLe
CZGSRHAC7CES3c39rWWfuhykwbMPoMGFgpt+vdP+OD0kGia6T1gdDWh9AL4Ydt09
JnJot6WH+Jp/tgaFc7hdTBbCEX8zQgdaZh37aof1eObt+WXwg53oq0FIWX2bGt1U
Cqy2Gc+RxgDLOiBy3n4GKKVJcbH6z/PQivTCpAuXtL6pS6C+iEu5gf9P5CJnHPHA
6mYLqOEH50D6FssAr0UqrvwiXJOIh1tE4I4vcvSWAMzhhs6za5IwblYIypFDorbp
87laLVm2v3SGOERV8Is4c6IGEVVYSelOcsw6hggMVQNf0aZslfw9shmB+VnvgOOR
CNtP2n+9w/NFaW5eKlRdSOUJ3XTZGB+8MojCDAsOHcDEEMoc7c8nfAn9+Ay+ocTh
A7uh0X05OY2LVhYxFEsoyF9QcEW7zxA7wcm8wzoGjJARTLYka+7CgTKmxGPluIbJ
JeKHHskOfikdB09cPNl7ppsd+BdD6R71jqhehClynFtnkSBBg7I8Y/GUdhNaE4Uh
BwigEmkqSFno5nLv0n5Eb0jjvO226iNKhAOgjj+Uwz7IeoHcFd8xpqpBhEVowN2/
Z2trrvLxdPM+rQUpHJ37gJ/0jgHbX45PHJw/q4uBb0Eg4gVHpg8M+Dqoz3clQf9A
5n3OaZ+0XqPlyyWheK7RNz+fU5FmxdFai1/IazOXkQUBx0+dPyTvqMvdHn1h/Ngk
lCRCJGJPIHLoZNAiEtGRTlKB5DcVkSEzyVp1bB984Ky1wExrqeSOQuHrB9KQngBH
mBzf5685oUyFs3r4iy2QHI0A1WWs+mFSwA8BqbA4w5jEto6ewT0IJ2ex3InI+6gB
S160W+aQhDsA0xpiuzIgQoT14SvWSLiDYazImxEePBZMSUtEfc31ot7M43RS+w9J
aakpFs4nAx3cfgZpftWY/y6sBIcCfRNNybIlAKtDIR1lPRrnN27YZxitJ8pPB9UE
cEi4BhdtfaN/pVSAl8TeSv3KK4x0ixROpyNfRfFTKH7GoC6pfQvtzjDSQRQkyj+8
Lkr+vt6vB9WO8/NatC5a0RUDkl09dxGvCoeNcPTidtSpB6os38MAhUCl2FoEaldG
R4TpOVPGmiSmWYi5yscLce9M3KovEqY07Xtf6IQ2WebEukYuePZ8Mb9zx3Ec40gA
hL4mnZzW66c15w6cAzOlLcZUHRDnDeAapRwYGp7+UANQ+mGEwga4UaKlJICry/rS
Fc1oURJ4qkF9Xtyin3KmE02qZcREw+WZGEhkgNBeESfYW8igwTfbYje6fwz46d+n
NDhpSV4BftVVeIS0MPCNWvJbWcby5suNMA24Cfevcc+y1u7U7Ki672DwfvXt9TEx
Yz0CSXsJN/c3uOYPbQCBgGLZOxLEh5xbv2mGatwupzorlykBZnfOmaX90Io+7v6+
5gKyZr/ctuOcF0LceSsjha4/JX5ZOYr5p1oFs9EUvoG5BmJqFrZTXqr09qUNGZCz
1hbQuoXpzkC3x4r38ZCO39RsCelnNsMr97/QB/76s28KfNOk7d6bv/MnOrPIV/Vr
Q9czsBoOZqvxw1Oa+e65BnyQw+aH8Zb15CG1GrkxKXMhJfRnVa/z0fzclhSEoEgd
iwrdAkm6sjAOattaJdGrHMKt1frtoF76jEUKNaklWuPeCQ0fErL+qXVuxAdNOCzw
zEVWtVObGX5YGZHR+eyGr38I/IJQrVefU4g8Nvj6piEVcH8OxGOkaauVfE1JeyWb
6CQLzzNdV3YiXIW3vpQeC7FLBcsfGwRORgPyZHH+BRs5T/7IBmJMBXGfgBzNmkKi
uWFXdEF/ZFiSyH4KLClXErUEWc5PDzC+8GEcV0Vwn79dsYu0tpn365vVEDRfigAQ
Onb58+29BTmDmnLbOgmbt3pDdyIMPqaxfPhhM8lg1hVJwBiTaVtjGB4mIH/lYAa9
pCU6Q4oakguOz6Wr15LdFKzzVr0Ad7QBsIJK0UbKmOMSytgauMkXX7ooyxmS90jV
yBG88wwJyLFEPiQLq//4VoVGe1zw2Eg3EeGUr9B4IxmW93F/HmchJnAFGrcipTC2
xhLxKoIaxMUpdrQR66wh1C/p0evhEiFOl+NKIwr0a5/JutwYt6cmOKycXugELyiP
rqyoAMGOsZpoby+AUdzFsgWKnR8tv49Y2YXvutXea/r6poN+oIG5jPKf8qZGbHIb
sz4eqOfwWDNQUsePy9QBod3cajkURFv1YSJ6lo71lgLqjaSSm2VN8GQJaqfs9/i4
8UY0ztU8QmYDOM3SLznsmp1c4XWMeToDgNKf92LY0qBvNxmb1nZQGrH7WUFdA9v+
EmFxV27M3tTE7wKllxfLSFILqjXEj+0SEKY4zjr5gYgy6zn9lqX7+UdtVnbPRfPx
p2Uggh6ICQGFkRhfYPCNDZ0gug+HmSIF6Eux1SZYSfp8Hi55WFYHlJtGKtMGXKz9
Uj1U4mfSX4abB6htCEk2RC4nUgkws9+BX6XFvSM/ilpZLn3tIN4BJgwqppFMgEmf
zr9DxmK8LSWsrJkmmwtiY64MdI8fS8TV7ZxRz6BhbiGGsMri6PuY7Q1OfXdVkXgu
+Mempkf81Wm/bF43yx7Q2A7l+UuG/zGrQmMANMOSxLOctZSSFRB3p4kSbdz+q4ib
5Xm7TJp/cGqBVBlfs0Y8DBPjQDGwonT8qqVyiix9ppuqyzQZXOgyUT3k3I0ShLaj
8rob5ZLt1kObaqzWrYJjaknXzB5ACOZc906pMdsnTxUAPKehVuFnCueCcIaGfA1Y
X7RwrrisF9Ui/RHSSXv9rNgASdC45q6XvRCk2UnPcAN5vlOnRrBv563gIO5fs0FH
DWZ2lqk5m9EFAi07CuYT64FkAcHSCUJ+dthBOEECuVjeQ2Ra0YZdQkq/DwLPpoiP
WQHyTVZyLFXlOq8cZ6VLDhibx0tygjsp4BrlHjF8jg5parokvblvrwVB6kCbqayt
pvWSXKAynB02SJInbgFxTuQyXsNws7J7ks6iQNrs8gsy/nCwWf/kDV2vI0VYinNa
xOUZDXUqb9/u3tsoHysQed9WlKW8wC6N+dbVOWn55YwaOFUgTc/70vZvko+QrHUf
qF0Y6q6TOolyku3jbZVQ48Aas8/QAth+54f1YWm9fo8uS/aqYKC+XeaKOFJ6H6/b
+/3oZytYH+ls9vCccXM13qzvAOE4QiVZ9yTJiJXrjmuUqD1GnmxLND5drfFaKVvI
Aw78jnbAARtAgEvabaV+gov3v8mMqyTM5n7GzocF1io8zTmD9MNbDTX+U7lXS2Kj
T+WMBTeAJamZQDpNCpCSvmGyyQPLFmF12boWS1TioCEHr0jDzgUOKLO3jfMZ2IL0
aNNNvinqUcrxUtDeYjgqQc7aA9HwXE4Q4oVK6S4uYwT8cjt7Mu6Ya87KAUAjSJGj
6TWudD8dsWJyVl6k+hedXF6eKh9phyx12rkczil+hqvRxvy2DdR38Dr0Gcb4SxEC
UdjBS5v8mCNyhajIlObwX5zW/m/PKMQUEx5U3QeBBM4V7KIj9ikXstwm4vSrCXbl
TIGoPE+9zLcYxr3Jgtkp7NIVfDjX34Xwk1gipGBLE0chiV450+vf6ym9NVEJgoln
+5PYA/DVaHdrZUS/ql+UK1C52AW84NQ4znnQfepMLJIfNjAX3nPErsi72iBWrcc4
VskoTOeHRPtAoMIgbMlNu3qfjXSNxhiH8cl0S5HR2LbcNjABBVxwPyYtgEs4ubtV
1uZ4BjfEAKtFS0DcVlJS2+/SPx+Dpp47mQ789o7KZzomU3GerLxpSneKaMvwt3+l
0prKLkBsEulDf9cbjW2aFj4aKV32tc5hx0g1qqdJIBGAk+a3pdrMd+JpLZdAOR3x
oGPJ3nSa7/OuTlHQbf9ngViU3z3OT/7T+y0v6G6mVVZRkSNVRQIRIKKNPpmKJXhB
hsbkr3ME3gKSeyjA+Y/IVu3Ce3MJ4osJ88azym9g3ovnsNCzA7akIhjGmWPqunRR
1i9TlSJbGqpjud7QoPA3BgVil5Rx4ewptHe7ND8zTxFwKvIxHODfLC5Pt8JKAVJY
QL3fkLQW1RKdZWj0PDlZ82aKCmYuns3l/xwvyU/kUkKCd/sc8yZVVOjq3k1hGMRF
+qf4HZsb87ZCFDgEW3eEdwn75WkKW5znSWyLmpMwnigedFaRx9viJ9e+/Q+iV/ry
DK+cR1Nv8UpIU28jfi4JrFhZg3DxexRUtFJQi9uU83EbdQ32CrorozZtg0l8eSBI
aG8eVGECwATjB6D2ERFWsAt22pdbJzX92vSit0twg9RbudlCLeXDQ+hfJ8eDfFnD
Lan1QLSR65//oom9FE8zxlCRne9jIooUZsWR1RHkSycms98dljoOn/FjfjLPFxYB
z4RYhydy82uq2kRtLpQOYpS2vIeGu93dnmMU7bn7ZsKpICKvwTITNhVx+ish7vUd
7o4eeTuu4xA53i+w02qxW5VclrjZ+rQrs70+xQvlZNNov7HBnSdJhJuM3IVfsaSI
oOv3JZZDMREmWyuMaI0ExrjD+JCFfHoAnhk2y2phOE/ZfAD+PcGsVp1CicgQkbec
0VqXcqb1s7hNTKvOlvC7OzzYyLF2dMEG2RqoBLy2tbeBNImE4u14aFMVqfoHyzTZ
/NfoUjYaEc8jgMGpuuzKzdIZu1bxvOUnAlTGK34Hb4mXTjr3NZLed+KrmsrGvSrE
fSD7pp1OovcJEIJu6vFyeaSfHNtDdXCY2BwIfCeG2SOr00xIXx4ueAMkNFKiF4W0
euSBGE5LXfX6kSx76mZt1AI571XDZX/kcsnYY1TNOh6OKZ7xkFHegcUpgmy3tL0P
JJQ8rFlzINrM+IWy7lIA3psTB4/xTOc4LN6CRygJdl6m5r0DavB1RfMsRoDBvN8N
9J6ilcg5hPHBjgdeVa+zDpQz5TlYBeJTuj2JhF0Muo66wCaGkGwct3SsAeMLgyZT
Y/lnClKrEhOdQdDuQl7MnDLPqUgI0wZIh4uNNzf+HPgHEfzDnqXbxUJk6WIAjjjz
X9k8Uxm2EPQjqVGVL7R7ISiNYlmIMcM9by0YiRR7nmfH4NpfeTm9Bl0scvxsJ0IJ
of5I8ayXL5mpGPzItj7Wu2HhdSoJsTioz/rChcQYxlVReyzpQChgczV4r0xkuFc5
A7VE+aO1JassnO3afDNBr5DDNbwhwcyzHcUqYQ4Yti8zOyjcps74phVNeKGpn/Qe
R2InDuPulnTzcy4sa35IRFFj6gRS8UH0Xt2skBN/sXh3l8k7Xk7hDlAh4hReuOXP
3vLEImWxxZHdhmmJK3PbtmSfPgDr9tizakbm4DcUgrMFu8V1tlIrcH9FMKqcrcYD
622/yMdHAB8lCGs5SydjvKy+3WddQPdLZO75NSLTJotIhce3LDs53gMRWO/c7scd
pb4KfnBLzG7BhKlgYt7Sw/vZzn1zlZLiEu1Wu+Jf/qPgiY9g+DPJ5YxNfrxfPPSP
kli9krmO5c183lRPJ93OO1r0MmF0SB457LRZehws8Fqf/z4YnitMYw4MLWqTjs4t
cDibc9XhNshoAEnPnju7rfcu3GdoPVTdUbv5HRajiR0k8fIQiVsF93RXXRSdb7g4
NHhWNWjSi/sosEi2ZFioei8GM9Sco1AisT4fK5F7k2weFCv5eMPV4bMYg0xp6hdU
iwdnR5rm8TgPGOu9kISdfvCqYDBatMOD7kM6JbfyJoFlAio+NjKdPLDR04NmkAh8
dDToScQ2EIU7eE964zB3iY0cS9bSGmHNBL57BBoBBsJhjK42cufMsB69H0/SjGv6
DfQvW+a6WdWK5GSWN8CFdypKaqePzvB7d3FjWdNKw3iL4P1YfUdURFiQM+JINZ16
CXL6yWcpDmS/UQYFUdBo00cS7OHTlRhmF96UnG/wRUVTKfoSRRKFnxVz4xr38Uqs
6bw4/Okuo2pwXOC7zqNEZlUG6E+hIJp+TZ4qyJtIC19HKMLkPSI4fy+9slKc4VGp
Wd/sUz29scKF59aq9kAUc30HB75tMcawXMZspNxqXYWYyEWyhZ3nV5XWlE9qpM9P
nSooDwcpe53nXRzikLVHSBzDPpA7pxwW3dzdOzibmAWF+upI8/L5FJOa1BANeZeD
hctiI2XlMYSb8EC0VOnWD7iNs6hM/oA8DKMD1TRHUH7ppPO2p2IJVf8saUWcKtra
GMFnWGPFFCLYL1c3Izod3kqfVZmvMK93HX19IFH6fB2DDz3gmm6dFXwmBLknaNpB
NPKkI1oKhfP+W39yx5uMyMZ8fyvVBa/Wj3B5NIq9kXdQlgx34Zatho+jOziJxPG1
seuTI7WSOSiUT7wQEjSLBmNTXH2wBEMz+jy/RMnzA07MdRfPi/qkEPFeqm5YQSYs
ZsVl5Fb8xGh+yhAIcs9quqyWblrJMUD9bqX3mmUzgAr/lyNw1tSh/wIaQNcTfUOT
04iE5iI1zKzDSW2lSq7Llc/AFLQk7pmPRdJT0ogkg9EoJmsYjUUjmRo2bXlmBqzD
2WiRbLrTIeWPao9330gn2E5Na4GQIwMxdEsJHUwx0tXphGLSg9DSUufNGKt62E0S
NEoOUxNELaAo5MFyZj7JgNqm7U4ItDopxu/AQXOTxu0Z8PSE+aKKAat1o5rzsOrH
4i2Cvy5UKVxbWAM4uGlbo7myhAUp1QDhrkzVsi0hKUjC04jo5fgtO18vgTugtkhA
FvcPlwJwocpVQ4Lruh/71cvKi43bP4K+vFOJlkRSttbNP2cqTHiSILhdoLumlck2
873mHvszU+2dqMbXvTKh/7IlW84KLU2gUrGUV6TSH2ApD/+GPACz6o12Ty4GCLr5
Je2xabUd9b+Oqff0qHpNieOEYspkOpCh3iA4X6muXf/+fsAtIbErwSWoN2cVSvjT
FTWBWSTFMsQWSbNSSLcmtjaDMkqRS/28z8hyiWuUlmB67/9SmAWqziZh/8CauZgw
lqR1WgdnwY8fjHK+3sxfvYOtWC+nBOtFGj5KI/qFlefynYOMSHgxcJsbUdia5C7j
ao5BJX2MGiGsTqblmmqvt1vQ4QRBqTacttvFiK8muLpRk4mUI89jbwPtyySh5emA
qJdkX3LjrLnhMglZ+d2tVXZ0IrImk87HX7uxT+J3WLR77G/J0bMD7lUyrlEcCZUO
iNxio4w0alRoftHxH2a6JDHzcOodVfRBSUV8HZ5V1S5xPA4u4GjOe1VoEYlE4u4p
hxjAt/9cN11bxRFH2C53NQcReSfaBkgp3uf3Kvtum4xDoAllIg+zVwQlgvSYOnca
f5X8qArFoGzM9L99SHuK6EVXWmdVMojo/7lKmbxECNrhKPtJsBU2bg1XwA60SrLb
/VsqNejn6wgCCWNxzBjKB/pcuyCp+qRnD+7dq5dPZdG/LuLyCR0BBDY4pMe7GcUx
VUipZYHXBvukHFNF8Mm5C5a4bsFaOkgOLD7IRkLARvJMMICSwj/vAvZFilcA1xqL
iAH/gCRnpO9hbrjcivTHE6knTgX8wi3BGXFO0gMn8Lsg8Ea8yfPa2TDVGQyrz+ED
UcHFdz47ECzmB2Ta6m069S3zBFK2UeicnztOtyZ+P+/YzOcDcCQC5k2l3TxHKUM/
xZSp5faaL+xnYNhKqvhktlX70jPFwCNFNpX11N2UlAt+2spdIDC0ZzcvmC1TueGd
xFI5kWGzz2wo5tlKU0Fn6NxEnJxR8gpK7ifTl1ZoSu74vpH2dDJej/TmrVuu/Lzk
+rQOGaRQFedKgDpNcYqn9ycW7T5ZcMohJLFteRCrC2fJaLs2TryvK7FZa5LMDIlh
udO16Dn7oYjFzDQvx6TYQH5eAbMeJGmnzoXBpik0waRp9aENLwngI7ndMBriqOgn
8CigJuYlCol2eAyEwO9hoWdYr2Z8EsscvMuJy74msVc65kaX0zfS/EPlPpnyPuhd
Zx1xSwQbWsm6Cq3UmzAcnBylOFYhYvhMniG8Pxuvrqrk6g6q2vk7NEwPR1RlIDaE
eivuu9ncEaCafRpFPfzwHYbICAVh3irc/FZ0v5jjRTLEk66zKpNPWju4eZHOwGrA
qoI4J28zDgnxEJvTd6ayBphL5JO8ouWuZFkUWWSeMuUddsdSkt51C5p7/bLzOBRi
p3xwDxjM+qlXL9j/6hH2YJt7aFOLAaSV1dZdj67iURn4V8HrnmC636oI+phwwx+C
9TfGD3AhczZ2YzOEf8e3aI/0mBZFdvq8txeKpHZqzH0sjqWknEVGqrkngfGjMhFq
QTH2q0DzDcJUcR3UWcwJAVsN50ENKbgMkmqfWt3zUApY0Fh33jqhhR93/u5LT2/r
3qmGfN07nmOpsYfPGNxxQRY2Be7TUW4AlWLTQv8IT6WCMxCdNpnsXLAI3utSM0Ki
CMtwcN6TSLaceM/8Fdt+gaIF1R6NsHJdj+LZnlK3T3xKsomvQF+RVybN47fuF0fx
vXebNehnx50G4fMSK/RwSwhL2DMrab8c1e43umIiMt4C8STBGQAxam4mihkvKdk/
jMG3s7lVLiBSRZJn8zCMrpje3i1EXqkRXlfG9RtTRxGf4HhAGQeu+6OBVcEpxLFd
5S/KDatl/VJufA1kvhMvjZ3ANV3FJSPb8r7A7fNPWqnwYGsmn9oVVnoQwvi72sXW
XQv4M8cte3d93d5Lxtwl9f8zIgUCRmsjROechdSHf/EpsxmAbM5DDBfMrO/MzXLE
vQpDDmMYS5BygGQ/yOL2yr4khJTr/j58jNPsb8uTsPTPj+L4n1xf6IUNEK02CQbW
6ddcfk/Grugr55VHr5D5WnGrV5ZleuQV5aetAcXXueS/PTpoOokF3NQe1p13fTqY
OCCZsaooU/2gkNRcAvWQjWMDAdkvPBeGAWUeRM2WiAzv+0Ka4yHVC/EYTmbmpTHT
VECYm9gUbkVvEOfhAwkSuy/AK56XMkBHCC7DMlRKezmtLreDrR0hLrdnj5WOzOtq
M7AdqJOMmjlQEqSfInxm+ZWMSz7+BxOW9t9LtIgaYTpZ+zFge1fPebXDKtIalf8z
ESFyxrhk67jzK/jD7jnveWusY/+DhZiSU2nKV9qOFcLVcJmh3L/nCzad9DDfd9+K
udcOQauUXF+NS0Np+lDTPY0NKUQZqyT0cvkX8INTcOsgMs29E1FQ0yCkk1ODx7cJ
vTD5PaI2uYgDztAeZu53PVGYLveZ+QwXAaDnbxPatB6qEc/nT7EDEyceQLJ/Ridt
xKgR11Bt7QVYefgfZqhsp/HMP5YGAtv1kxbNeN9TSonoE4HXNRvU/jEsROMp7y+w
K2I2lTItrrQ2oYXmPgcjXROGiiuDEBEZshAq06yDbEV4y+PwyQ0GiFiCMNNBclRw
Qce+JmebmCxPEyRzJ+548pCJv2TTACc3NFmspY70NIUM26bOXUh484F+setq9SIo
uHp7OyscZnQtpZaaw4yrTB772IHYsUru8Jq/D+R552+wflvpMwGPJdT+FDudpEXE
hfyx/Dg+ueE8gtC9iU1vmNihgxYClDq59htCxm3yLUEniXOkBbhsjHy/9bowF0jN
3TXE8S7merbymveCreDeqrKkbUmYJjbhUZT7PgcCNYusPHnUxdjbXT2ZGH4zQiee
FV1VJEyDZkpmjhZrMM3VIWEHGvvazIm8Mkq6I7u6+CX43frrXvhg/iXX/DLrhK0h
2eMbmKzHQIBig8skhX6FXJaSqfqFOJcnOt+0S1FkpW3AeXx7QxoYu5WN3S08NbAP
N3+Ka/lyeU+eEaiZ+stdKqw2IE+RP2gTVAHG+mMZ0/HanzycjiQpb3LYiDKCQVtY
9AdiDjdizWzVlVQW9goFIjP/3XsIi0X6SsNyDXLxfmZqrg5zlxTQ8lVJKZ105WtS
eFL9UT6/tJ2lqCTsJYezpDyBeizfTA4ZOMwTmDZ6z+gf+cv2rCKqXWEqbowBkbK0
fgLEmJzlDSFIslatbqHKfyV/xG6paH4sdmpQQEVxGijNUPLpcLIRy1q+7/KGQBkg
jZvG+O8XWK/yD6upbyn/Tt6Oozp4mCEGKxUAc3/iFVNJzHeYWEpe7Sr/ilON349l
26Pivv5Lq10x1hL4yG3AgunIcXsbLuYvnpmnVunpyLRXoqrHoO4kth+PGaK40+3U
TYvoCkLNXHMkUYLoR/D4ha76j1kPydfRaChSTQ7W2v/kQeH4774IvGorxxtwAbNH
EhJFNdmhY0mrEhaEqY5LFaEs89orIqvxU+Fye1QeSI1XfJbXgxKJhe4DWlHBlgHM
2RSkeB2ODI6juwhfCP2oFsyRIG2E5l4PRndnvhMzf1zraSS0rPyM8MkOoJYbKqxp
J66xxtDEsi0zN6uqCg9dmeM8piuG1HTQ87TZMAgcV8uK6oDtzmsQHEr56lPnHgYZ
4f8oB9V+coD1NKcc1n4YnoZMSbebrf49MRYGwMJrdKjWzqqqkmrpqTYqD6bfhHI+
/LpwBHeHAI95NEvSl3aLmgooaNafOImJnU1soepLF0iGZ6IjH0SvFJVH8mFFeniU
WYWM6Mf3Zx7tFdE543g/8xsDZjfm5x5jfa/R/6XYlmnc/TnCyO5iO47pz0FNKeSm
`protect END_PROTECTED
