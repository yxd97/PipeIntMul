`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZdSRyuzVUlnh61/dfoAuIzO8760snrA4oPN2c+nGU4bJ2j6FTwjsTVXTzklsMnX
E+WozsNzpSxFHLXAxHQiNY4NqPZPapTzsESNCFbzzWNYB+gDdQey4h79yQsO6NDE
Jjj9cs4mqM8eh7ZbLCoVuWTw2uY2hgFOaHWfL7VtYA3RLf98RgU4lF+Z7jbiQehd
75zjObglzwUCtMLzxO2DEckix5XSKNoriNLdRelwrEG7W/DLhOA0KVHtniJRfC3v
vpItVysTGxG2J9uEgktevbse4lKVmdizEgg1FJnUBpNXIXCKj9BB6VvW/Qf0xjjI
oiZ2tntxgEN7KM50sXFGJL7UYZaHYdB3mxaDDLjYC8Wqt/yjmOmdOVnOxqsxhGyg
39AYL/GglzSPYKL1Q1303M4lGoLrd9u5/2DCzBd6XfL8P1GFy/0I4HWUo4WQ6Qfy
hP22CIysZm+jksAw3jX1foHJMpi235V1XIXcdf/SneZYU2UViaxBGMZCA0hmfqUi
VSmWex97GPlaneYeCwcMdhK+LFEj9qHvpz/P3F4W9vGkUBIVKQx8CBYhDeHhmUYi
8pr4WDkwvYWcPRSIXvGIz9vNM13L4IfpsXxHP1llC9jkWYegaPi2X/S//5Qornz8
J4pXnao2yjP9bo8PNe0qaPjtWc0KnWj4NoU0yy3KQND9gliSx99SCY4qaMNlX2MW
faIqMAPjiPPA8PagT0OxYBwNzQCj773BhNvLp9kapC8=
`protect END_PROTECTED
