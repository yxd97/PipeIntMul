`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Wb9QTwuaEEcUOR7y2SRcFc7oKn0tRngPV6POU+6RY75AMfEllVwc07PD2gXJO25
ADCeGeTElBeqpx7RkFYxnfLNEEnK9bduE4I8wHDKPQ79395Dz7nD1UxIotdRmqAt
pkengZ+ki//cz17JAnTnUz3j6qbk0sS1u/8xACWRBMKVvvDkauQ6NU0G8DuboJa2
dMgETriTZUDDkulQxB+dXdXtEpmd7x2HuVfdcDwVQKAPJhJinoRgfaAL73S/jrWV
Jf8nOf63Qw6mTCFrlbAPG5I7n9i0+hEuQ+njRb0z454i5SjnUG278QHjhwyNpyOZ
`protect END_PROTECTED
