`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oJu9m0xx7x7nZzv1UhMQ1gbsveF8KChnPP1+OuXXYBQBsLe9D+05WpEvhV0Sw0ct
A2wwlDQsUsH031RTCyqasWwdlgTxcTHMKkzu9eIB79miPtxzYeU9Lo8GjdB5c5MJ
7I/UPwpFLgKbW4HJMYsqEz4J9bFz+fUTg1vAaFzCwTZIBE0O36qQPBSUcpAZXjEf
78xp9CyrLTZbV13cX3tDlu0/1kMnybA+upWa0u+1LLDdd5+NFfVB3ST+7u2KCEex
o1uOyA7HBxWOcATGrx7+McnQ6Nmph8+GEg5QKN9EXWHh3H2E1JA4CBbLzvUh2R4X
r8NW8guodpelu2DjEei7epp3p0aCqML3eDSGLyAnlqqsHbR/9pw/xs9uGjcEgo/c
NovKZ1LkedlGimtG1KlHOA==
`protect END_PROTECTED
