`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbSOEXq3H/2b5BQ1bUDKnd4j8+ektcvBfAG955kJl7N84ntBjSseACRZtgsq9iOJ
Rgbaj9vh2tLoVUDTSXw3/bx93v4NFPSNlZNVzr1uS4c1Lh9OMY20YXhBe7pei8Tp
agotVcQK+vOUGcSvQFLMeOAF45J6KWMLfkUodOkwu08F11uegy63qeSSsoVlVf5q
c0ThqFAb2r8j6C8pvrpm0IdREGoISezaPcTcIm0O4Y0c/TywMDZyokpQAvF+S7LH
7cPOdupQ9tnFTxjMU98I9UwAQQ7Wb0wNpr2Yg+7gVKV9IiWoxy9HaP596xFAFGLX
VkWlg2+VZpglMC2uIaHGk+/Rh3mYQ44oyfk0H27b1+sXtuRFlGUYCLHaeVSqDGcz
P75EExKpbGvoPdxdS+XI8EtKmDS+QqTcLVmWfo+sHTQ=
`protect END_PROTECTED
