`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGTq/Wh00dKF+NepS9lpmxIRPDQwX5oB3XmiTFvhr7jno4cbxF2aBxMExiaGB4EG
iPTi5Mx710JbSLINxUGQZpdFSmlIY2w+GsTX8UPnA2Cbb6W3xeMm+q3OUPhdsH4e
9okFPXvkt5lIRP6AmNs+GV+RC06JvakP44ouwCgmGYDtpXWjwxIglhU1U3rY6Oki
hQJhuWcKGqSpiuZd5fZBB7QZnA7DSxAFEQkvCgt8bi3/ysn9oNrha/2BGEdE8mIL
g87XYrhOeOdszBcROr7mPWJ1COIPy1NzG9YJiU9DTcQbqlWXx+b47E8ANIzIGzPd
yvFx2QKqJQoFLbHqq/1mhm+FAL3csNs4OXNz6c2Cpld1YR4our3H/YfeiWZcZPQF
UZfgbT52uiS3QZTVxSUzuqeuKX20D4oY+ZPVCH0NekF21YMwPfjFOE6Z/mAWYIO2
AK9K6FUOMouOKitnw4lugPPOUosaMRcQeTAwGY04HvcTBhhJ8kCbtjOd264wRlWv
qniXDWdaBDTK73KDSci5iaJ7hUwibrFTwH1NK+wm653PDdZBx29oTDi6RjxsSj4H
4RDWjFQs+VI184M2Ti1RPpVfUbhCevbBXb+dVLtOn3k=
`protect END_PROTECTED
