`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mx9uNJDRCdcJqpZ3UBu/YBdw6qOu4qkWNoi/jiYAPsLhIwheXAseO124P79eDML1
4/TgAUiyF/pIx6vTAznLKTxLnyfwY2WbbL3gnqUAbUAOIJ4WTwliXYEYul2TV/ny
C2dSXSS7GBkYWgDzBaNxyw0R5d3M9N0Oszbe9H7mMywyyPy2Aarnz1Kghj34w/H6
Yuzoq7loLY3Wt9HXHKBq5cWpTdIub+i7dYJoeeyaVKeVzUXzquoEQsmGsR8b/w/9
mNVF8UZYGBhFP/P0fCb2uqKFQz5/+kgXcDQ1FR6akLvCiAPeHbNKReVOOKfcmHLG
3+HGCGEuAcAaqG5sfsJQtUC71l8p9g9QjSgzEycwR9Jxs/G8l65DkjT0ZP3A8uwr
nS0S47XbsYz1BHZpCNzXK3YLqzOuQWna9psYYJoUhyo=
`protect END_PROTECTED
