`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qpGp2BSBvOjCcbkIxkJN7RUWHNRbPJhdF0bZ2ugdZ3fzIWDxm2rQPc+oPoGuUEou
AAFJEu1qvIpDAtl3d5qJQZQFCjtzna7qYDKLDGCTY8/nUf/mkakEcmOThLkmxWmk
hA0Vo5A9h2Xwlx6LfAgiy/4Qdio4eemkqribpzaacKN0UtZSci/VNxw1txZTeBcN
CmK+s/YtR24xy49ezBRVl+xdvnLL+yt55MLh7uXVizqB1kUJ9nhHElcThnERQCtX
v0t5v9AwgiAB07tqpf1b5sQPzQJe7r9yC7yyzQw/uGqvoiWySxYnUnNXy8gQtL+X
k2l0ho4Pni8MeahCvqQ6Sn/n+F3ADAsyQHsfsfgl27Kdn+cTdQbioH0imAS5kdW9
WyqUhfvr0tI6C+xAxBnMvU59eaZs4rQsPyDDAjVBLtNYf6J+mFcuBdTSRVIAYeUz
ThzkqAxrUKaoExgcI7z3O5KXxkLZltRkgR+J4Wbqm7Y=
`protect END_PROTECTED
