`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DWuKis88Zhw4NgLxGFsQU0Mh5g8g/FiMM9wNBsC5eydrpfE23y/qdnFjVQKDHcak
jkDqU9/8N4wVBVHSsA7QSovrIUMvBLdnuqyT+FtU2nWJHX/Xp2WjTPjcspRxtUsg
obaso7jYAYvQtH1ImTpLsNl7U3VtTM8Tpjh63eTVVxYDyQ4NCjnm0ZbJaNALrlgh
AJqaqqBUAQRF6LTnPpFn+TqFBJRd+ckX2W4PZzvhskao9JscVO4nEd+kCSqHttF7
njEhQcTWVkVWkO4o3oy83DfnjrMgSwN44HN4pHS4JXAEmuxPZEwraFSUiNhr4Qc/
u62sjpteaAWA57uYld2wdqHgCKm36uOOWg+y9UF03Y7yVIkqbHOVTaMhULbC56Pv
8CQL2QKJKMeFWVRcrVByd0g+9xUGqDcUO8Jw+MXuh9CHQaci9WfbMMc+ZPCaevbs
bAtMY2yrJ5erTMHJ0gCYYD2iKUmFNEWzB/NQ7ILo97HCvy0CYIT12Jt7MRePm1o/
ufZQVC69BiOw26mkx4Flj4LpI5uXfPLts7MqYgHIT3JT6kb7sF5wJi5x35xqOvvM
Dve7qoNZQcDLHEARKcnWqxpX4DqLDbsvlI5kV6+4/B+hl4MgOwPwksqUTc0K4ZLR
u1JYl+SKWJJ4PK3lq254bitUlfke0CE/0Wn91NeCcedIo3Luu5lbg/UWkR04gnT5
c5KmlaGb28z7kYJ885UoX2Ua5PN0gwkGRQ8HB1Abww6JEFQYZSISwDp1cPhhYvdQ
rJmBBHR/0mRRnksvD7BgCU27k/d1pmTruwUxTnmjYE6WVkyhm3xO6YrVRYa8noLY
3wOKUDWqFmeg98L28Xc8Cj1NT/Vr7rWRPxE/pgEmZYGw1uwiTpaykN9xdwHK3t4e
m9ux8fjwEGM/kHbmYTv4EeH9/bTqe67Pq7LYX7AIPVdK6U6oI2tDlSnQV1bGoK2f
n3PJvwk1d12nFKXF1rko5+6nQwXwpxLyO4iZfOFVStxFoE1tJ/+jbhC/86DyypKK
P2aKfpVM7Qf0f86vwX9V/KSQdzwvPbZhFd9xIxikvwda7Ili3sWqc7c+NpMLOA1S
dsdCO4TkLt+4ojBfZeQ7nnRT7guZMefoaJMlVPhYhA15xmljWVZplmjspmdEajey
HjTSfV/v8l5PItQuktyL4HYKla0Gtf4mZiT/xqoibXcnmH/SO5gOHQSIk4c4p64s
OMhP9QPZ1R2JFGVKTX9//UIfkkl3f94foSZyZhijhuDqkl8a1hqDIXK9p20J3QpU
`protect END_PROTECTED
