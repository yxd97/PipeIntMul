`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwakBioFWABFHJC1asoUxM3rhcc6b7wjkbxHz7+tdey2db3TJzj/0h7uMDitq8un
1Jm8Okwwo+vkPyhlQ6Ynd9ptUdtCRG0MF6sBv7n3um8WkNWjZ/0cPNUa2owCMhwV
HIXYmnknxJKD7fCwAbQtQm09jgaYhPHpW7/xTyZsNuBkxW9xzeag6xX8B2dc1r+q
KzoIAAn0wKEJphBu71UY6tgkfXE1kSTSaaUCPUfcBMjVgUFKqsErCqJnVehqULMC
h6uQJCHyoYyj1a8guDXWtM/BgxkwNBa9YdJ18WdaeHg=
`protect END_PROTECTED
