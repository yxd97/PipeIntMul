`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GDpXCvx7UV3QXFKqDMnGQARTaF7P4uIWwKaxMn9+4QNlxz481sDzHT3Kw55ixcL3
r8AHRffc1FRNFPYM5ubbe1af0UQQ+o5z2POoNpCaHw1aueK3JWJDgg11mdemMN54
eMPvnWwLOEz4GK4xrkdmrF73m8aVVxRYoWueSOmHdVDKH1ZwYj/dhN10WVltmYv+
SPGoddopugc0jCyRtqnc8hIAcynWe2uygvcYmbdVqqghmr+Szs760G3sltNWXtyQ
Z8AURHNk9UWtxPNSRS7XOcZCll1mMUlLE4CO3mOrGDMGgw68fk0ZgLrP4NjChLfa
GYwiZ9ZhGwdhYgXZIQsiS11UNRjHZE3t7FoqBvKftjG1VNS8ye9sO8sCUX4BtxzK
Zyl465oSYUsFL+Z4MRWRt1HoO9m0ofDL1SbakoxUQS7vjxrQ+77vqGbmGZN5UFdD
AoimH8VzxUpH7n79DtV9Qe9bxlKnrTRN5N6vIqelgCFCY6SVV3K+GeI95be45Kr0
FzxGSQFzBzAxqI3PbcDXcV0gCTBtEFfQsncolBWGgv7cPM61n5s37ak++q2T/WJR
2UGBbbd6TAO90Im6cTzWaYVSYoZeARr/jBx/jT4n4i1dlQYH2VBlPj5+JARRMFvs
FK4czgKvB+DXuKUG2fZsd1EkNXZyayCru83z8rtGy5C4Yu/FGK58nAfAuqLqjM4L
tlcdrCq+8LjZ8Fi98sf+Q/RsyRTaGR1WPEzebhy+JSQqlzyK3EFxlwyGTA+4VjsK
hsn0ekwdkZAZbeOSY1Urw/yQY3oHGxpqEvmhpEYiO5XJV9StAJpUoBc6P0YZX29a
SOJlQGe+Rwou7RIy0grzLaGDwCJ1m+Oq1GZyIuctinNW1m2Lx4jmLRBAd88tovoA
g+2qrpdFZTjaYnygmFWUTEHXzxZnq+xq229vZaAfvjaxkP2QQ1Gn5grNQhC8J4ms
ce7r125EVLCM5yD+6qXKGSWl3u+zNdJbN7vq9F/O1f4d3lfndyJ46gaMDul53Kfq
frUqYzN20+bqkJCNHDPt1Hj2YqIZK/bKDUcnkZbM70X2DTjGlbC5AJYcwxLNeDCI
9MyIbqg13Imyc1g0E9/ZPf160CcgRa407JsLt8RGaWJws6rnErEz6VMiHo6epUkC
Wv0HHmwqiSlbG0p1ICqCtmoyY/G+rDkx9FrSIAccZKTX1mGZtpx3Ll08ugUiB8Kj
+JrKdlTTba1y4YR5Ij5XPB0R5AbFzZqGlT8N8paYnF66wWfPirOThGhFcszMSsgQ
Epumzo500iFUZjloF8eIVhVhTKNtfQYztArBRgqM2epqvuqNQsLa8Ws9bA2ijqW9
Cfz4No/J+2ZEAkYG/FZA/YAsOiQ9fcxEm3nR6WwShlPJDhbIjtbpS4+C80bG9R65
ppJfdMcffcTY8sPCeVhzjJmpyr44IV+pW3Ao8FQbvd7aq+wNrRc5qW20yf8M9deO
USB+7aGqirJp1mpJN06dgz0zX5sfyY2RsIjCdr8gh1c3BUYcJ65OGMhMvEsfPtCT
Nl1TMj5Lb3zrl12yEPzwZ3mVj05X51LqCeKABwefE27v7nuOsCmDJEaPcLgoIjqb
BC6oLwKbd/fRkwH5bWPmdkmqGZyPHCypCM+TZnSCbAsg9oPbfVqLgyiRPyw6GwT8
6swnhv4k19zgQM8IFWUl1uM/vFLeeSUDDOdI61B2H8+CPqFOfNJfttcBM8MatS73
5xrHr15A1Co0HKR1T9/BJNJ6CHO03EkUh/N+1yauDOiOmzxVOZOuIobj9rK8mOX3
HXOI/cxudHZxP27A9g20eqES86LlGjAZOg8GfY7mXSnGQl8Em5pxTGOts/FbLCSC
gKRagKaPogalSaNTFVTAZibr5wwirp9kne02HH6dvCO1QsWKQI2pxeAMrMUcN31c
yOvNS0gsSSAjudnnrfTWTUU91pxs9DDANgPEe/aS8FW2ma3fVlgkBd8PHRHt+xzM
NpjASkVsUT1Q4fv7HBXT//HRQ/JA8jIU2F5TjS6Yq/Ra3u8GSW3xdeHF6XNxpVPJ
9FRK+7nFyqlI7IztkMv6zwPyFEXvvIAClQOvR2Aap72Y+0s9X2BgU6W8JNCMA/Jp
lCE/a2rlOY7PcWsHwjMewz43rvO0tWW9niB09kl865M=
`protect END_PROTECTED
