`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dow9tm1gwK7oZAwxOIFky6EMntNkLvLoG1HzZJNEkqhLQwqu0VlrDnVHFsM1wC0M
81tPgxz59YbQDI2+J3x8LxlQ9/g/3quYb/EoGL/ZZyEGSWw1soxLkCQh4fCZPtVF
e/nixROaX7AGMcAiG1BHHKK71YmRxNEE7kujh+nqiH2Gl6beUM4XdfZ2sXv1xFcp
XNrdGHuvVCx+gUTbx97SVwUKW/+c0w+PdL5hMzMC/S0lGvoQWz9nlwVVQ9Pbkka2
i7ZGPFlUp+/ceqFlxUSGIKpody/ZhJe8aPkIbZ8PJl2ZR9zkoZbudikD8ypyqDo6
t9adYZ9IpYbm2LYYPFulcaRiqybag+ku+RhMjqz9xtif3Az+0uClqcgcvV1TYY9W
OJsKqd2J2J+5UaDnVRLsKz5iJdv4Hi7crEhatZ/myVSmrvEl4zv4UB+WZujSyPLn
1+TiWauGDDwYTH9pVcRyFePCPubdzv1HyrAL1/6VY+mfb2MqgdW7oLOvVAdFu+BG
CkES7um4YoDZgIuAAKeUZINm2Q/Cd5+MV07jxr06WnN7DBFw/iEFXnkgqnTTSuGE
bQbWJ3+ZmyKMzzr9m77JalqoCRC1KGUO7fDbPqdfVv8iQV+IsV35Lw16no3nsYcs
DVU+Mmt0pqDR5FyPPVUeb2UAUvFJL1TZTC3xBAAjbrQkaXVlv1KCgxQl5vj1dzkd
Uo7kDwYTKZP0SD06PxmnqEN2hUWqPrC9YCxdLTZSq/Z7MbEonISynxPIeGKVOCAn
Sh/sceI9Zlvf5hsNb6F2ugIzHweIMWHqDga+C+sLhuToWrYYhKL24jK8eVm03r2I
eoDvX/0MXeBRFjwP8YMPPA6caHorckuatTqnLM6Qp3c1g0inUhNEwMcjGKAWkzv6
I7fsTHxsQD1dOADl0J6cGbGYyl57p9/DlLzPC0jvcaDvNY1kJHcE4WSmOBhgYJd9
UYpO0l8wSTJIT5OFcU9ijjaQApQYousPf4e8wB5MM2GnLWfX3BKgFAReGo0TtHvD
fZ25tnsfStAGChvJcpRtu3MjRsxrgA+WW/IjXvLcQ/Kqpcze3V9l2/FnjVmLWOWz
k5tMm0u7hWU/wqlogYZhwGI0V2CgNS6Iv3qz6fFRCCwV3dMEVQ3U4h27UqRDEGwM
YzsyUx153joVoJkryDO4tzv8kFT9xsirQ0DwZK6fONd6D6d9zZV6xYGBAelGLSko
FzE1y2s4MfoVBZfTlWaMRBprMPXEhKdQHeBi5Rck326kzSRWyGD7GOoiTBs/wIE6
P4tfzwn0kLIdQYNb2eyngsoYkMXWHHo5UaLppS5Si9nS308WuQYo0KaDiJ++W1z9
hdFti3Lh+5bdqUPIcqOwHa8dFKST9jOcVm1tqkBTJJZOdsFffo6C570TwjtD8NLB
sdS+8jbCxQs+HFoXAyaXAIZ1buNRnHVjVRLtzBWBDGYmvmiFHXLbkg88E9mg2ukB
IoBBIg0clpT7R0mr9Br2MpbEDipwfwGh+NaabQD1LYbzxuh+22IJ/bA+2l7u8B98
HXfnUAHWo1u3n5BqV8a/fgivrkHLhXkXfQWaYjYtAG4BlRLsnDQb4Dw4r2R8kudB
P3/B8xA5gr8klbUZEfMa4vRKOJsNGZ4FMLGandL4gMaHgC0SxFISQCzKoLZWX+cX
x363hjKiAVzJbQgvlE5vgagd0zcwJEVg2eoGHDDHIpRzA5+zDb361+J0QIBiPHNc
w8/AXrTMb//t6elMVT2kcIqXGNpM77gvhF5cykp4bZtUlFg+PRbkndnFs/PsVfuN
9Flb6LxAdIUN8yYONIuTC+cHPV1GcI7HqODaQ0YYZ0p0TXlh2KndQSDPrpC+ncjq
U+JHPzG+f2pDggBdzAnLcbk6UUUnhaEOJNYTo/p5P7G21bSFoUAlD5jnN1uR1aPn
NLZ7UN/hlqRE0QF4aCPYEKTSg37+Jpq3vY1PTwmzxcyRnQpXIpucPdAKTkWB0jvO
KkkoESaQdvUxK5AZgupMS67jlDXjTn3aj4aXtsaLFYvY39D1b+9EaWT+Nik+FlXF
A6ofmXcRUzxlYbfkEXbmkmns/xw/OlNupUfogl7Pr9ygo9XUToKS62C8lg/cjJcS
ib+qBoO7+DNu+dTcZvL6bCapNOczYqWA3AnjdTtTHJWZRoj5+zIjhdZeXo8OGHaF
TwA8BOTFmrt8Osiw/GEVFFPF8rzDjLjL+qThpEby+lMnR7lMi8z2kwEns2BhuIRC
t8YiTlgsoCXiKKTu7YWt/2alL4oBFIlEMXVuwtuFim14yE8tK17hpwwOod5cgDxW
qH8oAA5VBraY2mBam5pWMx9BuHCUI8eIKfiXXoIfMBC3XZnAmCDvpGC7yZhgi+2c
mX5sNGhmDZ0aBAigiDM/rpYsQTzu3ldhRX253sRQlyU3glB4UjokMVG6hYGU14Cu
lkVTjK9k/I4CkDINd2bTmDmbmGYpYI02MDR/5uUL8LDFYr73mf0dpS5HLsLErEaL
48r0c5kfYDVGv2Nxz7CX26SEo2ZQ9P1FUeQerJmZx2ra7V1GjjWnN+a8Opc80V2q
TVKaVkfiSTtepuS+Qv5p8Zs3e0l8jFAqYmB90+c21phtMV0yhWLsIYDg/auJqa7M
I1otU7IQCWH1xniEtJwSU3fhKG/HwAVeodkPpwZruk7LkM+6t/YXD5+434fORQok
Sa0CMt2oZdqE5LAimS09zQOJoxQs4He3JZeW+CQhsmD/3OnEo5kz7HynqPUj5NHc
Rd/Am91iYlG5UaPheHLTIdePppDNMG/uu4OFPncNM0BCe92C7WiJS1cuAabRmnQN
v1yP40Tb2lNaqLPm3DePma1wG80lUEcNDgl6tWwBve7osHfZEfE1RDywEKPpLSbK
w7HiGyDSq4TBmbGPIipepq5lrfTCWJinKpXXAuaNkhJtf2HfgQf2vFtfbkkTT+Nf
BGH63vkAtnjgAlepEjJwcAKsn0h+/Z623NEhnUEeD4PoZSKUg+0aB/RJM5p0te1v
8IS0uoGXUnBfxWkv5YT/aTHn4ieiZur69e41KWCSzO/GvvB0/KRwS5xfzY2fZtYI
a6/mRM4BiwdZCDcv91pZa3cpikxF5k2jriMioEDIKoNRvPRNP+Kb9JqwUuOYqb/u
dxJE4hX9M0KhPAM9anNaUDlGCf8nfnqf5k5A9sFME4d6i39JUHTk81g5p64eiTqE
BFZD0HVWhL40Ndve33rb81k/ukFnfZw/C4oCPYyTrZGP2JAFnIvx6wCfTzaE2H5x
4OZCC4yr683g/n7LB1lAvsRGmbw591HkZnMWfPS7LMp2oZnL5RALnH10XFlBRknm
tfKN8gDRDp3dtALQjab0wpGbjyydZO7ew+j6s9tYuWbfzrVs7/StUpoxr6N8OSDW
AEfQOPoqQnnD6cdtNo3UJesSmUf0vjQLMgKohvZuF20umSGVAFOqDH8fwN5x3/rY
yLgbTteEzV1cWFAy4d6wc3Gyh8WmySVjtQSOzx2uNVpfbYJWuduXxAxSt9aGHpbx
GsWenrXOLepSdTrAt1EbCJhz243JhCceJZXR3y9W1iy0bodHx7nX1/eJlgStpUwb
Iu7MmNmEHC0YMb+jXXLcKWen6OyOPE8xUvU+ll8y+mh7Pg9FKVII0OLyTYFtjnbE
dOsV9qOY6kjy39EYeXNDc98lZHMnZzSNuoxBqDBg1vk3/9OBYKb8/3IGY1gh96lt
eIr46lURfH05e0aIfnDfDBIYEYARxSV+rnOWa3gYudHnnRJ3Ynw8YJ9MCj7h/+Br
3ERrQd9PSp+fs0YLZNf3L5J4/EU7gc0Nf8GvONpMfnzyGHfpui5vQTsZ5y6PsPBp
+utf5SoZarlUG0RcWOMO0Dur/WaB6jMKynkUq8lesbJlQxebpqi+Qi6aQ8UtMYQ+
fQ0L/eDOO2q7BiJh/4FayWFQnZGiVjowiDd3GyjS3PaYgydR1ZVcj2xYkqNd2me9
IhX9DnJdGKKSBMg3h4sSSP4e/CYODi+BXrCcyiibMuUibvaCdg7Hj9/TxfVIYJ9k
Ig3jdfMvBHrBc0SSONZRzJH5BtTZZPbHE55QZUnsvq2iI58HRpV2bJXr5jbY1mbg
23q8Ey/A4YoT9B88AJP7IdlDn9Alix0GwEVzXSCm5YaIU4dnAbBILm8YchRcDg+8
QZgwPmi5l1vZN6w2AgejrU641gcpO4SmgD3DGbVwbpfqGKDm2xwT5aU8OAthXRdI
YXbit4sddd7sqqz8U7UJlbyO+KdwU/Gl2Gu4SqVPxrnwqjNl/C84O9GLReGUxQd0
3wAxEoE3eyViJJb8+4PC69G7Xr2Z5dtv8gH4axUnDM8N46aEla0PBuMzIiBXmZ1/
qJarZtmCQEwfHXrVgnwUkLWDkFOISVrsNRqeby7JB4Bv55ID1SnbJHlXv8SZcMtS
3kZ7PxeHWCFA2UUgMAyV7paAnXl4SmsQYaJThVb8uk68G1B/BpMl70cjV4+dJcN1
oWo06v5D+5HkwV5XiNi4/Awg56xp7BvWH6vJJrjo8utGuErnf0UUUMpHcDhA1WZT
cG5zXTzxhZtl9FurD/2+uUapeiV4VvVWRYaJL7Gtsh8Cb+Q3TdpYCexCE5O4kvAe
jEM7fsZxbqFgsDODOGtMuHtfX3rUxddRmp2kJxZts+fKm97CzUsZ3plsp5cg8Np4
SJIYKnG5Bjxxtr9BG3qUbSfqK684OLx52sNyzy2nbeGCzSrSiUkekRCuhBkZoJVk
PKHKSgeLbUeQhUUAi+YeKklNF96nxGyoFHsNGKqzjTtjkyOTqSNDz35tRw8jEr6X
87XqsAEwA4TJQALvr7/MAyG7NIkC6pZhjj2twspxYET9f+ORazKR9Bl/gGcvD14j
ffuDINXpP2B495LKGwTVkZeQrGcZfpkSi9ozQP4yUm6F1SdK9F2EN8SjefJvwWri
Tte1LNa1OpAK6+NqovvQpC27nRGhGpwKsOXDcxZLLFnoDLTIJemahGvZg/Ir3sbR
IJiWDP+nN6zn7Rr5gkFLEvhDQG7QMeSkQr9euknhgAgyfk2YSzGXE5cBq5WGdtvK
b7MIPSoxN4s1B8M69+2M2ZBZhDaRMq9Yvr2M8ZZ4rDRZwUX0SkeAJuRX00WBHXKm
/ZoBjH8VzBKyaZ5NPqft04q+yXJtw8tdeNiW+sHd0IwbDSbDKepFc/pOGcmG2y+c
2zoN9YRE0b4CEw8ZWF/MdkVkbzBuYVR0KnyNBpBYrJ72z2aJ5ZzbyCWcyevh06hD
TrynpHaH8UH2oFMJcupNyK+Hf3wL9WONDgaoEExyvbcZgCgIUbzFbKmVzoLbsbrN
vwn7EdV32cYBwa5vVuQplWvGRmn9ohLlw9GdJO5m0jq9QnGxMYraDflTA+L9LOY5
m92DglovqWc0wMkCxIgYRhyzu9544v51UL9+89hrKC9tRuZqgTSA3IxiG9oGDdBO
yAM4q0nQUiz29l0MC6shZtCPHy/5CVn+5UkbTvkGLiaV0fpn0jG7wW3e6RGEDFzD
H9YLV7Q683fYFd0ujaNINXP2WKOJ2liLyU6PHFOF/y6HvNlAXbdZgQc6SkXQ3IZx
C4Mi3PmiWgL92edpuoRI945vbfHGH5/cd9Y7b50fnAniz7gJulN0gatn4ZNPzVsS
Zsv6w3/zPneIhxaT3FHenQdna6NN2glmL7Kdos7wwpKbehtUNq0r3fWb2ZfF6QQw
F7eBNNhGtpADsoI12OY9u39Y+8lBOngRnuumPLVoQXCS5JSTuFM5fUl6cueKibR9
X+HC6LhxvjD5ogshcahO4Idg+srBTTrwkZhsflkwNKIKZ0KUY15QHUwqUe6t4bB4
f5q+5rwsDYCbbrfXYeWvitDwUOt0bWf4g+YH2lEFJ4CVGJFkKOvbfAcz0mO9Lf81
rGsHx9GEmBFMWZ9vbuG8LWhCfdIQKuEs9CeckT8hx4qq9VvlEoqGbLPqvtHKTrU4
9FAPX5U2yhapBwB/TVkI0FWeX77gQ+KBfLA6nsCLYOYmNRXccclF9C6YzhCBAnKr
vo44jLN4T2uSs+DvWQ50RH+JaH3fj1WCx0JkYaUCJsMXzPNLSCFldjF8HFPYEZWj
7GCxLRhP1T4outJ6kqg+qsbHnZagYgwUrCoCP9MZQYh4RrF6q8jvtzpVmeBTiiX0
sRiHrGaFHXEKLH6F87mXnOJ0qLAjblBYojVp7RSl/EMzs9oee6mtveu/sUDNImEh
eUMIL51W0tlhpTnowDuYZ3I4TGI13NmzyG49C9hZkjbXqJ7VwkhP6NLxHqa2Qxfs
NIedVxd5zB5kqOSBiA/MwO2Lxvq/hPk+TePUlCXKxrEa44YzWbbQ2lI3kpfu9Nnp
GdmI7VwM7t/pAw8bTvLxTRdoNa1mvF7ZJzHiVc/CrH/KdpQVDDpL85em1ivmmYnJ
D5D0F3U19Tn1cZKrQoWtyKJmmsFOFXHXeIZuMRWEUiQ+x0jwkqRYHaV3ribtDSfB
MV/cUFvkv+uel4JHx5VXCjJp9tHkl0BmpIuLBuDYGkLgywNoKr4l1Da6IxtPG8I0
S1xxTKlGcVjrGyglEEvSsZCUruSfLCOBLokGiIV/7eml2njQsAdxn4BUznW9jCDu
EvyNGDxyyQZwAq0JUitm3TQhxBVeXCMAToqWyX2xzbo7ne9Nq3riYCCIkieq8wKf
fXyfj0VTNlkc026uT3srioo60EBcRpklXPGvEW4ZeS+EhH9WjTxMyz4NpdP1kzM2
3mCKPl6vZW9enAazdC9Wuy850mClJLMLf38hwaZVwF7PA8pfio7duFpHqnMM7jcE
4OaxuTemSyFEljaxVbetO0CCMBJDVL28qzfkn92b52QlY31ZvT60u8SAGqGxvwgQ
xaaPE6DF+dHvO0YVVxXBcRUSg7SgHfUdsbp/0qLipFAJ2id+mn+t5UsX1OClaR8u
Y/P246hPaF0ZWVfHmOpg5iwOsRkVocu8SQraYua3E5UuCQ/NJ+HLO6QZbFBkUdza
nopgD+3xVptggsE2kSZyDa7S2xHywiz5dCoVQd9+sHaCzn1MZUiSIMlD4PFvokms
WtfLt4BKu5d2fXmhPXlSBOcUeheA5/Fwr1jfRY+A4X55TuBT0WWfEd/yod8NBo7z
pSOGy11mzz465aKLRnmrk5I1OOVUPAQi+sfQMLPvxdC+b9WNJA2I6OATyAqlUPjx
CDSvppmlKAfem0ThBMe/hxJnM1MyoCmVzQyEwxDO/cN09q0sLhzL2WU04dXj8K7/
1W3k7nfiRxGbxnL199V+3DqS82nAIrse4W4tNCBR7dKZJzEEPG+V3UrvmuT4KLcx
Ut+NpbTBWgGCV7vLgTMfw4HzCyTZ2L953/sVVX1GU2UxoyJDqRbaEI/1jA+Xc1YF
HYDKd62aaKKli6SK/fd61Ru4YDFCODIGifmlZR2qO8/g4kmZXKTMdrfcYo744w2u
cuT/5MtokgpI7yt1TtVmJ3ak8kX6bJ+aMbh5wx6mATPNySW8yA/eQh2By/k6Qoxz
echVAfioFY+SKXpd91PTEi5V7tA0aINgi8x3c0Dz+1FDmpDBCzUfANbW1ui1uFAL
gMMPJD3j/ghYpBrImCWacUkFukYEVGqminps3EmrfnLnMiqUK6CvUkM494nE2J1o
uLysnnQDI+5HfN9KX+6M8kF/1yg8ucKQDxl8Q+A7R+KJdh2URxfbRoW/A2qonZ0K
SjB37TV6N5vJPlCjHx3YulSyyQS9KBkjF9EwdjEmn/8kOHGXx6JjbGlkmSTq+Uco
Ha/lTRD1Ycov3RJ36ZHYLvGj7bFXnJkhf2Ie7BrpYSOHJb1qzFoQnW+kDM8MWkd3
UzmU66FHXrZg/mudD5zVRxU8gYO4/c0BPtUCOH3U+d1T1uU9ZVAKC8CkLotHiMtb
M1xx0ePmbW7sVFBSn1E40xTfTwzKBl0wljfUdE6y13gAiX8kAmNgWpKh2tx7p2o+
TwDArfHf0vvwEfA1S3d7aoCDbMKNXdR5kEwZP3KL1Kt5nh7FQUj0D8ApYCKSCaIy
3W/Tf7Igs6cQpzUjSFsyM64raTNLsleHu4EsdEY8nQuoTbDkrdJ4fSNOLYLwzOOa
yEWeXQW4f7OblzF6y+J223/4mdukSVFl2mzadu5P3RU5Q30DiPRKC+CxzK6nM9sE
iyaTbIziAc/xSQrW25ENpfpLbuM2Se2oSo7/6BXTZ9U0IF/gVmaGgwihO/u24xrQ
HHavb8lgqPol87noTXm9y+XFi/kcmddcs+869ElwkfVHBTfMPJfhKp+wlNWY9ZWE
0SOJWnLSSzjs+sf5Cvott7C0SmPjJIDMeWXO+MHnfUSkI6ncTkaUMfDmsR9N4BWh
0NralZ3uDorgHqRh0kcr8RBiJZtQvfJwjUcdGkir5ozH1HQe5WSscPGeMHFsBYfh
U0syC/TICzus1ZMP4WDfiIy6IjIQboGu5ZfQVfweij/GcGQHyWxvoD+OdiNr4UC9
Y92/8RQdLO4E+eguDsKl6J+qgyHPBLY3AEJK3isKZJcbaCQT3zwxTHOoku+4cOqg
KrarEkc5HJ3qRnTvSCzDIngpy+4G+zZb/iBSsRp/UDsVpJYOxDLWvwcXAuIT/JAA
c0VUmoyZSgLCeD+6N8Pyy/t5nKFU4p5X5+qG5x2kOcNDshgvhp2YWjPniM94LwTB
/aziU84oovlMxLqcLYhu/DS+2c+p3ltM2IPq1ro9gmg1OJB2/dtsPZ0shJUJjoz1
Pf9Hm4NKoxKm5rxISd6wT3jr1KddWuc74Ey2G9WNn1kcMHEnA9/7NmOmdIJbZVpJ
R1LmBUnydDXEev6zACdaoN73hdBB2hEnD/wPuGisI2yyWuQdkZBWcrfttS/PLs84
ypzufDWSDjWDWbpWAf/XgIiAzkXcryja9MaQCigt4e+RnMhb34z0Odo2Kkaxlp5w
VSsZ/cKh2HZ7f7tS4+2oHPduBwipjKeW7syObqERIw67zGwPiN9DS3m16bx+t2Rw
ah4J6MOVdcsmRMCrAZXY3xuGaH/++bEtATiZyLsRrRDTFdDm6m6oivADfxLZ0nr2
vXgqP6KNOMFXZRyGCe2XrLZdsgvMM1Dzq/n5mM/OREmVf//y4HIzGKpgdpPmgqFr
b+4AudeH6vi37PqDIoLCaOOl/fgtF6ibF9RfsKmYmfb8WQWjYurewLLm13far4o3
LhiQQIkZw/DCBqSS0Q9Mi5CXj2gh7ujPn3kmABUTOcyXIrzkqRFloPWnCYJkHjot
bz78tupjTu+1nlp118ZHoc62v/uHBGOAOUIoEIi9ARyuq1GuJ8110TDj4Trb01G7
elWFWEZwl9BRnloHf3Z+xYSwyvzlLciYl0SAKgAliNSAJCJYkKBkrkf5GUNFCiwN
gzYWaGNRJWqKvCPZZgmzvbL4Li6N0rxndTaSKeYv6wu20Ts8j34OrlTqbLB82nCX
36ARbEgeiOVrPEDei/5qcK+DzXUDTaX7gWfaxwriV4kPuDvMZMUcO3D65VOABMe7
+CNYaXALHKoRfa4UcZpg+QS7SastePJUlLCnp0WhGoGSSpePRyRA1n65k8yyK64b
uiaP+KOA6Soabkq+L8hSrQRfYn/dGSsp9z6JS9U3KHcN6GIjgoY2DZSEf2Gs29bR
76iGCbO1fZSw9hUhXaLRwcpwDB8j27InxMup4qVQdqAsXOAE8SEixTr7hY80bTbO
crqs5nNpMcN6KopDA42F53ru64/xzw184CKSztWhamTb8zuZWYPJjfOuI1IZeoWf
zEcWetlm+Rge69HywZrS18B0gTtvZfMUdMyqVZP/VCY+KD6Fy9ckvTYL4v7hRSOm
mHM2j54I2Qvj3GHEmCY7P/8Volb0E5zg5fIENeHgL0t07EBG55rePzFnnghNH8y6
EyYDHKjZLdrQj7akx0lngLJC47UDqo927/4Jq1UBo/ZdQLymsbb58Ab4P2gO8GV6
IMveclnXQAuLFHFFrvuaZGf0BCso3fUXTSFyJYZmBq4/NPnKhoZ1cofnv0MfdQ1I
AS/VKOk221ttLbMMrqxR4EjRzJBj+9VTPh0nrxBKpo8eOY+uRu5auXApoO6IvsTi
Cp6/UR5GPEuOPK4osZlOjfKeX5tIV9vd1wvq8oESv0ur/br0oyMkMF64tKRfsPTB
J5tb0F3kzDOFAqNiTwrco85EdfWjT28dB9jzDr5LiicoWUX8fs8fp/Sjcx+bXK2m
+XPVfmaE+/7cDYDcmWVDiQ9RsiQiTEyeJRp1a40tSuDxrYAij4qGN7VRFlCzgrOG
NaApRnIdeCWt6WOZDm8UdtU3TBPvVMCplR/9cmzeTfVPetDfHvp6Vb7yos20XaMx
5trKYbEBxyGuuoHMG+pFldnLVAiF96578PeZGv7u3w2AjVRvSKjj/dVKExKRSjE5
hHCwSkfIxepQsptVkfuz3G09QS0oAwJ1GGH8aLFt6mffrvJCM8Ev9WKQix/SftX9
65kIMdX56dDoaP7GkQJe09/10Dg0yRVAxfIoIfe4XKEoXn7dto/jLv+QairROgNb
RLoBjBVX5rObeMNS4jfo6Gg9wMEYhMsThDWfxKKVdC39pkqWzxocau0BZ/K/i76k
agDCFH16hafBxWuF89PbT08SMkX93j2Ko8JtK0OF0t6MOoSTK9r4tLkHt5HwgcsI
Id1q9VAXV0HEAYuugpapmqB/g3EWlWiJDVjQU0e4tPiZM/PRf9LkS+KyQnFiuAEw
a2Heu8ruSAMCuXugQfWGeFkK8C9qTDihJxl4Z97tC87dWGKzr4MX/Bn7GSOg3BL2
8cszC9z7c+w6D2fmYbES9ns3Aw5pc40423P+EcNDZgzfZY+5tVHRu0/YsTZ/xjXy
LqtZ4tV7lmgu2d1c7+mLTxPo34WLH6Th4EBOlU+0f89Y7JROJ64wWBFHCgW7/vSM
s6w+dqrKCAF1WIMlRyNA+pRFAW6gp3cLWw9qr+2F0hcrnH61FixjzTTxHOKqgXkA
3pDlrTArpET2rFNoSpj+x8/E70EmIfvLlL+dm01J/0u7RetFOPnz1vdF98uI3tbF
9+Yc+r7cvIit+3oR5rZMliI1aeH7IiDiPUlJBDo3Wu6MZIEx123KQHirbZ6o1po9
VP3VHDiQO7StmVlcADDnYyQr9mCusZj/KOVbmKU9mDGfhTtaFYPx+6qGBFwl17pp
3kxJNOMJb/6viSu66Y1iChK0daRHKZ9cvHzKPxXd/IIEl8cZaEEst/md1Rqe+wmd
bafmRg2DOi4E46CR9uPBfVre0RmDUps1npkc8n8OomWc3+ogJFTZp1/uCTWqBRXG
I0NX7EXata9qjG8p+VrCYvm3qV817dQo8mLjmv8jEaW6YeDln2HFRjNCZklpGoIv
3PFWepvd8XCyUNlQrK+UilkZr2vqcwV9d6LcSSqjdJ41KzKwGBTRsBVgXe5OFDhg
BlBVxDt13oknlsQ228B2/0opLT5r+IldS7lYkepLEsexo56mNc/wmy7JRvtf1UGy
cIzXQard9bt2gIOJGgpTgw0C3Y0phVVvC9a2VDwOjFchGXvroaCrH6LqJYih3BNU
qM+LdxdmBLIdcDJxR0d3eq7pLJ5TdBbjltw+k+XOL36R+JYEj84z+1hGsvMN7iAr
pmG4qjXMLGVBqdbMH8Vp5eupPZZl6AgfbMciUM6IpGL5tFCWrmdVEHPtj08p0rGR
H9Mw6G75p0LmVRK7bGT5NQHNn+hXjuCYdsmRDRpJw/xFr0o77gARlvVO2ezZs4lV
54dedNqDyKN9yzFiHp5m9eb2xidpt7u7tSdzP1dVNgXvFJaXdnKqXs/07BC8Go98
5l51YAo8lUgW76/Lzcf2+w/z0moo8+lelaOedTPerjFYYG5ep5lO/yTNzLUk/QGK
jepeOiyU8xKLco732bnIhh7MAQYuletBSkshiPZSmzgBV6dFnFiIpTP8vSwn397J
gQugRphXHgccnP7EmosmSCJAWfjmRmL+WzOvj6dwvt4AQW9mjryv/0ZAhZ+wtWf6
dcyYC0NdIQgVD1WwVt5OsWdEul/SRHIAZrnMCZA/PGzpWf8GexwJ5+Pydrdos5JN
LlOHZYW+1+MBi0ZZ2I778wDo5hMh2tkO9yh+ULY8/fajP9YDAb3wOnefyMz1c410
pOCCpA90EDCpvQT3MBTx7TJxvz8vtNthAjMPKM547Rpk9GWr0HV5NyR/ye9LZOIq
+ZQJ0APIqMJXGwTpcWh8W6JYXFvCtzd2c8XS+RkOPolGH8VN9W73tzYQV5wSYhW7
24Rq3MlSmMBlzXdIbMKI/c2VRzCz3WrSbllsnNwkTZOiyrcGBeKq1guNGJ+t9xeg
vZRk/gqVWjIZnHQEVEtqmgndMbNwdlC/tNyYsXDBaUMyRY3GyEC+3bRVAK3pX6U7
BF+8eIgRIx7YIkOujbJzhg8UBY8bRpeg3xO3S93hK+WKAviDF3y1Smjsw/qBAF7m
sJwLHzZ5u52uxJU8/mvHgzTDN4a5cl6FnAkDMqYZ6uKydEx/3wmd/JPporIyZHX5
BKLN555PFZkCC2R4kO1RLiVaMm/wm+dG3QR1b5GM6zKI4qDlIOHqlzsyM5cIwjWh
uwvxGiAkR8HN/a+e9WCAyRNA6hCNyxA2/It7z1X514HDaLlqj/bIGmWAlFXWWbRM
RMYMZeq6Nk8bwooU/bReZl2EjeGJt3WB5IWSw2WWGrpAEvQNtsSos+nq8aS6KbIa
2ctq6teyQkpLrNLrafuKXSNVRaMNtGdlLP6HUR7UlTgayUil/yfIJupyKwd1pcSa
8EpgSFS53+oSUP8YCl8zvLCg0GI2U3b99F9DUV4Gp2kLmnk6Z4mR3VajRG4h934F
pGhuKFnv8gvmpZxPG0mzAPxwzlJ9l8Eyh3WeSzHUmQFg7T37OMeDblpYqgddT7tH
HFGBlyKuZ4Hwr4reB1R+hFSkx1wg7xvBnHJitLCBwIGNkXe7wdqCOfoC6JOadBWq
ygwnydNOfP78uwDIK99g+HTjU+YgfMNOaJ9RfSx2ZySGCt/XS6JFibaQVNFPdQ7M
J3bD2mf3sHs2jELHJhxmCCFzeuLc1VGWAlpXWT129xvCixCOl2WC2vTtp2JJSByj
5AIZ1JjlPZun2yPJZ80WY26OxPxLOrgvFoo582uqqTSclV2Q5jgW1WOKWq4NE2uq
/8un5HWFkjK7QfCZ/0VnsU1Nmy+C1QsOf5eMRVp0NTbmJjhmqUwlu2d4ZwSMuzTm
s+8cfvpL2GnpM2leFdU250whmuc4RX+YCHf4LmkKEbKg31Xplk/1qALTl0LVnGE/
fQZwgxw+h0ylEuZ3QD0Xha16PfDcH/lkZxxjMBIoCf/n06aYTSdwIu31qXPCLRz7
Clanu5y5qjsDeRtyDe2GCRYQMrMy9XzMHTAxNk3HGbqZYAROmvFGOYim3QbpCQQk
rG6Wh7KcIrD9ydQfuRoBDpHd12/YbJitCxAs0fPR8zsmNtmu0twNUroLrVukSZJi
pdxc8kE7xQNKOUwmcC8UoFyjT8NDpQt/yJGkYEN1L8lpwnyJsAWQY0ftBxt9Bach
pSxDvuOTpc7uiNmCNxFQCt4dtCg9iv866ohL13+QMv2ycXYqvBfq3Vkn9blCi+6M
aHgdsVvjXs5x3sY+AesIJKDXRBK1d+LuY+djgBt2+5aT1CWRBDq3JNGYamqQri1X
LGNqN4K8/OGFcIy6BzZ+lAGilAaWZoya99spcCFsHmo7RZsSlEr7g/99VJv8+n/Z
XeBnXjDZjCYuKWs87I0b6Svjm5iSy+x3mY9NxOn5BuE0FqfhxGaLfog27N/JGRJx
wcfCNKifVwP6VFuQ4NcntRMxwyxYiK6eloqCnZHx22kLwUjjAB5Yb1IqfjIgaFvG
e5vQfmij2GKMEPID9TFbiXKBw1wO5uAevbslgV60arvoCcHq25F3HvTAmT4R7spZ
hf8e8GEiGTW2egYAZvNWcUE0dujaXZ56oypvYFfOWH9L9M3tpk53oZar0gu9t01y
VdPCDE5w7mPOiqkvBVYa3X+/hdj5sZXPW+8H8RICjYqR4Ti46V7tZqv5MSKZSJh/
4zKdvY+Am6kTBRmZa6/o2VymyHromqNyGc/jICVuAM9S4W0hphcqHHSuan8jx6S5
xgfZZLsCq8Xlp/rFMC2BedD34+YWTq3eAe3jtW0DbrNcwkBTH/3RW2wmfWolcoXW
b4Sdtl8c4+QgZMF/fLfKyG5+eszESNuPdVPv5ryEXlL2wht+2bOFFejmx0kUftWF
UU2LH/dUfG8f1aUmyiHcellUREMsigo1jOmC112hPq9gy8G5U6NG/2O3ZTL9Errm
EeRGavMeRWT3rolDAEOKTGxM3J9qLJ/Wh7ZTr5ahCAdNt89a9rBWBY5hfZJfcnPj
ZxZbE0nlw3p6fuBIITCDaId8NiNPCr3AQSuZ5KhAqE7DSXRoYmjIu8pSyK24NoRl
vF+LObE8jWGyNmmPfNuRiXJjf0HOCxCGHe5yxoAmKwnOHtpBOBVDd4IvV5wGUiaM
KaUemVCxJ9GJalNJ4m2mIVyUfGKn9NNAGfAOZ8lSqeJsOuIKPE4dBjU/W7Qj3Vtc
iH34Yb/ucY9qNoi40VLcUm3r2LJ7V36RSyYtNfBx4ezPTBUddxzfxm1TvVcEYLkJ
enVLoln4A9Sd50TaHBgQCC6Qls37KTBJRHPsG4AXPexjhKgTfaziwrey5JBbAChK
y9Pw6ro8DfUZIKURICiZsC0CsuKrjhXkAGneLnjgJnHRGyWleWcgrboCdEw5bnD4
VmQDI8AYwNPHpYWzuNZ/N45NiF4S/2jHkBANi45qNu+XJta4/GMCNcfYcIYAPEUf
8buMRJuRFn8HvZ16Y2yEZrym5Ki5XZ7mFRAwDYCD+feOooJHEdX3zwtm5i3HOOno
wFUELRXhlxE2WOscrFv/9IhatxYCBp0mg1J6fire3dleppqOMKIKvLDDF3B2e2YK
8SUFYqizLB2IVXBUmUFAPG7KOxH8UUWTFp7nCOS21jaIDFa12yt6+EOaA0eyYGFG
HY41/3RfQmcW7ge3rbzNoMrLq6ET4GU+MaLZH1v+K/ZPjOh2zUigTFUEQ+bOkITA
zu8xOtbmD8MxhF/FBJpXxteUwRS7YPKYw+SURa+o/sa/wtEMrsx4zJjkMvq5WtFN
RZ9j1g6FvsN01l3qIiP+rgSbOTTTbSMCWjLWqMv5XhiEPi9bJL3WD4uwcfEir4IM
K8WDrHxa0+lZngtnySlHsCzvpq6a9eMs9PCGG5Anl/w9nbPUndoZocQVGaImpyli
tFIICYMsoxqnb48h+uwiOwWyFaQmEq66hWQTnNV+z9oN0db4uFDO4gq0+64ApTgn
jboAX7uDnlmhXjSl7kNc1fY61HVpwa32SWm8rN+9L7EjB6T9+dUGGb5X0w3PDSCs
GAForu64UTsn12ucK1H90KWTGe+/8mgFP4q18ZnyJi+S+WczkVsJLMHr9z4D8UGp
v3W6D1gVD3SM89wQsrKJaRfbqf/o1Jbs3IPX77Kf3CXiM3HPMsQRxt0GF/1nbqje
N0d0E1eCY6zqvz0TcsNDBWgzGEts46AM76l12zR/6feqiRM9KKQWJtmx7v42zwJb
1k1ODPrjsi0yF3K+QtqhfVjS6rLUMrLmRm/vjEq8B39sx46AwkGVWCPzZe/aYu55
CD3SlBh+t83jmrWyUmBTmWSztcnMLD2B49X75WdnGmHSzM+Zkgy9sz5JKXYWBjrh
eogguFhVTMUAEH3VrmVPLZh6y4TTEtkfNnTRRrz6ueOoAwwDkUuh5dY7+JhU7G4G
4JD3BVvCN9QRtWQfbVhINuIjSRRtO7NrEfAVI35+sQg5cKwwMHbNxEOwV4u54lsM
I+fIp/wxL+6oFT8hK6LV3YArYNamiA3SevHBvCtv0n5nuKRJ1mmdoIGWz1FlvQtP
0TYAMGNzl9Sg9U5tCNvpDotkfjjUT3s0LZ4oIG5P9f6UdbZGMhCP4mpFypKvgpNj
cGrInww1txCNO3JOxFPKFy/mwKNtzbZnLxrDghNxLnLv8C+wk2zkmmTnMQxlcdHk
eMOfGgO9if6PqhNbVNEE6bHQlseVjaw2TgiWfs5+6Gchpb16XurBO+kV3GKcWBPe
34gS52kRXihRZ2LaZy+bdb7zoNsepQKDmLeDxdwqob5146wrYPWDFg3s8lu3SB8E
1MpAIPzDz4mkZuqG+XzOlB8m9uZSn7doJXx/5YtY1dkD87sSiaA1T8COXJl9oItU
9v+E2OvjpsY3Go5kwpf+10lUsWUkIZygjdVIYRcAjAY3MitzgBVv7CEYbJb9rUZE
VXukYk6QaCEf55cB7dRUn99wYpGv52vHAUG2WdzOoJix6zqaaby/DRKYQkEOVULC
69CTTjxGqJw8IHvvuHofZ/pxTsqAoHgmuicWvuqfHdlyk11uyNHPS7O1ezkCsiTo
c6vTeT7fZBIxoXmp/sA9mOVxdDALEuI0bILwKmmtXMwwA7DyrUUSSCjn6nsHsPPX
lPARpNMoQVqg+T3/Uh1stbdhXTZyNNfNAnhMkeJBOn/aEkw/b/R2wLxcHVVr22BG
kco+bXq7f11HSApFOTvGlwsXYLg3fAoKj1hOJ6RxCQCeFWEWnowaCCaHFP63n0jI
a9PTFx1gGp+KytOdMU8ZNOokOZZ/E5ZAHROvB7ePq+LowuZRuj+pNN6lSTrkGT6O
Aedt3bwlljis44sAyP4ypdBz+xFUG9vV3KnNVmloczvo3jzdCvvcKD7q4/C3LA8m
YyqxyNcldIeoKlMI4muRTUV3mKug7aKInq3uCcx5IJalaNiP5k+XubMFGRF5jc+i
1AOqD478NZ4oKB6cx3GvFrgxRHFW2SSdIUKmITgxpp9yOLcEDBV5qrUgJKtKSWeV
NkxHSvs7VkEN6heRZ++a0Nrm7AvbxLU5rxqzyWnINb5vVFh9DtftSb3gYN0WSe3g
Z4WF/mc+EgEyPaHdEzrlcMHkvH7296tjUJP9eA+Jfrbaq4dFj0wAxWbLduigrzdI
GHRywYcHf8FKcya9lXnqZ792qt6bznMJIin6gchAojoovxGSw4x0A+pRoUi3vTo4
amDLOPN7yXUaevvhg1ZZoLF5zPgKVwIedL+Hlc7vs9fzR8mKpeVs8zavlTdDMC9e
gSsXXYzsa9R3/K6+71PTtMu4ocrJ6S1IMkTJoE9O9pDkmxuJRnfyFrykhwnm4M2E
m+fTrFtsM9QOh0jUFxx6nuqV9yPNHDFwpvzPGNjyvM0+JTudjUgSEVtE9iAsWdW0
icnSH9rgGRpf+Mu7FJneH+qPfSq7rHTzWnTVmvcVUriPvxuiLbXKsbmjHfdVmWgV
nAgiumQ2F3q4mGEYd3DhB1isvjtWzRsKpZPgmZ2KyK5TKFWtYjn0V9zVT0T0C0dT
SZQU3QB8IoYCQ3pCayOQuQQBphkkoNPmakkVb0EDGZNB70q6kO3etHU7wV4QYLhO
N896A4p7VCcDOzPOszILpuIL86cl6a5Izwj19yT1V1vz6uGf1NMkHGmYY5cLLA5d
612dY6qGwRHBzZaXk2ZvGiLHfHepAGlgwVoodGMHbElft+fD3NAnlUF1mr0ohQPl
PybeodAv0hgnMy/fVNbXMZ50kjqJY66bXD0vVozEqHyICAsbLRha35G7XZgvTY/g
EHCHnCgSyggc8Ty2ugjQtf+GUZAHmIoTeQxcR8hljnqhlX3wH9k9OVdHhWn7l+7F
B4wCwxnX++WjPZi71WJgAILAI6Zzrj7M1F5xWPpCFb8rV/EkL3jPabJURQu+2joo
EiuIk8x+HGlQ+9BklmBuFKJYSsM8iQwibQo4yHwEDLO3c6cfOaeiI5Ig0hDsa4l3
RZTFkYScC7+Yx93CICltHQ2QIaF9xjrriM0yxNyYS+BDX88uPZOg6kC3AMVOofdu
5IdpK18gZa0E/gIHM8RlUQEh3ZZ/UhFSth0tl/x8ivM/k9KQ68Il8eofFMkE+UaS
ftTnXgE3dtc8xsciqzvfBiOkSHo4WyJwu0ic1CpZeg1GeHMJPEMGmTgvJuwc3f5z
54Ou+iQ1ZfPTXdZRkxQ2vJDgZ4+6HfYjHprw0wQpqyggsYTDOw140mYy6GvKMgqb
`protect END_PROTECTED
