`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tU+mvSeMx/VRTOMVvfSOtbJsi0/Lj+g5FxNeC0feCWV2VC3ShPDa47ilMlRcSoyi
L8t6yg98NsNX8pzVGU2g9rT3GJCqhYUtok/88HRMQ2AGVZmAjNpjOcknt/IzGs59
jZeIGMl9b9Ex0tWTEjyy51jLm0ux7QnQr8zuFzVyebM8Sa+XwJZJki2AIzGcLW82
ITua0E3qA03hiyqwotJFLNAlFs/sI84180lUNvWnAtmxt7wRs8aFQMOS5vjlwvI7
S6Ui7ntlXotcmoRNzdgyPAOu1iIPEOkJAUVFbEKpsmHvijtvg+JgPqH/pL9p7MEo
wPydvOfU5Ivm8QKXB8uMhjC5hBNYYTL5vebl00U0v5kg9Dukgn9yUZggC4Skc6/S
+fpeATlu+/KL4jvmOzy3xAlHZ1ntfnQsVIegFmeXn5y57HhBAcWyXMRf6xMnMEOf
KFZhO6kZ7goSnko6UlwCGzIupPHytCAl86CbEIWYUIEFN3m6os6e/WkfnSN6xAty
3E9AFTLP/hiaJPalKDptBDaUOvaKkRSrV3r8JCz9SpcYRwDx2ibdFCvYu4bYjBXo
7YPBQTjdaFxNB/EDwy1eu5oN4DAAvVoycVAM/oa4hBkmpnHIjCBdNBA8xUXKtkNJ
HodaoTU1Y+kq6K9J9yP0W82t1N1mwqljgkvcCmWzTppF1BkBY4jXFk6graV/RxIy
oUW0l2CFh/y0hiSnlOr4waySSvLiIpkorIPlk1vNsOyAfR9hmLTQPtwy1wiNoLFq
+24rnsx878tt4pFQJs0rGAJlqV2GI0SFboIfxEzsm0Ec0MTlXXoNTk82I3uOLvGu
b/bbx64i2gtyYwc1UAH3rhpQHuhXKZuUjLHAQz0rYN/NxQBluQFg5QP+EewMhWn1
OLvdimKqZ9AsN74y/MOVCYeoHlXgdOyIH+cA/L65lPR+R6xU9yL2Gfj7Czox4Yp8
c1su2gW8ygcZ00dhGkjvAelNHxGbH7hr8tbWWS/AN9U=
`protect END_PROTECTED
