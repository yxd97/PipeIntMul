`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OkPSxIOmVBS1VeZvAKatJi2Y53VbNKErB7/4N9uvMAlKbl8FgzO4HRGvISgH3zao
XJwGXNNj9NAX2/cb9SWAAzILohwIlcH1Oob9TyNnxEeJ3a3DuLFJ9gqP9WY2/Lzl
B893Mtu2Jbn+8McImdvJnsB5e4LFZBDRcrVHraLHsKh3MJO1NiLSAPBh7pKFG0eL
pFY0odA5qV6so0G4TxonaNOlZTeDvCg4d5qoZxOC6SrAftJJcAVA94D1Pr1nSQDl
IycaZZfYQqyB3EbzXxviXn6CKLQOgB84yAMPpR5bSana++9yx8VcbabdelVwNN6y
YqgYsFlifH6EnLI0k7xX71JWXvKy0tM/Cz8fI2GUp1Y4PGKTIAIrIPWbla5TBaJY
KFOfb29qh4/5Bh3bHeVZpIPx+ls8dJPGJmsjCIFewG6binnQOaT9AmvaALub372k
p50XA71GissVY4R8wkymEbpYUAuloL2CnuYvD+5O7lmuJLT9JfpgrhOKUsQn+iJD
sXNvOH/q+rV0i2m2Ii/UjH3RTlM+81dr+tXXG7jBijLE2XbAtx1d1e3zeEP4SRW2
5l4pJR9Fv8/8j2/FeX5u3S3Ej/FYVPGpJsLerUn9eyqketl4MS6NpQkRvxC+w7sd
jQR2i723Ek/pmcD6nF1x+2mB7tBnvcx3i3LJMMlongYSjk6LfU0/LqE+e9zShWia
/iPckzZAuz1LkhBX17GTXvGx5FsttcrgT6mK9GbeUrO13+ytrKEm51hjrUs78tU8
0YvaLrJ/jaickSnDOtv79W3bbLh9D+N7u+oo0Vo+X7nDCa4qOwlbgPsI3X+NVX9L
MmjrTPYdtSPMNP8nwXKfYn0eT2fQpe3uNmiUVmWb2BAv49rBMUvSfr8pNq3zI5sg
kaShxUZlpRqUZhm3VPe/UbYf2ih0XuuqNn/P3YQ3cKWFzChk77NAZ2Hmtpp0qgwP
UnE8PEF8uNjpIh6U2UZLytgNF1k16TVVf8Xxqz7Y/1arIhTTwVbKnCFMitxYkBP/
DJEqyCdTzordDPJVtbymK1TmXZ4fbvmNHnpnn0RL2ljyqj0auu8EvsdYTShNiBEA
U5juNzr8gWd00xkCKkynElBNSQ7IMTVkXErG0RoFhcXFb9pLxB27FAvzkgXfgTaF
MvyYeOhnN4+FzJu7VGw3cgsQygr7Buo54kNQX2Ido5Jb2bFfBC2aI0DRcIEykVMo
0x/t9E9Gkf8NKoZdvm/rTATPb9RoqTwxbwm93L3j3CQDxw3zWRaE2ZXIMvyH3pdn
6bnaJ7/32F4O0xSwhr0wWg98CY5uIjC1ud3Wkoea9uI2Yg+lkgQdFxNe6DVU03+/
nr1CW5W5Ya3ODhbt9AfCnGI9dCw0AhQCVOEXc9vaaWUSu5xoPNke/qCJJc7aXrvd
M+1Azv8HKXIJ60gOL5zF+2TLNzF2a0ekrub+Vi2Xi5KPWRY5rVPJmNLqCubxEjP6
I03/YzjLNe1SjhpvZP4czZ3XHu/CNNV4MymIFsAilSp3Hl1068ZvaM8i9EUINZAl
9/by7nHJ9a2xGCffnec2HiZ34mQr1m8Qii9/cmG3wgiIMeuoleE6vtKEemWFpcpS
`protect END_PROTECTED
