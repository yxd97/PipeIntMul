`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZ+vKyCB4bCatwOq9p/Ls9iaUkiZf8V/oKqZGLCtt2zGPU10bLLxXUYctD7/T/ie
iqisRR17zVbEg47qKKzQaGHBmXLPHcKNDuJsTsPw2k31P+VlsmGvsPoghy2Sl/E0
lsKzLbU53VPtsHrpy110pdRL93egwPNykVhAA2KSD4ewJdTzgIsBeuRIc7QcwUig
3on0tnFKEJosiALyIrW2XqqSzJalKB2Hh2vAFJnFlVeZb3OutP9RYeJx5C1gbZ5d
Z/CwoJNlwOkMWzeShCnykp5dmjHk5VCUH1o1xX7wU3vwyxUCKNxxm/rxtMkjob2o
8B3W3RUWQk5SxwuyXhRLRDqxIE4bx7J8yez7D9iqE8xs4JkYHnI0EzwFK+4ULSfi
ElPfHJ9luO0BkhQFmjEuXg==
`protect END_PROTECTED
