`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHbnw2tgDaLk5yNCE2PIQw0p8LzWB+dqU0hgIgr7MJ9eS4TAd0QHDrLnkMg8UHqF
mDSwk3JfT6UuKFTVJmVmLMAirfhlubwBjKMyPxDO3tGdc0YOkheDWKrp96XrgWZS
AzLfmNo0z4nFkG8Tc2xyWyl+B4cVKRslscqPJ4MWwXEVCk8qzhdtBkMUmgbFwTJU
tL5DECLSOjwO2glSmPHbYKUnrDR+mZg3ZYSeOiTsxP30wi9xsKFUcBJ7dfeQDyNl
Be0a2rzcQKDX7OLo82xSwZUoOa2WD3Y2+8yN57Qpp6niGctVjR9AOHGrJPvgRCdQ
5L2AgfaC+6pb7U47RFXyQZOX855hi6I9OBfBoigUfouqjs9rLxtpS3aBjbkzrWVV
/9SPL6ncB0ZdqI4KRUQO7PumeIMZ3cIy01KjV9akvR5pWljqfmsj2oVfsmNwC3kE
kIO4tXbecUT0gv0rFDNwvm0M7PtOOvqWvq46DgRt0A716i83+2Mo3KAWsph0/fpK
ScbtpjUs58GrL590UDjUALHIiZ9h4WYvWZOSsMFkEljPxSelncUohIM7/eoe5eg8
NU5ZVJ0hGx7xYxM9J+AOEg==
`protect END_PROTECTED
