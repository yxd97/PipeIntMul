`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TUqnGsvKiV0zAhhAFSiNBKMCTl9Myv2ki7w2g0HnVID/aIwVaEYa/dimlWARwwfR
5PlQf7TvMstXAkyymHux/aLsqqNZ2fZEB9tKVG9Pv0qgi+Y7KeSm5kKwveXCTdbu
ioqDt3HUb3svQmqfEuSO22Iw2D+vNhDB3Pz15baiNIn7BitCPWBuUS6oYIrO+KSE
ND7SMCpr/9eXzG5+NvPE/7pMxWVknf09fQ74umjChD+kS8cdV+Nw4/vulYURzo4Z
z5meUJx1ji0F2ULMR4Krw1Dqh4YpDvVS6hguiaQ00YiOcqHFADM71jQEHfos0n/S
yxQXymllWOkpNQmJ0vHkqg==
`protect END_PROTECTED
