`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kJzfgICYigs5VbwWSGcGniHoDsE9jrQS+CzPUKq3rSEsL9wvWNHpoAjm2Lbegneo
qHvfk3ATxXAehUUlN3zvb0R1eyurLCK34U7xrrsAWFDhe3RutZaskllul+mBIg2E
Qo1dDcrl1ox1/I28APD7Fqzz1oJPcD7mcefFWdBhWpnLIbzv1p3FupH92adJtyFn
a+NuyqbTJmRvuntclM1O6BdIXIuiOr+e/KftAYlEgrVNs0MNi/YUdqU4kG8aRvxq
KOHSJh2073blSvMMGCwXtd2NX4TPcI+yPBXC0pQAe1TAvB/z1MwJN7iIg5kU2tv5
Uz4B0NSXmfZrz+E9xoBwIUhfAsK4WM1Vv0bbhbjmbUaLRBBc+IrEA3/pCajGVQnX
UBrosxJAMjBAxdjXbWi/ldDN39xtdaumGwsQb94yl1N42i+Dz/hEmCSIjDxgKVGI
t89CG2wJE8JPliessEk8MLZm1qpMB0BVktmr4f1FMZ5R2rCXVK8ph/uAit8Hmjx5
mWIHfH475JAt8pKw/OuNKrYTa1DQ4xcJqAn5S8jZaDkSUz023iaLthQRmX59HzgM
MV5QulmJd5mHc66ub+uJs94iFV7wFlFopy5xmm1RKNe+04+yHByu2cBl50i2walO
cYEFOWTAGwvu4gXKfiK5oEYpsQinR9LCSE2+d5yihfSE2Gv1dLsfBjHVdgxR++I2
ZEZO0MAfOEwu6yXPJ3tWQ9zs1i/lAy6WWJRV/gaFKZ4=
`protect END_PROTECTED
