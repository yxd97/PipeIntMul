`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJYO1M3SZt7ubMCovvoc8aXGkSaPdDJ2U9O271a9Dy1v05CEeKfPiTTQ9J3N0jq4
5A91Jjmc+cKUwN/Nbpw8/+UAF2Vd1F8uG9Mk6UQ67NkTcErOlUT0wvfkEPV06Jea
5rlw+RiGTlK0GWzPuGOXBUEdUqABst9S9KY6GuNE3SNqt6Gwt1uU3a8p2Kde4xCF
n1PVkYWJmFTyEYNAE4VYeYS7C2+D03iH2BQboVYsh0xPoBLZTDKkXVDvTR7XZW6t
VTplgWwsH6j6s9sVZFSirvisUGR/SD0eCdt2g4dsjihMFRon7Xe7giHEd76LMr/y
g8fddiU3C6OVz51W3yBXMCoiwzrG2g1gi5DqmOSaLyXO6Ma/V1XjsyNlozqVzduR
kpbACF5iH42COmuSQz8bRqhWkOJEffsa2q33prVU9Tw=
`protect END_PROTECTED
