`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qWBaKj04so6VQ3f1LO3Cn25chF67ajY7D/LxpfwlKO/NQtVVMsX+pPHNLGYNgtcE
SG2s3TN5Ur5Fp3ZAHzXZPEXMNPlCX7ylP1at+djvfrS4LqkcVmY2e0wtNe1xJ4Rw
9c7ss3zrRUsAVg++4hEj2YgFxqMVVHFvsdxJX7pI0F8BpThmwzo30tpPS4onQXfw
VOtTOYDVj5wXj7fvs2m63CMqEdKqHgaHr3ZJW3AwJCfPOplG2LHvx32I2o/4aLsV
j3cuo1pRg9MyDRR3nTb1lx4uV1Lh17Ib3gjGiS6od6+pEN/r9+man4v08yudK2O5
7/8uVvgD+V+yDoe+C1Rh7MQQXPzkhpsdJDfAsYRqoKz1x9F2uKRr0P6myRBkAChO
RmI2Sps8dF76bo/jgM+zHJBkOX4tMdMS6bixBepHQtoEARqWS0oXziEknO+Ro7VR
bPbN1c7r2LaYAg+MM6K4TH5yXyGRNQwgJL4KK8BZSRKHYsdJIu1UWv+RXPRLt+zD
WGRU/Jdc6gTAQsvo+8ZEuzTDsHLFd9I8GgZ3ThnUs7nKQ5aJ8fDyZRS8Ptl92g25
Mlk8GzSPoGpDmdqk2Ow/qxP32Lri75pnfAWCBRtFXx8i/I/As0VZPygl/z47aCfW
MNRD8mVIIwo6gOeTJz6FK2iXp2zTeM7KgMkwyvjP/S46Q9gkbn6cl0V7JlHgfOXR
AOzL8M9btrYkD4tr4u+YHg/RbFrlShDHW1nM+TfaFHU=
`protect END_PROTECTED
