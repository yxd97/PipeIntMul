`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6FUS4gQWne3pVvXGeKZPzJ+hQe1HnfbmpaiNnuy4qatx9K1wS8JyT+eIeXLxYcr
5rc/lOMoSDY8bQEYGFpK48BLC+gOsk9/BQGXGbVzaWio8Mg35iNV7oDZBjQWD3xU
XtKNVg+dP9V4CRLMH7EIzqJ178eS7qEx4q56DvlSIX60xUrA/weBpl/Tw8lJHuc1
SK8lNBIt4vdbjCVRTviEzj3iAtS9iKJnp8ibx+AFdJjG7gh7cAQFvs29IKC4iZye
Ludm+4za/dMUjXi04nys8Q0TlvAVATDIkQZApVhFIrIYJ29AHkpDBWiDm+464pwz
+KGoUVqkCg5IsVwtj5/wuwB1KAhB0si0C5PbIwGPgCbCUNFTl+3MDvpKWe0cmrfL
G9mofuaCQCmC3P/oqlMTcQ==
`protect END_PROTECTED
