`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
idg0pTEfeKZzfu/A2wrWwxLJZqDDCLcl9IrYYWdnJGvfMq5mcDlyDnqXVFa+up5x
T6xPsoRJxNZyYwTFFV4M8Tb14ft3jYj9hMr06FppO/TpKuyeY8D64lJqu2zP8GqO
KF6pucSzH8bCzu3gfXpoheHImi3L43fvEZxOJI0H8OK2VBNDNWssVRXn61yYhMMX
SDKuOD9ilcVh9/QS1pp5r4lR+ANGe7hAZaKqQ3+/C79xtOsPYoD/TVcpMnyUlJp/
NEX6jjyFhxdn/1wvPWny/A==
`protect END_PROTECTED
