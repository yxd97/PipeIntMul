`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rvwj3hsdPvvBuKOfCdlFrfCwas3xKXztT9zuKqus71QqB7mDaLtYwW4lAWI7g+15
9f60pEniKNI7bazsxqFgqwukdty+AbYdubAbPe6XTTZ1dsyXqWPIeNyYScZvbsWz
EU8fN9TmWEGQjzh8vSjU0xdMCZENj3UwU0VjR6NU1mGdthugfmAljhahLpHfemFr
oTVB+9Q22BZh0FpDF3fRBcd25+0ULvVjSVN2Q+E5UZOBbG+mAaV0qFcumS7G1H4R
0FRRTP60IxncPqoTqZGdzpUYn2gue4JBReKQcjDihiA=
`protect END_PROTECTED
