`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zDzSeyvqYxUtQxQLd0+CJPe34nHBISUA30Ainyjj29Twl3T2sahXw9m5Zo8t0yuV
ur1xYpN5WfbQxW+Nswnk2dfuvLNRnrt+spBb/S6QsH3J+izV/DrMosBnksAfF5wy
kiaI/VcRjKVNF0RAdBbbrv7HPq4cCk3qjvJ31sL8OhJ4aXdYb165mV5FZ91FJBYy
2cPPBw9DPayBCYmvInCwzv3X8azej1MyoiuHuYAzzEjeEemcf4aw6uEO+pPoYAdF
PPj6mFg9ClAhXOQNgQG8MgLMW2JZm5rSLVtTnRa1l24CLxq9yGyxdMW9BPObSIKG
XiZa5IIqDMZjc5zqsBTuo58i3xwFs+adAULqqbTtxQ2lDki8mP9RLjRp49gOUdOC
wfdnfazjjnpateVbDuAvMl/btgI1soiGBSRAoH/oKSUY/9ZHk2KFMnCeBQWAtOsf
`protect END_PROTECTED
