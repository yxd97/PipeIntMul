`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+xI6g+NVf1ZXOZK2pCfiD6pUrzzuTnAYB3LUT8zgVR5cqpXDUDPlBUi5YSqWHo6
b/2foOhf2TTdIxw0JutLeXPLzMCMLyvCTxxArMqG2iQdyoa+yskdGaP2e6yUzlti
4gpKwFGH6B6XgY8g4th/9Ej8/RX9Rx+qX1piNLB8mB6L8HpyKwrhW9GWEmTBTw9y
Klt9wucqIaUYkDM3OyxNgDlTORhiiVJ/a5IJRjAwvcun8oewsQiIpjA9qB6cYiPE
407F9nE6o8qKndxnxOLPYUK8NnWWz6IDwke4Q76vHo6iZ0tVmsc9J9f5D6AaVbN/
e4OYc/ZGQeyBRF5IR/Qxi6AUQS/05/fJsnQpbJExaztTH58NOgMka5xRtv5DRLzv
JY7H1p4hrJdMCUkmjQAjUb+iWCUxbQXQUeR51sGz5vRWmL0F3yqeWFbgEZjIReEd
NxhTbwS3vIA6zcRdPGbbM8yCmjyne/9mXxZT+mWIZZU=
`protect END_PROTECTED
