`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aozCvEiWtZbfdnuXNJqJGg+/lDXYjOMCa+LK8d+rEY6Dux0xi9yGuIGXLeZoTC6u
tr0n+NRPhVtpX6zD0lzGncRmkh8+1CZtLcZJVWKkz1lN51gZKEiqi4rjOohdnf7T
h+n4+0zj7XINGc+/rgWhbOCTGlfde18nlE2anIqO8jnh+UcnZ+X9SzOWs2wQW/Pf
yljdw8M7x2FKS/1bHsFAePMWJwSuVQiEM7xaP6OYFmnPlTYFuH+OmkYzhnikMSsC
8mzejMaepjRrpk7mfrD4SqbEM0M3OglRz1Z0A5hFPNbEnJmL+gwadiSkmalbnxzr
GiRbAHnpUmyhw1v4rRKPAhOpGKwe4DzBC/no0wDE0UOMt53nmROLH9TIjYt1wPbd
usVtarEsnD3RQlDfdt9TmEUDmNpaOo9+w174eCyOjPM=
`protect END_PROTECTED
