`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lJ+QnuA44S09IduEFq55cksPP1IdwR1azP5PntJXJVwvdOH+hvaeaLvppwUvl/3
LfBLtYVKeEJ+z+WgamJu1roW+Fds2UGz1FtVN6f9ol3tEEUU9o6sZM9JaMgzFlGp
5QjHRQk8C/qwvBakGK0WUu1nculvl5ZFGXlyLElzFD4AgBvNJZgl2O4MpWVTKcnE
G096/caEefAzSEfk8SWCY5G/mjPKvAutJte8ucgS9LAxRukZgGPgCSc+e9j9PGG6
xsl3xpGTKIJqWT/4QXtdPYQU5XpwHMOMJBksm9fviyH9pKWnGz3wWHa9OwXgcHUi
vy8YaPIDKH2ynStqCtxxK7zKgPz3O2SUX9CVFa3cDTAzhB46fgj22ZiPUf63zIRS
7m6UNUxdp4qhKixTyEWYOVZ/jygMr2o8gv4UpZZfpAKKCsIUxv6ItJDz7gzWpBlt
+JZc0IBHwcumejsxtHpAHmcNFkYaBSISXxsTW7Vfbd197oVx7aTTyYurGKRIz1Hx
SIH+/UOzPauwuewFmq0sir3iAgSCkh0ZBheVXXrNc4Rk7WY5d1J42xZzYjYLZNpv
RoQAtHbYZxcZDUfvYl2AL0QJxu6FK4jRFro8md/EOs+LJfJcrxvQDbTcW60r3+/2
GWZ/4WigawkCm7A0GORqY/DHICWn3Fu+VS4w03j0Zqh4NG9da55JySc2tz5V+vKX
OoKnNdH9GWYAKDcOQViCB31uZcFVOIAZdlTN6AC2dc8TOpZ3VuqRVp3mG+iYfLJV
8/wKxtFetwxsBC1NltJlONtTKVT4uDVculPCUoWRwvfixlu/bWiP73iQMMaMTwi/
FkaCX1aYxAeJK6ltvI7xZMDXDQsdiiz42t+XzR/nx4h5IwCyidrQcGhWWaWqB3s5
NUVcpz5AqsnZ5tJnzP7FEg==
`protect END_PROTECTED
