`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fgHkpIinIFzJ1jeBfmPLWAfZcg9NAnTERS8h1ON0+FnyjjvvnyKkMONySH32xpq
GWYANQFyW/PCXhqgusjIL7S3c4FDDt3n9lcA8g+FThPmvUrw/VBmMUBJxmutb3A+
mzVJkmSyEv5fFo1cenP3oW4/EgmldYDlomqgEvXJAO87B++CMx5uWIPdXjHHHwuh
x9lv0A/Vos3/x+0N1IwGpw==
`protect END_PROTECTED
