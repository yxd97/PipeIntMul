`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cMxQEo1COdN6fMTl5uhN8hO6Bzkk+ZPh3uhPVsPKHDfuul53d6OR5rHeTPOCiaSg
wyaZdnhbxRJ6P58IUaA0cCVtec37CelJbdN6+eOpX3o+T0Q2vMKGJDXKS8wCAVuo
pSs6dUu3V8wppzgVbTvFAJTsWC60/g0ilZ95WY5eZntQJujrhjaG8WIbHm4Z4yzq
VQoADjbLB/92ofDLG077AQaOh/R7gGhuoTyxzBa9Txt3oCeUHnGySSfIg/HX0xTF
6t/zxfHddop6f4OK9KIV8wJgVpVnE8zHPgrMO8v/766ieyJ/zmOQwlvnyAbAbnRn
q/KWPUdsaeIeJtieJ27FyjT89h4ij99EML/jrT5jPBfmXRbDhVT91tkqX9DXyQa8
P6uIz9ygyw6TuLW7vEMg9vgtCwszu4euHnGDRsZNuABIH+Ac7vOnrYppqh+YE5+D
6nCKSfwP7/zGdiE/gB8rwbacV1MuQtUraxg4T7YaWRdM39k+SdDTog2Hi2C/zGkw
gqEpuDM+rlV378VptUq/iNQnx79AHy8lYbq/gcDqdb62U40QKLNNw/In8LrEIrlj
My8LyVaP96AvGCM5H4BGZa7VjUJprCqBD7gbpxlap9T9depJKPxYlPHGGps+ig7m
qP28yFfTsLatTRZyIGbB8CZbLrJrXxFXpNrEzz8Gcust3KghgIt8muGUB1BULsqI
fMJ5bqI15dXJRqquu0zIGvN1wi07guE90mJYVxGF9R+LZIeUcqArJ4kkFpt1g/Y2
/vYVsJiau1V9K4hg++7IK5jZdKaORJXmPzP5n5V8UJczcfqulqXAEk4ercdBouaf
n4/YUs8UC7C/nNu8HnIxPyO7uSWAApQzS1ahJJlddlQ3VP6VFuPlJdebSGBXdxBV
K5R7pLM4gfrvt07VatB+TW3zjkWKMxeNe5lLMxnT8LHH7LZUwskNCQydKq3AYEHZ
UpGKVjqLens9BWHqfbNUM1+hbxgzt9s510bZ1CkNTvBk7La5ZxeSJn53Hpx7xzJQ
yU1qyBXOwaKVXZZTTW48T/g0jMDWHHsD49vH/dPFfkDYk2JtdSEX/w+2XvXif/H8
h2cN977Wb7rDKz2Xn36bq5RwGKrkNrNHGttI33QKEqs+BPLNfHjlMX36cppweDyZ
TvGl4TJWtR/w5PTqNIrS8ReT2Aj82/0U1zhAQBivUcazpE+I0b/1Lwl5hW4C6jnI
05koaoiFOT07AAM1zn8GeiOCkDYbX3lhNlk43sW++kgUV7luIOfOA3z6RvRugXWd
To+RhJ0HKxe/4JksEU2YPow7TusAaCCTY6qBkXaafLlTsz2UqGF39E+2JMrqrwwW
wpXg/aGnI94eXahq3gh5NIXyiQ/scaYQ3dt2gac0fwSQ3/PGojhG2ocEjj+IhQ+O
04aSXBI290lVkBuMfJkk5MuibhfHeRrkuEmetj0sGL8RxT9wrmRY+kCzZmOGBO8e
389IZUt1VSSn8oYBtwHwx/VD9uaRCLWYfKXdo05nVnyNIv48RqJC7iBHFSm3JpLB
KTtz9GvKx2agbLULClYc/3qnH6ybu6hgW6y+OJ6d9Kky+YWvcTt/WLvxlRz/aVCw
qMqaWlLWms4I7r2a9oKP4xmrn4To4W6Xis4zY1dDUqspvQqNtWufVKVNuK4tn19z
T1i1dOhd5jbCsEroeRgm8CeGP/M2f5OqsOWnjWvRVT70H/faAK2h3NoCgoOZbGdu
nMSGjhaO/IL8ViGPxC5aLqXwwAdS10jNRxrpa7xxJusG537r9D/m87dnqMrkK3g1
HrcWwzZJktNbIco0wi5ntJWYQMPjzhMf3qDs0oJ+F47Upd9TAWGmxGHvvAdhraEd
ioBa2vnmXyfwEROOQKEhnlxXpAlID1cXGIGEsOqRhhXMOFVUXPHq+OSFQM48NWkU
tpJuWW2iFtO19ZRP6gtwLreiEYv+/MohajnS366JDuiyAW+j5wTu9My7oW2R1wCJ
dmMHf3u669TnYBf/tSjW+C4aWBFScmuVTeM4IsOj0mVA7jPoXD7LzOzHAW9IJXG5
majIz1Bu734DclJ6XJrFuQOlrsPtHOcTYjbj9goECqum60KroBVwcJuUbIL/RF4f
JGYGJagsUMW6HYYheQYJTLPOFum4ZcyRVSnYkEvE6cTY1G/hDW9kBmsYpot38+Ql
90/QwkL8dsusYIyMqSKu+Uczv58g9bG7yD0JJnGTaTi9DrsXqgpOpDDtmkDOABiq
MEhO+cT3aunfRIq92gR7Cj3Qj3/G8PZXIlTLBzYQwgWc3DZp8Wos2bC/9KH9Bgzu
NC+agRGLCaPCw00uY1Dj8teG9J6/lSIuJZJrgdMtuU4ENdTpfWugOG4spXgGV89I
g2+XyGmCNIyMtYg4nBA2dcnZVqRWxJz/hG7nUPbFMzlSuzftYyHUfhDz5D0dT5kV
7E0vPbJmbqCQjfbqNmssW7Nf7+l2l0YwT1zf93fP+v04eXJTqeoAJcnqteBgyY72
i2Mvp75VfoX28ZjOUZfS5ySYpEcEE6kmZjmyQ1FwPM0AqC/kGv2HvQmWZ3ujGnGB
l6UeALT/WBpJ6aCDX3gxkx49CIQd4Bzdzr6iWVyhMX+QPdDtEPpO3Yc7dQulWev+
jZCuZquDQ2brOf/Z9RguA+DIQ6tuiKGwnTm7nxJOPrHic9X3vg7HPmWX7SHfU/a/
yCpz2vXwUHTKwcB9OsRYxEhh+KW7opFKAGupaI9rS2jQL4YtJGTUt7c5PJmmVzRX
NMPVgurmQHop3ON9Rc2Zmhg+VUtfloONHMvHpVhsFzunMfoKrqLOn/pqVol2ownI
U7za/ffJLeGeYl5frHWxfuChYc0hrvVPEBnR6nUIwgTW9OMuCO0MDHxTnT+z09b/
ZG42WQwu6ltXHLWgidr5cq7aqAjL3S0gFk31C5P+yFDkHv4tRBbZpOiUYbrrOwyi
a1+o/LdpXpQFbaZ7gSu/Xw5ZKxnyGHU6HoV18FZCaZ8BRdPYQbJEEqikdc0dOljC
nuSJFhG5a5WgI+PWIig1iK181/8+ZZNoPMAj+GpOXZj/7aGOaOxLvsvxXkiyNWI4
qrfEzIAoS0gmUKZG7ltJyofMMFp6gHfVkBUCxakZpEvq1Rde4bwazWf29CEZ5XCf
N/BddRlc8/s6oJPdhkCqrn0a45YdMPjHOSy/Dp5htZVOoOHm50P963VnF/tSFndf
tSkK/EDfRlPB7mfF/ktIyTGoQLEyhosQ/yQXKclm2mxZ2tNEOkwsuRQzi1M+NwGW
DUjQpNq8vU6wGIo/6npDTXUCw47NnagWu9WrPmXf09a9GcWEOmRXNQD9hFaLYoRF
V/DDP5rCld2X4Dd/9ewBPPmhjqzsZf+707oqH0Ec8SXhBVocJLXsbobqDmMHyHNr
5fSTIw1shV/zNGsUnMy0R7LjFWWbBIMnesWwhQs4/PQtQ9bWxBj+B4bRb6e0npvx
P5dNwPFm0Mhxe0lBmAsli7qoBwk7E0W2DXupOMU3J+arA9P8jdNXDGyH0atd3ufn
BShplwU0NPf9YEYIXpbpYpxMT+XzzQvqASDLCB8llURR1N3fGuVLOSso5JrsCuT+
KulAmdQm5sr2KXPPyNzwHmghtZ6NfJjjqce90X4NcAXzMZClzeiML8Bq997Mc2yB
UMGcManWSEApLCx/FnZyfSIUKoXHt4J9iw/Yrn0nu97h3XVbSYk8slPG2VsdhOi9
n4unWp6fsw2q8/Y35J3KxKQk+7jMk9ft57zKDgBM49ltxwwLoFFPdw6jz+7HmWFU
rxOV1mlOW4cp80eP3f4I9aUpJihPPJlHxTmWrt6TzlC70H0S3+MQlDq+1UnSohTV
YMElZwJfwJHwGYuRsEeNM3qRJkILZy7SK4nKS+1HGG2E+YG9QFd6YbM+YI2yVv3e
y2bPogPjPuCIqxlzfJVA1KqGOZMjJkKQr66BIZN5dCidlvxzF3du/RP1ixxNvPj3
ZQHFeYW2eB+kOeoG/zs9o6A4K0HL8q8LPgg0Cipg98NXCbdUcZfthiQqJdK4xcHU
sqcPOOPbZ6P+KXqcTMRzNwpuISq6Gh6/81x709Fto9rVCa1fczz1foLBJzIBBA74
lP7vr1tY1C6ecITOKorUcho9qcFNam8nUtI4BrdFg/0mYuEA0lD8HzxKYcd/4i0M
E/Vjlqtqm48TNBOnMkSNTsf5wyeZo/JeECkSOdixkBVLVePxWdGLwpYYjY4urkxS
SJQ3hmS5ejx/V9CdscySK7uaO8LtFKkMzvcVaH2xG8V6ZaP5RocYI8bdtDFfTeKE
rCpo++7WRm9Y8+6PSXdT5I+DFXFtgJJg1sVwkjMQY+SAQ9zKnu3obfCIhYjGenxP
zxqZ20kJwxYRNShn8fh/MIFKy2qrCDO9kTNfXmX4X8c823U6dYmLHqoaCCQMS6r5
7f/YMAg1GxAVYCwEgnIBQKa89XyhAN/JNFvU0el4j/MMhcJPVwJOa3WrI19KaZ7Z
6hdWloh/iCWiuvdXmNeDxtRzlumn51kkAj76GXndUbmDX7n7fM6o19Wws1PiVBa6
tEzRQ5Oo0cq8fKG9SV260bTRNBKmJaj3CatJhqcJP27r90k2rdGtoBIqH0KvDuyk
pXFgtSVW+ZZ49A1dTrKHCtFwVOwa8AZZeOmmXRlYk92acv/Jv29ITbgYQTOl5kJn
CitvdMVwt2aWlko2WJU+wAdxfKb3hMg6u3V4zYagvW+NxXRcLQzt0bbefR++wAd2
ZTqEI9fZf55mZwALtfbjdy0pzClLMFd10vYPO5nX5oDb+Cmem6srnqXBWSWueEBe
pH9WD1/BvNYecAmUaDOr9n/MFPRauoccEUmAreVv76B24tr0aiUAQRj6oggGOfYb
6zoU95b6srdYhODetLULYUR1ywpY+/6SAXr1AEOYAqBBoCUjt/scY79Y75/hP5Gt
+htvPsAC/li8EykJBKw+fi2i5xKttZUrdL6kl7TNhpodYRIC8VqTy8uW7yW5CA0K
SKi2ZYYETVHnSDMhl8jYka0CFfqkm66PAg2eXBapT1YFU1/Cgf7ZmdLohvZFjV8H
QoxE60vpIm4714S6lZk/RTHMGEXVI4HLhsrDMcEB8Xb8cFNORxlVL0dW0gnoQbRG
zHIDrOt8+qR6OaekXa+4rTF+zWIC9CTgNaePDqwFbAVadoxT+bRZ+pJRzh5AhcXw
kq4ET1Ys6CV5NY5O523CMR0/+67KkEhLgVP70kIzDXMRLhCBZZVGICjg8+w/qPX3
9+GLIg/zbCkGtKTQAoN8+MLOZgQUytwjx5zDa/Koe21i+PRdjTjz05RJuGQ1j7OD
KFxlm9xUTpfjXcF381cJzSuA+c7M+AS+Qy8guH9iqMf81z2pLEIwSzYD54HyC5CW
swPUORjCDf8oa57NqOGrRJI9v+O1l5Di2mfUyX/WWaQj3cTr3esA4824QYEny0XB
y6DLPHsgznRah8PAB6PC7N9PF4uXtWFWqfEkrrkW8kDR+V6Z3KjQdbeqlTFExVZH
6CAMpD3XvOW8IEwIT2+tmE2/IF+FwMwSXlcVWZ5ISUe05tJx4zMrNgua6P56qrCZ
fSAXsXSgbXikLJPHaGTPEfuKZ3i2WevrciLhVP3Hn3I7am+ljulGrZqoZIZFEGhx
27CWp//apdMnWZes+YWk7kdG9FTXXMRwloAPx+B1VLZr/vPy1xXE30OvJvEHbXik
UNIaGEDY5cqRm95gBjyc2gvFhAztsRsuzf+9fJKPaa97Ot5rv2PYerk4YAh7hseR
GfRhwRt8M6C8w5kMSvJUq/MW/OyJJRM8sVcSJsM7x5c66OmQHPjeQjO9NROJRqCo
nJrpd387kh5025fTM86WRZjsqZ0FmTw5tgPhXamOY9mZLalN8vFEbWwaU6zYwT99
QwqhB8N6paNmkdLBk6m/hpeh3eJLyQtv+RBhGvmcWwRd6TGfLQsZld+sM1bOXPHe
EPLo95vGIC1ov2EF136m8Hv9a/GFLTKv1bteUFpbpcvjj155kmM5VXVOnYnPJfrG
Z0WXPrW4vy+XHDSBMs1+SsEYjH4r8aisgw5Th4vN7ktAXgMX8OJH6Qw8fE8PbhpD
g0uxRuq3H/LDkhcK3znSyad2l1qxYcNb3gPF2w/HSToVZD/12FqCSN8+IifBt9UL
/Xy4bAIvKBSBNplVK2jsD+2o0uIbsUwlA162+l8CBkbORfopWFxPMLKpvdc/HTyQ
ym4Dw5hfKA2jtFYCjuO4RWSuxoX6fYBUVXLCEaAYEIrvM7iI69HTJxPWRfH4g8b/
vS9fNsjt4Al5q4F2K0XlSR6NP0dYkJN2qWVTZgXRm5+1FWrt4nboGy9W/VYCn8rs
zizVNExcsIpb7BzmxFS9ef4lGtZLB4UjMH/fbCt0b3bZxpPPfoF7J69xfKu9EjlZ
0GN04fguXxe2RWSYFHalMBEIjfUYIEWvzVM/CB/j5Sle5o/6xpFwVnuV0Iju1Ibb
4pyg1BQ26n5rnleuSIm6uhnkKz9HqnNsjG2DOKz7U9cbgdMduBF4cr/sL7bAIu3U
tHo7G3cIhvWfePR18/XExBh1jXwYuv9QFtvgYMbr4mz/zXsGk8S54Zfsj7JvVTPh
88ugqkYS64J9lc/GsOjCoJl/LxMPHMvxMkxgeawg0c6V3JYVMlSwJioU1nxvMacd
Z1Q5cMIyDhKhbROFVq2qh0BbuiFq9Vevo+AFe8Wuibp2h0Ijc/lPYJvxPNFyfdwi
SQEVirc1oXpEHJhIjbcTt8jEkICYlcB8zrXjk1UEra2b4zqIDzFZjpXI2mrbmapb
yVZ9T9EZhWazTXsRUVY3QTqa0gNgz3a/1QWz1W/YEJwyiJ79rjwfFV/WgAaUTFQs
yMegvL2MJeDeZhklud3vryHnBvw5hiSgopCGas0my09CapAaspr4IH9RFv51H3Xj
6rgficWVaiRuYWU9ESBR8qEL6E5la7wMagquySBE5/nQkfnAoxkCMHcNGwChqToL
9SCK4aLY8gZ9IXakf2z39iUh+31WX5TR7yKb0Sj7tubEM9Fagt/XYZYFBhCHqRBb
rsOyKhd1aEAIdtUA5v6X2kKruXCLhjxlOcQSwsarKOIFoyr3EF4Ugk7YctlkgBcK
cuAZugjA4pubQytuFSltOY3IgbjWZi8YzWrFliU8afwHKpUD+mO9MTHUA9JXOxKt
PELspsbhTbu3fG+clyLHhfNw4cxGnk3XzY3Oj7i0PQSlc0WVU8k9Naya2DfqfJ5J
QtFYtwft96CpvrczNYBFefqISCFxzxsQwWMpYPMUCFl1s2pzusHPMjzGUD1Wn3zd
iBks1z/YuO7sKkX+HW/SBp9aMCHehUxL5v8tQnYkwTc=
`protect END_PROTECTED
