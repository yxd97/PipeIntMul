`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVShxUx5MafJa3QoZnhodu10cnrFGqH29sIR8iAmU2a9sn8KK9hSolZrM2+1Bxqx
Q/7e9Zz+vdZ/VJCKNufubxU8s749cLjLZNKNUtPnICJphzQ5wUW7HmtQnhf935oK
uKJqAcXupZzrRTN6GJ0dr0LKVGBjotG4MtXHbUCWghOB9xU+HBcgN7mYO+ybEDpR
PESZ5LpeVBd/gAr9y9akjCniAOWmjhrLncLGkvY6DxWk30gJ29nLP77muSR1ilr8
UjeLIk/q+f1uTwQ4eEPBZfvbkRHoVAl+BREkhYLAc32Kqcz1rmeJrufN7xO6mdm6
MSLKddE3CNiStu6KivtTzDmASQ1zDhzWDyr166cQSoZS9sNAkUXbD8ycscHuCQ3l
Rs+b+xyJVVb6QJr+zzXxba8NiR8UUD0xlBwSyHl5pwljuRENMqiPpPJw/eIHopXu
+ZF+MdL8DxEzAY0zyJyZ4DoqzV541JS6t9ILDvw1HZhFzfhO/Fepd/U8E9/oH2Xz
nxVFMt88GnvdAULtFGYp7TNV+B79S2DUmTxMrZTj8sucasrI51jIZ0VDObdcBvo2
AOKjRw0PqzHBCbXuPZB3W7gypioD0DyVxujdmcZGRgJuaulyBVdw9MyUDBBYSLFx
FYVEl5mIqutuQLtOk34xnAYit+yi1BNS4FNQY28saAneLmCAqdyTGjaxrqpYOxPH
b2sFqxFzzEJT+fxNRg4YHZHV6RhGrjwlXIhuJKWF3IrBAj6KUO7YJ923T21qnXoB
Zpx/VqJ2bDxiwXDIBlhaYq44r8QQxc1cLu4gUDv9+G7tToD+mYfQ7zV9JGQlTjYG
eseBJ5LMmu0z0BFyQk0x+W2cTnhXMyzGBELsMbwrmQucLg0GlFstwmVGao9QQpu2
KldixgsC80IZjKFQjZC1imAU0yXoS2MoROeb6nPj261GkDmeS+uOg21yIUYzhDbR
rgU5jqiRBgnng9fghNWvrn7Kjhf0YkJ/re4OMBF1rvvSrCHQ+JM1Wb7MPg5LAHMT
A5dNxcqoMpFofT5maffeohQCX2EqrbI/4gbPgcjbCUy+icMwVL9HfB2xrXmYeQ3A
2nXQ4xAvLp4nLWdSW54+ZpVanFW/wonFAJO1GgbNDwdCFezYc+b0Um9yrRJLBqky
WsybuJvsllEZUa3zZwjiPpqxUy/n4zZuRYjMQEvYLfjQCjfgyIWFkZoaxV4KhdkZ
cTKkqnpLddkVd/IYi3DQuslbfedVIEFlDrbgJc+X9ntXDAlYmlsLULKV5Mea5HO6
Z7Ds1H0N+HFUJsTXSN2PIB2Fkoe2vBPltPC7JTRejg+0lRSuL3Lcl5hiSqfM2ox6
qduaE8T/Lhu2UyHpQUHR58KP+VYDPN5tGAEG4zlLbUzlhc9G8pmYsXXBMOQDwuP5
U4V6soGcXV2dEq7WaRpxXg2k9HNexV+Qe1ZDjKnm7uiqXD7txOfk4oAmS5EsWSkT
5l5/GZs3A5L+n8LUxMM3EHaL7YyslV/ImoGydqsliEJPyXwipfiiLwd8whRIuFoq
tDjKKVJEGSRl8oHGii6pismBejypEwo122FMz7eUZ4mVwsj/ILvq5AOJZYE/e3LS
PNGGKfzSvQBC0hoF9o1VUZ9HvGuW/uGRa2CRxSkhEtNV+IayEtA/+s3CpeqfmZbc
c7N7XKVl5a2jCN8ZYo14rvU3ZeZ6cSETAiGyetKZuEiYpUPo8Aa9o+4AW455tIVb
AKYusQ8dcGrXspHGyZtVv+UpNNcWhdvvF7P0/oqBAVRZvMcNFG9MN+4pmIG/cPlb
1VMU7UBb2ViKEvU+dbcr+brEyNKZmZ0QrGIz5bZ0T/POGoTS3+RoyGMDawax5oVi
AqMmHO5Yj8bOp+UUSxrOZGyrLd+7ndrDBbFI06oV1NeSeAStkDP7st4q8UzGY7jz
azhbQTLUu4AglS5BZRADoFHPXsmynqvXDCFTqT3+PvnnCEGC/dgfw65Tl8o/evcv
k976H1ArufXlWbP11ecYDh/hWOtp18anxTNt0mM4M8S805pIHDv1Scelxm+PEiJV
89ol/OFv+cRShHvfJLergpnEUCqIA3cCr38LZTzBwvSLMGf28VUwVDrDIcCYIvIS
u57cFrcLsXPg1neGTqBWYsV6M9hlaF40LXXPTmsJY9bLwPQGZuPVsLaLHmGn7YB0
+Co7PQxLWCVp3zJbFM4sfvyX/h2+PQbMo/KrpXOGiqR4MYnvO9i8wvyNePJgvI+q
TI7v+s/GH7UnZ5VJH3EOeZvCWZoHwzlYhdm1F9dA9eD9PIuBNnIj5G3bmeZv68Fu
0Ztr3BI5wu51lbAAnrMLbbjcUPY6H7+kK3gJI6E/Mjkh9pVISQEoOZTRo7cmMSaA
gnlhfa081p6A9HoO5asSxTcSWRkLlnA3jZQcMG+eQX4nqwbYkskXEizXcnghuP8r
`protect END_PROTECTED
