`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iw4mFsJq3FhD8AS2WuFJcHpX6V4bxpLFg/a6Kkwnfq3B4UV14LLshUvK8nqqS9Tr
LZggNjzA125m0BgWq1CGv//MSde/uSzOmIwsAhush9Tp9lhNusoZTNhJmGxagZmf
7kObp8Lgm+earKq7WXGNbW3PJzEL2iNQtG2j4xS123886pzpeyEgoJvDPpTNZF3c
4iKy3JOcpO1hYriOx2XH3/OpX24uFVr7JzUnShblJM3u9QVMQkM5paMXpWwMPdYR
6eku4fZn0MppxWJKEz1bLwud2QuTjK6F9dC9VgXkSChHqVTvVIexzuDPw1lMw1Jo
D06o2Vm2lMPyBv/wsHo70+D0xc+Gwa9jGYSMxpyzHQw/cTJr1pZ2qUDhWxl6EY6G
Dn68Kd2rxhLdWCdyqgpx48kE3225ZmKNcHZsvkC2+SI76C3m4jqvfa0iFLhjCgwA
sikGcTnd/Utw9tppe+l7diiEs6l1Wt7ewMU43GrXYVdYJnhhfQysKTgOYNEOw4Zr
H2cU2kXr50sIKwqvBzis9/XfbqhSTJ3bX3ukMaXGDtSvYJBMcRafShSIO7vxjJBC
1eqpiOSvHBoXrpo93Ha1r0/U74nzerfYGh9IBApaR2Nvx7Mcst/nZ1L2Wk/bIogp
dZu8HbkXaA1yKVdwHG53boRfMlv/LAWDT36y3//Vn3b0dZsnW8HPl4CbEjkZ8kLh
y3e/mu0NLKahOQHSJFjBMzLKBrrIZBZqenO1YT9JuWC9oPlVoddhlvwCOpgjscZ7
osd2I9FvNyiRFeAuXqP4SqQG7sQpdscxUhQLumisBKxhdxP0uhUXZq67XEpYLlis
u5o82V6D5ShZDSOpjBYb/sIKDGjQq3kui0t1kKKmz8ExYABk12Ed5hTirwp5O+H6
b2vTR6SbmUEPJldLtIrvtcvPE/HV89mj3lNYtYAGz/EL9zsP86Ls0+eIJQZdZKQi
sLYF+Lw5DkryANbpKZEWv9y9c3qQDEaJ85IlSXjUa2B2M+7fJOB+Jj4rvjeEbyP+
kInU6HW9u+Ub1P2tYJEQVJdMcpP1agQeWd9TnkvDuatmYBmkFlgKEl+nTHkXPQyi
g/SADf3pAIG3FozLllR3hV+h837xEklOpDLqRcENem73r2OKpig0YRib2g4/xkGZ
fojylKQV34pHwwplvVPtrgsHlIcOHrh87RIy0Mzf8V2I2NV5pDLIYxYrKoNNCMiI
/zrHfEJPbXzHUFBvVrD/N/loV/bEZnmarjBfCxbYwMtdS4xtxBOOzmut/LPdI8Va
OvRe6nxxhYWmVoJM/T/NZAh1QwDTRRAysxKf8iSDgWniXsIpWbb3SJoUa4eJRtxo
YVrCvZ1is2zBjYLYeAtwRg8yX55PfNXrfCbvPF0cPWOTzUCXwJIpoKFPhy+KHCvJ
6fupdix9VY2pcF1lsdwkmEHbiK0M5UHXnNSk/XulFnFikPCpcn+uJPuTlI9f5FuD
ZFSKZNkZ+8A6BgW/wZvGXmQg/6LeP7r3d68ErQolBhfJTDFNhVhbqQuc5eTJgENA
lFh6jao2W9A8vBup5U/hR5gThPZuPTjB7Px5LgZfU4l2UwYW89q6HW3a6cQzqeY3
K7GNgRV36rhBTNhwxuGHqyz5uyEQfKthRPU88NvgyHg29hv08ujMwWhGKR4dp6oL
5zsZyoFmKdjfC/0lseugfHFRAx0Eq2uDb/Qb1heDHILQVggfcVRkZxpj//tephpQ
xvPVTPVbEVTs3Fv1i4UW6troLya+Q1BIeFI2X1bX+JKPmyKUMWgu+TLTUG1N4UWn
oVQ/XgZZkYAjDVzHwnkrZo5OZdZxPuUX5E+jUxl27vDEH3LxXsBq+EKtGD1rlv2U
yoMkST0NEBrbaApaJkAaSYNm7K6z/3x9Kl+YeOe7SUvpYNgJNX4fpVIaDh2+GGXR
jnIm61YfwtOWNog24USgp9xko0Q1b63VbEMBBr36fx6ETXOwUWvJWMzURrILk8YC
yYqnzNNk0dLmxS3AYEYTyhQrJjTKLAXODLzZlFvZCHH41TPA0/Dx2I02pn+vQnNp
aGSIdCDg2/dKb36nRlQw80ZUVmqMHsAfm4N/AV6COj+Fp9LIh2urEAAXIRP80BKM
7Adj0ZzxsY/Fxeci1+3QpSdqasVIBQ9WWtzUZuDHb6eRCJW8Z1hAZXlbzLPNhBAQ
CkimpA/sBt98/SXe8UR03aH9xqtdVz9PPAoFaSjzp33GFfcREQ5Z3tjbMQjd0sf0
BLlKQhhdZzr5M9Gu90GF4VKK3mc+H7t7zWiGIiW3JoCMs8ZLtOVpNKx8bpPkPxes
2K9cGjPjae/qlJjBZD1xiAAlX8Jx9SurLKerQ2qwX8HdDVDdHS/OsyrVfsZ/D8K6
a2anCFzzd1KMm7vTfoM5Nz2++6V2N3ewlUV1niRKrO+q9Sty+Q5vfvIjDSF2YFvU
as0y1E3ocCOVwZkUw8LdZaPEO/eHn7bRi6clKAQMG+q6EFS1QtWgJ6W2o1Bwjvqu
udNSY5UneLm6BalGPeoxmu+P43IJ13XlEPiDgzeY2ZgQuQvga4qqnyhOFtWumIiy
I8jUfcQ9Bq3cHBb7Z7YrR/ww3eEWTyeH33QTfSyZptVWGRYy9XxwVXPK0jpXCzgm
UkuN0KqjDNL/HPvrM4+zN5+vIK1Tch1Yquw4uyfmxhiVCyYfeYL6QbJah5IGIW5o
1KFH1yzLv0b8uBbDYYsrzdhCIVRxdro0TiwqDCZY4qtSqavrheeMB1zbCf9HwuqW
nyes9/oqQLfoRcZWs5lAylAe/J3kAvTXUsu196CQxyAgaAfQegR+xCcOjtigIAuq
+3HSNLX/iZ/gsY7qLI6ls9EFkjxMmOS2fqvKtY8mgWbjkUwGuQ6XKMMZteQ+EN4T
miWduovdzcnT0lu4LZBHTlhNeJ/Co9KTQep9XvkedcZ+rcevjE6NNFQaFSBk3/yO
W7Cu8vbcHgWe74xB9BUvbLn3qVxZu99+wWNjzb3sL4BGwe1HRH3oZfJmDadtDX7a
qHJwEFwP3ElxsfyOJBkHkdpfhletu7Ho8u69Cy98MxvCKjg5e7ScwWmpZpMoMvcL
QijnvZeHoccdJ8HE91BS78QXSO/ikURMjMUZ/WGXBaeIRl+/mnryo7oD3xwiYyja
+26e9QStCE9ZiWiBB3h9Ry8/2EJquvtOu74Xd5tg+dlNqxGWV/mgvAv2jg/zdKwb
jm95YMsfFPtcYID6vdwjOV8Lo/XKFHS+PUH3vqrXAb7DYcGcZfb7nmiHT//B0gO4
CZwj6aUHcNAGem4R8WZM26yx+pweabBZlP632WgQuZ8Z36zEIRJaJ4FeX9H3Wc41
3S2f7u/EYtTkWk1is8C6W4MsprfaauvmxE/nBwb9lkp5dnqe/GAvtJvQyhDDln3q
s0DaAItw19yrPxkrEQh12sWZQSGyKp9ZvpSp+YA8RcSX1u8UbklW+jRxlAOT+Td0
gU0O7euDbIn4xQgmZ3ajtsn/5J1ZTU15WUTkxp5pCEGQiQpmQwq7Y21upP6lnDJk
7tEV3CmprTN9rT3mJkUBRRENuhn9XEbzaUNPBt+V9YU=
`protect END_PROTECTED
