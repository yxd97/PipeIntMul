`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGVqE8xYSxw1OTIc2+LUh68c2LkzuV+emwX17v3l0SktvkF289NQhMGmMnTS6nP+
WOcmC9X6Fq1fnR5ELiMe5yVMSTrj7FXonxM9emXw0xpB30G4cj6rARk5R+EYqw4J
8wDXOxBuLhupj03xXAtTyPkkDyo6KH96YfCT7DCjEBH1PrjodIaUxSSNVWz/SMEX
kbBUZ4QI9VOWpPvasoogUJWn5Gn+QyWzZme8XTilepQ/0Ql1gtBZQsVHxDYBC9xp
vei21naubBngTt1vev/SKSpp/Ma3cSAdMu/JkSrhC/rNzEHbs0nomHWBErOcPKaV
zlZ2JjhRYmZO3pYp8yDEDoFmLdCWyLN6j1PT31hyXm3q744Nkow/s/n3zERnoZe/
BUtlWI/26WJZEpdm+nMqhbjqiXhi/sr46v+jw01TfICRqZ5x8QORHRH9I+c/mIoL
ldHiREBpwxW8KSGW6RVnE7Ki4i5MUCRDe2EJjmwvcNmQttse5eg2mKPZyiLd46oi
3yM5HWOkY8T/VVre7VB2/ZZUFkeU0v7BAzJ04bK8qfpvY+SEJbw9mXUUpDxQ9zdk
RLZ6EK7oulNE0qLBDjYMWKfEbY104G8OiOJyLHLGylfxBzBHB4Zv755G/4UEZSy8
qIstaUKE8ShVES5ELy4lHWNu7xOwEdP+JZp6dnILZDRfLZIgXvS4ysnKGrXnJZSu
X6c2FBGicdU8pmk5d9idFxJHLDM6wlW+8qwh63+w2sDDaoOv5+GN8lgYNmkmKzen
CEGSgOANLFAQXu4nBcHgmeiPA1ZHWsnJYkns2/SOZpr7vBZPk7DS7heTBndJUhp/
wnjGWO5OFNY4UM13kxUuhN1mzsN4RqtFaQFrS5cAa1aKedzwRzSIiBACguN129Tj
1w9yttGb3yX95yWzt17qBdTBc4jdhh2Of4t7LXSxWcX+XKngMeWMMVFcfHFFSoDa
odPIiDBRIi17cSZ8aG/2eSHXBfr7t4CGqUnx1f1ZjaC/0oawQ4+ULqwExD4EktYl
9QshGzrqUnn7i2LFQxlm2nuQI+EjyfTvwC3YfSKpkA6hbxANkFX8DgQxJ/iNBb1j
CiVS8hXiNXmHd0dQlGkWhTQohgwRyNb4fOKlOKDPtL5gpiHRWf1WNkLGWdX/tEJ9
ZtCPoP8StAPmUa3oGQ4LiL+YyZTSFq0FimsnKMEnA15AzRRyeiRRiC5G2EX2Car1
SE007F+2hKlyXKHoLzXijHTqRpEGbni6j63Ng2NXCCYt+zAFsUCpUGtCqTkToNz+
3Wsba5Vl617MResmAKIzSwNDaURh1xX7oK/nx7NDXoixSJ3U597phm/q4cjVORYU
AlGHZsdEQZDPTkcN7m54JMO+e2YtzbxEJJLUSLPRbL31/3B6J+b9v7O2vau7uCqL
MUNiOglSzt0kxpiz6zfJ0mznKwgpZDtTn+gEWS673N0II0ElZoCZWxdrYa4kfHT8
0KLlm0wShMCa94ZuYfzkHl3folH4qDKjfNyuShq5uV/9ODZdd1jBUxSoQU9Hyj/O
Uppa7ctsDfCoO48mCqh205yq9D3oXqKgLdSjX7h+jYDRNyPYOpeBAdZ58h8TOymo
kFQMYN0vMREI3T2oIRIXIotZkW2PMgFkHi7P0nrh+PyhckE2JbGZhRhPD4iwnO7g
6h4XGQDaIF/RfDwmu82NUZDf10XliaAPKFgkVeQ4GPZgEI3UTGU2EPmP7cO5pmNj
iZoCiEul3eFtHs79HrIO4QFi9anTwrk9qx8F9DKsVt27vXrHwmf/IYy/q/g+VbGq
4/B5h6/DKlCG9sJMdY8BreNHPDzcbfR9BWYAls7Lr+sBq7V1rCsaYAzR+SKclprj
DYfMfmfWlK5nm6XxXQj6+Te6hwaWyFOGjgmKdg4iqGmV8IfIt3Pi3+I7BqTxIika
H9oZGOYb5UWBPh/T1jFkGmvBxcK1ua3441rpKpOw8DQuglaSCiOl6Qt1siRBnIsW
Sq43Vx6O3Mui0BposIBCIj8tkvTnVkwcljEhEpjavnoSw265Ue7Pb8AY9OuUtl8I
xckjTCwkxHkMZceSa+BNavhPdpj/320SUZFO7KpeCR9jrl1OyxCA9jep2OncaTMM
pwDirLfEmRVs9gzvxS2KyyrapwiFoQJwyzGT1UtNw3ssEnkTeCo3Rvz+mb2anVIb
kP5ET8gNRG1yMjMxdY1HSiNtKiE6uiRHzHCXSrIjjh4oCSEEk8FZQvAWeaGagGXM
NJoWNHhIbEpGV44XJegKa3erKASWqriAv5TteSurQhRdFkdCw/hus1qgNKIgmj6u
bG7X6jOp+4Y4Fq1TWZdtC29mzaihYBQoPWhy9JHuJd37QVO+aSagvDCOYVbSGNbP
55L2+iarOJeBJh8V2cPegGeq2Xtn5449eD3xkAmRqwPEL6Q7drI6nGi+7G7hbvcT
tHdTe5ujA96MWBLYgY2FzpuCzCaBOGsH2P2tg447Jf8cBFEm7YByQ1AFEARJuRc2
M9SdtmJv6Ret9krJGCnvmpI1mq5rSnMwGK4U7GeYdQfk9zgD5yarV2hq63ETqodQ
7YQGZ28aoWDIxj0+w+QllpXEyr1PVHsBmC+Lmv3VQ6XM++qadkaSHDk2mHn4HypX
`protect END_PROTECTED
