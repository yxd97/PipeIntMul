`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6vf16oyL+tfdyvxKYr0CDCT1kMBbxs4TgAkPS7ZnAIPdjY7ygd9xz0hCtnRzS+0N
BIa4kWZoTJG6qipoYFN0rm+uHFuRLsMqsaehjHGC4MgtF2ZShHJo80VLfRBm5vKt
PFLHZBC/PBhPHJAKi3DpFJDhn4Z+Gt2URCpL2y/kxcxGKmhEx/tgaDfQC55Z2/1m
IDYL+eJna/DwshNJ1DcJK1bxj3+clbxpyDa2nE9Cba3gXqJz+aadIHdLGx0dekbX
WsKcaZgCXncZaqTX864VmzfPTdMCn/Qj1fkVxYufMNXGfv4EVFIvqR+QsZyWI2a/
cQ24xcVm2P0PFqIH3ssOy3OjuTaqfRQJPCMITNk1Aj3oLfTFpxX1xsuA19ql9Rrk
uhbnYxNCmBy1R7zVCiDDrI49iZrysua0ZIITn4lLuMd8NczoBXWi00YG9QDl95j/
qBZrf5V5/9O3cYpG1UqA4dSiZ4iZ8RCCS3XcsoIdqqQ=
`protect END_PROTECTED
