`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LzfqWpolrrOuvy9MXehczML41ansDgrGNGDCFaLgEzhAdicDQnXIT1tjdqsSy19V
EPqZ11L0hQubDDCeKEcP4OLfQE1iItZQuUiUdO7jQa0gTS/Ip2Caai9So0UAnvjx
O/0kiyyK09lqiWR0SqaDP+07P4/aCAO4tTZ1IQTIUMArczG5JJBs3IW0XTEQjPBG
eB4wakc6myE3F2Mao57NwjpQxZiU/PXrrw1hypqudgJbVSDiIKLNmYVnl91SEH0q
irgl8LwCdJlUfeXfDJ2V7CQBXOeYbnVqG+ZseSfd84A=
`protect END_PROTECTED
