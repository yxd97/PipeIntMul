`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OgTHnz3LfOJue/hRnKACutLoqns+UjA6lgi+iEKqaKuycdq0AgHNtJmd2v7jbQV
SXCx+6BYSCvHwoPHFhBP8TYxsNQbuImdupnZp55ACYvng9PeRZQWWSRyP2hVokpG
tH2kvsQPB0xGlrBPFJlaYmhuH99pIC7WJ6kEu2obBV0GcMCvItyTmPTJ+dvzG0sg
aFs1gY8kGv0ZvpAku/oguMSbNOaiRgd0PSZ+/aSwiaVXBsON2Kc4TdgjCQMyaeN9
278higU+I1VjxAXwDR9PcTKc2SqYudRVhV+VJrH3ZKL3d42ga6mSRF5xD1diMlDn
f2lii2lEVlTfKbHo1gR7JEpBxXrVAcwft1tYclxff2eEZgVl/16cxXrrfBD2qd8v
702J1LOt+xFD64pF3ZwrcRTK5SfnKKZjUMgnSO1qLk3TtQ8gbiL9r3OCkWJWJMRU
YIZG+oSNR5//y2kgdA39Y7uYy0c9Kq/9W70hWxs1p7MjSQ/vC+IUJeCP1pPj8qpg
UyBMgRbUUV8TitFURyeAfB0PXNoSoRGRISNCibBayrI+EmRLpSyKgs093o/xGZMo
PNebj6B9FQikyvtinDBALQ==
`protect END_PROTECTED
