`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yt5VKTKblX82IbBpszy9W2pHdIcyFdGjUE+pB0tcERnrkJJ7nrSmecdhVIzTZVli
Ut54k1llTfREEZEp+lgdf1ehgkQ2BkaUIr9afsB7zeh43alMs0fiHbrHkT1/cEFu
ZgVWMtwcNt+ZtFrO3jze0zHLFg9lsudcIg/6RpvVC3FX1I9Cf/Z1n5dIKjGH6zjj
nYGjiJaSSaR01ljjT2I3rdCot62Xpp38+L1vKyo+xY7aVx0xlWwI+RPPaCjxxY+K
bVBeW6Mb7AtmoAtMHki4QqeupGVCtTICI88poVt22WgdXes+3ZYk6OtQhagaujpF
XL2nfgOtqLmmVJtbSX7obD1oZQ3XyWajn/92+pMwKSU3oKH2OyKzIb5Ee9eDYwGo
`protect END_PROTECTED
