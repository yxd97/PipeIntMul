`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVeSAWBJqyv7CDQTABhafIfWffwsbhE+A6VRWqu6gGLsFwWDgEcqRPf09xDbcnLu
pst9QQIE5IehxYZ8SYLB4nUagNy7YvJOgghei9/CWRqFyDzStN3UQTP6V5NZjni3
a08H2BCFy70EUwKZIoYjRyBi3pKpLU1pLkM1lDy5JniMDXTqboDkuqpsgolrL83A
lTMo9+pKXygBj8QKjgpy1qpTQsuUVIGJkhEmM47HY8ZuuKkdn4Keda5XCg1udRob
w1hyYMHVPCg6NFE4Sa8RmB1eIpl4u/lpV/Y4WlKmzPg8KCBR+66GyLMBhs2FEt28
jHyzBDMeq4KrBqtpcTKJI2Qx6Tbjz4qYg4Nas11RPG3Niylcg7+yiNfvYY3QKKT5
MIeha6tI+ONwzaAOAk1Y4SS9U3ZRQnbvnklbUxO7DBmqYpAG+l2kdUPKk7B6iLOz
729IKXVieeYAM0aIfwP+Lel5kftoTmZ52eQBVJvcow3tVyeoRT729+rtJOhRjdHE
WxZWzCHNiAMg5TL+RQzMVbmbAwJDJOUNuVgS1nL3PNsZbOrnSXRO3qnpq1sNsmNC
spUXsfgc4iFPoNyCEqRQalld0zpIw0LHm91VnPTgRGIU2koHJUK0qD/W0R/Ko9mC
bPPlqpCjnUtTvYkAhdFlHxHT4MiMYcfP0c9ArlcMkJAnKZJTKHwddYsa2ZjHfKLh
d5x/H+4vwK5JBIITo2D838fVt+ujGf3XWOXgoPaDcaGK+O+kcBekGOh5WdUsmsh4
MOlmrb3Tz9Xt8IQgA6cVlFBJndGEvsaomfudTDmuHoz6jYJBiNcxqGDzChu9QdIr
CnIdwrMu32dr7ofs10mtnq67pc/Sk9fs1cMpBGyZ/PwnKJj4TTcrfGKnajZSwekF
R4GyYOx3yhHe3B8Lj7SAjnfeTmGbUMI3BBvahlZ6YcLokmJDqNCv3B42TI78SD6v
QEuEkPrAOq/wHi/PGq1l8P51OuYUnzLT0WU//t2zXngU0Il9r7G5IS3WEi7Ox8oj
`protect END_PROTECTED
