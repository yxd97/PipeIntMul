`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U7wPnxNmZhUhH1H+jvfzYOfF5EfBrntgxUMxXeTvS0halsHbjHkjiNvPkKUy8IQI
56wy7i7eFFj9K4s9t08LXuKLHV3GPONdH7hUGZkqSx6XVjlc9nW9MjoHqJt4BPoX
w9kb6/JJqyyiKvlcm70PfNI4q9BLMhn/WDGKcUM8z7vVqk7WkRZwVEiZQjQ+ql1M
0aKVp1W7MxbM9jt/H6JYpOaxIzhKjDW3Vyecw8xfEIacuSj4FdJ/N2Aziip4u29K
Qskkisyt9OO4BZL+zVWwmWPsZnCZpAJ522Yyc2kmbLo=
`protect END_PROTECTED
