`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fNf+hp9e4JmKv8QGvs+7pn4cPJIGjgZ7fhV/EbONRQ6IySSK52lvMJiw1u5aZCP6
Cv21MraIGfSmpNHimjs+7h7Px6ODCw7gwyZvIjYluwEVioB9m56foJlfTfPTGuJ5
O9faa2bygle3rQlDRkB++DYCmPUKTiuwvVwOTQU5253vlYomFb6WKxKmCd/xz+eP
GrNelW/QVfCmGhADlq+uxlh52Cp4GkYYQoAONYW1Iegcu+enRI018FpLzU2vBR/6
7pCEhxnw6Es/YTjSXLZzXVUHncgjbdSjljefPFH3NhFk2Zrv6nWoztZJZosDtsf4
W8Q5i1aqn1LWGjGLb91CRYvUJT9NqLCHZg1H+uQ9GdlN6FJYfFQ1ZZeuOpk3H1Em
KUz5ydCNzgIvh0r9/Cd9e85tnybi4ETQKNJM4f7bVpfTRuMNr/z6jlUMcTB5WseF
Jkp3HTFQxBy36DCeVDtiBgsrvekKwMqdWk3n0RRc3hJEAn1KRrIW3deJcFsj9t85
PxtfMJ+Jnb+6zw1pyY4Vdg==
`protect END_PROTECTED
