`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eehkw15FMrT3dhoJUDzpldoOfGZkSgFA1bzHSnpSRGaXyZZdFw+1utbW6/aXY+6+
4jI6h6slfr9l2k9Y0y1ITEhalWg27Bssv4y7d/vbefIipQEZxAckcJyH+dUzTKzb
rtx5tyBSj+wGnmiGGVzAkd6NMVPq5U74TH9v3qerA7E5g81exoHknXiU16ZhSvJd
FittO9jtr1V9+d8W9ota5CVSwGbfhgxH6UqRYyZWCVV2LVSQn7XKPWeOhpt2Snpg
QDbFD3SD5lCrQP7AIyBb29kK9vBSUdJO/b0rCWCtx8EbZVdt5O14PR9p8eHGFUjp
3ZiI7Ii5923g/Osp0vVJym4G84I9NCPqjjUIOFBddpPdIxJkqv5jl6o3nQUMF9tj
UNlzlYN42kE+fNi6S+DJZIMCzEv5mF7YFEFkru03zj0bKlixW+UcSeOG8t1tg2yP
nxhMZTldhm6N37kLAxJMzu0Op1FkBAuYZjX9VkKXlJwXfNwSWNs7b6FMkt3D22GL
ITl8VxUyaZ2jzwiS6+WitO9JBLk80tMlyt3YBcAhvBiJ4SkjOkPgyjl4xrnx/msj
MMB6JW0A6LSmY31hLmM+WM8tu0hhZZ8pH4munOu4akCGdNnIPKfKbZdjUO+qRD3p
ZtBiEW0FgWEXLO1FSrOMs0QYm8QcTgpr4x5r4PQhTu+tPo8vOiiwcFubO1fmH7XT
HqyhO3celAIUKPZ+Ld0QYqMQ/U+O/6PqYTvI3bYpgIP/AKKLav2JKxJvvQqznIEC
q+6yti8V4wZGR5ezUdOSCD9wRLHuD9bpDJyS/IobJpPJNTl/Aw2iLq88zL6H0iYy
cIl3/OP+Uz2PS6A375NktjudydVtJPRaE6BznD27AK/b3cUMuclkPyxufGmLVeYe
olzCr3iuiRrv4a6TmSoHWIQsXNjRzGr26hYR1t6D89WTp0GUBTW9x1VAhOLj9wYL
/i1g9ORKmXkSK5mZW7A/DtG0TW8CA8WJHBTlERKZCUqTEQdOvticJpUQnqIQVRmi
0lPzg52bNr8tdEEkJP1cqgjXUH2th0G5k4JX4ik8gf1gsQmUsZxvnxFDsml2krBZ
hA2MJoBwVU/b30+EEO08d1QoqYS2Hc31MnaRpOiTDicHHGoHCh+L6V2vO53eGzyO
uzM/gQdyV+Px3SR/PvJ9zYCk6iBgRg+V9pzZSwIeEKy0KZi9263WCnCRBDJ1XfoJ
1evKKkc++YneWbXH4sEDXuFPLQy7SXtTr0eXXEzu+RIOFyJqVTOn3NdU6kse8HnX
p0TVJy26R6TnKUFJgXzpPmUVnvh8yuMSRXFIdHVbWhMHUPFcIZ1rNA2lcvUt2bH2
tDuIy11XTrO8EoGh1klyTZT6c01BIIifo3nOQueFk934D8/vKJEzCe+zk5oEKVaS
+g7QgSE5pzkItW4jeMimWHlZkxo+pPBgwr9EzjNKYOoY71wOpb+JWgCRd3/zlyRZ
2mifC+grEhpc0p5grAUfCKqpKg5P+03iBEmxt0VSYSgGMBrN7Z2UGa2G2uWo3paC
h/d3++ljcWNqVH6tKZSrcH0Ycrg3dJR5UnVEunF72p8B3ibZEYeeLohkuWFcwn91
UtY0G3nnf0XmPi99U261Px/XNqUXIWw3leJMx8zFLkNmhYg2qsrclcyk3v0pM+I9
tEyPgH+lywDITd20HpGWww==
`protect END_PROTECTED
