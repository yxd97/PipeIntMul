`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SxD+hL/4MvFkKNiC3hbAamuDAPvp4asbYCAQSay6iG5R0iPJ3eiOOkYj/q2u9DMn
HvPzKBWn7go3GZY4TZ+RlP6aHj7lXbB7hBB+QS0b5zh/w6ZrDoeJwA3rLR4huI/m
QTcJhL73HVMKDW9g5heURp20ojF468RJriEVzXKXX0VBrd4/VljOl38GWt4+5Zzt
l2S4LECSbMGKPw2eb1Udy1L4ZBx9/0FrmKuAGuEnL3RRaPhWOm6VEOHORseeH0K1
7WjWMvWFdArv0ci28rae6l0ra/Y49bgJK35LzFKDvtMMgU1DwhVHgE66hbwMmSZm
HhhtJjI1BgPlI4ohB5yDVp/rCIZTPEYWoUWm7aornJiBB8y/ne+6zQwBJhv9/eB1
UdtQDQ90vWQid8+IDI7ykhn+6n5onukVHNZqIgCTajA=
`protect END_PROTECTED
