`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xvYVTL8KoGjxo7ziAajfYZ2EUbPmh25jnPlBc/T7tJ4yex5lZVy+fJi3MjCZmQDq
rbgkM3K2999JuQb++Ksj6XPiH0s+oD2Be53XqC7OyBWJkHeEX++o9dlas+pBrloO
NvpNAGEC1KiIStawTC2JiP/cguMXBvP2891v4jVdk26PG31RZrgB0o8Fq/ZSoXzP
bF0x4N4KwyYLYD5BZTyY+Nefv4F3aKEU/jg0l54dyAulPwIAcAkTjWAiWJGi3Icl
xuYVA+LbMldOUcdDibDSr1C2nABrzUjtjBMAOoht9N4EEpTPB5K7vLOgsFzgzaC0
tbAYueLJ5d+wFq8GvFgOVP9qXp/vzUUQUTK44cvkW0wq8byRiDR0Ple5tEWFaH0t
vz1n2G50GQJ1mgwTXkfRqBQ8fUnF4bEwQeWLQbVnD7WwFEWFdu/Ke8XsaIyhiMVk
`protect END_PROTECTED
