`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZE0H6za/Y504TmnbNyi/bZt+ZqfuTH+0Exb25R9ThanAe7Or7JsXFHoX3++BiMNQ
R/Ef4s8EqX0ieYF36meWubXR0TOIC4s0/WObBo77bx6VFK6GML+Mc31eFAmzJFfw
C0GHZJzXEdaTFZjsYs+2sh5DeJqtfWmSQ5jMG9iy7g/M/h54U8+3L6vuzLoSu5qy
n1cbCbR8kSJFjMZnuS05nfZPV6jEgObs9CpowjlwV/+hKA5+BDdf7UuT1++HFSI0
Wt/bWzoWillrPk6oYNS1EriW7PJfOsFaARez0+yG3IvcHIuemXuAeMKZUUUjoQTL
SpER9shWQTwbq8ft3EGKM0HupGtC+ekwtJJY4+VPbqjcANmmpc2IZ2PqLwsW/euN
bbJdPuGukpMSplnCf/4WAZMaXpvlqxPHFdWoS/xLQI7QbtILwJdiNacIgW7y4NPd
kAuxqztvwsDWom15P5kAsBJOBdA3AEYdtLFboBl7zUIr7QdB9N+d8SE0YCPvNX35
xhWpG5PH4UUIiDJnNc3rVJDsKptZ+8nMFcKOzyyXXNw28fxhzJZLd5/6OJbLnMTU
dGLYTY2ojbwJRdQCeF6WsyXQ07vIzGeleImaUV3FMAc=
`protect END_PROTECTED
