`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nerMp/CuaBtdGRCjf+SaqmBXJejGzWbhrLk146OL7MNzlNbh4zZWewXerzr8yz95
uIiIzKLD5FYnNyWYRQTcQ7YIk4mRc/02Fjw396/Hqwx7Z8wLAbaFrjltmCBmUbrX
dPd6+4NaEwxnoE6OmhdMmXKJzE09dSS61HCGsevLXxbuVGLdzz0FnjoB5gCBLoTT
H8qirRDCR+vf8ALjEW3WaAU56BMawJORNGt+RLvKTTgETL6M40BDN9xGIEdY2fK7
X37D7zvyF05Same1jOLtRzyRmxi4b2dtA3ujfdAtJS3P+e8s4hH0vW9rLfhrF+8U
521DccgUCLI6pqCd3V4RN14HSeBHq7uEioHvda9eQqoGeCU/ZfJra7sj/ZPO5KYz
FNGR5L0WcbDgke20r21/ZJMGJOB2W7xlDQDmHthr2oW8q5ygmaGQqGVGPpNejTtQ
il2TR6qfJJgEp5eDZE+hZQaILUpLqBD0odBjBLIr1Mpwo/0kes+mKvbh8FE+pyGt
Fsc1HSvJNApTucHHoRVqqboW08LKRKr2dRydX+oUeAGryvgcAYCyDr7yMg2y91eW
vfu7AeZnyghsr2cHD7NLZoFt7G6BIerWQxolUmHswGSK2NeCaIoZRLw8DuXrZAGU
FajLuTZ4yOlKUw+uUag2iNhDClCgK1ZI3hbxmc7WCTBT3OL/OB9YAXiNzjqaEbxp
mst0Fgk/XMvw5FeVjDYee9XQPWnGgxKvJfFo1v/HBNKT/d7VRblKZU7A1bG9FGky
41SeY2DLzrF0yEAJnB6z+jwM93It2UAUosf4+1HUemD/DkvYg2Xpb2m0WQWZ8BOW
VcH96GlIsEtkUXYFMCCFvlkwKKOpVBUEgUKUe5Y9XJLmrPxLtr9SRjpUaWp4bZ9J
Z2QJc31LTgIXmztSBKeFnrglV14PUticu6nSpL+a57c9zyOzfOalmicroev9Wy4n
PTK9/0Y29+uxTMTblBrD6WRU9fD5mZi8LnLNz46wEfXhTajewD0YHNsvWvWanvxv
`protect END_PROTECTED
