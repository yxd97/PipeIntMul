`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUpahkfQwGUT0bmFeok76+mX7n1M2zaghi4xYihsgxsSuj7lHN5Lqes74G14MjbU
svdMy4iXTbWJb/ioEc2XycQRth35sNGiS8gRkOx/ageifclQjqqFbH6/Sl70nZrt
fFCITI0OQBt1O/28GYYuaLAxUTgjoQUmAxPJajvHbyHTlQCnJ7X2bmkeZr7b+drd
AM1uujtCdC7EbrkYi/ISjaGz25unihwfdQmvWxwDujI1vcIOhVSVNNcWXPQw1q+E
C6tukUXDUfqzxhEw/kmArG0U3VykBq3bU53jAVLn5kJxFEHT1iKShN9kWXFQN1GN
SsI32uTbVyLyNou/VNET9H3yb+okhvM771n7IlUUYgr94G9skcK3xDNfRTrhl/x7
zw1fUQx1MXTrHDqrkLLCD7DGlwQYKRGyhhy5sxp4QSUQ1Sqs6myhmn9uOUXN7vjG
m+LvhgWTJWREQ0TAXIAe4gyi4trm3iopOuOF8Rub4GA=
`protect END_PROTECTED
