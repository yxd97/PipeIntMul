`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0OAeotYCd03xWx3wk8RQfk6VeNdLDU+MnvZDZhQ5TgUa2MnlkFF6z+1U7XUj7/G+
5Ju0yofXdRnu8dDF6tglT5fTzujI/y6AOthgAXXbnIfbXqrB/WYn7YXmWJX/4+L7
1b+thImrL7K4s5NaA5vShhBvzQ5rlSZPVYAbKVsG3L5DjOgEwNY3B3nc0XL9cFym
TQt32qXpAUgZCAlSvlVZUtcXRoYsJ45Nzuck3+KYk+/wQh7UVQucPduu6LcBMZPL
bfYmysIRQ6a3QmAwihuf/vAcCnAj3dSmhp89J9844nMOGxt8BIKGkqDJ/0+B9GLe
i+4xq4zJxFQ5iY17XKZxFxp6opJm47F2GdyqautNmRGU+USqTKZK1V2NTXtUCfH4
89CR8NsdGXOE3dQpK59SbCpjBN30MZJVPMHX8ntKWbeGoyEg+z4iPwAeTpoHmOOl
UiSE0GihPlsY9Qwiz+xWxKS2OvqsbHJpFtL/8JkiHdXeUaEg19Cdu8/LCbKKL8Pc
BeEYmDml9FXnuR+sZswM6MXKlk8u20c0M/klEPf1YnfBndm7dLF33Xndx4QxqIxT
vJfmbPqNdjETc7/LU7VK2ZFawCv3EZ6LMuA3hnDQcXC/5ozaFl3vClYAQ6bZzqpo
CqJw+iAV7ws4y3lpx0oBM5GnuXXGVYugGB2PbQkIl1rdNmlgCHUmuaOu24Ro6DOz
KxlcWUFfLSI8I1VCWofuWDQx+aRP7DdBaU0ytba2r6Vq1o/e5Eo6rugyY2D4CQNC
UVkENgmkMmvfHyHAqxRAYHQyLllDabh8O/K0exJZP/hj6kfMKNigbQeUTcOmF2tm
drCk5KcYW+FsCSgtkMnkizpfSTLcQTQ2EtHnxkfuTtwtn7CSkXzMZZ6VMsRQJidO
OXCCROoddkp2hgnXAf+a1E5toV/BiLkt4hvjfcW5ZGtcps+/hPhbuH40EZitIGyS
xww0+Y7vHPNWkY15BtOKKeCFN3OoGrRxZ1nZsW2snY7QkkKbrv4tKur1LTT/6BV4
slU5qlPN0JT5jvPlNxMLSZhejSZrEZeGae+heHUr3B3pOzNC5l5QO1wVUhmc3b1l
GSlKAVO0kjqVMVhXBwTN6KtWkbVnECMvRR+zuUIAGFAnPnLemG5gxnBKzKyQ4L5k
epoIaNUzq7X84FuGgIFoGiwhr8CFF8yzfNWt9G/vGBxws5Znm1Oxe+TLWFK8qijj
1Utef064QWjMXGkOlNUG4OzgzHpIJEA96l41mBLdnSmm8Ml03qRlpJTb/DsbFfjm
NbCyZiQvb7aflk1yNKZA/QKPOm1Ht5qQqrs3m/Mo8x8WS+r8vdAjAS9vPBKtz9Mo
m7T1BM7sf/xZlfGONa+Lc7Or4NTTmC/bBjW6rj/Tjird4H2gKItO1ez0GYJJnfE4
xffo8JZqWpsEcr51LFWe0NXYY7B7sOGkSbZyAnbzL6CbpITzIXc8fn42xLcqanZM
F8AbDhlrCyObnjeLIdxXiqe6GVE0m3tU0XMw5Klpd30X0CIqAsNV7wUYjw2MZ71G
Pr0LqQEaNX5qOUWaPRtLFvwxuYScBgSXbXNddxUc03F0BA+VKK/9g+6/ALLDU8l7
0f7lpHDPfGNX/9AX2KMrUpZRIAVJRj5qEjbKIWnVF0seuGiKbEiGlCpPteI0Lrbk
uG43/u7Tp73wmx9tPCzJqVhqc38FduIH8RA8dnif8rBbdTetsMjgt0O74gqn+kyT
A8vJOLp2tRNpViJe+4J5hoYfBYqHohruYa1CGtymtR+0R/rn4nuanUY5ZircOvDG
ffCPoCn96aabLT+vrErYruuCv817LxHMcNkJDErkNYgARbXv2hV2kzWEbDeIhBr+
hMu8wFq/746830MDAzCFexWX2fBqMNUsdGF1IeR+w6QSD+RzxDPMmIhVSV4Q3zZc
dWLOuy17jMqMpWd0DOCeBQN6tYjWoBlFx5s7yoaHfQJzKAzGXK2KKiolLsgXNs7T
Qx4ItG7iWQLWz1B4eo4OpL/Ju48eXvY5NGLnlQXE68Ve7IT1v1fQ40a2jAsQNlZ/
1rKu2FdN/iqkoNFbsHOTkAlLluzSRW1Cw2x+GGrJYtu7uonUItfuxDjp+9OYH69l
9ZslIli7LHzvEZQ3vKW9gZUXcwh8brfu5mzTsiRfoWAc/1O/lS3SVAbelJcnsqIc
kiFcLZ7W3y67QiIcTxZxKLG5Swsr4d7N4lHzhqQJDdkcinFgC9tquQ2FlfqZZznD
`protect END_PROTECTED
