`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZA8Foh5/OpM0Wz7Wss3WPxWc1PGDQPzgiODRjh0vJZ0b5OK0vtDTFNIDGyiwhQhJ
UdbOTxla2Sc0pW1HoZjGz/gS5mh2X6O4eEs+HEEn4TyVs4ueah/w82W+jSqX9PnO
by2VRt7K2nwuJ81PaVqaDxuAvmgAnF2B84yzGXh6g0zvV+zyUXA7slXR9tRsLMQi
qD9932BIVqclcgTfal0bv/KCMDjZpBYDaRXX7ID3vRb3dEg8ufuaCXxdl3Vh0x4v
jKeYQYEtG5IQy3AX7eiwicejqkcMTKsdU/f2wJn6C6ONMyQwDUMrboNMikqdgnCj
kuiUwFutqb6usGYoL8ZHhUWDGjQhUZ5cGIDfXpe/9q9AaizvM99yNi4LhGcq5fX/
GYhs/EfG93wSedlwxZKJIA==
`protect END_PROTECTED
