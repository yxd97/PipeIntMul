`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cXUkYurwbwazyXQ4PwIfoVHQi+x+6ZrLsdJy6G0L47C8N/cJjX++HP3mplxOj8KM
rovd1xlJAdUF6HTXj9/zIJTHDYC1NUlqCczruaoR3XBBw5ua26kWs95OKjfXy8Lt
U+duO50CLvxdyOG31XZVZ6ilzUBQOsuqPM7K0nQMiIaV/E+gXYuuq2Khu8NNRH28
g/XXbqFl1wliFAo2CNp4FkhaGZipkogtCD1YE1B9KDCIFtzbyEDyAyHJwxup/Gqb
bdwEe4D0oBoxuKgDgIB5Qiq0f1TBcPDBwXrgL2J7fZJmON7FHeCeVAkg0js5NPNE
6MGHbGF3y+QCTIX2UQUReizv48ebGfaV8jL8ecUAYwGjLTAlcC7pBQxFTGON45Xj
0p8YVBY4BUihmtAvdiT68PrP3OVITWxjK1B5QdpMpaWCvobFoXPR5+ZSOkvGzy4B
ulEVoSUJ8LHa5rkC0ZXpqa+BypRlGYYjuw+N3R8Inmdj1i9dm1xZdprbgGjUAqtk
7iP2fshGF0Kyse8lmxSAxtj+Q+tfPwJw63Mx5N7bxMjcyfBlrE2GBY9ql32w43ov
jCPhWKlW7pZ9Ckzl4OEJ1R1NDA4Gzg6S/kmOIopUzSorgDiXmuMuetdEsapcxAzX
OLkGtzipYA7qNWYa06uy1/n3Ztv9Izkxkfl/uV2kZ9v9yG4RzMFQTq5BB1T/T4I5
mmGsly5GNkzK6mtQjN5f1Rx3vXnE3EI0he6TP8BersVLcybXbFVP69+PCyr0wf0X
xUvgYmEP7lSQUgEZQZVK0O1Zo//EJiE0aE9dTyS2noeze7IvRPcV0AB+cVo9aDg3
QVqEQXqKtFlUroBkWJLUY9DoUAzzlj/q39RgtVU44dz/3hNYKrqkjtb5I7+KE5XH
XiUvVTW0l4A3CfUfz5EQCjsTu0dHpC7CNMtXC5lCGiMxqWas9xF4mtqV2ckYIfPS
8quJw0S2r7t9+jvLR9U0gOtV/gd61YIlMIe+oVW45TuIoZS5ouUFVk7AlqXwpBFl
Bine9pWXcVHAdp5c+ak6V3FC9FPq9yZZkEwHKCX6ur2Cvs3NfjAkRqAZLYhUdRE8
`protect END_PROTECTED
