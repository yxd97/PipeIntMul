`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kMUtwPx8AUbBCTUNAVrtjYIW333hcKBfUxkEyyrIMRkKFROuzfhbY28+oRFlLud
jzyeRqFkJj2dL8LXP4TZpYIbBL8Xe7Gs9cjVb38k4TWFTcslkCSKp5QB+XFv+Qlq
pg5Nj76zKSEA6MojJApz8l31HuhrTr7XWRKlC6qMrWe3GIDJO9NVVyIdD1ThKyoU
hq4eZ4bK/kMoPY2MRF+joDR82wuPix+bPRki/8NQxFGjqBq/xKfkPChwgsGKD+YL
vk0rM8zxjTQrqlp8ZydUCwXVTyEbAAE7ExqKeEyCmMb58OjVMXlNlXRXk8J/NOIY
mNPhPcp0Qa0YTgv0PI/eTOd8npEsUYSkMv48/W1NLuM+Jf8y5JF8L10Ma0YGjGR2
DZWTlPZyFHTn0fZXnKsXcg==
`protect END_PROTECTED
