`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZu7UMYmK7BJgmnSHuSr2NTTxYBLAtzxFbR2QO4q5veTdnYaMuHcbOZrn7kL5Mdx
vySaoB/M9JaqodqyIVEXRnS6jfELcW2kgTeqV3HcfWGxNSqy8Tee06YyUUoeo/ho
QhFN89CUNlVAHpVGbF3c2vPc2HYDxKIqUn5obURCkFdKhV2FpEgoeQqjvRa62Z8T
FIsLgJ6B26MJ8U1IEgcZIc+u6pasriILo+88aQSQJhInhrArV09cpbttRfx9/tbb
VW//WMoPOOOqnxrG313tbhzEboaLa3t4ZnFV0VE9q3xTf6OOpRt+zijMDLRppfCU
Y7EqVwuicf7jQVTMJC4m7ZGgJFxe8TGwYHHgOetieoyXSIuWn4TOMb6m8VKVdmU1
VQnVtqdHv1wuxwKgx5Lu5TCTTqWhW9a2kIppWZPgs1XExeLRGMR9GJMkERPW3RcQ
1m5aS+3+rsIlSQyQ/X2Cy56cNiMi98uYnAkMfesABUErVtSy2VCrGg3P5WdbuskK
AlSS5ZFYFQr6EvZss4kW6fFbvKOIxjeZMdljOp/r2XCeHuC9rd5v+z+vvbizyjqi
k5VCmobRmHejkSqJedlD4XbdD8AvbPyJRkbExlFNFvrSxvVQmgdmOj77uhbrVRF/
4XAif4VWWndbKxTLb/75AM5dZTQkn9aBic/4lvJ/jgch2wOHB7Eprh8/jnafloF9
dQ652abT7tDorIL4/XedYi9thPtMxcJx1zUfu4f+alpCB0A5z6Jkj8pJs6QXdinF
pPzX6cyq2ywj97TYTQvXqbERP+ET9/Z88KTvXbZuAMpDw8P9nrUSicoHvLFIag21
TBuhaDihtxXodSkKjAqKhRfOVmgT+OzKJBJqVnGO4g7R1wWnJzDeyCekWTTdRQn5
NqhFR1Xo5kIQs7GViBBIDLCcFEtAZGBU4Z/cpFCGR5Al42rDbdYLXIaKmO7LPnHx
0t3z+l5LNA1WXa5oPlrLbvZvJyDSIDEsfeEC/3cSngSYnrkLoqTbhFImKmRrK7Aa
JJLW1nLaYBGYdEK9QMr3nwDEIr8uigG5qG5LhM5OnPrZFCjO1Ovc3x2SmtTxxlnk
71iMrln6K2bQnuQ0OaDXRpITOt1q5W4Di/QN/l6mZVvdJOB3Pw6oygFbDlGUswPC
slJORYpXku2+CI3Lc9fOiQEZiLKksYurN8n1MBV2dj9JNgfYXHHlR3BAi8DllK0v
0tFJfzu3h0R82eff6gY4kJD8hcM9T+1FKz0gusxwItBy/Ko+JsW8d1uy9B+K27ma
ze8kVlnH2Sr/7iuW91IWgbdQRC6phA44NxLW0DF0aOF9CMlc3M5nF+SnKCg8NLua
uuvgMEG8kB3BK+AA+FGrmiYRBPzcpA80ai0pxVSo6bpNaqaTNA8ibsNaKqXN5TPK
kL1Rn6tXUAaZOc+At1PifFyV8UMMomEQ9bLNwsVMpdU9shX9cL6gmrAxJEqxm0eS
h3N4Ikr0HW8aFyExyHj5MbTrUipEMmbk1r9glp42M6RTJPr0boXaswAqpfP/4J32
WCPKwedHv4QTsVtJIoqMUDyIMpi5lToRwEDdJUlKaGM7P6jaACqTlQ7x0sq2k9aZ
B1oSVM6TJGBrMYaU7WdZ4uQQWmf88PJ/bHOHPoXwFzdyF+bCGKYQyr9q9W/D37+H
XCWDe6MGhSHM1zdwoIvasg==
`protect END_PROTECTED
