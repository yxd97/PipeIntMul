`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PU8K5Ez5FDx2N9PDQH6z/jt7kAkHdqJ9dnVsyWtgLfgzFJmXRC59364tQtyJJUQl
sTyb05hKhMcUQk4rNIiRNh1Xpq/1FguTY/XDYPKY/9BjdvoMnAwFMPP/+nOyeSRE
6ag1D4l6UBQ3urCw9E2sATFNnzaFdq6WXEmlqhv4QCSV1kkZ3QVTLWqNNOCVLNur
EAMMV8RP3FFMhspdrGZasy9EA/DXo2aOV6/Hnobllz3vi1c1hZdpxyjtlLNnFXBN
sUWInlbQCdA/5AnwXUBGKuKBc3H8lCX8AgBW3VINxYWbsMx2842+5ymY0AsJfozt
9MVjT0hSrCidCJVmd0f3h0C8YBvndyMnaDn6TrHdYE4Lfj6IjOnvPN7Uz6MHbYKo
nwRAaVUG1eoanvHWE/B+S6l7yL21btlon5EauPKUKMnwQz20jLL4IaWXWA5wj2DE
D0IldrAN9MsRaWoyQjmvIgMrjuScVKztpK6+95uzTiJG3EEjqDSnec5gdiT6LPOa
XsCogMgfAW3CPG6F1lwQLoT3AMRsz6x2qf118JYAESayRnDUh5gtcOrrhf0JbI8f
Z6p1hLHZSK7gGzTxMEb3mlvubfFIewpyXnN7cRLnkeKvVa7yX3QjdY577tzGr9bP
3R57L35q0IB9qbGc+9SJr3CCl5U7D79yWyStnMNX5j7XKIKlNTr+ybXC/9lLGvgy
Mwi+nj4ABkWSJEhGHEzxYQ==
`protect END_PROTECTED
