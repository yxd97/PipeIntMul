`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QsAPK57XbJlfcs2KWJFcidebsjgi1P+juQrYwO+deKtjDYpXVr928u2fERYplWzg
SU53VQa+wzjOtWa8UPcgFzqbL34YJ95Scwrlelrq8Oq4lag1Zs7LaZkQgAtepdOY
SXVxpeSFjMzBYxkolvrIOG97MCxhOJxk9aT4Q22bQPHXGfWGLcdFdkS0P/m/kqpU
RasxDtNKfRXiFTA4/P55uzKPV/qKRO81dI/WPYGFLqnu+mR7Zl/R7/oDcD0+RdH8
f2526w64rkiAXyUxWNdje47b3cJSqDUFXEU6iKQvhWSqa3XoY9QYbsk+5kyg6Os5
suiOJTjwcY8lC1dO/NVPja14UEfPmC2uOFvRKlVksGGrGjMJR8scdS/HQJQZP4rx
i9Vpj9ZjSWqzd0vxsNdb+i0MRCmvwT7QhPbFO7dNLYE95hCBCUVIfd4sVIenPzzg
4Lp5wHdxXxmUVgVdkS741GBWEGSy+mQgQ3SwiWtTanUqgd7Hgxmhptyf5MikQ1+D
mYGHKE6vvG069w9kvWTwkj8t6guU2vZdAieKZQcPXKYTdV7I3S9WaFRpzJVzzPiA
VOJvOXkYXWyp86GGymqZ7l/2dZIsFAhCvCEckw4EdvA4fF9OdCBJFFcEeaTELcJv
M5nWMKisYjO7ducU1duWaFSwY76avDg70pqRK3cro2mqvAwmutN0rLd1YUJ7kbHD
JdzYCmSG9qx810GD4476tVJzGnbYoJn7sttlJ0FUgbN9qT7eyTIw8Ru7f/Owai4I
tCou0nJaA/9AeZx1D0y9M/ZxC19RYHAFWJXutXAIq12J+vwUyJx2DcH/fx4z/awE
Osc+AQGNUAHa02FGn4WQLZbhLyjFVl4xapbVWrR1/hgS+MwzG8HNa8dp1LhPi1YW
ZDyIK2XHjqbQQMJbAp57rAiMl7RgU1fRt5ydqXvczBHVAzUVtlVT5elK8eilGwhG
eIAkvMrnBmVP83xrBDorEQ==
`protect END_PROTECTED
