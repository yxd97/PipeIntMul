`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3sQM3vaQIdLuMBNuTmwnFnB/Vpqw5CQ+BI1U24Xa85LEkCeUAq+EBq9qlSS+X6yx
de9AIvQhRJz8MIt2kgHzATo36YTqCxk7ORuv0xKiQHCGhGlhHrhvLtyelzQD889a
nJjOExGhHuHr+qa92mRw8HWvHgQoQ5rnhVtXHdwuxv7U0RNM2XWWNa4qlrS3fcHk
r8mty4k57+LqUPYGJgXHpKfgHZWptA3E04nptIXVUEmkWHakpbsMl96Y3JlKwfhB
lag+9bzZ57mK3yOFL6FEScDwkTIVyyOpjveP3pco/Tzs8kKCa0wtcseVGHPut2FH
VWhY2lKwGU8O9RkStOq3s9mA86A0z16xrSIQsEqASjKwAWVpaLTFyrxJPt4F7jYL
tV1L6a8lndBrfPrYWMDceTMkpYAOPDA1784TuPkNpMAwTGGolSJiV/sAXrAS63qe
2WdGrcqFqXS2JKWPtgbZOm0CK7+idoWa0yAu/rys4IetKcl3DegCC9c1dqQW4x3h
aKSQ2f8SmkTb4KOB0jRtyYu2OzzfVfbddQLj5EwPfotb/TEFlL071AkCUrOVSx0D
o/D3LT7zwSqpdzBIaSR4C5yZiuwDl22uo+MqcSHcleuLuDjSEiq2lC+6+w3UMPOs
05B8afSKvZY3UCwEFDcE9FRuWsirRZPpV3LVkgFqgxm6O0R73s7poKroOjVMseSQ
H5hZdlyHtEi88j9iEMT2XHAef86/e60jjh8yijvOLEHc28A4yr6/2TW8i1tG47xW
+1d1ZGSgiv6klPijr6rlifFT3XkK1KbQF2bnjJrLGEEbuyul1oz01PoMF2b5iDBQ
MjkfMLBr9vYaBe0bPejTB8amJ1fGN2oxun2G+cN875J34ulpkg/3VX/qm87D5OMp
PySnJydrjg4fhMSKSZULfFgxU0qF4jepWjsjhTYIDjz+by/3I+7GKpsWKGtYfD9Q
8eL/R5KHpkWgg3qCGNRHp6R5hJhS5tcGbizk7xQE/PWYAdjDe+N9hrtrtXbwoOsw
Lvrs9w/TfdVmZx7UtfR4jOPcQnqWeUR/Z68YiTWBuz9/1+qeEi9iQQ1aIryGKe0b
L/trV1RgGaFz6YzjeK8sI9Sw2Wojt+4KD0+ihV8LiAYMTke4qPRW6JDASKqSZ6mq
fzigen4DyQ/VsZ8doDsy9ruW1GwvAHjouY1qyRLI5fwvoz4OG47aLaHe791KKmL5
SLYkTKEy4wUv1MIv+J8oXRDiaZQPbcm0b93tY2EO165UMlotk8prkJ5GtPuS+GIS
J4CVdQ5pnAWc5c9OZpJ2dAh38LF25bK+nhm/LRyC5EZYDPcgc3GVGjvzXNatWkLr
aR6PiqVnolpG9xthDsSKeTBEfJYREWz20Nd27Ke002hVt9s+AH02W3p8qfVQTl1X
6J7c9iLQLNCML0r3oGu2iJwomzgDT2v3NISF3YEd5lJlxZaQ7xa9N2NyIh6ukRJw
AR9T9bXkkMx+U5FZlvbWuPuV/rn0x7hRg4wpOY7lHO6AJ8NKSmrNaod4YBl9npPf
b8QDHF+oXrRvyRu/jPuDGkXsxWPGUKmkB6CqqJzydgkHzWuEuDaaXp7658H6hTjY
edEWT8WDIUTpck/gcnTKiH4uHm8+2fcAtQ1uiGIImpsnF8NO4vBERW4hhGQkDNFE
8t36G5WvgJ1Dh+DMOgDdP4Y1U4crHnbwhD5AcAQFMO7FRig0ArtnyYRj9kP++l7p
uE4FtKzNXFlFCfU0ra2B9Bzs/+duX2cYjKw/QL1H9quuVu/9+ypgJketRbiBwVJx
GcvEMrjKPg7WQfK4R2bwdwlL+gfYJhWVZhFDRXhjd3PpziBt0S6Sa92go0v9FdqN
MdBitxDS9Uw1IlaUiZ+v09pl/M6jNtHbKMkLGfz4AdZVlRXz7yEKHamm/Ot5WGuw
gZX0SrEM80379LmSAVGddyHxMRSPd1rZVU4JAzi+gDh9sZl5c4cgJNwCnL+yayOq
Ny+D4lA8U7SaO15iU7hAwgteaSb6UXZevh7oAPKZafy7GAe4k9PdnLo3UZzJ7yt4
ekSpj42Wgd53VmRG02sUZRo5BveqwXi9rAYfmT2g2eNMU7UdRLUXAsEWqfvk30dd
Z0Ixbu12ZQSBH42pvk9tbGoMFYKPCz1jJTD/rfsNEGdg2CbRf9ViGGqGR3GBrmgC
8/YTUEXzu8o/sL2MJrPfIl/tCdznDC7DXHQ983jp+U4/4JZnFnSVO+Q6fUcuD28j
TqlQ6GXbua6Gf+7C7odHpNEKLR283OEHJ5rD4PK2tP0lnSW+yX01t0gTOeLMKnIo
j/Qr9HWewSlWKFEHueav8t+/ifZaWKxMikIJUquIZ1NfQq06MT9f0KaUDLK1SZQW
GWVEgwJc96Q0az+28X+WfGTVW+CLPI2UUDNpyKIy1ohU/zHdjnA58JPqEKH2599c
aSk2K4IQbMNl3QwhilvWZkcY7qa+87CIfZE9RClflrd4gUHwEnIxWmkMm7VgAKrx
6NuXRegpHSbJyGhO/HDHUHV4kAUgFCyrXv+SE5e3BT+87oQPi8nZ+fnYt7GnJEWJ
7K8otn4xtW+U5JDYz1DE7Gjx+WbtkBKJo6AoA6s5mDQJP2fBQ3MYrta5CDdyjgH4
eHFpeVPJw8ethsvb3Zh5hHz/ftnZ5w3V+dX1DXRZmk59WGce7uguVKGX9oeh/xaw
A0ChD4r9hK9nS9ntGvGMTs2x4QByPJDkZPibXosvz20DpSyElrr0bJXjbO/SlMfS
3r+/aUN39pB2jSwHc+FxdO5v/CmmBsIYBTtJLe3CjXVU2JhTGxJg7EQQ79f95YJM
AuBChX6UFBdUimOkvpilF5OQV3lL4zwkkn/Jx7va/W+TJvObPBn1LYJhM7G2DH1R
rNTOsArB89PVT+QwNbjPJaST3XpdUfzAgtSuuYCjmcWVD5OYUyNaW/OkhLqRElTk
Jc5PQDTVtRU8H+Ao2U+Y7lJQ5HdTqj6FHOu3EtXujFzJSy75YW/QgCNbAc4960PX
CGcVrmoqPxL62vrJtppdyBRkNYByDA6FSy0HO0HMMlvIsykAX9o3fSbSJVvtECG5
qQ4acf4BHS/64H9GnnwqIearg8mOMXrbZ9cYqwsHOt2+QicnYBtS/fW/tw55q/3E
HkI8soAryHA9SABs/VXEhI69nie3VRfKLX/rI8A95SCj5TCWIZju//a4ifVflmbu
o8owrKjGm7rbKYbxudU5BSxJhFEUriqCFFOUEL200N4dNtugCkYArlZTMuuR0988
j3+LJpKUElFqdVO1X1cZ640BTwyJ/CTGr8YvtFvG8wgLmhVRg97a2t09bt7eDreV
Wttq3cGZY1HCdqtX6SOP1PhtZdQcOiZcyA156ED7ODdr9piCfPVa5GyFNwzvbz41
+E/18TUCu9iq17/Nwca5F9q34HwsBcBM2Zm8eoVau9wvDbpRKzq6vhOZM9sAU4JG
l+mZcAKFwj5pyxgN8FANtuCDbJLuVUGnzhgUrnQqW+QhwNZiYjYvdLpDZpjxI8UE
SBg5FyS29xQgLM/p29BAhCTnNa9H0xwNRdydaSclsNgRYYJCse5zpUxBleopboc7
sooFpFhs3lZlHs9gs9d+6EqLLX7IYINoL420q0SbqQL2Q/JqZXbkKsFe1723Rs9m
AjHYTuJkYOrZyGwQDScUu0jtLzMuF3lJ7sPUrBzThCzNXH8AAnbXbVzmm0FkGaJ+
LoR7Bqq0XqN6xLMlJQboybHbCQti8QOG+snDofY3YltJTELLDsqkZDEvchC0xys6
FY11itusHdEhBxECESxKLttSYTHMRpV6h+qUHPuIwkT4DJkLv3e8vzUgjPRVmX5I
bqId2tkXR7jJnhHz9PPdVeqD5DgMC7qGYDubL9MX+cW72eOTBn+ykxfU/rxATN8t
Ytn9KC0GrWRjD7CX4/F890ohOy0rxBU2ZTmVQfNDlr3HzcknfdEYd3ofvhyoQtFO
ydjgnRafAvccfi6eDElWmEkJgd7WDQamj60soZk7A8Px+IsF7NEV4fMsn6LOM70l
4aFiwXhGFnrYQLXyI7lFxsbPUcLWlv378VDuwsLyAkAa+Q0n8tSn7praVecPO99G
vl4YQ3E1smFO28kxdRL2gSsWyZwlr7ozekGErdNXnqsvE8S834rBao3ZgO0gK7kb
Gj8q7wzc82kQHQMm5VlYWE4JEeXhCJ9zIz7OIJ+UwTgO+ap4clgl2m0KVa/x8sWe
LxSI/vosvRJbCgl5nGhIJ2q5/pvQAFj6vidULcgrsFzVFpQpOW1PulLLdWLurQma
QkJNgoab2MYznxkpx6qxZKqoavtI3np7nPm4RQ/urpm2NO0MGr7Y70HBOsGk1jMa
deiSj9E8121ymkoKh825c6gmAZroWYg2d9NoS3kY+0iY+YedW9mLGsazredZEhTa
J6Y2180xSSkxJotjHN2g73kJWtEbkJG8n1SvAuR72GR+Ji/w2i9wmWleiPfEB5jf
rJNoZ+cXwtEIWRbk4/ZB//bNVVhTRBTIdLhpbOatKZu03jnFcmnSQ1WNFHukWE2T
Ci2RaEXNBnvok0urYiROS+TjCjUO24j9Q2tJyHZjp4z4CsDwtVRLn1IJMHM+WGY3
/zF45p0a78J57U+ix1scctaVM5Z9ir910alFqRqmZmMaNupIDO6UxvDRNIIGg/QQ
eAb283geX2st0L+XIhARi45S5K08MkUuHT6rElFxFegEyYm4Qqt2howEhGOjSdFN
dMMOSfV5aHrxour4pzipXCb2bT6kMDbR5XY8uHIlLUBG5lPMlzrKv+xtSG+52elj
YBDfR+O7UIvXHIhkYJTrpefjOcY7GDOCMrtvv8yEFQJfaXs5T2KCwtxFVmoNFNjQ
/NPpvh66otpNzQsGjE+5osLw/VeMhWM5fi3Vdu1B3k7u1sVwKva+LyjH9+JKS22p
JdUORububy8YZsntp4CLjuORxPBqq/Dl80v36amfhgjEyg5THl5A1cmabmPzZkRt
kNC66ufRVEvuODbp/BNOANfl3miboogRaCBrOXLNOR8Iy2wxbL+NBDAFjkrUHq5Z
Balh5s1Q1zLIaHKx5Uta9PFPWPLT2r9Jx/rDqXz0G8PYYHYZZEnpewDxFu3Yw82i
M2vqoq1tPeZPF8PGgF3PFFuPR/GPCI5VioptWvi86mB/mlKb4o8C1/zncTCABOrb
LD4VFpWvLz8JENzPB56SWKHwneqbBMbtDoebxjVqtp6odsqQQcYainxK5AFTJh80
rWTy3WEN/mLsCiLIWtSgutPIUMlF0jJz6Pr9KqC9/3ovBYhb+o1NA8XHlxuPiHos
/htontFGzRgQgptucS75mYywFYBDi9Z2vAVNrMCo4hQhaS4GcEbFn67EFXwrLbvY
ebNtSaDvCwdnRSDmVg7s5aBF5zMrw7fm69LXPV3/6o7bWGX1ds+Ssz3C4iGFHBwd
Ds5dMf0Y4HH+XOXrW5G2WN7SAUHRKqnIfmPKYFAV/Bx70bKCiQKKhDQJGXXSY/J7
foa1c1tqhlxoeygV307QrLC44BvrMUK/knGXco/m336tjOTdikDu+6DplBym52FB
Ph7hj4XbpIOwMzzDRMvPAdMVtAKvfhXE60gizmR1mXcBRd4LIpSAi75Ze4QDc/Cv
kzYADSMb59E8WVIDw4I0hrbJCRiN8nMfIhK+cYo0ivMvVGpgp1yo76QjUnMG+plO
Vu+8dcYppxv4BxgDKoO2YNbCZB2T2cFlIKkpeIOpdgW+ePEDDxFMqybT0iDM6knY
CS4Uhr/vIJr/woGobc4tsWTP8pQm0Z8ouYN92iC56fgJonSm1P8c2HAFCCmml518
qT5S4pvOu35FSjOo6Ps7iGs/V1tJafR+LSGmqGLM+mMm8PeYZTyF7PlxOEu4DoF9
nNmxsf82/Is/yYCMM5yRgYrc5LCbPupq/6UFIWDuxhhIxznPndhGOa/0Q4/8oczI
HcGwDaaoVBPYHrdxY12nIQecP9Y2mjk2YLptKcX2xKICnDj0+Rxz0VVsV9dcMQTY
`protect END_PROTECTED
