`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SBMEt5wc6ORTct7IShMqoEk/BRIYndNpBtfet7PRWg6E8+Z4BFvtiXUrMXzvHSlm
K/4vWwLtjJaXUvMxiEE8F+4q9gLglQLDuLdsk23G9Lr875zn+ODAGVs4bUHIpIKz
B+HjVaUZjN9bdtTEUwAz8Y5zvV1w+Vei9j0nv01YjWuw3dcRsEDB0IjfVv4rroQa
z3RkKFo8tZJt9BKttkO0TVlGy109X8Z+wmDygXnNtc6GWMjGmJLmkbHEivJWpMbU
A14ZfV54jgqvzitNqgARCYsOystV9qJKf3kfdD2N+3VJxb3klNQhjWmuRf6I03L8
muLAJVziS2avJ2sfJTW0zpJI51wmU/2rPRuvesbiboYUHps3Qg50p3UA1FEnqWo/
woAuinulB0PmhAg/tckpzH5r5CRLwCHpCTwhHksN23Hwg/d44NsgrkRML/BBP5r1
UJpjyYonahGalIEDGkLx2aFdzRCM7wfmPoO+3pQaP5goqpFQeIkr00fY4BYddTah
K5hhrO4KQL6kka1JEWIU/QXes99ycF44zqazQV/kIJbHrFe61lW3arwyMEB/60qV
lPgF8c5F3vJkWraBhbKQ+CgbHDnS+YFTlBtg9M1WUfs=
`protect END_PROTECTED
