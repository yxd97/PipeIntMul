`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ov6dgAwdrkUF++llThtbg6IZxB+bRq5A1B0d2N1pRQlPioayomJcKfGvJP2xj17L
nrLBmamAGy+hH0TmqmuR/jxoSBBRjDWlrEHXK8lzXjno0EaUTf6jldIGQeEIIwTv
rn2iVyoS9RsC9NrNZdsnQ1QiAgvYlCXMkyPFe2nD4NoDTRr55p6xLqtRYiR65YWH
o+npKcoOHMHgYEIlu1HFZUPc2T8FsAQ4wQT+pl9lvZ4MkHM8N6PgSuHHYuG1b65X
C6pI9bBM2Novt4ejhvyQLJjtcH9jEo+5IYXWpCltbG62unvMruHRZcInRpERFBan
P5emdruhOUglP7XhchZEpE4uMk761P2+tgNF16lHpjr5ADEIM4h5K8oI7wx4uTXL
qDX/B6M6nwdh4i67HU8ytvJYX4GDKvr9HkWx162fCHyMWBfUQZ97MQK7aIdtz9Ni
bq8K9anf8X4XddnIKfC0Yvef/p6TczLaAyms0qsl6dK5YFBZJq+WJiz110n09c+4
AaQKpAM5Jh0VyG3oTUk+3lo3Oc+Wdx1D8nOFjqHvy5Im9foy3It+9+33N8eivk0a
wMDaQjyoYLF5oOsX/ugSV5OxzZTp5vjGVmQJW79srFq6dvKVulYw49JtTmTqeE5C
SSzgFjuiR3DJeZ9Tmy9TLOKESGwXdzAcpLkEisxfKniln8NuAi5eSLxLt5/WkOEM
hjUvawAwevf4nr8Haz7LGQlGTEHK91gyNXff6IZTxoGhGFF9uL6zeM7nRxRZS98A
ZSLSQxzjjWdYypSL/yAplF8Si9CUU9EcCaLKYLIlNH9vOnfc8eIQWK0D99MDGp4g
gXwBVsVsTxRqUI3WdL4MfCglmXXLU5qJhHyntMFnDz3KrBIesMSPloMFhwrEJ3/f
GxjYdeF+m31nuKACFNb9o1Ecp0GgVHHcjT7qsoaRMxq35hL1ORepqT8VUU9CyuDx
XY4Y6BEZj6PLWEdi4yZnOxs7BfBSXPfCk44b1Nlm9kzgNl7Pq/Q0dSNZBsWSYH4z
nOjjrcFZkbbi664z72KzsWySDRSyHcYxtTQ1kNIDvJdPdPCziVIR219OXJ2AGj7y
DFitwq8VotUxofOsgzbU+GoRWYx0uHIcIuVVMIXKnduiXr6DBVILbSEihhJoBDKE
/yfPYPW72Av0k81V1CI0WVLKqyKBSa4egHbDLV/RBWrCePPjtIZgn0b6GvCh2wxg
toFe5NnjVoQNK5r9LEs0UO1sGEGVMBAE4W6xJPYS0tIH7oPcpQ4hPVlDITEXgPq8
15xs9Qvs8sLBQzxAJkfZBJj9hp50ZQy4Pk5MI5BvmwWCrR4Iz77rNI9NWcO1D4ne
q6KSgUbOlvERgLop3njPgDKVPOCsHkr8/+rMpRu+m1Y9q56VRdgB+AWUYh8QFoGW
TH1cbB3zbtAr01tRKiETBnQO/1/MXGnkuswHTfGBswOc5DuTvvVQWsec/nMpRYwd
WU94h2zdRHjrdELr6A1GHV3KzpECaTmgFasmU5vGtNG/F3qPIUD2Xo+68GF/6rT1
4ysVTvEfd2crW4au5AKS22OGUhuPaRf9vAUbiYG5CvuRWJlmibM7279XbtJrTL//
ddzdaRDCQTxzOyhmv20sJRUEDJo70DnFk1b6wlcxOftq/1hTr2Vb3JypnGS3cJgG
kwe4yJHIYHOh4mCzza8A66S4MNdnW09vARQCQoBL+I5pZVn/WRt4j5yHIg5+h2dn
LtpHiV74UwkfULGCPk5sFrSLspSt1BnSSlHJIzXcJVLY43ll+imdGcydirwW1Opc
++wfcjfjZvb6uVR9Z+eyXw5DIXb4YEXwFxxVW+qIOWfqwKrTWQy94V5FW57URNoj
T8bS1OS7f21GXJvuZx8CMaZEzYMUJnEXORvg6bfkCrxLpIXYwW64aN4tHlbFvNmJ
KGcIrXuYsl3+a4TeU9Gla66ydMPvDiG3/Fz0luptKtGj0mtzVfXia11B/HSmKWzW
SqbE8OvE1/9QFPZ4lYH8WaqpxEcr0PIqcP9kzszOnmGbypap2/sTuWQnPgjXoC5R
ckY0XU/YpQa92ZpOZivTLrMbmUsybNwkivz7srC6vwdH4lYrEwP+2/NIGWHF+nOr
gZyOIhmIZz/xlJJm/8pnIPXHPZoqMUYUb7XZP38J8PljqM2LcHinY1pwbiG3LyuU
b0bLR1MFyziVmOHhkvPDFws9MIojjTrfobHSGTsNthPmH3ko1jqUwpTi33WU8guV
SQ5tAynaRBfYp1hgwpUDEyv+LpHRnY+UQqRa6I11KmBzQrgkaMmQiYoQa7jQxTGP
SFS2mskDOwdveLayCw06HG1LXFL2BqzQ5Bzn7dxxWk/q3U4kSjEQMZmP+fHNWCMF
4r1ZcDwDq9JuWMUYaGkIMCHjPb7hQ24HO+nPd2bMbr3GT8B8xKWdhoUoZM31Yg2W
ryq7EBMa/db2EIPJAiXfAFh+IBKVmQ+U9B+UH9ry1niI+xhkknRt0vJs+p9/DLYc
r/UUEn9V3ANsy9jTXfacUo88FL0VwecLML6QFGqQDbIbWlOuFs/JrhhtwIes+06V
oI9P7r4H2EMc1Ho814aYRA==
`protect END_PROTECTED
