`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BcZmL89NWgyUJMG9vZaUjabnrFsho3I3zuhtzLSGugMmjdUthyQWmQk79ipBM9FC
67MQTP1YyFzOGKiNG83DGXklmTW7AEwv2n76VT1jjbFEVkhitg/ebEHcEjLuKFoG
Zy5YBKvycrQEuHXUxhs0dbzYLYFLBAxwZdRoDwY6xvoU8SdBT4AHOYnpnBnakniS
3Hmfa4OpzBUD30p1VCOwCGj5vM6IB7WC465SZWQZYAgAPTMDebwlZkwntucOQ3qj
rHjzTnQ4JCoEPkXHNrPhk2aAajPgI+nzi/1ViciCo8qfQ4SrbrbO5xiawn7Z0nwU
GU80aDRQZ1hAXxAsP9JvL8JZkw2Q5t5bmfuqWUDZuAYY5v1e+7sbaFMZvFkcOU/+
neBXHy1AJ36KaX+DGRy2s3M/Lb8JdBM/PPobcAcyimhggNf/Q1/L8WVlagBqhCWi
tVxkYikxBJtt0jdpKwAk1S+jicrvpsU7pp99Qq4Rl4sFiaLyOY6C2brU0cswhLrQ
`protect END_PROTECTED
