`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ALB0vyCzcfu7o+RHsoE2Tngk8lomAH1hUU+nyTeRER8csMs/URclsU2AswmlCSMJ
pXB2PQxe0VWhu061LH6BMewH5qPp6dirdwrMbhYRT5SrbbO/cHFNs6qd1sM5AX0h
t6zoMXnRasBqNMlP2zBK6Ke94vhDsXTv/YvWudaDqnJyzlAnzsktO56EPR4GKUXi
XgE9ikuG/znfO2sfugEbFei/BvlzIZftqnKHhc00/3WjK2I4ooyEYce5OI0mXJwh
klSDjbx0/KD8CtYIKnvPhiv9uPn56HIMNj5mrPfCBV6m7wKnKxgMiglFUfO73mDR
orh5+xMh1nO7oK8v60mSdHmJfCG7qVeq/RsryFnJMSaGze7jI6GAd4bfgPxWxN29
SDrvmHcYpGiPsZ4LrirNICF1FqJ1YEX7PQ7ob+tx6fhSQwv3JPY3iyolgu4NztuN
PpugWbKrcYF72u0PXxWNsf0hmQtSfynOTwqpe2YXvkpcPnLTcctNQIbr9e8sg1nU
adpj6/T/S39muewd7fNZDr0+kjOB9rxjUx5gM6R9A4cPgkx5AMY146jvyQfbJF+q
royw1mIwlzpPjzwLTndowVQoBzIy72mwHrRjthYiywecgYAdQWXU+Rv0Amb0PGbb
+2ZdFeoc52KPnN2u86lv/5rXZ+xAcXqPFiPTIcHKfIM23PPsSzoJEVK13oeRM53R
7WPnDPqJbU/Yrrp8zlAS+Rggyi6XNDBLNVhTj5tzzlxB/mNq0UVfpGzMhRxxt8Rx
QCupZruRcguED/+b+bwUkl8QnDALu5z/LO2RfuWoWvWxutnIkcLtzcoBXjbxOGhD
WX8Gx07bIPNO+eNqOFVkCr6wHiCmIJa4SO2zbdb3jrbHY+GK0Gg0wejM9NBXO9l4
8Lj9WjOURvd+rbhRfyGTAZvnzEDqWnjY3TjlBn3nVxiKrm4/KDWIL3TAkpMMXPQY
`protect END_PROTECTED
