`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gNShnVmiYC7K49TNYoKRz1+MyCqxgyfj45tY5UKbKBVsOh/3p6J2dv/5COXLEBhD
bJT3b5JZ05AOlyQ/8WQbomosZKphjO0D869ETX8NK/VdbkDGENDr9CwNqltgKYJE
sgssG9ltCrvodJd9txEZYPavgp4ArYzlVG/QeyKQvAt19cLNuyR3XB1vhCtu1BV5
WOQKL39WrMiTCyQihHlxOqAoOc1to9qTSSYaF3C7tJ0mxKIK7z/vBw9ugyTClNJk
ZZUw8jeeYwsP9RjUlzyIVCmp/FUMbQZeRn2fTJYsb+mU5K1KKnb+m1aRcEtzbtH+
zPosq3vS8f9aMjjxqesh6wzGeyP2Vv2/QSfp6X3PYshycgb9QRNcGTuXYN8ABYzB
MAx+rciK62YlcTGFO1HIe0RXcjQeQZxTPLA2g4qk2AKGWhQ4iDyeuaghLUCi/hvs
iA+0pK3nUwbEYJB1T8I1ezGNjWcsXrPAZ0hWb9/DMDB9D7TPdZrA913D5Nu+drPn
bdop9WbkCD3C72DR7OtoGv+k3aekaO8OLKL2lCrXoUDbP6lP1xxviWu2xuU/SjFC
Qv5RPTIrZEqT+8h0umhRWjMT4ZjZIbzXFzNjiPDjTTxOKHLkVKWJ7P3KHAFGWK6c
oZLzjT++npmCa3A8zKqitNjRWVoygqJY5VAnhb+1oAIsHjOXlJSAAmSemg0CS/5s
lvtNXt5rth7cwgUzTSjj1/mwqFQBJyaDPy35S/L5ikLkczkXM2yIsl3V2d92yxeM
X5wjNegTT58EzsjrTRDmB4VWwisJfqsS+DPImaPAwwB2n53inve3IkP/sew9zHaE
PwdFwDL36qJ5z76roT2PFtlRIeJfTTtD3boLT2E5K9nou/GX7s0YLK2cxZCA3+pg
k9kOoIFBIToVnrlcZeNZIJtKHbkFAlut8cvdjtxWZ+Fr1U698gTBdZHJh4O/Fyvs
Y+29e8G8TlldKyelhpT8fP5gORQ+e/OJD8lbBG4xNdRsnHlTlU0GC5odTsKS1Cm1
CkhoE13rGfIQ4TzKK1EWxkNWEF/ib4VdqQKdmUloUwDFj9tpKKXNZo01PAk53eN9
SlgpOpdf6+PwT7eFyT6F/6z3pLsSMWQBtMcerYxP8xG3SDTksnD/w/hl7YucBoaM
etVGX/g6O1Abu5Z2p1qdCENvxSHJ471VdtQRy/KrBufWTUx2srsuqpgjoF6gY+oh
JjBXDErlCn0lMMqW99bFbStjyl3Pyjsmg37/NNoXBEIGTcOiepPJXPlqXP3XLBNt
UEIiXDZOtgS05sEC5CogaZxlwn1JYJ+kgaLirSX4t3GBWutPbhhm+/W04WFCpyTv
7ZLH2d5CTEGkWVXJ+NuDFQEl3zLqQPQDGbuBiGEsMdPTNEa8vO2X5oL49s4XWcax
8WCRloasH6c4Qqn65+u2YGku+ln01kzFqNqs4MNgzYWfAlBgjiBLz7XlHqBuoM2x
hbbhvEmW/9JI39RBUxnt19hGkYa5WWvUSljybQ1XgRhfBxJvxrCu6EsNexVMsskr
7rgKS/6D/DxL5ULlgl7s+RrDefHFgH24IBmIFcbXWa32XmoG/4UHUPKJ0ZILfVms
/9R+yHUJm3dQrpln6PFnxviwnJPPUsTgGZefUNrn391cB9TWJpvc7kb4udrvMGjN
pr2UCYtBbF0G+Ao8Z3Uk9WwfECmwrjcSjPpInQMm7jWqTt/ynoCWhE69ilns++DA
RA/eXURP9bAMmO+TZIyDubZgc+wZCa2rtR7s3kqIVBbNQdjOVR9HRxPGmb2gKeEa
67VQqJyjNQO+ERDqMP68oP9OwqSGVGQRTvWPAuzM+tNoZcuEk0mFjyknnDFOiipB
pR0CZJPrhjw5y58fRMQBFeZds01MFQ7cGR+zuT8L3HUGSmCbzqst0j2fMgw5tF+E
lgCEeKuQs3nTDgsrzEFYCHXAhPui9PZ0kw6qket6EyzmNY2Lxcxvk9+vHkEZ5cs3
sDFK5u+wTAsjWhNsowl5/yU8yc4b0eaqUDlfmdsGqJsTyG1TEROTodouG9Kp8+gL
3uNB5fhMgUnpen9FwS5WBfNeyeliG3YvgahpM+qDjB5HlmQ5u5J+Oxq+JWDe2Lqt
gzOQsbr115fE2wmObH8FDlTWfwz41eyHDCK/X3lUoRiIMR0lKt7RSvti9+VuxNyl
seBGYWyJtId2+RIpwrZQN5hMsy0g/KJM+sOIDSmSFmyO5Oe7hM52Mm18bpvRMIVy
0fEp64g8lx26opqlzxd2e20yaqxwzthINURTMCSnrZh+qEl+tRBEjMJ/teU2yJYh
Qre/jxstup9lD8m9rHsL3P6NVDVq7OIDyPf9wra9I4exPryDJvPqekQi6NBncpxJ
+XthvrwOXb5NeQCHmqjhxstmV/T53chUg9J0HiZpGwa8lcWHIXdPXyfmrWqzXOVs
LSis8Z68+J6p40oupX4zish1KtSY6Z05JczUebEioxEsDHOa4q1MFca42xhBNRZI
T5rlAx5qgeWBn2vGKKRIE20/rAlx6UMGBHUccPwaSpEIiv8KKEhac84cVRaX5Fj2
xXLix4PNpyFFIqhdLaZOldQ11LdIqBfE/gz5pVGdPshZdrQb07bRwHQGwbFkSLjy
GaJqwdRkQhCyTtANnpgk5Vka4JNehnoC+msZCE6KFyRizm9zQpd0fzY1ilm4fYy+
rcDfYgSD86cnJ2rWE9nqAiDL7uZ+FHkBKnGeVNxVC/4ncoERDOnVr7iaRBebIul4
VWiJuocuPdY0vspGP5Y4Qv41NwyHqyJbDlV5l5HReuKRH+sLnHNyYafk6kCsiQ0O
8Qv/bC7JnE9jCAT+wg1+eP3794d6dQskoXVolqUjbtsG9Q3ViV44Dr/ZprqZEQgJ
dHDLeLP+Sppf1gKgQ5QD/J8NfXpMzYy1lvOgU6jfc9QMMR1MEl6jd6PLXVRVV1CN
wkOj8JV/jsvYayzo9Si4QRaxr1fjGeKJiFlOvb4J/HDxZtqC64LgzDICGgWuDb6A
hWnuAI9eAdvLBaqt5q+HQk3PN4pKWyEm45hdOS2rgiBCGoQ4xSFQFpSRzm9JKsbb
IxIjtOAyTGUnGRdg0x1KfAxqmV+vuasNytP9UESsqANMjFz/Oha4TA2tA6WaTRZG
6aa6mPSZ422QIhCmrHyI7uiJDN4mi9XQBeWNYtYFCk0cv2wttbQV+qIa7Uh/SVbT
RTb3DJG0CWf33U4qQkU82GCpdLg94y3neRJB0EadJ2OIXlluQEmQxnrwrOccPKry
upb635j1CFQDIOmozH/mO64bGXVYiJTWTiqjz3XIFzD8+2P32Wofr2hlBBWdvHsS
xaFs9oKHBpMZQaec74tVw9Q217G6buCxbHcFepmBtgYaoqhtOiSQgMhaunUgftqU
W5832IDc3QJz0ICeVw29dVZbwWoIiK9btpd1If/2G5HwVY0yk88NSEuXGALO9/xO
331SreUFCoy2r39xLvypFxKkOtqFhX2mXEBhwi8b0oHXDZqiiFI0v5JF+cUgzXRW
+Vv+ZCvl4Bf8LXk6E+PJQoWRqQeo29JawECcRFyV3Gqj2RkEnr//8z0MkVwZ5yax
/0zhF68PKu/vhxYQMmDma80Fj8PzNRygy/GtoZJKDQ0uhAFJaPJ5BVgEj9rCvKmO
sG5Dxsjubsgu48eKL96ViqBFCoSC7rV2y1NswQOOnChbCncWcWL5W2HzV285k5vM
+Bf0XLxrJjIyrriI1jj64oYsH5SIiUF64UOfUGl/HVSmhmgJQXeCr79rHg+VLN1B
yK2stVaVrko/JuVcXDEsbfOkd1jAdGwz3Pb4zinwb1rE0JAaaKZ6r/Vj7sL6Rck2
OOd86sEH1F1xUR1+rDXSPMHHL2dqSQKX2d6J2JevGE3kMD/hWZGI9K5FnI/7eNp3
vSYFzVJzJJssumac/HNxl2+ygG1io0W2Hni5gAEdwgk3tifyV07xi89yYpGxnTUj
l32moWJ0u+hvnEf7fkHB9/dy7HE/wCwNjmGrrzlVYDatnJS+RT8AWNvo8aXwJVRK
tQu9RwcjtPmrWQuy5KtcRT6/hZseeinAMZS+nh5qwTm3odKfLli+0YSsuZa8/rT0
w+RJjM1RpzSYC074sWtd6ZHJzFP41gd6FuGVjY8egTA9GjG2POoDXE3BOoxHm24R
R+KzIfqtTBJ5OyUn0SwJnGO8WdFGYlX0x6e36xkeUcPR8Y5TFRmwQuWMPAYgH5F4
2k0621XPA5seoDVq5Csic1z4RcHUOecApNbHVwwLQSDWGM9+L8XEsQQ+YFe4bxwo
B/+yYxGqma9tetwK4YxkEkeCr/NQN1lNhJ9L+M0shSm3sdLC7RxbVisBY1ywrfWg
Q+uoB64E3KbYo5lFN7gHbHX3XEV3iVxf4pTfuC9WsjRb/YVxTkGr14dHin5kelvi
miqvt/4ref8LJiue6FLxGhVZCciXnZYnWHTF70zrVpqJKlbYU9J7xypDumxeR8Sx
dvRf6yykhm1+nxCmjJRebknwmiCuP5164O5k49Ynv6NO6PhXGa/lCs+MiWGpaGz5
iY3wlrv2O6MsNGbC2rq/C8t6OX0Z42BQ/VmME0PxhOPCVAWuTyxXitoZ8XyfaDgw
yyM5+fh/kbH4D+CsmREsU25NHaJmqGP8C7sqFN+2Nmiilp+hdR10tbXmAG/GCrxj
F3zYjnJVHwSCrPadUFC+PMe3p0Ukz8ZMS8KV/sQixjC8LLcz8whLl8fopzGfoKFe
rTnMO5IPQT1tsvWF/lE8fUtdOhssc+VjLbrFtpwMZr+61ARtw6xM84lQ775MHBQL
UDco7b39SZJgDlfsd59NCL96aHP6T3/Kxfi9XVka+5BiQOUHFXML4TbbLdMUpkya
b+pZDU0u6mTsSbF86q283YNhTYqChtD3cduOxdgFA0pQmoYU33OLM5qAV7i9RXYT
J8hq4XgCivjRCN9BzRaPxm8LTqdRRjFdG3uQ9ogs9eG6kcbh6EgQlQXq41kbZQ6e
29dA0hol1lmulcbq3h5iMQoc5/RKe0ofMTKP6pzJEZFVVTo9wZrypyWZBWLRq6I7
dmDPRcelpuxw2uLs0Eyb24XawzJ8SEwFpEMEYHLxx52A0fOKx5AR5bOMsPc50i9b
J4sADfBYk7FVRpHolvFOJaNQYLAx6G+rhFfcIEwSSwH3RmMzK2r0xIFR80BVvXy3
Pr7qRtSht4MaOzPj31Hy5NylWJzblVYC/sv2ibTv9dy1M6oD4mme2kegQjnYxqcI
X0JxAuJVSTSa91n/gBki5tn5y/izBDMm1GDC1yNoDOUXe2ZAygKNZl0l/BqLItJs
cFdSDdmpJb+6vk1SiGBC47+RD7n0t4jFDGwFRCl6NtUJ6SrRGnacUcINR0fyXT1M
JTyH6BPCDfSeP8J2GmVXzmhjl8h2ndSOMsQcffMj/1xD94KIfuxTkj6ocyBqYgjl
IGmCb7cI+OToPg11woutU6AL5zyw6OHb2ygpgSHBfMMKyNdKfOpojOhQRIbLGBdA
Nw5IUJFw/JcXR64h+AoVCwmLdaZ0+1YPiX7JmOmJzXHRmRf+9TbyLPA/yCeyIDqK
yxS4dvfhpxtsxgF5VqkSnDhez2HKEh4b1E81YSPsZ4z0jMvEg/0TFD17ptYLQ9VT
quUkR5r+027Z92o0ilkxaojZcd1i0LusQqZNnEjgfydI6Fu7iK0x/d5ruMHML7ja
3ie2e3bSem7ObAsbQytq1m5J2FLGup3bPSc3Bjo5txLfd6YAOJlpyVXwA8hOycQQ
vI6PPrI98WPqvTyIIitDW9/R0bAHdT+JNt+SMvXxq/xxNClHdPbUIyqsa3Ctrk3W
GV9VPthuXdh2/ybTaOMsnhqFETBTg2xeEWZ0VvXR0RKWf5m/AdYmuMA2YD+tZL25
H8MqxFd1NkxB0vRPFOk2apbMi8+mWupLY1lKB9MI8k6lxqTkOiJone/DR27wsXKN
xh1fBl+5FqWSe0jKjDNNTqwNipGjP0O2iRLNnoSaQ9bmqR8jrqlBBm/kSZq5eXUA
Dmpp1BfsIu/dI3EFn+FBGg==
`protect END_PROTECTED
