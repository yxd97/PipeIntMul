`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oE6dzM0wu74ajKSiTlSRa4Mlgh8kJ8tfhJGa8ZE9zQ9zn4pC4KKeOLEk6sSThkHc
sg09MLd8D8z/YN+vNdkZn7hDfwO/SfvdRwJxAyt6o6uQgT6HbXKI8LEcHL0i2PEM
RVPn2xHT4BFkgt43bqFlVWbPx4jHZndi2yTE1YUVXNWcNv8F798dfLvX5GZTz3lc
xo6ChtGNexuHn1xByKw8DyeoAng0I4z4YkQivQ98H/TkPlfbzLkVHQa0rvTy44+a
oJ+ScHVUur9pUMaT0gMEEegbE+eCtI3VcshrZtPft5g=
`protect END_PROTECTED
