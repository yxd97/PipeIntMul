`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AsOOOsKgGFcnZ4TIBZ290muvGGC+uAqzji/bw1ru1b9PNrfeEl08k03RrQHlWoch
Um69zpXV43fxrxAs8hKwTDqs68nBGy2XFzu6e9PJ2RbqcFMS1CkgtnfCEayUL5X1
IITlvHG0s1hQLD5dr8Wz4KMZR0rOW/CcYZwWPR/sHnV6+HD/li/OEMhGPYdVj/3g
1vDmMJKFg5XMBq4TE/yHEJFva0uJFloDKGsVnTy3ZOBvkFykeZLouXJx/IPN1m47
+bqC0d2W7fiRK+zwEcYHrYImDFaOc1gGTSOXmF+b6ON6YQtTCGoQx0WyHhcSVSls
ZuS9qrPStxvI+o7izyxWfkh4KAsjIat4Kr2su/xTw30eg0nOah1KOY37zNbFTR/Y
PsW1OdTdENqCBG7faqpETwtoZV482yRSSJ2Gbs4dJd161RY9YaC6J7e5kZoR/5AS
VdcjjGGIDnJ5Q8CCFTiovMOZG0I0GB4p89GEu7f142tIkDbBZKySU+O5Ou1CbBy0
NyAxkN7NaTNKCnK+kST/NtPT3wMtGl2FUzFveZjlrjELAlbWpYBOmITS4rBPU0MI
A1y7CkZIuJwFNKxazsB98QB0UCB9gIRkDdElXPeQLDF74Sv3AFVZomRVans9JfSI
QZZ5oiB9KpLfB5hcmKS2IAnCc7IxBUT/xCyx1dhEbuty0ca5dBM0tQGJTDuoi7Zo
x7VWlcAzRYyH8J9zKNiB14EoiLx9SXfMwAwvwafFqyckZXqHZp8dP3u5LA47NtWm
gnbhmHROlA+JENC5D5tJug3uYy5ej/lOvZtk9vsU9Ca0VE0gvy73DJTPBSjmouLM
hOPbOx5VTtyx6e64irseAiliXlfOb8cvJmGZr8MeIt9p93iCrWYrgfONhBK9qasq
7+ME3AcNWarvgPrGB/bQ26k4AT5/OADlplDXdFULiei8GGCiTmO2J0eXxv/tc4+B
TxLKEnDfxc8Bjdi0ZA2GNMzNyvNDjWiUPS2A+2ZHYA5vp4c1E1naJWYOiSw37w1G
AVtVGOmwuTjrRyvc5lfjCdSFHlLSVjsbjN3WyngXw5Os1zfyQdeKCYn7PoM7okuX
6Z58oZJDQIC3LDvGBMTOt9eMv/Q34SRxnl6olcDxBpy+CpK7oGByvAnLV6kO61Oy
+y9JZOX+vnzGNJ2ZPxkpFq1FTUY13EOcfzvIOv9rVgHJcfWzzZss59d/raCdqQyK
Bn1QETI7kEMnBSwmwAvEfS/80IAk5ZFOE0atgpGzcJn33J9T7V3PDg1U1PsUIq2A
UqPsDHDgz1TWFhszun4qMCP2yG33+Zbg73KuGbGSqUYp/mhRrGDWicrNfdL9VTBE
Bks8d/DpxSU4UeJhJuhLUZHDkNnL2HyJek9m3C8cilGmTg/0ar5uLQcaQjQAIEIS
n/VdwRWU663c26GlETuMD6uPQuITdjwwxsArP9Ev7myhFsRIpEvUEwIYcyPWmuYN
pQL6mC43wOjMckEnZZY06RB/O166LYfkgo8SQWfbUFKfOXXOwSNdgMWJABE2cjc9
2xJxQAy/IA9RniK7xil7erAmZ93CYz0J44Bknekcp0ISpAiV2JrDLkE6nfMhSi8Z
dMOggHz1okT6Y7p3PlW8N697OMifnF8E9GDNxMNok3ZloZ62TTALxfxRBSJ7vrUM
AVVF+Ahvny0CBRQK+OWEFENQ63XGBpQR/u14X0bfHshbLQ9FUEZzqIGnQicK7rDL
rUEfZXQlA9g6Hkslf7GAzR/jNDMGqr+eWIWjRsq4clxJ9SDWce52BWNHGxD1okUc
QOJKFI9L+nGM141VFNQbM1+PjePEgoWKBmfqkmGGYIUKVD7u8yK756uQnyMM9OIz
vrX+FNbXd1AgKcWnZk3Sct7TW9XuOOBeJU+Pc8XReu8z/EO2sCygKkccwIlzOnKP
9TTQRM7g1bsQbrPdk3IWwqzcexu8qyAHrnVBqqndsLRTaUgMo7jQfCIlBEt7v8hA
DfG38cgWpLOLhSh2a0X6aKcpx5shsxApyA+tlvmpwWev0C6LWmshuuBaFt81t4Nr
00fVFz6icJ0wW0Daw3ymt2GEJNWUhGHxUh5d/IAQi2O7o7K1H19l1ZJQ63tOeUqp
sGdz2HACjEkVmHrVpgSi6sj1CfVrP8CkQRu2x6mUuhe8Ij+XvhDnX3dMoCw2XID7
y4MHWNM8hIPgEw9KF8ofPIvBdAIj1o/f8k8KEcmgO3NMBHHsd+yb9e+WlwHRlQ/h
UrDOFi5BlaA0O1zj7qqWBJNK6yqNc2rFk1F3GgWPKNfMu8fY3cWG35fyf3XWEZDT
czd4M8+JIArY4IyJu+EfZkuS4pcGOagPg67rbIeVQXrOrmhc+4HniEXdD2TOfGRM
Ufq2Mn9tljAHRt0wIXad4aP5RNQl1pW89sNceXPfRzByc46WQInyIsm//9twv8+F
u4r/je/FhbZwGLEHtPcebZwZPzVTdg9oRfev9bdfOz8NVyDiCdp5YS6m46z7k681
yfQiqhKjwqQuhjIP8sR7luXt2cHJQdHatXtWBY1oblMOOJHmI1RofxBlEklZYv8c
XdugwNX823n0LIqTwW0GTwDyUoG30Ub003mObiXKL34KfsBLX6siBw8wWrYFpXvI
kBu3xGS7UnEBvI6J2L0hzxl4B4eZCPrS93UBozg6m4N+wI5i2q4J1CoQvuSWQ+9K
W7g1PqLHT/E8n5hGc86ik8/e0XOCWd8UJegjm2MMD0l6vdsyWebg1cW0O7guSsTM
oBaEpYV0XpcAwbUM9CfiyWJCbZTHNlJPXuOgTDAyISpboAdtRenH3niVcgyBdWS3
/EgBg1tV+780mu6yVn6GXVAc/8m6iOxgdPXAgOD20DwCr4cmNZRk8uSbVm9pYJ/T
BkFhQ6r6O46gGHaG9hCr7a0Vb6un+pWDpt5meTao1NZAF8HNeXpMqOC3pZHohn9T
i1LzKdBSrmUCtC7zDqJ6T5+5rmrakYgibpGFH/ho46DT9Ln+S3LwnkcWGGQs4qJ6
ixhbvsQsRTsiCiKvCOgKKsMfnxfhcFaUb7UXX4V3w+6N5DvkOzAfLvqUx8rcoK5N
WoPAhpM26ZJThhC5STNYlRtIpx8OZdZaVH66vpUtlOFjdc5q7iOmaJDN+RU/yNpL
DRCeNxL/qzaeSLtwUamf2xlKj/0ucztfTy3w0EHj6oe6E3v7Bbdm/KMptOgKw//c
+MkUXg0HbFlgv6JPYpJ9DE3JGeVzR4C9VqExHFH6T/coMuwjNl+0sxkum7msa+oK
n15L0GsJvuM22d3Ak0yjlPQonfkHyCAcoBQ2Kpl+J9A7foCIzPoI6LqUQytU9idp
QU87xmR7EpmmaIylM7MtdmECdWpWNUXhQe6cF50x/+odfY4WRxpJKepodTM0OJaD
KqakqDRh55JFO/1YrGtqr9PYeeP7s7s3jIJUAy2hOFDbRzuv4zNU6Dhk87FS4tFe
EL0RfpxGKS07Z3SHmh1bf/jMvdDyUDLIPnBwsrRk4Bgxpjwx+oyVyyTx0HWssBon
sJMhwmX21K0+6Bn5Nc6yQw4RDqwX/zXGT0iA7FAY15QVVOe+SyDCPBJKF5iE7bNQ
wVO8WqE4FkMqaYHYIUhFv278vRJgPlMF1GgsO0w6/BkvXWPA+g3uHSYgA0UpMBcy
Lb6yhXfAmeEccNyuHPgkf4g44wRiYperQ/LvZh2zf3afDVEIEmK8gseuaV7w2Xkn
YwhGPc/x4qIn03gIpwOoygfoGM2jouOg/9CaQRLJ5/ApcTqzKLKiVS6kIlzh7DdG
dXSbKLVDyUiY21kH8eUf+ByPvdtYI7vhvJ+Phpu/TtSrx2phxluXvUkP8vDsi21e
Pg+MA0FVQQoqGder3Z2nfP8WfYRhnO+qIgtRjV45wOpRt9ktgHl48xBYG+Li6jta
zvYtFh/lQBraxYJkysnOxWk0dJmjvAqk5Tr49V2dsMxQ/D52EhfBL8EdOcNyUpf1
thMc//mzY5AQSjBbDDJjk9vVTcDg3nB0tOKHB5xNw4p8Zb+6qVHDaQrflGdw8eEm
GpCiPJ9qviQxPoqTASw991/3bUFl/hiXCxiEMxXLsuEfk4vATheUiV3gwTnHqwKV
5f1ZtqwMCt8V5DFVlI6f8N8s6Y8S8Jz85WddKIg+9d3On1l7rN/OJP+zT0mPs6la
a20T7nbOTyn8/VGxYfE4izaiXJFZHRLGpGnGhj+JybtSR87AH8CEJK4Av0SqKGI0
rwiHzdss0BG+QxTHr+KwB9TBly5tecw2bXowvrIB3MK4hepEzPbz2gMFUP5tp5kW
h2Dw1Q0dfXME7BlsSZKsV+LU4tDuU72NxHLIGc9VNyJ/LWpyu1Bq145odA0Up4/O
tB/hZbOXlVW7hJqoQRYQLAPLaFPCBl3hYP+i6k+i8VpPo+p3xhKeKNm5rqT228Kk
mdhfNDnC92hkSLPXpxDzhaGQx8OADqfmj0s0b5sy2KBM5sXgrTgYhCLgbw2i10/X
NRPAUeLochRLL7DJv/T2jnnfRxTF99u+JQl/DYLnmFuoZIz6EZ6cWmZEwYyYua4s
CU/5d9eZ9KYdUC0Vi/6oJXn4pYM8uEO1/OzHzE6P9v+a39/u+X20NPU/lGCqK4o/
Lgm26VhTA+vxPM7sgm7NXozv0hCBs7twZUvktJT/ShU3DKQXHJ3rT+v4Ykt+Q5C9
Y6XKTxyhEREqN6VUJlw8s/RufJHrjfrvDI6/CZUHsHZDRxiITBZTOgn+vLnu1UkL
25V5twugby6lIFuoDljdQR6zXctWBqlFOpUwcNb0AYgbuAcfVOkoKjVcddbbn+Dc
uPnRPoAFkLlVULNtGcSnInBgmRAe0QjWzapi6sNdAXoirw7ozxeSQ/JVlT3K4Acx
l8C4e3mwskuX2dKdQ5PP6s6ysxGQnA/wYRLC1V+e2vArsvWVMdzpaAmb5mxFEKDQ
lorAF7Vjt8AtD+zCHhRO6mLZ8CMQ5u4LTWwVhJdRi3tQBw4b9HR5P4P4IK/3OwJx
8bhVZBcLKv+sTf3Hh5j0254xkFkv0OFEa8R9nP0wl4mD4hQELCdb1WHZq2CiWEf1
r3ye2lFRmiW4zf/r9l+59XOR6ETbiau92ByjfHUqYhM4x1w3T4Y3Iorqaat4DCPg
afajNYDg74B+5YqEl+28dgAVpzIqruvAUp77C0cM3j1gkMgtdbvEG/d/q1L1/mEC
/RHlNEPyV6MxPMfm6Rmv7vjHBIGSA/9scCjnO4jaFgBR2Pdp3GS8JFYDYyR6G9Xq
tuy+HsFOX227QJygLUaguVuT8DypmX0Z7eY37MUbLmMm7cg+Y1OiTJpPgt9QZ/yS
YKbGud099hRxXtrXsyjba6Nbqn+NSkbqOpe1fZtXL3FgmS1erBvNl8jWt6tw0CrF
X9eH659tmqMF/mnL+H8cvIXqxmjDXxKafEwYp5LzZsGVLojRz/c3VMR17BOoHNVZ
MfbXI/fYVR6GGUya7FkPo8YaCCfj7IibWldFAYAt2Gph8P9oyiaiHbhl8kl5Qy+v
8fbcLoojNRqAxnlltS5BzaGVbE3LVe2pphy3J5trBlvw+9yHKn+43Tp30BLzR06n
9VCsKxUGG5MGn10WHvBUeCV4jqLYurQz0thd1okCYKPDWijedwv0d4YSfa4BeT44
2ka+08q7lx7KICl/YJCP9Yb/Gz7dizU3iKODOvZM5pYJT0K58WGlZgS63F036Xo2
55BthnuXYA3Qg3u5tV+3vUHvv/KcJd1RGEC31QpYzy/evoRi6e8dlCPnqxf6DKWJ
6be1cdIXhjY+pxLduz/iTTIOGHNwQtlgC31vL+Hls0FGcGScDJdMz/C78sgyrn7e
JMHvrO2Hs39jZpVxSAjjoAuVPyWuZD8g44RSwNrvd8cm+2MBT4Qc1UMRRClf3te+
GOG3xqqoV2mxSRhnfSpZn+sdBl5y4JpeMmDjSQKdJIyUelLiMm433iLlc+3xJ5Fq
S2icIkPC8dw7NDsyCd7L1ca6beIdPEzLjgdzqAAAkr28Xnsc/E0Iuvyw4gYDYr5N
JUwziupwpCPMDBJGmKIPxRML9BD3f/cXVFuRhU2jvCN5KER6HPQPbt/vymAh/0wH
I7Q979ltWH/bfMcbqRCKgyhzVHbgNmyE3Aws1CYAp1jyfzXok1En++OhJRH5XXHZ
MyyDnntpvExLw7Go/3B5dW8HDIHZzrc97ufQygh370vPlbG0lmFSYN2Q7isjvATp
/RxH0CLy4dJwV1sttMHMwh43gm7V4iaXALJYfWdDMDDygxgHuLlHuVeeykV6bCE+
m4AsSmUMk23XFOLIwUYoqxCBFfyr71+S9yg1puj4DLeRRlx/1bBCKUlD9n404p5m
DEwQDLZmKTippOYSSzp4X1PHF0KfrWoy7upf3aQSMYSm8AgocbOBTHQkd4wIhW5O
c1tQKGpMqcfecUbig5xVJd641shcJmpKT5NnwUMJDYog1ur1bFngl7VuSARdciLa
L78lGTKSeF70LQUsiHx1a6SqwN3aq3BTliYL6kjTrk/xPNDexrGusvGuPREyVTEh
n0zG1JRQ/V7WEllw4FObVhW0oIacfiGTykneU6eWGtecp+y9Qf3tgq+hsuUvu59Q
yOmbNCXmIZDhAZsWhmBALRjjOCdGIAhVIp2G4osQ5ssHUxRG14PS7e+dttjfLGZW
46tobShfBhSqbwuoizZrOxtAzKdo46zD6iO8axWB82crzWkuJSNuq7BhSEgguvHc
yj57ahSV6Qwq3A2Gs7EEpH13uiqWxHKn3WqJFg1xrlD4d2uqFAB5Y8DG7cvBfQqT
3rwv3I5KczQmDcSt15nI/O+A/lG3Z1mU9oBmRNZeZVnFjYcDDBUaIczv4XYZ0T5a
tni+UIv5VqwfOq44XLnfk8UZBbG5qHnf9vPEQcomrAUOfvPqpUwlfGlThHdUO5S0
8MRaayMEEhf43sbVKzW4wvLp2MbnM20WB4NhpZThyeIyfiwGtZ9DuqKerfa0cmvt
3DfN2PvwPboTn63buzeFHf/T4enrMAsLP1FFgD+nRv3pn810VptDXppfka9TnzQ6
0JxaCFVu7VkqXM2IP7x3vG4NEWLQ0JjEt8y0YC7b71r170PnYugo+Ew7DHumFi7w
oa1LUfHu1ZapM1swADyd+nT1lHNYFEZ4JGnnm4T3V4vl9yq0kv91Mvpe8Bk9xnz8
94AWRib+eYmUgEbB64GwKNMWePfbsNB8fpztYhDGx3WFrwtmEF48f2i5DzEL0ID5
1WznvN8JnN9JbdljUNslixZ/R+NIIKBN/ba2BTwqlp+7L4ccY2FnT9NugdzKK9sI
TTI9bv+bQ47ka9ih3OzM5s3c8j3Fjd/8hU7YRKEzTwB3+whobW5Y1a3aV6bwFy+t
mFP6nnJCb9jS6hMIyLu/DkZdLTtMwoBVRwMk4L7+Wa0E9o6q24vrFe8u6qL8Zp8b
2fPUCzMD80XldpHN3Fa0s5j7S4MGGxlZd9MZSZmSfAmoognJo7MENpJDFpdZxKx2
yh9t5QO13dFoaQp2guXygrGPAtOR1UnDBCpwwCiOCQh5cLIOZlj6LEKq2D8EKDAN
9ofhOnBwj785Jij5cCelIPcKs1X09TUk/UEkaiREIzWY0xz2cX5hUpZEKSITO0TT
ei2hWSSBX0UHIQeeMC77ER8+cJhi9c+0EXKJDsNIYyyNstWpDVRfawh14xwOr8B6
VfGnwipxb9P5OcjVOgiybHNffKJr8Hon6Z6HJJA8u1o2J25T30IEvYVQArmCNb00
CMOqWQe1rjtx9k8yqkGI1zTFe8+A6yKZYQGcY/ve1S5dPhNoRZeodsoJQMAwxToF
sFGMb7yYizug/usXbftpn4Ignhw/pWri1DoDW6sNoVL+8saplXCx07iYAGc2IYEf
AKl89ijQAqt34qBgOhQF5f9jE4UMQdXC3ger3hq9c28ehyYlCu2ciRFV6Cg86gPg
CJIwNB/yHSUcCXHBHOQZbXlSYl2ypkOehbgeTnEzPgTl3pHD837eqAyNUPLDJ0AN
b64cPZbTUw8aOOWFk4oONqo3rYd9PJNNKlvUbFSxIqLkfE8hp3EPu3KZRKpge4jk
QjXtK/9vIwi3ZyGXwBWhoGcr5LvykYiwoyf6ctL+/O71Qt38NOPHYSA/T029box+
KkW8QsNmV7WvzJpR+JaDUx+TjSrwnfUlIbdTLpkLGtyxfJbBMWmhiwyxTLIn4SFN
TizzKf3WxqJ/4b4da4OGqvnehR+R0XC+TlHJhNkxFzJ/MrSdz8CZ/5N1u92aLwaf
dFNi8ggxQDv0cN8WCxlJuRQ+iaUlIQwwN5Uc6fSgcHY8fjkFomyZOub4ZYijADBV
YWlHH/zjGAYMwoe0UWjere34dqv/oBGXF7YSNUs+rL7uHjLHgfwA44cfYk8Y5t6O
rWK7GYhxh5/3HxS9i8NBDkpc3dHrYkUhIsOzPAI3JbaYlHKH1Il8FvkI4TQ9IbVV
F+2pDSUvJ8/eA4gHhYAM3r4ZY/pfcjJIaEC0wCOLXaDGZ5P2iLov//Qq9af43+R7
tL7SNaeUdDQ40P/c7Ob1CxaNr12pzaUnO76tJQP76p39N6OB9fMb3MUl+SAl2n7C
Ti+ipy4ogjdWOmEGTvECOIPxrKjmw5rVo53imdb4rQRJxHJo4HSsQyq+P+vHlKgm
w1EDlGRXQXlaDaDkp+QXJMEue2qS1+UOKPqEv89xjFIvWVPQS69EKLQa74+iPgtL
qdL14nJmjFHc/SowlkKIAZCK4hBHccZqTOW0juBAK4dtmZx5xZWI2DVC0sd57vbA
M5WmZIFsbtGaBPdWE/2bFrLxe4YCv/rmZaoFgBJz5mE1ifQlMkWik7bvAxvtqG5Y
LbwRO50PZVKFiDxea52792A5c+Cu3nuLWlWWBH3O8AvlPrHovhS3xtq5uGH25nMy
Qqu88HaGcgI1yGlPc9uf53pv/Byfb9TJTjrE40mlWYixHrKkTZF1yT3IH/5Kw/wg
2I4C+24/FZFHrRJM85Vn3/3UkaXBZejSo6FCbfC0VvQIjk9s9nCP0UnqchF3Bx0U
UahlAMA6lUbGpujHIGuJxV9lQNY4M8LMILhSHxMAEBm9mAdc5DDewF+tzv6YDWQV
XLHL49ZDKqiOOn74e4Y72Gf6p9An5IftzZGPvJ6l6dVCDyBQcNmGmQZ4NBghhnl2
l73G6GzHjVKOW6WOzKtMJi6idTF5AlDrf4XaVmDs1u2vZnsLwScNVt7zuntJGjmm
d5doKSsN/lFy7PpLJZzcKWgkGn5S0soCX7+yAOEho0ZPRtrUkNOQs/NTVvk+UVrx
LFreOGogBWQP5t8i0VeuPzMDwb8h3fqQr3q/69TvcoKnAVavcqF4Tmg3flVUVuPM
xLJ5AZspXgJFJ7n143Rqciz41wep4A2jwL25Ce2RUE5K5zBDXH0RyJwj4fT+izTI
aQ+XEg08SH0YG0kH6uFUIovN8bLwpjX7CKMRJjaBuIB2ZB8bAaZRIGWIbyiBl1DW
ysEgHXz64IlbeLZ9gyOWrdlSczwRo2v7Ou2F5D4CIWLxY9fdt+JUh7hF4TXSFsje
Zmj8JlFSm2umf7T8TyIu62i2j6L7bdFwmNykX2BxjSksxi5J7zayQByl1LH3P5F4
zZI4z7IdbgCJzJn/pmGwOVi3jcts5Gdgp9iyEq4FhSvyhd8aDjgIDv+ZhRY6R32t
FPaUPMRokVsVUwCgKy0UGSbeOf3ib4gce2oP/9MzkFJbtXOcNSUDxjnUuISlhacr
fEFqMQ3lgc7KG4fJnSy/EzAKy2XZokOFaE/HaY8BPjiLFNT2ocArw01N0CxP0gA5
UNhMBs78lLzBSTTpArxO3aTQQPUjIVALxuAnAfbHCDZo3/3Phi6px0QXBKRVStF7
FVqS6n6HptqYKva4ciUL0scJTAVl0CbZnmVPnzyROVjoOn86orlnX8Rj/eEgyeCu
SonT+M9ZbCJyOg90lRvhfEiIDEHtddDNO453H4nyNH+FB79urudf067kUn1yvBlo
CNBGzwx8JW6IBP1hR6DGzz/7CzaWun1U+3Bkugy9Y67+mU3vzgEhKJyUhz17iYlt
PByr5YjwwdB98BtWg0PbmlpdNRv2A/MfOQh5IO6aQ4OHt6PF0SPXGdQM/KOh8DHn
Ksz2l79IaE9a+XwYTR1StfXifkpCauLumeARHLWU7FcH0uyPhr8ieWtyEiJs/gDi
xtH6NeWQbsme5HSLUcmcc5m5CLvCd/cn6aUXpZ/z6L4scn1oZhU6GHFruENkTv2R
xsN3EF520uuUGb7wKiZEljSsai+7AGjxtm4iAQjrTORgY6rJzahfF1+bnCwHLE09
kau8ksidD8d52bUzgmc3swRng9+lwgNyRiv3KZmyTtqT8Lh4R9jZpplTea+xPx+f
cXxCikf2TMq2IdAOpFKrskzsBKa9MAF72+NM9g4RK7bGi8Z58S1Bv1okJX3zB1dS
L8T2cVd9FRwZZXd4b44O//fv6U2g6R10kwABMXeud01JT0+UpwJJ812QztytY+kB
eq0POCTNUOHnOvnnH2rDeE6/7x6+d92iXuFc3aBIKrb1HMAQ9brFZzKKAeZPvy5l
W4lZTCqspJUAlv3IdRLER1urE05JLtLtWNnQ/AmGlFZtx5vjflBjKgPra9K2dLnz
9aNIUk7cbyNdTlp2Br3PvotMu+a5NzrE/Gsfo2c6zUtjuQtd37/GDWyA+cdTOPa8
2PSiN6IH1ilzkhx+SqEjf1ywfu+FwgNucC3C8rz0S8LYx4MLQnoh2rz3LKoe+Jml
ITyNcHN8WBjEVJVQj/SXJzcp3MxMO9AqgupuxwqfL4PBQUO0jWHdf4V5MTWMxxQQ
TMfaHYOU6GaiYOFsdGlo852aKS/yA11R3QW9FZzea4jPTqcQBUgT/W8ERl4Ay5XR
XRP4fEvQwtBjYn7jF/N92cqHBccTky4WRGr2foHxyCXZXlf8VOijA4GIGv9xgL+D
LHRmCL9nXMol0XU5apATDfgZ1aK6wDVr3JIpwUJsuJu+P2RUcssWlv3iKWBuZpdl
NPW5sykirqPUClrlJx3kSPf1fAjp499IxO7bBVZ6nZsFuKHdDyN37WhTfnoEqNCI
4Ljapn72+k/HmiZaSGjSuyKtvGOd//c9SLrOLF8a39gFO6jCX887vxq2NW74ffRC
AHwFm/TcjmfchBCKUAqVNISTPwFUxh5OIPHqB8rqdzDXP3tc8EFETdVNZniCJqIT
fj4t3fhvDfA00y/U0O49moQ05TTYjJh7mqp2Ef2YITjzVVMjdv4+E29GByRRC6y2
K/BqVHBB2ziDUBfzix0w7/zRrfEjJAhcchwOklBhDbHEp7F1ypPqtP1EFdZCLvky
Wis6zYvLXJSIb+yN4lBejBABkUFF/XhyxvRNyHTr+86A/A6lIK/1dKFNan2tVoYd
rzarbyJKx3v3Q6KvWv89BL0xdtvWa495dzIBdVKn0oFZETQv5FCc1ysfgvzOUirj
WlR+74rUiZ+1CzcTHEUt7zgEeozcPpHrsLko530We/Jdcpm7oVE0k3DdQJgjvdXQ
76ZCIRScyqlmObFQ/aROgx5p2V6RjvEI8BhuftcudA9PfDHbDTjfJvnOojbCh2mC
MCn7N5qHl0Eaqv42gKmPNq9xlCnhdXf6GhXuHinKvndVXOR4AroqWXI4W2zROvOs
OVZ3b5M287qZNH5yPxK2LYR/QqSJ6jUKhwRJdVjFF8xZIvlGzZrKeZSfIpYHAdjO
O1zT3EeghjE/m+TDymNecdg2RxJkWMnclN1Yv2qxj1zH1Yvp2NRTdyxZgsLkNDAo
v4HmN36UcSqSRfwULMZ1H9LNq7/T1hDNXmTXoOgeOzjFSevZv++PkC9DTUsZnvgy
3GWYNHiRojyBAVe40r0F9wpz/2BBnCV0pFPazyifDDNmj+gQApPBVLx6ALuGeRC/
BdM6h0GoBaxqAIlYsW6ojwc+JN8uvy8MymRCt7voL0/UPCnortEv8Z7zD2kwr6is
CyTQKDC6LmUSfSpz91qRe17SGy+uNB8S3TiIBd3lM+1ivLtqQ1tiwoStPJY5+pTK
Wow8OCOJjIey4UeypwWQ0pDJynw5QhS+ZDmbE6VqWgXE07RZgdZjfaFFdBX8VFhh
AZDdah9VJM+dIWhd80Le+5IXsO0obdnHbHuvHdmK933SKeQJ+/LvXLyL0C6qkThp
WEjSk1gNssu275howddGcKoNJJhhkwdY0vFKUuM6JVinRNQuRj9qV1vULDaOqGAw
WEmT8Kf/i/rfGxeIaNRotUMyJwsoxI1uLDqVeroNL6/ekx75iC3WSdRmieiJ9S8P
uDxcc/NpXFx+LqN0718cH15L0EQngmdT4vmRIzWVgu0TMrt7L5RZ/+XLHTEIiYmG
cQUX0Ay42lxmmEWDvLkqqdifG86RhOQ25Q4NilBJ+OVmUB9Md151/s9/QpZ2PTHK
GF7yhF7flIzSLhT5hj049PqaImOfPExL+mND7i8BlBp35w3VB1LIjiapSx1RsnVE
Kzu4wWElXKxf0B0vzzyhf189vpWRmuPCE9oIk85wyULtvMKrn/ft1a12SbuteIm0
N+fVKiJH1X1ZP69DHa0uaKwZQsTtb7AyDH74LxY8PtvqqVAUFNy3CQGcCKd2orzt
slSxW/v7GTjj7IPsaIq9nnd3BRu91ExWMYUW48WXPOWkLSkyKJlBryJjmNyLkQzr
QO8ox4ZHYg5tjV6Af3tyt9lkJRR1CKAw1oY0ee9xa+Xf3QBd7zwGi6Y3iPZvNvJi
LKKn/6qTheXWh4z/xzDly7c8FQAhj9+eL6b8v2wdxq6Yx19PYL+e/17e0Ffq0ew6
Pwbmj8ZHVPN2WfLNPoX+uz8bBcrSQHVJ0nILhiKEeksFaERenBVK+hYYBdLHj4hN
FvF5Vd3vVRgyHc2UjXA9AX+nxMML9tFh3z73xYCBCiSHnV71czakDLSj7fQJaFdw
L3p3xTtEV77Jb3gRLrcpg6wNloDZ1fJBs5K2TVGf5aW+UunWzwDAPanL0ivlC7fE
czqwn1ZnlvfFmjAvHFAocD7eW1BPiXvYq/v/FrzCEmRsmEBxT9utpSZT/EMAwdLf
/owLOvaESmTR3v9U6LWBktYdV1y36uLTXQ2bfbkTMnJf7y4ATOsrMleVWg4ycfXe
EFP/yhY6vDOCelTEzLSTdcGfP3pfknuFwyz4ex1jNb8s3AZTu4HVNgB7iIIvFq8l
q+uSx4L/1mL8T67nfLHji012dbFQWufSgKvaebQ/Fxr3y4BZybb3NZ88t0cUP2Gz
zXWwDy+0AjLNgfalEvHWiD5uxMQJwU41yHWkBg0fnsElE9mP4y+pmT5BMXSfStrd
9GdPEt8NZmGudayddOeRW/eBak/1vQgKBzfAjcKDuD3kyJj87MlE5mMbLnGVasd7
uhxSTQ6Trv52u3MV7EL+EPjzbYDwdni2IHUMZzHoZR3ZJV+/OsttGn0dFvKlvlvL
0JJcYeRZpuMfBWxIGojIoFpis9GM/AG1hQ07kHe1/f71ZQlTAOOKiKGvE/s5MIX2
ItVNyFYymhqU+zi7MctudplxMmss7soToSy09DT9aEtigeUTJ6r8VQOWgI24wxE2
oEy8lsugnvohItsAsYzMLWtCmVwk5RJz7EIhoLpBOSd+n7kQwTnWhySL5WpYBg/+
w5iLFt0wc/QhvHfMD2kz9nO5fsQ1ffqUQSsBedSkR76np4mG42D4om2Azqe4KoUA
vWlji/jpzYEsbtXmoe93H+AqPreFYMljrLnxr8BZ/HoMXKh3Eb0R1n3bESbZ7463
8P2n1Wy/lGcNVRUUGrOX+z9Ct49nRVVBwfzcxHMqfnzm2QQVcpM19nQQKKAN2+lS
XZaTQVvT5xonfGpyjna2n+j0iyh1uX2yxZYy06N6hOenwoU6KiEzx4ThL4tlRtUK
4i5zTod+X4faqJBIylFGhYVio1FksIv8dLf6Jq226sSPZg50W5ytt0Vdu3XEm2u4
FpHvr8SD3EBqksiOR23Wldm147Pg0ibsn2hm+u2q4kgVNAt21DPevzWppKomEWui
sUh4/eQo5NhHfNZo5ASdsg0I8kDd9bst6+Gq3KVb9YBmWiHYeV3Tw8+tbBsRo4pe
Q6HhpWjJCFVa+Pf9IvO1fPHPsn8bFAEHQsmw2gouuB8unV8TI0ewrAZd/kRixGqx
BKDwmix9uAFtNM4Q5AxpJ7hd1PLok6/e2s39BoN/Ajnu+cEW0G0x8OcMGL36frVe
52OpxLxd8Iht0xR/vvUkFNlymGbtJYqfP1arn+oTKbMjHj3GQ4auLoSkyVWQuNYZ
Ypad+hEDZxTnd/X4C0CqqmIjNQj0BRE2aa9ioeAiIfBnAr5uSBNCjs9nxFODucMf
Cnjb03KxhKBp2uY4gM2wRtLZqSk5olP/sjGJf/3EkvXKEkkpgL6XhKbJvj1kfxeA
qoQCmvfkuyjeJ82vy6G+SUzSoXkCqHbL+yuecgUDufKeCZxnefGdofTVf7eNH+xE
sUU30vBtU1u3HeUuN899VJ3zy9ppCTVAH0IOAcyfw4dYZtCkNbsNf9aD56IK7+03
XBW8OTTH4U9R8EJP6cfhqVw2w6776SrFatadbDfxgj4WMTvqZr5BIBH3Txd3SJyf
uziD0SW6G3WffHRdWrpcfMOM3J/GHAvQmxFzHgNWSbIA3lyMpMLxN5PwN2id4oUZ
KbEFU84VOGSXWWsTlME0SYHdcx66AkN7jg+xfAV18cvJhMejDOcXaVOTeaQig0h1
r/4K3LHDfryGahJgVCtdZUO1wMUXewLftRXYKNyYQ+UxmjxEpyvWtkmRzhigkEWW
uBVwPhsVlpm4HDrWh4HjO3JH+WDNGW+ovihi1xYDqYhWGNIRmRc3t8RVcgTwv56s
Ri0605CGIoe0OgLK874vbldeU6Pdzusyul1wgT1opdQKhqbn9In024ap3Zif3VzD
/k/uIkSE3ETPzpNJOJ/zeH45GZAUsjDSIfSjVniFc4eaeZDSfY968fWIISCzh/wu
OeHeZjrj1+vpw5/OHfk+utupgcAal6TqhoX/o3elQMQnEMLtD3T8A4/b1MUrYwc0
2kPN3ieftdXrnlQDEbq5zxq5yefpiHR2jlmXlvRpa1mQJ+cPbAC6VBPRc3OJudLJ
gqSF8XGPjBKovmbc/UboZRKtDAe5Y+FK6HltMEGcS2HvePtWnuLrX/Qa42J1h1WZ
yUBKwEvVCIvfPlWw84ct2HF0RZNto1NTHqz+pcfGQ+zQug8IHx8ZP0e60Y/bhSF1
VhZ47dEn36DC7Blrc/QXx4yTrSfjXCHnu3HhfLFCo8w61YosYQV9MVNgnCsAuKDo
+Gzc3Bao5xvO6m/XFEWsA2HsB9lwpN4HiTUNDpK+B4acxNKW4WL07+kBh95BD9wf
C2f7vm9SAMtpQRH7EETePjqtgQ65mDegP/aPMS1xWp5emnjJvwdE8ozlnTJcFGN1
lf10NlM7E2EvvbgPP0duTpxsoKzV1w1ArHSgTBn8rmUFLYY4p85MPQSjlkzMZ2Ld
+KIL/tw/N5/qN2u29qJKXQ4iqhzO4m15NB/hAouGOKfsxYU6tZMs+7uF4Ja10tHh
ej9p5UXk0HnlIPs4AzZl0t6SKQX5L8oU7b+d3X4XB4OSOGCs3mb/qQHttKqXW8Yi
hOe7UMiEx89ofxTcfhEla4ZQv9s/zTWnEA9j3I2SCDxSqJo7OdRHihcAX/aEd3J2
on9JwsLmvQNMpDeI3ow0MSGCWsCyoKgjbJUAERoDHcoTW3eAvsLXn5VAvPNsMk7q
cW8tr4n4sxpIWecynJ8knyHRA+n0WmQhQxYIZl5aWqm8MefjFgCMr3dnwGPPrl0W
UwUT1PncpZYJwbwPu8lYqapM7eYge6Audy7/WB+8N6sK1ZIFSxDM+7bChpN/rdog
1Bff5l87648EAxKqO6xVfl114WetAGziupKF8saNXuqFoTwzwIBFv4/fa+ZFYHfP
hrtk0fwPx8aVRb5bKFHnnS4iKhzr6tHGpP/r8e/gI5ovLZ1mS8+urrB/jEKxi6nX
CW9gux7ZCo6g11LS9ltlAdHfr+S1YxjP3Xk+zb+DnPSPDYcUtAJqq1HLzf/IjQDh
tIePN8ew0My5MTBn/sGsvxxFNK+cEfMirUnxFGM//SLqEB/IXik6z87/+1PPVQ4S
6YNlk+kAhjN7Ns3O3BJS7MCPaJmGfbDxA0tDzLEvTlxZv6z9A1Khg5lIbfyH5LM0
P63tKDj1jwydc576zGcnLB+WGPiJbCz06oRi/8BiEWEobHEKcS6taeJ+ZXbChvlq
0K0JhOkXSGSwXaaXLqN/tuMY3ggy1KPU3EcpPZn5rhC3bZF17tWUbixzRCgQ2XwR
ffl32LYt7daBjmo5/Rq0rVa6yU9NlMOPMx2pew/O79Bms9BinFeMlyuNDeDTp7RJ
uz9ZptYMxmY5IzaAytUWKtWuwvdzX1kMIgBfUbQfGkTzwsSWtUFBuynKJAqX9Pr4
TuBvk4GXVpwpLStD6GQW1pWRJnW4hT18q3dYToGYnPrmJW7JPlVS+tCjnBaGs7Yr
vQ654BcLEwxq38oT3chUmPk4/GxSdOXHlzbN8c0q7E3f3fgGFEzkMco5fETv07FM
j+O45+1klhdyNJ0WU/oDWD43/bdrtI/RyI0AjGdpwdimgBN4O0P84ffBHDbXkOq0
DNPlkWOmRwTvTfHUXTr8JFvoCZZ+zbr0duBdttdFyVHVfNCVwhwj071kpZZeiZU5
nowJfr63HIfhwgVoQTkiBDd+wTYVvDo4pKaRs+tw4Zohrkk7omOQb0SQq0jjIgUn
DmSuB884T7bryhxWKYzPIxxxnsYZbuWBl1uNHELu8RSzz7zg9aEJlMVVBm0NqYeH
cIfJSPVx9/tV1cMaOKx4vu7HsbDJ6FH2+0ZQKdN+oGsaHFlx0U1M9wxw+pRudMpd
o3gcF7Y4tFzek2zY4HQJgnIh6PnRhAXHHzPbFiBd/E4u8abrPgC/afC2dSC3jUTi
VVY/FOeQArk/JgPdt4IYc2CfNgQdbnKnEcPcxQnvU7/Slke+kr9KSyuadcqL4+/c
XwrHSd2eGodGlErnqEfqYx2dmP+Z79MQuLILIO6D6Yv5j4jFfO6rQahDZISNXT97
xFqjWkUuJjmJbnrVMMsB+e79AnKs/bYqG2TsMU/E+J5atA2MfKDDp2GbZoD+Vgkn
PHQhiuSxJq/hXsFfkZnmPVhSK0tpFrJGod+h8CHhukhu11ZrZwf3w3v2I8LA/8oj
4egrhZ/haeAKcCFviaSBTnUFOT8ThYWS7E+V92qPv54HPZcznSalGkhrnA4EDUVR
gtYZokH7mu9gzaVDoKwzl4z7fd5ZM8Pny5quSbgzxbRdtgx8aSxCZFrVCdEAJLa8
UT7JD+1AeGRtYZZwqHvmQkp8x8gYksZ14oL6BlAHao911E831ekU7N8kkwpRA7Gh
6XVQUW3VDoff1baluE6TRThOZCBsgbSDJGT9cxOgLGxAVxVNWMiJNLam6yh9Mc2J
Cd0PGQHlpv7VbN+Y1vt8MPxKpOSlMfrR2skfGkWTuF0G4D4nLQKBhyHoSgG5h0M2
Ykg36keyxJ8H0oNHJu+aIkxN9ti8huyVpSoybwyw/8RlzQK9qsDBvD1x/ECb4kq7
MME8QtPQS9EddELp2oz3jfsAQnVYSZabdaKaS8NWWC//B0kDrfhZfsUMrgTqbOot
JOBtqsYvSkvVjdj5rYYS9M2nBZJLv/k97gVJMAy1HlLU5A384nG5+1ZaeI/nR+zw
IV525fvhacYG4/T8CzgEA+s/bM/iT+ZbnKmIiZrGfGnRqjNGZfL4m/xpL4Rp388p
LdkGVdCLQNOmQKjRMqbqJ6L04UNIPW6b5mASeA0Hm92copVi5doTHkNeBENJBivZ
K1zKER8llSzDJOrmtnpNcclX7JxSYyVv8MYvWHzCX3t5xYPx9icqzi9l0SjRbg+L
nlNaJXLwW3BSY4ycGQSntaW7Wz2VRQpKRTBzeCzUhny60cUQEG8klakAbTwPOZHB
Da7oiT0iONoiUEb2xfsFdW1Eiy3dxVBChpUm6ZYfAeMC/ff41ffvgc7vEoilieIi
bOw3SaWhRKHk4GgwfmjGetYo958C3aJBmgBYmuB7894HAXiXTNpqj6YGSO2s4YJK
WTCiUnq41iCNzj5FOn4Ha8G23rEGN/OhIJkstgEB6y9iDuJEGRWermBBRNeEVLmp
iat0hZJY93AB39LkRjBu21I2Wzp/QXasNeMCzCW53H6lZgg8bZmqar5zWwBx/SVg
ncg9HOTmQZV8JAJjXlvsDWxoqLQldf4V5IjUzpK5Sgum61iFi5ikDUCv146WeA77
3ZuV7Sn7VaIRNmAdCH0VLCJkhz+m/ZVea+i2lwIY4lWDn1qvjN3AtP6vQcI/PC7X
iyDgdgpc1g3ZNPu43k4YxzIep8KrC2b4wtEDS02lVjKb2MnelONlCjWR1aQzpJkm
KNR5Q03o1fjNHImPxNMwjGJwEkz5yZ+DdLUZQ9Ehv3No2DshGvr9v4ZuF5cSGgqC
O+TwEqVQt88RWTHLzftKyT00+zSiJ+z39jVDjhtheJoazP8f5usi9q/Mum/w37TK
S6rH39eNJlEA1taGG1HVjQ+A5tgPGcDlEYViKOzADGOMMORsXnOlvP+/g/H67wrY
criN7J3eCqeaMeLJ7siTR1m+VgaLYD2SITgPEfKQ18dkYhQVjnlyIpY0z/NiVWac
HgrP3wTfvNFpy5FSgu4V2kO7TasHLa19gkHcznT6g8q+Ofshl69XGmNALUj8nNEe
gwd2zzzvroKZt+6AbFq8mM0/CH5BICX1MOkFMBpmXIzLlrkVzUpaWhHnErMpf9Hy
3OqJ64OkxrmbghCAZZplRdCmgrf61ExLFY3CPwQ9LWVCf5M3ycB2sTgkkEhEFd1M
4wG2aDd5hgjql3GrhLTeuvCfHYyVcEk9ljo7L3SLXp74u3Hh5TKM84K1xLTqh7+m
hZy3VU33Df7QRGx7PVECzCCjiwa40YlVd0sFpFEwVYk/OUJBvfDWYY8G3TXw5oKI
88Wbb+3/tohUWrz0AK7A5t93lpKNq4OSgIzNAE0a2OoEhYpYhICyXCJ4BG0MKzix
liTeGxTHuYqsIjQdhvcx3qWCGmrtWv1C0i8Umg/wRzT+mO0B/wyM30pDFG3yplpX
DLZeEhXVoqSWSQj3JwQ7DyFr9IMu+I+FHrf2tScVJx5rOZthS+gKXrW+4CdhgN+D
4k/Y0rpxD68TraK6XtXFTuDPJMQ1n0OfCa8us0BfpXcmepCpipI3AvXPqqcTTmhX
qfkkSRvYqLzgcUQVM7OLHsHwi8q9OszqVv/tdAy7X6NhgDb/m4ZWNYuksiaHAzTS
O49dbeyPDbolWCkNN/UMOcvCITNMcBszSCX4ea+Sciqhf4kW9PU2QY03QR3fIIoz
+n//bS5BBPBc5DJcPcE8F7YsYlvP+uozv0o1XNeOvGa3xD7WHdKeoRRfObQ8VJju
KsAv6QHYR+GrvASo1vevzy5DEtwDs9qX3+wxAXX02fFsS5RiLjMQNwNUYQMMZUrU
iHC2W1cbfLuFchy2YOMz55rI0sfKQbahvfTObRwoJwuI6nzHURKaNpaJ/n1y040v
Bkvq+/QrXSQtIr4x5fT2r5js0OVaV90Ig75dWfccKgnAjbEiDT3q+IA9Q7tsrNB+
a7n8Zzve+pHos0FwmLAfC+BVBNZVJKa8naTGYJnbqWShKTxlAQa+dqlLXoNSiNoo
yVAlEL+4Gvzbi5vDyK1DaDr5E9ShAYVFwiV5Srxi82TmdmbV4zPYHotsxOiMpgCo
OR68spiJZa15RsrDkqI2zO1TQHtZgrpt28ixJPmc6YaNnQ6jCOtM1jPy3Ikmsf0U
z6fNvLVXT7oImzCzxVVuoH54kpD+pweernzJP+MgFV8n86wzJX6dwn+8f9dk5AJn
aRPPoiqHlZdTJQjVGsqG5NBk6IqmT/Q81mxy32oLmitxFQG+IfvpyPQDjEZjI18f
frmSMKsg3cYa1CzNuYzaoGdT/lY+S/6S6qi/0Mf8SG7WfSI65UZcoEoozd1BhYuR
YqrGQKXqyGaJFJyMZRsepzEDwTRlJ86TpenxNfRrh9d1RZ5dhjslOzeTP1ECOBdJ
RtO9o0NGhc1fc5Ktqp/G/rQiNDqt3Gad4rrDrzYKwHUolhGvZ0XPe1npT/2THj6Y
RCWinkVtLg5aAVCC46BlZ7gm0BOvTBVvnpf37BCMwYT3rxeEQjPgsfDhkQxgkvW8
fpJkJU6KcP3TCeQfrlBHJHsB4FOQGrYZH/pcBNTKzv8COpNUiRaKY4iKTW7ppn+s
CmRrGmfLHq6VEq31VmeiXqGWKI+qK8cTCGEurR0pvKbT7lXWWXhs5LPhrv/60Idb
U8FLz0XCDsb6Ey1ZtHC3FefvK95ZTI1+PseK4VtCUQs094DDEb9utxSshOZ5QoeU
I2mF/mXXpf9o7GsPiVK4/kK4k2jEtcmI551aMrLHcbdBXCHTsu+VtZmy/YA3uDMM
GX9kM6MKk24dwTywFDIPO389S20XHYWy5umMOZN8Oe7JhtMOvSDw+0JVJ1XDxPCd
gTVk40m00fZY22qTMhLTe2nKZIKU2fuq7AHG99izshIGbtgVULzxXW+WByb7Mlsn
kJcOM6gwSg554OTq2qYT5rg6O4X1GhUFjAsl9dxeEC0+pJSxmFLYmYqUdyh90vBv
BnXxq6esqLeHJ6DnFtxT81fw81GU2DMs2P3fCvbYtRringrjuYwGojXYRUOXKqg6
9vrgtrJXWQRWkeCqAsXUq8zpkqYtRLdlKAgOJqX5ILhiMsrJEdl93aP+1tJJFdHL
iejjeOc/faLUcGyvlRZvsykjo27KdReZvtfzkHmfO/a4PHXcUDN8T7JySyHP17gH
oWM9+OWdAt4GwANYbHa+zQASQxHBf6D7iTppIJVVquL5MGsPVxUd88SMecmNIOQw
bHbTOii9IlyE/YPaHZLaXQezdj/yJspZOf2XG15mgDfAk+RakAFgps3tU2ANdlK2
/c6smUbMPDf4B1pg74YdTomjkEiGB1zFJWa/Jpynq8PYdAsmm+i1CnMntaH0Wl3J
p86N7X56F/id/C4KXGsKijtP8G99D0Bnuap1MvdYaytxfsgqooGszC5n+D/l237y
R6S7gGXPO3SmPgmulAeR7XlAqll+w328ADd422D7CSZBWvPig9WukKlpwpsw7FpY
A3CiO4Ni8eL8poWPCV2cscyzfQD2x+NJ80INmrB9gXvQ4h0/ORagtXNZO5EDI8yG
T3GVJnPxjuy/jwqybYpnkDsd564o/V8IIzKyMitaEmASAyBlz2t8CjM5/zYRd0mw
73bAkMJn4rwyJaZxuUgEUb00qVyscYn005T2G1u3+a1jWpMUf+eHXFrQozWLa7A1
525CevZuKau1Aggxt0Cjuo7aA3Iuq7HdAe4bNSLqqq0ohRgxn+QXjIK2h49SUl6O
C67dTibbRxe1MUnaLyWHngM6cD+8crDpZhxBccgulBKd1Gyp23m9uqEpb1gkmDUw
tZsvnoL8ezEx7EHZLUEdKR1Zn1iHUq+38vfRZI0g0hjHDrFv3Y+S6TPyWQOjBwoq
4Tks+Iz8jodNJODJc3RHLG1enzBmWNvRrbEG4c6t3q54vsFqIAvxn6KN4eyhdS5j
i9KmMpC2Xhb43qqb5aVQmHHzjYM7oGOspnnyzrR1hCncLICpPvHcHS7zRjzbv6Xe
YonVsDLFfzW9kymZKl0hadygPUjxj+cInXoyOYnCgJTpwBXWWFRR8uwF1X8J/j6K
CRb01pj9wxWbCXURNKFV3kAaWZoRMay2IR7saBYs6reU2GbBLj2obACRPhQeKYIc
idzrQPAoMAlz5A2AMKYLpx4FMqGzqH5OjbtKZacvIfnEPGO1auWjG5PNPC3cVCYF
Nl0Q+nuwpCs98KLWwsRdjMxUXNa3hNPSds4RUezBjAaCacvBeUPfX8+EbFei2DKE
LsLDVWOD4SfH8mdjvkneFifyZKHA9Ltk60CKUhAbzQs5pAwSzyV+C/gmP8BLVQGV
uYm7sZ4FSbaWkkIoOYwoYveBM+ET6QlPArHnzXjcuKGS7KrUZAzlf44PifxMGwqm
/sXK+QSLZ8Y2ZlQnEdNu0bhm7uprs+Ys6/1ir1GlIIK1SspCZOp7o0Dkg0oC3F/Y
Rb4osYmN98iG3gxreUFEAknRLgci/9MphScDuXfV680RHzp/jZfhwK85NWhQMG+7
MdUsixgdWEHHlq1WhwRQ5xIoAFDx1YZ2LQ9jr/mwkcUus9WnHjuSl4+ep8NetPXp
/R5EnftsptjVjnr4fnFUCOHaRQigkGdifwjQLJz34Lk95KxVX8neoqFXm0Sf2kmO
S+91IP/J9igUYKBRhIK6EjRqjto8//kikMS+igNmDpg951Gh6tK6YqAGUYbNwlQv
esAg7W2ZnJCX067FT1Y0V1KWFQ50YXcSswHEdeaJtnl1LpxOcAW4t/OGqFxJJqsq
Dj6o95pbv0wyZmpg7H2zv7kGUVrrM1+K005i5BEjT+wORxUlqEmOZCcqMKzf/rpf
uZria2Yyjir0rPgS17fAMFBbpepwhAhg3AhlLPos4+vMEQJMInVnX3DT+qF7695J
+Yh8BSuZXDD9lfVggUYGG09SwTYtqu7V1Y3Hh9M74ICsPMnaRlI/kxbc1XkpNG2b
rDaoaSkuZo2HrYu124weQkZDcMEhju2CAJx5jhtmhv+VFzgdnyELeviyGbbQrZBJ
1hvC2FwixpqdaWX+d8nbl/Bcv3LpqXXQDw6gxniO5PQ11zdzcI3i/OvGt0JNXu8q
pYds7B/+b2kAXseAll4TAM9f7bvtOMwcM018mXP8OCz0/rwx4niIMgGcMuJoEUeh
NEFabaiMu7lG4wdYzCnDFX7nNo+GtbGRD96DI99xkW0oMrMTVoxt1y9TlT7I32yG
ifWzl5vaVqCromPNO1Z7ZLVEdDu8L/bzKd7j0AENKWZprYEpnoY3UwHyiU+EzCBg
6GO5UkufL+O1Qun0dBJzslw/hFggkw2O2TXsexmgL+vtnZOtY5I2uv8guOtY7y1+
r9+cWHy58ESq4ynUsb1J6yLK1c04DAG4icysKBlbuvyaPrft+upxdXTvMaV2yogY
0vXZIa6J/pLDh50wNbVHcJ/J6Sd4lqnHHeOO57cP8camJaD/0e4qaaYsODB6WpzU
vpwewWqTSzdxF93cgm+mO5vvUwaq4joerzZl90jIZDkccaOrDAbe/pyC8MKnBPOs
2IgSTPKhkxafyfNthvqddXTqJW/p7Biz1BgaKpanaOWriXbYIWLTMa+6ajghl3Jj
lwqPleol8obTEy+Nn6KesrgJpav6PCA4cLKRWldsTEM7DL1RDLWDw4lHT68MGjxd
a8sEqxNymeQ2VdWxOZjp7Df+odLdCIWtCYJdRwnISFnmZivc6eUDdOWjFlEUqj8i
L4Pzg1sUTTtiXVwMloa7aPVlZWvGmZzGk0rYBrLPEB1GBdXRJk7r1fy31Xj9ROcZ
KFC6V/Yg2ChlNGGmk21rX3+z2dHjpkdAcSTvyL0dI+6U7/z418ES60PXGtY6OQCW
oV+TJb8bpxP3ZV1dIvH0q4j7ab3moYix1vyHO8lG6dblGlCkzZbFiLcfBlR25ZZx
DzSj37Up2eNnSr333/IFVepQnCtSKp/WKZHT/CLW1ie0os6YIUCMssBbf4yXyvkf
imPFZ5chWA/Sye1kXemq7G02m8dQDF3gs77gYmpL2R1MTmr04YsULbAYc34EP8wY
LtQEsqGjFhZF00pFHkq0IH97r3lyvDCNzk7MpzekLRA3gv+1bG/nrA+8PSoubf+H
PNblZpCr3jNMpc0jP+nnwnZFKuR3khK/cZoMd332HHR31QU0PFq4j6LZWuvySoTn
3u76pVxLC/ipL6fv82gE2ztsXmfyBZBDBrhj8edeqU2GhhcbBUjPb1cvGBYvmWPc
lp9K/yq8Et9XBb76LOtqlc3i5CVDm30OhnTR6uaScRkLEVMCkS8kc7S70Iy8kCZX
ooEJl2jjWNfCntkVdMI2g3QJsMWohmk/YClEQLKq04Qs+wcMOpthd8n/sd1RSUOc
g45NYs2sZGbUZLuZ+MqhMXCeMtN82DqsstQKDPiRmajWbS2+IphxPfq8OLv8Hjk5
QksgtKX9dX6dwDtKdSGA4mvE9+dMYzKX7+PDkdhini9zALyKT+oxazhlDHFWXh+Z
j8ZgcVHch7yZ4bI/LelgnOgtuFevvKlxGry7/Vy+gKuXga/zQkIhQkCLc2WVR4O4
Vl07ah836l2z2dcd8PoZqRdtQi4VnfzGxXWR90alkLVRtNd8UmrlhQEEIgONm51B
mhCzjwuKFfabBW3eqSZYqskKJGsrBqAs+Xi1jRXrHSGA3h4xGFdCKlIiP+jvRRzP
5i3sZDH0QaT4RLupRibJMDMFKJ2YdwiK6i1w6mFmnbkva/5XUVuVL+jvzhBnQ0Vx
80FwNs3hn88V2X8tofV2mI+IpmbX6uoos9BScBp5335XXUaTdf0IMnSbqfVWCm0o
O0lU39H7JuifU/A95j6pIoSpWpBKkHWfvvNlTORsLiP2XOCgemjYIjUQsyYwnp4Q
VrNxYsdG0J5vpS3VTMBcUd8X6mTAccKT2xnk/8qvlW5VeMNd5hHG5EZbBotfZLE8
jIbOjguPh7dTUhkOXXph5pt6FZn4PxLKUgXRiPEcD8zKyMi49lBMBORCWne5tc64
d4eWWjrZ3VWW0gNodRg1aTd9J/2tO/ODzvmiL0U3gE0wClhv+oFI9wmEa55T/Zt+
BFGz29wQPsKRQOwbWUq52ay4uVl7Xa24/kAfSg5AacVOxMm+pZhFnODcGzv2r8O1
cvpFaKHtGgVtuN4YucDJsy81t7GIE+WgcTMIqY/vJ1QBPkMYCP8lcQCLE25XDPs8
tV/n9arcxBZOJCQP/M6FkUwcKb8ZiI3RE1Zzff1bbnroi9vw9xxHRP4enyCR632j
K7XmJ9dcp81paeXO4KvEWVHirepvuLnk1DUTDQE3MJ4rJ4riviMVXeVoG9tkGgu8
/R8jDLGocbbWocTe9fL6MJQ0hJJ5th40tv3WpK8TmHFG/CzIIN+4GsLMrV1JT7ts
v3/QzRio6ndZLHGovICt9uYs7nMbSfFSIjYTcsghZVgcqVZJ2CBuSzEgDGGBTzW/
3fukrmDY09amTCNAd2CRyh3+NZI6cEbBbWSnbz98a7X5q3tv9W0vm41/Fpg3wGJd
MBn28Au7csKt2b0Yvi26OjW9gWL8aWLgnO9rpE2qSqiNokT7eee5X02qthVuM2YH
6AS7NDj8Rg5WviZufuBYzJA2o+RyYjeBeK0yLnEKIQ7E8WiO7invgeef4VpNrJMz
3BLP5PrhzFCq5GVIpSaaTQ43KfsAVj44R1LOo2Yx1Xao24aS4KAbpXquiovcvAef
psR772sA0JWI4HuZIRwIHJHxt+SE5owbfCddRHwR8gvYW3tYrZZE7JdOqpBUubjI
ZkVcrL4j+/6kH1dZe+GHHLxOwSug4OuuUITbLkIAgymmVJehHLxSdhuIGnORUNzw
rFb3UJclORbEVMRYIiQLAzP5SuSgu/Taz0zqlP38/80CQ51AcloNGXpAyZAj9b18
+IqGf4TBJZCOb5xhWvula7lApfD565Jwty+gkV3svWvZtWb+FyqOUNVkiB3cFRZt
EQsU35vGuPd35oBS2hI+BEc9B7ZuPpICHIXD6acrSarT+D+bHUDXvPIea4qLFkIs
D7OkH4FSttkC4ggABGta3MIVM+FVFlnjESWv1dqKa23rxOuUh/vn0qCIkN+yflRY
zhL5blV+8lJxNuKXnP7FFQsJhHd9+Ia3SqHjsHGE78ALivTWORhC6+So1PPUdQ6b
xG58mdQkrKOCp7bKKJ3CVPwnnm0u/OiY6nqAx2thvKiOwzJjDZTbWaICoXo8jz6Z
r6bacv/dsv5aGGeZpyILdT1PQUx0GVT4DPnSTBE1u6Z/+Bb4KktszuQjzGPnOeMz
CofqqZceZzX5NSsSuSd/Xn9yYXFzpDqFmgwojiWL5gFuSnt1XcgKDg9kkXTH12bF
9f0mhNcKQ+1Gu1JomN8kMqnbiWjjqVES6lhio+tfwR+SaTH4CPHbKflU6RDRQtbz
7rfYbn0bldnqxDU0eQ8cfqzgn8GLRPiOBwMziVzWmZSO8kfawBpJOPqj9yYOilfb
mKtCjyYSaNVYPNuV25OcnFc7oWv8R3tvKssAuP4/U1Emyr7Wyrk8fNwOeX8uTIm0
dPxI80NTVWvb/+Esf2DFk9MM/3r8NCZEIEkG1B59fN8OB6rTbG+ajnzpLRkCVHt5
35inpgwqOtpRqULk9C1GV9Lpk0p81BbWjRs/syzbygFfOJToD5JfcQ4dK79K5Odk
/MtpRPVaiG91DZxJnHtINFiSAOcEPYoqKzYxrjUk3GCd27BRPp3ej2Wly8n4K/BR
7VWPn0QOdNh+mzkhm4hhRKe2Ilx4+SgcsqcmmG2e0XQZ6C39GMNG8h1MaEOmqXcY
1Xyfv5JllYi5mSlR3Y6TihquMu3QOck+ZUq5IxOwsC65Ylq8LNPrUq7FwY8sn1o/
OjvZ3b2ixozmJy6cDBOuc4iko0Emo9LB1TV6qsGc8BPybd95GjZ8U4NbynIhnE7P
JX2FWG7A1teKyUOYVV23H615aTEHxkr/Kr+n4t702TanxtoobsiLUJjA+zDxHlDc
f5xukcJIVTfVfJse+BZUiNtQy0K2zuzpPtKuLjoyeactRuxed4l/OTI2cZY769Dd
GsSI7gqUbxuvhf+Xs6S5D/ig0WMarcpuXvgiAIfBIcO3eO/ctAURyfPXac+1FMlP
51dgKfVmfB47L5PVjnhVTJ+xh2zm94zMnVMGTL3Mpc76FRaoMVnF2qehyJVvKv3Y
oSOh8CNQIJz3089YYPDZe11Cjb2W2pXLOFxtLHEvFJ4dzSXm+29J56rK8pJW8jkF
olsNaN+D7S1ClBt8rZKgMOGljLyp7gXl9BFWngsB8UF6x0uRP+GZg/vQWLhjQR1d
hKqcDCEFoODnvkIbF1/3IR6Uk/+BTTWdzaeU6xDqFrv7EcrvdaSpHyqu+RqCUV+A
Euze5WrqXwORellJtXIkKoJxZMWxlZIRiS0GZeJYOApqjsiyZpZFm73RwfUS7Jtd
9JlqIDcUVMOseBuBvNjRdEBJap7Pdj9XogRNqj/QJLzMQHj464LkD6caSFf5OlHB
xxQvSoRtwms3mGWs1pbkSVZO9ts5mIiqYLOAun+kDp9E68w04NF6c32vJ7/6BCBo
HN6mYqbtWl6gPaLKdryqcmSQ7cr/ZjtXbmZY5rOk5UHIf4eqwwWOkq69Ia6ruuiw
zCmvDXO6+neVZI5Uf4MMyS+H1WiJeZdUfJ9ffmmBNQ7LKdqKWYmslAv02/11eVtP
kNvDUYMMBnaxXezB4RHtTBTs2cMMeRt6fEIBqXdMLQ56CHt/DvtFnf2nITeBdOmx
OSmjGUB0Y9iIByXCxFA+3PnK1w/uKy7GRYIFt6qmM1/N41t53681XeHYZqbJ+LiC
z1zkerG848MYI5vzxLM1WzMcseNvrX5wAnE4/QbFrAzeyk8HHLNlXPxySHPkZ66X
xS6kachbhFY+XupzRt7Q+byW9b2FGpVGpwOItt5qzMGbDRVaWIe6VUWCzat/r6cw
d/FWDsujSwUGlj+485r8O73mqdOoJNxZ5k/WSnsXvIyNgIMVeom6sTK6Jw11t8SE
Tvw1uonfNEZNyD996ybWWWNalooO5relOwz6GPxnrl5h+fEppgl4IDYPRObgIgvL
IpPXVu06JtgdA+yXdxvbHwUVLfci45gH7vXdIgHUP2bV6u2glauHgaKZsvYqA4tR
xcLElzeHe528ULtmYs71tSB7oaGOCwk/cOo9DHWWaS1FBGqgN/Ji3NbGqD2zKoK+
B3miD08t2cTsDuHWAbu7EhzFcCgHfKGfoVlSIEJyJcpgVhpcogPlQM7s/xqbHRwc
7lvr31ZPTDXFM8mzYvxLi1udl14A3MBzzHUZ3jlWSF/jMxiYkbHDk2eCIOG5OCnn
f1R/Q8/2cJrAIRRelXsGJyOspeVZWXBodwtl/2kd5ZSry+kXgTpmFasPmqoy2H9n
1vVsgwLpwBPytXBEaytpjyLxzDTU2IpYae5zw2vND62JmjIWJAOt5mFau4jHoXYm
0sADDk46W+OIMRlZz3HJukE6zNz+NpeSvTAqI5J/nDyPLHRHNV0zj7Btq432WyMP
B5D+Fmy1Gpodq2tBL5LNg+ziByvAKihWTNhoqOPOvzNJelmTvq02yweWg4wigOwd
A429Bw/snnnPbdrPsXeFQuRrZm7K/iJBd5VMNSlj7fkGKJNGHB723D6+TgYsCfWz
xVK9S9KB4wVxKdCNVg8USCIQ2J7PcaKScQfr8TH++XG1Z9ap3c6046wF48kyXRfz
dIZ0eoyMHEaBWWa+SaZZX7Rk9Wolydc5buP4jnQ6UelAJfkN2LK54CoSoJtpnfD3
AuUY+PoRQkM9Gyaj0LQlxob8ZgNUjomQ26S5zfqFQBw2FmJVs2xx3tfJURU86vO3
RVcmJJdh3cafIKl6IdBMEE+XRg6G3M4y4lWj3c5TFLmn0LKHmL/2v/EB9CwxiWLr
6llIrcyDp5Vc5eBJSM5cePv9IihwU6Zw+9lZIxJQycIYiv2x8WD7skzZ0G6/9BRL
BPSgeKT6lLuXsMpJO9LKCKnPaipur6BAjPx+938+tzdhkxR4T0OhPNzZk1MazpeE
EPRVQB3lNzTWWhRjiyi81QT5AZsheCPq9kGyMXyuxCdeMAE+2G/LvLM+gR/ZBPWf
OSgdSHOnICaKIOuVPFl8/3ClkymtYBXgTElce/2GrMRiSHOGUT+IMKDxQiwTMdeG
31z3J4stga70Y+qqQ+ZfEMrKLtC9vMOw+yP9lDM87tgJQduHqVHmo0waCoWNhUYN
zDFICztZ3JobNIpaeK7P7aBVOVxgoVYa3Es6LxLgzKe2PsrTYQlp/wXv7V/8heZq
FBJtsRShZVWPmeuQjKf0zs5BRNFdxOLgB4DTbi6p7KFfT/9ySN9oGbo2O2xvZe/M
bvKwr/wOzIjt3F5PPNfHMZ5RrWLZtCIj3R3Ql4An0kfZUHdHVrGyQFnWdygMFRuJ
6mCWM0HCCjBo+jMZVMTUQik++ukrLHDZkuc178vk6dmWIYtjDRsW/tFpMHjLZZ02
1FR+QE+p4ufzXPICAK6JRBq0MgOj00Ux0cZxTW0Rw4nwnRrdRp9fQpxQkt7q/vvV
wP8RLeJnHkDJraswluCJImn5BPN5Eo7Pz83XqnSDoxWNG9nxCuZEpsI1Y/V6GUBL
XP9BrtdUBYINjh9yg53widlClns4/1mSh3JZfaV/ot8uBG357RpKgAXaX0C+IvRK
e0ChKlepf+0RvxWUjRkBvnog+Mlrw1LapSgImfrqFrcXwjhsVqLeo9NZaM4XBGrQ
cEi3LqqdbcKUWL9zizx/JoATLhBBcSWSBEVi03kLfHP7SoFA8r5u5As7I5zk31xJ
bIsK94ONuzRejCU2ZFTlXTT2yBJy6MKd5r+AV6Jwxn5aTjH9jisLmvTnn2UJebAu
1Ts/JPEwhP/cscQ9z6Fe3lCUHxcbBkNUhCxfZ/SA1aVH+khA8pMVQvldEilNVi+U
XQF9P1Sqz4a1XkFrhuxKsyQaftIOEInu3O4Twp/rHpoFX0vIeKHymTLL54vaVesm
fOQCI5Hc1Y1X+JEwWfAyqJCqodIiN2iIv74C4ZO+0KRw0mun+4zwL/iYkVWFGWfQ
JWMWz8ngQ5HAK2O3Op8dhr/dpl1GxsEoT2Dmwj+Dyf/aCMOeK4vhooFWGRq10wBn
pVx0rCSY4mjEHMyqVSFKWoC6LqjYuJoI+053vcucN2n+D/h6oOOBqCcMD0cLsUvG
X8bRcrSraNIjZbHiyi+o4th8LMfXHe+3V47AZZJY37mRTQSSFIPe95zOeCXYEeb7
tTxOSP7MGzV5JYM1KxTtfUu81+Zn5CyvhLLg3bP3kwTFe/Jqd2Wcm7Kb581iLj05
gPH+0PFjjcv31CoO9S6n5er10n4ynORD3r4PCW6uboKSw6cfMdKBll+bnZWeVeaL
evSFAK0NnKZWqrGm2h1LEdRonhBctjEqaWcXjg3fGctZL9Xj5LhEFnae5n/uZyid
cgMdRTB8BhZvXJ+Mh2CicZhosCz2tjKRdfaPOMFzaN6GKj5XM9tYh/xlefyC4UIe
31iL+fYB6pXYvGW5fywXzN72rzBKVzvao9PXnc4+IpF7Jf88h9YTJW+28YfrrMNU
9UzA8rhoEJhrJf+yGRedyJZUxDSTa7j9J9oG8/1DvLGk+BZGEYm+sQ+3NLTJJg2+
+hb86I61k+zpWddNAV+LpOhPvDsHFvKoAD8NP3zTT07JW8rbuZHlM9yeHqHfKB+Y
Bk+XCDpkDTHNk6bqGqJWThhKUYhnHQYKgOYtcyVPjJTOJuBQoHT6BxzXT8wDuDHl
HoFPi7Cfs6Be4M6mlsU/UZy9ed8JJohoLGbl35YsePCQu2P44xxKbtGtr8R9n9Jr
JuCXhiviQchQg4hnUX7yCkyvNjuf1qq4zw6lW7ERR9Yp0O5sblMTfNNTrTITdkkj
xrxkAeN/fLg1TrvasbW+3bsdYHHpcCMoISKo8n47T6Dl6J6MWptTWjzJ2SRIThlM
4J/KERauw2mezkgCm5f4RW1gyZmIZrOUrbzJax7rYRo1GiGISebu14akkxByw9Av
C+maiq+ASEN6lHbf6Yr4UGMDm2EaHMKX6WdcQynZm4UB+hB56l2hBlrYtbmBktbW
lMXOb2mIocVvBQbAKzarRuw/7G+jgWVoqXrPd8fwnsx3nCThdtJYrW/5r1nCrFSX
hQCKVtWdDfm+Xde/9VJsZdwhzWg5vW5ILq4P8luJv2N/Q4REJJqUXllDhZVoAPr6
thq1Om34Lk9rJuk/HLm8thOwaPIfN762/Y1ZbdxdU7aUHrgleP4PsInrUrJMjzoV
c0cJWmocIOaI5Kl5ZTsBIWi5enOf1ViG3ztPZnYSqBvrkh8l7CaiubpliefQy++U
nejDa7qmRlq5qlXyOGXgfjWBZ3K6BGCTAIxBlg0abh/1oQa3PmcbKNB6nllMoJ8t
iQKSu3ACLt9I0NpRoGk+FodtrNiLyO7r6vDpA1oHWqQLHaMo9T/We8KMBryXwxuF
fhXYm40jyhOfG1KxbtS5PNo7GPG3s0s/yEtN142n3I/liZArxzYR10N8I8qaCBA9
F1jd8hvtxAVll+oiKg0p160I6hhQ8g99yGArN7VeIGc863qbY4+fAJowqTdtuqD0
YGhGlVsW9hrQLL11iEnbMJHz0wSE+s2D2qXOxgYc/OiAkREpKQJtdZYqpYfSDttA
nzm4fuuYaPSJf39YVK/FeACXGtRyqZu8yQlDnqgwNOvxRnZb2BvJCGQGN6jSVGqW
4k+FwKOZI8cH0KEIImNhEtj7yyQT7xgQc4GdIxIf5VqHJLd0YoE9/W+47/E3vRfG
C9g38Zg0SSdv3JlmlAUGVxN30uP6it8QpXL7BjCBByU69078valq7HuUilmdsUHX
H6ipI8JGbFIgbwTbB4zq8VqV3t3I4T+6Yfxb9qAelGcyTD74oNCNVLFykHLXeAMB
ajmE2NZ//DIlGP2mYyG1XjQ25uJB9rERjuOXoc/1ONizU0EnGVeQKd7MdUsDHgCx
tqxmpQ4HPZiAxUaEFNQmkO3f564PClljs2MiPCoNmumsI+xAmjGW+13Y2hLnn1Qk
shrpv/QkBUck0o+HG+LGkugAuKKbbi4MCGRNfVYBHWIkqjujjdjj9bLhFXaXkCFF
a+rJQ1lGLr+4Bizs99vHF6QShCXVlJs1avhZtoZa4VBOs3JnaSejvYfZeNrM18ik
zZwlkkkwGsnTOH3yKql1uZ2Fp0DGusYfbJB92RjHWsj0n7NNRuVfbd7WQ8TSa+4l
cy1BqT9yZGSoMapQMLXrkPFsXZ/QGbaH9otyoWap1gk3O04Fg7SozC1NSi5fNtih
YMyAWoL2oN330jTvdWgwJ2Qh9mG8gMRFsZvhJCSxT+eSGAF8dPFRP6GDEMmUCr+3
YUr5uOMwRUPO7patTbAeBXu/GZ/mO3SzSSMCvVDS1g4wHMNi0Ub0GppuG5x8ZK6V
Ez194QCQpW9qiWiR7KJiJTJbcAc7kWoNwIMXD1/Ac85fBldOlthlI0DiMYl3JBbw
LIVfmUZh97aF8z0jqnrUvPIoBjLi4sZ797yjFgE3HQwI4cNpav8Q561ZRuzu3VvK
grfxk1Af5K+rViZa8hKICW+G910gkzOBYH59jGoAbCEzvWCX5inbEYQF1t+OXhYW
7jfvBsK9J2/M7a+/B4l0ZoswKygwuCO3L2GdnNnYT8ZvIu4gDNE5jE58BeJbsQ9T
4v+ma9pBDl24DijG+OsPQVOEObUi3qptmdkGZ+GygyziUHGwbrdaFA0rKy1tQnv6
nFu+cJa5PeDzvbkYIJ/H/78lK4ihSiv5zSoH8EVVaE3uYJ7buo52ggUoFSWZOgAc
d9E3pKvxvYUmM6UMhSgVdmTLef4hv7lQBMwmx+lr4aQlF7m/QVkXI5uBMGZE/Lpb
VKcQUH5UdCmoEBvIfShqxhAZK7foL1Jm12mRUOxGbWNvpiW6k4jZitCFBfNbyOAR
vzUn8hHb3SOyVDHmF+IzzRyKLUQRxqjNdpRr0+vQ1W/xFW4R8bc2t+jHdGv34cYo
aArNLKHE1Zn0nUMgKs4BAi7SaQzUvlcF0vraYJsIkFjvCfkVt93ZBp4Xl4o6VqTz
prUjeHc6XOSE1BPDH4NdQZi/aRNydHvUqSjVmgNOqxWMM+uDYABa7g6DCnjJnDpE
Rs70whmtNy0zEWxZNV4etm8kjuht8wodR+iisvdwp4UFdaP0WcYG13Tkb9KVEowM
J3YTTS7tDtj+GDAOxiHQhwsdsJ4UAiLFPc3J0oDKWZEx8wFxwMsBHrak4tdnWjhV
FXfl4afkxBXY/yWYwY4Da00SfbAN7AA2hTRCLDJ3y/4QxqyuoabWTvb5AWsu0FdZ
KCQDnrRXYQoBjWOearYzChe829Vz4sHEYbl5Cg6sTp7ojj+TCWt9jswB7934w8Ce
EPXeLEExl4QHTsJu6yz+19A4lVY5wDtyPSpbSJj+nDzQdPTMg2U0sYhkd0F7faAG
jt2Q8PAAiF8KkmV4FzTtqFVC6R/OnmdcG+JpUDC+PhLLvnAdXorC/o3lBa840wy+
+V9n/CECkok/m3Nu41yN12vt23+bWKXrtroTUYIoanQZwmoPIXICyGLEo18tDfec
ube9Zd4W+Pw8JAYsVj21ViJRQ3+l1ANwFCAhxTpwVEFAjmm5HXa4+x4eUih0faPx
gQe8NdxBBMGtBBNtop+mNLnSx+bPFi6iCEz6Nb8yrpeubr3AEQD9QBjWqn8PE0mm
uAZ3E1EsCj7kQrIRUduCzNZX7nFDgJqV6XF0dq1Ns7NrCgPfSvSHCNVsiE611Uwp
lplfs/YY9cOrlyUDxP0e1K4h+psaj+1iXoLEgpE652oqNNqxBwpB59hqJW0Me7Kg
dMeoEnic1uDhiqG88V1+KUmllpFP+HbDlz9Rvg+JEqASaOMs5tle+SetNxnMVV/h
z2Cj1m7kL0xzGLdyVzSLNGNMw166E+gmQ4V23GP6DKbVh7FFojJq2fy/BjDlS46U
syjVZpqMpZadKtP3nqDVyStxT9xUt5vWynYfwyroCafKTbPAtx3itv1oiXq/2fC/
OijIoCL18F1Y9uMKxJttsiBbzOawun1i7DETWDg2d3veskcnSEq6CgDKehPkS5SK
CiixFGClk1YxMmQaJFEwcPvvjpCndpp5RqPQ88/5d2Y/VhqYLmFdZvcUIMX6nGcM
C+8Q1ET7Mf2BbThMIZjmI0jwOdKviRozc4cdErbgkjTPsYy1WANx7j7P6RvPh9fg
oP4FVdEJbrQBviB3oPr9euJJ0ubm4j0ArW332ngMV9s1tJBRF9vrcbTbqzsX6EXD
sSs8GzGWj4TneWjzTVWTmw/u7V87g35v13m0Lz4fr+RzkKCrrQCMxEF3ia6WlItK
Cp9Uo1/H2xIY6BwGJR3646o7r2exylEErKRPts95dZf9+9fdLjxEA0j30cAQsUgq
xccjb09x/k95ciKgXBsWTc7oWmYnAa6fJmd/q4U2UObII1Asp2AawWF0aJUSQ5iN
v5ZD+F7bkBX1Z3LgdrcqemRrC13v+exdLFgj+SIprf/QmNCy7Z8+WyN9uKkAXErm
A+aguQ25Cko56U0eMCif7a2vOmTuu7QcP1TKI8SG4anHibtYLG4foEnvu6UBkKb/
GAVVviBHYhMHISg0UkBic3nIX7MjxhZQUlhOLc06y3eikUHSHpZJ23xFVwhcFVpz
kfRpOFsVhHhlceD6FSCnTMSi6G22wOZYxM9kbj17l8ed/lq4kSsPcWtxi7suaUGk
8HhHmfOasAHZPm/zhzc76ruveHfadxEqyCz4bLRw9sfraIs8jgSlLyV3cmQFiLD2
DAHK+Q45VxgBm2SF3fcRI/5tkaBFuGTzsOvffKGWaUzqrj4sPd3HI/0Zcexb2h0N
cKlM7Vr8K3wcD3PsIBs+0Uo9qcnMM7DOxSwuaKjN+1QAbMKeUFh4rPkt/rWcUgnh
niBsSLCQLOYHC1RPqHv14bOeaWzzxDUy7ZKGT5dEIPbn4N/Mz4UEFx6z1lUf9sID
cO/ksUF4MgBguZxxPJ6uTgGPbbCQU45xPPG+/+aWz6EQY2HY7gV0pk00PvFdngoN
Y5OPRx63cGwMoJ9KWvaBn9thyqvNJPRLaslDvalEFqXvO1NctDfiwNW3DcML72FI
aD3286CPC8gT6ufRGbOWmku5gQKBzjHknL1Tx/rs4skTTIEFa6MbLTxhqwLoHrBU
4drwtyePBFpYRtHL2xRt0EII/oCX4DYF4GorlI7kgIPBm88LS0Pi8jwO7NRMa8+Q
h8Xd0K9dTdDlEnUHM0cpAyNof+U/prWE9cPP0DezP1IoG9A1NAEr75GNkebgOTIM
8R1PiyAPYqIrD4w1Xf2/m+941MBgYxsHwnfOu6wvZyzNcecliEc6Mjh9yv7ig+m3
OcYiGZDsO2XsOKFdWwqZLKbfobFUzp+xGp0WBR4AuuMbUDb6yVdS6xS6rd5ZUVZ4
fCr8P1D3yfTOl2Bc7hhstQ0O4rUm1G22UKuRhNa5f7avK6dtVY+8cBN2EIHpOoWY
o+WSwHrf80e1RUS8+/aW0rPCoSY2ZppRDqodzaiY8N7S+qEjThe5ANoc25arDtbu
deAZn03Z0Loy0DqP6h/2mSbkKcIXa9pYGo1uvHSIO9kgbU5UZbTP67GcxEWjOtTn
l3hQYzI9Nx7i2W3DCpLGK9YCN0J6rQhp8al6B71GlRH9UnLdYLiR8wy4W3MHGrMv
3Vsq3/Zb6lo9mImvXMmdklFn2ILG4LZ3txh6XIEWwn/uMveUUhk6y15mYY9bCGxs
QHU9o0kWjDuAfO4RhlApP7KvSc1AVBihx83yRfwQhDxcWGuA4E9PHqqIhglhPSUW
hvWdwfZrCsiL/UDWIkPRJ/VAnFJTjLAJlReBQDRuF5oEBWRS1jI7elg/eq2p9izH
oONgZh12e0dSxoh/k8CI6H6SMNoYlvW/1q6uv1pKGT6h+16MmkomyuFww/JxtlME
SmZgyVKs+fMeDXqeSX6fTmZWEcfIj5OEi+n6gIOn7IlxkVwXeoEpLlkzAovF7b/7
IztZELjDda2FGidFQhdSRAbdqOJw3KDrOLkLk+Ur34LUFWhiJlNWtMp7C365ELyP
CllpRuXK/ss2kpze+3VLuIwEI+ON3tXnqockkrBthTcRLV1TiJIhYHHEZDkKwKJm
LbNlSHPSKZuwB+u8jWRmeXpbUu37JJjdYjDdOyDnuVKi6SVzpUwmvdRgeRmHkhMw
s6dGKlu2I5ebIX2RNx8BZLBJI0l8CcvUzixQgRDxFRmT+aTCYO0b6vt1QH1i6kFY
a4tMkMttEbxgdrVobJkIsGv44QnPUmxZmwBZeZgk05WqCDJTqalcY0TIatBHLDkg
hd8vSl1sUe7z5JgO9A5fTh5DBCP0LqfQS4BEJdqQX2fPf7TuCwwnMKG5D3ZP9V8g
Di1I3AOj8Tor5Ua5WuyuzawVs5uQL8Dvh60LYM8NXoFxeDa3TYfXKVzlJPsJNgbs
qpUeo0IYGvqTzEl8VAye9NzmYzOA3pv0EKhk1eQWF6eu6B6NrwbL/2qBD/ZuAqW9
KwC364Vimf01uJsv4ApBwUbXjzMyWwGDNcKpUIBJ+KH521aupNVN9RWftFx02o/u
72rreA8RvZ3aMwG7QtRKHSK5Syj5Z9sUdmjRv7Hc3BSINAPcwTYwa1Eo9Lizc+xf
6jGJmVvfgdSmurVlPQwKlO4LbSjgdfF4ZQYLatdq/EZ+Mh1T3rgV2kYva1+nx/vz
d49b28epSWFVdoMRDS7c5elG3WGPxrFP1F18Sy3d0VF/Gbl9Qx9fNPsualSjCVT8
NmzVyhVDPaOV2GwAYtoHIPMF+3kbw9Ki/Uj8WKPie5T6FObjqzYZJRIEBNoG8tVv
NrDmThx/SheKQKPt4KjVW16bG3e8QPaqllhFqfAzw+Ni+YowXB7qIccNNUeOq/67
Lb6OBz+VldOT071VsfePZ3mxcjXZFEAnk+uYn2VvreYm3cc0Zdn2BsdrhKnF8lN6
VNoqpRm/cSupQWDO6+xiXXoj4YmfEAuf5cYYKstMmInOghNTaeBTzeLewiB7Px76
83Ju+JT4Hlb1ZjZTg9yYSfKSUdRjQSnx4UurlQyL6mFbE8+Kp7ekcEwRw2lMJsOW
2o2WTc8RwR3XUMM7h3ifJQZWxzo1R4xFVnfgChpgZxeZBP3xn/gGTEtIneR4zgvj
XfZQo77XwfVQgpbGTNGZ0Kji8GK904DIC1HWYyu1b1CR2f9YaXTzWdBzpAqDxZY/
25yUaaYx7JNKtociYtV5nvLM3ydNGEqCrGEC24kIDZXrl5c4OtnIOWpwHEOEgUX9
/J96QuDCpm7jfqtMZm6HrjddsWTt7Mw5tOMAuxJNb+J3XfVTGOU2CC1SC72oob0h
F58+NXZ/NGPr3a5N012kX6x2r5niVM5HdGBi3qHIuw6m089CmqG6UTfVH18kz8C7
9wm1y9Gf4hDWBXDPcBR3N0crYd82fejL0T0hSW6aqM+qtjt0722EA+n7urlZOegD
CoBCftRDC4heZh/nlbLMkZtkrW9ILbMZX/F8KOf1oAHHTv6XbNDomAKzCBe2c2PM
rtxs/fjKHF+5SR5EQ+7XXNMYhdSxhm02Gg5A+Bx4Cu2z8XQU/yuihUTvBIjsveZq
/F3iQZXFdp5o+IYf6+5ips1BAkeJd+8gkTalDL6ZzgxBnEYhKsYryyfCCGdVga+2
PxL03MIYRCPYabQOyaOIANP+ux9AK4LOH+GkEmOk8yDHLh1u3PzWRW31rPc0VF8g
CsQ/GwTqPVMQ8c93SumSjmNRSg7bsxMW9Y44wX8ejPPeir7AEJKk/mkm9BslvIpH
ddlLTAv9bWcl0+lva5HdRXEZcxpf51M/2a10Vj4hEv9Z88hEAj6T6h1FGd9NvwUC
PnS8nd0Px/jeHb+YjF9lC9y610avTNNH1i23FFMUYAoKfn4iChz3jSfqycPlC8BT
J3LnksKlYIeNFP6M7VZS5CveyRvjPxMV1FAVMkpI2r2lKiEDwnUglwpjzT0mDafm
F1a4fnxfxqHEq7bKcBIloKRwWpLXx3O33C3mVWaNgqVDGAhURRD2hfoAat4MLXU2
FhDdLduNh4qnkOgTtfyZo1VxcjWkFxhGvtQ9Qhs0GBIJ8+EXr9LxPm9tHg1W8Yba
T9w+1+B6MiiYVhae1bMCxEd+B3Y51DsVUgPcoj5g8n33pnFPIopFPSWhbadMJE5f
QxOsxdE28vsPKThWkIbDol5Fvfq9BrSLokUpMnwNnfNgeKlbeDF7pCyKDzaX7DGn
SETgaezovcuF7uIQ0uKZbnE2Txah1VS6u/qr1O7uQDZvx25JgmNmoK/5dmA7UkWa
ZWtHguSaHchn7KD1mLz/MZioPaAVxZVyK2NnBcIadPr7QaJ9vF+vJ5Q8NbYcabwb
oY86qBrjIskgpGEk+SiT+eh9L+D/2hXJPqSUKzHeEoP2oisRxJKjZdKVK3Uwimvg
KHUalnsX6PuI8WeMotVVlz2H06nPBNkQ0o4ybgblTkdLHYYuIphWBMAU7qfthraK
gsSUMUPIaQc4X0p41zS8BYIH6VYn+K31xAxKuhNL5F93Ds4d6TvYZ+cePYDUr6+6
UPcFlZTQhRkIQnbJZ99/DxdgQqvj0MSr6wIZmarg08Y8yBgAsfP8oqDlAurFTVgJ
gO3H127MazbJAVxd0WZDi2A6TS53mhSzTctDfFUrIlSGiOWDEp1FO6wJ9h6fE4/x
97EZR14M7SpRxFBeiWw4vJZhQllelsH8B3OtwaDoWNNZpgHnhuG3sHpTlvRwJhrn
5izGyzODLBVd/rcfExjbEbBOY7dGI7QnRPqlYOliTlDK7QCG1dHqpwV1p7LRUKEm
VbNc5iyUzFRJzgBuZ7Rm65q78+Pj1Pi3glYEDIVl8UCQ4xAkYPfer18GlC3+Zuxr
8yhKkQ/awedZcQJV3dwtr/W9fqUGmIIucJoyU+nnY2IXiSU4SSmB/iHeq3rJcsp8
2uL64dclvHDaj3XJMp1Rkpl/YH0UxwiGNIvKjEg9rfibgyEWdXSYgNbv0sSX/HHY
986HNfteDcUJtWqIfrESCJ/TEVgBAkLSrP9ljibpU7ylK8bvVVVmphaNbSwDw4uV
BhTwC/3LNmC/Ftf+RfShW29mtWkvmxb/tSlg/G01unH63Gz2me+2NjcEJYFb5ggr
ZxAgm9lJJNQ9eAN0ocDLd6XpJzjjTPXtNmxS5V8k8urR7g80gmwmmCcTDyTUexLs
kCN2G7ALHoEmrIRga6KWHzTO3ETC9hQ+VigQlenDMMg54jpkmQ1xj7N1nexehuRU
gdv+hbmA9yBzg9o9gVk1wrt7FyBQyhhAI5fezT9JZuGMNwpBdM3MxFRQcW3XnU22
sby8VP2DZ2bADyvaPTfLmiYXiqujQo3LYM/gE0QUlHVXGGodBpG4NdD7V0Yjsk9t
1bG9eH1vYPdlBAuYwB9E9mlx8Nt6lFPU3cGxxHPAl0l8kIwzStubPPuQMzZX+Y5Z
0pIOxGR6lpAxIhWBL4jyYmS9cDrq6fKMJlMVDHOIagcFQMQ7z1FjEnJ1hpy1e35/
+jSOpauIOOB2ArpGNiQ7eWDQfd1JsD0tOuDbN1rxngqdpqtLDVbrxnOjD74lknNX
57037JhNEEeuJthyBXX6XYLixLNgr+XGJ1J7R0zDVA/wBS7Th1nEHpr4d2xwhp1H
oUFS7kg8MPhmTDmAPketH6LDsqctWDCFpai0+JOWMHWbX3rxnJliwfNtJGDEO34V
mqaVRSA9GP7Z8WiQNhsuRkEv8wgVPuXH6KPjK+yUxUkI9bp1CMG4U6aoBdmtVPCu
4/tZK9cIwSFT3ha1wAXSkGfnGfbqVEQPFYbWnECdGWn3ucNBwxpaTEmdJVmtxuQX
gSWXEdBvLpbZRG3Sg/5ws1f9U79GF8MqV37f8aFP+klYzwVB0g5NXYYKepuo2eH7
DiLX2JcUhFcSO5PKuRNDiQ7nEsveKXWflgobDvg3nz7UpsemK//lZgLLctkhG5JT
xTQpG++cfCsoTnMborscp7xLrf/q7EXiiMbkl9blMiKa6+LJ1lIgrFqlpTYzu4yM
QzXhdLPpa8gC/kjR+CJcvgLX03VdmwtlMN6X3Nfa1mkXO5DRKVgMPT/MMo3VRLKM
0RANKQUkq7rikaS1exf1kHuXLsw71QDua9XZYhERsP5usSUTgifOWk1UpdIea9JZ
zdn1UPKXp/vz/WdXCFr6Hnv3mTcyVtuIjTB3BK7Mluye+4vnKBsOHyXgWVlKVelx
2bzyZSD0NI+m5Wb2puOvTnpM1l73uf64bf5axbyvLfu1ljFdF/bar5CloIvvPqce
K/rJmfE0CF9eGDR1mSTBxnJTSG734vGViA911y9p/DBNl8xskkoDQFzEtkQ1TLTO
0uhA2XsLucbohCNHE1OhN3QWu7h6vfVeeaf8Fz5mzSuvUI/YxLiBj4BIKEM/li5d
fFAS+6PCbJcTksMkTzIZ3LCANmfhXde/TGP36cpxVNF74FtS40YyjUeGVhrWz6j6
7uzn4ca4waV8dE0U7FgzwYA5eZBclqNCSN3kQr5ejQFVDJn6hJ2rpoXJ05s93adX
qzQPfZ7uPxuj+TapcJXbBNyoPl9vgwKXx5N0dlAksby+VL2lrS9fk336YBbzxTfX
/DmPpzru3ZVgeVtVLhHUBDcDJtiEQUSUx0HRzoIRrOAw9TfujpgQns1kBJK2HH/v
in3nnM9blkQhsmG/WdNW0Rh/FQFARTN9KyYwY28K+ztux2QQbnHL+cZF8ndlsPQh
SBanzP58ZCFeF2J7JpclRTLNT78aclxy4J33zO60FKnX9ZCLnTI3O6Dcr1uiXcRO
SN3oWhRoBiH4aTi7i7Sz4Yj8QHUJ+rVyUK+Uddkq4GNnHt6yXgojmrMsyeDVu5MO
1TkZrAHNspMKsQO1DllZf9YfrO6IMFzziian4/XdpzO3bHFeeUHf2UhhtAdHbQY/
ixuLawU9G7LTaMC9jBJsL/ASZS8JD0l6j6GN6BBJyPSNeqD7IHcUHgB4Kb6Lws88
xijYioSMcD/ALJHOQBVGTqsBuVtXxWwYTemtJ0s8aXfsFoT9gEYnmjCyKF2SpJ6s
GcFJA+kLAs5VaoZ9XPUOiHMFeRqisin+OrsVGO2qj+kM6REDMDo4ZYcOChuQyU1x
MPIBRSEltem3F5Yn5VtTcid3vF142yvvCvUKxCTkQlU2fKYB/YfiMbj2l9aULvob
7X4vc09OyrtBtN+Q/VjvbNTDBiKf2k41Ab2QOvLqZRGjbGhXf5PPuOhj3j6o1W9F
hBCFtmkspicgh1n/Lb4HB3yRRxRu9c9RZ8rygU086xMCbnwiG+I7KMppy0UOztg4
3LN4kA0AZZL1L+WtdEigP1LFXe2Pw6a4qLq+cD/CMJHQDSzOnuyG0YcMH7brGpTy
LhkZgxRGYnnkdIMEtOgdRmHpxGSDheFF+qKf2gQV0CTdD2KfKqM7y0FLP9/TMntv
/nb8YqhYWUp7FdG3qRojDMsfHH5tc0kzAoE6HjnjMbqVB6VmCwMh2EeNkqxRfmyY
vVvG5ybBTYHgMi+bEId4trrY2Vxzbv3ZRo6YZtRZnEuVkWVUq0aIRh5uTfjkkGu0
kr90LrSUVLYAeyei3pE+0R3CEv65zW3GHj4OrnJiYHnY1dwCsznunQEdq1zw2ZWn
DXbVdY9AUQ7PSKVaW8PDW2hK1iYKzKhk3UONm00NzrMjHp+r5bmCha0/H5+N8RFQ
LyOmxkK5C0PM0E7blPaKFnbgfkY3vkILdTMwWQ8J5BoiuEO2CkmuWn04eJgnhAZI
my9BOjtyQQrIWuM5/bg9V6mjyag7voCeHOEW75ihnSIuK3qSLqmi8GsSlCu+uATW
A60U8OuWrOfQzeRbb67b9Q+Qy34v77lLvbRcycuf5X78CjgtDp9qR9OM0FMjHuyi
mxwKvYX8+MogLm/Cywzg3pbdl33D/FxGLuTByb1reCpc5O9CSF4N6eXwDh/mdK2f
YUhfQc/vahAGa6fypPqKg+i4BMeUvjk5AIFt+p8IRtkE0xhdJO6ApZXcrM9dmSJl
uv9NV909w9o9osEvU31M3vfaKqo1b8mV66KyRgXT8fM7fMIOxzqhxX/P311C4dVf
3h0MS/lTWUQj0szigzyVZ6K/XiiK4MW2i5ICgPtANtNo4BBcNzyRcAs9hsgh+yS7
b7+LODMs2iIrGc9JqKHfg79MvJb/fnaapBiqy4oxB91S7oQPAru/GNkwpaqvy7ub
tY9x0ucLFd2oOB6mmFgzppf7SGyE9vv0cazkXEi+ggda6sd+9T+u5isizxy/zUqt
ACGV6PNAkcteVZS8lWP2Ozo3ywismDet6KAaLBywKE0++md3qAahOXq9k5RrMSME
DOfD06zWzyBb5Jit/8CeV39L96MM98+BPbsyOon+zNjZD9YBLEN8MWuGh6Tli6FQ
qNqjVe254KRb2wniKABmEE9whck6CaQGTiy3Cu4pPvkR5XfakVKTQ72eOcGm8RgL
gnxWHCWZMfbokQlHrWXjGjXeOurMPukVZQYX/WO/q/m1HRryklCWOqzNzB+bSP3s
kjFLZAqcMQd0+kgtaMeDXwZTOb+8wstxcHyfJ4soq1tP0O/xZtwjerUsVwzAeH38
0hgIiaWdEJB/wuKhn34xMoq37xphJDIvXhF21OMeTDihpiZhxau3Je73CGta8on1
Wkq2dENaKZ0rKIQUNdtj7GwYyfUU7B3zRl+9QY71bJ8DCmUktvpFKS59AlMiVa/H
4IVykRm0Aqm4JuVMO2DWoOedemu29YiQ0lNMCgbvb5ZQ3RH1yc2lLY8qCcMjDxu4
sRgSSyRWI7I0+gHQNENEU6izAPajYcOHpD5HEHOH8oaWB2132+z8vB4kpXqhGacR
WbJ0pDEhCoRZmO9eyAz1IWSj2OT3sTCAfOSd+tPU8tz2JLopLTQi121mxqsMHmFy
VxZs4p+x3+zaRRrg2EJmPjogkojRxYVAzF5Yf7UKUfJMaRNvGGYlYlJakP2H99Tg
Vh5vJFTVqV6UhHFbf1XnFdYLO514OnDlSuAyaKi5ltGMQLdC5pZphv9NkWhdxBdk
jy64GXLzSfFcIQMfgdJMrtacKKjgxKIQN3jHf2IBOuhqtyX/RUUtB9zlgIA8MNh7
VW+CwqBQkhCbmRqqyqcuDkDteS+GenWQ8biBIHDXfizso0FGjMpbBo0HEnowQQji
84It3vT4GSxWQzb6egCmZle05lPPIEWennEeEEckalSIZyNf1joq2SbvT+MLlKYw
113IUmqhQu9mtdtPVjsAi3W8dq3x0W/f9KwJXpx41OGmgdftDJbG0izJm6FfucZX
0BetgsX86IBuhK6PlzUei2B050m9onw2SIfS4JOETqlQfRBVXBybpZWc9zCd9cbs
H4Ydtx+2UiNBc8mBmY/j/LX5eanQTTm200qgc5fAJFP2TFebd7abS2PuPzTb5dKr
2TuctiTy3SVWu6lAxg5/ifXvGv79eY/cun8TBGuUuN8Vnel1l5wevukGsDdYEhu4
Kb0F02To466dMwxejGwbTfm+rkEd6Ki92sGBN7Vbyww1M16wBQbr7A8PLos3CIqz
jcd5LE3Uk3XD7ugLmpYz/OhK0xZag3+gem5Wsq1VO4PKA0tArqvAscn9elDVtUzG
1fxhBRIeL2MPsKQvAYMvUCVsD3hRT9gdmSpjSMbyJnFPspUjRB67Pwo3ZwvwIptD
M2r2lwLzxMFD3VEhQLTDoxnaJxcZtCUtJWUMreL/HRADZkJ5ioV0vr2OctWz5tFg
V+ngrIRDPBkFEGEnZkRwWZKOFHd3+kHU06GczAWB+dVtwKO43F5nHb5zLP+JxEyi
br7R4aeG5otJYU7nn2WhADKZpprOytbQ6BaZndT5cSncsXj+TlbXw/IcJZnB7nuu
v5X/IQE8zeX/Aqslh7+ZmMpOG9vfjYx1SLGLdBJ9p8tICIt10VhwnhhHXsTomEpJ
30ax+pnmdO+pPSqabichNC7bmB8/UEEvpQ2waXnF99f//AktKxk0KmXjdaLJLC6N
ChM8fVyytzw4/bROH1PIzHZLutoNq6SNrl00RRzszNXk+f6tux1X6UsnTqRQmugs
1QILC1qQfQOzio+7xnw676vWljnlr/6yu4Mjq0muD4g2GrvJaWBrQp6DpifyLZBf
kJLqnrFGZxXXBbku/EzPb5SlkbIR9zMJF4kdF5skIJaBIw7OgP2EB1r+x/pJeQV6
thbjINx6HHWPWn5zzJICnjhiKX6TQVLm0kN0kXWqH462eS0IkjbuubaT/SWQ8mKP
Kiws5V6/MbHGfF82nh13mphnzdaBnJvdqQmXVfP2uBmvUmDLtVjKJA2E8En38YAy
fqu8OQ7oBeCf8pCOryAybQ4sdaSKlXk1b0yZDGWX/5ppXPtiLkBdonR4eobQKO14
S+CYtWIL4756xJm/Bwqe4dsRQ7svH8zOvxG5mcjxp4Ai88tvUOV5yu2BmPbnMvoq
ae2n0Vgaq0QolvEpD3jiwLFfcEP9LM0f6DcaZQH2S+NyzAd7k9wLJgrgXD6lZ5gY
LQdbG47tfKfe3ISg6lsjewKkBfMb1ruEolZlJGsKRxtpTPL48pNLOYsC/lleRyWA
QIitewtnZhLXudu18TZoDZJHGiJWlBOzUtsNJ/ri1NfwRwRETB3Ba6HmhfJpxGKO
B748tKnHA3EHTmWd7TCI5yLmj9z6wUwo/aqYRsIql1CXQwueIwZ7xzEdFh5rRgg3
9pw3rf8/EqcW/6IhKmpNMSPF5aemwVkfP1sF4zdgLcfx8DbLQ0u+RmH+RH+HToN4
prMBA+pYKhTZiB7CVOjOJJ/zvr5vzvziZRHSZzoL7rj31DKd/iJES6TZM0eMBWGV
fEA+O4EhOujvlgPbmLSpauxuIEEJhfYysXy/AwiigT80n9lqOrMGH0VyuHTlSzbS
KIFgvLzKgiJSTQN8hanhqXGkIlQtc1pGv11mGA5RMz5OuOA0VVegrsNFqnplf7Iv
jVXHKnUccFuAdn6fke6h+XexSApT3jebLYgHh7YyBV6Ckz2icyW+r5CBkWI4Mler
2o6zlLcNLt4n/QZAmqP2mMUbO0IuWTCvrwy4PkuV/VF4655gSEj2pEKaMALBz4oR
I/3ayItyRJHGrAdaBx+ZYXcQBAuoAKpGCGAz0G1j0D3v3cf709Hu+i8tRw/zbdFq
O+WQ5il9fr35WAql7xyWtZsAE1gHs1ewdXkpm1zNHCfAlmtm3UFbg0+ALXAGd15x
cmWjajkZOLxn2Jmgc5KUjZRoNoWKV3m17Agj9UtEPDwavwMnuEJ6H/P9YW3DKPUr
/agS/clP2gbgOqv3ImwMsj+56E8MXHDLfJyRVinWgxLctTYeJVyA4p88IB9IOduR
Je9wXtVXrfLVfySl3r0fLNVvfHVj/msbEAhozY5GrGGrWHk8TTMISS4XbNCUr5Jl
yOudjIhKJx7xwLNDi/Cqaz9ihCE1WvFtdXe2BGTpGw2s/gQQZajXDjam1zNKjWW8
wfdnBZ6SL8jWeufrywtD+3P5YEjKM0ALPrpf0jXdwNhngpvH84eiE47eFnbkCN49
JfAwgPXrfgfcQn+Xq3rNBa2sezNBhhmooY5DfU0jfHrnZkr6LvT/h/DMW9uQ+EJV
OwcMY/UhabaJPx4KmxuGpXP8KezRVGJuHPKZ9ZpNGEk/eWmL+FJf0UOsXdaW/xi4
r18SGBQV4k/9iyOAhLoQUD817D27Gcf6Xbs/Oy/vaN9Fg28Aq/3ejIOuUY378F20
KnrMpN8lJaAAmPwdF5bHFUxIaXSUZ5EAhn+aFp9PZQoZruPkXzaOL05e5bxxDmVa
0ti4AgTg7XXwFlcIxvJu0Dk99MJytq+WMsl+teNIP28k53U2CUUxspxpGHld/cku
s2hO+bgiljNtjbNlQNWuryQhg8PkeQqhXa9DL4gCvbBpbEp4QSujpXDkdh3YcE6Z
PbEPcd4Lz++MpT/1XLHxn7NHRtHFvivZQhNH0j+JR5UQnXSwcyrE2M6AlhORcxD5
nLnzea3VHiJV4+2NwGdA1Q8wSRKEuLCXEkMljWvTvmvl0EVT1oqmOc8+ibsI9lCR
sbdepYiSWDAtysjRfNPRLe5YMECkL6eTYzoC2NN5DItZb1rECtmbicf/BlklLkFq
xyntI7X/xB0MybGpi14Wl8vtQ8hjIhb6/o7l4llc7c/aMomp6CF0pTGTT7RRRvo9
D6K8dexZForJBfLUQWT0n5uOJKcA9Vcr3ohpVptWnnl8Hf0a19QDfILH68enVrU/
rtqj+atV3dh1Py6qnZZ96n5zub2i05W+janLingWhMx89SdtwCATLXm1AShiQs1u
6tl1nDW2fYWVIHlUsZ8TAJ1QfTD8Z5axeXzwfUOVfV1wz2h7geDjGaLaY1vj4cMr
YHW4TlAdE9v2HwKsriy+/sj3Xt6SzvOwH0nQoccdBGAlzzVVojdNDDrUPoDcyEL6
mrvceEz3MoLrEDn4NVvsEbmuM4qtbl8uPbtFcfEsxIKk0Sgw9q3kSDTn/VcyN18i
4+BGlzPP1f/uZXkQb1T/+ee8enp8TqO8CW4u7MqIMpAGqxw99YfDBpV5HtyJw37z
ttBVVu2aRupKRASCepZc/42OG0v5cW4ERPXVxBi3hKgbgPM2yUPJZm5s9ErXC2JH
CBUhcJMadP4/KPDrp1ARCrlsmsbUNzm9Zu/ajLnqiaJZs44uGYKlPiGjO9Nf4/FF
9qaxggW4kRTS4bqKW6kPEKvOuvSXz4RiEDiRYKTzBZJj65V0QRGl3pxZIWeW2G/g
0owO32HQPchoTAi5+mEEyAYKI/h7DAkVOhl3y/GbbgnrdtHlq0fP9S2FJPbb418s
6xoNofn385b12f2DlhdjTi43f37C8CvOd5Tdqlghha19zF4ZiGXX/OzdJaJa5B4Q
yRIyaVEAfNQJsM+OloEMLVl5aZFZDW41kC5ez1LMRoOYzb8MuKkb2UGd4u7RMCbU
vbSGNd5ji5PDyVzWm1nIsdro4Wtl9LZbDgegakVMiOWfSWMsgVWvpNlE3sdICJaH
bBqsEXh7hCpRij5BeClWlwZGaahA4S307GZVRTEsn28kAnMaseqiLm2y/bm9RCpL
3FNcRx0wjSXGD/8xXSO+QQaKy21G6zI/3eEigDdORiXg3JhN6pQvYPC8ESPE1bMR
l9irtug2tbfhfawNik0lQF/DojeeOkBS03rUwXsce67tvSwT6I/BPioEqj/ciCp3
9mhUAyudaNiyJw4Q83rP4qOCddtDaTiPDB0IHte0uZBqdnETGt3EiHIO6Wp9rnsQ
sahBTcG8svKee5aaGAxkXFfiI7X/bshvXLIuZSN6CWrNh7ADi/KnHLgIDjoivl5V
TZWXF9aVf+6+WL+lEDTTlFYON7s3cTmNnoBGS0Z/C5lRFQf4C1maSbhstduFmEDm
VSt44JhhUsmJO1UltGQrybXNgANap81kOdEIKvMiXKyY7IU65DEp5UfVlQ/C0qLJ
wu/BkNfK9jpf5IerS31k3jnVkh1kMVRd1dUgRcravvA1EVoB1DOdaDSVE8AdJfqG
uHioRckyl5MxGF6E3e2I/ZPvzgwQF6ssZIZpW7FDmVLUxC3aRZi+I/lNeBeG1VOQ
EHiotZf6WaswUQYaH5H8l8a+4u8FN9aPv90J4sOKUZ20vasYyLQi8zdy90BYHrz1
VMCumWK/BO+oOGngZMD8b2LUy/u6ya2/l4UxR24y7JbV/SOuOTAv0GkwIFGHIQFZ
ZfATKLrjkrdaPGrJM23u7DWA8fd1LNriQ2qCYz2Pqk09UBDa/fTgTF73gilbnZ0j
nT28xnkvQQ7WdAGpH+EGdt6Zhw6pfD2+duxFVKLy6RN/gENttZ7T7NC1U0+wkIyA
mMAVpq19t/dOuIjP8YIhb6BXicQcDKpW3+JF48sqZY0ez1a51tLixSFUPsY2zoHX
toHF8JulSOwTreLmavyXC1IRJCodIwtJAgrvbk6OuuYCIv1XRqI2uBhCanRpYQ0G
0IbqJFM28WQIG03db2mzX/8/UKfekCJwT2jzq2hFnr6rrRVpyZ5DCQ8HqlXQU+gG
HOLwpR5vxbxYZzIZjVdQEF1IUrgftUoFjMUvcEOBsvF9O1cPL19BBc5uk0IH9NPC
hwESW2bhPa+KWXdD3jv9yr91ja5MX85OizHRjtIQYRstSNZ8w9MTgnCUzwOnBmCO
BkfUdT+ff7ufvzOIsv+S45b6YZSXx6v7JK7yew3vNthedzYrfr1qsL0j/u7eSHJ2
evKRxzgqk5l9doHKRuMCmj+He0NfHp/QU1ndjCS0jx93qhMbneehQQbjluzm5jyL
b1cs5OHnedAQ9sOhlLg17Lqs6i7952wzQLfV0SWZunGMPHZq4Ribo16anSPA7rQr
9qq0kcl2koUe2bskbPPQSUjnK/fuXNbmi5pi76RTy86iVxEEUWMssBB0hunnpGmA
veFc4UT1CX7GKq+1S3MAQrBqCYjarBSmFeUUssd6QnxrM1QbuvYR4XhE+Q3mYQXK
+JJ5Uqbni3HSivYObFuE4u+GzsoekoMlDKnCnhMIFRSDSzE5a56xQuRfrvmjXWsA
ccB+xwfMBmlwH65Hqt/RD/MDG6tfbinIy+sk9iFVJLVU80KOjOb++XqUtU7fBiO8
HAQAyQB0TFwqQI100VtlhpSlaU/PMD4CLB4Yg29K7/kLhflmY2c9e7txcbE2vAw1
znscSfs/zQPNOayf18xmBfhxyKJ6ci+oTT7RHJiFu1hgS4PG5tiCrpPW7Snzyrxx
+g1ppuQ+Qxq0QUPlDatafscroRerFQBMy6HYubWee/4tvvxRPdnnf22RUBigbc4V
3vOe59l234JFUUIKQh8piPL59VUm+k2R6n+DdUa8SVicMoF5Vsk2W42jzB8fjHQp
5C0/FruZVtVmdy2/pJZlRR+WwQbOBlZkXcB4DWVaiL+JC+a4LEBxp2DC3IYYIGRo
/hoDtHGYKPmlpT/uMrIOTB2zYQGw5cZNGJ8Rryskoy0YWnZI2CiNKtkKS0YsmE2p
xzAV01bn5+2VpFkhrDU4sEPejptRegijCoRvlcNKb7BvRS730SCSACiYeEeLfAJV
/qwLwm9txKqBF/IAr/Lcd8AckplETwriQbZ6mL9rFjf+Pcj2s+11eYRaLcDHeFIm
0vu3NuBd6wINBXFQB2AT+p//ysctRn+EBgAgeTN8DNua628KQNGM+A3G9r61n5Wc
SMmwLF3Z4znaeM6EvPUgUH92d/8iV+g6wgM3KN+6tQCmKkfYqCbn020rg/LdeAuJ
Npp7rQqQjo2wIR5ZLi3KeZ7Ry+LiU2ESKsjKF5nqtedrjE8o1a2eX7qabhBS1E2s
M3PIj1nhcsbHJNSOgNddMHkkfEvPzSTmuzqajV06Dv7p1qCT/40KRiDAq985ZlRo
EhAY2nYksuu+d5HhS559QPjpRkMS2Tom5oluh+CIsgtWL/PcB+YYY4cmQPBllbcP
eBA6voB68SCuyYVebjtE+Bc9/h41Jdpflit3cdmdvmmzZIKwd8iM5yxg+0P2zRE5
QG1Q6ukXZxqeJpIpZCNpEgzFj9YmgmZPWmFZPRKy5+T/lBktog0B0XqcXnTk7Mqm
EsXmpMtwXIfJOfY297ymvCUwTg/MoYVM31GKjw83ahitfXsWMehAJl1QbRHL4JB4
OcmHXr9MBT6HFRlbvXyItqcS44vg75FxDKsjDrGhDkMKt3MRjca2OuiPQ8E10V2Y
vxfDbGY2p7LycGtSdbioSOESu9cZS6kcW8D7uax7b1h75UWPh4AvhVq+4Y5D6vf0
zngFzi9YYfKf/7k/9NQ9ipI65IQup4mErsC66CN0YWSbbwOZORoE0S+s9QZzAiAN
e7f36G+N69SDaVF9a+CCLYWvDLpS5Esv/hrQ5DL2tCZyOzfk9NGg3XiaizT7H8M6
X1YVJp0qUlfeiRsSqenlJEvYDuzrvWWvrj17ZGJdpZVSBFtGNykZAr4KL9zL5bwZ
HG6q1qhzm5ahSif/3B8JeTZpy+AKB7i1QUhtNK/KOvg7bFTNs5cOgB2C8WNvyHiQ
6BeUOmtRnUxZtmszNejJcX5Ev/RkaRofwPbb1N/0s/CXHuWuTgzoQCbn93LSlc5G
XCP35smfJ1LWhh5IV9SA7L22vidJdGcZnShgJ+kdGQqWiPl5ZYLwacoNMbtWNJvg
k8i23trwXeQCicIc70V88UU1MDdi52qNC0wRulQO4+WPg+vl5+Spo93y5y6xsW7M
BuJ1tmN8NZq14ziYjD8Znm8oI2CfLRdKujjEoTzEjXMd2E4g2UfMXsJC9dEarAD6
bCUnUBCfEdEzubjEtgZUio0UA/obAwiWCrRaIvLEZfGGQ8Yqrvj8Fvoo970BK0uA
adf9/K5Z6WIbG+jS/CCZHjA+xm3FEO8NQ5GF19IYnBlydExYYIAXnKWSHLC9p71k
4vNaFAh/rCABuVX1Ru/uc7aUjjc7C9RxAjTf+HLXPnLn0PvFjr3FBmHsBP/Uor+m
ByhehAGy+8NmYteTTnxU4YZIOVVR4v76GMn5+iW3yeL/f3r+89n8zIyt3umW0AT9
OVKPAZKW4pmxQxbFxZQiw/S4SqwDstL2+VZAPlxY8MvinERt9xQsErowD03IjYiM
Hh4wnnnzuKBERQx3JtEBJnOpCsYZodzJmr76daYdgHxnd9pol0s+wCWSZrXL+eOj
oK1zibfiAjPNYYt8HziqPQPGZLiF8kBmcb5+iBzXQXFRXDtoWLo6zW38f4/vp1uO
hd/mOrNh+T8/9onWrmS3TPsfHPPdp9lvd0ve6oBYMxe2GopJT2cdgBv4EiiHMfrm
+3S+9u1PTyD2+r6NEVGJNL70NvxQcgKIFrFY8loG8w358mvna1lA+GqVuHOQ7xvi
s+HIlkX+/AOaRRGvTOLR6/rGGA2uuoE2GOq9xfu+H4DM76OlKJDKysjFNBMuHECI
xEEmokXSKNg6Qj7Mp3fvOXiUzI666yJJxFYoMZlUyUllG9wApl2HlpvenTqDzfht
v/pUQsJ9wO6W5OZnnz9GxHG+h2wLf8kJPbMZoagMEEjZ2bO/zRcll+ZbYEKUo/Qh
YmGTN+FuitwSvHE1JeOPfuL9W0kQf+ymFAEghMWpGXrZ8o4kkQXleDzkKdjmw/rF
ojM0STAoba5alFDc9iawXwEgZjJyjYCH23uFPTESTnS3w8gVqefhvsdq2VQHoZtP
fBXv4cGi9UJcR7Y6E0cNm5C2Cj6xFUQQSOkQlWk4at8u+7mCimMXCJrLBwXd/SV6
vPcZw5vMJtH6QRJC9bf8tIMfUbkE/xozErYiflVaeqISRCpWx4L1hizd3ZpbPb6E
NHs2UZg6HsKxL9ROQcwEuLs7KH4zsGsEYeD6s1WdoreizoTyRsewTKYmlmaDxu6o
Cea7L25X+FpGynJrAgcxln0dJ+ra/IE1l5PqMLGBWLXx8yH1bVxpljUgZI9cvpU6
z41xTjE10baRezJLIm5UcQ/psk5oUDtZRWz2IEdhjkHse8obu1UChE/5/8FkLz/h
bGUpGVXJKUaXsw/yq1HjcMKAmqTxzQxuc+8jULZX+7hnLw3MtiwjbZ/c9rll/bbc
BGaTzRidO70l71wx5ZgksKBm3W8dfW4PbPe/zSXAukGhmEMmHwF+0wfQJH1W/dKI
aKRj+sbWEI69aff8/36tYDhXUTdyASQ2Y373390Xixb4w7Kr2L+EBcdcJ0lE2X1k
gDlxRPO08c2BW8QeKfcGefIxFa2v894jpJFaWBgNBP48mRp5LjJjxnvk752Tf0a4
N4VRqeAR0LYdPqPp4fro2YgmO945ucBEd3qjN4rH0xGs2eqzImaEjwTvkl4uJotn
ixzs90qN0t5juoUsv1z9E9BV9cvFeRhykuoitaxVyVdLXsYI90Qt7i3xbFrHUOhR
KYuQtOvKvKGkKI62MZr+OWzxrG3wspvehs3XoYIIOz1hxmrrWcgYn/N88CzuZR+j
Cw4G+OuGPdltqyoU+ON5dj/78L75YBa5Bo6PzbdePzi2LYIWAMxOMONGJ3PzWBRb
i7uwANKbtSESVJxRTGwuHLMx3vTEr3kfXIA9pQJsQciIjb9jzzWVRiv4FjI4r/PW
KzW8MG3NnSO4qWoN/WN6zTfEHOS8HVvH0Jk9wUMIhbiMT8clIRacrC08fYVKDnly
R8ZmGCsx5AQtVAjR1j6PS1vJ8dN11aXOdbRpC8z4uuJNGFkEbCFRhb0J5i72blaW
UMFDGgtLy1MlxUThZLpXIHl+391+Q7BfrEKunfX7fk1LAtlmllkkn+2KT6S/HZOQ
ecH9wv3GqbX2OsuQL89GiHqq6EfOmbsxKNllTpOKpv3HwCNMjOTHo0MmA+AEKteV
xZuc/YEQ8EP0yUPZahKWu0bk5cVbFK9XpRpKCbmGDg+l91t7N195htTkzhHAHLSl
TQ0r/T8CxoyzEUJayvdrq4FMA9X2Pw6PhLtKAvkD0mQcfhWfCF7+1l9JPi+Br92N
6RdbktdgiGXrRyTNEn/txkNobA8bVf8FQTsv3G31FGUji39uSGerQ4RFrQ3NmTn4
wfgpJqMaH9YoVdkvj444ID/irDGC+OpZIaSkukKigBjooivSnYjQ4gGmy36tAOdh
HvYUfkTwFaJEHmXz3i1+aOl/kB0Pp0aIKtKR2EK5BjP+PKoJ0gHSdMrFsr6l9qyu
IV4Q8JXpaThLppEXyMAl7AUNVR950UHokUvyHuARwmwVOjWlj7f3Fmrqs+y2TJVS
9WxwppLf4QtubIpWbS+0RCfywstaeHWeKvhb1RHBkPamTXgSXra0FBEbDaV6YDUY
wBSq2fXyvF9BfpazITbPp0t8wiqleX5FM3GwP1UG9zGIJ+n4j5ZIuMA5p59TN9Gn
spn3A68HbOIQQuYxrc+fm4kBZLQF7BUO+QgiiJDXzLR2v+7IXrs0hMDNSlWcHB0+
pbkI9sXx8bg2y0Vuu0odp7W6hwfD2BE1GtHqvboOdAt/FgN96dLF4wcM1pcQSs+m
ECcBHy1Z623bRbbNdqKYECaLgEXJNkuNFbdW7IlluMd71K6ip6z66AGD4KhJRx6P
3vH9Ty8364gO4qegtK9ddHWaj3UuP2IaLHyuLQOjVtQuSwMmXbHO3RznkIuqQOMN
HnOmt0ugJyaGuaxteDQp1UyKT/pKGcfjD5jJSrC16fzJAikZrWCLL9jRyRA7w2L2
CtBh/NgyDkCTR6N7IwecEpqy/XrXNw3A9urH5mOccxUlcOuKawUR6cNQIHq6+AuF
7I8iHwjtl+Lfo/c2nIfVqyzDqOKpd3Q3hBfh1sV9mBhbVxQScGjSn88ktq41AKXh
esDMu/1RvTBR867m/eusXRuG9CfxGqliOwpez/y2+Vuiz6vLbXS7lNKUPDi7zk6c
w18CLVYLFcKgIENTbjOTUps1B5tmzD/vQWV7qAlh1ZKuJ8O0sk4XvX1kXuPj5pLv
QYKuoVo/fVBEvVi3RZynj5qrKzl6kgeD1QX0cV6V6RK3twcVpJeYAplXLx5eDqgh
5uOueE13/Bp+936sIBPS5sHhRkZJzFGJ5jCx/L9OUDKkUE1gyo/R3BR0/gvk4zST
c/CKsgqSaaWVbeoi+Jx5gRVvJTrs0xZUr3sBEEGfd7H5MYM076Mc3IJHw3gh4nYj
uhWtqJPg6bVFAUGipSVvxPI78c4SUGGEdoQJdpzSe5v1vTxLWqKKI1Po27HjAwEH
88a94exKN0Bqf8gnCWV8q484bC/TRrW0m2iqoYH7GL6uuEO9URmPO8/YNJ9Dv6gn
qfq8euYeaVyUH5QszaywLEY3rpp4WuGE0ORqG6OfE15m49nNTR6tExaV2JtKJX0s
08vUqZKkMlp0iaybcH0+ERoHYhAtG8GHt4xVcfI9Gxmynk6iR4BnvbrFVUikyI1a
eQBFV2JQRkvuWEEm4Nk+/gOvHLVqU85fP3HdbrRmQ0Pm3NGj+cpvdB7JHUxXR5a3
ktXFA0shg5XXuA7xrs1oqFiG+y2xo0rpS9FViA9zMLzi0btxOWhroG1nXpiEHqtl
Sue2vnD96DSeCQhWOk5o77KVqrbDXZjdLzddoZ7oeaqWik9sVTJpxr+ryjO5qjY5
8nuynMk8CVAKN7QqAFs8kRC2CFCmyqI6xpGI5f2DG7b1DJrXUbXcmi+tUxDxORnY
7Rk4TH9aCHO7Ev9MWKfGwbm8g9adF8rkDVrCPewYlxKTmHRggFce49SMmyTdGxej
keMDHTqGeJ31YW28zQd/FofGsGPW+qWOFf1+2sf7C8VZx8QMN7iPwTO6cQUa/+wJ
+prIsozA+mKRACBwEiDrwD0zS6aRpe3/ojCom4IF0Ji9PALphvG8wbkQHWXp4C6a
4FFY48ged4H64FS5XsBQtWT+yvZlV9kf6HUwo3Tu/YA7zWUUynZDf8/mp/RQcLHj
Ez415G5bp7KvgLHfPXZys61i+4+UJduj1kXEpaVUiBbroxmfFXKjsReC50Yjt8mX
juxmCk11SfIVCJcI8Z6yiwVA9G6zouH0cZOjP2GRgAMvaR2vpwdmJU0jG3gfX26U
jsEt9kibfkazUwAouUpIbyrTW1eCKovr1ynTP3gDYmVojrXMp0sdqW4/t4vYFmTS
7Unth7/2SuiwjuyyDR88prhhrps2uI3V2jPUGFibWp/ynsgD4E+He4HJcnx3BGgx
VMlm3YC5nH2p0ScT+BE+IDes9ds1QKr2BaH9Q+qSkkWw/J8vbHLRM8aJOcjLhsBF
m1+RsmxFrJ8zjbxeiHO2z59X+/ykmazrOZNWRMLd4kQzUaNIBh9XiqBspynfSgRb
z1IIOgwznvYQcLugDH2LoFya7B6S6T87O8+cm2gRMSVeYaMA/DWQGF8HUlP5Gp9H
OpCP4VWzSh60DGLTywuIXwWgXqR1BKGSS1bsU5XnXxUp/aivSJDWfACc7Ov6+4xh
dXGcUTwfNgfaE0cYelhbcbMT6vgAXYvqaJ9IREBunLzZcOucB+vUHFXFBGWCyKlC
LE5FJQXHJV7KCq8Qt8HyfzW7sXMW6QQZe1FxZRgDWxgVSKdXwS+e5g0VbdybhFjR
oEcDROfGV8k4p7V8AfQEtLHniyFjTcvH7/SOfJSGXTLbsQ8hpK4TGfihb6VoKFT8
zKZXQXYe0XUwiwWX9jkVn5Jliy4f1rkt6RcXbEMVlT2cmjL8triSmPnh7FITTMMo
RtjK7cObBXDfbtL7S4CGu+1+Bqxt0ROw6VVYFfxX2LvdMD0WjR5GpxPhdUCtGYrg
szvzWAaoi6Gf3ilY/NnL4UmsN0oSePWLxMUOBXJ6fdi2ogEM7eArxQeMFDsvcsOU
3lsFomQPP15y75lZHBBaj/XoZiCEklXoo6XzKS84shXP1LVlZnMOpB/8R0CsJp9D
HqfqdbVm3DePTubJcn7bYjyMPUhBxqmFGXo1LcNN29Cwd8d/uM6ymyB9FYxkBH/j
6pMf1SjEDiJ6THgRaWnuvczGydYkExTHByOwb4jbTfHxz0u3vyfTKlcQWw8I2yHp
NlwsYT/bRJW+IY7bpONx0JUniQ4fqMNYLYmJDG2YFPgpA3Ye33afDLRQQGw8sPFz
Y/7nS9Z3fcLRoB9sJdJsHXIl48bA0nzWlsjDkh9csG3RbHEmowdeRQM77iffXDgB
Jl3jcaa+wdgO7KPyPii+Ny3tFrHr5+It7XP0gmXdIf3nPLVpNb7V4iT5P7oJiJbw
B7B5LcfkrlUiftu/fhDJEJzlEttJxSYo30sGeHkmGYZhoIPThtQsTNdl4UtD9NbO
tJH3/paIzJBb/bOh0lTQleoxHnbaePJRJPL51mNIkPgVi0AR1Ddr56hbQKH5uIq3
oznkSz/tkPlSxYrqLikU6fTbb/UEdwyN/PHCNL7gA9V3tVi4hMLzY0GNTbguyzlv
J7E1tlF3yTozWkcaoGL1UIoPiEkXrW5JGPTTRzSUosiY1qUUMYum6Dr507FaYEKn
PbebqP8cIaCKKGjF5ilWa8wyjVuQM5YTFfKvgNGM9NFC3g/KKci910B9u8DsoSbh
BqCCWjvOZRtVRK6QtsPAR9xJb/4UYox7PhM8Skh09Rnmg2QVfS7IKDRCrJbGH6Kf
oNdh6RfEOw6DAyXt9cuaSavwzCTlUteP5Zo2lm+tdUG0gBv5uVa8l45N8QKt0+Nc
dx32ZFzUhE1OTj12k8C46arbWOVv5rc6PsDCDBSBXkHO037E39sOQLZQehmycjqR
HuPKXA1Bp0D3Io20HFPqrvEUjiWEpKPuRaRoIjhkNOmSvochTXrRR3zAxfGmLwnK
XMZDDz44M94sQYLr0gi7ElnH5peVDiOcaOkazRnZ0GUzbnjsUFJJ9uEFjvmI3h3b
NTE8jSGlfer+PxXQmyK69/V7DS9kHyl0O3gprv2cFphx16/uuuQYMc4vlbM7/lia
kwloK8hauNIDzDDSf+QF00+MFxaCxQXKjCoSa8jAqSB4SqQIY0tHAdVIvl855oN5
8tpl/VUoeor9V7JKr8fOuOgMrcUsPLsQmF61n/+QwsY79/wzlwrCUjG31mQhcedi
poeIw5cd5cVOAUk7X0Rsjp1UpmsGDZ7KI5h0OIMCnMa1RnUWu76rwPjo2Uy0eS7z
8c2a/QQSfXgaR1Q0HAETh8L5MGO1hpLAV4K+3IL/SsTWq4TrVMC8ucNgp51Aof1B
iGIzJmEQrfkcnDFnkIMDocYfEOiAMoJji3f8g4NoIeOVj8lnH5KjonHATX63z5NI
/hQOzDsnJDDS5HtTypRbyAOCvPQxFMQRBPqBDvg7hY0FyYPIfjpXpIN3w+S6WuUw
I+lKWUNrvgoNbWsa/4V2JUoldoLMR4h4BEuOzl6nJMNN6ZiU+b1yS05TsS/Vvm9p
hA/+1b0ayTofBGiH1eeOR+uNRAA0w3oK5jI8kFag5MmR7sq9jD1snub9zYLZqu1q
wdeRHuQrX9n40EfR77JcRdqn0F3puuWcSDgyqUa0L87zBHFlzNzzDKcFyLx9uJ50
cyV+bWMlAWLWcZal0n5PD14UWVQ6bBPB0RUzOtHWFGc7zcAqFNRkQyVXJIRRL309
kWr2nuN5W075BNJlZ8WQiucI9qZxOrd3Mhiv+gA/30XSG8YQ1WwO8no+YSUrLK89
TxTT+WeHETvQugAP5j4rtJKBespC8XPdowiRYgUTsyed82sNdnvvRvgGsyP0O3d2
HWzSFtUyxFzLjBwTI4wHq3HM/mhgm5q2qasroy1wC6LhimeshnpIZs6ot6afak5B
pGITg1d3VUHwUaaNCMLjzEgI41DppN5Q6FMI0QYxuxOengWSDyecHu46bXdDTKTj
czn4zuQo3maypx2KBMNXjMb8IhyEfIIFM/6WRrrBqH6gfWqFnI+G4Zs04LoQdFcL
snrov5C8MyuIydr6UPnLzc7L8tS2b2fnuypjIja02JJFm+i2ukKT6mEYF0Y6fusV
Akw5GnwoelYR9sF5W9IOzZXViCVq3bcAU7aXeQ0jOtHRQ9sy+Re6pIGgtfMWcHay
+Il5uv5r2ZRv186OgkMdcqc4qnI6DF3o0A/CCYNnN0EbZhTFFzZlRgUaDg0VBU73
7md4QeHPzUxuyORkxklPYumv8+4aCpQkxSZK9EAbvyrnqPVnj4lqDJ+i78FVZRLO
lwtE2A8fizcROvPEwk1rxcOIsqh1+Erikfft2dL7l03rHmpcujfo2oEnu1a8Wzi2
6Nrhq7YXsqV6n70ijUk0Fv7cqVY49IsZFlp0tm38i2WHVeuP0Wx+KQ3aNZnfz8C2
iLb7PHBipsfAzx25QaJTcBY6DT/H+o+Lo1zDKoPn1YhK9gzDloqUo9ZPtfCG0pc0
skYSOiwUrQfLP+76gb0Git4eCb6V4YOjH4o972tHS9xu4aK4THf5m9Xn+r67AROW
egp0PWUbzbE/FdSwUmkOWH8vfEOloBMaGY+mGZUJY2DEkl57+RS3us+1/u/oUnrD
gNCVmkepI4VdF0j19CczVDL+7d4MpD3rKjlD7XaWUPZyn3PZ2AWR1+yAZyi6McV8
pgWQ0+fOl0yXqs7bBuuQn2xwmjP+rVOtn3o3/hq/vhU5jt//oPoYnPYhSPRxU4QB
oj4jgOjntM0snw3hU2UllzKZEw415ToKnWCHDc/awwuTcx3CaGTWWY1s9iDwCch4
ixcC8oEwdjmV9NPap8g5CezN5BOZXBXTi0uiwfnXzSA/jJv79za+tPyyT7kuZ42s
IqQ1LBI+KGqbsR6sJrG1pYBu0hC2Wuwz4ire+orV9iwyBial6sfFd8TdOTHS4Lx7
sEcR3MaM62yD98nKbg/M5Tu1UHoMswUX7dgEMq9hKIITZBj8IossKytvxnm4zkDA
57XhdoFPAKEKi48WFelndpBxby+OC5RpAoeL+44i4Fqdt0N3BVNVAitum9aa8jbm
UnzquHvgIE+6H0KylBS7uCvQoWyRUiGbYNQa2KkD9TJs1UyBmb7xur7zBPZUnTvI
05aPboNIY3Fn7mndSezGI7piWXrlTfry+Tctmfj+4Wiwk6KbK1gZcKZlvtmUobTZ
qYq0Ef3KgG0wvghluaX6uhYNJj493RLDttvg1zGkZINuS6nDnwQJQajG2MKTqaQN
QU+59GpbmjoGRhm32DTVlpVcpKebZ8lD6+q7fZKH+O7TGprg9cnwV/sVycLiG6VJ
gh+TLZvR/5GuREbW32ZTN+R+x5grcTnDbUrB5Q6wc6Bbve1vz/B422gI7WUjvnOh
S6UQn6Rw+mn25Yw9ObK4LE3Cf1KRTIkHSM4wX6J4YOuA60967hqJV+SE/1Z2OM4e
Hcna404drmAUrzefyn/tbJPq9242JwJ+vjklVSWS5jN3dgA/J3t0dJrnOh+IX4Y+
vfCIZK5P2iIkPWF7mOz1yPjB1gYqllwixYoQfgKiD86pwzKvBuqHfRldw+HH5Ydq
Vw0skqoDQEsZIZaKfGzp7dNAEzO+ylb24pZn07HFYbThaQwVIGseSRByDrGLvSOb
b828PHys6Yxte4zrQZOIcgb5Rs4xRWCV0ek96aV9VFp5keCYzfR2sqY6zsfAvOif
jpnKj3Q4rjVyjZ+RR3U4E9NlgyugkuV8kjXrBCviBHwF8GZgLsPyRIlDGwlsGb4e
4UlaBWibcitwGhGUXdW2ZiHtgpXIfCzr4FOswmdRC/emQyHOkNuKZ1a6dYCN0PKc
zYd1BG4RvN2uIKClE2W17lQNMzdk4hjKAwpwv1SQxfgRQ7ehl+SXfua38ZQVDKLj
l2Z56XbyM+AcZXxPxcbkJuGd6NraoORaJqmJNVK3QKUo1mDT4ElHEPOh4IZhMAIi
5MJ/S3Pct/toHIatDs4SLhNYBzbM+BuDmq33RqykYqIpCmtpigG2CivPV0NDe2z9
yndU/a9Z9Ex12UMGaVJHAwtm/4P0WyvxgOCcjLCyc0qmGq3boxYRowftnjBbLMMK
XX7Dt+Yq/DofyS9y8T4LltowKBVDxh5b797kiy3LoMc9CfBL10u7i5uaT8MsXYpo
2wT2OZ1LYK2TONsnuI9xOyZRMaOe1UYGxhGS1svtEfJvgnELdWhAeNXo1eGGRbBY
v1AIYLsj2yCXk6ClKIvbz1RVfJIi5yP7pTMHlfTib98Rz0CN+N8CJ5ll4u07q/Xi
C7CD695IcGIasQ5ZvB/Y9s0RksSYEAl0YUWYBcUV+BCGAJjO+Fai9b2FT2bNiLUP
HETZTMq8U8kAySOJCmixSBZoEdI/KQM18Bh8krokg9ZR3ARSfTT72/5BogdhY8xW
d/9VbPsenHNbJADPr0XtZLMQbNfYPeAPvNC+A5h5zZ14KWksqzNulyGru7O6Ny7J
lYlTfnX+HAVgPGYDtsRxmfXuVuix2AS8ZXlqU00tjv4Fta0uc3zpADOnn2FR+Q5H
qtHGAStjtFMII2o/qNqOAm+hbkzpGTJrSXcc+GvFBYX7V5hh3YaPmUpygwSswKMb
krmX9hyK14GWVQMbEdW3mPO8ywnTpPab0V6FjxLk9ky6MXqBo0oC1BKkxvmY6wCD
0H7u/78ieFfTMOW9T+/n3e5XJ3PfgLLyuZIPmBk5lc+P05uottFE9k5WOlgfsx4M
3OH4n7u9XX0GNCNbuaSIYOaYzw0VYZX3/k2iff0cHYzA4PlIfAj34/frXyHzGr8i
7X95A4npBpTOqGrL2XAxZG3UZudyXsVo5V6Upe50IOGue+J4Ljnh8DcRw/srD0Nl
CerSaqeNO8xRkSgFxzyQzfDKCPbggXZqamQkGUtLAdM1hcLt9J2mq5qMlprTxSks
NEUsVUfNVwbZ+/b5Tp6MkiDyH3k0VBCXoxiqFVIQifyNMU7+HbrkIsilu+8COtSa
stSZznOOphhxbu1oqb46flz1V8VuM6zLKbqWorEm33levQm+LJ1TnUxii8qNSH2U
eqmeHdjR8VfyoK1v3xbzk4sqN9flkXS22Cu7+SGvEM4WeWyIG77gc2wF9UwsI39l
JMvmibaylXcYqE1TgctMMnJ8IsxGIXEX4jhZ/cmEN6SV12eRXyfrwD1LvaENhApl
CzjTlmYS7/0iGDY6d1Uhlab/UKTFloeay5nJ3sphBPow6cuqnltI4PUqNXo4JExR
SvvXgtKKJIxChsd2xcTDC/B+wPi1Bdt5XvwXxr1l9xZGRyZ3z3AZVapfnVV8LiOk
yksg4rQvdV0EEPtkWD6O8esPAtto9HV+WqeyXI+wugvHWKjcipaTOAfHcmiHimBR
xwbrYXgQkcMsEroJRC9hWCC0XNxDIQtzdJTNEGEPomxKDBd8o2+EhjkDQI9wdyUS
aVVnxJy2QTFOABLmOMKHg8wQiRMIFrFa/jpQFe0Cwes4YRqTF6q2/9r0hKfQq1UP
2kPomRGvA+ChEoWwPZbmziZIqeDnRyZCpYn1iNWsO1nWH9TYp+0mYEaiX/h4Pi7d
Bt5gOvIFWWj6og37mfWAwKZINBjdBzs5Blc4lV1RiH1B/JlGvpnTcafCsOJMKyeG
eK610r8mfgW5r6orJCIA/l9dNO1/xGLInIEZazRB52s0D4s8NlFhQ/M0MKqEkLmW
q0M7UZY9v60j7UKzxo9NQLrNBxHhCxZMB/i0xDekcIN+sQx4l4XfbIYBZ43bgKqI
YKNLu/w3gpvyac1njAnRvt+TpqW/Jc5XmBlf/lAtrRheMwr+5xFAAM4hzSk2irgJ
95xdbuIozvhxU9Smy8xHfmQioXguPt6uYKlEehlQYQPFOLR94bbjiWcsQZBSnu8O
AHvz57iG3w4yKOV+2FVGtFKpDly6u33CEh/SnoJXDqSrjqwf3rXACqaZKucv8Vvd
iXRprHgZLR95Iwz37bfHMNP/jYR1B0e0eCLPnM5P9w6qQLuuRUEJs0Zqhy4z/XlP
zDvHKD3nMG1Css3sPY18FX0/oAKmhzMha6aFq8oGBRofQW8KkXptxyiYAKp+C/K4
Yp1bsmihYaiVRApqWpDtfbF9kIeApEydyFjkRDja3Pk6u/BF10wIoy0Kuy7ECdCf
NAx3LvdyxLNP6ljE5OUDUytTkw34HnLNxlITDwKcKhmHicD8h6NzEu4A6Qn8ZhIW
zQcneaKR62NHvu7QFhYKKVXucvIPonQugU96+brfYe4sbJul3kp5/FwV1S78R0mt
A6XxkqbYNUXmskW49S3RITNOj8teFUg0ZsaiT/9F4yLzdfGbVDMIB4OH6ZCSEfhB
lNBhFmtbHh+hPQD7kXWrA7+DIX/2RfjGX06MtPWGHCMQxfQv/nAm8lbD8gJJ3YIC
vB2rE/tL7TLmRorrRUIE9iPyfWIn+5neCU8g/IZwXk0MJ/fRED3DJFt/JaMPV8rF
WJfMtV0hWEekEfZywTCkvpB0rCHT8NtOITxJhiGkY2WfePIdQ9qx1N4gLfrh8ZsS
okSOmHqWRs2z6N+Oeg3FxcUePupeE5ywGkFCeXSlp96iydiTLK1l/IyKChjkFi5o
Qpyza+EKMtk+8+a82Ud+tFmeZ5z2OZs5hjCAzdWL8ZMHkwUWjaSoBPXocPgWq/dl
Z3xL2KyzJlV7xINgsmceJOVb6oKmVyQ5nVxdJm4QFfknAUwbLrc9CcVHY6kFbOKk
U2JaS8H7TNq86LU3IW/KByRqZNM4ImKniZYjVx+U3dCgum7nbYBSN20nDVBXRSoI
awWlV5NLgGYP3rdmmwdqkscZQhdG6XruV24WvIfVHnKP0SfUF8dxU0gHUWefASi9
qWv0etRyOemPPsn7nxEVYJsuU8OZdrU0LiZDxkXGcMJwVfN9Q7Znz9bbRiWWkCTy
5UPMHPGNanR0CiqVi1EGdkisHpfGFn5Jt03tQzcBoY/ZmjB7CMB0+jhYqBQ+yhLv
xZrNsqmWQ/ch7C+4vxfWd9uE3yRKntBYxmIqXGgkkWOXSyZenrPqT1mKYHhqc36F
F8NcMH6apKcSj2CAkZp+J/Z1G0CssUZVVLjfZyErbjkfZVNeoqlDWY+F/Yze304V
dxr27MzKhRl8PVb4pKnVPGa1QIUMZd8xmPpMnqqKhqoPL+Eam544+MQaNap8hOgj
nm1dpYRG62INhT4GfZrqXLNDaXiBzZIm+NNa5tyfigJo6DXH8MkI7XtzJY2jLK7L
BBcmoGPY3kxb3QEHRUhNoa4RNNrqPj2GLUyhb8jKFY8/ANlj4ZDQZyV90Bs7fnNk
NO6FW4rNcKEWKvU30SNY7jlQMu86nMs251z5qQYo5yITOgdbQSL35Uc3ExOTSk3y
b/UrVNzi5Crk8TLdSsC5e6/HK5uBumAoSaDth7ZXiSSbTCJlCjwGad3+XnAnyVMd
X8CdUBH7FwbSfctrqCPQ5Yj81JlMSy8XLiUfCILP//H5YpcCNaOT7sDE0D8prf3F
VDWUsho/cVxhK4oOj9HCXRt1SsCbE7RLs6XmRQZAUizxJHgxRz+N7Znw/u0gpL0N
zvA6grnv0D8OmYpIgMbOreyZEGjcB/VB4zrEg4rKz7x+prTjBwWvinziYdyjR4g4
BduM6cV9TcMKP9GTXcxTO2cHM+TTWt2EiZe2a7ivY5ghzwxVgj9tAvi3w3tSdynD
O/+/5MFqC4cm/VQvhWYedIRUPL4i92aLBlSJL9qMKguh1ujejFckD2FlvmyZS2Zi
skOPQXFgVbZZBJchxW1wk5Szx2Ef+2fPFzcwCnUGojo9YGvqD50ifc6fi0xh0Ctb
aBYLdbb400Y4LY+KzpIU3Mhh8a7T9ae+PC2YF1JRS241MgbBay5BwzIRG1naegqY
OYdD3u94sK/ez7UHcmZGGWYztZdPqbjLHebN3CTOJVm1CL7pBkVuChVS0ZEFA4nr
SbKe332XgAk+4/5lLm7HA/ysJtw/FRbxiaKnTeEyNFYyR3591uzFCShfp05gaZ0F
yqA66pTONF+Dm7JFm7ADVJwcupMFeS1QPJ+rav2H8bs274QX/RlVLr7mwGzRPt8d
IRjaJFzcPQXtK1DVBKpv+65fqT+DCxoemQyV8Of3wqCNfy/IJW8knSxMYoboCXjZ
wkL7///GapPGyyx0jweNnxUm+vQ3eZuFtOpKBDDqfCGzrJld/V/43Evqcv+Oqjv0
NNNYYUug3kGs3HezW8c1YVHvn6cJ+QawEEib6gxy7753aMMndCaOZ8PwJ1JZRF4/
vsKP9JOpNYxDNO98JdXwAvLNL0TCc4EOTXkqAXQPL1PE2vRcGUrLdJu9s27MerHz
Fe21VfguEOVeIXDRjr0xZbat7P/hOnE7vRea0YRisa4EIFB5VAgX6ylijWQtz0fJ
vHshqpUIaBFxhICwAqxwW9fmnN0GLQJbOG5dIzl2QCowXIZmUlM5VYMI5P0juTsr
SLw1SjVFLZOknqAJn6VCJAUjwnlgepGNOSWLXMW4mMb5QP8t2DuZpPe+X6JylWjx
jCOKSFTmZmyb0cgvFVdSHzXD8TMu6sKX9sRxN8vnmlIyl7mac9RK1nbPYyQzqfon
mgiLQayn9z2OGf9hLjYX/YVSPl7oPj5dQIQCtPr36fIVQSGlh9m4mGOLPLdaEL6K
DfPL+o+mO1UZZk2lioQJmTjKonZGoGwhrQT9D8P4Da8Rh8twkTfmUxl0GY0HoRpG
FaBGoHj3p43828r9rI3+a9ATC8gLzE4eQ6p8gHBlBZ1XbJ2pbztObfT4/2kvNJtf
FHsviizchTR9njhll7AngPP9TCzG6HKu5miVUQpfB2VSWnrI3NrTzLqS09IFo0+H
RsGG+4zQaY6PGRrbGjlyBAKi1qdi9MoZIg2uU7BMdDdYutQC2HdWZCc5qK0TeYhM
7qClv6Kq64FBFY/jZULLhWkSZuCmxvLLOWzRnTOeaRwXdNy8BHKDC6CogZw6Z37R
Wj2ihhqnxYO2uEQvEJCuPjjDA6AL46PWkfPrGQqaPpyI6+jG97wnPGgE4UjKPjal
dy5kRDHKQE8XdUfzHRdh02O0sqHkcLWDhEdDajIW7iaQcEOGRPqbOv+bN7MqYyBd
BqCGNQzEIRTb1oV0HRojEV00A7xjh7VFBDFjwaqXYHQ1rvUW71/7gAOhXuGC7RrN
9Aw9rAwc1qaxzlJo407rbdZU1wtnNJI/+YaS7yU45OyJxpQnroyZwjnsXYwFQsy/
pUs7SRHe7RvpDiUZ2v478T8eNEI1575pDSJBx12jQRv6O1ZMBB/HMIKZ1sKDkzQm
UgKiuEQCZZ/dEkXalciZFriitbwZ3wX9oZ+x2AlOuGhpr87SvwmOQ3Y8XyNq4nxy
oMhpNx63XvDQy/6mRGvgObWEINK0VjRy6NZryCad4BvAt8xX8/2T+GDqnzqlVJEB
p7pmFFUPAjLUTkFsprqJQ1i393mASAl7MiWcwqUVQI/L8jouhIteCnMZA4eBOjG1
H8lQrRIu8Z4KweFwIxHv6qSVY0e63BVFnOzMVuZbohc3A9CEY59SP4fXyXeUY/hH
UkN8VEBFTmbE2OZSRDQrAyuTlAL20BFGQcQSAQttxmglDUKnF/qSGGPaVgxbum39
3Ob6qP+I9oh8IqWSxpknCZKjWarHtJda/rpC3nH/BYUAZBaI31v0bVJq9S13UiZ+
sL9Em5yLbsuGNQXRGBjpe3l10FfBG6P03YsD8i3SiTsqRTA+ENAzesHm6J3diibI
pPqSg7XlXOkoU/93Vnqz9MRrl4kILdCRDBFRRxc7ABS9Ahj0K/ZfkLRZi5toQB+7
MQZJm602kCBhUTAIYp0DPlpizY9VLwKsYxmdQ8KC64TegZIZjP/OPLjbOQExuVyr
ZsEa0NAVw1nQsIMWobrXM5PEqIg8F1uQ3Ue4DPCVE8WAJPlM8CplkpLCNYt0KzsN
BKVBRKcwoon5Us+5nsXwJ8JXB9DhqmWdkr4VTKBPXGz/RQZPIYyqDato/oBbSoDx
1BP3kA9PZbRNY+5eOHjE4+GQ1rQ0g8ulqKCHe0zVgJ+58THmYrTxy1ozeeEX4sV1
DuZ2oSo423vjmrIg2pzSet5DyyFJRxtPK3310cwgVTauMeSa4eDQeLlVFGzIIX80
513FVBp2Y6mEWP+77qpUMThNR0rPFbyFwUT+9X5WkifN8uUq8b1AvtPK/nJg+/oF
pPDo5VzlsunzRlgnkU+y7KpDx1aq2G+45TnXp25p/j74H4pjmWgbMMTY4AApnh9c
zKbKqyLfGLTLGACsDN0Oq6UNzXihNLOg3cfgTEBnNxdY4e6I01rhHR0mW+QFYbYj
J6j6rzmrv9ZtTXMcj3kL7rdr15lFaq9VBSMOcSRpfDPLImRwTppRnYSfb1HjkLWP
XurBzVkYgA2BK8R/XtkCJmEyu3cyHkFWtham2iDU43xiiJLmMjbEtRLNP48XnXlI
l0WjcNaq7znLrOm35uV3yl5BVvv/rr9rFytb3KG1LHkj19cbPsek+jAaSptqDaxd
DoZQNxYPLDrVVNYKPUe8uDBuLW3ORgWNtOTd0aYPZmbynSnyjeyGFPd3VfgwJUso
bBrmbckA7BibRZCS4trJkD/DMSrnTHNVptON7BhCxogXWbbV9/JRE+nh11TVZNZ2
Vs61TXDGTvr6Tu33uC4mFxaZ/bNwvVsODL1/NrddzKqmlQYshaq1D8S4a7e9lXIC
ADNkSrE3KJRMp2ewxt5esayH8wfv1WgwcGqvgijwZdCzjYu3wkeztYd1IG9C1JRz
dwm8RhuRhQkF5YSD4nygibJoWAro9x2J+WbjCu/CkgZwGohvmY2c5kjU43vUt57n
7MluYyx9uI/A4jnRJ3ttpEmq2LGasYtPC/gMNi5QoSQY1RQvHZTXlt+vhRn7e9Ga
4A+k4oPZStRkt0BWDFukA8RAaDyfFJQSd57yWGWbfCpOvvcrm1BxNUE9zR+taGt+
SlCQ7/JpBZPeSU4fLOmM4DTwaiZ6v/odeSPMEYrQLvX4ELVnTGelBoRM2md/v0PI
1BghzJ4ucm1vBZbO+/lKgMGn3yreuf/uvsNjnTO+hHgSwnQ8OJh8cIftGExks1BZ
4dp4FWPId4AVNaWkIE+XlCMgan0YdOud8QCwsk20eTEv6yHG3X5lm4+kiPiJPGRY
Il5C3zSpNhfKGjngDT+OipJi7dY/7mD8iNf3/L117TMgJMjDK14JAiXhPyyKDvOK
LF6eJd8vmLMJ3yQ6wjhJLj8g7HZolqhPtB5miQHLscRVwTudq3C+0PVBDmHq1ZpK
oGzwUqQmyWo13ns3uBxk7Vk18jvey7PByzjYPy45GEEe83XG8/FYgTCI1paTQZLB
qdbuqi1ReiaCsi1UbfRyi+EtvkFmqgB0B1dpp0z8RBlLgUml4H4hF1qLSx6KHiYn
5foACP9b26WRK6ZjeCIZkfa2Um5yntrgtqFa3g9vaq/M6hO1HsYMkNLetU+c0Vcx
SqfzLexoaRGTj/G0UJwfjD1iir2H7VUif/ZgcawOCDEPBUqb4wBZIX0Igqtdmhke
EAXMLCWmB+i6qfSWQIiNaE6p8Azopcep1dxLJBnwrmLO3WJfPVqY26ObG6YZixSa
RJiZjZXiK6r4VjBOYZAi9is/Lcv+3BYFyezuvOOA3OjNa9zyAyBtvUcv+d6Fa7F0
HSUYXgOhuemtvgOXYZhWqN7Y9Z/WWLmyjw9OdaYiW6vN9iEcYqLWD1KbnKRWuTKz
td+UWWVA3qwrZyfBBQxjyBFthXbLNbx0bfXjsphoi1+lZpfcx5i8c0VJe05v2RHl
K3UFxJNs9KvN82gKuM3Sp/LcSIblVsEIdgZt0mBOqPUd8TvDNajaP/WV4FscoXVs
ghictOntjXYKLnKnLb/WMiUzMyHmsDMWby+Z46q2O3NrCb3iR/v/KpdCoH4K9JVu
8VlhkdPmnNJyXntOeDo6lySNduunVz1keukI8Oi2VKlmXGy9xz8ZhLWdF9mHGcht
gwBin8EDCrsPPYrGLeJbBI1iHiclwO/q0LJi/6a54j0R/bZvhdQXGLlCkzPRvFde
ffQbyM9fcj9VzJGS35PPYPIaQSHSxlGBRNc7yTru6NO+OUrczltl1AtFjh/ULSG9
7Msqqu/jivatcxMJAbsoYUIw/1aw56C/dxRouNRWMcj3DhZeJk631/8spuhyk9p0
Ge2BpNDYpB+fR9Ll2dLSnIXicIYBFKMDjjfY7viyyi/x8DehNHU8/4R5ZH5d84tf
/IzyqIx+Dbk7I5K13hAttEsv0oIS6txoEV4ztlKnQLgSs7YGZRmUsPNiNC/HnoZw
z9Ve54WetRerFez/X/y+sTtvJXP7B7N+Ui/4PokgWlqfNt2fkyI01fdcrbqyBWo4
Ut7LtbK0Ri7nQqZTtDeLIzyUpFnSXyAeoNh23YIAr4CQgBEDFD/Tvvmq3bCtJAFO
gAkIQ1+EuJhR0E/tcv38hpVSiNc18CdbFg1X7cUYrLGhLuiCTSawSOcXZrrtSpNH
f7H0ms3VW4enfDCIQBydOgLMBHv0+EylhNiJ3Vcy4lZ1rNikuD66wW6Bo8mtzssL
+cWy0+QXL7BDUQnshU3l7/oL67uNzbwqst0Wr7i4PUeVhL5bHwEpU+76m6LrO23a
yKNR0Fls7TUUhgJnc5h+EVhYLFs2zPr2Kylf3umrHovl0XR+RJ3OrZIoz00cGQlE
dLTCgddre1SavV6PbVKVOb+vpMUKORzQGizczPibIa/GJuPsniMQkYRm8LJs1P5r
9VU1preHBuhFIEXxIBl+dMNJ6OR6HSQkoumI8cNh9AhL4odhD4sfXjKQCszOYNKq
1CWzMQENZGCjRruukLgOlVmkGlrWlWcDhnxYGLjaHQgoLLnW5odyHvCcjNpwJJen
+gNyZvRkUpYuqfqOGCzEl8EOsucthNbtp5d2BdCp3Ns8QyFeef0OezBYRdA0n1Ka
zkfpdjWZSySEb0rAIVYdpAuqwt1f3CTsEK4/Kakn8HbseRM2BEY9hsIwcBMpQQnp
Nx1NF3mZw0/5IqoSNfTktsxdvMVk0DaOn2qbbRgcgZI3h67BCF5Ad9n//mcUv4VN
wXysdEbB6xuVdLTI5UT3Vgyzfj4podb66LZ30yQO8Ohhjx10Y/HaO1fTPm8JIXr9
zMhZ9/FrJRn94qiiARLKeWFeof6e0anP1xNfybazB2bHmHURAbLpsQE73W5vHKuK
q+CsDXf14dmMK6vN7SkGhXJOtxT9tV0OpiUhFsCKexpZ7ETCcA7rqAH+dvjrP3iS
+lMsp49feb6WAlmIkstuZE/BRXCQKHOXNfIoNDbN5JT1SWnkRaKg5N63K/5AXwpC
u4OonEm5roGopxvXc6Wr89BNblljxDvrHI/7CcCdArv+ly3uycPhZiZXmxYps5y7
J3m1jOzyQWDgBmTVELbbBYSeZfl3JAP875XFMuQAAkIOjcwTxn+awHSd2tNez8bW
bo2Y8xEH7FEgnniFHxNUVGNpqldMW5bMDanj+FkubF1NXXW7WV6vCuljOq81tHU5
dEMbpyrejKewVc9SNMl2TeZFUjfuMSIPIQVQYbGvd/LQbLBCMa45CYXRCxN2e5Xv
KDpfQ17STfN3ea4/Svprv00rt9UEHpf8SESl3ts2ywQskBg4FtGb0hnPMYuC9V50
Di2Ui3lt11JRtCY8zwDi23DAysobIPLaoj9q+cORA2Sjq1vIXuBldO5+HiKnL3zy
L7eK5pAJdRysdqLpMdgOygD/M8taE0hg1RFx0+z10LXgn9MObtd7TbjakohZednN
jW+SIrDw+36YoTSTrv4s27K35vgijgj66Av3uLqhMiVt6FJg3Ygt07HYBtjV7e0D
6kP5L5yyJXST1PBrVKUF7UTW8LJ3mg8VPfAAnVjRfxFSwOgJVDE7Mzt9Gd4Uv7rE
9QKKVhf6rZ+tojUH9c7TyyWRwMF/RXhJ+dIgc5BsQqDs63BwSZ+TvLI1AEB4wrrN
7EwzEjlDSpyjpNmw3/IwqCcNZU6lILnCB7VWNDtJwUc5ZDq5jRt2bAh4y8zyPKvs
RqQ2wHucf9SNd9SjiOM+51RG3oGJwgA7/W0GxOilSEsXUYgxTYGeNlnLnqbwl2oX
BVp4bZUqnc4QcrK5uhH2E2gxa/rzpHDNUgT96QC2RQdrsJWQZTyCcYpbVqo/mny7
GzaBMc64/czGjWzByyMdDGhiz79J2gUIMgJHkHlvNt5dQEggpVlJx+noa0yZMvWz
ya7VNiFDja1ZJ2YXpXGGE7RfvldPWhhij9aeDIzAgbNb8wD8Y9Pv6RNytWooJc+e
SKvOUgpbwoC+lcXONMI134tHFSLm54luF0tQayY8eAfFXDDnWu+O8+sk0Qkus15m
tAxM1c77V//HPwK1TOLsK8GFkOyfXAvtRRPKnbXIK3xoM7kNhvgZvM2vxtPT/Jxy
xSNMHgxw6ji/zdzwcETdQB1wIWM/pbOXULQMfiCOYNC50WfhxuTVlBUS14nsUKJm
V5XTacH/4RnH08Kzd4yoG0S53b7yMkoQXnd3n6pGtrplmCKI9G8Z9ewszLCv4jPO
ijq9RKzWBBLl+/qL31R67SzxazO92T46PJPcXUdogyevzglNY8S7SzjGiRFd1r88
siFMYUa2SdsIR8JQw+zcpCZ3ea7B0YBF2zKBJ91QTd2Osi03p0hkLspovDlFc/4s
Lxpq7cevGXyKb48igSBqr4QwGbLMYwEnqNHafbdIoIbWz++uNx5icaFyONu0Ti4l
rcsjO4fH3N2w/92eXjL/qsG9SGn3t9UBS+VQOZo6v5vyj/Tw/1A3ksQiFMiYIqxM
NBTdF60wOPUdzzak4D8Oz1ElwVjtgJj+bZlKawwu9RTB0BnPo/RqrR6yk5ZvNB5A
mPZ47yxlr1wYSICygvNcG7BbzIqUf4hLSkUuVxVmmaT33U1Lvz+Nj18XGabXVQVF
PIps5GrIfTO0uLLJvvt9Yp+OgualgJ1boGFxWosVXvH5rde4Tt8e6Z4myHMVaYbY
pjt6gbBLsc8VPEeqmcK6xfO1vALI/UR5sj3ZtTizMhdKwbIY5S3Ql6aDJhJU0Pu/
HUSn3ZPRvgHe8OKS+T/+9NMgtpuOBDPvCarw5/qyHZkP7X0ZMiIFeTczz1Ips0fF
52G3qSyFCixrY0U+/wPyHoJ9YGHhLzqfOZuks8oOZUqxsoOzFSq9SkfA4q+gf3by
LI7ttrDZGsLTy451ySH5Lfw5BfqsVC7QOneV7YCQHZstRaH32FTc574JbprDSBj5
Rphgse2+gRKax97dv9qI26TTe4d6v7+A3S9UhYfl5FyU4CnFCyvb3bQwbL/cWFoB
EU+xRaUXhTjDuGNfsmUJjut2u+pKMytqvU5he81ZUkzlJrLgZ/j8qCXi0JagLcdh
iqGDI8U+PrH4i1XPMEbGsmcB+u5wp5J3aJwPzHwpEFR53MjM3tgmVwjVZdAEPz3z
g24LCQWhzRSXC1Bi3JUhIL1l3vceg4bQgNXqreABPd3F2vVqUi/u6EsbhBQh1PhF
G71WLYabbskpiTvxohILpgKyS9QazrM7oXNZqOF2tQtvnWkhZvat+COAYd3HEful
OCVrRBINDS5OMnv63nc4raNCi8KqKc2xAnkLII260hr4JkEEjjBmeJplC/VpjBIV
VEL/+XBA+zQcqHbotrLWo/tFPz+i3EzPwbZQRcaOW7h1sgLQf3ZHIkfg04gYiqsJ
BkZRMpmzIchbJ/9bGzfyyk1EdWXv/GnhiNOfdV/yXhPSyVhA1w8qZ+ebzaz53Rhp
mfU/YzzmOMrZJtZUEyIHTClaeZgdv5FKhj8S34pfZUkhD0lLlQpTtEiNhpKEzsQH
Tx3fIF6CLhm2iN80oK+j7OK3LgxthxZ0jH7V/rW0Nrw0CL0ozF4VUpCFnx3aGBEh
sIpTJ0BmP2zm21xgax/uvsOC6/xskuBEc8so3O4QrxiYz8cXYDMG5Dtpq0KN48Wq
E4uhH8r+6DprFU49KoIR9F7ZhMlQqJsnQ6J3/V6FAVkzcJJMBqUObWVuc7Xp0A4h
5FtPDkYbv165E2Ne0xZ0XJ0+OcYsR6/SQZWEWdoDdWiXLs9Ty7GLANmD2Id6WcX5
c29lWv6rBiI0O+LdhEbvLxXng0q7dgzyW96pg90sTRD/EufVvD6h+o7aWemfEmot
Y0zstH5BCgBn8ulCejQyyemJIIy8Sziu2rcNbDqxBUu3pMe/fHD7VJLOHYl+jPJf
B9pOi+i1r5tfXKxgQC34Tppxeb8jAjdmONPuIXPCpapfSzMq7AyIHNSAvjkYhdk8
eqbtGr/bU53744Yt4RpaIETGU1v62Awvrb+ZcIUtub+OM8OSv+9VJCS3gO1x4J4v
uWOG9TjoQdCAS5gXYlmSI67crksc0nGW8KIeQRSePQHarcoygsYV1IVIAA9IuRq5
tcpmF/2cWTeDCxy50NtOItueYPDE3sxxQz5h5S2gNhRvoNMzEp1MzNGq6l1ZrxVI
1nA/3ohIfbbAK8eZg70C5GuAr8C+y4a8th2jIbX6ArImQk9doF5yztSEbBvRe2t4
1d55gI6RTPy7Ypm5AbPY+sBz63Ah36ObKZsrSb1ZOsyQ9KQVTGIsHOLmNb4JdvzD
luQTQKsh34RsrbKRScEhDU6FOYzbFD88TFKBaw3ftx5fsRR9JQEJYFavKIEcG+W8
QEEE2/jkSlIF5mvh1vvoY2cZFIfc+M3vfrfYT+o1jpZ25odPuYeKfILfw5zpJ/Xv
BKR0o6xjO5CagtYbsPqJmS39QbIprhnXCu7R4k+i07Zxgf59H7G60scjwuDBSWC7
GZ8r9Ikq3E4d52kIqYODY4bwOdW+vPJONmnyxb9WMpyBMW7dvNa5ZJznPWnpUjiE
w51y1ZmkwNBN4td//iAKluiNVr2wOXC3lS6JkKW+Rb1UUa9L/WFA5fE2Gi2K2ef9
cZb/KSUnxvv8VZAu8DRwlwCP4BwjTOxA0HybhR28+h0yohJL6tIl6MYsMCT7GytA
Zwtoh36v5F5PKSOvqwJwKzSS4KXazELf6+G42ZuTQPy2rOfVuzd1flpeX9MOpQ2d
PRNMrMh9W6hHtY4JFHRIqC81QLfvfYa0Q8+fQW15ZBiS0TD1iIOyfvi1fmFiguDe
mBVVJFio5ETxMhy0J03Z44OmOG+e3pp1ZUWyUQZiGOZ1CCCOdLu/Nmwl57rNXlAI
QQNinjLBQv9cROwGkuvtwt/O7di2UfukMyxRYV3pkmDuKroyOOXh3G/so5hDKpuQ
r7oRkSkjhsxhW8zipK4NBIaQQBGbNWUxkzD/vaPE/quF4Aa0+69w6ssf409xvACP
JbZ7C+6pPhQQaUtAqikM2cBmE62OYk+A1vQE/pL8MHAwmssuXQ3e+P3lg2Iz+PRZ
5zf819yRVWPNtBDjQDXk2maftYFk4EOP4v54EWbdodJz0or2pzhLDzKMPbRG0Tki
YRbSsihukAEyLWFYkFDR5/xqp3iWs2EIjNif8XG4aH+1OHG77yVMnaVX7v87VZkz
j9aZ+WHFFXVhiJY8GLRyo2aWZF41fwjQmutXyDImMaebMHN/asd9tJZidFzGwuZj
2NP7fMc3OHZQfOx4W3fz/vcWJQJlpI4iIXWSoDJ1Vfm6CkijxU60hTb5SRwnnXjD
CQ9k7SnpMi7hoqDpfZODLQp71blcv64bhtllE8/Jcg/8zC7o/vU1pjkhnJT5OrOn
mo91xSzCGN2IymWQdKxrq8XXwAzNM7oiSlIQOCG+YriUcJdIaPuMqaSWPmSld43u
Dv7qcWb01qyq02kBCHa7GIJhPxXWrYSHBb9UQFUVNnLxMbm3bfaYEiwppsqHoYg4
j8S6xyNhml9Vdxm1Var+ZnVJsYuy35k94lbTI56CTfQuTOO2hXou+cGNjEL72205
net0ZM3NFFcYSH5Qqygw0g6sr8BdQu+dp0nW4znQ945Xc7A59UjIw83/cFqYbXeb
hYNbgiMwLZrqfciAoFEHsmW7EZEbua2qbg2IVstMQDW5vBGmfA2v/3WUoKvr35oH
HK0liGArRK3DlFXgIvrwlB+MJmm9sS8/fItNoD65c3zShettgkUNWDEVZaTkHQQY
fMzLoIz7eJjsozUeVfk4i7TF5Xtt6RTimxFBvRnGxrYWl3FzFGt9QyMxW5Q2sf5/
fP2xnaK6nvvp9umXeuC8gXEki2GUKieAMSZuyEd6Cxiz+GfkWsGmot7IMwZgOdmn
xH8rC2z16uWGbogwrNI5BoZYeBbraLEFGfQ/eWhFNrkOGoLlJyezr2E8tvW19cBU
HGHFOtqH0Te4ou1w8ByqJx0RnqIov2TjFiNDwxBrrqr/ucvQK2Bf/f2NzjxG3YHc
mlpBoRCuxAKwdAqNcl3Xv7W58dj1CnpQ0Gj29bHFrCUCvMexGJpGnybq4929xQR4
PXo39Bd6E9lulO+WeZh+nJTGBcoJ8+ulyCANnsc0qEQqWbjL4oyLyQOTwakK+7zz
J9Y5WxpDairTFtvrWhg3VAvxzbDCPY0UM3pgq0nZVEIEvXX2/87Not1d5y80XvXB
G0swyblyCSgfQFbBmomFsgBsnYOR8zAF55UgBsLM4YptHR2+EHBm0hs8HLLEqBqn
HERqpQErAyTTcjYxKmoLHMTEYTdKzATAu5Bo11Z/zlE9tRrdq59brAKbjPjRmC0O
zs9HI/XvQjI8//V8eWw6jy8/lrzwbbYwmMd0oyOgFy5PDpRvEkqqsfURQ5ZC6QQ9
SJCbTtC3TYq6MmwWEdt1MvF43v64iiWIlHDHWvKEIwK3sjG2FeF9tIvMvGSC2MKC
sT+7LQjFC2giqHpqCfEgPQUtZCFvHXB74X7eK2wuNjAxtkgdFMAmncqlBhe+00Hg
a1InMhXjtvdnsrTOK4lhO+olXMxyBrNTTrcnRa5X5qe/KVKEJuKhTFMPGzQKXcTa
ZMPMXCd6QX2RhRRaEFMp6Gy8vFTGULllDB3cuORKdkAqD18aP6wQPmyAoC5QoyOK
d0Fx2NZwjoUJh3aTMnhQWjVpWSdKdzkYIMB7TndQc4WHbJNyYuoI4LZpMZalanWh
+aiYBE9XiXfcEwcwPiEIS2/2IHIIi+MFX3r4IWnvlbIdjomTfxM8vEjoKedx1+vT
3Pk7/ErUVw+uc2CQF70uFV0KtNOtC/uSZalvdLFi0yM+etEn9P7REYg+xU095how
7P7Yli0nJRLhwN1D3Vsn8Gaxq2QolHF5EaNavS1A2+qH/yJzHdigz49DIto7s8t3
Mzhu2eiImO9uj80cwaUuWZ8cny/5R+pGlUtvvHNxrh6nBsWqNtCqYYmjlQj05w6i
xpiGXAa0uMYqGJgw4dhBWeQb0RdyOJ0Qwx9MuxY8nNcz0kaPUP0wPhZce1Yzi3PI
He4q0TWw5kZokbJZO2uNTAr7nYAKGTFLBU4pN1qwPWNYdgygWATuBqYyZRDR2ZHx
ZSt9oqda6TIbe8a4OyDe73FLEsrCJUhb+mhyHWwqW0IH/atNoV65FpS2+T8jNp0d
/UkOtsP9CB2sRjUUifoLPVyaHzYkhqce6o3pckQMK8/9fKttmW0T/UQo0usDQ9Mz
1l6yw4L7MDVt3dBlgb7aO/DKHWIx6TRSBMnke10F16Mjq0GPnRPZ5wRACGwJ0DPL
Rw+aSQgypeqnSjHQ0KycBOBJ9bgmsynoln2thHMOqwTXoqHBwSKmnImKlcXV1A7F
F6L7ypCTcv26Br1gbW/g1lfLzycp0I2ReJSBdxzeCOvD3dw47yvmiosSZg2Q+WVY
tFPSQoZu9rwF/Zwk9Kk7Dpygji0h5Y5nPIJJQYNpA5w6bA3B7ASteV79Ai7nrUiN
cAT/XuiUnbiYWsBWX4NUe1nDT9dGUf7R9H9LVobtG4HVaU1bxQVufVVJQgVrz4fa
plMVxP/VbxUEVaFlN7nHXgumbvOVbsMPV8Kn5YcJFOgsiemC7OgX9gthmCKxyv5V
nJnEgnezk4a8d+t8lKOxWqGFAWycArqb8B4ggW4Gvps8X9ceLpXskmUQs/kSRBsy
CQLND8V3iy/LSVR8621MtRdPXRM7rvhwf/E4raiTfuZ3GxngLtzzP5PWaleLCGyL
XJD7Uk1aZoI9Vh5akK1BU7vFRzOVecfv6nTBYrO0kK23plxur8RhZ3K3POBhOIUy
acZ/zzozCfPUQyDqF0s1dDlF2/6SZelSuo4sQ6h/w6WdHftryUmR+iQl76hyEr5Z
9MthAxbbUH/fTqpiPiWxDr8g6d5a5d567aLu1QNHgyRr74CLVKNm9NP1S/IzaJB4
Ac5MDWGgqTnFv9Sjmrpnz5Ccg1EUU9VK26NY7kRww8dkWUvZSuK5iZb3z5jd4s7+
oyRQGgypzJaZJWuht6UUA9amioyw53NfHmRPaP+NK7pQZDIUxR6zK0UOwpUDHb3a
Yan3WOV7xJINXsgiWJ29LTs6xZ8zRvgyPPGDbZI1tHHAZ3tTarsDeMTu5oiIDn+J
bjwVuxdw/F0UHnlng13YOQgtkx0lA2JrKEusWqS0b7mJxA0kLGlEnqGiYs5CGm7n
hESFLlKBqwo9dHda5qEALuJo7xMblEshjkFRju2snHoO1i/hJk++Vu3y4AA9Bsc7
z4Pud4ygRn6bmXSojw+L9d38WACuZy0KLbmaS3yQXDFW3nTvVidBX0CfUsPaEqs6
VHbAmzjqI7zrZOQT72s62DvxCFnvrMZAifAubM5xyj5l806DHOIcnIXo3QG4I/s3
Os9YxnNqzjWbHBhCkjF83NhZQQMsQ0crjlsauwyuaQsmpTyEN4LNXzs99c6B1LPh
Jvn+v15qiVf615XxlwAdbvJHXybUQCZGCZ5qu7y96D/2aecZun+z1C8dcVHACfuk
cnbjt/GqcJ6pImgrchD9nT1V7BLec8boc5e/NcGTNNxXkCEu8AVu8EDAyLjKnav+
FiJma9GsjPT6WXljXYsFfM6TWIc8WYic6NRNfcic4ambAVfboiYAfOm3WKvW7mf9
vqTWuO1g3Iu5ZXBm6xQ2pDx7jeDdNQd08TLFgDn7JzoUMVnGKoNyyGV6UpW6yH/j
aL93NSePL6pTp9O0Z87N3IAh+cSqpG3K+S6NBGngj44R/49y2yDRvEuVTSgpFTl6
CCrCm6p0ZBa+rnDdZKpGEWCC619y5H6KxNyFDVAQnmrf8Q0lGmVnfRYAViTzybYI
9lRgCAPb56JO1gwepq2l3R88t1NQdkw2Uax7n3kap+FG3qH18scmE7voLheTPTwF
b5mesDiyYrOJQv3NByDAEwcCwBhlVmhQiLktMO932Z+5pTBV7riyQXqMPSrZyV5v
uu8o2K4Yu2coooJRH4BA1U70WHpcX+9xMU8ZzbsekwfIVgTZ/g+AQB6+qFytvr4K
0cMLkZNVqhyj38h7F8lAKk3zy8LGb4+l3nmfyJ5BG8nX28MUk8bWGfujKSbFrNHD
KxsgeHIel5iGUe2s67ix4jn+SMe/kJD2tEjGgRsCve1R2HrTGDRDAtfvPrDI5g0V
98W9NMucr862W+LboPmItMlNFjbC4Oz9JxpOM1LwrlYS6o88pTE56QPa5ad6mWT6
E+ueCyoWLW48rY+xkIloR/fOTdQ0SXWyPFmIbmXYqgngRGg31eiYeK7Ocjq1zjMo
6mu+ZYICL+DExxhfA3AOlrjT6daGK5+6O0kfDeEKMJjW7jP+k6fxHwy1ZbX6n6Xj
8rj5tvwgGQXMo8kEoxktmbPSXoh+ke3qA98qsu8rvVwi6X2AhUzrygFn5fjM7aTs
7EgWERHBeYhAUQDHqSm0SCCVd24hqB0bw0UMjBmMGca4w8gFVz2oiM0qieSuT5Z5
yoJS9hoq55Aihwgr66ZthC9N8hPceB7zmzu//m9Jle1guXGA4JNuMWyRtZ+se+N9
8P9mJqJE6R8PjUNMwBFWt2KJvbgYOUd7I6qyd2PK1IiAvYin6rDmfuzHd0lxQ19X
snkVjAOLoBZP3hlklwwyftouz2SK+QpChCBK6pTycOoCqxXJINjMbQk8gtKozMNQ
0dKEUPi/lDH9i4crHijQ49eMP6C8iXCAvRkl4eAyHtHkt1EHLIW3Q+NWK3HHFYut
C2UAUGtQqyuAK4509rCLzaehlbKBk53QGUHAthamfeq6Z3bsZ6AzcG9uGjJgm8pV
2aLUpjeaSEhNxJL3i1vZYCKFRZCDfNNPaMYsaBe0cKZQoxJpcbxZNKC6u5n9oYQX
8gQX9yYZBq+v85VjFUyxxirS+C3ecEY3QBVMuFBB7ziJ4IAPWk75Mdilr0aGQFBs
mcqMVgdk5K6OFnVknjJJRBjFLCvhHnYY0cTpEu83dEko/3+L1CWwOyJWUHvxGkKw
4s5mkEKUMkri5so+XbhrZka4FKlxhKmKudzpK41JKqmlKz7X5lkukaBLpXCbNQXV
xeM9QgjyP1hLwZMe0A8yFNyEOBwj67EIV9oCkLDDqKqAh4+gp9vDqDBe6P/JVy4V
jcY4RQTbBc5/igDt9Gqn02yPpUWArNnfxZSEayu9tQNthxJRKZFsYV52QsmlLDcc
cGvK4+3iiy/DpwC7OaKNdDD5M97XKsS+2iZOJgo8RcMd7jeBftbc0H0CmZ73P7KS
OQTfw13Sn+1oLkd8xlEhnhd146GWhxW1/LjH24toMPsNkVaUK/X/GCD3x+i1vaF0
5FHGJzvqyefAVnQuCQiPQU0EeOtS+bclh4iGIRMtW813F9DvBUlc/zK0cv/ov6Me
zNmIOxsOZMnVIg0naIbGpusGSHpsYgwNWKm4lOBiAIn2DeJy6OpNnJtI+zCcLS9r
qg0YFrF7aa0CgW/bTaOpYa8M3mSr8xjL2AdhsQ4pKQENQ62mLatgKqYM4cRdPs77
xj8RNYvvLgL4HWy48wd1AbpX4phMLozHygswojJqWX3XxSELb7zWLs67I53i34CU
FqBtQmam9lW+6mABaMScB+gR4o/wi0SSCQflqQJR5YMNhhhJlGyhL4nt+3z0LAQ0
E0uboLU8xolduQu4cSB8GfniEDjMF5DJrZbVRgBgKPS4PPqCoJGTyuYBWFk9bG9A
7Us6Kpl+gQXEW0ioCMoCqobCAJxt2uz1LSZpL/O0x+WR5fydI+iALcLnxrdv27KX
QK1jvqi+6cH3MlOaZxOD0e/kR9eWzjnzz2VyrQsYhpbBx8qIrtsanqPdq8Fupvy6
sqO6GjEaMaTm3YPUhTAbBmjK2Tp4PsHHd6aOyoiMvqanPNqVA+gbGhynF4eVI2x1
Mndv8DGkj+gGSI/3Sah/aEr5eBNFYp0yaoy99OGQrkYjzo86C1RwDjwXWblf/48X
pP+DRfbxuZqFbRU7fD6071qNJZUoJLVEqa3z/3k+JgsKjLvSNA4Yc21QDbsP9nna
Xlj82nR4wd5Y9O9tbI1SoI7jPO5lwUZTYi1/KJe88RUL4MdFDitcad74KZgDuZQs
qW+NiWXk3RqQps98awnd6ORg9CC2hARPs38UlT90KitQZTHN3RhPtHhq+hAaivnk
YmQApG3gwtWgx60BnUBfLLsXnGaq+xEw86ZdLmAq0hxuJLc+s4MRUpCLsMULnOCK
zBcNUfYnlY78W/PImlegakQ6uVHrf70eizrLcxzyAEpDIKlTnEsx5a7DNOuUJKUh
6hOcEtrypvizRAVA/i6ISa3YNfLBqqxz0MlqPLeyE6bcqFIh8nbMKnEV4H9qyuoZ
YnUeM1MCgGtpNnqA5Hf0CKpd3BF4RJXDBLFLgtjHuX4N0upY9Fbd69TmOQcujptm
Ot0zeOlOD4ddM0G8NcWNiKiiR0s2qntLZ61Lh94/4GwD/pF280X1IeRpBQFJqZc2
YXIGIy6UCbjL3slX7nkJwp4jWNlLf4jBGm9bJRAmN4MSO7lM4dkhDSy4Z4nBw3K9
8zfTGAHnBdMgVqcr0FQvVimvEG0wNquOYkjvliH10ZNFPGEczJ4sRlSfEhOYSD8V
BoT3DJCupal2BfcBwGHFHz/iXLUC7CfJXcV0rtoAqVe+9UxJSXi5NlxrnvRIAkGf
Ez+6+DkmwGTopc2ZVFIb+aXlvkE3kV02b/jVAtqPF6gNdovZmILeve23RFTg4U36
KyWEWDeYrl+WhtitkJVjt7lvAUPdkaz+MX73vr8yJ6DcQptcIpIu5Neb+RdL0bxP
srMstrfIvZTlB8wQcIqRBFC2H2yvqXoFffuGYGfuvG9H1eeZR2MVpD8a8DVwxGCl
3xsbf5GoZxIhzOZIExd8jHIGvOLZSUiC6nqp4zw+ncBWkJ86736ljjrGlCVL/Wbz
I3rWV+2CZL5Soveea8x7pwMuer7SMxlLcrdKM5OwRRRVyzBBK6n2tI+aVcHnxtsi
6w96OjC455ar1rJ4S74sH99HFNUfcDXXWg8pKRjn1OaJ9UZcK/3LN/JnhdzoChsh
h1ysYJi8tylMAsgV65qgFnKKHAWxBncl2QOxAbUS0yEZ8+BRWNdbYS4Tdg729iPo
39dtV/+1BtxPFkJcdVLQzsuevUpAnbX51fhPx0f65JBleCYdwoLsHrST3/QXQE1S
aHpqc6HWGppAbfrEzwqJMP5dOjb2H1Qk37fCWaO3kpMAtChkGYAfddrRnvfX4kmS
EZlmE+qP3hcaE+hcxSgzA3Yc8rWVKXric8xBNJbxgNbCfcYWwLDx/o80y55l4CPq
am3KqdTvcl5hO3hWsEQLCKzuAaduEfbk7XT4BH0eG+WpR2yHgjTDB3LNEJ3WJa6a
p0bKM6o49cYbfa80d/jYcu1/07vg940+U3sjQBIEG70v4HEI7caKVMS77AVTwc7r
WsePJPnANQ1a0ktSma8utoTkrz81d+cWIOKgT5PTqDXoHoBjXYZDCbbDX4FT/aQ8
zQFzuDS7Fq/cQvxQJpMeh60+6Dhmq0qwd1rVmesR1NRTVMPFjjlSftXEljEg5g/V
HBodMTA+3ckJk2GwFxi/nsxgd7jEZ/Lofq5YW2nQJCzucovi4QuijV2IiZlIsPqW
0i0Jui0m7FdfJR4OglIaOC1lwMAtOAtzReQu3/+R6QEMTKaWah9G63cCZfDYzxFw
hLpC2UCfsnyhJLfCuQrRjmjlfFUGibuNDtyyTJM/yxCbkNEPypB2NpfjTXknrpGy
c0B6Ex4BUPiJBGBVuXG/f94gdWBVYZfswb//blPxN/iqiUYxdUODonwzeZMlxck8
4Rje056bF51+XgvZPEe1vNHDxQXjAK4QcOCjklAll7H0xc+y+6syMWHZ370GiyMi
yurpiRkg2upXHtQOtMPY8OHSE850ddPkwPImCoFsVIxmGeVj/dPLOJI5V5P5QWLX
`protect END_PROTECTED
