library verilog;
use verilog.vl_types.all;
entity IBUFG_LVDCI_33 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUFG_LVDCI_33;
