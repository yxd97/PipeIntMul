`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QkbkT5kLobTajjjjdlI0eCsaScF78SH0jnBnEMneMX9bRIXhz4yglDPIMQKW/r51
v9lEL3R7AbNz7ivdN5C6EyGveuia2cOs2PqmIBBS64/kl4z+G7ibx9A7NTrZ/EFE
MLpAIJF9YcQZVJZ94HWMvuFdbJgRGP893puIBqmUCtOU3ioGfPRz5MNgKgsGhJJt
5YBRWLV9ohYa/jdK2Q1uq94grn26/Sus3eYmnKbXz03bH2Nj2WZ4zVOTuE/YzKa/
qr/J90ASoxTKxoeb2yN7leuPddxsStY+IxWI2eAQuri7n72NrG5T2UDBUGplvDpN
Hx6nI9U3hTk5fJkZTWvYeLEXS/4QRHOh/np6o66poKyn7SG5uMAjjKxm3UkV4yof
DHSj+eo89A0iCuxxvasTW5yi9CKmtqoQ11eA3lCCo30s/zeuw53xNlzjsjhbqYpr
QY+3eqorY2Q8hc8RsPrYs+XtwO5H+vAiM5fe3bBgr/ITjlr5M98nmZci9T/7/2dJ
ph+NFONBtI2iwmtgqt/OLdDq/xeJI/Qu310FM++bdzPx89OiWVREXrNbrtm8TgPd
`protect END_PROTECTED
