`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cAAni+ZrLb9CS5CviKkR0F+7dyc8LOczgew+aU/EXzceMLAK7OplkgzZsdRX7w4r
5WuzhjfD/hvXn2dkMrm+dYRq1qZTcFIrWTljSAjdnYTNl5Z0E4afheClUU4D4RIM
EyePCr5oCA3Q19qu/GE6n0bMas9uaVnZlzGdW2A8VAcMKy1DyIjY1PcqRBQWIYOV
J2T1w0C3CWc9zWQvp0dN/M381q/xv+oVW8e6rFcS2VNIQW+3OkiZ7ueD+4pTJJtc
inN0LKa44z5/OJnnG6d+OKJ+AbABOeeiw8By/pcrAt327ki94d69QBrfELvKh4FA
t1aQPmPD5dTObXOooaqZxeOaxwIFFRZ4UIgSLLVknTiGGcrHgchCb25ZfFLR1Fkc
5vUG/l/rQCdLTO0TU8ARbg==
`protect END_PROTECTED
