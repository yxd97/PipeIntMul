`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gaJK0IF/fbjWClhwhx12uIJjoNhKkv+AYVLI9dYOWF+HYmKy88LrKOBxqN0j7Fo4
XxUxs9kT9zp6t7YE0G2aHXEyff6jOo60fE2eTYU7jvLd++SuX/s0kRbK8ktAFPYj
chyd4ktYNnBZf41Dv8UeTgWnKhI4x6M8Hv/+B8gvKQRsKqMaUxP6bBCsqDhc2n29
IK4CwNmzUzgHZVw8dMhm67VseSqsAQQBRHSS03R8k6dpOl27Pey/DGFwwNQgYizy
jViJrs6mkieFy93+/wHQ6WHjhXgFxbeSgDKVttsjy8Kce7OAG3NoYtRrwCj1EOCg
/Ns8U0YLCXgsOS4viMlkRHOFr61yJJHzOsbtuMPHzDBRncij3Hb5be5ZCQtw1Vob
w7sfUgQCLEUbXTN8UJxikWADOdfbzNIdaPGC4MeyH9w=
`protect END_PROTECTED
