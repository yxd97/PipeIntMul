`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GdrITKPD2cplEcM/P3Irw9bEQiBLYwqOcyVR+1yQrj48TJGoBWVFcxyVCceRjKby
remDbXfDEHvLSpEs3oJWXgX5RxDJE7onwYtR74HHvBewTEAf+1msuK6G5y0aepWy
4Z2jn9xB+C8SgcFaiLwsbg2mM0JsNKIpd6g2Q58OGP/Z+D7eXrHNdqlSzt/Oyccl
lyQ1EUAciSCQ99vxICEMLIaHaOhSYhGSphQ+W/f5LokzzBcOFo3aqv5eqc2pgjUE
M6YfcG6Hg4t4uOt8kTCuIB/blPCmSlVmU/8HcttfPtaFbD3+HtXlZtvo6ktnofDA
iAwpa14mhYSRsPRWdt4VYatvvtf0/9IOtX3ACk1tP0eLVspi9ik0w6IqglihP8vI
l4oX9JUVTcQxlIIYvw96yUdoSWvS5LX5mXEWf6/jJQqWSu+2WOIoDUjPEptE0IMB
M+98yZBl/GoqU4u0VxokVDb0EFDbOHOZ7DU+JJ8vZqRxOBsSn8UVRnNPvKgfMN2s
Hr0l8Ph1zeGPfuQKPgSZmKSPg1/HBA50Z7ti+nrYXRwbng3D/tO7kebPi6gXYhTt
PQeWQyKMleb82I1+L/jTqvO19SthragqpAjGLfoqPYcVgkP06EkIsfQjLgSXqOgS
vv9WV3Kd20wgpSPZR1bVU1jh7CSWCTYHsplpPwuh4RDQS6j0hNC6NclmqhBv4jvD
aWNd9VRvOCpKNP1WNyp+pnDeABEJYs2MBs0G6XBd13ElLtobl3yTNUkU8GGxCMKA
T/qRhunD4cdJGJJH65OXeWJkylFtcGViFvUsEa+QXZTPQO8fqXONcd5UwUDnMG3V
Ru3xI99IWmfy38s7PvN9ZVP1JE5IZpbciUVOPP9UKLgFGzGIAPiEYE2zNMFr9fUV
4d/5s2ExGfgp8Oow8ipzq5USjrDKdZxUPYogCWeq1g/z7ake3jZaKbF1rUHn/4Hh
ghbBuLHjvpyzg/UiM20WKU+ir9nslMn10GaEV0jwwhzjbmkb4mCfNyGL8xo9K8dX
JsbZtNca+Ok5Q3t9rEiinV8h79JRNL6/4IohSYDJjFEu6WUEGRsK+BTg5geG8SQH
mnFbl09TfrfDSbi7630bUIOmKgRV0+zg8pntCMOSOyNkxZDl8jvstTEsZ5M5auPx
JlKzOkgvRJS+t5IkLm5d048+qVs/eJ42vM32c7sTd8z18u2lpSPDK811Q6nyIXeB
How1pYzoqs9khzAxuqnZmr8rzf7h9hWd7cAz00dz9OWdwr2zktUJIbj2n45NWq0g
Gj10wHRNWlU5iDA9QLPpVyChdtmsDrcon3nDoC3tZetlpCtndfRqDkYtIeaDHhjv
qrpljZQu7on8+qW1rXJC0YC+oKF29ZYTIz4Fh89YAX514N7Sji+TkVr2H92G6q3L
wD0duur4ii6adcSIDhNL4OXZyDPet+Z/0cEk9B1A841a887bRA7peY5gnqGjra9d
LBMNp2ErXsGkDv8BFXfFuSUWcd7IlSxiuknKMQKdYKLUjz2BDgEzAnZgFDR5qRcR
NvwH0SQjqa/034A86ic7NOUgngIHqF659hoPqcSHhAslQa8xTLIYZoOJ7+pkC1ga
PorazB8rmVaCAplUQxt7P2hLO/lre31U9kaW0EASeoWMiYVeAQNinMx8NhQD7qXr
IOv3eUrpqCAWW6bwbBqq/QM/DnS/j1M1+/DdvDdaJfNleChiRFo1iyjDpHcpmCjX
wu+55n9h0VjfVoL63W499VaBX3XcJplgctHmoe1B13KYzfzSpq7NWpc8Gz0StY94
uSoX8m1lJSGGglfJXEo5OwTB9ina5LpUxv2l817NPUZjj+PL08ovuGH5O1wrXo9/
yFajKsQZ5/bNgljDBJzycfcBogeq7AxM4Uq1yJl+RjY2NazMVPDb4ZexWyZPMgsi
DTe0/b6p9/kROsndJSjPwNl21Ob5StQRqgC45LKQZnAfTU2F2ErbSQzMrsdmujHr
7JeRyIhbMRCkJjWIFGxXtvL9aCrFBdNiSB687VA/2zda97axbPL1+qnfP8MrZtSw
Ed1KBYGSGkklW4NMySGy8Qy0vOpLCCOXGHUikKad/JAXpsW2kuGmOo4HjSC5td5c
PwOUCiP8Hyh8ADGFfaXEB0EaB0Yxln86LSDR4gbpve+zE49hXHtnqk/UuMbOEmxx
mnECMmnurrTkCx8S2G0E3K3a6hf677pfQOy7/n82MlFqv1iPEC0zaAmkpJu+eJad
s0s9Klx/M4oAO6CZBwE32HAWsuSybIjsz+iEOsitY7NykrG5oOET/mNUp4+jlp/p
KieIk4Wmw1rTjNGaAT+Q+wMHk/s+LFnRtcIPY+YBfSE852JK57Z6U1M6Rrg5MYRp
yRpuCRjr9reTCm8XFwoACZoGooJgI4KlHS0wEdlD+ErXw/n1Xy4/PwogFOSgEQCz
CrT1doZyDzLzD4vm0AbiJxQ581pk/dvosQT1qFP1Mm4UuTt0im9aBz/2d9AVIZhs
4QgHXhsNoCHoNdU25cWmhoor8suyi8Ug1Fywm62rOb2TkPW+///KQzdgssDoToSG
EVernlmEerqMnFT5DyWjHDK71YS7BEbIYcE7wDVaHlVdb8pvU7Q1U46CMr7RkNB1
Hfu5xPfjHSyItPtoXv2wOeU3yrubfNqCSbvGzqHrf8aWCogsHcu12Y3VdJU2UN/A
eJ4DgRu79rDXZfwPbKzoHfjrKX1RBnJ6j2XjbvhwppCgEuuHGmt4DMjTxpOcwjGB
0F2kKODpCsJfvkXkBmdKTlwKV9F9Qxn9YZXJU9UC55beoQSseDXXNhvc+FQt2NCs
PFu0V3TyFntuYff9pA/G9e6qBj/yeYNIbS+7lu0jWe2ANeHknFk/3rlWMQ+1+6PQ
EO2GuschUEan6FcsgxKSARbewZ5YMI43hAL7bN8wI+BQGd/viiGp9LNKwFHApXZT
5P34C0vuKXV447aWuy7Es95jGFTdcR42vqHEnP34Nbxo0z9zAJTOVGJbmstmN/o7
clOZnrDsxWk46hefX/hcG2DIXcQwmAlovxP//fyGc4TbF4Llh53PMGVNYW0Jhocn
G3mioxSeCPwRwVAMrQS1nz08tkDCeIBkeyR/U/BHNW2NWx/BeAuSZilwFZ4vgRKw
n1n7Cb5g7Dt1Ok7VD3Nhuni434o1FlE65sqWWMKhs5MSb4tDHRW53isQkcbfnzxe
Iw5foBA73ggU/hCFRLaff+Zm8scwH4Ow4zbb52+YXLijmYFWwTVNxRi4cpDWC8+q
ihv2RQIF7GO+WT40SakWzLYNIVd/1IDP9gDQNUNWmyO6nbcpYT1LfEua6lZAvPbl
vq8wn7IlK0/znG04YU9jidFyIk854UgUyrKOqZS9u2vt2kdKOeCRn0aMiVpjrcXj
pOOa2agLyiD9DsDq2wDX2ziXSzCmKM6LmAdTV2cQ6blK5B+omv1IqqszxPT7jnPC
3CX5iNMc6ojU3ZMkI9qCBpT1Ms4r6/O3tvoNYs6jP1W81iKRU2JyJV5VEyqT2bsm
qjTJjA6yzx80PMEHeESmX3w+A+8OYGin7XKLTkZRfGSJy1oe3jaDBsCBkmGkWGFr
lOpIYNSnFZkqrzMsUrrfNfOvQfe03BIdMQyMt0FTmPTL9bAxD5rWn/N2iQkcBnkq
xi30P8h3yyPcQjEO2MGo+PyqxHThcClgVybAFdMwRsDy73I8SwuQe2avt/ficZAT
/2a6z7GCzbxFagdoVRq0kTIUzllNBRyseC5ve/9UPrm+PxD6srT7LnT7VqiYHzqa
hzMBKE5Kjm+B+rYDqr3L/ITaECDnc4yG/EELLf0Q76FjmiCtvg3EtVEBONaRtHSj
aStTLkyoO9dwv3m87fbzRMWaN2H6q1Yi/CpoX62L6/3dOev4ZIQO5WfYbQZHvEXD
U08I9wnWk/dG9QtjILV5pS0eBE4YmBfVVnaK8bPR6Dj67LzDyWs+KjkegzPxr4Y6
6yKxRQ8FeORibCANsUJjeuAbVQfj9k+p3uGMDRtEx29zCErVVfwE6HnLpxwF+ZZi
9c6KrwFSHOuUaXeG6OWi2JBfgV2A57QdTnTJJEYxwL3OWwpDuyhW8jfNlTwoAS7L
`protect END_PROTECTED
