`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OY/6Rd5qJc8CVJoB5MxDqEPH4ewbB/X0SOgUlquKPolC45NeNucPctFTt81FvnAE
RlXj0HI9s2vPsu0zFM8VZkoBkA+3uaoY791FK9HXqNz9gRB+5FfI2yz/NwE1EPci
n5PJTe8FhXO09Oib5QHF9sLjsxg2QWcOLraSuRHxh1d4nN87pFJas7d1APGG0jCY
z0Ckng8750qr4Kgwl4vczWfTQyNfZgd6fi4jHLbDa2/e7kdKyUDFW1YQCpTc5nvK
Z1NAC0qqGD6QroAoshi0beinqLsysQfBD3U4zWuuWdAov2YJNN385pAgzT0V0uCO
pVOP+gzopZ/5QdlU4rBF3XsVoFeMELypkzzYSO5cAaOmJPH84IOZT0XXu/po3mfj
5TIDyUsoFG8+c9H5s8g6MehHzQOgCTg/30Fan0aOPl1zVyULF0hyFPoKXWxTyun7
i1TwezKZDFApZImfXIJ8H46jUCW6jTPuYKUZsBpl1C4=
`protect END_PROTECTED
