`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4hEUHm0/K6VipWkuOv9LLUNQjgpFfvlZp/UjJk143xWsF4BFn94ExX+YKlDFMYFL
EaNVkNTIMqvShx4L0XhCg2Wy0awH5obVfANPhtnUNgNeuRzIycA8bt2klJ+0Ca5k
jAtO0Lvg6jF31jd1b+uGDW4pYbHKdu/35/izisfrQ4bx7wLQHeyPDR07wAemHu4z
spUGmjuMI4bgeOY0EwHWHiayYo0iLj0O/iLbQoTXJP4t8OM3X/n8gPy+c5avblDe
kYAd+0lwN5q2dGXBLy+9ssOGlWYLZr374njMPls3in/zPlMvngNh0P/w22BXp1Wl
Ag3WMU81Bcb+Hyk9LaGbckEn4kVUiHxgCGyMjTraj7thjkNOAwJmmuXLnLRZ/Lc0
i97wwb98iGVGUPqvNr1TGfF0BcoSXKB8ER/8u8MKhkhLhAfU1CjQuua5pwHUL0C0
EIr5NXMbNZ4f2QtGc9vtWL6HcZ995yJ2akbwBlhIymvtmcdWe7PXkAHRwoPPIbeX
r7yMc16+PnFvAklN8ezq6ygJigkygDwilo0NEmvP8WuU/H89A8fz/YQTp9TwSwzx
0CqnJHnTTbdfP5zylS+AFfxaT9H8jE6iAG23JwuXLYpWmrcu1+Co08ZyE0bkn/2P
JVq5rLLjYDD+S2q/F8xyUHpHf1UC4uVnsxm/pJKdY3tr/C1FSwZl/Bco0ZJ1X3T3
iW12+PvGqXnwHHYiR0mgme9SFdAly9FB1ni8P+LiBwntzWwP7s8JjGNXFdAOVc1G
1dOV/HVMpszfOCr/fdyM+MfCNmhp1BCzJITauVs3xEWybZXHSQR0qGxUuDY8baWO
JavxXtWsnOe3tIVwW6QAzL1YI7R3b8IwWabXO2bkiWQX4Xeh5PAgr7IShJKIzk3d
1pr3Px1W6OCsNCatggxISk+iF3GZqfDnb9F7iysFhyBrcwJvRDaaNaDcy9gtQ483
hfPAU5nEBV3ijz5r7MN2p+x2epTsbNkQhddO4vmDdkLZYas0gAA0glpT/+D8naGB
ERFzj2XrqBUtdDMd1NNg1nb1FxiFyx92wx4jzfDyXoE=
`protect END_PROTECTED
