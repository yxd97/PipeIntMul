`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAEdrEAPmo4yPUxg7va/WFEGCu0U9NrExxyTY+z1GHRLIzdr6eyv/2lVXYH/mFWf
Ox4rhHwkMDheSye6d25E0+cxTgKX80louD7M50F7Mvj3xLqRyhkPDubQcUPP/8UP
13qajdFvFhZHkxosCrW9bUbAyIJyNKwed8olFjYW+xyD/xA8i8K7iv3LhfEUTUFa
Ve+kyVhQbELjjmDY/QFl7OQaNUqc6fRW9mbiwCZB0JGX3EyPmmBD/z81BAJFcDOF
6nSc1c1HIs6pRazAm1eZfPICvE1d0jxD94G0qr6kBkiF8ZWPPwuue8XDtcZ/btyi
idKK4Ob3YUxQ4Eq86EIdZLNMPEGlQ2CfiFaMU5KEieOYOiilIEM8+yfNEW1TWtnZ
SbP5/h6CtEz3mxomXVmW+qC4t78lu3QX0KriPo5JWKo=
`protect END_PROTECTED
