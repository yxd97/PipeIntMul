`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxyAw7uYHklbUSJeByGNiDd+OzKFTdw8JavzqkrHWpx2tdlp2XmAQFHPJvPgcq3a
glDwacobhbqPTG9vR8R3y5HX7JEhDDyq12DThQd5hpbxZVzkbd557u83lYLhZLoG
DTWEzTYMRII3ooZIkctUcIcK7psOt54xcf4bpj31CGMeEaHUrZiar9ck4GRocgm7
m9T2DyyU5+gpTRRUXwBJAbSviw2Tdxc10tcJCQutlCfnA2jnsnsQIEBLrlOmoohN
i6erev45sTIbTFadNbMbuPn6gnzZ23J3iTKGAzQwVN3Io+EK0dmJaQgYHmcl9K/i
qfc43kzrLnEwm/JEkQHWE03YPE4AvrHEpVJspQcjQlmdjpFuwN/0Z1+Uqe+HuGod
gjMTUeptMI4QTURZ3RVJv2A4JXdJyub+2VMLQL2cNHEKS1d+SJiQHWkUHZyyZm6m
wFrixsLFLasWI7RcKFBsf0pV+we0dAFhGhdLIl3y4sTvF2ZKUACExxe6XF73WZpG
X4XbiGRNXlDEop3vyc36mraNq7RpvAo4SD0Mh1tLjg22z0wpIgxfgRskgOyjxTqg
2GxzPjsyVSPuife+VDs/cjrqE2ALULw5kTvubAb9caEJWsAyhEUxJvw8TBTN3Jjo
4+6kYTGY6IZ926oDlS/ns9y1TzlCYLZnQgtKRvnbMMlGK9lAyhB5w4ExkN4KDbaT
FJC5cC9tcfVbQlIYMfXh2fO2vRSJeWpDKc68jVFCNVtlZRqBxj2/z0iP7cw+TXjC
MvDtgQ9qE2c8xS3Hex8gZwJ02CwDG4d9ZeCb3T30uRuBlosHBzJkiaJ0yN+w6lHv
p+oh5NbdGKpcE3LOUA9WrkPfSy1Bdhp37bDvn0FH7Dpy67KTAvWFH/iyeTKMckCR
ReNh6LZ7tXMrTxpyhj2P3A==
`protect END_PROTECTED
