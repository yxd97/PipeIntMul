`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWuJsrrksycQQEjr+llUZ11mXh8fcv4v0UnBCRQZR8g6bP7P0ewaehU0wAlkwAqj
zVcTLcFZBO/5/XJA7J2ixHjwevcakAfcd1rdjkSreWc0fPRv0KK5sOJ+0QyeXC8G
EVXLdpp9QYX7RmyxyzB2Qa/qA7KTbud7a3SwVq/zSA+wGN1qVUtcHCfdX9VF2s61
Xku7BBsuM6ngAPRkzRH2jGrS6/kGD0Ll3CY0IU2Kyv0P0IN3K020I9/FgD0vIpwI
KAbmX82vgfln9xA4H8lnbw==
`protect END_PROTECTED
