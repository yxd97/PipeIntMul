`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SWKALlkqNLWT5y9UiZQLAPBq8X37LFMXBcKZZYKH/wI3Z8NQSfUhe2Rsj48htnJD
8cRxVb9i7topmx1dqMZ8hc13CLvjZ0RoXrrsuQGzYIvd3unq7H4nsAU+w7KstnCI
Fzz98W4nOb+n4iT9yb0EVsDpYFJCevaRn/81jrFvH9cYHatZC4wKT18RW3nD+L+z
Y+UJJu5fOoLTrNrBGn2+AMzJk5MytF/6l0ILSAttJJJTJCD5jH6SbLJfRXm1B+0F
CFPWzLgRQWM2ikz+N1iJFd4NH/gcwZd67+6/ZoSecqqFdzThFWMKO9itk4Tnrlrg
Mm5LxUEXMQNZvN0KcQci4L2DEI5qHHPrsmrTsbqINnEwbePpuuP1J0/+QsFnpbfY
CkIWO9CjzcNsTia8BHnqfqlsCaaDgEVetdwLc+74oveM8ObhVjzKQPedH03+kdV+
i4cG+dMvVIIU+g9FOS9jRXqlik9OGmdvtOi7+t66YJW6HjYZD8IbbqW1d2HtPr1z
ahWZw+afNqseMxVmqF94Huac+8XuUQaEwkjZij6LcPYle1H1zKlUCpwMCi61ujpt
J/ZIyXAFpLJoINkbLnieSwwTXD1NlVKGigEyg716lCc=
`protect END_PROTECTED
