`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A2r5ZW2L9sx+g2fSugunMHrs2LZNTw2sZlZ6AQrksqD6tvIr4n89Bs3IL+CJm6Y+
V4MQJQ+/gg13XpzCzynPuyLhfbj/WQNfqXlpD49gKuTb/Y0go4PeTvzyLSIdWECe
fpcV9BG/fIcddeMJxLbAX//+FLNltj2rScdIwg8/fApdLnAVX0h4H2LhWq/i9fn1
1zwshBLZIKgzeuwY95PST9XHZdrxDCtnsS4FCdor89i1Lhg3tGqZYjlMk1cMkUNu
I2WvaLc29zUDAi1Rf+NoiA==
`protect END_PROTECTED
