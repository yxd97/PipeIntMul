`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tkzBaWM88E6HOQLP1BSgM1EiZs+BrF7Up8/4qDuMKpV4lTFy1oSpgMk7S0MXQl+v
B/AkRWCOl/NlSJ9sEE5AqW3BDiDfTUsTC9UNqzWwRm4RgnQLchooGlTBXG2HgXCw
HjEnnYxTWZiJQTRjHEQIpbKYZRjdiIgfOHxGoIp4Z73OXgqPLIbKXljuc0fI8Xxh
djTk05mIkIX5Bhz3lgla6/jqKKtjCaybaP3Ya/qoTN83K3ff0vLigzz7KyiJDkei
oH308lsoKbOr84kyYrVSeoHD8H03WFkb24vEL7Fq+gz8IkxBYp/HBdbHV2Y9RXAX
kiv182fXa/hwIbeYqosyXnHCm0xZSDimCHSBEazcrhMTv9XmLfxZH/rdfYlVv09o
`protect END_PROTECTED
