`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
02xDrKNUYYHUCgeh87ojkl5yC6U9PBG6RLhUjBqQXDyaUBDRVwfFVtoq040utq2i
5ivt7+qx2rTep8G0k88gpRipIPRlCpax/hkCB3KVfuUffMj+o6MjWG02j6kVnX9/
kGwXAVoFCDCVhlX/QubbMF9Pk7PlZcnNHlyl8BbyW7hjadNhy/jKRCqIHaZugSqb
X2SNjU+7rrgWma1HrDRiB6F4bKsIRBmSX3J2EgPQ/WZAW1TxK3IN39gxWK4Co4vA
/2bsdAGkEluZ/aMAb+xB19cep1tg7pcHn3OLgXA7rXrdcCPcOWVmc8SxtbxaMsru
GlQXA+PIGmkji7d33EaR/Q==
`protect END_PROTECTED
