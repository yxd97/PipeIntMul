`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
goC0nEYBnh75O/Z31ZXDrRH6Vo+REcZR5kFx7XvauXT7IuYq6sF/VUNhGsuul5um
gnB753R6U1HnCncOBpPuGji39dt7TqDOjGiaYq16tDYoJV/h+ch2N7SJPk5wHRfF
ao6oI4KGohnEpPfHFi1NS88n1dBvq1lYEylI5xCvVxMZzaI12JrplzaYiUZyu2Wa
Qeo/NYcGVwIeGjCa69DvpxUBPh5y1AEVGTy5/Tuq5qdYEz1lNMH05+GtWSRE3rPH
7KNUm80mcOKeuCCVPYfIHzcrcrzkYRExZ1HAFg5uHd0GvkD32tCcmfJJUH2zCjDF
zeB6McBYr+sO+p53X0r6p9/FuIV9J8uE2Rf6XUcmxC3hIi3GkzNmQVxKRd6+QHzG
gxjy3emwK0HWduI5gY4we7LJsS8R1a0DS6Rp/ElKS1DiqGiyXUfQPsKxBKS11ALA
pavm3iTHD/4UgafaJdi+MPQ/mtuBUCci/7Fi6qvUIMVEIyZJFeNk0kzhIskxh0+k
gM6IzFDLvin7sac28UXR0yMo40QDkQyznbYgHHETiWgSmLUhVyKX9dmzlBAgtIgw
TaoCpJxv1tA7mV9q9Wpcv1y/sNv93+QWvO6OBwRRtHr3VwO0woQBjogyVKlS08Od
u1Q9hlnreGoN1+nKzP81vXqnmmxDpsCgAr6CBO0TlrIdCuiIIApg0Ah9JRvRQQn2
8q3ll2F9RQJQuEf6Kiis9XUVp1FMMiMa5zApc+A1oeM9vTmWIXkTPgX1pPZLrXtf
xTpfVScYkVbSrGDPCN8oEaztNVG/VD/k0YB8rNZcYhNDkBVYedFWnHXNo8wk7TA3
5Tg9OaMfpu7H9jNNuzCRaOtp8dKfjQGEynLadCcdgUccGqqBeqc4+L07CLE1M8/Q
iH7HPPEJClO7umJr61BLtztFTCVBCWrYJNCLvWTUg7aaFxRc7/cXsu155h0JO8R3
MJ2jxgvLzstlXMwzpn6OHbHgfWCjftm54khEsZ8+GzIL8axvtdaoGHZdAxOCC5q4
rU196qnvE+AnKFT/OX3synDsby8DYtVb75MY37GmhCMagELsi6JN63AaoAunPY7g
v+5QX7EjfLcW8ecpYpez4A==
`protect END_PROTECTED
