`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
13Y/xNtizVIqpbjbZ9Lntpq9uAJ+wwlDBQVRSgy10TY1rvwBakNZRXx/QuOacQx2
i5YPF4bqCgI7kdc1qVsihivvdfywr1UPjeQTe9vHeXZcCuxWzbU/ic/uQqWXzOBD
g8kLnaLkHjHR31WK5gK48K2stiwoYd/WeJDQJklYpfA0cvWFPEBX5Wp3hxtaF4Ey
sM5LSKQpjPVNjYU23aeg7CwG4Imm+3G3N6Y8zKj2z7IMck6kp2dwDqCnWMcaNVY3
OXtgTn2usHaTpQwuCUYM1aP5yBlfQQPoBH6mOvdcqGN9KnQbIAHJK/YudGNVKmGD
ZLEBIZ12NqBUWEVyST2RWXVG0xSTx0j97wiihylhMAcgC2P4kEQsG5OCmkwbs7Ku
TSAhekbcySKVKIkF2Z7EgVmiaZwNPqusLrIh6HUO/msTExTDFJQx4HOj8iqcWa/H
mH80U1UdBLU46+uuQJqNagqZ44YujDapRFX/H7LJb90=
`protect END_PROTECTED
