`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UAC1HYKEDyn+0rmLXok2TRjZ36xVSdClJvwOQiJ3K8Ro4FlKIk4NiLuyv3bi5kpW
tkutxRotL2zrEj1Rkapw3ZXqkZMztpGfsaQpnoYlsKf+HS9vdE6ZyViLJinrbVoj
eIrnKPkpwnJ3Mc7ASAv7TH7SY9ZR2PvQbyA1b7U/cHnfwo6qteDjJOJIZMSW6Wtd
WWmkkF5N40QQolicQttVb6kISaor4wniZqkJRq01B7lIlJJdweXGQiB7NHgQLkp4
SNFmO3OoQyZrCQY61o/Pw7QddLE2ZA9bO4GjtagAcaVh2+wBy8xWzC45u+YyTyor
2PmgZ0SAbQ6vlGp6ReThVds/o2wBKPgELqnl4YxVfdwaYklkzLgBKrjn5fKD2Lw8
7t6EcC57dSGPluvAFnGKAMO9Phv3e+cwPQQ27fbsGwAw/KAIsSW5uOzpATZyF6Xw
V8wtnw3bv4YNZVEJ0viEjDbjSoPIN/SeSYTlQ2es3/w49sp78326oFavwtt6dq2M
+FhdvsC/+b0Qc9Zpscys83hXPZJGhDtq3BTHP7kJ8RO5kxwb7FnRkbsb5kYbmdyZ
IwjwWVB2vJtfO6xwJD63177bONgLUeQiXOg6gcd8CpzWdGEd2E/K0P36mDow+pMC
pkSzVaJkJi1kuIdn/V5P7f7u+n/BXzmi1jO9jzWjB0n9fuhfRGCQ6D4IiaUxZTCf
YgMzQ1oYFvnh4e13IFyqSvN/7Y5F7iKpPTbcOF5btV8e3kh8vNRIDwP/glu883Mw
xtsYrf9UpulrH+0872KLqZVXX1uS1AsScAR9AZ345hEvepUHQcTAbYoVtk1tN5J+
g4h3WXekWVWhnopDUQBdrvpKraSN6Czoqf32b7GPSG31/BRzUDzB2tHp4WadZuvP
RkYxol95Dyo+a11PfebPwgq/4Tq8JpQgxFbzt7pg6GchUC9hXFJXqJTAdUE6HdsD
RDiCcKLG1zmLG9xoATDXFe2mEKgL7qL2fCtSbCo9LuW/Nnx+B1K5+kYeTsB/RCNd
F4y3uB7oOQt58i3+q5+BhQDg/I/TGyDDY/0XvpDAmbUPWKYbkw+BShP4uXOXmk0r
siaC/I7SW3OzCIsjMAExXHEwHFgeX8kADGX+VNgvJ3aiVDv4ihb5v+TMnEkaSigL
X57PSlDAFPALLMDHXCO/CepB0zfiStLrQUiB4M0hG/SAudqd6hAP2d9rcnB/OvFb
gkYTGDH72XlO0txhLvO9Zu+31CzJnMToIHeHTHFMEYc=
`protect END_PROTECTED
