`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHygh7nf/LkMD9owWvjK74jYA/ExfBmxEQTkeDQFOQdog29fzFhqNQHzPvUbA0oX
lES0WnuUiftMVd8ysGwso6i59h7pZdXaI0L71mbiFA9X4OMGS78OOHF2anjOReYD
tPyG3x51cfQKj005uS1Yzeix96tCx7d+/NV3jVc+7URQpGCEdmiyVeoKteiytWAd
VHCpum1iuPlTrBAUEai32qaTL+3V3KHJ9y4Omm6V5iura9dm6QRk5r6GNAoZLYrL
aYvmGM+zahJjcnREZDrI+GfADgm1c2IbtYVJgng9TtcJi49lC08XnIhU5wiVU/p1
mFtBIZ0gHgnttEWFFR1S0kl75WxShXWt4wqsC7Iq4H8NEzYf273KHfrD3szLHbSA
ccAs3afY6lsVgyrpp3aTq2JuVT7atMcj1yKABAOAnzukvpsBB6FYYHQZ9Uq3w9h8
/EB6sOEtCxk0gq1b19nI9xTmFTsQ8/2mIbdF+skHfa38h8F0h0xTCAn+eeYkGds8
OxIWiNDzs6fsHrnQ1yaK3TsKIxb+5dQ1262XYw2xVqCi2CwxU12xRUWT/NVe2Fer
r3DtLKmMD+mbEuaTmcSyFy8RfkT7QvDjJeWbPsRGfSM=
`protect END_PROTECTED
