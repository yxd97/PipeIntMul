library verilog;
use verilog.vl_types.all;
entity X_CARRY4 is
    generic(
        LOC             : string  := "UNPLACED"
    );
    port(
        CO              : out    vl_logic_vector(3 downto 0);
        O               : out    vl_logic_vector(3 downto 0);
        CI              : in     vl_logic;
        CYINIT          : in     vl_logic;
        DI              : in     vl_logic_vector(3 downto 0);
        S               : in     vl_logic_vector(3 downto 0)
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
end X_CARRY4;
