`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8zQVZev2hjh+aQiCdAFh9EDFn61yN03Etz+kCbJx7tLKz1maC/fZ7JAoBs0Zy2T4
/u3Esux3UDMAO6hnDuKewyGF6tUB0rsCkQR29+kSxdJTCCGVK+Zc4TPsaaENrTGa
dEl8vhUGUeNPYZHMhm+vlAK7r+6yD3/64gNezjABkv4lMl9a/rZ62WekGNyLCmqG
1PC/hi+mFnma9j/6VtuHVA0xPPUNSfGwWIBOooa+FCH8O5SmNbxyv4zRLO3VVlyO
4beYGcA/Oyzm/3j0UB0IkV8pQQaQN25S2n0ohXiKnFPQUM2F0xfLFXIXpaIP4Q0O
QJuvLoWSgPyTjryd3yoIk/LHrY//orj+29ZZurhyO/KwmmgWIoCy7QmvSXWZ3tWW
R3G75eA+wjmDZp45Pw86NRDmnmQxJ6u78bnxV6DGAG4mdpmog07X85XGAA/m9JIF
+/dGgnx4AZ07P/ODP5rYOuEqvfJt58U8ZwYjOuQFbGUHEPj9nAPWicTl6BZ0zfNf
6v2u7d3zD+1SUgM1KyPdyEZ1lkr6oQx7HvFZqgZMMdIFbuy3yNNUWtMRzwKDcL/r
9S5BKYV9vyil86aWbD7KtPmPYyGR9R8WiXhGqm3Sb0F20pgKBP7FMFBKZ5vLIDFx
8FWSY1utgRqN7b24jrI7kCyUqjoRVwiB/3JXMv2JYUT2fwH5ONresO6/smL3y/md
YZ6IZmetMcTZl/HO+PrxcYe4DdtGiRWxdXqYIG1038U=
`protect END_PROTECTED
