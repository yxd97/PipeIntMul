`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+iYe1K8K5GC/smi9YI1BoeIbd+09iHYXQ3toVQ7QxELZ/sbaNXfdq7hw+uEUYEA
pGJj2mxX/FaJt5LnofKLsFiqeJK1oNfFxl3X3kLsI2LgUa5JH3ivGnMs5vts19h+
NgUg2RgLH6/EbWN90ShSKypZ/REiB3VPmC9trtLLFhzTjjOyT96M+YaSbSOZ1d6k
8KMeLqXuCmBgKIEOwpR0tgdgyZvklwng93KAbgCUsvNTDj+y4PHAYoy7zSq+3SNW
WLQN4ucZ53lVUQ1nT+EOAZST1Sf7fjqgTdm7/cqfygzhmrRlEYPAikZK38U8lB9+
O+Xbx7GJKp0CHevMaieujurqkWbQkeGgbxF8PCDCxZKhvMs9U8pdInjoQdh0DNW4
lYla20N1+eIceNyQz/GIkA==
`protect END_PROTECTED
