`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sEUDTfjTLGmn3KI+6nHLYWplsz/Y2imLivBTqYjYZyFX36AXTQqYSLFlpzXdY/E2
frxyaRg8cLYE/otm6cMbO1Kd/QLBqySFzcvDvn8InvB5eXjjdjUwwu6UxYALQDHm
TcnHyyzMQ8Yak5P0BLsnrTRbZZw4QVbf8F+VG8H8CkLZqNzHNW4O0Zk121vdPysU
urC//q1hhGnBKV+QIklLqtHPnmUbxyBqySxp3g+3bvtazmF535glmoGWVW74x5A2
VtLQG/kEbC6Lwi0WqxVlckko2yXOBvBGcZfca4/dSB/NzFzyNtsr6yc6LtvjGSFb
O6Ji4J47YdZeEi4EOA9ws7+PGe8/CyCCS9/5vA5gQhnYfHJqGamPxgNXc0mDZFyH
PX/9WR8j7Y+HZizdsGc4d7SujC0RM4byyawRp7l2NuLmhyipeUzW6VMKTtgvL9h8
`protect END_PROTECTED
