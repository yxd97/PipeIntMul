`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ihdur82sjZjn0EW33GoKA4VLBwyUSm/+ZO9kMY8ObJGolOXc9ROA16MdttZPGXKD
uVzR6t6922R6FYuYwDeA6tcDZpKxJBCCG4bVka61U7jB/WTWXm81eeG/eafkbeEp
jZuXqJ6flT8sU1z98paROMN2SkF//2h87RaUkSwmvp7YZzHbHfstiHL04tftTXeN
E4Q8kt9ALHqoUL2CCVbcCosONgviwb529qaUftR7EfgKZ5+t8VODvog7xzCurO7r
eU6aaCk12+xqXENHfLYJpO9F7Bo5DoqvbRldNb6YW92ydwlwuqIFGw+HS70BgOuU
PRbFAHcNiv1/3sq9aNHHHIkoiiIbYpVH93eYqcMddekp/RUwInIChqGhxSMu0ZgA
5rZOEH+XIEWa3kcBF/NFZ1yEJgvJ4nBN8Bh6CHYL2TDif2NLvs7Uev876knAeAlG
3BzCiH8NviEyi8qElVf+1VZGywURmq52l2jsvPG96q1AksOKz+L8N7gdpSh62Xvl
b93PJZ7OYUc1fyIhoLfzsLJtRMsw6mW54iwC7SE/0+xl/Gq+6a7wKIvWLJOIZ+Dt
8LZwHqb9wLY+K0RqRQl73lNkxCwms3kVltuA7FFxk+bXiIvBlAcGQ2pixtOBR/xM
KYCfWTXB95IfPe/ZRQSzLDh7/iNlw7Js463oXbcBMGwN1iXfva+joS9xJNzgeySZ
Ouabdf77C075Jv7QRYdaTqD3YRtojh15k0ZSKD9Mtl0vh7jiHh1cKuZBiB0kFnn9
3x63jaHhR2V1b67NWQ+kGq6yzy77pQJaNvPYidmQIui0Y8eRZIlTJlCh2wIv/YLZ
HSpcq8aLP4AtvYonaoqf0DmvanfcgIRoKo4QjE2diOCSBakcgOU8GtC7QnepklIf
QXNcxVG6YVlAijrF4ndorhD6GnmIVGniHOgDOxsTuV2KyAqSkITAWzDiX8H39OyG
0LcWT09HGYq56EMKPUhYA/jQwy80+XANz8uMT0qxieo9QggvJLO1N9hHT303RBtq
J9Ue6mP2LYZfKd72UPNwSA==
`protect END_PROTECTED
