`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xigme8ts1t3UAOuNpJg01dJFumo5WWmzHCRQO8VZrR3NxwSL9cw0M32l+TNwnnk5
ad0Qklp3Y/Dqz6NDzdB5lj5hh8OPr6NlVsw3yNNSX5YfAavoUmq257FewpqCdpVf
n6zHawhV7bf1ub1Oo4W7I2WCL17HxdehOshvYIpx9LaniCTAGXT4eHeaey5eLEqf
pTXG/TDs06dYdjFYrmVVvtAyBQhrWLJZfLc1zrfaAIS1JJcfW5dzHqqhG0ir/Z3G
2hUJwzkVQ6iKy7UTS4MPK/Y4k7z9lqmopmABcZhaO6k=
`protect END_PROTECTED
