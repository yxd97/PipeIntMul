`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7o2j3i6BashAdcvHM9GSExdrjdDXkSeLw81hmFZcnsRu2g6gsClckVwIy0a+3hqC
b0S3toA5IVBFA9BXGiPkFy+0xRql1unne+hhf6Q4B/HJOT8wEzJLpucvCUXVzpYU
Zq407XSQ4vwtMuaVApqXQMJIH7FCoI/CBM+wiMgusBgk52AifRwObtGrVkoaw/uc
Ue5SoxxzUvEDocfPaN1u8rCzBxupxjeM+cG3nnXFVI53dYr6MbT2tb5lFCQtKmTw
K6l3wjEZ5EL/yetHUwU3c6Iz6sEgpEBXNE9jfYWe3AQM+o6iWVmtgVvTyw9vXK0n
AqMXDeOeRvjMjLMnCT952F4DSmbryKlX5jLRb/8JqA2qDP7Ijy06ALaDNRMdgfsn
AzFOpYbeoRKz2vRPeX9SXvNPchya5a1xHMVDXdqd0SLgR/mID1TMaKdhkm5PHJCx
Dwi0vHTt+aaniOBdXHCxqHHZTniANl3Fwx2vEC1xO353afO72SR85zV+3ij2VO4m
DOdneM3UDhuYs5F5e8QXHWoPAmzaB/7UHqDyuXI9Glrq9SoAxDAuRyb22CVtsLMz
5fizMd10uKzaLw57LdojlHTQ+DVN7rVlqZrL73PzEurR6grFaWTDMoe/HCDMMKg1
pUr2D2WyEzYB1qEx9JgsacxxXtrQDtTVDb5pTb1PzeL3MGd3h9DTpml4WUtDhZuX
d/ryhfWevBwGK2TmkNg6DsNnTRed0V2MUMgYWPYdIRza1+XLaK5kyAK+QVsNGAvQ
pJmMldjt7OlFn4xeMEZFpZtL+BVQt4Ihskaz8GxSk5crtt1JmBAsAzcu+Cd5kSSs
lhCrtwcwc1WrwRGa+bd46fsAdluDJSPjiE2X98C/mFjlAUdxvUc94yA2W9JWt0Y2
tjgJxEAMmq7tcqlfUVMeGbb9yLDK2u367iOuaFeVsIxAkGXZk+ViKpYKDXVboFmE
DzI2DaLuuzeiOLMDsMxjAlttol8i3LAlEku3ltHEG6gtE8ui8hmxWl8licoxxMVM
Zj6KFz1ksM/VsM8dlEYJcG8QTTLuQ2p92hubQ/afb6LdzP0zkr5yQ5sfv6k9iYDd
n/fcWwp+ItAlPLrW/MNgswhCbFl8BWDoRsj5Il8kKiNUIb/EZO/+pKhbY40N6BHv
01hRR/iP3wlrIDKhEI/jkgG6ctQ6ZtGLst4qiEHnkFSt0S8/P48V8s/aGvLbhlM4
UcZU1FBHDqp6oTHhxalsX0MSa5nMkuUVqLzDAFUOFicM9jXJ4qbBg/WubZ2I3KPU
ya17V1u8NBp9PX23FV9eD2Z+SVDrLtaiM58V2hsjQiJULZ0AMrD6C8gsdR92mk+a
L+9XE0tV1iEG85uwl80y4qjdkOVxnEb5WPKHdPdoRc9mwN8RemUjYZdnGocD8D/v
YqZ2vW/GenCOede9Z+nHE5yIg7gHF4HMQ6SvquEUr/N4MLU74ZZyr4+fGfpwDKGN
ji/RxiQVACnyamuDyRgj/YUBC0OTxCEcCZC3FkSn3zoxeYH18toNBLmlyVpCOWxV
t30q4prhwDV7bHd7OZIVPmpy5CP1VwSdQx33cv9X1QtT/qeb94GAPMW30PX1vnJv
k8eabiNOZ+3Qkfgtl1sLn/zhZEZbAH030aNmONfOEqWj4mTWTwClPOltq0+d6gcd
ZeFk42WDbv6gBr5KIzjU2xke8sYkvAPcoJy8jZZWCijuPdJmkQN3mUqH03Bl/w54
wAjBAGeyI5jOlLoz3bPLUW06696zqJO7ewBCa+5Tt0KAmZaH9uJcFWqLuNvecKlu
HS8ELuk2yRb/yNmuQ/osx66Tgb6FrsLdata40aNsgyt6iyPXl6K9E0QDJ5vNrR1q
7HiCB+0lhhzjgMaFukItleZoFuGveiFLvjmwOKXM2fcdX10VsHvhtb5D1TWxmClT
Sc8xipcY4/6pZqqjS8PTUIVEciTcspy5uHg5WMHjQdXrpvosl2X7CaCJn3KIhWdk
CG+7IMk50xefneIU+1tZGCgXgqUQx2J4d5sljxj9zpgKMyncTezeQNAHzPFMca2D
8iDGtG29spsMM1INAKgTN5NGM5OfLaDHPZ15SZdmV3LVNRaw5AmgflUo2XU4SlEj
ZIoAfim3gIX19wWt2G2b7CoxAmA6j/Oxpniu5nnWgbj8ypw0bTkQtVXsJpVpbprO
lmi2ryiSvXvrssjmnp/hEgN0pNuKf9SqrbU55bZGQ3iKpe8QHCHMZDFkbIBd40xS
zfDwvfq1Ady7in27dcDprkrYqs1LayF0vpQWnnm1G24zNfOdciXq4vbkiHkcv+9f
NkcMpwM49RtKwr7rSsGx4RNbDsBmUJ8WSS/bQW+fItAFUDDH5CSB2c2A0yGtxweG
bnretodc8Zi1nQ7o6seTZLO2oCTMxDnS53eMjdqkQQRo4eNkaAwUXENXR2snXUOt
4xAOBjxlyZ/2nXsY1I2MxBdC50mBpPCVP5a60XJTwudryEzUTC4XR+vn+baLFdo7
qMaPRhJQXJZbwOMi8vD5v0TqRjPPs3j89M5SG7NjH3fhO21PNJBJiAteQQD+eA0t
n5x7iSUGuoD+JRLQqOHD4AUWSf46NUEA/oQ+iGmX8joRbRrw88fH53wmmSxin2pW
6v1ECvh6EcUf9Z25TVuaLyS4h3zManyBNNzRH6fvb28XZzHeoTwzp5PLTVsoxxww
Nnc8v0x+uA436ZQevB2ht6er50Q63QDC6oJPT8NzWNIMJlJ90BaAoN3i4I2tKJN0
OYz1LGOPXBeE9ZjkegsTwNDtzcIBGuDpEU2y6OUtKbtyOLCqChTpv8dvGu6n9EoA
eDnWSYntQv1xGw0YOuu3l80dmXHl6tsIsShs1ROze1CoBhleln4cLcgu2it3vsoC
AMXz9xtolxScgNf40GUlj4ORwi8qCCrvXHgG00eaZfPFQPmplUH0R9uOcQglksgG
JsHF8p/+9kpHh1/AbB7v3W+WDdK+wxwYLqZYUtLUeOfov0XwoFfbAvnW1PMbz+s4
ZwVIFd/hjzl2O4TnfU6Ck0kLV/zwYy4BBjNGpybwabdRVBjghjZcTnLQwapFtaXB
0kH4vOtPuFrUJkdovHCIMIxO8pHxNm2OOoYHEW3Dxd/iGO8CEM4QkTbF3Xvh/6Nd
ZoQq0mHi7iNIElhQeSw7OpJVLcuYdahClKmPPtm8oxzcv8l5jh17oJ27oK243UC9
gbQtc4A9QF0xI35sTaCPdehvI17VhXWC2oIEmZUy4THc8Tl9NXB4B5o6/FRjC8ul
fN/4g6Ak5ltW6xP1SaQbT9Nj1kJfSmNcHL0qCW7hximneuMyW1DwOfS4mK/OgkEe
oiH8QcvXvbeIF+ndMErGfn+e1uGT+iJasylO70VM1iE/L42zLkLOf13ObpENDrgS
HvgIBDJb/920i5ErzKhehje4HIvW/9OUHFiR9zzrjYwJxJVuj2dYukqeKC2nn2Yc
7MBZQu+KCIt/HvygwqN3mKruJ+Jr4vJl39e390MdT1yt+zbNWMm0fkACRV1zaq6W
bhTzbxOPyyV7aFeo/Lo6iz167rrpNCBdV0Zmpwzb4EMw/kJ2E/laMh5RjjlGrB2J
9/TDpTfwyN049+ZUXcuhvVSeTtdFWWFxZhf+KuwnkyG70br+YyxMKWQcHiQkoRMZ
cUB7DS9LBGCYswNq65dMlGlXn57B6SUbig2lHKJ76Fui98lINlJQgs+vXrBQ7bA+
VQvuVOgooz08yYv3QBeMsb4nqeFdoE8pwIPKgBYdPnvJBt5Ay5iv9QubC7b7BQ3z
UBqEcMPTZhueai4iosB5YLMZggbpAk99ra0H2t8a/03CUPgqaLJgKfQrIu0c2976
lOQNI7WjpoCIfZkIKSwvxfYTC8khnP1xvHKX7exxHIczUeVPMc9b2TzIeMe+VlBZ
OnNlXGuJ7OVCjuJsGkmP0EInRvonqNt2qx4vBqdW/pVauimOhcYUX1IN7AZxU8Kb
RjBG3vE8ZtHk6vweqBK2Gh6BUPLo1rgDp3i+6HjRVx74jaDY/pA5wRx9Gyj+EYJD
2JAzIaVhU33VbBlj4uIc0mu35GrKPfkFEuFBIhkwHn0/w0YqU/jLkN+6Pso3Rtzm
IGv2O1zrfi37kMcxttn1wcoMZERcmBz/8Ln83lx72snkZ06QTic+YyTAIMhgiZub
hSrMVOqtfTkK7vx9w+wcuzT//MLlLCZHXn1U2MOI7wMwzEHi959HCwhOy5Tn0bPW
Og5lHxdBHphRbrxpNMyZKcRK47tJ2LE9bvjWe99P3/QUvM3O/9owqUon8ysilmZX
4Kcn+qzYDIuxprxN+eWSkyynO8FcKxnl/CbyqLk94iDaL0NE9winK1O+Y4Y8EoCZ
LjNWkhsUG3l7zGPWjP8cdh74qW+Y2VT5zvYCXnd8+eWUJEo8PRSjzGyVEm6naN6g
EOwxMGvEkSYiS4kw5ueO65G28336Z/T+Vwoifhb4jsH4XsSOoIGZax4GjpJb80z+
nZOTX9E5TsaxRSpnpkUMU6sN3w5rC0L1KzHwx018BTAvt4lcDLYySjZQFbnkOqIy
R4u5fSeiUIiKI2DaORWsUQ==
`protect END_PROTECTED
