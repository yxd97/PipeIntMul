`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KwBwZhR9a5+Fj+2UTyb6MFAbxI84iGkO1DTABkviAwYxf4WdjGulHLzQbyIQDKp/
E2WqmZUql2jtO+fUMNPy8GxhzY/sqINeIZY1hz2WJPAZ+5lcQfF6q6uDr5OETIsU
tcn7TwH9Djbo5ry4rzloJ2FgI+lravp5qWYAUakPojaMH8WdkHglfu2hZethzAeo
bYt/kElzSS8myaKIqmILkmon/A2RosIzjuQf0FBfz1oiSTCO3NEyzj4tNljLLhhD
xIpb46cOhR/0SGSjQpMxEpXfM7al9UsSdUN1QGOe34Y+qFk463R65pSCyZbaQsh3
uDBcGP/PVSHnC+CV61uaxyGp5UVRwBwF5U97TkWAF0sOvZ8bYM3s4NFR6cewDdoz
fXTwkhF8c+0YElTqh1+4627dFI7NViuICz1LGDP/CFX+rf2Cvxk2Kdx4XsnGW95p
r03s6c5+C/2jKRv4QfFhZojVtJVvv7+VViuQejQxntDqxPKi7TuE4RlLsbu0Fn+L
SJGHEZIKzfF3aU1Gl3fnoq0vOBsYkZt2Z5WlgsdTqOFcwhry3tSr8A+JOdtWB6oK
D4gAbolqeCyx9wH8NBrjpCPOwJXwPjj4SJ4NvMiwkpaJyRPPDD6FVoKkahpXnPlf
UsSeh7vd89cZyqY0tpR7bsn/YlHKYs8/dv8lSI8YtZvvAYU1VpgRg24oKxpYsDgu
Fe0sbj89V0NzGjBshimsBCt5fH4fLfNVIqFO6ig02468WhCKblCEjI61xGG4oq6f
VdoSEO9rTOudhSOTYIpTKKvPVrrimo1fwHZhUBqjQrB23F8nB3Kmbq6VSXMgROLc
TTcKQ8ReNJLnbAkr3eBGZFe1csopxmdoHcxN/LYTVvquxGfaccK5Xq7uIGwsNurP
h96s1igawi8VgRgvGLH1ppDZ20Q9l5L0BRprjhtrTnZptvaBVHGMwJSmekEIfKR2
XVQJbEg9SsIliy4hyFWByqvj4nI/tbv5b9IitqKNuP4=
`protect END_PROTECTED
