`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OldnfBljgWYB5CsiVyuWtt/Qo7zuLISiGtC7F2iO78DUpfwjkHP7xXgfFIkap1bD
nbKJACNZECrb9l8VxxutBegijEKUUKWusPgkXFEMCK9D8c1SCtbAIhdOQfFny+G/
d7uggaAQCJjMYl85OlZyNfvTDZbKZ8oNrLgFC1OcADsDjvJ9ta+aEre0/fCq2/lE
0bRfqke+3F+VPSwoBEFD1EzcDQAW1IvMERzL7Xecyg6cEMbPm7dc5MTpehYgbKbb
1nvXfoEXRzzjpodTm5WSR1UTh6qS5Bv6s5a7hn+2P/19yoORT5LekrsDJR+o72I2
QWVAv6kzY4T1JnpTGQwW4A==
`protect END_PROTECTED
