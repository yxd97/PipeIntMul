`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
06O+nvjIjtfiEoC4Lv8+b4QGa4MWkUhzktNha8MKdNUf9FQzjAmelbn3c+2dFc56
03yrewb+ITnO0b82FPsPm1xdrSTa8ETtae7wht51QQ6P4rDQH+sPYFJPUQf/H1HL
O3TGZRrcUdTz4jcM3k94I0cvY+W2Mikyr8v6AxeTnVRQLiAU2dQb1iE4SiEw3pkW
p3xhMryO32KjLuNbSwDJT/53xrDH5dwrF38fiU5B1n2uq8+sd02B4hab6eT8kzGg
v4o653+MbAV58y5TmX7VRyeGDdHdqSSN1RQgo6QHuO2cm0ffTigen/wDn7AU6m65
Vk2nfwbXXR9IxRJDdru5XFlgoS8QlkHW/Pag9hEM+wSEnPzB1kxeaQxsghocro9o
sB02sRFVJfxq8ekh3jx/Aya7pRS9nbEPppdAnDJGa70gF5GMU+sQVo2D2LPTqIcV
DMmIizcu22WcXzfWiOkWqahET1OOWBU0E3mKsqvDj0AFvSwkB9Gv/YKIt8aALZex
meDuu11kHQoWOHmWj9mPK60ozbx1B16jrntbqoEvi9FXjS2qUNTQZhDiqL9IdXIx
pGsfSQzs7xIFJ5egyoCVWtDMUEinQ9HNqZf8M497S7VYf+tR1CqBAxZNfhwKnbUk
8FJ738wIzThVJ/0wk0ADq4sM84IliFcnNHE9Ts+DkOwmWWn4jCsiH0d12wgzXUr8
IT2z3zMhl5dYbOPPx/ZbkkCrIvQzCK9bIipCuKSPaRSwjgtK8pnhVW8OPqpbmve0
YV4/1ZMHSoKM65LBzo/swg==
`protect END_PROTECTED
