`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZGudSF42UulX3BRyIwGVFprBwmBPI68u08Ccc21VfdQhQIq68Inp1LoWuE5Wr9kV
2ma4SOonNd6ToKuW2jTEBe/MRX1UZJ8naCqZtuFHTAvIZ1XAy3NHZfM+PTF1gR/r
UOZUACXopO30h1ezTSAZWcc4luAFAeD0X5rX0SK0Gb7iUi8ctCOJ74vRFsarPs9E
D9Yxr5FH2TY8DWS6n+9rZdWjt+qtfqtXntII5r7zFzT8Wz/iaNXJ8w2DxoqtvH7w
W6VgkOu6JH9cfJ2+H6+j6qTkrSB8TfvcIjOomcgSSpk+JRlKA677ghdSKzuW5Xvg
0fcZv/1apw+9xRVTxjqG6gum6yZFUKaiCHXfvFHSm7gh5pOwxrOp0rmWw9yrf37h
0KJQ/0GFQHcj10h5jeiWkVG32qd6QhWAnIMlXVgdz6o0tn4/Tf38yyxP73oOsX6r
YW+m8lPRvy4jBj+OSRJHiqO0GgwIky9o+ba/649KjZs=
`protect END_PROTECTED
