`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w4nbXlJpr6pvp7njPfR2mw/6Jzott6Y7+KV/8QRVeQKxFI8qHm0Ibzwfl4zA/r3W
aX5684iDrg1H08tY5oV6ojctdQawClBXkZdQvmHELbTFUTn9BIAfSCI3evlEdLdL
P5iiShYPoKlcqqK7iTMZJqG/Xkw5Ml1DUN4/NDv4BAxMPNmcmJuYLRERNKeDFF4K
+8HISEYzBwoFpCRvbmHQ2SFJOff8MzLpUEZgcIHJbsyuY79FAO5nUdg7thwyJQBI
ZdwKUkd1hp+Dvu3LgnlIfB/tBdchzcosJ2fvrlxOzK/REwhKacnDUVr2ORVmva2e
or5+LQM8qam/VK5vBgygyNsPQl7+guCV7owVuqsKZ20qHMrZSyi8W1YSq2vZiapo
j6g3RsMklXFAkL1o6qT2yA==
`protect END_PROTECTED
