`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mfhs2Y9lCHs2G3qsAi+gi1IQ96c3co3TjxJUsHxRlK5o56ynKlVxumjuUnWzDxIZ
XJcdd/P6HE9KNwA2MBx5U/rq+6KKpyrFMje2jJR8k7GKSJL9NC2V11eru/in1+M7
PrrMCS5jffEKAsgyI2SG+gF22sy+RBczuD1SD+9W9g5ppXTvjA3ga2T9ZemAZfCp
1BSt2zP0StLvXbMbvlC9I89utE0x8Ks4Puf/eoKLQKamBj/OEZPOLHo760C+R32Q
WXWP69K56XEvdCyU/bAjaSlUqrjw/Klc2HxqR7JPJ0xfB7hlLvNcLXbaAa84P0fZ
cdp4jRVbfqP8oPtiTMNfg0ZhifiVBtAotHkPDWhosPQUTQdpTGRs+kyvfWo+jkiL
g33fexE7rY98bVS+wvAVdP+H3yqfR2fekrUXUazyRz2C1/H59ZcOkF9WRTik9edm
NMKzyz3kYV8FNHtSxBWDKLOQR7NMnkUPJMfAfPzk6S3hBHJsPET9JGzpC0zXEBBw
qRKlxl4oSYKG0ih+Rw/o/w==
`protect END_PROTECTED
