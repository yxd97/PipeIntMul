`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CDuuqMYSadJUFjRRiom5EUGpWSJVBPiHbkZdKIRnzAvxdlEBEHNIQg0kfMb8CDgP
fSs8BDG6Q2EmArkuLL99m57x8WjnQ2oK7G0aVRjGZ1PPilMQHXROM0cmTROf32cg
gia2LVGMYkza4/OreLKbLo2vDfpUCl/p+CAy1zPMZU8+zakO6LL20TgrGj7NfrhR
HAVa2OxsM7g8QkiNGyOiIB62cdgsiYSTFFlqRw3ft8qAmfNSsJvWO/aZLurAmjTV
pHe8HmkBgnOjLyMPq7zyBA==
`protect END_PROTECTED
