`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ccnJZsVFXHOER2U3VWiB/IJ/JLn1ETv4iR5ekG6PsXzLwXhtp0cMG9VcGvaEKER
hVmuSUHPzm19rkWMhLdkKvFC81Nkh7HVeXxrqmzeXvZGGxeUSs6JJZv+yNRrYes4
ODsBdwWYUt24OcfzsP6rrvA0JQGl5nzjGGyWkYGtvyO1AN+XtqhSIRJhlkQuSEYs
L37GpJOKZBY4boRgGLVmFri4LFZeLqpWV5ZcG4kqye96pa4yGZZ3Rij3WEkhTEDI
2MST4EU9xw6pyT45AyTCkgGs+WehLPll+2XspzF6Qw/QSgL2Ju3P+Fd5OArqCgR1
jXs6dNfhwpk5fWX8NRHGxmU+E/yjK2AK/4KSWt5VpVXuMzMD22kGuWq3jMnnV1QD
uGmXkR6PLHkOgkMpUqw4Vh0Bv3YVS6vHuwsu5d97NklWEytR+B8OxA9bO9dCBLoq
r3T5vRylZ/pJi5kCe1boyIdcjzo5ilStDyEbAu8guvB7EhdqQRtpBBD08K1TBrw2
fDMMTarv40gOVnej3WGravnVqOak+xu8jabtOb84J386AHjGeCX4DFxQtAsusB9+
X65y9OICq/GIDhM3KHy9iGOip1Ghu93ALhL5teNw6KKpM0W4gls2w3LV4QAmFhqm
WiXpd38o9JKWHMZRI4Arsf6GOdeyt6lyyLbfEhiLXU0yozJ2qwOu5Y+00tivTtFD
7Pxak8QTpePJL6iZYbvvyPlqsz9zl70HHyPGpnF+RjymxEEUx8sX273JA4zIzCpi
Aiv8DMow65maxG9PGdCRSD89A5oSYDEAkJ5yaavWe/oS3Sy1jW9ZwJluO0OZ5b6V
Ch5nClsp3VYfY4z78SYf+0xIsLIbcsvQDHf2/n0OhmZWB1UU4+PLGtvytW/fsUx3
Grh6K30+Dg6TVEfseRMifxoseq6FWS5CDgndNFfAZ4q2Mew3EZ5m3fmEcYRujtB2
+A/D0ckJsQUMtdpDt/Ia98D/xSSUS/MbyM8ACsIzlwPFkF1JR3imGt2A7yAXlRcw
M2DX11agJWdogea97Bq+8TtBzLvOUzDYqGvXwIyuUSfIPDfWkh1aO6fym1mZhRee
VHlslMonHJFCjt7i9IS7otPJc4GIoPSWOlfSvko1S5uODLIUMvJLhVLWfL3v6/W9
RkWq28Slx+mpo6p4AFdqtfAVhqLZ0P07Xlh+bEvxhR9ohnJSBaIVwYANIuXAFz16
s2FUY4uH+zWTKU4Ti0BxY5DViNZLvCj1me1KEWWMW4UIkbJkecOX6qfn470b8nvH
DFroP4VzGePZTuxhBCWA81ePuX2BOHSxjaYW54ldJBU2Psl+CMHXa61i2Dj9X8Vf
Ml/45d+8QvyYJehR1wcIrOiwjOpi9JX8pAJtGcvqExE+VnO4poAquiIKP6szHjwx
lXnv5cz272+JMBQ9lSSXcw7aLdRdP80z4Ci0VvAamSmNAPuZRvSDCTEp53KVbLnQ
h0GYgcY+aRAX/qRHjtFn7TeIerEdFwbBCJHi7GQjYlyajIZBxhWrI97+1DmgHtcM
tP5rcNB+15SV0AoHl8lc+6pmtd2l/Q1KDIFHwQ7a0OXP9MJ437FRmxy10T6eBvgH
XaHhvoOi7FiuAGv6KyJ7SE4srKMMnaE84iqbgCYEkDy6kX83D9qJ1ICl+UKt0mtB
pg+dPM/jeui0LWGL8uM91/04VwQYL0aOauj8b98IGFUj6QCi14Noc7xFg7k5UEMX
zZgqjIKENYraQtAk27BTgfQtAgGXzX9obAtjhqq+knc=
`protect END_PROTECTED
