`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g6g9KLme6EH5AKIpFi/VxdA6Xu0WISKCnC0LvTUt0boJXOKJ04ScTWFOIXcD/c7+
sCs4m9mmSSALNqKOWtYH96J96SgUX0NuRLBn2/sgHFLPQOJiPtNL+eYlNWMyc3j6
B3Sj1Tu3JUBpmX4uv5PT3OY/keE9lCqkWKmFtqpWiqmsLAWboD+ai80ZbP+mrasV
XH0k8rR1ugznaw9hEyqfvxwN6JW6x2wdCIwHxsuq99AVXNl8+OU7OSGtAwbCF5eL
X0rx+OT535Vs0/8xQ0dRzgXlMvDelixWLjMb+eeGAFqHhAp62iq9V7WgQWskNReD
JU+lk0fH0HuVSlHkm/rGU6bXdPdf8ghr70xLn+XjHGOKZtZty4VNzN8wWE+Gb+gz
Fz3NDY7HvGxryzAC7aGWM8Ki5lT4XFARunjsq7PkC60HLBDyQKrXN8OxWApQcWFq
aV9xjQRf8h7dGx+C3rUe2ig/dysjApcgigkuNKUyOlrozHua0hEKRnhrIHhxFkv3
QQLXDpjWgk4T691N5UYEi//s1uSoSox0OzyP6vGX4gXUQUjw3Zz6RRZ+JFrCxsDW
AlZxtOJ01legijmt1EOb9VnOE3Kt4FjvR/x1JKek9kg=
`protect END_PROTECTED
