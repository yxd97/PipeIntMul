`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ealFbMmDaw3knvKwq1uSgMenppTjEjOm0IeDfl0x5raA4iCTzSNVuVIa38Hb5KP
gYqo2xsPtSJ6Lujq1/fkomN/nTEcHlaZJ3TgC84bzbuBKY4GJPNjDxWS624C6KAp
yoCR7qknHMKtIMDn4Mm3h2sqIM1BwOnkd9aQnDTh01LGYO60TPPCe7s5VlbULQq8
ePbBxjdXjOtAF/fz0XJWeYKaNFgL7KXbUCMZmIXxuvxgnio8Z4CGiZkc1tUmVwK+
l/2IUT9HWOqYsFiuJIrrFn5ZAX4aQPeu1gN1p2kp5Q4hdqVS897T6jkQ5pAIU7XN
Xj7XfWnjLUXYnZYiMfFP6FNGtjHR4Iqfp3+UTlgAHARLlVb7wRTukHQDnJyhmlBd
JRpA2So9xx/xLtSaxuLrouYH+c+1Sk5uDuG+dxaa4h4ifMKRj0ll8vL+uC3TeUKW
bj2yJ0WwHeL5mm5JFbptfSiWVN89dhHY9O7WilcuxHOb7karDjPxSFxZkLWqbeNs
DetkKr+9xpsw8UWK4offb9CieQ6C8fWw8ZZcVlmV/Tr8RoiqBwrWPR+Dwy/Uszf4
3uqnhGkTY4dnhYiJEowKh9gtVP/bI+edbQF+KAlt4KorItgRfq/eC19GSm8ui9ol
ybi7FjNjmp7VjRPplOonAo4uPPcdZqKfjPBa9H/wo8RCpXMIK//CosjVxBrcHi/v
yMo9E8YgEbLtVZKlMT4CKUFnMzSnPzu/psXwlw0hHbxuZ/y6s9ydlyeVOc2xBQFu
/J9N1Wihv3LnlPZ0IGEdZmOGDT3G096GFTqWrnHcCDHtS3G9hV/ZAi7b+N09N/CH
7+OxOkq6LGtr8/lPIM4koUeLCBn06bL76GwNmq5petBpJXoPgUXNAQX8jqaaGgjM
sbsLxlsNQBlX47VpKnElchGrc7Vj3Fc30OcL7rLiYp9qXmAR6+wTbTHbzrvbQqbU
2C/+J0PuwXzzb37RgmFMsMTN+amp9kFfFbrci5cHC5z4EvdxQmIy1bBV8Hm/AM0U
ceeDRDgNv1s1AIKM9re+xg/ejp9TXYM3+auusvg/oG1N5eHXncFqXQWptZQcQKpW
pMBzx4FhkZ2hMceB7G+KpojEYXKe7flAijSscP2Q0+A=
`protect END_PROTECTED
