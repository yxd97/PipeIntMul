`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CpTMTBNNDKyRuDFTeT0kyQKYzRxdX8rTcoKRioN9lcVPwJiJGm2haiuZ4104r5n/
t6CLdKKkAK3amtF+nucOWpSr8etAeaz7NYSWotQB8ZJuN7VI1EDj0X2pCiOcWNXO
KXyUVo4NJuOf5KJH/w5mtR49A+ImsAudybEdfSNUnHBqiLYffp8NxQ7OK/XB4QXF
obK5srio1b1niz8mmcCfm3F0V/WOYHjargMPd73Dy5Yxgtw4VZGT5dep9ZuDNar6
7/2NE+8PkwJ/e2+3KD5Hd0COVboF4PNbyFDmq9vgdbReKTFdvSjKfJa9bX7/zhep
P7CuIYDNwsNORPoq+ye8owkuILjNATIAmgChBD4O1a+HEm+pKQyDL8ZtvYo1d4c+
T2OBoHdekXhk413ZllvFQpITLgkpO6/VE3Vd1UgeBGcj7hKSghMrSpdtFBKX2Ub+
8vTt5OCqbb4uXAO8mUMnxZvBvey94yq9+t2xQyZqzuvqrfes3Df0GIbNHlHHQMb/
WmwTP1+yWY3wQslDVaOCOYF63If5Z3WWiop+CS6PwP0Km8MAu1n0ua4O5N5sXWOu
3F47BdjbpNlzr17IN4X5KhKP1BUycvK3/EWqpCrnvMYw12tWVrhjuuHpacRz2Kbg
Fw9T/4Z+xIQvLyXrPkNaRZsfkAte4b77bjjjEvND9gP57VjPZNHL2jNFugJBNZF1
qLfPVYyrKG2AqayVbJ0DUcGQPibyO0ajY03QfZn+/C+zr+nD+bXWMqYilBEa+21Q
duF66jAjhgVwP2yCDcoPHZVrQr1v3/yDRu2WZD1eZe+zMEQY35c1V4291hph0JgJ
w/ibjMLf0Jv7/uCP+md//QwLt+RUicJYP7W5ZLecCLvkRW6njSl7rPmv61E9S9zy
yUXbwkO2HhwsuYv8Xtl4Ovxtur7KeG8PiWa6Oo7g4OX2Bq3NJ+dZZoOSgB48leWw
`protect END_PROTECTED
