`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
viFKITug3cfW0Huuzd/G2XjEhFobln3htQMpLVh6h9hOrlo1OK95l+VkSVFPewg1
jHK9Ncnptq6upaPk4d7XA5iH0nua2xXwQBQz269DMtwqbfkkgQk0IM79VdRkHWIt
hsQni9Ut4LsokUGSV04O9ORXlceETUqfG17fHnmywIGw7dqQjiv7VBoStRyOpnrF
mEpFedJdG4M+9eVoRMNh4svRtmdIRaSF+h5vVLXNdjwfnINLlmqDEtCI4GxuP903
M8tfRbf6YtfNBme57x0FBzDflbI84+s9rjtar2AiNLrcWS1B1F+iGpWsGTfZBEqW
Dfc54VsJzT0bcww63+TZYFb7S09A5RUc8i7UI99S7vk5UIUHESqKY0chtHEw+teK
EiunmyzqhhgyFTdutJQcS1JIfpyzbriYhudPMl8cmxPlemBAz011cCPxe11L0q1j
mNHJSqaZ+w/0KVBQVnTQdGdTHHxyZD7CD/TR/Sc+sAB4ZygKS0/2NvMxANEx6Qmn
/X8zxgl4fem9IC7t8PUJ6Y+1X7xEpZi2Vrb+i5zUw06c0H0SHlP3e3p2PhGcb4vo
`protect END_PROTECTED
