`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRveI8WnEeFRPP9P2fMiwCRtg/RCOMYlXF6pOwxt0a981j6sEuhZTDA6hAb9XsP3
0+ZogF88iv//863JGpgrr0D7x0dk7N6+efqBFarSElodX0AcDSfyeb4uHhyeyse0
7EehFc6lC+7e5W8pXT+sN79XaFwCHvcmQzt+iCF+UFVoucluPbvJn15MKJbAX9ry
H+Grg2q8v5HkzT9ki7zkAjoAWaYTzQczqC2/AUiyJxBOOUCRxipQsR+Qb21/hAyr
i8b0kFkRH57RN3+d5sT3RDqC59HAaYbbI6DxDS9NYVygXQYzjuzUy9P2+VJ99SjA
jvjrMwfHfQVRAby17kzVvA==
`protect END_PROTECTED
