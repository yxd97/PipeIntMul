`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RV7jci/oXUEbzgQhAhyRhceh+ra+xvIPedD+Xv1483G8gwb+S6S4nrX3P/leSmUn
H1IFWYyDFz36bzk+rPfiXe08LpKzCHn6/kwjph5ZZ7GY/ULV1AOND23HfVxfok/l
MMI+TQiuU1/+GsQsiJQ3MPhvksKXT9EVmWP8xoAHycSmDwYUl+js7z3mNEbfu7de
tv9a2b7gUpLpIoe2SxtEMM0yARUlaFpGvoh49SdTHJCiyGc2YFfV+3VG8cNGHBUF
JdJ8acng3MQUyzt4Djx4GdGaxTGK74LlDqRZWENN6x0MXbzqt0pNY312dpEkf4ZM
eP0FHl3tiv+o45Ttar8xxYzcmLYAXxCPcBOEUzu6JfB7F7nFNY3Xpad1mRezaWcx
3OKOPXjJCJ9KdqNviCi2yQTsRsnmRve1yW1Ps6M3aXyByzFgk+h16k+4OZDGy9Qx
`protect END_PROTECTED
