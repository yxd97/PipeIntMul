`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7Oh77JOjKdm21cRBr81qnncmkcIxy7RVJQ/XiB3xy5yVEHNEK5jYAO+IsHgA/1N
XRZLstN6Y+jqg5QZZxqUjQSLTaj5HkUgBUzDhvA8KM/PKZhGEV4dCUbNa0ut8uRw
F6OycCd9vX8W8TUXclxWxz/zQ688Wm/vqGiE9p7HCYT9Ts0WiaS7U9/IvcBByuVx
MYxow3DUxBxOUVy72oHh0RaaYVzpb3doBzYvWlUexVF2eMsnAIzrI1ARTu6Y6vxR
bQscIspq+iP8Ead0QL4OM1q5EqfrT4hSR7GxFXBr/XPmrJ4qZo4A2Fl3B/zBHtP3
M7A0acOAwWmXBTEff2029R83Ny8NnR2in8wtu29+XOA23nWagzvU3YzhT/axLbKS
+lP/FkzVU3ui+uL5mp7Qsq+XMTw6HJK7GuYIKoHjUkE71LGP4RnnhucA7KfKHje3
xVNt+2/0ZYcJWwSXi6Gx51skyI/hQWSe5Cwhxc3TvH2ByDh4UGreFYoG3l/gt0kN
tXB5448QeZZrvCoelDiz3ydoPZjuH11HMKX1LkJss/cIeZngzqaA0Fz7YPLV8iYQ
oEnzimBg2L//OInyHJOjBxxIzNDRfUSFJ5dTKHzAvXDkFt+tnZMZdCpGA8OuOFiP
+xjRQ4SShQ+6JByQV5oeZPkys7dhH2iw5sT+A9sDWbl+C/cQ2UcQPrCPVkOUw00e
9729/OsNHNOOQnirFmyQo7uDBWtisqO0oMvubSbL+ThLDk3N4XVVSyzrs+tMj5mE
/+yKKN84jA6vXqiohYorNR24GxmABlqJmIU4Fy69u5dtTovkm75GCqt0K7bjpSgU
2nzbu914XLb8kFq5dlgBI1eXyBthrvm1s/XYsjujGk8LWwEmWfIt3fORS8n6S3aC
raXtEOml8J4a2nJPDbad7GztDkdOkx6QCsFvUFxh9Q0=
`protect END_PROTECTED
