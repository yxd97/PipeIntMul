`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t9T2tGCt+91z35K476Z43rfmPwnk0q5zsUXXGJwB++ePNVbGI0mP6tRBTyfuRRzs
2fP0dowUeYy2QPLbiCsw+NLkNNT+FFE2XaMX84f2NTkSaH3q1xkqUBrx47DmCWQl
aXXME9fidtB/ORiM0D2615zayRd4FfuzhtnASOEPfe4nzuCdhALEMv8kTRasgvZ8
Y00bZUzRB+SsJ+VjB5nBsMx3QmMq1ydmn0prBC1V1r2IrqM8SvYOqrPNG99Hvopy
qPI0FcAyKep45Ms9IDTxYFG7KxPObh1wcQJDsUwU/O3GAgnsBiy8jId5Y+r2newe
PbpecsW+cySIiYs9LzbBA2hWWYpD1EPlljj8AfluJGTtmL3FgosMozwNJpgM1bAC
`protect END_PROTECTED
