`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ozKU0wGgH73qOddkecZcwo8ywcx2hFJxmvawr9ZPUTlfkG8bDVJj/TcZbWzFLv4W
o1wPYV32zf8rPCZsEN13Z0aDb/LdyXfEYOC59cImt/cIjsrktd2KA7wvSkJNmAUa
hcSeU/Jj987xZML3rcBvOutDI3cxhToGpIyVwnwOuyQSNcK6LbaUOYqtNgMy4q4Q
ugSjeTfkrijWhI35AoenpeaxLjKS/wMz2+zKN9heJGKb2uoyxbhXPG/WDrnmdzhW
9xfZHFKpMfhFaaTso40IWnU+DH7cBn4/j3BDdy7F6sND7V00BPavLZvK2VxMpj2E
WsG5reFC4QNlVOxPIbGm9WkzkPHZHt3nS2dv2wlG6KIJDt+hFdefpXQ8Qf2IznOQ
OdF+oq8oTRO7xJIQU1hoOnSE57ou6rg7TQGyDm6jZaF+8W2UAZCWuKwVo2o1bDCm
LYd2bJ6CtvGkl161FMn/ww==
`protect END_PROTECTED
