`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
//kl6qUtbbbln2v7n54lLLbtMW3zYPhGoOkku7apP+hsiWfdl5QUmc7sFSdKed81
fTPMFz8TWdiXtmUN+idpgpRzqOojhVwcxKhmi9bxM2U8TtIsQYd8JPdDtVLYChT7
QufxHu3Hn6ZovWuVtj5YfX3f/WqTTb+EwawcW2mWHaN6ilNLsin8HOQLrHw6/bV5
4GKU38mwtF0xQWiL0OSAfSJ8CtROMG2bXFZNbOHsfKc7et7jvfXbm7P/qWEV3ktS
KdhxzL5KTevBODfl6uqhZvu4dr97+5Wefo5IcT7PeRSczNYieJYakShB42DN2kI/
rJS38YS5Nv1thVgz85SdzS0+kVfpukMWoXYjsTRDY9F1Bw54fcWI1l0F0k+XNpYe
WbhzVHh1ZBBtjOGgGu4uaZlNVQaVcnvZrT5TOnq9oy3E/866KgGPwpR6PiBgC8Xg
v2w1tN0uLvmqbELtuh6Vr1DZUZYDpzJbL5R6SvOxqdxhoVCBYXC7NfrxcVLgJK7Y
myIAnitOsCjrJrwVgJUKpaSS3OpbxGbIWpV8pz1RQGABoylBNsuBpd+ovfaW6ojo
Pew10JnlrKMn4zLVOOkdtaDyHzGUFIfRj+MR4osVCXy3aBWwqGwdQ/oHi8iUjVnB
vSqGgVmFXGxW5BW5qJlBdN+OceYAAAk6TZG8NG5dh6zXZ3P+2K5qMJaLDwZ7H+op
qjlEQPHN9JTjNpd5DQv/FIXHKHErDONsEHEhWy0TcT7LdEGqg6ZUsltWqcRMOWsz
CuC7z7IIkDnGGtem4I7YfEzSB7dQI+OW0TzZKGkZLEFhmhs9TPXFWZf/2FvihJ1P
ZE+dhgF5h7SPbK+IqjI7WzCywhQQzBL/0oFBYRbHJhLa+A+IbYj6w3w0f6v4ae4T
CfMwwCCVqLR+eOS/cMXWi9r20JA0z8qNQGPrkZ5noe1no0McFrSv+6KlziyVnGWO
T2AOjSU/dRsVpxmMdQEdp+RywOlVcoYrG/YGMvF9tRHm0FI740GOsWmG8+z6KRMy
Mcso8e1bLIqbpo4dqAKIKgG2OnGawdby/Qw4Au8NAhG2dEGkeJvjt13u9cX8N/a5
K6gNCI6jx602hP9pVywdxccvY2pRP02hn7GW5bX2UYNzOdZY+0WEunPWZuS+snoK
VjSuYbtLf1wt8GLWFUCi4r0hZU61TW1HeqM5unxdJ6OZPW3Fb6aUEIP3Kv/6TKJc
OUMAM2aQoEo8Nkr4ITyUbcH0QjpJ4I6oXVOAyF6O6XvCRsA9SSFnqupKaLPxgpfp
W5PpS5LxrtTr3Pt8JyQyk5F9mgsb6zHZaKcm9JWXGqhQS6d99T8uombtdYgdYz+0
VMoctWVlxdmt9Zh13qvsFEH6967iIo+x9yHsuHs1OZTzTvhQw77iRjkhMEVURE8t
aObPG7Q0De7xnsZFcCP7XvSI8JXzWqpcRZFxceyXq1P8h3wwwXnXwLdlLBJVOIM6
ASSo3HzFV7zoPyppa7wwhj5FVk4aC4XqKkB2UdpGPAUYFhWTf8aBgo4kzyWvamam
VKtYzt1/YmTcnj08u14wk8IRh5peBaaOZWRvTmiMXoHGOCYXafAga/ysv4HNPhfn
YgegXEucPHKDbhCmnkv7gifMRgFiFz9zmXCoTzQUweqMtbeW0THxaCx+ucLBYx0P
RJBvfxfpPjtUrewlGy1xDvPG8TIxtn5ROELkogRxSrvGaneCOWFFMriDvRsI/I/T
fPxLaqbDVHBMUb9xmVIyHyi5rmPqcWtSDc75N+/U56rBLIj6fqF4R0i3ByLYw4mr
oyrb/SoJ98gLEm/BRteZ/7OERMN9c94+04lxNlWqoRmBUfnoNxcs8ExgONLzT8l0
sux0hzc6IYv437h7h6BNpxE5QS62XFK73VOQa7JRNTWOrMff7Lubawlg7pCjp1am
MA6KodHfHjJLABEyvDnqe9rzV24Z+WwwFF/nOSYEvhzMWYjPjsYYCTYi+wWYJyz+
dtgT2EIhATnfaVm1RWJfrJhXe5B0xqN9UV3w/wXm2FObo5bP/xrE7D80Y/2PoOL/
LeqSvQkH/gBzRzW2IoeJIw5Zv+4pvS5URKVVqcVkC/RalSwiMdERYPjZn+JNA5+5
EgnfnS9oBfN4x0RltoA/q1/X8L2sOZlM/0CV6S95S77dYmIs5xYv0DbMBCGNl2sE
FlYFbZCF4SensAxlIF9xHtyvi3MFQuFskRBD3WRqsBEbE7DqjsEwDi5ex1fXx9tS
McJbiWhGoJAwNMzJKcnPBDJ8ENnuwafO/cNvNpItppwsmqRp0j1xepZTLqZi698y
qPAgu5nrJNA4grXANvKp7JRrhNolvNnxakio5yAViBactUsYxBzxcVanFRKpHbO1
eFYyELdEq/fhmA2TRJz4NMospIcicnN7x7S8CsCyEUzHKZlyYiuo28PeinG62nSV
XEIklVfCV1WTfDEax/2Sieqv7BlKqx4XoobH1tH44+Ika9emZKQGXIbsXNwaVGkq
Ptyom4XaCjFKIoBRp2kftNeqhVwOAW3+pa7geQB/GFu+OQ9LXqNrGdO+emkjkYro
h2+SqK7hJaccwO4ukCcecxiZM9VNv79NVGDrqaPlM5ozxkiTCa2Rp9B4R2C4ICHa
hqFeRvpuGaw9WbRgBI4jWMgAqHD3HuxE2YwlEOU5rizTks0oKvr3Z+ajZhXhoba+
cuL3V4+2nRMs7Az1FX/Pqb2ie4gsjTSMcDk1ltf8GweQFUd176GF+cOm7cAW8BGz
b14DRWwlnuFQ1LUoehClQwS9uFalfldEQeq/I3UQ3x2P2AAPvScDkbvIa05Lxjci
cJM3uQwBioXFFnMOeEOYsILUwQEFfHVdblmLQeM7Q7T4g1yLNMku6bOhhkDH93we
r4dfyd8mQX16Ik1C2mg4asBgqMUeF3b0ocm26mrL/7EWH/w/r/hCzEfssyV54eiA
AnBS/caEaSdn+2sjyW9A2pC3ytTsR+GRoOBnmnxv4+xnYz8ohmqpM2zyUgAkzOLw
CozD1p6M9hvbU/1EI6/aRi8QTst5xakR9A5HqE+mmT4zR9nRsg70LgiWje9xVIS5
QIVnEYvQ33k8C/sowdVcneKzxdvHNnl7Hli152h27PHYNwHDOqKkHNHNjhZwsGAT
WbsWL0Zk+4OnSZo2sRZimW7Ouh0LES844YE9bW+Cjjnx3JhQJejgKj6/NFb4zRQr
z+01uH+lF4IpjWOczcQ1xxu56UQ9Nu6hK2wM/bnXPcYM6k8kZF1qeutGIKU0rCIR
4Y3xvfQ9aj0AS+m0y3PmBHcE+rRoeTtDc4TMpP+SAb3NvaxztblhL1Lqxv38+wQ5
cYdGS3EWZZPgfYwNOrpAq76+lY0hJOa/jP3G5/E+Nck8tUGx44apU377Ni2BhhCl
JBY0RoOv0qKJJGkjcKk8NpLlJRWtWDeE+82pUS7ExVN5DwlEWRZCaKofO5/OAjyw
THk8BV9rBDxTU+NSyz918wVvaQwKigGJ8Al5esNuJ5q1I8WRKlKdL2r6BMA/NK2d
ubp0TfqyNaudkARXoDIvr/I12III7gHCgzoITSnPNC/gksmqtp7TxWraIqJ9sYUq
AX9DQbQg1AAJsU3Y1esfF19MzN89Zkqp1vSj66myvca+ood48U31uyoWLngMsjqx
QT1dKNqbDEkk9Y9nLvtQmFqNOrDYcHaLeVGuPivss7tNRqr1QHo4cunZ/NgTWRx+
yMzpYsdlM0jcLaWdn7NPDTFBaqk7WnXYpRXSVd2bFu/K6AMAf6GFaFnFiN1I3wKE
kT1H8g+cdVCLFjNXkS51LdIkXNJUsMAgNRciD5yZJ7uqlaU3NwBDt/F5Bi6IXUVZ
jSKpumbqM+oHzCRrAC4jyr7Tswyif5bO4zp3Wx3UtRW/p6SlbyvnWdsGdUXtPNCb
IIx/FaUUWLoCz2D6dQb3DZSijVMmCIeH/N1miJ6Zu3J7Ks+7Wn4NTaTZaZcfDvG0
/RcAW5Uy8zyMTTDIhFMHQawKPTWh/QzyhCEmytBCDc+ak2k85bads1sOhHXznueT
zffJ2hVuazxkZ9yllteGZWeR7AsGOZJD1Asn3z+ZbkfJgjgZfgMPTskW7RukX6Ra
AdZ/c5k/rrmF4yEGxvTAhiRGH43eUSYfT6+5aYpV5TnDYcP2GgKsWxOuckt37ryO
gQYzg1zrm/lPelECP5Ar2P4CNTVAMERYhLssfBZj7pkkYk0JjwZi2utER1TLVS4P
U3QJofzyBaNaB+qAKy824rqgHUhm+RUfcomUXmnuTHgjsIHAmYjnvVcT+537XGfM
FRPdoW5kDxII2Tj7qhtER0tWpS2HtdMFA5BJcuW9kx1M8y6s16pvpc+Ubbo2Hbga
3TPxgqydKvC87RwpwRmXHdPD2y0VvqlVJO4befpTyrWc6fKYTv359KsPIsPP3KxQ
OOui7iqheWsMVykPpR4sql9Qii3NmhI2+057+mOx1aUGADeacYuK6sJO4MD1kFVV
3b/jgFvtJ3Ry4efWi80/y62FsDmxnmxPV40TXfGDvwzWdC428FLtFalrIFMTkwnN
vDkMlQbRDJ1lBBpZQF66WPkpAKKSd7LPmQh4/XDHelbh7MfXEIZuulcdLRGN793i
Z/GyUqotffFtd4nheK/2z9qt55U1YswvzZvDMm52PpzlwZoHYKjp1KB+tBuP+x0p
qzzfuFCZquZR138NpTAVkemDqSH2frPFNPJOqKoPI+CTdHRe00shW6s4KCYljzPU
L93YzSu9xIBAeDcUV6iyMA00b1z73Lx4pmWnDD621HOLaKDADxJHdSEIFI2ZQUiY
S/c0lf4DO4d4nx+ku9kdrDFGBz+Urk/3Hk3fzTDjXpjAaWV571TbpMm7E100pk5U
EEGkWMP5Il5pL4J0OOohqupcknrFE5I4rkGhNXYA/LnFujhg71dIOHhANIJiV65N
rAcmizVGHdpnOfYVQFi7lwpJeiRpQ0o6MlNCYr0QQIVonDYx0X3pmnbIIPHis6ma
bOTTYF6pPECo6l1imgP5zHyz0fcvqZe99g7W1uDsduzCG/cO/vX1aMdvTBTdbNg8
MWQhIaM6lTxobmsyDcVL6ChZR85Y2JDC+Zda+NtajyeHqXb8mFV1bX0zopKhyP4N
ES4gyFLcXoWfPqCb92Sug3gJZXfraqtkh3YME+W1iWX4yw6X+gRCwfDjVdXVnlpV
LQdz2pgU0Bv6PuJaqPmYRvPaAFkR8lh8HQPLohFADdSqYxPR9paJq26zDfNOBHY5
H8rY74QR5cfwhDH20a/3BGow2t/Bn32l1ZA3KstWUCN9K/aP8I4P1O1Z0IsGOgKR
17mSWSZPz+ZFTV9+c93u0jB8EI5qtZjvI2UKu9mdUI0FmwFAfypoQu3rlXvHzMNG
GbYSa2tb3ClqjO546BkiAoBR4ojNi3FdAtPZG+pzXhR6e4yBH8/hb6aAhDbISWNj
u5ymy1Nb365FydW0h73H5IHXukm+ztM3bJTiZIgX9msqqFYqumMsJucy515SQYtm
kQQzivderbm9H+Pz51HfDDXE2mKZ32hXaU8OrwELytQmtqvJhpaMcjse8ebqimaW
SVwazoD/Qv3LwqazSRfjR80lvR+y8VNcZblwuzv4bStH0W1+2qXGNJiJmPOJvFHA
0v8pAdHgsySS/aholobcVgz5hdDQ7q1KqGBiZV4PrFBKH/l7MxMT/B/vLNShdn6l
/rxO0Fjuqw6x599QdQXylCG1ueZ4G4liS5Gr54yXNmdMIdPKnRit9hnSXPZJYiOK
MFSuHRHy4f1UI+MubauIQp0ZVv4KmB7WWM0Kb+wPI6pYkWsn9sgYJ/P2Oa4HB4b3
9uS95efUsfasA09/M9rimcaBT/qzbGtVNgWwZgCngYEmydjb7tPfgB2fyPvRzIw8
ZO6nhTyk9PoiRm5tDOTraWn+nb5C2zMMaGQt5vNaWjP0cfzeMcspsLuW+EXZ/QsH
GEMuRCRCRtCtuRkhBv88kCIFgitVAodAl7aWBRKRaufe/y4cav+X+6dIU6VkbHgm
L+IHIpopY7Pi9G6niXQmeki9/gYVtbFV7AihhbmjskKeUyHBOEHPD3paqDgzcLDn
T7uDD4SlBNS6vaHgN7ZXCOqc2LhymnOGH7lrVbDzt8ZPEMsWY7qh5WV4q+R7Dujz
k+t4g7pH0Fn6bPovN5G+SSd5xwKA4rFuMB2pkbUI1CZaPvxVh/TIrW39Uwx2bn2M
o3vYYs7COUj2dnISdl1V2HVOFS+8sb4Hw5+NyJ/7hQHQC1W5tnIRlFkFnbqRPJ+A
wJu8spX6bh4Ut62ORnOocw5C2rh4mMPmStxQHC8zEztsjyWhLS1hDDsKwvuy/kRz
nP+p+tNf3gBkBKuQHjJ+ufJcv9sHxaC3zscHHTwP/047hNzfXYkoBNe4g+iLfUD0
tl3JuMda1cXGz8vwV3EoOgfY6dzp7fsSPYpvaiVY95GYX4A/R5gTylBbwZrijlLo
DTJjVGWQIIPA7yGdd87Tn0HQtzJ4wnLYZOxKls7gz5NLvhoaFUQDuTWuRNgfx/HY
req1mzKVVcgt3lIMMHJum/rCYPUsFfT9dLNe3IZqXepz8ASQxEnzwHsdxCmL8QeV
U2FZ0MvF2GF8r9sWtbEdOSxYhfUMZNWVill41/A/Xh7wLTViiDHZbQcLXdOjY4lU
bHc1hEsq2f5MNjMiw8Dm+aIdyNaijDJ7k0qNuX+9vsyeChPV1LJsr5F3cKYulZRN
ZApCFiQVTXOBHUar7IuBGkFuVq0qkqIwy29p7Eh9lB7pKFdliQzQZyf3mwB9YTSi
26Pljm3lkE7esf2EdLKamfjkfC5+Q7KY+MfUoQDO/RtnA5+X6I/PeGeHZHXHGBO8
y3Dd+3YQnSrOrWF9O0NibLB1X208NOAKg88GfbV+O5CKfdQ8U7ZC5iHbQCRMDf0v
dTk6gUdq7z1BQJCl1OzmwLBpKj3aEKRYCWsJJ/LOFyeq0JEFx10RcPgVwvAKDf+F
veW13ie/uj+C2dEnj2x2LQlCjjghvsyqKCMBU9LNgYTlSrcSJlqJYYB7pR/yFz1g
9RicDgo5RtFBWot0qh5ElNOYDSG+Je2/cynTsUx3c5xqutUHh3selNG7ckFj/ZVi
PuO2+NroA6LLR/rOHEty29GWMLbIIR5sQ3tYAD8ckR0r6kApwT6cRBtMjdeRsXND
GNZrF1iJOxuYm2e76ltXDfXy/PTRFgsxn7rRkTeW5KL0jgmB2Az7SHsVW0HhJFVW
fU9w6OcVKPq1QmxfVgUpwMwvvoLoJNQhHIUD30jzIij4sUdIkE6oK/oOOy8VIT/3
uP1IFmjqPoDrtPpJ9ePkRPiK1nRrMoOFJ86BwRa805ig2zUBw6ZQZMABIvONhgnC
r9oulXAvQWXVXv7b9g9fnwRJH7/KVMM1r9+xZbPPM4aVDij8Sjyn9ubGreCruRlG
OhKeH/nHZwRjuNzAlpwSR0LdsgtBa/IGmaTkb8qFbL+HEVrdxSQdGmD14yuoR4bT
JFfIaM8nwrYo4/UlQL+yMlJeOmfq/vmUKgz03y61DaH+5t56ttOcopXQP9Axmaoe
kPebFFssqC8zhN+LHDECs4lVXea3jV+SUYort6mBiNXnHcpd2GrE73GpJKPncNUf
uBsRXixxluc9/ZSX1rbwFhU9HXYQuKy+xu5XMyAd6As1IoX1lWJeELcsBm3S8BE0
SiFiOJA0IsYn96MkLBeC3Jm1iMRkrIR/rpInnPyygSEnmd2rNFcSt1mhbzpc+Dlx
cUjN5mckgmaRP2y60vPPO9nbSFJODspX4PxkmBfsrdwgLfPHrAT9KV3eeB118iQA
FGllx7nj2Ram9iV/vn8U9A==
`protect END_PROTECTED
