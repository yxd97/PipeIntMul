`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lmyghXaImLpjntV1dvbrYOtVGJ1bgMkIDSGMdSzq4BoalN5sJvptkYrLiPNvODZN
fY5EETccQr/h32u5hjtPnsAxwY/sO9SeF9fSHzORVmxn/3uzRQrD7i+Y0I55F1na
itm/p3cpvkSJyDj4eZe/6aiYzvS3zdMH9OuYrxYrjfnT6f+92BMoeVLVo77b0xPW
gZUWwVnMt8obO7metIq8i46b69mud6LtJDFCgwrPKOIJaKzZf8ksOoOwhbVeP71B
MRYK/UtKmSijTl5+dgYKPeM5nIMoqe3N/oYBpwB98f6xosrp0rqCjJQG291mQHJK
oMFi70BUZMRERe9B9jJwHOvk84FU3lZFjeJecCuRK4Q/zf7U2qC3cRlv1MqGqVxP
sZAaJN5rhG81WBHFKOabvkugsme0X/qmnPlWDtZSsB6ih7UKu3CcQ3Li6yzHMiD6
PABkUNVIXj0fW9gilo5LK41IfMyelQ7Y+kiffMobiZnxkOBzJEL5Vrv559JOBAQi
IjjfyBsbXNElUUYt2RlczftW0iIY5SPpzqH1b4RjdbjCjNw925aLuXy/i5LRY+TG
CmR7OSxM8idIT1INHd7oBA==
`protect END_PROTECTED
