`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I4DTQi+5EaXHyK120PTu1PCKEOzEs7jNdg+9EHcFkPF2LVc6o+6oiag9rrWkuA6L
aJp+j3QiZC44IVXPsOP0I+Ur54tiJHXiqj0wZ8A7iE005gLTHmhz0EEwqVbGTHvK
kcCzR8gsxZUHaOXyAqkxQGXh/9QHYoxnYJRCkWp4K5kOFv3hB0H5fUjndty/F7qI
Nhvg6dK9f7uu+8Z//duY0o5C68fwutzhDw/B3AkRSIqWNhO3AdcddP6WYRAalTiL
qiHBqq6d8UiFLMuli+c1kqyA+biJa7EB3fm4vXY7PakMTlWbZXlK8/TtNlgpqc6/
xuRa8p72JtCQJ4iePETvAAURB8t2MUE1Ng6i2RrMTd2khAPtBXM9NqSKPXTXSRVT
UMJNSeeik0Cqe4WXXe4er24TWaP2a20AIuRc/MCmry9VlRnC8mMSL98mh4w05Bb2
DB/0HToDM/YxyghaVB+7qAs2ULcYC9zWrjYsF87FB2yV1xBit9p8xrJF90bCh1NF
blqHts1VRZO18wSXNGsF57UHlmqm2sfgYjdrfM1EUfJDMccN9D7K6UC2ujEVfivu
SFwBgS5j31FxZQyOzXYC1C6Yb0Ltwwq/IOIeRnjBKOW8eBqfQovSL9tX4QZ40fpd
qEhmB6ySEct8gJkPgXdMuWDbDflnABScskB+jUtt+GJEE6s7ua1SrI229KGp473U
WmvCbBAwn3ma41LahxdGis9+XjVdttaAAHQFuIXsGtAQBvYQNhu1hhk9JMyRr8I+
3hMjgAn6QcXXABl4zB6Bf3cnXCmUeJIXxw/9lhcTHNmCubGI7rkdvOzWifViiNTG
jQ9SSGi6awtqqUdAiu1/TILtoljf6aW0axCVvSPW4TEpzQjUb9H4/hRbccTnu4N9
gYDJ2/x6jbn5GIYcuysasCvN4cWOo5JY2bDnez/rCAnal5q4UJMw8o6blH6MCwJ5
SAzZFH4fH0T+Ea8KI/p7+8pkbavtE4v6pl2s6b6Dmg2D/DGgVvlUcCM/S/+fyt1L
MvRcFyEtkpAniBSvoMtA1h61kVMDgzJ0Yk3u92j0ejskE7jhut9rZBxCuy7BCtdF
AQHioM2jiuo6/gDJUK77UAoFfQbOjkKN2DlumqRmeXZb7sG8eLRYFTc7aL8Jektt
sZK7mVleuM+oAPXcnmc0+651Pr9uwOPdm8+Q7QkpIl7P6ZGfMAkvhOQzIvWtBXTs
GKqWbcYsoEmArrYC/zEbPA==
`protect END_PROTECTED
