`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uRJfj2AUJwacKjVmxDBHzN+cVNnk3UnW5X3AamFaiFMJHyNXiaU6wy2YxgOGGklx
WfhNqYyPm3wkzvoP6KQ6dEiHmMaux20BvNCVKPGjX0amopRedYs2E0AIHTdkmdQa
7g8cTAku4wA/2mPYhdkq9OD+zo+Atrvv6z/Mw5rO4XYmhp/PaAjFqnbvA0BFlrtO
bpTg1rYY22Hgrta9aT4etRtqOzWJqlF7I0HT03CUAusZYZVqW7i4CG+gTju5uX4Y
SE5u5AouliyYuPesxLKJqaBLyYKwjr4dRWbKGRKqBsja+99TdB9E3B4daWYZeQpL
E2t37ZNhrrACMGXGiylo+0yNx74o8Nmrpdwo49qXBkL1ZJVEBPsqZJk6DTzPIlTU
HcJbraodk5SRC8pdhfmAAwaSAmeyKqI44JiaBWKf9SQl7Fnc+8IzgwWu9LD2gKNH
2HQ5CxRN7XJ4MgIEseDlhlfDbYG1+VKykKt20a2W33rJNPAEBBne4S1Pcg8D7/oy
yS6gWA34egLe3/1bT8TRpDn+7a5C9JPtmAtyhHpByyJ7UB6Kz+X2qeJcNG71Op2c
+OvxfkKtJYraJEWkx7ouSpM/8jY5gNHCwYGkXqecuwDKl6hxw5nUFMf3cFtSi0xL
Dg+GGKw0f13ZtQFcEjgwWi7D77EUq3QYZlzvVC+6GlM=
`protect END_PROTECTED
