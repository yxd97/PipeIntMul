`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TAyhUD9thYaVYBtXmKM2ZGx907tKFfaGkYgYNuyoA7WctT9Y4CnhRogwbqx1waWX
SLKOx1+kiPNzwyssQhX1fkzcYHgB+yfgP9F3MsGez0J0eBt4yv/8j/lFSN/awJDd
wSeQXXeyTMUpqXxBoKezNj7a8QquTyw8lRzsD5Hlp0J+iTeCb0179XqCHC67G9tD
CjiWWhYzh7p+WlFagAYW6fEkJDAKH/asS62CKT69ACMIaXRRKOQOw08m9BQqKvex
GUeSCzX3OoYGgX+oV1d1YPb7kLoUK2o5EIJ9L/fK7HMh4Mea3XTfHKBqZdydpKh7
Zcq3yErQkLjVCiUGkyFvt56543icJTw0/wH9ESgnoAlK4l0ShDOuQbbOlhiaWTxv
DFzwkvCfh2Qha6FpbkiUmUPVJGQcU5MOzBnBrVqLc2YIXcz0dFU1CNSt4EpP7N/u
XjJmU/3m7LGpyICqjCdHaYmVU6+etK0Kqw8taJEHu82h1c6I5eApB50LvnVe/8Mg
`protect END_PROTECTED
