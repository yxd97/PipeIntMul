`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zOxqfHaHaJyMqFg1hJdb/LqqR3HBnDPg1jm+pVb8qzGSSwyIuB6XfYFalf/ZBoN
uWtdQP7ryOCYXKesN5tySqyHM6UoedC1UmvekxvTcouLsCucxm+kEdr/NnExiXWx
a75ASO125pxrkPlqkkesoiGuBi6Wyuc2vtBT+EIqbmHwwNSU5xoYc70dBJTajLWE
FH24bVBWjQw3YJ+8PbLX7unLxjkq1ae2GHmeDQzpJClAbWBcK87kkxP9MkskXtPt
DPUnsgq1m/MnfsvoWVkpKAcy1YQjs5OQKWY1WRnK2kU1PKAOIVdfK6ngSs8c4ha4
DVWrpHyC48JyPoAvxKwS+ex3SOxfEPVAu5lSppVS0RsjofKxXmvHbyxeVzzdRcwf
enTYShcdTjdMxrqhspreHg==
`protect END_PROTECTED
