`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mex1xYFcCgM2WGwt2W5dfmLYQhm/vTpao61/wL7Fk7hQhZ8b7FMHSHNK14jk+MQv
0n6MHKFoOXMmHuugC+dcDLGl9g6bpaBS34x+a4UMyxiYllZuE4RRb1tSPVNQ6F47
rS8xT8bnP1OLPunbcGbemDhFyMiKV6Qu+IHHivWybX4NBxCdg1t3Rt+s7K9daaLF
PdPfqLlp0+9nakfI0QF5QHUeyYWqPCk5xyYFezF7L2iSdrnTJC81GyhUCgGEHtBq
fnkO+IoaUGSbX2U0nFKt9Jyu4kPxPNxEheC9hPS8X25EwHToJMb1jvvtHLC87gMj
m9T8SkdlMMVg/aDV8sNgOzXqhXMe592VsBrYE75lrVFuIfDesoZC+Vfi+1dA98yk
W0wN1UTrB/weM32PlbTZaA==
`protect END_PROTECTED
