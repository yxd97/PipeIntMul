`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQia1q4MeGshJvM5WkKRCWR83CkSn/SW3bkoagYLDUWK5atbGT6xOXukP4DIl+9m
ldvr7YstCqUwI3fzdwfbXCc65JyAwBYxJkOHWKythgNdENcrkoUx4XX957+Go1wd
/VUo13YBOnkNGQNacRC8CQBNDtaLmJU+HCaDi53MSnN3ubpA2JbvYa8U+E/s1F2q
SGpILot+XKla1xCENvCBtFaVKZz8FCU0fYsVuzMTNOpkx6xxLJkVUzhNWPge5T6r
yO4qFjGPkpgEpIBCKgmncLtqYeSlyMqDUbdeZs14lzl1tFP5i22aXdDfdNWMWkd5
+aNtHG3sFMsDzMABjZUoJQ==
`protect END_PROTECTED
