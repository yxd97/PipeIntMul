`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cduZJKxNcLG2hjB41m/s2/D4q4AiSkky8ZRZ3VprVEbYmuuBaCgK6eWs5EaFI5wP
xyqTa924VB0vJtczOXxcs4Q8fNu9+WgZNaNr+ji/2Tr/Qo3hEKHMQqY4mJMjbhET
JQvycJjerlKym4MvCcM9WFJ+bVXjUMbbcU52mOn/8odAzU9MTQn2oYcz5pLBAAp9
5BFX7Pb8fXb6uWTXG9RrHvF4W4uXIZL78s2JOP1lvP6cZMIDyC0AX3k2n+iGFW87
KUlsQ0IVzWXs7t+DdKeqXNI44rSkR+cdOEYLryDVIriipgodciECX/K26nu0fkRg
W3CHEDHwReHIeBhL7WagxiNlQBIKthNljtdrxEYlS3VuTU8iSVJ4/YN+kwPdoLLL
82PeknE/PiLo/UZNt2EFuLPvOWArstUCiZXWsBJkHihQC0D2mEprOJcPO+kz78n+
fwE/5h//M/Yr6Lh9kniUEzcDWMqcMVOWs0SCdLq6vzk=
`protect END_PROTECTED
