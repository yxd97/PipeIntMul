`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bezJ8lesyPAzSv2w3NsmNTGeXVYlEvi1Ct07WVVpsVv3zZz1qOMEQOHKtHAMFzyC
1Z0TEAy4RVrZivpGu5aZlLpACVvvcyVCc+SCPg/ZOQweRBDtSBCex9f+aHh4N7Pi
OyTjLqnmOkiOHWcM37tBHZ4RGAtOd1fMYF6DcGWG0OX5GdxDn6DbSkTUzoeElCGK
Kd1Y+rGU21b5haegKoaKCG8cN7o98zkjiwQvWTZPNPoFswM+lW8pd/DshFWiu2UY
X7j6rVNVZE/kRji2XESc+/PlLSOCorqjKUA8Xvc+RYlhPMsH0++VlkGdr27O+vz4
ROszgbe2kI/8t4wODtv/osUyOUhiihnZ6/dPbnAKgRYRnji6S+wQDHZobWQEizHO
y5HbxXOzj+Q8iFf3YcB4cPv597K4SmfSsnY7WIZnK8JXFyBycG4eOlCfp46a7ILc
l5prtg13DEW5CmICE34SotpHHn+3yCNJAJRMnrgotMna2KZhZVGNCUGw/qK5mSfr
g4yWEWUA+kfeUEtNVY7+xkGfasiw3oYBAfHtvG2d14r4hln+NlE0BU9oVgy6FgNd
nYZ6rn6M+ArKmSGThq63Z8tKz+6AFymWq8TjCsF46ZP1k4AWahStexHCNusIrjX7
TpUMhLi+njEKZuwxxhLydVQ0exYqLwHKOVHv3ml85mNK78AoO2HDVDpUqSAVsgoe
p/b1YVEa9alwAUb+ehsaK28ehCNiDi/LuFc4SKIEhAmMKsL48xxe7zBMpj48g9gR
8NEUEYDiuG0I1ObVOB7+/VqYy5bkt4MIpqOQxeoNl10SgIeV37G9/257btS6AQIu
53h5kth4Oj1wz7uxsuobW/ZJsQtnnTWKVpxg+wGfzbURE+Okf0KswKUMj2v5MKXS
NSDusUdkv/+vtG2/loI85KWIWqWbSwdtVgIqcDKbibSAAC0QP5ot+HiTcv3DbJUt
oGn3K1A9UCb/DZXLqsKkVUjYA4a7Aer8F9NvSD/WqbWp8kaZUXcrTaY+i42jpnth
3R7I7ImxpnoUAQWTqw/njOVGuFtVUeCRYL+borNSU7qxuBPr+hxiK2zmX94CBGZ7
3Bmd4To4IGNsEwp6HdC0ZxuNm/doGAsnfQSVkQK8XAR1JHsTc+GxiG1/LpyQF+sy
`protect END_PROTECTED
