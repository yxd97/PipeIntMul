`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kkl7iFAWrE7g6xp/27kIlg6G4h74w75gbLdzUkN0bv993oZJ1QtMTnaOtZ0N/+A4
CHmiX8kS26GFZ1eJZvFa6fzGqlu1GCFOURMQPnZp9xuVRpopR5JRLUgGArZ/drjF
CRgZQSeRO2KxMoEMmOmzL9qNXX+hIM1O+awa2/NICb1cTKkGT2n1MRYAZbqh3zF9
QdMH9R96Wcvs0UsvN+Qw/G8kn/9uYwk2LcZELfF6W4qsLiLWqCXTYg87w9ZNwvwI
we/deeivwS7iHkqYYTMRbRfGJXLdf88Q84m9H6ELo8R3L/DSQqC7Kg934ujhfMA/
eIM9lsD9k5ageoqZ9TqG5r3kWWTU9hHhf0kJxb4fkXXhtFk2LYYpLsEgKcn9rc41
jpzSaP1aHf1cB0HzmGe/GvhCl+BKXGa/EzGqJtVssCQG5YK+GGbEqdpJAtsKFHQ7
RQfL8kLE58g+B0O3TUX6aoaqCBy9aQO/IQM/sKjWWY91j+7Iv8flMIt+WU/kgr7T
Ftu3efrDLQHAoQyr6ErwA4dLrt7ki6VhhWEYp4oRpPKT/akWTK+YC+WmNVTIx4mh
HALr3VetZgDvf2V2AMOCsIk0J9jk3OIagO2031o77lh1MTNUbOiH/fAlNOZL/Jkv
r3SCcoP/orjHPTTBGfD5zg==
`protect END_PROTECTED
