`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LpWAsjeLRLy7D3Pz1FhipMlT5x7Sr+gZBXd/NPPaTGXGpa9pmd3Yr/bi7FVwoibZ
9KsseJeUAEqR7F7IHzgCBiQkVYSsFRXxDudJ3qnw3GHiETMPDELKdOCnWMVl+Cgu
SvGVcwf1Aucu13tUX8DfW5kky1eFXFBj01hLdkqTDrcYHMQtq3kL51p1RYpmS5YT
XkbtTkQHbvJSRsT0OGnVZFBWvzShzHzP7KbOujVt1ztcn+1wEvil1tvQrEbY3O/O
tlGWP+TilqxRdRFsPPrcaINYX0OMoIMmltpmj74y9+QUtbbdXzsIv34hIu7ElQOn
Y9NU+mWi9fIiOGnL2X/kn6cGpaKPq30wAKWim4AdW9k1eaxGtNpWPK2vyBOYzR0k
Z6qUVeNxNaOrpO7UdQd8ieLmfcP7XO9GXY3U+ToAPvwXHuJEtAIo7HHIwoiB/TbK
VjoLsf0M4w0nF7zX8me2ePn0gbLshetxd21+i/NmAYiVxWJ4EaD50ZH/3vbUqS0N
7CDMhd18jzIr+h4tGCD08JNAsF3H1BBNnBXsSQnWdyIVxUPKaWFKyXIzkgZ03s/R
///ENCa4zqtq9vgvyAco+5eOfpMnyLQmwab6SqAuFxil19OOwI6C6hqRGxQzYwjF
H1LOdXc0kqQ/nNOA15Tm6pF3ItT+Qf1jS1PPLbo9J8CGuQblzQyBxULRTgfoFnxw
u42VgVh9kXQrc1uPq6Kkh1vchm9k3uiqsFVxMzBNFDycISaAiBMZSjJ8cl3JOL6W
t/VX5EL027svuKI1nmEEhp/DtJauTNElJ7HDixzI7pw8suvHQkedDzIlciYHxUZ9
AX+gw150T3sDPtObflQnJk+pZmGuHVUm1fQ2aHC3xdOh4dEtaWh1ajwTcqox7CoE
EXdJtepd9/0cRkgG+1h/ninDjDiZTJD+cG4r/hy7oPgQnFD/Sar4rF8Q78J85ulO
pSL06+5hv8Gbx98KCWfZY/cE7waJ5GNE9OgdtHP4EpOh9dTJhU25tUIdcOCvt1Q1
gmMBR88+tqprPKJD4Q+PNOXqwvEFeexLiONTT+Lmnk/gaDtzfZmVkEy2r7S00giK
QI5T/jtVykh5tu7jVQ8sCcNJEgoi5PUnd9/HP2PcWrANtxtM9KxY7HMK/aZUSde8
`protect END_PROTECTED
