`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8q3WZzuRuWihUZAedGEghaYRt1IfF93P44piiEeF2cwjdxSmyUETYWV+XLexeQH
bYcDbbIqD3IjXbi2ZWUETfvny77iDnRetUGmpZM3KVHZAJaN9xdGucRlX/jHLpsF
Zl1BTPs7UEFeXMGnzLuWqAKtNiPnXP+8RF/1IoUPADmOf6MIAP6RvBWuGLlR/9tI
WCruWUmdeJ0Gj139ZwQed4FjNiCz78/hMgVD+m4K2EHLFf3biHTOgh6CdAvkxm0z
FNV8s5UKNHUkah66LjESNY9SSBeOoEvC5E+IoAkUSmFdr2mRboNy+nNVByCSFbjw
PXKxCTrekkVvPrgvDSq3zI/tnyEPRG0z62/NAeJi9LmmwV/Mxr5/s0wxL48kjOvV
6Z2eC7ZuURQ5+5c+YU50/gItGsPeZHYlgRazzWLB1oWjQNNiQYK+rhHQAg04R2Af
mWvTw058YNU0rVZ7XBmOhuzeWvVGSuQr3gdQIvI9sJ0=
`protect END_PROTECTED
