`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L+qhVIuv+pi3vNiyFZQ84R1hC5p8XnYvcn9OQGwyDXtaByNbisFTBql/f6c97ccJ
K4wzEvkGNieqv1HZHt/d+i/RANOZQWQ4Ju+XKfMZneikU5ZQa4/66BV8YXKo3EaV
sTj9iwsFT2EMFzdm28qH2s86WW540kbRKqevVr5J/KFDgW5lm64XNoBdTimGTRZv
gcYWWTGxhCV4aEMCfxv7VCVYj/rAeIT3ZxA7HLJ7wyeFFwVYYTgTE+3wnnhD0uXo
fpLysarHhILhE+VWW/9ZY0bPRPhMNpEQJpGKR9Xf30Y6KnsY3OXy5vFzC1OqUBcn
AlaxJ8OvauAlQ8zR2uyHMXGJkKeje9hkp606d0PZSFyjjBYYPbaG1tvci52lg+RF
9E7NahBqlhTHSJrCcQOqCdblhOopVQXrmVhc8H8GbIsFl5MPCv/ec17MlXqk8XOW
Dc8iWCQ6uMc/V8f1woXTRx5nnVkD2iBPqaKfuqZp7vDMc0qhSz/5ap48+IfXHwNw
Eof+U8jYEc/riW2LqlpH6Bw/TD+N/SQg6s/+QjJb0EuykF2YvtGs3bgeRVinEROu
bED6N8tCc4HFIjpcF6M8IfsK+Lyn1YshllBuFUuzlE6s5pXXCefiCvYhgg9FfXvJ
M7rGXGagCKQMnFmNvQ6Wc5FRuR6R/Y7FwNV+Jc/N8LXI2DtzqyIkN4hJyeFMLLc2
LbSjhOO8vkGIsPepEn9wUNiF+zKCMvm330QzVfJfh+nGKN74jWygcGwPn7Ml0DT/
dhB3GAS38CHGARHSioLZj/1nq8TUfrJUm6fLK+ViphSM0pP3UI10Zg+1hsQqagJb
Fg4yYHp/oxfWDlz5rWDG91tJLpkrXSAG9g5kAxBLZ7tWp5UMbLnYLp5M653d4f89
oUBIKekRNHasQTbblKQ26xVdMpsZwuTbsoe2wQkeqgP01QYnMBDbMSki+aY4ncSY
`protect END_PROTECTED
