`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jyjcGpUqbwYJBmCd0knBf+JqXCQeW4yUF6+ymktC+2enfPvzD31AZUHuGD4uDWOS
tXtTb/2JDhUB1EZngSQ6gpQd0bEOpMoRzhkbZMWhYmplv4kV57+f7km4sXURjw7u
3CEdiiMifSNmuUpJbL0gxwM4fB15HAU5fiNZ84RAsjtH4YEmnAB8vZoIri4SnsV8
jY1LHDjqYsjr7IC/FBMrjcxWAsrk4/zhr/KyjvOqaSh708y1eT4rTPYfTccogEje
JCRYqDs9oX1x1NitfVBdEIu8yUESZHRlSaF4tmCAG67ZobelVvnLuMK2vjBjfCx0
0Ohdg5sJsZSFjd8bdC136EMSIR94DzQ/9UUE9e+psSyDz3eIcg07UIvUO4zO0OEU
QZ5Hz2aOh753dErYeT2SdCvDuuivwXgGYuklYqyVPNspCr1xOWPXbEYtXlHCeYc6
CuxoqV/DIQaFD/9AfxNGNDRBaxVa0HhStfb/UUoSX4ORABUfvDuiMLzpyB2VlkPj
a1Lj+LLlfgK4aTVLv41PaAxhvC0OuoK7ITgfAM6VMAoxnpmsQ2jIc+QtS5zXLRj+
sErm0JiVClT33OwvrfO3PMIv0h5wXHbN0HbH7NY2ChP3X2U7loJMDhS06Bu5kCle
eHwn4yvoI6Q5lc83IdXb8vKcbMjNAR9qDyNFBjoiUW/LrusTCotjWKxY9xVxRgL5
toS4WidIS0TUxVsaZeo8Q12nHtAPVtzgnIoiNynD0y7ExkdTMfQ42DO6yLCiqKNk
lHAzfPO/Xp4S8hFj1hDHhwHMrG7VKGqha2437TzD80S7Qd1k1W8lxx+S5dEaESan
B4VpVz4W4ZLE/yZWEWqHKro/o8YGKQJOa0h7zj1ZuSQB1ysNGalqGsqn7msy2AnM
JdpuWyp/FZFYFKzBL6qNvgls2TT9ILAMfZMTAd/lzEopZyMO+ECCvPzNvcN0j8Wj
zVy86ZTnTkUWwXd2jCUbXxZLkRsLOMkr1nA//E9IH6ODpUXVi94MsVI1QyiI0LAH
E/ZQlH/NfNW78HhbSSsMtMxCfTvVGQc9qQicRNDIKRUl/0WXnDymJDTo6HgjxqY8
zZI6ZHLU3TtXe5tBFNCCCanlso/nspYClhXF77q++v763SOPmtyWoANoeEnvJkXA
6gDOffN3W5Nm/k1MXieyVGGT9jHQvcjjR78Rr5OkcZCidNFQ66wFAmeUTkgJ3KSi
`protect END_PROTECTED
