`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UWRV9D8gbNoJwFvLmbSYYqWTezZpa7nWJe1cLFfvQrKapbVvCsAb+WuKnrTNegBm
hsNmxCJt85ZEdPQWGhdh+ZkWB1zrL7PVHawahyTnA74rifVCODkYQj2BCXylNziw
aisKV18EE48oqDRGAxU3WuEN+bBIDaeWHVrBJaAWnOMPIYczCtO1+SJN+sBUTJHv
3Yrc6YSMq2xlwiY+bQi6efss9yF8BlCfYBkiovqewLhzZXBQoLQFWHSjPLOufCXd
p6qudh4m6c0ZFLh7cMcxupCdDzrwxrJcnB9Yw9jpe+A3QZeMTmH/obl/xWpXKEbQ
iLZ7mHHovW6HAoTlYczjEiTCbV9nJHgtgKJZ+au6Dz9N+b3LFFDEaZTP2VTYyiaC
KDhCSYIjMEc3dPdKmhv9gHCXG4I4ZJBQH9GKA4I4V0Gc2TQNIwd89wbue1/0ljsk
eqlf/wnJ7pxnDnqs5RKAy15BKkdu8I+0rAo9D8vfDTiKhYkVHimbLYkDA7gqUPTu
RpTPBqytCDwjhZaEnKy1lnZPKbZ//Rt4zH9Ep3rz1Vx/PiWX76JM4VY9/Xp2Dmzk
bkKvVj1PUOE8DbMMmkWq0EXTOFh6bjAZztiH7geJV1URf0VQsXgZjJDUmQl/+7xF
KLD38dxlP+QhXZj3hzoZ1/xdCfd9d5MydBSgNKYTyavtX6E3ucE0DSoV54/O0Ctp
`protect END_PROTECTED
