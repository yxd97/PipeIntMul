`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLrnNA4MSNXz0ykDRJFViicxMDA4PouHXQtDMHxkJn6YB3yI6zBxDONzzcI9/WAd
T2koCCH7XG2+4z+7ngXW6iRKSsB/m3nAjs+vU79/ix6EquSDwPHwICnhKEE83qIL
5EIAtkGT3i30WqYWMmAV8t91Z1LcLbNQNiZIijkXNcO4aDW2nvYf0Ofqn37sxklw
Dn7Tw46+axo/slRF9xR8eWgIWEYMnuP8l9gkRhjGNrFUtqz37S982xPHvbAp3nbS
Se8DTNPvfW2pYtOIAHg3ze0yWrt9RWf4O57oLHRWno3hBcCZCzfoXtljzHtC5rqt
TRU66NaCk9RUW0x+uNg0xnrIGLql3s/6zHyILEAWp6MmLnDoSXXgiRCSMXnhNkJ8
olmeZ/KBWGNI0EbL5XdofdgbCL0PEFlARy3cITydd6gYky6hR0qKLKIwB9rYEbgF
anGmE3bg/zg1nX2K8ZGGvPDMB/2GsKgPg9cMv6GWT5K1hVKD6foiF0shUBJIKqta
AOpiHiEFZ7PZ23fJxAIfA/GJ4hogr7fzZTECxT4LfstO2X9moG6+FvRbDjmdrth8
/CVJyxzoZfS9PLlp/CtiGW1QSX6kBEo2BnuYleZC6C4=
`protect END_PROTECTED
