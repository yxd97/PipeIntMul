`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEqgUeF5w+wKLpZeqxQUa36SvtfosVKfRDe9Ynv0b4VqB8arUPB7gwo4NbaJ5TEE
OS8VJn0w+eO1TuqUUDR6fJHfJFFbFVje0nj+idSSpt9Lih8Bi3nqJGi9P96tZmVf
I2QQqLsRWzqasg8BSz8Pp7s7boBtO0+wetGrcRQzy115ZKuSvTzoZ39AKZE/SYwC
DN+KGGOpYwmZCyPYwJMwhd8IvlUIaFo5vzofu7UTK8DdPkHiR9v14HwuM7z8x9SZ
BzrM9kS/7h4+P9YBoBL5WVDpEw+IEgEjS9WaObkgReuGODCrgBlPcpaU3xcI+f1M
xQG+bVXyPzv20fnkb+AlBaOz9UmyaLyp/bBogIUx708njZLhiKA8+l51dHQR3jM7
bpJM7ERNbw9aZHBxeRo/kDliJe8SsS8QIEVrjDkj+3kOgOFfdpwpCGzeyK1yNbPu
oS5yM61Vamqnu5ESDcAnZteAIm/waBAlf6hhEzGvkDd+kaK0tgFEmkWVhRCHMHjW
`protect END_PROTECTED
