`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQ7bIE6uzLPXcXHah7Dyv5+G6F0iwfV+PQPUhgAi/FzfT2qEITV0x/uZJZc4jF8/
rNWHc559B5LUGg79cgd/x4m4Wy2CCrYVt2qKE4TaTynN8/vAy3vBLiQ9EDCrODDt
ciG4SXoinBTbQaGblSaWF/Ivq17osJ7EwV7uNWrnjh2DTukC/OeG7vnPC2k5Xfxw
1dvjhWQf8zpEQj0L9ycPndnC9GGdtoKT+CBQUNJtscJYFqgFEPvxzd7X8XoWP89r
nRFEOXqxMjnrekXAtFKrdpXs9hW/H2IqXHA9llora9dSAHAFEUPiX0wFkbWliOVR
TzBnJHhZ4rXS5jnP4KhjOsZwYkpTcNjEChs8i8lKTQHAkupb4aoXxTl4bnrVv48B
b1V2kmD7GhqKYCACroD5EPBTtkuAmIJKt47bk3XEaQtr/xf5Xoc3Mxi33wFZvdRf
SBsTe/f4MC+3Ld8q3kA8TrU+D8laagyTAI+C+QW79GhlBf7pRkxrnwB7gCKPJbkq
L9E6X/FDjPkFrpw3Yj90+mvQRhzBsA5seJJ2ksH3Hdo44hJprJzW27EM9UP2T9pZ
cyQuARWrJD1A8pJkdfDCEsSktRMbx8PBH+wJNOAzx446AluFVcsLyR9fNi8NeKSJ
YdlyGDTX5aAmf0KtOy73Q/wKGGf/KzUq2OldKlwYGDf9rukg5dTIcDx4lHKA+nPK
ybS7RYyaoCJk7goFOV8FG77h0LbYvvHIoPxLXIZVm9OutbIorNH0gavAPmwzLY8k
+ZOsH4+ctoPRwPK64HQtOHA8u3oG5TN2qKn1Tbc5H3pA9ILxB3OtdlPmyavQH8hJ
0nH+Z0rN23jh2yxei/SROtIXwoxtxTNH2avqXjsX92P4BhPFduwaVzGrYSntGDho
Yu6Mp3oA9RCESt3jhOJjBknjVPWsiJH2ELCER1lfgy5WbE1GFvh1hCCTvojPJZIO
VpXD+ttl0Me7bxL/h/YJhfN3egTwRu1Wyz6qf92BzXOCpHY8BeLHx3IyHM/rlNjp
kV48+vbg55EftwpKTlB64aG3iDhm0kJRoenxtOlfWcw8jJhnGu0m/IiQM+oa6fIe
uciocz6UtGGM8STKh4FqmTEDbyoFjlsN8KCkMne3kua4Z3eaYrp6Ja1+3oaRKhtq
WhIAy7zwIJjbVxcIW+8J4ujvLkiaQSEwyuaHoYf8yrQ=
`protect END_PROTECTED
