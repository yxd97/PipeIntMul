`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T/kTzAO3oGfdsvFtJXZ/c5W7zq13cdmyP26zPr1cEjY7k2pktIc0Ur+krmDD/8NQ
SHKdtvw2PsTK1PK/GxMUD1c72UWtJqPmMrq79W7+Cl7Z9Gd0PcKD33fVJfdb3t/U
2WxA3oAoWcxvW55jy6SF8i9dF2l6yxnfPVqkfUw4U2yy+nnF0c1TV/wT6tegFZNP
x8xg5ltyqoTWAQmLfg9jTB+2XrBdK49W43zR5lZ2W6CmCZm853S7R6yix0/DuD6o
dfjVxl9Rb5xB5+Gb7qzVRFeD6w3/2ja7rPux829zlcMkOCTLrZKNdxO77ALSzw0t
mO+2Ag5KF4LSeVMlXeoVFU559upG9FbAmHp7FpTejLmg2Kw+/4Tn8czD3PxhMQFS
ILRqFzQ6os9aSpWbJPkMbvnaQ1jn/wI807yp5XugT5c8SpYtZ5VryHT2ZzpT4zPk
J1pTtqwKBlDIRkXo6qczPSZzx8Bv8Shl+06Hsw9lqkKwzLK5gTSbNnJUzQlcMt4Y
TIm/+LlXzbQ6UYVvyGorpIU+WbjEoLk6lIqQMqosR1yG5zlPS2enslIkbC7Ii9QV
zpz/8+4rBwhV0bWqALwKV3r4hqN3rRfx1zCMfz92pYik2FH24vL3x/CM1i/YBylq
P+zfIetp+MsRcRKmlkP+jkUMS1JUDv5KXBRpAjGz84op6pW5+fbCWIrSnS/YnV1U
YIR9tqYB9pWH42pHSQY3Q16R1VXIaPUZAwCX2dcKJ0V0Ahsadi7TAxVv+ux/Mes0
WTcupD3OUfIlujmQPth8GNfngczN11vMWv64FgTHrL8=
`protect END_PROTECTED
