`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pcfaQzcrdC8R6wCoDG0HgDr1mr82RdEXcc1rzFXUZuYWSy1+n1JAiBGM8aedkEWE
A4AM7d/xcKXRtAk6voEMPHO7Ps1biDzCTPUy3vh+xYjvivLhHKKTURXYa7A5Z7ci
te2djX4Hts6XgaXYSxik+bnTOr6ULqGFETVLc8UvasaUvrKFACpz7DS+WVKDI/d7
OYte7L/ZUJq/D+wy9bFRDxEfYnJodNKgrV/dBVjs1VqoveRLp4O/D9gsAuyzThsa
DnZ4XJMVsKO6puo4FfWHDJU2MnMJF7usIRi4e1HZF+WzKsR+3WnsAEF7aNJJcZYY
/AQefMbBHiIGcnUSebHNn6jbzll0wsYa9TVIGoQ+GsLbwZulEnEf1MrtBzyK67zm
8UMbXkKK6I5/eAZYrn1ox8zxbRQrdq0kByIVzngbjIeALhZD8gdjQsdCTmXUpiu9
ygC6hau7JcOnAKEt7U0+dBA8r0yOV7bXOD4SICDRxwt03yA+enfv+qM32nFQ0e2l
b1KKuAfsjzsmKNMorMsDiYRRImoTqkSYUqUVJKsKr6FHwu8q3yyRSSEgpEV7hm9n
v2WZgZOqSVXlrE9Idqf6/uGDe0ziRQ5NzWeENr/ELtv3u23A8F6YPLolisCQ4S4S
fd4mwUsTLgL+Diy3y9fsqo06y3E/5iXAzO/wgrA+5mAcObdLTRCwup8rgYQ8d6sc
Mi7gmXfxTeQlijDo85PMVpQSoK+5wc+1BP7AsuZH6i0AttwpFR6Pi/EwzvQ3/tj0
ZLRohPxCP4aZTOO/1dG0xVonoZfOsmBRBtYubiHRNMEzkmsNitW4/vJwlXi7L1nP
hcY64S3pQ5GRxfH/aRCAM/nsFP8+bOm3jzXoGI49lVN7UKmS8GRzk3VtNQD1KizA
QXRpp0/oNDK5zt7z4RyCkMapbnOhK2HRypGA6IxvRhNQ80EeWlF3t3KAlTNRvOkJ
ILtNrtP+BNc7RtEw6wSKf9p+0/px+ay0i9bMabdjI6Ged6LXoR7BDDQSw5G2PsBt
E8A9nr8lyzLroRpz6PkDWlkPtkE83dSw6pjHibh6BXGb2x+j0TW9MBHyftb0JCWg
Abx+vPaDp7mXc9R6SvZQkSMs4aqP3XNER/c5rLzOubiQbYKoGceuWKD8ogSYJS4b
`protect END_PROTECTED
