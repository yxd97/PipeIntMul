`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xoMTKPI0SpuRDJhYaV8Hhpq/RWnVD4kcl0jrQMLy0Nj3rsNSCKWI97cwg4G3+gk
06La2UqwyPetS4+pqfgYDZ292uD11Tsa8xMIAQZQJ6md0nWMDCU/J0E7wyuRfLPE
ZHIH2LsMajGOHtQtFDdk92LWpEPVwLMsiUmRcx+MKgrco+n/JoiopXOV3YgZQ0DY
MdMPWWbjNrvm7igOvP8el36lpjSxslYb0tiVhqdnG2vXjzeGcWkm92Z91bOUZgW/
WT5EUxtg2F2OgvzxoZPjV2xTa4XOdh5gMxiYC60tthCyV/WgDQPTfyd17Jcc7Rf4
T+9qMMbUaRDrbGvp9aiz0XWnPeeNmIzwf9b2tmOIIkqljjSvOxbGF0ZnuzW+Wsgd
drPIuYlEENRkWXc+Glcq+yqu/WAmvvN5JPSR063TRR/XVXlCXOX1cFBzl4EwaaoV
3XG6eMblJ+QkGgei+YnV7g9nzjEXKdCh6e2YQ8bhW3R0iYUD8PUsMvpzL2yxh3oV
Ftxwl1/J1lIbx4wzLrz+h4nLtVpvDrHFe15lkibXjZN/l6ZQS8VqgY63Q694cL15
6rBjEHVEPQd6KaKVXc/DmNLTAMToED1ZIbzl4fzeeineV8yh36i7JKVeqa+eZFfh
PwLYzaCpVxBrFQ56OBTRMx97JHFsfM8hmgxexUvQs8HGKMw4zI3X1phIMem/t0BA
9tlWREBvxcK/PGF4ESGnOrvZs5zykhZFuWVAEYE/1fGofttrOQtqq33ObC9Q2CVY
ul7hMzJjLxcyXB6EZUJITzzedxc6MwlUM2Bzz9zbFQcd89qg9nWgMt0OiNwjRbMa
zdk3zmKbQGhLbYcgEpPUPqD46po2CkMoA2rSqH0qISxzmvI7Eit6QZBjcYnBAEs2
6ZbTs5ZGDPjAjNb4G24ettox1Pow7H/ScUWf1y8BduywvMCtQZrNgHa3QQ3eWOXR
/BGfNwmkuXPIO9ZjjvpiMQ==
`protect END_PROTECTED
