`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
neNyQbia9Ygb4YDvRfE69wSPCuGtPm54YDr/t8djxmNN/8i7inhGypedb/b1tc77
iAR+6bflRR8275HDCyGE9/9xdnh6E15tbz0wqF6aT+c/KSi9uE0XtCBfglUciKpP
VEtpLZkoa97cfo56sbzi51ORH2XZiz8TWSg/PdweAcb++kqVIj9Dpk4hbwAV4aKG
IYHZSc5ndWxVuK5cbsyJqqX4L6uVyMl0n8IRbENfSR9M3msTnhny+Ty87rmWcow6
Ei8s86XZwRN9L36KsIz/IOrd3C+VLZKNjNNxxv929oT66JE6SlEecIw0B3gl3DLj
Dn2w8CVJ0bpt0knxz/8SSghMmunlK1QnHP+hwv+2r5ZJJ6Xm1UK+XlFtlcNeR789
o5lNaAXNhASCfqI1D0gWvZ2PoPY1fOI/BIcanN3D+GD3yVXpOh38crbw0Fmdt0lH
7nOfklJ85scon1iXc61byaPStJlpJCUoX1v6mBWCCI3+Ro/pGrQipMLtq2dMSrjw
tMV375RSST2qupUySONTCOnn/I8W+ycxkqghzS8zCt3G4jng8MN2n0qU0pB54pFD
ujTWzKN/zOEXTepbjIGxQQe8wHVqVEJeZgelE2x97dWgAlyPMKjbGJS4TeZkYUuv
tgp77lISRmGE/oGm/YTXcG6HVyj/ulFQ4jj1ufonYgB5Kbj4C7tIEmCtsSN1RdUK
kIuYrTbm2qY3b9RN55VVXoFNZ9WUIONeABRwJIjxg3uxyRIGMdCJ8gtIMOkd6DrJ
atG16D5PP2CqiNxgDfgLUfUHI7Y7qoUuIJKHYYGSQ2T/ldUBK3FMmp0mtN834dmp
yYvNBQHWwOuZEAJPgkodvWEiuXPPJlN65WA0l2Tvw7zWQh9yldQicsopghSOja0b
6e5jq1eArZQHvO4pEtUyAOaxdTSy4WF7SUhX/APpA8FCivTrOyLjf8B0pgurxete
`protect END_PROTECTED
