`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DEA+WTuYEwDhVKLUzdLWI52t9DXTZuquQNUPkLhP3ak0R3SPp7q6lfKCBWGCJMqn
52i2+E7bC5zhoNXWLvOq6jnQcYC+FGSlOOKBnCTQ3s7pBUcvzT6IVeepnamehyBA
KGDs/lx6re/ottbVoaQ/qfhxVOR2MgwnezPvO75csf7SBr5NAmdaxQjicHyYlCU3
YHmsY0JPWpYvP8MxrtyACk460R+SbouT1nc5tXTZ6nCgV0EULnHRBNRewx+2fVy9
vDx9lhNrTm1t8ddK6nImYFyGs5aPv1ETlwvXt8I+g8f9mfK/qLoc/NFlksCGZD9o
haSX+dUOAzQiI31zsLN2Uia70DE+7FWvaCCt23Kmfag/CqABv8a4Vs8ggs3lg4uU
DeLgnPkdzniuNVXkTAlcZd7BS2sKSyHiHqOnEX6ZeaSmuqHag3hDbswdNETG9LFf
fXdGXMLcDA/e/lonsVBMAyBrdRQM5rCI5iCVpy4w0axZ/v7lY2wHMGarFnI3QSSe
/lm+/jEnBTOlLBqst4pVFKuBKdoHtkPrLyV9tHkELYQ=
`protect END_PROTECTED
