`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgfpLEhP4IUPOta4VnigNyUseEwTogta0sfDyNV0QrCC4V5QhOoW9SwWkQG+smtC
mJlpt4A+4MpaEkXY4kSKPcp4YDlZQetpTXjPWdkg9kvDKhekGizJB3cC5F/NaEI0
0utOhKsQ1qbPnF+eP6nc5If6ZjrULac7D9cPfBfZhd+cR41DRZbA33Dr2Jz5Z5t2
xbxZxu6mTcadQlYxhHn7SwDI3vS6cqk4i98JxsNjxnnBc9qCITak6XckMq6/PuCg
QAPXcGjvYy37BpDA1SXD/6ZXwbV+DXu0jkdpV6NdR6nB4/rYiFs7SfjMaGVlicks
E8P/bYoW8Hx9f9InoXOlvuNdAkQ6Zgj8vAH4/+vIUzN0nhlDHG8dOCxbKUIT0HEP
YjkctXkGvB/t7jP6WqhIjtsleBsXDVPf6RBVeYDLE4HqQZAE57z2WsndILmn5AK0
ANRRN3PKssPt4DM33NDfKfmJcUP6XjCmCn6perCE9Jiy/byB/U/QsGS4A5hQTobv
3yyOkTIuRukXLDwhTGJWNlq437kYajiVXpvnGkD1wzPywJIvKJZE5y3g12h25sI+
2uQ1e1s5uGNUh9NFONnAyvp5Cf9iuOngZ5GOWIpIOrFsBvXzQtzu2QmNFGez+KVe
fRXydxFbkzkM7+Ksf/2scF6qgaq81v0JZaFKjWYLKoshvEh3NLP7X7UJgVFdYK8D
XA6x0jUeWSxyfaMRXTfnKxL5hvb1MhfsHliQ5kNCaX54x+gy5cIR8hxXAgkauboZ
RVTYFFI415OxwW+oDlAy2llIu36kPoeXYzbbw3k1LuNBTy41fTh0tyKQjgFc+nvv
S9UuZFi/HYwH4b04lRu0OC5ROEc3MAsRKMgpBcSTbFG8wtOnBrGpT+ZmUjTSi0Ol
4VK+GoUDdwU93M/BzHxuqZgoODtplzU9Asv/8R8V6bSxKDcCINS1GAdnzHXTzu69
DFiyT+ZooQ1JQM60/nk5kftZ0Oq2W1cPQ/WIjx7pWi8u2faLw+HT4wkYNjwq0qAq
3yloy6DrM8GufZUHgCTfWKKBmNjkOKN9CrUUuBVre8s1X4tg08f/hsSuOWPJ3iBP
lvu/1o10E5cnn7hUK1MnRm/UFnJwkzGdOWa6EC/rafTLZX3MZNqsgRTQZNrt47ld
7qvvrgU5bMg6sccFwNYfReTbiU5QWopYKbpaNayf/hYiS6Vyzm9cZ6cBVO+afdoO
a9y+hugB4HITZG8QxB7eVJ3kbKQHaOjMmRDtGv5Ko39xPldTYLkDozJGqSCHiiPc
QAOLfnG6JMpZSPO1q41YnPIb809CxsX41yqIg46jYrK2TALW1aIjQ1TMTrszZCq/
6PxXqX8cL2Zz+oPgI3JqhEg3DpPZe010445MYrqA/z7wU8nyIdOVjcfoMamE/N5M
108xe+5O5uwdre2dfFKwDuWdOZitLWfpivc0/xCAOHW69UD5/iBJMpmhLY0Tkjtr
6WHKpo+unfjx88hNbA9YTqpOdpbsPRthat4y9mT99FU=
`protect END_PROTECTED
