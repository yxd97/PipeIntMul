`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOhOMhOTSaqYEy2drPKL6e6zubie997HNmlmiyfz+oFzDeUgJovDxCKP9S7g3Nbh
UaTBYxHliU7o/dOTXahEMWu9MqRbc5NkMJf/PEf3J/kQ2UzyYlm5FWEGvrrUIxEq
N510Rxdhhg3BvH86uyjMNAn2gmPTvOroqYohWK3HGY9O/wGCY2hRMkANuSCBPkt8
2iL9oyzlm51d0kcDNhs+PiniY0vKQ1k3FKR1XwLtmSSSvNy2a7gnkzJSCcQZNGRs
qcTttP7CMYNAyi5HhUzaUqrISaFPPv4JebKWDITHqUfFmaRALyfQ5bZFO93Y6x6c
Sg+SwwKhMDanyj1wHgxdL5YHyfAv0sHeJRExCDPEog401TMiiabFdJrwTEz40dfe
1MecIXMqLhWzC8hxj50A+OMovOO6U6VscddkQihqWXKHoajDnNHIVslDL0o6Ljig
SBhUvtG0caY/wTZQwCu6XsQQ4zgvVCb0Oa7zYt0sUjPcw+y6NS5QzP9MmAiFvKeu
aUvip5CKxe9dS6Xa4hJi9A==
`protect END_PROTECTED
