`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PDPuerYb5G1+jaCaYcvk1msAERD56OFlOVKsEE0skzqJDG8zxtYPZUQeFuYzB/Zv
qbVsvLOP/t3hXRByFHskqsLuJdRuTyLvJDyad3QNGvBcCfrW4LVTKg6OK7DnkiY1
45+GBTwErLy0Mr7/YrXW1LFfFuxzRCbbd3ZcJnAsxrU7Tl4h8ECqc9kJvTKtqYVO
ak9v8hNcHqr8nKOCaTG8pBVedlbX0/JDgLe2RYYZrpM2fPtoAWuqX2neWBmpxGvg
MnaDT9DShYGkyBKD5gKZHFED5jVxIS+gW8rP+rjGpkEuKWHSZJVeFHAFQfR2dz10
nSFwre2CrKdlyIP4WBemHFv4nDRHdcnRze76lW8XbVwLSBnvjUeOZeD5Tg+p0ulU
0lZwE2Dy7KH1+JPo7FGLlg==
`protect END_PROTECTED
