`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tnPnzK/y+XHnA3Itm567CoYBxcz0ZIgD2WyrRRuCcf4JgouNVjgbbBZFnfCMb3Bn
qhihREMea8KbKF8V0DsTa8ziA9t8eYCqoF0BosXFcDuiDuBszlbhBWRDFrTP3j6E
E9QiMKK6tR1TbO4YgiPv1URyyexSR1VVkrCqHyI6lYCArVgWjMJTK5zaTNdf12gA
ZhUsXSynCcU+75mU28FSqVe3Qdfxf6PuCnumFwX2HnrlurBbIGCYE2UBufFkLCk4
`protect END_PROTECTED
