`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v997Zynzan5F/TEjttqHM3xAbXaAt+82WEJBb0ny3DE2ofXTr2YrBYnMA8tj0VWy
y+K15eJNJ59pIQPOGF1NKeSSE94WsfblcF/sJVqP6eb9uf0rp27TiMqjX4aTH/K4
vOJ13SXmxDFPYTaLLge21dvl13YRinYiuhzq60EVEY5S/qJJeL3ZrcEM+mGwhJ3b
8+QeHqmS9SY30nQ4+aSzoxSDrGIRRxjDX2OdwNq5AprHdEg9UV7xihYoJHfFY5nL
P1lZynY0N7mThnEh+DYiNA==
`protect END_PROTECTED
