`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tlpwq4rTKAfeWtfhDDMj5h4ekXOvwAFPep5TPSbAUxB+915d4JZwWFRNQtfffuhs
ZT+slnCuAiA6LbaH+MayAY7W8PGu4hoBhTfEHFjosCyD5SOlUX23bp8okzJjcA6P
QcitwK5Fg/vc9rqx2+b1cl230TVJBq9t7lUsvhADLF+ZlRvvsQiqYxcbDOCU4VNQ
6NyMdrhdjnScKD19srQP5E5Q9ojVMj7/0d5hvUEsfmMgWMTj2varWBMsF26jz+N4
SBJbOMJzvV3bcnfIKUZ0zaDb0lKPEX9H3FS7zMv518a2sqbPt87d4CJ7FDgLN3DB
49fGQLVTfYB3tHPwqj6tbRDyKdDfBJWy0AygWTIDgr4+iT+BP6vQc4B8Clv3E6Z1
kIECc4v3psQ+m+igVgshxWKFB59WlPtpqH+g12SuCAfSUoh4jGijfk1so+OBEmoz
Qn/b2PhIMFkvQnZ7eoxPvIXcX40OKmMUT6duOAVgrrxHJb6z1VP+b3uwOGLCmf6/
tSRMvXHfTg4oVWUIZC8gkjUe+chgyWzBC3brOakzC1f5ISytK84rLcajhA4gDKP8
28k6WqVC8VbIuife/DuJxlNGxhhMmlT6WWIv/ywkaMAObtzbQ/MnAcjzM4ZMez0c
Xcf0kA44XKJthVmYb5bZmHANyBjVoeQhHEeR1JHhF7uGDs7rcXlnJUgsuPqKnpwN
`protect END_PROTECTED
