`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfA5+8w4SxBvUnNka0/vFf4KlbGsybEHepzRbU76v13pKg1S3ayVSCv3ib+Wv89m
0XAo1nNbOgpn/vG1mxQvzSaQylTB/F0aBAbOzSbUQsZAZbM8pVZzDIOrDQWfjmYy
yxSnVK8YDtk9M29IAQKVMmL6QaHqBFo/qBUB+KQYQZtjA3uVkrBacHTv8YPmpjDd
VHdptbW7UtVmKlWUngjVXfO+GeQ0drbIOeIWfal4q0pk6WNwGRAf00WNy+u5Qsb8
niA5NIYRyLapEgB4s5El2xbGvPEceYQIOpikjOYDelDlSHizy6H+RBTOeWAIBsm4
gcuW89zkcnOrGodW4H32ag==
`protect END_PROTECTED
