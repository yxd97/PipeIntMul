`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QuX6uJoqPrfaWiJr7yjIbMm0wAB+PRTUDO4xxTifgf8DLn7ibfplTa3tBkhu+vCx
YO/MOtGqkNyh6Mo3aziDI4VrTwAAfryYWUY5t325/Y5qCBBznav0oNe+XfZ89bb2
ATXF9SDYtyxcdCQPuN050llDz58DJN4yJAUNlvBmPw9D76X9c1ZvNcPTV9/pt0br
savo5Mr7U0Cxt0fCtvnlrxbfl2J07deyCmQ7A92d1NkoJiA6zyhB5JJfs3QsuSGZ
ITKmyN7/L+JgUlu+u6a7j2CRXysLLeLZJF/GAeaiRW8pa+i9BV6I0PtGn1cddhyl
VXumF5qTnf23BSDJfNNMYlXXJnHLYeIBLSu9uZzV2CKZ65K5PMJD040Sl9OUPAVZ
mYnrujBwC4bEak7fnxHA93khtvQtwoQJtx27WooMiNZa8YhpYar2ObZBxIduy1AX
k5qbYnFN7Njf5IqL0x3Ge/SMf/7zzWTwg4BW4mdUdawUGwC3hhB/9LKEwjNsjD8T
Ko8Z7D2M6O3DmP+6JdAjLZfZYvNhI+LIRJs2SOUET2/4wd2BJ3WM210I/3VNHZvb
UTotrarSRuelp4E311Z/ZG+wW0PwDY6PE3u17Ibf03UkcVLZ6hNERgnF5C4fjQl2
Bi9eGajVhBwFEqorwSFn+i3XYx1KG8IV0sjl/e0fvSDQUJwjqq2fkLlD67hRQ/ZV
L1TFQ0qRH5r5PL/PuBwSyGWLIqPC1rYLiEyGWidj1i/fTPZxvl/nw7QIZva4a4PA
pQSGxYY9SOrlmoIqaYbx31NhY+D0sWtSMuVwqX+D8M4uPYw+S73pDxk8t9Hlamjm
eogsTYtfEHDEn3/FWY0jQWnFbhOwIS7g8Qnm3rikvMCD5YllegILevQfDtESYW8A
SdiYrKZZr/pXxjomW+g2g7g+X68GtUhwXF5seBKfMNYzHKgyniyrgPodgK663XkE
1WzCjEOFC2/2vzMN/VCpvLTARgNjiJpU0RFxuPXhQA8=
`protect END_PROTECTED
