`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yo8uzkkk7qI2wFJO9+i0MTeYDwawJsIaYWgDU1SgJUPCLwRgS5aSgwMPIdcpYpfT
OYe9Nm+AAP/KZTqUCgM5EC2Gri5Si7HCIeIlnOJrEZykz2CYikyXKhwZUoeiKlAl
qW+3UaV9GpTp0/7xUrpiEE8hwWZflgDtu7XihHdeM63XkAxp57H5LbR4AAIMim5b
QbTowqba3wh6K0lwUZCPKJhWy/Z2e7ip3RUN5l3jOhHdUU/ipbRTwWMPA/swZll+
6lpEKJFXHRbTqiCIdzubOqNmqS8PixyL1w02t7ScI6Wf4TfftyoOTJxy79gHIPrR
O/B9LrCxwVAdUOdMiEXanpDjT8acBLiMIGfoRoxLF92a1kCXeaj/in+pC5Td9PSc
E5sVfExe/ZY8KDTIceV2YEMSUDnlWMxIi4ww4gtgoDrEhMQn+6thMzlxPK5tHgnl
kHqJWnhtTLy6sdXZEwe5H5nN6RxOZyeryaV+ohfdzLAjJNMAx1kOzTvrrXDn/q2L
`protect END_PROTECTED
