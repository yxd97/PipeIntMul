`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zP+CPIzWo3gPVpXgAuhniBe2ih48MUILosoTRAltjvbDspstWNIw76JrbQsNhSbU
VlwfE/cW0dNMm/nC1KcfevP+uBfy2xgURVjQ8pSvy1FDC0F6mZ43Er6Z2nfhyltu
Qa6W3eIN8OPZZgQsd4RFiEHd06GdiSKvXGQvpKbZV/91tXGho7138GvlqxeCxZMl
xZbDg6WTGl7rQ8XDpnkPQBelG2ToRbUMrit0J/PXyV584rB0ErM/tKJqOHkaSj85
USjoI/sHBYo1K/WMxplwh9+w0JcNlRo3qMB5gKJGjgjIoWwr1VcmbtOP7RUjuAeZ
ru71TEO2Oc8oM0gKd3mKKIxfC53jxFD0eTOTBDQW2y2yslZKtRghakdoGRhN0w/h
aftrl39LF5NwmA7/LdUbaGBmotsGk2h1ZegTm5MeT/xjTokAlN6ayVKHPCUMwDRC
J1AraGz7L96NX7rYFELLFtvtDiBeokb18+jgbHDzXvUsKPPFi+CRlnkeLB6HX/xL
`protect END_PROTECTED
