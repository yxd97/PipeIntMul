`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lsIfq7AiWZv25jkN6bsPF22Xj9qSB+L/qptLa6UxAo2ffIh9d9hOiD7g/NoKKoU/
6zjmlQppo8Co/eClcUgU+lY0zOWtLRGd4DS7N3WhFXBhUDmoxEpMdYYXGq53Uq4Y
wkjm13QwC72t6Sz3+wBxRjNc2SydlOsU1cFcWyUwTChT0FdahjOQ//v7YmgJ3fR4
qcNauWwQyXldvv72KlvASOq/NUj2o5sKgjBTy6YKyN2Gtu52ka+dQW5DSnWd05Fj
JZc3HjjU7iU94CCVcs41eJPc8GGgQZsQ7tVAVEUP7iJ6WuleAhJHrkH/kRY9p50t
i+XXcZnCIy+YH4INQNFMBQ1FbLnhbyhZyEsKa+CbiXEyikDKdpcAvVkUIdAmXyov
vNNS2stnPsYxP02VkDTsXk797IwBf4HxlXJi/OLhuqtcbde8vQnLrnsTdjIYkO00
FxBC1HDaBj2Bw8yr1Ki4MXzyzlfv4YOM/eukjvAggGAauj3Hq2FlKnGgz0kbN+0f
DAMSdlj2YqtCtgykSLvMf/qKPnHKwH+c+KMezGdVRRv/peomBaGTAu0iqichG2nq
oyweqFN+KKKlpHXNBvrORs+PD9e3kjYxP8RFCwJVOl85H5cESKiahaHp9Lgyn+YC
DEK56x2U7DsbEydtigoEDKUJyqFz+IaD5LVDAazCIpk=
`protect END_PROTECTED
