`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GilDyaB33toi96YvdGUgkDJo5msHw7Xql8mfskR9VLLgIe1z0A49hea4cYnk6aOo
HjAIvMVOKm/THmKZzc46BCM6moRF0ELAN0hY9qEvvvUq5ZN7np0dOCiWNicwNxxL
3p5arCcsLB4CalL/W+TF9+tSg0EO1CSx+/QkDeYn+VUc8c0P1vRwWF+7NkVGx1r+
CwYFihqrVNRHV+3Z1fhOhJZHeAWupNrUp6FUSvGtFD9KOD+Sj0rwH7/NybdsApvX
t+fQ4tnIjOEkrt1O6zt3BUmRpX4C9yEUHYBUlNXVzzk=
`protect END_PROTECTED
