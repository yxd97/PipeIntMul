`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmdV1hoAapYlvo6BgPy/nhxL3Q9u3xfWqIskQL5oJqoGows5aLia0tpYtGrVbEjv
41bV4PsywEJyLmHkkyN5vJ+MLgXHtQuI//R/Nu6Q6YiysAasReE49ogxvMSIcOTQ
2A8UR+sgfoeLyuxLu7KUc+/cyMopCPha0KYO/QOmjBut0suYyGm5nkMVLVvYfmsZ
grLf9WKzJPsi1SsDrpD/zSGR18GeiCmMrcvfwEUUS+8m/smF200DOoHwLEPWJ8TN
Z+JBluNgZsBWuttkBRdb41hq0oi2f3SR7rUjCRxESvOs2mtPpTdEkO7kpnF0dl3k
9AGL/sCqE79UsWN3TUyptK08/RcdY4FabOYBq2Ea41sc0wcpm/jP5rPhVZfa41+7
4gRPEYOmyJpR9PzolnPU8/ogvCWPnXVKZqUP//muSD/XnsjKgD+aO4tXNfjDSapU
I6Sk8CM75LVz9PbsY5sP1w==
`protect END_PROTECTED
