`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuChsVycEKQuskq+vsWGcYxmEsJg14Io9s1twcWszOaCNDn2kAW1BwhaN3rkjtVt
jk0f9+6uSdOdh5TqcFxBVHqHZFrASZVD0TBL5zbj+P6EgeAzcQCTfdrLyhqxketF
hvJ9Zky0ph35nokdR4GYH1gyoDBBfq4HZT/hQNGe1Cx3p35PtzxkY1SnPl9b+WSh
lOSHvXDYsmUUeW4DZXaBOaI0otE+xlwnIdfXwJos38vYYb0GSk3CH6rK5M6q0JLQ
iJeuKVfQfLLokXKTnaDFJplhN/HoyU0nSBpmV0eW7os=
`protect END_PROTECTED
