`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UxEssKe0NJCsrrhruRs6YBEAQaXA5LaVlVvuN3hBgYabTpUPmc+rfAlop+7qR1Bg
n4RpjBOOJUVwcUZDJ9y/eN7aENuD86lEsKQCNSFUEzWF/Ywo4HV58VstLmrh0hzm
JK2CG5CKt1VK0UHobOiQmj2gMeatShR2exodffwJPoMPfJIqXIFt7i2Wv5YYk34P
fs8DN+ZWag4UkSi7f6v8r5RHPETcePRZLuzj2LJbX7XaIbLjB8jX0dM6EIs4gmGg
+RoLobX4LOaHZTUvN9pPU05WBARm2fTwKAqaoC9wMMXg/HR4nOwJt5YIRtPeiGDQ
sgYLAnhywhpbehXGpgpVivIC/OAzChMjKi8WmWHL2irXSNc/u94WWyDLVW7XDyNs
MuDqlFTW9C9aYmtKbQJJWyPeXPPYlB4njeau5mUfQYrXeyOFQIOqitHvvU384X5K
Qv/mlrr9hfiDBVtbQOpWW+ovrlbscwVL1rheABdE5SG3I7P/T2TF2lhRU1HCXYi2
y9WAVyFsx04cZ5FkikgYeHqLtdMLi1rD2O6UScaMQisuSC+ks8Q1FRf53aytS8te
5YY18h7LsXbAnvhVnbiwdQ==
`protect END_PROTECTED
