`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
08EoyzlM2KDqEFB1HpenjLAzZUu76EUQCL7O9E4wnaqgPS3VCAaqyZj9runaHome
4L4tCreZN2P0cEkGxrOG476iq/G8FVxvo05t5UaOi7OE1JlnSYe6bJqqtiY08NRl
JAw7AzvKPeFnPp2WODyh7PATKmefx9z/cSn2PjqMONdYED7UhY1i7jZXOQpzlpTi
KNmbu6dSSBDobX8gblx05hdAyZBKtGU/mXFs9N9Zt/9hv9PV/qUs7aJt6lysK+YP
rWkZSUhwYd8ePp5245l32VU3XNpLXfW/d/txeSx8sXuVJH98f81RJbutX3IX/RdS
sqL1tI1KKP1uEFqJrZj137V3RSMj5zFtcOGRJb1PFKgdvgf07r4cHzO80WGbn2do
JXWLfrzM2qVzFblPU3DJAPSmd0CeckLCqedHTojXz1mf5lOfmagbyN7N9Nc39MXc
O7HDZBLo2+Bzb/OHqaX5jzgkYBhiSSfWR1+HFI9J33BTY52fYE+mTTot2a8WlP4v
j4nOBvQfWnm0vrh97d9zqbs6/e9VtDBeY5JCUyCvpMt6o3fy0zt8bM0OO+IlRkyT
KE2mnvULh0N7sp5/lVTF7egAPV7qtVC9H2hdzH+veDIEZ3g6naBEE4m+5h3msXuv
Z2HYGCCHkIfqU308FXDXsSKdIBwZu6HlBkcXkC/JMyXe6/vgaa2QOVrAY8kT7WmA
66TDDeO/oleD2IovJ05iPQqWFXdgvNd94ZiAjiWm1BnRe1E/ObW38JhNmAj0NMVY
nttgb/Z01SaCx7yyvVtipaAccgYt7HZjNilTci3Gu1Uy1CE3RhTeAEXm93iSQpql
Y4YtWhY0iDiy033iHnoSTzXtTTr6I2NBe3AIw1zWk8Y53gMXkt8RZniDzmykCIas
eIbq42OW6leS1MQNhFl4b+D5ZiZ8HGeB73HfDeW+B25KsHSe7esa1p2Si/rr8HMJ
pRZCgG9fy10edu919xvHdNyrdMxvx3wL4nBFoR/JYkQc0WPU1CRkzIEZ+a3Nhcld
D08h5ms0SrdbGkhSX3jHrde7/R9beGu1/d9jmK6yzRh9wIdzpY5Onfsm9nCUtfZm
n/hZaCHc5TD+OpfIaDZwYntHciB/JdKQ5lVvqif+x70y6egUJT0EZNb4kBT/0AdX
qppNg9WllIclM0zqUqjnAQ==
`protect END_PROTECTED
