`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvfmAuSrohRxhcupPgp3ymwLFXYKJkf20PyXDG/yftb6RnWmOKVOiP2EM3xvspu+
BcfAVIJU469OWXelJRmvUBlxGoq1NbyIYE4JZk1kdkTCBAspZ4ZHTm4O2xbh8mxK
jgpzDgl5EwVBxN12n66RIwkI0HW3hptYr+mrU8kgEoTRPMfbWvqg91ooLqav3ook
l817QcavHxunh91bBIjq97T2OCTLYPPcwONKFlZCoAF242NAMzotBj+iR8V6m1o8
LH9Unvddipq6340wW8Hy1/ziEIydf3iKDjkGk80mx7f10mzfdWegh2Fl7seLyhPx
eD+3hv+PCWWUMHPJwlA72wrQXokZWBNHGOv0z6/GG8dmBFruttB0T3ItjNHwEQhp
uC6qE+Sy2UAYyfC7F62tM6YGu9kMNChZ8IWSMVf7xhkFuZmZSyXjhTLyVClXvpcR
RkP+WWwSog2AKBACalE+lEwZZR6ybCyN1K3yDxlFifZo0V2GmM/z+Z1PalJAU8uD
Vr28KJD/uiXMt8u7PVKHhlbWXhOTxInQbdGhV0TjOkhoTjbKsrvnsBvJYss+MZqC
Cn0i1rMSuylmYnGk6kDCluGJelBU2A/9C6bpZxnLN19SZm08dZadM8cPfxcyZcKh
EGGuNEXmFZxOPa0HW0iGMXRgMozDlppr2cfzsO0fZsYsP8Axa4syrc1LqRD+Z9Ox
kAzIhhTlyLi98YrzFU8sww/kJqdy7EQlNydKYs1LKRaFLruVWKdjCB0FspQSDDDc
W+VszE2gWMcCOXjlLLzE13KWXP3vupNkXQQYanLxCXhKegKx6nE22xvpT+4AWKc2
A/WuqDtTolkF0c3Nfv17b32R+NAJ81kSWpKgwMV5G5pAsXcbdvjIJzD8CAxkvn55
2XQ7A0/hIC8s1SqydnAxJla/W4SBmxIK9LBsUQNtW5Unoo27OxaVEmLVtu4WwJ7k
bDaVurIriWM8aSrJTg70N7tCr7jnjzX5Oa3O5SA3BEEEER1CfAJfmdEkvZ+LNSKx
qcdbbN1ZKmbNhbIS0Xdh6uJlBRYOWNW0qjbdaviukd6w/Mg2vPqB54pj0dHgDQ5b
2Lb3K1IsFqegIcykAtAbmk4ibM2higP4O7R8A7j3iXJqCB8GcCxwieseQQdt7nAQ
5TuJI4MGNIBqOcxiq0oeYBr9wsFOJ6T/Y41H52JMDlWOTRBAgLHWQ0XyDI1L6Aev
+n5oF2+HPS01X0XaN1FYlm7WvSzeziUl1agOeLcJ68ohJBNHEOFXk1lvVMZFwg94
YjlVjTLHmFB+EDhRLjkMG7ewJmnnvKSVD6EqZIyF7PWZIC7Svg2XKjjR5vJ47lMS
4RnmMLp2k5ybm1kToeKE+rMJyhPDbgfZxliRSI7H6IC4A8njNgnQxPixrE21GdKg
ZedweziqyU4D9jFslaZirOVmFGSgkMIrXhEu9wL2W2VqXWv67bYHeP91GxTE/HWK
GbfGBrYeZJBg+klhBM4dW7EhKMqiVdei/p+crvSDeoDhSYg8DH7zCcL/6j8BioMY
bxRUawIjS4foj8lnrXFGhvklvHGOQ3k9ELb769yzQtBPfNRD7pHvnxUJGgd1UAFd
xO19zI+w4Gcrv9Iehx3ZMS1fCcPIgJPOOW6pKv18jBHWNEf7BqDlb5y3LNNiB8qB
3kuSQML9mg2Jx7y678BRlArlldwbHwoCWeApx15ZlwWFME3T5rC9kyeqRyMA31bl
Mul4Yyap959nEtm3BNllb2IUV6ZF4pKUxKSzNBlSFl86opaByxisI7t1LMFRFPix
ZbD+HlEfOCdRAOwsfO/JPrAi6gPqFNiG86i3X4+JPlGDxFN0in1FZj5TannChSkm
l+gAvG8JTAFUdBRxFBspa6K+RxVkNKGkyO757w3BYwHiuUqrWysMYOAS89ZBhuFv
NLCbNbW4mK0G+hJOtetXpvARS4kmEia5uRbOB0dstCu/ftCK1ofyyJ5/TZPPNaAQ
veQMokyXlG+JIRYk9OZjr13+D0ZW1fSmCmzBUdD9dO5Csfhk9yeMJJamkIfYVTsf
ZcWlAePJYz0v0hiJJ7LUlVFSVzJnb5gBQRHqdkbuaYkaV9RB2dv3wWwx3wk35eFB
fZsHpuyYB2786UJXGSOO2QmNQyPfpyNpZNLWqlkbTOSqTn7TM1LuBbBreSvFUsXB
`protect END_PROTECTED
