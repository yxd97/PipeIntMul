`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EZ/RtTUGawIOXx5k8Il6hoRZdxhbFVkMgwTwNrwjiXcQzV9MGXiRULlCSQntTczX
RcGYgzwUWUfNEOP7y89abMLDABc53dVlhIi1M1FN+9/wOvPCR7mktnUfSVaOKFCS
9NKCEOh8JmUTX5fprN/tYE3s1EycZyRqWfvu2yYO145VmswkfREkWRsvijLUsCUl
GU/8zsLL5PuPWEOfwNpDs6nj9s2LjX8dwa6/LWK+PoaTBR7Ww53ybiRFj1O4q6y2
O9XXJSXrtsYJZFfuaBnpJDJosEyHjNGLQdZKL5vY5yYUTJBVAvLyEwDHCstLCTe9
j5qrEpEeaL0iht+jLWuMRg==
`protect END_PROTECTED
