`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYmNn5xtERvWPAdml/hHK8HukzkuoUWzMqM+vLx7piv8+pNN6qIN9FA0LBdvmEcr
CU+DnuO9xLtTNYYEgEE7DM8er3NqJ3wL+GLITbfo4HbjMFgkojTrmgmBF6X1N5Xi
4f2R9dsVV9Gi/7/ak5yBKEMPHpR6DO1wpgorCQLRgJeNGL0ZL7N8BYZHoDJGF1Zz
btLv7785+fUJEcZxTjtAVP1OEqmU91Uoo9ijs39Hv3jtcfTMkYLCpP/l6DNxxy+e
yAcHgWJZ+cdHfIqhcY+d0nllccthGx1APo7rk4h3T0Iv9L+vXX+Ad6OnF5hqZdN2
eTArTPzumGMdhvUbXFXYSFluKoUeuRTMTaQ41xFw3IbCwSSelZLuLOzoMegKbPPF
Al9NPhpugxLPqO1xWJo7T3ocByx5xLxBZOEMwOBHnG7WAmMplP7tK+StcbO+WHu1
wFGbc3iK5Wca4bdtB2tpcgLSYGi+odttOcZp9TzjqqA4My4VSeC28tVrcZamFSA5
MKCsh6bq8j4/mCeXSVDPAncMiiC3F+fg+x32Gspwn2+MeEDU9Z5WIY3FC4JqdsNp
m1FVyx6L25iJdrbR+KoN5oQopFBORtu3mrOwaNMBp800UJlMEGVC/slcp77fY56C
EEFeId6Rjv4u10nGNGTFM3ent2LFrg9MUGezKXTe6jyyfjfM3cscUoO50ZHRKcOj
embRCRHzICqjvfT+b0fB0ZVqcUlOOvRA4jAy9NewuxL+5XY+5j4/dobkbRv2W3Md
xiXeckjEE8+Xgmxg9bw3EQ7M6rZO9630Z2ytS3CDDGjhSwiIYWc2O/+zq5mUDghz
0yIG0zmztOrW6mTv4BUO5yYHXCVTDkxpRjMSUU00JzRYHekEpsDGO4+WUHFS47qZ
2m3ojMjux35JytHwR78AvGHBkRebTn9T5VGS10Tw3wmQR3bOpzqRqsnNx/sm+pC7
ElBrsBvMPGhiQ4Iq0LsHy6Jf0QGSVlDgahauXfH4DtlI7xdhjf9hsDcaWPG6KQ9X
VpaPbf+I6smBNQItPNf/HZHiyB/bqQZAIvQuAdbKiNRCT2KQeuQYk1YcoN9lRLqq
Ieg0dex9UDRjXj+4dp4uvg==
`protect END_PROTECTED
