`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCM6pdriER40BGTrmi+TvD5WKfntlc2xScPffAHJJNO9qiLkJePOyJczwYHpL17x
qqMPeiXCf+blwgBUMDpINZlzchqps+bbbiyr+8GtqTW73//nJJ82ATSR1ULoTiQH
4gmbw0fOXWv+Ih6ulvx+eTZUV5F2O9pA/+ONzlU/mi4h75WFCLVgD2XdPgMyuRSp
HhSWIi/SxSqNDUjsm+rvVFqXuKiPFjmuAyVFTO6IKn/WhTjmLzeLAvg00kvzIoFE
aNDiW7HsZRN4X70rNk49rY1p3TYBSQKhEA3bnquMcWfKA2je98b3zDCUXS6SVufJ
vZN8YvrMiMNkZiZgKb5j9McwbrdfWnwZixZJ4PDWeSGUk3ETCf+Th8/EYTKN8H5b
RQKxeZi+hKbgU1plZmM1jwOa0/LBzYAW0A/erJySOzPeIk7vum5eRPle7mASgTa6
d3CRvFhEidoraxIMmdGGDo2Jhv0OwNdaYNzkbQYWlMRe2ZOzmBN2lAWouZObN9VP
Q/nOvu1RxJPrwPK6/7luMbfo1RfIMBL5gokJxAoWN9MiA/aDpzkD2eOD+5OGF/do
fhWQiI4dEftb9hX42UZpBwRtvT4vW8OnUY5UcaTzgcZXQWQ/6W3XYTEyIETu87f+
cT4pLWOPG8gxzn3F7G6wwQ==
`protect END_PROTECTED
