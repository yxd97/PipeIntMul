`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Czwldso4xURyuUmzLFDLKfB4NJV+N4DcA6JmmTgt069VeK7yaiwjxZbbRcIzGAnF
UJlY2tBwZL0nNBTucJV0td1p9Sejtd1KPkGqdgNPTnXUSaXQo/LpdjLJgK8B9Xch
7zElmwpcdzjDavLvn04SDB1Wf06y/5LbMTd3gHdlmehmZo6gxu4sdol6IstDltGq
E8VHGSyun1w+LUUFC7TNSzOx78xiA1SlBW8BUUnEaO5frKYGiKlhw6KL6Xi8KQvH
gPIdrW3izz987wY0vWdJNUN4cvBZO0RowLgyGP/NO2GMdqDi9iUABpudZSReLoGH
HS2qTluzH2u8/Kct66EOtb/VpX3cgYJyavml7uXv4aN3M4CJFaEgSLsJr0F9AXAb
Aaf4RbRvyJOmY8BfUA3KPejwHZF0FsYvQQymbABrbFXy0HGbAzN/gr2gJbf9j5jx
3k8gmSux4950PppPBMr0xKVjFgTQTUXZV/y1RdirupYcrGtPSk7b9ATeseYohD+B
Mh93NUWr64rxGqKDQDRpP6vDhW/hHCSvl+ZHGoLZmc+N4e+rD/3H2ZclEG6jlb5x
`protect END_PROTECTED
