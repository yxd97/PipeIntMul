`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Fe5BJ4trSgWS4J693IT7shsDTtv9ElcgKn3O6ElUVTQkRv08EANmDLVVH46TGVv
jr+RuAEWVnNSNSO/N5cnsjbMJpbXlLx1GQoO8CuVWxim4anejKgFBnTnLgtxw3bo
XeDNkRVt4MLhtO4dKDmOpMjymv/0OR/amn9jA2qQAESGCirGBqGwzgde6zftaQh+
f99STriQL0pG0n1U2xeCzRAU1Phw2SmOGeKWvSIb3nas6N3l/ogYeAF4q+ZIwJn4
o4ZT8J4wF52CvoGMgA6D70F/GUbNMQk0tKeGhcPTRHPbD2ZmxMlEobIhsq14cl28
rCH0uOjK/nZ4wG8hFXPQJA==
`protect END_PROTECTED
