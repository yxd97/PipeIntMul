`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gTxW+pPGfZgTOZAP/gelzYbP9ZLPUDVk7rM3ABKtLa2CvXAMX2QtTt12NB4wvG2j
0N7v0Em/+3BQ4N4M4TECiIJArUN2cp2W+x+8MjUpFltU/nLMA1raLBbpokVcVxTX
Npktel7ZFF2qb3mfYE2z1I4GgMS2SqSc8Qz9tSdcay6STsQ4Ny9WOQnFSUnXonaW
Ij6PpRuBFHjyCgIpjdKPgLjOmfsquvFgCM1dqyitMC3sCCClsVuQfG3tSA6yr7Jm
UArJcjmXBm75gAHXddPFxKAgnB2nEZFR8iXMK1/onD/pUsU1KI2domWmEyz7RQzN
0sP1gLySLdNlvSHE/EPm/+FQ4Ge3uIigczu3TLpAUh/RxA3n1GNZKNBTfSQpDtYj
ZlwWktPnTor62Dtn9GhrJHJ3gSzlEsbTwK5ktNQcrPf7xFuIRi+a57ia0FT2qGpF
`protect END_PROTECTED
