`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jxHCHQqxIA6aTfBExQspqCYLHz+b120iqjF9DqUnwcLKAgeXPfEHH12s2mn7A3oP
0/LNRBSfQwU6tEh1hkp1A54mBI61fhG81LoFTwvNwxYNCr9DkX3JSrghD2/0/71V
2Ut25bBJQxupwyNx1GiN/4Tz1IdmhzG2HehK+AQ1o4Rlfet+xrImtLnAkSoccz6f
xSCLeIukacpUnDGJDcHWMoiDmVbKjoKs+DzysrdxC43Kh7/r4wbTj2GUvZGfk2y9
CPSzjHBjZZbHnOOL/mt5DdCe+Fn12VGztS8i2VgHArPctqsQs2OwF2si1kOfHqML
T9FUx8yvDU1a++t5LZJNAJrtnV/zpsDmHPL8JsJD3hcT8KpVVG/S7/32v+VtGYu+
C6wtwJFWyoGSpYqMKMUlvSiE5SlD4L/Lkk8gLt8+JIADYSVZOMesgRGAkuYFVbuG
RnOxcOxpoEtOpGe9VsYD3GxmBe23M9sUJA43IvnfyYAifjMXqZ/9zeldXYKZO1Ze
5/UesZDO8Y7XvDspVQfjfnwhbHRdttHZL6F+1LzDKlIeALmkp2cUadEAyyu6ZESG
ZV1Zw1TpjaZh5xxU9HNW4MB0zKffglp/Uk4KJMrvoopac6QSunGM2/xHBI0JZ7Ri
wrMzsBOuDDpIqamZ0YAnEipM6vq6PAOCywvbj3aiHgMbwYdk3cBisoAYLiQXtEuf
z6UB2Ne3zlX2Aci7Rryq0j46lMyuFu6WX19ZyHfV3akaPhQNtn+pUMliikChfMpg
UddiULy0CyC/+E0rkE6zkZuc5bOEHybZSmzgCYg8FnI=
`protect END_PROTECTED
