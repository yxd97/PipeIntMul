`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lYaTI6mA+x0GDmUC5+DoNBhbyloKhJHrlZkgQ3FYylyq2WMBLqBovhsqV6gl1DaS
//SHl4Q8s5LweG0FaaMrDCV9cJnnPGNTlqmk9igN5WdbH2L4Frfi8TPGIZz1Duhw
IEEB9MdVQCjv6YKGUj08yNy6EDpNIi1GJ4ca8ygj8SUlaZMDBCzf4UszwEqqmHMZ
anq4J0h5VeaWQtH0edbMJNdMG9uLQjyzfCYHmrfDmEGKpl50sZErIYoRx0LGQNgp
0MfFWHVCCwhdGLOyB2SbgxRA210UmQCHR5rTRezV5/q8jjwEoVKXavVec1XCQ84n
KNyZZhOlIXVwEFMl/f5umpaMu0/4imqvgIK8kiO/PpwFn7vsIUAQROEIeuzxydop
KKeeirrB8qNoX6dZkWTZLPvUVQkWtWZzTe21L7MJh4omej7F/Y5lzmZC2Be3Spj8
WMFje92OY7jiCxHgcrfPRIIzmoDZJZfSH6gDeVEL77ecYtgqhGDyxD/RDG27kF3y
Xs7uhzM1JxlND40nyer3/6Hv0WpDoU4d5PrwN8DjStSf5rc+LIF+uWEQV7V0UP1Q
PPfgIJa+h7rBVonKKQlp7nlOqHpZxbtxvBt4AllV5Dp/4CUCHXXljffXvbEaqKdC
BDpKYq0SLFuuE8sopHNjPDhhw/epxWnc1OZOtyLE9KYU0lQgLO6/gPOJ9GAnydxf
JB/St6RjdB9I+Boq4OJAyjyMd3185zSMT9vVt1MhVXzGdEumuZ7HIOTqB+VPCDPk
z/6Edtnca5JLx0dX8R0ahB/KA0QFy4w9sMHEpBy1f1SkuWqjQRKE8NSrxD45g5UM
GhsLp3IGY79PxqK56Q24ldMIf8Vy6zrA/5Ko1yrEOTb3/K9SX2d3D0LpZG+HPMBh
sabGyXvltoGKNtZf3zF4q0ybKbCKmiQCHT8HN1qYweU=
`protect END_PROTECTED
