`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H1muiaj70f6GCwNRKA3h1yUqJQVEqCKM6a2MZjO3EIdzaa/Po66l+/qt4NrAq4F2
StR/cQCSxqGbMGLujy8vYokiG7EANH3DO6OCuEYmWxw/39zgZrpMgYNinjuvK/5a
yWnl869WcLYuaOZdsodO3AAZLLeXBlazEWdiMRYENsG01GDLkrK3VCHXfN0aFLhJ
q5QytsoUmsTWJC5eGy9L2ufZWF7gxVFeYrhwn9eMdo+JbW79SgrvGWDrSt5JM6ec
DPsKrd74R+SF5GVEaN8DLiU79AVecUAMqn1N3KpPuUODWH/qsvJByWQ0zNg4oZvo
hIaHrrkJC4wdgNGkYE+68cNxSF/kEayleQ4M9co/DcV6PYyAsTetukEU3d+vDYdj
tvNjZ5piQD0DYb2llNzrSiW7n8e69uP8xFPO+/BtWvcwr19chWXenJs7MCK83rab
6PBBjiNN/zujgLq646/657emftrYGzfTpgWLDV/7F5uyDPU7UyYFivhfLBjGePxt
e5Sz1G7EW8IAVuAQ9Bu/HpGD4+OrC9hptEAJrCMxLH4auQ0QJ75TF1wx8WnPzkXy
Nkubxm7QCaFfdSDXzWxPgWLKp2TV6vTnQAUDza8DOy4oDoa1BytmsjFydoqpIHBJ
xjRqFbjLlYmFIpivXLzwOHMnQjo0r/dS5tYBHZQ5mDIoWDQn6xDJxXnvta53K/nj
jLUP5q+FOp8Yx5wrd6blry1nQHW//etOaTE2e3u/PjdIIwVsQtQji0HQCcKtZvFT
jw/Y7rMmWwf5U1Jq+rbTU+hypa0gjzR+MO8dDTnJ0yeLmN5eDUuN1cM9NqjRVQru
qtPuoZSWNC0BywqMKG+/yp4C8GhegYeW7BX2CCyDoTQaoyIMQncEW1rBPGtTmyLN
OL1nTwNVceDs9bKs9bEAqnMxxh+RhuozlOUzq45+2qErokJc5iDwoGkvei7vAgBT
qk2cXYlOTQXcCYiGM/4+2RkP+JHTUWbhW5vwyf8NOnT1ufOc6K9Dp4kZ954ZPk+H
iS2LhBzp45aoe85tgIUFj3UH91fV3eQX/n+2j4Yiruv61V8uV/gh58etoe6/F3M7
xX/lCn0wWukFbXur3nfn07n+Z9byMW12McettPu1Z81/ptbByCFXQzkMDVQIotkj
mL0+a6LkqaOvyw7qRN0dke4pQOCWjmg/z0TPhansGu4ZjwAqWSWjtxldupysuU/r
1G2aAg2sYsYS5u9FX3Re6V5ggT9qLTu6yevtAw7JJoaE+Y7n6YTk2MRuoAkmFXoW
B/feEPx94VgEbmewRHvKe3ASS18vzXblkt9Ym6OgCcUZpN3WWHij6ChM/yuKH303
9+WXPHleIHthYRpjZbm+hwlUssncdz/QBKifAIMnBtnh0kncBuxljp6Ft/yscSaK
0cK/HOB0iSBHSzjla9+rSanJlELjbAancmIVh0q4gQB9X1I95uD5oxVpuzt7asKs
X0P1XW9AUCrQhjthedZqUfAaV1GDTqx6hafowQF9/MMnpOp2N/H1j46v/xK0+aFU
+ranQ0BlfC2ch6q6rDLroJCk2ELYsWyU6FbtdVYFjoJg6E9/a8ZMfJ0AFP+gMB/P
EMKNSQJOqkB1QIszU7n4Z7EeUdstkkV8XpMnGqlTS0ZQi+lANSjHxGy5xyEktbli
nz5IxvLOI2YqBAJJRpLUbXateOpIyDCBI/4cen+FhMuCfX+bIRaHFi4xshKqYrFb
UpOoVhdUOq0jaJvpDh1Hepvwi9ACnbbeWEvwusjhSaRNegwM1adOBrMElcr3+vAj
cUiuKYOoel/6V6rQjm7aT7xVujZuK1nJS/VIViJ+nG5+QRlI81WFMmYwCyDCS9Ae
PzHFjcGJO1khzKzYowaU/n6MDXOyGOxNYOQTPp3VRRXfrdNaa3aLQ9rYPFgeAWud
fdnYATS/Fr7kCN/7YQ/D5z10mjdocbL9Z+CXt8HyMQ3fILOoixeer+LEdybQ7HcD
s3JWLmh+x6PqqGC+OQYHuRP6gxo0WbHVLQ3ujbq8zQiiN9/2Xkwja2axED+3oHYG
otPJWhFGnSWDfi3ua0rjSZJBhFmoSMFYSVYoVqft28MUWuqly9SRLcDJO9OnDD8B
pEpIGjODEMEElEQEj1IwQfbk7J1t9VtcCDj6zeTg7AtWVyTHWH16baSpDj45zxgm
15lJ3MHKgE7smPcPB0rp1fy+09x4x/SytfKE6fUs7CEh+TkBY4H2jZlB+V3ECTn3
Wi2IiN0UV43LvkGsAH3IUA6vBdXOHKam46I9QCR7/NhWIjsuSn2Of9qIuZdc29Bc
vZfMGKQ/jldRz3ItAdRQld7qK8jADNoUxgNduw5uJ/Tvrg/nHI7xufUi+YMGVDyq
cXZKUUYe7jeM4Ym/772E4rRsfF9k779PwX/3JDDVN3ZS/W/7rdIZxlQ9dtvUoJVo
5eHjro1TaAMDFQHZ3vzaRmvAdJjnK9O+ybI6wnd3DusGQjsENP/mVRpCDuyH3wZc
YEsDHssVJ2bmF9Hm3oCnIOL+2KMPaEuYtNKGQgn4AbhvXqHHhMLijUml/JM/CDlb
SFcdw5PbGgthSJzoPULyU/kbKCTxprJKvRLHCmF4bqRtL+uPQXJr3ueBoqlLEDWt
jE1QBvkiRdddn4FEZWOwVbb77JIgc8t97fpFrthQknb+tcSMjJcdVNgQ9x6C5t8B
INq9eW8PpptoTQ2CMtm/bi+8tVu/H1Lr5Qhe5xIuLAnp37piJjAGXWwEnnsfPJg1
+WVGYS/sasMljZbesYEqHPzrTuMKUa8WnZqbBoORChv8dLf7lbfPfM2DbShWCbXz
KLgWteb3miRqDDHCL43aYEDQB/eLeQvbZPL22MKR2BvljTLKHs482OhZYH27U+VA
nnETsgw+zOLFkx6GNFbq82CQ7JbyGWaWTUmkL6gNFankE74dqD6B/4kqW5/v+TJi
2ZNtw7hZ7Rtkg461PmDBjvcsqV+FunK9uS+ebgrqleLoWjStbQlyrh54anz3IDqe
7nx3a9pynTPJZhkwZbRQldg4y6F26dvjbS57uCq725QFx8h52F2L7FZbXdA/7EZV
84ZoqXezzlLKeC/UlkGxjeGX5PZPmfSNux++CUY/d1EJuR862Vt+rtTHW5ifmqpK
BXvkqBokijGWZzjVePHqUxpdTJAN6P+izGScZ5lUHZ8a6UK0oMeDRXmQSAJHRuAR
rgsBw6QLkRwgyYPuY5JdnavZMautrzxUxf913ZoY9x12cRmhDx09aaTG/KgGhfEK
+RpGFxRzEUC/qgQc/82sYmH4iWfNiggNV42Lz6P+cSTxnlRWfFhycSZRe0AwrrR/
72Bfv0ZZLXhcKGstyh+x83pzLwhzpXeuFEIKncQv+r1Z/QUgcSVWCRxUf2A3407P
7qz/BOGzJXFtXS6tJpLTwjgo5SN/gWeHX7DQWSQRQp71/7+wdVB5J4qSNmwkkNfD
+5FZrJBCZD3urgvsUCAODrgThrrxPkLj4DWYnX3xNme+2y6JJVD9HlMlMsb7ez9t
4A+jGnmQyLG3eXrefIbIu0lSY/T8YupE8YWsdwGqjKxoWejRClhbHPtFQx8f7l6V
C91S64GhvTZd3DE/ZgyQYKBVgIgoPNs09SpYpkjAytM+qetEI3/No05UWJw+5j95
rqSenlcEjqLLHdn6x433xIza1HIZRj2MpZptGfbgZR/8ttVdc9fCt5w+0k4Gn56y
a7JOj8l/i9yUcFlgD18Y8z/EFddECU3oxNVhDQTWgESfVqM6B/3+cWoHTVtH2KVA
VgllJ9xhEf0SaEx51XoOcddke2FdHdCJd91O4Vzb5vY3ZrLwSL7Euy/2ldZJF3bA
PaP8QvuIFNapfAjxEpSBPFl9mK3OpEt9ZMYXhBj5DUM=
`protect END_PROTECTED
