`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cAzbYgIAae4c6wkNqlDDF/9+eyv4oYYWFIm8SeBieng2mOzXiyZLs/HuNyEUTLFp
28Ind7JSwcz8XxAGolHkigGQVYEufAJ1VUNKuYvNqmxGowP5oYWmD/NheC4SQABI
jyrtsNORghwUK0TSiQKgY5HkIoYOrkc/Vev+jxKNXh5Cn04R2+xXqJauUNkL38jI
wDOna7eVW0++VOqhaOeSqLk+bBP5GN/Q4JShzb5/iMHbOloqCifwl/Syi7vw0plS
ZLBxCDI2mG+XbB8fEPFX3kS+bpQTU0SLwRkhIiUyCqb42qJn2h4i0FKdVtOhqge/
`protect END_PROTECTED
