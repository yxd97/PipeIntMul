`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ywL8zXbKj2Gy8G79x4yqidKHHBNAjuC0YK5a1jw2jWK1fdymyBKeCcZubZ8vWI4S
/x/p/v2FBXdVOrCxutkV1A+O1ubd2XZwPPB1rdXAtjX0AmVETWBS8bB0dFDWuIvV
1w+TVHhWCDpxDNCOPTUZxn9I6cNFvKkbw0XEIUkC7vOmQoCZtpMQy+dhBajc7q+J
JNqy4tFvYz2bBulD/zUbl3ovKHiENhnv/UEhK7kuOpYTz9mm3Y/kjKCEMDqC8/V5
CEzRYYi2IKyZ+5UGUQlwPqKSK0smlm5LxqluowP55BpgkKR5RwLP0ijL21xYqkN+
mcSNWXgpowysH6SVxHv7xLVto8f3WOC/Cy8Hr5rlkN3mRJyvK81Rq67XmoWxvGJz
iO3Jq9acdHP5G3xgcHjhZG26LCKhnqP10uJb+itaWF7eKGTZItVBQW3lBEYFC8In
`protect END_PROTECTED
