`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nWmOAZzFM54YGm+Y7szlzmwvLSK3LjGFAajR0ws73rGnSizjqoO2d/LmEAqJdPa5
S4IhjE6S2F1Lpa8XcR6EhB51mg6/XLaodGXdGMg1W8rjjfoszvxiole6O8h0P/62
8oAbhunwko0y8mYvlqRqnk+jei29t6pijjSfApam8K/ONfoHd8Mxl6dPBDeGESOA
E1SvKaDwsld5VP2XEsLz1jyYcaXlTJGEG64FSSu0kS23vPthJauKKcccWJ1tlc2S
nInLeshC8z1ESAjpOW9OBHWN4j+ddw+8hIgvVatYMHMQ7ztc8wyR3mVx0n3Rb4YP
Gn3UdIjDigttorV2/JFuKgZNAPdhQLDLz1yNyctTKozRXRCCKz8KVWJRWN9DPeYh
RCnIfEwJxO8IFG8sRKXKRkzYtCLjVwVM5ClBFVZAhWwHBlKjE6T6PoAd5JmsmgMk
UrS9sAhWljM5KOx0Y9VYpU3LMOzABc6NzNry9TMRXWzKzVVEGOX/Fuf/cF3VlHma
rmV/wjX4pfTW4IcsetJnDvoC/vevm8je4Kk7F01qYNuX3G3onVTpb5z37exJI9Da
vd/ZWp/0ww0znfdVVYhO9FvuLLQpOii2TGFbIjv/8ESJ6f9+apYwNunUwT8ySK8W
wjDOz+POagKJxcW7TcY6BFm9wFNdvLJqC6CnAQgBdU6UdoUIr96SpjBBaRkhpq3D
GokPbKGujdFj+XSj/OqdtiTQygOUXsll7HZ6TvdGgOapVIlJJbtoTnkWaboMpoMG
hu2viYE3467z4qg4+YjOXZeSy2dhtCRocUYlJX2kRfPB24FqXJHk7T09DcN5TtHY
8nXJof8GDY7osMKNljE8dEt2Wi/zmAUsfR2uRNeCyEYfkLaazDBRHQF/CyKgGUYH
lnkrFmpDGobinSISjDH6pw7d0ojUlassUqwgbL5tolYLK+U7sVp5HBLUdLn2cfnO
C2R8VObgzSr7RokEb4HntxZWr5R+hYicE64cSRabLCJhB6pkdOE/XrhcqvZxE6Dq
xkubzXknpQfYqSJ8tevXsaNdn8EcsAKPc4aU0BgBf6xpE3T/S+2guDhAu4SEGrAX
BdhbWMb30wSlBFFYRT8onAzJtQIbSdXqYGL0BJ8O7jy7J391099/yVSSCD/Xp2Zi
xMrVdOzS6HUO6Xq3pkwjwDpzMTj2OK08wheBDCWZf1Ir5GVZNfAyYnV1shPOgAW2
xmribC37WThvYtfhe/BBdz4nx4J6hK6SjVV7Cv7mDI3juQxO4jbPXuh3/XS5GEPB
r8vsufIPRipYlB+Sc4v8CBIkFmkDqUX2wEk3lhmaTYZY6Cz1nhAxOcorg7/lk4J7
r4EHLBUqZGAwBzw+WOKkxMOAbKoE1Bdqhz8nOxRGIBkjKOlewWkdvDXwQkYedidM
0F9LZs/Z9vCdhN0AFb5wDYzfhCc79m28UVP626SxWNz7cRpb+lCHFNg+357BVEyJ
t9xQm9KtebqnF8xMHAXk1stJtc3n9+mzxEJ/RknDvLk96o3S2nMCTH0lzNvFHY9A
4QIOBT/h+Trc9k42WI5jGrndTeEYoRt3YSoRhDdB7691cW0ByPwjI694VmGBfffB
npYIhvd+JKBwo3uEiqNJ1TXIXu1QzwwU8LPR9d+A/SgkbnJrB1lXBRnOikTW42L3
uOKsDp2aRU3jZO2LnbGmpg==
`protect END_PROTECTED
