`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
opjdEeu65DWxYgM2/adx2KOH34UilBtXQaiTz/IFEFW1xK2sVsCmqF/j/XPYTKI2
XHNReBv+BOFiHUQRXVjOCuomfJpW2Y6n34dbvQZxHJGPS488XVDYnT2jwB98jFPi
TPDKDxliU+Ii8QUlbL5kPSdahq0xVkfRNIx8A9bGkJMpMNCLYnn6n1/6KnFREvPS
KSAwXgxIDjWgdSNb3hCqhQJDjXRVGltXDLtfJKH6F6EdKC+i3Emb696BoXzzTNAR
TrKfwvJXz5yshB6XCPB/M9X/XtFMO3xE5SZTXYEE7dpAZiYhFT8OG1z1ZF9g4Fwr
Qho9DqGu5HF7QEZRGG/Y8emkHGqY1nVtyFJiKDCoDc9yXl+0BO5rVW7eqcrasezv
3tzq77skTrN6glq38I3CRC1uO6ctjOwDScB3xx6aEWby+dx053dc1FpktGSiizOv
Sybclu6TPl9YhLxFJYDkJKxZv9/0nbVKQ78yfJrlCS+MSqAfp4A+8NwBm+PlwtB1
ayjPpT2FiY8xIZf8W0AFMi18fJp87wZGn27kkyPbzdif4V0T+kWNSJP3ImSx1bSw
asCh2SgRfZqB/XvB6mVPGr+c8pbFvUdu/Bc6RVCSe6pdp+CwLqWQ8uOTb0aOHJ+2
rDbAq0QPMIYBYo+VLGXij+n1lA+ngShmuj8JGBusDgbqWTfrArbc2bgvfyRVj4ny
MIgcRv/FHDcJjDfSrAOFSh906nl+iB0GJ/BNP/P5NKigtkxJzQLu8buhdU3/qg6h
lyfx3IoE8TwEb5r3eqFkN4oWxn9VfC+OozGGqqU1SZO3o3VDoRtJybdPAIEMhuhW
LcssoWznxXfcnSXmQmlKJXS7GFaZmY0hVJ57Ao1hrtVwhySUQS10SML2voRPHSAS
2d2AT2CF2dqyiwqKe7UT7qYm749ASWmpezSl0TPDzEO8r+IDe1aN2aT+XwCVuuWu
mOqoE783BuiLYqKhsd+5Wez7WYPPEwIkXSudlYFNX8wteqKtJSQLLRUSl0F7z/eJ
dgJDdo8OLt0OY3ffqPzl7DJM5F1sZJ00+2pw2fYqmJpJfAqeUidH7NYCRPxnXDTZ
UMN1vAFkYC4vhQZQBljtqf32SpyzO/cwjEsZ9/i70DcMTHSGBJBiNllU4C8V46Ke
PZVXAqFrJdYT8MPZ0rqtcKrK3ThDPR0VKsdYNTThx8u9vWx5iLJ3fn7ntT9N/0HT
eDTxjJC4kWyJ5u5/LXmHY5NPInya/sD6ikGIQEfMhcz3PMbkil8Hy3Nam3gdpGNw
ta0FkX2TmK5gOyqq0XXb43ayoe2bwVAsevTH6jE9d+Awy/hwNZoDGAeILZXwQBqe
d54u/P8ZRidrQDZOtYvPn92p+rGs2Ng028/5C3dLFyO4ewkFNRQROVBPSP0y0zTJ
8l7qCY47AYyhk+hdFuZLZDoBsOpuAewWoeaxq+qGOtTd7cKoHlpw098BFPwBACIw
Hk1l7J8ueim/BfEBrhHEmHf2JQA/MshBx/0nkwpU+CHDHIg0mFdyOhhVmfIwjtL3
wKj38p1Xhwmu93FZWPccXtl1NN0MK8KxG5kD1Y9JZUMAMCMlBMeG+gCEkBxSzTic
aKF5hctzTUmpopTUgSXwhSfM2IaMM/wuEHg8QcUpjzPq+QIBhVPpHP5kUdEQRxvN
Rklfu2yjwliL1i2C4W4SRLqnqszJvjS9aXEcOoOWIinDBUhquXs1+AZm7RkE2Rz2
x55m2+eEdcBAI8RwnZ60captVjHHmwDaBRDj8qVofzrPfbKkPxSTANJcmxW0dRi9
HW4ChJX5XPX62i+9jL4HEmwldQg/CN4B0YDZhBnc6SQVy1NfFaAYzsm6yB3FDpDR
jLVmHcpU05Rqkq6AYopjf2A4nHiIZhDNyZGT04bbeeuW0FcyByzhORzc9zCp44vQ
EL10IwYKhPY0lCXwlwyeh6VDy9VsCG7FSQ9gvR3u8G5B5C9iIeUtxSDCBlsDPS9h
RoUzG5yqBvl9dXzNufEP0KRHbYNDn+BNNUhMC6HRvXthvRZUDZCdmzOniFsH+u0A
O9QEiDdsDrlzb0XEhoAyFLgpem/mZysuLXn+2ivisHB6x8RrWNsaJU1YzulyLnNW
E4gu/CTWzFnJ5T3qwyHHy9aUZd2oO0BvBKnjFiE1OsI4OwzoPZeN4EObYLL1AY6/
DmEtgDGNFUA0c7B41glLd3kI3Woz4GJSOMmZQ3c7W1bzyG4aV60TRcVcL2EIggHR
4rkiomuG56AfRsMvXeY5uAqa6TETPXoJSIqzifv7EFWTK24M2BFpzGSz5xoFaO14
TJVHBEEhyv+IT/25d0RWV9YlSpeL7IhF7p1neffOx6NPnt6RIzPbhK3CP92YeUfX
bVd/ALljF5aQNAHXy3IBSVZkOEvjCCezdQP4pkXfW/yeDmlLkeQ9fEe3LVDWy8vJ
vwn+9n/moJMyHZT56eY/cJiECNAjj5u0VIuU1Hj2unjAmGvmY0L4a9UMMbMqLb1Q
yFwR7XpJI+gzN/rjmqjJcztRcJAw4yyfz2Xx2qqhIRSEZlA0CWIZQrS/vHO30s1N
w912yenc0+IGcr79SDlKV6ZZfM2UHrpKv4foeXv6qEvwzxT2unw9jv7WhBtSRTlh
GHYYx42wGESGEIt2Bdc0bHXTlQEwsf1gajeLp1ojU0yLcu8/66p/6XMkPKpcXWis
UxW1l9/ybuB0h7AEl5EEMpPjXDPaKd1z6ZRg64nL4Pp6UDXi6ddV570eHG7OwgLv
aCsj2BXH3OHpqN+03O+UT04ORHv3+AcWvklT3NRhQ/+WtMH41+tnTMgxj3ZgF07r
1R/HIGca3Vsbk/C2pX5wLmMjxU5U0PJWpbJlKsuCpMGrB9MTbBillFJlld7lYKvh
xy03zQEB+5CFThmwtQdEKJs2KDlp85AhMbsRdl0/Ao24vROCUpT0f5qZQgCNQPZA
3ShOSxW2Zhye15poSiF9iCWLuSGvUsOZIPzbvgfSBkmk4+dqrJ4sAzcMLdEwb3TD
Vqv6Liv7CQD15XzAb1QMxdG95BFjxhsFSrYticOBH5OqXC2ifKFYkosOGac3cCvl
5p5RvckQeJFXRmlzjBUs398S4dVj26EsXFybAGhVtvQjpt36OcICYXm0FNgr2ft7
71wH0UND6J5B1GNyuD0JY6NEtEsvrqOe3GUbkP1WUydATU5lXX3XmrZ9AUZ3fGYr
ucDPGxzWydtcO/ii94RSzpAUUBp6w7g7l0fwkGkI5Lm1gei2VYZXwLP1iucW52nt
ux+ucRiAURFJgW/LOiOLNKh8RuGx7VhZzuri7crbliF8TAhwJoF1WH1w+CxvSeCi
gFsTYAmS+rSnXgqYVSMB4txBKVa2Dle6DvoXJ03f8LrFkeWUL20P0uAP42/nqXCO
Du/Lx6Fp5dWd4sv2O1VurN8/zq35DIL1jld88oTKPO4V6UyxUEiNt7zZxcxBWBLy
Mrkdl9yb+4/lBM2vMu3DHLc4iZ1bBceNvErF3DQksohLPUtUEsbKjGQTtVzP/r6z
DRm5/YVe6bW6rvnc3FuZ5IJE96Cj5yp0a/K2EZpreA2s3pUnzcIEMXD4Ow468Vct
W/SOxuGRcDbc7hGndUIH/O5tUH4FHDxzbZnoM/1HK1HAcwg0FTLSa6LI4usHFCvV
uXLghzadZpQDjuyF49691LSMusPHxnuRhhwsE09Hgl9b6y5HLj63f+J5KAtw5RGj
41fJbDI+5vuQZOAmNkXRMkS7yuYstdmaOkN862rWidG0MAADayjxMAO4yaQ5aLnZ
HxEAMPxDG+ddAxo/1NbHOx7Ooo2+NisGxCfNWyQsv+plRehtt0SvHtlwO7pudySi
uN/Ovfwhn6oLwCnP/OM9eMZuTWrOt3B/70x9KBZdJyVvFxiCtfNaUH6OUgcuAAb9
vHVlrf3llEcVYX+HJu0alnGy+5K38ba4KELbbWYnGsWnCHL7OaOzgMNEdImK8x8U
ULqhEkJERWJcExwdF27ffgyr9NL4/MiKx8pMgF1T6LpS2MwKqWgYovcZL1R4Z4Jz
HnwyYcyY7yuDShv/U0i9yBnIVOJZrZXtg95UHUMyyaYJ6mZ2BykXetH3KswEo3Tt
PeNM0/T1FcqQQqjXRu3a7qwVTYrPjY0wtPwny0BQkHj4v63g5om8YVyn5K8K2LM0
Lwd5Q5ArU8J7e/nkQduSpEkVyc8jdT5qy8Oq3rDv2u/uFQnuYyRFDPM35mDUmgbx
QhN6W/dVOy6sKpo5PuJKLe91vTShpX5m8H6eYl8ejp4JKGVQvXGqJGXckzdjG5mB
xp/ouy0/qC3cur5/Pi5BdeH+T6CXU7gZSce44Wm5VB+5oslXtXpR9d0ICLxxSRkS
PvkjWNhTrQnMtjsqYLT0oenxNSGhWY+VwzIKWaMN7xDS5I6V49sF8stssSzUWH/7
hmXjSA4xRgxvBHFQw3nF39d/+q8OBYn7B3i0t+AGb66SJlxLJ3qCh9P2EkI6lndV
ygW2ZnMZ0Hjv4V7Lph+tYKGyp+t04LZIVNgvksRD2w0PZtsF5XoW8bC7pe4bbwda
i8+4p1u1HBomfKKtfCkXXQRi24Jvpn9BQ+lXhKykbQZ61k++hzDricZJH6Gr5TuT
+cfA/oDC930/LULEPQWMqsQwjw8qOkynMGtsQ9z0rUlSbrVGxdZ8ln3xdqBKna5B
u/Zwc7pkfTsG+aH4p9wCJ1rUnufx2heDZ4+FzkeJZ4Mmm0ig6iarnVGJ/11uBiqR
CrXpUfGRTutOHI9im2UE3mppLiVbKOzCEi4RMPVbb9bYCvFVBWtrVsUB1p/PNhjk
fmXIzIf4LI+GxkZmQQD3k3dxHsPrNEy5mW+Y1ElGnCZexFq2S08/aW1OIxS84zI8
+Wj6CzIlGEarmqy9BgwwpiWYO60pVRVuIu70FMyeIGiaTnVZOsSlcxfITzKqr2Hf
iO9Wov2qe0wYw33J5tQg4f8/ggGQK/+cV18Bxt4VsXRsbYSS7JcPdRoPSOtfdkSD
8ets5jELr3otteY6r5KoUhIGTJqjNRTSekmQrE/DdpMo8ii+zG6fe1UPrx6BPRTu
GCXSKBhMctuHTBr4TGB/go2vnkkL3rsb5MpvT3AI12/pHfmZapuordf3xUPzKs2W
EyYe44eq5SMS5fyJKc6nWFwC0GMbNJOZ0FaxME237WPT+ydgB5y/2QfBZhQJpKh+
N6jP5VzcpVU6mVCsMov63OngpZa7XcaRCJLPFQRVkSdwkD1VQdYXpXSxVXdqaeOi
Xy4sPmpcxt1a8i7F2p9Ndxvq/TOoopWYFzuYqQGPHLelyVlXjZuMLG0cLEWOy7hW
GP+ZwRVAeoWRBqH+/jFQykqthDR41A2I9b9XmovSJH1+eKkB0dsSm71TLrs4sjfK
WsAKGZmuT0qg1S4VriL9q903XP/rByTBHxxqQ68gTWmGTPqQRHNSOqRRhbPnsf9X
aKAizvdDdCXVzMSVOhXuRvhp6a/m/p9/Wrp16IsetpUbY9PLGRRVeZaucIircWFi
ACqmsJZ/zwMBu8SqhQVGX5ACI+ZbXqDavNsmMKKzC6bIPG/GAaHV58TzYAxgLnbT
rpqtMWYu7/oEEkQN07Vhrw29s38hBIlNeq3FS6wywLb35EMIo78UnClWGfRCha3S
CNThR9hV7jX8bx60QIdlEykpoezcN4PSEodEGZixYpAUXz7cJDZ5v2cvk53G1VAt
XVEdo/DK7ipoCG6TTmX7iaXH5Vk678Q79In/KJYG4aFpwmKpyGLUErfCznnjUn94
eapLU6r7zoWG2igt1vCfj+oAyAT5A7RFBK3Q5yl4zelFFDxz3Dfo3ioQyD2oaXmy
5kTwPoujgy64Z38O8wWeVbgl1YZag7FXJtO55reEEY8uHcGTqxawUV9TNbRXhStW
6F5s6pyONv8l1Sh/3Kt2XIZ0jZu0ZwB3RrT4BnHsyhMFR8/sz61kt5C8LXUggRG0
hbMOtreLD2x1sHcZ/BCc3yxKoVOgzsT7M0xoG2p9Vos2Pm879E2Cf8/gJhZVaqMH
2taqIWFGETITgIm5u0iPPPI9BofO+auTHfWGs1DUkv8kXXUnxF3E2WbU2yzLUl2Z
qTyjUPS6MbcGve1JXfwR0O5RqfEmMN49jOQDTac5A6Tt/Obptt7aa7S6Bbvi3Qm+
UxbNY5Ig4uMBMIpWAj0m8A5UO4z8+PkZG+45ctv1Qf4AQGC/pYZFOz+k7Tfhj+64
ohnfAmt3L0xOzNr/ZVQ4oQ3IBF8zGTV6z66ZrsKEHKusmOkcADJlqd4Ksw/PSq0z
NtS30lxc6kYk4ZDknxfuuAibsOMswIm8yyNsvulmeiJPcw981cmql9r9J8f9OJl6
9+jUwjCe/iQ7XwoTNdz4KdxPMZioCjVU7bq72gMcQgBuVK+EkbW2k9Znr5UFkUcG
XfcOcXkQomvBPmWHkzj7NaCIe8Hj6YgvQOETR8ur9GqXyCLYyPgUdCnvKftcjBb7
G7MHUBc1wuEI6hgmc13d0GgT2MU9l7DaburXM4wpW6SUGZLBK6K/MCOYAV6eJ1rF
vmYOpsYC9fSacUuYBjeJp+GL30wsN7dQoHqqiBzsI1QAmFeZbUMfG8qxEEYcyqz7
EVeGJ81XVphs/3CSHStvRGf9DYyUEC8o+LMpbdjFibpBaFvqTdyVGywRGy5AjtBt
coafIKN5MUnff0ocULuLgcTgOqRVLmz7LRYH/3Fi2u4+ryjOSEkNuiIWOsijJ64l
d/QZc9OjJ3z18qbFuXGY5GpmClAE8XTah2mBK8FnKp5sWnz6SeqQZidsAM9rkSA/
VMawMHgSl+TbV48s2zCnTrB5kpM5P9V9AHmTL+Tqf0RKTKOu82bHJBx4ZiAlsF3M
Vsr29iAI/RlnMIyA/0AFXtTZxG/R8Hn1VU6gfNgrnuuBOOg2CCL6Wu9VOpKerhdQ
ClgbymhJKcl9DeVPpYVDY16TxbtjO9u0RG2PBZtTRxK0qe6heViSgyr08DX9RYuo
UWh8qgSVvoIHkBcpZLdGh+H6Su5SX1qVePMP3GCFS147LypDFV/vPJryNkki7dHp
+MU5AMhumwzpgbvbdV/YoSWRTYhPnWqZxue/dICrHmspxj5grcSEOKAnSpjvfqyw
Dv5vbRiynohrBPrTuGSpMNaaw7fpDeFeHZaRZrJrz4fpC2pM0r99xP/Gj0o3jdzH
Ai5/neKdiSiyM+2rhyVuvDqcMZR+ZEFssBFgjSZB+ilZan7Rtx4BabvwHn2DkpQJ
p96SLux/hjvOUh46sPQ7+f9BwplqdGQbd/656amDuOZmx4aVSO31HepY3POVHUYF
Ahsg/77rnFN93XJYbIxrBMfg2bXshhyJLX8aW6GN9M6HLlfHs6LFMZqT1hgsyx+8
g1HYApP8Dt7lfwdTeOqsVNQcZev2H196xZtgdKJZ3JYnQqHCV3ETyzS8QOi4RYdy
KtbyLYNbeWtKVcD1JtyDVKfNUBUtgvONoNVDMH/0oi1uQ6PmsX0+g/gx58f4kAk5
UqWVUyqxQ54kR0AtU7VbL/Zr9wFUuuMo1L32K+HMzGF+jq8RdjP5OTZ+U/qqkons
8tjiWz/7uqqRwd7gO3tsBYlnEoiyyuQ/wsV08lYA9TNydGh5xHFVvF5DK9kvtRjg
xgTZG+d27eClqisG37U4nL97B35s4r6ZhGnwG3SdVITvXXf3vunKFVOZfVTQvJEm
6Q3QV2/Q7wk32f6h9PeVWQy2u+iBuNiVbku4ggXeggM5g/gHDzdgEra2PvwksVen
uI23YRSKRwI6HBOlbPG0mwQQvvRWfFeNw898aityXL2NOOLIgonq+m399jxmI7Gn
yqRMX79UQXL/j8mB447tfI2SfxgsWswe/oClFp6ELFR1kL6XFikrBk7UXq0Cm8Y3
kTPLO2eavaBBP8B2iC+Ty6hL4s4uc30zjsXlZgi1h1RDnPvTiu59qcqty7FuZj3m
FYPvljdLSg3BcMJm3o/apAjqXTquO+bTvsDajoQUbyyGq/T7aEOsdgoht1F1z2W4
9QHcrsOcjEtefb5by9BVKRVq3ujvdG6WX1CCa7hNZkyT4OJXl5YDMQywQ/9/Uxct
ONssTil6x4v+HChTrOn8TKfddF7Cmb5YIKLSF5lgoyXg8hSzAJJBETZzRA3iHV3M
Hqqk7bTx3tIVeh7Bld5NO5rUwAI82Pd2TKUWkn5gDA3dLo1OXOyPvPAFsJZw45Fx
P2WiXHEFB62b5MSnV3TtPUZz+EiZbKEqSaMroXdu3De4dWhldsat65dItBfkJ89+
5lBB4uXPkfGphFIgCbG2FDHgLSMN5x7AZtUVxOogbLCbp+GU5Sdvd0CDEBL+flcz
c4cvHO/lh2fIoOB2yM4GpXHcV6GPufspgIMDtG0xBYOlNmBkuw3d2hfoJPV/ln7+
5WnuxPAkTK88nNWLmoi/v8q1QQDx2XrFeVSV5+XeiQ5i1opYiUI71c4JStPbawM6
Q8dBmzsZs+LO5oSo0PZ15xzZ5eAtUsvi1MlAWq/6neE8yEG1vuAgm1wTlJhJgslB
`protect END_PROTECTED
