`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oN6jfHxASUOjlR3/phPnl3z9ogvvAZbp7hqhiqxG8XjWHAT1oiUucn6Qt4wcxY++
7U6PI1Vli7oDuBYYnraVyjCIUIPgtQ12+AJxgx1JBP94EahHm/1rdk8/iw3uKQsR
sfR2E+xJeCP37Quh0OfQSS6RamXb5pbNIr7iz002Tb23e8fHz8dxQSmejV/mLaU9
8PcI31TY5aRV9MxMJEl+LQD0bZF7SypwlRvJaEJaxvixDZQr51VAVNkcE194ajgd
`protect END_PROTECTED
