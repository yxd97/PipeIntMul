`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x5WhKDP82d6XM9MLVjKIPV6Akp3EWeIZi4YYdSy8+H+Kn3xEi3AbrFNwIgqN1q3z
8BLlEU8Xj2Ys0HHkwVZlgcLEDfcvReJMm29qDcBxaPR+YZusl9djjiutm4ZM+6/w
OfNtzLraq0fnl+VnjXhC9BvkoqTm39tPd2BK19LDs2z1ikIhWYdGgKYSG5GyeLM7
akTjRdDK6O/srelXiyBu0xbXp0D1GbkGi+j6T70GeSYy8tPTtc/v4m0+RHLH/pIC
WFwqCKrv7shNaaH0B+Uo6WSKwjTtISsa4+31DkY8Qi5liMvD1SopE6WE3DDoUTAd
hWc7jmn8IANMTOy+xkgGZtgWtWXGgYzCRc5KcvDvKlKBz3BbZgiLlhpYBD61rBE8
kyHE7fIJKohROa+fx4Ztsw==
`protect END_PROTECTED
