`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuzNHeK0c4p2Z6QHw4woaICltBCPaONjWIfmrnVyxmraG7aAV0J0WV33ycpsorN/
sPub43EVrzStLZdZyuV3JrPjmee8kqkEORT1M9XsZ75QefszsUyyWRQ6XEzVIZvP
O3JDDrkFO4YKqueaFW4bfaW2E7Qd182HBZH1+rmeiITbGYZ1rXuBULkTTHswNGXv
v4E1SgT5eBdFnoiGSRx/JRhty1sDAJd3y5PiHuZt0NIm1EjcclH3V4pFGmHvDxsv
WWNUTYvuGxn09qjygPfwty6fop/pq1ygRpB7Fi9ocXCncvlS/EdwEUGCeiElecap
MKz3x/WGjBFMWOlN+tcxUJEkgP5uedDnkhJ6J+LpriDQrO40VUcJwXTfa53WLqk7
C/tDk9OV9y6SllkkwNPBn2DK/yQ4usKr4vFCmUt4J0Jt/uo6HJbre/DovCywy/pa
fVr2iV40cLAgNB3jeiv6u/y9YvogPmi0Rjoi4VXEkKLJxkD0+XbgpbUcIdte1I0X
s875yKYmEp2x0bhi4mUNAnKCoSZlr3D4+D/BIgDMi0FSjw7Z67bt/Um3ItzA8HSn
i4vtr5yZF2wRuBIHn78FZ5xd5tQKFiyKxaf92CatcYlgjJVnIh/qxf75d88KOVqn
mv/rbX+qUh/JmDA4jTbsP/VSJZ/5cx7vAhDYn07IuR3ylu5w/aXRCl8gO7hmxHNj
QdmIUVyqMrtAUW0vd6LixIHFVqkkZaB6Wqs6NW2660npMmtPX0zrxiocHQzaHvFu
mjMLUcqTbmQJU4mG5kyLCutI7CSIRZAUE+e2+A/nZTvwr1aZDcj1ESqhrd+Cg3/W
//U67CaMg9iqjeIFot4HgYatJ7BhU0NghUb3VXYK6sXafwZGnZmHIR+nmdL40M3c
wsYVpcMc3z0RXEPw5DlVm6R3WmCAPj7Ms4C1pJOnWldXlGGsu6yTQPylF0KJPNgo
SeCeUWIOBkBn4Msns6SYPWVif71i9C5/DuBowTHH0FgbXnMnxn4dkDqINvgyXkse
RUlfbHCNVdhri3Wbv94VQay7qkq6HOROw2M5hq3UIJ1fLFJdXcQkAtmM/fa5k663
Kz9Q+Ha5l5hhSs0xs8mcR35AMaZ2fC7ol5UPfZf0eiNFAkAjeVAeARf3MYJbkkhW
FEJQoowhRFkga3Rqu/FNFNKu4HN+4XhFBbJXanNCqR1Hw6i0Zq45zYx69yF5R5Ls
mrBBUH1AokDza617PSmuRndRuI3nYYnc0Od+d497AF9b1LITF9cMymDiMZva+KzO
Ar2v1W4y8x+Q2p+m3XgdDnEjMAbzuMv96nBf37qfttTm67UmZcyx7L5KV7fOMaie
LQUopNBwVSn7mbwFGezCwblbJMFbpQayiutZAdsBv2AvinmTC5sH41Lth1/2pb14
klvjpPPTUjYd3Yqu4iOGFeZlEFH/1ynnionOndOap1fCAnJ/PxPN8vdz3th8ngwU
OgiWDDgWn6Nr8W7Npq8zWA==
`protect END_PROTECTED
