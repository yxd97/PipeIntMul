`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qaJ2YW1xMoJzMRTZURNqj/lCB450ImQVt0Ju5KawjPpfpotwVFoMqdhkYn6bxq2M
oMA5RIoHRbfkxNvy2knl/wvmhG0ytwpopf8uhqmcKsX7dTpWXEHpeBsKkIOQuuBj
7ggPzo6FRWTfAUUCdj0kSnrtYYEvb5b8FnkkECLT+xcOfOMDsCNmnUvXdvsAfLWf
Axo2KohVdUhoov4/V9AGEHRu21dOkn7TRww8jqTxS1MPdIHmsjq7nwf48JBLUEEc
sYTF7+ArLErwcQ+U7r8KoNdZ5evSA9vJ996vld+16kQ=
`protect END_PROTECTED
