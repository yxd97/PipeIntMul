`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+r+E/OMYkAHb+EBt1iF4e2ISrGhxalWKH4mR4pXagITeWMurgb4tSnBU/eq9tH3
j885rQgY6oU4R9Fq3NF0ghhYpCfgMD5ssDEg0WfmSX4knf8XoacLIb/WV4uW7eVL
pl3+DI3YngMgdC9AFCqtN7EHqFRCLFOHNBdB5tiujrlk+Nr+OKkFXEzPp1GtwtM8
rw9uLry2y/rxOVJWF1CPO9PkShxs5CgYye3xeqKT+UUF5CbP1IFLGN41+fRdD8K2
Q/bPrXhQp6n7BCiQ4WuksAC8dJtc1SeC3TUi2exMY7CIrHvsUtMDRHoM0nBYdsGK
uBILRKRDGpBb5Pb7tcMNtg==
`protect END_PROTECTED
