`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiLS+ZuG71MAnt4B4mT++gZEXJlBeYNUklgV1NW3P7GPKyPlkST9s2R3x9BH6dx/
cZWT2T6PWlS59fwS/vnc97mnAvDT5Dn1V44+Mu9VXLGRKfeMtHYlZXyHQA66jjZ9
mcEvi47RF2Qfy6zc8mvEL+X3jDdDpf67UqsUbt3NYp1MHJaN4KdNJ7N8YmjUEZSB
1J0odhve1VcLNlgfQxdVbYQrjmO4PPX9F2i3NAIp/dr+AfEnyNk5/OGNZmo32OWv
UWq0dG+GGQ3Fca02n8a69DEWJ5VWuEJPOh6gLAvw4jzbUTReJqN/w41nePK8tZ2I
LZApttNt/xGNy/xf4Lg4TVc+377p+JatRfQNzBneWyGxHzdZUPAK2sG2WZVVtf3O
eMOE1/fSig0416zd7gYHLcgLKK/MsEkAoieaRV/3nBcU0REc/d9u+F9uuZgYn2MC
m9cqGwNmVbG54x/HKLJUXMdeUdc8WUbTnTepoxBOs/6XvfVgrPL9ysbg4Vrav/bZ
a/+GKRL/+64zRvonN5/S+VvCXeCO3piO/jCu5OfC/hvOuL4eUWA6C/CIK7mFYkiA
etSoIE/AVEG4LgrKvTlHlnwn+WkC6NTu5mjllYtws3E=
`protect END_PROTECTED
