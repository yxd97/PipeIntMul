`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCNfyBOba4hu9CXuy/V0dd7YHMkPcp3lspgYtTUjP6+0C88o5Der8uPl6eBiEOeY
EiACp+Dmh+BMzud+iR+LbmskQKmdva4fnUD6+mABFXuwEjL7HdbDc/qMVjI4fYu2
KA9eFCGoGiJyMv3dUu3dY27UJVL9V/kILu3PCekrL5fozJ9+7Zkcm/v89kVUVRzN
YKaDC45bvP/LjQhtSYxw8FzPUtdZjQsGcI7HbgdiM0Ks7fukvwACfDU40xkHpaCE
ZfcTNH7Mly9y3aY5QgPhAIdycQzwnIFv99jNxJKeWk1MMVdgcN4DldB/Y+1xE+c/
0vThtEfLfH/OIJkZq2CD8/Jsv+IbrRj0IDy3QQRiUt3U6dLxlQDchHp774L5URpJ
83lDqftV4CVfDU6kHahBR27PVMEfVCM9RnScrAf7RoQSza75uXL/IwqUfj9p0+U5
5BAoWsaxBpv4AZyzNFDfewQ8rWk/OGNW6Hyo+vahBm3zX3kH8ZtqzNURiij+mDsd
JFlG52LL/iimR5k3WTsEZqiCOTCSfBc1IRLuh2llCfLnuJfPAUQi8vVl9Tf/Kt1e
oii6GJMYtuZ/4ftcscbVuJ5+Js0TFRmwc9LLj7KygLI=
`protect END_PROTECTED
