`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7wLGKI8FigGy6WQJ0Hfvc1hWzgmDqXAE5xb+yon2kcQH69C57Hf5uqWIHksVOxgE
MF2muX5FiV1zNB5FVjxkECitHIVY8zAiVuLtZiXy1XUd0q3l5ysjHDYsyxkHzpWX
YKj98YZE6Q9yMtRH3QIgDUjAm8dtvUoLbyDlF961LPYUA8eWPKMPqJNxAlM2g35K
Az72pf7hTdMUn/C+kl47DGr1/YmTAsLOI4xAZhjg+Wz0xiwCiAjT9HjWJkRII7pN
2ouMM8vaRbLS7O9vqkXj7B24ANUOEGgwnLM29k7xljE/d8HduTUc857kjz+BKZzN
6aBV75fP/EcBRWndKaPBdmvtqjZXR8md2C8cvUFUoUQGADHF3a9m0sur34U8ROc/
5SEWf7SGtYYHYmfB6mXuwmf2jwBW6FVhjNc87Uk5gIxC2pLaqwQjnaWpIIclHJKh
Igcc7PuI8jQ2koJCdohlWBnWbeeaKWe/heouXGYXI3QUm+u18+D7v3DhmkrHV4Fz
H+8b/s6qsWerYkL/D9PPrwMLLTXWKbW8KUKJVEmyECr3RQjJ3EOdJeyD27OTXiWY
a/miOr9JIxbNRz1JTPYe8pAnhY1kErjvTYuMqb60atb2zOMc2ThSOeFXcosm8rdQ
v3XSrqcL/pcSdfb5vA+3cseZAjHR8LQu3VT1tYcKgawZAmp/IxsoAuipgML/Hxjj
pHetZRGvLPCOVvsdLcCYtOC03TUwnuCCI+0OUqQYef+C/am1S+uKi1R/QaZirLu/
/H9lSHaXcQmMLb9KvR5fnjzIeehpTjX64GuXqjybbatyHJa9ReBliXMN4IVscKo+
kMV3y0zPXPK9ULIuPt+bj2EZqDa7JtWmW0pQq7gD3+sa+sVthz5Ftb8B9xpDdcGi
`protect END_PROTECTED
