`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MdPnTx6yP/yEI12fpYqx4M8l9V28ZxydU+V4abI8LWm4m38SFBQGBOaFnRP9SX7
f8c1nlQVoyMdPQZTyBCqIQr4pdv7+ROcGGB1nfk5L/QQ1uRDOXmyUKGfgoxdLr9x
mTwT4LZZKml1fw00PYuPXqa1eWzSuRdcXwW9gMA2ScNn8XfPdqV/eDK+eEgK3YMi
F43xHxAQTwGW86zWzYzIkV0qnk1HgSR7zVpkP+iN2Ewp9Z6FcLST9HLeMXeHF7Pq
1uxisG0GzhDDHm+M6U4xOhQJ7sELP1H3FGaC7BrijJlplITulvhSN21AgMY9auvt
KoiPSiUfCMEnaJxPeT9ZKKGo4Pku2dCaM+Xvw6xu8v08LgVGadnsPWqfJzl1oW5C
J7y2k1ry10iEeMvi89MAj4jHfVH/4cd4pG7hyNdFZ+gg/P89gziqq71gIejLh1AK
WPrWxJSJvI6oq0qxX3WwZgzkfUUIcC/mJS39jbpvoMg=
`protect END_PROTECTED
