`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkdC/4nPo4UuVuxZOOzQodCzm1n3qOA95DThVQCpEbjFXW49+pLqOg1jXmi7zSe/
d3LOz/IH5rhW3ZymjEw6bacvEjKcStSmm/hBKFuqCxR+5bmUtZJq/Gzn307/upRq
Vi4N6kL/Lt8EbxxrNNIyyI11/6MMeap1IRzVpP69HP4Iws2aEN2Sx7EMzC3HgONV
sYEHUc00YXHvEhzPMKRxjtEawNewNtuika5M0Mq7iL54qJUXHcEbaYuitobYqRxq
e/laRq6vsoteXQUEhtN3nlG/EOx37iSVpG2pAZW1aUGF2u7OPn0aO5KHumX8YkbH
46lk4eXM8sivHAEwciUBkLUkN0iqQm2/K/QFTyBddn1QtOuQkX2jDgVhlsZnLi7C
JnV9UjIyNRZy0pB9kJv58fdokCIg52HpLsxA3E3SR5BPhRt8lEGz2sTi89pC0jja
qiVjizqAS7SfgMX7UubO28gOASZIAw3rPaDjUTfAaBFjCL376D955AV4skPQm9rR
`protect END_PROTECTED
