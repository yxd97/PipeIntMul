`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G1aFztugz85uWf3xlR3OWr4pfGio5ckinGokWk6pNvHGglNnApEcU6LApqEj4Kel
321jtCcVFWl+Kt9uLzAYq5lhu2C3SpAJ3qtWZnLvUdWTGNUkZp8rBxwGItpA+66H
6Q0fY1YG0XUjYa4F1x5sbpt/jpJMlHmQEKVs4tUVD/lw/A+p6hUwKer+soe8DBJA
3ztQLfU0wqg0nRluv4ozii+ur9PLWhrzYw5jGgnNlFw5htW1NC8THIe97jKiIvxi
m0BkaNDhDyvkuO8cJ5UBsJR768t47kIwE/WPYsUmkeUMRU4w6o6y8Pju8h8beUPC
WGpdOzuRRuXPHcljMM17kWG/tL9ZV4z4DRhH41Dq42lYfIPS/hAudsurTalmSpgn
v8AXgstpPQLqH7H/IBMzBnNcZaG0oPO3jU/nukzxl1VJ/nqwXfDrx73rqo17Xglt
wiZG5HWdOQsQixKj7jhbzAmFRPjCNzSPCl2ndpRKcD5DnWcPyf1Rw2co1DqkupHr
ib5fey3YT935RHiQu+AXdyljuuAr9OZNitn2oBvnw0hAxva6tofM+wpBaRJnBrVq
6xHADYbQRzrC79PI7LUipE27ysosoY7Xu7I7z23pHMhL/FiwgQKOUf1WBepS/U6i
ijjxhOegbA9vq92Hb+ihZin0+aEavEKSnleS6kfiQ4A=
`protect END_PROTECTED
