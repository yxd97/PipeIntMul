`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qZz/+4xidPUsc0ZFwOJXzDor+hAIWWc7fre4EuJeC7MzePFvghJkLmxpFv7tfs+R
h3rB3patvtrDTGzShGaEtPlGkXKMS7ecTle+W60hIi6sXXbl+7ZFO5M7XUzY1lSy
EdmbEOWengh8uEtrlB+QjharIN9H207AL/cieSSBLKAQLuf42YrrYT+MWhEcfMiA
9yQvHb1U8Hui92inHYE/if4oAxeUquBYphLcIn+wT+DRPA5x3qpuLdEmCZlfvOcs
mZYEIkipEHhiBWtknfsvnWo6K3qQ0y9s0m4Q3yShdMv1T0IgO6u3eMlt1aBSPrqj
EZX4UmQ3qb9BTYGy5duerLGnxHyOsXYaz/eQR0f7kxzbvYUKPxpggDh6l5eW1z5V
LufUfcYFVS9SS/OrsWDJ33IqhWxH6UY/hkMgTcfVvTo9BV0IGq/WSazszamaYuq1
EJlCqI4a180ZSDBNXsVNUDWYSfGsjlkmKd0jGYJ6kGD3BLWmR07a1XsluKZGW2jD
OGgZS3/FvMg4xYOC5Z9zurPityob8sSmkvuzRi+7/4EHb0b9EHnR5pWJfTX7f+ex
9JHl2rBPDUCczIQvKWiMsA6HsiRz/ZYQe7P1ekpyd6i30F6Nl8dBqaw3ihy7NoCs
K83ANIyrwFZ8kxiUfNcfOYbyJHgA519pEjVs6CK7NvpprBsL1XUHOrRwWWWpWiZt
eXNtvOzVcu/NlQNrzLC2zQ==
`protect END_PROTECTED
