`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmRc4REHw1k3k5PK1u1w57MtPt5yDfxJXYy5E2WkKR5Odf1GmUZlG69EeLZez2fR
zDrHANTx821awkNO6Zchcy4bTeOqDgesieMoT289WJFXh//CwLIa5HWnrLzm9khP
WtcSSqvwBciyHE5gneOpK36ICwUT7i+bBMzI//iKgyvp9wOs7OW1PCUqHGtV+jCh
D9cSR/XIWft0NrnSgZfnYi92UWooMQlgPZgzIVbo0HP3onQDPztOz6Tt5nmQP3in
98b4OChfqkmlIYTtPYA+42csq2GHg748zmV365y9W0M0R8R1atfpOqlDmYFC1QLf
oLGa6CQZik8fWBB4VRd7lmQnOBGuy0uOJc/bGjre7BhLiyvWT2lfmmO2vu4xN8QL
AV2u7HxR34TvMURUZp0OhHaDUN+LA7Ypn8k/LofykI3NGJvLvd8W6wzpIIi1BprC
Ed6CnEq5KK269yIGD62wVT1Zd57NjKkOpUXg39y8mko4vptvSn+3p/Nx5zyRv+Ue
NF/94M5HT/NGyJWDpSEWaNaB6o/E/gIkFDU+tSh/Lod+XZkArjFzV8RoQOswZXST
M+kQO/wStpuanbPt9tWjg8KxHRebGUr5iBVBU+W2ba5W9mWU/0coR9KGzHoP2Evt
rginAqgEYXFNDPeo2g+ux50zJY180TzWZsmVDyhzn/X7FTs2XaghIIPxHfNkyVU0
nyTSaYBTHjqomAMoE8y9dfPqQMHNngV82vWC6V5iq46wvILA2v9cl3QAmlpWZ2IA
CZeOFo0TwrkWv+kKb6H5RKUHU8q7G5BSG3fxC9YaFDwlpvQvIwQJDZpnbugIXY9r
bndViVdYNk00FldEa4ChRpTOgoRkSFsI4ZdEOxBJnJY6KsOab0RSZVY5aXFstJT3
IlKB4QZ1TcZk/RmC0ThiblwI+ig9F8tDR5XW06uXXbgmjI01zJb8NRv8Aai6tkxY
PsspXJq39Jr8QT/GcAxhADHcuNGt2+72RIvPl5xeJvnsmtP0ceAg9pTZhi9fD1k8
i/A+IyDBP8CA/0QYWUO/Ztm+VQZQF7yanBHt+qqXOtmNZZ2XlC2a6UH6839HiN12
m6OpyvN35bTULfT3EcfOUw+rBb8PCWGYYyh5z09cDHItGyY1GVjI7wgg21aYxMEF
mq+QNDVrmSI+NmUPEyKe9nWvyVBfnFQpOoJ0vNCEVw7WrizIk8oRsRn6nXP0qCIk
wPTwUBofGJHnHGtNPRJMVGS78v/zRdT2DXgtSMClFs3KcsZ+2lOnBv9/HKeXjpr3
3Drjz3pAU/I7pDFvw6s8ItXM6KUJwFb6FKsOaQKloUyrYXF0tOcwVkFbbYlrdvfB
jm70J6oEAKHeM8WDN2Yxgt81jBVY/zhSTFjS7IgTIX8NBsM9ZBSQGRfZ1yYbSOMJ
BbAowAJ+SBdbJyjOb0YIVFZbYAADuod7555zVrk6MSlM2nCrP2Cu0HX0BJJqcXFo
vS/i9RcYfsVHPpgMPJu4IhTMYiESh1ZqZ2Kt14tVaDDq3NsAYYX6nvhg5PeTxJAY
bsFB0ozUoL3uaAljdwPK057re2+lIh0MNzIWjxpkAckte6Q70jQVF99TbkcYaJOQ
wXzjAxy7I/yVYWA7xGwobAYeJScnQTUqHAoLrNfTEwWwC16ZuYdwbW/wGVnk7pr5
WY0bUMvdUqOPEEQfHmGJnoMeM/jY08zahMmfheY1YUC+J2l60QU/BBgBUNkZBJ61
mhiXGqV3l7uE1MyKS6V0mEkCCXMZaz7M2Ijjg72Q6SHx5YxhSs1ZTI89hFprzU6x
OjMwSXhIuxiqewZpIzqBVgccha7JuPhWu/mNq4jJv3qJn8PTUNr1bMJ54EZ8ChNe
Ql/WLINMrI1L6oZS2XukAOs1SpKY7Ohu2RO2vDP1M+ZGw/xzu9LAdlhcbdOXaoFs
XFP+kLd6aTZu3n0GHYX2Ipd0k2CfMj4EcL0b7uDJWXHkGS2Ga9cpBlp4s49nJDtf
C44Hx9EP8wh467u+daRZSh6NQmP8O5tI3dVLjzbrM3GThxzCE0Jl5OfVOJ5ArSA3
UsriRWKpJsotC4D3Kz7aCtBrHBIAxOMK5RkIA9JNX+KcWzwYvLtB/apQ18lUovxh
MnLO5kX9kUFoJbDobHXcsvOhY72nzvGwdL6Xy59RNjweVxwfLqJ6IhY5ISAOcRCv
NSFjeLzD7XnNoI8FzniOCzskhZgr7/fwF0fa91V1LYN09WPGre+6JcsFOTzf6FC+
8CVTjYMhlDuQe0P5my+PTaeam3FkXXU2iM2VY/SeUe31ASZ8lZR+DeEqvtv+KWJT
OCG6SY0SEx8GQHcGl5nMlAQ91f6sYaxMAwmcwh69X+4cucy4bAOFlJyKoZFx2vIk
Mbk/3adMkzWcTD22TgduD23tdbdSDCDRbB5+HQ5yosXfjyvxbRleMOt0+gIav3N8
RAkPALhpRjpwEUVmCP5bSrU2CkCrh4MA1Sbn+isKwlT4mecOI/dRhGdu5vtPQyxw
yo3JiOlMRFAY1t3d3W8jIIUMu7NB1LKHtZPwW87QjWC9epQJhbTXOOPpw6ciR7eZ
ZEqjmrt4LN3d4l9QBzQFsqjYs+mgaWgXhkWHXqAp4hpwtzJBL4BiyGVDKqitA+2m
c4FokFZEZsAi+MeMPb5oue7n6VaI7CDNkZO1HeLPyHtwl+/51+OCeWFhgK3d2Khq
gLtRnJcVm1tEBJrzSOZNvXA/HTbmAhyOulTqLTr2YMVZ2GRWtT26FGVJyihESOhO
24hW5R9SIsVsJ8LoW1QeNhR0sb2iqlI/TxwueEvpEz4ekeDMjwsbIhLRZPw4eWQk
9fWwUik0dNQdXQURnyaMSdfNPnXTXQsxc41tkHD6+xJP3LlGXmS19aNk1t/vCkIa
pnxELLQrbQGYJRJJ7jTAbrEiZ2D1Aym4FetalfWnt79eJ/apSrzqs4jz/AIVfIVB
YhzVWVEL6+0xNNzhg5RA6XmDTScSUM6y2kKZGZbZuJHgf9hVklyJy4GBIyVvZBdR
uwFAOYEfDwqxjONa6ankwMm/AC06Lpla7bkRVoBDA/I3ChK8uZnWQO2UU4ZR2yDG
yFju+XdSYJKGqrbcJMp9fwOix/z4ZX9QNdrWewri0H7EJ2Na95wahqFnqvLk/ZNv
rMdD22s5KtQYJoohi985R4+6xAblVW9IQB6XIewYouhHoTrtoNeRWZWzg6j71heH
gwiEo/ueIjS+woCfdd4G5M4vM71pnjmpYQ9jVP8kdvNepQFBwN01LDBDABFguHBm
sA5basr1d/f5YA5pTONPxUd/29Ktm/m2jjmFE/HQbRUvQRACCY/spgrXnedaqfl7
ECkdHGn4qdVj0Ij19mwmnlVSj+MH5MfxcKBkoTEP3eJPgPfcNm+ZM8AaoQE+yNGL
QHkIWPuvZubDLrH0PW0ugqGBtUrTJWJSlWA4rRE1EC0VIdjaQqNEzaEUFBR/f79f
7df1ApPm5es+MrYeEuqPMk+EKaYCr0QFcvJKZMbJb1ZRQKuJDUQeBdyNrL8Qauqo
CLVhL5DarWMxESMKNWmQOICnQf90RYTcbgdEMgLr7SZdm2b8SpkKtBxY2dveilDx
k6JdgtPKtKZvb6SqcwSzVoOovHEhM+B+dvk+lz1FDxU5AS9afMgdSzaLq0XDOViu
1VkkJSX6k+95BDHj0pI9K7cMK6rsd0L6Y7+NZkMGTARol0pKgMcawuA+MYvmVvDX
p/HoJ+QtbNiuoyd5L9bjusH6lpNErBj3LuMTWvTKNwtIcgXQHZKDQafNzhs+NQL6
UTxZsg8Maj10XLz1PaH8gU1sUwdnPI2uSFpYceQDtZtdu9lZ/E9D5Wyzb1EDJWAG
G4X+suqvp7FIP3qnAxOsnsecVlgl9nwrSh6qVvdDS+376sfsbMzqARwIaC4DWWdN
yAUUuFcSn2sGtpwrowBiCoBA9zXkAA7hrjksxC977YBEM7WKzxYrzMGQ5BsEyOk2
6mbaq0cJRT1JA4Y/kBWZeIM3ecTedZi2OaojZU09xWQEJBZhvJnoX7AscgKMEUTf
H2Q+xlrDk/aYdFdkufPX8dcgJTh+bUOWfJGA2wuvUOEDLo8g8fZPH73ERE9OA2rM
Vx5n2nTmRUvju9niZUW5bFv8MvG2ELidi5RRNIChiXDuP7ETIqqTQnEqju1nU6rS
9otigHW0x+3m87UlC9Y2ApCUngj7lY33jl20EPZU28PB8TJ51qz/RZyos+fYo/IX
AftT3Sdn4SLC8MU7qbPDWuiTnoFZdHRqThUHz/uFKqHw9kghSQobY61yrgUBpv2/
Pc/izn03iW21oDOWaaOGudkuNM154wR/LGDOpZffqbkwe4EdNiznEm8a3mBdmn1s
klmB9S0yHcoXQk/XtzCqj9YJh4uJLslIXNmJZpNCu8Ibl+9X/SzUqjf7waUwRZK4
L9WGzn+Cd40n2K6//6HMBGn8eHhvnpO4Kvw2+TmBOwYO0pZgUWda5Udp65Qz8u+e
8xxTBD6O0x4ZqySEy/A2nNQP1br6dsgpnktrgqnbpLk+BqieS4og4vRiVDGaoTzV
EViOF/peTmFxX8MQwmY1a7R7PXxza6NWRGEOIIg03isFCZgye6/cK/FJN/JIXDe9
5i0H5Hrg+CY+De4lJ2uVLQhr6Umm/wD08cku3sSY1vUl/irm+KuwvyxsrCTvYov1
qkofljcdEKgcCvDlsdtMMAiodwlOfCgeNEMj9oVKDYTOvdhKpyt6N6nMmRDgkAJD
bAiDLdcM7XRHsUajMvsOsHPIqvRV8Iy0yxCW6+m50tSZTApHhbzoN5MHum4Ats6x
g/5iELm9LRLyyWJ8ac5oYWZ+TbrpVEomHJcvp9yOnSyJFBdKAhaLxySvwlwtvQru
4xDb9C+pa6kzdoB6j4VwX8Gp+H18DhsSFEAW7ew8cxb3m/K3ESTRt1I/f34uNcsM
it1nUDJeEBlzyHVHTcDud1TMDiyachauBhLIy/2uw0hNQWihpvtTcapT9dcZsqcL
ZoBPzmGubb2t4btkqtuxz6ENmmkyQJIU+BDxu2OlWIpt7tHAriCs77XQdsnVjKpG
u+fH2sjhcPPtHrMns6N14O36aVKN4EJ5dysq0czjicgb5bT6V0I1tAohuN5ydb54
9blqax5Gjar0znBjEZcHhipgOTWkrARHwgbRXKFLinZNIentFaVrh1v69RV9e/0G
FbAOcUbMeJEYY995Oq5IzTK7PLLutvWZsLUXkEoSfHMPUC/8505rOlhOt3dR1v8w
vCPOfi8dY/eW5pLrjkF9qL9n/dfq3XUqyLgD0pSugn2RYxiC6/J1JvA9mLefMcBb
YQwDt7IQ70lj6RMg6aw/IXpOQGcWO7FmQuovEKpkkVR58OtPR69RAig1a6bLe6Tg
6gV6meEgsmvdb1ySJwvY1tMMoGTqUjbAYzCOLivW1iTSCup9OSoaEd2p1G4u1DPu
kleJkXfLx3dXHEZgVqu2pUuL2WbCHdgLHnLXWNaTsPyLJvOtynb83bIRENYmZPRq
QFqf39gS0rAMMuJOYfR7RVrEomKKJKfW+5+U7vmxqxHs5z3yTK8rnSIQfPu8+P7T
+NIsXnPJwoL6LERcVYaKaANp3JuNkTJ+2O95i+5fZSdP9uIDuRuO11bS+cixIgI+
koT1Js1fgCrSZp+TDN6Iv1/qGHcK2zfwPnqswFZh1tb7zV9v/fAPi7TSHf8QoKq2
O87N6/u0y3x9ihxwH2u30Tt5mj7AHj7RRGMwS67/9P6DY/rflSMpMTPhPPnJVL6Z
JYodo9UKjoSqHbNKzMrMim+vEQJ2BH8lNfGO/bVX+OcVmvmiDINRn+JsZOoIh5O2
LdjeiTqq3oIb8QVseilYM640dYybbjQnS1Ff2FmhsWzbqzOWNc8ecpBZ0s+tXWyF
IeFUg0LcuSEvXIbNclOSQcnZC/0CXowsK6mREEsDJt8akh4/d5mdF6JmQ2SuebFL
Sqjxl5g3hS62JiEoYQPRehMm8VEIn1ZdvduHgiiiDY/JvXBfVRPBroqsOT1lRllM
ERv62WM7zlgebe3l+NR/UsArFE+xKfUL35JVZ6Zgq98aIe9uEd7XWdoudUwTcXAm
gNepfGhS9qtlbKhOyRejiuk681ddG9tRnkfELhuVoRkmWDoGEd/uOF3x5zUmqSZl
HEE9TMZGN08rwWQx1JHV24hJUPr/ZuCxMX+Jk9o8a+0K4+2523G63H6/PgtqjWuO
nq5Dm5SqOhfaT1yR1Kean41XZ6pwu1ZwqlQSRcR/sRRD1GSfpnBACC/duZOnBIE+
1QxpT8XjUOSmiiAFU5La/eSatFDAD0r1QUp2RszQH4asM/dQoBwmXqjwWG7m5XpS
FTqZYSRmKuuF8Lf/4qIPAsVEMPJzke/cBfslG3xKmJSb/I/rq2SMj/sNq1NeVead
B9BmPomtZBEM3/JatO6Jaoh1gOB52jEGJ3HodbspVPdpNj4pn4PvlbX2z7dKKkl5
VwDsnZwBtQ4e8h/oKBv7YAwC5tsr8Or8OzZ4sAV0k3IFEt0pOwFFooNVEfZGivC/
itB3ZOVDgniX61Luiwl+GxveA5iy3DKOEZDY9FNZAmTt5qwmh96XzbMnqhiaxrfF
LyoOTC//r48Ql3rH2vercVFiHWAOBDyPhxCPcgBYoIvYWB8msO8aI0ks9Aw1f4bJ
8FyS/XNZB3Laj2q69ItUqglLzMqxFM3VWYvfVtcU/aaAZ5Y5i5ngjDANKT6hEJx1
xjvqyIuBy4cDfNBIvHHqO/xumhCr5y3iKo2WrPoEwwxs8ZH/sZ/y/lx1ELAPgiCt
uOfmSaPvOPC1jvUQ1BX65/uwUWdcv/xhkU20V+EIMQZe5+ZFtscDkUMq5B2IA1Kl
29GBDs6w5HeV4Zj6Fnwfkov5dy5eyhwWLNsXF0a//sjtasJ+BIxst3MpNq5FxBer
3TmEYhQZqhCqxqJpt88XIuIBGmuzNjO5EsWyyW+/xcscusmTIXyWUXzGoimDkpG/
Zeyp/NOvY73aodCnU5BT1fTo2ZsZzT4tCMzUp3I9DCSP0xPYgZMyskzZz80OkNmd
qQypggfdTzxwDIdOB32htVKSKmJX6Egnt/Gia7sqGxz6URSpMq5c4gex0/t05dDq
0aFdYqtVJ7qopuveE2RHZUtBPdU6OO1/zZO0fhWDgB7oSClJ202Iv5EXfrNBzoXq
bh3NKNEselqKJ3AW2aEgMXjDJ734lvoj0u5tsa77D/R3axu0qO30xxLeEK+bValO
zP2Vj+JQGszJvK6YYPaVWd0GKCxsmTbwPMd4kHp0EvguiB8P/xUx0U3SSjGtAXkf
FYRZ5OZMxxmJlX9I/HvA/f9CPE0aPsDWYJHqDM3hvkWcc5C3h8fibQVY4+X/Ku9l
2VcMrCXRUR1tmBCStoMKgLIs5aGqq/ra6enb+UXpjcyZ42qvEO1FkptrudcBauuX
wXk0ig5IxbcZ3NRnIBygM8CvAsmNE/9/ubQjvodu+tgmBpi/cQVFJSOLMhdmIRpF
GL0/9/CSyF11gpbNBoEHiOq47pmAuTX9j4haXJ1+Kk8zrdtfCiJVjeCc9xdJFGMy
9K/WursVHfyWmTCbVc7UlRzaq45K5XsXBiHOoeHMcqe/DxRHIs+Dr7lt/1L18jSN
nvEVXGDzCwRktnIq4IOnQi/gwbVmy5R2pM/ndU664y2Bc7g5JSataKxHTpXlExa7
ilJC5trpqV7YKwEZbc985Gle0ficlAu6QhxYe9oIQKHKlGbirfvk6+ovhmmqgFgo
hZxh2vFPYGbcGLXL+wHPuQrJ8BDyJhyxG6m1FQQb/mGaEbb70Yi44E+Z19aE8IAd
JfVP5GGFlk0yOUOIb535rn9fRo+IU13lfsqI+Js4szYJBcBiWa3DaCNRXMH2oHPS
+7tUseN+z07xzXb+4oSSh/29XxQh5M1BPWgH1Gj5khfAVflXq2A7ODruzLP6AcnG
wplwtODyU+nhPoaihHD9SYwWMfQ5k5JAX6iARBIADbedcxs2CJCFAIumUW2RwiiU
U/NXK/c1BqDwxv14g1KzW78w4xA8d3Ntz0/aoe+WYucJxjpl7RBY7Lz/CdF2euM6
FAcytTSZrItmuNBhjVG72ngg8hLeyMtl4UCtTEHDPLTcqTFk/eg2FQeF8IUnCQ0b
i4l7XXe/u+kkoJL+NW37t5UkOxnZJ64MB+e2GseN95G6P72Ai1fYPthOuGZhKvfI
ajp3X7HsS6VRklRASutgGYJFf3kFP8h1U1/x/P88npFCzmDOicDx899RJtPA/S2V
sq+qfvAcqJlojTdmTeyrdhFENdgVo4p7+rdhZgBnHIlq5+7kARIkRnY8YgiV7qky
+wSfduP6DY8r8lq/caNKHuRy1i0SUM7z89HENRFWapDFdAqFEldSxQdVT0pAHGzt
8RPoau7E4+wp94nkC16B8A68wBp1VrjFUi/D1ruhxUn0Cx9x9BaflbliwP1zuvh2
62PEffvRME6yHfyck0CwYhZ+qROc6+Hac3rJ40YZ1Z4gh7vELVtsNTUqWa4euFZh
XiURlohGxHc2LQEw0qtIthAsFXZrI5h2qpiUu1cqHBNZEB2QMqiKTrJzROAwrJvz
balQLyp1lW4JzUDJJVBjLubH3pY+/2WZtZAoOTirQl9n2hOLH3MkYFQuQ4gWWuiW
fSTRyxywwwGFvZyZ2gr0bPLo/NzzEBGkVC8Wfp8QZDiph41yb9IfTVKRqyNxhp8/
g+Ow0Iw9xcMnTsEIg3rXNbhXTqwM3ogDULActge76nzgMEq1FQ6ublxoRQpD7fz3
YywFbIg/qDYJRSPY36Dh2tsi4wyQ7k3MnlEQLbhktnBgxAz7KE7NB5jAsA1RmZax
XCObRWEdTE6AfaxfDork8/EidRdqxKx4/L8f3akfgB6jnH2GUqf3PmfW5K9tMohz
drNNMvS7hXNYKB38Vl8rM9nfkSXuDEPDnxYtO+V+2iKKJokSVHDqKbrpX/L4yHAA
Cs6PgN2fYJXhTaZr1bGrTLxF73q0IjWOHWtNc1IzIccg7fkwLnnmQXGLG83UdGup
xsAHyXoudT4Khu7aSreezkTe8pBq7oXRZG3nsf/vxmj1LlLylN20K+DCVi4mO2fK
UauRhUytpeFju8Ix1GoV5tZ/8bpTdEPd7jZGAAyxNPyTFuuQ1YgEZt7snJHcmSY2
2vOFF6mHhJA0fEoEHRenSNFvkyxM0YHQGDByqQApCSdRtr2XfynHRUxA0kTPWCAu
2uVK8h5uMoTii9iBoNqa5AhA+2RAZCYYOu7e2pz+gJV7B+6iuehCSlsKTDaFWUsN
V07K+cxWpUKZ/KvHgTp5LauWX/Cpb8hBIWwnzVERzf634Fo4dgvesV7nkmIuaXD7
vLZQPVMIYiDXFPjTRPW5Q4HdKNZLbrq6t/WvzE9IXWbP7+hBxlWy0kiYX296xbso
QngJSZeX263AwQnsL/bAtBLkXQUhP0HLzmnJxzmhRnO4tWnFOgT68HsOUOvWhDsd
5C/cX9ZnQKK1givxLERt0f+DLaFcHoC6wtJaehRQUS38gVszjeBLg2PUcz5mxp/H
2z0wMzlg4npuZRK3ih44Dh/exq3EsqaqHnPiVRN8gv/BcB4ZprEsT95n/bIpCpvx
gMr8oDSNFWQDJk1Btvrg44UiolFLxewj7XNc64LXIScQR8bEUmzoA3IpSTi1vm0r
BjUQpo+koA0fWguv2VAi3GuS0Dv3XjbpRbSZ87GNyjgyHM4sU2Jv5FDOjfDhlkWF
aFffF1qd9o2qP73qmR448MCNhyLjxGwJZYP1NAZweVtMDMee7W3Mps8XJ7sVUJNY
UdXZpSB2tapQ2wjizS1LD/YoH+4I1bY2aIFYCLNAKMrr7uStM3Mf1xPE5TiHgUYc
Z6ZGcdUyn330uSAnwZN9cnvgdY0t2jXUknqlZpXsHxrMp0xy0n+Q/Tf3eNWwNR5a
2E6V13h5dTuypaG3lgeV55JaKok3anXKxycnbRDKFI2aTDdGe3updtSPY+qEtWh0
Yw/oKhV832hBSAN0oNK20Q==
`protect END_PROTECTED
