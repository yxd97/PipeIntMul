`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k1IkXlodLHDNfL1WOXkoZeIX9attBNOVcV3OJVJYj6uUIY/n53ID/7HKf4XPtS0w
0ywXIJG+D38Tt/SXgd3mpaCxw/FsO3jHJ7q6zIgpyGgRwMRMcdgKdkPudirT83UW
1piWmCcs/GBNkJxTeByGq/+OEZpdgmbMkToCX3wxTnF5tppeR5Fop+843PCUt0P4
vQfYASXBzk6DxjCe2l9LT4F1woLTCqZvC8cUdZCtlXc1nmTvj5JqYaVv6BOJeD/S
mS9B2NWRAMw8P1yKAD26ZzUpgQkl6Wp/kq+KT17OY31lloYaM4N2vdnR8u4CiMVa
NrnKBS+ZumU/aU1puBsooKC8kKqgrcxRHzrhAGx9yI8i+Q+lf5jz3OpIywH33u0z
B21TuTKS887E6WMA6kwLu1ouDxMvLq3tXNViOVIeLbtkr/pmoQmzdlADIHCIRIwm
Tj2/JpD9BXqjwJIVYtWP7r/IJKPDBdkCu9nHCd1yzLWjiDqQX+ZW/9OHLxm4ARwO
PHWL5kTi90I35GhaMXOGFca1w0PxY2EAZVZoVyGa3iRX9KH/RLb8MUd/3OBd7aoF
U+9ndCZLxfkVJMxlC9E7/96k3uKzlbrzjwtZ+/+S7+nvnFTh/5jZywW2a0N/YVhq
YKpVFteksQwjlEvuovba9npKJq1LQ49oGFZOgDfYFcL4n+9bMTbDVjqmnSdRs1nb
gZSKxEj9KeJ5JbsvupUQVhvvhp1BKAgdAxYrA5d0SFLnE6NtTaWLpVy/mlmFhC4L
6MtXf0UyiHKrFg/Zwi+4zptBLy8oZZ1bzfuSdR/hz6eCOBJQ1fti6kFvOyIgqcPN
Hp/X6Cur1QG0xopshcTXZAzCcwuMnhw9xrmjL3EgMRaz7iNIrCFdQyMsB2N6AB5o
MqsntJSODP4DiCM4HZJQ08UZkZqHW/e/VHtwdUg7gB0qZasGlXwVrcqzfyqO+GlT
bNt4mWUNKkDrEzSuHU+96OKoX4zJjcvq5KASkKYmZDitoZSU6lVbS+V7820eP59e
`protect END_PROTECTED
