`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/M9AU6NLUCHE77yuGr6wA/F4Gf82CHbtEupqe9DwusQNpuOr6ns4ULtYxbWqyYHe
8+DkHBoeW8DGFiaoy7xcZm0WGGBCiI7LkuwbgVKO1X9mDHSpKqGDScIK2NUE6xVw
6x4rooKhnPa9BUmtOUzP6QpUuY0x0bQnbC6pgIih0CrU02BvHJOnb0WqTuvg3NMu
x8zkZMK6wZho0znESs3R46MGHAXwtPN5FoKqXeuYi8zlKYiu87n2HlG31WZjU1zE
+FkE55F1d8Q3lmS6gBAcrrGmBcidBuu+/8XlkY8Ssu5B9Zwxz9EcRoBCkzELIaEB
hSZm04tyXfdxVwQh+sfswuQnhkgmfuaQDTChqSupDByS4QtHohbVt0Zo9oMwY1ka
CMPvUDsTh1Gn0Ixuoi1WLDrvq74P29zdBMDhgqLSzjw=
`protect END_PROTECTED
