`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X0W4DpTd+Q9Yh+9Sz9S31mSI3iDog+H+om6nvmXRtQeNpL872wmKvXMcLOomoy/9
Wqk5Ko0E97E3M1aa6Vfh7qGtZQW/s2lml1Gl6ISRv0F3fzuNoNTfJl5vbLn/orQ1
psnajI0iwozarAh/f8YyqbOoliX0BlkzmOTffQ0FDC0b9J+2L77x9y8vMdpb3LMq
tAuGL4GXcCSrb7g66R9OWj+juL83CEWsOMOlBzZkrFng/xbcPdn27HI+50vRC6V/
PqqW/ATv0nVaWowm+y7+1DzKZoFQbzI75wyEDmeNKLamb/KSAZb6Dx2/KFbghe/W
S40rncrBWMAk8D+Qgjpwjy12BRtLTaRWoAJAYoujh/Tpz17UTUZttRfPcvJdN5cN
IFXtOHNnq8/cnLelQ97nSgEnskwfil0UVrPX771vsmyg37Ie/FL5j/2TK/TgPLQo
wW8kt7QXSVgrsMrN71PByuxE/De4oDSJJGHNdXgTGtfI9RPHuf+0b+lFex2V6wuV
R11QKK2XRrC6izM2uwBjFRg0Kx8OOLlmjjYaHTIdQZXzEG/rkf3D5kcLYmpqtjus
`protect END_PROTECTED
