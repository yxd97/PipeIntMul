`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z1TqPc8PAhASKLdLlMfRsqxArvbqYZOaHDoBvls8QYx5oqbHKTRNyiGwZL9mtHpJ
he+vUUyiFb9yLl1TT5Yju7+tcL0SWPmVpjVhFKkUNMLxoZdEsylnIS6Dg+u8y4n4
CoRzhXMlHMSxlVRV03v8Mm+LqO8FdMdj0Rrl98JLKYLkNkXp17qMLCvmyLIMkjO3
pd3gd0Mja4b4EgSpr2UCmUQhesL7IUgU/4r28fvgehpZMIbsL3MWBsqM5jXnXe02
rBpT4Xedz7H0gtN+x5jptqqanePXRIYNMlDjukAJjTtsBkUp6WzHQuc0v4kAnCES
mGSx7+yzTciqmeJ+kWT49J16UTn4DTjnUhVgP5LSXXKxlwO5xKaTC+jTXpKQq1va
hTaXMYeY+509YXy6/aYya1xaYAMHvjZNokxIERBYns3EeNDoPiH4KrDcXmXsfkYf
jV6XmY0pYaA0W38l344TfpFelHGct+1yIQcYpnktZywXr4Y77pAxGpoewnL68Zl5
p7x+oV3DAREf8+Jwhk989wLCfCo4HkMPooewN6w62MTliL8AvkvuXAUJYab7U0lv
SU7sSmMY+VCGBzXq5CQkNIKVJ6dsv61QzL6pjAqAIcajrt5js9pX67JHMRWAWDEp
R5NatbyZZbzDPBiAcyjbTe5cW4eKznLVyRr4SpTOhuIcqWEol2jXvrlLwH6T/80I
kAAwzLDbx79NsnYdVL0fx5eib/AaNRs3RKu96GPrbVkrl5e0y+g27Ct7BGc3HWcw
52MreOmNCOlYcSiEFal15iu9YS2mMB6puU6YT3MKMexpBEIzoLLjtgi22EX4c+Ge
MCYt8T0i3obHE+2AtOWku0A3IiB7SAD6TktuRobf7QcCSD2voGbqhJRwU3i1FvmS
mBept9QXrmLtYMcPnzDocCOxTosp2Ya4BpjfjoDDfc9ebxClLdzlOuJOuqGbBkzg
HXeuFPm2QK6iwj6nXiP3Nuu1ZglEdKT4gcN78TVvItVuVC0yxNceycUBFZ3cLNND
oogLbgSIFYAQ/AUwy90VtLxoe2RRInNBs27H67vhLNkUf6JJp0e29sf2wFxyOx7E
1nW9rNdw9rnlDUY5NDq5vXT6hZnw83dazDPA42TfjuOctqBc6k+02wiKXvveWUCx
19HgFPiOJnJvgkcnMxP3NX7Qa5Q4Fe+uktTnkt7A4x/FukvKbShYfISg1YiwUq7O
XCPvz1JluSoRtC1Z2cjghJxhNKGB8CkJ1VOqFwv/vyEQiY9D84S9xXgVaes+zT1K
5kkPGnqd0nXkAszWyNfCXbUrWIsdhnqBhAD+2Y/ENNULgrAYezAb83VD97JxlrK+
jGr+oy6FQtWrTXvAgHQ3fcIWpujuRWAzHieHKwZep4vUbP1r5IofJCSJ0hy1ZTs2
GIecC04yEQSsyEI615O0qjUpQm+P1xGqjOL5CGiVsrzJHYK0xMGp+LfV4S7nOUHo
Z1mdSG0XDIBBHnhjPZ0frA==
`protect END_PROTECTED
