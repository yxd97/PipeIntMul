`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+3xtwIn70s6DRAHbdGguzrc2WwRmHPwV9QhOOL7qA4bCGHlhh3hXX00u4wmELowE
/mZAvJSaUdNLlF+ZA3Ns8PmUi9KSc5aPpNFjNlkTgecEuJaLwec7pQWw41JP08aP
CEb6xRrxsYM3/8va1BBHVC5OxM0+6nTQ0snu0Cl/xhncce7SxC8qPoOWVuL6zioM
zlr9IdIYMGjpXmi7fMZlBBXaNhYVPjLZYe2Q3RxduZKskIKsj0apc3UIUOfTEiFs
JsZhq3gmdIWxEyFTiREd4gwHMN9oQhoEQUgYCZjPPNeaWQwspWUuE29YlFPW1E9g
F34awHyREN3SVhEwuweA8Oags2a2l7kmN61JWbf1WjZfZ7Q8m16SHEfN3hqAFqaW
Kv/w7ZwvRd8m216geSLH2CwnBz+XZHupkUxZjXmEH59oMMMBrqGLGp86DadB/ztM
6G+CcNjXV6CSqpAWU4/m2D3U7HJHPQWQlrCJavGBuPYNoppw2jt1SYue/7TpwvQT
2T/dzwVCYbN0WgD9ey/TEQgMYcHt/Te7ZoeVE9wrrs2VZTDKIVqgtpOdTeiaJi/K
SGcYsIjyfXQLeVRRMBac+FHLrVKV4vYHIvT8v0SirKM1M0hqp/HVUijIHPc7Hdbc
rolAIQeF24osg6J59LomSsWAl+ihfHK/9ucJD0qwHp4aqZEqWHyZzKX+q6v8kTZP
MgiRhdH7hCwzfMFB/tXlmUMk7lZzku9XaYFlinkDMUQ69UcTGG5BYX/NN1gYw4hm
ei9j4kNzaTSEuupPQ7SkZQCJNZqP/ZO37xeLRU2lgPG8eyKKfeTOQHOQNYLPbVKM
/GffMj/dtcDx4mHZqEfW18fEwz7Mn1EpVUVWMgFAjowIs3yIo5q7UpMiN11OPuRz
dU8LfSZY+k7A0gC7MkBhaYU0g1BzJZEaabseAeHcS8Fyy1hwnWAG3Ebb/Bj01njS
w6NSTKwhFp903tZKanS6Z0HqlKMhZAyU+wc/sLP7ARShF/6HDbkB8JouEdpkhVeF
NYQT1zdzWx7yMl+rsk5KzvHfMpd0agpkqYgRxj5QWiiAQYH95aJAfKVbs93yTg18
gWWBOZYQLO2zv2+WTraVL5GKSBR5Z13O38x5wExw/uRGdJlKoFecQgcSc5m/5RPw
cRgVOKm8vijVq1ZApinxDlHWvePbFj27dk1n9LEsNE3TjWIVcCbVePsmasWxbYDA
p6OEBxXJ49kvNrvy0v4OBxrBFD+6A9x/2oRH+QN6GGpTASRnY9UxhXr7sjcHdBsS
kknm5V1Upr1HJ6Tsiu4zioN4hz20+Th+2hjMTwuVh1yTvGwtaXl4izCrGOx8nXdm
XG7gJG9wzEB6Wa2b+sIugx68pl4aJF27vJQ7qpyWJcuDMkpyznBuIXcxwWIJjg1C
7fGrWBPMwyjIIlXn0BgVIyelZzkidJMwLvhr82Nxr+pyrmWrSkB/zrTZRqNINlD9
01Q6N1apl6iKaDi01PoPKx0NIaKkhZS1RyI7bwFJaNpJ9fKk8zKemkjDDmQgT3ct
ZN5jkgSRtx1GUGVesH4WnFW1BNd8qvinbvEpkBai6haWfwCo3V95yIvYzgg74zKh
9s3U7pOtjwOd41qP5TRxVcfIJOyMDJeWkpA0i9Yoq0Fj3cuuPT71KoPxyoZMGpe9
ymopXewOdrxohabNqq9Gb1yBIzr7KyCMMGsmN+6nA/N4hPO9mB/J2GGKqupFLdY1
C42KWEoL9GQphxJrVWzUd44qU47vwdUfACIeBBOnFBMHhzE4BnYDX/+7c9Zs/OJz
dUR/MwwdH4lp5NSEdGiQuPl1CfJSoWpZLLJRV7WbfIDkBC93G5+lzRB7Ko/uwaMX
HXkOZ7aF+7wdJ0IJpdQvwHn7FgJMHnBtsPjPoPbQXoyWNeFg4h2u7IzJ8QLHRDws
ufNKXATPoQmeO4nX0Y+v6wAjq3XkfH4otimS+bTpYbKbYg9pR5YRy/kgmBLDn5xF
9ljhhLUuQ881Tb3Hw7TJG+KhtrmXxQl38e/B5ysebk0yv8GY2+59BMo4Tw13fUot
jpkkOLF2Cqwl2fJ49SH4ER0mU/Ha9OXOdPg2xq8uz+Pet9NGHy9ULWJar6l789Ll
UyXPhiCtfQatFZze9kmCo05FVjTxIOOM81OwL5H7WtlTLffFjZpdPx+c8+W6xNCQ
ceFCsFTvJP2b0WZtYxNzhbMcdiAd5+4gFdiNUyAZf8gzaSJ09/EbczXNZCWO/TEc
iLtuT+bSS/eLdm8N8NApKdJAUv43CHVIeF099uwiciiIPZItFDDyMuTg7rAhjZx3
jL6xEvAjDlQvDIibm1746OUMKll/UyNP9OVRH9thidkQ1wl4tc/OPbDkOFb0kge+
RavL00j/YyHO66/rNYZZBj/Z3p0XcP3MBO1Cog+kRyScQZP3SDNYXJnH60FMI1BS
`protect END_PROTECTED
