`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUBKOTH74OT5hteh2NTW/d0rZJAnAITGgGwbRbrjbmGTXHjjp+J2H5+vAwaVRtLE
bqhEdEYkrM0jJJt+1Vm243HZqSZgXXLBCwntTx6LYUBWQRY7ZEXkRh+Wb6flZU7y
nrqS21NrBYNAG8gBdcSS/d2D2FVcJZDXxvCXTrP0IKGE/KCjrJ6+uJdCKICIqNXM
PKfCueFut32iLwqb3YV8cUchAWjy3x1of5C4nthEgESpM2pMLnQEurU3IFwt85g3
bYFv9BmQzvfPe8yWadXMCOEZ2VRO4wKepW9SASiEr8RfdCC3c7mmiJq09h1d5B0I
hx0g8bLAzmWe17+ZYx3Y34pDs4FY8XLEPrKDkA3a4NzhVyytFrKK1joOaghqbGwc
SukDa2b57hcErmcjs6hE4+QQz66k6zQz683V3wburfd6coK58CGspiPUlpvpYrGs
kfLIqqJBPDqL2GO05zjQdtSAc2tC4p8Gr2XSz2DDdCYYasbwvjmvuJn9AtmXmyoi
yP0lgI2wN3zn7wG2XRDe1B0lHp8h16LVYEv+qoCABPAbF2tO2RBjJq2rEkXH1JPB
lYAUyKHhnwmoKuIhwQcRztNV1D+UeeDiyOR0e1Z3LjgS9F8aaRIuAMpcZnZLlYpe
Tw34ZTNWeJMo9B0pGFJgcd2nZs/tz7k/g3V29orKNjiJltIp6DTwdGkpB4zeW+wk
uI4FDg/mOIKx+R30YiB8Hty8XAq4tQQ5oajMWOcXjFrTpNY8ux1AEloWVhQ6+sEk
jArvChGW96uCzwSTV9kxZ56nP8UiY/9vzuOvRlTr/tsUlnGYC1JbQ9zy3kfq1hZ0
gn2iTkwlhPd33lCqCVIn2b422tBljSpEz6NOvbPmf37Qozu2O4//QpJ8BLIaJuiW
ug36enjK45Wr94ETD+xWomWfvAH5RjW1wJrBrOQGgVRQFXuUoa86XCblHmijG2Si
F7wcEjZ/6PbkI4vwWb4SAiVlkKyfuPYxde1GKESBGZOaZ/0iD3TBZpynTS73+AcJ
`protect END_PROTECTED
