`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P8QkAkYoR2OQbDyLQ6WwBoH7sc++eBFE5P0wp1gP9G9w1d0jwtwt1jQan6/d/7he
oGtdRebW8qaS95AidqFo9FQfuUizoe6DzaLSTx26tPbpC+lwniwcjRgSicMQXv/O
O3W13Nr8agN64oklvvs6GYByfHDd/u9TKiIBI8qBC7GY1A3ZgnZPuEdsrO+OwkZX
yVC6DrUo+s+jW8GqIBPEPryuSyjhl1K1bh6gVyle8jbUJ/Wkn0skJIWSBoJWanCQ
Y7ut2/+jFnS3CerECDoB4IzMvhPu1zsiX8XN5YEzphejgGfTn4/Nfa1LcxQIaV/8
51Pqt1EI8JUsmt7t3kILlDTzHYJk99IklXi1dmPSkVBb09rFI24z7tkpcs3wfjiD
DX34/dn+yzWKp7dPGiPngivoxJKPEB7GqwL2Nkxyx4MI3SSgw5JAibWO/NG8FVNR
mW7uv60HvQR7KHNkeUrpFzFrTfAGUqourVf6qBcFLSY7lD9JqLOaNVmP6UNrQkag
yVvr66qNloM2cFjVUtlBBkQymNWuQRKAmY6Xzz5OVUSjY1YLlLbZl74N+NNZVIHk
MU5iqEGXiZn8rT57zSpqvLTUET2cU7NjxIm56wd1Jp8RkAsszqK6BcLAUJPKdhk+
5RFsNLzZ6YKcV4SkU8WmdMst2O66ALXLINRySI5uEfbGH962jJ/XU0ILTqMH4pH3
zQFdnQpnwOdTKL2LO/oxLJXbSmGSLbH0uximUJ+PBr75zZpk1rQ4mznIr45fJFhm
r5DKaWjVedwFKTq3L6aqLYwV5dM/aYwB4LthipDIaW1Om36/laLfdRVTES4LzVJ9
U1RzXvw6rGS5vAPVPpEzPX+QTh2MFlxplJkYxo5yy5W8QiK60LTCRLqWzG1XVILH
oau3IZH9ybM7vkb9Wu76yNAztSpvZ0fvBRK7EdqESUtq3k6oOWkR5eh3+PdoKJmr
0zQYC30qctLM3gd0CXPu/37aFImoGi85cqf6ZmVld2JjxY9L7iSleP4MaIVapbFZ
`protect END_PROTECTED
