`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9X8UqQYYAZASe9M6zU47HCydunskPOnV+HlbS7iG2ygyVWusD9lfIp22msW78tvA
8BDXybb+FffM92/dIkZe2Pa3QyZj0xBTyqrKF3/X8wwWDX+zZlOZQ4E+iuQvETEI
hiOQFQRM+UuerGH79Zzrv08bvuwjWZ/ejv/bTSWmWYsfNTFleUHEX54X0qb99UuA
xBa79pRhTFhStO5NfGyxEcJ6wRbbpy947UgeifetFjtmA8ULX4a/vQM1z9JZHK2b
Jw6vXkswvwNr05V63eE3R1fY876ZgqymVi2sbLXDRQ3mSYtQBVoDl5JkMSs9Pq/X
mbP4yrlDR4UZRgecXxOdDDBYwVr0cZrEU4dX5QoNlHu8C1WTQXDwOS5xLmP2siae
a9JGTOcDIJ7hdYz7Jxje3qYej2mxXyunJ4oN9sjH3M/mJeqQHcBdKdiuYDGNQUE1
3arkPNGdrX3+P9nac/QRKXA06SlW74W0GawsU+Oxwf+35t4WkMKL2bqG5qPW5e5M
IMbuOQgEF8lIxmjjwmhyC2npspmTVFMc/jt74LOsW5g=
`protect END_PROTECTED
