`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gujypiYxc23cr7qBuHAGJU4pvC4J7ZfZ1QUXcAMK+WUKeT/YtkYVYrvXdztRet2x
8e3da0HT+cOWscRWcppKqCb1t3kQgqjmbXuYxHEXu1gzpwNC7IZ+0N1g23LJ5C5m
NSFCiddxGyy+r6VoaLjNTGpv3TitCZ1Zb473Rk65hLJ5qsnRymGFTyh5fwL/ScZ1
a4MklbkxsYZbIqX8AgMtzo3PrSteW1AmFbbU7snd1b4bszYFWVZW4Y4tAuSGB469
RvQAew5qKeZ/hGTg3oyJybqwaVzKwX8evJA5IIBeDdZk3AFrmFSI1fwSE8Fn6pX2
`protect END_PROTECTED
