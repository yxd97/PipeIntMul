`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vjbgfv2/VUFUCa33nuSeWarp7WdXl/FvmvRadDfi4IEbf6KdtnnvLbfs0VFALrGU
rymDKUrU50435CQymqwmftbw5f8huhoHkTbRllyKt2BdwtNkX+rPsEcsJzR5PG8S
3wFZ1l3hE4G8N9yY0/QA9hXCKTA6RwVdhA37AcPYq8pq4aDgBM8ZxUgm3cbZ6PI4
jYdtUfLtMJCtm8khFndKAW/aG9u6mTrgxwtTC29Wb0woiIf9grmtpKQ7R0PWbg+z
rqdoZdejpe3VrSjdcjK+JWzU+sZ6ehEhe7NoU7h23Q/WJKd8NAqZjXKJhN7ahLTv
FtuBAwJOUh6JFEOXbYCO6wSVv8QMFmSVp+6AaCpHox7hB5HJPHdfboOOHLsIW4mL
KBFaSrtpQJOqWP4iE5/CHyuUxtr/AQCWB6b7Cy0CnZcgoHJ+fz9xAYTFln1VEXkm
0DwH/gbVHrW4X+7hK4KcjMRwtambqxmUMOVWzoKZob7pwL2cRGLJjWkCCOenTSh/
dwn3SgmPLXNGDeTjuymR1obbnguA0AdNyWjw3w9oRFjUbW0dvgK7g5KVn2SjzLvT
KnWe3ZEEBrw/AXkGUVfSxvYNXGH+kB+LIQmIsUJj1CEPz3VL7dlGgwXfTqHSdYdl
hUvGHXmU3yEnPpxUkFqSn7SkcHfxD7cdWL30u2M2jhrBnuI3q+gif5zRmzuvZXIC
226CA6vdNB4fT+15ZicswaOTRlYuFuigu+z1DJxWBnadGRLmYaMr3PqLbeIID3W2
Ph5jA5ggt+NMdrmq9iafLUyatttdYcHUW2ZPN75gQDAoKUPklc1c33N/8yMAj2X8
eGFJSaF+FqytJx6P7aV7jIWG5NA9dsjpLOYDnRGY0D7xkBmkz4WCMGok+TDR0Ym1
Fx6z8Hkl4+4rq5MsOUXFs577qgWnRqsFKq8x3EIzdi64nOqdVwyj5OkAnSG0Q6DD
H9qypQagHOOjB3XcrdYQ68GYJT0DiAmsjdYKH06MB+67pvIJ2UizsePm0I7d1uul
iFxsi7JaENeG+mmInLVWB483zyjofRrys0CCsa3CqgKiBacJdbfeGveRfN/GW6un
fB8GllgJw9yby70Po+YG1egrY+d9mPIiSxfdyadEqRFeR73wRHYhXnMaxrCozxZH
ykHbwFfcISrUsgxcZtf8nUI1Lwg5t51wP9bhSG5xDJCQmm0dJBXtvi2Hm9Yje99i
M+FFa11rt3IihdE7+XHiu2wkHy2A8300xY09PkC7+POnv9UGcIiA/lxnWFpcPxiN
eK1FRJoruQD3rJM/zNCCVqBXrVm8+X4btli2S8ntJZu+NWJn777DaArYuctGrDLi
WI+z835j39HRarNrh1WEKqRLB1LGqDYB8UQSxkk8OczBx0qe3yWrc3hnjCgOxE6E
u6T0Rot2GW6EPobDLfMhZtNtz1gtepwhwJ01lY6Ba40XTcFBAc+q8EjOMyiym/N0
fU5Hz+CN1/rMadTQzrQmOuBagEelbdv6rr2FKxcqpEX+3aNbqR2fWeT3HRAZmSO7
7nwVLltMODYvbMUSQxU2XWienTcM+muoubeFrRzCjQOE1EciuZ+OGtRoIV3tIivj
hAPJuzI1cwYO+IiFmR38FfiR/NbyCG/WzKWl9BFMK7gS/FKlc6P+SgtM2/goreUp
I5gUDe6AifP/qO/vOqkHJwe0cVtvZNhBYWIhIq44bU+13dJMQD2jVsjnrF269j+y
khUmF+smpNNzY4P5ruPkRZGL6k2Sr20yow2sED8qXh9zTk9Ih+lwpEBjxn0t3B/y
3XV9zSz/jopRv82zrru3TA0Sf75hHsWRgrx/wbk1nbr7cvztIq4GVhPK/WVaOXh/
Jrsa8tIdLumVItzPnDiOPA/Hi6eiPgsBQ9A6FeoATjk2oPSVrirXY35c14ZMFh4K
pbOIfZwqdE/rUTrA3ovpvscGnvdjh7uUZr70g9hHSFtdGx9zhDktwgvU3H8AGYU8
Ccp9ynqHpAa7o1XFdxQlSCizQh2cM0CsAFaw3vxY0HBT5+k/40LCneE2f8vdNf/d
27mlgWEgdnAYgGS8KCStI9J0PcIMPdiWWDeA3ABG2+s/u2bg8QB2ahvwZ04wQre+
iNfSLfkfBvk0rKouesV76sV24507BDr880zKwv8zPSTevT1t8yb1ZdoYJGBmy2Yr
8+x9ebVBc1WfxSnvsVxd/6bUGuETjmqJQUHKxk0x6dXKCRrffgBW6nxl9QyM9Ehb
VQmU8aa63NpFQnQMeTz4d6unqY+We1bKS7ox2xsXsIh2BkNzlNiQ0gQYr9X1Vhug
N4pddVik+6HwtIonL4nodbSLlOSS17VhDNwFWe5e2F47fdIegbDr8pXgZ4ouf88W
0qxWlshzL8SSUJT34tQ2ETlEx2lNzA1GVE5J5tsoGxkD+MuufeC9BrVZxlz/XGzJ
ifoOjipK4CyzhUSOeG29ZqOVciRHtJ/gU57QT+KfnGmSkmZRm+CerrIJGVwv2frI
x0s+FWH8Q8mpZx386u5ZBIgU1QcF+awREyVH05vPiw0tTZcCzZfHwKY2GINCwS4q
GPKlIgHU8U9QepRiIymyGEpjsUNwdoJjXnrX6+Yv9846YkL82gV4NHI5R0dP/OY4
fP6PFaBf9XtEhWDI93EHNsjPB2qFqk1CTYZWuj6du7SNmYEcpLpEfuOJqmHn/4mi
YX/p1doPjI5Tu1gLOINZc/nachiKU2ogI5fcJjA5cNm207i4xW4y3nmh2XWUlAwJ
MOQPv0IE11ojV6/ASKF10aP6KQp52MneAYKckJlNe7bg5URjvQHKVkcV/ze3x5TW
GrzgVNAjTTqKVkZmqXnbKFfaHqkm8JsPVwpGU3yB7KISqBILZ3pieY2GpyfcTvMY
qaNKno54dDgIXO4TY4aEIhawBxapHpnNH5eUK3WHyXyT1+n36OUMG2abInwYcwU/
4b8tQHLFA5nCox/2DFta3HZTXg/1DnRrYKt8Vq5guOszIIrf2uQh5jjF4utdR0qZ
+zWnn8YvLRawVHIZZuVq3gv/kn0l04BzxZQQP8aY2zkQYKPKiQPV04aCygPRKt6P
aj4qSTt5PuDDsVVPm4P5rqhe7fgP7ajO6J+QjocDWTk2yDMJqjsXsvuVhZnRTbZe
Hc/Wty67GtogGeckrie2ulSsBGP5gp7nHgjhLH54OAvQopxJLlRhjhVwSD+AVdaR
SIY+/JM6zudwBoSuRJkvNUoyNy71puAX3JfcjhYpR2p0jAKNcDN+QOQ0UYa2Ha7B
sPX2at9Vb3VJnVnddwwA5IF6EYZ3caDpPy5tDQn+xyCbZcKDSotEEDEF6FW1HyC1
JBKILpuJ+XqEXNSSjbrf1sH74qH3IZJ1ZBuXDvAjSF2jXelej2XgntwBFaghMdQC
2Y2CEQE8lBQNlsQL+HAnRmnJZrxE7qVRAplsHbyCGOtUagWlfgr4Y2rWn72F+16C
n321KkdyKdnph4LZHjuf/Es8DFYrTnJQSDzNH0m4UrN04bwiCUQCR3X8WkryGV2F
cGi55st8xtkTVeqsQLPLB+k9qsVb3uQEtJHFkJG65ArNoavBDjbRhBGw9PziYtWe
5+HkFvDWIqclh2S1kMTzYgiaUn24Q3/nUG1XhlG7Smyqa4lp/bVr88+YknmJUlgm
RRK/2AoACci+K1UQKgttLwmk219qvXcT5F4FC/25IK8/M/6+LD6hAmFJ5lESviSe
9YcS0DMj/TT5+4sLaT9AFYYxCp7l0xsTqEWCI4NClmToe62E60jimKpnkyUBicxL
MEV62EfLF42dbBLzMHvs7DtCfq7x4Hd7YWgL74R/2AdK/otJwQM1IJY91ytRaDzl
jTSbeKG+Xl0je6QeY2pjNIdanpWGkIqkyEG2hgNuienxDQBi1dKefNlwvAomjjKg
UVIegZRk1DhLGf2NTSmk539hoZ21bKcVYQKVbJApP1wE912fE5DF23xgnxagzbDL
CR66WeOMNhmTRkn//OngJ1awa999yzH2Mlqo81VGs8Soap9rEkZTHw4XcutmPtjB
ncAVJnRdgmfo63I1QHs/pQmeCqiCsKDtoRPzvDnQyan+Y/ykItSz3A5JhCbmkUR7
/SVe8RJcfCun2m8Vwr4mkXx6ibf0A59+VTUnPftJPN208ief2pMh5q+jgCZQW+Vd
NR10aGikdfya9igLR7tn9uhRBQ5E/kOQB/1QV0zj8b7refXhxwTcGgWsNuRKqUzF
GnGSYcZ20QygzOIRa8SyFPMeUnqYZXLcFSI7Pa+9GxEtA13DLDjc18o3uJ2FS1cY
PIZDgQAH2bb/8GQULs8cu34/SWEa23PZ8HlXj7BF7Jc+NrQGsWk2eHDQNuOUX86l
nL1FSBetpbcLmVXZunAK6JBztiuymATYhRqECuCzMZRu5Kz+ZRcdPDqkwJ0SsovT
G4puRww9rfBmm9VcAiVtucLnea8ENd+Yuz1XxieCwlBXGWlIbBHB5TM19XvAQPeA
xd2dPmwg2VpdFhCCw7Cf8XV3INnuFCKLlqIOPvg6E4QqGA+Q1ZFAnULCe4YSu9Qs
fIGunpxQQgF1PPCJqzNguUZ/+O8cx50GsPloe7uLA3mb8f8KlwJOB7vhDbMV08rr
yslliiMgws+0fm7UdO+ji05vgAcExwbErsiD7dG5iBI3i7GMiBL/UlzcjbSwNF7J
8tCqqgKvJWP/Rhlyq+w5S6NKNB6VvG1ka15x45g19SitaOes5sZxnZM5v/VioNg9
VVw0HPiIk0P01azePO4mRpSt6cabaNimqn/etZxPz52JiFc635+v2wVM5dCaM4FL
4tbZVp9tchRjVYG3IMUpmTZu2MWdnsGwnk05VT4W5/f6okZEyPbih27bDgVJxTx8
nrDkw5wn4E/eaaM4TX+ArCcufTCDW9vygnavMojc8ksVnxjAi03gKzLdJT7OQ4Xk
JgRJ9eEK2vIo5UEwR2hFoWt5qMe6g7m0H+OszrWFtIRAdkks5cvz3pD4lxwHHmuF
ulIt5PWm7RWD6mkinEb5610Mgb3D49MNwbYW6wGDfpkA8lO6X0L12RkbfIbhGjmJ
gMvY4Zj/vkNHXpJLmGwQ7K7tIdaMSC7AY2weMH7dqbBU8zVjD8wxPge/ETr/6pBb
6N2gKVUVEdVO/HAaEQ2eTGRXUXm+itBTs7CV7/Exa+HLZubGmRykFlFrB5/e9RtQ
uM0iL3CHbAVBN8vKmaN6Wwp4l/uvcHF6TdmHEtm2mESJGmo2mIp9li6iQgd8nw9W
Y+XG+HR43yIONtN5k63XFpRiRh2Tpx+4divCbd1Nssj4X67AvexQPqzPtgoqy4db
fWTGNCDRJu0+rAmoMfewOxFedod6BWqmWrk9zA6Nrm8+z+F9InWy2yZyVrRAY8uP
8HPbEpTsNTPjDuZs6W7z9pBt1DblV3S9JCTIQDOWB6nvo4XTjM45NZ3/kS/c4GCJ
b3lmm5IzLBGsPEsPwHUAHi4Lvo7o402JEXothfIleGr8+H8/G3yQGxMWGBwPtKWv
lELoHFwmBWMKyLRLUiYt3lRo/B6seLo+vImc3zo0aLiQ7GRP6xi8M0ChMoGahYsL
4V5bD9uYaiDSYoymVxe4F5eh0PV2KUrRGHesaBuZcoMhfBw/tbeZmqlOCyJNQ/u3
hxgbKH8+/3Jt2AaarLM2XdNM5zbZseQ4Xa7NorEbz0lo65HfkJkKoqobpff0IuTU
/hTY5fQSa1eHUYgFmFu3ITkqARNhP3el3J1KFKxtXnOfyjDk6gGS2k5BUvDt+b2F
gupt+lprBBurHNUjFM2ICuGyh4pyvfYejIhD9gnupv2NxkaI03NjNkWXl+TKhLvd
2Tn0/NmCaH+5JxqpFCMDeLmwSFCEn44ijS/S0yPi4114IhSp04PGpa1bxYhoIN1m
adUctQtyUcPPxroBXtXZD/ERvUz76+lODBT4yuMmhez+QlhbxnuyNr31IhTzFcOL
tBI29UsAs5FF2+HzBe6Lu33eoyX8UROISmKmotmVR7ZO0yfAibCKXiRy4SxvCpjF
8uq3OOCK8/JuqEXYH8VMfYKu/dQI2ZJ3PeHz9EJpnU3i2mFTQM/2D45xNhCLO2vI
onCQdSOdwUWDL9kW1/N2UQW1f6wgdQ+sQsVKub2YXTRS62Mvkkvz190UzCWsQJEy
FkS/aSRJXwJ19pwBmm/HKIxP08a7Ty2JV58wl3sqp18gVLTUGxRcww/mZkbYJ9d8
t/93URRlzlrvoDQvnvYhKkB0fZ1LPNB1MufOUCj75Ze0GdKVaxWn5K/vIVe694vC
Aq0vA1HK2Cr0PnIBuzGcuBje/nU7Rw4gc3AyqlgTyfw1gWun+KN79uS2CNFPfBg4
jZtOmdPdB9eACnDcBsZJpYB8FOOa1nDKag2GWfYJg741EPd5w1+CMNy2/HciFGmt
WR8wHYrK4ealqJiA7DdWJr61Oswc38qF7s1ukrQK9gLI/zOdrwfUXEmmWfQw6CrG
2rAdXZiKwMBsu1cP0vVE0flpf846/bstmOB+Hhej381UBzv6lJYPOvttfTpMhOFf
8nBi9dr/ucteTmMgMt/XVANtBDE/N27cDUxj7dgD8X6v0iN2O2Wkhg8IUesEhSbD
pp2EPas4ADMXmsEpkwr/gV5ymSy03ADwsA1MNF0RVeESnOJkKRVli56DQEQxLV92
41lz/cZY69LVdBE+MWKBITgZu8aRj0WRubIanoGHSqwrHbpvjE8Tsbf6wZlUydDb
dIl783mVUwOa+7m7LwrYklxFeYOfaeDM4aEHIx9BdVEwp1EnoHBQ22MkKSArzAqL
bgxrqrY/W7vaS+GQveZrlknuX/b6BcDz5KaghXaeOMGVhao1ocL3PtRlvyE+heWu
j0Y0fYmzJ52CEwGCm8DIIHHfkY9yDZC92Lt1/ch+JEUYeMzzQ6jCTcT6CXwb2VWT
imT2lt3uNydbhlDYHzZcsVayChrkcrQuO4tTSdbkIdRPoTJuUVwrIPXaSCcd49ma
d7buHVcvJexFcYHD0daG1FQPiq/muLqf4XW/I2d3LRmt62UR41UA1f1ur4q8y/tH
Ojk5qqSi0YVTtePuLnjpV1n5ssOjJmp0LSejrtrZf61hQbKk7qODTssazK8aZlm1
R4Bg0no9vx7rB4gEC8KRkL4EFNSqlMfR6q8FF3i1oMI6kqtZxz4n3rz/y3DdqDnp
IeyUYGIH/wgel60AVFbkGQZAZrSFCsvfRjnjY3B51BQkx3qckICSXvmFupoWK9WN
+3vIgOhKBIVuL20kuRPnvT1mhArXrCWNqlGdrzT12wlMp3In62gHyKqtbjYC10zg
OhAHfjBE7d2W9tFXNeiBop8JY6dqM0P+80DgmQ/6B51hwsbgh7a+Ja3XGag3Chmo
L1Wz7RQ6oRVSME+llIr3PuGQGO3rw7/553K398JhQoj7PSwge5qwF9xK8X1UNgaW
XamctezJpwKsRpr2p7j1yEF4hbpest6Jo60O4Wmx7CrEp5SXvY5UeDAvebyUT7Yz
oPl6alpmrAxcVK5yaxFmhO1YqxGeWDX83/KqlmsjcPXcF2klUvFh+g2Uy+sySZ7y
DCdVJ2k6rhnbF8fdNJjgbYWDh6CDU8yrY2/OrFfytfEGx9LN+yAi6diSexJ2pnvM
t4QRqitCJtQF14P/8dBpRymtpAY9lKaYlSEZSObdphgK6XLRUaRtw7AJo08mJ42X
WKZ+xc4MezzxpJJ0MpRSzbNu0Ysch9tNWukw3pQe66JoJoKxCr0AJMmmcbYfFPPU
HTAQDsjukyidY/20V5X7sIeuNQ7z6h/+GsVsW7UNtI/FX/pC4Sj27ZJX0yval3cX
IuI7LiIbaZT6SQ0QoG1O5LF3RxCzX45LByDqsFZt0QD9E0hCI9Btuc1HXXg6zYQg
utrhLLKFsAQUwxKYLHTwNMnV0XwU+xZNucQl17EL/L3CfKBIwn96dDhmgsQHZkQS
/H5jS9BJLKli+GQEObl9ZVHr0Yl1NtxKGxCvrnv7XtHaAszNATKHUX0WXBdCzGaB
ZIcfovcR1jNHjcJHqw56rUBc7anbJUJn5SygdNV62RQ7aTJMVNcybzqUjcytrdBH
kGQLZEWhg9lUlPH7W7iAmq25/8hlbcnziY4HDEPKY74GvQvafql/qHvqVYVKqZ14
7W3mKS6LeYqSGpvofNkTf4KKXPCkvdUyHSKjdYseWcHPCA33BpareUEajTG2P3nU
8kzrZrvAvqKn1f+Np5bZXzLhUFvKm+y/gpTqLHum7mWyXbMDc0ynf/INX/xh5NR/
AKlQlytkY/esRDxzrO60lG3ap+WSoHGzIJfJvfxHaDEanVDgCf2bYjY6E3mGwCU+
r4aSM295E1kmUJQjKs5ZxmTJ6krHdDG02nXa7fJxh8eASf9lfXvnu1szNybNCExj
vSRvLuxV13gbUQDEFeWe58lK6+++s8K/l9j2MnOb6/FfZ3T5cCpbHojnM/0D9Dcx
QFTChcxGP0wFWhM1a2sXfzd3h3BqS5wiAo5lTjWOswSJyoaDiwHkK+QhXnmRpO0Y
guvV4f+3ZIBr5NKmBImZeJq2cAhcwsmWIrRDp/PuW98FN+k68TvIzCaeRAOxUeA+
wrgsW/++buBEb1W+1mN7pcQiW7mR2PWoI/C1+e80i8s6aqY8GymwuBzvHTRN+33O
XPN5/QZsgJFuPOpUmvTECWU1cNG6iS/wBtmCqAomJVFoGd47Kc/h/Mq3ohexFwEj
/EPQfXg15z/FaHsvNeGZs2PLb0ELJgadShjIfNYCsrOOPJbmKL46tDvvJSjtF55Z
sSsWvr+hVhAgirNusWrIg3q+xY9HI+eet5UYhZDiJJxDxAFJlFeB7RD3KETA1Bam
4GMUaurQ6QuaJE9rsHO5dz7HOmzRrNYGqnbHhY9f33ulzGNa6A66WqHWFyMjMh7U
C8YemNQwh8JRVvfSMelaR8iKuyF2OlZF5pwOv5q85vsjJGeSpwdM9IbNlGcf6gVK
v1WmQMVbDbZJaP7ZDVAUl26OR0564HDzuKDhE2d+pTzunU5rCDFrx9VAFFa0yxXW
uvjHoW25o1baag7PEsQ4HMgyeTXHo0gnhlSDCsKdxjdh0RsXXL6+vre5GshlmLcm
WOXi08IQEm4nt1gGAN7u1Ktd5jg5smIU3cszaXFruQGsvUhD9K54K3imnRV6YMQw
F7KNiH8POY20+1GUeZIi4wxdwwocD5aqaPoHpF+UZh6yBOebvgEEW011OZ6+3H5w
X4W29BR7go7OqC3Ty0sKVCMOmJx4RL+PeyQVnHEx29Ff7LrkuFziuHUEhJfqyE+E
Zm77gRnxaLQq/N02pxzxJFiia2jAgLNd9+rQEnc6XpEd34AUXvC+6ax+GtVFJ27l
doBBS/xLZnhtLa5oCbKWKN35/Oaf/08jqe5nGCOk43mzgO+XQEHMkekOJLlv2Hiw
qPfZbYHpLU+a2sc0i3ZqMQWEphkzStvolw8svXifLvESQdsDTCrZiZ+gaIM+phFP
S7hA8LeO9VDa/ghstAYgPwdbVUZXhQUi850pVf6zGCIu/XFXqixOii/LrdKiipoM
hYmlC7S/aECTe+9G9qdKgXGGFJreqJUglM5OFU5XG8azG06nJNJMjBkfFi4/ldIX
TEFwXgUrJSKX9AHLAZTU6difM7KJkHFc9ayZ4/MjF1CtUZhWxE8HoluQ3PBiYpmG
Mg5GS8iBz/odjTi8X8bdW6LIQQxzlGX2DmcClWcmtRTFD2POD4kWIzAkODwXV5G6
+mFys/fgpINYwnd6YEY1tcEb5Gi4poZAlrAFG9eo/0DcCVe3sTplH4eYzo6yDCqV
+CZLqPad+dJFISbgbAMPIMid9REEnNtp4fQ8/TrssQEiJtS6TtqG/bHQC4HY0MTw
oYPwujY5MnyX5Y0zSdlzt4Z1wibNuapX1H2QOpp11akt605jzhxq45AkeiZlga2P
RPb9dh0Z0sKzSO2d4LMkBW9SJCxaQMEpohb0vM9erBUc3mauvyaL/bK9yduqXeIT
x9Apjme5dviqExFVrBY4tstUVR8LnkIwIRSrAq7e9V6FNxcTDCPAYJc28V0Jk88k
zGv3ZbcPdUvtVL10sq4YHw9ZlJXcOdxoj3ezrMW9JfeBfKI8sc7Vov4JmkuhfnSo
RfRoquidvkpJNQ7TYJXkCMUpsevdGSzbz3UtSQ0ibXRb4YQrlUyT8Z0tOO51R1SP
ZxOWN3cvRj9Gkn2KmRiXdy8nkdxBbvzEtAXP2AgeKURGEAoMuvrbgVa7qBMTLFZZ
zR3v7gSJMg5a+lXi6jxmmPP5Bip6hoW9OXeiJupzbjrj75oQJNAVDxh86D0xMTmO
v6JVoOTqynnuxP1eXhhvpERhvkmGdErUmUtM5kni0gkjwRvJ/ZLAM8G0B4NmBMVv
9TUKMpwop4BLScu/S8jnbNVuEYQmo/SbItGfQhk+oXYbvevpEm74AJAnvj02hnWJ
LPF7qcowe014VyG/jufHSWAiS3KhBpu9gNtoIg/7EugYH7xwBKTE5yO/7njLR6+W
2vsRjm6DAqGXUKrVgVgr2sIWo65V1dd/ITRrgLjRDqycC5LATzlbHIfTxcG9D8+9
7iLnPuY9IrEcMzWX4x1NjC5B40fTZOIE8h4003zSrXQrslqF6E4xmyKrbavdfGYW
P/rTR0yrFk+ZA8enfwJXsiVEbjPQ+g2LMT0xcoUVCRfyoUhlwx+A9EDmddmu9iNb
4LejxDGWBy7fgf1WFgqn+PkQ141NMMo2HkmDVw686odoFEVFhmrZcep6AhCx5PEO
j3uDkcliw/jhvbhX5gfMrStPzzxh8vFVbKvsidjBZfnOTb1RU+/wWL0ODzUNAJ9H
Z/fbTeR78yydTX+NTiaPnnvSq/yPhTBOX2E63c2gkL9EaiOuYW+Y5NIOZoZxMuxm
GFqB5hkRzz0xK1HHlQ2XYCd1k41m2ImYcnq/ED2PE3934IE9v5V4ACviF28T+DC4
iRSA1PXB2WC6ksT53ZWrizO/ZlC2AHK4lJDUD/LoDC0d7+kYZjkK/PhlqM1hcsmU
4kBnzUe+OEZJMnCyp48gcxSouhFJGRGV+TC0hGK+u2e2fXKBqCvyQLk1Y7TbHCKk
+tugjhOFCb0cw4pV1kDsx4zkk601onrIbzNsNMOD4L5NSbp9es8rpQhois+Bm2mC
J0mnuMC1zLvB7NRsqAiuMrIxdI8LOUCQG3QMzR5If78QcrbCooP432Qt2FY0ZChW
/IDJCRMWRxATIYtJC979kGKHkNJQJZfIGW9UWEzA1cyl9hBShn/ZJNHfXoMW13iG
xpQ9CegzhxY9p0TX/3nEeA6S9EXo8ra0b+/d2MMPWCdD9GD7NwS5PA+AmKDBNWNG
ry2zGvUvheuJCuQtyNYmjfQDaVM4LXgOitSGfyY9wFzEt2vzcPJGCPFUNF9FG4Wm
i5izGCm9EPlrV8UqnCrFdpHng3GN7y9rQ1kFefuidYVObHeXn/ZKCgnU5E2O2v7q
TzGw7H/TrZgFTjZ/pzkfSCd8auVPbUg366dZUy1Utg9orQ3hqNL17VcJsVFqDsXL
jm7ykkAIAkPn9fg6FMP3e7USSkSb6NPXCvHrWpIhqTSB/nj8uOZL2OUR03UpAn9L
iUAi0GYtNn9w2X46ZsLM1CqHqAW+Cv4FDgg6Wt6f+jqxVRLBIITxokUlRhwxb4yI
WfQc+qt2csBVsS5shWsa1ADIkR+fd0HYQx3Y9pkBfYb08k8ZCDi6mBWQvwyJPFK6
6HzqgWUHO5BJc1GenqXUYpxpaEjsR9SJkW0MG3smVmcn0F+wGP8hvJzH6ks4D+Iw
whXArY4pdmM8IKRnBoH+RouqTnYIt+citubMXcREYhtoVJ+NIh3oXp5ctyySLlBU
ib9eLQC3KUzCP8vXROt3e4P4nrAiHdg0sDK5zVT8eraH3lzfGxSQvzXgEbAgHrSu
8YSId/u/62djX/oXH+xsZilQgTp8dEQlrxPfL+LIKh+UbbmFo9N2CwqsM7zocemr
99TtcvajzRKEL/DDuKGbNzmn3owSIyj7Hyb/5HsQhZqdpUWmaLjZp37bXSAyU4ET
jZjYRQtsT93hq0QUevR5EGbTL/0gPwZtQBNpAkEbJVWD1pVu2QF1Zl7ZvlrAyrvy
yRNlwROK0WdH0MtWIPhJHq36HEPaaUvXi/8coESxYALHzoclk3YeaXljXISy1yQ9
OS8gRD50QsZBA9a5wo1hNkT1yQwWmynnBIxEnpVcH4P1EnHahx/OuboYp1hh2g5s
FmdvCoCg2aBZ9qO53RUmY2Tu3SPQACSKbGgJDBYVv1aO8EBqHc6WuJIzMS987wRw
JnrwbTj7JSk2z3FmJ1iWJSnSiQqKsIh0Dj+hr++ItAidaIeJOD9Xj6gIiV5BMinA
+5sFYpc1PT5rV7vufyCHIwZxn4bzo84X7rRGce/7631nXeEruHy2yceRjA+FxSqS
VkyDaLPS/N8X6FaT91vDnWOS2xtJQFTxVZZaS5wHiyTxY44Es/hbAE32bRd1zWSo
CBdiZixA5Ut/1oF04LIhiB/L88efy0WeGsGS8MBlvlfwU3NLgwxk2Gwy0EJXvb0b
v2Mvv2Dt+jVhC8PTis/+I8t7V7ZXKn4f35cY9/q4nbf6BmuHMPfWqTrZXOXjRojM
AodzeDSBPxxrh41g9vSR61qKL3OM0ZKNb2Z3S6It6d2KO2nGy1ZIEn4VpXzYaUSE
Nn40gknhyYcVCz5Vk7P1thNzF8FP0bdVoya9u3u6KsRpwEzSvF2yBKW8V+VDkjcu
Dwxu+wdxzVm+9+ETZCwq1kk9xVsUEfCkEx98GMgi7LtImUOUCj9rqcv3moV5SYHq
KYLQ5eR4cHiuEjuSGUPbJW5+UtEkpQAjS2rQ8ivU253lflqEceJx0GjCsOzb6gbJ
01iQnDBwCqYJXW2JwRB5W0piKqZP8jviPWscIKJMWCTDFE6xEo3I7148TUdHQRIP
C3MhMFjlR/IfDlgc3VDPaYbDzxRoi2w8m0Y3UAXhSAxm08Xnl0pLJqrossyiwiA1
hLeqLSnVj5/LduqWp5dzVhzDoekQsVPOSCSTR0OiaQozqY9wtAkxnl5WyTZL3bQG
GePkWYgBEPK6PlEoqD8h9C6BkE6G2cdPVr66gXM1gf6C6QcIyM7UARsB/jvdKP3h
oSx1gWgWbK5vQcJKvrfBFZcHYcXuCF3WVhSqYf6jBKcmodGEwa77DAweHywvwGDn
d6hZZaBGoCKW3bOEWGgIpVY7i6nLjcw6qDqCRKKx1r3+zkaGZg65nvlxauL4G0S5
vdzzMqaIJpKBb2CyG5ZBaqdqqI3jilmhKjoHQvdKKm5/tqI9by4ueHzLSamjSIEx
ipAlOPjcMQjheg2iUkY6GoTw0HDLuEWM8TKM9lFM+/hJfaLbgmOGMjYeYW2t7fCQ
7MtKB0Z+yc6BnUOvnUT7ANSB4W5vauew8bqga4897nWgEdPQz5GqRtRB1ZglKU7i
loDoU+DTjGyCyUioOFXbb3twoUBBOa43dtsJT5Zjh8LpRbfOrp+e5infXVHqswJw
kyUE4a7LRKqsNlox9wuALfBaseashjXe3HbVULcunBPw7ZrqhlBE8xTee6x2SEZ8
buVA+84LsY/DjZbO94khx7dC03wv5WkQY+CMupDtsMRghvXe3mVyR4vddsJHV35A
B/4ToEG8ATqQzciK1O1c4BwilrSxuHxghtxZAgjKNUzlKSzSSLgiJzmfCKroRJaD
SrD5PDsrJ/ZL3SML2liQjsI3XGIVH7XOfEmX5dPEsh9Tin5YXOT2lKhv356HkgwL
cehlOcOl/M/aRKAbZjqgInsjyVnH/dRtr+hrMtSbbHEaf2pHzhV9rJ23LvRS/aFA
XAV0dxQp16VUxi8trnySg2QfEnkic3XR6TI8D9I097FA2TBqgjmUI2gXVV7Ef0o+
T17InOMOMneIPlFF4VRcMw73cVbgFFMYkYOkR8q04B9uHE0bdjmysLlJTpv6UNmS
Wzfs/u3HnJbme9035pIbKmmfUxmVYhPJig1qiLD7MUyVg52id1OVqgwUhJo1gg7d
0H20WdRGpXJGH5z63ZgW+Cy1brnCaRVwMjkCX5aUANq3MCBuLjJZnbqHZhGDdO/p
LyaNn0Ams/o0LhhV0fEjFcEPbMxfP8mVxEW3iarsv+WqvukGYI1S0JsCG0v+ZsyR
gdEXS85Cdt/iIsxsHSTnrFTDjazHkFWodhP33LpFtAaDQVLWGL3pO3lEEDeX+I5u
i4E56/dw620AWkXn/fzdTYMViCOAWqO8WsT6h0naUuzLs1z0rwXizZ9isNJ1K6p4
7+u/Gjgi4QahYwaxMaznviOpHZsdjIKpn+i0kauKIus5rx66722eeFevjr8SMJy6
/QnWSKuIkP9RIkRAQj4ZVMNhYDYXDdxlIf3L4M/KhvEtJptoM1oHKzcpX8nnuofR
mqGOlSkj17XmvyE0MIvJmOdD3AYpQ7xqjUb23w7fHPTI92jM8pL2Rd/+Ka0FpR3r
R+Nzo3N8z2v/C18ZLjkStLbP8atawZUKCi7sD4mWtQPgAEnqwqH4I2l8xlKd3CxR
D2nLaOoWFfKQK987S7fHkR6WnD7mkHacFXOIPbzvIX735FgNjxFWDLwOAsRbzKd5
4iUreFUYqQ+u2SskNziXDpMTcgkBMiqoY0u/8sRIzZrnWTvI3LM67yay3dJTiOse
wpGMCGi4IIlcxIwC53k1eg==
`protect END_PROTECTED
