`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYAdku8XHvTxSULxfEQ7C666ZQaSalMqCQF3D/GvmqL1keD3DikNAaCj4yxme9Yu
p7Z91BBpZo4loIyQCj57a0H7+eIs2v9je9wUIT9s2XRd4514tIELwuy2BxBSg4hJ
3BpGQnX0nIQfJMXkQbOTKn+9b+txpBoSC2anMwUUmaJ51w/AxY/Cn8k57IJcOcfh
oXFI3DVVs14w1iCdDUUE1X3zo18YkYzg5PElbWcfkwb2lBckkwF2hbTMVfdXaiVF
0VMszSeeC+rgykhlEQyEg4HGIqzpQqe8dtvBij5JTJyGXuuWnvf+ng5kpCWLcs2T
y9CTZCVgTV6qgsdKNSIPRDsisaadSNx90Vf+BNzokety+5eJYDpSdQaLHiqEshqL
a3qtPuiokx09pmOCWEhv7UhsuVecGgC8kJ4IyIuhfIzW4/CFUrbPKXVFG75YeLbM
`protect END_PROTECTED
