`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jC0RrdixIWTjXbSF8f8KTcPlc/ArIZwlK6RLfVxu+oAM9lu7pM6JRdMUr53sFjiE
eQNb7MxRQFZBTzYQgkMExEzL816MJCSTsKpfvW1dbzvMfQe8Rx3K5GIpqQOhrx3l
0FV8Jx6S/aqornvI3QAGsQs1+M6PWd6OLmVGgh8+oZ3g6hEGQGWgaAu9K5JKNHzf
YHIypXgDuY7o/fiuoHld7wwh+Rwq4R4XeaSafa1acmJjo5sByZTt/UnEBwpcbZN2
CQoKl928xgRfxt41dh0v8Q==
`protect END_PROTECTED
