`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHfx4g2F4XRBRGyfYmm7/m5t/rWgp9IskNPPxun+MSDEmJzM3s2JnIxCvgpVXsB6
sbi6matyo6t8QNRuaoLzLfWLs75d8omQiwmNgZ1QCJUeNKXZDuVMBcHa/Kt6QCIQ
4tGVsrwPglBxL0WUv2PnJEKIHXd13JyZ+eS7Umtr/7t4DuwBytJjG0azYFZEWUXo
hbZV9xBybu90n6XoZcGWoprvOckGsU7wDBVKPQn3bunHbM2EOcye9LROqHutMhB4
ax2e7cFRarTjo+RCWARCUh/s3/S5BPYSxAJZZHhIhqy70PiD899y8+FyJ8J7Z4Bm
7XAawMiYcHeQUA6NkAwaFia64pCITlT8dLeqokXSmbTD+L75utLSeG3asUYGDVYH
Pj2nOjSg7jW9xh+muOPMil63IheYj4wA0Qi3XumAqod/jzaBmq95VuC4wY3iGTje
`protect END_PROTECTED
