`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixTLIkavsVlA4AjXmKTg2ZLf+md7NnwZKSIjKIONic1CiN/H5ViV7XLjsAm7YSi2
6btlVkVF584xL1XjXi+NzMaqKlCK2RRWdYfMvoj5lpXISC2vgFf5sWjDdKqQOE0A
7z44kaFrrFKs9wZO3Ye+mdxmn+JjXcUxTAPZGW+tjfsv1Tvc1SR2rlpttEtQ4m0i
mstwLKH3pIZfO5928wVFeS4mhkche1uIuww2FZ6nS/bP3viqjCG0NFWKrB7TJ9DJ
rM7WU0nzLOi3vNTclfxizz9fWkzdHskKetP8TICAsySZue7qxFwISbHhDfAzvciF
HamX4hBNUr/qyOxinPaDxghHmzfV8xeNPQzenrCgf2BGCK4XX8M4ukwnQ7r7kVny
aq3nM9wROqIp53a68QIJIMakoExKznfr2VfUENtjkYJ5jqIQT6ak2sqtPDMznrlU
ir8ZtlI77PFbSG+9BDrk++q1DrKYlKT6LY8QI1Tjn+I=
`protect END_PROTECTED
