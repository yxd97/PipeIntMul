`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hqzBZ53M7hfvQ2mj3CBxmDOuOM9U+dHqkXKxebMpk+s/cPjqTumbPxAGk7YSM9It
BfxzCbiCBMT+sDwSTqEjeuQhtYG1o5BLsP5Swx9g2Ygnzbqrho2kDZqznbZyJVG+
tWBZGvYcHC3s1abckipf2CgClESf4FS15ovNZwbtOWfqPiJnnMlUUnNvnHIfTgwx
P7BacHhSg4eInuRHGuRR+xpHznCCSpweE8REY2CTy+GGJO95yiHnQnsn7JeAkYq/
B5Hk3m91jSqufueouqCkzOiqYjQqqYAGcfw5AbTe5ydHMSisu1Q4uQHR26Pgi6yR
fIAMsVzz8J7ixthLq45JzyrUhSZUMmGvjHq+Qs3zvDlWdXtSbY4+LO/2TlVut/Co
xbnBceVt3dqGxCtDh8RjXFsB930Sl/c5RQoffc6N/3e16WMTXG/4oZXuobliXkyg
`protect END_PROTECTED
