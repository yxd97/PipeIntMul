`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UF6Hsyf3sXP1osDYvDEeELt4VL6flFk6mIsN89tWqXFAv+BU4fddj70aQ2cThW19
XyeTXkCNlo6DB7X5JpiNx0aW82lqgDiQ9ZgcndOjOFn/RE1MXIkf8JrQ2EQXrVZ3
r0puvYC4ydNb+o+SVPoCkMzmmU7ZS5BAm3wLt0f8fuWjE6DcYbj7Ha+n85mLdckh
8msGc5APv+zwk45yA8XwtwRw3ngibQAFU29IvOVvS+fx7Q9mhZQaiR0qrXssdm/J
iomZt5EBmoQ2WkDnbdESMFWZdRg3V1HHesG3JhSMPSvfCT2zTPJELkyt19qgGNZ6
69KCT5wMZOlDUItZknOeZ4cZ31DPe0VV0wrZBSN4P9RPTgzui1Vif1j2YEuIMdz8
lS0b3jvgFGsvqZjfmxM1GVzsfhI0cVkwwTl/OEVxx4zeawg8HHZmrkpwtMoCFOq9
vFBXS5eeS+7XPQ71Pv0flx18v4M82Vvzjq9Usey+c3aFt9WjZCIv2HToGmsuEuB0
ss11yY9HmBT+GzkI4zNrJ7ANzYIwToJBP5mNV2zo2dEqds/NCHTsSmHQBwZr0W1G
eYqsgL15ltyiiuZGd0xOawuvFFY9POHvJtcAI/RaFJ3dGLxb3qcgMFw+IX23fW+6
DawssEg82L86/uBdTzCy113u5o5DGnRreiMFiTRb1EcRe3rY0aephQao/PkPD6BJ
N9WuTJFEMu0yAwcBLaOOtQP81sRC8syKFwcZbjRst3ig56QXNc6K9NyBwWpgbiM7
M1HbZOA00LvjEFmyEHzkp3UsUvEIpcuUNCyNhUBEFkEdCIgfoJPJQuN5xleH7A9y
eBPDCEU2GJ7uldfALSCADCHknPaydSnCe6q7w4fk+5y43vhEqGXfDM2arqOg43Ko
AxN6houwGsNHwuwwW3ZNcjBpQIirq4LEj3vyiM5ZY2og5yHKqRXzJnLtgTUEWAzr
NKGZ7ky/n49ALQYc4YbccbHW0as32OgGAjgjOM6iuBYfo5WgRRXx3zsUGEMiuBBg
yBsdrbBfMmjC0beS1gZmVtqMOpMeUCQ/sc6lVnKSpdH/fbluxr9ju8WKDTTepqfA
PCPWs76pb/XGoq/tf3qNOHWEd1cMIAsv/jRt6Mxv4P/ECrqzUP86qGcm99dwf1a5
T5PVnFG0TqnDHI7cyN+tmNOCULRK+PwJyayrzetkz3OOYUt4VPOatvJ5XG5/4lp1
tlKcnRyqZvLIyRdmA5B0V2BbMxuQN9xLIHDhYEDA4Mtq2aQmCgxilx7KvarLp5W6
EqDSpPHt+nHP9TWQZIhngo7n+//6D8nGgR6gJv6Jaxv8KM7WtIhqnyR/yJ5pkTFU
0OaOgrtSdzzWBVzT78xAenvKt9/9iljRyyRxORICY4jlYSZjZm8H6Yavuip0eN3b
8RYIBeZuKXfxVTzmeA9pbWiB/4hiDTElzoOQzHDeST6v3zqclI94L2Kh2hXdTIeH
ShH2OYSfaM1zwV8CppCIsPfyJOGcRZrXd0+i53OHXxp9IsKRrxtECfJw+yirUtvi
QGfPNZ6JP1qsx5Y5G/uYHvkmJpMGk4WbDnO4EkIrWoaV1aslRJqmckeEq6OjhEYR
uw0U7DMzkgYZrbbQ3V/1USnTYAGp9PoMK0XZV62WR2QGaB1LBWWzPb7f2ungHRdm
tMaILuCoLzIXiZmKgOcUew==
`protect END_PROTECTED
