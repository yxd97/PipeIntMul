`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mt3Tw/aRcg+2smd5sTvFSGdf1ZhB7Q1wr7K1perKKeBriryk//VkfBAosSvCsVlh
LZE4E4qc6wTr8ZiWnqmw2owWFvGzmquNBZPN8QKAUwJ5EsIEyDg7uiJRbjHG028V
SHwPhATxiKhGirQFXaAlimHXXDbVIbfN0MXJnEyCFxSYKhAOJxQVILorGQUIQBo5
02QfeVJKHnp0iX0Y+mWfn/ZhxqYIwGVLAr69lIG6NBtactZ2WmlK8ObXGJNLExGR
LFuddqtOyv9L0F7uxXp2FFSBw3aEqgZlplrB/Y6sLuWIEmtc/h2w0D05Mf2Xjyfb
tBbGKWU7cILoO4OytSJv2lBcFmOUEmLB34og9v6bh5ZNiADEpAao2emuRBZ79M+A
4D/wTjpsGOovqlNbI1SCHBYXSvOCzCxx8Vg/l83dkDM=
`protect END_PROTECTED
