`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lO/FkpJVqRxkgf8+tQ+nirqnhW+AUVFaKjA17kj+SZFtAeVWIb7VF/sina3CYIV
AnVFrz4NzTFFCI6yjtLM3a6C7QcQrmr5gxmIp9jdRmfE47sjgTkVk4AtvlmfIyld
KJtGrSSl2P+xoIclhV7TJrmaFaE5WPV0tey6Frl+pVkAhYVtrGMnsAxs0Rmj51YB
+McJJyU98oEgQqIJx2SkPLPmr9n/UaqNUbw4Y0PPkRk7I0dGCmM8Lj8bDwbb9Lxv
6FR2nvWWL1phG0/Y7/tTkADj4bYDxFxxysEuQCK+CdbOJ+LzU2uE+JSoQA5+JP2W
Zx9r/hwELdE6G7+bZjgnuSpo1lcSwtyti9fimhqA7B8DNU2+9Htk9cpyhrc2ZzZQ
/uOugfm50Iz7vz94O2ItKw==
`protect END_PROTECTED
