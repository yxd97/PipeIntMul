`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWkm9UanKBq+mnUKxSlNG1VjwrOUbOcrZtL6EoeAubJDS2IFO1uPzboG1lmTjle9
j59yQfgNKehzIqnkgW6UGD56nh+7K+H4OIRdmZN4GyMet67A8j4INFrFxjJnkghv
OcNWQRWj/HeyL2DG1+bQOuaLkVjgiOUeykj8p+R/K/HDAl3PVR8mvUQcSG325YnM
tNzEhz4wqDTVW9UmvCvuOb/HuxO/4WYKLWzbdZJKoq6SZHNIjFAj5KAV0R2Bibe2
nP/X51h0aSyjhxt8lujJEunWkuPe0lGIxkDgiYtZL75GkwMEWnsCE6SGBuVuricY
eOg24CxRa/KGS4ABQxkTq+RYdWZO9L7UZ8fWHjUR4eqsDmjIJ8NYQOgC8AFIhb09
+xaXE9iieVeAKat2L2PfXRMS7zwY5sdo9rRiEglj+/imUkO3WUFUXXnkN6ynXjQN
vrfUHv7ZBP75tdzGlDGIax3Lom/lhRAEfKFWI+RhRhW/KhpAJbxemYSAoMtSSElB
r3Jhl3PckUj6TYJbYkxXiQ==
`protect END_PROTECTED
