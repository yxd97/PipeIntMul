`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WY3v8m94HHXiUBGzG2AZ5+dspdeBpmAZP4ZRlzQOhvE2gwAc62whEsY824IvhNNC
HyvCTeVRyuMnvU3rFELa/TYE7X0wc+0SjkCN10ek56ZI1JAf7x6QC1SWJzs6kFlE
kpZvc4Nh1V1z2ByahALEKVyc9siQcw2bXkJrVD44vqVYZhgnbLe4WpnQiqWT2wAP
WTVGEj4gahU/UD4IoSEQolJzk+VTSa/QFS2SQZlzIlJnfKrEjZSR9LX2qapawaPG
cpEKvzhPdbSdbsOJ7Ozxy6qddrSMqplLntYOhZwaWS7AQ2ws0kQIi4IYhQzn8zBF
BcOVBE6DIEPET7zEDGQIEcVtcBVH+Q16fGdT7hFsOQwFTVz+AyHvxYVshpSvYbts
1JL7HCrce1AZ7dlgPoytSshBn/304MNGYzS53npur7mSc7g4jYFcxnhTqI1P7U4j
28vYnS/Zql+PQcUMoBRQTD/rmXvkY8gzXT/pPhc/sWMNBA8bUsUuNDtfayvsqnfa
7L5oLT4577f2Sek+mlJnZ/2IPcW6aPirydW9Qv8KA4LFLPmLH+SEl0sR2TNEd9rc
IHb5sswMkNcGLAQ5B65LxsKFyzkcFzB4YCj5ztW06Ohw20Hzz03qORITlm4h5VUV
E1RuXG1/JDo+9P5Kc6aunlFJlSsunXpRdinzCRyYWvoxK3rUsyDlka3Fxqfcs098
qA8ZsJx2kf9nKfjlXy7BHHexj8mHIdvcRwxn6jaX5JCbMbB2b8i65OB5r3DgsfeS
Z++GSgGa2V4577Ajk1kKL4sOUDEMcq1D7r5t8UXN2IzqY4apSgXrQUDDr6S/CaD3
G/lb09Uj7R/Fjf9Q5ExESP+TMGUvqBNvP88dGN834PgEVq/fFn0EdLpk/eUudDW1
Xm5o2E23mz2at15bFRSqNft7gVHckDZHUmIQzcFJPtH5FFABscJbpxeOuh3Rtx9t
T+XHCBV5NeRMBHiqwZyL87dLcpdj0W2X/XVHFEdtuIwCp3XS/LXuWoKdofYMUSnn
NYFHtx+QtqeJgLR+RadtcgFUWXrr5r1GunQN35Tch5dowbXPqhH1Cej6d3WPs4a8
I1q8QhzCJxm85yvGDTRKUj6O+Mk3skFJvRY2fDzcjLUabEitWdT1gB7p73ZS8jFJ
OmnJMkKkRS+2Hq5k4ta1B3ZZM+2IlTVt97qq6CYYSknp+b9nEx3U6E1zJB5XX9C6
qltho6iOwLGckS1KOPyt5r+Hnh+3sKLo5dGq7nZafgg6JhL4d/GcAMAj496uSA5o
W/X2tEubwskn4Vu5aJ1bBMFlFeGqB19AsyKoWZ2Dujf672vj3K3+Vri4eLPNen/4
8TljepYxBFALl8fhld6nf3iuPqkRsVu1Ef7pFwAgM4BDZJYILaq9qmKo9dhMGmUQ
zYOtpaQ13kIXIF3AB2kZgHS03Gz5uTUI1EAn+/K7EeYbIZ8t6L2mkbz/b4Bgt6Dj
a16Ftx5r+qSGsj7AxVzeBiFlUi9aWU+Dt6BsiancOzFJKksJMl3Zo42RWIsYHUiV
30MYQa+h3qkff+pPsswcR0jRMBA9vvX3BkNixMCtJhaR3tJpiL5m5vC+GPE7FILb
h2/Iq7K6jcmH1kBlMHVvuIbflhprqTLytucDaDiFVaj7yHgJkzc4Jscid0RwbqxT
ociL7TrtygYzqt+M7dxRqCi7o6WsHMdsyNuuV5bC4dy7uyUUUrN0qgwJRLI9QjHz
wp/KboVk4X8Y64okQnyt3oCS1mAoRc/U5xHLpeRBHpjlZpnvI8BM5TfnMxr5prWr
wFd58f5u6g7BIJSu19CoWW3fbP3yJbBsylxRB5vWm24lSVzq6HrTqc7cgWwO9hfJ
O1sQXjJ/v0c+XbcnFxzxx8sbaFP7QClKVEsmlh11gcTSv4uqkNl/mV1M9XKxvC56
WyqiVSsiBiIgNW2S6680p3h7/1JyXIIf7pBbO4b/sT/82oNA/5NOPcK3UVmGOf7g
InrKp76lWS4Tl5bi5cNy793/qRYmvtofklcil6TDBcACQlOcgPTJEyyye/fH72sn
Y8KMUjDXAbECjo77816pJPI4U1U9+E4e2eXQnEQatnbK176rYIqzoQ6X447yRujF
NQXGweTAzaERRYttAXgYgLnaCcFaQ3x/sl8TOxrnHRB2APrcQ5Cf5IiMm+paqvmJ
DQgWhoWCnDwVsRMcqBhLsCnXYu5Uch0l8vx35s5TP0TMnRcKb4Dm1fvOwnY541JK
cXbwsPZv/4szd00hgLV6cHTj83IKgAgRVqb/sl7/zdk7xt5KYKTCSvQTmu3znm0M
uJxnlthfW17KdBTSuOeK1Uy5R4bccaDvZqG9HUCl7eaFdYWv5Er2+SNZ7QD8mvEw
cNPQ/OrWbwyFn7lNaiiykp7Z6UGVHL5N3+phZY1DzpTCVkAlI9j5rEjv2DyQtOEz
IV388UqKxj6Nl6jfW8pwQvhf/YFxhSZ2LY6RS1bHYOVswPERQ6vLHUAxKFLPIeeC
zMAjl4Qm3yjEZf5dxP2oJMNx78T/OveIPY5dQ3c6sG7vSckFoi0KJOI6eoRDiuqx
NnNXNWsr4ymmbp0yjOoRQ5lcZ8rhNMEgFS6CUhBmnOE=
`protect END_PROTECTED
