`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cn7EERU16pAezSLd5EvYUR01wgd1x1gcwhhdh/KaJ3a4VahH5sYWZ64c4OKnHN8/
F/sdYEfp68DK+J7fDc2KxwvcOAS+5s7sGO74vkyV7J9+BvWCflc5+8z9t5lBwME9
pUfo6xmgN+MFGYnHp5KbCJzFN7Z3sWNCa1uPAw4MVGuoAa8r7v6gu6RGise46dLq
GHIianp4fVauUb/rDlxEKxEClkJ8GEx5/zQfW6LBREaunEMpHC6bwJrSgweRcPL2
A+J+M5G9SqH1VpR0/LbYe5EVDHyzlonhDhl2/BQ1Z60dMVJzC+1CuQtQUQEluAEA
8BDkrQmVB/0u/X718ZiU7T1sv+DVT5yQa48iyVPiKvSClcWlfmlhrwNTXs6CUY03
`protect END_PROTECTED
