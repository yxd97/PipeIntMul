`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMK1vYGWIDGHBM97TnZsht5TOFqaf+C+o7ap0bPzj/v/CA57I6sHOrcLbmnFInui
Kn7eMgzCqhHDAxChe/st8UsjeBJMNtjtseU2Q7uJsUA4kgQXFz/w/2UEiWgDy0Kx
kiomi9Vq7wofHTGPuzGXlgt85J7AzQpHd8latO7/yPQ3XSdOujpOLZc+N6QxsKe8
Rn71xzJ+TU4Gz5KLh7TdtUOAv+7usdKEJsUqSFzuSE6nnx7zZZfk5Fw+W/zpUM2N
PoSjl1t02EaUW6HUDL9N8m5ekf2nAbgkhSR7MkHYXlc=
`protect END_PROTECTED
