`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a1qPHG0Bm9x6yt6tqYwlIQ00E1QoMF4e7Rt8TzZjYd3yKhIiMHtzi+1+veOsGiVC
QKIgFZLi0VhkEm1QGeTvu9L+sWmHOx9Vw6FsoKyCTlHD2yilxnUTc71ZNQfMyxRC
g8cy6Vf9ATUkJY4yahV7o/fDOt58d74mfOmSUcqWVOcDvVUiMF/3wgd/s4XgtXm4
qdMrRKYCR5ikp9WShF03Mu6S/I02AIdeHlRHF31mw2yOqhmT39o4zyfUD3V9OBtP
6Ll6rkd3Pol3OLmWQ10BZ74p7ueOLoZ+rMszrrB1eqeDJiRK4+YhhO4++HCCE0wK
JESiUyF2lhKM+hK5NowKY/eySaG2NAERTJXLDm+4GnXHKEXMPk9zHb2K1M6um10b
mQpL3KNPjAgnUIRQQh08s8K9xXMfmGVzm5ui9M71+gxSxRuZiFXqKutR4qJZGEHi
biZ5ZrgvFBUOZ6RC3RddPftpPUOvUhkRZH7PQg6b0+SqOs0ASJqI3iOre0R9+oPn
FYf6pQ0S/gS9LC366NThhEmo74FRG5aKpe4pt2i5xMg1Dh0AtJo5RspeJcFj6XV/
Y70cbJuxGgHa4BS6k6kCwNuu2gxknfL5v+QbYIUhNv8lOZfWZfVcsPTjEySqy37J
ZecC1h6MehUYQwVsJMkngM/gHdkwUt/wkjPhXHll8NtMBqtVc3pL9/eeAY7em8xJ
UIV3GQpeURyPqvjJf9KYhj7s3ziwD6i/4tzoMdiDJ1Usyrc37VVye0pDKsbImu6a
tr7TfNaGLZUlbquXg+U9S1+uyonLBhHe44M48zP+CPkLqbAwXPodJnsPLcECyxa4
ToGqiC0gm7RzKXP65XxEIxo9ZnGxwSFiG5r1Dyxvj920mK7mqjh+K+jgorpHNupW
bMd+8Iv2+DJYViX4Vg+z1LIproYTmerNyYPUYO87G43zUg88vdDFJa7dktsCvsH4
Tmz+UCPSID5ntbalzWft1wf3+O9fjsMZFLrTmoa5BOTRXz8VsTJAH+OyiUOexGZK
AbXKp9nBQoC84eKfea5B2paLZ7lxdfCm9w7d/jvA57mDhT98yiZocKpzS9TAnhOn
YMwo/uS9fWQyRHBOUnRCKM7w6WM4CplB9jri/btDqBKQdtlZWh5SXFnZkercdL31
faWglMnStEzfoDjG9TPAqQi4QtQ2p/9+GXXLdKb9KyJWwyDBBg8gtxaKqshm6cjR
8cRuF5mDpk4DC3HngzHs5tiJB2bNbWO2X6Grj2A/p2NYwgdmwFMZJgpRxZbWSDG1
qnUoKXXNwFq90jhv05E69k02om6CpIZvJ5RndGL7MAE=
`protect END_PROTECTED
