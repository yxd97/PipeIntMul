`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OlYt9A8jKKz7uV4fzD/6jAFHnRH6Qj4MIBLUwDFKAMopZLv6pjd0fBG8UFPWfRak
UsZX/wiT94cejN7ndGS3kMjGCBOP/8SDzzIM0HunrPGZaH2/QeNIEHZR4QHtdul6
T5xOBfTf/4ucLkzJLrUo07LI4g9IdhK2StAOTL/CVGB6LHwNE84PH2vaXHhAmOmp
BSKZ5NNMgvzFMj9MUFRH35MxD/403xSy/3TiwCFXDcA7m6ZjhsfXovU1ohHbFGvS
jVvoQnEHkon2U43RoeH/UR1qiAq9zr57sGf3ewrdu5GtRCTRtRW8rcesUmLPl2J2
DnK7bWOZRKJf283UQ8Ryit8tjoNL3/+O7HCkzeSEa7f+jNfzi7fpnZlqsrl2SDdE
RHNhGeo5aE/s3VJny2q1xBJon5/cGZWy6j3FkEg3E+INWCHwcYmCxFXdkhUyGOeE
wP9bRhut3NwK+Gd6bkDLKXtxvMJqpW2jFK5uBH42UqAzLTb3ka34a0q4wdZuIsiw
Jyvj2iaUuUoiuCs/eROZhG2IwNnprkAhUWl9EVBzI8NAWzy+cqu6WdCyteZzm3zd
+/LVO176RCc9BfQ7RYEHE0CMlo4Qwl+1OcEdw0Wi2+lpVhe8lhC23U3jYdvRZOYJ
0y7J6cGCurhJCS6UiTHclMRJGFUbEjE5tjJlvz/uOMG0Ta4Yd6r6HiBXWFOGK6WA
6IIL9YyyCH2XRoe09qpRifub/j58ZNtUpDlokek4E1lznwtEd/pLdIBOGUG4maQk
sRxSJc+Dya4StQEPQHoe/KXCo8XQN+xNkeMecUeTaXsYq2dIH4TV8ycSwNdTvIaK
Br9suQmy6UYu6jNOioVYRg0dlDNsMRtsQ2sKR5Gh2H5X4rskX8zRIPcgH+0ZYMdC
RNlMoxOxxIlbRlPi1sd0VGl/JU6RNfZy/P9+JbR79DXolLt97dKtPa66/7xNrBxa
IcdrZZEq45/l6CAU8B+9Dxp8Bkfnq2lcJWlzx55/OCo8Vn0EAsDcsF5uHXsH7SYP
M2j0BD4yVnquQrKL/pLRA+rS9NhmNZyESPc8t+UVVD0BXejmjFE6Ri9cImztncE+
NDyVA9hC0YAnGIY/DNFiSx4IImZ/P0xg9l/6ran3teSakCFjF+96/1fq3rVvT0IG
3Uw4tXG9xIhLXiuW+RxAoSoqKkO6oPErWZ8i5LqBuus8vX3sVzkk/f5LLOCIayeC
4mA7m7SkTBZhBiE4Y8h9V6U1jwln90p7Kad38NvkRikQTNhbmry/vgaac6c1Sycl
SjMcYS9ljYXaGFyCygRSo9oPZLiH9RBOyrYTz19TfpCYEWPTV/styOP1JAqjsWzZ
C2bFrNN/PTUcZ2A1157ltNm278wjhhRJ6Pl5McMB6IK0olGtPaMbq9Ov2XMUxKVN
UQ5gp8UNZQpZVVQ240VRFVs88V3sIqhREsse9D0j4Q+NGNKwxKkZYwH+kyfZFN6V
zMSzl8whM8qLdX/64Zz8TnvqC3ozVv+j0aNFh1GxH2hZM42WYK69J0NIg5N+ebRz
PfYVDcLq/16WxyXnNJCpt805UMj56YcT1S5FOWTOVN59KEfWmchcgjzLDdIHiUJm
puMsuRRZbkYvokyByxRorGAU9h9zOSsSGOK+xIxt9iCMz/OvtG4/KmQZrrEH8/4v
yuKTyRyoj7zi5V7y9NYc/s5cYkj39cxZN0acbWL/20wS5jl1IMWSC9/z8DgI4ROc
sOUsjGPwh3CUgI8CPBZCfPXNQDUqzlhtoIoqaSdYuPM1JGVaXIa8ifoMgWosyz3l
Boq4P/ndtgDbcLTBspusGNJOvjketBc11czgg1D7MA3TYq35pd/c71Ec6LKH3WMz
K7U6im09MTgZ1z3q48/12IM1eVpAQAFMz3xRA4zdJl3bX886K6oJE2L7KnA5Q0+W
IUyAl+oTl7TCdRTay0xcy7cUTAPQToQAJdadimsDJQ8lW88oUzZqjOQN6RhLhVJW
6KlgDYSqTW8ukjZ97RiwqwA5cQDqNlynZeCvNEYZ4BcJTrUmDuy0qtHojDoLnVq0
5zm/7Y9mW5gkobzrIF27EUDc0dcTTMbphAR1a3g6SlphNk6a9H4fcP06/w6aGz6H
eNTllgkznqJRBD+orIS09vMbx3mdx4gIFr30SObqD9+aWtkBNDrIIq8eOcdKgFjy
8UlZTrOad+uWMwP0WPwzDb8FNJ0xY6uEA3SDIWXE5djzvK5UoEObqi3NBMxXmB7d
Hv7z3CmLK9xMc+wabeKt4GknlLoJWXXn6Gui8Npr1EOf4IOIKWSj8LfpSVFVODgr
3MJ+ttwst1EThUWbSBhMNojmQnBTSmwoJg4cdCSZec5SWHYW7OAEQTLDK2z2q+K8
a7agSFFF+DfvNPZ9GeAjp16oeWYCpkvYnpi9CrOFTk29AkhgvWrn61/y1TPLEFwI
AHOphveCHkJOZLVzjEMxjc9BhcCLR+ILOCAU41iVkJSCtF3Fyt1E16KdbiwTDqv7
G875vZG44vUsL6ayOqrug7UKVd+aUXOvn2E3KkN64wlIwppBA2w39Lz1/HAhnHKM
HY/p4CvUc//aw2ah+9RdkbGAQ+YXKzvxmFJL8m5oHmvZuozooBCzXh0RFvGCdJOa
1CxZ7Z4RwgOmw3fHIW8NVHAC+rAaAsaCeObcJkpI0UB3V/wpQZwLYPC6bO05YZw5
L/6C921y1gbqzDBzMqArrpsylf7+xvWdiPUN9yYSctURGjmNzxB6gYqR/RJxXg9u
Idax73r/BbYYPi8u1i8sRbkDZ7o7stpD/+eyZCRPNeD+++ev8oES3R4/IemZh9Xf
DtZwACRW2Q5VIdydjzhh9g==
`protect END_PROTECTED
