`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+7qWuIwlwrGE/kbT7ezgh9V6drZfrH1poUAjqLEbnZ32QZITJJmGBxpwX/QT3PM
fGT4GZ/1tS3Q7KYkX1DirpTss16EpneAXaK/Fi9PHpITqhvGvLfrWb/Fm7ib22pI
je03T7XkUjfLjYOm5gpMdpkY9+LjMCRSNajDvk76cAvsPHLwUOz3QBU9sYAWJ71k
aEa/Yp8hLbGfsqzdh38BikCst64ApzjQCBA+Y5P0+jZgZ39PYc9/n+H2gV6vhNA5
lpNjviCi0AUUeMUBR6hxhElgnauMbnVF6hSobxenE6rTVSQBQNV2WHxv2ZPxKYqs
AsrvErBPpFeX+EdE0w3v2GOowuU32Dnev9FkddXPGIHyXQc/5paK59OxgEySIi0x
N9CuPz5JfBD1H6ngOhULafdJIL47/8fWCJ7pPbmxC7rVqxk5clWtpYOlCiduXJr9
b95USzpbpvMKuzvaloRvwBlcbtfU6J0oM9CfrBJU2Iy0ESDXIkVpVWxCelOrEA1M
X3KRuPavXJgoaR5tPVAMPNvPtR2H0GH+gToRBy0EH5yPS+2t+/gRAO/QHqcdALKj
g+GjJc3P+0ZWRLay5hIvXmxBruJrM10y2vIzBaKDsxQPOFSufn1+XfkndSZUNobm
8yp7SMvSqRYjuQ7MCT4DShutjMKj/YTNWolTtJBYG6lA0ltLK4pXVPgcDxXDJz3G
T8v8hYrIW411xcGPFUNpdGuPLLXJLm1NbGfZq+Si7IQ9cJneIU81Ad2WYsZcwwq0
2DSaPpyOIqhg1qWI9wAKNfXnUecmEPRNsDY3skdbaXagqvA/ISx5FVYeKG+LZt/C
fCjzlU/UO8YWrEjty28o30JHWrPkojVRCR9Cq6SOTPHXIVdesZA9zJqr33Al4CgZ
EQAn9jvs8XUE/vqYY9/XV+ThE3hFs+ssLj4MZX3Xx8NMn2vA8XdOTHWvykB30wg6
w8PrNF2Q265Ng0t9LijVrscddZvhxoZCEGyUGNbULGdiqjE22prIo6aZM9lxJb+0
O8aBBewuXIoaWAPdxZYZ4fXCfaRXv6wPMg4A7jAC6jIomdK3YlshNkhVLAxCTepZ
E/X9J+0TQxbghmG7BzPDCGI3CuWGeKORH5oO/eSeX+lla46f+GDse0p7KU94TAyr
9x4Qhq6q1o7WQAsMcfrq7mnuMMGI5URymBjFAonM6bBnK0QMxYI2FSORkg1W2q93
ekQrsKTD9QtsSBCE2z8y+lmynQai0XAn6eTiTOLK0mI=
`protect END_PROTECTED
