`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9j1MMNy85f68+eTLg4p8MlPa3RnAIMaHwAaofTHQoofzCmebKGQnYImZqHNxK3hC
p+vOwDOLU2YiDNZXqWdp8HSelx4lJGk9J13yV1DuHOhdEy7WbS3v9w0xb4810HTI
JdXTSSFIr8bbkYFgg9ARMEfyY1pXt3b7a172L3URKCj8uaY8yCPpiHbH89zeF+dj
FV4jW9p5dBkJCMcZ3uE6LojsiYE4KVS8Vd4ZLHSBAATWiGYhoSrEo1LabzKaxmg2
gl0QrJLCmym9ryc3hwVyQih/OaB1iLywQfafJyFBu54B8/pQvrXAnNWQlf8699Z/
IR3OpT+Gf2wr25QbcVO2VvCd9iall/c9FQOCu+2+1eC0hr/rZdcHLimP+ZWRBkJU
PZmxUZesYw9EU9mRH33N6hWkmOjlHMiJjQwbL9120/R+/j7D0IT6JE2ipSOBRmgC
fzsbHl3uw0cktKWsAdFJ+agdQ4dLtc/yC37gQPdOYkEjJtL2icbMB8HUjV8JYIvu
kC/TquKNQPjJA69qOLNltocHa7CcKGYAeDre8k/Nhv5y/eGg64CCkvgAKVpEBmiM
5FPRSnRHrlfvHNLRD2ULqX8+qylOdta/ZtDAzE9/YPR8m+k5vpBQbxPud/3H/NYv
4eGrWYb6NaOsUMJNoKcFdGz9KKJRZy8zqz1sf583ximJTt0gEmuEBqP1r/NqAyS8
kFLp9oqMjAd8kRHfiPPMnbJ6qA/x7jrYSsg/RAaBBNGA8h59fd2K0fzV2SKUlyt0
sB3FopxnvFdRZzSohVWvisbNRrKHvIx2/StRgagODaTTIUYKtjYWvS+aVUZl7ND5
Dc+H3I2XsADEN4Eq7leiAr3hY4LMXODzjCAYFzj/+Cyxku8PoYTgbN3HbQxYi1Nu
uahvCDppikMWPyEIdte0WY08BhUvKH3v5VbXhdou9WRXzkJlu7PzXxdanPbVrdJZ
gsRCj6TKvdYiu+3BKLZh5PCMjyhY2cfMZjCPjil1cg5zZ1byrWTwZ+rSZWMCGahi
fHaHvlmW6yBt8TrbsYwIBvxFxTvZNupqYB6+b1MErXPlCFoLvWpLp3zncU4uavmu
VP+HuI3ddqdvIvijhnOYA505c23U6r14Fho3O7zQ4jNenDZOIm0/ZtEQHkEsL8le
vC/J49lLRr/m7qKtjLN/yPOKnIU0D9Lumxiv0Bu9yUVeI5SujH4GPliZniz5K1LS
9HId1cigE+MT4wY3+aiwuuDloh3RE4DgXn8lsNHaDhCj8+ns9MjHrP0iOl4Pwgm8
Yh94GbeSLl6YIjwJlabzR8o1ybHtbQbsiHuqi3yyWkEUNAhQbkDLXSxsOrOcC7T1
0jkxRfURufy98VXfn0EfqBOmP4WMzLuHgqaBYQHewSRLVMG+99G15gzCGpBB8KKL
Zfk0u0U1Z/fvL82Z8KMH1rXkUlut6yZbR8Nsllup8SgUwjx6WvDLUDBh4pqICpqF
LEDdmDKR6jBvKD6OQSNDmfmwAD6Oy9bV+v/RfHQe7SkLsLu/32A1L8m7bEQMRK0z
YP0uFBLTDEcNbu/GQId4qYj3ENjGMkd+2F6IVuXywLDVwgBiR/j2ePKYR3s4m0rO
PW4qWUO9nV8eDN4mM15UcvJSMuy0AWdK7E4URVZpO8lzGbsiy8DrE4aFVmcz5ail
7xrAAqYdER66QxbYv6yJPHZrFPZ4zC0PzcngXcEgSaa2bbW8ifEQ8Y+jBGrGWIn2
5DrsNmpS4kNjtEJ/KOZ9ba7ojbs2hr5+oT25u+T16+Nde/icXprbRojte6VXh18V
B1n/2sKE1YezuFnKdiC0UkWlr3rdR7aHntfbswon663gVIQqvBWrawroV+zsqSy4
wpw0L1wkZH5SzYe0e4Fl6tWgaa+Tga2/LsUKPIi5WkLB/j3vKTnFYVyMiRYSIVdx
I0ZmToB9+3FqfilHqrL5jb4ZaDQ5eAo+0gUNg+hsG4BnuYiQyHdoZjmXCiC2+kAn
oTS3a2MXBdMRPxH6FyaKuCIz6QgXXzDiXP6FCxoC4ZjZRSSOSB0fEGS93M7+JkU3
jgv4w7bkhtxAOLIWXlT7LOAVflGfFbkEgq9wua2PJjNTuvgap9aECCoKPQ9D4B1t
3B2IZmaXH320aH7bK8tRv1SO1R2BCwA+Hg19BqKNFoqz9BCqvlYLCTktL2uDh+wn
xrhNpOKu3MjJV7y8Os40AzKjzAm+cFMwgd1CADiT1trNzds/nQ8ofi6HSUeNVyAH
vp3UjmSUPQRZIf+nEooylR9XXFOyxSbC3KpSNqaHitfeCr07G1uh7D2ZmS9vmwQj
5UBHF37yxhjuXE2WK+MXwlQn6qjeJ+wI7qscUoI/0mf5iinqmZsgXNrL18dStbDJ
C5PbYGVRy3JGxr36meDb8SF4Pc/azh3GKRbgvXCnXuAFQ7gMnDxbVqTtqMpVV0df
gUMztfb3aYTJxH3goRCbRbmifL55A0RMRfz18xb8DDIZAvq2TBTcQHJ0p7VyGTXR
zDX8Gxj1Go+XfVkH7BPLbCFBoDplT7g3ovHGXMB56IBxLEQ3kDsJmpB/F6OX0cxY
5Gv0fhIp7zM/SDFUZwMQX4TkfxEL+t/rZr0aqfHrydTDcQ62f2ruyj5wNQ9CaDkg
XQxwOxwSIKF6C0oJZ10jM9APoOW9CJmoKiWBHkapPhxJwLtwLQaubXFF16HYYwfB
lN0+2aSNK7NOocohzUgUQJeX/2Y1yGJ0g3c8ycohoEcLGmhObwPgEkhokezNnKVo
dYL6LcAlrnle+BtkV8968mtFEqMMVWtzFvd1znIOhM6Jdi+tTpJtU1kec7jdK5If
/ApyUUiTgKm+tVUqix+1RbfM2FXq+kFEN5VwaBrFShTnWwXWuxD3yRoHRUEJJEII
hsRXFEW+w65/oWemL9hzuwPN9abJqFwAiEMQSJ4B84hUWtPnthHfWNxK5eOin43J
CV6sKAstVKFY2c5b6yPS+c0Lw2I5CK8C9cMy71a7bzln/goO6xYBjUcDubKPRgiU
RIgunfNGZBRablyTk9qbEA72qpnS2ht8hl/iemDHLfdGgcILpL+7GosBhitMuIF8
t1M8K5b/8ek0INg4dsuZN0KyVC6/qxuuhjMEH7lt9C0BVf/ek/pw1u3RWUEfeT2t
5YBBOWyW8emM7wssCo0mujlcj2rqu4qw4Mhkn8Ho0zD1rimur+lpQDY6/0D0ZA4E
rbg5yUQ2GFnGVV6UuYudgIlZFR0vo7bpqUXqkvzvfuwC+0NheLpqWHXCHaKhQ+4S
064tJUI9+QtZra/QEQjAqEju7alSaTZCtoonrFTLDia1dniwWw8v1jaZ9UfkySx6
NEDCC8l66ZPhuWiirmRXv/OQ7YO3lZf4A73SrnBZEMHjO9l/uC2eLRtPTpN/HLOf
xZFHmS2lyCpYZ3iZ1jzZQtOEzUwCAqie3aACn6ram54vfBoFafb3wmhlSklnott+
lp9XPTIt7fvtlcO1Y9srZ9RtlTjsVJiiFFGm+jWj+PgU/FjLNFnPJ+nOqtQcCJtJ
SsVo5YQ9N0QLumzjHbsFcSAgCa8lde3qNrAzG0wuuAtqFwaPX9YixASztFi4lYnQ
wCc+Oh3Kyh9VyJpwmuNQDq3r8TdT6nAonONcZWc/JwTEoEDltxVQCOiTDBQhQn2p
xj0Jzjo9jig4Jt7DFCh9KaFuDzrwmAZK/KcM3etcrYWTcZfHQV3pW0j1G/0kmhqN
n0bFd3Ggnzrmqxxt5MV8nwt1aKt6FVN5NoBzbJYJ80Bv2/ceBRfTmyG1avMkxUph
m7R+T7cmxyqkOUmWQMEuquH64UH/GI0EOCGWZnvNk3FBf+/SVV/HUSPl/MyU3/PK
6tD2qCNpAc17I4WiblHHyJEtSbJwa/664chT40yH0pM3GF9flhKOqfwCi/diKPlf
OmTISZkw6E9C/UKeSAgfd0rY+x6QH6aEBwSI6O1xeBZ/bkxfGYGHcwhCCg4P5Zb0
ebThEk4aX6151IHdgbN1kOLHqr0KT8cSs56HUgBCbeM3/sHZN1C2efqdo0LQ6VAh
2X5uyP1w3Jz/zAkjJN8BYOJvnwe27vgQ5u4MR7KaxQ439zAkWDREOxy3/Va9Tw4R
gYP4ZAZacctx9whgiMl42xS7ok37keKRftKRAlz4ZtB9Q6lmVMzLTb8uq3tQ1EOy
6R6ZW7dcpyrU9/1bXd0PJtB8FxuWz5J3F1XW5zB6zpk=
`protect END_PROTECTED
