`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AjfXP0hZQUettt6cdOqVpWn/QS36RyZfu1a0A01jP/aYthB9NBNGhgaimYIilHuV
1k4RGd2TgiK5KoizqQ7nwNgoNjx+X4jMGYzJEFMerIRuiFatjO10POOf5FF5RjxN
wgNmqNiszJ7GtcMiHkjaJNtadc+3hwo7UKvWo8Og6GNFNvuhZoO5BBzLY/yLBPan
Y1T06H1fVrUZL9HjRFz0lPC+grWjr44s8j0CJeGH4vqj8O8qn9H1gI4v7zswBumc
c/GgalUVh0rJpc7t3HLtHIU14Q5UCXLRav62ze8sw8w/gGNpwGB+6JgC2rYmHFCe
9UnMLOTfKFJjOclpY2BZToyh5ii5IgXzQeR62YrMM58HblSFa3lObLDk79oFi7xO
umVtmw+CFrnfVUIYuwCus0FGjuDwJipI7sOhw/XdesyZnjkiaXR/lK55XFNqWeuA
uO2R/ZzfarRGwGDmdgOTVQxwM594Qt8HkjGaP6sOLzw66a3FN5Vwq8ER7je/eQuD
x3tVD3CqzJPc1JuY39tHPTFmDuSKwNEb4pdliq3rSdTbmqvuaORZjoRy/BZ6mukV
ttyrlwyiC1qXxVluJ99i4Q==
`protect END_PROTECTED
