`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9e1D954Hy+hYACC42P/28CWdsUS0qXIS2fa2LY2h+jhGcfW+ZVAZr5k3cKBVYDcK
ZgCaValGb04x8bEMVsS1RuuwTaiJ2Bimf3UF9qbC3ydoIxz3UtD2uiG0lB5aH+LK
ZQ2tnH0tvbSKwBkfyI2gix/4J5fi9l7AX2PWT7PBF13DmPzhLmtktOHd44pghjQL
vDqC8EcH46LGcY4xsy82LUYV3XOhAWe1bQmBwx8rlhVx46fmJvib8HYPfAitrRzM
+tmXdA7yluAQuCkfe/8tD282nyWUaHHIJWGqa1L1A3uLequBulllBoP0mhch83JC
k9iq05Io0fL7jRGfBmvbzwwoWMV94f49PCy1vY7W7w8Tt4V9WsaNhdqt++c5vPrC
p/PvB/4uJEc8bIL87DkP2D3RuT1lvrVtXYTOn6uPvF1yusDqfN6ifhnjVuVXHBse
cgY8I6SXxThJn/nTudYfbzqe575COwxbC1zVtIgEfqmuiE2IbcVJIBJbvEpJUKcw
hIihjP6PUZOt7JrL2VpkTvOv88wOkRkcl9f6mtx54vgOWlqY9Vcyt6bac79w3w+1
+LFNzVK0HwfM5o9TlCeBgr6QSJ6tE+Qmj4HhYGE2A7MWYde4c523HH/pa9tgjFkD
3SfLTzgEiuoyDNGIpWUcKSKNpgAGYtbQExQa80iBxBOKFa7YtB0q9+4agi/XyRPg
PBjxdEch0zvjizghBxwSeKKs3/+Rt4kL0NswCv5mM64LqEerJZHE0H1JVGi16Baq
teCQgQPbAmXVbuPf9N0foFArUo3Qz2drqVJtr4EwVDLhc3TTUuaaD/8hpzsofJN8
ahN+FWKsjNUGkv3/8RJHKG9HIFhXpMboFlIc+3aE8M3GpDKywRqSch82T3/yTPob
Q+77hBxyqDUtJ+xwmLlnRYKpRI8xdDZFEmhs+EEI/07Z5l4sgRIyYPWx8ur8dhDj
gtIoCP44GpRoo3/fBRXvjS6AvpqgTUphadb9tbhVK7386T6cAIXI+OQinir9fSpN
Fj5CA7j6Av5syEadbmOQXvDdpU2AzUQNuZWtkOK8dE9ZxTNVNoIMDRXLW5o/aU+k
eyiAsclFIZ8UpdvU6VlvDd1leghgDKiRjMlbRfvBrC9uf7xjQniPTSLbJuTEfGji
tvJ2q/Tbe1v0aSzPKbO/umnTAZAfpTDqR3jVtn5ckGa40FMbiDilv1RA70ZZyaEs
B7p5s+B1mpCzeUzWS4xX+XzYCGTa9Uh7TGc/uTyCMdvJOlvoIV0mOwAvdW0aiIqT
ch2y5QxYIx4H3OjZuqE+aBMsFlFYOksLli13Oh30FFih8n2x8OXufHtSatN8V9Wk
65X9lRt4EET9UoXYDCfyvGbevq2k0kpG5y4Ck82P0qyaVKr8NM//JSlzAUWePjgX
rgf3aO8QdarJYBmn2STITiOdUCytZJV904XPmqRWgHBu14qxKVOhclduSLEjlcrF
MAKrxzZJ1nRcTZTPuEYPoSSXQ9W20XkUbTPUmGxckQx/IWze/D5NHBq7BcsqqaVz
75nOKPyYLm6ABxe0YTabAlARXdvon47jwoXf/4bNXCxk3A+9P+WHeyAG0aS/QcQZ
wCICiuMGIGyOVPY5a6uA7JCrTIb+wqxwcEjkdTcBbT3cHPO3m6n4kfblI0sGeB32
LDTS/CcUGvsg6s3VznYYsEP0Da0eA1IRCs2IU+6Dpy8S9Ot6N1s2e0mYiJEFPSyA
LhrDofqefVErBmXk2hyNS/OgaeI0ExNrvqXXwBPJvyLOiyr4Qp4rvcnfvMw676RL
vd4ZhG2ybDizZgQwk7b0PViVIRKtEWKtQyuP5AojY9L4Sun5DXVQtfAgbmFRon0c
xXZLslEYkeW7jjkobzPoa36h8xViYpBfIT6MALhsbjvrFxFcOvzbaWK/62TgqEZE
TtSMsRYX4X1uYFlVwLL0rc+5T9SfOUSbGwnHsssdCOf9q8wiOwE05h8bKiUEApyv
M/h7QmPyaOEcLwQdS30nI2uSADaNJOAgC1IewSL8XOnL/WR6bW2Ipo21oZSVzVJc
yHS0R5rQBW2sAYLYKKDl3a1tysi8leQ0NmlGqxQK0uAHE1vwavt8EdWeoq4/HEQf
L9833dZiXtWke+wxZ5WusA==
`protect END_PROTECTED
