`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQ4S6U9+rNULmkLCddY2txXsXHjAbsezrzIaLYwoG4MAssLwctqB7cPdmN7JT41N
VCMSh+8uVL9RbAH1ptjUBAqmI82F3oYAzV+oqodXnSic8MqtUpo5Nt78KVXAy/kQ
KLdJfuKTvApNUGf1SHZGdZ/KO3PjebEYxGF7LUk8rrets5orn5i0JfQTP4zXnH7a
jN9b01JVHiDax1vXmvJD49wCNuz64fuvX3/YbOTvk+1dTFcSWx345vEa2AUCS+Q6
2JLXhHyH318DDhVVX7CgGSoFxm3zNPeeEzvVVxkyiEV1s/PEjizZrPEC/ag5wtw+
VHVNgozQUfI7XXptfcktfU2bRkttR4qKVhTiPqGaMfvc1JAlsKOttUHIyW1lUMVt
`protect END_PROTECTED
