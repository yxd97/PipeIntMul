`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ITY2G+OtXENm3r8sxyjbO4afuVgIaEtXbmVnPZeUmJSeAhbQkKcJG6rz20mQohnM
Ilhf9nTkom23/LY9QJC3N2O3/FMc6blyTpUdNn5pu+BBGMb364QldAlc8gCv/9qN
apJ7bi2jqvEY3ZhZMgUdQOGNS7pLbboHRMrOxCmDDzQcWBHC3yjeR9vWTiHRPsqy
oWnEjQydhDnJk2ONbJBLDTIlDZ8clksdufSj7ZHOkNILqKEV6d8Xf2E4fsiPnLif
tiepdMR4RygbFgT1zt56cCNzySFAumBSKQjKlZDsoPM9bCS8ZX8ReQqd/LsbRSqf
8KyuaFLqCP2CK4yNw7+mU3Sbn3pRNarq+RmuUOYa7c33JxniHX83sPhqd01FCuxz
HfkCdSBquZ3rZhCajMjBNLY167L6DKYFXDKG+sGU1u0=
`protect END_PROTECTED
