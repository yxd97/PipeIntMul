`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYLbrp71LOskxuo+5HCO3ABcfFecc9UfuMFskz3IjjHL+aPdBZ8WuTXkIqeYmXRH
K0rW/G9rsFeVnIWbpntvNP3y30waWhlOJN6NPJowPJWJ43Z54r/96PRYKQ8WKzMH
kpRW48zj0y/Ow2srvie5kfiUHeWez8/6wJmJRtFnNnV54JrzNKbg3fXp0qc3eyoN
inRlUY/b0KglY34i0ux5lzkWNZjjdksagKEHOYbx3xzYVkLIQf6i2LYWEVJPU4Ko
cFlg8zrxV2T4rRJ2uhNFbCLz7CaokjD6xl69UOpOZH00z9nDgJeEU00frNPazg6m
TSR7uNWOVTAYoNmtizcKp+ZutGzLOQSRx2sAeuUcdxNPDBaC3gWuP98X6t6P0s1D
duLMsWoZAKJRMVkpI7CAIXS1IBZTllPvk600qEm7UgKfEqbCWNLw8L04U3QNk3RK
6TC8YSmXqjHZxKhXBI1J6sfPEVeddxu/hcEzgtffNtE=
`protect END_PROTECTED
