`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXvNCM4iu92zxotnPqaMeq+Ny59sBb6XwOvGhMbbPII0zlHCx6PjUt8FVzX1mqJq
AZWs/xicr6H4twZwnyyKUKCylk1HvCWgwj9EPEy1q1Ck/GI8827wx+C4RcOFnGOl
fHvtm+xKig3skLT2jVTwqGCYnIo5MgSG0ApXhJpDqBEVm58n8mzL5imMUDBQeGtj
sG33LJ67ma2qblLpnu3cbf8Je9r69R1w0muhn+WydVlTIQDysIAwT7rEXjh8ovKb
HBJH6KkvQIwOvSt9ZaTBntvVBG24HUvtx5A3dzT/Cf6AYBimDr2MVul9E/1rv81+
NKhnGrju7GTYPcUZgealWkQ+iiX5MsgtNoopWL9LqTAy3TwOmeU4jy5nq2SnxoxF
RjauNSCpsIPxHlHG2Lspj+myFhwQfCbntnVUwQlz8ReNn23YEjKIf7Tf7XDwBuuL
QKDmi4qlbie7b1cLOfecs9h3ddO/hIxsMCBAdYSoyASfO0tqzhpeCW+KkBNH09ed
gqS6WRFlOHvJqdjc4He39C6Qx/mMVPXwK6yozML/6SX/LLchKerJTu8mQvQruHg4
5zO78h7nl6yBjcqptYR9fa9Usbr3c1pW2tjSMGFWcMBbs8pXp51LQ/4qCXCBXWGK
ZAwEqmCJ80GYUfSkvvKyxDh8IUwjr8QmM1G3ZJ9hcImbun0aFyr8QOXKeUH7u5k/
Jj6EtW+IeQAFYASD6bGt542fbzX+K8L1o1H8+0LQ8wyPC49GQaFSg2kPrEHQpQ4H
nuVWfFs3QozQ2wtYdDWMlhM8UAod8Smxr0SgSis+4VE=
`protect END_PROTECTED
