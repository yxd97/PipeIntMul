`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WPj3ONdTRQZ3sCk0CkT9fd6YPAoLdBjxeijtbnQ7W+zKuAUSA4FZxEhdbrXzQacj
M/Bh+6oRpw50cb8BT9cl7VlejTOKxqSD2o6UFATh+FV7mc+GAY+lOIvlY270w4xz
g2/sDac0vvj4Mo9z5EPa7t6IpwB5IbS5l5Z6f+8C2syA8nWNGZHs2D7raFtbVt7X
U/doTTT1Q4MDGXraAVZ2cBdt5oY58Gpl0SQlJ2jbRcnkqDJqc7cqE4cApluiEweO
QNcZLzalHhhNn5ahcM3NaeMRcjUW072znyuWKSJNRfPHEq7knM9NFaoQP9fqQ6YI
ojBpQi1v0YVFvApEGeXMNVObK59vRzSEpNVQro0MTIH2tJm8JaFFaMFOAbma8AKp
vicOcv69ME1AcJRxBKVeaByINvZoAm31zOX2Th/3NN9WqDVS0/vaXE5FVwJeBTNm
R7HfUHxY1y16q1S22iVP9+WQ8foW+Sh2hTeK+GHF/kek2fQnGRB0RBgLApEl2wlL
4LZ32W1gdRSXM9fcbIEEBTGnht4nWxx/AK8OLM/U9l/EBFC34+chMRSAB4zXKDCc
2ZDOahYJFD5Hjat9Vx40tYlC+KWzxRKe6s1KSRtCDsrMR4BO3VDVFyKNVTr1j/as
ABaxQOaaXCC84IQPIoYV35eD+RblTegIC46I7NQJK14=
`protect END_PROTECTED
