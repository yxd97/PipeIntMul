`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y1aTHQ9I2FrBYlYgcSG7XAREffZ68GYkBxTZMfVcn93Qpp9OG75zQmzjoqDNpkC9
z8cvAldo8rzhR/vogshnc1mPcaUNQ01deOe5pG2BzWStFl/Ptq9gZM/h4KfCCMTp
O6jqB6EvjYps8KVRAOQkL6TCThNnjYVnVyzqnHpLdSOqFDh5qAs7HFYDI8GR/F6/
4QndHJR/Zjh6Q/AGpRCKkwjfwzdGAuLKo97kSKjerVliexI1sKGi4aeb3ZGhPG5Z
vKc05Uf7k8JctpWqqHWFrp7XYTomaT+plFaD50p737oPpVqKzjRBhB0nmlNaqX6i
wRIiSKgc2PCY/lO6ipRl7EPFlo44DR1k3sh5kCPA0o97hifqFzAxsVs8T800XeRT
w3aAFQ6BX7+sWR3qqRyckMdsJt52KCh3kMKR6v6Mr2lzJT+Z0i1TJ33fXjzYDgLM
2Wm7tja6UazNW8gDlN4ndDokIiAt7zatFA/ksdIPtfbNKVS8gNZrYcffo3Pa/1jk
laA2Ka9+q3Y8tgzTwpq6pnygzNtmJa3/DNBaN1yWF+Ho2D9Gh2nPg14BRNwbAGMZ
fzGiCHFZUEGOZ1vK3NPmoalcyuB13K5n8/748Om4/8aRDh+Sb8ul0PoCFN0VOzso
rDI9YaRKTy4CshpkUY/IHK7cdbyfFDsJL5jpJTG8TQ8T2VCO/tnfPSe5tWkpYWVD
fv1MtCRs1euY6rVpGEYjYZcozqoDJZ1E5evSuQGzuYDmzCW9+HjlZR/6Ia8vZ/VC
4TrSZjIkJjBZdBwh4sudm5FoYXORHkRMUMHlYTYnxyfbaGW4qvt+hwAbo63uGftz
4ev9XMDJz0t49NW9l0kJUTmvNdCvLY8fY84lzEo5pbKvoKYPYtx8rm6qg8m8tlgU
irP9n9ENhfvbA9cuZKry96arO4n1ZmJTHUheM1iHWcwAw445RGFyBCViqhOcsvJL
KPZdQi5OZfm3KMw1wKzy5rhE8qjFTtOAQHGWEL4Ho5KrF0xCQJgdXaBJBcHvVg7M
Hto7HvVuZgLpcfTidhoQwWmEzq/AtA9QICK6Pe9UV4zjUk7XydPJzXmq6IfFnAvT
1scbZ8+S5e9lBWBkhtrjgQcRxG/86VvOS0Hu+IxCnc6nPawucSU62054+G2ojMQD
L+fE6gsIRiNaXVvKdlro5eZejdRgt66bnFNtvqrqEUN3k6h1qWkslxb234nB9kwV
9VPu3pTPHK2Zc+LsZ+VJsrgurALNqfi4ecTl6vdN0uagC6uWEZnz0UjgFeYoqKM3
OwPOWMwjGGZ5COLJp+i5cusmgEPhsUs7YdYDTERPN/Rcli0o7cAunnnnhm8c/RYe
f4XPMcMX7D3qzCoxidAsTEepzlt1qtFFDW1nc/Qjgy+xJz7nEKjgYZ3WajUN1DwG
luN6tRHbvlH9tg1MhAtH1/IMddK1Q9dQV/4dMFtkL1+6HOXSGGmemTFOja3FfwjS
nTyN/tc5XrCB2yyrjv4brHEaRPUuZpn70/jA0qBhuGHd7sf7kuhcHbKufSvnSifS
ee/ODahQD3KXwAQHr1HPWAkn9G5LzOZRJDDRCsfzA4C+kwSR+mILL5lMYzcjKybO
YC8TQKlkLM17jQvjt3xnLlsVooiMGkfZDms4qq33TfXiGAU1VwSSW4XpOIqLrsxk
VgFsjUbCuflN+8wxa6u7yOqGca+MEQOtKV68wBllbxk=
`protect END_PROTECTED
