`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AqtcjJTdwTPB8Hi5tSSb5HRRBCvOvFYUvyPGYq1GQ6YxkcrY+BYc2kpVwBRvG4Mc
1GaQ7b9fuIWPTPT0Ul0djHxHSnBcafA1UFtlUQ+NTVM/HuAyGeGEJtPoCrp8upWq
iXEQiduMYua2v3MSltGWk4j4OVNKKFX2MrGo3BSO53ERinbfypc0eVmxLzBY2222
nGB2reg69De2pf5k5e0lkkMWqzbegUGKqKqXMO2uTXXIMvMfsOSN3/WTCvwTDhWb
84VUT4aYfKCNTQ29x0urqaqwOXZmzj+YeI8y9pGqvT0mLb938UNildVsCNHu0M41
yR4mIbKo9gpOVju/qGJBVzykVrMfDmJSTbzYM5EaJiyJyTfqZlpTvl0oUiFNrUAY
TfgUrueAXfbMAIuaaQMc6pbyl9xqJNjrl7OaeckqfA9aBrRoM4Sv2tkqCsYOTJou
cmzl2i8n9D9qzT0Ek7QZEzhECuurQpqw5+YSAH5Ke3ij9nWPSY5Vk8ZXTU7oEYNC
uOO+YVJWLGQfchXwtdSnMClXaSZCNyfpeyptAknX2HrVNkMQ9fxNGls0iINoUo9q
Ad4cHlsSuDXIVijQswBQuZ/vMuYglz7gBHFGf6dkpsvkLp23XkqBGIBNyWeu4ru2
tHgeeo39/3sxo5C+muTXEFTZjWTUgWgPSj8iPD/Bw+FWRYdBNbOroDwHLkc0Qes9
aq67MMYcnmZMo6nZnlJqIkUVwshUzObFTCtXI0lehh4uGAXnLpWKkdwGHeEEbrhc
EydM9tlI/LkHTsnnXB1FIUY1wvdmW8cwaBQCoh9y0pP73wSVAd6Z0Llk3IMIeob5
NfKRcfaW2gyBUck99Q1FVJW9Aha7YZlBflYj2PpLmsqHgI6NvLImLKLG8mT9pic9
DUKJOI2iNqHeSnYnyKogJGChjkLhzwbD4EMATcnFSLyREMV14+K1uKjYwyEEgawB
4szbrOClx9N4gkux3/PRei2LRzb/Bgin6/AFN++zVEWyZd9SmhA2Ynog4pnjFRR1
TlX2/TUC/erQyDZZjSS+z8/mprEHGDTSjWw+UJogwUmrVeSYpE1MXy27w3AY+UHL
GglRAPTieDXQtrL7Fgpg+fcVdS93ANbvZmAN7wxVrhj/ve2n4DjMa70RB9dxP9NF
P43M764C5qgAZe7BLRl5fF5UpnkBRWeN1z9OUBPWwAP6y7/PW2a4rMiHg2eWIhV9
VQ3jkHchGrO3Uz73aXMoc2seQIcHcHcsPFZg+lCQmX1DErL8Xty2hj/7muNJIR35
P9TVPHS+UVzqE4TjLGQxI2b2luc21QtzdIjbpjAgqkc0S9KPQKA9Awx0T/pn1KrC
bvZhk2Ng2l0ZTBZSHZg2QODfr6MjX1DjdFHFYy0sWCSN8rZe0kV8CR3OLG+W6DXo
ao4FSbrP+WYyoidjPbWJAiwmIQkCsw1rI9vsDxbwLwmB11VdTACnPWD5x2HLkvTD
Rs6PbXXgYi1E92yzbARTPgxveILAVNmHnq3BXHgftPdpODzivQEmdluVQK8/SgWa
HSluxzVnPUxtFUd5HPgh8hftxetPtfTl2K1UAmzM/B38y1TFCHQjd+c7x+8/6Yf7
D7IkkuGzIptneaEo3IIPYZJw4L+x2VkfDOctVwUtKND5qTqZjiHSGdKGqwwc8Q40
pMmTe13b+nLxnkAsL9DJ4aq1zpbWElmLKV1I2YrGBwzOXAXBJOnL5vb56+234Guz
NtKfP2mSrzTalGxgWQTK09JDFNm7E3SnCZCTZYyEzY+gn8oLB1eD7koZqS1Yr4xp
JY7oCve7zHPUQkVTY2zBk2d1OHQHwKe0PxxZSSx86WDPU61zqEFYPhjSmFPWI15W
9fyWE+i16x0idUVM2uyfLOtQqqGk0oBSUXu/woNyEOrjJ1AgTMdJ6C9XYnmUFUOa
L3gca1dGUtSJoqEHI0dpgxYBFkfQB9GcPRDeMGXS4bcoFLThH9tWRjsXLCUGr1rn
IYzqlOpZvCj6NFXzwbzzdCM4SUEbdUVn3q4e+1LWM4e0iyVCffIWS6LHFhZ3jXRD
ACL6j45CKyanCJDlX1CUhnX/PmZVHRTiqTLhLvJY7d3X9EvDtgkjsseB0XUkhCIB
yuw1jtLIhUl2JH008ITQhP5C6OT1wMZKXtQLXy55eOtiitGNMgq+QhLiEPB4j+OD
g13RmYrYobrpWDj/10l5U37F8aJoKPnh+NoUdtAykI5hfzIWLPdLQzCqiYt49Git
X0661qctm0QPvIcmyo0FwIWy3XFEHlMbI8yf58fUpFNGwsy0oqIUmYEuHz32d7eS
QJe6Yl5AXkayq0fp0uRLbQZ7C+OTcKKzeaI6CLMeLCyh3NhY5g9hAv5ec0kcD7xL
6qTUXNj5HBI57d5bzuAioWfpKFFmwj1UcrNIsl5vP0A8O2SS24YxzDpg5yJBcpN1
SHbKlTWD4WnVSeOm+kP6mlKzQWCGYjmdzw7zNio9j/Nl2p7c80oBsgYSLbba26RQ
ByKJBz3Hdh3WI7HyMsM/Yxlm/WKBRZxVVdjutWKRkD6tGgWD0D9rmsVwS1wqqIUb
WCXe2y5t9lV97X5jTkhe3jVg0C9QzGfdehePy6wULiT/kJ477sIe6V91YDO03gJj
47E6DbaQCkv1eVv5k8oBwu91Y3nkAxJBkh9p41kJIi75R961+tn+JhNj4uxGvkTs
NcbO9//QQyOHod4NSg09QRV4zL+45KEXDdjLnWEX5MJ+ALSdDr5Co+Rydj6DDzjt
piUGs62fC8dv44ZBL9V+TSB2zRV/SWd1URo7rccu+BbsYLQ7lgSHwO1FuKFaEAmN
a6ZJ8X+2pmt7i+IpfiyOq0xvFDW6d5uam4TfhdlT70RzPsd2V7sIftI2Lmj290rO
RMSOyj7aUeye6XyAmOG2/ys4WHN3nksSqLV/gP+tYGcekcS2LYmr9BXB3jo3BEC+
reks6dN7zdxh1H/Vwrul3RQUEgPoGqLh+jRlRWSCusnEy/sJ+146PUmWjgiF7kUy
k3Tudsc9tQiQc1Ah5H8KlSlBCOG7hj4fwV0UNoCZGmywGjXTU2syIqXjPu+Y+rns
ux2Fb3uL8/CGweRHTTL7lI+COsuPYhIIFtUb33/T8s9wnLENp+gHLr5mszMyKS5O
m1oJemGBs/Pus3Xs8j783ZJyAuD3w3e450cevGUpW/PLrjPDuASD46ep0nHrV3a4
lJB2p1tVRocheelUfII7GfCgcP87XLPlWcWx+34Ritpz83vPwsmokQAzCiA0J2vc
9RePZb9D8oJLZNFbHBfu39nRA4hlyVhprejRqRqhNsGnerprhf+etDCJ5bTbbrm0
4itWQxqVPwSvYv1pe26N/8miX+BFHzAL/qrlRGigsxc11uAR/8dWCcw9nCFlVq5M
sxw5l59yvPJPvfMBM8hxvkUyM9FJ9BfVZuDbOjizXGI=
`protect END_PROTECTED
