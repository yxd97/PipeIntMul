`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXK2OXNYSPvu8UYi7Ydv8c/XRvW8a0LVuZZCeB68Ew89EnoDRrmYxZH5NukF0nS3
jHPQsMvrmBWoBjQ29abAZIYOFyJAsoCKp9HRLVPBJbdlJaf6aCtIaGxBCIOBgQcH
faaPEVpM37VbuD82idI5WvU31vktFdkYuax46Qsc3HWNXayNu2MEXS7Kk2BW4eXa
v92T5CnkSgSMUHxTBHu6yzhvth+FXrJxhXdvPJ5HCkvA9rB4YhplBgX0OlphKFfz
aLuCPf9QVM0YeWLkcNNuieU4aSX2hc5rWeiUTm18WElAbJrQ8gUXbi1A/d5WOaBo
w+N7kaprCd1AMwvPcEZWyvvzpn2Ow7xjCf1QogDbIK2LL6Csq20/fjbhQ9he11be
sTiF85524jlMWsOQIHWTD4MSGkpVJoHjNTjlQIwpoiKEL08bkY/HBdIDhlXFp7Qn
zkj4aOi5OaWIJH1D2ACf4lNqxPHH/ET1+YCuT6A8i4U=
`protect END_PROTECTED
