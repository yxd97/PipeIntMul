`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/LwI8G9w7GkyV02elGighW7kfRpSCUcQAmdDgtpq1kR4StUxSCUmBEDKe/jAQ8S
R9VKj2zNK83xEuc4Fh0v8E1UbfNA2EM+DUO3BQdBqexaIP32Ht5RKoHFtQaKSgO1
ptMTwbwBGU25TNPVbN4WzL9EFU8KDGm2VQVvZW/sw9BOwxrKtvUYFEsBK0mgo92d
rMRcsx+qUvM/INtqUyD6nDwj10L5qbPiGb/1yKznjgvlKp3/9/G1VPYCnT8qRo4v
oGMuhPrBosGavxulhSM4yNTwqtqxa0ZqkXtwbFevtf50mc0SXlh0/0hP2qnyExXK
Y9AUqqUoJxm67ptrpp/SOA==
`protect END_PROTECTED
