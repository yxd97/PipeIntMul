`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6YaI614InJPIlcD4DyEGFoz0DctCSP1lYM4dW8GvRW//sNvqjqxSbK52vdzsP4X7
8JLezsQocTQLys3jCsOwjjuIC4JHNrpFzhwIYzYEO9tyZImL9F7v5wbcLqdEGzij
c2fYhiYFoNpB82aj3W/YC8rTDRLspK83lOlck4dq9X7csmSLbgwRAomW5ruDN8lU
2ESvdeybj8SCv8nYFEg2ECF9asqgKuM80oO250ENJ/Oz3948GnQI4mdIOte1U1QX
5taehlK9S5o8YDgrzKAiwZNSHixwNT7Dh/wOK7FnX80gBpo8mm6Q3Ncb0ep7+cT7
ByqKhBuia1VzzeuI6DOW/qiPvjD7CaP/9DVuDVKo2mPKF1P4FHOe2SprgQdUaPRr
k5CW9MtIHV7/hwqSOZEF0JJm2EAwa7SZ5vkEKgHzNUkuorWqoEHman60Gkp12Sja
`protect END_PROTECTED
