`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58Zhm2UyoiC1LFOjdIlQ9IW4xRGeBohgSacgx/NYn5+EYIqUaFAjV6IVNcq+UGQG
uO43Va9PYfToGX6SEOjbP6l6UW6rcxpdpI4LInO69OUDJgF8rZdQ+di0U7Sz5y3j
vKmdKIpvHt86y8Hh9Frw5p30hd15k0uvJN3xLfOxCdfOGjvQZoZthnyZIeQtoLbD
+rmOfHK7LnOybrsll5wfZw5Ks3gtylTX8sczji1sXnkMbvoSpCurhnbZEcolldMa
0nnGJOLm5ehUaKlEBjLybmxyFxAaDzl/ZIAVwQ7qCuJ6bpwRhx7HV+42blIiaJoz
mHJKjpbd/mzBIGwhQbj+KxnFN6kgMOREeK4yOtDrenIr2mlQLWTv1t9Jd0t9U9LW
tfxd9KSk6ERPIkvbjaSQEgxepGAhVVCGHG5JKR8jji7Y+lbqhn8M48GKVMShOg6w
DqpJN9c0UEPDO2crxudeexU1RXGJ5rliUhzuH/oMV3Ba8WWLO6GseqX6kocbz0HD
Qc4oUR4iXZmaZIbGSXq7rW3MHELUi3Xq2Ghoq1Hh5iEJHdc7fwwC2aMU8hsLZvEy
fCyhdDn/Hh3dEpg5DOCj1FxzDhhlRJaMEabZgN5sVYsNPBtD2J7iolKbCImbpNmV
E+fBK3NRVxIqJBQuPRxmx+6f/EQIXuCki1HNoDX74ZEmgyF1WRQxEl1c5DT/S0aB
qV9UDAck9l0XyA6wXS3GqY1IkusbYblKUkirzRlE1e8cW65ZOOFjLiE35SDjxEJ4
`protect END_PROTECTED
