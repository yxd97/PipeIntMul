`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1zNIOvx4AsYlBMisi2dJCcUhjSi6jYWBWgJR8SbMXoMycP/HIpnHZGMXJzax2siZ
hFsHkJ7unkuqKk1lpc/Z6kF+bzhYFQId8vzKTT1okdIxjzyJ6Xs9Od2crWguSddF
U/fRnay9ooLiLnsQsmsqB42O3yasjIGfGjjHnijm8FLF9Mf12HPiueq0fjovCP2O
8F33BtZniZjkytMhBwR3enllKqFo23uz34apMTo9r5BfOtAS0beaQJQ28s7RYj/r
k+LXQYv4SI8ZBLCRjwiRlu4u2HnClf4b1tGbr2cQVM0=
`protect END_PROTECTED
