`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPSIQmvEfnplLySmklMWAH3c6l3TrFn4/K/HTIIvzpZBstAkDgChcnRIp2nMqMlZ
AjeqQ0L0up8qlJlgfDYbuVQt3/G0xWxSquS9641kLBvnqeRRN9utGQgG/TjNPiQJ
dCYW93n+Zt2cKLEjPC7MeU1CFuYVAWih4+5LOAA15Eim86XHaG+ymX0Y6jD3wwLv
AyH99uanfvQXfViG2M2PAM8edywEH1bLLrTaEJRSqWA8/Mmf8+qQlZLJEmNrwAYQ
EYog6hq6sdo2e3xntbrzHosa57jtrcafGsWhBUxO0tnEgusJK59woGLHZN8r14HS
Pncy0ksRqz7PBVTNqpYopsQajNy7qrgglB/i5DbjxVzZ3TIsM7AhyHZmPenOyQxt
z47tnGXYHGEX9GlCXW8ndtuvSW8AUZZGz+su3/OjOMFRYJHJmthWrS/QwoRygwbE
`protect END_PROTECTED
