`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djJV5VSfr1LFaix2G7cShJUhpdxv2T/4LeIqczp/efJK8MVuQ8yZLqCY51bYvhnW
5drErgQom3deKu32dgkKd1/cpVKASUKbAFJWkJ/P/qY4oXnCaoBStrjX2z08rg+n
Fo1ebZ/GYXSScgXnLXgEPtOePXdTboOwiQ1/vhYvbEiPsz9P0TjpheLffeUqw/Ft
nnt5blWPsbX13rJOuoCjiGl34xMbeaLqSOV7kvUNuCD4jJykUSRP7CcKOSKfMIIb
SPh4cdUUWR+H5aNS09TJy/baEwW+WGc81wtLLnTfRvs=
`protect END_PROTECTED
