`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mJedqt6MZOhEt+ArZ4Ut9ZNuGFSY8BfSFcOQwQjvceg3NCW2sS72OPn0cUFTzCMQ
7YUEqYBst+cmEg9NMvZpSFHC6qY2RRg5746heL/i/miKo/nLt20JAVXVwqwbdRbM
LsnqsI8ED+NFE93fwOFvFMgK2qLTxT5rY9zMJDT8Xidej++daGvq6w/oOhBfgQyz
SLjpbFgTjF/+q5JUBws5WFRw8+DJofGKbE+75NdnrddG5LCwjaOOhOT1erDl7HRO
ZpviSNC38cd9Iakpdz5fF6moXfSi5LSZ0U5gdC7eUFyQZzKPiSFtZFrWenWuAjih
VFzw/nMhnosvoEvnVQoDRQPEAvITyiO02b8z2D01/xmrOlFYLG0UgYQFfe0xErMg
PCXoSJ8eql8VlrkeRmsC0/waNCwRl6eqnS1krXLrAjpWAI6DFCTH1wjG5izxx4CC
`protect END_PROTECTED
