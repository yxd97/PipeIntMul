`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6V4JOu6ETDO/wCaZKF2JVZiZguQvV3O0uBT7jUeXw6GMVFYbShgA5CcOFA6sj3i6
QkmtndkW995Lhm7tyiDywodQL/ly/Biq7CCKg73VBSJo+dMqiWWxuNs/coww6rTI
BnC765Sg2nf41/7vn74cMVcpziYruKJt5v6m4M4S8N7BzoYUrhxtMSKooWaJAJ6Q
8DS2c0tq1l+P2HLfXJfM0W6dPHX4PJKKAUx+UQYYN4Vb/RxmvdfSVaJVIWWXou/M
x14J4u4Xwh26nCfQkKad63xCNKYHT5Wz2OBUpvP95aPfft7qv2zEpq6PdV5H47MZ
tTaM83gbCeNCYuCI0B8Mq9FhDyKxGM8rdn/l4SQfy/sVZvoInOJSR2np2/uyzHBP
ZTLnIxJfVrcWXwxLH9coiRKD60fNZ1xh3sDSUKvD1e6GVVoqgKXa73qSC/ER2nhJ
eHtOq6Xy9JXUYbRj7IRX/21HI+oYdd/qOXQRFumWWZyzuziRdWMqi2A92H43i2ED
zYfN3xcbY4+60qfnuvBF1g==
`protect END_PROTECTED
