`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GcEN9HTfCdWs/nNRTwkGG5cA/lI9krRVW6o7kMkgZhRsvqRpg3NlWO6TO+i6enLY
8xTUdez5X4Yv4EbMvv6oXXzeo9E0BhgXRlhpCcXXuJQ3Cf21WRjNLADflw0MW+6p
uEkjbHwBEw3ISIKOXUSlhEhIWHcghxoq63ZwhrzliOpqzgZShLtNFiTSQJ5Ma6s+
i8SSs2VWRBjKGWBa8dGMM9OLDuVjjWF2myobQwVpQ9f1J7Gw1s2JGtpmjea2KiRw
12EvRv/88MW6LWBV6Mw5coGXqa3aRJfq9czdZ897pXGbRszv5pJyNpUtLGUhgot2
gWox6LjNcMsaqQqhBteeKSTxunEMg/EsJ9lfSTrkyYc=
`protect END_PROTECTED
