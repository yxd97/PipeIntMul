`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cQvtfGc6nWN74ffkw5fj3pOqo2tQFBQKg+S3Qb8zkldkB5PBzA+1m/XF1hwK1tpP
db1H/hKIb3OIPJujIoX7z1UQK9aexy7cnSh4TLhE6KPM7L3FN9NhEJsH8kmUx+JL
Ur18vLMiYdMCUYPhtvQaPxOUMH9nVfCofl5kWG8MgyS5hD/MsjvryDqq2+Z+3UCL
dgDxXSnrjnHXlWpTjabPwUIsZahY7g7B2ATCjNYAX3bVOEBE1485B+gZl6sBf/4G
Bh7Eve4J2/BHyw3DExw5cjFCK+cVyp7JiF1iXsmUUnhmbJ4zpJdlb92w4tBO3im/
MWn5Pa/ZQ+RIsZOSXKtq7WlGcyQG7uWJuJvY+z1VoVbH0eUz+knOCEN4bSOb6pWn
vIe/OTKFRZ/lK4VP9JMA3LN4pKv8Ejpw2P7yL32RdLrXhDuxYXvl63zm0a+EUSXV
gypJDn2cyD2FlENv7ni7xe6lgt9cJJ7/B0O/Ui29+RJCjbJYuqtRMdO/qC5XUUFX
C/RJodR1bjhmOajL5QJZUQ==
`protect END_PROTECTED
