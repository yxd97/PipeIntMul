`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UwCM50k0jQmMYUA8EivwTHh7x5PKFHj0b1hfZI8jZkz5OJPBTUlvMzdzGRM3yfcJ
huigWnqmW2SmHFLDaS8QdP6D58jGgvphGnsQ60ic6dzGZnQqZEbvBdnmr7Pq2Yh2
G9dQARUNyZKoXFQfXyksJC/40vetrypsBJhibriyWJhSiaCnAVHD9iioLT0klIM/
4HwIAlKn/g0/tdKIww2VYl24LFs3YFF1ASuXHE6/eoQM8VjtF0pPn9TWALnFCjZn
fMGB1X2WOzkdW6ElyTGu940AfZN2KSjPB/lRx+yOh4YpDCm7BuTS50gL1hiC0NlV
dzpDOU1sfnNVj62lgxk1qxEGgF8/kQR/3dbVf+008Y5MaA7FZN3mHCrw4sEOeX65
g7dcUDpF/Ju1hnSDz67aDw==
`protect END_PROTECTED
