`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ijuUL9AwKFF45I8bzkcV+DKYV1Nhw6bCc0Ol2GcYHhqkI3dt6fJmnFrxIdL5GnOt
2A0DJ6cs8m5mRdu6ZAA5q9c+CnqC49XnKMSqgFGebpFH0n1uYRdsD2tR1DGUpC/m
qVcUNcXdw6L17AQIqr5tyotrtNe7HNUsdWxSPttW8bstm+wyUGH9YBBQmIbwymL4
32U/Ij2vXWnWnKdG+rhM0yns5lBglrDc2tdoXUgbEB7jVVpq7JD/3N9t8csvgKNw
KXQFIzcegJpuv1qr+nZ5xsuimnqB85UblbPfazNUfIMGnaLjaZqFnlUmJvJ1JdTl
z9UAfLFHXmg8L/vrrQnWcYhsgHwhdUhWeQunavpgvUfl3bGo6+Pgx2NDQJNFvJtq
w5oe5QgC8XnG/lDdhRyB9FfUA9gS4DsjjMjnDy4gQyfKeQBdFBTDGPIVsicV8ZqZ
vRu0owVwRIOVWQZAdp4MefuXfEv0PNVYfzfIJ1D1cID2wsYGvA4b5i2DIC9B9XVz
DAKYC8Gf+Vg+TLtWi0YQupzPRe4LRhQyXOBUoIKDt9K4idD3zRbjdqqQqsw6KElo
JWUbRtZwme/SzwhlF+on8BJnaQaH734j5iYj7ybh8adb5Z3KFZOGOlu+PXXppgVH
zDdmLXQfnLLZ11nc9FaW8p46AeROsdlq9e960pyYKM5Y1zZQSkfiEuJQghMksuJQ
87yThG19oy0tQAaJ3dXbOka7fnkD3Q5dbW+2p/W/ATL2B9GPDVI3C6HFF5Fuqz9V
o9APo+YWRXeiTStfuSf56+St2MlV5eteRbuZ509PK0DYlD1mLZPTiw6BlMDfC78T
NzxvuXHQHWJ5tuZsfAAysCrPHhWMIIO9rYFhiHHRWOCpOw9qehx009iLbd8cXvwp
2TjWc7L8xB2w5wA0W7G/F6O9pjAc0Imdu+8uBIaR6vtmXZ7bmTaCCGaRpVDUNU+i
HQ5k2moasWCX84iieLJ5+bX6C32UMGO7ZnJK8TZaQGSbsOGsoYL1jxSn8lchueNl
6lmOlZd2YSu+zVCVprRvwtoEBkmUizvz99a0Wbu5jMCqr+xbODK54ijbmp8ibdvv
44DF28IGC+9gds0OklWQG/d17vUnCCw+KB1EM6YcH4bs4COgZauR47vR6CcdF/gO
wymeS5wW+rbHM2h4b7G7kEpB9dr9NcrXD/B4otzUMno9+o2Wa+82VPyTQ7TICmnY
giZKiYy5HjTnjsySH4uobNAG6Rm28yI2NQLERimWkQU1ecv4x+HEeOGwh88sUGoh
T5oe9JSzNGALUZsyC0+Vtpfo9Dgrwqa0ucNtYVRngU5DZJYgjFNGYtrYplBUy8T/
NO9b3lX2pHUsbYNAD1RQKRwkBBo1vfvUuqb1hSFlxSoY/NXWXBKLXOK1z4aUc4p/
GjACklLafg8nEtd+FIJATtw5UchcPDh5IcRHnP8v0Q9Y0v3k4JJxFu/B2qCCslXI
s4Tq6Y/YHUItDjh6hvSR/v+V48mILjJeQ1ZFM3+6DDC2jDMllB/mjQEBa8LBe1Aq
Ab/gDQ0aOS5bK7m5mDsmLXhXCJMAd2Oc2f9oNQl3l2lfmEIhHm2rsZ756xgXqzm6
wgl4uyp5J64L5gTJl5qvIyvuLVlcuN8Yh1uyE614AShtH/FX9OihhzkoU4DDMjMB
Z6QhAUdba6NOgZjpg3fxIZqSVmSl+CoFsDiQ4rKXc9rcX7sJcTtMXNDk4HxcU7dF
UWVUHJQ18r892+zUe1fEwbN1/TOHJWQLB3MgGJJ23K+yrthn2sfh8t+5vLu9HRIr
uO1In43RKPIAFOeF5BQ5kJ6oyAYaqbDC5+jvxsi8R8xakseU6pZ6O8wEx5Qo/ojE
anu/G1M9ukxgaZQ/Udy3Q9NubwfN+N2Y8BuFDdlgr4Hli/niwv4BW36LsQKo+3X1
AdYK5IOeYO8s5IsVZid8RDcftjL4X/5RTU4b7+BlLiypi0QZjrdizSo8MhC2dYjN
9EqunPEpUrx3TOFYaZh0YnDgBHUvbJU5e6KSrLilQnneDOfWqCB679/YYesGEOOH
tZsCJGB3hpWkWxiCC3CNupvxSui8vQS3/bLAopYbcSsqSwN9CttopVJYohGpq4Cd
kJMz+KMTXDddsG/Vf1+VUERl+XTPKP2zcVpzK8srGIi81k7L7ZE8x3se/zJoEZK4
kUPsnkuiSw9717IZEOfgIIB86WSr82Z/Kf3sUYp8DRgLgrLo3KBI2PY+ABxNjdtf
dtY6nm3M20vGuPjCb7+mAwpOt4eiw6ZeVeTsXCFxKekkgKXVzLlRYKKFjLabzB+Q
CjeaiPgqN5VquBXrW3j5eIdzVgXTmB9L3drHSvL2vuGIocfLy9h7k/S78trMA8MX
hcQe+4Ef8+ik7BJqfxpYbnnZRPhCTGScRUtTP+TrRsBw+CZEoXfdkqyVK9f29ZA7
ZG8icIt3M9GA/uO9tVnygpkaxf6jrIbJQ7rbCEpj+sTKlfZxGWSkRxsoqaMpU5h5
ybCyM6mixmVFQakGYXhQwFoQtSyQPKZ9z9iSDd1I7yRx/cxR0Bdth59IEeoxzwQt
sLZWcIulsIkIjWZPuC+PUChvuxWrBuhHUqG4fanjdJ96JfhnbS680aR2pFn4KBq/
eVoFXNGdDM47pjuvvzRHYKSnAVeUa8Uk9YSR3QeU/NEedQiIq7MlHMao+mSkNhsS
yeDYqE/m8XURB9k4ruRNpWfHrz8K2VnidRbZQbKiGp/9hM9g+YfU4e3ro0L6HOrP
DNO7NVI9ezKyVSfV72sNbdW0r5lE7tII+lOlmIUCaUvPK+wE6pp/9rpR1RARPB4g
jlEobWZpjA3GGkKVsULAB6BxPefxpDUyxpQLT0oJd25vSoP/pweLYZXf8q4PfBhl
zT7ounPEDXQCz7T96k9cGsv3du0ocIlekovaUKsQtHTZsS5dOjD3Izp2Fy2iu0Oi
OyC+lYPyVoT2zaD/LB08qNiNmhRVuguRzREgHuIf2NbdTvLynOP2UTAbCt9eaKhX
LoOKHKozw7UKTUzEjyTnBLeqyCiZj5fzvVh6/kFTWWOkHu/cZb4nGYkv0Cujm4xE
OZklfrqoihIObrrtAS2SqMUEEIiGE3jd7phHtmdaZc9Pnbv6cqCHRWMZFiOo+rtA
TCtYj9PYhiNwG1BF3sqlA28OHw9ikZXroQWOAm8fML3hjgVkTkU6BQIw8xl9ZS/x
5zKl0fysHyuXqRViSNnRLKiyrNtWKiS0Jgf34VvRaGPDhy1izTBvaxXCug1h/MhA
tX6756oVv/+COUsAB12B3ml8lgbLIwfePZTKWwK2OdrJWyAX164iXHRbQMKlbWze
SRd4ybUui/xpoMPvfuhb4BW5ME1RenwtKZ4dB0I26nVYjPyBX/8olvwI/HoYiDv1
Vjsj9ciW/B/aANHJj1edvKE+8DAHSJvAZEaA//DLNWkrGKnveoZ+WbPVzigkthgf
LqlSw66/39TTUVywRtjBEm8qoJ/xS9bTjB9aSBm85ENErtUukWLVr+Wuy7vR050S
va2yKx0X+zRpanmDwOrwfMKPeohC3rQaO8aUiS6ycrylhLJTl8Zkx74yao6CISRO
6Ai7D6gcA3GV1iKwqRootaiLF2OY2icyftUozkX8FIrbImXb/e3l2hCdMUBIVX1x
GPG29TrbKYOYcNCLkUQOtasqadH+4/Kmpx6f6RlK2PEszPqe62/y0rGMp9W3SB6u
lKb6zq+/VRYD8gplTiiSZb/hN5TUE/h9OEXPvDJ7fDRyrXDPkVhK6sIZgxE5PTPO
07cfn7Sp1MJbkaPkUapGCQwzFVHBNVlaZLemdv6D6p6BL3LmiXdLX/VCvwnzVZJn
9uesgQ1nzMbFYPHaj9kD2qA6BH7Kp6EnqiH2s25c4sAGRUwhRsXen5RoRG3YK5jv
I4rz0pPXlbMBBm39EHM883Vi4voTzHh53/aHl0wLyX3Ru551nfrxf1nubqCCLk5w
yjO6LaVUW2BKxhKOprB5i9yFCOn/XBwiQRUomJ2U3I8VlftjXMC3fEMRw9Ica5/d
z0CKfBorsmBpt3GxOm7OaXNcaM6o6K6CMsL+zInS78dAJTXBxSSm90PlkRcEp/9g
yDGzQNe4mBEbJADbKUmmTGmRjSsCqrqUznJo4Ye++MMFbRmx6we7qCkkRxWyvIeC
BzEuIS1v2C76MhbK9lUH1XHo5mbCgqzsgUDwHXAXcFwC0s2M/xiDcjaRM4EKbbar
T7TjTMGDb8ceSJC0PqQYrv5l3/GAz7THKiYD7SqyVsy9PPgiFRIm6PNzMT8IQgm/
EeyeTmz5xB3XEJ8ePqujabMI8GtvHawM4kQo+eT8qrQ5i8DVsWVT2s6Ul37/G/ZJ
GKKlVLX1jf/sVtZFGkcM9J1qhTRwQLrsDee0aXPdzibehOy8NsLHV4ErU2tXoUsX
bDy78VeLRPU2V0CXsjwaXZ3RhUKsbTii74L7sGuIlAeqOycT590b33/FnuQhvWdK
Ra0MkZ42/gR8JcD2nOcT50QI2cJkWXOrFGv4Vb6F/a/SmLdesj+VRJYv0D6PDJiC
2a8JBGBWQKhz+t+EW8Q21VA4umWOtxSc+c+Se6vpXCH25s5XSjACtQT5YqBpl8dK
4aJLcOHektOpvmwUu9Vz9ONZf1JbBAplGHX8ops80Rjkp5aCm3aFDGeuoHK25RiJ
OAi1L14Wih9bQ9IgLSpuriiRpZ8IfNEGna9sLZNgJqeMk0QcPoAtaud91A8odhcc
Une1sc+Lxundjzv+ltTu+dPyWHWEWCAj7kCveK0Va4OdVA83Ij+4pOVGmUrmbfFp
wWU5kXE/ecpTltgy2vgXidFXiLQyURuFfkiWaYKEOjL/D262+xuk5atuoZkAhdoi
32fc7TYD8MbQ8XfFqghSYV7zZGCX7W0EzReLnf/yNg5w5oGl69B2wWnCHF1sphTy
pLkOHcXYMDaSl2X3X46cuOtonwmg0vHgl553qjE2jzbbM0fzDd1eskzeov/lBU98
MCdqOZtOACmcyjoSwzlA+HnW/bGSFlaa7FAXzTRUm9LRTcEi2OGUGhs9DlE/xmTd
YJq9YEC0T6GZHq4+ZLJrFVFxtKJXxbDtGeWnMtTXtVQy/YRUSkBg4nOXJNbWoPfg
loVGwtw43Ibe/1UBd24nTZ4wtq4Sw254QOW4ZoO4hont84g5p1zBsGsbY0lwW9Qb
z7veUFpU6EukqKScIfPKwMtUhmFHfL6tUE/6AP5grqjMNVAoYDQ4aU2CE3vDC/QK
LbYOH1NuVEZWtAB3uBR/ArKTOQRlfgm38SJPiQSojey1YP/87x2p20oy7sjWv+aU
YTeTHxWlTf6w6/4LMOcIcatKb9KVnkGR/+RE5W2iFh21dFLCn+/ULFYadiq5ObV0
AwumBQLyVzftjN9wT82uHn5icOBw/4ameJNFQ3tIMO23ZaKw5dZ5734mJhVpbr03
vrEvIP/oBADhO3aQn4NuijI+yBy8sx7/FqRGyGD/+0xT5cGqTSloMAP+IQU4e4kN
iHIIWDvvRwVC2I9adEA9/oCJ6I6HMs0P9EM4hnW/HJMgzeZf0KmyKQ81M3KZ7z/k
xw1j+tsXmKgQVoYtVQq9uCx6y++aLUBHxZ05yOpcv1Jb9ejx0fhlmVIjmwULgB95
xnzE+t48rg+KU8GEzcRVp5r2XWYStko2c/zM7LVf+yaZgKZc/7mdQc6dubGCToIb
t8IjdRbKwQ3zykwYMOs5p4jsYomzImMyndDIBPdJ6ZREHIAY3imBSNKR2fFIzrPi
SA7EJUM+C1zuWnvEOXPIpETt3rizK/OIgVeZOrAT1HnxYiJIKVmjDK6QA4GLkgj1
RYxvT4edZAr/WV0fByr6eik1PgWEdoCCFFAsyVpvQ8krEcFtt+jv8YuIjKRhhePy
LmWmPNksf76Cfkx1thkfE8Ef0NnX9wKwQ2RS6AhTXrn/9fys7op0v58Fh0fAAtrr
Q1qKwwSbc/FByiMxrWZf8LXMtMRjej+2uAEHtpY58IwRbR9GFtVGxv3suIqLM24x
flxFuwiadjcXdZP8kETnxjOwjCsXQJgg81Kl/pJBUB+tagppk7cN8ejLBpw9yFrn
S+d9x8dLatIusH/TV/j/nMUgMG7NDeZkxUR0WwgZfhkARqPEC7NKzlGay8Jhs5KI
6WXpYM9L0Fo0DzjByP/JU5JhSExhUh9+5RLE7B98m2djb+UQ20aHuDUDs7sB9THB
u+5vd8CohP6KTII/Iknp55xAl7ucgsRDXsw5w3iKO3Ry294J1cgzdRk9q53U2slU
3uMia4IYIt094mrJDZyt8jqktYUA+jDVL1wQK0jI//Y=
`protect END_PROTECTED
