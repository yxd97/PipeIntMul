`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VF+htzUv++7o4gYA6rkqnd9LaLQjA6VlPhgLAp6CPEun8vcUOJlsySRKeV70l5+0
vPJ3BqdS72nhxWhhTK72IuvaMHMYpRpk9aXU7Pz8Rn2yaq31o0/ompK5YRZhfyBQ
ZY8oEwS1Y4kgabMVt7coyx87rdnnzOZZ5yu3sdVBaLTj+0aJBkxmGILvW9byg8iB
F8ts9zVNDUZn8hZ9Q4fvsW+/PZJC9qAEaMKPf7YEEJoc9Nn+TWRLrB/nM6AHpK8X
Xg61vstsQXnMyMvq+H7HZrGmMlFAiXjhfu+lEXDbMM81rsaKUpBDB0opwvt7XJhP
6hA2yDkA42IvssfbJ0QLpmqDxY0sRJqCi/3OsFdbv+V5FCjeqTUHBs3op5QrfkrS
KmVFHXjmKwbQypFF4CKGA44stq5PwfYuOoyA1I6ZG+vBOcL/+PhGlZLp/SDn/bpJ
H+MU8xYlb5gB5d6gKWKr3g==
`protect END_PROTECTED
