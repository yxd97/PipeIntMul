`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/0Njq6gZNEqJsOmhC37hANaXrSYtklRgToDZ3EGskTcdkNQhb9Pw4FzAlL7wpXzi
MJVPIG8/59VosT3doJLvU2LbxeeGwVJLnh14Z7loKtAK9rw1k7FoklXHDo5/67yz
/VD2z7+9cT02qc8+kiWGKgP3Qzd3PAjKHoVurRRX5zRFlzrGIzBJagPejqSXF0U5
K9S2zMNObkPcmrk3oFt6X0YuKjxdl/WUJWG6Mar4UQuLJRgpfQiJTtLH6mXZmQzQ
RR2pof9P4YsCU1SkVXXXuw==
`protect END_PROTECTED
