`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tnoo5OKC0LRZcxXolGg+/PFQ/Kp5Wv9jV2OW2Pl7F9yMwlHJ3Ah0vRzwOPfeqe7A
1l+k3tmiB9RQQdaUHBWiPT7Ox+E6TqeaDo5HTg1YfB+dDZIAKOuv00+rvqye7kVO
lW6BitZsk5vxDFYDjOpHTVxqwBA95RNT6kScX5ojYBv75zk+hlLM/+Yg2ih4YK//
BtO198sMp4FIW5xFi9d+tzuqUyVGll5E1RPxzuV/M+9JKMV7MLHgqLDLgdH6MK+L
GWZQB64Er5g2UcljZP+Hgsddpbtlsm41ezCufxyEdL3upva3T9ztHWjodS7od7vs
Unc5wz5VDNUyRhSmsTpRgA==
`protect END_PROTECTED
