`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CUc6hnC1v/JKMS3aTb2sBtFktXQtBtM2oaJmkVbXZZeSOlLFe0AyRhds5weP/u79
VNa8vdwsWajpMYjhIFUuRPdbZiiyLR3VotyZrcFgHGF1hSij9Bq09kRR3RcUPwBF
VWpflxhOaPAx4e7kj7HBKd0ZqTUDf9kOScHjXZFYjVUPgcTCF1VLkMAKbxZCUsH6
CD5eqpTjFij9GIfN0yJSW0/HVM1pVFd92aeNIKZgqPQxS6vRjmc47829Y892Hq1q
2BbtYRy04qebQ+o/OgVCEv+uEVk8Qz04pXyNqYi4/qNZwAzPg0ZJf4kGIiXpuUXg
UqkI6hY6XgqfjkENBAc057KZUfJuKkXNsukRS8hSgIpdtwjfac0WzzV3oWC39GFf
xlBdqbOaBBWxZi23STSStnCyIhDSjn3zVA8YfgEb44y/9YswwPLDuuxRV6kQqasF
5dpzU10RnvtatMyF0XTlvU1dOSO3u5m/u5lpExapWj2zbrz6IogAMcb6ByITYeC0
WTZHXJ5fS0Rm0xu1kqy1BTJa/lj1QWhSyXS7w3KU+3JNLuxZ0EJUFF4rXBGX8CEe
YOspW42t2sgydhUw84EpfsXjQKp+QsJNukdKdES9/bZHEq0ZWgftz/xzHdp45f/Q
r3CaIvgRsWoB57SP67plNUMR+Gkk8M7yvHz2jS05POS8GfC3kO44ZAV5oYTQU9t/
dT9SWZBvSTBJuTiE2BnzrKkDVjm7v4zZguNemvVpW4Q=
`protect END_PROTECTED
