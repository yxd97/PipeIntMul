`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0U3ioUUHCm7gmQPUBOI7a4q/DCfR37xsv+Ow1ZFozyOkkVjjoD1nAN6WxpbxY2ES
CJ2/b0o6ph336KGbNf63O/2oKsPKPVKWsOOZAI6RjW6EFPfMu0KhAIjMlhwtPd6r
5/+xiuZk1vOkSIdpBsnVtWKEJPa0+eEjcOF5gUt9iXZJFvZsdlhchjUxsaALnIzc
zFik0N6i278Q8xUDa+RY1yQv9p+vrPH+/BYuJUu5ibtsZdEorwZRLd1MQ30cF2S7
hLoZaxwJ3B/JbufDi/StO3RiY3HGs2o8Pbvu0CeGWlGlDuTC2cMAatixBDhoQwSB
C1QL4d0g4bdAbTk1/OIqu2/qGk+IfooU5tZzte+YQnVnFZrMKFJ0x8GQ76zAz93D
70rAh22AMvmzhLIkTs4pcK6mavzke4qd3CLxTwbScufnHrC9W7JxbosHKbSWBCIo
Mo651bUV2fi6Yd4GltzfcbpJYeDOfoaM668I00w5nDLWc3sDT6MdTEHvkzpSmHLO
RUtgSSD6BmtqoWpHZH+enlIZ6/NLLHvcEKsJfAOahBpJfhtSKNzkyBf11e7TQggf
oZmaLsmEVZ0R6xHevVEWHjZFOMikyIYYEBQ222UynOqpvZbPv97hqKqqljW+u2eo
rbouDGVTguneah2/1o8NBxChd7/mGxfaWBn6vsBo0Se2yDBD6T27antvC4gu0cos
z/klMC/x5CmAgraQAQxrZQ69fBejFns33PELUDWUuIEmsc8zy/DfvcNcBLaPAfHR
9NjjTtYpUHa0MlgwIRVPDm4v1LWJ+s1l+Vtb7UpoX9a/pFMO+wHp4dR+tloBv+do
oQwjnbOlHQdW9wXpU4sQz/kOhm1zbt3da1yQIGj0Yn/0cUvtmxjkhJ9rxaEjI+Xv
euVYSDIKMuDWMJ/cRe7lJ+vL0RFIAgfmJOgfJNQtkhlB4U0DFrWdJ9qBhzN4fQ+Z
HNPWT+LC325vo7GNjMC6huJTz8FnpgZ7lDLpb4rZQ+HSxKGhF6iM9Qakjxps60pB
sN7I89yAxal2Y3tGvUoGO9VDEKjjrG/JCZHZAuYjy1QynTbf9bS1xL3m2w0kIV9x
XrK/BZ7KRSBSxm/cqhwU23K5A34zy7hFI2oG8BCYlY9Jsfk7mYg34CKexZPmXyA7
CUjqhjIjEv3tpsrot1rIwlGSeFrBlDtLupDDGltlyqsBOsIepqKKM/ocUTwBWDFI
MswJDrWy6WAj7ySTAYaCS8KZ3Ol1lC+v5h+8coBBZLdmtyZJUha6f0lZV+azOuYG
AjOStCgiSEF0b5sgjgQnFtnw5XNJNO5iGIi6SkiTbAlBwwdP0dzP8vjSV0EORDBj
`protect END_PROTECTED
