`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xad2vHUQBXoBMPA2lZuBAvHrruJ6by+kYZEaD8KXVC44lB4yOx6oP3XNWwUzCED6
ewgu7AhnNoOqYbMK58f0QFCqU6AFUH6T7tOmBuU04FWN8S2BoFyhZDXFPKqbv+be
l+hhzXDq3QRapowCd+B9r3z8IYoS3Q6UwZCTzumT2qMhkcsaDxmxyC9y0iYxt0uE
Vdq342jAcs8uX79NcSjEL4fEKHpQESasCkw13c0/H8bIauzM/BwUmvTUT9nVUqLQ
NjoGXMaQlQYSc7+TiDs1uMva9vfKsUzYgOZiVv71oTnyyGr2R6PKPvzTEeAggtKu
AUoqFK53NxpoD7njEo3k5sFF86dh5nGlXl/f8foszQDa+EY/ifb2W4VY2QEuuaRw
IQzmOLOkf3MfEeCspyD55StB8/3IWEUNoB/I3+4uaE7/hHkhD1lEqpIxpj1NH7TA
ojTN+2oS81q+x5maJRNsHaUKJl3ACpxMvD2Zyooqkb4OiX7RMfZgOWKmUW+V58NO
fp88QHjNJvU4mbxdTkvnDfUBKxyO+GEzX3Cv9O/+0GHDdMJakrTeVMJoIx0iCPk3
2tN6oNmrS/6v61mB2OFCdFJ4+b7cIyF7UU1YARK6itDUBPMiwkzQLOVT65EisXdB
rOEXjVjm7r+dP52M7qxT86APwcr3BA5finwh+YbcTQAfTl4hFghtLwXBtgTJUm/N
lM0HxfXv+NDX1+rC5v/CNU6LWVqJo+9lirDmXuZdnR+fMh65eiyXrzunTLTV7yCT
DPWwPkH8/qvGJR3VVkFihL7Fs0tb+C5exotWomoz7lHxku2JDjcGoAdfxgDw1qI/
PRP+V5gmNZ3YrNM0CphEcrF1T+ZCHAG9T8A/vgYGLlcyZct4jCYgA8aX3JKUpwMf
DJ5DkWVJqlK0NaJ5GQm/lXmiMsF/NDap9IZJk0i6Me3cmqSYf/qQMGHrTejv4TNt
eYrpSq4RLdsgV71SJGw+sw==
`protect END_PROTECTED
