`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rhU1XtIz6GLXmGXkD1hHZSdcwi7lDttrVueS1EMwL/4neJB6QZcIDESgEdAvCG5k
8ujAx26g4hpB5E4q+Mkk1fVmUiluq7/cId9UD5BHtn/J7xPz1njR8cPfxVW0SLZj
WttGy2GGUiXMJkGOi7gWGm2OdU3WDBEyQrKagIlcfVdZUzMLu9sMm+bMFP8Cn5WH
WQ+i5+SZj06lOUwaOmrlnDSzZeQuQ+fpIANpjc1BphUn4efDtDQnVtalrAjbQVLQ
A+iV/DO7/CMZVDG1UWh/3VhgjBMfA4aVET6umQUUEE2GZ/KDkQ49jCDZu/kEk45V
zDHhUfM/dU9D8PyMzu5TBaTd36g0GfOMOL2E3igBoqnDfnLZWEc/I4prc0/gBEwE
+Iu/Uz8wYoEomolk/w5AHQN9OYtYGYadsRxc6tN/1d8820h+bm4Vha9/ZgSyk2C1
16xz+yFMS8/mpFkhqF+SLzYaqJA4IfHDeqmTf9URDjNvSpPMfSMynvn/OnmSyMCE
xt1pGLOPwCyNaqqHZwhBZf8z0K0TI+k90TspilTQ5rJs9gNnQn5nAkwYXctG/tJF
N5sqzMtKW4bAZ5h8h8w6R7xX8lEyiwrM0tTcMRMP9cQxuTvRDEj2MlAFWGeldaLu
k/FNoOk88lLgnwx14e7vHvTxtCzzSIs4LB/KVSIGORF7Dv4jkse/lZa2ZqIGFcge
848TDA1CWQd4tnNijykqYMZJApS2C+oj15VurlHI36fpGNwyUdf80lml9TGsG17z
H8QcGj4t/kM2PFJjhwXtjjCumFKlRdXeAbCOSmhxNI5e1ZiFm71WVbasyZuDeBh4
6qzTNsT17ci3qg0/T79kWB6OKJK+ZfZ0qxLyZZGdiGWVOjXpvf7nTdjv2SMoi51F
0WnEH1M5kx3NXzy69nwdGUhYsTrCRrQ8skk/YvsmuMAbrZUZ5Puw9l1Gfip1MSjl
lKMB2IylRh0LEY+kEnYhPzS1fEqSyihCUzBCHa9Fq5gGU4zyGsvFBicXCYyacmJp
7NkgWOvaWS6rCWk3K4FHek8xV4/0DTRWuw7Phr7oGAa4oA2pS28+Ph8Mxkt5SsyG
5YA6AXmsOtTyGg6VepFk5oHPDsZOboAtVRQI/yB7IzWAbPO0FKnmY6rMMCDZXTU/
Ksgz/vDGpzMNvnR8TtiibEPLJ8lXlCDi69pZ04WImuvFudgjhlHHfeFn9BQ0tKHY
oaCp99aJmFbKHfxD4bAQ+zhFjRkxJ7IMHFhvwpTIaxAkm4dGR5hXR7MQKyjJMwTA
mx6dYbPAoWYMRwfiy6N3gG3As/ZPe3r5BHuwBgaiI+lQ3BFT4Wxp5PjmByLkJeaV
nrpBAwXL6nzhTO74fHhwcXoikl4C+ES/iu4Pz2KkWbw5YORkMfisw7371CdCxla5
jPjIObcdQoc8haBLc/r5mmJoT594DH1q623s9+pBuNwwE3JYjsjNe8oPxCtxquEA
5WbO6aD+8SmG17Iou2ZHIcc8VHVER7KGocnJZft3mlHAXJoKuNVW7VmUFmU62OKm
RawflCD1vgdQYbDP/K6S09GLzqUuz+2teV5u03YGOB/qMikzNe097+otbDVucbvW
CbftDEz8jcyUNHyy8ojnh8+UjumFIpeBUwld0KVL0E86BfHQksHNHqTI+VSjZv2B
wDO8SyrqLfom49kpWf9BMOVK1YiIiUiJYXBtg1OuJqo6GQ/uk/8t2m/Qe8N26/VI
9FXaWCNq8O2n6KljSYVF4izmooUMZNaNje2I9cnSn4IOCMmhaMtLfMxyKse/9uYE
5SpY1xOyTAJs1m4zUSXXCQCHD9V4W08Q9szCm+tIecLxekVAOT0TgGDjteAKA+nf
HdAeIKSKHbmMmkad5wmVpV5C3WzIBGOud/Ed1uKmLC3p1dlELQymvX+xEUS80+uL
sE2gNzYfqwwJ9RDMXypKpPXGcYQYFQwG59oebLu5jdAGSzMBAvBQRIsywWerEs+u
5yuHwmjf+z37hjquW1GgBpPzJ6Jr1eOZyNz+BvdZs+LjzVbko38Loc8OGEaHPuzi
ZYXGmWK5PHF0RX7zsPl8KVrqkXDsYOnJ0/IctNCRywdKV2VXaoe1rM9/auST3mLn
jGUEh1F1mA55WkVPD/wG03eJ0cHSiblaHfwtLeGisq0Rkq9HMaAda0rUILbaQtoK
Qcb42Om8/j0W07uxyTrKMiCgkvbwJ+uniaCVomzNurW9lmWZQhkGm2EWGuEq1/BS
Q4SovGEy5uonNAMwRqMpJ5co8PrB8le8URABl94Yd8L6X7t77FLE5zxgmpMFY3/p
oUyis50DPG48prhiCQceJKWcfZR9tVZgMRJ5i/9bJIDOb8Wx82Q4Ojj9U7sOrR3c
gLoRkiEYTXTvGL8jeKNP1LIYBJo/hk7xk2sYR5UaUHiGN3UuWHFYRknzVWzRWDKk
B1DJWIvN5X00v8hg6LnLCrnfGX7XVW6eUTmu4rotZC/DJ7xck0jSLkysP4J6Tk6x
oIE4fo/oSZQIpxl5syVCaF8JxgsQX92wQeQuPIszoHpz+xjTRYN5DEa6Y/dKCKT2
kx2GYVQTS9Ks+gxDaoD1yvCqSt97wr6SyLLqwbhwiNfTKPrsbr/2bJzJjMcOUsiP
WXu6oFpCyRBsRz/Aag7uOSwVViVdscpd2D4qk/V0X3BvKz/B3R22DI4toNpUbG9I
mRqq4qNxvf1qe/v8fjQazoJlXBZyoTXXbukUB4sCOuGPMryXTxq4q2x/RiYraNPS
8zXnOb9kCpeO0duFAZXoubLxhLt0rj3/yftb/YLs/6IXPgpCANDCB1TsoB+XbDFz
Wa+UwlhOVXHrajT4wFDYM9699pLgSWIJqulPMoFQXEm04pU+OyTe+m2EhbIyA2+2
8sDH3TeHOwzGPU9zQvY72Q9/F30FZSH60UFKfI07b9QjIo5rQWP6iIf9vj//e+yY
leCmAumGp3g0+POAyXJP5Mqw+yjbsbMn3/1giR/Bph2oSZmy5udzBoNLz14gEo+1
6DdYJBR32R5VPUcosbIxAwmXhMqzg+FcfaKT2VfXJlm7LJxFgFieUiSKbBYMigA+
pCKK/LZCsHtvaNDujj5H48f1zF9lFVbTmtOmdjkzxZq/1bNSLo/4/9qLp+Poj0Tm
8PY1B8oCgfSnKEYpZZf2Cle+kCQmO2Ba31516umaLK3fh/uy5C0ZXvMGqyhjdu5v
5/g1KKO2JFzh0J41rf4PJyvRj3Cj5ncPPwzBRVI7f0qXkJheODo7cB2m9YFk2vuz
wPehTNfFfiMZA9Dtvyru6SfzfvnTWY53TTRs7pKlrRKL2/NO41sJZKb3Wu0HytgK
hYOSmzXJE8r32X9BEkTWR6sA51Q+Jt5hZ/VNX7avQl9hn0bcVnTbHmGD3HnIhAmz
O1giMG0UNHhGWLSQtgakEDU8/u1DrV6GeZcKUP32BwJ1TyZdCetuesWl4/arDcDx
wSezG8pV3FhsGZKp9J4D/kBkse3QhYcXBas9pF/XbZyABnaunRPFLIqCqrThzRYO
VxvyBlNGNnN7QwxNfmenl9lYXnRmY92mPg3S2bLha9hK4apmeIvFhj+7hwaG1Xxz
XoCBF/egwvHCqZmmZ+JJc8uUxVZ7C7TQyrVrpws1Qlt6aUcEgTxAwPtfG947+TA8
f50X2GKGXUuqntPRYXuQGyieKUtF7WyL9tc4e2AZYN3AW4vtPgz12W+PghBCsEW0
ry8sVlQi1nMcgCJ5/yMWInAQNTXJddwErVc6Snm6Zs9YPqMZwt+n+mogmZ3GAAcG
oqMOqEujAuj0Snrd8jmibo8bEwdbsYa+0ISDNs885vVEqCXsoKeUzGIcICHaZDXH
MvRiP1Dk2Qxtw1ZxbaqR3GDNHyiMw7xqJVkPchmWNrOsD4oCrJKa8qX8kWCNt0WQ
72r0Ve2YFiVfKI7HgunLvD8SoWPVhHgPhYGeTGrWFKQ+JWHqZ5ts9ELvB+yfm5CK
vleg8oYvOgHZOwvwB4jl3z0Tt+QZCkjrQfUNT4N9v95llDwhVrBKYbuyf7oxeuWc
+xnwY3OUThuPywWaGhE3N8XIFRMe0KfXpg5Xl5xeS4GPP341hUiL/8nST311fGKw
YdP19ETcB1f8vnUsMC4yJPp23NVmAwGaiqu4UjgqQaxI82amsxa9qge8MPYbbgVc
1V0+NfZkCGaxTxCoIk/7cpy2/fIJWHOXiV/0Ps/mQlmc82CENXQ4vSq95eKuMaJj
5pi2Gf1b9/OmvN7fImtqzdDOFnzvxqThHzaPpeQwdj5c2VAna9dHIwvl6ojhRN69
mkml634mAs6QMPiX2ne1LG2szK5aGevVCF3zEZaRFMBh53GzjbjfcipmRGw61Rlz
SMAYBg1Yu/lnlWfjp92bnS5xj49xRuN3VdEGbavBhZcGzFauQbbM8SIFbdsFCL3t
eLWcz9UyKKSSpFdVeGPSIY9lOaBq0BpE0K1nq4xmo2MI7yo559gvO5WMtwUqPyMA
MsjxDojbNo/OEyheHqOSTiQcKQdE0ulZMU2cY7/mHEV9KxOVHGYXhjR/3ax+xH64
B8EeoCOGhJwH4wMhpURb+Z20fFi4nnp1I6GrimG3Am1BZmhUfz9WRdHOmZGaYnK0
884LGpOZQ2YiOJ98WWMRYptrpjutd5QUij9WHPDu9QcwUibZ9KoVAivN1LKy3Rbo
dkPU/fgxYcSRIPNx/rl4/+jRVjMxjfOkchGGRl/UjXjjnVL9rJJw1KW0fDG38ECC
B9wi10q8U4KVQUDh38ufLCYWaml44AfVxlqrRUIW06LnRgM3l0eOn+2drk0FAH4Q
JLrWuzeYDk5LTV+5PzPJXAaFvn6yUkSK7Ps+CszDc1kvtHEfCDcLfVa/W2YFKbWy
J1xsQonfPmpA40W/g7e+iSYn6R4GongwODJeKuNLRWtMZI2lTl10+561JNiJum80
mCr7WdSe99rydlm5AaLhEIiF4uYzYYPLbbgUn9gdUkx/69mVNRpO2kyju1zxShlQ
F8l/o0GQNv0jx9aoHaMgDNrjaEEYHzFUGFLZAjAiRw2q5zfPejFYQngS41S46lih
uZS1nkQqFJ44LDv+qPU2mv6mKw9MH5SD4VW6V41+ipLcA0oVwkkvqiy5hSeqBFbf
CeUYAEolK0/y6DZ/Sh4OPCKKpPjYMi4XmREbNLeK/NvmmDQB700XH2p0a2HVDzZ+
LQIeDAmrY+7ics1lNokpM98Y7uq1CZz8dgcJGq+lpeE0PieI1I6MQmlSxW9Lpq2r
rfhiAczreyWkBKVEAxOMpqpXRPsjes9TfaPoa+ZPCNlDRQoNIqDNMfj/yfMuBWrH
16j2uCePkFruz/1vS4RXDFQHQfBwk7AnE/9YoM/hThjVT5yAcK0ZGFX6FhdDQ20Q
lHDLpkJSD/J1p9LSvJpwrxTQe+R2HYVq49xu4eAb0eKhyMXI3za1Sh9ccJmNUJwY
4N2Ez2020IdDtB/LrCQWX3YMuKShRxarIfuHx8hX51NLCuxM7QROxOvPeumctUeh
1NvBnJOM3tgIgS5DVfvpRvbTIrp62EMVINgzHc+kP8csx9sRSNxUTDmsu5DPQl79
J+QRT3srsCc2DW2hlqzK6oPNWW9uFwQA30olhqeq6Z9svLE7syFZMmu3G1jjcwp3
QB6c/V7HzTh/GWEetb/IpJ8h3EAleR7VOQTvMSiJRrNY1WPPHt9j3xOpw1Xjpk9i
Mx/mR1fkO/O1o5yTC+i1xB7yAT19HFpfgmwGTZyguO82RLml07R7maMTZbt62u5q
Ek+gE72Rkxhx6+k3MZN0HmnSz9V7nAQRfrJtWANp7F/Oyta6y3l8CsJb4D1kTTXB
/vWdR/+AqgkFhMVR3phwhcFt5wpXAudV5kLtWdT/WHDBAqcefpeWJXMUgEoaZmMJ
kyccfhrh+rHXTFnLA+vvwTINVvUhqnLKTDv8F3yTzLDjqOoaFkV07kqbXMEZ1OXv
RTyRXFqfqX57OutODg2j89rfs909wTH3GGqZ/9yP0TRJlu6ISWF7Kqa0nwntzgKg
RHuhBlQejZQryRb/q9d03/2V9csXP97aKfXGcxlv9ZP2wKb1nyKZhOt272NQVf8k
Kf8asPsnPR3hlDzRiUaZ7cviq03bRo21RfSJeDTF/4+s+34fQ8MjaW8ws3xowQK+
TWktHlHt8O2+w+aZtTdVQKGTof0OdFm8zaN0MCyIp2RerqLdUufmxIXFd+RlBJSM
nAX9f9ZC4E97/J7bP+RFQMtgkZRrhyX7iTf0sr9UwC1QlR9MxNwZNfuBU0g9gwnk
4u05W1+pwAbWMDZYfu7Yf3gbUo8rwT5Lclwx4IiQpcI+xhAlRHlJmv8A0QnC46DJ
DK4D1/YUNcOGiXjHJ6IO+lauM43hPhQqzBLlRs3eFtB55ial9jUEKhXoBQ8ufs/Q
Em6Zg3YwqHxAwgOzMISDoxcj1yHhDxxFmeYfqbJdrGKFa298sV2586Wrnje+rTRS
UNLoe1OokOtv1VKu1TaWum3mx9CMZhDc7CaMiCucrs68lIJ2qY/6PDbsuaIsWHno
K2uBGYm2BPP14S4fGeOCYO6HQLEkJsfo/ZLdmx1EebHs/4KlwuuX2KLDxXUyJ7bL
BrvrT5ia7lHaJuTj3HoGjS1p6qLzlJtNzn+Uo2a6GZJ9gwC3lzghUpS0iK5j5U3+
ZzagleOPQY5kOPkAZrnvVPD41+JnGdeIS0jC9Hx6ZDOVT2PHU4YfKjTd/q/Ss52N
gl1n+rMNGmqhXiKi0bzM979WGuLwhWtGXVdzybMc8xoIWQpl5nx6mHzM0bLQP1oW
SixUUvrkVTUGMNubmcN+4LCojdD0NZTR2OXsV4DqfD6kWhC9PqXNhSMqNxTPELeF
oeEopSUKEvj1qD5EaDFNFZE516hA9qFQQtgYBwjR13EaHio4NBObbwuh2sZ8sV+c
ySyCfNQpbufemYsmZAjiRNHBTxmDAWaXG8sB9xZeq6U2rOD1n6spd3UJWDA5TXE2
OWXj9xK6DXoq1K0lm+dd+rP56u6ARe4TVNEfBgkf01axZQptty5t/g2Tj0lu1QWI
ByvBetpN//QNILi8ub17/Om6X/IGdxk/uzkG2wFv7/8zHA+3hOWo8iiFxWWzQR32
wBXYrrtN+zUSpEX8OoPWlPhrAlqv7YEVapWHcQNsqP6FCRWlsMlcl38TgFrG6qpp
hNdZ+ED5ohtdSCyTaAwgnoereLgAHYW6csZavtziE+LKSTVZAVX5BV/khLkDz2t2
yfZXkH9Dqv95rWpXZL35o3l14U8kPCmcOcF8775G7Ay5/LJBHP/6sjvydTX5iubr
EX4lGCPVwYNN1zOBfQQkod1nTnOfZPfmh0ivBwsfxL38sVvUjQsLxAcZGoYMkSg+
DoS3Dj9tCmnp3HqveuSyOiJF259oqqZoodzUTium4W6xjytpVcNB+yC4laNmaovB
2ZNu0YSCSjL2aoSDJLPPfPCiTvOUjSsSVWxZUOOApu5Hv3s+ZvfOaPwV4yIaEmLt
yXRtGbIPj3Nb63YTN9i8JYE7eAK/K0iT9QlE37CoYPe3ETJuxg3INig3C4qWDpMe
OBsOFsp0EtO4/0sni+0G9HsVqqwUahskXwsdz/v7pPYd7iZdt+PSUPkJv8lOKV9P
7Dz79uC+Xh0W2E3O1X/XcLe/Iz3seekGoW2gTICX/G7NVA00h2egwX009T/zPLvF
r/Ij9AkBYWVvH9WKXVvpwazgkNeqRP859VTjf+pe+mNgLdyy1lVXTfb/RgE7qe5P
746lOGWt3xedIlb8Q4zluDOEQM3X5o8oZWm4rPggCSUMAD4nM69ls8yhXVgp2uev
ccErHPyBUuEC5g24qaTSzdSYIRrnWe+XdA4Jsh5Zv30xt5yGjxOavz3r+Q0ux7/R
RG4qRedMqFzSlrIpePXiPtYNsZ7wHFxCCof8hYTgdGvPdD+TOt66RYeymf3j6us4
NFZ59cnG/NJ2NZsOZBlVaT67UYaCMNZG1G8Q74wLFA8FuqoRPVN+yl6+XKYwFYtx
eC58Ozivj4XQWHOKsh4YZ5vnrjlSuk1wMwmSgm4ZBlam+JQMJ+DDuk+N9HXLG4z+
PwdxkIX/oS0Oi53l87JRXNBiPU6ad2B8SkTlgYp4U4hhVB2B4iyfDLuI5002ekx5
EwAQzZigs1MMFMjjDQ0pkXevmmnnvgIaKbi2e9yuejoNBWog8mll+TqM2G+UKTTw
nN25rA6PxgNUGCVQ5cPh0tyWTPKYs7ttNz6FZnjmtH9yxjuRxKMOGNOs33m14nbS
sSSGPilBgxIoPLWPUBlwCzfCbpUCzRTxqzIEAtiyGlymJS/IvS5Ke8c7B1CmSVtC
9pemDG7LX2ZU3T5cm4IMSYj+iQRoz3Y0HPeyGNNWRLzNje8EopTKBm/30VH4WaPZ
3qhJvkzzz0rlfWSXMQXXwnPwBYXGI9ypEpx5gvHQOCyvj7g4cB9OhzJaYrVZLK9B
aMo9FVl2HidhJb9IGU6IWlxesMup+I1bW57g+GqiJRWm2Sfi2M3wcgZ5scPhObD6
EWKNKc3lV1/kqVtMMyZWOu4N/JcGDF0EyBWqajT/A+fqeh3c7vRa487iHUYydKTW
ptCtjYQY8FSILh8Ha4ykyVSlWBJyWOx2pqoz1kLn70sdWRlqI3q4UqFiJdJxFlj+
Lk3cshM0immd7MPXjVvpEeYnVcQn+OfhTBlpFm631ytJzqVYcpNFS6K2lqf2U4Wm
wYViZg5JnkwiQ5ryE2Whb56E7DBTHLFHUf4coCDRnjm/j5TZPo+bNIbGTGWEkUHI
fjYIk4Tw/AZQYF3qnELPs4zCgM5boK0+o4MhmA5az7ewmbD6cIAiO4JFjDWLNpl8
2JwqW6ddfM9369yYdddJO+F2BrFK1LZE8Jg6wu5HZX4dR5GxExg+ZwohezvAJCVo
PMhTt3avu6rXT23Ult2FFi+EUJM7BoZulL1uZSb2JN+fv1c8WT8Rp7H7T6QxZuK0
x5pjNb34j2GMXvcI5tcjCaK01cTU7krvvACiN6F1W8S5yX+Iif1p4uZ2Hmq0mLoS
E6N4E8c0cSkM9FpWt5z77Dki9iqzpmWmJaXmPw2gbmJcDmMYxlP9e2E2gJmFD6en
D7L5Gr0q01tBG5CcnB6wyZ3IjCkMejzmUCqGf4usXfwbU1PmvnLZK3LwEriKcelw
iOc4NYXTZojIBhswounB+ik5nU9kWm9RnUgrB2Qg/DG3c9+JJV5CaAhEBNVRtEpo
Y79+Wp2qjCQVjO0Dt2IFm/5iOKpWdy7VNW9lLXYyYr0re9MCKexgs7kIFWalXcka
OV+DVL4NH9W/tQoaB/ZtTmFSe4bFoALWRO0RjszUAcVAwxMdBswaWj10Yi/4WHje
9B3Y2lCFYJyKmQmpOVmedFmf4jd8tT7rSix7gHfKk1dHC/Oy+QDnjGHLmXAlwrFS
klaR+H/pNbotRLEpERJxpPZl0sOJXmnV2BrR34aWXA46g1/kS356GvNg3MCYLlWt
6StnUb5z0LoWJDEDbbijgDVFBkJqbj4MHxLtmqDqbbuj4FOjvD5482fvBVY9XL9M
YdFEgLWab/CGcvwnhRtobhJfjHzQ6lr5A8jkNs5n2HyNsTjD4uw5K3Vlb0r233oX
fa9xcczIhN74LcauEx+tHEJ93m2z62s8u73qRVa3ONdHCgPdQkh77sd7XoyWTmG2
1uCMo9jGLn1pSSq6f4obd7qCWl/SsxMAMhErt8I3NzgMBQOKLNambiK+O7x1KQ/C
Dv3rTzcGg1sSZCWgzdpPqEVMRnxKzN7nBxqni7afu5QyGJDJmy6TiD5qtVraXU7R
sbv5DBbiFEUGzpeIIq2Hwts0WTEuKk6IX2fk/B4RYYaLbFP1nNfG53Y5DaioqNrw
/Y3b3WPP5kZsZkbNgb/rGiWwkSQ5FHN17u6LS2L7iRyf1/bcKLS1CK0hP+2ImIH1
tPAzzmP72XahnfDSauwzmqfC/nMrS/bQKYA2n2V5ZxRc/AhF8FY3hcXJZb4GC574
5XMjg66RtVpFwd0s66NlTKRFiv73amFroWeaLlfQLSwTEEG6lDx2TdswtWPjtL8O
tIFehnsE8T/ckIbqtAOKsjTpdcnP6ufSEl/qZxsNygy1sZFfutbn8m1JCC0pqRqg
qOhjMj8JotCmRrGIW09MEMn7jlsEpdr4A1p5algvJ0h0KSLekD4b3P2vwdF7ieUT
ge/NG/nIq8ua8ryazeEgyGNwmScgqalk0i3U1LP1z2Q1GuaPLwRXNl8YlII1LOtP
V6amFL04DDxMztsi4bIIqesn5/akm6h+x/40CwdRaElYJVs3WTRYetffRoVTb7bI
HImwz1hPsrj2gRCGGAps2ElPFG1tPGzZl4b5Ttp2b6xpUuV7ON4FuLGPkAqExkEY
JdA4UKFx2bKpKt5H138z0FkocIDfXqSTPVKRc14eMN2DJnxjtclcHqIRRlQmRk8G
htOJSOQqmVguISV6GUv7jKGrYZOfsN3HpOjVHjj+vkiAZjNewISB36/LaHwsa/a2
SllpyXD+I8qHtHzLnPXE0x0XsxF1FI/IQY1zb1x291o22zroObWxGWidI34+aZbm
1JRKR75TMvs0P1ob0r9+2KxyDXv3fAsvUPLReDEXeLf2LiXG/ostGplZDrcRXdYJ
tORWBzcT8QN5gdsvMNGdC69fLPEAtN0aEDaGaiZ1wvu3xBj9eUYgF0tii4PetaWJ
LiuNZpbbcHiAo/5+hqy+6jHnTxKgaR/tJ+xQ0ie6vB/Kc3WHbW9BNcsfsmXKHBbm
kUsJCZ4gYWZHEA6N4UhYEVMFZVa3Fw2TDobll9vvFKW7gAaDMafjayYgUyT8wyac
Nm3vAM64CPDk2uBEkLQ95owv2x28JChkCJ+uTp+O4yFf99YCNOIXemIzxBLlHcjD
VQ73bVsOoraO9qFvvm1q5idw/2MDyKUHXUhmJvIcs5Mzt1oXeFLySPL7w4GxcJv8
E/Fhjczn7Ix5SipN4LTOvH/ZefC1Lc9Dda11/f5mY2PFUXj3/KWQdLwKExaNBKMK
5zvA9Gj12oIXV3zkLerx9ljep6y2+n6xx8OzpiUWzZafx88RpsipI3aXFYHFg61a
3S0/kXCI5eClWEE1p88j9H2pGb8bPO7YSZrxSfHwx6IzgzCoyV1wKe3j1HnO/NIb
jZYmNb/zQm8tRqbjJBpe3cN3yfdgfKa3s0V2bVBgpTVSD+vZ1GaDpvuQ8ARcoQx0
vItJxG2s9Ye3TUYVKVCfb8pBQSET2zLYWPX0gUbxCvuAcORdLja6nFx/JPtfTQTn
0CcXx+S56iLMI/5odWKFtou32me3NPFXBd5jq6Kz5osCVpl8t8hUSsgC9hZgoiQd
B+bMnJrwmF9N/sQeMIL0ZsM/2LriqacLcP+NIgP43bjPSS/YVdqVwNfm/LKhJZBA
gIojMoKo6RE2qCeAMAD9xFDxJ8MB5GYy53Bux/et+GVC9WXM6yI6tXTq5F4/ElQK
S33yfQScEpNgsoq5h1z7Ytg+TGlW3091QDhjjYeUCw16uwxWLtdUeAXRuOkZIsIE
7AuEQ5LUeaHaDu9YktpAEGtLHXGxjP5Bq4glRT9QMx+fqI5ZnrvNil1NKVwLR/jx
v5nJQBnQj1QX1ExYDowwgKRF83bNDTGs1PK60Luouo5REGZwuVxxq+slJLRHAw3P
T1roM9nOeTUNSIxKmV2YAluXvySHVyC9rcGwzwO/qDAG8/zaKZeDuU1UhbmNrIGx
whr7TiLzGlOgbTDu1a2C4TlYd5cwmWaPfvzQgo3oWPM8Mja7t6F0VYqMfGwmgTFD
s+l/fcavDttkyEgnpMHKgp8XeugaVOAXsYI5hZG/Su15Ah4ETDXtqCyZwoUDJV5/
YbX+S30AzGBlcTaGdwxWUX5Vwd0Ce1rqBC4Zru7tNx3thg50ecAmfnhA9yWYEt93
NelxB1MY6KC14k/vg/wnJwkVkJzFbXucH/utb/aoup1PrDRYoYAuJELHh3Q7Nq1y
bcYNbvClXH0m7RDrcPSS3l7/0iDZ/X2jxdr2muUIcG9V05qZvmgNDu5ii82CLMgb
Ln/tlNKGCkGQ756DCy8EbXbjkIwCuOzdI3cth7e/KRpjd/mW3hpGUJIM3+yIdlBi
2c6DMaCGUCJppEoXyIVegt7p7Vv0ce9hInv+3SBzf51019Pl0UrnnmHO08B116JL
mt0s0cbV+gUGFq0FH79GjgVDuN02QHL/ylpTnwfRDL8dO74cjKX87PChEam1KdiA
+3lWs46ejSyaQPGPK70eOR+X694IqBd80VvmBylFWNHoDnhcG2YCmazTIgzn/j3C
CS6Uf05LRBARB6GVtt3EhD9AXBh7zWca8ivsSfmrGa8S8Ax6Pr8UP2utKUpXmCBA
0es8dEjU/537s165OgQrbhIYKiX5FwjeBGSD+OQamR3JaqzYq1+76rTPmuDD2okC
FO+kMmFQ3QoJurjW4j94P0dlLAriadEjObXvYsvIxdTXAOOZlpZMgEKshIlw5xzT
hOOheA6H8LCBJwRFVrRVRF0URcn5wPwDn1hc29Wxrf/R5rUr6Sp/QKrKbe5FXLWy
a9TvMK/IIeG1yFeRLu36nZQKCEC5IxT/+IqNxmoIOQXm6BuFeqyiMI9g1YQfKKUp
GGHb1UJJ2UPjrZrHQpzZBSifwZ/sNvmIa4UoomqyybLmpBNSh620zWg0IOo7Zt/G
cuaCHF8usDn+8KBmXBnJakUC0s5Ei/c66RGCcbdUt6DTL6DCfo6Q79KWR2FpahBx
o/fqrCJHId9rG8CXM1q55rvRp3+QSkIzT+mnhL8spABJXFNQYiH5vvftyqf5Nqob
uNfBXcypwvxTKYaO2q9QCgkJsZD9dJ4mm3+5969G3XmxJkKlM7z6r1ef6HLn/b1b
0EU4PCyRDOLxmZMmzhq3QemSGaDMDf58Onf6RWOjcXUWHFTh3EQdMBhCSzkr1OpQ
oDq7yWN+H5W++S6z2wDcpPh/OlbmpBCmtoqnm62farKGSqGO76KSlVUMz2Q3eAk9
2Oo+c9WSdUMMlfWUvBezAos+dFr5LpzH1R90CFiu1K0DVAJaDjkmBdbDgKlEfhFB
kAw1na/rmgXNU0VJwxmSm03pW4zbU7B3vv6+Mlqe0UKgQJ4KRefwPCxc66I4XSXY
8kMk93j7V4kocH9x20U59MuIqX2VzPdpDpIuHrUieh1jwkTyxY2sEe5iWXwmlItj
BeQP+kZgaK/MCNiXJgX+e8DbXHuzns4b8rNUMUyCbUxpcHki726qKTh3sV3nxghy
a7ClCGEPq+KmHv6LER9otz80Ssny79O3SnlalKN2Ebr+NmfdTi3GlawlBdGKF3pl
rGczyvg/k5dNylfdd6ZSuhXkdnDlc4u519hiXud2qqe0hqi+ut5dGSYt+TywqGIj
GzM2G0Tpzc8NpYp/9whmxXveeDZQtmmNFPG/N1XhRaRvhP3+o/ViuWQdM8B96iP9
zlY5O5FlsBh2loo+10uMF5y/CCRBTUKxl+d+og+Z4z7Q7UJc/0CFOZKm7ieBw+br
LwuKVhkuBdm5ySScmJ6fBHnm+MLfOT2bMSc0Pz9GnAYlNe0z323Ov7oTj+/AXmvq
lGK9Axiw8ku/TDzH8XL7+vxoI/l2n+CDwJeIiTh14sO+hSBZdLPhdUlfiN00diy5
y4d1DW9fBwKI8XKhJqwN38gjsBOKtdT0E+j1oRq/TB3c16ZdIrUvvCof8bQBdCra
LWgApHW16enrAUDS4epL+nAMByA/jkXqP/394nlkC3V5IGQ2qbCbcUwm1b40YoiZ
KiK208bz5TPnOB/TQ3wMuRmEmAthmQO2liCkos75h2O/B7njzM356Fq/bE1rLwIM
nG8IJ8bAfRBZ9ohuf0SRbSBef9RPgfYt8lLx05n3/NJhOhgcXau2YH2yu39tfT4C
e/LBSLEb/KG0JC8Lh1/BNrCK3q1D5JBMF/W318fE45aOkzyPTeinzcPZgbb9LDbg
9Kcy4iKR0Day4HhG0CKOT+1urOWOY2rClaeCgk7RGpMiAjqJhw+ysGF4O4P7tGiz
Hh21ytRojlvvh1lxZl8qlRvzBazeebb2ZBPgSMg8S5BDePJgHBK6HBF1+B0X9JaH
nc7L8kONh8wu5RLM4cuUtZI5xzwUwit+gt0OW1Eo9RjBJnSgUShy72m4+wxO3kH5
NukrN2mOmRybvcx0pgG1nFTszzqEUabtmSndV8gu2Vr9UAz+0L+cEdysk9BIvOcV
ihYYHOEHwrh49N6OKxsJG1JkpnKR4L9wiBdWvS1ZXKVC+go8gjsQmHxuxVMzzkU9
dZcao4O7okjaqB8S7Qyli1DBFIxUSxJ3jxV25gyn59VXNCbex4iIdEeoM7MZ710Y
E0yjp8wdam+zfy7rCHyo0eGt2ZakeeggXaWu+y7N2FqFZPPxZxjjyPlJE70sRwGX
yFOoKclaGNOxmw28Xz2N96bg6u+jVadr6JG7LqN6Geh0e/pTVzz1gRvCtEsreSFb
XoVKa2EHOBfKCDvHZ1wGVpQc0O3SVKJFChLULsj52MdmJV92MJhahMZXKFLziwZY
zaU7/phggoig0bp8h/dopp9kTiY9ObvW8isC+HA1X2V8JzJ/E+CIA4Jp9zgCNlsF
WHdAJ3Ss+YuLArDycP3cjuAAsk7dF6O6OtYNGMPe55ofkaLdbIlZ0x6ECyr0AcpD
NG6BVU7cYEZW+fvXmJ7dncwFkWvzsSPUgV3NkXRhC4iWiMMlFThT1jy2XFHbBbKS
wV6kUnBbbfEiWoHNdctgsKkdXrNHO1PdhrFlsI/EKnv6TSdRJcjuztMPssyQLadh
hzTIv9oh9R12UOgjQWL/p07Gj6yjj0axjZpu3HJ/V3AE2Ih1ezTFBot22YtWnAtn
1sjwv4ffVY5EtKZ2RHoI7lH7jP3cIH4zwn050lxOAyelEJ0/AOQDx4gBNXlGFhj3
dToyqBNEWlS/M2kf3SUYowaJ5WkIusI3wVLGgxzyM2iw0ym7oFc8YrnLpXab3Qk7
HudEYfQEr/ux1ID03Cf9C/jI6H1+PwX97DlGxcmAwwXQgg/9Www6QA00R7IXWFgG
P4PiAhCvqiPzhD5jadhiRtnM4pIC64gEqKcaJ8yAFLO4e7WJutgow60v05x8kt4K
sR2BU04wHeBHaTowKeHx5do6jdol6+whp9M5fL2e4WuMAKr4EZut7xcclPZS43cP
feY+9aMR4ZIlBngUFfWGKwm8aoxHbR13lHLjFSrI16poGVfKvwbPdFDXq56Fl2iS
h2zNukyxcMfZdH+3fzxrlkvG1KzcHMNbw6TT+Vm8y7GVmkHh53TdrM2HyMI7H7xZ
fKZlU8nkq7Atda307V5xctwjAwg0oLfEw5r674cSuUv7QHqbEkZexQnEocYGAMyb
L5xfBytIO8HCriy3vM+Cule2l3mGGoqGN1xKngjQzBej+P5YZL/PqpMNa86M/Nx5
JQlA/dTjAyKBXR/uCIb0gz1OwqEHwE5GVwYpxuzXbomVNkvJiqdT5B24/bHdeVjF
0XkIoOcWcuZbT1gqUMFI2D6gdKqQpzB+kxvHR63CxJDiA+7FMLAXXXMaNoPQDzwc
Z1M8s+jl0M6jHxaAjqPF7j8wF+2x2F+hpFDXaIm3k91dc7mu19k4H3tEQVeKecug
HspUvZIeqOG3sOKjxvLVbns9ZeQX8fEN5mHh6nfXH96kocv9PVHxTpj1cBET6pOR
vjYFf0uQ8rDjTtkx8npNsgKfXD+ObQTe1kzFliTyopRyoI5qz9zGJ9gs0OlJke9f
5zQno9wzbQaTn1ZmEb5GmcK2aXX3FXhG7Ztx5if46lA2cnrHlge3upAXwvHUlclC
9dyw8q3nV3YZMcuzteQokAWb4HPCoAeho69q9jy88MT4ZVcOhBOedlV7TRFI44p4
MsDMKiwe+bMYMkYbCDiwalvd+yHR2i/sQVvSUVLGrfynmu8P8xBm9WxR1eDgyh3L
CSIpr6AK9CxHEvRIa30Odcjf6gXWwM+Kdkvjm0y6CzgQ7czVdSZgXgN5uHXUHRbe
m7yDW1s9S3YYJTGgKjJ0/cy8ElJUC7desMWqpSD3/o/P8pjVBtgMFROYgHsP9Zag
WBOhR6tlyPlOE+T/KsTgpAn+ZJEUsXaq9iARZArERECilh6UBeNiy9cz5Dn5iIYT
KxLjbSoEaFeozExC8si1vpDyEZia/84q8ZSkSdwYix8ybmI+Sz6YxGL6jV41/X6b
ke6aQEGRMBn1HbEg7ijmuXQKuoynZ/Wrz57t1bLErpHjewABEkwiJbYkMimhnIRv
/rJGWD9OJnWcn2bH7ZobM1NoKmBzHkkfrYmxhwnPFKalbrbSwDYRiuqRWqHfBeSC
SAr/b4CTG4rAvECTsWS82750osqyuyIj1vq8MO95/tQhBd478M8AWkSaQBuQWj/s
m3T7tiRSjypH/yhzJq6DFOGJ7YFMnRK3sWnOorXJ6z4S1NvtDwzfHL4oCigSqrNH
K0xryEMrsqTI5suLWXAAruA7zPlSVVF6SMFX6RIZRYLOySmQ8+dQnVyG4IC2oGC0
wq/iBHc4kEZ3p7yHlGblrjjV5bSqW+Sw5mDuDsfHF64aYbBPjUDsi7VcjnE73wqF
xAj30EiqFuwxjNU4pZyLpim6Aof0GK9A5NKi95JHe9xe5V1K3PiavdDco/i+QPak
EAZmw7LH87MO2+eCVG0/RnNY56E9IqGj5o+4LqoR2oWP8+OfPjK1E0FY2bcqZ4j7
8U8jjGaRsxR2eYAFUgiOHLpxvm2S60xqMvg2gHW8/bSzza+3l8Y/hbULmRYSbpCo
yVx3fvtQvhiYHhSJeSIL6q1W+2/WDMcVEVmIT0yG0FFBtgxnPLmtf+CrD1jGdR6m
qxrOeX6JpwDnycD4wdj7G/lyFnFrAWDmPHz/6LARn66CVTBZFSNYeDGl8hCxBCZB
sX1wHLOcSeIvZXazuv/RAhlfIWP9sw3j9rX3sJ6Hm4OQC8Y2Eo3RSwI6RIYOO1Zn
xK+R6We34by90SrR3F9hG478f1K2H+bhAiLWZJ/mDVWXLM/AGqlWp4dTfp6woi53
cJ7tD6O7baFFoZIqstRN+YcIsPxvKvQBwEArRyDMK1LAzm6G3uKvNn4Y/VJpfFF1
+Os5f65BqJ25PmF40sJs5UaEeqL2N3U6rPKKFmrEdLlgcN6vHPqDalCVmyJSFdT7
D4eNt1/F6gFyKBlazpiG50eaXKyzwODUz6x73ZRYpHKpC6PYt3T7JfmuSK/BJPma
EKP30Y2N2xP13vXyWWo4pSJ367E2ecWdkOsDcZmsrFoWhi3+6pfOfA74E8I+psTG
Nqqy9yWBK1ZtOuliXjIEpjM+3CowdoryzXtQfReBJnXwhUvRoN036rckmHQFuU3k
8z+hWztCMVm1jJTDqnsCzfODcxqdHsqqUowsXNtkOinBFNp1tY8tEj/aHIRcEZCU
WYDvFE0FSK+qnVLiNaoiHYku8ao9PnmUXTLbbgX/H0XIg0E2EoC6EtnDU60Es+iT
k3lv3iX9rLdkpYd6i2Kpc/Nn87BofrnKIAYtwQCY8ioHLXXFZ1OpafxckRRpwFKi
JlGaFycbHZWV2ur2gi3sfOGZggv0hnzfwvWmgT7tOGnkdKHTPbZ0bCIyOyuguHYO
QQGP9e2S3VhnuXIYZwXLoSZS5Oag30uyyJ9HqtiC1EcRqFtxzoWd2C5NChI1GvW5
VloRz78ixIXEnlW7nQuPOJ4FITI1NlC3ATx3YDoNfe4ybE6BASPXUmIqKDDXfEyF
jccsooislCEDaw3NfEvx3H1wXzdriSWfHE0P4pUb8ho5SbsAu1AAK36nQ1xkBG7A
W9eCUKt69Je9S8bgMTyFTMfvAZ+T63P/7OFdcuuJimc4dNTIEa8pIKaWqok/rO0/
ZR3sJTNFpaJ8GGmDgRAqE/FHUUtOpjtb7nZnDp6eSh49zb8IP2qSquPwjXyVDz+k
Lkxq+hVWluxlUqj7EsfZ89T3hTe3x/LUPbDRq1EDtKW/yt/lpLehQ1F6WrHV/RBr
C0C5qkBNgbR2jTHmdGpha76auElCQha9pf5fsOAhFpqXBEw1BtNFp/AmPfPIkip+
QnAEioUf2CkiDKM4AW1sxF5BO7yayxTkLB/zEzGfSW4jiC0HNr/vzvN3++cGcSUu
090VBq2DR7E8IOHXyEk5k3XOdMIou6coYxLhuguOPKjP+by0A+SUO+wZZq3h6tyi
XuNFpnqZ9CB50YdSCxnzU1Drzoh9/tIFHP4i5yBuf1x7GQiI8ioDPd/6UTAtR4jq
LMveaZBXgQj0S5W6E5tIoTTaF73viIjP6hj7RjGJOz/VMeworSOkP1+ZeyZGeFVj
vxUV8ZSRy3PJCSCdHhmyrK52juYrkYMYrA849V05EYcyRLthtAeOPprMvi1lq8bt
adlj4ErF7EvE8REAcHk+qMUXJoRyY75UtldTgl30IXFyR+TJN0wDgYgheap42IZP
nBbDRGzOhuguZsbi6tgox83pc8nJa7u9CdFBDrtm1k/l0DxDKbJGeexuk+jRMk3R
D/jvfVFQJk/gZHcRS1TxmpTrKhQhAswrYMG9f7sGxA1NBwcAx44p4eFf6PI2OAbv
4sQNezkfADiqfDsUZ65WZREt3JWE0Z/NHaz33mRubqsXk7+X56BW973crREU6ZeI
DE7KTv8GwhZwTFVEuGlLpg2RLIZbJsQ3CZqKc3PokMVR9K0mF/KAp2jdaA6xy13p
5MHp9IZ1BjxuF58UhAsKCjzF7Z95a1JiExA1eEH57Di+36LJXIYT+NhlAFhLq7E0
1kZHn4nQZAMqW8r7RUDHIt4en3ZpH/q8fy9ggMFL5Z8nisTFqp2pA89AOEIVhRAA
A/h/DCIEVOo+Jv4tf9+3/8Rcff9eqzbC7dJ9NHnb+Z48/Ud4yFE7tQWLAQubFSvO
T/Zx6i6Dgz/iExCTg19gaR85fpcRMNttbYkGJ/cJA6pvKn5l0u/HWapiIFSAoxOH
L/9DBLsXYS49dTIANE7mAr4PnvfLpBVCUdOeb5ji9nHLNwcV5o/d3p7PRCYGsRem
E9NVp9tUGQvhnt37ObfBeaoSqrmosmDiNh/O/Ee1iUiHdpjk+sNuwFXZVltI43jV
TqY58CeG/LcMxIAMbmK+cZux275IC1Ljh7bhcpvFLM+6k0uZFUbKASy0HqW8YcFh
MOzSyGieJGA6oRZK2sUh5LX28lGGrpdTtttsvcGVApBEiB+2XLBmqPRtnQdA7NsY
JSCcRpxDmF28EnO3aI/1hWiXJCuC35oc6qVTUvAkv9ZzM83ZzBY1V/XUCOZioh/D
J47duL8W8jsD2wOSpZK6JPbnP6STT2VLcxrFf3lRL5OGLZpE0OrA71rVF5r9pSRq
AueD6438sY105KHsr1fLFaT8D53tuAJgoq2Jqq6HyOLJQpnnyB74TNqjrDw2xKkZ
MzJzzmCnLXJQHMhTajEl2AvJGW9reypqDlhlbTx0K5A8xSkJYeSi/9z1SJMFIH79
7nJD88o57bO/i/pcK1MsfZZneCJdTU8HyKBSkgR5W8BfjUvXt7eDM4kD4pIK8wJs
QnPFmbSF0JdhXeOMYbS2pTS6Yn05GpzrTsZu3iOXCuBu5Lt2Lg/gTNO/ejm8m9bp
dxKYVIeSuJH/DWsOjbanWu4OhDTiJ8crpeAOd81F7uh1g7FKh6e2hy34WDLYVfay
99lBErF37+RXR4QWT3h4FbaPt23ZtPRK/6lVoB8lV8+DlDgwbAsWq+5NA7ULQnSg
AGYMR7RCuiog3lg3Bf5AeNPj0Cruaa8xLekgQNTTmEptYZVCKeEBvMvBjtAn2+WS
4Qp15PYFObpbfDAcUpZIxbFTEDfam10nHM8oBwB46iGubQB4fBb/uj3bd5mw37uj
4gLyIuu1QnNJmHa9sUXOmEcbvAoR+yKhMn8N7OLBErbxivtcQP2/BZI9hI+v4qBE
Lzp9sEV7w6yGqQANO2BCGIq9Ceq9xtiDOsD/B2z0XmcAFRH6yYYykWzJfqLG84St
BwWck1smapW3jf6VmKC2DMWvhUl67XMZsUGCoVQEGJxBsZVE/EH6xwMupC8fwn7y
+UOTJOzSCthZt6G+GdAeaNH+KzvO7P/CAxTg7WR3itWOqmGk45hRN6a5kJ0cBJha
wlVF8De1AvHadc+uUwF1IyQ8dlCQytbvuu9q6fAsBJ2VunChrTq1AgqsFd96nlyj
ELPvNiAAxYt5V6SiY9v19Wl9jbQ30qqZoKuZy+LQNDzhzQ0yiQnCF1aThD7a5dEs
3ELtLK69ifXEno2LDT/5MiuOcKscs4JgTb/Cff4JMqY5gwDf8LgFXmkMjv5DGlrJ
Smx7GmC41z+f8ILyOm1obeCbRurxyq+t8SAYccsI4B5UQtItPxr/M0bb4M//8Nne
JGdY9Jx5p/BKCFWKz0d1zTfbniRXUrXGGhI7iNHD/y1dD9/j+5zSMg2kGBjW/0lI
TSqFUsWADUrEeiIyJ/sJ5CotvxNwWEjSf0yP2w6pX7ugNPsSELUxHdSY/tTSvxyi
9z+IsR+pjhvWVpqgW7nRvfpriFGLFFRDd0hrGEypjW8Uq8daJJOMZVtTJn0AxFg7
aLFE+LwR+wkrqZUpyDHstGODOuTOzQshSYVfd9NXUs00hjJUKA+iauXcSwLPlb/u
3FVBJO9EpMyJwrsZ/XT7IbAMPOzGAcVrEropLJ+JHJMxiew3bjYI6FXbaD8nxHsx
bdR9etQtkOuT5zWRBC6ADC8845bSjoNunptpYzM8DvFKDf9IMCFYGejW5/N8J3cF
xKNTkmgWq0jK00kr0OhUDLcJ69snhhYoG2aI/KQ/NMGJy/uP8ptZInqwnsRKg2VW
ZDXQrS4000tF+iUkhM3RVYh5WLzxXsavnuusXPUIMLHIp101WMIQFon4A1dpanIo
Bq3tRcQ66xiDGZFQepAfiQvrpzpqiGisoAAX9h5RrTZqlZE0hLMLU79nKPFic13f
Pz5wa4aLlQeo6fwfSAoegwpAJ8LOmtQ0BAiU7kgNNJw8CSsd7WkikmBUOpwPYqAA
28VIfqgynvZQULCyoGSBlIHxd2ULF6mffAPfaa8rITifMMKXNtoJJmrd8lXpe5MD
eTSKz1PAC0w0hD46QjGud+GrDzGvUpZAMKG5W2LTFcENEARJoo15VhfD+zb1MZJQ
IyMhzZd9ikMqiHLIkdYKa6zOAUiwnEHILhhLOB9EW7j7K2Juu6VktaBwolkbxZ93
HEMUaD2rii/18SEIqab1yjnnSu1KOR4TscM3wObeR9zjynHXLtKk7nU8f8es5ujw
Vwp3LWFIHAJumPp6dZPqPuHZ1yK3in/WSJptN/7Hpx3qxZ5H0deysLpyTGcOQU3m
NcjYZ9oITTrWA/mc70M9sidvdAADepoeBtwp1yeOhmlWPJqjcbv0t29pW42Jz1Ja
1mVMzQjRT1fuUObgQj3lHj4nWLlf2VWtTS4MFVZiGNv5dB7D8RH4hfbPUjzB3C5y
lUQK7NISLQ5bfQXYtHlNi18DIvGYdcVb1iY6jZswIr3Mksf0wXtVs4og5d4seTuz
AVetQarBmVAQ3kHPndXxI7yudIwbvt+WuOQc9pwJn6kHmbGfOLxqz0uV3collo+e
StLUrbIsqMondSd1AfAcyhrSIkThmcBwYYejcaEZWGnL1iDpnNRQSV+p9dF9ktGH
2jDudC8y3SG1ayGU7mFeT9DFhGtqvbRzwqIOUbz/XigT/FEmdw2W4zLNtvQMqap1
lOJf6zrcnFJPcuFL5N8zu2niDxYoESQKPCQ8kaGQDRbSaLBtUMLb9zdgXC3GCOiw
F15k38k9a9C1ZDkzW2vG0vdfJJXiXbUREBes1+q5gniZ3rrz7f6Ua4hudBuRiYOq
DhjpPwnJox3Li3gSiQfL5R0sLZGmKycmj/KgcLWGNS4YUiX2nnWEzn8CmBEVyDVc
bEMa4kzSchjUj5oZ+VSpBWfheqtDWz19XHaa+x22DHs6E7rL6OL4ZQShLEb0Q7NQ
tkuCA3jthoswyYx5tHdLyWuDdF0RuaMklbStXlleJ5JLs0ScOMnqgywGEuUZyR3h
LzR8zss/8dEjNo2U6Cg4YMO6b4BCwq7dksSkLGguk6ltFSX07LYmIRWygtZA+vI8
wkV9Uzf1uRkyzOqbjq4HOgGhJslqVMsJbcwg/3v4+pDTRnRDBIvgY3Jfbq5ZrsmU
xq2c/KvA2QbZM7cIrj6AgsgESu5AWCg9vKxtMW3RM6IQE9rnXDXYwpS8NRZh7KZy
knOo9eUdi3PPFcxt50JL2rQsg9m/DGP9uXTKf+c96gsD7W9AWRrpvg8RQIJXDRGz
vekkZhvHc6IEL3Fx43ofn5YzvI8nNVc3Ktf3zHDvMsF3Xbqds/2D6aBBlD5wNUPI
Q2eygoHrP3KxSEHaEcFb5owZkxNJhr6/ew/9oJXMOsyqh8jzJRZcIuMJx0m6L+z6
gDvosA75c2EgInBhNv44Eb5iVPWHS76YEcFUxFijni2GDHMPPHFIOouBCazc/beN
/i/PJFkxxuksDlRgAK4MH7W3JuJ/67aWL49cVR7CMbYcyAv48eqac48sHkMxhyjD
eHcNCGOvCReEe9DE+EHWt6ob7+LkGLUtckekRd/E44VFP1vvkazMSI4ZYkGe6CwB
AUmbFSSLUdFMJh6V+EjGb6bUOwotLW5XmXhzqDgt+weYdAnvbmKKbXu1GQD5aoXl
woGMsInWfSlWqvrWohEcSF5jgeHMlevXXHo5I3SnUpx84dJX11PZDu71/AyBfbga
k2sjmKXMWmVQ5ooi2YP9w6oGUBaBALW9062T4fie6fVx0PZ6XwvUhWBj6BFneoUi
drrJ6TNDOFjH/n09CWa0pvCtrCn8Rxrk6fmzflVqnnosMUnxaHFZkl0+Qw7fd2Vm
6/JptxEeOYlkX3eOKVRnEvfpgVwAiXdXHXacjxzj/fMQCObCaH5t3g3YKIyobFCT
wCmeupmzA9yh3C3UHPAHlkeUUoS6tdOHHSFXwCGl2NZwTdKt6A3hOGItQbSSk7QO
6hTZNqRsLwziIXRVaxVdUbR/SxD4iFqTlQAjZJFW9CQoJT72n1IOYyLKR20K4rgA
Ra2ybFko3kJ58ziKZTIHqWKZVUwRWW4RLSx2GHFd1KxVEe1+xYKSYRlGCG23tPmW
yKwCRMa8NJf4pAQJ1/Rz899F5ZMBulvK9X976YpbeyVePfWHrICqCLyFBJ62Km7f
atc6t8h6UHNnYchd42B9lmshZ31kADIZwXdHbtJltcj2PhUligoJUBwsF6EWsUJy
JcAmt+kJ3vQFvS+5QaVOVBuK7utyX9/EPgTFXu1mbF/X1WeAtNghH1pzeP0Xi6LJ
InoAsPF8Bg8bSq+PV5CADes+K0LjKButIIcSAPz74FuC8/2yykcEdhr9oN61Ei3v
AwiQCVHxxPDJAMInT9NR8xoO61MxOhvdn6ZmeGQSn0DrjVEhB0+eSMCG7N/1gV7t
LVKVT57b2dOdOT9Ozv8HAqPlvtZGvVw7J4ZE5gUfoJu/kthzUQpDLrbwpobZHSMA
AGG2h87NfMLYzsd63BWn4AT7DHwXO7HHoRhD7Gzr7DruaX3MV0o2LHhKj/vKXbXo
GHi5VVg8OIUGGP1uGdT5RkFyLDH7DWRpSLW7CjePRvlhGNSx8AeZms9OALFf9Ppp
eg6dRDx0hg6JeG11UwqZ/rSRLHI2yzFuiY0AEl4TYYGhxajTtAvEw7e8MJaFyAMD
wVKULTxunMhwiepstIr0m7olGSTZHNcHdQo/dlxHBGe32WwomePSv1NF/XntA/wa
ghYH2otHg/oUBQIYfLWQIa90SuJrSW7YzVI3PHdOOFdeWKVg5TEGLNsViRZm7V20
W7PjX+Xs1w3N8XGKM6mq/1/kYE4TZPEkTIOPOq96g8V3q2xVypDRqIW8J8HDgRbb
Vvg5Wxp2xPPPlmjuo+frSNe5w+UL3YQHN4eDpGKpf4UrAfxfWtZC1NbyqKijKEcC
u9iMNqCS4T5yewxAuR47wolyixm62fLN8Agtvrblc95qLiwVj3QLFsyJB7eGKJbr
45MsZOOQ72yQzbe7sREcEXtyU3gJtOcSawlqUrhEGgCk6YzWQEDvWIgwBcNdyrzx
cGArJ5anyTTtlZoNo8u7uGO13LFl2pxrIWrori9WV7R2i3si5fddi31RPtSm8ec1
th2Cf3zmWJAKoWqK4Dy8ZKzTebmXABJrL454wIisMiKuNtkvlPqD+vJYqUgXKaix
hf0oW3u1eTWvxZg61HPhFUu+fenRt3LNmC7BJ3XZw4kOI8h5yPZTFj2GnyfAO6EF
ahuGdpSFcw/lzo2dJgChoMCgLHOJkS3MRvaFIw/qt/z/+YZhMoaLC5D/uWB3y+tC
7BZOsma+OY6ayvnpXpiPxWUFvyvVYVMnguxqIQX6oif8JExnQwgnJWIPF4xQgr9X
slBS204L0rAAWYc5EEICDUQedftDCQPxUk0cWN/Q7ufYTI3LPtpZRI6PO58oBGmz
ROIcYkpp/bodKVQnvsDF4If/tZxJJVjBU1FSOcftmHCgY7VNLGjegyQO7S+L/VCV
+AIRxFncKXx4PH9xBiYbZaNnA507MyC1Cp8C5B+NQKLSmVkBOxNaHJAWOwW/yhLm
vD6u+a5H2+WDG2TMF+Ut5VPhTRZWHb3YNIY4ZCKOQ6az55F/FURMaiwkfVlcxeGl
TcoFwiYo56M1Oo/+v3PwXKDxSJF0pCB8c7bLYV4l5MqCi60jGFvXs2rTuYpOOpOk
d83GuCyKlKqmJarZqEGUTpZTHXEaZfNkqgVcufXZZoc0XJMliGRkqk7wwPd+WYEj
cgNWJkvhwT4fkwjQqFk32qGkIiK6xd1gWdPgewrPcCoiB7GiLNsZXYZizxQ7EmX9
oTzYozv8so3YdbsGOzu/HmX9lOCEuEJdVvTsw6+Tyk4EuWoLgV+GpHIVfiKBn9QR
npOr7rpTiVcoeujDXpw6smFMaGFV7xnMti94D4Gr+F7vyZleFKV4d5AcVm00h0GW
m2GDrjUaKiHRQxgAkRUBqUNP7nzVVV3pfBl5b527RYOONDDNYyIBQxTEWVqTtUAY
tonNvXUnqohzK/73fhSScUlCCk0lhtdrH3nKO4zPBp/aNzep0tno/0rdJS0E3w4X
fQaeMjw94UwMQ1dDZmeNpq6p3KF/Rm8d7sqgL6UFyLKYEa/lcoSVgopa3QF0Rjm8
DhLeMbEpool+V8AQG5hNjcn2zXvi/hnnssHWLvJK0lPVibs5rbl+SizB/2hRe2ao
UmN2t56xqzAsU1WDt7CasXXVblK4b6vBCMo/GocdilCJTErJiXpQBZADGGFu5bSN
LLYU6oFii71ujb3YJBf5red/108wZq1eRXBlIYicT3FjnaSMraBbqvSGDlINFtJT
ZsyfKqIRfocTOliMQ/8dzchcQEDOtTC+/yCKZa8hZ8U3+byjK7hN/y11IKKzezqz
eQBHAkuz8Zgla49yGfr50AbsItWo/H0CUov3eTZkM99eKPodZ1JwL4NcmbUc4lOF
wgaTmEJXLYaVlmiCPqMAddZ7RgcBxLe+Sfv2ntVUovEdyLGHpqQkPQPH9TWn5+z8
ZlFM2XqZYzAOHEVibK0Smhmj1eOR5I8EE7pGxjP58Hp9QBAlJ4xxEUjYkAUIolrX
U/dGNmlJVPeZoSsrFZK2nooanJVNaCSNFwDxJAd2jRfWL16YlPg+bUsGHrT4wrvC
sHrhWh7blwIjlniVb6q9mKlD64w2LxFAsgnK5ooPXo8f5sxiq9JfSbT4T5pkIqkN
IgjlnIaj5dTBdLRyD8gKbxCsjntZBuOjLxJ4x0Px41nJMhdAD1fwttdUg7tIvB6/
07hdh6tB4huj1G1wu1KMkYrXV/0nOLFRENghdr5ZIYo2ju5p90mS/5pcp5Vc2yTy
39RPMYG6LRcsOBOSVBSXSZhNQd3JBsB3DIi5WEA46IuU/glriTNg6V30YF7XC9EL
AWjn9HapsosfSm08ZqPkiBzBdPMP9v0SbHcbal0/F+0u3K2bweY6D1Yv2xVmV5eo
0+cvZuKAa4anq15/3w/vYNWexKfUHu79ntwsl9wElYe7iHBoEnJIfZSFILNbyAGZ
o461Fg+ZNrn2WggJzEkaJvzToh60jqyANgakpvRGSC9CJDLn3oADE7G5cIcfiqLv
cri43Yg2txFKeP0d3v/Iyh/5b1ZsXMVCMC4D1YfsC/zBNT6eWTtrxKr6+m/xDETb
+DKwA0FEfuVi6cug7pxvj0N6f3Vde016zuoeA3E06DilsIrKqY0o0VaNdvKRBC2o
vXxn+FUQoqKf0AnuKf1KEZBg5+vC1x/V32JlKA3N4dJy8pAfmdFUsEiS0H5nxz+k
NlpoJgHb0XyhY1rayGHvonKGAJufwC8Sv1P9Yv0gZZmzBB77MmmroJGQIloBRFQK
V7xsr+qKAt7NXDkldD0mCt1uaKqDEA9sTMhP8dXTWCVsDauVDHwoeTuY2c2n8U0V
/45kVmO0PuoDVeuzBLG0sVURO4D6Sx5ytoi9Fn7wyUjFHgZB91yPIxseOpoAJesA
Fnq4RAT3fE54XZGtuN/4yfURuXnWuuJ4HXHyAzh5CcViHa3+7ChY1XHG0HlIpeuG
ZPXAaDaYw2j3+H0SXX3ab6wMOvZPShAnC6Zf9mAjIB/lyrxCF4UoVWfiReG9MmRH
aCUs/uE2zrSaNA1kqfnrV+SsbTgw5M5NKz901D4gt8pSjoa0zx9hq8isG8dIdCPe
SG+ozaMPsacxzuPEJab2ZXsFAYYHsCBvqMs+9lOs6OKYmfKe3o9P/Abu157BV7IA
J7IGU1/JdmIAmfJCMmffbVdza+OKnfY7jIlFKDHgjmqpATseyWbk/qi6WF0LKrN8
pGCRzbq66ek3xAxqkDjW0wcUwwDPm5seA9JsdcP0XTVhmxlgAW22fzXOjvmrNXHQ
uyBceLkVr9a8Y35Nc+ru+wQF8qqtPvaG69ufL6OrOuEheCVmMsplwlwejMQInUL7
HQ9UIbBiIwRJEOqRQ9VO3Yu6Ua1ZCGsGuwCr+CM4PY+YTgE724N+E5K/NIhEQs6e
v5vDD3uZ0Ys3EVrfnxaSJgUzAGhEiXIfdeLN9MrABkPMZzx+g2DyR8mSyDiwJE8i
zth0+y/pgBLoV5k/EZjZuDnr53jD/HKFOU2IyXc9e2Hx5BtxQzbIemv1u26xGzWt
Zexs5Q6nEXucWTgTsRsMQJoFIQqxB44nJ1RstG4wvVk7MepR/E538qO4e4rGGGYj
PVFcb1SeuuVFH1TkVhrpANGmAn/MtpzvV4iuNBO95kE0ljkHhGPmVhr1PDljOg5+
iQRwl61eZnfXzXO1VQbJg6FT93SyU9Qtc/nIlg+LgrPhiaYZGxoSa5RqvZAa9QJ9
FJhvZnhYNFDLSnp818jRim1l9wGXt0lmS963U/bOnGF50UAARiycPIPZSU7gkxWZ
K0wDW8Mm4QQajj6fa30/xxyeozYfbC5spQ766rw0SJyAOcqdkavqpQ/GAoG2Avw3
ZSAG2Ru9IuFcRZPtONkzrUJUEUb/h9NvVqjyTk230vFncLGQIcjbvsykAx1irOXJ
AiJeL9waqKxUqx6T1A3vlyi92ah2qzyqe8E9AUUPKLet0l81ebF44HRENE332qdc
ykcRADLojaUkfpgPTXg/b93K3yOnBh1g1Ti6mRTeigiWbVqMKrlheh54oE6UzTxU
28FMPksIwd8887B/u8ibAzCpSPCDgCWqf2rtxMvr+XA+DEIAr0K+R4ejXzPaRph3
+r498wzYbUkbDf5wv53BqynxtyZxF6O35iB16JsZtOISzMJPQdtH8db63m4gRhEq
4Vt6zBI70oNMhIQiLeKjMGk+60Z+Hpg+E/xg4NnPtuZoji/boWPC26KosQZF2HuH
oIBwqcvRVudERCrP1ZvxyKdrdTdIjKfykRM1T0Vbxy4aGGKixx8GeIlX6RxsXeP1
6Km7A6eTrKemO4cKTgTsMcqTYl2NZ+ioJpCtvDeNmiYEApyajdV7wqUJOj+LTYCp
003M6rpckKXVK4atLt+eWXWTBwyhrIaD23nkzzgY3vhLu7A6Z0EP/RmvPPqc0oJx
i77STyPKA023gMxh3pzLJVNL//ohTl9f0YNozRSxQLfX3g3bMy/ABsimx1l+56Nz
eNwOnQ9gLCZcMtw/tfwOlHO2KsJROX4iG11LKzL9vJr8Q/2jqBWBtJjCktoknAQN
Hdc5q7eUAEj8x6tQEuZYP86I9yhqkJXowrMwqcwbdvNuPcBjxFrmJE2wJmdwBok4
urA/rw6Dqr9lme71mhpFbAP8BwkrF1F05Jiw0Zj6qOoiIEcTQGEh1HiNuYFVG1eS
aeQApqRXoh4Q7zRV0uaaX0eN0V7Q+MBO8R03Uy3d0htXDvZwW2RL425Ovqd4aOuI
5tNh5MswdSpI2NJSnGprSi0omyuXmPf2gT06C+pSw8Y8TmZKFEZu/aNw76hk4HUS
rQ7AJ+GTTmimagNbQ4P45GhTWHOKOB+zjW6U/xeGVuPBOmx9YViDbHlyPOho2ym5
TN0N6EgVaJvOUAD1vexviDLvtKwZKnu2maw0NdpVujJE2zLHn9LIBaeczm2ELuBC
ttQ8ogt7KkFBXcBHEpnTZaJCFjtImgT3xvB2hrbF4A+IuS4259mK989aHUjZvXSK
/ZHzlMA+jGP/UTC4sBx21nSjd4FF0Ck+LfXJuMrKtHWjvzVqmQ0Y6ctG+9EHo0ik
skcZnGOpzQlcaKUTewiCNV1MjUuUq2abZKO2H4mWQjitG1elO6xUw69pMxHJ02y9
7fvIqpj1XGQ9P8vG+TpNuoT2j0p9JqnuU3Y4YwLsR4uVc7uNRl20db/gvY0cmn4S
E95ax9y/Y/ztTN0XUB4jk9ewVK45TLrfQ32nYN9MNWZi7cgtIfTN43tjGOXwogn2
5mgIT3lDkxLpTwWgnKqGHczhrHJCCFPoN8tiJmmPxxR0FLR9joQyWOJ46grPTCbz
p02EyYwn79C8GaJhkw9MHrvfNs4IyWwf8a7CKgBHNKvN/OEX2LfAovPymNYuFm2O
aO7ryz5/FWfscaCkq/rP8dc/x4IB+i7O4M76K1yH6N+n7hydAV1x6er3fK96hUsh
S5Rxe3L7PaP6IGTRHLIaqourNemsuHpjx01m7acP1tL3krfJmY/dllEZQgQIAAsf
sM88a1BLLGOfTlZZcWKtwUxDPK7ZtOP4CEcjUMe+SHorRg6jKAYT05BcuYbcdIAJ
6l3A0SfrWmZ1mCJ/D1z5tETG/FMDvtp04WcZ+Zxbwn05Rv5e5K3d6q6oTD0jl+9f
GvbgdHsYNog7pHDTi4AsTvhP8QALwaHa95F2NKG95hsTwK/4DXZItfjp/5mKJnjK
wQBmct+wYLH9D85WIyvUSF4JeaFldpjazyVfbVXlliduJsd5/wWNxQdHMz9VrWIv
eb9GXrzVH61XdrXJX/EG+YTTdyGBhUEx5EHBkx5R54xoMJcyMX5tlsgUUuq7zPmj
Wv8jmpbwLkuZ1XrO7N60+Ky2n24UtWMxeM4mtE0wwR4R9iJ4SMd/Aju/OVKcmJaT
AStgWjkdUNgPdQ/CdqwQP2VjDm8wtcRIZENCpWgcxdvtxSp0edW/12nPN2TGC3nl
hHETtxcmZPGvrmMC3zI7WD5IG0wsASamTDuhQmDdcFbErHFnrAudtuBdLS/K+uH5
op4J2dz4MLuTcSR4qk+6oBL7SiCb8MiuoZOJlVlw8pnfAG+onK8/fw0s6yfG8eoS
iwnQWtnlPA4VwagSp+ubfZVCu1xQs+F/cB/KQ3eWJ/BO7F5ZEMMUbBNZm1suGHOB
O+sYbZ6sSD7Rdx/og8NtnCFOdG5rJHcVLlrN2JNP9TQB6RihpDPUCRGWbocqq3mr
CAo0e/JhXOiVwumAbYscexXg03/dy7OfCdeiupKiHDwAKmq6iF/QmRoEkP8+6Qp1
Qgr1yIRAHov4bp6C+pn1RT7dNo34LoX3+LG5cyJ+5E/lYqHBJe6ie1BHFm6F5Na2
IzkT4hiCqyk5BAWmgOaCWC4+ctFgNm+8+aWl2jPuyaob9vJ6gr63YhszryEqE13y
/IErNQP5h/EIjCMrJtyhkXGEqIGvz+Cc+8J/9VZLpN8LhyF4VykIhTmLn+VDI5zG
mHguWIfROjXdNrc08vs4PZZd0gy24BOtDXpIgNnIiHquzKYgqSBLWE5MyccAtLTK
V+BTYrP9zv0uJV2ZnuMmrUBqH+FqDUQOY/TIY6XaHxUzgIGwK7HvRK3eEwCUqgGb
Euf323mHi3WK1PMoPqiv7ybSs7WpBLH/o6vuIvdEmcdhkeRNXgk4Ig8Htf6bvS9w
dE8UEAGzTYTiHWfIo5ggn4SZUChUiJHaKfcOnqAb60iZ5CV6jU31Vye6NfdXceLL
dbjQoJ1PYVeoxnENEsFCcAvsMTFoMGy6OPN/ioj3VJU0squWd6xW+aRNtzYzFxmN
0HBiE1AaN8N0M3X7WWtzbZteUeJdYIRfdT2R80Gd+L8QQ2JZ5EPTWONYovi5NMsl
+G1Lc6+VENPFc1r5JlYoYRaSquRB+Oc1oC674ensmYSGIt5tS2296dXcWkTJ1Gci
bXGESdgmQC00xMTWUhpHdPOC55qJB7l3oDXTT5GKun5Gsdzy93h7cdQ2jnWC7eLn
rezJBYPdLI5K91HsbAwzAMfjnZoWC/H+2f2GASq+pQ3xpd9vMHeZZ4M3/ry9WH1T
R4kEUC8gA6EoTJbYxxhwAY466Hg0qm3p+/FJzFGDZsQZOYUBj0okQMUdha0AT8L0
LrMUBqlWGtbMvs218KVEEAR/Gky6b5JK6G8IqwS/CVYgi9r535E7hyaY1zsHWsF/
ZaJYKNzsLjD6ZOFCkF2bsSfOK1UIifywVcOwdJknXUgdRm3jeVZcFXL2GgrXedwB
mQ5YWNV+Rj2dnBx/PmrGjEtCvcHbE7yjW0Z+j//AnBD9n6t1JAPO06DmjDxxYV2n
fbFI0GC9yIQ+LaHeI8cYr6u4dpCCXLEHBNrIjlfVDaNBbsedvoeJAqgfMD4j0Ss9
f/ELb7vsXFzDIN1w+l5CJ1jEnhz6KxJS5rN0Ej8pVqd4jfVXw8bz2hcPTqTc2f3B
QTmJX0+E0OaFlUR2PVXBF7lJlrfVJx6dWV6DY3ERxVHwNqn08WuOCzHKpf83HcwX
S258rAHRLt9vBqV8jzYK4jvOWwetfxH4jM4SHwmcIXSesR3yXWQTII8XzQ0pGTrl
ovk47GXOis6dfT6a9hfp1G1BqZmj1PWOWiHM1BubKJ1e587NooPSynepjZ87XUGI
bZo7NyZTGCE61J2JVL2Bi6FhOXZE1c/DvasDhDaMFMmN63ICdO3EOpdIrL7hpI/3
vZIkkTMoBNcr/8o+7KimzbhR6jiQVyYhPcDHDox7kn1UmDjR4nxkYZdIMDgukLA5
EquYtYxuJVebCWfKYrJmtrxKcSt+XI15tP0gQdZlGl8VWr29r2IB3F7eznitG12e
bXGvROp+LjPnTCZjqCgjr23OF4LjxMZGgnqdUNadDGG8votF+XxjR3u70Haf1G8J
JsjepXo1VNhk5kfGerIIK01i2nj5jpyL2wjdQupLd0fOvQqvThtlch/lbzA9yQGk
kAnhnQRCF1AAETDT6ypt0GlISgnmGDNW4PXitwChfSphdyNuU9BXxX/SiQPnwG/g
qQqmHMniidM27ipyMaBc0ljBds1a26hBS+v6iJt4dHI64IQEiH2ssHx4XB4lE8xT
I0JtKp69RyM9kXJ3d2AxLyQw0L4Yf5a6paJNjM20gS0HrbUErpCVDClju5hznTT4
juE/iE/9XEMrcj0kLXBxFiM7zD/RX7RzI0t3QcsmZWY0lfB8ZS+AT9OH+rotSbTc
BYPTg4gp8hvwi+XW5GHvN6nlAj363rYNv3XlAu5XWUI1Z86g5quEQA+KquBheR+u
70CQtszv0Aww4YAnMoruMIFxMx6FCe45WsgLncIiXSt8yAoaS4Wpz/9va4BK1TdU
BEZfma/4PJ41wzn5Kl/0V7ctYNfvNN+g1XHa/pAsbGxmY9DNprMgkLYeBbfMuaJU
wbUQHe/UKtJzfw5McTVpE4KbTUCN5luUMaaYxNToiXJrKb/hZLdOEiIhkSwVYs2C
prHaqh+KQ5X6Ko+wvkWcCOnHgD8CcVgu9BCU5htUWvMMh9sMTtZSl2kDRGqoVQbM
HLdWU/PVgt03YEbD9TOADHihgx7+OvbpmnX9bdFieoEUhFErp9PuCAfYEF47AvxP
ju3B1o6Hwr8sPBDM5P/X3gHwezuqBmdxc/AeVir4Ugw8Hug0cTyISE8gNkN/+5Qt
xu5H03Xf0kmzdOrnhXAOMmTI51WCuh820+huzWxKcRLFV2JM56TuvKQhNUXCP0Ms
JzFHoxLZjmasU3LvgegU7pootqP/aySsltjC1vMSUB0ovby0swXo+1nBch0GcgtA
7xr5GVeWEG+LQ41Zm1RX9GcubEvU0fbUujdI65kOlFltlKvJddi2I60A8JogboUX
cAhnpdJfey+O1PmcyGzjizPtBRV2jMEwBBoqGosXrP8/M4i4SQGUAABI3ZlczLT+
rj67VlyHfVjf2Q8Ro8GEn7iUCjvi7YYlTCRcxeD5UkWTIshZ7MwN6JpIoNa4ZhxO
dliS6ogDjZG06iSRrqHJvH6oLTs7chi8uKYY7YMuC/K6eIZMIbZqADhljXqGQMAu
/Hz+S3v/F+0GTBSMWrLqRsSo5DxktKW8W40Ee1aDrEn5krhgt9iIUkotphT4nTCF
NjIExn1Ye4fT9t9MOjPORiHjxC2M0ohH8zxz4p+mAgdMzGiCka30ju65Vr4P7efK
IKPWPibGqcSSlBTWTGAskpfgjXWaUWN7VEEYwLOPub1e1DZLggwPlTnhdyHPHdyE
/ryxQAO6SZFC5uYo/C2+XcJmF3u7iHEykFJPlFB1X1ZrTRUcqaaPrOXGyTuQaYxW
gv874F73LgSQJzhpuOwhgZr1FzNt2VF9sZ5HKsR9GNwqO15JnKdRmb3lEQQ+PQCa
HFYpN/sgcgz+aqbg/+HSa3z6Ca4+GVaNNoMqAG/CZW0XZTbGdbCX+rN/fnecXztY
IMOWeOc2QhaLsqW30YZgBbVL4jXVzrZIvD5jjjNVcZ/B4YnFGenbElAhgZlso6dS
mKMsG6Wt9Uvx73xmjAmCxeax/A2WRZlBNYj9vr8gmHJEe5J3UzD5FCJdtNCeJ1iC
CS3l2uCzSzSaEyX0bBR8MXUn2xA+PCxXsQ/uqueSiwndd1GmANxNXT1+M/4np8VZ
vfJGchCwVfZ3YLmC17twPgXg2Dcxu2ssl0156K5VflLKBZ+0hqMPu1tKshnCJF8B
mVsk6dblO/A5ugz3iSG/WLudvuCa5u5ta1tS8NtxvAUfHhOVdMg3ZoMbETkRPbab
mY5dG8ewpQVj5RzYXojl59LnpiFyl/XroDL37nbY7G995O9Y8v3zSMigVZYQF4kL
Nh09oP0BSPbzrXfpbU7GsxJzeHiTPOyAn4nbzh1Tn3u904C2Ggj/nxgXyKXJZfjs
KpXk1XcHUr8j+qRLPmJ23aHQVgEn2/aHmXMzRi/bZyNUHKQ4B1b/yZpqHUX6MdI4
7TaFv4E7LacK05uFDRzlfgJOAauWildWeFyfeLybkrwFBVXP72+t8qPVd9etLXOB
Zwtbu3shi0FsYbdN/yw4WpMRoye7sIfBOn5eKL+N2Snb81JWCkYKPzLqCu13jiez
g+J+lM/drLJwyUxFCzLbXR0cAavsr7NccjeHVHNzVvQA2PP2CllEmnbeovZYpUQs
DuXwe1AqjXIE/QqDG5GVOecE3RBF4F9bLHeeh8RlBCoS+r+z8TznXLuuo0ah0C09
n2TLvyBmsQPKszJDm9l0VdmQVt7+VnkI4LjniMDlIMsSiEndFamWnbPF1AHfgLCp
qi6+ckM82oI6FeKcgiUq4Kkv2lw3gncHErnPwcLd83gycEPCZW8vjA/oaO1Tg3AG
g47BEpUltrXNsB/QfsQxBcCr1TY7rJ9n1NyhRfGtlUp423+oPxMw+EsYzAw4HvOY
BMc2raiQzHMlTqyZVHMTdB0zUP+zYtn2sfB//HqxHETdN1oWWlfZuS9u+CEpl1K1
gILOd/+2UOv2MCHiZFgm0vFWOcSj81mpgzuycie1a6UZHKoOEFyeuGLpM+ShKKZX
L5PxnJ/CsTDpk+21t0cdJUUvDnNg3XH9xcDKGrtdShFcWlUO9Ra73wFkdjRkeTs7
4D2D8XldvNZPAVgoykB/7D5bTng3sZzOpan8qq6hmqQr9IO2ZFulLfnZ61NsYca7
qlxtDAf9BKAuQexIJEvczJSdUs1hyKXI5pTw1lZmQf3wstRSbLCY97d0TzYmBI3B
ZExseHBMESkjtDClDUU5FOLJREGx2hYOuqDknMXhTYiZ5wD5qj+gHkIMuNZegqXd
LzQIwkUJNXBYsP1xLOhu2efHwza6+PY0X5TXk9etAphsqZTQSi7ADxxmJ/aC+FCD
e9XHFcl8zCKEVvYSu0Eb6KS7mnRZzAM7/GNwTyC0WZWMVzj9SoTXCgc5MVSOdB0o
H12NE2we7tdJmobSXRv3w6ImC3/8ownj5FMNawAlRoZ97LbNYAGM9JD/Wo21VaWp
w95ib6I4BSQUw9dD2hIvto6Jtx113L9xH39ESuhAFDeNf2nPPsoDenrql/Dinjx4
1KiYthPOkI/fCTOpJ/yvcutR516AMpA5eoZA1Mge2HlLdRz3/L6AY7oCTwp0BxuC
nD3wOFh65GvWIhvLTfU6IkalsTyyW8ywijqLlXAWilv4aG8YdjVjs/UnvbQlBwZy
yxGB4mUdBw1VXUvMHDISn8GWeP1rOpdCydgx14e4cHlMapcm8FX6JSsBzsIqvcvd
HUAoVktLd8z+ml0tIFyIgSfbCQbmetYcy+WnfjwFculpboz2h0NSHpd7ANM+gEhN
r2FifWiLwb834WtWoRdMKx/CAHtIcxP2pkUdXjUZe00a/sLjL/NwWP8a8kAZwT1r
oY6vtbpnKPFUjzY7MM9nr8pmQeDsMO03sMsCyPATceOViVn8/TDMHgFEMAHKH+tb
YlSuHCoPEnpqJjJJ5VaRtqQ25uwX5Wu5Hiy3q9CvivIlbpiovzwFz4Hqxcvv6IOc
8k01WxRPd/1a2NCnui/2NcbnIXg1fekJiWGyyxJvggkTwPUTeVN8NG5BblE6Thrz
wlW8Qt6mCirSAchMSK7RAa7apB07USi2UDP3+Hzc7jwDAXywH5WpEjcyi3W45jTG
DhrsGBSyUOhGV6cNbkoCJvVcD2p/Aneq1bk6tiSC8Pk21f/4CBudgnc2RkRGTHpB
KzKf/0f8phB07bT3LK5PQLF9vie51REBQIznBoFAsvfpprk9Tz6xzfcezOBLSiIO
R/RrSW7TpotYcL1yNXlNUpZbfNx08ixB4V4GUQ9pCgWT7EXgZcK72Wtpx5DcgET2
ZMFNzGK+9almZx8NIPgei3M5qg0Yu7W6d8YRduU7rTh1WBW7K5eeOaeigVbCaHo0
waOmv0D0Uvqs5ugLgNJRxHZrYxSqc3O5lk5fPtq2+kQbQjKg30ihPRDrQXIswBHe
fh2vm8ENJAMVvKJR9b+Oty+AJ2dd/J2mi7LDilGRqf/dA+sSXMfhK/unZVgsa8RX
YD5GyCeafg3FyKWRnjTWuKJsxo+fZs1S0ZaSyUG30BIgkmOZjYmJmVxRNqAmQzTh
5CtjJkDfQ917Vw+w6d3YPZU+M658OySYC8t486ysNEY3E/LrryD8sbt5ZGE93swX
2Qm7IA3+CAZ39CjSZI7gbAfHXg7aNtvKQD1iD7OFI6rbQx62QPaO2w1oK1J1gdlv
B9VgV/htgjafJedh99B1LflhqA7dVwzy29VRxzmTOWfVO5oEB2RM9cuimSCIi+Xh
EEh8EkC/jGFC+eFoqrd5uV6plbdhlXBpPiDJpfTyJis+Cz7NAmMRCMcuT72ta0WJ
s8FnGcBCfgPBJ/c/6HYy61TurxZerNO8ioYxAItjXvwcYaCfwz68fOR36nSz+jgt
n8K1mQYg+cCXmwcg6r9j0mJNHjz0BDMoTB8KfrfiG5mQ3So6qEoKuFkacSqIZJVw
+S0berEl92Lzq3Il5SIK7W5Awb9zVT/LYIer4U2uCW+hqdQnlEo0DcDlhexX/uUB
IawHdwP15xY62bxQ9qDrNnNODESAQkwcDAmoYOvk90SR79gjVAQWn3sdZOcm0NO3
RElVkn+Tcv+SUMcVVKG+p50mPhLp9S8kyLvyV9H8y5y/sbNfCBGd7DeRj/vxYvTj
w/r5cf70knfcAjQHE/T+k5aCKWe82W4anq7Ld/cbwitxCNTAI/3OLVfLnL3CqQLC
Ja4tK7tFCDKfBq4VzUD7iObdFSkJq84nSdvHwwRkfkxvIs6lgvj6cV4GD39N/Scg
dOadGWPCogAGi8GdR0V8OaOfmYtf7iJpEc3FxOXU96x3UxVKTryVjxWIYR0CdQhA
ntssAWiXlkXhfsOtPfBU+TmHrcwBYTwGp6ilxkW5UMQ3a3PFArS/NzvPiwI3tFho
GD2QNd527RXe1+JvWbsoy71PWNB2AhqthRx9k/2ZgBay2fqftrp8TMkDcWnOrJmt
bZqZGOoohB02OBeU1PcxhBbTOisbm4E1oKa4lB/fIPR/aI6GOtJNT5+jxsv5X8Z8
vVOyxeyYAKOxkLa+/h3vwKkZjfKYk+5yEWSo77TRe+kFXq+xGjGMEdyaf5A+PBlL
SljxDEqxpXgrTB6w0hk1QYsGCN/PwTdOzrFI7CfZlyg6pZuVvYw7rygmxG99SZ6a
0J5ls0nlnWqiOcPcrKqOijU8ZmxznEEkk6iG0SemlY6utqFGCnZyGbpstSr82tNI
59lKpMkqr7BfnXnrwxanIuS/9I4yt6+RJuKjAtSA8kEm3tvghWI+hMxtO1u4Aqqg
q3ZpvZn1TnEWL9ItnF3J9pODFFwm75wEnZ42oyvvenFaCy2JfZGEEYNbgudUGoAW
DEeudVkiRqY40qFh19BZHYiluGBCFss8qy/NrxvqhTRcsPCkdgh/v090E/ThOy+e
sjLYt0+dZ15dUu5osWUQFbC2EXPh+kM4qIjoancVmLuanf4r/kQMyxbgy29Jc4FP
qS02gdge2apE7JI7OkunebNj7DvOkSWu/vMQeANK/KTjRcDeQS/+uOCCKinommxd
yQizVtSzW5We4n0hwAD/a5mg0OBeYPxhJt9EOKiaoUETmDZaEbq05WyTg9ncTkSH
8oIVQKiPtOKKMx6G5br+tGx3T6vKZSAg4vE0eeoGigbRTnAFU/TvMvYdkht9R81U
kQxbt8wGj//fO62w8rwHNG7KbqN/v9xfUsoOXM6qpz/9RvEcQzif7IEgMnjonqML
5SOwQWIDm5KmgRrOqbFMk/3fSpyjpeIrr0vM9ezRW1V99ii4vAiD3ZhU+ciK5NHc
2RIZdwGE4urB1cxe/NkVssdo9Nzi5Ulx5lFVcxWtHG04pFnC3NypxO6AwsV4yobp
UZwZd5pi0LGK4ubK+0JFtDQ7cbe/65dvhofBIf2jZylRJhswhDbOuCcSYphV3mfV
ufSVT5FL5IfCbZaht+sFFYq3eTUi9m6h4VqROQObb0nt21oMHQsdRGxkpIMmyx3d
Kd2gSt5mY+1/8g3gh7YtY3sDZDpdCmkbiNnwPlL54ByCN6q80SpiXVNGH6Gl3DM8
SKsK5nqRF2ToSNooyczY2UoNStlCeLRyKD2XLf+WzQP+gkFdsAFlgNq5S1Mr1PFu
ov5qhjn4GUKWjm07iL029l4fCacJ+wmSDNDKNqaMHpRlaGHO+Qpsb+kB2MCjxpwl
Eb/z768WMqGQfKVpf8r0nqe1ovUAhlMie/bFZGLsjiCqAhoBTK2JRu5b9p01PPjZ
yOF+Khl9rernJs+c2Dp4T8ALckdEv/K6KBOcmqTM1gtbrLaD9W+rWgq0kzmCqrz+
izzMbYJOsT9RmtLuabuIlL/0d9hfMDSdQ6INYqSBcYVDf3cm9C7xUblspLKrdEEO
f+4uWGpNOZR8ZbIAiUf7oDmp4csrGPgh29gB7IpxzfL6QdfMzIkBhvmjo1AgFueK
xY8QplE9dZCzVGvXGT62TZW6FOKmj/Lo0cveQYga0FGdXNoJKOHqHr7v26cjskcm
9zRKPd/DSnsVTRnvtzuaHAAZliD7QKeE/mDXpdeV4FvgtsS9UD4yPlBnLuB0bJRc
nNVp8mKaz9KQxDDEdXCVtfnwJ4fhRl1Mk7kXzInNX3IZgjNdClvTgRryRz/Jvj0q
h7TwvzCwgMz8BAMFF3CpE29DjoQ/KgdnOHeHc4V9+FKgiomDfJvvaCUqGCmZxnfp
Njw1GdiiKYXmvx4NXuNw2TJI5OuP0BqQSUjCLYBV1aQ4apC1XY1zMp+z46aLZyQ/
VPfvwsE3QOG4CfiA5OsPx19ud83UXFeGI61bqLDBnBPubwL3nHgarfyQOBqgKFSv
43If4KHLb+NJUAZpe2sxOtMnwhudXsS2QoAOIhK+8xs7h7c8ktbizQQHyS3xagC8
Yjl1OiVmmyVxAcj7liz2Xt6yKOCQZAMVAgdSV346Sr+LmkbfbfQAQoecFmPWK8Er
Bz24Tv+mdQobkZXGefL0dtLnFBhzn6c0YGCCdLzgM8cGNCa14WDC9YDDgk3TaiSY
WVl88c51HgjteMRwkfPQJ/iTBEYMTVK3mQmfRRLSeEmUe6SuQlx01AADtNjIrqt8
A0yRronxgpb5hoGgKqa1P0ACyweD8EaI8XW2vEjIDyENEvEgXcxEMxS0LOpAoQdV
q4+OP0Wb3i34ahwPM4IBGWCDTAvKidfS8lgteib7hmTU54iAfxcCIwzBv4Q6HZxa
+nJ3malG+Z5Vs8V2uwT+YKJQ6V/RLq2e/GsxwvBM8AUROp8/UE4eKKNmuvYxFqfb
9vBl8qbkS7tEgYhLUpUO5GaTeBGRR0GYECbYXIzpbeps3rtkhnISE0SJwq/o5K0s
7qi/4mk6mlqGk1EcbWu8vhucATXLU63uO82tquuQ2vOBzsA4aWcBBMVzTARWpo9D
Jpnvn5ZfuCg/pQZ3+cKjQQlu4MgzK6W4jmALVaBqoP5lYKf/NVGfFAm3Mgnu9GrW
CxmXg7VVdlezCUyfHIkxbzqMZXAlrCMwX19dRmA+VXoCecEZnWdVYlxRPKZxzN6t
NNcllTlJF/nvh8mePlWWTiKH6n9+WeDyme/36UiUgy9VPYZA4MgCzNZlQ1J/EK0v
FIbPDkE1PPvWWwOxvn7BmzKd/ydOf8g4PV+OPA98ROWox8l9MfPxz2lqcT+PFeHh
HYMBWIzK6bHk2WEwPMXQhy5e73cmp3Uymx1Y45v0qxdaQJspNnbi+/zvI6Dmwu3M
bL1ioU7posdkUdDI4luBFaDKvLqFUZd55p44eVI+Esm0DRaHVUy2pmMw3aq0a6/X
D7H01kF0bUUV0lyl6VonVG/LbRTlI2SMFHiRs9ctxac6lVJzs+u8YCBExus7vkVN
h69/DAP8N46wUS6L69l8z+B/qFnV3kWiuKh1nNaPTJM6CSdqOqTKGIbWC6D48KGw
rmHp4jXfTMRTsZnt//bpE7Ajf7FIeoTZpx84xJSwBm7BxYxs8UmF0Ks4uSq9ezTf
vRyH1JswryBpY14TwJBqZ++MCrix0E3r599qnGxA6R/EURFws7Cah9Cgy380mONq
1VblG05CVGSJTJDKxcDquVy5WwrAxe8zZ2DuOqnGQfuWHP6UlsJAOr9neim6+2wb
uUYBCzbsJykAIsQpPzuT1VktmWnvO5JpsD4z01xxWbbzZzh+989TjTzbE03ZldK3
fKBXTCJAET8KXFrKqRWA8Tm9oH3pMDPppzBasO4bytVeGgAS1YEiSyu3e/UDm/Rx
Hh+Zv2an2oLm65RC3GDgBFDl4+LrvPqi4OuunULZWR1+BiaCSqCwZpQYvdW3pZ6G
06GuZUOgN6hISfHmD5uWtd01EDMQgluVxsf/dHc7jKOX4M2y7bvs97Z+3Wx2oMn+
e62Hc/ZsPikFS0laGpKwJiV7klrjwyvPebnTJb84Me21aPNJIm2gIFdglK4pbWCW
ojC3gVgvXnjMo7BAvquYNMv+FwirpGr/zbafKJJSJo7wB9ncEV0lbOP0Gxxtv7rO
I0kWp0g42HhjiiwW4ty8/h4pkWvjKLvIBp0d8gella3pO3hdHIVt/lwSX+3zV86n
lhYX2RRa6hg/GgCtr3aWwfsZrJkV37Qhrj2bceEZJIWEcAYH8dTXiE00/ppk/YVf
QSSjdS3o7DlHaUnhpW7fgvnWnaRTxjDh5i6uT8OZQ4kmbnRSKfQv2LpSiI2UbF+Y
TXFuKmLOUibSifAklKP1oHqOh1ANJqSrpkF3puEisXOnngSOfTGJPKY7SMqu7hDL
y+27Uxu867CY4I1kce9JowUeChdsHdSaRzAmUESmwnujizf6ddlWzHXAd+VEc1sw
vm4HBzOAqILVZVzZGDw3aya67li02InWU+FhMSE+1yw0GtG2VTgYBlMsERLSUOnC
CddY9SNmZFTefkHb1U7wGEQeFrUk40i6CTgkphuK4kxjoSDDIgnQpCKLpY16BGOI
oEadOddgYO724ld4utdw+K0IAs/K8qo0+H9KX6JFCgLKibB2YFeoji8PiGy8DHSo
JtPbIiP7xlCU8rfKxCdpJviVTZ2DmVQh6WX0NJ0cVzi8QwKk/C1B4YNc5Ta9ofot
NkCBSOH6zhS5ytYe1SyA6u4PDST/QXI4wg+IdyjOHUhaBOI5ZiYKXI6qa4qK4Bjn
u8Uryho/5mpnX5ErsIyPQ6vtsUdet5nFJyoYStoGucfSGHnnsr8XeIXigboUXVNc
YYPI1DidDYivbLD2aOYFUb2h1caYfL6CWNwnhu73TBQOvrGzu4jj5JVijdeco/r9
FsgIqzt7pa/LMpsDzWP44QelA30fUyj9q/pJ617gFr55k/StyaJfyblEHL0V480G
oAW2pXsM9YFPh8EGa+eGGULH7yHaBckleJrfmNbhPrYTULc/zc0N2FZG4+pCmbeX
P6bnB+5sAbWpgKUR3v+bJfx8LnKekk7RMOkl57xFoLlANNs7/uXUonuw6k+/6zLz
N6m6lcDeZGqLjejCZX+oXCvrzTNb4t9XL+mosK3iaX8GWTYv1hSR2tMoc2xMAwMu
C6pSQ/BR+yv97BAkbZKC2XXCwgZYT5hAokjxQbk/DZoo3WTv3n9APW4+gP8nm+JD
nlexJtaGgmIf0DQqQ5c3A4NQBikQBIIOquuiBpUuMS8DJn8I8D7TBTgTfvS6ZW/o
jMN/owvILnlhmyglC1PXAbYrnQ+M8zBpimr8KiiSq+R60rAlCoblC6/ZT6OXXGys
cZWUQkBdEfRif7lncK/zoPzpIYlsVLc0nIbJ5/JBGLj2oYhWL01Is3wt44K+PsrA
Jwfq3YapLKXqauuPaZYSh1s+dDY53nXdpOKkzTgaQNVhvFtK1riHDUr6hRbeKeID
yYmbsl9jL/lCRVd1IL/VxERcNBnCe0Iid4p50mKV7ikJTqosY/u5X/EgJdwBAUHI
2pW/zXYHFN+SCpqPNaUbgqvQRt3ybDsTpxb06+4wiu307btaU197g2XONNtpMam5
g8ngsUSwFgtd7bJjplg7KYZaJwNBtS4jMwb/xeIggPejrKuiCf9OIGpnBoyAucbu
Y2oLzFuWfmQT0hMhrtbPVDGSKCggrnOsYUDv8gMC0L1R5ByWd3arbWO1oG1f9ViE
xdQdmgaZQtgV7CDgvK6dJZ063Xsh0vpZrtbbjWLJB8ilZjmCYCoqy4MAYN77yPmx
PoZqvTkZZFoOPUbGOq5HvLir/x0ONPiedlpLH+tk5p1tQw0s8VIsiwTMrHLLNOFj
DDknXgmMmQMtQxP/hvCorqZq54GpdcWFyyJbt34qhBSW0e5LEixt6SJpE20JwqxA
c+e7WTuspLrl9y4wD4ndRpFWVoo7w3dKSR/hvzYNgH1OzQYHHMNKCOIhd+od27rS
OAJ6GDFmOm6aHh1SrG9nW9rwBE0aodNUYAcoTwaWLfvOmQ01jlD8oddRVSqi2S9J
qpdfAB4BPQB8SGKm4llVtA68ZH2rI42m1ozlTo4ACHan2OAhOrjwsHBINfYkj5HC
QjubN8nPjZx9ChqDTfL8++V9TW668wFGdhyfqT3edVUQGiuB23VfMuqgvbPQ+O6s
tuAOM//5KmXRZ7R/jgdYGop6y2myFx8HOaxO9p2kgTkDq+REVPWKFeubvlGux86O
r6PG4vh0jtv9/vQhTQO6puT/qAkinZ/nP4UFMvpGfSKqcwQCJCgzxDgzXAVKk3OU
9aUp/xdGvxg+IJTqwppp2znLgSt8vyC9dbrQyOGBlMToEPFykYa4qYVbBZcS+fPw
unT7CkScjlYdQpAsRSUT6H6Y2xN3oc5nl6AeX8VMtL4E3gpSKq434ne63la3toZC
WoEPkW1N4MvhfzhoTFWkgGsDKoo4izrQmhlXOKiIsGbYJV6lR73ReDReF9w5tsL8
8KND1rgd+U0qUk45FIdCFkp3hinjRxTfz8H/mQO6lY8j+x/tC1EJ13rXxa68kZaI
ynIoQDhhcBwrSXuxJLRmsMmHLMHBu4ZAIV0xYiYx+jm22M2F6i/Fm+Ak9ePAAzax
A2fVbCJyqD7cqedEYYZKy97H6IGbIQAdqIOHOGGglQt9dGF8v6/X6sOzk89GpuaL
YhGOQsbNUlPmE1SOJgsMGgLKMQ0z/7Vw+kKWL3jBdKWpxntSnNSuPe3qPB4QNgwl
w93G360UjkB4ssClD/zg/AA6yTo+HyKLOLu+5h1j1MtGXIASKNF+PtkOPf0x9dii
DP3TV05FuotuHBGvggXLuvQnk/cc8KfkAPgGAoSmPXrg7+9P/UgTOfTg83mftmFS
D7PdHxgq4ncCrlJ81PD2txzHA4WVpA4B1GegHOsYNwFZ0pcFlJ2o4wP5/Y3DaKrQ
zUr5o5raqfkZOsNzNjoTsU2L+X8IyqslZYV6xrWwwTraOBPVNCYQsie5oozyCRI9
lR93/SNJdZeWviWVhxoM98O7h/quXRYPeg/Frnyz9COTxLPpN66ITSUHlb7sMlKp
hLQulsVR2ZXZ5wMz9zu7lvfQRhOGvJeDRkkps3kY67GQp75gOAe8fGlulaOO17aL
PLS0uPMUMeM/quhfpFapdHh/EBUMU6j8xspTjBlKCDienoYpknVmx4xFbc+QPOzb
H87l/uaPg+SPcc6blGY6+DpB/l6S9e5W264leKjVZyZI3y0RjpJQvK+cU0ZNGbvq
Rk+oNVBp9IYGG4vQRyLwTPfhh1M7wih00LGclpLSPLMjIXJ3NOdKV1vmQ19HQqCz
sF+U4nG9gKzFiNHkJQAzmdT2TmtFm8gvVcCZUDW66PzaV8Ao1GXwKLhkBoS8aESc
qdil4spNduw0Yydpsw+UTw8M3ubR4CDYYjJ6MTHKmwGS19yTnm7qHDrD31ndSLPU
BOQtq2kGyEcfIeWmES2zqucB5mhfvGfwxyjKCjUh50iI30ByxrSEiRdWXIT1UMzy
7AVh+9zN0YFkkGkfd95xpKsPRcUAxIShkMHRpmzNvTOYrfNpJvuHuI0aV+OmGy7y
mV+r+UdXrcqtLvN7+Rabia1mRvMVzE6rReIfp2P7CSdoNsaHqUUVPaYcKklP6uTX
2I9tsDqysPXNkaxTXp2O8yi+s8CQw44F1bHMIwDg8ygCJ3DKQ2VWlqaratj8p+6s
20Mw/DCDzGgI2T8sYnoZFt2WTOCURlR2R87+zKGW0F5fxZfHCZS1QOCeqoHAfp/M
kW5lxNgzfcb+QX290rPmvZPEgFOk3yl7xaH/BDftTs9bL8wT6IshX0wSIvjt/U3p
b2R91CwrqpvkgMZlCZHJSGVZOFwVNzmb46vwiS4pYtOd5Ohyv8Z4aZc8ia211Bl8
KeblKqFnFa5vXBK5uOfwoyVXygVNfiH9v1oapINrVCVnASoQ1JJmV6RRnhkt7rlC
fvEidtf9Ukve4O68CabM4MKjO5uKN/L8SppL2njBg+ss7kRMZX9TKMYw1BPlEraA
8QoGv/jJQFIIrOKVMJCFHPd+dzsP+7PPscxMqoK/l58pp+aH/I71nJ/OmnXoukjv
gKrmcYwkvs6PU7/9ZnpymUjojQSG3X7HjVI4qOGl4ny4XYwXPa9B9gXPL/H4zwxm
SrcraB4QmpHlgW/ABNmBQXX+YtIpgEODZ/+Imo1LTXVkg2hWBKupe8hAgXCcmHOB
V/5xAUEWZf8oLXVF65VYC5CUz388N75lDBhEfkhWUyHBP4DdW6YHVLaT8fke3vHX
crj0e/MO0Y5T+MnejkGeF2p2IsVU8lYAl6rCvqFVU+FZFdlQccfSwhx5q2JUjQ0m
aLNknWU1S5CoIM3pK1yO4aY0IjNFuGvFfCP5axzXaP3NltoGQZatsAJl/x0jXr1L
3WneV9Sox1GXPvDVCNJC//bRsS9OWfdW+80B5KlfzQkUYAt+mP7EVKisFrjGzvDT
gqRQ3VzGAP049l5vpDtqOyv8pBKDyRxdRjvyKNDi3KbHf4R3Bwt1s7w1jWuI3NbY
KRLm50akwMNndcdpj7dXQxHl/YQDKHhx9o+5fdDbPjh+hRC139BbxD/5XGutxtuC
IX9cZjvQaRrahbHSVd1wrL1xGojypt1nBOeuy8uTQAuRuxL+Ozl1AFuY8Cs0u3jz
RsLeJFphWz0uutSWBNm3fetIERzQCEjNKVqmm7ptxlHn+br/QjzQ3Pl3yZVs2epe
dA4sAcdcG2SvQDEXG9qaMqGROGMPiA8WO19y6e33jxIX/0+jYWA2xjAc4gybYRhm
sGS3ij+cu4XA1kI/Pn4bWhvqQi2ZZjyMcWwiZjooH1tT7CpzG6NogFbbCIngf+MA
kmAzaxjj++U8Bc+XkJIbm/Fi4fkPFeUabU0pSaZWlo/A4Eg21OY0TnPqRSj56IM8
kwXQ8lcrZy1WA5CwunCF3fogSBm2D6mnlHHoPJMOkv12MBj5kom2fjMz/QNXgkTB
djy5v43qJQhb7E2LCGq9JMXhL8VwwZHhmu4Mht48Nn9GlJoodaRYroLCCG40G6d4
c3xNsqPMA3zewxdEWCu++apffdDHeDPe9yzbEqYm8uZPUCU9fA5otyLOxn09WpjE
gzn+qZRAUPOYLzECB8oYzF3AX1EaJYJcHvetS+516zcdpeaMd3Q9LWKxSs7YYldy
frL9FEB9gg1LrR4ITYIWlkOe3oo/bSdLTbMCsDxnfw0Sc1Rx8wCZ57M4p3qKsRP8
64cZZH2I1Iax2JDVf9KAXyD7YheXrq7K6IpDKRZtmptgqlbM+C7VbkTPaKhL4vSy
TBDBpB8dyTf/6Xe8aKGIkJzNek/SSKnNfuNGAfZAwqgouPXO9dyQUNGJXcnc0HvL
uJjeqfJUh39bRi01jknNQ1P/nDaSO+H9/XFIia4eIeiyx0UmejsZQlKAqxne7Fas
8lJIN06ExIinbo5R/41wyFQA7vtLGGhrNE2HzGwy5m5H5ckJfhiQp220GVYT8GML
/9U//pK3qirRN4Brf/dTNhlMuMC83Je94xGE+Z1kZdGzS2i42dC6iznVomRHfTXi
uczjI3YQ0bwSsnxCbOG7intlzQVm+RntSNNBl8zxGpRXnbvlXW2CmIc8Um7aOwRH
EeEp6AgX4uV639sn6rzqzYRl37LEviR9lt1Lfq55rWw8uR47YrT5IKfHxSZD5J5V
B0nrX9J415sdQesx78SnfJ9ufClc01j2KIsC9fqkb+NYWnylpXM8+z8rtBMATR5F
tzvQo9ji2eJfHHCS7guJSW/j1Hl+Ao/4AQhdyVy1VUz54jH/bh5vDPh29q33DoBL
KAiwgN/jJH4m+UGko7TzuG5MfVgi2Tf9lFhNkbXV+Uc18WKgrABbQppn2rry9ndC
fJMdYCRMyDuKCb6f/rhmV9RMzRQE/Sn8KjJJZoRmXnk3uD53b53Bldjf31kKsnEx
8aNfVnJGC9+KWsSD5FPjd1dXgaP5Z2G+P0Gf14c3WSGFbcCVf2P5V+ZhpDYoarc3
++4OkTyXH9f8a1YQenVjUZBB4mfPjRDSr5fLIAmTuZnaNdnIYNlOp3eM9MDhZ1FC
hz+vnVoAcTW6smJHPsCNj1DApXjPFfFDYavr6d1GLwO409CT96j11R8/VFo8/Qcj
tPMGWlbC6MTX+XYS9crVeUeGpFFDa/FqcyC9NCxE9A+yAXQSf1bKMDfno4A/uA+F
zwXrWjLLizEUca90eXW1kQvm5Zo/ZIQoFFNVUlTBe0nbblugqsp3lLuabk/UxZgU
b4yNBQqFv9mlDzbIITd6axaTZY00IijVRe2f/Zsflpp+oXPpsBp84a/QggDDXoYu
6aBBRfn3nhOzdxoAI429mBY4+phBPhcDyOMTxvi6QkRC9wB6nIBvwLZwxlirkLBD
4D9+XxkAY/j4suxX1u+Zr0QVt0Rk+y0BykwbmxdCrdI+4SAsfzfMYY0mZ4kFlK4w
7w0Rr8UU8A1U9XzRFTZSateYYa4tcNql04qvbFRHQmL9ZH74aEN+Tf+Py4pJFbLr
DtQ+tE+Si4++n9K4D7bqxTyPVHCqc2uCH6ff78vW10nekJSByaERuOw7CDXm2Ukj
A9dnFwWMLAh/WBHSt72IznEO5C/qGWpKQ+RxIWK4OptrSroZr/xIdpFw3GPHLfwd
XIAvRUKBJztzPtKUjAEuXfCbYsg73C0+7BtGQrTttl6jG2AlKM3d5YPByPw1mCUo
Je+TIgaHCtqaaIDnyZbd1D7e2WYm1mDDOycBlyMsIydxZ+fSFenCv/PKc5fHUv+o
nDp6nH/7S/sFpVBFbOw1kZfaXJzRHyHZ8WMPUSGLdxxfYiMUYLce672hGIKx/++J
v/mCZphYlSkxBTD31HoaOc7E+806i3Kpx+gDNhj5EJa0+vzX3kEBpxWxi5x+C1Gz
LSJQVA2ncL+5pIKvvEUEB+5vICyLCFNKFzkhmfkSH6B9KiN7BybN9l3q+iQ1xhq7
KfB83FR/oTZUreMW6z7Q12KQJYgqoK9NOr9/y9s+0HP2Rcdh35bavm2J8p0bP8I8
TX1+GjsGbBQcPbAWcjnIGOlkObxHsqcSTHDvy5K4zHlZKfnDLjr6I9UxxdtTffm5
ho6U0ZLGA0BLf0VolSa/WChNM00ddstnrs7Ldt40M1r8IccQZ15tQdzgcG4Nlyss
7UirDfm9bA96pBpV4ea2nIC2j0mfMuVl/OUNGpk5AhPrQOvDVDGm8HbgfzEw9Ovm
p12s8V+VAprbscMssc5VcQM3Axp1drrIG+IN7J0JONiA5ghEmsE8b+OSCnE4V0Y3
1SNRhppeJot8/tBQVcxCRdzBqUzzLVi+KoBMbcCbdFojSCZW0RFSmA0mb0FA++Tm
5ShGzNCpXjhJt3ElLPoCrH3E2IdIMJ1q2tLOLNQKBnR1t9qi0+w8APGNaacdw3zZ
aVdyDraLPSsHf3IeNtwNYaIjaS634FQDVB5A9OM5RTclkBR4BChzDTpQ84a085sr
IuI3cYfX9T7pRfnnZ77p0HD4KruFtzayuPne97WAyuSGqgahg90odtAp6rBaxCDl
0A3A3XpJ5xQ4QWgd/PKA0SJEzzvj+Zuh/cUxP3Z7IxRqkiqMETmK34BBG+STRE9D
ECsgGAzzbCxiO8RIziMqHzIP8hKsOiwTHSyUa1kcg2W0l8vSc7ly8OvSQYtJl/Q4
51tux/0EeoW80jAp2JS20f2XdQe0jhxphFMsxN5jjwV+lZib3mQx609ANNA+0ZNF
3lQ1sTjhE8zZRPfLS/pmFWEX4wwo9awhrGZwXhM9Jrd/2zbP+zF+tsSIcJf/1l92
p6uLvMVru4z5Bzdksr+7eQXoN8hA4ZhsNsMtNaY8rBzuxo2FPK2Fhh2ffGyWQtA2
H9zczrzduIzvlGV7G9S50f+bhVE/QpgEysDvg3yVQctM1aqnIphIL8esQVxYb2ER
UeJUh1IbJLSk0c1vIK+kULYXGy5mMo9sC62debXj1DfpQU69eXbkX15Wn06IVcrf
ZC+oFO6jIbmduE4nVH7sNylsnpQUiKenBKvoD7BdkLPJ9SnfXDPir9+PG3UdJW1t
oxFmsslMXWoofsdzp0NFGwKnY+awYqaP06B7L5+YBOMHQqEZupbAk/K8Ish/yknE
pqGrhoAh4BTz0n5QFAm+eB1CAwRw+mc4AhmZ4fSKu8Riu+U8BebXemlbpNk6pZyG
5z92RhZS0M9N+CqPPR71fOR9lYb46ld16ul2qazSRZFN8ytsuwScRwnSPMe+t96K
oS5viM882uP2lD9H6vIQGvm8kJ764o3TlJWHw1EAh1xP8B42n75e9C5Qhaefzjtr
RcNl1GaKeFMQai4KQjL7Xr/3GACDM6N3+7qzO28pkSRKUSQafMWWv/zCDtgn8zGQ
J7bgHzkZx1csDh583Ig7KbJ3du1gJdvBBDhc5NAXVQfW6b/T8gyKBYaTDa+NKx8+
nsx9bobGVoR537w3gG+9/QXyM9C04gwXQ3+0sy6HfLX2ffU7LtIk8hSoF5QTC3ki
YhCbc8exMtmaOKWf21laCJ8x3PQ6VR8XPZog1eo4lGkgj6VGX3LzbR8f5JGnV124
l8Myobqhns+2e8kh6HCAhhELCOHfbZG6+13gC7dTs12tWfKElELoGSEmx1fUIsud
jufteT1OvX6UjMzIr/sdM/9P+FM1XcM9IuLTZJuNUSXgHr4mKH3FSl5GrCv6cxcv
BOc6mefskuNBzr+rf1ecCOc8ouW6VCpm1DfoddeV+LQseUBavCnSyk1618wx1yfL
YIHo7zBS4BCAEsVF+z+XB4yIx1lBxiz5IQ95pdOo557s9XCuZx0ld5xnqYQG96MH
xswN5rRY9cW+ZqUmup211HdDzxCbqifRtdlZKho19ZDXvWOXvuU03VLV5V3MhKI4
UYeNpgKzv6WD6bN6Rl7ch7M5AIsFVYpzDC7JWj/aewu6uU1SPBZvOzLviFaN3g2L
FEu9s7ScALyktk31DWrFX3hmbNfiBDOaNlZsS6DwLr59046t9zLSrR3qnTjZ19ft
0qAEbbjQXrqF9rOG9SJbaIEmq96VAljl4fVxMubnrtV6qIJ0D3C0jEgl01msGlhk
qzcineCDrAp7l6KCpEog2HEbcCYEmqs0/rNL8/aSoD5n3ZcrD3tJ5QdB9+DD9Tp0
qHFhEhunbxdTUroLhaOxLVkSi9mJUo/uQhMph/AP7YOt9UxU5nh/gtvkLICwwjhY
Q0Iz0BX1O5dnljJHk7hZqXBBL46/bmcq1M9/+w0lTrUJSm2GB4lyQUq3CPnlpQaC
XGumJEbcJHSnI6Pc87jWgG1qFKq08AyWl5H82b98yEF52gzTTjXUizc6DzHDUs8z
4+80qt2TDG4k+IQvqJ1qlUA21evQi55/tZL+//e7ujtX+3/BQVXySqos532+Ce0D
Lh5ydL4J5tAEZ+eK5/Rv0rc3hNjHeMHrVC/0vYfYajrTP7jMtAMgF+GxQXDrm7tw
hdHRWAc89qMT625ZVDAzlZBE/mz7uHl62noONGfqoQCktVVIej6IMONlyIbJnMaC
W4xkDF087tbNi9V++p+tpAIfNX7ZAV9xzlllfce1eeHj92qeOO+1q5bJGJieTDrN
a6nworNJGLFue2OpAdCkSpiSFc5Q/YuZWgvatBTYFzZEWWeTBqlJXpj0KtRuzz08
v3YC1LTTWJmDxICHPDr2y77tSDvGHR4R8EyD91/y5mtofnHHBA5BkyyjmXur8p0N
uZHOyB+wCsVFl9dfy9PqEf3ApGN+cred20GVvtHWHRi6sgrnc0Pl8jhCrqQKuAPr
w40Rvs8RnRPyeLfriORUYvrHcT+bSy0hM/WJyPG0Ie35BEdKqUwruiAmHq7WnBdE
aRCO71aBjMGKBehHluV59paXzG1grPhCderQouayS8zULPM2rI48NPcFEdfrRc9V
6zabpKbPIywd/c62Ob9YTEhr1pfMddLAnNwLe09wOZHqZOdoQKpsaYGu0LwYrLZ4
SdeYrMK5Q+naDJ1Zp3OXdXSfXIlMd6N+x3MWD1Kqla71KpnQunZq7xymp+iWFAzt
UVUaCAER3uJa+wdbKh4pVmIGeyhu7X8fDYwT2smOn65moICTWIXOh/AE+oP3EJt/
05Q6gokpsss6Eond+7ZZ3Hyx9EClpvjUR6aBgAt3lqz/97O584P75Kei4+cyDY83
e6KhYonNmKn7LvDRsbu1bIU2RSM+zRtkasy8xW3EHJlmobLb+7D1JfeAxVwHSuRy
x0gDcH0lw/9SoBQZ0QnwCSG9tlHGAL+mBe318ZBhCx6Jm65StA5aTlgISywxJ9W3
mGh9sYz+W4HxiMo0vW3JGzCIbFnhPCAOLTh6zcCvF1vLOoCnQvKzyvTFRL34K25y
i+0igGI2kRwfAilsQ9IM9+arCThmV6Gm+AWMDo6OOIHw4B4DhUmLfNqlboPGwaN1
7NBFM7lQyFuYtaacS/aX3n1nmDYVlzE13okQ0b5YdcTBJ48yDh63Om8kFJMr5cOB
3qYXbmMg/lvvud7tT4DzZxc5KIcuLsH3MlNeiRxgC4UPnw6uXlbDbA9upT1VDbNS
bNVtFyAGmZzLkpqS5g4db5X0yK8WP4BBNF63VOuW0wnOeOj7uanyb0qbKXoIb/59
ou/ouDrEScBQqi8YBiv8BBxBfCbx+I3BH1/6OFPNeuhu8htaazc/tEN/gfSpU9Tb
IURIKp7aPG/akTCCGTuc0fAQ+UFJH+YmT0lTd7/U4YsUuZy2SiNiP4YFZxjo+TlP
zGSTc+pysHkJNwfKzfT6C73zGJGwlv4kh3dGRa7Hf2OFs1CBtn8Hsd6bA+jWx+sC
wthjRUglG9hNc2lZlMmJr0pCJTD78vMm6P35xdrwUiiq8BsUsaQx824GEx0ERZGx
tlEmE8NA8gnCDGAPWT2ZL3c38u3ZM0UkSfMX4zAuBgyhGimqU9gFYjdGexh1dDxv
R6vXp12Rj7Scp+ZkNZp3KFO1lP7XPfF97lvD2t6h3dnjJoq2FhFTDbibPyfrT7iq
xFMq0V0buEoFml5e7UxhYXUVWptefcX3Yfhh8NQUM3cX5sTuNj+Cmtbvh78RKlyq
+0tfvZ0IckNkTYHC8+m27JtyUaSFTBFeh7GIkvu+zqollYmQB3yOp8SxwhzxXOD0
MQqaHRfHBHCbGd56kNJk+wO7bb/y31bNPBnUfy1nn2lZo0hLrRvXrw8deHkd6IGj
qeqEz68l3r+5s6esBxhH1DeapUNfBzB3FsK5QKFxwmeY/eg+mpVcHW6IZKYndrUB
+DGUgMZicNf6mJmx/zo8b/FoplN/AqEnCknpsu3XFq5VwgF3Kv6vAF9vSF/zbsFo
E7iCcsROU/d2jWqhNnY3wPkE0hq58crUZ8eNvjVQYoB+YPyGecLAuVchdHJbzV9a
JZxYiRja50C1bbXozh6n/UNOU9H2uuZ69T0wUL1798Xan1V7tq7k3F9yjFrb7UVx
W1fh562LDd84mTwZQkb7QxlkIaO8zDJUOxLN+/Dp/8nEQEXHtsSfDYyt6Tofz3Kb
shd+UpAKy2i4P1TIp+MaqhSzJNmxIjk7GOicuUxCMCRFf79oq18CayXm0scEdcBm
1Tg32/yCOXZRteGOw8tvkhKQdfWIisuvpUcT/n8Y779zI4dTMQKJe7f1VlKEePrN
+jCBjDp/4mXMatp16PrrW8oYettqIyV+Ge/vPclQGEjvxi2jDQkdaAstvtnkFVZg
zGyzeEgI1gN66furhcBWIs3pBkzxr/lob6nu8gSC5TDLPY7pr5PflSOMrTUtswCL
uPpna9HEAu40SRh1N5zUMfidZQdEcqL7FMLC3SL39BuMtoI1D96W6VPZWp9uI3ig
WwOOPKUzWteXOBREbpvEW+Hiw56+UrRRvoQSkF2JLgdOJUYDIAB3t9RgHykMNw6z
MmxGXysFAcBv4HnuxxfIYTBDAb386JJ67tJOWtjl+j0xJkriAn0A5zXGhCMC4oQ7
3oKo/1AblJoaON7J4tR4O2AxcaYbAtDDdApO98wS1VypcluGM6FWNc5mpt7iKNY7
cNow+7/3RkV87O3q7nloxpAZWIFQqhSnZlEJUKXHtE9z5GV1wwOigyripw2SToYO
U3mGj5UXte3HZScrvSmmyM7pT4Eicfs+THVxwv17Fp0pKMkoBOZ/hfw+fpL/1SsP
eVGu5bdWrSsAsEzgsdSfPe48rXat51nn7ljaq3ZPrSpdyFwrc766zSDh9YiegOH1
eYmY06ItoyBJt0MVzYaVx1vOZu8z9VqWdQNf8TNeorWxOqaOLisDYEVr29PW3zoP
it+tCBJe510PriesB9UNy6EKwxE2eZfr3eKmqAMbLjXZxRyLGGXXejd1MZn6kX+t
sOeBLWtSLoASwepZNznQ9OupXwiIeqc05KW/UlcLW7yr1nO4XGIRT/5VMNaTc7Zb
QI5ccgA8eIvUTs+rQmwjR1JEt4dUVfBHLmQfTMuYR4ruYFnNoGh1gJanuEVFH3O6
JtT8cOHQlWBo7an6wU+bGEKo3HPEZDQVR8ROdbqQRLi6EwtCYQK12imN6Wq8oJpa
+R+8ANktaNQjbh6U1dnggQLtbs4Qq56/GBb1HS9p16nMqS8/Vf0otJwGTk28b36G
gFIntmDWuqFy5HfMPj9lT2jmbtnjWec7lA8PDflAy8F3bNf9plIvbiV8WCAE7Xnb
2myYUvLXuz5YVYIjYJuRhW5lh2zarNTMx8qEaC/sl821Mnxm054vDx7oIu/s8AoC
MQ/JAeKHSQgMC8Yom/bPPrmBPl2WKwPad6Ug1HYS7Nmp+Bsl0SxdJ7jMGdNfHLfD
RFWRXwjX+j0dQoMkn2GsQjcB07c/graPOpQGrNXUvqHwvqirOF6AdAliNV5wsvS1
iD90MTlWvflk/VUZIy0y+YdGvmh9Ch+Si47Jra6wAwbgS58YFitrIwr6JrGKTYg5
31CQkJSvME8e+yn8yhTvNAumvK/z9IbywrN6TiAhr3Za5PyFBOLlbkE4qfKJhGW9
PnU3zF3uswM1IbXBQ1SCJygCJAw5xWlvasc5TonUcIxKffZacvoyMesxgZ7R6rOQ
bkU10WVHXRTGB64lGiVDztt7Ly+cGhPpkYnicQyMwRUnoowaCCK1Z8xI48iz2kWC
7nQM0HI+6tPlu5121xS5Dcwh9XkvPIea3/1Yhr5Ked4w0JBlBIYDqhp7uG91nL5m
RDYnYsIY27eXdnBDAYiawUXI42EjrZWXtMHEC9iRBhBNGhJTWVmhVZO3QrrkCaYS
8m6t7uDyCQda7ZIYvFdZBIemo6UmgJ6oDZBZDEWQWMAA43NiznOmEKKPMGqM8w4o
uksUVq+vgvB1n8iyd0IJczecvwfljsrHfChc92WZPE/P99Y870TfGeSvqcv6FWcP
wnG0zm6Bf6MvZrjOH+2GSWb3Cf0QHG8k+1zRFT6gZGwDREgNYoM9hIFWj9ww18wN
PlAiFskUPU4EibMxHlNlhrvqVx6TCs1RRaBeZRK4qePOXqBA/tz7LVAFNYfFaBv6
LbZ6//Zk49xjqBm31u7imQU+6BzsFSYsfXdYpMFGsOMv81k5KuKp4QFNcZTFn95C
jXViZ615Ov+A4feE/ftqIgLaajZF5e4a1rPhsvWkZ+FYHbrlxao8hYDiXxLp7qnF
8bRU4b1zHrtzqXi9XhrB7/JhnawwlWx2cJCrihp+Ko8rOCpZ9q56HmTBlAJ35cDR
O2C2yq3VDCqoFCd+fECtnlegVrsTsTh0dBnn6MhZPbPy6xFKPrI0eYQDorg4OmNT
nsmIMcmtckHqXybdKYztw5pfsHapA9dAWtxQWNv2/Jx6y4QYjznxIipZRV7JtXRT
83GSZLBzBI5o73OXT4qNOZb43IGfJH10cvL3wZZb+bMaXLRK9/fiIl27UbFvxhSx
CF2f1h9cV2llzv5431hQJ00s1UNmmw7B4+7aW6YNsZKS6PXQcjDNtnFXSqTnNRDr
NEuAFEH+97+Jzan1zW4FXSTgfJIm102ZFqstE2bKHO4PTG0/ax00t2nlznvK5g4A
K9Agx5HhtcCfyvpq8wEbNO8Gr2VmFK4dMxYrs4C4/VbNRa3rANefsvbhiWiJghlK
hQ3xjTGLVQuuRbfXxfuQlYFLRod4Lj/Bkh8/rp4AQkGEEcViDHikSK6vq+JcEAuS
/SUcCIUa2xh8bkWHxOq9AYbHxrAd0gCEu1ac+Jvl0XPERedcYb9h9m9V/JEyqfS2
RfpOHirzkQ6KibVvoazyUvgLfuLsZHUnbBsZYxF9BEDhxUV5bVt4gbbZtQmabGYD
bOr0ob0OeNXJ4cU5RB5KZ7cmyC8c0TpGTby/KDz43dhrUc4qvMuezbUCtl4gcJbZ
bl0IsLJ5wkH+Z/jsZkys3zTtFA8QV457BBmIveHWkW8gjC3xDONwFZ5LjeibhT+X
/4ELdgIvrBCfvDuJ+Gm4nG52vxI/7aFzrUzM3TYxcGp9OeOMIaIGUPt4PXuRichf
BDWNhGZLs1S+/9rTvZicE/7cRYuMrPGnqfB5vfyZcopWD3Scu+mtQpnTqoxXrTpN
bkcqZYMaObwn6dQYydlNWt4YHe0Q9DxKF1psl3zmxTgSo1tZEiYDwuUPsE+IsGdC
B9O9LWmHVPBrUilT42n8IDyUoXBWW07CNDZiBOeEM3yFvSqbRvgXIx3Kwa7KOGcw
3kt+8bzYW1kIzlW5LZrTj4loJl+UofpBiMxsG80ZscxwVuSkkFkjsXI79FdHJEUq
gFdY2U5zjgzEpb92DNm6gllqR2LnYJa+jgi5qQAHG76he+pKJ3JTydXCI+FJDhll
GaVIIQ+DmT4yJmWEUbwOZWw6D+8MfWTNnbflXcBnphAofskkTxD2qTN+mY4mPmv1
BUIERemTuBPjQ9gCy+afTKZpO/Vdw0L8zCDPH3H4MmkCv62eg/cJWtKQt3OZwv48
MTmjRBwTlEzYO7Mnu/CzdMAcNo4bKNFNtRasJTmK8WM9VQVzDpUJfEM/VSpb0Nki
4+gR8oP1bM94HZUZxcCySkHjRbkVhIX4MKQkzBAeWCrASs3dr69pqSf26+uHNugA
lyLTmUlwp6eQHHs2S6SjiTL8HgBpjHLcuJ029eAcqwJx3k18hgsItfJOPD8hEvn1
Kx6hWOPF6IbFg6v0UrlU5nLDEWqnvaBO1deuA2qRr/LpgHTHthwlILcMAzKILsEz
jW8LY+fpZ7NpjAZjWVmJKuA4yDb7nWTKphDyPlw2Zi0h+It9utU3JmxxMEBMr6F9
J4/NEXw71+6E7SmJyHBB4oJ2TIMdJP1leR9nlqEVfZAThXlK8wqG6dKZJW04NzGH
RGUwIDB8+wPrLlaxTJoJuxJzLxW0f/MbmfGywc52TlR3Z3Om8mcc+/tiXFrYXBnw
ez1S5dftrxrp5bJGp/CUveuQilEpVg9r99uqv8ZEiD6FaA7C1eCA6NlG4G/QnFJv
BG4O0Q9qmxIT7ylqrnzvtTrNv4mUuni4r7kGG6mV6WIEEhj54NOgZEFUG3kBJIJx
8BVKsCiahbK2JbYX5nW1x4+DpYTZ/8yXVMstRMkTzXXYpbgUxHRrSV4wzYtytibH
I0qMZnYK1MlyJ/U3XVU8bD/mi+sQBliGYIvNTZHzoQEjK49RtMkmJ0TY+kXDVl9h
UvpLpE/KgwHu30mMb95VGBl8pMPBjJ4IbFV0R13K3Wg9Po6Qpzz5Xxb64z7B8NgQ
mb89eBtt2BJGypBT8LkMHk0WsuCF7si53AP1gDjNyRiPcguwAE2kvOf8zOGFLjGJ
iKSisZt/HLd07+N894WdNmjoJYTqzCxvmuyyA8+etiYJqfF46TN0xQRidYXURUHO
QvOiY4uhawnU5UYIkVMm+8RF070QIWV0UnRqFn2HB5oduke1A7q33gUikThQNmmS
v2H5DOEUmz0ohKpZW83By0QLShbshgh6L1N4xkEp0uzlPf/aH4xqm1fmgjEcCA0j
taLVtOH/Pq0xGMsBrOX7sje+reH4oQFEg22Rs0/BrStNcUukC3wo2ZZdyM74vgUm
v/11FNe+twpwPSAFmcV773K2PzewcERAlTdfdUfbEaYQaTq7yErhW1/tnUq+XmSu
SFqnCi1Fj+FfM7zEQ4cKc+54y9Xmu4Mn6pU361DRpn2Cv2yX+Xv+oiJdoQ4Eevm1
HJsrC7W14r2dfJsS9hBkiOxso4K4yvakH98uFKSff8n0iQ6E0TdK+pmOi+/B2D4t
MCIMU1q4cLB9+UgWAbKxtqvv+JaJDMeCC2EYMIGzZts2pxv6+kVu4LBfN00D0RNA
CBYx40GjWiqNsO8nB7uZTrfyjCf4KDw9sCMFv/Da5uyPCyjUdAfTe9PpLlVV9A2O
5cwKsiMCEY2g/owU7IoEQkEefvjbM4v2Tffkrts1uVzAvThJDjSL/3Z5CKYwD4cT
pk9UG4ut3N9TWiJsHNdC8qKV/n6y+d4T4r40x8eU4dI2ZtiKrLIt8ll52ezmAXp3
WUaJ7QtpejZSJin9wM5Dcv5X7/bzJgfzkI1gi48eA+AocYsZ9sWaJoWIM/yCJZxY
JLFcnskv2ib9H/ONKg71DCJ+fDhjlKYyO2QsSNQNNa9xpwnNeqvrW3sds03+aZq7
Ag67PW8kJR8ktiP1gGe3HS09zb7SY0JVO+aH0+4XHmibwdF3MQzciRUSETuJEdcF
o9GcrDPRKxSN4FZFD4nGRR71GaNN+wRhCjl1ijrByG82IiqWudsU6q4edivlpYIw
k9oZb8e+j4eQjFGGuo+VH5O4J284JviWeNdFgEpQ+2L10NgJgAy/lESaIS6AmIzO
GqXhI95ZlzZBplh1IkyCfulR9Sl/Z1cwlejVfkgEprIZSXPvWlYuumKDSnXwHPOz
zh7anwfjioLl3YmA1Ed12MKgEqKubiYsp4rt1GBVraUstpvIKgLnWnzggs/Uzc+r
zQTCxV+Qw+6JUC6TsgGJFqt4Er5rJvJBHbHqZOYBrA7GeJuj+2E+J5nBxfjPi6E6
hDOERa5foDRhep/O238I7lt/UpnUYDqqpkk337V6unAYBjoZaPUxtRcQAqLw3oVO
Je4Uc7u9mo4zKZ266Jb7qb/DvPJ8iH0NIwp0tMmYiIfBwXUFKVLuQZVkxPwQih6K
bptc6wu+HvB156cyIUhcntjaD8htsvGA46spH5iUAOC83ljHWWsR30qyg8IvRdXG
XUYvCDN3FyDUr3J7RxCkzkheH+aaRtca1CX3umYE0JjM/+igkIRviEm2HAQqCU+f
zCrEI7t1YXUZuKoGNwwdGwqaP7eBCl+rVCnf7N33KvP0D5qELdvKwRIqhXCPRafX
euRir3uQ6uv+ANFIG4QNP4TKgFzZicej1WeackWkO+VAw00PFsmqhTFuC2+R/Osz
Hg8O0HUQmu3U9UpK0YZFpde71OmZjiO2SIeyoSWFdj4P6OGRbg+5fkBlFUgD3ZBn
8smn0oyGqtWouqpdUfcOlsTvL/9DpgEPBgGf0wFFOi3nDvb9oHJlW+y9YARsQwqY
wcOzcmtPEkYyNLSjHRVEVfu9FVPUaw7Hwf5s33FJ//IBI7hxbWwu6NL/uRH8FH35
ASX0XnyyNvq6iQEriUGqmqIZ417CZh1g0TrKveNhW9oyZDmLj4ve2oNw2DX1LY6T
3VIht5ZC7Pg9t/j/SLcDU5Nzf2UvGApec+vmv/md2q3ITwX3D8N1F4xQAg4dZThx
jTQzJ3lVXY72UMPudEedHOdJbuh+Q5BKxIIYSjOLrtPSJae5k6JHPUPFjYgOEd/Z
OzKKzqOnTomrQ0ZYqg3F/64pxDo/+aCx8XJ9uApqCT5/6VTGsqliIGuq3KTNhP74
/UErLVB5IRct68LM4/qS7h8aeeJ93LN2j/NfWQTd6/0zoNywCnbDLXu6AI5+91N7
XOJ/3vrQ6lFZmE6FtJKPqxLTMMLLGe0m41lhrfpFj+XsIOdAKiNdh8+m8gfSGwfC
VuXTx4Gem5FeYYidcdl/kv/vSBONYdTmSTDWmcCcXvxljKItQ83ryrC+MZAYXaTt
T+0VL979efHHNevZnjnZ3Deg4spdeWoF4+Lq3Bwa6P8bv+5at8zj36lRahgfqDZ7
NV+7eCp1RdXM2+p7bceZwBelcVFiGKeVyI8zyojpzgYJ/dXumHrc33J0NWN46Rl0
UAyT15XxlOC/anRzcyYRtD08/aWCG46ggqn+eQIWqFFS5v4oQ3GBmeAWnR5YyxYo
KkqxnRNB3wu0CUk7J+yIa4yC3R9203E2j4sIbE1FKUCDgaDysMtZBadKv3gcI12c
QFlbyWXX0LWsgedVdd7O3Ss4S4cQipl0WqV4ND7pfUQbRfAANxwevPVMiKeiNKgX
cE+3kOJ1c06jPXvcmDQWz0OSsHhDgqjLMM6PoPtKV7+Uw/HHjzi8YWvdVC9c8wLt
dSJT1YF022kcivvGsZ05YG9rRO2/uklGlDSwUuDxT+JjzdMyAOgXn7F/0MExeOsl
dP5yIedpAtwfQXS/m5z3y+PG4ub8yKikVi4ILSOjo1muXOS3wgIzH7Yp65w5Rmqj
uPRe+uHShQM1Xn8CiOaStyqfKT3Ax8qJjX4Y+ls3I1Vpy2pKJDwPi+HoKYDX9JTB
ZK4GmxYNIeAnY9fj3lU3iDFyF14TxKdlw47tQickAQA7/1vriQhJ6p4kTRCcawJT
FwjTHJCeF7fTACSHVY/osOCAn4fZiA/WfwCGc0v5JZFTtedZVCq3sSwitxPimrsK
F6qOvncsGOUv7bMJ7obFkNJBw4bkNlKLXeulB+PVv5xKhKo3PL13awvQcvoOUVsv
cq1iq3lKlf4BfzyHSblV9GzJnF61a1IQn0qZORzN8U9ttDhSFsiwSzNABoM2sp6t
xnmVmlBZvc3oI4oMqWCUec55uCNjGXB0TNP1QDXRD09aQs/9ysoeWG+FsvqnNQz+
aJr2nBz/zxYVt2RfVXIltU0/rJxHWpZgOvMe3vLwOAuBiZ4RTOO47qeN9QAR7im+
IZY1w7OHbQziq3hOpYyv+AdSPw4pQmhk5XWFUYrAyilU+OLcUsS30icloRPU0ciq
ENa1WK4UBzijfQOlkIRR9D/YCCC3AEzePBOTEwejGKxBat8gbb8MjjRq3gp6Lg3U
EXmLknPYKPSvhhjRZv6gE5rOnz0EpZX+NrQbUfUqApFcMAOOjQ6LlI/PZyLTx0d+
OgSrT22B8BeQYkxq+Hq2+VxksaFLfrpcqbqSNxl6iieRnrfEidA5Apzi61/EI79s
rAz2b7vxDigxCxyP+RzNbshkTnFpgS4ZdvsrMVNOklTWvXZU622UbqCngp2XiYja
i9RLbYL2Obc2Bm1wNPAH806DUTOyBRUfkm1503RJv6AvPk+gtzBgVIz3vY/mczom
3jjINJ4prZpNyGMMsGGl43JiPRpQ4WFqYcVTUQ306jwYaLEk44rm2fbE4Ur/EZLu
wt0wfYsTXT2C7pfMQ8mN0whnRvkMXnBNY5oYYJ5fh2w5DRQNbEkShHJlhDFFXuWx
Nvs8RUXkBhIlpI0xpsn0Cu7pHxvqDCOr6O6Y/tq5+rCWKEhjWj1A2CAkywfK6eWH
lChvmtDTrxJ36g4QxMaEeG5V52WFTz9aIPKG/D3YqEjgZXjUo7RW5yW+AaNf0KSQ
8aOqEfUsFgHww1ow08RaObGPSRznDPVIphHkKxhs1mBPLHpAmxh5EI+mPF4N/iNh
mIFtijQEVleM/mvL8dcPySpxHKVdo9h4CU+UV12lJB0E7YvHXuvSmL2kMZa2oJE6
OceAsUkK+opFVMRap4UEb0TMHmuEom/I6UA9di+IpBZLLHyWKihQjJRxNMFKVtvw
6zGFFLgh+f+5EZ8lBDCz2DqJnnTnadsXuHAWbzNC19VdyP3RhcsfeboAB0AutQn+
xZ3WqoSHkia91YAls/HY1YSEX7SOozo47u/hXMOZ3V4bjwoeLWxhRCZvcwO67Bao
EWkG+2dyHl/gabWj1WdXqNWVopz/VcfUPHI6Q+zy81BOU7/pxgNPnFALufIhc8gB
doKSbX5jajEPAD086IHtq2m1d0nmB7Aa54jcx/bs/6T643gvutT3himj6XY8jIQx
D4N7OR2wuIqPJ/vu0h5oxY4dAJl6lvFHrfDUbcz4l7fs+fKE9hhhZOvxxpDmhhTg
qZ8to71MRxmf/rG8bB2n+7fT+y/LQz93eVb6S94Yb48C/dHXbp2GkAN42VsfBul9
QE6X5VWFTYCz1KzZjb5DrExvYSj67MDcZQg/SoPq5xLJc5onfEJQIxN5Juc4ZUXx
7n2Em4paS6mPuEWvQmpDD29UemtFXSDNsVM0Q9KsJfR7cHvZBwLGy5qSzhNjIvbI
s8YKzt3KZczqyI/SKPSpMUFUVfuUSAyzwFoWkvX0RcFDlh/R3r/EzcLkjF0hHyN0
UL6QCvdqJBG0y1dlG+2BpOD/4ROGk4HlL3nrfHlBY/Akvmjxw/z/uk+csPXdNxro
83p8Cc2Hf8gXYh6rFsgyjlTAPnheShjEo2of/Ks+UQfyvgBLFG0Qcas/SfAEDqKt
vIS6JxXsCIp8/Gz4pK2xGl+Rx81mxCK1iFYzNJXyZnTZoB+KY+hK4ELw7AC5dgyk
CTybxLShvyW5HfsZn59JsuAh+ScDiVT5EywiVHX4+3dz4maU8MyCZ5VgfShvBxga
y5JE2Mbifs9UhazabTcnZ5dLJBzRBtljphCCyXnGnZtnhFSkqsB2/RO+i+k4GHPO
Mx7x6UnHveGxz95SqvpkePLVPIRWtpr0cpugL+AZXN/It1WNAUqJfZRUzhAWxomJ
ihfo3b0GFtJSwR8dfSTBhk4w+KIhfMBRyePhrdwkLfvf6h1jgqxDAJdDeXwrKRdT
9lSQLvIzfd5SvciHwLHclntjDhZ+SCMymbOylJIfVA5fWcASk8K6Am+iagp8MOTv
gDhStnE0gLll3mwckJ6PdlkXb7E8suqBu1eZ/ut6Xu5b+mf5YA+sK4PxMEO2J82c
As9PytNLQMslI8jJjY5bSVioAVw2v0Ygvrf8NcUk45wid0mkWdYYM9q9rx3OFA2s
Q97Fq8RfIT+O/3KJQatI6HG+Z1fzuW5rIH//r6gP5z0faewxbabXkE5oeHFhX2GU
irvNojEQCHnnGFL585PRyOZUThjYzSCfdXhttKoDmaDl7I0TsydhmSqDX36BoXZE
lnQDnaSHzA+Xz9M1g50LvJYjrypW5yFd54kxFhe6AMTQxCAZ1vg0jh7FT8XJZpEu
j/g6R2i5jx+S7eoei6N2+54pbaJZ7MQByGJ5+P0VjESP0vOfeiXDj7fqpRLhWzIv
YRBBRYMLQwTA1SxXChl3t0HxlDFkzO3D7vJPF32E7iw+PqtNI+SxzApr+FLYgrV/
duuR40rBEbJKRa+RKkxOQZkZ+Y+4aSpY+rGBSc6sB4OCinggYCy+VBmZmXKRzuck
gM97wu+lE1vb+CSIv4iS+k04A5p8Y0BeN6Ktg8VVl5zdwcZ5VAg+yBBeRVcxe8FJ
vYqF1BRYnlpleY0lCqH+sJHgGznfCshuvA0z0LplXrKu0zREYTD/qDPBeQ9UD/7s
I6CXkRrdZ+aWyvVgdQAm4BIwE4McoBoAJBu1LWfBmVSaxBQIUsVPQFontt8Uz3su
ledK17Sw8UGWs52c3WcGFftUER9jwlJDS8ngx4pviaGNUpCil4GIkfKyHqcJFw70
t1wDbBLy/T1a0OGVkPFHylaPFGRkVJkFz3zJStJFdfgdVewDHDWZcbQoLcC4nwq7
/nrzef5wDMpnmVvytoR+mCqg3k34IUb0qaSqN/VqxiXqZkHLS+9XU0lBFajtAMUm
JhOdAdfDGfOJP7MTxHVnZbNh/9C3X9Hb0d5AGGG3kQEbL6pshAup+9ZYwG5UjAEY
b1xJVLLd7QFKkH+qC2niRj4g3CZ5QMVUfVmH8dvSsPqpyymHw5y6mVaKYpi1LQG2
G/CvzNznaberTz+9a4fjMnj/uQa7VX4UGTJozGJbhy2ulae2aH0E6aMZvHlQhtiu
94U3ip0hl/VVzLOvG9hAitofJ/CHU+GgdGj0hkDPPzQ1114Ph70QG20PvT8lRVmu
M6C7kAtCQAeSVSpJBxVghGE1y7AOwREsooGx0aBHs0xlebpISS3QNvD2+UWPlv7p
eUEq04uhYWvGcVj6av6uv3nqzcdi4Le5JsUdz+OKD8jqg65t3Y+QCq++0ZqpV76+
oFTsapdQXPaEPpClEoucSKlcHA5gSKzf06xlDPG5a59P3XP9Jea1ri+ihs0EVufd
ibR3iEtxz+pGt6ypVh9YDjKyt60n/RQCHY/X6sYTee2bzBNBoOMxk+5LExvfpHBR
dyrklOxMr6Hwiieg81E+l2sgksCMjfrjKum//DCPcIsQBhUyILGCP0eKFwt0kG76
9hkNbKHu49nOVI65j5DMXHGQqBtHzecbFZ7NbrGNJVEHTatQxja2V8nhmjiyp3Aw
KG+GjlTnYVUuJIJsMrGt1P4yzk7+tHJqOKP+OY87vbPd66fKY/GwBoT5xQZhkcmV
p6r56zqvpqxSgWiQbR4qarMu6/zegmimqqsMfdvFGUoSuECZNk2bKLnAcFToz9E8
XlwUKdsqK4HZpDvSMwQ+swiQvt4DNeJJQVpe99ZZb0I7iN9RuUl/l7Ck/ZHK5rms
TWEEfFtelLvq+jL1tmO5NiQKHDeom/+ihxrNhjn9jz1mplIl3dHy+3ZYyjPJM+0v
maRN/JDmjqJE6ZZum6oQ1fLNzg5k05cGDJ/kSqcfZb8QNt4oE/4XbpSZauTv35Uv
IXLTOrmpfW1SUtAXIPqoN2+Me1wbhRs84VBitdPfPJViO1mz+ZmhnnfbVOmzTimj
mLOqAjBKoI3oz3CMelhiaWHzLpCvgkt/Azf3Nmw/GVAWoMgxj2sjkMAilM0xd1QJ
FeVdXpz19c3BEmqeI0wSvR9eEligr/1g+eTrcn4+FwKr1XfB0Yqi2oQswT5JNVlx
PaAuwaUdfDw0UTiGwShjTRqaszM5COs8OjCRvEKeEGywHE/Mz+qSNb7Ldwrf+dXh
FaD8ooRCyBGUb5jVp/AtCdDireifHf8jrhlcS6J0ZA0ldDtnFTO43sViqAwDN6J7
e2sixphZ5rFQ8Z0i71PRizWyfbOHMYssBNfWaMjfM/jiG+SczV5A4m5mamV/epxe
7nmVT9kZLZgIF3wmnyOeW7b95OAjhFLY5TdrTHyOuuX+uyctFv+M5e+YkPbXA9iV
c+cpw4WniJKkaOkUW5WVkQr6PlIYVw+4CoM8eIb64A9g2CBQWpmkOhj2exqjt4j/
ZlW+sZ7kxHwm9T6AuDJRjMvBSxs2KPC6r1DnD2H+ID8gXzaLr5+yDjiPqoXUqgSk
7+Z1PH4YL80+e8JxA/dm32XYvm+ybPNbe0WvnZrJAlfbRdBmPIvKVR9ZKmT6CUw7
K65onBT9a0z3UUpJ4c6Hk3+lK2dkDtvf8wTzUtnfYLJ97CydUFMOy+zbe8EBVn1p
TWjNQS5Z8a8D/7+G0ZLh8pKWTV5sA5CbgKx4bA0ugyYl0oq7tHJ5fycqyuwC/ZW/
l4o3bTA2glwAeZ4zknJDp6aN/XodqLbpZGhGMi5YBTRF1y9k3JdP52NT1Y9WSvSH
COcpN7h6clBpyJY2Z5CFnHJv+RcOoMuWq7Owc4bKdd9dWCHp1jtyr93+ZFBtk6Ir
/acNk2cji6MoM/BafFqTVI/5UOHTqyzs/sk/g1ziY7zy1bnGei/kkZ944pYGrzTg
a40uLvGZmvzegn1nD5/56m+PQxhXmAloZBFS0Bm+WjEmOfA+6eYNRERCeS2zE+08
5N0BucKwAiQQSCO2dCjDbhh0Cm2M+wq+ilUdOGGsB5vbX1GUc+33YYzf5rFotqPo
/CnVxvvWY55xJrpG1dr3pkzhK3AEuJc3g2y/bY4ydMZ3R37HaFB2Bz7WJ9/9nPfP
pJv73BnHsfDaHESykJMI7PjgNHxVaKoWL45buLP05hh013VvlHqBCQJK4uKsVoc2
KsOYoXKQAcvABVhsCL6/Ru/lyrJJ5elgsYDDfDHGEYqxntcI1B8hF/0wb0WCeR68
jcJJemN8RINrNSfxDHRCLHevqA83rE1zUuQHO/0LVJpEWtE1BT34pND4nEziIPiN
gOheoNYno2yLNiE9E7qgCiDT1qIqNFg8JTNwK9KhdwAog2BCQpWsvDScZuCzD37D
saMf+6dDDscriZ24IpCKBXIvzqe6Xwg9/D4S1Oj8NA5q//sVczNWjnz/w1xhy12A
epXRaNtiYaU4kMgL066JrSokAxw3NsDiuKtiV42L7o+cfNg0ZhAfRXJ2wUFkAfFo
6rec4whXXlyLg0uNH8oms/DneTgKMe3RclX36mxr1FYTT5jiSBgUVuwn2jUPKy/e
wC34I/ly05rIH1VmZAZldw5qdiaYmf0m+ihtC4+foA4xYnZgrqg8XHbWBLz9lNhA
LXZGD3vEtE/doAnFE6I0qUuBU1MeUVS6ttVPYKte8koBCbRtkpf+LHynghoZx5kx
NImBI+mo0j9XZTdcbwfrKsY4gnRsvGNYph4VzPLuqx++24RtNmw+7IDisI7wb6+M
FjeYarQ9ljjxL8bHf5lK1wIyPkmUAKs2pkw8M9Bq8aHdI4btXn1Wro6fW1IS7b0g
kqFSS5UrI4IB2gdKzm2JfVQFni21H8oXOiu+JNpiD7bjsYK9yTXY3spFa5Sl9rim
lZd8eah45bADnred/UkPextlc1lGADfxlnJYtD47z74ZZmFZUKd3S2DGwewT9iHp
CkLyeFXGXwWhith+I3kirEujIYhb7xG5JQ0mh7SAjfJ6Uld98NBAINqo7H5SYbsV
yQyuCrHJvZEuqteL3BF6fyf+LPR02Dick3SP3fiFJAQ1OQuQPZfjCteUK61AoXuy
6RuTyKYZMQzT7RS6GOuc3bubsgNZZTdK8VaafOjTgeP9Y5BW69bPfpbMGWdsw0iT
CMDeoKq1gHnag4yAOIp0nRlbNRdthi92cxyBHS8I+uCatmk3TO3TG+Y2pikH7jPc
jMobemHjRDMfqWTihwy92bxH4n85Sqr4lJKR7AhCKz7awCH+Xno5EqqfdhGAuARP
04O9vcSy3IyA3W2tPWb4OMxt/+soyyqeE67J2G/8S+kLlZo1f7PLa10e/1nzVmAK
Bhab8Tpcqs3oFji6hSBzpNpyGVfsbQDaDll+BITXlJtzXycFBkUpF/cHBDr+bou9
r9rSXCeDINTYrSi/du5LjVHPRzl+Dc7V09C0WHBPHryIimn4THGG/ilvUOr5SHeJ
2THdNsVdU3eS17s3RR9U2nzo6qy4Gg0rMP24KG1kE+TFRYfp2AiB42cGSgmM/XLF
M3aEWZFzeSAow4/IGyMNhh6uktONrm0jly+/aQ1KjybaFnDpJ9ECaiFaItY9B1zT
HX/OUoDuHzOeVt9tpvwb0Gtf3G9VRwySTxR+Bvlm/XVRliuYDaeySmMCY7RIXe17
XCORMrqXiE8Pab+LpqFqI4EeayfuVe+28vo0nk/SKzASy7VZhiM6CZz/aP3QU94V
+80osYFeVQsIhChVmSEskyNs38NUQe16FYXgEP6IlfB7smXCSdsKbSUHKzlE+kir
zEb3AGOsP0+JXYJjycrkytBOLrPQoC8g+E1tFwcKye6ORbTu7z3o5AvdbcQhXI74
AzFfEeth2npXpLjfTTtNK/EMlpCF+0j3I6TQF/tM2QHQspV/7Mw4wi/q9x/2ufVN
5vosgJFqQzoU21bvhhdhC0Mt2eyZGKMC5Khd8hj6dw6UMqlKIw6lSwD8qSN3ufvX
p2Xg1QoSTFrCepHIQQZ6KiEmlNWKnwG5QcLv1iCz9Mbhgu36sQSF1tuUNcTMaMrs
Ty3QWu3siwYGT0gRimOD1oQGZdt31C9Z7gCevXxP+pFqW6R6iWxFmPC+stTNG5ce
uK+o6eWVMyaSRwZwhGe8UFf9NmxmxswiYEjkmD77UQuRQqpOK038u9hPBcG3L+ko
kefjIdHjxRR8qacwpSUjLumg0z4G9SVTqEcoR6BZkmbaeogo2mkdmlSX2ZAEC/XB
oedAsHE0YGxgcJ7TjbRt5nRLtnGF0DjImZBBGQc9uA7RT/MC2D8Qem6Vt/qqxw4x
gmD1QxLKurvuqm8+gpkSN5oJda+FDIQOo3fZQgdi4O+mju326WsGeruO4EZYKMF0
o9gHsDsigeGUaVl+WH/Kp/FRv+tJUdPvVtTtYC2Gk3qlLOGcG8fLYV9AYjlHChxu
wT1oB0CwUT2g+J26UbSNcvxePzkPNm0rIlcwfHfzhUk/dTGFWYbFr2+Jcwrxlcmx
Hz/ruzHxJceFJt2vPD/mbEpZ2InD1L1CfCdC/6S1YtPHjsMG/2xLy30kTGDinndf
8NIsmU8ZEDEXZ3TqHKIwR5zPCiz2gTUPJTOTtoQxiL/EKwF9xIP+XCTajkL/MQxg
tJwuBzbmj/CYtfi85eGDQK6FYnjBRFwMwj5XjPLRYHehYvacmiaNGclE5HyDRxeP
+xgVUj1CYWljQxHOLadvrcS2OOwAYTDPSEII9tvxFDSIohUqd/lWPMn/4sEwvEIp
j9RPjJRgO+rY09F/TpnZ/rcV9VdztVWwkPV1clXGn0hXeiPZFqc6rwuKh2fKNMm0
981Q//IXUKC914il1iZPSbt2KMmftnSrBlduBj/iBiXpg7i+AGdSQtrEyXCJdF7b
0rX2xH3N/caja3nZ4SeVvdrKmEuNK2Xv08t9OwTtGR0MEX+7jqC1yMfpRWRYz9NO
0Bpu4ariCLI7iLBbG5wRHbM/Sl5CxHfviNIV4R9SwfrtAERUIRjlYDJ6M02b2tV9
p+iauTGn0pVlhddUbSTpBioeC/u8t6Z8GDNc8e7mvC1ClX/43BhG5Ej3EHLh7RBD
EfoxnhBbRx3teFp/PxuGEYo8hBUwJHxvYifugvNc4xtlJfbIQbssTnsn706oOFfs
MFkxs2ymPJmUvOVhmPRDiqnAWUVAAXhJorSPkMvydkjU8tP1w+X/rFR45DuXwvqI
729B1UOoWv+ubCLydpOk/GN13zOfr2OZ5I5g7j/eu/0MXKBf7ZvqPik31dxeMY4V
kW3m5kgBwqqZ6G/zgOvuA4Yr4busqgb4sLB7JbSpzHIYqHQYtP8I7ATV5OvvY5Gu
ZR+bSCv8hF/UhE2YyADC8a4jSbWwF1aQhUFmdwKCBScC7B3OWdg1zeBfvTiZYcyz
SLwTi9O3JMtxdyNNW/UZqydMmrpmBLtjYP0Rzbp8QBVWWsaywVLVUOCbh9rAiZl0
CMr8d1gh5GfsS20FIJI9Bv2qTNGo2REO2e2rAhA4qAe4zBnXnu6DoKvGX1miFvAp
vjquxgdzvo9fhn1AlsT6nZiIHD55a9lfr053dHfFrm3eKfGvk/E4NT5bRB56PMzg
baV2caQI6De9YKYFslfLoGMJV4aRl0DgZL1Ad25Hd5kOAnEKw1HM1xnpOqUNHt+3
KzGSIbFK3QLTVrqZYtXbn15IWcQEv8jX2ehqmSzlfW4JGic9xEew1Iueu8oQI4jw
bkkFs01+81QH3ak60v3I32OGAMonZfo6pWbaewuVt5ajnPCbqUScMoUVReXw4ebB
driX64uvx8YMddD+CGD6t3b22fIIePRke7h9Zbsx4cToasP6q2DPbjP7DoYareF+
XekPR6VYR88h3M8r1+9f9TUqwVrAPIYIeUCBgJqVH7NeLp5h20d14bHAHTshCjXY
5Xk1LTOGBOh1FnaBUdnoNAUrzaCp/X/IwaNt7I8X5CEk+q8JVmhU/AHQH+vrGtJ/
JD3/T1JxfL2jI9n/A65mSr5N+cu3YwbiZmunuVXeD1lHHJ0wCLJjcmbUjNFzVYc7
+1usoMm027V4qa4P2qKL9zldgTz1D3JR4nLQbwayYUZkZOyBCsDSA5GRe1Pf1iIk
/fsbcb/npuWBsLiCwbEBqcz8CHPAaeToQ4Zxwn/PKOZjJe9B3pdh9sTWSq+k4A44
xs4dyrdwOw/+gb+eE656Qp3kUJzZxNVEbROKTrsWXCup8rrDOKWWKhsVpas6SIUp
grQDIlUyMjZs3vgo61ImzDf1V1UfnbZh6+Jiv8YvumVoN69VYl/9p5JqEPZpE/Av
tRCj4qRkUJgeIZLw4D9bgVb1vCjOPHc9hO5vxpM75m077wij07696et1m3zR08tk
tNOfb2WkFXw5lUs5fsKv2xg6wEMr47PN86KpThB/S4rM5zH0sm/q6TmViK2nm5Rz
q89OB7H3e+fRAja4zO6RrmllFhmOyLGq6Z0+n6oVEMeScaILIYe/52+LS0PirhOp
HOD5Vdf5dxCQYwTKnvCzWsA9zZUTpdWExS4+uANfFweG4URKEuGh4q8iHFsEoalA
apWaDwpB9uOpgALDc8wps/aj+ckCaMULxdt7xzAUUv5NhkXfOXahsYzVsTkOkB9K
mYnF/9ZeCE1XqmCFU7NIaVoprgclGTWhdRp42RiwsjAfeZrsyQ2VO2NCRHnZxdR6
PWqiwWAnD1U+jM40Fgxz6FUNsEHEEmrwTX2WJBNUPJ2ndGsjnsvseKEo1vU1LH/B
aZ1ad8tLtnNurREaqcjFmrhx/otm+s3zoAES9XgYDBM+kMczadcDUqbPw0fPnLpc
lG9V/yctOJArLTb0gepoptI9xrN8o8GllTUitsJxvlfC9P5Y853do/JeeX8JRi2P
UxoKLzGm1A9slPmuVIiSZv3XuVvfo3DoHUXyMkUg2PLhh8w7sj8OcYj4hX/GiZ9f
hxIOHGDvhJ6STx2KSMWxnM3RpoaNQe1rPq6Xkom1/8S3Q1eysm2pGGgJYMaZcoKc
9hs2Uk6FxhMDCvbZzQfyedd+TwExTo44l5cNH8Dt+8qsWGfxhCQbiUDcXDCdfbA2
C9gwIktZMgdOChLGdhjzNazuUTAKdPw4CCcROmz+oC0NEmTRxW3lihyTSV9aUu8z
vXywTU49cRnQYBaQO9qHiEMwuCAS0Mzpw5nwda/lzDPHuK+jlWlW7yk98jbbfu0z
JtJAIdW8pMs/303jZxeqPuoaxYaO1M0R1sJpxjXO6gWeuF4iKE8XHl5B56qz4qec
cAGKOF25FDzgEoLVc2G5yft6q/TrktkKp66LexxHb+U8xm6wdlssFE/NNZFcxVmd
9NFTfYrCyje9RHzXdnWjovInVcpYi8SWxkzpzn6w604pWvYDJpEgRpB1rhxpNh1F
QrgnGWrwondoHQDjCKpTGGRusq6baAKx4B0o/D/gSA1VH2CKFjVIL/4Y9BTNswZW
FBBoOv51NL3Tq7UL0l64dI8XzaQgoY2HE5k1mwEY7cICA5e4gDiaxDMb5PdRKmGg
0+NAJdh1uZ+dRqdlhMRqwRGf0F4UTXbh2xOb+tFD6zpKQF0KSUUliyxs4TshZ1Zu
NUC8zaq1XyfyjEZLYkZ3rdZWxYz3b2WyePgsuhxYCeeH8mSaWzqGMPtWX+kAw6ck
WYwr2Y2J2O0SBW4NMej4/qrIorzjCXSy41UJ4f/MugPEJiqDa0pjrxIxI09S54W3
CdVoJn2TyWzHzr0yPEAtilveggUzoEOMq+MYLBcuSWSID8z/TZYoH88F5Iylm0S7
ssXdXKt70gcnPUEKMrVtfw/k5JlBv9GJF8SkuPcukyIjcR2AX31rZkqgIeqTfo6Z
obBKGH+qPwS5JQiKYo++Vy//yzPakCeWd0OGjutCmFegL0o4BiC+6vp6GUaB4Pch
bW4tDmvOmCo35ptAp1AAA3k3ELxGWNR/KS8+IdrUHoNrpk63UkvwNXkOLDSs4v6f
r+/oppQLh9+Pya/HUu3MyCfdsD0ykBOcPmZ81as4L7fz06PEcwZrfoZRGPdypKgh
8VwrmK2jn20V6cQX8QTAL0qt+iqp3Y1C/dvsig+HJM98sz/eCk2AnuJQdNwa3wC6
CCyKMRNymTkGouGnZX5zwybRrzeGhPnVrPLedeIvrzwscxB/+p1nPbYf5Iapv8XG
Shf5PUzP83v6Z92gXtUZqN3W4JXORHLd3z+Mv72ao1sNO28EVUJRUA7UzSAviCfG
PTP7tElt2vKecIPkYL0VzY9lmJek8yxuSjzQnYVDzfVX3vI/bUqIQO4LqIUDBJbI
Lyw7uvB6qiqG3Bj5vHZzl36UO/7Aob+SxcJZo9FHHWKkqWuU1mhRo04exnmeFE/E
b2VQN2CtZR/WCnnnPsdwxUWfAgEFayFu2SHAEOU1eTAHSA+ZHwcBUcxq8WO4VvRt
1Wvl9lowHleAdHIiHA7IG43aWj1oHQfoZv0Js6b2oGelZP/xCtuab7WogSTpDaHV
zdQsS0EnQgwgSnzE2dS+vmTI4o6DQIvGS7Vl1wv77mK8ehNBxqCJyaiZspNaZ2bs
3oYa1PM5alOqZa6ITsk8m0aXw53zEf35J49VoQURivm1e/LJhFG53jZ/qVQeWHSn
Oh6dQOMPJK/k+0KYnVqNcnlwSR64JAqROy2MpufnHVX1Rk9D0qR3YRF2/qbTLo/H
6SPbsVioSLRXt8pyDVdFawDMCwfcsApsdjwmaZ4uDV5+sZYypWHAIPrNvzlT6XIN
HRLA+cq1NzJotiGX6CNpeutzKJ8DtuZtiL6CLsADFL0pUMm8fE3bR3T3UXXbRJ6P
qoXlz63O9QMCSAvCOWo7Utwv2AJK1ccpd1joCi7p9Pn4VLjPtKiGdh7GQ55gJpmI
WIBxas+3BII5sr3L+5k3MaZb18UWVYCvraw/yDymdnaNQk1a+UcYMG3qZtOD051L
5Gca6TViVdGfSU4CQxQ6dg3jwATB0lDMUL+Hr5kFdy118lmlTLSNoFC2ewyF36hO
rGnIZI2rwVqKghaSxHEFIC8PG3jeYL8I2mPnKSpNwouKyGMSlQPwKHcjnTJqP+1s
vuPRUqiIIR7s/jmlD14Csh7wt8Rgbf4ZTFjCdru9ZXg+5wcCtXekVnZL8omTpz3f
fam5AKfC3HUwaWqDoXIIskaWARTRTqogsGDxai4GxMhfuf8dlUQkc7Nfb0Nu+b/U
4Fljf7SC4+jYNQBctbnOpJZTMY3ApIBceRfJJzT3KfqnrnVEXJzHbLr/JuB75Sgk
JUWzatIWuaVuXAcM5IvzhSFOY7AkkmfpppQEqEYOYgZrg3hk0eVaf4C/WRnrIdqm
NPoSOc/DTCbl6wzukLRz7ee8f6s7DxLM+bp6FMNFXN/7+OY1oDPI6fzICGvX6nUu
ayonCoJCvYR0nwqLFIsnQx9W+RJpH9/5O3uiY67vv3LxaKy4DOpn2duyIXati0w3
9IdrZ8RluOrpR6D4DoY+Ve8w6iWlRX1yppPa68eK9COoX8dQ3Vpas16MIbrQgRkR
sP1b4xE6gYF5EVga4wjIBo2ZCpE5aAWyaccDfBMkJ2dEfJm5j/dnZk2HPIN8Z/eR
HGSof5dwkWhn+E/M3Xkd8ndqBNKfF1gZB9Wixj74nvkHewef2PJ/8x7kaCuUx3GW
ywE4uoFwgec6zhjb+sFdLdt4yfArfroEScHogp57i2vwNHOEVho7ffqJwU7NOMS5
VM+w0MPrlR2K6y2CGQGUVPkkX7oc+dQAz3nerWlY9ucVknzndBLCKKRoHu39qHFJ
2/t7SpJJ08Zr4aeaqiGfZqARSx1Z1QyjsXGKunY6StKKDbgzbtVNXayHt58TQnaw
Y6f8LnnuxRprIPnLgFUjYon1TdH4NMlI70chL+eI3vcXY36MqmqBUn0w6vX84Yr0
AhZHnmsM0fSTyTOKAidLyMhr/n9dr//Z3nCnHmYvGFUNmByVBjHKTHbGKOfOkcrQ
IfEY3HFYXAWGhz3L/f11FrMqDaDGcNCnu4NZOaSeigRg5u4JD9QZ/9WO8Qw3Ro/Y
eK74jpo97xbm2GZvHQJXBDekq6QAUPBn6mzy73t3yuf7fEtj5IkCe2xquv4j8JFI
l1rrVTgb56eHf4IQDmV8m/UbwbRa8H0Avh/zQ8iWQ8R6Hn9xg+5IQdzJIebgDXLM
akdrwCm/O8zWP6D28Y5GCiF4VQNyfptdPAA3xLZOoYk9ex5PNQdBncK2gnKbaE13
adRroEYC2YG6Nz2PGqqttQ==
`protect END_PROTECTED
