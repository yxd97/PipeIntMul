`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8NAZV/2TUOAp71AL4jWm8BiY+SZX1i2eiKmTip1PYoeSnnpC/65U7YadM1qll4Dn
rExo/HNDvHs/mCZon1sQU2fEk/dWlub6ogSRTbuTrkzpBBvdxtluRMLJrlJfYEiR
Ca3XkNzZvQI3uapK7xlbBjWUatq6iUl2RcO7SjXGQ849GOovVFz9YzR7kJBmJJKJ
KGRNCEf/ikXJQt30Yw9X0QoxXkgoIhX7hQFTf/XvEX5J2f5uWA6+BBSkJHREfU7W
5kwjl9P/avaM/xcm2Wxi4NUqmX6C3ZHYASgKqA/wghPNSKc21YIDECQHOuQJkLiY
xPUno83pnmIQvk07bBOFipX5CH20I210myLwYnJSGpQEIe5ONxQwMnsyz38EyRj6
DBDYKMdzuxx865Vyv72iZmQWremuxJ0Vtic90s1GIa8=
`protect END_PROTECTED
