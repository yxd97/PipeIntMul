`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y0zUtByOhYKatUvrxMKm6dhhiFt6yMMv5+sQyX9Ya2Rt7grx5tSK9Dua/XeijFoa
qOSp4PlY/dC1wWTeaDaxsmhy/iUeNf56JfayBc3BO8eHee2wMYUP6x/QqXCnHqEJ
DDqN2fbpvhty2qZ1aEOr6VVRCFsRuhYLE/1FkjfWH+PpMoXOtz3RfdSZkT2efwY7
pn4Kn9/lWTWVjba1qlchc/2/pnXl7v5upzHNz2qvxWpaL1aGRgXKBw9A2xml3nxM
oToG79CfPRceQapMg8wJSe6DYRiywIlzbsEI6g70Yz4PGj0Se2uaEVl5xsWhb7nJ
A5+nTu4lRsC0mSwx6ppIOK4LfPiPGYWXMVfAf8dA8TlzlAzmbcR4x7QXvJkMkD+n
0f8nXiuIX5lhoUPmttTHUFYdjsIv4eWMhQ+oQoBq45omHt4NABfKP1D7HKkJDuBi
vM2Gd9xMzU3XTk94uLS9Qq6+Lq3Spf54j9kgfC1clh3e76oWQGgYF+i9XckHpg5F
TvG79+EduzFXkmTf37YR4OltRf5KOMPcMnNDXd4BN0g6/ZTqwKyIzI+nu2ju1OtR
PG6CDj8CCCo4P6kKWUYH7Ng/Co6mQcoq6rIrcStpec7LMZ5XjEmFaa6orwBdNjvM
64LBY4zg57zUfF3eKrE+hnOqNjVno8HK5ixLds6FUKfL5l0b5h7GQtFhSA/E78wt
4swUiylfCvAbRKXQW+d+QJNyoYixVoL0AnlKnGRQbiiT7W5z2Bbj6SiJOKQ+EdXu
05bOBhy517GlvhwPSbxSWBhMdB2VWCHPONT5DxNX9QukOFA4rcwp8K56SgAEfFCe
5v1lMDlFgz3Wkjxjm3ct9S5uYjh5i9xbmfTiMKuHJGIQJf5M3RRowr3Xy320qoZb
zwLDmimxzK4NY5+Y38EVPRwEEPusZOfdwH8d+zL+7Do=
`protect END_PROTECTED
