`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMpbQHfN5aCIj8jjcdQ5pOJGu45HVYeLaed4Dk24FyY9ynrAh8KuN6MobX8Ml62u
x76sWy0u5NokzXElvy5HPIjxN2AOMAaDN+4WYz9g/plNrGT/zDxqn+zZvFTrt89X
2eMmAJHHjO7sKPgsHFOR6kg509Ewh9jRvgvFnNwgf87tVGwEZ6YKTFanN/TwtE5A
zOsDHPGpkXOJ2tqODRULTq4Mq0lDXn308iJ9SbK2dqXA7W4x2OLCZKwR0Ggpg2WN
7cjlUO04YAJQ7Yw81+fc+hDMlPSMDYPFSn2Yt7RvTtWCUe9bj07ZRi3WzHL+umvT
eTtUkILDRRmxrKuscZp68BzYZsoAkqnpAMFxYyiIf9jgvaa9URIzveIeOPKsiAXU
So8j6zxuz9PHMlluxlQ5SaMnf8lEQEyU3OR5rvxR3UKDT6mR4KLCDgi9t2jQPnCo
drMO1QziZYWSUr0GKTXYHDN2pmQubC++XRx9hUYesAvIcgvDhOKoXoQtVTgBYvE6
XQQ0DXrt0P8li8VM2/bLNSO5GPeShSpMUDaVgEELcKR0tzUx2D4RtIB0f2/bN0OE
`protect END_PROTECTED
