`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YukWB4LKlChxgz57JVV0iNeLPlXXVtx2NPoeK+MUOhZriCtUY4f5U/WpxxH4xwi
ulwdW6mrbxtOG+9f9sPHptLquUyNCd7qc22nGk6JgatsOgXURYBAuCTzoLb4n9jt
+9iUFJyEi4kjprrwCws4XLM1gmtdlMS0wrSOP0cpMJBHNg+OmvPILtJ/w85ezYh5
vHI6zFmBDCI2Ki29CpGpdYRgIcK+ty4jsGi27RMowsIjMtlhoTYRW+AGAeodFnqz
2x2eyK1Ku8QGHdR9zMeHRon7JlTdrw53o4W1etDvBewkZV+sxkZh+bTBKM+ZXInS
F+iSzfn/sBP9aCC9lnMeTS2hBrDb6/u7FEuAeLYL7qLeIgCTWeVKUhgVkVd8vDAk
keA+VuX/AWZaOGB1gqJqCz+SYDm0hpZxRLoa8bRUk6o=
`protect END_PROTECTED
