`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNmvUWwrsUluInyiKZ961icX+pf3P0cy+1ky14VUcIPhOBqd8HmZJOm4R5oWwQMy
/+t2vn7GwkYTM3Jz6f2PCqZ9SrR1eL7vmsxAGK6EkV02p6xEIXMN70zrS9+nSj8g
2bn6Ub5ExEH54E2CRgbgUQ/1+7WqXRKB5uJQAAV5OY4VTUp2be77hSgZyo6P7LHP
HGOx/BosV/GTTcxRQyr8BdTIIdkPS/VpVCBwPUbefRzhIlGoI2dZutsMfmtyAkAZ
saDap5ujYF+OFuRNIB2AGzF+FKKJUUwOaQUUPaWxl3I2rux2dLnyd0Fx0FVr0CAu
inRUaQiZw9SyOq8YMMaufxGFtBPfr2V/URkF5N6ZTpC/ZlDCdxjhBto6TCmekDkt
lptBBLLeiiWN9q/dACfhWQ==
`protect END_PROTECTED
