`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MHEZMBD/32/3Pp1LHmENEYg912SbIipn/zzxEgAf+5YVzQ3FidZYCwF/aZKCy0I
Z7yarlZzuzjHT1HDSo6IRbWJ8VpLTjUrxH2Q5JQBLCIAqlnjVX5/w4GdTQ8PaYRx
NFAWFqLy1iMQKBT/VAN561iqmwZuEZxnWIQuZnu4ArlJiJOxPCSiCeQ6cecEkU9g
E4gl6kgD8Dtqd0dcCpj/zGDBSCvnw9m/GZwWx/vu64b1cIAecegtFetBep5pqhIZ
vsmq/wmLAg60r5c2dhAYzF0xtOHf6xcKDAMUuZ0S9X8HX2A0riBp4hhrQaVHGcP9
GIo0tsCVusvQ7ZN8q9UKYldvWJkyzQ4xs791qL8lng//hWyn+WWejaBYz1ERJkp1
YhmUYy0KbvcsT09Eru10elwZpodLlbT9tmZ409rw0uHBZER0+lmDX1cVZ76CiHg4
xnekkv9QepdUBMvANpBKmjCv6mQ5DdsD6gLQhE9fuIjS/49ykNpvtLWco1HOV0hv
k8qBD6/SQsv00GxYSmtUOyKYjxf2eEsUmqk07zWkM2/Kj4BovK1OF8ASk2RzMdAi
EIQjw2M+NcEcflYpUbWSjl99L7NWfS4E+Z3nOiNdnV6Hfeps8z6aLMP+TezTGtb9
d6Aj1kYWNAAPoRCGQEAqSSUGe9onAXAAA6C58r7Whi80GTINnKnL7tmLjiQl3vSH
uD9+ucfKKHD4MHEUYMs5ovQd3R4jOuc29qCmOoy7RR/QukZEi/H5+KVWuKzBLp53
Q5nTNQ4n4Ungt7U+Mwl0Vp1iSzXULhur5qW/LE7JK7W/mZ7r34Fa83Bh8qoEruL1
ENSbKHim5qYPjDfOJwrH1/qBf0jgpE4mJqLH8hgFKgPbOO7TkQox0Y6IHJlQqL/W
CChFh8zTkJKdMujpTk1VT4MGYYeNepuZdoj2dSVlj7Sq23PZmqK7u9A5Y5QVg54E
+tFMfwNXt0PAMnX3q0MnBeyCIq04GAc1JE8HpUMDKobPFDVapDNZFLAYfrkXlOqL
OXgV8aX3eKiz6IdL7d/kwchHorSspUsauvYAm2e0kA39mUqaGvosLR1vzpjLbqKJ
pC80yD8DW0MOp3+Bhu/v/B7BkMTXZqBUvkuV/0NcNB2BRXzypMar9KoYctIxYWtS
N4O5NGmnJbeB5f1Zam3VrykZTliKvgwzyZEIabtBF6+NX3mHCUrJH3hSFEoHMSJ5
rRD3EQ2b2WgoMEpFavmETm0Eicy+yA1OHUrUIwS9UpPbS9V7uWJZr3kdDx+7IIUW
QKaGvqmNWDdICAvZRNliCuLWMx+iwnIEWAQk5zAq9P2gSNOTbdD5MjDD49TfNbW7
TXpSMGNR7ucwyzQLLoPuKKuIU54buotejlzR2EBcmiW/I8DR/C+IXl4rtitdSYIf
bf7x1prK5f7MVV2HcZ6pWAFsMLozkjI/NtMfxG4fmVkXXq0e6Gr/lw3Cu26SYQMc
zzQIXs/CAoxB/L/d6zuW1bxLNaiBcdl4Hh+Cb44MibUxFyOxhdnrnipCbHfMceFu
GpkHHeIETzv99AP0u2DKL5iXSrM3DotZQEx4Ntaw84oUd3HAiVTfFtLTeyhwZr9+
siY3vYUkBc45KB3ki9n3AjSurxgOM5pAKUmfnrzPoriSUqcDYvjkm+0x5Kq+exXC
1cJhSBzV0RnNSoURq7EMnjnydzJ2q00AT4hIzJm3C+JaDa42ojyhmsNzFOuo7FKW
sCfty1k8wGsTaG6RBLoQ+uROTeiJo+RXlupzvpqLKos=
`protect END_PROTECTED
