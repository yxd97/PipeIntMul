`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zhr5awfn6dJSUfZ9gSBwVy3k+1I09zptfUhVDiy4PCqhDOIX5+TqUzhWv5JZBg78
bB32fBDRVDGg1jABTVdKUxqL/fBgn/FVMZsXA1WIvLkZ7JjFEL6PKFIfYCn+yDXN
j69zoM4GTq+Q2h7pd3Y3wZRItlSAJu9sV5YzETknC8uz9bbQXcOhlo7Y5ynD4dVV
Lb2yHwbLY1Cjp+mrRIh5PRtjdzKq48k0yvwNoAKU14twY/mkt37VJzqRDIecgHUM
LcAc/gp68AfwoGxX/Q1IXgQeEKvUfx11UHzJZRafCP6S4nhwKjVnR9Y9ZHgGDtqa
de1tgMxRTR0xGo/PQnPRBaEL5olvSQupsWAFCjyW5S50AyBArnw4ypppVh6GEbKu
Au2kQnYYYdQg/Jyqy3cXYFesXAhk42y2N65Kou/ODc6WhC2slvidpR0/fbYDaKm0
BC6zF8VmFv6xWuCvEDm805FEUULOtE3nqHLZ5jB2x12LkLPre94SrnnFyAFKYcNW
nKMBBRlNEE9b4FIVaB7DBjHgADZ9SE1aynbE7KWlYmDxR/kqQrkAeF70Zm4/vQaK
wvNTZM+aTERJqKjz97H4VYvJsQEA173UOGqKJBRhXREG1AtM4z2AXh13sMW587qX
hPljtKQwOZ/MZr0WGquoAMj3E0JTe7vsUTjkLSUsNvUGElAf6h+so8PN863C4CEY
O0fbBthMZONXFo+EQvQKSX7FTAA9rIWpLGgYrcS7JTuyrN+6cHD7jhIPZ6YFchos
n0V3GBBWohpZqSRkAPc1JvNjmuFfwWeflOhYEnZlFghyhS+lH1tkSqk9rwm/D4Om
A2tmcNHWmWlTf0jjPgn33EpedapvMACNKlZ53+XWj/Yle48OK2g5PdgsOvHadJXJ
LJrNQC+5k5NG98KDlHAoWdHsU9Yy8XUxJfH4i4qC0vltJiZXBV40PAHrutE/qS4K
SmHUiY1R6wd4qc148TyMzc9YditBJ7dnPBkErJ/hTujsQX9T6Zot9GYi+aN+9pxr
oI7et392/U+Di6PSe7vIOoKb50BmdX/m7AWCy+S6sCGg/CtDPdZRDcss3CU9hAUU
+/cuIxYfBVrjGalYe5VQL8Fa0STLIaZ5foTvi/RSyivgDX2UFQocKKJZNzR8y2UY
8oLTkfGRvNOqYI+cd1ZuXJYd4i+42afg2g5ZiodGqD9uR4mU7yL+qAIlK1QiVKPI
8HkJPZWGB6eUeI3dnGTHyOIUQJsC95hCQUfObs2fGuYiqIMFK7Lbn6K2X4tIxh4D
iSEj+mjSUK+X7EdTIQCAO543kbMfvexyGbjg64ZTn21R+7LVtnotsAmiEOtUG/o3
ytyl3/N8bEFQ12Fn2cb03r0j7wENROi94l10ctViQjUQFefBOiV8Hek+vpa04d/i
TlKtFQci7J8fUWQOR7NOE1Jk3wWoSHvLY7JjUNMcZo5keL8JhFD5v6+kETZGZyWc
gcbx+C0B/hATfYq7Btu7XJ2OyPeSDuMZBWsUFKvu9sHpyWVWnBRum9gdxCR6nuHP
lye7UfEgTw876iiKBfFgDEa2DH+TGBanxHsuShgVP1+lgZFC++SPnZawXxY6zoo+
xBQNvQsF3G6jrbcchR+0Wj4dfasvBnbjWxHhXoUE6Fvft/7gy7S+eK/9nosejXfg
6zhLQc9ozODrOACI1YHAKD6r5I77Ky9ksuKXALlgNVRNGoDw6POly3K55VAxvvcd
U8QwUxVPRkVRjlUS4LWHlL021fuSRme9ECWpmlPuwhmxjfw9wdVHqpo3Pb1/aHMD
QQhkvf+VWi4ZOfEGcmny0bRySN25JXvu7jtJgFqGNlYofK+Vy+ld+vqkNMn50xcm
FJzu0vp1GiVlWlD3MiNmLNXoQqAymWAOWhIH2J5Xb29r89xP1P5J7AIVHEAzyy+S
o85BVUd4QVhAr66osSdsie8mUGVWGqRpiDpyOSEFiQ8doUVD7bzjfvExOv+xAnRL
29UL/D3v/6N48rwNAkrgaVf5D2z+BBLDWewGMEujzM/lfhJ8RhvRkyU+roJwZWKY
txl2nVlV9vO0wSLIUbmKUMQ4ZhfLbhXQbbic3BG2fni34I/81y7uGxpERF8/8jQf
/Pr5kA9eORZWKYJlEssmrumTsbAlFRi4NDlVjwiuspC6niDoRRmN0vmxBsNyxvTe
P6TBFVrPLpnY3prTD2fEvINitNmt6BAno/FyeKJqddiLkdiNO/wK9akeB4UcD43d
XczQPPJpEageTdcohnm/H8wuCsIfipzmmjVgwxZjhPQ/UqPGAv7ZBGlXkAEpmqj6
oghkF7ldMU8eNLIoYtHVodoPC5N8LMAHwQ4r4Er7y0PdODe7y3wPoz4ZChgNXwGQ
45ph1biR7tzAO8w2QnowGeuVnN+2Ko191rVTnQVH3MAZiQwLxQguNni/7lpLSYL7
++pJ8toUERkevdxXTj8+JR6O2rQq27wguvSQKjBE2Xqz01pB8J9P3pSgfNGK05Ex
F7Oxh2RcTAVNCTmZsfqyCUxRwfj/Kk/Tqmjb+PhtMhoNq6q+QWAKmsZ0nyUfNasQ
Jbfao8zcsRVH4NbFBLwDi+ltJVrtnPPxPiYz5nVMHUWzsQVMqMNyJMXAxxda2TZ6
+aSjkuRa4HFATi0lGFQ9w4YrTt9vvANL25sGmj9ZF3bFseWHosH54ddrNV5DvWUo
fo9Q9O4el4Jmgh/dac0jZyAgDpBwSnsdBUgaP0RkDk9NNd0bB5CnaQETMUs5DNBk
MCArPnMagaS2lAPS29HbQw==
`protect END_PROTECTED
