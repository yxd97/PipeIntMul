`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqbZ8mwwaYkstq2jQoprVheDRO4UvogY1QETnk8oTQnlZeYU5xLTfI9UpABkkwcv
NApklbmsrmxdtJSbiyRAWyI96hsktVvGimPN+CIkEFmmP+Z5WPHGRZKjjzrD0go3
EK6MnkDtRp70AiYq2dIvBqKZ0OeAOBkIbopvSiQpqc/xxfamT7us9hiOw/PUErbO
BO3l82tkOdWjWsIbWy6scawbtE9/6y2jwPN2oZZOS9PfBLG/Xf5MImlxDcY8dhWJ
y73J2OKQUMaPV11iHJBZTHQAe0LnTZ/Kpzt356QuB62ogqJ63Ucmvfxq74hPD7L3
8QQhHCsIUJafY293S3iXsxlN5qNNyGk0+nHJOQQCfx4x9ANOKrGOEB7NaDlaFSej
`protect END_PROTECTED
