`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jrUmFfWrKfh3ghxmtRolRq7jYlOlKEjsMZwQBAHU+JReJseQ92xklXWKyoIjJS3j
XWMS9UfoOoM2HLAkmpXht46gr4mbQD8YtXFPZnByVB/O1Bw0tanwdbPA7gEZJOc7
wmTJZBjj3x8uFfN9/LkGFaiF9kc89gUiuXrwdTO8bOrhcqCVCW9a2QwU32EZinmX
PA/Q48oM8r98JC7gnVvrCCRKqOHnzDsTsytd88EcHwvmrkFJ/q+RALJ3ZfLJGuiE
WuOJjmDbXTuyEw3tOuptDsw/FlnwST+txsN0KDb2X/E=
`protect END_PROTECTED
