`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z0kHedsvBHhpF4LPIma1HWU9qHJ3DX2c/ePNQGeC7Fa8jfHqiOK+SXggwg//hKHw
bQLHAkVcxIxGQ/1D/jFoERZ3e3pTOAV2sEvXNmwPtHEyVKxbtJtPZxiIdQR50WeA
JLgigPVLw0YZwp1QC+xGeZ+PvUexJri5ulszAso0irrZUoJbSwdUch+UxStj4bki
FI22YXDWj79waP+xjNuKzMQwUdjVYIn5v1haIfOLC8th0cM/bTmw5kQFtlM8FvgC
kmoIa0M8YCFHZ+qzO5DMe4J6HFbPUr9o8T75dpMmzbOuHCHWeUDjxEwXBrQJlQTS
ux7vQjqBFYR6ChwJnPrwqqNvnB3H+yQ/kITWi4IEuPGVFhtU9xoDECaGYDm+Wvlb
Ins3NOkpfIdYFYeXcF6OuSyeIpfKr/VyOd522lG6uSA=
`protect END_PROTECTED
