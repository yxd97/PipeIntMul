`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9ELiEypDZd4SiuJ49mz6iOMqgqNUiVJ88hDD+n9VWc376Tpsqo7mWEuDKKslYtA
GkSpE5uY1WtL00NSznZINjpPPs5uvSOYvkv+aE4bNP2zO3O0DvBLLEAiFJuR3BPa
1/Pt5+XhONXja9G57OyCQChg+r5vq2FvbLcNCJZ6F1gAN5q7NChBTFygftqXwLcn
u+l5L1pY85EkmKBE8MXGw2Slq3SToABgNtL9hVJUM6GuNOZt323IKya2pLE8iGuk
Fd4rMNju0myqBkD7AOr7YNtsUEdDOq13ragy889GjCaBxlUk7glY+2Qm+wyVxryJ
5YuY1rCEPfESl7wWzpoy9ueD8+IXrWLofXf8CEmV7UBGoILaQIkcnPIisWmc4qii
sblKl9q9CcedWiQY9zfECscK/a5WLlKIZljEXzBNTcFApOmxUQBd36RSLKa9Qk6D
O9PRJOm2Zv7iZRjIRoJJqAsmjP14PoxwdWEMDDgFSHw=
`protect END_PROTECTED
