`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9AJEjepHZhaWQ6p6bNmkepHRSMaVrSU3rAhXRxUY4XZpQtC2HBOdCtjG6EYOogK
JEALVA9Y11U0qfGkK0GuE0fLrqM8VXjbAENHZXQJM4MvORjMwip6LtSxHZoz+Hrv
Zy0opeXCuOB2LAYbYArty0A5IAqtQnyk/m6rNdmkoHuPJbuxRDwpcAhx1erVwl5b
li1OOdhss2sL8AtosbOJgz+sR/rsw2qeGIZFod2oOtfr/3cz688lo65LIAWeROli
0Snpd3JIcF4szujKUkYSDAwbxJgyWfgu7b91MKsZ4Ec3yfK+mER2D9OoFi79HOLi
pcjwAdspmielc+P5zcRkWN6FMRje1BsgBUawrjoh38KNmfRO5MB6A6NGU0XnEdSd
`protect END_PROTECTED
