`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sBzbze9k0hVaqNDMKkVAa1dMhDJ2bg7qjPaCEpTfNKr5ZeOBnzcYn0ETMy4DMqxR
3LeBEY2mM5f6LSwthEtFvVjvsTbrkyg6oHIJJfVcURrPFqck35hwshVbmUwbN9yt
ge8unjsN05hDuN2Uy4TKojrmvds4rsnMFvA5GzjwD4oewAE9jDznL/e6nxDjVYc8
fI8Wm9bZxp9q62uvSNy497juKCVVT6Fe1n/HJBWA2h468D0aWDkX6bxxXv2j9ZWs
nNvSq1RveriINYtVAjnlk8DW9jXg5OQLzbsbSDnQZJro2hbyIMjVNf5rHrQXN2Lb
Fc9bxPyNtF+vtZqeX7YuU6JvhS6nLZVORbKpneSY/riY5WAHtXUHCsXipPPBHyYg
iWjulMN4VN2WwgJv09hfNXlyRt1iEaEyaz149rWIDfkQwzqbSje3AJSMeMvkmc8u
XBCDg8rD/OiJKxXFlh2AvjJBtBAF+6ou4TvJW/7QSLrdxGklDIlwRwfYbP3PVuij
VHIHNaHCBhM4kFjhUObijOEIwLhLILoos732kYrPHeFZwoFUB3lrSXyMpLsMnvv0
`protect END_PROTECTED
