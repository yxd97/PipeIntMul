`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHhFEIxTyFRiLyD98boXc/9K0p0WySwvDWRtQ8znEm7AP4yKtdaLg1//JdEApNC8
X1QH2gJ3rB5rxOsZx/2tsctleWIUXiHRUJrBhY4hj5D+ZX7m7VXOO2GGVDEhNAX9
pXmQGDNQp4fqHhAwkvKWfR0K7l0Yg2/77NPNN1EoWn5xWUdoR2ILF+HlPozumiMf
5dD/eZbIVEspMT+99kERYzaT8WpSdNn2QjCZSUf9fzwO7E29dnzb3JfxhyVT7eTl
25oJ6S/5LfMVkiRpXi8aJRjEZDa4V2ZJI2LDw5H3WL04Crvt+LZ08fPsttFXcrNs
3UdkhtlFe89sgw3y06+vM4gaPkSR1oypqllV/TEja2gp1Ph9pf/2dnaEeMMy6YAr
HYje4ZftWE79k4M+HYVnEo6MouLLPDVV2DPnWdWpzMFICKUSZ168VaaNWoov2Xjs
YmHXijcGL9dPZc52JkxLEMZqIN1Km/QiYugLd17OfCecYXkdcUWZ4Hr85nvKh25I
lYv1zyQBaX8pXK/vfaq5XyAE5YXS5qz7wb3Mj5OjvcgAyfPCOsUV66kLFEjXqs5f
mhflxutBpaflDKk7jT9Ugi6sA8iWOF7l7/9tlIvy+lU=
`protect END_PROTECTED
