`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MotjZL8j0Msz3N0a+VgUsXyqs+UQpZ95OqSZopKgpApZVtq95Xfwfl7j6VWoWR2z
f+QWUwLbTny4N1m2bmtWFaGYanJlDoCsehN2rFn5HIYNfk5W79kge6oQ98wnTdvA
LZARYDpW9z/jfIPEqB2kFNz7Tv68iWAtvU8fWjfbNGX+SbMVtHlHGzEPFtgTwAOp
AyuTHOp2LcOy4YwFgUZi5ssHq2pYvcoZJ8o7C7rUJ4HR4JsUYjGFGoSPSPGHIPr+
RfKogX8sw6ZVrBI0lpZyJy0uZxjcByqL6hLcthB5m/xWBqHnq1E3O+iVaNOHt2o+
7KMNN6c0GFdiDVBeeFugm9adJ2gZe5gc4MlpRT7i/SIDDroazMNHp9Pa0xkaoGIV
h76HsX6ZKG5JgEHcOZyH3q7lbn1a5SRNsp8BwpANGCEEU1AMb0RX5ZB2SDs9cRVs
vuhaLN0mKTmjdzja6llWUzSc5qeQM+A/QzeLDXRY8vi/fx06NmXpC7bOgC1Mu4MD
`protect END_PROTECTED
