`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHXj1LFon2I8rb16GDKapIYgzB8fzPlfxwu+7fng+ZFLdgm+cq0kqCIBsplTMAOT
mOt9hAVfprk94rlX5jJzGsvP9TeLnYkK21G9r6LZIqkRJj/MBlRf3+INHW76RJqT
zd3wFSzRk3GUU+jiCmczya/9eHc8W0ZdtHl7RG1aXqTb2SieS043fj3cvor9HYIH
3ueWdox+gjz7VUYcPbSLRs6e1I3ZoHuSRsvCVUZJs8QCFmZ8lIesoUmJ1vsdr+G6
ZBGWk7RPl67tXP0UFae29kUkyYpZE1EwYWE5RDMKG4Ta1Fb+JjDbgsZoIJiEnKO+
3oX2W3ocewVdTrJkzU9unnJ3T1ldABR9b+JhUK+oV0B3qS+I9q9BMUidwawolca7
4XBTyJU2yI1ghUoouO8El0RkjTADyio1HwsXDhOgimoFlut0fw7vPe6mvCbg5TMq
9LSH0VUDCuZcPiwGb+/1191mxAtTnN8Ma1RUMzoin3KXP5F3KfMK+ME+1UMQSZ7A
tOWsDLLyoWJwxblzqs8Mxcgf6areMLCHlV4vgJrIm6EYTPYzlSBOJB2u78qgb33+
unM91hnp71ooDGRLoRUJtUOfD5nnM6dqg8DVHybbhNILeYoAdoXiR79pPLVh1DM+
ccCvTRvKJ6cRaN2hvcOwwdCEFaYD7w5VGj6RWS5g9r6aJ7AL676Va+TKFlV1nlCQ
fNieUMy6nIWxdZR2/EilVFecywmx+e2grhhh4SSAAecCduRo8cn+hS2uQiwsu675
DQSojBGZzgcn51qLWOf9/uh7z1vPRv+NqdJz5f64AGMBM4fGPmNBbyYRLp8j9iOg
uzYKsilvgoQuY1J3kDoYow==
`protect END_PROTECTED
