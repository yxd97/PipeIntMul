`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UUXGdS782eYGtl5CJ0UZ/9WgdG87XMt65U9TiCC/+sJl4b1CeTirDmPXfPD7AVun
OAHGtrbCQL7MZjkBcuUqhiJZw/cmRo1XxGdpiP8HTB5xto5zml8Z4bQDPoUHWwix
twXDi+t/ZnsckAup2CGzJBILFp3xFWwkfbNK4dlEh+fgFnjciOl46sGmRggC09/q
i/dYCbJbDNo7MOWKcjBs9FbJ68g9Dz4S1Zeo0i/TaI6tV2ptoYk/J+eMpW4ahMXm
jRJjO1lzeCYRioEdmjnKmfs5NujEFqSctKLgn24pANqVipCMDDaE5LOQ4tgKg+Ms
U47I4RYC8ZkWpX5XsObFV2qXkOYBtTmIDXiv5YJlUJCoG4iuq31vTKUklusWVkJX
z2iAgQBmRB9z+eVMB2PQOrDCIoMgKbbHfD6FsCO2HaFwcAWbOvC5Ek3TN7KlqUeS
EdbNERa7qcCzB9jkHU60BAEU0Kljhh9jSvmgpNGrWLXPQIArEhYrVJ8YeXGgAC2H
JZGmAAMwyb3H0DeH/wUabRNVclSHis//X7qz+s1lusnODFY+RdrkFGXsTtPifi0I
J+unxLLPbsIIYtk55rL5FA==
`protect END_PROTECTED
