`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8FzdbRWn9lgnFOmNRDQu0UdYqdI9vY4ob5F+HecncuHlHBz3KAWX327MWfkFT676
sUvysKkPIPdIZH3BljohRcLcVdetrh8hJvDI04zP/S/DBkDHm3dY8/sVFc8zkQQU
LCAW6LzxtnhWb63mnbSRx276/ysRpseXoE8zpeW/prag52dFpIdtufhvsbfvCSQw
zOWsB5IFqiRUpjg58s7RJQzX5IrY8dV/D8/wP/BpFaJFn0yJy/D5/1QTSzBDZz8k
M1m/aOvWvRAPueVfyu4dG954hkur5keiO1SgbfOwdvbTGipE3xo6o5UIcmf3x0/S
glDo9Pl00jEaLWyPrY5b8+6boq2GyIa5E7za8oyr2niyl/YbW+hAD19GNDo5DolL
OGiql5dpN3RqN6ApwjRmC241QfT3REmrlhZ1lm/vN7AxG1UzPDGyDfl1utB52Dkn
PJ9cxHuFOmDBeGUqIIRqy2PEw9gwx0aUkFbQSs6ko2EP62Lk9j4SnizsfqzN/rov
a4T7Nd8Prc+1ujdVPCztpnTb+C1jSqrN4llWbtKAkzM97I8pUqm5UzKykWUS2eOQ
`protect END_PROTECTED
