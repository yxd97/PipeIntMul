`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RgkdcRYUteKjts8u41gbionxZAThIgj0s6+ikE7EToN+8IKkOot7nS59VXCGMiN+
ON/nJGnMy38eatim7y7vptXB95xBW5vx4Uy19sI8q440QlRmBrHyBH3akGXi61ag
bVC09HFShJQU/S5Ra2uuNmOxIW2Lc/cx0sm9X87lwH7ntD1nH0ov03T1FnpM7gnG
+y27vTlv9mb5nCdZ6qchHUTinS+Ov+sPaTVmVf6EoxhMgbW4iHygIJHRuZwcTNtD
qKyC+PtGqLBHD6f5ZQUIIqG0xJ240kCeUKva2dTflFB690j2Fi6ygNAfaGfokFTS
7EdR78U34upeBE8rx59g3S9r6wgdInEuIphZOMa6GCNYqdt6t8Tv17JW99TYj5vm
Gt2kNVr4iNGw5D8J/ObGmE6MA99jAH9cArpxR3mnbrX80PoAZJ8Qnsod6+xaxFJG
Gs3ruZx/DwvxYN8J2odguUiVW+uY4hv9t36EfQASeSXeN25wpsIF8ajKocGiOrvu
dDD0drlDhwI2SVsW1E2x/pEV7+ZzOLq3Ue9LVLcsSon3cuWtARVRhM3XhGMO29SF
Q2pTPzCd9WfiDzoAEbkwqrAxqxFsazob8jq/YGfK/sVSXilrvrucktiDGMMe+dBa
64gnMJRBR2V2LqY97g+jCKrAhRvaXU55buHFf7zHNrPhWCpLdXufWNL+WavxHgzu
JYXwuk0LFqdYrT8+hqBdq2x1CAlGP3gbWDzjKTKlLEeW2FXQQRAiPnkqhp3BXbNf
qBc4lqRa5d0s+5JZPQ2E/t2R6bjVZJ085q2hicV7w2kegENTQsGSsfxC6CkCtwti
HN3gVg6zaZoo4sEypc3Dj46hKB/76465+Ce9Ry9eVJnF1SvUa8mQ50RXehiB7Az8
SdEJiiEyUnh1L0+d61rApYL8xUm0nWWeFyy1Jg6MIZNeA9N73v53bZhgKVMJmE0K
PJc0NZAmOGGhDiW3HwVu5MhrUJF6DrzCnvdtPg7rQf2rtGRw9ecLkW31LJXCQm5G
YIyevlgtosVi+ayjgmyaHTgtnKptcWFd+Sr4QLZifua3BFDJyte+PU6zRaQAPB8g
cgkOvgaKgxDy7chr6nnpRBhSZHVWzu3kYEXy/jrpmEGWMA0axmbwS8PwnH39TCjV
rsHHLqUOzqSfqp6oDIoFQTR4kwxgwLiQMnsahy2DIMyFdqtXrv7k1lfZo7Cq8AJ2
vPKredlyRzI0sWEUwZAyPuVRolBIhouBFbFzCNU+zFM=
`protect END_PROTECTED
