`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NUa0Zrk1uZewYEoF9mo2o8a3MDuH3hjAaKXP5FcGBDWOHkw+e/Gp2ME/y0Uj/0Df
tGl37pgvKX0f1WpDNXMJQE8lpsTJzh6dUveGBDXZwVjQuWcaFJMeMZJQOox8qfb4
dZLF5JsHJg2CC6ghoFZKP8FiEmXLR/vEFJy8xUpou1BY2MbnLvRk3masmffhGEHB
RlyBOU7QMrbkFLvdeQ+gwH48s1DZPdL8qfXha6JbLi0g0xIciZaiUqt8msDB+CPa
204q8Wd471GfL1a81CWqOWG77qn7Ys4LxM+ymgy98nU37TwpRm4/06t9j5eCrUAw
K39nL5/YnTp3bGWLuGd5J6d9nIjDk1p9B0o4hj58wZY549CQ3Sg71jj3XqyqVh7n
K6l/a/NCQXRRn0a6s+TvF5f6NQqKrU/tYaebLgr1KLr6EEZSg6IYq6ouGbRgwXfw
`protect END_PROTECTED
