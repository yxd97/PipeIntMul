`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Im2iuyqE7i7zUzbB7Dg/1sQzXJRCDwZG7tRQmZqvZ3gQzODVavDYC4hYs3rbILXd
y7BbxkvbKlWkYxZN3S06UoEIKcGX0/zGEPOpDKq4GBIF7c8pCXioG/stWie6awn6
FV/3cUIhzCDtPOLh0lK8a1ko5wb7B1Jviy1S8CUC2ui8XYW7ysWYJ0gDHeWSxP1X
S95jp3e6f5mBNRCNNjHoP05DqGgPgDwkjqU7HbslbjlTicB9hhazIThoC16Gyu3o
bUoKyKF+SZa6hTLHZvnLtbZr5m8S1bM/zHTkxFtUa30DHu/Q+FvRDokBZmTfqeCc
PJsLxjgW+Ck+ovX/FR4BjOov1c2135FOeJc+Jgyxte1m1hD6Kl63rI0FGH1ra+Fw
9JrEoxYmv/w2YRIfmOZ/Xd7Itl8GuXwn9iHMu/WARbA3jkP7Mqxr0v4tQCHW7Oyw
`protect END_PROTECTED
