`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ptRSbJQQmh70ugVo2AT/wUPuRVymJ6UdknNFtMrvcPTBXa3U8qe6feEZ9zSXNpHr
rMsLGGttZe21EJjrXrCR0EXTCcV2TWOAihMBz7MC4m2UEl1wTMTxSVstglFkxuhu
1JJ45Tx3jSNlH1wQUeHSIv8lL5mvSlVHSUQhuUu9X4HG90aFeuRNIE+P74kdHDla
hZ4FZGBEdl/bzf0oHuCShl9H5NzTK9C35UArHVsaBUL1g7oTx7Y4ch7yxPzd7P1K
9uvuUydHlv2Pho11Qhm2iQ3flMj4ak1/BaDSTwwL7pO8OWd6oG/+x+bA1LwHVIX9
7t94GIqsuUr/J+VdPOz4KgmYJvBj7tnbdREYvx8+hXKdIJnnB1I8xcVVOUcrh9aF
`protect END_PROTECTED
