`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jonh2cdL0eeZdTuBPYHCEmt6q6ufKQGrdKWJkO8knT8KHSy+GRP/7BBkqmeFNjQJ
NmJDQFGLSXGAOBeyEBFkfEyTaDAmuEAET0aitiDmtpRMMNcRfE5jEtRUFOYnIPFW
GoyUx3k3AJhaKYSNFG3863jWjHw7Z579Hn5/NrpruMxQ9zJH06Z5S+VNjzGI+uaA
pBHWJ0Sld3vcl9EdPNY6r2RHG2ZYs7u2pb4NDWtl1pMpE9YBCrlqRBHQOBytvNHC
W9OsSDqgqHdu28Bo0TeBPueyhOcseibdK5QyTWlMIMRPirTM8F+A2z+BtA6wof26
maH/+7y4wtmGb9cWNXPDldfMu5qIAJJqVwYUPnhqiVDundNMpNWk7ezWccyaLTgz
XsFPp/GwmfRNNKbgaaB5su8R3PK92kTwmndJ60ixScxm/co2B8EqfpEhTOawoxsG
ipFgVrQo/xunXBSZCDuhw70n0JbvKuwPhNZmxsnyMU21OPZeeA0jXPXNGFOQB+ha
nZIPPmcrB+OUArlDt04ZCEhm8/SLJb4czj9f2xCxyYzVqGg73BtZiG7qiohbkd4X
`protect END_PROTECTED
