`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lRMPaCyY2wxq1smhMh6EeJEbIwmpcilLvGAKFi00oMFrCHwMuBT+nZ6f51uYWqq
NaXi8pbTYyu6bhsi5yWy3v6BErSLsIDA6Dj6y650Fs/TVEm410hptYOWyQddkiNo
XqbeC/yRQg69VbgN9qgCaYq4JwUAUDMVjoDcuzfz4uvDAE9l3Crc5kHypledpTBF
7+R6B3c4Zzs6u+ejWRp0EGyUQQOM2A6l9YDCrTBib5LBq5QPUp4HD9jgWm5niV6G
s6nKdHLWC4dymPz6O0GAcw27fwsoYe4VZ0XcFaAEvHjJtVgrdUX+5iIa/7sTQ+OZ
`protect END_PROTECTED
