`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmFCjZ99iVI4UKnd4pb5AtPuKoA/K1JVLQ5gzZZNRhQoM2wPLa8KgO3Up/sFaJe/
Lfoli/npInCmS8+WYG3hEtp1z+sp0HyhUtsJk7BTonCOmv/GPq65qaVRBRq/7g7y
9dKYLCZ6vxh7WBoU5HCy5Nqtio/uSIurFbd9jgvhQq36t3iLuJlGrlJW05u2385+
26gLboQXUk9g/jQHVnhM6NnfQLUjV5Bi/T/SV3Nke8pDlp+fdeVsNPSWK/vXeNrb
eYNubZNAAcuyp6vwwP/c8v1hFMxWMw8g4EhPj4rbbg0=
`protect END_PROTECTED
