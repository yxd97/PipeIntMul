`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2A2WV+dntO6cHzDQXK4NmNIzVRBkmVRk3FUFssHpSGinn4gdDJZIpo9iWPVpdEiV
t46RMGBXQA7nZam0TlbZU8wkX5lkVgeL7TDKYlTReRna87TWgFFqhqdpx+OYxmgM
JVK/Q7WLzU+8RABeIDq5nBp7pwNUCMvEyO/c8PidcwnzMON+aNpE27MNcBwloGZc
XTFU10rdU5NxgUszlKNMhri7NgjnEQTRaonXU3lBOAOrhKQ8989wiIJpdgT7vmLU
hnwyYIp1XKQWIEmvq5dpntAzOp1Behp1C3r28k1WdoLGMDetNQ/YYkZzPCOC+2l2
jxeESl/qCSGKTOZxrZxGEneFotfgDygauYrmWoaPectwkPzbSVnrIcdsP6H55CnS
WfZKmkfbFxRYK9ifwzPkoEG0nfc39s1TJyLEaqptEBk=
`protect END_PROTECTED
