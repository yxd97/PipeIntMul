`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVOzM8dIWfNHUie17SrYv2acWQwEq+EV20+9v3D3Gqfxx3P0l+ZTIXNMF+eQogyC
KRTT5IHKb/z0We1W9wVYwbgLRs+hyjIdEnOZyHxXZA14p7sdx/ddpbVlHcMHul56
Bm3EULorCj6YMKH+ucRpsW/1fK/bTleqTssr4Np+3trW9mDsMbPnnis+Go7tSbtp
BahVp6/EfUOGckry3R9TCvJYxSuvASym6AFz2CS2yjLciCoZTHLvGQrt4h+81Wn6
PLK7zW3d2UjGi5FZ8J2tbV8X41Lc9p4yEgzLUD6Dv0txWUR984sqEaSuGG1Zra9m
QNTtGcF7H46psrKrgjPrEzJcndeom37GAgojyM3vNwBfk/2Si2wpjyvVGRLnzhHu
XAOau3iKtk30tjd/vnd15HyVrRdsE/34sfy0tvAPGg7KszphxFi8DqhzxbAe5QqJ
`protect END_PROTECTED
