`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzfKHhfdgseg5sZk8k4vTTKHfHJ7VJrEZuXhsBzTPVi/GWuDXq1oO+08oWMJuHg1
ARm3qQ8P7FCbhxyKjwXfDYFsNH38K7AMhHsClyo6k7JzrdlXcBuohmIOMQy9ND3n
PfdDnIkDYFmCb/E1NbEj7e2KYS4JUAeCPICxMEKyRw/0IpWwgMiG/YgcmZVcOiSX
Iz7+KlKmiTlEp/0Z/TIhkS108RZaXFQTkHAsF1UcptX+l300av4IDgoEp7WJAdY5
wpuoL9BRrHs3KSqwFXLAcWO7xIA3pC6b+4lO4YrVfK8PKmu4aq0Dte2yvwptXsw0
wEwmx/wgyCXlGc9IOyyP0STQMsrMz8qqsa12dD4iFLlV1Ke4uaytnquEulMmzY31
xBMZryDUjDt1Gt1/057sjnTa7MxwJdgoVLUO0nUqV2JPhw7Aoo835kmVVCXCxhp4
wNwdpH1FVcaQ+D5LvEDBq//6ggqGXtOJNuBsQibqK+NT44/nyKwQ/RN/QBpqYDnw
ZJj5nOzVnyn2BcJh0EoRDQL352dY/FJK/SafgOyP6u8V1CWsCFzILlqVEKJNgIdJ
n+2k35I8ox7jVI+0+yrxivGC9hNjCl9LsZafKiJwnsx/5MYESa7aNaVcTiNcHmG2
KmqGTl7EtwUv8PxZA98X2jklbGpJNhkZbPp/lhZdstGxR4LHnZA/TEtbPw3yiwt+
3tK/1JRhXkvPgoHxLY6x5uCvK/eXJnU4IiQo6xY0L31S0oZ90yu/Cs4GSjI+PteQ
MBXKWWD6syPl/xu3QWO6lHeUpAMbjQXLk5gLuyddR6y7vZ8J0LGIRnNSwOe6+V2Y
s1rMDURZ3ouchV+51dVFJHFVf2NinvFEgb2KcwpiFOIjz+a8iImtNF7x68RngElw
rImMrn32dBLr07jb6av5bIzgZge7OUxd64TzZv0AbFnbYFUep2U18gkSc1rhmrM6
xVsb8Ta/bg7aO8QJAVeOuEVdr2kzj5KEq84fnAqSkZNKkTirfxdOha9iZ/bqrsI3
ovu0cFhs/vkb6wK7qKmPLujTxpJH9y51ePk0Yy/9lzztkWLSAWd+Ymd9uqiUjf+J
8Xx1u6AmI1hV8tus+mv3oCqgiyRydUGsB1BqyebUjDCKuHnxdJwZXP1h4mzqjnh5
dpuBZGAFJCZnEBPMgeVqdGtZ+ztABqgzUxA0CXRBJyzYvDohMU1MH+aY1RXuT7wW
KdFb4fEhxGj0Bg5VSfdY5gCup1PQgGaeBIaoYdzVKvwXqrPQE8+1xQzrHwypF8D2
d7ez1g0K1ieFeRmpg5ooAmBxH8kmAFN8gneopnkvzPuu/Gincvc4At4CrEYrLaNO
k3tlCoSKHrFMEU3AUTBpufbWEMTGSxHADKwGm/fgHySRjcxKD0a4UGEHExIgHjRX
lbXNOPl1+BUkapIVIo1mxyjZ9nVycLyoE8muJO+xVp5WGhiFomyp7i5ROqZs8Gmn
Bn4o9Fvo+4qRuIdAyyzV/gZlbrkxusja1CtMQPv39/y0d/G0LvkJcr0pNyiciIfe
rMxuHjOzh08LqiowrO3bi5Bcdhps79a3Bq1QwyAnSODOZ58YEJkfunfTNbHrPFmd
HKdD2pNp7G0wGYu7j+GKsmeXRtd7UHV6YRk903oxIPBCegGGBlx+07QHydXqAve/
pR0g2sihV9MGNznhff4IRm3ugJtx6VoCighbSFv5DQVhkfXAguzjVcUl9UYKod7G
lNvG7OK/4T6KG+Mt93PaGkR7rAXIUm5IdD3yP9Dc6vOf+LmRI8Z/TZ+mYm5vnsVF
kUDKyMG2ulEJnK1a41UCgITD3MLWGMveq6rs+GKaCfcOoxpxznlxvFrKtQVtmSrG
OjCj2feXxPmUzNOG+qduBx4lHre22O3FLoCimnuDNbLRNRKmH+J8+tIUIM8o9LQf
XT5F756pCaaJkAfIsmSaoeqBGYrQTh4V21tmjG5sE2ebGu76cKeH52aZQuMUVAwK
GvulVSWg+1LV2MW7qsC6T/bAZh8fd4LkOfz9MgWKuN9aoojQPmAbij5EOHTmWE/j
1KKikxAo1znOSCU06rolHsiCHT/xwu02NVIPRzgi8s5/nsq8+sozJIHtU5chcpTN
RmwkkhiPZR9weIvKLjqfnN1gMvaoyKWbg1vX2ndUoJ8H43Uu9kCxnCNr6ZF2krX1
+POJuPXhUt/7GZasBoy3J8tS85NpMZjXCfJs4+PlxNKsIjSgJ4Ox3nG2Vl53TJ38
N1iIvE4Qoqmrp8vqM6BJfB4HVma6EI5dwPIPWzGesfxSyVJkZkYj0gQHEdBcABtD
vf9McwQ0jymG9KraR+erTfMybiBEibn93r9cz0VarZ/qeMXVKb45Oh2BwWh6llZZ
E4yVYeaEaOXgeWpl11+f9QnogT56G1AApsfqp98Fxu0BBLSsUE8JGkJSVeAGleWR
PHr3tjcDRUWUnA/+s14jGPxLA7QXlDvTpH0mtxBRwhC45AEMvePyA0JghHZwHtyE
qOpkYcDX76yhMJ8EHZiCLFQbdp4WabchkKooNSOyHyWtuK72lIx/SrGC21zmjaTl
H67bLybSUmKpx+EQvLzGLb8jb38zjx1My34eFJYqpTG68looTD/ctqqCUetH7GXO
zWeCbr/2TxYtK93NlEG6kqaTFRrvUXAMqw4FDs4fZ/K1dN8BzY6AQ9x5hsuRcTCU
xhDFxJ9Zpo7DtIdAh0LbWUnalBne1nxTvC2SOEiuqQcM7x4zzXrEnBFTOvru75Yh
gMvt4BEJs+3Q9sLLDQBt1/3+lHHqaA6eH0bsWiFxuEiorj0cy0qJovS57O/kljHr
s0YzaMt+TIwYa+yFzC6vyCeKvuLiUnXV9Rizz24M46xELKNSBoS+ZnqksMYxwA2c
9cewbEOr/cwYyuFXwhLLxi+imB6CW/y81Xe5kd2VbvCbBDlh9GLiW28VMRhOst++
Aa+tOleV7r3W7W/ZsMTAwgq4FLPL0usIlz7i8YpZbEipQt7hwM70KtEwUMgT0Lm6
8irvMTv9DTrZs9QA+ZEoUiP5FfYBO6lvABJ1VVch93vOIz2OjPZAlbU7haEJBJKI
RsxZ68W9cuSev1j8EPXror52Y3o72Rz911msMktXrUV+om2zW3ucg6n6pcfmW887
ePsE3Vp0PmUSwjUoH4ZoWvB9TN92i9BPyulWdfUzfu8AvZ8PjWSBggPCc/YwbR3V
oYc5VPg0blX2h8Jq4z6oSLMnfvKlo8l0UGiR8ja9TL9jx4u8RkjzGAW4i/OD9XQL
01exi4EgGILp/XkkQPHvKoalxQ1GQI5uynCRzsxPMRsZ+0EkP7nDixh/vDBL4+wL
UdTB4UIvJe9zMuey8hw0XUeDKk40auCBWSBciRg2cKFFQV3JMsZUQ0Dj//TTI3it
5/V+ucaDQk4Ayh53LTG6sSqhdaa/pJJs4l8xpIcVOdbnjFUvPp74w0wT3HZU4622
JNe0oLFKvxv7WSHx5xWaesn74Iis7JDbkrqiRPHVHinjGu43O9/Xejp+Et6kyzXE
PuMOARRXwKbTCyJHkjxf1OhX9jcxUNEDpOvmnxYStrJvfhTjDhIaepH70lMmHGn1
BwT9gKoqS1PNwxoCHk6JYD5qfW6esbStQXlA/jAlrJxrvuhl9UBhSbxd9DjxEHXK
z62ij03UwaRy/RZmHxdEycFffFtDv0h+ojkhAiGBnpvIhApXJToBv1HpfXZFqo4F
vSpDzYOAQAnZPrSB6gLMsHc4Mca7ZddSK5ZgODxu9i/dkqhitaDiS/EayxSVOERA
kuDD8Pcz1PC+Al30IP0ui9Rkpc2EOVGrYWSi6LcLnF12fhAcMB7VUDFxJg32awFN
bNjfOe16he1y8AGVCKCIL7IgkcZrZx8nJ4IFts1iooNRbk92EuASeIwGjZfO+TJI
CciF/v9K7jnvy8fw6lO5bbwqHn2/HkyhJ2+KWU0vyn4PfK7ZtzYmDDVI6ipGfCfU
w1eSmaUPp1qutT23wODaOvOmQ0n6E4pxyravZGj0nNm6cwqhqufH9SNPiCdP3iVJ
q7bKcaoJDzjvuIdmpxVP8uk0CV3QrUVov3oWqwAQP9UiEoBlJdR69MKFOEzmq9Uv
dD4m3TiE6LJ1zVaSwMejaoaTTwfOkt0vTpkdGGJzDustguRBpzj46VoQWB5Vy8Xw
ILmuTHMJOdUCCrqK0R6oXkuXfAjCXghAEzdyU03pMrMpq9P/NjjfcTVEZtTC1TH4
dvCISnuod6wAChxYoYHjxl5PO7BPCSoW87WEvJTQqHWFWe7p4Ow4lT4P20XrcDDE
sL3h7GMTLAwJecY3WDDPYnIN5JeFLRRWaGPlxfDvIQbCd70UqdPgnbtw1Vx7Dag2
+MUAkPA42vecfaNvPYQTsH2qcP3CfoyADWAEF5gPIyB0V1jPBHcoeQXrefrDfyIX
ILBHq4wNTFf9sQwxhFxeAzvY0dRfjO99gKwIe0hF736IjBVuVO2tsu8EVCfiRKlK
tzB2R+2THUqXnujMpVIU5FYgT0nZDiTS5hugTUBJCAOzfg6x1A3h0Bn523qYSkpV
8MN5wTDnMdB3RE3TXMvf3I2tIpKB5zjQTsBQ9mF+Udyt1hIht93QzL7WMo7v/aBI
/cmeLjobmgGPginOFVa4FRsXfzITHlOK98z5j/vTOE5ToiEYMHpTQ2ki6gVuh3VS
JNEO7bqC7ZCz3wMs00MfrSVDD28EBfCxBx3+9DxGAC0EeFgpUXXnS+iiiU3n1ua9
sCL92qBXcbZ3AE1fQfBuQTfAMMLlaTbubJml6ycxo0jBfV7ZBv0ZI/56FlTlGhdv
dC0aefmN6R0/qaRIC7yA/jrO4SJQRQBz/V6gW8J1tUffoxFg2oZG5NxfrofrOcQt
5w3GJFl0LQx5ipVPpTwbEpnRiaK696XzEqzrocoZ/v3NK0kPdwDTPeNwvlqidKwz
oAIhE/nJVHFkz9/lNQWj1Cx42nj6YVVq8Odk1LAydSEVZ0rdFRddip9JIS95WzHC
T4rkGPTgrIKU1i9UBL600xdt3+spFoZPtlT7ArtWsF5JMkppcb46F7BN8bwZct2E
FkDwt78uD/qWY9+aioJtRxw13DHY/O6L66+MEq0PCqPwZButD2FQOfJGL61Dqc4t
Ff1+rqaZGCgXpgZ0Ra46dVjFmBnN6qqGSXXRNhfutvWvPte3FKJ3meGewhgnhPQu
7m3MMPWS7R9RWqPUnQYC6IBpkFhR3FLdkcl1CqEjWSVJm6VhP4GbLpNWfjQoxUUx
8Ls+ZzV/uuAUohuoI4DiFfXE467lydDftCu1F5LEUZdy6FxisFH8v11fCPPzyKGH
fiB0TaEw1uVcFNy4d+v9IejCqQeTbLS4rlRzF2hAblYLCTPVi/ozmbowsJ2wGxna
yD14C6B34FBktUuAMduvMN8zkU7HiN1cb1HfAwMljec3GIyNG44xXLUO7PBfMbmC
+OsJRakXVv070BThcLN28WoHsfJnPKNOhdggByT3GpU26q3fwr5mBS5a8YWm6SbO
qbs1vZ/Kppj2OHfJHWageWnAT2XJDyqUMkE8OkpL8v4NuzISFlWuz7fICXkfr+IE
Ri7Xud0LNb1PfIzVNoLQRdCKtQ2/GZNO6fEgRDTaSlx0GQ/A/9EM2Ab4lbuW+rwl
+oP0Xx+fivWaWMnEfAGVv+hGWAUyBzO8VFashd6oZDiuqvBNZzd3LcXu4OWqOYi5
Ebf5qe+n7+pq8Y21U7oP5b099d4Ex4BlW/KpXGVmUaIW+0dzqpINUwQPJij/xK8y
njv+mf9YIFMKjuLGe21cErhqVY/eVn4uo31u0A+YrvMgpbqMWTbSm1qBGZlvFExx
3Goz+fdEtqDyV/7GefR7aV8ohvwPLby4RF4kDHFeg1EYsHc6/Br4jZ435mXJNKLs
PVkPmaGtQEBiXenboqLfwKoJ4ysDXbM5YKvcC8T7HEo61XVbsmkhvCigv+v1xxOE
6In34MpXnJZGYpbUos+OYL4yyvYorHasSWcLynJ801Tq7sSb6LXKOUqbk78CoX/X
QQ+QwUgh/Di0u/0rcjLjkvl+82JzJ7kCHSNSHZEJR5km1rxfxB4jgvACkJWutamZ
om4KFtWhbhVYulroOluiIykORiye1Ec5S7ypGx2IBFHSDIicBKxbYMqIMkW9LAqm
bMEDo9WpCyqkECm3IBlVnvMTqePSKrbYqyYEl3il0hXuw83lH7KP/59LOOZhucJG
btoOeVcYDxxw9ZZPoXqAJkHtm6G4DVoaySM+7EP6jxBqVhoiK5yilWlSCmiscEYW
eYXGha/lKaPfN4iFVwjZnfeaVuUA90+Aus99NdUoapYc91EopRLDIFr9b2ZkxCCe
X2IbZY65lbCTBoafSrW1rpJbGvfR29bY/siFZykKLF68U8mUdSvmT23zzsRfhUlQ
qLkyEO9aaguuFEIzl7eWm6jGgLllIexwkknsnORACCskMjjhl/3yGtMQeruZ2TWf
H9OPyq1WpQnikoFieD0uFHfVWkm3wN1EXsTLMcpTlARY94XyyaBRwINPPvsToEXE
/TbXLIiWUVXP2FZLbCWOJAqhkJAwtE28IOpQ9csaJJPNdkwkeopaSQT8PVEa27yc
CzSVgdYwkCUWjyWQbHLYkJAHRESMY07scB+8szO1gCNno4EBAt44NsFYXS2NL1d1
M7JgOjbKvoZJ/nOkB/TPnV8oRoynZ6MrqCQgiyHqtimEjo2/9Uq4+hk2xsgaCIOB
J2xywqAONAITyQKAAWD8LidKdsrzKQFdHeuKCp0UNiqCTmrpQ3OuJJXr5uz30OeD
1Fvg2xYaml24Mx8+PNTyE4pPxkus+IZGVi2/WevGYLWD5CcEFHDusOe52HGCi0wf
7FLXuufvZ7nl6+zfYQDrrbPEr01dBc/H7EqF4k/OByGgZZQAkos6jOe8o1iN6Wgf
57HSM5Ol9LER0F34Juy3UeD1xDqWmA+BCvrKAO8En34/IIcLtpmpWImoQMEa74gR
1ZhnCqx8Uvk6EVtVNoP0AFzNgilB8CfaGwCzPvSKFaaYae9Y6oX1kxIjq8A7qNux
mPSAtxV85CIU62JrwTBdIdq8wZ/1pf/K9RnNli2WxZHSjabbqxOL2Xs+rC2SBcU3
+sDt6a6cqjbHQNYniEVjD14otQmFUyWqx9O8DEcg8oJwckKL2Mn76+ajkVCLokzW
8O8EM7Gscm4IkKi4k2ioGylQtzkxSHhfSAh0ndE0utdfCiUyBrtbKrfUm1eSwlo7
KHTPG6ITq6ToC59wkpAq76Nwz4u+pq4zI0Pv9mMOvfH4yJO9A0AKiB7yupoHRri6
eKxfUZCYQuXFdQrqr7zw9dI90TOhi2wfjEXrx3loUNlya3j+eBlit6czJUJErAE4
gW86L/kPctyvHzOiUHV1tY5BT2EYBF4xhqaUQCCVGRoayDl56q+JY7csZPVdL4oQ
+WSgkIg88MSfrfd2x0YwcsTyltolQfviYRdOx4YsILNKPmbbFixQh5hWHbj2GuOo
Jf5xilbKpCRHGO06jzziEKxfCmUrCId5qtXJoHN3JTSdk8R2vnk6VF076y6eNdsW
7ln2HvD1LSAL5ccxzASjIMCP3+QJtcYMiRgtf+TWOei4UZxEUgp2jlfVx4b2zWIP
nDedpNrTKs63MSJgIPICzBSwVvwsMNKd6q7GyZEp7uSQvOgfY1PHw7KJfVBue6rc
+qaJRnGMw5xNlY1hGiHUYqLiEPlAcCaHwJAZNuIZHhAu8jMynDrO2kMKQwUx33eI
tSe9zi1DQKfRCVXF/WgteszbTTN2jZm1E1Zd2uQOEtXgwK9RCL6us191bnpVgEc5
j9BFQyxlSq6BivGTiOqyodtOnxS7nizsQiX8zdA2jNqo85sHWtQsBmoIuv8PvsuE
ojTjkcn+WhUdwiRWJS8o6f5rc3csh5aTyHHiyrNLsXjrDuYrxQFz1TBBszM2Otcf
lN4dImEyynqoRWVKdO5R+ovrUZCW1k57KVVyefCJ2Qjj1uyFFqIF7UoZFMapV2TN
wT+9RmzAWeIxhuTRRNjYdqyRkpWTSml781MN4A5lzSdAUQVBL8rCq6NgcZVzKJWZ
EWGuezaPNeJ7zFuTRDElclrFaJrQ283Fn+2fuoOap62WdbPW3BFhZNpWSi9vYf1Q
lbN+FhjYgpyqknj2g2r75uUnCqtZaZP+SMoJNOUzjl8tT2TOrfFCJFq+hWHNGMPA
6L8mtkKkQ1n/ZmCHio2wHiwuQuZHnV2yzs6IvJyjLTq743VV4aIGvLjdSJQpt7ot
ay/wRx/efEx4MviFiJTJjGY/EETgk0xTmWj3X6KuXAvLX3rS04yZZkcxNsJKELBh
H1xbZEOYyvZIyKkNXLJ+P6VSNnn1JWY/yUFs6gpav+lhUo3kZ9da6zQ+ry5qw26o
DsV+k6P9DN3n0QbRA+OOo8LiNimj+b3c9W6jRKOfyRJDk1EZJoOw3Bgb0+Yy5aC5
W0nxLTuzHFIEC+HRtrfBRvWCsqvTAVVy6hEBEhGfOc+PHi85xXcD7RCv4IyNELZV
OpAQkPZpF0minNbcssLIqtHdZA1NrKqbnXX1i5y0c+KrrszTWGf927iXGZA2vEIt
7+JbxgzqwCAdhHh3nRxj5PGh6X/VJNmL+mEcHJEtFt32xr683btlZe7aNQ9QZfZh
6OX0pRbE2nqLh1XZrPj1kk7dpQGVX6sDep+BLpbUmUJ/4s1eC7bs3YQKx0RKc6Ns
HXkZ5fPhH7L4Rt9nCX6dg8YgpkigEiahv5V+IT4dpEvcB2Lm9gDSaXfrSuSyy4VQ
2hGzZ53bZYv9zExXNa0bbsgJG1E1xbL9CoGv8SUwAbr7LhLcmye0CBVDmKmOuXhC
GuiLsIB8nneh/lY+t6Qhrtv7jvzZbUBPNAWEVUEO3dAgaOR6i3cC2BHqf8ulhh0v
AAl6FfGUfxSX+pHcMB6ECQdglhTH7eq88T2ZF18UHN4YtHMnf8DSD/N96/MZliKA
4ULycIJ4FcMtKoyXBspxW702UeB4oqEnfzT6qhXe6T3taiZp3Vi6bQBQ9ZksHihd
2sCs6RQJdFnaxEB+u9Q7N7E3VvxRr+gOiTR5E9zRQ1geid5kQtvQ4O/Q2zGyFA1e
zLch4Nux6X+aJFS3G03/AfbZmlvi8xb5YNLoqpf+bhqcjBWTJPwQwjJhqHWR8nCD
AloNi7U/jrlyNyqkcUdZhWKU+IDiZlQQ0Tfb5jivAdM+krT0cKudPqU2Bn20Rbrk
2nzNL6eAfa6ZAwzksNDYadrB2WX3ev7Kb1AWDGhFPY911vFczdIlW9OcpRoFtwCv
k4zPxiEXrBMxoL41zSaVlwABKZgN6cIhRD4hYijwusIs+aVYXvYlSAlwNdTeN7r7
JwFqX3KMqu7lxCRyif79e47+aJHTkScEKURvmgYE3zSJTy65lpERraB4+L4KgOdp
eY05DGXaEs7q+Ovka6zzrjCMGK1EzJa57EkEzfxA06kSfgabAPa7UID+9N0E6Yfh
yYQfRw2aHFWd5p8j7sJ65ZPzgaR8fprH5CjuAti39Gz8F3mgPKCVhMd1H6yucTMr
Ve/pZYUGAck5WnM2w2tkzCR+1ykIBfoJmFDsG7Q8/MDTmgtSwLvSBLW3QM/rIDbS
W4KHi2SHzHZGgG1QEy1ffjHKWuco2me8/Uet+2kWBqnkwUkpn+bNI0W1eHPS9y0K
6U5lOnqd1rT50o0yS1iC0zawwyEml7X0EwJVgNYJkYsx/2XcSlKEAmaXR4I6YOIb
B6kGiBgAcot6uBF4ZEVMig==
`protect END_PROTECTED
