`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70+d1wp0t8gLTy4EIVnhH5j2M1P3o4loOv34sIiU93HbcggpbtyPSKxx0zTw1Gvz
llWjZDZ/IqU/HvebrPb3Ma9Bt3/2BvhJptFzYcnZaZFz4b+ryoopWtA+LW1Y5oox
vsj63pggF/H07HtYUTgj+/mj3gkJLTVHkQzA4T6hXSD+2pmoI4KBtri0sbwAEmol
yU+bdLYzd4xPaMARmDDGi5XNMxehKBn9Y+HgwGwma/0FkCBKwnsWbMjcGPEsRPBK
5OfKXC/KrVz/a6jVTIyYFS98z7e5guwFj1oUwbqsinejTxDaaO3ez59DqLCzMNmf
00bEIbSnYy537QKMvf3DNnzvzr4fs7jFqJnnMreNfc+rY3rQYk0G4wUTlwyEUz//
G+HrHeJ/3g6ALNuQfb7N/Q==
`protect END_PROTECTED
