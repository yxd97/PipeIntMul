`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4truuoGH3KtC0nfZl2lxOrRtrK++9FMfki9Ycb03+l2bAcUZesakthAYQ4vVoi8D
eq/9yO6E7gJIyqCkJWENSNuvZXpkAefUVa6BGlznbZzxGhfhsyVsfyQd/iytB8Ti
/kX8OgP/PLeGaNTPiGkiYBQ6ghPlH9CcTgWpHgbS0tAahwv6ll7VCu3gHU6TrkBm
3G6l7R7P9mf6Wa5hqw0R7rEEk4iSTVanl8rKNaWRnBSjaZsBJCJdRsSEqyl16Vqc
zohzgznFNXR09MpkRnMpNEGTQ0FTWqLNIQxs45fDSi/Ta4lkpVaqbk769hK+Hq8F
lDTLiFj5w3md3DiSsXoeL96klpHJOmUtbMYE5YRzbfQOwBA04BrKNKblp6rUt9kW
qXeulSUz1QZ3cd9ctKsMlNmfG8n6bRNXcq8oxlkYZ6TZxRMpp+D9xsCj41Avkmxf
mL2dTayQS15ew+rV8/LzdTebDbckj/fj4uui7F2gR/OhBzQ7wfuExXhuzWvHsfUc
fYyg/KsOJAd/tONid5DlSfZCDumPjDJ5BjDsJvxzzbWcfIIn6Z/5Qddk/LjhIh37
tyS/VVxJUkfAzmk/u1Y0Jw==
`protect END_PROTECTED
