`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NjbUmA5wBpaZV6gqUOPDaYJNfoPBA3tH3qkv7F2dlM1itCTLbVVovUuL+LdWyT00
2P87t8nmNka3wp5t7Y6LZ95o05an4bZrfMySNVkgP1SwH8XFUaAutqJJOKCsr/qb
hcGEd2D1eU1spS56GnumENGmpRIHptSyMwYx/DZ9+5qLR/rtv2qZR7VngEHR+0n7
XP8Zuh2syqhM1wV52JmY1Zvx6IrNGqMqFyTJHmUM9iHEi/KTVsRYqj5O/ELNt+Ij
M74b2+meJNYfZ3sDcyXGPGVJV5wJ6pVMCrkjpRhG6h4=
`protect END_PROTECTED
