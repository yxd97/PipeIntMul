`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZX4zVIGIPJfYr/dEXx7qACEeYIi9mZnOXiy+/Zw5Ku9c9K4SZfVYuU9QF4LZBZUL
VcEXk5BQG4EVe31OvA9SjZr7C6dQlno5NQpI/t0unF/r6pWmhgjJO8FqJEJ5RYBX
Zc2YkbKdjNp7+isXpI82aSXQO8gv/pAzFsjijyqmfiGGrZYn3F7x92vCvQkZVP2f
o3s0/u8IrrQdtxYA4LNSA6a0/tBvGpWhpbCzRG9ixa2UaXLLKhkKufUQktsE5497
U+RPQmYY69SnPiQ56ZtUlrtVcIgtYKICe7vRjzHObdpABEK9rzc5u6uA5CNjEl2Y
JV3+XUt/ohupTihLyMznw9tNO7/hzBXXR3l8Xx04iJgPENbhnd+GeAJspeBDNo9v
qdUwv41nRgS0xq5IcOftqg==
`protect END_PROTECTED
