`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WP4uQrH3qmNv6CF9O4/wP9bw7CupJGUbwXtjWxzmZiHK+pe95ls4y4KyIxhtWpYV
GOcU2an0D0+q/VB8/cLvMWf+xXYbfg9Wa23HOqgUpmcrx+QmFqM5O3dpdyAkwJXN
iFUW3dNWhDngkcjkRn6ZkUjDySe3JUVELWS+XS0xraO9fv/mQ53A4pZhk7EOVE5o
xFsgUTjR3eYPxijp10oUIF5W8roia4DdT69CiyGhg28JxnxMEMRr99RuVVHszNzb
YezTZQsrBvS1J+0krt0yJf51t4dBrqcZKHt9k6hoaS8ELmX31YZAZ7TBvXco4rM1
`protect END_PROTECTED
