`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59YdnGteHb6mUlkvSsy9v0MGMsmEn5qpz8gLgpJ7tF9Vk1dIdr3OzGzKoh7tzczl
XUsEotHH7pqwjSs5/3J4K+Vz9nuMiUrZ0Cx+T7xxS30xrt/xvb46JlcSvLLvfvy/
xzxwpU5pjlJ8niqNmqVxSJ2pxaOwqCWgQOc2fHONDbOBlxAmjix5xXrYagmazWEB
2eb57Uk9pN3a1vrg72jyjPfesjvy1uLv74PyWvSF+4pdU4+oWlWif91pcuZTJ4ZZ
Jtm0qvnHRmdgRQATavJkEBjULUWgyjmqtXMgaWZoP40=
`protect END_PROTECTED
