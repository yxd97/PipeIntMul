`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qF5FG30OHazcRcLuywUysGIwU7AStllqc1XLaIt+VJAXNegDQSoW8aVCXy/8nmIw
vtkcLob+eqVss/VwEfNbZ2Xl/Iw7f2Bo0TnA0CgVhNSmHItewGNu+ylO2n0OopWt
vyCvSU1neIOcYyko0YPlfqHQm7DqljYsu7g6iLn2T0P4g1S5/374WkvIjA/bxmMl
Uj55wBGiTLLN4FX9zvs6CDvmDHLwm3l5q211I1RlZnIVk2MAra5AbCV9fxxgat3O
AkiJAFoYALHuWPYVF/hCcYCjEalwZOkKlUmuB282BoPLSMiQXXPgzqqjyIF/I+NQ
LQfYfxAtFA1f1bfkEPOuZs/+g0G3TxFqJqTKU8jX1WMMTob4wjILUZqs7J9t3FJ+
ItfE+tvcB/jdW2IUVe5EtaKhSeKLIUSyIvNiuUYXKhXA9yB4SfE88NEwVR8LdQMe
tU5uGei1M2YeYUNOB4jWfkT4kEfYGJY3sHs+swmPSjB9psjwX/XFzFbg+7tBUkxR
ClBUFSCvhfZg7lLbd6YUnFz8zSO+RfxEMgmTa211xlo78nKKxDftQsR5P4ogI2Aq
12vMnNVC/vAzohkXj/GmjGHqoq+w7zmCgdvtjQ37KMQ49nwmGn/IaIFy5ivGYNAs
/cOhIlzT2eveTEMRlWaNGxAEAMp5nOjtx+Fg6eIwpdZL9qLU2MjMFu+A/IJfQGVQ
QjyzIiEfPtzOgwv+BVxiysXJx22buCv2sY9wNnzXY9RtOvRrjmWBWwu1jSUP85FU
3cPar7kKh5mywt7nrh8u02bNOqBwfzeMVN3LKtQOzk+56zJJkfno1igGI8z06/ZV
2JJNWcFi9A+UM7cLhBVGNSq4I1E7rzWdQ1rdRVxs4gpW0bHOgv8G6+PbJbpqHReQ
xwYVOA6Hr48naGZ4JkY9kdZdYUgei2bsv3hipyeMQOaiFzh1qQIAc7nSJ4WfKb6j
D1I9M7sxnG3J5hpvGKfAsQmn6Os8j52+ZnLMDeJ7rdvOIbFGtYKyjjeX5TITNrV5
Fugdc41VkvVrP08uTWR7RqkSECJhIwHfpt2dAJPeV0/sKRLbvrO58Sr+ZU2esybn
IuL5YawioIJ4UyLTcTcGtAP1zwxDOOF3tvohTAYaP8OkvqbUtPDPtcQUZYfSmZmf
rOe/roAEXxErhcBpPSD4UpYs9Q1vTLzdc9K40FpjOFSu4NA5vlP8hhPK/ZKuoYUI
bRl885dKgmufT6OxMgrg7FiRkUkErFxKSbDTUxuJaMPELL202Cnm7dOHZ//9jxBH
J4ce7evl7aSIKpTWxkqx6ZF4zZfmQN/oSBpbHxEVf/o1nrNvKI5h0aFQidARVscV
SL4M1Tnh7zg2t4OiCmYWn634GOsj/SnNCIs9g12/Y3ypcO2gZURNyAlFpLj/otjO
P7ZdQtb+egD0hC/y9TuLMx16YpzKUKTwEKm+MxFB9VlbFE1Yb33t4mk30C5oM9f4
3ajdddsxmgjgNptn8/7bAepuyVbJdfv6hXLvrHipZzmLaQZpaSHcMh++HihaCDjY
KcoFFB1Zsu5jyJ1XWQ70bgvw4nn1w8jwcFLPIVvlHo9VxBRn9C5FWwJvCkswncJX
OQSUYFhMwqwiP12Qlg8GfS4I82E617OGfSSi4Gd9nLMxhYJY3T8L8u6qSxpCyZ2B
OMSoq+4M6LQqEOOeEOovWBPgUqnQ+vXuUrIeDEKTTYdZ/GMBs1B8wqXXZFj3V8BL
YMhiTc7KD0CYJ6fHK+eOtYKbwRg+9vnNnwy1O5r7yqmyvDg6imM5wG6sdyFA5yc2
witjpwC2qE79QgRvf9/RMf+ISgVi2jykfWhhHnexD9fyCk+X5lg0AbA0OMNanKSa
F33Zwv05TkXATK4IKoEhIF88cfUixOi8fgMLZlbsNA7n6ixlHxMZBV2hIq9MoQ57
azAQNBlK21XZe7jocHsZ7fWjp3+Q8p22wATxKNicDwl8Z56IAU6Of/tUt8cnaInw
NQHOJFAO9dF2Wf+Lbdsa2Skd0enCieTEQRs/ytOPitu0lwRtqr/K+RmXLkFtJv9x
5OdSjts46RN11axn+kD/uIlwHBxyZF5BB+AmdNCAfyN5tna0MpxYDrWFKJj17qIQ
j7az9dwZfbybNh6/OXOEiN6SWeiQtsmyA58na89rS+F3v2QqlVAbh2LeXlADz5kj
h0tVE3yuMdMwjHSsfcreuqAob2bGQzF8kH+/K6d23SpPifHpjQoml6zGkOa1/dVh
OBiP/3Zn3q148X2kQTn4gpgSkqa28zuEPOX1srBFJSKnBJrajvhRQBS1U3DzMlp6
qbGuLmstcgIW2L0aKfN68b9pLyKsWGAGAQgjmT1dIavwo0mxQW9tCXk3G//sguAx
s75NxTJ2Ek+nvrFwhbfUBVtY0kPzXg/GD/CdkapW/O3raBDE7vQE3t43VTMXFf8i
40TswFVNDIq8kbudpnCeBeIjblabNtxDvjuOzdIViABCae2EozPlh4gIH7MnuTqc
FS2ZqHtPaXXTdWwe7jYC85qhEExZ4wt+TLFx4n/rX/ZiLlfYtlDf0O+epJpzma1f
7i5Do9OEV5KQZmOhiPb7ESwrspwzWxBo66DvTYGb+aLoVYOgMxZkaPteLkjqmOaU
Nf4usAQQadFBUZ5VbGJRUT0Nxdy9JI+hlzm2NfTcJVfyQToxPVEO8OTIPF7YdHc9
Nlndz+4wun4Mlb1y58zi5yiglTS2Gb3CT7m6DlsgRPoqTD5SI3qvXUCLXa7+ynmv
8xqcqOsGow2xlIUnz+AHHmVk7J63vXsGHqLxQqPtqBRu20WkmCoQTUMCR6YBp/sm
qT6nMrLvnVD+YTTl2lI2SkxMBdRGEHZPNmgS/nEJST8igef0m+Dhr9OjzrwYNopL
UAccrXySLbRifocLDnoZNUcPpEMR33lcoaClo/HCZ1OVdLHAaDDYaukWM6dkztyY
x/Bsg5x/gn1RXTECJOn9b7eBIuahF13DaGlDWR/6Dba5YhMv+IZNS9LkhS9mrxSV
wnAIZkU05XLn1kYoI4VLvHuC6VaiR0JdkQDWkoUyC9K66Zc0M6ya0vdtMgM34zLi
6Hc8XLD4JOztpeCcYmVN1dIcQoEbH0lcncvd8gS0YzfNAhxX7DAr4UHiv/AQ8G8K
Rzk23AAol2hSMlL3GNayWBwVdP1W7hDNAoS16EsS+qFCF72/MbHZYNKxWcSfswxQ
L130jZCuvCKXyTJdWHh9YmXr+CS3sY/LaGsp3tVElzt8cAaBTNWBzwvAKt3qfZWT
0XEshy79z9JUw6NDtLfXhh3qYrASqmzUYBxD77j8Z3/iJh38DXVx1zEEPtTzUDad
cP/Xp6pWBWOngvZqDYGdMaOycKG5WCGDLcQa5Z6z3Ol2qxFY1Vfz6sEUdCAOq6f3
LeILwF1is32f+PvMwygANy+dD4wsbzt8XS1JGiSwTpC34IhpbuPAA8lAkjDQUPUn
U0ImO0aj3FrcUMSzdRXJmV1RUFz8j69ALG9JRulyTlqviRzDC4Pvj9Gz48DP+d9u
AqJsHuYUc54qGn50C9ZFZR6ixfcVl5ldj70AxHpjExzZbfrIsiVfHdiRIa0/OPsG
xn65NHpKvlU1gD4P/nm6jXpIrO4kYEku+WClCxlBzjUFHQCGP2mmvUVRhma3rGpj
XiokLaFsaACcXeMTZUzVQqsc4y4LusgOJ9sb4mkYg8DCItKoL8Vxi/CYA8+Pty4k
olZBrVvLf/R8hzhF79Sjdc19wOuhQ2VtoOyoe6CMx0lmLcpO8iXrLEjfxZuTRiDX
EcLrGMyN1b4VJGt1bbVL/9Vr6TDC6odyqz81quVKLM9TltFiOBlmlGk6ZYVwOKbL
WuzOUQnCbZ/GXZ/QxB98ScNnIj41UBsb7pA70TGUGuBT1nAoHajGW/pB2uU0QQVs
6Cc5c2UG8Q4NELVKQV08kDFkDi8BqT59WgdAyMc6XJJAchsz+sw6pkLflg/OecIU
t/kUKCA4VkBWkatDATJqKH3DRRrU5rkLaP964QCpMCRxkDHD+tz6PkjKYMOMFpCP
dJKgahzztLPnSu5eivkzvYjd9J1C0KwQLKsg75mgA5aGLuNWQ41g9FhGspl8Yv+q
trfHeZxKFiRAAG1MvPNgWbBCSJdLv5JSJVo9K/26TxbyD+jHtryAbUY7SaZzRSKH
VHI7WZ+S85K7tKaGePED+5hF+r/Lgw5NuSJPL9c5YvJU9bDF1/prKYLL6WEPgGz8
kMIF8l3X0PlD9ryFETct7rRhotoObxRRDCRGHS0VN6i9tvTYZOV5KyOCtPPZNdUR
ouvK/GkhslrrF25wqPb9gTkB3/iQAKz8WGKmEua4WKlinpkOUSfRZBEomFr2iBX/
Nly48bbJWnN4Zw6sG/32Claxm7ZWp3DFdBY9IJ5uctIzIC4afotWhcn8zmb6PkNB
xeXZulkTPVghlzzK5e5OSsWtpvhHlJdLQbI17u8oqPku0r6Xf0Ed3aGfiOMExOLo
Uh5Vr15fsTKGsIFUiTHlaf55KCHKvx0DxXgJUOWkkmImjGcmz8fEuelMJgsUDBQc
YTd49kKw2hRsp20bgro4J9lmsdXG2fbtEylaOPl4nMt/9vHfdfjKUM9o1gXNcKY6
H8ZNmvkaKm7hl30sx3M6N8eWX1BkBny3GzJqjKNGpVEHbibP50ClcAyhaljNyuH+
RQKhRLbyiPuw8ud4IFCc3EdCVpQOppb2t6kBofRibK5CXZlkJ/8U+Km4XbNtybmP
MggU0LuIzozR8zj+tVHpumlmnpARgrrXMENqfmzQKN5AIpMBk281C20GdK+hKJ/s
82ti0zTFZJZLTFTzUM+qc1CCf0wn6mATm/cgA6AOz92DVgvGLk83eW0msw6mXeK+
mn2L69tfKixzMvfPBaoPvCvyw9MG3f4GsDPHkXQ2wpcIFbys8x9lat+UvPHo8pdO
l9eb2aaFvhYhCwTCVD5uraNjCiThKo9ZvkcTQKeYRCfMbYGFx0ivq2HPYAn3L3/e
yuCOZM/UjMtchh+EciZUO0isDlGnXduqtKdr74jfr1sL1hfBYC7k6mDbWlGHJO34
7aqovFkPeRn9//U5wTJ/ep4/TU0FzwrYjD04h9o3n2y9C2nl/pPNGo0FyClLwHR8
SG5AU95QBNwEP2pzHi7RHKiJ8Go7lBqz8HyL5kWmX1QMge24722xPSNgbQ83v2Q5
ywyT31apnHN5v38r0edXHnEEfswlOMlLJPBud+vgx90KXRDL7Gc4sg4ckJVoLGB8
NOE866/OXNwWxx+4rd5uVPpjt0KzACZ9nB8kbfIlnDcDg2G9b3SKzYjXwwZMpujl
s/uxMI5c2mSZeeMVfj83DVJIQRKwPY++44Fr/wWuiq0FRswfOeTuj3pOztdno0uh
y7gzL4M2PGn/Cf3tkMiS0BYN+eKDHm9sI3R9fCqTap0jsRUfn7/B6gWrvnvBY3av
YwBs+mC6yiTt8fRKrXtB/YU0r1hPBqEis60MpJAarz7OF40fPF4SsKI8N+2iq1Fs
6bsIsQzSyDjD+xvDYULILSa4Q3FY4FYJpV4avTRjmaWF75Deb75THFLTExq1ZHFz
PaJhnQSr35BEc9u6zbZBDKsLffBStHkO7GlrsjsPzAKISsQ/qWsaE6SjokkRvLd3
DwAVOmfn7mIOcWWuUCUQCINHqM0+WFTqkYkQk6JNBCaepI8wiOiB/03KYVyp+Szm
ZR8EZH7F8yoEf0MGcZfPhoTO5NCKeUlmtyYduSC60R/LKjg34dM7PAiJGck4kt3N
XajnpaNQrBrnYuiZwqRodZLgh5UAhtS0I3pbeLxGJIuSXyZOVz350J6SERNq7dHP
EoRZi+mxgmGQHHQQQLKQxtbarfASsDJ+grMdjJ8BySiou+0avha4pd7DvzZ3HmJZ
MkPFrgB4YEQiswbIG3l0hbRqdBVGGRQokg1EfE2YKrjS07HmKWVX5k2oe7zEneqm
/YtPffA0DbrryH8JLRZYHm7uoei7dsqZT3AX6mA6gP6wadN4xz36w+wUK7ZFosIU
7rJymoCK+Jc3jXHpeNH08v26H2v56t9FRP5B6nxwD/97fs6BP5LdoGZFWKAdKXcS
J3dNKdRXVjhX7euJrLl6LAL8q16qyA+EOnZfOBxPr9uDgsDsh3cGVLUQ77sf5TsH
xk7SPMc7+fBwRHwP/aJIshQ7de36SdYPiOtUJnWN2qvfkZlT7dfI+/gUwZHVVcu6
kXu8S2o1UVrcYEwBGiB82isrSo37bFSFCQW1PHb4RrVUwnx0DYmUsX/AYPaYY3mm
ihIvytv7fRokUfvi0OreqctsR/DT96kyGo5Hl0brm8M2ntjHvUBrRnpcyBLM8HSR
PVsoN2As0q19VHyodD47BuphPvKfmyFYYa5htxaImgMwTguXyOrJzosSMwei8Je2
TreVY6Ex5JErMT+zplBCAWMWA9Kf/VeV6q/ggdjPS7zh/mGmjMwHyit00JX/8yVr
A3oyuEFPl9xZBo4uCGtrkMR/AKB2X4QYJoMbJF1Z+jePccMlqDQ2V8kmbExzRuuB
MKk8qCkdn0zO4L71+S2jBag9JTEkB1fnBsHduy3gn42p+w2A57jXEW/980OvBlkV
bZgyp5F49Y4Giy/RmCT2slKrEfi4asSsv1Tg2IMwi0CpRsMcyeacYTGKZTXJKROs
ddf4BO8mA0UP4Vix9LczD5Ph9wCTLeODTEC37fb4Viu67cSwu5uGBiSQL4PbLoa6
TDoBhKykhp352wYx8OkWbVk3o7wi+FKH3OSAL2P81Zubh9KpNtrsGaK/krU6t9K+
MyjZrCd4SCN06pXU0M/0MHuTWsEIbm+QAykduH9ogoL27qpJsehD4XLIPElkBOyp
g4WMqYolAe/iz6njQwDQxnStEE9hp3AjGJwOeKPtjDpJ7hCMs0LhXTbzNCYxj73N
M3xzQDHvHdR72AHyCmQa10Qdrc+7WMYxag/sE4oTvFEZW7SPmiZNtemVS/Dys8DV
p1tl/UE+8zPDNtAY0WHrA9eWdd7UX6DMhUf+WGWxzXvstaHt1VFRbkZZujVF6ioy
yGJa3+STu5uXMbSHtv0ewVXpz0eMHH7xyIyEpxTu6/RflOs9dzweShe0MXTBQ7aj
UmdsQe4Khudvtpd7RWIviD7gxxX2uSP28AnXzrPswyrwBYijR8vtsjKo6rLMrlha
c1xujAku9IEJ2nYNBzI1AS+h4EugzgWUBQnLZutGR9kAqnNy0K5EKLe7Jt4FS9y+
e9179gzxeOz8ev8eB39c6Vj5zbGbAJIxBB2/oMzGnl5rAH7D68tBrJX5Qoq6VE/+
Cg/mLL6jUyj5KYMu5qTn02lTNqFvyWsM8g0ujcKvF8RsnHwj5Veqy26bjKPvQulq
MopCEMcP6ai56Ts3N8gnbSPrbDHrSH95uX0YbxG0RXZJVolHmmhaYJRhIKW9RSV6
ll6fF8F6Kt7QiVAYTwYMrS9G3TKTEIgxBDG7uL9eRiSvyaR+XlFe3NLmcwp+Hyku
7R8WAgBlAvp2Fan6Gs/HYPWrDaZTVBJK0Nl+YLGMhXMElOBWRS7sUqotN4mr05Jd
jkxiiaXlYXktNVfuWYXTFg+UM8pCcYmY/AOEuCC1TTs8jE3EJH73CHZiij2P7+g1
88RlAtqmM/yrZsCtPpM0M60auGd8m72BWBsa5g4JYUzRjDNfsEBmColFVIFXikqE
PVni2bI4amsIDTKtsKMIoG5KfCx7AEFitDgV98AaWZNVTK392fkLUhQhqMDwfmah
HcvMZF4NJRJOvF5L5/d12qA9WMlwsjRYkskLvo+Z+YTfuPQ6aeNNIF5NqMFZz/Fk
cxc6XzmB0u2ldMCAQteVA35XOCYbtLIwNJjGn7g3fQwLV4jO/e7aX0If6s2PFyJT
ZF4nxvG6u7344WUivOi1I/0QvBkLKsf0acfmSXA0Gt3Tv6vUVZGse7X4NUTAGP+n
7FF4xMjiF9X5XwQbP579Tu++VPxUe7tH7RW2sqZYGQqZa3Fjq74M3Rtp6EX7nAmJ
0lscLBPTf4c6AfMmy2OySDVYqlBDUseei1eyr9m3F5TRN2pNbEseK/YYGe3HwCyL
ml/5ScJnlEOmdtZ5Ad95wrnSOVCUTqail/UqTXExHN6fmQJHGScMoaz4893dgC42
abAtlamdcxzAQ6LuVkhcv6BMhjttcbM5g6PxmvBJcn8SBvAYPhgRYHE00bDYv9S5
LUIPKntTDw2W2vxA7GrmflUviN6sXXUSdLgNvZKwkR0ZAnye1kQ8lNLZ/5EJjL6J
bpgNngM+fmr+ecdM2raB12Bgtt2/Y/PtBr1u5TS+Jl33nDp5jV6rwZg4hUGU/zFf
Sed2tGhwcWkF9cGZjzwfGZyl5OcVnMpuI6WfQ/N7mK8qBhZYv5yJyyzc2kntVFY+
whQ2KjLyhU2kAEricmNEAORFAuwjXctOK61FZb1FfkKdUc3H1J3/6wXXNrgPCtYd
aoWJVAd9yKMyJeVzY7H07k8aJbNcZJZePjE0lknR0mCoJ67VFkKbYK4Fwmt9hWl1
zpUpU8kEJrK08hbJ1w2n3ES1xyKtQtbr2UPcrUVj8VEMEpz2VMthHqSwFoVXAlGF
gjX96JN0JoFf06wMkgQGpiQucjQsAA5CFfvgFIKp4xe9tatxmT7Ff5pe/91szC2D
UeRkKr/ZHh+ifL2On+bde5IEl0f4aKGngfAHb93XyJqmN02/RzRb2e5OHeRThU52
olJNxRPjwCFaAUWt5wSTzOP2135SiMVP/cUlb33y+w0gsONiV5IG8CjUQKzlhM0l
EhzdwmeZrz+Ya5S9Vx4qj/SQ8Awk7K86pKa2GKkEhQHYaI8AJXXZ1OSXuwTNcNZb
hhcyNonxgXiqzC+sy1ImY4wxUgyLI3ZgsH33qOJ/jTAtceo0VXmR3JXO10mCj7z9
z6vwZ9ZIWkESe9nR7iw+/H1/U7DMIOtkZ4AlMxxTay3xDgPKnGvAE/cUdmOJpU+7
0LlkAtGxmd5mCfx65XrJElpKj3G0jGcegj/Wr6WA7yczXiKImWe7/OQoIGVCh+n1
Lmj9kJ4ES1Cc6jKAAURp2b6NJOcUBwSfFvTsygmcvJhYsWCgGzXuvX39UhZdYXvQ
1dLqyzleo0B+HcPzPhlB1LbSUeXxvs6pfHLybIV9bAbDSu+4pLeiDpoeCdEIv9Lq
03Bu0SSanAPVeJEvUzLZKk10nt7bITqxm7pq/Avs38OB1btCq76c0wENk8hlulV1
GO38pf1q+Bhuw+5kCZKBjSGJEGQ1LL3+qaawsKXG4GESzIj+WBGbZzjqnUOz+L3V
hpn4LVJufBSpkmPb7dKmr5t0V22K+8J8dcM1+/bfghloz2x7Er3CeyTdq2IWsegn
VJ/6maKJaoPut5e62OLalek7MSUa6IV7G5+HoxqSLGC92KI8dFUUr9vzb5JzRjc8
JF+q5E7Fl4ziGXG/tiNjMm8RfQHmExJn+jgXQ/AIOIrvTs3cw00dR+BsIJdWHOIm
Gy31Nk+f/kwy7fq/s3280KfCH4P0l6LdzvUsdvDIH/VVsV8G581fV2KsVHHk+0CH
+lD1EaW2sPaBRfHDSEh4XtXu7E9aV34P9cmh1plQk4nLup2vvlFGC/+BNlLgj3yt
O9UUdWJ+lIN6kTPR7R5bRvUSg9uiLvA4zZwPGa1CO/phQYZfZprKYt+fOZWsmCeo
liCo8DRYBThksg+2/4UucdDMMphPN50A/qIB32KcUMGVltOWNCzb7/O32Kt5u2Ac
fsHtlwe40mTVEyZqsQanRIfg9xwJ40eg53Cb/pA76bIwWk7L1yRsG/JPOSyCyagi
8EW+PXlOMSPnEPS1TOIwgwPfrAv7cQpIc5aA5oeey1n2iNnFZjnQFGvRA8YXCS9m
cUaE0AG9eZiUoh+sOoYTi+0TBPvO72znFtk7+qFwzj3b86w3p6JyqFzeQICMw2IM
KcE2//xoZbbqCP0IotglEMrB05/oEO2dS/tjzF0E8QY0UKpsQCBkuivwJyg2vv1X
vraL0imHhvEWel128DG13tFKEq1RQrIWUUbxhbvjG2JqFigsRHNzVPb4pQcFRffF
gajuer6+SQQLvzQFIZLJxyLLgFgfC6W4F1VOSQfrjbYjdylKg7S/ZZBGTsheyYLh
vHGc3k8OfpV9iH1Ic7SiqfPTkzCzGVRZPxx+fBW+bsI3WDBIrN0sk4fJqc/VO9Xo
FZ64Xsd4IVK7tsiz6F6fzse6FBHXt5MDZ9zfxVs5qxCnh1sYnkXB8kygqDPkKNBE
SlxxxFYcQ34VONTkdAtrU/WBWy114T30IKRMnCLdC/+nWW1k83n61KNLqVMfd9Yd
8s+TfFvoDiMvXGNP5knWOnyXa4x29qQb7ZTY5b31wERnhqLo7ttzUMpLEGOL7PCo
1d6xiJ/F0VdVE5TWKoFp3w==
`protect END_PROTECTED
