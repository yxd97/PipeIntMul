`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7lGihG5dAq7wQcwFmVoEFqsbPrLw872NQflvWN7hv/ahzmtnIdVaUQW7s+tSl3f
jtVsSC7z3Q0TAulLwcfzOd2Rr40xMVb9aS/BnjBbcaaxcArJ9e3/lDgx1D0CpQMY
L4i1hjXjfEaNq0yuVQ0mLE1cCXhFs/DK6pk0RMFl0vtahnoE81LkaYSCxCAKxe8Y
KF4YCppqotofdJtBgyIo3zSF1Zmzd3RuyVmeVW9x6Z4wTNYDWienU6NaXGHkxFdA
AyRRCZDjsMNBnV2tZiRO8EDmTSgkMS30dY13d7JIFuqzUIPrczi/JUlPZ/z3POKh
bFpFBlKByNcIFyH993G27QHXxwmBsH1cpnxO/Nl6ayoUqZExW9oZey3SyvHVWyH/
Wqk4sqbMml5VycZ7epC3rLW8jX8zPndw9gEpaPYF7xjxwnP1aoRWJX11Nz77ugHh
mQKb3lOgwOOXDrI6LbHYcpMWOKIMS1/BL0jrBVrzfK2l6pcIwAXkOBP+1DbhqztI
tm3+8XbteveN/CbDNlWrJaEsBBXmp3iuuX9uDP7aTQABncGdJ7Bv47n9eWm3O9hw
FYAI34nPDCGyupj0i58mg5s2KiGxwf/HgG6wmQ78NPliusOCmjvPKystfh5kDKAr
`protect END_PROTECTED
