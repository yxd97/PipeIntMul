`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dlk0PWm6ad/pyD4UBRy23OjvFH4ObEXDNnCJTGcCtBZyLo/vrgMqATiEfROJONtB
wWGpkgN1EDaET6oR32698tEB5S0HSdTdcS1RWg9b1yIPWQFjdq/Fe5ru+9+WYM9O
oalPaKTFm6UMHDRJFy+HRrMp7N5HF/TwmXsOIeWc7hoiBFfCLkfV83ag9mSP1qY+
2Bd/2fr2ymQw/CVPX1Lk2RC6lKn/eReqLa/D0cAE2UzLkfkMrRpNOTeyRACFFG+w
4xUgEHRrHNdsW0fXLH4K7s5PBImkTgYKUYMIbFr3saFZhCwkN3Bxdc8gVmqKxc3n
i9PJE/60ha8qS2T57c+Tyg==
`protect END_PROTECTED
