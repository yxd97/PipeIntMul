`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UexDUkweNXIMHVFRufiVd/tHji4qXRYs3L3GBcQjH2IDVqRrJtLHWB0/w0yjQMxY
5bvCJrJGLj4V1cxkmbljS4ozYlCFS8I64d8u1qsMfZO2Nm1ZAuMya9JPCVL2C7c9
3beJXHogNgoP7kTLk9W8L/42T/6DjD9bPv9fYL65Kj4VReYc2DB0EMxdDOJnjmNU
fgqZH5Khrg/XPotuAn6cMqpOIbAF2asn7XC7tN+pKXmBDXXxBDVjResiCmk5Ripe
aoT2IqttB333EIeD4aDxW+M3SQPZsJt0lIgVUO5H4IzQwvEUkNbWA04yTvxEtON9
DjsnvqHQ2kcAzTGrLWEJrNG4y9eNj4pJiAWCaVYiCrdGSjkmE8gPxzNXBjYxDr1e
87oXakIn9KVCxHaBwBNDmUPf7SpIsm0jsNJP7La5Gn+eamvHsEWSGRvOAE1mIdlQ
SCcAq8qGOoDbHJpeUdWBEaB0Px9cDf7YytzobOvuXlbiB0OTbVR5HKTizycy3zJ6
XavAGLtSf5N3NHAAYCbIEJf+L4BXX9knZ2mHqBSYJg2CT9GztFISaccjs2h2ZVZb
ca3SDP908RQoUClzCGYGVbbdEbNWvA47uXvo6D5i/jqKHG7oc+hMZh4d1Kr0dO17
P8c46PahNj2JZuBIhIM1zsA89rQfKXO6Kg/vWtyuHdcSt+xN76tcvhhdt3uRRwuX
dpcXay7n7ZSB6slXrSm2iJ4omDNuyYCQI7EV0AJyyrodKv3WZFmkBWcelN25bi4j
ayMY3wu1jif+hApdqcs6JFiIXdMBDTnXp6Ky1rx9DoJJfEZwtq5xhma8f5v/DGm2
mM5azgANsiVx+y+1tVvkpg==
`protect END_PROTECTED
