`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X1osxpImi3gtCusVeS4TSPVBt9LdFsVtAKCWdjCYWS7LSwI09zVM4iE6YLSHe/5x
BvJJ7p6yhSJ53al1m0/kP9v8iB2gf659SaucmiPpEiZdwrC+91EbbDBc5625mD2y
1XNG9gD3eyC1XK55D8UqupRXtslo5ybdxszP9pbckJiDLPeI0eLAHuM4s1c/i7uj
Caheg+EEobsGXyxNNOy/8KwlByLmD+FKXSFbowUJUX9KdQf9ExzrESSS2lwOOXK5
YePGBOV50sIwZoUiuJ4sFCp3HzmkGgrhJBLbRoKpWjZYdZv/Lgewqr4Lv/RXqufx
TnHYe0dmMXbZyyfOKi74HIu+TMvL/4CYv5nAu5yZvR+nvGVzsG1PgoWJLyy8FpoF
rOJ6IZBG29NfYI1Y8yY82iLoqiTfJ4wofvqTq5korrMjKdmMD4YF0LIjJYuzdcZR
EgZ/rQXHuf8W42Qk1vE9RteWXw+i4B8Q2+RD9ZgiA19pXnIwP2q/enu8TGO5BuAK
PiVi8FzaECuNXkzVy+q7veuGwJ5FtuCSHiGVI9EOt0AWIdIqXygz2SWEOoZe4THn
Kuf76lZ4RkLbZZNhV84g9kUcJy6Tfk5RhptOQZS80NAIUOWlKxm/jSGjlv3irV89
nUxaUNkKQJ+cen1QOVMYthnvTL0I0r8Bbx9Iu9DL+T7w57WkhwjE0J9lGcTb3gmn
ai0kewHlqlGo2BLQYTKcFNZnCwa8fh+0D+lgN61NiYAE4ZwrulhcyqQf7QRf76Tb
ROn3KxCkFAKexLCHZXiD51Ofk/6DzAxpThHaarOqi9FUsquYyBOdWwutt3FvsWbk
JUGrF3wK1p2rZW/S93WO/HabPy3q+owA4NRCheus63DoJe61M0hZp79iTStlvIFv
Gx2WOn6nkMRv1A2PXgnK0dX5UHLwFA7GWZIylYcR+XFeRO5cowJcE+hbXSpWSmSg
nCzI9m8hgUPmWRJVvwR0MN6pYQK9fi/WBO8j3VrwNpRfnUlRASSQxisrEIj+RYF7
k7/STt6iNB5+ZE8TxtcjHvtMdGkB7s6hogx4OHbVkOU=
`protect END_PROTECTED
