`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXDxrrXFcdS80KDrSpoh6eSmrd6KLve6Up1bSkwSPey54fyrIaGslx59QaQj2tpi
0CG4+syFgZlRHWAh6b0VyEwz4lSv8li8lW4bsxi6CbY2qxuRmcIkUQ0XQ7rRtUb6
XKwp4m6+mWrs+MiSAoal04w3S44xsDiuPQAo9Hx2XuHx0gFkEPG1oGl04X1FIvtB
VS9LmF2Iw4HECRlLniTBr8Kv6HvN+ItR0AC9rc97DMq+BH/NAtTBHRsQ+puzjFSK
0+H0/rcvptJKVO9Fb5VYTJ8Y77EVMDm1Z5L/TsHVYLd9psAe3RiHAYhMIr6KDTXg
8SYcUszSXlMFemQku77hDsR+248Qo4q6BhBV/XxOtP3cCBxmQrDPibZFxzQNkZq4
sjayAvCvlx1rxrIz1/MK++X0xoLvMHnh91rTpv5PDKI=
`protect END_PROTECTED
