`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEY+ZFoCDWY/JCM6BTXV1ma4YlSD16QRJ4YIKQkaTK2o8LaZMtU4fR3zSKu8KHkD
MPbwmV9liV8bIy52uJPb8+ZggTvPenYZXPHf9JVW5mYfBr5Y/3g9kx1ZWU014352
FaZGjj1grbdRUJBAe/nY4vXCMz/hkc+gWXaqPdqk8Hc+cdEXXE5N9LQAyb+5cItA
uuKiorEPWHN4VHQRdUF9W/XNpg4ZuGhtpSRSIMJqfMTN0Y/L7Wn0Hty4jd/FfWE7
5URienGmvTqP3MPhkH3bjgZPmNgcrlCJuA0q+RzXJyWFab27XbdqnvWQB25od3Ad
PonPU13sO3qhE+rONkgOa68Tehm5fTECP+lzWhsVSOgydOgQNa/DGQrxZScb8Izh
pp3B8i1yQN14onPgeWD08Q==
`protect END_PROTECTED
