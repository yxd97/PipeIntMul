`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8KGPeF9l0PbU9a/+QixzoCGXZWe+6HhpIXET76u1YYwZ+swTdUq0JQ/zI3TypZ2R
kLz9jlx/7RAZMNNXOJd06YxkK8EPvu6wfTKcadkFG+dEp2Ml5jY5i0LNq5kJBBVa
mHkBupvc1f9hyep4RrJnya0Wo74+q0Esx9V2khtMaMf6gHrGpBBRYUiM5bF4J11P
AJmB4/kugEMJW6M9DeY8BqYfKAlawMkOkLWpG1bYh4Pzo4oe2lIYntUuYmePUT2S
`protect END_PROTECTED
