`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
04ZHB+wEJrLBh2VCV0FJhSzuHT1cYnKI5lY3/xy9SJRIJM0/a9f/zIi+kotbwbFt
TCYExhwMMEeqgqcnIuc8DaYq2Vr1lKNk//yAt8bBUrPXockRtSXfv7tRwDCwpCTP
6vefFo0sanZUoH6iqDeg9PgNBv6oTKPUv/uhP7cy6NLe4llVq8/JzK7uui9koTid
B2Y0YqMapQZ3CE8JcekJixqg06vPUNeJQG709H+W0opBfD1YKfecMb49LlyE037/
hPXBKcOEBluEd/IWWobqtKOhGI18kJgHrWzD7LrGT3Ef3FOS9TqxRVWzlDM2Od3P
6GrgtW07h9juUsNlMxbRDBKtreJBCO/Fg/BaEXi+CVJYkgRpwNRAxIurfVl8MwhY
wydXBMXAH39q+O4iS9Lvt6iG6YGMjGcLVOCJiVCMzyovMowWKlfRcdmko/x2V7vt
nYlZs9y4i5684WDk5sXS3Ygr+t9E8sKJzfs9XEwtggo=
`protect END_PROTECTED
