`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nU4KqqNatG9e9fGL2TT/ru25t0iexayrRltT90b7NM+UuNzdYGQX23QSTF7S2G5K
YgTkgoy10I2lyF16PtZKiPM5Q2qA76KmSFt7UCTdvGI5/5RpaXiuo7Fp4yJq21wJ
ZxY55ThMAonvxwd1YGf7y+2dwwMt38iHfF2BHaAC3vI1OpN/Xw6BWLoW+Yh3MiX6
EaZaZpoJcnCtYXsvDyo0Qb699cFuv5BwbME/CPkZj5M6R0/5nRi31SpAQUc3ksNI
pfSSahRgyz0XVvlLzso34b1Ytts9MbVAFGF8xENP3Hd89PZWfmrSOLae6y/mScIr
OSK/yxXjR40yMBAPAg1jwxnkEwvPj//Ker1ydxCZaG+PNCcHUhTR5DPSKkzaXY+H
fOx6zKw5cgQ3nZIRofz8hQ==
`protect END_PROTECTED
