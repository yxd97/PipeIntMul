`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tug1N5eUmPO/tBK9rY6IaasA7LAeHHgQhWvcfkks5prXhkLWEOPfKRqJnNGkReQ2
BfHJ7OYxBuAvPwl7jPJEw5uooweettOh1pdexy6C2VSAvNL5Up++KZn8D3G1gx0D
T7wKowupoREzQcaP0PFLf/fFDUWa5xNkQFm0R6aakLQa/SkBzPRoMjiRrRpK4+YV
jDYUG2u02C9+qV+dbcVu9RAYpg3U7EQypEaJISJaDdqEXhyXprsg2eKvnZj5s+Bn
nsKEcVjcJKQksReU6nmJlLR8cZLcdHbd7GH6SVk4QBaGmVVeN3X56pgVcxSJWgwb
S39k9Pniv4Gr0W2SsEcON//I/iAovxdNnkgE/dX0M2vt74PcjhwJQ1lczx/sJZyH
G6NQcpgW411Dqw4RARiUJpFCVbBECnSyci2RQtL5JDHJgqVoNsg5NQUmvVXB7lgV
ggmFPcK8i9na4xKv1ZWB/wEi3prtCzw1uc2xPKCGrnH8wwTYUPJQmiky8+baVw0j
2G5i98n5BvlmqUSeyVIIEcdPA7UtoV8s+7Eh+4Sn3bKay58Q2xX9k4tKI5F9qi6K
b81m+C9ijTNSOM6Ho+LTlNmyhF0l9fvEcp1Jt0qUOSw0K3TJjz27F3lcDSpw2Ob9
2bXbiOUaoiptCgYbOkRV1pk8scBBgkhI60IaalC7jadM4u9NMZhuXGkb9xpLDjsh
LpFAIm6MHBVlxYBiB0WZ+QENwZ5gbV3RwjXDyKjeDv0Td+34RFvUgexjuKVyJwlc
wAHIdKQq/7lqvweeif1LDnLyR6iHOUUoGiN6+8tMjQwzLt6yJz5iRQGDmtXC59rz
PDfSMcrWEQ14cLSc27Ck1UGofwoAHwFz4lA4uPe4tlB7GxbJ9GwBKbWW5e5+xSJz
+j6PaxYuCfnZBm/tZUPBVSLExrWX8dI44v7qOxS6JswqTFr2kGF8NaW2LovjPlSD
9kyw3C0xhkLSjwq952hVQpilKLSOFmKcH0Mx1qcFeQNcaPACX/CIHBWRpKhR5wU7
TE+pwWbc8IADAtPKoC2GcVvnODuvrP+rPqivkJSKf9TpvDrY8V535FaifG/5dflp
kZx4Qwx25LU2kHyKp9s7PhKh9x1TZpeKQd6iTdE4QCOxlV/Ru9lS7V+dD4ak+V0e
QYoJkBfBHmg0pKRTrHbvjr21Rde+Rq6YYQTxCOwiZ3gCUZThN41J76HZgDU1Vn2G
lH3eSPp7aUBxkwfBnxkwWjs8HWOK5zbltJESQLzDc5rOkeZPwkk9Ez+5hWEGNyKe
9Viq5N0TmKo8KhxB5JlvBOT5iq/X3WjzwboEUJcmFvXAOyr8JHTwGQvf0eZ1qbxX
PAp5SRrWX+sp1ksOafD3g+ZB1YOn2nqoZHdnKQRQS95XmF1xo5Fy9aeK1b/VrHxJ
8VVyqMY74o3rZXlk5Y+fctAjHhgbVqfbMzzm1yRcBRb50jqQGeGeAJ6G1mDrtkJ7
mItmxyzK0qdojlbhFGbUaA60b9YvEepdGAecKnpcO2nUri7bxeKdhMO2kHqsYvLA
h91YXVZoSwVmjzP/3i5NiIY9SOS2tv6WCPJo9v5kZuCzpa5iGY23plIAoLzIjQu8
YLcfNfsMfKGRjBTfkKt2MsV5QZ8KBfsqKMGJvmVbs4tKmxHZtWWbjGOWxsryef40
adQIkegQf2hn+BUtKx9KmiA7FuIozX5dZXshbx/ormwluSkwBmFY7Fay03XDyF6A
X2Rtww090MHtCLdw/JGlCsgs5Jakium6azjFtz2hoCI4QUSmDyN9iWDC8KCEWBc9
EK2RXi4FQdHz25iajMTY1TzYUSy56tUK7ERrA3b82SzPBrzN7lllrrCAHF3Orzdl
GF7aihTeuiCgc1DF9tmqyc6rhMp5w6pZh0mtQ6GhuEEwUU2enFVHrQRJEHQvHrqG
Df24BhlCtXcxLEILjKR5XMGfa71R3trTPQuAnZrhNP+jQbp2gm6VE4Xz3BrYBWxh
bVM+tQ6wE+OAZBSdmtQuV+FXuAihgxBNRRgDErUyxQkIDfE7Dxg8PQ5TOl1i9hiI
d+4W3mxj4Pchc+oRvQBX79zKMRYH7FPGsujsEl3QEp6xNyuZGL5IOLtVz+WchroD
mhwmImSxAJa2ib1smZ5oh+gQ9i+79sMle7fZvLvIUSr0/8n+fGuF8qZ7NEmeET5f
rFQRQxsGRN1Tj0KHLOGz1ZQ9NkJfTpeTCj2JQWynY4KMn5iBVTReh0oCbnz1aIQ+
QNd6wkjpcnZgdi5ecHbkg/IAKOa6I+Kuj8lH3Jgx8gDgYF0m2UfW8pLnBMxqbaiX
c0u8Gofw7GeCvK32uNbFKdeQaEgavnXt3pyXW1b9sz0R3JwNvRFSPPBWldGZaOO9
ctT9R2B63JscAmBJYQda7X+ojIEDP+Y/WdJEag+dn/0eboT7N8geOkX2AntWx+Y3
HfsCmN0GoFFMYJWs5ul0J8CF+cxshKXJrCQAREbDjFlnGQEJByLWX/ATM8XWInr2
gsl52zqekXzgzqlbpJULWdpv0SgY4sOHQJBXc2aMuVDnTC6RWqHZQudqK4QeP+bx
hcrmGE4/mECMqSARGIxJ0fLK1KswzTNy4qm4rDvd74PdwKlNIKsqbICJt7/1vfcs
JZc+essU7iDHOYS3NP6QitXEJMhapDNj4ryljtUeUmHXHvkyoYq9y55QCfr8rhBB
2RamrBrispSLkSdbX0fpTX2/DwKVpJ/7FaQh1TEYiEAOmBqg55UE48yNhn1zIKJd
0bTF0FEOh52Gza/zKZFm5BI2AoiP0tJYseV2SLJH7yIaJABrKRLFxcWXqMBvUz47
ZGTms9jC1qkS2gCfLgqBXmePe7TfDKGonONL90MatplT2n5kvrV9uY9rLE6kPuIx
TiqpM09XtrOrnq+Z/uXfvHaRAeZhYMP8vGcAIHZxhjs3VhdTqGrdOiTugZnZGZH0
L0GYCbE2uzjdoO6Y3EJqF1LttdI2iMAcBOH2xP3reWMbsQmBZVSForHJWgjUs4Er
McThOH33LCNthduTcGSPzHvKR2invwwzPYqeXBIpvwBAvyZB0zmAFV47gJmqk8zn
dwiscRIisSa+AXD81/uE1XVZihn+KJ7N0HdGFgbYKmDeN9QUS2pF10XIQbulOKVu
eyutehuSkfVCMR/dGDWhNDObQV5NR19+QI7KRyNEAxGjSir9oMBt8jgcVJxPuNHW
k0kSk+v0jvR2JGcoQO7vg5naSszdnbSClHlxqzi1yKwnL6TMYfq9DarkKJOLr8jm
nS7URkr7YItCi/+wKzBNBGHfaUpyW7HKoRgCEixR6wYh+j91Tf8bFyzTM34m6/t6
k8ZRF5TK0m51P8b3RMcfF6zYF+u0nrmIPmt2V6CNhEKnXymOOw+/s9diCpxryduc
geEGO5uT0+F0L227xIxlzUSbmzGhwI3JzbxECARNhkPBsRNg1IAI4dc4nO+DnTqB
Un/kA3IFpuIw1Vl0T5nQX8R0g1QyAF12peXPFy/IyBLPlbaZmQEevEZG5Z7GCJhc
X4AGzYoeBuqAxQbKlpvtsYdRjU7E8g9dFGBiUH5ISjAtJlF1UCUaDl55pvSF4EWw
DptLfm10qLkOqspbx0pKLqvt4NmxkqQ3hHG0ABHvCwDnvkJ+8zSz7P0wsKnJqzug
RyEgRo+V/OR3KJEjS+LA/NNezpSkXp7ojksQLRrHXaQmNhneL4siDvp5vTRhmkxi
/KloEKIbDzHyuS7PpTFCM9Xj6ZsyMvaWENZY98KPbSSoA3yQ04BpRLS/rCUFqijL
AnkG9TZRmrsK1RWuiOe3GlpjgpP7isS/XxreukTrNBfNVFoTaXiW6zeoB7zl4zXr
z8fuufDgEO76LqFvfQjfgyIs6bFGc8W5rU3HV3zlxFFPfmAeh/iBxIEwRNeCS0/g
oA3Y6AWKkxWCpEjLR1gPPRGeBE2j8vsxlz52iO2/BkSDzu3kmzbDbCBo+NRnhLtl
TQ93oowcZENMgRpL2T3oGrCPEM0bjPaw4dv796m87jO91IN7SiEjT11jxXUhLi+H
WFcHIeb5mGsb9UH94+aA1CZKRg2F+2uS207ygbwAUkT91OPJMPnCkR96yKA6MybJ
apttuzAqFN9jIaNqZYbtLlK6+pvOR3ugMseeUGehy8Z6toCp1Jj9TiVhqtL5Mj5W
JVlQOizcr82Gz6cKKxEo0HgRkhKwPFBvpXVqLOlCcE+7K/kBwXNX/itymLPJBs+F
m2sroMa5XpQUR4g5vm7rARVSeniFHz/8/eBrio5lIKlfM3bu+SXfFbjGK+2Z7zXW
U9ubDX5eKH5BH1sbHGy3cZiyw5N2fBoK4Bof+0+J9y57XFCYkWBczjcJJHWDAaag
K8EUPJ78tNqIn5KXxhmgtl/It2dAM9ZhBfOkuFdbX7JtS03yOqyYjz20nR1D2Yd3
PGTYutpUr2+Hy2VViTB8MWG8eUi3IRXMHeKhzM2hlVrgbjiK53SzI6x3+CX74cty
Elj6Usg9AG2zAS2fTb5jU0Ywe3gunZDrLp/7Oqvdkbtvg6nrnuO1b+1FC0ceOasS
B1mTQZrG2kkzKIrnVUTseRU9jkwdZaBod1lsDWDy9Gd56QpqPKiwsvkgeGQAcS6x
Dr6lQmJObu6OsfvRCyEX6SP4ulmFCceT5FdxsnZ1ZVfye+nPKR9oBtltaUuwRpOj
QM+NwgRHQ5IgIjyisSp+67GDEHpTAxKIEzVs4I35kjmuo+AfTmaliK4BF3aIJtnc
z4l5CV+HuOV7loY+3LzcRVCuIJkDfbsYYEoJKD2DUBsv/0rsBoonoHZxWtiP6/hn
UdamY0qm9mPvBPuVYwqFHq1lNyisuD0mdgs6ZdXYKlJ+EfZVTVE5EF/PedBrPPI2
Gs9m48K5ncEhuN8sSIIuDNSecDULWsABmii4B0fQJbdPzGXphKa6Za6nv8a7pHNB
DRuT2s6O8vRWsUQFtrCPSjMaQzmrKAGL1anH8B/hke6HZWdL68ZkWj49hWrnOHku
RQKQIEt8LotwVrE0I7h5oYozpx5U/Am4sen143qJXatoDlwSKJhzAaL7ATmqR7IV
Fyx4TPpn96gHMlrHSWEX1eJN1MSp5rJH7N7JyG7jeNOURjWsQkbIMCp1Oplm0q48
5E4/FTn1fW2LZGG8vDhKkRe6NvXlwViXGFx8vxaDjFgSTM+zSGmd8TbX7I0rC9VF
v3xmiVBmcjj4br9Lhg6sFBRyxV7a1OMOLz78yk+VVC9or/3zR1shAVlWE1SW7R5z
UuRYc9Kly49wq/TtUozQjZVms/um+UOqD+c1rgMd3FrHSmMhLLPt9bXDxEi/9Vck
25YQNaOp0ZUg6BpWSIcru5O4AX2+CYSn6U79Vi0JcjIxRwp4M/f6YoydRkhCPtuc
YTKJCYjzAWPHtHPal3kauvJ4hWDokMMAEMH8FGl9/pDUoJgZwkXd025XHH7QxFV+
Ekh61bM5MlK4rZXzeqTAD8Yu2e1grIlq/BMJja3NUpH6Obf9SxGkDdWfGmuP0DoD
N65fbhCsbCQwbRQ59Lp/oucbjuYVGF4jzgC2cqu4ENrzWLpljvONQKgyA2ApYTbc
ydfcLu0sI0TGquH4V4PBJACsmLGNx0sZb7q9TW6y2Eic1S2YVy8wpwZ+1wQbu5Zi
J8SKo99IcLRw1iM5pl1K1TShEgHYq22Jbjc/Bt8g8qi7ns9r14LRAjOf4J1PnMfz
hJaIWC3bTszG9dyo+m2MaE8NA4jquBoczcWKtwbHUH27DtCrHPXwf1UIStUliOjU
HMX8HMNaREUWtHpOAZvo2XnjFWdzUGseEmxXhjbRffjz/0Zn1g6qEryMWHDNsCkT
E6EJ/XRohAWbmV3fJL9uGMwa30Wxd0zIXxYs5B7878nhyFe+OMGVZDYxtJBZ5cnn
jPxElCuTIfXyfOzsYhb93fT20eqMp6wi7cVwS9pDCNrCKXgaikxNnfuDVYUL55kl
Nih0UByqahEY28duCyPd54Xil++o5gLgRxz+DFpL1Udf2YOEboU/aRK9XnOg0aqb
K8vP2Hn4jnf8zVtoTZ3zVHxB0aAmOdgw/ow0ttKWkh8IZz3HcUNNInBVkrLnD5XO
dLDZG2v0zahzmnNoD2CL1bS0bUvIlDnZv6x0ZH44Blnz+Z+GkxrNekMS7LSVS19c
hQoQHRgt+tdUQ4cRX/1J9nrYAHyYWQGQzwqNVj6oNbxN/dH/RCHrA6OtG9hP1L8L
Mqc8yWcETpywhhOSytGNnu+ipZekTkZ8Wx6qukTZOn6/3a5UlJJ+7t2ggeu5PS2v
TtKhpFc4G9qAE5yF0UZdqM7Gkmm0leREZNfxIiVA6qqiy2x/2CulYlvBvwqBXDwl
UHaZ4S+XgxKJscAbQNyBW7Dbz4C7g/yE04RGaR/lgJiKXXJIM2C0xQDA4IgPUDl1
vDLwp61+PR3Wb7mnBTnu3AsypNZvt0R74gdJpsYkC5J8FkRIDdnXWQB57mF1hEUR
d3uj6+Yif0I8+fIUa7h26ag0qCce1i2wUS4TUoOFoWGPvSaOc6bBQ1/kxVHfd5mC
qG7fby7wqTEZf5MeN289kebMLfsfTucYH5/eZKgaYgYgq3r4hxtsC50MfDgZbtZG
5uOeHnbExz8xxq5aiuXtrZv/5FY3JAAZlLZmmt8tKkdRowYPUQay+ZuzAqX5aW5j
k7MFdlNs5+5vrJUGIpvZpa3YkdWGF0KIEUZjh+RcsCB/z+PvUaEXkW8w6qIQGXUe
aOjMbxbyW//FTWn/Me39w74Yg4s0vFWUaLAgDdZxugaGZ99644A/2DPxnE+lvQfM
ClBQ8QmjyJW2R7rUIP7s7CMaOFkfM2ECjS7N+Th9Oo+Zgt1YzmWM/MoFGrX58ZWf
FAogzEoCRHWlOjrCFzlr1iqr4kqI9QeEQLwdHObLy/5ByTyddvImqq82xRz9c9Ra
VxE5pZmpIJ4qFRBOq3ZlBgs9SjSl8fNXUx56iqyQ4GH6aI08D8sqPIUt9tSqF/ar
v+9SYXer3uOeDJ3po4XO5d3IULxMNXqk5+/c3mH84wkbTgoXpDajt9TB60xAGeTq
tACUvY5KeNUiAG4K5JGxf/RJS4T4Sy1lLosFrvBKYVHO2dzqunYni3/6F1NnJuWa
PXZI/1K8lNFcxsRCcAr/C2jGBc+Erw4Tsiox0HFMDD4W2TJIUl2EfnFq6le2u5eT
+ngZf2Ng4WqKP1GhPeglyEvctwkz11Uylfio5rlDPhriXTbraTozZ2+Cj71OgSrR
BKbFG85Yr4EbOuVJJeoR6x9lP91nxvPdKqmISlk/XthdnUF67hzb4lgTYVoPDzL6
NX2BjCuOkGcFr1XabSzgRxef1vQswrPRnrq+DPD2YC5e/2E22UCj4jnYYBiwG8mv
+s1GKCBPFXYIF/6l5sgUk8WFBdOYhyHnUz2VBEbq/opkLjDt/Wu+X4k4+v0l/AfA
39izQWJX2af79ECYA+P0yFiNwZG6dBQOtb3Gms7tKlPbnFmlK7VgJ7egpvbjRi1Y
ZlfykHm52n8aLt712vFiii/OEECSVpZ9RaKmp3jqGA5oF2RNcLtFjXbhlSZfvH01
lwpC4bCE/lptndBPRAV+e2z1Pxwf5Z2xIfnGVPiYYKasUhl4OPjKc0YVHKoMmvAV
yRb3Q72RbUsMUIgVfjwry/JeYCgv2ljHwF8FQbyx3SDvknoCQ4DZqzOptG7kDPgn
C5J5JIHNIJF/rggtZ+wBU2drhm+lwEl6+ejhOkqYdj6hKaX9gBYrxTp691ONi8jD
fLBGhsv/XtHddISes3n9HklXqYgawEnZDho1Dg7t62PAfhULz17+V9R9R63tSPLV
NIZOtkqsFVzoD/8CkvGiIBiwQVAwJrnzoSHdyIzSzIK9RRvuYcl9HItGBJ6mUJcE
cdkFOWFJrqnL7JDLv1VdWomDOlFnt4LVYpr2mhfgBS/iD9Xkrfo40HlTQZL7JWv8
kPC/kuDOCesr2fo5mt+0K8dtAT0pAsugL1TlhBBIp1gYBJNvujiA7HlrXxCrVYzH
WprM7FgxiBoGXLTKE1pYdP0/UI93OgGBOMmZbOYHumlQXTsXKkLVU/LKuLtSsIGJ
WYnsCWSpZxoXZN36gvHjveTI/Ozp+pCgkBsM2s7W4ZUVUWZmAZsgp6W1sGOqDMQ7
O4zL5C8FWQjT5tzX89Dgdl4Nx7hCcGGVoI9sy9PCDb1MqtmncnGGjo6hxRS2Or0Z
qYhz2xKyfhneDtsgWXhBRJP4fqoH16rrcQoijVOZQ3J7swgCnIozXIz3W9fqy4Pu
6xLaAcbIbKoKlLRxWs8G40aJ7CC8xp5DBsZ7RoDi2SaNBe9wTHVLeJpmSUFvj8pR
Q0q5ISn+RfYpV3ovcagICQ42EVO32bKlEOqG0UR2rhz4CjCqBXxp5i34s/S1AQyw
Y4XSopq5AdCHGXrS2TZd8BQqyge1tTs2W/S+UYJLUZgsvN2oZFOiKgqfQLphizN2
4/YNlUP3XYqNDJNELXM7vrXm2TOlIg8U7S3oBrZoUp0QOqjT6vntuvdQ+wE/Q31c
S+fAzm94OqPDEi8GSMVh542sgj2OfpnePHRdJu0qY1Anhwfbw1pvypX3DySR1MGa
MssEcpL4sSd77OP1NKDFNuL/Aelj95iVk9E1HdVJT8TZA0Jn+ow/zblrtHKsvr3m
qSre9VElXjGxlqHnTK+lLZedxrTXbyHKrPhrx4GTvFgTF5xsFmx0yBrhGgCDFChh
4yrNKfbwMB7LtimYgxZRwNaoYbQTViZ9gqs0veaMIv88vG4lKuUn4U6Fg/ccXf7c
V863f5vkZAfaG2ETdEN5fT5uiZQ5+ImBdyEddoSH13aJ+7sjQtLBKb3IZnlJKNho
pkB3CXCqkZQkW7UqMsfn2cTbRSMNmuhlxEshgXSHVanqaMbgRvYmrYaoOFJ7B4jb
sBaaMs1DYhAV2JO0HmBvdE3OsgDQ8bouECsEXk8/4uiUFq4w8t0chPSf0hFZDwrI
NZ6e2GG6H1y0zA9XMQx3jVoG9ZOIHY6sE9msqHs09IQq1bUiQcw4d74yatFYbkJS
p0f9C0cPSR4Prd9o5vykL+ltER9MBiIacLXSBGyNOl3jP59vlKhLo5nUt5pC1f6F
dUPSG2F+xKXnP5G3WWwqzc5FSFovE1f/OLmdjUa5hDB5844z2UA6i+016xIS0MVQ
IJ5TEPXXipJBfKl8u90UhPAV5mMH2JOg1fzGg/z/9QQpuajzmpypgkFFxr2cPPCk
OLDv0L36PWq++JIRni4mw8HtxP9KEq1wKp1OlT5dh7Jiurdto/iMdkuu3/1Mgxh3
H7VIOjMbPutzntcdKHdVkrcy3K0pmcvcQQ07Ta4i2jWJUg4/Qz1HcNSroee16RkE
NDs0oZb0dviRloMfm2iaFJnihf+81htlERtdjpQmFdLb/IC8RgAJtDWk0+NhGTgB
ucbkrhJGpE97OAE8xEem3FJGe+UePUvia8tIw8Cp4I9B/NCGrHPSMQYwMUgObt5W
XMUeqKetdidssKcUewJnV7u2J2+Nhz/mXosKraparG47oK69Wx6sU6HZw3zyOIZD
u6KblLdKgWJWITBI5RlF5TxVhKPvPxl4GIG2tOjBzra7HtOn/RFCdtZM65Q44ar8
yyGYvumRa8+n+eIGI+mBcjwrQUXFP8B4INebBv8imcfkjTYxqYe+UNpELUvmflTy
+LPMGEJ7u+OCduFSh0qQlT0TC+CcLX9UIx9ezmiikU5H4BJRB1GIF7iP02ZlQgob
I9DGTpPt81SuVb8DgD7fBLehzDSVshT+xcAhXoOWLOzf8QqpknWxeNUIhb2O1QZi
Fxh8bU2UpE6vqD6M7xp5cVcwpNNNX3ep/mLQn3jFzr1sCZ1Vp/0yc6KzRbS/dFZo
5RFbt4iE5OsRxKJYkZg4oFLQKU+qU6A4gDiVfj/LuOR5a/mXLnIO11/7fDp2dEwL
RwzNI1o6R3TxEZ6PGKDNgc2pfUcy6plmocZOerFwtMtrZ9McopzLEE8F0KzJDYho
JSx1RHsO242ryLtdBogzsV6rbv04akqdIPktCJUOlNppxbBjVMNi0UDHnSEITsOA
/Hzf7OzQ+fxlkh+YUo9G21zmViWyENFeKe3WHi0eIpu7x87OYfTuaOGtfSp6qr5w
3ErfF1aFWUduLXEp3hgVMNysxLO7R0StMDO85ukNLD+3hZheqpUA/lYq2AGGl69x
9fUL7JvzXdl7jN4L0NgMw/TBO8lNnzKuzE4hU0i1K+awO1V2HOuj78mUd5k23jyW
IKqBhoB7UtZ6fTygUCP6HpeaUhC6uD9625KhhRkNvu6CzQ/qJYT7w4DIHbPnM0Tk
GR6mVfSJzzfV9h4sUGYAu1xp/4pd0qvoEPjhWaue2Smj/htCJWigI7Jlhjjz9J0G
2+ikfVrl2bZSheZQiSTFi7hPBNi2NwKNdIudwkeNk8lO+RE5BCCTLG4hbsZAxy1x
GYd4XEI9hHOwADgASa6aYZT8qndqhQDPydPzktskmWoomaYj9mA2V/B7dWM5zGrN
iKmHcpDTXaAgWedLJAuh0G/V1G6DPn38QXJdgBPg28ePFgzoAQfeJcA6x5saB2T5
3245V3+kzML2JoEtJVD8Vy0bC29+SUrln6g6Zule41/TyYQrjfze2HBLRO6qx3Ft
kxAIB4HdlREXjOyxMsWJgz2ziHqllfo1iA4l0xhNn/bSgujaiTJ1C4NMoYu3GZnn
IXhLv+5AlcXMMVApYnDRj/r3h3itq+6RpMJCy5EhVD6piCZWYuV4igH6RuXAJdN7
2Iqy+OCP8k6GNPjFQfPmdEpulFqTO50RizY08ORKuudMA7SNEqZdIKfVQ9zNKVIR
JCkGufGlEk/IXqgcX7L03pk77dU6yzAatHKyq0pfw508qJW1zitgMzR00AD14su+
y/+NOxkzvvEu07quaOaTiulY6A2tR2Je4U3JP2G0XE4lMPvPUS4ANO8PhH6fclCC
NvHEqe5vHV8EURRro5fN6KYbklkF5oft9bqVYkx/WTNcilPXPaaixGUel0FsbEM6
bOrE3XRDW3fduaVrvtWhxWEN5VU1udF/b4uxu90K6bvAzIUttTRzun1NZi1qNkAK
fL+QL5AzUBt2iXYdhwNxS4DFu4uon2Lwm9aMgXz0k2aHXW7qPewDUY73YUeU5UTd
/JKhIDlzO4DA+TdPw3VP2q3q20uMInogEord3bjtPIf/vx9vpZvFnqnDzUozI0Xq
NzeLq3+9VyNAC1tG3qMPXWAl/TtfIgp+s7lppDRXZtzVAA99cXmCkntxUveDCVFn
LGHeXdax+GtQPpyGwVxXr/UStwJW5b5farSzYx4a8xPuGwGJU3m/Ul1124odxl5l
Txkc/UQzww9qmY5Lod4hxf5IvsHuVdcpHZEDsbTlJv2N/JNZdYG7b7GLo6YlA12X
jI5ArSqtYIlGfuCuA53VceTJaz4eAMtqXyagJnIU+P+HeEswUk0mt6zLdFHVr/4Y
q2aJPF4Y5lDyfp7Z/Qn+CQo8iTbb17JTpHIu4LEXg5MbXistiDvy4+hAywLh1Ao1
gSMB94wBAyatAlkhVRCkFjUzwEAU6/FkWXYt3jU9JXvX6jXgPPf1jsKe/UAenOYj
nVKkdqOT08YRwCoN/BsVkvO4Nv4jZ2xt2nFLleUbx9Y5gspl2CoVIgGtPXN8d/9d
tHZU3r0ymaICaS7a1NzUW4M/NfPQDfEYioGxLGcn1R1XJRBkeKcNMEKlTL5rS4N+
v7cO37ZtrBSGOxueFCxUKDFoUcbMwSJt+P0gz9J4Sd5upKW5mnNkIxPkhT0iIQSt
a2Cxbv5G8cySVvIncTI4iWGCawdo37j8Tye4Wb/Wbwxks0Q0zKLNDEAvBd1KKAn4
bqepGl2tVL13RsRI9AYwtJN0IP+OUq5to3+U0M/aO3SWiGDa/IwqYaJj+J2mLqbM
kpSb20zKEjVdz0BVgVKzxdYr6js45Qv1BwO3Eta07penlRlLAAyRYTqTjE20YOz8
dUt5zi9lLwh237fR5EmkrAAhdMVk8jzjl3hf42WeNo5Sn4U2WtAF5HiZI+vF5owc
4SANEQPuDQ9b3Rt5ZZrK2vEapwvH/EsQi9qAG6D2EqSZ+Nfkec07On3/b5tEN4Jh
18hzVEavlt2B0HKoYUT0ATAP98ZEthjP1WhtpUA3mV8BCdSzbkzUBdJeoavTURDP
Wb5a11bRaRErH/ad6z2nsyCVjkDV2V6R+yCoR3a67CKkBDyEGjljZlISBUPAq98v
rmcLSypi9HJsPx1Vxgt4MpC3XKXTJ4EmZwPCd+p0kZ22FtWmuvxjPbjFE5vNV1zq
or4va8BPISuS8FS2NX7T62i8x876sErDJX1G4GkcC3FjwtJiNLxVJALQ5NftEBiA
vw7mPylJKYYLG2soD5ElDMYSa5aV+8Rp5CvsgCdVxpyBtL5tsBCK4jeInGpNpodn
nQS5h9t9fPff7PFWYpkqoXjqvKuuyHoaZZrzlinL7qAjQloQGIXah5RAyJKrBZQL
3oppdS24qq1hedqCDHtqALhM0fQSL78wy9OS01AdAy0HUdDc4HsCqgmd/UWHLAhl
lFRmw2ANut8LJcR7Fbt1LbSWljLmOOCb/cyC801pJqnkQRIw8w7ZOvMwxAFpQT21
irpc6FrqGM3EhQyjUg5MCCZtlQWBfN7Y8d+LnsYav7dda5LFB3zRBSPuhJhHrc9c
2k/CfyKYFYzP2va5SCXTXoSZcrT0fEL2jF9Jm6/tFpGW6anAqu8b1HJsby1UW2R6
frPb9hER9L4Bj5xAvhkHGktMiq6teNmg5S+5g/+LwVQCNy6e64cTVUEmfgBjLcyc
+3N7JFbrFCw5AmZKgv3yLEk6w5A5vCrEtMw7pCbqi1nH2o1pTDbMhZRQkwjLQSAF
Rf0UnLxkciIS91GISIfFaAx+hkjrlvrn/ueXH2Oa0iRpqln2GMgXaacvnP9ZpB+E
syqEI1Rlfw5XxUhGR7K+T+gq84MSJ7ksZzMigp5No483DwbHJMvLew+6R3+YBaK/
MybipIjTxYRUybfBKyigDEN99or8V+7eOMzLL8kK97kSe9tALhRczj+EQUnSNPtV
ie+AfETCYwryVLLJ0AAr2CjJmYKCV8csJSVjxNkAw+lX5kdJKmY7hd3WWnxUXdo8
9jwMI68+Jvjxlk4clkafHn0kKoLWN21IlYbFBpegWHa46z7ubKWsbhGVKWrAXwny
xNKw+lVw8kyQKTWSwl+JBtHsUs4V0ptwv+4nWVfVEq5z7G61q14sKrrSpykc+GmM
TyvGCm1Q/ph05qLMcU/40n+lF9sP1aNIWbGtfBlwEanFMwk0/jmX5X08YSB4EqMx
8KgyC6uJZw/cTa1IT75M6zIdBrWx071+K+0mRQbij7k//IhqJpWAJG8qP8AaPADI
x2Hvl//8Hf7We/cMbs1ho+kcB+PPWjRVoaJHwYtRrVbQk47sIa/g0/IVWYypTMAh
sGRZJOZRe6w6cn+MjBdgCKYcJfsNKXgTpKcgLAZRf7HYxtGqEu1uYseZEVxPLo9v
OqNsoP9oEW+uxJJ5LlVj6Xqh5zqK/S0zdFMTrXQZzfL/EMmArje5AVVkmit02vqB
+2wxH2cQmtbXlLyrP9u41RfVPZPQyvDE2PgxEHmzF+gZTYEw49juKdTEpq1sHapd
0VgruCSDo9ggKrWoI3SQy1WclnSxUsmftbQJLTjnvvTrxA3Yt9phPWYc1dMkUtia
STz/cNk2VSEEt62DIKt5dW7yvF6nQkZb4/Ofelq1O0iFu6/CXKDN5PZVyWsk6QXE
p2OssqKCFKEt0Y3O8HVsMpWeHwyxcgAvUJ28q0MagG0zj3jnDct9aiyNCaFt6YAA
i7oJXhP5cH0EQZp2i+jTP8F25dhC/2R7Rat8sfESL3y+mmaYcbu3Wsj50X3STYtL
3GbF4vSVPngn8A1pwWc46iILncCX87FMFX4jaNBixUMSfsyHEOnFubS/lOSY3sQD
SnRLNI3FnBJYEiSNBDohVo7j31HxywG0CUWHE70V1rTof6bh9k4iayScPTy0ZIX4
osJLfx1hHNKqElcR+WscYTeLJSmzI7wTfU2qJNaQZ4SyuF6K1IIhIVP44rJ39GTH
vB8OmPNZQFnVz4V8p0Q472qxie07mkg39JrW+y7YeKl8cyibjbXi/UcgID8xXgAi
s/KcHIgUSJffVNUv2UcQONkrgWa/Xc+h+5ZOfXVo3xHap2NbhZq1AZJscslfbUDO
sMaDx6mXvNLgtpxHizozTg==
`protect END_PROTECTED
