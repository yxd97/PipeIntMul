`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2mRpBO6ChwCIB4SqvBc46LlOdlHboPUh/yUAiLdS/db840SB6taFAttKOaVJnZsz
1J1VjVmXVLdDbwOoMq7haOnvaNZkI9TU1FWhx1UNECC4LMY8ngGBnnAx8/J7aAz5
KWo2L2kMtpWngKWtTVUcrinJcWuIkXbhIaIxoL+tStfbABAXwFxq7cCbXl0ThEP4
tOetOrDE4UVQ1e0FOdu5Q/6KIJ7bWTMdlw2Gr2o/rM8cbwBtb6UzH37Ya+9n7Nwm
JtP5JaImgfALnBqiAJ4JsvIK0G8WlKV436kU2cCz0IKz/QD2KGbBBt6Qm2ECPjS3
ooslWZWOsIc3elE+2BYYijmXQCovq7ZYcYvcntbZZJdHYL3/WtEbNOFmn7lwMa+E
2+n08DjjUgcAy8b8pQhdinIdOaL/txl3gUEiLswKh5JkAYvl7hDRwxigmapOzjJ+
X4kSt/gFZcAR2yF7G78zy8Yhdr/V5uSji8Zdx6SdNUJl9glm2lTM1V7uS29+RSmQ
+QMwAhSTBmZB/o/4v6boaBKWhiLhL7jEjaYrsmn6srpZSOnI08aywWtCvwoog0S+
T6opcW9ZALocFdpwAH8Fy+Pw+ZiNutU9zspdbcPqHsg=
`protect END_PROTECTED
