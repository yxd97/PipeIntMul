`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kq4LsDXXSfoXsUaBKlyrf67lt9lIyEg7lZWtatflqS3kg9M9LGgrPh7arDR3gJm8
lrXjexh9NkqNLEjzh9a5PiUTwiuqK7z/mLHy1zz7VlO9sOqw9n+A4R+p9vPOE+n0
EhPBygbbUf4H6C8rjFl1lhrmRs4XYb8sRUiBliRVqshV0mZW85iYqPxVUvAH6ZOh
2a94Kxz+vH4Pg4564PiBN8249ksuSxRkIlekbXPc9JhG4nDonvK+zvzKlPY44Bad
3+d6ns9orPqTt/0+oOR8ONz0IImMMmWumd/XYAXjOhtNjNLqMQA4LWUNox7Uoa8P
0yJfN/Qp4+X9Rc5SesuveEQEKyhr4sD4dKeM1W4nbT5a0YsZiGwz16ZBZ4P0LwMA
6AIRA1VfST/WUke2xJBLC2wQ8O1TumqeXc5yLlQhy+XWVcLAS3KhE1+wh828s2e5
toVLKVGM/U9YtXo5a4cIfOqfYqlItm4NO0xWTLEJCaGJ3MdB7UMS8C0k9D0fgj3z
H2PuxfErP5fV6G1Dt0JgwEu5RYStxg2yBAsoQzqYx8efA51nNK0q0f3hNKhJ+EaD
2tiW0SYKnBnr2kcsoMqnOVjLO9ck4v8XxLrWUpNs5eYwE8ymZy+3eJZ80v3cCxry
Mr1rur3kKBCP4BCgqQt3nwodWeLOpAaTyuRrDCRXKlEdc1pZ59Q9pofJnGMMtmeN
YKXEMpyRSnJE1LSyISHi+A==
`protect END_PROTECTED
