`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8xKznOJmk4rpD/mHujiaBOf0G6TCLKGFsglFjfYrHfs6BCfDo8GLvbBTvRmaUC1
gxvcO0dwYwe5FEOoOsTOJSsPFmPkecPCdw5HwHkJL+E848CazE8ZzM/ppZzcL1HQ
Luq54j1D6GnJZALbycHstV4c2aqGOg/u3wtLHPOkwNi1mchZH2Oq/jBFensH4wOs
yDVcauxr87gEeUJ3amQgbycvkb+h81SzzzMprz5bZ7539MyV/2ZzX0jPNihzXSuU
IfEcPnGShZ9yibidxLImoKrGj567LXvJdI4E7cDwYSpQGyl5n1DLVgLB2LTSg9iU
arkmx+qLpecGHjCG4i7pZ7e3bZcVKch1/oVMT0wMvBUcga+GbUhlc6GAPvD7fiaK
29IeFT4PfGD5JMOTq7NlmNmwho7qMR+80jGaazkhFvbTfeMKR+j3xdZZqQlrI7Eu
U5/X636rmaPgUoFXn68u1w==
`protect END_PROTECTED
