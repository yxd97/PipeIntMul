`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2TSHrOJX2D6WUUgnBP4uaKYyYib5sDsoFjiJunwJDoMjfHr4FYaikfrxt0C4MhL9
GYdD+C+1x3xX9xyOGK86N0rUzuH3/uLdj3/OKZAouvwU6Zk8a4xagBUymSvqXp2s
FREjiyRYnlsdhA+gk7iPu7iVyrTY5z50DYMQdJOAVOl5QdHElareAsQENXHKtEy3
wb+bpvZcBYo9qX8jfEG85WueLFyLOV2nSlFUhxowxd/KgBCNs1GM05t6ZDnMXElD
JXSYwxP6SyWbnOH0fhxbMh8Y8b7WL30Hh/DAlb/qnuxYANGU8XGRpxCRNFskNhrA
DMkj2rqLbOiRNb6A0XNtO0c7/DsRXKvW7En6JSSPvW/XidwpSbWU868tunZjCQi8
Mzo4QuPr65tWT2BgXxxFZoXbTEH5lp481puDLLdokUoOrmKbM0vIpyjJOJi2LQfb
VoZJ0aN39MF6uKkPPMvr9Aq+zJW9OjNadxYIEmu6jksAoQ4A+Nun+i0vMUU+DghA
SMYF1e8VVbqE4O1MmeO8BjuKJ7J6SKEUVa1SdfeIoyua6q6eTnOxOdkvCccqyIA5
Ifk/81KJqMrG2s/cgHr/Tw==
`protect END_PROTECTED
