`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k2JOLcVFsLqzDQ+82NwVikqxRIakvxbi7y2xPSJ8IRH2x9/qslsENYtBwvYVsZso
VZMNOebCncUyUV19HqrHvAHg/KOM7mUVhP98siRH0M6lYy6KXMK/r5syyl0b4P6A
1zHCQO9yfR3oXZ9JRZRyAwFjOfuFPLWoBlQcWVRfwdgXNXOrLw0BuZ+tNQd+B4ZY
cGyY5MAkN+4kn6T6KDW+KUX8OfUiunPORTzvVcYIRd+eCmrURVi2xiPhYnhpo1GW
aDkyJC2t29NFykyH3TO5MHi5Y1oQFBMAxtvO9goeGIUHLcXc17U4rrzYBEuJuHbM
0OIegtyYoNbKbQ1XIst5xi/z6VyClUyfCkEl0HqBqLbC3Qr+TSMuteu9EpQN83Yw
gx9v5b0Nn5xbvPKQg1UrgnzTekNKKbBE6Yml7TYXVKm4sIT8pUr3EqMzZgSPJUj+
2L6jL4p3CE15A2VV7erN+xQ6KCeQXa2GyM+cPrlypiEE8CidRtuP0X/p7FCk8Boh
`protect END_PROTECTED
