`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sSeMBlUdBiVWKf1159kf+LiQfAPimCbtoMmbBek762iFEsMEi4dT/3iUfMimLPpe
fzSAyuNKUz2xWafh/tY/QIVy3rQgsy3B+k39m8fxYW0ObQ+Q9hyL62vlwOwBvF7r
04bdpInd7skQLH0mGc/QsznvnHeyldMlRPS5Ojh2aOQF1Vt2wCHzOgNAvd/eJy4j
wa+s3x4L6RyMgV2LkX5vTq5Sj0TfX5o9nWiD0g651Wi7denTWtCdsGfki1lobuFX
bE+UA8LsHsMjJWgjyLeKvDVESZ48sVAAaUz+Reo8lDfRtYIv4PN7SC6M21Qs3MOf
qnDrxVmv+p8ZocTSVhy/mnKWB1x/erMbjJbeuju2QaL3TArqfAhzhdt7RU8JvMsG
OJvE+KPFSpdU3lJG6+2dJ2WwXhEQge2JcB2+0O+YOF0=
`protect END_PROTECTED
