`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uy0w+Uc4G3MwV+S/ltw4hmQsin7hUxRusstG0yTlWpvxfqwVKsm3QX8Mxsvt0nwj
SNFXKpy06x/18mWCpC1rBcl0ULYKhXvymrJAaMus4BldkkEYtNnt5i22jY+GCPKp
xVjbRfgNdGKF6AzMGj4oLjD1ikdMxhNPe1yNDTnDbHWnZoA+tl1WHUWbqjqKXwVT
U3YRk6mgkNPkS5ZLawp1O3pqHPr83vOd+cUQ8MCVDj1dyp3DnEEdDHsOdHZNqhng
vH/WFCz2tXAdgjSxHwrLQJuVP3u1bhij0ByMOMrzY3c2TZ3C9fk6zhNphasSHgni
IKkvl0NHKjXgcz2RholOYqSX3zeIesrOunhKfgiGg7EfjVTof7YKhV0msfiKBEil
h3rcgHkkc8pP4AOaVoEFCoeSp0ad5P+RWWTl26fmfQCgqn0YS5ZSkIVB7eihwK5p
7SU3s8E2cg1juE5bU3Fct74gQt8VnWBYdY/ceM3RbEdvsdJdU+iSTZQD7Y/OJ0pc
`protect END_PROTECTED
