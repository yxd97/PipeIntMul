`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OD5oGxoRjTIlYmr0KDzNzEtrAqfYWnuDoz7QdHtzX38AlIyYSBkdDJ7aZzJXMctl
ugPAU7PtlBJud2g36QRmSTPFVkO0xjbT3dfM3Z3POYlpp4nDJOtRIkLF6aIm7vOO
I3VIrrdnkSQUchYmm/Msu1WcWlRfGjJMuhrLZEkYWodMysvNQ6cWVuLEZLuAm9iW
QgViefke4jBGDX4GKefBFJFk1Yph+WSEXg5SljwSf2kFpZuU745YDH5fwQMbLiwH
XK0GgrSO6YrD9JcvU0h4zz4sT/QXmmHovSPfSET6yjlWxA35i2cgF8sjMAsndJVC
zX4jNcQ1qSjrDvZsZDGAY0vZMPr7NTFvRJiFaTBl1bJ/zfbh+PwJeVrG4UBDnDea
PiqJl/6dYJ/ktJzAwq+GGKvlvumDYzyEhvS6U81RlgHQ0jUa5VI9ToUGtXRDgq2S
eo6XhyQZ9YsX3OAkQoVIZGqkkgnHFnpAQxLNquG2mGrrbHZqIsCEUdyrgQXqZ4r4
A1kImBUnRcCcRXKy+2AuiSU/Ds9YgXr4UvwRNavoJWP7Ck/bqivrCxHK3s3f2UU7
P4Y8uTB1tINLN8j20+/PTfvYZlTgBvUTk2Tc9GkbCJObr3x0zDyNxW9hdPF+GGBK
7BYFuVHvDIeXXin2EdOhXSIDSTH0HFwpcq/2//Fy+HSeDlpzzzRNyoL7kA6iJMlA
7Zkvi/gZH7tbyyNRqwl75gDJlW1Zc06Wx/hmMyo5gy57dLVBjwpRQvZak+8jz+PR
WUYxFLyK6sxkqOA1oDPCYb9gBepxNbbnneP3/d2Zxqqn4MnbeiQE31eLZxn9kdJ+
7XeofGiqE/G0rmS2mlrdLqMEF/Yo2FvB0jLLtFh86WxuqdwdYQXD0aov5eVhDEhk
4Hqnwzk6yrYVo8SmuDHfIGZ4hkxblNKvqxyurEzysWdy7BVJFGBuS+WniBfBl8EP
0enZ6IE0LqeEJfeCQ+wo7Aojj/dO43GdZT4RtNw1XDztwO81Gdo0erP15RdmnLRW
Z5wBzMr23881JqPJRdn05+f2JbXgCr8VrjP8mZezzqnFXSmhEbiOOkZ/YlIuvf+K
3s/I30C2mKH4IbnNgJqmOT4qPepT5kfzQPBHD2ebgEQKuZKkN6JJWP6q2LfqlBES
`protect END_PROTECTED
