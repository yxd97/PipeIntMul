`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PP34YwkEXl28Af7h8C9eij8zvz55dS8t9N9evbYYKRNpVbe/Y7f8rbmblCmhWcTk
HoSL1xPnBPMTVHB5MzDrjksqzrxCa6zV+QHa3pjLoxQUW6RSJq3ujMnmPxYY2wBB
LAhpKpMvUml7CTPhAP8vVchh5ZF9xvcJSj6p2GVK/V2GmOTzcd17Tp0Hecf6tzDO
sdbXdI73EdS44M8LtgrBtDKLQ4lE7caLbk+31iFWfWLT0orJl4B9UfUvPgRdwPKs
6BJRSWU/+ebLLV8WglJng47Vv3QgtPP9Vf04TCnCRjqMXgge2XkELhdwCPgqqfV4
qcmGTcsRQ/XsqLfPWPa752VzZxF/eBLoPv+T4krMnKqvbAsjxm36ufpxj4vTfoNX
WY6T5JMdul35r8r/nAd5eA==
`protect END_PROTECTED
