`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B71PgPpLLCsAQuwhzi9Mnv+mn9eK0DxhEpWau9vhBrW9QdPcTydguDRMPj6pONmQ
KXRh3e3unuPV8DVZYZCBBwebuW2oBk1C/9RulhYxHWwIws+qR17KP0djHUJoVAsK
WWwZOYzBbvsCisgCOAp3K/uMvQCcfMqqgPmHxKSpVAGqxXElGTvwkf54N7jEoqom
0osUwR1vzrK2eOFCH6tSWqvM+YQSKINR5GtJvFhPOoZ0lswYdOZjs8ta8ODQrZ2J
YCiHEx7KNvYHHnich//V9rgqNdLtCfIIh7LqTPfWL/6wexRWrKtw97BUXBJEnAta
`protect END_PROTECTED
