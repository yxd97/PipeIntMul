`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6W57twwtuiaaHnbZs0G2tG6vJkqUZbw2sS1abiDnfaYj/ip3gZkF0Qv+nJlIy7QH
l0p0fvRO2woktHaqde6wc3Gu0cddVkFHEaSPuGYJMJ9RwiuoMqNSZXSO+2HuZBaw
evu5M9CjT/t2DzP47vgWtdFElpw+fYDt25fgerztPJotuwnfIJE0qiNsuRIwdgOR
bkhInMW4zwxSQibX2ChC24ak+xKr/TUOZEhpNlznORRNy8cafnhVI+SW2IzasuiS
5YXnoDoDvvQ9giba29RmrpguMJ2ADD6hg8Ra+8iu0OM=
`protect END_PROTECTED
