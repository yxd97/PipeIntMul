`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HH/fdCtmJVPTKJMWHeqwfAVdC96o8+qH3P6smAVxDDYMhX6rg/Ry7sOhWTypwrFa
y919yYbzK6vaxg19I0C6OQ4zZZHWCb84dL+kI1qRl0UKOJGgIZVpH65zvCy1OaT8
p3+v6RXs6nEL9CkD/ZQj2QUKe5foQtporn8hdmd8ZjWthv+yqqAIYZbtE3h28nwS
c2sG9CqhgPJvJjXMXgfoXkdI8dMNCp3jNNdRTtzpYZbJhC6N00Qrt/seYRJrfUls
MgV58rs16abOml4CAOhkxN+F8zvlqzFsXyW0Iy6y4pEz6I3sNrz4ntisyMK/LGJj
Mb9y3lZIFfCl+zUjLeqIa67wdgEgacDG23d+PkLLtolOuxf+md8hHABBJCKdCLAH
3GjWlu8NCJ8hXRzOWSvT0w==
`protect END_PROTECTED
