`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DpZABTJ1FA++3JXV3CxOgr9duttREo2bQAj1B+uY5MttSDfqxEIeYGRULDeVi8rr
IwwjxdV3emp1ufr1MU9NNEqnIKcv17ePTIlBr/uKYHkIIybTqSZ2md5OVl9u+ezt
VNk5x03CntQFIJqXZYWkko30GqNtyAEKuGSI40wp1LIQkNSTUh2UKB1xeiQbsi+z
IRo5GM/2uFYVam8uP95ymV9VJ1i1lWDivhT4GOGseVwX1jV4ZLHb+Q+V6cAynpaD
8P/aPlJ8Ec+5d9/2bszsdWKPip8VKRW8IvtdYGDwG38=
`protect END_PROTECTED
