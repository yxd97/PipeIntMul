`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKYYN5sFoPT4lgNszv4wcOQFmJYL52H5YmJq2cGfb5fQdzrwo1q4dNVEewDpGxre
GuOFdZ/wkkMXzL8AndJZ9Z9eBFkaJs3Xw9x/jcfEvucwZ4K0Lezqmw9sIgmOTSvS
T3Wdfdm6GxaWRDv9fatf0J+0IHOZZESsre92bWAal+du8KaOWvNYsTPXscfLODr+
XnnPq2uhewLXxPZwX2NGWs9el1hkkivNETmRE42R6j5Vj7dpIFZD7F/qa44y1K4s
R66MYaEeCl3c1IHNWtBAjBMI25R4y9pWvonb6HhZWzwuVBqdq0und8JgtEtza7bN
BwOimQ9568QIYB9G9Zx1DuJ7bxH0HxSo69UDeZrRW9SdRf/M33zvzfjcAnV+hSlE
9T8LRwDnCtssB1duhvkX0LdJpCfxInUt5/x0q8n8Kys=
`protect END_PROTECTED
