`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZ2TpIbyfkusUVGtZ9nXpmzaL75L5DcN/znX0gl104Eq1T2r33RF1lQ2EvzxX5Gr
3cCs78QPJVrtc41idxrGEAK2aa3ZnkQ0sky3sv228n4lx0tA293CIXHL7w+asd4/
c1SqxyJccCg0jiROU9g372nV8CjjrT/L6FEPbP2rfeLIi5ZLHugwUU2+upbUoXXw
JHqN8GPc9Tv3otuCdTiPZBC0pEX+gB/DXqHh8f1Kqk8K/GQzB88Mf63lhHUjL/Ec
jPaVge5WeafIq0oEijQanJCbOzbncs9JsCO0GOeSPG2Q+LyvTUAlTOQZgA2kE6J3
vK2KPk7u4P6qMWXVLsfgxBBbaBhAd8noq3GtdchvPs5T+5ZBV3X7L9NotMmfbehp
oH4s5KdoUFhCiWiklctgcmVYfz7QQYND9cJs6fbFjd832z/NqtpQao0aoZv4fTAh
xzcdR3HzQfsEtlEEEec7ogBhRcJscZ+Px+azj7rqXTFKDWbT7h+x3ijHfhUoS8AW
c4Z+VTYG40ZTNfKQRSxUazdbTl9Iy/VEmRi1lvn3A6uDe/sHm2sC+FRzUaVVsHo+
+X1JwJPqc5S6+dMGtwOsTcqhvxxkjp966lfDCT+gmrYgIdxuPjte1mVnlMxxR+nK
7nKRB4w7spAwASDhSIYLPGb3lJm2nM7bfD11/1CTiVsmXkAtd0m7RvUcX9SQcZsF
dGWL4RDQmSQQo6rgUVeFCXCzJfb/Ud6qngUL6gFCyUuJEo5yp+edOLzsm9Q1AlCi
FNx8WvLJX+wxHmKKed9FiMkibVt/RKdF4DZfeW1+lu6nbHbYE+h2Q0Kgv5TG4pzX
TnAR/Q1C+DPZuDj259xxdFh54fWn/d1kx00qD7H1tZM=
`protect END_PROTECTED
