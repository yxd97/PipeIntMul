`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f/y7eQHWvry9nV/QeZMSH7hKYFtTLNln8QlYEzCQZUDm4JsFxaa5VUWMwzv08YSo
zdoZrHs4XyTiv7M0AGRAzB1X8XlVVaGo9gt/iCJvCtZmJR1qJfxZXwUfAy+6uORw
O/o+8JbmcGEPDV7tfjFcdwT+O6H4rZDx56cZ3KZu8kLDefSGhhZhGPmmIxAKEOkH
iRMG3/FbH/ZiRHfa9+RkmpyqKZdMD2bO2H/HAGS8D9MfOahe6ZHsX76T35mMFYGj
3VtaP6Owfx6sNnG/gZivNOhK7xv+BkmgjEDeHAms8F5rKTzV9OM2PDtMc9b125om
z/oWyDfOhjt8zQwBtZYguPfVKo2DD0Fyk3w4ijo5ARCRKoIqGAcLlDKIs3mjwEjh
f5Su/QbVMj3lFgTbjKzeEqwv7wK404IkZRQ0SYwKvxunuZkg8Xb93ND+5HkVaqhc
iFMDfA5Cx4puZSiT3tegS0NbAG+uaDxZg8jOqLCbbWnTv29x2+82nHVuI1dLuLcW
DozO7AhGODYdzuxfyEyRJaFTVXTse9mEBK4TaDn8p3mrfkugkrhURQ9fUtJwJBLt
EBs6SPT0NjatFn5OB6XUQaI3NMOW5K+OUasBGYEHwHPsePEfCEKDMYWmFoNdHOnZ
zBrIJGCQwzBeIc2/l/so/Q==
`protect END_PROTECTED
