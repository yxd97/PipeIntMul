`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gvyofRD01+rUOHqldMlDjgHytVly3QlxgzhHIR5CB0DJPo6nmQMQ6JqA4jsFTtxG
t1fShLj1pLM+UQKj6mx3+lry+yQ0iOIf+4ok0DYUoT3l4+POlCiQGBxiwdHHU2vv
KcEwETmmo6pU17RhMv/pdmVi24ayufAzwtESL/bQv7ovtntflOZXPMM/b5u9JsMT
A/voiJZP7BPrI8b1xBVeerA3ErneiBcIkMUPl1j9s8VDG27upIEdavBCtc0aZoH4
uDXjqR7PyhVE1LL2RlBZmTge5MruvvmhMGIImm/t27jxUsnRI/u8Vu/2k0LVYdYp
THRMr+KkFxvyEDgurF3RuW/5G/pM11mBl3i77vgaezIfq53q9ybXvpgilMLwFiJe
Zs/dq4kzjYa6Q6iJ/b6eRA==
`protect END_PROTECTED
