`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfsZhY3RI7YIfBFHBpzdUOzokuO6bbdJrHFzKHxejiBfmakc2S2Ko4S5UNrjEl1/
9Req62U1es6xLh05qjZrQ8OUv2Rz8Gtyg0NJvK0gHZsPb+o8U+EOhQOVkLQ0qwS8
VJrSSHufVxyENqb5GKXQUSfcsgGV9tqvzrFyySnfWrFqLgP2Z+csQTcva2ANSEIM
4yd5X3yoKFw17YRqqNDnoDzjoonmabf+qvNBWNl3LsW9Dcp7r14brhVDFPmrSVMT
JBAHEPw17BbjoBY1zNQ01XSiQz+plir2uKQ7RQWZ77VAHk60e7UUwp6/l12LnGba
++eFb1EHcyQKzmDZh/qaLaV3y4xQ21QSZJICExn7TwZNp4nxEW9nBEKrQusNp/sI
+wU2Hx8XCS0iqJCNtkPoxTFeaQoJ8JqpV8DUyxIx90jTMsqktBgNegyqPFFlsVRN
umohYeLha8f6ZpVNzuW3zQ==
`protect END_PROTECTED
