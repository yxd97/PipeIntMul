`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
csy8Akv7+GM2chcFYdkruh9uhuQB9P+WJgMgfeu75y++qxS2XA5IMcZApb+y8lC8
IxDSUn8L/zqHs2C84JkVi6+2MOmeFbcKX/itkw1q/02UqaWvaX7NUa7JfnD29qML
IHf/wrCgJRx+UjGJVwiYJ1v+G0WxND+8Jdsu5GDSKxVH8oQmcvq1Wxx4F2mLGt83
zFBlG00geTAYlMIvqyfscsfGA0d0yg2hHVv0MtsZgPkWYjSwiRlfmfu/BMq62Gqf
VWK6ZOOUKRMmIGl4kMDb1OE5sZxf48lKdPwXXlY79qFgUsaE1XqmjqmWr0LIh+Li
5pVdXvg0KkxdZUFDfEnv6YiVDf2PLiNz3SCI8R2W7zw8s74pV8DM64NC8HeS4Qwo
Supc4OA3LSCJ5PFjyZTVoTJU0t8nNdGruPTXsvTd3LebYjB+KyX/FYOW8RvxkGPS
KK10+cUFizAGQFd0H2kIHc5y7AibGUHqUAoWMJ9Q5Y9gmQWHP6BQyMRJfY+J2Tu2
zS2N3Wp+qwwn7gthHA/bvSuWD6IUCtR0ijhhXNHwZMrIQNS5Rf4LREpAv9e22gWJ
tePyxks7fh2zz0T2zDx31mGVfQCpnE0deWZfJqZFiHZq207/Y9uQ0kJfXBb32hzV
AQT6qemqDYrdTZopGHsTWQtKm7xfNYjVPZcXjFNylTRd5sHuwZsriEaxPEkeI8zl
Vcg7LVqw03udIsJXEFgNTfUsDw2In6+oGfow7PFBV0P4MzfIyMAS2rzGbbC5Fpjv
spWVjwVch3jzKKOdpJx7bDuldGl2f5/X9jlVhiOtDfYnleqNSiwRC6QMd85Gf4AU
EfvFZJ62BQS7W7ir/pQs+PzQwgw+1iruntFagn9++1PGBU2LDl53fdSn/2zObXST
lzMNMJvXG7zP0bGUmMOf/72KECBsjp5JwDfvFJdE4gBb5aYr0MTqXQhmC8a9HbSh
tAbSaUXVvf3ZUKDpvTbKY5S79gbznRqJr9X7M+5TclNyATAMTRobNaYU42qt4yF8
b2Duat3KDkp5YFrkFX9XIh6Tn82uTp8seCg0o/EfgB0L4fbpjR40AdNEi8uL8J9Z
JKVBuooKpIt0NLDHicjzPjxxdUmH2j1eHJWBHRXlJOhAfPFbMe1KwhuSVyFYZlmn
Wvd+4fIwfyt0wlaAO6Nmc2TgsON/+V2cry5+Jxp5yLPZrnvUghTFPHN9yxLCbaMq
PFmwFUSqZvDJECtm7zPjfUTM7pc2pagwoXJq2VIkQbFStW3ieeXP+TvDZrsUjw50
38GZCBPfVoWNSSwP01WP8fT07GnIEZ9n/bhdFN9WskN+3Y5OZjwdUgV6UMTuC7pt
cP1eoo27C1pK8ODSzkd60TZWvmgPi3ZTOXajDkdXWLLolDN4YFExRXz9ov8XUI75
qq7fHAOpnJvZQWMVTfe6q8bH3cj+wyS3i/dzVxY+OyKDfIDe7gqZliTVU5HvzB+L
tK6bYRo3euHSt24T8nXmNf+RxY8x1ynNwTXrwOuLNOT9Bhg7zIZaboVEfpNDjDKg
LbaAFKl3ivy+F5Qq/eRPURlmzp2ZecANlWVBdYArDKbCTctA8cJPazY81gHEyOV8
rE3bKUw5hME0i9oD2DmZLkVjH88xYaMLFxJxgXofAcycQVt2EzleEKYz3ofUNUOu
ktTftwdq3z4hcecMKUDpK1+t1ze5xzsELdKqKTqK4esoyOYiewJMnzV5vDvJCj/j
8fvz3PYdyKpZ6Eqw1wsW4guDNaefb/zPTHQaeqYWkgFvXEw88q9eEanQBbP4HaZ4
qmvTeSL6ZikqmHxQclT2sldKFvU+dK52Nnzdsw8nlE580jFXFWoXiKctTtlp42Fn
4TOKZ5dU+D42C6GeMuN2RXqAiYv1cnKdfIa3hzNClIztjhXXSIoiSINiXrLEYdXN
ZV1GiGjmJcbEFYIQwbqRwZngy3rolv12KxKPJxLOr4RniQfYzywmDfOv1JcWjam7
KEa9eg3FUwcvlJO8iagNoR7TrVxfIyXLrU/z7CyQHXpxb1PHaMH9PisnOZdbsgL5
V14WDVP27EDpJiFRsgHpewI5cEPjI8mEE8+t9cps026D0dRl3eVspj7rsJPQcaUy
W0W7g2u4zIwxgUXZ2Pkr3Te4HBm0m6iVIQFaIcVAanOp/glaJDFdQ1UuUEPDTL85
Brs5m/769QVo7NYnYM47Ip4UumDIpN49YmsQ9J8/TBqq3XKlQ1aLQ7F0q3PPCNpJ
asp6oHnmn+KpO+oaUu9o7uSL9hxdfo2twQe1YaZK1JirN/oAuvgEDOMpSE9guPim
z3/qBJgRy5MmHkukHbLNHy3VwqTGYcK++wBRn2OmZfELnYhJMDNFi0+H/edkXvF0
ofivaVcKCoNQHyKK62f18+OV+E0ookLPcfz9Y0uxNNDRPJNF6s4uIG8WpFUfLyYU
lk7Tmq90jt6t4FSiP80UQGAz8ZZqSgiQZveW+E6RuYMhndpeiKYmd0LOzzMNmmGD
alTmrHSctgCM8c6F/bL3aY46WR6CaYi8de2VYbMLUMhbzM24iNSayCKVxLom/qFP
4mREa+BxgAo6AArG10+gg7xDPZMUILFg871yse86KOxMN0fnK4a60Zd1twDjieMT
gZAwJg5AOy+HD7jHsnyNOH22sfD6IDJKoazfRfw0+8sTnVEM5Ydm3AYzxO4W/t8c
+U21cmgIyZrWkyfzdrabpmj/0ow4EzazsI6J7cGvIfvbfl8bKYcOcGXqUINMMR8/
`protect END_PROTECTED
