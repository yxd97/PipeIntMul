`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOySKDIzeOjWsbLV/XBBZYJb8xm4D8eVwTzQXdYXsr1YImg5WUSA7T6hWWiQe4vB
voGy8qzv3lphMRgX94ZKbV6swTPyDOI5k7Mfor1v3TBbW9RBFA9V/f8yHQ2jC6Mz
29jX2XJiIThsZ+MJfbi+aJdzTiAMHNFJfLuq3AOo8lC11qX6llMKk8pWKR2GH68M
vGJGvJJxPT7kFL4giVVMoRowONR7z7CbyeFLsbET51KKR0xsZRQdraYUTr10ojqp
Qk+sBnwQOJW41rzzHIlukHgC78DUqiJYQXqgCFFP2oV2W5qoAzP9iua5VWxlXWDv
bmJ/q8dWWy963d5K/s5xG+XWZXFFuPuosB6jj1RkO1Om29IVs/bjHSzA9KZ3vfe5
3k64tYroFCz/YcmJTHyjbYsQkko1GFArI+V/bgwTnb2limbfqaL5I43DqRCJA3oq
CjfP+hekRyaRumYd31iFuC3ONMqlwLnynTcmmetC6JZpTIBd5P8WoxW4dbtLDgCF
+pflDKzzTjxQRQNTGmOo03HdGFr80DQ2cvr3UjtEiTPH7d72gjF2TP0IHSPFFD16
7uS++dYxNa6hdfywtePAZA7ZNO5wqSvEHN89VmMRM8heg5jJ65e0X9dQAmJAO9iG
TCDT7zfdD6A9eGAZTxruBS/FrQ98XyIjtIPQGT1tqeOfgcyJV1rsvPGRbEvfv/ug
/rNeYJ5nY9YAIlPh/jrfVa53JpKeZOn+/QesCbqV4v20K2AJYxL/NFb8GTBzScSy
VnUaetsQWIUk6CD/pntsqqylfDqySRx7LLR17IHDMC3kuFmvYz+BHlBZN5yyPHDE
QgZ6Ubm+LDepHuXSZavgEA==
`protect END_PROTECTED
