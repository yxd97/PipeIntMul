`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gg4VmstkPEI3j21yRcFWPqx1W8KsW1gj1UdXQDC9nYAKNZh8qFUQ9s9KwXHmtTlv
d+A9XLP6/6l5ProPnLP6ykWZjH2LonL3KjqB1jNmZiAiRavIV6UFrB10KMXKXrss
qT4TgqB3WGzeRQa++4QVEcux6F5sX88m3tla5iVR92IBXebpK7Cp5nOVYB9NQCa5
iSM52kr2gfDkAQ0imvRFu9wntq4hDQHlvRjpqitB+PerVtSMGzzpzxQdRbS1OvOb
6o/pPcVq1hdyjtUI13G1sJm84wUaeOkJjxYg7l3LBO81CG5w6AtvZnO50bWtwMCV
vcpchfPGcWKOIQeJSLeLOjKRx45UheqzmdrFHab74qZTohTyhnzF0Bg4qAakDlku
TUuyMvq1z5HXDMtqkA60LvY4WAd99j0hagMqoW0f9YX2KiSnyu6ygo0bVXG29UbH
8THtjGKCu5zJLoCnEMZmltRP5q2R+IguDXoqn4nO+b09RRdG0YoLdqhaazDMtdNM
`protect END_PROTECTED
