`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIjrXdEqaCXppfLkVFkg608CqPo44ZwbuSn8NbitkX07NVctu/fX+CqrXadTPtff
fgY3z8CLXIMB5r90ZVGki2W9bQ59p4+Q7D5BbscyKDowg5oeLKDTzy6meZtSwDAJ
ljQt7T/TDc9mGGHip1D0JM3naG5u4vDvBhuGYctU2gGl92TSorwP2WaLShBm1cx3
9X5Y3ijVT0fe/qILYF3kojDVZQ6NcMDD8WLeAanh26Z2WEJHy4cCZw4sIcXmEwmy
aqHoBBoRr6iW6Eu+xXrmPhfrur824uxWzZvxIVOsdDV65MxHvKFztze5MGWHfi8v
8mLSSNGNnOdq7cv+8j7oCUEgOuUtsQtkhXBSSOYvsSf94UHyp7b6Qf7g2PNEl8MW
ZGxdLf8d1AwNLNOSXyXvfCf8gSetG1EjiZhVE5Sx/H1lphgLBAsKk/q+lOtQn+ji
XWZYSfJQ0DzOgcHRpenuhHM2xiUQ7IZrysv+ET4hOl/Qh11bMIsKGo+FpjqhpOai
d99OU06MuL7n8Z+WRpn4nSh+yRr8hERzZXNvRdoUglFnwLTdoC++wC9Nn4trqdz2
EjMaxvfyk5roNlErj9A5pM7TDDmrofHJnPwfkv7cud4=
`protect END_PROTECTED
