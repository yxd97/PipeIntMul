`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SVksXrtrUduQ+hCpkNtNLsXm5ji3yOAsrnHYDE4i1Lpgfti6/mw0zV7wHD0QOfGr
YCT5rowD+ywJJLcMuS/XIXDui6rT7DPiiDyA22SiRdov4SZWDDWrnCnj+EC7DB0i
/oehXbovaDbFbzCr8CRWeM+QBxm8ML28VlulUTNwRPGerd5VzlF6vCKgkilj4wcg
NXUoh2tLYPfXxBRsfCe2X8/9Qugfy28nTzUC0ukmZGOkXCh3YGIt/uDM868yHGaE
60zCLnAi+q0AFDw/qGY7BWfDT69zKDCLptRInu/Z4fiI4sinMQbo+tgLLk7hHpNa
Gnon2dcf2sTIf05xifU3M8ylhqLPjoYoTZ+YpRWKmqyiPbZNMGOP/8H9ADS0bqh4
Xs0lM3nTvmpyUjRTFTveUoFZZA0fwFU/w8HEta04jJUu/VUGjZoj0hGVJBSnC/C3
UF3ZxbttS9eFum6R+GMEabebCwQEbzJzc77RnrcrtvSmqLvPeVsulj+Aa9OactIN
`protect END_PROTECTED
