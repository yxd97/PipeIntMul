`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLNheg49KvdETRLnHEWwgsW1gVDga1P8EmJVqxm3MqcN8lBoXM7ixg/v5Uup/iEx
jVuWuFSiWSBvKbYm3J7TfGBledMDYpLvQZw/qNlXJg+QCqnxmLOXxQwuh8NzBd+C
gW3CWeDkDsyqWH4Eo6kB4kJejHOyIGRfMPmIVDRq1wGEpa/GWjUlz3ovjW021iKY
35/2YlvQM2GwPKfqcLO93u0G72dyZHvyoUykIZMeVkGSavwkZzSHWJJ7CEp0tNFA
iClcJwcycXbMbzXW3GLWfm7MX6RhFXGX3WKQY9wLq8J3R+MijjTDPvONCYpKsfUZ
SC7C/TiwkjmSo0gKe8tPIJ9IeaoHUba4SXvGj4f3BhAU+EPxUOly2tiCqRXeAtFU
S1QY0ATvZ1rx/5jQZ5E1elHLDA1f29CyIdMFgNEgrQ8=
`protect END_PROTECTED
