`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OB3wFn2K/ydrZOBddajVakZy6k8cTH+vrjbS6vjbgo3gL2qpbGSqRAHZy9mwxt9o
NGRpyJR4dswEVRUOCDgDkwo/ING9YqyzEe44t1XCM1SN03l/QndesphJdGAi8YTT
b+KK+hOUdDgqdpb8FVUDH2ot4TnAW5Z+A39QGt7k3TEpcheDpM9umAWNDSueBsIq
W+7qCdfBmDn7qq1gCdkh9hP942BnLpAeyl5JFIz4UsYmIzOzEuFntmGV4w8jjWSV
w6gudaRW93qdwhdXNFyekBRT7qvEnH/96ceoXbmvxmcicf3tEiZK+/irkpgynXLa
djP7FsUivPWFWW3L1S88/5ionbZJQZ0qNx6vJwSmr55yL/xNCEKOxjqoKVw9fE0O
M4P7KJhUNAfC7BVomQncYw==
`protect END_PROTECTED
