`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5gBlYy5i4vYwLptAZbkfd/mGfg3evdTKpfgwuQ+j/gCo2oU8d9Ni3am5uJglFXbq
iqjYRATlCwcowhmIrZrr9OyRFcZXEHWSa0SR2QMSXBpfrc0YJbwT6DawkfumkVDK
hp07VyYUA/X0PkO+b63k3OLnYe8oot4utuq1etktod7RDrpMAqe5u7SqpHHmnfxw
W61SW50ReP5fCNFGTulGdvf3McqF7iylRQgPZ8FEjC+0fN7V5V7g6ENu6PMKHnlc
YAdZxiFn1UO+ZEPZG90CHumqGn6BgOAoYYKrLLFz3VaFjDimHcQM3NXs9CCEbtNw
mBAM9JQNrEEcezVdxDNBnw==
`protect END_PROTECTED
