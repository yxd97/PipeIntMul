`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9LVSfvCoD41Ti70Z+wvUEBhZeIQZiWwnHwFA2WMfVn5PZmyG8akBvmBdjrMvATbM
1+TAKepqPVLaLxCBUHywEK8U5w6D+PMDHbhYjP19gVrvMMTC8iwqhLC0vUiaIAE6
WgtQRUW7WzGGMl1lZUDZzdddDywI33HckbkD1q9E4rh8/cykI6CM71pFh1BEW9pT
ijLbk0MPVzhWMcp3iHwuyMO7rf0Xv2uc8VpeIBcf4VKEIlrOJ1lgESUoHDrqdgRl
FL5Er6v+CcirEiqDCHjqwcXk2LcY/EraY0qhclpjxbtm50P/5BwQGgnkYCZVPxRy
ILG/k3qJDOE/aWkub9sw1QTDa6swYXr9CT3P83JJ0IbVNcOBH/qcmBtHnW0fyW5t
p+S+phk9dD4ZJN2JRtv7KASRdWXrKJYRo4sxhfULhrGLT1ktmxzMu/h3V8YLDaPi
JPmeLcrjGiwdj+sLmPNv04hge2AySp/es/CBQf+3aH2dAnNQ63AGWmuIhcIOXU89
woa0zpMsstVGuWnB/wMMC2/aOciRH+a0RLm0U0DYWxNUUOtHpQrh643pClTmiHP5
O335iAlrf1N7+1ftwKMW2AoOr8Ky/EobCXqUjjTmuPrkQqooFKJoqtKtQGqeV42i
Diy/gVDCOxjlSXAArHH7vg==
`protect END_PROTECTED
