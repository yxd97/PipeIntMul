`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7N9P6Rh7jgDo+87694ZmAc6r4U3J1uBIFDenLsPsXK+ZUUsn7vzsK6QwzKxMU8mG
a0817CV4Ak4DigsZmGot7BeZVKTzOkChu1dVzf0WkK26PKu2upshmcE803QLsgmw
RtTVenu4PDLgb+UBDa+XEgDAyCzrfWfjzvEatVjFC4pYpCQiUbQM9xZRefA8IqhE
Aen8KN0hp3sNVcm5h0Rx0GKKRIkhlkgx6k6Eo0mq1QgVbWghn62172WsSxWSudlb
bYsaCjAhJkKAndjMV0d/BE5XOc/cD/Exa7883jmCIE6M3cA9nhPERtn2tRWtdIhH
xmFOoqPMmzbTEalNMKPa5+YgGtS5628P8z4crnGafrRF7hXuzjMWWN1UojM6sg7Q
2TVrK9pKC5bx2MBFhaDHitFjG/08EeY9VZ5XOtQhvMcrXy/aDCnssSyD8MnMtF9j
6ApNIxq+pO4uNLLyRFY3oJs5Q6SavBcdFtXsubuEBc87beYhmyX15luTr/nZ/aj7
a7q6MzsG2ScrSFLCyQIjl6xI5yt33KdYrn+vmevksQQ1pwSTaSYEQx7+zJ0CYwXp
L5aTynfXZ2CgyXF8jH7AC16rc1Qhs89w388iu0H2unWHEKVGbeviRPFYlDWEFF+E
uwIMWoo3NE84Mab11305mQ==
`protect END_PROTECTED
