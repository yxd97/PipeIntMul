`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HA/kNbsqObBpDADLBJ2szv0eOIzI/+KY/CVPstLLu0+WYcPd/tPAf9NePP1Xq3jD
19B64skaydGUhtI2mXghkTpO3xvr/RBeO7Iyu9cVcaQMiVu6hyUQZnVlUhRw9z/t
QbqPr5QEgLQeaUwN3oqRKV1o/bbLLjq7TenB6u2tI91rJMWVrLtd56FwXBjyCrAP
TJqj8J1Vt7Y5mFyzbP8G6ch2uXXdfOfCkz+tFJtFO89A6DIBwfEIaLXmp2iMmlFH
FJ8xJDT25qvDpNMew3C4ibQbiSWSBQM1OrpAItQZjgRQ+yIfRSo1SxgVQj/UgU1s
Dez5jquVWqo7IQwcKb2VDKMUcZIW8/t0mLhNsFmKd5ipLDYcjuEu1m+8/UVA2mBV
4SOf+s1cAtf7Tk4smSOyBEVPo9/DTyhDe8tY3a+6NcMdCPqZvBRecSgNIJ151fdO
7xJQ7MwNuIY03KyIwSpdMrGLz1KqWit9avMLqw7E7IqLMtGQ4n5FaidbSoId27dM
AUxMIkkQqSgpoRddn7S1a9W7XMMDU6PjY+XAgD2PAmwrygpY5ltpa3b4P1eFGQOt
QX4UEX34yGtf5EjFe2NlyRYZCc3Q7hxfxppr6H496k9HLus2Hk27N3BzkJmVNd07
myS9k7/IXmf52I8nar0GyIff/4KxoKMXf/ZtaNwCYn4FyF4yiTKWkQkAd3UWBVTG
khTwyMP4pEWfOZz77I5jKhj3noeIq2ijCd/bKNGlYI4Qw2BH+O8kZ+AUZ8dlJvIn
fRIMtY8C6zDKDWe5kSGJlNHSTeIA9OPdXr8sjCx4A15L1XiHCRRo+3nB2CK1w2ze
fyjmc9hF2iiWwlGiHl9/md6lCffnl+1JXOJ6Bk6/xo8eFArCivKJOvrAnjksodmN
9i6jAwx1l43xuZgTGS/T2qWi1bvmg1hxMeSxZEkuRb6fc1VSD2bCHk4LvmlxkjP4
72MVpS/l9EgPtZT+/DQkryUlSF1vJrVc3oX8K2+mCQal8KwwPfG55xVxUf4ssh1p
9EJEOpHXi4aslvzDhlj9htQ5PIkefwgXhf2hySq8wY3P6hEk7ZVQh1dDbSSKVNN4
Ll5wjM202wEBUO1Z8YT+UNGVDazSZLfrbHXWzsOXVQ30wTTjc22wcw6R5WjDB37S
pG4zqQrbVFMVxwWwzbpui9R0Q4Gv41nZ5/ZJIQuUZ+I2a8XzYiktEfBTlZLcixdk
6KeoaBWuzlqxCmVJTOTiV2zOFRuEOlMx/y07TCGz2Kpo6XcNcnJjP3xGJ/yJmIS0
+c7qU8rDerh8XqTozazQfdLluBXOg2I7IH1TFQf/K4NGvIPRT3SuXLj1maSBpNbg
lAmFime4Yh17KP/0W5c9VzAOrsWhtOG7Xf5NOL/bhDoxWpNDXqckFwFrtiZNpPDF
a8pWTPZtxVngxM1ulhs+SEE/kcEhFahfU1ta+Tpjs2aSV1drD89Gi9plLCwsx6nm
6fMstzJBW1dUUpUH6iWrpKGt4xDx/yFcszQQgV9Hm6zlwyWxMprWNBOLDEIvv2vd
wPooihPMoCbOWLm3d1pbaxMSik/S9k6DS0JHu2oPEiIXT5nxFNKh7PiSFY8+a9kx
PLnIHnrMhH09B/5LPv5Bvg/iM6PayyjZlNtdVfIEKgENthCxlyVffryTlXrpy7G1
d8ZDlhvVDDigTA+BKnpF32TD+2rAzszZPL0sSyQzsNUjjQGKJGnm2PAU7q5aodOT
oaogabfqF2w8W5gI/r9g1BSsbVuaTMVyCf9OjNAYpQL6kz2L+si17R0AZM8IP4Gq
vrOhlCTD4Y76hmYpZ15C2f4lWkChC1FqhF9CXENEsOkVgpmA6JyCz8KyOuIDKs22
2c+OunRpsYylqTxc2vPP+0UjY+q11YomnPRFyTeL3q1/loq4tBgEoEqe/BdrebC3
rNpF8r/qW+HeQ/onvAdYqIxCMIxxGh5Mg++VEJwMzTaucvI8K8E3UbEeX85WUZVu
mGJbewihPF5il+kolsoE5WkkgWOFlPSMPOTKkNkyC4rTspH7RdGGRMnVjIzGtdXe
XEVuQ77klRoKv8v6P7P60AjrstiRmoPzUnyf6kyDNlgs/8x+gxX9l371vyw3l9kK
KwB0qpMZya3KxIjJI+Ag5d2iY35VPgiVQXJ/Y0v7n+Khe3CdWSL2qaMjRQ/7cFre
PKbnHHaF48Kf6z34UwZvWb0Ym/lOR1tviTumfrZ0Ze0j9YQApXne28f0tN8EKLcW
38r1P1BLse3Hdwun4O3UxDJ2kiBSOgtpThV6QcZ5yXYc/zo4WMh0jZp9QO+rNvS/
/1XxRa5t1qPCQdVIgacwt9+2VR/JsTbWomhczojrcmgWCdKFJTXas0I4QSV2HuIu
O9nLhFPYmfn9Vwcsy+WeBsg4hDoYnf69A7zFUdKoSvvcjzj235mBje0kGzBVgAQi
c8R69YP+fTGnuuSXRdiOHmjLVLAOrXRety/H/WxpasbRhCrL69zgKFWHxJucJlC/
ME34JN1wSIO4NATqAufP5enMQq1LgMdkF/LJrRL/x3MzqpLzE0rjHrV2rFpvcyZZ
TjvNWn8Rn0wSbrsLJJV80yDLho4rUzmjca+Th52TpOXWAFISTqZcEF856PZRW1dR
PaUlecT6nbN/ej8cdcTTwyBZW7gxJKFJ22WfLn8+bJ7kyuAeLtfeqmYXcUpNoSxA
qUGeuo9vlLtTUVtn8U0UiVLHk8guLHHfEnu+yaq0NAZBMyFVFjmq/dDZTDAEEN6B
7RS+SRAtlgH20E3PQqcSzwT9GT2cgMumO+/W+q06Z38EqW2vzx7LBMoCmGuwUB/R
MX7W2X0OAXKzs1NdSeFJbrWwXY74lph7bt7peMzQVMPkxoTUoJkCQVUxX3XzGcx5
UrQieZvuIDBllsZ1PRsF3fpj5u4tkKdoBzfRDLC49RSq89/NCqiSWA+ht+F0CTKX
PfZzFy7aBqwztDQHFTqei61vJ3E5taV9zSU8VLNCcX1wSf35wgmwAER4RNR0nwwk
tIxIKd/2sj+/l81Fvw9qx0ByyPGqAG0hFxRN7w0cQtG6cV3usXRB1PG2hLJfLkcU
OpN0VABaS0lpfDZWGdeSgZJpcMB1rWpfV1/yVWFOWDYjgZOJQ9fhOUSU6x6iBXsU
njvwkR4VRMi4cigVRwKjC6W2a0BcOUZtAuCwtvSaGUD6+Lo2SjqL9xnEv3FKkkcL
rKVkm9jmH5GSNg40g8eCE7eOYMwhsIoTrb9HvGsLjsrag5vO3Dtzm7GZarpaBOx+
v565VYXLu772LpUEDPxVwDOQiI63xdpfuEizbSdoKDfaRl+2yurRgdxRDZNADGRM
W2Plgh6ECyE6i93RPvrANeKSY5vPYSi+LPK1R3DXrGVKZc5B8YQb9T77uv1MC4FA
D1gNQaDizhl7GYyt+sw44im1HFxjPHOz6CY+wE0nVRjL5HSGcksniKe75WFhIVCx
d9jmvBrj2GMKCuhDLQqFV1l4hcisiqdoCdXXEYOs+AIiDl8Utj+5k+Tf1XfQ6izk
01VXZ4HKbG53rz2Jd1urJiJSdJxdSKaIHDj/QEH7ONfNVdjfSLEQetqWGE2oPzGE
wPJeqXKrZMoXUenaDIOrBdTNY03sM2eZIJwuJgYD5TjO/kaxtz1kZN3kNjKFYodk
9LbqAvOvNXhV/4Cxq5/WtW7+EuP0ALyJuUrSKawGTqk=
`protect END_PROTECTED
