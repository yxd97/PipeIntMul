`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d2w07SB0v5Q9V9vfPR21snNrmuO2DAkugwGFL2FV1vVDaRMNT+6dYaZ26BQVWZXY
eho/N8Cs2IPdb23T7qv6ixcTzp22pPHm51fY0SLGXpH1fJg/L0z0jdTbQL0sVol4
u0Oe61GZDlUAXB5T/uvCvaSwVUU71Ju4m1+r7ZXCxj9435hiN0bsmbaVbgOVgQaQ
Ouwadf1dHHfxH15iy2RXOVAg9DoglFC/yPTRGMLnyJkV3rtF7+11i8JvMumJK0Ys
fG2fw1vLjGMcLyoKlPadyhrjdYmeV4zCPtZL0KlzIHRbSigTq6uSF4wVMsYTo1dc
iUjfhR+ZVdSpLk5e+kQD4Ivhw2zBibQpWeYNCETQoIlVUOuMnVvW+kpaTnkJeBUs
NYiSctYxSRPSg91JkQw/uaGyg2iH/cGNHkxVqJcA2YsGnmoDWzbhHkCm2YvuwwP8
JohPw/5Q/owd0tyAO2uVc3qWh2TuiM/rO6UhhetHopBcaKbDo3BhyszkDt9soa+l
N+wT2HpnY1xCQHm8m3ziiromy9qG9gDVcTUkuVC9MCkjqy+h6SAmVYfD7Yi69LpM
PjvYO3lMGJ/1+zdnG8nkKNDHHKoKo4ZwYx1tI6qqGQYg4Lg/YnEUg8WfHB4UTaPD
Mp8chjFj9dGKuZgkf13HeNd1teY3INolk4fIaHNQmfwDPpxQfnL0BClI0DuMWyFE
rVsP4fsEYfTrY9hIrn+th/aGsQsOjghbucX98bzsRmOBldSq+AZ9HPIOVBif4bsG
EYmOw8FjaU63NoT0egaDuDoMd1PS9sNplmLDQEDCoRMecdfEjpyBLwMoTXTpdiuL
xBeJzzPNjeXr6RX5ST4VB9jQtxvzOn+dFgm12GMq2/0wn3tH5iaSukfu2EcMUQe2
cwHZR5gt/ixB0WtlhmFmg0Xof1Kt7aO9WMJJbK6LFBkFRRpxrv+SFmNPHjSrSKSa
Rm7rvlHR4s9pM7gSt7yzetAASrqdi0YKbVU66qdYOc3L7wbKgwyAW28cSDs50wf3
eHthlssr6c9b2hsu/n8zYwjR8OgaM/TWFl4e1PpvtKyiFLiA62qFWRv1d4QRkrit
zAnRr1+fN/FkRu9V0m7gGdKN78ghjvgCBQyaGiZI/52MYp6J2TE4dkmfRXtbLV2z
EsDNzxQbD2lwnZGu/6kCq7QrGLHVqBQkMYbkn/y0M+mQ+VgKzAW7BqksR9mN0k5Z
+Z8jb7i1AOm78PmY/HUxwJnR82eubtrqQDk5LOjanIOQLyVCHswByKHYUzHkyh31
wwWeWDHdIqBsMPnFTQtFb2tXIPYla4QxcqGcd6RvDAJWQEQJ1cNdlRIqom99oxxT
6d59nn1G66LOhSkm/nFlJRMtVYDXci5fhWnzQLnZykDQlX6M96w58tX+KHclOAaB
+0c+LLs/PYuO7pdopRANQwVAHa12r+dpidSZsCJFw4FM1DEh2NETc0vy46mDnQ6p
7Bu3OsIG1USpykjvSBGwGTN/Pwiz8ltHMQCkm6Ao2VUPFySiHOgroL1EYYkW5qMR
I8DpmqzNx2SEDkQD6Orc1Qr35+654gFuFiNF6etE7zWLW56cjEiVzbtxaSm13POd
oJ/V3pDzA5eQPS0Rn/8S3QfomZnxisr1HtscNoVPFSYHEM4w5dsoHIAMBnWfgjFx
NL9p8rNlun6sJT96Z+YIoyNut08kI7CPPm2eQO5kKvuzNZu3tolVdQgwFlIdL1pN
373K6TYKFoOtOf6xZaV64dSKo4vgVQ2HPodHElIdYvieFNGlFW6Sg+d09TwaqeWt
VJQU/M+MgpG5YSv9CfZR5ZShkjR8QeaTs3tLmlzpjNkXF461YNRe/0MdtjgIMb9F
vg2GXHhXxsFnhQ8NkD7XtjiyrulK8E1NxAtyVysydxyattxdAolMyflSucK2Mh2h
9+IgKDgAKj6wSuTvyzGutNjoaVDQ1fmSab73ycUXK/82t7H2z8U/yginL9KcXjR8
2azGRWQmuLWwjo8eGfuRgMs9aMVujvtoLxduhAm60EhKxk0sjDo2n6L+I7cdLkIi
uUVIsJtHNkKcmI810b7n+7LuOtpw74qUjrqFMjLZxQjNmv/AK+6K3+jKFNixasEn
3mD6CWDLsxF4eI9dKOjWIuAgZtSoQCkyF2pkCDO7V516LbcROksqowUttI2t0TfL
ukDvIR5weoPbiPHEp0HhWG/QqYwCeZksukWeTKZaShAIvoc2WHYSc9Wl5jNrcLmY
rkIZ11fraRNgXnFCZNBq9GZrGrfciwzsV+IJyhKwoXbeqtz6pb0W6o+fEJLr+mOt
sRRWdQvgN2CWzBCNLRdoixyRPcHioXlfg6M5j1xbORYsZ8es866iZo4kPggg3uoX
Hy48hRJ0plj2i7YvuK8zSs4ycZ0+1QoZkhv95J2ewOz890ZNhZ++FjbZK6X1QS6u
39LwIUy+IvCpgf/HedMcWaabB4zl0qM7GFJFfAtH+U02JBsCTjDaYUXf+BLetnJU
qXR3QAK4uR5MwJAVzvT9VaqyOzpLtA1dXnxQtOMQj3dUFotORqRfITqqxvek/Dln
4lbzlycNE29aRAwX1ZTOvt+9L73Wrp6L1m/sIYG+adAOVSZ0Q96S1cTnBFljpQ7/
OaOOm30h7FmeM/VyCNikGuyGVRs8JK+et1oJaflJVe8pT9iWWaetZmEsJnwk6AaC
W3ybdiTkzLbbN5UO9kUSE8TpBfBnuUxlTNduEzPCXdmHpVtunfx4lpDq2xtLdtLU
itblSvUw0/Wosw0mjv/xtbTvD/nSyb2NQ1DrWpptL7C1acyvx+2+4SGUgL4oi81s
2ZfrTsOaeYtTEj8QK6m4kkFJuStgvKVtbOSxM2FuZ+FJdHEluJfhkfRLL5hTvhYL
MTsZlq8sm9VNwu2/Q+Tc4WLNR7DBUXwYnOVICujIj3MgzLJdmn75VjQTYnfpsOLU
Z1jdPEFS89/L5chq3dXShulXXZTwqTii6VTR1PZziFz9vXL3QOVzik0KZyFGaqbJ
Ntn4iAp4MKcVQ0Tr8JpyHLaQIzmkttzlRqi2jS6MJ6/ICAWuATcIEYd6WlC/9aOO
uujEPElqg9nZrwlJTn7D0nzRLPAx2o6eImE4ng4xSVp2aFSaxWDaMj5uFrEGmN1t
YQvDDepz5l+if9ClS7t+/hzIqPee06U+PWRztEbqRH83qSmsEkM0xBJQa4jwBoxO
eM8RTAJrTukow2E6gxwoGtHitfSVoswLUFJV7BsMhPciNnu+wohv1CSF3tdSuyeY
IHcyOrM/cQLYvqd1aNm1qLjDXvTyUgO27SVbt0IOjsn73Kw5TD7hnnB2fDWdByTt
dT17prBvcpLazxb8EghIQi7HWZgT7Vx61bttacqsStvr9LNSpoEYDs6bNyYxixrm
xRQRgpgvrWK/gmP/wwTskHb142i7fxBlpLTVBATMOtWkNmRWTWfHUF/511GSkDhB
QjoxmBMjHrGzDaPcKmF6UgXxVVml8q9kXDqiOkV7aOwSRRiqTf27xDZXZwHxdAnu
8236WG0q+m6DYtwu8kpENuAX6D4OSkCXiM2J60l4Rysb1z5zT9X3OVUl3mnyJzhf
efCqTyS2EFYRJ1wOtyF0dh+2eFEsTqDJxi3bPSDw6qP3n5xjQ4sSIHPHQD13N+pj
7cC5RpqU4LlnedZucrGjPm4n2iGe5n2aVBh1lU5wVbTwoYAIfMQQ9NLqbNU4EcLA
9+Rjw5baViNiGln5uGbjVgJPP+BvPKka3Rh+McX7y/pUyvZy7DvPTeh7G9C/dkxZ
R/AMyrHstpyvrCCZk1cR0Dyocnu/VhC8G73p4kI2FMPv8oSLDmp2UsG0+00fkOZG
Pz3TRseTJiy6nlHju+DIUrk03LCUrBT2frcJ7kW6YvrBtq++qZEu8xiYgYB0db/l
kxdHrvUBAKyHMxljuy45bNqPomka32QspyT/25ibuWDygaPRlI3IqkeL+SQo61w0
tpzM/e+QmqVbEKfEZq/c1q0Xq4iOqMQWNQ9NVAoHPa1AyvihSZIkLWGcO2u/oDXF
XgWI4Go+Q8FwEiFdJBgVxWYqVySIgtW3AIty4jBqF7JUCZc2XNlkxk3jUGLY2iXd
lq1PuG1hZUZ7QIwKSW0oB7MfHUxT9put6Ho+dD23gVh4i46R2rMikKPYjZTYc8+D
KPxAVasWK2e/zCUdCI7Ol6LkKNZ6WLNv63fTXYQOh+rju0Gjt2tOqrWJV5ihoVvp
5BQMxL9TskyQtPCIKVPO3SkTxCvVRB89IkEFQTJu/5S5uEB4ahjwlqfKy07rm9jj
56J4pCVAL0NbYocBC4nHXmBSGZl4vlPGxtHYlEJ0hIsbvRamoQETAXuy2QyXvkwE
TXowQkLWf439fLKTEV2KuBogogQxFV5tguyl+cekZY4ZvncZXj0Ejp/aUzM4Mm9M
BIl1Yl5hyt9KmI5doO9DpNi/FzeT84f404m54sJRHDS7dhghJQrC8K+DvpdnVGdl
tPnU16oOfzjKVV/aF4ogqqzifJJUWwLIyLoMwlxwPCkkqcPB5cg/jwiEu8L55B1a
5sasupy1SOpASXa9g+SF0va1gmsabp0p67O5UeJ1e69c8PPtC6dHnsKWSxXptK6Y
WWYR6Uq+7UP2gonA1KyyOCHZJuWTk/nQfgCvNMV6/SMZcjIr5xqPmm1joY2Y0rJO
HGgdJBYNqoA5Ec8A/m/jzB/xpoNrNA8Et8embyKgz5E+vGXf7L7dXfqI/vn62N6B
WNu181HfmaY+HRvn8wpL8NvbC1ey1WrFtXawerAh4Xx20FDu7rESA4JK7LDTzqNh
JNZrajb50GjI/krZo3iI0FZRFdQe5M0lwB4mK4U8H/avuvqU18S7NVwHqSSVYche
ZkVaz3GGTiEwSPxfhahYtKEj9+SI03IGKT4iV8WskBMILVerNxtI8sm7x2lf2AXj
z2VVP6joYs6RfCpFs6LuawvtmDcwUtjaFSmdzUvq3db5GXMTCrZWl1iLasoIaQvW
qpxZ5V0UDMzSxB7OeQF0xLV4TJMsPoVbVEt+ADbVJFzT/hojD/qURscGO+ovCUiO
uPRkoAIqRsCvJk0EtaczqO4CrBQIC4Y+JYzC75gOoO09GICfoOdS9lGkvxoEEXBb
4W7JYbJJCOp0nBeeMBt9N4Q10uZf3mYZlgVuvtaXf3WRHBkoGTYQB/TCEEMTTH1r
Cpktvvn2VJWMV9Qu70aAhPyFzvZP4no22QzU7HL+1Vd282bKjIBXgHMaahgxl3Zu
ai/YQf0afN4PrSVk6sxUkopvEYTlu54TdxrBFjyjkdj0Sh4OIEOH3V6lmC52C2L3
yuPybxdwYJ+YEXSPSlxDKRCXVulN8miDZzImwX7cz71geH12cKczD831t+TzMHJ7
PabzjTVE2/p+avQkJjaKn89cMRn4jR9XGbenQZyP2j8jYgJGypnzZKClxxGsE5Yq
Ch2/UeU4wzcB2vat7b6rfy+H7XgCfqAnVG7c/cx+eR+B2nNEasdnle0XtFkVlTCZ
Z5lOg5nB+FTe7n5hfuYkD4Xy8VA0V8YC/vTHkJca/01+XtlEcqwE6D11bIf+aOso
iVer0JO1R4JKphjgbi5QUIFLeiR/BrxxoQKe4XZqlxX6rxh4N+biNeM7czTvJp7G
QASB8Za3f1+IgSCVQpDqxgPW7ZTaYZip/n+SMpz48YbVOrA4Q3hF/UDVxsNNa8Hm
XZTMqmAfNQU6gls/D7hpk9WbZtgXD3OU/F7zAQBesZUx6xyj5Is0wFCGJTDRVTaq
6Leq7Ys4nTYCLxZl/exCA4c+7bjdXuv9P27oXtnMrPLTfJBTAaLrukp3Tn3267h2
Ek7aDi5uTzdZmt35KIHzNvRz7b9E4n/DFZ/Fk6Qa9bSWOWnv2DbUjZ2WRfH/LFgF
9dU0C/XxN44PgGZNn43iV6EEA6v9bt+742jX64E7ejAdHj519oWEDz4LgkpU1Dwx
2f2kJm85Bi3YsyOccHDHMjLw68zMrCwuU9L32W++zEL1Fa4L9m9LkAOf+gAoa+2k
PfpGmf034ED+Kecp5zK0m/0Dfy4oTmfbb2imi1S8PRB6MqUrPpNBi/eumg8TqStg
ZaPilfTPaV15uOO4KGb8wsvFwUkHGIVsHWCjai8ivvNFW/x3ovyMomGTfaQwWjkr
mEQuicDVkxT3DxiCKZVCd52LHLmdNDf/oyPoQW1wayQoZSh2177JITdMM4nBmsVb
xLXI/YpkC93QjQcEGY2/M82RcmF46MAwuU2RX5sYU/KeHmJBXPNiGevNcXsY4DCe
Eu+gPgwTkv7gaClyiBj0xCuZ32ykRtrwi/aMB4R8v1kxqJPo28hqDorjvTy7JQrH
eGIDNdIojzrQ84uXu4i4nlRhRUkByjEWQLNRS+iDHfxI/Zq1QxTdYFVslylQZhN9
aIruxaWoZt6PPziU1ucseOMz6LaNbjUYNxb8TkzF7QYfmCENnF89HzyGQKCD55uz
W82hGbU4cv5PXZjNHSURqrQfOHguCAaK1ZEmdCX8X8/+m2ApMxVplrUFU0r9hV20
NbM68l4NOrakb8wK5qu2MGRmF19TslpJysXCZIQDNqjbNMH7wiTnECAlKN+bDeut
8pqhEEZVdmBhztAj5yDR/2I8WF1dNNAeYlKC+ZfBKk2DYxx2GSpjhDE7AiS6+B/2
jyM1rtad+3nOVLEv/q6ZtZTmK5qAwLl6rpsTsG1EE6LOANc8gsKkmibsbag2hbkR
L34NjI8dX/YPY54nGZTNaw==
`protect END_PROTECTED
