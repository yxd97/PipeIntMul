`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Na2KHGMVRnUkOVigpgfDKM5M+B5i+26lZW3Wa3Qj+37/NU1hkTKNhNV+Dzp59JTn
HsXyTeXKSRHJ2NPdepxO3M1eu8asp2Srs6HFQxb9oa7RwGV6MBElIloKHMPQqgZS
L+RZiQ1DN4cYsCy2PXLtctfXjb4JildAbM0Dyi6xA8u/7UMf2JpqSk3VNaiX0kUG
7X06ZlccUnc4KED/ytSjzEzEFBHeB8PUIxYeEs31+eTz7ZIKpUgklr+ILEDVjlSQ
N/FcOjosunWot60BeWiaI4sWhkNImS6GDk+pVQ56Ja+vv3zLXLRtntp7NeaatBLs
b68qLbFmkP5ckvQ2Q/u4rZiR3n0XVBTcdmbli+Yf+KuA479nUn9/MtbwZqrLY4dR
qX4LIOtVn+cdzZpe1jGG+L0It5BsAkZetyH/En2/FQ6uzbeUmpik2XkvZ/UgvcsU
+4toqe/FST21Rpmm2LhEGpvPU30aQ2XxSaAaGDcJQBwuUz6zSpd9A5sknFzCvj+F
jEwqn5Jh1oqguHGi6fWZeQIDA8kwhyl3zOSbCAaYMNtQ3e+1Prd8WPZYPF6IIbJq
0i8PyZF/EKO7CQcbxeg7IUdw0vDUIPiM0jhO1zbn533LXjRk7FXGOnRIRsdMNM8y
5nSA/BDp+iYtIJ7c8vdi/0fw5w1+K/bxVv2r/nlAVtXzpIw25mPmBLrJ+2k9dRo7
2E6uxn1ict7KdCVOtvQY89hMM8AcTCteKPXlJwD2B0rNVmQCssBYEa4c+/eALAu4
JcjEit3V0WId7YI0yzhyFCdQ/LrDSyGpJYruOuNEssUcgEl85JJaIsstOOeY+eCj
T8vYEmwQw5ZFaDdwvlUEAnI1qEH6k3CagNGYTfCXnTCMlrCyrsxj7NxTYrmPusyH
Ey9LUizflDtIud4JHuSMe6MXKaI+oO1a1thzmAj4CzsBNiDVAd0NIfg75Tsh+ed1
`protect END_PROTECTED
