`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Knd/W+kBczqiGGqdPU0NOJEeu75KhXI4BhwycG86FUPvtE/7/Sx5mBbNvv0QxuZD
8SWbbj//DIFEysdI4Hg0TI8qp4s4GMs6E2uvneyNPSO+oY82kOtXLXbOqVihxzg3
HPT7QeRZ2oNAIpx2M8B5mSUAsp71GCLYrSgMRNygGHRQMe4nUNIJhF0GgUjJIYMt
2DrV34hY6r7gwnKCk995hwCccRmdgFI94temw4SChbnaNf9lsa+qMEo4Ud324LeV
sp68VbyfXT4QPjjcu7umGch6obKu8jHt0OQMgvEcfUqOaC7xNhe8S1dw90oDKq2b
j7EQp34hOPJrNdVd/ciBFIvKUQJchN4R1ZqpG+xgIKYLVI2sE6gtHEWMF947Fa4k
HjYk7Vt+fbf3om4DHzqy0StDh743cXvDZrDQKMDsfqC8VH4+IdhqFnqBGVdFRgQv
`protect END_PROTECTED
