`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9QgQf2ZMAKUGSlsFohMW+aWOfZMKKdEZ3Zx3Fc7CZXmfcAPc/XMN6KRicwWGFciI
6bOyMrVslftbdl4VLb0v/y524MtGwLVEwA/aoQdmYxOnJzL0wz7EMe4uDdvuBra3
muYLL5wo1FJ9XOW0WHSyjAq/nvinWX9V8pXBRcpS1N0H2HC5W9JDrWTqoSw6GmYE
D4MuCA1FWwlvXHbobw4VdaWAh0G4WCP+GPPOE8RiHnBiJ9LRg6ItZgDMWXiF7gkv
dB2NtXeEMILLuSa84n7PfnF5NpM7yuEf3xyme/x8r05dqc+KoqbXaqXgx9hiCFxY
JHlxIrLzehoIPkh4hCbJLiEJaTiPredLuP4lPFejaeAbJ6h+Vo8Q/MEi7Rqp6C0J
be3RXgNOmg1lNqbqpj2zmjEENCKw+wq/KfDImM71jG0boUT9wJPUeLHixQBg1efE
rGEM9ZToaQVSQDsLhCh0jFMz2h/0JdJwCKfFiUVup/TVDP5nqcPjPVfyhPnuFB6q
kM6OwnPSwPADxYRIQGH1p6Lem6PESSGC7z8WEETrBPrpX+65Tn0cwgqp9KUFO4ZJ
lxpHGYyE6nxNAdXmimF1uyPFmDJ5G4nWXgIW52jlsMxjUyLMgJt0bf3fAaTZL79U
LqMObSFllTqQzuQbP0LUvVl3hJbBxRL4DUH72wO7ubWQmFoSTctt69wMzXBmIzjW
mnU5G7SaUaObY19DEPPIXf1/bxdnmtodHgLO7GNfdfLUcxy6bsrgVZwt/fj98oI1
sqDJdD3FxjkkhUzNzNa5ll8HEaTwWDLSjnY7tg4xvLBn/aIehbAvYuf0Mn3t+YJ6
l48X/od11dyV7AFAaEowaGWrNjWX43cL7YrcG081snpElbIyyNuIJ7zuM0T/DPzR
q5Gbonzi1EcJZhJ9X16gC1DHqkc9tiBB4WF0XcVzRlRscjTFG6ujC5Jar1UcHPU+
e4vp86uawn39+jP7HC0bO+sCRWwwzQz4aKDmWQWk9FIydQgJ/QzKBjzJDuKRPdQN
7K5Y0OCzEGsxwwHYR8D2sJSarmqpN7NNqNEr69dRR3rn8a31UodjGqDSitF4NeH1
nxheLW24GMzNQEV2RAueTgDZKzxRC2/A0hyn+N4MEJUmy/owqJEP9JRvT8Ha2Vv5
g6GlTtXW3vCG/RVtvecn75QUf7EhzypNPXp+pKuEci/Gr0bWdNgM+VPZNZiKdoCc
gs0ksLSIXoFQqEeD7L6jaFlCP51THf8mZlQFJnyHMv3E5yQ6mLNzucI2dJHh1tXb
Z/kBlsqgQE8cH5mgZZwHRIyMY8ZUOXNBhdl+vui6A5MmShhNDfetIGz+FKNikeE1
8afSEoNuu1Kc0fsTMEO3NZwVrrOw+icyQRd9bsxGHTE9i1SZ/M1Njb+b1fCoI23x
VxM/QCuxETcxS4aWHCiEwKaOR1nx3QbVYcsSTzbT3G5fl5eeYeIG7BvFFxISBw3T
w8lY7P+ZjC2i6WyJSQX/EahU4vVQYaUWcUzqckOhbHcwPE1yqcHtxTIDzlROr7D3
ALgyrev9niCXR4X/xZ2k81ksYsQBooRCy1HEKdZGYqHzvF6Wtg8hnDxLKMw+nbsM
ATZbopgWukJE3//c4GDf4W7E/nDjoiNSY1gmH8orvet4Ut1g8qR1lnhBXI5nCMPi
i+Jggs27fr3QsDmUAA/WuilonwvBGJE04jSy1UQfaMoivjTvRvV7zWGOvKZ6dlCo
WrzVWYz2e2W6bD+wFhNyhx05TzAXgLCls7GZ/2m4ak0o814TfMpoVW3EYIZIQzi2
1osr6O8gn0WCXSqD39kL9IsC+LtWOgHhrdC7wJJ5Wa3k9EN5a7HeBekS5mscqFVv
VidKiCK/vbMd0G2gVnF0tGLkaLl/iS7ATWS0GgXepn0ug01z0lQqiKP8ZVXUVngT
O/pne64ozcLQO4PnmWav3F26Ax0+jgY3B1aPkGMA+xW2MCNfpBkYUj0ykPwu4Dqa
QNIBeu95+aSgL/x6v7qzL5gt4fWBEZ+PzcO07CzSdBSjTcUsQgT5nYLtP/M2ThQe
ZCxlNUuA1JLre18OvWJU3t/Q+Nv1Ar3sH3+XN0wuRBSjIx2SwSdZCdCxuh+dTUXU
FsvFIty8RibyUlrDjY2Fhgz6tSPUnIlmctNsgIHDSQE4AwL+VaMYmyUHImw/5sQS
82wjKzmvOa+uwBjIjT9l8MEcMgv6bAcR/uUHDZFJpqvw0keCXw0qWn+ZMBoToNvh
YUiYsI0cyocDv9Jnhp4H2X20qUQD78x1vYsBj40+gXsehyIyVgH4HiMEMrQBdKA4
RxByKsrFnHVbelYIWkdDeOdXO6JD822FcutkxsYmbnDbMdWyz2Wy71hHTAytsunF
uzukPfG29nEJCEmMFk3XtdyZwH2sCopjm+VGcNyVa4bxaTP86VoQbJCc8Tjf+xmn
XfTJsvgXEJ7FTDOzzW/Y6CU3UL8zDl/cgTkpMDQyRLY=
`protect END_PROTECTED
