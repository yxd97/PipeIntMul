`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhNXrdF41usQjYs1T4puNJvj78tBSLVJtWvEoxpUoMm8tL7C0+VCPNWtBNhxzlya
i/sf3prMXnDe+1N6StL4F+nOtu3dETLqlbfo0S2Viu26JbGD37TuqJzXbyHDgG5V
r4r21aqaL/9rGmwtcRwameXbMmZfQ4Z6/IsMAuUjNhAAjJATZHj5Le5XbCLJRSow
/dQ9ftFMvhYwu60K3Y2PGOMxPY4g1kJ/gqy6DvN+NTTI0IxZa8Y6Wt3AlY+N/eRY
FtNe8M+5tfUO46FwTKQbf6jf/+o5Web8uU4M+j+A5lQIJIS/kGC6PRrfJVJdshas
M6dPkumciprjiOldpY+yhE68UTSUrSHJwGRvJJyAh+41QDuKEGxCfasDfNFfiIJb
ax28xbcmWMzG4racY3N7CRU+3blBYwgMZWfsPz2PPyHzXRLCDMTFe5m67Gv/5Ot1
lHUuZTTn7neti7F9HgHGXLeCZIQOg0RjpRP4XsOVX5tluE5OoKs80Ac3/jNJLDTU
LrOW38p2/ZaR4xhcHTVX46SynKM7bb+Yt/2qXGPsozBetXTfDImzh2jW2m6IT/Vs
i9IriQyocpaP7hHhrjrJ/aMYLpcHG5S53W9dCl0Ngbk+gmx6atmdj00W8o1FYIMz
HWdfMXa1ANdlwg6giFh5zZG6+pOwx9/gLFhIAVR9FGGsZYUpDgfA5Sfc/DDPdXja
nsHNEYiUB1tA7cVNkmz9nOafG0kN/N3fMDy3nL+D2o9PmKo8OHUlw/UlOLA92uEf
hFJY8Zgln+NcIE99L0i9W65WiT0AR2LAjrAkvoDsmcQZDNZSmZS2rd4GLVP67pP0
iajCYnoiABxTrlJ95Vhiy/soScE+JlGU2/JRzJjzIbvJ2YNbOgT9iHLxP8U7z1UI
FPrUsYyLTQMyhUE1zYntDUfPF4xSpfjP+7eo50rNc8Tr8grJk/wx95bnq35KKHFP
bBOHkW9ovu6SIY2iOhZc7ow39pZcSpnkZa+u8nSHI7GhY9exb4qnIdw5rsMOqjfn
sqhTJdjbDRWPT2oKailTdKEvexV9lKETwxbpHMo0hvcLKRyLuGXcaNPUKK2sQLye
ZC5EEte3FMN5lpVNiKNV4awQtaniS4PbTYBOlS2dv3Ew1qrvrz2JBx/AnFUskwiz
Q6FIAXZ7LVfULsn+MRsMg1zxgAnUI9oHIK7ca5LM95tP7qU2o05ghqYMa3I4lJbi
y6FcyRVhlIxv4d8mCOERK8iH1EVNeOCS/wiZeBo4SkKn0sxmpExr8QVRSX4APVag
M8LqUM20mz8rl3PEhhCCJj5Dl49K6axuKTQTkzfo97TG23Aj6kSNKmSAGxbeVPni
`protect END_PROTECTED
