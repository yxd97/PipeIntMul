`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dA5mum1ITd0okf0n3OSvAzY6tR9lyXX3RZkFlSl3xWDS0P6W9mjqF8euSt/agL4H
zPcP2WG6MTQMPUAk42kLBrB+fqpDEp8F8HjQi15AcO9kuuoo2reyv2K1GwkfoJgh
YhNQ6TGTIpsmVzAxT1th3xxteEreNbg5PNUi9EAPhC8n8gZbpRns/S1z1nE/Hbrp
L3YJhTMgo3t68CASrmCfFYm3dH0TLDWP7LvCKqTNrJu7BvgKIAErf6IX3ybP+cDI
HJNoYfpWKCqM4loTGRYg0IkJriI5qwQmpykregnqkE2XfCEgUyiaKKnGuOLmM894
GgdMR1KpvAOyi9M3QL9IdHre4yh/EIdIasJkVB88fJxhbjnF5TbqtFdELHxwxMW+
i3ApSoXKxu4Ys3HVbVC8k8jpoiM2P1Cd2Ty2Nbp80CkcCY4L89WbEihDUEuDCoH2
NQmZo6yfIeGPaIEcBRlpo+3m78ju6lp8a5I526DUmEoI9yaAg8LAekGF0YRc0XLU
GE5ZlZqZbqAYqSOjGp2gPwfmDg5clB2NUcUvyRQNfXDiF0elyObTk1RWT80yn4j8
dUU+YHfiw7w7NhoS3iZX5Cd1mX7GLQM2wJ1JJv6/X6+c3eqaw/eoI3pXK0kFqB4+
PNDWDJijg0cJHYxg2FHT05F6wip4erEpZ9IYMm1N6Ye8N9JtZAg8aMcGOSJjgRWC
p2o51Sy2hSQD0+Km2r9PjX9SVQvX52wZXthu/p8l228=
`protect END_PROTECTED
