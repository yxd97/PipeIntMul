`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZEgeYN0+EwitSwfLzW/7sNCD561gkEsEMuQ+FFPJyN2OPGfLIIOwTselbeoq3MVO
ppWylz3ID4yhkiyd9GgbfHJe6cEAw+rR7SyyCxD1Dz1dpEacM4eVN/6aNEW0Sj6r
N+iLkw+vNe0K+QCJIEh7AeVE5qp4gpfPitaa5O7a9FGcZpD6iDKxx4kydrAOnCN+
T2F4SYTFlBCSHs8OqS5UjN3EIqmpy8xhdSZHihyvG18tx9yJtNy4aI6DXo+foJ7V
`protect END_PROTECTED
