`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1+U0JpbnpmWPbKxM/KQ67SGzr6bi6hn4PMu7xgIy/UkorZE54mXa2lw17+MSzxvD
tOGXoJinsFzFMAfGHBo3KLxfVVfNrr07iliU3ABILOp/Nd6cCxDB1e2LRKPm/UDk
ZYHcMyqLfJjkvQ4h3AFLgwOzEGuF0O9NsZ/sct4r2/YhkJtIq4LCeTSiTIVfU9ra
aIGO81ugX51baiZw9HfxQvK3e62/KnXEoRDBbKv7D4PJno4V6lEte67O40fkRaNl
oOppl9gb7K1cwHsMkhF5Sfm3UcZafrmfttPHAEtaMf1bMx+NL8DlEARczdrPHo/x
B0CR49y6gHZpxrb10lK30i2qNyoVehU58wk5wurzwcwhahWGmQAOqUx5Bjg1Lfar
jHkBk6uO68BIvfUBnv8ohu3EEyTjSA0dAyhmHAXod9Lg5CDgZWQMkyWcUlUssOj9
cw7l6lOOTO0D2ypNeFIuC0ZrJoS9h7ysOuHvJ6Q0n8qiLYzISHdhlu/F2knVtog1
pn2S9biLHiVnOlRMpVqxolIyl0NdgWNGY0p95OjoIs7OycZCnlsLHg3rz5HT9j5j
pyilRlbAGiuh5J4nd2Y29Kg91fhbOhhfDNMDxlHfiYa3MJmpXTw23OefEFUGbF2q
agNEpnsbGCZ5kayY/PQgsxYXyFQ989KWRYigvbVUZ3ULjGzpilVqMGGJ1rK1qD4j
NFJ3x5VyhjTBXXFWqNeD5EqQltzqSgXXB8HzU0+oYf4lSJzn7O+oacpoCqJboztn
VSXKKtGdxpD+WLy4/fxQWKFnzWZs7PJJw0ichjawhC0eHNOqMHq/mKZXiXuVUiWt
wvxiW+HD8VLP9s1G2wJA79V/l/AMaCP31Kow+hht3ySFT6vDzGQFvihNhZ9xX0Yu
81TON2nrPfmhVVNdibTSVD5YJqlXC9nkrxodI4YhR4nEHr9VSlmgsWcUNPUrLtX/
C5Q6ep/AzoxfMOeZuAPhgW3t0GdPfjrOMTZQQ6wuGyTp3Fa20ZfntkD98t5QMvrA
4xMYobtPbyX0Ymny5IdPWfUwklY5FDT0v2GIXYfmWNzKCKc2kD2pUJFNEItlDDGH
lkOKjgmAPd6Z297cLtJYDOmaJWAutixFPnBTtWSvWMMeyDO5De/zMQ8gYfRTMQFE
eOHNwrrVY90+AnTAkmyYsjesttNDN9mYsqieA2/W4QHT0N3foGkFpbUGd6iWsEA7
zLpyisxSMUa2Gs2umltkf9E74TrCLzLqWVu3H2tA89Ew4RRNazB+MeuY18u+tStp
Ch/BQpiJMBMnN6e0TRhQs/oDSW2VG39HQN++/oFD3Rku6lXV9IgG0GB1u70Fjh1k
s6Lo6Y0OItBrQuNjgfZWx7bRERGxTw5sn2UKxSdjq/G4he0RCWOyGShRIzKM4GVg
Pez4FNLBAswXjXmcRAkLSrKI7zL6v9pG4MHd+W/6ObSokhqMIg8SK9CB2GjnTXNa
TZXOfyDtsAfDsvILeO6ai6/nzsz8LAYfNtpxvfrbvTJDwoC+Ex8vssLEPuwCgVXg
YecNEY1V7HBCd7mpKy/MWvevUK8r94YKdUuLqckCJ4IpaeTWQfaDpB+o4XJdySGA
TkX2u8DhwFBU+7SmmvpX9tj3xmmPYy3/+gseEFAKKhDSCrJxsOJp8UAAaQ8mWHL6
BD3bivOGwXqHPQDOTQNxnL3/0qpRyBk+pR61adA8w9JX6rQOKlCsFdsZJE3oO0aZ
vyIcBTZucxGZP3xD2CqPQRK6xcyKBXsqyCQDZ5q7cV00NRB2fefcI7EZggn2M7S5
cQTXmQ2lgEdU7SRRvfp6jpr+hsrAVxqrRlFzW+pQ9RI1lqtXToa/1qDakef5SrOz
I6H9jw5vQkaa9F8Uh+rPPetJYCVH8XwP+rvb6jB0j4Fnxo6zWpqaQRdEjftv3e5u
hDPcjyUjbwVLT6xCZaRe5qu4T307xnjCXF3xUH7Igi83UEsLpDFnhrJLLQihnROE
sCJV/t9jtSwap2jT3QY/Nilk9BNAj0q2lGI/WGm2fxvnv/TkuWxkcRMGZsHx7Qz1
eYpmfJsPbI1abjylU8lLZ+mZUr3UG1HwHw3tvLEz+R0YjnEHLFBgS0j9Lt7CjACP
6KEKpcY2CErM9AAid13Y9JRIuBLkN34TZTFsJYf+bdHy8WRD/wWA4r7TGt/WMb6g
+mWdavRorMKSuDnePbh+jCtkymlaEJAxgtbTppyKi0gFOO8N4Hie7LXgKS8BDiOl
eMxrv/8Ul++SiaxP065vVWgHog1xdbczBcI8h82S1CCG/+RvMS+cMdmbnb0ALnF3
DcvZ0omE2A0m8Zd5cH9+dWremMYox6cdFwAlC92Tg2L5WcqUSAKgfdvQCzBjn4xn
7y8vvi3IyUBatac8M2ucs4hXzp6N9tO3k8QcwAJ3YBL8GKzVbqbyX+3laW1LYEiW
wKH24HbQlTarG9NDylggteaPksx/MoqkrNldLjyifRDexidUpeXOERmbcJPM4Vun
VI4kxwso0eNcTtR1aBAL5QZ2KchaAe5n6YdwF+i5/jlcMtBWUDLLyz2xA6AUjHzJ
HwvYiksyGAzFtSLaVfibo0fpBcLpen3RL2g9GhoDwhLiASzVlCLbR/1k+FvjJUaY
P2sQH63FuA6zxEb8JSk9s9htG5vlFxKWQoGIl12TX4AsPaZpQVyF0Dc4RU1v0VLb
bDpIAeRXWP/YWCYMeEbB6PqXkCclYmBPkQcrTEbkGqlXGS+5KDZs+sptPnkKatmA
uGH8iVwFeeyOheZxlC+9p/y/BVhLyl+uGcefyigndClWqay3ECZdD/zYPGmUNzUX
9FmfmybQ+UluuPt8WbhaD1LZo8fyRlIWscN/idi0aZSc2BFdaCOpFgYxPIqw5CJe
szX4IQHfWAuEG6QBiyl3i5Zgiy7Ky9yDC2gjTjHB1VCXE591cYCw2cMGWfuf+6jd
zEmlRUroSu1/5OYspLzZL4Zf2j2glPBVzZlmt5i05DFnPk00SDRqmzo7XzomHY/V
HQNUtJrcuVqXAnCEw3MV5cuSwXia6CdQRWNe9iEt6BAHsW9D7Y5ixE4/KNroc+EC
RCEoeRiyQgWhRwH/YbKlFu+KjnggiTiIn7Iy7qQkeWLir+uG2aGEiiT/Czk1lpeJ
KkY4uV9WW6sVZtoq7abYCnLHESooO8aoe0FzcFyM+NLHSkrl5aFGnNTzPohRCHZ5
FDDXglgjOn+dxhsRFbL3Cowkjie/hTYgFwqVH2H/Z21K1PBj+m09URbRRdiq+Pb6
OcRkeOs9K+p7hIG8uFHlNzcNA0jLoX+bHXJOLHKV6RE0y1TQa/23fYrWWYeiWGyv
DkGCl6xP4CRe+kPmPGxGKTmG9/vuVPuJ/asNIWJyKxtvdLFcAsH8gT4ioCP2UXCE
`protect END_PROTECTED
