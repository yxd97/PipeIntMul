`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tm7zq6ETVcatdx2gFEQySHCsyTJ9ynoCLyDyygnGG05uLPa7Vp3TZBxztJJL3/jz
8ObLBmbMjTKdP4CSYnoxK0Iu4XW1nT4Rw+bswnxFFMpeAJnDGt0y6cqXkJ1tHv10
Ng66ix/gKr13RSsuZzQv+mplVv0KrwtMHxPikRFj8ReuV7FTOda8RpHvl05qpvCz
bAqxycvuPbMA85NjJvAIsfS2EVLlmMIsA5LpW+4NHzS9iyXXMaBRZ62ecX5Yhm0R
L5oXEG9Psg95svJIFQkRDZvj5QqCqMW0nUVllh3cwdoh8XkfRBOBG8fcDE7fTICQ
VMRDu4Ma8jaOAIbt2gUh5Uioyx4vm3oqZ4XY0joUH2hbyl2aSStPRjogulD3B75Q
fSM1dpdfV6FHXv735TTx1/IyNX7I2mspz4vJU9qjRVX/fP99sHNwraKbTJbSI709
yQsX1TQvZtUAgHGPHu1yJ9ICbgaHpBJ0mV8Ywsc9PgPIwYXlJig47DHZv8rPzABA
cnxJmZaOBKLk6QXxKQ3i0Dq22LOYL4scFxtBOBY6Elx//xukOMyrn7QROKB7EFiR
22Bzoi6c344njtYZZksPA6Dv2Zy+r/kedBQ2Dw82aLEjT5kOvzEFrhdyjHAXnhY3
yjN2dVKCtneJs64sBe9suy+9cnYlLqntGLS2I9ajTSumRvumqDlS8s7utFxL37zA
yAOPKIO1tUuhU8EanuFRu+CZa5sOelyQ14zf1YEEJu/Sw9Hb4+PBnexGZklgcQrL
0np8pg0OEz7S5laJ7Jn8sE/amfrUtS4ueHU3hMsBckInwSZ2dloL2cHYjJcPwt9j
/ScB8CM5qB/JrRiTQaPV/ynqF+Txl4qI1SsRTsqcepHVhhnThROIUIXdaSfBgE1a
gfR/PB5gQlaMNr9iPhHSa6fSdl+UayotGIvLMBAxE9rkpZ0QAIQmz4NwA9zY8tH5
Z2OW+kRnps1f0zCNY95HNzoCXNfdwJoLzQ14J+S5xMFsoedqZPBfq+bY/aYT6QAW
RTMp700wW8pDawUOpfMwSkhpgtMgV/Kjr6LBf6zc8Ri/U4FQ6wpR566yZBtIfyDD
YWW77rt7jNzrZtX/i6fk+tWM4HOO7wmxyLtVjkaFotCKZXD3WCCdMZySPWyRYCHv
`protect END_PROTECTED
