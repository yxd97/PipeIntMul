`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wHIGYKB8v67FpmuTmB4S/PSbafTrz/qidJqt0UtTnqMjoV51aK/UL5SDiUYiUexJ
7lWa1Kr2f68UkfkC+Jnd9QhKRxg0zbwePbbIdDXLqCfQ7LXJbtyPt6mk61pNhOHB
w1fbpJ2raXFlvHYrnvztImXu5WmZiYvEtOIH2f+1yqD8F99oxOh8N5prk7Yax/yV
lgDsuzRWq9IHn0TncIdLV4BrhgswIPjSZZymZmsklTaE+GbZerC5aMQpgM2dYiOl
lrW/XF5OewIHXAq40ThDOrpSR4EiC94iy48RSQ02LrqbXPquX9P7idcf8ewpn3P9
nNkJ2ShhzJjz+BlNvvaT34S/hcjy95BuMe68e49Vp/fR6AqzU6jfZRc3cw6T7Nmb
CuDJmFfhf6Q1I9dHqKnGKTzvIso/gjoC9EDqY/AcMXE5So+HmctsiBtS42pyZ1Kh
`protect END_PROTECTED
