`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T+T7t+j8SAh2uZ8i/A2AWjCWnxC0Fp46qr2makIyaHSO8EDiK3cXmR0IDEgynALI
kJfj4a/hZcvLQVKeTSASyqZyRmDWAsbwLmFrCE+xEJFqf3HO56attPe6VugvQiC0
PKwcnryP4TN24gd7YjLJdyGfRjC7Dpxsx3imYOrGEL9RDUXZNvXrP+XzVjRD7WoX
D4+5yowTQC8mx3MmpJ/+TVw22xnm3DYIkC85y10OqSOY2cWwVLfY0IiMmAOkdi6t
t2lumBVzD3INfyWZnN0TBT1hFMjxa2M6RjRNDpE9IauWH9d/O9Yto+JS8qGmWF/M
4ZR78pVW3lwKwdLfeGHmp9EnyD+IaDJBrw1tIiqIBdwmEO5i/b4TKD7EhSZOuU7l
slVhcINVStVsFXQVzlsev3LMgiTRTh0WPXw6FEXlBJQoTZiIqPXB5Zsdt5eqYeRV
`protect END_PROTECTED
