`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0w4pQKDngjwh8cSZlVPsSICXSDw/WSA1vKJLXdA1Pxpd1OduDbfLxzrSyyVW6WtI
btrERFDyf6KB9xaftiCKS0yjGTdHjSWs6bNFIdAzLu8trTytWaxwgJL1uawkQSul
39rKOIRnO5ugglAENXWQPXHdUxqU/oPDMZb9PlvQLDrLWNYI6OFSbf7UAWd5tsgJ
1uV/lNI6qeGf2Z/mQbf6+8NKE1ad8IefwGxCahx3f9d3HYzTsdGQ4fnNEejZH5Ps
VQzjYID1PnJ40Tm7RZD5t2G6DDab76ryONlfe6WGFnU=
`protect END_PROTECTED
