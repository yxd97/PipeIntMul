`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZOPS6oLzXRXCmG1h8ce4EW2ScmkX35OEX604xusW5CzhWeU6aHkdkX+/RjjRazF
Q4ol3KqbUKIxOur/mtWEnIekhoGOABwieTIJhNjHmKAKI0sFCP9TK0cgMHa6yYtd
KKAAzfbaTAoEXoT4q4zpjcXcVUVlM42cigXBg70MsMhqar6hzYczYCvOEyKI3Xe5
PZXC1nv2T45lPaALN2PkL4B1rx1o8vBXsDGeMY+1qFRE7pwUvybYvTBeIAJ2aQSR
79yreYJipauCCSXBnPKnq1Fm08I+UcZaxG/ke3XIInI=
`protect END_PROTECTED
