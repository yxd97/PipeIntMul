`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHRAl+x5UmBL8AOS+ZEvGYdGfR6gURi++3oMIwjiBnVkBYYOM+EJG8YNTOVT8bKN
MuhZIsLZwsbyDGE9hTDuJT82s4bfM4WFeQidBUbQ+XIrmq4q7duV/GZ4UMrBAUoV
tT7E0G4CEg2pgYjvU72+a5nUfJGsfStbfSrTYZ7RKgq/KZCcE1gNRpuPYVK+v1AS
hkI/iIAvIQmBF2ga8IQ37iTOj42kJh/gDGNhAeJ77LJLuqP9lEbpuoNb0OBBWHGn
bjZzM7WV68U6DRf6fhxU2ZCeQPczjhP14H4H3zH9YP5jSrvGdOjD1iiMrgcfHpQp
by+rloC3D0W51cpO0RncPx2EYQ8uH65/iIiioxrTcEOrxbMQZ8nZJHwq7lN3QSUS
CTicUumwRDO7eetQvAcsyfuGom7NhEP4rDvB5SstiMR5Ekk2nwihADfyUF2J3Nqd
5FFADZCHaOvRsm1AyBnQHJCMc/VJxuCkVfEVHMfpkZUnn4lsiWG/rYyft1dPQaJY
ikdV4s6a4nw697vdOBCUL2KlWV6w/sGbmAPAv7cnrku0Yr0QsaKk3HPXmKbOud+J
RzqOhQs4cnkzjVOrPO/TuGK6BU3zfdS/ftbccsRrPycYK0eLXgLYd67eY8GaNLRr
gYhONNJ4B0VjWPrlFEzYG3GUu3eKwetjH9VaOjHRkFqfu+DAoZgZj6+aljuHeDO0
/FQ1r7WxRJ62OxrTALjht5d90dbd8gbk1LwO7aUSW4a61ej2zq8NH7OBH7E9Fcy9
67fV2k62L1O/s3DHbQldf9gxm0CrPnAGCFc1qw4NXrlDAEI8Wdw2bg2L+uLYz5Za
YXtdsc3Yssogit3bJJdiT18W1RkklXRRRA1OoXrdQO2dqxm51Ob44W1rZJTE8uJ8
`protect END_PROTECTED
