`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vi13u9AHd4Y5afZvwMITJNjoM5fjmNNB3VqRP7KTHR/E+CFkFhbn1qtLHIf8cv2l
tioKRSjC57OWnUk/pS+2Lqcw8Ll9BrhrDVzwrfu175TKUCVaFErYPEAHm1ilsFKj
JU0lJ2x7RgGchexZnLUri1spNioc+gFs4BGwYCEPgQAr4MwPKUcmHn8Gyc6mqnRH
vRxqHDu+gR5k8cVyII1kOsWSWBXonIPSP7t1Rx2snGZJ4rdh1q0dXAeUrXH+MO3N
hqJA7OdNgfaIB6j4Ay/mtAWD1Or6bHRMjVOWTPpMKl6FKW21uI0e4ebM5/U21fg3
+B06SozrrOpeFGCp5kT0uZq1rT5+wCaaTwYIvxRSQOyMBcBKHwfxeGfcaaZZCFFQ
hgY832lrXnadCAvCT330AVdN546bvj2M+QzURsvjLwUST0jSASh5wG+vNBYhoZ8b
C2xa4jFsitMHUWWI2eMPgtoTfaKsdAkNV+NTYXXQU3Ae4QUraedViLYvXM2cMgmh
3V7eBsUPOvv2N/PlkD9Bfrayf2hwx4bW0wRt2MYTBMy3U/9dhdI2Y7QXuumU5T2H
3uFgDJuIOM7TT2HBmrspYcahTh5F67qDl8AIy/9AsB3tp/q6agT/jagJx8qRgpRW
bvhG63IK9NEyS6HAHDb7qzSKyKHMUCfs1J++M3aVEMODfibsh1EurSImrePm08um
VyUrfdKC6Sf5/ZuHl+Ps56kXxmNDHif9U4/wH8J0XDCx8eK0KwUWypBMDXNwGicK
fPmLemT28EylRy/m/Xk/i1uu78nwAWxGk+P3D/4rJdLJ3uyb405kU2sGgGagdm77
yy3aCLp1qMnBao1omvU9Z9hslxo9T5F8Y8+HpRrtuY6h04Frey+/OmztLCfDjqsO
5DV+nl4hTb6e2j3jSraG3ypYzIOETNy2gDY1wtcvBQp13IpxFlTS3K+MY2dGMF9N
/VrbLfTKN9pSvs/uA2l34o+QjphDLKRak6As6q1XM0b3QHVQaMBO1a+nsgMs7AD+
5jtCZPIZnf6E2kiG7aykDpaQp393VWsZbvvN9R8GYJd40sl2q9w/9DPYVyO221N+
FiHcLArHu5JCNBhKpg8zDOF+hjLtEtusBqwBG6wiEHI/IYUHMQT9r5IVNtnSKaYY
MLoxfiQBZOediT1oGr5RlXBUA0TB6xvLM5VVIuH+tq5yl8II9V42IBJR3gfsPd0d
QEWkmKrNfm3vgF5vqbT9jiiQ7xis/gad8H77+3AZSfNNNfWNjIqhgvIZ2LAntjSr
jUpPGOdBdAZogFKl7F0vW//aUcARS5TQ2m6jDRdULqYKrnfNHbj+1UDx7ye+nTqJ
fI1/ORMW9JbnF7dqQdi814EVo4fU6JTJUSvOXKHM6wGRZpN42e2YuKXGw2nVIyli
rzdu1GY9rRF+w972voEIqaGBGEBVRkaoG2QN+LBAiJ6Oc0Kj5Sz7VonoUR9l59Cd
x5Ldf5fX3olq7qwz8/IUU6GFAuu9pqLsK/LWZjbm1T8AGzTExktJuJRKS+eOTPyo
OgzJdg1GNH5BhusQDnWBrwf3WSmWLgJRedwg2IKgjvbRDMULvWxhRgjVkcbh8xk3
HA8CRhpDXpIy3OxRD4u9m8h+cDA3KvZSmeBoZVM4ds89V/EW4kWBWpNcZvmmhPUE
gUBi3osQ4DybSUuGDF7Agr6qHWjIVcuK/DC+SM3Nxx0cf2GBirpkHjgrs9EWbRW4
84iZWbjZhZHDBQBiCWPC13pqN27mPR9EmQnrGyGzeiccufdHnG2cnk77GZMBe/It
18kHERW14cOhViM9Ew0I4tSiy8NJ9xEGp09cIgG1x7XXPRkTCsezs/u7FavIQM3F
i+B2HHyBbbydnOZ5hgr2ecodTpdeDWsdIg7XlkKbUXmf4OGLctWSChj3rd0iFXQA
+kG5xFnvLLQOPhqLwxUK79vjQIORW/fcSxN55z35yTE=
`protect END_PROTECTED
