`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0IYXeeRMQAMs+7pRMDGLhtkiMJZj5U4ZwMaNkdsJY/qsV2iduw7NeFzHu5NfeyuL
Hec2sGzr8AK2H4u6sAQEPbKF4YAhI7Mb/03A90HcD0ABTp6mEpfuPmKcRMhWpX76
Da2bXrIW83NgK2vh099G1DbOgSQVHL4eppLt65tYV5ohsO9uUjm1OUSD57PZlctm
Vsmy+QpUsk2mYUBkyXh0tXrp6fko8IUsXI6pY7WrGpE/5FQcHzH1oT6qY2XSafxX
rugGVcSpSRPZayHpblorxHDtFRRJgVeoz0xR9SpevcxF5UpQgBUwiNqmoId8mIvP
x0MOyy6nCbeU0V2xeXvBmuHrGCIu/26iWaAO7W8zJeqM25N7Ym5/0+74YcdeZioO
eOwo8bF/T7G9g6LVU8YEMpeYpWGai5/v/JmsDqmGxYEYnZGFdZNRqIueWZBlKjwH
PLSKmSuvJybxJJGE6fDYbu4DrsuL7t/VcNH/suf/zKYNlyRl3kToZbaP2xbYg6X4
698fYUc4Ra8la+D4SCh7/pZxQD4XGXJzQ0+61pPHkADF43alJ4Apcvo3H851EO/9
pJBLhD0UipQFy7TFLe8RksIYnfUwrpkISNni27RONYYn60OXgCfW0RqyNxqbHFi2
FVNgbGwE1+Je4hX8TVpifa71lS2A/WRQFUpXR0E/wLQuQkn7cCH8ivIYRH48ZBDh
+kYpnoEy8R0TW5ZfMUgYgEh9JHL2lt+6umA6Dce5v+zoUNxi/KPE0BmCcq4qKBIo
tP0P3xb96eioDW4hIiaVohE9YdCyl8nJ0owO9tD8bcu5EVnDqALijo5X1HjB5d7S
23kyoLMaN2rtKIzOP156LQdSOnZIumpc+y1S6QDGoUPpKRLHGBOUvk0H9dVKVlNg
VW/JbdU/CDX8LhGcjbTG7RXTMZzUeWOQLVltGqMSsksiCzfY0rvZgb1S2JajeaXz
ZJqEbIUGP2+T9xQbQyZnxV+TjqgKQBIsJxTndiEOZ8oBtZVmYJsjNipa8X8EOmLy
1zwJOJK7NrYSvHjnKqg8q7XldtAO/h/2SK+P99/vL02v1/QCNpd+2ScCdqHdm85f
lS11ysWMpVs6rilm/JFMzD59XLvP/hHCpU8dv643G0TQ3dO1N9EwmAX5KbbwcGT6
N3ZaAFeWXLiO3iY4zG9Kf3zVest6FNldXphJj3d8SLqG0TUtd/eck7FU7Sc8cAfP
HkzltCXhaHEKLyKpG0GZnq4mArwnvQXpV1gZXg7QZpmDmAdxP7Gne+7U4kNW2v9M
iqYYT5Tnt531F4Ng0YGH5bqZHezvvGwsA8vpN88a4OVqb9oX1n3dfQCftgNeq27L
zU28lPG3kc6K57V4p40b8orRH4ahuR/u8sY/9hkGDXwJEkY9v9fOZDD2NOPps7PT
lhZ6vRZu/Aji078mCh190N3333n/CBMUuauxxi1gQeGV2jT/UBmpUH/xIQkR7IvP
7ausAAoP1gC+THDN9MJrPB/buGI9BykAzhbGlBNHawBDtY3rFh3iUEXjqehagZFu
t15+IiHjkqJ981YB9jvxMzk94ASkf3TvSz8CEiniPg3MWnXvlHJiJmVDrcMWlJHj
Vh7UqE3SA0dLbKqY0yIqVPw2mG8fBDRRiwtoCsYEYOX6SdRsyJw98liA94+8JfR4
HOGKwp1FNnW/NTje/O6zgI51UARwfpwUjzetiYNAC2/Ld8AOFz3Gkrk9Ws//y60X
0IGYhBVNS/kd3F2tLu6Lg+pQ+JaZ1LvnndzOmd4xFKNKwGgSec567tsG1Hl4qvi3
nXb/HL3w6qMQfcpCVpCOb6TjZqi23POp/A22zQ4xtuum/+6ZMymz4RNUhyaJUlo+
J4z1ICNsVFv0FKZlrlMGu9uOPj63ARsjqdDwBjt8GN6EYThJIUuLe3dwo6hY2CCD
7Ncm1aUOKcwnK5AwagkNhRwGof1EwwNvYTmB+y7pfyPfiJ6uJkjEv4queSezzo01
8hrgPq0+FiFZ7KcIuzA58sgguXYCbiJW9ZodDiX8TFf1aPc4kV6YWFz7OYktnRMR
RdNqjc/FUymw+ZSoOPOvmTyFIAKxNzX2+ZwILRiQahg/MY0dP0bySzakfV3qtsfB
VpmvTp3RFTDvDKXe/kSMvCLX/xufQbpOlf7p/4IiVj8ELsWHR4Hhe4qRLTPYCQhl
U/XrEGEaxOgxEKSOSdAaPc+3VnquA51wCD0veOXhE9rEKXJ7vjYqvz//ldOlrnvg
Gj0OXSHbhaLVy1pqfFmC0m2kFTQwCR80JOheCYtLIpI+quUJAkuW8FLGz5ZUZjB2
wW4bPBi4TJW+bDOnnk4ufu4mIiC/PTAFJC9Y/peiNP7lfGfKrB4A6YBcwRCjAnuz
+/JNo8AFeYK8tiJnYxX5MxdVe/Ip6EJDgXramWeUwR43HDy7kqrD3eeHMwV/G7Sc
qvZnxzva/ghZopv1Uq3UgSCFWVO9TW9+X+AJwp2ptshazGdZhU27Qs02z1j3cKR+
6X3A5eLY2g2ySOlOLlFYcF+JnMbvn9M/Iyl9wWdnRN/ukwVW7S8Rsuswaq2IaQlO
iBhyMJ5bqMpEPdT0stldv1LJQqInUJK0pp5ncQ/qRSnsG4b44wbb8N9gac3t7yGg
iSYPn4hwMQsocCyosLJwPcUHE5Ywdfc0T4NHO7HYPB7VHzvtFVzTmRFZ3JbWtauH
2VVd8mCuLnzv36q+c2QS9zKXHT7Zq3UPnBfr2bgAP28Z2ER9wmAb5SqmgjMuZESv
dzAJZmO0JeWABDIk9WiA8qnemAujBaMZGPDEtmaBuWSpVRZUuQXPTFXIMRscr7Nk
w93EbWgBcA7UYgeZFQW41x1+U+WmksNqNwafEASXtuHftoABA4J+yzkY2mIzzjcV
qQpAc3KGrAFBYZjAKNSfd6VqoNDiMJvCCAZeDeIRJsBha0SJJisTLmPGNvFXOZ8q
90PKuOOt0c73u8bsYK1Nb9WUV2LIBp0Ksv6yZ76i2WieX7BIB3X0eluM0LDKYCU0
oHTJITf1iMoOMGgq3XRkRNgcUisPRNlu2YtDF0gtPFMFNdPLUyGotnJqi0vmF9zo
E4vzi1P18auY1oDHLpeW7xgWO9hx7EHnSFoL11FBUnj+3Ctx9cAK6qjy67NHw6V8
ixiEL6dfRoZa1StGfqBWo3voRXaR1e9I+ivEAi0Ilo2yqJfKMKGl0oAFjTbPzICM
iUYmbtm9YUKnCuIS9u/TTcbcgKFeb3sMHCVQpTX1+DT2mf01ZKbX9Kt3vDFgW9Xm
67ESa8xghSNF2m3hF+Xz4S9gI32VBURQ/DqkPCSErQjrwJ62hJF6DXD/aPVqRhzI
5Eo+NmWdxEMDoT3tRVc2LrzoWd9sw1hU6NsVmt7Yrk687TGhVHRHq3e5QA6PO3y5
vdljmp6zPqkbyBQjjZdYDKHF0jiY5pYjAr93vSnhyvm2pwfJUf1LZmGaarRusW1E
Z9T2YxbpwbfuofkUtveeJwRePlhCN4THeb1Ptbljlbh0RMwi5k2YzqNqFd9RZ3SE
NTkTxNkVBzNhCq0Sn+1oH5Ka4AvhiWr7P4YLZhoKXCgw44ep7tDb7SIXPuwGPKH4
zq/5T0qSdxnRPNiYKCdk0bd558UCv0FnSgA3pKyZJKpbhR5UE25ZjnHRBdICjDut
GdROrMSD7hWxguRoo12m0KwAuCQuY9mOHdP9oerCbumun/wWxMGTC6yNnkOZ0sDP
rYPqXHf+NG0ducGNv9CdlViwuO79JXeHVwGIji13awDWwdzVjfEF+PsIW6nj6B0f
qT4OevWg59K1r+CkU9eCsA==
`protect END_PROTECTED
