`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kfJJVMUoq/I0K4b1QR0xNFUvw/usmHRDwwBxHIwqCGrOLmTECULSjhC1RE3HNUnz
Li9oCD4/CTk40Cs22Vyprp3xBD6uar4emCbqycQKs6kuO9E7VwurEVeQV9cpDL60
Xo0xhg2Xo5HfcMYfVoZCgMIii2a/VRwnfx8OT5amdcjx0cYZ1VH3rYKD7Pz5cnNk
Xg4pW9Azp4HwK2iwWqkppmlDZx93ERxHD89vn2dg2CtB8uds2U9+w7omcG3oVxMc
d3XWWPZJbZAwlpDQMCgq1A5C0iACP7QkJiJa0pITzbDdlDQlHqkuh2HB9/YGF59s
o8xsiokwgPVBZJb+Ibd0vWf7shXJ51D1IQbH3UsEWLDsK9NI+R38hFyAbgB9aY9t
jYv/2z3AoT5tPt0RfW1fwHiw9LFCLRXclLpcDTqbO0qA9JKSOEssBwOfAuhbAs2z
GnxsCkzu0AalEzd6ko/Sh5gx1gL4Yay/2wkZd59kMZPvil+BpzFxlZBkhZaODzVY
Oegp7Wo3Y1niLpju0u3NgSLO6DGNBene62c2/3K5Upkeo5g6e+Fzh55ychYmPIgl
G3KRyCz8tVjBSir3QZTJy2hIqE9RJUpL94rs1vUjki/4BKiEkjsxa+ihhU9AlKBf
UuJYqsxRJNk7zxvEMiXn0VjMbAfQv1hnQBJ0vBqhnD+WQuylpkwiJZAi83thSSRy
gmyOREHsf346ly139W7Yyw+zGOE1dsV95jOEnwbXurtJ4A1zgbN0lJtMtfjPjQNk
YsX755sbK961+j5VZo/UyrpdpPj9BZ9RJkHGD5pm34hDbiNPKw0RcPxfFf0fOg5y
8VOk8ZuaTdMx8n8NuZoAwyHAmfADH9SZQLgk9zFxd7t4uaumg+QVlch3WVc5ugfv
`protect END_PROTECTED
