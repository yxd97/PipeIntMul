`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NyhIrmNSb/fIjy2aGDeCzrx4/qXsva/kMflUCkiawbtBSBowinQiaC1cgkA2oxJj
G9g1s5PDliuos5VdrgFMVs3V99WCX/rRF8XXwqeirOutqtXmGl3X4u8Mqn6ZexyY
DJC2yTipTkwlg0CWO3GKvcSp3Ui6HubdPq63npDZeg3uz6uj0I5sgWCn9rcH3GTn
XWHzjPPbwzevBGWPwA1nU1VYDtc3yQShzGwzVWGu4jCSVnjApZ9EgTDKNhdktXM7
k6xQQz0YWnwvzbARVyzAQaXlTe9bQXBdQV3mTooTTSRLNoinfk0th/yd2O3Y1rJD
9lX/bbnA9GNwDKZjC6hXvuD7myRgZi2we563gzfnWFkLDNB7Qy9TBJeQikkwK4lW
9SKL9GfMWerqCZoEUBbsyQ==
`protect END_PROTECTED
