`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1m+RVxnHM7CFPzY6soHLlljrYk1JXnB721utz/zmom5VdbC2wFDAhUJote+8L3N
lWcSCNm+GB65DIsKManIfhqfg13C+8T8XORJIW2sRBirFVqUsxSou15OfFKZkxXy
h3CDPhVR9CIXvyqdeJhVd1me12Y3dVxDSNqwA9baBvqtafC5v4E7FDoi5jIHZPWh
zTRx7WHfIshste7aiKeEO4eCkO+7NthbiF8aEGoCQzilVRkZkWqwMsbUun5jFCIb
reucVJIxqsAyYsukH5OyXA==
`protect END_PROTECTED
