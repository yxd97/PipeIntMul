`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uHyEWmMwcmk8NLx0rHNuMGLwjeWTchGS994yJ0N2JCZwY8lfaWBCuNGJHhyYEduO
x7UR1Qn+7HzlIe4TklrAAJ+4OgJgLA0xsKC8DNUpTRhDjFtepeTXQdbfaFlzgKWH
b1NDcHa2BziDQHoko2CPSRAb7lf4YQgcFfGSUEU5Kz3RCeGsGMOsoDa1+Mo1rIIu
QKJfSZ0J8HTgtVMwWMZMPiZjUg/PZCo2z7INwGYudj8uOCcR5MMOoP/HKNyyT8I/
7smmiWxCOP8MwCALIzQNUT3w62QJr+2r1RCGGcuxMqUZRF55Y4P3c6PF9OKuzWsG
ZFe/hheKGf2Fjvq+ydi+p4A2+awLSdJ9bDcq9TAOGRu+JHkxWQDceWbobfwOgzlE
yBwkA3EWD2WjTl5V7JbS0/CUxZtl1+QxRkmnWnZBgaMYSollAuQo0hzYYuqTjXTa
qUW84CJsDcyhgwh3w4DF3cUxr+2GHW9yPpP9QJR9+kPxVahUIPo0AqDeU2T7Et2g
oaQV7ZZJMXIobEYdqBmlszy8Dl/GXTB6ui8XnhkNX7QV4mx8O0Fx2+r5fj8FMqRe
wzZ1jTwJS/YkePNG8jvCh9PQrpgGrWTYtfq0lg4fPDM=
`protect END_PROTECTED
