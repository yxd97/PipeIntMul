`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6wGwlvcbD8KAkUq12C6Q5EbOzPUmZ9xDGAbUnWLv/5TxwrGzhDpDrQfR2pxFhCoi
2uU/7/6lbXjEvyX9G/bM09zXeW7sLEwFL9cutNGsxFuO/Rlc87wcaUgdfujtomJ5
4BTDAcaM3+q+Ai6Pg9A+Kbbn+vYqvzMJcm/UcbS98vmaspugOqFs6e8YhLzMCbWw
I/eLr3xECZ6vs5yzst39pT2hCMwvoElc0kaNm7dyKNEprhC3Zbnb+jOEg4QP7tg9
76BTr6ATmE9I8/UrobEPA55Ka8wAz5r7WCKsnX4qA8gAt+RtXP3KTZDqYvafPQks
JQZPX7uwyGnah3wilY8Z5T4KRQtM3nCCbjMhvICIo+olQS7lLpy58FVe+3vFAk8P
p9EyLqBnJTlk2mXm3+x9Arp1CkWaHimxZjn10H1x/SntTVZsRuA/R0Orlfl019UW
a4CdDDGp097EINdUbe5da1XMK1MRhJfdTTbpbJk52BE+5+CYNM+XUpv6wZ6Ym/R8
5+6anLVL9CTIpOzQ5zFKfjA0Lip65XW7p0fD7XM+RPQwF7Qx0AWExK0mLoi82yf3
`protect END_PROTECTED
