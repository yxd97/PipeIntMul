`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8b31ueYBNkzmGDv1hUDtatKyN8TyVoKESQKDfnnms979QrHKppxuEyq8WFOoZzq
1+0jGGjlx7yA9Cpsbp7R8VqB7nNkuLV2EfvNa7I79r7vuPWCfXzU4FvvH1Afhdjz
VAcfuDBG5Szu3JZMTMZlc88MST+f/U1jNY99jFEUNeYd9SYiMmyDrqXxboP3c48P
rwkFYFOJD3P+Olv4lq6tQmTv5QKrfUkrD9Pat2H782qebGLhgg3DkEI93mfFRxWf
arQPj+e25pqoPWJ0G/uX9D7MHR8flaf4pjeNbnriXP3JeIQj8pb4CeVLTy4ujU2n
4a4pEtM8gaWmzyEadGp1QF82CexicGelha9c7BWsnqf/74HnUyzSHBlhvj0Rc3E+
1WCdCftZE7YXN7t1FHy4nEocvl2EkEu9S9H1ohXisM/m3vkxoKb9Se9TDNBpBtcr
Jzw4SSOcWFStnIq3qK+Ga2brI5eLxTpR00OHQGOtWojAD/3eqPlxnI4DKzjGZjiS
bBJtKNeNSCf8h1J6DV2QklZsZpS4Tg2ODuonTJlcGttxm4mPeW1aAO9rx5MlvGM6
F/ZpA++jz9yMey/1jvGT+NWkzTK5rX1EUfTb1qivgmeeHxrfnMRGzzlWIXR07cwJ
wmNv9FN5oDUlvWmc6w4CcbxEwhkBM7XaOLJAOLsae7eMORctIQgJe389PS2ZJ1yI
Kt0wcP5o/kJ45Z3mDvoDXB/j0th69UKfDK7JV5qI6QNKtOrxxVixdz6YH4GIb7+J
xfDPYNv/VnKysweP0e8cwPGBvKuPPlyBLuc1idvz7f5s4Zm3ny9Qv93CYx7uQEoJ
YsgcswKK2XZZQLdgvoRRRtixU89RW7qyTYxuvlT4gwfDpvF5F+jTTxbx0e8wK8Cv
`protect END_PROTECTED
