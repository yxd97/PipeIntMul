`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOdkrIH1Ns/ckpvDO66asIew3+30o98IaP1Ru0z57Ivc1DOPx9LlkmCZuUMqkSQC
1Sy1C7J0KFJXNKkmTn2j5GrGt9t0uQIwN6CxHzcpVegwcCpWsnYNN4pyMg2GlrBO
jOQPcHrHvMQregPtMjkp9QHR14Dau8XpbykXHwFLSJVXaHlae75SGDvAsz59pn2Q
eVi2qzENN6Rsqr5BNUUMZ4uwsO4LEe4+5G1D8cDbOS8klWQLgFiRfRmSSu5mjzmv
ozqZUq+gtVqlf1IbefapcD40WwlJyH9jpjoAUCazX6Kc9ksUhI32vifLTyATzj5o
LfN1/qoCLS4bj4ui8oZE/FyovEIdouAAkkTckuWQ6nayt/7HbgyoxeQpPv5v4NsL
uud1QHHgVU3vcxXq6WfTosQov6cO2pG3e3kTzFazDZBIuwrqXYXNI12BreG2oUox
ow91ZwP2LskplNlZIQMHGt/ZWTedXU2auhdN5LC19z0qzmrYrIKBQXlsdDcVW9S0
Plnc7Y7Fi4yevB++IQmpxXxryRGH4UwN3zhwvHYvHR4qL9Yh9itPjGdRca2pEXLs
2Kcd4iued08HIXXwkRCqNgwdXYHRCY75tdg94+4rN3oEfk33UMGUzSsX5Hffzx65
k55w50XsmsNFiT9VKGww1Ui8mZmMp8mZqDCVg+A49RVBAdmXgrPcPKCz1jcL1GR0
dZ23zKZrUm8LxK0LuoGXQG8aXLNXexJ/DUMKaxUViZe07ouqDwK/XzzcGdQTwe8l
ZdBNjKGJrTAZM0Cc+MBPMG+IIEVXonoYUEgLIoKJ4yDJSWJWsgmxU+J9Sq8efmL8
EsI0ev+U5SodVBBxWcHkHdnDmVlbKts/a+sj52DZd/nS5QHznEE0XKiD9XzZQCgH
whdw6NQOIsig3JaCUIOOIzK//6SROvQI9xe0ewokpjh2cDseWrgbc0JcPUfgYBLa
AMucv7PtqzHahISJ+oecc3VMeY76pwtH5Pdtp2ZCJPnGShAbqfec6dC05JVe5oCK
BwHLFgBKDmyYwWHud7ANwb3dhCdr5vAnjkBMMvJqUt75DKhCxYhjzZGeynsprsx0
06hCB7JdFaM5IA9UFgFXsZDpjj7wtaVjiYDnPrtyJczXDaw9MdsptVixMbrcc2AA
08gfjQXxXItCShZIxu3jrBx8puPxELO3UztNdNqZMQOk2e1e5efHHo20vAvCMlO6
MJTykv+nIsgq/Hr4N1vWcybRuOr2dm6bD2Euz3cZD3XQWVrovVe3P89Bzjof96px
ZRsoFUgsJan2WMOkArxbU47FvQE94T1AKIxDyvIW53vTtnigEbuhpnApaLjn/XdX
bj981HRJAqv6uleE+MP6B3ATKwmWCUR2IktUWjm7eXgTaKgIZAbEnCxJXBwurbSW
opNg2KPT5wE9bkeLU8g7/Viwm3Tx/I1/h9l9LUJuQs3Z5LinU2KldO6Nx0PY6S8I
bVaZU7uiYt3yDPbdKo+D/Fd1hPslzQTqji8vk1+NlegDqs96RdyhtqI0WI0d5gGE
4pOmTZHEMeH3LVr4dqqr//jeX6OZog5VAquPKeSHXSrCyV/ExnFcrVNBNTesIVLn
`protect END_PROTECTED
