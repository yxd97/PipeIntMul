`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AzT/y2oWxq36Ka0YZ1u6Uk/JnFvg1EI8MKgxVhEyWQhZ/d1Q0bIU5hyaHzMSfRyH
ra0ROVYzYMI3koQXCqB5Pt794IbyKMT3DM2d5Kn69K6Ai2OKZmehqIlchHlactT8
WSC2Ms+resrRBMVGcaUv6SFSZGGHaAKDwTJe1hEg1jcMg6WCVx+etV2fuF2zpJ18
BANZ4HWeXUbgGYffqVzGk3Zvmp7RQlDD6MryMlONQlkYdhgx0zjsvlHKtz9+ZV5q
AhbzRfcMx1g8uQlloUY5AEC45nv+8QLKFObUJxaiY2U0UmBW3nZzB+3LBTjx/OG9
buSssFh6r1SORornmXiQMletpgqBuAY+87VeZ9GO/RyRJhY8TeB3o1pFj7rNkqz8
3Sf8MQGRJmYVqFRRbcbKDIkS24AMphv/ubXGPG/FN9XaL+i8nF3Ka71nrasZCKJ4
/nr5rlOZqpOPObQRPZaYCKVFzIrFL/5Sga1H/Hx3maat9roVN4SNLBWaiYLjzNhw
P8YDucBrDUeIx1kH6Pm+BSZXjoCo2/FNZSMH4pcEJe6AUAPW0gehfOyLkn3Is/Vn
bcgdx/IvKlnuQgjh6c2GytckJtsbcMmRmx7IocPbq8wTGMIMJoYPmZbzCo/YcmjF
EuBUfOm4G7BLsqy+Ar7OGW/YalnnhHsqozQmYltw37/2ZRGSVzV8VWGIrFsErjDa
jmTJMr2SP5SgiyZLLlD7EPGrgvqF4oALDUtoq0TaJTPAe545zxs9WcrPnItnwNgN
dvy6f6zuPpNwf+1N849/2rZG+Tdl7eCiuIGde6UhiJT35VGlBwmMm0+jTDhhINJN
v1EzqxFx4yrEHHCRHisgo8UdRXtUSlercRiTgE72gwq94oa1ChUukjnNzF4wab8f
ubCTUqbnVnT8L0kkmVfPm7jHiLG5FdiKGYF9ff2gMxCLmbeC49jtQVk3bxQFnwAA
G0Eis+biAdoetMjTUYvMd1fdWyZ2sfonHlDAanvd2/0U4VT2X7ULSevtguiV6dbv
aljxXShej1HzDCKvF3wcpY/rvmlb5bkJSkJ0F1x19hYn4lOew3S1P24oj7uU7Qdb
RaxVX7YgSZ0DJO6ZYyV20TVvU5rGXjoVbdHiVnZJ7NOE5t/H80Mi6BsKDy9fe/VH
ro+indd8d1d+lB7i43ulWQfp+CJpTwhEnrQAXvEE28P3nM4dHRPkttmy3UKjU/gE
fBJx4enMRWdJ5pyfO2XWLqFwInhZ0r1ESctHi83g6CTdgqFY8hbcfA97prQtcTaR
RY6ANXfeJcUCShhoPQsBHSx9rM2ZszZC3A2TE/QHU72GTDJ8SBWZu0o+vSax80h+
jrBAnWjBUkPDtrKGiCbWweaZqiuW9hQdKITTDOdDsOEd3sU7nxxlMkiqkvgXEHop
ZpuErmWE2USBC02HHFaSBSUzm1kocInQyXmefCyg+ftb6p4jdHV6UCtGtfRnkZkF
F0Jh6TfSUx2aFSk379rUermLvhix9wj2cQKCcfa4lhER5WJTHc6djz2Kq9+NwMvE
L5YrCG2koWntrhDMTMipWqGf7UqtrqALDp40nQh/NsA/931vkeWU9l1OeNjdk3de
iha5cBEeE62zpCwSjLJcqB0rKGH5zWnDot/vNnYW8MLeoTVDx6emCkH0tyVOKE13
R1cz5YElXqcoN9sgwACos2mvQuGs6qOMZeK1RjYE3Zjti3RCwwGET0bSBNAAfSNm
faWQFJRwUfJ9CSZPk5HlpYErSVRpP58f0chGSM9j5u/vgTW2BNyKcqyriyuw4oTa
nFAS7j0FUbzZklww/JX3sXt0Xd7naDIjQ+4knFVJ41awIM3vo9WtKQ1kg3w6m4dZ
LPmGPGTZQeFa7EQr+Jv3W96GZMkgChDEyM7dH+1tQZ/MMslLQ09KBa7N0zW/sRDs
I8R0EsKEMTIsx3vPfGxzeyGKn7iXx/6DKJ9zeJMBnI6wf4H8c7vI/VzEkQ+sFUCo
dazWxtcc6DpWwBbSxxcaEvbJa9fdsw5BXOWHnyy/n4656E9vjCPsgwPRfOc27DmY
0QyyKvrSLn2sc4ZpfEPaNTfc7o6SQIx2oCsxQxk7oN7BHNIJoNaTKfbfQ0a1+iEM
SsIeRxpr6tnXb4YDSSM0fVbw5NrAGb07bgJ9rM0dGzxHKqjxsVgqszCpNAFJ9JOi
jszlcicL5QyyGiD6tJr/iH8ProEtKhUL0vr7Wl66xdIku7kPch0dxGDyFzuWriMg
Ms/VQZdchlFWT9rTMSlz6PejyabGlhGgzuFAkcY0S74=
`protect END_PROTECTED
