`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMGH928jjCNjBBBSuSHUPN30gCwZMcCbdkBZUNu3WdcFZe80cTxUe9M+M5tO58as
Jrivi5RNnWjiVMEkQXQ/3zoU0bk21sno6DAWuQifiBVoJz8A/v9Djg2XmdzA68If
G8mT90p+5VGxgikg579jvyu/Ql7QQ2QNhDGMrO7dL3spB7WcSaUzgdVUeG+WaCVS
xB32g8tJ7iKhTzVO43x6w1x2ANpkm0sU6YJEqEuL1LFIJcPoN+AEd1el6/+QcsBl
4Sf3L0hzhH+jXNwvbUyongMUVCj4QuG2iIr7kblkSKc+QsrGya7usAfwUze/w5Wl
74BH0HHZszlBXiibUg/65Ee10bAgL3wisjht3B7hrtUGtWtjhEW+sUttMp91B/7d
Uxjd+Cuf+rBY4NLxsUXNCgCZFy76KbSW5b85eUehrNTmytaouaIYZoL14prhvYG9
kAxoOaApl5k5plR8n9RaYB/DLMjOxvI9aOBvPxyZ4jk=
`protect END_PROTECTED
