`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7xlTBOpxo7U99Sdi/KU5Up100mLhjVdTHy6ugzWjMhqYK/294I/K5VXZf2nrD2Ex
Hy1R7e9uAveawkn67jJ+2Up7T/o9QVauCGVU5uYrnJX9nB1M1WgTklRDpVNDI3SR
qnO/Zc9oqOfLSivb4NDUYVsTyqRkXvzfZbZuZvcBKLrnAV2a6XbZjB+Nbz7p6Bq6
n89eMNVMNgdQK5l3bqgAEVzLDn7mCNSZjemYY7vcqnjO1UIlbjDw6CHpxnNWXENT
iozc/SaUqPPjksUGHlHyXZQ2NS6rb2DTuKveQohVOduKdfD3wlqpA0qLKgx0HbW6
YPQEtIb9gW6yTHT8IL8UvyfCLWqrWGyJAUlMi7KMa8nQDKCM6Azmki2tsffk4VIM
AX3jbr3ZBUnlR38W+EFRGg==
`protect END_PROTECTED
