`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoKGFGjlnubfNRWVQ9CIdiiqMaP0Ii73A8jaKYVgrcOfBLePSh+zjFOZM27AFWy5
xdpBrg9ugBUKcrp45l6P7SVfEMEnPnZ8wcm0Nvc5mm7r3mG/VDtfbk8ySyuIanDi
00L+9l9cUCDKodkFYnVzv8DjWmwFDyjePdx815sbkPSJ5iEwcwrRo+IwNQeVsrf1
LKzgixgbK7YdFZdOezpEHjRS5/B5JTQHRA5S6L6c6ggOKz3XgHkBkoXD0PvjsjCK
rZa7PTW2sk3sYgufETAoT1CMCPAHvCMAX+OjQjbVVTUqbTtTnwD5LlDHRBd6EuU1
hzMQnvvhGv7swSLXHWTGeboTSyABARj5o+bboKPYwVVYmxr++M1u0LfJeadO+OmM
gaVVpWFNymoNXLI7MDIpEVRcv/Zv6/yuaFtBmxNsX/wrFM/ezMDKP+uHfsuLj+f9
ASzOZIN1ZWRVQX6b+wV69IItiyH2YlonSJwOZEYklAMdGw2QQuYlooTqDxMZXOqM
30Sz5SQXEKnzUez8mECCT4sElOJwy3iPGBxNipffdmvstSQDYzpLlrh6YFr4V5yQ
pLX7YUXW+Aj2Szh5zgwk5fzga2KFlxYpgnOKxLlKuFwV8imz2r4XHaZsLpU6wvei
uGXfKlhQFhLnVKXZPprRmUSbe47e8Vy1Ww8STSgu/VZAzZGGJClzOBKtE6m8QWC8
+DcIa8nZHl3hWjAgujKbR33yE9MvnhtwfKdNSt14TXNzJeSTK3mpLTmL0fYv8Hct
NPHNuK1AEB1Mzpuy7RNrRxELiXHkNcS0RXWcn97mm1qwgNGB6aO32h8pdP25BB/j
auELYGloX0urhTxDED/cdKC58pmKE/3Gxs7rFZEkc8vWBydlPlycsoW7sU7O8xzw
ygshRQzr1jNxpBdzRbNRtKXV5kF8eoJ00nQy6+AcjxGaq1cq2Ga8VNKq3c6lLsHI
brdr6RJOHlRzJg2kQFzCPUFAd3Ybo150GsHMdPtJgSzwwu2eMVPgDEh38Aw60bz4
r0TB3UUvzgPMYSyP58DqR6XhaI3YtnwyrgHu6FacAHGKl3s5JcnHNOMO1KQ1KaMi
Qt9ZFSfAiTIEYXXHPpvpGTNaRV+HSDIbH2ueh4EkQ7U=
`protect END_PROTECTED
