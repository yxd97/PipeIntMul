`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wcpF/fSMXW967yQaBN6vwjl+5zNfMkob8KFTMk3baJzTGIn9AnHbHCsZ89lLAkCb
mRTStmnn82oCcZM1EZeUGx+fPY1xg988w4A6wDvzXw5GcOu8nBIenbeeRPx1KOrY
NOzU6qSGE5Tk7FVK8iexcF3FJEAJ6vFRxaG83N4oJxRZ77wHQleyZytT32Ar09Nb
2ldkjbjDc82hynMxx4tdvx1DwR1olAictGQ39gI43fK6OIvgzp3h3qC60EPDv/rA
v1AC4zliG2jvb3+lQGWijIIrmwbBqVc/0ySeJcCGkxhPF6CM/zC2kjcLQad227nk
ffDTWJtHU6YinS9HePi8QPbnpRW8L9t0ENwK6L1oNR3Z0PxBO0F1Sd3OHf+oVebC
x8c5J/S8huEdiCb1kRdlBQx84IzJOYFfZfhPUxCX/Yf6lRRD5v2UrjTitMIwYgk9
JLR7+irnH49eE+BspreygDdZabnKm8krjYO60f8uXx7ihPJZbbrkl2AmacxqgM2T
5Bsv/+7D9EciYbuyTMoYMTLUzbonZWAnmxE4HKWwgNrF46LVL+z/cBwXevncpXAd
2lWm+F3a4VksiOUxXQ6LGHKCTk3brGc/toalNJrQm6U=
`protect END_PROTECTED
