`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AvpVGZVImBoi1h+gaBTeK2HmUsUOm7eCeIeU5MCqztPKAmpfnrPlKfdQTBDx33WI
4ntm85L4rLns9AEyAcDXVPXr88kkSPWRIo3DYYMM7VDqfYPsz8lZkTFL5dDu1Vq4
jyl38zw+KtxFHZI422zOmuMCghL2GC8W7agea5tWTBRxOQJlbW8frZEWp4txjgFE
gqLaZ6kCpfsCly/n59YnPJRN7Hz+SaHCh6OoccxtZf83P15xjiE5P2p4yGjO3hLh
GfGWQhUGFnr3EBPDjVsKBRuwX/tezQz8qpiHq73TyIYVZdVNRFatOwRVbvc+xZKI
IPGzMRT5iSkjKOu7WR73Eic01beryMqB+X6lKcqt4ggzX44+W/bay1VRh79UnV9V
Mj2LRXsUqdVtBfTXutzeaVgvQ/D6a3fuQJst3+Xa6Ps/N6nEe/IDViZq8I31v4Yj
WuNHhqAgYPNy7tipdiTW7W285GmT8ZDaC/7h7oh5WVtt9fuwcWKtZnVbmcyIer0D
rf1sU2WV4QnW/5Vsfe9FuQBeRblaogbu6i3UwuOBuPNF0F0BuPaobDN92xcxBPZW
oCqImZxO3pv5r/gQ+Z0GTYJE59WJ7HgsXdlT5uDyLNuAYs8LI4hV/aZQoYZsbvHl
svcIY4wR5SX3no1PZNRMdg==
`protect END_PROTECTED
