`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p06cG4nEbJL7cO39CodB6ya/GEd5qVAQWcADk01PVoHIos16wtV9SUG07BPiBypD
o60VTe8Q0GgbF/9bxmnOmBFixWz9jyFVrpUiAM4jHDwRWszeQJLA9uGG3rCrinor
dqRJbvaNohS4muQ9j4TVlSyfm0l0EuDT6YieoTxP1vgvQuehlj8GBuVjkjWQpDaF
kxs1+K6ieUYPT7QIxGGJK5ii6N/Ve2sQg6tRwYTqB1/TQemU93OdW5/QNpjSyTt0
5ecK7NGsyGTOjNnDADFLzeH6pegs1xwZyk9ZbdJ2J5b15pEWqNWJg6XQEpNbuWQ1
ygVdIuk3j8aNI3V8sz4bQD3kzGwYQ/9z+sbcJfewSQ6Li6UZRTBVjLZZjkWO6loc
srgSJ4AdIo2oxwngujBFeq3a8VF9Ux8o9rAvem8yZKb32pHB5df9XQHJ3ybxD7N6
BjbcT8mspRCF5oe0A+uBWRKlkf7iRlb+GdrVnSLbjXF1uVsJDQwapLS1twJwS0OB
U4wjRNz3vH7q3xksNnIEAd51PklPTGC2oWF+KdtIFWpNTGvrueekLxsudgv4rR+h
izPlvDrLH5Mo7oPAe3Mgr0lNJsQhvyQlFOU6x6WFtYc=
`protect END_PROTECTED
