`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlFg+AkVJXs3320siYjkYgPXf1HjE5zoa001Jhq1lEf9BqgiEeDn/8SAPKBJJ72T
mkg0VZEHDTJ4kWqFR9lW3PGWLNKnXffezMK653dNstXRn7Avzpgi14PNHNG0PwVS
KG0H6lqcAH3AXPKw7UnDjX+eOCEhzXNXgWbH3IU3HMCiEXKbvmYmoS/gel0Ftbaz
pZnPp3nYumpRRT8eHQaIeBFNFUdJe4QwKJd+NypxUJgiwxcaI/yca84xlMGLMYjh
iv7ogkHgyjvlBxVuOz8oYb5pYUCJ5UvUReUqy1EGQ8oKgs1jIF/zPPHSNIEP0b2K
2wSkoj1WibGCsIjw9kZBiPUXMFK+m43gfuwB2GmeIRmwz+lhjXI5vfcVH5neA5c0
ovKFEKRQJNBeQLmVH9BzjJuGOCpkiFT46ZwCmuf5OoJWhnHRnpJOkQzs8O4Z5eth
8Rf84k7EXYmNdIRhNK0WZ63VgdcFz0T5aQ8Fy73M1wLmBS6fEw1kul6nIWVIG8Xq
`protect END_PROTECTED
