`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gntQJ6m2RHRXJ+rQU7QAfOv79ejTC60LZZHfO9HX9vPgKLFrll+gHzQnSvCD/Y1M
avX5L/c7MnV9bSwmQmRytGK60dnRpdbeyWwippl96Ls8nNLCwGby4FFOlu8fP2Ah
xD+UCSULx4uI7v4UKWK04nIsHQz1SUMfsexLKCEdK0HsYoest+z51hyF0LE9BczF
DiqDhEQnPIa4Wq72Oy33IBGwV06MjtPPi8nm5rkMFf4rbp+VHBFtGrFUJOHqW7KT
Y9BdcWOrSp4VJSP/+J8fIZRhGxh0UNdhU2h+VbObVBZjUYOnxCOYD98ugzSLDb3U
AqSxX0nDZbhhD9bTm4DtjONRdVc46wo9MSbAW2EJGpSURz9kOQJ4B5ZeRnE41S0Y
AkZ1o8ZYsJl9T/RSkuiQAxFbxG+9n2ONetCr4TFZwxDOZYu32xgr+dPTt2r2nFLj
pycQCeA2TcF3Tr9amXpI899IQUExJyIDb28CmoswPqqbo9J0Yq/tKJNIIsoNHFgv
GLb24i9NyCZf68niXhnVqY/3ddQ7oVEpAO6H+pDy98AAIzl9nT6RZNxXRy6i2bl1
bobRNUynl5H7oVGnRWp3qTvHIcZ80/liCXTCYNpXcWLkeArfuURXmxj+WxdAxzZR
czndqLhSGEAKpl8Uw5ZYIFxaijle7n/F/hyeNF7YXsjVkpxQ/SpiR9mhxV9YVBlJ
vD3wS8yaB6iAOPLTJPSqMXUkv6Xw8ohDbFZUs8WqV8EDsgukLK+jT2Xb2WMMGjhg
p1KtkBo6AyehfQUOGLmr52wnQZw3x6xu8twvpWpllYJ5geqaDibHRpPhbDYKl4Sg
TLmEyH1ruXCjGJcuElNFCblVftejMZm0QkBTcFaI8Mjz4ZMaXL/Nz4mkFjehGX7w
OSETenoY+3wa4omC6eECh1RLR1tOscPCjDBF5KSX4PxNUG/wuN3ypKM2ivNLy2Gs
jG/d5EXLTo0EdSNnjBJmBZzvveWDlzFeTzMnYSX9ti0fb8qfoqvl6JAo8lxd7uLA
8zaqpFWYlBkXqa6HCYid4ItkCCcdJbIkyIQPftqbvsHDq5nJZkdh8bgOeEW9+DqB
sxni/zmTRtOwYpbjvoJJrDVi5fst/1SeSVBVlk8nvfCu8T7OXGN8RJ1/+103kMGj
Gr/fwd8zwuC9HaL1F3RZGxS6pWa0AkQSWdWbVdqad5LWVff6zMYANZPCR92sQyUc
rpxejfyLayWkUoiDGwtI/a3r3DBdcLVdxNAD5dgzw0vmthMFFlXhSHL1CKgR7Glu
FsK0xd9j993QpktBO+FlOQiCSA0Sxt1sNFxAKi2IsgaVQjOHJ7//tOOaJglwVESr
2dgE6/houLMC4Mnjok657/BH8PxNaikupR9b/LOoJ7hye3adTtSWXmPxFwiopZ1D
3KBImzFuOVWisPd5Gr2OAU7bl/hZ7XKXqKe9v6uY/JpvVU3otw8EsS0J1J4+1GRC
TFbDbUvWYQbR3CIxPWEvWSzCKtpNuzUCu5qlN/z0nShhKa5/u1nb9s/ehh0khK1i
DaH59ZRJI2QhAVjuDd/OL59Yh0ICWEnCDMAGoofbRAgu252il2pOESUlcN7BvIvv
/su6QqHM/6VBRdGPdfJhUqEJYWtBYe/aoJ6yKao7naFuqg7SYfHPAs+gaejT/Yeu
baYBU37TTZMpu6mkiyspiTroW3EXVXsKIdQ627S+9mzUdBWF7f05bukgECxJWWls
VkHXLDfhUUllzIGV/GZeIXHX0PHVa6z4s/C/uA2kvc5xWjPVJFC3Uql+3niMyD1E
u7K/55782xs/qkPmWIo9+/qBeoK8mgj1xU5rpOZwODADpTbeAJeyHPE+gbzedYCz
MnHKnQk57vVDd40sA8YLNHxYa09SIw+JNLLe+EkOt1Yxc4JWxHC5nSnCGZjvxwm0
qF5nmA+bRZNfA4Tv5V1E+Aty3zOxq7hgiMDCq9XLo1cFBRayBKVAUINEYlVWbDXw
Yh/MvQSuWxaGw/g0zmIp9QNytEGWyZYHHipryU/82omjmD1MIoTcb9ZjAjU/y872
+P5b9Fvh7mCMO1j5h8xt9T2AFNzFU1/G1kRxuFF6MBf2kID6Aq6S4m6Cddr/rzzv
Ub6duuXw+Of5LSdxV0iQQyfUJkwj2xJHDZfB0x+js1Xj3reiXuStgGZjpLq/oJoQ
uFTDeRBO6MiU5yYG4oiSRVwtpecbwkjXnyg2vsyDs+WOwshUbiRcmPRp8r6ybc7N
bnxbUvGmIfa2ywRoxOCsJdtm0qJz6gSmiXRk6swaAy9amkdbaEtTWbCE1cxKDRyx
Vpehpyi7K+gZEzTf3iSijkeynz9eFGgKwpIQ2lL4fXHn7nDfFjwoqtZUFS++Gux8
jl0Z+hRWATA2lH+lz9q5r4BU7wRtd6UnNVHbgF6taTv97BqyTC8fGpo7hKRcb+T5
R6m0PZxfcFMhHq1DI6GqdWwdkNDqwWd+W78Brby+zCUrNVK1qhnTUP4C1id3UI9q
A+AxIEoYwsmf2Asx6EU41QLsUZ8V5t+NpWeGZhCDyBRLjZYzx8BspTNTIlqUymWV
qAShxZPG6LTlRQCjqJkJmC7maezBfWb8udn8pY2U+gLKOXl/+7u8yculWR5HWOYG
4vR/qds36pEj5CI+5KtmCrXL8CKJzSi5Ct6zkdiLnsVhmBAQQoQvAcOGw5ctSG3M
IxO/ODzRHO9KMsluBUb71UEesIfS7Z6bJ12NdlcjssrtWZ9+5i7BmSeHap4lI7Rc
kB2ECmX4IQHPkNdIvbptHbX3gNOyNe/iDfi2HYV6IZnhKrQFolR3DhOpF6no+QAv
cJvybvKK+yZkNRCv7QjuThrz9IxYLywv+DP6lJCRjkASKDBPV8ACBVVak0fjeWyf
UTJy/Xyye41ftHU/fI1Hnj7tTpAvdx7K209Jesg5WcTXSvmKmucdc7nb5myr2mMa
4gD+oH7oak2BqEeVFUHh2t86Sk/XmxHX36tFK8oFnNqh7fa/JI4MMMYMBP/t2bb7
yldB6EdKmSsW7L/IFwcd3orKkdjDKgAG2iMQvx9njAQflxXSRRmQLdeK+P29q1re
/tP+eWN1jSTRlTztt/K9Pk0XVBZ046pOwHEodqRIDEhRooFOGBS1+13p8jTwHTE9
Ia7C2bISOvWzAvIVu+6Q8q0ZmiwnTUp8lybT2BPsu7QmR6Lthne4sgfOT+d/aVRy
Nt2+ECAWDX1XlVsZ29MmvqbX+J3cTMS9I8XH0F8112gwiwv46IZ2PTi/neB5IZt2
NURcWw961JIYgxb3NR9x95KI7x7tO8KpYhejxZlOEC6kt14Eyy2XYVc+DmSwBPMq
qTYfkUbmVtq0NLwkad9Dyb6RfY1YTpD06fvCPcpa3gFJYR3J2M4Kdx+VPC5P557b
f6dtiUHDvlW4rBCAUSMb9vyYRAWVD7UyHIOTqltMKHQn/4NbotepSXd3h3ToaBbs
ijR/UBcQOfSUdh7/Bs2eKYziH6hz0Zz4VFcSTEzMW9orkdmfaXRxTdXk65NjTkrm
41jHd/jKrGgpq2mUNr3e4uNRpwJzKLMogi2Yqdakv15ewx01/UWeJXrOOV8T2QF9
wmK89+r2cf6zvy5u7a6OpuLsO0BtQlwxaWlv9Zr05+evbgamnWrx95cIDxbpGR4g
WMeKsgVGS/j8YdQBymeGz5Bf0iylvWPrQLAXmLfMjnaqA0PoiTQSYLHwtG0vs67f
2PXQT+D+dXuOe66PS5J9fTddVJuGAIBvF617PoLU+tJ4qlWACZzN6WCHgdaibL73
sG4a0tTsd7sCg3Zmq5isLDBJ9qmyjYl7lweGdfCuI0C8zkPCqw3jL3DE7H/xeIb3
/EbwWxOOBrIGEKeuHVjCKhcZx0s+9Yhkdj3uNEJq5gYNhGTx9jA757gZ0SwDn4k3
BpmJPKNtsJAGavF1Pdpgd7gYf5F7cPcFdbkkWx0U7yPneDz5mlr15oTBUJCCROEV
CG0J3bD2tysqDKMWFVvcZ9JYriheVQqpjkx+fQ59alDo51ZlLEy7aef4MXgdyAMx
BU8C7FdyMfrVOHdHHj2465Vgq7ZplVbPrjmNF/KvRTDPfxJqCs1RGpI6yI7LGnBP
jg239vQ0zpaE2w81bFP0SDpFE3RGZdosrUcnsqCOfiakz/h2pLAS/xQ1iYDo+L63
XGu3GVRv4Wfu6PzTAeWAZrjD8XO03/bh5E/dhHmkVTbulffHMt/qdV0U0l0skpOs
JdCid3xKhSJ7G2RvDQNGgmcRkgPyfldY+TqFz4hxVVybEV4oJy6HZOfG+Q/UsvzV
SYDp86ytTjLUaEnT0+TGZ1b8AQIQtj4OYlyvPpkZEvZ3Lej2KT2k+Tk9AGs62tXj
zctWxMXDdRDbQ+7ApmPMxd1ihca75Vuolm7lEMaB6J1QVHZvjvbZrxdDS+q12cpb
eJd1VYwbA/OuRgN1VLLJ+bze+Gy+Lq8DPIFoFXBp2sitE3bIPSc8IvAiRJbsINcu
EKMOEV9ZW//YiWU3UqhPZ5V651ALb5SQqJW/3JvNqPHxN8Q5HSKJ+hdpt7vZ1wwz
N5homVaEaMT4uziiaEez0ZAuVNvmFDavByJX2o6VG64eJ4dkOHhe26W9FFDmEX2P
D8K5o08Mw8prT1DxbKuSdLlFM7qvxOztnRsWq9AjG5+itAkXNp+XzjMshKoK1FJP
eOe89m/ynthJESfbUoiyxyeDL6FUBm66i5gN9wpECoRWrJppMqR7cOBhRbLefPOc
qCUHFhe49z7d3XlHBNC+Nn87FfnjFkoL7fCqxANIaQcZ+hhOUReFj7/PLTuDxf9i
VgdyFGeyBvEmbBljCAfyvh4EuDTLKIuLTE2gCYaCiR7GjTGsKurNRTWcksseo22G
KOZP+R7NUgXpHYUXRjFNBlvnZVEPip4fG67DwmAOlxoabmjp1r/pwDCSryPRwYc4
oTQDGARNNNasFxz6wdTa2bZ48Yme3g6UGGzfNe1c1zsz/sQjXATc0blg1kqzND13
8c02yU5lBHWmwqvwcgEbYfmfFqjXXY+nw0sJDfFbHW6/hqt88SIkCq/U3m5goLay
JgexZ2Q90gbgNW9+qRs32seBNE5gouscs7PxnbqckmrUV5SEB85WraAu60+jUZrq
hzybLvN2PmUgkk6lett1VVxB60ct9s5nOcOf1MgY/Yb2GxSImYAngDKuIhCjFH7g
Nx2HqRp4Pc8BAfzYL7wM6Dcp6fDWt/ZHIyF/6zro/ItIuKMxwCJ0e1A2J/+ohFOM
067+4jlaAGBNgaft7MGRHXxyAAf/oqR6E/Kctw8MESvP4LEA0NZKYOiXDROYtYOs
QWgUrjuBUP2opVMv4FmKKtJwZwHE7PgnGu2p3INsyH7ZMuc2zO05zWA3wLUkPi9P
G+tDrHVn4IEsDK2OrnTfnStGq51EpGDc099h6Ffe2QZCCW2a0a3oB8Y4O1J7cDQl
vWAkdyv4LQU5C8Scp8m1HLWnRrVW8EKPfOD3zg49MyJOecLfUTsT9GVOQ5AVeF7P
w8Xn/0P4YsnZfjlhvm6oHepv5UAr5y7ul7HAfALXW6KFTiPxwSww4vL+dEaRkjC3
t4soSqKthiXLJAO9qvF1cn28sIZ4G/48Vj/Fgvs8In8BeDTa6533kb5LREBMr4zb
IAIbapdryW32mFVqIoiV/0WXIAV8Sx2v1kjVlOY0PNV+N6XBWY/uhUcDCsbZWgv8
5MD3SAWhdNj92B7SXHymtFJuvAF5mqmLq3mH6DM9rgpsATVYLRwyj2Di7kvHou+4
25LdnoFS/TbKkog1GwSK1PFu9s/coGCEapNFJ6p0gQV/nCwjAgxox2Lw76KqE1SI
79YA+fmxT3oElHPcQKlbDDvVDiMuWO8tUDNL2DHZPngrJxzV2zRof97XwMdx3uNH
Lgkg3St5kZR+n3h8Cm0ddb2QUsWVEwdNGpJJxfureVgxDyFduU27pT5Fc/pvmMPz
clcfrO0T9XtRJAriBhT7PDmbKClue26BNVa6cqJ93Z6efEQTJ3nqoxojreuMvF4n
gLUpFGwBO5OvSIhq5X+t7YeXwjUV/7aGfZSdIPt4C4t+koz0yM/Ke3kqC4yFM6wc
d1HZum6AaLfkq8yaF8yxB6WIaXYba8UkU29V/YeZI6mX4my9JnEbqI5rGANhOdAO
n3gsmNT4EmXAsFsXASpwYDVpxHV5MFWbRvh7AxWcUrwJ9HBJnWomP4dkHPpre+xC
1m6dRjpSX/z7OiL5/ePBa4Y09hH++eE3UgcF5bXKuW4CkS8Nd0e286No/pxcSHPw
sGaUqEwzjfJT5hPXrmy6wIGOoUOl0Nk77+SDZqPakkColxpvbXJiYPfuC9gn/ZnE
C4W7Qq8HpBCnx5kwhrETwALRH7C0jCc+AecPmGKNfGXKhEYF/Jjd0SPKMmBunZyc
/IZF7OcF7AfFOgT07FAYm4yDBrmzaaurG4rq7DRlI9VsDqBGxLKlo/jlmv5DuZ4j
MyCEofAtkUfY/aa4BuJdFZDuSfAXYa9rBkvFlKfWDyw70W3f+BQCqLqmr6As9oD9
KmMZpsqH6Sb9g7AbyvfJRopQVpt/W3rhVejmvjTsdwLaipMksuP6l2JjV/NOLKs3
LXkOYbg+BE8fw0ZaTsoKOMAmn5RjeMY+X7MyuepSclMwDjjX5JDuDTtithnWJaq2
LLLhbNr419w3byv1tDGtODUO5aTM7PUAgfnPQ7sxtRwY7YzZ6/kX0nUS7tHXIces
lR5ZrR+k3Qn/aIT/TYp/CMZ2P3tKVo2Ikpmc53GsPioRAaGwgXV74lMPKdDjj+TR
kmyWS9D+LtS2skzwlI67/kEZkmE3d2gkrSsnr/uAJADS+rWiZL1ZCxdQGK3/Qr6H
dikuZp4ZjrDp9rF/tCj5O11NpYiFXm7m5zBsO2jZwQ+SUC9cUF/9z9If9cR78VVN
LyqWB6X4DNhMCcJcid+uRu9RCmfVDWYx35H83QCSSpe/VbdJEo361DDICt4MwtMf
4OAx1d5P/pVhtsDcyYQl4EiN2PjOwwfV4dB0iQkkzqZ1/Z+B5x+R+GPmmF6ZhE8W
Q2jHfCfkLt4lbGCZAFCE6IPHGwkKnb4iOgPZf/MbUYbz8DqSMlUF9Pq9GbKdwM/s
Oo6SlwsQEvMHMOi73C3tMly9JhMCzuvcsRLIRI2JDHTewtnn78onI8I5GFOn9GEn
Sjk7u5NdM/h/sXw9BMrwnqvuIcCicY7GawxCgWP3tACvIcDejqkp3+4ZMJVZlPf6
5WvExV4hAMP25Bk3gTnuCAuiJSJe6ouL2Rlfsjcro8g/uxaElS2TjWyAzCNHTaV5
UXrYCa+U25F2gClDoJ4+TBXTSISGUfmmUQGKOJcVEr0v+iY6dy4dIpZRfxHzlyK3
EUFIb4uz/44NOYyUqSU7nUHJaUrxvx+qRA26sf9jvFir9/4dMv2y6xEydOwDsQR1
TRdLJHNtKxOaMgojg9Qq+vNhuw/NdNcGg8jGQw6TNqjDbXUKnf9CAfselj3WWypO
NdHzvKICg1SnyC3+L7CKlH46W2cvuwodEk9stCsBcVZ/rAIzADvfVeq8mkWSmOXj
ITLduXDowEQIuc3Y8O7hiu9v5hUEtyk5eqBPl8/ftv/jHKymnOUw83V1V+iAXzuL
sUpwMmmv7JN1wZHAeMXzVyax55gXO92ZUxcNl6etJz5IBn7K+r19AkcAI5+FLxGT
qJ1I6TlPyxYnfrSm3VOFxxzfGQO2sEf2oy7uck0u/7Am410H/eTYl/7VxUetXRj2
atCI/T0sm5zG0odo6+Yf0mMoHj5ahNynlB5Mwsxr1Qih/h3a+Q1JQNsBRysYmKfa
khF2T34+duhMXgCpAHDf9o04fevx40D08m+/siBVLGx9L9dy7+NnBBRqAcFGhKTb
jjjDAQ4H+RfmDN79aRXNHr/NQyX8+6IKNIrPbpa0gQbtoV93WQtcR85A7AInP2Tj
XZ/8ZyI/3vLW8vJYDk2GMi69TJWhqcEJuLULjjGkv8oWTNshZ2zauAte03ud3Tfh
tlUFujwi9r3vsX99pHKUeWuk0i/yeR7JmswsK8l7tr0psiMf9LiKctP8avAmpW9t
NDzStlfB5pN0pYC2J7bOO6LrWXQMrhf1K02I3CZZCZV3SGPd6JtlV5iMWHVgDW7g
sLdFJOXo7fwnkXTN7weYlraALFM1tNllvDG0sVZFfTW+NZxQ0StaG1tV5+iJSIUv
R1EGqQG3Z5iHE3oxX+n0V0/CNwjJhH5uVP0v1pKf1Zk5eiVI2j+9gNWYszzn4c0Z
qj3a8Eqly0qmxc2LP99GbRT7z1kUA5TGCHhK85MyW855HmuylhZ+cgUz9ZkC3q8h
NnOzVlUFRyy9sv0ZkFWgfJ5d3OcmbHq3KlyotnQh8B+GJEQFw8xpPreuLZoIYKWr
2cx+F8x95f679+0qEazSvElI6lauCVtkbJov2lqMWWK2xNNqK+rCSQrUrsTlz06P
J8kO+oNPFyk66b6lMtk9Ruh5kZWbKU1gmwpV+IuRToBbdjonz1kchGwvpcSHy9PD
tgXtD/2yk77GZTyWB7fXU0/pj8Mpw4+F/YD0e/efupV3dneNbSIZiBnStEaUT+ft
No+0S9888SUekkADUupdXP8QZlkRamw59DW5T1LLhYZCBrDOVWRhHS+u3h4apyIN
wsh9+ThDJWBrN9bQ5zdmi/m7wOHMxW/KTO9llmZcBpSVZlBAKj4GtOUYzm+PY6V2
8rWFz80xSpkMpgwaUUbToh4BmMAJuH+CWJfpYIQcHIUyN2RUO7tK3OP7C8TsdXu/
oQH6kAn0SNW8IjSmBrlOXXt6URF4Ak+fPUWp05hRgtKFH9sgAuXFg+G19V4wVWlc
GOp0P8QV8x+R82CoQMvE9hvD6GpdOMxf4YwMRYmarbV/u/ncbUZ2ZILUGupMMepN
UzRPfBzAVZS4vvgp9Eq0U1RBRuSO9Nfpyhg6O5JnTJOCmYNXe6eH0sBZsn3SwMV0
AmFCBnGJhSD4heuFzZjJomp2CX9UPp/opR7Jdc/ZyxfyoGhshdW6lj4cIagVsdfy
T6uMTaYXCMuXRZVhQgrhCYna7UxdgFz2+b9pLQgeF5Ts4+Xq8u6tERDFpBn2Bs4W
Aum7eoeGp/9G+SfyYnPtiRobKpkvxj1D80z3bfWRts8vpT9atDJulKikmhBg8Xw/
DMdSXQSlI74a6T5FVJojKCBM6Z8p6ovhA0oVYwrhG0pSlwS6T0KX9SUGrhz+U8v4
oKVboLAqdd/EvawJ6yVSMtPL1OuRuMB1Gm4GQJjfCeCplqMVCf+ClX7KQ5cYfLtP
L8hlnh4r0T6TPyCQjp/knmGhcK+eh3CDndJL/xSzeMm7KpjJ/AlopviDqQcWH+QC
ECaZvyirMzQ7mrrwlF1FkXjXcwjsQExi37k210TLr5B6lRZ0ugy4aoxBM1T0MfvY
tZCahCF9NytdCqGm7lauxC+P8+ICfyBPtxK+sbViHDCKFww/wr0mWNdNbb3XMDnm
+VqMjRzg/0SrZQYEudndcGsCjZ/6LL6zN8VzEo7x0XFzB08jXNE6fpCvE5sOT6Y7
lIKj7DCSPB31TthFq+lsFgZI3AB24IQi4j27kIBwfrPMR8jhlYqDbK/Jifv48ukJ
pVC7rb7cnawUMVopxdB+Yum3436b1G/sHE+EMbGMiiu0O/EKgVsDObYrv+fa1nsA
CC/a4Sr3w6So3fIupIuikNcAC/d7R37dgOMNkb6Kgugihf2xyPDDZeddWcY1QqyY
Of4Mu64NOB5f5jR5zK7BDu8TL0e3nG23qVfggJ/M+iDGl8aovTGSx086kg1I37TN
AryulCQFqZ4eMrVodkJr6MpDfTJ1G0HVD94iVYUiaBfQT0JbJCkD3A0qoAD0zUhr
AMsyim4af2BTZQCggaX9uVPvcU5pB2I6qgOtT7jua/WBTkBlgvGGhsI2uiFECEo2
vHgLR8uD/Ldr5smaxDcI5/tj1PqQ0fIEw4i5ABTx6yqjE9CIY27tr7SGu+3MofnT
G/Sq91gaFOi+DbRJmolvmt5qwrZIUFyV6pGyy/9HfP0xsGauodIxAR08p5fi3Zo2
ZQ0qRImor0p8UgDnOlUuLYfEwW4TS3vw6psWHJLT+s98OsD2sT2eYInZ5a00+B8l
mUsPQrKtBMfHkDf+fk6XrItHAGIHYaiU6lfh6/ugoAGmfxAXjBrZnjrzIX/VzgsC
+CLwQjybwjLPoavH4bWtvKemEFZL95UVhjV1akE33iKP5+Kmf4T6Ev8pTDjw7jWG
`protect END_PROTECTED
