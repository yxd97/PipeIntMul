`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gApJwm3qQknrzNWC+h+hMjyHaGxF0hpRiv453OtIirZAhE/VO/bwRXvtLiOg+6wD
deTKOp6lCWirNPazOmpvxB0U4Y1z+6boVygVEvjj2NG1R7CMUuf7tCpxX8Bp3eaJ
e8e8AnEyWqYwcPPYfzhYkMJ6r19bwamrPBWXLWJ/wYt+suHKRG0j9/RVux9FP985
HR28dg7M9hnwiSsdkFxUAveiutCwxPdQOaHe+mo3MSNzkIxrXoVZpbMy539dgBko
`protect END_PROTECTED
