`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dq5jz2/0flhwTYhu2onM07eT5+JxPttjFmVUEMsZuWcSZVLkZtg+VZsYAZYcVZis
vh4CALrlSxi1gkXDVluT91PTaAMLkMMa+5zdXfqWOoCyHR3K/8hMcjlhTT4dGEpK
fbfgrQ314vX6XX9nN2ZKRf6I5EaN02ohXXfqPW5e4Sl/EYGlWkLJg+uLotX8R96d
X1Uo9Ubqg+g5zPCMhU6Kbx7QtGFiMch4qnj5HEQ9qF49h17WIHfyRpffyDiGOaKI
52HleE+/Wtxwl96Zx0NorBTx+zvGZBLFFNdSOIIq0V5ZrMV1m7M7nHlM4olMY2+/
R8L0Cuf+4cTRk4hZAaJO6F03sZAfTPYsRRMl/KQVQZnWU/sxwv68FXyJjGMOLA1G
gN+bjJ/w72i0FxBPAgyID9dJHgrDRXOaFVpdfPeXHePgR6L3B3r638NJcU0xWtyY
+MWXhy6APufQJcqOIZV4bIU7lSXoEX/wh1ZwEWnETZWOJQCTLr/WveAwedI6kwxS
Jb6nypfj+cVizq1M+EgWT+sZInr1hcWW4R4aOg2JHX40ZY/NeqZpAO/kCGsHZ5qA
3PAIixje566zbnqqupWYvBz6Yeh7UFTlfc1u4grcKmP8IFjsMUMBj3F/fqk1v5dY
qMl+gGIdeTBFvA5BtoK95dcCehZ17ay+ioa5KO0gtAakmWy/OHSALI41LnKqddpM
iuVdNZWLc9SvzufGmmrcUZbPL3Nqvjt5uCEGr2r1UtaO8s8+oW/q8XSE5+47r7Js
ASUUelcSYs3oOdhzI2cmzAeXatyWpZwDXrxRtcsPJoOoacskkGJiryrL6ZqbEEgV
Uf+sjXXqXa9QfqXfyfPoZZt99K/AKJiQi08tAE72oJTi86++tDVSMwY7/khCEum9
WuWuSi1OsefK4ULcuBESVH+vlIJCUIqnyDl8yOTgTnHylH3TFpWeTGTGhBK1di6S
5ozipSVqQJscG2SSzd9/uiIYh0H7JgHlODNJXE6Ae2m58lLAD5N1HlC8oIZTlgES
y+F6xflUu4ZxtfodLURUAW+iSaqd/mX2SYd+hhTxxCqZuy9S0qDVGbo63ggo39ad
fi5bR7kK7a+z8V6z/H4J7S+ltx5wudI2BC0NyZ7kuTith1BAjBs6/QDX8/NewxHb
2xSuAKLmd67v6fP7hXCaItTEIVL2p8F5n/CdG6shT70FLLilbfVXBN/wtZmLKRgb
dHXgj40nsdDm7fE7sfnwh0Z4k4uSIR0rE/LiB8dH+yqqHjWnvfh8JIGIikZQwGHt
/ZAvmYUANSlFR6tCq8y5uco+8qRCNJN8DM4Pd0yquxazgPqbKaocWJ2zAH4cSfbI
sW49gPMC/5IwcGr2XZFV+x1HB7oz3zAIUYRwbL7t1ImVuEcjMauPUhMcu85KepnK
4HeqB3NMm0wKa5xNg8iWjT78wnVpespeufAWohrAHhfLHjxb8g2bZOvnoVQRAQ84
NNqQBTP5FGOvMBXjHVlcdsqjNqxxAB18RRuKvniVPLiDtS/EG5ofQiurnTNO0QVA
st1TadSQAkN0K9n1mJn8EP7G/XlbZDx6vQd87irrPkBg8GVHdPXI2HpuGfCgOTzc
QHGkyxnURGl6D2EEFTM8sj5+WLHqYaEKm4SMiDlCtUcewS7xRiFx4c98SSXEdILY
4kDD83WBaNqsISe67aNy/K4jT2a4t2EI2qOO2E5RrYt/ZB9QzVymQys5LvPoEjnN
MyiXQuCyyF7lHOMyR5rxHL9RLf8pPmoC4bnw9k/DgnxQXDgxjRZRotG3Wk6ByWYz
wMva9UXLVZUrU4cLiydPfZ9RUYc8mTGAs/auOsVceXUPJr1tZqXgKq8iETvVMmaz
XNG7xwGUpgPDK7idrU//NsYm5kCD+o7aYuyLm37nCoRSiub3483o19SegExytTlK
+A8ZJwXbBooLjMciw0sB9Q==
`protect END_PROTECTED
