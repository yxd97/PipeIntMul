`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZC1MjJcyd7UsUT/yxYxFRglc8sF5snCGc4HVFMdeNnyuwO3vzpuqxteRF3qixBq0
BfjH6NPRMgkAnQ8LrKRwaNmAGRRP2jJpPQWgPm9hm6KiiFBWmhRNYX58yehX0035
MscaEg5sglnL5m2nbInqPg3t+hp+bntN9gPe4p5X8AR6Q/Pqd6Pr4+X96HXVE6ea
ww4eMQHE/42Tk4AnC94GXKLUX81uSTC/AKk1Lnqw0TWoiJ5NT0qZWV7s2Tx9SWvo
hErThnglgnTnl+3Twur5zQ3QCiX3ET30W0dumDXFG9SAdBUQh6GU6Cf1qZy3Lhlc
Rdcdy3XaNztxi1VHrzLfFgvxmrcDlNLcJ0hwOwjLzPPDSYccj1G61vv2/XIAW4Wh
HepNwiMhEM2eYB4ygU2DBAIlr+0bzo5pRtJIu3FpmIC7IgTMQ+CqrF0PCxs33J8o
`protect END_PROTECTED
