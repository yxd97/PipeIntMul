`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SsWN6mxNZN48T98VDL2FntdPId2Sy9siDYM0TvMpOwOXWnfwUQnymkIB1EZcb+UT
ea5lJbK44m0lWQyyHTsegfJG5fTNnK7OH2y87lvihOlrQcUzLyryhBJerlHExUQF
ooMZnsanQk7WXTv0EKpU7MV7dhL9SqUQbFaslkC+lK0n+jGD5kl8CLJXEP5Xq4Fb
UJozbVldHRu99gzylmeDCwNpG01DT/I6XX/0AufL6kl2QNmzPy6HrnSk9AwvG2Hh
CCiHmc/0yY/5gj+PtDcBLrg/P64vFVAAo/ZjogMLplw=
`protect END_PROTECTED
