`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kBKOibBDsbEGnMpHSXzwsI47cdI5ArLQaq6O+tS3O3wJ8DbdVnQkT2vnYCzzKlcY
GuGqTO0tMoAsrdDgacIlTohbhGDmTFltAqRPfOewVpZ+Ikia8pi18xBRi6PfAgdV
huw+DxF4S1KxRSnL3PXAMJgJykFV+Gx+ATftcLwG/BqZZB0XmTkVTrsu9cEonIkT
gQ9LI6/IKngA4SiEpjikfKyn76/E/lZRnkU0YVgKfAr+c3VGhaPWI5NoPQLVNIDZ
4e9t4PUatQ2lJlGCVH/rSUCenwAzAUAP076xiT45oCwD5xnKHzFnK/qg2ZE1oJTv
IJJT5kuUdViaciIEsQeZdL8c18Zg1M/YadnmC+JXVizO2F/yARNTCaBocY5WXOr0
GJsEZp3S1wWWNeXcPjZKQgmeNjwmYeO+W5lBiHgUmV0h3+FVSADQqLW48kjZHu4J
`protect END_PROTECTED
