`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iphR/Q4cCt80Y61cvA0glODUTCeZg4sVzkPhHa7S74NS8p8+8bn77kvS/IKg4ud6
PBtq/0qT+XW51U5BycPDyrwJ3uniVIw/DKifNRo6iNo2fVwPdQa2OcZatVQNeuIg
5MAugj7nj/RE9mOVBKIzFianz8/ElFRTN2FUpENzYqDt/paj68cWfI/JmOcvVxcu
ZYHpybpmdg29heoYtpb5xJl1Y4lFdhxC4iR1JVlctyyKFQTcvNTjz5/Tu4aZx0u3
xo5F9s77zy6Xy9NUmNdzN+w06P5xZpL0I2/aZgrktJ0Vx5W6XeiKeyoxcbUbgTkO
l6C0vS7A/trupYsm1nZwbglCU0y3sIsWCXIkAZCr4KmgmdMino9nTMeYQ+HchM9v
MXkExyFgZNCW9ijn+tuGf30yzkvMRWbqBqlf+DKLHrLWdkzVC2tiMigvKmBx1jom
3xjnVVqC+l6kaTjQ76m8Xq9PqD6Wqf3TjDPDhjx3TEY=
`protect END_PROTECTED
