`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRM77UBqJvs82xh3cL9uh7j7U1jIc2dtKaSQOubfOLGEcx1l8Rh3mdLW70AyDESC
dpvAqLM36pmEEbdvC24Vf6M6xuiCkbl90rqQ6lZD6KnPYQ5+d7R+nr5vEXQBLoDM
SLr8AWOiLED7okrLk94w6d9B/mgpw0ARZ2sV0QBoHdgDRlygFtnkf2/B+diXVNG+
YTFj6cr2dkqozmtKphW14N++KF9i2LT+tDG78lfJDvkLS0Tuar18GzlIsQL5jAFy
mpOVgJKzNOPYpQAdEyKDOR+ijdf991KW7WMOIoNcbdwjZRrneA4MnA70Q1mY1bCT
XTj3H5IwpGZ15XUPdiKe8JNzYUCA2xsSFbUYdPmG5n9lSWzKxtimTIKxy5ZqulpN
ed3lPFIVfDnFl96sh8XBLr/i7U5wPTXWFPTn3cd1LPU=
`protect END_PROTECTED
