`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vr/sXpVyVISCQBhExRKxewNQZPKLfTJUVx2x/Irl23trSaYlvdlRL0V4gcW7W5bh
xefSv9IdcYMr5Q7ekt0Uo02xpTY1R7RyNrPfnMz1OZCGbXFhlJ5rLAvBDwm5XfLf
jtjhCAQNZ3j+cKVRoi/iNOAmlgr51sltkUUjS0/hMEAUmVbQ5naj415lVWLRPWDt
n4DR9h0HzhaFwf9ewpOJ4sMS7tLI2A5mx6YP7kj/p+0WJYEyJtz/m2fL92oX0QwX
BDElAReWTjs9o/z143LQpJbIGfPNadavfaA5DZMzlC3JLaP524H0e0rW3WVXk+r2
yB9VC0H72bXqKO3lzz9Ks8hfNwBm5Lqjd9QjCRs/H7HlSYeshg8n6/8G9fe/wrzc
Kd3mTiCGFA/0JHenh45/RjaW3g1lg7ICu6DLGxlWrCG1Z7Kgifl7lro1JX63IJu8
130EcFivUtkANoWCNnNX8VaL6N4sjUa9yrgvgJpbs3Yrj52yBAhwE3/CvUNmszd3
aOgAKoeUq0u4do8mUEo0Z2ObskxAx2tVMocMGXQYERIQB4dFN4h0CSbCAsIXdWlS
2u3h1gVgl/UyqLaxqThDchp9eRZnLKXGQywWYg44xX6H+87rlmD47y9IeQHG8X3D
Lr6JxqfN19EflZYkP2bRjdTd3dlvlSqupk0We/15xjE8ikYgcxAiWmNipvMAgfB1
kV7W4bhQDwlq7fqwVzGHMbeG2lEKAj0ikkExEJBezBZLqzWOVm/QT8eqLUs3ooQm
CfdhMEIxPUHyFJOaItYodA==
`protect END_PROTECTED
