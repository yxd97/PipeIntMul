`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BHJ+jJxVlM0NBeJz26119EhEwMDiHKyk4nlijrXH1imP4i0Nk8/dxYrNWETMuuy
LynN97jyA3J4YK6hLQaGaiF+8dCzn6RKgyRG+PiOp4uB++glEKR9fMjNhC3MEHZK
sq6gkTO2yqkK89rxPgFQa7oQKOhIqf9K0vhWAFwcaKnuZ1W41XCsiy1VzhJKh8Gq
+XwvfbsTZda14ZjWkV9QFGkGEY/rXBG4NaOLpeDpv6HHmkoe0cSLK2mJFFMfdzpS
eyGeCcKvRiWATgY4bDHstY1nsBlq17T48S/xXqcs0TIIvBNsZandgCOZPcxduOet
OL1I6S7l48mldURv9YIxvL7niO4fqN4TcdUpBh84HK7P8xzbqr8ahnHo9+Fik+Mi
4s3Tx26oJz0/LDZbrXOKnVm5edemtJL63GRhjtgIjdT7HtLxDw8CpquBSjpMP+Bd
pvGVJh7Ticzz/SkNhr8jMXD/X6qodGxTfJOQh5A+iZNk/9FwQgH2cyH+AvtYVYX+
Onp9OC3R+wGs/el5r7TkN2GJX5b+miAO7tqLid0djObZ296urFw1BNLST4CMAWWP
/WddqAVBlZKu9HlP1xz9pYCc4nzxDK8sU8IHgrPcM2hdD4HuXjMtfjuRizEn61HU
HFdz+GPjWJUolMH0uSxWVYU00UhuQ9UhmyX/Z9rK1BiST3CD0h4YD5Kd98+SYzwr
rev/66uRTszvgqLgMi8wXZ1Vs1G0CbR3OBbtJ0waQbDhctuqE825210tZvoaHllM
F1DFyb8/kaUZkhsUfH6puYr4YL1TGiN+1NR0C2+7NJWUtSPCIrwUS50JdSDXIBH+
R3RlCZfad6u41FiglNOM76imcskylYUKRymL4IJ6ozOGZyo+bV4a9TgbSzOmKOSi
NwDpMy8Grn5htAXQOqgUux2HRqTNaDUr9FxCeM7sWCsViOegGN+cLzdoyLhdTGmu
yZofXR/gHcdwSR20y8NqoofPVxEXzX5wp8/6c7ikTO0jsDXzBpb0ZD8cYCyxu3px
d6EijLHdu9yvJdnSB5hbYez49fKgwjjMUCtjh3CHApGo80nIIel3B4XoCmgncpTr
x1ZLnhQhzALUu5iSNPKKNlVoG8sneGzru4xWpOQthJCizePGgCt4/+VwtnWsHhjy
AmNBXzma7DU3geN1o+eJB0Ed5GXjCNIPnyLX5djUcPhC9Q5g8b1YSgcSZfV3WBdT
susjiuHBcD/VgvkUmjBQYSV5WyWfNR2OJaWxSw7OEk3Km4OCKwlXw6cPjzYxHnu9
0+YTsbRi6/mujfcaY/HJBnjpYDt4EUe3H4kEJrPchYPNpzd8RI4hEG7hukAc2sx9
l80ejy+uNut06T8bkMXKbMTuGlNypTLDbK7uX/Mgc9LKS1XwUOelXfXJmWZQnxCe
cxjRYG8B5FjJaffQHnq2Ldi00VEA8BM/3lWVlf6BXi4L46iiOZZtW2AnUlP1yzrB
l7aj3QB72SM8dyaFxFo59ZpOWQhK+0isHAciKI3Sgrna30SEeWo3z9hI1BNINtBl
gsG7Biwc7/BrhX0UkWwt9BSTuGgAmdbV/WggxIhtNHvXqWEY8yj4nVXLVW4QIBe+
6Mcy64mL52OFvghG0PbGQIzmRxZ3+ygsu5FP//Q1hZTf/LnUSJZxCltyEe5g4N/p
azs4PHfwqbNeVyYthsgGsl/b6CC2RWADdUePbNQBG9WUEs5bdt0DQdyBvHLg2u7F
g69skw1g993yWcKNiDlkdvZcdsi6ssNZ1oOF1eQc4+ejEUWfM7oLoiCapDYRpowS
sMuZQQELKEEtmOxA3GT/jxg4W+xNmQqrJt/G4u+SXhtWC1k/n+M+RlqdadytVDK8
EXl+uBuiOSJRlNmSDRX+OjBV+B+/RHcuWmuqXExI4ay1mSTaBIdT+rJP8+Kg63Av
VT5tNlvXvKXMB0l2FpTmaaH8OMgRngMRSEr6mEG/QAtWVLHPGbn8OveYOFOhSav4
LWQpnHXX9vHfkYB7dsSqB4IY36gqMGvLzdkAMIb04EORm/yNQLWe1wZ2Iymxu9EG
jp5oVx9W3B+haL9imab8WB2/YcBYJoC2CtAkbG4EluqmwZvvJ3EqZapRrSEJQXOK
MfN34S7aPL5qN2LMIorJDXNfpshkog4SITSq3X052i+uK0v7f0m4e6277cr/w9VC
laz/7oFI/t9nrWy8Gw2JQNBrLnw3xNi2c0SBPhm/cuTSBpgiC/SIj/F5esE6DuAZ
riHixgQB+RPjESF2mgDTOv/x7lhhLpSFkrasayV0JX99AygQzBGFvkPJLV8+rgsU
nre3ZJSruAbNEDZ2PnL0cw/M7RViJyTohC7CHLoLZuXi6cHOKgXqYiQGFjW5Fhfh
Zg1FJSePvMRTc9RbZpF372kHVwfnex6aY1q0xHaKNeuJhK7wXHtFhN6lUDH+TqEc
2QNqtba4h5mLZGRHmyBt4ATpWLWlSKVyVT5jj0KDQZj24KP1g60v+MoqMK8N9dcJ
idtBedX2zjyr/6RluowYY44JGjMz1CePvC8KNSqeaaExwYjq2pffIa4W0jFakMYJ
qFh0Wp4xZuHZF5fv450DH+I2gB8gw9mCJauFsvLayhS0G7NOstYdKD2pb6KSOF6m
aBdzuaTCqVdx2Qu9s5ETBQ==
`protect END_PROTECTED
