`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSwouRxxgUsJvK34xTZ4e/PcjnFtBsB6zwpAUyyu5E/+HHxxohtNYe+T4sB8VGYU
ZHQut4UWoxEs8VAn4k0lHVkYfKiv/oXLQ1zhJ+wsq/SD9RnPfG8BJLs7LPOPhB1z
8D4Q7K8P/xTvGATdULednrTZtd87l3HUZjFPs5mJEEh/sfNv/N9AbQGqOGnhT4YN
SLUDaITGvhX1s6bHo/Ois/gQXZs0KeDgll7+Gm/GVGWhbKJOjsb2fkMWbG1GwDMR
Jxhn+On5TFsA4BNq7F7l9XuLUcL8qEl5kmbLwwbHe72u+mT5xmL6L/lekTLaJWiF
`protect END_PROTECTED
