`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tT1BsRuigbxhuBP07aQdxV+PwswfiZ3QSCB2OYTCQeEB/tT1MedC4byf0Gayt6Fv
KQ45vB+aPTLEVB7rfoT6/Mnbk+uomxGo0T5d1Kj+ztXzcyrUAFVMTSIhpsgBbsBj
R73UayT8eDugTZpXxrHtzKQsz1YdsKcAkWmrDJDexRFFsQFYrj8ulDGZK8vQ1LJc
oFTHn4PMwBOoWdYJAz2LYKzYx1Xg1ySjkwjqMU5rmYFXMUYd2RTNd9UIbtFFhLTr
PY/Fc77L3t3ETQ01gy2etyr5VBp3dn5unaERAZmM2kM8Kp3Mu79UlElUFWPMhqiL
vuEdVJQNdsrNK27OmyJVPGO9gt4v+UfB79/5p45tXQjah1Ui2CwPcZUDZe+hFtTm
NMg3ZJKAjI0g/BX5CvtaKrKXDiFl9/0NrUZqYt74an/u7/y5XX4U0gngONnLO7Y6
/nGxYJ2CaCdG2IhiBHBS1JTyCzQFEQol7FYh0b2KOzDsb4VNyVgWQC2UpX7uCLei
+kRpwA6/jUe1SDaP3UhA1G50yL6pFfHphdVUqiHuBbmnUdGU5cCn5r3kMHub73M4
2TsaLm3tUF7piaf2unPCWum33FGDAJ9vJtZtHCe3SHgwEZLjMGPslJ37/to+ALXT
kZeLyCSU4MNniksA2TC8BNMDdEu/coD+KJPJmvW4aK4j37PnT0DFGK3HDLJWukaB
7UAzwPF5u7tKQHKdK4Xq//yJe8tdmi9W/JL5F8nkKuSgam2JqsmDn8hAAImYszBi
5Di14oA4Dih07lIrJAfD2lV0iyvuv/YvzLSKnKazdQDj8cCyf+3JAgaYT5Z3iwFC
0dvsuTfq//FGuwE9ki+MvTnaGeh6Qie526+3oTagA6+6RUiMl/CdeohKt9chRRLU
6GhmXkGb0d8gBAe/58bJDQFT/LAnXJrjPS5md6YQnzVoVFdrJ+9POukdnFkDIhF/
oehbmldkN9UNrMsp+7JnBzHP+1crZl8keq+kGOVh7RVdGtf6SeAJG+ZKTcCnUCgL
fDwYcaFzR/vwDsV5Wsexfi8mkkrk71vjkYqQ2ZPk9pLtNkiMCDoRCzFowPlmA+ba
1Ve9a6TdXzmtXeh9u4PEF4xZx0C3d4cGGLIkzezRajiI7ORmn3ToFpgFjvW0Mt3b
EanivVyD6Q9hgEyDmxgl68Pqs2gvksn1Pc3x95UN1+OnhSGR1gc0o4/YBDBzbaDf
ic+qFlQzubgjYAjopEffnwVsw4k4MNH4PzjZEugAcd5+sfHYR7tnGB+wcOpaoiN7
w1gETMnzjL7szfGuEohjQ2xfNuP9xzY/hmk88NMndnfw8+8vp/DAI9qKi+qn8Mlx
hallrho5+UPBfd68iCFRmZu+nh7OH2iKrtVH9FUIVZWFO4/+SN37ZQLW7sEqyNzE
3P4zoJh/0IsnmWD5uPMbpA2IJyR5lPH8kLiUMmvAJ4HonhhuEgJUFsvy1S3oJF2/
qhLkjYPBBI0dE/80pmTlfvHq4XP4yfoh/sDEqkYKZBxUB8miP2NELaclNvqVsa3X
/Mv1K8RH98Y1e2377NsTGE/pttZSPfyRn3tXqZeF10iMJ+1S3vWHfpZNJkb+QfVy
skkuK//nnA62Y2DuFYSxdBjpVdzh2yH8c5VVPFmtTSJ4fQYrlNhvZNGr3sj/EHoE
/0T765YRd8zzhurYnnvprKABPwEJwWduP2YNrhf849Y3z/HM5P3+mIgCIb4/qgec
2myefl8IOb5229n08XEhsJYc9iDulw7x21Yys0s2cEnCHvR5QEldLiR2FlPqranc
2Ct/zPigkqwJKouLoAdSTHWeqM8KL7OvAbe6A0ClkI3+G/bJOQcwd2wOjtArXB7c
0CIVQt28THf5jWsIktVoidEAPYRMjQylVR/nH0doLE5c9pF58uYpwrvGOkQHb1TZ
P/jjnfwnkZwc3HzMtgQ0Y2I2FamGTTsZRM0DKawTazE+MyF/mbzJ3smestsVOENy
yThVuS8BuKiGePWr1C6YwKqdGtg+Redy6B8X5N8XhEEzF81uCnQLrtHiXif37P2k
cJlZ+YRvM1fkdJnbGzKUz7eJZR60FDd6wVwK4UT3bbQ/3fAusVcF+Zc6HqcwOUV9
DnTxDBow+JrQTYJp97zreYh14kJlQ3UKETW2K3uN6jJ9UykpkWgYWVWVW6rtQO6y
kllTgTYzyrjdbBcdAfdJ9cGsjUH6gjz35hsLsvxSVx2+PyIR+w9nqPvOwDsBnReb
6umsVs38zhv2l1zmfr2nfR/2vjydC9uluoJb2gG45dxt4jw87++XfqqXoBe5rdv7
iEGxlB6BSIbDO10Etq7ozY2/4rSbL3jlsQKB+M4zElumiJWTIa+1yoqRqtgobA4d
EAUyEivkEZjRuRJR4+GdI+mo9xV9AixtzF+uJYH81AiRoVNYN0Fzk9stcx9Mgj6E
bfNDa8lWeuZutWTqOjFZZ3U5GfUyTn7n37+s7w/C/FGDhgQxqIIup8OSPQg4VWMl
2V8LRQhn79gLs3tcWaqO39BlPB8NEQ9I5N4Zd7UEAEaeP3Ghcz3UMF4MAftRMTyo
kqQXTqgEV75IVq8vW70wYHwKMY+Cm9opaKKGQcMuQznRqscAm903v6a1kQtl3iDK
lJ7CoZs/WAS2H6KqfWplriX29P+CrnVn5VfVzuLRL5cqPUkec+fFOKE0rIv2Gygx
vOu+YifNPlzxkcOQ7Y1hEm7FlpYLJOyJOGSyXoqb9QORsp9bGchtN2QM3yNG0fxa
tzDpOblNXSosQRpeIRb1lhOv+F2ZxzxpgYmb3cJo43GhfLUYQa/+HsF0UlhnJ8xg
cqcllmLpZhPEvSQqvGDlmgT3ostPf1KNhNKdEJfs+PEtveGoC46tYeGUlmicX8NU
JFX+0gwI2U0Bg6hoxXmZOz3737E1EFLH/OOQFZgZlVeb1JEObmzFhUOsNbxaPzYH
RbyAaU6Dt1sR23CbGYC6IjLC0VPz/NMjVgQ02nRJ6zuyveQ24ecBKwgyW8S5s+CN
`protect END_PROTECTED
