`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oOh3M3G8xW7mukRCdbnwOg8zVeda3o8kjYVa3drfkux3MbzhlD89GL2x3OkRh+xR
aSbBvFCv0vq6e7UbTpjHEktmXqr9zflqq9HYZoNIPXom6Ny2RgHGjAjnJ0Wtec9T
KEaOIEl0YnoMf3cuPlmULUI0xC9uwPusg1xy2evHf1Of3OsLb/yam1WhQ1av48oa
AtKDp6vOzNpuuEt+4uyNhwR/a0CwuyNSey+9mMor/fHoiEhvbpO1VZgRLrTX0Wjz
4uDYago4LnQHFKoYIHYWI8FbjhM6YxYru7pD4P1LpciSzJ0XeRqYVuXBu5dRsGrG
ey70+tVmBSdMnP30rjNYMelRfjyIpkUciVhL5/ZHQP/uZe/7VOyskjhj1cSJj8vx
SbHlqMSHalDequ8Dno0JgmXkKQpFFBw/EKhq0U5TadpWC1oZc5O7ElNCjXcObXo5
V8hF4vOYPP7vaous0S8r6Q==
`protect END_PROTECTED
