`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HX2cs50DdgrQad6voESzO1HxTYpbePLnv5KJl2RGB5mCxDi57PwAW4sVaQ1XZShw
XIh+cilUtX/qtk/kz3B0PoJI+sgDpr60ippNiE5pm7s/NlCjCK5g7YkAF38W6gyc
EbdI1ZmMGWvbZPmK3BT5cYYabFhjC3s5IFMiq4pMfO/8pt496Knr1PDq+I7O90jo
NmwczRNumFK90hxM+dHL6Y/jtCUpXfKOQ0HqhkbH9S1om/7ovVicIDdd/AkCmN3T
qs/XWksIJUsGOZYeDN1FMfAg85Omu/7u0yWO0cZ6jrY=
`protect END_PROTECTED
