`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
It1KERzUnGydWye37ZRMM8fUO9YK5GI9NgIVHEKVHzTjpQhWqhYvED7a+26qkx2H
1ap8Cx/9I+BQwM7HHHeh7nm5XRdRylqzkOaAI76TAH2KdKZRNZDxWQM1SW+pM39d
3qPxgpGC7OoJ4pVoI4caSEm41HZxzzG6Z8KUGMeOi0C1MPaRXcJn7i+xksHCiuOa
uQVcQ/ou+J+eMuaH8+HpBiPb5/yEd+iqNHEd8Q/U7T4QdfBqx2+g8jpwbx6qCU1A
LRFpmbi0r19eNNTEAF4a9PVjhyKDY8Rtd6AbO0NFQLm9QO0l8FrjU1IKwvwgLDuQ
`protect END_PROTECTED
