`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oUWopF5k/dg/vZVjZZxG1y/6WUhCsRfPCBveV0K8ZbzJ9dIO3ENZCk5mmpdvxLLH
5z4TpNLPPBgJkrjEg9tYk9AWiDW6Cx4JTSk9E0PtNtJUcbpjm+qOSy5Q/3oNTx3/
FlSFPV+V3chf9Hb3ZpfEpFFi/e0L9poqeuMPBcmSE+D3LtL5Gh0/XRZGEWkWaR6q
gXAhqA8LvQI7iasHR7JeeZXBBbMyBieSCYqcrmLjNACEX55C4Suxjd0TOR6NywdA
1qR8ChUhIx1KqF3jVXDgajjXO4XA2W7IplqmdZElDNFA/DGb7B3qglJWyUbwW5VI
`protect END_PROTECTED
