`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PBv3dgv0ushPuNIEe+wUgw7ILYOM2SDpQteGXbdW9qJM3IZnvtWWEIGHVc/aao5J
OJjJpww9vP7Sco9kaRWtKEix/r0mlsV72zcgzh21NtmmTJbcws/qitQPmYyhFQp5
43c8CScQ0Lrrd0/fxJ1bV3Cbd2oYTXD8eNE0VPNZPfHg0dM2iGDRTH/e16aJWLZ5
aBnISjtCMezG2PrOted4KK8o8WNZUkQ6XYxQqJACa3mCJtBWkIrP0oyin8LfMvNx
My3wMoKFgqwA6qyaJ8C9HpeMI8MCoWjYteE0MF6u0UyAc59zSlQu88bo/CpDXsgP
tdQq8RRzJMctvVBvk9rP6TriS9lx+7+6I2KNyEjPrbYEkQkxXYi42AKrQTXBsr8m
dPAEwro4wVvgX0Hg10aKuQ9edTbedQuegtsseyavL3btJFoeRreiB2l6uLif2p4f
kdFnp5QLaZzRiZ7CxE8jCsqthvsCD1dVDSCF3ihPnvZ8UuFFF7Y7n/ycvSrXd/N4
oNmCV0kH8nXWxlSxT1GxlT60mYGYtkuae1ac1T/GSgz6pNhQHis5qzzOvZ8ojTQG
SndmfkxlRyBHtUZnC7mnSLfF108UKx2roXMYmfgvyhgwwo/nwuvm6BXcDsJwupP4
3j05DX0AGICwWeoDIMj8DOczOlspjKHtKumk0p4zAvUAqcYcYSE2bqS5RgN87KIi
F7AUnFAd01Obj2XoYyC6nJYEPWm1wmdYsvCdThu1YiFWuT+ceeOtMD28IveHTpfy
G6tGoCj9m3JewJRqPVAvlIbJu4jl3pI1FeYPXygq4ec=
`protect END_PROTECTED
