`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TyOG+C2NvtCjD9CA1DXKXwQyheg00HEFLt0aS0Cf04BjCn9ToNU48I06N1kq1BHS
djamy8ptIdqa1fSa6on/0cDDavjEw0m40zvlD4bQYgLETTTxfk9+S0cdqVf6BH5q
Gex1/rrHBA1Eu7pOPFJU/kBWgKkwVgTz41eUDdVigBdKlj28UeqZYlKZtneqaxQM
UxaKrp+SMsUGUhgu2RCQN7a7D+kTzxcjtC9AZB/VQEegil85B3f1nV1TGk4GzYpi
M2xrYVr1Y0CRUhEGExQVW9yr1yKOfroqC+t/qNmeMJqtZEqDNjrI6fwxkUQD0Bbz
sv8UqudCzVgcKgXQdA/8ho30VoU+L2jH2sI59ESzJJtuPoFOZamQQ69boZCTpU0C
CcXzZeloYMcbblyFC0Au+jDefg/Mbim06gcCJv/7TP5cZs+1s4nCZeT59Y39r+Tf
B6JAzb+OXMpxV6RJssMVdC1tT5SlW7R6LTRfxJo0a00WO6PK1qdYlsu1Ru927ODV
NpOcjnyRuT40RjmdaPmWW2dME7hgjXWVYTbwBTkogJoBZR8bHOx20Or61ADdfIHF
QTGNwnjiZ5ESGsav/UVRuiniWg4T+Qy8tV184PgJZpsVA0kTLVzOgGpUNh9DU1L3
QlJHVauQGJ6rkxTxoqOQJiJlQ08QwJAti1g+z6O6BF8u9wvbI8QSxY3x2NLeNVX8
3daIYYVXT+6QCkCwP0UXyQKhkAG0Qm1x2S1nlx1MfuF9XYPPybTJjUI13m6VPdZX
aQS8uiMGHuVxtdnFWDqUJ1Bvqn5aa7nijt3duj29sEWg6CLauNIyqQbaM6hTcFzH
ZHStPDDb6ItzgO6KYJ8Pm9ArK0W5XaQ53R3C2hVsP9NJyHVoyTzbNbGgyYduw3p6
xkTvkYnpEbO5GltMasSI7w==
`protect END_PROTECTED
