`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jp/G11BzPRn6yLBl8YdJUHuwkh1oONVsSYUf4PUz0kRxXYC12Nu+dyLTWec6/OPB
EYUfsvHR3zzLXj/mpFvC4q2E3gEaS3Nf4SmctIu7XreL6ryv27Vyh/1r635INqJV
NTh5WTknb6jeDLPaHA2GZxxs4fd6UO0fTNklfUQPuHOAs1zXPRxZ3v1yZduRq3ie
k3OxptmASQSyeI8KobZBqc2e+YAr32riqVAPKKFqcvVcKHCGoMfhPu3oZxDzXEGv
zsTex5IJCI6OCbancAz5NF106WSu5gn/F1O/FSogi9nUzBDb8lDOrzXQOGYRNuBM
yO4txejU8WwukB3n9yHlX+MDZYg1BNG6/aIweaJXxs0BfNlCqLzk+dJ3KTstDGcg
fgAXRwGQhNVNJ6xz75ME4Jl2Y7wOxuulRNzYZFr3FY09+VeHt6WVJ4j/hwXGtGYr
d4H5YVUYVcU2aMoQW2JSGErFK9bYwOn+RYBG7qmY9j+IxF0hHwm9prMsJ1WJFWEd
QBQBkumZ4hbNP7vuzS+UtgBrfLtAkeWYlJj17Ikp8EyaFcaTr0saYE7spLxbHuGZ
haa/8lNZ43yiR80xeVGKiA45o1NMSHnp33MrhYqgJ85w4+teBW0adVOXnIGQoIwD
aa8MyJfImWb8dsAJLKEijT+3MqCEAX76wuD74pyTqR6DGY1cW6hoglwt7ycbpfJb
fvL9HfP1OC3PJBuwyZop7Q==
`protect END_PROTECTED
