`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4z5+RbYHZZHMgPfa3kbvv8a7Lc11T8BNJuGhZ7CxtZk1kuyGAj96iMAuEONhB29L
tqRUHB4H2JJf2wRkPlhG28ftmQbm4xVA4u9ylKK3broDlK2obmlgGRQeE4FOffqe
ChTDWYEgPcKCObJ4AOMj6ywJCMyoZ37P/Mw486Df0YMTTro2ebVRzy353I52Senr
2zxFkZnA95k+9P1rwib5L5jyu12OygpAtcRWkPuz2NSMcOgCNwdG59i1qXbKsgc6
mWRohes7DHBoq5f+/EsPvRuCqbNYAtpVeyk+4IvLi95mXCjOX76dJnCBhFgZs8IM
nliQRuaCXyVGoiumFWSlT3OebF4Q3gx1JuYkJ1g+50qdTtGpoubYVs22fUzsYWjQ
raiR1TMA8jKgz9i3uuS4BPwfJHs+iN+pvKYh0BArhYrBnXxT1sHjHNoEklERufSx
RoS77M9WnMmG3MRT/OwGm+zKXgVCmE2LYks0WJdCO4IvSCgvxW/Lm5i5SovOvbA1
jd0/VvkLUrxBB5zY5uhUCMc05YM4vdgcYuYWD9OvWu3J7dNcreyuV8wRTvQR8Tv/
fy9LBWD6YBEhs4DaW3GZl2ASX3G8/28lzsggSp+A6BcEv6eXolK3f4OuC+3gehT/
p8jjd/9Gp8z4F/YFq2JmRIvwqPdmpoTW0pWjhiKDU8bowRY3swBaVwlbBm2fk+0G
gt8Kz9Bl0iHtl/1tTPk2Rbtfn8Zw9pCUiB7rt2f0WNNTqjxRr74lR1u3df4xMr1I
AAdfYFSjNN8g3XfDu+ktAjUqz4OGgEpl621qPNaRTmUrM4PWOX+NLndxab3lGqJr
1naSNdk7rK+BVw0meVrg29UDWeM0DQJFhlOAQkUweZEcBMOD27LfxvbRLaT4PbWk
8tVaU8f5S9agnOfmOD12f4mrjy1o3gaVO4mlb2UwJPanYqlC1qnKB7XXOqH8UBWY
uA8ZM7M9y/u8tq7ZBNIPh2COuAIUvwNobyYZuvMgmuCrbwvBKHqtGdIN7Mp3oi2C
GHouNYQqZ7UDa03IRYKBL0ipvdDHfEgzBpXA+j5QdVMMRHnmJS8zYGZiBRgNv/Qi
Aw8mOtqFeUh7A9hpq4qeKkDP3GcYnXRssPtZtHxqaiFkpnH3knrGUAOc7VUx2tNi
Z+MtuGj5Mnj0VoNwr5NZmzawBSjw+HN0RfbgcLvA5p2q3ybALoW5CZLhTD8Jkrbl
oCJg3wbXm2gBbebir8BuMZwPBX+m6SXL0ja68tllP2Q5+baSBZd/ELYkjARJhK7D
jTiDkUHFwzrQpTyvqFP9Kq6HYGX3uIbi3gHfkgqSCDlM9WV8ZvMeYIy8+ZuqXZSQ
cU1i7odlceLLXdYl4sOmmN6HtM933fTr92cbjx+zzOqsu+4koikQ0DQlmNr62qLy
e7o/ETo6sOedZhHEn31L13vgi12r4ZKd9f0ssZn5G9ackDaQDj6GLhEu0Z2cdHUP
5jT7f+NGZICOj7JxiBFFt1Rof6hKDegvXHYHv1rrTJ2cU4uLB54EmUCvmLnmt2BU
nAFZEXYNehDY7A1K86s7jWfRd2PUKLptFL2kqZJIy+1f2B/Y5ggTBE8Ef02/XTwa
7apBSL3TPHkdTLP/XSj23DoU2clZK3YZxcX3SBs7jzhXJf8m5/xk89xn6JchdD0y
sOexr+/ANTWps9ZCH9/0zmOoMPFRZAMUfY2Lea6NbWgZAkvnmQfK4zENgLMY+9PI
7sSURAmIwmJHvzJVqGlIMP0g1YVJtsdZaEjvS+2kphPIwWyGdFasiM3cip69ISI/
6Su+lrffX+4tRr+v4t0F0cjhgKGqC7GvMjY8J/LWXGNSRcRYgARTatjFkf/E1KFW
hFkHdNSdhC++DTUPCf0ChFuASIIHfs66w93gLniPEr0bqkK0+lFfH2v6zvI/g59w
07uv6CaXwCHY1eioECtIZtoBiYLcvLrG7LiSeYkwrYzaAS2EmvwQdvUKBUhaOLwB
FyThDRLzKlcBD2WEr3uEvwXpT5T2bmkyXywiLVmVcYIjl5flbX0t3ZCUMWF6oTf3
tK6W0FR/Gl6dUrLJsUQUE6iDnUHJlYh9tZF42GVzwYRuTjsK5t/iqP44zK8YtzLz
mbcxgFPsfnJDI5bfNYFcWe8/mp+SpjBD/hTTKeHEvfelbqMt3C5psVg1HizR/wLm
zpj76Yj8jpPtgUWYqFP9gbvrU8bHZakjnJmfAS3zCvOpV6sp79vN5dTUIHfnHqVg
MDHlMbG0tDeYRnxD5QlxcGchuGy1hsK27MN4yGdKQ4CsHRfR0ow9NzSIGlfnZTQN
BiLbTqsu1uy8Ipz80JLVD8PUCZk2Avd3R+u+aKJAU1etXN5/nLpXNVzCAeIkHkSd
FPyEhutWUF/2i5m44qfSCg6Se+DgKFECwoX27bm3MzaRJNkL8roAgYPVldYGqgpR
Nq2BSKP1qztw+YAR1kcEmHXx5EQOajhjeiLnvr78RBiGPehQQNsMgTKcy+pkboWE
+Kb1KNwm8RArsZCjwYMl9fCjkvhfWfngadIzbpWKTKTLcWHET5CV3hqXRHOSO7JJ
hzG+igBi4mk61V1iE18QeoFMKkBKfHRXpetVQK9Wxgrr+0fDqtCn14//bKVVmZDK
r+Iirf+DZxa/qbSbwpEKH4LFCRue2UTHhmwtuzdSxFM=
`protect END_PROTECTED
