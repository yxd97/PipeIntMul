`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FcIjkKKpmQBFSPYEVltYzbqsNQZoNov9Iu1mIx0WViWekgDgPl0FthPV0/Jj3BWA
9vshyQDcyL0349CVSCitox2uTOB8ZqWQeg2jLDDEPP82ewL8qQfUsWdCW511IV4m
L5N+ewDg+YWCoHWK61Go+i1fAe87Okcl/dBaMZdK+MnYmKP35cU6Nr7LvP3rY7Ny
iFmUhXO3Lnv0CsOVOtWLTRxiI/pmLrrg9rKnII5QV1YtV2ezY1mIDLwHAWFfggBZ
EyzxPstuhoUW9XH/k6Oh/yKxlmKKJGr0SU8EQaCj9oW92pKN8RY0QBPyPR9LFqG6
2gL3ZHSAP/TD7fXyGTQ1vpjRGF6t1H9BzceApvvP4zBStJpBSUtgXz4Tnb3c+5MU
Plw0wH9G1KbxSlWhUnXEqBnZsMgWWcdcMzjIm1vIyXk=
`protect END_PROTECTED
