`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkzc7oj5vBRk3mN+YgRCX6qb6NLu4Nn104wfrmk0KGUtvDGR+LN6lFwPQWMxS6Gu
2qatTkd/2uolKItwoLP0XeYIM9T31xCyCaT9fYZFcXzMr6jPXufLVvKM7r/x/m8X
On4S/v6Ms5u5p0o4UcfdzzQK3axWKwIHE3fYftNJmu6awvS2Prj9UZwk2y0tzDWs
gxPx406gO2cLjom3HDYRKsfx3D9cW9W5DL5VSvLLWRQ2vi4VArrmyWycSMrppmEy
wgl13Dc/MJbAyBFYI44mDsS7bOxSl834diLoPCnMjhz0vFSfQFAlpM8Fq/xz3DAi
WTV26np28NhTLeK8DdRSVKstTRnTAtSR5ErBn9zO75sWD0O5Zdh4+k2Crf2BrOYC
qQdDbtxzNijAmNj1VO/lVuO4ND08ASTopUkPbCQ1ZRTW0J6WF2qVswuzjCCrn+Pf
cyDKjH8ZgZScKcqCx95EYsgtZIqLX75rE18gW1/QVKuwkvE3a35EzKOiMtvvOEXA
596oxvArMS+paxjpZ/Tnonj0oMI6n/RloTilInomN8T5Qz1xXc3lLM8vMtehV/Fm
GsywkN6iA6/RTLbyNW8As4P5qGN9RSwkL1gY3/5CMUSqIBNt5ZD7GyJD/QgWyeLv
1AgXWke+pINIsryFv+dMfATuLmUErnbqi1uXEttGn6j3rPGx/Do+I/tPeOo9cEMe
`protect END_PROTECTED
