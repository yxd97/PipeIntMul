`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vkWxMTjq128IDoNDkosbzG24rD9gjBXF8HqtDQ/seGkYpgzdVnOrSozacNQTXGp
M8ngWQ1UNRBE9JLI+IBKJIUNM+3xO/7+K9ngy75pq5z812uVh1CfgCpZEWh/8fNG
0lRmc/8f7Hr+psaDViOIDe5ix7AlwK1Dyb3rzbilQubcoqxSgfgBTpu/DElUjyUS
0qGOXCS8pXazisqKlriASYwRaBrO5//txuuNZIpqjKqeI0k/M9FzvNSOmFnJS0ML
O+0p1XUJT7FTqa5JYdVypvR0M5nEH+pKW0RzeufJlXcqzVxB1H/AADO9cWb8KFr9
GDPI2Luw+798tbeXctrqi7qmExuc8SxCpwRX822r8YScq2aXjwr38H2gW7IigdMb
CWA8LdO3lsvsJ4pMwaF/VPf6VYw6yLo1quSdDfhBhFGQmI2uYbKSS0+Vi/ET8R7X
SZXav/F1P8cja7Td9XsHh8BtM54mmuzNeKGNgUuGHCYQ3PA+dWF9tlhLc6ElnQKs
3eA9EFGql4cWxvaKEVje6QcdqTGVeRPt/tOnY/H21Hz38e720K/WEeAH6EfgYih0
93wt7fJIgSdFyBg7V2X5veXELsYr36nL6qBlDQiTG9MgjxY80bRTScRfH8yP5H5y
wfULeS7W5ls1zYUdXwwj/cCSTCNKZrGJo8uhoHh5LcneLa4IwAmBWGWc7NLS+mdM
zkju1wIMOTIABzyEM7DTeovDlZITMzoWtcvh8ooD7WnIyF/Ik8T7FKkFdmrzQJWA
KO2hEys42dgeMh2kMMEoqIZwgZRHIHbzFHb2fRQYSZi05D3jXPI+1lLsEMz/BmeK
93kHG3zi7i1GMZpadJKWXm33x7QqLKDqcjGCwGpsm5KJj7vJNJlMBKK6CCSUk5PB
fAeF78fmqPLKDj04ditJ1AGG0T7yvpVo/gfLrr9yDUUkmykRZ3pnC1JsPp+iII3r
XW9ROxT9spuqAwMleUnGsf6b1D7GgjlQQC1igu65x4ylQAeGLgAvECZ5GHroJned
xJkcawAI++B6JEYRY7aYWh+Q/p9DOJEZheFlqwSDOpQjYY/Ai9bf3vnl1/sejtrE
otiDXN0eOroQSCf6v5lLp7romVeFwFhADZ23FQ0trjpx7C+wWfi/gXWqxkaNT721
mkCk/9xzQu8vAPYW9vayS+ys05YwhZVa0FwnkhuA9uwoRR557owk/Or5eNCqW/zC
AzPseOqq39/4s4/XFRxuNCVeieWkAfhnML9Oo8u2R+zi9FQBfQ7E3UVEoRY75y4B
`protect END_PROTECTED
