`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aK3f+TVAZb0xWb8j/MTUIzgKbTq5dsw5MCrS3VNhgj4ljg6eO2AZMDxBiVIBqEZe
9leT1QJmPTSmqgmgmtx//KBHbOeRUJLW47GRsn7WNCfOS0+88nge6Vk+599+NrXp
9hgi19bd65FhOJfHXTIqHJzMNvCZHZ8fSU4jf3CfFBLahCw4+dlsi52SvjArvJRq
LsCy+KQpyuk2dsdWTqpIV1qAKL69MFS4RLj9KaJph0rUAveTOHtsWCVIok6Nmdd3
5okv4+B0Bel9cT8zLIH0OOGvRAqIb7CVAUxkr8HnlipN1Tlpy93gSykdpax2MXoV
U09Y7oTBkMC6WxEguD7cmKS+ShnHlRppK/GXqj3a4opzw046QuNVXUDM/R87xmdb
JR4QaWOw7NMmfoNPk4DO7vm1Xp2KUlxckAoFwLYCqRjSzKT7JcscQAOOb9BlXw33
vGveZbDjS3IBn16rr0LU5syaI2VzYLkWwFdoVHaud/c=
`protect END_PROTECTED
