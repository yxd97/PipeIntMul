`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QJOwNvCBkP/XYnoy20YdBU6S154raMd8C+g9nXVoKNbQb+pJ4/wHYLVcBlleLDJ1
M+jCLnORxOOhpFqbQQbHGSbxCulbtgeHi0SsPNwnLoEdmO+uTwDjOSzKmayzw0L1
2tv/HR5/QkZaibB4s+YVZWPhKmSyYMihTUaE0g3PfnFrJ+QQk9E1iujkNThe5Yvl
6WhbajfVzHyh/q1Rc2FxKdevvmf1fwDxttTlN6CgiEx0AbwPcrdLzUElxubgrAWQ
FM5JqG/CK5u9wgMZy5U0bCyyvwKcbbo/+Fc2EzUus+c=
`protect END_PROTECTED
