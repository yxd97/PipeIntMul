`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4DUEwjFEZCDAUwKdp48rBxMveMFFMiICXAlYmkQv7DONw+Z9+dDgO+AFrkrXtWJd
MEkOvWZ6IH1jGMYA+pN8J2Nc2NDCqAtLz9vwhmKU/i/aEXw0ZPeUxmRXXJmxMpOW
TIRTdA4Bq/kH32MNP5N0TVBoZ5O/FXUHieFb9hcbRt+6Jf08szVuK370OfTYgoux
B9gBcv6Fx6kyUJBKksfuJIhMKtXFvSg+l6V5SRrn+8aefu6GPZ6tMnV7UB2DIMBR
5kDX4gJLtnITSTy9Pex3BpNxtw7HT/YhvfOOK1ELpj3clijPWga8HHKMH9k5TTyn
a9Q3DtV2rbiqCNMXHawulYU+I8+ZFZWXnygx7XZHxex/VNlZ5+aZR5zMW+V3II4t
QI6huQSSj9ywIkf+Wf1bd+DwXNNzF8ehKsHwZijKcdwq1NC/Vwd3NzdcUjYm/lgZ
4KcYn8jMI7vIO2Yc3mS1uf89uV2ez3maBXFmpQYXTorCoh/d/mtv2oNiqVlrhPtj
sdJj/P6zgpb11AWeGBpsDth0eicOG0kWE/EeZBqkN/WmOtuCRQ5aMsWbLp3Qwast
3u63Dx1lt7BTM2/OeTMpJI5ElCZRzgiDFhSrCKER058c6h6JtlvzWiwVkelUkVWR
GU1nmkif1pWDFQz7moSIb0zVGJJHpLiVpzYgndzp1USNXF7c64DkukFK9e1FK7li
1VrceSpEG5g+/brOASdmh7DYLATVLYYb4RkAXKau9unKykX135MiEjByidzziOUd
LkyAqgKTdaruaqa8pvzKOfsSMEc1qClpwNMsZXFNgrLhLb2OGiRfN7LwQ6f6FeHb
C2KVbSvdq59oaQCne1qOd4flFI9SoxjQDpHEqEzCBXul4jQ7NzjTaufkQ9TqBlsb
3Vcc+53TQnBkJXGSERdy5w7o1oK7LI26KOE5apC+AIZ93faMGFls8u9eRJdhuFsv
O17JcpwGK4MjPBsmyPEM40izKKau3GzRDnyi1B2YEUWD9szw5TSfMKjEnIusRD+u
U7x/eUMhENCDlyuMmQulPwo8RUtHQ24AmUU7a/qsSsvKhLZFPO7dzfTVG5sCuuGB
YK+2pj13iRlwH2DdS9cAEX4hSwLq2AmB/XYZ86+xPF2Vn3Tkzr0NiVUDiT3FhgWC
ikGQvMqGeg2yuthRYhieV/VgDTmGgLOugFvJdZoPYME3hDKwyumTrf9uVad4nq0T
gguM2c+DFKaje/SlqgOLphJcc4ZcymimhK5dDC9hcmfsV6dtVhO6Oxj8JlFo3uQm
SP20iRvIsKc0+tqZoKixS54TMtws9RXgc2Aci71SMPJaSbL1RImRaE/FdUgRpSgp
NHF2V5TS0GBfTiFTvPxidvSVEmtPDMmAJJSfWf28VqWGzH+kFlE/ubAeMgvubFVI
NInEkjyjJ4ZFQTT4ZO6Ngf5ZPS9tAnhCTrj6lYxsoY94FuPWPq2mqP8s/8gDtQMR
WPsC6y6qPRi8Enja4i8Ch4NdAQIhL9kAJZyT+V5SjMr41lL11YP4xMIx5SvUnGsh
`protect END_PROTECTED
