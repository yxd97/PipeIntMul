`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T53556xbk4JX4gnedvI9PSU30iiTRE3K2njSsT7R+EwC7ZBeRYUqLILK/W7D3Ssg
pXHRdQtCQjN6Snebhl1IgltoVOAt9LBL0wzr1yXkGEsRBGsf+Rrf4bIBpjRM4Up1
41/MoubqiLfMDM8sa3OiSKBWYTh8v+5imOV/H2xUpV4HVFuK91CAU3tYRi+pkAoK
P5iUN2wIuf2vTbktsKSE3JprMrYw3Fk9MF9lbeRw1vEw5Zf1kYyGMxEXvX+r2Xxl
WoX2BhZhe32425OWsprXOd9oUaWPvinduK7q1yeUM+z5UWPueC/7inZd2/fzMtHL
mYeoN2qGdmkTapwVNaplS0nr22tK6xnJ8Uj68MSRttzoxbjd7SPDzgmP0YtYKaQv
oN/wM8v96Teu4gIdTncBvnlDaBglbnAgxYSw4BapbXbiKAR5JFeXliE1/PkL0Xas
zAi71pkgwx4V6+T2Q9I4rFI6G157/LaM2UTjPOF7NoQsFYxKYnE6cuNPMg0YrPp3
8FC7TWXMWkpQzVZmCbSTps95vR7Kx7neDnYNl4xd0DgEqPlZxw/kDr2tFTb7vo/i
`protect END_PROTECTED
