`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aWxurGsq1hbXU/vzm7wzLJXWIXiaCrM9ltulVvwk5Bgi5bdNE0F/61owuiOBUxHd
nocEltUbkcxSR7EsqT2Z9gOoV0NSWEOdzAiUY0gi3gp1PpxFxEdTr93KjshpivXm
x2ad2NnEFNT2Y0I+0xN6l8BxL1TT3iwCWyCMMmwK5NI6avwHJPmZm+T/rmxCWoqZ
T476hPINLYNv6QN6nIokbCFU4QAr+jkMXOARTPEiQ2Jdf6IY1T8joGW594Q9BLc9
KgNVJpQL5epS9wuaVId8vpho/jVKbh77Ithiyslbylh5jyia3uh2odf2OvHUZT7q
iEeZAVJwf/Nk3kTZy6K0pH6TvrU76/6SVLbnV9UUVlbwBE+L0j+v1Kt4A9nIG349
8iWe1w8+FQIszsx1xQ/8M9SzLNoirXfCLbYx2Tky8rI=
`protect END_PROTECTED
