`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CNhQQGWUloxmy0C331xhyS5+8mf3tjG2xjVeCTnD5hnexg2rUiblKxN29doLUEN+
6nginU/yS7jIgQGHqqwsk6d1MsEeFelleGe+X6E8JUiFHZX42FdHhF1zdNCW/etU
zavDC1AnrmcoymeOJZfx/B4DSRWvzXVewKOqYoxBPOJDF3hcMPuG1kEeaOuJQQak
sZXrNVQPeISaNvUQkopQa0MBl3D+fwcZ1TXmhSvcgz++dQNwqjaSU7Ks646LpJUQ
fGp/JHkIziqcHuDs0sIpVwlAAbfHBRsLkmOrwWVDNqtRnHUMS5AElWnJQlMJ057i
lPLa4RBvx8VSigrUxYJPu9qVLvMRN1OlKTBrpK1g2/d93OdG1LMEZsTEkx9j8z1S
fYgroHuZTNmvxpboNS0bRptaUf0fKx+FdWXH9S+i+tU=
`protect END_PROTECTED
