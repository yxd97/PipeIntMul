`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DUy4UnQ/fOHnitLGi/9YMuksy9zGB8HXOAEBFtO8SkwMNvdPMvzFG4Gv0fTx2ADO
5W0JPCdIlKqkixVRrG/j0FJLA6YqCBSlvXHmxqo3c0miDSljl4SJyTKI2AlIulT0
bd/a5TTuaQnDdvitUQf8HrRkHLtAraGJ1LbFV7AqosqZJ9M9cKoxE5nnl1rdyAlg
55pXpkXCYzks5xw8ZZ6MJYKLRxp7jpHtJV04y+iHRBmQnZngtL/sgx9Ys4JZoiwx
t1y49UA0fB8VmAeBd0YZN4aGao2N28Ag8Y0LyC5SAYJ3GrNo0c6q9RNWBahDNuIb
lzg1ZJM+OVGQhDd3s+ScML4j86FisiuGLGG0qAsLeZMq3Qve6SThcdbuouYPFWkJ
5VvVD0d7Fx2Dmi80tavzLwwqBiN/Gdskuvy1f2Y9O4orJ449Vxcbo5xs8S/ZRmYy
KfL8vnG4nDd6UCxGFTKgjw9wrGKm93ZfwiSSED8ajfBQxxtPWZ3it6xVFJQrZWbi
`protect END_PROTECTED
