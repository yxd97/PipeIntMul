`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tJ9GMO1CRHY2b2VvvT393OCnuvOMPd+YUoP5gU+vfymIyBwkWFVitDcCtOM3agvy
m65rdUQaQp8YMyWW/zhWsU4U//Q3JEe5LmB70AwXE+4LCSJVdH7vxAT6irxhRvh1
y5UZV8MxHgOc3WqLTXfCjzUa8YqC4Y+z0l2X6+dJIGMGORnu5H/jdW5upBnA1e0u
yqYpDl5y1XyqgmhpsABu+LKa0vxmgdgQgFItgDm7PK0zq7eLcLMLBKLQ25VHbAK1
3SGt5evUM0IPGbw60XueWnbM9JJ6nB+jHeFbjbQbBcisL83AU0gI9conqIXi/rhb
qSdhkw4otEszdzihtXJ82cH6+uLmjAciHJbzFtzgzdh6El+nl3qKbhnMXfJ5wQKM
la2VdTvRt/2zAgMA1kYvllM1e0+z4SJcDPnnaFYyHz+P8EFtN8bSzCCuv0EPruTt
kOGfaI97erkXMuwgQDaB6YqOE3yokBAOC3G0Ok5kmnmeEut4oXNgZb0LQqosca6Q
+N/4W8Dk/rYeCvqcYu1jPagScYC8LK5y83v8mJJ+1scJDtptPIM+ao+IPFDWyfm9
OTwnZdS2dDa3HQat5gNYRUobDCXDSen+Y6nprtRdZMegJv+1gVJc3sKZPAZVLejg
bXYV4hPS7e4RBPkEu4PZz11GpKlzJQSWhejVY1arGlCZ6BZRkm4yD7lsLx2yOF97
dXEba152YNTtKzv2Kx3wtQMOxflSJt9HU7ROYI1b65mBRVcKyw6MmjSYcnJGMw4W
jZv+J8KoqSb+NxJeRpUjOpOzhUv4Z1tIqoQlXB5vcWK4OcZ0jG73fs1A9361tSN4
3DN5YShu0Q8KtKGVXjeIKBKvsKKm8zJRlghxzCeZqOi2MP69knXvMblEpUTOdu7U
jM+dbR21p98nJfUcg+X9uDbDFekkq2DSG7b7rvEAe6dN14NrRDFK+niGu3EVNrxY
h+xYuvK2e4kjdooSX1FbGNrZVXMEmgo912sJN9//v8Ej0mxUTLAFTMMBaZjOwcdK
RZB8CHH3hErXvhJeqfzsdCXP/rI+TeobYPzLCj1g4uGPsv75h+IYJCrbIVf91QcL
qGYD/mY9yU4k+4QOKcjM6xYXSiVF53xNXuN14EwEOqmK2VTIN8D27ELYsQfI21x3
dvn9Sltfl/kVSeU8XGE8/LyZTNigjZqnjE8loVUu95Xf9Cps2djgf+5LvJ5ic1za
AD2BAj5V3yPpIlWI1cm7syTkidLyE1efT1ZPzS8rtIinFgEW7ZxIq8AmMnBg4+kj
+c1KDUAHj85PQ0UR2Ej9mHoum2IPb711ZET4SjBOOklsw7XLjcOso1/zrji7SQuW
kAKS9Z+cFZ25Bq+x/PDhZOYyyCdxtIrW+p4bjUHRZmO4T6B5g9PDII7sq19+dA0/
ch7kY7jOTxx2diUcllTb9OXl4uS/yW/4CBy63280VFQBQrd5crNC0PB+EPc8lmGC
2mqbg1vObLb6XeNGw+ILj8KeDocEsI3XnMzdfHqFsABGLRMeRAmHibHzkjDZOMEM
wsyKTPC4fk7khJjKHuXkqKb9P+GlVjqkLKPl0rEFpQUYcwq3eJAdhgh3KBNsSX7o
menvArvXgywug3sxCzdyToB37CsvSc4R7C8qNkIIJNeAmETPqo9BF/aG/skU2lLH
EAEWBSX7XUwXLu018Gl4/lwP17q6AhJZKYYEhk2vf34yMwxc65FQOq1hIDgJK8JU
LoBAIgS2IAEzp/NiMnHZObZj30e201L0ATsgEwFYVNiEVzASMH8hLm/wTDA6f6gl
FhvhkP6PJYC1J62OtXUHDWbyl8tJX52d3svTRkGnXOQrcSJ3pyLUU61b7U0JDBDp
ZbUTxflzupkvUt+zER2Iai70/LM1CVrTI0vWH7Ijd/4EZ1Sm4sZNAMro/RcHoLJe
Q/rSMaEKzAJY7sT6VflurDHSrFU6vRXX0+tKhz8pTIA88MIdDHOd78Ng4189hnyM
LXqBfkuSC787b0ky/leArYdUSBdZUGkEz0rneuIYQIvveo/GyqsUJHDIW7OWGOhr
/9U1qzcnyVy3YnqhpqcYjQ==
`protect END_PROTECTED
