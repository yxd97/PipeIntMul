`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9xboWC53Id4FRG0AZwGzzw3A9ll13XT/RIH/MF61rIRpIDrjVZQDYG2hDJvcKhbq
3VSKc1B+VWNIxb/gMN8T5MSyvRpsINZujSHzlSrrPOSMBGLlNZQnVHl4VNxEFuFc
9FJBMYK50dyvYfyw1gDCFS85m2J34fwDDkOp7eooX6OvUnN2uKh9VyNrmlBqQbHm
v6GQWupwe2kLgOo3KUmdVEI1vZh8XFvV6AZeUKVoY+7Twc8iKtNvFmeN45lz1/y9
omgoi1QyL5w+btFriK2hVeHb2/XdeIPgO0mGtLgLuDqe8bjVo/uaTwACZOr0kcpu
kmB9gXjyUZGmWe/ExPmwydLEn2MDO92qIewPgF9m7riiPmpK15SekyPRjYeeD5BU
f45qGJn1v8IxZ9obSBC9SGYwWyk6RzfYHYx8SbaeuyRDSmwJy8vhCkhYLPti30a6
dst1vkvzOcF/W1zPvthc5hiOP6bdKmHUT8TGH0YOKtJOKK3KogOc0i1FSs7R8ZPC
IYocfFOSeYnXnfynA2LsE+LJTSEFRKjFEr8/Bo5etxj8ez3L1Cn8JnW9HxOM+061
IE5CeYflOS71i2CIpNWjoQY+TwRgdqsTGk9aVRTJORo2fudq3cmfK6pTG+obEbXI
LuAW5uv254RtfS6QW0AM3U2lPdG0UHeEMxBm9ZEa2sdz/ulrUd80ZyhMsMYf2peS
IfF/QpN4IUGv7UYSVO11mdup8ziVaJ+vNpwxgCi6fXD2z+4BhyAcu9Z4ShVdfWRa
BmYLOml5oKd12GdJLwKrCJtbMJJr5HhiBjAXl41n/OrQb4Wf/G3tiqPsqAA9QKXm
YwOqsl87RrdwfQkaVZgdxzb48pETPAtfkk0RxCHxFpP+oYnyylskidhlQ4uIKZ8W
fyjpdZTPw1RcajxI7WEmCdQ3LnHHYZOtv7m1DloJ1zvewpTgWvic3ML79KAx1DfW
`protect END_PROTECTED
