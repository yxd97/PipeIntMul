library verilog;
use verilog.vl_types.all;
entity x_lut3_mux4 is
    -- This module cannot be connected to from
    -- VHDL because it has unnamed ports.
end x_lut3_mux4;
