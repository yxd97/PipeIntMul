`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6lJtiIRthWKUHY95/03bH2rDSHc2CyI8QsAVVnO3yN8CzfaJxV0xVf0a5/txGZak
u6TZCGZjLqZ/Ao5LSEE1jW+srdtYhgGdaX2gEYBpB9clUaUcy9J81U7DnPRzXiyZ
66XKSxjFlYIk9us/ZTZo3+lzocm0ikXsr01ABFeT/cuYLT77lyH91ewomazhjeAD
AYLyNBFFMofB6QkFqnJgTH783p0mCM4wx0vJvys+aZIiWmitCtVJ2kkcJD42EVSr
ocp+u8nBhor8EMSuu5016l71OzM2r568dpViqJoKhqTc1M1UgQxvOqpZ7izy5+EL
MfTI6i8q/mJ3hUu5BhYq36T10/UuU4xTDkoX8NdkQKblJxN+U5B2tzJgz60IOJKE
CtTLmXNYjmoQJ5sEjxwlDg==
`protect END_PROTECTED
