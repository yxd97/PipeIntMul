`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zXXVfDCRMNAnUxSRHs0P3v+dunyX2ieJULLasgzAyGWN/KaI2WPlO6lyMhHx+/L2
HnmDRErHbRHPttNES7iZlmGim/LuUkBX2Gvu82wZxR+mm+2MlnGnYI2+ferTlFtT
QrSQD/pBxLyRCbfl5NOXfWWkhQWXwl2ZKhkoi2JQQMGIhZZ8f+dofqkNFQuvRAU+
yT7U2D7WFoG1gcM/3VZ/eVT9CmtgZPGgmqiMSZFqNPPLmeZoOkkHKUKoTOdqeKKx
M4ZaLNM5xj1pr0WOa5lMMPBDlHjk7ZKmS28SSlcZSlnBX4SA4bjEbkGM05K5Is7f
tSJNYNF4IcHaj1sk85Uhj+X4Gu70LArCfemXm4UvCSe/GOfF5Yln282dT+g43dtX
kguCw8OsVK870Rq6k4+3PDGNOBOsjwbEbxKP4Hl1ZZzby+u2XLi8QGaIs/o3z+jM
orvi+VbIcsqlhC5SK06CLYkxiqsBV/gUlm57j73+knMnD7tqQJaIiEYdkVDC2p/E
sT+pKw3HIKUqlIneSY+YL4q4vmVqbgGb8OT5HHn0xpB2Bp6fFMHiaJJWd2m5LXqL
NCJ9Rt49vfze17fGjg0xDDQs6LsHTfSmMW1IoN/4Mruplaatb+ZX5RAeUft02vch
Tjyapm0lEtmkWX8tRTJ3x/sOy+m9KPijLibOB/YZyMNaPwra4v12bU/AWlbwYRHg
lRZcjev/WRX3aHU1QHuYgxZWH2AaKdVUkQXF5n9QCjbGjZ0pruhfW1t5AzxhlzXS
+ypfydCaCU0/S38ZN3qPFov9jCWMpjQ05m4sLwL1KUkX/1oklR/IaaLOWlB9RNPE
8meyuJMLlLdDx6zmGvpNnu53J6Q7Vx5bAK820vQgNUhaP+09tyRjikA96Ptqd+vS
cxsMDN1keqZGSa4eY0eYXHBhMo3FRufc9maipyhRh9vmQf9OZGhWHxx46J7njwD7
GeHdulyg7UHPvRYxC56gp0wX8FnMEbPRCeKqtGKlx8IxjNlUmRUuWc4TUGw0WNQx
VlZg1o3BZuF/VTgaqazDkbQ1LfiBYpW8RgqtFWpXPRz6WewWt6Q2aBFQMs5pRR+v
9G7Bozk31kdy0umSARon3f7zznu6v/BeNC6P4mQVHBvoecYXkUjmOXFODGw80GZV
jSD1WW39yx0wrFB1FBfJeztM8c99twDhSGuPICT9H3+uRFzkjwJ64ooeCw02/66R
BRodJ8Gcw1L0d4ECc7jhrnS/SfSa+beWYSS9pRVg9Btn3T+x1RSzomYnZ1WEFbUl
ZW4Sx7FJ8FLN2MwMwzOlZWwY3gQfYFoXf6Tdc8RZavIAilLk/1r2ZfP9eOdP1Y6/
4a5Qo2vN5eZEoN4LCSE6/CIQFtDPxULHN+iBZpiPTRSZ4XYg3a+yJrz/ZTOibSmz
T95g/gvFUodTZIn8ttIDrXvOPSk5Hu802mXmvsUxOqs2MRhP1ttvQ8QYIUsj/OTJ
XLBqAS1MC8lVFNDzXIN94iPs3LnveNiuK4QNKPSBzvbgcuQsCc9bl2q/E0qv/b59
DdpKmwvNn65UhSCqLadONv7sIJunae8Qi/cBLG5iNIC3orkYJyOpx2afqUaQN1cb
veKq8nXR+4h5YCeuJAvFEQfTp5I+iprBjSd3r7N4pBODO++cNC9ODg9oQnCpJuEu
Sxz2/hwRtmgk9h5vuHEGTYbDdvvIagMEQU3H3W3w1QEyg96jm2c9gkoz5aYuSuuL
0HFO/1CNO7HNTAgiSJsFQel1LIQip958jvs/zmO9MbSzK8/Pr5diMqtsH58M+Ucw
U5y2310d9hNmF7W3M0syhgokK81XSIW0BJuBG9okUp57HSR+7ni9yY0dwK2lwUDu
B1mbnO520iVOrKtSj8ot0NGHxrnXM0dEaD8Ts8StlFMx9V74lHl0ZtkyN7vYHcKt
TW2UzlCL11uiqjNB4aE6Oz2uUV3eXHR3l4YR2spqqdgzRQoKrdduTQHOvbAIwsw4
O6OQYp9QfwL1m+N3Ay9dNbSFtPr6pUao451hbUSV/8RIomn77IOc7xTmE10P+FIF
SswRsNCp5l/3a4Ilcykl7kwkjVsC3u5nZ1Cy4X7Sh3qNAyvw2VGmQp8czY1eX8wL
wUUiHkN4yTAfB+v02evunjPOCV2ljZrdT1kdUefI+n5xaD76wd6EplZUF5UmN0fD
GMnlLhzaFqaRrf9SUVU+FFZKJNbjmsp0eRMQgsu5pPZFsAzxu6ZPW7si8uBc2dLl
9dBDk9EJxKKFkOvMhvM+O8TNgKj0n1/Ocf40rq4bToVxlUeKIJdYOAgaqMOy3WMM
5IvR4CPkaDP3FvPENInk8W5tvwoI6JEsHW0BXimOGjbAus9j0zPn9mT9xChK4noA
xOOPlrscqLz5xPquzZMhVWo0aWBnh8Rzy2tzTKC98hffGdeRU0dbRjO6nZg0ZFNv
s/zjNNyujZ+b54vctdejsbOnusoLpqbxhHK/UYrs0QcvRlwCNVJV30TKSQlHiQbl
iSzyvYvPT8vzN8GZuzGuieMMu3HQ/BBS+9zuBgaT4fqICwG0gdcd6LDatxAnPpdP
jv/QHkLbaXhEUTpTRnn1c4rVg4iOIi+Jcvk8PnI4QpS5u/04em7Dg/IE+Wt7FJfS
GNeUuiGFu1tnOby1H6MSGKb8JuPR9N6Df52ZnQweJolF8Lgyx4D0Lj80z3ZOo4RI
gqNjfLTzzVWE0irocZPNuN8UOCm9xv1MGaKl6Xi1zRZ7RbSJM2Y115Rkfn8pa0k6
kXwni4/onkoLhZYCREdTlvRWkxqYYxDpVR480dco2z9ylXHfvPSNA+wBUwnHQdyD
XQMChmxQJWXtY11biJtkT8A+905700tFNVcwy3pVYJ3hp5U8aNJA1dVtnxdJVLN3
CWnGEZONUpT9+cHVYet1HoRY/TdzRtwydh8sn1oBtC6B6biyeql4i4BLNOmq9B2m
cUjAr9sbk+fxRH8YYyvkAV4BX5xuIKCFcO2yeFHURrRqJ6rK/YR2E1XhVAZnhJJZ
IG2id5SD2KJzUCCEVRH3i6tE4PK6Cj3L+TTEJCbjAxVHMl8Y0PolrnRc9w2cwrTA
p48NAYkeVqHQrEldjOsMtjyhea2G2IcLmrHw7/i0sFlldihvSJ5/b/3b6HUnESjt
MPiVauhVX/0FnP2LHDFGbEI+aikUvnU1AlXronTXX1gzzFVFqmoVE/8AAd2a8Lcw
rA9/0jN+EO+LsOeuS1zc8YA8xVY1tYdwA1Q6Uywat52JWIuwJ17beiuv35i/30Ij
86++Y1yaHhoDZTy+uVAAaXxRxG7mu4MYbna84jT8lt23hIN+x6X2ZIPyfEInymKl
g/er99sUqobm4T9u7FJM6vvS8Qi6qC165p3BGJuWvnfYToJ6b9Ewj87tp6RKrW0d
x8hxX5d89isf870nn2w6uoSeQgZZ4JsSyLxnPeY+zBVAop40M5x6mE7lEMe8Eso0
8h3HkBq0KUEiW7X+h1obnk0dWArOd/6a1caamIi5Rqm8NB/Ali9KZz6ByG/zQDJ7
8OY6BuDTL7DMlFfEE1BhORsjMwy/Wk/jgQNnCUBax6CHD7VTy/L9f5nIxndpGd1S
EbhewTRaQgGfZmief2epTuwmbkUVbisZLFrqByOk7XPNHqE4CsGl8jktEUmV8tp0
wRAMkg6H2zgxEK+gMdLclar8LqeY9hKtB2nrBE01q+YsleTGnSdqgIRxoLC6jrbw
w8Qu6tU4mC0540/2eYspl+Pny41KBkv1ro9RqMO4OpbSCeac3QVnD5j4hgqJ6iVR
8Qp40WLfvlOO7IHmBInkCcNV/dyUURoKWNI6q4asqi+7BrUVsipkaXz1FIb/vRvM
rVC2MRlfTWomT6hillimcLJG3iDppgG0ik1J8OsN7ZJOPfuI6TJ/jNR1B39PU2dJ
kg7ctUEgeGQiGY42rkJVMCmq8e3C2ajYaqAeRsrnYXpaGcjn2J6dWEGbbB0HPjv4
F8k+L8NJwjPHz8GS4WRp56DISbL9oMgAlny8ccAlYTyHMO01TiBu5UKov/vQXtAR
THOB0Y5GBbq55mdIcq8fsKOUAN0CMkR2FZjRGc8XYnn+bpOXOdHIFbrW7EuK75hO
FHAS9+6PhZp4TdmdjJlc0GMrTuxT1ddoKgwlVP/DTuvpyatn2KvojRt1wwMUqLFd
Mmmk1GxHLW/aWswnVlq/Vh/98N6w0fsc/6uWzCuI4sDL6WAF5SDZs3/cR8aliJMx
ESB15arrNQJsPa1i0pZ/JzbUb6lCl92SMzNQBhbDB8KaxImg97R8/yN3I4POnU/Z
c/eRXYcArYNPBWhqsmS5rGhaB6YIcPH4Hz0spvFKF5TYrBFbLedhU7v/MAOjeWAH
Fgga7+AXLgfm3dLhiZ5fDE3c2/BipF9Yz7xv9ssckX2C5bvR+6xCLlVyQVYgG9sp
SKvqkBvEncPLHmD/fHiN5pkiFFPG7ZsNYgg99VysNxVWfqMaICM2lzVPWXN00+B+
PSt08t5se631TFUw0QNewH/VTyLZHvYugNHSE+z3KkHyTun8bKz/eub40EBn8dzb
WQ+rPV0ZcTV2oJXzH0l85vEg1vW/VVLbt+/MVxB9STrVEmwIlshGwvj+8XuKcNu3
CrBLUvQ4fGSV6/HDgkWlDnyCBHxLwtoidYPK1AGs/OVGqiKfxYyWSBYkMMLLi2ZU
0qbMt9LFgTSaXVTZ6S5kX9gzMZc/z386aRldmvk9i2MpjOvpqp4AnW710c5fVQYU
HHBfdg1Pxg/P10K2RD/tfA2HwNLlUuNn3z7oQ2rTawVAj40NO0LPSWOOUVs3umoE
IqK5oXjilqGid4D3WXo0sCV0ks4SYI8X5GVn4JaWRwhnrIHW48RpWjTfrCEP1YeJ
HN6uljr00/7l2Sbmiq8EqPNHEJMW38KUGdbrI+39ZqwkPzoN5+oJk3yTWzFMXsR9
RFurSmsJIRl9TsFaSmn6jmQpjPCK0AqvJy9YxQIIHfirQ+MIE5lRGO1kESud22e0
fS0lTCJoj6U/2A+isEykzqYoJ4VPJe5S99m+I0x8miXVLVNgGTb6vgs6MA4LGJl0
fuIKOACWGlxB6nQOyb6/b2bDx1QtWhTU3BQpydL+35UZJHtJOsGBKzOjzNshdmAe
i70Ml8R4rxusrBAWbR169Ye89Y6czcdiXAVJsICsdw+MPSAUtcxeVVRZlQAU44UB
R+GijNe/r3/MxRQlUOZaW+jG0FubO3BzTI/1ZUhXo2vDF12peJfE5Du5xsSDFU3O
70HAcozRszxSxvkGkbsQBU7/+Mo0aWgOdkicpVuq/C5nyZ1yqcJQEetbiMUzAT2z
dPNSm9rmiIFBehAg0GYuzwl3vBsvDgeSAAdxpkRre0uM/1f1dmHmRs4PD2ftZi/p
py3zorLCoP4WCktKWt3vhCQIFQipoSwft5cpuk50owdf8Kdw+Q19HEJ7PQTz5Waq
Nsmvz/lFUK/FhIalcyj4JwJIVcuW6U0P6EeYn7ncmMNL8PPcw43X6TOjvpBudwcP
PLBPFFu7t5uO5xf7eq45Uvt+xSXboPLX6I1zh64IZ7lWgHXS+gfqu15bN0da+t4q
9HPfbc/GETE8LpE5agEnWachnoSEGV1/uTUUSKdu1Iz+fxjWAv2QflR5jKit7V9e
HegEk/MawInf9/r/unWtcygdRJm5jdQMWEbta5eKKAUyX9xSgj/Imw5OiH75y6qY
zlSWxRflVbHhAkqnIk8j2UWIIWtvxWTYI3TmmZUxXy3rBPkpFGlomFFai7t0h3eQ
zBCIjbLKeMXNYA0j/HjNf+9M6AlDagipUim93wqAyLcqjeN3MMC7po3JSwWR21x9
NuoxSQkN5NOKXM5wmzrW/ZZno0Xcks94qp8Z/+NQXhLiylnQWnXbdWwB8S6gFtr4
GD8ibkHpnOxkPsMOsQ729xHaHg3d5DwMpeaPjSvWMRBynmisoXFodAIa2YgWKBy+
teSbrWYHzDYU9FUYqEjrVM2p902oT4NZsZHms1Es7UIs+ppKCecK9WxdmtzyKKCC
hc32gGem71UEPwFPchwUTVqyBLB9zNoJp+D/zGigsgiCOPw/cxeacgWgHLEq0PB1
XOuEp4CBqhKz3nrppqTET5gSHcjuysPob4ghuDOlHdy9a2+70WRSLan5QHPt9J9d
dJXnCdNUnn7xT+xqNckKgvULCOM2OQ1J4MFGZpuVgwpxQGfqtquv3F23DrYWy9JT
zBWGKFOgOUs4mvuPoKN8nu3yGuARmNvlvwMltFVUu7PT5mII21RaAieK9wxlhkFL
E2QYxqdpW0rq4I78ImvKtBKIlROrzKqe+9iDykwBmobQXq4EkZkLCzv7HwedMD6G
BdzSePuC+HO4jOqAo7KA67q+eWZ0MlpxvVLEByJCvhn3hhM23I7sORgCJgx38sqS
4XBLYL5UbvpXzWw6fndjqAU084rs+MgSw3PVx1JJFELwGihLVsGU49gi1BZdZj7I
nXM31BCvRQw6c8rJUGamzBHqO1kOMVjg2hSThwAXe4/82aX7AQPINCjnVsm1lnWG
xW+hhctJp8SLvoPWaYB2T+jS2h890mR0lLarsR58H683VOpqFuNG2Q8305YxFEPu
BNCS6gzCJHY9SV68N7MWCfo3PfYETohg5N2qWUvcXJCO+61yikbVtqvPSrbE0076
xiuuaZDMGZLDeEgJrWVBnGl9PAYSiuB35FqKoSG9h9zlL5inf68/ISBU0FjK2LO1
mhtY5gh2coMzOydIgyq63PWw0oAxluJao5o12BSKaVsHAqIx99jq5ZHNMB0QbQnP
BtuGeZCOk68tL/FvbinJqkIDiNqkez2IH2h050YzeH39XfeFtvINWPDLA/2GTAfN
PZX1TIJkT4+Ga08B/yzz2D4tI1UTt26aC+S79FJZZ1cGUyGsL5jF9qya67Fj/aH4
dPBYbbNkrAG+4mNVskN8ZxUEbDa3XcxUWoJIV7WX53/698sof7KXSV6yZB9kPx9Y
hDbba1U4S6zzZMifqI13/62lci7njU4eWmXn6+qqETjRJvqLUIjjFmyVF7hJGT0R
EDba3HjGKeMhJnLeAubv6BRen4MWbHdVVD9mikdbTZkOXKOam7lM2nsf+uFwNK3c
6bBAWX+f65HEnfouWPjpR6r8XxiI7lLbIYq64zjBcx5TcL8a4FkJV+oeTJly/2Db
RmZ4a314ByZu7s5X+lewopCFbQAJdf8+fvhQPG6KfTDUZAfuqQEZR3M9wPCBKnTq
Jd/cHpRRnOIZBXpez4PiiPHB60kC3d7seOYZ3s6Fw22WM4b5j3Ui3Fy6Dl2dHGd0
os2BM6d5EKvx5yl8BvIsiemft8TLmUuwB4ptWgX6jIPax0BY6Tq5/1x+5XXyxpiM
m+ToVbJjSk36FmaHAVUVG/2hvstNfq2T6cTfFU4A4OgV8icw+stdduUlKTv0lEtk
mdNVSYkdsaC7DZ7nitBCFThxXRtu3ldgu/PYvsoouD9GnEGkCX1/EJhAQr0mcvLJ
IsYZuewwSpFmJy9qAnavPFmiU0H6KuQA3GEMOWeGx1o1naJeYcp6pk+KG27uJXZ7
Jp/mbYFmM0ZAF8oOUZ/B14cVSgtb10TlZxcPSCVQWTcr2zhKV9nHG7TuyiBiknTJ
1qXVaSTy8yddeEwmiR7RO9VM8g1VfNp92259xxzF8YaBwwfYNaIBRu83ialIwTvR
oW5HIYuhEmQuo9mn60VWOckQ5Q2rEkVZ9QVzUSzFNOMlR41CXUgEve4how3hlruB
zpsGNU8wsBawMhFh3Y38MeGmYzhtR03XMP+hJGMl10JzhzXV61V9hpTqivo7rA11
4qrRuC761GiTer7eXa0Usm4iUtUEWHkXZ+IssY6qout6vItMa27F6kFP02iR/ssa
55qNuFuPaSWiO2aQ8GV4mQDR7W6fKQUGKaU++v0AXlAqGffBFendSNdWeNyyzEW8
/F4WhIgG6nRsvowNk1+plLNEkXnfMHwej9AGm8v+lzhHa8VIId0S7WgEO5fxIaR4
oVzAsUfnZve975Yz8pYTMOzKFm2GoTov4ED7JCuP/tNGuQ3znOIXbdWn15tC2Hlp
eYDNUfGh14/msf7RRgbqhrxwD+FAvICclmoJuxxfdsFJqmwpGId6Asd4g9Dht1no
dDtlCWnwS1PQiv8jUJID4A+A537AvT/upHk6Yaoc2NxnJMSS+xU7W0ItYVa0C5HC
gEgnHeKnQFfzlwUxLxm44VQGHydmeSk9kP2d8gd+FTY4GalELFI2fHjisPZbzTU1
+U/yPRIMt2mB0ywZCURbwcu/eK+TyF0B+kno96xGMx29mSZXDXjByNQ8N6N+mP2M
YwcS/L1apIHxSkGB9I+Q+8R+Yvicwmys5O0n/ENH4jY3zGETQEDAOJ+RJY6HteZU
t8ik6n8UM4tZTe0p5kE9nK/ZZ6dluySK+wplF3AvmJ2DpmMh4yE8gQp7jlSAlRvt
JyTTDkjtsw3OpgSgDocgoJ+5Gwf2EXC7aYQI2fL5H/U6A9xeoXZK1qMNF8G9lCQe
1y8BIVhAGWNUarfsUz9jwHDqgqTZuzsHP0AULdq7YaLfuVCTqpYwrtlwTbpAqMz9
5cn6SDSlxluIAQcY5n4TkjX0iuAFhckiheLm+dQc7z75vrqfWOge3pyKhDy+tko6
Nqb5MZU7TvsCceLjWLNHkWugucpMwN3uDhC50VLexlccmbHgxN+AEg5cmIqDFheB
7EvGm7elTwVKBilHDfsgOAw1qQHQzK44niUJklRvI1ZiVVX8lDWbocz08aGc5jPb
jIiIlvsW04C5bgkZBAMmWd5uc/tdzMbmdq8SnIL/8xEutU40BgQancFJ0XyDTsgm
ePAUzoJcbyh/e9bJH87m6D17m8HhSFSxmGga1ms3XfczD9AS+p17FVIzMOgnYQz4
XnNf3uhyb0zWdN2ZCGMI2tcRxDHzStTMyhaL5sWgemDmjNGJgkh1ac82v+Yy/PJQ
VZ9zQtcMxMIaIspaamhNqH7yR70JdiwjNAhsiSZ0XsoZSGvS82hSJuG4dV5R5eQz
H7b70udzxFuLR5qfVoQ8ddAV5GAC1vJJSMNpTJ0V6DsAoj3sfiegiWK5rbpY+8G6
5RFR+KnXvszkJwp5C4WzT2XSOiGYcEGGnQaX77rmFk7nYQC2nrKM/v2dy4Co4+3K
IoULbvqYu+zHLwE08iFnDXpRdoP0GGWK1QYWcrbB2IKd0d/t66JqfiAVm0PegklK
QK2L0zjM8Wr1/S7vzfSpsF+KaOFaD7a4Nx4e6ketb+JkP8THqqSKov0Kx/w17Axi
T1RKYdQcH8s4mZaS1MOnJcU4LLDsZP93dHrjHWecqa3VhyjZVn9Ja9AqUh88ZZ2w
z/PPayWN39hrncqlrBuqsMXCijAM5V6cjWO0/zI87tPsrvHEO2myFCmG1jPooUv0
9zYSGYkS+UknL6YkgZQjLr9eNgEO1Sx+JkBWA++Lsr1+tI/7a3r2ZXRRrEHIJvdf
eziXqP2dvkSQUNdPABb6/Km6UGAdMaXu8cDHMbVUjdu1G3CABg5B30V4KIzxIbf4
94AQFcNijeqx/hmf/7jA4Rzi8X3RieVKG1UuWfrhuOA4bxnYL5v+bEkRNVtoPrMb
4gUoQ9rNgYfUjnhlmiLvRtuYhw1gy+hA1biygVq7ol30FH+rEgt6/ZbtKhTN1jFW
6DtKj3leLoutg+B0t/niLY/0m0X7w2SuiZaofObc5VtcsuISz24eXWGGzuuZRX0f
Yvm+y4+KeNjc/0ehLDSYYLBJL4IsuMbPsD77nwx0t8fBxScBdv3zbECUs8mvsJFS
0wugWA7gxMcxNX/iZGs3W8fwS804CEf/i67sa4GlciI8Xn1Zf43oKlnvV3c4sGrs
opCn1SMQD64dKPnW51aqus7b23ip+D7hJFz80guAbU6mkrV+vhu8BGOIj+PlFKmE
Xcc6ssyZMQeNuVGeGAxE+Gj1uuxVWgKSvCb2gKngAssFp+urO+pdQUHg/Yj1nAvY
HfGx6cFoYM368u+tB53SquCFPYz/Hyiqh90ekOT0F3loN/lcOcNk3BHR7LDZXiMP
ljzDZUDMjuKCxhtBCdBL39kqazFEnrn+ZeHp63LDGgSTxoWyrIP6tfm/LJk232yf
NMmaZJmrRjDWfyVA0qLIw6zlf1HUfR3BumVd2cQFA0sm4CDA5mbEYVk2hb1V35Pm
QbXWXcWxZh+yG58W5F/58wTUGdTDpgMhP+ir4z4BcoJv7HjPHY4Y8eMAFpJEc9xH
xsbd9aQS+xrvH2hBx6sP+QD5HhpNImUSvljV4zSrNNW0Ok7m7gtJzLLxxklYLEXR
Z+2EoDU9BMmzAxMKe4CTZey6U36ORhp37da/nRqqja0qb0o6AWFpUaHxuJAhzbWy
JryoTsV3MVTkTrjTTgm0XhdalwZDSx9ksqqbBMk0+kd4zW/u3gpKA/iSmc1WfFY0
D0MpyBtttJRXe4khpdSzX30+N9uXDNT745EwzhABYotBh2RbHHhpJZ8pPBfaV23G
LsVg+4zx8scNJ0uzSHrXVzjmB98aPF5+yHmoWQwXdGn70hUumXG8cYPCl0sEv4mN
3fmPoNMn+rWhBq+nAQEQx33l+HTdx6O1mcQN3XXBJT1zg2p9/rsNNYLSeYRxIk5+
q8eF1EsdcXEXtSvXeThEivoHthVX+tJp9cbc1682+eZCSluRT/xZefs1dRq3WS78
7qlu6Q6XcEnWDV0AcT/IzO5GgdkGS4gMxIjaeLxOGOHeJHkt0H1ZeuHcbZYuAMdl
MJEKAUhdS8+g9LCdFXLvRvt2fC6zp8PYGFRlvTYAQwmC3LH9GVdM+D93FbGx1SZ7
QMwJZTYH2MxVIMUx8QFqvvlLHUSKAhIQcH7y2byLhN0WsCros+mUnbMUfnYTQUWN
fcwbT4pMSbpDPyo74BRhQe8cLObdwhVaWydeuUUOQo9Pp2s40xPkSkYMWMxVLvJx
cQatpeXFk0q95yCpiOtAqvNC4OFx0DyMpaJ+YRAmUjFtj4oJcXbI0eOseetLZ/zl
nvbH203eFGeEE2Nxpc1YoYz1mN56UvqHRxo9ZtAF6/11E3tYcOmpO6a1aqCiFs58
qmyFWYy7qVCcxojzBMNRJinAz4NgmijUrF2L5W25Dd4S9H4kXp7YhKuNKTR5Y6Sk
bXa45RnpQuEmcN3lFgQvNxFzdAKQ1/DJmN0vjFz1JwjawGBotKp8h0chTHJLOiU/
RiSEN2nwKOjzhYq+KZNfInLUm9zM9oLkVN1fDGhrmFhY4sI7OpsZV3u89vw/Dx5y
2oqC0BRW+rMU8qdT3Oh8eds+xYARLAKYYWFOqtsi/58lwhFRALaxOEKa2injCC3u
iEkkGuBiixpMPlu+vVBv2G3xT4s1QbDNcmnGiFUUj1nWiwSktQEMFc+wsIHcPr7w
PAEAYRbn5XzgS4eNL24WG/KIgheCaJtqry/UN6YhettApw2M+aRaY73VH+5xVWik
QlBNFt/Ijpp2kqi6bxzcaWoc9BNVYRAA0m8haAzflzi+L60PWt6+bpKIYtTTSl/6
0/gf5uBk/O/JwiPIi47ibRfS0ZcndFgQTaQJbUPmcZOmbIh1y0Y3KpMWSiJtQikm
Rl0Iwf7ylRZvfpu8cI1b86BSHQLsK6/xUyrIFhbkt9QXrUxWLaJU8DkdbnpxF5mI
gLx9fUzJtZYNBP6PY6BP6Mw2hyaAB+uziua0HfabKzf5SfgE9bnWG+DQuV7tyYeZ
lx/QQ09g/jM+xVz6AFYXORoNJUjPB6KucxHmWeqKCmpdI7wswrnjqp+WEfb84F3u
7oaJaevwprlovLUcRLhoVc7Jko+7XIkfCInLqEVNAOPQpgHJK1vcsrfiqMV4AXiW
bIH6LXPtE7Po+s0kP38zNfAe06J+XFC68kyJZv8G5vCeYnuzqJTgrXOLsu5qzl1i
zSYEL9VDnlVW6RP9tbci9b+iDaTlfmSZEfCB2mYzvrKLFo9xhX+dj/4Wl7fvrNtv
JzlMo7qMhJvAKR0/lPmZt0zBaWezNs/3hgWznOg/g6n+wZW5SbHWsL6GOgv5rlVf
ONpJOtD7rED/L5IpjDCHLClLirOUFednH5Mqs5YzEVxbcF3wFmnbRhRwXQ+S5J6k
Dc8SBfK4j9nRpkRE1vN8AUmPcSAlOQ6e+UWbr6cfmZw4RElxmOwVr2XYWjdv9Ndx
jteCypRxia7QKN8tR6mAeKGB9vOKG6Tj/64khDFFMityG8bGvF2k2qklbmTcDEbf
5UPPOSTU51Fx+auZt58Z0tGNPRPP4ZQZ3kxjWifgfMafTjCwHn5HdGNAZboIOrB7
466UXSnjuZT1re78IGKyBq1kOsVZu6meCG8KNDjpTqp3Re3ov2Uo9wVbbAvb9XYQ
EooKlZijCkBcE1mbQG0U6B+oQf4mK6wRWUrJ0W0C4MwqUVelDZEut38aQ3jGxm25
sFwvnO5VceRwE91tJp5/VUJxEnVpEz8sgkjykbEF7K7QHhlcy0l7yqQlO3y+JiZn
j+iLL49rPXT+sEqh3/m7vTMI0UJkmJqCNwknDgbbMkyryA2cNzLwhfUyov3N7Mar
isOeXoVrmOjTX0qCyS6IVYSBrti6DePeeBwidmwjJDeCduBA1Z/nBZ4XNg+jw5Ug
VnxMmNJLxRYjd4aaARVctBXC+AQdD6yrDJSgZ0u/P0RbdHaCD5PahF/XG/8XZJdS
3vwjGxLU0c9lezo0O4Dw55hx6xt88wxuAhgNdgbjvi3npgip8QjezIdnImpN1gmf
IgzuPTEhQlSuop8Ch/IvUyeJbT3+B0JrgDCMXRI2+PMLElCsy8U/UJEw9yBtsgHo
9iibm4lLqF/T3iZ/0WpkYia1s/zSTv/Wb6kmyyOiRX33TInL8Ecp9bAryeJlQR+0
Ff7UhHfiqP28LoB5PAqXwI4+xOLB/ByPkfRri84XgEq6/fEkieU+jekJDxnJzePd
6FkaInh5DCAHMemUIbYtZuGRzE9bg4a8u67OuZyOZ9nQwP4AbGqgnZtVWbrua95J
PNBwih+O4WeeCpMYFJUcHdBcMqO76FRyi73JoCt/PPp/+q/LfzKGxCKlcAF2E1Ku
/Ba2J+l/NhJpbK9qyQgSXDFdXJtP8HhAWj70wMT5BBly586pvKtC1IHRFh5cooCM
6cCSidEKBurrmxBjuiZyrIXWtkH/g3VaGwYVRIFZKxsC7umjCu1v/q54Cecjyq6R
NkE9EIdJYKVxbjqU7aaogPYS5aTc9TuxA4XnBZfg6rFdp4nF8LGR3aQoMTeaOAJq
p4kNn0Zb8FycVeJUClzM9PGLCWPt5r7t4JmzIF04G8szAoTtdj7eB3IQhFv+iYQ4
f1joEOrgL8y3lCQUEofT2CINELCMLiJs1G4GJ4YO5ic8d2NxEQzjtJd664NKMOp9
g+yVZcfaqqdChfwDyrE1nSHFpXe6qtI/dq4ghN/4fHvNIRwdDH8tLbJ/J2VrDAVl
WgivgTs449YpnznY1IsH0lav0X4n827zOot8z3V1iGvtsDHFwu1/EfJPPF0BNj02
kY7Kco/zLFkQg7dicMkthUtXt0UL+9KBdvVM9gqZs6yYxx6xTbMy8KMwMqpFuffi
/Lb6FrvesZ9r8k2Gql4AUCX5ukbH3DFtVHbRvm6mN5rT2PqpUCYROUxbugNHooP7
uUh7eysAND4Skg5BxrQ5TcKLNcko/ml2CKVaF0cOiQy9av5MvfMKtjL3p3bx9Inr
OoTEMd9qzYsZuzQsdS1CYDZ8LxR52/0k6rNQpGB3jevdjNIPuJxUDpgSDgXBmq4A
2hXz1slcPqF6XPG9tYh6+mI0Pe5HqpsTUHoO4Ijosm8h/JzfYtdDXE0x8jbH6YeI
Iq+kf8bvTCSt/+7jzgRmdEzs10w0oBWZvGoDwwLLjk+L1cEGGId6MaHtqBCKuwgr
AQXXSlJ4R1aV1MY4GIlv99EdWp2KMOTaiP30rAGdsz2eCwNvennZadn28kQsMNTj
XFZkYzNuH4j/zZNf/1UVxUYdOgzchQeNsnag+0nZHRYvPRcIKdpRej3+R5M8FpgJ
ugsinyAKMKYMdYtKNZLs9lVCYzKJ9x9Q7shxSCZNEa+en5oA9m5l4v2Kari7QjUA
PB5nq4NuImR9KBvhCJOlyHFqff0RvqQZr1w+m5UGzg21Kai8PycoYzpx2ztq1JHl
lfmf4NGixs3YC/KNewpiMITHACl/PGKXOgVpfEareDOqnfAgANIywMBIqSAVVgAw
wjYBPP5LfjZlnFFWFkoNH+1Pt+Gf/nUSH9hd8y0mCZErUp3GtHGf9/r4REV7kGel
OB7/pxZDMJOBwrPL07JelGyvE2QURXkEQ0bfhX0fUkTyA36hMkAE7YRshmnhPIfe
/O/+ZmNo6vJLfWFoCI6LiWbcsmBWPI/JPvd65Gqq0/+RtrGybpzE20xPkgfahRgd
65YEpYsgrps6px0HslyQXcO6BAXZnhjBVfooESBSIzdi350pE7OtgT/v+s4MrDVu
/2PXiz+klfodqhIDc0XYLYMQVrN2MnbFPLuYvAQyy1TOYKXIoXPNPBvWNr8S1O0s
Zc+HFCGiK5ct1jT5MMZW+BQUSsQdekrIK8c5Qhgg00pGLLJoFazI3uIeYf++4La2
lymllxG67ZvzVkZP0MsBvBn5vSk4181tG3c6d1CdUrDLiqPeSTNw1b3xFHuDys4A
nWsMq5y96bNAPU0+KeusxN2krNzCR9eiD6hLLPoiDvVeynhJQfDLZy0SIFBytJYV
DJ7WNcewoR6nOFScfJ2horvBYGDue7DU1MsgRVJ2xLscj/nk1X9oGYSbyXyqmzjV
Q0Dzf65XOCA5x1dtiRZ7wsC/QezLg2Z6hgFYvUvV22CUdjszHyD6vDw4Avv336kO
9CQZeEpQFlKzPG7yJGxGMCFmh647zcPoqU08HkHgekdmUEvUI8dj73pRlbh/mVIc
JnoUFweNfdYMpXQiaxylgm+WseFZtcwL4Wkc9Mh9BrGkeZjHfUao9yKf9o2i6tju
x78iDw9bq3I+GbkigWtan1+rJgd1Q0mb9Ke7mGP/mjyVUlcFj1jicU6damTlmMZ1
ufe7bvG+KMshj0GBBX5//4WwXwi14bk0T+mpykz+H27GoyDrk9rvggIxHTI+Qmor
BZ64Hc/GSIWJke0JVbijKAj5WRaqDq5AdaXB/ESBuVcEScs7/QC5amVR9WUfvDpO
11lnUFeJASXGQUp9rSxCD7ZqDorN7qIV8+YJdv9Hgubs5ogC6SZFZ8PTFEwgQ/j3
Nf13FxQyui9G7Cc6SmVMm7dDvUgMGHEtVIhnfTNyCUvAZu2yXDt8jIAG2Ays8ulb
gWWHndQESjI81J/tXY9Vq18tA8+oLx4PUtLvxkiuFFUtrU35JWyp13IADfl4R1W1
CWfc4mW8+R8OYkAHq5LVZ6aknc9WhQUCwy3HOouZZs0xawwQhgSQtezcZkibKdvP
Snh9O1fSTsbDog7rlO4rbi3Ji3Nv+1i4yMy05GV+Pl5S8ZY9WTT+l/MTdPiG69h9
r42ll39p4C700UIqBou0hBXHgA8PDJKQDe8iu1v+05KHhswbfPlxLyIFs7CjLnhK
kw/P7BJcyaSzOjICB92eYc4PmBKohOV5OU31C9IwAcKVo++rGcfBqMa36Y4RC9Ib
32YnIFVLruZ7vUJAWykRafIy70fNNk4lamPXvg6IgDNVLSWsF+tArqGGRZ14HNhb
hZy3dbfdXvInuv/ci2rXjJC8Vr2x2FgrOJ6m7pOETSKzCuYdXXSafkUibaTZJIdU
AwR0i2IfR0HkvaLdl/YelerxQlu36K2Z8jHI24ByBItZ4sd3dWHy8SYlrtcThdbo
OH6wsar3E2Jm1quTzCo7lC2GUJRzSbpHLv5Gq2Pl04Tv5fn2S/OshMM70Qdtf7L6
qmzXeVwiqUdQbc1l2A7z2VSKWjgLYPSfQJHfXSUQ6ERThd+qiMqI3HvgX1YuFbpU
4qI3XU0Mxr9L07q6pPhv7tqXgKCZ4jQb/NI6Dc7+3Dzj5eZtXUm2sYKtK0EGN8mk
KC6+tjtHZ3C+q1KVHXPuTLut7FdIDyC7CejAVdfYd6C1kLcYVBPwSqQ4P8FTBV+4
QnpQulWqVa6ocbumUQ7PTa3fIDkYMuCuIX1njB2NIziKsRc21zWU8Ab7gRZI2fwC
cAPccDK9HS/vSYKEf4XQLZ+xlMWxCeuWDjl9NhCCXxUqmg++r1V0ELKnlG4+VyP6
VrU8CPXTCON9LegHPgc0wNNXYLdIUJxr3sUZ2pyFcq0G35n2aSgmMu1NADmtwKCw
2yOMSLDy1Hd+vGkmccsS8Piu8wTMmIEvg8a8CXhmWYQcf6gniNqrYx2vTf7K7dY3
tELV1RVeCpc3qb0S6F/B+7Zv00yuaKZgldKZzZiYTDIeNYu9N8zjzxWbLy2+qFuZ
fOssncsXlN/jlbxaEck6R59xSLmlodWjSL81r6LjB8JCJ6m7YPH+dEoNaVoyZi9J
YdgJQRbi6rEX4FaY0WLHo9KJdeghwfQqgX4GSWBqQcyGUIosYQoCiHxav4fTCwdg
QewMaUTfvGdZy06iaBObjj8/uJetIAazAWQCDKzCwadvhvqQJrIZ+h6dO10NaRtn
+FPXC/x6Ky/SEhJk7FBGoi2b32tEYBRZl5Xbkhp39aLP+rhd54qJgoYsQ9cXjzx+
lvH+Dl0TYiE8IDb9edvgQ9dN7HMX5x4fRCvwYJaGmKnoGjdAbh7BVEX7UYCQx+TP
40OiwvBjMdKwNy+2LmcIEaTkDCVCb0wrdL+i8PjGbXexXV8Tl30LLj/TIN1bxKNc
2zMDWXfOlKDgabiLALwQE7xM0K6wNKKF8EO6xpnaM9fSq9FRrZicVkuONvAqO2Ue
kdxmZjNPI7uArieTu6rpQNAmDRZWkio3+//VWhgmEqw0tU1K+ZnrWaTBA3cNKTx3
PtfwyY7Vz0XVoT7jKXVnk2knsVFsW+tr7mrxd2r7NaVMInJ8vCqAl9ZmFSNTd9Dm
4f1Sv29Qq5gEaV0A1WJmmsHsKvR92fU9DCmrYsLVzisXtEaiOM6tJictSU6XqREj
PTY2AAH7xEJ50nI6LIMp/m+1pgGb2lgjX3qUDhHup6lsiMk7wbvao0cGuqMsViSU
qaE5rcfBy+F/wnKswdh9z1u+TLvWpNxbTJ7kJjBj1EzEE6SmDpUuaY9OrpYr7zhU
A5TbPFvoHOazpqARvbSFyOjSzIWo4yEIySCK49hPc9Ka8s3vAwwwB/MLZM/5MaZw
oJzxsnFOEidVMKqd1Dbaks9uhgPbj4vtT55Jl1TY1Yt1gCPGCkuRWU81m4GKHJwc
zRwmM0OriIy5T3PvRZvghAQEH8CqzqXBjxfJTrOJ7mArfMRKDN0gp8kHlO3VyvNB
DfY4dUg6qJxw82mJdEy3IraZPldxOMQau097aoUAz6SNfldCIC83wmKDQsFkYfix
TePhx6OvkP6rYlwNBkR/8w8lQum4QOuNLIzorFxkkScVQasF2vEf97lPxx0R8Xja
mqcPQe4I6a9bjMeD7A/5OeNcMOF9xBfcSdWjlftlYawmNTwwjABOI4J/i7AWFrRl
6AM3sYri5uThkA9iChu9CTtjm6Kx/6lhXmSgKl3pcbRLFohdgHmkxIfKWM7slcQw
RkuBNCwr2siZDclYPWMVk/yTm1krANZV/cQxJkNawe8cxanqj2JfsW2evkRlbt/r
N/jDCXBVxIK1kC/4AF7HG4syA+Wrhb7nYucXk+aH4a6/hgOlmz7+OfJfy4V1/upZ
eEuD31+lmrhuZ+3v6axNXROnv/i8w7RxbeaLHWeKcg95hAlm/D56cLzJ2AdApnT9
jB/sP9zVM/Br11IVwvQeYcpgdx32bq7UyGqabGOE1YHAGefHxKBLrpJ092/c6jEF
J7LJ4uuffrAwn2pB8J23TpHxFiyuuVm6z2p2hZsl/GRW5yXJlLY/TN/l2xEBPsVN
xfgbhE6RgjWotrhS/8frg9U/bTykBFrWUb3IDpjpNUe1+iNZrf9WMGDHMVYaa05G
ibcS1Van+ZV4IVtIV+bUCPHTPsUxJLZxJjzfV4H+p0ogTJljr0sv1atlOoMHlrhb
1uduc3rGXcTtP8qfin/Kvwp1xA36pJuj++g82qCqMC5/K2R0pc3QDCutydpgY66Z
CqyDz/xu+AQpM5vVQEjia4/WL/SA09iI1CoBHEceZQJnwMWdtVngbLV6GPJDGIPL
UxPXyRNS0K5tyjlq4/cNA2AzLL4bT7C/T6a/EEnTEhKHP9JdRfcME2hU4mK4Wriu
vqTt+BiIWB93UVgiY7eotzOgQIOmVO/KRT7xiCV650XW3BX9ZLa+lDfhPKCvBfRH
dvZQQqZzXCzZrff5/JFAFE+DBL96v5933lklfnell7jIVo16DT894Kh7Q4N4I4QX
IdWTdKzPcIE4Qbgj1CzQ7zzWKuWcziMrpLfrvj3Z4qA+Wft4YypDWu7iWHAQJ9XO
lwPEYIN121Fi5As9YDc7grvB+8x04wHgp65t4rtZhcUa2THQf38/UmpEJ7+HRlhW
TIJMhwY6xtRAf6sxkPGrTADBdHxOIC6j4g2p/509gKlrptCJlpu0avJUM33dR5z6
MhlTOo6HuQdyM/VlY04KfgkOjcc+hOjPeAPptl7vigm0YlmI0/zwdmzKP1A2IvRW
OCMf+iqN/3BH4ms46vB0HEywivwLl6zjm9D1omJdXq5XB1+oqq8wKZEv+LMzeyO5
cr8x/ej8SkOROr3ZbVNeqKtJK9+1he03Wj9522DlYvzL2DMs1q5pZwEde198/Df1
g2WVxV6P7/0lK90WUnLZksj0wqctTp/lLIe2rPnYX2nMNLjoDSYHGhx53QZ+OU0j
x9p3u4L8pobmwscJcHgy1gK3eN4X5djpa8atmTZvMsJrAvIvR4n4Qy653eY9fNcd
773HdOUPL8ojzXrtYWMaI01nYNOHApK1G/5OlFS8OCYCJoGiQ98/QdiTsZdfGtQ2
BXUuSAqrlAJGkqJbyE1UUYgoCFkygbU6jzm5J5nPX5VVWGr+HblwDHe3HCEVPdmZ
FLnpsg7obZrppBwQYvCe41AyEOumi4ASRu0nJIt4xTFyGM/hcSyF8EoQospkloR8
ACqzJPGM6XKuNGL/25pTKdO24f+d46/ETvsOvnePAUKnNYR4PXWnvqREoFz0Rq3A
V063WoF7l8weet3ekp2861fu6TPbIe042PrIIGxwd3K0Pcpdh57dxtGj2eWdLepT
pMaqi3i9E5avjQmLFYAu/lju+bZb15Qr3Fj4+e+NhF3GuKCAT4HCBzEPvFx6rdxX
KUARJUCAJvNn4MvhC7lJl9tUuuAMKmV6dBx5UV3TMUupSRrWGmAbNjRJ66UuECh6
CAY31OsMS4ZVDsK+cFIEJiNBz/nzZ10wKcHSHBqtbVyU1qr3k6KVkaFJr0QGeY5b
4acydIZ1ueE6agIocLHvNLmOigAjJ/8BbEknmln1qdSP+yn+wYx1YPPS06qY2ApO
gIcQuFmEcpGuIEhueNN2hYYkkxQ4wfFXBgp4U5hUIsD9iE346SVmkhtB7SSV1ohx
lmfyTSDN78MY+R2yVVAlEjqnB8O3ckAManbwbCI1H1JIVMl92NzZpod+1LkAGMEP
FDGqTL03ix0X4ees0a13v9zGV9emIRfmd8WCYPJ4LVVYULJFfogE3R0FDp8KgfyA
uhO0ZvzKIIhIAT8xP628yQVSc1tL1ewYURLWLcq/PtT0BF9pGz9ImlNiCwbUUjp1
fgV3CP8hs0qXxiMiYogIwr/pwT4YA2dTJYh6CfdgICkc8SZuml5LZR2XcbsXPQ3Y
4Phs8Z8/NIvy9ljsoCCvG37FQM5nMUY/+2LLlevyIfID89+LFL0dYq3B/+dwo7dv
t/24bHd3SexXUOwg9+R1EBqTQJHBkbLuNPbXWPvu+zLXNzZ1YP2t8465D47fbvVk
8B4UO//kP3tNZhzkWHnU0paK6aP3XCIq0s+Bf64ClIMwO9V5bwrZlYcP/CE7r+VD
fRDVytkWLsINM2YDrf7T/kgXRFWfVyNDyuNosVO10SyZwH+cLg3HMP9bUutf3GvC
PdC3NprQsa1U5BddLy/x0xKFYp0nzHdNZaCEeldxeEXyZtLfR1318mI/Re7xhz/m
uCDyPFbmx55qXgmcUxwIlwCNjfY14smmQuRIO2eJJv9Rfloa3AYnTqZ0pKvNv9oL
0HY8NDiXb/Ayk05oDAFEofhDcWhLHfe4OKho/jBMfzMyzjrCsrYIZRqhYWst4AQA
Olt9bwSKpH1/xTZ7p719No9+vibaKuT7YkRBIcbXivPGGytf0AC234QlZXAPWWnD
fwtYh5Pz/iG6a4W/I7pxpX0/82OHSHDdA+ZFKJUp64hiHPAwQ8rJ9jXtE/kubYby
3Q+uywkMfNvTL4GbKxGxvnYM2jL6rEoiHxNy7hYNwaunWGBrJ00LqgSRlSUtfHW4
8H+VzwROKxzzYRyqzZC55O3pohTls/WJkO+qPtoxMewuSnDFVh50PNFuV8C+IfVf
uQd/R2xEf34ZvWO1CPpqoJo2ax+1Xc3x3Wf0EpYbBThRsUUuullqupqp3wxJW0zc
qIhZ6iVTUmHBQtq8CIog/pn+DSEjOqfkblWoScxVGb1GDdgqQZfDaoFEY6/Irv2J
FNj+vmjTIQ6Vq3+Al+311OI8xUCdAy1nT9JiyDC8BfGqHW2JiZidpdozmw8K1a/G
+Sjt0FgtYVU7U+7klpGZ6hXA6vObXzpW2BgroK11c8cKA1BalHwfnO0DS0Q/UfgQ
i3dp68mB5hg61twdo+W3N4e9rf7Uksb7eSWwfwfk2j/BYbHf2GaOPJJMP0f/WGD6
/rWgeeOi45tIaILfAMVFQgyVoinF5LTeho6dER5ZtfID8QENs6SQv7jyNjKGM9K0
NNUn5nZDxSbV6MPAOCciTheAI2FP6o3BWBVnKgpV+tzgysFhRaQhTZMvqpzu0YLP
ol4gyofk/EUdNPjrpLH5TcrwRHs0p29XWPhJRYkH4skgV3YN3Ws8vewsJ2zjDrZn
hWX8jzzi3nKrJd+4cZ29SUyPWij1Qpmyk86XCtCl/iooyGNey2KhasLICzW6Qs0N
7Nj5aK5wjejY1ZkFkx+yO0GLzv10/smgmFrm4bflh4aB3xf0lQCzglS1TQbRY5Or
bvU9JIT8xGgwd5rv7syecOE8otiWiBGsf7gl6KtrfbYhQVoeOVlbHNIbd0SFaZEQ
9BzFAMvhxFVtR4kpxAZI8orHPsHtIVqJNXxSp5FPLoRX5vLQPEYTvQycL9Uhcrkx
jdOB+FNloxh3lDcazhYqfYm2Qx84UIjppbQQj2NqGcN5KS9wRTccn8fmGjtWEaQd
XmHcQJTQ3CKJH9rEyjUqb1itIFYAPEqecd5anAv4PK5nE9ifu8aJ/iJizMgPsYwM
T7KtyNPJD/NPnCenbBvAub8YhoutMu6iAUQkgFEVSAagKorSzlCDbFafuR1sMZB3
UFV5oBeaNz94hm97rYYBAwqFubOYFr+KDttCv1Z5IiaYkAz1A1BYwp5/PbbBEb8C
vhL054x/huhKKeUAJG9zbg==
`protect END_PROTECTED
