`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
112vmU+Ui+NiwBWprHiw9jWV8YBujDr1TsyKEeYPe2sYUvjT3gdHuBA8BkgEsoRN
uho77n/yp5601YjU7f1JUfG1691WkJY6cyGZSvSKIinQKfXbdMxKmtNcC80z7yWQ
oB74H9n1AuokdggFm9IUMxwtW7DhF6675uI9VrfE2Agv8bqOJe2DbICGFunFvgjY
f4GRsrBA27kGpt53UV1NV+5bh5t7DsJzX412sVaqKszdC7DAcVj8kvyihwkjFvD8
gPqp7+WzXW4RZ2pzV6n6ocdM9d2m2eXOnAxlnPrNFYYmJahBIXIZ6SuYLuWUrIi2
gUjU43bXDBi9svkxMlmCEka9TofYhnNxsz+y3mWsFC8eZg7bD15HnPzMZYW8QH0D
r8Q+dlnq3SIL7LRy6g/orCJKhqO4L/cUbwdW89FNNlvvZdNqcp2g0VKuGaddOA8Q
iV5CzYpVrNS8qVrctt+cgbfg5vntUJJPi8eUPReklylcSblsu6Uqbf26N59cNF7A
rEpcvoxUBz6Ooxqnlj3SVGYU8nSjJAAZ8MSnCx9Hj5VpS0c/BUoxCX32VKdGXbFR
px/OvoGCgANIWMGg6A1QZWA7V0l1w2P4JDUdPTiriYg=
`protect END_PROTECTED
