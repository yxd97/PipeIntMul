`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zvmc6Sas0BGWE4bGF6ztrtms91PqkZPoxkl2GCrPrYa2dkW1mjLyn+Zbli4VQCX
gshmDL6YiZFjZh7jHoUgvwGJ8NnSKCUlNVmboljM2k65+va0mhGPpSdzNudsI8Zq
ji4a2nYyECGl1DZGOyZus203TelPgcDbesTGTQW9g+I9wdFDnt+XhSlEE87LbRIe
vlEZsZ8EpEKo8t5CHc0UTZj6znJNNtlGeYUpNgpyxcvbUg3DTBfM4Hv++f8WFpdo
CM9U1bBK4SNJFOispYNa9X9jG/Q7ZtmJtwqtk+1rWed0D3h808/BWUO2qY+FwUfs
O93K8s8P24JRLVam6ut0bS6/oxGlwpXjBOpF0NM2vG5i6UQd++7bP1x8brQYLGbs
55k4wt5+fl7S3Evy7ThaHW+L376LkaTSwc8OgbP9Ilk=
`protect END_PROTECTED
