`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eITEPlMFjtAczQFvUGS16sGSGybPUwDU4Ks1kwXPF7syYZQDhAnjz704XX2Mtadg
dVldrMWaSyl9ujThKSsmTsODNhO/fpeDaX3OxbhuuSFPbCzLKPo/S/klfSNL82nc
YKVXns2pxXMhP3wWe3SibLrP+vNplKw0RehQsq4K2x5ZXR0Ibp4tjKzmp3dYEYcu
40ZA65INhadBV41fCIUK6XP7p44TLujZsavqIWPIAAPo2BGzLZWH1AxwUuxxjEfj
p9Xa3wJ61yzf3M/tt4YmlRIobgzHi9ZaLH0f6qoyaLxIBFdaTLT1CS1CT0J5ezwO
VvCshVjqYgHXgvjzcwTcXg==
`protect END_PROTECTED
