`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xdhKGvihBzOb33vgw8lDjwAYJpdLGpa6lvofArg9Znx0Vnso6PaD7ZpL4fUWrK0I
AmeBhgU/bH5V+4O+nJdoJKN7GplpmW7JoT6mkWxefXS6M0xOJ4rYj1Wt8f3x4iE8
CBFVWLRhJqWZAUl1eRYRIizYeIrbqVmSzN/9UrKzEG+yMc1zr/IZcNPTIEpWV2As
tHlSrCCfimbd/UnkbMbOOj9tcM2YESpRHBALDEHrgIwOhy2JQVx3DUoO1+ryGYf2
52PG4UgF0QcKe6M/Dh8MyGc60jtO5w6vAv6NDDNYGrPfs1PU0ZKr7UDkfpedJJnY
5s/bZxz3NOu6cB2vipeTKzwbQv/df8eR2Vxk5usQtJ/WXfGGctJSsIZMk4qxrikM
D5SXNIi6bH3MnNYTg1UyiYO+CUHTC1R7iMmy4iO2WYCi92uRSepFbrp/oy45IGjx
eSY6wILvPtQOtbQ+HBIvy1ICPiDZdKVKHTo/t40DbubWi+chELgT3dZ7FA1HOcs3
j2iyjPOPOh9X0VriEmfi8sG6i5dAqWDCtAiOzdcTblGag3e5Ux3Xwu0fs2VNxWoW
avcFOO8684+4wuWWAf2ACHC1ZI5HvlNddk+EgpuFNz4pSZSplkvVYdqmJZAqWXPC
YFEmtgPckl2BwSos/446K4BYAFTjX/b0mu915QchLodEoCXiifbP9bS3LanLOM/y
VxA7in8fko74dkiDdTkdeA==
`protect END_PROTECTED
