`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nAZn3QfS2t0YN433/UIohquPR+DJsc1r97cQGzLMRXVNuJWGH+6VEewU4hdhysvk
t4UTVWirUdCDf3mRXc+DyC4JCzOOlgm322wRO+juvmg8GnGdYnHhiGJeTXnZYQ6N
9IsLssxDH+zZy3zAqV6Jf72eqEii1BxWSg9KeqGioKBCK7hIXF4NgNYQQiNBOvfQ
XjG/WZHhaeBJSaePwz26bqTS7HtTK1r6FRbaYsvQB3CWpFwrG0ScPm5A1hbqRr4K
125Ud2K3xkgyX6f4BIT5fuLqdXA9A42mG+HyqZ6pwoupFnR1vWqUK2AFOE4Vzrq7
t9BD3rxV0oRPAaWELfP9sou+eI0itpIJDdHYuk37to0iJCgr/LsCgjiTRblx44gV
`protect END_PROTECTED
