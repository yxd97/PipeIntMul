`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yLw5N3dXqKAfyJTeG4lnHIAIL76C4UO2R2foBKC9xv+/wQi0p7bQPq0SmHgN1yv
gOLK5yboqTmjdPmpGq2BghxOea45CuyR2qADRsdL5BeqLydy4UD+hTZ3Euj5OG3x
kt8iBi/I3BYvzKMbb0scdHHmxIShsIdr3AjiasJWMVJXaGT/NFgHO8BH7fw4ENRp
uMRgY4sB22zQbl5q2LUia8s8Png887x3P9wwlyRMaFMUsnRP71X5M9ous+8kLER7
LoSojqAYZMUqq7lIARRr1W8jy7GsjpfvwQFi+UerJZ0P21FxoiwlAmbQ/ogv+tQI
XylHbomjUM2r53oC15Y6A9or4D0Lqd5oq3Y6Uqx+tN4WwVLjZ297zvxD0k/sOotB
rzMdlqRPqZkM5AWg8Weqg+11Q74N2s0pANbd8UmSBnDX5gHhY3LP5DFvE0cKRmeI
Ay3+TVpSKE9B8n4yo6wqB5Lz0i6QGh/zbiBDWCEOINgzHZt6Se9xRes7Y1zefiQT
M/Mu4YM4vt5CpJJVDgvxsCUZqY6Pm4pKfVtf6M4nd7qIudu9vjid0d2bhfblqXKL
rqVZQh7HAdV2813GpA8JOA==
`protect END_PROTECTED
