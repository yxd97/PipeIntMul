`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yfUYlUt6xcYpT+33MxUli5Mf/TnjyiqyodZ7M/H7KUf43eMKqxXZgqyUMp6ZqGVZ
HH1zTciVR5YviShnQNtAA2UqpnXk8D6pDvum/Mql50UQpDc/N6rWsilPsCATQlUY
SlgmOxjgmV7+UDbi6DHF8IcL6tM7p1Xd3yYOwfWuYa50Zqd3xOP3WmKW3MgedNep
Sr38sB6zOhPtRzzlUFiyYxOt8xn5m9fjVx+jqfgLAD0QU0IT/R19AHkybCzHnVON
/t+93tV/xOPJmrbC1cYTHGqfEQrag2DGych1J/hEpbLSW3ITFUoTexvaH+l/NSL2
a9XZEURG9yykQYhWH+M3ivXCglmZ0SgYatKK5E38P57+ypFx5nr7TLiMYNR5Xlko
`protect END_PROTECTED
