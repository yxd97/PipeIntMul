`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PqWo5MKyQvPY2LZVfN4bn2xoGvxUnO7JWM2ofnjf3f1yZwncAnY9UUd2q4oLSfLA
2yzVenF1OsI9lW/fi4cq0N13c+RhUz5/Yy8aIB4BlVagJy8gFRfw4XEzbAcqMHt7
vAbKCQXXFmQ3gRjcKT/tOaygGEKQp2VZXcBsJdeLpQCePyg6Y3YCRZI82Blt3uTi
+eBzXm7hvWe6IxymNtg28a0UnVBcZ1+dA+TKZPe8sRk1fkl9QhYidk5fYtDmk253
5/H7dGnuYtfAsNtjQ10/EvjQN5KGk2N7/jr5Nmoss7oUcb50VDnZdKoorEyY0EAR
zQywvNDruhJ4dzPeW2/tqd23VYF0azuQoD9B3i0ZlTfIyykQf7TW8KYy65+lqZwq
2webktl0au6gwGDzWusv7PfqTXdM/CCKlzGhRyLRNrbywi7jk/O3FqKUouSrrF14
`protect END_PROTECTED
