`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZweH9qCCP3up0Ksr8BV0OlR4SBGti4AsBaTYcOCJCuMakxUH1ELm07Rm0XXmEW2w
8mgejDzwcu6EB1HunPYTNohSb9sT/8d8CkafyyY6y4PTgnuJSF/rA0Vc+L4f+hWZ
tTicCZexDfA67Z7JcTaPS1xgGzvvAlMEnu3bjwXRsV2HnjYIkajQfzVobpjlktEv
PedzdIT2ECfIBZk3eGjgFWwQxB36Gc1QL3rJpoyhiX+nKHoH5Hj/8rGbj302l6lA
LhGy9mjmWwEr6nOjUHuy7C5QZQd1hZNdQ5Cxhm+nJegaOi1ru9X8M7maWvIrIqGI
HMh9WT70mHeCR3IqJgRNPvZfjLEmiomtaLQMQPQbDw/WS/21svDDVp9hQFiJtHTE
Xq2s9VKNGHskBLugH3N3WszfQo95u1ZODMDzA54qA3SIkdKTFdHpLm04DbPV04ep
Cw1dPE2rVtmMV9q2DIZPzCN9uOJ0yjtpw04928IE11gK33rOqzDTbDGzReo0LXOK
OMK/HkkXEZRTcHm+6BemOHgjHxx6kbcGniEq0Asx7ymul74ze6v9XQCU8MDRgWOA
qDiOARREBlg1YGZQbrrTYPvnbKD2k+UWuXE/2mzvp+94O7JMalNcmu52dHd4vhBm
m+vO53gmwRMTSssB+1LlplirKQ6Tca12fvODFtkKsUdjMPTD8icugNU6BPAooSpN
wCrgutWceU51PSvYMElUuzRMeSZwhb3mHaJ2x2ComW+6abHXmaymC6RflkOwM2sZ
wXRP6syTlhU4qe7Ak1XMiGEPYPAEFuXRsb+FoNBeygS0FyvK8/e4KiXhEAtkrQ7f
RrLLWkGlcxHeU0arzc/raRfMUVYSVQFpUECDIkkoyFjCyz0S8OJYVwEu10JjS26c
5+DaWFa+BiaiV58ngzlNEz+E9cczGi0abixXA1vvkk3P04wMruqocXG0WLDBm0MJ
4WdS7jlWB3W2jEWzD+xlg/SGIz0jjMuNxL7dURRue5EyhEYf0pP1zjdYyP+VwFmm
`protect END_PROTECTED
