`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HVXRdYhhJ2ltXyM72DRGoKaizUbivvCEVesFFr+qIlQOD8htqLsTsUXeWG8zKxt6
60QkWQtn6HfbzfpE0hF9XgKp9QSXK9u30hAlJbcHUTNpXYgd5xVCWeEx3PXHQFSc
HbG5TuGM8bMFJ64fkPkStU8Nsj4dCI4x+xeOdjnySRr5azz5p3r+FyWBI4uL7NgF
oqPwh258MuBDP/kw3LuA/d8TlPwyMUkQkgqLrttyIITPIPAXqhKA23Mc1hzw5qCv
reF85a+Olx9tLOa2ZypJIrhwH/NAQIik4QH+zYdDJxBKSVZLqBLoTH/r4wMI7f4V
UktV9L/qRyJ4DF4rSTTguyJKBchWc06umc0qMRCQR6/vEm8sx0aNJgw7PPJpAvd5
kpV2tvu12FX8CKKK1JiY5qruj71sFPlWeQUeczzsGBSM2DiaowW6N4vxR3vKXZ9k
aFfo0bH4/SL+V8DDLGqUOJJwvZpMjVUVbYIECdBSW9Skx1tOGE7NMBiEKeHAV4S9
VnWwiSx7pO5tOSLCyhG+5I46bzOFEawQlbZ3y7DEyPpqf1xg0KzHnEFayKLGO1yt
`protect END_PROTECTED
