`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hXqdjILMDHrEDWl32dWCY5JtikAzx7Dd0yxN2FNo0q3KGFVPVaG6/g1kSKiMr87K
5q7qkRoRNW2R26X2Ig6fZSHfiLboIScPO4Nd1sPMPTlmU6I5ahv0WHoD28UtET1y
n8mP/g8mQSNbRxiCzsbUb0t7S/D/Vtzcm/CENNWHm+Rexz6c5n15+zwrty+5P2s0
sfUGAQQO0/dRWRM6GgMCG1vIeBzgMEczslwFz09THHrdvnRJMwRl2nhlD1byt4t2
h0qnbXKBSSg6PXHHfeDN+7pDJAg6FUBBsraWb/zVOrkkOscOXEa+XUG4YF3VlJMb
f20BqZ3c11eHWeCXxMN2Gj5lwJb+XUWmdLNSiPhf99+pNq+hCfaAy0Nd/fypSlRI
km9EmxE+jidcx5B/q1AmOzGKRjSWh3t5GF5jzP629szS83Yp8WZd7SBIhhPg2ZVK
EyZYAomg6bkP0RJtRdSkjTJPm4+lzgqzQQLFWRGHcAmf+CBk92cYvXf2oqsUYH4b
DzPq0eP31DXkc506Gs5D9SB3XVV27rBtJUrdJfHeD49TbLOlHh7aD9QhVTLTy0ve
hHvVJDpDBwfuwqNq0hjTXbzQNBH7UyXb2PEIF9BtGhbR4o2fv2fD6kwWxaElEIHT
gyr5sS/2dPgqGnRhkMLkHhBYQcL7UGdq/4a8WZ/WVEOB0Bjq7XA7FChhYS68cpHf
5xVxCDJ5rrtUCmON68VNNq7UaD+hYK60bwuiDcesG0g+cnZ9r6mElQaFwMZfOcsj
DrAovSL3l1xHrifbo5PwkXhacxZug4NcapqKw/VhObHvWZyUc1vcbsmutaL3rMqR
cMb6Y3zMOzvsGmz+EXqN+taKUNdX0BOrlhyhUQnVsPU9rIRF28raYhZunY+A0Z6k
mhZwR9OgzPwchIUqOqNhLg==
`protect END_PROTECTED
