`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gm+kZj5FkctiiXAw55imPbp1BiMkqiINsWUl0zyLIiCFYlShNg5ajtNlG+/K3Y4t
qAQWtshPomh8dZLpFj25Ku/2b7lQ0+LU90e6p7ovWiTWAulxF+Rih1cFBmhm0/kO
8Or1D8ExQ151/5mPYxKgsyY4fo8uP0QmLPlzAVsfhD/NFxISqTmB/OJizyPPErRR
/eEclluyFsv0wLRXYveqaOf1nsDnrEDT0C/aIv19dJssH5OWfP/ITjKJmZtDUkdC
s3MRDEExB7M9eZKy/CjIww8L7ZTNQjJY/k86/2PZ2rSzmh2f1iAzIw36N7/mNxRQ
lAmyRvgYlKcu0ExbdQ5Fxw2VSBy/Yc8YrvGivSB9mu4BqbI5ZlAfkIYD12VIcDZt
8fOvkM5xPRcx8+HRbzKkdLk8n4vHE+jJ67sMEljZxHi32pm/nokG1l5MRxxPnibS
6zI4Q3FzC0TBOFsaXds1LFgh7w9f4WCeGCNBfElHd5T+Q6UpIxHqvc2F+4cXo+6o
gAevT0gf5D9ySI2ac5O02L2NnCEBIiJEzXWTk/29aMccz3bzCZKJruBAhojlMETE
VqAZfB2B0K+24xMC0rnh41dNm1PgVe3jxj0mjomS0d49rcLG0FsimF0BdAbjHNgx
Zu3kUeD+26ek50L3rFsngpVroKjdJBvkQCTY5+hXbPpDBFdZcv2v44iZ+Oa/m1E3
lhL91IuGYaKImUKsMFHK+FY8q0Mxl4caznF0iA072chzxG3ehd7X8sJp2qpVtzNR
a7heJwot+sXQNQr9OmRubhWOi/ofjtkrYRpteEYXPA4yuYRI57M2FN22g37EN5cp
n8SvdwtYtnhH9hZg+h5YYUO2PSCL/fx2Ifoe2cMNQv9Cbk+4n4ZtCzw/Y2yzXvf6
/aWGnn4Z+tIqpHAuPNqxoRsWdYJz9u3QiZFwHaXEDFBK9Lmp3N1f34PVu1Xzzse4
qssk5zixqn/VJS76K8kU3DH1N5g2wSqkcNn+mTKlUI8x5MHCsyKbaQIe7V0ZD4lW
habJ93xRzXXrcVwDfoJ9RCuWeq0L8H/tSpDMCKY6vnZ10BigTWJmFvnumFiEEKaG
cRcvZfz1t9dYoaXCrz3dbzMcpkXrfV025sGbfcaQW+CHgsTyNJ3Lh2Es6HJCHOPM
NuyXh4R0Klglm/oOHUaCSle0U/c/yO6tQU425o9UTLl26gQd7zI9a2memf4HKE1H
iHFA7XRuu3yXmggw5QQv4ocbV7gU/YKDsIIfgaHTp+e/fSRqkLkeeX4TwIemuQ5K
`protect END_PROTECTED
