`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afae0jX1lFyhSgLpD6bZ2gXHl2s4b0Vb/CvzorLB5wGirLClIxqMnMxN5wwMnwfx
49pq2LQuhk9nBJCWmnXaV1Qz8IS5sO3i2hk79+a9O5p+axA2LWtoKvqDWAxn4SQv
nN7QofvU/vomSYG67GYgq+w0mu30CzK5SiD57obBn4ZigjOYDrBzCDSpHdX3VBTY
xlJjWh/eo7VwdG2/SfSScubBqA0tNfvsF9AxjQESUwmaor9clyQP7c0Pbw7L926o
HZXK1Y8oECme4IG4kCshEzBBxWmcypahBOdaja2S8OkPElCKoylvM8hIGZ7zGUm8
YglE4DKPMoCBJEtuZESorLtCCqwAsofqNFfz7L7zgaheOpBg6SZG/LKjiTooBhrv
04fl5Ew+59rvJjWdUmx1bkNmlyqj/e/LN767AeFNU6wU0a0y/u3KgRF3T6tAycd0
9KETkwNAebt5cX7/8eeghXfEblmHU4rRw8y3M8qPSRkqXnlMCiTF5EF0KKa+lqeY
PHUL2jotObTJiApZBYekp95H1DWbkTu75DfJ7NnQE3co0BUtB1yQCfrS6plSksnP
sYffmuk0IL9Zyp/RznH86whs3v96hfv7IRP2n00jUrxdrX3d3MPMhqFV3c/veNK8
6egmIrl51ZqvEwZKnYY8xozDNpx5jU7KbkTl5WKJ7nDiElSrUqV8pwxiL8imqAPW
Nlom1DQfHMtxHut8xAiJ74yhOtSkMaPr1NQP4G32TRyofgCgbJ6TJHg8zNxwpv2o
XgFmSXfPyUWgMrfRnFm9Ef10jTGqAj8V944A0JLWZSEe3slbJ7MUm1v9elp1II9n
eQcwVC73sFtT3GkhGYzFCO9WlloqUWWOzoKA6Ec+ggoYUEaegYBzJTMS5IuALBmJ
OTKFJ94y61gQfRKBq7nvYIFiKRkl+WMhEcKB15m7O1fSO6RCgpTXhwA9kYn+PM60
kIn1SkP4SnwC8Aicxi/KKdIVy/yCIIyNKyp3+N1Sc+w3+MuAMmHpSLmiv+YStWHw
Y2IGMwvFR7f7SyQ6xTUFaoTW9VI+qaFcs8dd+HLZ7GsTZi+3wDMFPD9Mn4HmuEUu
y4tCmVypV1g05ohvUgmJrgY2pi60PPXIuBi8w1gnrdh37iGXNavEC4llhck85BlT
duNN7jomRcpshJGhMD2lp8aNowj+luG6JEx/qvuA6k6oq2lwZqzpSBU+ZPizBH2n
YVIMxvpqc0fCrL6lku6AZ6g8FuCF0SHVGXLHnlzWYQHtwrS15DrnRr1kKl8UFXAS
AKPz4yODKo5kHeDuNhbr45ru+kLbya/ppCqC6G7CuGAnEu6lS27akoUtQjWvThjl
i69wx/eKxdSwtsaC+QpYY7RejPFqEETrwLm/Bnwx01ZsmB74S6JYul4T21VWU3Lv
uQwoqXYEA6qy0u1xs+V4AdzQPQvX72WhIklmgagMlDXVBXzBGHy8XwAvJXHe8n/F
w3kaw+wCsjRULltiIRixp+U7JNoNu3bJQzJuPFc2O3R4DLmxaB3yTwIOyMe3DWEb
UhixImKgXkBAjNhON+MB+ba35/sDiiHbm4W+iRfoeOCLtRVrSTMYj5b6kWC3wD2n
PjzGHYuO1HBSFWkaCrlah2OeMAfi8fF9RPjoIypkfL/iOMYCE7qvGJmGjLzF1gY5
Z4zdp7Iewy+Tt32E+Bfec4cCoLVQf+9TGFzByvL/g+rxt0/wKXDiIcGkfJZiBVDs
V8Bcsk5HuHCNqiGyQSTzUaB9HL7lhmWrd3167unGK83191X8ggV4LcWrihgqLyR4
bw2F7I+OTgoy+7fjwvDe8BqO04MeIehYivQJUX/qji0McE5nxX2gH9Gol8oWoBjz
X7Zl8K4IzJc2Th42gwyCfo5zQNFUfboCvYskR3cOiKsVvYqYf7rFH9aBwcKXZl/Z
b4YfEu4A3zCplFU8s1LoiJvsTna+UPPTC/zKMaV35FBQAlfZDSAg93Wv400nECle
EPe/XFg/wUJHmKBPR1V6Wll514XMKn1R9932ikXaxMyUhyvC/RCtatIH6vL6SGsc
WKE1xiICjBIVG/kM8SHo/SwJFwC6gbWN3U2ppYc2VlOJpeG8fCKv0wtF99LKvNyH
GHQppgmC/UI88I8tc0AQnYXvDgKhGz6Hixow3XNkYnTRzmXHni9ckjuxQSR7Ssgc
ddPVwYxmp5Dr3KJ/S/ehfplSxrjjdiEPKooXMwA+YVm7iuAOo0rXSJyrQwlmb82L
noBN03aR2t1otLqC7AZzG3QIGMi9dxUUW+cmyfBMsBTGMcbLi0Z/j7Aomph0luIH
aQaaoCptk0BE0I+qn4o33AY3qUyyK3xdouw/xtjmfvh8JJPOEi9iT07m2m8PmvpE
l2UnTPBWqG2jW0t666pdIunL//kwLTfT4gj5KasCPDA=
`protect END_PROTECTED
