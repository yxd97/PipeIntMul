`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xHdSZOIE8/YesObkOSs0x+NcijzduxtGp/ThVs7oRaIYVSA7P0geBBEewjkXljfP
XtiPgn58GzeL6KHe7ipxGtn2kBWFZlkF+dJq9JzuQZ0CzAARPnMn7etdwJtZRjW5
94yaW2udjEqRtHfSUsRCJffxeDyOhy2LkkFrAIQJLcH0iEONNdDC18wDNzRTz4Gk
wRf/YDiteCPn8N75ROVlnYQZ3N9KsaY7BCBTLIHSwy4ORu24ycm+i8htnaAaFptE
UNzWCKm0yEtaWPvIsYxdc5lrYgz/wFK9tn2q7YsgtyNjLbfqpUbhFSjXYboHkk1w
4/UZEtw2fhRZhQ1p+ZzhgeecFwDCPd9FM11nHGeAQl9lu3uk5+cKvJXlf2GU13pn
a5jkgBvYEitJkZCitY8AXM7K6KsGV0iOyeYQQxHQ9PKAF1WkIaC5NMIGqWuyIZJS
fBK9wkjfrqM5cMdE3tpwWInfE9fEn4J3MHENIr2GtPkuc5HN3pBeeob1dbgjh+Sc
FnaQpg7aFbI1Fgiyk0qjNw==
`protect END_PROTECTED
