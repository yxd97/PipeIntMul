`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
szlQHLCtr20ONR9gA8jdgVsxV5RuvnIE1CJ42kvi7/w/IUqKGYISQJxN/Xdm1X4x
a0lm+QDpG+oAtZYDyiuOTcmHKvU5OtbClNkBmuuAWmn6HGYOMsFz68w+S7tB3H+P
pdS7Ylwp0b7tJbKdmSCgk6Vmtv3ryfAKgGk9HXtpJTTDUB2QzeXCp59H31/8PS5w
Gdb/qO82Np2MXlu08dRNo+iontXN8Z6pQiuCxurqBm5CBR73Lr11R/uB96u+lFRV
kTAJTRoC3cCIh6HinrjaKLmlKg/j3/L2wJwUVVYt2XrzMCJvBZvK25vWqxwI4KqG
dywILIanc3IsHzuXYyhOkE9WzmUeuzBSsPs4+M4XIIPyJTYz5UCZYNKMq4unsv6I
ZqZIwV3Bum5coLxUQcc0N/HYhKplmZ8W4X+58Jpg0wyoDuglQwBy//BIPNTbCJau
h9rpJwpFXLGTpwfKVJvfu8Mmd0sFeZt/GDZBricFJWBlwX+QOcOu5yBe9Q4gkOWe
ToBi+30JlI0cVkbY9d4sVSgq/oOknHLtyhlz4MjPpL4=
`protect END_PROTECTED
