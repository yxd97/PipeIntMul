`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
asL7S5iU4DJYF9WdjkakWQsog7esgpoZCZdiRuxcgBjTg4XxkwXnq4fPya123MrP
zINmk1FybGMYs9i4UnRfhGFjRUkd/NmZ97GIpKSGaB8hs5+fc7r2RGS8Yp1T3KNW
1vMS84JiUmovO9kjT+ajcE/LvnN9TUmY3JAYEtF3qmeVjUVWK5P4BL7PyOpeTIQQ
2SuW+qjz4bD2XIwe7FSCsjtPX9IJEQG8E99VXTt8jTM1G6sS2V4USE51BIM0j3s7
hAjgCLHH61dN230llzdRSGFNflVfbE8GLNbRCTjFOS3lphL0UAShS8tEFnVr2I7g
dG4vZL+3pQKDFI0oKcBEiV2D8WXPXuV2EOA5+rtlJMY2lRkiy7pdCfJHkUTSIeYn
uSvdeG42UljAeDIFDrZ4Tt2xPpgnxmFJGiUadZyGEcn8iC0Njhc47MfhT72C740+
ixI/o2Z+lfQyP43sETB+BMbUkCFtBDNhsKmvLynftf75+/QjNJoofFJexmfaI6e0
Y+2FYmHyXTr5/5nVRkAvBIKAoNLQCX9BC3p7cdKbCs7Dt/T9WGLr6j7rVuq2qVXi
/Bbje/uGHyvHWvctxWnVOTqV9H31+bszlfctk6pxwtI=
`protect END_PROTECTED
