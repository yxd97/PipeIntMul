`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gaIrY4dq05H1xin1KKoHOAKDNz88Y5a97pfXrEgc4BeOUAOHIv0dEyRwZZxgcTwy
t0YlkfTrtjJ+j+CEdH19U2Ttjj80FlgeVixdAYnZrJqa1flmATWDZsUGtrXFSafI
GVPATKMLPbQKUrXnFChTdZk6f0KArLL4kEjSelalIHxdOtYWW7ArBEQRO7xU1Jc6
rkQ5vGW2b1gaPKQmhgTRhWDI2U0iomdmvs52a/bejFvtGLbFQqy6TqltM7UzFY6G
jX4yG6LYaHMu5Kz7gbQspVC+XWt1+M+EoEA4I8Z3G6YBw+q5pnihC7DcOKk4kjBb
K36i9pIOWPvX/WhUJ/A/MqHw0a7nAZ8E7N+1MRotUt+U7EaQ185IUxhJZNgW9qbL
nIwPOg2BnpZ8SDsXRU0JDofQaC2eOliiV2Vuu3so5euRm/jw5lJXHdQFEec4w4sg
R8et0aNF9A5BIXexc5JyYdnlxFpmlF03fYP8T46QzVxe9HYZDTn6WABcwDxujsHx
`protect END_PROTECTED
