`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FDrhv+fb6tVPfZDr6WX9M8KL5cCiUM8HxP66FVux9bwlWp2B3G7YMkse+10tF2SL
DDGh4pVR+gdDk1Z9Cg51xYwHJ6iPVC4Q6j2ZxvJGJu7ZqmOgaD9Qt6DXE6M+IAqL
6cnXMT0sKxiGWna4lsj7XYBT1MaqKIk1gNyY5NQisa5DToUdvrdDNFzhB0SZR82f
/15w8nBLospq94PYeXydcdi3qLsCTJfwoed9998m1Yf9x2aehkKXDH4u+l5Mj1im
ptU8T4isXxWnfkruYYqkCfrDxnvUUGkBVyG7g0eu+r8y6dhqgnTInEib/Ki8+wnI
Bdg1ApF2VnhUMMmzX2J45tC3kLEwsSmFXMCrKjFc68dPgvmWhXBlsiS3/seHozan
m31N8ua64CPAr6q5B6scOzZhLQUf4ZS7fdSkSFAbAxg=
`protect END_PROTECTED
