`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wp88ZGZWklaj7K2UoTNFgl0RW3RLtKt++he3fNeS/neVz60iLCswe3NYzNh4QyxM
YyTmtw9jPI/VINMwnt44NxnfYgRfQMUX4Dh613prRp8zT8VmsEv6q5w3KRmpVEja
1Kydsx3AkJ6DF2nf9NV+XAOsB6/P/f0gZdUWXrfCZ8iNXVoijSrHdBt3SHAMxTXW
Qi6MRJzgnUVGQpWnVMHvu5+qfD2tJDOFLDBZZv4tekM9Ous9D52g3QTKBeeoTVgp
ovf9qRk9dWVKiELuvU+dUEZ2YSSBhgz38oRd0SjsPWuWtCrRPLvTOtj8D9UHUt0G
RFJ15Liw6jrll+GdFxgAyQqxxfpo6YtjIbhd/n3FzYkEpGmcHJ+e6wFcgdhTmDrh
rUeqmeS3pXYZZQUGh0ODBWKZMKmEWXLsgGHZYVQxCTFR7pUklSW7l90mr39rkmMR
`protect END_PROTECTED
