`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jOm8HWC0L8GmxFv5k3wJLSJUuEdoN1ZNllZAGANcLWVDqnSvMQj5h65GXV/rSbML
IxjI6lvMWK2v7thSkvKG+t+D8VDFrj1NIlpZVOz9zHkTQdXclxZv6Ri/f6lOMO36
Sf6Iny8q3mJhLRwEprb9KqjbDxc+efT8YZZKP8RNmtt/a/LBaNm/TA+/mKJwaIlc
kbd/N9+7InA5qgi4V6x0VPgwmC3PeZOC+QVhEz/GBuGXp6QzaR1tiX3D0vPqPf6Q
GFMm74uCmHk7ZeFhCYtotsvraBQVoxElm3x6tJEvZKVQv+y0JibkSgmkrO5uNJJd
BS1gzfc+xs94tcynGowT1Cq3x31sD/LavqLQYYgj7T+0wiSWzQ7hDj/8BHl3Ikel
wpzkuYfmeYjYs6u/80Ge6EGNwRLjSgRaXBlccv6wt9o8oOyh0ECsifjPaNsPsOOl
GeLIbjiIAvrHv6DXt09aQajv577Y7ykAFwZuad3HVoixQDIPGxJUsiCcsnk9ZWVC
veVaPTuPeqp32H1Fk9dmFZjuYMlWhLzZp7SOTpjTGAU=
`protect END_PROTECTED
