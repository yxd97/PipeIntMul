`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRJ2z6JqCD0Nv2uxGVltQsPkCFZejoFZc3E/o/a0wRZXTZYHfLzBKQR7didE95h4
wPsAbZeHYmDc3oXKt7g/FcAvsGNr/ab92k0ZbOPTqhMEMCgZtTzsToRnGJRUXMfR
LTml6z9SdaPXqwCQR7ISvzQ9Ksw0cc8fITaVrsvuaTyZq9IElUlW8/+bs0qKzGUv
LPY0ZHhBpKZlIGulcqy67DlC9Xuy0IdvgtPgcxIQxgUMf5rM17lvDxytK9SC4Y0P
xEHV/+hPlGJjNokXgf+/3c+m6I6Y1wCBHkV180Mu779k+4uSiinVpQlBLeFfeO5Q
7byOf1ZgYKHaYqrkuXtZOjq3zTwych9wD0fIXDQkgu/3xQTXpk6Y8gdL0jbm1x4K
H9eZPTsDXzrNy94ZIcp4filVN/8dd7Ff4orQvmYOcYSfGwEn5dvkAc/vn5Y4t9zr
xu/b/4yObhd26ltLLzXX2fEBmGq9iWov2ToHlYMRS7xIawh18IqV9HCX3CCvwGl3
Jb+/XMs2h9Jtp207pzCT85hSwAWxTBUM/TOWlKXx53l2kelh4IVh6r/IWKNv0dLX
3k3LVPQK+TvlD+/TLWVem/SW0Ppj23e33FtrzIVXqL/uW+nYLyr156Kziy6kpKmx
3Ab+Y07hOYyYVpMvvEb3/VILOoBF4Y+GGlBrxSq4ptkNC+gK63QCnoV5uKvSr1CH
gkgN7QezycrV55k9LajDPxhnGx0UK/WhnansQetJDVNsKnG/pbrb5c9Pt1rEwKFn
ol05yeSy/oXOwHi0M7QTIhBoWX8CTSkg0a21CnZ8Q5/DI6Q66B4YwYPxvRbL8kLm
OUSBFl5RXvg0nToe0UISSrKhvRsZQeQGOiJnQJvY/aNh2UvcyIsHSSOQqMO1HaC+
9/fy8KUmKmtv3ZmkMCqB/+M3YNfdhDVy84f4iwcOwBE0AqjEb2R9wto6gcVholz3
qfUIvmQhUXkCuZVb/YNF9tCtRr7XV0QbhrMo90sZCpDYv4fWP6TPbkb2McTrAVhV
KkCJStZVV4vM1xI+LYY3xFZIgrwySk9qlkTpR2/pUaklq8v7DgapPQRbYRJ3zmod
laR0ih20V6YmfrhMzN09bvGEJjG+7bV5dCN4a3lUus/EHeS60Kvfv4E8wEEujJu8
7lSdPnwTXHdDHacDUiiE09jF1GUnFor8cK3f+41F2mIu2McTJGVFGXY7QAnWI1M5
FCLO8liU2AWImDjSUsv76tkcF5C9aguiDBKWDkvtDHHW50UqQoZ+6EcBrq2W7Gv9
RYZK+P65/Y7TC35UIQQyX+hp+pJDBFL7J6d59CI55TSssuKPw3r+By6YK0PdhMfc
rE7m8U1TdGYE9bKtC29D8ScX9m79zFIGk4VLhK9P6ihs8K4rNWWH9XD2i2xgjKOt
BcyLdMxgXbYkDos0TjjZMnWnebEL7HHa7KOuOzUGJz46vLwr4NIlC3SEom2x1Fq8
p00ZOukPj+mbSoCF1QZjPJNPFoxFH7Zq/CiN+nEa12G0HWTSr7KwbQz05qzPBrx6
S9J54Y01D3PFwMI5mr86oX5kwRL025kwdeCKoZRa9TZZ1XSw66dsqq27pbFysNp2
JlOcbGIGSFKrHZABpQybGcB9WhLdfh1pHLSqTo2psjKIC3OJjkdnLjRvVdTn0eVS
/3ytWjSOi6NhBwkQ6Ll0N7vMg3O8ydQKM+oQSZHzuHXyRBD2fVDbt6TlyRwPJsL6
roag2GrZuvJOjDdUFtevwMXL3f0o5Gl1L47e/5Um69ycM5xcUH9hupmtkWGqYXHI
R3yZk1m81A4befjHs+sVP11A+ujIlWuhZptCY6OJpAAjtF4vdPkpS9OeKCMoY/g4
7e+Vvbn7FXTns0M4cRPO8hu/KuyCVTsLRr9YlZcfCrnqiii87beQcoAwu5SQyZX5
x2enMQtXFfoV2hJeuolIfAjsoyY92G9sl7YYBOewwGc04LE7+8Krjontp11EN6Tl
Uh8/423fJiAYC2dtZGiQBqAS1nFzeletmm0fDn2gAWGjgtPAlpdK6/sxg9BkPyQO
9hF1ouG2nV0tUuHEAButRWHjaBQB8jGEqFpuHbr0HsAt/3riHX4VgvDoaauJ6ffC
VLqZP7ZfdupN/WA0bzQ60H/HN/AtagaV7RwBhCl3tbzyaxRLEQHweIh9V+mH5JuJ
WFxfEJiRr/QEv2vRKGZN4Cmt8IaMP48VfaGf/M0hDyRr3sYUl0hou6ry3q9XLYrB
R7nCbECvdCQvkad50N5b9hDhB71ht4fmZflxWKqXfdKqbN76rMz/vDIAmeHEN8ZK
U4E/6Ayx6AZBwOJKr3WQ8dG5MyyyTrrvZNFbtCN0YeNTC47mITD1j31NtAEBvXFx
rjt1AuqETFx4Ak4Cst4tEPhjBY/Zn21kEYXBX0uDaNfm9qeYt7fIX0jOCnaRXXcl
hdY9xM9rd8teIozj8AeBqYOEeustDWSdYWbLc3UEEK9pxk+w2G1S4BFI+AMEfyH1
7NliM+ErjdTcxi4GtOeqswx2Lmn8ugFVcj7A7Y1qPP4piy2Z6kjZ7iLF/pLu2mxa
p3ppRDVqZ5amhng5B9eCYKm0hoLtG0W3T8OMXd4zjZISFt10EI5t1qSb1qpi3MFY
ylXQhiFSTieVSuC1YzCh40NGCCdq6qjpnf9obHi/9sL4eww1CZJ8CjTCSSwjOWw0
SkSgEKck98h6oORjiWIE81lpOaaztF/tzXT1cQ3AXJo1WXViTU1pYds4cit0yaLF
7EtropxpFeWZnl4CnYdGdDaA7TKEogMz5pgAF1z6kjAnwlikoEYgUYMFgnmCgflr
OWrSiqCbzrVqYb/8rYicTLD7wABAEaj++lzyqrMbsRxS8FEHFQOqxnfQTx7ACXGQ
dl5pVym8JBSKlCjxl8EAoUwveuazElh/fLcPisAVJYhS4d0U7a7xFuhBNx6CJ3UX
R7tyuLyjDfhgDeEt3m8dv/QekIGZYN3TQ2YtVwKjcxw83Ej4T17B/4bc1VcHKfCE
+PFOn39GKzEC0jmwzE1tQwyriHLjzFkCD5IkwEA13HopA0d8hItEvzcWGqMAgQYw
xOUCKXB79k76IwQgqWpognjV0JeLCZcAQqhKpn2h1DeS8ppwIg/D6e1+BxKw+t9a
Rnu/MSHMEzG28SJTbyJoNFsoNnXZlfP5YReBVEkjLIwsHU4jjp3r3DbbD7Pf0bEo
RPBbL7uM14hKA1F1lKih3H30PJPwy5GQ6tUkTOE5CFBoSDCeQITvuX8w9ma48J+q
4vwypIxv5Q5X11I+7RnQcu3LQZCjvUp2TtORFD1WqpW+0N14BkwdnQgPieIdVvow
BjOf44xIlglUGeqLgJ8hIZChKdmLaI75vdTvzT16G7xfJZx0bboIv1er+o2FvoKx
FeBLn7D7HkcruvNmx/rhB8RGNhx96DFpihpVHcOjjH08dH7VhEGhIbfKhRcPjBQU
LmjgRUaj3N2Jd4B0JVIC6tMnmOQiV2eSlyqg0J8jQEfFr1yp070yTAaQQCz+Mxcy
d0H1mY1u4NGhpPwUyRIOPUkS7zmkk42Vcy+Vsr04ogmNLsAUPTwmwOJXJlGZjsid
/xDTBWG8/Q7qTQ9XRmDso8r+xmiQF3DP9JYwnwvwn2HxxsIGUJ0xLycgxX3xXuM3
klijjXkuUJlPpgOwEXtlXOcnnq9tzmZKBFG2qf2MpJ//OBT8s5jlDwsXHZrCrH5f
beiwV5sc3RrDT0rZdz1qEpblnsx7AHUR7KCFcaAymmgHBMUxRsY0g/jCOeZW9z62
ANkQnfXBIvFIVaySQ4vb2ytUVF4x4J0SCVdLEKcxpbOHZ0/vPzkXBH1hPnGCl11V
v0iaFf8WoGUa/xqXWf5hcqpPGzie4W5wcKFhP0KPXH/VDGogBNubLFtKzfsycL8m
FxhQ/rGBrIbV7D54I03UeGpxBMYKVm2Z2f6OagQNpqpBF5TELNyvwqwahEwCcQ4/
6fl66PHY7QQff83ROGVE+dzt6i3+qjSop1O3KN7Mrk3LVC5jgdzPVeud9F1bIwYV
GAwrhgaMyRiJA9jPLw7Iv1VWZ1Be2bwpT2d56fd7YSGdzt6g68VE9LNiVB8pOrBn
xojdm4HjMtlhYTwoj+9iY9rcGRcxHpICSNwgLjdxjjDXSeR3hl48PR6qgnLdfL0U
BLV4hcblYy0cgFxcIyp4lc4ja7H5Z17MDafNwi0fuwuIPglsm2WDv6hhEBXMGljO
mf0qtw7oS8U7l2J3HKY6aRIY89s/c7uB/N4ENu0MW5onh+PfBGn8u9/5KU9fIbJF
+DmcHW+RN4UxpdWQXd5cv/RirUowECH1ixTgK6mIi3E0dLJrxgqRIsvQZ1G3ase1
GsVLlC8vFcXBeTAEDLM/8Rf2SUeIETpmDDf2gsgExO98YMXzLLje7jzXKEd7cHFq
HrJu9A+ZMSP9EeXItwlZkBJaHWT6Ir2sdSutIjRX7QfUZRWvbiywwwgf8A4GJGqn
hVSWublTVFQ0aTfl5lQtZ/nC6J2poXg5TYO33DXqBY/UDcKS2tk/4lhikhN6kd34
dy4VDw3gShONNJPKU/7RVA+Q61sAWL9pcPG8zq11Fok6XTLhX402vJ2k3/32tvY0
zzTufnSlPqFmDxL9wpKuyefgaeYXEdMEqKLumtsq4wSHKmwUnFwG3QOpiE+MheLl
zEALpKfxkAUImex8PNVoHUe1s4+8rlv2JecZN/ojRGUh8VJoKIFxifOx0ZbgZA07
QCC2ZTKvp/Q+4gQxPaGcZseoNIvahnlYKlebdOsEIYar3i1xGpjfRr+stF423Y9w
5xmNr8uKNz3KyniDJDkqHidNjBrRYWN1ZPLYmUbUZR0uXxqrEL6V7NSBXOLSxw0Y
X15YOqQE2wcBLnuA42bKiXOd3jad7bfAHS6JwOPwJP94vFJ3y8RMQZve0xzfZAD6
Ki6jHTtPEB5mmGkzn4tzGssO8aEiSWsPkLT+QL/x1ZhAQLPZxtkcc2ixJOP3MM+q
iR6TE0rzfETN7h9ogDqOXpAGznWOZwvMKjVqEBEILCr+mYaogSG0/GPlSENMU3X7
NLA7AjeJ+OHjf4C6sh3SLcwhVE+foDesWf1HJRLVzX63Ywl5llz777YEmL69PcTy
lyw+KhhkvqZTddc9jW73DTwDNkc0GBMHNUinNrQflyzr9h5jvpatDq1PsxzbO+pk
1e+L9BfEtzNgpGtrOoAw8b6Jesnco5h/coQPxvBDVmo3VrIS+/W5mQ9l1yavEgf1
bsGm6g3Gi1vE/x00fuVUsc7FWOMHibCQIAIDPOftYI+nWxnrHiHZDUCEvOPcQRNH
7qiiowbamKTnKzq1TNoG62FRpnkWLvRfD5FlM10l/h3vVk2/N8eOXx/U1eX9eWcn
3KZbAcConJpvxBrisWBDmk7mOqBplRdHMaaOv7tod7x/37UQFJuNiF+0jDRgxDmY
inYPqxv5n42+4LRuCf5zUSgoQlFmwMtPe9aGRZBqSe7MqbWoNff549PTFFj5S23A
ohkrFRDM1mlQ30i5WgbyEtzTUdA4ZoWLsaq2MatRzwGMQhbxE3aKfl9xBkDLzxCZ
SSHPyd2/vzKso1UGQ5JSvBNpoi+3h1PBRseGeLx0khjKFQ8rMkqcXoY8/+4PKUVY
jpMXBLtFp6wIjSGyr5p45FsG2XsUhBCpuAq8v22Pl23bbql2O49869KvTXOY4w7O
kB8dHVpT50NoVv0/uFJpsWafuYVgSKvc4X6hlUPeX9Xesz/A6WKUeX8QNRrEqhXj
Qo5774fdL2VI2k4AYDjRVMH5AIYytfK0v6rOucV6runS6b9N0HXzqAZcxRgqpuTs
3OkxReSNRMAEvbah3U+jZaOKH0+i4J5IprorMVId/ZRWD8GRB5wo3fnRDNfL/SPU
YhtrklHWqBYQvNLxGd8zAzR/5jsSBh0QXnwpDnMHJIyvMIXhTnnWrLJnrLb7JWsC
Q+qPuVBo5qJBuXuxC0HxVGTzEwiR1I8uDc5PsCpy+2AGfu+fJQp6sLHmnrl3KIYR
abxZlVha/7X99cdDf1ucKU/9liRo8L2rX87Ddmw6oPI187h8b1KZADaMFN3qoe2B
U3wEsDihU4lbadS/N/l+U+8rI/OI1IP6DvankvkeObdlDb4stkTMrk5gubDU87Zh
UVY+72r9lvwer+PtPjgP9OdxDzMAK2QSlLdBGi5Aa2UBc1mF0cuQQ0w9U1rSHLTi
mWGbKSckbHFqqsAufLYFVmRMWqIjWmdmaH96MPSjjLThQscPROVxSP2vjAZKC7yF
8ZIDwL7e1Og/1fBgNSlRhql3HXmyUIyqk7QKqXWwIkqqSirqUSUnI8CgcAmWbVse
2yMweUJtcUan2l2ECIk2cF7W1YyCryaH4v5EoCiddRpMh1tE5GD9aROKuqREmhRX
m28vHtcT32v6oNauY7cA2Sq/rSMyACMW0Mq7ZfqzbcM2zrOxXqFA7JSHCxTZEzOm
RAldPrUzb+IOOPUSMVE4Rbj4WeyzusRLTrXMv99t5yP4dxv/3FhKthQmERI7F4YU
eK5rTXtpGm4VeaRB8lWcdt4iJc2JaOjYFjZvjuQAp7ceq1/hVGM4gTiQCs8Ov+ZE
i7LyigQ3Gt1IMIU4ic2/I/FfyMbGiDh8EyGOkUx8A7thNxcRHDVovJ5njRoc5Liq
Frnn8gFATggWNC1m9V20nrbh1M4gRz0aSVVJPbJS3JMYlO7miCBqZZb9+OI3EE/C
b12jlA9SiNVFds09WP364z+TJR0GGAurtKaQMNCq+o3I5OQa7BANpWgK4e8UTHgE
+ri7tojj6BYbjnqP+zbDpG9fjkgWUl8OlDlVgLFBqcbw/TieFma++C24F6skJArV
yxs6N7SOoAQHRNdAMbxymYfHQ9uys+YTJY0owCe+LlTjBZ8D71zS/jm8qb8ByGGx
urMIGmsiN8ZU9RaqNtPU32ZSeF1Zj6JOLHKAVzxmfxhW0GwGOf/9namp+c1fks+n
ZO3vAGRHqVWErWfqJE/6WhU0NfDuihV23n7uqS5C8LAVjAgO6Xn+1UFKZ3xS3SXy
YKNJDJobUoTc4U1LoMl9eTCSCPiJWROuEpSWs4UuWeplpvPAzXPke7FcTjw6fF5C
024wpNYpawFhycD3qZ9agc/AeeoMbM8Agtw8/8FowfqFZoGUtAchA1+z7nqsppfk
4yrCQilCimAmbCDxlO5Vv+uFKea7TIb40K+kNr1K5X7vfispH91by20+U2sQtFl8
PfK9iyMyKPb5AkdXrJcMcucaC3pwRfsgv0d5rk1bc1V2fdaa/fUzqw6m2aR1Yx7f
HMqawZtvF3+Ex++RQIsTcAjt2ocTdGBAje+WGBDOHcVbj/mbdeAtVLNpm4aNsTV0
rYEsGbfxGseHkIYOJy8cNKNaPhB2EAFsb2+x50Hj4gjP5Lc8uSv0sTeRIh9kTxt+
a+3zNHL12RXv53biUVa5dvFGI+i/UGtNAYFc+rDkLACuQpp6+0dsI9Wsz2ebD22J
UaNcsYWjs9hsLP5nkOwENYdVNePOWGOyQ0HWVg4bfwv7XklASVfUemgDnLHc42GU
9CtU5Fc8OiG1Q3GtdBZwEQ+CR/U4jX1yIJpdLSha3yvbBUSg1zTul35Mp5sZ4NQN
82+l1vqcOWEsEuOQbKota0jTwrvtwngb66QtoWQAJc3WFOOPT0hjz6rdgItYL0on
5QwPOFiN78u5mQfayrAwmKg432aTz3KIjzRzo07Z66IkqjhakEA2bxNjntiT4Br+
H/HrETYwYHvbYmEDkrXeTWdwtIcXUkqd5Z7PE2r9U4Mtr4FEwS+xRHdJmkujz6Aj
/AEk+oZCvJm4bhyy3qq4+Kluv3NiSUdTUMHS3Jawvkj00MU3QXJTD9SwNWwfZ567
FyrZxx8k3HfDDt/kqcsksrYl0MNJSCTC4sXlL3aUXZzr8vSYXIGze7mYsPIq/t7p
8XVGQlFc3akVXMQ06ez+S/pC4orkpGGV8dY2k1DYZayrC1Zv/hO0L2cyF41ptNik
wsrwIRm1sEjI73xQt99qSF2vI2yUYrzyF5m+STPx7A9P6BXjeH3F985dHkYuIuwf
juRwo2/M942EV0YelSzjnQeD5Gw6zPLGEn1HzK2ESn9ZvTB4mH7JRuwB1mvmbsJL
b5fIbxYV/vexhXmPujeSq9oyX2XfJ88JxZLd8QONfePQhyWUyobPP6Gs8T0ksY5h
lTssPVhUDiXokVEBClzWoOh90qcfKcFSE30OLDIO00gbjHN/YVFUO2ZRciCGXZiV
l71NmDWoPjWp/HMyLsYRrG5hYRhiBAvhb1M1QOKNx4WylitVffsVwitut5HE0ogJ
A36O10gv85DAz3dIKXLbbqbZYEYijCbvG/kAe2F3KutKRGF9gJYDVA5Lbf3eAlhJ
deW77EKh+/9f5soEcVGZuGtQdvA4VeruPKwwNEztSVOoUCbSRGgoMSbz/mc1ygJY
FT2nB5mXHlA5VrMM3kJinp/S+VPLDzqyBscwT4pqm06UMyNAIQQwfPFNuAhJEMjo
nDbCybo9Eri6azhTESESsQzBeykn+tnmpn86X00yqIU2ia08dNZJulKcceTrrVNY
WnJjxHTlVE4VcMqsSQLRdJgfBs/EFPKZCrWLWxS0awF0gEUla2nHcWmt32EPLOqn
SCOBWd2tEbHf7P1g5a4IpVpJeuoWdTEukWq+b3Za3IpAVnnLNCkg9U1B2cfuPj2l
3id42LztJAPTS+o5by8Aa0lA6ecU5//lminedlDQHAQK1248a221QAnzCZ8m2/Fi
uQOymcc/dzY/9izGeQGEQgnt/RfyNwkN3QIAU5tFe9WYtrLgRIsR6nozV0ipa++V
1EAl7qZwtOQ5Gr70Bco6p8CepoprcG9JL10z3gwnL4z3FcKLb1NUtTXlytXZOkFB
/W4LGX/ievCyLpYnuRvYqfxTNIaFM1iA46VDvL6btMvR6dgVtYCQO8Du2DnZGj88
yCzVW1LuczsjB2zGEbFshFkDhouSPt04KtaUR6KfDAhBA07Ratz7eedMzus6xMKb
gZLKO+a6cDWGA+M2NCYBL4c6wqIVsE6yNqH2ITPUG8G0NE1cbRKHf0ta+tVWA1zd
JkeRkwIbG8oPY0D/Eid1r3QiFuMYV5wJ/tfvsIS/DyIXkG2/418SDjTryW2BFXBX
wJjXrLdAaa+9xVAHDg1bzn++bw0L4550oGgToCBT5Iqg0odhWIFSq1GemmFdSFEK
PFlePcveaqzOtt2ioJQ8J2P9rsq924BvgmgJljP1jyVLxhzmvLpb/VegCKT2J1Mv
zJhZI1oBxfsq6Ea8P7hJ42sVu4JfpFq/ImXIgcKMAzVnomwZgLW30ajT664+0nZ+
0Ox2sblGEkE51VrASrydTGTB+VG2yGPMJpYXIB4j+Jdnt18B4prZr/0HoJBR4YZ6
WbmjkFNexOfGFj8OXfANgJP1GJ9oFcE5phT+YNDNreexHCTYVYIJ+Cds/zx6NWSB
7NEy+xWALdl2Zu1DoJcaVi6j+G3BxzEiZjajf8yee+ylTvJQlbqyTTKb9QePlkyx
7csl66W/oiGXh4eV9+NdxzbogtYw7GVqu2zxcRgvtlEMJESC6su13WMgC6aEYt6k
1NZde87XwjS6Rw3R2EprRZCwyGyao1tAChaylAXfpB4pY3xaKT5MAU9akrjpPQz/
YbWX9DLAFOFXtMBEG5T0RdbqHaqdE/1qHuE0DW0VHD0KszIS7MHfI+tlfeVBuYXo
pnqZ8jFJ3+Cqtr5naZerw5Q7JqPe5HYXH1jSy5YR+A7uNUeW2ubCyyxNc45IrOYf
BmxNKu9zDDC5K28at4CcE5J1TNm3J5d0dieE53dyA6PWUOWtM1mtveSPurVKO55G
sNfc/TRpozRTaC7bc8dmb8Ya2iTOcJ2H1vQleeN64VsXf4hxZWKUwlktzGWZ3CNb
Lqxf+MIcyYaHVulUg58azFnRxQm9NEYiJQjncb3uQ3UAfilTCpC/g7fPnmmcc2wH
o2wBLVHPay243WDJPYGZG2KgbpjQRgKVeEaFhN5Wgyi99yoB2Rg5QFaXwWJv8fqZ
fxbiYIjESSX8dAPAGNcYDFGXFWjQcqcV/upWT6Tw4n/9521bkfKNpfaoiCYW3l9w
bxyeIYBl5/B69TOLDi3NQPpvdKMKNqosgJKima9YexjA/n4kXi6eeh79gb48aIAn
vaMpQgDosqufmotMZD4bmOCHhMpW/xbbIuQBaEgp6A4/pU3BSkPxiu40sdljGaFd
cQsxBPjVgrXhAOqXrMYSYQwm/qXuHB4rKt1RDdLB4lBQ1VwwZEy17nTw2l9V/KGB
r+CYz9AwX94Bp3HrU2ZZ0S4nxswKeEpiNz8RxVKrwmbBD08B6tIAv+2r7x5/7ZId
3pez/1ShwY2INTewNvuhBVahGWHuoEmBiVHMnrAVmA1k0U03rDJtArheclu9J4am
qXXzdn7jEbFFZ9ed09hjuxHC6Nsg90ituA/HioC6ZBCtuYv4BTKnFdz4oV+4eWHw
QQP+Rjp6c5G1Lay2JihrArsDwtiHaSqvMQbPA8qK+6+rs8+nVfcnyicI8pzR/joL
iEhusj36b9RWwpNdhF17pTQbnfmA0L0sb1gaTGBH8QZH8ZTqaXGDdrqTAjztIVTH
l+UAJTXOUZuBE7LZYV+p/wuR7R9ponA5gnDlOWcV2i47lqto0WgUtbG5Q4i6tlCy
pDefYKwo9d/qgF7c46d8vfZvBqxFErnl3/7j7W09gdBanF/iGRjcYK37tRAt2fAO
AZDKjT8iOfDE9Mxc/FQVbadB3D507mp7qKSFGkEsV39ZTXatWX2pa6Yp87z6fRJd
A0ynB4SZvzyGpVuMN7qzHnWr4RUvqQpzMEfrThLp5Xa9tYBqiiQl5cRZYePagqSY
MPq5Rzt22ZRDWQw7p944QY/i4tpJryWZaYLvJBwkzb56cxYBOCEBywChGVDnogOv
5t6ne3QNGcg/imaj5C7jBXegmzSOyEXcmwAPn7ZHkpm+zUXZCu9b1Dd0F9/k8lqI
y44rzL9HR9WnLSIbB/LSXKmH0ezVnnSkxgVfTjnsTJu0TFL4ueCgpOx1QQvKeFrS
YRMIRyNgVpWOgTmKMqLtNexfCu3s+DQn7xPbijhpw1K3Hqf1r+DJ41+YCl9DhCYf
F10hYKG4OO5dwGkVyUJOlDDNMnMBDaTiAfBE8WUoDMjBYITwTBruUtFlKR67ByPy
QSkAHsUj73EK59hNhDhQLrQsqcUETt0d8GEWOJi7SKXi0bPYGtyvnQSUwGaw6kwY
5Ts5HXgnEgN8bm/6s9Y/vYJPS6sqRn1Ey9w7auhWIPTGdM4gdcPHd8Fg2V5o+8W8
eMILEKPJaeQ0leR+lEyRI1Y5KRqbjZAToQTaWGRO69UOowlylrwRWj9pZIC2ClDS
zwmdpV8yKGnL5dfBUE6jAIRhc7YehWduH8LwTqR+YNQFKVSRGJd+qpceztiKwMsK
XQLQdSyGDM3oonfxetMUbrXZbWejsDaGzIhQNzhfwUhqpAiYox904qFpXBRixURU
jX7oSP+Yy90aB181YqXPlghjIK7DM+jz0mcZwFCcUU4VuDJtpP+5JJbkYpOLwBJ9
TgxsTzQAMC0+GiImgkU99+c9YkZD3NxHhmkrGRUGDPZfyRiN40uUNL4JEJaE8CQ5
d6AZ3qDOtZH7ge2G3FZk/5alTIQoBiULW+6yUzPRqeK7YD3D24K3pZvSm7AX+rXj
yijlmsmUcJsWXUuAt1PGultflcDpRo7NCjwR67TXTDIP8N0wOAQ8+Anwal+FFU3/
NE4D+e0Ce0Y4LbOzkW6ixhXitxWbsMUkgREOnqMJtl23uf9lvdYqv1EdlfXt7xdh
bew2g33MhEOF8bICWswavOeRFoVpLl9qS3Xi8i1cBWmu/97i9hzXKsBKZ/nB3hdQ
fKwvmMtdgB3cJl0WJrAOxltZMP7i/sEa9husFjcPr6MoYOXOCcgFxkv/cRX+kbgB
6KclytYUvgbKm0SLXVmVQO0jizurmxfVBe4ZRpVusNbIvi9B9S3OIUpw00/mOpZO
i+M1uDxKbFY14m3ERJY1F7sGCO1MIcF3TKB9l+Vh8uQm0cuUnRla7j4R0m35WdK6
lr31TdbbOfVnBqQlXeUCy5uXRDe2gkF8eHxD835vKj+alxEfvxDhZwrgii2Y5g1i
72uiKjWM+r2YivihjrQHR+UlOr/WOid2vwN/7Vp9+Xeb00YmFKTmN1NsvJlxULVZ
c+iqBV1SBn/qfSU3qOkpeO1gBqaR0oX3lgO9cxyL7dBYLV2qFclDXZh6YXMLhsHY
Spq2JEo4/0lr3K7ZRno3W9Ybcl65LdvGscUXYVUg6RGkK/9asH7wDeCUlz4NcYbg
b3x04Yux4lSJL5DwEUTMOYRwHSqThfOeBdbMLF1f1Xa4OvoWFR9sWuvsTK92zK7A
BeghCkO/xldUyTtS+JRXfcHHjSXWn8o4bIR1xrRFRtlY9K+qCT4MLaaoHyKM/Vz4
u25C1m2XyNOZFBR8Vags3fsVkpAxNuWuVzlMirL65+JDPIfj73S/rzu0CV6CggXv
tZl+F53PG4WBRc4UHQm8x2ojwjt+6wQk8Y7hf14hLNtky7Dlc6HA1Uxou4T4Ikpm
RGwQJ8gEJgrH6VNGAPS+GpQ7yYjm1ylKdTDwZtso1XsHx3fmjOkmseZjMmqvVmSI
RfTQilvAlIXc3tM3f2vv5iFSYz8BTH4In3x+yWSrQoCzollRQ8mrXlx+Zu1i9fP3
eOJoYLra07YjjZdizpApwJjtH12GB1rRnqO+cGZzu5hOFy/JZ7NEtMNRoWg5Nkzv
0MU06DTQb6mLYUonkDfrjZh2BRml/3CaIGrYIG7He2+GzGSC7ORRYc/gy+dPiiV4
TXTbT9oCUypQUigYGfzF3wgI4gfMTOzM2u1ghzAtANqQKVgh2M8pMH/gG3ijE8Yn
DUvvO0LNPpp8OaBZm1Ps6zVYU/swBnKLvVXDaEUEg/zOGevtRbwjQA9PEvA3MVtL
8/sGQijbbq+T1tz0WKt3MiJFMPDxhaWHHp3QT2JLOJ/9VmJAqF9h0ULjiVoqPd7C
GWIOehSFNWj5MDXY14G8Dr5v+senHzJtbKYUqV85InsRJC5B9CMk8YzR+LFR/H2b
54RguedpLwD2kYIfwR6q/Bv5V+py3vXyx6eFQeTRTiJyVmZE8zVHHvUc5zbnJ9u4
Ip7ZPQLn/38nGdlwjmDvQ9kYkFOO7VZKa+OkNDWZb7WLAkep70HVjzifM/9yZ827
D1dKzLw/9WGl9ViHisJYllBVkKipBLdjsqhNzHnRHIx3mmNldbbPOSLTalhdgKKl
QVhXY140X0pPh9iSSrULDomBOwqCCYYOVz6hBKSL8uNW7G0nCEsbDykPFxDzws2Y
mzykFPVIiZ9X2MbhjI9rO07nHj8pajFtMuSxpA+7kjuDVVjZmZfbvC5c4PFJLmfw
I+U2k/GkbtcTUud7g9xMJaP6Q2oqOxLAsDED9QoN/ugAUxLqGT0zJBWD42t7w0hd
Sex9n4zyq0u7U16H+8oW7iuI4kYWq3RoTlohkRzff/IPtSpH3VT6JdG97TFuIrFF
J0VJfTvzwiPpGH1tSGj3t1Mie711erg/AtOQDLgR3qztCHmmXYUlOaEeXIg22Bp9
L/ukFvEZLiJFZB72Q+MjS8uJ569YDfYxIzKj+NptB7mHVWheMdFqrdgY3jCXwzX+
tP98DRIEgwzyRIdJSTMANdNXHEjAQiSN3PYmteFnhkmKU/g/CgvVQ+J4GNwU/Bg9
QjU8rx1qcCGWz71czcxgwNnT9/l8b2lNJnz5Pq2CH5FF7p9knQTYFchBitajNxtN
ltnyPDGzNQTweoStJTDy7xhsx/srRKhuMYoDnd0pFnb3r5wcFaeDClBWboBb9thH
Aq/r6Jsk4x6lB3K5+qnZLH6N4TFS0qe8YrWpQt17BK50mgyFClBElOEhEpJHhb8X
uLREf1rga5vPt8NGZbSIwNLor5yJiWWB2B74jz5JIIfgCz/FTesmwhM7kN/4PrVk
GHEzGqxcHFLjtBDMTbX9VvWn4LoU0T278lCiACVGKhRqON4Ee8tLM7PmtWH5KZvM
nRRqQqF5AI4+mECd7ppDihrMBLP5aMsKWJMfOtsZb5tV/6MxQ1Nr9Np4K70oNiTH
HYrwrtsCeq1iLiw0+bgIosMjwexp4b+ijAtuNBFIkwMflQPqHY2gU1VwtleB9OY7
Lhk/rf26kYw3OxnNyb31zgjKUCiIINg7X/8TlS6JeAcn5RtZy9+EYR6aYyrF6GxP
RZfz07hWTYenQaS7W7M507t1fvAKNRse41dTCKMANZt7tyQUYEkN/A8w0ggkRYxp
2O/2K7gJfrJdxUeWG746AMQpxogNF75O4DkVsCvH7pmfcJQXj6YeGCRQM4ouDGuL
iqqMAuFDGRCx72KtCIO32FB/fCIuukMcJCNHpiUwa0oI4pH0XtAgeLLkj6/Nf9I6
tWe7AAQtRx171quCUgrPZc0sVInxvcXkY81wxKk9//yKtvrBvL6qABZcOFBKydAx
O+r1eJFvW7iNnOaT/7z4gmx3JOuS4+0qYk0b65uSs93m/b0Oq9RrItcKlM2AKGQR
4xiLGVSqo90xZPVZs3TWvsOGiNCrf2rw9ij3CWCC0KVwENMF0GQCd/fbP/Rm7q65
KedBSp5pKXovPk11JpOzDX/Ry6TFycJfGd8RFJaZdEkRl51BhfO/aQsAO2QqIcd0
ivjAg+fjXZSTtlUva5VL2RyKcFZ55nv1rafRMWUUoTHBy9pDooiy+otv4ZLjzBkm
oXrF+hew1rgAPBgq7GdfEZCzZJU8Y5xjSfyy7RvkSZJpC+/nUKn/K31hq1+nupwQ
D+sdm3vj6kL6NzFrYfrZyJpjVnSrrgTBf5B8/2dGV7/ALGcRLySPtQ9WUYiU8ywA
TxJAZpyPpOnxydOohcr0zVAsgfcyhQw21W/QD5L3U4s5BYO/VdzPo31DcBPYlDql
LDmeb+30Lpnql+qkP9G1XRAevxL0eNpW2DR8TrZ8/gWCHQC1lv/hWU6DHVgjYZL6
5iEi2RL+DoYn9v8AWR3IiF1c57src9o5WLYLXHjbmIa5QIyL9QL+IGI6cJS98qVU
VSFgVumBX400YDbWEwTM6wpq0d8a/lhL4W9rI3Sdh+HEkh8gE6QWwCt9/ftGQ1cF
lLendrvhqMX12elroQEFmDdikZeuOkPpiiZVDBrwtkyzCVL/ARBI5ARQMJy69N6U
EN4bNkVbEKKhKIeD2awx4Hu1YapYoOeSheRTlz4kRvn/PEz4hgbGgNjAeeFQj9It
3TTd2/1tzAfUVKKe7mQmJyZu36sFw7AGuT7FUKUtfVugyN/cZ3AnC8YqYHDmsDhj
RrDDaqFh6aXgt5Z2x4ny3i69iN9/Rx4UhRsCxvGCzt+8S2cdRv06znbUCZKTMjPd
DzamUtqO1PHU7dy2GXklYUlYAxTO7uzOhFOJ61tnVqrY7dVPOLzeDhh73fuwtp6D
5OyONN0fv0a4w3drrzxRnbTID1rFlx9e1iRE2M/yjjTqFDw9W6utg5xJk/1H+fCW
plu/+JpAHw4AcP+FXMoC1i/un7YrmLLxC1O7dnYq25L4YMsF+eG2NKzjqhxK7TQb
sF5QA0+YWRRJn4OM1Vuk7eW07paMsFhyqYp7KsHuqzq9QhOY4wmS1H4gJt10Qx8+
vqgqi3AydmOp6fA7rbnDPINe6WBvdAhGTUWsiMRySM1RbY31a8Zj1tc9Shoq+sos
yBNLdIcEoiSajN+2DM/d48Rmr/6/1cNJlcLGoSKZFMUjtaYfZj6MnCOBWOpbMyFp
lbmTnBLaOUECrf2huMWcUjM5af2V48FKGHy0JWJ3/fLrmirov+RF/5zJ6UCQ0kfH
8pVFw/oyRtCO0VyvkTRLG7KUjcgc7GM8mlaX0LbupOtxGdfVypJttR8x5GgViy/i
MmuFTA1XsJo1emB8v2lJJ6NU5JoBXs5lk2412ft7etgEZITIbhrdwvXBoEadd/Ec
+CeVhn5YZtATuu53wo2LG9DaKkPR1s//1rpxoylDCmVhRUa/wbKKuaCGf0Lqf87M
iUHHELOa3H7v1qPXyp6COQ2AhqpjVbGDf3pMgotFo2uMQfgbeftbbqE75hAxuQ1x
S8XGFF2g1jkP+Hp/bP1qgbgfSao+to2wU3USCUI4KWunpLg0CuXZmT45GPLjLA7Z
dlKl/cfxbd5OzaMuei3SDgAYahPXSMzaKVbXUXw2KrJx9xtvBZxwhj0SYq4/JEd1
vOg0QdgVUJQ6itzxDqA9FTdcmZP2AhEX4OL8CNH/NA8UIcrnZ0VeuS6YZKPqcvIK
5jul2tClwMBt1cUOma0VsnCH8Y6XECq02w6MnDNZqoEj/t0UKObGJvVnjpAzONBc
kAxOSKQZYXIUCg3s9R81KwCnlsAQJREPJqMn29bywWpk7sfl6uewHbapz4F2Ro4A
qbR0JaioClCVN1on6j4du92/gvtbRigDo6MB2U7sdxguD4pGfqDMlTuDbuQw2odO
zlJ7NOg7YXrWNXTj2LKroS3li9tHaHl3SkhUiIAoJaw3K9WKL/rEIOMJylGlr9F0
NlJZB6uzGot7lVip7GHq/qd0SFu0tmvmKUAvKwdM7gI482iFkln0P3lsmDVMQMO9
FJf7CMgZcPvZ/JN6qPFnWDM2m2PtGq5XICxkdnEbEpRHnFJLxx8HuN2cTROFzvTd
YcNTYY5JF2ZeO3TX3ahXfSmnVkyU/spuR9vBC71E3rHjBNdSuI3VSBy1tBUVGA7Y
ngR4+Mx4nZtwlV3lROAh0QHqUBiJsI/V9k7iXrh5NRORndybyud3TQyi6nmguzu/
sVuOeMAv4cxhV8b2OPfusRLB57O783j01AM0/l5SsCcsScrmg7IT5kyeXwlHxtCm
kLU0siIPVxyAY7OXFwDiRA3coCUZ8RsQUqBJL00x2Azhl53IL99JXMBfFt0G1918
4k49HsxGwMKV+luedHDt6j3YrEtqYaUMAjRp+jX1alzTpL1NdLIO4bujCUcvXY+W
IMYELAQGrLTjk1HmTMsM4aLhW2tJG1qR84DZaACMmp/D5C2sJmY8WR8PUWnK2fEA
OdSDnb3/KEtnV1rfmcok3yHLq0MV7yOFuYBFucGo+ibolCAMvI25mnqROQ0GsqIw
zCtv30JcuG5/iwasJ634WlcKEPbE58+IlIQPcvFOAXvXfcXJI8Oc6E/T4zxkmXBo
v6ZZRwQQo3jv1Xuv4RTqJA4CcAKlqisL6v0v8T3yhbwetj5U4bh8PU24DTtm0yt5
MuM3T47kd28jb/q3YRwLRNrVE6Qe2ZiX8exzfxDjat1X7J4V0mst7znr4g6KIYwX
dghCaVWSEOxRz35ACetg8Cda+9aVJS3l0oUomZECMwg6SdB2oA8UYZj0kWXfYXif
TKeWroaqF3ccOBAj4BU9ESyelgOjV2OBbUDr90jiEs1ytSvLsUSoTydbY2BiSmB7
XPOrj4oHWAVVFsVvockDadHSiX5dSa3oGzAn/sjeO0PLdYAr4sTVAEmCcaDnDPl5
EVSIAeOlKO7m6SvObsGg7cVKs8SJQxG5YwmhDD1h++qZgkSX13AJ/BN/9iJuVc3d
AFG9P5bHn7nNelPpSZyeJdKEQVKqr73U95AuH3cUpuC/h98O8yTDDOAq+pYIvvbL
FzLFcLVcowTqoPwTfx8wIdqfx/IHzu8Sh04w9Ft0KNJe1tFaKVjLZFvlySAi6keS
145Dk7YfsfmES6vTmncS91UdwDSaUJB9jUgRR1u+SsanC+pRVFsliJ602z/UFh6b
VNt8DURFyGYB5DZBC7VBgp/qRijFQQBN7CaeNlvkdi8KWT4h3f+ChcePo3RQf5pU
yS0FPEa6ssbuEIXJE7ea/1S837pygyqzi0d2WrGJQaWO7OzglVzjblkD/IHwj9Yx
VTVjC8PE7OR4EWiwRd874GXNBaNnsyS4kV60yNQJX3z2so8YZpeSivi0StwWCOME
iFv7Ik8MoUsgjgPrNp8Kr8J9jxQ4OI9ywcs3qua3YK+gqbiBCEyEozn44Um0QvPE
tNRyKc9qYONeTbYA8kHrRxudv/9NLoX9BefEIVc9ghO+j29ZSfgx7IY3eDRNIjJQ
CC2Rg0jBXL5ZV47Pt6TwjyWsjWGsH3yZP3DA2LdEWFw8yYzuakaZ+YQRV3kRPwgZ
WdQWlVaetVJZEJ+6svF0Zn/qClGe+rczbkV2JCI6RFNg3R9SRkoB0UhjosZVva+P
4Q3H256xHAxQvcEDN+8iyRl21iRPE0bzHVhO1CzRcWo/7LjPjqmo2jGJou12hUM1
H0Qi0Gevpg64H/IcT4IWlNQ5N8xa0ogciPjJvdNZb5RtUwrqf0dfquB+MlC0GsrW
Q9BQ2NjIWryy420Pc/cl59ZsZ6Oce3yJ+BKUOOcun25dCQUnzHyakuJwyUTHpQVX
+NU0GJrkj/LnE5Fpzub02nWmpYvaoKWPrSxR7K0+gxFyiQAhVZmbOLPodH9ET9kY
qqrU8yZUUwYmCZknBM4i0xQ8EM74+3FppvRIYvB2GVRb0bE77XD5Zw4taQSDJE2U
GtfVFpTDoDn6SvltoqBIJEcFpz/rQ+e7QZ6DZSgQ/AZwJC3fJLTQaQU9g2Ceu7l5
hxQJrhH49Cv9cntLPIG4YjE4TOj4lR3iicEKNPzlayoOHc4pj4/cGCbn5QQNbfHf
A10m4LOe3esxL0GIkAT6mLBzxoIV8TRgV7xxfINn+wemOq2qm6H4gDB2ogYiqaGg
6tRZGS2Ru0obIPptgPYJRqd9+ORh9E5+nmjTzz/3OWrCH3SXg4mqPuhh4fk/rzvb
hvtBI0gubYblYsCj9zBGpn9Iz4VAsySHx0hjqkgZG5unweq/V4TZWdouTVHyM+nM
9WPvQiBaw0dNUAHXT14TPt0uzLlyGgmgJvuVKDfhaXowtjFaN5BdD7hs2eCcyetP
tqhOWZBqe2yshVNT2/88UkOlr/fvL8bMiyI0/rYsyZW20qSnClaZuLGYin38tQld
`protect END_PROTECTED
