`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+EwuibjwolZiO+4VtYx4H8UIyLanIw7TOHkLGG880ncRMdPgItswck4qB0hoKSu
l85RVlf+7u9h2OYf1xkZPiJ2K6F7Pu9Yh4h/1qopBWdUS6fqfPg3JUb9dgo026QM
p+woXbvZ5dPAftoha2CVvcDG2HFCm+8mWTMAa/qCsl+K3wfw0DWT12gagXoKp6yz
evJ180fWa+p17WBs0hRCHYSnGLTzke4aBOjFVxlJevcb5m30EHSR8mATGd5OQ4L1
0om+Sq74DvxSkiO4AIyiFpZnhc4rYjykx51zf7MT0vJ64nE6uq2TPz7rCbD4+xaZ
4iuA05+8hMexJKwmwQldLt97oko/szqNPhiI4Vln7/YwBoNTRmdujfpH5m6AwhIa
x8GhUfbAnYS622jUXoaDJMUHyL+kI1eXyW/jHt42J9QvqS9ggtzEb9JNEI3rrIpX
yCWa9n9k7mIkgqB6/vlQcoqQem6RM3fu4x1IuIZv7M2CfdUzNRkjk87cDRTSGv2D
LpC7S3cRsRmPJgnKAzAzscafOG2CyoFL6lNUR08GeMDvGB7Q3kuBZ50cACEjDukI
5KAi5ybIJ41pzD+NkpWnraeTaoQCIOk4VeJJwH6LfTI=
`protect END_PROTECTED
