`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4UkzXP+cuw2p2Z16aePdtGafGKxJQaAaJgn5DsNtUZcorT1n2AiC6smk2n5sKJ3M
IALixmygZxXhetEF5Y33x4cEgpGgiQXhDc8vpSwHZrRw2vWW2hKL+hMqAua5QUu0
WP5QowXRyCLv9EhxnZFBP3uZIwTIetm3BN832lTEr5WQvsqCAKYfPhtv25+IFe3P
76rTYH87zo4tS4JNFYsJzd/+9ajZzbIlN5+VhXASEd7laV2D2GrXF9FkP2/Zpycm
CYKA3fTzh8GU3zvStPoczA==
`protect END_PROTECTED
