`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PGnBRFmnHLRprFPstD3ygUjjA6TJnABxlZgAf1brGMlvx02NEXXU4Su3qwya8sjS
7vWWcBVGND2z53wjBnoPv4btmMK+q7VgLGKWHe33E7DRBC9k6wBk4M+gj/p9kLSi
5JuozeIQF/jUmczjT7d7dkp3cWPtmFRg2wL07BATWoGVaCyI0OZ75Lze2IjA17nm
GzW7PzaHYPHOqNhcYpLOoIq+n3lQMuisXEhJkYg2gM2EYbXpaic7AxQ2NNbGDsBF
MY4zolKHIYzOPO5Hk8aPOA==
`protect END_PROTECTED
