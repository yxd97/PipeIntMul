`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FJKu6Vjg51SElT7oD1y4Iu3+JJPe60JCNH2nvlu4VKTfSGE8Ei8UFi+FYumHIsLR
45H6bhV7F3/WgSwWFfa5SuMyH3s/1bNPbM/TFOiGtHLlokiUbTwAvyBUXI3k2MSo
91Rt9rxgjsfiz7c/4y0gsiq+tY3SSbqoXPMVcsv7govBM4+TvBDWhlB8Bbvk5oCx
o35tbjmshgSNlXmpjptNH7ys/pz77JKE8VANOfqqf8ZMJrugrcmWC1+cHvizky77
kkO2PE3JGu9RS8EJHxDJ0xd1xABxY667iYzbn7SjNhyCpva0CWlLr6U7IqWGuTZS
JQRAQoixzFB+lCwAIPKh9mGNeAQVgqsyCuyMCBs49fO8FRf/EAGTnjhArFj3nGrg
cOuz5KzAbJyw9oBJb8ASWvR4qtH7LI4A89+7HY5SZxA1P6W4l5x2cl/Mw4tS0v5s
Hk8yYRIBFutR7znAdnYBBKu+nOC5P8LtAzM3gXYFarU7WsOpXKLitHos3MDENTHZ
HoR+XiVOoET1xNuueT6MNq1djc9ln47PrvcVd6McYtU3pMHTq8Ym3b+Ws8Cn5PVQ
/JvZRkaB8aLrihi5hPeqtjqvQmVofoXh3wRFD1Wmsx3Ml0gdW8C1KF1KwCwGdoQN
wpDJACEbCBE3Ao55Fl9bnfLaISILQlVUPMLZlFxJXvBZ7NtbQSp+Az1FImCRvO2E
KPtzSj0AmS2D0vbEXACOxrrR2hksXFszzI7Pf6bYbBQ=
`protect END_PROTECTED
