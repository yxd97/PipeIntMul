`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tiKZ80RhG12H1m9Jlo9/mcphpFZIHGeMChdYDCgd2qcAfpv9v4SRYvQrca7IGzG5
NZxsPwzAp1U4npqOouLBv+mlYdOpt/GjhgWRm2bHIbmi2rh4PvBBb1/OOL6r52Jp
aYN9Y/8XB39Mlm+yicpCujVORyM5FaepCgQcDfvbWFVgQ50+dtShG1zI1j9732F4
UUVymErRla2kQaK/aQHNNZV/g6SXfC53Xnry/D2T1sNigKYLUZOt1M2qRVTf7Skw
2m90UjGcq1e/jwzLTCR1lNDhm/x3/BA1qXAcDshelYOl4IXa8uiLt/mo1g2lVVvz
ySKDCFxRPOhOTUSyvk/2EkFCLTMZUoy9Z7qvUnNQep0p/pkyvfqBvjZs9qjRo+N0
Ma0i0A7lsbU4DNmXbt3y+73zru5P69pk1ar01cDvBjiT9uN7APbG20J7n4WgpMFz
2/sRATL4lWxGZ3nMy/54NggCzm/o1/Ecx/Ai7/e57rPtdGFN6uP49JcG1zAP8PA1
RhS+a9GYEkjCEv3LMABT+iJhr2DKp9GrMq2pdAzAvc/aBxOAMCKxeLiZHpRK1jXE
0KeK8Qaez51iwjvLE8YWnWkdXYDeid5IYyZMyhBK/PbdOhqwPIBMiM9rvf1k4CfU
Ss60LfZgisQzSUgkk4nwtLvVBOxxuiAiTv9KIl21CDghI1KzA8ecr0BBHvdwlp+9
KqDBTZUS9uP3/cTpI6e1gRsayHRzplJtDX15y9f0AwUS5ZvhEmFPDhGLwAE/urHr
yYy0m56L7X99pnuG2Rl2Jj9VfNTvKjBfxe9r2LT/zddHiDwwy1LObESiynGtgFIi
ZBN/L73U4l9fUpYS4cFHaSXn5pNHCPbQm885BY+hmwOnQWVEzY5gxgVE16U7z+Kl
Z2q7wFiAhA7jHHAJhffpOpvkadFk7m3cVjJDdCUwui2b7WE74wjSjrKB4y6SmoQk
noaNdwJLDhy9VDTFRPG55B2KreOcoEpDQO0KGCPTh9vH8aySCRDg8LbGOPK4G/Bb
w77rwzm/kcGknxgrvut8U/BU+3oJ8OLxCRCK/g8qrGtyjzTtEf7vttkuvdE7k7Z7
NYz8uuNGj70noiTWRBnfNE3CppRJ6zWJGLjlOF+8jSW+qdzjoimV2WJ3Cyep7bK4
08oEc8iiC1VQI6Gs+3WwZBmBvcw2IDz+El03bH7s90IrfKe6U7og2mbiX8vLPcUF
DJIi1i6mnVLC9VDDO48UbvuVrAjWiOQhhxFn95Lww0YkddiuQcBguuOMswtwbRQ3
jJo4V10/V2+H/Ggl6j4cnecRPMDSg1WCd4ri+yi/yTrpF3t+Wi66TwcPlLr1XLoN
iMUr2xLn2C5Erw5LeJ9LB3HCMkQVpQJSxHdxOEsUWgbJx07L2XV2hEO92twwvPyj
vsMn7DoVJ1bVbdiDwnP/1FzStk8bnbqlbYIvv4+rIMnCMTpdsjv0UwKoW+ob3d5G
kNNR8p/7PcXV3ymqcmb0tRxuhMNRmGfuPwaFW9cSc+Wz3oP4UQFZlvoyi5/agrXu
L9LUJZKWSYkG5nuLM9dzcc8Jk2qQravmPS4xlvzOiRwRD2diJpb62gFCmTKo1Ug/
/epr62oEZIL0n8MZgDaz5wRSU8Dur4UbQFCcHXJiPEks4kuIHZxRNhE7cJ+UapvF
GwWLZq4hwL/9WhKTWEp1hew5iaiK0I7aBVZZSnwUYo6KfzH4AYERSbkonCNUluUV
Q8xr40VddAN+SBpgkLSt9R+ntL8SUOC8v4KiYj8kdcZuMxbEmN1DYEXfIpT62lys
rVGIvyeHMlsZQyTYGBjvkO4L4ITfZPv0HCWgRJpd0gkJLih65N28FZC46PhVAufB
CvUDMKTMDU9rq9/9LHvO4dOZ68KAmyWrodGS2N9PQvaBcNRtmJEVnYCErloGuN5g
CvIn405Tz4H+mj63Q0yfGxV+hxHRa8FUNJQ8RbZ1v+FRBDmHUPeh3dDSw7NVXk/r
gCQGGqLUfKvlw1q132Mvg5hN93ppulpzWxCBBeWv/na0HPxyeyYXDdBy+38vs/T4
6jHVkZKcCy3C/nKgHsY6HPnPYUeYFVA+hDnWzhmW4XTncScRBbhQPmpSB12qMEXo
NejHw2jfp+kbX+HQ1sM9MhfW9cJbcBGuYvWwAJqeFOCyFyXyrGGb+Q+x8AyViAfC
XC6GMZ+3FVwkMwquHYh2J7/i9yXbPYCWAQ5nWY3eGS7NEgzQdxVnP4/tAEMPW3NH
8rvKH0A5Dq40nNYhdGvS8VI1P5tQyByROkCZTYoQpWYlZ69GW1/SRL1qC8i2+zwX
XUMKV8QFhJo8hKNUGKj/f69TFYcyLiHudT4W04yor90wx4N6Xm5lSW1mYp9yBjOC
0R7Wf0LnRhQ8LBG9TvfrmBRW7v9BdY+brPzo0iE2i0uQJT7tHfFvcFDF4IDXB3Lo
HVXLUGt2XNveBrrEHftyKEa3WyS5QBf4WfMpYHylJqPWoLen16PnvYszMhWWngIH
oFrcHg+Y688hR0b0SqiuIMxf0sKQffW6e9gpX7bQG6i5yde7xKCvUweih3OByN4G
0GnQqDhwk3hvqNKzdwVVW+c6oApsuOXikwAVoDaddR3NrLQSwngWuzhrT8a+7ux0
WcxLW5GHLsAe+X5z6AQGycI74ytVHUPZsVo21n1pP4t7fJz8Me9x5vPOFhzjwWjp
Jgi1UU6dqoLVfXghR5GEPKa5b6Mcg8d4Gcq8enlcGBsbeabT9bn7UyT7WFiylNMi
fTIV2ZUzTVnJaE6lRvP9KQqYI1g83QnYimA0pcS9OOIwgIMfPa2QWX+OAxpRUo8S
37gUPCfXgRmsRsZxI5ugYB9/rHImdvg1S2x6m8Bt0fDSEmFo5lsHhwf/il3KSW8V
zy6g3ML8MYDDz2nU7mHsoeELqRyvbcOCLBNkEegthSkoeojSNmDFd0v9k1XXbO4b
80M+OFTmK8NbCZB82A8vfZJui2HYKt4XlOgx5IXssNzJyE11WEDjvosyJRzYcS2h
V8RAnLXEV1SABvTBMoOYA0TEBmvjkTDixFH4lf5KDH3IwRo++7V2OdY3LxxMSjw5
ZEZmNWm8T7MoOXv7lH8oszTRk35xOzjy/t+/zyiWGavTh5racYda+b0bTRtdxeA/
f5yN6xIJxfaSWou1R58ufMZrb2m/FjXkfnAuaJmlDWHHDKM1pXGwCn5sR+NCPjJE
g4pDistIw5o6xI4hwTSX6ahz9Rhx7kifyJGLtS137+yiRfi+Hsp3MhFy4MsfleKk
ATkw2Ow8wechOEtfm2sdSLJJLE6sxlCjn+1V7jeaVoPRSM0hWt2IJ+sEmbZA5pBy
N2z4VqyE2dhdGlt+sW4nN0tt+mOM/+phnVzgGIiR2oscbzSZRYoOnrXtiPMhVFzb
A4Ol0WbZwHkr8rwZ7kzO0fmgVkxjqVuKLHtWF35Fz013+yimSNoKETA7IR2GvU2v
lTTqtbr0W5C0Z63srNMeKVltK5cCsWewBHVo5W09aAnvYjVGUWqBM3hfiN9wA6D7
Ou/fonPEggPM7qh0R8tSR+uGL82dtn4Ig9GHlLWCEQLd3bez3K13/8lbL48dB93j
XGSUGoKyOV0041BZ7ZhrV22njmKweSjYSe1TherxB+NQmdUfTkRnnh0PZR6f8DRj
/3WDFXCCwpqhTrwMG2flaasRaxTcAFs5R5+xMiEDsspvqtI/LTQ4CuilLXwI+Nw2
NWIb667YT+IIiyGJv8oseDgozfq3p795ur0i4GNofTtBwS4nYRWLA16XhrLRkSYN
fHlGCYokNLwP49y7Bz6Ad5qKegmMIo6Bms5lb4E/WGzCB3ZrF3St8AYKHevVHPyq
Ma9xSIb9b5RXXs/TM4pTgUgyNJHFPFRd7ujFN63ydEDj7+UGcEBMLC01b8PudDj1
lF/6tQeoKQoWWv+liKNpgshmtAQanSWWbZ7DEPNoC93/gQiZMRpr4JMmwXsddLvz
3/VW03Q6A7LSNm7YUZZLQLM4aUXaXqUoDjtT27aT3t+9AtxoqA6sFE71S9pEb7RY
BIstXFpKREIjQJpbC3RiAf1OV3n6LpjqiQP53MrHvBUP0iNShcYZvcyiPtkMj7i6
G3eM+Zzatil3mcLymcMdVz7kycGY10sk62RQQ2L0hgtHC/RXwPQC+74aqPVqeMna
uUJP/NPCkSy5QRVFAmw2OyYSSnhenpJXVsC0QamqZD2WOVBLjEAqArN3pEZAr7I8
mk66elpzcHxISSE0RGA1TtjlePWKMygxHhp8ZATQFg7IR1MSDbrLzEoeGwOFYgvE
znqxBtCANQrHO3yYMVxl488+tgHsB2PhmnE2MNM4HnY7hqgaXzTlw/JfX9VSHeaq
D6eyw0FQDsBuvDZ2dEtwx81i+/p4ekdB24K1WRgf4+g6/5rE25mb7qaTSckC5F3P
50QID96RWFPzOGqXwmDO+vhGyc2Tb6s2K6+wVuHGTZivHCIh1KaQnmRDC8ZCJiii
P+IexDc3halaZUHyRYlSX6epI5DEIeLGHjxAAapNYJ+eO2rP3xOdymcSreijsJA/
VHn4JzhgbM+jNW7kyxYK3oNovfiUdVMHlgtiwEpG/cy5BI3pL1yxr6Uj5krKpvA9
y6+Wshs/axveEC87KHImtB51oiXoWoaPMCrAeddrtRZ94J+zcVQUGB5iuLPRdn9D
OXvP8XaBXXmBgJDwrnCSSgz8SqUugIccwMY7NDl0P/M4mH8PHYxAZ/pu/tlFaXf/
ipay1KyJiOc8rAAbA5dl4RxDwGRUnUw4XaxfHtK2ryNyA75eDD3hczYzrAF9GTYx
0jTFos/rrvBqePMUPaFgveA4Zy2oRzArDsalPS0tAa5xLITRclrgLVMNDNAjCvez
oSqxorn1p812zZ8E61grAghV9JnsAjb0Kg31oBkdB1U03BbimHuyCAGutSrSRjtb
YWFHGM0p6GX5/3APy6+17dpQJI43RaBV3MDI6pT+A3furIGaG0AhqcwcMP7qFOKZ
90msxpL3jzaAyxxZALI1Ui5v6bfgby3v0FRw3fXU3CI=
`protect END_PROTECTED
