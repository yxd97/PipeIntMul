`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dyw/bClUQ3pe5mzResU5z8vqfxHCvIjqQyzrebMUHq1hccjNlz8eb7VEoOkgOd01
YjI1JJVEnALbkEEoyWx/IxRrp7s42CFHDk83WdpdOMLbN4cI0IfgLyCqy0xMrZRT
Y16qfgTJXRpWGtC2vwzwOZ6IhEts8iU4oqcJkV/ZabODfDZsksiZIZF/Jn9ETAjT
7d7U7+y0JIgIiE35ysntAOfRqzFDwYi5e0pVpPK+4srdXxjued3y6zYpjPbn4z9S
aohbJPgozZGJh22d8q34XdMfNLfQxfw61PW4vPg7CI8QJACnmkP+y0oB2dJVhacD
eZGVBMbgNB2+Jp5E4m7a9+iOAgQp61npa5uRlvrXaJylz5TYuVMWTw1S4HcIU8U7
7vEKzBCnhijnP/+AAKTKzUN/VPP+2upsTDRppXsFoC1xzTeZR/5cz2OeYakyyFgy
T92sKrPSa4Ysnpkzpi3XW1x5fu7nefASu2SWPCkxGJS3cKpE06aumLG8bp1txThe
lXVaKV0QwchvAZCFSUVgGd44CMhbSXRBwVA0v79vZKedAI2Dr7tHWXt7U81fS0v4
YTn6MY8iom4F5G+9Muvuuod99nVN9DOEa8qzrwIE+xRsBOdgbVipT1e33LICC9UY
rnI/umtnu9Yf67SCJ+CoiXFb/Ir6t9J0F0Ipu+qpy3098tUoSrLLchPM/qvmp0bb
q/mexvTmLzashhKmjyFUukrRA9SFdELN11guzePO0dA=
`protect END_PROTECTED
