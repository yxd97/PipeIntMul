`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUR2SN0A5RjJzl9iagM58Q0amJwddB4B3LDQSXaqdY2WCoiv5zh9XlPsvtqFfgpg
AputFexBwZmZiaOW+Stprk50g0SB9KzGQhbIvm2wsF43TGqfg9/nmEgQysXUOx6k
v6t/PyFGw8IS9Ei+FkduweeJ/IT6GPYtAbNJq0J2041EGGAmd+R/wyEIopbv/b5v
QJiWWBhXe39iVSdxj7nSNBqbePM0Kp48gpbRIhlwW7N2MJg7WOqigCBbJB2nTUfQ
5Zftup8OPxjVio3/FFsA9qQAjcUtHe7oAkeDuG0XUNYRLjmC7b8cU4LMZ82OGSg9
FcenCnVodqUdTm4L8hIdipgvhnZm56V1WwXzIN1ZBcl3jA01C99O5QnSpXyn1cLs
jDiVbI1K0J091vf17B8jFYj/iVxvlQmnDoqNE7FqwbQCevOypU1rWZ2XGaZ57fA8
mAm1Y3bsdFlR1dITWQN84Ry/NbDq326ECUWJMzCDroPJ/l+2vW/zubWiHn7uD/22
P9MAqi33njNlQAOhxwbE+DoXUo8SDOMzM3cD8C0wvbh2m5dNDrXG8BfYr1NXDBT6
ilpnK/zT2tboCC0ThfMNzDDzHE50u3JKGM+aZDKJ+VlQupQnfyf1g31Ub1Jv/rgs
X7GGYMJCz4cQG4UKX2c3PvKm9s74MdPPtUHsmIw8jph17XkEpQ2iWyWgjUn9pU5T
8bzURRaHHLmLN9Y/gZhZw/xK1fz7/s/azGai55Qa6cAq/R4YNhrSEAPVnEmUL/7B
PQEppgkNxsC0aahqGWeJKSqI5MXp0cHFfgzmZjuBlxHqlHvngtNq96xX0d7Cz8MQ
pzOISV7horCy2lFg6KC59cth5CgW/gTJ9ZlBKBDTOUVB3zlHrXBJ2ii+2Z0JSAHY
DmvOu7vEJ0z3bqy4yUIO5w==
`protect END_PROTECTED
