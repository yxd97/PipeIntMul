`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tuS+pYVyXCbKAQRxnsEee5iC5//4kZS1Vg65c9VkdXFB0kVdLKIdP7YPd35veGOC
ZgT4p/19wGbkZsjgomRPrMF0vZ2Ka1B+fwRzTmaQJzW3FUvL5ILAMrCpsdQ87++E
4XSdUmrwACHydzG8ahaidwdGQPt/j39ZR75vFlA7jAhJit2T1NK1KsvlGbNdKdbj
9KAGJGzTVG+mF+VLWXwGl38gwYmfOJVR2p1X9hdrj2dMs4miwNgGBhUaXozBEJ+p
gCr3M2vvZE0nkkNsdw3VcQe8FrZC8GWl+WZv7xzYAlMs+JMZ4UARY8CGntM0eLC3
pOCVtCHapXxspk4VxJOcL5chuu7ZMb1mwjICvhVNaMaKhU9Luhe+FoahZVk0civh
b0kST3oc8HGPXUTAvgx2JOWKLdZIcExCNMeVoSlVOlkOkHkwWpY7jzYfVfNLHGqZ
9G842ATp627q2kmZUN4m3MhhRq14aQvbKWduoCQvQq4rVhEhc3aizCPgfJEmdx2S
`protect END_PROTECTED
