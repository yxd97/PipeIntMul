`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8x+BSG7xsVFawN2quXmr0l8QYqW2w6tvsikpqpvJ9Flp22Xtl+v60hj/sPzUxJm
od/4C51veNh2CHSOLrmfeMLffPTNeCnD0ch2Teg1GYfwI2dwMDpVjXVVMyQgiYSI
XPZLl7tCPPUqtFg7Yrw35GmBsyCauMBlSc6K94c5oehLWdYql2U6qx6Yb6DlOZ/I
Bn5KdXugP3lcW72TYfHKY3WEInYKjfv/oI838Fg1xdNxsEFoN9kuUqI0zWk6AHak
7nJljtCijAAwLmIVMizUe74VloMSaT/qvIAunaQabAM3jyAVDhIK3GQ1aVFKh1rU
tonYd64T9JXJBbobJurYeZvy8+CGiLTKuTcD94RlIMvKAmQyDx8/KThwEPEVO1/o
+VhUocvHLIMcJMfn2cqU6zckfKuiSrvPh/MnmbfG/QyauSbVcTolCsQr4F24og/D
yELvq0Y8OdjjRRmB36/F8SBJ14ajZ8192ENG9BA8RBHOj5Cw9j2IHbH+Y8n8lANB
Qxg8lwoZ8yqcdU4oSe7AHcsDuZGe4e2hqG8rca7SjOOx2EgaiI7vlVO5c4Jj09JT
nABmCeECsh0DbCgWOyKJ6emu1sYJkPcszziF8vwdXtXLhw2x8meAfGoU75qqDjFt
VmpFbHPYdsibiiYQ70xAe/3jfiBzNlZldYSvySdhkinjuSpY7BAGIOyAXO5A7L4Y
Ru91Nmw987fnVZRjGcyTa7VJpZoYW3z3dkgPbWuey44J9jZWAeQuKneKk+aY9Bzb
Gbkazqj08EAf7mtVGdCPPQcy3e8jigBoP9077eiEseneU5lLdLKVh4rOKt/MHRkr
FQCJ4yvjdhb28hA9zXVwdsi61WhLLBY/jf8AOXvLw+vclt3vmKWF+biqKCDvyMS2
0gsRzQcLDOHXB7b7VDLNRkgO/zQHe5s74ffvWLy+Pndq+syOZGlFOzdEShZH5aNH
6iIgBK63z4qOH5imxSvAEn79JU0nm1zyyKuy1eHlA3EVtIDqua7jahKkgu0ygw4T
m5KiQ7NUBOF4aStNBpP50Sx8AXdwf9XYwXQV58GwjhnEKTUqcSnRUENVhJsv7tt2
dhip+dQMhG54St0DhoF2ubmTgY6I45Eivw5xWnCyha+7DF/mKHJpW+QA8q/Z70Bw
v2iK9aB2VPbNDX4GmQ/4XHvU0pFUWjSceu6gfdcG4Dqy5CLBaIUkaO+BDPxyEeMs
LqTsZrnqIuwws1xUqhXrtNAm7/rnwta3aXRKpOaw0sT/Zn54CbwuAjFLSuY7cywT
pZnRlP6exYmREOZvVUAsL/feELmRxSF9tm4rV2WEv98R7jZr2htRzSUkPRL1ALVf
GdONJWW2JG7oyzL1PNR3byV8KG7DfYiqd1PTnqR5KvcMvscWiSuTMZRuhFajyxTR
iFG2YQId0lKGv2UjnKteJiXjDIuQM9P2ANXTYgFvIS5L3DCiYWuR9IJH9tM9ofJh
TZmST/4nys4gmqo7nJOJkxVhNYFpA0oHLDWJOawHJtux3sFkzPyxPviqBs1JVSPw
fko4BKreF+QezrhDMeNTL2YUpCIDOVCw4VMuG72fB0eP+Qi7RnKnFHhlBpKdTfIY
/ORM+kD/X4UkIjFz3JFsI9NFcPp9QBlV7ftaoUPkF0ZlrUVHfU+42qyHCVfTZrN2
c3pIAtUr3O6oMyIMupFAkc39LIW8UA6mOFDXp7BIv+DgE4ppygfpWWhmUZDeiBHV
8MiPyBGbA2COEbyH2SukWWv7McrUZx8YGleMLPhjBF8wSrn6c3IG1y1U/WJeSBGe
YnBudc+R10JjO+SsdgUPsqeXEyLzEmj7ZfV/+6MxYE5wvbZwICV5tVwmnOHFXAwK
CDz4vA/2NlhIJJNBcAePjnloAuDMWafcGPXJGn12kpYDWSy9u22f+NJWNmNnqcjz
kixYrsWnp+PzzllGLJf65R1yuoejHspqsbJmKLsPgeskWcHIGJ5Goy3j7TL+TNTH
2O4DZSFZXcxKsnk+2yRag1GoaJ/RXeYifYGJi5JCuGd25Gn2Lh0jhcIct3SQya4I
VgJ3vDZN7DNdZ8OJFXN56xvG4d+So40U02QygSSoqztilrE9pKQ629FDxRy0fjIl
eRXoJBWcag7zL6T36dUXnhE1N1eDzTWNHcxLEJWEqF4JuhN7w6mKTpRjXkZdnry5
oxnlpdPjkofg/OsQb08DEQzJon0h/DMCrh0zyHav9+HYVOKEY+vAtZqp7DK6uP5M
YhrjznW5D7eyvoaMgXHfQTckGd7/X8XUJyc4UD0hBiog0jF0yTN2pMmD6OHDgKDx
NMPT1tdyNJJldhrCwjI7YL3cZmuVdBcThSN2/s0QmsVgXTDCzW0RNir54cIsGo8j
CY56gPrXEy5PeUsSY4bsQ3whYHeb1oY2EiDWOCHwcw79R8d7mcE11B0t3jmL07W8
bq6SumndS+tmE11dmBHJDSjZCgKZw/TWweGCIqNLgAGjgeHRQWeoIiNQetT6sEOV
HZZXqC+iqFuFcjrT7nD2BuA2Ttih3bwo7OWqmsLGSWzbz8m3pFftBfaig9yRjVFM
1Hlt9zcBOrB4Dqrnw7tHcLwOvUmDLMvleBkQpI/aODj27uODoLP9neMtkIyDLV8i
s9L+/bJggLnxgzJnBNHuL2uOlVvx8VetKJsvIRtlj0K/ecbCnxIckPt+aWjygukB
wJeQ4cHH8o7SOXaPL9LknjEdffYfOmT1TwyBwfPJVLNmmrvO0fJKS5klQGv1eS75
rK2nHFrvFeMUzi8KZlX+O0X5dtTsT3jJgnZLkKvS7C5kviwuui1P7/gcW5prireD
a9NGgNLjIHNSyjlPVgnaQAk5D98vGluakWIBHzB7bCni2s0B3ECZ+5pdlcuE8S1c
/nisGsVz9pt5me36C3xTULuqz2blb4r6onRgRGMB1bdu+5OHiHus3e0d9Q0e0mzx
mVqTxXU2hrYslXUz6i4mwME5awAodcb3sq2njMSP8HzncLm+Mw/SwC726PjEVN4c
p7tHYEEVZurMydWBXoDbfLE0cPJioMxAddhypp7HCJpISzfSq1hY1QidBgIDXW/g
ejbLIquyyTaeYjZchVDJhP1RpTGcNqFgmnlN8SQg1WTrV1TnlsVgetFnEOqJWp18
nSm/DXb/3zNv2XaQjshD9xxjWvOZgZGB3nJfYOIe9vgDfPKJSH9aP29R8ZvB02bK
fr2vh2H1uv2tH8XlVaWGxsZeIArxNztjYNPaTLE8BkvnqN3xoxYT/qNP/UVxNaCp
M+ctjDHW2KTnFcrwzW6pbeByAHdr76ra66LU2Nfa7uWo73K95KAHsOb7DcMIj4IO
f3S7dmiPf1fYAp1u5Hi6hUedlK6VzN+x0vx1LXDBJH/QC4/tme24+tgCbFt8GoGD
NyEpbpVw2XCyO8ZNmPld3urtn66re2tWnqtAZCpdtgryZt/4PfL57L4pQMePh5lp
NRovBPhT/kqpFz8La8lm3YPsgwz+YZTm2+yCV3vXlqI2RTlfBkTvnhlqsKtQg3wm
bLqrnvyGQR/ZTiZ617a4mETR50T7rtB0KlzECbpkc7g8OHnhIUCHx8Hr4KEuqVz+
3ehITZrGDdDjx/rGXyqOya8HIzWsMdJ2hUYxv7aImksDazIxhOZAQsRD+0MZWVbB
BWNt7MWNfaGKICBQ2KgVDbkjIa40G3C7FM64TeEd1kkvAreV+oMW2tgepF9R0zMK
G6nPtJ4L9oEwJ4V+Hjf1zMwSQinaY36l96G/042RNmUr2GBFEuiE6YdOL0ocAsIA
SLegQsYGNfyGva7PZYUP9DCfLKCkZ8fGE61llMpdRh4823GvAl0K/YtLV54Dj4eM
C6d/vjW3obZPeUu6PmhthpFZv2IbBOWon/fqhABp2yr9ZZoQtFXURKVhwPPBa+nY
gE/0kQxS/qaDoi9pGB6xs6MbIiH6VuQw/VGeeBw5Eu9neA2JxhozDEu8ng2Bi9Yh
DWumeuCJVfcm5sPFV6g1C+aKQKbqNmBwgFqUJn2OUY10SQYnbk2PTdXeRj3DJu27
QnYL4yXY/LR/79YlRzvdp8sLnyubKgCCbTQbDpsESbjM3x61Q77LrIZG2WpPKvOV
v2K/Udmk7VBo8WuDnf8fSjH/5zbvNH6nCDSuYW58srFVTZf7+uoNfBpdJCOF19c/
Wpy9vFrtlF9qrA4yDyN80wDTTo/nnzGsNAh0GZdOUc+dZ6miT+oFDCgrgbrvW4xs
zIL5LwQa8oaQEIJCEan0YX178F99LGu1Z+fbJqzuqCqzYqGy+fHnP3f/zgOrIC12
rVzFyh8vDnCp9GCJ2alorz6IXee9sbCedM3ni5wZCKf7ZZhRpY7+G2ZtSg7eX9gb
koRj7XIIIr/zQdZ28LrCO/vwVkSv8Cc8ZOqN0DuUuxopDtTqyS82TAPVZwC+fWi5
rDblyb4p6cGL5KgMQhOEQE5/UNDmKBkkRqqUtFLhXTA8NkvDo9SVSIkoFgCrHZUq
f9wMMzzvyFEGBMvBnImHhpTY0+fJDhBG/qEc60MwhcAXHAsEYIwOQBiK54yDCWZq
M1o0/Wk9IO2pYwRlc4ypJ311RGJQBi7yorrLPW8FzHbswRYzjxOXA23mj12Rj73j
L0i4vh9j/8d9/JcU5WSovG4qC0NG8xfP5SSDepticbDMrWNsPB+zRam8nuojKoZj
XgPAAWqvg7M56ax4Z20588TXIQuYGOTaRug20OGsN8VMnutA+g4pPrYReS+iE4EG
IhWXG4AxbWxWyBX45fgImUD0yESNdc+ZxZA0SKKDqFO0ZT3ID/Aac7yB0iwbhaAK
oZ27ukGC1cpwJlkvni9cAaBw8BvNtyoPAPmIQ3RIMMlHKOXkm12qqhxi/dfTsHcj
FOfnzPEod9CpZQr3NtawMTA/DIpfQ2VcHUPQjgDAJsF+K+wfFt3/yHn0GnZiVpLx
1RVXQr4U+jmkLGDK7N2jYDKcKU+V9DE/+EG6YBrZElPRx3MnT/4oZDqQs+SVP0m1
5fVhxZRdY7q7r5hkTE++eIYWqwAESlMz0t0auxHdLv4ycYV5p0wVovw0YW4m1UzP
HcOBTFmGBpVEJDVzCYmvCve4aV2qB1GEBgDxx4mwj5zHNtMOpkJqqaRwfz5M6x3a
WyObr5K36yxH7NQQL+oPHpuaYrxXV/mG8AUc5sq1JNGj/NeScRczBSes2Bd5ALAO
em14fur0qqpmvI7JUinPuIDubAud5BAUMKOxu0Q1xiT+R68R2WCNMA+CXZ+i5ySv
ukTNzY4qIL/dhIw2dQglY+pbma3R5rDxPOl4AzzmbfUMG2Rn72oMvdEu/qZRDwQ2
F8t6OILgU6oETuVkE+tjpEP74vk7kz4mLRa5Sf76NrKMTNq3YZpM375ZO1J3ybRu
5Q+gFe/Yjxd/rYHVm+XAK6Z4nEpZ1AK5OJrhYfsRd0hDoqTYWEDrlZOedKVjWHSx
yScVo0Hb8zqdzWlvRvKqgzDaJ/om+AWaRAi0aUN/klnaNMCGFctCVhF9LQuPFBM5
m/NLBOrgg/CyzZaEIWv0hupaXulX9smoPZQOD+7kYnf0xdFYSnJh1slJQOOOYAKF
2MKEaneGDOAvguT+hTmots0PNETKgZbhyHg54YxNqHH67/mdbPor9IUcUK3Ka32p
Hn95VGJFO5KqE+spd1ctVYqlk607CCV52XNO3ebU+VGQnSuhUEcgr5qwpGzHtLpQ
HvLom9LJkdkzZHC7kXWpKXNhNIU/eYw+XQl1je8Gx0nlOgLm8oG9cRgIuAZzi+VS
MyKxK46MIp4o+09twOtWVhbFf976WqnifFIdo9pEl7y3fGojssVN8jbrt6cl3On1
Wb/e1cQdCiOSCXglHnFM4ftjhlJQxdi2XATkMFUuJwUc/JwkCB/sJwOUjhnM7Sg5
xl1P2WHseT6SFv/X0SGbb+6nXew3J3xk8AmhoyIHrRIX03xvAMQM7jx9xBq7iwtj
boM8YiIUUXPIbbi76g82qaTpe/hrliv3Zvq6PJ0S1gs+Lsk9DOtMRHPzYxq4lf/k
B8WGvoFqhlA93jFJpYpRTRDr3lt7ef+myQEq68Sh5DjBiGafsxO7zvaOvljj+k7n
hNKhbrq6+9Zrr5bOHoxVeKgtVlRp5yBMLohAkUGJTmxj0PbWo2vzPgdWPBwtmEu8
2dntwtW0K7aL8BA1YKA3Ib7px/83hvU20fCZ9ris895NvZZ6bWXAo9cNLFCUXzW5
E+1jOrs7da5KtJxdD+qatSuRkxW5cLrvNFs8x5W4rYhnb23f61PXHPXac9rCNTPM
UMtxEAUdwEREy5KZh/3eZ6vTHoG7smS8MCCmivlDZ/sNe1vO34eBOabAcaHVvwBf
TXvRyjWUfOgMeYXAA7ZyiTQ0EB/jJeEA/lw7elhPQUNJNmgb4e8vnM415MU0nej+
ayNxO+Z7hyOWDSvtzP2AT/xt6i+E9OCUbdQ7OzwSvGaR0ZbM7o+93tdk6/n9jfy1
v9ZhQiNcnDH+1Fyn2a/W/t8WYfm4qJ+Xq6Mc79/YTLcIOMU+0fFWef1I6yg2Owdl
hOKGbodw9bjjfQCIqVpSA3BqoDSne8lYW46TXiqmep7/LJOLR9rxNpN40TXQqmIS
M+jWzi75AsA0Ub0zJRqVWGF5aLn9sV6H2ax3MuYDbgz9KiygwqiwtmCs+zEu+UkD
S5TSKxzBersZ4m/pfCTsRHQ6O1IzLFbgM90qwlNLWOUx/4SqaiPBUdSLvOKoBycs
PNkIQjcbEpLJw75LkDdU0MfOKAnYNchzkN/e4zm7SAbtapQGqFiVjNoVcemvXdEG
c2AtUw32vmH3fjr329eBCKysT5BiQiAeNjZ90UCBKHh0sHo50Fz+eI8EGkL25LRR
3KUDEjcOQ7FiaKDHCIdCZDjeV5zTNn9onH9YeA4Z2zmKUzR2zHPEyimW2yLHkHKm
7xinnthsBQpqatdMUjI6O2jBjQNLPe2xLad4TwmFELL4+R8m36ekkrOdLiqSTAHI
a7QqFEPPPe4jG50gKqMXZbzJjVVA/zJgrnIYll0rGYI1mvpjHJX9Em0B/QXu8t9J
vyEmg5FH5iNOzOy32M8DRQhqT7P/QVC/FhTSeV8KJ38C8S6Kb9Sefjm1i+3FWr5u
86qJ/3liHkktwWUITSXbBavTq0KzVRe6053kPwlTZBn/3npXIZTbO+C2hNV7hAzA
Zt9lLDF21JCgvFH8SVoVocT6oB6WTrLGzaHDFRDCpxWmuDApdRnINnw6GAlZEsHU
kY68oLwyJfCb/zkA/290SA/QnWDLLBbPNvINbsAa7QXYrzTLQ6BHQ7iDauSipy3S
aU3pHddIk2ThBszMbopwYSRukEJE3qtqNCSHDA7eUWigR4Ev3LA43fl+HMYR9hcJ
waM1AsHmqNX5GzYKEb91mL2yH1VsnOuSo8AHujiq/YmHsfXD/KBrOTsJblnjkRu0
xzZzsdkp3P1AOzjt9GqE0CReNCh9i8pCfQPnLqAcX8ng3vWmgbhoRYKd3IRQHgPg
GyneGIE9oRI3gnIWmYgpv8JKkRkaS+Y/0JZF9CVZdZBLVuzNXdP5IgUp16HV4Cjk
QHgFwsNY37cmVyWH9NZyofKrEGA3grsykN/CNkjOtCMlgWJNbdV8ggcl19WGiIJG
rJWMA8myZ90kCEUvQEtjtsbY4zPLfpziBafqHgzPyCaVWLclRykGPoRG/KVMHf2+
XHM/pD0O1g1ameXcIp1fUGGVoY2b8ykOnB1QB8xudyR9WlZs7Cxe4aF698VclJE4
UFcDTcz9RiV7rI3uJEjuQn2uHKFXTJ1atYZJFKNl3X7cxayWuaezHEpxx1X/ateG
i7tHWs18JUDZsCPWWviXMmseOyDMPsKLd98nLRfltG5pAb3Rq6L9vAYvRPVGs1OK
WOrBshqqwDPbGSIrMTMEAkUqvp3w1Bt9VbZ3cZEtq/PYGdveinbW38204OvUJGhb
sicXUf2gnC6AEc5WOP/CUnQ3Y25PzRLrno+Vssuju4haKB82FZ8+KUWXxhhw1Nmg
uSuQxNlXzkZY7RngsJcnW8NuWXgm/zcjvp9mAbGLP0Li3ucxfP+kUURcFqKkRyxs
BIwjtTDbhp4FL02r4QFg2EdjTIsLrM26DfFyUgefFfKU9SLrRxnPx6AwTQA1nvP3
TbHn82ZOi/QOB9KJpGaYlUjGDaDY8FXXgJVTfN9Uayb1Gh72yHdSYMmSl2r3TE0B
gV/Ffa13qIJBp+BsW03lhs7uZpISLqlUVJR6B4th1a+eeU6YdGSWuVFGBDHr1O+6
By2NLqwrTq2DfTuGqSCFLSYCJKdQJz/8ZSP5rAtMQjzlUrsEVkYJk1jnVnbZUFGx
3THq7ejcVwVrJApZIOkKE1ieofWicogmvUv4o15tfyNckXM+uLCVLzK0PCBwYjYg
TEMhuPqRu+9diRlYhY5775OGXb7Zn0pBCkh84qdLmv0LCPjm06abZFiTBmjxo7sU
FnTB3LHVRI+SsNSCg3vRU7kpUt+ix9xKp5ovFOPHdNkH8wBBWL/qYp8UaBsugDE+
mg9E/x6qgHhP+Dz6ZalR0lo8nfwuiUBno69+vpg0QrEqhA4hizgWZ0+GtkNHtGZ3
OqDCo7N2YuLvNIud5U3g8R1UXqXT8fVykBTn3vtCpGdlT1yynYNQJoE4NALHxFuK
ILE95MzpqbeSeLVycxiDrd83BZ+G1adq5YIyjyOuiNSQAcHRMyZ+8B796Yvi2L5V
q5RNj+iaHbfWJ9CH0yVA7qg8GFf4QzF2DrQQCkwRj4q1hleIFHZkxxBLQdc0YMnA
pwyUC5/yn5orERFz8ahbZ2ua86xqru7jJOBUSTK0v6KOjXeA0wg7/f1gvxWhlbSJ
psvUhEWGCu5DZHzlUnly/xKrRA/0Se2mLLV7S3xj9K2F82NKwdz3HWhoCUShJZ1R
ge7wl6z2FYT+dEI4atQSRNxaN0Vh3tgdLGZDy0+rXqaox1jeCLVZrluNE5U7mw0t
y88vJp788msYzIvQwjR4L9ImUCoGh/mcm9clElcnJ+BP+kRqN5DxqoxX9HPHEh84
vqaNEdUtwKognoxApB+tyjhXv9h82LF0OMjBG7VKSxZBVw9nnPpKQBCdx3MFdELj
ygzwMagyhSkgibGnVONSj3LHJYi2cPT5LaAb6djNVMm3wWcWeFZfKIMrKVRP4Z3N
UDQoaS4I4HcBOfzg1v5XeOKftwg6CAzDm0r+yHsfZmaMvbR2YeeVh3uR9kzH2iGr
74Xuuqi3qNTMuq63nJfUaoIS9n0mfsi9slmA+1lcIqaoZmLyXKRdLRLKs+QRwmc9
oTf9AL0IwuboF0mixllqMcUr0u0rzvQ5DxTf7aOO499QxMrS4Ad7otKzIbTNhoyL
NLkBxfZtPk+bJ9Ri4ILy8BJvi/iMgQtxRdqB65frjbTnhCQX7vYCG+QJj+HeXPG3
eHNQ6e7Zfroh4AhJP5gwE4TiPTxrENLQkmU+FeZXUJVlHLH/dHHfwA8F7uWYVyO1
Uq86LDWQV2DuLjVBkJz80H6ZHYlXIQJ7k3AwJdkUmvK14YnADTeewon2byL2/zeg
mNCAb3b4cM87Gj3wZuFynPad/pnMu9DGGQgeV8Bdf4Hy3tYVeKmKmu21XC1vFUg+
60yS/bjJ2pWWIT3Cr/CR6UUDBjYrYTjghjwnidqWZ8LJvfBO5cMXj248YnzNdlTi
Jmk0VrjvOW+AJOCzEAZS/Qf8JIZaq3e+aasBcDygfaIuBAd7u+pZQNitgiWIZQiS
jnGCG3DJ7JWceZV+CWHt1kUONgAjPkEHC7us3gmJzCE01Om0J0kybfBJEvrWo58p
RS3gh5os0HpnL9PMBHR2BaEnqKdIHkIOOmD5Guv3SQkkhiLUc5Yar0In9zziKvZH
lDdBQ6zky86un79Xo7v8YATkXv3KW57ltOMVBnhjfSJPqqaASRkHsn/CHoY7QhvQ
o+z4eG1M6+v1a4nZQ98ZryyQnH8uZ34wT1lkd7JhXc/fF2b2ek1TsZS5V1ch4oBL
ljWXlmwAnH8fBjHgC3egMmTHYYH/bsLWqmBy3iEzGYxg1J17FbEQhufsvqSCTQo5
p8TGdyQYXCpvmL236hug5Izkpf4UIIP1XTNVQ2XkLiNMoRAxdxK9pdJ0rYwg1bcp
poVDIQIop8KKguTto92er7v2JqDFNJ8THswRrA3HINyqQp6CStV2o21u/0rxwwJa
504ri6aklVxgYJyRN8iRQpFG2PJdgPUZvi21Z5FxDGhTWiu8kvZs3TJFw48NW+7s
vrmYor43kUOSz1qOxOJ0OcdfdcM5fgaZ+9Vjj/0iR+BLG9R9V9GA+FGj/tozTRqk
sDnMWXamvIFrJ2JPxEQWXJoMt9uEtAuHHuPm5uovhYZmss8J8zhDti26llAoiqi/
h0h/NG8z3oa6dVH5Fk7BKP/mdLE9pg9hEwQ+2aWltmiERaqsgUuPIbVfFhAHbUwp
rNfhVzaz9nWXJoIT3+cRVjnNRQ1TI3RfiEPUuXvWymn7+PJ23P61VLyWBg/+UyPr
5md8VEawhqqmALKvabzhqj1dgszsmFbGtft/JXqx9EpMVZptTmNetb9quHULzJc0
l1KVsnMiu59WyZuQPpvlb7UP01NylKRyRFOiKXt02aSI4t5adZyukSdKgW0OnPvo
dN2v9gNe1outOzAL70nIisPidAgp1tN02UgWLlsAMGe06gOBkux6h6G8RCxYNHlK
XuBa3Lqcw8jA9I0Krrw1BgUgVAT4mZnc6nLfxbmR0Bo2AfgtgYtk97YekMi6CWSa
Wh0zMgvR/JnKN9GB+0DSvajL29tohjQzA8vu/vqjjGadJY/0/YBzVJSMqqNTRHk4
JADzDrWDl71jLtOrHt5RpydUH/FxmKnlTWxDGKEHc2ZJIph255nF81EaBch3CmRv
N4VqZNChCUqMvKTKGkz6BhykMlV+Knb9DMzLIibTwfuK8cGxORynZJK27M+xsHTt
rH4XGdDGJwmEC6/MN3waa1EVgvM2nHO6LIf4C/z51NNPXZEmB1rkNTuQdRN1ofee
gkjhot6gMKkXpC6oanHca6UD3K8lEkWUi7fPfCvtX9f2fI4Frl023elDl+8R/NyX
cGj3vpie/9u/Jk2TDzwPF5VSk1PTvEXA/1IAIO+ivmyVtX5vA6pAMUwevbBoJu+F
QtdPLUbKSkyw1gVmD7ED7zrpYay2iU69R4L6qyruJG+95ZVZm1870J0qX1FNUIXP
M2+4gLa8VZprUyGu02y2taA8o3kmDORwdBgCs+vZ+bCKnwdjvYCUbwMseRZ1U/ea
bYsu9sqFjXIRPKrrc/yJOjWYKPYPrCuFp9ZzFsUVuCjuaSqeYreJscC2SKRpc1QC
IKNtTVcML4Y16VGUiKS1unavRpdzTZB2DaR9foFnG5AYZpVpbXmTubU4EKScMTbZ
lp6zj55rYcvTCQsksV3fDmW+d6ssoe5iiCrU4vRrPws8UwfeqbnsGN0EpYO365PY
pTyd9HaN+XLJB8PV/QNY6FSXFt4RRkNKNZD0aldL90XUxJlky4e+Q4IvnzuozB+1
voxB2bdRxgALhRXwotuWtOcWGg4Vn3Xbb3+X/NS6WhUeVX52dTACAADguxC1uAil
Orx8/tgjhsYh7yRpbdTZb6FvBv2qBL/TRXdC2yRuceH/nClFb4ntCjvbDYDm+Ol9
1c+X/WgoNiBKWzAo2bE0gjoOwcEzs5mtigy/Q8ETiILEhAYbek7Jjf4a3Lh2ccAk
Vlhd5ZgPKDK1koDIOnjWxF8Uz2hO68me8xL5hO5kkLfLpovZ5tBHOSnKSkV7M1/q
Hqax7uA386M3NAAaCFZCPFbc8r6YG3zgwGJP8Pql8N3czDFxg2UzIbJlUovatWyP
ogyBZlFKP7vfk+jlY75/UHy9KgfLvHiWxcxAEjtR3Y36Oscv1IbJX1fteTjK96rk
Xzq2nnuOFLfI+Xx80bYM+utFTPCiLm4cmd/iV5q/fuPdpeucs4ErO12vWJuQUths
138kHaFdGnC0GbZi+dCP6fMjmAB3wNIbYLhqjbrSzbsDbwrXsGPWFAc2Bcs66cdu
efSmrXpKxOCGw0ljMjOrwNcAOXD013/vNWyvl8+x/JnV/k+nrNDtveRRnG3H62pD
mC+wlp9i34lw2ng1y2sBnQBCNcaQqDZGhmOmMqkjj6ogMys04yFKopQqqYtC+LOd
RBawIMc+TR8DZw4QRnNjq1dmMXTEal9dGw+mQf9hfCT+ft8sbVdkyum9bYoixq5M
utxRzAS+gM1stL84EnFdCPMZ124niLETjmR53GhjfOykk0QzCrzksUWst4lThGDb
GjH8Mmsc+9dzprsQGfhR5oMtt76d+rojiPaYVHoiKfRtrW8VTWbncGEvt+bTu9Yy
l+lGB/IdGco0HJpU5EUP/93s+FD5jNHBva0lSKQ22M//gRjkA84GIYb1Vc4E/JEy
qyEdNurpTIvqSfJdmhu9C9y8KC4oAYkH1AYz+8/1HNK+m5NuTnWByAstVQtQ/En+
Fgz1uhuqFABKb4JNZhRZwf3IFNBHJFtmocL1oFJYBWj12/ksAwRFrg38RwYe5Xjc
eOBDqopC1ydOXXQFkzTCaQDD2RHKHPMh0N3pyE6lGeaorVYFUankFU35hYyP5nHx
btaGiWTMB3Qswtr1x9RMTO5iCXMW8ALz5U+NFmorFoQcYvJJzb9DgadiA7IBiR2/
qJdL51/YnN+kwVtRYDsHogOnnstloJ2zpngbqODHvALLjMPIKm74bV30GgBamy43
fwQ1UAJhWxmbtSQRF8/6/s3tnHvqYzNARQa1qY2eVFUjgdCUARWWN19yKLSevTOH
jnZz6YhVl459dzvtaYs0OTFjIsSep4FLh0flOpK+8+TAKRnWmBPioDCsn+Qpgbtx
rp+veu7BlQQbEGGMYSFPQpAC71Dfct0fiCz07YZNznsCE8dlVLIv1jA91usXV5u6
JCqqrqLSwyKatX8XSd+ErWyeLvJ/c31ycutuR4dbQloIyb0ILsP99+s1N8hHSIRt
93josv1xRpVkqX+EZ6rWF4LGxCuhWpfgEEKBbw1Wlc41G4zPfqzcwHVw+cKygZAg
yO3mY7Sn6o2jagyNlG6eyivsth5XvaLzmwaUWGL23SJppi30fnHDqZTKxq1o6KDZ
0KsAo1ObQvGjPhvb8PMXwJJWGFEZb/kns6CEDxDU7V4n8obwYsIJ+BVUlJYl00kA
49DdWRQICThgCD+Z2Lx2jdDIYbbK1Yldfj+2OJEIY1eWgW45IdxGSsThcASQxs7W
wNdu1NHw3q8J0yvFdKWnuyFAUN9rezfH2VH30GeiuRhtfUdn0LWKUeASPVVLUvoL
ixowqSqTBkca4qE+R7gbVUo/42LZPbLPE+3qx4Iy4PIT+axSbq7x0ZnFjxBD6BZu
f36VYj+iw6ZlYGou99gaw16jf84dQbdLmXHoLYrkRrbBz5YhnLi+yrI+UEdFycbj
0bqdH01QeJKJaZC/XY/ByBtshSyuwoEdnd4kCJVQ/Gw/24hAKofQrWMs1guP/RSj
xGs4VCcIU9ltkH7N7k7y37AyLcsP5P7GxDhAE6gAl/CYN+3a6OWlqesV+FcUzemf
5TcQi3plN/O3en24s4ljLJWEimom8+RKOtN87apwrvaf0hCbWT6KF+k4otSsCqxq
oJ3WKAVt2pS1aoOv9WOokPMSIpN6ldBzrGibO4ZPKo+bHeCARxf9iNnRIwYdkV7R
KCxf3Jnr6bGOpSyr/xbMBweGuZanj7fGypSAtu/2z9KB9bJ0R3proujWv8IqEvpB
4sL3KEv9IXvNlp2Yz9cLDCzK/YnEyNIwDvLjAi5s0INr0cgXBp+vHXdFuV4NizWX
tLMXwzJqMBvRSaGADrQwzk1hGF2dCQRMRx955DbsZz7LO0MXwUhmVaSXVnyxCdcV
3y+uHtpz/uPHsMvzELRUvt2smtVgB5RMEIQ5z5FfGsctCTh09ofkHYfFIBFcIV6M
yT5i2RZOICLYJfY95Y0WAweeex6zpI75OqF8PWcskB8jvGHYW+5ua5cPxETW5tUs
fUzHg6sJqD6e6tf3SWbShP919rL7bcKTIXkYd1zAVgzelifluuHEn2yvzIP+apN5
T2EmixnMWFY8IrHkSd8oY4vkjhrymG7t6iA3grkyltsXoeGUNSnqpC4ItM3HvFNh
9PwaOZeW63sFBvyV1kh/v4ISqajhZjKiuYhbRVA8uD2FRvQYplwr0W4rUaJBJ338
`protect END_PROTECTED
