`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FiITmnKpmIAQzv8JyI2GE/bmSZpE8O8Eg5mzJ4k5EmVPTVK48h6k2UUQ+7KiG3HU
qgX4WKJbt4qiANDtcwr2hhSQQ4AaL/MZkgwmuABDkdGiKExoa6otzmuvI6x3B96Z
z0wpvjqWBYKSUHPVjpCqewff7CjQbUtNfnyYgpZaTtxOZr1qQJIue1cQK7mAHBD6
e8nGC6i+ZGH3LOKDr35GVT++PG9NuavOk+U1advjzZpDYh4vpMHJZ7v1grSr5ZVc
fLWi6SBH1cz9pqocWGPOQNPlEYhfQO+H9ii3HadMcran8N8qTACLBfaM629r1bbB
jiaI2XoaQKwnvwFnQcg9FKbH19oNq9Kp8f6+aS2cZoWjOkd9HrDR+RB049GrKz86
uXoN+GHRpdrKiA1mdUg+pmbJXNgF07vnajpnahDTvs+yk+b/gBT7yrDPVULrfGsC
onCdaNKXHLd2+knyfE5abvExxHAOMhwYYNCLeO0syXv1o46bBb6MAAlPAnpJuH7x
9p4AE7/HOzzVbZ0VGXTpXgOacvM0RBa4eY1lzPPHtPRb8pnq8a19LSqlSZPYV3J6
r0vhOxEzoUDYNyhcGZT3EiTd0KnoLNTfquOEetCM7JCJAtxF0WZaMb2S9Oj2LW/q
QCCu1GTl4CjSp6KssDAMew==
`protect END_PROTECTED
