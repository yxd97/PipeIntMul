`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oBkL7EWvxZDbXU5PEd2kF/u3LhOcmEVGTuCqi36Z2wkm0Kp1XuHa1crseLImXLNn
s4sL8+qWc9KvXh91MTcg3wH2ldj3RFSO3rC5MBnDZF5smFGJG++lL5t0fZmAySlI
gHzqJJ9E7HHyE1cE8xIu2GN5JPynfBIDPHK+38aSrfmhQ/qr7lMNVasqffG81O0I
mKxrmzSpNT47a92DV38OKsifPhLOHkQGnQ6YMukhuPHi/wSuL6wnDHGaDM0qlnZ9
M1QUARFbfB9LnzvHdGx45YS9MeBUF30q+WfffdufAg7qbvWx32q1VkrwrpVzw5sM
SkfhA/6KUojsyt3amZLIjXRUkPLSTrMWWpGW1GqkQJ4cTyyR5a1n9fphYUgGOUXf
Rc9UZUc2BI+SEfCX3c7TbItgLEhmPF/+3u4y8Zf2PywqOUOOx46rMDjJEXH2I8yE
MTPE1cSTBCsxkTBymwo4Zq328fpYcHclHsEQY+eYsh+x8xQACeNTE230tkf55kQA
XxUmP21WVI1tg07Z0nAUK290DJnZbqoLjV06kW/hFrMLg/YaHUu3+U1jfDO3Sdit
GVeRo4WFS6qma690JCUvqjx2op/Hzhpeif3n9z0R/PzODVshqvlC7hdEyu9p5Sb3
rRC1oXbzRtr2HX29JSH8SmE/I51wD/cyjIxq+HQx2wVT1W+3uG+76ox1yy1pThWh
lNMTvzr3x3ufLN7b0kyx6H2lJucshOd9RFRut1wQTs6LOEb0BL9TuxXrmqyywcQn
HI2rYGWmIWbPRJFx+up3nQhojPM5ozHE5P4K31FWC9rN2ZveMZG2zG1BTSWOTC94
YSBsB09QG44okFnmPFNfCo83wYFBgjegG1VmZw5tybo1Yp1Ozev+TcclkxBjUwDH
WEMTZJIxskpXjN/6a0blYqhvCrQWUFChdqZh5JIHByOMjIVe9Kc1UNYSOAccLEi4
Qd7a9cdbpVBQy3GUnQKcgWeci5kT3NVx18clZp15HiOCOIcBpDSTNnsDkFKQ3gDX
qrDbI7LKCG3y0Zv2Qboc31vcn1q9JWr8jxdKzeRPaxXxIy9EOQIaZ96i3F4VMfwW
XMvGXDhGOfvWjKO/grtpKPUfuHZb5E4yAUsjTT/a+DGYfELIYarLK+XwL8lV+/Ky
licrHGNR5sCnXO/I7CFYz9BkjemlzQLmk9cKJpQLpbirHhl3bTAGvWm4NDPi1KW8
FxQC+I+wohqQloXTQePP+3YwCJg30uuaFay4XGynO3NLS5AHr1MMeOzv1xU1FVZ8
qfWx3hrIHKY3DoTbG7/grat4CLgthh8PSRTt9UPtZsbvjdytTBtX2DTmQ/ZN2Q+H
EZk+DWKfqd/k3hWkS/QGT59qGXemB/FojeMLr2Px53Oqi8cZHBbJvhP2Oooy/FwS
vRZ3VBDKege5FUEf9OUIYqgP49f1RfOzYgwBzBLHRT82WTSGvRfbf6HZ7bZ+KE8y
G3wmgZYWVrzRg3NDpW4NWyomgM68N+TTBQlbkm9uGtJW4LmlxvFrlhycx50vp4I0
X9NAhZE3ZmrEUFpdqAqplb+4tCMuzkNr4B3DkrZNj+22A/o9j0k55EqOsvAHnla3
fpKuyaBJFB8Ioq5OyXXd3K+JJxDWGJthP+PiHQ4dYDqAoUL2FCkJ6lsI4Cy2HC1+
T+pSSEmeJomCQABtaUT0uNsrDHIvzU3ER1CPgL/cLJFtYmlCHPF7QA8e0ULvsSHS
cv5aje2WNiMs+UR3cz4pXQ3ab7NU1/6AbywC7w+LBvTAnA/fyzgsJdbYzZp4eSMn
hy3RCnMyRozxdor+vDZoBMOZsc5FggiveceyAIR0xz31HbrPGmFEtW15O5/Kmswm
9JSbBBYvjV9RDaHEATOv71h0tenFJIolTm2vhXAEbKBwbXdJ52AnN7J9gwKXppPh
`protect END_PROTECTED
