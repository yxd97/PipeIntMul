`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lcfOmntU2N4oKQoH7Zf4GnVrXLXfFaMJtmSi/JsI6TfdoBxI8UqjY5MskCWVhYpz
I2JWXvNfs/J9Q/waYoupu17+XgCOMiqk0TA5Cf9mfgb9jcbMYCHW0Imfmk8sERkl
DQiPPnjmEhQwl+Mw0zNcQgY9cV94NAT9GfZXvxn00o7PB+F3mq9LfCVHi9u9D9VL
dKUzBqtZ8fBur0Dexe325Cuxn8Z4mLTfOuzCxNQII0oj4zEuK1rp4icpaTfFFRg1
CuEsCNiFSSDPbjHzRGVBe7Z25P37nT4vLSoq95zHXPWSFQX5agNHh/ODR/qCwzmg
6ltdBKnok2GEbxw7nk6LqG4LPLXETQBKQb0zeMiwiF4VpWJrZwx1tBKLDczVg3bX
r14GYIw06ZphIeh8UnwQumEtvnMgW9p+GRvYgakar4HKO2dcXyiMNW2LHPk5Ie7G
`protect END_PROTECTED
