`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EKhrLtTP0tm8W7dmaupVGnoGR+nhy0QwZY2zhvIDPEZbTIbb6qukDYYqL6VnS3qe
Vwu7wcbWbKPLdwD/XrxZRTZOGNLokk+a5gKDADo4kpOEMyfQaHC/2Y6yeat5M24S
0wmTuFqIzVSn4rbB0+ykaXX10otTs0LOcd8zHvu6UOKmvn3XHTuVif1xw6K2iomS
fNsi6kjQ8bVFq9UQpZRoxsJ/dRvDynqBPwA/coXVpDqTEkgEHu0LpG28nnhnpJ5s
21+Y1KOWVTKOTYtu5VS+dX3PLo5JiuUfj2AzzNAITF34IviVbdyfQBSeh9qkZ2kI
fHRFL2IouQIFa6EnsHlbMfIKviqeXl+IYDXWGouivVaKGdWoDramKmPgkewWg5fz
aPygRpi5yxgIGs7UKJ5M5Rpp2VTZd2C715HNJ6I0CwB89s8GH/HYpKJEjl6Ps0Ek
eSH5fKvnJqkeX0LRxyiJ0fZbD7t7rCJLLXAJSU7Tqg7PyJvH3EwHEJfWQHqdkrmt
VPD9qJ9go7gjuCO0jiW82rKBJ5LuLwJMIgHy3VMME7czfpIvcyvTkwT7rYZvOYtb
`protect END_PROTECTED
