`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2u1+R6N7Ez6WbykDUQI9xM7UYx7L/RHAM5ARmZUTkT92Tczo5QvlMFrp4IbsJ6T
WQ2ox3nxH1l1enLtuFzSVSPYJ9ZAbb7JNiOb9gCxmBs3gD/QEKyddQ6d5fwWGKj2
TOdmHhb3kkU/3S+yVX3Q1/WcSwrBGF41yEEoS3+XXJ5d4cURCDjyZb++27p+vL4F
OsV21HOgU6CHKf7DPn6HoAVgEsAIRihdps8HlgyQEdATxAO0L2sThSDCsY7AnDnk
g3U/ooIN1U6aAZqhQNLnR4Xo9zyDvku8ZcHOYfM/o4iSBWF4Hujp3rMvHmWk93+U
L+w2MjiKayIGOdys73PFFA==
`protect END_PROTECTED
