`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n+5rWdKIPXXLaDFYfd37PJ5DkNbhtUfuVveWqKwW6w5kAhnqxRulVYve7XU25OVE
I+VEIp5bIjAffRwDddMNDPLSLLEx6k5/qP4z7dajIGBaQTk5bLdo8MtStmRXUv/Q
DzJpZ7FqX/UCB1d3tL+KPJgqhcc89Xt1B0Cr2bv8/69QP5LVxVZHvNu+MclI6XMP
cb9dojr0Vn4SLQlSy0ZDWIhsjw+J4SQDQGayDdGgIyI4ufzsjkWbA19XlLIjHF2i
Z5r/7mG/I5fuOgvtVmQTagI9pdE2by2QLd4PosRAjIBRqRFuI8tDYcesDRo9KOU/
k0WNKwX7QHbQGwQSbB+O7juL8xY2gvOlMfx7lZiYOtAnk1orIMwGhLmQAnOcukpN
fI2o+IpRezuGRu259G1F9XSyYPPiw4XoD7NF2eKtb+zTWA2Sy9s7Kopr44bOi4ZV
gHudCqqv+7ONIMeJfDwUs5JHyeM8tEn3Zrxlv9HHpMVac9eBrS1ahmW1KpiEMt92
lBVyskuUi2NLcPZDZQ+UNfG5AMWx/Q68j459c3FhFrmPnOclK6sOyEClh5tzG8yV
adbdG5I72axGwkgfY84PTw==
`protect END_PROTECTED
