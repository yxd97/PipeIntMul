`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nYodpbN5APMl99EHS1mTA+i20PzyRBtKk5wqfsECiolHAVRgN1+7HtSqDpHYDwHi
RtQZv8vTIcfwwi0h3jPTjFCp5JKFNJxJpdCKSIj+CjSanIz9mgYjtgWKeJwUO2z2
YxItJLPot7ghWuMUMgnY1ClmGgv9Gh3yhppSa4REdsk+kj3QzTArXy2L9fu0Ygl2
jFJP1TAfB8hJcnvmY2hpElKCxVFmzlpk3J0dsjr0rBw4QjIDbF5EIrL4lDFIBN7f
7asZNVoiEplkidLtVsXS5CuNSMioQIU1AlymXxcpo8ZGX5pDd0wZ3ha+oher4zvO
`protect END_PROTECTED
