`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jjX7gJ2wayjeR1TBOU5Pm8xWN4iBvI5rP8SGa2UByILBdlCSM9epZdMjvXYcV4Hg
09Tc+7LRqQbHWVvLAuz529YoTzmvC7kCK5sFuXDDHPDMrfdmhT9snc5t9Bd3PeMI
yDcL7kXyCZjYsCeP80oRhzR7kwxe1+/XdJ8HjmQonI+mxrtIHO8c8c3kl48cDPwz
57EDTmTvX8FUn01cNHJh1Vs/+zeq803f0UXfogVbCZKMyqxllUpWVhZPiiCR7kQR
lnoaqVCIM8p1bPp+tBKM/L6c94lex0IGEm8ShFLOU2a02wOVzWbD/lft00elb7oy
Ya0Ohdn1ZOubKYASN46syijewJ8gVPniDpnFjx1Yo1t94Hk/HJq9DbRI4OfdwmiZ
`protect END_PROTECTED
