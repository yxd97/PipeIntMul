`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qi4Dwc1lzYyk/Qtsayr4OaUaizjjymtw30u0nCFTVzPuOw+4wIaj7d9y2AN6DZyK
P3arQQKK8/Y2rpM45TY56Ruc+GBXIJ3ucn3j74xQ+RHF+DqqonoPT8hjJR21wSUl
0YjN8kpSFOyc7/ZH4kf8EWYACT/uyspZM7dN6h6xwaMVWXft+leT69zMZKjXc2uL
P+XeVaZzaF0ApQKQUlpxMIWJCNyg2c9h1lVI/LtGKLh1YkE0Nk3ZQntqLW2N8Uan
JyGFFeqS/AlV/42OwdZ7O/qYwME9i9X74nZAjam9r3UzRiNcq8hp9uExxFiIrH5P
dEPPmYRYsT+6QcWOFIDVhvqpMVvPtkO5CiIcj1wlvTbYFTLJPffpY3a6mn6jDf97
NQsnRAyi1iwg++mhmW8nvkJCIC49srhbw4tPXRUJYmqcmFDP1i3cmOd195DD/ABb
gUPgz3wpU3/8DltMv/Uv5b4OiRAxRHiMFuW4JBsvPmTmUN/ubxWbfpa8pHJ8/qox
jpGLEXKngMPBfze5+wHF94Wlrsiva99yYBSuwkame/3W/FEddXt2h6k+i8pCe6/F
+6Y6kByLAbupY2H/MfO1iXPwCoZNM1akfqY/JOabDSUFUl/zPFG5rXKxunu6qBQf
PUcS3c2tgQYni0SFt3Ag5u/yKdzpv/Fp4vpRiv18eH3e4TOROE6l5zqIsZoOIWj/
Ewl99CvFHxR6TGzmK6odPejbupk/w49kkDlkXIUOSyQM2Vu1WsAIjmHZYMQMwnJn
jQQ2XWbfuj1f83AdnF9foMFlVLawlczpYX8f/2be7TM31oOKZ7IdMsobaKmz6zaU
zpvsNYR/cYB8hHuEB7fpyBsTB/Mje7f0wi6dj9h0ASmhwKBJcrZljPyDASPKXlvy
bFbm5GjH3FTx4aRHFgI5fLNMOpemOdAPLY/fxhnMI4ENK4tFj10X0CA+nDe6PwjL
qltqg+TyFnLbwY22OXGwQ9YBN8gLmwxtvEX3Gz6RdCzJcF7EjJgbQeG20AWdxfH1
QEon617A2EmVpA/JowslaMnju0r81Y69U2dQwh03bG3QmMM1kOP24Rb52TbMH7s+
rOr8MA9ouTUt9UhZbZ9E1A==
`protect END_PROTECTED
