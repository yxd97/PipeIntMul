`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EYCVbhW0vQ3G33FYDstbl6z3oLliL5EkrHxk07eTqt8RpaMgvRjjskdrfLTdq1U0
NVibmK85tvdOCKcgXN1IENPoIuz/sK7kIOrX+T5hhiOuINZTg96qMmWxnzkv4rZm
fUUKjf2xJwlUD8dznuhbOI3YY8gHDA22tzYoKeinf2tVRcr++c+Gzm5Xf2wTewoK
ErEFIV7I6iONmi5tO9vDy3VQ0+PrlrLg/sE98p86sYGPkjfgZnxg+qwhG4bqYxQ8
NSoCV2UeBr5Z71p3t6xaGkIGiMnrtxYZEdRBVL+/yIyMqf6UiF08h6eiHW/R8E5M
27D1b72OfpRPsd5NTU9wwg==
`protect END_PROTECTED
