`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zSgclhDUZepwZZwmaXqErN/tf6EuN8iFNkl7hfYcEn0Ob1TftjmeX5cvrlCdkI/1
Loc+0QzDphAaG1oMzGbeirinnbJ3vxWr5j7uMkOpAGX+Fi5hWdD1fYshMo+uv6Pm
Hz70EiTwAo/55AdMTVM6USDTJ8Fkmj8lXXUP0fCVOh3RhSdt4D10iMQEV8WmMB+u
xpvC+Ju8hxSuKgt03qUufQAIFoT9TPP8dJGRB92Zc0IDXi0nA1M8GQk+KJ6bbNK1
ufeJfH40OD9ibPrjSh/pqU672mws3babdDfgZNX82I+z9EzgSTyWwqXEJhULYRM0
rRW85nNW2ryCvq9wE48aP5qRDotYlparN1FajIyKWW1QpSxuVtQmvKZLWYgrrKvk
N9f62NQyAb1aaPEA34ASt32vlIHWqucgMuQQWzraPZ2UhKOUMTcTOq2F+o3AKPaD
gQ6psZvVNnuorhVbHPlJgbY5eBc/4okhG5uhaz+d0er6wW034lFrLAKE9KEuvbAv
edNK8ujy/TNfZcsDXZf3zDxgEUqGN5WcTvJreHa7wqbW5nk0wL9wC7+qfBr1bxes
0PBbmdDZdMa/438DScIdek2uDYnX1Cq9w+m5tXA/Vdsf7CvM2UeHLNOeiashJDZy
iTZOoSkbrggHUCmXRpKXT+3545PyY9cJUhsll3F2FrJvBoQsfAy/rydjaPwYYeJf
56S9SxNTp59NpHxRISuzCW8yOXI70hcyAaR/kuXZcnGy5F2TwrhsVcDaAS4mDY9l
PohgyfdX4CkzdmllB7zNxfNHIvSCHBdkxsr09DXL5XxWpLd7n0mAGGa/dOlzJcGl
fJ10Tt2cI1fJHrYaqs6QMkRo4SI3mLp/X+UPkqqAj40=
`protect END_PROTECTED
