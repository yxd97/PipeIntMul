`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CFqDtEhR+rk+6/1B/gGDYTzi82PAP1cVYdqcYGNT4R638EzHdLyQjDSpfC3EFj7O
vcPkkhXHYlRrHQcagCp2153uepswVWPjc/OXwpDl2eLm3eG/LrTTydSWPqF3hbJ4
wTOL90wR6N3FA8dxbBX6DhNyTD66ZqScreMjjmJXobzqskXLtlYlxY6f4Mw2U1/9
xn+2cyP2MUjKo4H2WzsdpB4eI8kVFYTGeIb+8s5qBGjX0hOS7YQTJBtl8i1cQ1cg
Qhq6Vmr/ELrAsEuBMPMQfWXFC9Oq2twyzS3cWsfUDp24fjH2CCi6xa0Eq2ETIanN
kI8TXIxdQm5cr4eT0hb7y0dr/p1TeA8Lhqw38Yow16CpfW5jMqRe97KnIrao+3Qn
uDYEPxA/aDBOGdhh+lXLmA4DMHi2knoMNVrAHsHd9GxAS5ZKuB6bwpJkKPi3nQO7
0SdvPooGwmrJp+HI3UJc/9ko+i7UtjjsNhgh4o2rj70GDayOLFMBlhguVULnVbDQ
jjCi2YkVskoFrFvyvdtv65ifuTA7g4uGCEuDb9RY1Aj3TIvNZjJZ8RXM5Lsk2Xnq
By9c9z11C07K92N3HL84Az0nKcQkAdJjIdqinzoWW+k=
`protect END_PROTECTED
