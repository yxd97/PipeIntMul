`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wAPVjUQ7H663yibAralQgosOsnXWeSxQfRIsaK03gPU4sHRFFme23nYhfbZJKp/j
ZrBV6OjBziaVwVEsfm3eLaAbDIiDH0TFXnZ7YBAmxW3bzIJRGXwm07/tdeCapOwN
byxW7V8WPepaFVQh9Ywbck8KJd67P/cc2WP02LHyYcxfGPRsqXtIo4ZZJVn9onaQ
+Masjjlbduzoa8VksXsor0jriJglTHze1iwZslJf9tHfKAypCBmo6dft5+k33ugy
9vvcmmJxKAp5LlHz1Bw2B+H5Oxs9S6taq9kY/Ho7G5nAW5S3B/x5tBWy/lEeiuLq
lLvbGIHA8wXPuftAjudPFYGSM/WKp1zaZebiN3/80vusC/y+F5TdtVvmBvT9YnV3
XOk85VALiZbCxbn96rcF7q/u06dVAQTEiaGQ6vnSizZM5tsfHITUP2e4FEJ9jBgU
QtaHuHxDeDfWYWvFlVGLvKCtdBm+kupYYzCkNIs5Y0wVgMCfOQFZWLMZ+XKL+3vO
7EKtoR9zZpKN645H9sfufBwVwSkGYsQX85RiKTPTuQOmlLbwLr1JDXG9Jp6NVVrq
rQ50E9XsaDRFo1BdCh5CeSWaPCbOEs4OhebvGiYL2Jag0N8NcvyoE/YXBDmIlGvQ
HfSUr51Mdt/8XvogW/brP0a9kiQwz4ZLvGKJ7Wp0A02K7CWcR4M3GPGtS5T2F1b+
TfHQ83Ggt3rWee2VBUjmVmOXerx4AQXCI2ETD95B16pCyZtALEdYvoS01xodKsAz
2z1ag/r7Jf3E07CHunPXK05TsWFwRxX1FzG9usQ0Bdx4UEUldEnLneaiiFwWm0O4
ObjASIvoCt0kst6hg6tAgjRnP/1u6JzUKaNGF4Ly0rg6ruLP5HtyTMCJIuXVQlcX
yz3JFRUrCGJbQdV2ogfVe/tYJqxE+Sy4B2FB5rjhRQcngwtBhrOoLJZrFJb2X3JA
lU5WaaRrGVj4Uzw0pC3AYQYlzA/lTsRdydpb6BRNhopwV6XlpB8Uteut+fsmmCum
6f+2lXWCsktLr9fEgsxBNfyNmEQrckw24FWUwcd8ywOE6FLSVW3A/2rh7yuvoTAE
QPs8w52frRLDWlmmgTOp6P+DEyTtDci+uD74Wxh2XKkaGYWdR+jZEvNQD44Di/Pp
WXCjtNILQQadfA3Dtt2QxON3cxFOr98zxXDiA7u7HO9NCCHsv5EGmAY6uHZNDNJ/
1hKAtlVJgF1pf9y4YzyuIs4W0d9cy7makrpQpoG/2Q8PuRV/3HQDMVpyaH4fmTl0
e+p0jcxZZSr1LJHpIFA9ll0GuVMcZWHRNfNmVPrUJjqPP1qhIYbSOj32BlYZKNGA
icUw4Ith0huzPCo90bwtjHHiCDnwbjvwmv10PVTEqmupJ0qmvLxmEIndIBXbyERQ
cw8C0MMpzvvQqV6NWEk3aZnP3IFK6DL1hf25w2pWDLXp4evXqRcimapjdqWaGWRJ
e8QwE64oNMXIw9ohZjh3cNSiguMT5HTlIPtpkjUQbUx/Xs8gMW2mA8tUiFcxGVtB
fjm3Ogd7HO/wePbNR98iZxcz5cpZPah+GczczsMYHflFHSYiq/qNjLzSMcF5zUmU
uA++uZXeW1+D8byvNqtd/vat7wg9tbgKlL31lk70sqp0xr13Wrc0T3NKUpwx8i8z
StEWnYBx8fWPyMFZQ9HuZJ1r1sCY7XY8hG57wmP4Xso67nVbPsVIoP55bsJ/E/6r
huqgtAmCkdp82y99MkbRaTeYu+MvFSf1qQDqZ4fRmCAQldPSUuT04nz5JODP+j/E
1t60QrahU/z961NjmdTOYbTwlEw3LhVMm0a2Nr9E6p0deGCFchH81PqTK2xoLuuQ
1LIWYQzfiL6V20tZfExemDZ4K/zHNBZnUX85ZYLR87CBK/94dFMhgxf5LcrM+Mff
wGrKDgxJsC1qMxo5LUappz44+cec/WZ3hACyuI9rJGL/AZlenzyclFCLN5o96v8B
`protect END_PROTECTED
