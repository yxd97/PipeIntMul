`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+fn57lb9oLucxywJlYZ4X4zuRzzIT8rPOg1P77LjkZjv54Rxclcd3erIJ8wtk4bT
izrMr0zMwX7KlfJs0+6vWNuWAGAjX8dhbiOxDUzk7VNJ21Ac3YB2ytYUroNPT/RF
eclZMTy8J2kvjfzpxrkNUmk4msr183OUELYStyZm8kdG0jK7I17PZbAwN2bVAfuw
Eh/0S5dxmQTtjHMxTgCBEexTyvnozZ+p8XXpNpeNRebeDj8i4nvUzXJeDlR0YrBa
IF8a7z6liGlIFfWIUlcq5rTgWjPRkKvgwL+yMme5q+1D4bgKwvb9HmwARk5DO8WI
mFtGUX3iPRu8b3QeIpkdR08VPHCi/Wg7jP4xtGaPijw4C9kQ7OLKgQ4HpOIy026w
DzALUi+nFNrWia6P2zAjHaMscg0DSYpW+YQhai/W18Y=
`protect END_PROTECTED
