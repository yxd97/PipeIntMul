`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xCcL73T9X1aqeUEO2njXjLJnRlgNdNXlIe2iE2w9sRYJ2uj1vtxQNGrCaTR7NjQl
apsfwXrKLs0amClEBenEdFgCK/+7Z6E88hjJ8xWCtv7Gn+MAclAMiAxZlncVEtY6
HzB7tcPu/qHnCel41IFo3qZhKl4Ga+zpIDkOt1P8+MkMfeyaL8djqXLW39sploCx
mNVhvuqCnnyEPvKjhjt0MbKg0w6emancV8ciDwBGooD2xOs1Vd/d2qGBQGmVJ/Jc
bGExHjBabd3f8o/3CzlQFOljUmU5jbqcT0haz/U5hZNgUeW4hc52uIygZjmUJ553
hKsbxuJvnx0Fu+l8wyK5DMjQqHgxYXCH3dqy5ykNdwXPjKsTvTzH/YcaauHWGWdr
X2dxIMIxe9yjK4slc+6VvKH4r7ehIGKVy4dE2HGJ9zXIJ6fqv6EMcshNSzh8p3Sg
Uyos+NM/cfoyJS3tp/5JjA==
`protect END_PROTECTED
