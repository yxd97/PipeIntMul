`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xGEM46hzwQlw9tto+zBIsq1lbnUjTkvUfYVihAi+2wP4OjSfoFby2nKLSTmHFKxr
BOeD+WJQllRqPR2vEHiLsnes3TAt2ME56X5jjOl5ofoWsrjczCiKJ6F8ewjiCOAW
b1JqSULaweZ/WsEkzP9NjvFFa3DFSjc9RErdJokXZxHa0/3VpTQHRXnXc5bApgnw
MPvY8N2pugjS5Twzk6lTMpAj2tKSaDqOlQDmrnAmBobljmtu2hmT0g8AvWNxcH6a
OE2SZ7CqmghQ8o65RoBcOovzfcJBQlW4Dvbu6zVEg4hP3QMY8Ur5A81T06hO62Ie
ASmPAWiU1uMRZ1r4qo6oOw==
`protect END_PROTECTED
