`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xp2poF7xojuEF+R1zdT9K4ah+BM0EjbRn+thFmiDrcobCEpcMgL0Cf9RUAGWXjSe
7JgFSQxbdSsGZ7ZMB9OoeDGLunPGiTppW79s0MctQFPBFEgF1/2PQI1pqctDZ34d
EyidDsf8DRJNdFf6zJItCOghF4SKOEF1/gcR0vi0a9MQ0+lu4vPDKoH2bmvLajWs
Rue9/hPtGIZMzNEkuXMWSX3EZ5N3yS8Lawkdo9N33PJFibhQdH0FbGz33DkSjV6F
9oaFm1rM1o4UAxGioV7+1JIj0rDMcdjKWuCd9gVXntCSBaKySEZHxGxch8tbu3w7
kQb8C5qyb/eEMqmB/NdeMZGioexgC45KJbszGldMG5y8EMcAFpgpfcHuEXTUK6K4
ojzhrfP1l2DQACvxYVHKTzQKtyQPSK9D2ibMeFyxPiQuyMo4u873q9BiOE1nVQJI
Se6wwX9Eve6HZlxOqtD5moDXP9r1Y0+RiwsMeZxLTGV8zR342lG55duSChKBo4Ec
qxNm5MKe6p6gNhk6Zzhk3hjcIj/Yw/ibmm2erTRqQ449qoUD/zpLkKLd1agS1nsL
9wdk4/pGyYUM6ypQ57ZOmYkCj6L2Q4D/h+HUlUJYpJHw5y4POfxoMCpwZVCkzy7d
7Vc5/3NbPdZkyg62mkj1UMmJorS7neL+5KQjHS6Yiolz1prBbVY3LcUsNKVju5QK
YP+tyURwaBSKiWj7kHh9BtACdc5mSqqDF50/W31paomHMhftr2ITKdella0fvAKN
m7jjR9SqSo6PumHWX0q6316SHmUfswV4lCkNgCtL8PKb4eY3ZLsfvsgSDhTRU5WN
FQC+aWQK09KEHo8Y00yWiQs4u3+NKmC6Sx2wVHTwZEEzrf21gWlNgHbYVQlWfDgw
l2iaHPVKC1Vy4CtvkLISqDCuKDvhytzC8cuC4dwbyG44i57nZ/L5TzZOs77kH3vI
xNJ0igAM7MZQKoqjucj2Pg9F+o0t8RDC4ElaUAXQ50XaycF6XBkGvIrtyfNlycfM
7CIBcC9gIab+2xwmsVEPR6G0TiMs7aLhMCR6fXyHnx1psNkbBHAFUFlyTRpThZFZ
l1eagRCqqaRmaUKL+/f1LG0AphKCd+ysqh74rjS6/b87ERg67apUXyfvDncDrbIn
y58kSvuZ39L/lFHsOLcpxgjVcL8E2WeDvw78ywH33oPFGwWYGOOPnvmoDLm6jerm
ZhzeEr9HK8OPx3+9cLQL5SBdkaWSx4qzoqoic540QnwQBFnMOi8/IJ3mVPwNUwnr
qM5zVAEdNHCvC9Aqfv8dKbJiAkbqnM3GbU3mMLVF6zisSGYKL/8yOQUDIuOqaeKn
8RCn2ueGDGb/zYE+tvXW0qxXCOvKhRw+cWsZil2i3JCpx1OtgWl/9awwtzjjCQi9
S0LyA/5MZn7ddtwy3cYnqlUC+RfpNW17nf2kieBptMD8N+hA+ecKFwM5hW0MsBoK
Y/0iPI/215/ugXQWwq3+TWCXheqpceTR1WwcwMkBvNChmzPpA2p5fm8dCEPoFfTI
`protect END_PROTECTED
