`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S8d/DG3njfVHmCLutwiDwxa3wTFt6SGR4YOJuLTGqxa5DVvblG3Yfm6n7hvny3V9
wLnn6HMfE673D90A22KfDwP9S/DVe6CW1VucSl7GEhw3aUBKUT7Pd5PCEOFFJRvy
DXXrT2ReuV46Wa8vK3kpFs2EuFIgDg9m/rYUBugAyZvgTBD2m0mCqDCFLOKDI/wX
SNSetvdlc4AhUV9iWQJ2Ukw4Sez5fSiLf2xk/JkqNhcLedaGPT7U12DMH6A4MfT4
Pp2y+IF6hNDkBkSaunlFAoHlg5IMKP7QAOn+NV9kVQ5R9f0sTGb8+H0gf9HKqKcD
`protect END_PROTECTED
