`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pMqFRNW93KIEnqvvR6ldImLaiFQnEFvCaPvYVOx+yB0EhT+g2H2qQiD6yz4uAiaw
0p9ElfMfjsvEdjcrE+74eWn4+yFkVUp5+wd0gv8yaMsASH4UfErKq41GDMd/Yi9I
KKTmJ1WDBJ6mHm+TYl1ytM6bfFu5BJzrOqVUhssbbWhkEIpXQYIaNp10T39CwYeC
TDiqZ/DVOQjsIjyiPM5muEW8/rBuW2uKdtLsZhKRmdl71eShk83tGg4OfOEgIhlY
n7zA8vmwF+LRlDUACJh129y+Aw1DfuGXl1Ke3m5VbEriZs0NvVIwFmYznYf0hvwC
0M70SiPmvYprSJPQstaO7Io1StiSofilYDMrxPn+otuABgumn9j4CO8KC8+/436f
ijiUn0B3AvV7oXNoJ1IUOU+AsE3zuSw3lm25aGbY1bVubP81gMIeLW0c2DqYRruv
vLGySMsiD3nK1SV/kmUrhNc6WrFhisEihZVRdNlWU6gnnf1mVPqVxtrVHBauCYmj
UhLfLDCa5ZWXv/2kGBT0A6P9all6QlIAeO4nRlKctD36O+GUm31gagXZNrkEiYQO
iglpGzjrJOGF/dxI9nopEgv3tmqjjPig9bgI7OfNlRlN215vVsY/AJh4F3CQMSdA
CqU30/xXSpKu7RoBDv5e9H8f/jGod72/iKdgrt3ciblLSWD0T0wKmY0YabITNP7w
l4JCT50EZZzXlHAKqYDM+Iv7ygNF7pLale6GWNyDIXUh4ySXWaBf/Fp5xrj3lzPc
LOeHVfov88bf3wXwamRA5JnkQxGqs4TPQyDKNCC+/LelxuYkGQu/kwid+jqw3bKd
5TF7k7obi9W2fTUe/OPIN9A7UZRpZFNZ98Vp5b1LVcqtWIVeZ/nnir/nj96Lzdqj
MenTpUtWTYIv/MmyW4adJNvbCloMQ31b80Gi0rWbJQSH5DwQCehOWnPvpD5yT3MK
5/5ngKWs/V+sHf688QGpcx1yeh9Y4V0N93CP9xSJstUiASp3iSi35sSEOi6XKM4Q
kFKG1A7PSE5wmLaTJgv10hRlZsTI7Hg5bPzpE2ovRaH+yrRb4UB4qBoQZx9nF900
OikPLtj8uGUIMulOqZI8TA==
`protect END_PROTECTED
