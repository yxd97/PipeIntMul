`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHhN3AFpAIOMn93VbctFLhe6Jp4VK5R7kF60qSktvcsqbEz4c4mF9AtCC5ZDkhdO
6zhlFb0h1nLl/Kl83juPl+RSNU9DlRRwh+6eNoecnzgguPmM8KBYHDbFPYCzYq1d
ONHXBBCGWMlBDYXsumqO0opYzUX0jNKOCSSfW3/ZWc462DkAiw54/j40KouOYAF+
hKdHRVnhvdTSNn7AAOQKOfXIgAZEie0ahFu0gw1E8O5dRlFDUIzQKGlxBs41wtS3
+5L5/oD00ZXqoSivCuo1D9iY88xHRw17sU1Utg2eKBi9SfghSskv5qCII0Y3BKPH
GM0F6foz5mM9G/AcbTGkRxjsuyfmhQT8kAxg8eyTaMMdF6gBa/UN+HVlhh5tFPEn
`protect END_PROTECTED
