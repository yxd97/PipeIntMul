`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sp7fA7KYF6fO7vXfTtpAowdIjkyVEhhi+7WKnk+k1qDuugIiaDRn5D5rUZ41xwFC
YDZIzOJBicq1NYvB5c46nQo7Zb+u/3GB5X947EZP9T1xa/p7ekwNtuMi02LkLEk5
bO7aNvHqJ9TePVDrNlNvhZXeVK2X5/6Ir3orLE39KbU6HJxi9auRdssgBjVoxB33
2KsJJcQnV+iAWI/2VXz9Q2DsyAp2bKx2IXU2AgjoB5oV8iIoeG2LAw+8ucUUT5G5
QlrtyCjbtMOuVd3e3e7T+E1saKNQmp0mEzAzAHdm0zEeC95TUWJ6a0qshL7XNJkg
8jzVpZVTOP+qMNPziDKaRthVfY3Cr/2OP+m2vvQhw+JHySB89nUDOsQSBFQqGKYe
EmTvU41yvWWRMoiQkY+vw43XibTT42135i56FqydA1uZavDllSR/8CbLkDin6V+t
cFcMcgmKQYnY6RTSSl97ibwmQZN61TioH224+dwFVEZXosWrRgjaitoL4R6Ly8UL
9+c9elw3EyTOEraNmMtnsTouakQpS0UImILJKDvYF3o58WBJOzE4x63RwJplBlh0
Z5yyPw6+HHZbqo4wrvxKwtrll86M7KH12W814PTsf1gu1tT1lgQYS1p+MRGertps
iWN7xhsoeatU77Dpv4LDi7iNnldkxZ0QYGiSXUPmvDeEm/0QqKNekEkL+X2XYs3S
SCk9II51BbNPx8zJOygZB1/+qLuF/zHYFjlqkjHFADoZxjuaATf/JcIERlTbbHVE
`protect END_PROTECTED
