`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+wMwQZjm4Tta4tkxD+jmuQCc6O1sJOK6yioF2SRVXHDQdOxenZFdZ8CQSOUlQgSA
5f1Y6bLAw6pL8hGqmnc55G4CK5KlBdXZc6mgxLiPWpGQj3hEjzb7YlfoPjtvt5bi
966qkzM7GlVcp+grJiu7oVzUwKfpI78j5fAY6xCCjFtIFgetMpD3ALi8cTsW4gfh
Ek9aNq+tho4lj7UTaNzgzznLjnjpPZFSdrTiOnSQ0mq43xKU5u2uj4hpIOTXYujt
ZPx6gCRY190dNT/Faq20BUcaqcyiBpgiq1vH53dbipnIhqkQyHDqEP1sFnRmOw7i
5fs6jsHO7kkUoNasZ++ZqYMUtOGNq2gPE1zJIhF6mqwjr6iC0PA1eh9KpcZiPyLQ
XU6NoKwSz2c9TK0SoD6+4QH82TA5iLTAFSLFaFa1uPbvGVZg5D7SSkiW0NrUl2QC
diNICEzVeundacyoEkSfjpZVm8l8X6xTXUeOZXQfOeTzoOuxwGTb5EKS7H4BlURP
yrepAujk9AoDRxbvP2ncxLBS1RwxEd71fX87MEWTWHi84298cHujG5qRn2rMNWbc
MYelQBy4E/TarSB9CV1+Ja4Sm/8vvhXuvW7skUNI9p8V79rjBLPdwfkMTEHGBZx5
rgRBcjSlid3GmrByISPF+VqhLSygDC9zjIdSZjOBDedAijMuQRLe8n7bR8k84LC2
17DEYbUxnFyo/5XX149xVyPLynKjkPRraoMSi+efJ8jfNG+6EOtp9dmJDKt1LXDQ
NKJVNRIeYvTwTI1HlDtF74j8/qo9DcoBIz0N9dva+rSYoQg2DiKVWWOdMskXYw/T
XG57/ItwqHUtq8bCZL7mMNi14nSbcVMe5QIbYgIxzXAoXYujQ4OtllvOlTZ+Z2s3
d9sf4/63mYayQIQ6RzQEqqXM6j4zQDIFSGRRdbL2JsPmyE/iQWyFnWrGfyI7FSkG
yoOk1Q91LakZVMLF/OfNydn+in1Sq2iJr/0nx4ebCN4bYNwqmN28A4CShQl2QXA9
NJRLKnbIBYV+BYNXpqz5SQ==
`protect END_PROTECTED
