`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BWQes+Djslhh9biZFA4XAg4Z/Gg/G4ToksGpH9vIcf3zfEJUTlfjVPOsaakOdoj
SP3g8zVCoy0BLKyihPNjFJrLIu5NEGZKZrQVzi2PilzG17S6/LKAu7DhLYVKOjxB
WegnZ4UaqtVsesfRYuGo/pMdQUTMa+iFLSJsaUS/gOXYWmEgzJzUP5khk9boIA/W
GLhhFHYWbR+GgPnT29HeibZ2VmVNv+CdKrOix+y/Up41fRdIS9Lj+aKiCmL+w/vP
1v+AmhXHmvPSk56rAbBYqiRt5f14OmwQVfR0uiI2/KGDox9ZH8AW0w/PJ7usw07P
02CGJsmLQZefxzMdybww0BW+yjOsALhIL0sryrIYgFoWTOEFjlMGZ4S6kMEbNuMm
I2/n7AvhGas4tc8/0fEverNAM6G3NT84XLsg/2teAm/2S5R2K5qD8kgxqYP+xBNS
gPygx55w4jTDKwTiKA3V2XyRWwIueeQRmxvF1WbCAT9rIdNu6q7zBUWXH0KnGrz2
/vat1ts9IJH79iRiMS6UsuXLEruKt1ai22LT9GLuh/nvfAq7S+r0oJLo5PRQnrnS
D3JO6srFy/hWwarABYoSdHABUEA6ydgMlQcdsK/Rota4dgz4NOmMpe4LrP1mMFJW
MzHz05GqzezfHcmj+F8L8rWMsdGDhrtQJZTt7v3m6BY=
`protect END_PROTECTED
