`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gMHdjVCV129pgw6mwlncenDhjz/W5FHQV/NXT0vq4Nwq8LEVO2sARJ2mSu/PtUUK
q3wrF5+HytSq+tdJDBX10cBTKT2s6LpQABxUqz8HB2clHjtYRmwgYLr2FDLt++Q+
Byh7luPbpmZdHZlQgdRgd5MMQ25f/cutK1LXwGB7E7afzoHz29HaPv9Ow2e9Pqdt
QcJlhlf/BS7QgOXtZmM+uL0K+kuLTm6OWLAVXpEPY9oRrwV4dAJZRukDpPqhxzVO
1SVpE1SGczIH4ui+2XbFZ/8OcY17wDj9aWlbFGVoa2xwSuqgs5M2VWISPDC409x3
nGscJvKqvaiopRRxh3gQbKCLPV5XP5z6PSxluzEqq4KJyeI3jd+/pdnNi/QOGoFw
mv9uhTelSo42HItgWEC/nDkVTGbJNxXrU+JDJEyU1bv+sBjFKYaPblxMPCY1HXjP
0GAU5SRk4+EKe+zF04EMIIFt3ZFvSwkmKRH9SIQc9jL9u87grqZutIEg2KbFY9KR
Nvk+HRlLvvE7DHiRrqiCAJH06AkHdTl+1mraM1tgOJPtmSGl6yw/OMReGuH3sd7j
`protect END_PROTECTED
