`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqBY5rdpmm0l5q0ZXDsqBHh7zGqOtt9JYBDLEe+08TAsVldKUDgTYvpMLG90uw3L
olPfc6gxeuR8bJcEdTFvrpRYCqcqwigTXI2NpCtzVxm8sh1vFh44dBnZQj6jEwVz
ZTLd7pGmtEkHVPMsm8WkGchRw1nDdroxoioxP47n1urXS4+gudRzOgLFiCpCXXJO
Dc4tXXuc2ot/qYeyJiD4dz8Q4WiWtsnSEA4jXf/O3U7+jLbcsP8/dAIfBs38U78F
tFNvTrIJeqIY/5KLEsaGpITNdrkFsLJ6D147qtNsfbr4Z22jbZK7BwRczoziyFts
G/VEw/OITsP8f+dD4HGnr4+V2GYzMlO37HoVvsxIN1b9NA/aZ2c2uzzsgcwG8AfT
0hZb4BDibmGWqTbnkc5uRQfrhBS3bwL7rRRL/HAOrjo=
`protect END_PROTECTED
