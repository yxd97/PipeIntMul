`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KuA5eNI0x/C0r+AdlwlCUVeTK/SaIyWlygrgtm6Kd8kvGRuHRYmD0q0xuD7O8siN
ePi/Df2V6SLFJr6kB2Ed5gOIc2/yVmzvtc/sYWQnRbmQ6hCNZmr4RXXAq1RKdgcP
8umRjh9eiJWdaZ3+00vG2b85HGEQ1dsDt6R9Ny/nXZCp0+5NEed7Fymck6Wm4LFL
BebTTJOCCYUOsP69PfAxkYvG1208b0DN9TAfEUUUK6KzoIRdghH7FWRinTDLArtX
1nNhh330Dxe9DmD1majtqv8rjgbY8VkTCEzVuU6KAJQfdkT5Bl4MMB+Fezqv/kmp
vOpmphUmLJkIV4d32G4huMBFz+y1mutvVY3WG60gakuSIXv64mxamdjC12bJaxeD
68qPd01XVSHd5IA4coN0wCY2a49Yd/2bJ5W/0jxiVHR56K0XMf3V0pDola4rlucw
KR1Mt8VjhtNYhGPYRHu0PeiHqDmK45GGDJT39DtHHphqLwYWhSZfouX6j/jCwmp5
P3NFynSV/xzXJqAs0SZdjHrx+2ICalbJKxrxml/Dj0Gdo+7COWJqT2I/hdBjzq1D
+nB6eL4+ZBex+ndRLh4OgeGKvUOeGglJB0OUBAMx2Dzlv5L0NogkmuGQXOBBl/8C
Xm0DnuW/jkHe4L3SP0SiQ1UkkkOM1mvXf5NiS64XO4CXCZUeNpnQc0ssU9DHIQyI
PnEnvq/qVor+sBfAfUycOrN6T6tl34VkMm9gdP5fTYUaQ4CLSjqXCvWI1fSBxtrM
QMFUXbOakWR/LLQM7pw9XDjLrhzOnniP84nzyNBF8/Ln30EGLyQw+YpUXb7jRePd
/2+wu3WtXoh3D3HXPlamK6RjIXqxb8soUX7B8igmKHLTWrMZyHhYLpInUtp+79UK
8PTPQUY3iIl9/VmAeN7S9Z8slQ4Wuqjn/lMWxgP+1/0ZObiUSLL+2Y7/X4ZddGT4
0XwxP4lzLw4e9ZaD2EpJ+GLYYU4dfRIZuxUMDDiHHdUMeIgHUWnBosYUAj0jP+8f
MBbMfyA7K7EOTn4eam8AW4IUiApZ1XNfc9fC6Ix4izkx5guDNyJZr2fpS4911M2B
Tn78gY8sRtjgf9R7mcq/XPUwx8fjxgbz6wmbtJEQ9EJE75DQWr+eij1biASkzbA1
asuJsTsUj9dcUrLaIexVDJfW493IlJOwgAWfJgxkEqIUrOynppXD5bRX47YCvHNw
qNq4FxJlBjSUfuZ8f6by0QcYG4YUPOONeCDeWIq4xHCxgVok6Q1S1CHprjKhQhpn
QFf1u2wr41M4lNPGgx7p2O8RtYcwMbuuIiFZSJPhAMVojU3GRtuxvcY9vf9yd4SN
wBBMzzZBe1qTMYQBX1z1Wb6wjsXFu8foiwMFgQZJ9M2D2R+OeXmgL1g/lw56f25o
sLQSbNanemkIooU4BuUhmCIASBsP6e6xxxcesAWUAU7WDsJ2kVWYbJteTCpqjDyJ
hVIKNZVJnx+e44sH6+ctjf3xuaS0VSDB1kb0ZN0n98oq6+z0bNbuMY1xwORKF9OS
4WFtsHfQHXrmAl7gJZXHoekQDdBbMv+aOmcVB8AyuQu+N+dtl1/Il5coN47SNbPs
ubRr61bHVMXgo606h3HryiwYIozUETT3LCkVBz5nouYzb01ZY6xLFApSNoNQPDS8
Hb0G0qpKLLn9sqDjuym57LyZi4DkV51Yo22ajqW93tOGV1175xTbHB/lTnbGicsl
zSlRyqRVkwWHyPS1UilLejqwXCuRz1EmBYq1MioG8sUQKyj6+LaavV4suL4XAREt
hd+t7VmlO3lA8Rza0miWQnoMMi9MsrxMNwCTj5kpSljgM1V3PKWvD7y/54FvrOh1
G0/Y/mvJx49wyxQCD7SDSujSeCHvNuSK5y/injVf96SI3TaWwwhNb/8i+Tl7xOlO
uaFO7t2DtCuzbh3XFwZOnxKmd2fG2MoWbFf/YDt4EZgo/25tQvM7sLHReUO0m39Q
f721blfexHvW8bHSVI+2uKBMxGYb4P97SuBhdnO4InRiv3Hrj20PdDQ3tVGxohzN
v68mQOv80gBjUa4ehpjdkAs7eJ1IvXbVHEmZM96eYz6vFNBGJRvCQTesSnJ/5V5c
zUfEhid/PkGmfeobBTB73c4CNIZZU/EIW/Rqmi1AfSjDF+TP7jHFVJIMqYhNoNaM
W5J9hWF6hlbrwC7SKaPeD9ZTZSSRwthfUcpxitmdzhpqyics97OPUTngRE2J04rs
R/2V0amd7W6o40fJOT8e2zSFecGx5PpsI8wS1Ycz+Ui+ZsA/x26q0LZEj3k4Z16M
QKp2+wy5FbGshmuwINRo0TbeYlP5/knZSAd0j+d1RSultTDTiyQy6ToSUyD7q3jO
9QlQna5OXOFC/uOeeJZvkTd/GrRDBt22nWLgQdDaqjVD2SWcAT8+RS0KHA5oC5Dm
rBkNlGj0KMD1w08kEgeQubwa7uRcPJwaubfnZcqYnuVwiRvvDOXvLFWXuGqelCOl
/wumoqIYPOPrO6vW5nLDIKxePVDExILpUsVk17QEYO/AKJ3GcNesnDYHANkDn7Ze
72S3jFYaBvrrV3N6T8B34dek/1DD07zyNpxGs+p36LslITvGQOi+hbfrv26Sd1lP
S0bFgXHQyX/zRUK78UIxcgT4ZJLhYabYQk5JFWWBJYdloqw51KR3UyV2H+ElhRjN
jPgXckY57VdK0ws+9rbDJClRlNzm7b9abd2rrTH7qK2IKYEWe//BzaUXMNcMBPtj
z25bIvsOd0DcNuaB8cjLnnhvxUlMpvRu4IfSvXkYN8nioXs19gLmoLHiFNZgCxdR
R0Hq08fAvsvzv59+/qUI2e5qn8E2Qqxb57PuhJ0Je60nGE5Fb0fYkLSk9nr6xgSa
GEbVwakF9HUwbsOUVAAgzBi56YczeqS8T9fzm/vKSc+qH1pjNpkvnfP0VovgD8MA
qtEHIgQbogfwyf4Au+3rYmWblX2bKqu6dq3J59loMzTHOizfRxvrTZsvNANyAgdc
8SczktAmuiRfR7uK5teIn+ip2x1hps/nvDaybsTy+l8PKVfDYCGGOOGI7A3yXIN+
UTOqWEH48/8Q/Yp+YAN+qKcxokL6On59R6JXXikOAbQn8UN6eo3rVYOResrwOOTm
czb3uK+DpVf9zRp+q8vV489TAcJithgSWDq613t0OPBZBl0xnJdgdiG5Op/XBn3k
NZsfYGiK9THPtfnmyG5vW4H7TqqgMUusVRoqa8pnxpDYTT+gIPJUxcWYFf2pIXGR
R1VZLN4Ox1aWoCHLlnb0TUGnYsslE8LosdMIZeDBCQNtR+FJSTn1c1P07HwOptTq
wkp8UAsR6qldh4Vsgeryrt7RM3HAbIGehTeWw1giJpNlid0hgYhGfWSwmfqnU84h
KifZBq+Za7lCAQfypX0EHVtmtKs136Lorhl7LPVUn+dkVUCyBmAtFnF+HdHZcUqq
q6NwqhLW/OH8K+0F/HYmi+LSZu+WwDnPoh1jLyPszN3siLi7X0IiK9s5EL09GVCu
jebXuwLqwvZBIIQtLJvS3YJX5QexNjW1Em/X548x7iFZGL6gT/6TVqd661Wm6ykq
FpgwqGxSzm9tqolWlgVctlmM2moEO82th1BMtzX8/PZnQxcicIAY1zJ2PsQkeoq5
Y6XkSXAMXUNGN8RZseFNvU/7YyX5gaHaROeE+024qFsdGTbywpE++z5q8p3mmz7x
1elwi4kV75TsDEBYcnaNKr7mSBW6yIcLJbYzbyEhghYBaG/WcN+OfP6aXAboqnCV
1kLQAm3gAfr5XL3kbOy6u4/58EbL+XrKfyHDfET+4uMBmxBPMGBLa5luGwqnKeAG
Tsi6bviipY+qYNFZUbFPNNGDPIozz6KLYFTaZMh4ghZxOtYxJqUVi21x3TC/OIW4
smHz/yejj7pTBNSW1XSKE++JiLp1Oljut7vOoDV32hDWh7DG5sfxt1E0cCXZd6iu
iZwA5hzQF36ncufa3TJv+0yDcOlpgi3cU58pk170EemfVYhbx6C94HjkjWBKhFY1
+L4uBDRnTXU6FKDa7SAF8RTRy3KFabUuyZYXfH0uJ95cxhuIwCBrN6kRxA7GRMj7
RWQlIcqXftyOFNx6V3Y3FXhfgWS0KUGSLYb9APMQSmd/pMmxermylsB0LbHApYKa
Wx+QtJ6D4S35jNg6ONFWzJluX0uWTUsNwvr36XbiPEmOxUNZiRyW/JhGPtZeU2KD
f1BS+axM1u8/q5X1DU90J845sL9bOM/YjHms3clMJGAw4UR2O4JEIZ2//pCSlp0F
2H+VfWYVLDAHGjCsSq6jWdtTauWsuSs80b99hcabJi5bdwTZrYuqenXQnQ9GZuVD
xurHKSplUAXZerKIZbPR8ig3CguUPKMCQLIX7vQBVSwd/NVaRHYU7IjleKxdy4VS
ht9EZEWuDB3sfF7NzMsmCGlO/765Rf2aZ93yUS4niK6yzeR8PFtfA7s46Kz0Zx+I
9kwjpnKIYQi1FDffxIVzQKe4XkXF42VUJQH+ATgiHZYvKCtqg8HLcWnvRdM/HntK
UCEvSHpsZY8GkMWa0FY3y8WBtOsrR4hUhGZmjkQd6M/AvRojWDhoKi5Y2btvsIjp
WuzbGAeqIhR+aWMw/Nhc/o0pBvxgAbYCXtrJlYEjpR/sVqyhinw8Jh3Ufl9LSVwl
K46lTRY4idTzK5NciKwSmL+LnP6ivGd5cmi3KT6U+ZY73PeOpJ5KAvPbLwNZVUkV
aQE5aRPfeqt9iFyMcLt9rTLOd1c/fWDnXmsh+CL4RxBN3gegSg0BsSH5ypzLfnDB
EZLaWHUjOOaXkww0Nf9z+/SxiHaFn7oT9RY06pw4asKU7yc9//9+qH+APpf15iSF
/XsmrRUK3QSmGq03/UTjUR/hj02EqrF1T27aYQ7vrohQ4/SG6N4nSQt8IugO8uAU
1NGfL2c8oYPd0qGPNcbn/wYBkn5CzOEzaR502dK0kbipQo/cL9S65+fD5HW2RbzU
8mIfKnvcuICiGCjyUlDQqZdXs4xneyiCGqSX7KDrmTKsekhDcjIcmuNYYDs+vfQY
eR4rTH7YbBaiVmUdONj61Pil09vbWI/nTNW/qOqGrnmg/YYH+Wpds4BO3UanbSRL
bvAYe08EZwh2aTZJqVCOXSdO1bwpFyNZ2Gi3MIoaMpO5yEKO2mAjfIrsvjSraSsE
cl13NTPyFMrIj+NwMPyANID6AHB8u9ZKhX/v0iKJKHwv81zE45hmvHkwF/PWJ38Y
WJo/aXbp/wnYtZfytYZkrP3UmyaVDQEGURU6YLWjzwosCSGumJy6n2u16haHi6US
blv+fZYEeIGEnC9g6qbu8EQTvo0aNnvHqEMGz9uN/kXFqkkZ5nZGMa+Z9sF1/YTk
EUzGjRrHXQ4+u4EwzOrqCxx+/xRqWJ6P5CqvRj/tttoNpWiO9+9NvPREZZ3O7gdU
8A9nZOstYtN8aQ19J7xSaAMC2k8faUulviooKWMZjNYh8eoN/sRyTmt4qoHlljnZ
gOgeKDzYvPItRJP7gWRMQV/h7whDPlsCp9kcJ4Ggjk+pgEJ8lTafa8gBvGO9KlBg
zmbtJoOQhl6KOYy19aOilBryViP3F39n3FW6Ur1/VVgtrb9XxfjnjZwEhSYzjg3a
Co9sNo9eaNlf5MXFz3R79kLNvC/fTj8uEIvYzwqJ64PFfqWheiyeJtCp23CR6nv3
DctQ2QHnku+dfj4I18fGxyB3/KciGcsF+58/BqajS6xeywdjJYT8TBFmH/9wFnWe
RZUZd8afQtjSlUWvvVFqDLfDDOEAcg6f5J9OGgwg+d/HkJ6CsRe9Y2zUNm5B1rBi
qPCT4g4mopv7SqbIYG0/ZbOXueJb2PVD09wfYwjCGzy+8A0RSTwMSFDlhqvd1B+M
GK15n0sOBXPqb6k+4HsS3l1NOqLEnJgdWezTD7SbaHbcP4z3WhsChZexKkHIt1mO
+wZQ9FyR8psuuGDor2fbu8U4L/Qke4FzbdCkgfI1RaLyvZoFZYcJ4gRyLubwq8KQ
DE+dwBaebiDNdUnQaSX4fiJJ4wKw8h7Jf+X8PBIkFVnznWGru3TINl1K+KfbnmMK
dwK1TT1f1rt+2tB68uMD/C/0NvwEofFV0IEnAZ2YCi9nidem15c617H8C6c+3t5V
8Wy7bj2AHhrLivqnAYyBQsh6Gs2okpBfes1OQUB6hdIXQLyyhWi88SUsumQcr03j
5+F8k0Vnon+BuNK0w3hOTVVsxd5PrkmmRV9J9bMS2L0kB9IeBfeUeASmyVPIlLTV
Fy06BK4AKnE2rTS+0RdhjsZ2iIR+yaZqrsG8jmx2mu5jLObkP/OVfSVquTzJ+MEG
sSkCmgsIjGPZHl4tclLI8h8vOqcpsa2Q/sPryoXB+SynM84mTukGPJxLOb5Nkw6B
GpnYhnMdVN3eG9eXx2Xy1o9iH72rYiH+usEoQwJJvZi5wdX++OOq7g31v3t7bryB
9f0cDign5vI/FP9LRcqB68wSFBA2ovNWOVWbHL/wUvJlDSb+YBv3tWrnYDjvsrmw
noGfh1IfbYiPkPOvQFzRNjzXDYtRuQKrayJlkg3jEmc75nsq9h820ceNRboUqXrv
Wfg6T/Vq6eSkOetQeiQuN0GWeqL2GHGWud3PH4Gb+hJD308ZKTxPuIMCtICUC9v5
zMIbV4gS9WfxXNR2gD3bBkiKpnyoZTZ8zDIoPsa8JMqMMTyx0kDste6mXq5EK92I
Yj7iU7XXWeyhrVD6HSXCsDIWA+MIpbPTxVKAiUkOT1NR8KluUTPiyw+LnsitDWUM
KqAQG4ZeFA0xq+FAUlwsHmUiI55kFUboSxRomlPCvPZhCYoQK2Ale/QzVwtnhV7f
gH+HlFFjpnTb3/46w7qa5sQOEMxo0hynA/fWdWPz6LKL9kjF1OJklcDY6mI/vzw0
XoePD10xrfPihp1I7Wm6sW8dwTW0fRzyWhCta66/rS2Gc8rGQI6Lw/JiJPIwQdx/
kt9zMOQ1B5vpb48Sq9n2gW5/f2Mwhfq2DkRHMv6RiRKmvNtMIe/DzipYsscD/2KH
2k7QRb1qTL6XFq30eDTw5iSSW5CbrVZgxmvtcl+IeJtrR/F6jtkwmxUJt8zEIWJS
Ocb6UpNqtrs+ZYvrWSCNk2fzVz9DZ2nTIpKV65KwAxpP9InMYBdhyLKZPfdeelmt
7mTcUJT0AYhcGMUrg1QsOGN6JToTB6RU3jSj8Ea3nWxUm3R7GgISI+3G68LvB4kH
vuO01m5LnFgwift/7bHkP4vP+yB4TtUN2BRoUVRGWL7z2k+9PhIucwRt9TyN4Wo7
Aimc406Nyxnn3CtvSDAWJNDXeirGDkiZgJ8VKu0Jwctcdgv7m6ISfH+/sVx5P/V3
LAQKaBdwC/6FoMXcQ7I4ctOWwrQsBtMgI9V0tfhLfM+tcfIv4fJiZ4jnXoEumrD2
Sx16Nii2BMMsr13r8X8NTATdQSlGRr3uAGYbRi0O3+veglNds2t1Fp0Tho6MpIFw
MJGB6ARSp08nhirszHsPjDKnXVYny4Ot5tG0HvuVv/5MmJOGA3sopzg09ESjcSqT
g9vOSbdCVH/j+wDb32TUAJCyaBGKPgq5FF3NKeuCm9oZMcoy7cQUfoi9Cg7Xnaom
vuqiZ/SBMeJsVPf6hmLOf+pt9LrDhG3cAqgd5G2jc7hUl2x5Q9/FT0tG5Yd4wGz/
9gNgdm2dNXGiaPl5iIC3+HBY1QsaQpISv1O/lgMvmThRNgWbQMWUu7Fqjdns+ctn
BQd+w3pWBSJ9ityjCEzT0f46bxqfGSo8HS6QReuv2SaS/L5CyKjNtF9om5dQELqJ
XmDAh1ryMqFXysOsMVski6qyMMCpnAKfF8Ki0tdoH03D7Jt70sPPKEdT3YMdftcq
A7aUoQ8u3dDxqJSQjlbfXv84W4YkaBkp4wIVF6WSe8C85uQNExhr0FZUBUaulzxb
aZCRXc50C3OOboc3kFsbPBTPLdXm4k3ru4xQvaOudRFa1qkx02ES0NxxvU44Zvka
SaX/Qe8Kk5ZXs2y+EASgxajqU2Ca0H4R9Yh0YkpBpoYNMEpZBn1RprH1ZsHJvjup
R5WvVL3rwxrbaiYsWijmjgyl1jlk/rEAnxhnN7v+VF1NhvK8vJmSJjKazarieGpc
T2zRJl0KAkTQ49W461HnWg0tqvmzllPp/wVtR4fIuwQzHVQI/AkLAlpRzXEjTD1F
EeGaPaicIl/sfaFW0pjAJ+OkvxpNW87e1YXGtF6zwALnMC0avaCYtGAmhKcHHXSp
84Y+LxxVdlp5hO4k85bqVVqdlKopwlvwaxKwOAPWOW16HdusvpgY3Txo+BK5AnYm
78CaeWdiCTp9hj1oh2/50bd2pZYUc1BE08QICCgFVR3lXaAa6mghjIhzjUuXjGf/
rBGgRMghzBYJG1ybUKdNPOyosHwGKL2wCAQRr5t6nMONxd3a5rj1jceorv3WdKs7
VM8k/D8Il7LWp5NsLsOR37JgyPpI39/obheWX9towCopvop9HgdIO2ke0oPGEJBs
BgJiTw7R9ed+Um8IIqShOH71dJnpVOEQtdlqAYGgZHQc6LwxhCQ1C0dl/koi5/dz
QNP6C+8G6B5+ZEurTDoitjcaD8HoCCiXW3qB+TN7OsWrm1LsfrCTzPmxrwhkkBjI
fSuAFMqnYo66z3WitIGLQDW+53mZjFqteoSfw5A/6e2OlHb+EtI2lMlOZuEF6jbp
2VVzZ/QDAbbYpX9wRjGjQIdqrEkKVVVBpLVyzzt0WePLHfyars5g4jTMf7BiJm17
uiwiWOdAc1XjP5S4AePE4/uyRwbxn1M6IC7+0UdANwMwNbv5CxiRtH12yv675OS7
Ge4vtKJDBrvJX1SElyF/rispSmqgBzVxT/WLjGdNrH4ZCKyBvXMF9AnXRaOunruq
OQ0IqAfoozs+McYA5gekKqj08xnGlqslstSX4oq2hf+WwLCtl2pZzWxPnEc1Fuka
OYIMMhq1dFE1HOHMEYnH20unWcfrn87Zwq//n6lZBo0N2z3tTLUEKT1NRrK81HCF
ksbxP1bk4VaMeR6xjStkufbnWSE/vx+uBDssZCknLfmKDXXa9nSUgdTvkcbZOcQN
FVmCmRO80CKKkkvkZnCBvpHR8ihexMV5T28wfybA2Ip45Bg3jq2Dm3CB37f1S0tE
RVh1lgXpK7AQUrClw9SOs935RQE3Ciwrc6nHizNG8ACHf2V65TC88R4du1L03T3O
zn8TMBDxFq2oGLttkxEdTSi/79s5cpymLQ8Qc7SV8w6CmiKcJQZbTZAD04Ap4F2m
HU5ep2NnLfc/dxVRam26ygydSBtE/wUJy1BQ71a8jaeeboozbYOHT84/jr7uaoEb
nePfA2MCSiHhymbNlfyBRiilW3/GY7vU/Uu7RvcBzakJXVO+yfdGaJtlEkxi5OKJ
M9kDKXa88i+b3KfvEEHcO7gXjAOJfRc7HdM3WXfTcH+pq0WYoDSGW9phioaddbBv
Puisr1Zf18XlDxVLYbprvYTl4lzV09BZf0yaSKrXOM+b+IIKxlfGgJtWJx3vO0Ar
3wsSMEOedCh/q8W4uy5yYKjR3xbyQuAkjlkfySQfzBl1+Y0W20+tbeHAfjDQaoFL
+fjTfzd4tD7WcmWkP8MLVZDMujHF/9Ji+TzkKiosbZLKc8BRvDBtbSj5SDD8kLg/
F6JX7H/5gtpi9pLAf/WlRG5XRm1ZsPvV2/yzujKsUEiIWsTO+EpeBgac7XULsXIB
hThBUGz7M9xy2LaxL/f6QDpq5VkZppKIXs08vKc4Nz4fwTbjrA7jDhTAtXUuqqjG
Q5uIGhk+QAaJrJ6Zx0kYZzO1NThVHmKl3aInUlI9zUJ45msmM+7f5/HhMyyFm9o7
5Degggh02uIeWNTKxQUMxLXcU5PIxnJlPMGO6d3oeyB6SEG69YblS6LwMUlHfH9N
L0SstMW52JCRhP5A0joiQgMmiXg+vMlHNDiUqgKXprt0QC7WiI6yIB4KFfLoIKo9
8bF7Wc+EfmuhBmODP1GEH1+JFt5zQKS1TX7u8euxiwJv6b2Z9AD83pgPFzmHphG9
HXfVLKpQtwEl6zbnl1IkQiAI9uG82XStkb5yem2nnPGvFGznLNg7xXWCnD+9v6PZ
dQZoonjW3UQ3BxWhKlVNN1rhUzJzOc0qFve/nHvCvc/rqIy51VkN+PwB2/Fbbt1A
3g7ykV4jEEs5Putaej7N6wpEVkM0r7qHFPvBY5dR+BaGX5II0EdmhuN41otatTC6
Cw4Ev3YFuhcrTfBWgPdawYG+yaebNsS/QbWFGNwaQUR2GRdXNceMAB2XG9X+1kkZ
iamvsP7720AFqJG37EDUFXB3DhEuMcdr3WvedBC/Uj1shqCAOWP5sR4jTSSz2LAV
uQEvkCpo4cv3D2si2G7yv++CSM0meNRJSkKTyfHpeRvzf7vOaHYcrS2bmcTEQ9we
g34PpBp1O6IDRilTqR8wufF0oNBs/+bXylY9kM4wgSBlfAJdOnVKaE+Bncrje9LD
LX+ZY6U1XC6zztSNZwE1Cgb3dKo2FjbDf/zjFtBbqCxN86foI2C05jQrCWG7N3fM
Mlu8KxSAhfs47TQt/JgRygC9XlsfFjl823lRyQU5nXRvMU+mW1uuO/fJhYdV2gHh
jZE/U04jwRQ6d0HnwY5odNuo/t8rOizsbS470egJp+B6UQ8fQIKMSqMNN4UZcsxA
mNaOilc3KE/Wm2Z42ArmDxqCKfFsBJoyQkm3xNmPFkySmf56csKh7/u/gGUp1ilq
d1vcdITtR9Q0D3N/CHlH3MWr+dgqAtYrMX3tioLPLo5zyHJ1PFkBt7UAmazNAFsn
ulPZPHvJJL47YeCB8DeAIhcaDTVsYPhDTEp1+72HVskDXc+1CS0RZDtCz7R0wjtx
nOviqVvCFvCbc+6g4LiDJfBHi6DLswPrzIUzeGr4igv61d4Cpk15cLukVjVaD/pq
rWtBiYmyOZjw2LMqtJvaCllax6rBhqvvTv9nndqD0SYY+Ri/7a+o3ZMFtSVJuOcN
sC8g9zpA+wWdjhal1A8m/ncA3E2C2LJ57+hIiZQqQfZnEGNILMaDqPhxxYzTIwuR
8UkmzBLBtevtVorbbzr8xOJEcIHQSCOO8DxP4mWAVHWAC/wK1iwbn/BUWR/ZDzfe
aeKXrErRcXx+8W/8bKGUAryibPJVLRPgMTHNO31XMMPsCd/kAk7+peVgl8pgYD/I
9TI//oGI33IU42zx3Q5qV1JjT2LyrlbmOV8XYbtjLkliSeSLscCBLbs0NBDu6adr
/7mStHKc/QKFGb7hf19jNDvYFYr8aide8/Rz0Ad/nXw/6f6C25Nc504hckEhM4gD
s1qpLp1JqdPPdvL9qaAnlG3/1G2w7sfC0tPl5LqYccErEHQbve0CruWV/2CLt7IL
7gMlmNnvoYMur5nJTf1K+H6K23fj2Wmty3TcG2Y8C3k2gSph1qka2tstsrkV8RxM
CKv+WHoFdNKVXoiyVeoWm7Wttp6FKLmv7recbARet9tdvEqEYGT4vSbxyWSKDfFM
o9cDLl8V1GtyDcxcyMJzV9dWT/W/d3T/ys5YBZR8KXq27bw3DTqKkyxalPB1i7Rk
mrFhIZ80LkvcZAMifsz4EwtugFsKtXmGcvV2JW7rBgTPWqDM4Ng+uNvZRYfcjHhd
4ltM/Sw/4d9L27nM6Ru+fcTL/eGGVhSCvK0Tljc0ZOvsIcweG3GvFjBZLiaXyJuz
Ceo+v1WkOqYXKPB4saVnNcjVF7DljFbutH6Ffv6N4mxPOrhjwj8F2NYwNwZzfWm0
Lxem8UGAOxrhuS0/T1X8gkxFUY9JhUlQUWfg0K0fXdo1M1iIk05JJyEpkxKck2bJ
joJiJh4h8aK0aER1sJmqCFv+Tgo1+nkMV3+Q5v+OKus=
`protect END_PROTECTED
