`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O3k+gp1WPwxczfRSgvZ9d26sNFRd3W6jnjeeHGLgfkKNuAOEz2xwHy4FuDOSUrrl
DsICTxzDZZtb62Jgssr+CP4PQjGeNfmxf0t+A2ocBIxaA+UaDILoxoUZ8B4jmRQg
B4KonBo9fmjenlLIuFf6LTqOGZS/miM0IQtcbukTuJLBNH28yfuEMuDsV9MpHIr7
hsIcpB6g4Blqk2um/+iPfXOhKTPNA0+g6Yk+CpITB88hTgXO3PDgavY/389S2b4c
csplnaEyuxqTlzTb/uJ4YEkdhO3nj6/Y1SsiXdzyK4bDHVUi96H1PajhN/32sAy7
xQWNmDz6ZLPP88Qgwck/vQ0NWOxBVfs3TNXkA1RmU0wbAGWKFUjQ413TmXojy5In
XmW+A9z+giVme6yQbzfKH+CMSW4yjqts4ceqagnwcf3BOkfIOHR8RFDV3aQKGEmI
vYkyI5/PfEDDYOSksAYVkY2lyydYlf/LkwnymvRIpFBA3RP8a5silO4jvGaJ7KUq
`protect END_PROTECTED
