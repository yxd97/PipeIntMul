`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JuiYBaKNqbxUMzQ7rzAVFmN0AlNu9yCYeN4C2o5ANHS1zbMq/jg0YbLoGGZPDrmP
UZmUOTkzU8+7+V7M8/naatI2dT5e4sw8CnZG8+7Q7b/EuTt4LiLItDwlwTLYAvKS
ga0vAiFJrX9AclA+LcAPz+xw3XeW2jRnG8iAAsM7GhbHozgm5RcmZbRTTy1BKnm+
n8p00Wqu2nkM0BDzwWQtL2wdxlPlzjp3WUQHPc4UzXbLDe30/LDSKe9rewZOvMhE
RDArYf6SzIML4OJEMK6jaHTFQpXI7NIQY2mo8yaJ3NDwhGfShQvKriPKEAILiqlN
/ZGJkkUzYVryQv8ZzDfab9Om3i+xievQ2M/C0g9rwwrjtFmuQzwCURR1QV8/lZkm
XMwkUX3M7i9+GkTKo0BZ9Ws8I8DPkrwf8ZXEjl9i6/nYlR8Te88pkFMqvtF+/fhs
wt9oaczKi/QlOUFRdiOH76pa46z2Tit7jaHhD3tdwCuPN3kRfNc/dE9zkPDeiFEq
XN5vvwvcP+MhOBj5OZ1j6MaDb1NKCvgfdNiw2iqFmraXsX6OYGV+4U7dC+rfPoAZ
6AY4Fn1GhjOTGbFkCHR5Zn6Z+DHIwOobh9z2p6t1DHkzC8f8Xoj61/Hd6I9Gj8oU
ybMSiBdNs5p+5WNMYlWyOYCGWQSGuDQ0AcPa3BvAs0f7fOT9dUCbwBzu0hZYLCJ6
AISTh0SQH5J9L/W5LmRjNaH2bZyPJEnXTgl0OhTtN0u8EqqPV7nMvbhntvj+zDK3
VFkKfQkP1u8Y3tAzrAXXn4c6OVbQqLTvtWB754IdLRzC2gAYFNsjgmi+TYGt2QEb
GWOvSCVlVvtxf0/zLOCdSz6K/tGo4OajrQ0fF6olf0QhF5JZDHbjb0zzwQggrHKD
Xw4oflF11eNjuGePjF1U4Oixbkzt5lo7Qd3B+eBrlQtj7hqFb9VWLupNxYi17nO7
PH96/14laK0b5ezABcQjMfa6/DdHOBuQxJdyLs4GEfJxC+2D2rHdDKQfXadNXPbC
IgdJu+XANH1E6SgfRi+KTOxtI3hVigpEBVmmekbaRQSuKzRys5SfMYzHcNU6D1Wa
IqbiB2chSJez4DXxaA4PsOOqiUUr0PWF3r55eSt9lJlLPdfRUYTtlaUOyMgO7ihy
gIxvZaW6mkfxa2jRdd+XsX5Iee1yla2lFPSsjXUKEkJK7K99MvZZa6W5YfMfYixq
TChItp6pG64z1muHkpYgpSuHmTZ7BIyE3xr8jE8jdhP/lQcs9hjfMmpAqSTFdlhp
TRwssGt1N0KMJMzful+3138B6NuS4NYLulTLkNYk4BDptsPYDCw18qFqg8dMubUu
1N0t3CmtrEP3O1ux7ucEjXTG37YZLouLFfO4mnEajaWlVEPtVJv9b7tcjYsf2wgz
Gymx7wSX/iV94/QpTB0UTBqmn02WK9AB2f4ksfr+A4DRWa7Gme37i7hHt7piff8t
WQZU2NGmsFwYqdxB0ytr5t66FoCl+hPKHkc0CxlQ+kQbr1iXccp18SsATbhrxR5i
X7wPXCg9LfTzsJK5obp4KfPMLDXoNkvHqvUg1uewBdvYUXi2VaI4cW8vZz2vwmSv
degLhp6mxVsKmYq79RfX3Qg8nv7pJzzsyHeu56EJn9zJhOTutc8DM8OK7LIjiubP
Len748CjAIfZhakLKnxPIxQviX9GW7iGojEOj0CH4HRzzf9sarHs37ly6Vot5TFR
NVAtBliojVBf0ABB9qKXDSnNi+zfmUWkrfDSLQzXVMKeiCkoFTxZFuMv5+2jpLM7
9fcE8Jnx3HCxYG5M3GzyqmHjDY3xhUmC6KMTaQCrpp8tQe2hHSIHGOY/mgcvXb3z
5QAWQS8ppr6e6P4smDPSRW+BWzLafbqAo/C8uvNpK+oAo8WTf8M3dVHXpCFoenWD
m+nuhHdr0v3GSIHyhZjQLXLsCyWBeuHA6c1HxDirm2i63zcXcHGFvSD09ekOX+Xc
CQdPiaH0j692AZlI7QN64xV5czwP4ws6PNCsQJwkSyyvCt1eQ3ne8sm1BY3h29zT
04hsjQsyWqcACW8BmzqUHSEGcdnab5IlVTOXko5S/jCr+Mc6B0HhFmhs/ocPRv3g
OYTr1KncUlgpzDC/suz2LBXMHAFBfeV2mB1iEAZErEoQ0UpMyh7Y8HmIDMTaJCnP
b2sUUF0+yp7sSN1g5fPHj7zN3fNxhIbuKRT+Ts1EpwyyInIaZt707WLa/GbM7HOI
zeAKqHJ8gM2+Wojo4BuSh+tMQpi/qBtka+5A7Tf8YOUvEl+cKTrCnnXCLeHpPON9
jY1lkFO0Ptu5majijH7AwVGJEAU8LlYwXnxhMkqwv2uDh1Yqwwm2EOuzop1iqZmY
Kt2yrpNii7VitoRXkU2y29Uh5TkV9lCZtPoSepDLkFwYRSMwz4u8KJGD/gs33Qc1
dclD6enZMphMmf8wuFfY1c9BGFJuTmuPEpeJlpv9yZc5OxhS4kJRxkAzD+YVmXPm
lVxGJHp6z5crJh/BlGS0Vo+2zEcPqsLGl3rDzsvcixYqicgPh6CknSURbTOl9lJO
Y31odlkMjDg9DqNyp7tiwAz2AOFhBsHpG5xqpK7yEk5OyGSS1DqD9cZZYvxs/Qd+
iZSUDWsR6EjroHKW0+RymMHC/ZS31TFWtSKVFEU1noyoD33+NLu8FG5oszzgQs/E
bQROgGHz6HLBg8P65j6N1e5nX/mAXOWEofQgYr0qQMZ0bY3EZ4vF66QvLp+YPnyw
BGI+nrfEMIvMRaRoFiok7Hm/vOBI/1vduRITPnYcC+PxI2knhqMiGhUVzSuvE+Nd
lZYWyqLX16D2/dcK2Mo84MLbE3NJ0AT66QmCMjBALDDQ7ArEnQxDFrl0SYxodl1R
+4umrcdNL6wbhqAM3Dhk7zRxYEqwMcllczRdI99iy7fiLyx30GeW18vH5H1rBgGp
lMcMNz1x1a9lLeEEIqlfDl0YBAT/7STnmyW3mOWNg9PEyutVU0hTvtH6+HON0Ou/
Cnm8srp3BSSG/QelC8CebdE0E1KcZNBTn/B+dgDmyQvJpzZxwHTfK4f9/yJMU2ow
EgsKGYd8rnaP7kkZGQklD7GLnLLcvtvAxWnX0992MXIIStY0rRE6eeQUcZ5gQ0Aj
dr5+41dKDNA/xwjTBjf9re3XWEDHXq+ebSdWBO4w0yHJJw30PmT9zTH/W+X/Frec
i1jT76oGs1iZwVAvXvjHEktD9T6Du2bNYcQ2KGiPfQoTlfA3Lrq/kxHarZ0FNnsh
FsdPCBcZw1v7KMw1gU3l9ryTSfFxJOFVNdyMyzzT/QpIgHSQRUbqPdvQtZVYyDk7
W+u7xBGuWQJz91nBEV9SzGFYOb1jnCZNnsnfUm8iwR8/nr8wikRKeALB+4ACZUea
fZVfIKO3SKPxGJaPlOsKMKcV+UIOuSgDa6WgPrXMeEvU2b/i+FHN+YuHRVKDP9PA
6Z0kVZBXg4A9s3l0jp444MHN9FuydL43UDAm99hj+NOfOZELixroz3TqegYvV/6H
6k7qGF+2LaEef6MCt53Xv1JDRJKLCVmQjw1xZbguTDyTOr0L263FMCVUr/12ShiG
MXfivuFR3YKQDxre27oKkSc8oibu9tDRjiGtI9a6Y6WtBr3oRshdnBxl1Z/AqUEx
C8U4swk9Y0S1kmVFlawze7tBaNH9osRLJSVOu6LBSMpqI4QHu8qovUgc/cICRMHU
vNc6b1RF9tuxcbq7XBiIdrWlTUCJZcw2DaJ++TksPqRcxNVuadDGBz2lYSSu6xxP
t6EZLjbhxW1M2oKJxMMB/mHFs5rqGTFGrYkgIOPAjmHwUYw64/HePjkFWXLNP6P/
cBVv1hSzvmyjEsnCfqaYP5PlNk4Mf9t5kG7VIUO5XaiFfp4CGXaSPSTY7RdmIJOi
txDXcfbJ3Umw0RWOrzmixZuTqyK9YQ0hAt79jMTHWhuzyIqM9V4ujlzDaqku9Sdv
VlbKMsB30ZDaWx4SwuckQV8fCldXkSl6xxtNnUsFj9A3lBG+CzBYU8NKFGIzVlMr
Bl68QIJl83RTleNNmsVsUSmrmgQBX+lNr240zEbmvjJYJX4qmxwRIz61qnbXottx
evIs+zqtVoLecRM55PgFPWDGr7drS02BxiG+fPkE5uxri4TRp4GBiTPU4Fs38Eqo
VuoCVJGpADX1mTEAP6rXCZnVhOtCcn3dOQOBd1Na4Bltr9qk8fVbi6cJ2h/NCq12
+nEtzNKz1kszro1s4WMB3XFC2kAKzL+WHeB/DU6mt1FayivV1q4pYFY8BBtzTQxo
aU+weWI9yz4Qqu75wub8GL6FG1iPP5qk50k62nN6OwZYxnjDinKqQCv39mNGj+Dy
yqmKmgM6aNG3SXjLi/pu1GNwifBkTgPzGVaj33qrOoJ33WBKAik67yy6nJ0WosVL
X8QCqg0iRji0RKjGk+3cJRRzYX0LSD1J7hJbfFKQugL0QpDTm/2ecbEYW326k451
JqoXdYVGEyGaL1gpcVZ06iuIMc/GwA30GeIkOX4MqudV7pzUlwZrItHlCCUarCq3
74YeyJb3tYxKckB/iACPkvm7PqgdStoePJWCJw+JnjD3DZ8oZE8zeDzWMSqRTESa
ZWOyACd263kkNH+rvfFuvkO5TORTms86BixSNurFNDS+p3Z4yfhENP2acYXRo/+R
E4BSjPibj/hEnxQFinH14GR5c7jDSwcmHWdF9RjxVJuALXVeUTvHlAP48x31J4At
E0/mf4dzMVHZ+j/l/oQPKwFxouyHTyhp21gWGHzA7waPXsPmVjNVyK01pHSJr4E9
QjHcgTdV3idY9a1Nd3fRtEDMwKLxcxe8v1wRoJbrkI3eVm3t4uleHnAMkCOl+e4i
Z4j1VJ4EBHx3t9BDIg1YuJUffobVp/ibyKJ+r4vA44muxBMig92yBiHYfvdKaEhZ
CT9ARCrvGLkDncYEmyFQo3smMbZcLf75W7X7/0LCJyPu++BTpV0E95Q1grea8/+z
iykv5E77keL3TC89DfrB0dA4YnltQKBpKhgpnbCds91hQqUzY/qHoHUS51si5mBz
Qtyr7/WdrS8gPTzK8shnzkxKElepZEJBKcBCan4zM2lz9ble7yhuQ+EQnGRj4NL8
TgnlK90As/tuil5sPSpuEN6RQUW9hfq+CdHQ5OXBRMHwni29KVs+pUPXBi94xCLT
Zg03iMJYXFsroO5XTq/RbPQZ6qFJWtUCzfymmKjfVyGzpzb2dqbTlIY0HYQWMYpy
qYcHuTED70aGzqVbUlFXEDs86fVtcscELpI0YC2MgAggd8wJeK5CcvwMkwOxccze
zYv4TewBmZB08ZYQoyXRTy+t7I26hrKdmdoegO9whaDdY31nmsQeD4Am2tTlSWYQ
6TI4DboK6ieUhYMuCm5/qqEjDh3AhgxAHiLo65TjHJVQJvRW51e/ICuGhO7Mo6j9
KoyNFdNFVV4f3dZwEIFCgKazNwfozUg30t2qXCTqw8b+QUGBPCrIOR/KGzyS1A0B
JEV8HI+pWgf4Ca8k/3EdV9ojRckjwgEVWptggg1hKv5kJFlDFOGYt6K5whd01b+d
hPEkddg+ymb+e96uNzILfdHSx594gxdZdkFrYJIT6Sppzx93vT1jzwl7GADO39dE
ybdvx6jvGbnv0Hl9hjn//w+AcctrUwHG2f3Z/JFK0YE2rxpO/XqOy+in4h1uCL3R
zslPabOyhGg8/mJfbAnbx3rrlZnuUQofvwgAa/9GlpDw5Fmsh+cDHS9epEJC+elS
QxJmzH0iunXBXgdc3yIsFShWtfdIsDWGYKrtnWmF+Wy95P7nbxzrhxBwJ0C193DW
4md2ZsEM5P/e3YxrdVkG5SHpbJ+M7QAM5Z2j8tV3P7iKCVYkJm1fJnfm3m63IUN7
09X3qYfNxf+0LQ9E/S+MqHZFmA290GIICpqKmBYQyUYbX1ZhchHuBY9LsuhnCzsv
Em1KGL9rmUsIiV7Cfbr4BpvHm93lxdQVLhEvNzv2AoQEyLy4KMhIIXthOPELCZcI
qw1ouQLG6DCCncsSbtvu80gX2ASRjbJjVkstgYQaghIhnM/c/4jFQqkanw2WnPk6
6bEO5YOv0XzQLLTRE9jkGjG5YAbOsLMbYlj2ZW0DEQEOc33RWN+oFVkzZSYAjR0w
NlrqDCaFb7ksC+oc6/7fYvD1zOhDjmVdgIukcW3FPh5G8p7ZvdiY4pJLz+/EEGkr
BuuHpnJ02F+nIR/ZRJknhjzDqfGf3ph2vbNDVM95ifvwX6tYeLxA+dfhPnLOT//H
I5zr0z5Hdbo6heerVOFRG8iomrdM0w36H5AdIezKX8vGB9GQFEYKWS5j3z/deW10
MGfEtzdBcw+K5CB4kimax5mfpyWWkQdZogcZyp2dUb97qyJ6uUi1X5zeZUBM04wh
xV6vwNlB27ze52dpoM5EM+uvyv0Hytg49REoOVmceSaNsF/5RUtN/hNRiHHmcPYs
jEEY2JcU0XB+vyc3HnKtlVMPx1HBN3ldibVAC1nSDgwasuvTxIcHdDG94Ed02yfI
YWnwLJ/N4Am7E5RkS8E6SFbf2XqPcN5MbPpWCTqeBwsG2VXxB+h/hxdE0giOODIq
zmlXk1y+DBJ/DV/K+8xfmXQUjrK5diI8Q5epg1BfcvwCHurORgmNXjgITqCIGKeV
ucRDjl4ap5QtIyrMgf6Mbx/m0KxCB5pT52GjzxlXxVIKeUHFL6q7DW1kyCYmveVf
qgT4e7FvaKoLpdwb89Nuwt1hNex+oQhdrvx3GdRBz35B6nVHrkQAThhdt0YJwv72
HMVMPiahploDPNvaCu3AGdGYjjrKZ0i83zScQSMRq5tGiBeFo7c2wrCLldAoRKJl
qGlFW5bDEJ1gyyESnFAbZ3PB46LlRr4s0ZVS5z4R0fWhnvvXMguJ7Z0SOs6KhGrP
nzPrTDw3DAe/wA6g2GmpHkS5X+zZR9SGFc9+ZjnXzanXp0Q+94jy92uAGKW32C1s
j0WmgmOt1ciyilUMFqq6n1IvhjJgypuEPJvYasOWm+/2QwMH8LPUVpffNxr4fzri
5fJOCp7rt7bc5JpTyV1XtfhqaIupySqWD9hAoLredAD5FxZh3NTKSRhvt7DLNYuu
92o2uPpCBAmoJQV/V0Kha6cjredud4CgU2Hr0RtQd7KfNE90z8/X+I2uHFmWVdRK
/HSEyE496zhUn1bBzFZIAa9RB39ZsZlNE9e5gZWRXg33Pebh4d12WpI8mf/z6ih+
f+ExVM+7B23kZ5z7ZTsSsOC/G9C0qk1jMn3Q9wSrzR0+ZGpyzpcnyDlSxUD+XHWf
HjqeWGD4+mVptfSRogvUxyxuz3bTSmtUWxVMMb7iMP2IeOdSeB0rBlOrEOhVf6CW
tIniLtCcV4ig//JwmN64Z3+xAW6SDK3dqNONE32SGhZG5HyB013UfRRCRrRIxFOq
7SGUj/8ZmrgMPIiRJyocO4VQg89HywgCN4xcTKbVx4Ula7FpvnhZmZmAm79Fa6RG
lVOzuXwegH4TvHy5C7xTv/97UKTv4wOjueOmJmrxka03vgDFO1fQAFuBWFePijnF
Z55yIMU0l2KSnLaWAdskVY+/WSp2AaRX6v+cZ5/CsRU1HAoTpMgg9IeOuNxlAsnT
BY3UiSAj/5Mr/B0bIxwBsHeK3kemoNmcN0F3JEWdux0d5w1d/hlav+odqTnV1E4K
GGe00KIw8j5ZToRDZXbqhxzsTs7+NO/sYpw2C0UtgbhDie+QvvashpW5Z2FlWH45
WR+5snETkqXcz0U/P9s7HUkqZtmqW5npYKb+v/CPaSk/rqRj0HPYL8zqmq4ReCf+
uOF0YZUJk+/ZngEudbqLpR6EARksEXVyKFstewkwL5jugJWpTsMoKxIFCHNQvhI+
M/gfY85lYxtdjWcqP7Ymy6mbnTHpR/rTg4tU9VxFVMBCIym322QZM/MO9iXtBBWE
t+C6iNHgjN4LSw/F4xG9FMaRR/H/IHsAPsk69z9n4WTX1zP9XxMuKs8f5Tc0NN7v
yUKCnM9/SLE/YyMVtHucH/mwFTMZyE315O7Gqbb7m4DcxASAN04qSe6x7zOTByoX
BwH08WS2KLwYc8on7xlohd6Rwf5xjFpiaZvwGG/ZtGXMZoaUoSoT+7J5kZAQ1VG0
zjGRgr7zhAyGlze0knGIcXwHEF/4zNwMsfNj7+OLaqx2L5mTNIwo+K3rHmK4TDdI
2l/ixffUUaZR1EWqC0gErPoWCSHwltSo2JWDy6Mn8Bon2CFtRY1FTYVdb3nwcgAB
PK5UCLTFeXA1Dvul7zIZK3gJfgxJHkb+8fY7ElhWDvNdqPfzksqc0LS2rYCEsff2
gd/ZTKhnyd/kWoIzndRywNHX4BvnwNtMzOam0A2fOhD3JDqLnBXz8f0njby7O/Gb
N3txGp7afm4L3rRODFzVbEnlYeUbSqCVFu+fsxaFY4nNiUkXblk06eZrx4gmUoeD
bMafVwi8L6bioQl8yhNyTjwx0lpZn6i1qY46wYZa404tfH0k0i9VWbY+xk5gCfIp
oVjFNOfC7ucSeaczfLBU2AzXk9EHGj0WXSZtl7V6SA63AJMWopMov6qlR5kfogdm
jSjsyfHO74lpvJ3cPyVriysKLRfCE5v9oV3PYxJvztGgW+VBzods1CzH3uaBfeog
FWrW5AFaELbMQKVRFAYo6Itsqtr0thhKKVEsmkX6pnIPgKJy2h0v8KCnLsd1yzVD
R1RNyIN8FyFdf7cWd88WzCNU3YUNNLidot9NP7XZ2P8LCnO1lkpkiz8SBUKYigso
snn5OIxO1Yc5FNCM7R6peHj8Tgvtp7sJem5TUxOasOGLVivyzYFyu+J10TIhhO+h
bByKOPyWIx8c4TdWnkMgJHnkkfKti0PcQiVs70hVq/GDvI0FbVEIiAsxw+97PHU/
zRkkomLVixIkhdBps6TaGCZQ4psLTEm3kD/iDMvRi8EG4qRqpad08TrRwCbsz+8y
YqEAtsV3+oLeVlRUpS75RrfrZdfEfwpy19Bn3wZxaYkXSCh5JeRWeFI3QSbPVr7J
sQgmNEhvHolWht+rN8zsjt6vSbGyA/hFUhAabkzxtoerWDkx6joLRpbFN/bcxL0S
JL28bYBGlP6YCSMrPo6G52Qt2S5pw9S1hhC/R7bQHiRhulJcY0ceIiKe5xrH7Gwh
dnoXJa18Iub7wdWLOws5l0ZTim8YOFO98N6n2xM1spHrZy6U0u14qhZ9RnranXB2
3tDBWK0IbGXwXzG+Qt3hTtzjknqXN+RhoYYe29F7KpBJVwlyKgdviPJSzS7p64JV
8Mfb53cDXpM7zMhreaJpVXrzoM+XT3maqAKPjj9XgbtKIISuJyMrO0rU3Egmb5Mc
0uVbNZ8b3R8LjkhlXyqcL7PbUdE9y5kEbhgWjnYnJzP9o82zuW9Pf/KYhJ8jLJGs
ic1F7QpCimg2r9O5E88+cfJ5KkrJhY/1Sv/q4+fn+lEqpdVXTIQA8apjR2l5AUgZ
QgQbZsVZhdwf/ub+DR8oo3q8n4TVUZRsa+TQpnFJXEoxsAvoiNkyKXSoXRO6m4dZ
ICAhLh5r1P/UNjMoEfD2mvqkamqQMolVwiyzllpd/vy354GtjgG9VKEf53Oxtywh
ucZLY2H4s+O0p6dKC6UkVnko3Ll7CN+OzwH2QWFM1lygzM4xbGTBM9s5VejfOkHQ
o6ay+h66/iMtfwh5/ycu41sBvMpr3mpHSNu2JCls5sOsWYbcDX28+gIKd3nk5ylX
IJMr/1SLgoe5eTzJGmUg5YjykCHCcJSuLMpWiESrXh8r6OW6IjYcRK7o3DsNlnVj
cFIuqerzzXCbcOa7XGabFdYKtOjTJQjQh5/bj4xMATICKYRfvHThH7aPRXHiM5JJ
Q4i/T+6XcojPkxsv1QrdjchhtvBdmIcUdtobSTSS/5JomLv0csSA0b1LMaZyQ/Mj
QTdWEuC2T5Jg8V83FrxLSO4weAeg5c5xtisaIqZsBj+2snSqZ94p7+bFE4Zqs0+n
ECLmceSCnabBeXNufoR3UdCKgBddj9lJXOADtUW3hfzcCpZOxPCDvtXqNW+6jdYe
t4OQSWIbvxwvhcxZ5b0dEbtdGanHjjH4M0kknmc0EQOHQOiu2+l3qvlL3Frk9vlY
wp2PmjFWaPfyg77mbvcjiL6EGZfSIxoV8rx+Gm6hb6jLov0pYAT+URvdS4pN6BB4
Pqwte12N+UYejhgGlXhKetjmROwfKeEj4EMQ3VqOUbc0/ePFqB4dwXDGY1VZdPF0
equjIqOk/zYqaXFyK8SEJjHfeuTqXXmEgMmNFLlpmhruaNmwOAkRXv3F7bXgOmnZ
8NVM+Bb5uVgU5aDyJtptSxz3/K+gyHRepGyjBCqUpIWZWrB50bvnr0KdNXPGZ9jU
Bhqm64wCQmNrOZRfeGeb0ppge4iRboYj0TmvunwaQr9p4o4afRoYgJx0EXUxwLac
UpNd+Q/jYhKyiWFAyWHT2w8nw+3cR3kSUS0gWWPkbwNlapiFYNiCS7aUWhmUwIKu
lKx2Rho3puYVu7WuLJ/GMw==
`protect END_PROTECTED
