`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYnrLJij67Pfcgur6bIbF2B/hU99+3Vi4Dm+ymQ/pOIxqzlPF6YwDrkRSjNFulas
QUmPL3fEDqYUNCpZw4YtZjvomOQlgvn/3y98PQrYe4C+4unJ2UkXeP42q1JxBHQE
vuT132rFEkpvFq2QNyVOjiAI9GIejCFZHK1A/vdAukmMtNHat+Da5lDEhiBQnM+0
e9wx7CPI+2LEDXPAsOrodKAojG3O3TizGuy3uX1BxF9+wuKmvrYF9dLRqeUDl7aW
idHQEDO0Juh1oLn/jUaUC1/CXaXU75VY+obTrIoFoViI9cVMxJo3DNb2lbQRO7ZG
ZIM9e6G5ZP3CiOlpgJuklnQRlCKdvejg8lGUj9wadJdPy7fucMLncQ6irYTvAIqu
IRopIlr7qCLFntuxpJAD1GJs5UK0q0Du345Kh4/zAVUnlrw3g5KQtBRQEGxq9sjj
+0JO39WzVNsgzzk9PdNCyuVKXG22PHO3GDtUdp+po0v0XDrfN0UuhB0tvFHbysaS
L5ub3zWjdl3mheiZhyPgO1O1MIU+EAa/P2p8n3TZim7knGCxneO4KsES63/vBKNB
TSQaPKKGZI4ZtFttGJHk0NmalMOf4nTSerwzdKRM+zEVGnYsK1Hb0FpMJXKB+Ugg
zpCOQNCRf5b6vCv81YFsrH1Nadj4CpiVpYa0+Vz/WqmNjlIcjjL5XBU6Axv8oHjR
Mh7ec7Uq4NzXKW9IvoKvu9pM3m9Hp+hLIyn06vAqzEnlLrsHzVgt8EbbS7/ww/0F
7N2cVbvSTMoDFPqVJYJypTc78v47wh2tKkv1142gBtrr2YvWJY8E0lQGV506NXag
deiYTHOZ3F9WRFxCDVWgn5usLSlpMISFUtB0tQsqzQOQpffh9q9woQuZhq2czWal
mka6zNfXxhb0sgpwQuE7FAXOeE+bOEod2o93WHvFD5bEdaFCMMtYiuqVygk5t44t
BMqVAQb9gLAAFt0Jha0q4J8bD/XFdWlNEAVHGau2I7YCalRIXvkqhQfCCQgsAgH6
Nlnb3e5qKqIt+UIAcdumSWJYy0EToZpbfyCFX/ccL0hU6xn60hmyVjiOUXEueObU
RXg7NCkMMCl9H+8h1HsYNMP7xvicaIDC79Ctrx0QYW/SUVOVirhwhA0f90nPC+Hl
PSaxdjy3/UdTZ63vmO3ydt108m18k+AMLWfcF2AiZ5Inx+gAl5Jxq9qvlqWDVUgE
KqEubnG+kFlhmHNgld0gJ93tunuZQXFkzEoGN76EnulLy0Ai/GDUHbCdF6JZfCvW
hheay6WgEBIkGo466UelAGinMnButdV/rEBbhOYPSvMHmKy/JdujdBYFGu+Hn6TJ
4K6/02evuc5ggY07D7RNZzpvTDYcOhrWszY4Ae+BGf+xwGVV5/jx2X16PIDw0Ehs
3tA3obYsYSyiUURBuLTvkwSpd50w6xEl/p82NbzlEcK0j4UhEMfk0ymL4dUj06E3
gNLM5Z33dE5C0t4XcaIkDq+8HvzqQ/m8GpfnN5QV9VLwfKqpDsCmbBEq5fA7LGGR
zG/a9N/+vWgzUI1fZpBYTNfdUMIbnY9E+JMOuUmkS7l4kS08O95CEWSLUrN8XvdT
3WJL9L5hkyuAk1q6THOPzxI5L48TBS/91PHl+36c1vV5+s/ymRhIRuhFdJ0/lrL7
E7AjnyNyKqplA7V3JosBYJlpRv0wcJO7kaJEWAKF6k1+9eN7rhnnmUlRYmRIOFoL
6AgTbD4zeRF6aK9MAWA0+/SIoY288NLeIwLhZ5TpF0h/MnFV2d2xQrARhkBKKPtP
EZLuBMjnchBDzQCay+lY12w1QokCwlBr8a465H1tma8YIdawuz7Xrr8+pKMkHl9V
QEDMMfcHrBxgaF0ABHnqYDjmVcCppKzapxHQtvvvOb33VeNCQ1kopWf56hqe0i26
yDQAb1/Okj+lXdAkzmLOUzrXtfa3/V1EdypjdgqyaNoNBhxx+b5Z2jMalaL2RrY1
BYvAIkPm2u3l2wqUvL3r9KH+3IpfxM+JVNJ1HaTz7x8=
`protect END_PROTECTED
