`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D02qDBdF1dmrUxDNy0nFmG3J74vgkKhQ8gRl2tZnlAJLusLXu29yEhE+xnjEj+WK
0SK+5db89f4C5n/3EOG/rHFJFqEhnSTZtyM9uJ+5+fpyqCiwREnZnPWzUo1ZsExX
lTziOjIOg7Y26JSw3cFK4cBjLOru7+gJ7+Y68gTJ635Lam/rwCEQufcOvGfOA1IS
1ODLHOmBf5TuCFLKu8fvecsUWTiVHDrXrkVMYt/VPKY7wca3otEh/Z3jfQU/+D9h
evOzk14D60iShY14yST8tppeAzMHS89qC3SXki+tzzHnXdwOgGz7HSjXF5ikhN0c
jE012bI1RFFet8tSPeCr8xXF7QHjwrTylWwsczsEm9pBUpkwXJU6Jv/PZivlZY2v
z9SZE2vk6w5S+AUu+mdzFWBfNkYnYzQpKHLewaJid0A=
`protect END_PROTECTED
