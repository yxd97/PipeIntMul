`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uwd5Uu5dcDxWD2vKoa9uLj751+FDb3wPj7BdXzte4Xia4tkIJxVhnm6M+NJzJElw
svHnSjvj4B5f+QxDsAj0h5vqheJaQp01ldVWoBDRRDS8UDBt0AQUXAdM9lywe4Rq
Kc5gezE1mNtO0yO3AL+Vj7AY5fKGJtmzFcAMd4BIfes3fQB7L751YB3dx9V9JeTg
XG1TFH0GrHoePO67qJjJZXcBAcAZIkkV7NGPehWgqTNE5hDWkjMX/0L0eh25E/Eo
KkQdw6eUVNjJMO77/QVb1+Pa+4a1UWWD57G6e896hvyqLcqoosKmL/ZY3FCGedGc
lfKMCGGttJPqPiE4LXay9xyWYGzeVnc/qr9q/lAO5ffyYpHl5orXPno7grKo1Pxa
zMYq6Kj/aTkNPvBUYamy5wJ5czkkzHgfGNhHesJwqq0FbQlWkIW5VtHBGIcFnAoy
kiHNorTZUqGbJSghOy+AFAwLOSORQc0TpMdgdajBIGM5DhtCHcCujaQc0JEZBQTZ
2MEm97Hh4WBK+q5EUPCpLPbpqhXYg9f6oLH8PajHzQ5Ph+asalgBfrQ9nk0X3zzH
`protect END_PROTECTED
