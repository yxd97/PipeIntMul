`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2a6487Rd6MLXOdfagn9dAmfuXzCqokW9PjuA8E1+5hUiQMHZqqqVDywiQnmCzDu
FwO6v4sPx7HjIsMd3EFP4odxQpncJmWU5ldmLP5fRbYigLzUQXHFi1WQ6wqUQWtB
h+x8dYXl4mDQUOXDWzDCKF4O2bu4JOSAErlm+rYjnN/jMbQGQuZTb9Dw/ZQEC7re
J2hH8w4baJvNZnyAtHFjCQqqD4ol/0JvlhdCb97g5iMNRlKaIqYZjU6hp10G+E0q
+q6+qutj0XbgUxIwX1o6yjomXWFLmVy6pe85KdPpyHOs6sE46ET8GNsZN2fqRvpk
f/B1nH05ieXGnmj2jx2loUFXaGEe9iv3BdaZZddF2mUXKXlo/1It06p2v4uPD6z1
uZSfvBeuy9+g4C3fpKwyDqxczNI2SbWvu9tQuEiYQ36ksgLXqfPTIISKmIMh0VaU
CiLNOOMAAPAqRxa7jc2ua45L2Xyfy1iDE+cnpbJzLZDwW533GwwyHRPBaUtV3yh5
EJIDh5PxaSBtgDOQWjjdA9qncPYK4YZwW1UBgGiPnb8fWbGSN+vv/3JUX+9RHqMl
ST1BOPMcVfqja6QxaFyGJ2pxKxxJcbj+Mw50xQxVJvNLneH8cQI1QBSv3xQgiE2j
wu1XyAoc5l38LrjP5jUV7v3R/KUHl6T3ty/SyoefnA2rHm76zm/s8j0syG1T3lZz
szrKidu8CcbWm3gL8riRdq+J++W/8IJTIbVHWl3QL9Y8a3ByparJstJxCVFuRPgz
wsBaM039EhCeCD6jL4nRd5aIfvrsiX00aadVQr2Gy3B3aiv5NkMO3PxYT6aC/tQN
an3PRY+YCuzmQ7koqdMK+p+er621gk3qqNYus6rqCx+FR6+KSc+6PV3m2i/D2R6Y
oA7A3fdyRh2tHwDiat/L4XOh2SNvnW3VnD7hkfNVpmTyFPVwp78gE27y/VTR40QA
lJtsBCtqOEaTjwM6wh0nGzxhiHumCqu0oGX3vgH4KmYK2Y/dyT9w2zN0b9IoIzP7
F6eml3nTF/3IHoWLfrO8j0Jj87LHutAy/+9EfQN4I2c/GDBEk2/Au/tu8v4m/YbR
qULlGlzYow9fH6PImMTcVBUAjeOplbd9FUSIadRUNujkOv9SC7OccnZwGTSGEQqx
HlRCFSwJgQXbHuebKTwh6ulaTzl+RvL9in+KMCohBnAzw5nnKTkVMrTj3qVuriR1
UhrN9rsRb+P7fs3UVaW/WHIXW58ye+BSDY7NutbgzM+rjArPR0Ln8bfrI/4PSprJ
s4t5L+r/fI2J394hnL1B9xsIs1KugHaVNcrfqFTd+h6fE+6P0Pgr7BRn5LHinULQ
6UK0ol3CRsexwFqsbzTCHRjFh6t/0qxmLF4OG0flcgflDVz+VZ9PyDUqVXtMIBOt
wjyrkbhsU0pfuQTFIt/FAjBmJwO5rkZghAyr0l7Lsq7UDTLkQLcW02qzI86oGoZy
cnRvPhBNd8ZJf16poiloSThJU/ZlOIRjwvq3OJJegq0EeyymRf0k2M8iEB2SgGGG
WexuxVF+BJImUKOoVJ2sbMgFaqquBuSUC5HjRlD3Cwu6gUmV8D9gteOcyIkunNds
ddW1rBn7Nfnw5onfeCVRBBJhZN33NcZ+89QIyh2kIlWLRg3onw8nBXpdJ4Ws4HOy
mRxWrGutcnwJQgsL4mjkkNxCFRyPwVjh/Zy4TL/K9mKAJG7jkI7DuVX7k/HvQsV7
viQX8Dbb4jnwihEpsfn+kvF/thflmHHOLfD1qetKXG+En9dXdStGVcYpxQXm3MmO
hLfCW10VmOQOrYnJTiw/lLqvBwIvKjWXL6LxcpoPMkaeN3pamt/JKMhOpjOVd4tI
yXbEwREsHphYIHFOkn7dvXH6iY+OCPNkgjg09FLqGxyAO4IGjTfuBz2lDmEv50H7
gYJYmqTSFdnDb8vhMBTVBbwROxj3couT5T/HXP95e6lOau1hach8mSJovyLysh2N
RPD9ayiRGkVg7M/AeE5gnyJnqvAE3RQoTMJUG1dGZyqlYsTfm8hc5yaegqTgc6wV
JAPQkgCHMHl7EUzDVjrCn90qIwGvD3SHloQr2BnxOk/mK9Mt9f/BfIKczCSqum1r
GhihBhppoIp59wXOqK2gCaISbb8gIvMlf8aOE/lQdrWEQ4OTTa+CI/NroJ7mj+mb
d83S2GfqsWQsS5PbT2Ujx6UyTEFy2iTcZgXgjGr9BPRETI5qJc6WhJAXH005prWt
W1ogNxN3wQB7q6fPD93Xh3c7zG9S4EM/kwPqpg21j13tidhIpnGfcrZl3hTIh5BF
vPFQN9G6yI0Qhd0xzJ5aCkzvQST4uIobiou8f7pqZFjlNRT4CYLnR7ZANPDQc1Et
avAQupjh6dz+V9jRMVpljN+RznmtG9bAgyq+jnidnf+9HTK7l9/X+KNInU1O7K6f
brnAmF+JeXTX2TOYetr4DIUesGYqHv29+5reak+VNyNC9OZ9jyGAQYhl7x7/6N+L
nihRQqmnNfMAr9IHKHgR0/AqFYPyHKr/Qk4mLdjWjJ/K3s9zGFoNyEI0fulCq+P0
tesldWVMDPZdxEaIleXld59bChWikLXWvK3NB3BP9HZvF3xnBKCZZ4sM8D3QbkMW
gX6V58e6TA2qONgXFZjOGI/yQu2QrDL3xMjJwxX2UzXtD26HRoGtEebMbMBtWzx4
/Bw8NAJNw5NqU0/JS8f9i3HJdGbb9WIIMSAMKKuU1a21lhmqhRUv3smmcQCe1Zkx
S3GqZKDm73upJVT9rsDzjNJvCO/gZDOxixg0e4mf8UBrMnqO/6FcPmi3wink7mzp
eImBb3iiVGA8GKCIWo7HGQrRZ/du57rIj8vm64wyKzZORMuk0xx4LFhYzZonHLDU
ATeJy4upQ6pHMT55YXOA53RQs2b3mjfjya09ePUsqTKv3U6x6w1ehR5uYfMu6Zrj
qh7WmLfaYdg9+kdMX2LNWydpnixsXBsfED6f6jA7AiKteM/48MswjWk+LBk5l4ca
SlZvyZzTzwSdQHv+ZBdnMiinge+KxPPXNj5FWDAtuWQnh/qmxuh1NpxgdnnD70Xw
Pd2LH1WYX7Yd43h4pAmdByY2T/Bg064M1+WWGQaL1F26Na9/EM6PdRH3C+IX2ves
cjYbaGigT7h1x9xD35K8/oqcTJrUjbtHqPqSYY8QyDEgsjLTUX0SFJCL8NZ4alqj
aTE4qUB1diaGnbEt3shV0QwW1rK3ZGuq/ojCBP84LgM82qLG1v7CPm9dDcm7RAS/
K1juMkrxw/Boz14OOccZmTl3Gr2aDgIBkWSeP1ScEiZkvHCrPGdwgHGwJ+QPWZYQ
NLTE6tR3M3Yd3OoZ7sQ84UyG3rnJgZ0czZs5c8eaUEygZVycaNBR2LSj3mluCrDZ
jnLT7wFSJUs40tBr3FKrOLz3YMjUHSw3I4pBAUK2G+Jz0LwzKOMKbkWlpMoMVMeR
SuU3dYLh3OCSfzdEAm7RwQzF5M6rjo8lsWxwn4P4ToiR95CZzhrP8qtxHhiuP894
rcyL9uFMUw1U3hfzrDj4WmYoy2v2xpNcKcsghq4I5Y8CyT1RSwc2kV7FSLWBsagg
x9q+FcuEhDzEU7U9oiIKfhdf8f46uK76WFCRJDrZnkeIQJCf7u8kXE6W52qjYi35
uxcZoe5dgShEEQy747NpxTsMoRvbA826CvFWgMIATdVrtD3MVQwKl5P9+zVHMi7x
bHFKlGyq+d2HgcN29DTKzyzjv4QZ4sOrMAQkfrZzvK2QBSVAMvx9EQ+/Od989TnB
EL+bdDPfUTskKBoJ0ymRvfn6k166rT1eBWO7X6WdHpfsgL4QBuZGxeQQ9AbXZW1N
doe4y4ZYwPoZic6dI+EkoTGD+rXraITMRlawlVsey8pF8+lAOMA8rLG4a31xN50I
nZBmgn4QcX5yFDOd1gCN5rzjHtNLGzk4eSC48MZF+wszlEjt4QPN7860vZnFaXcs
1vZptmlM32CQCIHhqZwF4z4PfZn9HzgGKJTZilf+5H6qWBMBYJlSxsy8z81a1PGb
8T8Izp2x/ELBRpHsHROWBG86qfloB+dEOssjCQ6wpVIXFzR7MA8UG8gVH9iORB5M
aEcaXqwPCAkK9QCTjptBX7KDx0kWrOyE3X+IR4KHzrhkumquRvaCRvWjxRMgPe+h
SV/37u+yvYjRQQoHAevt3aGjX1sCxy2BgDvtudhkPS2++0tjtAbnY3P5n+nZo+9C
EWK09rUme4NOGXkg135OCHApuhQraB+Nx7JdxKX4N5uIFMK33el/LH0kAOH4Pcrm
R+fxePJpuSUJrMS5Tue0B8+Pir3FgmnPOfb3op8GXVGH9t2xFhvxUlpy7rY3vLba
Ls3+zzbXxu84qNME0anBaKr1DvY2nw2MqlzqVcT6w87vg4TMGnhwgQhC8UCcUkOR
6IXv+FjKRFCdL6HLAHl/ajzd6681SdmpEBW+5OawCtd8ftDXTS8VZJFc5o7i2J/d
dJhkqjIhjLJ6P0sNh5D+qqSaquD7KKTHK5BjaeVBYoLEHAPRZvox8IQn6pQzRNsN
2KsUDQ+Hhg71NZTn5F+Htmc7TF8BATXGKlBgHa0ccwPhVeVZDwejH0hzox6q4E9X
LkfpF9NCWkuTazbfSxr/mF6HJwCZfQrhjHBiFEtMGv1+vooFIi1b0p3ClqanMbwC
PmDfdCcggCLdpGUdMZ51SSZPw3angZktQiYvE/WudL8RCcO3o50i1Kdwejog+WFt
/gCKeeaixUd7T40k8GqIY/Hs+BXpegL15YvxIleduQ16ASEXUbnm4TT3a1uDsOvQ
NGoiaeFLLABA1UJSpHFYJSIs2q/Ir5ke9ItOAnQR41wTvktxyhShfwDFD2bBKy4y
aGXc5Sx2FdHOlXPBP5K+4UjhdNGIxa/J7Px7FsIZiCOjqJ4shmVLwaBdwQVNmVuR
Mq5d76WCgjHygRjKZHgiXvDoxyE3s5ZGkjekc9wmxCoNRcvihZqWl9n19CRER+vK
QsEMgZVlkJmyi9y24HiBP+64mKKRuaaAloIhhoIjJk4YP69uvbVFJXPh49kS3rfV
hgu+SK8vMWC469dhjLHw7hSA4fWGGyLoY+oHvkvF0QNH3KSDODlOw9a/w8tBPdor
LFtdkV+CS7QlpXuQsPtOl0CiGu+2EQVjCAtchD84zDmXsTvcvkq3E+NY0J0uZ4qk
dXePJGLGCqQ4Ysxx9hvxu4sDvvp/VAYuVYoPw36SyUaew9AYApXD8cnMSP2KpYbV
dcUI60O88O/PMaeORF3KT1gpaI99JbSHICa7zt6dvX+Ms2WP2hwLz7rVZlFtYBe1
0/8WRotZ5XKchKZCDAbras0jeRPM0iuMgSIMAJu8cOmBc/ssgUAuMDL4N9iBLAsb
Qr87Vb9bWZmfZfJfbHXIf2+IW9aKyY3ccewsgxhV/PqZCVuz9ClyUf34dCrzDdSt
tujprC17aOwDJYD2dGIyANt/gSbgOQxoAC2AbNIltHHn4jR4XknC9oNp9r696mog
UsHa9gPhgUynEudv2oSrepqH8/eW+CF6dcg3dLCnF4Tp6sNsUp+qsa6d17q1P8+i
D7mGMS8edSQEHboSdMdQd4mnPzwfIVpfN0HpjWtReI6/v7oC/PqNl4uIyugw97gw
zenFdarvUO2YRCiyNedlpxk4mw6oaIAW5zz5KwGK9q3NLg53vKeAraKgoD7/cvcf
WGEo6tmduPxJxIcFK6GUNsrimYpkrDMLOa16tu39x0/Xl4CF9KsBCMtLEaC3Fssz
Wjx3ihATZAwliaSYeKd9qAg7RTE7GGlRVt2eGdTUJ50FnECnAgsArNkPUoSZBkhh
eRGTjP4zlwoQp9sxaUkewpQYhouZ5FJI9gNfmwI4CXvy8QoridGp21qd9jErBBgt
vEf97GpB3iBBH8fqGalYCC9Zw+7k3nX6ovyO321Nh9L3vfRoMdJqWhM2aDb8FgL+
UCoz46pp5v38lQNQzeGKDkN87NAtEPLGhx7A3KLcAyTI8nvmvhSZw22IRfuRr4r6
Pgr7Nf4t9nClryKrl5bcQM0RQ5swGrX+11NwuA0X1OoeTzembdUY49ySS5oNoaDo
WGWBut3NV8ote1Twg2+L5lHLqSXMgUiJAc/Wk0gBcyLZQihwEqujcR5o5/6inyjs
87rnfFONh3PQAJ5i/OVhXDuRMNCEXIk7doW60EaESJghXNk6lVdYsTrAhl3bTyNc
V4HOjHr553angTC2S6ls3O4pYYtwQIY72n+NE/lusmOPOybrdHfwJZHQwUzPfh2+
A5h0h5DKP04qHV5hfx96gF5T1F7feQ18r+C7mCU/6oV8u0mVsBKx39WJ1/cpYxM3
Qp+n4sQmfP7Z+pYt+7I89AyKcROCCqhL8jOhVgOVkskqj1+P11Q4MdoNX+b57EqR
84h6BBjDSfDMrmz0dBTDXwccZSFMS2xeHczz59jvx1bQ4y/Xb+D6iTSub/2iZ6Uo
+lJZBGlnfwHNghx/RocdBakN2cA4yQwYPrNFFDpf47P87vuDyJNAdxlLsf4IXDP/
KASgxXQKNxoTXtnh1gVYNh+EZaxCCc3u3C9ih3cF1RAuK9c6hCxx3YvfGXxx+0ed
zfTpEoupwa0T0vl6U2HYSrFyW+aJwFeb/qx4awoqpiuywqJulHQLT4KyFoassLsO
PtE1GRrtbdbe4U4I/zToLgCfi9oSmuhPBkHO/Vu3m7AJavSnnqEvHqeRp8Apj2AT
S0O2v1IRU3ozpheB4BjARnM0OVtoxWSKLUVRsZFjRdMZnXpHZkdjtRulgwF5QVzG
F11YqRU753WzMaxXxiuzUkW8d8+TeRiUtbfGPpc4XCB7n/b+NK08DG3S1VWT7et/
kd+Cuyeaai5rSZr+0vZh+iM2b7WaaugB7ZR7ZXs3QADSRBvrizTlc5pdoHxly/Oz
Lg5yIaoUeGqM5iUd8ZOt7YQRf/EfYLEDI1yBuEphiQCzmvAhyHpO/ex2l6+yh9RR
J+4OeEJK0PuW3mY70mY5WB5E/PWbn7TqaJNQ4aPH4rP3K5e3R+LJ+GgB7pVyTRJG
jD/73XZaNSh0jO+HMPYFUlxQL89tWCrBnZGc3fcQcGb9KfgoPW70SqNOXDeqgYVX
shXSkns+Oh0UCFnKWeuKbRkrtu9uZBnJXTPyfI+I1sESQxA/pnnGT3xiKqOnYIRZ
/T0CF2pZoZpAKRVqx7DPD3jFZK2HxhvzQKRl1jm77KuUaZQi7+xdI9u3v6AenPXG
V09kAKah7gR+OAw9Dobzf0Yb9qTcz/KkOlDWTPT1MQbLA/TRQY8cQ8jWyXI8ulKc
8Xqhitt+i0hpDA/XSVQ9/HN5vF+UAtk+4jA8nYDatwY/9uM9WHK01+qoENj9bi1D
hwYdlyYvz1CSgBhjc+HYaXFZaKvOtsmociHB3h4HFtv/l7DCrvI3z/yi73/K14Ng
YP87pw6lwF9Yf2drzL/RgD7QtXVvNRKdd9JY0z1Qpv6+tJB2zBfGenXS1kxVdHfM
ItwBFv9j9j84Oh04pkHxoq5E5CRPzzBjNQvnTKnjGLY2ShgidiAcawTZzgAbX+gk
zEaJtgUg4Ur/6sTN1ZSLVDyG7F4jJ8I72DxaxgCO5KnPJC5lRIIXnPCD+uFssWog
Z+OdvE64m6HAatR1xG1HQR6VgUjEebYxH2JSxl3snVjl5tKYtWhAW5RMKyYDAygm
/kMrJwPQfkK8ip7uf5ZRzg8ntCdUo1zF9YI3ECKxe5O0zZF0CcF3C8/DfpRv6lwa
bPwfLgpqqMYFnHXxnIMS30jKsoXeN3K3ZPFjGlT5SAd38Z1y6he0AEIVDS2ivsZC
1HZcA60J4YiNLe8VDcWH1i6mOAgj/kj5BQ5jw4lpcVN9M9ZybzO8dqfDKsvMxSOy
iqkXOghJCQWLMg9BGML4qIxlP6ycKtOpe1Qsl+H9vEkl21vNUcLodMkOIGC0wh//
Glvm7uxMjGkryOjTff0a9QY85PMsEUdn1qf7jKURmINdS8f4UJr9ny51/D59/ugl
xHeOWAzqb+Wrt62dkMZlIRZ4Pzh5gch0WmmTV54DHk1WwSOJcQepg0zj3AcJrm9o
wdYDWp9C91XKxHLNHSPaXaQAC7kMbCPYJU8KoO0zPth+eC1SDru0p3aKVAgBoJGa
7tNRXFRpVSTSQOG+qwn5gad0w1fqglSzjciymwn881bPSLjsRauHYeD68m6yzfQ3
KvA+qiC1vt0JVuBW/PnlUunBdLDqOm9GCw+SzEfRIwTHUT7cOf/6noOg8MIGy5Ic
Cfy+BAi13Lsz0DAjvb7JFGx0j72eNVQ0Xnyh7qlfnfBcWCDvLLGdOe9SIVXMWIa/
BPdpdGEWxkwmEgkwRE+aVpM+4FWzErhj2dDA3Ai4NE3O5We6EiGA/Whrq6wFLjVk
ABy38VAXkPabMaj8HzF6EJePZmz6U5TUzZpDL3fw+oz0sTJjOuV+o2Geb08Zelge
HvDTmuqFpX9rNYAz7qXt3I2fdsMuExw6qzknT24fyr7U/ZsCS6v7/mGQWodTbSxn
h8yJlerTr/G8mIugoe0fIUZX+FKOpKUnw8MmuoCFdg2Lh7tsShWmSDRy4y8uTWMe
PkeLNOrYl03ZGpJAv33ku44DlBZlRVWZjRp8fGx+qXjGUqnm+ZXsDPtfuCV1cm01
oNbsW7OwuiQxdhFgeW5a02brX9zD9y52S06cEF1aYO7NV3o7FummE3Kf2GC48N51
801Z1/Iz+SPym2DEA0VK4wFxCdrcuiFoux2pxJ4ZAlTrT4EZ9bcqnTDhoHT+xSU1
cbeUWOxFlqolRxhNrZo/z8Zlnt4nYaQbYLYUJHeMQV0fHmYnfVxRKGGLJJqVquoR
UtmI3ZVh6vIJgwpa9s3B3f2SAJJBhhv4oELBh90otaXyo1aSr6uTLLEBvQrx+Bdk
1vrOILcRAntjC7l/l3QPk0WVDjSlWqY1w1eCRZSqd6bnp6Z0GJdfuugugS/W8L/2
1AXJ0JBaSF/2bqyN46AatixD5+E6WaXILy9hHyKvbxlHgDfDbxEX2K93oQ+9a3Xr
X8B/HWmeuFCTX8kjVfQA6mNax+tDF2qs8wfNqGU8pf9jKhoXzHEvMm37oMY5VnBS
JQCikTclHYMdLOa/der6HKt0KBX8mPKhDIFInEighphKYJw3T3zcgoRDP3b1syMu
KMnDmnVezp+HK/Ear/xCEP6Ju8n+K4dLKEYNbZrJ1lxRgvhmyF8B/Eg5hr5OjW6l
9Dt2kphVHTfH0iq1IKNknAodyFCxtL5Vm04tcDATAnmn6UrYe/iVt5ZRIWbv9hQn
KDZLZmgx0cugqSnS0LtjdHZ5UNYnhoILVcHQlaEbI1sOGgjoK8E4MbepdDDvzbAE
yKsJu8m9b2+N7DhReWX/dPJ8WEhjLjeM3p886vpUVJeaXo90VogFJcj5gMlBwC2a
6QYTNwc3iEFqHQp5CPoffHZC4Lr9efg8t0F/dFCGeRhw3jtKKenVT9O1ieEoHyZ2
3IyLuSqxYIxdu1v9g14FW90Za7P6E74NXtIANFyFFtaXfR/X4kDicEwRnH79+8GF
szFXiYt08diYLtTWsWICU0h69X7VrxcgriJF8MsCpyZBPpYaxSQzaP3/hiwD0DoB
F4VNzhqAKGig65oOeBmefkcrjK+ARB4RkLmFh/tzCAjOpqwGqpm2s2zVfTHCyeqY
o3R0T2lmi/F4cS4Xtr3+GJ8eOjhFewzPgSN9usjGxMSIn1IeNkT+Ek4dwWEDtczt
9Q5/tO0Y6LuHrPhfzFzS2de8EjPSVWXnEb6F6nOGtJn5iZj5GQ/X830/ouAxrF4f
Swa5hlLe595S40XObZ3zW+ENeMl62G/8d1ZNREicSzcUqrZIO4kiKolnHgKQbpSF
BGloMH2at/vvc06OAihGfviH7EX//B20FX6F0a+AIPpurMqKmetmHM3GMiY9ExQB
x0aH/RCC2+1lh4n1cz0l3+RqdnfwggxqioShFe8lbsC6QsrZiI9JuAw/ffaUqnzh
PwT4g/Fml7s8l4Ze0BmDklDMdwH2PErZexssnvYwPrG7ArYRab5rCdwxVIewz0ng
re5f2S25hiu8OI34CA3+7+MWziQ8L9a0SRrgZAEu71Y/nCNjP1ssoNXyJCvcKu3W
11p5OHDuA3JDRAJ2edZwOqIxv5QUncgDEvphMOnAfrVmJIRP7bLE5Xo2fxzvDf7c
nlsy8aF3PukwMUBgBQ/dEZ6hcuyZXwRKpRF74ZSBDQAKV2pyibvsRoIhAtFw6OFn
yM+uizltBaKZ6/rtlrT+qvm6PfUdhoJ0ITKqh91M1eaTXCfnQeQy73UWdoNtoXnf
l7ZScv+faSXe9gYx1EVdBPUcdO4bOMzeGtRnfFXq+SdCcOx10YXvMMfYl/0Oery5
kfK2k11tXzuGN2tXdIDc1YhdHpK0mYQ80kbMgFB6hzS405Zdp9Tzn9KgprUGkAwn
sb6RWUceWrrhy0QrSerVp3/UATQhgusYpweTcGlIKqJKledubgd0eOVENl+6pUfP
bxwLEkcNYjpQKsytiBoNPzwYlRrHO9uRB9rDf8mDGwDzhUaHxKOORdrga3BD+Wg5
6R/mUeMXIOc2JIMNwKtpv8/vq6zqeLdAWSwFFfr+JVLlWjbW3hNJCD0VcPJlLlSf
a5HCsSwRZo0kbzh8a6DlNoomktZ6kEnihp9Mni03n1kovk6xT1B0PrpH39uFOwRX
M29gGsGLcu6fXzaElT/HYalbxGaTticAbTcYzOThfo9DByE8kU6hRpQ/xChDDXRx
ImvinrYVYRO0BH1Cir03fNiq6i+nAqI0Apa9GkPycZkp9h3vcQqChDD2dsF2zcPd
xmKz/UObG+rHkng4onS5mVXN9HK3ddSIM69A3m75bFeNC0UCpGOLrt1NHKGmIqHX
2CUtfUwH40zx1xx+/Cd0hcG+XU5yaPg8jUDwyF6jT2k2o8XhSe5mRTWu9292cMIj
QmY/aLaO78VpzOQPZ9O/g8hC7UQJtv5sgp/ujf37CoPaW4KIDeBTlPe9mYwUtAj9
0WAgvpXGgZ0jedieOOsoiD1NE+q+DY7Q0zCC7V6m62R8S7mb5IiLqA8Rog8pQnmv
5EIyC3VOmIKcG9I6zSF5+Itvs73uW4ob61/nQcX60x2PzmvqMfm4UhDp7nc1etGp
IYQw6gRISnhfJ1jRM+r6/7QfiwPNVVNzKcvCAsoviLuJFcTxdHfw3ru6a+4uhD0N
wYn65dXWxwA/9PW/m2fhA/+/dVJWRAd/P9VuH9Cgyhjo2YqUwVu1aaywO7NFNfSY
/juzyIkr5CEaGXamgW6Vr54i/3aqQuP0zYN5ANJZr68c7x7QiKFUDV16fI22dJsz
E3O+UqTM++ltIMi63kT1dhLKkmG93pfgNZXnl7cC9r4hbPR2ECjW/WTYMpQRjB+H
KkgeleKzpOh7r/EEIsRxuj/+/0DNPH4iPq3R2VSt6LOWJbJON6QWOshSpTavu/8z
bTBqCUujZv4VWI2cv5biKOZNb2fMHZi24/mXxDYHRwesrV6vFGAfkeL4YcoTeuGU
zr89OCla0E2K8OnEBn/IKAiEUIJJZpJeKXpqEHh/AoxBR0VmSYWo8KiYf8QiZ2hk
o7SqQTABu6CjXvL57LL6OV0Cn5mqNBSfqqB0wAd9o3diSSZnpe6e8QTvMOTswaQq
J2ysJtClETlTm0kcWxHfrK9lKxjbcXVIxym3fdNSBAm1uoxI2fcULeIB/Wx3I3P5
DNybGBiidTVOiqEFKobdm6DaYc2ZbssF2fh3tRBCCDZikvPk9cB/ynEVOM4vhezC
aSQGAExk84iGoEbZvskZQ0IT1Un0lNaskPKeMDEkxr6tq5V3MghYgINBSbpf4I3A
+YRnxFC6VFrWSiPo9XCQOpSLdzE32C8Kt+17Y3sOIolr1j9fVaxX9TUMWzMB9EUq
o/czGUeOmBX7N5FV5AqiikJbof3oEef6xa0SuZIzyVO/MkCn5naeY3tONgtMe0JC
4a7/WmrkkDrZ3tfTMfp+omtmuJKRr/hn7ExgwCFJ3WHDBPGVC+gg46fRJbfLTRs3
uYmRq580Fk4Z2eLoYqS/cg==
`protect END_PROTECTED
