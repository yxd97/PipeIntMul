`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
47xpuIsY/63/avFCUPaVZITqBLVvEOa4VaejkYh2TZ4VMSUIT14t6/sEGLif6gI1
UfQrVT4MPjJqYoyZJ34JhQauXGxduQFobq+Fx8/ukn/k8OPin2SBASiXTmX5OAxP
8i7f9BZkyZgtU7cPw7E+ki1Bt7owRjoUwlGBxpiDt1kOMIeLnYLAfA2SjbQG4MYa
/yND5FlAdIuNGB/UmqXSpz/IU76NLcPRLfQDlTH/cb5rChEvLW1YNrwJ8ppzFy37
TXijEdK9ZjQrYnLy/7TB7eOK/eYFmqHkmB5CgEijh62A83MIbBS9fRZTAypKDWwU
58cjNyeVQcvM9TbIf5sthiL46gA6in6MxIzEAXxGNIdfelvLdWG/ozmvfplC4d4x
9PW6gvpEezeBUturrGWbdBkePkpn5AWWk9hcx2LbdfVb3aVUVhvaSOMqSxavi9hd
/agjDmpBJzu7wbTCRE6Oina8Swi4PCnz7AzXVAfiK2wdsKCEqJHO0QDrQPacPH/X
8nlS7PDxvtIgE4ncypWh37TSqLceqwt8znixbsam+Apu0L7sCbdrYbKUeai0f2j2
zK8Jm5lz0wNB1v+JO9AnFSb39nMxOXwtq7j/koz3Eb/ftFQEl/YO3UKyt/JeK1LH
`protect END_PROTECTED
