`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xuo3b9a4JdBRHNSg1U6F6MOyiIaduufxCeXOScQ4xxadJjnli5QmIIsHSXTMx2wE
M8iP3g92k4VFtHJ+99RCGahBbbOfwM0W4pfHkk4whCHbR+2fH0j8q4qvN/M1fXz8
uTF0H4/duomu4Mil5A/m/x6G2083nVRwE6fp9UVqMe1mFNGzQJZwWRZYbPsTqFHj
45SHWZo4CTF3MEdLzkM2yz6kYIHb5adZGjyTqEodAqBhTn8/IXRwqoGfAHRyHDNu
gIPfo3YELetL9Hw9EzNO5w==
`protect END_PROTECTED
