`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8Hec08+I2u3eBQQ4kyhKsFRt0xbH3jFTA8OPFRiiqJC7oOAN8eltdsfRl6dBNx6
1TWwTfA7rWdYqSu1vXkZWyqUKzszCK414p+QEiOg1boZC5KcwclCq/VuF/p1aab7
JxLy+09NSQSexai73lpKbBseKYkx6jUv6WvDwixhV460A/0qmRKK8xiy1YGSoBv4
Y8YhEYcF73zgz6ttWx/IuStlW554ReMwbtslDcXxeVVIeh2l774ngCjc89JJMJ4r
/rIHGcSXbSAhxar+bHo8G+htMYh6j2EE7S/u+yvuTZOOEqlBwyVBDt4Cy2NI61Hz
3MMTzjzye912xKG2VNy9FF8rqbVjMn2i2+YM4rqzrJ2KvODJ5s9maCc9Ahgy2rLp
thZqD6+uUy63CFD3yNvBIwoz55TuLq81+8I2477iiiKLNAI11nT6QCWpQNRIL9sF
9kBF0UuOnAoRmYYWaRq65afoFqAIOdx5AFYoPY3EL1EEBwlbRXQPPhsZKMT3hOQ+
LXKLtgmlwbwZKWp4hSgPgabnEpsBfU0D55w5axD2LqWatTmfmDSoyXg0jYyMIvis
cLYPWf9PMiAEPBCsDNIngHB91ZE655XvozOprlTXHK4lwhVrFJjHfzDVTOush5m5
P/KW6VhTYTcs0EeHprveY58ha5lOs3NE99mnHOiAGI4=
`protect END_PROTECTED
