library verilog;
use verilog.vl_types.all;
entity MULT_GEN_V7_0 is
    generic(
        BRAM_ADDR_WIDTH : integer := 8;
        C_A_TYPE        : integer := 0;
        C_A_WIDTH       : integer := 16;
        C_BAAT          : integer := 2;
        C_B_CONSTANT    : integer := 0;
        C_B_TYPE        : integer := 0;
        C_B_VALUE       : string  := "0000000000000001";
        C_B_WIDTH       : integer := 16;
        C_ENABLE_RLOCS  : integer := 1;
        C_HAS_ACLR      : integer := 0;
        C_HAS_A_SIGNED  : integer := 0;
        C_HAS_B         : integer := 1;
        C_HAS_CE        : integer := 0;
        C_HAS_LOADB     : integer := 0;
        C_HAS_LOAD_DONE : integer := 0;
        C_HAS_ND        : integer := 0;
        C_HAS_O         : integer := 0;
        C_HAS_Q         : integer := 1;
        C_HAS_RDY       : integer := 0;
        C_HAS_RFD       : integer := 0;
        C_HAS_SCLR      : integer := 0;
        C_HAS_SWAPB     : integer := 0;
        C_MEM_INIT_PREFIX: string  := "mem";
        C_MEM_TYPE      : integer := 0;
        C_MULT_TYPE     : integer := 0;
        C_OUTPUT_HOLD   : integer := 0;
        C_OUT_WIDTH     : integer := 16;
        C_PIPELINE      : integer := 0;
        C_REG_A_B_INPUTS: integer := 1;
        C_SQM_TYPE      : integer := 0;
        C_STACK_ADDERS  : integer := 0;
        C_STANDALONE    : integer := 0;
        C_SYNC_ENABLE   : integer := 0;
        C_USE_LUTS      : integer := 1;
        C_V2_SPEED      : integer := 1;
        non_seq_cawidth : vl_notype;
        non_seq_cbaat   : vl_notype;
        ser_seq_cawidth : vl_notype;
        non_seq_cbwidth : vl_notype;
        non_seq_out_width: vl_notype;
        INT_C_SYNC_ENABLE: vl_notype;
        NEW_TYPE        : vl_notype
    );
    port(
        A               : in     vl_logic_vector;
        B               : in     vl_logic_vector;
        CLK             : in     vl_logic;
        A_SIGNED        : in     vl_logic;
        CE              : in     vl_logic;
        ACLR            : in     vl_logic;
        SCLR            : in     vl_logic;
        LOADB           : in     vl_logic;
        LOAD_DONE       : out    vl_logic;
        SWAPB           : in     vl_logic;
        RFD             : out    vl_logic;
        ND              : in     vl_logic;
        RDY             : out    vl_logic;
        O               : out    vl_logic_vector;
        Q               : out    vl_logic_vector
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of BRAM_ADDR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_A_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_A_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_BAAT : constant is 1;
    attribute mti_svvh_generic_type of C_B_CONSTANT : constant is 1;
    attribute mti_svvh_generic_type of C_B_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_B_VALUE : constant is 1;
    attribute mti_svvh_generic_type of C_B_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ENABLE_RLOCS : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ACLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_A_SIGNED : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_B : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_CE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_LOADB : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_LOAD_DONE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ND : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_O : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_Q : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RDY : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RFD : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SCLR : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SWAPB : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_INIT_PREFIX : constant is 1;
    attribute mti_svvh_generic_type of C_MEM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_MULT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_OUTPUT_HOLD : constant is 1;
    attribute mti_svvh_generic_type of C_OUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_PIPELINE : constant is 1;
    attribute mti_svvh_generic_type of C_REG_A_B_INPUTS : constant is 1;
    attribute mti_svvh_generic_type of C_SQM_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_STACK_ADDERS : constant is 1;
    attribute mti_svvh_generic_type of C_STANDALONE : constant is 1;
    attribute mti_svvh_generic_type of C_SYNC_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of C_USE_LUTS : constant is 1;
    attribute mti_svvh_generic_type of C_V2_SPEED : constant is 1;
    attribute mti_svvh_generic_type of non_seq_cawidth : constant is 3;
    attribute mti_svvh_generic_type of non_seq_cbaat : constant is 3;
    attribute mti_svvh_generic_type of ser_seq_cawidth : constant is 3;
    attribute mti_svvh_generic_type of non_seq_cbwidth : constant is 3;
    attribute mti_svvh_generic_type of non_seq_out_width : constant is 3;
    attribute mti_svvh_generic_type of INT_C_SYNC_ENABLE : constant is 3;
    attribute mti_svvh_generic_type of NEW_TYPE : constant is 3;
end MULT_GEN_V7_0;
