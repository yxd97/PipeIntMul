`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICvX/3qYmqYzdGs/EjsEEi9RS7pVYVs+OjPwOdAIh9qwlWSLcw/eNNz46FNdU0xi
GiNFSx/A9+lyAjxDNhasyWRihDdZHIn2WshOB/r6PmZp3mfGvnXCD1pU72y0nLB0
8Da4vQIrJz5ASQtHtflTCtHBqM4vvhqcLogtuGGik0MIs7XwhhXLpUn6jQE4a1ya
sXQX48rVnXLONJu8Ya4yyx9t98c5rkM46PJkHc2aWcXZpl4CYzIvT8UYk2hGmMPY
lugs1uLKCBNu+GT8hwAdU+kdacAP49Mg5SiBk5nC15OitKus7G3sySEt6lvNQe0E
d/fPWUT54Dus+fcQ7c6M+9hzJ4wzTK24kQQy/b5ZZHFdxfj37TwGhg3ML2gpgdBu
n+KRpmcDW/i+u3xDa77IgcTGjq1Z4FafnLZWlpIUWrfbVLQHwZIgNBnRVcXzF07t
piFuCOsVmm8HmY4MecTfhygx6cwhegEgu6W2OgELBWI=
`protect END_PROTECTED
