`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FhERCNZ2288BDtdneAxFkVj6Y9/VmkFbnkDv0TS5Vtfw7yNH1yc2GSc9cG2dI9D6
oag5+ymJmr7IDc+SpfLTR4VHPPhs5r56oGVB57wr+ch9xosr94+XbxPNB2ID5+BG
6DlWG19gYRplGY+JJWRPXfbPh3EGe9XQZDlxZBT31/5VjAnhbIibLCaC9mVHSGbw
VmMSA1cZfR9v0clpdYyRm/CXpYd1dzqRM3TR+M14b8uJqvB9Q6BIXeJo+wpYR9vJ
CBaIOqtswmWWUWbGhGdFldjZ3N7iW1EG1ctnSABvOlAAxk055LXKhe3vQhQSyRxQ
UwPTbYUAXymGGnfcS1gvRRw1IhY2nOKB1ADNVl7sHRU+fmmCWA5kSjiUvO4KoNSX
FwsYIVjbiMzqlDobBW70yNcQVcGCMMNcszvxqu11jJK4CpBYSyj460RuWMJ9HKf9
IMMx9LWFw4W5sxy50cb2ButwZLqepsRY2B2YCj6mtyxT5Xp5nGCkaehvSxhyf4x7
gFTAs5//CopvRSipW6z2y8I9GPhTueAkMLia5vjaZVO5XrLWwmYZxCKKwi2e0gdF
ONOaw+tIzkyMbCj3c5jKtroRldmUUxsxhu/4Q/rWGPQ=
`protect END_PROTECTED
