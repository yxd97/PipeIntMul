`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xrRWunIu0rYym7Le0/j5kpYlHHwSE1wx+C8fkX9UTmLbGx79A0irMFz5BPD5B6+K
Tqa50YXPieWd1+stsqtimBwK3jqu7S6du1X5do/tW+Pl/OAofRhy67F4Q0zvV18P
HVNWElcuyTuoFwQ2G/+ygcDOVLfWECHp91ojtz5cKHcCfqiwr7nOulPXIVGIn9Pz
BG75pQIyWzAE49jPj+X/TK2/CsdJQoCUmrXcDLBrCpBrd7A/YpxhM5RS+48rDkyW
cqpqOuEQPleMjUFzH5Kf0qrsuwrafJJO2A7R36Px+krlJhveldKWU7z7jbdNVDJc
Be6q/KoRhyxtaFdqxl1y1J7qeQy19W82Eu3dKXoKZRcodTVkYzCHssy4di2VZ+Yp
ASAGdSEcPKUsdlACacBJVKHgW98vDEDhlxk4cFeicJCS3iO1Fi9x6XNEEcrQieyu
6OIBJxM18lHc7vSGPW4TtNTRxCcd+FpTrhO2OZoqA9oX/yCdxLPTr/kee1Ow0xY9
rTTzHJoXXDFbWoh5lFV/8OeGJc3oISRFyAnVrmveXEGIMxiaGBipQgXFu4Qa6zbQ
1RyfayBUycjy/h+eNj6lowy6D2taog/nRDnfH3bvp8WkivMB8p1UuUdWCRzYyl68
no20uLVLLg4XVRB+flI+W9lTysLbrj2BmRIpkboMDgyYvNd5T2m1F7acl8wO6JbD
+TlYhzwZSVMvWY6OvuvtcoaBbXFHJ52PcOUAnw5chVs=
`protect END_PROTECTED
