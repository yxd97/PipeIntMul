`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LX+V47IeWmZKEqwdOVhwgybFguVJmnNJoz6eRzf89qqtX6dDCyFM0T64UOV92I/K
YSLkyOSzDQA/stp8NgBd9ozNBKLH5HcHhKLSVfZaaTjK2V5ytqp9I/iLhH+BOZqC
sz1+XFQEG+xhV2Ej1ULGlbIZ1qHISe20RG8+G6ND8Y6DUXhjLCoXGBfKiGcDkPPv
rSrZZ55GCbBqNIQ6lvp2sD9Bng6fGA9Frog1FE5rDmKuZgtw6052Dk5OEHrN6RKr
OxhYhg1w7fYhP3dsey7t4v+9OXVCZp4Gz1pfqfXNerGmi807d/G19k5qtJ5YBbAt
tkxbIjHTiHTBv5N1ulRfNA2PqI65sp6FLSHsAZfP4z/eTG0PdATRVNdr4NvFV4XA
wed/lk/IyleEkUDfxp8YWqdUSs+tmJtpzK7kq+tOT7Uu5JJCFksupRjLmtvgxIik
90Wt1VhOqbsUJaNqrvUZmFLTLYilHtoyJ/4wJGha/5l/UdvGQ57Y2g3YIcRjxOwV
0v6i7j/Go0jURI0tPZWQlHeG0YiytnJM6NNtEZ3y7kX4OsfJV/NypDdekKx/nVmK
`protect END_PROTECTED
