`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9SJDv46hYTXbIcIQ3D1//+YC74nw9PTiW0SYJa4A0vN3brnex2xgHHfg7AuwsLde
GqdvqjM2TMEs3WTwMcURb2n6d4Hujju8uK1pKmQkhtqTLnSqM3vVQj3G5mrAMEK6
TiFCwz6Kq87jUm/ooUro2fnf7uSzBDi93DPq9tAeW76W7Rk+Muz4bGYltBDCCt/p
JKQuaKMCzQn/8MEq9v92wCMuD9FYqkH2FjO0+i7GAegkbK5jIZdUTZXipMCTTcdS
MjTpmToLSdscrnLrOrbmYpu6V1JVQhMhGqceolissrjD+L9AhwG78E6wpK0XPwNV
9CPbUZUzUkfpt/N6PBdUYvU0j4jZRTgJUPhiVbiWS8tJqoAOmOuEXGCY99k2soMs
vtmC1YcT3t3w3VZ0YQqWImMPhC7FnHkctW/9jXUS8BIoNHuCVsqcmIbRV/haUnq6
5TMsOL017T3FAHlFuYjdpWM60ih4qomf4O5SxBMtJzqY7EZpBs82clWL2uVfcqJT
4RLSlG8XrmAfBH1oC/isE54gg0b2bc1/dfWwa6R1Ld/QS41/WwknxptFZWlCRoc2
XKFSvK0jPi6o9JVt9bfYkw4QbGsep/+XoAkORs/Yun0ZWVzmib/obLX3AQHR+mth
3SjdghV1N8Ja+X7IK8EDA7xc2uYgt1WIrDp0RPSN4SFeHWBtUcIlES/jJBYU75uO
rrgDJn18r4AYepgcxCrgEF+NAAgtdRha0UCh1rqyJ6hPwW9Jyekh7HFRb29O3h+O
24WbSmBBF3dp1TcE9m5P3OpyF9QguEIyDjq3VaWyqIxojWp3dBp6e7cK4f4xI9CT
91Xrj2ZnQcZZxV1N+4csUVhzg0smF3uPLoOfwKeONQtGZaBtVtUGnu3aoTvrDxfV
hWBBG0M/ouO9cwFOyNiHLdVUso1zDURQqa5Bjh+DKfgBrMc7EVWd1UP0JwKfDA8n
`protect END_PROTECTED
