`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p9mrwigxfyGI2nljDsoAjrwqQo7ONEwxdDAOgoaC4LAk2tBq+9ltJQybB+Sa8zQW
Pm3BMcjiBF5zea3IyV38bF6HZ2ePq5VCNAyXXIfy5UJb8/NraSkqTGJCGP4LsEwc
9UdKxZ0T7utdNLlujBfxsLzz3Qqp0CbuDTe3BoJxSvZAgqWNYsRmiAjJRnDon5Ng
l4Ptbl4xkEV+NFTS6VeeJBS4TFaGYuIr+8bnm7YAG/Yh/VXHv49GBR5mMwtM5U5N
cAOQYjYwuSpR2gHS/iLPowCvzGfd+Wtjo/o5eWwZUk8oe5HU0jpuYm64TxqPOnpO
+S/OO2ng+8f8iQgTGFUYMbIptFgnmoPF5YcPR7hNc8a/vo/v1ZMof4+fr1956k9y
YVc28pVPdkKds1qA7IiVCZU3XZJ9fqz6oMlrHfN9+rabReyY+Kb7PvwTCeMKrd7e
zl4IUJr4AMf7c0M0zIeMI8A0E8Y0+w3ci4P/KxmzAJ9hqp4GAZyRnbw0S27fE6yr
DHMl44c5tvIr6c+AR8QT2MLs2AihJkbaiBbXDBEU7fEdPTFlwahDD4PW0qv3otm9
4BwqqAgOUEkiPTEg4pbrK8ss5spHvOeu9qU2TGLNFspY7IXer15r0Q3IfMdlA7ve
Wbt/2JizBNO1VLuVbb26dV0wfFcRYFaAAH/1FFjgM6/2UfyJQBHDfWYHedvHFFU9
Q3w7QLu19NL5Hxc6AibdZCv6ECqno2fgX/26wD6p61+6KvY85awF+yBAPDDUvMoy
XZmTYbR7DmWeyqKjOy+nocuNTPcOWfxQH4eYlHPFYpEjjYdKJdL34RWm9JG9Az/0
FDPGoapapK/XKmNeKmdVOfLItJPeJE67eQscMeEXf2tJEUQ8aO1bnfim2XX97Mey
A29IExLEZFM76ibqX7hYveWVLbpXbfU5+Cma0X+vm+D03T+2TnZGPbgdeZlL/Ce/
fjWtiDipE2Jvyzu6wc2+YJnS51j3sg03OXtk8K7FH2cNz7UbFvGrUH3j9g9p93nQ
BT1G8S0gvqXtmTHRaVKNdDY2W6CC49v0dHRQCJJccFmJrdYuL3jcJHk2yDaCLW1r
FsqBk7MTzkZliSv0bzihnXGio+qAVbBY0jbia7AzwctBP7DKftj0vRYro/NIZDP6
+5XnI5EMlwK2CceGNvO7jW8R4WpJizxyzdr2xr34WkuOx9rPSoGneAANOgUsYlTo
uHcJRxkRom468/NjaGExJTMjp9ezMh7jNnxqd8C7hgPBwYFvFmTT8K28vdJZ2oyJ
`protect END_PROTECTED
