`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8XG+Ku/CrMsAd+t7XaX9U7o0VtT3CS76HXp+KDuDJo5qPA6UJCw9fmw4PsU0UQpf
jlcLs1T8X+lz0x/sjIMg/UHIVVnprn5AtAHNsQoQWt7VNvhTjdE6VqmH7/karv4y
Q7ov4cPyJR9ZlRjnuIWWThRNZYvjSaA2yr/jSsEl6o8GuK0EWIRlKIya6rSiyLOB
11BeU65B3ziuu0MhgNmw+zyD6NMEDpmqVTBzenzjQkD+MKoWt7SHlDVFCptJwO/g
ZN+Ux4Dak3T2IwDF5+d4/l+U+DFxk6xNeAkCoXgmpIOxNHN/R72yWX3pwEmvV9CO
cHYbLa9cOpEuhIj2Mmyl7uLHnTX6fcwXptE0HqrrhWPce2y/BzpOmSSO+ruINh+7
Q+2lKQdM5rjaXiZmWSs6gO3Grif4gWci7Uc8GVzk3IYplgbCmX7oXBm+AKLHmEri
3DvgKadn7esCCKEOzyvj4ezQjF4fpZO8W8kVAENE1ABmIx+7tRcAW2fSslkHdaPJ
8mSoBdlpw0Yq+VWlU0GuIBxnIhKf9HFc48sQsbjFTJjNoJMNlIaZlZsJ6KL5NoiK
t26BVgK6M2vABgg/7vU5T97Y43WI2+jdSIBoXurfDLdj95KdKjnsM/e1Rav60fwP
0VHw4Zi4UFgSG1V2369CMXsWgtfJ5qtldE1i5nT8OUoqpuWwXHbGCD283SyiF345
oBHMGfapdQ3yTgIjlCq+V9fKpjoI4J3iSvFQhHdlvT/busXLHPgMJcoTFiAE+BGg
mgx3910qj7pFvBHKqGcQ1GdZE7eU7678ZSDu1vV3MwvirDU2hgurCdoUQIHjSazV
9/U5JC7o8jlQtP1SQRMCWoxhbO5YeU/ZGNM2YqXjKJ8QrfBEdzHwUyGZ/tNgjMzJ
OQnZj1BprSmY6rq1gSyIuUwCnzR4xHDuhelB2v/WOqRRHay5sIJpa5TfbV9rBS4j
ggLIMgwDMAlihj6aOw4MPfp12HDc5+Es3JiO1mEebVC+kr8plo/9KiYyhE+oy3Qp
StKk0rUJVMd2bK923YpRuUKfnWcnidvCEK/61DsgDDAd338YJL4k+yWWeS/aeQQX
Hxs+ZkmyMr6emWx0RTmUaVuP2OjekaknCPpiDT1RD864D0lTjVuknKOIwrgPMdJS
VA63jPbGNa92D2N+J8E01j10uGpkcIM+HiFwZAoDRTbBr6wiA95tnEfqA9uEN/jb
bswBIx4myiYuD0sOabBupXYbzY0AJvCMG9X51aKkIpo=
`protect END_PROTECTED
