`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i0b9gVFCndqMLBviiB2ghRo0tPfi3yzithVF70KMS5jl9QIUS7anMYgep7y/1IuY
dvdntF2jgMVbF0ZCnQlD2UWTDU+AHAnEYwYxNeKY9cbKjx8t+Yb9BLYkaomYCRGj
rpOzDVNooM00fwSWecBKbHjUxmjw7htsHv/x84orVKQ+4QivibwgJTEcQ6d2VkhQ
fJNfpR7N6ZEPuH/eXYke4dqDRrumCyMCfVvLa4d/5HxakfnFt8psi3NwNlgsp1PS
WR7xty1d0BkcvNL4ZvFagnnY85rykSENLl+nzRJIUrh46a4cN4gxLkGID1sZ4iAg
9RYeQ8+QUdUImIJKQrP4jlUyydLB+8S8IZKDtC3wvaVeTxUDH3rdwkRXENEabiOi
JgSp5RXkWdW1XDY837IIbci17rX6KVaaeivg5I6JySvRa/ZivYks2cHLAwe0VHFo
Str0wkqAF07wS0qhfL1mSu3qOzXbqhze9m9KxFdYBiCCMZABydy26Hjcb0oqHSzq
ptXN1kBZRNO0oV+ma1Un4cOMtLleeTryttYWPePm6FE2Hsr9We3t8Ke3gdHgnffK
z1rfzOvo1CvrT8suIoC9B4OSEIhEEUY/zpCqTJny1y4=
`protect END_PROTECTED
