`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dw9Lu8lbmfxWb4i7vGxqJ7RGJfIiBp4GzbxH/qopExVM1RGgFhod7078qx/kpG5b
ARUoMsiKkheBb4bqpeAy9mQjPrXWJt9UPOCIMvle7WgNNqJWzbM9lefNoiiRCVF6
GU1DIiwgRZabUl/2WZZLEggKYHMjBygVtJP2lhUhR9+A/p/vVXHHlr5hdAvba3bz
kcXcfVWcMuRqkdoE3r6jsQ+vPEdx/KHSbN6c6xDhbotmqURyBVsrVaG4l6TI7etS
OYkkBQp6dyLQV4lE6L37IAHIyMNHpVYAAp7QRuQMpyPxeQVPocmkNkgOPS2b/3P7
kgSVBHoTNKa/BcFvVP8xbpPrnc0ZyiMVlIDWrHz5+9dka+3X9N4IQTV1pt988mRy
gVZZWJuBwhS0asgWqqanV9XKfg7D1ebP7ZEyk/wLEKjkexw4L9vMQaa9GRtdJzns
swiF5IL9LRCArfoCkM/UMyqR5/E/bqqKLbme5Nb8FukucqLkzKeYQPNeMxBNbQER
1pVP+nWJ7fB0ryQMqxkVpqr+pFnr9yFgxUwmbXlYbpReKRWNJfLahXPggtBsEPZl
pR2UqSnwAIqTsaIUauny9r29spjld8q5udtQvIom5kO3FcrcO8aPXhTfPop4drwP
VvM1I6b7xiE3Kg5bCmPBZKD+kZV9CU7vYsFd30Kpp8GBRYLFOah7IzOtwlnh5WTy
hW2761HrR+fFNw0y2TZcFFby1+MMWCcAqRMRxnW/HGvhVqJYpFHFcoY+ufA7DWhk
NxG4dkNEi6hfiDNws1T/TXJBSU1G36lW++4QJaGxP5BWi5VvR/0H8AzvRGi48NB5
jdp96oX37a8I9OJxykmEguPmQmJwmKRl7b0wi2Zjpsc5WxhyaExpT4bPf3CwXj+v
7strsdOp7/licWip83pCtlC/BGX0XOtE2TMcgZ+bSzK3aph5GoHON3fhnwrGJbPN
krRcvqhiJpt2Hhdyx58C7um9lT9XyEpnENxWqtXFX9JFIh+jUR/pGBxqvpfHaIpS
R2GLFLPynxxmnNjmkfLQCi2huAkgBMML22uqs6426DB9QHIRLqvn6xGxBoH+2C1a
53efggKCIqs4+A8WkAIJOW+P1WkMeCSCL6xm5RtC336u8yxWQYM7MAg3nFlLWKjh
jZZZ/FV5S7DrRUknT550SzQHTqxlYF7TvcRUqqjar7Usc++YaMfpqhtI0cDj1hB2
Z7e1LfY5cbSpexy/iHP/FSBZHxEGnkuzPaU2+XPp8RP8+1/uCL+krR51dJIzctjJ
1Lu2fuOlmkb+uXe8Eq7n75zlo4F35BRQj+uPYd6DfbOqOz4kha576T9cJmG38bxZ
X2x66wWFu8d6X0rQfrBOpkv56wFMGzAEDZ0QZc6nGQSnudUVjiQIKHCy8Dp1G2bB
uyvd4YRpZvfVQ3VVdyxuQK7aCxy65nbMZ2bbA8zAN6AZOqBvQ/IxOkAP61bmxWVD
pu34GomBwaU6WiQskpzqKkOeGgkE0N8zQR45484qDmmD/cSnjrgoYHVoSORz0gyr
Qc7qpwR5OQcPcmFI6G9Sx/oUZpAJ/8Nh5p75wXxkgpRxrT93C6yQ80fCx5Xnus7X
T9RGdetqBGJviaaCkCx7QZixxeohQj3uTAhY6Eihiqt3Nm3ghVyIVUiiqqSZbkfY
+4mtBCAfgKI99LfrHRwuTKY6lbM3CQAAbztHGZ84PmgKmxFXIoq4ydyS9uuaO/OB
meVGxW8nr9ORUmPeopJ3r1D/Nzkf5qOgKtEBNe9ARBx2XrJ+GwVsIZF3oMLGwd+r
1G9nVWhh3mw0a9shisWG79Jz4RygWryhuFxv/y+g5WF8Bw1BLL0dJz3NKkTBw/2Q
Z72j44ckKKBVkji2GL4FdMADx6lBK/XgfvFCQXYMgJQ=
`protect END_PROTECTED
