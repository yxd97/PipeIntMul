`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9vUaPO8g0C29BUy//AjVGUhTN5Ig/vj4TIu4v4gqkMZ9k+xGK9anq5gLZRMsYYdE
UW1ANMBsCUA2c3OONsrTzFAqoNhlNC47XbvugbSP32YFBeivCzUMt7Kb1euFBF3D
pLq+cazEC4GiH+K10Bil6jAplGSx6XnPPZbg0kjIGbk4JVUfJQ9dL9t1v+FteRf1
USSP7Bfz+4wYsrS9kYft/tdqdj3UOBFIUq/PToHMPO/eFpOhsZ3nJO+lK9nk+BOJ
QmVt8Re6g9OZUvB9XVR7YdXx7P1teO9wPhosPkoUWgv7S0Q6PJFii7apJGfIaFbJ
1vZyo3+n/6XvyHb8ZTyqYsINmkvJmMEUG+IjjEVy32V/3Ie4tE5zrdU9TL9twI7K
NtkL2PUQtCXScH9zTAC9k+uXGBiygCLCEsxja3R7tpIYHQf3AS9HGk042qAgsaJc
CO30Kq82OBpgWM0UZ8OGrFNdSTAr1pdROmM/DbE4KklLJxkOI7JYSrTEhVfCuia1
0w5AAjVagOZkPyuDaDakwfxlf2Dnh1tjIjPvhbsNeiJ9G3OfhlbFvrMXWnk8ZVFn
9vXbKuLViVA+gkROQV5okcnm1+oYXUbdPYhhVcG3GzW+E/T4+bWcqz+N6ElVcpeq
03rQxsMxB3ZgSpam4tUsYqrSH6FygpZjDOle/vbEomLKJ90nwSZHIPMinTVqOiG3
vpeXwgVe3UqFcwwRUSBlgCqgHdwcb6CNaeLjcvIgRGJEFYxDckcPaDz/JOMhHHKi
FPBF/y1ma2WF0TVa6ACvSKLZwL+3t5HFjettK2GV7BOOZfzQMEvHAR5NjeUgu9uc
zJGtMbCfoPdwRIcZ2gyc8xvmHt+yg4QC+hArWZafJsOAQmZM73r4W1RiXM9yStgu
BdnnCi93eMELkCPogbiDlmHzbpm4ocTeNKxSyT0zwZdL1W3w8xIxKurdUKn6702i
Ics+YTCGHVtM0IcBnXgJxzut9zg6C7PLSnX27qlrBAX0dxCm1Wgh6oCWq8Fgrh4J
SU39Qcr6hi5oNuWGnXLbUcrubU1X4d/jPPLT60y2bCB6uVqPilAk1MVdCtx1khVR
YIEdj0F7vzluZnhb0IV+utAcy3tOykUI0SWbAwf78jdBC5dSvSF11TlchQWHnOqO
`protect END_PROTECTED
