`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/CunWNyivEuHWAt3QM+Naz9LnOYlFwFDgIWtDfsYIhoQaxMTbPiIboPCBqYMeNH
UUU9Al2yQpSlBlNL2R7vtIARM03MDwLD1WH8scGhHMx23RCa5o5jodERT7QO5CN1
oQQR5iw7Y6GIaltgj78YTzST7CwUPKcvFWhBfXxws2QsuIrSQF/qU98w/xvpidlA
by1GD8GA/tVeiUbIjZMrbmNDyHU+bC0RUrl0CkGBvVqfJBvqhtONLtNR1ZSvSqgj
yN6DQtCeTf/EofmrsuWRzrX8rcifxiEhnN0+eVqFoOw2/yeZaVfIZ4mmIZghlbRx
0S4qMKzQ1aJ8wKbkS9Eu0VuDpXANJNF4GIGUz2XltczNSDbmi3LO1zifP7PXEcLz
U8Z9OwEz8hikFVW27YgCAyY1hjUoUtk+BtHdinUXkEwIXdRXjleIKtkqoJyqvvLo
DvjXxJoXQiLWK+G2lLb9DXjXRNmLy66VAYH4b5xTontj54uaXxkOKGU1JQ+44O02
waJTVDMxy038mYsyu163V7Sb5SlU23A7pXo4w1jMyFf9PEaDFr6o3pUx8K3eFm/9
YVMRb5xRBTrZJaKPQmU+6DLiXY84fs6mP/g9+e1nxIhxcVHeZLA3DpyEh34XX9fQ
6sVnBjWoaYz4ESL81vx9AuzTpaqNHchHhER9OD7J1sWKiycEHfMLDrRhNi3/gSwb
Yq1LxlRBSlOFNNOb3vo8s8a5ZelYtp8taVsnSaMqXldRSReN0ujEJFHNu2vENQsr
J8kad7+SRAGyJb5mFUGhUU47uo9HrOwtdnmr1ookJktEDkbgh6Zzel7aaw7RPFxs
VChiREOfgw0sPRgdsspCFjBVw+mV3x0MSAMMTDBu2fbBBGW01/IvI5FfZdzr/o7n
YShtID2ucgEsVAFTrmlwGqYiQrsGxpx6TeFlLpCqQ6LPYilc5nksut0hQRcpIaao
l4hLe3RQwLvZk1KuCxvrNxauC8i86ZzTVMyoHU+gbV+iydeREopGFY58hsyJBOPQ
0Htcxz6aPgpNaeoZXcFyEVzEKNDArYrUG9L9Mxe0mt40uCDeZy5BFtAWinXphZEg
OjdX+P+G3MueuJOJh0fA0dISTqFW8DOg2QM4Gfhmlz/jLotahlAM1eZlNAiUOvGe
RLb6Lpz+nLqL1AcOY8BDJ0SfJfZaRfr30WYPR5Y14YF6DtMSGJ755/Unh4+9Iq14
VIYp3DT0VHRzj1op9iCGTLlZiRBuURZm/runjavCvh14wpUVl1QjGv92DE2iCT/r
5gETDLZsDw1tenY6hhsNJn+2EhWjKcPhic6i+1VLnUNO2ZPSzgqUdw9mdGAte1VO
avlTj/Ap37DYa8DL17ErWHqpiuA2LbKA34wPyn239IEgWmrTokENsfpIAfCLY/d1
KSe9ybqQpSmN34p3Yg7g+c/4dDqAFfPCxmD/o/+or9b/OYTLIgC/5TENl25wffgn
lhloWK6OOad5cth5qv1c/zWEMVME4ZT0jUHKzL49fSZLZjmaK0DkbCyw1ubsNESx
EkWIH94e60vYEI0x1TB5xxF7DsG3Hvf6OQ4YiZTBafbJsJXpz9wq47pVkRr2G7Of
n+wkewh5AsvAUTflYY+ojJeB33JWPsMTH2r7mKodxWV7ukvgyOzCwLsogycsg5jc
4wDWckL9bAGj0MqEJHpvqULPCI2JYCapHCV4ptW6N/cIgC3FZula0YPwy6pDS8rD
V6i9epDrEKfPE0CDUTGZz6sejmniLlm0VTb5FohiphI29Vin9NqJCkUAqStfPe2A
HnC++nbyYxp45pdJ1CgGcotWqMfZw/u0x5wBROLOkZ+/Af1li//lx69/gok31YnN
zqguzXHsIKViumeyLvGVq6pSOMCuJyiimel0dtsQ1m0jqu6ej77OSx1bvcZGtmHd
K4xMgQjjiBWzIo/NAkonYi2VKny32C9wvAeIXCC9OPb6EabJWV2EbZfS5v6LamM1
CLlCV9LDYV+MQ7N/21CwsrvtcK8RMlO9V+2EAd1yOuD1QiEtEMS5E7p3VWwrm02O
9tmpVL/gYa0oVl3pWf0ogSGHEDVdhK2zDVmV/A0VwMqHnvzLn2myZGcqQUtVcB3k
oweh6Bk29dtwdzZWFCNcoGGiK5muoA+mzz1LnU5W99ooOWj+kQcPum1iqmrUKev9
u8sPzso0+xJz8zShFwXNvtFKzily+qT9ogTtckavIw6dpdAZhp95qP0s1kJVqRPl
mUiobls/hrlweeO5eS14fhrXyQgsReyVoFJNsaWPamvBo3ku3vNEkXejLEs7FJS4
AvrSmiufSpyfXfv95pqhTyUck+jLsAgkCsTUmbkfFRJUsxPTJ2U7fPlUJO/ofiux
BFPbvQ8UcApS7+vxkCNppip2X3a1xCpSuG24ucCreopqx/zYKMYB/zR+fLlhg177
Wo/VRYxiFCg6x9m6CwNr2PNsddlZgOQcWW0qkkBejOyl9DpHEnbiuPoFx5e9EeiV
UKn1KcH1Zx5UKiEPNvleAEh7IW7ekCP1LKf/FK8yvVbkQBS9SCDn4C+5T07fi2S9
L2wJQDnf+w7Zns1GySW1WnMKV3QDn8q4UKj6IaQxbU+y6YWvnCC5v61H/TtT5gwK
15XzfjPkmWTdDDEfpGNjHS59qrkRPvoHtwOT0yu+BWDJg2glrfyVwbMXoWo8LfMA
kBtRiawUkLVegdzf15qweZxFhwAEJ6C1pMvOqZErMhJUGmAyzxS29qMJFurlDVwm
pMSILhHCwBYm/aBpg13cFRSCnj9fYjSBe+N2Ce196tbd/oiuFKnvdTjB+03wj1Wg
iI/yWSw2kjQF2SaGPALqqq6cb9/wJl17ZmRgktpMqd5Nk4KFsKIQN/my/5mFTNAP
p+nuRATgfLI5dLdLJh7myw2ZLr6kK/nAhL4Y3nOlRHoSdPa6Jl3iKblgaGnAuovj
sHR0OoWJAWA0POQL8uj3NhKK+S0tHFawoIj5GhTvuaJDEWaa3+Kc18WhUlPpPUKV
a9w6068+dwoRdSbF2OvHlQMyNcWfKFwjNewsFN5lwyv0PnTPIZ+jC020YrFjjomR
DZKE4q97NUfMV0y1CsJmLmMKjcn6wiegLQV7FChIVRminmea4bHu5P85nm+jgODf
YYPIzQQ677ROOk0l/VDfaJcj9Q2ps3mLSG1vcBTpt73JA9GNsGRDDwPXiKzN0dGT
aQ64LLrGOjF1vH/DDd5eL6wivnXdptsTcMdcHJaMwbI85eWQdZXw9S6r/4byQKTB
rVdiI7VKsqWrq21xY/XT6iqXbG/eTKovYfGf//nQbsuKi3UvidKPm2Zv3eoYQXu6
f/B6zyMRDD7GgxTCIfAqz1ZLo3t2I8dBOd9vOSWu78EmIHpclWZiUpP+up6ZBmHN
T008PV4nZpII9jSInAca7u8b2ziz+BW/6KdNFM2v3P8K3OtYSnLWi04Tv66amPW4
cSC7mMdvtagsXiWD0OyKP8tr+ftCAn4u2cWASsPjSivXs0bGgSfnNkU1wmSv4Uul
ZHt1mriWrsMGgMtloWk6Y9wTZVyIrB4j7b2l6eI0gUDMoep7BG2SgD7SjUi85pIw
19ZdcjuSeAF4XEQUTBMxnbwAPdVEyONRqueAgP3HHuF/K6LlUmIoz6LXoWG0XFr0
7UeRc9t3CIKSFTqScnWKjECbysEWTLXJk0b8WzUVPkElIW2SV946/ngQUqQxIzV/
QuxajntEohSvsbsn1z1RWv4mglxgbaiFW/fxZrLtHa/QQxdDmh4fIMSrXN8N1x4Q
4zvnphmraSy0avDi6YgwpT34UXI92BEGZdj1O5j0iXQKqjNejbOvdBuO5GY/dUHN
+GJQSjluIfQlerBGj8ngK7RtxqPbK63Wayzu/D1/Jt1o/5jCcny7+ggn+Od9CBw9
G6/oZYEncP+9+jMGOptRJmmYL6TzuhjU3Dhx4WNmYJjRgXfAcR01WcfHUGnGtrg5
256yv/XcrGZqgGb6QkJoxvvZ5/3lN4tWDPvRlOGIRL5ArLWyiN7t5dbfBnktDD0R
KOLAOXlxzLEy3obR04ScH41rfnW4SS21wnEJmd/kWwrcaj8MBdCtUz4HKDkkJw4/
LUTNnNBLgYs4fgFb6OWUSgsXY0knnMiKMWXarLYkURQtBBfhdvfEgw6YR5UH40a/
FARlv7O7zPaxlk9oYxx1HSBrRDesnPaPBmk3UbCj9WM84/gvTk6D/zXw/eBpOBpE
4Wuv3DRVf6ItIAMGgvuAF3DWjkf0MZNKHB+4g3SdaW3ag/wK4kevZE5IjYLbXgml
twGsrvbWy6PaQQ9d3IvyQaLz/BzMkXodsTesGEmSDh6CpttzjLOZjMR9ir4nDqpu
xBBaWqxUAwJj1eSdHandJa5+0dYDCXKL/+PklmdwzDxpaJkB2PSZp20xk+aL9D/p
F/YyoZnl5eu5/WBJ1i84di4o/gF+cYWBvuFRGr69BTChEkeqdTO05XIz2f77aPqY
6D2U+w7LI2PBXNp2XkTp1G93ZYfEA5jJsrdldu0lPybkPUO/vpObyjkkB+2/lOPy
THO16y7c7UZTt9pjT3MAnk9uSK3GTIVq74Wiru5jPpvD4dyY9Yf+QT+Az7Ll/U8z
8veKEgN7TlLAU+SLfFLXMxUr6Pb20IFMqtWSvAN6qpjIBNr1xfIsWoS5MD7Dq3cl
mu/3mFnv6ZMjffRHcWeDZw05n0K0q/vvqeVCbjkQon58MZDtIsNTzSc6NnXq75az
1D+m2VaQNpFhb9LXnoTzBMxiKVOPdA2nrtDrLGxh8xEVs72PXqNFZ905ZeO7d2zH
TG5XWwCWUfK3FPHlJ/XyRltn0Kfl5eYOSbDNBQjb+v1plpcfziGOnS2fcrPAfIxm
la1+z+B8z+z9Fo1+cL1QDLODUXpn62R/f/gds3N6MyNEtOUnNnKJa7+RweHyhbAO
dRVcAzFHKrl1Vsd7ZGroU2ZYsseF76XeouMMnBOg/vVa1h2RfwQiI4f8Ak3qtGAK
j+S0aWowxNNI75QUKkfXNG+GEHAi6baHJV5qiNBGPi4iIRRZeunxRbQ91AWcEU6W
Z5X5B/rfHdB0OrCtfrIYzyBt68CCROdBOXRfQ7BDkmnXstEC+SK68EIwCQ9lxpcf
jMRDVi8B1UkA8jjHxIV6QGauLASw30bjztSCIkTsKRgiZ0qujJweNr6aYO9Yz6nq
PjnaylAZubqoofVl+1K2qYQ9SwL6NEQ5b5egKm/jIxz0ftu6EaZYuYMGzHFGRpO7
JwLhh/6mj/EVHVoLqF6/7eth/BoNpqcwgF7QdFiVpY4uT+4tEa55Lrc8CivkW+jm
KZysjIEoAGA6yj2NKWeCkeuNfcpFBg08/xczLbGno0PzpRjmHQFTofIJYjYrv5xm
HeQlgwtOlNFYJA1p8wechNGB4Ir/7HNNwFxpxBEyhirdv3rZTSoIGsQDS5PtjQZL
gkIMt+v5Otm6v5pyrOEfundJHdqIOr8pkUacGmhpA/LA3+mb6MV2WgetY7dftkQ3
+iJQvbaVfQPQ309nlcufxCmDM1rn1GWsqfcGxHKLBoNUyRt/yT/AeBFbhm6752LW
nVK9E4izyKX/b4TCu2pA6GNB5P3zYCL0NelSnTDXzx0ulMnTcBug38dfVFb2KZG/
+evc3XeBlxjzT9mrjpNM4zRzvxyWT0QpZC2EJ+XG8+vt1myigqi5UPpeWJnuyOzG
0MKxbV72Qu9OWeKoRvMp+PvX6o6e426EtOAvFq/UkSXWybECVWZUpMLPuhOhe8Cr
4aaouu1T7yEImvNYKX/DQg==
`protect END_PROTECTED
