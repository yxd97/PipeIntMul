`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39eb2dOvttNcc/8TX4+iQevUghH+2ggvl4hbsefCh6EFGIwEnWqiPCrCwPzhVNw/
ZvAMLZrgRH53VE7+b+T1PPnhczMYwegB3UooWfGQi/UC/wjqy4TadKJrK1cq7LLo
SdfaHXxhA3DXgVN7mJY2MK8nxTJbsYF8JA4rDAH+gcCDc4XMY7pALVOpMyKTIuCV
7+xAJr2QgflorRALM8V4EfK61SD7YajUPl+KDtXT1dt7LyrFMCom3hEj3orB3g08
XRiqmr7gHYGJKG7/179EOOpEwUPco5qKHWpnpaHmgecUEmRVBJQ1rk1hJH2KeFas
R+4Kk13y7hwO3XfqmHB5beRlKSpxJcIlBRzm9eddOY7D67NyxxruqR7cBxhMoxHP
bq3SWJQxkYbWSmHdkgYz5gVG/SOE6w91/oWG7OMKX7DyJP+7R0LC4dVQH9rC+0DI
jg9tMDxG9UriCToyJ90YyDo1k47qvpTjwg9P3QC/n6eKjBo2ZV52Wcd6EjNjGt9N
Jf1Um8xPtGNhV9yFdqYQnS3N0ZWYO+WNqP0+O8QfXS17gFa9rw+30Vr4DobXLBI4
oT484urW+cibkAA4pzVzEg==
`protect END_PROTECTED
