`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XHhPcUOF7vnvCVBie13N19zLYH+7KlhYzHHkagGEp4TkMhV51Vpzb9QA+hNlDUsG
g8eSU1fZoLmGwsrkHhHFs2U3KCE0el8BLz5CQmGzuDwUFVKHFVQXtrFBafhV3AYQ
emMYs4TuQlJo4aYuj7RP+BwVnT8/S6wkIUOgUxNPlCzxD8mSTsvg5cVNSP8ukrto
Go7cp4ZpAM2aA+288kk+6Z0OVV9d+OCnxpyvA9ZaiqHY328+n2NgULdzYF32geiS
sr4ARVibxk8COaoSuFLpHtYAMupRl81s4/9bGWrBJ6S+g/0DVk7qPGybzEqeALy3
7+GZbACFQNUIN+ysH9DQSNV26YJNWUlNrbYpVQL8jwqrRU3s6Ev8ttdBHu7TjIG2
0kXuVFiDn/KcTg8S++kh5WVCD+YjzoMI198evrI41Cpui7lAkGus0KemWOeEdCnO
psYRVqQgcZC7soAk+MF4521cF7VhLdg2fshe6KHLLBRqpXrCNkxf9FR6/0M6HeJJ
UeGwOHhefcnSuQ0C+/WdTAlyLIpL9qd7tn5mMQtsWWtWReqz+uRH1gIB981uCiCA
wsgQQNJGTCGEVfWCvIMln1DUwWe2HBfZ6xceAuIbycEKknCPXwnWphO9vp9Hwuwc
1p2m4QWEQp47G1c9fGBkvrmkyYWZKjGFHYAMoOM+Da8+EmFoQWMacgQmP14MGHQ8
`protect END_PROTECTED
