`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jbS+jXFJnSnJA7YLYt0LN0TPA/Wehe3JBf2h1SMr0p1iuN9EWGtfxYE0/PrN5csT
l6USRPYgOk1xLuWeQuztYkVH9arjnMzuKG47ELKy4EU/IZTxjkDe99uXCfphaWGR
V6uEx08RZxpj/OfeTZU2lomzLM5uIADV2owFQoJ2X/MlYj09S47Lx4qMLQYuij+8
yyznjBQwnWCYLqM/Q3C2TquKUEyRC2l+rwHc0/1h1sk9d0A2OnsRzF+9fVc4oGBO
zq8zc6YngQ2pkq1m+huzQdn7Acwv5oK+f/lfKb1B+8s=
`protect END_PROTECTED
