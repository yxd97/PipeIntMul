`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iisKag29lHHPI1HQAgFaGL6XncXvKhuS9xYkp440lNX0CCIPyWb/ALlBvoCELqbv
3RN+Bt9m1AEjjXh08m6fEZF91KkRULfpJwZSXZQoAMFCOtsx+5t0PfvA1CmZgO04
ugCFiv5za9usBdwtDnOe8ZdeVA//2a0UqtvaI6WIbcmy/Zq8XlU1/bSG+mx2fXz3
LQKkzFooAV8cdKM/trJadt3GyjojO6Svt/1MyFMsUe6RAJQqgmnyEGB5glLyxopg
wcOLBzm2Gvhg/Y5zlhEdWrSW0degAGnpwNDlRzVjQ23KWYdIgiqVgzH3KFonabS2
1t0J6m5Kc8HDlSVmmEdIYIVu9Sn4F5Ijq0lnw7SvfGtWbCaje1e1L2U1NNRijOsP
d1Ob7AbSPnY/a+76Kxht/Jqnodn/twwTrmVm4xMbwvHWju8tzUGIuxmVf5mIuz7E
StLDobAin2EAlpTpdyx8ig3YmATv2h79TNABOoGjvzj9DY9+ifmIKyXAujpuYV69
BtapesMh4dlj8kknp9fJn3LNJprALloKA+JInZJAncHUbwkOfMTfSqq6rxH8DrX8
xWeyPLwO1cMM/FhkjM6ihZfieSdhAzFi9GkBUHmOhTc4/9o5H8EdrzPsUakWQWFY
SekPzFcBIr1k1QIL502QoKEOEU2hQbDfvQ0uRUd+MleJY3W2vlq95Xjgv91368Bz
dPdl8ctDLXIIkhhjZmdfym9yaz27H/DY89XQXez2olsgGdov8yILLuN8FiCgxUx5
ew9rCj8nJYisL9p+RYcF3Q==
`protect END_PROTECTED
