`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZPMblhFnLri0f5EgCf2Ym6D5EM9+yL4HTuwA1Y0KwZtESO0MLg9raylm5C/8Sb4
pwded/5D3o3aQK1aYoA/MbqqpNLk75ZPBbhAjUhHCj0jD4CHD65v9JbGJZnCHAXs
6eaMaMTiAYJ3+iS9rjlM2LOxpVD/+ucbV89hKKVpUMjoYId0yqf3jar9x3D0kMDw
RYGU8GWb1bXfCU6eybTXmgbj4PHTfiAT+kC8U4fTNUcDATes8UCHTwfsg6i6gNRb
mB9VYpDHElVScuLds8WOWueBQRmVjWOxciGXblByegKveePaB09pz8ochkpppr7q
FYhLF5+U1/LF/NAtTF8B2QyPLvsUP3fGKpSyVBfTJiaLCN4x8iN5y3I0UQ/uZwmB
YUktDaMqha8+j9iWwj9sczON9P0clAPfJO2fOX1vwuxphZxULxv+270dj4GNdAN3
b6/r2mx4GM1+P6+htCxMgsEsL6kAu4yzP5mPJWjOebAnVLmhPWuLAPDz9jm9Nmqo
KrdUvKSqi5d8McdVX+sGBMKTsysJE0Tyj9x4NprBsnIFVnab4CBdRpQSYCFWEE8c
UrDBOXTJj1v+7IDch2GhfbKh8Bi8clZ+KIlo6+RddASHq/VjnJHFr0dZVQkDnaad
cPlPEhRHzm9CV136QU63hoiQq3E3l/LniquZH3VNMGwVDTQHGzuMraQxms4+ssIj
wpZyPK/2mSnQNC6+WFrc9EQqm+ilT/rpY85it4r1lG8=
`protect END_PROTECTED
