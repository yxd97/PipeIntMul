`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UO8pb7ticRJ0fgvaIDyy/UUYuoc9XqA+UUtykjYFwprOCOx/Xb/3l1bFIH3N9DUE
nEAi8HvooqsY/mt3hxouvwo2clm7iCrh8fRgYNN9duwk9kNXcjBRNB4/cIiOnP/T
bjZ8Ni+I+/tnh/GND3otuPC3KdYNg83WlcVNzaoyev2FRUKDLLNLCTZN2LEkYwTu
co0M8NdsETxUqhnyUwMf4PZm9z6Qzx0d+3PLCF9Oe4nGGl1vAA4Y/Rl7AMTCPK3C
MoE08Wd/vVjJAfcLn3TtITY66+RwX1UNwG1zILfsvoJasck//kq7hGUXHceveJwi
FmQUkbjSqV4ILUfWqo6RXUzVNvL3W+Ow7vtcZTTo0mUEqyJsbwl5FSOspfZjP3dk
szIB20c/qvnaWs6Utc6hA5CM/yCFqnl1Azt5zswsivNK1S02Ks9HPMPZc2uiC2E3
Ml833+kEyzoKjZd3q7B/sqWGhCR8DgRZRUsMiHbtvrTAINZtta5R4QA8Axep0Z/p
JbEDO3F9oNqVnH65lpmflH3ikYmV+G6DdzUfZR0L6Y1AD3pEMrc/D7AfrM1HxT0H
zhCvnipOXvC7yY+s/CETibfh9tAdrjHGOMDxZDQSSin030NYbw2Qk0z7+SSgXCwy
1aPEAyTBaELMLL6SOhn7eA==
`protect END_PROTECTED
