`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Z7EhwLabpgoaaAZgZp8QgimS3KO+Hvk+Rq4ItRlb6zePPZjkkf8Wt9GVw/NPPyE
D8FxhCbS9KaTSc9oq8ZW0O1uEwulfXtQTCpFeSVAm93MZVjBKvqd+FynpUEX0nZg
MlB7nHtQBYLj5dHiHzPXw+4iILinQWEJnk05LoUoxoNVmgpfeDk84QyfHfgRyGkL
9weamXheXFJ0BRWqechR7nh2txX/Ya0CA+PgXuoL2bOIg0kUkoVB532EKq3h7eUp
I0ZDXGTkV6fcmdFKFvPZ2WxYRM2y17XyCyQ23UukvNJVpov3IGAyw6NRf40GAQhl
iJrZVy29s5n6b538FdDRJDeidcxTS9mpdG3CfarAl7cvrlTGjFawBvgUQbI4oDgw
DjSaFoSoxuwOd0JhcXYLilhjKodTUpCQR+FpvJ88+mh+lm+S+3L1e53D0+kH2eaD
tyrRZ+xlx3JfgKljvAR+kg7ymft/Ml4rX/shd/+7A/e7PSCWUv2YAzxNnTqReA9o
PMkWxlSNUETLWHPdjqsydxUaANgBjf0P0mTlVnOcTuH/wR0OmPqZCn9ukjyzhCR+
OIMMF3AWOChhd6Qv4B8VpmSnp+DwCeMBbtyYzqAfcQElbBgGIEA8OGHJY7AgC6/V
Sxg1I199opjyrqZyeab68coBbkw1ho+UjNJnNd2QuH7BU21/na3oq4GOO68JHSEF
tvKHuPd4x1PYBpwm8UNNaTNPToEYA3iAeDhPf+7TqS90pFTJfnV2n3tETnLx5BY2
JkVUMh0HqonF4xqFzXcv5+o1C0fm/Z7/JJlsDOhEkhmaRs79E1j+73IEx7oKW+7Q
/i76Yyfg36vJSeiN9fl4rMIOe3RHEnfB2S8ioCLi07SwC4JdA2G4xvPlcItnXCUD
2JCSDPxB6n6H97kOrtLj26BVeKWcrdVU1QUJ9mGR/1wZoOsO4ZwQsuks+q3SvKDs
C8pzeB+i+A712g+HowDR2w4NIo6Rc/wMerDl47ZZa3s3aRfkPOGkGuYmI14Y5B60
vzDVOjY3XK/FMlPku3MmkQRh9JOpdBHJbeCoSGs+7blUP2+OiyinpYLbd+z8QF8W
IR/EvR9HX5AzVnEhz94qYoTfpUnguMfkHZEaeIfrmAbFY7HVEBtTAep4LZVPlPDr
2P48uDsg5KIjuTzKxqnzuM31msmKGy5T514F5uO81SFtabcKMeSPcdhqVNJMbgLE
9m+WktyFN1XaHX59T9vG3o5rK2P5CjtWmS61Sj7ofubgl9zpXaUPIJSBqh1AzdUh
t3yIpTqvNogWVVBoUId11o1BLxkTUtQWeA2OaSl+HnD5vB3fG9Kd045eFJkQUoSy
sn6beyfB6/Hz5RMf+ha4MH05hvg/WouuFgSXbKfelW4hAzHLd0NnNLX2TAwmTN1g
GCZhFSb5EBDIWZq3ZhKq5ySAOYbz7hZSY0x87XFZAanjdIaex8G/pno/eU5hnTqw
4sQbKdSEhswOiPG17upqYvdSSVatEueghlAh26/rnZi0MxTFjJa2FbGWGj7CQSGH
DY4noV23T+CT36udZX7Kf8aQcFKJ4gzffRmnL/IHyel7UtCW1SmPtRu6HHETO1Om
BJTXCIzCfJG89CnG1ulpXFhRd2UoI/UigPHgZFhzN7Uzm+Y1q3oUp+c0MfkdMBfi
j5WKpcvNvXd6Tntm+dwgaOO1/XrNqkE65FL+9mcE/OQAmYx2lhBXoDF233vh6npw
8xEZGpDHVSW9tHOooIsbbVuP6c86s/A3CHL4/VwAzriIri6JUYu2ZySLZCGQiBTu
VUL8iDnpbzvA2TeU2/t1aTC6qIEyMQ1+OM4xn1MHecY+VErjUzUH9gP56jOPl3VX
eqR18ZTjqfc8bGTTzHsNSV439d6DyrHy9LgVzW/oQCy1A2h1Rb21oAghzyhXl39M
uBaMOjGoEK9VlI3pSn8KX5HB63lPy8RQ5IZ9VTIPPRXxpYWyBXcul0GqC9nWD9zD
MWqPWgX+MxQl/+16yFgn3Bs1n2U+BTFNog7S/wdW+0JtzdNnXQ3OgTXscTL2hNIn
/V0OrF2fPt4Xf78/YGJ2JTB+sXbSuoCr5Roo24KuzU2mYMjspE9YKKchs0PoDmD7
vdb8y6lDXmeUXDSuUD0ARcPI/NbB7pgMEsbRgUyJlwI8qMNJPheHWB1bhuR0D/cX
nvzfPAyavJhawQQYPl3/HnVYQQS+Vhbx/u1UmDLf1mv4OQBsc7632+EB9K77elyd
G21dT5rfcgT4FxLgDz3TedtDt05fkof8WHG/4ZH+7Wouh4paLmSzeGqdpRWmS84J
XKiWKoSg0R9cosAYRZQWxdqEX7JPGeOkKGBlIiem7v1KawYdGBjPgJ48bpABStYv
pRc6hcEWXvmKXgtsqyRtubGfCKZNTK7vfI5T6Fi0QVytLlu/U+DOidn+f/HrlWU/
PYE/51hd3UMaw2FWTe4d8+V8oJ2xUoDw8fIdXT/cXicwP6zUNWMGQjEVnNods3sQ
NR9oR0AZKIUgesUjFsl1qbzH23j4izCKcEhduSd9o4IDR8Ch4Jl2g20jQe9dWROx
m1gHBHOv2I2p9N3Rox0Qr7wbNYDEItG2+3cjhmyYE5nuegX9pDbpYxZp01QJ9NqH
VN12bOnAHgMIGpFIsZnGj+GWDmo6wxSqhmg5gfOI+mPkbSi66jcZDfsyDt1Kj3nO
GAJVWhU6EdpELEtprphLipIW32eMi/ebF8KeJ0mP/GtPyAILXUVOAEnRCv7OpAeG
za8sItFIARpY+TS/lhV6LuMhnxvyGtv4Rx8LUKnH8mIx/GpK5IFnhoCJGGETHpnt
FVU28ibDhVTuD877tLsc5YNAcHuzuQ91p0GQEOv3N8HzEWir3k1lnQCZ3MO/Y0en
zqaM8LSDtM8PIpi9ePraFxYxuomWhqzL6AVne5qJK+4ERwaW9a6QUylKqCLbnK9Y
g8aQV7DPQuq4z2ehhu6QggFi13eUR0EGXLS89JXzjKQcbhDL5YvWgDITogLEm5p7
8yrYLdl4qG3vd3yHQmXZ5fV7fC/20gq5iMnFa2flyitHU8gxZ+2+Zsy5sd/6RNRk
vkHdTEpJe4z24c5wZ0qzG4Md20Ya97SJlG5nPOwoNNmo3qpUkQvfYyaaxCa1fVAu
rcXdtQePl+8UeA9aMxxq2P/U0eq7/+87OmEIUAQ8C+bBZaN4H/Ouzds97OdNl274
hrkIkdrY/3pSRt5ZxSMpDCpR6XJpSFUFyuBZ2QaFpkOSo6+qCJwxSZ5MLMvFJGJD
QUh+9n0GC+RiDGrQfgwb/jtXrmY2rF839jAs34mQj3vA+0NY3eCqsMdYfx+YY2Oh
kayWwVzI4GgVfu5gtRkX0QMKdacJRHsfXhxZXxI729Zl8zZt+QAyIfT4Z+y4F/hZ
e3fnHsTJlMp41STgmJZm3YrbUoImvhITcfCQa9fOtpEvItEI4dmyebFfTPBwd+fe
fjbVgQVzIENx+uMUXZwvO/kKT/QNRO3/aPwQun6yDCnQ5APpzpyI7FlQC1f2mw2B
58ZdyUDwdxAXWRBkLnVnq0zCxWoCjsgHWZuCZ5BpVuZfuNeNajcHr/f8UaPeRh2h
R9qXR8IKTgs5z0DEraIjA3cCEGWcB2YocDz4KeNFG+mi0sBolCGh1zwaRRZ8QSVC
nF1uTZfdr5h/O1k0a4v9NSatvA1av93w4/SCTo0N0fj+XZ9XbBuG0TWP5nEhIUjk
5FBhmul0qdOYdank0dSKmBQklImy9Ln0EbtVZXtG70dNmDqJ4y+D5bOCd9Y5mdkl
iAy7jfaR8IDNPcO5GXsGqiGZBcseHbsAMyNoUpMRsD374iKaLmHdHaN0FS2P9oDw
kdWv+z5HYR9GWixA4vmynk0xrphw/AVl+IQDUa/LQDet2byHRKNu0k4j2O9K4nap
lMTOMLy1BKdjmELbW4Fe9og5RsvhbH01/HBHcEhSOZrxjfXXUYRi8KouXz/oJzIR
Z7HmncSbkWapBPniFZCmqpPVWiD1OQWT65fb2EfYvb4jlKJVHmZMwRUonafOseOQ
S/MXi/4SybiXvVJTRhs0D9P6v7Q9+nua0HQecUSCKdN1h4tqEvNQB5kjSmI2aXTE
96aJuIHgocTnhXwOGzKj5AxGfVtx1ye7JSffrGt/+b9lakLTpfAiAE/O3TQlunfq
e3Q304W4TYFgxoPkmoXjWFwwaC2oFvtg1JQTvkWmkxTBrm0EZEybgsaFXN13+RJ6
NlAHLPYiXbrd5qQLjMunlhoNsSvuD4i3r53BNqb+hnzGEETQ/+LiCWFqDcSfCv7l
V3KkoTftdgOKpp02KNL+BOzTskuobnGr9+3cGNmIAg4aVlVv5zVswqWBlkDFSzOC
vFgEge2ZB7g12RFq0g87y21r6grribUE+49sGCRuEbb9JwAMG1VgTqUNUoDjOrc4
KYUVf7FGEqzeTf0PQ9NE8rRVnG992CHAn3b8rQs+Ob1Q7relnyumaAbVpbIsu0Rc
IQCvXWA1P/c6YGVXzSnkmFNDB5OSguVLSxRwIITAufQj+XsKEZtGboPy71oe4Vby
uHoI0lPjap1G5f7FvCszIg6usHi2HxZVPjnoyi4QrqUogWBGRHHcwlfiJAaE0ypZ
S5uDu7nmrribCQM1ZzKTpvu9d5hTsSTiKbRaqbAa3l/Zf1w8+y2egtuBlz7H6P01
ytDV2uX5aiy7nhVvACqCo9BTyA+rjFyMznZlpg6pIz0eY1+2GMTgalkjNA1ZV2ix
w0P333W29dUWodLpwaVtNm6f+1vXPRoBdN/WQZVr8aA2+L7+qZ31Um9Bk6UA1hBw
T44sOw54lW4XTwLLuN7GofTPa5IPIGA5a4JLvAQ36rvqUpNfAtsSprH6VZU94Jty
KKoqtT+KxhDY0fSiTRiDRr/y6YZLA9+dburPc/79fgD13xSCrxosfTtVysoT3U+6
A+VgHiAIH1dAbP2tzGvX3KU6zDnBSgUSlzAxOcDqv8Zy2pmWx5CcHIwwqtHuEjOI
VY1T6BCESR551DYf9JALaMuJe6grzQ21cP6TUjabuGXwhVllRs+eupyYaPX9n2a7
5QnBPDmI8fFkmGIqu+Em45IuvcL7QdGUSqgSnfeFY6LaZSN5NDuH/YM88j94THMS
TiXMF4eRIc37w+Cyb24oIrTKHz0VwjXHzBZFJ3sEJ8Br4RN5p0G+1o+oi9zj+nY+
2WPmJjaT+AdFe3dM0h5ACcQLKtmOyx99UU2/OEkZ1CH8iDhPzmf0TpXegW0cqZGv
wwCtPjRJQ2rEnP5ZBlPlZwYRZkK3aDaLrjxfFos0ozMvoOtqBXRa25hQAbnTR9x2
sr9bhx7whRnUNO9zFuHeJkvJ2Hd66LLthTrOLt83I1ErAZbUkKiUKeKMRHh4VnFu
sm70gvdldFhvMNfQ7HyySQKb1skVUBbG3WuZFT3I3bJjxfhC8ZNKxsL+6YqgIMIK
VKEnB41VwrQmDWcvoFYMriROe6PoFiMDz/hfob7hGhOdNfQn6C3WusGiYA+6qLqN
/Q1vcGnnb6LfDWwpRr+M0vFYRDUcIlWqCpkT3fiSAtDX9ITliKPaSg38awOJo1ts
/T9kQY16dX61gnqkoVglI25aZsDsHqjD8EgPbGRxO7cQ3yvbu1nSfmp8jYS5sH3G
hbBaSZQpy463FQBHCZOEKDdIJye7BG1OII0s9ozdEt3MuwrEmjabt8HXoCyLNjvR
kizr5kQyYTC7sROfrsB/A6YPeL1uPzuTGIWG5N5s2QYkKlYl65CobLnOmw2fbStx
/yqjQoM8oLJ6rj/r305FhJiVhgHXFhE5x4OERxRI6zCyoH3niGLd9mwN0V7XzDdH
DjfUspLCi4QTX73222vANTZKHqPQSQs3ZGrnlbUHhFZzN1XDSWuXf3kMe4knKPMC
EwEZ6tGr1NlTh8ZZjBHcwgQgNujXwetRKhGu68PZhI+L1bqQopd591u0dzP4ZIaW
YKUB3RDKLsyarlhPBvnQ5HfatjSQBJ6pQM21P9kOFUanShoPn0wI/h2Z+DwwITsw
uX2z0Is6hXxdBBF0flB8mNOUyJm5amUN8QrNVoDq9pDjElBN6EAC3k3MCr+eCYpf
uMk05rW9vHy0WYVSVqWRpjuopRYO+7k3MzhQC6/pSr3042Vb6jsFs9w4rQvYid9p
Ur9ZBbWLTHtKKQ31dXhIuMyLIH6oUz7XLUny+b+BHF61A0HnE2KL5NfQjB/1uv3U
QBVCmz+XQf6HVxoTWpygUgUlm2y+ldWGSQPhU+uv3ooUHAWORsw+XpyCRzo10Ugb
HM+EioewEKEDK1ZFC9NNk0om7VoTbBeXjkNjjBGNXd1X7GDdveiay1CgIhINn6H2
3kJHncNAhgBAhomi3HIIueFftNwGEAHpUEAVRHV5K6iytuWYoIvVJD+hYqc5+6/x
OX0Tig4o2cv/fiDC/fOwS5rczeITLdVZjkPbmz91tLJOLc7x0BE/4Uu3eqEBI1ok
H28MwBLzJcUhZodqu2p4EC7ZQHVpwi+HxiJ1Huo/y77pWYqCzxZfjGy4uUCA3c1f
CPIyrqCFzSm1325bu5AW3AmdL4zBcxNIzJU5KmeiSwbDIeMw6UlRNZ5eymYP4Dl0
btOW1XoNQrqhgjzNS8nKjSRpoiXsVnCefy7I2XnlzjjMlPjHkRilKdlMt9DnPSEM
xrFQ3ZWRMncjYSmMadL2xL+kV7dq/VJrhB+WfUknXm7XW6eRiWJ/Cnp86irT3qsq
aVjA7gqUnpdMT7/NixcpESeNQCWl0tROpqZ8SSuQa1sIlbemAhd1g4LWyEsGJMQX
pJ3Y8xdHXwcDWmG/ZTRyLghMS28+OA0+ii8wDv1DKEjGAj5X/eqAApqu978LREV9
UGxM2ZUwIAyJR0Wc9URFgyhBR+9yewE8CujiGItXgRkqIU1fL/Vc/QVpW3yRTw4d
M3qbeZQOqwfrXwejG5gc23jX5aTfMnFv4wPrTcwNSiVctmRSTg3jYAAtCP17DN1x
HS7BtgPWk7e43MBcsyAx+SGwM/izOopttR/+uMrPZXOAa9xGGdOXpO/Lpl1XpKWs
6QfYWYrgXuw4FmO0IhWbErZJCgztjPJgmqGlfM3994aQb6X9QBJOxhgyGAlfOK9d
dhe7RUB2DXHNLvZurPPzC/gIEApb463qVAOdTowHzU8XL7MEif8Fs95UU8AJChN2
rd1wGKdH5MZ0J9QQBetaJP2SotKJRl59Ys4fpGWZroEDti70dMko1astQxR5QR9B
PxcyEIEsL1fh/XJcD8ycIk17AL+XsacEgdmVIUDK+BjfP+SRWR0S1m4mv6lXx36z
VmXBHue90nmDzrR8PCVhdRb/RmqfCuxigUYeJnv+7IiXEgIKFdHT4ozXxEp6lfyN
2CAfBfs3fqNLFkPu+uWQYiyJ+H6hb2GxgJFuIXT2QUFoYVplLv+xPqE71r6Rs1ND
oBY2EFDCrfW4cSBXWzsm+kRnSbzJ0bdZY+DMBUcwafZyx/AmO4JITLEoQf72qiQU
qCxAmUEFzMu3MM5wO2PghkS8GgBGlP6JtWU6250mesBEEh1ae5vKjVsQHh1HwRoV
vWN9+TD7Cw9dGQ/RFyQSPv51lWvX5cWt5sCQhsM5k4KpNvpElTSlQbpp2Gqx93r7
qgHcp568XCjHp9d4WuJKuH+DRBSM/NcL3wdpubBQPLwar4zsBEP8+CXLJsU5zTue
XAhvM5Q314IxSwPfxB5rNQZQVgtHelsPONX3f9lBTPaQPOiLylZbOv9VqDGzaAXu
6oXd8HAZ9+wS+yYzP06FiAOlgQjcUxr+KTnRjOceJAI7zUnhJxGFt0mAZ27PmA3S
FlCbsXxhEAGzgpr+LBJQFSOTN6Vc0cIU1LUAOMOL9mX/bLMcKjlqizyDceCyHs86
RSwnlFjD+mZjIn1jf42kmCHHDKFvPMcGsMY4Amewi0eKrCJIhyMYRqcIeJQHPz3D
RVp+Ib4chN6WF9jUEX2bO6GDFH398KXR3wN/X4e0sS5TBTey6EtTYyRbnv1OCS2A
u9pjpK3dY6OhBIBNJkCLxDteriBoAnk3cHoLFCEj2sA4hRa647F89RHxgWeqtZLn
m/Tm9uWzLLyzRHBTu0jMv3nyWQZ2LltnA3oyGJ36JPwL3ftniwzgAzBeFsXIW+jl
NMHIZdTew5HgwwcQ5kW9paWSnIcfFZsAoufRjQOT7vWxiT25BnLtLxAwZNFtrO83
FGeVOojjtNatj8bgvsfVOgYVVFaB0jkLIo8YDGkSBFZ/lDLGT0LKzxhg9ExUdzQ6
46oejQ/TV15E83eooAGrR/o7PP2q5CIPWdajO1r0T5D0R8sNiGOQ34RFBntqk67Q
78aCSEwdi0LnLpkdDb12dVn7zxqab0RspEIx1CzCTf+947antoVLPr06r1gTHMv3
B1PQEYUj8ngqqRknbuPYlRtUkXCKPuWZw+M4k6BJ8PiO5UEj/fN0qSipUfq32AO1
vGrxarojVpUx1RfycBPCXlLvVNA7ca87eZe6YSY7CqYz1zZ66wPEA6lqHUmbZEMP
72DzHtufELAbHj5rL/WMgKYXZdHY+hyu0c3n3TrD+YephWysbMETOuMglHnPIqW+
ntfcSpnkKbxp2OxQpDGdatVZI6Ttngb73CWMFShGnuD1rtHOAm1YeovXVapSuIPo
lhPcRH7pEd9XhlGs18OdORDClRI9xYWjs5TN6Z1soh4s+lBnC123NlWeS8LcHag5
hPBvJOhqmr/pj1ldACvCReERqWz4TYiCbmyrUZC1DP5RSl/ur+nmym6V2kASCogk
WsOeXSZ/jMQ0+qppj1Q8sHSUKJqbkVV7Uja4TLTQqJ6NYFLdDonYSgyZ+yni+3Zx
P3e8EMEMrHfOpI4Uy9ehubB6HGux9TJldhOYZQltGGbYfhKEbspzC9/rKISNL3rP
GXcgKDIQW1z3E6Qg/9/wEYQ4NGfmFqLVTCJi7lrDecA9zAei7H0E/8Gc6vdPzl/R
PZ6XkG2r70F6HaK5viwcfjtwkehJsS7pkng45fK95hN4k8b+ZG63wAPFCQe7+qTE
oD4boOHeXsB+zRqH5Dy4518FRwU2+bP/d+xAemHoAlbvkYE2huuGvddAyt2OKXSU
tLId1BhqRep2BODTih+uEhPAYEkb8OsmlEMXOD1Xxgb5QK4y9qZ7rJApXBn2VfyL
bok2d1rv3NiZ0I0X9/y+PNGIjz9KR2G4ZkLaMQSjhEj/31WUo5MqEp8fNmhFhbi9
xBptJYLbHq4dbx52iFu/uOTl74VodeBQTc1Wd7JwrdwVyQPck+qDspzuTAsmLCv+
AfGSZcXa+dufukdoZ83NYNh88EArPftlJrt62sWLf8slmPMwo0AMOia7h6BWGpPr
UY7XANKP+qNU1rLh1HhgOOZIIICUHVbnPpTw7PegdNJ8VPDUsBFECedJgg6twKuR
smzuqGQhGpSXZWLzhG4gvB5bwxejsSj7eKSPXUyPziXky+Dzfgz7jBZ0xxDRcyfQ
6jU0lXRSMRBjjqKGEy9eQ0x1dR4+GZJPZcRwkuQ+knxmmD13p5zAeYobQplFzppL
jZELGHC4RZdJkQJYSekEQ6/8xkbObO8pWv7vsclX+t1z5PAXz7GZRDpaMhC5z8eO
4tmUJltLTxxBZvjthBRloHdOktwiH0yjaJLW+G34segULFjlUnfuFq7hZ0cXy3vh
R8+OSq+vbhMZxAWBwfUXZxOoqfvsQqBsmUF8GhtoB1oew8lwnx/MPPWW/69kelsU
hSOVFiY1+R5GQtkXsjXI3VhKn5IBJ0bKL2yxhPoVAU1hEoLncEAaeQ+mwxvjgJ6+
S3imQ3NsiPm+35PVAS3N5FHlXpAF3fAhpTXxSUn6CfbUFpmCBk7Bx2x+1Gxvjs8N
e8wsj69ITWlbCWz+yQczoDowB66HqlYR6GtzVSEXULlTorQxYGZPKbaudqizb//g
vvCE0SYe0YA6nQsyZbNBueja9jzf4Gix/FtPu9yly1qi8agwUrgJsURo4cJh1ErI
NC99hrmh6IB0caA1/5gASoERGRQWO7cP8SGtBuqY3KicfsoGCjIJ/VSgPPcw14xK
tcBPwD27Pm+CZ03L0QBzG1EQ/PKX25VgxPSTMVKFuWyeQPt+I0nZwjXqNRZSXZNC
vs0aNZSN3nwArFWxKamkmA==
`protect END_PROTECTED
