`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M5170W+J+A1TkC5CryoGRtNxmQNX6AQe61+zI9piON8M0L3GmySrC3TOsYNBxMF+
7QnB3/0B3lviZj1Q0PJkv3PydFn5ovTDuHuEbeZrjTaEj+dmakB30CYc56I4Ffnp
yc6Q0HS+UcrlCTwFtrg0iivmCO8RO7cHLNwxTqe+5Yzudm0LoGe75QTBavYSEyzw
f8iKqo5Ye7Se9roLySjHfJtWQaM47Dy1gnAZUmCbYJFLsp6xx9SE2zu0BnZ/mV3Q
oKRBSXjokPj9Yql0B+STpadGRZyuFMVkT9hxO407Gfn/C9Dh+nbnuCrxcx0cYNiH
45yufG5ZqFyCrV211BoLpJFgbZLbYtsCH5lyere6ZESoMBpIhLPur82pzO0AoiNh
IRD3u2QgQ4Y1SuD4sLUd5F63GGVkEuRgVuvWpmQKuxSTIn2Z73K8D3icgX6s4ziX
yC8Flw3GKCPHPpXssYgI3ZyE67p+oJ4A1ZYF2wQ3eQA=
`protect END_PROTECTED
