`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gXc7rc1RYOO5ANwvFEwHU5DkXBIHl6sQQFC2fKF+W9POm0UNXfXMGN+YECbCMEHF
h+WWpf22CBiRueX19h4m/xbH3hRPzZ3AzUNumK3TmZdyk4Ti5Y30cZdXwABz87I+
OvNCF12QlEUJbwNnzyYqqEx0EN9Qu7nbhLtLtu2OPCd58g+t0H+zRrrdZsFrA/h5
zu2wwScRUCnr8lB1KvQelDuIlYARZCFUd2oLenk8OJuWsusqkCENWGtjRrGW+Aws
19KxMU23qCioGDCB7LQbKL6uJ1v27fsHDXA5j0QIsJbQmyEQ5p95L8Hwq1bxfS3c
3nhhfMJdWGrLdRA97B8K8thA/LZDm9nC8UG+wPOkVaUt4zpRUGSA3orzGEz3vJt9
kY4lYiY1A6hiJudco0wipTzi64yjjd44oaW2Uji3FBBgTHNjsF7XGbjKcPLw7cBd
yLW9haOcyPs6mbR3bf/5ZobyMtNAZwCWDInZh2sBUJTef2asRLZ7IltdH5ogQg+d
/T2gmscskIS+rdSOxsjJ0u/Y+QceovcAD3qOgmLb9ZT2FuFjB2Lbq0oDWGZZqVr3
p7BpjIr84CX4M4G0ev12wH2+ECUqsIeHit/LeO/zsosI9jMyeglU7PF/TffEg/1x
QxRIZuJLP0o8p2b7ryCiWGqpOQ03KixM3Qw7X4D1Z5M0yyJvnPFzWvXrnV65W7xc
Y2phyAWpuf4vlwg7nkadXfi5sQao6h2805WBieKl3f+Ob2Mrf+ZeZ0qF6cHpB4g0
pyCAGyaxbyuYjzsfp6upjxkcglcnaO0pyXtPc6Wmu7lecZG9uTy0IAcZEmeeZSUX
/USpTWJuZHMCFZhrXZc6F/bKDsj4mmX8ughXE+fq4Wiraj/bOaN13fgw2syButfV
J8HbjS3BgC5dyS+iexxwD7ZrQx/D4YrS98FPWSj69Kz8Ajl/1leU++AwgPYGIsBg
vW5w/cAXJ5HhOHx3WY7rivpMO3YR284b9ZY0zhTTHfAz5kthrnfEWB2bMpWrY2aW
HF/ieplkSArmwCKNv1oZ3Jz8RYWd5z1w1UqDTCivHaxgXc1FpPbOMejBQLEpNXKL
HAc/eNTtZhHlEK+yEsRZmCEO478uLlPW/dKv7FaWneqbJ90Jp6619jP2Qn0toJrZ
8+Di5zUpZRVVI13d7iLuHMSnGQLET72xybnOEJiArqtuZiM+zMTWlongbIGy7z+K
/YhONN46FLwJp2dVdwhJmCLE9PYNcHsZu4l7CO+DptB7sLAOaVbjP+j46c8nf88x
wqzYG0AUshz3vH0jm+cJJt3bfEAhfCqbNWCqJOZ+V0CYydASFIYwoOpdUGVShY+f
WMciTg2bWRZumOLT/t2ECf0elA4wbSLIW6uckzVP7e+jusx0KfeNwJGXXB+tsA2/
LApRJBCf4zgBo6tbucOZUBLA+ICcyRiF/LJnyeS6vj5rk91KMQbbIaDvJnM0ubrs
EbbSGCNQZRsPiCWIVej/rEDxTeNlqDNAtDIiwGWMaPH2iZX35D+eAXV9vRjTU1du
76hgLub/UWlkIxfVjklLnIisFA8JulOBoywr2Ti5xtHzXs9h75lGtq2nn9NsSOEo
tSDbNFiOXvbP0n+4Ej3hYTzCtJ6qLHrPKHRE9YqGlvc0EcKWfthLeUFvTT+nd+r/
UuliEz2LKPkDcFAfOgaQQue37MAcTZttIqvM9qAJFSW+avZuW84BrvOESxVUl0Pn
7iArpNIeVXcyP1cJvoRLpA==
`protect END_PROTECTED
