`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QTfDQsi46mU0Ymz9vBbCQP9unubC+4MyNvMR25wENuDQxjiUr0tBonAxjt4w0qZe
qkjHdA8FSZ9Yrsw0zUfptOQPswih08C+PriClPwwa+9g3KbmuhPMb4hMlTBrWFFz
LB6P3BDlPuO8+eZr1Imtoc5bPTPjUpAbKA7z0CDk0zEA53ZUPzQRpOwb0XH8/RD9
WggA3h88VwWrwJpH3Y9XAl+eproIL4Q46eD9PwKPOqPB97z8KIFYRNpSLTq21Zut
LfdSwtXPx9JpUzd1xh8iLiWp3WBP+bMWvKU2dJ09XnXCIWQsE8SE4kfSSjeKQhOD
RVfRh886lzmpyTlTJwxcRQ==
`protect END_PROTECTED
