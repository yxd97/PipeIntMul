`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
01OZXbTHu6yS+7AIWsvD0F026AFiZTDE/anHrpio670CkR8QNQuCg4jTTkUmu6Vx
2R1ikw+DU+LMhOr6iQ8C6NSKEOA7BubioJpSZwmJsnyAESjEU7uuqRF5acDbdfGz
mAFJsl9zYXUOJFOu8PkNrS3wtanww4K7TzWfWjHui9zx7UpxKaXphE9CDyM7m8DT
bJEfO+UazB7Rv3Uzxk1DNkq+eJYE6lUr5dOzOo0M4+R5kTa3ZLupYaV9oKpfhwwP
0e1iNfAc6zwTNi+YCOO03dFTfXW5l9w6f+qwppfvVuX11BsPjUM3mObMXd49YJvG
n9suBEjCetqCON2hAW5S4g==
`protect END_PROTECTED
