`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZIpKlFGtrr6aXG0fSPHpfhusMyn0DE9mpRy8jz1sh4r7mDheT1RUc+CyivKwpHr0
7oDPK9H47L7JUB2MhgEXrwG59Jx0bBMOFOb6BYv7XKX0sz/PeGA9Uvf2gGVL4c7a
oXFUX4ZdZRzMvaxKwcf/Rk/MVL1E6jZPVUh4qzPFarpqulZG5ZMIK/NiqijYSXLz
2jWZB5sdEMjgYWg/FDJPpbvadA7/9SFTvyku14gmk3BkPoA3sAEufJrgeyN/W0Zt
qSPcFEi5OttYDACWAZdlgNAB37E3Z1arJJUBb3OOBDZMBOYGIjROClIAxhTnWHTa
Sm7rHrfD1Trm0B/YM2n6yBGWPAw0r+WP3CybQAKkdCQ=
`protect END_PROTECTED
