`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6J/cz72qW4qXcdSFNCCwkqn+a4CSO7kTvSpcEEtJvNfjbrQl4Gb8qObbVxfzN8i1
7Q/egmMmCybQaDYALJOvc787VF5ayVbBSknQPkSyxtvOz/opYLuamdgVhZay9ZFM
oirviP/5bSwUvGzJ5FrucZRxJuUC37ceNe6xCha4cj8KVN9T/FVKssAGXDOI0PgV
WHqSK9eZgSul60X/v7mz8GIldDseptNiG0eFsFQquF/85kkVrBb0ShXO6s78zk75
hwxU5V90TH9zD4Q83tUgOVFqvnspvmcXWpcoXB+I7+D9a2S7XGGXKTyvySzcFSAG
eF2LENf7Swz0uQ4vCUR4SrnoyHSHlec01qWlC7B0O8P7oDLgkZ+XVfwI9PV/bAoO
iKn5kRCvkgD6B5sE2bTOY0hbsv5Cfdh5mxmOj4IWqKM+ISbjDArBkl3/jYPnJsa7
F5NmI/qECNEiV+abHjU3RfIzhIuKb2bZnFdAbF3jQQj/5ebcJqUwoCqTjSiIyRcv
WZvLj/pGxgjHT3MGmiiaNg==
`protect END_PROTECTED
