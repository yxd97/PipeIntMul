`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PHGeveS282O9H+IznR51+e2Gxw28mtoMgrCSsGYTqAZHb31bI+KQpKY7FGHuaVTg
349X4cbu+0/LNsmKyNL2b9KtOW+DBHBcWLWj2EnQuPTwa04vdygIM2HM0bTlTk/4
QzZc+clkPhENsMF+XCyR0tjJ8fzKleevAt5W5K/9JOaE/3sHGQ7kGwjUU7QR8VRW
vyND/5GI5T7abRWqJOeUQg9mpghE5iZdp+hM8vvbTjX7IFLxoLhBbU1f6644BCNU
ijwGZ/Jvjrgd1wXCNzH6u7cOdJoBhqZcb5zVHMxgzUDIdXEMYdFiSqP7hTD86rQV
4IIakUrlcGyW5gstrGZrtApwBj+L9eQUNxb/MC7BHFT6XBw94lLw8T/SbuQ30vqp
cmT1xp5rQVcMA1C62MDX7O2gQ2NQYKW+2yGmSW5EhKqceW303qyWcQ5zYBQ6tSqo
a95/8PAJWjU02Y6OLKbtybIcy/llhl0B9PIwmlmy/67/vb937s9/+Ar51WGohinB
`protect END_PROTECTED
