`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LVOhe7zRmkVQ4ssjWhUeeSbS6YSh0zVUjzCmolznvlYnflfCYf/zJhI+/BhC65pM
GmN47S0mr5HOlaJIHn3r+op4NwexDzSbwXlALVkfl5fZZ/jFEDwgEtH+230cxcrd
Mkko1JCcPm7CmhKbvo+E0jn5YAXok2DTVu5AFJCJLFON5oMYLkfC7Y9yj/fCn41z
VKljv3yHZCUW1MCeRp7oh74lcgQkH8NSyCSjmjD+72dHA4csWvGdiNYyjOXlIFH3
yi5vULyOlw0dg49JvVz3mg==
`protect END_PROTECTED
