`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0xleNuijJwNLPx8T7RQxSSghdgLWAo3K5+j0jwcOtUXYKcAZIds2Be2dxsMR46Zr
YbQaJltfdn3mHdoTYwqIrsdOt4Ertn/9ocOSpzhp8Dw2sgsINO3S0tXVP7dkuOla
wRfXpxp4uefXaVQsR69OeaVuCa3bJCn4f1zqo+QK9XVs9IL8otWx+yki9xv1zOuI
/0wRXcqQao9AZJJqNFWm5qWTduOLahg+bxLA6F+4ljogXPq/wzvmRyR4XGYzoRcG
LHrh+WzOk6KPtCzycfxwv0fddmibKT9B9lAJKiG5kcLOeYblPnrZnpiyTh5f9gH5
a5g5faBVmpW5++9MBuCylOeK9Ns5qi0tspS1+4jk002QA9Q3kd4Zq0CFDaT1c4fX
A1/eGWlMcSvfskAqVfKy+MVfyVaDYC32w/3weFPW22jfMjjWohTNil+n+xDqRqL2
`protect END_PROTECTED
