`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9/Q5GAIiCo9YQs6G0vc3Q6kWKROay57bfpoA5p+X5e/M1raTxrQatm6y831Jz3NQ
jq7t4X0ypXv4UGNcLG6k9pA33UhtZSXOZ1hvnl0E5/QGbTdAZYkgEHW53N4vPevL
CzifZWxz+Ejlt9btE1ntTTRojtFwZqBm0U5DAg+ieCoPjxkqUl5FheQBQBJdkX0K
vyo1evXHEmMZAV50Yqk8FxgXDO1a2J87jiaAafpZgYSjlJmQWaWif2kUCrk41t3A
nVpmqGIdjjptEKv1HPuXeBJQQhQTSV8QVyktnuyUlyNqbztmkSZ5kdckzsxsXp3q
uVxBLcUyzxj+oNSJUhepcjmQ/UJS+I0OGq1g12fss/jmcDjw7eFQvd5JHtjAd86/
2S8n+p1HyRhAl7XRsnLMzr37A7xvMx6l0s234q0edLs=
`protect END_PROTECTED
