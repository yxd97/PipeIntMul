`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3lov7MOZQlB6sZfumigTXeJ5KbFNbDdJUCBrdGdAfS/OmBKJTJaemJF8feuiCMbj
qYc+FZLPXXI+M4L08IkMLuK5fLRwXHLd40BFYkFi2ls3GR8DRnHLW1710l+TqZre
XSpmhifuYEUhnhJwreS+Y95YW17hesIBOzYPvwcqj2A8UdafuLEqI8miDUL5fSQm
//rVF9v7/ysALeZtYPFZALsmWf2HjrfHyD7Wws1LEI7WNUJsx/Y1W2nzS5++xemi
s7NTtGvt3m1EOYzJD2HPH7maTDlgu+ekffVPFObCazR+qgHzB6eZmtXUMCJOVuN4
ETrg7nPS+wmAf9k49HtJGgc748IITy/xdpWwgmFOcqzZa1G0+ktR6J561NX3m/RN
4OxmbrMn1znPToGLYlewW5TpgOX3doNaDGzqE0k4xUa/mEDtn0g/fhUqbxdEuqoE
`protect END_PROTECTED
