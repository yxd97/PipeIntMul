`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3P3JP131lTCITXAVRWgRE+gzyHuyykHiYlMb81SMogBHdl6RTUxovJKShdBcjKUo
m/ccVFTfv6mjTk5c+H34cSqKGBtj7iLwt4rUsLRupbv2RXY7Py7L1G5cl2pCFjQA
AnayZRCk3rIEcWxwTzL6UU9AgHQIiycCWkfJow5N2OSQ7SSL2HPuD9VmuD1/RAMZ
dSKr/+wfaOwvff1aRFVyWxqZtgTy+RClsXO8dQzn+kgvw9v5nwQWXlJAIjyT0k1Z
29lzdfbjQseL4Lklr/ZE4EpJ/9ev/ywdud+9Ke/4peR2Jx32NqbE8rvdNcj0dZoH
EdM7MRvBxJz77qNUCrdk6fP8gtsri7ejjXspjMV3pqH8ivakJJuPC7no7WRi52P8
cq8krnwXTFuowjgrbegps9CQVHIppqYJmubCT2pl2T0i1g37IhqRmtoMeS++Zh6Q
m4xg0SkSQz5fPnHtBb3nikGzLQHmDk477XvH6oYc0XQFxWvahqSftdE5PK8QX28A
TuBq7k9CuEyeJTSOLWyIiA9eq+3qx3sI740+dExy1r4QQnSIHdoIgyi1SNbl47Q9
L4O22vNJs7smREmqroCwl0TrkI9OzX7EEG/NobO9ei0SAI5sPcfDP1/OmbpJZy6k
KGVllJQKI3mpSi+3j6dlOOgIMZUTunfo/FlY0V8IAjtPRe3pnBd0DPHB2awVBfHu
vw2g4wcWz+gkD4ZYZa3X/IV301Bbl+RnfcVqruQGbN9eWC/2i3FbkC567jIqTp2e
BmAfrslwq6sXcJlGuX7k5hxDbq+9Su9vebNruPFtYARrcfCCMt13WRs2UuHkOgho
CrfSeGaf2yclSzCrz+iKT79Nu3msJIhgu78k/3RE6YqbEobqHCDyVVmhZBAFJoEb
yeSI7uwAX3EIdVLaIE2t5z2/vUCyIStXcfJafaK4veSmbZuFNjOSQuALTMVZOu1v
ymYSDGL/jGIcOh94oS5gjZ1FHrxbYg1+zAIBry2Dkm9X6ttC+aI1/thdA73yRpe9
XcCVbUzewwXOZgYJYCxyJVl8SgX2DuhWFOYXcc7wNEQyuWwrwQ/d0nbOwDneTeCB
86pNTkzm0d560+2u44I3f8F55gJeWKCwoHvLQ6tmKeTb3uZauPaSPwSYa++Nqsew
evlVoUGveleiTzFP8l4t9eXSIPO0GxjfT39t/yO2swm1xupxvMi5wRLxnFAHifxq
if1AenVtkCArRYrveHR14lqvI+/6EKkOrmzFM18caio=
`protect END_PROTECTED
