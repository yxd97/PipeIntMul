`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HE0e/L5wYGN+5LrqLTNZNfSQvpjqMhNwbfNd8vxKNFLSbFI8tpLzogwXXfDY4PN4
vRy7O03Xjp+c2GuZZBJYEboGR+/A97Pa3c6yJyaV24uhGjAwijK2BdNuC6s++pEU
Jpr3fZPC3+cy/MdO2z5hZgmNpnDRNz12r9NQpt9W+JjEMKOepriQmVZsLo+ZaME8
pURkCFRlOtb3McC65N2zAZJASCPpmq6w0juTJtHkWbmdBLYVZVhH23TDzRmoe4eM
HsmO5Jq9L7Ih7QmZzNMYYBCKy5YTyAiSXSHeSiOmRKDufVPtkl1ZsbKS3BSqTNZm
LDnFuEHKO9nq/eqPIpEVixkdwsNRQJ7zFqRD+mmRcNVDtkDJHroHL35N0F9pZT9Z
cU67fJEvydfImDVlPF3eJWOHO2ONojs7ogjb73EPB/eZI/D08NSU+zhXBdueagBu
cmPJxEypeyKMmlQiTQC/3uZx8dT0M0rihVSjmsir2II=
`protect END_PROTECTED
