`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6H+WHRU2u6vKDfgMytYE04Q0IJWYdt/N3TvPNc9PL/xGQMyusJ1w+hY6Zl5RRlQm
6lZGsimjXqUEjZYuZ3K1sN367X692xz1uZNU0jSzJsRq+UrFG8xxNjMUkhQvUq0x
8eAIbrRDYuKzHBZVPIOHPAFON/6oj72KuGfg9yeGoYwjmfvivN60UTc6lYyScjjY
/3rXCebKqcQlcbJBoTV7WjVZ+X2Jittr6v9jdRkvCVcWUoUk5QYhzoOS9EyoQkMJ
0ojubo52CaHm9MV1ZqPFAsuNF1egPG/I808qnUsdmq3KAUwgUcS9HOvxOtq/ZMnh
897i0cCvnlgOV1jen1zHSKTYEtK/XmpiAGe61IELiZk4BK9mCtnxDwOpxdYcjfYp
eTf51v6utGo2fIjlmVwEt0zPer/Zl2qMKwQJ39TFe9oGMRpE81fth6tbORsAgUOF
af9Mo+YkkDkvxd5I4dnEW2LJuHhrMhZLYm0dbmuFhi6fZQIhX82XYLK+ooejmOz2
LBjozhrbvQ4pyVGhui8jW/ZqFt6EOPwG48FuGiDX4xpZ3pz0c8TgA5wuX6CcaKIV
1F3x7B7OBBL+l8kFvCzlSrqFRJ3GJAihhZssMpSeq/O21egt7jOTRNU4ybcfo7nt
PidwCmSz64jzqOLbjG1+G0QqF09JMbphnVOBmwtu9VHmYGIEz12iF6tYwCzQLOT8
WBzOFyeAphn4NLEc1EkvYrnFnl2p+RQn48tSR6Cbl7BHQbbv/J9UfAnkt5EH0N6r
cjYkRUHXYoyaLD26ZnTjexveaoAkUACNeSMCy39N/LKxXoxb8lhpqZosrMtHdSs2
aXTHzSkDr1y2/da4mAFgk09niVxNZLi8f0Qrsh6Xezea/PdhNewOUgpsCf3tNUJE
f9vHliYva47K/m1/y6S31kvjxC+S1Qfqe034tTAZYHgnAFynV9tXH/YlbQDP6jK5
9Eihhs0AGiqaT9Hyr4M8vozRr8HLe4IFYX+n+V/H2UMK9DyureeP49k3pH667Ujb
rW/yeSZcopnP5FGdX9pgbnXxWXTmi4RUAJToQNzhCWiQWOJMTFRjXhj8cSFCdQ1i
EfcLqn8g2Pw1RK6DqhyFk4z0zA2Fv2w/FYlOLDbNCgxbLV0djK2fMHQLP9IQ6Ci4
ZBlQ4DDcXTsv7WwsR8fedEBLgzgrxXST3FDcHpo6pS2SP01vA2UtjAzVkxudzRQ9
F42t/mvWI/mKnmWs8OIxOSfv0jnRL38HXWh0/+geOR153CgqR0lXsWwict2VdP/d
FqeO02rh3GAKbJ/FDD4QHf++wU5nzVtwIQpR+4BD8xkWSEpWF9BhEbg4G57rdr6S
HrpEsbX6wHs8XyChg7659bFH6aQqQNCYQywBZI1hHF99+qmpwC/xGX521xZalFq7
cJSWjIM1I4REQ4tTOTxBg66aVe9HTGJcMcNQafZwaPIXN008YnbIphCx8SA2zMXa
fqwBtz8FfW84tRD3EN/+Hf30MFHVSn9LF2r0b3iwCS+kf7pYCzpIdfCi5Of7PP6c
KgL6KBfAIEWJMBRPlIt1StTCQjJuTcjWav53fPH/hT54TQLhNyp0SLkL3seylAfp
2oO92k79kUJ6wPH3pYiG4HWZTugIw5GzZ9sBuA4FKxo/j8wNRCEt6p/133FBLXoq
KF1d9S5heelXWlLT/ISlA8Qai8iQxeFAu+wTyFsS9zSgBIP/8g8qlauSPO7kY5ml
i1uSfmTYNpL3CRAY21d/IfSzPxGOerrbd41mEOpZn5SOfD7eu6nZzfslS5anjsm9
74V3KlpGBETZU8zOp+z+EKTApAbPdccj62hwb09+sH3zxvcd+FijHkx4/oFgUHlw
6bMn4uEBSDMCE6PdsL2NjSJJjZVrASbcelgY9anNaeOSa3thx8EYvOXob5VG1tA/
+wwJFWenPBC6tgHJoe0rsug0q5YYWIBCfd0CQtDoKhuDvUjeZAH8f2OK8I+E1Y6O
DDqz53LD1ZyDX0U+KvqaqaWj7yY+wXSmeZKLpBowHiWFdxrzwBmQTN5AQ1/RGc57
ANtHwdUhYGE9p9k838jJ5I2D+2dpiaq/mD++J52DCCTa7h9LAxisJ+qHwwjSoufd
L4ToHP4JU3dZhZ433x21k8yJ6TgoO2Hoc6fgG/pzGzDwucnOFNAoi9UhcY/LS214
fHPU0X+CuHMWt7lsSuF2jsmWHYOVtebCWLf39IFski1bC1+x4brz65an5DMzmgoW
p8HykDonnULwFQwdUSAFFH5GNiEYtHosOHzW2K8K+ULtIJd+eyXee66Jxzj1yIrZ
08gKYprUa/Evv1K4xMyzn+smAcaff8Y0NojkPb8UypXk5Ihc0F3JT6fGhWGVl3mj
+kNLOOSm3d0BRqm0/JFE1k/5IhZ9DWyCAf0GPRSJeySJEDYyEBqQ5GallOjg1u4G
3RtBEoWhRm4OvzudqG7EsiNEdXmZkzbY/45hAQ2BN0ySvq20nTj88CNkKEK//FGd
OXWGD3D0IgK5qyxLWlBkNg759FSpzmlqYjGMfc0Ncvso4cc1Z0rJZVyR4C1RoIw0
N6pslZybarSXWb6ljhS6nUDbu12vaFDXnizQZABeYApWTr3NsVi3F/zTX3wtrHV6
4t+DGIK+FwnG00dRdS/hpwrrEaCOuOqu88TnEq+wNmw=
`protect END_PROTECTED
