`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lq2veEXtqd9LQSPTkO1QJAdlZ6MZ+qjXG2wyaG802YjmYHo+FE2UYvttOmPfpRYL
K9GpuLYyiVnJs2VhSfgFm/u6tzJfTU4zvoKYd8oMP9Ty1Sb0M35RtK3jVuZGeaiO
3obHtifRezQ4A6r5pjRRSzsqBgXSNW87bu1W0yltDk1QBMHLL76RBXgyBTfOw7ZR
4vRLRGC4PKe/QuE8Q/r/cu3ITqeR20JmJfqLOzVGR4a2wcB0vAC1uJp3kda7fTOJ
qMUJtViUjSFL5YA9Hj8BzX0kgS+G3z1wDk45h46QZH6YKHV4xt14xqWwNE+6C6Q5
XedCaWMHMYIDyNQJozj9TWEpEJ2EmK6z9CpX1E4/7R6HcuXjnGocyvX8xtCzr7Yx
d61MgQMD+wmtdZU6Dp9oiVPPVu3ucPkiZUD6WdSjcMZREuiH/57hrM0/0uOH56Oi
zDI2nfuZBd3na9hJ8x/Q+D4bfzDjsdRjrgFN+1G5bNdbI2wm34Bcl9RcJIuc9d62
uZ5FzIahjcUr1MX702on6kZsN8X+qwAtv1BxoP2rqnVRlhHEWklqoCLELFsO6Ei4
eJYsdlz817+bxcQ3yc0GlwUWcC983FOcmLhr5X8TgxdYi5AQbSpYnfBRKu6qx7wx
4WDtBYxCYTC8lM4ZJBDUJLZQfG0D4sKRkynBv6dLhx+Po/ggU2Ld/2rO7yzgQARA
bCopa5Tqdc1kIZZ+tbCZ7RJWocaq3tl1WFZLMMmLuc3KagxxMrlX++MZTuSxwG7p
onckDAO7NfJJkE/cwiMOOcjIygDj+gReAK3aHmg785qrWkqbigT7X3ED4riAoI7V
yNJ+ab7M5gLa/wozb8WGGenFF52ZktDMKVx4t3a7DA2on82d+mXcxyt459uIBF/n
AOxVKQDZAYzMybwH7nM5mT2V4uH1mBSL3o1xZdsRmZJJDfkonQ6aJZY5NM1Aytcb
Zt0wK2g1GhzhOkxY4b7X1I8nsXfrBJ7CWn0ZuHzLrx9vtBG8wNfO7J5z9bvPznKh
76rGJoIOq6LIcR+hC8otLGko8TbuxK9UNz2AuE79WxqRAw8AslsKV+MyPS1N5sZu
XaCB3qQxkV1u2SqHoTZnem532MPUf/IY6amk0anrbIYfmnHIElUBbks2eLPR8D88
394BikHrZclJUgPVFV1UGNOlKGQml9HgtkFBoqr5TbP2PfCWz9quIY7PQwZc+C/x
NcvxuZfAG2mrV11Q0YDvOJpewsRFTQOwSusRJdfyXsNnWVF5ODoCETQx2uN1wtlP
`protect END_PROTECTED
