`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G7neGtFKIpW8i1WyLwehuNVjbpD7O1oxBWhfCv3sTnqWsNk5XqektKTNw3oTqsNA
PzHkO4e9qFXJ/mg0FZv4lNyIJqLdrStkF38BOdoWKHFmAiVpQ3y9QqFWxISR7zS/
jR/W7w3bIEvcOV0C1kmJph9zZSjBYOZmnLF8zZ8DmVgUwO0jwdXd4HqZuzc4rCN+
ZO3dSBsNM7BUVat862JXgWpTPLX02xc1fQ5xENZpTm3Q0deCc8AWuH8QNdzxz8JG
0U1/nkfOcYZKpLNrZeyuqUdLYYhwSfg9J2hMw7agSn+qM47JZ3LHcWxR1lpZ0yt1
8ALHIyOlBspKOSUkyOQ+AKpEtj0vgtXm/6KSKzvvlQCxYDFkJ4ER3Pdep/Qw/XUN
YaKbOK2WES+/wG1AHeu04PT2JyAvGHf1jBitjaeYFbgYLlCfS3C7K6XSRsEO+n3B
Qoog0htiA76ZczZ7fmHHeZgHACWN3qYN1zW7v8muDErTyRxB/pnT4+Zcwub3MuAZ
KLDnb48ZX1MFRNWTC2bu3pE0Dj+sO53F8G9CfSpA7QCWdW1MnbPEVD/a7wtYDHYt
aS+sXLrGGZkIYtH1Qlml2VfZhADp653q7vvPMoz7z55rDLiNEt7L5W44yX3M1736
UIkBFsi6MmQAKU0PulZ6lC6eVNLJ/8htjl062c5drjN35d2rPdXgD16bFHP0fwEz
T/jnKiC7NyQn6rySzp+AQmyJQV8s1Vx2yy0fyza+qBKDGBnCbxRzsoGpADuOu1Wl
0yvR/bjpTau49ylJMNZ2ltwXxUbKdaF3mjGDmJJcsuB/69wxHpYM0LxtreQTD3Kl
Ww6vJTckYKw+tzjVLdz8PWX/cFbzh/yrGf26SQDFmDQI3dsK+GF5PTQlh7DRHCSO
3/ION/xB6NhUmmxIjzT3zgJhHhlZCypwsWyjUSr7Iom9cl8CndQUIABHVQM1om27
gLFxAotW4Kg/mtOGeL38O+Vfu/ktyQ35GmRV3Qsn79HPVMH9SWf2FN2YtCNMNXw9
QiTxThBQTn3ArC5WDrgsz19wZm+wPgl85uaCV5AR5Q2/pfYfCkKZH3rCXPNTp0yh
KLLYPPk4KuJEdN9ReBfiube0ylQfTZZgp1Tru8/oaY358OeGdDpap5Cb3a+Zz4KJ
xUqFVJREj7JzyYGaYUsO960JRO/mTMCIfPw/yMYGhdJmcUwEFXv9LSJqEm1hq8kK
LCaxLQnimu6raBnBCfg67qQQfQu6E3+8ATdlfgy+IlQstWyQ/GZLGfwzNgOq2WzY
gkrg8O8ybbG+AYOjWPLBpsH6YIIDuxIFJUBuoV4cLGCj6QpRpSpYyEmpVundJgZx
buz2t20JMzwHt9rcWlfxMV60NfvUZYXxd1p8+hDCjzUWypNnZ6JTILPb2FLpY5Xw
M3Lf5dh7LQIWi8WWBYNGa2iTVAJ9iKgPOc1KUEazGfaoxy+l1uUw8UWHo1u5QasB
KoGuQ5SXfIWkyEdHrc2PxrxXDYatqZt7QiBiNoTwbg+hoLJpWWbAp6yKtq9V1Oi2
E0OAcbxvHm1GpgSjs5LtE5/6hcyZ0QFbAiQa1p3Mr6Tbr0CSAWV3y1v15yp9d1My
x3s7So+nERsb5G2Yr2SGqpZlwLi4fumFB6dhOss5VQuABJ8cjNZPBx89kWULGQ4z
Oqecu9VTer8fK1mo554mG4KQdkgMH7Zk3Kq3lyZONJ+RJ/re4FL6jiskkC3wiqgJ
7VM9vijuw8dWgWFplFfI5AW5osbGUvkyFnva4ilJTahY9K0RachaD3snEKOK34YI
Y3yYDXTa1FS7aqGZ41Rh4ulV650YWLwLLH/6qw0btdawFK3s3WnvylwZRTSGPUHe
Wgt21uv4IPM0qrARovliQzmeZXD56nItnk0i292dnvB04FnRbvVW/91Msdxes/JJ
/RcNRh61U5NRRY6g7j21GfGryFZkWojkzZ4tLcxPTiQfNHsMy3M92CyjS8NbLHvA
U5utDxMUbuOiZSbEDiREWLf/R+SJIJQ1gv7a272Eb06dkzTJr9Tt/B1e1IBofiuU
G8C8pYhiP6Ye6wTg+ziWVNnkNrXK8Z83stjOCha28ubi6Ffdc6N/r95LboB0mb4B
IwqcYXjghh35+hHgFQHWwPw4cD/DkEibIf3nwuvAZBtIBIfoTHmzurR5ZEhaR07M
DDMKXeb705TqfQXHVTkVX+x59TcBz/KzTogSReBYQHMyhkTu/nU94tizkl9O5OJr
OOBu/jA5Bk6o7UPTGxYTrE4U0kkfcsiWF1b5jLQL9Glk/Zax2RTbcihi26kJxJ47
lx6M9O2WvjiLOrcyUhoxUTuiwOFMXLzLZZWfv1MXs+ODms16FGx0zh7GC7FIt9vd
flgnnDNbU9s++niEC9N8dcUVcbpm7U+kt5Dfk4qXAvjxTLOUihnCEwUOcK00jgwJ
yGWhqxiQ0uXS50Z0T6jZ8uVphW5PXQcGMjAwhDWcsYHZHKDggWQTPS/7HxcpTCPH
SlIv9UKwhgoxprKrr1oc9pqhTtIPz1b5+3gpTZ83kidzQbDdZNg3wmzV/JhINczW
r0f/uxuw1rVkzzCE5P6229qUUcwnf1Q5GHrBFWUutnOwp1TnAEQlmCp142GbUpig
gcHkBjmuXy/p+cCgMevyD+/SoJPWgXWm3i0Fbvs+keoQXEly00XhXzfeCK/XcLnY
Oc53HEH6i5oNTWUWb4k27UbioNRbGrtGrXnEznaJV08/G/zWxdC8BM0fHYrPgIvs
tg/5BcYhVZdeQnoURUObzksuNwRYObs8DohHQ+BEvjQMCXUQzIEIOkn9r8k2mjuD
55xwZuk+Ic9wZOEyK+RtDiV0g45E7tZ6vVplUrewkQ48j6EriS/3mWcBMeHur9/r
82E5pOHUuHuWA8nz89ZfXpUxGP/YjgNK7Q/1LUSiN8cO2tFEeNcr++6vLSjvzmMC
vyspQth4OkN6rqAPK+A2V3k4hO8RIEIh9YbSWGCc4GWWy0z2nWkPwKqw/Ha62AFI
u7QmPTtVf73ysimEC0o12BZhSXQYo7oiqcmGTDO44+rNN2MU5Bpz6QU+VEw6XrdG
e/R+9s/LSrn9Wc5znTCclah/NOynmvdtD7iQ583Zqlqotvis1arQTc7IewIwaxqF
AmmlZPcbk6AZb+8YkJahBtqwsLe03mD2yFuzzuJA75RBiSP4Y5m6/wWw/9PD0Dwn
i3/q4OkptvbodMzDx7SbKQKOv/pzNbk+gGtIIa2PzDkUZKGll/DJNKoWYswe3tQx
Z0ERee7I5NyireCYobF0vdxosFl/wy916R7T04U/Rc5TM7uRDd4u3ytczGMuDgOZ
Guzh6kmCmfao15nXJ1+7ii06a8D5MCQimc28vKBRaiGQOQJy09/dn7iMZ62uEsfE
fCZ+rfBg4wO0GN5U8TLk76zsLHEUedmIachGUD2EOsDfuP34JVilxsI+OxQQDDPw
HDu8jpJ+CBlnAZczCueyO58C1QgwJYgIrpqFHdMQtbm9VRssWuSeQ7WGnFiLcWMf
VMpQQWu+IT+2YR1AI1/nK/ZrHlX7oqpHSR6I/QQEcjuRNAZ/omXncgHQYfcNm+Us
ERPdPmK9g2FRVVqta01LmYwWjbH0VChncv6Z4Fr9nVGoiDNjF1KckK3JdKrG+/Sn
3UBOf9xsxuxqOp6hWhxCnS6Uj0UYLLOgHEPTwAO5anuOjTODToOHVSe8CfIKWc68
u1CzaZl2ZKs+BnSs4XlHkuuaFevhxltaDekD8ShvvyQ8swFtSEsirQh9hFLKDbBM
w5tfYYGBTGZ7o4URaR/N/jpvkOZ+wlxkgjRvxUwbhH/gtWz58HhpsknvS+fbuHFd
rkHrZ4edt19rjut624n459vFOGayf6bMSe70dnXl7bINHRsuQs+B37ZG7KqhN59Z
0UVrAPsubdFMXw49p1dY7uUSCNAS1FXKFBvu9W/Hg4JHDdIjEzPCvrXe5iSV7SbE
0mOq59pSRo3QzVTDUu9QVstHrRKBs//LqUtinqsLnyXS7hEROOSiFt/JWHk4tPPo
UWkUslpJcuI1RwMgG2oCzyrKPIUrOAk+LdJciyURcyloFxzb5QQP1dIL9OHO/Dk6
zYljJcDTC9TS8964VuIihgfteR5br+AppBtQlIC1bAH/lJbAxMo7s4IChJOBFurn
Wy3BOtuNd5amtaPmushfMn6vjokPPQnEkE57krfwNK3KAlFQbevcXV60gsuBOETf
jJy4zUHZy8znKgz4/5DcQ0B+i8uURbXDqwI2imIdn4I85kgh1vuPpZdyDhZ7/AET
IXrR6I6pIiyVrjJrr5RQTGaZPts1i1wFW2q3JbLWwqYs702aX7I4a3RUOYrRtGOZ
6HkcylCzonnKEfr7QBP1S2CSGCHqcXwzQnDq/1/LtYz8gU1e2DMHDGgy/SoG5fNs
Cq+LIRThNNHJYI41e8ra3XNAKicBIn5EDz0kO+xQ+1nZ3L60ksYfrRTKtMCxL/gS
79YbLuadytDhCx9TGzkzAYmLv6OsQF7OmljLt/MddpK8NUaJipzHN3cTYiD68rgM
DNsFQ973V6HOaePQVVTerD/6aP1mqVhhBj3n4hVzzlI//PFUOgLByiXyKmTMr09H
HFPJPIPIvrdu4Gq6y5nNjTkT9co+28Fp+tlePXg+6zh+fyz/X5uowSTItZry18FZ
gE/YP8q4BAVrxgDw8h0RQjGnkb+udpNMkwNYQkfgTIhkOqeQPV8ZAIgZ7/YYesBx
J0GDxq7lxXuBHznQIGhg90pF/XMX6JpBEEe5M1Oy0su0PwdeuSWKLzdwiui3AEmH
YwTvtEJHZY338TpMwyfTRgF82xpji02SnqcBrp8KycZIiqnLpZziQ61bVx7VFZFD
s7VoaJ0qX7u1Uwvdhb5GLSKxlnmOF+zzSYkelTp9e9l3mXAhy6D/vEfyOTlLZi1E
5PyVBz7aajg5FRkW6tjb5kp+jpBTtSa6JDSK7OCmSciuX3v22RDOW669PB31va/+
pOA+SvFYfZLPw/FNMENmw/P7CIculKbwOAQDnE3TTs4Bi+eUYA39VCoxQ+Q+HDmX
Y9xMyEANdBU9Rsc/qwwJiZg+ml5cS+PlvkVa6UBdzJ9cBYBRkHa4dvUuuSUwU0ac
PjfWUuFFdj8D/JCv4+pDFj1jGVK36eOkI9vQ3SDAlG7L9Pd6w/Snk+JZlyoMo438
LKEb07TEDLkNZGxN29te6QbikYCNDP5O2HJygRKFeWwzPdDrkvp12AR6QB7gXhuH
VmAkNMxMlYjDtonX5Z0ovVsq0DRB9enPK4/mCSB9b1JoOBOrz1VV5Z/rCCSaG9Hz
PINCvNRQZ7nN/gqEXogY410tet5b78xPT9CkHUtpEcUrvbrJ61XkH71pCnho584M
pflegn8aRjZqIDsfBcxIddQuhL4m2/o9asvYfXFtVwWTh82bxSv03bIo3GvWPmAE
QWL1EXtNH35/OLDbNo9BFW6gyWwJYoBOv9VVYFuzxhmrGmmvLT4IX13EkCQPvz93
N0BsNQ+MbT69YBgNiM2VY3mx07HuiQNue0F7YL+GNK9wvUKPVxFEJTTMVtJiO20T
LshkpZ32f22VdA1PrSCllkgqhX2cuzFuEkZzxbVYS49NtGvJetQW8Y3O+SmDNuRF
KiI02jywFIl9RJ6k62Pjm5k5e6ScfoNB/Ldb3rxGuEtC32qRkPnAgBfy/uKT/Qqw
CZKR86Mzc5mehL2nP/XG6fnF12k9nVlQX0rd6XN5Y9tmpqePEBdnndYktogSD6NV
kILaHM7LVPccfPDfe4FCkvbbZj4zCqyeHg+7fz5uCVPy01nTODy3jgbOHr3aFhjk
gy8NsCJ9hc6g6q8C1qdy0WaC62SEWTBhEu5W4T7O2Yz/xV7y3emYWRDba7xFKrST
nAnt8f9acJR0dyXywlhdFu/iLyq8fwhPGin02073fofOrzpSLyYb1GuQ5iNWw9hF
1ux5WuDiYORbBKlOEszr0g/FUshBf/VAiyT5WIM5GDEG5sKG5+8+tRH7+M/Crgro
Ukysi2ufzaTwtXTsqotXWqGw1m/hag9BBHsvQx/c/AyILj/r2TZphcYJ6qyFrJ1U
8IZdiOrK9qiq+H0n3Z26uJjn5a2b9sOaMy3KgXzQhCpyF/Jm7eXVGuEleqZOlA5H
b3Yy0x2ogWtVfi4lDNAhSNyAVB9GLIIkXDHz8s+qzZQeiCV8nmLGl5UlQfYHmSes
DqftMoPlS79zFU+VqhnYPqTZTG7db91VOE+p/cQ3L1rW6VM7RjTfQq6sZYvSRWw8
N0PJ1/3JWdVzpitjjb+Rn5xUIfy36YU2qVKofrGdsClw843+1d8FWD4TaT6B3RmD
FdP19p+FFMTbNAPRJOfku1hDaG9yeLCh7HxMn5LIoC2kyVP0G0CIvUTyslqYCZCq
1VqUoXhaXECVCBZ6flYcAENc2z/oEe0sviSC+n8Pw7akLLHPemU4J13Rg9Wzzuct
RpQrwbpsG6x4EbEZnijy6XPgSvr6T/gqSY9+SMBMbiRLb7ONYxhza9+9JFJZ7Q1d
W+/HpPZcEtm0+rcOKZyBgHpoA3/V18zyNf8vinFdBHyWj0P5+YCG4QkoWVzLx6eI
sr3ZFvBFJ1k0Hd/VBtT57OFEMNAiluNFLqKzkgU7SpPLrMS/idgSpN9xUgHvRIAD
hwKNRwej7lplQiz4K8giDqAnuDRWi6p2z9CTGizBqhV3R0UAde4gKSTSFL1peqbk
7l+djTkD7P6TnGxvUByjwjrdlBfe0A3//GE4lz7kcEY1V4d/Ve7jR/2s0WdgFteJ
80bby4sLN8f3VjfSZDmbYcBDq2Im0BG6GLCATg00rSFhgkZ7lJc/InCbMh0G0b/Z
q1oKiRMNBpLNP6tK/JIZnQaph35XlPvZw5+bXFi9U/0E8V5QLI7a20tKk+ry9NsH
hWP+ytcUabtsVg5WLho9nRzVWwry1AW2RTB586GtUnNU4rIuOjJKZ5kttR3NMzQO
rs5/DCcjhUtKJ0qgU049Hm60ow/4QxCYWjvt8LCWlfmI5SEWiqcPQ/AbX/yAKMaU
4BOFs8EmlM6cFH4lqE5W9pEIqYNHaRWPZkg8Ou7Utg/IVdrjzpfVI1qxZB+h9vuN
IYgzaOB5seGOM4gmsoBH2aN0kgiRT1laogyTR0Mv4gBVwXyprHzlMNoh+8Hc3yM7
3sXRuEEdGLWu37JHQ7zWlxtRfiChA8pUNYoAZ0ZHkkrNkAncO2sJP3XEQaK0ncnq
v19IrGLG45wc6jeP93XvKGZfcWojxGzI0CyGRUPL396abGAaP9RW6nf5gEOaU5mm
Ocdxx0RgUQAzEfhMY8hCN1PNtSZTXo1XyKjtmmGXorprypt8WuMqBPpJwAERt1la
9b2oDOEBqyKhl1jle/0O8xqSyDhQMQNm3x+noNEQ7nHLUHpVxrCyQjL6FcNvSrZs
WH8XcRj91H0d38CSpn7AAxZTpkU/OaSfr5D5m30fntKWAS1SDlxYC8Cyyi92YXc6
o6tNTPUq4ySQIniYrgPD4nNnR8enw07Q4jcc+WrNS2JmuiRHi5zNlItlSSD0wZVE
q0PI8zOMOFebnT5K0DAErkjjXsL5hggRyu1aBnLbbh4Q9xUIIEaA88lnipDrs4aQ
j/LDhnMMmm252gY61WX2TIo4NGHP5XfH8WbmX659fdD3kZDoUPHbOfgsDi2BMO1Y
bc3u/m/rmU23dMVHmESnptmD97WI4ISqcTHXRi54a0dZNnjHAMIVNbKFTaI035sR
djnac2kuY4DOVWPGRzMxFNM1fiQqeCn2KqVuECCyiz9bsOvs+AZmIWbaQVHR+ZEr
0vl+rl0cVjeK+Nn/lBGVen9vpcxN3Cn2NfuK9vG+/ukyOTCb5klyVX4dZHRTTV3S
MTr702ZPeunEmhEjwlGvUDB31drtlvIeKDhCv3GceQhQNAv1wT0YCQUe/P8KVfSJ
VvT/lKRNaPpsQOg61jnyNVyxffrs4aKLGtx9ZXTMwADU/CDIKCL9WNafhmguKcmm
djLOGZTqoAYbilcu+bTXKNpErTG55l9k4PvcSW2JofpHa6wAwcix5PIrHltOSmc1
cGTF2tMoqGuBf70u+sE9XmZJvi9Jk4u9DIsashSJCM199V/F3Bgvy5N0cXt4K44F
SczfjMG+8W+wfzQqTBZXojRTLHIKQrb6jrCSPrTFWDqr9Ly0ddUpTohk85gs9EOz
dSOoFuoQ33Ccv9zlxmXGQfMV5vppFRyi3IFzdOHYOIjv4f2bOSJrGJhiv9HxWfR5
gFpwXdTmKZUYwk6dV1WbrlU5i7uzJye4T45c9Z2vzh7zXUN0HzL1Rjosg36oqYyy
hRTs4msNR4q1frKU1jiBg0rz2l/sDRCpiWgzTAr33pWw+DYLY6iWjxLCwAHNgk3k
3+b/giJvXXrZ05DGdt6nH6dV+KRe48M4OS7U0442gOXj3VlLkQA5CK86LX/yURTs
apjYBtR5Y80PLhq1jJXwDij+Y8e7esXmJ4jOy4A3PPW0sfdvIPmd2JPIEXnE3gsn
R/i/VD3C0FR+H3GJGB1cb7l99Dwnsl18hT4PymPnGjxV6nEMUQggEu4VnXrmRQdO
XWfIxN1VfFbd1jklcuaWe2DRI/2HVDvzmOjeIKHtNi5KPmt6KixMuPsSSiAGjDO3
9meQri67FnrTopcxM8126xORefLneUymA+kvksoGVk3INxj0HcGW8AI1aqY5EfoA
cGUdzG3KywA7Jaxyodmsti28ue3M8fB4FVdXGOh1ujGR5N/3hoWaf8ia5cFbTduA
Bo4HWsegP3iMFKpLm9oukjk1/hVnI4IkTNRmNgh14Hc1mldWy2SefT0Utrhi1KNe
a53/QC9NIR33r0B9qgcD1TBo77cyZIbsCEofHxC0+FJtAuC0TrQniC3TOgqkg7KX
y+F1gwlvl3Epw3kVKAWol0zffoH1cLSVnzm+lkdlQK2jLcDA36vJqm32+5q0gZqc
Z8uyJIMB32He9DbILxPwZ+cDjYXTASHLpgx0McBHxXW08MtBGyTWP/QK/lfXxcSY
SsT2wJ9BC7pYOMtqO+M9MYk6YuBkeEbKr/EosCEYPNPgkYPh7wu/IaxwQ/ZcmCim
9XCb421Lwyd5hbmvgOtJN/fcIDPs6zExCdBOVi8wrU788QCcXYdazZZ3NGXRDRAd
O790yoevV5q1XzAyQjSMhuld8ylF/2uQmiy2nRZJBDVXcL893Mfcm0U+olsQc/Qu
D7IzpaLNm2N3SaTlUoHn9dUVZJEQX03sGETHyQeysaAgBlbGgRF5YgWfmP8oZhre
a3aJs/hO1QTDLsgbUcmvY99R6acSe6V8/Nn1bmN15Ch3pz9K02+52Ogqz6qV+Iv5
f1wcrRQ8oP6O+SFUp6ckPqB3nghCL/FFyw+YtCYvUKXpvbAol3AQtbXnDKRQwwFb
aYBO5svNBxC9a4Y+oMPqUONpiUuZ7LxhL+BUm+5RvxVMuzuOEBg0TrWaRrXu/2RX
DR0MCCwCZa4uqcynxBVd/eoX0uT/BMm+n1R19OS/DLTF6r/hp/XrzpF+pOFAcNes
1CtB3zX7bRoWIeL8nm7h26MF6WYEWtBupVT/FvC8fNcEq1KrWbQejSoYAVapvJ9w
swdj3YZ+h+H7HQNrqp3B7pLdP1NIwR71iYWbe+opTi3SrJid62+qbrixz1yPIEPc
0lfyvYJpNWUbc0oDtdyJVtGSp4+skjF4IlzjoBas1d2noid7vx5YJd2OoxNYXMb5
Fkbmi3+oMdgy0w88LJHWj5XZboYkWDCpOrNSzC5a9tPmI96+I7HikmHR+tddRBTW
nIFf4AbrxitW1Nhu+KXtHSg4yzKmaMr7cmpDu2N6Oto4EgexpnP5hhgItBNiY/pM
ycrzRdMWlQa4+g7yTZmHHEagj5L7e9LpDK3Jeg3SPM4ObunPkyDWnklJ30NCh1/Y
F0Dswocm87Vw4DS1ndbycNZYcufPHmjKEdcJgJrV7xpAkY7V5a0/7xB4PC+5mEy9
/SX3d3XmBFp/i8ssgZE3JjKC1eI1y5wE9HSR1lRZceABmosHoxnU7HtW5pHNoIfd
rQLD3iCjTbFmuveeNRbznDuJjSHy6jy1IDjgcX57EO4jo1CRZskhnAe9RMnKpWSx
mP6ft2eShebveri/trGAhl5eGl5bl295uINYk14PXNWB7Ipqc7Sx76W8oGZc3SdL
tH9cCeUZvmh1HLHp3HTTXLGfWBGh2AbpWf/a9dHQLjUU6h8YFA/bqWnDYazmrEEN
lX0ApPwcSmw9txaKyLu3n6nE96C8aLf1LsUhZWYWOzoaNqVtcgt7Z416jXSp+iuE
skZg9gjEkc+MLQwp0wkDvzgCGow8WtBk8kpf8W97H2KzHUPggYn9JV/et9g/GYqn
uKQTLe75uOxOaJsI8mh+IQsJMPqhDBgJGSRAuL9Y8lSt4Le8pBxDJ4T3i+AEo8fZ
gLXW0dY+86/B/ty5s6KO2fmgbHeQV9mb0ZgacttC4E4ljKhn2wuUghTO1DKi5d2K
smr+Ku/871vyg213xrj9OtN4Bl0alsMwKsTkqsXQQaoAHcKj9GBgPXXAk876GS8e
lHa9bUJMLM55DpwOdZh0lOntPKUBNEGaEp0T4aTK0zhUHI7GPxzkPpbfB43z+knr
9BeR/nJUI/gBihS9MTByRrDXDpxfXjyqXW5+OoskpXULksSkbKqmCi/LSMNR8Y6K
tx56TKwR6VKUXn+eZ2Hld2VJ5TaQV23fHVDyss4OaugnLjZzttBIEE0gQ8wYImem
Un7t93q7fzskkd+jdD0015t7v/DWi5jr7JFv4bNPhk7pse8uon/QGVy32b41u1NG
GJ06SUg2MYrkTuV0+M0PsHzRKHskMxqBDpcDj8ioIhMx8UZa3/3TeozSiE3k45EG
1GGuQ/97k65iy3fEHf1V/b7vQDO2df9q3ed33aWbGqYezpu9gFgqDB57U9sPg/I/
hWIK5mMQF4gA6+DrjSCDZVdlmbhFa7nTm6PFi4Vh0xNC0SAhBwFur4nzqk963Fv+
nUwaV2wClbUyxBKq7ZPJBaUshkKQlrKxG3RIGyLRBxcCZ8Vg1XhbBNHztNhEwAoX
opf3YrmtJ8Ru5FgnTxFSF9hxm7RNnvktlrMZddqJFrM8sUeVnwmHPePQdrJGVaAj
HFOHxa/XVDzRLUo6svLgdFUueauS7eTcvPD+zEb+QaNGdFlxRHwxKcdZIyXJ57jV
5w8UQGd6ceSHt2guJN0JoSE172l0c1DjVnuapytnHBDUvpy9ogCl0KVT3q2bO6oT
nyo66p9mv1x09keBzAwAQaVf57VNZHJfXAm5EUDEhVo20wpuB2oCHLDAKgUPBN8e
4htzo1PvVRmTCudgTbu5KpAREdV2Wy8sWtiUyC8o2fG+R7NeNnechB8B9HBy3Bv0
c+DmFQ+Mkmh0HsHSg8syNf+q4KZMsngQnab+zqV8AVLzfv2f6V8oH9BBabvqUUuK
KYFOeuMubp5BX/8Th0ZKRheXSYg1StXLla9MpDv8GIweqz77S2SKahlxFUkWozEY
haqwAsigLDAFkZqrML1UciqFfPQaKQo/MRX0BQhZqQYivfdM8ytTddjBqGT3k+cQ
9RuYcYbp5bl2vo52EjMZv+R1g9V8jsLZ069Vc71g4qxqCJVxjdJ7iRecMqzbim+k
crLCsD0I1iZUC4CV/MCFz9xDWnHXxW0VcX8Q2OrTsIfS0BX1Zi74BQZcYptde+Z/
3yyTOcHSw2hIkoX7UcKri8LEdU/1Rs4HQqAySjgfd6PbMMvIDUSNvy4rKwunNYre
3iumvlESlhxtHm71heAQQTlSsOKnYbvedVkXNgStWayDjivcDrMPCRI3Ts2tdMzm
nUqzosRVr5R6kKjS2XZqXKH5F8kYqzl7gZa/1apM/6QeM9abGhH+ig8dAkQx5QbC
DLTKAUjMsT/Fc73eXR3buUItIe8425mCUNWyZIOOAy2qRJJ+g3SYfJzADdJ/BNn/
SXCJwDeQwbbekXavR16D9HB3rXfMkyp73cWEbxHPqbXZAXAJeeEOII38NKoa3dKA
ZJ7LIMuRZtQSdoMSZD3dyxSSMhAncdSO+7fWmmmrTI++yrssiVHRCgKa4UDqCs4G
gJxYVNgXY7aSadCBi2/FKg9nY0dXs9vAmk3Qr6YVEKLRp1MNHWUx8iBZXoen/iSx
cMfkK4qeMRtRkGXQiYwrMJFl2URP0dmMMokQvvl2yl1bgf498h62V4zJwpK8QKpY
fSn765swTFaM5/aXKaPZ2LiccTThle0t11ZhKQ9+x3v/kKcEPKkXvtAoyZ35xjd6
JM4W1gZdHw82CEi/vSTV+rhNSb+ZiaD1G8IMq4lA4SLYAk6PeJJhJjBUJbMnkfmv
EZsq3wcz/h0MJsFwLEdwFn8HHu4MIRdZzO/gBCxvRKUpXAhWPFtYYWM7gSpNu46A
wZOfny7obcvC5jMKeNA+okld5gcJy/Cd8dsiOnfyE3Fjz/7HNsxw7juqcD6+DsFK
YjTOVrMFFtSvgjCkD4qMEIpEQOWgqc7m6d1vpNct2PcqZWnVF8nWRG5C74LT7Cu5
ij1GdC4x7xyOS5KszHLV0sg9/x7USQOLRFD6aNo7W4CWdT/CDSX18WzTsCdRvfyI
vJT/+LAzOrTcCbNHaykQRs2tXaB4RKqf2WpHS2fv6NoMf34FRI510/bQXOFc+OJT
vQyBWQoSTGxRhsg8irbtOR37MX61NcgvdduWcW5ocUDI9r/4jmR1xNbmz0Agkgbx
QSW3JHXvLypNEjKdEOexmrU6wAgVaMQgn9+e5xCdW+7TGrkktdMYhgos0px7aGur
U5101+3a7lun3iPQmvUdriPpeqre4i4KaagvFGHG/LARlNZrF/w3/JdZX85rPBYd
5jXCET9a3x79xE0AT1MjWNJYGFF+mT2C1O7COP7eyPs6VlAve7RZuGnGjPpKeO6E
01LsKRMjDpa/Bo9bCzwp5RMcK5IKwsbAjPFX1xgWKZBTHcvNONpuO6nEV54k+Fvi
PRf8Uv2hMfAFRxnx6NP9Bd959Z0w5i1Jj5XO3lFeGehDvo9NfqaJL7V5TMmJZ85g
4w50g3q1WjIxOe4mKHIb+YUzZEpRDTfSRG8hUdkfFVp3Ix7g8DKl81/6V4a6Clpt
VLQOhZvtmgtxeQA1k4MgElntfPYnAXn0VWpEFkuXOP/PlQ72+ZeZNvhh0A/Xfrae
fipxead0COSB/N0bxRhu6ZCITrvgF6o8CVhPfYqQak5ZClI14qeSxpE+Dgmqd6ru
0WlZBrqRaip4Q83PbUT90vy2vN5cF923eXdas4DRqJw8MFNMgsby5714MY31NwBH
CXFW4gMmHrxY+D3iriHs9JbyfrGZKz9n31GOfzVWRk3nx5TwyXdujzD00xVhT/ay
8muNC0FFY7LyGY8Vm/52FMxo/dEbGTtDvPXA250eRYuWtjbBp2k67NRILv2mfE1V
v8q0M6tMzdOuWwI37dFrCgLZS6hQQZ4FIk+1kRoUiLd9GdxWbdzKw37XaxBa+ghX
1Cos1mOcnzjGId5rbBBnTDRwBSQ3K3XZO/0xifkyPq4MTsrhWqZm0mxi0vzOoh5q
x6eaqQs2J0jJ/BXjKv4K8RFOIGzQ9ezUGfg+1rrQHMQzIVgXAU1MkBf/7fAVhz9c
FswTCzE/FIXRVaFtr/QBkYfIpFwH5BZudXWpfz+m2XytR8b4wICFBMgTNVXfooiF
C70iwPLPSBAGakl02XQ7Wx13y9ssaByCfLsLlJ6SpLM0yEq8/M01VQfxyKD5S2eP
gtnlwG/O0He//ybwrIAlldcuk7oJTTExn3Qxzri+qGX9bPGBW21JKccziKzWegQI
Q9fQVQGkZkqu7JUNiyUioa6Qti419yBNcWzzdBiNQ3VmBwuvZdrQYf4Xgg4KWyy2
xwZs8KwhY2clBCLk4GuFuom5t1Jpo1LInBKm5V+Ld7pt8KiFZ2xRg2FR9BqedRZt
oxhxyZNGH6njLD0lAVIPmbkyNwVKAq2/CWbDPZisjlC6vf3eD40K7loSdFeMBSuT
qfmDF6Ox95hB4qobsr8beOIC0PlDE3xGDSz/3lsKAMwj9RKBRFZsOFCTfS9Tu5XM
trB4LClx/pg7GT0lqU5F+/Pxm0z04SnPyNlNSOL3CPkJVTD8Ah0CvBCLKpTluk0s
XaDqIe2jt4FUcQ/zjE2+0dPLZyAs0ekkd4DkE7rQDIJX0IQciJHFZsj/cq+VbOhW
hN6iUWzJtEgseHodFEbjIneiqBwQsREENMTgpO+hjPS/N6AbleEY5XcG/7HXWvHv
kRRUieeq7410hoO7vY/lZG3RjzhTVnQEh/5CyYL8sT1MbroBUNUflTTmpk4J/pdM
vqop9UL5daeEc69sq3qyu49bp5ySQYuK/PEEWDVAfb6lfqkpdGHKf333LaDfIOJe
aigdG9pvmJfiSMkaJce3mMBRcp5z76CZfiUCgEcAgDlomlRN12heXzGQr01ui1n9
ak1a/YJ1foYKvuxikNJeRKOZpagkScVenQcLTD3+TN1M2TB+u3J7OkV1B69QaYF+
w1jli0oM0EGKA8OuaqmlqP01X+KxOXy0SXC7SBN+vnvsn45/Wt3/YkHNkOEvfKoG
I2tr4WkvEUQYQcZK8PZK8Ip90AMO7MCD0tWbTGsvoUcIyNXGcMGF4lJ8oEeXbwkR
lXLMXTzxJKbryUgTshABnIf6vDaBUtuMiMgP46wqbgLxZkeHOpFOKa/wjlPMf0gI
D5MQSvzNmEa5rNA30V7KMp8WLwlDpNlOQsYbXMu20cw5Jh0eUqd9gw65KbvyINxF
yCTykxh6KcqEz5Qyf47IzQi5DlcRd5zIZ0BnHWRG7GhOwqedCIsYESn9gh9crZVr
dSsiyZdNbZ9RoOWln3smFggkYGamLJPux/YbMdCUZZiByrkkvIUSvWLFbtT5Y2ZU
wQSfkC9lGsUii0M4unRnnCcm1MfNpGJefhMBKDI2AkiVZP0jM2quKyI6yz+Yce4r
6Oyazyiia+BAm2AWWPlkZHc2dXIK4HVMwU7qGhjYd/zA+iuSqTYAA1XiLombIFLi
QQvzp5WkSSAjaetJbzISt39/+JKWRwYBWLJPFkPuue/8xBdEbhYowcfG1Y6mNVlJ
1fWnHZjpup6il930iWPIE4yoTpWshbzJA8FRftm8IzUE3h9j/+D/639bcBPYHOmn
GCWYvallummcpeUm51Ome6h5o8Ax0i/6xoHDSAsLBAGZd7cEcEb2gDodQUFTIB44
fw0HEDWYL1wYD8sMS8Nhcbu9iX7FD41/n52ATFXhSUXf23Ljjd2ohIvmKHmxMv16
0+ly92bWAnCGEZZxp2ugLAepLLk6cGUKCtOu4wwklOJUTU4Oqsuh1NBilC+6xjjb
KEQEzWVA8Mk7nn6PS9kEbZwmEanE8udZzd2wBZOw/g5yjtM1OVytxa9zc/3k+KU+
UrCG2UFNvPL2wlUeYIfFqHjBdQ+GPTzXcubycsuruS/zMV2BtPuspiTo6fi+u1eQ
qWX4TvTqpwOab1/LxTZt0gI43NR9bciKk2IYKqjW3+VuWZTQD4o24MqdTLT7YYT6
whPbB9M1ZQ0SBEyOqpVVuM3zjLRRRTsnv5DbGljXdW5BFwuE1Q5GGY+/l5Wgnlws
YpPBo63LRp6TDvC1N+REdK48qVLL0aiR6Qt5lPELPdjzS8u6+DxlNYF5kAEu31OZ
W580+nU3ZIO6d/XDAsxC/dDo7JRVjBR3Dp5+M861puFkorKzYxkvnhWrNXTmVW0E
uWAKQ8hNs8vC8xJGF6tFZPDuq1MlVttYYOwCrCLXCOAS3vZo9cNju+YxBVR2/qQO
CRD6K22iKpBdn+0r3OvNrDbs3ldVj5TICDIpXkESwQJma+Meau3MJy8CJpPnV91O
0cgHxHsPj0RlMcg7a5WG0O63hgYBQls5DJsZKAnUWGdfpfmMO0BoHPmUPcWtB14m
BLqGo9GVA33C3UDSBzDPFLSMQvMx4fYsSQSEbDTxS1zovM0LghMohzaTG3ZHWbNq
LGh7Bzd+hbd6y1H/CS8/KOqM/G+uiIpj5+JbRlmYVJ9UVRvvH9bX+5bctrrXvSfk
hjllSJABafGoMWmtjNce/VFu08OEFEtxBYN9vQ83xeM/tmb8JdjvGDHpPyU6gM/q
MSVq8MWhhlb7mkH9W6Crgp9iIh/pRS3f7UwMUV11pvWQuU3B/5fx8l2pTUauNeQh
x/i+/ch315jrEZ82lx2HEoERVogvbuKjVaPiWchUV8K9u4ny8QnTPiQ+dnqD0WxV
wirfUoHToTHZgB5YviQrqp3I73o4MUIvtiiAnfLkRr81TMvE2v53wgxoHCwAchNx
crDcPYq984pZa9/wMRsC5VcPcIy4lzI35R1QXF2k6WRRvDV4oKfEh9Y5y7bQbCjE
Qs5dbyvnCSRKhRYRQ8Pc8yaMJ8WT2X2eV9zUE/xofx2JezLGEAD8mh36HV37l7sC
xDnucW5RT53WyLuMv07zUwSiwO+hSv1HauQSTkmRL7g/AKTliZd0Pa2xu/Ldqpah
kc3J96I5skXqFAUAv79GAPMexpxqxngdfO8lNc7+pPNWY6j938sTq9E7sAsbqLn3
8sVzF5lQjMrDlyU+flYx/OpAdbSFBjlZ8RHw/q+E2iMXGu62a2A9RV7AhcCBtzcZ
ZiBOUuTEETlrrs8dF7ZyjhX5EdlrmprFsdRjjW8yvtpDKqlNaKdxhvZR2+RHnR7G
QDLt7ds2KGpy2DE9UUcr8kw0j9vCvuZ57nJgB6lMNOyJZEfDVlp0MbnX6RToO486
1Udvzy8wPHALCyPAahesF3QvUA8T+lKNfJaSdlcMp0rmQ205Cakyq8INq9LmLxiN
t91+m5EVnDncwKR8abGO3r/ExRpDZkXBABgoI4oALK1pewTZymcVdYQbTwjBmx/Q
6EaGH9tV7Gho6/2spyBRZ1SBa+TNkPgWtcY8QS5HUJ9Zf6HNoKTo1kKlsN7TVGP1
2rQNz3FDxauj7jz5uHw0wCWeVqRmscNkifdGMbH73gf/hCrrEeaOHyLIxO8LVGnQ
SLu7DXB0hBv1qsg9YwqFnbZOQHGOhQohJG255Az724vysBMn/8oga+S0yx9YHbH4
Q9MTuF8GLv5J0c9biQp95rtXfryRBbnWIYiTZ0OBRi/FcK0VgaLG+vDsmA0xsTnN
pk3HyFuMqk0eAFn+YRUriBHKlTPBGALdu7/p7ltBf7IX40/rD8ROzwjngGea5/+0
1HusT1o6wGRqiWuFmtjz41BbYR2U+B073gBa7+mVzO9VSXqQxoiYHC+NIdgLi7Ru
AVa6GE14lgJPQR1mSkTqgudzwkoHVbqpm6lccqGaHwlbZ4O0WtX2ObtQMueo6b0G
0ugFLxn8LM69GFBO8OAcP/87yzgAdlNNYZi2sKwTT9k5SHkkF35iHWzb/46sfTaC
TyydEkE37uc/mpESkaji5Iuf4lJPtaQycCv7Quw9sy4=
`protect END_PROTECTED
