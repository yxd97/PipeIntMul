`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bfCBIfUHEf9lFUQolzDhZzoqbbVEbYu4jkYgn4NLO53Rte0Ypi8Fb80cwtgKT/I9
AI12gic/P4C2+n/osIlpMedIvo32TCsDvYk1rQlKoIpt5aILRVGXlTRNTenZhiZG
Oe/wicNlEO148EeZeboEZcFwcQF3wj4eApLUfdcEJy97p/T35irE0XHYmrvbrwi7
y1ylYWf2jC4rKqu75waHITuwwI0ZDXiyvLMFix7O+0KU2DsS9fcLoqQoTguoPIo0
14X0vjZYejYtFpFxPkVNHdpjkj6xTu8/gaxjovSwkPXxTWE/RUQ2wkTRg18NTeqv
OtcKuKK4ux6Nu2wDa2MR+rdcIP3TBrM1gphdyLRHytnMIdHafBRTbmri4WBvGRZc
LOuj3UmK4nYMW8iU0JMmNO0Qdkr6SPhAVLA+gqn3WQggFNa6/gMPa/ClAbxcYZpZ
+ruuIxCbRs7f49WqOVpFaE7qyeZzAtqEHWeaeqba5xRxhp+ujvH4AatZddOGJZO8
3sGF0K5XH8tTUQICxmf5rvrF+ocVa19hhm7TSzFQuZ8Hi9sl7n9zrzVMo62fsSLM
OyQ53nYRfZuSwd9wFvOXihJ8HI0WJ7AfKn+eRyl6hYQtfnsidt++gE02UaqFvGpG
4xH335etIsvibgkaeR4H2nxpuNdtm8dJAwqN3fkI4hHVBY7guLqYAsk40P7Ye82P
OZ0W37QENOa8Rn7d0qc8mQb0EJREOrKHPXpRnH36iIAqNlpWPhltq4QWc7Cf34po
t5Vr53zWuPG/VcdABRQfDLK1DwmzML3SQnzfZAdC6GxItS8AumN0gJ3xfqsc++rH
RXfRD4HLRXcYWNy6g9f7h0Y+nuUjEiR5KHWeQfBGc4LGzbUuEzmQLXgB2GnCXtkR
6wnRMIxrj7usO2XztolUAD8Sf6sc1ey4uizSFBo/w6+NLq9tsTrwOxcMxvXj++dx
qZTc0dbbm8esiAA9dMRq1Q8edRmlyC47apm5WIxCGES31KBVKyr13160t4O5pWS0
w4hM4h/l8H9rrBt71AJTPNuwRzyqsm2nEafv6BMkv6VxnrjU2QHi60He3qQKy2Dh
w03HyjGJTt7eSGgq3mGeABOYIDj/6bsEN2F2DgDB/a1ZYin1wZr0QR1HwW+0V8O3
l4Ylg5kP+nY8JaFQQOS2guiALejxXhdZV9kgYNOcgYmiz1EWr8u4X+ePbSFgG5yw
8bKOfLfQDL9L5bAGBnt1YBhp4rPqsyy5lwgNY+Hl7YDjHpBN/FDYdukd4Y4C6nY3
r/yuUm7wKvsvhs00DxLAjhPfXo8bbhatXotJtFedq8aHGDRga0kuc8RLsptTzoP6
floeXyABH8bYPSEDkvSbwlGNolEsm8MuRoaPuC/Xuff9CYh0OJU85GFmUqgHuLjO
cFPqo+Z5n/i6Q5D6AeGWyToPE4iN2Oz2dYSJN3BDVkCglVEm70NpdDn6QK/975Gt
X0jASU43jhgMKxd1OHTWBsb02HxSCaOVwfCYhVMu7sYK8CoQgVTEQsZRqdXyoWh7
bCHk4K9UUMZ/jHmE4xdL+wv/6VysttfOOvke+he8IoEM0Lwn6QzCz+zbtsk+Nxvf
C5qYKEO9SPGxbiCU/r05WD1UOlWKmmzg8ef8RpVNxmf3rIiXvQT1djl7ZsG0o/DF
n2wup3T3K2RssMhh1J6Syn7V5z/bNWQuHrRDnjcuaOrjpP8G5Z70miP+P31t9AV7
7rOv5LiPeEVHbXreZGZo931yQ/BxDCzsFuHBq+9WICuwkmgHz2SRm1OnKfvPA4x8
zcjIBkyXbeLX4S6uqtBfZ/24Oc36XYKxaLkaeaAg2/c1goOxUH8K1J8mSIc6YsWX
hJrByeUN61zoc7Cts/fz5WqwHxfTKj8Z0tbpFZ/zK7gsHKHGylqBiJ//YEhIJpkX
L3sf1zWhDm60Xzl67NMQwfxf77JLiVUh2PA56bnUCvqA0MFpClS+0IYixi2h+4zW
tu+prMQ29DR1ylz3Jq1BnwhXA3BTBRGDnzVjKzPPncj5wd95QY3mEfVS0Pw4j6Wi
5tSvpuVVWZOupA44PWhugJoI1vLJdbkRxh2Q75WNHppOeJ2mqFfgNLzCAOBOMaUr
+d84EXzOhvwSw+QMday1N4YBrn3JrUuKWfpPL7YWU52phdmScn+d9kphdM6gZRUM
vO6VdU06WIDaHaP9Kc/QA6cr6UU4tNVEX6TkH6k3AiUUY2AKX5jqKdVuzCLVVImJ
gOQDG2vgAlhcqVq+7aHIQsQsISWz57b2LHg1NRmXoUmNfPOAYwDb+W55dMk2nNTs
Th6sIFC1xwxchF3aazIMKfqj0n31zAX6e1aR+3p7A29VImyZoXEMjgdA/Gv2fJf4
lObQdGLhqMwaU2AeUAgqb+gQO1Q0lNFhlO/azCNcHoRfsY3TwcZLvgCrouKNH9LI
IHkeVRrQt9QP/wTmRCZheahSMrYnxO0qpLAODeBi9UUQ2qIIqY6MMBajROvCVuDD
W8cG8UnudTE2hnOKoHgWhDhIe2S0TSN2tozeyKCErvqO0T+s3QrwhtkfZE1+F4bq
0RTfxTUBGTwIzBrxSW9z8SPMcziopbmGmYLqcmZWIKm8nApywFs0cBM4IYHtCDLy
HICC4LdFbo5lqH51NYEussUDAm5pN4kUls0xQ81jbfYewaG9yECzy0DDNW4VdEbg
fSU1givewPPDAVVmpGc5cxynzozqkVz98ttMHjFTbo88wAKB6MflzPLL7Po7yWna
tcbfM919oLrQp4BStqHBA/UOf8efYR4q9DIMixTakqENqszugW0nr63WZGqV/5lQ
LLhc+1TE2vmnuBs2BABkq379AyEfzNaZkIIv9CjjyTN4NGiqdUif+UIKMOPJvgil
B8kgcVE8OkziCxNpVpn+puROkzmQP2rxHnzSA4of8iZfpJ8wbAa73NJVuOKg7QWw
QQ1X6Q7zV9Gxv6pEZYpfb6myq9Vp05zCViE3jNDnFiQfevzbyp4l2v3zZZOmUXb8
496d3xghj3I+i98Cl8CEzPUEwbmXHfB8WBqs1kEcm5uGD6VqqyVn+WaWLMcV7eet
T+4m4UelX3H3jy3qp9sQf1nLRc9DGOIvBm1nEQjwL5RyMg1D1aXTf0Cmt74/YsC1
7mH+eYr6ZM/e7sU6s+ZJfYcVH0myb8LLSSRQFRZA2+NZHCSnjWe7PJ9oEkJ7OdFu
sT9+LO67Pm4bxaUd7Nqm4cdOM2xE68bN+8p7e4rUkrPqM6sjOiixfeTmFHCenHA3
D+jS8PoH9dAFZNH1MYdqZ9BzIR+ZpNjYf6m0yJsR0bvId/TUL93eGQHtNd1Nf71Y
1bpGd2VGrN04Qz1pHhyqqat/+Lw+sFakZK/BfdXBVFSv0MqXKxHfphCzg3pVu99B
fQ/lUNUaI0c8JEzqnzIRKOQooyAKmvjxNnSZ95h+Cc51k45PKyBdkGCkwbTmObYC
w2MG/IPiHfizx6TVXejDBiOt/reuoF5Pf9z3g+7gIr7ZW1bWj8ggFYL4sUYSfKct
xAUsjSoTxpSNVkivzNcAQY0k/YWFU+7Aao1Gtv6wM0llTbY8IvcdQORokW/2imS3
6/Kuz8OdGfnpHb4Rkp9oUmkWIfFP80At7yIL7QIeQR86WZs10gvFLGs0VN8fp0wL
WbK1TXyPGBv1pTw9GNRZLzXUbLaK6/pr6DR34drx5gqIcxgbLGj9eM3p3a1qfMte
GecgCn7NkRaOCG3DJCkXFRUVFGDvYgi4l2T3duYP8/Ky6XKISweFQp+Nco3BH186
Ol2Npyr/xZdvyWWZ9MOVBVLztGvD38TQYUG9Dxy6v9kigo++djDeVS25J23yK344
0+CNIn1SuUOmOF4cPVFRftykeoT+sSf2POdm1sPkRcB6X1tcZsht6T7EH8TaTWHi
+tbDxgShK1MzirljbtHrT5KvZY0wGMwiDft6vLHB+fu5J+YdbgXpAcDjggbXPvBo
O3CmdTTPLXlGRi8NxbBsS41h/TtMa5YdVcZzcThPpTXLYCFX4e966WdDOsulE8x8
JY7r7VGLcdhL+2BpCscsyWh0K6Be03O7npzj761+/5Z9Fnd+KaUT1dud5djYzeUH
HmeOWsVUE9GBA4bTdbodKV+qExVGhtVjXdsoyaUsrpqQ442RyFdN6/MmvL2e9UAD
G13fQXE8qWZKpsroW+DQPuIl0UWmz24vSK8GheGmgACcOeDoeM9d0B7XPHY1UvRw
DhxJ8e7droEGRUKBzEPSdCCEtGbfh8AF3jn+tY8H+GXlszHQnbNszRZITt6tTJun
tCKq2rmQ5MrpiUusHyKQNG25rOGlxdEetF9J9iVDHDAjmLE0fjQ8JhMSd26eUVHX
1MFtE+YXc/ByK72Ea+agXNoXZr4j1ydQiFBZkBbzoayhseO9tnvcP3IxBsm8/eom
rE2Yl5QYwZFLlalJ387WUYe/z9ve/mQS79WmqBIKlz4cjzXI7wgWaWfsMlQEP6/k
7GK4oXEkUnfTr0ADqlAuCS6oeON/k8kWIXQWqLkExpYqGpHyYfb1o5cc+RrMenZD
nicY7MraHUDrU32GOzDBN5jIoK3gCrrRPckDDKggvfXntlIC3dPf+QLHaC54EAG+
4gchkNjx+O8b532Xe8iJP5SN/e395XrkakjVxnr/WuiYWb8VmRcFVD8XCQKxTdeX
RdfwY4N+dnu6SrlMMJFwM7io92C2+UR+SkpaDVDYS/Q2l1CeWuYQCC3AMOgu9XR5
Wdo6TGYxGhEFTtFWIrO5KXZocouF/fOWo6Bto8kIIniAMD3ihirQn/1JXr5l7WKX
QJ6PpWPfIQBvHLQK+0LRy5h2OaTIU+3ZZpJko2a2+F5STdD1L2BUeZy/wABev8zC
WWd5sQOspt8oSbTaguqJMfzCkt+7nNw0WykNYEZDgTR6DoilQDFmrentJ6COz8sY
wAno2uypdL9lm9U/4rqC3z+qFHP5Sgu3dohImp9S+MmxdudPB5PDFq1L6kOKyr8a
NjcdhreUpUeyX1jT8melIyyLoS3Sbex2UJJneZ64lb+kDJSJRgf5+20MH7x6oXnA
ltR9abm+CHJdDoZmX/QPUT9Sk/WKRojk1ZTub6LUS+cGhtZbXnGRYeki2eyTCqNn
Vzrr+r0K+hqxpaZEyqVe0zAT/V5qEXJzseHTCI7OLUfi43QxEqiBhHFyWX1HjG5I
Fg0Bpm8JGdYA0+zuDpC3Y2Fqb74+JF/r2q0dFBDOkJqYavQri5ytpvtfckmdg0SE
1aLJDySRiQLXNo63GiK+EztR5Z6Pvf/kGhBK9hAqtFaUedfBtsOyWqNrWONOpSVH
E21fjGArqSsOb7m0rWmrv2X1DM+LSKUzSvc9hrM70s8W6h6xRajKZYQrQSQ50Zkh
u+Q/UV2F/1dHMRw+zYYblwfh1XfPsWgHogqV/BTF2+l56B1DXyJTWQ4UUT68IUBg
tb4rTrZheLsN0goZKm5hNs58K32ly4N6p/zZMmrHk4VGo1thoiwUwidFG8r+JWIC
hyhbJMiLWr9ZNcEcxFNZDKAB3OUb816XAaNsgWoWJH6OYSy4t4+2LavST6+I82H4
Dor7zNMXz8JuOiNfh8apFFqN/nOQKtDbL0FjNncLZ+9SS5DXeHtU7CuNQxqd9axz
HYuIZECRU/G7i6axCwBv2+NEVaCnVaux2NmR4SZwFoVqe6JxpKhaAUB4/mCpmA5Z
5lBmZFqXTxDshQGn6ISzDEB7J58FZAMzX39OTrGkvFUxJ3lBfwRGhuPHeTP/Hj/k
d9omJj1vUM52iNBUPhju00hP5Lw1jqr+pHfevAmxpdXymW2H5QKQLpQ0KkAgAv5J
v9TVdOTlZDa1OZ8TM2h9vAnsNdi+3V+8WwN9RwhVECFd/vkiDSJDD0xstYBWt4mV
mZt2ghCXGDj8BfTnQ7DVrc5xXD/Fexha3Pwec9N02JhZZYGYNb4q7VM2qVyURVTg
x/6oRV1U+LDqMQKAOTOIgaOZk96FvCLMIHkSD9S+rUveanqA4X3bFOqXfenoOgyH
4QdvNFrHdrMc+biZtTxYvClIqQVHcWjDk07h04nRQr+yQSe7sroZFyWJTjliqIaM
Kx9CUVlI8iVPcoE0lb2iAlyz6d4UxPQ+T5rc/MAwZPI7zI9/3Jo61kIk18AJYLDS
2jB3dRtMo5K8CX27MLOvZFZo7wHBqyVYVIvgctBx2iKL5Y7NsqowMX4WQHHqZxGP
K3qNgmkT8nK0ez89QsaslDeKAu+kVzOxAl38rT+fokXxNVi2F7tRfqc89/vQT3DF
NrSTtoIORebEROB/l3yflznudaxGWpQvbziR7RuvHJTZtFASEkN16MG8WNHDjJhG
UnerjyHIsljqft7xTdxtWuhjYAO++lO8hxPlVFFd3kkmEIMoPBLRlxEiSvX4Ts9x
XgD0B0GOASEEEuaDpqIO/NAPmaJdMoUivB1xQMHJ/ZkRjikwfO7eSvrJ5p6UjjRD
DcaG0J3qy2BbUiB1LJODwiI48i0+4MJMzHK/k5YfKM4U5mlaE5pwivUXt1yp3fji
axoaJlDGxbE6FmdJh9eL6g6+S/Qe3aWEE0LZiM0Nrj10/BwqId6AC949/Ez+UyL8
QPOPOOgVPaUzVlRWWyyR7YgDrcankAVtkyqK8mF1Q7s3+qK5qrEXByKgzkdfgBod
5nSCVg6XoV8aQ5FIIKBskbQDxhO25bQRVoWx4CBuJNVR3Ki2sM7aH7B8IB1pK3h2
3dj1BIRHVspdlC6wtfga1GYuNzAI1wW56lnN60TEdwLTLxKdunsHyCMS0IckTM1H
cwea+Ie1Qpr+tThQu2CQO2lL88xXcIX4evwBVhsBAf73DfdphECi0t8DptLoH2V3
oNctWThcmSKepX8QYnStHKKVbhKCj++g/DB7x4eswk6chK+z6vhmXOeZt+ifEPVc
pneyKYU9YcLPkGz+h344Zyil1fFrUR7Zu8RbZwSAiMFSqgR9H1yH6Hybq8UQtaBp
hGaxtzudPrkE1FCKESsl8OYHHyPgfSKN0vOgyGtwaZvbj37LT6PK9o0NUHrx/HJV
QxA2+7kG20QuqW8Q0WEN03jN5kKCGxtZpNuVA7fuR5ruDuj2EXfDOM7H2Ep63HFM
c6FSytaIXKzj1MZh3q6zYLeaAhUOuZXTvAnlKV66ubazJB3njlJZRk/AQK0Xq9V7
vgJdaifnxx5d1bsWm6RSFp33O+gkvfyvVUdjCTINwvdCR0/lw4xdInzSzo5VctSc
zObwIsXUHMnOGKxMCwRXJobKruAPi+fEG85sYlEbQ36xiUULHE/vwlj0Wzdn6wWI
r7C4uoDzvP/OYQX/7GNWLglgSKbykwLkoBfqkIt2X4eQGjSrEQGyk+xGU/sSPh0+
5tDNxqbpR2mVz4s9DGSKxroHcECV4LA5IiyrwSEe9BaLM8V/c/gi+5AloHjxxroA
/0zIibNlxxyBj6XoLkvbPjRJLQ6/S1FhgAC6PfPV3HNqoctqjkfkgx15v2fNUbeC
uKS89OhoP0NjfLKzV7/F+BrZBdD4Jzb73ZapWrW8jbBE/W7Q4OEhWoQEh4k4WNU6
5dvXVrSAK9NNZA46hl3XM+BfpVIo8eVXtwZlCw+aoVTt47Q5RPM+PSXm29R93WP4
e/CYwUaa/l7kwX8ZDt6uGduJRN4S6iUDsvysCOz7KeXHbxyfmC0oyQ/VhyLDyjmJ
gWLBgREi8dM+m6C6wMiU8UlEEribMPJ0+LGQFOL8qEShCTGB9rHU04Lgl1+q1tjG
+kw1YzPYBx/D8jrgIk44fL++EgtWwaiJOG39zFFvGBou0Tg8TdAbRl3eo3fztQ/n
Evuux7kLTWzGAE0AjyyZwdp01Plksg3zJJpXDhfS/d2XVCfEI6j5V3mA2rWQLy3E
KIMlcDqVRQTcMqZ6vs3SjITp2CN5SvFF+HLEPTAMUbQ05na+TdzycItPfbfqHovb
2snfZpcc0EIElinGCA1isvEVCAcBPzw3SSpWrWhHbc42QiFTZGdYRIRGg2fwGIJk
vJIbG6qeNV9ppFWJvFYlI5f91J62AeYbJfo/mdBQJWxS3DJP1hA28WErcDl9wvGZ
zjzOOVYYxvcOgoCxdpXT19+vvFjraLI22rJK1MfBbHJiVHGb6pOipzWC16/dfHJO
JyKJ9f6ud46mtQyctf+NFtfYkM4acQ12VKQ5woEk4jwEE582+vnF+wYdJFdlVaj9
2H7fNy+/vWJ1gzLKhaMfDPhCoy1dIBq9XrbV92IuHa1c3Qqc/SCuvPXxSmEoxy79
PtLie/W4Lxp/fjITLtG77w/twMfmhL3uqR7TJ3i6ZDsfKWd5cWYDK7XQYlwivDpu
0FcybYKVDZI4AXqwgliX3sEg3dTuUuN5zgKOdO6kPZV/N1GN7K4vzZJN2PpTgbNi
iBbVfQ9dKK8YRHmwrJJyQJRAmenbhD+FYLSLqsWosZ7aToBzWvv8XDr50kH4b1/E
Bk3AsXIOujeH0i9CpREPQpf2La/f1aS+vx4Cmu6j1vobtFff9GDpaTj+Biqj5YRf
AZK6YEeCV8iSNf0COJ6pTfnQp5DjEQBlHykLGsvqXXUq+wnZf32lkSF2o6gwF/sK
mXGupLm63dTg3kNpHtAI7TmV9eGXcXc0JNKsOUyupykpzEesgmviZYLE6Jqryj+n
ec7fH5l8ufPrtEQKh5xw4aAr3L/pg6m9jGbUTdtBLvmxXTJWXYygbunNVUyrLrbB
n8K9kdpgmu9FF1EpiY5Pp6hW87tmzlUO5MJon91OeTRqrFIw8VAqHoWxO8VEYB+T
kwkaKV0TtvGlpoWvZY1eGlck3rX1NN32kl2+UvcfmVrcfsFRS5ad5D9KsZdsAIue
dYLru7+7iDAT3wg+SR57BBZyem12ClW31KxnKAc44pWiCtGVB5YMSayzOhmEQ2TU
dQ5j+AUHt6r/pu2vMC2lgP2tfkq/6nqkmx75/vxTIjajFgT+Jo+xx8wjkQjlrGOk
fY3hr70+lKkfqkOm6KyOjGyDkvPABgqAD690WFI9uLq9NlDe7KwB94NlglRLUkYo
0S+tCnNQJ3QKL7cmD/tffK/5hTADy+37K4FR7xw8YNfUJDu+QcYEb5Gsek3/8Nso
Kv2rau7vrMIJSsNApahMsLNEECxzPoNx5A4h9JXhgLSxXq3ICchBGfqjYFsow2G1
jM4g383Vg3IiAnOV/g3PtV1TAeUSlplXQeWYnFQHpCyAuai5TT7dtzJBoMTynzdx
/Ox+xTre+gCDFG2/3PhFJmNWfKZ/+EeFzdfzJANOEQNo1FvazSQ6S+3CbIhLdVc0
7Pz0g70p/MjM6A7txHiuJAhKcnACE5hxHq/srKJpcohoqStojaySlAARckMz3JeO
g8Fhgxkprq5R4Dwyt1MDoxYr3Tl8JfmMQJl6GNh1e2A+IYqgyNjeJp2F554eYgFJ
OPgTuceZpD0uBWb3YQlhEZykJhHi41EN/Gepj8HFeS1NDNlestvdnPE8eZF7lWB3
x4GdSLaoKDMdQKhejPAK4AbDdGGsYtjREqoqIpiWMHxCCi9U8lkzu3LcKBDzKwqa
eSpqrwqv2kCag3yu6rYMn+8ljJ78n4qlJZLIudyI2NM+JqNV87S58bQRR7tAwE1y
DAB3YrWlOGp0+0gEYGiCuf6KWcfAB4wQk3AnX4xP+0xiZKSvccg86aNPua9oYHVp
VgsEyy0iMX6EyscLmtNhON5cAHt2uxzxhMgfR4UvHGvO0QrVRD2F+IgS94DgCf2w
ZwjvSl2YDgUnDrfIf6DwJwNCdc72RDOplf7AdWqJQv6vsOtok/ndthTekEzCfDMq
f2S7q/zjIZ2EgOlYlRrnkQjkI3yj9p1UmEDxIjQg7fJQc6tVZjIDLoVY1QaG0qqV
ec2QdwSgKDAIXWwPPLmBRDhYhEul3IIYL+gggajdyyIiHfinFrRFEtL+ferE/2gv
fPcNdlrQ0rLm7DoU7hJW14trG3MKtNUTHaUpgRU3MJ1ykwNMv0zCuGfXVQpM14OD
uafV/1JESHuE3X2De0uhD8ngq8o7Q5vVsviXESmbFmOChlZMABpfM3V+UZsnplNr
TF8zsptyS9nfNeWcw3uxGQy9ZLTr67OF0rKfib0OClFIpINZPVgnWM9rDUbrX0s7
wWoKepsoDKY21lyTgxpyK4bo1MXXs6poUzdaGfbxZzNGsrTkXTUdXExxk790Io8S
+cSduUYpluG4GN0zDUFEU82ypiM/K8AHSyEfEA1Lkrwyv0s3Uu0tbZsLjKPcit34
K9N3FcwDuJJgMNfzp97y/jD0t70FxdYo/KuqfHtvYmIebAhz+67lbN6H4j0IkISW
z4kQVSQgiOZIpMdG7zyABFvF8dkw/ZS8+M8UdDSceYh5+ZyD84Sl1Ih4p602e2lC
I78KlfK5u3pE72HqRArdsdvxz0NaXCYr9Q90ZgKNsrMeDYJeIbaH362VfjM5GHOa
HnXPqdbIBQEfA0YvAaGZtdvqhkYKTQhAiWn9oQ+RUjhHOeX6C3NkJGnzx8vLVYLp
EF4jAoZNKyKO6VhLSVvZid2M/TjoowTQ3RhuaQvKgCZ346YM19aiJ68UXjIrJ8f+
JkPwuF77+eU0cCIyxtfzciCKn6u/SXKWmXJkpTd50vmyeTVX8HESqcYl2z8l617B
lrV9H5r+LlodU3po7noRq8fYXa6oe8cF0AAgSK+1McC143Y1abGSuYWgyhHaeKrl
7/cVTzOIuq2WNJKPJJqZEmu/fFNmjHAPYrUCBec5CHLPYlveJlpQZCxY6ykzChNs
mArSeX9ZTohAyajcENzcyEc9mqxynUWazMeYnoP4gDxlQAipqR4LQc+qh5BGI3af
ZWUUD0UmqhrI3XDIfVerto4m4Q4lc+t3Btp9tpbNhF0u+UciL+KwklcuWv0kmUdj
01Hn/4zQCcZdK7S5jfizxQCTd0k0K42tRD5O9xbst1KmIBu1EVXmI9dl2marRPM0
dZQ/AShUIlCuuYerIk4u963haSxnEJr4qTs6+01ULN44NDUGX2WPzQCpp/WH+euw
aCVojR5YWFIfJqyt5NrmwbozJ4QgfhplV3S4pLf3OSdqIRXX2o/PeuSwHKoU7wj0
+9jBg2KpCubhyfUbNMVFH4YJRo43bPiwTXYqWasHse72AHRqo7amyCMUSa1XRvCN
62qRibTKJgZRyQa3kl1du6zlVK4ekdHxl3sHzLHaACsQRT4WXbpUJngpBKxV0/S7
vkW4vpguiI2LBfktvFPBudfeTEECtHmpQgkYd/ADGG45/DgiZ+qc/a/83+b37sOl
bX42xPf8tUsRcqfAvLNbgabGA/tSSagGuwXCQuYDN9OZ7BwGsIyarqqUaqoBegaQ
tsRFr3U2EQaMkuMxXCvlAQEqmJXTsZ9DkLIYKZ+R27uHz6cEcA3xqto9PaDhFp94
t35lMNbLEH5wBDaolaD2p4yJJIBHJGD648pTVRM+dK1mYZJtwrgFQU3nYPrhKRCj
XIsTdMm+zawz9SZ8qz9LN6MkoHJcAc3ef65k7xeGEoQ3d5A2Ydsxj+/NS12/Lj+A
a8JqtWCh4mWmd+KN61vCZObioFgdfWeVdykL9esKLuvvdP4B51zDQHbAxTJ5ZA/Z
o4frc9aFoS3trGgYx6z7ny+r73oNu9xNyp5QfJ4QXAGmjpgiCwxuUA5Fz28JbyBU
j5xKUfrd9lzMi+dKYICc3sThAg/SqiE+C8h+hARBPtuNSZoFd7Kz56NKtoiAoe6k
1D4b3QPCT6IE0KEOeVaNlh6BZ48fmNMyYZ8T8xQ2oHWeDkJHMBMFK8cRJ37YYeoj
D1eULjuWDeHQ5VYfe3xPT7TumEH5BAAye6kYJxlJTXORn3c9sDyKpPZGc5r9QdSW
aoKkKxokGp5VebcSY4KUElhNwy57bDViP14Lr0AF5XY97Hb6ZOy1MlhNYYEpkfg1
rktVjf1v6cv+c8PY8+bHwT/C9NKNoiTFzKf0/feNwdJeG1LmS3YW3hw3I0XEPv7y
NQ2JzzzOeHZpq31N7Qm6zW2F6UeCKNtVmQjd8QTu3VvfcXy1pcvfkBQSH5mK6wql
PyQdl7U8tYj4vo8WYPuYJFhLlfLySDmr/FdH+nLjxYgqMHsN9Bhg0b71dVEyK0RQ
6jcsKKwLjBD55+FYdoBndXXigHmLyuCoVhIcRa7KKDvim4L7ZjPQvrJeAri3sQxl
xmk99Ile1YJcAnL6gLetZudmh7rgMtJgz3B1R+XuUV+gRSDx4vYGKXyfeJxWfHE8
ksuhlLv5i5EgrmIghMadFY6z9D8cAKfwgd0vLZt8C5PA/IMkSvUdaKOZQXWWBn1N
F44huFLn4G3NJpKJaNIbNzCu1wwzX+126/yrEYDPvnGC8kr/LhdBmS/meYL997Tm
yZgRTtafTAWLxTualowtpcAbtllwKDUyfTaOK17f00mRi+/t/FBeBUFZ5NI25yMa
PV2BcRqwqvSJ13vzEQKGsIEmqQtankXHUvX4mKbikQkOPuZCBbwlYeMqTk6zN5pe
ThAzvAjbYhxXh/TEeM+Z5/cGNbjl0Ln+ZgkcN+Ewt/DVqZg772psuOrlyiVqt0cN
bvXiTwa3Mwxq4wsHa5I3Q4NWbkc4PTCmws0kwf1rTrYdjYCqVxoZ8uCVAlFlZkzd
R50/qzVpZHZvVnw3NyhG636FpMZNhUbGpdRMgTAEuXNqAF27rHRlYuiw2JiUjvMN
AR71a+miQoDYaSLI1kbx16fZnGb5xZPNcj4ksQ+OdFeYus0GWevIMd2oFZmIUpDG
CgyT8HURv4udaeQtHftiF+ljoICmXrR9KJpj+0V500kknCFezdhdvL37Fp3/6UMt
6pwmooQTShLiv9VhtlBVAifkUU0n2nlrlxxEIkkg12T8Bn9ptIkUXz98w4VETt94
0rCVsUTc64EzHg6sLGMtBurMtV+nMTupCAlnBVRPq2dbIECn38UdWPsQE6AgAzU5
0/cQIFxMLHXlwSoSxZXOhnM/T9PMECaKEZCgS8QdFPwYQ1WcoEJh91Sf51no2FLT
N6ELsI+jPmhAIoO9QOMUUHbk1SVPTuJBmBMx3bbMMnlYWyWj0I3a7Ct0aIDWeaNe
q6cBbwpBuH2MdQ/YrlDlmzni+OLLohTZIcxVT8QQtY0Eja+ar0MSNH2MyqQSRzY6
r+mM/ysmTbF7KsPTwLQhm62IzCTgauKBaLU8efC2UKbOhWJzVtpLbfta9nRtJBuX
DTJOz3fL6rhlIo0oErDGY64ySMF0z9j1/Gw5VfUyxqLLoFFnCDw/sO0ddJtE4Pv1
v0vkcS0OxjYKMndbsu6I79mHUwL38ACB6SrZ/hId3u0Of4xdktgIRKZNcey0jOFN
jugE8TZvwzw+5yrvtyArqVCjOV29HI4K17YVSQjbA/XMe/blkkb5hxvWAs2fX5Rs
Ork6PDjvBdPOjUHAQw3wpGdewT6KqEWQLhKi4LZmAelke2svQ+laidY0gaTLxTTM
JH7+YNWegEkNTPiHWZhtoJW8b2zMS8aIW7ljhQPG8CdwTQLj7TieCJZZrahBrx1q
aRm7hxwhd/iQWiL8RH/k7i+BkN5+WKPqI+9poJCfz92iXD/yJa/7+OWJdouuer8N
rYTV3qwfl9US7YbJ6x+KtdwnIveF2cj2Lb8xt/UO3+32YhUYg1+5zzlhf9iNn05l
Przix/OGllINBt3T7vXu+aKTst4xya9sVj7shTuu5d2wIty0TaGTTwb0tFUMX3yO
NwUUN1njF/At7fD5Tiq6S+EPZscqeG4TvcdUNOp97yFxDcY2vd+Pn0Mky0Y99wYe
hJty3ZHR4BY8v/4mneUkFCtAmQ5/rdLH45YLLH3dQschZ6dbXB0ENtrB6Xt0bxoL
GuUjIO72mSMPK66gBTGjOytw5xIuWqb4wd8ZvrP0QNpjQ9Nd9cZExw06jO5+/TRL
AVPTkL4/UvJ9xyq0CXBPYqHdJRWrj7t4jlf+HyIVgxIDO8LZL0F0PaZVIBPnX/wE
WVrDM95w45NeDre/1Jc6Ztt6x/6/sxDMzyXcErsXr9sgh7M5mffBpDzrOOFJUlvx
wZ/yvEMmt12O7xj2mU+22g0lq6PCrXM32D6BAJQbOethJAJM8bsy2MLmvsrF3SM4
b5g5NHq2CZTXJA8oz0LdKCGtQSO+m/Ql51HnJw3YGmDkc9ERtRqOGIygsJRhaVAa
tzbqRJZ3j5RxRBWdN7TIDzpX4GYL8cjMV7ukhGhJ/JL8ytKxOzrpGcB9DiUZJfyg
p6oAsSgm8OipRwicnGtMTqBY64z3kEsJHSVCBfPclJoFYdwpVuvvAK1uQ2MOdLD0
BVhBbyIsfkrMYxABsMw5pqhht3PJAF9Bq6aFWev/9a12smQlAtaHxIjDbihVpJym
33u2NBk4UeTO+gBWKsTB1OywE4BYdk6sGQ8oBNIAL1WMT+GIkMA+YoB6Pq8BRiG0
6I8UDzybMrm+C9fkVHb3RJ+RfJPM/0ITwlZlCUYyJHxvkhxmYPkrpRmX8YB57EDm
dTwx/AabVFilcgnvKOKRzxCnaL4E3jMmbhKaMLXzBZc5RiV9awrQWSC7cavGAK4y
LNbFlLYvJllxzX51sukgF2f9RiX/cGwP5BjaQWdZ/aHp6irwTVho/gqllHD8QJdt
zPoHpdDNoua4b0u2lMjhGhPEfAfjMlLG4B50NgLMxNqm/CkpX2o1FNJiVft/jE2l
8Fq7ccAGy0d616YEK7pgzUrd/LvV/7a0VVbEphRQnmd5V4PAwaLB0i9Hl4p3QA4h
TQK5mm6WI7K8ripGyvjEZcGgxX3fuhwj5Mw7+MIWhthmY6ijRNBtKCmeaB7a1gG/
h++n0gnvacNWodSEvmv4WNbRhePIJBJcpdMW4y4cNnHuVmJEdfbVWU++OZo4bSAf
HCdDYXLMHNzS0UuFaFiO7a9lIhSQhpv8uY208Idn92kSTQ1eKLaFe3biDFV9+Umq
IE+W6RFoWKo8N6vEwLeBQ9+6KwwtYT9/CYCejLPCFNWp0lJX757pe0/zRdl/DmkM
q/jYb5Eqol6oD4lnEkyGdNKKgxXTX0mrbarJSa2+Yw7fr7JDLnrsq0Byn1AIYkY5
9Gf9GY6lUnhwXGVCtm21brOZyh9odisx3m9Oxlq6f5vD8jagCt4VbguZbgcV3Tvd
/ykexKGSXguu5X4CKE2W7VRg5iXOV7ZSVslmeCQ5Hag03yYpvItTWHdIwn5TEWGx
8Aurq5MDB3c7qEPkua2nMxSZyqtNaWAhpnoVPP7YXY3oKQqpvKTDJMCHVqeOIg3I
VX9tuJzhfYboS+2oKBlE3SwVekPffaTZrV8KwF3m3ADO8WUv0J5j4SFgSAmS8tGN
tGRv1zQ1ofJiguqpYHPBnLURMzj+k1mJ0QeZOEiNWZj5NxC5iXgmBGHF43tqgvd3
zN5H11FALFwOcaBb3BsImYd82xitVWGgScwnTqza5yCI4Ib8NYWnEoQFTnAZGIuL
Vj4iihDngec44qsXO5LKHQCjtPisqg3C1FPFPw5kojJtC6nAn685++560YGBqjzV
c+wI0rVw7AGFYL78qhuwf1ij9yJoQnrNupj+bO6EWuIJSxV5rDS/hTDT/V/dL43D
f3QonE0y/CAag0b4S701u8PWpLpzX3HnDnJwfEVQ2Ocgwgod1cq6jbfMcep3r/Xw
bobP2kNJaAcdxoOAw4snNxNEjYBogQKVeOnXuhmOrWxEGSovGQPsWlLjSi50ryo6
VoSHd8qjYZyobSLgF7TaJeX2iqxsczepqeqfU8MpF8epNaslCTOnfyfrek/kSaa6
xpOvsBRlhQFs+Amt/abutU8WC4f09f5lTCSNGF0xloJGEnaNqo4miIfXVJglfAxU
+CpS65/IIqoMGz+OUNTyxFVz1WA/ZP4bFqviiX/MVxM2fFYl0P83rQlT3uMs02bN
gBKYUoI2bqA+12J7xQuvaa6eypuem6VIzSV9WQd3We3BP2WhAcVO/x+2ieauakHt
0SBJGMgMHEcHW5YKXDtvTwap/gPDn4xTtHR9GiZtI8tH4NrSmdwBmeRZix48nhyg
RExgBfQ5D0rcYQAy6ihVSws6wgCZOi44j/m+kGt4M+pHAHNF7ABszH2A2TXHhq3f
i0wC3+A8XIPtXFcttKneiJRWHPYMlqh9CndfgJ6zHEtSW0YEQP2iz0NgmemPOWZd
9xACt2E66KnvqB5CmnmjUxvWPAoq54AxhsfQakF8OaRJmaN+154v8h2v0OQD6KiQ
/r9UC6SgwjTkJtBhvlEn87zXRNKqRPrIvAkSzY+9ss9dyArBFtVP4uTIPAd4y03y
/1c4rkA3mR2opJx45XjarEQCcUPjTid8bNbWcOnF1psZizl1nGbeFirEkVD/pnyv
u81lXM0iFoxqvbwXE7srIUiR+BiqFMIIm4O92zOH4qN/gT+t+pQ4zFAMQknAJo+x
kLtst9wWpBKJQF/gDLOVPHVtLaFCr59scbzhbzv9/SvW2Mdd6sMWNvKMUO9FCChf
y6hyXeS3VwocuavllSXqW6rdFkjlx5J5b+oiYmUpP3BXufjHIT9YOtmwW4pfGr4K
0ga1LT67Ved5JSu1F3iEVdOZ5hTf6eC4noFxuL7XGmmHxTqFD479ghMdiNuxTWLg
IEHEyvq3swW7Um5ujGBaiKbBY5AqZrQgI//lJHrNZSJmjRtdHF+LrypqLhUnuTLo
bNUMUGrBa/HGxLaTnzmp3aWoe+6zsjjFkXUKog3Dy7AiprKoBCeHQCvSDNQc5fHI
TP7ku6VEKzeyIBI/qrLD5vanmJFkfkgjEApR4AfrBwmEvIZbK0398Y8bgYa52yxE
AuGdZASfH3Yo7NSXfrN7+mmjqJTh2SPE2DCZK7xHCgtkj0vkY/4vsHyNLeWwgga4
yL9TzrT6L0GnmjzZaHaL32zjBtx788CNWEaIPOiLfJHSzfNHS4a+KqwMvn3L/txR
alWsJF/5kv36kboVnV0JU/jkVH6l4dhEGMFT6MBLKvgwYvVnULKLPwjyfmVHV79O
qszCV4seJWXmWoQOorh+mwRay7C8eJWXgeNMi+Fs1cS7icmJFDdHBrWWwtnWRU1s
y9gnaeHlMQd3qiVa7Yb8qgVl6R3qh9mM/VZzNYh5Xl1QZxxTEhQH2t8WM4cROxon
yyLVNCFENTPf4fJ9WuAzJjNulCmc8FaG2yeexhb0AJcBMiTbLrPISrQZEedTE/fb
AjAPEI3tV2YFfRIq/g52tgVSFVRzKcqOmxeRnJjoHY9yWAdulfm1D8ir1l2StiAo
ADzgByGOXx/IN9enDqGeE11gjlVEuYgHXmmVllj8LZAzI/79XAqIgXyrDMtHjndr
pSTkm/4uGH6h55tC8hUBmfvrXxPmv9j4YPArrQ9L484mmiG86OT/inmWYZunyA3/
C/NTHU8rVi/XFxEdyZZKrrQCcDbstY/ZXzDgacjYgLOKHA04elIwYXnhi+HFrAYY
Cwp6WEwep/R+JxzRxs6VDG+NAsbSpSfykE30QRxbx3oB0wJYDSzuw/J71bnfK0bi
oWysHSUObKHgwNyEhtEHXhiLy984Si8o5qcTuBE5WcAXNPsohUR4fgH8oHkLIeXt
lucLO8IZmU+1k2Iw8FGc12O3J8j6TuU5fC9ARnWN7xO8vmrsowFb7kMu45AVW0y+
E+qaHzz/Z30rC8DJ6JvbhA5fiDOllcKHiWhq5ygTJ0VcOUzBa+10dwSTc0cR48Zg
KBZvOZDI8nvYCzhm/HnoOHapvfol6vEsesmvdwX4npEiN4fYDLC4nFEVnZCbaW+M
xP9BSlOpTBrNuVD2cLyOOfNittFMENb2vybfj4aOW961Nqqrac05v7jnam+VlnPq
wr76BMkIN779E80RsDsO+zMMLXM2BIKvZWj0VKgKYpqdvBklGzJDTxU3IHqsA2tj
uJkhv3NwuxK7PAD0fHbE+dO4SeQ1ARDK1KK6p5CHoLJsZ61dgoYtFY/nIbCUWwV2
qsZw868i/wrhcHY6fX7IntVlAuhCnyXF2BunSCy4sWTNLvQbGtHo96x/7gKZACj/
XiilIyk1qybcS9JrEjtOdSbPry7FeMKrY3C8gi8/h/I0w3WENg5FL8o0ILt02BZq
4+8CBfmhzGH35t772VnxH9EIR2h/r+FpOZRY2RnoNTbnBfzyn3EGKwvBiDBOjFM9
Mwyg6Ti7IU9ftvQ6N+1i0CdvWpc0voaXdLFgi0L+kU/OZdtJRUgr9r3fUSYHV95d
jzCqPKFuwqvmGScZwEvB8QmiSP1qO+yo/Agg6GyeNikSWGbruShCopHm/Oa5R+iE
lNRgljnT2xGTlJr6GSiPBfVZ/pfb4sIZELO33W6E8bQ7R2tBh+QWmR82Pdf3ZUeG
4DBgGbqQwSGverdkHtrIbIJcm0ZQYHjtam7M64DNTnry1zbclBEpJB/6pwpBb65M
oWNZ/uKpQDsIl+TvHsUqAXc1c2pKqEjUjHpCeRWRjB3L/wqSNxAJNPd4/MENdY11
gCWXux+K8AVUOP1yHy/pIE7kyWR2RXoFxaCkGPFBpJKTjF/ndmQX8tAcYLncFGTO
zh9XXSRFrcteizclr6xEEpFvoP3E+HRi8llkDqjlH2q+Nmk80ffD5cQqh1K3MRz9
5rIp24OnU0Ik4oSmQ3xbC8bj3buhl4sDhr3cIDXQI9BXmGZ2qpElflcRAE6Au9Dh
Ywv2oR6NvqbQ3/wwR082iqgkTgk93+6eZig6iWzBMhJn5lJ/6nEjl3vg6+PwdjzR
25sRUELo/yTYFndqzEw0pSK8NE6FzqxEHBFTP4uOwrRZ1VmwCeL/VWye9dAk40MS
Y29GEsFBgBKXdmYffge4F8qrZjAC8O/zk4uMO5xGUHIzSQtAxCe2R5CZ31u6MJbq
xnQ14u9dntNrcHDpOXk1pwIhwlrN4l0M1xFBagqa7z/sN0I7k/lAr+lyKt2LE+vw
n9qPAGbjuyQjVF4Wg3cgFDq1EXLz3CNLAJm2vfeL+LpFLJrlynpWijEH2h734MHo
nd3BmfXYpN4vxYNhGrjpcW+OnmkNnEPowHD6qsMfJviykMSZo2XqB4s/AsFBRlqG
5OIWcdueZ/Vv2YZBapNlKXTpdvwf20EklvQFncxvRfFaLJDkBQOJYervH5HviY/1
4qfanha4NxLJ491AePULweDB7AJKNomN363GGZERWfYrySa2DZfry7QcctbPqBkz
13H8Rl7V50yxdvg7JtT5wLhXoQs9fMjJnvNhcBEm3rjZDrQUuhpsRVl8Tofz1W8V
6L3EQ98a2wuiSQ13EZu8xSM9Ez7PEQBC1rLZX1GznUUq8pZXc0uhEWTcfveCFRfA
VzuCFo/hw/54IxTcUy+NRnfGPAYKpxJ2okSJ3UeeS8Gf3Swz/F7hPKINXE8XqJ6y
JTBixMn+HmqcyED3ePmA0mzztlq9juBavpOOPJ2d4M0+ipxFCCCKYzvWYPyPVag0
XSv9kZgLkpC1kk6UuhzV6NJPVrs265pabBSIPLzBqutTHsLWDVdP9r4ToWjp3QL0
clG1PBvDtM3dFtzpqqp9KSOdB4njNgkVESKr7827CFC9xQuleTwLlXRyicFR4j9X
dJNzPn18ZFI9QWnjBLCiLNGRJfv4yFGSSwPziGlPU7gbAJbMU7/xENgbkhndFVpY
hY8OISo12hWKLhRC76mhtzgkp+hNm/7SuFy1iV2bJSLg7zt7X0VOoYd8dqC2s3Kf
aqYZmt7Djqs+5fSOsY/McqFOhlfQ62XQ51j+ubk8oau3jp9SJFRHNn/eynafAdEN
QLoAtMs8VO2KF27ZgVrjYgDtPalkNSMvD2Lsyw/InQ3TlXCsh2rbnjWtEPVDlwCI
t78u/BuaLexbjZJLfkZZzM9xEQ+PNChYbiJoeWpQHiTX9Ln4ByEemu2eAG+xFfXl
S7+/czZOq/yGn7yRQrQGuWpIQ6v2ntVDmjHixZgBsbu3yBL1eIQUaxs08G2uD91m
r3jm/1H+vaVYws/goNQ8W3pHihrru0ESrkgoSBK2Q9beQckzVLnVewjBijjOfxsm
uNlV82rrz360yv/xDyMIVY1vy0Yahif3smxgjFOuWFuSE10h/J5K7d5eJH1Vkv4h
Gpk+34oTO9L0Hj85cV1Mg0FkQsA4DSOCoFm+7japSFHb3iRov9Yadv7VvL+Lh198
5sNX2+pCS07hS2ZYko1yJrFAye11HdYgWbWCqhQ0jj4nFdGOuGuOZZ31zkBzdp20
ERC4fq1g3N49eoB6524Yhl9Jf4uJUUGBTJkOK6mAAMgxCytuihLlUgFNw/IYgcj8
EqAcoDUe27R9MZsTGjJH4jUrTUkLgeVermr9AQ6gTjC+DVOm3+XqLnzfVTUTk0OK
E+ryORRPc8ujmSwA6CLbbr50IPulrTa+w9KBxMaJCW+Y3qsQywBfxTHsqNWR9qSK
oKiO8fRLSwBe96FlQH6jMTFyAUMEPNcsqD/MWMBIyjrIzykunU/yHtpl6LpZm1eO
xERZgHGAaxzqFZ8KwRiCivx6snGQK9akzIv+E8h4GMSgEnLsIt3b9tlBUvAWxSD9
LF3Au95JqQjadO1EM2/oMs4yb4doKPGBDDcZ2jTPSmLm1x7nRTlwAhV01EVurxTG
s1LExL4V/Vh1f2jL3+dwppwGg4psKWsnApYf4m4QscqrwoRCsaeUzzt1yp48647A
BwOT1qsg0II9CholM5qUiObJLMmhydasgkNVohb2wxGurdp20yy0pRTn8ElmMoP9
Mf6VJbGM6EpNDm09uu0orA0i3uaz7BjrNKYcrxICJZoa8NwM1SF3L2oi7x8tYoNR
XjzjPjS9IzX8uXPC5fOwXD24tieZHd/a3zgektKX6OuD1Sycf1zUrEyWdGHX4Ncp
8ED/NiaVeW/8+dPQkJiNkVg7nMIBZTqIae6fGB2aro0cyt/tzxUVLirYvmnmQzKA
I4opmRZXdde6D8SiAGMDEhzkFW/U10vjTXlWNE1I7+OtLSLCFhgAyRb1UhTAVZZP
C1chJK4iY1xvssowQxUvgi7MSnI0fZ2nbEbHFSRpAElIBcNvhvgyzz+zRcnUoWQn
z1tPzhVLc4WHxG+Wzee67KM9TnaIFi3rUJ2hKR57wKqzo/9b/LWhjbigi+lFY0ht
n4Ejyp1NZv79UeQhgeespS/yC1if5IMRHocikmQ8cgEj6hZXc6SGGrcAtrGOMfsY
VmKOlcjFu8p0bMxfo/4+og3ASCyJD2F0xl8gHmwxJjSkqW29emkWsUpOAlTjF+ey
3FaYRBV1M6IJO6XSAtx2IsbhaVWE9zxDyiy5y7BYvJzyPKF5Oi6QyU7OvPdW1qfD
eYotSpcWifG30kmR3auP3Y6vdRNHSPdhC85tYJonmpUUDOHsUWp2plDcYS4V6bHt
uA7xNiG8l8H4LLx39sgTEBMi0e80dct75OiijVJO6pjd5sCdDwmV8RquE6apFMyo
1fbDyvyxyubN0RLbcake4tYHsYoT1jtn5ccIqF2TUglza1nnMyKv/HGQx/2XBlw+
oFDVWrc7a6FotYNot0eQBra69RP305LogAn/FFbxKN6DJqyCL2MaVubTuct9+bm3
8ydR0m9Uvx6Xm+07N5mycQqUEyChQZSFgfEGF/fVCWHsqKKYZ8h6wGbVcKx07s+A
X076g+dIu3sdUWrb2KEGEnruEvPwc7nbb+SIQJbUSQayIoLBbULLtNcbO3h4G/AR
DXo4TxIe1clOOZ4nidpPXLNaymlhHFc7gmnb7YG7KRFLUgUBmAJHCL1a5bkv9g2r
FqoMcO18TJ4IwTd3XPt6V5A2dWZNF1cShcJtPS9E5Ce/AXYm+OTBU6UUMsG17wcx
Lw5zSU0czwOCul3TS3pRqBn+3afelVCcgFxWXFidByagxFEkwGPg2YTUPk3kCqGa
HSPB9ybCn4R59J79JvwyKe8YX/lAnZHvj8rg9sjNbAE8Q8KwaC0FH+PfHYpEJBB7
xGNm/UzElMOyHwrjN+Rke95DN3Gu5Kjj1ucQkvsoO5Dl0wlrbJYApbKPLOZAhpet
aGOEiPIHdyVT/sPx5ZseFGNvs9PgYR/tWifBpFkQcz9SkGFB7CW7zwn/YXVMx/jm
f2ZCJwvwv/faSrRWyQ7j0W2TzB1Vm7TUpyWGExreKEHy1JdxPvWyppV1klcTiEVp
VYnJ2VjJ2NDWN9NCfC74uundGpMAfAG48XEhUPCv9TJcZPVEsTjKMhhNyJsNlWyj
bKAGiIazUjEa86a2pVFO+G24W+Y3ZPtfZ0+H3MOAiUFJ9hIJvCRifl9pz8mBIIV2
gQUyAobkb/B6SKvQtIEdyIDCj8A/z2x7NHm3yZZC+LbxPl1l084lJ9b4opzpa1h5
U4Nm+oruz8mUsAeUzEpXDlnfa168eLeaLUiXcpo12TmFeVI2X/3UYvuOKtWFSGY4
vQ2K236yUjo0W+mbGNSQOu9uXaDlSp/qqnuTX3o7xOGgnnYz0yy49DxKtLo64Bgu
Rv9JmF8Cbk6weH5nxzeBpo+Vbqu6n9u/l2xbyyfh0LDIkZ6bBamMQ4IVEgrRoIlK
K7TLqzcpY/bL5IHfJjzyj/rp/8cMK7hr2QwQridl6StbLMhA3zSXftjDH5GWGOGL
jyJBbKgiB0qDXx1l1bNtHk6jsgHW8sj1N2Ry3U/LvmFMAaQ/MmP4w8ar/QurAMmZ
ApN6o/AxlcwK8q2L91wuLAuwo/C7hkYPlZvB+o5BszQRA6ddX5OKBOmBzuMTQLGx
Y99PwsTXpGvsmQdPHTE6I0ylSSAAb95ZZcN6TYb8nP8+i4WRZTzHgrytgGu22epu
OXvvOfYfBRHfxuOV95gsBJ0XxA2GWfJZCp09/H5uy+dlqQu3CvoEd7QpiZ0TIDPH
ARXiac/a+TDW4XuaVg+PRs+O8yK8pQukXP/aOglYEUHvE/0uO/4IlFNF6VM5hJgY
C6sBXPgStEBhwplOQAhf4rcJYNIGoqULAJf98EZj4yfuKZPSiRd3679unMO2DkES
IkF4PBvmh8mERvfvE0jyEtX1M0Xf3oSUfWftVI3nRlGZrBL5qiRiAnPwdXW6JZIG
pFh/5JIjyu4e2CASDJ7vt5aaO/oXm7/dwzO0w5DBdMbW1Z8ToM4oK27YLwiUWq30
huvoTCFa9IMzz9rSF4LiPksT8C0YYSPPioZ/sbtkTVVwxMUSV87t7S26OXlbJxOV
GQJ6piJevsVzAV6swUOzsWlqWBnXRdkg+M77fk/e40idShOqaUTjchFkQfH67c6w
sSmVnPIHWWJ0DBLUvoozVFWMkZgZNudJO0upKCPwjgnZwdUKnisnemE6UPA6Ssd5
1AYA6FWP7V+LPDO41Ilz4O/ovVgYrdu1Ft13KWlFu1ajc3gdVRdCqcnpUjfC2EWo
tQNOdRzGmM+D+acXvf+8TKd1nOkI9xfILjssDaFK1DBezQNa/UMPkSq01YQaO+2Q
kpXLsvFPJ1yRRXLQHOd3Z9apyNu575iKkjBDE96r+R+iKPhcpRR28a07B7sRTt1x
1aH8ofDPepALE9AySWFKoMuNgnmLkoFZktDiQPGlSxsKF7Ba4TPze86gvwohuq9A
+0Oyix7WhhfRRLNnqJswe0kMV9svinIvcU/6941n1fW5PbRo+EK7Oc7g8a3+o7nr
EWEN+lfEsY157A5RPTAGC7cXmdl14dnCptkqRMvEJwzprcd9NLRQH8TXOczrGNY1
jF/U1xd6Cuj6Qqkm/cBwemWUpxLtAkI5Ofi/CoXHCxpKGHIpXZLVYgOFaIbBWPZR
z1qUrf4NtyYBhDFbAXsth9LcB8yxXJUgeWQS7VXHMjqL6tey//dL+H5ApzNCuY7H
MPrmfWBjS01pGvKEIN7Lx3GvvTxvju6QyBc5tvjOgr4wfXydGswx6Ain54cibLU2
8QPV03b6Acb++Ow7qfipYjCDw4JY2NjRWMPa/tXt4dVA/6mniIbCKs5m9snOU6+v
CtMBqCd3/sDAHRyG3Yafmv/bUc2ZbQ6GAJ42O3YcYN3RUeZsxirfJTzZfvdR5l4h
vHDAYd0HiUAZ/d4wjkALKs3Xn5WmFqAjfGYguWS9qAluPCCV1dZwZ4jnYQTJTJS5
2HzI6t3pbpPK7lETWRq/2JaYVUrQ1kpMH38sWobg08QEp3AWKOr5VRuwCrKvinWa
uMTRouAel7hhpXMCypqxM4myTuKOKjz5SUGUNirkQ2QbTq37JBUQ93/OG0jiDbVK
99XK78e0frX+BKgyBrtTo5JxuXD1COmAYIX49xlFjYDhjIkF8AqJmM64MWT39kLj
iWgab7/tU9djsC6Pv6pJRBUZyS/VA9i2o1Q+3IlZPzm6UKl2QpdqUJrhF75az7MB
RzJ6YNC+CN+havuM9hODSqHeDmTR14FaDay08svGYuSglPzA4rYIGck1+tYvm7p7
NL7o+ihcCw3LlLZVTbBud/oIxjqUUy5214D74gCmRhwqMqigJ0TR4lpE/OswzShf
JBuYy9j08OT1q63DGuaqnPmqCnthlaeaWyFOjN2KE0FcWEcpA7RMMhakp1iTkg4u
+6K6+3Q0LY8fF13XtM3swqliUA9+g/g5d+vEZ0hu7EJoBNTclb87jfBOs3E8EW+d
uak4mHpQu9Wfeu85qUyfit3tMxDT6nYEgFivD39z/jJJuVPeGSVbuEUORbE1rUrV
//eoeeoLpNLqY/RbG/heEKHwG828hYHB7H6VOsir7ekT4uaQlwlx2kkiMwF7XD3n
fGUoF6EnOG8/7N5SiA9vMaeNLZsMn3n7Lt7YfNoT/UyBdRzmGSlq2u7eTgaFX42W
o7JbR79h0kSgfyQAaGUqyOj3ShnONVIgeRXHTB6RvAS0ZdHdfKmhi+Whyvft0rzk
bFtwknpXWJk72XIDXexC0vWXeSWslXhscmhuHe8uRFseizr4V8rhpMcejoWT+vr+
SPslIgxTes7lRevlStb10OT62rmokha9pA8NLKvkb/P8EMtoyzYRh35VoCcp5IFm
ai+5+PAEUlmcI3z/sA1dJ5x3yWCDl1CxYrO8Gla0vgGjVwL9Me0FHdjvd5MfitrI
2aTdvTVu21pnRX/NNWsNmS9vxC4VKpQE27yfEqGz8f+L4UWFrIldIO/XvxixPjQp
2BnYkYCmRcpHQkntB2YLVA3OIkYoYZ4sghvrRPht9QpVLxPmkqW5y4A5KnBW4XHG
Y1XZ4RpnceHY2x6ZI6mmv4bz7kiUTGua1t8H4y1LxmoTB43C7akMVXTgON+ry/GZ
uYPH92R/0nGg5ZuC/QiNSgtFXPTy2CkmiBRfbr+ZV+M/wacWmI0hLFwSMiMKgcqZ
gx5N9K5hw2AN8S0ivIwDESC04Sq5xlVyw2Hvw6Q9hDI6uW4S3Gq+FlHF8QBN59x5
95t+wYxpZQFVciSSR479yJYceJXe3Ukvi4ohWMo+OuPXDtZWXxHTihcFKI1hj8V4
Hq1/qRH8mpMfn47W5roONiL668tJRV1ae/XK4Q+WyvbhZeF5+Sz2GkypgiVSwpTz
0hP8umxpv+jPgtzp4LS+iLtBJ8AcjWN5z0fmzHnmx+pwMQJB0A/aIpz3nJC0gFog
LCf0qa2q9M6reXXQvj1N1G4q+Dy/DqvM3VKaCq36vE308+6g/SXdAA34baorCjP7
fC19jLlEmrup9hFWHxERR+n/P1ly7BVxmUU+0/vf7L4ptTlWksDnwz5VV1qJO731
8shM/oj3pnL7SpbnTGXUdPm2m4w4cbzavziE2vGuGekJTNCqYSW+T2QLUgJA+dQ8
1QsM/ReDIt+VGsLrKDIKQZSgNz/cvhfi8wjZNr3zT3DTMiR42SCPp3Ma1Z6GTFzY
BQTChCvv6/n1TUE68RhqOlX8uOj6g/KR0gr/0NxpiK7PXhrgPYjQlUUKQ7UZWU84
soApfH1qs8+6Nvigtc/8OMlJx9+V2eIDsdcFW1IjgtusOQdQDSnFoeEBDabETy/O
FLWWfjDZhKKLIJUBDosoqEYL4/q05SfbyItHtjBhIUN8vlYCXEYcrtRQHRIIkvay
8e5xsaqwMorm5W/PHCfLanWK3ZuUS4QmwRZJaZBf9mBwfHDl8JEjhbF5V1f8ZRhP
33dazTfd9a+yGQJcEchgcZ9w852N/392amBVW/9dcq8k75UpDVlwi3bWCk5TeYmI
dIdCjS6gdiAjltRWrUQNd+m0tFXOoF2JKKFjjlmfxtfJoacUD21bfXDvHcoJOoIO
Nv8/TljCK/WZyNZQwnvEDib3Jv0TewDfWTdgAah1tE9KTx1RIQ2MflGRNmvPXCM7
u8/ulwpYtK3ljikB6ehoEB8GaWkWqMA9cqKMAfFAMWdqdv9Qe6lRhLwriieSf6Hx
ytAYvT9KyUoM296ni/bYNX0szF7LyTLlmZEf6y9uuTEAPL6038y4BwqBYStOzZ3k
fVnwrDl+4zB/a6cv34HW+LsbYS/xC6nMYebiS1V7uW9AHrhM27fZh3CGY3WzmGWE
VbXsvgJifP1VDYe64kq36FBQMmYrNXVGN/ZJfttnlnPMYnEk+BKU+3jUXB+H6yyt
HLnBydBjnBx7zh6dx34vvM48JBAQWGsRSWRmbUtVNpjbBKx3xYtp7516YTkCBFpR
ZXAFYkIzPSXzWMA3RQidOdOrCYFmXevfinjubAd6eM04HxpEKgvzChyl8ktHJmPb
iAv8jntO2F9N/qOhb0X8Mtq/6Mw2dYbUslJH3zUN6tvAF7ExnmPcjWuDUFJt/rRX
DHCH6bZ/gATfWN2/LQGBiSBDR+Y7pyJF3h7DDf2gDNJVCirFNuMOTHi5dWbcnGx5
w7jP6Bix4Q6ZHn67+JBHawSI8jGFDhRuPcY6qVY5l6yNJncxAwwnh65QLOwRLN1V
CE6VzimM+DFHr/KG55a2dsCASdlxwGEzJox5IRerLNtSnlJwKm/+KEkGiluO6XHE
V9RVXI08Fiw8wbopba0t0hAL95SykxG4WYq/+vawqEvsLQA98Esigtrl4LbMlZC5
eqAUrh5yA9a71CVnS4mCLySE30yddb3ljRpse2MOLhVcC4V+xnZ84lySJhVRaZAK
1YIPQzQOF4Cr8PbDLmcKvj2iS647llqCbRFojsfGitaYcYt5rifTAT8KvbZE6fYX
6rK12nQUDW3gfUlXhmPa15A/D7Lo4Q7NnDyf4F4CkEet1LnupEJRLBFu87qCXC6e
4uXCZJcW/Zyzo+A40DQrbzHO1mEYA3q6w10sGvDCdYTqM7nSjYoVhBCpkwZj3jor
SXdz5v6lKesXcRAnYwkBh4RRcekHDEYABa+qxSNPrDRys6CtPBUfoKyC3MFEVd7F
1L2xZcvVFrnutuK5mRQLh/GwJ9SkOxjdq+7RrRw+gZW3FxF7JJrsHSSF7vctisEr
XtOYH9VxkAxtVvg2LyZcTOUp7JCZHJ533kpRywiJlEY6CyMfu/j/gd4z6rr1ISsm
FadG5P3gHRdRHYCkex2b3CKJ12WKTHESAYFg2m/km6pnT+ifkjeKLEGJpZ1M7VYZ
/KZZqTI9Vst8VAMgTqQGCyjZC3EYgLiNHVD8j0xKnvG8e0AeTD2/EVoTbhz6NIvC
K/DIYsIU32jwFY06XZHVoYTE0osMGOh/eNtW2npZoscwWPe7McZTyS8ToZZ79WYd
0qWGlUYgksZBMZpB/Tha23sXbkZgcub/qA/tY5Mkg/B8556xCXjr15aFYyrgLx3G
sdK2R16VRZqpuig7p1wGEcYkFGTiQ1/9LIFmbv9abjdZMpFPsxssvQMMhf7W+D84
buUn5584KLKRE9trKZL0RInIXXZ6xWz3UUf6/OAEJt6JAADWopq/oygMbfZZZp2H
7LFY9oRNDl+BLGHF3jolElLzfhadokYAL/sl6qnhrPkcAz7nOqi7CM9ySPwKlVKi
628QEBid8nkmBDeYTxTaqeCRofQ9+3JAcKJdL1tvtgzwKYBY77i77Cx9xq7GYzWF
xd5mnkIjL50BPd7pHRevb5JOTY3IRA055MMksl/vbuqjbl2tctKP3RTyMdq4nhjM
7VBkfePVvw8NXgto3QjDNHxxBNiqvY/NmBnlH0E1lC/yBJ83v3PWMUWQTlyIEvDa
QgVAXoLwxGjFK/yaSBt34BUVL7Lqmknt+1V1is6W62aTCuNeQepr0S4+J6+0aac6
W2WCjjhfQDbcF1zwY41ne+SUKidafWB1xAgTDhRvwngI/N/6sgIFwaPcMozjm9M1
Is/p6Diltsf8KM876+iWblUmsbmhSJDM7Mo/kspwoW9OaGvW5kyrrZ9UuJTeL7Up
5svjTyO8oYq2tiFUoHKr6EDOLM3Wix+SBetc+r6VfqHosMb9eFTURUGfASC3WTHf
i1EwkmH42VGVVbSlylrHb98rpExY37CZhZnW4DZixPW2v9O0KElB14jwhH+/uBOz
BY/XoINq4JgKV+ZE+SxaWUSM4m3hIqQxukMYu6cGawspSrXOaEt9qkNZGf6J/5tI
mUiim9xicwOyvz/TvN0RwGucn0y9XjApZXT97duvujWjSkubCSiwJF7nNZyzDZxF
wR3cCW1TMetEwDI/zZ/INHN7lKP/GZwLx0Hkfc9VcZSJZszSsUlCUcDjiQhnB+Dk
XUGuahVyvHuwE0QbTPsEMRoWE/Xww4YW5CI70f/9dEpCyNwUtYflz2/k8z3vykEw
cRwPRKlmqULdLsG2vNIaOHLaJp+rl1PA4xm6QCVDOrnmxiGoHp3zekf9hNKOLgIK
9X+4Nd/f80bWT87BDuh7TX8tqqqbUNNcEUxijykFjam8Ap5lt6xejK5gBXvuH9EY
eG/boR4jaaEk3dgUZFaOrmn2sMYb4js9s66957vFbtNI2pF1IDRBITTS5wWrlNSG
JWw0EZz8A/9z49BoRrfh6nB1rb0I7FPLK5ppX9BlqhhFGTZTyv6qxg+PfkvpFd61
tpp2eGxL4UX6lgilyfVTjwnrkqT6PwsTNCLkJFEVpeziKvNcVbpQfJHTbJGmHVGK
bK29J+MbFBI8m9zr4oASrHAcRK70tP/03Z7YLXSgKb8IOP+BzrkH66SKV5loyjn1
3gF2OjGuogq57zaeOSvqx/CS21PS/GWHni8jQD8+KXVOiHQ8tG29XlaYFEVOsrm5
6jDKZd3rAUgQ2B16l5ZFv1nz/d1n1QXLLZaCzGmQUBJ3EPMQNZIXPkpRPW31LHkG
TVlpPcj2SlGh1KK0IipFtmFq8SkJhKIDHV3iz+p10bHq91SzuSiqRX5MMSQSQ9L9
81czXu4vdTx2HlnQxy0GDvpoE3dsqALy8s+7GOl54tYQR02tgvj3v7SOFju3xHXV
Ez+NdxdWrcHA9+zPgGIFcHLhN+nlCXNTYRSJi59ncKcj49gEYKftwBIi2xVyAY4X
fa3R+dAe8EyOyGboQqg23rIvmb27M2YxzqbP8bNFY563H4d56293u9X+23pRmBoO
GHTPKalooujothSD8b5j/CHHmUYv2Xy9whe5Zz8I6XH11ty0MvKip1aXAmX8zart
BSe5VbLol6jWGfURordlkb3IaNkJN1uUlKveBnuBQZmSWq087xm9YbBpqmGpEtI/
B9gLkc0/yo7KMnFzwyTvSw+Y2GNn+ynP/53fzT8YAfgfcLoh83F/C8+JrorEPALE
GHA/6ZAV4vlLgX7cvJFvEiFrozb/JYkLEo2j5qnLqbGNA7ivLOpSIZkxXNvEId+X
EQHSEA0hHGSE3Kh2mozQaK6GQl84Vro6/ARF12NxN+JuQWRVTfaASBsr6zIckidL
npnXuJTWef28bv7Ko56+hp6y70lMsMeQj27kVnz5doivdooIGdUX9Yk20oxL4+jp
1DFX9gegKRcN2rkSwQWK0NHnV9ZnmD1fwp89X8sKry4kfiNVh2uHz0UYhFvfdX0n
46EYpQ57+jnQu+uz02wCN+JWe+tQrnCEAa9VbZaaFnL0/2r9CS7pJCLo5Jiix4fo
QHCsnqZyTQdqBiEmyMl2Nbi37+B1YoqiP7ueZGF5kxoVJ1bM+VdOBHwAVLW0k0rO
uRgpbxq83faH9IVLYA2oN1s/+UoWA8NTcqPuQ/+0tyOAyIPJwCHoJwl0dGPjePaF
JjtyttZIs/2Vyi4Awpx9cWNWd2gw912ZRcpEs+6+LwXwjEGyt5ul6ZnN4pf5CD+a
Ani8E4kWkAbms07ME8UFbaDc6nuulb1raB8IV0boja+aGniz5wmvi+KR0gr9JqrS
HNzEi5A22vGzMCAK77RcR9HB6f11T3fUhfMSdt32huLKKK6y8OBRQFqPguj540va
nO6K9xHbo07+VRPukjwUA2b8k099FGthAUxni2ZOOsUzvcQJ2fPdCYgBPXcEjyjJ
tlR1h8M0prkmDqaWe+dpU3ZSY7G7QdxFvzZlhl/FNuhmQMpAeC4aDHrQ6i63iPId
vTtvThByMhdeTiu5GyiV4h/DPbjlaICsr9qTXfk4NhV8Rm06FnrY0tK1yeUN5ZBa
z+Q2Klb8+cEKLdmMOLLZeQqGyQ9l3be1OHoNL1adsSoum+BDzJg5KNfOuttN5ylM
5DEbJy4WQFW/X/k0QnHWHs5qFUrLmbmwpnTaLXDaR29Gi37LnphMflydfMjLmaeW
2TU3kDtpJVjrh7lXF/L+czqF9HWF/FOfqzfFK35R+rn+/L7n4K2mEIWHO01ZRgl/
N8bxBX1N5T0LvSvqPRatd6cJfaeLuq86h56VwRX2jHGOdsRcUAB86kPCkuWLljDZ
1gYkzRos+RjiNFdQMsN1h0rAAQhdvShHCIeR5Zh6ELtiFaJGR6UZwVrFvNWIfWA0
9jmPe2Go8rcxn+WSB0q1fmW50vnLCEz/RoDPGVU2+pV/qAlUvcLUbQavD83Im4bA
yr2palu6URAMRxJQxBrAMXqpXkI/s7CDTLLc9tr0Vn/sL+qIOgfPp6Fc8oPA0nqG
+sY9I2JQI4DkNWWg5CE1mwLj1dbLVcv9R6eccWenjrnGzJlHBxYiD0YgKh+a+GNc
gaAc9wWGRKr7vK1W3XYIAzD269B4W06vd65wnq7F9d92Tedh6CAFADbrrLKaqMlk
JE26e7JCQ6NU3b6w5ao6sVTci24wt0tJRJkQiIMQvo7+R5p90sHG0gcBjp4diVEa
E8hJKI1OGdyroRpFewMv3MPZ2RU7l0sj8VjD82nz7EtxkMyI9CkjcGNHl5XyiDt/
if3vtrEA9VWk3ZS3fx+nWG1mCVRpE+fS9JWXLjh7tNiYmbJJjxyYUsxN5s+4TnAz
tgQa/9PiFJb3qCeo3xIgwFvaztH4eo7ZBLo/q8UK4ccNNuyAwiateZiJR8xAm9N6
lCogKrO/PjfEM07jl77hlaIZgXBKUBpoZWcBUPpAVAFy7bcdVWLv8PaQ7VA+aF5l
Div8A/0KY5+5yQjXe+C6nXGrHPMm0+ZFIY6pxb3n6PvOzw2eT/bgehk/xqP/AEVB
DmPgACES0cvmyT9UcNevdGNWgEvYwIhdgGmBxMKYUl+H6rci4da84p1WWmJmQhGT
T9O7OqJqDoLNE+iTDhp4eStinVW4gORbKZFED2D0jxr9/73XZib9TUiHG4MEqckG
8+NnQrIbR2CjZxzj9nimFBR8yFOVoYiD4XJFPX5N9qAOHdfLK3r6QmKu0h1ZSlXy
NqWiTVUeBbd4z3ZZcpRXwmvtUABlA8RHt7voCU/hR8HE1l+AP2eoS6HKwrRV8DNI
oT9dBdG8QQskQ5hUgtlo0lDbmWSdlROFb8Rx8CJ2JKSQIIBsal1FSS9A6DGpQ1Wr
366sIaNBdlxN+PPzQ6z9g1SvEMfNftv4tfGdNT59pzeT2DHbUVvjTfKTdEA30t9H
DnO9FOj7Uu+TaoYblZa39ZE/CdnbMJ42N3pRcKAr97imNrqU6K+3n4VSoavRZB1V
BaHU96mhZCn5IEdnHSTNvUh6AMa9sI/UA39BYVBko7t00N8bnN4r9aTNUxS/Y+qN
2CjzeU6r3I7QVk+gfa2jCSk7iVb4MRnaMi5MoWzxi4/kKvn3gBrsrmGK84Xs6gnQ
q3q2LO0Msn5vyEiKohC8eNOiMKC4+hvCxFdsouBcSjdRBmXk2czsRYrgNZ0Gpo7D
MOJSfrcaKzck8W3Q3Fm/l/mPPT4A0zl0SCo15zznuYUvcY+7NOVcWt7VVJUI87Kc
QbXjKpBZoe1K049DAG4WD9NZdG1MSBZlHWlr0BtV7AAiJMWrfDw6ltorrgRbpgdB
82siPwXter5P7lk9uU8JiDHa92iWyHeah6LV0DnYHjT5e8333c9WwBb+aWF+NDE1
hccL7G6rrtuUIDMazbnRSQM3MrwPaXh8zfJgcqJOfO7ia4dnLCzn/PQn0ihlCEXy
L0VIY56UTQwiFI9wscsfVJb7o0cMzMXt6zvOGmIYD/zuatRtq8Lv+XZsMYIfYjcq
SOQ4RibJ3Uj86Ae22t3GNwdlnW2I2DX/lGOJEowReEuGfzg7w+zNurPErkb9VslV
+CmokDx+kOIds5to4LeJ51MCf2isuVkVvDzJ0zhCHObZHKjfSdBEg9dx7psYMQn/
Z/enjxH4XR0V0BWB39zC1WQSwB8AzSGEGmroG3LCAjQn+nO55AcV3caPejnp3i9p
X9OIgpkW9LV7lXH4o2/fz38bek/Nv1sMpcPfL+xJSjsNV4/9BhYkh+nQVSajst5g
W2RmgZkcLgR0oeUY+KU8D1R117QTEdNw9kSsUois+KFP2rnQS/deTpxqbJKfpYX5
BBpCpwLStrTaKYRnGYkXXx8GzH4VGE9/LrMj6zrXsXiMI2/Cjp73hyviU3lkctHa
1EBjvmL6guSzxzVz0ZhYxOt1bd+A/LG59D+cTiGEes643iogCvhCXR2P6gthj5tY
NO6R64Ey3ghmicOeu+Imdng5KYAyFiytBbgWTOnoKaCIRWnUJcZRqHYbX9r6DpOu
RcVZ+0GJS5hPwtng7b8MmTASB32Zgb/KC1SMXDqAzIx8xgGdaUBRzPODg1IauITE
HNmkSYfKZrPTTRso28+znOWrrjc2HXHgGxoibrPhhmlYr2Ik0oTY8dILTUyfAJ5L
iXWKqLmrFrYWXiqf6JNUqwPGGPH5/hUeLF+PDETJeBPvlWGqI3AeY5PSO6zhlDgX
qkC+LvjmKAIBp4xa0CxPRoQ/1X/4gRar14er7wsTpMcPS7rEv7/izaXSjw09e3tW
4hL2DkTY/ptpn006hWI/JSM8QwE5RbkRq2DCIucp6EY1Nb1EzxcbGLN8XJ2+xYJc
rwM4uv2FoU3OnFFFOJOHgs6agBORVEKigZtjbRIvlsBZbXCP7tl5NqjXvGfkihl7
0CWUYUShnUbaPRDvDwwvy3vbK7wz/reXaDVRwMI7lQczlq0A5brr7JGkVn4VUkwU
+Ij9FSeJ1S/io7YeyDeJm3USorZpWK4dN+olsC5t8QXphONPkg2jIGW4pcv9P2BE
RvASvx8hcqf+1fSKqiA9+6JzEDD7W/8x69TrzOmsQTS26LMxIjCn4cIK+BjLNNEU
3o337fPXs//pRyt1RKJA0UXwNKCRM2tTY5dj1LVb1aM5oPhSReLd8Q+RWP16GR9G
lU9KDxAOhIM32VJGRcsatMZsVy6+WyCfebYAQLW6Y6Wte+qPK0an/770cmRP+hH9
ftVJmM6vv0amzJKJBZWZjLsZFlC9X6s5/pB3eeMSKWwhO/xais8TnfKYGy2I4YkW
jzBDpot47KWYj+UvVXgTfC9v1gnTApEBITs+Kt6TTHpQd7IAlaOzhrQhZ89/FweY
AzBSFidv+SnKeD6WuKsdCoYevy50iQVRRBYngO70cjcMb6QGgAGS7sPSilIJMuTP
b/1reEjxu92mWEM55sZN8IpqmYSgP0FadqWj7wtm57E0MoqF0BSfN/ZcpzsKMBla
pwX4HTE5cDQ9Xkd0nUZrVrs06rAKdQjyhDEDo5NMhM7WTxUg1mp8RmV1sOW0wKB8
aoH1I98/28n/FdPosbA6LArFqd37PhuMWnBvssNOdashc57o482piOKPyhOsapeJ
Zy134tN/MifwmLce9IpavR4llQiO5H3OZJYeLxnl0viNZtUjxRW/LJEQfqq1WRWy
2MU+tCK0NHbjWxgKONKPnwRvdf2/o1LPDgsFj7M2d6KU/XQrfJ1uKsDChVkEdUJK
39uQYcqSAk5ysi0kL9UvaB4BP35LVANaYKjQ/ohi4CUIAXv6W4L0wv8Lig3wXg6Q
bSSWdofoAzI56tIZh/nZ9ns42PkeF0VeIX5vuhBVG0IR8tuaCH0brd70hAldq+o5
2H+et2ktUtDQ7Apul7wyHb+NicgN71riS876iiYu/gJGrNrQ3eajlY6BlgHFhQ9x
2iDslruGRksT+1gpdwy/MDAkdTFOPebf9l3k1GqO9Gp4VpdLR2IJL6+9wqlA9LVr
iqfBPc7Iag1UQ9k780JEgSCcc6SQqek4u64gj+uQZq2/174xcfUj96Ulo5+THJbF
8mq1oZSUOu+eHtPEYgVn2EHANPVG8x8kSpfrbaVXemCElVPhmZZOCGWcKdfW3NjQ
aMxftri1P4eNnRYTX/wNg3B1x043iGEeuE9U8PGsFl8q9vxEHO8Pv5QgmgBo2mnb
Hql512pDcv+pLp2acy2CPPBJ4JDlGVb1hgLMI2RgeE8/e5ZPQcR4n2o9zdjiuOux
Z4R0o7Eyo1Hsb4qd8UBgAkxgHicw/FyFsHRlOKD0Mmk0rtYbV0NtjNfz1ejmH8GV
sAUbYa45yFYCPTtozwcNQ/SLwar9nFFxYYOCueSbiNbMQGD7k6Ms9mEVs3YNSpso
CKPaxjmpfgOJnzp3tF7L7OFoLg0xMvOXY9uJeTH6r/cMctQAtvsf7wrKMQf/aPGJ
iDj0GJ1Yb5/BOo6vFzvCNRZyZ2x9+tp9DqTESrZHnAvgCVJaIpzGedlGfjq4Xxxx
dNRZHab4B6RG9vnmqYdng/rBrwFFhvA0kFowiXSGfuALkZp/cgtLhZcHEJQYg44+
OhoBW5QJB1knDQtvUlEHpAL990MR9ezFTcq/mKthAuxzBXIt8EnDAwCrpqvctkD7
riuOYD4fOnX1vQkGJy4TO45cg7jk9N9MT8tNRpt9QPLVyjILBqLCpw3PmI77qh02
hU8t7kwaa+Uh6MjWHffJOzUvbB3YnkhcNKTLDiwKXQOkV8t5B6YMxvLFPLO8+muY
WLCUxMwoOCMwKmWR0VWLCtKaZYM82gwyXRCWqeWx9AuDOc8/U+H/WaBr/7U56U1S
ukbtLtkCk4PUB+eK4vAZhc9YopbCZCG3k2RdRsGrIybGarU96jJUBqmzvgVxYnb1
xrvoxWs2GZ2EMfKruVzDtem/vKbtjMgzPkn+cnFJt7r4QreXBzNlRTHPmWVgqyud
Vo5HH/zsECmnpOiqDPs6K0zs7D/JiwyT+Aq66a5/p7jG2+9iZRUC2lEBiGy8nLIU
W4Jz2mnFLO6JCOYt15d/zmriT8POV00o+T5+GgazZ+Q2TFN210q2NbWi5cgYvG29
Snig6zWboJvpR0zufmJ4LlWCq4kNpDJip71QlT2XuSf7R68qHClvHy2CmgA3XfLF
mkMlALOjGTJ/5FGmapo/P75lt9dtbmx5Ethzvs4eG9/tVRJoTiM4bNOH0pRZ4o44
74uMRDMGNyI8cAihUbsFDvegExA0Sk1+U6wl7K7lLXcecOZEngxKdJsZyn5mSKyq
KK88sucpXPyCXCL7cXol5ehRTT/F3CmKp5hZw7kUdA+3CsM0wSojD8C/YH33/Ccl
5MlBs7QPosThdycQNmOj+k7RSR+KB6QuEQDLZ8plnzihAf4q98QKKX/+r5twp3qg
WREGno+I32qVlKdo9nAYQtLLZAzZGedfcrIQJw9QdMjgXsaXEvYCTxG7LbQaLnUT
++zpvsgrzFr4UBUBvunvBziw3lDb4/plAuBGDM8KhJN2YD6EqBFrZXxT39+eNpns
UeL9gnGPQhZoerm9cUxYUktbsw95i/1NmUZhoubukeSPftsVFxv8Md0MizXFwTK7
JpiA7JxASh5Xwfrzq9FDRLdaxGE7LYrgnLQgQfibCZcjWPzsqGjtAv8VNtuH8HRs
DxFjQDEbhniCp3Mill94uSM3j3Pf648JDyfVkXiVKQsRxc52I0Kjwohm/mhOpofh
zmKy1kUNOXvbhYjfHyRe19Dy7JO3nxn30f8J91X7itzYRwJv3x54KyM5QwRYWPRO
IKcPHuOE86ahwns4KnIZaDpvni/u/WqoQtxz4eDjUW0Qo6ZdfnFcIaogYU8h0KRx
YnMwAgO1FzgAVZcv8Z5T5lHTaFKkfDAZZ+IAR0CrBC0bf8JX7I0I5qOqFjAMq+xf
rM1LCDDHryPvjCQUtvfTucQYnfaRmHl7qUdyQVKddjn7jmd92EAvexwFaXB7B9vU
Mj5u8v0rwxwbdQuGvyDL+5OuU7KlsRMdqbNCqqW52mFmhHp5PRXtTPUCKbcAZjhI
CBskeooE5kU0/gy5r/ndx97VeUSpXmr7rWngKZpxkURj/3edZduvdl/BBz6UkAWz
73W9mfpCmyO94BWjyFuL97BquTwKZvSSiMyUsd4avRac/d/aM0/fyin37o98cll7
E1MkHeyXnQp7gtQeCFhSfFDRf/YZe/BVt+FeIbHaVC3mSz6d7v0dL3MUlv8dYKSN
sgmaiK31V/8BZtTRGPvgmNrAspirfJePs3zI8/GevID1K55uiEDKrzVjolOL1wfA
+2PkJ/ug49fSaA1ZxU29J19QNu3CQuek6p5jGFAEqKVQ+luv67auhqxOADMaa6sf
TNpaQ5iwoB/sIhEC6QaWpTXQcEznQWUU7UIPmUV+uBjyYY77keS/Gryg1Akf9TVS
tHGAZEKHmlaKAeHpXEAC/+OoP9XG3xcPCfJCkqo4yy8gMpObB0iyUfv/BKdGhhfc
YMq10C7gLKvFw5EjnVJvLs72ejqv902DBYCybCkxwY1zwJ2lafPRxzOnDgkrErtV
2fM9J3SOAUVweWpmrASbUDy+j5LGDjiZ23lYClq+DD5I/Ddq49Q2jR3p3ds4MvV7
qaU0raJIm+xi/vO9vesN8Pyjn6VqGdcwa1Se8eevIiKqMWcyaAH1c2y5sGPRBNna
I42sZKgxhwXc46G3ov/RhmobWkaphrZHc1afL07oSL1pPYbCVKRyY27ivRkL6ugC
W/oxCdxvu79A/IR3suHegd56oHqhOUj/P/HrzBy7ihNXNzp4qXaCIesvAKHMotCh
zPeTpxQJYaLSPS/HU8+gOMAyPxcDomJ7cODQ0SKo2CDH+EFWJ6eQrJqGyDngGRjL
ySwQShyk6UWpZMAw0eNXcx6+3A+gccb1RKdsKoRtA4RWGuvR4rc8TsfZBhJGx5Y4
JRfkUcSQ/EKZDUZ8Nh8mHSZinwPaJ/qvkWmTbVGVbvGy5oX9U0QK4iYpAycs0g2X
bTzuKP0xZkhbNvyrQ3mGH1J30CqO7iMufXy28B5TQzQFAYyDa14c1mJr8lJi/5Ex
NhDtTMvMLYLbGWq+bVoc3NtrbYUhffuMwXXImSd5ZKJTYcbbX6Yh74x40lOS/GLi
ZKIBa/Ecbne9W5CiZFaVyWHGX1VMfEmn/FzwoKVOD4YJk+jalwoDDJMVpEYl07hd
U/NB+2y7lkCwIEE6qe/kkQOfumr8gQtW1GC9b9TKxZlzuS5+NI77LmguTHNYOCBc
uGjyIzZ44BRT6/aGDJDILc3+xMYw7HVjUj/frOLxlog7k9eZJItrcL70msMTK3bF
ngDbfyx7Qg3vb+SxL1QuFmXxYSTU+Dt67BhLKcBTA3aGjZIvpBWEfyRgBxBQxPoR
985FrNpgfUOlnm2YVH6q/fUVhEfpKGePoYkgOCqCKLt10loO4dEs/z/jk1sfXbjP
xACnTHzVnIZ+lQKXXENqIXeolpBDCO+mzD4vmsiylDyiNgCWWoDPEbbJzCKls16j
4bCqbzWvcTzQa6uolQBjJafF2YZV1Iur/2JvJHTcf3f82uWLS5cPBwSUPq6x9wfG
OnO/oWGFVaN4A5CJvJV3fQQCxAaokOCxsiKBXL7OeIz+6QHRYgImTkF5z0p/mme9
xJMqUL6Uz0p3dJSF320xVaMeUAX50Zu9tozCiXNOd8/ZEz7pF5oC0XYQWHko7RwH
wlCDV7ArYbJAOSFzVt903GeyGa8qBbhDoiaZAb2Bz9Sy8JYg3p8DW1GFaiI0x62I
H2KuZ5v9Z8T3qCmyayPNJWCU+yvG4nw8w1xawJ7/b6Xu+P97jNeS4XorNSlhwMBK
IkOnq1sfe1crf0xtsZniwV0V/hZYOY4wBS7wF1nQMMp0Wji7lwRVwhf+GlfpKbNt
zmMzphNhIwjKMgt83L8wEWPCWgCpO6sSXAQiC6QAMWpSsHVwSSvA+fUTM/6JFzuV
BTEpLnxt7SgnRs2xUAkuSuKogvUWEzrdJltheY1oofED3pD00wYWRPP75/KLTVK/
3D/dblcWQAlL5AfJtfoQpTtj08bjZDap/oXJkoW4juW5v8FdO/EiGysqJCTTYGHZ
05akPH936M6DuKaX0XoR0udJKij4ry1Mm3mnk0mnM97Hk4U0kE/K1pcJDVX5mPe3
7jc38n3qw3GFQQXgZEnEWogPcp0+ckgtxGl4NMRZzXhuAEF2dveUy1PuNxPkoWTe
Ubl2lQIyjRJ5xMHibXh5PToOVTahWAXhIMh1M6cFfikE8vVTIoGCdSrCeRvok88b
DTAHG5RROu4TrtQnAmEzarjeMECWqbuhsWMb9x6STwrIPIjlN2BCk9trFaxwrdg8
iucnHRQZv83jPL+aScjpcDEVYRm6XOPWNCkSEx6adE1eJvIXFcyfmhwJdn5wAq+q
DyS6VbQsBbvBUEMTzivQ+xs9YiYth2pDW/yeJT4iv0T4pQpgJQoRH1C6ks/xSAdB
U1Aq+vtfl4VPr5vjFHNdv4766Vz5Jap3iE80KFDHmiWZQqgt6R33LDQkbSbm8Rwb
qMJd/GZLPNThVFDC25rkpqied01uhqqwW5OsxnH1QMg6DDHofAwE46B2ghc4mVB1
aNHh3k9aUmxtljlHq5VlXzGUF9f/tXXcqoRkMVOelGFG4rUwft5FGa/yXHhdYTJv
x8kzKm3JHS4ls80NMO2g/CjEkUHLcnB8yYcOcVhGMlrG3nS87nkGlXYLeL83/Tr3
SDsrFqXdUu4M79eLY8G26BjpaXimNa9iSUeFjMLoGIiGQTuXnlk5ZUESlnpHBCU1
XZwXz+0qWk6NkonRtoohxSsRoymKZC4Bn9kDPay4UtxbnktLePLqGza6nhCUvchE
aTFpnqpu7appFWJpxB420w0rE5CXMc8KtCfYk7EcOsZJFAN0MeF3aqxIDQfj/tDl
tCEdmHazGFkxmGmy3pJoq8X48+XNuRRhvFC/02XuuhtoTDdeosmywuXtfTilNRLa
kpPvtyBcx1DZfCVO6NP/Wuta4kext7yAdRC6pxlnR6K9iCSPRQWCBKQaIEWEqbRz
RUN20c5omxwvks8EEYCSm1okeyjOrQ1yxEET50LI+qPne/+7f3V2/n1OsLMucdY6
JvJrD+7nl2weV+Eg0C09d5DK3icddrgRPLiXOsv7nybGiOd9VGHYAsZeu0+4bBQH
bj61B0xmb/9/shF3159jLk70R3xNB6gcwJg88yEA9QFIXqfKmsAsCGVo32mbehkI
I6ckY34r7XtLKCV+jCvTlkv7IIzvuNaOwxX4UcF/84oc40ZHGn2Z4E0O97qIJOvl
/rRjHT7Hhd+cFBgJqfZO4TPByjgLufmyzPJirX3QJOLwZ5RRucSHRkz9X0vjUxLd
pCch+pHiMsuhsxkomi//82Exqp2LOfV1KMApFjmknGD6JsVY8SuGSLbgK5zdY3ee
cKjoI5Y+uufO5VfwQUwE5QOAoB3s/aw5L9dTHmHK61ccJU3chwpqv3Yq+Y8joa51
Ar5r1xxQk73zz7sIOIItY4HKGrs/WFg/NjWyT0XsEIyMYIdARCZ5495zMrmlfn2s
JQhghr3hFiWiRv0iZlvDDq7QuwR+a0bu5Pw0mRUrk9b20LTAyQmJRm0ezBLXYWvD
A33ia2e8skWJjbqRLkgBP/MkvtxudWlwCYQqPwcWlfFqol4ZZmUjg90fUMCmzKrR
vaX/hwsqu7ySqHOhJ6R9uV4mMt4V9YsqZn09xPqnx1zn7u0FoToPR8AkKYVNYhqo
PrpCB8U9h2ryFtW9VTqnKPsQjAxbO3enT7mrVY3hMnPQaIvfK5Bg+bKat/iIj65Q
PuQZ2Prs39LNb9VhDET7fZeA6tXdlNnMqVl8ku4dm7Ig+ErKCOyCaUGkj5/zrd9N
jy9WB9B4AUwdn0OyfZegGae2ry370rg0ZrYAOC6+Zj4B+W1J5Z5V9nPHGZ6bixvY
vuVwqWWOvMqHVvb6fan6gOH0LTlDMx5AuMMZ3slbJCszKYqkWhTZs9CE9qmKmpB0
geo5+iD2we3VxNN5+m912OAdqDiWf6yyyCvHFiKJRHjKHV2gLjNjiqJyCCU8hrzP
Tc47nes4FIgNn2z3yMYpaHM5W4uR9NlAwSCkIpw3NuAiPahWr8oe8vL8Yh7YCNhQ
nYz8HEVq2CDXXuJLmNGnz+Mja2iA9CudPvMcKjzrUyOeGbhAKprNfrrCHiEsA973
T1oeCNDhAkSR4BldPebq254BI9dTaHB7voSdEBWjBypU1XTTdRyIEv3HuM3g8pQJ
WXuEc1rEoBXjSjSzSvQ0Gprh1ncc0tqOEnVl3TEtAp7Ku7E/rTWxfzUevYbg4KfN
k6cN24tpDWXGHy0ifGkDtBHTg4NmjlqvKPumsTLt2N9WCFmWVFqjt7xXYRkvqbVl
Mcr1dTA44GyxLy+CkRacRyFEPLhdqLE8tpmDM624yLaAgzG21MmSNRtW0nYLZcco
GUpi3iWZjGVLVmW5+ypVqTYdO8bw75vthmqU7hqawmYsuwX6V64wDnhDlW5iIVy6
lxFuI4PwSLv5rxSnqA4WRFq8yWmoKSvFnkUOGFghmE1dLCz9DbNXr+ywcVhMmBeG
662XvE0D8+fo7xgCifxkcW6m1/i6vzGqayPlwwghfMZT2ttau/OS017/5GqrFvjH
dYX8DNOGINteuYZnasRKGbT3W7/IRq/DUf9omd5+vg9ncov33gQ+o4LIShG5u/4T
F0AETBo3R4Cc0eWawaOekyfldgODf83RxVEexaPEyqba1ahotPasjoZn6iOD0ZeD
9pSFj8DtmPvJnod5rd3097Rzd9SNXi2jF4AnVXOcTiRMQN4pTHsC4L8KkNUTMJ4E
w9xuOJsPB9jJYzY7IyyZHZsUXnHNJhRaZoQ90TF/8bmcTzpZRglUiWBNY4167mS2
BuQeRegYLZE/dI8Kc1VYvs0z9rIXxJIxAnrYEoOgWZZ7zIer4Wy/qRzsB9uJkdf1
3FPrwk4Q1Zc3sqJ8a5xVlC5bO7EnG2XnJGGVomDI51G88ZbGKOIUCUdncCw68zkl
H4sPD3kxZNnxbAj3Y67TXkWKcqr+cBjcC2hYGvpdwTJwtjHW7/Fjre70UyaJsgvs
VnFerQlMpsGdfOVLNSClm7NafcC68qoPTkEUBSwOvqeytNwnw6ED3F0MPAoRwvVv
bYAZSMbiHPr4pWepua0oTpRdRfqNuUbkyvs13PuByk9PId1RZIZUMXTNw4fnsHxq
uU8h7qxGDbsUas5NI3+Qk05jzwHuqUt46yOSOsCln406vn2nPNU6ei3pYgch3Amr
MJNNLcn0HV61sIRxEdfatvtAvRghKXGj1ntHEeLU47nYSHoXEAySI1F571tm7Wj7
h/XiLUVjvHX1NzjEab8dKDvBI0io9O2GR9mqjsNE2mK8l2iI74Vkmt84I9SCO7KV
euFN0fdjbcAKRYh24Rnsgdb6pjJvnEOJewLzh2rQzT3tn6WYt0BHfilJzLUP1FYW
7smwc1sW55ftBroIlS/Zc9uRuOGFsHQG+gwwaml4W0a0M3o73cLu4V3HtFGFxMEa
rD2Gh2HepRohIoPRWV7B8bmJtQSeuJ2HM2pU5cf0ujEPltEfVUmI3fzvi2lU4FVB
fxIwCh9rvL/wV7Bdfc+rcow6lnIYcVegbxLRCZVqpqzbrTv584PjC6Q3MIBVM2KH
r1uE/LvBOBN20F4Rc4uymYX5gBkohZpF9pxdFcbu0l5vaY45QwwWivC1/RoD98dl
aUSDqCS3Sflnn1w1V10wGKUJ19jxfbtr3W05OZpU5ZHo7UeX51uHnarVDbPGXPsp
xPzGcejTGkUBJD/ZSZgjed0IERF5fxImwjgKFrY+b1h2KhaYxp6DJ5uCb4zJ9i0N
+zscP6nk/QGWW2uzkgqlf0e8p8PpVJsnHbp5wInih51safwKlZwGEggYhGYa14R3
oUv8fZSc+hqHx4thy6uxf2+811mM3+krUH3BuHKxAcVz1kwxtqfelOpxVmbVghHq
0RePqKgqxQs9UZZH2UEB81H+DtrIoGyL+HaYj5b81fBCBoqcy++tGKm+mKKHdZll
YMPGwAcLkS4KR0ITri3PCRxQQeWMWq9gSMC+DRkph8OKdrG2pvhedCv+uTTIxoWI
ROX4Oj78CZrNhtdAMCPJDdA1zjazW4wQrZJpNT12fba3tZMpXFBDV++3d+zzWye1
y4AX4bJtJp99bYsAK8KNbWrGK/4I+kvhtsu8U9NMNu7T+5PbHtWB04UPsTQQJSpB
bIY0z35asIET2hWcQ02/eptXaA1TsekizI2AWqIyhnAFn82j4rxHvfbL9UrcpTuw
RrPcjAaGYitPyTsb/SqciDZk5l7SJAtSxdVZ8IgitRfYNvkWHNYX863vKAGUbHf7
LysdrSuXh+DJkmP8VoL1ISAsSLUl15ri7YiI/1DIpsYyDUrTqLTK3ReY/XQcA8ER
kVHRpn63PLgWqGgFfY+OYjbIXN1WDwxPD2GT4sh+ORAPr/A8WIQhk7Z3wj0GvL4+
FnUEXL4AnTTHacDYSFa3G5RjHIXfXD3nkprgxFJL/xkeG+zxEvrXvbKrmJXRVPmE
vTQnSAQI+lBX1TF1zsEnKbppJ6+q3hOrwMV8Ef2DmUUDJ+gwwcVg6UKkAACJwdmg
K4d4lV/hpKvuDs/Xa3qmhnoq57CU42Can/r9uRNsmWBaFINE1Lm6GTn5chp8t2JO
igCziCPPTqsf7073HLWbJThlD+WkjRZWwl7HywmggSVXz4NPZmKZ5GNJj2KaF/E8
hCTMlBwxi1r2Z1NUZqWTmJsmfTm8apcK66mDOlkbOGFpQlqehB1N93MfrweUGRce
hMLjdaLblzE/5x16JfW42wEwemyRB/97xdQfSuAag5+QxDs+MsC/DnHqIGhyyzSX
/aYW8cFLpIfDarOuxbtsYa29tHAZC7zWIDOyba2v7DfmCgmuKKFiVT4ZwNwKvkU2
83eKOEDMrrPBPEVMPoiGiPpm29KJ7/yza1O3Vs+Uo8XB4ailS3VV5nd2IJ/X1y06
+CFQqy2TXTqqf/BtJWj1/NZ2bs3doONCLqfG++k7Z3R2ILxhJCHGGMjGsEszIIwp
VQHDWNKxlip+rDKDiCh/V/6rI/1ZqHs1Lrnv5djW9i9/bYpNwd6SGAHVJ0mZ9ujz
eKOFAOnUbOgDX0i5f7WazzL3epd9A5yaYnd82gpwfoM4JOub6tkEZQsH+dMqF/J6
orS6CrIM34cP/+c/h+hudX4tk4TCokyZ3MngT8gplW/llg1yM9dGR5NKPnwISp3l
ksToj5e+mKjUMZWPwPRqblZSDZB/Ji9d/wvfBTmF0S8FimC9XAF5XP+Uq8Y8M5+5
/gxT5LhoZKxRi5kP1H272xmxp4Fgq97G1mbwI9sS8tR5xmWI8m5KciKfvj0K978T
R+mngfJtkxJzdjuNlQeM+YnNBUxoR/1LM+egWABwh9uEtW2OiMKVoocCC36n+BYn
a8/vzG0vwI+WIgCXbfodSM/E3ze3VkGjn5N3XcMu6eY+E0pFonTNTCc4gWCK+zho
j44+WH0X8Mo06m3oIyJokT5oAW9FaPeVWfgk2i5GxgFtsdL1znuHUcEdaXNfj2uw
BFA4O8FD/ktBqZcmMP388nAIWDURFME/NddXMlHtNvoCIXwTqavvA4wrvPwhiJcT
pPQhkLnZ6duMpq1a0Q1GYFdaDk/0tDrZhlEl+KD98GdksDcQxe7dltFRTyuYHmTR
4Qv43mdbOImwoxEUeVfllEz8VdoOENMaqw+n13DvqEWI8Xqq2doQp7K9EqqmpeKs
HIpoLub/vMvCO5eN02CbwyWBBiJf96qGkOX3VEpQ7O4dIfvF3bJenCbdpHy24M4F
RXqEwdzyKLW/Ahs2qDAjnjF7/1rZK+sFd1J0cFet4Osn6XAxV8ZvmJqJUrg3csUf
T1AXu3e3hcn4Bk+sRI7QafF3Y0FH7VAEt/ARbLAjB79oK32ssausF3En3Q/s4AVw
syOVuWiShRsv1hHWjTtb+t2o1TSkobRk92rfyzEkSR1FY0ycmjw8zBlxqaXdMXMN
nCkO9SaVuCi+0MRRsufY5622AFjvS5Pz7eW/ZEfXjNlGRSafAqqbVYSvepZ0xJ0g
TVUYrqMp0qBgbbBVqu0+o9QZzKDf9yRSVleufVDf7Gbd/2brrKqT93V1iEvcXZCt
lYHwkqjlrD0ijjYMqmtCz4aOR3QovdyR5r/Tp4hIlIse2KPi3KpieJo9m4gY0zxl
cHCyk6Urkgt084MZWR1eBNltBLpH2KAHgy9UfHdFTSTdXT2M5I5bwbI6P18RJNMI
U/yzDNaD2+itPkXw4EUR28Uof115P9cdsVWOdLqtEgY9CMzgLp0lieguX6yTDJOz
p6QbhvKppsmESZQLatoFZy6OqocuMGKsGixPfQ25FYhEZqW+wNI+y/optga00FYD
oscVdVbtGy44TljGij0XV6EHYmezIUiPP26H1w+BZ83L+qq48wdjiIXtsBMjxA4O
5lFbbDXptI1I31g6eo3NsKT9X15Mn+onWOrVfHHKYhpKTYFWK6WLy65FpVW4UDIT
sSl4xnfyhBYo6+lDkuwzyI60fsh42PBIgvrh1QYOSUNzgPLB2qkdCnWnyNcvb1Jb
sK0jkG+OfYoDKcunAftaYbtpqfEmn/b8UNrcHN9CC20qp3K31hcycO+udxRxYQE/
mxKmDaXv8V4AdPZRX/9LaH/ixr6Y9wwLgFzGhRnlyzd8a/I1iqMkDQB24HuUqTid
giOFsBmEQbdPuxSmVe4WInDWXoX5BxoO10/Ebmt/HKBsRYG2ABQ7Yn37lw8BoVS4
3RFPVEXl8Q71R7gGm782KutV9E4zPGrmFDZj1XZjJnSDaBBVVilp5L24MpdR8OWV
4X7d23bSJoyr9TtMtRVjqTifu7CxSWOYvo22EMUCJEleHebRqKQakC2CMQlLxnPO
Jbext0TG1trpAh4pkAjnlK9xNeiNQGJikHcwBNve/UPFX27CKa1B6p7B4ZaEaiNg
rsi769J4m3kIMpVszIj3zzlFbsYQXuRZOxuWYnE2Vlh5fNChb3wagc2A3UveOtCZ
I+sDR9603DDB1UM0pd2Fl1DdqPcmX+bsiVrOMyHPll13wsGLRuCgbFjNOZDUuztY
wwuxoFaM1BUmr/etKkO3fx8to3I2cVCRtOPePXjYoGAmpbwIENiY5lGOIDYb82qY
QapkvlL6lqtzUp7KwDyEZv+fKE0ZB2uzuKMORoOM2G2yTaTr8oS07HdODyWiCfFr
bhVd+PXWantw8KwgzZLbDUP3MGZmWFzxzjL7FuP55jzNlUZ5eAVZ896njtqi/Luj
R88Lak3+FbDklDQl5ucLJOhGl83vsGhVJgmglfzg8i/sfeVQeeV1sh5qP/xnk6s1
8c+Uu1tPHrapKls4xsbOkkAkBz7EFAW8A7hN94/KaKA7fsLN4rnMn+EzOh/UaSx6
m+aZhOqWT/K7OqLjef/YT9WIHtTO2bBydvALO1BmKgTKE6e9keOHuDTnKskvOckZ
ll4u72v296UGDUUVn0I3WDjp8fOXoPR0m1Hin7QOs1mU4NBoyGNcYpQexIW7RGVX
ZuIqQj2senZCdqPS8q/+oC1RqG/igwSvuewfXuZlf2Y/Ixs/jcgvxz0FxXF4ZVcK
iiRMvVMtt2156XUIaWNBSEvtFXf33ylmxcEn8JXOUYu6/cjckGFw71Uxdog3U6By
b6y61O4KGtHOXbdeDPsuI0ZUpLnYXy1efrVBmJhANSdOHzySJwWvBQMouuEkFPeE
dZh3u499QRCbEeRebEfeSZpbx0C/xhLLiM6ke6lW0sLsQ1XvG+QjluNvOsUNXb6v
IFvXZl2iFiXPij0UAXZI67Min01Wfee4Zo09MNRoCmtlJY3H60zSND4gNAPpWzTZ
3mnOdYizOEitsOzcjUMVAvEr0J84NGR+xx1T0ZtZXpThZGY6zBSIw4ZekmVxIi8P
+wSAQExWs/S3TPjtP8GZaKjFRR3S/3UkVeMjoXF6kGE03FcShOAg6FIMPbIE+Wx0
oRcIP8jcAJ+Kfjg+jFaKrhsJJGXM8pDL5PdIgM1EVtsABMNq0sDbHVxntlVeo7aw
lwfzMI/b4gWu+6R0dibiFl5EB6C5e+pkQtTgNMVbsm08QBefefHTOKvyt9dxGcXc
lYjO/k7OZDMy09vROfvIgSbA/EvNmL0FaMcyaKtETgs0oBFHCrrzQhh2WM6WfYgz
RfhB88LWSXNRHEHJR2bPRONYdIg09lzFxPig8SP3MYrM0GUo7T05pVa+deduOIrs
dVEMq4tRr1ChDZlWqmOlMXodBJf9uSKTARIWw0PvU0jfXYnyx8r8fT1vpuw59wDl
wjROUPrmD4DlPqlxR8kG8PulxwxX/IPisaPlnJUO9btZexP80eHHmCXKIAMwejZ2
PxqEvBxpxjwipijWrwp2RkadlNfWe/goqYwS2wvdIpgi31WHLfs1ZxA3tBGqqKka
fGudQOe5x4NfnaKPdwagzLbgAjwqmlMRjziVJJCrSyPoylbPqOJWLbbkfpKzKQjM
GmhLjZdOCeeqdHZZFlxB9ciBvhkMJWcKo7XGT1SulJGYUZ/vJvZ7zN4f/BntijXB
OgNbayHXB994MXFx7IXv+MGeSl1VhjmLFG1vs3uB0qS9/NOovW0Ra615jfP6QTYb
fXawdH602FJ8BZOnsmpUCKmO0CDAg++S0slITy1js9m348TIB9qb9yzjburRe73M
fmSq8UxT0kH1t7A2SwpCoEhHTtbSAmwX5kQdAe+S6DsN/kavkt+rN9tQ0+lCX38e
MCLmFmiMxRJB4gqcMo8dyswPGuZDDPe8yIF++UFW6uO2dnzrjfQpRky4dKgV1yXN
qxElEHKWXOLqj5S/8o0OTv+aOxy4hj1/LVVWiCIkMNJGZhOH6abPCXpZyS2pc6DX
3jSg15gW5Io83McMUCWMkcPUcTNwle4YLdQGM3GoIp139shYGZHRCfoiB3ANOOqd
SNzKcK3W2ixuK6amwwcUVtD0CfPJoxau6WMT13qnmjO60bju0QRm3dtGp7uvsqv+
DhLz3gW4hus/CQqibx/sxfKD1GdE+wD8ZwCKz093WWXH6A1tRcWHz/e9B2rcT2nc
EnT1f0EtGWqnI0lzqzwym5Z1XjGkbEChkRxTOLiNk140wQOgIP9z4IMdcHYPwPge
m5KNp/eZrKFpPwMOtO/eO5nYH2cYcFu5uhE6o3GP1VhPNpPWrFwAr+ZpwPqj810z
A9KLXdjNZrddRrMjCYAnEoFkbkZ5bKRR7+4xNR9aNgfOeFYFXmWWcCewcIyaM5jy
LO3NnIHppX4Skvi1Z57o1K+mD8eFMNilV/KEI955GS0rs53IRSxPLBQF+Y5n2QET
B5vDqmSrcew6H/8UX0/IiAOXgwo8DlOlFWY7jbvoJdXQswD64PTmJ37Vk2z9FzNo
HTlpegiPgcLR9CfTBUltzFSMKXNc/KzUqmTtuGiCWahLrJILooysCQAWtczks3Vy
3KzPAJ4ZqSEBFObHtvA0+PuyiUADXpjX/5npndsaJhXbl4wQYfIu93WmpQ8boumn
sx07i/qVI0qv0D+iXjRNHnBUyw6VSoH6yapB5qLIWy2xMLtDi4myItj7yS/ygX2r
W9xjIpNjxQ4c49qHHdsUAwK+x3vWTUBbcjYHejMa4hZXaFpKz4MHRzOrmwYzkVMk
LVDxF/DTjGUOuIpZBOSUyRZgJPfJit9M+Mqr1C4J6fd0o/cRbl+1IKqMhOP2ADhW
MVv/ZtqvrZNVBRWqiaAcFcyTh9rM7f2LFTVs407QX/QkdNCPSnzKTmTxV8MnYQkv
wLQeY/KnKZYK/ryCdNVWIrCHS587UJLh9DOcYJ+XhOg822j0/hjWzY9MF4/qhIq3
Zx/oMBYjDyWvwqOJTOuwzlOhI44cwGu8JV4gPeM7ZMN4utAFmby6aG0qQlwC/R7C
EPODOlZXFHwP39HEVYMBxewOpvAL0Ki3IAzYVAAKhY3/9BLoDnOCXINs5sLY/Cr5
tz/eAb70rTby79bT3dG2Yo0JFaMeSvJtGwv7lXpp997rL3iknrjMei5EVSNO9lWl
ThmympcfPr3JdGZzB/1pQQDMxq1LQqcHggmD8hpRdOrx4+Mbupf7j0LspIlueZHj
P+WiX5ph+yOGoVexn5ySAMslbHiAu2oO3lalft11VtOIz9ks++mo49CIUHd8LbkQ
tAHkxTOSiFNPOjhNKLZrqAi5vdClB6ox2waQdpOCHmvb1rU9oGhgvgPhzAnBPDNH
7psX1b7/UOGqZTCKNu9P8GyCESdeEg+95io82BB6GQThN9duh/WNPgQM0LeW1wxF
4DQWdlVwvjsyGLeLE66rSaGsHYGylpzOKcHwD4Y7O4KN+qKITp34KSoLI+7PPWZN
bVoyq4M4596unFFcDZUideLQ+BoNi92VVEP8L6qWIdUCA4W6KhX/Q/fRY3KrDQTW
GFL53X6+u9KDkYT4hw8+Tcd/dPYbLskOpABlUJQsxhXsA9wnGD08CkniPEgk0mMz
rqqQ2PwXuhQskfQC2pHljL8w9/QiFL8ZA/09R0IjrQ6bZx7kKYDEwqIAsG5V2qfw
3hPP46PuunGP0bGJgfx1lNpK3BlhQ5l4SUzlbFz64WpShxrgseWG0pwEv2KIRO18
Cg4G4XSNkthzDGYvcidB4jb+yjdbHug7aw/NOn/E5+Ra9NA3TidJjHgz7kYGNgxl
5d8Z3um1TfM1ADWfZwji05rl7vqKTKhxfKCwPauyEhD43pOFucRHt3NfNoZEruFI
CqeYVaUAl82bcU0hNeTRhyqGLpSSqxnaoFQce2vah9UvbhRALgEqcsHqN2VPbsfP
aIy4YOJg3Qu06b37d4cdx0/nhE4fCR6p0mn2pK+r+eE70G2VUVNf0c4bXxoW7vkg
m0U/lCReuzdscFaNM2O2I1gNrRjarLFYJBhleBvGFUinBqiHdeDDP9d/gQv4ue6W
Jskp2tW/u7LUiTQlAgFpjKHJqE6r5zAtXNI8CSEqx7F12jFDkfGz3eR695Y/oIpa
hfGhgyLbvIbvesmFdWuRaBpHpnkLDOWDpK7T9MAY23PV9QtK/t3O2jihrpvRiUnR
cSlm837Bq2k+Y0F2YNVd0nn0Hum6004ETCMLC2SdNKe8488q5TGqYmzFa+/3Gjdh
q34TSAq/ziv5g391oOcVZGN5aQ/Eu5T8GQ4SlAUeb3I0bVpZy+xy45u5FJNd1h7D
yovkhGAxMGL2JbvBZsjPJjIEFjRt+DJYO/0f3tvVQdgsuJcpw8CEn4IGBYi4iJs8
Rb3xhQ2wypDgyKj6m7e7GZ40TdZddWHxxhvJ3FWZQ3MSXJN/kBweFH67l2eGw34L
plmFUWO+dKjx0JqivGHZW1WfqQjEfnblm5ZLzBD/mAv3pJNkESMCn+WbuDsSkzRA
6KE+haVti5ymn/LoGaIBHefAYjHrrar9kPlq/bPH11knfk7GUR6dPuiqy9ci5XnC
6sEzXqZznk4Y+VtfxuVXDTjzraGxy9Dnh4VVFhtUV9c9xLhttCRdgeKpp6f7Hhrn
k5GtU7vsphUUug82o6B432r7jFb0Ug+6AFKKwMm+m27iWRBxqFwh5Weg3A4Qo2NY
Ifd2PwDl4tnExpbFF8q1iaeTbaQXF/MYO1KUcRnnWa2NPB7kOfko0C4lha69Qqwp
/hOZbvlnV56y1oQTHX/7dk9Nc7TqceltC/99SW2r0wE4LzQygMAtUR2GsDFssamK
MgPKP7VhyCbH80lo+c0iOKznCbZEHbBO771J46urHjktxAuVJM+4elpfmU3SK6JK
zc6gPOYW9Cu9O7FlDktIGhMbPJ6ibAZymPRVez+F5XcZhqsRm0Y/H9KzMkjz2pka
D3NkXEpLgWYWlNzpd8Ei3fFW2UnJBObOlJXTTzltfH0xXiymLyO1H8dAAZNChufh
8xpd7bLUWEGxJvihlfH3yeKE1y7RYktdUL/o6UoZ3c9+tN6O6SbdJDYA4lgvjb6b
R1nzMmEigKvhr256s2q88DvL4uszOBo4TM6iU9xGIBvHEnSyeGM/+Ruc6ZNggvwB
onpjHfqlk+PDG+81uuEU5FLqAMaQLW6PQ16QJ4YLzlG5wdHLRMcW/iDA6baXrOj1
KZdUN0i2o6dU3l0UQjabCcBQ3VhEaHyucLDCTriC+eTdDlLg6zri90/QBoLWBFt2
dcUteDuUDyvI2W981P99t2vpM6mhbjbeH5KeUpjisBx4T1vKR+UIhl1oZ9pMUbc0
yhvzXy6JktYTJBbzFi6rhS1KtgXoRHB6/nsxtVRUmrdt1cfU5INXbmh0TrS2N2wD
WGnolKPCMqsTPEyfbkNVMWFal8mB3vvYw3glR0pb84HsYxkYoyEvzKUovtJbNjFn
eEdrwqtNIN+h/zwKTm+q4gS1SvWjavNo24/IgqFbLQGlh40DxteOkHSE0OjWLC0l
FkXcZMgtg6wVndR/DHw6nP50E6o62zk2B2KrXwal9IZmI6PIIvzpPD9eOvv7TFDB
HVvpqDu7ZJZfaC1O20WQr6aF7TlNpoydH0mO7Zx5b+DV8LoonGac7fEZk0U3Hbnm
iVN1YsvPFMn76YdE/FWJ3aUHtj1fa+6lz1fcHqxyqmqTCeB0FGH0hlH15sfRe78O
wC0pm1McveZuxb9Rpk/6qziItnnxEpF4bGXX56UbNGivuZ7BVrIDTjJoLN9Rid4l
ZIrMNd6YmVpKqD7UIB/tnm6/ugHhV23h9OaOz511cEHAzoFedtk051w6iI7eIXFC
ZpvyqC3pBdHaWYI3WTMMLI7NL41z/FikkTkGQj/bUoDlmKtirF4nCG4TevArzhfK
cMNTKCd84GIzRGDwByJ4jmGkjr2YzHoznA95ZKAN+7H5eU9G1nIzmHT2LXaj9chm
Nu3t0RazthI2Eor7udm7KJoU1U9xZf3UllaGMe+ZuhkuDRWjSYyzp1EqssnFmMAX
+lPyzH+LA2ROASQmKbxnzkH3N95Om6bYOgzRU9naSW9SxgWmkOksYMHASvrSOjds
HPvdBvdcla/ntKSwfrIs9xeThVtucTtnYy0XhJTlLDhuFkox8eUYWBHjWq20WejK
ud8PVTvY7icnK+skNELyNOJkAjkJYm/Z5DT4R3btpXScUD/4mJ1bkN6ZyTyXIOf7
cddETH8CnG2LI92t6bKNeJhQSD43s63oQwqdIx3Z6pi8wLPrnSMqHJHScaw05kp+
ll1Dv2uBwu2g+xe3YzSfbC8kJl3d4w/D7N4eGF2UF+Y3MGZov50Y9wWeNggCRX2b
DsCh/cG8ikPQCWK8xHZNcttRZVFzwby1Qza9iB5C3LZTU2yBe4F1YeJDV7qyD7P7
WoJtGriDGRh6GVk9R7w5tiG+4jBQm06JiKpnfTPptovM83r1jtE72HzSfbX/6erS
geTKfJWoruXMljT/IgirJikcUP+TW/rGyhCscLWnHkiWedGbdQ3OouxcYhiJyHIu
U8YkR9l8Z3m3ZP2y2yZdf1Hujbn/YisaT2o8UYdRkD8TQHOCc2vPlhJg98N6NMAJ
GV0u010Vv7D0PUnv97E2vIXtMTANcAwQwPzqZPu/6Zz1Nuj++0iLHTG2ob/0+A/9
sfDf4KDXZe9X7urpH8UhwEjL39jFveyoOoO6B7f23RRUG7KmHAnhYkTySA7RSu4h
D+YX57SREE8a2f21cL8cNrfAR6gWQqnylh0EUM5CpGtSQn4ZjcArwwTmrHT0CQaO
5nZGpPy63eujEkH9ckKNEiRaRYopdSWBzrvZvCTWdXFAlxCkLu8+cfKAAaG0rEz8
WKWk+IC2Wu8pCiWAQbdZN1QuKESTIO3YgzDm7WZVdrSjXteT0TYwQKgnX+wPVyFA
1JeAx91rdpncSIa1s/SrDUNvCeCwSozWtX/mx6JiszBu28jEAuLVUnZRSt3Aaw3P
ouW8Ks6aXhj9KoHIAxrWBb91z+qOTV2DQh6fNU3iHrX2QBa1nKMSElr4Z8Ttwaru
2Cw3q3mawkzQ5sfqIhdTOiqiF6HzdfD6IqiOdsXPhZ8ZnKtobEGVBjauQqNiZ3jd
aY/lvXi34agcCRDrTVJ6rG/7WLwnIBrBX5JmvBOqJWqAeevDRPUbZC130kHTwxmx
fsUkgU77Subdcfy6ty9puJ26cVdJwmqAijbJ8GYDnO1W7UAhLYgBMtX9rxRpyh+8
8Fe9D4y3REJtqSn1jtjokezuO1x2mgksr4evBbc1x4Xh5rmC9JARnlQEBhg+0RGd
vsFR7Eo/fVvndmj7saV51N6caR2w5Jvb4tdFpfxu7h0NvR8A0Q2TZ2+8vGr4kF4b
aML9tFqVaFV3awRA4pBO5rR0mri80eSL0yQ2a/HMBVD/GoW5RdtPRuJ1w0FuwfZ6
ssw+q2wdD1dB9AbYoSP9fTkEx3irDJRzkepfImFenpsI6Wn8ietzUnaRqDnxXskX
bkaC9h04FmCphB93LgseqMCPDMimXho3tiFMt257CDhSHBsiviwvQHNHKJZMlLbA
fcyvadtXn0ca871WIcOoJNgSk9RQxu4BpMqaxqvbVqMbSlEgssMr/gHa1Ja+2s6k
JHDp/rQz4psWGCKmWYgvzDoMRzH+45mS7jYXemvhp1vdrZoI46xR7pGLrzB6icve
D79rPQAba/41A49PJNX4A04Nqh92r71xNjvhcPe94SOumkAhh45EuDUQap9ijH4Y
hvSb9iBHo8cS6tlMSFHsj44EeNEwOBYa5Hng8qiFIRgLkQQ6eMB/qy9bKkc93gAJ
b6eq14JwqqSpDcYXVFwKjx2DHbNyW/Gt/asLO71U6TMM4lr9Gczxtue6WjxsJRP0
VH5+Jq93aERFvKm4Fed7EnKTqLQoxshPNBQF8g3GmRoCK/HA+NX1Bw+nR/HMOZmZ
g92hek5DJaKP9JxIx9yJYnJ0E7uowmUYkRAccmz5b6Zd4No/UOT9PcnZSHImI98H
Nc/cdHEA7seDgNcpD71Ipg0hHDp8XMagVC3AkniCkLwQQXdbnrck2h47urYyO24a
qUqKhgfA0YkiOq838Y4T4E+kFWuI3PZ3RSOzN2LAWJpXmzUCXl8wvh6v8KyH7BA7
TWeaY1r0RX3hAjUPLF2O1tfKiTNxs49roqPBog9cjenLY+G7NN1pJl07pY6EUgbV
2leAFjJk1o+mXpGxSmsaVuxA1bpiyypbF2P7PRjBGpR5xaaB4vp4OunxoAXIE2vk
ZdyHV7Fqgjb9QfO1FUXuyQHk250cm0md8N9a3grbG2pXzXE7b+N2mahuiHYPzc+A
wJlRaUzLzCxyAUWGuUmP8GVjNzVtYjCp7Y0u9ymB7sqrhIPnab06v0tgR8dGnmPn
XD13bpTbHft5InyqGcW8TqzATybfc9dHmQunzxwsiWfFFqsbk8LM3ffXvnK9cXV/
Kqf8RreSJqdfcNDhueuvgCJR4TQxswAk+8fs0kc/sI2jHmuP/OopD7dqosmRXUgB
dXx0K9TslmaOa6399oEsYGTuyhXK/aiR9rusy0+9bk/hrU0qhbixP+GcdkxUyJWw
zFC6wQtpSeaj7tgWP+QNKMRoVk93c2QHzmbJxv5Vf8OwKzF2Avt3GUgmId7HUvnc
bTTy9z2IJSgK6ixj+YXWz/o8QZ4YV1fJtey0N2vRA+WoUBoe89Q8fgq/bMhcM4Fv
HtAcJ/Fv7xz7RroUSXijfxKWcn/VDUTozOn8Xr+8xMZQI0Ku9KkynkFw+TCxFZN8
UXpDxbKdg2gv6KU16b3/nv+qq8l3cQsW+jg68TfuEhYO3OFG297SBs4s8zDojrzY
/kt9ZvAXHiqYqbWg++HqaE3qeYCWbvz2K1raB7wp/KBg9ll4VsuIqMuJf69a1d3t
KUjUiNf9SrOT7/JbcMruqgR5GBafx3d+Nk/fIZhSAl46wFpE3uQsXRQHqyavPCyw
2v0pcCLHRdfWQSsoKQFoqUSzsOQ+/biDGPgILoibTVMQBhfpj1GxsuU4p04L3fzb
CoIHvoJeGK/QV2hjcElJ59Ad0onplpcXzrgDPNapx1m6kjMJ1hG2BQB9vfbBTpup
y8Xc94YrbUQGdfmnGfgGonkY4L3aTZGVgiJCboIKkd9Y8cLTatBxV8A7W3zo8HhP
iiL9rJsNXdpdKsrIGLOgSrIl+OV5ll9LRIucoyafPqRWhuf08PZAAIgOp80E7LWj
hKDp+taIxyNjTLGeuTn2pOKwZ7i+omdW7cHeKFDv3ui6t6P5Kno992MJZI9HoqUh
NWBIPhm2a0i08B21Q3REC+0vTG0douYC/4N/W9X97ygqV+nKJGKhbTefz0b9Q5hi
sQVMz6dTQUkDXrnHnb59FhC2l/rtjzhBRL4MPJtHNClncVI+k1r3BCEMQNFo5XuA
CWOtXmGb8TZrI3yNbo9sekMPbsnx0y9Lr6TmBtF5CxqYllNZoNCDNyhpts1c5Km2
5RbJJiM9sB9ZVWfIgPl+bDY2Al6doMjUSesVL9KkkqO0crBMxB3RWhtEz2qKxruw
qilEqCTo7+5cYKTP95a3SPl2TeYRhF/42njrqCa98gNMnEY+82CpejMecDalvBK1
zQvrUx3lezfnzqsLQM4gRO7/56vOXQmtCMXDnBm3lzQJTJEkntn9C2EjFUiXvDCH
4bcPdEYcX7qQfkGTkQveBOFaaIzGmn5l7/vRcEaup7fGRPzCSMOvd2MjkzTBf/ks
j51eEHkzBkjwWLUprK3BRetO8t73PmrZCu908fwDeOMBBwtuKFv+M5jNeT3BFmx9
0wTE5Peh/wjsgnyocybYK45jmGth/kY82dDZuclaXFI3G3jDR52q+uM1GZLwBmTE
DBIcRDE4u+jU4UWbSPcHp+YB4R+G6rU2C30yfkQSCPoz2/HjbIpM2wiRh9kn5o+z
gRvNtmQLg6/fzpfj7rkDODW03U/lIyWwACnO2OgvvZ7Q/IsJf4jvpRAdDa0/L5PU
4DrN+mOYw9PuGg/ofEOQhboz0SkJYI0NC9ZdInTS8OOnyFVOc8CjfhUDy0gDQbNp
J1IMk0D3LRaUsDytzXHe/CuZlIYD6gHaTYOPMWsv0AsnvyRWOGEQ8tl43zK0vWRd
RNXE7Uq5cI7TRFRiCCCw62MA3pBrQAE7ttCfkKkcMIq7y1+CE4cuIH/aJnr2z8Nt
lzyP7qC4Ps+ufcNX3x3OY5oQK2cUuhBHU0/xZGzzW3mkoNk0OMeesBGva5tM9msJ
pYFtp3b4IkdAByUOrEBQ7y4Hy72Vw4klFuCdm2kq8O8qzRDmzK6eQCidMH9IJKHm
gx79eIK6efy2efXozyokFS8yIBpurij2khuLTw38FPvwLPmYPdkuEvwdvKoruT6H
g3bfMI7CTXLXDx8lyaL/3Zech+Pa4ckluZXWdBDyBCldvR5wi2dolx20kbZmtpkZ
SKAk7+ZTdKyacKzlEfEMPXToSbQzVp782gEfMsl/Ku3o6WdfIbupD+dfoE2Thilg
FahZWNd1E3pZIHxBpfnJN2epHl/Grs5gRXcI20wD5q2WGrW0eG8kpKXsXmvbFmMU
ay4aRq1uHa4rHQhGDkdHsnHEoCl4HySKAolar62mpEz2WBX/FXz3o69Z7P4sjJ05
fe7o/P+cm74+U6YJL6zh2crGKO5aMlWS7GNDEsjrxpEZGZ1nI6EpfkY9ZdEcj+9q
0KfJtyvEcTrxoSkch5+V1YugfGvqY0kVTbEaHgqDSZLEruUsuMWBxJeWjlrmtJFS
hiX1BjOn+Dg9hlCe0PaGCqNNl3NheFME8xmLz5JpO4Hu5+MvHqT8mTFnR9DDEvRS
HLe+iOJ2Ucup5or/0FuRagm+Xr/uOvLql6fz+V6m35LFn9oUEhqXf5+pF2LXcSee
aXf26t/75cN7P7WWuISOBlAJ+7scLYcqoPLkeg3sDBCSoy9QMUvWVNebJb6xPGEu
OMSVDOez/Cmfq5VRFO5bKIFPlfSYB1I1+MpO+yaShyACBNZU5JHbrPAH3MXyjyNI
eDAy4Gxjlxp55JzxHK03CGRW/miPUMNisZWdpEgKXq9pt7ipJUIsFENiC7UB9opO
VxDKho0eevYITwzl8fx5VxyFDoYOIanx+ZtD9tZ8mv8THKPku/RA9jFLqtKLbgyc
8odXCabTWEJ1lEZhBnD7otQdYGZLrl2TBKSfxrVv3W84mWV6x1JjyijoZgT/Ddpl
QeVeZEOZm+gB7qyDBrA6AtFx+zhyKOa4CU96OJqHG7RTQViOvO+QtuPZNJDKcEYa
/OEeM7JZDUdypiKwSjQIaeC7XgXDe/w3OKCXKLLNAJGzKLgh2r5/L+3tjWcYsG9k
Xr+w/99tAFx88KusBRwg5sJFsZDZJW5i1Mv5RHqBTiDes2UNmRE4fPLZc9K5Erq+
zPhZcVFxTyPQgHYK/AUaVy/yT2MxFvR+kSti2eBSxCKQKClLimTR5Q15lkCUtxi8
PzWm4D7j0PNVnTOff+tG8la1LxAglWA/zh7H9Gq9Tw+uZ+yUzfrtUjjOWuIBANHm
WkhzrRB8DYynfuTC+K/Bu7rL4aphxJ3NB6XMaCnUOYJIqX8bK8g5lYPyyvTfEHaI
ZJW1QFzK1O4GCMJnb7rYOFAXwoCG7yRRPS68myFP+cLt59tMQv/AFHzGbOI4/AxI
OhVl+wfe76rcwLtSMKXF+rojwBT9YDrP21glAgby3rCuTWJslEl7T2PBTpE3VwfY
VIuJm7mnauLJHz3iSSJTOAHZ8RlBFD/10aM2gJEbE7wlqvu+UCukVY6LGyzNc2N1
QEOBWUO4i7BTBN2dEqAPicgRrapzwXZf28u33sZVURzteyqVDc1t74KAmJBqa6ck
b4xy+su9YQ/IXWCIi55nCERwZKDFJElTad1i0dgkGWT8uHeUt5MSsN23pPTXI4t/
IlTiAhTLL4tCyO1S1qd2t76ouR0EdO64a8+7sn7Gj6dNSNwNrr56i/PGvDQOelon
TI7xKQnto4iVCtNbskE/k+n2VX7ls5uSWqGrINU81qOvDN2w/bMTeQTo32Xj2et4
eTDH2UVsJaevGu9WRNMkN0JR+iHJwyELHYR1qn5URXddO0BzguP6J7q7xmGCGzTs
8oWfz0HHqs3lH4zZl9cJfRgKcnIBcLEYp4md9FopdLK2FvYG4mUprSdEftnscbpv
9akD9ZHr1KvHRJ6eC7/IpMb9X1kl5+B3+KT7TWeBbv0abfpox9sh3E9jocAu72dy
2zTAvA1bJB//BYrT3rV2I7t2Owxetv/B+l0iYE8AaczLP4W+BdC+qUvbLMWwCK38
fIv9BzYfF08bXG/pdeN3cPuZi8HthjAN82P0eLJy9WuECflxyd71dP2YL3eZw0MO
Zl7lfNdytsLGwKawJuE+WfxXJt55/Qi908AEi5QnaJViS4Gey+dLU44nH2xVrnvN
2IeD8QRpORKOnJgnkXPo7rfDCudy7uHe0whJpV712duXV8A79N1TMwBbJF/T2IU1
Vbdpl8seDTZx8C6LWN2FsNpFvBPf+7mypRwSnVaO1afeyxk3A1gRvb7FwKCd0NQH
bQ4QiQW6cr4BSycMLixmmp8lOUm7ww7UYR6iGkU5fxNcQXDn7mbACQ1FVehxwwUw
c+L2lQDscHRxhShVMb49hpsyADeN3HxXc+LiuzqVAfDgMBz/NEVWRx6hIGrtbjso
DJSBWtnu7kBj0EvGd6U8KP8feuS3EiN6XEAf3L0gOpr2ZGYLrCFdWZC1xp6kftr6
VnByrMwMc5/9Yr/YRkAPqNoqFhD0c8srfasdEjN1OBR/NLC47uqg7PBz/IfeYhHg
sfSkVpI/YBJ2eWS56JiCl78bAmO49CRmQxdSjNTlmbA0jHwbXkWRlB88LYNekQRK
3FuG3O3+NKW1G3cKLjsuPZTjIWHmDKmcuI17DQInwPxgBCYp7HcJlMfrzuFLH/th
z16AESRQgHFit4PaM/pc3qRMW55tsEbCDFPQVcH+8rLc+MhHu3RQpd5ibJ+lr73p
VkeyPovC3lRdPjhT2bR4BDX2ol2fWRGmy3t57+ujY8K6mqR2nsP7xyZDNEDyY826
8vop8MVHB831gaMLvNbf6kR0pkp/xnLL/Y9SrkNsSYtzMggH/B6dsK+supP3yIh3
LHRHku/H6kHaXvFSg6VbE9Wh5BSw6SYX0SWX9tYzyvAmIksE4BE2KXfAJm8UrJ5E
J9/dCLIYSnHhLGciaWZd+0ddhshm4rb7PrPj3bB84ueNKTzsu5LMDgkkhEnkQI6k
OSvWvcVP/56LXb/9WjO1SuphUTFZohRyxXcSaIAC5eeGNeDdHCsPKltH9gGMiPmA
/Wuanzv2qHh4ICmqwroDbfx2z1mrEvrz9UQKCeAbeE/9+XAOi0xcS80Q0bAEx/Z3
BErPLgQ4oYu5yFj6UYIFHlc3IB40y1Deg7xMwk+20LmM2eiDl86Vs9amyhjwT5Fw
B3yhRTvs0oRW0abXqBejjfzY5+2d2MCL3+0ca6M1wrYLgikUXZCZLBCbsdVUN4MJ
qUrEjNtr0QC331QAgDwVDHQtPX5gSojJ9CnDhx/oqTGsPZ1IrLcTf91p5t1HBJ5k
jiakXnGHZh+wrlzw4cRAPFsxLXEVXiw4CZlXhY9HyjmmQLj62IMjvDcr2tfGAots
YWs/JrRSjZbCn5ljGPDhJgI/GvnY7/pVzhxOMrh/h44Ht/Chwr8utE3I5YUjTAb/
OoWKySlgqQKijORGmVSgrfgVZTqFko6u6GcoZGwMmJE3fZOefdFxmgj7jeCvr3wf
Rf19+23VcmU7BJGTcXX7OlaYZlo/cWIHobN6Am4e1S4oqxYwucG77rFfRyb6rjFM
MT8IoIKkKmkLJ9qdMN/b0JBi0HR2wd4Q75Sj/uTBJFPTHRV0fgIoEoyFBGnXIho8
6JBx+HRzso40Ee/Ldq/nUfUhcgKIHyEij3wXP39EhVa3nRSYz5NIb3Iz4iyb7BSq
WmOxD0MgrYm93By0x/OKOfWJGpeLau7ytoHf5zPhEPn+22fvhzugVuWIHjAaQLbt
3HjJukQPmX+R1irLcpVRH2DXyzNCyPg4QqBcCP5o7BHXqxTTAJW+UTvPNt0GBYL3
4SQAYL25IHSRoa9/KYkTzHRBFUamgyznaWAMKnLqSGEFb4TP1vTSNeLadBtTvMHL
9Cd90ppxLZsaRaijR9zPzvzkJ+7BAdx9gk/+Y0gMjSKlc8qa3lHdwM5tmjYS9tmK
R+oq6glRUXJkQVIa2t3lZ7dfuZmPOh77QcFmeH+EeAjM1lWgZi1krEdyfOOn9cHP
9PqxoIR7Dsoa39XrAuv+i7m7noMlxVghfs5fMMWiEMa/ofW1opWPcqo/rQVo3deN
MZm8+ZI8NhACQWJHxAyD3d4G5nWhc7pKF4nTmidg2jfJeO968yyGIHyrd1uXsobv
3mRC7NDTfYzV0mh4bmXN1iBsT6wz9vOxobucknrycc5EPeyUAO+yRN6JyvHUgc0O
bHoJll8mfy2v5zR3Pag6ebze5Yv4FSi6/zAGuhghhSQVqYvxRl3lGFtdAseCy2Bd
hoXNg1zaxXl1STxdlDmBTQCbaY90ERWQLfilAQcP1ZtN0Ok7oCNG6pnkgke1W98+
Hx9KQduxtwHVkSIwnSoG0p9+njv3R+lyG89aSetZFXDTvEgGb+PMiY/fkjKlQ7Zh
DMcVm6Srap3tWQgNZxTYMyQq2D5QvPGLKM5aGKxlg7+9+6KmH2ik66Ix/ekB3WOQ
hez6AuSfM8hBnfRcyYejEp1ABwY1Z/8sqa9EsvtoMwJmuMTjq2UCQ9ETT6tja+Cr
mXqavx8L4RmqL4ccmTFXUILp51oCr4CTk/Bx66xHBlf8GHMiuGZLQpeCqC8C+wjF
hVRT6QwJZwb7E0DPJT2AGz8RQipusNrSW5bYRHL1i2Y0wFipbwlnZkopcqJgyDUy
DIm/GzNsSruTsUtWYRP0kPRwni4kjz9m1rGa9XCY8m7d1WVMX7teV1gGZrcygx/n
V0EvP/I3WEXU+cY94j+SykPmOW8NjzmaVBjnLiRpIK+H1NTcIE+MXzRpwJiDHh36
2R/Xy4TvXVt2y+uDTgbRQd/THMMqZgdvyTay9sNliU9T5czfL5xWP2yK+gSX4tKG
IP/Yk3RGu7BOk+bPAFbFiUAgVmmJ5PFIZ5uBhjZmJO6dH04wABgwyZ519hHzXSaz
jR5xxnzOdgb1+j2TuFJqoT/jFyj1iyMkAyq5JnxnJkzQytW9W9Gp1N5p4SXzsaWD
mIvadUWGXRsMA8ADn3CT1EXih6rnzA6s43YmOCBi5MTA+EyVHTKBO6r1RlfXw+B/
RKHUbFWRtgBtznr8oTUn1o4RTyhpIwOJblWj/zlzwh4TCCXfR8yuuF41LCV5Jbg9
o07GXA5iO+ylewrIRze5T9YUzHu8cK61CY4BwUKQ9vhTFD0ovXyLrnpeNli0Ac7+
lZ9ftfbKRyZxT+q7ZDvxbjwWaBNBsztDFXKp84g4F4zEvLNmNH8NjY+PFGNBXShT
UQrGk6n2GfWSDHPjaT6tpteZ8kHRN035SGgIHtYfzI8R/PbyFEbQElXgno+WCt7G
G6oB3HULGWt5NI/W+tPtmc0bkEMCE+howwZ47Uevbn3gYLeD+/AsWhT5RaiUMWjQ
fLy+gbQND+SDUaowaZaEqWuINoaWZNGQIBSASk+wf27aoGvDYghtdUqsX+/de/BJ
hs8BPKzcrnrTDh9XM87hgRL2pmGd3U8hITPCIJF6jEJs7ERAhw67Yau2HDv5GPH0
eX/0rzVrnwFqwi8xxNRO4JpV3Czuk2JLJKOOV2m1w6Vk63hf21HeaDYLyI6/auUW
qedtRztmUcaENEZNauye8BScB119v8SCqZeDntsVmez5Fa6yswJGpGEbZ/oZmU0q
kFWrKFsLtLKWw27ARR9f8TWf+oYHRCtRPyrJQ5mBusoNNeDJ1FpLqq7L4cXAD5BO
etsP/hSeNwpaNZGD+gu1MCg0qtXlSeJSBb06Fi3POBylIyq9WQpz+ATmb9AEfCCh
OTfSX9h8cFjPhSXeBJBCsDK0qa9bdWeC/Fgi8EKcFITQbQ1LtpMfFwekImEsJG1t
DoTTXkbsozlVP1LdDIqrr5SlV6FE9ep1E0vFiLO1M2dZf6sMywtcjAbNljdyz0Iz
tS8GCecbIhunsLlxnKSReqXtMc/SgHrmhflYQU2Gfqlt366YOviVQObaUBUp47Ou
09BJt6xHKCBkBVguVGL5e87+TpQLX3VVp1Zo1EsfngAuPSYqVS50OkiQ7f5IeJgC
5p0l2PjCJg9TyumoODfUY9/wTZaYFevrTRmuQMX7By7fOewnPNppID/Geb843sdE
XqMTB5+02Q9P6sAklBsbrusET2+c5ybsAoPaomzSdzPC3/uGTDz09t82RVcPbz63
wx5cXRDaUkbDqGyO+ZASt0bqR91FopQPqvOAlxrz71KMcjly3tMACAN7HlyeUXa7
hyd35JjyE40E2a84WmFL3TWaxU2e9j9xaueiClLkZzkm9IP7eZca1j86xnKdsQYR
HOiqaZUdsZMxx6uapWF8Aho50qY+DOSWiM7ESfOHUuzw1qKRgWL+Ma8Ft4cbNTOR
LsUBdQDPDeb+vr7jsSj6ttB2gVn0PaI+EvVPAXBGHH6j+HA+OgwVFInddHxd0nnZ
2ypruBMUp+DMmjqgSpSJJJfK2eA9RuxsrzZj1EZsNXeBdvnefuQrpF+sD8D42/z4
PZrALaFjneumQfokHRfryyIDaqbyoiftCVQ1BP851rda7LchIONjF/3DASlgN01F
r/SMcLW8jZ1OJV9KOwX3LRoDqWeb/77pNPWd+pJ+KhbsebkKDFcxWfBCBOhZno+W
7mhPjz0XENyrTGME9hS6stHfNXN6lAalOFv054IWG0CEnMMHlrhc/HbZP0/ENBom
fQxdz6WA7AiPyT1Vec4PCX6Rssg5CN6hUNNplSY5nmbf0XVuH/0jK3FA/XjvtgoL
Se+XQEijolQLDefVOz0IP/9kk8vZGiBlsr7C26/jWGl2BH+B30V71/ep8syBz5sA
WBGb9qtY9yvTQ2llStFOwBTnSKAJikP9WjysyavcIeI3Ww8TediSkLa7c98GvDvt
ymp0jhfKeKwN9vRzpknba5w7TuRmgBIiIiPWq2O5yX79b0n/PNLW/ZlxAFqkZz1G
6rCmFkqacsTyn9J7wGPE9rTv1qKUGAPG59mXw6TcSHbFrHSqNolH1TvF/kuAEvZu
VdE8qCs2O57V/9pugKzDcULt0OIuO3gEVX2tjoWv34v1VMqi3KFjyLE8Lo2YJmcW
YzNtbYsZuXQrK/VKlpG52Rea64lslIJrix1AfWRYLenvU5oMbhsVVro41XVdL5JZ
8asktNPKvtfDZL3kmhIECI7qO9VjwQWItG76WdppjxrRedWAkqYG0ZmF59UOU6Gb
RDNrwqRmSdiv2vFU+CFPBm8xAqWUjHVWcmuNU6d3OTY2Bv3B0edW4zBTByjIx3i/
wLR4rQ+tiy1xfsajtbPdjvbKt6vT4l7tmuWt8ZlAMAbGQeH33IZILrUlytQgs89f
hOxvLmMH4Gq8zAkNxluJ1MUsdiF8X8v4bD2Xko9aJNzT1H1E4X4i+Ew4Q3Gujs6m
wlv69NgP1PPVAcO9Itw8OYzGuy3WqYzi1XghRKYRbfHgn0QQGY+1MZh+UO2UArHF
J7uac8UsDjknXDEt5OHsRZqwo95Z6F5p7DlVUiL9a83Xg+0VT393o/ze7bn803bx
nDFWDzmg/Aoa75LVy8Cn8eYN8Qz0wOVjRGhYXRPqghEgx7YdVeqdqbMaDIGfUURN
qyGDlJzs2a9T3PXM6RGaAJrkcd7mmSZL9Xuwb2HGuj4cDM06257huu3O4tQ78y6g
uCmpI1SnMZpsCawZF1vbXVOaHjVGr5n+dIKcCHxcsv1elQ1ZwixlY55DE1/6PxD3
u9ohN/XdteVGYCT7ld2p3a40CKHkYGpFoyXhCJVaTQYZ/BMQ3PNRDMsQmAnGYQZS
YhVa4LmpkNFFaUOTJK47+RJaY5akJyPGeC6EYimJyCAQiahUvqfn+GnMEk493ufW
3Iiy94RkBc2jLBdqiicougiU2eQQrXAB1vs+l0MdpBes1ll59V3izw3rgWy3zsEb
MSUDzd9yqBgzfXR/c0qjGtGzjgYilbcxW8wfCobtAR71DamPkbQz0bnlJ26VXkdW
r64ars4A3OBJPCSg6QZQcy31Ln4dzCqbp1rrD9hz0e/A08GWEAzojAXRAiDG9SVf
sIilAXPriVQz8Waao6pPaAyl0KV479gGg8GRwu9lNVUBp5VcT3hNadm58fZiZ21a
NoM93Zwfn4lrFaN46pyvDGRSEhNDVOSsosb7ei7ebuj4fg/s5PHfo7GotTUUvk79
rmFhBRQwk0hEXMZKuueatiSdw74Qi7yqRbI+rhrIF18He6HndC/hpd2c09gRQGV9
i2PBav+VJW1GVdDs9tVcvaYDBF+pstay9DENq+3rw0/LBQvfPTsbVRAWtDTthm3L
S4ITMFltyrEr7YLKjrrmGcHdwDqxpkxYJ+OrP/b0uWexy4KHeSY9e6RqcIKmlw/B
gFV/+/BPsOpK0WuDhGhcqPhbMrwv7kZLMSRXDVietbbCdy6vkbfBvUwZ+Yqtw4fJ
bwk26fKgiwIEgtynArLoZ6Dx8gqOMhBQetDf/+eotbGSUJ8JUZxjyvNRMsk/TPOg
TCut86UlGd/ao56aF/JyU13WjoU2U9Dpa4jVVrodoC9F7Lhqho5SmnBsUvDK2Na5
34eSatyXbyknMUct6PueyL6w0kHU0R8YEo+9tnndjiGINO6l0ktVLuxHhA7wuhIy
Puvibw2MJUGbpWxqmccLuMbWnUJWIzZap2Ij8AWJiR8zcsWXO+bHhGAzawsrOL2N
jvnWjjYLNWwn71Y58gWHV7d7deybzoW/IJE3XHLTJ+ojGCd6q2tvYP71gxwiH8Be
OI/NwEUb7z4Y16ZEksMwodzVHMjVONZtKdgGnonSN0ugi684vIYzBm4hCIP8KhIl
NhohCMVPUo0dhSMDac9bDt7k14LcDbJgqRsbB4q9e+clJWYEk9jGeR3PSEOZISns
o6E4bIpWbgHdxPOf9+SIU/bcIuqjJcM/qLRttQxaLx0swoUMwRb/SLZTFmDogVK0
sBcPaehttDEn3w77R7yevnGSQmPRIyCOyRon3XsW4oL9/BFM6KPdEp7vYLi1h9sG
Cs/fLPT+sPee2Ewt0hOEVd4fyT6eRV6D/E4JAxI7gIWqzjExvAOikCKVFHNQmaPf
EN9Djfc4xJPZ2mRSey5pQiTttRXYnBxYzbpIVfqaBUjwwQYK5h2g4RMACWIfV4F+
I0V/zGx5JZxvNRtWxKR0Jga8SExeQ7/B1BTMRGf4U3LVWoKI8Qk3LnuV4nKwkYBC
VU7l8Zk+vGQXmL5gENERcWMWfr8bowJofRzxKbZ43PDBpikci322KmkSX40yFjvn
B8Ce1bL9QJWu7th1CINv7TAz+T7ZKS0RqFYK6oRwKqnezenQTPDXHxdzBc8UzWHH
Zbv1+Z5L65QCrYQ5G+APZOK5jhGMz4U6jT0rARNnt+rs89/ruVJdiTnpFn4Ze2U1
+WpuCkiqRDUqsGZ57fJyEQuoL/bpOrT6ePZ9Xeyy/8rdvVEgEpgHMF7MXp5Ksf/d
nWafGTUuxJSRIaabl9t3Kn6q3VHPjEwHbBmJcIo2J1MTT1dYed8sg2dfnMUycFjb
yXX7/m32pGGxKCyRfMpnMYlyJQeSOztuqn7AK2qNNMb6Apth4PieEv7rf7juSxHC
hnusI456puHIGFDENBWmh2zn4jAsUB6eRekRtokF9g7SmtvuT5tS7NDxExRABYTT
EwblrU5uPZKYDWdDNVdwH8R4qqEUeArvaZm16W45J7IAKDVCJfzuKK75RHtDHusi
BGLYFLajWZd6lM7yUXFaIk0bAguZrMuoEjrqVDtpLVut9xO3flDHFJ896AV3JNTS
b8dyN01u8zJ346kai+rKwPvjP+ylxayCyxOF6SEcdKVyQR1ZPS9Yje03YGrE+AAI
msOeGvnVvuIrSlFxBalLFzdcVu9AWOgfB24g3TW/kP+wJqGzac6aN8YlwlM+rtsp
bCjapJ6yRxS1uiPMZMvTtOzf0QwhNOeaQyvEy6BLJW4abRuHclqnFJF2z5Kr27K2
OZMyMeDDWDuwQ5vrX8ICPc73s8XedBPwHQVyhR00FnEESmzGMwnAqnOyR5NYONjK
CFwPkapk/wJ+u2uAs8LpjoIp295R+WRMFG9nOLoUXwpv536+3Z6nbl+Mj5VpsJtW
51yl1doAJM9sJE8VERdxzFe6stq9JnW/2pVYSEtkWoBFfkeMNWCsDUjQGbkIwtcL
QseSrc9lX+aAyXdn5w2LFIZ07d9SblNb5QUv44pfZyZYQCgVEsv6xDWz4Tk9S/2S
/mhxht+ZZCVYldcuW0PUjcyQwOMaTeFd70qff9h4FrDWa5Ivol2WR6kD8iIm8LTP
2usBDyX0CTfdVWASxfUgiezWrMnYJZ0P/ndf4M64V8tcHoJsVhCD3MxRlfbbKLjW
PLKeBdnjCAd1bxQEt/mZzBxhOFBysV775NwuJIr0Mb/OtEGW2GZLiLZcz4tJIZRC
ZwNwag4wExaflTcPtJhZr68c0vdcGRt0YXeCAcOOXVimBtmWPIh8zSsTcfM2dJzn
lDEohQkUXjTQe1nAwnhaXnQehKxS+A1GmkPpbp3G3VNt2MuWRIKu46kRoRw0SemP
5lJ50R08cS4FbEDCR+u/EpBJs8EYp4jmnYaUS0//9z1b7LQ0Y/MPh06iKmmi8eZK
lB2p36wvEZomszTlW9YU0YaoOJ9ohmLBMfeaUuwfMZEBCluTePM8S2IDcif5kXjy
M7/B0dMrhCXhrKacRCu1FG6BbJKkNBdSdl4ZZWuf/q/IOcFKqlLniK96HbJWxo0q
/aDWCiYOXo4fg5dghXN+QpowwKOU8fUx71sdL7YCcK+BZyYZy4PtXP0n70VLiCIL
B8vVGjPOeOaJ2VOZea7OWNnhgI/s7AZJioFt/5rpVAI9GqsMUzw3x5waHJn7MQ0P
o5b/lh2lV3JaYp7REg6o8jCU5HJdnQdJ4tuKxshRc4ViNvQxPlegrQbvP+37lGYw
W36Gt+3R6TI+S9ErXAAsintt9PXa2U7RqNqhJdGNItFouktf37ZdeAjMSF5ptfLe
sItH/dk1zVBok5iXSZMRUGbRLJYW5HhGimv9Jq8W6irSbdIrJA30iatGI+B5sbUZ
UY6a+isoowsK7LXkYvhK7H2yZjM8I4luGlWtYgcT2fCEgB98+FMjJ4oB5AuFiUuj
8Deq3jKC8EBOf0eg/SfO/vACEqxazIz1TmLRUzessVTY3PJ/cN5V9bj0nNwjlbnh
PDTMWKa/ombp459xmQmcK3cJfjMkpLyCAoCfXrgWrS+T59bBAFohElD0K2hO659Y
XLR42gTIO4ajErKqf2qUzfJkeNOOoiicIAVNSO1eaKWKOQ9vc675QCW09MlOD8t3
hqvXsU50H5nAjbdPTsw8npJ8Agcrbb3Ai+N8B9BxZaTy/1haTAArYJshw1uR6Iq2
cksHXB6VSLk3xVIj6abdH4yiAxOLFGsAbuuBS9NtCnOat7fXmWplBKM2T+Tp7okO
0JgjDibxPcENiNA4NYVBcVFw3BHercsUSBLKwKNt3sMDH918rpLSqAY4YPm0jeIg
63bkySgOsPmeLkl6tQJWdDjXLv+Nl0V1cyUhyUdBqYwXBrKXRcmFg6mEMRfgNbUv
+CC+K/QHkV8pYbQOprYhVGtJtnP3e8hLUt5N6FuBVNqLhgwdt+Sn7Vq+xUDesGyx
1NeHcH3AASej9XeuMOnxj0yK7+7ldWCGIlGrT/iQNxh4lAZO8OS7EWA2OOu+vUHW
YyGREk0iwAWH53cIAYFG96z7ZV8xjKHM/+0X+YQUvTudu3r8KWZsHJl8LQ3FnS8W
11d/fAV8eC3kPsZ3la1++8bIYCG97x+YPZtDDftTbdgaIKeXQSwMz3CgmCqYPVCm
v8SSy0qJPG2fveWokrVBUq324XV2FUPvvilRCOkWhEHvZdJj9wxfqeZKipJyt6ei
vu2/UAZE/8PuP0hd3aLKnAgxjrcofyDTHEnSYRlSS6lJXj4sFHJ+rLCodCsoQSjI
QmJDbqaXwmeZWEY+rDvi6JWcpb2a4bgapkWf+H69gXfg+fHXoaqqrtx1auAAcnVK
UhBj+DnOY1UvhF7qaq3e1iMRx+4mtsMLSq+zK0EKrO2LpuSGwQvCF9Cxi1tBZY8Z
dAseaVRGftu/a2jpyrmz7nAv+xH06zN6XpBiPk0OmagvP+KQu1SqjYvC5FcZFdfS
XzPfUm87iULiKtYNTcsUZZpLitcHnV222+0kx+Zp07Td8TjUESz7zFrj3ni/+U1I
7U0G2Utmemijrg5OBsKLulghGUbFCvaf4KWsCqBwp9aZXQShph7LESA06yGt7KNP
zHnOjZUyKUzuPrz9E2KY7cbJQ6MetbXLMiKL0WedBj4sMIpY6J0V5Fj971skLaYk
yUZgx50kdHiVcDkE/b51GU4kCDDtivnJEc8wX4cMNdGn4BAlWPWvNa9zfBoSAQTV
mpONlmZ4FVSkyVcD9qbc1Koobg8mcBUiONg7jwJsaerlXZi+VNFniE7UexwD62vF
zrTZnk62U7ozZRQt6F5uA/cij6CPTj03DZyXLUQXX41Rkk7H+TU6O9dW3MSOwLCc
g4hUX8aGHs519oEMhOFBL3JJYIgR7YOJ8REeJapsQDn34IbL6bxDS6yOGmez7lAQ
DwUFvdD0pyFukPJSDedRkmR9wEZa2x8vu7sb0+KTSw2jOAeKPKe7ztKNmmxdwrWA
G9khDbH44MKV6qNGpbMtgv9PhqlNmH432HcF3JWK49mcJq68uZ5a1WZN7JWpeO+X
BL9ZMYyRm3BUfpf04d8jhJSqAKN2dOsRcCMNXuHdtvVp+4/yudQ+I5giVW+S3tZc
kubeUcNL7cZsUi+Gi9IfZAolfRx3skbFw7YmJcfYFcG+wVSdBqbHzMNVcrZRdPtj
foMkUiCYZRwvAgMmVOXY56/bG5G31uSvjy0vRUnL+Sw2AN6EBIAF188CixVShMXe
OIPvbsBPrl/l2/tjRgec8xW9AxVweB4sZfPQBNb08Y6Y9jjR/0I07TbDmksySHFa
1av4w8CrLZW8/CA17iQmTbasoVh8NzUp5mpMKyfWyAg33lFs565uIcPBNOYsyBTp
WFqlE39zaEXVU/UqSOfk19CBGx6M8v0B1VwdpCVnDACpM8Gk36DWuFFZTxhBblcx
tmE7fETGvEz5vOPZDzNPVrRdzsIxEG9F7IVJqbQVOFo2uC/dtCaoRdz96gxfdYyz
E7HJ9R+qwa8YsHI63A5I2nxKEDYjeYPnie4sV9wcgC/vPo1pzbTxyhM9KniE3N31
cP3Pd/xcEwuZa4Ka6PeCR9SbMzTYPEpZLM1zASsViba1Zk4vQ6LCZZ8felHCJBIx
Un27dil/iDy07Fqmcs8WCw29L0bgkR8Oiz4FFwrg10XXQpaXmZ5f1D6XPWRqTLiY
jPwPJCJlMprPoK6ZtwCZbIm3VibW/B9BfMXiLkDfB2pDRf2UJ76CYA/gdjQqlL1O
Mw+OUVEcDyg7ZP32xi8vKOZrHeTGVUlIOHUidDEmsHrVYlxDOItnddAeOGCZ0VRb
tK62xZ03wmOMQBFJTMC4jfpmquougB+im77ztbkkk3XUAGuozsK3rZYkMWYwZvD6
zRoA9CU9/0ws8P5zrybju6aFixzBDrikUP63ndAWMKXAxih5MLa3S2SxsS7dDVt9
I3fJQ1oxxtSHxeUM36S1PkL89wWGFXB18IsACq4hXZII7CaLuwwQIE9MD271815P
ZpGmiexpp0aq0swLQsknuKYiqKDuDSiH2kdobljW1MuT9jN8+ISfhLxDbepJ3fcO
wmD9+0YFizDoTLSrcg7mc0d1LxAew5e6KMstcSb2ZDort3CqOHCSkNgc0+ZQlZXB
UpntXHlAu0343pHDOu2L4Bo+tANZ0rNVy/6sWya7vy3XxxJatR3qO4aYdpeh5/4C
m+hqxCzl7OS7eCtPk0lqUIPqE0+HkL/NUYq8P8WlX7Hcn25Ps75rL4CYkBoTarZY
V8XnYuxGKMl79eJIizVtV8jtVHJyvv9HruO78vfSgSHWNkza3P72152qdQaY8sQj
ouvaiCjiaxNTMHPFkssUPSjM+nIUNUv9cfuMWurYtZjh+EwuiSy6meM8gcv6zRP1
M78DQctztIrVwKxcfakT8lVJqk/i4w2viPf5gaGabaN7c348EGKf5FO65lUmoL+i
53uYiD1c3PeLSI6L9Hh3dh0Q/5/nVYjnbXwABsruY7AH2FrtGP1rs/9IOx18Q2jz
kQibzLYcfCY5WQQS9aQ+HLGGfC00Pm1+GVSkW2uzA65q4NLB5zSQnpSsgNNwnk91
37Fiwb4Ro+SIyhsAWRwbXx2tfDt4PHK68Z2FOTGWYlsfjgk89OlqKuyNNlClL7h5
coYa2QbMMoadAor4DzSStgm/P3f9amLxHf7YFaehg/2gQvPIB7HHF4JO6E803alt
GByqv7LcLa4UNOSTpPfHkxNdgK73uPCUEIRNhtT/QuC+D80GbIeQu/31FU7SD/sC
meAdnz9nS0OJ2QRBvNZI3nCxTkRrwoJmugbvNSdg+RlnAteJwKP8nu9gy2wbW6Sn
hqKxrsSa2FAcWNazo4ENre6IwrkoyD6vpsbibFMI3YKYvupCSealGgqzZV2zIOXI
UEJZ2uvnWX45kSTHo7wrTgfEnFFtzhQuUXIPUs8HKeemySgx4N4NCd3eJPQB4njs
taAHrSthucqtecAyLIe9RwamPgmrpWsJpYhx8Az0OjIzjhramj2CbOWN8x2SsMNg
z3tUcJ4VxaVvi87ihIp4MB4d5tl2nAe33BuN9tKdveuzwoxEP2643yPEcasxWEax
R4RGtNA9YwNHOQD9cra6mrIJtRxe3sPRb5c6lKPrhJh6g0KTXriKANMdDyfvjXes
wx0pYOUwIOIlcYT59cWW27ddvhkSrx6XF4HEdx3urkpgWM3DJOZ8Cb1lKDrpiJmQ
vEalJzH3D5O4NicwA2ciIj4uDxenPuufUN+sv3TzhSkccvmutlPtn9jiLaNgt5+J
Y1HOyJWJCzLnzmGqCAjeueZIJESfT+KykeH86yryAioG6n/MfJkIPDZMNC7/MX4h
ro1xKNPZEJZAweC4V7ps30eLakBJNpLi4iqO/Zrssw6/pQUgYP1amaQeR98xaWpW
s0NhDM2Mf93fUCuOAyzKk+vKW45WeIe7fNxcgqo3DvFycjVcVAVGOruj2p712zMI
zaR1mNQ/kdsZp4+filJeZRBTyG1FYP9IURHuNxwEv59iKMAQlJ+wo7qqkTG1QWiZ
1e2oBn8R5dF8wsOBkI/YLUOuaUkCmM51SXOii5GYv3qWoM2+2L71EoJbVO2zlh2f
tUjbPdEB4xKhHrRtAEFBNBaDZZgHgZSyDH6KKjNUqQ7kPwzHSDmL3IA8fT48a6HC
kS9roJ9wJN+9UAPEhxe3+w9e++UYRMe3uG2IwwRNtjt7TQq3d6n1v6Bye7z353ON
6eyLAji+IT/RnWR4jfmJDg0zQ05A6vHysAI7IFoOZaBi4YKXwLS0ebjCrFXtpDRa
miwD5Ru3xDZBA8sngWNhGPNhwyK6Ql8WYeixnMhb2HD17Q+gKlqj6mcQ1Yc/rvF2
ErkE4h35W5OPNHTaYy7YyyUYgAvadJZt8C2IpvQYD6z7F7ZbifVquyTvzoYa+ueX
u0iiHzmTuYo/lNuFIMxTGZ4eLAMWA7TD6Cj45xjds73pdE8MSBSgzJVsEv1RVt56
u+P1z79tNyO4Z9NWFvFcHNJta+kHMNlxPprfj0i/uF9j+tdEsyC6lS+uOkJykicT
i4I77a8PuSbQVuQT2LyHTUqHY2Nn320LHMOyqB3NCmps6w0jRN0MTDanIYOvO0Zp
WEbaxZJfEguaXLnTjHdK0PdJylwHg9Jl3AX/9Cu3jhY5y09zmupOevM+mMK8RgCh
WO75uBk8Tpc1j0sYj6w/yVspOEv7ac/8ecXnMo3jlhAHhemzboMMY0TYK30vr3Wb
626eQtaBhZWMRsTNJH5mqKFjdXUpn4kTAhJ8i8CYZhbqIbehWWWkMwS48gYTIW3s
TtJVXYrqYjnuDgKsYtA4o4Df6NBWPT8ggEVszOJszgzACv+tRTvBw3+vQB57ALhC
nd00imy3XtPN3XMKG7bH6BDgpvxLUHKw5mOpmRF1BasogV29dHa5rqyo4m0i0ocS
UwGmf8vFooF4pAZWPmWsnhS7qmhFJ22zgMcqgPcW0jnEusXmRq4c3Nmv+2uMZOhC
IyUgSTOGhQQ8kstJN8JGPXsUKq6ZIDp6WFZht9fuLrvK+wnOGMQaDWFx3ac9nTa7
bhsIdOgQIFRJbZqHLFRCjGyfOF7AztgGTgGDrpdvNEWxH49frjurLow0rh/TGcZn
NaZmJbOW+twhRklv0nE+ZKywnGoFw8gCC3oJWuGwrfS5WEnWDmwgPrkwvUuNdnrX
M+gqDpUIOFD/7QrO9oHa0Mgrn3G+LWqV9M5pljeDaWgkrYx6RqY2lhn1Wv1q8f26
kBrwFwC96ECS3EnzxQx8uo9VYqTE/4UR/AnIdN/3CMEIKvAU5u5Y7bZcf9MWkPAn
/OhGowkA5XqzjN/kdHWGlJzfaUdOYhKmXPae4HNoMfJjbFUwv4O/u+l7tUGdnixj
4Q1pWUmmSK5QjjVe2eYxTWRfPfinEAPhQLMwL9EWoZPjvO69bhfU2lPDcvTXGM7q
lhQfZVXJw8GiZO4wdbLYVNyugdzovHfDIHue+v0t9ZuvvyT7CW6gtYOqddnNmZ99
OKTUmhWUrUvaYr1JcHKMc9XcDpc0TAELKBJVeEbXYi+J5x/3KI0M9VQQKx6VPq2V
9lWIZQxr066epsqCsaV9rHbdV9IU4L7QtB1wmuSIAeGb5wU4Juw5MaT7tUyq5ztY
9BH2TBU6vPIYjb0ov+fJp1M46W+o9oLdraOSZdWjVuAVD7/N+nVtzSYSeAuoUsdU
mS/tHzLxPZJE1sh/0I5wWtpROc1+EWmoPxtB0rJESscaSGyYSZ9j8WlGwuGO1zIg
2Hamu9hyATYbIsfAxLfSP9KuPHO5A92L/I9U8loZ6/SHMOBAopRAIh2A5KwLccxO
RwtO4wrwa0gC2Q6phBzNCtPMa3B0AHjkSRJaI0VebpwYGTgGDkit5uVhaEBjya5I
KtkmiKPE8YGOIbBwMfgRPiQhM0VEqgZ4r2y87fP53E/Xcr/1BE488YOxs/9S3J/d
ZHS+TrVXwq0fR06mNlrf0oh4CWDHRaNlJSiOLsZC6yEFIIrMQ3GwkWF8VuvxlaDN
3ZIA+FKWQ+3VTsHzDLLmL+fBLnRsiyaWyayAGTWz75nOvjgICynPoe91vWkVoiiJ
xNMG9M3n9FmsMVanjNT3M5QZREVxHABYpiZR09/k/o1Ay6hsq8yOjnqxtj/D81Mi
BQUIOTn49xkM7uO/AdMTJawwUvE/wDrtHfM+ltook7h0B1+ya7pkn2VxBRhXO8tD
apTabREPFG5dCi1Pt1QAhajppqqJJEuJTyAAFILgPJu7DuYG7OEo113xuHQDfX8S
G2nxX/neBx15LSps4z+pNcPeLuFmZEJ68yhcmqkperMcaRHpSZt+yDgm2FwGdl5Q
/tcp11MtZ3jVWFPjYSpLcHW8VTaIIeUA85UIRU6AjOdmVzUvWK/cpH31IvTonSXg
jI6CHYAkmLvg64FsOOXYZ1fzxO/gG3cHwaAAZ9XsoWFb6TDuqg4TYYSp9oW8+37Y
erasbmO+p5ZiMT/pecmNYeCri5Kt8vupEeHQEC606u5NVML4uxmxU8kOQ4ytKmAl
t3Evzmrqu6GPEjK3gWKhCsZjmG5zh3+4TyDQtmLyOYN6qge5llPNei6zJoGDcAa1
oj756/jev9zqoGYLN5Z1BFLB/k8vhcTQGcJhK43SERRkyozzwGmkTCQmIpxfMcqQ
uDxSpRo0rHD3D2rExmDs83qmG9ybIOAq4CLlVHHCKu2z9vMaB38kqXNsIK34ernE
cfvQ5V6Dt2B+pbN2FPcouGsdBx/oSy2JQO9LFnVm7shH8ia8O6wkKnIQ8WmgzRJ7
JTO8ePrhCAaUELL3gWBeYnFXz0L21FGFSKw5tDvqV111wHqIeZmhtBRuU6KhHZee
ok3Dwe8MpnvRId5u0ikB0ex3CNVCkLbC6nfi0q5/IErv10LA/yjzl+eQ6Hv8QrSP
2S7NJIlZ9oBFbXjGIFkSq2qo2Q54+e4j0dMfHGQhIjoIo5yobuc4iNxLrSJORwOU
8Jwn+/1yz8CqAH8tUAX1SreeT3xiXoRdwUeAqZD/Te4E210aA6jlSvMz+i3yNBiS
qqg69WQlBjsj+HBWdWIhwgMNynjE+DW6zRxYqulaCi+R74QXbMkDNyXg8/VWagFe
9eLoz39qJK8hiVWxv44amhIYia5RQyU2g/ayS7EuAb1OLuX/+JerZfVGVSHQFUNY
jGyVBAooiMvuhLuXUIgJQ+lC7lx8ZVoeHoFagDX+yNZy+BL/0ShWwQmzPUkbwSRZ
eQCTpcuvMH8HdjXFFN1fvBNR4Ebh1ohFGGx8EKP1mzMA1JkWlY7CCeLTAYgRWli0
YkDMi02C5giWD+aXXF28bwWhGOo1b2QQUGvtYlaLtTzrissm/w2gQJrIocT1Lc/B
96sjIHuCH2Z6c5DtmXgbdBXyhDgACXLH1875yvUvlDoYF7o2lgcpyrgWRphPL2Yb
G7DF8zbdU87ZeEqNct7xoVH49zhSOpOU8WuPf1Wx6zoVBmhEMgTYmnHRQSCe/ueI
MxGMMmCZxk4kxCnMXw8cT8wml2Aw+iqOgWBbrVpr2nAiqz1V2J0aSYhEL5AFN2/Y
NW6DZF29yslb84z7B1+h//P+k1fGvB2niiFCxoNrEV7nOGU6NAxUlgoalj4f2Scd
iIGBoK25pp+iW/oLGgbXJHjUBAz05LrTa8AJlhNfyF5zNr91o6DbDcUpbCm+9sJK
bOSrBlngMkTuYdb2yHl5TmQAVVIvVr5ox+aAWc0uxiMItGq1FEEtfo1M6Ji698AQ
AXtgav8A/P7glkkSEcTRmzQx8h963SpbQTMslwOZoFiXcF0SXFbK8R88ExjFmq7y
duce7ey06l6Fn4kJZA2qarqOD0sP8PYdp0yohJWT4w+VscphBwq3832xKJU2Q7Ea
lxHI4kgtt4rwHcOGDO6gJXfVtCrcTH0Ep6cE7/6l4e3250f2Ed6LqR5qYCJjpQDY
3DDrwf6P3w2b+FOlN85eLy+dJqZPnyaZD97dBZMlzOYfnGoNiiXFWTn2vcz5mTOh
Il9uY0garCt/y0K5MtYA68jU5KbN+qRf81CNM19LYcGbUX6g/yWRm3dwGlGNGYtd
CTy2TjOBf7IwLbHCNUcfAef48Y0UZ99pT3pspLsFu7F5tIBhDeJUoJ9Ap0K3hhBd
IVWOxpC2uINp6UWNx4PMmRjWKVWmj/uNm1eukiAIxv3An6u5kAe/QIhLZ5V6L2fh
HJo/HUre/EPQXj/M9CvmrL4ovaoiNFI/u5e3ExzJYXZbB8t3JSGGORiIGfaCz+/i
Vv0WA+q4fnsPsX2JWdogDVgUhXA3yzfvuVqYUJUAUi2AhvwrXtgu+3vtSUILg2je
3lBNi/U0xPFyd7ZV/DctkpmymoZ2NPxj5ZMV4piF31UulCPgkb2Uvk3nZuTDm4Kw
TeHxej50p5VGq/ZczyKEaFZdevEGBaIpb7hXcvTI78lvRuT9FqwQV/NV9OswBW+2
XAlnD1DrA/Jl4NF0CSNwEoVz670ZZArkqgsY2DU+mv6bQTwjjRB+4OGb6HPoRWVo
wTlBxpnRxSTRS1CiQqIW7qwjyqQaKXT84jgXi0zn4qiy/paCmMcsnEE2R945XgsA
37BQupIZg752xHvNV+Wfvrf8ZM8PER0yuyPUcNhX7DYvrJborhp8eCXLSA/5g8w3
0x79wR77AK4FpVNve0hDzvhquFAOGtirYHIxGDhfGr1+YwIJXJhrSYI5xTkKtQwQ
9gCTE20wU7QJ09fwAPhbidMIbpMV24c09iPJg5fgnfIZKD6bEsUDjZnd6PO/rREh
IV6c6Esy1TSQV+HzixTYWHf4urRCgfUr/kEEjnXDAK1pRkxbaNiYEyqT0viTtVrn
o7UmcLCStQz6TVSKHQXNJIVUC35isTDAq5C75kvLM6qR5UodkA+S5hmXMYMFPTdY
jrkuKvbHqU0Gt61lPwQA2lPWfJVox+ZdgnrnQPMF5FXhe8kBli7Lf9dPX+07jT6n
fF7vTvZaGKgLU77tIObE2HOLrkugh1eOPswjPVR0SaNVlNp1swrQxWoih7Ux8pKj
ZGULZRp8XWO46SRBqQHxWJPIB1xWIwza2zibJ4YClynJ1qg7CBfEX9q0SNEgS6s1
E3Eyzylrk4fihHTrYLRUtShV+xFzwn3PkYryu0TNX4MaOtsCg7KLBQ66p0FrxMbM
ZjEtHo1a7A12A2XNsxH+NpZYmTb5Fd7J/INzm6kdFfIblquNjD3vlZxO3GPM3iMW
ZQQYl/LYfxgIaN9wiX05DlOcmWGOWybIwKwV43Demz97z9XJqI3ZJfhnrxzNwSZ9
W5k0yRxywhPzC+cwvvpEuE61RjSX6hj1Snt/Aq5GuYW7vNGmiGtuxeqDcvMpWuuR
8c2Dn2bjp3OSYjlajUs/Srt5+0Ht7F5IVy4DbCDPv6m3TPrQZS6zpgjJwPU7EkLk
+jccmT7D7GIm9dy+agmZb8pDgQXmApplL+arED7BN7+DFHcgexzeQ3ToSBfUrnUj
BsTengrRCIHz7gm7bRiFQR5vN1nVQ9imnGvCWfTQ1qzJpLzXWuAXSPbcvcE0gT83
XMAOOUicOIXOkDuXM+y8Ah6xlR5gbVIZlZNI6rJ9YANx/MzfvwJ0cWKEMEI89hrr
rbYmgG+wiv14d7Zk1cWBJCWYGyp2gDTrHx5xnUM2SLQMLiyE2hj4TmMShA1V3KQo
2o3IS8si0dubQyOXiLMqZjM+6Sa/yw1TK2nA4vBB/aTOrxY5YQoaLKmLK1N6Jpft
hZNK7uWLBXn2FLoqMO+lqnHfRR1xe+LL0VWLwTVVPMmz7VjaBP2QrZZS4TF5fnwO
55rvYPnva+3lV/3Fz+fwvSwvSd5L5iskPGR3OxbJyZRCuXoaOM28FnpQzRbkByVx
zDN3t6csgxDrrRaBKV/p82HFu/lc95EOjev8DU4VmfoUFmMpMBctcSfrbwxv97ft
KGtTQ00D1ok46SzC3i3wxlz3IrWPwwcGiOGZQ6FUQiUbWy/3WNzVWHBRII0DVSgw
vtrWkRvUrVOjZI66wi1yHuSN1HbIYupBzH7/NaJNl9I48iueVqZsce9sjWs8+nVe
wdqJl1wuiT0Vmmigj829FqF3ic/I8B/aTZYkXAmMAVPR7Jgv35Bpoo4xmaVxhhyW
q2KpFj9hXh1TBnFRap3SZutaBzg8JbPHqjRY5SHH5EIXR0p5ZBVsNqM2LNh61uSB
CJC2hf582z11hNF+K3FjEpl5OsXfYzv/OtVulqqWtK9VDwXlLU4AoNjQBGZFqv0+
YoQD4o6mBRYWepa3oeo0Qbm0Eux+Vt6wyetz+KUrMqRv/ghq9YZP468Qad3sugYz
yAjKQs54eLINojvu85XHbFXAKlENiHWMVcjHHTW1VW84bSGCQjVaIMchS0ghTUFW
PlnAQw859jiUO1sUHzpBpvOHB44St/Qz5qOlpWUCNxDodsnVofjl5ZpJc917dVSO
7Pn9DhWtTr/gcij9e1ka3OJYkrvVkWYJOxKUTofEhNK8NaTmYqSDL2ru9B4W2JNR
kOevn940tSxnmdU4l3hnxTejs31/SqpvArU35DFKN3saZa3coo4uCMD4yVq395Kn
1yleZfIhUmA1rb9yrIb9D0/9M9OnCiM221xATaQjkjC3DHpohK9k9A1ECWw1Y+tL
lEppUy3VbAoeOUgx26RqWO1hXpYcVvnYuKnCRvey8AodKctnt+x+AqJwDfL8xfqO
rMIiJU2bOomVhzErRLhb+OcpvRt+pnx9j1Fr1xvuWLwPYZkV9hJ97vhYun4dh9V3
0TxVKZJXOpV8BhWf9dhyQTlj1jqX+2LfoTpQIL6O8SeoXnq6Of5EdtBdLIWnFkJE
fPBidTodUfMBL9b1/HHgRXPLjQfkiOyyGBEe3lHLgP27eZT5EpKztgbeAqsr4cBE
4CDIuuP1PsRnf1H7GVXvxS6eI0RbDxLbT/iVlFIsTMRR6SQNLGsOwR7e5eVkO4B4
0wNjLtwZuQTPEga9TeWwZGoQEnvIXYyT07NIt2DeabvdVxqlI+THPC5T+xaBDzCk
s101GDr6KmqeUulX8IqDVXq/IAlqsINYjBSa3Hz9gcmr3ZelRpqKlOgElJy2j8Gv
JJQz+pCfF4H/25uYNINLbmscN7aaALBicQQKHGVHAcITPe6NJfJJrQH3GAnFKzbB
cYgYcfONC/10o99giZ00xp57pzJ5F/mi2Ys3SE9B5U6fkT72GyYkT12JXyzXJh+g
QExcKWp49UpTNND2wABoxW5R3t2rz2xJ/6F8kyvGcfMY2230fc5D7CPhiOUM4Ric
9uX3a1mx9xcW0msr8NdEetcDRfFaZt2zZFq4rnLJkMVYJaBnfuexQqSCMk0PEM3q
uS6P5sKuJICZBTxyPb03ff8ZiMtYsi/Xys1RnupJ1qPTGOHq88d4XXXQhtQB/Ha8
cDlDM7S+5W4sgTbBlz8FZ5jRkulPqMdbqu7zpsrPo54OBHfrYN6HWWV/a8dHmFud
BrYdXGwAJ5Grvi71u0cQX9HFMPs+FsNpRFh71H/Ymn9J78+T0pCiUuDO9UJJ5V/Y
/SRLjUb3E7hMIm9ckDQSATHdIvtj1iaGTEhAeRsljdPYBqNjX5rZqSx/QvsjIJy4
rhI6N0TDfTiyuf14EnOM64tuySmPZKOur7+x+/fmFlVq2jNLnN/+0/t9qvpJVEpo
NS1OwMH3e8R0Kr8bD0t436djKYVnFv1fZiUeluYDAFoWWJ/gc2/MARteuSPkqAgK
iqT4Tavub+Wta7zHGT2HSpdbH1Gkj5lgxsdfPGP4btpaDBdgYAqgm9t6TVHdHe1e
lCySAdPFA77INZWmBeGjlnc3WEyoz8JVq5QeqXSCqkIB4Ftia+0xIalnXfEAevA/
HbswaXYpe2r1a39Cq73I0Y8ZAwWKiZhdX+7lqI/iNLrzaPbopNo1PckNg7DXEvfT
3LwzyrD6E1Eyq+0h1BXfR7+LdjyAX1YdQeNsm0oLSKyhxcl4Ih2NRXVD9pbzoxq/
3yMfpZAKnU4CXF3rSOQylOjEjB6O4JU0+jvRdrz00jPOiv81sfNk89kB4EHxQyg7
3doiAAfyRHp9S03WxsvFoqH1tgMhrRrfwg2+IhyJYcR+LU94+wJbkcWL6XJsXvSK
2Yb80vSON5xzJ0K25s3TCqjraU4cBFxhAC32+4vP9UumOkC3nRf1W87EOejxqf+t
OhI+Iceq5Q6ztuJ04METTmhRiWYvVsFYGk6XXnB6nmSpwF6sRAFU3ip15xLeKhwD
DASFoOvfwD48GrGIoqKaMf9egpoBTZL5Mm4kjryeJNQRlCN2CI6vlaF44MbrEGw3
4JvfYjcXwicvI0iI3CJJAmRVsFcBzStM0koPlkb3BhYnjZC5ntkzDWglZOC7XbDH
yLs/JvLyHo2etr6XU96UZV9aI/orxDGht8SLrQzlMkpqJb9fZ9QTWdBI39Zma87j
a0kwuSk+zd+8VXc9ftaoFFR8vAHbROqDbXZ+at23gupAzoNOoJrIGE52oH6UoZkz
K/alqvASAOByHfRrtb++T9TjWLlPBxbciLKmSnCqTstVv5sJ0j/av4NWUj0K9QdG
Ne2S9m5z+CCo68Cj6YrnstKzYSNxoUFAil918sHBGkAPPD288U9wVGBkmO1WdtQH
G4UR1RPNkObAg1e281irbkdknxt4trWWPGchK3P17sfHuzmq+gdwpiHreyVAmSIM
/lV0ClDZtuZJPcsGmzMZrZWpjdKNWcIfdp/CFblTrRHFV0g7cLOFFuAX4Xun0EWF
Ar2Xf+fMZ+Da4NWa70UP8n5Xljr9w8lh1XjXUOdSPuQUSUXBfsTle1hzmmFmGFkS
m1y3Nx9aphrHuroLHLXgWnKipx9GInKcS8dGdxGxswUzXve6FQX3FjSzKcjqpqub
qOov3JjqGsZChoHWilkjVtjZaFH90slfp0YA9q9q/89TvKByG7JEWuoZf0bcQZBv
LPaQrzTwbEAiAEhW76x2iveMSHc1B9C3H/ad5JaZKuChD4AIo4DoZQJ4F4lOwlD2
87Ym0ovYcfrX0wm33eVR1Jt3YwWTGKFc/hwTo94OFr6/5YQaTLMD0qUQCviulBuB
r8XZomfsFFU13qejQi+TGNsjsvOZpGkCXHukl4WbzTPUzzz+qCgIiW+ffpCkKS3F
V8ESOUaWhc6NrjbJCMQTl1H0xrzgLZ9N8Z8GiaZhiwnus2RdcPZLWWvi60426g5W
THw1/nSs22JhgDayFDfjwqkFKT4UI/IuS5/2X8Q8Na7NDjV7Sy1aa8MvkHCxEhol
9wHiD3zXVV3yjYBLcffBDD/m/ipavJ645vErrwt26tpCxozAwBM7zXYPDN946fCF
kYfgXjtsTackBYeVJbMmavPYOdQ/Ccvkyik5wJU5g1AQ1XhKy/LdPu8YFb++Ar99
hroygeGRcCcfm7tV21R8YtJr7cGIKUUxIoqMHuNYyKgHDAhF1CrONjJqu22rLS3n
pjJnyRCYVAkWfW59S5Lyl5CXaYIoEQh70YjAKdLd6uWpFaN6uUnasZUIV/U07WOI
IGzgtcJ0E0pKlVtSzKsVltFfFuWKwsmPkbTqza7mcMsVMV8o4iPAtvIa9iPUJB6j
EAaiMsm8ei8v0sLEXFf7N0O0yKs6MIqhjHuaPNWG8MayvtJa9olAUJnUAmhiqrYJ
wpIzi/cMZz9j3Pxz7ZFnl1efB7Pm/eIt1Zi8BjJp0YiQnXx3f65y1fZ9vK19Qgv4
j+0neCGrMvAo+yzMWzWXaMnxX7MW9z3XrfMNZ9N3WDHOGxJ29PaE0ZTcu8lSLTqp
z9e/ir3kFiC1mJfxQR3UVMSzf5xhMrXAvN5hQPDHcXQSHRciRvuAdzLgNcv7JKlt
vAqrZzC5BXVek+nfz+md92Tz0Ah4+CEh/ikiVYLgyw3sbjbljqoL8naw/5R1Strn
jm7NQ7VsP7hLLRTFaeAcySEPcg7j9G3mMlEevqzvwcVIqyOdAX89dAf/LjiEG4M7
DN16b2rOd1T5aCx7ERWpbHr4cZHwXETAf/LuRvmiFvrDoxWSyik+hXmhp1ql65Kj
kAeu5DuTkG45UzInqQaXgWYKsW3ytqk9DhFB6XkI6z547F+XSVbwmL4U2a/bcrq6
+c5NCcHtPrp4O6E8pzFzuo2f38ohy/nUvhiPhcCc4dPw0z4hi6AmW7a9bQ3WAND9
vGnDBuIBkOhnc0Ybbvzv88OcnxuvPfLYTT1BDM4LmQH+PhnMA5EcN5+f75ZDMagW
i9jVVhJKeV5ceQCpnScact3QqToCoxyDRR+0YKjdc5zRoQw1/GgEkmChea6z1iVu
xAYU51soo50eO3nYwm6ultnkQvCrWkGjkVpFMyXxLMtilNLqs68TZVreQrYJn6s1
3Qur+lKzc9Jnj47Baf2irfo1A8BEx4YiwJoiiPNX5g1laAghq+DeKnp+lgQ9yO7D
pexm2haenFycwOYx84ChyA6ugyCiJAaqLtbD8sF7bOuZiuP0ere9iZzl4pFBoVe6
K02mPuPqHS+d9cHKzwNJnD5cReMrT9TOGygPVNrAZ92R/MabKfp0woBEWzhEScg7
gOT8qd5V2zU8icwHBYfupi2qWWEHO86gUCYiT/4virTT8Vh6D89BzD+8qlyrHJNI
ir71EdqHZ73M1HA0EMGNlBYvC9Q/8Q+pbClsN2FPdOdXAGYXBMkrJ/E1orobPbY2
2E+2ZGUHd26QDngdCuX8hEun3Yd0D6bre4GPKGcVF9PzFgOuiGGgBX5m6zCMQbVR
nrxcl9+WW6ZnV8EU8jpRpksLqNVEqPDGx0n7H+0BQ05myqL9L4SEtFGhHRfwW0Rp
cRBOzV9beCr480xJtsxUMr8TK+CnZiYVXtgFbKknFu+dgantr4WojWP6Z3UtRaR5
NSdZBC3KYt9VXEpBljPQ9vLNUYx1RnrqUMoHmUAjJy613MvRL1wrr6EXV7L3KI7L
rPPrET6JY09AgPrwve4VpnPvSzUIEwXLk5BpNuwLv3aLbFiGfMouSnG/HZ0fdsUl
MlvSydBkYwceXSHE3UvDQSD3MRzOt36gWX0ibixvFsMtsRo7fBQ77so7QpYiobI0
1kp2vc9Abt/1J4y+6IltU1bLz+UGc9mTsuxNbyyvkw0YnGypT6h/3lPzw0txrOAl
u1hqgDOPi2S3zuOTgjlu5PGDpZzY+BVfvX4SGhoVX9H0VP5tEQ4SepQz9GOz1Bis
5Qt4DwL/q/rFxle81hMtYOgcibOMv0VR2q/FXgqLkg2K8r6M/KKfeNgRd/2qgeCv
rHtNULDcGHS26zrkck1HHZ5FhrL6LHyAHip+/8gAEK90XR5+2VbSRpw90lcWRhQb
htAZSH6Whz4hVDhmy/jrROde0KH9Xqj11jFRo74psHpLf91ZOvK41EAvRO/EphFJ
P0cKUINC3e8gMZIDm54PXe3zpM83RdNaGN79759C/0tK6QpVmUU9LtECrHlcu/zd
jrd2CpcZ0mW9EDCN3DXsoC7U4iH3bWHBSmCZ/Y0c8yEzntTyeYqAk7IdnSbZ2qt2
ysTbECv5g6ELIJdD++cmU8FxLs8hCcGb4h8vSawRJXcq2RAaiX7L9z8xtOK2Jp27
yFXFk0XeuUkbTQnyav1FcJYrWRzGMct2Ar2kAuqAotc1PczE0UEbZqG4sat+tXsi
UYppp9LMd+dTdnBbFxLVcSlPF8UzecvTjrxcDoCjKRoFL9ZDvexH5R0AYV6o1jWe
0huhiqAa96W7aZeUW4LZ0/7EZ8xrMnWn0rwBcDXnytKzS0geaBxHWDONgKRJcEUo
uVz/Sk9S3dMKXJQDbG6NK3g7R3IePt8V7O/gES1TMuDccNS1Fx4PygqHm5jKnmys
D1vwfEDYFiht16Dw7dMlu6RC0Y/oBgEDvWvpXo42nXbNYMg30OQ44rp/h77kEQk3
iOvmj7bwAX/BO1cpa3Y7BoujOZXCwEzPq4TxSnm7hjK+xR4v7AmdOwzDdQBcugOv
1ODqU4aGM1GD6SWt6TjYThdcepFTRP5Sl/a7RmRpkFZm3gDlz7wQ7ed2LLUyyO41
dqKqH35pZpVk2oQUhFI1YzXGBT+6/pEGwnN0LM05DZkT2Ettro3ytpTfCVwy6H+M
PslJ0qwKuW6lME2gM1QHdU7wt1g4wnH33u8F0kyZgd8wLOcQYJVKJpAvMa3Ev6wB
053XM3fE8IDaWGoSD2QAiFdDtDj6Y5CswI3eDs8kTrXlAsldDJfKliQUR/yS7vmX
jmydT5nJRvl6X2OvO08RMXU1auXRBubHTPdgxJRZPXYmoUd+xv/LJH0yDt0/11EN
/NpeWdQnUWsOyR+K13YE9jtCPrKSN+gvYG/15HOU2y24YkF5eUEfli3Yiwxpo9tA
iMR59FeWAFZy4p/PBD/neQrs4v5EnduoVShXxolrQaN+Ug33xWageR08LHdicjlJ
KC4gkvXQx6XQ1rX2ffrXCwqM52Q9iVJa2zk0guHaNeRSbynTsHgcCv2iQRQq5H8u
Y1cJ/bQ8rpu3AkNUMPZI58EcWDQ8GW7I/biF7DE4BosqtN0jQW1dgFukoNgdXXbr
HF0/fbTeoZSKnWQB6jbxkdP6Y4MG3Cttzqt7lvsqXJehaXoj2clXeyDJJQmbdAWM
MJGhSi+feM/F5ueEqlGVkzctPHD0Ap9aLRoMWSTzuPu+LrgyBjfBQJHtBFI3ycGt
vqZPxJvPmGVhvEx5wBLLHriQdvzLX19NOpnNMXOVDkTezDxzjohaukPifa5B58G6
jeDAJgAZBzlSLaMYQAksSCixsPHAfHQQI4uzfGB4XmuaP1NhegyTC3KgrEXj2nXP
u24OqhRcaTERBL5WtS4yeD5CxEdGVnEofrjwndcs64Sg3clrm17Y4GtehYKgiFDv
7jzrtrPQq+3gUC6Uo+Zbk1YGXDonlUz7iRbF5USNEq37tpiIW/O+8Vo3Q7W7zoQv
+IFTsxCriBwsN0BMGC2j3haQwePbJl6PHTwPh7Ro/65ks7+cCRJ3RLs/RVzbWSWD
8q/GSIv7wbz9+rWPIz/CrxwoEC5lnzOHhWuyZVTfxDjFR1YYh0KV9WuBt7q0K6yk
2lZVuFs4aTQhW6+LALBnP7+RYhGt2wzasSNTHbJNw+tPMoQI3QOzDo/kgWRmsDMg
kRDtUiNvKrkXH8vgyPeXnNViJI242tDYWwPMpb6RCNCUUBFATG4wORVD0cp5i3yb
hLjdDh0AhqfoasUsJ9PUJfeHgsNrAn031XKu+Fo9K59PGrmHeNsdJnvaV6Vz73jB
XzPSQBql44iRu0G1JibaiEz5y26lzktSrddvhKdDxQI+7MBn6Ll4se9QTBLDL9Cs
eofVvVQ8CWmfZDhUhOaARMdcoP2KPS0eIUI6NQqtobOfd4y1cQ0UQzGJvfj3JedR
DFbWyXCKIP8sCs+JKTb2cHv5XWyPxtYFwmFEz460QwTIJK6KmQ4F/WPl5fXWpxnL
gc27HnuYafmKzl7VI1cuivV8eILVdxYMYulEmafJxE0J+scLawpnbytYHbKhXeLV
1ftHc87fbvMbKY2c6Dw0KPuSVed/s+ftpgt86lC9mkKfgY6fYWRxS7T+IR5S5yag
PRU0UIPCSpYFhDbXIkLK4ZLcB3Tmp9efVSBQuAg2sJ8R1/IBctyMH01WJAOrSIAk
4tr9onhcGZiFZux2a43otpZYo+JVuJ/8wrHkBz3Hk+fJjcTmed7iB+2LeFwCKPHp
xROCGFM2F1nSQd43FZ9lL6UGBoNs7RHwJTTviWjrGtO3NHQuiT5HKJkbd/dhHNOU
a3TV6a0PNXK3srxi5VC5TUJd6gzAHQnyssIZm8JRo9I90DvmUo0hfN2CbNGpZtra
D6aE2TIgh7qaWuoaRElpDyN9ZLdBx16QWGwDnrJWgoZ2JMYDCEln+MqVaPQbKGat
veuVATWHW683wtoc7C70vdYCpfM0WnKLcIAHw5IGYesIBy00gPurSAO+bK4zLwpl
bzplsGMnc630WzTmx1cn9xiDCR2cwji2+vGPOyWf4KmG+mn6p5NfGLzjsP5RF3au
+cgfX+oMAUdvVDdE1HCyHt5f5IWQvVySc7B3Q1fYURwQPacsRRStpr2BNCOVbiE0
CKnFtvz5fjv/4a4TVVCMUKWWIYnY2z7/PIfsFdaXcwKIW1M1C4zaPbpxP1FsXj2h
DqA9Z1lBhmoBHrV6goEP6vKHRscsvRBJ8nNnE0bFcbHnIGGBKGJQ0ILj7VsKhtPq
lY52V0fUR5moQ0W6a9jYF32DsEGIs4H0tt8FVdpIfuOenLf9+SnVTftKRDVQCYR7
/YbOb89ggHK3mfiX7EmwTQnRf2SgjFKVV9H5q7uS95D2GDcRAFvhZYT/9MaZVhIK
ZKp0jBWxflctY7sBJFj5oo04T5bKg29Bs7TwBlcd54wtUsaEy538BsdMk1cg8/4b
ijU2tggFrgzKnNjqnxsPSCCYgoJk/zKrNQplSR4v3dhdpKlH5DmxnkE65VTMQYJ0
SSJUqLmMcFf2dyN6+V5+7zsYwaKMpHWRM3nwUbsVSk+VDao/GPJ9owozzqEdRqCT
QV704NWu9RB4r5QUe5xgWouOopUoy3tFef6D9bhom59K7Xi7PdLXFtT2Ot4AjnIB
Q7wRYRpOq25ud2KUPLA2Dk8DzIt/DiEKZt45EyRxcMjQiw0pZiInLDr8da3bXvon
z+6n9RJHWPGZOcmrGgAeXXwQGJkYW+zZKvSlcwfF3AH9vEq/w2GNTU9Y+h65nXfK
J+HIybGGQ/v0O47rzZL5WSg8pI1CKrjyggXiP775X+zmW58YPN0AVDOfMmA2OH6c
u4dfqZLjNNZS5sKELQcKMVRaOvPyWXeCmYZxlxE1vPd2dIOEHsuOrpr0+sRyj7De
zSFh8TsAacWYNg/oIc7dtC7fqx9yXLqzBlhNmyb59LdcFzpsCATretnGfk/it0Sm
T2APymITc6iyKdcnNeOO3ITdyYeAR74G3nt73E8DAcJUD1mtLHboa+AnkHlul/6q
89gg/MdIxMcoYYZ3DaRDhfdJsY2423/UvHdwMLFXfCswFHHn0CLh4OVM+RNgbfRc
Q07RdLNSFJxQaP4qFN1wFwRktM3bpEEEUha4/75PuUDJdvy0cV4WSUmi6MduvcfN
zwqUYda1DQYQegX0G4/kKWglbAPuOyMLpzd25f5W3m6U4PGWClL0C+zWApIRWfO3
yWUr/FfYB7qKRAUKt8cRjbRqNaa5BdE73kHX26rZbGZUodYRllLf62aEwhcAVDy4
ZCbbvkE1Z/key/pg7qrQo7iFhp3YAv3oCSx0EOjyOv0Zm/zsnCfFm9cCQ9sCD+Ow
54Vq1jNxr8GQx5unRUjBK7A/Awwj/NBdf4RS6FJuvjHStMY3uh62vXELl0FGZ3/6
SrkgggbkCONTpqLoNsxnTw+iX8rBxPNOi47AnicAnEhE2tFsppwSAbOsJ/5NDus/
hfTLH/AEe0c/5zL0cupR+B/hC+gvv38xvS2B3Wc44gd5bm1lXjaQHV+m3z9VQg7I
px9QnuCcdFPDhAek2JT7XWl5idDKoHBCc7b1SsvWPdX1J/pbVa5tMfQaL9M9rAWX
c26vYcp+flUnsKDGKjZL72l85uAKbEbAsWvOUfyDr+W9EYjRFnPSGcOIf2+rwZdb
NDuIb7bIx840sqIEZk+eh8Ue92cLouvpoEzKHyepqsXORyhOShd3Ff5ZoDIaj0nE
aaVrnSjCEfKiWSnBRT5knNHzHiOyHQm3L5mpJWqF0o/9TvDKAtBswH5uDvl9tXRa
aoGaBf+XRiWzjj/RPSDqzYDXClhDzHmvXfRpsVtnl8PUwb1FJfX+WqVnt1u1Z1B9
ouTfo6e/04FI4WJ8499EEEsi1HqHLVBweGu8BGQ27RWO8yjnqWW+NwFvduaN/w2D
Ol893RVUKugRcHYcoFYspURW6gUvuwbH+GgX5DG2hY6bRe89mlNQe+o2fjzdUKMQ
3S9nKPCoGi2sWcTQlsTwGECZ1YUfpWCehsoMXnE8uetsVYlld5QsG3s/ri+TWsM1
ugnXzqfEjuSz+GK3SDs53Cqn4nOFxf32keq2p39AJqnK+Ozxnu0fy0W/x+z5hdeu
l/w/01rU1+RRTYYZeeVkHWu2HFi+bPIr7DxXJpzEAeYh2ae0nKE0XdyhBo/3EOss
Px3KmCXrMW7mRmLmuwQZCjbId1zeZl1tdHxQeysproysvTvV5042pu++tLusyMn1
3pFv1ewZWwG1QAJJ2TCQdJfNP9mPa/x7Y3eksGKe6M2ZmSLnEbYpiRCD6nEamly7
/c6QaXpYoMpYVdnJENydO5vGhWVI4P5aX/YB0iM2Q2YIveQo0BFn/fnBHCyfqeXc
WbDjPJjlqZFzbLPjglMjEBbQE9Q4HOnpefgL90Uz32uUsswU89kMBnAQJ5PRRqTR
VfYy2egnsQsJapFqk1x3N5L9uqE951FPaum8B+61Aa9/wXaaxl/Ioqme+pfERrxC
EOzEBtgjN1p1YTV838LLUd8WaNTrJow3VtHOuvrFtcjmWyPtV/wMHSX9YQQAoyXE
SabLNegTgqPme9ry78RwFZKY1v+PQxgDDpcE1xGJ7KBBCX1YvA48JrlII4GVIy0J
fyfX+ZTrACHuT5tp8sL9Imy5wThTnJ4i/JFqxEnQDkYcAvuwnyWqE7uRMfmuhfhH
ShRDt14bwhRXBp2I5fQvkbWzegtEpt01Owj3QnlGU57+coPRPN1Wf25UAnEcAb4m
BHNuDfbKKqwFms28sGKGlIqdj174QbXkBAxgEvJSZbo9+MEyOOwYidcCRPq+NeEI
9pO3LjZZvO1EBPlpOtxDndbtaTdoOO2RThiLHvn4gpgwFZ1LGgoJEN3t42r1pMaF
HkHYzCWQGUv35cP5wY71OxDyTGq2YcnutkTEzuOWwRmM/BZ7XcNkS9uGanxwUpOj
W4eiPPG0v+/qVG/dcDG/asP9kz2wpS2zRV7nD6fWZYwoadEkK0aSNQJMh1OQX6FU
bW3fg8rCXJxWpsAaCLRqbisvEGq0RMH7JlnxkbcTe32S1XoxBeSB42kc604RE6rI
Lu2qid2vD0BmS93UuvdOK1AOEejLvxlAm3pw8WFPERMsoOMTBCSbMPW0G8D3ynNs
+EypFG0ZnzqOKZ49ZitNyw2EMFrMscg4a5sJWIfT5bT8mG5EAcdI7IF2cHai606W
mryiYP/SfFx19sPuFz7urV+nP5VQwHEIgiBwfN5XaC76qghkeZmOQo6yJ6qZ2DX+
yHBLGdV8PAEGUQtF/IxyQljnulRaUHLKO5LL/cpaKrGar7gpVqjyUTxVOJoOSnXy
CAjjlG0oLkQ7YF/YkGzygGB7aEpmmDM+y4rAbcTircyCqrgLyaKGS2fGy1+swlt0
vx1KwJ4G/rAnTm4SUM6CvtVZWMQthV0EweC2Bo3X8SUMYltvR+7CQEygMrhogFCu
HjrdP3KijDlacTSrocrK0YHwS+Vs9b3rKZ/NfZoyJsvDurrTMyF6MoDoCaV5DaDl
mx4WmnaNVnwCx/cX4gVDrlPN1WWiuctx0IsFg8RGoq9wvrfzraZHukB0m6qOP3ZD
N8pRH7worYwAs4tFpxqLd253iuypyRCJhMCnJy1ilIbFq6mSFkJRkLHutoXmxuSN
atcjM9lZ51le9Q+AF5E5k+blMPhndHoH8/a6RaRvw+UZiMq+jCySoeYcLxJ7v5FQ
YYm77BdED4ECDJSi0uPUuyWESvPXkcJX5+mISKzBBYnoO51CB/3fqfNSC00ht7kX
7OQb/WE12lSNXeUVsN4s4IZFnkvhJQXO558YAasvLuX5TPhj82kakQBuyoXgL+5k
ydhdMKy67MoouC95F3GzAZJMiMG2A3Y1mHLcES0e3FXzIgc+34nvjuSYgm265I4g
6KFQM+NVVxF8biYKTo34WHIK6oBrSy8ASGGTUD7PJqjcjVrmhvlatrhY+kPPovIW
ZE4CnOE9jytCVpFyoQZPeuQS/webrtCCzKg8d2P9QtyDtwHEpdzy0/ZACKoRaG0p
MgzXYztZHKCen9XQQHP87WRs5Zn99B0D3pW+EgmlzRjAgFCRDv1jgMO0twC0Pm1I
5vx1e8MJyLppp2HUFfPVuzwm7Z9sGN3X3L8iED/pEQk1Tcy9CktfJcvjut0p5qNr
Fln7i0oz+Bl0/UIunsTV19UTv0bmazvy9JI/JWj6dYR/dM2EzEArQ3OE0VGyBBan
kMk2Zd2M5N1Pj/tjQHpoqKb9lCRLRbI3XYrx18j8xYwoyQxoXiPx6tMPSwb+Bw4m
rPLOUbBhpzXGhpRcu84EREnBH6MGbgkBCjKZ0rp0aX6zaWpr2B3/+sbiVzS5iTif
G/glkvxk9t8EFciZa82ROIfsTAXmGjwSQNY/1SzjZAyPKvOFVKdnTD35UIL8wwu5
e+Cea/0XIu8kxmYsAke+z9VZZbaxiM4ijKiAHrU1uuO2imG/KBPwI7pYW+bcozo1
HPTrARWZgfLE57tsKsRfbD3U+KmWsVRTH8L7keN9SzEBGwRtIBKaGPRJrmuTNmiv
NGrfCIEIyDcMt8qYzOC66LXdqqcRLWHEoRh1GLckGkCjphf3Pv90BHnLeXA0iOMb
hQXj+m9dj302V9R9HjF1JrScET2Xrvp/BUrztEvQzOSUG5pGmWmyd6zyZa4gbDOd
Rra4uC4+HJ2VWWIKRgDWJSx8s8I69c4P34RRAZsOY03rszQA4GhKwQMrEByWL4Do
Ca0toZncBcUTUG2C2x64F/NQcTjVvYtHF8dJwZ8EO5aI2aS+JsMGhnhLR5/W94jq
P99JCTSVVLOuqhuXgDpYB5JaGmaAy4r7H2bdvCT3wG4+PNWVVQK07bYAe6ybolJ2
H3ySXl1q+BTto6ac/iV6lSjs8u5ZxW58gv9mm8MKTnOsTN4ji1JG9ZNE7yi9W4/+
+iuQI+Ov+NN9HQDvPmAMj6Xs2hzQe6CqgktknktMZtd3SQtnOYD4X5tm8lfV0Pda
ddaEdC8A16P4ObWSqgAYTZY2flJ1KDjrqOS73bFOFi8PhY/RyRMEolJlCVFSG7Uz
vR/Px/IaECDiXvjBMLodalEbvpREdIJyeH14JbNKF0ExBaCSnqCUfW9nBNAwjyuM
Qv/uJn79cGi3Gt2l9HpKEOAbaQa2hcsuC/KeCjK+xkIlbndy05Kjy/qvJjbGZCTO
FOaXArx2VvxnxoGbN0A96/M7hriHUUKaz675BTQpp3d6NepdCjmlxNBlIcyhKNZr
EizqS8YNtLrrzkKfjrhxtgiReVS8myM5kAGG5w7INShyrfI96nxamuMRAtg15DPN
utXfzKZjldtPcNppyKeYG+uGPwAf8S8o9eq6/QJ5z+6Vl8jvN7zoai2/Jg3wrvZG
/AfVIr9FWWM4vODv3aWpPb6Ps4FIROfuEamUFbq68/mKT12B3J0CT2g2yH47gax+
h3GuerOwouW95qDkMOTdrLh5RGA1hAVd7HS76j2cJ8Ii6Rnxl/Dbhe0+QHfveVs6
ajXvaeqGbVRdT++Jw4OxZTlSxsrxWQtuuSDI9lxVq3IgaZfoKJPpp00NBBu/Aobl
9HA4Vw9gcTa47eXJ4uug7zAM1THFNiNXyw5JOWgO7Tad9AuuZ7nZICUw2M7EYTPA
Fe6uVJGW6VndO94b5YhKBIxDfaKTOBCXmetOToE/Mc4xKKsfTnYHcq5SUKAgrzMs
z+5YUkkcagu1nCqWWerOmn9DVyDHE1eD9T1hU5dCsw4I3DwQI8zA69L03Lr7H7rA
6fwBpBUtUOSg+qqs9dEjBDXd7XBL1V0U+XxPdmOdf2OQGr1+LqNMVvWgB5OVPz0w
5zkBF+625pV24S1w/TixktukRQFKxaEOatFTwUjS6Af0HXLp689iUqC3FBgZ9434
UF50+cUFB43Rk6Y5TnfxyxJtP0x4OmxSe6+vORuj+oTq7hVZeZ2j/7v7LlCm2f0t
zKNo0OiM4D0Qy4i6aOzENhXFH86kOYBhKqiXxhh3KBtF8KV74LwTdNRQoxlkXquv
+sS6vikjbsIZta0IraNoGOFPCCKYIQINKEWDP2hEv0a+yB+VFwGKaoyb9ksu2rxV
7S6DmUnteVg55KBsCfa3yfZv8O5QNQYmz3T3zvPxXbLWV/Nc1T/mkK7gSaUGX6bd
2qWreo7tv84fceff2eD/DCq/Bv0pO5L5i2pHiimi1lK54rGvRRjxEktLAK0qZHJ4
BD4NUhQXlVQLonVcKuJFMV1xebiwVjBloq7tjBof+2zbQzosqJ47oWA3XOE7L6g+
IEfD0rh8YmuzXBMyzMoktMBUxb1R3nBI4Mk3SXGfeuItE0jjY5J9yFpHrxG+m4gQ
prRCINJ9JQ3kq0zpxUqCZEDeFYXJhLkoF0hsiI7kowevzHm9ydKX3te3YkUO309k
cWkoOmJkiYf9XbyHX8zs1YQA+KcLjgjlQMF3qj2kB3EjtW5l2MkxYKaI+0ep3X7i
3e4wILv4+fQJ+km7oonL/Wi0T6biJaBHvNFj37PxNxN0v6HipSARweST0hp+7Mwn
vdQqmVLxzHhAPHCeGxy5nGmuLkH9typ4JM5k1QwClCn5CX1RsnTWiWSsMkyqNGO6
K0Ckzr9ixJz3FXHLO1cVCDCXuOAiGoZt0+4hXmSZQsjp+XIT6VctuZrQrq75Um7G
U99AsO+SVZ924LZSZxG2cRgRE6mN2LG0yUGviMhkDDtyaWUGBpUg9V4QjmqF1Xz0
D2CegaQIPgwfwjfScOs1KRlDOcp8ifDKhYWAbZN94IXvVZEHCD+V92u6LO4DrFuA
nqMSiuBOnPwVkbz95jUl6FdHNczeY9WfRp6bPHUWVqsNokTYFB8sGrXDXCSGxw2R
AHnngTMFhpfUb3gcjxvFDN2fnzpzMd3I3lShrYfhbDuPEql8sfF46+ggpy9t6X+G
Pv2qX5AeR524sgBr8gAzXaV/cJQGtLyLKYlUkrQvEVsm/a1dbwP/67U51m9/wM3s
wOKx9WHDQQXwJL1qCphWwuhvSUNmLwCCgY7VsRBvyXQ/eZ1bSkCdu9HvfWiv8OrI
y+fr9ER6UbabBq92zxeZLKknrIFyb2kn8gtLTkV3fksuTn9ZiTpD94TpfqnVYlDD
CQBKO5Jg3MfeuqUQxFweN9Wn4g8iE4d9pVkf9qyW3HMzEBxCYyL9EETVc/F8osxH
LC4np0gt5aWx7MVSPBA+5ekAucP92VaSiGppIif8YEWO9KoCgOB7wNMkZdy6N1Uc
+FagRJv2LK6G+HuW79HDy2k2UV6yn+2qIAESNNjY6RKpGWQKZsiHyOzcBk8I8y9b
byNDeRT7sztniHvuXOiVyC+d4yABRG4u4MHvMzT1WjRVjFJiDSqYQednverJgrap
CIdPkCpB0CB2Lt1SJY/xK/jOJQNbLfuDSXiMObgzpq4QiyJHrnYy+7LvlFGOum91
XEazktmhKMTobgVWlUOeh0ivmDb/PaB/AmWT346YoHBBOMhQ72fOPMBD+41Gee7L
x604aQQPgkPK2+J4S4a219wZVljKwT/EAfatCw9iwmjHPloI5jMuu8C1vjK0BVN6
Uc4WUBb4fJYueb4nllwcrd089G2PMPGYq8grNCH7YBcCTmqZYe+TY8FzTIAGZj3Q
UQBIsO26zVmAoUiHr/nc5EvkHvCTKNc1fkwschZKFK5X2ROmFHtdO7n7Lu2R7i+h
jHKEa/19NGRqySFGoMJRkcFlBj7QBG0URMnXQ1aPKae2t5X+Ar/aLZLC0B/Pgjka
Ug/T8RGm68cS89UPFEXJnuN9OGwOUbaNXkrIaeglHfiHV0dDQw963EJvRKntYaba
mQHkPo9Bof37rkOq///yUEhPTRimKhOdZhICaCup7W1VzMuztAF+pYcwBcbmxJqo
US1Ah3EU8wTMvA2VmA6rvSnuiO+ulPy0gWG0Fie1hSRHrE1igi5qyfifERbaTcfP
8jUa68IH/Q9WYf6E/7a/QcE/PYP7ftRsiUJt+sJxRtBIyaNGSSP602hlmyV0pA9E
leT3aTySR73edj3wHPON6U0NDDLJG7u+9tAJN+eyFz5KmPj04E+iNlpdAPRTY1G+
uqyu1yg3Z6P6wBrQ7zQAYhtCjhJ22PVfxFLPoLMS0vPYu2jOBY92JIWurpWPqx6G
nBvqCGYLnka1CB5BR2HTVo/1j70KICnIe6PAgGOteITqcFS0uNWP5GS7zMRImrXf
eu/bfzcaQ/ojilZP78ysbWI53j2LclwvMOpvizlkk1Edw8H/LHthlQy5WvIAqYl+
upHoD3ENAWeKlNsULfszPWie+0ETjGt9f9TYrV87Jb3CZ+1seoWeGauRO2vZcVJk
cGiPIuBx9GdDIG1kfWUlgqTpYYlsAxutBsFhawBln/8XbPRaCGquFDwVtJRSXoCE
gkr6SzrxoYBc1lpmTHnH5aF5CPyRKHGv8UudAtqP/UZEJzrgo1PLos4xw/GBmpKt
SYMMarHIW3R3KVhrZT4rbpU2hVp2SKXv4cgP/A2nNjxizSa0jFHzhPrYcfrgsdGb
gSczVesKkv76bXBbejsSViNqvfRNh+yhBYBRxkbzcxWcOzCKRfXB36IhoAJm++Mo
6N4+qXEpofodMoIrimX1WqrwlDYqrNMmiH08EHQCROOXw5ylDpSerM9Fho3zV7vM
bb/Q6ybObM0NwCxqtyssyfk6xjk0XPLO7BM5YDHIbF7kPhwYg1U6o5SMnXfQqcqe
+LfEYkKXv8XKs7GKgWuzLYtjueLBKQfYY6H1DRRCIYCcaYdnn3da6c2f0uFEtf4Q
amuL0x9VE0OLcli60bcrHdLYIifUAgep8bhc/pR0OVXhk/FDTgCrioaIGBKjb8Le
HgOCnECgPQX+Fhrc7Xo9pX3FMkr9IajC8ofXNKI8G9j4OZzaUNrItDKGBwKxaUSC
/7FKfHtx7KgA+HCTLuwvVWOGyFlQ/rsbfCocKBpusPHZzM+vAp4k5NaWdIKucZd+
+knzPZn8Qoz4gFIeAhNPLwIARu+Pi7+VACAgCP3MbX/u6qYgr6qlEbBSURLClbpL
t25S9BdlvBPTMmDagf+IB3kxEhMUVPfwEOKTr7mDMSHKOIJzhoQzfbKwmDiTYX0Q
zznx0nkjW6U1SARSqVWllyRmH/3tWG+dZyvIrwkmpIetSYy5hfFGUIEIJUCH5gJo
Wv0u1cz3KVf1NA2xWjog8vO9wpXZp7sEQ6a0pVRnI8ns3r7k2eAFzLz0E73NoFzJ
b7sxbm+5QeCaWjv8jBRY7lTyEZFiwGhBEG6nR5ejjK0IdmQcwnojrFqKc92lmEoJ
bDYr7dzqFBFKnwuY9/VDNm9d659Yvk+LMEjdwFVIQzxUkNzb82kiH71YMOvU3hVe
QYT/N5rQLAUgkVfoUcW4GzWLUwdFGbSFytMa6jsZoOLMk7Ppro+CTOQ3FK8Io18j
LjFqzJA06NtiUl62aQrWlNzmFmKdWa4FZW++F8kXH3zb0r4DW5QM2I+9i9uXOR+o
VNK8v/q96AraXcYjKy00/AZn1gUrb+DkkOJt/GEs/ExhQS5u5nC+MMxRfhCGOgqe
nbll9vDtkcLzyLMiWaMmP7z1hnTpob/+lxqerRgYRgNZQLzhcJ9Tk51Ld0CJvjco
G8DbmZ+Q0t9besOwd8eDH+QQeV2zUKtfZ/wGNE7rfVrElQlfrXrKAhTajAvsQsP0
i7UQivVyysnxAE/Lk7ZF/mD57YJS1rSoEyN8FpUcKkuI6dwAjKFtRZ/n4GKQ4N7c
adY5bBXnO63LXeXNpo1o6om+0edJtrE7bxjysPGpPvneRYU8mg7Kl/1v6HhmoVjq
UF7K7K2MnqmkbIsUH2bDR8QmrfevrsFXpzCMAkKlgmv40RMRMOke7DHaLStW6Hdn
Xm4r9rBDvHopmaCf9yb9lcU6WqdiunEbKU7L3UBsb7RpXp5p7X8H8dkAPXdKiws1
i9JzkYCL7ARKoOQnoGT4wxt0b83i+IhRS71DXXHdpmjY9oHDtEot4lxIFEMCr0e+
Iym4qBn2sGTK3lAVBiNDWWCMskjokJibX0ltltSA75tJtcuhCg/NC7eCAN3Ucff4
bSYxlr5LEKqb2VJzMGRo1qms3hzjcXuTdSl1plqlhhN6xhX1a4l5Ol9yTPHWdaLK
FTkklus6E7rkb9hxa6EK7/ygYRjUqNubNE2oNJGzWOivYSEOk/56ii2JpPefsjCl
BJcdp37hTTpScK4jS5lCSWFUwJPAnCtoIACvShP/nvxzsKIY8WwBqa43gOxt5P7W
d0OvJ+mybTmuAdBHiP7JDwUJuwKEAh4vsiKwsWeqEpgTd4hHXfRJdsgqgSSm32oH
j6K2Hm+kWjg0cjZ/OP7kYHP03OaVrTOCEiavwCBgF1TdlwZBYdSPUsr6AIGi/GRi
SlHp8PGy55xCC4TXS2nZiL86KzxEYphzKco6urzrvlh9l7disb/zizFchkLs9dR5
IbiH8mg4z9+HcypamoLpRV7JNjfcoR73Ea/XalaYCuCFCL8DD5U+upfkOhHfcbOP
2Vm92iBVjjJfukPWiCXbXCGOc4Ak2nz5PktJNDP2rnMIkxoG9nwVgivTxpFPbuRo
ZkBSiPTvypxnjmNRKyw2TEXQ/dJW3YOFToXXl6khkUWKhdEseOEJRg/xQ4b3vz+/
3r0EcnBQXC1P2g3cjgZLqdX9av/0tqKtVCzigYjtLTVYDA7Gq2ut1W5mLa1jgOSJ
+aH5sIdq5yOfyWIKQNm/GSwrnEmzfHrUbYOAR4/nnJ5z3D/9RV6ulOGcXziE3coZ
m1NeZlUBJ0TPP/kWgrQzaAwH9FqYSd0357U1UZoarj4OFhAK33FiCTV5hc6yBu0m
d376HNMQZX1tsZ/b0dmIcza6iXV3hWUgUsvH9lB51xLNOkRBaCe5pia+pN9zk+PP
aNH6fyX3l9e5imKCMFjMX96Co4zDZ7bSp1yBdK2Pckz8wtBAkaB0xlf116mz1d1E
VOa1p61uzg54Onn/HuF0tpw5DdqVKcwtGXbKqnhATSgyY7YDU217llt7EZ6vQxD6
9P7xnhanN1Wozit6c26L6EjVeAkAHP9tUZarB1tYEkD0NQv0gYHjmT8WTWhmuLTL
hiNNznDjJR4aDvlHeefKG3l3oueHMoTe9f4NNuK0hmHhwznK0d7uW32N0DdW2AUt
4pbNevHAvh+vkT1VAheRNZgW6EH9iR9vfyD9CzQtlWa4f6dTDJezUdzWbgtDqEx9
LBcz/lWAZqwOrs51rTRrtiSq8Xq27mhF4v1/KtjbzoP6gotedl1MIM10tOkhKWSi
Mf6gE3+HQgzE5hvKInHm9hWp2So56Oazsdwd29afp7Ua4zy61ybl0Nq5B2AptPV0
xCE3dk4gfXtW+tuJfd7XAXvLvTGZJH//CAPq43J26lqFXjQ03WimwvANYnoIi6ri
uF1ccHBR5+IaWCFGIw3YtQjALooV09WNtDoCBL/4AjgGAo6GwmAhlvm83RPt0NvK
q13KpnPNcV51ug43rt67RPtzOcfs0GPiL63RwG71OHV0jd7DNxoO4baidSJwROgv
T9L7Visr4zghd7rZ1fEF3WD/KTMQtIemfRvsAkeP6zmQSlqfSxlbgieV5a+k85s1
Af4qbeMCeDX4vDSLQ4y8kVLLqJSscKmmZvTtF5kZjbmAMiUCAbdCGd5CK+RsKZME
p9BxW48UufNlQZwNcjmkrKHCRpzB/Ch8W9fWPcVxFuCEDJG1EoqgQVucphHjiiWq
50ngRaFutYwq81jwu381LzJwImafJQ8Ua+HjaQ57wSQ1+h53PQPVoxVEwTcnVpD7
caVPjZTW7dGTF0VhyA7QWBkt7WzNaV86ZpsSAQTE/n3XDfB07y5aQ+1e0GyngcsZ
AYxfN95OJpVQ0CMuKojJtZDDHgY+5h9vPd7GhSRnxhEeQU8KqLv55ZlKg8qh2gGM
xtkICOYCtG7CwtCmzoT+UnQGHrbrIFSoy1Jx8haQN7de75M8umTPOnKjAcyTvSFH
mWdOu/mE8QA4OjK8hIGVKCr0O7qTfQkiI39WJC78J0q+4iFfCYaFHqtLP6jmIhFr
KdO170rRv3n4lq2YeeH7ExBvWp8/3Xf1eabDD0MvRZJw7vyih4rvtank9fNntkHF
MoZpP8cpCtQ90yhusBmLKxwWhqlOLMiCahDnFgGMBPFJZ9+g53GpVPaVK/Cu4hXC
iWRYYnvp9KEOgUJp8yFn22R5IsDGPvczZSqkfHwy8AbL+I+ser1LoT9jsid5j4Qw
pa9AhvC/G8iJg0hDYigw9eNakFbUtqKYgKhr0mHu3sSYwHxIM+hmNa1dHFvKOZvb
7hg+V+0vfP0vC8BAE8uClO5z3Rdfv1dILe4ztVJj/QD1aIfVsuB7BIFf2vtC4iGj
5H2BR/TlOhxSydYHfqTHsAedjw5/Jn0FTxKEAmNf8XJBiVaAOSlPIVpiC9yqbNQI
+MfjSpMOaETgXIbUxtBQCC914U2OSqr4VH2q+7h9SPGJx1SXseoELDrlorX2/M06
Tk6oTC9rWMdKinXe5e1vwuEfoGbhRThJSa4U9RnGcTzQ75YxZz0g6LC0295DWSq3
NdHkjtyf3w0VTbfX2G5c1AHN1YucEhs0J2ZsdzL5ZCXDE+nxhmh061pZHkp7hDhf
KqKm1bDkIkx1bvSdDzSqJHpsRhmkbHVi4bD17ew/8XIZ0lwXTv2YqKwizcJ9ydif
O8TnS4adjYFsGIY+KZ2jLiDA8j+d/YH68iK9fC98gMnBUIF4ucHHJ4mCYFL7CGX5
f8JeB+9ZzLEpHmtp+8oGzj65SzoA7wj3aR3w1Fi66B6nfVVFUMNrCPsToP6bwYCI
QST4wxDgAB8I3DTg4/qa2nyf0PZkqY+jTq2t+oNOGxygchtEBQzBePVYWhDc7ejn
BFeyWRRIShpVEeJOQ3NUP18ZfCzFjsTQh7bLw5z/0bYuK2s3fWkAxItE19WfBYUV
zhh1H351/upu/FmFljuhu89NktJ65KL2YyXG0u+9p3KHfak/tjfbM6/jsqOxc1OY
dwQfy7fISLvsjTAOgA+Vj+v6l9PJpt+ccYP//7lykY9wH58LiUUfsZxTHyF0ACAu
u8rr/LcJRA9AR3nSZlYzOO/WxsEG8gVrjdR6zEG40oppgCBhwF2vy6tGNkjE+cTQ
ARlxyNTETZq43G56kszSI0jU/bbxagePwV0GJPMCqL17alO1oY7el4slyeNjly7q
5JlNioBpGUCAeWtPxNdYh4NxQjig5UXrEFGcxzk+cS1KkEN+BZbsD4WVXqg6KCgh
oMKaAHVtbz8+hlSUNuBRX6UQbtbTF0GY8pB9+SnKNPjEkQ+m2gUNN+jfGJkz6/7L
tV1s844D2WCqQDjcB0U29d/te905aNHBE0hQ/QZGvLIRY1SDJTpd73XULJ8ms6Qs
ME9mA4YPBQO8eZWVrAa7wNZFwwUcseRtfSHq5WCJSc9CwbypXreLAV8ks7qqu1uD
36kxseXDLGqjFm0wh7G7uzjp1woFruuCQbRLqk1uiDo3IhJtlaAj1CEUJpqur6fg
ouBbTcvKlVAd3SV6BxR7ggWI/dsp/U+zsD0LxfAqfv4FcRlhYfMg2g70K4QPAJYc
Zs/l/8fv0F4eDFicnE5OyShyGltqwB/ALJocLNA8B1Ulsb6j+j5Mt47Wh3O6rtC2
ZJA4I9kdNCmy0o80yha1Mv65DTY8WdL0j9srJj0wfA/dHpJL0tHE3HFT1iq0LiX5
b+mxO2VReM/DsRtIM7XyL1gHMuMAgRulomHq5dw9baKhmkqCOaVbIY1OBVmTRIfO
P/wBhoaJ9vQeT5LCv+2Qx10PCVyNijRDk6v+Ao8KYnv9DPUIQ8tdBhxxo6d96iyD
iwuOx9qRwqJKAAe8ssLx7dLDLRJkJAinGgfG7BYg/tmezclgSW8nfcXI6Yp6YDsp
cEcv+SbpS/8vxn7/xMjstJoznUuDTk08BIXK3uTfzopfh/fMGaIJbZyVo8ET+h94
NcaAD1x4s9UW2ccJIzB94+mQ0y8tHMnYChQv8sc5Wk4hlUFLrh5cMuVR6vo/5XXq
u5xHQsjLGdZ+aZN2XxP+/beK0coR/oEusyZfpEMs/iAkFW5PeJ1XUuLmzKEe9Cc/
nKpjs92vRNpNXZp2hwaQkqsJZE9kUASOONWbdhenMzFGepnnEzenlAILYCh+R9kT
b90h5bCyTypl/haCmemu/qtmsjSUBY4mQGX++scGARnO1W0/XOYNO7lL/yrrHMCr
Nad6yftOGc6P90IWh5l5oR6oiUT4LzGr0cn1LM8csyJh9tkvh+FuFp1NUlHc4ssj
blmBNJP0G4nQpoG1msO/b0rNUkkvPiw79q2o86pyM1fTEMAaECExdrcICfFr7mfX
nroY0dTU5AXI0QSshH7Rbdqlit8f+mHkhtqhEQmAMQlVfHKzskwVx0yE766HhOrM
ZaJgEUuZc7WzRidFuYXBp+pZM4xMVQBbOU744POAA8GMaqH671P6sxkg5y1C5+/q
dW0izs/8pTSJ81Nyoepav3wTr5IrE6kWFwjurjyxiEULDj/iKoawSgnZrFjhiHlx
Kj7jUi5YRGQj7F6Jci4ANpfCoVExy5TDfl8LUp+sXi/dnsyZraOg1sBptakxiAp9
Tk2xCiN4SiYekbezSbHAi7DsFkFrV05ObaOMjMH+7a97aqhDqU6syfTC5lp4+AA3
jXCNkEZ2N9/8jaudJ2bFDp7jYLf5EPu3+gqCS21Pbid9sGNh2ohmmoM1XYBEnPPR
BP/5MMpPP5f6pIXAuZ8fW9g6h+XlD5NGGGAZeaH+8pVn04QbRhcwfMALirNjwnai
MX8fCNWkRmSooXwu+EOa4gMFc5qM7eps6cx62eYVMn+GoXL47YBYzYHJdsXfBZ4p
xooPOKLyhM+EkytlNlfT1pUzsiZWbfMBd3ELDPlElYoIEsBhl/3ja3G4tgeRYn3L
NgM7QQ1P7IvAr+kQChxibyQldVq3M0rVg5494Oj3qeogip800OtomfLyI/cHb+wa
Kg09Dh1/rp8z6ceicE6VELukx0a7YldA/40xe4U58iKbAMYziqSRMplYkLM7ZNwR
DI9sm7LyIKmzB++DobPQvz1/h3cC02Vcj7p4yusS0Tm1rJ1vmMU0NAc8/iqMIcUu
EZDDM+lRO22cE1np6GBXqZrGeexjbVXIHQfX/HL98JD48lWEkiLg4gWpxtT1h86l
rM25WL1YGGZcHDJUnlD7/P38oOke+BN/ZRrw8pbzmNCdu7DOtqvW3BTr8yebxscW
UASY0KpNl+y4KWGeISq1evb/Ut3y6H9xOuLzoqMoCFqYLVmMVLuYXQX+UjVEgtNL
s3dh+0EeoLcIRHstvgyEiQeHEVmkaTfMuAvrvg5a6BlT9DQJtAuW4+d07TEfDIIx
K3V/uRnDz+SJ93KxPDI++s/CSSriUYMaVNnhOjZ99ianwHQXWaRSRw7bG2tUypm5
K2ut4IESa3XIN+HLAnRu0SC65D3iI742lW6bRqFmgztKHeMI/W9xU5sEnHcgHjsM
Lp/CShc9b8rZjwFo+76qv7b3l3TCYbPqrl9XKo0gTQaSmAu9QpgrVJnwkANjTggd
B5AFsGQ+03X4iW7wf/yl3ItsLk7t0yY3TED/bdHKA8OobHhXCO29yP9HB1q2aeeI
RlkjH2qik7ZB3duL2+RBpAIIxcH8Up4TovbfsR3wq/eKl9If14HQqKQHo5Kah4m9
XkqPSH4t3G3aI8iwkHghHQdYDGSA0mMXcPIWb3rmEf6CFyEz5spjwICSU5NZzb4b
qCp5vcSFVa+WENdLJt1O+xX4ppdjsuSXnsZ/eBNCknAfKigcFK6fW51Uud3CP0ZP
yVGOWR/J7QWsfWYNfn/4b6DJld/8S7Pn3MyfjIe3SoP6TvRuXmg0+8qoeLQ+DxSf
KyhoRJBCTJZP34UoEnVZUsyAT9yM/KvMWpu3sUO8atHPvOjm7UZL6evHet2CLIGE
O9QfGUT9/vYLQAq8/itB3hc1/coeT15Qr9XpoSTVaAJnRZsso0K6nBDRQ3eisYuF
x9mrGE+w66uDtjMFeM/RCoT4ws5jCojRUN8p+utycMHetHAB80sqgVg/tkVY4iNr
Toa+hoEixZIZbIdHExP39N5S9uEaWDMX8JBjg9V5imcO3wc8Bq2P7RTqlNcnfA+K
6YfDEq+fmkIZcUSdB8RfSjnAARpjGa6M4WuA2QRdtnr0LKV+rARQM/yDbA/z9ZRw
QCA708rxii4dtKRkbmdaH0inNHpmk7yFoV6ComSoBdpd09wMQchteRs+o+RlN1PS
LdHv+iLhQf7SfB/W5v72El37aGTmmPG98MSu/s3Dn2jjdveatHKOURgqt95+MmNS
RolcXoO3iRXcxbKhtflun68PfKzWP2vySfBAuIP4rySik8s8opr+K/848hHHaHyy
Iz/L0VrRHgT/mVDaPrDUbOsSQHX2JnkJAQnZF13r7rJF4nGW4RKts9jTei4EPmHI
3c0gtQ7ASTT2Csf+C/NhgL4660IbPZd9/qyLenyg+gcaF/S64BQWcZJA9cyrhYli
hMvSm6aQydJeNNbbe6GcMig/ZSFAzN42ErXXIWFxztDvt8NBF8x5g2/raMdu70a/
G32ta6BeQ8p2eI0XA4cExxZ1+USxZgmKr+M3lnfIMWWW/AynZDwvFGAk0d/DeIHm
OjtwJK4bNp0wzCNMQOvLAViLzlCviL6dqdm9NqIesJFVsMiQw26P3ehhcd3ZFA9c
vBNGUejOcMRh2v67hq8/+FWH+9Xe9q9/hT/Ur+faKf8OwA8CAhL9dzC1QZmedXYU
/Hm+5g/GbppKZjLQO4c+gsdyrdU1gTgIvKXTYGUdMtNWbLRy3YbAgMeweD+iBa1m
LorP2wBOpcOpbKFfWfL/9ikMI3IpmxmQy2Hmzl/WKr89n5AJV50alqVrjMa5jMOI
1jtDpD824MsbjMaqCeG6QIle+2/VVdlt7fFb0RGihA0Q14Km7xf52yamHPoZ1Bu6
e8otiOVqE7XlBNTCg1svJ9EiVrpp9WyHruolpIAqOuZUZ8CXiup3lSwQaENgiIrT
KOpkSPWShB/Is5QSDGVV5lU8KYJ75fbLozIGDJWZQ3z7NIy5NF574+1MncQSnqfv
NOr+EU4+eRtq3QpZHkxNUlNQIfQdbmvI7RYjw9/Xr6Q070Xje6Fgz/ufvSgEZKBj
YjK5VtUeC6QXBnXTa9MmWb8H4jt8HM8JCT1OOVr7wX3Rw4u+O3kDh687FLNE6cgP
ddXjaYzVSFCulTUD4X3g/rUnW7TOdP1WM8gLdHl/xoI9JNU0nli6rqf6lTQ+4TPp
K0rNrqGV1c2qnGvASsol3JJ2PSNrrxELI2+DAEhY40GvjN5aGzVEqLqzMIMe1Ysq
Tg0aiTNAwf/R/MxtoZ15r1/fX763NCkSpNUlXsBEBz6f7E5FNZYNXYUc7WKBw+TL
G5BnnRqVfN59qrXsr8brL7JP0fqFKUqSkQAmyVxtG6QtDXbrAiRKhXba1ByRwTzL
DOqknNy+eaJV3GgPCajHSCTezTLBlt+Bpe4sdZ1o838Ak7m3MmrWtShndlaFFXv4
d7BhQrsec2jYHaudNFcV1cOQ29iG523dj+OkOrRR1OGtazG/lHRz31jm1Si8qI92
0HZLi6gXNnZzY66S8ykvCpswprEuotoQ4tQu2ft4D6coq164jiG9BJLLnvsvRcx0
aYYpFBlFKJw98sbbJmJAU35CTCvFlujddNXV1D8xsthIOXMS05HYFeVP5tNuw1w8
ehRTb6X9OQetlsgpNmOLb4WsvoCxxbnnfpBeI5Ws6yKWL0LW9obOs92S+uRruYER
HJUroRRVWUFXTnHbgxQLbVmz5glOAUUKVVTvsMfKkDuKcVn+fhvxxe3k4bkUPEDH
iQAvpEScDWca1A1Q/0TX8kpY5nkTKsjWsXyjJitzLXszqMplW3siydGGLiOVJG8P
A0nbY3FAWE3odwQSHD2RRMX9dVNSk/5exL0FxT/cEOM0vnliLlB91Fw83T9KwhWH
3BFD2zC+LXTWj+MQn2zeMWVPWb8gYcFeaEvI4IehS8uQ0xbpksdrUSQeX+NJi/u8
VJ7NjQjYb3lvRHpevNwGlgZpOdm6Ap48Hc/wjqzr3qmlhlQSV4oyRNFQBfWdxinv
VvhdBZBUyuO2MHh5y2i3U6xdBmkHJNOasEJuvl4rjTcIkZcZkDjfbXVZLWE155KY
q8WDHTLNZrdudkYo/VPZ8wQmmLgevxaGq9h4BpYif4G5OpR6nk8x5d1sSc47Z15/
q1uj00UX01IR+m4N8dB92VeJqa2rOeA/2OlMd6jMhVfvcXQ2ewiBH5gfxiCcZpoc
53yOoVTKIvOjosaJAIWZ3rUUaKkDmROBQGFCEWXsJblHgVeMHkiCB9PNeDfOXLPi
AaU8QEncuDzmLpO+3J0B0yIoUgfYkWzxBhNSbNRJiYUa909Uq+TwZwTiQSP4RWuz
DKoS6TFO2Z3CnAKi6+nL2M1+cUz+FFZjgBozzvAkEKnluAju8CUfPUxr1kp3tKbY
YWG+0dUMFss2XMlUuzbdLPNhVezyRQXy83CQOJKESziUEwWCD2+2ldXxgDRaN4No
+XmCzuw5fibQPmiwiI9hPFZRjNvfK0CpTn1pa8qOKZZT6thpajVapK/SKpZE6Yme
dZpXXbikbzjMCIPkHEbB+/lLDc15gEie8GsLLg1fW1BoBRgpofFL7fzGrNnsTy+5
iPcUqk1C7s8GGNLgQ/WGmr48a6R4MEh4+ilQj0craqdYZnfViMgAss/mWBBWtAOV
7XXz3UC5y8jSqxrD70zRkPFVepKP/LyLGnM2HIW80TaWTN/61uRqLDcHeEz0fNG5
p3JxlLiEBZcOdQ7iYQkgb4mrOn4lRzDYvWVnvwT/RG+mLmjlhH/gGfFJCNimKTki
Cw0q1cPivVMI9xBKvKrrVa0t7yGnP7gxOySaS/FuPsoplZGgPNA6Ttj1vYu81hSI
nfEMkaE/hO7YBEol3ay8JxCQMxAHp4mA+74xeXVV+YTtRCCNrc08nvEHa73RIPM4
H0j1YNTNYtHCkGJlWpMYS8nHtxKnMrUWpq2jC1BjK2k4aCld60nKBwugRaWxUGZ0
zGyuMV85MWCuvy+pJTCWhjh6I8vmHrmIaYyYZ8Sxs4MNTOMkRZG0b42GowNI/tzV
JAUA0VrkuAZbsFwh12xkcbuUU8xkVE42OSoAJyZjyDto9UgafDUf/izCoBRwFdeN
7NW4e1/CvZmvhQpzf01/Tp75szq4HWxp42/S8zOW/OAjjJomdJTNbPvzE8XA02d8
VvsCPVrHeECidjs7kqyQskJZ03HvQflnK/QR8rBJXe1xcXr0eRWcRKXdoISaJaxo
Po4KrzRFSt2OUcBoRg7LunvWMNVPdSVgivjWWkDD1BGvMRdVoSwRT7JzDQf/Vyjb
0PXnFDTT+jZh48V8nVfp2kZBGaalQQWIDLzV2eKYdHGtw1UlFSiPuj8gkTEm8c33
7pmeRVIpme2MEuD7XHsO9YTbYXoK9Xn7pF0EZqAyknblN1ez3d+CSgcoKyGrzkB7
dem/ol4LgjrOzFgnUeBf1dOsnjhXGOClJencG88dIivI674m92txUHAktM43qm8Y
UhNQAaI8ygk+wUfZnTea5cWsgkZ6QbGiVzcvOzhgSe7F5imti112avsXlcGKznq7
959sd5nfV7KtC+YmtAPmuhbtO4uBjXg0PSZcc8O12Ckbj7uBkJ8CMwsoFdaPwXcU
uQ3kr7gAN0HN5CpembMslq2YMfuw461wwxw8SllKbyuxVD5cL6cD6Z45zE2c4i2i
ESQYjDQnOimjVK9LDMpaFs/llxtLwF2LzlnUsHe5uL4MOp1G7sykSdhOJGbGYue+
Mt3v1bOVheLCg6NkzHQZx4fxuNLWJqPtOzc1cyzkpDCveV6lIt+eaePSDYm601fZ
K5J1eJFRJEWboWuF3Wd+XkvHWMgKIxNm8rruhZaU1wAmK4gRDG6j3pX2qa5lzveu
Ijuxxu/9n3gYGSONliy3qnSa+2qMGrCz8HB6dvslVVTMK0u5/7nzQGqCFKVIkiOg
8VQlq73vTmmjyOwDhBUrrw87TiIV+8m2D1XbNfH2Q8m4lU8s19Gk88V3pSjaQR5G
dERQwuusV3LWcgx0qV48GT90e5bVSwETDVmKWEUq4XTNm+IcKhmW9Ovzn7X3BGni
HxuK2rg0si82oJFal1MmSYZz46IC4ebYnqwi0qR/m3pNqLkbHUDfT6CTRU3Vv+rN
wV5agppDv+/YMfzNSIMmFizAkBEr6YP3wD6Qdj+PAa2UdsTlegdQ9xJEccGI1E/P
YNvcoHxe6oJawQKi4cmBwWR181v7pGdygAo8GE6jj6h/65nj4ka0BjY5EE0SGzn4
ZzmTAk5lU1jjf9ZVn4olHF+UPiK5A+1nb2Y1OoRZAPJZ5eHPXpYwehkWCmiuMfez
o+/vrHtRtVGCtvKEPHL3X8JQVwcR3iz6oyiRbyYAYIxAnuI7+DKaLW4R/D3sQFta
snU/5XUoElmBmrd4HRo9VA7Jz0wbG/kssB5uvKzTfe9doK2oN91bSBjvbXMU/zFM
yG6ql97CIRIILgMsz4k2/xxiIyab8HepRBgONt1XOTVV8oL+OGzGIfvFduiJumeK
XJNAF7n4ovLqamaNzI7l2VEkikirQCOi1UvrPAYbQozrBPcnrKm5+5GfvQMWt6Wy
iL7dxtlhDj3hyob0IMuhHDa/yW4j/rOiWnwvx12AIBHjjkRlZWMF/7C5gjthPHn1
xzq1DRCmIeGpKtgS/KVZ6zJZzE0RB17/B8shBTScaeDxoxuoB2/cpxWT1qd6L9xc
uzi3deV9GEyzFghgum/2Kjun8rX4a2ihdqEHSr7xXC7yO+uVkf1vydgpZPhpMkpA
QpLcMLiuxXgN+09uiew7liBJtlWEQZtfM3+JpXAzK9PrQgOf7tjhz3dCw+NjU3hY
aFSkTJKg9oD1XjbhdgHtjFdLTYguxlEPTfOqVCAPoRXnSCNdRgZYvvEe2zmjWUJp
V9C/lxzuACcKFqg2kC8p7xz7fT/YY/LLqheLy5vDyuRURN595vKE6c9/x4iDXfgN
FNzIuJ90ktWsbb+wiCqMHbky70bOSAEI1Bxa/OuknyC2zf6Eru7oNtTmcr+OiCnb
35Oq2EV6szobxhE+2wbsHPxzq+mGtF5DJR2r0NzTzK9Zav5sRKkku+eP/iTQpMff
OioiFhqd1tRNutPLzFELJt/OGoRuecTYshXGZ3tFcJqbWVSf5FYdeZpMsQqkNEYS
yegbX79BeHgtN+9Bb6KNPXT+MlPsAyNhK4UAPA9u/SQw39s2/K+dXSWJcIyVHlhR
wWuBwKzdhhFYqQoiS8XqKMXgzzQ0wRgsD00BjM1i2W3FhnTdIpUH0T2KGXYxGflx
juWsfp173fjIcRFhtQWo78fk/Sw9gGUi7NtoTPj5amMzG5T1AAjVKo7n6EtbmvYu
GLuRoi3QAtrqCSwXiR2pc7/XmioOS+fCm8JtvI4TqA2wRV3Sk6914wyDKbqOqkZK
+PflC2vRipj/C7RA2mviNE/fqXPIbrvBDJXYYLL3OeG/0ABeYobKQ+lzCrRGQuyj
7BboAZrg+9WJaiSrm8W+K41OqOEZBEQ5bKff3iIUmaivgNKixFFvMMxGljxfoCYK
MHs1iE0Ai3vlEdu929Z0tPbnP4dgCXFPKyt3IIQ1s/jwfdoAb2j9czs1N3yLBYGB
iiYyI111GavJ2sZefv6bzGvAtf03OrJ0T3ean/mXcR84OftIjvJnI7hrQAwa3IwK
6BUGNpK8DYfQy5KU8LjSpznf1T0tjgSoJSTJeNw8qTBxPv7cZNfmIZfU7+55cs9/
1AQ5jTo79SDttGLzM2HBSNlClcgWCFUJaJ2m0HCaoh/FXE6Hf6rblNWkg92pzXfO
xFisWQeaYjLYTnOEldpTW0qbpD4Xb7qxnsFkuThVpU7ZIhPkOI2XmNYbnn9nOqb8
K0nqgNHKMq7TKIGJrpHV8V+K6w7eUUGyEm3h5bQB9QLC5NF5qvxSN8vB3gZVUFjY
AKhpujtqHE+mpToqDEe/d4xbuyZDMDXJhWllQwPwkA3itVBBYbmyXEUsTfSZT/n5
WylhZmsrIdhHUVZnbmVrkGLcw8J0IZzW7Jp7maz2r2H3BB0YklccIXrp6rNWcAM7
dw8wuy5H6Ny6hrSmcnSFlyPjJNMfow2VdXpGCZy1I53vLV51td5MLO1fCZ/6BaUb
XiGFPJiQwRl9FYqoAsaP1wNdPoZeIin/NT5gSSdmQ4vmDZpn/NgvBOkVl03DnWU6
SglAB/um1kIPKEYS6cmv8mSAPyG+xmbuJzoS+MS4GV1lWfPgn6RlwWbhsl2G37qO
nzME5Ah9iXR1LsY9AME1b8O1izGTPb1HFKCVLBKMEuM0bzclRrAGmh3wYREhQX68
nNrtD1g+fIiTJEHXYuVTp7NlP/AmkeA/eFRBESyEWP6nVDKuZa1twri5+ZtG1uMM
BR09qV6FK3kGnUjr0UcNjnt7eSDwLEJVv/rX4qbjgpFCUG3LyHLHEt/PvtOPYu7b
uCP0ji+UJGkRLIZ31XA648wFR+HF2yEWTFE9BZQf0F4OoYxOhbSR2wUewEJfg6FH
GTaQRaa+/3unRbBq0fowE0I8XjCw4Kk0yofdyJr1YuO7TwIaed76+INnpPyu8MWM
X/sA/3djdNcYZ0BlkKqRhCkKU0ajxoHViMHP8gJrNzIQW+hldKSAiXnE/zXyq9zo
ju1BT4NXcnPpGwId1Nqe1DkI7odDozIoww5sdQP3yDaBo1jh8hlW4VD8m5K23X8e
kkkXEzqWF3au3wFHeF90YgFJm/Cqyvi/ez33fJs+mJf1MOuxk95nh5Hw1qp715sn
scRVQMiWTtuO3JXgLeeKZiOA0ELabOWBkMe59+2Za0PqdtBx/yhEOlPu7lBvKXml
Alm1EocY+4tfxLaI93rAccwPEI70VD20XQtFwReFH6yVAER+cucSkvLQ+lFENnC+
6ytVLjV9jmz5m16Kud+ynlfIbAxsmvmza/N2A8YBfOIiYMmfFI/y5PNJ8O2twf2f
hOPSvSv9MdnODUl9LuXI6meR84Yb+KkyA5mwpYCzW8I8Apvq7fMMwoqBV6QIUZaS
FWdhL/vRmBCvIubky08VOcg39mgrR1akk0dsDsF9bjw3pW0GRhzvgyGf+lv483x8
PiC20s0vOU5vVgDbqozJHavswz3/Fh0+31na7rKf60JW4U8i8M0yDhqXCEtjVjK5
865UPEnWaKhB+/V0hyCqr/bkv7WNZLascDSUsSATn23AJz/uurHNzX1IjCJj7mYZ
C5KJ1tcGVDNYdC/bkcCKrMlRhTX90Fr7P/qVbZTx2ferVlk3L53q3zOBV0u414f4
9dR9zwgmdDjT0OkqWDT4PwChOnPBlw1ygkV6DqkqoEqtucxp5JW/12zGfkye2g62
H0pe7Zk2eEWs765UxcA3b8RyycC5lqHwdcVNKJWAB6fEWiDRjYoQUXllN/jNONkD
5KRJnD7iMis3tXsazHwfNClaVPJGKzRkdDa7IhaZndFfmDAgImQEb23ybxe/pwTP
HiOMq10Xf7yLvY7zJPdXAhCsUC7hyN0qsaRM8lGMzj/IsRCfD+2zGm8ZYKKFOywa
pEOpSTYl6W17ehrp6xapr1Rf6RJWKjkqZzmDRB20qXuP6TrA/uHMKjAyA6aMcv+R
NneyBCwa2zuf0zKo77ElaZDGK+zIrfXxW9yXe2EX8RfF/ycaWYSati4Z4MSGPCkF
jC8X1SpCN1E49htT2aNpKUwgMzYMQ/mRS070A8wNGDChX2fih/EOTGmOF7LjmWHB
I5IsIc8Q63xBMg5cMlIRLzDcty9RsMhSg5F5EOXrNo4QnIqlEezQ76+qCTJ+MdjG
RsoL/b0m+IwIjB8Dg4srkaGXC8Xmn7EAZmiSbjBg5L2JBnqs2nMvzwF3v+JZT6zz
R1BD5F+Y2cHUFAzAPM0xj55iA5Pq7bUKpm8JXPrYAvm2UGRd7151kKj3k/St+3OY
x44NpW/XDsbIu2476WcHeHNkSPPG/weyiSiKLogz68R+CMqBz+hB+8ruWQ3buoje
NcIO+IKV8kEHORMft93Xi6jRUBkLqHnJ1iKU7Q9wQtTk41aXpWhsFoLs7ZpkggZP
MuyBP9C4uwvj31mIsCglYRHdbD5/RXkdJVns73lzol33guga414Yt/VG10OXgx91
BMQ/37PdKwsqGjeU1Eni2ewCJ4oktOM0ahz0Qmg4jsggIw1XRDkE++MaqM17HMGK
EHWbU6oPXPxKyUdC/UQU4FOK90kXCpKBsdD9B64EBHr5BLnpEwikLcp0PLNMW0ic
LXSICnq025CNVaGh6KCLjUbu6VEWIkObPVUA8UWAVVdfe/V8z6hDM2TxWoTREXH6
uy8nTvIZJWQb9S/t7TqKJpFtNRfzKlKWlo511KSqHFrNTQ9yogsMld2EEfiRUBU/
iGp9Jq1pWbhRYBkh6Zl+FBhMJrbXLK66zoHSP/BvhAJJb5eK/5qBBPxkGqsP0oNL
LbFYE3bba0n4kXlxKEtnooC3vDNfA9KkaNmHmFkUKn5qpASovp+7tMKcTBridM4N
k0YsACJ2pL5IHq80Rc3OusE/jxM5tJQR48d/IHCWWO6GYrsKRnvyNP4UG4e7ddIA
4QBF6NsNO7K++Z6uGEGu/NhIFONHnBCny1NQBA/T4kFzS2QN5xPRTnWc9lmUAjrO
5Je2dXjm6qsJN5gTB1fF4YUudWoe7Dd3j2unyNC7ZKm2bVJ+rUc01z1zi6Uxqv/G
QRWbJk4yhJEpBXrBRiKwJ8CQaQ7IUaJuAnsVhMATeI3PSn0NRfNe36ebfeyKWiqE
kNQ1LJo93shbHLyqNRecefA+0YCYNwqkf69CV0lEq1zPsfL7CwTfjnMgbBykX/z5
nZwPlSFj87/TlHnSEJuLIdADcjNp1hU1INJ1loiummJLFTwrl5ZmV0vBSbZVM/tb
BDVMkDPVT3uPDkQ0egQNUfzA0A2Rpwak6RQ+U8c3lekSIEzBmgu6W7dOdfEpE8S8
efX9JGgn5o/Gj176wDbNqf8MmbSegArfAaMOsn1B/om+/ekHDSUheHjU9bMXP7Tf
NcBn43Hr724vloTvlMRLHxO+YRw02wykPD63MKT/I5VJpyJzMhlrvgDA5j4CDznP
CE8ScPjo8uVvjQw6UZHsznT0F7RwpUP08GZXkcS//2K6Zg8/Ugxr9ZkvPk0PHzO4
iHWF9nQMX3FIgs/7tzA6AEG5kovQ/lcvLCPtlZpusRhN6LLlNbSrPKP89nhVBYq+
S5HCNwZR3aOIWPMSPEI4rzrqh6VrBer352M1tPLOvSAWzr5QbPbLkESYJZW5Bt69
ulah0dRmztn6tkkGlW+oqHUT3g4iz3BO/4vEU+RJO8u7lwSOkahNWC6x5ga4EuN2
3KuRQswv4ZEWIlzyycoA3GyLRrsOXLs1zPmMUQoF+dJXOySMHVbtQQ5IbGkt7bNu
CDsZcJcBtUy4AI+0WSYEp0rqeYxU4Heo5pkeqBwVvHrlMwZoU+LADVITXhhHhTqs
g47OGBNXkRGQThqw+0Qp/9k6y5NE1oL2U22S79nxpZMu7peCqRTra2n3S/bxvtrd
Z+3gbUBkJ5RnK0xd1TMqxuPNr4KHGHh/xzedDSQI0gmgRFcfqxHW30EgyMRMite7
IDKdknoNwMN7on6eB1I2IcdeaawPN0TPyitYp2Fk35rVO6CYYtgZ8tuqoJnsY5s7
M3p4YrkJPTahN4MLO9CmAKDIerc20eZ1fYrKPdVH8A8omRZakrrNfc0qIr/Xkx/s
PQA1VY8ICnH7ZPGUE9kE/0sCha61EbbX3MI2CyzkTUGzWbXFuKDt/2UWv2k4RAxx
5JiDk1/4OWrBsO64ZI5zT33TToibIVyE1T0f5o1NvY86PrCZ6wX9az3ZcYabAk1Q
skFyigYXoASI2R8dN01uH44CRZeHnqaLevqlKgSWkP+WWglyjPxlsUKE/4vpnxVA
YGJAMqjx3rKE8mgon+SnZHs0tZlbSMZIHR4U6nIY+zUDq1wz3dg7r/G5mmOiR3/O
9wGV3jywouzOGOo042x4OqaQghN0xXOqdcVxrzckzcDMEkjSH6mHIJs4L0+A77To
bqTzGJefDW1RxzE5C73wtybKot1Gvdz8Ml7cSnET0UKPKIvW15A/apgH61EU44CV
U9hS57dZBEIV6eD28/4hD6uQ6YTk3S8uAGCFY6bh0+KEwBS5iiMcTY1dUMp46apV
mUVZmhqiloCXsMaQQN5xj6cT9gVixXt0vCGfIFWN8pgjYH/BEr3x0jiMSOAQvPS5
WVt7MZ8gdreMNPRVMUCkiaduSBNfLyFJp1vvXPmssSvwTA23lhcObSuJCqWBAr9B
/8uSrfF6HVBzWJv0kG54a02qmcifVPM0WT/if2UDdw0WRWHAolhkctH9bPNqag30
rGoasFuxBap1V2Df2/6LxhIrQZmsu59XRqzAJaS5oHJPhixBFcHb8lLiLx1qD6/o
UAojnLX9k/xfG/Ycso4s+J+n/Z5w+Iyaz7Sy0s19BVa3em5CnaD+Xtf2GIBIIPxP
L+wB2YFYKbX+bTAlFoT/hij3K3nmqGHa6ODA9wilb/4CaHA5g1A9Qz+rKpGx3r56
yeuF6BeXAlW+bo5joCpmjYGQp18WT/8/XOSvwZk3SFvXr6DuSLc8Jk89GnMtE0Q4
7BPP7atlITJA7O7KKLcxVOqhyO01qq+HAhmvOeKztWFF9M58AoOPKjgAhFkQBy0r
z2lXG+yt7Ril3HkLGP4OjjXoLzjBGSVXvcDIs2WwFS/AhaCuOCxHlmQy7g3reB9E
Gzvk2+Z6iMjdFYUW5zA4U+fv6aN5jK4l0OmT7McnYqxl/L5kxCBXMAERUtoAZ7+y
aAQJTR+PhmiPKkea4xgEd3dv8YC9KIvrTd+5TcZdnMs50TPGNSfOFkt0wBAlHte0
e/Y3DZ54SjPhnA/vgISz5XtSz2aPQxYarLKLQXuadWMPq3vhDgRAVTAisN80GhbT
AQ8BJNSoQIoOzqRG7OkQHVVp04EXGbn8peQryXbn1w7bcipxRNsU86hFYIr8wx9L
itY2mM6mLQv655yo/+qsrnOpNISy9rLuoq37WrtaDVHq9bEd8n+h+zse8ptXXsQh
HobVfQlEQk+h965IGSNVGKFwYerYuUCsz0ct9f+KCnOGToRmBz0h+X/Bzjd27ZWC
8mRwVtDnLhIMPwk5qTXXTkjMmAq6vbJV0smRSe8h9mUGdDZdCckrcdQfeD+PXO6Q
lOjISJNsVxY7cjfmHqA5ZZQFjNj5wIus++gARmIau8bBoUepYJKyG9zh0hbd+5HB
fI5TCqicLhCobdm/jNJeW9PXgOacnlGZ6aoQpUW8VJWn6MXmeFoI8HakVQNZVUeS
fnN/EyYTxH4Ygz/EZIbT24GcecuwUzUGZnTg1tMB7esIBCr3UkUyrOtGqbvZswul
xJAeXiBEAIaLD86mwEOseagDc0QQ5s1NmVB02ul0jV8IqC3REKIg16NPJ50IToEr
O7TbAAlAHqmMaf4i8TBzHsLfmVI2hBhAnQM2CAUnyqWKKRPAXY5TP5aUkE9NsI/5
GyV+2ThnvQ2wEkzFyZEwqY//h7UDLW5Et67FNyPmf5F6dme9UvX+C3fxXv8DwpK2
gBIKMIC4r16L/sGI8eEGjiFsAFODBkvjLTncS5pAZOkwhmbSTW8z7LPxCzppKnve
d7AldGmMI7kh+jQCcN78fDb2yUn2kqzhDfO2QuSJq85iD8AgGtbplle07VfnoLAN
3Fgpp+5V4+ecqtzmzBCkXUkm7bw8/daypAVKSmkAS9X/MDxQVTe3vnEOlCpKfIaS
7N8a8MvFzCD0huFVRGuOaHCSdjBeNmktbf6VUOhMQnGN4NGPR5kHVFi9o+IVOt+z
gKf7hsahP7LSJCX7SGT68AmqhlUBKKgqfigi01cwa92VwnBmwH6cR4ofsycIn4iG
pfIT3vQP8hcmhaQoT/WQuTHgIgruGq5/THfchHi58wRtKQWNSq2gVMdg5D2gvg+n
aK0RgdnbI5SJ2xjkE3ZgQ1lHd5mxProYJNmGw8rHXyULu6PxJ8Wq53CzwD6c99xY
AoPjOGaIsxSsJcX5S4KiGd8OO9bzlWXkdgFGwLwS6Is1RmmjFrcDQpWba5pP4nrS
buKGljv3o6iE+QEl0rMkCcZyN1ha/+lSvqw1/Ae67zmArocBmyX2xgA7m2QFsCO1
Ld2EnTk3o1Q58eVM0WPWDTiIAOXoHqF2fKps2Ik/W9PGq490NEPvA+wwURWx8KP+
RW2pIQfNyplvLFWtkYfy6VyNYL1ShedzELDkwxRtbBdg+HTVLISHbJO5tlHobWjC
4RORJA0pVPTxca+E4HUeyXjChYXN5ZdUKj8e0FWUhh06NYJ+8giUEhwN2uVSYGFu
hybbmC8CLqt1hXLSXc/LFc8LfgqCWSFArl9n5u8I8ONUic0s60pmI3ywClvJ0G+1
13ElFTppzUm9PfNU3B6CslfgHchwgK+AWR7Wvh3DGJgHN+xCr3+0l5dGReX6iVRb
spIiGK+risrCtumrgo10UWZfQ83ELImsxnoVRQV5eK0Es18WSRkMYzsXpf3zR8FN
4DAZC10i8pqa9z4D5lXTcubv4EibvvNHNlvYn+xTqVUrMkTheK1DTYCOu97befHN
Q9V3gSbVeGFyYMc48Yaqaq14UGRQnINt2ksHG6IRG4VjX9wQdBiWgsRSF7654yZm
xoDsyflciD6RkOz9bQzLWOm1aqIspAUjnjxOvjsTELrgJlosCeil56IIpsoO85r1
3pNFZSJYvGVrIrtP2gUhl+FdMI5IxiKWrBA9jRpOGMrplmH3q/k+f9qvXRP7yglT
sP4tOeLRxayvDvBBA/J9vcMucJmGLx9rnEKEDih6guUwoxrYSPihYiuDcHb0nrlK
Op1iHwuZdkij5lfUTbvtfmcLMeFPR+v2Hio9ivHAmz5EUFcWKt/vjO7F5NYWAhUa
LnVXwt6+l4lMj5uL++p7LrGGMINrEqkqMi7617lZGkbReYu8HMniQsYWl6/z3smZ
noeVM+KPz5ErW4VI0QwbIq8WUedK1Jtt44egc7gZGvbBNn4CoBoYxFcrKNftEeJg
KX8zc+rdk/z7nImA/KzWm+SnQRQCgLjWtLiUHgNKvDlLqHSSOoOIsgprTDagJc+r
nXaBO+cfwkVG3cyWrJ3oe5wDPj8h2IZrmdUl8j9aEof2idP6lDSjbcEr2mrfS4Zn
0ySMN+2PtSQxnNdwJHD2WX5Vc9o6glU6I16dVwoXJlLEBMd4qNJv+1NCpp3AablH
r2zvw379N88aurozbgHQH3up3XQs7HW5l0A3lGRc/z+cEqkiDc9c2cRxopdQa6zZ
6RTSnYlXlMjsQ3AMepQ2jUwS/55wTXaf/3+u+bvk+VOoJ/F/lUNvaxq5sM3MxqoF
VWruYj2cgnf3TMJsf+Pzdd8PiCN2fAzFDeBP1AIh1thV8roJG6iAdL4rqE/JGFKw
4I+clM5efrt32Bvp+sipWK7TnrwAWa2SQpACbA+jB4SVxpiP2vo8r+6rJVRCUvZ8
sXP4SJQe/QIezWYLHRcDqvOvW5HF9iE9iwfJRkrQ+IjLmw2Bo3A/bzKhmk+2pxUJ
i/wvndfk2z0yD66VIDrrUxqKR+SM9ws/jwJCgzMilj2S32fsUmHmwLFfyTiOvwPy
syIoSV/53/Y91sZX39/ahZGKLWMlqkWDaAoJMwpIE9R8gSOF9mH5YM2pMCptcOY7
ngs7uH+7II6cBUV8ddyf9BbpcCYoX9SNvcBW3PU0o9x3dBT3viCRxRg5Z22p54VH
nNmm5lcEKi+Xl7SHfSYRAOhLl+INXX54P8oITco/RCR8d9v7e20TkennxpRuRViT
5UwHCaKTZvD9Dro8Tg0uKd6tRKwOb18ainn8jpnjMWkmINPw5MEfclKNLp8RUx+U
iD2cwm7L7I0jbDzSdfeCVLldhH5R1wlgH/2a7hVZEzpG8pzQueIj08sZv2+IlYe4
JQKZISodCvAILlPrGMV84gBCRh3qfo3OVNHFVqzfoVFARTYwV/1fYYcCKAhThhnv
sNtxkQdWozMhl/ENhdYPy6PT+nq0L/IUAy9bxtUP/dJm0/3ivEv8jbSXxMY5iSxZ
Ym8dhnradbIyLFgp+9lFiZS5z+oPeDOFAKBHGnHaO+iTzB0rapZRXsb0kURbAqg7
YWwEDG4AUqmreyX8jzOoVgskivWEwLN+PyyLWbVoMRP/SKP3Y6zutsERTTeLsn7J
1UPlD3vYKUxVmirjp+3eMv57gmACX4KWC3V8llzy0GUEAWnIlH/fKuviSzLXmzpt
AcS0YCZx8k/srRJ/nhGF3JtzOVkJGbQ/eHGVV+VmegG/IRXS3t4ZhCz670qOH4Gj
2Nw04mS0h1DXUsBZYGqwxEr9CT9+ufEGIdxN8Z1t1FIW8ZlmqY+m0aNhNUt5cycm
Eh6/qZTVMxtnPX40yeGmP7VOe4rZVqYjyV7zpw5tmVdRGufmeDrUBess9D8EWLeF
qpKafyNDJMtuPA9TZ2IsLq29Ax5SqZsbIfmnkKKBeUOhzsN79JK1hurOFW48JM2a
9UKVAFbdAi5pg37tULaIhZKaeHMWNiWpa2m3MC/3nu900CiCfhOiMTU9T2CD5vP2
oh8Tm59YckMLT/OgLVoDg9HYlRQRTvnfkwa7uI7d7Iz6qb2mrFmW58N7zO8tuOqo
N+OiCxpiaoclX5JhQu1mxJl9p/vjgVCryTavhtbGAMNvTkax3QnD6vb7Dvv/yezR
IUMEQeRh8pkDk0TsNlgetieeaol4+C7vzAI4tXCf/HvzNcIIl/nn5NSzRepqN0eG
6WUC8928uruhibsKmV0v7DggsJ4uInb8/2BgPbSApFXHYmXwYX7Y2T7AUry0kSCJ
LTAfDLqzbtmFGbBiu3JXTgQMeEqyrDMyRFsPYLgaRjkjzVkU0yvJoMrEU6rbo6Xh
6BnLea0qPBQ/+BQatsJORTLFhCepDGtKENvQLS1fgap5qTwyIeJd6u+wYAaP/Zff
TsQxvNR3BZ4M+p/yDEVDNp6ajCQ0zBIFaB7QW6ZyeK2vZyCMsOe0hmsKUhb3/WUP
OS5gghJKfAQQqS9ybXnob8e1SUoJIjYU/2JZfOH/6BxTNRwSP0xpsNKYOzPV5+rl
6dd1TfWXp2YyNG8J9Aiu53Cb+7dOpA8kboWPfhA6xFS7lZ7IXgd22EDP18wyQnjB
A3lmF8SKt85Lp9ZOYa7MQXAkeggrPiW26GggoOtTCw/v3PDNr/5ACYzpOxEx9qtS
U0WnTkCceDaGUXH22zu0czgQpCNNUeGD1FFjj/df3moNMTw2rX4L8jijo3D7/qiJ
FeXjQM9PaIcbxEs4DLfmlXc0v2p6z0QdyYTTQJV6VNOnIFfE7rze/O0kGlwke3SI
K6DSYHRsCxo8lbjuntvAMBMnG3CYVznfDAoIEDH0Gh72Q6kMOjrY8PSIAWQtU+/B
JMtdIzVfWNd5R8VIzb/4lGnpWwWbnrwENptb+IxEJkT8XW2gji7xBEiQH1WMVeOf
OeHw526/yhLkR9J8AU6OWlZPHGvJEa6Gn1ye+QO3SL3vdHldCeR1gVSECEXStQwh
8n0KSL9HpTsisROjhH7PzLZljeAHUPyqZExRqiBMaucz2L4lTuSJVrduXRbDB3JD
BMAy0LF6ZEZyvnVOpONvdR9IK/Kt/uGNJZznEOZVr8zK4EUBka10ScL9+nyXqfG/
BjmP7Vt9w/LY7PLdhPYTdg04i1n7bW9XM5rJKL0bNMb27GS0ekq+0xTxks3o/dRI
z5V8pQgEh/8zd5DRuO/5D2Bo7UROMyTGxZe4ovmby5UyA9V4y55Mo+ryky4uIh6K
g3Yk8F3kjGtW42mQiKtUwzdcwdqVYIBEdf1OHIKHPbbdt4HjwDuD4lbxyx3plGW1
o0fgqKtjNVs8pAMGhxUI0oxuBteW6Zk6Pt7e3PVc27uvGVATo7Van6J7RC0w4my+
X4QnewvhXsmzSSlz0y2g5HebrVDjNk14WlbjgGcP5f0K6/LUT7HyKq9uC0uodnZ9
O2GIEB2xHa6tD1EVn0R3Vf9GKUMbA1Yar8BamMVIWzV0FbAhU91BzGbO7a/sLx1r
7yeV9I3Cxxs16FNqjqNHoeTjx7T5Hux9jEFWI0/QfY7unVrf+qnaKzkfNRqZ1NfT
8vPSvy5XiARkRIAfLGtwaLJjDAV5e9q4T774Vw7v/vojGeJ39bAd5h2sgsiaUjbW
vp10YwiLH5pHRWK8pzAWel6g8+L9mpc8qb+H2BJ6mtxw8AW17xYE5b9uoxxIsUdQ
5gpLNSjtxwivWohPUme373Oucc9VLdgOblGgfE4kgouXlCs6Tf3CK8IXhICFTkNo
HyyXze2kh3oLSif6uOloAJOnwjaZsG2P0vmvPx4xt+cRE6NDjSppN/ssgGCdzue/
Gzi4jekRYwMhjv+d7OjQ68bpcLEYBcQ1uo/8heg/k/2C1DH0eefkwud4V2FZ7Bkw
ooYh7U7eJhgggk04GQIvc8GjpD2o2hVTFMtt7Av0oAfT9obzOAtuxzT4DrHB8Xod
FVGhlArfxd2I/QBiT8TzXJxk2p0zFJ7jZcYO4/SeXy4v+aQVZ6ChvbqYLXdQ6pBv
bau408mX482j+0bzws2g241ltZczOYITkPK8CCPpZcd8vTOTSZIyxEcrIPaMNEb2
xA+ggcPxc1EdUbGNWzuMNm7B8LnFSNsjXmBtF4qbkaUTUcuEfOoulHB5M38xP6f1
rVWZ+nXJcCUlPQLUy9SI0/aHBlCI0jwY24e/66ZdrBWACr/9uT5TTrdUWapDiyTs
KW/9TFh5qPGimPbRQQrQilgAED7kuOzafiTnqGVHq8GFmqEVBxxfxuClvj1yvl+d
RRxNeWADhoHF3p6Q+oACIzF8gnCfaRnbF2PxeWq2QKbet80gcWbUDernKY3X97ic
t0/7ixro2LVYiX81QeNE+iue6v6W8sTdLi57/nAQvV8Q/O17YcN/8nTucu9/uWHj
mTwQ8hN1lRqi5rnJVSx2U5kC6Pn1fn0rlCPyth8xwM7ilcfJvCfqIlY8VJxuFJSV
Ze24Ad6zeDX42y3bM+8h4eJwIvDlfk7zx1em+f/imCBTx0gRGHrAtpPnDqwtv+Q5
DSBlx4Moucc4Z4gQ0mSSA42sdwPu44Ij9uGHCnsLkFhHjV6kmXzdPT5zsLY20yL6
r0hLGw8iQu3wlgvOJOTFsMK8HjrYLk9kqAjn3wrhy/DHbc9aNyP+VzntQQ/GzHhM
XEZmZyYbjWc1N+OxFxJnjGWA9bhB3BaVWrzNOOMcelYUi2kmIPM1i/vSmv/y/wDa
JS8JBfP5YZeNQsY42sZ9k7OrH3Jmn0paynB6bbnrl0/tl7FzX4l9y3gDKoxMPqFU
VdINFZk4Y8CFy9/u6DMk+ZrQj7deALBk6Ofi7jk/x0uXQlrrS48YtZB9iVaK4u2r
LrA9jsjxP+2POJ+kh7YrP/teHkbfz4y6DGNT1byjHgwX8+6veY3RP9FkSiQD7rk5
jLtguJS/5hMBy1KqUEH3NVypwHPxWQwvWLcR25rDKEXAx4qNIsMmzZ+6Qe6i/YPF
RriUcriKn19FiSNg5Ny/EiR1hDa3JBF55+x3jdommu+uBfHAK94X6moo+zOJVGed
DXg0wFsxBf/m2yQt3Y2DQRDvZ+y1RZOecYkB0PB8uAxI52wicLAOvt5TtFRme9uL
yy/OrrcWbl0MqPZcP0nhNR4ZFucu5jLIJtrxV2G1WClLDo5j/VeoJ5/UDclkhmyA
m1/FCccs5EebYv1R9h6CUuIZfIins9/QA18dLG8wYrNTMtlStOUUz0OsuP8CQYxe
9xyLzgncZvSYuTXCGgseuwRmpfg7yuu9i7vQH8F5+us7BXjFL2i843rJNFVJyAw+
iJ/kTyBs5ZtFFXFDHUE1gt/58DcaaMHsN/t/1013f6P5mr0fjoY9UST+MgWxa4VQ
elW1xDDxccGnZPXqRpEo5t3MZ7hEprby7+g/GISfC/3YTAl0+na0SKxCST3OeShR
Tc/aDQHFG9fPALzlWSyxuX6jkT0tskAyzsNe1sqGAIQu4VCAZaglv1/10E6EU4DK
UhSCqnuNMb3XDc0yS7qtXDjlLW2GhQnjwdLYdICG5uA4O07YELPAXHQXkRX0HNsh
kwv7Ssx+zawsfZtDEtoIe5xTaQQkrxs3aYi7ib78PYErOTc845iLCy4WYOt3y8KE
CORTZCpfVZbFoCOIJO1FAIYq7jQjB/7uovhRr6YXkIueMvhuowXbVansi7fyxu+v
0OMkVGZZReBIMs7Vavpbi3SbyBj1iC7c+3JinCoD4kUlVbXhks6+UFBSJUCcgEPI
qeWDtHUz+uS68ZAHYqv6PXWrDePv1bU/tks24KgZjtbiQSupqn0ul7suoYl9oTy2
63+JaECObXb/Y7CYuSh4ly8tNWmZVuQ1pk2bI4NGcPprM4GzvNB1WT0gfEd/F97x
ARatebB7vUcpTmN/JjpoE2iD5GcgLp1ZyNsfrC3163pxS6l3HSNuml9VHVBpT4fK
OhJhEYLKqw4Av/+i43aVW1Gdye+k7r2fdbhKOQYLQLAuJuV9rY9i/JzlzN7bzirZ
/tTzxWdF3KJA4Z8UnBoFLKW1HWY2yBoTdSWG46oSzYrOzaM07bV+i2v2js1icnTl
XvdAwbM5CFMdj8Z3S+sb/w3aaqo4GIBKuyq7IfGurxYe3icWsK+ynV1RcqM1J29J
5pYhe2dBYrNQmSVHioEMWUZBluUx+7X27Xy0jGwuCdtV/MnOFlCuKPJeA1gcu1kM
PuNZ6cuSdqDBNENbvEwZIjehaDvPDV53K/otZUrQyYjnY7XOTDPN/ygfMlkdgGJL
dXH7TqSkKkXpGa2wOiqomNtwo310H64g1u0iTIcFPSDcD7N0ay5t6nVsZopQDEWs
a2iRET3nV3AMBK0Dh35Khc+PxfHsjbiFs5FvcqipCgwrAurF45WJ0kZmK+r+9jK7
4DvmTSOnqOf+3D0W5UyFBtU3AhWNMJmH2mz3R993/CbcIEy5IyyTNOBNOpIGaICN
xegGRdK4RjsSXaAU77uXoohEJB1CwbaHAi6ai0kcj+TDOq10OdsUMrAMb0xRfr8s
icQ92P9NJqOutXFgs5NrX1IeMSgTriTnZI/7RWqFGtsFAfKngk8+FfkWfr85f18H
DSEa+a6ETkIXbqjP0C9tTA2gnHlQFKji/tHpCb7GHj8yJimIJgOOWRj+UfRHAh04
PE33kaqqPOYFQ99ookbluakYcttLu7NjyoBOxiT3HhZju2iWY1jA68GCT0L6Ig0U
wxcfA6N7iy3VGdWbIP/bKmmKxoCP9LPdd7qd7s/9c+7ZNft/tfkRkYFwVeIivNnZ
gMMmYGJgTGYdrLJ3TB0+5DB/eDGFGro6cRijEIXhFRAAtlRVjVDkVRYsrH5rCGyA
Fdht8bUjbL72SDFzSvw5f61Gw5dngGalGNalaVF0c7Tc3+LssMAI3x54A+l30zU8
nk3Fr6Fw6aX8wy7zIWNQA396Xyu6o9qmlfB+gKODkq5NoV0URni8LG4nL/oMeJ7e
/29VNwlFu/f4CM1FeYqvf7NToqeFCiYl10bFF7jN6B4t5BLFE0K2htcu+ZY58zlZ
8VvB9FetLXFnhjnWkbQW7WxrDbZ7zkPLbabBv8K6RMglcnyWaKIt9m/v266+ZMeq
Axi93GB8RcmRl/lDFO9ob1WmMmhdzgoX+0R86fs56kYuEMcN3MrbYdJK1Irinukv
Qujl/QsNJCUB8T1xTYeF3LW2ZyyywBOdhLGDZNGkqZtLLv2TCQGf0NRP8T30MYBB
5NHYkQTx2HQ2KD/N/Vzrmv6gVcXkaYwNkCXTetKo6PvdJpCd6bDqJFepYagJst9B
6fP34wc5M3reVNg2pQrU9XTWH3kSO2p6YDgxuAUfekk/FpqH6TE9H94uEjYQ56cs
sxbL8567jqujhcP/t9dY3L955XSwYqaqzDM3bpq9U5cpEpUQDQp7+KLsBo2/yKZX
mUEw/hYHPv82qCmoheYAltpK5Mh6smmGMPahOmbi3V4k+MBlpsmxaGy6gWIqFGoO
4vSLwFNy5NvaU/h4GcIdXH87hwpR1YXWJFw/wz1t6D3DWqgH/onykUsRGaNKqdjH
kLoQPQ6L3wM9pcgvqK3sq8LONpGIQuAToh9q/pcFCwfiOVbZPDYAqRGQQeoUP0Dl
avh7eshadaHYKnnsm+IcFtIC1RaIVTW/NZaKrRD3ni+5zrbnCi4lqf+FrH/gJfY5
N7D/PSdZrJSmiNiSyZtdHfDGfTv9Wj19ij5RyMVq6EkIAq6v+qwH7PSQfTbR0A4u
+zTwTG0f/Tqdy/fyF0loJ3C+aAnH43eEHUFllkHowIVfaNyTOH2T9uv0/Ej6iHLY
N1RDXVKyphJB4RZYSKY4/56EZV08vNaJ+5nU0cHPS+bXGwJCKyHjkz/2FJ4IyhUY
tFWSH0V5aFDfRmVExklWSG19fWlJ8RPjgDRXDMOeRPqIy7wzCcrdj0OVknXMO7Yv
854rTlzin8Md67EyxEB3wsWtvNFJvRVhc9+kq66qFSWqs2REGTN2bGR6TMCrXkvL
e32JIY+LOF1jZ4/9ByCtz0jYuQCCI5N+kan9XMggrKVfTVMAUmmuOFYYWe461ihj
OM+pgqMF4vlJT24spEyje9LFvHR+5V7f8DlxHF/jKVrd+ibCaAytIJaAcG1Z2RSn
GKCuY79LzQPn+MW6oM3CgveNYSbt8K+O5KAanjjdMMeJGXkyIjXHAYa9DskBSWBD
t6+tQ1vKqEkzRQG+59KYnQJ/xVK4Qrp4dNKq5Ho7a2qXZOrvZEMzAczOJga8lt3E
TU9KOyLEUzyE4TasbfU4vm7qIwZ5QkfAk+H3NV5qMZkcmU+gnA1gCUcEyrPZvaiJ
24+jNnae92+MM6Z5l6QSZq/ExjvGM15YksH901vi+VIiACGIuOPU91DbOcAh1yst
jhXSabpoGay7DBGQVuLig3pAp8g6dKPjTwEgDbrXaMnqmwdFdtpPqKKt/Zy8XtCr
VFu0e5A27svVWqw2KOwdiItqAR2L72e8AhxmzEbWacgD3cgNTMZgEyzgKXbTrCXs
fqFyKOh1Vk44aWdRk/oPWe7v2CCLATCmI89AlZ65CdyPXPLY4WJ4bvaipc7qUJ9P
kXvTBtT85D7eCwctTmizYjLsHYmHdtXx4oO7ev0gR8SG460CoO/aWa/dALPfoHm4
vg25F93J5MhNKludVrJLoGUGZQiu8dl/LkQOAOz3fqZnrpS7Jhj6c7Dok+M7G2o6
LUFSXwNU0Qy1PpWwbp+Vs4YazWe7tMnBp0D4yBMlfxfHX13Si7PaSTNWjaT5KN/x
4hgtBDp+dLfLRhEU7PEkgEHkevZ22WsXj4buX3dMJD1fof0OqdqhfygwmMyYASCA
pmdFXXnAoeDdqLr49FXo7AAD5u7ySs+h4UyFnV+O0PsAhbSC0471biTs6Wz6C3c/
OYXuoQyrQnMTMeHeeeDfPsvgqQaYyRuuK34KCG0GK8tOAsFTl6QqNZDDqJSio37B
ZPhHSm3A9+o5pKyeexRncNKAgDCE6NNWfkMPnKRAzv10Fvlq2/rLmq+qTddErVtT
3ja2SA+c13lL86+sffF397v9gkSVFsVLh5BTJyHbzpsQJuRt2Edobzf6eLTsaVrX
b/lBvtfUmrtSDPSasbxofROXfYb0QhtuaeAvne8H99szb6msLE0WwYOtkZAtBx7R
7fQZFGDFxppAlwaqyx7uFOFj9T9byAe/AQzhCLHP3jvY9eUxZccwVQDS80vaZ+YX
GfC/qTrN1WVeUZKNAnUDhqHa1EDX2rZmal+nO7c8rFWSjsYP1uHfX8sue09yph50
IvrlL6IEcxXXXhJvxaOqk8sU0iKSEkZY3vK3uM10ccbqXJbV1y5IDiWa9mSPX1ps
0SechC9OlWFyiHzGdA2e0BcRy3r3B49/O1pKyCHPWMuLVw7KCmveFrfWPBUxbdYM
5isOUYbuKrmOwRaTUGuXME026oBpXXIQxpbhpDLnRfx3yxt6nyqXE9HTyRG3XxkW
2PmBihc941z/NMk5JLOLU3oF2YKJlVCrBw8TCpGpxQbDo4nVc7ujlew1LrMG19Ri
6XjGcJTWW6CM/NF3fa7lll9R5A9Ug8VohU6TLUr7EtqkIBrY/mYzpFm72+0QTpjf
8eMxP8mKnQHCefVwtBLih1qThs8piwlFf20W7DCoBjgkedkwG/bqc3a3nt9Q8XVV
Qun+s6plUBRVMLsO1qhfQj/pfCWmcO/IbVVVZcb7Vc6MUwM8SRbtU6qQ8uAzAil6
ts9S7oRLor4RLCZ9cpPJgn+pqDBkNj3A4lJbLUP/cLlmatFg0WMDsf0jqnBSLUKC
FI9qZwNDSaeOP5DUp/e+zGPn97D6JxtHHlHnyeVDg9Xd44V95TEhAReEAsEVlza4
sAm1YMQey4LA9uynoEF0dzK7c6NL12EazDj9tbgjyAd8IPKy5bNwjYzGJq81DRkZ
2/KktfZNRCIb6kDDjM5xbDhfQrOqNe7S5cQQeoIrUFy7xO3VacFVzhA/JU74UpVp
TeJiofOY0+lCMZF1/N0iQNOJ1m9g+FmaqFy/a9EI6+SCAHRArldcumIcdvMEErgw
jvrWI8T6pMmof//uwaGFGwq0Sr6u254X3auok1+Kufh9SPu68PRRAF6LnV1rzVFL
WmKbSpbLxSvk3Bxxz5a8PcQGq1ogbL1M9FmNl5dapTg0mSFpCCili5VuU35bziJ1
QLdP7A1Vpp8oQxITfuWD0WI8CgOcbn4ve+L/6io46hlP6rN9D+NpcStKYrbnq2w1
Nobtxkuu7Uo8b9vYvfkJHERHM9ODU0OlMQhutM4baBM04CsKCw8dPy0jajo9z46O
P1lLgKA2tKy6pUYtOLLXnktl9JFh4BXSA0POMKuOBgJEvomdJJcUUP+wLnP7wZsp
+EQOlVciuTPpGWvYpxZ1kicFjx/7+Cv/qr/DxAM3Glz3JW08gL057beHtOngz5DW
vnc/hzg3Ox2WauqDcRZ1KkOryilg35XE920z+TzfK1c+rVIwZKFKDxQl9y4D+h00
1ysAob6s+FUp0X49ZgZm83y8MvJv869/3bH1vn6zzHOzIKdvNdtHbAsJauRAdB9t
KZEmvZJGfuzVtWutDCczHpnapKNKBGBKlDxorZm4ZkQueu12tCDKl9nf+G9cWod/
gkfLb96jTRnxiEzduV7FRhvmMUU102iu8sb0nkWbAtK5X2D4Y/3rmH56QLY2hQC5
na1n3o/Hpj0/axIvYSNntA2bHTMd2Tv7+j/h9/90/yXg6HKrf/l0PPu5iksUykUi
8rPtHZuNXbhYZBbioPIS9KqriSlfilRWIudhxjHhbnQONPlvvJlUF9/zW2e4KIpI
WQDnMh469NA9AF0DsxyojWFuHE3Fq262MCpIL6gJD9i4EmEKggVaEcKvmHUbvfkw
rbAYmFZsieYcfPlut/HvaaRDwhf74vx8lO1xwZFmeUdJJhT3K6UA/wTyJwn9YCAy
SbyWx/0l3MdDrdQ0xV9VuiGq+uILs5uPReHroom4PgWkOkmLuqxq9fmReo48Y0wM
ICl9fK85QGzoatYoYzrt6bUihyIun2xRQc5obuxqRRH67/RLmuKT18EU+JCMqN5y
r04CxHu9bYw2Eyya/ngNS8BWWoBxE6o7TGblqI/y/XCg19wak107XZ0m5heia2vu
58F8d+HhiqRTiOV/Li3KnoIiZnWmYBvRH9DQV8L4HreMDXPgx7dmpLDfIvRDedaI
DG8BokFNTmMJ2Zg1cJXtZ+dwWlyfIJIn5BtBzM4fmqwLjhWYS8znUYk/7A1O2ii7
XVag42hSeGkVrOqqcq1C6VzOO/znmwPYlw0/IreO3xnUU5b7ZmPwr695sTd9iUeB
3YXdIhYlVVOwtnbXaLJYmmjF44X+XqB+MjRDW27G/5mEGYyM6aCONnYOQF90ut1+
Wds9Ko3q6hFiu979/b9iOEsIp3Os1BqWIfqC+Gohp3/TO2htg3a6RkCWRDm6Uyds
RT04+sTGaxXzjZ80uxr2B+O3y1VfS7gXA7fPxM4W9c4/kHz2T0V9dg2HI+414AJp
Iq7y1SRXQnRC9Ff8dI6ngHIS7v9xea9stOyUXsfMEosNypKgOgea7dyZCWRdFX5m
3AP8H0b6+eIgvsXh+VmDWRfvYTONIIfmuaoYdE81IqOUduqIoEz8HFKD8fMg+IvT
uV6f4ViC8gCM8Sc9bub4lpkN7wgtaTQQTbNczSK2kYKncGKXVuRlcD4yRKdJFqo/
uLDomxFS4rWIMw/DB+VZAVZX0XADlhc/e18lwGSB3YpXgKAlBLfXNsJh6EiXqeQU
Oi36CRJLvv+OUO9NgwcSoYQPRxur/TjwiShqo/AO6p9alsrnaV5H875Cr+SxgLWt
/MQXG8fLDVGVMxb7EXqHtDwRJ2vqWO/+2Grl8vurpnyZhiRKaHoSVVnoxBCET2NF
eMstS+3ef5tyOb4FfnFQ8hdhQKfAOTj7UD+rdKFnHGlCAj8Bc7bACVohWSB9qLR7
Ny2/NTy1B+V+Z/3Hy0EWjnjuZzhe/jPbNplLjZgdFvVrkEM5TM6UXDY1dN1CwtMx
DrmitUUYY2v7Nr0hfJck7VRgVyYKvY+VAqRPvbnZKe/DL7D0/OswOKbi7zKPwKcx
jY4yslI1IkSOxRrRQ1yOEnpga+tjlDuorWG9MQLVcr6J/RlM8WaN1D+lXEKYIM44
tE7LG7dlJDctl5FZcwEoNLRpzw1OARmVmJqR1VaYc6A2vrbLQ4YZUSI965p0coqp
g7wGmiNvsMSjsW1149JUMuFR8C22B7i3DBpZcZmOrUvmzhOu8m4OsAXE4qxde5k/
sywx/rpuKUxsHfsWPbKUURdvFsHstKLDmSKrCjSG7tj8zYh7ZIq3QgZI9sBHV5Pf
0VkGhKBwz1B7rkwoz5jCwWrDivnRUShUcIeOLlmenM6+x7W9WRwY0TRGuQSmGpZB
4873hUAMCvIsi4njXlcSO7o52Yo1I5adBf8mbgiHBD24znkjX+YfoUxntYJkXgsA
80UuQMiRpWrQ3JekFqTI4ZaRZKMiDAI3Mvhl8c+gA4SqUI8UY4P2YyBjIwaVZgPf
Lk/P+VV5J6TKUE4immIaRREdhyc8+Vwojss0QYRKVsZdWwjZ7geoVnA0XSLLIzGe
q1xAv0bRQyCmjXjPmb8kyyURee7uxyidOPPfo4wImfd2+togXcNfE/oCBPbm6unG
Tn3v47nsH7+x0dMoDu0Vs9j8CFQConLFCzAbhx20oSTAltGQmnayT0wbFLNIJrLc
Ezl9fKJCvbYgpBUYf4zi+dkgWME5svZFVv2qJkEBd0JzsA/qQKX/tdodwX3/la6Z
6IVg6EVqbNmGg3PX6GYpeCqTWe8ab3BUxFn/iSxyzSQ5Tj0OUk9K8unz7zTNJUIp
cBPpTwUhHF7d8dqcQJlXtMsLI6Z9pfrFayXCBTk2dQm45qx626XIfTX2sm7CyvOC
mY5KhPH275LmnVk0LlGAIeOPqdkjqG0eAFDYTdf/W0pzhNYDe9ywfTkqfuZFFyLK
buNfWExAiL6tUo+Jw2fJHv2vVd5rcYStBn0i18Nb8zgFq/+X0bspi1CEcYH9d/Or
+rfkK4MO5zy02iHACg+YhYxhMGCWtCx4LIeczMKGuR1mJVPdzid9nEmWJe+V58Fw
vWWcG5oRSszDQPTH9cm8JTGjdT9GQF3ptnXgTUSWkfUtvdC6S4GiONyCVsmieUHt
/DcFwUcu2YHjk2GQuaKlqQ8c1udPYWBA7YOvt5yPjJy1jdiaYjT3c9knBVJwCrJL
nXTpmXjpPanw8Hg4joXbcIsUe1seyFdJOC4z6NEwzGRFfOlihbKiC2FiTMk2hJHt
IuG+7WXQH0R1/fvw6rZWwij0QGz7jqhoMSYd6XrsDkqd12fwnzEUmP6OuBvbDM+w
5b8McHVqZe3pqbGAJP/fFbebJsiffsd8nzI/SKl3nD8murJMD813H2Dc/7uqWqyq
FLoSODRSqduvc6C+L2nWcu3PwWNh5/ZItFGPX8rgo7GPb5exIQyGR7c6ImZDbbox
yDqXHeqtdfwwkWkAdxxOUULQ7ai8KVSWhZNfaD5MdatHTXQTEfuYIpEw5pOk9gLQ
1EJ5ua94029m5Iv99+74qU7JM4VFax9cL0nt1qDdCczZ0mK5lQBP7lN5nEmDESPV
K3uiLmFuJ8MOKR76VXCOH1r9euKrSh5i+cmlcD0WItdLIvqJ97TwGooxX/vNsNg9
RgzcVfsF2U7c9rGuEDOAtPiq4zz6uUgtpIIWEw5DyqlogDuYvOkf5Vl0WCEXoPY3
MvZhVnB2EpmjEoIqulWIBnvsxBd3Fpmx98jp7OV+QHhICBfXup/lZ8H06uPrBxBG
na1fcDhQJZ6bX43bwgfU7XsLJX9SQMxfxUTeqQUr7XkjGwGDqL6xQy8JScKYThrB
MZEadqBzwJA3rR0soWj7KusBNQ91jnP3PsSxNIAl1mvOzrdM+JywR8d6u81FiAkW
gEwdGtZ6/h0u/aDQSwfTFFIK7uTm3AAWdu1FGocW6s/MAo+IL7B9QWZ24mrlC5lS
By2HB2cYe+MehwlKuyZ2qU44KV+rn3I2Gtdq+6NHX8bzwZJOneI5nrD/nEVh2QS5
RUO7tL9aMUMxzJA0t2pygjqKm7pA8ybjkqZ2Leta/CfQbx0tdkZHY/yIIK27CmCJ
QxJPeyLCM3jmgRmKf3WiVBQdkDqTmA0IM4eE1Gr9USL58w3ahjh7fuWMtFv84gmi
NpDMFNReI6E8qUAmBfYaACfyAlIutjhqAXc3HslU5Qhg3+hn/7Vzl/N0TIqKw1oD
XmlIV/gyGpDSp8k9YrBmZdbRWG6486DIt0TB8w3Xpwb5Sp0a3GiLpQPTVgqkHDXE
qElo1RcD4Ln6Z2qg8m40NVn4HbQsmpsppZMU28fYPiFKRsnOBh9LkSALjruFT5Eh
GNtJ9EpBRf/wOhXCQtbMp6jsJb/ivBuZfsqTwfgJPqzSwuauoHGmDHmG+j8klr0c
AyPMsbZ2oIKJs50WILGH/uHdFtuEceDgKROhtpe3/YSYYWRsVf+kQ0kxIt+ot/I9
2d4og7Jioi2XVmbB7G53kjsLCEwYWLzqlfp6evWVIb393iHBxN6snz6DvohAs0SJ
aj2cSIfpzxZSRPHDBzZC26wGuQwMnL5hcp5nxNz7c9aS6rLNasThTulrpTEY6oIO
BBnIsMjNHvng8fO8dhdULFqUt0OxbQ1ZlXLAxIqByqW6IONjqhaM2xtY6BkEYyjM
UVx0P0pq+HtM6pUKrlgEJVQmFwq+pKVDN8jtvhKu6SGZU4wuKbkcDmmdRAQueveb
1f76f0lE/cKTXOvFPgKjSLl4Nv3QV0cmskC44rsVb2jr/yrgJrdloi6Otl2TuzVg
Zje7J14/ZCK3wkePmtnZIK3Ga8KcCBcS05ujIA7Pgac8OmS34u99MgOBZqs2jZlT
GwUS+4H4YPGDMgVaBwreOelhEXbnmLRhT/PoH5JpJ74hWkjQaw39cvlIIBKjlWuv
0arfSN8X6rwrrl6xrizVN1HnDecMOdwnhcGwFtNFDfHK6vLwBur/LaMKhHcKORXH
twi4CIKMUHhya9O/yGYdozljQK9uGIa6HvZz0DrKNYh/zyDsru0tDbLz2M0RmN+5
mgT7yyzBl7FV3/Y+cy+AjV/X3EQt9r3Zl/6FeUiito1YdlCFso5U/pslov5PhaSn
PdBmLybuwr/QMgTm59Wtj5foRi1EdoOJAWSymHD2iRvB8kpo+4Hj4mOtqcxqoW9+
wWX0jIDckHvKb4zBf6uP8uXibhz0meNBwsFtk0PN411LPQFVcUmhve2qhIIXHlaO
niyOqLzppJciG6+O2wqjE+jOYpoTDQEN4cw+LmVGFa1vh6XgkXug4eHeE+4T9KyS
vdfwPA2Y4EH7+US1Fh3poUO6+fmDywLDjRxftFqNEhjuiwvzAZSEmI51h1G5fSWr
O6lEzuoLfia8h9U8FX+Qe6wDlV70riR/5I1rX/2yvAg25FBu1ua9pIs8yF64ijub
w5DBY5es5SGVKAoXNuDDQv3Oy1HHedEAYVepLuk3qLi/Pvx351O19ulCadUprLyG
w+oFTlQfct6LDxyOw0CK7vFZWWJ3s4qaTRopb0n7b6LbUSBaYvrG/15l1hmuhe5N
kVfLiZrpiaNk32Vy13K5NfPLUnfB11Ud5iDZIxgS2xIYhB/r2FTDklOh0SJ+6Qgt
/hplcB8CrkL7YHGHpTkyZApHeg623sjjw3YD+nGeo9UjPT5VbQSk3icom4SYnL56
08aUtvPl8RfxhI/wLe6uuf+GO8kkKWjpRmtnw3fQbzZyKZdpXAxMd3F7iByVvG6V
rMlqSaZ0bM6TOoDTRFpF8uZut3RYHg0veIC+SZ7nBZ+pWZ45YBiN3on3SOn8n58s
n0E99gc/S+BkWm0aVwWY7IH0lGiHNFfXVWZsIHkHgVuDLHgf5hg6VY9nB89XC1b7
C9n6etEUiHRQHUn8S4d0IsitC6cRziSsiOoU0TfbB2f3sw0dBJKgcg53yDRQNBhN
iSlLGTUYIALItVqp30l826Zr04UcptmRsFYFqmYyJ0UZ8j9LRhY9abNqkZqsR9yA
fsrxawlF7+GSa+/oG6t2kNmchpPbhZJ61Zm0zodsYOleOpUQR1XCka/unVXMiyAs
v6gh/NTuFSnTmmTXX+4e4c1bquwW879LBqzRxzvobLWVYA7YQkyadmOpjUTKXYKs
mia3UVvL/MN7R0E40YMOITGZMCO+BckkwG2G6U2jVd68DKVwywMFylIa7BQpbgRp
vOUwNPqJNQLZt0x7zN9gK391FHFrF7Qf2kSEhPptRfRvmX31W6aJfs+2b5+tS1It
0kho/AcREaIeLpqLs1rweNFcVzN6FsUw00dzK9ErGpTRfCrDTtvnh5gkh1rbPlJk
iAQCeMw5j/Kmk54+q8geFlJIX4cCaWz63TMRG/8q4P+b/v4vHeId82zCXXf+DFl5
o/XeUG46zzvYKzATLUIRZ0Nt21CU5KN+I96r8p1jeYXSvd2vg9x2UL6IvRblbsTR
qay8ct8vA+bqQIEECq1TiLON0NOx786lYrDJgD9Fp+IknaKHdxHhQTHbpbP8XqD1
31kPPDiVaCRDhmy2TMLLHDzZq9DILmyPUgsqcnayqxmFWvUoc796c2I4rSK90Dvl
IcBG9fMtDiDa9lFmHDvlSdnuj740evKHoCYpOqCywHEfUQtODU6S8esGb3cLgkHy
MBrQZ2kd1kz2aKadfUxN01xIHBBQ7S0y1UUBYdWJlRpR4nA5huzAks65fNIDghvN
h3YMiwef2aFkRvYM8EGPhBFNR2CJDNFXdiis/l2ehSwG8QW+UvvqhpTDG37m8knN
TSUqz3rrS3lQ+VhL9k4DmoZlLNJ3DHfxfrYQT8RTEpqwczX2bIEQgYcqQo2TP77z
zvOV3Y70XvDYzCGQTQXtzIFenkD9GMGB5czsvLdvcRA6/7YilbrAlkzbgNHZpmns
mOGGziLieIs0PSA1l8sFPNl2DfYrjgn/dcCSehsKSJ9ycuqMy22qCCiCutFS8MGR
fWNqGt1Fggty3Zw46O5jUdtwbJgRHPHE9+qyrn7YDcmIpbKVfQKUHwQsDJ3+zeI8
9Uqc62q3sINnun/MXDLGHDEhSm/Zf9X4+2ARZwMyFE+F4XEz5vcBgOCta3yvTr76
Nkdf8m8VGJLe4Q5H1bXGwRORRz5Ui+skVl193L9cefaxXH97Th7rW0OOuXlsTxXb
1Xqopsd/4flPrhgWwdTkcsarGvNaoTZOHWCNHKmGDnYC3aOrrCTx5kaKAfEF6+mk
3WogCl+TC8d4vtIMlSZK3330e1uhU+zbaWwjS4s0gk8tWz1pWbutmYD7coe+Vr5B
mlyQjUxWDH4N6RM8ycQ0d1IDJind5hPvNqcqHEZx7aZWr7JAyvUQ2TFtLZv/Wyaa
1DTbGsdH+NXfLyg/u2wZ/dh0RJmHjupJY3wGYXWC0AK5xNO4TDjR7TKVwT5BuYWJ
BqkLMvRTle9WWQFOsxT9Gj1U2IgpQOV+4sQHoYm/CuYat2dLe/+cIMTnKD+pnX9M
Rf/JkmZvEAmxjxXSGS0TRTQsKuU3JQxrFeBiT/PMoqCpk3Zj07LLWDPoyj0eM/1k
yA7GJ0/598ct5ZeLpwwnwzz5PoamQuGN+TxABZav3b0J5gBJ1yuPLConhE1jc5ER
j239IqEepe2xBe1Y2bbnYHKX5HbzUodQw5NB7VlrZECnC1OGJ2RfN2eerFq0WJDc
v+Lge/U/x6vEb5f251xtgtyvgh6bwaQUakZo9q5q9PXATtpuNmjBcbkbrDNYQnZw
yq5PkuJtxkDqeF5yVVoIef8eNwaR7jFXMlAJsp0nLoC9nmSIOoOfd0sVIHDVFu13
KrA6L1NPi1LUAiaxahGim1aNobegUTKXOHyBxezbJMMusK9ZjDF8bpUi5MZKOrD/
wffyXbT72eQg7paOunonlww/j99iYnoleS0xDK4cE6vGtyLDi/zx40tpNYvTPszZ
F2nx0Bx3SXDJ3xLTE69W/RSwfyfZZIPd6VVJHbn+pfhhfUaWoR3VOB49EPBh2zeE
9t5327WbMFSLtEd0/MYqD/z+96S3+Eiufu1swLk1/XkKrtvJCnu0rD8EPvhOmZD+
pi5XVT3L0Uxx6cVt9u1YIhXKgGIXhxtA0p1Md+wnDmeFJhqxtWdC0j18fnU3fZXD
JTxYaQxvBJ5k/r9uFu23b4UWWzE2nxRWBFuU8QYoVG4DWHBTd9w91jNwiMi75srQ
8WMz7jhiSnTo1ENtxCw7lONDSoQD9BArU6gWjxzVoQObUZyA6Yn7UbJveKQeYUpg
qTHTTuKk26h2dsrt/ZEgkHbDwoZ59wQBZn9lO+wuTGWWLZzG8DUW4bognZk6o+HR
CxV1lz2kzBcxGShwh2HH5ZAxqGVkhvzijJxzB3CFqmIyrf33zJIcMTWSss261DcQ
wBlJ9/TE20LGVtryu627cxmtxWyKwLukNFTO5JYxPfKJtnwbOCyJVorBKboGe59u
2JBA+zt/5qmJ9mOHIGsqHQ9QwRNoXKDGR8UAQNtuAP0kcRMEOfNhHjJTj076pEJv
87oYf23sYfuUhGFloqSUGt1/8t1pXse2m4ouTuX2WPI7tEu2zbaHvPrhqMQxFgu7
ASaDH8k3P6uWHiAqTcGlLCuSYxckG9+IQkzfLLARVU4zwI43ztsRQYNmVjjflkVi
gUDY8i2Egoxd5nDUAEMyGiQ2gdbnIvJEYAp99owzuJrwQuCL2NYzqbLnMDaRuSO2
FGgiYDalqDqLYsVXBRLcxJ2VfAOXtFd7fFgItKiV8FqK62EqlWu5z5Hoct7LAMWL
yaTJu9aD3RrG+KZ0Nho3X4aqd4C+PXInXIl1/YQs8SkIFvFszcZeniZV1b9Z5/S4
9i3P2Uk5hO8W/+uIE0gBaRwe1mRQaHbjdhPg2AeCEoI+NjAvzJPThZM1YXBkqVWz
Nz8Pcm9kD4D2gV5lR2/WGko4T/iE64ERJF9+m2oZTVObFU6LNByqsqe4RIfjGtzT
2mptR0pJJ4vkWg9xSZzqhH/MYRtB45R+0CcV0UjE9k8+gCEWtFbMrCsWrRNSjosv
IV5lyEhktRxx2rGvai+iRaxUrEF184F4M/9eEB9lY93EETKjrwouV23s6xOXL1P+
BkbBdtTxf8W85+9j+mFtusWwsYW4ffewt1gwXK1VZntF+upnWLHTvpwvPImfeaUc
wHp8xiftXi4pzKrpncrc943KY3T7KN6aldLvebev0nqOSIRhBsy0rh7BMYC47ljO
NmPgFNLACraIOXAlU/O93FFE79tD5qCd8sUDUDi6WatztBIzWPkJQU6/KhtTU3DU
wOy4m7X6+ugiGFY5E8Gdw3ZOjXN7zU1vA0gYNGRnCsWOg2KeP/KDUMOO9OSIz0v+
OT6c7N0GL2paI+mtry4EYOjkWjBU06UVFy+r/1NYu9cRsbrNwsgJjR+8CU8Fns/k
r6YItCdJMLE0C5Rx4p8lFdtxkPboqlcQ+3yge9J1xJ6Jlye5tmXY+nWc4CNK9Sbw
NLQD8Lrk7hz27ey1LoFsjrLyMRouXDf+eL5J4VGZCG5h4TToXATULFy+r09rUQqx
plak5r8di7TyPztT4BRAzZA6WIfBzTC4vf1PQnp3UKwIrQqE0OP8oJixhbwrXdBd
pYAhDuGf+dLsM5Q/HLQFCGQqJU97yAvPuuamaZsuybm/1Q3qX0t3aTR9L2neYGcb
9xF+n3vVTYCTQpKIcw2pm1RBTmiMQveZkdK++PtoKqw+CIGMXMk7sGc/MJkdxOrh
K7bgkC6OeZpQChtbCllQBw31EqpOXfb4YYXyNNAHQPdpGxhUNMlAMYaAQ6zgMoDy
eMhHiMS31oMBksunVnG726KKR06463SmBmPWTgTgdo/3541rmVIOhQWZLWNqegDK
WFATUUK9BR+/3bMPJi53OKpj8GVXvELQQdXBE02AoHJhjwjR92Yahi/zysFMNpP6
IjL3ymrafnQ2cfwXnQZQUFJ4EgRm9sq19BvfnvxqIuhqtME+vLNVBHu33PAgnth/
NITXJDpkgJO5gU/sRNWWoYvStkMqY+xaMUVbeg/jjtkB8ud4Vw16MbNr1LeohQ//
f/c0vat9xwxLrzAC7iy+/j3pogjnVr88i6qIKhSWlujwW0BA7RPtDSJ2QDxOjokj
zF9aJ4eEF6Pudt+hklJgxAJeAD1qwWhzp03pdzqejNWqk/XGC3joCsDiXr/BVbmO
+w1LGbbDj5hUNI/1sDWK5AR9wIS5td+dM2/X1jk6XUH5LZ3uP7OZJnmEqWEIARL+
J0n3uj1SDWDzL5c5rTIyWU/c2sXJjsepQ/MhJAKDc233AARyaKHHZHCBu4rc55I1
A5RrUyxiEY0YDZWYpcYtAoLxgT2VabzXeluxy31uN6JUFCIubRYhThPfFeDv4Asp
E/Fs0bqfs1tVP+a4a2BPQDqki4jMu8fNEqtY51xUNnYDyrO15PMWkEbGXR8kucab
jLyqqd4X5cgAGUsUle7guFQ4Xs1ScZ0b8OSncDceUUeg+1ohikbDEdTLlbeBkDNP
qv9qdhwZvAI2ZlEvbQD72OxdDpLv4y8SUXgISgmi1jLPpeAt6SrJOnBikznLMaWz
/5i7UTab4q85hGuI07CSUPYhlv3iKU8SNs2I+rIt9dDeEcrDnmE2y+cuT/XjOHiI
y7IrUooHlW1/UaMXZkEZ8wyOp7NOppaTn7qooIVZ/ikDy7iBL3kDMUym7pXgBbvp
q6D2Aj1T+jdZmj37GyBZNOZ9CIKiItqd05PC4gOvDyisufwexPsd/45lEFF8bH1G
6Iquy6/k/hBHFLx38eX8xL27NdoHcdpAYy/PNr8GH8bsLDIxJPtQRAkIRnmJHVvC
SMGeWFsaaRymcymjdtqw1qwaXxr3r1jNrlGN3TDsBGVPXvOQ0KDVjlTjrzPQadZJ
Zpo7HWij638bH3j12N3oanlpT/B5o5tE2LFPO+PA4tsG88RpNmilNx3LJ6yBLad1
FliTO+H3uyTfhNGmxdOaYNkHj0cy5i2nGf3oEpej+rpndimyanLCGYv0f3ra1PGK
d0Y3H0bAORZ7CsU+OozCK2FaakIoV3nIm3MzMi63FbFtNM5QtjikXFz+4mDepe95
f0b0Lhd0Yavx1N/ZPPmeSBn2vwEPpsBHm+lbTaIz+umS04CX4Kj9UZAoPtFHZ8XC
5P2yobcbsLjVhZyf8Ex4OrWop1WW9CzpagWdblmmkO7ocxF00fwZ40P72rWKQKbS
I5sXUkM8AlE7FS/t67fVLGthKXgUbw26suUXepx7NiHxxvGNyjyCY8xpEGS4nFoH
ZAB5BFW8tHW4CHt7bwRMYS93EFgD+BT0KiY1hQ+nKW5BzQ2WvLpkKxKl09bPy7Zf
WDZ3Z8vaCG8utK9357zyBA5eMqgKY246V0x/eTeIK7buSDSajnr3njf4B81hzFMT
Ww1DUJsRM/fJJd20Y3F8zb8Mct5je27dxeKFBy/3lbFh+pAKBo/Fx4+gmLXGiWE0
YMEs9JTFq1Iv/zuAwKRWVPg+pusPvCZHW8tBT1LFjkOXycCx9aDIJMYd7N/w3gix
4STAQmAd0s9iazaYW1GqtSDfa1VUZ84e93ujzzaIsXC7BdzsaGe6wLQpq+7iZIti
pvxj8tbSCqJWlutGZEo8Mg0NIDxl/D8VoMTrpOqAo39oWh8zooh4t9WqV5RQfTfc
tU9kVsOKCAmWyRBvkOao4ZPvOvOHz11EpG43ACNt4DPH7S7BFDkTnwGlirZ0o8RB
na6EplRy6fpb/5t+txQvuR1PW5z0zjRXDStWyFE08hbYPg2pUtuI14XHY0h3Gg0z
WQHjppr4rKDRr0y+OsJpXRLj4ATcTKHpwAdJdL4oV2+Vn1QAYXcc+tXM4Noo6D4z
/HDFnnxT0WfBI45ruwB43n7fksTqLiJJG6doMLZJ0aA7SyTFCbSllDpyIA8W3MEs
HkGG/eGljne2wVmzrDk4tVy/k9Axh3d275uDJ3+llXimUxguNCtIoS4ykCYP+X2j
be4mT/7oKIePYVlOkaclUXszm8fk0iybEfQ45ezL43fNd4D2fhyGUgN6xMf2v4GJ
6E1pPulqjVi0FR035+gi+2bybIyWdzyaNNm+efoyh7UJ9MFYDbxlLW8ViA9rSzgA
m27NcPlpl3FKY1uiEX9WYn/ZfKebpkj7LaaXT/zHAtWam4fuUvesfdzW0kcfSMEi
6ty6jetR5OYUfsM44NqlJALWHVTayhSuyf9cAfK9wugOctE0QpSbbhbgZ77Bpk0W
kfRXjQ68k99C7MtlFRU+9O3u+tSDmL+eZ1ESwSkYb979rpong4XHV6j66W133Yp+
FmYkLVMC5pQMVBjAL1U73tOwyF42BFg8JdKBVodTqtF4/ZtkQJ4ogaQymJsCsWsj
UJRSQ146RydC9zYXSPomVvD7qxJOMYfYmaHuOGjlgHET5b/EFQIE4ypfNRVs+hlk
YfQgSmYHghOQgyJjP4PbOSoeSiuk7qdKO7Hp7Jn7h9F6cFxvKvLptsJFOZ8zavZV
vH7gbn36B0rwxB8jgnuxkPD7BiO3l4ekMkEznti62fcVPc1gPiqkiB29baGZHM1h
IU4LI6sg6eV68Q7249odHYeYNUSgC32Zc+//gRh6Sv3JDUV14o9I5yQBufXxUkj7
`protect END_PROTECTED
