`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cxrSn3p9lK5kQ+A7TaPoKBEMgb0LaQP0fEI/DyybkXd/wXvOsDpsUA/MzDxYMhiT
7t9v6+DJjle3HCu8KNe2m3TagajONMKbHSsIJIP3NqRBNe9aw6xMH4tVpFwpt4+9
6DXaufS/ipaBrM7d7+BvSCT3IY4T7alB3As/mqYTAdC1jKWUNq4zAdfutSXZBUiN
dA7jgFbQicWx+Wy1KQ3DHcc/CKtwE1w2ie6AT9OwN5mypUvHCic7oNl2hBwm5Tvs
OyifjaKPC7UwbgY/C/O+Y45ZmqcZOy25wThfdwBSzNhYf96ptYJuU6hqBlwrmh06
QR6YSfakyrs2igaIeOzwZg==
`protect END_PROTECTED
