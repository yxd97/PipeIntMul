`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1rfcC64qLCJLTph5oFQaKVUNsBR/EdQiihjEuMBcpiWSR7EXvLYwS1cNcth1OrmI
y8iUjgVGgaz/YcIJFYfbGTw6yWrRXnrTJ8zGIktntyB+ynsOa9QxCwV3vefroEEI
qY59SQkAeiqT1WdzVqquM92s1meowtnupOTBy3YwtKGDKforBiUZDYaFwaSWhYap
Ts27c8v3IztpCdecssn5BQSyh9Wp3eydrlwinig1uaLdckH7O/Hell8+N75WifX3
1lfRnlYDOeTLSkSepqlmqWP5lCrOt7U09/1InxhFyqbSvJAgVuZ6td4dW5pFNbeJ
4cL3af9eAoCm6XvG5a5A0MhBmZ7IFBp+4w66n7pQs+CzJ9+2bhj1TtEnPDbpgbJq
6rwsiqWUBmftS3ioWPvov2vzFsRtiVGmUkkCqgaerGndJDt9affROS4TIYSbDfyu
zFgE5aRe1tV/eLtkxp+mVO6HEbWeE2Era9fzBTI1ZF3X9p4qB+8IEwdz3JHCEAvu
Ahm6nrUDB/WT6rpo3UuF7NEZZNErAjRWt3bymg4cwpmhRhZzA3RcOtf8kkQb+w+H
NktF7rFZAXsP4wpuqtTQi72ycfe+Z9uAlX98T2CfNa2YIDyNx7W7dJMZ1rHyN9pl
ffPXcEcDoHQB8Sscc9g0XOeTLBAJaWTNbD0rnFWWCN6lR5uFzWCH2kgcZo+8w6/Q
Y2p0fvZxeMFvnXusCRqD9mBwEQBtKqWBDgjJwoxVsCAzKceQGDwb0/v/MmBi37KN
L5wBTnPi0UwMNSqt8O8yZVenkbZ5XzeMyqAB84xGRCTVU2WejIZH2Z4McYLnmm9r
cDAxbLnKr8YQpyP2Sm8E49tpDf0tgJd8NaSM+EQs9fNtN+PSBLMmG4ijy8Z9ZQzX
Uvz3TsejORZi98gR23kj+w6J404gGDT9cGtorCShN9Ox8RXzQ1BAM009dEyunYQ+
fnBTsX+SGTqpPSnG7nLtQHnp3KG/p+eHAYxPwDXnnaoX6rb7kTr+YNVt9g4SGsTi
+7uYOZjlwx6djBE7DO8/j+ZN64E4rJtxca/9+qTJRDW9RmctZDAOGP+Rnub/qlo3
RELX0y6LC9J8MmJ8qwPYATND5KrzsFw0vKMl1PY6alYru74llNcFbicPU3BMu8fM
SutlS9TaI7+hK7BJwn8IR3UMJqSBN8vjuA/zkG0wgAymJRBdiI49AfCPshAg435U
ptVxo37QvP9vwLGdNZ21GMPREaIl0mNk649k1fHLFAcITswdDt1I5ikV2xJ9t443
Mb65tbWqiOA0qYRS4lHQnL5SowfnZZtBUCpvGRN8VT1ENWfjlnvQn/hKzTtapEDr
gKCt5iPZzVQy2o5lv9JsTrsURePaBLMY2PhOK03k9Rx8Z09fpLkUg6OPv9siI/aO
uKO0J2nEHMDi+ejq6JR1LkPiT0TNZZnH7qz/EIk5SebmBbEhZ81kGj5NOMTHleGf
nlU+pXL6HEUQnK0NeOUnIKKwsWBNcjeF4/a45l/oTf+KvL8kz442DjWJoU0gE8Li
svbmizzyM56WB09ZX7e1OdLjUFTtCOzvKtkj3GXmzOFmktntgKCvglLnq0wwFNDw
P/CzzrnNurh1/3nEDOZ1DsmIoRl9o2iNoTAfHkdXswNolSq9iaWJ+wn0VZAOiEMb
Ihe4iHzhbGZIugIufnZsCtJIO0MXAY/0Ipqp9dhjdKxZBmP6ISHk+DF3obE6LbJn
fFUvfslrfrEaUoMb/hOA8cYv5m+xDV1FjzamW4dk4xmw07s78bI0GfjoRpYuoknw
Fj7rRDMeB52yXypuOmSsIyJ3W6RQBZEtZ5tuBfxR9PtC/R7aicH/5ro4k6aAaSmJ
bTPd1DF9fmhuTfnGY0f5+4EDI93rGuJDZVIfOr1dv3+eBKVmIVlHsM7/hwRZFTLT
/uyFM38aeA2wyEVwmOEgYNK/15ywbRniXmxQl93s5TVpivnkgO7/KUN6QFSQtcgA
SOavdxNZHJOWGPVp0OLecqVMK1bq8lti+IDHrwv2n2mSORSvLIevY3qEx8FMVOnC
IQ+M+feYjvK3XjGWswZff9Y3By/JN+Wf1d0P4wFPHwc6fg/hc6zarhqTAIhrTPYm
wDGSdt8mnGyCAT4F/sFcMIldcE+lxc4t7iyc/560UKhVs2g/sH62V+4LfJn3W+RN
l0PArGGl9qOqfRkyrh61YihChF5ME5dvOVrlx1V2K+mPq4cSB8duc4pO1ZNW9gv5
PqLBnM1UYYu8zVnR1Um5f4Tx4ji15IaRNtAzjb/+3e+vInMIPfO8dRp4vPDLCcew
xoHv30KdvL8GN2TUYYvnco7TRQVRpJSPF9GwdSfx75JbYJLTfepu/foZzEb/9596
1WluUZiDEeG87W8AjxGkW3XomNPAWPTJczD5jjipQ6t4HTCdllMw6pehY1XW3PWL
D0UzLAF579RAEwkMHvMflO5sV8kfj9wohiRuWi8r6XTIC4ID9Reb9ncfpogsfM8K
SXZMb45SsjCYEJu2mkqi1Z+6J/2OXPd8QJkkkNFl4wj9t2D8/FMa9GwyAPuujjhX
4FjvbcDBs6UfvyMz2CnR/qL6GRHdVMWMOO2KMaXfLAwhz4kAugwIes3x3OBOnF8B
wG4h6KbBNxbBKidFJEsr1n5NqGdOsnzmnCDTOlpuAqgRRb/hpe57cTMrdUpgKYIu
znpBoP3qaYGyNHgvP8L44cXnDBEm2CHhn6y2RVkXL8zH6Qy273FtlsvyxRVsyvcZ
o3rnhM2Rc2wNNXX2BmDfkrfc0pCPuUvYKVbuU42U1pvPAgOvms+wdx2HBozNrAWr
HIKu6S05GNjC7YaDXw9Ox9fWb1LK8Xzofcy3fEAbkkLj8R2E/GYF7rouHQW94ZaI
MWOsSXlDpAZtA9R8syrCSJoSF70AMSy9Zyi1E9doA5I0r46kEhNbbdHHmMMHN7wB
gynt3Ws3Z9l1p3j3r/qXrCSV3xWIrMhqpmAixJu5lPRzIHcegXxL/LZ6POqYSkLS
N+N47RZWqmus3Ku62Lgd/rJ3fBauC2H15S2PNF2bt0bZsbTkMUkV1CvRcSwYumtQ
MRKKDG6k8A9EoRrZZavItH3Z/Q7IiNq2mWqiRw7cvlUIlxdQRwBrrSg0f5fOt1Il
IobsigUoiH1/Fr/3LcJaLIJP1AtNa/fdBqP22H++Thkh12rZ6/riV36gaBqM+F2T
/CxxJD75aLkg9u0L50P5U5ZkY8yYHkvujb/n7got7g2gqQlMc8ZxOxih75hE+oUI
WChZccF8N5vrq9Ud3utydLGca+N3xnEUpmmLMYKA34X2kd0VJ47Cb/kMEXN5EPET
eEp+C9VmzwD2/O5I2oMWVgFNV1okMwzo0AvgyIwUslJnA9EgRLMjKLiVP12TdRGs
H3pzVG0RyRelyef/wG4fmhWrcroK3wpoV0vGU8eLsnC5BJ9HgQUsr36uMbbQm2dI
onX5BCmowjXK6gDFKnl8J40rvfeKLkhqXTaEDxkc4LVq4fKqBaSmJfqzmag5R2Pr
pHpXWucjdAx2ykZ6YfIn4Zb2xltDjLowcy9tXdTMWeAKGQfdZTXVXKT9pOYBC0L+
w/rjuFf93UPdfTwCBCNugHszK8zsoIYlDip9h7GIwTIaOZEshtQGS35lsxRKRKpY
uL/dMLzyQHna8jRSqRohb5uTrFvZbEuyqbBN081dRt/7V+mmGZqMT7iuG3jDjnmC
VMBqPFN4cTFBRuRPuazkgVhi47nQaUUS0rFTsGs4KniNH6erIS2dmDtxeoPrnL9k
hstzlSEW/oQg6hllXEs/GdNod0u6WF5mzKevH7MD3b5M7rdq+pNPuc8g42fsck2/
eImwrmy3yEEM3yFO7D55/m4DVOfzloVB9m+Pg8rf4/rXUALscl/W9ZcJRM5Kt37a
D6VCWkZfAPAagQt53OVZYluChjT+dzB7v3uF6LTsGSnYqtvpO+kw+hdsYjQqKllf
r4KE7GRQgxDAxtsWjcwDJ/rFyfsj3cbks8yhiZinryntr6a9fpKwF8gIEtD+oBx+
71FLfKa+khf5Kv/lbeeHQfOiYMgjkT8CckgfBZTxhdKEGqjkj7PjkukGtMmHUXxh
AvZEq75gnUObyT9vM5wM/GjLa3RkUTTjFBmQEHkBbtB78k5AJ01vOgMlUU/PVdUg
jqnCDr3F47h6Hl65DgQ3oX/o7Mb1NtCVd6voYic27OfH5g6e2FgV+GeXuw6urqpM
0GRHF6IIvEmfCXE8VxiOIws0RKapZxfc2Roj7912kxb5rTN3jG9TYhiRc6+/7B1E
TQpwMep9xEEuboLMKBSw9+fm9sP0ODJV/BO2d03IxE5zhncCFv5LpbaDLGVsADF0
skRfhhg9Mld2VIW99mwYoQtJQIkrl4NllzE45sPSJexyBp/WulgeF2Ow1EZRYtC/
mGC//ATYDe58yHb2kQJniexiB2Ikg7D2KhflTwdlXPwD0laGVJt2Kb+HFUbfK15X
L3MVJZKAtAQ+Fggon+JzS7t2PMrVeIgvBWbDUtB+v50np4Z9bE/mMgRN+jCbr4s+
VXezVmjXLRuR3jEGArdBZ4UVJnMkyHT/JPf30yAplFux+b1P+7RghvH5+9NbculC
jbUH4YcRzlIGaeQAcEqdEHExlgkQiRP2G91vTX9dSMjA3EtbJenodnP6Jjqkowwo
64ga7kPH39bVeAEXd5quFo7e7t0f7leJMtv5uDtLUQkoQxElWMeMyqvnQiqF3GoJ
UlbhxM/+4eTQFiSOw2R4P/gWnzYjQ0jTFKTEM8wxM1hdttgXv90dVNALXiLb2g1L
CxtGDWsD0Cvfl3uTCJbJ/CVNEKcPOM83XAMAM5HyV2kTUwBmtJCiV90wGTxlGjDN
btOzw8R3rgl26uAz/wlfVrzJd/LbMHRgqcTJ1480UuUBz3hCGy1PhTqfF9Ps0sU2
LZ3whi1XuES5mSiQQQo6mCustcyIhSluhrEM35L8Hk6KQnWHJr3b2iA4+BJlIyBv
F5S7Ala5CcU/mUCdf7q/K8/xo+R2dGtEVPtB3fLY5J8AlLg9y5bsdBO/+tQ41qoP
oXS5jLK4WcCdNJFUwIaiKIbsyQBY7KKiL0309yhshnm+/qZXDlimmfXOhgHbSV2V
GP00abH7/T7VpARrszlu8tj/8TE2ViGxQNqqVZWLUA1THlDOcjrjm+dqtLgJLi/N
W2RBjnkF+zke2I+tyP0GzuLfFj/8plvFlgvFQ4J/NQqMbHwACfXv99aZ+c10OmXi
t2boGuQ7VutMi8/Sjo3JUioqJJPWZZsWctHu7dmoRh3qUkjRXEiYisL4RpJRfcTZ
9J+kwmcCAfktZLseXOg8dtxFBNMcfV5jb9v19gxGnwqPgRImXF9U8GZAT7H05Yqo
fnjRHt2t7MCyjVFyIH4tvwRe2Mq/aQZJPOKwHrDUOoZ43ntRQN5hcs538DcufHtp
dGprluobmQkvCTzONLdNPLascBp6y6/aKY5HLOIlSDT0wCeALYPynJ8azS0ZUZYy
cpalpQ/g0eRfNmTOfEDWO7D3UfUj6bP+1IP/PVNNCAig05Yff5QHkjD6cfj8YYPS
QYNECoWoqjPJXaHnxxHurHhDmyxSwtXG7feaC8wqicTd8GkvdV7FLr7YF67NFaa6
S0z5r5yeILx86RVrJ3f1hzy2AnsAY4Rirf1Rmtnd+Z6lsfYz3KDT6ikqpRb/HNyG
VGQXgOaaBFmUybjNGYcAEIThfKCqF5D9M0FjCATSa5wnCBTvze+U72kc7QXDNKgp
Na+NNWg2T+HCQXng3navUF0STavP54BDXayo2bIHjpkYWELwKbOgMHjVayMLKT2y
RpHB2wPTgfkckX7SEfQizDQ2iSTvjaOaXYXByAYqzbGDoclw4EbAwMiwAYfBnx+K
pJ4DkyNR+ipoPhCBYXOf9uVOLn884S1ulrH03O477K3Tls+K7fdbcmdwD9hbh6mr
kNcPmm0LeF7W3WdLffE+HmLmqMC9XRuRTimXNBhaKPCI6QwcTejYNMsgoHhlcTJs
jtUqyNUX2q/L98x82f2tzKEdFVnKiiZ+Gtpfg7nBs2NLmQOK3FXM1ma7Opi0n/hS
hz9FS4b0GadSON7aIwjYut8erng3KZRXzS/xhB4QFidlb6pZx0cGZnECp4/+y/8g
+KfrqrCu83N/wn4JdaCOCHtRl3SuATdF1hXbUW8+Apxt0HrkmOM9oIAGkexw1pqn
WxQTTVmRElW37ClER0gKYQC9kt/Zf/+oUeOhVf/38+CYmTUVUoZGbqrrUJA+4aIi
/lRmd4ctMkOXjiEnsaOts9v4+DrrxuyedKRamcq2VQywS9Mg1PFmC8zzX+FzUdlu
ALa4nMZlhcNfZXiI+ChidCuABqbWyYINnEiQeWP/So750ftjqK3llOdkMAV2erf4
cgApl59cHMCDzLbpo5FX9YiC70S+wC+yyKwX/Fq43Elzfflvlk+8Lk39Lqbnqu+w
su0r+AH8KplAu3pzQtGRW3ZMfqtPnh1deEUUNcC1/Z+Mh+r0V9aWcISPYNIGkXx8
bfKh6eunNEF0+FSE8KjRQNY0qWBHD1oi0x6Cc8ydi3EKtyWKsUgD4G67mA3c5p3B
x31uVzZRnNxj0poTzdtJ9Pc8AE3fWu1jBO42jxbUFKdbKxth/2AzGe37EMT0Cpg8
IN2nEpxgpM/Q1s0bDE5JBpkK8gqPDKxH6KqHzVeu6sb1RnUPnq9lkcLq2PKjrJ3C
HK3DeMrKAg7Yv1OILf4u826OyXHGaIxDqtXHwiF7V5r0864/MTdR9yGoF5NHCkJ+
QEn/2YAgh1fQKfuLL2DhLwDY7+6WQV9IFZBrFvSZ/7aaIocQ6h5csIkkjEhg9AjQ
hcUV/zHLcO1P5HWq4EQfdDRtBukdkKcEjUo0CWgvP2i+ktYbepz1M+qCWD5ZNINS
2/GFSIBihxkqCJh7Pa4b/+5y8mzqbeRZOqsLF10ABL+uV9BCsSMCuXL2mnPJqCmy
wOXh8bo3SE3bT0yP25lqOKgr76DcCeb2JJmnGQm5tFc6WrWtdoRJENvlBILpPsOl
vJiBzNY/gZnCMd7UUcJKuFv0gMRaHWdax7ciP8k13tGtwN7WxPe80vXnlvhyqawj
LQM11Zs3FszOK8cvV2QSvjLwcORpkrnMnuA6E05twlr0DntHtmdZwvaVnSPbmQr8
zlSbpN53EnJE9zExLZO1qi/tVEHEpuAcTmNpkCizg76CV744lJeQGR7i7E2ucY7V
cxwlIFwcKlwKa3/+ulzcekemDeZnku8HAG+aqkIGsdxf9fJ0tH6xafrva/xq+bFK
poTkLt6KMDefSOAhlhhbX1aXAewtIvUgUz/Y7uKLkIWO6CwNVQ4y5mMVTSCbVt3l
w2ijsdh1ZfWZ0Gnpt54nE6bJP5py1GePgRY5JUqj5iLb71YM+JQ/lNggVXYNyR9q
0QkAfqTEJQ0e+geBWDDa0qyA0zGUOxkncn/uz7DSG8SJivKkjKlZntepHYESsigb
UuNjkJIr5g+nYEQWqTnaSFapxVzOVQbTnblBhe9yvkcrL/J3CYWJUIPK7i08sDFa
3uzSPndV0MIwZGqlB30l7gUWdac+xZc/hfnC2LPcyiLe8JmS0AAL7fdL1StAXiCc
6CqzImdNIrnTftalvaQhWKyC81goriefDD/ldsOmIWPt8Et31eadsLtwnHPVVNHj
z0jSqsmbylCWZ0aecBXZcjUQa1hdrr+r6ibPo4e8TSp/zwUdpHIJ0i/VnO3zkcRW
NFX1JioUEG1A2MD+nFU3p/+ai7EZgH+xYmtNLoQsRv72o98a5VyRbxo2AKi3Fkx3
iSAiUM92ZkUyQ7PYotDMXNwFVEV1zzeTwZRPgzAlHxSMdEe4IUk3axGkXTK9hpuP
fWx5C7TJjjBkkoaxxWzCAMpn6pLrqSBmuY/QKsHMOcszk/Qmwzs/PZCNaHw5AbwV
zB8oB9rdjJkJQ4/wFt7SkSdMxhk0Vpe4xmd6vp9htzhmPhWT2sL8zhOaX/7hUIzq
RUaRX2+UiYry5kHMgrTtT3Eh6HFPCNaD2X6updVxgkv9ylaGLct+f890sfTJwQPL
3cgM2VlGdfB0M2v1XIy2AKykfqlHeuhVOZYU5oDiI9NYzeFuWszdbG2UwIt5eqG2
jmZQDLlQW+tHsmTCjIDMf8XN8w9rFLdokRS51JVz8e2McOWKS3Ho1S/PLYdB8B4e
DasK3rdMfFxmIZa8SsMz2uxpVZzgsEkjqfmhzBTas9eXwIFa1RlzEDmo/4tUdM2I
HBYaq9083fHaTxFsWelXqxyInoFyzhfGwZTfkla91A9I2aeORBstUKBJZDZq5Ps/
R0WdaEUCqhncuTX5shAYvBrz8D7SNcqo1LmV+CK9lg7zUIOyMXbuiHK+vTPogti9
6aVxBr5d1Be54G6azaBkdVmSYiTtaXeB9ms4n+n6iacvYPShWCGt2teQbzuEE5HP
aCZg6A266OtHj4G58TdzaERMYjeMbnwd3394rNeizHGdOPiM4Szn31+67oI1dXfn
N4G8ntvdIOg0WsXQnP2MlZ5Wl4AGtaDSC1ViYQBnbnaU+c8fdGbaamc5LkjsStsX
nvcZdlWfRGGtnVCJgAqF4YWD8NcEoDCM/1q7ikHsbiiDAO07AU+f3aZjgVw597s9
7S5EYCZTTJcwhjGV7GfbuPCCO+NZPsP7FnOUwJW+7+csIjmp7vShFuN5KZ2beyFj
Mvd+epzDNlYPYej8+PZ5xL+eQzftqgedaLBho6f+mA2cHNLlEjfj9sRWVhTp6/Af
veaWc/PLVLLSRyjM9+xh2sBUrPcv9MyGW8yuStnJZ/ceI43HKN/B1D8n14IZc7x0
jiD47/V27u/ky/+mcFmdnpddjgPDH8gghqpjq3jY0TTLC7n0Dq5KsGYjZaVFWpNx
MnjdpVYxcdt9cgoXdCfEjeDWG3LwxmoHsTIy9I7kKWx/HKPjNgaTYMZ00fqUp33k
oJGK6XT3iwompktp9ThNDeOQB/mfs2mOxUG2WsFRcVuZGi3aFb/l4VriMhnsT4uj
aXrLeWVECTr/jJfdW/ek3MOzQWAmrmDiG5oPG5QzBjOTjdCZciBatVIrtsAAA4Un
j1NH4EWBe+fP4IMl8200jQUemm8HQwEEMMF3Oz0PgcyHAFWPEACZ2lq707VR3Fnm
S1q4//algy/4ktK0nQfn49cNgfrBuf9Gv0WKplX8KVqPHdLuRM2CWRIBMti+z8kg
abcXAt8w9SCjahGYWDLCfWtRt5HEtgVtmBQhxbfwf9MTKTGju6ZUVL2hnptk6Pv9
G02F9gTwQhkdn9uOapmNAs4EXstkvjUtdjyVIrsCxj1y0gxjqCQHzM/KlwX3JQ40
JAjUWuxQf6AkZGVDWs1fPkrRyGPTClplb+UPgRnPhFd1nw1xeCs04xRBz1sjfP/p
2sNw+fbPORTR7r2zXmqBhkU/7uY0tnL5jUFRl9ltBeCi7yshQkwMmTrVyqVe3yaj
owOq3cyeDvaX4QNwjhavc+FtDmdoX3MWaw0uXZSkgf9eCBRWtDkNwTsO6VzoY+Mp
RCfHN5PlFGPDwH2rAWEZcDlkKKakbFbMTU+MVTbLjHIxq79kFOA4ulbsRdaH++a2
rAZnm0fso69XCz2LHMaTVBgMWAoHElis6ULOZ9agGPCkPP02SqRVf9qPPESpt7KW
hpfyRAi4mxr2hKKiQIPNLWOx9I+pp/1TKy+qdIboQUsEku8PV73FFA772j2o9lmJ
2Z1QGuCX4C03RCgdi9I6GLyYgSR9RpNh7E9gM9hjBljpR9EukFABGzfcljwlGeT2
Syg3bTFg0jG9vo4kTEGpirhTi8jWNLvTciMsfWKFMaK3GJy9g6whgM3pe6xItC6P
1eX2LWd9k7euNk3xrS3CRzcp2I5U6ox9aE08TGlevTwR6eeU/0UKULIAFM5kz0Ml
Gw3u7w4a0pzEtY8jnnyjCYJWFWotQ8vjbCYRFnJGRbVgxsvkRZcB9iXx2Oy9n1in
cp6qQw40I6SiI08KS6MC00xgw2BNMBu6mZ/el2QMT0dWByRgnqSZ2Y+DxQcVVPZK
KQmW4R/yorcNAmIOoryeMjysxbO3Qy8d5cDDU5KbTVgQQ5AEqLCu0Ilz9mFQnIrM
zMWSAQOSFtshn94iGpH3Kc4pXu0XY6QYqe9vqhurPmpkagtSFFBFIDajFcMmURjd
6YmiKPIeKnvqREnbFEJ9cNJSLoydTLo4dZ4q6JNGslKDP/qdJ92g2v97z7C+b4fk
NK+5VQT653UaBAaQD4CT92OflOa/CrUpXt0rg3L9mE8SeGhCwCOPY6iIl+yy2jUU
3Ywnkgp2vYvzO9Soe0+WZz0wyQ+RV/0iVVz7MKuqeQvrMf1mkfuRSRdMGF0ziROx
hxcb95AQarNvaGc70/lE2GoL1s7JcxE2QKQlBP/AoKjqZvC8sR7+I/SyDqFFad8H
k/OXythwsLqm7ZE2mp1jcwNbFO6jyzHtkHFQVYiMIvCqF7+jiIbudGy+RWO+RECO
lPVHJ81bM+/pMKRsdQp15kRW/Lp3iZccAa+buTSkKXiZQ0p75ZOW5dzjBbaLnX0+
JGq6Fe5gRPK5eLX83ZS3FE50HgrX5qiHXXu7m5seF7lqbO+nvib7MijFgOnUBCIH
CHtRfJdIWOCXt1ba1sShfjUT9vIC6xMz+ZMBYkIEjk8bxNorxLudO3LxPyrlswnc
jqZKV+QbQVTwvhvMF0wdjuGWO4O72KRdQ9+emzOGJ7ZGsE1ukEfyJWt89Ul8JVRB
Bw/f4VzJy6eToh2S9XpP3VqXmRLI+atjo8Bh7vPLuT49+MHaapkaaL8DRrdAYXsN
fwxhinahDPd+nnmWTb7b302b6faqgyTjbMfSLBGEut6AiCfcSsiV0Rcei06jTpf6
dwV7lSQEaBtjXFqtsNISNNk9Ju8Wk54X9xJ/XpDgrpnC2ClLzLU8o7DkDhov9GcB
dj7fv9VyniiA9fZW6Wrj4b27KH4ye9ALywHoCGApBlzJCY9dZJxvNv1YhTAL4CX0
mNVyzgdUbME6UsHvHNbh4F9cmvRfczMt72hW6khgHGoVf/IgB4xU081zcGC2b0tC
VRKKXuBGH5izphkUXhYs4CdegMWY5FFnm9uAhIYyBe18gr5ineUNWI7SHR7FWE5F
71IEyO65DhLnx9PPkfNdDD9W5PH7ms924B8YiApcMMNbQfEsJNanoxUUXbbZt6BO
hJYB7EwM8VNG90wDoQFUu8bc/HI+u0BUtsnCTW7c3fp0pZyYyQeAc17E7+H2k9Xy
j6GWFh30slc5wHxHuVKpxh/NhQwINf4AuHst5B9Ma3uLJrGgI8PBOF4orQV9vzns
FqqN8YtD5FchCPWX9PKrKVgEDHWpQ+0cCJnGE3Gn4XVS3EOBaQ5TYL6j9fp9A2In
yWKHsgy8+mTCdZ8P+vh+UfvkIVBVpVPch0PPF4dWlvcL7O6DlvxVBkGqXutQobZN
owHnb6ySHBHimq7+BeRU5kpJbx0tTkYEgHyu1lQEaJd4XCZOenKB7tD8gvjnROCk
Ot7fX8mknfjg/1gSeV4gp0degDIy/w54j6OTHV5V8EOOQv3jn4sEkZlCThnxv6tx
vGx4ymT4P94m5Cjg1/Lg7ZhYByHJqXXmevSVhbBppdYvHqIubG0ZnSKuhQSUftZ3
4UXXq6Al3NX0pEOrOWvwFdttvlCLwD/j7CdxoZD0/FnHe3gPUv/KrHVxmnYa58LG
pxo1BgErVJPednOm+hibM08MIQ9JN4CWyIKYDCGpwl4kEr/nqisLzw5tkrd5ksdB
`protect END_PROTECTED
