`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PwI08HkQqCxdldHO9MaxMwMZoebfcaL413advOL17XR8DGiAR5VJKuVt35uViTVU
Q+0bH57l8WtghaIcqSVqnCDVGUA4mJd6p3q7m6L5A8FiB+aV6PuagSYER1D14OJT
ncJkKg032nle6fyGNKet0zK0Szt98MmUoqtR5+Drwwv9jq9WsXYMfOHww+3AtEjR
NdbiIR3hzqjynNhmVuSuqim3uvT9Q54pkXBeYM0f5GkwVih95Z+EmssMbxdhqh2u
pBehLJgRsYrVN2smETQqDaUCCY5MVLgO951smPGR2sU=
`protect END_PROTECTED
