`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lMqc7gm/NT8vnvrIMyREX023Y0SC0xgrZjwV4LvdeR+KEpEpi1LFQf+D3OhzfLMH
qdAt6LELWsesIhaS8UomtGzQuuU3J/OHNOz0dcNIZuV/e0K9cTgNj5HnYLFWEvVi
b3UwrdhdrJSfZEohnuxfZOe6OsUWvNmmxjNoqJr+jUvFVukeeGjXecLTPYvM9q8o
35ADbRThLPCkLbu2ugSzWKRuP32Fsili6DWUFW8LEflmk65UzcD/8+7nyjnHrZ4v
rKyHMuBCA0yRs9fNLQBZgCgvaVrsXCq/Gr0TdiPN4QOV8XjfTE/8vIlgP4v94ICz
NiUSfyImWvvaJ/p1RSlh7XXj15707fzNFHaU2hn2SINbsP7dUC0jX7dxRKcWSg5i
EqVac7orPMfjcw2YlPSJAujTqxuPG/VtC+E2Oo24n7DGQsH5n1vFgarmSDUm2Eyf
dinRH+8Lml7Kig8yjMVcs/rlHP6xTzaukfNQV8+TbFUnBM+JcZMfIvFdOPz16mIa
vL+zHC41282gfqKgSlT+muHzEkD0MnSruyznunzdD8+r/wSuS6bN78uvkVGDJcrZ
O1jxyid9p4dNxWCYrcOdk4R+uC1KzdBC2+SvsDLYx05bO8Hh6taHJfg3PFQtKoqh
fM6/BmaqBHr+FLyNQdV0spMNUjU1WbAlJ6cOgv4inJttsc109tLBEQNqd71VBM3E
rWk8tk3CUrr8U0iMBG0NQf5DKprZqOolGUgwH0fL0B4=
`protect END_PROTECTED
