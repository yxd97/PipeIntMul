`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZJtnGqyphmhn3jU8SCXHERrkDUMAHvKds8c0wmWJYeHKeThhiXtueKejjS1edUry
TnnTf/ZrREKhe1X9NT2hVXEXWm1bzL1hCddoUu/AOO6kz4MGxo0FEbsbVTL1jh4e
YHjGdJB/E2zI4rUVTJJnEW6cyaIwWxSpCrsBOS33VDC/vS8kIhBk9yOyF6uTo7vN
bRpzUJsLoRVOMtPf+H969J9G/SCvrkRbqL3NIYVo0piFRzw9YoO27UVUnv1L4FK9
GgSZ0vBZ1/e4VWzXbZOkzNtgw5r39cNMyhJ5k9EEzSE8Ooded7BkPvXKPq5uOMSx
LDNVVIkpJxsfCi3arSZlHQD7aJMTnmy98rm4YF5DFBEn/ggfmQ/+pSyJAI3dFQiZ
QaoTHv5kWzxiZTES3Xd05llstSy6hmsLxVnvDpvSpjYS+I6TDP1t7ZGq1YwEFEbM
WniK+BPCcAzNoSf64VzESxBDbtE0H838+qCyW+T/yX5+jwXTdBmQSmffjw35dfm2
`protect END_PROTECTED
