`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nocafkiwfMMhEuLLa2o6ovUpqpZ7B1/ZCIjXZxuIIi4TxCJ0CmqQ37fEYvQGxTGE
w5h3SC4xJfFwk+JGiEC9lJ6RQS8zYa070D1yqWrwTzGEQFwRscnwqwgZVe219AHi
c4mgvzNoeq/8jimhb9ZAfvvjyx9fkBrHSTLeoMXvzo/sdeBkXeG6bLt09tZB9yqB
B71cKyyCZtnkaqLqk+WaYUpALBSFZowMBGNi9B+WpSU5ZuO/KI3Ce+mS6+AIbxSc
ewIHZKb2+s8ppeLH2YnU2OQaryRkepp3gVtm1uTvtAKCkzQjAmLx+vfYAhSNmw46
9QNHT7EVqecPZAbl/49xL7ToHd13sMdu15crZKVRPporn30aw59uY980aR7anACS
dcF4Dk4ZO19m75pUPUb/Wsmg6NCnJ/wYpN6QK1msFnrloHFx+HP5yUC9Y8GQiPke
5ELuENB+klUh9fNprV0JqjIl2JsbUhfQPC34Ixmni8DXfm8OUNSctFit1ce03oUC
cSCMJUE1gq1E2x/sNyEeAiUOwz9RZSY0Obv6c+AT1xMAZ1pXhAybjd6cir3gYX05
`protect END_PROTECTED
