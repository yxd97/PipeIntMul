`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bR3/2lkmb70Toplhzb4vr9RfuTToBK75fVunH7F+gKrUjnN80WRM7CJ3kK2IDEFO
b5coj8RdPEyuw5SZxY61tkEl+rWraNfwR4qm6kmaPXhynEOUTm/9+FsD/G8X1VTi
AO51VCNTnewJNrhWW7/o1N5F1Jvb+ZZV+JE7nZyQDYFGrtfhOxp//xeyBpKlzWN2
ZhQgOVopg/9s5d2YyCxbMkua94KeCGOw7s6RcqhlGp7VynnsZ72fVa8xN5/A0dw5
YTzBNHd8PJ/FtwMAnotKtbg9EbuGgYORuctiqT0wtl2qorXCk5ohZ4z3Zy7MLNzD
IIUhzjuwRT891AWFjw2bGH1oK3y7dN2I762PdRR7niwHL69iVuyfjD/5dj9MzH/R
5bptyPfI3IUfCTR15VS6WA==
`protect END_PROTECTED
