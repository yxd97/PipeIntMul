`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgUZYn9J6Rr8PiFkTpTi8lmGoD19lxuZ6dD0FwNnWhUM/+alh7kjEuK30kLuLkXE
OV2+tA0Nhx8ERozSDS5gmAy3dYxIaIQHaLCxU/a7sN2zIg2VfB8Dr49AiU9n0EQ8
38g1RhOV3Suj0rtQvj0GjloHXPANWO7OZ7ac4mWbtfIa7XT+9er4Mlc83Pc8jYZI
TYvJTgx715ZYOQn54Ipbk7jj0BOqP9d63mX6sBj+EPLEMvL8ib/jtQaVopqMo5MI
gq3jtQZGXtt+yxPbKlvtWl455J3fxc54MABON4+IelbMSQquvFMr1zxo4OSJ6DS5
19HlBE1wW5n7yNTfE5dxDfwaXCuGk8eNmHm5A2/3t6GxLajpW5lDrucGk8szt4y7
jd7DPTPDioaEa/W3+j476dZ88+XDn04UOctRjTeOGpKNV6ndEYi2gJjeD4MqYLOU
g5//GZPqgpMMGenpvZZmy8rDCRJv01WJut598AAf4VgRR9pUZ4weYac39rwMWu/3
`protect END_PROTECTED
