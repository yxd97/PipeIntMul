`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZEKNM2CPWYJt85hUKB1TudkR8GFYl8WC/SqiDYZMburjqdccBPJy4MJKIyCHPS2f
CjUauTNtHyY94BiQtPyEQsI8wVn6KsgJPAwL2qSaRTMKvxf1nv5aVlnCwjnoCs3A
zVLKjAVNi6Vz8M+U8SvnoT0MMklAtu8j1R94aty0UEqFDPYkBmK5/ur0ufh9jktl
LILEyuczOElaIIGpUG7hCoF/pae744HD3TuOZpvMxmU8fUjsMHtkjvNOGDgxoXYC
2OxQIJxjZ8a6cGbbyf2th7RU/UPFfvNd5lwnNPAoh2ox6mOglDkWZ3KVL/oUjYNs
AEEt9Nrpi3iMIu+nVIIXtCY8hbK0+EEBGUPY7lm6ZqKrxhAFcvyNKTE9p5NJ72Ap
mmCNERf5p4KZektlRk3KXY8Tz7fIqtIn63PRkXheh30=
`protect END_PROTECTED
