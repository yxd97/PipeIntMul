`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GeccLwCgjwIE8kp55aIdZsw7/Pl19+dMzKrtv6nR+B5Le6//DwNkV4eJkQSR8F7C
vrD4p/ejhSZlj/PILrTT/Ma5hKIs8rxhcuVDsHBnLfe5DViHfqStF/LEKq2Np1t6
nSq/Al2AGXbbXq1kzsfC3A9Gpuicdoq/14R+yYaBb9evcC6/kNU3d26J2nIErgTK
bYOlAEQKK9VPfQbc3j2tODgzlz6xBMid6BFz8f02wuwHZlEj/DksSybGN1RBOD8X
Ztfw/7VEl+VjpG6JrjgQu5+WYrXIkNUXs/yIy39pGlCKTooaXYu8zMQdF0IZeE4I
V4s0xu6SvA5CJ08tV2wNs1Dne0RUwVC8jLyJB4g3AuRvsrO4FgzZJMdS+WNhS9Ig
cTS9Ml8DMghHE+mzAO/2e999EEoKmoWkvZhRaaoYDdfRLrzGZaAKTxFlh3etFaZC
K5d0WMSigQarlGZYCFeIG6QgAdgfKGbd1y13SEeeW6vfWnivktnm0E4bYzn5noUf
`protect END_PROTECTED
