`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFpr3EIbKdi+sgeKsj/9yXXu0oreu9Bv4moSfAoscFC+PX402YzeGLxE0JH8GP0p
DJsMKKGzUSPKJ+4Vlm2kNS3Sx6XEWLwcw4iOcRXE/uibPcgzjn5rH7SP36Zicp0Q
5qt8TVz+CsORMCK98cgovk+4KdVq6kLfh2/94YxobierSPoHlqCvHgXMCposvYXg
4mJHAPhOEDhC0qH23KrfoFCJeABSrnGlmJtcwaFDLtee8lwSkYrhrHPob3PuydTv
WbTio0m2ua3ZYdfaAuZMRloUZfQUGtY2x0m2GKDuULBt+aQ0BtLqhDrPNmtxVa1g
3/WkY0QuIexMShLU1NyDsX/qEEMQMU9Qe/SrGI9SVCyeIt8OV691u5hI2mME3tUB
1ww88y9awGN9Uvsr9HM8/g==
`protect END_PROTECTED
