`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qxSYfCzzdn2RokDOhiZ+QdVLlhrcr+kmMihWoatsq+nr+BSW1oMAz2dggn8qrIWr
FpgLG88uAUyQf/SklJpmdjQQVNMq4W9xX44Z4Ux6AP9utN7bRJmoCE3YUJCEjsgW
wOanOGWR5BFH6YW00HXlZOiVny/R8p6u8ag+pviRj+eQsf7XPo5Kyu7uOaLfq555
eDcjJUJQq/ordREqMR/8CiqooWMpSk75vOHpYktV5z91N+q+SaGJ+YVDzg6oin8L
R7LTg9GBqn/eVpHZKfpQesSEd6W+ll5xUy3YywzYTjdBktdx5CaUOLzJ0xdEdqNl
JvDcHpuz23oF9FM2gS2bL1oNp0LjTaCR/3Q58sfNJVQ+sPd5AqQtsmCxYhdjsMNa
UYHPuAk/iu0Grh59CH8DyXTyqHwN7f1N+/u/mRYI1kEJ3jaEleXLoPcKH0g9+yw7
xK22dQe+OyYHNbyVN+BDVxg5XvlaWHoyMIMBRujYjJjIfj+3GZi8DptvgbEBgCLv
39WzZxMVNQ7te/wmYf0tJ6N8LP1ViMwP3S8Ga5bUTgLEkgPMRIa5XA4yLeuHqLVP
NTTwW/X05/Mf6aN8cGTIFZz08pQWqAq6hR3Ory5Sxl0Si48mm2qvJ/+eFV3I09/g
z8b6xpKjIW4Ysv3u7Q04Dhd4v6p7rcgxRrgf8JMfOqQanpGYXxMBlIzrtzUt2TeD
womvL6J2ExdTp3VcbBSON7BnnRXlkhr04CeiLfK7O5YJsh3+Ia/ArVS6HRI+xq6Z
dqdQwvE9d3qdkb2LN1yfNFCwv0INMNpRkBRo2fV7/O4jow0YKa28lZ689H7+lRPU
8lAz/J+CCH9f2CNl+wtKOZQUsMlP+QuFf6XnGMK51FN6WTdjfUy4vty0uAUpucot
vQZd+msB4bDliSax5yF7IP06vk9yozv8f1mUSkl7HIjrbw6sv80jMPdOPM6FQPL6
kgZfU7Nxn+F0vYyYGQhmhN7w47pCYM+3yYxnPhP92k/VSKJnWFzfs4x3PmYKNBP4
5gfO7FXeffrH0Z92npa/5hi9pInFwy5pfOiyWX+VsKr+Ztw5BcANV+jzyBiOPnC7
arOsJfzlCdxUMRXhxnzxPc1raUyqJd+lfl2lfZWEEDLwiwxLM2zWyYhqp5Mr5mdJ
0GOfrJ8FwPu3AOScg6sU+0hk7I0GQWlTmI6wjhH6NdPmOHYxK+lHLTcvNagxrWHe
NczylUUlw0FaI0BYoeNFtEWHvvA46JxxJVCVxVtaTPVGMUYaSpx0WntgPbGEgRFe
QLutUTycRnVeft/yv3XV4mU4jB6IWFCf+xLWgsdb8lAdZvr1ojx3k9c76Wm1ZgJA
l0h+XBYFvGeLCFd66JeXH2CdHDeSikmbachCW9W8F9p8KpwfyBKfARiKORIxnpHx
Urkjlv16kU+KwJtVtuWwLA==
`protect END_PROTECTED
