`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tWDKzDnn6la4SHC25Kq7vy8k3QKsFVhlcSAjuQtgUjMiTJfyxKrx+O166zU1xTxx
WYJzlZLutTVnw8FdFmeeyqSqa6Bxd4+xJXPQr6gh9B4l3nDl0E2AOPVyhOWwWKys
8ylQDF8v1eHxYKqGGWpa+GW4HAQnb+ZX2B7R+pdJkI7ugALfWf4ZX1KDVvVHoJFG
8UuhQk8Oc4IWZQoICCAfFGniyN0VLDNB3+Yvu0y/5HlZqgQFNM/HA2nqj/4Hqw92
JF/2F5t+syXejM/uKyb4GmAe3Dra530zahPHGMkM4ryESsIxXudsKZTIpqZQfRQM
F+kByJYDgV+0HwqARSR36946F1xoIJT2AZLiL9LX1c95dDH44LCg8IUrZtOBcWdW
bisWFpmMbEkIVhBPjL3LRSJRKNtKVzlP+Bh6dzpIXDoHzWNOqDnS72ooN5nivEGB
soYaOIOAVGz2oV8OLOzFzB2IP1nKwksMPl3od7I9PS3Fom02wPZQPdZ49wJ5Q92F
+jAnA/9d6cIS6R+IoSWvUFeQ57vorKpQh2VguXd4SwTBEfKnaD2cjfrt2Ys938gI
mer4kFMuknY8EELPef9T5izL0lgYAsFm7OG1EfVXWts=
`protect END_PROTECTED
