`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2JmwpbTr4Z32mTReBNVvFjNeheNqDZPr5bWsqENq+oikWwCh98sra1VmuIHYDkY
HBAW0YXTHmOSbqEhYiLKZPQ3i7Akpo+VnzMNFjsgQoiYOaJ/Om95ytpXB6oo/Zzx
OW95XWJykkjIy3zrX8OnYYot/w+ayPEtW2IduCp2pofkQ7qP+uklvzCfctO/hygR
ZPOOZAxU9FnJxGw1QAr+pGMI3iK5jdGEKTs5MsRp+RFrh6ym/0vDVK2xBTSdw4vE
Ykz3/9tkebljwyUrb5x5Vf67bEoGIKbvrH1dC47qAtg=
`protect END_PROTECTED
