`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ADwjD8cO7JW87nhlfHzQ+uf0I1PQTNow2t/cDz/EoHfYLL06+wRqV0u6tU7D6GFo
8c0O6jLcSMaIoNpvRqd7r5BFZKEhBvKxU2/xIDOk/yfKChnb+xwC++YnAZbrDLY3
jwTTyLgeNAh82ZjdlErJs/Rh1WWYzb8Yvj6gD0PhBrlf/9SeZLgZx/Vi1tazXjzq
NGT/+TeGuZSpbyPSGDGCevGCQ/s0034JdeSX8nSlQbtyHg0oXREwzS0S3IxHewrK
dXK9wjVlrR7no5/Dh2exBQ==
`protect END_PROTECTED
