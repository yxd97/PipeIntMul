`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uI2IIRymn0u1zppa5d1Oe0K/1VC+viaGvRZ7qAffDjTmAduaOtMvWjseDjulJTOr
az5bVDSWG15YixuFwKdcR6UtVYY3iiGspYe1okPV3BN39PNh5QX8tY/zy/nhjeOj
XUcG8DRMH5yCVnHAR23s8zvoukOPvsttAymbwRuylcwIUHGPBwygQcuGjjMW2CtU
l3AGAxwfOYqkB+FBllgeaJEM1xc2GO/nZScYqo6U7ix8hOqZYa2uhp8br0P0DUzZ
MiXkPbr9UAIiuKBSo8+nSKetsiXgGiM1Gbp3iEUMZOZg4ivpZe4Z+Xl4EhsjbjIi
tL+MkdX/IWyp4xLYENmq9DkmH7LgzdmzUj/DmeBcrSd0NdLQGaBDetT/7ABPhvDh
xcTgVE8PhXRArYn59wfL3D1TNd/IUMKhqVsXg9ifFsU+UV9n4QP5AikMa5wbUE5G
pLvKSkMkgkPOZlOAMUzotZ4WJ0+VbuxoSaTuybPfkcrrnIYbhb3OIeXjk+b4KWow
RYOAJw218bknLjcg1Kj0hHKeQJQsgBOS0raevzbPfkGUFni+zacAYWUhVAEKICEv
hj1FXMVDChkRVQybNOxR2RogaFcPSW71eoSO83WYeFKI8TC+oGoN/Y4vHm9Xwj1g
cLDRQlp4m0hEC9j0yld2Mkxd15AaMYU3te2NuqdwifJgBGbN4HPAqFP5PolcDjj4
CkqyG9Xxs0SnAYzz8hqu6b1y1JaZcya+g/tGXyaVsNFRjN22xmacJ5kQ2f3WQCaD
A9lBh5S6/aMDAkjqPX2MlOJcc4P8x5mMdG+6Kyeh4mvL30l5iLR4yiHwnAUOm/Yq
pPeBtA/6DZt0mXzlkJLQ+AbTibHgsPpjEWubKDVocW/Mvpi5L774jTV010qFdeJY
1VKE8GA9Yhi1Q6We7oez2mHuBvBiU43ZhaVhIoqUM4Z49dxm34oJgBz4QoWjzNpm
/JjiYmfFML4HA18OKoDysyCdD3o4eDySrb9BwqJ8tBkJpGraYfSAKe33Cq7sPxJ5
UvdaW+DFGYagW/7TvJqZMnYVCIB5lbf0v1YjlL8eEvD/WSM66TuM8i8xKy3csw1q
Mg7es0LUcyeGplOgLhS8ZQ==
`protect END_PROTECTED
