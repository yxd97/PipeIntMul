`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9zJoAfLs7iDAOro9WR62hYDWqm77rKhBV6kf5zmCc8/uL4DWt3z6vDneCLls+jDY
/g8TX7zK2RcXoaHlMTEAI/bon7Qr2QJWsdJBzF3iedBuQdT5bpxYahulohhPpc3K
OYbEhihGs0aSE/uzktdel9xlLEnidos5xb9fRAIw0Jb7JAfnVjyfU0wx2i3gvnQZ
5Tz+vDA3DsVPRbC44R2x8e7I8Nce8HZwIvKPoR4S6t1X2RBKyQZ+cRVdfpr/rJpA
HowJHRYxNy99lc4p2LkULB7C0w9FLiUNONZo9pks5mZYPAFkxJg8XS1JnfQLs3cj
GC9L0GbooduzWIj6rBoeRGqI4Qv44PhyJld9/kW+JcsqUJKyVEYbM1Crm5IxS8SF
/B2EjyXcmWXOzllvG3v74Q==
`protect END_PROTECTED
