`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AwBtnbmSfCpxKxI/aCY2PQ6ToqacpwkX0Dj9nHGGgaVNRr/erPln1dwagLJBU1Qk
vDG4+q+9+tixM1Dm0tiBw4wVHzfKhzHimMui/oRBr/K2H/Vhye5cqj3xEzQdxVf8
WL3Kr2YsBZVOXbp72bojWcvyVXTNdBcuM/MRcGM46cXiFio/IlsjLvObo3bbGm8K
t4LiPCLychbwdbg83zzfoclWTszIPO5o5qRnyIa3Cw+OhH7qP/J3DEXK92upgdZI
IiMXb91GtWK4xiNZ2lpN9YY0nuJWD0YsZ5n8bdY0Growe9vXkdWqC7QkcePSaDq1
+zpDJ4yal4h1ZfzFjbg+VG8Mh/nwQpbRFh550Gt9Vx5aRZgiG/32d6hYlEqNIKNY
ChDNqBpPgk9Knc+DAnQN6Sop3bRR7nvR3WUfd2st1YsVpsMdzrW20BGT5VkFQq4t
JlSDoqA6GnzCM6sb8CwX2hCfqqhscVPgCh/QLbtvdTe2lBOEB5ziuZgpW/O15UhL
gk3uyot4m5jVVcGkWxSClmN28CUp7NODbpFuCs5IlXuQMG3a12/MC6Z9foQrrzhs
UVdTFqflAS/YE/hQuLEVQEMfCWkz3qZSBXa5wGxWaczjW9FG8fe6shXZlGIdwFPJ
ksExy0NljoB9LH9N4BBtHA==
`protect END_PROTECTED
