`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fGjCdmWss8DFy3X1A6dmBk7RAIYDTsQg79FMJdxUl5NErCyPAWZiCP3ZWOtzW0WN
7WlyCUcJDXZZ03Yvg1/I9JAcRN7ysJS7PEab9p/B2G4LGS0eTUrRJQ4NxTr6JMJ0
Sk2/mMaqeEvV4mJ1M2wMwbs4R2zMlqypXR3hKR5MkTVnSupfRF3O/zOajYrEeEv/
2oB3yGAHQm5FoyCCasKNYZo8744cjNBjsA5p+0Xpz0PMdZtGkxdgWdMkNBR01VVF
mMO9Kb7Rxy9Cl8ahPiXe/CFICpwTzVU8E8dQ7xUK3YTeqNckrvGX1iPVlKcVSjIi
tR0WsmILk8xClylF7mphTIiEAzNeFXfG6VQseIcuGG6TpH+juzTbtaY9AxIozFXR
FWbumnmEDZzm8W08HuRQwDPq8OlbC+r1l8I9udzunZc=
`protect END_PROTECTED
