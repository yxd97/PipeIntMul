`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJywewE0gdgPwVH+BjejLQfgMg1jxImIpSCzJr8tLO5m/fhTgailXmwxTlzPYWTf
piLf7AxlBcUwXbYRWcJv/sVAxkYq3c/2vonCHdaRiktRlWv4JJkX2GDJcuC4bQUs
xrQa7I4E4Wt/QIs2WpVtrAEwMQrQnZtFnlDTFeXLyxGtq7zNyTsyQz9VqoGP7x8g
6XoLl5aqjlnVzKjIB5KQBbDSdLL+luyqAJgBqO4LXOoJCPX3HDIF7Ov9remS1Z+J
dJmmeUEjvxGC+JxFMwEUbWnTDKUAtS0RyxqlFzkOabGgLqW8Tjt0i8bt3c9ks9Yt
82Q1yuL9U76Cb6dXoWkPgpK5aWZtyNg1ccvjru63rKjQB/IH6PwaVfj+bZf3y8pK
s42yXw5Syz95GNK/eheSzYNTI2jBtxQe6DvSALYmMpTccvg0erTHWOeRCvoUDlyj
2x1YP6FvKZ5Tjv+C5TSCTu96A5QhYBwhJ/qRo9ZMO/Fjy+hzc96TQLc71rgb3MY2
VvpUa9F5Y/Yt88ZL8+6cqaT/BAx5qXtQYKJz/Pm4pQ79vuVQjSIpCMraV6tOdrWN
0YIX1N7nuRuFj415/O8LOFTMujafypyDk6W48tqinBgbftfXvbnb6v3hEWP2LRrD
v5ejQ7bdgh81vEwUcZZwXxU3TxqgAwAIU57+gKwnLUJWt6EDrzU6CAFFEHdAzVcT
3p6k0NV6SKbnWoBHVO9y5DlljvtDOylI4lf0egtYc7qQyCJftVayo74g/VqhTDTl
fGQiKETXYYxOC585mec44p4XcgInRrduXpWwT96PCZ50iqGNf3taQ2gMcSwrby2f
NnybIp2Cr1KbGdbi2DxdaJUciuwoczICXhhJtw/jPRpuagod18uWwyRZTAv17CF6
CP7RsXKjVzdSx6qohLOE3uPSfKVIViotc3EM0h6EXhE6w9/aNETkipEwuT/SYUn9
xRAmKFRGESYvndeWiN/bJFVwu2KMv1F+XW+CryQVUAdLBhKejgIaz3xt715jxkXC
albGT7t7jzlt98iHk2STMh6OCL5SidfWpS2cp6SprU+ahx3QJFNf6dqFv2Zb7XAE
STSUvs/qF6tNUr3PJZK7VdgocVfxadX0YFEKc+F1p81MzKaoyD17gxBjhavbjPDJ
i1EDYB2Dd8TGTYMBaz+6jJ/yEzbDcO0mR0wtuhqF15kHCEzXQ8jZHFBdFIMuEfG3
+zMZVmwwLbii0MHfRW98JSF4LEAearZYsNxuRLG9hNCP4SM87AMBRcv7SBXaHyjl
sntf7mqXzqnrjz3Yx9txHG6F+F0K8ZtL9adUGNP54BZi24qLJHK0BnLx1QCruj5Q
OZGzkNoS1SRXjs+hLNbpq0iZKBe48PGS+Lecn5V+ON7qMiGYGU239Mq16b9RZnew
a2EEZbTZLsc4od82A9szl41NGwTxVByH0Sc9+LJmIoTuK/1rUfzyRqZkYpZrNU6R
riS7AKFtGrfnhXEZiACXU87XGbRyCIAfb4lA81/tB5dIGLLTRIaMSDHlmdFUPGPy
g8kWHeDC1jaUM0zOEQWMrmcmR9ggIQEAGcpLaLcuAYVrBmp280VdkGXO3oN19AVh
CfDEUyXRCvRBVo9NkpCM+Vaay7pTVOHseusZHNoiogB1KkMrvIrIhzWBZdsUxVmx
zv7egAOBYqOMKxS9GBpKo1rNXQo7buNwEhABdIP8FRjKO9m7Lkrw4yb7dT+xQ004
vLT8KfmPfbsxqsFIiJTYcm0xtgfP8C2Rw9BhueuiQYU1aoQqZd9hXwgXIF+Qe/6R
v3GSN0pOY2uUeDgn3bzp8OlCYy3p3jKdBtoJjopjy2c/nPk7JxkYtgaYHoYEmkBP
vwO/Hq2OsZWgIKetelcJ5+ojN3dmBbJSyv5ExIGitiO8FAOFxID1+s7PlQV7EvpV
Bjmk/2mFLQhkxaAoI8RgqrFFpQhGtdP3f8HPv+r9DhftVLqRp6K8cGTf8QEaJb3D
vFRGPCK94KZKVAknEkKAk3Fk9/q6x7kVHuIkP+zsxqUmpgnH0ppZMhoCxLukVxSG
9TBpHlytG+39L6h7x3V7ICpYZ13S2OTgStNHvdB2EgCKkqm4BCg0kVJEd8bvn66Y
EJimDmN/GzW/AByavIlmy8Fd8pzDU4cC+nkPKT8wyuyPM+LkZaFoDH5beNZoyVyu
LPMf1/dIdLoWakxybN1lrKtZTcAuwFV5rrhqFoGhh7FdWJMnrxKQyFfEBGi4CbK4
aw4RP6JHyChvE0kuGSyNoEpqUXD42pB1CQGEqWLdGYa80X2WG43gqVoXMK92LWFc
xkM2NvfP6AAvTVvBJc6l6v5Un9hQjpBFO93EvZlo5P8=
`protect END_PROTECTED
