`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N0M4EoMy7CaOmeMraBHGySNZykQwzTCruKuisjARfpMpn63FDPfQyyMWqxsyrh/8
2QDX18NhR7mzV2QP15lDnFIj1YSjKxUIw+5zbLjsJX16Lb1snjOkO69hqf0E/oW7
fb8AxfiGGnY/ThKACzOBGW48P/LhVEjDhtYWGSxtxSZxbplGW3Iu5ZYcsLWBcDKT
NI7jFkshehEngqEEx1xOCA4+VD8kfNSjo7mxeg4M0UbJWjY08K6u3ICFybUukvbL
96kvTQdk6DS+vv5mIF2+FQRiF9n36KgQZsNtgiTdzVETYlASCAxIwRKZwk0LmL5O
7OlUwLvcwHnh+KQOeYRm6WJ4a2tNulIZOQr/+lxQI7R+28qI5zzNd9+Z5VYPHBkQ
`protect END_PROTECTED
