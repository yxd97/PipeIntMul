`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TWRFtIx85Bcb5Fap55iPFh9F4LxkDNybNu4Di+y8PnfX1hfHY8AEK0UA88IxSpVG
wNfE5pOJwNNMtkv4sDlzhl9hd1pDHd6KrzvLULBxbNu14v1EKV2kZ9mifS3hiOdo
N7xqiWr5YkbCKz6gQsgI3pIEZFrEpL7F3/jdBPwCBwILSU07geOa+yg+oz/WpNoR
AbUMwHRStsjQLpvZbuyvQQsREPxxuTEyKd16qUYQkuVOiLAbC4mGLTx4JfG70XXG
mWg9qe0Ea4Pw9sBGpjA0NAKRD9iRtrujlLW3s1xYfW4IBrHU8Dbt0hTKPpFSSNWl
`protect END_PROTECTED
