`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kx8YMGzclPC8t3LKlLuXUJmV7SsUjNqZR+L1sjCLCW5YKNc5rNlbDNtljXAU3S9h
IahooymH6sWkBPZmRk1s+8FlEsFUsU6qx1btcNd3UZtXrlOL5h9Gn+NdVcDxq+C1
KzgwwSvvG0PM8MpoXLMYSo8B12OManxuC3EuUlJ/f8gAza2uSc8dJukYOZE9UrJo
ig33bfPfqARrOxeXErNz1ULS79VgJmUPSCuxUOgKaVqLqu9O4HfEBs0M9doQEoPS
bWouC3vzDFbugckevE+lbMGX125crjWSZgMEDdGvEz7RH/PZyFEQph3s3sw6gCBp
1RTP+Ip48kFouuTRsoHerSuYEGGyLv/sDsCOwXRD947rj+LtZ797FFxK/cuoLQJj
mepAcG7TA/mhRA82XzELfw==
`protect END_PROTECTED
