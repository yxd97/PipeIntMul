`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kOgQh37lGfkh7Gaa/d2sQwsxDZ8J/a7lk4AMYe5+7in5uG2KhBUC8YJczLXW5nS
Ylgxe2ZU1nqD5L4MHHDdPnMHRN0tUl9+ueCbgqtp/SWcClxDT3fRArNp2x0kLIPP
RFmseL/g9ysjLxxpn5EW0k4T62+rq9QLacwAloCHwQsqMHgfZ12WHc4/UWRz3M7K
iFHTeVjFn8q60BezauEfHXx9jyo2Ske6CeW4xWcblJNzGgQIkNYAICFsHTqEoFdb
OyCtfDq+hx3UuuKw8+LKHRm2xX6Qrr+aqtFdIszwnauuQnQlgJe80Abu31562aAq
kCCJgviH0RksVmrU1jCm7bBPVSlEcAqG7yn0nEWTLF9LIloHUkihiMVopjzkbHya
b8ehxwb0ZElGm8LhTelXcIZjwoP1R/XeCc0bw+/ZErY=
`protect END_PROTECTED
