`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pIiIEgDeDjHLWNSsM/2D+uVKT/jrFIcVpZbWffDN1uitgo7E7rrqLVnIzQvGYuLE
/iUOQTII0PZCAK8my3b31VeoVaPmFwC+XnLGAMDWcQO4WG0pclZfP81xs2A6Bd70
7Tgop/jSWIi4vW71qzgU+hCRKqD7irIvRkyQpH7IjMZXHHylxF0A52WyDzX8e9i9
J4HO+Rvna4CHr2peuN3k6mzxGjVS2SQSM9k9w6zI7l3OPre8PaRYY87hhTANGFVP
2d4AVEMpPN9TyqfCrCG7qd8iB4s9ubLaKtPtC8m3ujEM9aiipNs2n9bF7WbVdIhu
gucZW2z10aJG38dCBT13S7RRA4/8Zn+xFglXiGOL1y9BDq+VeXAgU8VSmk6hC0DP
6xtCqSx6ihkO/1mR4ISHMp2+ScYQLuyY83gKOWcjg/yaFoi2HFcQTUJDV6yeyHEh
t2zj619jf1sDzEqPmdQnZ1C86t4OuFf4cwqg/vAJa2NVQ2uv8oAnPuwvcVwr6p0a
//EBWHXeEronQ694DpCLS8TrpBRTpOHVK1xT/Qdr5+um2LQxFcdg5z+WXlZ9flwx
ouIAtiO5JQA1Ec8YrVwKKw==
`protect END_PROTECTED
