`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hyy2/x+RJRVkVhmG7mU+VjbCGTPFQETvflUUvXSkRVN9Z75dH/DHK25IsHb6OA4k
tFaygzcQajywEOZfVcO/9i6xWp1dtoRT+EiSNFGiJkDnpdrDCIBtpP9Lc1ws8q5i
/PLlPTqzCYiuklBFy65OSlB7na/T5IbENoZntvh9yARhGct4GpTg2L+pS7i+DQSd
Qz2l54dbNAYYp9oTk7c5iZhHov1q3L4QpdE63IJ7eWUexkEXYyZRrDG36aSuACQ6
BZoCNhVp834t9NlFXJpH2E2WDnZn4YqVDjnT0vvj2e29gGBnBoNXKI00oC8UH21+
L46BXbszbGfWYDJWjExy3DevibNS9g+gVxLucL9OH//S06cMuGrWyoQ3wmvLx7YJ
F5+JDRBGYMFcKKLzbTGT03ov+uwfQuQmMVB2+gJI2V0NAb6rtcTTrCVnhNW7ATK1
4A1HnLdLBNPOKUSE0UFbs4BdOMWnSD/SPGWd06fHZf+74jyHFW/QX1kvZjyO2ARA
n47xx5dita9+mkhUawnEqkXQXJys16XXwQfePde+l0rZjRPJD4NA5CbS8exMnWrI
5gRp8g7jm5I0WZ9+c89f4gnyQ/fP8Ar9RRHYr/jTVPSqrMN9XWf9z07iWOrNQ7dX
ExVflyKNrhY6mPxjeHrhwQ==
`protect END_PROTECTED
