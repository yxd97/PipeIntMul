`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fh3WYPZDXXIcITQAk8VEo6dj4U6iUpnXgSvUTV+IgnKyUCt7hyqFGzG2BzsfUlxv
MDqz9TxKZpg5qrwqND0nOipnB5AAzl7EcRLUI9s+PBE3ZpP5C+5kPU1DAOXvfYTV
RSs16oW02VjUTh7HQ5A5iAe4dOLsiRDE3AQwzRFZvaA2HqXiJ0NKlg+TzUUu1YOU
mQ9SZp3XaHwbTSzj6pE11hYHLdooJihCFhaKxbWJy6g7kUuCR9W3InJEk8Yl/sGf
Xg+ZUxZdpkcHqsFbYR4FjOEv+yBFFVOovA0MLNU/RTwSik9xfzilnhs0SS4uYrIN
uVlZKmwIBd5P/HtWBUm9NNf5fNCbZ3wk3az09+8DzXu94R4U9hjynLqV2pzqrcwE
6BgfiHfbIAtpRk8549TtLNKjvsBLsB0tYg2MwXkg/8sPOLX2bM8dvH1Xj6O3sNKr
ldIoSE/YvhKz86qy/fekhcfr5vFlC3H/+Mxb1NKrF4QnpgKAq14Vckurc4iEx/MA
uvs02UJKBPh1CJLvSct8VdtQBVa7eULyZ8xzAdXprHm/CbSt0ANvCYyqaNMuaZYJ
U4gs3AboNUnq9Uene4cRHC039Wp/DMZBl+2/NKktt8isxg3H/29wyBSicHOQsBeY
qXkkg3PNXBmM5DN8JjVfAZGPocdF6HQIVrxDWzqIG3Glh5zZ7t9TVeD9Q6A5y77r
PhnWBWKQzkCSzSBQjkA0uwY+b/udayU7AHP831y259rgSppQprAppc3lRZU1l6hS
dtczlNaY+T19RlC2CEOwAE0Pw1vaVyrOZyqRs+bRbdiMdqcjD9ZwpWL9Mf8KSupU
nKLik3eoMzQYKYhCgcSIg2mAZRnsQPB9t4Y/SX8PchcI0JqJPzSuRLyIY1/k7Egp
KAiwNlAVU9bHQJ3ImOBmb/xHM1GOH2UW6FrLAHQvO7DTLDCuH1F3XTPlgUJCaWuf
4dbNpyyMFNXoVYkIzSPSKpCbbotBZGCKuYp0/KV9a3DkT4nyFye6yz7HAgV9RDNW
GY3LAck2/DcVDqxaE7G8KdswXy2oHBduJHMuKIj7EtMtr1HLtwDvPRbLpIr6JJu7
l6vsjcvCLgSr3kr1VqwR7a1jboW98Yd5PmI8ZMSn11TnmP4pekCymelvBnIvZpd3
9QbgMsvpFBLNdTwKMtpxod7Hm3pjXWodNsiWmFYJhcTAJYKrW6Rc5GzWQkCQT6jy
twjtekTT4HNoMdcdJdSBgfbxEgGjv8ze3Qn4AFR0P+XzSs7/zjlqLi20waOvD9nH
cAlZD2qcjjisreflqG7VoNznzOHHSguqKy7y1LxnOdJpPablnQqgqEj4u9ITLZQL
l4J30GHXnLGyM7aOjOMmlj8gVc15tcwUVefvdqnNiRcs8IQCs9psMIAJNcnnSrl+
D4ZISmJdT3J/Cu2sAUo78R7wkXYN3stMIuZkBBu/wjeVVZbI+HnNwT4vbcSXXwsb
KSOiU61a27ks/4KndpwpLoAw6239bbkYm0Z+rAHEMDi9uzysR4P90tVd3kjRmuuU
JT3PYdqPo5UmI447DBtBrgVPpQ95jJU3mIJzXWbAo8u4c8NDRYb3SR/xBJgaLjOz
xzn+nwo3lEqssLGK6q5b0VarwfootDNBWBbqUaam/njT32kmTkSC0jyENvqpTou8
v8dBEpjNXfLbHGg56Q/ZHSQxPGLuZV/r+1iW5O2DD8ufUylVEOsZBtheOnF7eLPO
sabWhyaR4OZLB3HRa0GycYjkT6isrqnxTu/q+iJP12JlQPBA17igCWG8qnYJHEK0
OQVolffcLDyDafWrT0zm/vdx66ySFyh05/kAHF7oPGoqW4xAk3zRI3HUMkleKx9E
intzFe8Wg5zypdWp3CQUWy5NdLp9cgSMyDqHREqxJw2ZwPseYJ7z3iVtKpiArvrB
/yGTyXRn+D0FlQS6lITzH/fcvn2Yk3Gpuje71buEE/ezdecaz5MzX8WJyTNMnmTM
e/JyiBzZIh9sVHRzbehrzOrERohZ+pSX6uHOFgqO4boUi1ipkXWS8TuHbTrBtgSo
6vR7lWTyS696NHCTEDgLlcDYaeRC+aCNpUWYYTZjOdO3IXYl4Y6bxbrlzy3wS44o
+2UWCD/ZEIChSeFZ8N7rsOnavfn4sXfIs2M5uaRp8OCZHDMs3Vk+Dr3T9RmhZ09j
OEmkToOKsmbEQRULC1RefK11m/wHuv17UQ/OM2Vn+yZMogSSMDJnT9gZI+0QJF7o
j4EhLbP4HDvr+VTlgw5/WiXTDzW1v9H32tIeNQwUJjnWSUOvVGZAZKJWT3KZuj78
5COtMtpklpufxEz7uTtMxsYqKS1lLfRMdm1IqhsQOma7i70artZNP3XC3hXAjA6f
vRiI+RzhFXX6YVh6+YnerrH9agRALSQ4HNV+I90xc77ftsA0aXXKO7e6Do8JyVmO
BPibCtOnsZaCjdqY3JKV/Tk3EnMhs+QNwILw94J3ZC0DxVNWfvt3fuSTR+lUGhWu
Xmj5/rGhD58ZrG5R5JH1DsBpMaP7av+Sqy3cpkynwXl7ZiRy1ah4ggO0OoQu20O0
JdtDHpacHhAVIvJ/hUWT27QkK0bWyG8zNL7RTjkH13Fqa5ubFR81F+Fsnxfy8dAY
ZDtPI+3NOL71VZ2mWNHerftLBtY7VLa5diuS1L0WT+WsB+ovnhsQHm63PMLV3SSj
AhYmga4pjYuZ25fQG3esl2RsnKCaeiTYdHDsqmDIU0/XJoK+4RTPWHKlHy2aZf3p
Y4DkCN48/QEex+u5EJ/V8QdxYqsoRZi+HeeN7TORQ+yDyb+k8AenoeB2OI7NrYEH
bf5ZAfG61yfLtz9EzRzhYK57NTfYz4dnjkUbxF1Bb5nkxYOwFeDCAbzlfXkhgO9O
Td4hmlsgiKIKF4rjHAsqX6r+B0FbObRtuDk+4yW6PQlGXsfLU7Fb1W5shI6k1YzP
AmNFyMZ6LQQluFUfMzzZxvpfO20CaBSSFKw/IzkqwXQM+PMYkJbbgrrKxQx/sGxW
/JlBF4F4ibk/Rs6GUPEMLRiBdlMoLcPLkeSoHKSSGO1tpOtca1kMyVw89Avq5Qkb
4L6/lIx148k4PrN1mREF77KHlzu1uD2pnvKdvva6BuWM1vhFgfBHigXLUoFcDRp5
ZldcVHUYOG9AzbQMVz2WqmOyBCUNhvXijCU3NZfEn/mSkzGtMUpdS07vVC0e25c+
uWnW5cadyLfs3G05tIkFg173Z4GjKbXYhWKvjlL3cNvapGDHxRyLogF6wvcKwcx6
ceERkqI7Tt5zVKnkonXudZE39dT8ljYmK9S1p/V5hVkcHnlk5cU090onnN3ZLAmp
PiaKyZ6+0/lFmqU7Je7McLEu7vYYInZq22AMhHZvS7rSaoqMPtXFFwh1HKfUGHDF
fatj9O4All4n46XSmuOnYb/edP2VAKdZSRJUXIoCw02emos/TsS+ijQ8IewUlD6d
/NPn0/CpJiXyzls9KJba8U7UZsjSMec8jBkJUuG0cCyee394grzqGytqnlfdXH+O
e/sxyFtCRIo6DdiWuugpzjLrTG2wKLvv/JwnSesDkOtepULlhLT6RMkkE3w/vrNZ
dI5otFEmreEW5SNlfbFG7KsmPIik3ocs7zbIHiUH+AdBK+8rFMS4cZlVO0IjkZXx
ogtX9KkH7RzbwkouWpfmFlfnUivw0rR++bv5MS58Ivjopf3sKvbXzwJt3oz/9p54
KoQmJ6CrxS19A6I6SdImti4/opkoXv/LGxE+jpy5bkwv/1Wls+FbpH8IQesycaI6
5xVpvCyZEWATc/daqqlEWz3sn37jkwlKbuOuFVWiduKAw7yi6gvA3iCLsazf4BSR
zW0vzyBoKRB61xe2DZ+zb2fOjNyL2OJAZSSmNSzKFs6AqWReALywm2Kwp03KTHQG
noPJPvXzcrKnjFL0m3GZ+JkUnzvx/z95NNw/rSnGxJFtAmFwm8xfFTPAaedk5S7J
geZ0nzkIGMF2w4ALdxIOBc6pahJC+vaYjvxAwShHV7cUmTT2dCRAez6xubY0tHvF
D6jNaDOu/ypKyalacZAOf+156Rkj8/pqJfb+7I2S4RW4VKjbsNuUF/H+FDCDXXj+
GAR73210SEfRbsAH5hAIxxLztiugCnFcPnCsB23TAvKsY1XBZOoeLbchgSGGF2ll
TRLGB0GqD3xda/VmYrEx+U2VddLbxboIqu3dcnm/KKpKu8Awu7eFR88vy5BKq6wk
a5J6PfkQgVYx6CL8QoAJylGG7WdW6se1DqlN9HTSyAy/zuKIOxgpu3VUP8wa9bNp
5EmgVa6aH3TClkGFrUPjNnaNhKNwpni6hsvmMezTPgBh1IxGq+9dP4nwGZla0yi1
n3TyN/tLZUdPoCBd1L4xFjzAFhu5urSODHrDoHBqHQgpqwyVy/rV0Yl+ZVFho4j+
QTA+/smNnEqUBNwpCmFlXnoB4Bguc1+3faIb8T1GBR4wnQH+mpvgrivQxDrGuHQS
V6r6VnkiJXUPszYVfwC/rnOF58H+T6lL6lML6ZIY0p6T3/dgpRzabW/cnj9824MB
3KFWAqfFQAM7rXeYJjU6j1W/hHYR5CiL4rbz4E1QX66NqqYY7CP7L/4aEs/mpu90
tLcFs5kCxlclqItfMCwFudLGm5nkSWa0n+wyFc0Rjn343yRp3zUKD8usg6W3Kqen
agh/yuOksQmSUWODEnhwLg==
`protect END_PROTECTED
