`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yL1D2WuzvIGSR5DsCdsiR7Y56/EugGzo1wXY4Hsl3lm9NBLeLcAjJZHy/HTdeu8s
dV/ujdIraQZmdU4Yfgt5RaObq+1zlzxfOK3Z7egh/seDCuQevfRe6Nz8nm8OmzCd
A1kgNvRe2/7wWgWupH/PMs7Vl7KHuIDbwlzziRCkK8h6DdgoXJ+CLQR++zjz/ybp
1blqNIws00winq9nyHUm70pYXkXD5JjsbxoRv3xqhst9AK2clq4ShqAzpOagvDvC
EhqTapDyzRuGtF42GU0bgz8i18DCEMD1Ha5gJrVmk+UTgiDuT3yKB5uIzMv6qjM7
0mDATbpcwAYCXPmLEbto9rilQl+d44o5ZKSh9vvO89xGQCCpEhi8j/2r4TsrBEXi
o24J31ULY52zy5ieXhF+IoXU7Tr1owY7unFkv0jEefI=
`protect END_PROTECTED
