`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2XB8S9vxSMchQEi5DHwH3gUlzPTa0r2MogcFSEGr7WPQwySrxJS+irC7FJDdtcS
LX+XeyV7ngOkGtwvi6+/TEXC0ToUNHFUWnuyx/c1J1RBjrO+ZVvyDP4ypz6TyBFz
0/qoSV0uCQAts549BLCn2HvJs6Awj1VDbHxtItwwb10+tDK1HcodAV8YAsM46IrR
O/ItyXXovXrC6a8u39rL7TVRu79d3zoptnIiIg6A565B+rkCq8qGbdtJyZrH61Ed
5PkOoHMh6hZPJTc+1HKQUcXe9kH8kKm3i9RO6YgS6VL+YCUVvVHHBVqA6jFDUakX
jF4Dic7QJEu0Bx6Be1V+chZnAUKEOtzfbn9gSjEWPyDJU0a3A/9hEaJdDqkOUvNQ
lmWFs8nH/JDEc89nuv2RA7eXM8CGkFyLjtEo3XBIIB+/Y1Rn5OBOnh9SqjDvPTgv
V+xHmes8Cl4jqRXPXz2JHhVkRrZP3GGmEZFNOHrNl3U3cW+Tz73Ax+2kX8PeQ3Vv
wfndUn5NGS/08YjyQf1w7u6Vpj1iEBXFEXI328yuL185ttaQEICbDh58v1LmQLZp
u8Adi90s1snDxuDDuTX5yA==
`protect END_PROTECTED
