`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N33VkOiGe/F9pJA5oiYVh/JoZg8qXwPygWZYAn4pEUkamJ6nq6JcAOqP/x31ovMX
bwg44fVCJm3DeV9wBXRpvj7bqhUIZaJzSNw0ODhGQhkz2Y8Ki/KlS4/U9fztMxOU
ljOfhgMFbU9N/sEnUFHb4jYEKVKclT10dndtMbyea0edg+Ka7npi1XOGBinZKYW+
RXncC3vEdNNpxU2Q2gJvIR7MPxamTbZp1d8Xj5BySxChJrByjYXf0M4wmKgRCOML
QHe/2WG/gV+0IaomymV6IZguFL1Hjn8XAar16RM+sHEDb26yiljF2DHjdvHU2emj
1WbrqMO6V1A83nMBqF68pl7prXmghwr54w8J0AXmW//s8GzNb3HpBroUs1maLRdb
4Xje898H4R/v4Pw38/E4/LwVSzCD6ATRnKR8coA+FC7cPX1DKEaecNhig4+f4Tei
QmSHl6El2aAJhkay6N1T8UglIFrv9AkUu6aoKhWtvwpR85dZ15K/n5QHNOwZkM1R
kOkj/zvg+8m6LnuATs1Y57Nsz09MzhmrBV4uU+VdblASwFa6a6YXcjFv9JJ+wNeO
xTcUgzBFZpXssDhUxbZ9PqVYwuZtgyYejjUBrREu1MLfF5NgacKsDTt8GMRqpsEP
RVDDvaSCgiA5XMcPWVK0MJK3n+i9jvnp7PiOSBvenGftY9Bc5QHlvCm4+/ufodiQ
qeHiKt56G8Qphc/pP3NCinEz/cwWwBhSnrzb2VRQvXuNKLttKTLl/H4g8OmOAsWr
ZIHskqGxKex1VIaRMvcphyHkxL9I3NfItP7fqVvsqW+qaJEPf4AD5NHSEpcSNfyY
yE6Ld79ATx2jpxi6OoX+EvDQql1kxN+9bQwQTN8H3My5JxNnRGTLptbR4oLcdbh8
dR5ZeYVpPx3CH9xfSwNs0c4Bhc7VNwRHuLhlmC7OF9nVIhJntxeIQOtGbcCxM/Ou
hW7SdyzzZvgrFzm3Z55yDQ==
`protect END_PROTECTED
