`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U2FiqbSWoKIZ0Nsuvh804ay4kHhQpMHsU5vndXUVaCPxRwAlsVhwFSJrvElDd8aZ
5BM5VWGKCMGdFO4ATUhXWPlTQYYnC3r5Xtgwt0XmMOxeBapyso2BWC3EQzVGuWMf
pmF9S+mxg/VYaoPRE3//PivFuHBH8/Y5XKhGGf3oeJ3JPnqFyUV3mqXCTrcozzJ7
FTXXHxeXmfYnT9pVnu/1fM9VU67kOo4YiBWUi34BaQ/ItGMN3gkZKCzL6ooQ6VTk
f4qOp5UBTvAMa0U0vYI0IQLLEqLQih9CPnDpvxhO7HimYlax6VswZVxT5bRtd8P8
Orn4w50jy7mHt8R1rR1Cd5G1K5UascVMjrCbu5RYkUjuEEdEqVO20AULtZpDAVen
fInfLnKjDm9EJW0MFlTWKShB/CeEWp3fYUtwFdkX6pyQeT033UlGjFyw98l4nKxC
WI/xjXtcnQC9/tNXuT5VFgIyvHqgmMY2XdCj7uMzR7U=
`protect END_PROTECTED
