`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7DWeAyQ5dLgNpDm+QztilF18xCpnzXeNiL9Lx3IX8tQPgCYPiqI2W+YP+fXNRuD
vpOxXaMzw64xKV9YH7Pwl6YC20WpmQ7UxPb4qxUcg2QfGuoa2nkuJJEugCyZerQJ
WrJwTYClq9x1KzpLq04GiVAr6lsLvApZjf5nzUcymLab3SVduHdd5IxF5pe8xRil
48jyIbHBfzci7OXOgdIE4Qhhx/qtQiEUtSxeIfNSWMjvWKtK0UhjEMnb+oaPy6DF
TaIuE49m6kIIVSMDWYcMRnoSpELGZLvJje+j1EYLG3WuEjVrRqL8Vd5u1UWUzWDy
Zji/xePVH548zvXhTU+AGr6SdsXG5HMUi8rUajr6CC3ci45Fmx/jPK6gEGNSLnAs
vtbgHD83U/JfnL7fO/ZdUZGHB9DAogEIoKQjaTHqUjFiIi7Ru4I/Fj16Yx2c6cf7
6PnSReoBxIc00qLHY433RA==
`protect END_PROTECTED
