`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tfhyh/5Hi3uq0lLLp9zyNF4YjVjKNHEILmSaqwTgEAPVF63ja4Ph8q0vIbzPWUwl
vn+vhSBoYo8/13VScht0EPo42tldDVtvlhwB9Dhx1GdSo2i1Ejm7PILTWxf1RDZk
xxkTy5LBjPSEN0s1hOYLN8gPo1eEyAMmJ1dmumA3XK+iPBxqmURW5FfYMlwhqQlb
6bi8ew21WVGbUVCO7/MkPrsPPkhHPT+z00cQpmc6kFsRffV8tf2zG7XLMWBksvFQ
US5a3bHwV9zhrXrthq6Wvj1O0BHBhvq61ES6+LZIJlJd0TrtqUn32zh+hr9vwoNa
dnmAFe4lVwytdwFr/t5N9fLa5FmazibdsHCRK0zM7V++daTW6wSAt61soDYvride
xqC0IXnzW1ihEJD4aeuYz8wz1zH2m8Iwmw2+O52moGCZ5TrkyKyzJpL62iWvOugM
2pRLduzbCPnv3WZxSsEl8aYxBtaLCxp9Pg8GnM5GgugHhXbp/CkRaVIPiXu+f8Xb
Kr6ch3al9mVqnfEkztmAQTxWVcn4ennXeAkiRaq8fAM=
`protect END_PROTECTED
