`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ITiWx0RE5iXQvUzhR/BhQsZlFb2G9bi3UF4fVGOLklLNmGbMEirgBa9VoKulf+w2
aF+VeSU74v70TyDdMhhShC44vs4sxFNjqkIFABofnMcMss41DafMsd+Ibr9h6Vr3
JehpRxYD8ye5qCiygLED3lQIogfC6+acZD0oUsHefOpOWiqBWLgcmSsxu7abT7Sl
jdSpjM68uCDHWejoZ3+Zyt5LJbDvcG4tvysEgMqsVzYFhx36w7kQaBnE5JSifzYg
9KcAY0tFgRyIFqoaqJERubO1uTEaXhi0zyr1087zpbP9pZSfPiBcmDZ5imAWbj5J
vC6HcMLPfmGkIRI3i7//hB2qMvpQ3Jb2eUhLagOQSngC+BBaEL49uEcptZsW061v
YM2XhOc6ndfbytagswUF7FyPFFsSjmjzzNIQtce2eaV7Ud52cAm7i3WUFy9DadCh
xeQkaU+Cl0/TBNwNsEn7SUm0HicFLOtRJP5uoCMLDUmAqLnI9JrZ3so0mLySbCUg
fQwQv3rzoODDLZTUmprgkXMN9vWxQ5OjQLlLERJJFSH/pFA6KPxuD+rGhJm2LlX6
X52+rTxwxiYQ8rDrWHWUP0z6pF6u4Y41Wyy6HE4vrTC3tsn5HDVbanWNz7beBo45
XwxBQN/sGGNkzm95KxTh+1EYlyfXxuyJOT0/afbZRvfRIloCc0R6wWmqO8Hqe2Jh
rgqR22xEwErzCxAQscezbe/n7VVlA2S7XR+M1T1h2SjDDSAOIyIJJAcLO1yiD3Mi
Av5HVNIuLMAgSlu6Vus/4ld6TGKDUpVKjA/K9Yqu/ly/Fh3FSC2LMBSYYDswzkdE
EoYL6d5AwVjk+deZiHLLSinMurPfvJdlbHIs9aB+KnCV7s2IC/T+bTJTwHXA1H6O
CiI8dfYwnnbMRjGid2jHwvieSpHIXjEpUkWm0s1TWSc5X3pO729IakQCl1DSJehL
ygxh2ybaRBNKF5RCNoC3goni289YvWZGWPaw9sOC5oyBAffL/e0gQeg1rkZSDxIv
`protect END_PROTECTED
