`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2gIB88sWtMvXXhDrioBBaZ97cZmlOsDe5dzrC9emsVBGZBY1NR2ChISMBMTpl6EW
8muzRNTJDAAXbXpbnkvWWbmA3f9E/fxrFCJlPhCvszlCRxcVKESks+56MZmIyGGc
X6WS2+Ymz0QeIeIB4BhAIP1Beqv8iGSngB50AEAFrdHL+B8tEOknzbzPAHFRqq++
8/TGLaQG+Z1hfM6tHSYbrWFxJb5A5YY3rpDBasW8CjMmoFLVJMqU3C3BK2vBea/o
hAXHb6jf2+Piudc6Xjwv4plaokv75fj7T6KI0r3A4+E=
`protect END_PROTECTED
