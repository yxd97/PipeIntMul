`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dxOGvt8O7TnmFgozqVH06dk1Sp/4KR7Ope8uv98TpxWPmweZ2yz6xqAKfgwEO+4Z
PwpqxgeIDjuop9+dxRK4qx3bvPDvql27pdTavuXtyidRZXqGhHeNkvhJGP5jdiWM
QUPVopPaObzG/+FE+cPylAqL7nBXCxttjjg03+OmFMb75TxbPO2o+oR2AIqofOuw
hirGqL1RoRWaeB9GBC9+I7f9Cf8pSKWF4PybaNEUhdVwX2ejdyamdQZ8RYvm+m6q
SvWaQc3CwxYWAl2kAMhtdBAdoRUpQ2b7Ss4duJaNe6NAXTnZ490rR5W5TmFxmt50
QjgLL4Vh5kjfM93DpyKkPqb+QZNfFVQlXdG8mMVEc90juUJrtwnwFtwlLKyxs+MA
yW9yOz/56idjPwVIBi356Bq3IDwexGTPqHIF7AlwotCCSl/jZvjzLP+wGoVXRHw8
3Z9Rbf1nZHG+hy+NdXjYf5J+hP0pvnpyKpCFhGREHRwXut94XS5CLkdHDj2N4hr4
cDd7D9JcuvJbnfoYVfIHMlyOGEPVvMJpJy2DbUhBEIf46uhacZ3zAGD2aL0YoewJ
KxnrDuB7TdgHe9KrIQfwySxh2pwbqxGwXu1VV01JjVhhaFT7AG08DpbUxeqRF2aa
Ep8SQTenDx5rptchuieUYgg6ZcKpASAovEG8SgmWsSRg5BCU6R4hdn+dpWUpAV+q
k2P/czosl6tWgB09q+aOos7jMgkeHK6OXQw0m5p3Nx7Y1IoeKSly1+NTxzfsP0M8
Iy2k/P0DjENrmUsuquzYFZepk4ILtv/yheqvdiPjAFkeP1ioHZZb21iM4bLe7xw6
49atVutdwOTGEvRN4hchBDfNmWMmkefikZhiiiFMo36iNRreQeG2SP7VsIRRoFoy
1UwzWnaNWSNURhPYZjtBobpTO0NCO1ChEws2WR63CZUaEydImf2OYoThT0o27bjk
8VBA8pa29ohg3JtZWMRzPg==
`protect END_PROTECTED
