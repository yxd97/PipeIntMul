`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1H7SO/UuGS/bwUS41cEad8+cX3ZKGmmjYWjdNca1udo+bwXfyIV75iwtL2FBo8S
6DWsHRQsv0ihnov40XThabUrZaRD8BqKn0jZmSYma20YTysV6iEFcz8M9cuireg0
44RoxY7bvO1o3AJsHAXidURQnqC7bRaBuzRK3BdfWDr+2wgVBmy5+GSpNWnxirdd
xzUXy0uKhravtoyDCJ6CFYNnzBUKcdF6+8mqBhUgQ5oHQYvQwDufL+1PTwTt6y5L
yvYycVTfWO213ZpnAmduUPpzsf/2JmN+M4v3K9N7LHRdGiRTl4vRNWuvXcojOnbp
9ObTs+LQEY7w9BuKzPzo7FdEmcUJafR0iNVOwzo1nw6VEN/xxXXm5r7ZFfI5XkC7
`protect END_PROTECTED
