`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mO6UqoMuVZonGJBEFa4zNPXeuXYP27zPF0KZWlgUtKYl+88aVZtAJk8smPuizZ1Y
yw7ZunCII9nWSl45GFiIqqc7kSCPLJmCPnHd+Ja8xfcIy0X5W8+GlfBejIZsMHnn
fRsgoCX+toBAn8xrOUH+xwotAcHKeWfkR1z7SrUWwTFJX8IwwZn+sOI5kIUkzX66
awkDVLZHkjxuBhUblPK7L5kRaItScONH9S7Tn59IZB6napxonEKO47wABJO/WGPA
M7WP+x4v1v3XXYrmY0KCS3aRsqni1x/ic8EadrcgvZH9lynVgE6Tw70/ibrURrCC
DYOuyR9DKxPnPBKCpfmmhuNa8neLKDfZ28jd6xeAlj7BZegYCmmbHTCrr6bmzTQf
/l0rrZ2IakVa/t6sPLEI3engoFIr0ue9Rqbvjc+sL123+232j9hIm2I6IMW2+AB7
vk0ySc7PlOzPDoK6eArutJU/l0OuTNXswPq1UdHiPuIHObYjcAiAN7f327aThgqL
sUEsv/t4vV5oyy4Y3smtcH09zAD9+miEUtywuOFNsTAHMuaD4ju2vNQJpBT8P2Fi
Hhk/8Q1s+qI0JG4Dk7rgVQUcuK7Dyco9xVVrRJBXNuzYd2p7q7CRM9gfgqVjBFjF
qzQKMMrdl6HugUBTVLkd9XcDjohkotl/QVfAhQwhD+YfUfG9xgyrcNx2YWGb/y6Z
Pmt0aUN62zNMJz81EKE1CAwjO2P7poDjB0sUgu8DtvxIjLQrbgod6w5G65G++m+7
3Q+fWyGN7QR4GTz8MVHOr58nvmkVd8ZGlguxEeDWhYXI5OuKbyFaoOu86Ng5a16P
IuTcusyam2weQyFFZjZAFOJLBqMlqYoHVXsieOejB4Il6tdDy7NQRVK0N4Ag8iSK
F0BECDxI1wyHdFvOADL5GnktDOcNt26xkheAowQOWYTmqyDvOQNG704ik5r132Fw
qf1r5AbCrTFrWe/TgNcmsv0XVE1+svIJq48F0tycJQ1crcH7ZnLSFIiS8/1T9pMo
bkwkHZk57XNrHbp+mV52m3jUAZULjp3P7TGWHaMgSCeyIpneqpBLn2WgVvgUjeuU
RXYdnA474U/MurhdQE5eyEQuMKACLS+e46opBvssXa9alFZ4YwOx7Q7qeGgO7qKh
vNQVlwst5Gvrl6nPMCCVXx3WMJrD3yS0qeUFuT32FMM22JmSarNIs7Ta7ZZOooWp
DZhIOxgTxBcs5+0kKdkXGQQdwhYlJl8L0dk18IGB6rWE6LaldCI7D/CsOMr7/9Pj
7x5PvT+Ls1KGqn2GgpbyYwbrRQrTHQDiX88iW5SiO50zzIahUIJ1G0TeJU+MJrCL
oUtAlPk+6gFhpbsCcTEVrFqrXVLRRoFOELcQs6iEqIhoiPbyGxA7lKsO8SLu11oR
QbIkeFd+5zPVrg9/alsFvulQucrIHDu/a70EhfRBo+SDbxTMCjK0chgKdZ/hfue6
fruaBUQT4CINgrWGJCvzLUhkHaL21qPQv4Yk/dgWUKh0F3M9GNsOs1jCz1pab02i
4a8omICMQSUXThNC1jPMMbzv1LjBUCGYmldaLKjfGvMFtOSWhmWKso9DdPIHPJlf
+t5hAIv4qvyer0eskOqx1Qbhu7i1/c6CWpfVhYaY/QEdf/0NBFAnZPXgMNCsF+tv
9TAKZbycmrXuuVgH3V8Lg1AYXpAHXSX7xtOFQK1h5Cxy330OcG/DKF5ixh9x55eX
7aw9mHRjMXs3olqbjduPtvpIHktZskDRQZUU80eWgCMSYeJW0r7OC7ybghTXnm/5
5SQzTIY28elokjDdvFSAO3rC07nIkpAigwOlpKN0Aqf1rVMLXq85CC8rmfDbPF7q
RCvx90SYM8ecd15INrUI5PFWlVWOQilOz1FOWGwGw9686qBQQ25ONCZq0C40jUpm
rxkStSTMP2orE1RvxHA8SbrD/mWiyfqdnkedsyBbSGycBDBYvRqOn8QnOqoljQhv
+MwTbDoG1nuLG20z+q4qOL+ZBMRKZwqsrYIGP+flIMx1yDvOdmRMA1aMHPKBWLAu
05OsoZ6PJwz7oicq4WGywGwIuHI13PvFU1hlkFvQeX/rX+/RPAL/4XrXDWy9FQ+j
StbMm8LFZmVg4dW3ONi9d38VcHT0/AXez5KyOHNJ0eSQlUXxiaipDmrDcwc8zN9m
QbqQgQjU+tVJteQjEmaUjdvHH9+GfA+BQ9+6RdoiHA1N6Vs28Uk9lh8VkzGJxeN1
QiQqFFgQFXYShgVXv1gkhpSzmsXxEGZAhk/QdtJADpnDIPrBjmeslOACFLoqC3SH
IdGyMOcEtK4Npt4WaYFKg4+XqdHYMEDILG88Pmi2J2TKpEl3MAko/+yDOpjySVpw
RqilnI1tcGc5s9VHHL8vWEfP3gIx9QJ5STw3+eVLVvo0gVwzn10nKZ8MLjrDbupH
pDMblPtco1gTsl+WPi5/Hew3xAfX5VEWg44O4TZ7SAbZnZlQrEhLuzuiGDW9Aqsd
Ow8C0y2jGGH7LQekeFZZFmmuYdSneIKrxagqvWdB9kT3EFgMjcBdWkpePR95uQIF
E5uSaaPZFNJniODzFNkx5QO9wM3nu7ezTeayx8o0D9WIN030ABuOp3w8WiyipT0o
5RS8xVGkKLj6rWk/BcBerJERDcfDeHwBekDAMKXJh1avV+48IzD7jdBKV2Sqf4U0
cNzuII7gTejaiUxHzZ+YWHb2SscD5yuoKnF2lvhQ3+tHHBUvNVAIsBg3Kju3wwOl
SjHddpEe9Kw8b3qFT9sXTw4HPv1iH4Ko0iWSFTE7hcxaTOF9ZEmZcakcneQwG+22
rGdzunKPq2K0BsAmeDKMZZl/AuxVvAfT873NgrTrWLo0ljy5JWDFEscZUOk5WUBv
krbPt9v4Z/I8agCKE2FSCiOpmfNb7Q1sFMhGArrZmsZR2GjQyS9eHDzbfhJMmxpa
VMNmQuzMmfwP8knTxm+V6alex/VSOYLhUE6xTpEyp+gLGYb0hPy++Lky/cE+fSHj
oKy2FtkWCdsOZhSsjnki35D77pKCz0WCCaD5qsF1IPobM7R9qBl0r7IgPtCLhyW1
Kk+BxtZ74IqgEeRZy1lUNdo4WcHaljsErlLKD7MwyZCaAmFp47hg2dn6j44n57Zw
otFCpt6eMlP32s+2QpTRxVJaPLvH7CQEoF8pOggCbQX3N+3Jby84vdlIKukvVs7B
R1COiHDFNFP7tYs94QNh16OyPTMoYBLs4auOSnc8eD7UcEN1pmzxO0+fP6OwNSSL
eqEKaoxzRX+uqAFyZhGAnPNGY84E5u/HpXmAxOKPGV4=
`protect END_PROTECTED
