`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NqJvsXiGnKaLP9waGCpd5BV3eP+v+ZyJuPANMn2B3AVMCUyJDFryTg7dKj9h0A9p
AXT84qI2bcqLbzN3cCFcCa33puf6gB6zbTGL8kW4RLeNn7VCxidUaJmnjHWG5Y27
eB/6uXuvrvePC7/nGPxmSOkGnRiVMp3Iy87u6wRb6wifm3/KwN1v2h3z2wOxFoTh
Gstj1NSRHXJPo+CC4Ssd0lgT6Qpx0FLlvXE1fISyiXlCDLznFsyUD6wtVTd1cYMu
9wQKG6TxxIc9wAUuVwBMdA4/0+9ohS5NTufqoPYGcds3ljm6n/fvVOvPFCu5reEU
q8SgR4vCz3i5wvTwesZBN+OH6ufDi2kxVBbEH+92p5dEw+L+UIOXRwxOaFFslq5L
`protect END_PROTECTED
