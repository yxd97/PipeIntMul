`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xomQs8/BSKez/SNfO1ld1s0RsosmMGFSfT4dPjaQAtuiQnahYGxQf5vrmX1Oyy4
QEbKnBJ/0+tcm0rrAofGiLu0Z9JjE19C8IxScOnMU9DG95tua8gx4STIrwHzWKwQ
VQOthjPIanx7bJNiqB4YDScBwqS5K3ebop3ZmZsTJGcWF1VdAtw06I+s6pFushEU
DwlD2e0n1LpI/Y1SgrEYayjHDpF44bZOm+UWq7nQQlANQH/ZdhTYejyqhdDZ+a4p
7rpC3Tqrq2bEoxI080iZsqQmCgbg8H1oMYdwmn0ujr3NI1hFEAK6Ld5IGnR7c8zr
QQIbHwMAm+nR6hLeG2AlC0EJNun7oUEjfH2jY9Np3DlOz/tE0Oj3HqxxCc4PXKYL
fDg+uOR2WQGdBEVL4Lbo9iYRXFP8ohk5zZZdF36ZdpE=
`protect END_PROTECTED
