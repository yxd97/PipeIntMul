`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92eQbA1R8tPGbLBTiIjv0ZmaB3k08yKFSgUpLT3w3AQIjrGyNbg1ZelUzlXp8BMT
IVt4GdDnwe8f3Dwh7eUL3h1mlPYqdeahftnV6jok0OKBxbk2HlK4C9GeKkX0p0Lz
Wk+ZDvGSMiUjClio5I3UI0ULc7tL0RdfqsU9ZoVtFftdYZpcSkKIEgLUGzCJK0Ce
wE3aMvb3CRzy41RuaMWsThfjb19hnD0TnaDe56y4Nu44qKaiGTVhhDzmk+P4uq79
ZOEfAMmYYVHOOuEgYWbiRQ==
`protect END_PROTECTED
