`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7SAuxplrkqpl9ut1vp3P0LGABq4fIZbFzyFu/Ay8r0UqlvJ3PCCUvj09MwnDaqwX
59d4UQZIKsptxv9QGjdIVM+X893WxKf0BgZVaVpRWXSrbgpShCXsbrmnYo0EdVAc
mFRVwMGYG+llKZNyff2txcGOwvZg2rEkNno6DSOKnoj+pfnqReSFA4caN4aupo3R
/plLQfF8l1E0Ln8S8+UBlO7Hucs8AN2bjQXZWzRsXazZyp/Dqwo0j7ARhgVO4qL1
G/HP6GflhRFP8kl4AK2i+s5ed0mwaqU0ndiT+erfskAUmnzlNSsmd/8eUK8qrgZW
9QY8zJGAa8ubdoN5ADp1KPapgY3hCn6wSBDWMmM604btHANShq79HruRu9vPfhC6
Q20d6VkTOG79/C3e+F0tCBLBqAmw6isDHBeZKFWO8eCstNYCaY4qnv3zijzakBnn
Fbis8FEy4du/7abx4BiI8sgE2O23ZZmYmI9M9p3kRw+KPqrIKjRm/STawX5RmOuu
9snBarcXEC9GJ0i6f+QyugJTtkqkim9LLRcB2ajhdeC9fEv8kRSbbjZIFfmv1y7H
tw2WMP1fnHMI95jqRW3JJg==
`protect END_PROTECTED
