`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9pOHOJ2mdPEwmoIY6EGnvPeVjp9oLG2bpRcaKL1bu+rS5/z35mkJOloe65i3QWFV
bVgh9ETtt1JtweMSEvN1K/0G2uY+Xz7teg+lvfmpwk5q1GHe1KdFGcNX7bk4akzE
lqwtNsve0auVXGMjqogGql92VOZN3uCCXY2P+5c7jLmC8RRHN8AonRQGj3tzQx6h
/q6isWRfXKN35+cnVfwc8lD2JCfXGvoefZ1vaREg/LcmKAOB4BLt+D/mv3bhSF4F
zCKT0Pl5aPqnEWvgx8lgFxQ23iJRsxKC8aG9C6NEO8UvjsBHMA6+Ay1um2YpdCyX
u9lD5efvOUe2GUnidVH75SwyKcnLLOEywrr3BpH3np47ThFzeq8L56GWt7FEzLCT
sBM3fjpye1JqsTiqWVJio0vSAznUU9VHBz7Alg18Pv4/6dpylHhtS1tCsMWjUIZF
8qewjNByaKi9l+Brl0rH8oBCu60SpKxeRgdQtrKhrORv92zKD/dAHW7M6XbfX5tM
Bfp1wkpPnEfATWqadkTt2zw+lFsM0xqmGkyvpSDghZ0FWighYEm+hdI6vbLeNY81
vS3GqC3PS9xDa8tRgc6J/b0CrUG9AW45Dltcpth6qRNhyp9WEAzbpqMHqgq2uMfz
pSNLuAg6fDsXDzYdogvkMCSIp3Yhweo5oTSCMzWDa6CQsWBGq8QCUqgaIXweE3IR
oqG6nOHUxOtiCwkbLIC6Hu69FutAvFEZi3hUYUDHMsG4aM1ZCWZWBpDNmhakS+D8
/tsV+FXRcu+f1YSmNPFe43TyrwdLmCiOPmS+BBQ7yeU4Ow/4MflcFjpXTfkamGff
gHTgY9PRrW9+zQ+Chz5+pL15fEAUPz7HnkVETKbx+U8xUfvEtYUCouO8xFG9dbGv
9WljJjqGej++D/+MA/Ic/npaS0IvvPxTJtf3CgoRZ//4lJQ+Q2WhUWT5D6n0Z2hU
CVw65HlzCZeQp8wvMhcVfj6WHfKaszq0LnjdpNYc6VUU+xb43U2wELdkq+HEdXkU
tR/rFwieOsTUcPxwczGFZlBdL2lKlx+i0eFCuKA6rLPuQqY1pnp7pJTLXQ6UD1nv
`protect END_PROTECTED
