`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyPQXGUOcD7b5YpOQUQPFTLZ+DYS9adl/bsLZxRCKbinIddT/1PW0juNFvJKtXON
0DKPBKqPkvqSmJqd+YqnRlJdISV+v7SO8A7Cg1elCPMizfDfl9WyrlwHFrGZX4yP
u27XRZpKHDa7ldvhUVRBVHsLp0/aKGwdf2PJf2EEVXnG6kPaXy5cuCspqFhqMeVa
6RTS7grbCxkXWExVPm1Hj0Px2NLcHJOt77IAooJeUVWbXiwrmVhY2G6aKJecIdtM
C8bDiikHjMkGyi0FzR23OYuVrusYLelT47n3knG6oyqnvydoqy9KprTUHF3E7xrK
ldl/JozzRGb/f84QCmEI0gWcKJkV3oQsnMEaNvS7aG5MQLhBBFFrLJoF6MAwpd95
Y54bFHUndlieLQE0Knz3bfDWavpA05ZzuXskn5n+YZbK0ul1alQ3bl1cZT4unFAC
aRocJ3f9AxDuOTXisqMpcHCIw6C9xfNkOPM1Df6Yb3MGekNzQvkYa9g/7rORrkrU
8YHzBWngDrXYmHUHPJhOUnqmzu358pBn2esHLLkqCTXfYSCmstZSTjMEaeyh+Eg4
aVnFPTjA9qZHodrseWJsQFY5Lzhc3Os/+ewXIB+vqkXeRgBYoHVFlVw99h28tkHc
q1hSSeDRHEvBP40+PshJmYQUBcyoF3//Utzpve5m8d493kUpyUV54SlbwuH7gKvS
amDIv5wJ/w9f5VE+kEh228bYX6KLIjC13A97nwH5KaAHeJqOUam7TxXRiNms4qL7
4OWs2CEJv6kcKvtAV3qyFWrUzkCp8earFxfO4hQblsl8JfbOPJOnWBC1v9Gk5d9j
xrC6qb4taZDY1C7WIs8oro3NZx0mzFh65m9513DM7uHrzZb4bYS/98G0ft6bGGCu
Dfv7jbrjtyDYRJ5o/gdY/eWnBKF4o2RqefPl5M+9+veYuHpPcT+lQfpMEEl69jrs
a/OD5Orhy0KvQ4bK55TsxcFxpx6qGG/U42ujFMl/Zl1apEJrYFCxzC+euLMH/6Ry
L/MhqMxRB+qF8/8k8yJEEnR+H1wBLaSwrjJdemP4WJcfHWP9bR5WEjE8wS4tEr84
zqOcT21AoPiodvZr6xCOFz9U4wVeAsD5q3lktbbdkQuMEZgAE82IXIEDvXvPkHbC
MrkHsxkM6LdIv4YkvmvRqwnDLK6HoWDKTgnbz4mY1XOV15RoObRbzrsFiRh91ur3
7EajZDk+J40FhI/ibvhpwjzUX3Zh+KJz7ctXhRqIKB3m8Q+IEfaLi5aO2JCd1Xbr
U5/qpSoOzpmTh/c0PYwtkbANKwD21s2pAE/2GenKppuBT8wGUCTBPKHiGxP1W58h
s6AFc12Ip5Bav2pggiR99vMaaoQS59mGi92FTZnfWQBXrVjdtS9P4cA8oqlq/qwM
VvGyUdpodSJDgVKxk3jhOmjaqA/HcQ8KNl79cF64Q1KkSi+KAeN6CunYou7K3Wzx
6LUVXwuWFSU0Wc1FoMyHQjOIwogAqB3ePUztGuQBlvNhN7CFKPau2H63GGwOKcq5
G4AkOstzpKCiA8zXNYeOP68vHiyPAf5fsqsAWhSjR6aCr7DjMtT7mYYeA+LX8+Bx
9hKdBX/WyMzfks5ndDtzLypEVMoTsCAgK1sgLxFLpU58AXF+3Xy1CtLyk8RAMMop
SklUT3oDf4LK/cnF4Q6paBWPDSsNWpXicYGkwSN0usiwrTMtFtHr/UfFu4JsVgO4
wNlgoMD8ygckZmnB48orAjA3Wkhlu+xeL3kw4ta3h+SYSoKL0hBkj9HrtDs/Cd7J
`protect END_PROTECTED
