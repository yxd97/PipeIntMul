`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dN8DjyAUPowDTvE7hFtPqJyLqeAhmInGYgn+YvbE548ffM8kMq7plBXgc9bESQL9
nYlakDE18Mv36T3E3LQBbWUr1bOFGdETg/DAl4g6MrBtqHjEbXtku2ylsPkfPWpV
ItXLQpMzt1OCPcjWGr6XCA8TuTnk/l8lfMnowS49zONrol7diRLUmXQLJT/YBBOk
+rZ2WN5Lr7b1Xf0INscAysr6XmDZkBTvKEHztaYDG3ARSG2HJxLWW6ZQ+8wj3Cin
3Z6WlJ+8ggRwQMWfy6JaqSszjtiDdF/nlls3aewXDGBB1Ekd+0eZwS25Y8O5QyVD
9TT9Ua/gD58lsT2njlJHdw==
`protect END_PROTECTED
