`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
exHMgrmXWysGcSo1Ci2svrbYFcLJ7poMBDkPgR0sEy4b3Qeb4MyUonQQwwMgNVHJ
CPfLYW6iBp9IyFFRgnykrR9umbFDqwC0EvwqeqE0CQ4vI3sWtXgcydTeb1bDv37u
fgf2f1/nkUq39mhoovIxnylcyRLYxlxyfuje75ycsFeNDb/LrJSA7ClbDfil1gsj
nf4J8vReBI+bR2YCj1nyF/yIQp7NdGRwo4Dlx2MdP+q7R2sEY8BXOrUoby4jN6bD
WEiFzP4mVR/oCLeCe+Hp2Trn+mv3ukB4tBKZ8sXElGXGn/L/IfVLzcwvUyF24Egl
GRgRpFm9QSu+SEeG7DrMwJsuAPeWvkfHIOXS3rYfAYiiqpRj0Z0Hv8goDg4JblvW
kH+W5CoZHLBKLQM0eytwH8THeJ87msNUse8A9TryKfZM6tU6HLNoXGp3PhRTo6cG
kLl2nK/J12YZ0IUpyo1jbeKqIy5t9p4lPBBsvsU7nXW4NzpCAwlji8A3xEGt3dYi
HcfriyPB1+B9CENpNOdsingg9hPhXZ7RdL83/xy2KQnuRF0Fu+W0s0U0HFTgqPZI
9vl3iCzTQ5lbDtHGdA0SYb8ylHHMuef8fAybZGU+VY0fYM9kXnGqEB3K+k6+JCx0
L3aWD388z7vS/q/a4qNLYAPbLZPS9GaDu2vVE3RexmtgY6qHcZtNNOl4mrQax6K5
jRktAXufRp0lrPDrVzLsa8azfLi3M7pkBYa30p5VNuG32K7YgUXPKCpMGx7V8QhI
O3noXg7DBDA9DEmj25VlNr05R8ktIeS0O4P0BwSXFQyE2tYsTk0AEm9Nhn5+0z5y
ItoFPrFOESp2j5dPJJ7loQwe7oRJX5GS4K2eUexdVWy1TaLDDVdhC7qb93XhIyYM
Mo5QUxMATcd9yW5fruXuwA==
`protect END_PROTECTED
