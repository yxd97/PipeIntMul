`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzxhQrMVEan0dzJvAhzhnNBarwxRQ5PrMvy0exencA9XbulG0LD5GWBn5GinQ6HA
h3I3ipvY4NB3Lu92Yv/Sw2OqLIiCNkLu2BtKlNsEsa2PKRTlFcPyZWx4x1FDrqf3
AreTRhIRsi7Raofl06/eTPEMRtTeEO9ls22JMdxP5cv6n1oWhEw65MAPgynOQCP0
PjFOaqzHodkcfIbQzio4x79e5ZadUz+K+tBepUnf5W9AcZOmllI2msILUe7j9ifu
Zt/LAyt8eMRdYwgzOLrpxdOmIdZSmgCvenAEdK1bmdXnuMmt/Lx60s2Cq3v9HTVS
kJPuRv16WWQjw1u+nH+wICDFshg+PQDXVeeSrJgBkhYWlQVfCVF//Gy0rliiUPew
YrPM1j4wkGOX/sfc8vIVHB0Oyic3zDYVBGXYG78JzaVi5StDiPiwc9D39StBbJOb
0sNPCUkgUv45wv8lxEQ6fdXNbmkuok2NY+7J01qjCOVNUORDty6NxAf6bOvfsM25
56s1fYBEOHEhMAfaMmTRShPWuVdSD1HLI2dFNIz7ON5+9xa2hRwGa61PST7Veysx
/gIe/WMYcGcPNkcS8OfEg1KEjthX8lVh+1NCsKx8tezZ2EA4eBklLwrg+RZLNJEB
b4QGf99r6gTM1NLIEORYeVQCfEB/xEOjrQv4D6xkIW+vf4l8wOPLfEzxVWudDUqQ
9Q6Vd2YgOgqR0c4xg5GRwnNissTB/HI2bpSGl3W9WuhK8tww78LBzBmEKOqLWq5S
1+c9lPkumMDOM6txC0A3MU1B/VQYHvcTLANN66e3ebjVz0b0DlY7qvLrMcAwrW0G
WTXYSEHTIU69lzBBRv8uLXDPnFHiD03RhdsDEId1jjOR2HlWF+epbbzQbIspQ2t0
pBZv3Ao2uCVGDGP3HMrpfVAqbfpUzMeDuxs+FqHOXcaaQ0s1rPOayTUwc9Hhfnlj
km2ynxCx43LT4OiR0qBa1Ll7nuXSo/dFNgKY9WLPgPOz9lujm6RbOZKQ5KKZ3+pA
coTmlx+F/YYvhfVS2iG8mgenZGF6CMYyyCktfYaC4+pDdIaXNWP+GKXt1+hiSHrA
l+gCX4JZ8cS6HackEVq2UJrfMWug/1ZaIXc4a6EX7fvcGz6LPs9V4Xs2SPfZhgIR
qxRFz1lgPvI9apB0ntRe4V5KOqzKfoNeG7t/z5PjRP9kVun3tZFsNVj1xWPH9JW3
GL0oaFb7S/2V5Rv9/MFmPQNUDt2br/6CHGwU0MquyNSnA9h9Zocrw0q4tGpKIvwy
P6dxPmgAr6kYWdHPGK4Q5PDRScW0YyAGPY6Gq9BRR+IEgQ4w+r1m2UQuQZWqPFlm
YZRCSZdE8L43kTd864sUVq0OpIhCbiIpHQkgH+rgv3ELkB3YPma5OsmQc2wfC8gz
h0FJinQN5TIVOZHAIfj6ZJWDbsBRzfdkAyb/zWxuaw7+cGB2l+yQ5S83HtfPU7mH
gYTptuzBEMHoj2EarW/ozQm9UpqCIz3BchWKngPRNNulwrIJnEZ+HW3vz5m7HdWJ
BU7+JnX/RL5NL0qVTbDDSK70lKPe9eG38zDY/hZySjSU815Va28PWeYqogHF4wAY
VKo3xGLD/16OH2Cf410ekeoZtjqjCwkfgKqDeGmN5Ldzt5SmvnRXUaiigg+m0gfF
bRtOrQOX7XXDQYz2arKHv+5+PQTdhtoNulnyb0FoLQjE/bsbkBlaQcaBnxWpd4ea
ChVbYbs0+PV00/siDWXUEl7gu55TdaaaDHAmlQqrYemsphtLCDpLirPeRyuKGqeN
bKhoN/fVZeFPRcJ0jDxBeo/CNqN+UzvdJhqYdNCyH0DL2+5DxUY54Eno2swRIzBo
Aw/nGGWjDGHv0kqBHXxcmNgxyfnZTjE6iBeiGX0SWogi+CbsnIwrEjGeL/ZiYuV4
RrkLdlS3cTe4QHJ2IN+95Ci5qtBzrU8UZe8C3/DVb7tvGpCpbFN9s8DpHK/xZC5d
bgRB5tE5lmCs7dDAJj3IX4j++mFodqFxgzJ1SY16/rQ50gJEzUQtR10PiKxAThp8
2FDhnvQQ2mUDNK14ubE3CEOMp97Tb+Es1VClfPGPQGlM5zWpq+pem9ftOJgBHV60
nTJjvlGTpxMKNF66dWN5AWlKXc9IqVSCKwzIOVaC41+7iOCg4cyta6PhPqGqfxwL
70VuQwD9DiSurkqCan9FCQ2t9HQnfG1kCnTWH370XP8B9LzQZDwZ+JTSIj1mnzC8
mnxRM3JE2zbhj8hbCBJHUct5QnrBMu4jNVF7l1VppLNZz1Fct2Ql7JjqJ6tTx3V9
wW6Nd30gviDShxtd4SuXB1QktI8+u3Dp6rL5qaO9D1KgwnTO2kVExdr0n4uE6TXL
SgAYQVDhtuCVdIXgEqsG2+Fi/YSeJHHtNL2ITBXObCB20sCSuljYvxHozTu+LMB0
BUsWkh/G1NY6zCrQ6Ch2rcdjP6AuP2mAVrcHRgZmB2evrpK7A9hnWQbbMBMoqdTU
usge2aL/JabAW662rEQlfnuJ9JHejRs3WGFhNZ7BIW8rpEYP1RGe04r4/3piylb+
Nb8aFjjoRkNjgQ/THc6nnH1ktJ2+8dvW9JXs4KZLzzwPERLG1L0o+44k60KvFIyq
t9bBS3Vqhv7CnApt5ryVlTYQE4c6ndxb50PQhp86k3tiWejlfNjPDqonx7Mnv6dp
UywL3TRDF9zkgXZG4xTzMQjT1Eu//05KiqQf1FX9GYPCVpBZRIl/GRCiiEgytBWS
ifr4okTO5A1YCJ7e5ZYde9wcUaq4ACTQYwhRd02FITq/HOarsaRC/u2pZImY+GG0
WE6CFIcWXM8Bq22LQwJTve5jXG161DkWA9Y3Wuo2nGR8msSB6W/QqDYoIVpX47e8
KUyUdAIz/2Rg1ciDmdBikbbfkh9wd0as2TAApFLZSHpo3FLt/U7LRND5XSZFwPbC
XsyiXETyDXXB4NUkNLCcW5BRLSorm7ApmXbQpkGEF/XGqbN7W1RcnpvVXvKLKB0y
iFneyrglKIGg0VZ7aG+9QX6+Hngb2IziELEFlYrfMEvzV2BzurazujH56JBLW3/6
3UU3GhGgL8Hvmgq0BeKzjKt4nwlhUGMSm6B0ENEa6BWENK3QItjCUzFwU2vGQZ3l
QglLLZnMZB9pXxnFo5ecw9pSzQfk0XgnWnSs7QKG6d5SWSdBBmWC37DLsGf+Fspr
XM+tNCYS2eBLUXubaSXUNg4MvlXQsBrCIeuUaYy/xMR1QbPB6UdAeD3tBChkRtoF
NLYLnHLFz2dxJcPONmvlzF38n3Hcq7ZqchuJLBW8eD2fkNRomDpP1erWyBI4PV1L
jR8SM6tGbVLWyeE4Lx6n0RFnTultRljXKUCjNEqqIPfUGyhFZXv8VxS1rvSIiFzb
rHg4JHvyzflyDdnagILfHED9k59ax1doDVAea9dSpTsJgScPegiFW/0rvisTLEh1
bo5YH9wDXKM0scDP6Jz12glJhvvyft3UVI1iPG4NbdVKWpdXwiXvVly0OnQwZ+Wk
J2sxi9AvPWGK3i55q51e3OtacANSb6Xz8/C8H/CWmG1ty6nKYfhVgMJgBtw3YocU
Kzd4r0/8v54fuqS4S/IHypdVeEI36WKvFyIZal0Drg2/nrcCoq4fm6TxCw4TtFE6
JeuMNg20v8Er1Ppy1GbZ0x+mMsPrmowXBOR3KTfz8Ry+xaoPs+wmFjS1BILEQzFw
DnsHVoe3jHNz/rZb5Csk0UjrEYb87w7vomA6PAJc1/6sSCao5XN5IikQlYLDRk12
2b9DfBNgy7cPUdK7pI4vTF8IeTC079jxLhaunCLvkHTf+2SZF+CbE7XFlO4UA7qZ
dCXk3/uoS++osrla/T1Tfxc/f1P5bFyZ4Zhm/2EAvM3Nmv4pC3ECo63FjpU2QSNR
mGfddF3tW6TI2kdHiYwdAIQu2/aSyp7usLjKeIClha1JBPJ4f58Tx6CBjhCc9ipL
bPCOm662Gq2p9R1vgz3Ct8Q2KzxbmNSLr5NAG2ycqMrPeJdT15lD8z4IRpWbEtmk
JEd8ulcPNbpjL5PoDK9erOIfSHpYxQTJ8kpVuzCDp6mYJ0Wyy16g6vkl/BOjF0i7
3p3/MaCP1srxH2rOI1bhlR40Wikg/Vp/vftNyveZobndiSh8XhNYQ0QcjshxM3xL
i8McWi+g6AeqWZZQPq4iov0aqGeYtA+g2LQvUo0XW4dfD4P30Pb/CarvA3uRBHA7
t9v9Tdoi3KAg3l1c+0HgDroOLneMzO352a4hEq3G97x7TXaegROb0agJN9GTvbzt
tKibaLbKYwgzDwNmvifRDBE9uddilrtC5kQCabYXscAxNrf3/TZHNjm0SM3l0vVN
nyAPjEigtdGoflnxXF6T4e1yHbisygiPhSRjVjszcEgy3zPrymjLEZScAl0z3xSr
FYwsHilvA/Y59n1trxc2lQYb6dJaCNHf4CdspAE/Gv36U4morv4A3VuthfRGdQJ1
IDNkSLtJbXTNdpjIRR8ouW5hIq8dQJzNOfqZ6UK3vamuuvvO0JoyUzwf7ShXSsPq
8+pO6Swxb0l4etuI82aniNVcl4l2a+qnVYvu7WjH0mAegCiUUBPL4Wr17rc6eYEo
uhgLU+n+WM+wc9x5gQGh0Do3reWmjrDLVe09atk/1Rbb9VlrjJPOaiICmL+hEaa7
5VjhP3U7V2FBm0FiHE+vSKUR8sdcnHaPzhab4JmSE+MnW/IlyJMENIoxVzjVtG0R
TTFELqsp88zBQ075t/YbLK/fyrNlYUjrmVD7yWpT40GplP/k6lEHHMnkTXo+R071
2bIlmSkqECefdqw4G26Zq5aruS3LZkzrc28TvgrQfo7Oxit6OegYRedOnBgnkIbA
o2xLzaiz3Smw31JSO6hdR2AUwG1TmYrw2ZNGKJlKubkCqNPVsu1r5TvC2knROcs1
UyLUDJiVDSZ+LvKE13htCaWRlVJfWSJ0OK7W1RVtN97G2Vp3Z0KkbB5gO9zYZ8Sn
bXAbL+a0Eu9ukG1chA+7X0QWVbb6bP+AdRzBDSQjiN+eT8pYD7QwDNIqzFAc2W97
JTvVaxW6JKCSbMmKfEeWEEZ7XQM0Z9N+zf3XDu9mXU7T1xkyEcHg/SaDn3/Ll+ha
/qfs8HJ3Kw71aoPq4t16gJNAd0e0yIP0Svx0pV2HJFQnvB9HSIj8tAQAE2UcNd/H
V02ulMSxI+CPFA70EQ3L93e7A/9k9rOSUA+AwxOmLco9U9cmp9F6BKwK8VdnAr+r
xK7RpkJpbKIMzrXnZXX0Ej8uvoSjv588gn36EqcBXkWOvMwhR4h3iBxXctEv/+wt
0tviwDwZ/FsLdyg33ABNvfPTjB/psHfui3Mkwc/1GQJYgJI/7GESOa3uXQo5iPVX
ctEclHolGWDH4chrS0m0gBFrOb1FZiC9OLNuGQOdIERnRcp0O1aQW27iRA/+wFW+
xZqlkSP5+xulDoWRNDic0v3wz08X3OQemVZYzk51chuuvgXHsjmwXGEi7WRFyuVu
DTZktvLBGKbAjcwzBaP09l+N9nKzv3mCVBcpqRodhXNjZi/U7XjYsnu2wmSEoylU
QbZBHvNwDZSN+Ejtt/JjqLbS0PwN3n5P3B9HnyHm80G5/u8QkelERXrSc7k1oScI
IXEJ7SqjYI8h7rNzPrUJfB9rfeRw+ZuSYBS2bQ7GO8XFclknwqjP4qKBHSL9zmSg
eRRjj8aiX/lpEJ93KR1JFr5iYsju+z9ZRo61O0sAf680/bWgS3C7W1tXhcM3elQv
iGYy1mEp53G38puufCrQ1GYKm7y3Evrzs5SBziWmEcvyxbrdlzFCZ590676ztOE5
Gfm1GfOBMtPb/DOxuzDFSkSeDZuHoHW1F8OHV2EqJUqIjYzznwsCXm7w9lrWamPF
qtTUVcH6xE7u5pdQRFSWysbAfKUAka7B9D1XgmxeJ/m3Qy0DPLaffLUgUe8LKey/
pHE3goE0InGTeKT4Jzy9vYM604ogBVpxZOpTY6iJtXJk7nFk89EDFshMf8btQUp0
DWQvzF1Gca5C/AKC6UUR5NkJHscoXQgE/evKt2XQrnKX1NiZVHmCpyqbPDYRdtOC
WqxvLlenwfKHbHjenNomYCWsg6u8PtYDlRM3URf/eFXZbqpJ3m1VkNrRazimK0JU
B4SawVfkoKZVr8gLYTPLrHh+eV2aWbGZq1joENbiQKCXzvy89omZOL8Oec2hb/59
xlF3i0eS9SDY5HfxLc/34YLbV4avUEBGgplvxtriCWlrXkZMtE7VIWEYFbrilUBG
1qPVlBViOwsYuGd0Fig6/mL3KF4wyUIiaANcAV8d03eCar5NyOzVZvqYrMzi7NBb
o5SkSh8JfO03DYiivAHrUa6Co5vst0RjiFTz064jYB+WbfkXk//8T9uAx2QeM/QT
Jknx4LwMiT5sGuwavc8Bl19a1Bo+bZP6wep0hCvfJBVKu3QuQioI8XJEmgyoi7os
PPE2dxr7WexYUZSZ6KMIjUzFaZbeHL8J+puB1S2iNv6V+4wJzq+qlNC1FYt/N957
BcoSTR+IX6wDm5QJxCw7B5CHRagzZCFnchLSjWWsxROKucF0xed8uX08br8e3IkA
/ixDimQVTOL/7G/is6jiX6D5PfFsPemU7w7E+7qvNlsPDinc4xR6ejjgC6MNRzJe
5cehU+mhluZYODC6Ae7Pm9dbWK8EiR1eIVfNpHGkN9/QKUrSvSNFgFNID43wjkCr
8LPtASgM20KYclUBfbIC1ESjoSbzrpPeknS+P5n75DDLYh1rCZZQziQeHooGOSc0
LfyliqmsVcSk2eQuHHVK2+7jyjLhFfh9cgSs7ycBUfKqk5QA5VfN9iEdWxROPxzU
xgAbwigCwwvdIbW++1+ZJ3B0pKx/qA93700KJ6KZDIx/YhNTPdTAzupOzsT5floi
ehDc54nyrWmsjbNpWkQExPKFj/EDIuK+M5qlSa82T1zS721a96S7DpD6JoSZNCJ7
0qQJyApzFhkoJOC+DTpClnedwJ+nqJQ9GljylnEiePH/eUjMrMTC6TAQ7DNWZKNJ
xvp1Ij9j4soLjLpiejS3eM/zSsAOeFtrDsBBI70ETY+m/4oDfZM7NecMysCRJUhH
VpdsXkCtFT67qZ3UlC8C+Tr7dXXzS++2aVz18QNlrbn2FmogEIn2UtQApBGK/wqQ
6QdWDlPoPkkknRdzmAwVMr024yHSlJ2qTQbU2JHKQCxxPi6zWJBYPVBNIeAMDlZs
7CT8pn9CMbRCFIOLoEftLFtwl9+eM3AOptSm0umyEWGvH1kLevC+EPMwHZ59Xwac
ap/ZIJcXZdFk2XxYDgAzyHJkVkiHIVsjJqOG74biiWTLtiFYhN8nqo4UawJIqLnt
u7jqwAt9kIoVYB6mXPvtyqeEPwiJlMAoFWe5lG4KNh83CPtfqw6aa8eqmeYfNr5/
hXOKbQ907LHHTG16/w90G20irOS9yormsVhsLYTKdAPUZtNrg7vfqIXm29zvXUbI
rZd7DSgA3QfZl8cQh12B3fJb/mwxvDP5ZEv9ZOWqkGVnS8xiQUZV0fFtz12NBwCD
E9TheukBmkbUcJbemGKXXe/94QNdKTigD9nYex9a0BrrdxAq9zuivXCWpc1oDDRQ
UpgV7zKug+4YkTRqJjtMvgk2vihawzt/ZhpYzUHwRqnXMyY5bebflL48fu73R63i
VT5PFSwueBXSWI+ZxowCOA9IySUQ/xD3ClyPdJYBDjZWwsHE+ryztvTSsfK02IRj
MMU9LpHpaM3Ve7MlPquXIclOFXdrVhwhWoNqgBJ7Sf0Do5rRvDHMstcYFcvGaf/g
xZRwRx2U68HbKRAhyBQpFdOgThVt7IFFSUikzy0cOhBuTcygN0LT6FW4bT33/Uv3
N0/ODDvvJ1BpRdUuR9WfGL2+IlgkRSZEbA3MQ9BzXAgVShgmkAuy/O3coy4WbwBl
2EmdULgoD9L5Si6pcPYkZRXAOxGJGKYI3UQGLe3a5RlrUHLJv031QSgZv0Zdy4J9
zNHL/11jkE/n/vYUHUTs7NSdmnt2jwQuxs9U+/jHIUVByfZQatzSZBzFzzogWTHv
k1Y/FljoPhUAqgQrYyYiZJR4oUSBHzDyD/HUbrHhUvzxQSxwCr4wfA2zA84oTQpQ
nuAQqLo0E6fp8oYWnHywgxEBGpeHOws9hDszXiQnNVbhBnkhwwGwoJzoaYqFJlM7
TqiUatzRUhEFSx2R+pv7bIfxtuY3evUFOGwLLV8tbc+gc7eWJTsYUmdSytRBoFGM
GqFKa3XMqbDcdMdl/jEA44LBtJEn714Jk2rqqwyG7dkMbPL+MCT4FXPxiw62CLfV
PdvSPQf4mwOH3BKeQ0yJEm8X1CH96V4wazk7kVTSqAPVjkUatlyiDq3xczA6DUfH
Yit7+NDBSX8U2FmrMCNORlhzpx3XGTE1b9+Y8XuGwmSfo6Gs5zOevwSkP1RfI2Wr
v7fFSM0nYoGqC5zPjM2XjuRXwPy6fvYI4ExsG8xAaX2kLH73YZFGoY1aE5QuehV+
LhKEeZXaV5vp3/DUCWRqQDao6N49U4aAj7A/4Db0o+W5iSr2bRNGTMYmLDDpbVoK
R/pp96bCA3L4VCGi27iekuuF79GdlmUKQatmXF57V43IBOh9AZblDWaM+ii/zmiZ
pZR1LCHLH/wmVo8KiaJMRs4Db9DTYNNq5V87KmTk8mmROwT60K/UYDMB9FnYh4Mh
YHx9Rl4EAPS3wAh8Cq14xdsoS+NdvQPEpF0vqJy1usYGf57oLsUivn84b/Wr3vlc
34TYZulLEQppS5F1gSsIq4XAFJZ5RiUPj4xjh4oC/IQaPlHO9Klu4GQHcD+2EJsi
Oq2Zao/QKsjSLTUa/Hl6ftMw6H08Tgd27G1KF4NtSlPzK7xzDKeDhaIIkS5hZVNx
1lMQfBbIaevb/c1aBYfuYXNe4VxK7+lIYkDk+tJR0vTMoPa8IjIQOht/Ye2zsQw5
2BwPPulr2GWWhRMzXV+WG9BhJ9QX8E9cHcoQ1acrUoOAOIfnmv1nMdibRoTabb9f
5CDzXweZKnfvV9Ugyxq/8n7FoCoa+rT6oJFAhvFgu8FgkIl/mtOshL0JJxmt51IG
UGDq5Z1RkUPwo1aOfBX7MI70oDYMBaTluNH/6qt3IvIIXQHCqFKAQDnWrph3Weh1
oRWs2S7JATN2zGEBXB7owIkB4TgCZ5dPuz0WHvLeDZGmNdn55QfyXSAl6Vaef2+e
Cqv92jB/uxjHl1+BY8D7P+c8R+rbQ9Q5GreZDL8jOEv7NJKtaqDSfRgJJbUH/Miy
WMJqfyOeQYC9uIw8LXwpiHdHF7mn/L7xyuEIn+/eIS6Y+HFHTuVnMCss4nNHlHJd
X1Tqu7QoS53pIpSDw0uHRuccNoXcTlmgRlZnZFKsaovGrJ9k7NIFp03se56D2aPY
ZVEGnfnu7MIUOG4DrWoT/y929dSdhuU4owcY2ZASxKukWNmrN/FYviQXQb2ft2X3
YwaiJCaVEj79rnSkbIZYi5PN8fgPunoNlRHCJ4oOyeSVIKtxTl4clSbPiFzL5XjC
cMJUGigUSXrue8D3Tpm/Hl3yYQxpDxXlC9jl1b27pOqQuu9Ri4LrXbM5R2YFri8a
C9WHAKhTwOwuoFbv91NmcvlsIwJmBV3WyJlI7ZUN4bLDdOXn+u1EC3FqCp4kDAX7
E8mycYVYy9VN2aMrk33t9h6+JI1D6UQvDORlLcrLjQXBoV7ZOGRxBULwRi6iAPSw
RjWdiHH0bnNWMXkETXRwl3EEq5cn91SDwv55nAyzR8KwQT4X18w8mvftW0wuW81L
Ymb6tsdS26IRMUMhXr8UhVTgjaqDeg0ZbPrrMlUg7z1nz3wwFhCm6UApg9rsmdSq
kJHIMf6oD1eNQcqJ7nyiRaQL3FGo2Uy8BBa+/mFGg7s5Llg3B9bANzD9XkomMnMY
SV+LC1AbYei0hshFgaZBohRURJOaCgs+w/XTdkenjILp5CD1z7M1u48dd+EUA6TZ
gZx/VdOdskL49Yrp7d4KZypoTAO6/+6YKIJN19+qSgMxQOF/0s4Z6qU/+wOTbNXf
r/C1yhmf85ARPCoJj1YrvwwjXOzXhUqd8fZJYa9PhOZq6oMjnRnHbly31UDrVE39
9mKg9PFGwxJvANzDBw8N2B57OUIPkZLza9PRmRooSKQePbCwfnDGLgtD7gkB0RzC
E88n1pxSn8dSZesPArsmwWvd+3GRf9MOxZru/9mQjuFucwJYSrx6v3AnqJ8tnqb9
o4RX9zUQCP0r5XBM7MHdfERx9HDYJveSdXlxAmbufZAC8h2nrwxWRX0g6P0UPk5Y
7ATXuOfftQgS1htwXhJdv4R96k0ZembsvWp0VZJbFJJW5HEy6E044lEVS5xiaMkB
LvrA9dZ+X+xmoTWz7gVymL0YIR8FheNF8ja2g4b8PJ6ZK73Gefa81bWuR3xUn/jN
obuO+sr96lp+7UK9P9pXnxvU/DAQZE9nJ6BMIVZWZlMnqozX/qfUUKhZMZb6uZSL
kDrL6RHOcCq3QDh7MzIVKEk+mcfoPKdbi4VzgJ1r94ynqjlMrmLwLrXxImpjx+/8
l9BpOg9f21nhpGgOEFHV5ak89EgrfOex/En4ObncQhkSMVbvZ+kmwMRpbVFbk/3l
9n10RQ5sDbGJUQtb/rWU1izbMClE1wAeUTFQihXHKlLBILMjZN1/kAMenSx4Nxse
69ThvX/8iUBkI/dUorTEY1bcL6MmYojjN1KrHN88tnmkamfndlm6WkAznWp1G9et
ijjDDlWNtHkFOzznkZEsvk4kmXDEyg98kTs6kx8YVqeXznaREE4IpL9DgIbwXKGc
NnLT1Dbf69GufzZpyWjyR0WZM0JTehYQ/4HQiMnLikIam9UREfkn7X3KvkfKC/Gi
blq67uVaaEpFWR45A4HSvHSqHRYaXoePospYoC4aJg1c2cjEybIIdAB6Eplme7JD
ooi9QbI2NAyU6iMcsBxMHfjtKFYiTwy5Fsjwpdjj5787AfcfcQXSsdr2IourZcBK
9xV5MgsI7i+pay1xJxdzaPc+oeCspepYBpRCtPMp9AH6uSJbYb7QvF60KcCoKaZl
iUjwxoHBf0nbrrk2/hyHKmna6sLJjK5phgiFOGgR6rcc+XDKwxVW02TiqUMCD1f0
fzdRRfUFfOu2TeHvVWxjaAaf0Tv+modqtq+eC2hqgcRgQqRvJD9nO/xnKsRGTn6Y
Ghf1BVRI/D/Exqp5UoKy4HW2dar+o19qVODK4M5Hg1kBYvgwx+cZVxzfzsWhJJCe
tvIVmSQtNLNnaZZHZX1ifh7j/sVNC2JZdwVe1nZzmyEGspDQhvswaPjrqhMgVQkg
7Zj0XOoAh3fZJPtdYz6emRF/l7uG5oEsbbMYdYwnUp+cTL3xuIacLJFv3OwSfkP8
5zjUAGxxiiiKVvX7zzPthD4YsNqOU3tqK+Kp764oSDQGBhBmVtAqOxPN1Yx1mvL5
X0/CXlEi4p6dBTe+TwHfGU6t61cH21aDfxSbktJxhVjCNcMLF3T08hIl/RkwJJRV
9JDyMFQuk5KvPFb+oBHbKLNFbZ3bs99eC3BjrrGTtjR/urdOfvo6it8HjoPqOW6O
W8Szma2hXvHtf1noJqjDDJww6sqjtRCA7hXqI5wiGoMmlo/jGncYX+CVK277nDRi
FMsb17AdfeBhSfWw3vDxQjOY5XkUH/d2zM+jlvDfjH++qtUwuZlqhQ8sMOrdw7Hx
Jn8Df8Dharvsd71xNh03c1e8OtTJ3NfZQ3rgtw+xoaNOeEwXKXV4I8whuzDz2iz6
n5dTXg3ni1chjjIBeRtl+fkAvuJmafGIbJB0grBELGMexDvdORavY+44IIr3Lxyf
CQiRO/Ng8azqcs7bgTiLKQXw6BlxJW5BqelupuwHkQKQPh9JGNJ0/szxAE7yV3rM
T/XWY4bOs/XVL0G1dEAfz7rZMixnUWPjVg0XxgpZ4z+GAwWdXeSNgKhBJSoburGa
+eSi8yUpJIrYhbKLSXpWGXKs4hWNUADV6D1/y+4xbR+UcCs1yZ/Ii57HEVVDI0ve
KS9VCPjTNDk1QrNfYSMbHEQiXDbhNtku2PCPsGHv13m4mszdmtMCsRSwxGt6vmV6
VF6POPXcBd17+0bVjNlVifKImfsXbIrlLx+H+w17gOwqD7K8WPDuxMMvcLKpEbd8
Ju7sGqjsznbSKo57qh8I/oXujUwJENrVr9xEffW/7EkPPdlw+ZiyQD3mVUASKlyj
746t8ZfOie6lhIn2n/8//JtKtG1ek6RHoKzPwlG+igMpgjBMg32FnKVl+l2SRN6n
167CDkFYisdcwVuBXAx0ytJziRQzUuWlisD7K5RA4wBxl5Q4AfNpyhR0MJGICndX
xvJFp8sqXRtMg7RVD95FhGISspSo/y28SMP6RISAe/V7Ub1q8Cq73qKxU94hd2Cc
Cam+6Dk+rs2mVCl/5R73AuYmRRHTc+AN18KUMOMCViD3+1Fszy+fMZH9NrJt2JFI
FgjJlupuejbHd1aw44hlrk3HEqQQ9eOS89M9lwcRIhC/59s5nVIlNY13iL7qmQ4A
lNDonuiawjG7C/wWOeucmPB0X8b4Tac0zcqZvTDP8eP1WWkSQszrYEaYTK1BrLOl
gF8AjOdtDuSEWGtjka4spolWS6GVRqUe5KBWpbN9y+LM1ferjyPaR0tie0gDacHL
lsbP/J5ZgaYgAjEDWkh3gv3BBTnHiAYVELUgFRrRwRMvTMHVNeKSbR++UozVRlCC
YmOTS3a+feyCYky+KrLhVgUoQXGtsBTXCZSwn/C0iCDgAY7DkLFqYaO0Z4xEuxW8
lRcKk6lWQT7p/zsn6zsMENw2zTFHzhcjyZfoP9d6Ca+vw6RsVNWRShVzj+BexeJq
pA+NDb72/C3WajIBUxg15KhjFCRyGNWbjSlqwOkqDwZb95SpaO57W+pWazsBTolH
ZJlNpWBdzZYRNw131zpwwCt4T2BLqd7Dvi46+pUWRJhOaFzhwq3aCRRS4T8p4hKz
3Y1hi89jpu+t9YdsvTihkwlhgO5QOPviMBAe5KbnySI6s2GkA04Afu0p4Flh4tt7
v8ZX+RmMiYOmQZJLi0Tj8230pz8sTNUbD0b0rtlxIF6iyaNS3m3BD/l2RSRTCwLC
5CsaFaq3KY4bUgScDAph4ccQ6PF8w4vrvAmRDbzKqy805FGqOeKBgO9sEGZ4wSV7
mnaNVpjlRrq7KbPtJLQiv1HWIciAbrXvwTGv0SaZAp8jSjMdMazM1A9u6LuoqCvG
bG8FBjWpbQN4d5zP57rhiwkbth/i6/Sld+RmNrtoi1H06MJTb2mAsZP0EQY1CONi
8MY2skeqwpWM6rT3wo9Ru+g8ol2bpIdWYFvb7YqQrSJnU2C9tGlvBz4bUNzTN1Mg
hkdj3mbNWMLkqjlrzLjRVx5NA+RSkYBqrsnGPD88jVcOnzBoWGzNiKB+s6uK9ODC
cIKIzZ/rncckBWKwStCKNw7JP3e3anuU+zcspCbW69JgnJLM0ggpZ/les7WAg4dh
//LQDYr/iiFylMAjqDaFeJ1777pzDJajFTxOhrcX35FdT1v+tdYqL8GkLHg6O+6r
R+BbruekyjsdVURgujxFg/PQm+CDRCqqml8lCYeOBg4gXptYpTBnXUOernxX8H/a
1C5K9nrGsrkw2DChWPgw8Kmaid/5X6PlJCrCSmsPBapCA7++Fm+FKc9hPVJz+Yud
YZLVBxI9zo0i4JR/g8WECNJV4ozv4m0n54pMr0h1RnjZNRSTa7m7HPErDAYQp48x
Zw8s4PBsHrOGkmpdin2/rygzsN0cFwlV6DZcrxdpeLDa+WF6YcI6tb1U8Cb+kqoT
2lDdj9UOl4qtGWi9xfEjo9KBa3sTHehflTxDg+ASaqLgZXkBQNuHVX/Ymxr+KjKp
o5j+vBTJHz4RTj8hxbIwTuU9UQ5f7pXv7bxd1iJjgVx0nEfgp3ulxUHZoV2exXfa
gNIxddLnJk+S8zXMZXZrHe2X5OW7r+6W+Y//p+6pOALYAgdg8d8SaA8+sKBUzkBc
Vxxk9dl8yaAHond0AsE8meRfBGkNz6kIMkA1PSYynQ4qnJzTzEPR0bbPzn75DLqd
+BCf+jUxcuOG6P3RraQ8B/oSgThLz7djoTdSdgzHuj/sBk+3K/OraDvYkaeHPZdr
kuVgRC9TcLBS8yKWC6PIsA5aTg+pm4Tmkg7VGaHyPWZMvIo6iwTCPQMKGzm2KgVJ
bAc1fyBqK1al2DH7ayZEVnZ4Rd2Lw6nuuI6clRX3YxxMW6zgSsSoIQQDX0nMY9H/
EvHkbTTqRiLdgSgV4VTTG0NxDl6bGNVEqVs9Hs3+68/1K1zjWLFlC8AQpzsytKod
4dpdDWO40TGVj1wAVJ0T+FQ0uRTLx+U5ozVBNamg95qw2X3gvCZpsfbeEaoGg6xw
/ToPnizgqalO+oaAb8cIo+XCjmPHVpFW8bozc4GR4s45V9ITiEbDK21EINbosO7n
Vb3XzHSKc7Tajvmv8QB+TyHN0bzAO6BiM1Mp67JGv+6qW9rhqqvyPUbrLxhXglag
4KTDeknLqFbgd4aDw/YY4WQXxgsmqVmtVXoS1t0W6Io87vdm6tJ7Z4rhxVCMxFsn
LPHeOuImXSboaoCNy+JkOCJ5bDPS/ZAekt2NXerzOkagMcsihpt2KnW7JpIZjyAO
AW8/4sszu9FnBUwJw1yo7uDSA2nbVasGZbDL4VY2ereOGIE0Qjh5ibr7YkkS6PGV
BPDq7du/RPUsf/QiHygEby3s5lB3uSKmKRnRhbI4DicCH75sGDdU7pN4ojBp73vg
/E7odPfIPYZ8bbLWHMba2fit1lO3YjUq5664j0tUIIMN07ZkMmJsV0Jc/aRL5Kwg
Q1tkvvfvD7d5AhEntSrDSrpW4/Y+4pj0XoqB5HrNfDXkQ/JPBK4JKWTReDCznLPp
cvONdOQmFu2NJX/QeoPCrx3Po6dWqHHia5j0SQ341M/B55d9323Mr41s7c2Chsph
phXpHTunlERnNsz4AsrGeLrSeiOvvTq3gpXHOjmJgsRZtYeKueVCMdU5D+/5S3J7
shj1df0DhOHhICYEiGn9yEgAtZpmXSlbns2b2GIlxElBW5goFH7MDXor1cDoMfML
ZQ3E+/9XGUm+M9dY/ZpvOGzmKdF6bHWa6xQyw3B2emKbHvJbXRqe3zBulpl7NtGa
HXkYOEYDs+/BaavRbuqjhJMeFpn35WAcBSCE3wKcorq10ZH/9IdSID+oo27hEpfh
abI2CetKTu9E3oI+ep5vXKLHwUwtYfzfgKS0b7CknkiXL+a/LnPo/oNSPxdsy37G
kMnzG4SMtVl33s5PIGVBhrPGBCJidKP8bzsgdysckl91ntPF7oy1XejEqPdHdoUQ
q5IJ11A1gWW7O4Co4KQ4EFHb/2kSjBz7NEsDJBjFvnFV+EDRNNKcWkwM+zZIIzE1
actYvqmK0N8u15IXKWAqpzzupp+r57uo19Yv7lOsyyDqMd5muve3OvgghEgnL+5g
WGkXuWGWOVTDjMBFR5rUKITbZyX9mne8uOgbY8Xe677FpI5i0okoTuxX8qFHxvqD
GsaYhiNbkdwuxS6SgUKnqmvTw+6zWG2XNhRJxG/tJWj8p5nlpNa7TlQ3xScEa42y
q5+tZtwgjhS70equSCUf6EhgPwfkphlNXk7f3ZyqGb1Xr8WH5piulEVQqHIcBvdo
LXNun1y9raF2lUbJ4ckpmlIKYSnuw8kPMVaYYTS3W0anfBP+5hgYCmTBjniCnGJj
AJufyXc7NmxfyflRxIjpiH/ZbWm6Ej+Y2ZXTs8nhO1/he3cr3NulXaVlMgdP68LV
5kGKrHRP8YxH9uEji+rP5Xv0Syvq2IzWHpdexuF/jr16BMfHx/uE0z1ShY4ISTOD
aFJcfrJ2U58p2icoMcPOt82NVsiy1mnHSYkZUHfVyyAIqUt0GzovgF7j6GtVIVb2
82Tpl0nXnqDSx56XXu+RBaMSWTIxOAunxePJkgBCdkGcm5H1maEys9da+c6lnpUE
gYuxGxUJENx+ZZXo++QHPtiNZ8/Cf+Zl8KSajHRwtEhUl0V6K30pkyCuvTveJpxU
7EiGXGrRpePUJBCPRmQqcSd0/jGkVoo6SRTiHpgIqa+qRsgusEI0gfIzZUjO0huX
VUW077SY7hS7+VCPquXHlWrTAUhbngFwEKuAabqdgi7V5SeGkfyj7hLTHIQfzkEO
Uhs75qmJoDt3uRSYFp+vl3/m+KgWiP1HgGJSKm1F4dYlgFIwfO0ptjzVJZ4U7tM2
JSdHfiDPPjtMuPE07QgnJyLSMsU8nvkr48dikVbOVSdU+n/XsPakQElN/NdKiqIg
xkETw69yoYSLGF/EqRdrUfAyDAc8Hl2TYncNSio58AYGtKZYnKy0H4IQ31ha3fMl
kd1DJGXdGg2bRNA4rfn8LktNxZPUdj8oT3DWLHE7fHLqgGhLcEKd15BPVwk2hvDZ
hdQiAc+buMuPHyqXjEkhRpInneg50s3hseWpy7fPhBbM8j6wJTORlcN4Rs69WcPs
jsDrgjjhS/Sgpt9Qm3mWUKB+tAbnOlthGNaN6JxluopUDMIo8SvjWiXacZ7K9zHn
O+dtF837XYNayyDRvguMJ0nSV5fcwecr4b0McL5HjLee4swcurwhWVgfMx10Bd4m
gyqeRCsVwGvIgSgqvOHTW05FhV3DGT8lAh3Z74oRsZYcaZ3FY4NcBCwnGmh+rjC1
y9QTMY29WvigDLebpo/Wr6PS9IDQfIBjOCCHyDcgEHdwhF1xNcAYTVYzGvUJ8BtH
kJTVK9ksTYKGcgvAJWyiEL6+WuP5qDErUv5chX5lkaJ1En1vesGT+JUFfpfmPwj4
81L/WFnTvgsCnxy8xv3VLmpPnEbNqD0N63VRKIh3wj9ihNzxvoHx2cdpsaaHe3mZ
wuG44pxcu51Bt+rwgg+MYrYzH3NKweNHWg+PCCE+jFWE7GLShx9Dwq92guOIX7VI
odnR1FHOieUOAG8NEIMWhfx/yI5nkyrMvohvJ3MoxQTlZFBipb5RscV/tmgutbcn
PvPML43o20T4SaYWrEFez5wNIt2Dsrajlq8HAFQBgCBUCkfQN5OxmDGYCdX9ofsR
pOF6o958FIh2WpsifpxcLnvlEILRCM7Z5wJMUHFxMZTXNhuB9xxKIKwReEGioSpt
1MygnFJI0o8sbkD4zWyIkvVvi1E86+ghxEpZZIiMTPVAHasN1FQvGz6vqI6S75ol
l7B8sQEtYVNWFwtX1E+mOUCcGmJiCYXM0G1equSxk6ijt/Niwhy61mSZgt9Wn4ug
puY1cFaHwtiY91jt+r88ostcmsFvg1PaXGuAgdupaUZSGD/G/EtDNEKYv0LtXMcx
Gj8FZSpWGhFOY0wOi7W8V1loc4Y8e8Oy9b9/IiqTPziQGLJ9MNK+3hXfG1O7zZjC
IRhgjkFhEXXKe2OgoJBiwGCudpZQZ0JMlIMkjd2A/8HbVfcw3t2uLeacG/6hNfuh
7ZvLdurwTIcQVmwYX1jNkYb/KMzg9uzmnviS2Ur4vDFsRcaAfWTW+sZPKHHetDpy
4XoFc+HJFUOX9I9XSXXOa02IGma573bJUrRprOqBn8CGbx+nV5pLkeggHgYuJ4Yu
yonlmpGsmmN2pKwmjXATqf4DoNpAzyeX56orBwCayL9Qg2ArCzep+uLw8VLAhwAO
8n8YMuwbxR5Ppd9sIW/abWrWm6K2mAnK3sUPUVctne8tJxv0YRjrpA2y4QspJF7z
NiXkiAtY6GTJYE3simGD2TkupiI9fA6Vaw+eCgNHLxpHQBEZRLzSTYl8DDJihmIX
z5IwByU2Q8wfTIbKYXoGNgbwXDeeK3wlC2zfptzWwuRLafkh1e5370L5oXG3Vnx+
4Ginv+r24mJhG1SqAbJ4iHAELta2TloD0mEVX1ouWLYDMW5OrYStjLBaG8SiQnZg
z6qZxt5zvV3k03rJ1Ck4GWYr42UrdVXP021+oJ6b3JZ0LfXo1nQKHf0H38av6RtW
Q5CZa7BlXVYr8Lf3TFhsvXq85H1PkGQSzlZ74vBo6a0zRBw0cP1FkcDzRaI+hPpZ
Qt8neRhK4s4Xe8wmqsOWmsrIjxDlQwQvY4/ChB3LL6av17fHt6VyMS4RbwrK/t83
/LhqHqwIWa9e3FqO0qzUseLYW8C1kIEUNoV4DkLCrW+rRvTtuZ7Hia7uKLtlwzge
weepfrUyPKpjLVLMIokfBm8WjoI/7sOBtiD5PpvEH2Eft3qQaxwkdok+KN2WsNJ4
gI7G2zce21PNLdNTjn1PIxg6TZ8Av/8eDm/clwXhFbyZvJ4x+Uvoyeq6tK3V7Iub
jJi/Q0nFrRbNCLG3CH9EGDwaAKYl33b0n94OhC/SaPUjqtvOcvrOLnrWLw34+CvH
HCr2BsRw5EI8KPHHuHdUdpEkPLq3M3rD8gHMKKRIXJ67qzWbBUFV6nG7zsZ+2mi0
j+WQSd2UQBC/JXOOeP+AT8xlwYKQ/NKsRpwyjqjkAoCtlfzYhYf0ec5zHzkuKCov
35iBab93bxMqsei+wSfGvwSJYA55Rn/IZv7HNeRtJfTqOt3naRstE1WVYtIxmM/h
ku3XAG5huy/LD/S3YsSNoz6ECiQARdukxOTxaY1b6DUJAlJrFlkl7yFu1cp9wEeV
wf3/oihB+ktmOlOn5hwEjrVxEEI0jzYz6Q0jYbp3nzUP0MO9o1I0smJmlnrM0f1T
+ZLWcLoJdDHfBne/wERMQdRtc2NSegwTMJNsRhwnpKUNes8j6YsuyLV1ChjaepSJ
hDA4PpKIV3rThhmtSIJhV5Qq5aCVumBdD1ftkRJZixgNjiNr/EmzRwjgo0KBfB4x
A2nUdwTkworcQVlBf3SIeu6JMo7OlkQLhro4FLopXgdz6h3IzF+y8jhs+xbbrZ/a
Ubfj7G9gBukrfx5i3AgM6cDdIgOpsMjhQm8Pisf4T4z88fOHerIV75m5kwnkvNvi
CFGgsofeu1+U2px/dRXRRJmn+49KkJEPXyql0IYwkhM1vwS5Tiu3CSB3ONIanrhC
bCblRPTVow6FzJbHdhHWKcTUQvlQ7ULMU0O7Ho3WFWWQZ2JjcpTgS/T7AuVHT5sZ
pol6semP4G7LuBSR1F5Bd2DiQ9giWwyZyFeEnNCi7OdMPMDhx7YBv1xR6caEegy6
Ttk5x4gyPvXS2SnmF0JrDNmeOk/JbdwL1gu8ge+WYCFoNztH4XCxuhDjkji8E9Sg
YJAKyPyl74vII2Vg7v3FnCyLGKCNvjQhCLEgnQXBLcfjdATaGVI0CY0u+QE6T0J7
gQNOTkA0uZ7Gr/ngKv5Uxl5GgvQXsonis24ShuqpStVk85B178iY5nEeIEWnfFPt
VpZmnDRg4+cD5QIdLTKjPgVTpiogypP5wD9EwziC11fK8kPGiv1pEv4qckmlrUl5
bPTUMVrZ66NmX2F3MRQwHxU9EvYFGn/GTXuM+YD1W5dKSpUSyM5W3+d/jKhYf3TA
t6ILbRg01t8b793E4YYQz73cZ5v4R4n5zM3KgVbQMrzTnMZa+x2BuyPObdqKZzDq
nHDaWnO3316jWcocTIsNQ7XKPUWUOKvj97iyybNzXrSQg4TnpCLe28Y4WYqN+LX9
f+pfwlDsD06xE2niqUwWRYkrZKwlWQ+kyzpigi/bCBpD4CQKEW3cZr0Bi6+y6CQT
p5Oqexg0A8ttf/aC1um2uHZszfZk3Amm4DrF3Ah785ykgjPIrBVtNlYKrSHgBIOL
rkB4SuBuHjFLYiDUfGtWZElGqINsU3c60VCLbuXklZyVF4sP3s042wNJMEWyi+cV
IyInCRM6oi7Bj95cdKeMQEILA6V+RSFG+su6xqiie1km6UkfHfaMZjdkIk0sNmYJ
II+OnYIWkL8UYMXSB2eKfde7/jyuqTtUMXOYW4L6LlucTB7gP0FmM3NcPYVf3vyi
C8uRe7NsE6iLDQfOrBru7Q+jCHcMosLDH6aSKO33huExEMFf0FpF1ECNUMK5DTHZ
fy9tBHhgFzeF+d8rF1acrgGcws8vUtpGMs7UlWx6wzq17wg7Gf1x+UML+gPDxX6q
eqBG96MMZCY9tdBeLgZuAwzQzaApVpx3Son+vg7TktVXo/2Wfz6qqyU4CgS1vR1v
gzQIo/TsJ9dIDRLys5qqBqc4hBvR3izrTZs2me4p/IhA8IO3FDRYSCmOwK6XGJ4p
xL8o+YyGwPNdxT3ZDLNcGIVevDBrixx63koTnLhGkYZUEVFKg9SsjuGZmAt2rsyn
GAV300n/JMKIkL78ut2DTxxu0q7VcljKZAlhzczkQEYFeCojGNfvjFd7ID4ighbQ
D0jTE1qq5qpzTAEgzHMTgik2sfx1pvV6YZZ7dGoBoFy99s6MJhz8X18eqi25OJE6
Jm6RySBJvMNFu5mlG0SdkLqbtKWllviDjWXzgErkf92+QijWd7+Sq3xJvNiIq+0m
sdylDorGm9z7wum15NihRML/ZnjuBGTE9PNd9yloJhiZxlUk1QHohR9YAiwp4tGm
AAjrvOb1VUZAjXB7Mo2u6tkUv6BjHOYeycpj4i5s7CMF7QvV4WzyslWKHj9pUm+J
qALGDvRX226PKhNoHSify42HLX4/dA8daE7WQHGtRS7Cx37iDb/P2r7cD8G/Y23v
7GJ13TITjUFYO8Izw0JgWDZUmXbm4kKo8boX0ZkikvqPpXCwGYr2KYr9n2XA+0G+
ZCPoXDFwUlixDhXhyLX5W8R+Qn9mLLqkIlwQxejUrXWyLgSiNRKPTaEmvFTq+YdX
aYkb2a84v2DBOserfMl++0+NrcpE51Qsew9dJpekcjXAD9Ue9me2dQS7WP946KTf
iQNtKL1fnXf1x8QwMVUi5AY1kiDhttCAuhaF3iwBBuMeOE3vjDeyHCkgWAZLcvSt
ualwiqq7nbE7lpesx2YUWfNZy3YaI+CuO0NLppy//eAX9SGopmn5RD15sIaitR8j
yFCljGkTOd7EW/QRrYiT9x/0j74QGVQBHtKQJuzduvRIdf8OkgZC60RQdqf7+lFq
Mz323SJ3O3g7bqZBuAQh8JkDddDm/gVfk2Xfg5Sz5PYnlMbz1hgOv4aYWsO4FewA
QyZsVY6J1qmPKrvpukc30zQ+c03Cggnwx1waYrDgda1RfRXOj0ahvISB2i3T3Vo2
Lr0k6Ei0MkF+0DKACVt2zXHTjB3DGTEGvXYE42XTVk87DOGlRdNIgvs70o/sNzwR
gHKHO61lAYGf7ylFn/3aOWXVr39R4RWiFfqaV4WQ40SG3IZqANbUsRfqnd1eY7G6
Fxwa8MBC88NTfsjAIJHVXYElUAVlsmSaZvzRcDnaFEB4lGdr24mlszGIHyESPw7x
Gmfx9TphGxjSPp9o4bUw5xFtQpidCAmTpL6ea4x0GGfotaEUUEj7r8fWcz7Wvtrx
BFqBQykJRKpUw15JRIrYvK6XoLcv21x3eHmmWKdg6VFe70VYotEy1raRmAHVNcnM
vzTiQzv8l4+RVWMg8lWWMgopgrmtIjEuEeKEviHKH29qPre3mqd70Ze3R65vHxcU
6SNyMQb1hex2j16WTuQXI+u6kmIuB0+4ObdtrRAQaBlr3M6MQSYA9hHxGa7qabyI
XwqcgCpEf9WE/rZnZtNX70vXbJ4av7TQgLFTAKQd5P3jVMA57W/8M80r1QBR8n72
3Zeq9P5FpXueb1W9Wh2yUdkZt2PewNl7FIRbuh41jj2ktCm3hj7AuGUXZHk1qkvS
uD++mpVmPLH+1y79UOUy1GzMl/BVDcCHDs/nbWOny7uGSs7/zgeITAdM9FS04Nvy
vJMb5sLxGTiyGeKeL1PNTtcRMsb1vyr1qAFeg8sMk+Zpkmh8n1lvs0Txmyn0rTO0
C4tvEoin01f9jybWLtk/JWT+TiID+AW5419/RAVCt86WncOlLVTnUaxhj7z8rcVa
r8Upr82qTSAPat7zwgbH4bbbPfixDe8S/5oSnrhLL/rwetuMJ2MiGrX3/5TCItj3
R+STO9b3KCD6h3A2l02+z/8jSZ5RTwRk683BBKIOIpjzc7LWtuVAmYAs3w9xaufk
v3b3BPOIM5ibX1Q9U6V4HnJEZj1yw2F8yoa9hkynALFWpZTZrCTxNytyjhR+zOpJ
69C18YB65OErZvE1Nx+zbR4+Mqo9zOwfnw0EIIkYBENoDZrzGyVHqjNee/7AVAzM
jNqoXRZctd3bKklK4AUyttMcxhmgN29kqFP8G8G1Upvfz8K7/weI6TUtiB0/bk5z
K1Zq9KSxmyGls4pYCD7Rk2hb+/ZKwpqIVTzeCZDY1rbMsl4gWHWN1Atjl5P61Xge
dkm3wvJhUKFPmHSltZ1GvmQ2jScxFnx5ydJ0oYElmKWd5FgYtpQB+79crcXqgajr
yjCO0cgPZHD1eg2GHvOl3YkCOJe8sVSQc80kO0074Wg6Jf+SzYBrqBHXZ0uTTsZs
NsqZiU0WRMiDOHWbA7MkaR1ZI+9HgVAbd47sj5zAC29bGTox5wme5UMuem24pgXH
qu87lldxqj1pULLTLzQ7GB8ryebH1YOgyLXTP73VtxMiXx/S9IyiAvwvZDbp4Lz4
va8K+YfV0rAYax8Oadhk2EgO7UcwF8I+iQ5gyHPjJi6iXJY5oEuHkgQjXgBj1Ga7
MW6Xlu2siMH28lsY0Wuln1Bp8oX8RpLhNP6G5WEh3BHld0bP9yb2R+AAiJ3+JpL/
OfTeBtmDKzP6kShJg+DtkivKKCQeeSOOuXzPIC3+3G21exQlyAA+0mbROHIMtch9
JYIbtYQJWur0Nepp2UEOdzo+w0vKUO1OBfiGrlnLGFEorWybXyeEijL3Zu7Rt9P9
GIFqIGiiwkEE9sFCDv7BmQs1jSiknoTrN1ZLWCvp/pSH4xrqhBpxJXbrV649kIBx
rjCeqJkD259TQQlRhKvdaiyD7uPxjfryGqhdQCirHltxHesWK+4bCQVqCLQ7VM39
rVtyp/u++lb7VFSYzSewDlBKprtmZJuweGzs1T2ugWHh6NaFXjWzaRVX2/r/o5O9
n9v1F+3lLCsY+7TX3/2AamrOrT25rGEdNI18zav8r8QJ/OERe+K0ezIXImexW/lP
7puO8bpwuAi+TicqxEx9NeEpKgUFfFnW7koVN17uk8m1MUtxU/LX72hwPI6Qji6N
ZjaSBSJOUqt8Xk55xVO84k/gWkmQUluegy9hHIvLMXpokbfYkO/6/ilztByE9A9k
Q5lEMEpuyEpwcslQtP6nzKnHvqrQjQwkGyDN8nNX3MnBorB8X9/8ryLWSWlS0PXM
8TBBtKTGuJfO7gYRenQe2hJlYyEw8cZKis1GNi0htJ/MVh1a1ZXoQTZk2YYkxaBK
WdJmBGXVVyKBB7iCEam/LBuZ6f7vUUvMDZFx/1Qq4o5ba0jMajV9G1h1ZIRUQCyA
h9k1uDjU7pVwr/BRm2hlHWsHjB18BTRFogjmC2FJhKv3ig5Ehmvvls+YKdn6YEJk
q83twVjJCPlT4fuHAHoozA2Nun5FckB/VJUyyP90wLRMUZfgWrqOmD3u2mFgS2SW
Yjduf+pC/nRWmtHEqLzGYPHg5prVpL8iSw0sxDaygnqScPTeBFGpRKoSufEdF4jK
AehLO2szB5y+HS6HMj6reZLwJoBdWX7AMLA6vo/f13VqK34RlsKb8uVa8QNpbOEx
aDT5IqTihSsfy/P6wTtGMBBzxkQ3MN3w2TteGJbF7YlxhlTET+IjjMzd5tdDE0yv
Ydc0ipw2xKMeFZ3W1nC20gPcIpWNuY7jUgBl8UErijPxcWkmwSU7629IhInenT34
iAjc9nON4Tg3Vr1rsHRHfLR91RsHZYi8iZDItKTjnbval6RuW9WG2wR+NWcLxv97
pm7sr1ebvYlqjlL05Hm2lfHG319r0DZJ+APE0YoxmIcgK9ryqIjAiA/baeg2zgc9
fNw1rB1HrBCtRWlMj262QSvoeE3Bi5lgkWe/SnCp73d5NFFrIn6dQpzuAfoQuaZZ
KvzyhjXqpKKJodPsL/UaBeOxtCV+mldbGK3uaHF0z0Hk6G57btESRBEjg6GjJEKP
oh2anNE/h9Eo2xeBPNWqeXkXZZb53MaguQEC19164EKpyxmRsrCY5oywU0ZF9X57
ogAcYpvz/+wMykL97sq+Y1tj1DEyPGzUaCqL29pTKUdM5GYdUrlj8aU9B5pX7RQa
utMr9qs7ulZrPPHw5dnAL+sv4fa0TS5GsaxTKcIe7CXKdIut8XgvLo1XjyymJHY7
STnDhNzBbe9IaQpWh99jcTTYE3+3yeCPw/P5wUaDFRslsPVqdjO4g35hsbGXdCaO
X5R3FF+L+nvSpFGhF6ez6yzP6jq0N00w95lXW6mNeOVaF9HjZRVMMIvN8qcsuSXY
gvLUVghCwFzokMrLdMV7S8osM1w26a+EcHejiVUczyMXuLmLJHvt3zwS+W31+wSL
+7i7QbO1G3BHr9gqp//NWme9iPq5BWLL1hKbpTYmGJabCictq7Mx34wR/cZE0FiH
xXc4WSTsYN4V511pJEVdN28B4YgLxzhMLNRC0ofeAdjItooe3MfeqWun9/NMctA/
wXTqARUM00RMFKG0EEt8LSAKYIS1cupmFF5G/4iOyRAanevsInymoHmdISuANulD
Rl2CtoQcbtM6UUiXRjDMFi0V8Cn24lJjp6ZzIeXNA2C4Lye3prZvujfxMgVZFMHM
urKnvvrjZvBwzVwOjAMn7OCmE0ps+D5to0iEafY/udy9S6hgZWNe8WdlsTHOAZDc
YaaJtgkKszY3SYfuwF8hHxvkJwTcJuMluul3CXG8yMS49bQ7i2Pt/iRMHh7ElUs0
q92Ii0+nDKrzQa7Bkc+ioFcr3ZnZ5lQORIxhSMIIM5l+csckCxb3+1tAiUsO5sZk
0lV7S4s4+jgC1hsbZT4bI0N+AYDEExoGUeSRBJ2yHEYFa1E5dK19XJ0r9FxP+l6E
h8K0tq4YHjWK8CsRrckZrDzQKzJtKJIcUBBH8PPFvnKTsZf7c+CjZXLM9HPDiQ5g
rXeldE/xjNIBAknhptJ3jxrqbaVw3Vvt8xeHa9pWXvbG5LEGCi09sWyD9zyx9TCE
v2mBGM9g42wbOG6UccHO2j7lPDnZw+k5jj+kZEAD21lTFQqXHKieUtQV1vhqHuoy
GxuF8gxX/KwmsI6VFB8l75ii+CY0dp6T0h0HgK8kuOXSgkuiyL91LxTh46SQDn/7
WDB03fm4agJjpaHar73xuTgHisCgnxczbMt2duX33AE7VOR7rHVA2TJA7ZxKeOMu
IVht1D0cMP+C4qZoWI6CRhODpvvvRVDbtdUAdjgFK8w0/ixtKgV5Zgh7d9I2+keU
axbsSGywYQtaeZ11cniZUj+Fw/jPKwO/BQJ5KeQpycWgciET2qNQxDbuggr0t+Vf
r/2HJiN1RhwhbD7zOXs2PHmVMiW6F/0ZnDVmlJu1rwKp6RwTufOLcz2fbqS2rHfx
vI4ZgA5L6YcLzvZvsAX/xxGWlRHAhIFU9CpUV/eVNw3Ira+Vlcl+S2yZowAOkTmo
/V4FxvuI1R/oyWMC0O2O3jXDeGM6/Qzj/4Lva9ERrAm8iBW6+KaIbTDMFypQhk4E
UF00LHnkYBA0y/5lq+PVUCTFO9/b55PCHvIr+tColUtc7BuaSZfDCX0oxgaoyWqP
GP41hqHfzbALWoHG86rQ3V5GxSWn3+buOGsPqeh91vvX/lVFiteX8WdYemBzq0ug
v+1FitAuQZ9sL5ITEPd6B5+5IAvSyVf7mLUVfkmQtEdNhGCn9sMIWggKO5XnOZ+G
Hqcep+HUKoygp5zKtv1zdalQIPL6Zg/ryBa0Qg2YBakNT9jV7s+5UVVsrkFjSyfL
E/8xAzXBRXcYtMUunRZKYmPrdfP+Lv+AsQd5jHQRLM2vTtmvSVldbXHCcBxef4MY
0vSI2xXSJvLV/YmBivW3pajdEUG+Eex2GydYF1BiGiiXF1V/tWZe0iHr6YFwDegW
I10ylygaYYfK2eSoBbb0r8DcKSd8k1GpdC7rC63zchdzTBJvaJ2fZO/7TX+fL/1V
J3Ghsksg0lIigThVXqmM6vPbGA8zO9ois37KDhIs8esIL6dxyI4XrkwyljGSxLKL
ur2OZEbF3Yz3gSzcKVKgQPnr8gprI5Q4cJzLRl5mTFdtMgY5fk/tMUgLZOUPz9Xi
G8k4GMQhfIkGuAF2z226ir+nW7BtvEtNPUjYhhFQIL9A8tmoa3bCX3rb7P4Dp8jJ
cWbiKaAsICKsPCnexaOEfnagmMQNGZJodUFUnLbl8ooOsKk7B5Tll3DPcTNaNjHp
fEj9qPWmM3UgMlpt3o9wCFvDMs8OHkXA47qVd/KbMS+UqXN3BLsWu/toS/Pn2i19
1OE7tsgA0Gt7qvc+F7AP66W4kP4nyze0BeH40bUp7kPQ8SzUmceJjKURR6lgZyMO
RzC7zdrKoBWFHry6iV5VCsF37qMROV+uVT6rC9IYbogLSLYsNbHJb/Qxr1lvHsf4
YD4/APHu53jNZgzKFDO9HXgkTrjTyVDmucBLyx+Edm/opSZx+4pvOMrP3i4hOD7R
CYG7gpFjoe02O/YTNxMwV9uae1c8+wkUlEt1TrPycXKjpejH8cln0EisRKEOrhBF
GbqAXn4w+LPoAA0vRwirjw8FWEX4CMfxD1DJiAu5eUT8BeUrKa3hTg+h4UEdrqoL
NAmjnHtF5+8cD6fJOEN0BD15AFO315udTJar5qO68175JJMaRnB3jAltXNcu8kP7
F5dGK5aeLIBwX0j/TTGXGO3fET4x9uTfF37ulDOmjPlnESVa9Nc+UDn5DyHSQMxt
2vAj52TdKjm7P0ddbcqEOftFg34lnhXr2OUft36XO/vau1gRnQeuAunXjMOVwgd4
wwExd2tZP6L2Pn2SaL+2FNJ8zHEGQoVLicdNKCNjR5uySxNYwbKttfHtaU4bfKeN
Tax1u8owMUFYew4QEp49YO8rqtjdIzf9CEChaq8g3xBmJpyOcGeWQu3JyajYI+kg
+auctmzT8dMD5QAetZME6YqLuzgpI6bF/YsBXkZVgc9OypYJjHmJdqg+ScJ222qG
r1k6DOhZzL4haHBBZrG4s5QsVUKwYfHq82iHLASnUSqEG8j1LbWihX3e+Ybs6FDT
1pHLwFX7E8+chNg7JJLOgSRc0EzY+aFkHoDEe30hjujV6euIwRH7Yh53qlBK/mSZ
2esVQ4POPqxYVeQXim0ZX7voMrQ2qxNaevvD7NlLmfvoyL6jKwtGOAMDHPSHnSoo
hndnv023of1WdavaB/9zgvUnvfXYEJyLL3wfKeyqNhkbunxJsNQ4I4W52W4WxfBo
Q9m+WTU92P9CnBqU6WlW182RUHJNvEDisHJvKe1h9eENzcCaC9E/wMZvtMvMGGwR
uqRwaya9wnIDs5cd5GWeG7GVCCKceZfNr3TvlI6Wr+4MJrPVDF1M+uZyfZv87W1p
k5XL19Nx+4CmseONuxV8nyOnqaqtuY0BdfdPq6jyk9heYdO39K1EQHlQrvZzRhA1
6C0IuEQJVfgffK/fvcaJIR2c3vCXgr52sutNuZFsxgSDCjtwMk/GjxQSqEzJjhZ9
98+5WPnWELIhQdZq7ah3lRx2A0eLd7RWtzJLRLffEhSfvQuUHfI2K772kzAk1IH/
LiZw+TRiOrN5JqdDRfTNSv5IU+QvXrtUfH+sRL24iCMpVquyMbcBGIOcSZqxM1VG
9RJdgLQVH7NABasYCvBpLBIb2jenU1+YvnXQ16uZDjWf5GWIAPMPrQtaVBVRP++D
q6ricxIK6gU27PIvoCj/K+5BRAGrMP87fhmomghLHmh1gSBJH0F4OogxewYWi3Vq
bQ6MF35v7T+08sfy08AK9GzCsqqF7nIO3Wvwi5X+BJNwggw2nyPTs+y+a3NOMj3a
+doja7X8zrTw80zopmm0s7+xN+IrUCcRC3xc1YjwI10+4uSbCkUGI2PWtyQLZnqf
D15b2/PGKvJ8VKroU/9B923k5mWuZ8lyKVv6ukb2DKktGkdmZz/0E7SkSWnOvg4+
3HMOty6eZNb3xtS6LBPhNL6LqxVFMop0YHLKNaZ+PS7cNVxiDirRgu5PSjhMx5e4
d9oGKA19SLmLuJFxypWFEo1WUhvCVtTB+sXi5mvNrqZ7eRfjqh9iXpLoK8k91NJK
PcBpUQ7l7sNUsEAZ7aKeyvUqg4+Ch9PKnNTTP+R218XjcbC512d4BOd6cSu3eiVi
qeLZc8a2y3KZ9ByjUgq1V+OWfixURgBupyvGJazaalGkYa2pL0fPcy5Z3JHE4aDZ
s1aqlvyuoPanoyMLy9JWTk2j3EsSU21fcZvZ2ee2vnfIc+GGsQ/Vzi56jJhHlMA8
CkSteLL+x8RM5mdDqN3xOfiDp+F/NXaVZ9/iczeC/Hpx9B6dRMp8oh2CI+9Uf1Mz
GMLIngJbIPHLlX33njzVBtJBh7Ec+10pcqMx+c/jLPElvCUKXJ5DJQ5Dyc3qgjOR
id0yvgLeqZXc7muEOTia5hxRr8VyX0HbZY7aSqpE2wa9b7ayN7DmnWodeXAtidlj
Unog+vHng2EMeQ4aUBRFCoCVcUA2qXubggCn/qxczj316UA3kCJRzUXu/M+/Dkkn
/FmXlYXERspPy82GSXVBLBkqagJo7JTV8QdDU97rm+XbGyutjD6v6wNuwnuJrOyH
U4Bn8R43h3Cqy3YRPvB5Z0+k8fYnc5ZIs1GyuTZlPdpIt9oUJ+/iJy7P2BWLdUXz
MjVi8Nw5vqmfx0pybj9ugrlyGevrnbsxIf0t1HNKojC/CkDdndXJhH/kq91I8DPx
eIuvWvW1KtJiT/VPrNn33XQ96K7QnSdtN9Z9L6Lr+ulE8oPe7gAp1YwUo8p9mzAK
YhcJip/NgwG5am0AK0Z/5+Gp6MTgTjnbMcsev0IFP0Zlz2QqwKcOMRlYmPrjQOMg
83DmJxVHbbqUi4S6HvI9/CItet/Adkx7kVCkqDbhO3Ib+eZx9r2GL+tdZV8DVaZ9
gdxfmmc64Nxk1U8O+6RQzi+XOCPZC0tjAzsKAkF0UmzMj7tvHIO2dYDZLAE6gQ/l
gC7lBOudEO25IhsCEdrBb6g0A8D/Tk38IWNIzdkp8HKoOgnSmr5RSZ1Gi5kow25B
if3uokhjXOd5+/C3n/BWZOdo/WbmxoENuOVeVr4RodUp3q630BiHOI442/calgrs
FGuANjswsgs2lbqybrnUH7x93Tvn1wNt0Nh11NHwFBW9nxcbmKzIOPMmsOfla5Kg
1LEENW06TPi8y2IBtTONMmbfKlGHljD2DYHQwjGtqe53Bv/pUZHyQ9MVJO4KO3wK
DQ78teIdVPqKHNJ+fdrFuSpsugUBIoRvw7RbHzv4YzWZ/E8RZEc3LqAOixWU5isj
WeZtYmUx7GWsLwi+tbZ90Od6J2/orFtHenNRzeFPW30SDwmpZfqDPLYSypBh/kst
EHJF7Dydau5zCOBcJf66PENkFsqF/HBMX3FW3F52x/Zf/nr9I4OMjlCT5CyJ85Mz
xPs/30O8WfAAqrfFT9jJWl7ya+4jCBCTWqR6YwqLmB+1C5zY21bL8I3QMhQp4RNs
ek+azc+9PvqsOqh2JcwtY+07JYAfVMcbx3SoiJR2ZbroE/c4n8Emr2TOtggk94XP
ZoqoPZXR7StiOgX7dJ+38EujpAqHlKWiME5uGzMXpGw3AU9SFlmPzkvevlIe8DaB
DDqNqgTjknl8P7Myxxw/y8H4b+pcxaERlIX3Bdh+mcG+mBvZB58qgy6uzo9UngY2
+OUH1q9cWDK2g3KmzSz7cs3hzrjSsZhhZ99wATnDZb9Zd1eW1+mSaSYowF8sNEWn
T364ea04ISrkDrdNasvAs3jZ1lCStCfy28aJLHeqlFF3fXYjc40GJAq96edKszaE
ifeQrdPxALoiVFMXAO3B1d7rNrO4A7GHbn8Zv4B62SWXzGLBhzlXsbprdRD6XT6L
FfDL+Oa99CUNcLuPeGuZ/bRYbvAMZFSk24d97u+osM1wXPmjd8c5rgjHjWvKXJHE
PDJ0DsG9nfhC4LSAbPKWq7tJIRGHNHco35C3zu9QoPQx22QbbA4oYn4ZIJvCiZil
YlY0ePpOxICioUWJF/xxzF7blxzOGwi8SqWxspFQ+a1EPLPeAVTon93uDAyHGrqB
1LXTugALGI0R8oZJRX4EluJyX08zqCFyIb4aVhnG61t71xjUzmMa08dkLD5IxeLx
4SPiWxjdO0QL68UVhptfKkuioSw5o2XtB0NzCB6RSmFRNDstatGbl1kXvUE9nwz7
MuX8LNFiwFpzi0w+2NcARizVgiRrYPOvZ3Ej+iMoKklFxcutmVqJ9fDojoyQDl0g
inuhn0A1YqqOOzGs8bNNXhvkUl5oSdFXblVpg7GkxIk3jR+yJge7v57WvGZ/ETpa
R/GLbWDmuWY7wsc4vi415Xx5X0wc2L7W0F6Ac1hPekzpzBhMGNFBL2dE9QUrIKBK
PT3AvCQWKN4eYo1oyO8dOcfqc9qMiQh6jpGHxoidi+03qtsh31iTV5YSkOeS9nq2
GRI7UDHCO0ArstuPcXFJbV5YV1k4zDLE63IHRmTV4nulELB57/s1B87b7Mb0ZLtr
ceX9fJATJEdyhaYHVjdX+oRdFkM7G3IUKj4LgV92weSgvzFQZFXpPfyCNcnjFrxp
cjOcAoqDIazkFslOcfEglwiZtUbaap3UUpApVUg6Y8P7mUQzglSRyIeVyDH5C7FV
5KsS6WbBF6pvu8i/kIvbPNxvH9setKqCWYGDnDuCjrOkMGF8Z1hJXb2komt0lnSZ
swc7mvn7ZfZeUgWf3KeY4k0KEJ9fkdDgi2lgUPpeA4r/pFHbjBGArP4VYVIMgPzQ
sOFoLzQhvXFVNHnwJxLhWwgkBlnpQ7ES9OGgaSlVG1LZH+/JP7EjKhg2dlMq5/wG
cFKL9PLjPq/9Ap6eBWbaVxidHMVtnzXeOV7fpTySY8ikUb46/jgUIA5rD91wSZ7W
m+C6DLWBB9h36TV8dbq8qERxD+JBg2FvsaVcLzC1XpbJrmgYqT/s/vGVFy8CLoDw
FcDZEapBXaObsfWWlpmRVY0ff7KThcV3CkorDOLAmT7ct+cMpsZ98mctVevZ33Mr
xitMykMSSss74ESfa5U73KdVrlcQsWsOm4krYeG6oa77BP/tvLp7Gu5et1AXylMe
0XXwEQdSQfGiR4UOKrfhSJ1OFfXIRbCjNGDqPP3B/rhB6TQD8hFw6a4YhnqG7BIu
DK7gvBjTHHbXFnF99FoJ14HNJ9XB4EfZ3H5JZgynFVxO5wXu8pddmjsctsqXq9FY
AXU4gwiZuBk2CntBXJYTImEd+6yapEM9n5WjU2BAzcPWbJSgqXR68cxeFGWcqKhx
Vt0iUbAYJgGvnDLOdoBR76jLcACzGtogsLO5kmbblN375vN8oZc21zQOTupWRGW2
tojVLt415NjcDVH56P7NSWcJTjvBSgGEh7hvGdchjcNklFnQopbR8lQqfcOvOnFs
B2sGTCmb+t08wLG0vhGe5LnX8lSH3FaZMX1clqCO0h/45QxuqcX2iNvEl+tO4B6O
zfPyaPBPMwsDr3ozVId8JUVeYPuHhDf9tgwQxZVaQ84NR49G1gNgpRyz2sycGHHC
pr9wyRbCPIzk//ispjWt7G7Y2GTG+Z20TZwrx/l2HojiG7oMz7Ij6k8eO3nAZcVs
VL+dBrqMJX1TSnuNXkyWwZcgARCk3kcv+8yGPdjqE2fLXYmyGnS+mlaIq/kyYyBG
ZG1hG7dzEyT1Y49jatilyN/sZgR9ke0l6tMXNoIoPz5uK+PWEg2aKEq2kZWCTxY7
F+uxsseOPdgV7dc6ui4GOzJpfI4Yghd7/sZZeQIt/StsstiEjiveKbY1MOuw5LRP
6aE5y8inMxYLonxeFbR6L+hNePx0ydbNvQvWug0VmMDVCMo5i0eZMB+WJ2xuyIuR
nwbz7LKnkgsroRjDi5NXH0XkfIoTiAyvbaioio9zP46jdBktQyIla9NlXwIXx0WX
+U4L6vVqkse+TwQMromLGsftM8B7U9GGlIVjolXgHpAG4Yl5K+KYsehkssXOWzRn
yYS7mNHzHgfSyZAupPvvtjVboau1scz6PLND5tpp7b/p8o86Uc0JbEgNZOMdE5zT
aOYQLeOkRNZfWWEW3iNECDzmJnbXEDxOv9tC+m5p2v4SAxgdXvOgtIfZU5OeN4o2
caSSdhvwOiGcaUOMc34V7/iQpGhyLmXiUCl84iIMsEUubwBmnpfOthzbPEM+ihAD
Xu8FR7yLJma5G2UY7kDTa50VwDltk6fkh9wRqRGEYJ4hQwLRyfbFUCDF8QY9nF7q
KX1fzLWt7kGGxjpK59OAQ/ZueecUAeRphr6avnx5YNJiXIaUMfvMhEbo6lcuOLlJ
Dq7qOJ7+a6YYJWpWdPY8JNB5itWbe1X+lXr2ekw8suHQsgizLLqAWEzubPoBJJwE
E7wMqgOpVzLtIg2qg8k2D55dz3uTBW+MyLJK4vnuk+l1Li2zlQJTxY6oCHlCXwR8
05LkGvDybIjmxKbr1BJbe0akTuNbzRPDQjX9WqO4iGXEKFdQCDI/0G9m2n7PfJ0s
/1qMVMl8C9MiP/54pT0KsSgW4SbIC4vdBtAj68igOfgPFK2pXBNxckYXmkKhkM+9
nQqSluNcWYhfbBmLqElGmUufgYY95m0Gib8bMd01iZfszFEv0jBpNUM9jwyYRU1Y
bcS+z7lYnV8mXrO2vA4n3EFAUdQ89jiOKVsOeHFt0tYY4F3XlcqNjW0Q922czMAX
ETNPhPZ286+aVr0lWungqUNAyibGcGWwU4HbdiwtAIJhZ7ps0TGKFdbfVNk4zGub
56IIAJKnjuDpAnUJs7DzpH0yaKa/lyVM5uDiZ2aJLrZlPd0dVJ7oLuJ4Z0jBVdOC
lRzltovbJcB/wwFSXR7Ak3i2P5HqAEZS0oK8uwxv3PBVStX1zDzF9vCg948mbzLB
QPAvpH1VZursPIwvT59skOwgFKQ1A7GdvNAwlPOiYdhci+4OG0P7pdDmSX+wAKXW
jrrv8HbE59m8eK0dtoJXVFkpYArSbCe3qKWy4P8ivnJ4lxdYBT6rQiVwJxMRoV2P
//KjqPtvcoU/foHFKGDwVzoCtWRJCMA7Lzt1tZGRxv/sLp6Yfjds+jAJv1RRZ+TI
A/LlzRP3m8styi1JU1wp+kKgxw08dO71A7hUqbdedss6JAg8gW5OdUA8iz356kqD
K+7i/GoMl7WcDDjLzFavOvuaHy7dhG02xb5dx0pJoesWWhaBFv3rmPFMv524vQ7T
NKyDGErz5KLa5bq41WZ6LhtpOjatfMuavToDp4mF8+dqIF9EOm44dpdY2pc1fE1d
IJEyIFSHmyzEij9zuaQnMLnHM46cDPPWrhQCvoXcdDTqyLVEFXDsfDNVHu4CP7tq
VoT4M2PM4Mmv66SMRGgINgTma7AbzWZ9/PIGH6Qx0iBoSPIoc8lU0UzsK/COgFfg
VgHMAday86RX55HP2u5VT2e1znkO532x20/5wAwGYZhN7p7qJMdx/BJ7CiNrJ9Xs
0v48PhL/0Ekl18tiznQghISDJGWTxofdE95Bv7fGM/15tE8g0wRcgUe8erQuJi59
zqwRmpC2JSb/7AhqRO7pB/qWcACFo5A+UrbnPATMRsMjOeAgEq4wdnUARKZlVrXp
eo+nDoQo/XL+MghYNkSGxHN8PQWzNRftL6GIEzVYcKNlDEGdZf+fsF55G+cYKDkW
i7fhou+J4RzjAznIsn7MadARR+S96pHVohhMJXPsGdghUMPTs5VJJFKeyFWfIwY+
w5tRvDmOgsmqecmBF+1xK5RTa5WisI+j8YByrtuFV0JP/GZvxYsqlKTZWN6bAn7L
639cKojOXeTSxBXjbYKo8wWGnZq0HPII3PwnOVqWN16Bz7j7LlYECHhVpp6u7EWx
mqwKPhR4JLMchutQAy933vuMncUcqMM4DEcOFcSh3M12xtpAUL3EnznET1XpJhPh
6WeY/7KcNNzdB9tMpTgOusvY9nJ/EudnOqR1k+apKLRaUFEHTabTmrTYFo7jpXRf
aS60m2TjZ8pIuZf3tpmJCLjxJ4i7vaqH3T9RYK9qI5CtoBQgv3zpT0ZvsjL1cnpL
Pu7KpUToBfcc2v9LvxQzhtU9hH5BzxYHCZWN5qzHf4Kwsi20XSAXmuVRLYp0RhUk
MPYLmgiFxFhP1uDADrH0v1iTahqEkceWqtHmW1vxbpSI9GpJlLAr/izES0JkANOH
8U9FhJLYHbZohFaHx7fUXoQLC4ua7qg8x+aWYyl0JwNvYZ7WIyzjtj4l1TaWWdad
vTMCWWjaZaxcrHR4NdejXC+xcWytD/bqOJAHaOu3J30AIEvXBvmjSndK85xAJbw6
om6tkQ4fyboE30vr/2OIWEyWeAkVW7XCEDs3gcRN5TWpJ2geAdQrVuQU3Ok+Lj7o
Ei/HBQVz8UpSWQ32yDj0x4bLBep3fmAUa+kqiHNKeVZP6i5pdnZYg46GxlqoJEfR
WfnCbwOkHzTvJVuavqkkWHTKwq6L19Q836N2rnmvhZIDXLeXO64BStxsLwlFYz9p
4v4na/ZbcSXlBGMoiKBtVHUKODkZk/DCDyN+XuY1baKFvyerrky3i6S2VVLkrm9E
DJmZvhyegx0+b6lI2Q7Rpc7tqgEOBeHRzZKZ4hlq9kUw6mnnf4AR9y/Jwnoq0OWq
guSUFsAUxj42evS7NugjmgRusjVcrUA2BRyrAbTuxj1XHcZ5YuuhaFtJZ7lzm0Tn
wAdJckfb0m8Xx1CgaUun73z6XjGjmlmA9XMsqS9mqHLOoKhBpw60Jz2qYrjXnEum
SuCN0sJoEglwMxJ6+BCFr+Zmd9mg6vxTl6tPGWkqDPjNHPnCosYhZlTrpi2I1Bo6
72QeUYtt0ocK82t06PLOVKNdCJLOzZtnZpp8M48k7lhob5/34ykOWJAM7kgompQO
NyFuafTla+sYdmxQw4CyVXqEnJBhvwITlId7Qf32mchn5Ez/hV04NSLzy5HDclz3
LQAFqN6eF4qJBCPJWMD+1Vew8dY+OciKEMfhkZR/PS7rhJq3Vdh3KkeSt2/Bv6BU
XiBfj7uhe+aKWqP903dPe5qKzS4/wqkt/OCvzAnRjos6t6m3b004JNnJEOMdX0JN
y7cHgvhOKTVmuEO8cQx+smFFe7oG4nXhN2MvCEa8QcT8xeQbItBPoOvAVOsRjtG1
fpFHIZRneMVKY6P0CFtU3IyeBH89FVh/CtsOWpa4j++UwYUtL+bm7D4kepcRZIKW
faClWgv7qa3Nb1Wyrmuak6rWlHJSayoWzWkM19CabalQ77oaLKZNSbdFJ3UUYluS
HF75MUFhsHzVp+OKM5wmvWSEL9URkipW+gWrak8feyfVipJUxlCgcf9vPz7Lcsn8
DgoIICPirRxsc6ZZYPODODomtV9PBisy8yhLs3KvmDkuSrP4oR6Y8QWiBr1IUmTf
MyeVNp05EUODLk5oGJboNa2JYDY1a4KaFNdHtVIMPpDaEu68GnvmtTGv79c9A2L/
YKi0fQ42tAn2a4swFoLntNWKDEhK5+iW/yvsBjIM76WJr+sBGk21uVGgzkP9D3aL
R9Y3uHnNVNZjEj1IexDfo9weRGYBHnFRScBl5ZE3Xrs4IvUNAjEtB0bJ8KvXfjZF
wYpFUIsU6VbBj3q5URwagZBpBLe6ISAXDuDCOnrv+awAkhhEJ3oAoVhjR3VX0Tgt
XAI7X0u4fAVKrGAh5R88ZLXaaypDy6/ZG2ifjtn5UuNHwiDSVTm+t0/fanjCVGy5
IsIjQjAHSD7CEZhsMJWJVTi+I+5/3q4kOxCYhMN79L1d9K4IMW+6KUaOR3CEzwTh
yYRtpb5MZb+9374Y0Rsng/QZFtOCgcoeePt398Edb2vyRR1oQ2H7+5GBAlQlYEMf
btEmSfE9s/pvJeUGZJdboruAfFQM5RBzEmgKWh/6kOIPx9ggFiFo6wggnQvGhlPU
8az/CpqF0LzFHc9zpCP7Jx4/IkbO5XsoZyplkdXtj/inZPLhnoJFGJ/o5M6sJhNi
pxe7P6Br960Kr/r6Ec+eAPltDy1LbFI+1aWjqGWnrUafKTjkEirCKSrb54CioSTh
JTucEm6cnQJlDq9K7iv6CE6XUvHA1QA/AXUFMltPltJJflZMMc74C7QARkxhyaqL
3kg5QhT4XbWxvY0zdNhwd4QAIbPH1WFL11F1Drkv2dBL/LMJbNamwM2JnZ6Yz7rj
cgEele+5k5EoJGAmBUAJ/r0NvEBAvmwcrLnC9Py4iMpaga6bbM5M1Yy63orWPMnh
emJcRmsxW4udhpSzPaR70FV6h9tK4N+GB2mEH4xNS1GNpXAKUgZa8Uh8VaVXxrIH
6t6A9PAchetJhI2MxuALWqJVD2gMhTRMS6dQlvjVHba7u5BT4AH+6VgulHu6i1gE
mIG6GSeI2ydDLDpo6IUUR66Uw9hDoXzn3tau97am2Q41huPcgRT7cqQlHMXk5K/4
VtlPzGGT7zqEI3bog2bcanUbLF1k0VQkJuu0XDY5fkMdKHREJlFLT8zZ7JGUIPZO
3jUS+OpXAQVS7NBaxGRwCk1VBsI58uDTriabpVfuBb53hrxVB7JgTVVrUi30vwAm
0W1GAl15rb0K8eCgdbh7OCHky3iZWBbOaaumry0GXeDHQUUUKwmhQ9ahmvJ5pppR
uHsQkv5CkCVBW1BMjfavOGqKX95YvmV5BU4en+4xKAdGTuCvqWdJACSuIQ4pI+hU
nQaPWNNVVQBGmaXQPiXvg5zS8sGtLmzul8rQ/tIByfcaVvMsnGL6OQDb6rZwJvVk
eHVXWnlyCFygDyMnJrOCd3eRS9bwiLwy6lTWXLylWe4qUc+MCGYPGKXS1Ysc0sv9
87kGlxwI8Cl7IUkwbmS7fE4ARoBo6lHKM4j61YHOMnlBjp/2bXKgP3EJmjKYYnGX
hS+50a3cwLVt+7+EBSHDtLj2GBExecvpWvAjHjepEbrkyqMEx2T/889sEgu4Hb7E
qml9X/oGaS4xU2YQcUS8zVyzh4nqqnxBlJStv3FhyZEDu3FjfeSR6GRPYrm9zALE
wJLFDIyxETc9sZObs+U7f2UzOCKJRGPOBPTSiZ1CRTsxB2pF5IDcHORIGzzw+mHD
FUQCx+dOZkcwsnnlU+Qw0xUSxA+nNbaJ/nfa0NJzSouDGrMK7+VzzWsaT+Vgwyq0
yKEIuuuPyDL4MrkVyXlL7GhYtpouFuAFjKx5EqAmYW4X7mGA1rww4rhhSe5Mao4V
8l1v3P3D3Wvb3sPH9GSJ7lFn5bP7J/Rz7JKxz24jkyLKMIUmvZk81loRfvc1Oy6t
sR3bfgY0ril7lHoUyw2KB8SGMHbKlmo4vfkpmOLSxd2aygA/FG1Dilja4eaVF+Xl
ZoeLxtal0gH/jJ+oSwfnAwWTX2Ub9dgSvuQTKxaE/s7hirBUt8pxH1JPA8fATeaH
95d0VnRDK5LIw+2/KGp3MJA0UHfuHj2aEs57DAEWTGEyikzQIx07KQ3WiT+5sTLo
TWLbkojL1eL+lmzuJWWweVQ5SqRPCuOTuk2OJBYXeeuxfHOV6FiHmTL2WW+S3Yi1
g62oLUBEhyFrKyKcA76kHp/o/hCt41J5TTu6hXvcSc/+yi0yXci9jG8WJ6MOTNSL
4RFV6mmxjJdOXd1c7lMqj7GgOFFdvPPkxLiY1IAjSa41Ys1unY2h5HaMgj+CSss1
GgrwxdzprmAJd1GRfUuvVOS66cNBpZquhp+5I6AEHD6wjDe4kXNiZoaVdtwzD87K
LK+BaVEf39mDSs66bi8jzo+nnGPk4bDVS+IgDWgFyoAj39rahYXtzr8mDrlF/nie
OsL+ummTVnevhwx9bvRE/qf44MG1/2VxeEioAQQUYlKkrV0fKhElQYlwbk5bJcgw
yf5C247oX4Y/dLi2mbVFS5uE2yNLZPyABHBD7ABtp5NWEfhgJ5AEaHC8fhkYvFt/
D1DUmvQUQtYu4hhEq+kMPf1jDSAQQ/s7TOzzX1j9tmVTUSchgbOpZxbVbA0NKQ4V
OBa9B4OckGCh39wXR2/m6kbxWvD3BKlhXoJpHXcYu0qm7peiczwULHsFNsdKua/l
nqycGe9GRmJ/wtwV1z0EzH5mCCZDomcP04/A6k7MrXnky1xk7brPhb55tMrEqLkP
kWB91aqDPxGEhx43l2EZmCsRdw8BjspVy+yj7iWcxr0QgwwZfVj51MFYt121sucu
mwgbS2FBUWUX7ODw5WO8MtEuy8V68R6T/rP3jQnscTw4JRf85wK0hHNHQUytBr87
sYM8WA6HPVKLVRamhqEZD2ov+vgtT9GjtQVjNAEpkIl8RcpGWjMUimRZikxGC1Cc
LXGEBVVB26L6RHA3BHFz0JsD0rKQ4KlqU1YVsOIllUfEDjr0buWY898rsiwfMe01
zb6u28gJgGN6pIJm5T8cHQXUB+STkSGG87Bhc9PabhM8BdxB6m6pRV9wb6bDUG0+
SyzQYRCdeTaXPij6KI6hbqMD4cxDXssXJXTDHbPI+xU0P5NY6Xjq4+m44Giy8Fdk
rd9VfWtl+3IolUp5cljOA76y7EyDL7GPP3WbWCCjqVVb6MmYcwS3drPamRyaINW/
KiIPsDa3wfwXFNuE9/nbNDQJm7N0Ya1sFxGyAAlSGvCTUc93GItHQONWWktoQFKV
5ysdCca7Y2h/mrWYZGwW0D9YtKQpTP26w8bjtjYdbIfJ6YfEzVVUIzCac9hfFoIk
NL9vFoyElZsi1m6/nGcdfBUnZzQMFiVe7DW1nzsvUHVzl4J+/TbDMOBXDG60tgig
lHppxUxO9Dk1Y0dJvha0dogvwlMxXD265AG3XQdSgINhks7dhjE0Q8ZFftxHRKVS
pYogEv+FaJOv7TWyN0pg0kqVt4MRF85BgNf8jifdNHUfiin1sqcaUQjSH4jQiOuJ
7DAlkbdkvwQ+hLlxgmyUgpscXLKjWI6zUlclT9VVKi1IyCR2rtVZan7ua2eqvqHR
GbZ0SFVBcVaPSOV5SFHyBUaTTCQm/JcnVSguWrMsdsSeTT4Oo+z5QoXXlN8Afo1Z
6xf2lp2B4LuoxBGtcV+OysVTmqGSzRPZTn1FwlwSR6eFCFh0yn0I+/ui8ueKOx20
dtEta7ytFNtfWY16R0NGpmWmweT7sG9yhWCS6US2NgU8Kvj73i0I/pZlYI/gLnHK
9WgfT2TOJk3tiOs9iO24tKJu912ljQrTKmaY4gY1gA04CgH+GkBJZbFcbNpLmJH5
SLVWsYt05IneNPkV5sbOta67/eJmPtVu+fkmDfzHVbTOmiJT2ARR1mep9Fh20JZ9
unHSI6CM2+LhlvPTk3WP5/Vh8IeDvtv2FoPgtBjqDI88C/mLkH6wF+z6+V6JLn9h
hL99cNgzZR1gPSbAoMDWM8tOl/AdHZcYUz2vO9BNvTgGwRRW/c/5MUWbjSEKtS4M
n0NNZQcDQNb4PxvjGKAURIYBu3FPmd2WYRcXWINpXeWJlAUQnsuJeND/PU3bBdqy
fevP0LZB+Umc1FOWE6ZWD2NO3FT76V9Yu1iUdCuzXgvd+ncv08G+F11MbfEu1nLO
kGGRnMyOKy57vfUKa397Hi9D2fmvNv3yZpYh3dB+bzkTiOHC6R3QWcKwNOZFjJjW
2gbNg+4nfIxtMg8UfCnyoje/Ee4BgULyOnLbZQaEVbd+kihf7+nOQkdpZrPjYjfC
OIzSdvl4r1Fi5/DEhkt9jSQUzlLmTbkJh/BqSUx+chiqLXbfyFVns+1BMoHsVbrz
WmlZK5qK1OPNtbxBmEXLoqOTJ0Xtkd9ZqzPtTE8xy0EXDyBX5leuaqe0CRVga1i5
osm76e1KCuiE57tjl5X9fGeGUu6AmUU1AzOQjUqXClr1IiTPcVoYGd7Yu/SRfTx/
G1IPXmhhKA00NxKfuZjROO8HiYUm+9sVi8+ojd7+9GuxIbI0xcZwdmb45YIIsj5y
tWT663iq5ME4jfC+TRdbOzQV1Kn8WJNPeqlS4P7G7VdamCJLgeJDqRnf58HkO6aN
TMcLhaCjnkG1KzhyP4O8cXJY+dazps+5KK7IdA2bHeBM7UurEGVgGo5+XXqIBETF
1OdgPEb9ZUk9AXgbUJfMaiv1lkdq5DnLufbaUxbnUF16puwoA/0kEvobjVKy/R49
DKbCRtR9vtkkVZi7jpZ1oAff5h7TkaleOWq98BKkNG2vBGM9UJTizOdQN9scx8Q5
Q0Ed3iVch6VQ/2ogm9qkt14lC/ry+zadvHRYgrR6fUDLSC4n01s6B1zls8QsG6cI
IIbQ/t3/BDbi1CusL7HSAfPSdWSIeX4c+l2IlZoahb4yxajgdB/SPlYZjblzYnxk
YoJ+ljMLzX5T7AqUSQP/GZmK0U3R2sTk1mSQxFHNHIMsEDPAGRY+TY/AbRRDn4ak
yEji5wBuf8FUgNgMbosKiO5xiVOWNt8DjOHQPCwL549CzuD+cBFFxCY/mrtwd9yr
lV0OSctm04scq7RAS/w51KLz324+p6UaS7CuMtxL8lOurjKp/hevGUFqmNQqnCUN
c1m4ERNgJ1Tmi4QP46YMzlEPTjUQQxsWw6H+C5eiAwE1wvxbx66/Icq+MdEvy60h
lqhLrfmCYW2+4pNKXktZBMiramYSTglly8f63ri5zvZOg0ti7yaZnR6aqDMy5A2d
tFkHt3+GHD02vz8vOL1krT7o7IR+geMPc60bRYxmJk5hbd57AiupVdswgM+/+uDP
UD96HZwhlpKEEJqAlG9xLcCBQS0bg/0tQbXQ4yeajhitJAnv+eLCQ2NQdk14V/Ig
SenbOw2Ox+2/zC4P403/bwdm1Oz/HThX8uYQGTNIe3E01aRmy7KUGb+NdQZSrhe6
5d8AVXxSwodD8cGd4NVn3E2lFcBeyF1CDvySTrfOdL8ZNxp/ASeV4TJj8NmkXjkx
uihO+1psYRtMYGK0BZAU7rdj6UYIHDKSq6II1ruQWe6D8Jo0kYzbME/r+FFCrB3a
c/qnB6rYtz2wR1Ee4GpPolWD7KSgIeKiJ3uSKo+oifSp4UtjjfMvQmahGQF7QXTU
ic8YddAE3hbIx+7hk/QNBvMK2mZ7C46con5SMQrk5446AAB8dWlwdiJEi5BXlJDg
9ClnXEEYNZs6cpIBzM5QDm/LfTAF+ylwXUin78iyJGN90Iyl2hyeDqSHcmhnE30A
64KNe8gKYOx+mwh74wMI+xvqfy0lKgDjS33mDhvqUxw1Pqe0gAIFeG4ap/ESvlUR
Rxwe1EAilIlN3Dpp2aDzTMztq7/A2QkufNABw3HMwCOEryP7TzskGLWgwqtOtaeB
vA4n4CDvmHKqQzgRGrqDcZQ+1zIsMaOGQGaqJx+pBikBsApY99/pgSMIjLn/ibGn
o0PAsPq/DI6Qf7r/3dFsbigC3dkOFkh4XCQlx8+dcnQSLxmO+cVa+TjfUU5uFZT6
P30z6HL5CH7A5uaxlWoX518Kl/wrz7Xk3i75UqalEl9lK54xtA6W7AmpKq5QZ0Qe
WCl+uhxqlG3RhC8wpmR24uCZcEN9tzIq8z7umgAIhmqWmDD5tqkuIVyunrjsXS53
sC04Txz1sKSeyeg2El1/nzZpVbaca8M0kuC+gXl0aLuxVTe6k4kW2sV3jGplHif1
Hed2fvgiQgjrObl7hZ4svRyGyyidwM/E01/51+45dtI58115hOS+mvrP8p16PxeZ
X4BixCUrM7JJyHr9+0dBTpnTKb3bdTWVUIBTeSanWFokf9LJ+euy6jK30/zDXUBt
q3tEEq3jCEZic9xx9LthIXDzJjsEUj8d/6ZrFOwcD+ANU4lYQx+oUa44VeTzteu0
GX3V+tMV63k8BZAbHMhCqoOZ3y3zK8c1EOoCvy6dcGs6gwaWJqyRFGe9Yl/hd22Q
DlV+C9HfTVZeNRqvp4JH2I16nt6TD7t0Dk7nD3yzYs+lOiACfDM0C+OufiIRJRsd
L00hsJrg8y8ng77ZjjvzUlvRdHwY6qyCzVdbtngEV0WYqMP0zy3IKWevuWIyZMDH
jWZG20gyoNdZFyi111/Z7hZr+ejGXWOmzlZN7yfE36IuoiQhFTs0+4DmGyEIU6C9
CcyDRdfXYrHaK0SJGOrtlwJJBUfLArVqivH+AhvuSPG/K+J4t1iSuvFg+4UP36zx
liGg5Jt623JnIWoXlcyQHRXYc2sHQ1MaKcJBauwjjBZVmmva9DIWodsRMR1J35vn
qyUZd8Exkrb0xCjqXx54PXdL3iV5M1LSZvczGIeXPBsA4VlKfFtubF1t+em3Ytnu
XPFekrvfxy+atE+dUVOWHoe7ARdBLeqrz/LkVE9ddXcCyqtg8r0XaJgqgVYcpBe/
KjMyIMjqbi92hB7EtoPSMce+PDjlY7sjUB8qtLp63Z/SZUZhwSfe+zrqTTWBLwyO
qZf0yK8Hem1a9IwbntaQ0DJajOOKL6vpWRmu9Cls5GJZskVEIFN+d1+OSz6Kn+cY
MHHLckWgNAXuYb3S/48csCpEt4XEgiRrDM51/zXosMl0jnZFaGt8sB71PKqGnc+a
KjwxA4iQruoVO3z1bqfcfU1xT87GkyVS6gpq46YaAxAcInANKzOh1BfPETJyZwCP
UI80HQYTwbMhuqJ67i0CpreTVU4Jb1Btre04Q25wy9nJ0jNx5ai2izi9QQghXO3c
AV3c1sshyqdix3uSVdIfbBGuFWBHzTmKJRa0uHlF8QBupk2rFcSdudIYax82uTda
6BntMrqCPB+ZjtdmbQKzh7AhTpiAqcd0BDH60XFdF7O8Aupc7VnbWo+ES9WPNkLQ
7HzYHmrx9BVaf7NLdbSnYFMPwV1WNY+KbG3Z9SX9jEIO6KshlaQ7CIPy0bDEeRnn
pCx+99JCGe/yktulQ7GPP1El7SPpMcvtFXTfUZIFKcXaW8q7VQU7m+d8rFjco4y6
x0JRWudARxEDHa/2Jnz8Ajr86yuCR71TjNOOMiVNI9psDf3XCfViRBUQKf2AVwjN
wxgC9qEPHPIiLw6VvRjNHYR/1g1ptfkcqnLGBqGrMqmtAXJpj5smN+8a16pB/LVL
LBKDivVA91FgFL6n2O3/DYZ8EKlrEt3UPX1vDlrWfem+cL/mn4kO/I1P5bBqMwxy
Vj+ZnPVh1q3g8/2+xPcCXk1Qyfhj+kDyck4ENTYrgJgFMLdpRB9xAK+YubGFe4IS
/EH4izrnBfJPS9kcX1OX0Ujw3NapVCQEKXHr78HLtD7InaVULjvQwHnIgx68lFWY
kQi8GqnJaTUmhPd1HKlgu0qifBfLCDGqEX+EDjOgUV/PDuhVNzaasRP2thTXgi3n
nODT85krIWmytDK6WYB5vlTugX+mZJ6ByTeBav3Uf1BubFcLPl7fN3FDn5ajjFS2
OKFTsSJpUQXtc503g1gwKNQu7cH7q4FqF6y34NCFZoqkkvX10mVwF0Y+yJb0OKgp
EwfXw0N18m4+fMsmzbokqNF/mi7k19RTiFaswOnCzCaV3G+SSb29nKHx5+7wg7VP
jfxNdgL8mcji3YD/bScZdXqgTI5TRVS6ThF/Twi0Lul4d4xN8WnCSr9hUZH91YG+
kjB5YeqnE4r1/dSspXVyFtUOliUBFMI6cXDKk2NQYXO0PvtooHB4s2B5w1g+2S0Q
TmVa1WAGbnJOMRD4qsdR15xvBrrKYHJs9/o3OGWOg6m2gGP3tAzB/eWyJ8Q13lK2
bGgcP5cHwvg2F8gqv6s84Q5HI3rJuPensv2gHsvs3PzYoALA+WjVvPJVQ027Zv7b
v5BK4HySiz+/4YnUxbiLyuqNTdooA5bvYO6rBLwwjlvfwVowaIdRbUnt2k+exK0g
EWbbNoZtD1cbYFnLlZtTrTIZIn4rYmG+miCHYGhNClp90HZJfThH8ofjM1r2EqN7
yD6iCtZQJjLeOuittMT41CubU+zKK6AfMkJfUSGOiJci8GrDBeqRecZXaMo1qDUr
QztAmpxu2mrYCcDjpBJXsFA4lQzwuOcg5Cx1+rRMgz5AwieN8IXGd9GrGE48daCr
22dmjn0cdFkxUPPN8hSQL9bWBLp0NhaNRgRnMVhQN7lSE1fm9ZHTB4ec6XYsn6Ep
oJ3sb4EQZRfXPLFz59bAfno4QwPL7eOrqrle8r3TqoR09ZCzcBVvyDivBD+a8XBL
y3ifs7aykvpfPVfJV3WEvIfM3RVI6uZzVaHxjDk0xP2h+gD13r/QyIwOACsQBa52
4j1MZeOojZZV7vAFvTsXz/9INVfHsM7tPY+ZTLg+UmulHse5mFInI53ma/9QXwlc
0HXa+QrBmi6bcv8DPt1laMR3GbP228XQaAV5P1cHi5vIjzJKf4wuwbxc95WZ4iP5
MdBYX6MHMDkczI+Kmmk5Nf+MKrI4Lyqi1KurXAFbbT2/UIQxHxwP7nB01Wn1nCvl
3EwIZVTvYrZ7IKG2v/4O91XAncLYH+naCjzURyCuVDdpb9B+TJgTQCeTW8qXf1/D
NLKU+cQc32Z0pthZlC416WjdMFc+cZX1Ip3A2kYAZUEqKk0kGn9WcJBBxXUr2uUo
64Iru3u9Gk3syLOhZ1Fqa0EPbM1jj+V33cLbiGHul9KkliBUva3kBbGPt1kC8OKu
efFpzXWg114VTVD7BwBbRAhYZdFbDtkf5LzF4ekuWHxcWUPmOqSoAnfLdwQ2Lehb
zMykRRURcI6NsgWtdd0d8e1755uexORi54LCwiWpmTdNCv2txl9krvLjjbc1Gcox
gAd6BYEcMtubWTDumuxDQ6oX4kK2TfPbNR50gA5gh1lV7TDnwDSF+myKv8b+AYUu
WEv86X3fYDbYo1tWLzVZO5hM0faPwNnD3y7+fSpWFyaouqMNdFcrAGQhO/RWqFcB
3ukD7YDmwPV6X21IbSgJ7nX0aREu0zE8kWT27fTQUn8yv9WUFE6xI1us3IB36dds
oEUkpXGQUOfL7vMqoh+lQEDh6auB/RnHMokzHc91W7ZNgwsWN7DzsCcTgp97Ef+R
HSAT+Avi7CnCSynLyOqe3fG0RP0QpNPvrc2NiIcdMnG1HwBklWBCGHEo0oP/RUln
uTiJLAbXkBBjcXZlOfjsS47Mwdy0W+JbtKvDXqV48SYAbbjtuxn2cXj4vemPYzAF
5mYYEWbSNoOw5M9tPUyyyHFOAGzMeamMRdoao1PTnvOifk3QSe7gvP5JtqhCnymn
GZwT3jSKB5cZrtO/X9qPMzQqb+eee4gAXDFeUU361whCBuPkT3VFbD/9+wavi1yi
AhxR9uoUwTsUDp/zqaBH5chpGJDbcEz7Ryqz+tauy+4DapeybR/l8v5wL+J2jPvJ
QFiOQQOyc1JM8IH1bm0+cP/y3GFEVyPIswxBVr60fjbxtTGrt1ZgDJG83UdNblgg
T11FDEn6f2VU23iGHz053t+oFcG6V411ki0TBK4TvHh+rZocgIGFs7Trft5rJW77
aQLzzF87FCRJgbFNri0WmBXUsBMOO6Jz4maJk4hFa/RdGcytb7CS1X4A0fi5JcXs
0xvvEdNbf/nrDhXQjsjeV+00d/e0y6lhGaPShuZNCd0vxJ6wC9PVdsDyisu+KYCa
I2b6XPzfZyTNoaYWBN7gLEVRF1AjnmErHO8WQ7nBCvtflUMASLbeb48PrzyL7FRq
ryxds3wrloCzCUoeLkCOrqV9eaLdXndDNDI60msUNbo75e/nJ+TnTf5G/r3wSA6+
Zfdejup8yxWYDWAjgvzq9ymWrdWesppqRYWHr6yipeU5URqIF5RYtBOmMPkFEVVG
HriFNfUf+hr3y12jcc7YspAduRAcx5aMPOx/U7l0rFmFDE5cs67/XF+kfSS7OWFw
RBkbmGcnQn/GEuyOLVvOUhiM5fMtInGlD2Lt9nuRYMaTsu7MTKfe3L9F6RNNTuti
Px7g2QF1Ux10EVoKam5cEY0Uq41PJIKLz2Z+Wy5x4yXBoq3BnFSYv835E6UEyCXq
5EbVWOXCUN1ALIy8tJxOlOAojA6IN3Um4U86rJjM6AbNxDnDjP4aRqdkMgIpwep7
WXfugyumBWWmWHfHoD7Wj1MlUojKnsg8kap64H0hZ1xU8Lm5e/cgok4EFSdwaMit
ZZBNoTlhE42lB6ZYgiLQ+Ut6EHV0kIYH40FjyxqWMfiVK6BRYLyoHDC5L6vITTSY
2omHigX8yR9ttTeeWc3qox4zGvjfS0JsEGFcS8ShRQcjHtdybBNS7TWVMHZ/TqdH
j78n7G6W2YDjqCWiUTzDdkL3GGGnoytfeNHjKZH+zsoU+NKn8s4RFxSRa6zzRE3l
7DhJJXYX4BIQCH13Khau4gTB1obo9vTlpjUR9ezmLF+OUuZJlJ5DYdyBKUQPo6EM
75teWxZzutiLDVGegTrPUMU0iDRw47KQPEEPrT32dlc7x7VedyxNMrJt67g3b0iH
0S2heeSKJkDWsEZiwU38PvbI6rEuIHNeB6I6ZCQ8DCxyRJ+acBH+T1H79C+/EMyy
6o4BdpUOPesxlIYIHS+UXjCDn5JpwVCm4Z0qYmlx7st76T00mirh/MLPJMXajuPi
MR3PAKyz/y1HDDWgyuSMUJXKE75DYTeploJdm75RTj46YE1k4h4Z8YQCwm/GSWGk
hNVKFi8uPUPfEEBjuyX1hTYgwgveVm7J/eYjhhWf9PSfV6Y5dit/ip8BVmxH9yDf
CGlqcCUre/BLnUH1BjZDfaJeCAu2msN6Y9KedL8FvfGQFxoFH+F+OlnfXosBgrjv
SXcBw48kKfCpNpBST0AIHKLPh7eKJZRVo2x47u98HtDjGnjZnabtVgxWza8ek6KI
v+g+0/VrL4S9UgmgvXpWQRUAM2v91psUeiPA37T6sxYRpIfQG4m2OP0PU97Nk4NS
7BJmhfj3kBkyH/kDAw/L73kNEUEucZLMmYxxPCGRjtyoAlf+1OncvjXzM+IMinWa
A12mu/CZEG0XllOZFOQtm0o4XF/YM5UaEIrRD/nRXwWp/XCUmtrj5HkCk5FQG2cM
2SrKXRH9UoQL7HyTLfJFr/1CaqvmJhhbUcoJX9/mmP27tTH51u/4/bOcmhlN8g1j
E6/3hy56iz5Vn2NquWsESHVUMUxcXzusJSBOKAfykxULBE+/EjVkMsyZm+yRlC84
XwubfrllcTcrW9DYDOmu+qDxcIGYSXt+wkPNnU52L9qnxVAA91iNmpJoR9V023Xj
t74YIohY4qB1zPZxBeIXGrF74IFHh6kMWP086A1z0N6D9elPC6KatwG2mT/Td0Oc
JdWKs4NkBr8D+2cQGb6ti1tjDWDyJR0huJ5vz1xeqaX7QrFYb8roi8EivaWbu6Pf
oojBZEvI4f8f7aRknq6SdQsGVvdfoi9WltpQjfV9HBcoaZXTxq6dLRUfPw3OPoNo
Qc1XoaVEh+7/tnFGuhMlKmU6G+Fc3/fYmAnxVMCOd5wdkabo3r0dOR8i1KJRo13+
VTaq+jcNnG95gcRxuoOpO9XlmG+XCGjhlaUoYts0UAN837w/O3IHLpIcALWtc6Do
lm1mpPUkHSHUdXdK3vhWNHgKfV2b63ktUFYOMLvGoUdpEZvedaSEwitbZHrXsnaW
FMhBVsoMoQSBB5N3cuirlnUqOCJtdV/fET3XWeNMOYah4ha3PMvE7K8/ykC91LdF
22gz0xdXhWpdrfwQipiyuFUv2upmA6qCX+QaNpJbAjmtFkN24tTSVo9uQdkGXxXM
UpL/mksrzORrPv6DB+98Y3s7grsFiVZeAQQj9OMEqrye+9422xGn9BbbBTE6wryA
znwUy4RHrv/yhqNx4hy3eHuwVOmDpq7H5Sl4BzhOsS0BxYgOfDg5cfWrhN7IAdOZ
w65w/5GDa9Iryx3yCtKm7t8j7Cxisbv1gNuCIC6gLXYl/X5aWqi5KMjibd4T6R3Q
FEY5UusevM2jm55omRNdzObkItaimue2uM2YKzl52b57XtDHu46IoWRe/6pAOZw2
PvoRUeuHkwxW02zZ7At4DfYfynzOCCwmLN6Uslas1ytlv6U1nVGUtvX9vGugqz8b
6RbwklYMc2kC6TAzQAsBm4CiZ4l/PcUhN4OFXdfXJJMVmqewCPwMMuzm+/ZfRNvG
hBQDEn35+XSWRFIfIAzy+KHKBMEsFApNVx8tlBlK9h4cG7RUgjBQH6yQMhqQiKIA
QZCRT4ojCFkXeN5LMs3jy9XD96EUdlF1XBIcpagZNELBfmh/fntuhPDf1x8b2vLJ
Tps7p8HlF8Cdd0v85mgHcL4A+KYMF0jHogok4imDQg3OBxedFaWG0MWA8QC0hrhr
aX3DerzzkAiIjyiXzBAXWjOumEo1rrriM0IDg61Se/w8oWR4hX2Wk75ofK06gvOS
Wy1yWggtKMEHpnkbjf9KwqKsMboZOfVhN0I+JN9+Z0BrPH654a/hYAwQmcfPgAO0
FoV6QaB8cPan4LWK6BIwHchutgwlwM438tAnSfNKHtqvuxhdhm8+Opu6DtvX9/dJ
+SDRoagcPNHrg+ZmThgeLksq3ZleFfY1mak7CkkKzDHh0XVbcHqK/c6UuFneJbN8
5KYLYe/mKQoX0XYclUS3/fJ08uZXYIzeCbcA25XduxfCDgTPz3qYVXW5ZWJZbWEb
loYE6Oj8wX3sT76XJsVs0qP3fuhUCZE5RIyxHQrVARaRaR0sg1gtBPp3aG4tkESc
tOVBjFk1KGcHljdYCGnt/Wg/jDndgr2WfT3Kc+e9oN4sCAJ+IYtiPv19p+Brx6IH
2skIW8TN3m9NbtAlwhAhShNcANWGawDmJ6FyrLVb3qXWMYmde7jiudSyTkgfOLf7
N0RIoT/2Vn+bR4hA6nxTIlI8Q4c2v6gSkwDR9mBOWGcjrZAXFUyckUZ9y1CEtku9
sYmB4wyW6fL0svUyMMgvOzMGZwvyoPMPntUBkTrlYxyK0kmSEke1+qksvnXECL6c
V4JMWjhY4dgGBrZ7cqOtenIIO2Kv/4nEIPLQfQJSkm00f9Sz/Jnf5urB15HO7IyI
hwH2a0XtVnQm/fxrFO/XuDlyobQKCFeogZ19wPaXh88mqpFTYXzfkcoJefhC5LKD
k0hKcl7cMpThvJbYPyOm75zb9BR0mJsQm0HP2873wJxwqXIRU/H397v94z60lSHG
AMAI3a6OhHylXjsFTJHXE0y5bJd2U0+G2ZmGWZWm+3gRGXrwlMJxx8BI9H8kDGwf
kfrolUbbRyXtKlUbUngI7G7dyKO5q3QTJCIkH2lcJimPCGk5J7BKfDC4Wombqccl
XYJTfTuD4TCuAb10EwYPUy6C2eOVuTRd8Yzi3XVz+JAiwDpHv/F+OXAb5taNT+7Z
4xPq6nClk4We5SZKRHwN72hu6YgI0JHoReBMGFzb9VjjxBLmBfAfOV9T19MMSpPN
KDfOh6OmGFzdsqsHY8btfTaV7aozhcIgvtHx+8P7QSks9NmDLFyetN636c0cCiwk
0pdrYT+KIyYTdpbl0aka+tBJGuYJd6+6RS0S6WcvSO4AwuC5mcOvOrbnxx+66xOe
86qrY1CZaXasVcD7zQnhSt81V+/ZwuKYr6S/Cy0HOVjYZSDxRxcs0ui3+59E5ALv
b6sD1PFJ81ktCs8zMDMou2/JPUgAJUJutJ8SuWi3Wa4zqhE1BySg0166zv10Jk+k
qhhA3YEgYMFZj37rJXtlNuSqjF6onk2DeL9aec74qgeIvECBsJokMfQUTbFPwEyj
Do/ZYEtaQqu+/V2F2evbYz96a+2rZxQkEhuHtv2dkwg9AAt5WKv5z6/KljdIptiX
jAsCaRkwg3tARuoKmS3MUrpuGF8xQcPyAAjbBU5eO/+yg1OwzvyXYYTzcghullkp
xGocG4vzVlwDrlhjNVU3/P2QTB0odPI1e8NFkdTKYNgfwXtxbFZKLfsMmiTc7M/u
2236QtKt6WLl1UtNw/IncgUWVjbzW1QE+vxCFtthlVgJNf8Nzwh/Wg2NkgcysxPA
hJujyEWcW8Z8UDFgVlQpBrEXgtq63iZq1M+OBuX1UzXLymHnSQr+C+7pVFD3cLWz
T+7/Rx1yy4OZ0rHLCozBlFX4cjt0xDU+9dfeEqV96wa6EUtAEhgmhooDxVJxZdBm
ECKUwEi0OD3BCP3qe3nMXrhlBrw83HKnJPUaQky+TXUX7C+d2Rs4h2UK0M5sdhpY
YFltGDkp63LBPSEJ3l1oeOYqsY4psX+QgGtGbmqpVHHYyqMRjIaiEihSUbbKDa/y
ZaZrnPbMrrGjhHmpuojrXw0/xmc7T8H7sSy1n30lJEpxk99fexc8mWXPk62We1qe
ze1ejZJUJ2kuYwY6emHQuAYKOZmYmnqKUd0hg9un3qKwckJkzP64nmqyfx6pnx9N
WR6bcDeQCYbZIYqI57cXTFeT2buTuMn4OXd6F6t3mFxFUyzjX/AIGO3vk4KcZgEv
odcK357h3WonTi24866h2Lp+mo+qRQd1j/hxZ+g3vT9flGq9Q0qcS2SQiqhTlXPL
NlbYjmyiy9UBdMXBkIWp0DYf7Y62yNQPrQQo2iSh3idjYHsBbeIShQq6KY5mgswH
pyyhTqnKC5AnVdAn1/jnrt7VxttBnmH2LK/1Sn4RxDbAj9LvCgeqnuzLSm6F933V
QQd3x94q4qJR14K4ekJGRIFFWKEAuCXHfMo9EE4spJyadvbTbqeIdRFNr3ImL+oV
YN8ERr3fKnJmGx43juxOyx8fci/LzQNrgb+cMaTQ/+TuRL+ayxPaQWGkiQzh3BcD
VF2cOFXSudrGFv01ArY8Cg/wwCrAx+gO/LCWXnF+DhqIwAGMxwVysnXGtoAASkaT
1Gt43ChMTVErE+eEcbgzQmMs3m3fBSOy9Qqu+Ptj5O8mRVN+UiJ+JBCCXa08Sd35
Wbz/oMK8iTbBaLv8DjDyhhiWHglyVI1xtNiZMX7JJ47MI/aPz2gVz7ji/taR3x6a
lSI3w2xv+uJGnpqRvIVq/oOIcfMmKueAEnT4c0VKnaFSYU1KeQ9ptH27sEubLZWU
BC7jldc1XMYVhDpoe4gcT+r6RR/8nnujh20wJ1WSWgbKSlNwRAA9vyPl81nRJaK8
R0CqyZaeSJVQljaheRJT1uFK/ugZr4fVUVgI45Q9Yk0EPAxJS8uIU2tyMpGtiK4+
vpJ5Ou8Dpptfe+Km/N0CsR2nuTx5/GWmUqekCCNHRl/3jvcz3CXw1gCfvMUxlFn7
J4IdObaFS11A0G0cdMuFJQ+QJDBxvTMTY9vSX5qI/BsMkX8H9CRQZx3cpQml1OW8
Agfbeq1JB3mjM65ZZL1PW5mATOC2JFHGvKB7lFwO+rUWmHWwA2I6PLV1qSDWBYi5
jIDGFZTre34ZCDjAfe4DdS2WAOrWzWUNhXphg9uAjL4hgFBDgJAvcs7EMY749hbf
KFfodS12aQocES5B7E/QTKn0Ph9HlUFKyPNUVTyIoQnUIJxTxnw/yzkg6dxcvHFy
dVhktWB1OhltFSi2UhPbhyosaxn8rxnMdjfnBgT8j3B5xHrpvv4XCW40U3MDDU2M
MGPE/BYFrEy8nwPP2ezh5gDcf3OGIUfUEbnJhdyTuj+CTiW/a5L61HKDSpwHcAn4
Tccb88Z/jm4AlbegK1C7sYnYZfMr8zczCavuQ4NuEkcD9LyE4cr8EYPLn5f5JMv4
LUmCYI6/kVo1DRRd1jqeVWyfCWbsW6nT0okfb2XKrNsPFe7RYKu3La4+0meLhJQ+
OHC4AJOYWdOluWRwaB4hlYN+tR6CcuwblnHZSztI5XBNwdbnPMN9US8JSZj4l7mv
touZFqG4pDr9XWbcFTSoqDFQP6ncKAUsnN8Q8PUwGYPq3Fd5FGla4ts4ko2rS8st
McBrqtwNHaBABNwbD3IsAOsstSp39dOjsXgCP39n8acOQzQccSVOPXog1Oz4704c
y+4A7y2CgQrvpGwU4QDgWFS1ZmLlQYFbn81K/Iz0UWpRmrhFDiJLwOKpI8r23rqA
mEYn4g1CDNbqullpqrjmf3twryrZCUWugTuXAj64670yrPM270xCEcGAnPBDTjlt
EKt7Iqtdup2Q9XyxcGfHKARuUylwWEaN5dlHYZZ/NlmNGCFq/JWkjLYdXnPTi7tM
glmXq1PfHlX4fjKavpC6sTi6RDvyGHIeK+9plvb5y/KBnrJmeDqdq7ignVxiepyS
UFFv/JPV8wdhFZgiRYC+zPPW8cw3vSribil42eSUniFfPDz9nZGnVKl1n1PTWwdl
JBUGVeFsGqX2HV9JPlbG2JZLkS7mJwKGI0vZgMdC54YXPKdNV684nM45u1OjvZWv
NH7m62706zPdsqXvTIZH3O8rlaQRAMjKhE+ZhkMWecYjMsvtC7fJ4sllc/BGT506
LJAJPdV/EJi4N1PAgYF+RhVVtx0H5qgOZegP3w5EQNwtOpAZ0z6Fu1AIpbleg0xk
AkWpjfIAXErBR19yecQ0urDhBeQTa+PSvpocLGvx1h5prxbpXh5PJDXHaFmhRpZe
VMtvPtkO2J9mSJER+XdWaNFdN7yqVIVRcKVgZa/bd1/ej/8dKurWEYezJmbO/arQ
R2+2zLrOVU6mFQ67rJfzOAXR4tTuWs0FQhNM6m6bhFpllW2d5FJ/h+ibx8JfBGbv
YdSt/BYTGIQMZ5ZN02vWkEmG4qEF+Y01S2St7d0oCtY7ntPs7K0VFtlFASKaovUh
MbP1hNxZMG2kTl1+6UMwI34nIKyuLbPzKWo6iZqELoMdqMN6TTjUOQgytLxeeyIk
YZ1WAViUw8FKguJx005yicmkgccIQTVYWhuAS0yAReiApple4EDONvM436baeyr2
gIz+uCpTZRjpaqo0FYJ9yVDqJXkYF1rz7w0GJ0VBJ93XmxRloMsT1Q66gJ87ZT3r
OBVMN8EO8E06NAz8tAwECvegkyEVlT7uMucLv4UmxDIKfC176lHUeR6YEHe5CLLe
QwcgQFN39yLM0JjpTgnTwPJxDuKD0xONMDdI8wsRfbu9ONJOUG9gZFy7418fccYk
wyLNLftW9+cg36042ClVivZ11EFNnSDY03gT0D/ie7pAqfqckX17t+UUxXiJTzvh
stWC5edLi+Bptpq8pvbXzFh9XrpjeKxhqt8iUmsaGTTysrRwRtv5H3B0ZCVs/rJp
eGmdKIhP2kkCkRPdNO7D8JC7Tayslu0RhkLH84Ei4gHlqmUsYV7DnJLDGnmirMzC
enbSMTGgu1ECK3ZDMgn+iF72vYykqnzkqei/oSfLSxMkr5B+BTFeHgdtS2sxRu0g
In4lklJXWwJ3Z4DMLIB4GMo8SziRt5wDMzZiQnc13HQ30i4/Yt23JyjFBXBnEoPy
0buzBCEiJBgvwqQ2SjrcCvbKo9ar5kcwaDsCFQhRx8zzYcmSeKQYPB54B4RoY6hy
O/b5IzPSAaDIOEUDIqYD8dPH5Ma/EX17Fj3NMGM0ftSP9pLIPKYxV4a51iRh31jx
dwsnabUjNTsqw1SQhr/TDgFSEZpqRuT1U6ADLEMd5WgXVMzgJzd60Vu/6W4N9SRE
EOVz4QftZcMft/53bpBE0GbafB2SjYm4cm/35dOXUBgfbpu0bfi0KArOzxTEv1Tv
UTVcFCe50pS6B/QjW9haVBLLm2FaVac4w6A2XfXCioiF4jjGrQLPy9cS57/EgC7G
EbAVlqsJlB9MgdE45IHyMiwUxFJLclq6+6XwhpzRpwXtPpGKnG4LrgJfqLAkghHR
AUmVCcrdO83IoiIMyUrBeihOvDTl1o7cCjxJUVFLGBOLeSJOKHYb7COBYYa8M3VO
8eKy8EWz6ZUYeaXPRSmlMlNinR7fkhj1mdzByeBrTvgRgFqprFzXmvIwPFu0EPNj
o519ipRU2tcirgZpKstVvr7sTcpZeNPQDMEg0OYgoI2UVeCD30hRx0uXzZz2itQi
deDJHOA7Cf2Equw4mYuIZE/m4pOO4uXBIRE1FlCslPAxbnYODXxjhkkR/XQ2ep8a
jvMZMaAalAzFQWeWb+rZV1iGYvajMYwpRp+/mq+o+rRbhh83IyK2va+1cjqDRJqt
O0e5f0+N8ioHYcxJDp2P6EdOMq8N2GLuNUJaVhxqJslV+F6+blB8u5UwkOYCyiHa
4L3oNkTxJfKUW0qeUNdMrCicGV98PCLDyNpmprEGuX1VnoWtQDdwESSeTznASix3
JeaW7MXC/OOybUDCijbnzQvqHdyJQJe/K2izmsd+jLlnsHPjeuJFjK6hhFi5pmD/
8lpqxO4hvL3pIDmRj0ffWrOLYCSlFnE15aRS9+ct201DBDzn6QDX2ai4wk2dvR2S
paGqJb8ksYioHBR3cCONavdFs0b61GP+WSaWK5+COr+IWG4iw3vA+xYH+ZitBhDg
rhgJANdkQrBpYjYs5cNF+Igth+RTqOFnmHWmQR39Guou2GrY4sTMWhygCGw4hSL9
m1da5QwOzb2l5beGBs7O6UUzfMis5J/M39oClbo5JWwrBoy7lsqZJBGEXCcEbvJ2
V14Fmxhmfx1TgMRwHrlZOV176ZUI9sc+dwPU8lI73UkW18fPAlVYgHfMeTtxjDGP
Gu9S+noxznP4SPw0ADF2JfcE19sl5mNNfeCXYg9o23WeP1Bi54xmcGc0c/5KcYja
+gSP6prRm6MJ+iIlWpsFswH2eck15/rIsPZTGjjgk923hd0AmdZHSJ99S5MLAB1W
OkFj8yX5xBBbkciBWBpMLLWMgT9yBSyRB1VZ3hstBe50G+BJgWh/UpcBVQYbicMa
P8L5cCLaF6EJpbWDNWa+3pQwAeObkrW+uKZIHjpTm/CXfk55sT02rPpblUroe2Lp
bbmJWAxEGY9MuF7phi1x5592P1Jn7z11iR/DKtb8V7P53mZLFP3sdvAgH/d4w4a4
sJK2jjuV6Lot8e/Mf4dsYCoU9lm+OiSg4X/QCKYT1cwtdg2Ge4Inq+T0CWb67Y4K
ZlWNtDJdD5leFJ2VMj+nmXvOeOow8SPyNOUkqsOK9Tull5lJqI6BDFd5dGjD6knA
lFtsZXiei043Vw/5EptHfb0AJT1kn3QsKJAE4dRaJB//ySlj/ow5b+VjIo2svoKf
HUmzzuNpIFFy6RL2HHp0QGWOOipY7WFe6PIaLnqCNRB5lEmVbzvBiZv6lMRflL5A
EerD8rBpkUG7uZ/kHQyc8b1y0PCYzDYVNlu55Yd4r5J4e1ASJxmqPwBZtug7KQLB
uRLcOXiP6rjpeOF0xqcq4Y91/5/I2ZXKwHHznW0aYo8KhuNYQ02kL1o6Vn8WKQ52
sjOZ7QlrCs84OGwmX9R0sAmYolRw/TLecFr0omWMdSzZEsxu0qLHz5nTxFx/leTt
S76qXH6wFUytMsXjAxrfWnOmHiICthFtI7USpiMfNGnaL+R+nrwkoi+VPd+4+6/k
K8OiEaQe6C2H5rRu9row0bdIz24Lx3T2FqHYbiPiPItKDing8Y766QF9QyIpTMU7
LlFSBK2N/NZmu2rKtTWroyXB75aelpKATJs6NonoZOmmkV1EetEULqcCSJWASJFe
ouKOptWM0EclkNbnTxEad9EvIu7Qu3zG3g3w0OMj/B5rbSub+cZPktvFnRIlCCFQ
MVpgGQ8RUfG4TXpVV6J1BpXObo2mlPkUyDmXsEuR01LyZ9usZ1PUMxpN5PzDIfoa
Fa0s6V3UwfKYs+/fb8crhHqiLyHzqaX8WTRBgNPjOltBmPfOrtTtlCTa/IP0PaFy
ehsTmE4H7kk4CANVnvw70QgIHuuLr8AKYGJDaTIboMCZ4x3mfSPyJ8FLkaLPM3SM
QjtYU1aw9fzEi4eIazjOzHXAXF3B0Tkka96eTT5Im/3EbRc2wIStjldPG1kBedGN
1z6JNCbtUtixUrJmDmpkev2adIX2n/MbhlrrNAV+9HeddyZP6Mvep8uZlKq2PXaD
wdBAijxbBMupOIAtvmasoDiZe48Hsn4jjj+p5zEzzvm3y56FkO5rFunq2KCT11pz
n8B0BSJJwG7amd5QC7drNBLIX3eM790V8W+F3VNgqAz7TR2MCPOzMOh835Ke2LhG
onkmXNZe0UnbZT1+IKoazV1/UY5Vzx+9IEl6D/tBUuxSApZ/DOmwF2pwhWER1krl
L9qrJzxTnt5QLNQncgdjBFOzkgkAKb7I19LaVaB76Bp/eXEN448iyopaDQYLnuyC
D7omGLY/ElH40KsbEpASWiCcsJkwwZnYW9RJwSRRULOUHSz2GZno1zZgLNZjjy7h
aU/DoQbpOYRhr8XivBm7fQ==
`protect END_PROTECTED
