`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRbhw3eLOYDJ24RYEfOzyTjJr7ikQ5wWss1KevKLvkorP4DG1z7s4n93qsFTUho1
E60gZ7ZNMhW4GhZDGXMS/hjZ+nC5aSEEfzGdG3XALl72nnZf5pHQA5vZyK1slZPD
zXVuOy7PyxfI8oHu7gNqRB4tXvT4m3x6qlO6YYL20apxHM6Fl98tUrhTKli4C1oK
R1iyuukeP1q+qLo0P/DLWIPJpk8BR8om3LfDh9ffZlGlBr8lndf0z6AImR7KejbC
eA5A161YuEw+pgEmMQpdLv7JTAFplaQtyyUX6b/7C/SNMfHApDMu3PdKXNDblMc3
7+0kr2BWQtHiZfLFkxNnZW2P3WE/ZwqMhgg6sJJpATJFuoXy49ltfaIi1SfRxNdX
xPLrCfBteCcx9a6fYA2yL6OpL5FtEnFMNFYkM68y9fCpOpb+7T9Nnv8G9W78SHYh
rWg+4M8fPMpvtOJzafTqDi7J+8w2ssnYSVBUONUhql63xsMqZvd34ieTf5JW3Q1Z
FuS5AUR4oP7Ebu6kwqPPiLNhP+cr5bPl2+6/MLoZGDyGw9ar7Op5BM/qOi3U7ZEr
QNnGWm4IQQdUASmaVqAvt3wzCXaiZA73nMgHyuOUAR8=
`protect END_PROTECTED
