`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SpxG0ElojPi3Gc6InEbXfIOpnSQuJJNHqphzjWhQQAcXEpw6+dssx5COWSXHDdaN
0oCM6XiALzHunyxVEce8x7c3FMAVJK03B4H2sGito8eERTKAjUBoP/HNnA/FELlB
PsBy40frKaSQiODgdDCcnECcSioVVajQ/Rd53M+sf/rmq4IOu5n9aORod1ic+Odq
64Tm7IrVhUuQSS53rZo3sXaglHhL0QvqXR/011H1HWYLdejacxBQNQ5Dqkklx8IK
ZyNE4dH5gL+yArPQratPaq4zRhRvRvWioUb/d0n6dLFSPb9/6lymJiXDhPShBDba
usW8GWwGwkhZUrK+ZYvo+weyiHwjaReGHOm6gA89kuc=
`protect END_PROTECTED
