`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XKYKYAqVvRLO3V45uaveYAa8K7EktxTU3XS98SMadY30ILM3+GXU13w5bwOneUAM
LrhVqybgbNYN5j80hxwaCAx4MPyeFu4ZDDuf1O6KoJHLvZNFypecE+C3ATC76REE
WwFMLwFuA44RFoJrEed6myeWjpEB8nXwT1JRAaG/NWeIrVLoDHXywtGI3/S+zDEs
M7T90nT28LlumK7gLbLoX2MtI5tgM96zDxYDqy0ZEg+L6TE05ZszyTgTjlmTND+k
p/SaW5864nqwdPcbYBcVzA==
`protect END_PROTECTED
