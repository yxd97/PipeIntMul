`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9NZ9Ey9GGZUKd3TDUh17+Str4UGXBkeY+o5PlLSIfEcC5UWs+mR+l2WAZ1klfyC
5WBDruc3/gGDRQzH5qsTlK8CoTVPvh1XDdmZ/lk2MqdG36ppi+UBXggx1V3A7A/S
FG3WH9u0u0YzCtnZpu3GHqJFOEFOf/Bm666CgIo1PrPivusGXn9LkU2CZj4u07u8
BMSymop0Yy9qHN9iCZ22LDjCqlAzboi4lceaDQk+r6c4n+JtgICIEpw/+vfpb2Q7
DRpQwvp9O6OA0m22IQiA+vwcmJ7F8NPNK8mraXTbCKmMjDfbu4tVIMoPvlllxo/o
P1/4u1ZU+xuEEM+wRfe6TppOPg3k7gyp48DP3AfpFznfk5bhUCZ/Va1AfWv8GXaO
VGPFNT4MCGApZkEhbYTM4gL/oWXOInZqN6a2iqjaQIQeORfeD4+WSZkBwZ3bsMDB
zyz3jfEIFZ8yRX7c5zuSi71aa7cVjoB7+3tR9aNL5fef+PVgsYM+rxixtGFeAxOg
opR3Y9JyHu1HJinimmrV/1u9eJEKxt9Ch30L9aT6VWURsGyiYHb524ScDTLoELl4
vROnoTbJ6W5zXiK0+2svzg==
`protect END_PROTECTED
