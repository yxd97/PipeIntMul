`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eR2rOS1cXi29KtwqS5QeUc6n5u8C4+BC+FqRsZ48HdTlfU6Ns4e3Hr989AOdGU0X
iEnY7XYLDmK+qJCC29eI4MvoXphNbiqevrPju93uIHCtnaeHVsM6uHxk66q10MHE
nYJwp4PLX5EqrprTuIvqwVpi1H8B3mILjYkDAZqndZE8F97bfhX34DVx5RcdUaGv
F239dkD8WLDgjieTNv+zjhm9GjTIbIlDI1oc/k/hXXvx6bx8CDT6CeRG0MxAsHG0
Lnh80P68CPPrJWLTiOni8JsZ4romxZOzlsBHWWlBieHvMCiYF8IRT03nPxMgVg0b
qNWsLAyJF6PlQ59F+XOj5pQLMDqZzTjCOnt8GTnXUitd5xhKMEi+FuMl55wcXQk4
B/1ZNSidtlbffwTFbBIeKkgrv22RuJYa/aRhjl6yLZX1DSHjWfWF7uclDnRnoEkW
`protect END_PROTECTED
