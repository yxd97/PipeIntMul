`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXQPMLKKcHOOwOVJFUe8DvkL9fBQuYP3rla8vwkxz9MgSyEUkW8UhsjHxFVnFu3X
t2J2FMhfAz+TxD6vHDBFWpHIAkFtDesqQcbuSp9PGY+B7Fo6OaZ+up0mCj2lb8pC
JLn0QpqrrBVYwLB4KAYNtFF5g0MK2UCNFsfwYfh7YjjZ1R+KuHAnpJ+lngRs8XXI
lET5nBQvJUyO19jT3uiVhJljV0gboenvbRndn4VYsKNGPnLgx+MDHejMSF/Z95xe
EkB4vkqzxrH+XHBt0DpzOKNxemRbfT8thTtjqWgaraeGazmYfLEsYt9Or82OcJaN
+1lFdIfyFSBnIIG8j/4LDOF/Cls1qqtwLTT9esR4bBMk1fUaCbsZhhtxHsHJwBbA
tXrvfMEVvOpc2xLP58hWK5LgWC/FhX/a07SkokuQm4nexklaqjgwpq2wdJ+aCZLk
rTef5MQVdH++j6zoTV8+/CGfH53c0k3qMFoR2Iu6E2jLqZuqpHZ6xTyTZ6bjP08C
`protect END_PROTECTED
