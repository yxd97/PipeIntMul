`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+KxE2U6RnyYYiMLwOUUR3Ez95QvlNU+QVRN+kjV4X/2W73VZ9OvEYWLTnkl0Qp4x
IjPPJbnWurAvUgKmwx4BINFd66EuS09r+kXYdDc69Az4wWgoMklTlQ9L0fATl+YY
7TRj4jTrJAKBOxzW1GPs5pualnu4ClGXaJmvUQz30ssQKJSoMR1mFWHlBkzJEJb2
XDH7CAdhPZPjZZw1vSN/1TZLz4sdOGs/68yWbhTOXyge6XY7Jk37VFtN7uTqkF+H
T3A6SEWiZFF7K2x6mIj1E7c9VUEdYeHX0iObP33s+RcH+hM2tzhzl/QZiR5XOBrH
XDNXy35Ouh+k4bJjT1v8n/GpN1U6uDeefOYqjwrSTlPeiFEF3iaar51PIfvaNqEo
`protect END_PROTECTED
