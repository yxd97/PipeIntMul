`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PFvkqKbxbzfsUbJgyrWlTiOZ65hq5hHw406BPnfI8TMQt9kbOeEEW1sJAtuYUmOH
Oz8hIkjMw5B7uYmVhsDLt2ZHgCq3Cw+dNbKrUK6hgYP4aAAwNoqTiyFc/knsHBKN
X+DHe7NhyhRCrDMPSStD14hWWUkLWxlWK6tuT7LAC10euTxsz32QM+DxrmlQmLx8
bzfKaUy8O3AUlhNeX2ge4tb8YQztctFveLAivRggryVuNHmmY6yW/ex/kzzHcPiS
NDdihkflKMfRmo5mucUkmA==
`protect END_PROTECTED
