`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FdW1Chri3gL+JBkiREcNEXK4F0Q1koW0zDE7rtXN7fy5q3gZw7SDixgGr6O0kihy
8MqVg3pelWHYxfX1vS43N4lqxy1fBZ1z/IZ5WEYjvffBKpxfksbtV4V9oImIs0zn
zLN4lBkWHPg13oLwqqXEreCp4M/YrROquP8RmHr2pKUKMn3lWfi8q2l91ngAT2lV
qWQDBb7Vfr6wwN4CdDITveQDybP93bNQO+JAwerbe8GJSZk/jnkXfeFNoQ4fuO8n
//qmSM6UzUB4U4+6SfTvVZDfgw9QbhqoMY2S73TPo3Diqof0kwUNSo6A65yyz/xT
fgCiPr7VijIJ5jRK4u82Jrsxw7Ute5DFHz2ranbRFOu3zLhAVGb8Z9ZrRq7bDdQX
aqWGn2gu5Q6IwPbjTfeeOaW73Mt2UUN8APwIfxo6/gke6pKLqwBy/Wi4FVLc3FRm
ce5920HIKtaWOxdJMxNDZF6NWeSGyas3Xbaxr2t+iA82vIeyFXq6VB1qhybKaWpU
K0qAyPp5rJxeKBUX7JJnVx+HpnLIRzHEcVqkROUhjUmdeLY0L50Sp2Hx59iGKR+q
xQymoeZ8gk0WF8OWPS6tUJvkViMXyAIdC5TNQkDXqRE3x/uG0qfXmzCi14FViTQz
8iwrnzOWEeXqEKSjbJzz+AGE9OlTfOtzg2bNE1e1juXcXkmxSYTYGnAXydvffm1A
kC5Tuwy/zkUz7n3XeHpmYre6GeaVuNIj8RNK3BL6tmK7oIu21LoRuACznv+tBmwZ
CVeCwXOGvSqlcg4b7ydl8feR6wBSXa5wN+EzU02GhhhWIGLkfwHnx3BCs0GoUNS6
DBeyjlXJaLuKy9rkXKkUEnuWgHFsbL6gKp6fRXcEwaw55PE/MDkM6BB9fxJb9p/Y
VUdno3ClefEMon/Yz78v4JxCKn+LAIqqTvbnJDMyLiI63A5+KqS3Yph3RHXvfAk+
2o8dlnBXwa9iKiTR+WLHw50mt28+5W4l8pjV74IpqGhsJ1QmcAeActXuug1syan+
40qWtjLPIe82WOw2mxWJjYX6aEj31BdRafBGf4o+4Kh0UDpMwu8Srs+rnSO1rd9Q
DiSbCjudb4jq09OTgv8kNiFu1wLNkiZhyPFrZzYkGOlEJxc39sx9bQsXgkfai6EC
ucCmwmflrJ+Wd9YM0vEimj9Iqg9ES7pQMThq+fffa9bnFOcvEDmu7HYWJgnaoynJ
PubbLjcZslVP00XSEVT6dbOENlKiRkSsOPywvVM6oah6RxPwY6AFnVoVMWZcZYbj
MxBBjaAaVLZ3n4tjy/r3M6tvq3HUlr3AZkj1jYOKMi7aBEVjghmIZQE4zxtQbfS+
hG3sh2WmBEy6vqqQNv6kuvDJDwYvibRPH0PXhtTNLsvW6UjXyk/laVPM/YY/BDJo
3qlTyFxs4OCEEeOz0kmUHU1B8+7+nnduckUC4kVtdPi9uStboITGqzAYhn1ZufiD
EnNJEzbIWWOzviyG1848rbfHM5zZZetVEIpL7e+0qUqWTKUjwSEhs4E/Tm1oNjEx
F9Mc52687JgCFGxWagAvyg==
`protect END_PROTECTED
