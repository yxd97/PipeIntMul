`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nS3v/bqhQ58d1d84n91FsjYm+F/cFEbgocZWXydS6/fmMQH60tSHRhwupAu8TsET
EIgSGaw9PbKbfkzgpwjHUkyUMdJ8M/XkUY1jRxm8cmsNHlUS26L0suJWj2+Otvx2
yT+K4wiaoABzOtX5ub5zsfGqcqmm8SqQzQqqtrfH5M8K8b6IKVr6n8ldHlgryrsR
ChLpiUDzLcId6/TppT/+yAHDPNFliRy8uKNSrbvY+41OfQsn+3yiaVzcx9FImzDL
YibMcgL8TSpRIKR150SXcn1/YQ3WVH6pg3a3B7/lhrlQRI0nhg7txiORchFusWEN
irX3gsWaVROmgWpmUA2zJpMmTZMXMxVH10/MNNJCyywNj+mP9YmWnzYyXdcyv74I
N8WPpATsUq5wPcUaM1BgfMiBAFlUQDSQQgHwYml0EFiosENBYz8QQVt1lzjBjmhg
Ecc23BwrLsAoUBQLSMgBcNm3qOTKKTEs1B0uao79XC88w7aiAjdfU2xNiT62ZyUU
sr5Srwa/Hwf6iih8bZkNyim1W+XpjEJbwr8Qje2EgrTGEhIilYvHXBGNwYS78WEJ
TC/657h6T0rqAMZZNLQHi1xbXLml+ysndWO8yLmW0WT4eye+oMUQGZYRmYzn7yZr
`protect END_PROTECTED
