`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KOqW1cmDx35+6q9evHBagfZSzgqihd3j+hSyWC6toMjS6J4z0NUwBLGyrtTfrUTX
Nj+3pXTN1N+oto3NvCpIfzdCiNbpaVfqHUXNOG+kBrOre6vY88xhzErJ6y3B0heo
5Tz4ZeJlsK+6JA5sDPhKVQiGAIfarCf4wlxa/4IgjlrXVUtS6E/Xb4MPfYUdFzZl
XngU/ACx49I1VMWsWrmOrtkwgO6UP55hMwY2CJomdy3K2bFkSPbkQons47HdJ4fH
Fxa5kWln+E4FrvIp7uSb0HeSVCXUk16iNaZITXKbWZlGhveAo+Brrh0+YLpaKOFg
bYAjw6Kkjyyo8/AJtZkvExnrOo3Qb3BYMJuftyVw9YNXHfIIdpYKaS+vRuWlN99R
Qsu4be2/CU5G2KdMBQ9cGf/FQSz1HzkM9TjULslZ1cc5k0IUEu4xuSQg/R8Zff65
fBTpK5C9ksBc6E7aGdk9fE/aeUHaEAxcE68HE2LGBR0=
`protect END_PROTECTED
