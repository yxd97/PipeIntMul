`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIHm0v5tgOTwR+0FM+wgcuvxFsoFvGVSffDRJZy2VxBXigBEDsL6/sqbc5+knj7U
inL1g6meqaWz2ClXOtrGCikM3z3OjJc64/QMCi29idOIzjKvss2xL58jkhRCCc0A
jWmwAURwczBoacFZhZIjY8ZkVPpv4ux7PpmtT/mkZDVFibxe1KbFr1pGNgRe1nXL
HpAT7a/kMH6rdacnrYlj5n1gli9Vfx7014dxn4Okrv3tMGdOk3DxXA/nR221rHfX
0AhCYAeWHsU3M5ZNmYUiTS0jN+xY/uwrSBzJceOo0SYZipzfrCsFm3DP6qxcaVMX
UMr+7AQtN6lsafuZf66KOaXIo+q2AoYml8Z1Gt+kMBMMQroY2A1Id24eshZG8vpN
rc5YHdne/xE0m3pccVWAcdiGQGBgGWtYeVb8YWn18amLyM6lZ/viNCUYG9P+qO9x
zsCz0EsR8hY0AV/SMATwNszjh1/akt7jmZydTcYFacpXm2irZcRaBVD36cqDZ/Dw
O/QYE+db1aIpk/D0qG8n3t3ENCGZfMZ3LTU55AuJrdcL/KwJPg4XERMDmWMTWNpU
In5d45l3fxBdjoO3s8oikYVYilGigpOyXZp0zAnm4yGTNzE/weUbhKKD6YkN4E0s
4IJ3h/bcP4bRTSsisLUvb5wc7VnhadEKUUodnDPMof1wDXgaFlhfP2MkiyWGlJQJ
`protect END_PROTECTED
