`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JT94LGw0xcLeOeQlK1kmklWsTrrrIdjVMnl5XWXnzsdaVYD9+JYODWUVBDzNMqTw
BX8jhWpxAQzyPTeyzKfpmRJf9hm66H0BXsIB5pGEZNNKHIV8sLZoJeXXcxrdSLTs
S6THTB883KIKiQskuM4VeHo+sUtWum0XEMPLDb+E9c1To6IbGhpSUB47/r5yP+J1
6vUsYM+rVbX4wTK7ACkX9ylwYPFc/VcU9BevO6KhhRpQS42FZysGeb/QpNmudOta
1gFTA9EosWdQO4fhRuBNUpMR1T8Eg9R+CG97vakiUdPVv8Cec+a9RGLlJnd37hiu
aVHuffLEi755jLqPk7aawA==
`protect END_PROTECTED
