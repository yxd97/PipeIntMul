`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
76DI+AkNqputHcyvgmEQty0OF8WqjDb7aWs7JGzHNkoy8n83hPKq2GYq21KA09c5
6QxMGdjIDmcESLzyFglLsfj3FeETxoIojdcZITngSQzRAsdiDmJIY39j3cRyaLOQ
2355UXGXAe7hwMI414sx8OkLIzx7H2rxOJQgkbh/zN+h+IZ8JnTrf5nlhkQrq4gl
uBV6w0HmtbQCl95VQ0uK2lneihiBr3upn3FHpPtpVWEzjVsJ9h/auEoNnu3mOw1N
TBZjrRpm5HxVfeA3vo4TcfxGe87OrtDEpIhGjZY9oal6CUyO2oaI+5FODQ4QyY1B
dwmh6+xdBBZk8iC6JJx/jDfmc+jsUDwRqNHiy38qeS+eA2TD631PJzOD1/G8GhOv
wh5UwYAPMD7JO22TQzAZwNlyvlktQBmVGHrUIx6IiApxM8X1p02WctycpgoRIUO9
SvlbQoyd4P/HLUFJsKx3K6b+0UaocliKQZWIbZPu8Jj2Gu6puHPWwXeYqhKqDkWn
PoRF6c5iE6xGpeo1AVI2PIfORuFK/XiNFWAYMKFWcX8=
`protect END_PROTECTED
