`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z+7zRmht0jxGfbkUsKc4u8c64CefSkZydEwY1KdTTyiEkDsDvHsdoUwH+xeMKOXL
s18Dbb11tCAYAeMcPPZWLoD8tEJbkyNyb/g5l55dd06nrRfusHXJ6iLUsP8tZToI
iRg3Znh5moVGkieTVGapWJogkiPvo2t7ViyJ0i+mWn/OSGpzUbraUHKAxta/9qtB
ppv1BYzOeigMV1/UlXR0pa2ryhYHq1ksFSbw07lWezhGqFiIWpwv+lYU4syQ4tVC
FxVn1YcBgJGQU72G7nJ1kjc2rC8YUM00XR4NCio+ehelTiaLOCWfJwAjjpxcoXZW
cE8JaEn6uMZTa3ifxR56QaXjSDSz697CsDRVvVswF5aBPGwqRpGNs5pqx9ekTtPw
RQY8UCCEkwMa6GmKJKI+KCQ9ujycAd/7uAOw2AZu2SEMwdlv3/t4XQgKdvXtUBW5
bcFPgTWCxTZoVEZlLHlsdV7u2nMnUkwqUKywCbCjxZlRpOm2dhCsQ/vuhExjM6Qm
`protect END_PROTECTED
