`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zwrHRK5MYr4UcfPfxlePwx4UEQi8LtVOVl9rw80XOwLTSAKZuHP3AskyzZ1acvcf
m4VPIuiTJR0iaCKXiqkJW2oe7jrNtEthkkKpr8Aq41HPLYgB63p8XaN0mmIgi2Eh
gPA9KNJBaNismxAZQbhepwv1ce03mwk0shSz9cITdjPEVZrZ6AuLaR20LJouN8FH
OgfKSGDqY5B9COycSb6hjzU7ONV8XaYAM8HgPIOK4219gZ0Vi0hvuFJituo2KLaN
QVjZr3TYblSYmwSro1Nbdspto3C1lDlnNpKeedz3KneBh/QiZi2bCgOoXk1MOzuI
h21Wson3YWMgm3Fqq2FFZHH7N5KPJgmwQgr6uYrLoZ9Jhc4RuJAM8+re6boQVaGL
RsRnTCEVOBkutGy3lIKOFWWBvQNItB8+Ot3j5V5hhsm72jYgmNOfuBH31ANvS8Aj
WUzB2WyFU83XeSlAWFK0UEo+dlPPXGJvgm9r6QmL/06lOwUcretijdjPO7lPNQbt
MEWHSngu6Rro80oKMrxcWq9K32dcEcMFBxUaiSwnutfyXIJ5DfClzkAlncwVljoz
1bTeIIpIM5V5a0tPm+oNMmRQh57rqnA39C5mI4JAMyc=
`protect END_PROTECTED
