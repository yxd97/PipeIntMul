`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0rB1g7KwI/EaMUIr67K22EIgdXUZZRLzBuKJ7bbkPj2UnuFTKZy1xnZ1DqAzyOMA
qCIO8QcxLschaNb1t0p1So5G+TTrrGxw/MOs3ioaX/mIBf9zuFRYC0GIB8HLQIAM
QIBqsY8KZgJH2qMXse0Hc+P8NJ1u87yZdqvRrYIOMgTr9sKAsOaKkay28LndzMd9
oz2ZqYKM4NTykPOucn5NVuYp19UrXbz+5dFEHYXqXIdehXMaRaZTuIKqN4VkSxXj
iE1kKZKWSRibxkNq2/tcz3cNnoRtCdGHNtncixtyUe9VeyuK95BczkMuNZRgpr9G
vTWWJ+7OQnekYMl3+Pxwcw==
`protect END_PROTECTED
