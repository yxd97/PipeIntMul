`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Thvs61yXM56EPs3wCLYd6ScX02UqDMChHhTFm+cHMG7hPFb2MQDIEJqWQxS3Eo7g
ZQBtRZr49IjoIHeWL6D5ZzwtWpjUH+OLwxpO5Ubp2teq7cwZhQX8nF26H18CUfw8
HwLvFJ+Ch/m8P7nOG/lELrPtlhButUOTmSbjLG8WcpHP1gb5EcZkcLHoB4b7flUn
va+KPf+p3free9HqeBzHh7cqZz2XbtqO5i3LXA5zRM5K11cR7a7/qf9jTRAFdRML
+4Je+LJeG5DQJ3SbrG1sTNUQ1px04RVI3meyHGZx4CtvIClJyz/PAi5JBSdATqwb
xSE+yjTacZRvcTr3SHMa9BJ9GY3rSH0aeKt5E/LYvn01hM78vwTanRMJ/M1Mz2/8
Hy4gV6axSPChhlZmX2sNoIkO0uhUeloLTAzdOJmLnqnL8EmkL+YzW4g9+Zc5FyDf
7Y1dQtWSsBiuXhCNXlPlEADd2U+p5lsHdxmwJ44FHMjEeFnBVq61CLy7rkvCbOsd
h9X64Xq8mBFxdq4d2RF3yPDCPKX3CRW/eCBF44kb70uStyQXpEG0zS6IOgWu78/4
JKMkVtdeO1uelda+pKeGgrH+lUHGHysUk9y1TPdgUVcG+jm2h6+HXx44Fdv/NM6Z
TC6ozhSWpH3WRPteY8iUXuY+wgT4VxYVrM6OFnIxlKo1huLMVpsnznXpLf2rxWeA
3EQK12nvYCc7cKBaTsffuJUtnDpm0gRug4X18MYjhX3ifXdUJG3uUxD5ARncsRoR
nt3kdn85tFcn7/6ta49clC6ZqYh1ICc12lqcKfJpJ1iaNGvnoavw4NszzNgiaw6E
CupjAgw9kHcbsbiLOZQDDIx3YuqfES6N+ufATogPzyCRJHmlHUpaLIRTRVvkYxRd
2x7sFK7/YjVQqhLykjo6eSJ3KuTkMUpBBjk8J+P1ijfxaLIVTo3aO7uxRpWIW9bJ
V5emXsgEYQ/pVBBkqkzsQy8P9Ah1qGwRbQe5W3R3z37cjQNFc9xAa0hDk6VRc6Vb
tlGT/aGi3Gh+L6Wewv3Krf0J008u6cqrAXQOfl1y2ym8eQU4mX16jPOBiApyHaZ5
DS+wWwcl2O5Y7GAI+r7qjfv4oLMs6PFRVeyus6MwPoOLW1e9UE5G6duq6pbLKsA8
s0CGO58AHxcP6w3TpGSUy/1heLGS0VLA+/iCzI8xceds/ak40xjxEDFniDCKuFjp
6qsESBPAwKfY9/SQ9TAhWQ==
`protect END_PROTECTED
