`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xlx+WpkUTbbap66QQg5MBhOqbDQPxso8kbI7XQ6mK3tqH4ezOQn7ycA79te7YNJ8
OO9GCmaCAxRWWzEQsuDdp17turwcGBxTPCkCcxESSgJGazs1auC4H08Eb66wzuCw
AlYk5/PP8MxF6p9ZtYGlduSTyTjYPEC1tJDc35kUM3C/NPLYMi/xiTuBoXQRjfDv
r4yl9jHg2pH3wlNew9Yznb0yxkRN0jgASUFWpRGz3lhoJepTPIrS+dzzhJ+EJYI8
NnxzSjMysR2eiRrT/vsFfglMO879Jfc/5Xs0AIQkLjHVylGM/f4cKMLbFuWW76QN
FW5k65BWbkyTtqa5k4bfBHJwcuu/fS6y6l2g/ZbzUW9BzDu3xyEAhtv77ia/giTC
TtXZjFOoyIw1jbD4v2EbRtsFW8gvW0xtRBHklKeOkJfLAiIPM8pLEcnUHn3IKH8y
0I7eR8BClGjp26QXhEcw5GzxQii+l+ZzBDh3pbess56vDsb9hxPuq/QVFsF9YAS4
zoM0gH3i5hSU/2LIfTXCgY0WRU6Y2ZeX52j4RrcYJuqMK5i4vBTXHQrTwYyhX65+
0Id/9GxKxL6qDdZ5Dq4PIa5SlF9+MaPH1tNtZpZCUImRAsKCHKx6zfpZPi5rOQcp
jelu9gFSEWqrNdctiKjm1rRMZ3nqzvCsUrFUNk/txlkvYK2mb95tqyfo802Gs7do
GYPW6HT/FehhXLyukVZYDGDlSJDHEHVTlM/VSWFxw8h/c2yGuVDQZ13IUd9/vR0V
Znc9fUzfQJZpEnD9sY5R/1E8ZM7ZqQ3xScSh+wN5Icm0zHFZAbDSY1DPTJJ7EMMK
uLd+P+MmzEmZrqUb77fbzPX5HDCCZPttQmnRBPoJ9cgpQKYLVdr4muPzfvFaauIY
I7cNuT/akhas9Hp6eYrue2pKc1rbrePxGRNI3T++GmGZcvispCOjti3oLrrKx12c
OK90nzLewB0hFSASy6ii0MHLuSzOo1MxMiEuug0Qv3M+e42PScTay9rIMr6mQrOt
z4WQtp1zT9pQ7QeNZ6w07dq08BwXuiIWC6HLq8O0rnibqyWVdqp1C4Y76Wr7ODCz
CiUHHlF0SWdNsHonjInSRWdoQIG7bCdPjRjvu0OV949+EopEySzM7Nojeug/Raog
OqRtNYcjifK1n4PhDKm0rpGsbQBXfE4DNEjYaeSa6mf6Ag0CezH9k1g5tJjhPT2t
v8BTrEbJ2IdUAOcasuVkLqVnoZJfFvqeE3LOQ2IZ30D3+hys3KqxTy2lhYdEwnkd
xV8c08YDbkT18CvSjKibSuG6U/+tFZRvzV4Ez1cpxHVEHik6BTzDlBmDY3a/Zfu+
l2cXBpwSOpQl1oPDYjP89cxcI9SaxSsIu+ioi+H5kjC1aVddoOcWuZcJ8hFpY0yR
jLc1Rd4aNG5Eyv9JvXz+puX0d0odm1ldlBGgPJPsVwCCswJyXMOfZFJz6R7pMeKy
nSXQaBPMB2aCe4m29kkPEgUzo4L9IayEWBtUlsNJ9561iAUajaosS6d0ODnLrFhk
xNJBRFPbpoIFleSvkrzuPlWNgy1JEggwLRQhXeA3WeR38OaKUlyq7gPr7ieRaFdv
SVMGxppB7OJG7zNCH7GIEInYnJglhGVSzVP+l8+fIh0b4WtzvEwH2djehzgMCXVS
fHN+D7cOTLDWQ54qa6gHEIr438gN3LuYYHICgrl9eeWVhrEVZXJ2QhZ7YdkCPNOR
EujanTSf57Z5KW8dHg+U2vpuFgtRMqS9Pwv86Oh1pi6dtb2fSxFaeGpASRwFhUSj
ifhQforZ6BODamH2cuYuBCnPBMWqqaaBPlXxszozOK8RP5Nlz00pQpF2eVVg0aUW
9Et0g7OtIfEi60QupZAcLOXaetUDKcIq5p1+RNt41WLX69LcYiBGIptAMbQNxwkI
m6IMWUmE8fXwEw6XMedvx63myV2uZ8zlrXs8Llihr15uOAWL+u+/EEufh3cHW/x8
ZzLBnVcIU7XVecRjruRYezwdVpIqCCP1V5xpG+cmeFPFqk3029nWiyStQ4E613sz
FKjVeo/AOR2Yf9XWD4j/xx6ZkY3wfUDBWK4c/gtEgfoCJou3AWif+ZGyRQEzkiwk
EpSMOmnjI5RUbl069qVTf9n6U/A5VYsiy7C9VXchtxP2ma8fN1SQdaTDJfVuSSw/
PR6GWC/5dc5pYXJUBr/KhGlXHyRMyEU4Eb75oko8qGFagjb/udGeus4Mrd64nr5y
ATpVVrwXrRASgqdNcugqNRDuDPq8EpM5y6n38AnsxTAfCewZvbMae67MMdXeWX6u
L79w4a3XWkw1h9Rkffu7Og0ruirWgYbTBEkW4LXHYlRvgsR5rqlF6Hr102SSKPsc
+/F1+t3bTkKP7DF31gkR9HTwNvWpXGju8RpTUsl1hpp7XL0TALmzWWXZ6AUbIUIA
l7Z2n5ktRsH4qzd7n8SO+K4uvWguU0FQV/XptVgNdsiw3+YwvMoJM/MRkH0zsMR7
jF+H7aCfwY+cmbHSJGCZd4JINW5KoI0kOx6GQ2F8LIFQsS3sgGHl/bHeiBFDIRkM
te1wnk3D0O9lx9guFxgMBSOfryZMWJPGj6juKEZFegV73wjrNm5Updtpzb1DLUw1
geggfB6AmryFc9FKu+BFqSECF0IqzFNdaUYHM1BzN8JS8sFZ+onuhC4QKWMJl307
7x+OTrxBRjKC5Uf6Jfw+wyK+HLahWZGufIXonjP/7Dtax1bhzjHwFrkHZ1WQl622
dU6GC3rrny7wMGrFQDEbU5pvOuYa1+p5g9/AzLX/4JD2Q5hTNR90LbYP1ANJ9Jc6
szaTAEmMYUfMmPEy1BjoCbU7Al/xfIQ9Q7PBKoEe0YH2/JRDt5utIu+5Pna8RfW2
hgniTl6GwgwwA191ayESMkTz9ElGbMmWy9Ph/Z8M9YEVkyNktJrM3/HQ27KjsjAj
BVctXu5aKSJpdc06BNFPFfrQiAeNW8gup8EkhbbmY6CWLO0B9ODaDyMT2+a0Xo77
DYhQ0g3ERdyFXZAv7d/zjfJaoX6kbZOOFssSN03oYsCGwOiIU2BmX7PRNwknIe65
oXQrC+Ji1iQNtjnwo34D17CTv6QGVlTniWZbjcn5MYgTUOrccGR8LOtNjpeXsM1/
J3X1BpF4IEqNy8bSu4ecul5UZ02Oeyyi7RKvzkstuT4acLerbnqzwx5yB30mPWNC
Nva0Swl0Z3LBtujV78N7KsJC1G2Zr8hivwBNLOaE/PxOhSLopZAZYjjXgCqXbU5y
35JWMVsNSnR6zwTAlfUBvWHE+lMUFBkgL9p8VkV5QgPSmzP0/d3m7IzvI3t3uBZf
FIpC2d4JyKzQVVgWGbBAEoACa0kxb1nDiDFRAerKyLEmtEzbsrhkBbUDo2txqHnv
jiyEY7myw5MYeM9i3/zLlJIrp9YOHSUYelGC9vqo/M3fvtexGA7NUya1okjItRQ4
Mc+2kL5vJdaV91hANX1nOUNS1kEADo0wZN668TIwt4egeubzcgK69ARA2DtwcNM4
Z9BWCzjr0/b5lsZhAamq+iOVirCPTeLIlZzErV/SANhFyhgyQ5YgOKymB8wNfBWL
7gnW20KwWyqUUlGRGX3u9FiYwiNuQeqzSVjxT0nQ1I5hkcpqyiNEmrN5BXL9y5j+
MfLC7xg+v/dLiNLBfNswo6ka7gZTm1C8j7FziVtcIUmke5qWiNDjMxDT7RyFCAyy
TSs6jhgUJ60kYd1dDuu0bMTr6I2wscA1zmZPQOoA1KHp0si79tad6h0vVh2vY4FH
cFI7Y/9C1D8Llg7x8wAveXCj7yEV8fGfOQF6k2p+08VufaQTTKZeMZEovi7ortxi
xD2pe9nRdGNMZ0997pRYm5d8rjAUVdo83ehnuxIEJDcI6hbcxjkD2oVtiVlQhQeb
3tY74NsZP1c8nxfmWJ9TA7x6nwlyI4XtsAL2Sa1bDGgYsv2f5u8J/IGSnasHRsvS
bcV/RXT52shJwoT9mbDfTuHVBjPQGhLVKVB3rProMraBzbeqZEWtUTryJKV1lB+B
DHKQKqmbeoAkTQPU3jkNYc73Uc9RA7C8ZNRK/S/29VbYRcupahzo7ZCG8vcTJ4aE
VgTdiSHRiSIx6Oly+lHiWp0ifFRkPP2+dpeIINudAa7fzVM7ZmQUpgC4wEfKBI1X
wZCjuNVh5UXDx5vGgKDoscbwDDngfZ+WVGVkNQkBevapTJgxMKuzheqQSeVaC8Kw
PVSJm0qLivXeAvCs+cE74qEwo4Lfmf1EPNZGsgFzvhGgYWa1ssX2Mhc8xq4Zak/k
DSGYuqPDWLKhUtKPZCgrrnkePrxWbu9YuRZXvR4CG9K3sMZvq2GPpSNR41gDt/GY
xGvaKg+R6OBNfY4rghb2YjHYGG5GR+M9xVGO2gcNGxUR64sB445vCfS54MAMkaP6
aJtjwBSBpcgEgrNYUVop7/PMRk9oRceZvDE7tP1bmNde1dvfqqyLkvE6oJGWu0TK
UEGTXDnTjysdoex8jLrPepmmvSEDgm3eThgVozoOnSwu0PkwWoJqG4ulEzc5paCY
RY3YUCHmbm/zcyfAf/Tu0D3LebZr8eFVqUNIwWQQh6nphbe18hlBMLBD0onL2HjO
Qmomv8+PNU6jxlbojGGGaO7V4Bs/leWUFsImDg6+SgCzPew8bIl7VFpFLaJK9lkO
F/mtboJ5hSb46J0ih5GsMTdeVFt1ymtGlyBBmvG9z1bit+Zc5rVb9Ccg0mxrt2Ej
+7YRkoxN9QwC8TSPiAXLByetcr/fCffJmY8c9XId5EG5R1RvwjgYZtCp4HwWmSfO
qLwotn+TDJdITnLJUqfp+Pw5+dXVHyYH6qy5xrBeGrxG1iZDH+hx/83ARi4XdvoU
91xzTTJ21EM3nifgh2PH1V3LR6g4YOLXm2vTdedSx6OGOaRaOjM/AM9g7HQssc2y
kKSrvMSo4f3j+IXco78HZGEsQqPcik0grANkJdZfTVO9Yhf9hGEuDNTqQT31KEdU
HUU67WjGOiNlidlnrofFhuyPKKIq46Kie1HGaAVkPdHXP3FgXMKVfH70hEajSHTK
tvdJ24aPxFOrS4H2QOtnWL3Wf67FuOnctAU4LV021lDqoXaYfFhPM6MAq4cgmGN2
BAgvIwwRFTE9ulrEBhSvxAjiQUyeZaXtrvgpiAV/sVQSpzVfYqEs4ufctyX130tx
aLMScvjwhj60Bfz3/ESi8nNz6aNInGFjZvrRFyM6H0wDsO5ux8S5NIFCDtbuzOkM
rmJrUNeT1U9DD7HLqcs0Qn3Z/ZKz9wJBZGa9A3/y/KseiZtFoJwRlGxGIR9b8Zpc
hlHLXRvomfmRyo5NeJ/TTsKiJeBF5mKO57O+gXYe680hRHBdq9Q0dObCj0HY7etk
1lAZPDFp3YpXYywxOeVS0qAfk6zOzmXP1qT3U7ZgCXTRs8S+cY+7QPR92TjnVeoA
2H1CQcvvUGdqYyLjJHk2nW50lbi+SJ2sfFgKtqFP0BYtzUJRAQfNQftk0kRW5xU2
X9rQK2HE6v/BLSONh+Z+OB5B476KQUvOBBIFMtfwIcw5YScmFMsRIAaDNwVyjH+0
kY8K/yjg0zQiN59ERwo+mtynUCZf0JlcG/LIqatvCzK91+EZdJYB+5MQBZsxybEG
w6urjlFOgV9Vsir2qv5AnkvlzuooVcsZGuuOB7ncoIDJVYE7159yZh6AtaYwefJL
lN9pG7VaDWA8asABNmSksH90te7bQEp3MoJg07xEtNIOEa4s6xxW3VfzVUO4bDao
B3Sp7vFpQIXJK8yC4huXlWCcLD0L4GjMzHPkPzpt/9tF5a0xqHvJAH4QnnOAZ1Fr
Z5pcLHqgYEjL7ADsczsj2hJTyh9ehGy6Fi+ew94zwHKN0lnUp5CeEp7JCZ1dAVPI
skIbDiafO4x4BLpw4tU3xk+TJjLhKF1SmYcY5QqMxCChmFBnUGN88GRVu4tdobrh
EuQtgh9hzWmRLVvV1iyqnTovnRaugYocrW2dPHynyXDqRQTfcyaiiCAijaG8iiWz
h9bf1imKw/t2V5sgufS+ho9CVD0TjG7+2iu1XBfq02pxxSJ6BccErhS9flVjcIWl
GPrjjqtitiFUtT2qrXUfwohBVzA2UDOY8KTSWs1O+5JnOuyF8qiz+63asM1vNgNj
R1kmAmaBcVf0M+tI9gXugRj8hvsFhe/wNqNFRr1G9h0dHT8hRcYN+yv6oEhjtXPQ
/pPHbd9rt6aUxnbtrHrL52wrrw7A8eTKWyq2upnfo5tgC4G3JvM+TSry9Puk7G8q
0quOkaFzZtDeoi93kgQM5EnpyxELdMhrId2IGBhyHWJHqzxjR8A9KT4jqrqB3yzO
MLchsZcH3FF/+nRNzNQNewdurzfFdGstQ3gTYb6DMOefgiaxLsfH86wM7gOdmtrC
55dIETZcTh4+vq0fXJGxn8PEvF3cGUjNT0aM1W9NcVzq/CJemf2C7DT8ybslQip/
/1ZbthIXqtQyzQvhfsC0bE80eflQVg3cT6eAgc3v3f0WCgDtNKOaMq32zNcwxv9v
7Dmj4I4pSaPBaIRceLn+SU5vjPjSy1OaN4hEZqSHIgXlrpIqQhGNwNadz93bBMHP
z6PRMBFAqVvIKFnhuCarrv5gEO++sPe/IEQqRgsIF9JzW0gqr9FAmlLinUlouobv
pkxjsDJvj2lx2rNf3JZMv22jFmuYcIkD85hMO+flJRscTGIi6dFeao0wn0jHS3CK
t16C9NujD4gEszcaOIyBg7K+2WyhYAMQG+Lzp0vl0HOfDh7k3paUnAvg0RrcrRxt
J0Iag59n1n1YUrQ91NvH2uLQEGuXPzbI+WTuREBwB8/oDmbL/2PeD9Y0nZ86mI/U
vfRmKuUuEZGL1bZP/PUiJA88yCbRpzucbEwRABnZqAwjSSE+t/c3+VMdyPmhDly8
ZSCsm5GOPVzKjH2biZBQ+jDcXI0siEvnb53qWD24crvcALqHFqomN/HURnLtOiNK
yoZlq+99vG5BrGEJkVL+6Omdg2FqY/49fihh09vS4zcTYI/ohStgksuNmnjsmq8O
Ppy9r4rMbgqEBkYG2v7N2L+7U+1H70VwT9v7D6Np6eZ620zKpspZpTJNLs8U4Ckq
2B4LKxqMARuADvQ4xlm5BT9xKzyQMLMw5UWGDymn4S5dBTo20VdU14v6Gtcmr1WF
hDeKhGucy8mTncZ2caRf5/Bm+5KGeTYmhNKcVfI1epIX6YRvBzKCdEceUdBcBzPi
lNWI4rpJy5IZS87018yagJ4qF2v34jdyWte6Lz6e9q8uX2cm3/wOea6plUaug/AU
FEfAKQ7CP9+MJmZz3n3f+xSsvOpbN643oIalxHaCzvuwj35OW5vxqr2PNS6aOhL0
Oj37Aq1UtCLS/dLCtYI9ZQ==
`protect END_PROTECTED
