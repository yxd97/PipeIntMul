`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEBBEbLpsIU/yBtdocuCvN3M7pQLgXMtZRwB1dnaS99BkaA8CvCi+wXEKXKK5A9s
jasJ3PeQrXvDnZvv7H9JSv5ILLjmaxoqVsq+GL4frB3tCY9xS/A0CQq1iM69PpnG
i2AR4su24894eETMN3X/zWUQyzOCHV7i6xvQDpXgllDqD7Buuw2F4pW5UcxNBnsc
S0iSolxnUYVNc7P2Dofjya8r9sWACxTSj0xyo/DXvhXEsS8fpyyyfg7YNFjXsCH0
JBPMFstM2B58331EMjcjFhnclP38DsLH2f6HsRa1ozsINHMluZ51+HU85hFaZKW6
v+uGDaUzTpnJTI0nVMbj7yCt6a4PNtaJux/vfAK1PevNn7cmQtJFSX8n0gYT80V7
5qF9dqzEFOUC8pLMCkyBh+8vpDh37nNVW/tK7wIXre5gbTT0iiE/KAhbSE3wQCeH
PhDdQjmwNUeVISScrgltfG96t4m5OtTn9TocXwF33FlJsbw4axzRuHBkaqTjfiBy
2BOP6BE/qXbPAbDLqEScaC6+Epe1g/FYZnxYzIkwVsrHo5YLBvkZl7LVJE6L8UNM
wDpjDLy01lgPFpIirHb/IMklXKj+diYEVstL1OFSJMlcFvZ0JiToj/fLe5Tv43S/
DOv6RKSz0BJfQP993L42rhgYZB30+Cd2Yms8k5Fr4uSF3vWWcdNK3kjGDx9yNLnP
rEagdYBxB7F7uo54YWXB9PQDV7wod6E2DLQ1YEKJ9livkQtwr3Z1uKQMBK4iz+LD
QiT+CyIzYQ5PR12ik5c+DnfIq7/Zh1AOkAFev9tHBztrPsS+I3GNtxvL719hi2GC
djIA5SjISzQ/GIEe6hT1VSZ4qMmDCbzg6Gexh+mNBw8h4PlM1erhGjw2ICcu9mOM
pSewLfa3Z5g9Qod9MMJi7g4NlLCccjUgZxUSOPKA6kWDQJD/5cntPXVK2uwKEJ4j
mPZZjA/iwbtItz2vXsidKA6nPpmVp5jk9rQ4tEIfTZqVt4S0tSfs8QZ/fi/5DT/d
fWnttMtZSlRklLt7BIGK3POJoPzKnysTdlmDwac3PJ8B8Q7Y21it8W52k4ljVVsj
22YxzCEUlHPEjokUEgw7hA5cV/X9UqTIyAx9TmYfFYhnK8OW320VXN/H0nIbe5zd
yDEgXmHwjHHuk7nykBGkTzDpCYBmNFSe3Hy696iYFbh8DWbikTKypXQTaoCJVmll
2m5EpLNk2qru8zaRjdkIzn7JKnDPW4ZIO+lPu9sC4ZiSerdX2q8XsOKFfTr+iOra
gpIRB18zbRbuKCVUgkz7x6uMItZ0T+suSpV8fbxFbE72mqFv/kWcHYuIJTV/frEQ
yTlJpIu1/t+iKutEUCmV9CRmeODSi5qzP2rI1bThF/OurcQh3z1Y7LiZECfk4riH
EIg+EzFHItmnZhVvJV2IaE0BAaTAPQJxohvWM6HcVaQaVi/Pf/lGVoxqWfvLrmaZ
b9oM4ArAkf15kcZDyrMzEdqC0kGJtgfAXXvw9M4IX/oygjXXvN7mDAlWyhwQnykP
FPG6vBCqJJE/kITrQoIR3FaFRdWpXf2lb7k0Y3axan3jvDfjbt3wQcFsSO3PseF7
H2Z4hNQx1PCZHVJPex3seYHw6wfBmiHv30nR9IPi2/qBjSYSAO0+AGbeY/H2AJGS
+4OmeXlkUqdWqr/dP0x+S6f5wqFG6p3bmEHUBTOTA3C5uq0XDRww1OsUJC3+teoT
mZM+FOM6HsrftL41+LL0OVzSsxwUfJMRc1TDwmsqMp/bn2R0uqpIo8JidpZEf8Wo
E+zauwC2qbaqJFIAw9q5q4atLD9+HF/EXMlWUOm9xyftUxA3/DUwPEmqu/kZhLa+
q8PmMdZJyoFc0rcHX17HgX2CNazA52wuB+tYPQ71bE+P6ZgQCKBV2peNdUw7CIh9
uepIZ1QyFofonjoPQBU0ZT2x/hNXu4qOrloijLPOaTYjh4AOmcPQMgn6Y8E/JkAe
//eKKs0XJjOnk+8Q8AlUVLiguu9l5sBhaQ+bn0HpymyG6yrHaV8o1+p56Ro3bkmK
mvY9fhXnmozoYjgUobk2PBqcdVu1KQHE4Hzi16ZtAnnPOArq2GHGPhxmjH91MgKP
MShdBZrUcnph8OSx0xPbAFNgSLgt5klzX0g8idHt4y30+0ggAXaTJg3o0WJOOJO+
hFTW7DOnFWk0PAbhxVD2JepE4bnPHH8XE0RXhrBUNpQqIRrYbZ6cGQaGZnJkIbhO
Odr3/GHvCsHC9i4FBSPZXODzIidFAX/mSAGHKVHMCMARt1/CDIGwmvnSS6oabR4l
Mb3zvrAIo3C3yP6RD979y8NNt0PGzdVjQ00nfO1QCHPff0dhmVY8BevXIYqr9GBU
55J2PSx+7ocVhGa6L82lrKBTyZOPKWuyWx40G/pp6oiXp3kwe9uogXki8LO5lz/f
NXvgCg8DkoTgLxG9Bl7WvrecED1odM5p02P+7diO5zFlCCyHV58F2byAYcAe2NJ0
Otx8j3UFOZ7etk8eFLrWzPYYeFEqK5u5GYf9sR55yRqz5PHAHtykJ6YQSHdwHkyJ
DnFx2h3XDGuJwsdOjIMaczmPM2J8z+8nEl4jZ4MBiIf8ulsjoEwSR6TZK+qbhfXb
vMvys2Vy2g2+DE6GHiejcw==
`protect END_PROTECTED
