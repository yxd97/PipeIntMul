`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
025lPRJ73jbVEHHe0HDlCuYxx5zl+a0g2fB/r25fQ8lZKffUxG8/LwQghvuwH6Lu
wQmdU4YkhgkWAm1uhzZXQz4cQMfhiChxH0SGUQMvMAcISU9kAoS51vBc8aw/hAKu
rDYihqnR7zoi1G6hr6oRuf+vhOrdwcho7ipyvKtC697bEwaXhFjRk+UZKnAdMAL4
ho2OY7Vno34a48Vf88OcEJHNMwx8aJlYmihBmWWeATWuiih7L+Kfoej31CX/idfw
TzwiLyH6n2plZigAIPnyylSYcI8LORLpXu93LPuAdV5ewA/0b4a6omtzJau7V+1k
habFJycZCLZvbAtCe6ZlPge1bmix46yvQefnEAeNTGf7g9vavRb0cX7FCaZ3snW8
u+l61L9oWCMycwcXb8NZGSnUv4Q3XGV/oH9CnXY+YFnkpfyfFrVdwjbjDUsACERM
2etvYMH0bw/jcxYBZ/TT7XP8jitJAlrssUxsupBef2/xjD3o5og+qSVDDEhxWCgF
NZPRa0S36vpPhKd8F4E3BVTPFNGfaYTKYhnlaiTmC+ZrCyr4DPHDv6V3F/zzoXcI
XG3FAFk73k1yHtdoNUHF3casxga0M4IaAi7/auYkof+HY+m4rQ98bxo9g7Qhedn8
yGXwkeEgkCEzPgUuh6pxnToHeVV8sKmyA/tLZcjdbQ4InRRKUyx5+OdV/bkrgnpo
0i/pLQJOnVEj+fC26XK2JdTaukhd7Bd+S6dd3DjJ+hT65x6E0VHGhqt7HNn340ak
YLnX/m+WEZXT/VEWH5537OjZGKq8XsN3rdB/gcrwgScB0XP7yCjBxFF7cyQIpiux
n0Fb2SEP6r8w4dbk2WdXZ9adU+mM95qdf8ySvFs4CkmA/PukIGvqLGcUA7gPPrQZ
6WCb1y5WXiSCz9+5Yob513fjy3hNQSSA3nKhJ2UP1wVwL68ZREYkMfvMh2aQ2brv
ltvf8doA9wspdXv+JpHAuhg6QMjTylpSLWk54BGppNjvwcIWGueWz3PMHjDX5Be7
TBgJd77uflQtskWq182xaW75LlCUsKMPv6ymHVvhLnf3T3Hn7cTYH0upCgbh8Ptx
eKGlH7Bmdz967oD8Cv30qFFkAoxnZUi3k8nWHWNti3dCkT+Wg8qrytR1whiWK/Tv
2PL0kL/7J3dSK/2qSDSQaUlvK7Mr0rrQoGiR9nQbdYLYIryoQSAtof7EvqEj9GoB
BMCsPYiSqNvpP5CdXbe3ZPTUC2eIyi3H/hrwn9tLr6SLQk5+SldN7WTsiQz5+VVt
pPhUBfyb7tfoqy9+cHi1aX6sRRtOe0yWPGYsHwjLrG/RbcdaI0YlExv4o5gFuKVG
`protect END_PROTECTED
