`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZLGYDKusApXolTyq3zA7f6VcG71eHS1F+qOpuSZqw+Bq1/CtMFqwvyZwBZv7kt3f
X9ERaCylxt36M5tOPHbOqFLoAV3Gn65EpGBVOMgwqR6TFrcPgtBQlONbVTFEEwBP
1mHcCQE1AqKd+DK7LXxP+DzoXuCi6dhL/PfTdg6I2nSqlqKoyra9iU14PxCSiNjK
gb+NP8mkySMytR+0breQUi3GnlUbBbBhHJ9xlWwD9PZy6iGa+SVFrGTfoTIhrFS5
5iOJIPj2MhEKF0pNLPxFamZraIk3/jRoIIdU95Cpx6U4YE3GQh3lHm1XW0AJUIex
iWKonW4eZtwbOEERmDe1sj0qU5OJQfSh2onBV0lesSSU7gDIkv6jBqrT9ECGCAm6
6VIbnmdrS1HcGqv6+ubKAxmZohCSGzoxNEVSIAHjqwdWuNLPA3XLCa54d0qbBWTJ
Dqf2CVKlRyGwQWUW1XMRivk7ESmrdblXtUGLYzCMekKrGVkbKf/GuRiB3NPQ7mtd
6HhiiF2GjWRzEaZTBClR42gN0AHjk8bowmFxl5KfLFsQnYG1KDyagr0PNxkQxNND
VNzZlfuoJrcsE+Smz92eLDS3E4exN8Hy8FFkKDV8YOBE/1EC1YXHrduvqTD33C2Y
ZTPpd94C2gAPM7K5uOA5+yiGh0DsIDB94fMrUP6zKOYSQjyjjitsP3jKwolhblCS
`protect END_PROTECTED
