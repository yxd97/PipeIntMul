`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Ry9392MkUBmOiFaXrN9uRHyftpqV2yeyvdZLPho37Bm+easm46ftEkYZvQbyVeQ
7P0+wA2QeH6dmrYV7Qox6QYyR+glyTBb9/EDKEAuV6wfHtGi25HCIZvDi/InE5vB
awYUC8KmUhzdxPo+TcigWjphSvA4rYb1TdrZo9963F1N5Omj1RKlQl6Z0ygziabF
7Nql5Y1nf25AFToZ3YhQM6LGfGiYIY0gUB4h45H1J8CmOrWbMcLkItzy60bE0ppI
mAajSRBg1fhcEoaS9yfdYFKnnTSz6EW+p9dsGnpfP7MpXjPgndqAR+c9ayJOP6Cb
Jmd2dYXh2lYgbmttnT6dxxA8D+9eKQnV+sZYNc+3ilDhYROjBUL3Wikv/VCswB9H
ZmUyZxxZHeepRKu9H9zAsdWXP5np5tEilInZxXlOt0whVUQrl+0dUUnG8UrXwqZP
RYeCQ2v0S9X9p+wrMoDIqWYFjlXbHei3PUnAZZQC2pqBpxZz5gxl+RGBV1akruwZ
cev0ar/xhdbEYmAHg5q/VDKRZ56J8u4Co8JdO8Ygb8uzERz2R24CKI6LsCwyLnHu
KuFoxn32lAmO2uEbhxT1awUR4xU0YxDVhEcC4jKh1K11BPq635NMkFtCk25V+3qm
PSsbZAloa8DpnpnQEzK9j4ZV7GH1wsKXLh15oshnaIcNA1qLh0HFgLYcWt/u4sFM
sPnx7RIqVb1QIJNoCm7YaDjJx9L+QdyqpkIyk2ROtGuJ5vmimudAbR5crU+eElCV
3xggUfnRPVSmnMsb1xDn7H/S68jOkiooKfR1JRJ6VrGuKZTehwuqYreWazLs9Z0b
np0WB0FazPKhFfLaNO85qJHf8O2KqLXs7nJ13RZszxUz5gUvj8dXQC/r/Eya0C4q
`protect END_PROTECTED
