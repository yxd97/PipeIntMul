`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFJ+UDApg5eU55vTSPgzDdjoGpo11v/G+6ABViVxI9tfeqEPIi1+YQLVfFtXS6Ze
HRATRF5SdYZ/YUndriW7lfD3NbkkwoPkVKUBudmqnzixCiVrzo4kWmkEsA3/1Bse
i5pAuXEngEwpOT5bqu9WXDOqfUQGToaCMjF9aAlTn3yrkXnPacCKi6kvRrv/1ZYk
e3fr0elg4stSzOhBcnBg4zvPB+Gbjy8qE1ofj/HaKzpnIgvKA4vp30Ia+cPLKhrA
66LVG1WE/mjMRzwtSxya/I6YCqxm5GbPsRvPirG/BaN/SL6u7SlUR7HzwiibAoNK
HEpPkO4oQYx72V5xawHICeYXXXZRE7fT9yy17tbfuP5DTEZuWhNhfMAHkt88zE7P
LHQrBIHNlS80SfiZ0V21PJAdZJMvPVgAThqy6AonJyIMRRP7zGpgTX3mMR9J/SUw
ylxeVXXgCZlDKOY56VIPpUa9hwWzcAn2PiwOXkmwO9pnpTp0WDyNcEj4hP7X0ANC
`protect END_PROTECTED
