`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hjy3lyOFoB8aPfzIDXbaH2m++sQZtbDHhg+TUCcHGR2chfERDpnZSfxFq59Wvzdi
86kRlbOEnBG9TNQmX9QtgdNKoid6LYuSAuQGf5sK6KagdQ1HXm07PGNHXr62mO3I
ptx5lK1Y9A03bySKyYTwZPJyobr202VLDxd4uadtSVSd1yxa7UckCrAbmaKJIPrV
XqwjhGqICvAAIRKYc1QDokEgVxMFED42hogV9jALFwFhA9lVw44ZdMX15i0gwUbI
KuskjwWmKJU4gk9DtFctN06FvlGNgt46RRxyAAJyeCBYujeeTDcGQk3zJI0l5shu
OAxt/xTB3ksFN5FwTWiAL/OPy57VMeaKz7UDr01UIkUZf9dy8/IfdtzTEd16+Gsw
tI5er08gTAewi90JME9aZucYu52TFpWUL8uNXe2VSMD7oXG4d0dymcDcXQkiuJfJ
ygPh8MATY6xGJMV+X2EjnihoTYwxQyCjc/HID9KJl1UC+6ObiPngcXViAClOJw8A
4lyXmTX0uZAPnIKaU2vsFWV6BxqHKsE3tNubQKoMExzJpEe6L6VZ3izglpZK02+Z
YJ79jl2ShQTzDDTw1NCogqq5l6W01xp85FEPvZDwQOLJ/rcnnyVGqq4t+9Oh0TS7
NJRJi7B6FbKlrZ0UBgIzGZVQuVMz5t10M497YfX7L1rBjQTlvxTZ00QXZwW3f/Ll
SYQaXuvP60GL7Xg7Q5jKrnoHsjOIgQk4kst1KNG76VfnEz5gg9wFx0zpqUsQf7M+
2DecF5vWdDkKJUFRni1jfNxEMV1q+eCx2D3TcenucOn5/EJYlFK70edHRVCnraLS
ZiC8kzum3svK7f5m41PeAx4oSZvSrou/DRFJvZeRieo9uQEOQ/I6moUICmULEode
TmKZr6M3jIAt7dBs+YbKfB7a+oSA5YQbs0gykCjdPgS0BMT0LzPvaJf2z31aV5Pd
Fy46ACgzKoYeR8G7TTMts3zW2oVZ+N+LvyE+THTbiZ3J6WTpgyaDyJuO2Qezo5Ff
SAgZi6DS5YYrxlB9nB893Hyygueql20ZO0mJzaZpI+04cVBq42ao9EO1Fj1fVECE
RFNFmjiylrybaSfszHx/kJ6hl07XA0r+z9Nip+rM6DV8f/cxyckxFoa8kbxxCAYU
41NMV2ZgPmvR89QHp1qHB8vFq8Qdn6HZj0OywkFK7vyJdfhwIiBdOeejEjbjpJIe
4PCOAPdi39cRHBZvgVqUMeYEvJLjhlCyZ1S37+RwrNQoztmROYuUOOtXdZgv4pGo
mwZ/IJvXQef0wqT8amlTlxDks2mZo7AJE+VARYE+k2E1X/zjrPTqZM9yUwf9/6NQ
bvItKsZPpqRyPnKHpeFn8FbAhxLFuGArynoy+pmO8xKBUjB9m2LwTS1wYZdL065y
sIf/eomsEKhm6nIqsGdFN5wE85ai6a8Bz3BbwDQQwxXQKKelA/icOTiMdt4lMckt
RFWuftX1E++dnZM2vG04W1MmuPsIwozXqzAFVBR4Y7r0s5GUC2BToOfjCIfkLTON
IMFH/peGDciqgtlbTtOFwFdEUNZaeV453lRbl+pZYObPvMbsH/NHgQiniJ888uti
`protect END_PROTECTED
