`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PTqEwy0q4ktDzU9BtDLAqgGvYK8wkPidwr82awAadkBrfBElhuzuE0DkOimq3C2
8YkLaxoPuXEnP6P2uYe+0naAdxS8ylFVmpJ78GjdnGtMUBKqhTr24rBiffXUZ7gk
gMZ4ryAo2TW44hzI6nSf8gIm0ZaYFqNRKPPRMbV4up20VDl9Ar1bWCVTbx0fIaV7
Z6o2AXkWxRspCcROIR07RJntN6pH6S1LePr8RNGsTEr4sJnjxgC1zp7dBCknUoFH
JwYM2Gg2FwUQ0r2Ovwwhp3L5C2W7YlxXEXBxmlq6AcjehX2hUbpL+QK0QyZLYH1L
yo+WCDit9OL+gkx3QVqjs88gijZ3rxxRv8x0WYNu15crNDo66qPfW+daoG/RHI6E
fpExLaf5ClA+l+dXhU1hgODBRPdI8WlLx/FLuKPj5MinsA95IPpAUOZHuzMOOfoI
2RyEcyMgE+O9nYb0+3WG0nf9hvpcQRhW3b4chppIZ7m/z2m7hdOvIf8PlcUSp5/3
f1dfICxzzLyAmRhCIuBkV3Cq4wiGQxU5nG9dv7MKYctDFTe5C+lq65wboBRSzqVn
`protect END_PROTECTED
