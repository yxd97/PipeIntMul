`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VRUZeRqOjR0Luh712z93hiWQ4kqDWOc7ZS+Nw5N0ahfwOeeU6ojNV3Z6D8qot27Y
Dy6pOmyzAj1hPWt8idk/Q5cp9tAnplRhEb8hZ4/ISs0o6fhw7M1WlVxHi8zcOOjL
HviYNoRSQcxtqR2ssrOov6BRiAkBOpKafIEfu3YB/UDdlScfrgpBq9Bzsp7HIAWx
qCEP695fewjWZiOiXzVW2Xm0r8rwV/rUHrsaMBWvxdps1wXzrJ+boKdJnO2xvB90
5cXHW0/SnUik/kfZtxQJdV2loXBRuOu1vZjSR/UKg/It83mQ3DJufOPJ/IW+ewnp
rdfmlCU1EZnDR8Vq9WZarfTq1pTpPMH3jD4e53itL6Hrph2OBUgwXEHo/aot/SBk
HbMeLBTXF6Ml2Ml93oIk/p4d09vVv6WhdpHDzJnawkSSw2lHPT8OsMgbkICoL7Ph
`protect END_PROTECTED
