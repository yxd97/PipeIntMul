`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBnlOzhlSjlV5Bb/7XgB7n0J4mHasl8tpwjBLVtg0sYInw5bQlNJpZ2FL4UPlcxP
kZ3FmgiQJif/MjJn/d+HevJ90NJ8+FICiXmkldDMIkR1mrJmxfecKgRVI6C7uBa5
nv6yob4MWNy5oZnzNPQqjygaGnJ2QjDOPa1CE8rRaC8M+nfzGJjQW0WfiF303fKw
gyoP+nbctg/1NFUpFKev+Ni1cbhAAtDkJNJtE4/FmC1+x7jAO5b4uAHVuLhEMhG9
csW7lkmptL61S9eAaUVexpWF1jeSZd87bkwkixbKvnw2Z8rwi0NlPtCU3L3koqmK
oHhpyKk17N4BGogsrOO1kteNMDPTIrf9r5/GnJ/43Gmf85IT3tIehI3m/1kHgNWo
IulK88yQoK/7NjGDztxj7lQ7wyuwt/JFzO6hoDCnYwA=
`protect END_PROTECTED
