`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IRoGb/JJJdO2bfATA9Q4EhiUd2cyVqOyF/VTLsffEYh6jos7+Ae55Z3424ichsJW
2oPKIcfCTCSBv+d2bBHJcksj+SpQ1qHUGFjos5hgihA/gzxLSFaFvVNauYRcXP8U
8CgxHM8ijfpzCH3naVFUzgarPIUPmZ4JETlDRfXpPAO4lNjbo+pvKYWwBTUQ8/qQ
6PgSlpzzrixolCUjjBc1R27iMcmKVqV2hkMeB/AWcDg2XZq4yMyZ+G/RCLUKqPpC
821w0z1S0kAjkgdg9WfsZ6yIJBt4yjB9JinKE7pWAPxz2mFq1mFqzggqxuC01i1e
tQ3TiCaz8/BiiNfSd7AsobHFq4pBWd7/slpleRYyCscCS6aPRHNivRKEJjETxDSe
/XsilvprRo5H3dHL8sHBgw2R10EnSCTLFEpXyhJ4tsarcIfz+bZWLSrWlkFxZ6q/
xkH3YCJRqafRlwrDg1PEkKWXZfL8HIamk3S5MUrYr1B9u7pMIaeqhlcfayO+B5Sx
LXd4HOU2XSZKroirOBXP7JAE/TQOpx/FzmlwBs0dKXmoEGV0oKheK0+4O7oBe8VZ
`protect END_PROTECTED
