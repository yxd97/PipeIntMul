`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvihfDvpnozLLV8+KtVpzWuPxhYOLoqvSCj8BtGJ+817GnLS0yuEDTwjOLcs4Xc2
GODeY4uw4N43bSUV8hwQclzLofzGe9gvr/wYBv1/ExyueXwu1ZBwbXXdXBDoMeOa
Hn/7xy8dQ+qm1D+89UR66+q1R7cSZ4n369zNGAScP8LdEtF9X1hj3ap9nY0y+wSc
y3/kAEMwLClv++1O9tmFD2IiVEYYkP2iFEodsxUD4zZfjOsdBKz89DvplihyIn2e
e1XhAGqDY7zubTufi8drySrxYZqygTcxQ7jk4HtG6wS/W0WtWa8jxz2mmvic3o4M
+l12zuW3MRPbpo3AJ5PKQw==
`protect END_PROTECTED
