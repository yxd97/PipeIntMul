`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JjSS4ZD3xX37YsyYHwZXdfazyP6B99FG3gwhaZmF3NufzDa7tSFfRaVa5380OMhA
CktrhoGWDGrGvXb0UbeX2K1cMAwNeTjukcvQpZCDAOqn684gF+gmopEtqrgQUFGU
1Qg6NFVWnWcR9TUU2hPSXviq+ZbXUSnq/My4WbC2isvvc/VQLmdrvwH9lZAG9PIY
bG1UPOQf9GQ8v8FK4l3QwJ0Pme4Nfkx4QdPkgJjjCUReolrRJUE434MLUjkL0lQ4
zl+72eMhkcMsxzYRmYOcHw==
`protect END_PROTECTED
