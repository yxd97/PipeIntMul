`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NI69JyMYdjRElUMQFMUhKQR3sYIDp2tbz8h1BI5p2KQipCVpuwhaeTV9Lq/z42Nb
SsxcevIOYOMQEdYBjW5+YATQEtVBcErj5GB5hl9KS20CxnMU0G4lH3yUT5EwxsJJ
JKHDE0eFrGXYN0RWJfs4yroiUhJRtE5kNbxMoXUfwUnf2dqHPUg11XJpe8qMgjwh
CaUmeg+MY8psIRVlR4sGXW3WjMchqXdh/82Fj7OLf9PVaqWwYMN/XmMMDj9Ytmzw
jTyxmPUClyjr99DPT+eZ7j+acbPoBIu2p4whcGd9rPm8n8jPzWOUCi3ayPDS4yl4
4pkFvMQrxyF3HRDju3lCWzZO6Z8ZOtEmv0KEXaBUozCg4jH5Q3bKgNJKjPfFESkT
/McGBGPvbvIsstpR45pIwkqYDxDNBfT/pg5qr6M1Sg7ZBmkGcWmYUjBzv+ugjhkM
2NVpA23QWN7CiJxAKjTlwtilmOsnuR+hsBTS1aGKfKUNygOSHOrDMKqPkiCIVbT2
9ZoKU4mbtZbAahajm1L4UOHhAw9xobd4YslvCd6EJ8/DqdhBjqc9k7q6c9/kol4M
rG/yl53Xm3j6WibF4RcBAKSE42zbJwi5p/rqBp3s5NdpsBlbdSKcakQZMwhwobzg
KRayIi21AghAX8e6Wo5nbXMOkTk9StB0LHmcNGpZfpKwGPG5JFMBb2hohExKt0MV
LRfNKgd4dGNy8PflNe2jve77+pR+sPpL+chs7iDVmANY7HzA29N5gGmc2DlmyKHX
sC/E2T8J5u/Z+RFD6d44TvMaOElLmh0ng/ZMAiLCUJW1CcYAhyzPHzn0PtCzIeq8
k/JQOoSNnpoXdkmj5zGPEjJK4pLNHMPuE7BKn7gb0ghE5ppHMoYQSsIDjVaK4TEI
D4ioOCXFZ9mPe0AmOsHUw+ij002XPUah7Z5r8x0yanuRrZMbz6u6pYxhh9U0pYLZ
L0j+3B0/2fzQCWkghTfYAObDbnWq26I2r8BqbxLxK3c=
`protect END_PROTECTED
