`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EF/1IW2F5LZs5ZdN02NX2g6a3Bzj4Z60c84SebDVpeubke0TLMhliRpaqr7R/cVj
I2Mlr0xKh1qgPhhIXGkn8+WF/IeMbtufS0w0ia85GXo+A7StgSzLFfKDfVsasAaO
NW+cAmY8Br/LSyxlqcpd0O4e/JvaKnyyjvfgKK/cFRXwHbnYZqS4Y6TNobCRJaDo
vLdUamqyjBy6B5Vt4ImWChjMTxwvu95VGOAR54bUJzUUp0+gC5BNphUTHJFdK8it
ExvCEZIux5p0euZSD2JjLv53oDpL0NO5uyNdLOzGPIKiaegwdBHj6E7O9J0KALaJ
BZggDditV7Us0R/Gvh3Bo5v1f3Yq+xX7ATFPnItj6KjeEDcWULELcedmrDJu/1Sq
rWvEzc2h+csVutOGmJj8bOo7jw8Ybhh7nxjKzQwTC59tB6pCo/Lez80vpjo8iZRW
RYjiCySqgUB9dBuyAQjtqmp0XiUjZmhyfhZG7cZ2TyHGhLONHrPZFCdBEfV0BBJs
aSI2xqqTycIL5f0WdYSn/MZGgKdFmIJ/QrSzROicgM/aweZr66RZ1M+SIyH90APl
3PBp52tjsrDBkrrCAomBIMlKX0f8L28YdH3sAdOi4AIXrDeis7eDqQPx6TunGdK5
UH9gfhAmXqVSRTEbLGV3vVriMTnkbahRzFgSKZhOeeZPSIbxBNcF6gXSjhFf+tMQ
1viry47l3OBzuJ3ZB1ouRfR/5lkfR6z89EJylPbg1Erld1scALXPWFUX11ZB+hM/
sfA8yiPzTF9A99YYi7wc4ZPSeiEBtGRY4F/EKdSWoCieODXjo+xHplMp1d5btbfg
i1F8DQsBqp/RAR5zCAXUd2UuQJb/EymxfvGmdCnIxdNokexWeyGwY5+9splaakyZ
qrr7kmAw6mOOrFo9jM5nynVTxXUXmsrQ6JdnBX1OLSb2mJKjJvKKt99g0Zf1PjYA
waEkOZOM5QeWtT7As7a4DLNcXAun0JDedMnIRzZFL2gyw6Flmhf4+VJ29EDhh7AI
RGjLDmEIRri/y/LxbII+l0HR4eLELQfuRs0hUZLuqJndFxcl3taP89U5YOdn9x8q
g4bRLybNz9brohxF1Anq+7urODp45IfA4brucLqUm5Nffb+reRmyxWJ/9s15IXoq
/6tLUY5SG5DY0cjQo3o51J4ZS2FfcPRHaqNnuEEybzjAGfKx5xRKtO8+IAUhOGTg
wp+ouX/u8mkMub6dYut0h9oJaLdU87fN4/Mi9ajMvDHqCCAhDc8njszoVWLTBANd
MFPZNJADOUVNne2AOanDGk1z3IGUrIY8K2e+ykzSsf1QEcLT9SdUASV/hfDuDT+G
ccJ+9iibfxajdK+I1zmrpnJmLIMjgaoG3dOThVu8pW6B1VMuT+3YqRTH+wGQ85R5
vY12xGmr1mBvz8gPjjGcRcdJ1QVjKSlHPZ4ncuaW0s1sDzNsi2PstN2xO/QiCrDK
9r+JtTqQW6KZoyTsNPK9OcqTSPPlY5IUfcWvDLODi3Ewc5jZCbQ2GzmDK7lqHgf0
39wkNQTcwd0eChJv7dea90HRmqI/UYCGTv3MG3nTRJj2AxgW0eXaCwvJvo0l99b2
dXdiOIv0yNZN9Wfsdubve/+CHkMnVDRuJdPVHhZ5gmB8n3QnngMbgahdC9rsc516
S8X2kJJjMz6ltwDpwTh9bfGchNbgH8suaN+xHokdUXwjapQ34+0mCO4eL30cV2Qc
kcEeKOviQKvO22bXxRi6Jvzz9yV39FJj1+buN/tW4l8pbGbYfoLzoRcBuH6TISVp
E7ECvAx5tTPuKSEm8nVL4y9Wbj4Oj5DyqIVcU8z/LtIMWsGd9rJ+59bEvHJNhGoE
fHHmhxTTlGNDm1rxqG8Pb+piyHDP1sTEWDLmJPG1ldp7BxclxPtL4PObcqM3ukBc
pX9q+RWotss5prnrcS6IrbZfOLVtGeSZnlmw5+5EYLvJHRPpJBpBuU2rVwJczAzk
`protect END_PROTECTED
