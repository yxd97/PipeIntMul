`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eCKdX866c9AW36k4HONI6CfTpxG+QcWlq4ddI1UFgj1CNT7bNw8hK/WVcY/7EEmU
Lae3IqX0zTCfj0000O21KcY4GcpSkFoHqNWhcGGXgeoFJ9jFPCr28RqUMxzphhtf
Qqg8bomQ8uFOB+oZXTGo6ZFSayrrkSGisCF71l5kyZVgSDA/aLGgt26iyKrCEv2h
b5iEQJM52UottrOC8qK30vFb/p/iwN7eoeEWnXeZRZ06QoUUPEuGvWj0RlRI128g
4IKz1tO/dmNm2vsNYxRGraoqvJWRsI6fBOSXHJWOVkKW9t2Tc/s3P6pIG6VpYr/S
IiGUeCYUmLZL2oNSkzzIsnfr8kAGqpkCAq3MXYEUOXQJnLzCMYBjkpu3nim1yw1H
hZdW+BFxpPqDmBBK8PP3ir3D6IOKJ2SZr/rPXNoY4BwpClTrqjPmChZh2LjV4w2i
gfxWhoNQFolAvz6yEGNOcNEMcieZRfMxtJ3143fb9vzdaeeJswmsKbmP5yD6NvKR
rgxlmxU7qMTnFAIWfZCMStBP5j0vM5Xd3ETpkl7FFMTigbyqG7cK1Ta78oaryWgz
7XqhuBy3Tjgw4ronoroSm4BERHcb8YYO3qfGG35PrynGwOQqj6PcBWbcuwNNf1yE
40CSHaZFkPXfN7KO4BR7mWr3Pwb3DLzO6VC+t1YIuww=
`protect END_PROTECTED
