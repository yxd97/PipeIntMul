`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
InPNsFA9mr1M+BbP/qkfaFBxdVXAYqEepHTxRvh/fzNTv+r3ga8qs6E9MatuRghU
Hd2VqbqemhAUATwm9u8HwwWu8C+jqXMX5SCRYPtaCTtJuw4QcMtwS15CgWsWwcxR
e3rzE25EKvBUIhHEeDVIkdUAl0cngQGJowkb0gzXiaG2B9A1PU2PMtWwINIezZHy
yzlxGcGeFE/HVyozxmDxDgLI/FuTyKOj+NqsL/aWqB85xoDETrDsXUP9lFpw8EY9
56B4oadxqLQyFkeoG7mb8PQOK9pftzlrgI0ArH/SmvjlrcEhglZqhhngCFEbHFnc
`protect END_PROTECTED
