`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QAlW0d35KPEFFlo4KfJbs//iazpDNDJBeNfHs/XkpFZn9arD06piflj+URmISZI+
VqaYhnF/bdj6Rs/UA2hRpxDzNH09n1Zz79V9HxlzFq/n5BvzeTUSS6LG6ipy8Avm
uKPzpZFxjsMRR8eXQM2uKXB08Wz/7i3mQZfeScLIL+ZW1Oxqccmf5WUPMeoKG17e
Dkm6RFd1lv9+i+aE7CAtVoyVfJeliSEjpzpzuTXDMa2P3Ha+IQLOQi7nGsYgldR+
vVpow6YYJcMfgNMA7w6mRg==
`protect END_PROTECTED
