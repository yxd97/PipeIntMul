`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K3Rl0KyXkAYhMsR3SzzBFRSjhT2lzhMc7ZxoHKREwkPWNBAZ0L1WB03TQuE5g94h
TouHHAxHkMxbMfGILenfia5pq1BO16o5oTv3CxPwp0dHAYFTa114TB0x8nTezAqo
cE8FVWtoEqM8ks2xVNyiD7aL7vUnVIDXMqF+ZvVHEf0WCQ+UNK5e8HHBOGW95By4
8PzF5EBcSHvUJA76sj0rYoL/dWe7eVoCGn3yypQa0bOSoCDTOAdwAVeqLWvF++Qw
yuNsrNNPBLmFbVqMNKNCZsDtLGG2rSEyddhVzPMuFD+gYQeXPvh1E3TJfz7AQT93
ESvFrZk7h2q0GwoDF3Th3Q==
`protect END_PROTECTED
