`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xd+6bEDTuyJxEXsKgyRgYFjw7pRxOTHoLYgbPhHMvel0atITnLdUF+rXrWPyrNJM
+VDQfF4igMBPN7hsggltqHLVwHtYqj2xLcaQ75jndguaehHMWYVxqumfyjAVmTw9
+P43i4WmmlDqHZlDzI/nmLYUaArefbADXLicDB/rwRyqitEACZmWPwfnc8Rzu1Bb
pRwvHG6pEiHii+zDFakHwl0ufh030OXTXNT32hjUqQ6a0k/DdoYxjkqm/pjXUS77
FLMyx71mV3QvPubPTGVwEA7mnSUAlnf2euxzEMstcj0YHTFnRY/Ut7aTqiVwnU8F
gMTmcz5oDSTSchX/InfVP1G+ZZqcjwW9ftBTlkNA/EJzMK4S1D0c+0aEpIksG+UX
LCxtkoQKGCePFRNQoQlGhj8Wn06rhbzdE/ZA6QD0nR47pCTGQ1aerFBOLl3hC7Cl
lWbwPY29802RteWEhEMSHZ3YHP+0LJWQ+s+RaOgmCxCRR7jJV+6GtKRTiwIx7T7e
QgqMbJSG6jhAvTFmbWVK/cH3apd6HXHkVDI0F6pbePceeZ3N0CsG36ogwlcldHwX
VXS030Y1IIyQN0s1+5wYnJr+1zQnDPeKUI8r6ShiMaC7uJePIzB0GuNR90HjHjX0
dxyfWi+GGCcW8fYxnbQJ3rdL3fGFPA5jecLrRgpTHXslxKQ4+4/0HyCzvob5G04t
ONoUE/CgwrWnNAaAOYaz2GWSIFlSvdxiDIiqw4B6VLOqwE7Vz+iMlwsXrNgCNdck
qaOO9iHoA5k/edeN3PuZ/FYJHdBiZp//OEO6Kb9bQmsxkiJpNcrZcrJxjurzy8Gc
70wBGDUtwqjK6JYrFRcCPEuvp+Y/IH2YMDj+6EbyUp+9+awH7X16BfElwAAuAp8C
wahpFj9+l3KAMrIPOxDj2BLQZpuVnncQKjapmJ3tAx0=
`protect END_PROTECTED
