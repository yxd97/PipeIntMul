`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z7x2x/2gvg2JER3QjfI73bvfl9Yf1oQIGyyBQIi5gXoXwNEoGY1NMompm8m540bl
0KzLSF6bwchKShPnCwY7oldFfH5xxIomqaKQYLKrR2cMUyNKIeg5bwiuk87ILlu+
e7nz6gJMDfhGCzBHasKQZZcikB/nshsYwU986sZ/VHil+Pyi1by9zHcvMhOH1Jpu
EAJ/e0teS5gZlnOF5SzhjEHScwBTAvn4B5uKQHTteTeuONrH35MEUjm96vEE9n3M
tlJAlNFShBTgMUtgrHXqVREhK/sUH5ri2Tc1K+Vismq9dQiVfsdrKMvIyDZOyrTq
FsgbDsSBtEOH6H3v6Le4fw==
`protect END_PROTECTED
