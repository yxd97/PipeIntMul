`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Krx+v4KV426T/Uue9Dd1N+WGUaOOFHxZ07527eTupkVpc1Hxrl/c5MCoq9ltiJSB
XVZaEoP/5oEw+kHTimyZJ8NrkYeIgaLKhJ3D8hX51iC0TaptqlrqcxN4rqV3KP9u
CazeRwQ8JMRY7HqPgaigQuzzFVVhMI7EqGdFGnQ/baXy23IBEsrRTBMfikJR1IUT
+7SCyT7q+Z/iDZpmhk91SAM4d8leT2c4g+ADx6PGSzIAllBHhBf139++ZsENFwz9
7WsExjKcsaEBp3YYkfBkxGG8R9LTPoe6+uw9hhaNFm8v5/WrtxpmhIAYSM171uRt
as599v3jPUPiqZI/tAzpkqE4zeKQpasjRAiZg/R/oHU5fdXdXDS40WD5s0OOK9qF
OL5u+rfXHaXGpkIHWbzZEEoqnSuIh1nDRD7498F3xsWkmv8ibVWC4D7ZMCbasCqZ
1rs/EGuN89he278SBqAAbNTQi2gwppbx9+1pR+Gez4Bpi62llvqGI7Qoe14dwdAb
`protect END_PROTECTED
