`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NX8cHYQ2xDDQ/Tdo6LoW5qZylJkJTffyj7Jv39HTyMfo99P/uJZhcg6VBbA36PNu
wYz4dq6KgFpmbNLSIx27Tb6K28EqpIEnwUdPPvvi5MLJXzFg8O0+B/CT12LfEHsP
gl2rr7eWncW5F0MGoEaQ3DZOf67HaErrLmu9i4XXacIBW4zBH8popZ/Oq4lIEWyr
LOAMQOMP7qwDo041x3FY0XhLGMvdGM2NE7ZsIIPSQyI+3gwegRMhUIiy7ufgspGl
IzrEBrGPJl0GvjGeQGQS6Z+qZkCujUvb209vHQODyYP4EteAxlNG2qgYHM1fma1J
VgkHqW7IysibvaHm1ZUwNDzX1V7YunHWawafsnK1JfW2gd8/KC6RIb4Cj5Iv2Uyx
Z18K9WToHbnMd5PlRcS8S75dZ2WnQkkfexRbz6Gp96LttMgLun9q1vTIljjFxb2w
eLwTKD7NeVv1d5mKB/a+eQjtIv0KSuFljvjP/rEAsBd1nf54UzCC+UaXfead0KzO
9vB0dcwtZuDBZbpKcncRTE9Kr/W80IZeCMV04PMxaZjWZJ+llN8YISoVwoWAUUYc
X/P9/Uk4GKnlBGZHTric+Q==
`protect END_PROTECTED
