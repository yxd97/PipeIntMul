`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s559nz0Jmr348x0Yc9IqsYIfqDUYzuyPtYCsK3k8TY7oVFAfmIQ86W+gcws4mQjv
z5nUIjdi2Tq22HmK/VpEF9mUpCg2FfW0Si0fRyX74vw4yzgrRHE65ez7oKT9wyaB
TLA7O8KOuMvVkTrHZHhL9VrKcNvIc8Ml1h3nmu/AZ3cpheuXrms5Jph9gFfPTIlY
8jF+PXH8N8vIwNIBYACJjCAc7Me7MyNU58SnjxAmrAXkwOATiE783fTC0R9n9hCg
lsnWXO5SCyDmeHoGoQRnug==
`protect END_PROTECTED
