`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ZdaSYKQ0L2O7O9Ae6sxwW35jWRSaan1jvtUn4EBM7EPpVd05fuErNaI5gHRcVcK
Rb2cM3VgZVRcMe6CK6lCdiIf+KfN9Pisl8qvZ76FDKaSBVp5q44N6HlozPY+PlZE
ORg1pyYH/EyO0AEmtQrh3cBOmwU8HDmY0JWmq1msf+DqyYD24n2NfinFPdZaGmUp
KVT5HCdeXWTpCraa3cPP5EcLhdBy6noT5aKZnoYyYYoqPDflG7ljTsTVRJQ6I8Gk
XsjEi+iaNOWjpXHy8jMGNpaleQTVSb+BrlShdSpeqMytpq9y2buLpCU0S0BRgOmk
akZ+a46dxZW+mTRJvIF/4zH1miMJU67xcTtN4q5ScT+mHEoYO0zaGWhgsTeVFTXf
fMMbcTTLHRInlcFh5RPHFFAeW3YUth6U3wZZ167beT4=
`protect END_PROTECTED
