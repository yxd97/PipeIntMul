`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXvOBaKuWYDLB4MzmhVLpVoGmagmb+uorlP3XthEhuBPFx3Q1XHkrmZC2F/0Cw/3
qCEQTaKSkqZ5fb2NMGHpzitPCDQbWcaZ9SIQrsAnH4xXE3Ez0Hxdvee56V42KOrs
5Iraxyn5CL2Ws8RdmdonaJviWQG1e4plO2KcqgNwykiCsamf5Jwg1CNlFxP4TloT
rHTzbrPB8yPBBD71ilZrfeS8BmgOlL1hXZcIk1Qm/pB9IrhObvC74fZdKpEgsiPo
8dGamBLOuU1e9tJ+cD4ANVYch83GSVupM9GYoDqKvk++VwopNcIT2Mq1bQ2x04Ap
M57e3dwXyNm+ysnrKWhc+I4kTEI3wGfLI8hgs3npfibBFu8F0Qi8VhONDMISljeo
DQ1sA92hDh9DEjdfrCPNHqRGiWRyOcdJHWhkFF5i+gL+Mx9ZCn/cNNz9DCj/d6FH
UVBnxqaxVlL4mUXHGb2DUTD5+TSqBHj86EvKHJA9uHErH4ZoVE5fpgBvgYBMDso4
Iwt37BeHPM7iosdR8mrjUGxnPnibX17MsirwanfORsNXwxLUjddVwJqOWmJA1s6m
f7xR+XajzX+9sIy/7FjYgVj0Wz23qeVSrFJF6seSDDk=
`protect END_PROTECTED
