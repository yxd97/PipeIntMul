`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/+BG4A7Sho1BFJRbFAlEHewUJPohh365wkjMsmiCF8Geq/45EO7sfuxtMA/RMMI
O3gkExcFCkCUW8hmsrq+zdSEXOje7EmmcfQS0UxXPBb0bfxydrwoWK9UgEWkjx9d
s5yosf0lrcwW4OHxuOHQYBi5UdSt959Ixp3PBuCw4CFKtiwSfq+xT+2ZXHZHL7Ky
TJ45icgqljVSz3ARsCPxTerbOBEskk9DqcyP7Dv1T1e5tnAoxsttEDwqmwwtbbcj
CJT0uSZZYe+7rw6+NF41YH1QIdM1+T6wdjEYh103w/0AxJxVUE7vzGDB4JIY5/HY
1oNth4GVgbbIZKOK3USt5+TgHO/Yk96XWfsh1mNQLhgagmT0nzymT+oc8XO1PpF5
ipkhxn6ikt66sK7N2s+CDHQ+sd0Om1Yg72TvWxzDx7w=
`protect END_PROTECTED
