`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o4YaKKfjHYx64qYxX5pUk8lYSiKFbFiHkB7mVpkdOl13akCrayB01P87NgRAGV1N
6Lq6it1cYPCEtLMjqFS8WekLSvbHPowtY1WgW4eNfdiHjkNgl5cXv36HetpmHzLS
OUIK/FdLHmON8PXPn6i2bx4vSr7k5yQGadx/QqShNcGneWMRuPWp4bLMg7Yq5pNx
3SAhymHjD7EcHWyV5JpvCRYz1KV4R8NWCy16BaX1zxioJkxHSakIf1+MAGG+77ON
iJDf3K4xNEIkJ3dRvhPIKiLF06+BSFTQfIWe/ABTbhvrJDM42++Oz+QoE0K9TTqH
Z+ItsIqyS4lJgL9tIqqwUS54vJ8zdo+CAjr6kW7Cfd0I00GCEHU1PG9CASzO+p0t
cmu2x11oNkQ19QSOePXOjUgbUhfsljCvuq7dol5memm6eDKDLbGEAL/yRQzNbHoS
`protect END_PROTECTED
