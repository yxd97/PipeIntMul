`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LGJEtXAv/P+Q9Eh20ONuVf8eupiDJuf/N8dyZzGe00mLZsVQtUkPDB//MmZXp3Qy
4qw2Osh14rAVAu/hN395NMzW7PF40OxbwB2cCGKDuGrMuUUDCzvkqN0h5jo5TPQ7
HTM+JID22Um7ef2lmgJ4+Ulp1gie8IPhlCprgCJ7XtJl2N/g1Yzz3VT5srPCz6jJ
mUPdwgAxUiKlre+71QfxHTtQabW9j/4pw2m1uLrUm9iQ4zLi06k1RnIIPgKpKlNO
FskDkMEXPvVAJv7JsbXi113BjajLvbINa7RPPSjpbWXBBIiv7DPDZ6dXJmMHe1Yb
fgprQ8KBj+lagJnUPETpMQ==
`protect END_PROTECTED
