`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D2CvEb0PNUSI77PJ5OFh/M8k4UcMV1RzU68xkthsbjBxUxeobmpK92rjPRUhf0yS
gATqDlD1nOpTGjX93JOqft6HvtKAhmakiICl7+sEM24Zrv8DKJfoyMu8OiY3Az14
ufoF1LEOZ9mP5Q5HNY2OnF8cHYb25TN2/xZ2EOhsYTzs0+/FPqH04fgN6hSdO2H0
fOriPKEW3I+NrehfYN2OuMwjksGiA/ge9LMAoaw74/KftIuj2xHRQAsBUg89BgoB
RuYvIP7mtZf620ymk2H5KPbuqU+2lVUL+TCnajBBeC7EX/1fkmNkQ2gHqs921zZh
KpEpvBhN/V5L8rA5+kFTB4wE6HHu/4iE9TCVChtLutFzuVEW+OeNQ7fB6+CyfwLC
JhIxrYI8ZKl/5ZffH/rPq8E51VkrGSAlfHMPk3UzYP1Muc/o0AJBO9SPg6y5LocT
F3pPW0TbqpMDLAM5su/UlA==
`protect END_PROTECTED
