`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Pd0diNnfWaIvjpUNqHJ5IQImMm4urHVXoVDoUaFGjtKNVRpZgbPONFf0BcDkJtB
4nq5TNkVcEkrxujg8NPL7UaUChONJ+/sEzAwFvf8pJUe9HjnqLKvhiNnR7QXgmAo
BpZwguVVKsR75oaY+dmWjwr3JIxF+rjRJoHm3cY4qbuVtkWysedfPG+KA6WpVlQs
2rUWI5ii0waSRODBwN6pSKRQjOs3vKb+ZpqpSN8vXMN9yyVuzN08TrPtLkeDN+80
pVqQLf8iqht+vFEUoOLhBU4X66n/5+0gGZxVG2Hoc6CdLSfUs6GpLM7GSyLow0aO
kPPBx3BOYP4drETNwViMjPBCKo8QIfNZYMnrffUiRWNwplz1cTn3xo6rwhC/+xPt
swCfSlGZywCGjZ6o2wccv2rejXMmxag41MF5qr9/sbI37yC4ia0JaFZ+BiOL6pvB
QAtPTFYogtFLhE5F5HeTueRJRh2/KVbHBVqSvRxlEbmVdvffR6rz9wM08RPZiBVx
tMfRn8CQdxMdCuQnybFngp6ArkCeR/oFTcrHtBcIlJJGDn5AGIuorIiQ39C/Vgvw
`protect END_PROTECTED
