`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LdD5+jAlDU721BFLQFpvtmt913hQYxvS95kJxQ8vlMl3NcuzeIUvB47zcKUfLSbW
IS0vaPCLcyXMayYcO+nQ4UKM8G7p2WvWm62zf9G3oM8kZncw7N6/JGFqoxsyByFB
Eb8VL8EasZq+hwLvbiVSTmHhidncdmavUYGHYmG9qNZsY+MQQCuBVcTjoiopU6Dv
b/RMdVN7WbZB2t/Mzjb9O6fpT7bpJM1wQdCx5Ld6RFGeaR/Od2EUFRcA75sggt57
CY3TD96pp7Y0n8tBul1FdMBo1gQo2TFJI0jrBk1SM4EnQtuB7gOzcgbFqhRnavLH
`protect END_PROTECTED
