`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LNFbmjmn0VFuidlYJLthYllRXVkR2fVt2RWo01wnLVls31Vv4aHL35rniuv8bXya
TUbsNxCWxesas1hzCztOi2mtaymZhrWl1v+Ik5NJ4l2QnNFInJ8is8l3URgjtfds
62PwiTyvkBh7+JpHSw+2ycTX1jumrTmPolJMkAAkQYRoFrTcJ/P23ZmIKXlza+oT
IsbjUdz4W+W+8yNhbZ7PmYp1dzKouLo4+BVDei3XhvDSG1G2HHnw+514gDcPgAkR
lbWzc0zDDskMl9tS7aSBuPJ6fYOE7K3a+T0L2+LXQ2290Cxl+UAUDyP8wneNAvsa
HIdh9r2tjgqbyPOwBJ9dOrTHx+SvNib0g3lYyZrEB/iDWdt9lMognCkQeEeOmxKf
b9KjHxZmmG0P/0y4Tl2hbzltJZEZU2Eksrk7WQJfzbHKhpm2RVOMPUD2Q500T70S
vidyX8vQHcNF/CA1tzy0V+CtM9GlkakLIVvrwUcdf2UMcMBLUXRZZrj5CUowfcrI
LiiOiIIyW0MXPz5g1PTJUWLHRGo+L+bk7nvFZUrv628=
`protect END_PROTECTED
