`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV9TyYRcXDEMWLg0itE8T3wD6UX7t+FcvTjbp6k/hIygnsQDRjb8QyjQaLHGOdOs
/fkQ2Z8Lm9W5+MauAsbI6ZM6cyD2EV1rocpc+1fBt42BvylM0SR4d86C9rx+7TyZ
LwPevIu2lM/hXhUwXejtWsMsxZ+dPM7jGcoZYVVKM07F5YZ03v0IAoDqxplyRHBb
6JoB5EUx1ged+hNL7FDnozedX0A1I9NDRJQyiBzYKLKOitAgX2BFa7/zJFAM8Aw8
izp5mMGVeHoSRGVYnEyUP/Ed4zFSoE1A9uMQ10VlEs140DOFcZOg0rBsJSvcQ6sK
6B/CegIOsZrppCBC9NZVkHdr6Jj8Rr+L7Cqe/d/+9kdTMapEef06vYkW+gEFhddS
ZmTMdyRBf9PGD4ZdXO9y+KVpxR26cUaW2oc1jegMBxMW3V2VpOvyJVPGqZb3eLNk
CGh3Yfxj8iXOpaoT1TF6i0TgxpAeBsOP1+hfzhDjoUnhPGOMJPQqmvuwKc4+snBt
c7xZ2WtSyAisc0H4kcqSmxiKsVrW7X5EvbUP+SHtlZwdcXab+U6vWOJSibpV1dzi
3OKr1aKB6ZuhU1TBtSyvMLvIxA2ysCz44XSSGG93cJLndz+UEobLkvknwOJPqucQ
0nnOGYGCRan/Gykx2WYkKmE28SmqBUwt17vdxYkjhuaJ2FGwe0YMU0pLpdQcqVWx
MswDDQdNWnYnSU4jr96peTvLc/etG4BDbz33ozMWYWpw+pG5iNKUSw2gVLUdzyPE
SsJNJFNa0COvN01cN7pJFbC2rfnceJHLgbPcOfInD1Qw3dLDO7lPwVQ0P5deP/3V
SDRU4Dak4y9lvpsTariv16zbuAufyhHxT4f2qECjVFwgIq6xPY/jgugjNd+auaNE
TZvykBX344LS4IcDUOVWEKXQ3ULb3+xbFwD6A0epr7mviEGTEFiDPuTvtbsw6AWN
Bjg0bAtX7YFGxS/7Tkqt/LlbWicv3sjVma/5LTx0IfdOEmN6HMW4j77MkeP0NqVf
`protect END_PROTECTED
