`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0O8TZ20AqfGOiHlM67XW2iDdw10X3zLufhZMfPilRgXoA1x6Hg9FS3hcMp/1QT0p
6KPQkrYvY9yWVZwflF95W0Xznu2puYY5yGbscfD+z2FSgX8qGcpczJBEwcQTIyBS
qFwhgiUY8dgK9YI42xCJvQ0Sdq5PNPTEbwguc7Nd1v4lWJoDKrGnEpjpue8Ic8TG
GH8RzSOEPX9ZoEL/iGADjuw9suKCmzRdTb5usOd9AaOPy17nkOmdEmQzgrs6mFjm
R7iSxjvn40arBAJuQWwGqrWYSJPoD0T7SQyxkcfm8DgveZi7Mm+SiADcIrQxMflo
O0oWu6L2am8N48vfR6DJ6W7RNE/php0QsAVB1bW1VLLFWWvgyKw0KcsEuFlZAOJg
EmmX4tgmZedOxBmSYXTE4Dgsn+/Q6Lk0VG55UYjziV3lYEvtU909pJ89pJARUN4T
pNWFTNIARlH4/bvpRmV5Zu2HTeXE7pJ1Eh6GYd0tHlUaDTYEWqjkOwZSNAfsPe32
R+NCxn0NxX1JxO8V3Qr5bm2Q70GfCKnRlCMbj6X/Tf4YeVjVLbWeB4A5vCPIqAqz
5T+17LbAtBnIxyZsoCiqr2+wgTxKeyOLmNc0rm3iR7qMMGEbpTO7TONfOPH0zdtu
/tuquutu301TVIotIACN0/2o8XoM8nSJxAYDu9fF0Wsz+4iOHfSkiQd4qy7+r39v
pGtoA1Z+bCNSl9vuwgeM4QzXVo4nsTlVsP716pvzkg6mm0aCNSkTKQSAwWOuMtX5
86uCueATCe+wGaQH9/90iMfYhBXqBqcKaRTmNGOj3wX6guXP0iw3sXxM7iGBK2Hr
L/AcltKLwzhkuMP71mIxyC+t99nSkLHMgMkLRxDuxbqWaYOS8Yr7F+Gi5eZka77U
ApocUAEgACidEmZwgE+wANpi5X1LNBFXyxkqJbYf/C8MUjwlerk+SuwQD060p4Fy
vfK9bXxPrx+2CumDoaX/9DsyM26AyPGeg6KQ7iSsQJV03B392EgTFzOelwAJHoeI
rq5PUq9vdW1sJwTx7PtMxz56MDoUrMbo2tIjGPCcWJUgWP/FW0HN978Jryb16zv+
dQU1bKYxMo2VTNkF7kSgzg==
`protect END_PROTECTED
