`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AuVHwr8PS1lJPQV8a2Xe1lGp/mA/YAov5ey97EpkieSPpXTMqRXvemvzGiKr6Blv
H40K5ODW9Pt9x1AfFWJrY3yg/ONvjWWyldY6/l/OYVylBjWrDrB1Y48l9ORfrKka
UOENq+u8H4helcRkv0ut74dG5dUvt67RK7J8bn4oksYg2cFih+7bll1rVB7vkGZk
sT0YKjx9RfU1i1yGpKSF8+zu8BoqFH1WgkgH+gsmxPs1W7kmy8dT9+CKToLJpw+G
09kwvBkBD/Qf/7LgfzjyFp2nYrnl6Mh8E9iRlOD2ZUid7hXrdIQmfY87Qlmu8fzf
AcV2rZQ9DzJoLeRHw5dgZUS0Ec955zE3bASQhBruu84SrZIRbCeU3n05lBfqfdiq
uQsChHbge0LzGqVIq17Zxw==
`protect END_PROTECTED
