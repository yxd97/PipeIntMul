`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kNFL8lJPPxEkbGsO1Fq+Yew23/tM/4NwWbdgnEpsZFJQajUfmVwGSoV0ne334nEh
5KBJrYSWCm0ttiBWz7HBe2WGcnJHdjJyJdVXzP29SH7ZeP9ac6VadtELKzgJbpQi
KxiI0guhHa3hGBoHAapOZP7Oe6BNpNKhiUE9NHa5goWNyRmlR3/XmZLUjTzs/OPK
akZHb/hO1031yrCy34CKOTLZX2YwKjx1aSlsArIoOX0bYLG49urIqoonMCpISc7J
Pd0US+C6Os2Q3bnkkKTZyeUgoqAs5uWp4c3m1X60TMuf2C2ojQtbdy6aiBEDVYaP
C/GcBRieiuQftdyWq3EkOA==
`protect END_PROTECTED
