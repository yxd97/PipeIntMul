`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YfdwK2X3bjXD5rAzK7A2vARR0P8UngQ0V4ynqC92w+lW9GTeoWxMLND5SURMA7Sf
S5W2K0DcOxlNbak/iVe6xMhDcX84pQt8Mmqcm2xH34mjUiE2ZT6sT71hsUfbtvCB
RmlKZ4Uuc8UI16ZrOECgYQBpEWdgchQ5h/zX38OIAqPG8fgkT2K0G6Jc7di9eYnG
BPryDehZciLYJi4sJL04p4IDvSK4W3O3FJJbkWz/6VZpfCJLRpT7yA/Ppzf5tVo2
j607arqtaWE3FqdapGvEIXq3ywL8SkyZD25TebI+TEn4AkMx9CF+buJZKvE2a5T7
he+FPN/pDFAGkJY3h18tameC4aApnwIiATlG0yVdXkjfkIZzfqculY052d5oXD7v
Fc2AIY2dSA4B4EuBvrLqxg1VkjRzUk71MF25b6NqS9UEIB3jWvvoiGGzRg3liFyK
q0YFt3LdIP0c7GsgFEgo/rUArRJxi/A7TJONeJOzevUznV7lwk0mZMJs31Op99qS
zUwdoPPz5mQHWB2yUsIvve/+rN8A8mJqm7Qu/cQ57pqOpjaxpESiU4XlYr3fl8//
54WjmV3Uhco/oABmIvfr1ejf1dc9p62B59YcGNZJFFuEQCXvUfyHziAsqKDCAVhg
PkBvZzWgUvriBfIMiSCUuRBDkTHddI4uzUTlpkr9qBXV9rI3s4cd5F1q2jxlYw5G
xUE0Urqsih4yBxfGALt9ct7IugMlMrVzAzGIH3aU4i3X1oGt5IM9HQIjfifSBgDE
dC8gc/zC5O1CUX+iIuNugzeh4Efx33QAoF9p8WAFQ6adpMbIK8yOpmrDshiz9jRy
nrEKDcqK2Fn0GZFV5MVnFA==
`protect END_PROTECTED
