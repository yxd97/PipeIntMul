`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQfLZ4dNYAumH9BiFzGHZqncymjU6dnXEcBoq4gHTF+vZyEJRPVhUbuZkXWwBPNX
Bmic7QT1SQ90OATvRsSWlPctdXHpxIsf8HpwHWIXcAREyFxqVVUjUO6OmddWFry5
+vj/wbNlt5oL7R1/6N/SYQUIWFHaaHBgh3O/2fFPtA/fIIvsaNQlw/jueMl+RCt1
slb2BmNlgjsFxfbBaJSRThkkgbp9gy/eqbIArbrQlMIfhjpVHiXjb75HyyMwJabA
MV8pjVzS1wXZ29ve8drEom+VIjHxzuHNQ8+HVJgxe4nv+OFPH8oJkNAzT3OoRqjf
F7r7R3eeMyglqBscN/bkVw==
`protect END_PROTECTED
