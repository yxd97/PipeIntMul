`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9u1eLYx93sCTwqbKmxoSZa6oVc1DVj0KklSCo0bHr1P/MfIxJDGX8Ful4m1H5l9F
1xDY4PmHkAZ8meR3oUFkApvwFRINzc3Bwg+5ctl5QssUMnkILCxg6tIIcAh2SQ8g
j2tPzpvUJuQCBUbg2LVHkch/V+vdP/SucBID8dmodqIe6QwonaBa+wDhM29Ms15e
fmBE4PsbJaCk6OZR+dzQS1fg+PTLjyeekBPfKDn4MPL/+o3J4p6C1OeT6tO/6SAT
ySBI3+pxhwLjPDGHkwKWUcHJHsZ4xw+hz145umOOTBEGNVlBs8nXzf+fKvPD3xBV
icH1oYMKcJxH94DkMC3X6kaXm76FSj+sQpEFTqEX1Es=
`protect END_PROTECTED
