`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSDeAlLjNHq4joLIBbHOMSjdaZ35gAhHzfztg/UPTRuQdroMQAnNAvjaY6csiFDH
Okae/0hrTrFEu4/T5u6XFVqq5wcodlp41BtK07yaIhhR6r+J0O6ta9Im/1brFMcn
aL4T+wTfVzigMXC9OQ+6Tq0XkdVpSFOwVQiyZqFJC+8mugva0SOCZX+V7pJgd2pb
u5U6bDttFsh3bbsVEu9duAU0GwyMHRFW4V5Yi9q62Bj3eV40dKC2WruZEr6Nfz4s
hFfMBwwmbX3MOejZzlej2QB/9BuwS+BtNKvGO96YmgFuq0Py5Vhr+ZH2UBdE2+6M
ZR7UI9rwYaBr144NEmXSsxhF40pn4HERRFr+SnV6RmkUHNBtPpNZL3LHeu22jbWQ
/5Uw1bQ8zT2UGD6gq3/AJdhB63mx4DNzlVTEZaT0JsNdkSeWH+nY3lan+s6WjixI
KNjJ4a9z0zO+bE1l4yZr3Wnl24f6lFjUl6migmBOWR7YcJHL5jsI2+cyvHdRGjPS
YUyk2O0qma+PkKwcHsUbmLTRii24Aqa8afg8EK1Cb0qudUcAQigE6WIn8XeXE2qI
xtEsh1AnUBJMTJdF5WtzLyXi8fXYAxkrBdyorissPmpTDDXPKInshL1aW4Bs2J53
n6okFVoA3Zsj6ApNNF/DH6ePiUzCiCJll/iKcJm3ai0CA/ep07MzLReNvjAKhsHg
CLp30qmk9qOpuK9rH884AgxweDZcEMKiQNj0zZQ+li6tMBeFPfixEG8/1RtKWyeK
0AQDF47hUZvG8gj2OkhOIpEWhrLUQmhtEAmcb0ckLkE8PDUjCQCqQqfGMkf6anws
yjmjriskDgWLq5K1rT6yI6bgoSgwlCw91SejdIJsNwitQXnHPQmhiubLGJqLdlVP
1TL+JrkdXLisVcqP4PskauFnupZZcoXwccBxqzgDUkkezROFRnBg/zE+/E61MB97
jNygqXoSDHkXC2fyygrbDYyGk106FH69YxK0/1rotTXtDCF2gzPJXAgKL1e4jgdi
xg6CUb/Hx5MXModuTA/gXmUx9TlEfWA6gBTZPNzsnmeGOjXhqNsFsCbknH8Oq4cy
BtYwLx4lSVwpGe5evr0W9MqGnFD5wS/Yx7Pe5O0S0ePtMNEaLaK6uX4xZo5h7JR8
J8Sws5hAaD4ZWGGCOwOF4YNabzBe6zNmdqDS7basaXqw9pXWwd4fjqvgHc1w11wP
e51jL22Qv2LxohibIhpbq1n9aI1FTwc0UBfxh/ILIV5p9GO8NSI6PN03KZ+7MeQl
06JSAcm7voB0b4QsjYKxX9CkKCbp80WPcePO50gxtNkVhdTiQtCb+5bhpoouEcqr
QfYQ44hR6kI1ro9cc0Oqqq0aUwwRuDQRnreSiZJkwVtEcQHWXYrM/WSa4jR0Ba2f
FjUDrW4UTwr1AfEwVp5QpDz0cDYKk887sJ5o5bX/fUXn5Vh04gGQ2yFVY0by3Cfa
bburWV86W9rnm7yfF1LhxbkeHaeINHyQQhq+2ZOwLVTwyBymF/E/f5Xdc7zdEDhC
GJtc80P4qwIoB6op370iPYDDx0jNwTRvYDJLR/sHHsQogLRmCwu7m6W+yRlu9XQC
u0VfrLLPr+61Qbww9XJdr7CSKQl4TaZvt+qxJZbAuA0hLB2NgwBfeno7ukuucIzg
vaFD4BD0S9+HNLAEbzzPeRRkNyxv/El1UnACm5H+skdd9Y4Kgkhmemqbb9+OUOho
bmdCoBLVIKlW3To0ekX3lIaMF1tyMwO1KelASo53AZCcE6nO3SByO0l5GemTloZe
aay98wnupV6X4lYNi/mbOQa853x2cI9vNnL7X0ZsNoxDzSH4Bduq8x8Sg7MVnC+D
IF9QDN4JtBZTLq2gaxNjWm+3weUESNuhMADacGTsw9Gq/mWIqn8Bk1eFSC9F4t41
LZ1J53S/FRldFxe5NfIvTqNumpA/7+zSLCoK6Yb4opJxn8ohLRtJ3kNPhPYFAifr
qgnXy72jxQHHcle2+kIWPyJggLR6eDk2sfaRsVCgIqOZvP+Zz6L7Mov6j0YoHNlq
72qBMScekAeAEA8LNIvCs30fv3KffXNYRNvDip5/w7IPaOzIApKB34niUQQEE9OS
LHtAEwG1ka9Epy84kx68/gEKtU+8OvS44xS45BZbTzlUyU8JPMNw5yEE2C7pvZQ7
aQH91r+Ql3BWhWUiW90nD47bRbB1yh1Mllb6rdMUhs6hNBEhNOed6VKGUuawhEU4
JEf5O1e/QXL0SOiF6L0YsCUcaHbDuorI7dnW1QUZqiMqmrcf1yagZiBDcUOoLBr8
XcfcAqL+lOP34VdEWpQzX6b6E5Q5rZgeeqvzvQp1QnPjU0qRRF+uboIL/uV8UKiA
EWWxMfKj2TTk9suLozDmZ4RawdqzraecIQtMTAJ3m4Iy7zNO1uI0RYmJ4ysemVnH
/hq2Fb4xf2KOy4tceYjcqpVJUYDJs6hYHCThLTsALVoARsTm1VvoctVGR6xRs6WP
qcii/N9TADCGweDlnkEwznmke9x6qgsxZ44oWb5Yx314CUSsgLTCu/eHxv3rc4aG
XMfRnNbdbCb5GiAF3udraM1sVPMDJEABZOdw0xinhH8zyUoNYOL3hARQNfHeDZxW
0VpsFRlhOve9LAm7eZSpisujqwLKj3qzlSVSeRpqCbJNWyQMjGyncB5z9vwPdaHv
9FW/FP0rYsuiKAGu5wJZkM98vzh3ZbAa3czECgS82zNr9e6xAY4S+2qWM/lrP6Wh
2o4pUmoIlvPXm8ECIELQU7PrLmskmN+pSvQ1DzS+WuNzSnOXhWusxngTWGoqmFXY
EF5GG7Pk0x0k5cwc18TeedN8lCNfXvfhKZ+h6M4gmVKMa71gisPdWmEFe9l9Qk9c
0Bl/VH9VlKw13YPR/qtk/PN3SzqX5qHE0AvT5k/7UvQRFL9RmutXEiG/XFrX0gnj
ldHIFRj9eNpPOaL174iSj9RJNPLffmEM+726ia4iNdw4QeGnr4O2u7RP7hAQm0ys
hgeYnf1w52Hn43JZ1b2Y3oHmSqVIwQhCzRyXrC785GaWB8C3kA5LI/t4p6hsXj28
J0nwBCMzukjgf63Gsasub77sSOCCUXY0H7KLKOF/OQo=
`protect END_PROTECTED
