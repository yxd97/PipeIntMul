`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbBDycv9TGFsSf2fDi9t2VAAXq3GOHZsbDlpwZHgwhyvUWE1s1MU4kI4C4evx+QS
shZfKFE/+IGPYdrErtHU8ak9963w0yZ2q/SXGxmU5P0VjTkTfUdA3qrbuC9konid
qYfNlPPLv4cWW44blHidOdw/8URR9mhF7chvkxBEeVAI8rc4ZVdppsnat7HxAjnW
uqPkLctmcmdqadWzjXf4AGwt1oN5L4wvRPRLWxaHXCWmzl+StLCo7SjXTawMRXap
j1hnbfkdTx4+vEq9IPrj73OcEw7NaUtWprCAzrLwyFx4V3DDL/30tz5Bu9Zj8uKp
AWvQZWI4mTu4zsVwa4/w8hSt5pbGloceds8tfqgjs6P2YAjqwd5u/mT3iDCzO1YK
`protect END_PROTECTED
