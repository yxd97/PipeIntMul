`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZY2869skeQv8NZIrx+tYzn2a6Nip6OJwy32bhbftHaK3sXKcnKgeDGExeVDk/kL+
lGRgw4sYwr6lSVDlrQ33URNHuZb8fxgn4O5mlwZVdYoy3Hg4vdfljkonf1srRNAg
8b9CB5I5eynW0M2QyIBUWWaoY7gFahTTNBrROdD7mN1+xtN6wsVj5tFjviVR3Wcf
F6AUr6T7HzTSQu60okBimhohfycwUyV7OaYVAIdhLpwx0fJV3uzyr2uVTqhxefpw
MLVqjFHR+TSk6TGC6xUFF3mHRSd34IGaGM/fzIo2SOE8D/b0FOX6hcJI8VfF/vBF
H4mYdEL7Vh7R54jGRg6pm7u1Qzn8NQtC/bqi8ALhswxEmWDiImxyCIbWwM6UPDLi
qjno46qrpHlOR+fbOgX4PAyvnpce/4QRdNXP8lljEzM=
`protect END_PROTECTED
