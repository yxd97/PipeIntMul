`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C7zTjRXZwXKOepJtrHNtGnrIfJlWaKrddXhspFUCQwZPRLknfxMMBrtcz1fVwnC8
WAy2SqTMZF3Ww+ySbaj5Jhi4B56SA+30SJ782jW3t3O3QlHK1ADjmLvcRkJ2o7SU
47IrhK7U8J+smXNrx5SSs0yRTC2z7ixIj1LpIfwXznpkcYbYY94UCaT00leeMjhC
ii2u8qWZexUPLD42e41oKW4H570eWbwuxoz4r76A9nq6/hLLsInwRLVQw25wR5Cz
85zcekk1QHIw3uo1+tfMu62Q3yACJo9nViYlfxQovJCeiL33DiwAEqtB6RJN9VK6
OybQ16NFk7secc8tFEIccQKZXjYlLr/rSpx3X2r3f1xS49xOV5dgi6bJQLPFBG3Y
Z+UqKSeEYzLqCaXoFuy7f6vUyJHIIYT+L/lWF4RoQ27pBuJEWS57sKS38WxPLwQn
b2iBPvHV4koncuxF8Tf/FB7tVr8QJkIwB0DSJgeYsbFdURr+TGQuCjkUq5ZnyJDF
QQM0rwET81RTtoVOGyb8h5flye2iYY1UG1W5ZQ9rI0ZCYaVvP/IUtaWnazf64vXF
plnbrkt5u/B70/q0QPwZkqS33fMz319B6uqJH3wr5gM=
`protect END_PROTECTED
