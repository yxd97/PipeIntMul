`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xIjPq+pFXPvEW0XjJRAG1SRe6LcdeDy5K7ytCBYSAxrlNLNKErSoYyx7rIlW82IX
Gjo9wlhpKRxdgh5pjnsS/yy6BFXS581imnh6tlH8itF9R6x2VkkXlRiGwknfXG/o
MDOOxKZXdleUtgO/xzlRFcHCRLIEuFHyCQE9g1+FO0PeV2202D8LIEzsuvVn/CUo
NH9ilWFf0ZFVzHvoufvp1O/lkdc6CjqaD6EGODV/dWaE4AVUIKTQMnzZuCxn5n/e
/9l6p2ccV2KhPDjPFikPmQ==
`protect END_PROTECTED
