`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
spaqxGUT1J0QkFCgc7yEVSYSJ+FCoSgIzxaFYwGfwaVuBDI9vbrg5EyJwsiVN5C4
sUQ1zE9oId37X1vLm75C39XbsshwrJzDCpoJx8E27MJiVnXMVdm84reI8NCWd+5H
f23yUfR/NJ+ht+Ybi7p+rjzHxdBX1LsYNWHmN/63AxEUO7vgPIERV5YyCd2xeWMT
L4L8+E01ZWKCJH7QRNpHZQunDRQnlMr2kr3TDbGn2JNfggzupfBdxEMZjlygwgEW
gxgSoPFBbxanMsLPJotJsZyEdOsd7CAfhL0oIJaMGaBMUer5XXWoAlWuAHiVJrBX
yIGFbDDJ/Gx1wBCXhlr2p+Qt5IRreMk5Ylc2lqcHN/nz1ADptG2r+pXdJANZvMA0
pIobrQDn7cyyXUWxEJzF4YCX1U3OPFGTqFA2dwpZ4NdzUuLvRsI/HQxtTRZCtDmt
Q96AUkPZ+PdNmzuD3Kyurjx1yC2KUJ87xHld2hbnZilVTD4DrTkIROXvNmoVIuN6
UZfDGOlPvNz9GtndsLXJ5rxpfLIokNo9KqeXUp11pn8=
`protect END_PROTECTED
