`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3mKiBF8iLb1PvdDs0iB/9vsQcjDyMu7PE3f3x4SpM6iSHyAM6EqCLr0qeJhikWka
AqlPqYD7cKJWurGFmnNmiPUuhHYTjNBB1b3BNCZA+4ww/h65KRzK5Zr9AnBobIhc
MweZ2V1G6YfiILKymDfGIhCJUCPo4ua74deW8jvJIW4r+3izxJiQzsQx+LzEHmct
khlLkrUzVvue1VHRWGCd6TIcgciXxZ8s+4KS17D0Dkmq1h4VzDqgIMbJ9Z+wR33W
cdvycFqBs9Tz+5zLFSiInPhnB+2ArW2fSPtHD1Ux6jIxNrU9P00StnSLvXjy7+27
PjX7r1YzkjYiRSPqTkTrTbds206gBmBJPOP8XhNLj507w3Gk1ifY0+AY160DJQTE
nODYs33auz90QcxRXaCzSAeTzslZXb41JFOmhLMo2YNF9ppr98Mr0icfcI4zdPIX
u5kYmk/wSLqwFx7dXzF4ogdwO7DSTvdGauY21HpYKgzONofNupcfOl8FM1eeUOWM
V4g7pjInLvOdlqmZ9s1c6MkTTg451ciWXhM6/d/nzaOuXSjd1KlUjwEAp5m0Myy1
QQqSiCjDLsiaIa/M8+LSPGSE1KpoxLlrgZXPcniSGfI=
`protect END_PROTECTED
