`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BekU7UtSaT1FuzbI6ClnoPodMnh8Lk+Qc1hBiR+V+iCYK7jWSHUYyyn74ToroGbo
YA0oqHJf+nAs2pGzlfmnJ5G8po7Uztzhf4z3yW6vo1EZIKvc5+R4rTuPa1ySYIbZ
CfZawbgautFXIJQdM7VLSbr+DI1iQ71vFCLFCHBrC0zkjvp2n2KJmdkav36DO9zG
7KjvSoEPbxxKALk1xZb0/U5+EHO14VHYy4GUeKusdrxja5exQ2KYkD1cUq9rEBCT
L9J/pVZrUulw9TV2thwv8uDqrrwQVwh6MP8IVfxqCS2EyPd1hfI29TynFxgKoyG/
rLtJH+RE3ga/dI7l+xHn11j3+wkiEJ0hPXbUowOtqBgP1FsJYWQzqco3MftBXSfL
NlaOmB1IWGzDe5yNGJeUJcHe8T+rLLzGkZY8inu6fMISqVMZ44fsm5odqoUHZz50
`protect END_PROTECTED
