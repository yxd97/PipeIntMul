library verilog;
use verilog.vl_types.all;
entity FIFO_GENERATOR_V3_3_XST is
    generic(
        C_COMMON_CLOCK  : integer := 0;
        C_COUNT_TYPE    : integer := 0;
        C_DATA_COUNT_WIDTH: integer := 2;
        C_DEFAULT_VALUE : string  := "";
        C_DIN_WIDTH     : integer := 8;
        C_DOUT_RST_VAL  : string  := "";
        C_DOUT_WIDTH    : integer := 8;
        C_ENABLE_RLOCS  : integer := 0;
        C_FAMILY        : string  := "virtex2";
        C_HAS_ALMOST_EMPTY: integer := 0;
        C_HAS_ALMOST_FULL: integer := 0;
        C_HAS_BACKUP    : integer := 0;
        C_HAS_DATA_COUNT: integer := 0;
        C_HAS_MEMINIT_FILE: integer := 0;
        C_HAS_OVERFLOW  : integer := 0;
        C_HAS_RD_DATA_COUNT: integer := 0;
        C_HAS_RD_RST    : integer := 0;
        C_HAS_RST       : integer := 0;
        C_HAS_SRST      : integer := 0;
        C_HAS_UNDERFLOW : integer := 0;
        C_HAS_VALID     : integer := 0;
        C_HAS_WR_ACK    : integer := 0;
        C_HAS_WR_DATA_COUNT: integer := 0;
        C_HAS_WR_RST    : integer := 0;
        C_IMPLEMENTATION_TYPE: integer := 0;
        C_INIT_WR_PNTR_VAL: integer := 0;
        C_MEMORY_TYPE   : integer := 1;
        C_MIF_FILE_NAME : string  := "";
        C_OPTIMIZATION_MODE: integer := 0;
        C_OVERFLOW_LOW  : integer := 0;
        C_PRELOAD_LATENCY: integer := 1;
        C_PRELOAD_REGS  : integer := 0;
        C_PRIM_FIFO_TYPE: integer := 512;
        C_PROG_EMPTY_THRESH_ASSERT_VAL: integer := 0;
        C_PROG_EMPTY_THRESH_NEGATE_VAL: integer := 0;
        C_PROG_EMPTY_TYPE: integer := 0;
        C_PROG_FULL_THRESH_ASSERT_VAL: integer := 0;
        C_PROG_FULL_THRESH_NEGATE_VAL: integer := 0;
        C_PROG_FULL_TYPE: integer := 0;
        C_RD_DATA_COUNT_WIDTH: integer := 2;
        C_RD_DEPTH      : integer := 256;
        C_RD_FREQ       : integer := 1;
        C_RD_PNTR_WIDTH : integer := 8;
        C_UNDERFLOW_LOW : integer := 0;
        C_USE_FIFO16_FLAGS: integer := 0;
        C_VALID_LOW     : integer := 0;
        C_WR_ACK_LOW    : integer := 0;
        C_WR_DATA_COUNT_WIDTH: integer := 2;
        C_WR_DEPTH      : integer := 256;
        C_WR_FREQ       : integer := 1;
        C_WR_PNTR_WIDTH : integer := 8;
        C_WR_RESPONSE_LATENCY: integer := 1;
        C_USE_ECC       : integer := 0
    );
    port(
        BACKUP          : in     vl_logic;
        BACKUP_MARKER   : in     vl_logic;
        CLK             : in     vl_logic;
        DIN             : in     vl_logic_vector;
        PROG_EMPTY_THRESH: in     vl_logic_vector;
        PROG_EMPTY_THRESH_ASSERT: in     vl_logic_vector;
        PROG_EMPTY_THRESH_NEGATE: in     vl_logic_vector;
        PROG_FULL_THRESH: in     vl_logic_vector;
        PROG_FULL_THRESH_ASSERT: in     vl_logic_vector;
        PROG_FULL_THRESH_NEGATE: in     vl_logic_vector;
        RD_CLK          : in     vl_logic;
        RD_EN           : in     vl_logic;
        RD_RST          : in     vl_logic;
        RST             : in     vl_logic;
        SRST            : in     vl_logic;
        WR_CLK          : in     vl_logic;
        WR_EN           : in     vl_logic;
        WR_RST          : in     vl_logic;
        ALMOST_EMPTY    : out    vl_logic;
        ALMOST_FULL     : out    vl_logic;
        DATA_COUNT      : out    vl_logic_vector;
        DOUT            : out    vl_logic_vector;
        EMPTY           : out    vl_logic;
        FULL            : out    vl_logic;
        OVERFLOW        : out    vl_logic;
        PROG_EMPTY      : out    vl_logic;
        PROG_FULL       : out    vl_logic;
        RD_DATA_COUNT   : out    vl_logic_vector;
        UNDERFLOW       : out    vl_logic;
        VALID           : out    vl_logic;
        WR_ACK          : out    vl_logic;
        WR_DATA_COUNT   : out    vl_logic_vector;
        SBITERR         : out    vl_logic;
        DBITERR         : out    vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of C_COMMON_CLOCK : constant is 1;
    attribute mti_svvh_generic_type of C_COUNT_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_DATA_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_DEFAULT_VALUE : constant is 1;
    attribute mti_svvh_generic_type of C_DIN_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_DOUT_RST_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_DOUT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_ENABLE_RLOCS : constant is 1;
    attribute mti_svvh_generic_type of C_FAMILY : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ALMOST_EMPTY : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_ALMOST_FULL : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_BACKUP : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_DATA_COUNT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_MEMINIT_FILE : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_OVERFLOW : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RD_DATA_COUNT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RD_RST : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_RST : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_SRST : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_UNDERFLOW : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_VALID : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_WR_ACK : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_WR_DATA_COUNT : constant is 1;
    attribute mti_svvh_generic_type of C_HAS_WR_RST : constant is 1;
    attribute mti_svvh_generic_type of C_IMPLEMENTATION_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_INIT_WR_PNTR_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_MEMORY_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_MIF_FILE_NAME : constant is 1;
    attribute mti_svvh_generic_type of C_OPTIMIZATION_MODE : constant is 1;
    attribute mti_svvh_generic_type of C_OVERFLOW_LOW : constant is 1;
    attribute mti_svvh_generic_type of C_PRELOAD_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of C_PRELOAD_REGS : constant is 1;
    attribute mti_svvh_generic_type of C_PRIM_FIFO_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_PROG_EMPTY_THRESH_ASSERT_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_PROG_EMPTY_THRESH_NEGATE_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_PROG_EMPTY_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_PROG_FULL_THRESH_ASSERT_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_PROG_FULL_THRESH_NEGATE_VAL : constant is 1;
    attribute mti_svvh_generic_type of C_PROG_FULL_TYPE : constant is 1;
    attribute mti_svvh_generic_type of C_RD_DATA_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_RD_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of C_RD_FREQ : constant is 1;
    attribute mti_svvh_generic_type of C_RD_PNTR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_UNDERFLOW_LOW : constant is 1;
    attribute mti_svvh_generic_type of C_USE_FIFO16_FLAGS : constant is 1;
    attribute mti_svvh_generic_type of C_VALID_LOW : constant is 1;
    attribute mti_svvh_generic_type of C_WR_ACK_LOW : constant is 1;
    attribute mti_svvh_generic_type of C_WR_DATA_COUNT_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_WR_DEPTH : constant is 1;
    attribute mti_svvh_generic_type of C_WR_FREQ : constant is 1;
    attribute mti_svvh_generic_type of C_WR_PNTR_WIDTH : constant is 1;
    attribute mti_svvh_generic_type of C_WR_RESPONSE_LATENCY : constant is 1;
    attribute mti_svvh_generic_type of C_USE_ECC : constant is 1;
end FIFO_GENERATOR_V3_3_XST;
