`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WsEB2eb857m54QHTg1XsVvg0D71LrGXRegq5DdgSvjmg2sgOQluEgBD3tcA+AprA
P6iOjKuIPBVHX5lDxg5F4XgWzT/AWv4tQpstl4TljLnkTWTEdT9/OOXTSiIZEV2P
DhjgA8WUqivMP1BdcTwDvLEQtBPXbUOLPBM61MHL94r5gVUNLjEJzUtaT2XbasM3
1xEGMJMQLE+6rUlHtgX5MlZP7s0DY4Bk9hicvq3VRnhJUf8f6WR+uxItdHuW+rTs
vsV/I04nVd7BIjoKfB75yrrLxgbFQgEzj7PeH3MFCbAt6b3YLtinmo/OgCy0QP3F
nGA9XInDixki8d6T8AbhivUogsk+cRpMWegBb+ASWt7AQMa1VMTFX63p9YRGM5u9
GQAaN+HDdJqMESCdGywcaowFWA3iYNbqa2EVzDoSr/Pwm9gzfFcGt8U6AdjWor7M
ZfxbBGO1u3U64desx2i6wme7FoNiobQMEMtq9eruqZ1a3LtFioE+8TJSyKkCvVXM
XSqCiU9EThwMq4LW5Q42hn2lULaAUDPaWY3uzqdzk0DWSBM9Fvyb5GtBENxCujSy
Zd9ANFaq11WE/JR6E0loHk7dHDz0ldM+6D8jJ2TyYZHNuIpI1TA0hHUL04pal++C
5jVIY1HThPp3KP6AnHXIS6A84Dpwwv8YCV5MEo/H//VdbdjcuV+ehFQHJo+p4x9i
O7jeXcfYbbC7lUg33pUlOg==
`protect END_PROTECTED
