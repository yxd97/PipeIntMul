`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KLJG1XHj9eadJWTF6wHZeNigAPAh1Ul2gTCyGOJu1sBVS/lInSG3HNEQMnKGcAX9
o3avtKKgjktTT8hny0Y2QABbkreXD9vKqpxozY/cQu7ozW5oFIaWF5fZi/ySCjao
+EvexUCby4EGCLqKPmQZTF2d1y1yBhbax38PvEitSUdD66I3/0CgLU9Qj9LikgY1
XCwn56nILBIbbwwemh5rK+dnUKy4wXLFFkXT+T7S7cLPgdaFiCuHoub6Y+0NdkGV
brJwkPf9CVeJ7iWKQP04PQ==
`protect END_PROTECTED
