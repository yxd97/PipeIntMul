`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVk+YblYBBjAPPbi6CcwOyplHXk+cVcDGkR3TE5pXo/zGjtWanar4FeWKRSxezvZ
wpNLXwaatv7hXXStTF+1Bkk2OP5ArMXeJny9gWF5QD/Kgz5JpLsHdSY4K+zeIwms
PKxd8sopPnqkJHozXjbkBA0HLgIY1U1VTxGOslJwzrxQIlP3507Y0/WAHg9TFJ0p
zYGrkU6rhcebrgoOFBtjSss4MIZ1qNv7hFABOViG64Z8rv9MeIMlWuHFsTlDkWPw
f66ExxDmXCFdzQxhSnQyxcdxUsFuvL2iRV6NTyGCfBg=
`protect END_PROTECTED
