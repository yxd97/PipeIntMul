`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oW8O8ZLk/cEgwxBw7pGBQsmC4cGjWJefyyULhqREiIuqbSpch3I8oxo5/uGswFE+
aKrY4hQYpC/xUNzuiRjnXl1aSg9oErTlW2J3QS8dDi6+XbCZKIAlgIjXWSTzorRA
HTltAX+LHSWYH6P9shr1E+yjOKGrZMlXfj3RJQIMY7pSnS+G/5wufJUyB0xgvn3f
f/RbXyWImcswGsOvz6z6XnCdWfv/vNxcd389hkslY1vClT4Gaey3ecN2M2Y/U3m5
V57OPWxtfUpOPQxoo+D0WjrnkUAzzP8WQ8fNh/xT4d/t46Ewlng6PHD5JzT3AGId
LeA12Dv85kztO2lsc+07xGCnc3YcjyYqhXa0mEpLt5hTEKAeS7gaOM2CAH5izdp2
aVCEhikrmNEuLJ8VRl50SEVlcQ4WAFtjyg9tYx23DjbM1/7WdqZbKw2PFZsG2pdt
w56Do7TMEGLxaCPXjW5KMVkrEXAeP48+ImDXKIjt5hgUMNcGprE3TJNE1BznTOip
0dR0hzfo74AuzQEvdxvV5W3BuZojd6tTAziN5l+9FVi9AsgmNMZFazINcC9LnQnL
cXTTEz+BZ1V47yUUdlTiJZ9GC9BdFlIiGwq6R1V0954=
`protect END_PROTECTED
