`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZCJduxEma4Horone9s/z2Feynn0OqnO8y7i2Eoxyok9SKdJzxk5xEsb4n48+xiNF
ZCC2E3QLt/hnQ/GtCl7MKit+rjhyJeb2z43Y/0mAm0Imeha7muiCU2VLyP3MWfTh
7oT/ap7LQWi+wtuLNygBlIQ46PPwJlCtKbCsPuvpFAzA9vgwhbAGyxx0fXc1/IC7
GaS8mwe4526/R0ej5sDin4+3EtHwnYas5aOMOI9MABmFzOjYHZyr4TwOz7kKnQBJ
1Iut2s0+NT03yKz4gtrChnlaI8oVnrvRs6vKDsc3A9N2gqWU00Sx96AOf15nGf23
XW6RY4JBcgTXSQBI3L0aRZ/si61m+DTCoFiPeMOGfGHqGpSb/lSo66prgefd+/Di
Q86LBiDM11zrIX7n2vT3DTX7vUWDyxohcTzWPTF//o+Q9QHW/HPhi7p4hI/UR4eK
u58MuC6dX06ckg86qoJ1dz1hvwWag/sKKHxapLAv94uPM+M8EpsTWw09G9C5ONUM
BSzcL1CZqECSczuKk3tdnkJdimfW3la4SGlSAMpTZUbtdqoYDXcxKvYI6g3Y16ZR
pRAbRNcLqWYnhZJ2tHVjE0tEF5z+Klt7My5SfTA4oqtM3XyuKrjmguk+RRoHI0ok
sMIZXYQGXKaMm3onm8qb82xYsSP0sREcCUDU9ma0vX0+exfWPtYX5M4rPl52WSod
sGtC5Tsjksdhgx+lESdYa7dHCvMeY3W55xrhLA59tUV6/cA+F0ub2OEeMb5/2voN
l4eeHs3s9Lm8gzFc6qbU7zQrWlC2govwknMVHC6ZsDuhMvHWjF7raYk99ZVqgMkG
UehLiJ2LpnLCdw3z+oxIBr3ESPPu7LtnblvcFwhVzFMXEAK5sTTPTnEdghvZ0k2D
1fzYPI1IHD6HCEWIvtqQ0bm7peblSUEFn95va88B/T75QOnuK+45oYCc3gE8/2De
0q0eVAyDpfw+GcZ2VyKlYohsDxRejxVkk+/A/9xI78NzpOqZxU9GxWYruqDshP/i
PIuyl9wr/rOO24dgAoOnu6mHrdrPbAHIkISP0VDLneTFj8iBloLp5pUsQgyDzxMs
Y0dTJQrOuGjay9J+53fAGy+U5zrWb2tyUvmg3ATHkTG2GKntvXiq1qXdC1TYCcGQ
e5+hkqtG9yDjPGG3aZmQpk9e7RDrz5wprvot+gW2HLCCfF9WzeYwTMQ1s/7sojQR
O3hAQ/ArK/pm+gpIXHMZZoFkyO7xKXRKLLbQxPcMCCg5aTd8VK7VWoNJxitOEY2s
O0pedpzHqrnqsv4Ui9LPMnEwMhkeeV0U6hoar99LqCdoqTJa2f8yi3KMF8eGZZD6
7pfqZqSUn7SNkIYOP6YbJ0qAFAVjA6DE+Cb8FjpS/rIYAk2vEc8S8U2GlJmjs6Pl
+Rg/DdqcTvkVlWGjF/Xpb2bMKWsnVXktgKD4eW6ypW/1JJuaonsDMSdsK+hJhMgS
xosPMS8eI8LMQmSdjSO/6j6kacDtSHHCEqaQQSDIxjnpEQ+ebOfVBZ5Z+tQtk/9T
7In2Hynj8LbDFOt2eCgR1ML8kTICur2/Y4g5n1CtdQN7J84PhyMg65kP4OKHhQrd
FRRN2IvxvN8BrdaRQNvEVaGQI8WlJXbMTiXfbHGcHCdxnnddQRWnJgWMeSoJJej5
UqDGNkRzUbd40AdeR1wzYFX5lvDOJhBEoC3n02qq1XrkDbgg9yv8Tt0EaMtkPtJT
iJSEImnT4mx+DP37U390Y9tuGOav3rf71EouMphXk4MtstIc2Sdkkr0neodws7C9
ftErWAJValLm6R01U2GogIXC+wM1Dxq03p5KRa/DsZ0p9E3CVCX+jW1eFgG1nvZd
dL0xutFTKm05vzEn/LZJ9pGDLBhxX45NnoBSC9y9vUZEa+pjBRBt1yWvR8Ioyph+
pywRMX8Zq26bwbfl+Ar2XaDIRGrA2OFf0HBfnjtKce0VG6djH02ae4uJDw3AAFC1
OegjwnbxT06tbnAAOONRvMjqRutUvPIcD63SrOwAj7nII00D8enpmFXFRecd/CKb
vzj8s7NuR9lmOj08qMZIc5ytrLTf8x+pxCuLXSYOvJYSTXGHDlDaBRiJJgxX3DpQ
J8+ldQEOanHqk1yJBIByc0vQwseAZb+qdKLBxiyXeDTDa7i72QbHJBXJKOhCCmpl
Jt+Dwu0ud+4UZmNpTUQy0C6l3yBBmo6Lt4HILpnQPmwGfZ6m8Uj9LtJVvxaUBTMk
pGm477HUieM4EqMU3cC5IcQN5lAqmNmRYrFOkw+R7iSPI2ske81nxD3NxOrjqTto
Vh7Omynj1tm2X860npjf2aiiy/t6RNLeAr2qFLxNmuJd2UH3/PdHFVLqgMxR0LYY
ktp/TW1VOlymoCORgjbeFukV7RkiksGLR3ChU5T6W4SBUH/jxGLKbRJinIyMa1i0
9KiH+xDYhE1urgxPwRJmL2DqQLfsTJIJj99ynLpcaemVYPSYGp9tWGMoViPoxqrR
39/BGkUzHvajbIP6bZq/lGQtPLuv/64Xcg7Vy+fL8ZyXN/+OQgVsc9MqHFYOFeYm
LiYz9o8gBRScdpAAI6AuNmG8xqOKvhauM+kcoKuo/2JVCEl9rRd+jnn0jvUyWoGg
FBKXwGMPBN2FXLrVRG1cfz1iLeRgrbJgxAUeQ4B5hIDjU2bWiEkTqY8qkLDsZK4o
pi7EfUfhQixHsfN8ZSDtUpQ6NwIIzFhdLpNHQLvkzeOLiUaSqt1JzxKm+0n0XNaJ
IMb7p6KTXc8POfzCHCTqpiyyBl5/5FMpPHeVjK8AYE0SXrHtsJd7cM6ADgAnXiQn
woaNzFZg3JPXR6i68/b1/a+MUHzMAwKXKUcVGRWLtebbaTQ4ex6lRz0eG9Mq2DNm
Uh1QR3MOWa/RQwQsEUQS6DGyDY2fskQXDe2ba+g7lDxcwA3IrGfzYmF7/hKS3j1e
oRrB1AnbtqLncWXH+xPxaxP+PkBzqmOzlwywibzLgmnLEpAkfqc6dxdgZCoaSegy
rBjuPWyfHqC+zz0DN9Wg+DfJMixEDuBO0CAa/FhNQWUNACpc4/H97k5grt1wNkUz
Rs0tqQDfGGzRUmkE8NsKAnqDGkvLlUsIMUA1CXbvm86WlQFpahkaOtFxNpjXWVn5
rdq9v5B7CXFakB01wNlKxgby5RtIrKmZ4DrOHDZJSm45yu/RuyxjLVScyFAbF7T7
jU9bN5PfuQG/cg6Hzb5VFSdeiVvDlBzlYTPFdr8C5uHIy0wj7N2DxgC7gkFdUP08
A4h67zc9kTH41XqJG1RhBxyqQupLywHNnqkX2TAi2TW3K26Du4tSmkm7wmKafxOp
hIRwIMJ5vkG6Dk4G/UQrA34VhI2IUiPW+Hl7rhWmb9gOcA54DbJjqG7h0KUvVxA4
KCTxAiNDxGbww4uTu3PQ0talBDW3z4MXejxofo2dDi/0NlKIHWFRJNXp9wTwkswU
8GuqBQz43MgpzbTRDpKnheLYCHS1o7nbAXZmIqY4ctZEH8f2rtYhir3qZWQMzcOM
8uHDpLnVU3g7EU0sgS92B0kP6oczq8Rq/HTzwAaYyet+aX/Bi8uo94NP7ChSEx8m
OPlAzqrGpm+hwvvAaX1fMBIfGGkZDDGCMcI+q8Ko8pU=
`protect END_PROTECTED
