`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yxagm1Eb2WOD0ojVr28w1arq0WN1TkB8CtoShBbeYTUchd8CcK/17hfZL3afp1q+
WEyXgKT+nE2BBPAP4G85wsqS/qLMiSMYYjXPZQfijmsLSSs1/e7yJQ+v2Z9cOhPt
MBXgvRPtmV03fzL/prU7MkmJvcgqcloStdwwiPK29cmz3ofHnbb6nGpaVxoHB2+q
r3/yobxdOxNdalXGd+bjBNA+B4LU7wIGtntWP0CIQfDProc8cdqXPc8ES+OvQqLI
9jJavIfl4Gn69S5pyAankQKMDia/VRSpOY90xMP7HP0BBZv6ZxC3f5Y/wLwvCAlG
X/PqBznDprACttZuflF3Zqm3iKUfY7Cu6CmVvefa9PrI5se/JL7oBOPGcQGtLKbw
EF4UrfQMh/s4bJ9nSY82dIxeqk0/eR4l2K0apWZ6Bi6d30HdV58XZsZFtz9SlBJ9
SJyFNhK7Svh7ONpokm+ER1s0n02neU2kxrHJ4pDCNRRafMrBYgfL0cMGSeNu5Lt/
Qi+mpaEEl+072d3H7/gC452XdRnQo7t1q9ey5otuRgSlFoSZoV8UNuM0Ih65Rzwp
ZFFHsVMQzd6CK6TtKZnI1Cb/rTpRuaYS5DkDWXWLFoFQt4C+/QS+W04Qu/wLSKyA
G2VP6/Gk8B4A7hziW13kTQqMWI92CrsbiW5/UcR6Zg0f1WFOvPw6zRMyZnZNfi2L
xmTvUMH8AT0PVnBx39ZYUAhmqrpj4ys0owfpCJvfXA2k7dzedlOkEKoioY2HyArE
sQW3tcsIuyM7QQftpS1VvBlDQnEW2cr9PQ6M7gjSptgHwyHhUS6mH0SciPxj95Yw
J2A7aJ3pvdkg8VeQ/M/9agNDVWU4t18GXfnbIDU5AIBYgp4XoujThq1aJncy7W4K
c48B7zlv91Qjm3lnKwYaC9hIwD9a+qggSkd3/BIo+Nhv1D5EllbdtvSevUTysD2y
3ymtHHxVYGoZ9GZO+zjoaKvsV1d7PdiJOVt9KMMWqetEo+Z35jwCyTEi7mkFaFu7
aQUF6rg2XjDRrbSiHrcJo/HSpzYlgCs+AY56tScrq1r+k8FGslXNCgESi3SJTCn4
c8J6Qos9aOtWNU0K4A5LsU0M0DOR7QgCwg6aRW4+pwfIORWqEF+wXIWNDSJG2foT
20xCiiuPHUT99998PZrst35IEKpCieqds2gpVyThMETcBbhEoH41IWne3/QoyXJg
oElSE+T7IPSWBbXipLEa4D+JVMrhfK7FhXyr5vVkWVk=
`protect END_PROTECTED
