`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNrgHKJ2qhHwG07xR6PEuW34DnqNoH8PcuyuHmt1Bj0OR24EY79DcxIflvZUblA3
Fh+/nOMNSdyYjcBcxGgkLwd+LtyHyr787/j75/3947eMn1uJopRr2uUREikuUYUx
USXMCmLdRE4IzEBJIu3fIebcTkLiFvgHnI5IVEZCRL73BaNTeu6pt0sVDTNB1MnO
WMfS4EGQyS/eR3a0L2lUSFpqiBT6CyxhMap/pivDfWoHvCeGj/R7aqN+jeE7ePGK
SFAyJxTbiucp36kTzz9qPD5wdKgdDRQpy8RO5XWory6wqklAuoq1ZwqJb86hVKsc
WFqHbewz2tmR0EPGYak+vNgl3VZJ7NflpZRl6eGRfDN40svOR6Fr1NqAFUB/KrK4
9af7sMOCgayOFN/gKcJ0fYfiMY0ubBeLeDFmukt8zNWKmKyRUACCYxsrdwJH5Ut0
XNgxccnvoqTbdhYm/YEo1PcTBdnlIL0BggiulUIUFfE=
`protect END_PROTECTED
