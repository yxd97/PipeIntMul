`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwVWTS+kPYtjzsO01J0y9jB17aEqEgP/nMUk93MGt4UPeig+96f0RF+jw+WOzqp+
lvu1Op7ogz9qnP24dFQwPkBrp0n1LThJ/5X88R7qpuyh8KdI0ofBtyoUEhh3QlvP
NekRGZrNM021MMEDHj+fe7u8OKV9g8suvYMGVSlHv7cQW7ELk1J420subKMDeJkX
w1V3w8jHZrhhTR5QzaxhwIzLFd3OcXALq8oyzpjcohzjLJFYfV98b64Lv359AzDW
MvP9yBFcQtVp2uYatYp8jeYSBtQCae7TZAVJ6+yNC/wUJ0o8vKhAVoia75VUMzhz
kXITiI5GNgGuwufUIWl9o66VezgQT08EeLFFSH9YbjpUDijKweKo3tICO5PdCh4G
Iiobd2fMrtxNsRBf73Wj1H1MStNhI9bDLMFBp49F+0SM6Wv0cZe7wW8virlVDG8x
WA/3Y6pVATK5fpShSVtB/JQVDs1/HR//RRqH/vOJOr8=
`protect END_PROTECTED
