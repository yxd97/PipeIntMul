`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5kJ2YWqqoU+vMNNkthZXD0WfkTk/RV+c+S3QtHiu1Oy2SRT2jaxT8MWvKmR23AOs
QKTbfegAyh3gDZ3QFah79WDW85Ybf6moydZr6JOFngYoNPJvj/jIY7JpbJIrLHV/
QDg2e8qjE75eEy+IDDmB4gCMGL6c9mOPJoJcthe1L1BiXXoh7pj6Y3RfEmJZ/NQm
wFwBOL8ICxv5JLmqsbRnMJP1tV0wYTCGftZZHlVRE4xGf00JxNRJUQ6u4VBBuf0A
rmaiIO6a5kIledjpRTbk49xDwa/OAyI1ecgLXMtlImF9llKBbMR6uzcTTX5M2UuQ
KAmasM2z7VxZpxHx7JH7AoBhoHhrJayGgQYIizdnEyySR7Gx5XpnSV/zCWVr6y5A
wyJtwJpdq4JzMTzqrA+GDg==
`protect END_PROTECTED
