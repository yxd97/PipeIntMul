`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OQwTmmiqFx+P9bhzQshgebl/yNnC4SckhRuzWj18xli2K6uYz+h8VitbyzazisQ
SjG07i5EfGGHWqCsbhRs6QoAnHYBw+F/pqhUlygDlSlaLI7RJf5SSx1kKQDQvKbl
Teryia0MjoxCrxFo6Bw0chbSZBZz0ds7wUTQNQ3kRAmugT36r9CQAbZCJX6f6x7p
kbpVHoP68xrqZ+WK7u9h+pCZ9v/Im5VoXgkbRSOCpWtNst4ozcTuMYnZbh9En+US
keG5hHUsZe0bib1ktKr3qjwCZcEBuuNqQ4JVg6ed2i1dhXGTtrRItlQumAFk5X88
r+KjkOFG3dl7NGtS9znq2NNX3uhTJacAdM1CkSeIS4vbnl2VZaZQ+8cF5MVpnil5
aJFxuxv0hxthJ7r98vzd1NNPyBlkwm3N6ttsqFlt6xWM8J7bMFpyhH5Ztwf9sKyh
a8BG59yZT82VIrSrMOMD87jxiKDs7nmjJy47lQKddgzxRNUkR5O1fgA9p81s9KCY
5CuQ+7UFOa29thQWq+wXs5V/VrXS1F+lJj0eUPBELI45Wrfau0BhUoEEOuzprZeX
MVtTWupz02ctH/J5R2Ziy8egWw5IcTG8u8spPoLCrbGiO1f1buaYhqDXZ96y4GXL
cm2vVjhWDlGfFQtAX4d2snofxKHoniOsq5kdolX5jlt31RjXxd+tgP+AOM1dCfmU
xQpitXQIcCm468IvCuieze19IUb4EH7K+cvETaLqDqbrFaL7mnEq0ii/Rfs/ejyc
vmGIP0xtTlpg75dutjmdL0PccNnw3NZwTwV1BH4DFMBT/QeZZiv6xmD72z+CLG3N
amBwnVO/C3+SJivW3wpwIuG6jFTrOtJv0wRw7BNVPVvjlKO/NSFsu+dov6KvtK70
zvYPJgz3hNw0wOw8lSX+Kcn5Ol09iOpQUK65tPl8Xiq0ty19bb98hqObhxdu73zj
6YggFIf8UEVM4O24dfBq+5yvF2PwaNonmZvP29w7zp1T1ZAp671iFzPIlm5ePPC8
8QPgisF/s1dr4oG/F5ukHo14wwlaMXjau3gGFXMLM8QggDPwaI1bLZfBB4w2FpIw
`protect END_PROTECTED
