`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwMhs19g7dFd7SbNdj471BEyzXnI850uMu9RlTi451rIjZv1vZJ2b2WpuDnwGNdI
1A2D46r1C9PBo+Lxo0ZLVU8b7Sl8M4bcBIOuVWycfpxcTJDShM2dglBENBE+xaH2
ihn4GjFKNUHNSoO7tLZrr5SXEttdQ1hHo1ZYdN1VxoKWF3buuVwGzJrgutScLB8p
51YDn9iKLsIxAuaCsUNzwS0k3jrnaXd60JSjlsj3R4mWhPkXc1JgFTOLFjOqDn9r
7oW90aZGP6cbfOKQhSfA/fLczq6KalzCNbSfUi3Bg65bmWcM4PzVAl3H6LZPgoyS
qGgyavp7KdIeCiytiD0Y4AM1Pq2/JvrgNEH080ZG0Rv2MIokuvRE55MiDD5vYA3R
6+xhwEz4cw8Nk306OQU5E1FQTuzVUpFtBU8hMpHkkDZ6nqmkfTXa8bovfnlpcuGP
SVY/BsC7XDM8a2d+AG5JOQI/MPto7i2um9b5M5ZPQ6A8pUY40yxFgJZiGd6Tx67Z
1ff9a2d6lcvKmPD0DVEfhEdjTKdBFzPeSy/oVmiRlVHw5qkiCeJvBwSOmmVZ/8K6
N9Nd4Df22My7wAnFxAwN953LlCLUa0q/1O6OH37DT4CliVuXJhAOpt68d6CUfCK0
o5BdalvFmSyXfDacBl9gWKE+u2DurPDa39h4wifXmSDVEpbaDoWOjtyg3mVe7F/G
ljWxY+VgpYNb0ZSQQ5Zz9c35UVekfEQ1WDkVC7tCGbcqNf2rYrw6yvhII9RcKqex
eaTuC4DQGIl6VEFLWja/Fku73amVwb7GjHM3DXvXkL6FrLroBW+KH6N9LNc68nGr
eNAoyB9Rn//qVHu7SjAW79Rf5LGIeJ4sZtrmutSqIG0XYoo9gS0KpzSIMUKEDDHF
Ld5yt3AobNOI1M3k2ON7GLjNhtv4884qfNkWrKlGZ9/A5cASypSB3f73LKS5Q1fe
UqhWoRCDPaN/x0mOAcrr7wWdWHa91+FOup4jMqWZiPnP55TlUnr6X9n9A/UKDDs7
WAgy/qrw6KZPc+0qD62oZEQ6WyRVkTvuHSV+lTBsO7XYM4FauRar414eY6Qr/EbL
G4ATb0PLIVnH8SuNLj3u1lbCPAfgmC/aDQd2wQMkPJ74j/ThEsc/kASrI8muz/M5
dwngYXtvtkNYGUR2Mb3hrg==
`protect END_PROTECTED
