`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXkEyGeUFePgLXRTCM09TBcMABKTLyfuE2aSgAkwxIfULQOaYIOlNhQUKVa5OAPR
vDVwSiO+EeiNlbHRVISgASLmH/C9tL8Ejc4cvcMCV0lPENOqjSJaUv/tIqGtoWAZ
w7IZMH0ZBSXHad3HXW/TGIh//AMPJYar3j5GGJ8Vd9LcJd6PEfInh8hskr355EI5
m+7hjtwjroy6peP91pyxF29dlcGc5RA6RC6UjTaYzE+hFyKwVmR2SJsI7ofcxVcl
9y0rU7hcfTlsx+zhJXGgfoI50CH8I5BOg6B3xHo/Q5eIriC1a5xcHl8s5iNBNy1c
+EFLCM3i81zlIZSy487sCBrx4qJC9z/U547BQcrzS/Da6dQSxY2WmpOS+1le+YSN
dK3IIXnoint+7/4OIHvYxPkpni31i8fIHcUAMSTQUQnO+MZ6gunu4qkeuHXmGtpo
`protect END_PROTECTED
