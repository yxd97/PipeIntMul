`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KEuqEKUqKkOswcdUN22qJy0YkFP67XqHp+UI35jXecMReL97+l5ZhCOkOYy2P104
luq3WpWk5raA8nyv+A79RYGHJj1AvOyZDCudGiTRT/dWbwnGaCrL08Rb8RILcz5o
hFtnHMi2q+jmEsTyl+sMLgXpob4AAsMD+Q3is9V6ehE6zqo+cQGHIo+A0lkBYBe2
vkF/ai31UpAYadqQeoCMAR/Eg/yLy4yYsLXfw4SQ6O5fVTdVAYySRhLrKgML1Mhk
wqHr0FKxPOWf8+snfsWG8tlT8/uewIJXi3tPGQWLSDz75TNF7h9AwKhaprT+zI8/
2K+XBc1q8iZ9jOd5j5gK/tf/w7Oie/JB6BiOyye/1PUXYyyQTbOUAJvravgwiVkD
dexnMrrvsH1Pz6a7zBgXWhs3eLx+9Q12JMv0/LTKW2tqZQjTZtnjhx6xn3i3BWre
Gz114Y8sonAS/fd67QWqXOzRkVQKXrF9zmRK2FPKELS/bVsYIE6rzevEWhPzTFr+
myvh0gpaQOzePlbu5aNya+srspaWG2tPXz4wu8PDdQN2aqXpAshFZRyvhHyWe3TW
4l+DcpZRrnoEZ8iLcrUWp0ILA88Q8i2jBfILMmhZuvzi4jRELctzMDXfwPL6HZkd
IfRWV9lZ8ZQ6E4E3SRGYCycB5SCQ5zUVfHGtnAUFpxwj8/r7zhd3i/7aqVeVe9AY
UaCvaMcQF+IN0JpUgMSirZh9f01zZEYKTxEJ9GQuOlf7XDYHX1iFKtfouoG+3LCn
YB0sVk69O2dxAVFGh0Yh5vxhbkjnZpW2ulrRRpfzzwAOjaBzIwVtc0SdJ74A+zfL
QvhOy5VZvb6EYXMCKxH6B1bv1uszXgrGQnteVE7U9crH3ge7MZme04d1BYDHsWwv
9DM0xu66n9d20+7IAIClyAwH4Miz0f/I3A5DWCnBEda3WFSwXHrhV8E7BghjnoW3
euRbbIlaEywqY+7XpdHWKxhPnbRjRY9H1T2IbhNTAGX1PIu2dH4n4Xl25voFwJ7E
FznnwMfQTHWxacwZwO9TJAEFkyvU8j97CChColEOVU1R/VYgtSDrrYnsXgx+FSUh
XNyZm+z0iE5RVbaEsbtdAIyTzdpQWDFbnr/tPUBAhm4Vh/qH5GOmtYTGssjSPieX
dLP2Uu3KTYIrGrExS7KZVY4DjjpWEaFR1nrg/GG+ITL52NagV7WpXGpduX0280xz
QrlJIMoAr4wH0C5kgCltjY9J2U+ISdc9BT3pFTbF5KUxXcFqAu+zdCSlA0S2wuMp
UcyIA7qosbTCtbOTKfllA4o9W79vX6vjuP3ruPlT54z7v06wB8sIaomTmuhJRNVy
0/8csRgM27XvreKPa09AtKoN37jEH47l/WbrNri/tFbEMa3BK5JEaUyOj3kdqDCr
HjSTebBChNaCrPXHx5Z4HcuvlE2Uw3Er3sCp1iTkNuM038aipHlxY1hUkRkV2xrl
VUdDTjTGRM/n3udJTu8FJSX058IasPyxRa6X9V1/d6PnnjUAShlk/7VXvQudokrA
IBqAGEjcDttP+J8YeoRPTlxM7z6j1PBjYCVpfYUgray6nHK/i/NXsnYi6PnXIR/f
gcFTAECt2zu/xlRz385WcqcPliF9d/ICgnhcZ9v7bUOjPr/g0lYl7pQrUD4u4h6X
qRsSrGDKtQIlxq/uZFoIZYHLMtxBd5RD33NcViStpRl/hyoNPywStRKDGAryJMDz
GYLHJq0Qw9M3huawunLfb80vRbfBezlo8vwQIkWpIecNSRTFsqr3Jpg3RrxBpZeL
XH68ptJNcpN1bVhn9dTLaOpR38f7yD2ZPRbhXqloRb5LlokLORvyY4gOti+LKfbZ
T0ZKpfARTEwPoBiDMJLr7QlsbajCLNayS9jZDRVpzt0UtBLH81OwsUSESAfbDaJp
3eeNTGnIyoxe8cYz7bdyUJ50uXEDDFvgKTG/bS4STm74ET/D5nRb4zAOivMkAZl4
OULxRf2YQm0RfRqgBXE0Dij33BC+WBYup7/oiDgw7wH2Ix5R5GJ6pzjoe5AJIoFk
/nrr6RBVPCZ1ZgRMGQo0NLGv4gOCM9T+WaW/T3iSr7acu/aiNnpyTndns2hyuB1w
a5bFuiGyxEHaiwvcolGK5pfovC/8gn/mCvjfqyoFHcSe+GC3pP3mySQGxWA3pWyp
mgFgEb6x+m8sMNeqeTtqRn4k1rgMw/B5fI0a/bJFev/VRCjs0DorXfLlo0XzCOmR
JxICXdObbOVvlEcwIuWQrf24nQB0b5RlfV/7zlIq2BzCPYB9PxK7swwChN6qnsuv
0jvvdknmDO1z5LqC2blRhcvWlw0WD7g0mBOW/25nEvZ7jwjEjEer20mkrB1YSsDG
6RhvmW6TunBm6WPlkzr2vF/BDFu1A17MLkg0/om1THfevUM5zLRw2k1L07m8leiz
PhyUQSgFhWGsAX3xS1fVjDqFxjyWjxJkSh0h80gsFJ2chmnid1iMF6Zs1tEZ2seZ
LfUz9UT028r5HrEljiypypcHvoAu0qY2nIryfAzuJ3LjFz58+Sl1FYhnqEiERNa2
SHN6d6NRGD8m7YyRecqakz3QDxglV4waUe4DtGhxy92YYJC/3qP4tBMEl32mUh0R
Xvy7lAZlS1xjJYwp1HmpjCnC2jzM1+uOj2dl4z4Ge557gxhXZH6F9NA8nD1VY0u6
A0gn35Gq5w+ELkImBk1fs3DnLZ0aZGJN8w79tOnbWZPaRxSru1LS9jB6w5Y2t4QO
Fcctd6Z492vS3PwTFscJQtyuc1pJI3/CyJGpB7YuKhgZm49LU6WTmhP7tUOvDASI
/+fP3+flLPgO6saShKlqa6883ZWGHcx1vHZr0yeK3TS1DorqpJ/EiMcHREcj4RBp
KOvwvy7xaHhY7UujbbEpkmW+ZDdpA1ojw0bzmLFpE9RJ/HoG1arkPyEEc0XsrZ9W
8xDA9JYZwLsXJNeT+ayZRSUvTNWV+x8pMPhRv7osdbB1mCCg8FqJqrHTUWbjXBq3
0gbTZEkGu9A9Wz5BWbdp7dPEcMaJbUDQOjF6SFjkA1FVj7W3fl10wHS2FzVRZ07l
tafw7nhUisfslnaNGeTH0BJIgyOLvOlb+eSq3eohG6apksaBxce1Jl8FaJ3RHBuP
z2Lz4WEeLmCIZGN7PKgcrcM1qAMWpJd98N97yZ6pK0VrEzaCNjXAQNG2stqPKESC
mNh8yxjO74fVIok6svBkHXp6Zo8OfUgl8Io32WRfgP0YN/bgwYVF96AEYn/cU1Ue
y9tQqNUmTzY3Pug2cOxMXAcO/rG1G4qcPATEvh9H89Ne3LePU6ziyS75NGOGmvkZ
GLMFUNdHtEZm9JxL6/LXp/6HlHk2GeFe9BsDIoIGDbCYYtjLBzrUW7TJAV5QxspL
Ogu9Zrbxg5JaTkciEBiRkzCgbUwN0DVeIlB2N4+nUNZiePook/R9OT45v7/qx8Wn
0xW7wRKURDSD4kr4MTMtK11tp+aKmRSf1GPd+KKJ+TTzywVsKnIwKmX+sl2zhho/
B10wW3EDgxqZMMceZyNe2umv5i045vJxFfNnaHpqARRTg3mneOO+Dwe+Jq4AFJ3k
vdcm9IQHOhhA8shzwcNOSFClNaifSFCcOgZ1fGNGDyDSQFKkH6vv7hgLU/anmAzK
aNpV1jUTz5YRXw8CC6vI4WXw7SYLkLtxfRYPf3AwtdfDPrL/7mQE0b4qf91T5pJr
uWoF5DpRbcxSu9xp1VghsCBll9tLZRmrsIP1FrJBrLBwoX147OOgUxjXz1vrn8bu
S3KBYK2W1IWuiTNKBLCq1r5UXv8d6N+YxRZZfNX4Tkx5exu/eH2yNUP2sg0MAop3
0U88v1B1mcgihPclY3OFRBqS4gpQYNXRD4RjvAwJvVPmFgiDaq6a6CFReCp8U5Ac
vlkF/a32E9xzz1G69nkgEpWFp+bxx38cbBlzQ7k34dEpfJcs1vJ5fSqJj+KcBC4s
A4miDLMcVQwyaiOMvjNGjOQ2ra3g2+KMl5Q6c8K9cfMcegHozF4wMkB78SwIxiw7
ExldfHinHYT2T0ToHJvqQ3g6w/BD1oA2kzf6AWmCvfX3ELkZOY+YpZA/tlJy94uv
1n4BdiS8DiSKcCC+OreBMD6o4ZcBbIRS0y5Ysp26RG5xuRyzCjAp2s1zMOP2ojM+
HYPcgKIBRaITMj9NC6tThyGexUnDjE+3bqLGD95vcVlfnSBziMW8RIITCnCDqiBq
fhEHkgNV/ZdeZKc1k8b84E1c988RFeajN+pYwfOZPLdt6O+2X8k9rgnfLknLi+tY
u9luNHJ8xwrPD4IzlqgCsfhp8PzDrFcXWazWH5xjZRzMbaGqk1SjDrozhaWZygmg
OFfb0YhEK+ln3+Iubrm7jSYi2mm+hP6jQDtVswv6iBD0KNJqsHmYJ0a+M9umK2po
Dz3ED6MsbatjN1p6DEei6TQa5/u7rA988LsCGt5q5p8jfMZ/o3JbLZ3cokuWYcfN
Tnl6bR7bISGomAhz80pfrqJeV2FDnRC8BbJ9xP2Ytg4jAb3n1A9vGG6poVqUYRUW
wNkpzcO39aUtttDyrtgp1LpqWkiZrdoHCiNR65diOuFBOWjetFP7XEa0RK8qJExC
u9WKvtEAOsLx8U6MEYgHyBXmQO0C4dnKuArhadRdjti3b7JfPG7sYxy1NGUYrPpN
zkEnawyhtxEOQAxYiH+lTKCZEHbya2HGJBv6fFU/1J2pb+c3W/rgSDswwrlGe2dA
oCNgFE5IRI8tHe5+oWaK5qKfHFiESII+7IurlPVEijL/55rRD8ykne2dt5TDMPt5
HAh12kIudicQ9xWBgo3Wwon/aC+HCRmTEqUb8+BE3q9z1K96RL54+QHQkp068Rw4
2bDXJRFJBFowVE4gAK3l1piUDS8dOYxOt0EaAEm1th/amMVGHt/l6YWyPwB+9NjH
V5mUywOmCwD4zQ5HyxrvMOyFhQXxksjhzWw1t0bBa9arL/bV0FudxIC2Vq38ObRn
zWQsVYu07TPMQcAJ0PwJZHSaPRpCegty6tJZegHELKwl6+lESPd0pY2A2pBosvZl
wLPZBUl9aIMCy3v+BFZJ4DUwuHftzalrLBC3MmemJKL2Tte3d1s5ja8LnZiE3V8t
do5MeaE3hec7UWfGvLZN0u0frnz6xQjbfWAX+HVBQQO0Ckb0WOJhdULcbmope/Ua
568MeujnH9G2iIob7MsgxuHkniVC3vBM+RswfoOHUAFiwKT2cFjcylDji3P24i6C
PS/E6CXQcm1Uf9R50JcGiOXdPv8qCZ6XltHDL6S1iG72bXYMQmnvVtXIhX4OEWKy
qXTghTQ/hC9N4OsSgg2LVs48e6821pNQ0vKnZNXXfKYxeDbYKeSrFuf/Bhab3DYV
IVhIbJf5kwUKa5l9UKPTl6uPEqBubz0myNt5SEmOlhyU2Nl7TvuU3ia5MwGnZxPN
lCYWIM62gdD7nX5fG8g6uQGCf4FitkioMRH8Hz5ak/A+QWrPOOgf9JD8HOHIirQw
tx5YsojuQ5E+MuToJZ/lu9YCKP9S/VDUS4gUWh5Y0bGE8dvFpPSG7A9wtPUYpYck
HJrsqU6TVfVTHyFEGZAzyQYXHDL2KETTGXrmE/cFkxc3fa4KeEWApjLp2hcB6JwS
vS3+vtR70ofD8XtbARPTJgqzQ5+7u8dbyXNISxk692WNfg5F8eJJVfesqLgdR2SR
apROZZO3lK7ZdZ3SPR0PT4EBMsV5zTZQ+aW4dgM2IDFjQXNsgnmdT0Zrh3a1Zezh
qx+WmQgI7LbhkJVcV5fw1ycMa+jfapq/Y8pMCNR1cvmZOf+oDDqEGEOuX8XTEm70
OtDX+qrZAkEQSCEedrxc8RKt5W9vigVGv1SI7J0glvpp36yQZ6uPazxpm06WYQq4
+uSGOzKXslpDW2qwfcPBQ+0ghUlSFvaaTaQoXt+zQJKYP6NCrpgbYGFX+1ugmZFv
N6njnVACBsBIhBQm7dAmefKhlYdEmJsuD3jtPMkLNc5O+lFItjW5z6jRyk8xsxhp
ewXVkyBRhjrVux79u7aBxTMhKZy+2VZB2+hqwJm2YLYiQ7hn7ONRHDfGCrUa5Efu
7nYd0rLmRK+WsGE3NEpz7KlYPtwyLKByLMXbIkA9bb0LRgcRSVzG/qamJJuHk70u
TN3Bv26rxz+ZPR5z/wfRH0UoW4jHRGeQvxPoJKxyRTgiT+IBapijfRY7KwiUjSuw
9ZMC3hr2+9fPq9rzdnFSL7hZBLuGpfeA2QkLE1t3a/lR61smAvojSr0c0VhjkI4p
8Yi39G7H7+xgLh9IHn6t+SGzkdmnOikwc2l39bRJZAKX99v+WEap8rLEhNH4dIuW
4bLNA3O9ArWRqKwm0m+7arBc23wqQcBr0Ev954/d75G795JRys2Ot+sUQwqonzqk
11fcOnUlJp/eXe/b/LN3QbIqD3hTMRpb2RSyVlriwBeaH4iQJZCuECFpp2bLyzCF
c+itFJ9bS/HpUY/necRQyAi1DbZeezx+BU+w6DA6JDvj3mNbAI0aIfgOSeMVbdcW
JNaCv6COXkIG738LShcYTQMKJP1Tgs/ERVCEMBGFSEpB2Vr4Xagvq0GwwuCiseBe
63Sqwjh0xL+9O61VasNsbxlVJw2019mQcusFJuvqXiDdyQAxTQPutMjGeabLQAjd
9p+tbyQPUNQuwktzGI4MEzK/MY79IHmHK6IqkYbYF6zVTCGBEz/p2guLvonlBkRq
DJ+uYoBkex+1mSAsGLgrONXS6X7lTKpUJ+jywtHqlKiOLkOi/80F7bbPEs3rmq7g
BXcNOiudQm5Hpz8PJZ4Y55WMAPjkYWLdcnCZ6gZ44sKjsvH0yMrv2j3FZoqkYZwr
9S0LoXAZ92hbFMiPfv0xvT9Wcte4nAuyB2qbnZvFYzuTEBwh2M+RU33dqve9CYl3
J1CS48mIbRWGERpzI2JnbRTM1Sg/N7G3mDQzjyTrLFKJfmVOGk2x97PSQxE/Aj2R
zxreNqBVJmoxw9h96Mo208AFfKxVNAfTJ4KpCnkAybaRfOdodtbtPfv3FDIVMxJA
9e7BE0BMbYa8h+HUrFKjXhetB8/lF6BbA22JSr0rpo3JlBXxoM/PqglIImGnzxYE
xaby9mcVYm+vpiR9vFBkLvjUSTpBTwFU8I/zbj/PjJDywpau0SEXSTZ+pxORsBNS
p5sIbo7Mcd63pQeAELkQty0EtkOu95uEFtehn9PpcUwOlu6/+KUVP0p5UGpQWZ1D
vlwmSJYHo1/noPDFp5t5I7nX/vixnM+1n0bo4fO1H4Sj+4lzAojNVr8QZ/Of8qTS
0mgGt77JXeBrQYUT/bmQ6i/aRMYA1uXGm1XIRqPoi3g3GL0g+swzmQtP02sQ9biT
y7GcRzHEkZJPrentLdzqResdgPoyEpCc81KJx8PBQkDFGCoWhqZ5tB/UK4lK3JDN
GJa8+STE5bi50IOWJfQQ1m+EDsLc6mHYAN4hMxrUnZnKEGuHpjyndviI7tLryOkB
ef/Jc4uqesKKVlAE39lQomICNYJfcrLIvgvChEZhLOakjPFTp/eDNwMoie/H8fBn
wzHljP4u1XedAcsG8zJbzJ1TuXs8TQyXEdelAVDIUEm3wEhPURAx8duBYWRtUMuW
BzelvLuD6NzawQYZWPsskMLGGS5vQe+f30ALvlkQlWnT35MaqI70chEaFLlfXIqK
qpc9CkMJ0fx7lX4zFdpBGy1+KmGYV8y8TuU8jKaKYviiTPvlclmfniUlhXtssUvh
AwgLZQyrCk1aE7clgkH6epDn39KBgl/lqenHaFd8n6OPHsTNtveay8ubPr0rPEOi
mTz68uOTAQY9kw7NCIuMVV/AHOUb3jetVxg9E9AMauILAPVlUiasm7lNOJ+ch2bf
VJ58Pq0Msz0+D5eo4rzX+Hsb9Qen5YE/4sZmZgQLeH240p9iEYdaFdA8g65nMK7l
3x8aYrdiHcoXKxFYB7XbF6Il04zziQG3aOCKdccdN9DssC08YRB8OGaK4ygpr97m
XyKCmnrxHTruQv6p9oMzUsU85z/FMYSjjFLUL8kq2cnTBP5QvTMiuBUXLGUMNgaQ
ASpgjr7gRHpCftQR1jLCcfNSRPovX34BVefUsGJNBD/befbVX0jTzsuwd36nuq08
lCyIN+78PRdn3ys7B2iLHo92eb9NOT8XsOI2KiETpoNgJq1TbtyqBvmMXfa4eNg1
MOJ7YHCr7PjasIY27WsYM5qhfRdGNJKkcE+kj0hyoxcj9spCCkChtEN2bxdaoXj/
mu5ApTvcqi23/MGcdCwBI5qWp3FmO2Jr/tJvL7uuFdLUDzaQWjjM/Kb5+V8rLFFo
1hCkWIqHj8ewfCkQwMrdaCeR8KiGeurOgEFUsvFthar6klqvNsOfG7sISKQ6Q0lZ
hxJdc35ukymKwTIVJLAYYdFt03nW4NDeAcpUs8FirIGXqls8AWIWe16sBawCHIAc
jT0fPJUcNHpW8B9TWFK+KNY8QlEyqSFFqifSnyLBUDSYWwTdV2eopRBREs2IE9r3
xHeIEzalf8H7+r0XWMFdb4AhcyKXNrBq0JS6Wd80kkHQUk+5UHySMM64CQZW54h+
ndQIEtjIKXRSliN1EhthOkm+s/AY9mVChVKqQfNHlowCKXPqcGW+sEMxpZ/1ZNUx
9qjaGJJ9+5xIM1Fff8/7zYy8YAcIiarSvoQCDq+0cm635YVFIhwVzaYdcrEWiDXI
zllpMOjFKWpRBnrJqifRWp81b6tJOw7SJ41RRYe76i1ZAQXAzqHZ7vcvpH6r2ZGb
0+xh9q8xQDd+x3kwieGRasXq5b3id4VMu3mF88TJgm1sqZB5zYngjAJIt93L348x
/2sh9g+gbSoDqLEjP6T5O1OtPRoZpfPN7qV4xcziS2bXleYqTNly4nUyDcMG90iD
ETNP2ZX8Zh5WshSb9JxpAGHpqfP2o/NsL8aaUjUj04wWtY0iOZK7szaUBOjn4KGL
ENZZxAxuJPqIbF3f5oefpC2SNa5AckDUpOie7B0Eogdb/cq+HG+pxO5GE673Xykx
IVztGD1wS20qeTveOtG3c1JSfOIEz2JhveYf9x7emUoikwEbsUbO2Yzkt3vRNc8I
wtCbh8lOcQVmuQHDArakE8Y+aytosQA8MIUt+/gpcEkd8Ck28mEjZw3D3lzdj3zb
aZkdomxa9bcd24CtlgVsF8wZmIGDdO4redmhEMh8g5unjmwy6BKGT676Z6kmEFhR
QttdVzvEXl3QAULDRiODOfoibH8c5nFo6TmHwLRq815rj6CniBHqdK7MABZKRgbD
8JD0WCtXjEqL+IXuC6HYZ/PUCiwtiYMHt8zLG+XO1i8ck6MPbvBH0QOgZw4PvIqp
GVfkPM80oTlSBI1lhZs3yvxKnbqVWs3g/KhOVUtyeyq6+K1SK39iYbGh8g1BTZiR
X77X8OMdJfjJTq2t7CRKtYYOm2RJdEO2k6oNzUfas5BY3MuP4PJvvAvzJVt9MJy4
cpSzK8vt5Bh7kGc40X1Ot9mDrdBbRhIB4paw1B35E8nyX24Wkr87fsGPPbTUM2s/
72+mexlGA0Lu5EvTmKDVPVKa9r7E+7yYO1UWiZIFGGRBU4oe4RzsyZN6hdEfwr7P
6zY83MGPgnbsoYAOnPFh0rKSuWvNml21sWNzNaTSRP65ObZsS78Occp1KNthJRQC
G/3acSnXmhi2bnwotpMuiv3cFdjuzgdE0GulkcunwbtIQK/TJlaotjXjZk95lBTg
4NXQMc6snMwj8gd/nY4AjNlQdJ6VEtE2brApcXNgS5/u8L4I9f273acjzk3j5Lz3
tVresSjHTum3ddJqd+TQwwYnfkEUmPacrVl/np7ZSbaZWZNyFCib6EVjVbbokBGS
fY6vTGhvNpDmFdBmbRwQ/MXkCwu640Da4YX3P3jmZLTInQl22AOFATyBgiinREUH
QgKH6VkdRKJqKdJ69TsRzFszglPC3BDt/DvlOko+rHHXAudoR0mwisomOzq6XQ0k
eySQHDRHcOcHL9QFIX3mULL2Cje0fZRCqaoL0IZjbRr/CeRaC3ezqjPNEvQK062h
UX78bB4ZhZJtxbDNq4xkqwL+agkzSGo7nTPXEeOdWo7OZRqadegXc88QP236Tr/j
SP6bIEdrddvqowPjVP4vCgqiI0xCTIPTGmvCLZdOSxpPYbCOZC1VxNL1h7i0WtsT
ObLvPH201jxNauSV48tHSSiLCwSmLP21JeZq3d460tL8+e/v2MFXtHuXP6NcG/Iw
NnjzloDnJXwSLs2vUBlQCtx1flZbP9XV8mQQfrkMcYNsIkKYznzgm2MR8cq8MHyy
XbakZ8WNLGCC5qYocuqozGtRlpvGBSRQnAHGYJdpDLo1a8K3wiD24dEeBytWspYw
kU5yHeYR2OsTrbaCxSuS4x07WgiRMXnOUiUbvaq48ijuDIbT+k+X6xmFZloqHZSO
FlPaBxyU8IGuMfA+UNas8xFyxYs87grpVCUGGATJWXIp7EQafk+E47lfChaK0n4Q
cT1Zrr1oEjdYdegE8l7uQ6Rdm141W61UjTeY7Q6Ak0LciYgxX+g8CwdbFJV7rtOC
tUIvMx/WW6dr1mwocTC8Ru70TQC23b9ENuQuqxC+PnMMNWUtcpB17R7kUVvcJ3fh
q6ELP7CX3F/lJRtMlA9xYSVQeouARDh3UFF2lqqzHTdLiNL40gfR6veQJ2MJmLjA
`protect END_PROTECTED
