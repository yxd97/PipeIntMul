`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FQihP/hJKZDvialzjZSXLj4pPlkeCzJdMw5n4GcEzG1Rzs7S0d1nFw68vDleaqIK
K9EMtoQA8wXDWtFj5LyN48TYL5w4xK6nXVGKfQY9mZNea/k/vOFCj+sWZ76XSw6G
Ntn39O8oFeDonXe3Xtlj/sle8LPafdvrbF096SqJv9kG/owtGy//nzng6HmT3FcO
dsT4Rm8O8ok/QVTJHJJ5dqN70pQrCaxjyWmWF7RaMiQP3nhJkhY+zJvK/iu5owsF
Y1HHNIuKDpuE2t2Bpbye+zoiwLnhtb+hcmdAWFcoPDgz9hnyXd05hc9t01dsL+gd
hm0Hpr7X0CflOd9ivTkA2LFsKXorZOW+kfyr+B8lghX4U7DYDAgcP2odsftXMntc
EXuxAxX/j2t65FcQbVVWUNEK4X7GUUU7daoIUoNPXfGCPC/AbcNpNYkQYga0PjtX
ssZs+dPghF2oMAHkleu8ETXyjyFTmrOwjsM5A2vGOTPwhPRgn1ciodh+fqPwNB+9
q1TkhiKCSv3xTSC9Ll9raoiAMP3xqBri9uUmVj42Lum5cUvA9MaXDwyYuf9el+72
7qCFHtiAxhTgP/HFaTwvQhBohOGsMLO3RKChrXjcGiHuOaDMTCmqoCFApAYPGHdw
lr67nA4wmXLTDAkwsiCrfxMcXI3cOzzca5RTk2WXINr7kHJBuJzxxrXW8Kfs9BIy
OEHb92juqLkSzmztI+PXS/DFVpxfKOd0bPK/kP3Bi48=
`protect END_PROTECTED
