`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hVWF/OtBuXKUFNGnlIveUqyoPEPJTstof3Moq4xo3WxFAxookXenKfy1DH06p7mz
dRcP3IblqCHALaeoDqKZGoVYE+91VB7GuAcxERdxE3iXi2p6vEdTwMmBiLbZtCCz
QEVZFhSUaKQvU9fpYs0obw+h/t75F6mXTM1E1co8VxMgTiEqpXdYbmbYfmeJHd/R
eWE1LiIuNxjwyfZ3VQpxddWI8ACFMm9beu4Blk2IWZMNjgqmd8l9xq76ECUuezZ7
fUlxRJ9mV4UBbxf55tn1iTBwWKnZME+VWuwR8C8VS4JjyyhiEpkZO0guSBj+xyHE
see/9d651rBCs6pTwPLo6UTFlTYT2vYFLprleObea/0rXQ+jhJWqgMjegzcSYdbf
CWgb9pssdCVaMV2/J04JJ3yS8yo+mJRmNrb7QdcS84yTkh5r8HIyK6bZDDd1mnSk
3roMlOgzr1Cgu531a7tEQsbTDVG4bCiVRP3W35y6OJP2l85VL3hWkT6ZQgifzF51
dUusxz6JxUGTC4OI4l1Qcw==
`protect END_PROTECTED
