`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FMct14PJq8EmXr50+4QCUzTrWSHJt6NFgVoTizn9RhvFHPrtbSGQelXMaIBF+9df
nuV8sFrVbUurX3UTVSj5KUof9kkP4hiSROiDzrx4nMW9Iv7oFWKM4v61/+Aeizst
v+LSMisabMS0g0ARF6jdVjJsdR+uglr7xswDOJefcMwvhXT0+y8CrUbeJaACNvKx
jrldJr3b2XLQK4YLsLF+LBuJAh1dIv/uhCRzNpfJc6SjpI1pJVXico+mB7aqLwkk
gy/Hyxy39pn1zoT0s4YpiNXC9VRbMYWIkjAlzP5WWW6+AaPN+hb68ZvU5QfwSSC+
7F/e18nE1DgymwL1a/du3jwi4MahTBCWDWvQ8VBYFdFxLDVYWOExL1J+6pxkOU7L
VbmkkJ5M6oxbppoW3bZ+curztKUfOKCAYz/eUMFUNnNwPUDMLWtg/zyELvUbhCIv
vNsCOgH61ouyvRJGTvsz/kyaI7K5FNavZ81nYQUZozZHfvZRsU+z6EqTcGO9Bgex
EaOBVeAsDtwSrsKVTs5KJ+Zq1u7JwbBdE6VhRTUcIg28gbD/mP4WswL5Kq2JUTl0
hZbH4YpBKK4EgKgW3zGMcuVSQYIlvHxDPeM7WfujSyegHENr0xn5BmKX/zdfpvuH
WaSG8R8rh300+nxXppipNp4rB456Iuv0rWkI6BVWkPGEMWYL2wYdCym5sYQag6TW
SMzSEFIwu35NmkZqDibA0+BaAFrQscI/FlEs+ljJ+4w=
`protect END_PROTECTED
