`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2aeOPfuVff7Tp1yJ2xhUKzmgX4W+7TLTYgj6qiUp3tnr7UFqQ/n6vwlj377N3/Js
ICsaOr4JDElXOC2b5tdi9F5nx1WxGjVTVJv6/WmtBGNkc11WeC8SueRz9/XsHrsn
nzdzSc3quFXs6E4ES4znAVzLb8E0cqzXOE9zP98iQkkp1EeSsWxHkBUYGWIhjw4d
rPuTlMMw4yWcWeaw0vVnrOz6oeJ4JghdvFqBcJwqltl7lWRdge6E0/NczNxgvB6g
69zXxcWQ7DFDQMgZu0UFCwWqWSc0l7TBqxjIXZtWDDYg1fb0jsTO/E7zQY0SN33P
4sXskU5OlyATBDCWrz60T6KCQkE10CcA3rLZ3Y4jMtOeAajYlb9oAntGjMGUB3UG
Fa+gCIJ36MtocyW5gy6KpLVhYlMttTxykb7VDWKoBgdlI5yX8bu7rd7R9TI4t6Ox
0uVfbT+cZJVaT67a0L97w1swfm6j22ijUILOQ0Ge6eLgpc+1iW8USywY2uO+tMH4
EVBaKIQDsbj3e5Nfy0MCi+2zmGVftSmVSQU3PbWkjKNifWA4hmMehMcwvYPP4lwU
c8Qu6clz+OnDhFkW2g4/+pc4bRsfRkxov/UdJE+SrPOJG4kcxUBKWyL1gExrPjoL
qnhBohwjE/QwZXaYhaKD742WNiZMIf0MVMwz7ns4RG+ekb0VYyJ50L50MuPZHfgZ
X8YHBl1YBlidCiEIS1KJz97EHK4kt0RVDbqZRb8j8EQRPwn/IXDUm7/2XSe9ybCC
Teljof/a3D1HCo2TvZbukbL/tNxlZDPQuv5anQLMpzi0sTYMicYGtzhE4P2lx1O2
FZZD9+gbfe9F2JPpxkKw/4aHlE1DgK6PGPOv2fDEvk8mh/RhUyLF/A9RLW7GnKcU
b55HiNMU04U/sBOOE5Xbfklq21/WFxUxBd4oNN/nhzZNSJnokZatYIrv6q4u88qN
wRvO+Q3+FXopO/znsQMdcgbf2prRGwXvV11PxLHPgxCnU0fToJOS7MVLW7512cyy
j0peh+4yLM/WdZ3N3BDx2leffE2k9OYWSuEUd+Oo+yaFYYZ8FxjrixKRsfX1dntp
CONqbphOZB8Ylki1nnkPdcNbLIdUU/8nJ96HZPw/ImRP550rQvsJ75DX6Qt2a2Ha
6/P1Z//ltwCKOQpuY1w0rLBss5AtuJJtz8k3GHsQSYtEbtDEnPx1YtsJDaSNE3mt
gi4I/M7bSs0H1l6hxQz5L4TcOAqTCk4gWraG2zwBQyExwnuPKzM0QpQtnVKH40JV
Oy1a3iNuqVIc8k3wd7cJ/OCioDFe4MRTw4nLrnJVgA/9o7QVZOCM+jvuKvPUtSce
+ZYt9Z5r1ra074LRBdUVZu3qyhPyop9+VelR844NHB0i+FJz60mSA8Z42VjwB5Bk
`protect END_PROTECTED
