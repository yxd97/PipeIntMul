`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fV7L1JO3Y2raGnGH0gskocb+nZM8L9LxhNkC1RfjG1mz01m+gGD/91js3CF6s1Pp
gTRtZ7KKkkEzugkzYK9w3oEovAJQIiaZe+bLktf70s9VqEA8DRDE1geD7SwpXkuS
/B3zMx7Ab9HDTihWXqIHMyJsRf3rzKnGL6XH98yW4fuyNW79JOYxyYrKPOXMq9+d
c6jckfjf3D+Y5/GBTEOaKyiCp/dZkYEoX8u0X/FgxNRSJL5VOSZ0ej+7HJZz1A9v
TUKKZfBg05c4DFWkUY8SnJJM1VQC8KSRPMV1vpmskfQmunb3HXclT21CP/h5Oyaj
JXrN1sBqornEA1UYJDrsLbHEhdtPf+B96/iWdA7WyrQO2vCDaX2gNXAa3vX4hABA
8hWY40e1rH6S7p+G54KB1W0XquZelEzsVTSYUYEr9vURgl5geXgwXjDi/YdCdHMj
782+M3fRtnSMgLUtu0INUEi79OuV3bjEEXCQCgzjdTKJFRC6aFZf8ndAc9pF3md3
5eymKiN6DSSgkNsyrKWDgHTAvelmNUSNcKfRKvmMiCoNpbu0EkIQ/gy31gmvIFUe
B1S9d4HakSTjVRPlqyt8lIGWI7xT3MMaBBGK/clzNntW8ur77/9WE4qNnBZmO5TK
44L2yfbeLiBUDH4hN1dCDFzRAzZiNJ3Vaw6cGIfBsQrkDEOXYLpXBGf+nw7dMKfo
QCiJdqzvoUivk14oendAdMXLdGI4ZxIdSq5zkcS9/a9amoE0XyEvt3Gv3AB736pr
7QaNWH2uXXuxnxRGQWikQg==
`protect END_PROTECTED
