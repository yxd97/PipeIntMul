`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0foF56BXkAYI601zN6/H3sL37wtVDg24vM6LHhj3yddWer3tUv8IOWYZMN4yI/aL
aIJRaOXcNENFWodGkoOS39e8Qz5TIJ9dAoKFoxrwN1GlB6DtLuxM+8zQ8+MHOIBR
FQJ+zAaMGO/ng1SV3gdT5DT/czpsI2aajm4ep1SGZx4k0vrj8SOaQ8fBkptaUzo6
/POtKi/8MShRsSTuodnxtxHc81C0aAEXF+e/9T0eoZQw2QP/qVDW1nwNmNZ1wptu
pQZ+5vTp7MhE1oLQvIsb3cRHHp/nny90SbLfWd44cNyTmZUxfzkNHvxreOJ4DD5J
oB7Kdxl0aP6F/w063nUzc7EugbPN7xGp87XZqe2vaezVjQ15C0SRo2dZdmtkhOp9
wP+0w8xFr46LPoEg1mLPHv7XJNmEWv+h995nMKmdukDvl3JCEYnlCM3LhF9A2cWu
Ndn4Vw9J+RISyNC6Xdc7ID+6gAYEsvNxnOxo+/qosWM=
`protect END_PROTECTED
