`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NQN5a9mCVVJAv2GytKzUFnHF23WpXbbm0lBwkBxpfsf5uSFOo/CDl82qFCuFDBtz
WgBvz8gA6CnOTUAFQlLD8hSEqcWytF1woqDhARS6F12PLNfDmQsK+0zRGwzVSjh1
5HJcKCPAtAGrev6aCFMB/gbOROHZbC6mXJTNzVsf04oJR8TEXyOhwpGAYXcOfN/C
NZBMI+pas5Gf2KYD0EcNQMwMi+9J4o9hveE0YWKcfwFB55ohT6MrSC35Nmv7IuOi
/U849I37WsYdpxW9UAgHprf8aBqt7bVX8NK/mo9O0m2EHte00AugIk4bU26N2/qb
NEJ3LFhmkyT17ey2X7nV+oWgwnCOXjABct3dGlYYF7bLKAw8IJrararnkVj7VWq+
X8grr7GyuRPNgsXS7MHGF8e2jey9ni0+HSkXCojVBoUBsJ9hS3ImOANRlBDB60Da
SnAGeZ9JYWFF12PxJn80DD2sgHFd0EZRVNnpDAPY3wB+p9zZuW1X4FGFK9wL39Tj
f16723kQOkDJbas9Elyg4nokGhQJafRtpKtQw8CVa6ad1NrajwoP54/W9CTWu0mP
NoOe1hv7L+6JbA8WiIFpBAF4bmiZzTy7q5nVjvkSp635ybVRkV50psZ2W35yzgrl
`protect END_PROTECTED
