`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4HiujJy8CIfVaZHTboAWP6R8oF7973Mqa1iyDkaEpHn8DE//+F/PTVd4IqR638y
5VnwFnWJ5itE0slwIYfTL3VaVymkI+YA3FHoK6Dyz4K8XLnkVOKofQCft8bc8rFP
N6ncVQ9jYTEHjx0UcwEbNlmtaauho4WBy/pODiga+QnyU5UHf+ovIXMFTmuuyK0L
2HyN1S4hL5kdgvtj7P0YTYB1DqSa3OnfVR6PR7CS3Sx50IhONjJA9JF4z6yghqCV
J0c8mx+XRCy65QoKxVHdKujKN1SJFfxFpH4tRQgvaa15OrMOp7eOeUMf2NupMCz9
vLHh7s67QZ+UDl1UdGZ8nyaMXyYfEPEh1JYSPqWNdBdeD52lhXjPFU1ysVdy1YPS
HFCmuI7WPUtoxyoA29ldhHIMPCm37rZ7sAWS4j391Dw0U2G29cLpE6FOhtYsRGXV
ws8L9WG/tprFx+ja7j9TinkQB81y7Su9oD34B5yxLhQ2XxNqP7cx/V4ks4M9xEwz
PpWmqhYrQvS6zNgACLHRyhqHEE5UaUnWm0XpnCwXNqoLNLfxnBwnP+TeV4alDR4b
wlNIceF2RxYuHVocZAbXYWzDg1MSO9ZQghgpCMVJCnnklSpjgBRbQNd49L2l+ZFa
rLqzom53BBXU67UVp1gAil3XKq7S7mVHuNeiUE6qp7GdXt7r2AFWQdq36bxVZ/1V
NC16WCqPVIQ3jhi9KDhUGPYD9yhM0tUQZhLmuJ6vTHh6w8lKSKgOZaDj6aU7eakr
K+6i0W3STW7GGlgP/o5qaUtcACUsSErhL5DWPgB5K+Z4g+W7rnhG2iMA35rfkCbf
PhyZ+z4P9rg54fsKo6wevm/PScJB2jTdVCNtQy5T2H7353zWXbE7jWhGpLU8dn99
hn5254Sii0IE5ZOHjcRP+ViMj2d17sr0tZEHa5skIVTh9DyRXkzdV20qmiWKYaLx
WiARjczqj+KaN/APJJ37Yj/UNKWfaPFec3uGhWtwN9rI9qkwJqppwsHNQ+RZYgL/
OWIRXO3qi3UYDO0TDqTI7MBEgdwl639vX9OOLa78QeABKq7/cShkAl3bJL93JRl6
ym4vGUhBfDRX/qVDaDWW6lNc6LsEunc40gd7cKjXjh4/0++t3/Ypn5bcthNkgdRL
4MpoyPM8DzERdT0IGrnMoN4I43kjW/+W1FczCRQF2z2P1bvD9nDRy22fsScvszUD
iow9SmzRQZvmfdyI3h6eslpdRBi7s/v4+cOAZ8q3Kfl4itheL8DtHodtKpR9otTJ
fWgYWHjh0a/JHMCRI5h88sjXuvi8fFA+GAhTrlbyVt3RcPEh81sEqXMUWA7i3Dlf
Fm6+hcfPJ0FxH8/PatweWUaYTSu4JHcLyfb7CU9OMkfZBa+qqFG3o4dEf7Zo9qrz
7RLAdGnmAiXxtZTbkuQYRxiOGq43UdDg0qa6o8xsOOcZ8sf0AL90YbzCCojg1S1P
WEdu2UulDiQFUiLPvaaUGS5O046XxUrS6cYV5bqKmoJAnS+8nOrmJWurNJzgizLV
mfFk0ZyhS2aLQoDosoBmuFK6ocisc7xjl3HkvheF6L54M6iEk/agbhQwofOJi1u8
l52oLp7epBdVktzyiBi0GaOMuzINHcWvO1mxb4V5QCPgkjKNhmxTgBHnx0r65bSY
tPM076oFw3tysC/tQISTMlnSqTyudKFi6t0MxC9zZSxFPbQCIGyr4Pb+Fqju/g2S
aZWyQZ1N6LW8Ve9kQVR8KUo2hV34p41Uk5mOdRNjxUNe1G5c5khYwl9rrDBoF8Ku
0IpyEfPXCKstAjTIipGaXwt0gV1dAcIfTU9VCSlCPo44Zm0Nc+nP5oxRrrbBxtHk
7SfK3iGBjCUHmkqHMBExhToq70TKe2tEyfnnGdwsdcsBnMznn1jzT59VGdOwcPgC
KxD9uv2BtJkp1aScHI5AeyeUHJrUleUG+n0SvrSSrGKXgPg77koH1CIxMtwaLjBD
pzPKlUOe5WLr0rbQ2d13UIfURrX8lMr7fbI95587DX3a+9DpRGAunZcyAT+8qmS8
FBWZHApZJJoLlgNwtA1wJkUNmj9geYsor7YLPKAPD7lYIu5nb/u2FK8XGCmf4TL0
QLQ4UP9/IZ4Pdu02QWZcGNBNQKxikA7rZx+1mZL2Zud+QXMnTlMT0wpBqyr97rHD
UxrRw3jAqDnuQ66McC6u8XsgDtxulo3EyS7vPvg2OS4skM12C/jI77YBnXVh8gj4
7zD7nxh7M6NIbIS+byisocLclhhBnTcLf0+NbfLax0k0PR2WmTcXZXybrjnkEDNT
4gzWRljvgRVOa0EapXX0AAOTjoX/hhhvczTbxaiaU+WluQLmHuGHct7cOfDOIz+k
Ttv2rG4N5AFxaFGZXfOfiLxjYOwYx5th3yzWDir1FFtvVwHHyrL3SCuJhWIcHm0j
ecYv7jBgUNMLIoWhtbC93FILhxzmAq05CyFSv9807N70Hgdo55Z0zSkZnUO8bFjr
R/r9YmJjSso8TUFHGhpPxNZZeu9pzGnUDuWb/pK58HHZAHJr1JLvOjRh1ihDoU3E
iApAN4Sz06IEuccX/r1JjEBoIhC64f+lMkX1TMegCT6yN+Sum4R5Tnl0q/z4lJhq
lC9NqIGPMkJqFEFT6T4/Ooa6pdZK8FfXljxxuhrvlwb1pqm40QT+sGewpqctGNgr
1nlhA7RP2bGD5RR5tdJwzG9EGIanMP9lFb84FpH/SdR1oZFD3mAkIbaPMGIVFSQb
4gFmlK4tU9CFuqu6gZwk1PsclnJhXaCOQCZg6iIpydf7HOkd/khtCk94Vr8YacYl
3vrChkHwTUK132l4aHvdmjdvUvoCh4BPTU+0Rrf9GbZ1e85UwuC25NsGZ1B803VP
UWTPMF4D5fXCs+7f6oBs5+ucqDKpCFekqpYOdbbgN390Z0mdIzUs4ZcsCLVpO7tH
66KZd7FJiiD7omg1KyZlTnZ8RcS97VV1bFphJycTUx+UswC1QTDD161SNYsNzMWM
JO6zhGussBLNK942J55NGY8B0znkM74KIwry7N9MkQd1dEpkYfCCqKg2Oi0WTFxN
TrDOJfygW3f58B5tg4z11WMCt+0mBhCpEdbzJp1fxD0Z4UNhnQifRQc96zT59tBk
0CNvZxKNRbT09POOW+aDS6NZNWahkdDVrPJRGhn06CalUmFkOg1SLDpKffxYZRUs
DAzR4BFrTuHdRvcIglQabnMBoFEDSmjgXpWhG24+oyD6m58Cuzr5Jhbcx8jIUubk
unNYfZbgg8o/ISj5RCn5bR+cx7PQcu1r/565Ct3yJy5f+1I9lgxON1/zRdDzk7wm
VYLGc/k7G+T+V+ENYF+5fwwRa49pTICkDAGRNRfzz1DhRvhMKRwCYHuq2Gfq0luU
yALHeUwJNG713mEkfUBm9eDu6OsU8QfTwwGTY8tRo0+LQgtuTIHb/+jPeMcqT0iD
HMF3+HCHdkUo2R5Ktvh2g+2ECpYrpUZmoFHvGnOHJjlpK/RtZrRJC9METvakdldG
aYuiMnCmXda5wLFYU6Nb76WdWVspZwszkQeU58QlmHvl2HxCkQ7jnxBRsiN6JHC4
dkBMKrlvwziYw0YSJE+yp+QkfgihQW12WUUZmfksA9oWQw34UdGWMGWi1+yA0jxI
3ZP5avbY3u9jU+HjJjDNPI9uK9SZGuqx7iGKU/PVZHaMNyPd0hIpUkQHo3K/QW5j
M9HACf13NHs7xn7z8arEgjvZ3ADiAj+oxeS+XmNUCi4DHvYx06AW/jFkIhE4sMFB
z5Z01NOSLsbitZee/4+IxG9q2xthIBpPGINa9JxNz6JmcbqVU0l0ECBKTiukCzOp
Abj1vpOMvlHRmQIWYOEXvAY8JlnqExrYuDd+nY23/ySu07crrqumuqfq7mDBHYRg
R9dFvLNibM2PrqbWPrqBbFbOi8n2A9ogSTN7E4+raNRJUPtU7aI9kUYsWASNs8pZ
sbK0ZEUzfq50Hz1mEDvw2m/YtVGiNKS/yZfMPUBYhpIOTrA34bRTjou5g6+Cb3SM
E23J8ze6kh8tDjA/fwU0/19c6brmYQb/g22pVIb0OLGKcXxA9Yfl6uEvNVkuhyN3
8YNKa2xLFAV4uIva/q02ehiVCnwWAb/Ws9afAwQ4wk2t78Dy8x4ntFwB/ZQF1yVQ
wBWtYPwNA6qJq/gCc3Gv+tr7P23g7sFe1SvTExprMZVNOhgK5rYbdKTkJ9G1XV5p
GwscbQuomjVYDsizSqFpT2lwF5x/26Xv25Qzafpo4AwChYKgBF2rJ4aRb+fECIlB
JXBDHDY+N7+3s1E3FMaZbeRsoDMlW+rf+Z9ELjPUM7AGigFE2cXnjIId2i7ibLEy
Ah0rFx+dqryCl7Ic+4fKD4PghksRkG8bRzi1gmfHQv7olkKvymAA2tj1OXwq11IF
UN6ggN4edZJsiB75P4Mf52W6KmMHoZFmUVcvxIUMLz38vgtGPL85JZ06G3wjyxwX
pQyAwp3n8uQyk0AiDBt+aKM4N+6NCWbZwHaLfdXPljWp5A6IDoNiJqdxmbZh8XFJ
v+hwvMTC1bW/RGZdLb/+v8SP1fTTumu0+tt4hN1An6dCu1KPJcmsXU58wG6VAP1j
rzuzljq7ok5ZtMJyg60Y6NBSGmbHniZ37cFR4o8PixxGvn/hgQBdKbSnTsGhlmje
JB/eKYx4IW1VojaGJZthYfVpCSNmqz8SukvSLjEBOrOZsRYBjEvFoo0eggQUYQqL
E5Cy9+T8mc0RymCT3Q+UHhKkZw62pisFp9OYVVvyiYMCcCCakO3eu5/DJq57GWzs
qY1z5KrKqSS24IW3Zy/3XIXOZ3Rugn9EtG5Rnu0jP4dGnj/2/CywMZ5ZGOYs+pDX
4ZyyJ+j1ALO13XNXM4NYEKTYAeMb9wwWykxM9VWTlXB+MRC5/rUHdIU9j5x1Mlw8
azX5bnqxcyx0htDxwC8ZDThVXZys8/FYiHWRBaxJRLU/oT/oncfiMuMQOdD4A09a
b+VQlMQ34Txa3GF+CEAxNlfJ012ATDxp5o7Ew+5sMLeXAxqqDX38A7DiQP8wFirJ
KSSWRIKgn51aOYC8EHEsvuAkLDWvLfc9/HRiP1KQ2zubpk01Fzk5j8jJU+OozhbI
IjE0jEeH52CfuFbG2DTVuAukLDoP7BwMyoYn4DJBs3zQdg91yFs027wF8nLmvmV1
TArX1mQhduktBGdhLO12oJ+AqVv2AdCsbTFJ+7DJOgc8JtnoYgzbZy+YKzK2adxs
loiVDdEBJjwqw8W9tywr5142sMqu6dlGjl1YeIkcaTKhuxbwwtz9ArblhQfQfLtO
rNxI2eaTJqmfp1ehpqgtmKzTSWRxgVwGlfNRSe7soTxM+U3/oxvcNOqGa0NkSRug
iyAY7zOKvlmaULuRA/He6/89zKZ6CGXBWyPO7Pq97woh1ZkrP7oZI5WEcdh7pyhW
CwKIQ78rVcb/H52i/7VqfvHotwBv0YUrc0G5zI3zDLnapbDh72vozgHB1x6MJONA
iVUflWgtdNrms3BT07F2Eo77vjZJBO3FKYIzPPOWVaZBlKRtqTXNIeLdefljoxSU
cW/5XC6iC/16L7K+5e1v6iKcFQaSpWvKufCctuYs+Wd0fKdzxyZ3CU8QuojSLh9N
HwxNjbZ3ibDKJSmuCY0f3C8AWHrOaUPKUV8dtfvNtm+nmR+MsrqFpZbA23wEc2BE
kJnSbh/VI+OzhVKh22NjY3zecsDiKMs93MhVt4syhHuK9Wk+ajBi0NTuPBbeSaNg
NlTQc1j4y7pPx9XdoorDflIukWO8Hee5hPlOXAAvWLhUkalZUfi4/yzjOWEZiAxs
FB+gzJ4qe1uVBaEPhjZ4Z7ybWqFhEav1iqcVc1Vz3IsBpH2HeGXhuNNqfbGEWVoC
2AZl+gOrnVS7w7N2tFDdjuyUSyI/QqznS2bpTfIq/aHLYE2ejMx74f3ksjIGMN0Q
RBN7JDHeGl9JDU1d+zJc1DUde/8dpNQf5t+V6m/g9WUCaPKG5S1Xfpp/4ohhbzIQ
3WIccWyAcDXYnoPjZ3A5mbaE70p7ViYh7vGd6NBGYWtEH4NmEplleL7hMQVadJfm
q5y9ko73MgpCOwak20tb1pCQhLTd3LnyjhTXjTplYhSd8SrdPn+lpPrfy6TPHeyM
Xz0dydIR3f8CukDEmr/Hyiz4wnRXmO8D32MVrB8thBFiPu9K2TT2SF9AY/PDPfPI
vX7yqOQFxkDyIIt9BFzOzff1a6dg1fOzcTKqCm4UrM7RBB7yRqAo1OTVOvvqZit+
FbcNpqa0cD19eaPxBIGD8IcKuD7ttWbPLcz/y0ezQTGRiGYo0aMJ9u4cuA5LsFGp
cvJ4rLcCJOKwsmaGgMVupXbXeySx05r66/4hMvL7VNhDLmiyaHAxgLHTEY7gggBu
IIe642Pf0eRoe3PRJcuO2m+A1+AlFjTFaeq+UPHbpv4R+VgrUThs9FsoE7LkA+yP
ysyS6VfBRFMHKv+R+Rf4EUeBY99MwxSk17aG4ezf4DwkJthzUmSkXDmJctyyjsal
1RW87bHmi6SVg7MWCXcdbhvk+mJacABrQitWN/PjA8tRpTGWOKCjdmMXuzNmv/Z/
c/GjovWEKkDpC0l778ebsGjRGYbo0WL0joAqEMOk2DKm9ofN/95oTODpDct8OqVZ
HublKgJO2cYZRjEx3TVQ8iWI77MUiFSlN8/1YF7cYW+amKRp1Uen+A5bSVDw5b0z
gG0WS2KIzhc23TjnZ1zxnQ==
`protect END_PROTECTED
