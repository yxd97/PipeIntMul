`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oh7Y4M26ysRwAc0ne2an4C3HhCPHgFv82ezBWtZH93HUpzQrYfSA209HYSR/rN+8
4T1rOFLtQcVXbKtExvIuKN7zyUFf1q2kCCAwsPOEGvxvQOsNl/8MoBh5Q3bwWhOP
q/MBZqg7octsGy9MxFqhbcCiXsxb6IILuL6MWOVjjSyhNg0UrmTTZVffIkUZUTIG
1XKAI4xs8CaCxJQBXiAbiBOoDrCr8GlkXE4TBocFkPXeMZaILK8q7cOoDTr0IkPQ
Vu0gUXj5P8vfeeIdSEP3gHp3LAXWHO8R8ePocYoBdS+zULpjZN8JTXuem0oV90QF
tJmkEP7Zuo0Wi8OVv3SNyKFWJBg0tx4LO7RcV4skTdMJs2a52XAWi5MKU9iy5iP6
2+VkEU6LnkjJAcTysr30CtPeRxryLhn/oOkBevF47zEfI2HSjHdD3uxB1ywSYrDW
V+7YehGSLyLOx+eeoP267jiDtt0s7mE4UeGCjOWh3UA1tf/ub6cmsoz2KkFQr8Dd
`protect END_PROTECTED
