`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oSVc1gGo4oipAZMk4LKZghzlzp8uzoF93er3uswxVcrtBHCxOiIA+FwSHXESbLi2
EEA+6ag7U5EgW0MJ7LAmtnrtnPyrb0oTICiidkqJUw+g1c4nVxV3Lz8ga6OHb30F
/+2R991SkOJ+B6Hyt0xpIVWLB2WZYVzYECXO+nuUtYh4kXYU8/Z8XTL8Nd+VcsSQ
WS5HSuwBq5SRTX5rKwSyIXjoS2576hSxQcPmFqSCjlUYLN70PHwTcC6dySCH0+io
XtEXqlFErfk6DU/3sLD8cdC6hcdOKdqd0+PAJmN/5IlOK8tx4YHCsF5+/n0ZXvaJ
dNRQMOSp2pmUUGZol1pTng==
`protect END_PROTECTED
