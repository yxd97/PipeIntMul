`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/lPO5ZeLoN4Oi3Q/vLe9ZB6R5dekkzbFyPGLhOPznXV60E2RYpW1JCg/2OFp2ux0
XHb+B3RI+bFm3uMTcFrqSt8Y1wB681W4k8JzLN4e6SQX8k6Wp6rnszdTJAEpMy9o
l1ju2NOf+MpqFXEZiQW3VY2h8Ezs8Ndc3BwoPmwq2DgUXcZw+g5m9VY/9vy9Noqt
nN5N9oQgO1onC+TOiS3FypDBrpSbUkTfflhoySt8cBA4pXJVSSl/OBNVz4x0t+ku
mGocauI1zeEmmAxL+sfC8f7aOJfqsTei0rezrWfUlL34IAcI3VOivuv2DNftZJh/
jxLHMg8fedRmM6McXvkbcJy3LjrhxpFsmMweTdcUd/GqJ/D5ogpp6KVnwdYWtE7v
pwsttVc4pepbTI6bUDhkEima/agVV2mkcOz5av8Ieuj+BQvI5IvdkcQzFCAd+gCA
wRSBS47UAsZ0o8s5XoNURoUFA0omj8VkZ18TSeuFccGxJr10y7dRJiHuZ4+p2zfA
wFK8TxQ9RWD0q48455OKpaerKyUBH00kJMMjbitfahu9K4GDDX9N+RaFk61L+/qt
nBAdn1D4Sp0NbYuy7FN4YtcC/NtjUYyZ0nPvyyZ3SVlx4un4xRCbsBFcXlZDDGMn
CFHsE8TdEGgLMJysF16mgzdWTuHj61g79jpGp8VA4kS0UHfrye61aMMaefFyq/Wd
hv1IKD/WMivfZxovWEZSH/QYkqcXdt6i6eom51ay7Qs+CzU03KaaTsXDyohhD1op
wasWji1Z2HoBfCGO6i2laFbm46nUiy44HyOTOm0mQqb0VWX/ojdB0aO6pqKUrTay
MAJ7FRQDcpBMaSR9/TknWWmwXfS+sVbxewyw1VfDS6M/5hH5YkkXamNJ2PeBix0q
9Sn7PyMTTtmXU4SqgGEjPGXCjbyou7g6TbUsJ6vNKv4=
`protect END_PROTECTED
