`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFXHi9tBWOdSkLWUmUmLLUB1bE/meHOagpp0fKUPb15S7ucnPhKHq5nHkGiE+JqJ
XjBN4N6xGeYkm/krdCdOmU/hp6NRsGLMkY+z3fWHsrgnGsOlyobAJBm7zEnt8YPl
YQIW4fkqnPFXA4DcBITabEvCIeoRHIWDbJTQMoTJc2kL77XZuYAWs+HuxC13b8SE
bi7u8HZuqFg3zKb/vG/5mjLQobJN/lobJ3LdWLo1x0qsNkOpQgk0kI6ARgq6BAa2
YyVYgb93rvUTEifGBNRTfnJJafn+5EmDmvN4tHihXm2yTZy57yLZuXtgheqaLCj8
eZCDGx+3bW8fHX1OnK3tvqtl6cJlERXhPb3vWC0qq1uLYyr2M72GZ8pVr+YUuef6
qgU3lQioB1aJRS6dH0vKfBc5FEfPDz0KzMFUYizZexBX883AZTLy2r47TAayMbyN
K3viS98CneTVc/uTmmT4jejD3UvKRvEupe/VdMRxBSKCix2gFyPm69W6evTztrE5
aSbcXwlC/zyOJ2tmeo/dv/1UqF9uzSwPq95o4x1UDcWsLyBo85GCPhKLoyYmM+cs
`protect END_PROTECTED
