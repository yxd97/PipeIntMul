`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvOlfOWf2JiKDk3hHXMbpBgv5KOi6Aswe8QlylSAVrK+pT5sK8yZ2JsXgEyDcgno
V41GRUYmKo90y/nmnqIaq+pYepOKGWP7FyvyvJzHlbWr6mRq9s0P25igIe4mvc48
o69y1KNA8SEW6Wo4OrmuG/2eYHtqdtXD1JvZSC6OhNjwjoSfv1igSSaYrgK+zLtP
qDzlUK5KlyRsctmqxYzRJAEu+Gzu/zND/8Qr3OTKe04zXTGg4gbHh5N2ktPftZjQ
hLGrbfGyJdbgf2Wj43s64OEhP9Ji9hJQ1Sd29OrPOMclTAYVBxzOSBn0wX+OxRxQ
BAsJOC04SIrBAACyRUxo6bCFW2W6RreyAhFFopKXP87gLDXiGH/ZankvQpILWkKa
IvZ3KCS6e8vVZ10sqg5G4OowuFxXlWHYHiZI64jY+l3cbZs7QNv7sUr5MvZZiozo
uS7105IIroC2SQZsRZn1sg==
`protect END_PROTECTED
