`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t41H7NeTw5sGfO6iGC0muYS+d/oinXIG7PMJ1Hj4RUiQYNUN63LHPewNiedukgOt
wO6mtcgOIm6ZGSmVfBgrYzjXa/Zm/cdsIeQepy7NKCssWy6Sut17W3svloc9TJ21
t4vGYdI/WxgGGbxHqgWQuZYNHYMqh/oA7Tf9Hv2SJftjjz3uPcXrK4KcbWiXZvxf
e3JZw1QvKyMbz2ncOEf+dsig+zhWCFYcX6zYgC/WLr7tPmommxKgFI+ejufxeWDK
wINgVksjhk0lydD1rk/CRnoK9UawjRxSWC5DlV8XHCtmXvwb0pyF+9GMG7wwYYAh
qdy8ifup2fjBq1VfI+l+d7N+Z2xaqfZMBG4QBCyooqowyrZieX8+xHYO3DysX4uQ
tc2DYaW2GWGYHZ0RqRFXXwHENObC33fT6HxqCqtYSzC9IdMneS1T4CW6MOjvPRZS
YfFmtBn33iszqx/b3wPv408ISybN9JpLxdBilpTTvH3dHntgJIdF7Bez1csCCuH2
+deOAvYM6CdqhN7WJA/zBcz3T1RC4uIr33kV1OKkRXazejgYZ/cvogunwVC6l8vf
ZJVAKZyhpET/AjaTtOSPCCekoVR09xxmhJs/90gy5dqK4lGiHJIQlSV7kiMrjTG3
gtu+RM/Jh0Dw480/C70dFoSnlv7zlaThlL9V7iqqkWat4WWJSnELzwaHgqq2UgGx
SmRiE/+RP+YvHNVCRq/ay2PARS0xmbCnm67nfyReOdxyoAdEvm+b0e7+J+n15xX0
2zJWOW2cTjPC+p7LZEd/khjIVXYaABvuMl5t9BMngflo+p5Q+J64AQFIbzhni2V3
6F+G9HtpWh7qXX7xzxQmKtcNLVp+FeBKm+7nAJB/fXZ0OaZKYESKLZ88mDkDngSs
LmWQ8VldbdG781YoITZfIsijfAmQzZxwccfKK4GZC1cchz3fY4Yr8z06bMfI1nRQ
DDThc03f2sJ6HsE+pibQeKOb37MNZ+B10K+PfXDuRIG6FBa0iQc6UFuFVo4A+OLR
5DdLOypUGJ9b9G6/UT2PvNf10cHWTAYJvKJh0ArcVD+9OJFgwg858sXAHmMgeXTV
YCjcH0lyrbdfqi40NV072LSqj4srJjTGqL6LvNLPJYMC+1WwO+W5hzTGHLG4ZFRL
n1BH975AQu1ZeZ3yRY/V9GdzfS9cRpbuLkkI7RKfA16LqLdbXWQuistOR4vZBYej
MUTNOlJw2uRB+W0SPx4ZLuukqVZyPr/Epj1hqGji4neMQLLCWqurQJ+tf+tmGf12
d72ors+lTAqio5mgYEhqumqE0z3UBWfMjBqM/itiJXveDetinaglvMvxgeFj53kO
qbUzH2rP8k8M0MXClyDS6lFtAS0+3nJwApXDLUhEbOo4C+w31wxhQZ+JMkwEo7x5
6FzEwShfnBLKN+3/M/s4bFmDfpV1aZ26FcEnHCPRtr6rY83O2lwS1jqgBdrqkTZ5
ulVUrEsgi1DPyXnTuzZTN0iFdt+Kqrv2cu8k4rHak7Qz1b5ffL9t5A0rbtKCJ4JC
57c+WWKhI0HFb1RU8lCVjk4s5LiuMluGcuHc9uu88XWsL61/zk1r+EB1N5ds9GDY
g1R1rjvlsmpe4m0fJwJu+UJCrejmT8JwTqISFuilfa1Gt9+hFm9sNG0HRZNE3Vc+
pAEYvM68hxWR5RgFpEHy3ZF2WdOXBTA2hitMYQfdqfJXrhQ9+jKMqRyGjOuBV9pQ
1+nUX5KIks/zerUWwy52IlTHgylGU1gWoMzh36oWSQN0RdIs+yiGopcKz+6BJHR3
5S1QH302PCYMcAEXKWPeIFUBMnQ2JGgiHbXSLLot+E//5MZQU7oQcldxHeXy1Nn8
X7h0Hr56tXbg7VWraH7J1s8gHq8Cn54npwa637kWpP0w12Hpw6m86LiDF7FYaYem
kEoPfU3hX4r0m2tXkMy8+GhoMmtSkU1da7b4dghEctwpf3LtjbIzwm7z/miayYbV
aLqzeqbZegFtw4RjCMqrJ8R3eTRTQWvqYpXcA0RkWUBE6UMrUz7wvft430HANjJP
HXSnVPcpkMsl3iNogy15+LQSnNCJSXTwPZ2LbfVyh0SrTO0hKUpBGIhjdVQ1YJhg
ENVLP0FyuYWz+bHhJx4wnck3nzCs1e+gkUD5KP8uevjUprFbGewzXxYe6m97hUzU
`protect END_PROTECTED
