`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lt1n4upHdi7GLypcZ1VExm6H0mi7uiGJOLcId/5qZNiVfLVeBjgNjcoB/sVnSl9w
xpAEsXzr5pYSdnHkfUw0CNm+negJp+o5jD5aAnJrFlJyRJiaFyQd/gtVOQgq5jy7
+uVC/2qXcOwfiSJOWHW8Bdp/tuhTVvR/hoAhPfw4iGBKV7N3WtkdNLbGNIHBro3i
zWYokPKmbpdJWYKso/MXcAOHcpHxAq4cj1RestpDVmm5K5wB1kijBp0gu6jlW0t2
paynhVj0OQIHI0+6pvw6oUSmYkWIAph50dK9pNAAMMnI1gP4jRhqnY0UtvdqdN/z
5c12y4/hTS8nCYthA08mDHYXKjpXcCgGI2haYV3UiaHQsK0/s8LQ8HsoPMh8JA+K
shIDu9NKWth3+oYXnaSBXnvrfg7Zrw8OZ65Z69r+ApsMp6a7X/6EnIQF37F57UPC
cX/eyJM893qec5ikM37rb1mHnpPhDRzoQPkNVAmsuwi4ZgtDOh4UJR1ImAcDidAh
LUYwpmY/N4r4YPCvNQfZFch4I4rb0brA+Wl31DfycmGWpLnyEfK9Wt3EAnLtTUx1
EcJc2s1HxnNLfUxGQt8o+NUXjw1CRoFot2cr3zFRAJM=
`protect END_PROTECTED
