`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1AO/kFKLa+KTdW4uojvE0QgrsznrE5JBT3OZk0jC5HGZr+omx5ZcH1DmNrv2FQKd
OU4z3X0UcaHghGq11MgIll3ObQp969ja7coAAHdBb6xR6hBJlLyT2UGCjZIp9BgH
cSUAYB8rinRh/nhbfnuTij4oRIM1pmRPRTolWlb/Ur6XRMEY/pdhQbzZT6yqRPRi
zEPERMfWXdNTjvap2d2zsKkg2xA4KYxGX1qZcQnaUlFAIWvos0t1FQlSIMMTanMa
YPaaFpN6YPPgQYmhXPWRYmA4erfQ3mGHUAcd4KnBEdsaBDE0Nqj0CYRcjbRVTzrD
Rk2UsX0l8A79IzhHOrnvPsmZfz4e6AF6yclJ51TJD9J1yH7m4vWjUmN/UOtMNuZi
SfDfs4Nq9qWbhOoTVmgbrOaSx6GyHnQuUV+pbYE2dRXPC5+pgQJ2JDaIE18WsTEM
ZWWMpWfAAvPCFiL6ReuYtA==
`protect END_PROTECTED
