`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iRE4uQPS0J51qq5lHZtG/lHpNXW7w7VlSIDoWps1F/Rx9Tdq4DrZdrO2W8dT3yUF
FtmFbuo0oBuU68A+d/L85oXLqWCvLtCCQ6XprHMrn5P0PSCg55nQCnYyh51WBpmc
T2SCCsKQAJuDPC9fVdHOUTSZms6C3Ek/ZTV6wnoTFFj9Q0Y1LjQwnqgt1GA0Lk47
SQ4GnHSVLiooXSivSvwVKmtG7Fg6qnL7fD74jSLNegdE85aTaBNZ1FNmbD/0Cyld
gn8DundECsX7He4tcaS232jo2t+iR5Yc/3DEiwyYUMtq/PJmdlGaPwl9zcrZfNOb
+ZoyqvT7qevh0ej7YA4tLQ==
`protect END_PROTECTED
