`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/OM+zrcT0MGQuPhwN2C11zMIUYsp8UFQDEBqOCUUM6562Z6cuSQl1Lb/Riw7qrB
rbwZaJz1e2B2ZT9IhxrLKIYtBNrpEfmFTz8DbgMKnHbFcsGTNA906EtFYWHD3jR+
ADuOZaSB6WJMNB7EJTgsnjMpSCdHPXuQLm+MyNnmOOIbrLYjwAUSq7RPBPDqsR//
Gjz4NcHgcFIl5++Y1ct9Ckw6vKDbh13EMepdDK9opr32NDrmoMD+uIwzKbOLNFNw
ao0RaU1j1XcgzJlmsI2yazTH2ZS6k05nT1gIXtOhexjNiTJiKP1gp1XLS8oxcGYK
xTu5s6NetTu28RSD5iw7+lnLpHV0AmlntYZWzoov6d7/yrZ94PpEPo29o7U+yMHJ
3m0pJgSlRKnd6FPuaJ6sXiBIbRc2Klw5kAJCE/JjNEUlFrEPs6dTslrQcVhXlYGb
wIXkud5GV+jbjmvhqYvwb68uBsrw6DB804x54OdvjZvZpCSM5iV6X+4KX2JvdfRb
rgRyCIznhY2IZB55V3yh1ulF8t7uOoBWHDik45OuZ9T5jTyKCP2fhuvOtHrflOFC
fjHsroMpOwkC1ixjEv0awNOxovGWzLffXlYZ0SNU7Pw=
`protect END_PROTECTED
