`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X12e5F/d+/zkNMQmGIi5Fb5H8zYeb7zKQ2N7K1KUPUhGtZhxneU+86W94T9AgGPP
2mVc4T0i7sUhCH1d7VjF98ZoJv85xmpKejiXKJSJS9jdZfG/I2tdOklBhFqlK+sd
G780BzCs7mNVouNUPZUscJ08E3Kra39ENUBbm/vyKzHDmisTm73rXVnpBwEU2U0n
TKVdWyiOGa5JMz2OoaxJ/uVfDLAq1lH6JkAc7NVqCrdKtEBlUaR4bdH35ATSEggI
7DnqinTujICBM7xrCKHbq1vNfnUbNWKWuRT11FEZ1dpC5PPUkElc+OMyPalT7fkU
rbJG6uEc0GZoJPMg1GEjCqxKSXosttityCau4+c784XCP2e95gBHq6T3shIDxAYA
S4AAcB8VijR80lvIKNOxgEc1pPlH9Fz8n9ENBFYqfXUXcVIU3U4rSNCmU/05tROf
mijvf25VP5zPFmep8WSLjKnOu8ZkS+PJQAHhNWQ/w0l9aGheQWtBh1QJjaCHA1N3
FqEE8jK0uTrIlLkoHVVbYGH3mCVdpEXD1waBh4cGem59sQVvoTDiLPmX5HjDKvkD
403jRpp/ffhkVout0Zdqk3P+JIUZ+/6If3kUkn4QFxWfnEF+ARopXD14LDxV1EmI
stf4pTOSD6ceWSoEGmiIpGolALGa1fkOyKnVNBFTyYlko1JMy+Glx7zOJXR3nhDO
rCLF9l/rms5UfMApujvlx7NFjpzQT4I98q8ykkBO6SLMbEy+uNgHg68WEwtFwISc
qjTJcsJwiTbmifSu5fHigWCwFBlwZXF8HlVyFuaQkoQtGeMY4Evj4aRrcjaWhI4Z
Ycs2ShIpJyvpt+mHOKCgPXFa5DXxed1Nn4J0z5sZiMrWgJh6obwICS6c/81E2mQy
RI7/E4SvhgckaA+H8QRiSIf99iaZCFNtT0mL7cf8gg7zl4cLTnVqSUtffRVR3TTL
aQ+Aa8aMje7XhVJw1JAYahAWL7sFb04mXqeYiydhCGpTCmiIfIeLUUr1l3gZCnUB
4Y39Q7iv8kFSK1q5q++rn0va46kZqc1R7zoOI9IG0iRbPnyw+TBLZ2ogjRo6a879
IaW1NqGjwxITWOYmqQK+jqbscfRu0d2RuMW1yGobjx9JXtuEBTkHTXEpQv7KDrio
VukFiU24HeSqrjZ5m9qRDGF49XxtVdNNsAhzgGsMTr/OZ34Gf6rtUi+oEY+sjPc1
pJe8jezRFhi9q2zvse/1LFccCLGgdEasN9jaqw49ZuI4RRQRi7pd+wQp2w4ZkZLN
olggeEYMVSsnw4GkWtgG37XedO474P6kX83pbEmml4dvP6X4lmrpCakomkbNQNHh
l5YUlFOjM5CnVb5GDK/KKhzkLacyFdWC+IIJe7xcPg4m2JiSJBeFIQJvTIL4KsPK
N2PPWQ43mKh2AL/DNPzjMfrNjYQKEF4qBAgyZ3nUoFAyy6HftXqGckLadWW6hIQW
WunHKbUrOvek0eXkcvO1udIik8WlrMrk9nToorm08VL/PntvtYmVDA2K+6tabsQt
nQFCMAkhyxpTA81prO44f/8MJTey8+Zf/bUDwDLG21yQLt4uDUPODlDdnQ+cbi91
vvar/bb67f+/6hPZ1H5pgHzPAWrDZ9HRh/xa8hJT2Y5OVWwA355wNutpWsaavN7T
HhTobHyqen2xi3890nCd4+B3M71NY6OXyrrl9q4ZeSt3ZV5qN7dWN74Il6KbsHel
6eG2Lv05e9KwZx+4i1bDQBr3dIJIguwe/kUynsjnPlXcGj6xC5OVX5Dp776VzuLu
FunSzK/76lCMMEMRrQ5DJHm70U9/JkzyxNcA5HAQ3koAH8PA9cEi65a+3dvCgWlx
OMN1b+Bwlx0deWxUqZJTX51lTYpqUvJTZmyThlcqKkXOMFQWuN7DmtCD9Ta8E1dH
KgEJAiZltWJVq3TK+pulwU5pS4ojE18NOQMiQCxXGat9uMZ8qHdpz9XaZmhtkMGN
NhbPYlXnwpWEiYJTeCNx/I6CeS+6AXU0+nVx7xLlQ97fJK1M/dTTf1fOcC/RY3pJ
FDEI1AOOGM6BjI+MZaBajZCZNWK/u/pgbyHtcH8yev8HVbAvBYu1yhGbz7bEf5+o
qIuW6Znc0pbwI+UUcKW8sZM1uQqvhE66RSoX33h14yjXroLjomq4gR8QWwqLWSmX
xi0VpOvBju+yDoBJk5vmIRdddGevRTmKbGBMIqoRPma3mqMBOfplJmioOco0BgVX
Dc9jic64jAwkjW+iTt8Rk9IgX/AhpUyghdQsAiMvUJYFjdKRyHwdx6+E1n1T0sgZ
pP+HknO0Vs3FY/oHFBItNI5NrtiS7kSZlTApQfJAGciuO96J2EMwxROdfOier9PR
uP7i4J37oiJRdUNaLer4c3C0CvWYCS+PdO4f3AYgVaEPoYbFnfqthSOs453zgkBh
KI4mj40Jjbv3pryYyIq9SoWDXV492yt8Xb4YHEnQnb3i5gHEF0vQRkyGrOTWp3h0
gEnkyrdMi4Vr/JAH6GDuDZQToRPVcBrLpZ37uOMS4z85OtElNGIRbJee0CXXdfhu
s02drOy/gMOZQfdkFeNOZRieNUfTBhdtyCZK/gS/lnUtDGGQhHjZLOHAK76TlOex
jfU0Te80ujzUbkaOHROfNGmXADZFt27QVFUL4rG+MuXggZDkV3bIPFaufh0smnD6
TAfZXn0GKOBgrEJYAZAkU/wJHmYfB4ef/rab3gZeCl7xPWdcYwWsQXtuJy6Pq5GV
NlPkoPJhSwXz3hKZ9n7plSGvdDoB/6tBYj8yct2alYOSfUZaNaJVORcXISPnAIoG
p1vwMOKd7t9NlFRiEpr1HoUxNeLbvMYnMrNtGmOHZrnRlBoH6hWDfG9nn9dtkRI8
7csYSEhZ6C0NDoWHWmm96A6GZy2AP7RN0hVQq5pL1k8+gXabNjMLLY29dH2tfhBM
0d4RKaiWRHlYjWh/0GB+KSmSPsY/Ai2bp0zsezJWTONcncWddEeaeyqCTGT+mOBI
tK4o2FsPuxg2PP7PfwTrL9X9GGwX+FF4Ij5HfMY84/0pvprQkLllRGLzq9YcSf7i
R8kpq4ac33H0edB4ryRsnBcYBL6R+V+fBliRhNtuQLBh8wIF6rbDQW2HRSlfb6o2
DH0iBYdrw/hCcdxzK7LPjLzVjS87hYSSAaztJO3AX9VhQsfjwrKI7MUhHucBg7f+
RPGy3uS2tJPag0F7lWP3KWEvTd/TIqLqYrlAFIxnWcYieZhCL0UHJO3nPJryPtAQ
7DHmGHaquTRxP40GmCQYr2k1/49n6vseIIf4Fz8WF5attWIGIhmEZioP5e7mSm/A
K9GxxdMXChiPQgdJD/BhYxt46WkDV/BIHMMjcBXYk3Y0cQ0XyJ0U4E9x5CC6nbV1
rt6VRXTkAXpuAsSgGduGuX9PAnDeJuHouKI2dthB6jxHAczKAt1rjbXC3Ita5D87
z25ABTZ+Yp72YwsoZClti+6U72Kan2qrhUkkDjxr5W/2SPfjPjJEiJ9Jk4mwmWyY
H1ai/Dnj60BT9VT5rdh1NpDWojn6O+6UVKL2kS0x9HMGjhf9+2VGl6vnEw7vCMDB
ZS7Mb+H0TxSGFMW+ni1q6W+jboa4o6tfKBFhPsH+6TETkZGTJLnVkteSoSf/RrXV
j4TC1/v7Jrx+o1ivdnw95ARGlMZqcQVWDinh7x4h0cqwnp4UDd6SZrb5uy4oAwhP
zGOflooe3xF0EqHlGtw4483VMG2skxgDj+Bypa0oxsQ0H/OaxtuD5+dIxDgZHLAo
`protect END_PROTECTED
