`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
danJJyXM+FL6BI0bDaJBZ+M7O/VKj5sMF8L3bfWFYrs7eTEjeQnGLptuF0dIvxOm
CSfgXovgVW4kG2sRGU6vPJvBSSeRzuLIgTsWxOCf0vSShq++e1cPiWz6/AblUWK7
Mks//4mr4m+8ZVJ8LGNY/MD2tdVIX7zgLYZqHsx9fU9z8CV/ZLkfU4quX5lnGmck
+XO4P5X5L9l0U8a+gP3AtdVH3VLeUHagDDp0uzluN51vAtJjAyAHnUcysGCWYg6x
t+uM2bUKqjWcORo8SlU9iix/4xwiHjJIifWzvycj/cOqV3vW7kjn+bzKTUHDO9lp
xCLDiJzmwUW+fhorio9BYAUIsHY7aXyutF4/h7dcANlwSCAWNGscILwsvjQjItok
c7Of+NSaCmp4G/gU0FBnUSz0Tnpds5AzEa+JROxwRZoHdnkkKSvsJBIzz6fMREej
PBxS+nJ4thbj5Z7ElR8BGjTWLojNw2loRZe4ZAnTn9KBpbb53OYkDHRLr7ONtpZ7
4d/Cz9Nh3Rw4jg7u4OtDo8xSJr82RxzRGi3I/RjvF6+MhSSH+YWkKt/1e6apKOHw
bJv8m+ixtqPOLVWehW+yP4ykE0D0pT1ThKjQXqdDasb1MaTFNzkPmJBpGt6lr4el
g5FgmjZgQ2MEG2Dn0XHQb5Rt307vKwO4wgcwhcni+xhcv9bRHGzZ5QCA2sDqt2Rf
uoRmmjkL3sKzykXifEDBS4HLADshZI8Eubp51rjUxDkAadSsyl/biyWZJNLVVzln
p4sXSpljCsBU7gdKlOywo1/9CAnb9Isvyy72jcTWZzEQbqX8936ikhe0wSaSFnqv
QbBTDPdR2QmWGwPowTaMhbeQNrhE/fhWABUnWFWxQKwmcBaP/gZaMsX4/LLlsuaC
4D6j1mdSWCWhYjnmacow0O2bJ+MJt7vlqvWHwRXKk7v9MvVJ7xoOIToeNguoWe8O
zswWAwCkixj3kFCyoZCtAAKK9RJhSxGku4QDDUPu74y2BFaWCKJqZctowblq4D77
OCq9QarTyVS4skCgDwA7h1giTs1IOOzH13NeNO95+zne+COHzDCDKTX6yJXzAV8V
TVtxhU3EMyChnIKnDznf/KHL+MPByEy5bhryAjD7CUDXQi5UyobhEF4pYSzpu98e
dl2tfsxvzSaWXMFlE4TEDirjY27PTyT0FTNU9DKKO1K90Y3T1pRD2yjJueRXFCm8
7B+UkEkdS4DNiSQ6Ki7v/r2g9zwf7tLDZnm9KVw0io+Kzb1xs1QcYzI3eXiF4Tdq
Oc+QlaPZEwdRoHNeYOayd3CK2E9r0daFAEKndV6NQF4BFJLp1GiNMobacUW5S6Va
tmE/JF246P4VWd3LHldHSVySq+8UUyAJuchfcTHDg9WVrUXLuX9plfwdqmX2y0Fk
thoVA0bPy7WFSJrfUwKrrUvPdy4jw958wNFwVj95hsBfgxVZNvVyIyG9e2XNkh38
8TRDvw9uq91ZAAfjoVAcgWJ2FSIekoWwlpTTRAVUNHaWwsYRUzQ0ve91ReacIt7M
6jRohPEWSoluEBTe8Xg3VIRLx/jpo/Tcl7IbqE0XmWaZHiZWdJIQSvrPU2diJ7bK
S8Vsrqm7PB0YHy5Fz1vXP71PrnxY2j9UtSCuHlaTyv+4tAo27H7otxqTNQJ9b3uj
obucM7iCJj7dk5eYy5RjcgIJLTHJg+ILJUEd3mcy/Yx9X8IGy+C9Frz2YJ5B0gTs
UTmbCDRghq5OcaBTg7szfuX8gOw6Iy1iVJMkMUemIEsdjiRDf/i1/9KE9djY0v1u
crurcGXyNDkc3NBCZlaOIF1FzAea2MMYpQQlcYho9r1iCQZIoCtWuUUqqqhYmfKi
ppNEd4WvHCPe+M14+V1eHSri4pnlFFqO5LQQD/rJKN9NCvyXEiLxRjijkHSHqk+H
u2pEf6t+YepmH2deXec6lW1pqKlvEPirnUjw7ZcVMm/xTVtcFxyH9DO1EsY5abbf
m/RCKUPf6ykLpD/xXwsWRg2URRJzVnOVlt9Oj6wLC9JzRf5VbPYzolotuwS2gzM0
/B9nf4KmJg4agiy1OSurl/tY6StKOU0EgmFSH84W5MT6Wn3iv9mW5mc8k8FYfNyo
NMx8T4hXfawQ9Uw8nMCK64L09e9GUXIpgRgTU+iiuKX5W8+4ROf3grvye0d/o0Kh
KJkgnC1BQi2JdQ8fpsR0rfsb/2xqlBKxRdkst1a3FUhoU9zPNjzjWsXF7Uy2gN3N
oIYgF2JqcpTMqQiRRGAy2SQl7dU3ZBQb5PSzMs+9DPeS9KYzyBQjeVlCo/91Rjj0
TM1ZUbgcTINrafM0cCvQo9M46sYAA4LxnxLarptHKCmyoghnLGicNmCL+hTwjVCI
cm2PWvrQ3IVQSXWE/GzT4+D2JfTwoIe9c3b+AJ3p6IR+T7mSv73OgsYiKr2/ByDX
Ra+3QQGTwwrEc25bY7fgJ20ZkALuBrys8ChomsDeDnI20LA1o208CUi2WTXb136g
z55P+OtxC8o8jaawRFySf79joDTqvfpycuibERUNfJC/xl+nrqb3tfqaCLgB3d/d
UcEGSU5N7UDDVmnUGrKpv5UzvYzh2f9+MO+EPsQDw3mZb0RKIOtoJLvMBXIO15S0
VhPc/b8rNyZ5vFhdScYLjqjPhBpH6RfCxFngOBXTRZnWckNldjBRMUmtttuiIgTB
HwTYvuuFvKh9HBrHi/77ewPp113iHGl5DtRoK3i0KCdrMQeS9tozyl3O5HzWiYbV
A7mPs9syLKot9i9qnLkgwFrMBcHLzT+xz2j8HjGFIpkj0lEiSFus2pq7TqVi2zHL
uzebhcBJMBwz0T5Wcg8dQbywAFtqbnvWesV3KE+FIwqBl8x3bUGu5R4FUKBvPdu+
gciYgRiSAPvddtf6ZpzhkYK+eHIFr4ds9uolYOQ6fFb4ezUrTqyD86upYG92BQua
xzmWEKfh+/J5tPHOotubBOuFnq9Ce0cpokfpcACCpfPfd6Ng0ceQlD2zsBFCaKhi
bxIjKRYVbeERz7xxQCkJ0Nc6b6hYUFJ8Zdc66V+lCmdMMhJw9A/cWc4ruq+ozNib
U1+bmhodq0apwDxV2gkdlBWwvETC1q3XqcTwdyAU30p+UiExb/U/wRgeoBUmiOe7
q6XtbkoMDyzoY6CG2tO/Aq2Pg5tbZcUSf/tKCgYKQE6VRNA8J8fl9qkoaA+ORs/+
QxPC0vuQz19cSYhGPNb95LxfU2yvQnEEFgSvz0bR0lM2jLZr+eybEw3n4J9bNg8o
oPU40mAJGjqUaj+rEFHFTNTJ/eUl96Cs+uJoOzM0poE+tUtglfGllZDfQa2rhga7
AZQdl4vRZ5hy8upNtANoUr72YA+CsXGthP6WuhEoCIvnYG29va55fYo82gyIkl7F
bd4OXwzsJCdoBYbbK7Rs9k69I2uXFNN7tgQaXWMd/ee+gm0jGULk1E0h9An7pia5
MjIyAVqSTNqWNl9xAeUBsPexOBQ0/xXCa6TRgYHW31WrGCfXn3mSwIluYyjoy6+e
QYD/htIBzFFRgCSutDpvnX8dv93DWghyYeeaq596GH+DdO6RAf3WF8F7ecp2QLKb
1ZS94bLiGXSGCSScDRegHXswMrEJZk3FFe7X4iNbn7HZPEkrMwfts1sFJQBqlsrs
xnwOyzazboIxXkSkY8oW97Wm2jhi4eL1UKfQoOSaOFPGv9my2bFX1j0xjad+lXZQ
CskQGsLmGLQDoTuwThQXJs5asR5HZH+N7L0cE8gZfF/vUcOhARBWdryoP4qSY8Wx
57zq5dPT81raNEvruSjvoNp2TNxqYMHZZn6cXaS77/XXPRZR6wyePe0sfJBDC8w9
2XIM1SfHf0yiA99txviE3KbxgzktcihQJcb+Wxh25fZFruoDHEoTrpmZRu8lRmXw
vQMFo5t0EsDZWjwFF4fTqJz0+yEnZq3F6sp/+OFF8YR4Gx1RsU+NXi/IwJnSvK3e
xvopT5Ru7lOb+bhwqBi/orLkoEKSt3eAG/YE0wNO8VS239TJ70BPL1uAyiHaw0yo
`protect END_PROTECTED
