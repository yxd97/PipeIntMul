`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ODZ0mS+AOQutyrb5Q0Dh21A/Qh+qW3EvE3XWT5Eunf5x/TK7jmThfLJwviHuiw7f
ntyYpuCfat5vCYAgx7wYScqvwWzNN28MhGC+OrYYC6IpXO3dCvw9SxdeyG/OXQha
sAD2TUFNBfiLf43CvOHgFNOiw8DcCaOHKN4WUbl6ElvKTBhgJEGdGfy7WhDv4BYd
wTLng8KNpIngsA63Vb+GuZXbK1LzymyoXb5m4vZ+t1vaNPNjzCHm/SC/ggoj3gq3
0p3h/GFlErvnnR+MNVtPwDNZVRYe8NO9xmw02mrzpBuDmRRhEuTRMS8BEeaWfPTD
W4fkwOfKC0wvaiIcL5P2Jk0yhH3yLy+6RSjnM+wPARzWDWCGm7JqeSVijLKOXwI4
s9qDctOuM1YJS7e6YwZS0jE3/I7xjMtWIp94FLe/FOIewaI87aOS/Rrefu3yvasT
c388E7VQ4LwTtwyI7WilNX6Bc5lYPHYXV3oYSPSkvFY=
`protect END_PROTECTED
