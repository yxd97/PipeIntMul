`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p3BeSAJBkpgsPtAn3ZQUlQPT6rLHdQSt0wn+fR3kJrFBSkZkKK17gyOV2FTecyrf
Kks4d50mm08rUhysNwa+MVxmn6ayS+OeIA6arz/DigFpuGWefewl4763h76ndhZe
5lKSxehr7ciWr301trT1EReA4xBZFK2l6ekt0bg6q+VnUGFtVUOc27POrz8/dBsG
N2AW6lad3Vwkhzt+J/LLEHlylSPVEmDJ4zl/wuHyFW7vsAglFUq+6kKN7wiiR0A6
NJRYIlFdPQOrU6w2CpfUFQbeHRnTDZGJ1xB+dzTVk70xlpZI9wM5KN2nFkD9n5dI
v+xPKEQECc1Qb42jHUALXw97TQ0TONF5+CiAyc9qHV+EaiLT7fcfF+Z9zTIaNPNX
VTt+C3QInPRA6Qd8h7+y7q0zE4v60FIPzeW8GX5LnT4=
`protect END_PROTECTED
