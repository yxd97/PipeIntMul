`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfrmJcI7lYx5TUiHH8DNyWvlb5ZT1l8uukhbDr2u49kvd4LU59vEgGry1002m22d
Y6/UV8/ZQh21dGUjl7eaxqrNP0T2T0siYNkI8+Polv7rwgR7oN2XNE8e2nXmN1Cq
10TIMKcgfhkcq46whVXLRV6gAcLuagSsb2Ue4o1Q1HXcaX0nj1xXKL/rI05KMkpG
/D/E7lDH11oBtg2to4bVBa5bhZK312TMXqh2qWhQ0lzjItnu2nsKKtX5xQMqh6y2
ZRKtEw5S/Bg2dxVpbTlOlyiG0Fb67L3qkk7CMdQ5uHpk/EVCyHvlTX9eYm8JNr0w
SrW8RYLknQXEMP/hNcOlZ25WMNjR5Sck0K9GC4UG6wTxOvcMi5MAc1vXzPio/ehC
`protect END_PROTECTED
