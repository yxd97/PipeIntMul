`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w8Ugq4wH/b58asbMIAVUs/Ig1+4KcNce4Jv8UjJazqa3se1NfNpE8XMl46liND+f
j+HoDJXFtO/DGWRPkyEaYdpZDBuKsNJCJ9eFelyImRwP0nhJc+fLc4OEUdCAJ/6u
QeUdKpA8RpX7Wi1ZeVDkptZ39Omzf7spRMAUK6vn7Lf/l5xkXYjprT76LqjtcOtb
TOwNB+K89+yWlnJumaBG230il5Gkop8KsCqmlRVy+M16xUewFKV9RuPuokWR6Wgt
`protect END_PROTECTED
