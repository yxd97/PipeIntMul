`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ptyIPG9onpnDGNyff+dU+palZQ1JzNoE517pdgLMOYyNGhIEkatpQaxjkBP3SIE
nEav7UAyHrbSqAJmHUI/MIBBUuSmFkuLSpQHWkSe4hmVTcrijE3dIsfWMc9eY6Yx
13wpdndbSOIbas0v8xuxZ2B1QAm8MpFRqzjZ034YY8k8BoMxbUYUb3xs6unnOxqn
3pNlR0mv+DhuKMJc/G40WQT5p8CbTgxu7A9Wue4ok4oGc2yKAVOdjU2mbXUhK21b
n6zD6Ei/C7KNtdxwT4/zgejz20WG0GrG6f1HeEyFWW4BMaze11dVrkzXIBNcvXz4
3I1pYoNcfIoV7ksCvlXWLkF/Qx2wm/Vk3g1dgfPkCFaSmkJdFzc0wFqtZHuCQU6H
`protect END_PROTECTED
