library verilog;
use verilog.vl_types.all;
entity X_PS7 is
    generic(
        LOC             : string  := "UNPLACED"
    );
    port(
        DMA0DATYPE      : out    vl_logic_vector(1 downto 0);
        DMA0DAVALID     : out    vl_logic;
        DMA0DRREADY     : out    vl_logic;
        DMA0RSTN        : out    vl_logic;
        DMA1DATYPE      : out    vl_logic_vector(1 downto 0);
        DMA1DAVALID     : out    vl_logic;
        DMA1DRREADY     : out    vl_logic;
        DMA1RSTN        : out    vl_logic;
        DMA2DATYPE      : out    vl_logic_vector(1 downto 0);
        DMA2DAVALID     : out    vl_logic;
        DMA2DRREADY     : out    vl_logic;
        DMA2RSTN        : out    vl_logic;
        DMA3DATYPE      : out    vl_logic_vector(1 downto 0);
        DMA3DAVALID     : out    vl_logic;
        DMA3DRREADY     : out    vl_logic;
        DMA3RSTN        : out    vl_logic;
        EMIOCAN0PHYTX   : out    vl_logic;
        EMIOCAN1PHYTX   : out    vl_logic;
        EMIOENET0GMIITXD: out    vl_logic_vector(7 downto 0);
        EMIOENET0GMIITXEN: out    vl_logic;
        EMIOENET0GMIITXER: out    vl_logic;
        EMIOENET0MDIOMDC: out    vl_logic;
        EMIOENET0MDIOO  : out    vl_logic;
        EMIOENET0MDIOTN : out    vl_logic;
        EMIOENET0PTPDELAYREQRX: out    vl_logic;
        EMIOENET0PTPDELAYREQTX: out    vl_logic;
        EMIOENET0PTPPDELAYREQRX: out    vl_logic;
        EMIOENET0PTPPDELAYREQTX: out    vl_logic;
        EMIOENET0PTPPDELAYRESPRX: out    vl_logic;
        EMIOENET0PTPPDELAYRESPTX: out    vl_logic;
        EMIOENET0PTPSYNCFRAMERX: out    vl_logic;
        EMIOENET0PTPSYNCFRAMETX: out    vl_logic;
        EMIOENET0SOFRX  : out    vl_logic;
        EMIOENET0SOFTX  : out    vl_logic;
        EMIOENET1GMIITXD: out    vl_logic_vector(7 downto 0);
        EMIOENET1GMIITXEN: out    vl_logic;
        EMIOENET1GMIITXER: out    vl_logic;
        EMIOENET1MDIOMDC: out    vl_logic;
        EMIOENET1MDIOO  : out    vl_logic;
        EMIOENET1MDIOTN : out    vl_logic;
        EMIOENET1PTPDELAYREQRX: out    vl_logic;
        EMIOENET1PTPDELAYREQTX: out    vl_logic;
        EMIOENET1PTPPDELAYREQRX: out    vl_logic;
        EMIOENET1PTPPDELAYREQTX: out    vl_logic;
        EMIOENET1PTPPDELAYRESPRX: out    vl_logic;
        EMIOENET1PTPPDELAYRESPTX: out    vl_logic;
        EMIOENET1PTPSYNCFRAMERX: out    vl_logic;
        EMIOENET1PTPSYNCFRAMETX: out    vl_logic;
        EMIOENET1SOFRX  : out    vl_logic;
        EMIOENET1SOFTX  : out    vl_logic;
        EMIOGPIOO       : out    vl_logic_vector(63 downto 0);
        EMIOGPIOTN      : out    vl_logic_vector(63 downto 0);
        EMIOI2C0SCLO    : out    vl_logic;
        EMIOI2C0SCLTN   : out    vl_logic;
        EMIOI2C0SDAO    : out    vl_logic;
        EMIOI2C0SDATN   : out    vl_logic;
        EMIOI2C1SCLO    : out    vl_logic;
        EMIOI2C1SCLTN   : out    vl_logic;
        EMIOI2C1SDAO    : out    vl_logic;
        EMIOI2C1SDATN   : out    vl_logic;
        EMIOPJTAGTDO    : out    vl_logic;
        EMIOPJTAGTDTN   : out    vl_logic;
        EMIOSDIO0BUSPOW : out    vl_logic;
        EMIOSDIO0BUSVOLT: out    vl_logic_vector(2 downto 0);
        EMIOSDIO0CLK    : out    vl_logic;
        EMIOSDIO0CMDO   : out    vl_logic;
        EMIOSDIO0CMDTN  : out    vl_logic;
        EMIOSDIO0DATAO  : out    vl_logic_vector(3 downto 0);
        EMIOSDIO0DATATN : out    vl_logic_vector(3 downto 0);
        EMIOSDIO0LED    : out    vl_logic;
        EMIOSDIO1BUSPOW : out    vl_logic;
        EMIOSDIO1BUSVOLT: out    vl_logic_vector(2 downto 0);
        EMIOSDIO1CLK    : out    vl_logic;
        EMIOSDIO1CMDO   : out    vl_logic;
        EMIOSDIO1CMDTN  : out    vl_logic;
        EMIOSDIO1DATAO  : out    vl_logic_vector(3 downto 0);
        EMIOSDIO1DATATN : out    vl_logic_vector(3 downto 0);
        EMIOSDIO1LED    : out    vl_logic;
        EMIOSPI0MO      : out    vl_logic;
        EMIOSPI0MOTN    : out    vl_logic;
        EMIOSPI0SCLKO   : out    vl_logic;
        EMIOSPI0SCLKTN  : out    vl_logic;
        EMIOSPI0SO      : out    vl_logic;
        EMIOSPI0SSNTN   : out    vl_logic;
        EMIOSPI0SSON    : out    vl_logic_vector(2 downto 0);
        EMIOSPI0STN     : out    vl_logic;
        EMIOSPI1MO      : out    vl_logic;
        EMIOSPI1MOTN    : out    vl_logic;
        EMIOSPI1SCLKO   : out    vl_logic;
        EMIOSPI1SCLKTN  : out    vl_logic;
        EMIOSPI1SO      : out    vl_logic;
        EMIOSPI1SSNTN   : out    vl_logic;
        EMIOSPI1SSON    : out    vl_logic_vector(2 downto 0);
        EMIOSPI1STN     : out    vl_logic;
        EMIOTRACECTL    : out    vl_logic;
        EMIOTRACEDATA   : out    vl_logic_vector(31 downto 0);
        EMIOTTC0WAVEO   : out    vl_logic_vector(2 downto 0);
        EMIOTTC1WAVEO   : out    vl_logic_vector(2 downto 0);
        EMIOUART0DTRN   : out    vl_logic;
        EMIOUART0RTSN   : out    vl_logic;
        EMIOUART0TX     : out    vl_logic;
        EMIOUART1DTRN   : out    vl_logic;
        EMIOUART1RTSN   : out    vl_logic;
        EMIOUART1TX     : out    vl_logic;
        EMIOUSB0PORTINDCTL: out    vl_logic_vector(1 downto 0);
        EMIOUSB0VBUSPWRSELECT: out    vl_logic;
        EMIOUSB1PORTINDCTL: out    vl_logic_vector(1 downto 0);
        EMIOUSB1VBUSPWRSELECT: out    vl_logic;
        EMIOWDTRSTO     : out    vl_logic;
        EVENTEVENTO     : out    vl_logic;
        EVENTSTANDBYWFE : out    vl_logic_vector(1 downto 0);
        EVENTSTANDBYWFI : out    vl_logic_vector(1 downto 0);
        FCLKCLK         : out    vl_logic_vector(3 downto 0);
        FCLKRESETN      : out    vl_logic_vector(3 downto 0);
        FTMTF2PTRIGACK  : out    vl_logic_vector(3 downto 0);
        FTMTP2FDEBUG    : out    vl_logic_vector(31 downto 0);
        FTMTP2FTRIG     : out    vl_logic_vector(3 downto 0);
        IRQP2F          : out    vl_logic_vector(28 downto 0);
        MAXIGP0ARADDR   : out    vl_logic_vector(31 downto 0);
        MAXIGP0ARBURST  : out    vl_logic_vector(1 downto 0);
        MAXIGP0ARCACHE  : out    vl_logic_vector(3 downto 0);
        MAXIGP0ARESETN  : out    vl_logic;
        MAXIGP0ARID     : out    vl_logic_vector(11 downto 0);
        MAXIGP0ARLEN    : out    vl_logic_vector(3 downto 0);
        MAXIGP0ARLOCK   : out    vl_logic_vector(1 downto 0);
        MAXIGP0ARPROT   : out    vl_logic_vector(2 downto 0);
        MAXIGP0ARQOS    : out    vl_logic_vector(3 downto 0);
        MAXIGP0ARSIZE   : out    vl_logic_vector(1 downto 0);
        MAXIGP0ARVALID  : out    vl_logic;
        MAXIGP0AWADDR   : out    vl_logic_vector(31 downto 0);
        MAXIGP0AWBURST  : out    vl_logic_vector(1 downto 0);
        MAXIGP0AWCACHE  : out    vl_logic_vector(3 downto 0);
        MAXIGP0AWID     : out    vl_logic_vector(11 downto 0);
        MAXIGP0AWLEN    : out    vl_logic_vector(3 downto 0);
        MAXIGP0AWLOCK   : out    vl_logic_vector(1 downto 0);
        MAXIGP0AWPROT   : out    vl_logic_vector(2 downto 0);
        MAXIGP0AWQOS    : out    vl_logic_vector(3 downto 0);
        MAXIGP0AWSIZE   : out    vl_logic_vector(1 downto 0);
        MAXIGP0AWVALID  : out    vl_logic;
        MAXIGP0BREADY   : out    vl_logic;
        MAXIGP0RREADY   : out    vl_logic;
        MAXIGP0WDATA    : out    vl_logic_vector(31 downto 0);
        MAXIGP0WID      : out    vl_logic_vector(11 downto 0);
        MAXIGP0WLAST    : out    vl_logic;
        MAXIGP0WSTRB    : out    vl_logic_vector(3 downto 0);
        MAXIGP0WVALID   : out    vl_logic;
        MAXIGP1ARADDR   : out    vl_logic_vector(31 downto 0);
        MAXIGP1ARBURST  : out    vl_logic_vector(1 downto 0);
        MAXIGP1ARCACHE  : out    vl_logic_vector(3 downto 0);
        MAXIGP1ARESETN  : out    vl_logic;
        MAXIGP1ARID     : out    vl_logic_vector(11 downto 0);
        MAXIGP1ARLEN    : out    vl_logic_vector(3 downto 0);
        MAXIGP1ARLOCK   : out    vl_logic_vector(1 downto 0);
        MAXIGP1ARPROT   : out    vl_logic_vector(2 downto 0);
        MAXIGP1ARQOS    : out    vl_logic_vector(3 downto 0);
        MAXIGP1ARSIZE   : out    vl_logic_vector(1 downto 0);
        MAXIGP1ARVALID  : out    vl_logic;
        MAXIGP1AWADDR   : out    vl_logic_vector(31 downto 0);
        MAXIGP1AWBURST  : out    vl_logic_vector(1 downto 0);
        MAXIGP1AWCACHE  : out    vl_logic_vector(3 downto 0);
        MAXIGP1AWID     : out    vl_logic_vector(11 downto 0);
        MAXIGP1AWLEN    : out    vl_logic_vector(3 downto 0);
        MAXIGP1AWLOCK   : out    vl_logic_vector(1 downto 0);
        MAXIGP1AWPROT   : out    vl_logic_vector(2 downto 0);
        MAXIGP1AWQOS    : out    vl_logic_vector(3 downto 0);
        MAXIGP1AWSIZE   : out    vl_logic_vector(1 downto 0);
        MAXIGP1AWVALID  : out    vl_logic;
        MAXIGP1BREADY   : out    vl_logic;
        MAXIGP1RREADY   : out    vl_logic;
        MAXIGP1WDATA    : out    vl_logic_vector(31 downto 0);
        MAXIGP1WID      : out    vl_logic_vector(11 downto 0);
        MAXIGP1WLAST    : out    vl_logic;
        MAXIGP1WSTRB    : out    vl_logic_vector(3 downto 0);
        MAXIGP1WVALID   : out    vl_logic;
        SAXIACPARESETN  : out    vl_logic;
        SAXIACPARREADY  : out    vl_logic;
        SAXIACPAWREADY  : out    vl_logic;
        SAXIACPBID      : out    vl_logic_vector(2 downto 0);
        SAXIACPBRESP    : out    vl_logic_vector(1 downto 0);
        SAXIACPBVALID   : out    vl_logic;
        SAXIACPRDATA    : out    vl_logic_vector(63 downto 0);
        SAXIACPRID      : out    vl_logic_vector(2 downto 0);
        SAXIACPRLAST    : out    vl_logic;
        SAXIACPRRESP    : out    vl_logic_vector(1 downto 0);
        SAXIACPRVALID   : out    vl_logic;
        SAXIACPWREADY   : out    vl_logic;
        SAXIGP0ARESETN  : out    vl_logic;
        SAXIGP0ARREADY  : out    vl_logic;
        SAXIGP0AWREADY  : out    vl_logic;
        SAXIGP0BID      : out    vl_logic_vector(5 downto 0);
        SAXIGP0BRESP    : out    vl_logic_vector(1 downto 0);
        SAXIGP0BVALID   : out    vl_logic;
        SAXIGP0RDATA    : out    vl_logic_vector(31 downto 0);
        SAXIGP0RID      : out    vl_logic_vector(5 downto 0);
        SAXIGP0RLAST    : out    vl_logic;
        SAXIGP0RRESP    : out    vl_logic_vector(1 downto 0);
        SAXIGP0RVALID   : out    vl_logic;
        SAXIGP0WREADY   : out    vl_logic;
        SAXIGP1ARESETN  : out    vl_logic;
        SAXIGP1ARREADY  : out    vl_logic;
        SAXIGP1AWREADY  : out    vl_logic;
        SAXIGP1BID      : out    vl_logic_vector(5 downto 0);
        SAXIGP1BRESP    : out    vl_logic_vector(1 downto 0);
        SAXIGP1BVALID   : out    vl_logic;
        SAXIGP1RDATA    : out    vl_logic_vector(31 downto 0);
        SAXIGP1RID      : out    vl_logic_vector(5 downto 0);
        SAXIGP1RLAST    : out    vl_logic;
        SAXIGP1RRESP    : out    vl_logic_vector(1 downto 0);
        SAXIGP1RVALID   : out    vl_logic;
        SAXIGP1WREADY   : out    vl_logic;
        SAXIHP0ARESETN  : out    vl_logic;
        SAXIHP0ARREADY  : out    vl_logic;
        SAXIHP0AWREADY  : out    vl_logic;
        SAXIHP0BID      : out    vl_logic_vector(5 downto 0);
        SAXIHP0BRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP0BVALID   : out    vl_logic;
        SAXIHP0RACOUNT  : out    vl_logic_vector(2 downto 0);
        SAXIHP0RCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP0RDATA    : out    vl_logic_vector(63 downto 0);
        SAXIHP0RID      : out    vl_logic_vector(5 downto 0);
        SAXIHP0RLAST    : out    vl_logic;
        SAXIHP0RRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP0RVALID   : out    vl_logic;
        SAXIHP0WACOUNT  : out    vl_logic_vector(5 downto 0);
        SAXIHP0WCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP0WREADY   : out    vl_logic;
        SAXIHP1ARESETN  : out    vl_logic;
        SAXIHP1ARREADY  : out    vl_logic;
        SAXIHP1AWREADY  : out    vl_logic;
        SAXIHP1BID      : out    vl_logic_vector(5 downto 0);
        SAXIHP1BRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP1BVALID   : out    vl_logic;
        SAXIHP1RACOUNT  : out    vl_logic_vector(2 downto 0);
        SAXIHP1RCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP1RDATA    : out    vl_logic_vector(63 downto 0);
        SAXIHP1RID      : out    vl_logic_vector(5 downto 0);
        SAXIHP1RLAST    : out    vl_logic;
        SAXIHP1RRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP1RVALID   : out    vl_logic;
        SAXIHP1WACOUNT  : out    vl_logic_vector(5 downto 0);
        SAXIHP1WCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP1WREADY   : out    vl_logic;
        SAXIHP2ARESETN  : out    vl_logic;
        SAXIHP2ARREADY  : out    vl_logic;
        SAXIHP2AWREADY  : out    vl_logic;
        SAXIHP2BID      : out    vl_logic_vector(5 downto 0);
        SAXIHP2BRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP2BVALID   : out    vl_logic;
        SAXIHP2RACOUNT  : out    vl_logic_vector(2 downto 0);
        SAXIHP2RCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP2RDATA    : out    vl_logic_vector(63 downto 0);
        SAXIHP2RID      : out    vl_logic_vector(5 downto 0);
        SAXIHP2RLAST    : out    vl_logic;
        SAXIHP2RRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP2RVALID   : out    vl_logic;
        SAXIHP2WACOUNT  : out    vl_logic_vector(5 downto 0);
        SAXIHP2WCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP2WREADY   : out    vl_logic;
        SAXIHP3ARESETN  : out    vl_logic;
        SAXIHP3ARREADY  : out    vl_logic;
        SAXIHP3AWREADY  : out    vl_logic;
        SAXIHP3BID      : out    vl_logic_vector(5 downto 0);
        SAXIHP3BRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP3BVALID   : out    vl_logic;
        SAXIHP3RACOUNT  : out    vl_logic_vector(2 downto 0);
        SAXIHP3RCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP3RDATA    : out    vl_logic_vector(63 downto 0);
        SAXIHP3RID      : out    vl_logic_vector(5 downto 0);
        SAXIHP3RLAST    : out    vl_logic;
        SAXIHP3RRESP    : out    vl_logic_vector(1 downto 0);
        SAXIHP3RVALID   : out    vl_logic;
        SAXIHP3WACOUNT  : out    vl_logic_vector(5 downto 0);
        SAXIHP3WCOUNT   : out    vl_logic_vector(7 downto 0);
        SAXIHP3WREADY   : out    vl_logic;
        DDRA            : inout  vl_logic_vector(14 downto 0);
        DDRBA           : inout  vl_logic_vector(2 downto 0);
        DDRCASB         : inout  vl_logic;
        DDRCKE          : inout  vl_logic;
        DDRCKN          : inout  vl_logic;
        DDRCKP          : inout  vl_logic;
        DDRCSB          : inout  vl_logic;
        DDRDM           : inout  vl_logic_vector(3 downto 0);
        DDRDQ           : inout  vl_logic_vector(31 downto 0);
        DDRDQSN         : inout  vl_logic_vector(3 downto 0);
        DDRDQSP         : inout  vl_logic_vector(3 downto 0);
        DDRDRSTB        : inout  vl_logic;
        DDRODT          : inout  vl_logic;
        DDRRASB         : inout  vl_logic;
        DDRVRN          : inout  vl_logic;
        DDRVRP          : inout  vl_logic;
        DDRWEB          : inout  vl_logic;
        MIO             : inout  vl_logic_vector(53 downto 0);
        PSCLK           : inout  vl_logic;
        PSPORB          : inout  vl_logic;
        PSSRSTB         : inout  vl_logic;
        DDRARB          : in     vl_logic_vector(3 downto 0);
        DMA0ACLK        : in     vl_logic;
        DMA0DAREADY     : in     vl_logic;
        DMA0DRLAST      : in     vl_logic;
        DMA0DRTYPE      : in     vl_logic_vector(1 downto 0);
        DMA0DRVALID     : in     vl_logic;
        DMA1ACLK        : in     vl_logic;
        DMA1DAREADY     : in     vl_logic;
        DMA1DRLAST      : in     vl_logic;
        DMA1DRTYPE      : in     vl_logic_vector(1 downto 0);
        DMA1DRVALID     : in     vl_logic;
        DMA2ACLK        : in     vl_logic;
        DMA2DAREADY     : in     vl_logic;
        DMA2DRLAST      : in     vl_logic;
        DMA2DRTYPE      : in     vl_logic_vector(1 downto 0);
        DMA2DRVALID     : in     vl_logic;
        DMA3ACLK        : in     vl_logic;
        DMA3DAREADY     : in     vl_logic;
        DMA3DRLAST      : in     vl_logic;
        DMA3DRTYPE      : in     vl_logic_vector(1 downto 0);
        DMA3DRVALID     : in     vl_logic;
        EMIOCAN0PHYRX   : in     vl_logic;
        EMIOCAN1PHYRX   : in     vl_logic;
        EMIOENET0EXTINTIN: in     vl_logic;
        EMIOENET0GMIICOL: in     vl_logic;
        EMIOENET0GMIICRS: in     vl_logic;
        EMIOENET0GMIIRXCLK: in     vl_logic;
        EMIOENET0GMIIRXD: in     vl_logic_vector(7 downto 0);
        EMIOENET0GMIIRXDV: in     vl_logic;
        EMIOENET0GMIIRXER: in     vl_logic;
        EMIOENET0GMIITXCLK: in     vl_logic;
        EMIOENET0MDIOI  : in     vl_logic;
        EMIOENET1EXTINTIN: in     vl_logic;
        EMIOENET1GMIICOL: in     vl_logic;
        EMIOENET1GMIICRS: in     vl_logic;
        EMIOENET1GMIIRXCLK: in     vl_logic;
        EMIOENET1GMIIRXD: in     vl_logic_vector(7 downto 0);
        EMIOENET1GMIIRXDV: in     vl_logic;
        EMIOENET1GMIIRXER: in     vl_logic;
        EMIOENET1GMIITXCLK: in     vl_logic;
        EMIOENET1MDIOI  : in     vl_logic;
        EMIOGPIOI       : in     vl_logic_vector(63 downto 0);
        EMIOI2C0SCLI    : in     vl_logic;
        EMIOI2C0SDAI    : in     vl_logic;
        EMIOI2C1SCLI    : in     vl_logic;
        EMIOI2C1SDAI    : in     vl_logic;
        EMIOPJTAGTCK    : in     vl_logic;
        EMIOPJTAGTDI    : in     vl_logic;
        EMIOPJTAGTMS    : in     vl_logic;
        EMIOSDIO0CDN    : in     vl_logic;
        EMIOSDIO0CLKFB  : in     vl_logic;
        EMIOSDIO0CMDI   : in     vl_logic;
        EMIOSDIO0DATAI  : in     vl_logic_vector(3 downto 0);
        EMIOSDIO0WP     : in     vl_logic;
        EMIOSDIO1CDN    : in     vl_logic;
        EMIOSDIO1CLKFB  : in     vl_logic;
        EMIOSDIO1CMDI   : in     vl_logic;
        EMIOSDIO1DATAI  : in     vl_logic_vector(3 downto 0);
        EMIOSDIO1WP     : in     vl_logic;
        EMIOSPI0MI      : in     vl_logic;
        EMIOSPI0SCLKI   : in     vl_logic;
        EMIOSPI0SI      : in     vl_logic;
        EMIOSPI0SSIN    : in     vl_logic;
        EMIOSPI1MI      : in     vl_logic;
        EMIOSPI1SCLKI   : in     vl_logic;
        EMIOSPI1SI      : in     vl_logic;
        EMIOSPI1SSIN    : in     vl_logic;
        EMIOSRAMINTIN   : in     vl_logic;
        EMIOTRACECLK    : in     vl_logic;
        EMIOTTC0CLKI    : in     vl_logic_vector(2 downto 0);
        EMIOTTC1CLKI    : in     vl_logic_vector(2 downto 0);
        EMIOUART0CTSN   : in     vl_logic;
        EMIOUART0DCDN   : in     vl_logic;
        EMIOUART0DSRN   : in     vl_logic;
        EMIOUART0RIN    : in     vl_logic;
        EMIOUART0RX     : in     vl_logic;
        EMIOUART1CTSN   : in     vl_logic;
        EMIOUART1DCDN   : in     vl_logic;
        EMIOUART1DSRN   : in     vl_logic;
        EMIOUART1RIN    : in     vl_logic;
        EMIOUART1RX     : in     vl_logic;
        EMIOUSB0VBUSPWRFAULT: in     vl_logic;
        EMIOUSB1VBUSPWRFAULT: in     vl_logic;
        EMIOWDTCLKI     : in     vl_logic;
        EVENTEVENTI     : in     vl_logic;
        FCLKCLKTRIGN    : in     vl_logic_vector(3 downto 0);
        FPGAIDLEN       : in     vl_logic;
        FTMDTRACEINATID : in     vl_logic_vector(3 downto 0);
        FTMDTRACEINCLOCK: in     vl_logic;
        FTMDTRACEINDATA : in     vl_logic_vector(31 downto 0);
        FTMDTRACEINVALID: in     vl_logic;
        FTMTF2PDEBUG    : in     vl_logic_vector(31 downto 0);
        FTMTF2PTRIG     : in     vl_logic_vector(3 downto 0);
        FTMTP2FTRIGACK  : in     vl_logic_vector(3 downto 0);
        IRQF2P          : in     vl_logic_vector(19 downto 0);
        MAXIGP0ACLK     : in     vl_logic;
        MAXIGP0ARREADY  : in     vl_logic;
        MAXIGP0AWREADY  : in     vl_logic;
        MAXIGP0BID      : in     vl_logic_vector(11 downto 0);
        MAXIGP0BRESP    : in     vl_logic_vector(1 downto 0);
        MAXIGP0BVALID   : in     vl_logic;
        MAXIGP0RDATA    : in     vl_logic_vector(31 downto 0);
        MAXIGP0RID      : in     vl_logic_vector(11 downto 0);
        MAXIGP0RLAST    : in     vl_logic;
        MAXIGP0RRESP    : in     vl_logic_vector(1 downto 0);
        MAXIGP0RVALID   : in     vl_logic;
        MAXIGP0WREADY   : in     vl_logic;
        MAXIGP1ACLK     : in     vl_logic;
        MAXIGP1ARREADY  : in     vl_logic;
        MAXIGP1AWREADY  : in     vl_logic;
        MAXIGP1BID      : in     vl_logic_vector(11 downto 0);
        MAXIGP1BRESP    : in     vl_logic_vector(1 downto 0);
        MAXIGP1BVALID   : in     vl_logic;
        MAXIGP1RDATA    : in     vl_logic_vector(31 downto 0);
        MAXIGP1RID      : in     vl_logic_vector(11 downto 0);
        MAXIGP1RLAST    : in     vl_logic;
        MAXIGP1RRESP    : in     vl_logic_vector(1 downto 0);
        MAXIGP1RVALID   : in     vl_logic;
        MAXIGP1WREADY   : in     vl_logic;
        SAXIACPACLK     : in     vl_logic;
        SAXIACPARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIACPARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIACPARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIACPARID     : in     vl_logic_vector(2 downto 0);
        SAXIACPARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIACPARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIACPARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIACPARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIACPARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIACPARUSER   : in     vl_logic_vector(4 downto 0);
        SAXIACPARVALID  : in     vl_logic;
        SAXIACPAWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIACPAWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIACPAWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIACPAWID     : in     vl_logic_vector(2 downto 0);
        SAXIACPAWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIACPAWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIACPAWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIACPAWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIACPAWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIACPAWUSER   : in     vl_logic_vector(4 downto 0);
        SAXIACPAWVALID  : in     vl_logic;
        SAXIACPBREADY   : in     vl_logic;
        SAXIACPRREADY   : in     vl_logic;
        SAXIACPWDATA    : in     vl_logic_vector(63 downto 0);
        SAXIACPWID      : in     vl_logic_vector(2 downto 0);
        SAXIACPWLAST    : in     vl_logic;
        SAXIACPWSTRB    : in     vl_logic_vector(7 downto 0);
        SAXIACPWVALID   : in     vl_logic;
        SAXIGP0ACLK     : in     vl_logic;
        SAXIGP0ARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIGP0ARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIGP0ARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIGP0ARID     : in     vl_logic_vector(5 downto 0);
        SAXIGP0ARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIGP0ARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIGP0ARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIGP0ARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIGP0ARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIGP0ARVALID  : in     vl_logic;
        SAXIGP0AWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIGP0AWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIGP0AWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIGP0AWID     : in     vl_logic_vector(5 downto 0);
        SAXIGP0AWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIGP0AWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIGP0AWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIGP0AWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIGP0AWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIGP0AWVALID  : in     vl_logic;
        SAXIGP0BREADY   : in     vl_logic;
        SAXIGP0RREADY   : in     vl_logic;
        SAXIGP0WDATA    : in     vl_logic_vector(31 downto 0);
        SAXIGP0WID      : in     vl_logic_vector(5 downto 0);
        SAXIGP0WLAST    : in     vl_logic;
        SAXIGP0WSTRB    : in     vl_logic_vector(3 downto 0);
        SAXIGP0WVALID   : in     vl_logic;
        SAXIGP1ACLK     : in     vl_logic;
        SAXIGP1ARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIGP1ARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIGP1ARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIGP1ARID     : in     vl_logic_vector(5 downto 0);
        SAXIGP1ARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIGP1ARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIGP1ARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIGP1ARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIGP1ARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIGP1ARVALID  : in     vl_logic;
        SAXIGP1AWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIGP1AWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIGP1AWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIGP1AWID     : in     vl_logic_vector(5 downto 0);
        SAXIGP1AWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIGP1AWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIGP1AWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIGP1AWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIGP1AWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIGP1AWVALID  : in     vl_logic;
        SAXIGP1BREADY   : in     vl_logic;
        SAXIGP1RREADY   : in     vl_logic;
        SAXIGP1WDATA    : in     vl_logic_vector(31 downto 0);
        SAXIGP1WID      : in     vl_logic_vector(5 downto 0);
        SAXIGP1WLAST    : in     vl_logic;
        SAXIGP1WSTRB    : in     vl_logic_vector(3 downto 0);
        SAXIGP1WVALID   : in     vl_logic;
        SAXIHP0ACLK     : in     vl_logic;
        SAXIHP0ARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP0ARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP0ARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP0ARID     : in     vl_logic_vector(5 downto 0);
        SAXIHP0ARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP0ARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP0ARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP0ARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP0ARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP0ARVALID  : in     vl_logic;
        SAXIHP0AWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP0AWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP0AWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP0AWID     : in     vl_logic_vector(5 downto 0);
        SAXIHP0AWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP0AWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP0AWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP0AWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP0AWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP0AWVALID  : in     vl_logic;
        SAXIHP0BREADY   : in     vl_logic;
        SAXIHP0RDISSUECAP1EN: in     vl_logic;
        SAXIHP0RREADY   : in     vl_logic;
        SAXIHP0WDATA    : in     vl_logic_vector(63 downto 0);
        SAXIHP0WID      : in     vl_logic_vector(5 downto 0);
        SAXIHP0WLAST    : in     vl_logic;
        SAXIHP0WRISSUECAP1EN: in     vl_logic;
        SAXIHP0WSTRB    : in     vl_logic_vector(7 downto 0);
        SAXIHP0WVALID   : in     vl_logic;
        SAXIHP1ACLK     : in     vl_logic;
        SAXIHP1ARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP1ARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP1ARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP1ARID     : in     vl_logic_vector(5 downto 0);
        SAXIHP1ARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP1ARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP1ARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP1ARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP1ARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP1ARVALID  : in     vl_logic;
        SAXIHP1AWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP1AWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP1AWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP1AWID     : in     vl_logic_vector(5 downto 0);
        SAXIHP1AWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP1AWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP1AWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP1AWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP1AWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP1AWVALID  : in     vl_logic;
        SAXIHP1BREADY   : in     vl_logic;
        SAXIHP1RDISSUECAP1EN: in     vl_logic;
        SAXIHP1RREADY   : in     vl_logic;
        SAXIHP1WDATA    : in     vl_logic_vector(63 downto 0);
        SAXIHP1WID      : in     vl_logic_vector(5 downto 0);
        SAXIHP1WLAST    : in     vl_logic;
        SAXIHP1WRISSUECAP1EN: in     vl_logic;
        SAXIHP1WSTRB    : in     vl_logic_vector(7 downto 0);
        SAXIHP1WVALID   : in     vl_logic;
        SAXIHP2ACLK     : in     vl_logic;
        SAXIHP2ARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP2ARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP2ARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP2ARID     : in     vl_logic_vector(5 downto 0);
        SAXIHP2ARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP2ARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP2ARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP2ARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP2ARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP2ARVALID  : in     vl_logic;
        SAXIHP2AWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP2AWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP2AWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP2AWID     : in     vl_logic_vector(5 downto 0);
        SAXIHP2AWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP2AWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP2AWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP2AWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP2AWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP2AWVALID  : in     vl_logic;
        SAXIHP2BREADY   : in     vl_logic;
        SAXIHP2RDISSUECAP1EN: in     vl_logic;
        SAXIHP2RREADY   : in     vl_logic;
        SAXIHP2WDATA    : in     vl_logic_vector(63 downto 0);
        SAXIHP2WID      : in     vl_logic_vector(5 downto 0);
        SAXIHP2WLAST    : in     vl_logic;
        SAXIHP2WRISSUECAP1EN: in     vl_logic;
        SAXIHP2WSTRB    : in     vl_logic_vector(7 downto 0);
        SAXIHP2WVALID   : in     vl_logic;
        SAXIHP3ACLK     : in     vl_logic;
        SAXIHP3ARADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP3ARBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP3ARCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP3ARID     : in     vl_logic_vector(5 downto 0);
        SAXIHP3ARLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP3ARLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP3ARPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP3ARQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP3ARSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP3ARVALID  : in     vl_logic;
        SAXIHP3AWADDR   : in     vl_logic_vector(31 downto 0);
        SAXIHP3AWBURST  : in     vl_logic_vector(1 downto 0);
        SAXIHP3AWCACHE  : in     vl_logic_vector(3 downto 0);
        SAXIHP3AWID     : in     vl_logic_vector(5 downto 0);
        SAXIHP3AWLEN    : in     vl_logic_vector(3 downto 0);
        SAXIHP3AWLOCK   : in     vl_logic_vector(1 downto 0);
        SAXIHP3AWPROT   : in     vl_logic_vector(2 downto 0);
        SAXIHP3AWQOS    : in     vl_logic_vector(3 downto 0);
        SAXIHP3AWSIZE   : in     vl_logic_vector(1 downto 0);
        SAXIHP3AWVALID  : in     vl_logic;
        SAXIHP3BREADY   : in     vl_logic;
        SAXIHP3RDISSUECAP1EN: in     vl_logic;
        SAXIHP3RREADY   : in     vl_logic;
        SAXIHP3WDATA    : in     vl_logic_vector(63 downto 0);
        SAXIHP3WID      : in     vl_logic_vector(5 downto 0);
        SAXIHP3WLAST    : in     vl_logic;
        SAXIHP3WRISSUECAP1EN: in     vl_logic;
        SAXIHP3WSTRB    : in     vl_logic_vector(7 downto 0);
        SAXIHP3WVALID   : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
end X_PS7;
