`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6W8NadMpXVL0oVF3XMaL35H3iK1EllmZGxhJEg++p7NxE8X3W6hBctvgIlNkpOP/
kxClkzyRedc9/qU8wehrdKhVT5IcEmqWtP9uk/dQg2Y1Qeje4aH8y87QtiqeR9nB
IPm2Ovp8hf7liCNR+cWK5ju4DavmLwVadZ/ZM41x8ZnVqZDXr4l+0BEgojIXVIFR
4V/t7eXuPwR6gMtt2nu7WS76GreKoQ9mcp6+ELLbo4f/7yGYYkAEg9sJmFOhd3iv
O5AfFJ4hWjRSUBz0aH1YQkESawmrh9g9YKEwxcQg0jsKBLbwTmTkH8Dt5TQeeJ3b
D6V8piOX+W6PJrYxMWLRvUdS74KWDIAcs9h1uzDBn23IFQpiCaNxW268beG4FHUm
K82SD8EhlspY0xtLIyoS/jDIt+p1S1JSJH8NGjO3in6zv5F5ZdwRDyeH5D7qBfjH
vOSP4EHbOc+RQrudJ05GaDZqefUbdQBDj8ssKt+L1u9fvDcEKqDgWCTCYlElKpZj
xi3lJiN+k43tdWBhH9z8KcsB4XzcGyhh5w6zd7Ugi5tyjGP2U5VBYUeBsMokHFvB
SIJRs85Twtq6yQZooR6C8RBo7QKvyfqTprD0GxJ/5VYMQc9eaBEi83wwYHegxgia
S4LkCyRF5NWNkManuUFk3j7LeCQMJo/FPRR0RvQqmfU0UR+aRtjpV1AKc+Iui47x
/cdBlH/BhAgfm5PlfYB3id8frWiOtytFqanAxcNN5gpTQyQdP47NX8Ggj5lXn8qf
16majPBzJN220Fwbg6tUvhqIsEkrm9OfKrPmLKyQUDbLFpcfgvQkuoE3Do7J9Ra2
2UEaCOH7PEG+ddur+d4fzgFgCUk60vWI2kvRJ1VP0ecTxPrL+O+wQ66//65fbUpm
jZB2S5lAYKJ6abqw8f4WEXEeH3Z58/Gn+laNDp0nHwIU+3xA3skBYvSZ/2Agtvr1
4pO9z1l7ePsawzna4YHWA1YKwarqwxkZNb3c0fdWE1Cmt06Bsb6MUojicGewnWxw
7VE2cdoT0OolicUCa6PPmR8AJmEpmBefI568zVkZ+Rn9w4Y1YvLIHqFonK66ch7F
Byzn1GtqRIBSPyEFVGaaaixjJ6D+fcIqJTcKFNawkNEndpT+abXXYzQAVKYsAS+C
0K7q4mNXY8hDcu1wEC4sBXTUp5Ou/b64Ly6kQz25jqouKUpDUda2ZlGpV3qT9kpX
qGhoy+BDw/fuxd7+tluYm3qiw5MhQUy2p8mbSq7xa4VhdT293z+O2srytaYS1/e7
ByA0bAc462RblKECiIVLS9GGh5BF4IHVGzGzASsXqKNvR2y5BgTrsOXYnQtrilbg
Pw+dK441hNls/W7mysve7CE74qUFWmvmavyl/eqz/qGyB4gt1KnJPcjOg1DYhFFa
6kopWxYObpzn/P34pO75zBeWf3jdnoI361bgNjGR68hTCBVUlYgJrAA1D1nsyytn
eTmu+Yid9ien54I5bq0tgNxvQjiaEk0Aw9CoNkq6Mn/VVny9m7eWtAnS9XCkPFON
c4+QzJfyFhHDSfZa7bFm0LtIla5ZnRA+x6OxWZFwC4hosqzfRGEo2OP0+41rToJo
suhjyg62+3EjI/lyA2VExb7dF2hhVu1Y4XoLBIQShG0I/Eq+LXwIOHukR9aRtzhU
KfPWnv7K0Kb291IQDehBsq+fRT9pl3BKjb2oLsjR26itytdRXUiccPCD9dzrrHG4
1jJLprm5s7pCocKE+m67xY7pMAsD5e1it0K8/2fRI40J0zGME7s7VEZ83USFGf7V
WCcu/0uWrvZ585JyfJYCNT79kSJTW05ivRiN5mXMrX32WkROupIf4UjduHPqs26z
opsWL+iMikE9GYzFMCCDoNCzM9CA2iRoVjgexkqranw9TDgSmsdh/2cGit76951o
RXuHmesWOQgtGbP3Vkj6rjhzLSbT8mhHKONMwfDh/rdKYrVQZFZ0ObOXO3Ts/eTm
YmGxszDYVAxyW8wXT2qbRpHOLuNG63MdOKrOneaM4NLCAJQjuL5Q7mBNh0q+UUiX
e57jRpXivB9Jvx3TDvKDLRkBssfiRUWW7n7XjUpJfWR9KSXGNEnkhyRZUbnM3EkG
C9aRW7ZOXPxQJFadHlupfacvxRWb90jC4TsrVKqr1wPtH+/9KNhiG2An/VPlu7LY
y6NvtkoOkKjI3KYcGJMUdn+Q2pfH3o7K4FnJ/zHLSmJmcxtz2veW+ZN0jQwor6mz
5Dxo+9vTXcghVNNKnmlqvjKghLvsWfZtkdcmRTqH/XlJ8+WAKZ9vwT6wlq8zbqv5
uqGlHK8JJB1bL/IFAiBvY0bxwPyVRZgh0xaEbqwA1pneT0itJ9bBEkIQ8w9RB1RA
7dh8ULfKDGExRZDRQgM7PjF/sEusS6iDBvDctzrgCDxBJg16ZoYOPWFx7fNrW6gR
OYYopUEfoSXSvQ7ktKZmNOIFXmWR/anZvVXuaCZx1I+kEFP/vJoz/62kpEQ0b49F
yb4YMQFSPzF50WmDBp1imQ==
`protect END_PROTECTED
