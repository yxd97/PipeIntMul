`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tc81ERzKeQ1CK2RPzqEGPBmI1wVlKUtVUekX4tzMuAQ4tb37WRaGe9vVZjyF0DYy
79AR/eXv2LLADj8G9+F8ttVogp4SqmCofIMvKF8rTE8/IvOa9iBDDZqnAl0Cs3X6
OYjyuVv88b2va4H6dGrmKTytakRmIVQZntpnMWWhp3v9evZ6U56nMkylri+EjVO0
/D93ysj7A4tdB87KH4Or/6SvaL3/U/5jLL1IjjkY0TuyOWUqivSm5tghC2CYZwF1
rRK4dXsjsVGr88FLaCDFJMYKamKwpLkyhU1a6P1CpK4=
`protect END_PROTECTED
