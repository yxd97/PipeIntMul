`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FyP+3Bm6q9IsByvy0J2f8L/6LOi0/y4LJf9bMfB2Oot5XcGa0rdqrm7dPCpdvNWU
goZPGiXoBJTw3LcBsSa+MarIq7rNxZ2EihadJSkixQOYY5fmc6dZahHG6yYau9bv
lDT2YRplsP1tbzgfWg6WzJfMLykhbYHOIPfuyZZ/LXXuJl/xzAf2cmvHXzKII6LZ
3dyy+whaY+d7Hffi+wIQvgurQF+AxxTjkKWtHXkIVV/+rmRWW7NDEEOhCAm1q3V6
DaUsGcKG01seQp1AAvFi4FggA5+Jnh0Pa/bYNmLGP5ryp87qFK0DKIcfed5sy88P
w5e7BltsdNSeXn9+zQEKdTRGA/uJnwBulxrEMDeabo8=
`protect END_PROTECTED
