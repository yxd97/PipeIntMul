`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J90AFMmUUKCIf37yTP3xwcQlgOVNejGwltW3J0cDsprlunjXWz1kOs74dNtIH8Ph
qzpay1GefV4rdyLTB676pljVBQEvu3JW5gDGV5k5u/sJtH87tZv2I8zeUqaG5GQG
mOtoJwZpF97GdBmMSPxI9Oj5atOWGgMFk8kBAvuZif8BD4JaaVQ9t9wixSUXjdpe
P7XXlRV/YPqJ8zv8Q3BfoEEz73RGNSKanw00LWyBMg6mqpDhOwn94vIY2GEz8GeT
UXxoOehDEcy7TiI/fyyYzuMw1sV3sJasEjCuFtRED6NA4d261Io1Kb+MWJwkZ8kj
jMudnDSB4B54QWr/CcnSty19lUNsRYkc0NUwI/Jv2YV8xziGle5KLqAmkeOPZDP9
ubYRmTxcotqctvPuWTuGsvA7fpZmwIM0wzcxaUgkza55cQbKPzQ4c/16l4ydeSz3
/NDUmuv69l1y2yZCBDSRxcHLA1mP+wdxrywgjIP5SrWO7R36cyEoRK3eqqXj3sil
XcfnTGdZPOaCuI848L7NYod+xMnv1GCKSluuDAFE3j21ri+2dslyZw9IMLzBlRfT
WvPSyeqGimqUOEyzdnxo0s84oeWZyloExFB7W3RyLzpYdNUvC51pdjGJBMXCrLR8
IOgh5w+78s+eya+q1XVLJPfUWnvpup3DdxwDi2xe+EfQ5HMjsp7QtYM6b6qG0LSW
pcJHXj7dhtM8PoMzeB4uzoNA/Jg3BBV3TZoo5Z+J2yXCXykg9iXzUxtyt48FjLkc
rO5xPiAqac+OgfQSIo6hzhf0fN6FZK3YmFwpRf86wxmrzAhRykuHUDUC980a+tla
/JIoFCxgO3d6HxaJEJ5oI1msldj6b2DcNm/nEZWNnGODFpRwLisDo5HMZsuhAWhq
qnJqq2hcNBBDTI6DfwgmH2CDTdGI+Gp1D4DvA5QjAiQNtg6eQltW3a+jo4ECezE0
IlMqqnBJhlKc1uHzGitHunuetuiOCmVPoAPsywI24U7SxYwQCPqG6owPlApGPKgg
W8jWIrMB2Dfzzm5ztmMcvrHolDLEnNY6Qeq1C4NTiP9ygZJXG54gkHIO5eun9hOo
8q3GPh5wWIRzrHshtDoVVMS62f2So0w7xVHY4j91Kl0Nn44kT/5BJSTG3RtpNotS
pqyv0cMhmiqquQV/kFVQZhQRO/zefh/5lKHOukaCTD0kTHorizauxkwuTzL+55de
o7dTtrpWNykQ6VhVh7UMypaHVuSbnAO3RT1QW+DB7KStxV7w0sR6XxaSz9QhDWB5
81WIKl8ZAqLc5qhVD6Mbk0DxREw+SLAkRbhLO5yu3eGD90seROS9V01ckU3ZUBfA
ZCWnz4RAu0sNHcHyfs0dJfi0rTCZAQoCOgnjSVFLJVFo1bEwsI0YDY+ps6nzkgpY
NCbM2cnaH4jbF+i8tQVsxznI7sTZeoes84+Sw1d5/6K+4lC+8v5/jJub1PKmv8hR
NcQ9mgkgpD4e+lO7hZreh3X2hCY+4PxgnizhcyFZfHlZI0rhJUfpVK/1WcRDtein
Cmtvx4a1AeelwwRY8Z86xrYtsIFciFSgsOluWNIUbcGny30x77EqdtwWZU7G+Td6
u13QtH84vsJl69UpU0YCWryu4a8it3OPj/zvYs6JgZgVeIO9Mpn8X3SLVUpMjFMN
BhcDgX5H/fVLXxUhn0r5qAoVUuy5fvIlQSlE3HRODqWUeEJs5I+rPlAp8XKqSY1+
avY4fghJ/3L2oDNZbheqvnLK/HY0QKbR3ZWYjTOSnV3xZg7/f7vr2JdZN+hxuB2N
13E4tSp2H+3P2G7Yh/y4m8rZS0H8ooGbZsAhmTsqeEYrhRgzenVF/YByUcLJCOai
akkVrd3YikHlCm+KwzfpAY5sTLXlnnUxoIPLSvBEc/03kc+8sYyuJ8nG0SxZm0DU
ClOcboGt1KrHIXMnNZTn5AYHqkuh8Kb8O73kMkJ+nutPqyFlDoytC9miCGwJbZJF
O22N95SklZrUVeUUk6uUuEV7s+86bh8b2Q/9nDQ0JoG//MBSVYgvCLiY3bG9gm2E
XMcXFpkSKRxxMhjkR40bv6F2a3UU0WRM9AJTM7yaIcpovM5QM5gYkBnIXohO/GDy
QhRjkQycWtXXceopHptc9VhEqD2Sye9+TAXURr/cR2H/KkXN75MzZCoaSoXRXutg
VYNPWd4xKGUBEeC9MsK0WQ==
`protect END_PROTECTED
