`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3xCnZUe/1oBD3n1LEnbEhULA64v0o33UkkPQwehQLHigoXc9fu/N6+ArU8RaGndc
JPpCWUUcy1sMTXG1mVf4pVvJLWbOim6TifOeBCXY2buvvDOE6438zvbeBnBl+9nN
RHXGx/nnDcpAk9F0vi+3502NNafVBLuJvVHiLzTKuie10urOgTe4OI2PzqPRca4v
CcQB0sgF0KrYMmBHQKxt16Z5J4M025Ah7jma0IVI44K9udxuNY6kGL5337FgKuLb
JgfOFCojtrtKxdgUvAfrmXSebFR3vnJwPw/KszbGwyC+DxjBxtGqNqnB3JDyrq4H
0F2nIQokQNH7gVWYpnTxqRKfa49adT60diVGtBHsA5puMiktvdiYJwUar5DcyX53
gOX8T3ahbWHMr12bQx/7ojA+amt4Kg9o+xgiRrTdvZaDX/Bfc/mca3bYv1ZqwORH
CuTQORQRTMHHyaRtR0EDkOZU8fkaQ+ViMgwUGZbX5qVWvI19gf+sG+Byo6pM5nKg
`protect END_PROTECTED
