`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y9lRIaAXyyd95/VTaZgPpjOsk2D7jJN29RDpK3x7EQDcmX/G+p1VNaqQfb1u1oAA
4ixcluYI16GBRwdwJLUoSg0oetjguEuhrpxeuqtXORZZWHiqmmd2xR/qSfE8pEpf
Yk/8/fvmT49KVxd5Oyj4NJCAXIQDZf3jUIidqSyJsIkpJBJntJOSCxCYIKELvpUm
S5B4hPYkcwruU0qfX8Y3ayOVYO2slELhxXoVtxL0KcqVV2uJKwttO/yAc9xkUEdk
xbPPAv1AV/bjm9PVTq8arTJ0zqLRzG2LZuEOCkMEyx47NjH6IdQecLD4y+a1vySI
gGrOhFwr1G1FvcdSUqKFEIwvKwFFc5Bl7aEIPyDVFKCz88Fe46cYL6zknlZoezV4
mHHv7QUy1ydVVXA6L+f+yjtoG+awSViwgXMayrMHZP//+JOdRwBBeBlmSRMYjSNv
4JQIOJouZ7t/vn7x0utQwC4aRU5NOht053XWcHmBxm5PNT5WQIfa6EvtlfFuBDVx
6cJkNvBe9Q9MB4KhV7evMSOUT3ImfUR2/6IziMgARy6BF+h2fUnX4MqgDBObFTEh
kdOUbn2SLUIw9Rja6Z7P36mvkMzbra+GBoKefzovUUpbj3hmA9rq2LmQAvPfnspP
0R69vj0ltJtDquC0j4cmSBPAhzZFUKBLIBjbopKDhDbLnTL0T+OwkjlIWOdQaKrr
mRCpX5b3ne1KeU7f5esGMVXsZqYvMdPeT/oQt6a9JlWejRafr9R4Yw9AmNLRxWL5
ykMPwtok29NhxKyrxFHTutK7zG8GvqWtQ1sj6WcbwtNHcMqETRio5b1zDonwod1C
0SZaUCHcX9Gnkp/+j8vmtYRqGd0n+bJ1CeEfXpanWc9UiqE2NKXGcr/AZcrZ8ZkA
tFOlry7Ni5Zr7gF8BRGtOQPkfPo6r6c1WNncoX9dIU0oiA5VxbjyOn1j9ZJQahBc
Ofhne32fobu3DSTahRcSY+wM57Z116q2zDBzaoXmHyr9jrkkaLoYy2BcmQBsk+cc
yNh4CqYOj0ZA+JMnZaBy+cmUZXK4g14w3+VrVUolunWwtvftfo2Rnan//OEw8wOm
nN8pg0GMfCvW/+rIF+gfD5gs4UrvRLDOWLCrSolvGRC2IyixOz0DDAQcP/hQ5HrX
F0Jwg5JBbIKHxxCmsYn8JMxz7NLNveKcX8ZeG9JeGKCNSbc40jUclGVpBU46sLPG
QFHIPLsbUQLqztvJVFNmqk3JmGdWMhSl4/Wzvj9WcLj8l+GyzVQhQKkjHEGydt/c
GPSZaBWmxRTYbHb4toPmLkUl6KLX0WFGMm7pxHSHxbR/4KKvrQSUdkzPypoI7uf9
Olg4YSVPT0aiJ7J/2Ab06FxrDDz6jhgOnm9RLvsbM0p0Hn3zZHA5N91C6xWuJqAB
`protect END_PROTECTED
