`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMqLUPFL7kAmwPbfY9a25q6T2ygoEGmsaeJZSVEaPU57NKBjyZZ077XwKLiZ6psj
o8oCS8Bl7+cmXvUGk0Ygqebp3yDIqm3qM9oMuCM8nwTHWhg7yefpK36zCWNILev9
l6JD2vD1rdRbVDOuReu6mMF/RyLJO+6qQoUXFdxs47xQ86gnVFWuuOjgi4T8BkuG
t1aKdCjl9myFaa8x7odfcmHgv49I5V6khDlOCfp6Rwdjx1knDkBNAtSbAEeolMhJ
+x/xIn3yulq1bQLcJPzC4hL7JPspOsY++1Lm8blpi6oMCKwxICWMv+AcRHKQAjku
6X0EHMF+VNjWo4aIzCoAexRnr8x1w4aRzKWNcYdgIts75LbyRIZwRSemw0Skfs7B
/QKqDqj1qVPj3z03ZimzPWD+YzhH1VKpTs1YC7gxYHz/PjeMOGjvhyY3npFXL025
WFUMoVbcpUjfMR4MKigqim1GT3QF8TRLf/lFYofnLv0=
`protect END_PROTECTED
