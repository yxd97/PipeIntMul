`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uu32P7ZimvrW+7/3E+cbzRCiokV0Nje3Kpv2Iou3u5dcL7z2Ir6z0kFTEwZfFvvP
xbqk5hvOocGFz+83MEQDkZ/figTNUDYJlsV4Rcw0FjH/bZlJJdHKT7BZ1LX9eN0Y
mMieovG2vaZS3HZS4Mfatrjt7R8NSlFNBNweF5idMaYKUGWCx3DE6sXN2Vfx5gKP
x2NT8icF/XQXMzstdw+LL05AMcZ+AJ6+DW1KH/E+41lm0l5G8nZ399RytZb7WciF
foaIxm0F7vajoeVSjebSea5dsOLq5escjANdKG43mmOw7o4cQIspNxQaVKif9PLo
X5jVOz5sJu3KM0fR8syPnhYIiEp9ue6C+J4VANuCZq4D+QfEDMhcGTgmPl4w9/oe
qbQmm4fvKf/MF72kLt4nFsGjcaib4+IcfNzIMASf3y8vEDCqyPtTL4cviTRQr6V6
TSmzB1LC3iOmTHmwRCvgBHBv4q0egWZLTbuv0RpsFegmrSKMqQnhoCp+P8S5f5J3
gR4raTAYwS2nMaPAgritInXcCDdTGPgt5vlUJIsvjV+N7Ughw4bF89T6azhg+UpY
IsYlt33Aa7ihxzxXnbBel2snGzlv9xt3/ZBmVZ6bEqfG58gWGbfYWcTzMyO3Bw62
QL8y1MdwitnFhv+npdBbWVu85cultUuzVQ/cKRlgA57s/LzZh7Rx0jhli7ciTMyR
wteix0mHZ++8RB9OQPKNogo4KBpDvaDbO05yG1bETN8F1XoVpN6Pz+K3WTDxPSc3
i3nTfhxFYRV6P7m6/Q8lVpKnLUHN+Jc4Uq9wkeHLJaC+8lNpbJaCa5HHImeYS2nk
JStpDhC+1ImFSG6lVbCNAB2Kjecbwmg44KUdXO7NjCdFoaWG/rtuOXE71HbNK2FY
fb/NIKIbKtppq5FtYhGVeSoma+37B9VxW1U935LS3tYoTuOHhcNRDaNHezNi0DJV
ZVB6v+sXNTjUlf7JuLwVr38zxnyUfqG4dRfc9R+6U8DnlaTCIk2wrKRlNAn0n91Q
L8u37soFy5+AqC5dqLFjW015NfXJapSEL7ItzZkhoyjdasyDvUY5HIE8bVgWZ+BI
n+BJOtk5tLB4+xgUCZxf1zd8X1G24HD1+MJR0bXN1C/GCaSV+4zHDlmaJTGqZ6H4
x2hAeDZCcBIHtMiUo1JIGzhWKSgD6IhRpLdBiwUCPEoCmQlArQhhE5OOw8UnWFXg
GyUEXqU549ldl2XAMyZ0s8L++LsL9PsnBt/j3iYCqutZknw+w+RE9ud+HDBWdEZD
PhMnksPMYbTiVP59ywhQd2KWFAttxiWnSE/fvF2xjXNjxt06gUBH11qT6jYmAW0D
VOHxiB1Fq87Dp0ussHEX6zAqoZPpegj2tjVP0uzwgc/wlhf1igO1Ejc/6DOflFxp
kHMP5MWgxTmxahur0WdgIOH287pQDTFayFXNyFu2j/fy3KG76H6e3pUeHObM8Wta
3GAmUGoUA+Z9OiJcE+OgNtj1idWiXsvrfn92sAk/CE/dtX02bejEffXnt9m5RGVT
Nwj9saMcz9o+baSZ1R7KAGaxsy+5/n2m+0W+HUh0BYpKsEqdL867CeRCy1w1FThE
j52H/Gc0Fi3XgDQuLNhBpYKPorRrWORbXx1mTaM7i2REAuoiS12ZCfP4gq5yRivc
KxBXwRR5mSEbH5LqmtIH0iK8WR1uFE+1G+J6+NY89xwxrDIcdJ9tUKLs4Ja1LSow
0xfvFr18G2HvwsF+9icmpdY79kWIy0rdjKaKlXhbdJLT+guIqowBDR+VW+jBYUJK
qQcIGqDPlLorVlCaZy/LOa8dkuJ9mz32k+YuKxsxlBfzOn43lh5s3SROt1oC/LKO
1iH9n8URvueP37sdvkKBawxRm6fT5ynHahC9ePaRde1Qb7evpnbfAdbApCFjRtNz
fyaKKypv6/g7tFcRFRdNkHdrKxuANhmBynOG/HylucyWHFsOx4PHSzZzc1fTt7kG
oW9VZUS+4OZBh2A2vzq/M6NzefGAmevyaqRPu9USO8g/iIVz9o77DxyKK6pWqIMz
XhiJXYHv1zoRXmolj3n8l7ad5pthaYP5JNxCXXITrw56GAuSPemNdrIqZ5gxpPty
kzYOp+4OUhMP0QKEGbq4QS36HzXCITeztMDwj9yGp/Fd20RT7VyYwUnX2FnfZaam
lOEDA1GANxWRVn1P/iPbtZ69wys3RFRBFplpn/CtOl4h/YPfVDT3c7mEY6GXO29D
g+4sqyiCrMihcp4+C3CDrhu2kXdFd6BO+ViU2BRAJADJxXxu6ZRir6xg7EFwFLNg
fSrpXmDtLEiWApwn03QAsdx0J65Vdv9q+8tQNvkpk8twEkrr2Gbpum/YFQYiTbfe
Y9IO+zR3D+VmGffxmSnCnV1wt16kVIgExUu8u+D2h9ayCzsLNrihsgeCp+Mr+d9r
HD7lmZWsFuTgXDYrqVlPg+Zr3xTWGvY2EmGh5Qy7xOpO78t18MDpdhwnUEKr26w1
rR0QdhoXtAnd067AkYg8cwIOsRRsNbLcJcmtERl+LThMyI9whNm0SNHDumIJRDm0
O2lPozhUnXAFC7T+TP2Ao4dtD0uQ68tyQ2NHLUx8y/JwmI4BfS7sT5MqRIyB/0ru
mu0pjm8L9Oh3O9WKOY6k2G9d7qUi+kxC08Do8UIYabrxyejosQoxICVq5vd0x7Zu
PrF4nZ1Yu7Too7qKELmVcHpy+e0rqFhoJucsv+j/RoXENEa8FBfJeXTjwcUVhgcf
Cm3SgWEYJKOu6Nfej3GcXf/wf4iTWWEOyhGjEAMXw4q76IMPAd0w29X7FBNyJexe
ScOKJXFUdKn64TbRU/vIRBN37wTapmbCVeRiPxMdQehtAefp3lhqDZDl06f9nicA
HEPDSiZO5rKyZalgCNc7udBPAoWBeNnuFiZ/FtkRxLOIhHlFka/eNbwynRHKMWOa
xWMXTmYnHCczgzwFQTSdez/4/W0oJcPp5g5WijNMVV3fccybfyny0jfam3VscqSZ
nRh/ZMuKmDy9KREAe5LHsJruPNJu5pxkGZFirtWc2mD3J5sFJhY87Y+hmhZ2Q+/B
wZz3Ht6YvBgthZVttmfw/va9EM6Otm8lJSUC2QlX8Z2hydx+hFwLzEtEUZrmJgPz
PFN9isVX8xbHf3aZ0gn6AfCQwlQ+o07AFhQnaLnRMSdF8rvyXej2PQY8Jr+qwfG0
lO0n3R+aLMtJWB7kAwZkHD8tZEW/IpouLaarCjZkhPCjlMUpxaWQz4RtjPdFU+Gn
cxPNVqLmS/tivw7M4atrObm/JMQE1vneQi8clRnBIJVOs6Wm9DKfUHCeFm86BT+X
gtE5DVrzNCC7oNwDDvKF7gaZPkUmW6VH1vwAatwAARF7lDmvbzV8+OJTBKgaL5Wv
CED6MSxZB+cRPGyl+83Z21I/NiAH4G3Mp6PNNiPb+clCwvLyRMJBYgHtHZhe+Y06
/hwsEZNJ68oiMruIrtMjfviG0s644//Z7Q2vwHsNpFAxvnKlVqdl3I4z5wqG6zi1
PIO48fOARH2135BbbPfIrLkEjPKVlJMX7NcMsWOi312Ekyx4q1foDkLTAfA6T5j7
cLmsaDO0Kz0siUbBSP9VKehE7Tl3zmfQXjFRIQg0kYERpJ88toMQ0y05aESTY0OY
Qh+iVSmYW5ZrEGk19OIenaQmSQPXJak8bSAl0EnSW9oTUoZsR8GVyA5AL2Fc3Ukr
pVOJl7ls5OQb5NEK4NTBYlSPmGfPtI26+GliYuoW6nddjM/JkZyMhDf90ZsL33cI
4gCiD2ZKBkGg4tMcQEACV1cn6gTt7xhKeDUP5j4yMie4It/xmS0LNap4V/I3R4nN
vYxCCPvi+EttZuzFZk9Bz/wSpClvGI1ndxqarbMUBnlyZZahMaPPJy1w00o+5gEI
tiLWtQ6b5gdT0fJ+CGlBB7ybcMe4xnx6EXq+qEFqmcGdrBzWKY4RdP7og1UmaIUv
sXTpIywkj8RT/qH3I9hn8BI3v0xHPe1uccbtP4hVBjADawONglil1vuBcQJ1IDJj
D4U+OosOnRqADHd9roNdqvxJa5xm05kvpOFisKN9lHEzCLpXcCQ56w1p0mIbg11V
xcZwgAFJfX+rzSLiwZtBjgKWDQa1iHtpppxPAdFIUxkk2mQEH0y7rK9HFDGZ6l8M
U7E44e1div//lcA3mPTXaPtqEkEDm15cwkSzqIQTgPiadk6A3GS7TAOg5YkG7EaE
SnC91DUcr0WD/N69lNW4VfDVVTbuR437fuUxaoMSFDBNF/H7g+y3SrPHbrBWpfYC
wv/IdLCb+yPcsDlPDWklCA2k54WHa+Brs8EZtGzAnaAEUxPFrvxlQ2UC1/+ac2t1
5u4SPdqDx23Pc6/naz1JDTS1+lAkgHepDEkWVNvX3MiETq0rii1Hwd8khB6K9YnX
HJ0F1gjBFIyUbrmQwLLvHhQt+ylw04ebTyLK0mHrxbvcN+YYZAIptPQPvp89I8gh
74nodUDp8f3R3kNtMHXoClOzSBgV3FFQuTFWnZgaDI4=
`protect END_PROTECTED
