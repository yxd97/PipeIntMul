`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gB1MNT3nSVoWdzT8gQe20EUOcM5G8CSXJd7+/iiRYMiveMpZdfsnBxdSFxHWNakm
0nL5ZorkiIbdYBthzLTbYEmMQrXJgYNfW4R1xRUG7QrniBuXZxMRhAWMF7o87MPo
XnpTMGIC1qi7vOwGVKBSEb5JuZqUWptcShvzqI5WW/Fec4Q77TYQZuJxun8iu/jM
rR7UlEdyrww5lkDtuKqQvgD5KiqOBA90g/+CINs74bO4nbAGSWtw9ixO9BdV4url
PZbkb9uZ3Y0nMAe2epH1BSmkRoN8Z7doSH/e0PcN9NbwCn6fdLg/EfPWIuDxGlYC
ahtd1xjSNPJpBq3sTIq7+o0x2B9IjUDlEb8pM58nbQ31hwfWDhBL+eHTQGAH6Vo5
3L6YQYJTonvgYsY0koQxy7rVkj2VV05l3TjZYQUDD66rYfut/dfXyhLR6nrQo3Yu
0CptMjkNawoOlc2HLb0KtxK/lpYlmOAl2xr03sQAFLx1CZfmBQ7m1yznuOCFf6bK
yyfGXdyQVr1XZIwxztOwTS8jnasb/xmuSqVXy4r21SNTEQCHSFcseq0EOm4JW/AL
yRolVz4ikrE2PaicdM+H5vRsqNdFAcSoX4kQlgXIFkF/DQiwzKUiPe/Llm6iamap
8aH9+z1dcBcJik0Z+oR4qQ==
`protect END_PROTECTED
