`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4SNrTKiKTmczwgCSqMn8+27GSa1PIJgOhWxT8VCeeBIlUhttWKWSbQA2DqWV7gm
fWTwtrkGDeK5Hb+EfYhmnL7wCXxe/1+y25gZ9w/m0HC/p4ve/HZi6HIg52eA0EBR
bLcgVsEs5TlJ0CMZtS8XFlJ4UiUZTlIj1YGQjgEb6bJLoKxpJzaIBpnh29To4R2x
Y+WJDsdAh6r2ZLsv69iXcYr7wqn+YKYgpYg9YIbBvAL454q0BUTNLNku9k5UZTwy
d+2DxUucCxNcw0kFClhuUIbJlT9B93qMrt86jamxdyGuBvDSWI19ItEiTHbKALEQ
uLD7DyBrmjjGuU0f7yzZbfHve9SW0AMOHAipZq824dyGDrjQr0u1DtxfS2mn6vlv
2+NgUv0fnxUCn6z9V542Z6S/rX32ARPkYpquasfWUqg=
`protect END_PROTECTED
