`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W4XbKS4CKjUGo73FozxpOgAQDDbeMwrKUeHtcoZRpsokBpKKAMM7yaIFiD4T26NP
lxk9XvSEjqY49aClNtZOJ5M06M2roRiURIRYbIK2X8K7m1gSh1fUzBEWYnhw+8sy
LS0FPYv2H4PLYGbTNB/AhP0yj37Jn84u5IH1MGlfUOERj1ltgrbedRCFHUyOaCKt
55rUfVRhvLSCV2YEyyITBo+Gz+tmj7cCeC76xMTMBfNCC8xqeUPNoyx0nqZjowCP
dZEGJb0vc3J2NfbpXtAoaM2BaHHa9kkxUkCIPET2F3bVoJDW3W1RJ82cYmiZmBRD
9f3mCqBUF7uIfYGS6ylyyQ==
`protect END_PROTECTED
