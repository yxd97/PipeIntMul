`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQtYJ/iOwFZbYveSSmkeLpzwkZT1THXgpepCWC6kHoScz/HOxaCnAdGE85BGSc8R
eQqleKiIpU3S85B5llnASvnXPiBiUELkAlf79xukwox+VbVvOGJS0HR687PHDGZy
Z49QD7W9Fa9je6++opSacOuWh1Ijsvp3godGovGRMnufGr/efpPhfehEFi0lWXnq
aj53ndy/crJprVVqhAyn4clK6fzkGW8UPO0SoIdTG3SuJus1ubUrJp+hA+CCgKS7
OZV5aTKYIJhtqbyJ5i/+NQ0N5W/ZY3k6INETH4VekTly+H3UR/d9GCKqsPZ6BIFx
GIFfTFOUekDzLdOJoyqnYg==
`protect END_PROTECTED
