`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u13JWa/BfRWQHNl/qUqAt9ELUOp2dj6tCk2aw9kmNG2DdLNOTOy/L8XlOulABRYV
orsUZQf5/FJTRzJvrDZ2y15JCqO/nmop4GYenA5G+EPtdic3JHs+1UbnTul0Is7V
POuuMNa0INu2SpS+AW6fG3EeaOhft4o7VEyPBKm0XNjRBLe9kS+7KQpIY4uwToJj
atVPLIlbzaM4fNTonBYXz8PEb6TJ0Q3i4QbF00soC8R01NjEvWFKf5KImkMWtmHJ
GlScB1tJGyNOBcMpsrVKBcLVbZ+RlRhg7MlhBa7sPt+/WsDBZ201kmBMQsLdFErl
zstSGnr9buV1D9iGtvwDA69Y8EmKZ5W4gIn7hmjNaU7p/BJZ2rOusMKYu9jtnClG
89KVq1qQM9LUhS79IsGwFFVgkocf9ebbF9cB926BIreuqrNKkaW6CslOegLVZsdA
Cmkdw5MzIbcu+3HYp++t0ta5TKvERdyUoDB9JkZFDLTPYfihYaT1f9RW66TmsGea
`protect END_PROTECTED
