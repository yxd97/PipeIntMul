`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UAAWFUFw5cDodZYcXpmvl9NZoOq3BKw5PAUIUji1zxn49ZJaT02fwE0DTMBpwu+C
3Y8PE5VOfMGi3LnTXddZCtagFnHgpu7TkQrDqYt57i+zCQJ1bMZ0wLIvkHUScP3w
il/XufgbtXGZthM1FQdaKtoKltq2k2Uz50wWZmxxQM0tFZNmDWPyqHnsAwSny7l5
cSdUqE8lXyiWRTe1eJ+XDu6mop7po8ZazBs8BmnKtw1t+LUjh9io93HcFnvePT8P
jMjCBsnglTAwwAK8b8auRA+U05r5Bzy1027aWnAYCpyHJG8qWqSJNrni/kUbiS4L
ALTyXlNhyZUudRH+JwTgcmIGzpPVqNPzevjcH05eGzYhXycchmlRW/thenQo8Qrs
+IT4Kb9VZMcSogj/hcZmZg==
`protect END_PROTECTED
