`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwD/QJAVE3h5PQp0qqf4tJmARYqcb8r6zAiGYmT+PdAq8EJnV2yeKw7ozuToBy/D
XGKGx21ldwUKwXSwVjebZMCAcqR4MwDH/E4v9yVW55giOwJT1DN0XZseXI6hl8fV
PGUboaUruSyLkgltVPGrqExzMq2+6lmQydv4FhPVzDGbuH+DZw6MrmU4eV6VW9Vv
gToLbOGH1wNKS94L8XloWMin7deu/Wyu8HKneINdRjgdvNuZoN+/JJW3m6TXTk5J
POiopcKTWPTkkDAuSJG2nf4OsMGNlYhSq+8blkQbFMQzP9QTKz8KCTTx/DnAkUpN
JZWsTRAmlSr5i1imRuWvAQzJFKygBfhbPiF9JO/DgohXhgE6+fv+HPizA7SQ+hrI
7YtJEdfimFMcNTt0GrTzDg==
`protect END_PROTECTED
