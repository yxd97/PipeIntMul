`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YhdfqtmBGUWK1en3WBEKpVYb1zAfilkxGhhO9ORj5E4XBPQ6iGzNjc+I/cdPR6QH
XawMaIRsTB0OwEfHv+lIXpXwAcBNu2bWFz8uiV7aB/WUYg/1YHXxodr6Zs1YhI7r
lej0kt2SHDtWzdISaPScP1X1jj6Qp7UvzPIV+yasgSlFMHmLix+B0QsbmSnuDnG3
3ydaDmwzzeuYbnX3RJQFVCPw0EiF7sjdEqqXOA14tnmuG7JjhUqh2jpbFda/Q4oP
RLv334EmwA0L+GMcspQwNGBEZCb8E4mx7FKoVTWMuhLMaD+APsaQ0piCn641DZ8b
cQc5aUmpRl1uoVJDn1HKv2HLwRycDDffJCkWEO2bdqVOxiflOsdsVegZl8Iov9kO
zBfg8L1xbudZe0iNXGiuycJXQSP2Cv7kb0HvEsrv2IzgmAkZC4ckf97alSErXdr9
j980Bjw4CQrUTa+bbH6oOfwHHaAUiSdlFHm0jRHo+2u79kRtm/nPQooLS3nQMjas
`protect END_PROTECTED
