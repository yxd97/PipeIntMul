`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OgsRRllmf+lpK+Kdfz+fh1f5lYhHvDHq7W74jqx5udgkPHf6T9LcrFSI80INYMq
QKpQa3HLPfQtnT5C2n+OSFWtzXmi04WurkEmqF2DZGm9UbNXsdWJwhx833eoCHGo
4UWO+KxJQfr+dWyPwEBX/Y5vR061rAP1NQQ0LD2HbUWZpwOjlFTAchEllkS11PDw
jdlERXIVM6GGgAokx7bUFp8f6kFXA8+3cpdp4paCgt94IByRRg35iDdMxfRrBhM9
lv+UITgIyrE30hOmX0hPDhOFADZIA9pGj0DMFgSlHBoobOPIRrsTdwIsV0eRHwwu
WpyYLVUbD+1SjgOZg2tVhop/bncgrPAkGi7kuqfbJH31U3FmdUZdBEX1CEPthgxT
yq+LOr0u/1ghi10Gmuew2XBl0Tfs92TdNzwrfCdX1Hdl3pGkY5p9xdZk/jymdWu5
jnC890SIk/T97dOMowTDdZJA0xauuvrfO+rMTMSj43UMkdVhuhrRAXY/T897uQtM
YYReUdgbjS6KjriCCjfSRzYtssEfejuMLUh/JI9anY8WMU8RCT08x5S4HQKDVFWU
+hibwCK8UgtTbwCd6hApaUWqYIWpsPWA81XDTYAmZfcc3iBrBryeaRDVrHm1uze6
UEgybks4HJTokvdDYnRcVSZzWW5rq7IfhZL9vdVO9CKanF33ED1cJgo3B2SPO95V
`protect END_PROTECTED
