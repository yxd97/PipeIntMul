`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uN+ca9OylxySzA0c42RlSdmuxFo50a+xdzQHPScH0Ed6ir2tAlyxcSFqQW4m2WWc
yHLIgFicBW8ougUo6HzAaslemV/q0ormX77onZP7t/FaD44FmeDZ4w/u2YqfH+qz
MqAU5XmF18K2BDHLGcwWrb+DUZzdGPDdsuq+4+tqv5lUbz7HpZbOoYuU8g5GWuEb
XAn3I2LgCUDgBvV1hLhLf47f9tLJvSrVVcOR5Gpg1lRMBOZZAU5/mcvwSxI6/zY8
QaXsnFKeuxXie/oJK56wAqtsIo1yneBqiOsLmIyjcq+RpshHGzOotnoT0kpHgd/R
AGsdz7QdE1HrMgZJrNTBnjACkiuY2CswxLyGo/JV9CyLIJawUXLIHOOlIFHHMtQN
5EOZ107V8HyJMD7Ku/fbbvDmKmGumLw6xKQEsyVaX6Y=
`protect END_PROTECTED
