`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+PM0l3WajSFxqAl0vLs/vHLW60tjex1rJ0eld2rRJrpqaZ2Ced1IPz7JjoraazE
Yxc02SwcaHhRhwspyHjxLu7w4vnYHgU7JJfcH/aqZcAQ8zkPlntOCRs7qc1IH813
xont9C2+2tqY8x25so60ocbx0YBwLABBft7Dh+M1EJfxyBmsrpW9su+Tn9JF4bqS
ves8kC5Yf6DQP3GcHzqBpFBAJ5eZ4szPRIXMvz8SuWqar1+P74vYqmU7GYxwTtDf
lUuAf/Yr7q0XhP0NEKPU7iRs3Opgjl+MS0Dwu4C7zPj5HmqmJiICasXl4U9lvwAf
BnFnbXReG5Bkr8cMy1wh1w==
`protect END_PROTECTED
