`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5U65zfnyVezNC4BJ2xGiQoYYTh6VCZBTqJayjCM8tsL3CG48+31SAR6L7aPh8x33
MezpUFKSKtz2vKtdweTWB3RnU+mQAi5MSWPDL3w6a1n9XbY1vqcGQ1ZaBxH+ULjz
ecX5le6dKNTTIcz7tWzSijalMWqJ1MHULYAxA2scDK3xNlCGs5y6bZ2oq862pqIF
oulN3tisyYxeA54O+fZ6+scoFMtV8I/rhwVi9fdmSIp8thqMCK3Bjls0T77tToS8
TwAb0VB1mcOgiNkvvincShaqo/n8iIZNJIhpwTUTMcW9Z/IX8Y8DHkYiwQERWu93
`protect END_PROTECTED
