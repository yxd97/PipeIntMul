`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3ZyaeYyJLolJ8ad6eDvCzS16hyTDgmwSIZZsJaZMrzHMaimZmzmb7KJ1wyyf1Mq
9+ZPUkxGTzwDshZOxYeRORIHahLM4TUXWhB+ao0XSHeoeKLQ3jS2zQJrTthlIvIX
jiIiEUp3T+H1p4dlqfyJSs6qTfPQTnG/tXxDz+PGSFexDaX7COz3dQ+FXAaZ0gxv
wcp06s77KFnE4JnVSjMpVmuh2jKosg8oLyDI2wVwvgWKjodHSxNOyNBOabMowZ+9
rJ3rr5yJeTLyhPTZLgabos2XdzxaXWXTlz+0IxBtG7REvLFyrlzKtQtXb68vACkw
IpcKMknE3DZQSE/L7SB8EUMxXornlSvHYlCo624riVqs9OVqqy7H4tpn8r2I7Sol
Ef+YqIwL5pxxTCNMRf3evWK/aIQ3oPTLXzqbR6dK3R4ZvFbhdooDtdxh2xVhq0+w
K+gXZE3YPMr5zvfhI2BDLJwMJmafa4hsXj8KPGGoty12Mj5sJRpMPgYXML+8QFYE
d9RoK0mj0flBQI7K+DwS1mHty2zfhw/Wi1+GGyuRGY6bOfRHuRlMvdCPnOOGVlFu
/Vd3NQ5ROLboZhq6/YUA5yN1855PyEY6gumyO9hW5XHfKjIlXJhAwtB0ytzoEzQ5
mgIycm9dDkoDtJ6X9aEamFTp/JJVDy6/q5S6msyQhGM4KJKqqUd+LdH9xfot4dKn
g118f7WziKlZ8JtrBFUkjMdM6bl7iN6jUK8ZOTA8B2wVHqxpwbI7h+1I23RckT2x
VfAYxvCJXST25x7H7FSR08hoZrg76LIa7qH7s/Sq1++NarZ929pN7YMdrNTnEZ7P
2TgA3WhGLhc9kdv+pB7tUSOTt5AgpvJnY/f32ItTv0nE8Zq/0uGGgjFbgKdqQJ4p
cTCzGujIRAwNCmqlp7JfYE2pc3JSP581SqMS3t5WKyhjcbErlQJeba25+muqSf7Y
`protect END_PROTECTED
