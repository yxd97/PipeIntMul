`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IwFhChXFKII/5/TeMqbd00/CvDM0xZ3jaLoqpcQQjPvmmtfUJLcDH4qa7iG+6OIh
Llk3P8b1NuLVBUeunyW9XHDXkzsF3fDXwkx9yeyk8MW0/Tl/g/hmHobhh12MWmxc
nSsoKwANG0i/IOvufhmfa2laGNDKkc1eW7x2Pp9jXlLTWoElwxbuCrouzdSJDyuB
w6Lm+TIJNncu04Flnpq5jcXyTvq3XfGIyytx8pWs5vQ2BlBpKFXM5hhnGSZvatAc
H0/aO9VFLzBXKFl/zzyC49eg61xcZoGnBVbLvfOfI9sczUv5Ne4bcK3OBbhQPxid
JfN5Ro5AhqxJcRnBEllkgzRbT0yjJBPwq7zSa+JR4XCiBgB2j7ywZp4pAVCD0W2f
Bpr81wDqfnoupIM73JnMdXJv2qXVNMde7TpKztNHNLoNgdWSu29kw9Zd07JpJI6z
yY4FbkCug2wWcnhLCAevTePTjnWiw++22eiPfB6x7FandwZJe85qIMEu2n59OAkq
NS2ivUq9m8pRU2BneoCkCW7tZL6JzyC2wgHdFelWCRd1uPQW9yHSv0iQXz8/Md7J
d//NJQhXFpYZkk0DDdsK3AkdBzX5Nh3pxMviGG/a7+GUYBjllxhTSxqsJP7emfuU
YfSI2CrDYbfQnkOJkKm4ENt0Xhx6wJl+P/GRfvyiJbaDWXjQYu4uVqPrmJ8TLcjm
UloAlGGT/0ZPJdFAQenD1XLMDCpJYy+bT+fzIkWlCZxnIw3Prte8XnXQTOJnxhuJ
cG9Y0TlNWf5NHJwAYrql2OYItY6ErZ4DKJgzJ1kU42kqSq/J9Hu+LjpVPu179sI4
ZpX3DMs4DMKQO1XQtoOwlGVg5qNlt+MM/WZ8tgdkZJT9AQLeBLv0AsQLmZVHeAJn
knb4VIfULOMGDHTE8qyv1rIYajevSXguvVbCPZGhw2KAo3wh+1mCeZu3KNfIDCv9
8NDn8meidS70ArzX7qFfQfhB7082sLB54su2s55cUeZwQa7us8Y1sl9xkcuSZ2/S
7vYzUsoDQ958zs3jzmSyIaAYZeytAqVJpKR2pMShQBCE4ipIuuN+lOcnuhKtcsqB
tK2k0FU1m8iR05AGZRDDhWdE72OqKMLePwPU0f0cTS6SE1qFVzEO12YQFh1tIVFS
9+PDHOwQzdjzk3L73IoMbPQSgD7aEpaaZfBu1YHH95KdxVAKyeMwILF105mKxuvy
jfmJt4fh+UvWI5tjeLFqWLE3ZTV1+XjQ34TFrFWsDnWe9qo7N26+dSxT3Q0Oi7n9
Gp5yGvkgQg6CnffxyMMHosirrH/38UmqsA86tZDB85zF7r/CaA1ivjBXYhHIVdxL
fGS+CYT57D8P7J5fgxNouqQetZEb5pQh0oR8NGAFNNuDAh/LzVYmxemopWriIGse
X4QOrV2WOJxvRF25gnm9PFInrKvp4YiD8sbvzpuRFJvhAnADmBF7Hnwx1/9nyzOv
K6yJ/m0knIO4sAeN8816yE70joWPDevjFVUciMNdbF58lF51hhbR9ZNXOxt0SNvF
iccpoPU7c9xcPDarU74Q2K4oKjoiUjGkTqB+hqvUcuOw1JQIUbfFJaHtIWilGKtU
vsdqQOnOaaY0qxR8Py5NNssYFgJ75eDQM7dJrhrIz5ErHvA9yT2FAcdmPAEI9lrY
PjRQmh7jYQq106KI7Kwxeu1t5SIcvKTst4bS5VZK/9HlVjEVF5o6CH2JKU2QCaoK
amnP9+G8M+zGNMHsXLyprglgY/YgM4gtn+d3SGDmCUYy0bAys9zq+y70t9/j8z9K
5mlGL62hySZEVctyFt0dSgI94R542ubSpsmBGdglTMCz+a2bba4f6uJuD64fdwGh
KYyDWCKfPBH7cyf+Sc3DIrXKx/mHeDDqKu59acHtcd8TkKfy+LVUFFz9tHNs5rSH
ZKBg5wKqgPJCtlvQ4nPQ2eJhayCj6AiqqxzkNzAPnbJAlYaWMa8ndXvR/2+KQyYh
OCwn7Oxhud2PUkQbRipazuUyp1aeXYEurfJLjbbPHbnfQsbURp/xbAwCt7fdb0+A
7flHqq6iSOSVERA8fgbSTBiTuyO5hR/FxYudyfhNpevtjN/qDRRoZhCS2iTOO+B4
dOTkRXosP4ThBdlTJEvvQXhhCyfiWEiqkY5BUAIBmpEbw0W5N9JTqN5z+TXkqE6T
2NsuleI+SjsMyfJY1lwv2PR9AwwbytT001j9zhpxCZe3Ncun2KYVwhO9Of5mOD39
FuRGv9Z3xn7st79UcwWCctPmPNpIh3tLGEqlQxdN8HdwjWI96+1oInGxSxrLp1Oa
63+a1jkKGHXqOimmNZp8MlBf6GLq8LO0W748ijzz+M+e6Q8BOphW0MUE44PkcIVK
h2tk6PqDFXhN6m1hJKbxfrpgyZS4EdyDhob6G8Pzy8fHTdRdkSDr9LALjeuPEj+C
Wt2ShbVe1IAM0tR3JYnoGar7umvVxFFo2LWuzd8dN/jCCFCd3qzxY23FM+lH61/j
jb3z1Uwsb3RLwBPCaTMDMy1Ls4pKhVw66n1Y2yxCTcjGHbvmNsWsAjfNJnweSZaB
v5eJJDKSGPlFWujEV1Yz4voJfkTYW7AXmfpVTJhnFt/R5uU99e24xx5M+noI2vCn
sNkkGBfBaT7JcRjXXyKI5A/kbwi0KuLOtcRyer0JulfFrMbw6OJ2mSQ+Q9yljeps
vM0S4/nwB4leXyLfFYMv3csW6DS8N9LVSt+cZHTFg8BAh5kb/7wweE2kfGtztr6y
CoE8jMyYP25pyVlxveRYpkWQqm18vs6/AtSOmQoFQWOxDgExjwfrlVoeTMujOqry
t8Idi77LiR+Vw5jZR1KdLfD6y4m9TQxMoR+3hbhAcrFNqeDtxMR1WHkwZ5crEbiE
8fjC8fdnk5mz2HY+zkirFyX7qFcuy1GGzAIRGBGLAsPOhSTY24x/bucNuIhhUiIS
+sPe45T1wwjUQGQPFLmdxVf7CPj5vm9G6IsmhIT69MPNaeC5Y9lYWuy7nxoEtZBg
pays/JwVTrXhXVjxgVtgEn9sf649vnmR+L/VuwzLzHnLtfl7+qj82z40FJBaaLV0
k2h/nqAQwtokxb5kaNYlB0HgiOY9u5RwQfgPB3BqhzkTo06zGcHgjwKD/+S/C367
QBvEwH3r4QjVYZGnC7/hyJMbswWmFtslbmAwasvC8H66Rvl0FGdadZqlo3EMCI2g
sYKZbPa3wGXiy8gyLlH01fyLZpDM/BtS27ZtnICqrhbtYfPsqEcM/zrZD/DFS3VF
G+CsJuwaJ8lzV8HjSD9paxNoaln6yCLWesQKINmfgi3SURRQ8QJtoms6f7ktlYrh
m753n7tzVST/xZyjTf526SuhGmur0wfH0hoG4cXXCqe/jQ7N6h8yvnC5chH7iVu+
WTm1L1yzqFc8bCDVwDgd/DrV4u8dMm0FQ9RqfbFUTsGowkS13wqq+Vz27t61QXVd
Q1gMc3ID4GL1nvmqGsjrEQWuCAA0rgR+F+2akhjkUdqs4CP68BWw8u5YBagMbXf8
aMuYZvLrr5Zqh1hpL2nW8E6bvZ1vkP9zMzm1Khz95b4vDu9YKzBVOMT5AQPUn0wx
VCB3L+KtwlZNn7AT5K3vqpFRT1MES3G4BOZgR7kv8K0hGfzkeHAgy4ewmJq2SmKD
FdsoOkJ/yzqTC0CMCHWFJMecjKNCRqO6kaGGn06N/6Gnfmy+CF475yFCqfKnY5Ta
sJWU6ZLy6p8WlQ1Az+EGZjbeP1cglbwrbDZplUN/bEjPXAwBcz6TVBCrBf0dLe9a
TztH2ufWNpjmr3Adb/3Kws266vsHXBvX+c5DiWwhqpWHDz6ILsmoPFgmpLmfk13k
c24bNx5Yss8cQtHNUikLh7cPwv9xfCfk6K7O3raTWv5SNmIGNbnVetOgqd8EUuV8
siGPdh9GlJiITiAk+gx+aYZQmb7EKxJKYXUqtoLiFhqLZTY+6v8M73VitpBLEbOF
ELag5yfii5mx8tJ8ISyLsCQZDhZMcbSm6C+Z6BVuLgxGxgkyz2S8Y39I/TOty/d2
7MShH355wvrvncgBHfVahOxWlgjwZOEcMYDjgAYCrlgVB/87wKy7kqVn6Kxzbqge
beGRaoXXwn1/jefzxoc/o/JAHTTTo7ktw2d7zRr+pCXHao3QnDPXGIIKC9TFFYFw
pX4sPdqU1aVfNzMmaT/uqF41tnaX/v25QUI0jZ616wDUHizXue7/TIJP9JaSoBjH
nqSZs6fgnT0xqP7LGoVLPMDPLiedqSSBYoRMuYWzdXvLhDZq/0Jf68vcUGv+ucCl
O/ruzFUjDObSzX7uUm7JdYKiKmUdkGIfPxb7YUwJQK2rekTBHDO4bQ4GsZz/UoSQ
eU4xQnAvwU2ZIcetpFhf+PKypqOlGQHpaMMV8ooEu0tTQwZ6kgUxoZmTeP7PPYkT
WspOZPIajzohmoNUeCTo2bvKTKesEbnvnOeV47pvSfD04dXctH7Vjdhi0Pt721j/
OQzJdx3ulPMZtPLZ+tjLYRgQcA/QHHH6sQpjoq7hnNro2h/TAvhvT9Mv7JUJ1NNv
duAPxKzSj8ZFz3lKybVlRfIF+wURFzgONr7W6r/mCgkrut7WtqLo9Td/JX7WI3VK
NeDUrNnL9rbe/td+h9TidDFU3ZZ4pi+TeVVKw4qNTJWZNU4FGeyQtTf7zbdUCeEy
OA9DKzZpkAPTYdsPtPfO41OcuvIf52PZPViQWBFd9Tces/AFfNA9e/k2xh3EhlMt
1AGjl//G64M8fMCdZ0CWqwHcvDZwOJ49Y2rq16Ae4wSQKeuM1BqU57VWp3VahcgI
Cbot9TSSuHHgHPNRF431N5cysRy5fla/2Hh2Rv325bXogIEdCDE8gJ2pfC9orfVZ
JqRuLnyvVof6EXuwENe1yu1kvoKCJFXMdG84kYBqIEr4Zxy+8h1R7UKsFZJiyWZe
p9dMLjsNNM+ofhL/JjDu6NtDm/+GTFiM65SZq5oV+oIvqfS/BWShCMU7TjYHo6zI
VI9fGbxbZ2OsPyaFGukJTe/dIMO9Ulq4oMOxZ0pD0RlMnaKLh0YEgEOVnbGsZ4r6
Sx/GbR9NWvYIf+yYmcp6qnObi5BWRq4TrHdUBOT4SlRGNr3RcexH4yH+WxanNdSo
dvZP1LQsIxMKLFpJx1Immp95Bv0C+N0iSVO62BwvJGGFXmzjLrxJIa+OErQqkjJ5
lnKYy00epW+5RyU2g4sHSgVtEDaETjL6WzOWkjSZjM9SPoGkK6uVQdxkmDRF+wvt
YnZu5NnEVTExvIkcFEVqIg+tFCgeOhsO7SM8SmnHuyoZyVyQ6kegK6ZSNCajI+tt
/+31hHsQn7iO6qWwsNqc01AQnCby0IeSh3DUPg161JhKXjJjSAeh5TLzH3NAq9pt
6/rDjfi1F7eSNqBH5ylEY1INMhFiGLVKE+8qfTtC3WarC5mkN5V46Yo3Mn2Ajx3R
xbu7pxRlvN3zyrrqqStlARUdxEW5N9C00XHHsOcPZskrnA3BZB/3G0W+BGTg5yyJ
w9jV4z0HYrEIg8COfq6JvTZKi7TYtahJBXgZxkGC+vpjDJIIRmxvKMzPI4gqW/80
aAKWK12QzzrGq1gIHdwDIX1izWZ7jXxZ9yXOt3f2f0KX+Cc1eU/feQbz2yjF/JQ8
9QAkgPQ2A4etN0q91irasHlmxFqFQMDHPvnv/YSoh4kgo0GKaB0IdNEH+G/IUJwb
GZHCS3rJmsYphr/S19QL+g6ImB69rgbR/QHVqjP9C4QmJ7+UlhKL+GAOnv1X+6vg
ai5DmIbccC6WyRxxsetoHYHEmDhfaI4DPxfyM7JzpSDAGBJVykYotwXFWdLQksUT
zT8yUzbcHieSEK4L1x34faSnAc0XKVsaNjnDjKZ86g3ueJJD8LQ2W+VGJA2ot7kk
dE4LQCz0DW8/O0zXHUmKbwEjkgIRYtF8mjFnLFbhx7Izzxxhd+RZG7w4cJ9EN6d+
hePGET8hBAFUuwWGpjPLpyRoR8w0OuXrVATZ+ZkT32w2maR09Z2pjT5GXDwdFu24
0vRoobhc+1ygvhYJ2bOx7T8kpyDzGPsQEdnGraxSrOeMV9rGpZOeXdnA6VahwwKT
WuBgOYfAbkah2iWqchfKf2Lhkg5F4dBdKH+ke3SliVlvx4s7KkBpE3XE8iyicfdB
YFyLAo8LGw+3E4uZQCjuBAsMjMlctS00FMSc+bEsMnloIkOxuVbq6h8BegUoyd3e
1kOJL/Yj5auwW2p8r98eomF/v5LM7WLgST/e5ph2vqbwN355CP7DkqPMu+aJYRzK
L/Iw0k3dyNtI+Tw9CUfJ7r0oFOHcJutxiQr69R6PtvCRELyX5BVAciAvt4CGABks
utUGDJQFklfkmzf4Jyh4KI0Gw5jz4ildyTqfJ3Va/IBM7cF/mlxuob6ZHLeM4823
8PKN5PercwAf1l9dxT9ToUWwDS1lj3BTo3LL7XL0PL4zKI3DjOr/Sy1XbWShA/7L
4ZHibk473iZfqlyEnrS/mmOXny8U340g/WDBaz/ZWB8m5epCMrnt1MbxUBf/dzNs
soyfRmoJDTtYBQZiUE+lP+FEduIXtaRKGG7khrjUhw/8IM2iGwAecI0GsEE1pg2k
0wv0fbl6uBJX0F4nUvF59URmkWkJrqe8BnRXqCBU5xtNnHln7AKSPRdkJMESqeme
ZmLdOu/2i4bxyJuJGrsuoZb+ota7TRhim8ZLuPrys+25uMsk+UO0eYO5qu0R/E2Y
MgyaFG5jK9puUfUo0f7cVTtyU4RuyyLkjFuT8j8NhgWpJY1iZxHNO1Umm8bi1ieb
jB9Ort08IQJcSFLgrOzCeU1ivFgc0t4azotF17YwW1Rs+Yia04NrhuFba7ethaVX
vzasu1D8jcYVZZqrP16EqfjyVzTPCfNvQLvRfpuOGxq3iwZdQSZepQg3zZGQDa/p
TmEdr+eVj0UzhoxqIl4W49WSL8A0IF7GRyxe3/JCyZi12diBK87nKTUBT6x4mlUX
/29QoL4axkDqELX/+AIulk+PoqCzsKseUuniPvDirumqdeUq/XvBHwrzeS9Ez03O
11xdqKz5qaIM7EJywTFGsDJi1WB9W9owMHVi301aUt9iAqx1784T6Nokp+DZD2ai
5S/Higg6QiRimF/vADM1l2K/ScYtoMzrsWSffJVPrAuRItXCwoOq5Gfezfrb44R4
fW2TpVOC8J/xg16UVqnWI84sBsalcKcvf/Y+HMcm2L1TXvHFNWOAE+HzkjHF8TG2
L8a+rlUwRzm+jQApX/nEWHgArMGn5NRR3TRFwc5PIQN0+nhAfzXL7X9iCtod7wCx
Gl6g4voWvCwllasTciag/PJte0Yqni4yCjqREIwFv8Y1aeOJTB/ywR3OTsGNW8pc
zNzIwowBBxGQbs8XjbbV7utr22SMWG/xWF+336jR1+/J7sC0s9iTLBX8vFe69i+j
TLlcuiNFRHstUtDYkkEgnaBn/NSc49Nq1NMJY2iQB4Uegl38opiQMqcArnID15ez
cNI6wGj7Q+p00g66BzWZAbVqkdhXihI47K6v7oTPZO5zGLWPCEICYrTLZWqgHY/m
oRerWeJjfUTUlkwiI67Q23blOf0WUqyRJMufoQ5oYesGa3TtDQJTL0XtOYItpxOX
BpZuDZPUm6nLJQUIN5xvLHccltBJ9fMclX/+8PoLb/9aaxI3BlNy1u+QnNiaH30z
+KvUn3rH0bwFY4lPXif3n9obtd+31nQyT91egRJkx1s/fnZbPMG6ptxGPC0bA42n
5YPbIQ6/0yKey1r/0Oi0UCsQWYmmxyJbzqTuOLF6BQ6XfBR+7IH4ubfs5s5j/7Uq
USqy3G/rKmlvG6p4IXEtldTwY0CA7pgdYTzMs7GFBy6aqj1iq4OE01DOPZxrm2s6
1KTCBiVSPBkcu1JOkR2Tafxe8DclhNMJnGWdNcnEIt8qS2C0fQc+n/y/2Mtjnu5c
B9Aa8ABwAiOKW7FA2KyrwPqLCtwvw8tt4Grez8RZTs1NCle/A6KSoP3Ro8/pxOuV
U6rHoJV58JNFKVz/UyRa1FLJO1zI/OTnKMXbywWezqMikU1vYpxZFWWPOZzaywGI
LSPp678LT5xHj037ttS9KT2x6FVP6omb1K9X5oNFHXwRVTLLc21v+hnGzQsuVxns
evNoS4peynhNnSwXuSzuJOjn5WJNUt7XmIsrU3wJNuH4h3/gKFynqbgV0B/UZIG7
fyX/KDHJndiQsg/HHcTN8ZbmWEZpJj5lQTR1fBg+67is4cyPRzBpbo+YHe8f80Iz
0WPg0tOnCZKRsmwrsORzcHZV2klgaIcLCjVALc/JgTvMIZO4VRRZxvcPAxRueyhH
7R/8qhdLQ1qGMZNZweZtgSx7tM9jtphk6FVczvGfEXZtp19VactGdKWq+QF4Mmay
6YRWVzLfJaYNXeHD5uiNjIv0dMBwpr4kr2C7sS9IVTc8vOgJh6rrq2ckw70JCesp
8KyTZYAFAvHo+PcesqQrFggs3CyFylvQsZ6UaiMylGnBvNDdEL63kZRRgQsltPLg
zFr5lGlfG00E/095WmW+nXd5Eo4cjAMDrQSyp9IiJb6oAaYEfbqD+tKXElsDZ7gq
CzDKzASjs6vHuLTmvoDucHqWrULjN1dYWTwH0k2ffMyJJafww9FpnAc1ouOiHPng
76hRvM2/xi0F+JyiGIEQXa/9JTk2jEcVIFTzscJJr0WGtyWis6aa5PUQpF5uFq6y
l7Y4v7iuDMbMaZLKjd87q6byRt51f5C5JjftIVIanNvEeZeLq9gqr/wMkgs0h/68
rE8UMgvtvTZwd6lNPEJ9d+JdZoXeXXZdvBhgidc00Juvosvw1oRk9VTinhfjo4yY
0f4MHa8drEGp4wLnRNiICXAL22UAgB6wPEtpCWg8V2B+pRG8GA19fAcU0FaQk79e
EyDVVwqOYyqM5tN0ne3+lfHumvwhExJl8F4Pd9qI2cFdOcUna9Ihx5Bc3k4sbKBW
tXyA/SL5pdkHt+ZR2jzzZAlwNpoVDr9+GSk+6iEgDhgPBA7y//3cmE0VmAp0N1cU
zXoucBvFgYX3gyad8OKhyZaBFzZTGCtbCxKnEFNvQCJAQlAvDBaBIe4cmwU1XAO+
hiT2QGsrIaElnvpMUUXoOZfOrv3MmutQMkUVJwoVSbbegzUGK1+xDVOQL51P7lU6
PW3Z5Fu5huiBcSove2nrfPi+ASNaTcrWQKtphZyyz2xedJimwQJKLzxJaG+13Rhu
evMrTmtN3V0+Ev3NeV+oyeqDkqMIz3q/hTiVWcciogB4PG08Ot1AdqhZi9r6gZ8p
fLFUHsAT+zqUIR16HDqdKccAyOxB+M8np0W/OeCmeYqcH6mPWF19eh/EvPHZunlb
iaIRoHyiDRcfz3RiraOOls6jGUIC5Y9KvDDeJbURqXFTve+Rxt3isgCSRNCotd3F
aZP4lT071j1TdDCEQDRJ4CdHP3aOHtvHWLGEthKrlUWUGtSpopeuy07aSzJ32Prb
9rs8XHcG4aTMW0OZ/huN3nD6+dY25c7gaUQs5KDgqlh3Zuz5Puz57wzBLO+NK2A0
W5meILXTLhnBrShouL1+v/iLeBFSgUnzVy+hrRb7dk8l69AQ5J8lmCniO88l11sw
FQGVrqr0PfyuNHoO9l+QyIwGxt/yTRyK9+w16/5/36tJYe4Y88NPKKCQG17ZCuSc
OV5b0OexzJfaX0rOw3pOEjdVqghwEGQHk9KsEeW75QIPg0Pe020CdZDUuz2XMHHW
MqwwpcoPKF8pgXS3rmFw6wYcLc8TndJ38BiEE+MEq9wLDZ/Gr4WzehNBCC6lCx7i
KfMEL+0sx++pFmv0Gp8wzrVFjItiYN92vMv6BCOTDbNSgf6ayQHw4MoFdh4AemgN
RRlVKMQBr9yNEQRa4SnoVGYW9cbujBRmSpbRafkKG005pZTQYd6Fq3Z17vf4EQQq
GBun6ZeImW+Q7sJIElhAN6Nam1aq6hv4swXs8DpPC2Vhkg/dEfC04hzfZ0vepiC3
dOeJ4SwNPXKSlKXYNiJm/SMtmKLyrfvwVDCRktfUZp4T3EecAptKeh99qtDe4cVy
YYZgqFRxZxOWHEv4oxdERtpgy3SROO49hY3HSvqpz8qFu206sm8ao8sCeQV3bmmS
PIaV6fJ59wU5Mw4+LuNjY7I6MXIVJRcXU+3UMjIzO+1f699e2NDCSSgauC8gmfas
Qv8ARx4RUEZRY9U2gTx7ak52WATfDqX3EkqtyA9mUCPiO2P3QfVFUdDpvqdXTD56
NHQ8o+/shjY6BDlkROp2hqU474tqdDCrRJhIg6r90DYeA9bPMz7qMXUcnE10Na6R
BBLEcdunQT6/QEOuHnBseJdx3rIJU5W4zAbP3CDlXpb5VQwfQN+54+NNToE7KG0N
hM5uXAYxzt2PnAoqxmt/bHIGMORkdOJIjPbLGJsRwi0pDzy1EIDj+3mGAHoBwQN7
gndncjlhzLTfMI5Ce5c3FpcWo6gsbH5OYMJ5WA6Hm7J6Or7CQcXKAB/SanxjbwdR
XZrtzbgX8zJcOSk7JqtqLksr04YKbyikj116w+JsHbG67OfU2SB9QNkJe6Vu383b
/lIZjlm3Ewdwfw6r3Nnj0oVjvNfyaOcyA7zx2cASwuGdMxJTQAN+aRXw4Z+DafIF
LINJ2huW281sKO3kh+xNvCExlaYwHvmsBHmI789bjEuFUTUQHKYYrq99CgVfL0/H
milieIg2haEXwGXxIyuZFA6r3+SeIaijSh2IKgBpu57hM+xLOKoPt2kyAv77Ic5G
wpwhz0eYY9zuQHcjkpMhU/BoADng/bTQUGbEzyJ0wfv+gI8i/vfssnDiJwkkPBCH
tD/y0g5alUMJH4z7eJX1EvWv5B2cqgKZ6jjfyJYrd05xt1In5+yFDniP5pseWg9l
p9vrOorfYE0KTvQEYa+Q5tBIGmTIZcsSfW7Y1BYerSH0X8oVYkhpOMyINb3Rayk2
mClQHbSEDYp+Vdw05oH+osY9v+YKNT8eCGQeclbXjwta1XpSMybI0EJ+IrjWtOTD
/kwGyi3bapi6NcQGLGP0xIZbFo0P0Lb6tlgB0/3sZvuPUtJ/T5Y8calBWfR1OQgA
hhTFycIvG7KiWBV2JfG7/YlY3xWpLwcq+Gabie4WADK/ZiPzeZ7lUdBy67U3P+kT
dVEWjNTdcKEX9shymfQbTMOZYpMkxh/alQ5vfFOI5ZF9/+fLpBuJAfWqwKzLP6fc
gAVgwNmN+KQBCAHm28DCuXPPU2QY3L99B++Cpfh5+lO86WynDDeux97CnLhHgcXB
ZCfGMXX398dp7ItZx+9MctHx+pKAEAiPw/BnwBJ8WcGbqTJLuGsPVvYqfUGvq43C
6xNiFnTAdBMLn5OOLZMBVQOiIGpBtNmCwfYCnDVpufgvFOnTle/apIjkfDbDKfNR
yhJbNhAIE7FpHoh1lqwMopGjan7fiQ/RadAktUHp3k8MrUhP9Bod7BCerbri6kQB
Fj8MedviHcHpWUKA3Y0R8e5Ors00lSFqrzXBmTtyOMZcECGuCtnmv5brwutR1lfR
KbIwz3K2Xhy3UOeg1VdFS41fn4iqkipN0xP6OTCNrufBxJERrbAjQ0BP0kWJKwXD
k1JiVNUDpzHhProZRltyKdckZ9nrTlEcRmXO1QpDXsDQPG0qn9tigaIrVTUYaw6P
SgQb1C082BikA+nhmafjpXMkfPa+kPXkIPSVy1fwNc4M6QBnS1p8sVVhdI+2MShP
tgJxBT1VeYsF7oOWgMgcU+lGzMqj7fNKahzB3dz7xKTWlGbU/YR+NRczuaAv+IOC
E0NUFw5vo0CE/FT3QD0TNefQN+AqpG+vwCj+Gqw5lZ9pTC3Tx2nL8VVhKDkFmbmR
A5FHxSelqwhsB8Mf47XwI8ONXs+UoPlr9ovRYwmQhdnb+TVo0QIv12zv7WZxVCI6
lIHoE9ZzfizQhPA/Fa7boQhqkV0jNJo5jIpJyuLYbk6Aheyuc4gEVVrx4fxKcI7I
czYBD1+kOOZdNq+FEN31mq2MW3koXh8+AjenOyNa0+P2Dg3NPLWt2Z8GTilwM6hA
+woNX/GQyl2ywEEZAJRUY0NAZoG+roT9F+W2Zn3MNN+ss1Ed4+WfF0wbR0HkY5rd
9H4nZzjZhkoYxmfoyLbBGdv24Eoz9d5cnElcfeML/JY=
`protect END_PROTECTED
