`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M8JbGwNx+OjBinZ7wbzU96ntyFNDwGvoXhX/aJVy27qm7IRprT2/XhK49aWeDxMu
1jt/NBymYXTGBSKrjnljKYxixTu5JZJwqKDs8LFlyQjjkipVIA7fl30wzeDqY5h7
tIy0AdwGXAVf4WDw3LE5ogBpsHJEsTMlk28w/zgZlS2wng2rlFD9PF7mvH1kiOwg
z9WMBQjWxHImbfmsUVUdQDV02/+ifBs61cmBdMj88M1370JLP5q+dJJkKrmRZX/o
5i5T5J1grETKNZ17LzbWgnwfH6egOceNt59VALkayehOg2lqO+JGoOYZw0MVyUnW
MCuyVTFn2PNXwTwwbZJkKmf1WCel+LmdInvQgYZTVkagdQfHgR58e/McMU320iLi
u28/0Pr+XdwxgFTgrnDqIcxb4xGDPtsRwevPyvqgMzSvc0lJKPQujpbxhH3WVW8Y
v+dglAGDs+NRt83ARsMcwaG6fcizOo2iGLgrmkrkVe2cWDlWCqS+X4kvbMOiFY5z
xuaXff8MSulQEAnCa7JrQ6ZaHzIR5Ok8jbM62nXW1/BSskgdP/Jncnf2d5NqLE9P
KBkTRv7uzqYelaooLKtOXnyL6FyQK/7MOcAopUwJ93ukAzMvpW/EZSXxO7yQqsKA
XZbTOFUivOJbS/KW2aDwYN7ajBeC9a4BDe/deYurWdv6GvHW31VeXJfBY94f0npy
Wkt2WtrprnXBb4TACZQtRDtFZQXpttAS+dvzIH1bBg/BWmwajX1k9y6EEX508aQS
ZfEdjBUFuHa4P7chqfZysMjP0dT9uxmblO8tGMdsj/zEE1REIGz+Mkx5CsPtlEqI
MTPSs/uY9LFBJXsuRQwz3pZmuz3Bji7k2zaz+OCtq2TSg/9CZ9yzRrLFSuTPs00R
t2Mvou7N5gIJq/2m2dUIZDP02ZHbMIskPAE5FAn7cyRa+n6ZPEHJLjdM8Uvjz18e
uBSeKfiQZpns2osaPO5vxRD5Jp1jbAFFudkmKoK3q0MlDLJVIKiXwJocTn1aC9Qa
HoJJyc+RoR1T5ddLVT1R1R3p/lxAM3Oar/BYM6MvM3xlj1r6W4i6kAlGZ7OaNFmn
guDr/OwB/5fvplKkmFmgfiuQfIgfT2pjWkcxH9frSIp9YwSK7yZLH9zEDp3jf1R9
uMo8z8q3w4Raib8gDuWO+v+Ya6jaebcLcg0V+AaOAYU9t2JQV3Q+vIkW8acWQq47
CJQjbrXE0w4NgILcXGZpIShE6iIYxRRaW6RddyC1xKy/hdH/3cc/GSF95XiYXy7w
qMczClwTnuH+2P1mOMaJrKUTJJkyq8QeFQAVFepE3jUOPwwuWRFTCW2qocSfCAsD
ndXt5uqtuygW1bPHm5xJlVK42BfFbCUbzET4Jnw2OG7G2vqLE8youmJ029Dws61l
hAJrabdxpfv1/YCEvrkObI6EvN4ex8atcoycrb4UZnrwVIW05N4Q6wXEoBSpycb2
YCmmR8Hti5JeNpuNPs7Ow/A4m59D3RNZmq4Y4yrRXLlsrutB10sdecRMk2kbzN8H
GiPajkS2D7LhyNhoVQr/O1/ZnMd+dWRPJnDZF7bU5wiHQ3+o8ubRfVu4/gL8n6gi
FHukfLN207ScgqJnvOs6ZU9b8RF4YkXmLVuj3GqSb87t5pn7gkOIsbKVihzioi3p
xiWmUeNcukuq/W7L+DaHntm731JG7Qpt/pwDIxd/6ytQVYlAjKO1RA1a+8b/MGEU
M5l8ee6V8D5lnlbDv97f8hquv6SmcE2TUdY6GLezrz6A0drishVXbKlxqKWCGLSq
5l92YoKhwU9pbbpz2pABKi9ulMKVW8pxImpqXbB+GmGG37u0+2c86hQXgvl77XXb
3lBrClVfV9rG50TlyRgJAcoMtpmNcajiaOV0iaRWqnD5KC9eJRdqqcgUkz7b0oqD
MpySGFmNbAuiMsIfFMEk5LcdAbkDRX6A9ZGwtPJNTnkfE9Qw7BJ4f3lH/4L4HKAr
X/jwpezvqPanF+60gXVZWzvavgb/QqngAGVs2PG0k1mj9WgRndkU8WPeV2ubmcdZ
zAuBgLFUbJZOitcvH5neZqpVOkBEjfn92tdxtWgZMiyerkfz7mf/Z6R1EGjHHI+9
pKxcUlEsW26QFn/mJju4nN8t1kVdahvhtax9VeiOlGLz5Dy8XZTuzXoeWJyqdyQ2
h2UTqHJVafe64+rWs5ljjciQk3CLIbHQpUeKcfMM5eMf+CsSA7+JF410cg+tdja9
q8mwxa6Mv/Iqqyur++wJy62L9lpp8D8QZ3/hukluJvd1s97yFLKML5hd79MDI4w7
Vu5V3zJDdsstvlyJ0iKLEIfjL+xeE/ZVTMA+RJZKNMQAotgphqid7WgZ6WBvgxBq
cbbyVCEWZyxs86z/DXfGEYiDeu/priHnzkUCaeMBosJ0bIndW4tCor7CfpMxj0xB
U7OKuChd0sPOMe71ybZ6nm9WBnhlm3ky6pzvLcJ7qXsvjLPylOl08OP7hfJ8syKg
Ahc5H/rF6XRKryh0I2jbmDWonj18S1z8sb1ivdfCb2VoQzM/kNS2l5AOMPGma/vJ
QTsLjgvwq7Kz+Hkrpu5M/0LBZE2AD7sWAl8QVMppCekwBuWRfl5WXkCr9JeEtxfn
FS2nY7XzF3jAsRQT+P+bIstiw/KXgURZUUHF9kPe/qDaAHFko9Yg9NkqIUHoUAP1
SbRdR0ElTohrTllod6NruTro94IV5jFlqqDKCPTZp+Lft2S891OXpEDSkQJtP3XA
6pttpj5dMfSddW3Y9vcJheHC2NVJsCq7ABTccfyKJkcR+9pqeoAVhGoqF+sZuOlp
yDF2ESBoDoMsLUzWonsFNRQHwUJJMwoUZEg70yrJEA+1AfpKBb2YaoD615YXzyEq
2FdXIENtDEdnrCN02G7xzZBAPjdlhMCd4V5yBTeVHwesQ7n0pwcba1dzwQMKmSq9
/dvQGlgnezu62BPQptA71F/zNvj2DIIIIpZT4FycyvrwZcv5HR8T91Eyz+0up+ga
rQI1j59rBw5VporiQidlz9jvKS/BEgwy8xdO6b3Rop873pXtqlrEeo47xcYkOIzp
ldvAFJDnuyjybq2w8aqakzzy2swq4EsDLADp6monwrFBXXDjBbVO6+9N/lAvgzpA
TICctMZUj3oxdyJp4KzlujAQTG1f3JrwBl1nVw7ob7tg3tRymaPA5bOU97ryp4Eu
qkse0tW/ZK/aovclP1P05LlkUIMhjTxOO1lJJLw6+FjbzW1wkAtjkSxQHfzHEmGO
vMyv+pTzo/fH8SrhAUIUQYrFDImpZ2ykAwXSe5vJJ8b81Dz5C+PHy3ij3LDUigoZ
N8DTIHG40UduAuc4pOc5z4XFz3S1DtWI7kGq6n71PyT0+rCpOj9I62E2/qES7dP7
QUU9IRuPLNCF0RefnMlidwlqnhjb1LAFxenrGK8dyrAUzqDBgNwNycUlqv1NTxNr
CQ67j/RWcD1uWGbLMuxM74tBkMin6g5dvmuywOlsKeQq0yIvhNR4txrnubFyx3W+
Mr3CoYFoAOt9MZ1u8Hqy7wfZN6P7uY8ugrV3i1tT43+MXJm7iUf2HajZc99GdR8T
eilfIgiz0zj6fBR3+mBccGNdRkpG3kc7ccqrvbibJJHkGLbjPHk4d03e523farkV
nZHYH9Uhcq34rY/V1D4qPwP+T0k1KfpDHzoDm14gIHXuFGz15uSOaGRkDJDRtFb5
oBXaHomjnsU34Y9Cdh6+vBziNJ5fO3asgESA+HhQNhSIVUIb5hrbRQMFYOU6Telj
GBcxsRfr6HTJG7xeMD11458gEUfQ0lylPmDHmeG0i+BXPsnOhgOVDj3a8jDWlBux
hNMr5AGbgPnKf5sK+LmD7mLzj4Yf/a4qFbEEhdJT7okKfFBD25HBubjzA7qDGAA8
fn3wqyVshibnnfraH6DA8oeDd+Sq8x0HR+G4xaJMv6F7IdZ4ofVSWc35fnGXncnu
741XTb7TVT84xyM/8SiFqwCMVM2dHkwcYDKq2ufOBsNqfF8JtOz+1Wh366NyXQy4
1klHbsrda9uZnXtRDkBdmRfhKKNmnOjroP+mPieDOpDXOAWiXalZ268A9VGd583I
L2HzwyhDDa+Yyxrgjuq/QEejYVeUbeJ1zhSaKKf/fGRoBPrwhWlIzs2OIiL7b429
WD1fkT8zrEinwDv7JNkA02btDX6ajuE4NCpXNaoimCCKpRLVn8znvuV1wMma/mhz
QQCH0NokAb5FwbitFCITW8he+rGNH4jY9mN9GHH4fjpDsC96sXe8miG8D/26VKvN
M6IRs2576gGpRr2kMadd0mz/HEmvN76qZfFXpTNTiHPxdqQIAqJzG2E+qk5ytMhp
k/BKdGPXdgh6xDSDhQsSYmc0rShhea/xgsUDDEloGLkg+QDEPpvnOVzRHgdSSHAM
Q4ISJw446qLLFE1HT4yhHmxHAR+NKYl30AeRy1HlToRW08cy2eVi7YWP29JOn67D
jKx2zklUK8mPtCqEESwQKkioTJj08WjNfD+7OlH8yoGcwHFvLedCRBgcK47ZUwyY
TmwSj7NPqgRG/SMMwFTCfrL6/Z5QoJQTCeEP91qYIAt3rXoRc1MHJUCHcD+XBbDD
Nki0XuqW6vc7/Yow+HnvJT4pvnsSOYhg5v5xDR0JZiNVanz8J36YQHNMluvejZvM
ekigkYLhvyoQZiTcZ6AaOhhGd3HhmOeYkyZXXB4df2mXDMWuV6aIuXuwyIGLRk6b
yQKeXhQVFKN21KwrwiLt7g==
`protect END_PROTECTED
