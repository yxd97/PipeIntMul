`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B106DQDYbOMzqmblDhjZxDS2hyuYLsRodPdxc0YuH8Vfy3oc6jgOPhKsomZW2GSj
MzMHkJpdVSoQd44B4Q1iGoA4MhZ0nAISiY0LcOMg+MT+xKj+GWj9jpFCqD4bOmZU
AZSeirxfW6fhWNmXdM/WDja5o09pgkyAjHXxshhU8RBZO+wXTCX6Ju/EmUj9MAW6
HoGTgyhXlZpDvU75tmOSRt/N7lY2wD+Sgra2AB2PsAftm5r2Vvp4r+14A8Wi7YCh
/TpY3JBT1AiQYQbMhu2w5lEV6TpmhSyZeOShgs9q6sNr1BXlSuJCgYavbcXZDX3+
3V8GG7lJOWSsFu9+1ZmppurumoiUJSf5i/9/krq/anvVqwFbyKRoG0ATUCbHfnGe
TK439fEmZMerptUjr/iJlsN03TsV8E9NqKwL5Gkcd1MeI9dAGlOjltfZ90k4/esm
Mb8dTufE61UYL6AN7ep4PdvhJ8t5zgoRv1P7Yr3+ZANBmlX9/e4ZAGQDd0z3AmvN
fgByjlm5DJhBKLde2+on1Ds6t2fpODOy9VJnVUEgOvo6rplUs71/My62qYNi2Bsb
FRD6MyxHHEeXGkxHb03MiR5A/HBUWf/6ZzJ93DciAHME42NV6Qw1ZGzW6tCKa1kb
msvEIZCo0UQbmE/iOZaeLA==
`protect END_PROTECTED
