`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFq6t1ZFrBH1RhEFhwvWVMzKnRAp/sOKb2HEqcvn4GOjG7w2WIgO7dBGlXJRE/aS
QcNDIddrzVb7B2ZyC8opjly0ekEzrnDSvudFyrECOn08+k8n8jZ9KrArbzN76hCz
+pRYmTMTVgqQJ8AtyO9wNDFaDE/inSgrkjWv4ypY0Hf4PFbTCgon4WhNGA24gZNl
XdhXxKjqFDVRyz7nfkKrPccWANI+na0Bm/sc0HkLLSoNOhbtCvMWX89q24o0ElqE
2e2+hr0/HzYylBYmziY6UQP+Hbj7MJqs3otQp0cm6DukmZF+ltGbD5QQxvBD0FAx
gp3Y5f2/02D+K+r3frXj0pJL+lYBRhFi4gBdYQJAHu88MtALHDj5K4JZVg5+YiEF
P5cdYlT9POuHj0Fn2WDqI4GPnLO/3JpngOQM0IOb+959AnZfTYJDbwvFneDox2ij
nrNva879gYPew56LjNfyPtHOwUIRdb3IC/GLGLnurDekkeuHWgzMCEnkZvEy4wXW
CcgUSt3PYZ633H5oHW0MNXJTVagittN7q9uFBUiN201iGgaAoTeCMpFh8sd3lz6O
yDCnD2BYebYFiqipGjmo32E/Emfy9xV1xgsq8DksY5pERwk468YG6GpUieuHZQrD
d4OXV8ZfqUoXwNGo/n+p2CkLb7kj35ENOkn3ksAj1u5+EIiaCE5W1IYarL54IP83
5ojjNfDgg0bxOq541QY4SU1ysSdkFRglXtO/DMsaxOhGoHDZEO8vWRE8NnPv7ZN4
SxvYEyrQ4WpUtjeXXV7z6z9Bl/i4ptio+cOtAEDFFq9vJ7oCWD6NOTy6CNwsrtIv
q3ojBNofTZiSFRpNKmghj3S9S2m8LL5Frd6Vfv0/65t+uqxdR+i6uf5uve2Cr90p
+cuvIHy82+0e/ReCAhwRlqwpo7nhJDahO5ZeHY5xjd6K4UrPYZ6dAKfzr3FVRdHe
LH7h5MRlMJ/gKfF3rh+9Tfe1nZ2hksG3hw8DtcPiebgJ3GXQlPYvGDQo1hHn3QGB
u531ByiPCu4u4YjX49JHvwGQRX3eZvJvfkGSn5inEB0Fk39zdP4OkDE9EehsitMQ
EnS7mt/0RbG/7tiabu3xM4dOGC//9uWPFrCS6VMzfKdkkfl/TW78NTaYhdHIK8oL
n1dNw8M+HQ0CszxLxOh+nhoPmqwCtxAUGZCiFi6GiRm8FNXmdyPljBcbajbEPeuE
4tnhTSyVToVkYgLIWIW13lAgHbyf25vctflSk2LuJbKKyovCaoJS8XGIiG6AkLrr
0I1Crq1/xdD3BijRKRwTBiOAJAxUQZnjd8K8Z7ncGEaJwHtxSuyYBhEtYWJoPoRZ
aSLi18k7NYpwT5ULyYMcIsXJ4NP/WU3c7Gfn05ClwgwdgM3vqtrauBcQ4Ejp2ILR
CAMl1rdOyZBx0YB3eMHljX3UqeS/bAxHlCiPDj/Qn10/oeIlB4wWPc6uugaMKhDl
y3SZIq/GVYfHjg/JbGedO/3oc1+lskZRgmxsq/gtDEkFBSUq1ibJRhB7ux91ESPz
MKOcu5Jw+J7LU5BADU65T7hRx0gpNiTUwNlBxwQgsrS+fy18SreZOJdKpQKVcuEX
eww6NHFnDw+b+H4jynLIjxPThsQb7PuHiEAiMzDRW0tFqQg6zqTMfcVJfxul6hLW
WR6Fte70sy6oNB9DYfSq9Cn5LET1g5xXXGH+focaMN7CV5Bwr8cHddgsXYkKeKqS
ljIiOPED0Vn0htOXw6Tnoyf/rzquaw1HKky2sDcXKXjMG5C01gURCa7wBoKFc3H8
`protect END_PROTECTED
