`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMIDnwN3mjA3C8zT0pz1HkqwwNcGsWR9RNLum1I0kMStYFxgsJ6BpsoK9UvsDw+Y
MeIwozrrUAXAf6eVSgcp2uheB4HK0U/kmK4+RX2saxrB5q4OL3s2pGUb17Otoy/R
CRTjG88yD7Z1AOV0eskqjRvZkmG1rgOhA8UfvuLg7cyJlxloqDL0FTjMqtWQIVQA
axJq/4zmhc0NNJlKNco0CuaVoxhEzHvxFhuEMnK94LZMo47upowk5RK9jYZ63pep
AonQN1LpxXfjad7ElLEGnS8VYAC3kRJJu90ucdv0q5s/lq2+CbuqWn/yl/gS5Rqu
PjuRgKlBnehmhVGX1Nx2/grHQO8HctG++XfcpCzlFqqqQ9lxlEzwRbqMKICuo9Uh
ApBpTru4M5+t2yjlfr3DdahQQDs9IJE68AyFt8o7pUWEVtPDG6iAdhgc/CQEMOb9
kC0K126NxkjKrf1f0CS53ZYvKZu6AFcFqkVmIYbV4wLnv/TV3pfcLPFx3BOPdwZL
vpFSDqn3HadwpxG0UVM7d9XGNqorrjYBTctfHn13yWU2gHXlGOjHeZ2EvAxyjU6g
fwd+otm+nKjM7K9eExcMk0wUj0F/hdgU9WrC1vkMop6iBjnK1gHa05Saf/FA1MAB
Lc04R1mqw3YOuzDtYpSkc2Fg1nZZwWZXcmaWLW5vqfUSoedLbwWmZ3hrR2dY0nkd
0DTliWAOHxIGtRj7pfWBxmwVvabHVxRs1wsqkjwjcHpyiJmUXgJdbbVIfahbYTD4
eqpaEXUAvqU9qrpAYAcrokoAuRVIcWq8jhLh1I2lqtE7rMQPeD2FI+gGIGEipClQ
boxtdcSrm8/3Nm8TnK8GJJoo8U/MFpxIUu91AHlQGa8Gi7bXYVaoLqTmD2A8N2/p
m2kOvw7r6/sr4UJaygaaosnnPmnVxj0HzJeVbj6q+nT/n3eCKI2RGNbX/8+d0LU/
fr6NvSYujF4zdJZJARe/S+QwyJo4+1KCKHtsyGAVDGf7l4OniiYpg8O9U1PXnWkx
MJ/FQVtn4428Q3HXOGHHDrgtGUPlw/4w6KJAn0aA8EPkandpKbn+oc6Lnwly+iAg
PEsJSPdlnfQHxAH2qOd3+1qv0+Ne6F23AbNMFqKWnEnDHqXGLn6NZO381ViEGSY4
4nFB/g6mw9nlEL8e6l85YnZsImAh/41qBhChuxyhL1rmkIC+SypdOmM8Pjbkc5l1
8w9WguYJ5stpKx60SZvLXsnUbWkfPx8eHZf+tsHJmw8pA8YrINc7HHqrxDCF7T2h
FAmMM75KO/j4LeDvxkK7fBFySfql5xHFWB6PUMxA7zo+dP0O7cSmMNrViAIryrhG
NXnSRQdtAxdcZFkFmXfUBkjE1lKBj4/zLEYqZBpWq4Of9KwLPw3IE6ohHTKV203c
djYOVJxtAA3Gs/KbVzi33xVs6D+azBBZwEgwtqYSfCOwtahBFqCjo58Q+ZTaDUAN
ZZ0nih5I8+rKCLK1tKdOT4+8heZrxnS3l+SjVpvAMmP+WN6Vm8aXKtM/p2QqAKws
HF0yEtmxVHuCxSmBQ/dMllv0NkzAlua8X+IUqOI694y0MqvlJB8pnWEQjm2VlSuu
8wi+3joYjqxYyrua5pgkdvLTm48OwS9BQBP0YRwF3IdtA9IsmEPrPNXaP7/ctTkT
h6IGLd64D3GOhgKZKij2EQeurujNrXu+WcctKSWBtcVFi+zg8TyFaz87Tm8FABqz
J5D1azUhfWdqI+tKCTHrV20+gr/VzG8lmGDvCFxqeVx5EVQ6DNYjPEawHUn9JSwy
Gfq+WEzfETo082t7rCedo6Aj/uBwHnLRE7ZnFD5fzNRpFVsFAF2YHHhr7DhG/Tab
r3hZz0jyKDpM87CB0+51OCfarvrTzkm2sqEm8czXrEbNbt4RYQSxggA0yv5apX4X
x74Gm5A71GN6W+OLB/NTHkOKQbREH1rNjZRSio+J1s0skZuiWQ42J2rcmLAEcZKF
ooLqBmXlVvdZ/OyNVjIQjTbZkouZDgYf7/OKZO6abJhMoZ30Ekxkxi0glGJF+r3u
RemSQXafVBySiZIQuYJfqJ7JkJjDwcvNlDx+NlF4P/F0BC1FO17bGAdhrpL548Cb
S2gh1KW3APxWUkxNY15p/ntQ+RjKZliwqUXZy32pz4SqHcZa76s92Qinv4bN28If
YndmTCOjgWPunpR+c39YRC/Z5fEUDsBbj1uqBy4Ji0wdiN2OhjxrnqqvIxmLplk+
KcQj0Lyw7scvzIr7zXwYGFgNeESbEIheZeqJk0RIe652BD9C79cqIMpCb7RVzrT+
Ce24voEYYJoAceeIaVpB2ORQPfkIC37+G+tjYpxHGq6DvrVJRu4TA8iFzq+PPZcL
/kilE4AMVc8mZ559+xmxLUYf5DbYoIJIQCRfDJ1FwdyEDkZbcwEI1va2Hj9n0x8W
V7E2VgZ7V248kSIi2X+BsXfn0KafCt3ZgODXaK6eB1m+1RWgsTjLkMfGBHc4mm3/
IfNtc5UD5KigMR04D7yk8smu4UzTf/dEOF55WpTGwGZAC8MKfIg68ppRK63iEEHc
PV9TyqQfk5LjgeXq8pqzbkewWuIkXhOEqOxCGfV6FKaOOL5thumpq+jh1lKVlFA5
z34aKPzJthcXRb5zvQqYbiTQayHoRQxAuiXDG+5J+36QZaqje33Jt/1H/leers0n
04FzKciAcgp6aqyfQ4zVlxBPjSrdPBOtjb9e3iSS9W7pjnj8hve4muQu6K+XWA6x
TITm0MYLKjqmx9lZsuGpY9i8m8b3RRl3x4p6n+FRo08/HupDTd5Nqxu3ncD2zMs1
m5VDxvUbECAswKoKWpsZxz7ocmvaOTr/V6SenLGIB5p6l6Hr3dg4NdxR7BuO1+66
VzVy9JJZkft6ItVUzjCuS0Xq2qcUT1K8yiJaBUAbMfrMWVrR17ompFWZfek6D9tJ
nZ2m2siJMRq/yH2sV1je40CrwMhkMNp92LHYTqMtN6A6JwKzIS86aToyXJ1qrJG5
nC84hUnfQhxySTcF3FUXKV0x0Ob4iECMyCMoU5ZAafrSWzuqnnZU68MJHv6rJWVo
v/G7l6wKAjTKuMSpSaxO3GcY+y3C1TKvyLyjyCVyzR/yJJB1r8njWa5UZWvxKznE
6wfofx65+5uPyj126QzadKhOvA1cul+KS9ydZgQTrBweOHvYi+IlinQnp+E4XDbS
7XjcNqMAv0JzAW6VeEttXZ5yroCHMhJtADKy7jUiAILkOScSFl3G0/zi11rPOB9i
fCmY9kjNrvvgLHimlOtXKHO8YubSJUPeTVPLfLUgPLVgew0tF1NmBQCoHXQ/469E
rUXadSeiF/AfkDywOnaUGRyRk3bQbie/fC3LEfVvvR2DKf06+AJReVGSKwIFBxOR
i7BxRspz8cW99MQX/gbogenbBfpTNskHsiCwYAUqToCnRSz1+loH/P+rYwNPn582
61P/moSGpLuUmEDwALsqSUA3JrXN9O5THV6R4SRHDYzavL+6QAqjjsebXlZXFsa1
vzcRCTZ1IGSdczWtRq7dHZmVMAernOlxF+O9XaJfyVzRIGR9zRj6ompaNyC4dEdI
AmEvKA+vl4ebwd5E7zcqEQC8YQPNqbMdoglnGWc9zBS7VOt1mfFD1VonYYiLRupu
2mwaV3d+ZrrHz0jB5+x6GH78arOATdGqoI9Z/t28sb7VuErG6Q6ym/pg3epg+477
BCgMh749FvpVE+hnMZOmCPePdvzcLnDaynhPaahr4nN0ylcejbNIhqJnZtr51WUy
2OCi30OrZGVg9cxkdfpiXg3JJY57yr8CaK/6Zj4+ELujAKX9ETKGa2xm4knzl45A
9lMsLYKVF8FRYiSTNF0SbP+j7C4aMUW4Rt/GCdJNDpE+7SHKyD+io2Vx9Dw5KX7i
xHnQaqVOEf5EnzKGnWmntznUcWARPLKbqvLaW47Ybd2VmgfLD2v0cKowE2yWx5tN
QBOi08msd5/sxYRRyTzI1Uk3XqeBBrlOd5LI7XbWOhlbq+iuqJHvraFqx8mQV4rI
kI23tMhLU9C46d8pnJzU2hu/INMOR+MMpf5PbcDIJ7DF9asD8QG1e/tpsEv7Jd44
G27RYV0zNGnLvyE6KhLk+iwQ0t1gM1cmY0pWtZ3XUYoN/hUFHHt7jiNDnm9JnloO
3XnWPhpwNHRMJMQ2PF+UfWUSB7QNojTsqUNC1t9AYbmFHB+bcuXrweOTzuLeYJ3F
BBFE72+bhd5kRF0lC1oeDZs/4pe4wO6k6Tj02ehKVfqF8FAw0oe2Yov7ovTWnL42
VdNA5mevte1x9WSBeC1F3SOCKU4qmXPhqNzSA/HoEQZKo3rc2eCQvU62TlEi1zwe
9ckZ/yQk4WTXIXejVXrYp3/k0JAv2hxNM7B1nAfAmODTpg00x3K65XIkV3ckt2UJ
zkKtWB9LhLDFM8opdWMytZMAW28nBpStl7scYONSECETHhLdSrZFHf+LLPU55/Eo
btvhtsz98+oDXB6IWhc9Ze2VWf1EPWy2JEIOcYc7i8LKUjmowoXqpm68JzW5iD4Q
+d3xEmFBGOrwbY1I09r1vqI6kO7hyq4DVuOp7FnypnMQuUZpCbc5B56rpoemZoNK
IKHpgrEt5Z4y2wAVNNcQMeIgfxY+C4z2dwZdHnEhhZbvqG4PIqtJ+T8SNJtIY9HU
x6G22BeD4LZU5DMy2wpu2glVraC7Qje/Qj/D5GfqwgCgOofy7e+PrJQ97Uoj7OyU
liEuNlcuFRlM1Gu9/DLnzOWbvHfh+9Up1PirIvrYKT2PGeNvwVK+p68fgWKTOlsI
perXopBo613WJKs1egDfbzaQekNIeO7y0830QonMAfTihWw6R99Ia/tsRpyuLAVM
Pk7LAk4sq5SgoOBG2JVvYoAbocgnXnXGVkTKTQZMLq+gF3CSmozjC7tZYZ8Iwf93
1znBeT/9CTR0etH5QYupt23IP8Ud7zA8sk55R+50CtMZ34lDqIqaKzh7FOrhR+Vx
MdzJW4pUFt01dmrSlB8BYkIsBiUIC5dgQhxbCVwcQOLMD9pE32Qff5qogL2Rx6u0
zEwe/qYahX71Np63ls6FmhWa9hPuX3QxqYDIJBpS33VHYNiqOxyNW3ukPg2QplsK
5jXORLrdbg9uz/Wmic3rKtmhVfPV8KSOEozV1U/ewSOyPwgkpaz0i/SqbJZIuKcl
mWz88ZaKLsGBCgnvzHsmoNgSN612zItMhqZPPPE2Z+uH4w9G1/91l+CnPQR+SDFK
mTtOEOUtEhgOIV4yjFUkpK6BJOFFMYUjO331JordfibEq9NAk5tif+ah7cPe1m07
3aXlMCLX8vRRcI2gn4V3XPq3AU4HdKYL1Kn6IqOG2jwbyrUvrjYXjFT7wjZqsz25
kIEKj8WtrL+GPM/W2i11+gEjcLPsqTQfKmC/CuUtyK4HEKqRKkt0f/rrbTExLJQL
qER5+1DXP3DaPFspMe7svoK4UTk5/2ti167eWvqRzv1+Sd2Cmo7TabNMNUeHX75u
WbXUNRShUcdHF0ZHAd61+Uv2o6S8wsTLN6bEODtDY240zlWZiV/P3rphJ+mNyQT9
2FmXMxMVNIuKHohWUcaOlhqt3kPL+71xRxi1FAyrqDyw2XR3aavjpNcx+nMJTZeL
AWwxX5fSr9J/41OnbXuBjsjY9C4FfBAKb1daYqWPrbR5V6UGA1B8USrGeTu5PyLe
tMDDtBFQ/vaQvxcNWeRAozDIIMHICXsJlSPcVVRIPeNI60v/g84RatoXJDJpP8EI
92JXAAI7JersoRuNeyOrkAr+hHuI2/Y5r89sljiIZkFhFhhwafIHZCJl1Z4znHg/
S6Qz9AEwIdyHlpyAIGcxoypSEw38znvXWVphKzJWldJKMASObxoZY8QkDK7dCi7i
okQ02Vq85RT3jy+d1BePO0IQJ94gIE4Zw88odsW5uv6aLekfRsLBRA+d6tpccwO8
9LLZJyYugEV20toUDrNrpf2aUSAwHbfZbbEBWJHtnwbFNctmtVMmf8sc3xmYmlTV
82H7ImVkyFAqrh41oUZ+y1iH1B1da96b/8O0yA5U3t0jN6LpcbSg7ehwLRM2EiHc
USThh7mSFUQIaLmKYjEavFwxbXlluazGEtdOcSJadJysPeTQNbZUq4KAZdmb0MX7
taO3C0ZQtgMrdAV6ALIjaHrDCD3RQ0W6rnxtXFRQHvtdU2E0zAQKNQXE0HQSqMz/
ODfK1urVuYKRIDCt5q5ccLXOdZnMMI60OiNIEVCOcPM4RtADyRVeCY7h5O2CxUpA
A2wvvsV95YSaicbzZA8wgACvJ1Xsp87wMuf99xdQ6Qv7Yg3NatkBPp3kHVTmS8eO
GS5MOFiTpySEoeyH3d2yn+ixCeIC6LR9kwFgyNz8zJ5MCdZUhALs2MbpJ4PmSBKR
wke2ELASzakY1Bgzb4Xcu85R2fVxm0yFwcYRykQsTn9hGPFSw/WL6F6S23RlXgkl
xLZx/vqurulwhIO34KOTy0zMvMeLJcdw5abrRl2Th41ZH6KSbwvTIQojM6UEM6Pf
jEii0IefQuF3EkYDftnNo1kJOZ5VhP7MdR2r9hNjjElH/y788w3duv2uVTi6LRIM
ObsAHUKZnlxD3MymHtH17ADUyN8vo5dcSRHVGDS7C44NTrCfiAI12o5S1zJdWO+l
qNJiR+J4LFvsLAkZEFFyuZDlNEX6p1yv21H/3Xf6IJDWJIOyzUAV8Xo3KdgrRAEU
aysJqvxFMXEGsctoDUdkOHZI6G+UyUa4qXj+xIcD1TkiwSKnBRZ/6GJZq0IKJT8q
PELfFhmEoMTvIAfivWVaoHwwwT8VP6mycBSITtLoPm5ucnfEmFC27gHl1Ryg6+Bt
8RNIhmsSTWS8QBqzm6+SxGKT59SAhnF0hLAkpUACNRGAFz1b+DleevZ8Y26INhQL
zdgDlE+IFvhnsx624I6XpXo/gyjpXFolssCqfDyJBtNABTszb3AG8oQhdN1R/Ms3
OQbx7nJoO++xbrWVWTNsvRgtwGPq7Wfb9YjTS1/ahsnc6pTZ6IiCZy/sNeNXZoTR
ms9kHtSA/Q3F3SA8STbMagbxYPLA5zzhwXZxAbxN3GNacYOvUKa2g3SBJ5R0WLsL
X0lznZlCKXncsMmPr//wVSC8dLShYJQr/Jp5Dqn77CNZQRdn57VAOCZZEScnucB4
sXxA2DqcgEphQF+sEd1ZrfBj4s7mFVNqHnai1hPg/yVDkR0lDmt8ktBHYmoJh8Ua
erIcZIVb3a1rdx2ugiLpnG0rQXvMk0K7sQsJyETVANqdstIQxXaajO7/DHEVWs5Z
C5MO6Na2s1vXB9twW2+hgAKSTy9XeQfkeJZ/31iSqhnMX5vNj1KIcKSOZBEIgyCj
gOxSH69kXX/OFuvCCUsHbmkOj8W4GokjsgIAjaknqffscFpmQKP6dk24qE+x3Hwt
fb9zzAY9NeXPSUz1hYRYasHS5wHaS+EtJqdAIYBFujH4BqQNOKXlT0uchKFkWbNC
/h+53N8AyiS8qg0CclHLXMwI3rSa7pGotwnjQ0pFw73sLg3wabOdH2rKDTcQA9tS
bqE4um9bCuQmhm7VdnNY+V66B5AHhcne0Vhzw+wWdhCGQck/bpfKR1EIZIE9ROQY
/fE8AlQYqpSgDrtaxPTWCtsb8dSoyrR5WmGYIKrvutCkd6YnujJH+4ET628Acd1R
fUqKeMIegF3cquGQfblACxcopj5LyE5DvnxUZh9/U3qv7pzevyYk3A0r36fG+7PL
6ud5R5Qgyx0jOzoO/fXEo4uZmYwCcKSDu3+7U59NijnJrOK8kzd2O61V2fclgjuZ
R1PGf9POUy3EX1/w+RC6l8k0nHsNid/K0jrDnPZN1seyXQtkt3xuL7vZMz4dB3u1
fSExa5JChrJnB8wxgNJlvfjOJ979csPeaMuXGeS941fu9uP9lKKVkrypfdgJO12Y
hQ8eJs6G1FHlvjd/f6m5gC8yc095Q1ORUE/OUNmUOwfIusoE4/K+XF+ma16tqJuR
jLUfcztAWNrfRvi79mYCty7TOWmm8mGE6GC9OunQ1ZxXOje0aobtG5ivXt+/wgW0
eDDXjpbpXgBZhr+pEclYuw900o33jcw0ZH2ouX7Dv3VgXAeCwBJPiJz1TSDRUDzq
LHqo/rELlm7/kXvNVLmyCIVv+BkfkoBLX4ITWUx0LcIG+IJYOK0o2OI8kjjQFarL
QVvPO+3IKYSq2OHiFgEwCKaXIGm42pBfV5ka5F5LvsgDeRMRnUIez+gGqA+H+HsR
i1AhRdR9kVWfrJUo1J0x9rBwnlmew6UPU46vl8e0XjEE9qHvJWxa35d7k+mtty+a
v9tSvsv/NCEXrzh7hy6wN6I7sebwLEpZG31N+Qyis5ZIDOuAlZhMkniNvM7cDvf1
/GfwEunZ5MSNd/JXR49vkrnr7OPyVBe+Fd2bekl5lst0dhvOBYJk1tk7XxTVA7dJ
4dM4RXIeSkVfHn5RxqLJ2tz0+Vx7MPwMGcqUQVb0f9fAaZtGAkalXCHIOExdxahE
WVr++z6OD2UX4MUruCf5b/DBAvk5iY70FiMqjMoGxMCoIGc4fOLtlCeq/9oWfnqj
dAu32sr+bF8nLTp/I3eyG1ljtOVyPkH+mUKywY4tj+gzbRUA2u5773l/hkZcG9ed
S6MzLs92RxWKzL50fUFiHJHDPxXzpCYIChqgCv6Tt6UVM1MonKow3YO06GwBmop7
YSgoacyXVNR9d5qh1RKFb7WDfxf3+HHPdic8+CQBgUCd0qXQFuo96TWZFbMLmm2A
32W/J7Iw8LVeZ++Vj2tI39ZBKm+UQh8W/SQCFf/IY4JMIxpKG/hMLDtl6rPFizoj
pU8YyZGBxOrF29CMnqwr3vZujs0IUJ32BEI8fLzgrEXXjxgcaHxcBEhcJBiKgggy
8ZSVe6b8+8+d4L8XK5Kt/zmt5Lv57mrhlV9nPrkEjTy5knvhL9gMTjyMd9H7GhvP
aFyPwmHR7HJEiHoKiOdXXyCJP6pYHNv3Fh4ovlJuM968Pb1QRasT7xoqv+gFtVC4
SMFqcTWgTcCYzHoHhzuYmDe6Gu9/9pdRUxNJKBCwV5tu427uSHCnC7LvD1avlm/v
e2MtpFgrZDsjgpMcQCTbwR4NxVywudDo3FSScI7tfIbPG3QYYhQQo99YEaLM1Nl6
Zg1jAhQxuy8zxWvUqZu4eyaqw4STg0ACg/wSw3oQpO6CduwsUXFpvCquaoEGLMvC
wTIetuguleBEq5xFQklQ0r+gWi3+v2A0H7JyQz6/md9evJJZfy72nwuUZwqYG55t
BPLDCisug/vvEtxmr9AXurj5KZYUBo59TTIjAVOlr81mQL7O3LlPvxpp6H2nfxsU
LWsQzGCLVHsKAT2CbEDd+kU4YpZp92IWMZa6M0ySvgv+rZ/2gtyeszkrQEXu7Ihw
/WB/Wp8fKj19IIMO7sK83snaKggdlZVBb9hLiUJCJeVQsm6kY8Ax83Qbpbj8W6s2
9P1oJ0luSQ3/10VGLKYswFWoWJdGuw0YJ2pyFll5LTcmcnmX2v86xTdqSA5axhcZ
qSWXHD8F0VjhDqLLciZWoUD8xB4Dc8+aNg0zcTDqFvKAw90AQmeRtOF06xwmzwqH
fhroT6JRIKmn3TVNqIPEx7roZp+ntQR1s5fu8xYXr9pDsq7WGicy9xMk6/ru+Mw2
IcQIszYt9h+FmeIuGJ46dm1yssdAA0xpsq3SRaFsMYX5namEBlGBTfYNB2Tp8aah
1p8ZEVJ1DSRXzks0fGiyY7JiH6Q4rV+zmJOp0LMGn0kTuWmTJ2dkTZan2HqVcCIl
PPXwy0OV+J7ZM5A1cwL1DFNKQgPZdULejAqyk8ETGlufMecSdfJblW5ac0BWv3el
bokpooc1Xuqe60XfasXLkL6Xc70D3DRDpA6ptFGkH6uNM38n6iP3a4+uQWk9oQL0
egVsXgY7WN/wP7K2jk9z1s06DerrKY4kj/kRvhAQ7aogPfrLLb/PX13DTqbImNch
FswRcuWtBw7sxok2SH0G3DoiQ5jxyhHUifCbTFpEGZ8XzRiHpL3P7nc9ythH6dnY
dTL3TxOO0Atkad9yPYsCt1exdDx1dIALh/sux703ON3ql8nMyBGVPWZvZqIZDLiP
Bt2zOoVCREF0oIEQH1ERV6wdjm+06SB0lnyH0nPv9DApnGYaFIhJBY9JwdeUo97K
PvY0vQFphQ00lYJomgHoZLfGyjvGw1NDG632cKFCilpnMMkeVmxT648n3O1AjyXx
5tYnHiSfoISK9yNbx+LxZkRCVgjjlBGk69qdQGef6nYrKXE/Jevsglt+BCpUQi2j
2L0YHrBaoU5AK+v1oW2ad41sC5vbcnP4GloZ5PyQ5fcSQ5oexVlO7JafctQ6k5JH
xt/qIfgUH0JrP9YJv/40EngUKqmvwC0+j6dZQxKVKU1pd8yZyj0RFyncultbYtoh
7A4ZBlFvwQJxOud3bhpGJ2uwBLbQiWhhtV8aUuYnjzsoljfkqWb/qByrnCDmF2DY
xT+v31GXJI32QRjVuAE0G6fV5V/NePFAPtEFHXoleRKrxkYo+7X8QT2he34zZy+b
a0Wh6y80lgfZeR6OCoQWLK0cG0Kf0qHS1AYVlzgHASsLTDvudsuA7kxRZdqf30gI
dyB2XxnFXb1h+M4z6QWqj9bZG0VF6s5YugBW79syUlXX1MbN2ga3xOJ+VyR6uR/P
W47N8littJDZRgX7perJpdIyBPT2ZDxzFSVDISN3ftSNwCt62PMvQwx342TrnWjE
DXoN9izeSV3LThJdnt+Umz+e/FtuKj7oYf5XGWoXpdQuCoj4wpMhZn9bqcuX79pA
lDAkRwgvkmBuCtLhxoHLjX8iR05qG6Pd3pzPwnZFiigKJbox8kVJFl7+YJbghjx4
jX8GWlQFhmoKSm3sbAZz77eVtxGgocGelk1rx8TS1PeEuPe3pgg0Keh3uSO6hH4z
w/8T5Pw9qxSQoNK8VACFkaXxO1QvKNfs1mC/7TBsZUdTHVquwtbu3cTgS8qQMq0F
Qedm8A0rexP4oCw2VldOLY3srEHWM6r/yRnOXrWENmcE0Mxa8K9ahRGg8KVLczWT
NWSFUMpZ8x57toIr5qmFbGVcgH/dV89JPvSop2GPh4M3QH9oCsQdT7zwLbpYW1mz
VBwwg7ypsVfGi1rAaxRjKpArVG4B67J6KIaYG11pNKWYNtW/gccYz9mAW/buRoLQ
3QVqY1m/FYPSGMMnhxHYISlf4zZ1bvCZuNg0TFtxiX7kOT/49Hvv5MNLcNPb9+6Y
B9o3wvk4e5jthyo28IOk4ByXue3oKsRcIS4qOaLpa0vNph5mYXGvxshVpgBXFNJw
ccFOl9ft1tSP0iBNGA5sQ2SMqgZgK6CbrrjrxBgCUUeDpVZxANw82nqw5J08Oe1p
UWYlirzmhdF9V21D1XolhGYgMciB+PH7KbB7lmS3Q1fY23uFfLS/raePyhkOKG0t
ZrfCySt4Q7PmJXraNwLHz8hI1x89zxYaQYUvn//sPIyCFos5N3j8zlX+2Tssm6dU
qUDY4YCm6EPiqp4VwyRUGHqFussLE9bEGOdwo5r33kNq5QArqSMpK2ZKghj9OtK5
bhk4XKBAxsyekXBAJ+uTyqNyK5yKkAeBnqEDZrju4NvhW5FOb5HLvGraWLyN6ooN
VqRl/XTlqnL4OefVCIMy8/Vbk6DrS7sQ+9rSE2+gPMhKIDRu0jb/X6uEmP7txHd0
Sky+owILNoVPG++V3o5b7gbPUJJT7FXmIdG0pUbmWYhFDh7PWH6AzFw68AqMD7P6
Z4tkzMtsCwq7Mx9tHDPSLW2Jp63BpPy8GzTAa637EAxVyXyljDrE4ZgF/Ge8TUqy
3Rj+cWEuJkSy1k7oQFRQHBzg3XMmNmc0yO3BkF5WVi1aj+mo3LPn3KWdBIgBbtCZ
imuRTggfQXJoEENlu3bZisvD+o6Y1+FBW9gjjPyEn115luTDVXjczsVxLrcsYiRu
fn403cxzUeOS1ivwwJ65qBgip0Itoc19PHwddgvGBy9sIslA4yIu5xHBwZfTuIjT
V1DI+auJ665YyBM1IVlCm4/378Ntp8G1IRTQwsTXw1c6WSQqRzsO6rX0+DseJMne
UF3/1d9VgXf/thMdC8sApRr/9RWwKlkXMA8AC9OWZ8W3qixK9ByrQJ6X4mwyNfs4
oV7kAJ3PbIXe6eJxkLOiI20abm5tsIsiG6E4OtUziTsqN8wxkaAMBQ1GfruUzVyk
bJasDRrOJ0uEd9BgBMkiXt+STIskMA4hYOlBcZDQKhr+D/zMlWqvHz3ZehBRenHE
bOT/w7AofJwCOZk5akZdCr5FlzPSbJC8vWYbZhvXfZ01nq38Ji7eL6mgkC/WelFV
JWNkRioEJL5XDzGKWc5/CE3+cYTrvK9gCPPah340YPoxjzJYUpJ2KiQC6OYZqfkh
7DS2rjLcR6bh4b3EOozb0izdzceLLFHzWxX/o8Labb/aQ8KN8JhabmTkCdFPnpDd
2NXsevb0jd1asUwf2+/IayI3GaFb9fAqP0ZILFBDFBVHpvzYscRIW5SxyApFx8Wj
0hq+R0ALm4rVHbDuE8WxylBI7GVqqA7rV5U9YkVXTytlgeAnFSEl3t9UFCfZAxTQ
jDjHjkwO3AKtP+cqxRRkBFlJOhdsVqBFPwdWMAo1cVjJ5z9kY9fvvpe8oAOGA3J8
jP2kpiZzP790hT/2zx8xZT37j6fT3g5HPm36rdlTKSk0NgCKMdHVVisVLWkrf6kq
hRTAl+MkU3Vr+1jLGSE7hqYjsTnsxDCX9OF2xOJG57FA8iU/QXs+ASDnU4Szmh3d
m+x39kyJQF1rw8ZOHauBrSmyhHOi/dX/bN4YlBqFVRpMrpKsDqBOkNo2n/9JMsX+
mK33TBchOOFhpQNGcq4SDAZuIoZNQGdzE9VzfIic/hWEjvWweh8/WZc2YnTHQ6NX
Bl/nSJCkfWOKzTmuNdCwLR/q2E2xzXbhzrsUAWep+quucra3Amx8hyHd8Re+dgdY
8MzuWEU61oGs+uaU2CverQASEpntsEgZAlslwc7rwQEBMZarc22ucDJfjK/rHs2g
YSNYhpgyaaBpw4kJa05PS4XoDoF01rYCu+IPp1h8IIcfXAg/U1WSVd6Pzr9L5bkE
NvUpXv4ouDZ1hzpTNFAM07MHPBVLq6NdZe0FEu2Cu4fRrYQVYu3hYIBCI0J5a65+
`protect END_PROTECTED
