`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r296bnosz8w8c+xUUFfMDp5F6Mn/t+LFTcDUJ56UfgsRIjCkJ9uU8DRStjEvtDxl
w2twkHGqG3Egz3kqefJrZjYpoNSz2Elw1sGFaxYq9uRQBY2HZGRptcDZhDt7m0wH
3KhPw0ym1OahnwlumixBEgUAOYhj0UH6WmvxMh/HOGu1IpPLA5sxbsrNBt9CM1eo
8bEp0wtZAZbZ/tPlFee3NR6FVKoKophrUlAU5FP0yM6QLkDvuK4tBbl8jyl9AZqy
SZW5v68J4jBSjWjR1mu61+wJieNz4V6jUnxqPY2zhbE+PQ0h/WXURBo6fYbFR14A
o0OMZyYho0Mr+dYwtBXgB0RtftuLx0lz5hraH93hWUHD3qxkF+3OejVOH5vk3V9m
/UOfXmxBDZLx0yRoWIeJn4YHEoAMxl6tq2p06S12JK0UXwCwAP38bx96j1py3AqC
7KvY+oxVET+NdZ7lzT3mnHua1FNkakls62KAGFwPhQjTDM9GBT5VAwUARCwJwIjz
Dxij4YYIVvn29p0Dzc9V3YDr8cbTBe2r4ywSaxsLdHwjRsTySweeEGm48JI8UWfI
lSFt/7AyPPYHygS7ky4JAbVRJnnnXx4K1fRZts7wdRC2mnKnfolTXzv9i0J6fdFU
tjjbCgNeB08oqQ8MuGI04I6AS/Wg2HLts6EwGcnW60aX22ckb/9MNsAXLG8C1Q8S
Me+PiD9IHdrCYmZJpZ8bstF9wgSaH6sloXc6UTVjggNZFVeC/6H7iyPAgubKCfNO
QJvBh1enyHxlA6bkjtncQjLEwPDKJARCo+yMElk4NST5GM9JszT2T7Ie1YChxQ9V
BH8VLHB2WpXaYcaVojJlVEWvKiYr4bcorCX3WvezaMMuCJ7s53FQesIoPlvK0PBq
INDHwDiKCgBcEdgm7cQJgYg9JOlVUzxWfQTI7o7AWWi9URynK2D7kxHDiwPfjra2
8NOFvpITS9b6o+e1qAh6FeVvuz7TdtyR4lLb5zl/GEE4Ofn2ZbQBkkXPvDGstALY
bMdhw6xVNb/d2iFQWgdTuCaKLx5UpdyoQA33Cxm0KkHnVEq46H6ZOp+09V/xeFDj
CwydE1BWxaNmPlmoje/iRrneeTi8Avag4IXRxLvXG+RTz/RV+6C6ePZWcxgHQfO3
QY30JTNo9C89dv21YboKSVFw1I3KU2/H4pK7GMsxcS/9oKwlpgAdgwiU9G7rnugx
5AmWAltxE04e8iwEax4h9d6I44ie10zeWDWz9rh4HuyZOq0caxzg3aiEHRnIElJm
wzBl8GDE76z3lpbKvpHKiODhJOVe6/Lxum5EVzxHXRJZLTsTsa6o239wu+4I6+BA
eKquKAdA888uvikA49Muf4x3WMTgG53uiv9+kRbQkLZOO/tsyMB/ZEYVLiwkWGHs
aU2C1LD5s+SYSTqi+yztZJIRSTYPKcEMPEoTh61AshQPTJRuAVr4IzREyXLgx1ap
jmo7RrWk0dmCL67dsBXqG6vp+QAmeGc43NDP3EPFLIF6pxbiFF4ORrSCdiQhxGD0
2W+SFg0caAwo8HWo158u/rm0G1Cwg+8FApCXUUohd53ozkCwac/4jZaX5C7lxwpm
JadmdGUOy20o1yZ8mksBp7kSN+VqNX4ZzETVCZGUX9kippR16merN5NGMmLKLdRH
n5DTLlNb+zWkF2TOub/Caph6A+byjtE1EyiWvkRtJjeuZ7pNjkdQnRbs0qc+c3Wh
Lraggh30btA2jV/uM6coyLXRq4R6mUxsau14P/b/nKky8UHWn9vdS7kqvhUE5e5m
L7S2eRlJHiULa0ZcMlZRVscqGBShyphJzyCHM7gcgjV1RkuhrOq/EzXIZPAgRTIw
MDZybb4fgClPj6PnWiSV7K4jo49nivCWFANcizJIcT65N8k4hOJ3r0noKjhboFYf
2mjVN6KyHeO9d0cdxH72KmlQ0b02goymWhAYTbvQr+PieVTe/3ARYToyNaYV7HVF
8Y1Ffe8A6oN3ZvRAt5/42iV77dU3358QxYziPKv4n5s9pAvTBdDIf36wilTwi/aW
aDXwllgpYujURWP49cg0vYcJkA7wqAV5tiCbL6eiPCcJuhdY5wSESKu68n/yMVCp
xr2XSRdy3LerYBFoClTOaMLbmc4OTRvuSf5TP6z45Pj/2LNIrZrIN69hewuaB7y9
bqCBf47d94k+2/4HQ8143mZr2nrU2iZB2oI4pYKYntnIKQxYg9b4Xm+tLGwdZLfw
9SuS2LkXhhIwUVJRrioG+XK4xxC834cIErdyQtyw8AblAvXsdkpndN/p8q6Dl0YI
zfP4sDAj0GQpzxKKjyGgfxarxdc+MsN3BTx6eJ4SYffycdMWecCeXlCgP4d0+17I
Dt9go//chugX+B9T/UnoTO45a0Ug3+s3I1SU46xDIKZXN6u60t6QyuUapCjPtHvE
Sx0LzJEtPvDqj6wxstBtLYnTkRp2cS8a6Ttdtz2N8qY0yzZOdRTASfkouXgMckdj
D4YoftVkEurjIVS4NavceFlw2lac7I91s8NnOTRP7pBe3DphTXnwc6rTIJSQXY6j
Xi+/1KMdQ5jv7BrXazmTAYhkSD5/HRYCda5CotMA+RX61W+9wX+Go534RGjyxExf
3HUCPxF7qNJhiq0KDeFybveXuSLcTCYJJV5AaF9BaaOxUyN9qlO8+zABRM5uArYx
hPBjCXnniXhdaCMFvXZvpyjihc7kGM+5hK894g7B95FLdvjYBkxqwvmrTSnW/awp
Vmca3kw52FXyCI5j7oAIsef2f/v2Bx9b5FYnMMCO4HYXi1DU7aIaYA2152RH0DUf
/L5PVp8oQwp3gP/QzK3hb4wE8OUU1KUURSKKxBCxol98lmoVNyq8QFipO8Dr2Me2
IJjHOt+PXwKOHXPP3aMYyGyClF9wleWcnhiK71212e3iF5/vTFSS33VBKfP6fhlK
qRFZ4fgfkWfhNcoxFUMMm+TCMgb0ggH2WdAACReViZiNKY81SqRwOLVIzsf2w2T7
iPJc9OW9JBWMOEkqme9hDWZFAseMy7l35X0tHSXS4hAphpHeoa+h/oAcY1RbIWAO
OYXOQ4HDbxtVkaK5TD7L0X6viutlx/wq52mEVwajb2ZxCTecTWY6NBkJGjQ2/2CU
DlKkJHMbPAtkuE47ptK1h7J6wFFUWaDXG0iCzP+sn3qBxpZIyAxGNlzHHG5EJwZb
e0Ta8uI2WzAH6tsZfNQADAOvn87HAAkCI7W5h5I4Q8pr175kbwCq1tqvazoZEBRa
2y/9uVi0BrghQXXJE8qx8NWadEUVJMfF41lZ+EsgVdNGGy88N2pDQnXxKWxSzRB8
6TlhMXdFGGra1rkDSRfkAbTLWe3twMB1htVc13JnLYnQ0q8YxSIqiiztSO24Sc+H
iAoEG/0zrW0ErGXxq0cgadypbrWhHiOek0BFD8psKXPqpnZPuPTHISerm0pouuSR
rPWMmr4dFKkx22aOu6EfOFIngisUfxNhlV+1PgFxw8GQfCVhdnYixXc1RBhDOJdV
PK5F13Fdw/ZdWM07jdcw+5DcPHKr1uPrERxMBQpoo99ohGD7QSTMIBagDsLSE7B+
DHEd4z1VxS83EENOYqHppoVvFT1zZn/1BygojzNtnlN2dMEnw1gKRpKRe1bbfLRm
E/gnBU2l4lSdTeDooig/WOgaEqURXvLfAb1OSPYdVq00xpBYMocrPoN4q2mY/vs/
el/4Ov3sEeksLBNQV5eqTzyB0gL9cBLI4S5IS7gTEdDlMnMmsYb1/1UHE/kUxOMz
EeSq0eEVN67JiYwF//0AtuUSRbTDKHNZPtuA+Y9E+3cAYvwCjW2n+YKicGJ/L+ri
Fhf8DYFeOgTpeTfgv0m1WKkL8jojI3+DoRA30ayeFho=
`protect END_PROTECTED
