`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jg3KNBw0W7h4G8GWUtJiQa7RoXyZyTBzNgMfx/XTjOxPrPwS7o5aaYrE3eP5kjjU
Td4BJtVhYgyD0faAYzqR1wr5rINZ3zE0MTD+uI0caAEPPoOBJ3RfEJzhTs8EBb68
mtfMHN4OSIBQeY8HNjQSdeju+2BISIBGOL+wHYq/bsfpmYGxAzivVpRJ2GaWc2AQ
9arKfD1I1ov1GlD2l9DucmMN2hEb1dqzdG5tsjE7C2oMYWaOEJ/4nuaP1NSLXEP7
yV1eDkldMNx9gHxuWsa41fyvrbPFqHK2NlkAcaOhakw+zt9b9MmQB46t8Tag3p81
k8Gqhzq5tbO7VoZyrhNAwkI3lKG6wLqZV4SAvwEZuHbj7K3QARC9yDLn7/vH3zx8
lJgS2AHnz1LTxbNd54sgGdmjmivXE5dsKbgJzkSDL5A3aw1feYfiTCNdUm+7fRvW
Ny7cgLcTm0RibfJtNz+e8oJugs0KRrU8CBBM33jimznQu2mY7qKnDJdnu8LOnm39
A7tn8PdiLU6TzB16QdPtNPm0e+cwbKrN7yTy4MNwKv45ETBlxq9czTBFDziFD6Vp
E+b8qxt+Ev5ImizzicujKSu8V7aFxt4wKye/W+QLNaGeLuNsqRgG9Ea482GNbs9T
jEiL21tXbEPYWI0hfXGVu+sFTdgM5YXrILk7CFHkUyDQzVGhkEvzCq0zXL4ZmXEt
l/LcGLwbbiQYwQcqSGXo4xjJFVIj2yBLYDdbeTxRhNzmlP+iPGZTfHoCZ7s4pfvS
+CflCBHMgktmb6SEChFQOjiZo/qhfBTatEge2iBnbUO+bkOA8D2D0Wl3i3GFMRjw
+YdQg+234HUi6LN+p6h2wqBf+V4b0bmwF/376NJwQ57qyFH6Ul8C8yG07JpkA36K
n/VlQCqJAKAwPMV7N8DM9i4OppZSgh03wtnWLW5ZxFxzRuMt/z1s6vqC3TJByPE8
`protect END_PROTECTED
