`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6i5Vq79eyXRlGa7ftyjIl5HdQSlI/ql8o+fpycqGyCbbFCYUWvIQ4cBJSuVX93o3
7CJzogJM/uWozx4mIv4XXpLu02q8gWId/CkFtUZZyrKaYlLjut4OblgYDEbdSDHz
ZgmPNw0FxGmGX1uYl3EfvhLmnZcYaoOYQG2/wMPuWEKpJiGtbMxsJnL/pGir3Q67
BPILAyUPOXmZSLQfIOs7Pk5IP1woEHnCjEIBzneNUGLwMo8NdkWVyxOZoPrwU9J4
eV/pfhUfkWfbWX3OH+dcoSn7NZGQNIKALZ/lZ6RdUZFHgnQfqVVSkgZnisadoiFK
5rqprj7FmQ9P1XmuWIb6WmMGqTKMNlTelqFFyO7rqVXOSPAhDlWwcq/J9bLKgHH1
MypoyfxYcVRL25Ww4YfdzyMufISiTNZJcWPjNLNOYK/cS414N9ofn654plFnWLeV
gzZ/yETSI751YsLi5oMhtmm6BBMHldJuJHEF6PeGM+Y=
`protect END_PROTECTED
