`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9U+YtBJLkXnAzf7rupIxCBFV6da1KLhyk/zoK6bqSeP6LCguPdYzbILvHSp6KaCr
q/yqyxdYSVPJaYX9iF6eVH4Xp6Skxmy+Ax9rC31rryh059p+w/ukITR8fsWwRixg
1o4dghJV8Ftzd/dfdmRH8HC8AKH9YVgFW54HeYrPTXmrJtLB1jUHWoWvI+2LspMm
MuPZbCzA7CpJpIXf0IMiWMJoFQVMr0OAgK9VCXowgBXcMaSD4mQgqJmkCNNHSn7w
LcOVA79QUaQswdcwtsn3g2jtOcU7H396Jv14M40z/nB+gJ+GTI/Y/9RND8qkI2J4
LGFYvmHojQdIw9fHKnKKQZsxfXedYfQ0ps1kIq4ac2jLP3NaynwomjrDkKj9lyBk
isiQgZMSAqkDSdbZbP/0Lg==
`protect END_PROTECTED
