`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+XPwq8kXMMot4ER4XZQIQB6on3ftBou6Q5eXsHQ515vGw81BJtRxCH+1yFFLhi6z
NDFoW8ki0tYn8kt6tq1pOLFF7eW61TnXPZlMFpe4tFNsUbzh7Bd9mKkINMV+w6ph
JZSm4mLCKAk/oXRZrE5HMZcpOW+pJtmnb8of+qWdEFkgyvBnZSoev/98ylLXUOjW
DC1YsuErfHkuFJb28qeet4QRAGZ1q9fhuS40yV3CJ4lky1siurqkslyhbMK/crTM
3srXOYiet4kEK+HCfDsBMeZ11iykd3tHcIDgeJgF4F9AHNhu1hghNAHYTnIF2iwe
H8VcVyl1x3xgmX1ZPO73PzP9RIliVRmr3+UyRwEQbAMdL1gkOto1yL1fjm1cafqE
nUk7Bns+6IffLZovffdpJi/ZO43BsVjonurxa2uIhx301U2kPWdRAUgtMK74ZETd
oq/4VbWqFmMh+rgWrSBAsg2EsMd/tVUrFLprTIZPGqqe5BZXypEBaj4U53JDQDQl
cAVyITZFURJxoEVXgFnRBQyxvupirEkwd5c/shTgDtlKYqiD9N/ZCvSTQ1413lgo
2jAc2fsTGIOLZ8YdTqkvks5+zscTl15wpI1Tvzd3RLzZHfLDhBynPuUQxv5jgxPX
ljhZ3B5VLQEoi71ZKbq32UnvKllGPydX/wgnBga7e/TNKpxRrJDJL+3WNQJKcJve
`protect END_PROTECTED
