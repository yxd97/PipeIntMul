`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gnUFTn3DUQYD6dm4HxDXoU8oAPovAFfL6tgGMevikdF+3URl7w+6MMSN07RXXeew
bQJHxV1BKE6uEFZN1wz71WwS5MB02oB4WZdS7B3ypJKtzHGddaF0HqWneL5dmFO7
wVlMYFkufIBARbRRDNVgWvkbUW5AnWuiYsQsGwJ6E1PPuJidpAlRYId+diYEfDzf
hcwpMiuK8npuyse/lWVHZXE8kkXmd/Q0THcLlVCsGCSz5gjAjE9ch/dXv1HXxKQ0
ekxY6WSIGitaaMWS30P1V9mLpqS/FdN15DWRiqeP8Y0kqP1Od210HChmSPBDV/sF
ougdusIr5YBlIJyu3ahHrZ65x+OwMD2ZvaBXlfKAKDbTmu3SkF1qBILAfPHRWiCV
41/jRG1eebG9BcfyGqSmIry+odCil9ZcUByxvJOZAYsxGELSKuSGgmrXaPVgvBL6
`protect END_PROTECTED
