`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ScijYC/e1q9gejDGtPLMy28PHsodKC9sV1FXE8narVyWKLT/X6VQFAADpMwR3f/
mfSpY/eBABaTuBdJGoA/Fd+iibq74pz3pAjvHt3dJFhCCWMiRq/9GlHXriA1ovDF
jjX3Wl77vq1QojVdVjRs9zj5dtx3xSC+8TzqlF5ZJOomQoMy5u83XxE0Ii5O3vE4
qWMInrAV+WjUl1hkbSJTLaP59E2SAv5FaUeW87OEjkpEOXcHdCWB1cDQnN13plhU
/DEO0AtsauiRE7M2dc3OrE1lp04FSoEbu7YvXf6zi3ozjXa9yqYViPlIxQAmoLin
zamEhbTkJRef0oBN+MSh1fCwGVIETxr4/ju/0EVp2iMSk0duqUNWnQUT9Drlm3CL
pVdK9H9qmByZzjg2hCHCt6sc4jmLexUFkVw24bZewGtq5W3x39Owlv2P712S/t2W
kBIKX4+UCEb3BRVl0G8DVE7xzourk5qlIwydJa9jmOnGim6zHJ1XUsF61mawBv/a
h4HOv6aWqiuIGFRkVBICWXZOHZBiinAHTZltCKvO1OVPSXMRVdpldI6n88+rQ7kd
8Gt2MoSSsdQGteXGDGsBSHPsjK2z7Dq0BphzCR3e0fsrIJ1d2CVyLsLTXasmLEx3
0Vex54qI9bFAPtOypZBmrwKWdaHBA3n3nWDHJHacfee4kS5Y/hAYADkcwNsEi5Zi
BBpE/giDnvAnLmsN/Jnk9tZPF2WxxBFg19rzS/iU/9iwWDemS7xFd8elGVmR/pGv
+NoN+TxloiMfrLBfqjO/YA==
`protect END_PROTECTED
