`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
42zZv+WOYCEcBfqUyAoJ9DjTk71li97uTpDL0BYCx2v5PFGiIjfpOe3/oWwrYtak
vXDo7SxgR7j1QkoJLw5rCLls5DLTL5aYczqW6h3YJ/y6e715kI3WR0fQ6AEz1KoH
a7qzSq/dSzCZfGWPzExBlEntUio7jGyT6pMB0Pq6XV3S8akVRQ5RFoB6f+A12Oc8
T+PMVujEFC1pRR9tTulTaecf6d6wGL/ZbVa80y9hxUrU+KewNx80bGuTlu6LVf2x
hoV2Zb2I7jQSx+9I2HDWVtcnoWyKD62owixqcSS2o6Z6SapanposNRh7MVx2UVzy
jY4cj4rTvitdxSPrsppEVJEVNlpziM3rbeF+VkkxGlAiyF45L/Qot3USbu93Thpp
1vo2FHBntpwVPp4cM95C5LUxiDnHebTeaeJOGgjbBglxcLpI6lCZ2+K6lsNrr4+x
cc6494QDSdf96XuQM8dQgFGoPnyANWMWtP4RpdfSNmMruuy9e6hJ/Uss+NWRZgVO
8AuY/CFFhiZOkcBBm1pE81GVc/xLk6boxBT4aTLCL3//Gf1ERsTu/EFX8Hh7J0zA
drmN3eI+vKn+2iwVeYOCIc7dSSEm2pGoQrVg4pop9+wCakIR0YiW/Dj62Tng8PYb
38zsL4UHh1X+k4Eh1hmnqqw2GMXQfiNAqgGWhqlVtfO+OavagYiD6Hx+doLpAFTd
kMyxMnAdAGwlkThrkuqs+KOZm75Y5xIqpiJgz/eJYzJMor2GOCl/n0eRpZcn2+ke
M/HNc8++Gz2Y6aXx/l6mngxQFDjKqVq6fE/ccij10U+AV1v1E+q5kPSzL60QA8nb
ZVi5JbWND055xm7Z8xh9stSahhIruq7bochpHPvE1uhpq7PcyGMO10HtjY2rd5w7
iUbg3aVtUgGtOKffYpU9gDgFPVZIG6fn+Du9829d86Bj3MYOz1aJ8FicAZft1tYf
PCZGXlu6bbXLhR+1LrbFahOxTjrXIZeNK+7arbJZRANpLkPTpReghrtVkFsqy2+e
QpBPBV6qYk5+38Uqi73nhcCBzkNqafDWiG6mkHHhRgmxZbmjWA6niGN+d1w1R+Ss
XZue9m9lTMrI3KBAfxKWVkSe101MDXBnQlC/bPdwnV5NygrcZuCGwwemox7MEzqx
0+ocjo+gc5DGeiQkTQ26QO1v61YzCgcwpE+QcSIW/Y9pjmNj87ztt8IUmM3GPFVH
ZbS/9af/7dOpoVGtAgk843hZ488e+VrQBmKQmlHd4SI+8idfsXHfzcoszDSt3ZFz
SNQQTZSwndpxKcmRRWVXoYSWQlECBrO8svQ1ZUzBO7cupiANfKPghwIt2d8YjGBh
dpm5StE9O24CqQdZIlG14WkCyGh6P/BzRmUBW1C517Buk0YiAzh5djIlNPpa74ni
84LK++NWULZkDgawrzYy2Kn2V8b7rA66zJ+rKdMBVM3T1NHaP3HTB/xYSlpQnevu
aKETpRXp3k5hOdssd7PzNfS1sn1vYrJw3obPiFOTCL+9PuuIBplFHu54L47OuVII
29cV+Dxmegrjw+GFYSkGhsXbhQzqBk0pe1F26f3NJP/L4T8FdUp6JXXgBVAqAw89
FyXS5BFpTDU4PgIx3hdShSCK4LaBo6E9AK3/yRx4aR6zy6kfNietbs91NN0I/ke1
V1f2ij+T4TGz7Ot4QREgI0cIfZ1o1p+w2+q8P+iVlgoosNXSBwuOotGLoGuECVRA
qKv8ctqLrCILFLBpGnVuVlivL6eDV8aNGbqVvNbKN1ykMWxhcYnMFc9Jakemtnm/
V1ZQjAVlwI8IhKLljKgQH2LsDkXqrV8HxUExBS7u/AmU9e6zIiDmlCDSyEcYAXCT
QzCEfvGO1Y2108LFRzO9+yaxxy8JS0oU0sWQvQ/Qj1g0L7PG3P2W3Bm+vKoR++97
JwkRjCFZPCYoTS5Fwy3ht/r4mzZSyACNncKznZ5mr8j8W86Mvt9p2bm6twOtEdnG
qSh11HRhBGAeWKoCS31D+tYUNZ1KGrbsAgXepzPn+8xIEwyZFQ1cHDRf87X+Cwxi
Bbyk6d4fcMDk033Xaab3t5h59RLT5fpR1e3pD0f16P8ALxV/24J+mcJy5fiQU3Fz
6X1Na3xb3smwlk7lG2pfMNvUvvSdolc12F/F2A98JQlTML241oLnmSwbM8fApRBE
QwOMeZgkSuoFVSx4+BRu0g==
`protect END_PROTECTED
