`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Df0JYpVdQ+CjcXIxgSA8wsSWhdLFdOmyndzU3lYIFYvQAIxipia3fiiH0N5kXzPp
0CPpsaLtMOSRIwVFufMRobOlvG7mzTGtTAnkvbJeYjkFwGEHMGOaGrK9/Bes7Thk
1hNKiYoZCodNxDlrGt6EFu5poQJHstA3n/muAv+UTP5qEJdfyzCmkNKqwx25CXl6
GgTRs7GI4jdfvgxDXLYnZSa01eV/wGVTUYqUDQOuxpV4ohtrM1qmYpa3rentY+Ol
m2MntH3hF9NhIUVwJMuF8rNYpIhcazUBVdDauMIGc9mdzh9fm6EqMSGnKbb8M+cW
vBr43QPYrQYi00qSWUdOoruurWla695hdHRMi3vIrqh2TvE7GTFUU3QbZHeR/1kS
GwXGd/l7X6/pvzSVhX8XJt27hapZt6UEeJ9vACICrdySWt0xGkXOuR/C90rP2C3Z
7UQlhhAm9eUTcVsuLh0F1buj1eBC/8/U6OFWJSf6BVffyeTIOSelEs+5xVICeE/m
hwjCFJMSHU5ckb/KjkUsuwZGcjd2JdqNJanocZILUApPJ3Z/xkq0IUnqC/WwwFew
y9wGZn9eGZ9K7QmMA6znWUnlfMXL+NJy3xhraP4P8gUe+0MgLZdCZwqga64WCUZc
bKKVylUdVVGiS0KmGZMWBupxlepdnv/YlvBq1uVzMxV3KIb45emWTutd6nraHIxz
P47mscUNLWIL9tihcdrdIgEbNiGD/2ad/87OblEelLtuQv1C/ZqWuIYAC6BctoIh
Ut+2xo/0ayj3EWGFBh3TEg==
`protect END_PROTECTED
