`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PkEuvv8N7voNCpUy7TaGyVEH7R0M4WD0F8mtAjHeMN9xmNLmzQZ/iGOt8Gs3sriP
64cjAp/IAzs36L+nAHiUBwwud0+qweH4NLa1TYiRoY1TVMEgOuXsYf3QRWnjrQC/
lrl+jf16wtXVcBxmEB5lSn0WKAp3/t1gxlaPGOqZB3uMqIWv1jgCg7KxrC+Ui6m0
WmQrFdQBhQM1inMeT+Xq2lQ9EXCWOAgfdEommVGaTrmjRhV5LdmWN3QqBkD7lUVL
8P/I+dzGQKT0vfirZR6UbztS5Yg8BTLKw1EfYZVfMRcLmP8z5sOTGBGr6nUXDdkv
tbuz/MsPprpVR8F0ZTuZpLKkrajcnLMfkpnio5NXFJNv/Y6f4ojui8vwzacVCPwP
7JVDWlImy9zda49mczvz3q0vgweZmgaHzSp0ISbYxCZUGcgUViUf3mjiIntBEbbF
fQrg+OXNKhvSee6KFsaspCAYAEmzI0BCr5W5nR0GF5z80NAg8BiEi+c4KijO5aQZ
ObWcFY65ztQFn5eeCUiVQKIg2JAowoxNtaEPcVml1K/KN2hQ5p+0BiP0UKtLMvMj
A7t61EjMLYX/9BYVTw8LZGvsD3/4TLu+WR8Ewycn5WCG5YPVWii8ei9VHz3DduCN
7Wbg0FcTsrGHO349tM8U2PMEl4RCuwTa36o7qPnAnUnuEOi8HRsmC7Yp6ENbEeJC
`protect END_PROTECTED
