`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPEwlpGcj/e4KGUSGLxKM0oDbu/4u3E9G1jvwZdJUsYWIYNDn+6upP9gn8f1UV4K
k3VaAVV9Pju5zSii2WdHn30d7HJPXb1qwFxZQ6yJW6tirqJigjjpSeYx+BajG2fE
H61U2E1CzQJltDJLc4H5ye658WSvUBwfQsgjQTLITXV8VFg/dbwFZX1Y2sKvUpbx
vMC2ZDlWRCqdUveiVm+HEZUkTm5QmAQev28HxRCJ6qSCdA1TgfEQvnehgVt8uU1k
PiRnex2HhHprRNRmd0MSZRlW8u46RNSz149r1uWn98iZbDKoeHGvrjDeKunrrq6A
SBa0Q0epVFfO7xCLbWeB2LkhwEB0UH+okNYWUH7b0ix+8C2/OwTH57H2MT/EnMdN
ZFELvg1+VwOSJf1cqCczhohxGFvsdN+Hjgx/z9DIMshdMn5DS43w4eM26b1j+fRw
`protect END_PROTECTED
