`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VnLj3JsrEvKp3Dnkwn+bEN8zT8mXZbnGeM0TYQmGgV6LcfEOcOIzMPY1Mk+syoWo
sYX8V1awd5tD9kM4Cdvy+r3+KNixDtQMNtSp4nrMF4LOuInyR9KpbwAbDZ2+mx61
ZlMKawoUlsO3QAFQxIG2joZephxhVyl26o2deYNlwYHTkb3JQ6ON3WRPaqn8o468
+m4R7sG2jwgoIxqsZcOd5tBaBWLyM7rN/Z/cEl7aA7bou3z5LagfvjmqO2C18kCY
XXwi35HGRerIE14f/R0uSwpOjBzDPPdxQ6YnzuWumj49/EhN0tHWCYYgrkHdj1vQ
d44G3Tqv13UPbyV/6lHMVIY/rGkuQWvpfRImkdcDVVyY1/N1BU/yNS93Q1DzPxZB
5RK4omwOcwSd/KtK4DQVj4hkzPCKzgJ+MPAUrZSvWdo=
`protect END_PROTECTED
