`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8xQnndg0aC+fE022FSJw9qJJJIyBKp1rT/1HRx02QNI/PhAwxRY63Za0iVHgXf/
8iY2N21Q6F9ApYJj9/pysM4UQdC7Sp/F8aMYqiu8vfymD5c3c+6+vxPGmjkfjNuS
hM8D6wmQTxVJxGxcegn55eppgjhtHtU5QivYD1RZQ6QlKx6zQb7mEjbgFbGAA3oA
K7e5cLMx9y5QekSeDViWK+VX/c2RP6vTTU1//n4qVPeDRymQRJmdFfMi//jMZGu7
sWjJRML2krVfm4IjL8lnRqyE4kC2XJLykZbb16tFDPDi3Ds/G2yses9+ggp94FD2
WB4/cgMzJXRtZXr8Mf2UEkNuMF13nDQFpAOKjh1IvY5yG3Yca+6ZBQAWzR+M90O5
Tm0vV/M3mcgVBVN/ASbK0Rx+K+JPRLWAvFCVXIIatk2SK+GgiFErW3NMNxf+kBy7
ykZFWwQeX8F8YWhIU63n1wklliGNhKWjbA+Gfv4Myyrj15xhTEKc8RmFwZMLf6f9
Jb9CJIdHRWj3m5es/kWEfyiPURe1jWfDagCgPiyKTftpz/5OgDTIX8MS9wph9jOK
jZ/6F7ssnmymQWG3qORYIoThhrGOGxYHGoquFvNPZn7HowB/Dj0WJ9KsALhiDHLk
DcU5WB+f3y0OjRlRzXtLzo9OmDCXfK7b8ZTVi1No2rKxfGMWRZqtbyHmZowJRet0
HA8San6HQYoz2sA68kHAIVqJ7bNO62q5Ptv9VyrMwFyBuE82vCJVpqE+FyRuUacm
GB+IFmFwEvKmlCII/N2YdNbZAGUgGtvSgC6bZKDoW3puBEgZwY5W7mAfKATaANwm
2P/BKlcw7ynuku1cMjsYgZDSknyhAASrIqmnMULf6yMIWkm5eC74OxhtbI0WEzwg
X92zIaPuLbN/GG5h70zoUYK5/hK83F5hnVuSF4ZTCmUFcHOvtoNmV8bKVi2OIAvc
u0tE1hxUhodFPKIwBtM3crhh5lb9BEDXIJ2KLx5z4+u+LsE5FimztnHw/jmv9lUQ
0E6RUxi4gLHv7u2zABWxI1sAsSsZlobgwqKUAS9DlglL7UeyLpR0Rhn33olq5YqQ
hvoc7U+XIyGTkGSze6Y7YkIohFgXNzvEOyyDmP1litKtr8DdN2mvHBfhNy5NLKtz
p4okuO8Upr+D4mByBaMDXAd38xqQSH0wd3+4r60/CIoNCfdUKbUodDsVYRaXpKTO
ki0WJcXhAnG02jM7Nu269ECYGSye5vkPhnMFldiKJR6Za+4u8RV4RCqarFtJSYY1
xgrNclvl4nTC1oORtDjeB0oX9JFxIJg/BA/PLZneRsEePLlTHrjZSkKT34Um08h/
F8QTT8j+wb4wFomxP895YdcDSu3N5Mj1rBHvHsMH1PKm1+zRKFYE1gmlIE852IHk
A4+NznZoSVvz5TJ4d67eoQ8TzveZzacwW4b9bXJao8MsE0VqpropRQpwcWDmpcGA
Ck0hHvC6yzoPEL/0lM1UXM+7LLFB+rUmO8TupQrdBm/MphjDhKDvppGLW8bKKVA4
6vrzemnRprUNwF4GHCvNaLX2eHOinCRIbbmF4ZrebOkMogOrxqWOco4JO4VwVvAN
6diUiS0280qvcGfJTgX3uRVrVifvAHQXSXWqx2HgmBNc/X8GhIPdxtCyb6XI8jyn
0TohINTCu2aTt2rB5UWUEtpkmKnfW2/V/EkGqh0+Gn+z5MB/V1ILpzYpyHQHFmyH
Eaq2Nu1P4jqdC6MjR4sGmjMXxD0YqqoaZYwIpZkHDUwWr+G6YqPEZM1UxdaIWpJS
VRdtgESS63hE2f2Dom6F/2W7btWArVTnY8DwRUp8B+LnjlsBiBXf8IStsfbWlMdj
vSf7v6Bd5J7/y6+Pc+ZetIskp0eJgDMbG43N9Wz93r0d7XF7Uw3WhRHmWIuq2aqH
k+3IyMKYFSoCewchocN0kYOO8UN4Mrobt2K4DB7dKpfjsFF4A6xN/kAdEwIKL2Uc
8zoQWWjpc3p2bTILzLYhigpG6dOJ0BMlM7Z1J1Q9QbRHhhZzilkJy3L17FjTwX3T
RCnJflQ0XqXMFygbHPmGjTHDanjd6OOTV+JCUInulkKXgZd3MUGb4RlgSXy1xIMO
yhyIy7uxB9zop36KSCvRxjqSkCxQD8FQt1rKHWoN07lD4/hsnRGL7/ooZFHjKgr/
yfR6TUOOVSzqm7nY/y8PaHPnirZRcP6dHEy35yQGaj3qy/HEiY75nqKaIwX2csBm
tNZ2aX3WPoAHL63YjUoM7pxM33r+LI77yxXtL96zoS6FPL4QvG98YGIpmgtl8jRA
iTG8r3N8D3DTfCOR6r6C+9MzrKTxNzTNLy/YYZSC1wG7Dep1eVMnPCtM942rhwSu
CKQp6J1zlD/1m7ydR0ZGuAwQBavl+LA7dhw2E5Kdq/UQcomsjrT3fps2aTxDL66O
aHiM3RcKcEDPnsen6wD99Pe/GowWAioyv5GGUkb5QJ9/KCK3DIbXPQ9klApyvnNQ
EuymOYkwVMm2nFB1+GktT8IkMFlL6cFMbdJhUhgu+GLlrKR8447koWbBBU9zt4I8
UHbKy6+EQqc+4VfK/EKrkWG+sroQLH8YRwmpT6i10/tlYMg5v/ZplI5LTP9Ql7lh
4B6u0dZhRcOmCgI1WNB4YkNnCoriBve5AdF4MwWWyNYxfzvG71IcNP6XeueKmQXw
BEo3EEJz4kYiKXelflkDEpGW+4rgSjB9P4aJhJdtmycl68+kqveva6zCyD/0hTj7
rIm7YSWwvz5Yb9PGFNLtIHYCi/L4d4Yid0aVmgT7dPPn4xNjkfyR2pVbo1uaPLLi
UfRM3DtwL3VKzCmT0EcsDI/L9FWqIMWJW79mba6uPbi4GmQFh4k5RPtPVPnBc4Uf
IxHJgTsOQL8WEAo1daTfLn+61a1nPSwNxErmC0n8EnZmXbgxSJhIepF2vTpHnoAz
MCKtT27MqhfH+IywtVyJ1QDmcmzZxmarf07YzK/UsW2MMihTV15Iq4xsAmoc+Lo1
yktfDapQ+xVWZp3Ow3YEej16YUg5/w3bKePw0PKqVnhhqQUXv2NopoaeILSQqo32
dBby4zLykhm2ID34ToPLiLVwHsm6fnF3sEZXrD7W2cD8YdFwCrZJ0KAhae0MhDXr
7HDopYXA5kKQWV0ZVnz+AEyd+e1jb2HIXnXpEfsIW5bMltVZgtgX/CWxARP/B06j
H+oqTcv3dxoWARFUSV636Cp/Kg9hKQHeYEXfoEJiX7/DIGxk7l+Bl2cL9BQNjsLw
+3pbqrmPHrobwOCqiQK20Q==
`protect END_PROTECTED
