`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C5+IU6Q3eoPMJfAaVBiN2FQirVanhFdc97uBj7ViGRM5vTwY9XVrFgvicy2W3s3h
XoQmCOLATQr0BNjMXJsuH0J7szjsmp29hPkuImbbCGaCXNY6ios6kYxs5loPTO3S
6bbYMCpQCkiguZfhwczI3qkNK0Ljm7U02JQufTWa6lJrlIxomThxesPRhcUKdLiB
TFW4RxEVEgYOCb3otKDKY+FY0olOxKQywmMe/Y0oBFRWEPZHnNLl1aGg4y7lzwng
6CUOUwwV987VYbiAKUBI9TQGYAft3qWpRK/8udZj/BqhkFQbMJJ4jrE67NRD7k4Z
R4W6Wl/LBk1xbKcP/ZrErDTSFT8cXyM8stoELr4frXkDkLRZpG6Gg9QJvHACgCxM
VCp830CrMvbahdouRZ4nKeFRH5XgpTZAyoqD/gdU5yH1nqEDmj2WQkhCdFTOYe+m
M6bYCXVlOe9rO6UGiW3uUQUgCH2JVYY1YjoX+8vBR8BiFL5pqag7FjzyDSPT6EBz
9v6plskli9OwlZyEDPiBExHbz5XlMq1Adh0olkdamng+I2up4jwQ5Jo50lz6SwDj
jPNW8znytLtnYIdmc9Gve5UYLbUuSqhSPP5FxGRHc0eIPEa7bMVzr6jfRKnQJvqV
kld7gYzI+FbtJmrkqJl9yCRlSsIRyAE023z26UlP4EKlQVSH6+aAPDQBcs8j2sr2
1KVBq9Vn7erIPNxrIl6BMjYH8fd94abFBi7/PadaN0W1Jt+llzqbN0Vhre0ivaRq
KxoO/lJgzgKA3U41n5rTpWk6mjP3EBO93tZfXDGxs5pROVJaWLizwAoMK4PVdGiL
TtmJUGXv9IDPQL9tWgMoGzFZCdr6samx8Bt+EuvHdczvmMWKGjdo+qmD0OWBCdGH
z640QrxAVs/gigVQ9sTqJo/6ZGMampwASYVHJf11CJf/ZCxRIIs1TKcxnhcFwCMb
zjbwkwPiEnf2Ly+V5NX8yLKRVMyN8Rm4F6dqHeTxu/F5IZqF49eAWsAKj4kVuooC
C+CR82LmJjYTNNGMzkl41Zvp2hm2ld8ZaHaWChYsGXETTtHAAHwWnFKrmowGQErK
DzBGBlLkKJTCeJ/pdybghHQxSa6xwvu1K6/4nKyP2U9tfGBL46hKyHZ2Q1kLE+ne
kc/BQMj8pGYSx8mWeZrQEQwgAiSklXdVr3u/ZYri60iyZgzIyIkyVopuManRZSN1
wTkZODxVqatm2TIqmr/j3TCnO3JROw65edcyt76k6sRrMJBWQaXthCHiN4E4+gao
j91UVPJtwU448QY90Mu0O7dh3qhHhAgX8VnhnFFF96pkqddACPPCmdAsoRBSh42U
qpiYiv0C3qJXn5ushM0ZImLpi0vKk+KrBJQYBCOUYJ8Iq0Y8BfY67RcmLA0QrXHF
X7q1/5LY8MpONf5PffcKwZuki/jspour1NZNb+LvVmiLNISjkLLWkRDGsaGQeTZ3
KwWNlwu2EIudHOIa18j4fqHfQxUjU6Hw/3ooqD9vRoU2PVg0eVhEJvYx5InceIlM
SHI6QFYAuk2s878egSr3Lsy6dihBTFi286NDMNW5csEyFsyKY6Ecfhtt8wj/sFYL
iWpmURFzRsAGois7WtPsrgMUkBzdlFKtPDPhAO1iMFMiVFv5zqaeRyWinm3HcMf/
cR9lwI6FYGC7A06MJCooXG7NPSF2HMZtfIyuOhL3bkEJUYIztwy9uXh/ilpkkcPY
SRmFmXocG3RUb22c/Qfrj+UM+Y6TpSqpjwXmZq6aBlvhuqUaiC8Vn4m103bGq/3r
jJMhl3QIPE7kP8GTl92cNE16li4UGPwUqia43fAfoNSr3kWuUF9vD3i/jYK7kHhZ
g/J30YshwML9sB6YlghDdN5dlsPiQWC3oxkqxWPo4pA=
`protect END_PROTECTED
