`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cOr5rKA2Q6uVtoOc7t1ND6piYL6keTLNyqMXBlt57M+cx98Yqg93hUDPjakPGHlX
M+PFVbh6i+8XKVP79AuuefeM3284Kv2VSCNq+1SglG4ywuLzC3CS8sSOoOxGov0z
scOtryMqHiOh9/WB3hB8tzcL5B8MLrTFDOVby2McylNdYZcrjaeD2jebH4NpZUPm
xV7oufemTNf999oFhNBDI0tVzalp9quMDqGNhFO5uM+LDwa7ArsE7NATvec9D9qq
41heFWASiwWEMgE+e8xiDX4LvgfD1X91EknhI+KgM4R0ky6ma6Kb1jpmNZaKJZcH
5pO8wBE4LB+QbcUtByn/Prxw6tOiySJZ4Bsdqv6scZOv+zgx8zDoOw4Z96gdluEQ
1oQwoQehPci2OJF1Y6CSWQ==
`protect END_PROTECTED
