`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
upD33Axuii5PP/RDdV6lwZjW/lb3kQ94g7mCe0ju71UToDWJm9zp0RYxD/JORjKQ
htUuJjBpnX+c9G37dTmYnwZ7SYl5YKXnwlPjzmQEvL5Zy6z7y/9eSx1tCfd75ir/
I7K3YeUWRECX4uTJmknw7yodAHfMVOsk2XIlzr1JXYPmVqDYxQTSdsAf4deSd932
jLYPxdPYViPwD7iwXoMUTeL/ebYieT4xRzC6+E7xuVEirXX+jPQOUfaHg1dNpKw8
t5zDQh892S3NP33Z73XxIzg3H0zs+i6xJCjmfbZ5z3Stoa+c0gQ2e5zwT6rX1V3B
n09R6JKod3OWkE0g34D46cekmX4m2vGqxO0XcSDcGi6+1Z2qW5zmWGPqDvA7NZKy
pV28rGh+XMscW83fKVwnsq8dy9khNGT/ehmlF5gbd7aZO/+ke4B/fWi3DyHY4GN7
CLgNwZYB8N/nH0pfXQ8eemqZy6C+vAoOfEviOBg+mnHhrdiVmJFnRG/8H2tbw6kC
orGSqEBVw/kdUr7Tu1VBIP5lhR98r7SWOX2jcBC0gzOnZXapZmANH4rxGgw34yQr
rabUbU2C8/IjSl8EyMlpojcJaVOrOTV+77lt2HyCD+rylWjOfUU+A0F6irf1s+oJ
wWZtG78hBXvJVQXgTXkYpM3WrHL6C6n/hQ6OUJIK8rJk3j+WC5dnh5TkpKjiw2RE
H83vFznKufGlvYJ7RxR2n37ux63iGiEHkgbvZNYIApu52hao/b7tARNyUnilII87
UEKY7E5YZIaDVGjH6jyWDrCc/0zWDoGcHJ+Qo25H2oKzs7W1GqW9lJHk7SsNBmNs
ekj+UVEWbDFGsuSxeCTHx5EX3pVusklV7uOk8qtq5G1pCrH+FAlZHm2DCd1JW8u5
SQKpuqZtYPn/tvRwt37RNPFAg0AJAanwrt3EULsSVRw=
`protect END_PROTECTED
