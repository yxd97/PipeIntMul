`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KXMSyN6UDO8al/tEmfcYX2PKU2V23nW7r6qWr2qDCALrZ3bFffWzwg5lonChkj8N
G/Ivn0Tck+rnF1PQRxKHh7f8dXtc8T/IPRQi7enhsdt4eDkJc/HHvbFr5bs3c7FN
MRt9FXPrAs9Be321M9qWroKWYuBMRdts9fnAFb82KS0GHQYV6+mJCmdK5ApWzkfF
bOPG6v8xDJ1uQ3/LKgNLJDfbuCl5OJlSpbBEq73jMdsfssoXnkQDdRqUOzZI00TF
3IEdvpYNx0fL+0lSqqtj12y93Ib9KFunWp5Nn14R/eeG58gTTRKmEBg19g+xYGel
X/z4INuFuc1c0RCZxnfyqB8qhdv6DudCcZo1Zy/4INggrYnNJlTxVCufM0l+envi
34I3MLXQU8g0O4Z9mXSD25OudN2hL8cgqxJIrGfDFdfWQ4hLS10ZGJzMdRXoqKYW
`protect END_PROTECTED
