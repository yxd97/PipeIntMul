`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EWYH0g/cjhsm5ai0Kp0V51a6hXTw7JgpVehHHAvFeVsXQV1EMlLQEu1IaDTGvJ44
hFGtqSQvJ1DrpvyMSLGdtCLIDaK2qul09/yR73SRZI7AKuQR3Wod77YQVLSOnV7Z
kJQGsU8tKdymRj1VKTPDoN3onoy/5eQ4X9hbhk7sTTvZ96nTKI13G7PG6E7mYZK7
bvoMVsX61T5W+AuDpScL2GC+najZ71RROwaeTULN4LJI0Ja0rsG02QK0dGpzR+zA
2lz6pOiFNpNddNykmwDNOzu7/IpYHb7sbFt/neNy4Edd/yx/W9JwQu/rNpYrI/aF
FyaGd0gMZTmV4VwlcfOOVohdh8osZrGE0WUojCPixwlrCaiJJq3GqCLmwz12hoGL
8exyFOOj3DkSAFQhocseheewd9o3ZEbFHrs2Bwujw4Hpi4U/8nsiHToOQSHSq4b4
ncHUeD5uvMivPifmGY82Hve/od6f0/IyWnSqZmFG5dkb1zTCEMD/x9a7A+XA0QLk
8a5kyThpOChFtnbb4twrVGsj8ubpspnLlb0rMl7873PekpQnSvTMehi5+N4exCm4
L4xK8Q8d2VMqpmSo5+u0uu+omSLpS94WGIcwIzxWrjc17brnUBKCgLym6G4In3S8
9YiLBjAz+CXDm3QqCTgvoWs+LpvTgM28qreNilWN/vy/hIopxjFFbd0CGra/sPHP
pPuf9RoJpczCQSSeuislozvlgqn9UZfK67ipJSk+dUeVkc75C0y6RRjE9BmTEfWw
q3eX5/T057B5dTw+LlRUZg==
`protect END_PROTECTED
