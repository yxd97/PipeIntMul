`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RV72dXvqPaO23VJvZ0Tx9bqa8HidSmKTvL56170N4ZtWFcMOfyZMPKOfyvoh3q/E
ut92nb0pUG09k+OTXsudygIL2//FWdfeNvHMTeMSNcMhICJvVxmed/EDhHphJoWt
KJM69GZQEyRCi3DCQE+QKGlaGaD5kaBr5qts+Bj8Rpfu9potPgrgdwk+QYM7v4Ko
azrWdcqfyAUmpnhuVctTpNjtPKJ4FieZqGwlsb5GIZq+OAvu2g1qba2iMiQDfdhr
YDukj1x7U2owoiEN5Eo0g0IWXuuCyu45Y3Np5vVuayLeBVoeKoBQBNcbOEoyhWmY
xU2vJvw3rV98U7kNFwESoKYR0v4SR8H4dn2gFiKW30pXEXBR+DP+iS4Xvfy+TSBm
yPfd2iqvjTYCLfo/oLOGIg==
`protect END_PROTECTED
