`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bVmzomLifuAZkj0UJvmd5HLAdfY05bg6HQ3GK/QLR8/AqZxxC23xn0D888NuwnkO
v6ra6EiOj3GZMl91824E5TYRkPLqZH5feesu8kTJRdGyr15kjLiSi8muk4Z0H/wm
XOzdeHjIaVfp0XQ9EJAfHF2ynxvjGrJGFUe0x/CjbB6YuBWTJVOASR3QV5NAUMsy
Kx0HaNSviFbFRtR0LOfMWuBZCLPxZ4iH1l1OUo8r/3+OrQQhMViMbpzzPYQUvAYv
WhFcvpigzkYw3A8KYJSNVzlzrCH/c3Y2V1m+tq0zzv3On+YqYR30V5g1udUi0+zK
yrwE0/yIrkde30FqPUv4J1xp98FtJCI7Bmr7GZNrXFMnivLp9RtGHKX3UErb2z7K
TRMhfnzHsK+u61ZhXMVC9RM0wGpvOxVCMctpLlF4x8CRFWgsipMspgDgIlWuTrtV
X2Yj83GlIZ4i+izBSpURr4JHAOHmbbdd7Nv0457m9u46js2P5xoOTSGuNd5nSxJ2
5Sznd/F4712m1MGjIY3CaTsB1D8zZUOBdw54jeN1ZLNTqBRHX4kiHQL0kCFzDLOu
0ZsBAndi3GeTmlb/lNalSjQZ4u70JxNZqjPKUZkIkRtBKk0KuGORs/jTKgGrFQmc
pi83VLRb2qL8+VzlwdmbFQ/DS5MiK1mYzP51bVvDdYLBPg1g34HAtOaAG2FVMsne
ZZH/gjAGP0n+H2iAPveGAGEmwoxZbWh2Ja7RMDTjn7gBzy/C84ynFvBiBjxh6c2s
KNyrYxWl3ImOEpVXAN4nCTH0wJYp/QrQ1kA2Z7LpwVoVTC21jLEWt5THA1wmXYtp
oeCU1yNRkcJRAZJEhtFDye4BvLJW3WVywOivl0Y9OrhgjBLkO5lchiCdgZxqa9NM
atch4PD/jzu9kZTefp4C6HYczQ7hQkUjcKP4aN82Q8S4jVyJaUHWi+U75AODZuaB
OmRut5mfYG2vGcKjM66qjIrNq+2jj3bDcO89C56qG3i34iotoDpmWjN439vKAuij
GMXkzxYX3d4M0godkYAONQJtWDgJR68Aob3kIbQ5lo8W//IK2Verxnku/SdsHNJ9
XjIJJF2ySyWIhMEDof1qzc+dGFFN+39xFdhEmT7yEx293aisD105qI0x99/Ap4/j
3F2GryKsVoJqJ9r5/7ucc0HBqH14NjejbIOxgfToH1O0l7JbUqnmZJhFAELA5uDv
anxmb+tQM0U0WrwpuArHgRZECroeK2ijLFv5rxbjCkrAWlSFrt2in5Aadbhos3o2
EgxhM3/p/YoRFAx5MeQlSLa8nQeIaoi6B0UR7z0WbUGhCTuf4SfYNePLa+eCdhei
ClXlvXwLlEH05uyM3d+/CKWRW/KcJbDg0ZcAwgCK7LBOdJPzjdHIi/0OgoLJKO7s
wKZla+EhEBNtD+ONRO+4vMz+hULR59QmcF0EKlrW7ma+Rh3ZAFG924EBm3v0jrIa
z/8Tsgmc7JrjNvm0MNh6g/sOB8M1ZOIW2TK6N6WdJmA2Nth+p+1c7mRF79epSngy
kmnjNAt6PqnVIcEDaUALuQdoI7WxhsSa6ttmRlP8ooRAQweTRrgl43Jqbqi6J4Gz
fHOyjb2Gg/p0GbGs5cDx0U/PeOUyYgeG/KQVbRAmglPYywb3ww3CXF8cvzOsVfv0
99if4Nvbr7tcXBxQKP3AwSyVe+ODpN48WK2aQjAGD1EPy1IevmMFWU8Mi+D/c8kl
FxPiQfR3YL5rtg5zX7UvFigbLEQxRWAzLVaU7ddTHuCJrmQHeJUmNlrEMxvY0MEf
tgMR0dasJiRy57lR4gjlY5flccLL2Ub4tChPBPHdZ1a+ygiLAaljG5eHGYGFzJY9
NYrZMK99Leee6VP4SPrBj/HacN2ko7CXhj2r/pB4KgBZpK/xOPUf262pte4UaSvS
0kE8ptkJbwNTbD6h1DtLQn44VGP+CDSn5cxQDXzgFw0J/JwiIfsjTaaoFeogT6Tq
MwS3RsNBWC//nVd+bGL64TNylmQYbAA/RVBWMpJibbQtzj0JEkzNbTwL/SAC+urZ
0I9q+s6R5ihjfQz+k1GTtmBUp0N+h0oa1e/mkbUS9grwjY6E2OzrkSK1JbSAwrh6
dHyrZk6+uIJnew1kNnc+S0TvkpJ9GR7CbYW9jVk1XufoI2lKgfWpV7MecmFS0yts
/OAIJFZ11/49YnrrMAQ6NV3oMY/gqL+Lahlw24zq5/0s0jYLPmJa79YP3uF3FeAT
QKW7M+nrKkxNjkbHjFVyxjyzPHuby/38Ikwd3Ax8+2GEI5hUI9LzDpLiPeiZpWnB
qqQAjVsTm3KoV2pqNecXRNlbuZpW/ek7oYjyABklwWmuyxBYmf/TJ8EuLTwXLrgQ
uxbzEpoS+6n17FqwWcS0OoNMzFsP8T+r6XL1jRMkIhO9k3O+XeYYr33qqMLELb2J
AsVC7ykwkz8ZhESZe/Z9nupEieIqgfWJR75s6+idIQTgxh8b3Os0A+9gdU4OUA3e
d8pFnqR9Yc5g8DQ5+eRPX550d0F3RBRYVVJIqWJhRGIvdEkBOK7f8uk8d6mSeslb
l0EptQgsHHwRKHpYGtB7x3fCjYh1AnIZN95zsbTmsavXeorC0KLG1Xq7S+wuLqjE
A0cn2IzWx7ZIu1EccLs0aXTO8c6icoTxDHo0kvWPesMYCvOaH1SpFDf4MpXDJA4q
TiRm2XTDjQ5dvT+AadW2xoqp8dO38lplRUlKBQ2QxYiLe18hLl49ZWA5nW7K502H
n8ZU0LiCySqRV/o91rU/iNovDvHxy9bp6O8VHvKaDjRdWPBW+S4pQmtPe2iKmRWm
+euZ/+hfklhGn2MzjQTSpjbkCwzwCAGeMviLvRHbSIlK2DH7W4IExPoBvrA6BMYp
AziM9Z0WrNXvQkFiqGlkgv48t5/0jJQ/J22CDka2HG6Go89dT57mhNVKK3i5Vu4E
dHo3ipbZx10eM3p8yx52xL+w8gkcSWtgelrHBmgobpmI2frMOvLxqy5P0NgBVsxK
BUT16K8UVvgubt11NS5OatT1L+aTdO6NiWu4TbM977rrZwSs4mFxwQCmwsLtBrUt
yvVlCgbrShMW9CC2idR14o/dbTdDQ2eZE4UifqeS43tcDLERmwuvmx1CzWcIpwEv
W8IJ5zg5B0deLp9CuEMJJOmAPEsz4G9jEtUEoRzkCU3AknWl7IMQmIKo+C5wJ5bh
QwtIeeO6O0rxWbtyxo43rIbmFnpui958WBsfxpt0+NTd/EUwgIBwPy+IX7apnKQ2
UvWnsZA8FGfzgOVtVaAYbQqmsNKDfmxzBKPG/D3eCKI7l9roWatlKYRKqGektCi7
HWr14rI3usk5o0AGrrThcrp2Tpe6B/28DPm+lZir7TtxZk7XeplMCwtwM5Antw+p
5axSEFLbr43Dq63g8E55nJv/pyrAAqG0B6DxCUSdc/g7oCrbIzd3G2mPOILwxIMi
b1uxwETh02T4FfzmaZ1REd+VgwJgH335vAYo7ZSNhnCMi1WTp3dKDudUw2gb+Ob2
cDQ+qIC+VMyHeTybfGSKnHRwSbqFgWbuWKIFaXdKgRPPtADVuvjCvZgjPPAzfB77
F4MS87Vn1AegJYRS1IB/LneayYIMvId3TUKq/5UuvG/iLMZdnb6bO92rF+8sDG8L
XKm+wti8R4ll+4jsc+Q9KSgREfNn2IVsHoMGf5zXZm3ge325q+FByRVdtfY1dhzO
x+3tCKCpBPGzCX6nJm9eWmgtRNNYCtSYLabUd/DFNhP8dPeBKYrsadMOCXnD3ElS
ytlNHceCaLoShnNJsWyePqff3XtHkFvwe66ox2HZBlxJ0u/zrhtCa0/Dh0TDoYa8
aebGyYrQ98gNk4KRQpATz93xjXB8e6PP15TNM0tMfPuzfvPyrPrQqHR36Yp2TQJ5
yT/dAk5zB7Gaj0v1fNIdhCq7yPsgrIR4hcyrzbGhGqL9dvVtISvH3EOzqXzwxiWx
DD7OLBDUgOjP6b2vHiFJd37mAX6IBlrWkBejvyjTMTbiEzh2L9XxRAxSBN6abvw4
8pQMT3vSCEHnlcBSAjFQzzj+foqaVf3krfgQ8it32xYB5Z2G9sqt4/yBsW6+pG0B
BHg86WYUI9sAn0Yk6WrNOmQvwbqP+lksnr1hmvHlV2N2rLa/VlhF4OLT1Y5haLxV
ol4ZTcrD9IXWqlW5blKR0EPKUGt+QXKceuscA2Ob84MuDOtk16EBq0tAHFvzim07
IK4CjzSPZxoWNOOKbmZknCug4TDCC71sp0MqdkvdTv80GpKW5PYfC4kW5IK+BZ9W
JxZm8EEqRxeGNgGsrJxrOuJ3q6om4Eq4esh4fys3Yfk4vgRQ9wk7gLmzJK40flN7
IhyrQXNiaFhrr7PiHmyBJs0b/KtSFjuBCal1+1oQj9XIj0euVtzFXTTKdECgpk/1
ddfFk+1/DiJoYDAiL+qy17UdqhlPOFFHOhtKzJ+TmDRg7+jS1Yj5QDcDsoUvrXqZ
aX+1OHJrzQNpIZDEpg2uKrxvlGZG58D2e1BMD1whE8WFbe4MbqWEFI9y5SAPWUCf
xfQzTaErbWEtaBtjVtbX7lft2yT/f0b7UB9RM86S8EIT2sK5IjUoUzEy4xLIaqGb
kOslSaQOB1tuznCUEG/CPXrHX9Que7UVn2+WBJiy+NvQPRIb/wgU5nssq8KOG1gO
A4A4tHHZg6OP6aOmxt22TnM1LF4JwAHDlr2qw4QUzqJh1bHKLXKqCqqApBsIRFtT
JOpy33jEsujfxFgmAcfeSD8UjRjA6532f09gkXfS2vp6uoirb3KsWot/sEzRvl/0
scAgRJEe+ArQnArSwOjlU+2jCwU3j8qQGBU9Z/eoVc4jMY5jhU3lqIdOHBuuP/9C
9b+N2gCB/JFXKdF/Zn7m+fv0QFE4zFHe7MAlMom+TPQGUFJV/oy7IiXL8x39B6uq
+3DHB7hD4KhdkNbluOEXwIR0ohJxTgcohg3kFJWcewZIOBZPCvtpCEOsO/oSGp+l
EOAhX/ipbtQWg1reAPZKdC6kwSaE5e0gdoSJLvDhTd6YN++o+jxLUk97TEcubiU+
BgYClBY4znr9kyl3DEFwZcOEQTWdGmH1xhgXlLfhrspO8BvBw2kjDIW8oTNrP2c6
pzBkkHZODZ9evrMiakK+jvO85ulAFgngtG07TT+nQxQ9u2lBemv4hsLxxpVhAuUE
Y52sT9ROPvnS9vG5Hq/cVEjMsLLzSmJDtMgkxLR26NMPH7yPNgeJeIivFJJAchYK
l8MCJW9MigXI33Pbkqrh55yadyOhEEGwMiK9+n8IvC4NL7pxNNPYrklm8uBKvUwt
Kx4LH+DAjMBpZMMbvOMC8WquegocFVKSZ6mz+JovehbogFCC9cgCjeRvkvzEybjw
c9TXNjcCodX+EIjJUAX1bn4O4GTV6nY+/K0hSbeCfEn0RwkmJ60oKFjzkxVLZ4G8
PsUNK9gbGo3LMOazbfDwoHMmxIst5546KG3TqXwO0a4o6wg0KJENupLueL4wJ5Ir
yF9gZtN3He5J8fplPHJjk+kPg1gIAymO8+6VQRT6ggtkVcHvmrJvqiNmG7hrC8P1
XyLA5PcHpV73tB2O9R9+n9DvAEUK/dXK1vb3WjAkL7uSorBsdQs8LxrXGz0ASWKk
JAnrsXWl9f86zrcIKrv+RfSCtBoPhpK/sBvbDn8Bi9k+pk56NUvqIbbaa2y8AkCy
sWwFDtEwiVvmPsk/Tmwgt25jgxfJa/SakhvsrPS2dx6Vcbh2q47QhL1xr8wlPMMz
ZGLI3fTjp6PZfMDPaOK26to4FGN7jTXK/5jifT3jsZbNnR8o18JcZsHHZ8B6FeQ3
QsVJH0kYC+JoQe4tmo/8MmSBfjuJDyUyLNjcOHjv18WAT4HrHVoikJ7h1onTXZGd
/5tPJmHo1pvP2yE3bBdnX3hioTDYAg5EyTceJw0gCmMxtysDpQGhyWB8fFeWyjIG
UCWXVfS2oobdCpoP9bhk5yZg+k/ZshTaoQou1RGw1waKT4SnJjYImAxuYNf6/OYE
X/9JiLG/T6EVA3wi0GcmST830W0tR2AHhK7wvpizG+OfgmRlSTIpm2XH25Wu5QsN
yAsddL6NPToXVB3YrJyNe88vogBBEVX/4lccs0TVq5nt5X0w14JoRVh7iLhC7dDM
+NWYasWMtKZ25kOrX6mHeODIpe9PGKv81AZ9zFtxQRIsqaJTytBzurP0mCIHSaIl
CsaS9Rv0E+dDgqpTwF1P9AxZ6YFYlycYL+1sEodAVA+duz+7bFBFS3GIZjEOaCIt
i2DVuC0BuIHgq6nEjp1nW5cPDkViQ6jP+zuh/iudPW4PDSvj3ph/dfMYWypdBVCK
FDHM5s42iiPYGVAnL3OB49FyrOZEsq0Cewgqj3TdoRKpLHDefnYhdd5ylzt2v6KH
I6ibh5t3Ygm/IKGTFETiL6NRrkXzZQ+xKB3wMKUUklzS0V7DHF9eXAdx8zRO1yqT
naOXoDfzBquoAQ3vtrz+bABu4XhfKWCZTDFeBBpKV/EPrbwUaCqP9ux0lig5kLgk
RRvex0tvRxdsfmIBxBUEVSGm7rOKZkSsFzmrCPjz0jSRdQ0bvJ2TPCXeeDbftM1v
wHbHAciGR7rl0jc/oR6klILaA487DcNuRjW/+7IEEcSHbOK0QLDt6XxEd1gmtbAF
ciK5vxM4TYuFqnZ3ZJPFJmHut+fBp6gGcgeJlbyddY3HUC5/1mOKvE8tos0zzu4r
QitnF3+b/30+Zb3yfW/Xi62DnJHBC/ndLIzgo5lXhK2xZU7u4Dy9CLW7uWod/ZaQ
Fv4OnsgkA5pGhctDGKhDSCB4282JOIe3JqiL/RNqgYPyMnkE4kYUqD2mVGbDCbBU
sV1sPmWTjy2ZUEYGXyhLDFL4NiS5pTar9sJt+VKbcZtA5ZGOD5bjLv0KCfLIB4QV
Ii11iHtLj1UxgW/pudysgd+MyzEOWtJtydNWovmjYdeoljXrtsmA7Y1nUT/CXa9H
ucl9COzbd+uw19Hsu4ubdtVi0LZAFV38XaQc7x3ufmScBhlrCbJZyw9F5x6RhM8D
/oWEYpIsb5m7pYxLO+l0+uz3UxRuXg5lf4KrQA1+w5ck4EXO/oNruoWZG8C7Emcb
p/RBG1iAKJYvqlRc5I3h94lXIBdwETJ2nCKesBAkdNUKt5pVZZ5Eh3Bn0JhxPrY4
eR9htK+DXi9aSpV5XVVVK9uFNPobsF25cUvgJpRRcIqEAMAwisl63N1192MdnqQ5
7OgMjJR8RCuRMfhhjWfRJpGi+NkUuMN548xXFkfK1zyG7CjtzuhzpFNy7gCZn4y3
gZx2eKVEdQrhOaTxkuUIqTYdVkF536pI+0Z5XXo+tqXmHsh3Os37+zRXjpObLUHe
/TGAPJqLjGmPpFk27aWysjOGChzsWyS8ti0y6BLPjTOWDkAl3kKTAL9+mmgsWXw0
8brmSos5/v2hG75ydjwr0FmrE5yxG9IBOeMTy+nfba9NSgytVJFJlnhVSibbX/lC
7d6e+cWGmb34pMm1c3zUOIDi078R3qN3EOXFMBvXTHq8XIrwRd6JA7r5k/QT+We6
8Nn2ovFTdOQrYWr2ux/kAAXYAoxESAk3EFtWi1YA5Kcu2FeyJLfStHsXfQdJBTWQ
WtdjxPQG7wsLTruSvfH+lzU4r3ufSf2ZabHyOJswU2DRVkZMKrF2Inf34f9Su0oe
xNhp9ahnnkhat2kmmEP10/fDBBLJsdTigkO1uYjt2qddgWxkqnB+ul8ImnFxQI9C
fi8zWpD/Y6MnpqqueScF+hFUqe/AqaMcxbumTmezpHXOW4p55FulHWsJTSZoiLpo
wcxMkr+HMVtXA0EoeXGALJzE+c9GWOHR1j4xmwpMQw08GYl7Wqfha7EyoFy8t6cV
qZOlUg9x63FswCrbIJF3F7biZWismZ+PHf2HeUGCPcXP/XwqPULHKptZ7K16Jy4c
jCLlC5QQhso21KQu++f20rAhLcEKhcPMohPP10bvELVtM5ijcwZYMsrZvjLdV3Dv
4wGg74+TIdFZ++x1yqo+qoanoXOKDBJTev8lboNNpWMcDeFAzyPw0h0tDRQu/y9L
Adx5IpI3J9KT+bCHUeasdCazWBTbI5fdgsirgzAIWeWzHZxatgtl/MMANwVoAbAb
oP7sFHIvFkMoT7S0/oyHFf72GwBnoF0DlzfO0FhCdp+fQBIEGi3phSLJSjNvlD1X
Uv/pzIKYNQKv09U74x4HAqEqrqLg60VMSQdLpcwshM+49kzj2fHRZ4yrBI7Axvg8
MXwBeRz8mn1HYYrIJQoyS0Z09EmMqmnMC5qoDOCDREbYBgTm7oBqx2dwBrGcEq0K
bGd5KZmnaaW3YSI0++ke8sv9dWxc89At9jDkL8QRCwHrLZNXc3M5hB6SyME6y7G6
mWXS3odCD5lNfMBI6pOU9qw1S5GtDbGUnF+T4d0ZoJFutOjTmJv520I8ikT3z1mh
yEr7AWrGvALz92GGsIAANCMRcwhT6hoIiKbi/Ka2bOU=
`protect END_PROTECTED
