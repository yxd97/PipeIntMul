`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dz6H8nZ3xRhgVueWaNzRLuZSYw826fmtT4VhOh5OPgA2o1qah1qUWM9kWSLeQTR5
xd9b/KphetOezjNFbqSwiSy5BECOeTSKdJeiYNVzbsK4AMuL4cEeZa4d07mGk+Ld
pzrQjSj+42QCeUB7BnwgJrEIbFaUkAILEWbCSxpcnBWx45weEJXD0CgkbiJutoLU
jgM3MsoIkl0AMwslPLNLOnMpJ4V/Uh5kPTC9qRJI6PFKo6F3WhSZ1m+9AvvxjGXj
HSChVScPVeHASwCJBXgpODaZsSlU/GUt0sgakcHdb5Apb3CoWbcu2agAPMSnaHpK
qPJsy05R4WgtxBN8/7Cg7CF41taZdMyFUILffOSdVm/W9bCV1JZXr55WwYWa0hRb
N/LzkxscZd7OBy85Zw8XTgW0c9LaOtzzIgst/XVHQSR+zzrwiqanFUJR5WFANciN
/BHzp8cxgQSmWtRKuaDfjPodcUNK2evqBQz+1hBib8vFYJth0CO0bvinpoAcoO1Y
`protect END_PROTECTED
