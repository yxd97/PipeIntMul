`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jMRTAHiiEIPVPlURwi7UXPQMQ1u2AgQ4i3Rh+bxN8RpglhV2voh31J3wll+Xfq+4
wvMSVOxbMO/UOJt5aQ0JCu7pfzrnMoilXp3XsKZ+dN60dHhDjzlKOD3AfgTYIlLM
SNeohZNxfgahz2SEHpVspfhSM1EtuBTUujZlDB6mBBuLO68ghuZ4Bb5e0G8OgC1T
uuZnZMO1R3SxG9QzP8DmtNEUv88zxUIuBtkOwArvyjJAZt/VF//YPDfvm6uNZTDB
kchEM31mySL2KMe7WMZvmg==
`protect END_PROTECTED
