`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EI3T5FAWLyBz+thnsu2EP14U6tQgOryEzcRQfj+nOTWJkzqFfDxMBcp859HOOOry
eqsG9o9mmV9UaxAXpQ/+nbW9SdWj0gVSFDPdv89jm37/Ce1jGbwa+lGsaMC1IajA
kz71qrm80038PWaRgAb61UbKrYCAO04f4dzc9nQmg2kzXtnrkPPC/ZnN9CNI5FrL
J+4EsPXLYVj2FVmf9A0bAnlqStvU9ojzoJsck2c0gPTi3z6kz/4a6NBZgH2aHdcY
o6aCCOO/NkitgqXTp5Po6IE4vPw2VHboObS0u7x3RM2mnsVYTG6nx+kVZTfEwIz4
QOR4AlY17HqdGiMX9fuLMkYubYL/x6qw1IxSm9jwwh8=
`protect END_PROTECTED
