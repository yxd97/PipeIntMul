`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VD43N6tvbBbr7i/vWdrIUVT4v5fabT5UQLRQEnYN85WdFLF9mm/k54xOJt8H9m9
5oQX2J1wub89iL5Md3x1wJlR1l4xOfLi4WfpmhmQwLg7ppmeMYA1aknZf8FX5ccg
72BGi36fQncsvXMiZztV9hShknSTN1/CvghUywEyJLgfxs4UEC2irOILONj41zMt
3OmBYt0HeX3ANo3ieCKgc8u3zNhsf/pa+ac6Woyq7GRKpzfGNJpAkcDFYaECzeYy
ONV6bMbRG+Tr8HrYn50Ryg==
`protect END_PROTECTED
