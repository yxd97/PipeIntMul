`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMXztOVnA+bPIPvvBGZgizNTjLICN2ou/vDDZrOXnmEOtyc9YLEGYlKcvQJ8SNB/
9QzMLF1vUPBM9SAzA4Bq6jxXcNJBmUuZZlmuF5pBj12Tw5Z5AsWGq69AOJ5Bz0hl
82Yf+GpatP6IXZSz9ZgETpSpqsoJbu43RxEC3ePkuPLAfAwY4KwmTA8pzwkZuJWq
7Avq0d9b8RRh/dbSuHJYWc8IpIlkF1Z34UbLpzTrwzDU4YGXyvpRFT1E3M1lTyyt
Zs+Jje8kfVeTb0nrUt2vQOV3ghTgOSGEX+sQ67hD5o+PEn/a5MuX2oG1tcMBnMMV
uYxGIK/PsUZFkSWswZfVtkLFc7MG2+jYEZqYnIcLemmgWd30Jqb1EbQ5O52sqIPb
pahSY3WL+2xUnMkXLDQOD7p6i6WawlLCKGb9O+zVhNJGIj+6966t047q29oskbLt
0uyQgfoMiBPS3GBwkTxAnr52ogPeuc5Z7X1F2AcGtVSQ8lLGgCmvGLD8Iuj9YjE9
E1ImFpgZJ5B9ntJdG3HcSjGlpD5LHKrqApwxUjeQC2Ls6I9mCmmKMebnWrq0aHv3
2un3/wZiUPP1SU8A0lNVQ/dzLztN3zgeHdf9em8UNKvLXefenzhJE3qJEUB/Bc33
+RJZp/vu4YlF3u3xOG2yDLzKCOoffhKwxtCSpdssDztquUzuCfP38OdWENYmY+/s
3T0+fTL257hUNrNvzOwEfg==
`protect END_PROTECTED
