`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NtoY6xg/1Az4/I7KMlArF/0V9QlKAApn03mOOQygyC+j7oUwVk+NTGDm5huwPw7/
WVPMWCaNkPrS690o/AbONRL9MNZa2zZtrsiTyL3+e4LM6RbPGMu3lD0Kz7eUzvYi
GOEHYrd3+66mt1m/d4KaD7QmbB56izMRj5YeeKVoC4oSPT5uizTYmkKKTrZZ4+jr
s4/At8uziTIZQaR2RECn7Jq37yJnTmt8tYpByK7RTxS3nIoCT6vD4EuhaC0ao7F2
ofWAg+gtK3wVT8qeHBiieyG3nhmSm4/gS/e2MfE3IBuiL/FNTpvWuGRzuLnRPX/P
KBNMBQBPCM2vanyvOz/qokjjQenUNXvcnAGunu2YeyEv5y2RW4MAmzckc+2FlNjr
g+i8d+9agZWdqfsl+8tzTTzadLyOPEkTDb7pVMTlHznLk1iJDJDUFK9fPvOzT4bZ
nQi08l5SwT1LDd30nq31NP4HRhv5xwEYCdTTNCkZ7ghuWtZaWjnmTgGWPBEd5ADy
1Aru4APgra3ClgzuPBJDHAFi/7IpTf0mdFpokak1BJgzwxzCLC4mXVWfXso/Q51C
eQ3uK0rG0W/fYCMUiPPXEr1lQDv7EBtsx4sairWejJQ=
`protect END_PROTECTED
