`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y6YZ+7uMKu3zgEME088x9f77c12K3t49KT0hFhmiG/YXmHrU+nmkSSMRmzjDMyVR
pTA1/Wn1xGyXmVZNw51eabhBY4G66U3m/JHWuMMBabTSQKgTc1HSa2oanNfUV0nu
DtwNuBif5SXNrvb69whjpA7MJdVpnJ1QlIRF/mwiOxoJkdCjORBdXOenFU0No8ZB
04cZGa8Erctqh8m1RD5btKPM5y7kgwmJrLDHYsqceF4mA9Rcxv53XGklA5bPyVpI
LdB/k9NOKF10FIqqBprrdtKgxjUHem/JB6hilsUnWccyGeZhvcpLHq2IynnuHqVj
Cp2G3a+H1KjrOFQeec8aEyO8ZINmuGmpsIRCaHEjLYUwvxQbF0s83VZj8Rd4DqNE
tCyaWAI06lzE+r4SqlKdvw==
`protect END_PROTECTED
