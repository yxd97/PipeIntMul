`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWDy9Lgu2N+/2cSF5Ui1O2UbVjL4IsOPnYdknV2kEN9jKkFrVHbEDOLFq5g86dBw
cFHHGECvfdkWn7FTLiL0VV00WAQllQxxEsEH6y5tCEHK8Z7SprqWDjNJ6vWY5iP/
Elr6eppjSDIDH6ACS0GvQLyyl3ep0f6eyyR1iSYuP1oAPq1PWMNl3JHZBgHb3nxO
OWkMB34oo8WwRWH5mBLi04+ftxNMVaITJ9ApO2bwzzZgBHIpfopI4lje/rTqxgPw
UjUSaRqGHbTFLCIe6eyKaVg8uDNtrXX4LIt0p/4WLEmvVa4bmfU2eJYpLsNfvzkX
A8Wz+jK79lum2lbS/i2DYNktULdILWh9M7RtxP3koO6iPyrUf92D/FG2/2jF7KAP
+h2t+RCKtfvbwKshXnkH4seifu+qHmXOpD9V6Een2q+94jV6qIqls1hgOYX43zkJ
yIIruIITLNop7pjfcbGeaQ==
`protect END_PROTECTED
