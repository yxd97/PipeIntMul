`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GSTL8xnwsH4NqicokiytguqFy874KMc9xTr8L7iUa9UYwwrTd3pCUbGVGRe7gIqp
LFIyza561MeM4V+GhpIyYmlsqLJUUQQ6VwElcQTfvlyNtSGysysN9N4A7GRWsNDR
O0JNjuT9gagd8fHTeoYhNxzgrsrpJ+YIpfDyHas8bU6RwhM4AzjH1eCNa/FOo7yQ
pJ8gJhDJeOsoLQmHNbL4U6Bm1UmzgS8aAYct5J5Gel+1wHPONO/ZQBpxiBe17Tn4
GCJCuuIMitWJm1wH2qpd4AZz9xPy8Qt3WHmLWjhhBC5ZdnMkY1LHydXe8TEr78DM
6Sd02mDZJLLfBJYSQKBNp9WYSgEgnDobe0WtpplnwXocxJ/+TJ+3wBRqh0FINX8M
FSb2Anrlisx+4dok7TUQgbc8/wrdVNooUlaP9OPrVIG7LsHhqKiN6/tpxEj04TeP
JoAnGb5qg4LY3ECy+wff5DIRGfd3mDcIxnar/lj7e35VdckeWmYl6KCfD7X+97av
v7AeLCz0OnbqNc6kdgfdGgMsMWVHSAgMrI/NUD9uTkMxy8HuvWMrwOM2aDA3zILC
ssj9j9DU7kxoB24vNKWTvAm2VfKZJ0DmhQpYcvQVwtUUBRfg/VXMXOd7UNg0a83m
8lrIS/OlOP09tirT50uP4oJeyXDn7+xfPXkG2b1hvTH3Xp8/h8SGBrACrCtam6oX
0D8ZmuGrR2+boaPqCoK2E3vsxf+Z/NNI7wAgTwnt7vheNc3/UspVu36eNeNwWWVL
aCONg/WrhXP8YaUFG03hZn+xe8+gjeiR4gQTbNHKR091cWLOYC7zSSkldf8HzrFT
+6r4ppZn3Luv60W4OkGZZfb7DzF0RJ9KeGtDosfRtlC72S7ZYJ4PdxlAx6qfgTpV
A42lLhHzgugLcv9mdMCXxjDLT5LlIp4prP3H9FLZrhE2PMVkZzp0NwTqjcJIzbD5
YxCmZVDwULtQxuE+Y2hBH1MOyAEoLLdgucgbZiZvR8QcTzojIyo/6CdLAV1lhDEX
VBp1sjV4nv8XcUVzKDacb2JLSttVG12+753bHJZ9s3jekzirhiHgiDryTYtOG5Jo
AGnc8RkAVH22+yPV8Who6imOmJGEpwbiwoID+la4+BuLztXE2kEVJ5DXJay5ELIa
ur/FR+3j5+LMxzQTZbfmvJxYsBRfZezwRZBW6u6wlgNJ79mHYLEbiQfvvb5Bm3rw
q9C2ZC2nYXvvockcj7YczlT9ypWWIYpiNyTmRqm06TB9EPH7F8rU5fqQogTOD/K8
8ROJbp8EvN1ckS2fBf6qlLkXu0Y+pYsduUS6ZbYdORoafcXurz4q2Akl2sA+y6Ws
jwIRcJiMCucFIYSZgw5kH8eU8eZ03t+6c9bxkcLTTZ0lZDt3PfI7rIzuVo5WpoSm
5rPDCMwTR7wBeXoVyhSnw4pIjQh7PbeO/EYjm4KoKvHa26kBa3XM/X1R9Fvrd9NC
k5fUAqIBYZqZhuHaj0SgDqx2L1WsaRExaxjV/VXLpFhc9S8XiCebvYAa0h1wTjrJ
PAX40gAA0uMcwwEd0oSjGs5NUwKdtH0WvqiYnJdT42BoQ9XUpn2dvdaC4xyxKEg6
Osrqdo8D7z+Cq7EoJiW9Oh0MNRG1ZRT2/GuHW5yrAEYnEwSsmMT3QpQweiRX1j4o
+havcoRu65eXRassdzq6P8qNP7ZudSFiXxjWF1TaeGmxH/jnb2cIf8PST6KJRPUp
9wr2/NnCdB9XIbxg2sbrcnwK6QCe6GMp6FxHkC7tXexRbS7tDdPw52MdvToi34zd
AbuR9XppFsZFG0nuPiQetLWD7DgvPc7KmLdakz1jn3RqtjRMuajv3Wj5a4SyEzP1
pGfwI0FBGY+ev+jtG658bgCfWZq7pd/UVDNEuO1vCtzOekiJxLHIDVo4LYxrIVPN
h6gZ/p7mgSDOdmxDZXCmCmvUFWAcRQiQ1aRngvxDsc3m+HcFfoiBEf6Me1GleW19
cEc9MKU051vSwGQLieB9xRY75N6V/yvcVsdRgaog3njqrnbS1YNt8GfxjsRcjNfA
zJwTRmnVja+cWCSw26XHTj8VdcNFHn/JCkx42+r+TQdoczAhB5h3bmYJDMh9wgji
6zgXw6gZrGoR7Z1QFeE1cXij/4/zKpkGWX2aD+RbdvOiyERhy4LW1YO4C783giCk
zBidi5mox01ZVcwLYHBx2id7IP8pfhRYSdvqr650PImSlzZGxbVJ1nfVaQzdQFkr
RYO9R6/JbHOeHfyZLDmUyQK9swODuRUPrTDWut4EWvdMGliCwixRDjme9o/VNeA4
jayw+OyiYl3osF347oQyOY16F2vf6GhZ63fK+RNdD9JsynOjmIRUwOLKmx2QgSYH
zWvnD1RQQ2RMUD+pwqdHXenlemxlHqRTrhatTSSndWXpM/VGu5XRjqV8aTd3h7sv
O2gmwb1JoURgpSCMLxIPFDr7ubSAPCjM0p3CNNereU1BEclbOKVwxhj157RK6XBl
6NObq0+fCBfpNd4ceSAMCU8Nhm73856kKDJdqYZ8fVP9XBg0neaT7ujedNf1nz4c
XjftGJCc8DxkXbbih/+dB2p9aywxg5RzEKaOYgDV5gid/W1rbRBZfO/1pwvpnkkv
kTdBiMyAOnbqvRwGkeDxmAk9ejj0t0tFivDzLPDKUYmI1XzIK4zr+z3pDgg9SrnR
IkCfpfwgQJbHn0rMId1UBk/o/3JYsU+U39IUCNOpowBVEMbDIP42Zpfs11DXjJbw
pCa2Ey1epHa9nxSl/2y0/uEp3dLZlAV9HLdXszGVFq48dFv4Tn9hcHCm2A9KrZdU
uAl9sDBWwPA/Y0PUSmddqWeiyD/dO8DZ58P7ZdyjV7x1lUbial+tGhYGOKcQo+1W
AXZ4iT29DvNvBJsOUmyMCImL5h6eHqrC8I2JjCEjEkVqtwvd9dqDCC9W0dqqefZn
TpVwGls6WAkJL+n15pdZJJDYFhMLlZO7zppx7hE+WR8LnIOaW7IF9WeFBujKFYOX
ecKgVq7Lq+w+uWWr0HqL4ujvXlUmUZcu2MQHUZlcfkm8a3zrGutnUgE8N/DOjmnc
bBEQpqJ0XG+UugzQYEuEMXXt6XSINleAQND5r/MK2M57uK3JTdIRRsUJR60g1uEF
bB65jHzNIF8aTHh+Y3oDmcsm+dx32o/ZVCBvZ4L09WxNYFUdXrN5u36rymT1/l/e
R/uUbHn/y1c/IZvDJ+fEAEm8FkbXEqb4cXJvJ6CnyyPnsSqkdrckMjjL39gxXqIB
NrpyYwDDRpvZR9D+hC3l8IL9+FooG9876FI/n/5xeXymdRS52IkQuXNYJgZGgu9s
Eji60l9I7uBS+QJv9GGRuVxGQpK3aMaAIBRnDmHvB3ZtITH4489SYhOkZ8zFYC5V
ui24ST8fWa3KcYFQUaxmicoJWFouLXZhYCuFdHFoNMy2wX0nZLiDT8XNuESBcLOK
9Yn9f+WXYFHs8u0wEivZS5Bje+aPS5CfHhzxRbnM/26bkuNBgBVGLMVMnXE8rG7B
9/VJ02X0sUBw/jCdZA/XZRtImoBohzmHdlhNjBR8ztfN6OA2wXQikD8eQHdYxyT4
/x6sLXCMIc1K0IY0pH1Uf1vCf7tHlV6htMJll0k1UcM1Uet3CykiRyVL/yEh9gE9
UDuAbGGc+CilFBPlfom+XOifBCgxiIOarTCxJE8wyVMM03JEHionoWRhZSWwboFY
Tz5r1hULr6UC4ikU6RSmsounD4DioRkGqn7N3UT7F9xdTTjYnQmDxOCBQeL/qI4x
tOXqmTJk9fQ3eobgHcdi0a+oOvfbiblDjfL6pPxP+KgUNAw5gc7OhQPXoeYnuAL0
FfxgR7ZfQ8Kp1gM7h35B5BEncG3Mj7FcRNoxZPeZizg1PWB22msehzBccGTVgQlI
JqJd7YdKsOI0KKp+UgNAFLUh/Px1WdGF76zmnNI2Q0VEOlixvFg/RN0/wY4pKoDK
/qTU93+R7ekvK286oJJ0WeUSqUiZMJiUs71x0qP/SKHFGERPc0KBuPs1I4zFYAxx
WOwOVIZrE8eQTVLGSTpTKK5+jYrz3J0UCpHJTZz8NwrOb9J76YTlORB0bS9639HQ
d1C6RUqFdFerGawYjJ+DUdg6cdLT25D2+cKrb6AauAELAONFbaW3LA20eDkxRgE1
1im6ClAWdeqUhF1nxoJzPRbvgPuobGWqF7UAh2Qejyx3h8W/QnAZu86baT3o03eG
`protect END_PROTECTED
