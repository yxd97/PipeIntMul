`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyDLa8iqX6ZU1ftK5xhviRC7R97XvgMzkOsZDHlaStiGQF4+vOeuMdvW2M+qP1sK
wcJtAyg/hnUTARKzkvyqSEGEr7W3Q5g7wOQYk4DAct4Jl2pTUdX+Ln7d77ZlQdBD
MwiYDswnLDx3L0x595Wf5V8ljD48sgvJeveOBR8Poy5qpuBbnAH2IdP8BygzVcub
OtkUus5nowBzX1f8AG+6uWeEH6ZJ3m8OwSytn0cGtG9QVvUFBgJvqu9pPhD1RYyJ
c2N/MPWn+vzfUqM3pCFTkLjCBRtvOv2/KuGXZyo2lpfxsErIZo7LVoU0oGIUWxSQ
75OVo1lVSbuhbZjaEkA6UvlJdwK6yHXgy9fxTnToUjacsGBLPhCTag9Co+G31Ig9
l8HJFplc6JkV+0gFlw/PX+e8X8eDwENHkMQ6Li2TkBb0X8FPYFGU+oT9UmMCf0ET
Ozt8hyUwkimGFFVqOCRcFO9pZG9DgnEMDtagG0eQxWzPCIQjG8K/FgrWSA5D398e
usCcaW+bNRHXV1TpR+P3t3IPWENOYThncZKeIRu/hVffoDIIsAyq9GgZImM84N74
fhNNO9/CoZVdcsr7dd1M3rAxJcUpECfsODaaODF6GDiOJyvWuRZMRNqivIiJs/PW
n/fVQvRfNdeF/D+MmzyikFc8La/tvED2VgoBUwkAZ2FfXeFPTfmxw70xQaUglrIA
RcfHo6pLbvA723iouDJVC4tbiBJ8OUvkNeCmIUHLc80DowqAdK4xY9LZA2rAwxK5
SZjhkPx05pF0zQDjYg9RueyvXvOLpRcLfxl/iqwlbbC8XL7Htdwrs/RG9WEVJ8O1
c9EJJ3+6Y3BzobAKHK+Z2gMJTi4KisN4gcgnGLqQdhPC6wHws1NC1zmT0d/fHzPh
VehLWet1FjjbdqgDNBDZYus7HUxs9rsBd1o9MNAfYWmqbp7/1rw5Cj6hCtZYtQYE
iQG2RwrkGUisJiIQl+Mj1/YKSRAat6wDHMv6EH2WKdNL0LCSKWplS89MBfyruxyI
eeV2BRbkQ6U8XyyGFY65CZ8A08RPxztqijs/lLfGvZEn1DF6l9xPalnLAQBrvWHA
ozBVMhka09uwubmEqid+uV9dbTLtBnEEbJNtYGs1PKrk5UPsiC1EqzNsBIILa/nG
KFiMJzYzvLm+0MCYR6LWA7NvEFn0emuDe0J8HIHpogefp775pIRxetctQWvcp6hm
jGpSsTBQlqFRzmrtJCrLOTaHNL8XKxcp0B9DfODKtSzMPrNjoDmssGSdrIafKxhC
C2glDYPSVOa+GiZyXtg6y79/zs4O8ja0qnTYaPCfPTSy3LDCBDWU49rrQ8XSQhxx
CWT5iKRQh4/2TgRfvo0o3EqLgPWs3dYjyrfHwvMNV7KTFzchWt0EFCI7Y4n9ZkLo
dPIibeCkXTmCvL6jreEY69cPuF8lfn0n9HjQO1efIx58QA8DE80KyMR4mYQ9HzyN
qWlTWbnN3ZKe3TA5w96YuN9GwpwmYn3WvtL7rg5w7kB9N9k7E9I1O3ox+0kR+n+/
TuQ/DUirCQI05X1ztax9Snh3PD7vUrwYJVnvfytNHl9cOsSmF99efYfYnr7vK4Wz
DUh5L4xa1gte4+A4dAXMH5RKJIcq/0UfoeSI0ArnayQlBOICy+byoK9IJJGVSWJR
io9/0QyYKnaEHib5phfQnS88wn/hFmHdQLyE1LZww6+f2lPJG8t3jZ9IB+ubCzDM
x6U/S32f4yG2XD8OJPYGvmZph3vzWJLsEdS3Ythg2pxJoLisA27nj3bi8Kl/MiIM
kESCi4aWz9iS3iowWvH0TEVR9AobFKlP46VGLruIw9PMDn/0jUwgIBUule3VRv6X
N6rq2r9B5BcBPXwoudqtZYJsKuY0bjO5/paGUVQra+QTPgj/R7sckd8906vndUoZ
vJS/qOjkE9fjQYA6fDzOEm4Q86SLYLooG6YD04ULP1hvuCoqfmYK4g7MEDIfezVF
Jm8Vyddsa+BHgKeMAab9c+mqIjyyf65MXZv8zNFBdvbXqFqhZIg/LQ92K3LAHq8m
qql40FCG9oFmojYTtxK2gQJCHVz0rZJchBbPgySwzVX7HUewv767U9d2pEcIpEdX
dnXIMhUPD3nyitL2UR6wlF0uJjGReewq+D3GdUjahrLVtCs5vKHIyGc8bhsA0D92
D1qawBrxOj/6qe+duFodYvYTYk/aNVTpoBTyps/r9DKq+6DINvaAye+PAvVWDvYn
+c9X2CG7do/q+oCNnOknq14rbKvMar+gE+QjfCVdsVr+DHNNMp8DPwJaZ+v7Od2s
tzuid9GFJUr6YiiyrGXLfEcOJ5Lz6ei1ybfUYWWQAE6S022WEXdwv28HDHPgjOcX
tbEo4oefKRKDJZqLTQrTqNCPu2Jmvq2wgdcZxMvPYV6wVJR8xGP6P3kOiIJtJZLU
DHbg3gKzpmZ5hT7KYKWROP2IEqtq4YaF+uRAhg/KPwX39ntorQ20nFfvCbAdJgPg
UQ1+zFrkMnxx4cahrzMvI0kBkD+CAV05UTM4T4os6GrIGKuTgvIz5f8CCFL34JBp
xUW/h3EOFENrpDeSF3dkE2BphW9oz415Wwa41m8IxX+TxOJKwo3BX8PpGvFCYeHT
mEBzvLSCpxb/DJDzkc8y7ACV+ALJPXA/YbYxopIlMXp0pWj9PXPm5/EC/MgaQsSx
6/dJHrn9Kz9RR5W+n3wj1PAId2bBC+BqV2qRUst+1/rR52n4cfl4tyIgFx3MLrRY
OgI+m5cdeQlUo95PWAH93rJqEik5k83Qo2ZnYof4E/n5jUJufwAjPQavof33dngy
i8trGEdxPPCTILVPuS4eXE1YiB0Jkd3XxuwLlbQaXDVFnY9ksEJLbe9ZhLO0QXhq
sy9KK/Bszn7B5dgeNQHEbxAusj1xyQe5cPRzAmoxiukydJF1LT0vl6Nu30zOsbof
E+n5xTF5jMIt1WTRarT3D9mHMxMws6FBRLCzeab/LX2cwoloTIWdnc8xoI0J75HW
UNDT78rxIVDMYr5zqEljDnVFSOdCIt1nTvq72bwgF68n1YzlvIPM86X6Aj27BJX4
L7Ls+PL3uSXlzgptok8H7InvmVJplqJPlLdRqx3ghVCoY6xyXCmemgfb4fAUj/wc
CeXKOXb31jzzQcdVswgA1DOZh2OpS9GVq6gjXCBQWmBG+6dGVmSsqAsUwmFF7gT5
JfAKyhPhN3TT7iTkmAwzzI5eEQr60gwc2CgdMukHDk0QWTVelfGHKBYEFT8Ea3Pr
tR35ztk4/LRPFjLX92KUNjAuTOi3rhSXmGEDpF598qugCAXdvC1tnJXXQORoiq8R
RuVoqMhLNIGFYF2SfpdauBhCCKqKRCRwiVdIyhWv/hTTVIGmlbsduR70e3KEtQlE
E+2UTbl9oFrFoN7vRUD1k4UGAj9I7Az15wJIc+qyk+RME0plg8xD8T37AloBGZOP
SWIsA4FAOKm+VbY3IYZYfKhKdyUmKy/G86JI+aLXMULfPzah/fxo5WIKvOozOLg6
u62krnk17ot2E/mooWwZuz0LGsxccrt8dv5ZknL/kLg4ZV8vDuyNJvwDDtyt+tcC
JhiGDlPtxydC5n2tXrmbvBx3bApWBY7mVkV/N64xR+2K0Fp+9sZMG4R+0a+oO4in
NfSyabwmcWZ+JeqDdKFBgYaQHhV879gsqcpYeAAYQGTDKwCfhHwYPE92IQNHuBGi
rkQzRl7WYzS9PfS0EqzSbFkRFIIUCQAER6sroXWQWFEznbk4gwaRNdGXKOkp8cGg
P1mXLYQvqaQNbkTzRWI1AnQFFXPu0dWz4jkvzmJhhtg1MAbeShTt+4QaRnZBZWHU
NTiIyEDXxNP2mQtzexJocSm9mFnY7KYKKJwacsGmWAzkqYb+HkaMu7yTmT6mciMt
C/wj1c5EQUTFQWzKLlKun7zZtI4ZqmqIE3QFVuBXcMGdS2BK8ljXsqXtMY35uAET
WB1UmfeplyM9wQxhDSRWslfu5GoisgnWNFrlpF3KQjOQL/3J2qVc+8bwi7mDZY6u
+ZyvbEVrtjFbMPsPcFmJ4IyEwpkLF4Uzbtuv2Lt9a+GPdWwWqUT1BLXwimOYKNIC
F746Od0YwKcg750tEo6MHgDKft5fC3J4UbVtRgTIlmLbdyoecZNhrbVYyEtG6dSG
l5FgMZ7z2Bk1bD068BA4pwqXJNizxpVTRlHzJyevmkHpr/MWzEwTesE+HX1JZLqY
PqVsA3grFWOcYYqdVV5uVip61McezAdfOsgWYWx/y2rcjoHFDYDBC85kG/8di8dT
wObQYzLfU4JaUHDVpY7ey1n7cNFaW4rN9kiizli6ZGo0X+MmDWYuhGUCuwR9A1lM
YcDbh5M1MEjN2ow+8WVNi5kVBShfA+JdKXWFJDMWvjt68K4TPkfu97WcDXf0cuMc
E6geNmJadWYmoTNthwOUSMpND9mllZnxKDgdq6KLX3DzVxE2nR4ummD6UBipPFl2
qg770fK/LNS3OQbV11eIcyBlABUKXrr/qEsyY3iHOdZspv+bvtNDvpnhP07dnB+E
C0a/cW1ZrNf4J8WSAwdF1EZgUM3wAUpJNYak7NPLks2OQFrlATMFqx92aV0VVEaw
qM8Nl1ggnstL+L356SPMOUDidpIhnjV6P5vQaQIlMmOM4KCWI4i+FhplG3H0K1ih
tXhSrKYX2WVNj6NGSnsmbd65y2sLXATR8GqA03bbUMFE6YOxuoeH//nEV1k0Afu8
lDDano9DLGPdA7xBxupxRPAX+J/oQ1+PsWGX3KIQoWjG2Xc2d7FId3IfiiO2RoU6
TiUfRNro7gDSnqF1u0lLoGzkXC8bsv54jZOAm65hu9530eLZx//tZpb2T7V28S/I
k6PtmuoFRt+CcetZqAmDjmTN0Hz7wOGtA5kvPVZtHiQfMybEHrrt7ppbfadNGKk9
2ef95diJgvHzQs+iQcvy/USCv+0UeZRNzucA4Kv67La3DM7+NiNatnR9dd8mJEzm
39vmYnEgWlrIBjYixf4pHFhRDck75PrVSJw++rXGTO0cfQUxbE78pvBrk77E+0hh
bOk/K4xcttixG3vmyz2j3/zmZ/0UK9//BM9aku0UZYZa/jItXwKaraagslw74IFo
8a+EiWL2NP3nMVJwUBRtTx2APQ5o4OlRsE5vyGDLvj0HjaPaIyRk+/oz0WVhE9SG
a+a42+QkpUULWY22l+PFgX/5dgHoeatTVkXb2suNOSayg7IeG1THcM9hmcnXFBW8
DLj5c0LJfa6NMJyO/6TrjumnPdJlTy6AKA7dKIjUrj84g+uRluQi9Ul4EXiE7yLn
jp0zZ15IKBzJJ8RTPGHB7A8jTT5R0OomFM+GV/Jv3c4fLJWOUA5wKzPzkcBiJ+g5
hT73Bvb4z68XNXRmVHtaGr+VICFc4czZa/NnhJJbLrLaza+sgpZ/Nglgnmvg2U/4
k45sZ3peqhJulLw0Z4lorGq/goqE4Cq7FSoIuOq0EuhiTwrgjksLFyROKYo2qZxp
ZdeyI3sHBNrlUhYc2y1slOC47qtFQTC+8NqhMGiqZZzzOxHSkdoHUPkvgEtGgtJb
MFtAu9KNrPWRZ8PBHGZ/FP7oGCbynj01FAktqq8+mv3biQPLZKDbtUL9WkXMoPyI
cVidE1k4lo8FRc6TbizNHE4iN2OwuErvU+hBHDFhPryeTZ9UAN8bC4CmNFz2H1H5
Lf2e7KsnP/4TWaY9B+6mIC49TJSPC15wOlFnRPm4iCi5TkqhwsCUo3VHecc8h1ZK
KFQhshFLm5J7XOPnC7YeALPK0aSGd8JOxXXHft86oKlSTxCyOaMRnPbPxyrGK3K/
jEZ4FO3aYmSfiQLby7iIi6sz1xMROUGAv5lQEiTtQXKg27DtoIFO32pMfiEtgMlu
q46txKH2fptgPTX2vQF2cDvm113Job4WxLU+/Y20yE6O+PSZ2VEXZQptJmoruNrA
3o3hBOiahcilzdPIx2KEBduwuOEEBXKoLdvgX2zf4JNfRaMK43TpSbe491O9SPKn
OYGi0fKGEmXfO8crWXfXGjyKUUhGCnxxEJ5FR+slgoxUtbnJNJt8A6geIojEWhe1
fb9+z32zhcXqgbItczmLN4RiJdkt8VVyR5O5r603X5zM/F1eSLiCjjJ/sFCgRozK
LHSKOpga4HNOX4kVBaZzlMJftVD5Jc6uYogXXeih++jBIDhKADBqTDU/PhpmrbZl
X3DI0S+8GOhskpoVEAuFoMm9ca1apKLo6RIzEzNqSj3aIjQohFC2TxqlLuwCymK5
aLWtvwcN4D7LrxnRALLj3PFPPdOMWBcw0aisAYnIXtaENRLPKhu6NtJrqjiuknuo
iDxn2HsLL/hrTeKJ5iPhwXSf+DBoiGWOtUnEtZLV7F1hGfdTc0fQrzsOlZ4vDB+2
KiMyeDbWXWwbkN4FJu6iz7cZ0ZdHSHojbOIba79b6VfKFw0Gs+QUwPWAkAkp+ulZ
x/cCYQsjlagL+XkO2ab3k7iVmZ9j8DhQm9WROtaLKtswZEQdpy/DgEvI8eKNBgHv
jmIIMRAvHtmWgxJMNLlJJMemvrHiw2CTceXUxS4wB/WdujzkVRn2VvLwDaAHDr2Z
RKGuLtN8qn2ap5waFIJdwIRM/R6VtBqEAudl7tjLgkR3i5lTgjjA44+ybUop6AqU
lccZyHDqkWUhsCP7EN2oWK/fheLVyJLPPgkTHh/fBmAw+hnGfPeVCyG9oN7KKx3Y
rEnZEWhfD0b/MA7s/evRHIu8Y8j73bYyNeOXUi7/aKzH75UIsG+1CHDXAUNWCwVc
uayPTVOAhxSR6FyHah3KYT1/6FpEm8TEI1gmTq0aB4ycIRN2bni4n4tWPy2EMvsl
ay4eqiVaLbEb5CIhABRcuaaMghtgK+JMjvjn0JC3N2Fa3eGkpOtQpNqzpEnh8hB3
BnY4rspEzv6mZLPmD7PbS5l3vre7vzhN6aHVYc6WFx0DJV4m6/5k0pz+rb4lMsBT
B+YNYtUp/bGedYzyjR3m6CP6i3590WG95jIESaoMFSOECaws5FomiXgspEywrfHl
B7U4ET0PBXIviJ8/WVQAdahF6T6x8mU1s5TTw811IF1yCdAK21rrdZ4FpVxtKxxp
T1FB/zQixnzTSnRFuPd+VBu9QWGJsb+2ZIPCPZXFTPbFGbnJsuUDo4/fDJ4oFgAZ
QXLTXhW18Cj015wHKK8b0+rpieRA3wxdBbXZpPLr8QQXkUaAnSZc77FKFMDKCQ7F
Pe+PZp2uqr9OmJRKOf0+3Y8zyw4V0pI9DPyccPxggOvfFns4iwHdnVVevfsQy0pc
JDx2gxO/3vAruObWsKWeRlMFDAUbXlSN3+z/Z7HsOzr0p2LJKfvHYIpAmIIt6RYu
RH1tOPToFY4/oslf66YRxN3MjZR+l9oJ8rv8Hu+Jv7Ym21UEt1psTIVtvx1FnWd6
2KAiWWDvZKhbYJyrcco80phJy1ojfzuvYdO6QC9C8nyUK5Nm2kcbwk+hqJ8KgjFZ
TJw8vr3nLuin77bnHujbAiuCCIdgqvyEQ2kFZMigR0E3wxEVx6NQYc7ZWs+Uv6e3
oE6F7aR8wclrWT8VVGhV8GFVpu0fEbQXLG63NaIPda40+NX3NnU+8QxRVILjusB7
BxY7MQBPwLFUiN0RZseIQVPzowJG9Jr4GFpOe0jogDWkijY3/1rN+kGkOB/lW/q/
k4EVZUL406Dq+em3c4pNaHoGaw0vF2PYEUzwIOiMf0hbgafg3LTT7rrDxEAZXsfu
ZFKDSqAH3hCDKsaNNg+pWyc/0c/b/a1VnBVvknnTEiCH+WSs0P3ntzG9GK+h9gha
McyNp/I5ukNkfXjbyI0HGXq1QwoIWgrrJOSJRfzPBTOb16fUlHIvqsF75/ZKcfne
yKvP1XImbvXJJeE+Znyja914O+VrV+OjrrpTsyxiT1DH0otsEShh0hdBv6/wWmWa
ntFqe+BKhNdEcGbHHn+bGUoKPkX5kNswrMtZOnBC1KcQIJNQyqQk9SkQxZCuXcIX
AwPeRucJN80bvIHxsIq4UPBDJfHwhmbioxQ2H+xD7vvebvUhixA4F9dqaSwNzP0b
Eb6UTlgBp4XsudSWYY+6ChYH5/eLOoPebhSOiMTKS+aiTHHDkXfCWA00TypyPInJ
tAPnEP81pbCB0kqYmw686+UtRfkkVSOJ/lXF/4V2LLkh4OwytkZYO/T+gys6hTEh
duvxtyt09lEyEvfO7PvB4gf3sGt/PEwKLpAaRFn7+wjFc46VYAiocOM7YHSLwN//
JNLERH+WzOdwc/UxJJZfkBy0cKUPoeaQOCsRroFOZX8O2osfSF+9NfRd5LExAFWa
wOwo7kTe13XKt+31z6VUDqyeGkGv83imRiCxoQidTUB7tnsYcVDeiLvDzKJ+BFGC
13DqjZyxF6fKq8+rTuFmjpPv6CbYXmp13AbrACFD+AS32RpwWT5S8ww/jyaycW0/
EBrSr1MWXeUrXhlPeMM4MeCPSwNhyHx27pcg5LajF28DgDG1ezUIdY5HN+TnMbmn
J/P2D0YwvMZtieSQJy8AW/LI1Oeg5VKA7C1anA8yuKj7DYQyoW9+d6TIIIJegWVG
oMKsSvRyid3mHBi0ErADYTbVYTt+6d3q1msoaOyCH4jwId1GWoxK5pTuCZG9SuY0
YiekhvbuDlnPI4SLpj90BDqg4QPHv6O+eejbg4lUEPAEx2E/B89D7wyyCnL0+za0
yY3LtGqYINMggwx57RAAsPQoAReggbO582QqZ4GtZUxB35I6W/dpFBcszI2rcqZE
youPngav5Ry51Zcomr80Nh7L4RZ2JmX2SC6oWSW9c4S1BlH7C4ylowBYFE8vBrGb
NAfAbux/alpwQlmumIyTlE7VEhro19kOm4Bz6PJU92aWz0/DBwEwJUYTyUoJBD1x
Dg6EK0eWMYwYUd1JXcHzEUSZ7kTBlw98rYcblP3Zg0s0/pxht1Hh2IKie4b6Xz3q
q8WlWcuyX+pEu545I9oM8+XhvT07sWxNe6nn8ES0Q9H+xGpxvR0UKx4Xuh83yW8i
DtO4K4iujvjfhI/cVgmifUEsmsr+RnRPKOyM9JeU86y7N8r0T+ZemIjSXcjTrZaq
wXONGmm7I0pR/3Cr49kUWKO2XVhMzcB/kCVgpmxCoBaU3eMB0fVnqYx3WZNeT18j
QTebPM8iBxFqzm7HoQCoB2ubloGSo4rEYnj18m4ewnFSmTF5G+bjNhxifP0n2Lcc
vsO6qX8LgWhIQL39IvezE5IigCE75UZMalcFAhJdqWavZexGG4+YtxGLQg4bNuw5
NeHbd9EerHA27l6Zl34J384EZxk9e3IfhbpI4jYyE6D+FZhNfB25MFQ+5eQUHCl5
XB6eZczsQhkmyRnPOKL/Cq0PQ1tCAgUr1cVeRS+YCkikQTGofRNizy4NCfqXyB8d
yy9b9kCoF6THUtOcp8rxgzydR72S2HCrXPDxpzYEWui5ITsBsvo+GeNvFKGzsHmw
nQcohlKFrWQK7U4/ZcyrXtpN2XYlGs4DNeMvx4M72nf1Cu4Hrdr4kcjSrV6m0Hh6
QKcLnYYg5LQeMVEDbR3k359ScShyw4GFUr4xlKai898RmhBTUVjM3eBXlpMXzWGo
gRPlGSkYKP46pXl2XesOq+6F26i7Owvb6YwV6LzXfyUuyi11J3ai3VMveEXei9V6
PZQ1JhkoY+5Nq93t7oC7bmnm6Tx3vNcy8HnFrI93k1qdG1ejQ+dZgzoucq+mZb+E
AGqBjWPs9O/SNwZzV2Hc0Q8PXsA1uFylEOaju2d3ZSblzsk55SgVjxrMmzx9/f7p
Hknf7BLWmF6QxQZubT9bPVcjF199KXYWhE9JPA8Q+ztv4aHlWKJ4vB0QMYvBL6pP
KPxi5zbECdM1bNvGCrH1FJIq3dE2HaTixa3gMRBWnOt3496DjQIkd0tA/nR/q07d
oaFJATaY2eXq6M+Nk7XCxDuTEvMScMvu0WSSHjEmUeyTpZQZkSMWxhqUnKEWUKsN
GXFVdnusqwgMKrq/Y7U7SWQjx+MPY6UK5MyoXEl9omCXHimsV63P8R4Rei1ICNJ1
IF7co65P6T/rD623djb7ZSJp6ioRPUeHUDdo4fbXpqNLVtrfI5nDIzy4UmBsm9mn
Zzqlm8LRSL9/JIh/BFgONMPrLhlxPNABX6fVfdZ8ZBKpCX3l66E0Gs+iva1EGsy3
yw15CkPqSrnYjLNXL77cHcGwby8MKok7qr5v3qWoj0GR1laxp+fKCpF+js/t13Yd
bGiTGxJ4bCAG9Z56cI6/awX1hK+9EiSGXh/q03DEhVMNVcIK7W5JemuzvqJFcYa+
QMhx4S0ywwqjz1cMc9gHm036hKutxl9YqRLNA+6NjWjyrPGr/AqgJCde9K4ZAm3o
jQJ49Rvj+e4EEyfrw/SXUxlc/AnMJWztIb76c/iGsNHYHxjOK/gO4bCdKhNp2tdx
edrht0uuDkotDN/UjBa9hj+h0QjFHNbSlQRMCNP/LFcB8fCT7icnAfkc/doN/VPF
LRwy2VQ2UsUBTg6LCiLkpNq2F2xndpT76h1hP8TXTf3PixUR73l+ZuzV59BVF+Ox
KMOsK2UYJ6KDt6KTtFsONfitx/eIBFVN2x+0IJCSoHWocYrsTEZs5bRPq8MjRw5O
7zdAuQk0Z9KiVCFK5q1NG1Y6IcEMa+l4nIgnvxFaD5S9QrqAafK5x+VmTYCgmNDj
j30haSDnfcu0GTkk7qJHm3RBAWHQ8v8Y8yjKdvz7a4nQefLBBXAWQqZS3i1o1Soz
8gbytVF2uTrcufF05mmpZz3OOgStrLmbchC9uGaSj2ZAOy21e/BWY2IC2O/1Ya7N
FE4ZO+jJnFYUtpBnzhRXqoDL5AyPgoYotHNAGXClfj58qs0lUcWjjBEYgFevLAg2
na8e8ihgXmMnPtmv2MEt5wiA8xppugsH9kLjwSyhmnKPoJE2oJYPz6ERrEJtH+Rj
DppHpX7EzzYLqBtGB0LTeKtHvU5oy4Bx09UaS6XFLVU0EDm32Tsg65HPO0lnKTz0
54CgO/TxnhVXe54mbKiuFUTJx55sUacUWgwp5FsSxOrqySU6fXAilfayq55aWl2F
s2ATeYWj9RazjFT+zYLeZup2rkqj/gVLLIIINWKQcUHVvXLy/7AWttLbh8kXSu9/
Upf+lZOkp1eIc4sceVFS5QFmDcBeb42mWyyaW9cvXqzxno+bG5Rbsmat2RyGaceh
qI7bbe5wUj0Btiv6tYojv7sE4s/cIk1D4jsWXh+3L84kexzqHN2qTZNDmwMzAE+u
su3qAQoAEtL6kFpuRfkpZ/7ja7kX0bdgTCSboWBJhd+Qhadi1RwOp7LEs35CtGU3
vAmlcRTIQghS/xa18T4ffomBcfJfAgNNbgPhGTxGiprp/vxLB58hmvUUuK5hx9xp
NfwuUvqILOvEy1JnHsKuzbPJ/zayekmNoUmIkWlo4E9/PHM5GgHfnJ5qhIappQcJ
pIXxyVta42UCyg1A5fRADD5BLXIhcNiRz1rDHwVp2w6oPOo+4M8t/oCeLXeK8RU+
y3W36LRaQpmS0zaXVEszrzdgQ8PwdCtF7KMy90D/xlliVkEe5lFTGoSFPreBgv0f
/Vp7rrn2sg+/5HmoYamr8uRO+QnkjoyobRohXxOsuv1+QZMqiaZ6GhckZ4uknXgm
Tq7tYEOorxHfsc90tEvsM4Kt4KM45+H38IkczAiT6ARMcKusPjtmV9UT9d+LJyo8
hNWP8WpONznl99cLb5i6P4GHSACGeoPfbQHoKrEWmJUKlaSTITI35gRJE7+ARFCr
QBhqPAvLQH3Y7WtmifoGASdx5Ew48kXRkuvSUAfRPZSXnIKC8A1KginceElhSbH7
RKV/eYSPama8UGj3Yv9G4hmVd2tl1LUgbc011p6iYAu5cBYRSUm+tpI5eV2PGjjI
edi/PLDxlPRSerfbjnH4j+LnF/Df5ZIswynZgk0h+M/CDTPnY9eFYu2MtDTVH80Y
bcQcqVfJfmze3idk8wZaW8o0OY8n4YG4j7z/0sJkns/c7h+2NHT6FoN3zq5gSrzd
qDyMbA+YbShIrXp7Zw39n88GEmpj41jhC811ZW3ylN65eBSz2ic9pr1C615hVIGM
yqldvVszJbWduYgSti2ikODzePSuUFqLoyYUpo7Kk6M8FXRls+xtTQUCk1VGZuL2
++apolznUj6UNO6FMcmprL/+fWy4IKFQ9xXefEuRlW5hoSCLqePYGu50H1LmmXAu
dPHGOzdEIlRwECJQCJO8THd4wCb1T9wmuz0bLlS5E7FOsDD75Ct6mUiTMnhZRvFQ
j6mnI7P/7o9JSH46y9elgGEPLJ/iELhY66cDzd/muqb6SM4OhBiCnBh2FSH/7aVz
GC0k3wR4qhBkxgSqM+nJkV9TJTIk4bUPhP1bSvX4nMeRFB9tyeiGjCglxIapls3m
iygnYxOsNW1Afwi3QOdPRN6p4vo4ROcL8lc80/KhhGdX3Eg5mxX2eGfiLyN5aeOV
Bw2Ns5Bc0t4H0thqvyk1MmVRN6G8JS9uNzj69oHHWE0pbGPj8W1DeQKrV90q+40Q
n1ypeVA6TIBGN2xscOdpgf2J4b+f6ASamDeMLw3/pwyqReegwmrcXqq4F4SgjTID
xLCbg03DLVk5l2+TmAMtubGE4iaRB456nkOLaG+tTiiQ6nzRaT12ukA8d5HSmg5o
Np1gx6dFFtHtjuKTF2whYJueRi+Hd2I+BvBaxkVC+WqybdUSWgzRyaOSFFmxc2HF
s+hqW5E6o+A+blPy8WbRj8FO7Qz5BcJoFxL+mnwPzNWlopR7820sF8tHcBjeqPdt
Eh93y8JSynPZB7YYHytgxwFnmvCSCVTLq6c8Zs5wEm6riTk61cRcnnRrQm0/96FL
C6TpvnTN4P1b73mre5ebxXZDz1AqzDxpatC2meyP+6DqGO9hO8lmp7Q6BtNt+eGD
9bb6w1Y8HSNenpdCafjD4rNL5FtVlrdhx9RJTZRFUnlzevub3IpSEudlfrfZi9GD
SzOi54aGpI7MHEQVcZGmzxeo2ywjGQQPDPbWEAHAbXDfu/cTOpp2MuSgW1tbR2jA
0yaVjfQAbQSVenuBCOllGGLQV1OiL1PCBI9kHgsMn0up2XmfSvVa1QWgVtQocyEU
FLz0j7DcwoEwjnKJ4SIObIbWFiG8qkdCkXEz9JBI3wdehb+2uhcs6D6vyU5a0ypn
G457yOGdY/lpIwcdnnG01xjlWHTGp+8onlOQ8omPevrcBBLX8p8K6kiClwmfF2Jf
iQSUXjUVwz6wbqAc0kvAYRyeLHuuk2Qs1kWjx5lQzdSvRPl79GnsBdeZ7dPLKPpi
QQSFTiToYcjm4Y7XqqZjqy8OXJktpEldpRa28XIjyAYZeqIl4fxh8DUWzk3YvkBb
Y5COwg5ejV9PNE0YGyP/CyDjFJVAt/FnxNcYvGo14iFqwZPQLNz/oCR0F8OzZ69i
1lqbX3pV7czWw9+BSYhA0lwa2+SJTTtto3zEo2e0XVSqZHA+2QyhhyeXaYwfHDQE
be0Xw17wnSQxCG88Nww2XvN0OeBARzTH5n2DdwvJ1aJB0bRcOVKaXjeRmwsXhfn4
5tOK4U+nNFlszIgydZtOicnWvSELX4t6eSHVGby+A5tP5FWbcGdYrInYHc2JhJTK
hgfF21SkIHIdEV3tosvostZH9y0xRvg56TE5uXa3D0g8IP/l085f+c9Vd3QgHvcw
ugW1Ce/vHNr7/973snEVK+C4+kdXrHEbswpvZI6BEf8sqfCh29sm5S3uSTLptEiX
hCpfTwRMLmnsh8TZ8eCePtUjt4s22cAH+WUxGq4Sy7EZi1dFySc9jBCTgp1U3whZ
9joexIElSJjtRdrxnPeadj1Pmiw+vAO0mObhVaeJMO4zWwwuijleMsPAbHMiN5AR
oeEYtnz0BmIvHv1+fpFzer7QxEs24aF9VbZ3tboH2Rr0St6C1ItMfYSsjFLrw/MR
tEwB7lWOhSqNvaFdb6JQhscXjQc/Cx64mWru/NELIYDKS2Una+XVkbHip1wpa4JM
K59hwhU/aUbymThDKcZypqUm1I8GqGdQfNgp7ok68jlY1ML2WHL0A51SXPp5i9wM
xO7LG6hV/2og01XF2zOebbGG+3ZlpOe0Uw1/AXK7RDdEX65taBkxLQCxEtLXkiY2
6UnEuZ/n3fHVSQ5bi6DtLvCcpVOhzQF+bGiwOpE8Bofjn6mnWUQmcNY+tXKh0r4O
yxOsMWOxGlUZUEE/IsInpPYCDh3f5umT3WH8lijbZwPN+Kuqc6hNXilLPAC69FIc
s7ivGar7geC7chMDtKzZaTCNoQ6cHrRQJFiJXAvGIx23z/tj01T3oqj6I9wKN6M2
fUkaeOcvf9RMiXGK1a3+5xogGrSBlQJGVxhtcE5AuGsIdliQF4O+g8OWUsP2rR8c
5jYzJu1CDAm41cpMG7MGC9rYYJi790WUqKiz+9wOil7xv+9bEO28hACWyFdWGWiI
BdfrFVwMfKjmUniimN/QCmoG3hpirAlDnKMZN93r14P86DFR0Npne4L8wkOy5UKN
yZSEGdNvfQyl7cncLhmIw5mwMknizm+xzpn8JnBcTCWrTEdCA8xNFKDd8UVVx/uu
RSWoo1TuyZ2MjfxCHSTBycqmrPTiAJMF8qVjGKWDuoGN2zCzFE5jfxaoeDo3pYO7
kJOgoccdm2qsbUjdMSF5IyJJoij/88UOZn4nAHOrKyemnjVISMAZro7efxY6J0Cq
zBgCb1tc7ojEiH/+TrOgXwqmQdRGG+MloYYoW10+c53QMAcY4++DZnK79zS+0rNt
NK3CDEM85XGnYDMhvxvanMVENAd0R8rmMhcuUOdsKkNL3aQdN7jCFuja3sPhXrwx
TiPMWQItUN6LyG1x+s02wvZrBg5SbN4jtA7h3q6IPZiJgB29xR6KmEuwnQQw9flH
ff4V+IjbBPYYNw9wRXP2QT7D5Ttdc0hbYz1+tao/wteNpdwewRr8jlxBK7MTya+g
CDNuvMeWQxvW2A0tUitWJDeruWFKRftRR00DB/l5wXMlLkF3Hy9aBuOtH+c24sQw
YDGAQafWHBM3P9iNhCcu4Jd5GHoaZnT40UfTAknY8TLrkWeLUK1G/RSbZGuA59WN
ojeoHf2U5AwCHJaBq3K8Th0KAFnLU3tD4CaW2drOkEtrrvBgZLYm/38S6a5G98rP
8YbbIn4gJ7Z9EgpV69HpNaGPmuvpkEO+M+0/8Tr9DAbxPwr2H+//BenwWGOrPfce
GGoQnfde6iTVnHGXxUEgFjox8mLAwlQ7DA4/kWCRvRfENGlaw9lTDX3bQG6tEjKK
T2qkPaJgjqBK+Cvl45f0ImVTn0B+7f1+HuyymvTjAs7I8/HODkp8uq1S2jZ8ty+h
9Tn4wIVFlOmDoxEykOaszadU+FimECqtZFDOfUUwy2Vgpaw++7vsgi0D5GP1lQNV
c69UKKlttlCI/+BKIFc56ONeiG15/avPfOP0wLIaCdpZS/8z9ahXImQSEXCHJ2R4
NuUgGJE4R7e3nq8KcswbggoeiZ4jfkF0sp5HS36yfQ5G0aToConZcPK6qMZJhmrG
ZCvjYcqqSMfEK2u+usaooS81t7ot+IFv0509VWbOmJUWWqA4ISOxzkhEPUzTx593
5LQ32N5V1OT373Q5RGvFe9q50gr9zqyqrwgVZ4SMfU2ZSyVUi7m6unj9qqmbQyiw
XCm9VNoZEeY6n1xXs2koUfjh1ZabKOkfO8FF7wZoy4FgwUW/6R29ANQm8cHGkvzG
4ptjLwIU4jWNSd9M374y6bwS4gNh+Aduyb2AxNFTs+0ysMCVF9QhgW62YSbLj5fn
YbCBoJkOsxROWgEVOKbNrCh9S6JLlQpM9E8hOXPbpj2iadnyiuLomt1HHYOvooPP
biR0emU5qevvr76ykoVZTle2td0wSG3EEz97kehjW+fyNn2t19UiEMc3PUMKWUEL
f3s3M3JmqUmQafgAn3vBjQDnggZdD2PKAv+n0gz7L20lc36xdg4MKaX0baQ3asW0
CcAB2XBg9NsIvnI/9xx7eN4IUl81iypQt7AHpasCmoGePqtWGZFN6hR+eFNyuPfq
Yu7v8fefa6F+GoLFs0REDa+eDdOZjd5CIlELxZoJjnlu24Ws+5F0UzJjPzjZD/oE
9dgcvlwDEwW9BMRKygwJD4PITLrOxM4wqS3QLNf0PlQ8RlThH8zHSWFHQIByYxla
Hkc15Soz5nJh0dmMGo2bOaHZJSjcHkIPIPyRr4RFxqb+Z+TPsz/C0hEOA4UH3y6h
7BNP2O+jyNRNKHVeG01Vg5pQpCa3RkavL7PGzB1JG7tRqyBbUYKFrg7dMNn8JbNj
DTH/Je7Gz35Oy0v86XPCjqjSD6gFQhojarwXrsOJoH+8YVW7hvSaM2K1f0Li0v0f
KvI+9G4m/YtTq8F8FyuBC9+y4fVtIqNlkti0mqW8ibHx57qrZsj/ZEInPrrf98CH
RYeAOJiT8Fvy6LhwLHxiW+GwaAs6KuFrOD0i82xqWv6nc3iwr3JH61sEsvW932Uk
AUTkciUs86/FEXbb/WfDcmYRZ5I/Wb1l1GHr1m0fxQdcaYmM2Yy1iMTOGopwn2/S
CANWan5HTOl3FDccQ83L4aAtlo1Nw16zAcihuG+WFxe3AIJc4gr/MQ3k2XC6Vhas
tGMupQRh5ICIb1O0VKKxW9hLPMhjr9eihKGzDHLZQ4Pe1/RkjUBIrjCiF3r2zFNr
rhqnN9ZXfzOivI0S+NkK5BCq/V4PLQCo9wwnUGcuvPYDsBX6Tu9anEQyvPeCtR/1
4tK5p1XHZiBH+C+ckrdW8D3IlpvngkerMXsPXJ4x1zApglpLnWlOTPujC94Fnrn+
0slc+Q2rMV/uBuBt12hMvYoOUVurUS1el2eFcpJ7VF+/O5db9YDGgOxf3uS96SrG
xS6EVF+PxH0xjuKnHB0PVZT7IrF8jsRjkiIzQZyBcolsK4c+cY1ayrIhVlzb2Ecu
ZViPONpRLGeJeSFr9IIkSo7++CrFYoknPH+mvj6aI96J7Z3yRQjuEHOt59Y/q5fM
7Zjm0l98/gNMK6t0xrYQTZGmFkusb1mQgkiBmOZ0NoS82yTIF5SrPVY0PmhvFW+a
OxF9MfO5WMg1KloquZ2u+Zmt0Df4ZNAqAh4EDHaO9GUaSfLCeaU5jXLwMS5A0fq4
W08xaqiXXlqWnY6/i0yshUJE6gYogfH1LGxK+W4JoJZV/99sYY6BjaOfQtdEawOU
KEo/VOxXAd0W647jtmm/0cVa8T6SfWQp2y0zrYUF/sBIVXVzGtQcPA4WgC/sVeyo
2SqynGyFgSPRwGziEEOQjmb16HIw9dOFkuZEHJNZAXKCby0pwubcu5amF739G1a4
CWe9JFtZHNADZRmitx6gNXGkpWakkoMLyGchHhZDOSjzpcpbFVOVjIJg8fz34On/
ec1Ad+XK/PETQ/2nofVhZ8MVEHKL4NLARn2MLDnpvzN2s0WvEIWTZOyRXSXXxqF/
9z+Uc3deNjzucCL5GJZbd7p+YscsCnWYInDGpeivpz0DRt2+3KDB12DM9JdqX88A
FWCvbf2984I+hTDGvLHAOe5T3WMDMGwn7OtlPOZdyfxqih1GZ2ih/fOJXEqPSHr0
Q2muoOqxZf6f+7+ZYVb5g0epUTWSsl90REKIfsAy6gha6VVgYJKtI49SmQPV3u1T
b2D9Ji280JgBwjnYMmCboDY6tIRB666lVe0bSsHxyNMzg4xoSgQm/W4ys37c84GN
mYLGXlqmM6y6DEUfDtVIoBXUgFIXvXdspt8AjA4NpI1op7XpD3P4gsURGFlJGHAV
+2p4TNw6QRr91RiEjezdbkl0VC00v5J1IL8Op4vDQQd12d4BHsHo2Sm5VQmJDhY+
MjP3xvgsrECEDCuwGmUrxBXwAriOxaCXwZp7isHmA/E3u8mPiDIaWu/cXqZOIdEq
Iv/E5zegBmsx4DN/7b+vnCbjgi6Ahu4u2xRya7pVAqL06pa3CxyMI3g3KTTRd7us
imK2NGO/TkGEMBa5Wrt2gEp66c/OD5J48YwUEaMKExfUNAepxV01DSCwn1QwJyqz
6D06I/uphctpeVRSkSqB4wU3Ka5u9NGbcOscyFx5IX4E+TMhnv21boZ42+0S0IFe
CCxOOyw55SE1s4uuxAaF45cjx5hgw00z3OSPBl9BuEa6zLMVdlFPQvyla4yaKtZ4
Jf1QYYOd7chSHodB1q/9WXnCIgnsekYSO9EPMKFzcIv/yu5yi8SemzYB5pDaQ+2O
7V1h96LzWdM0uS/GveHc3cCcmZtcYSoY2t1H9truiaWGPwu5CtHqE2KhbptUWgwk
vOJvL1OT737zwVDIBa+csMLZrGSW+FIgDda24eQpXQ7F+mK0LxopOSS14F8VQyqY
e4qLtmykkqk/PPTkzr8LEMKi/op0CWDHPdUA7zWtCoQ1OQr4BCefbCVsYxWJJ2F+
zify2I2uHpLebGj8ENZ2xaocDIydKkT7gdxyl3grGXBDLghPhs8fE+34y20fHCed
rQ662AuL31w63I/AheD1f9hEqMklHWjF+R+0HcDSX+EXw3Cg1K2hs1a9mWWQ4gE7
iFbKZxJuq7ueMxFwKavNKXdw3G/f8CczevbZ9fOdZBbYEc0ncIh1PknfGMG/fa6i
BPjdPehXNehmUN02bUupRMDJzsHe78z4xaAtIke8b+Ylv4Yjkccy+BIYg6rbnuv1
KbfcrZXSN+U6aSjNQxNV3mVc4QB20KM0eqPRD1e38dX/LQjeq32ZJQjYuvBs/X6G
QYWUJvp6n0KftDl1TVpbckMVQfMrx9RoGaDALVi/aKgJnYWbUHgkkxzFivgi0GBN
Q32ASixuNZbzLy9WbgEC7AyN9ALw3ZU8ufPgaNthHgA/8Pc+sNNorKlUnFEfFsf6
f9mlYtKNzdA1+9L+/SvW1hPvKLf5R08/pAWpkouKEplC6X/MsNBBmgHeb0Q5yzqR
/zGHWYOSHjJAQDEsLbb9ysmqiDN6C1QFQIqJDbJDHqBqEdsIBpozuqLZYZxYsUsQ
r3MHEmuCtQmHr5MY1ndpAwholtqECnJLsOZgOeLhbji2/+l+G6OB6edM9btF4DHL
HEZKMGI5x5o2EZU2UMQ0VBvoTAs0aHVwVgx1Lf11lCYTlgtDivhWCLRiLy7Zznix
LA665MOZPP1aCvs8Xh4DulPdj695dh/K9YKjPCZJLF0J5sfcC/tAQAbJ6mGRv34Y
qLoQGVhQcvsS3gRP7jn9/TYsIUJILTgh8WmEaA/q/UV2IERyHedRMqH/Q3IqGbFf
eJMg7L2oRpsDN5W2OHWYKn5Ft7YW8zCKy71YoIneggroXUMQSfN4qDMv+VCe+V07
GtS6cuYen2N+/1JmLJR7N9lyEPgmB15Nm5QSyCC8PA0zI+ivEYlTNViY3wgpaADU
jSDxEVN7WO/dlCtc+mpPhG8DVAmjyiN+OiQ/hcL3JTOtr9BwWy3Vvi8H3xXJWpcf
nooL1YLDIXr1SWGfn5NxUNrY3WHhef1ppgsyYMNj5Ff/ClkHRwmTs5jg3Uz9chew
VLJQq8wXxONeH64xbWVmKQ80Pl29immpf6mWURHWmh42Lj9Ch1mScmp7n/i/W81A
EI+Iy4lO6hmgCnjiYBwVZ/Axq7sd/PeEN9w3dp7mW0krnWQA0P+Mmr3csMBpqqcJ
clGjewqOFMG8EsjZhqu/PN6iLzxVJw0+gNjkA8+n+tNSJpuN85MoObea1UyjR9sZ
bcgqzO4v6PNAeutWxZRhurmSfaAmEb+AxprCuLNp2rSWrLYrQLtG3piC5g0OZ2Lj
MM2zymZjkE1UaipbxmckfGBM6YtaF0EtNEVJu3NZVIBdUBTREcSmWyWOyxzi11+6
iIc32RKU82B0InkcAmVTCn0UTCWNcYCKD4fTkgCCjnyAiMM6ceDfMseFuSaX9z2i
JU/+6h3t+FZHhzKN7DSbORsf5m7DbVdUSTgAqFqol1CImzWADtV3ROsEzTzJ3xhz
FD7pwwEzrD8gUnv7sC7MQ+w1fJB6te/vAOWmZl0gV5yI3DuUkWlXu+WaBHnYoJLJ
v9zLSL9y0guN/Z+sVzoVMQ==
`protect END_PROTECTED
