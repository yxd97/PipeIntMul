`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1BEGvNDY5UTDx4sm398KtnR0nIyyKYSAfb01wVkS0MtEM8G6uOfV6nk5NifthPWg
gEz5auEsAqucdlExD18bWaGt9aaM6Wdyud0KSElNg+xRpvB+MOKfgCE7CVv+BsF9
DQa57po7ruzThvocC4/76EIDnPEeg3tyQ5b1oh80sLaEeMzbRMAbVtf4ktZ98PdX
lDXpH+DMB2XX6S4jGkGYbE6qa5TH499jUFnzEWXR+dTVHaDLHFOjlIz5DvhnT1tV
f5LnNhX1pZ5lPbxLEphII4TNKOG85EoSxnh4HeqJdk3UH69ugp0ScM6E6KNXJ9lU
D4+gVAuMBxHjYCqGkJCdfvmPA/0kncqS5aOttqmENwOYpwfR7aNXP4wdz4oedj9w
3VeWPyz1ZVu8bB+kUAgdK4gWtafc432erJq2u5mZmlFpigRNLO3Jzl63TTLOBlLB
7vDsKexbj36K8OZAeOrKqH8X3RnMbX8xg3NDmVJA1YesYvzi3SBxhAjnsEj5xOAh
b73fWM54T43HhO8cRLzkuEkse228HKQdEiTbcRdlUNPXx/sZv0ppvwnyGq24eWIw
jFfCuLJLemC1yxO+2fMHRagUMMd0FHbv0rrg43VjBhPU3nFNxCDmHy4xh+T1r2OY
P5zU82Us13e+/b2UJ/yWatkC1Y9dorLDMybqafntCTs4NojNhTh6Xj/s+hffYyh4
E85NeEqWUjFnVWZos/1pz5BJoldQETA2lpmb1hBovQ52BDWuOlgYXuhGb3S6BEzb
lW5LVUrZo5f92cZdT7vGKz65bWHjr6237snpHKoYCJBFRbPCYHhv1z6rWHGdjNG+
s0w6aVqjoAtrMaNlSmUxqGOj6Yqimp2UnTukd+xRPsZwTY4O7xkdfA265/rMPfOx
OuO0Pv4y3XkB4CPkQXIfrkyqPGLb1spJ0bNoO3Y5AoPux/pePo/IOwZh+Pm2ApXx
lyrURTLEwVGKevj/cQLnpeNpuV1Mrdko+6HF+7RtiT7gXticLQnyvkyzgVTKbL+C
Xd3R4rj8pdF40ekZpSQ+XciJcznoDtpyftrzNu6JWQoPGcZOa5CuJ/ceioHR0oc5
et4KYIlQx+o6AHBwxIzm8Q==
`protect END_PROTECTED
