`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uQtoZZPKOHL7BhUgF1CQDhXHfFWQ49tqQlEFpAvLuNX7joNSbprCUzX2HEyGuBX7
BozhQoGXbwf8LwVdi1oUdtw7JBcU0OFWFeIVD/Ru67QJlJi7w2eR4Uj7ICTOlc9h
ul4olJ3REe6+q6Uj8F7eJQzsRVk9oDi54gkcJmQxxsrjmXr9Fwy30rIQcIIkVf6s
tefIbV1+j92WNvVW0t3Yiq8TIun6xtUrxczkr/yZqmJPf4fbQtIZLCcGmE8J9u+s
e4m7jcaJbB/bsAqrqfxsJP9HfiXKnpQLPMQwcZGbFYjefoXNCedZef+sfBRSaE/v
6SIwjOvt791ef/lUCGpEWP9/5a5NnrBvx4s3k+shYSJIaDSQGzTx+7xiAr2hJlqw
6NduPNeO8x5iZpqV34K0KMmE05ob1TDBcgPU5ZCm74K80lKDuOoifkORtg/v17tJ
MEYPwOSrRuGrCOYYmqRT9KzVPjIWdcGsa39W8Yoc3sIMGMIQuN8O6JU+7e+GwsgD
37AAAaqyLXJh6YoaWFgpgbgZEtXVXKsO1k5NFSo0rnGtiEwcR8p7VioDwi54Q5UY
kPRNmyVbHc43CQg9+70/jmtwOroPqUPl7ckiJB9One0jVpAIkCIRCmfI/wsa8Bl/
x66xaEV46OGAfc1evVps3NBz0QBJGj+ln/+fC9COYN/OOq4PpZSWCueyzJOAlv8D
GFs0hQOEwXreFpggCBjup4aBpzTHj8lRY/ZyDt4IZs7isAU3ZJXfQv9d4pREv5x1
O3vMKpS+tE8M8hMwyFw6H7fxLvia61KqD51jjRGllRdw+aCe6K5v/7zK0xKv4Qlm
qA4f0XrIg73xHMbi5uEwFWQ6z8C5CTNYwJ/ptKTuGuNbILBMx1qEbYCUekpYYzXh
slMcOQpGOU1+vGF5mgiUyHlRktjvHSUOq/7ERw3w40p8J5OMv+s0qz5RZDoCDciI
TM3ZskS00esjeX3Gsl65+bwIntzi8q6pReYV/tFma90+HxX5HIEERYVm6xpxqA4t
4rPzbZmSB9NtumUFMVWRsIlhIH2WZz1jZH43cDiGMBDTFHN034pvCiemy0/kFkzo
vy+1gECBQqmeMo6YAg1gyPXoL03dEyrbpfv2H0VxXUexn1UhNDCT7YywsL1DFFb6
oO2v/BknfijfYufX1KGxTvcEjiToto+BRTJ+/QTTfoqrGUoBR+t7y3EDGaGzhJ6i
S0e2f0E87iNVGzYMFY2LZeao6Hi1M2MPmu5f+WOYD461naJatYomSIiot+I/wQw4
JYjHr2he8toYBNoj4rOWLv3vi41BLETn7LyV94XHb1DSuM+3VG6haqBKPnCDXZc7
mMkUbWEXJXU7otyNuXsJ2CgWO54lUuAC6yZxHk7g4PfDaAa7K3iWCzZLkCw9EBEE
i/gKLG6aG9j92VV0VV0FaCLALYZ0lDU+tJnViDN5gtz+HZe4NdOjjniqKVzyU34r
l8NGInMVs7vBvEEaMr2jslRN2YF9vZp+43/idvwHK6d0TIzNCG7iszk3OLTeK/8f
/HLRRzL8d/jGdyfL14NJ/kWfVR8RyuakqBGmh8cyefI73NgXupJsYZghMJlQJoEO
8+5m8j7nIe8xEogoO5beD4RkDBUYDQ/Cf8nkTU2uC49ngPerm93KAlV+r1TZuoEa
2Xp0oFUsP7H4Sz/LmcJEMwxmi0r4hOFUpvifBq7nQfBrAzJr99scoCz/AsdJsy0r
8bbeGtglDQCTqfJkHS5PtA94pE0vDTfUDUGQuW9XHcflTAFqhmJSWR8R/huP6szo
shNonQGFMSDR+eBY+9mNkNqx54wYEfyRj070MfPw+lS1cMdZlZzkLw+DuyjaZwms
SJO6MJAVwu4NMMaOA5EMGW38q8fmKIMr9A64CcSyYP6BtDhl17OqLSueGYxrzYN8
`protect END_PROTECTED
