`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PZ8G1LKBZ7Bm7O6Bw6kFv9QKUUDuquO6Xhl5tx1MpLUEfDTo+HDsjmlkGwZB7uXC
3b0PuYmR/odmFWP5vyrIdCqp09xRWX+qXr3Skjw4no04ec1n4ztB0uKEglPmHIj3
xjmTQRhpTE2f5kfnC7kWPUUBgRqfZqtsUMlKhk4dbdbNCvnrIbL1JiUTXAbPgWT1
8EW02yLgR/weUhwwvCVmsbQOuXSjMk5m4qbLmP/uJBxnNdoFyYcjLE+w9E3y9UFr
njuXS6iZlzO5990Sgf+9vpLn5OS/2KUWxWflEaree+QJASBsjEsCfCy5HrGw+vTM
jvuLOmp5N8C1mQWUB04jnw==
`protect END_PROTECTED
