`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GaE8vi/c/q6rxlw2Ahy/q+tRMKMncQGbY810DtyFYyDX0FNCpLMbsjGfXaZbLsl6
0UFg1Uen92ouE1Ihydf+z6t+H4bgMvLO6l+qX64lXrTADDdpIzoz7UYQF9lqAavP
XRY56wIstBm4rwNvNg8OXNmlooFyO1Y2Qn1nkrh7KINaCfV7TPZbq95+Mfk7ffMI
yk7kKv3RHrOU4nRLACPIFaVaduKDbsmLTuZiRtv8ovRmyk9k3d3ypVJOHA2Kw67B
p2UJ7r+tWWaYx50M7PsL1h9/S6ICHwSO+fSgpgOkj9yX7LMtJ+ighenysvs034qB
5mGhzegJw5ErRf7QQKcsNA==
`protect END_PROTECTED
