`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xqv6KiF7haKO2krX5sd9xSPSExwUEAmiHEPWnXoCReYm4QtEmjzRf5bkwwP3GTa/
J9502dlMdNn4+PK0EMFYDY0FgFZpZhDdXGY1oupnVJlbOEB7HNvMyvFwe66wvDn0
wEb6P+THg4oxn3/u40rv9L1+dSi5i3Z6DS2uRMyl0FtExTIA6Fh6A8peBkqW/Td+
GEubWnI9ORTPNSdGyYU+i+jJr1gL2cvkqoTm+4rmCP2uxi5tTXfyS0ZU91Cjout0
6k7K91+MVFgyvEd4Vq0FbIVUc1MaP6PVzdBOqetNhOaWzIE9o9+1H/bRGcRRRq/K
SEaMftwwaP554Q0FD2eOzL8/H1OS2GuwfOdacwM7aqcXj5FGRFSK5R8a2GP3wli/
`protect END_PROTECTED
