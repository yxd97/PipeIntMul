`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DP24aYAUZfv94auFmwix19ESKaxyPGXlpDXYvlhKj5TW8w6TmSBL4tNOueTMoC9R
BLxdOn3jOdWAcDI076bkvvcuVh67DXrVuN8fHa9UX2aQTxJJ1c1PudNmt1OxkoCt
CCbzTcfXpTsA0SUkRcuOWBMtRZ4Jm23v3ymk5b2msShVP+xIuzcN8wnZ4L/4Un7p
6EgWpbz4QXggphiXCOoNdYrg9l7ADm907+iJOVZPd967pTxX31wlaVNFvAMDVyUc
+0pW86jGsHRklrRocT7RAyPwVcIWxfguVdKddBSEsK8rAECTGi+R7kP7XHfAggdr
t/XCtg2zFhxPW+LPiNGDLbAnGGxDYcREGNwjsAgdCi8slk43orE1y5sC4vj0Xq+2
ASSuYopsPLR5pvQPidgMHFWkRczIYiJJDJhqced8eHjFLe4z2ildHBkuWGCyMM4g
Ubrmi0KaaxBebgnPXDtCJVAutOIFi9wzi9/VYQApNyE=
`protect END_PROTECTED
