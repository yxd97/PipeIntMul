`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9tx1tBpxoy4gftaKd/o7BVWg2fuxf5ihChOpV/+0t/yXTsL200PlZgviEJMcjNH
Hl1WzL8DO5acaoJ8QfOKv9AS9YSvtPNPQxPGFOO43kPi2Yfml+E4YqWVekqF7r6G
p/V6GyiOGTFlg0+9rXoN4bg6pzYZ4a/cXAcFas8EPOPigWvuc6yc8+yvt2yDFL20
y/F+H+UbEmS/dnwmcYI49nKEFxGCGzOkqIvTdBS+tHZ4pZr97YUmLI+GONbw2T7w
502Dx6D1U/BMlV6oTQWDw8YneaVsetdHvU191gcXfhMUv6DTc9nqji/Km2O4jU/R
xi9EMTcmMeTQE/aUDiBx0GyTXBFjp7G6isxWg8kgmUhnXzzU5fzkYfdNufeilhzz
9e5qM0nSZIQF7obrTGEWlmglvDsVLMCNhilUouNC/ITtfzMyaJVYMN7mBBQOl/D2
hiJeBrJ1ZpCyPvJtfGEWgdbUayG/7/yqObEGYFbqiBiQ3zzFzujbQy0s2L6iYN+/
vOY6L/NibS18i+ls4f5Pnsxyrnm8Z3V9X+pVSBkNkSH286c+e5xIFcCtdxJ33gtC
t05TlexuVgFQRdd629ekePL6YyNMuAi0optLVGQcJZjchobfB+GiBQvlvb/rOPV6
CRQdRqYfqyrO+V302zm5b8nO5TyV5Pzt3BI4yNyFbNGvTfRkbKRnAnmRz7WxJ7yx
gAnd4mXOU2r/kYaGUK3YJGYXKX404ZU2v6JtrpHZZT2SH1Wa+v81kQ2oP7YUqG3F
sGuNJuUo5dRfMewL7l+bvDy1WAbT0CBohMpRNdnHmvINSturk5ZMjIAkimocj68Y
DagoQXdpEIjGqsJE7x4Lb5BODC2LTptnMRiverv3uCEC8DKKpSwB0sVXgPQSM+Yt
0X/KF3FW9EibEom/qIEtZtFI40Nmw6rGGt1eQc98RjTV4fuq0pV6Hbccs4WeOYGh
mQfgCVqU3WialyjDlIPM1MKfIX+MSkJlHWS/8W3T0tKaF4ZOOsmMFyGuUQs9UR/y
TU/pOvwMtNp0ftDdxhWw+yXg/OVWjGkJUxezDH9Vm2+6949AjVrSs2gbEKlcB8EQ
fjnzGKyd4iQrYjlgektqhD0WAZFPn79Rry6/KGR3vyPIVjizz2ok6tLp/fuv7+ml
ZZ9SoQ2yvxxFrHiw5cTMV99No3GL5ZWlmsEAvh8e0Ah9rwQEQYSH2Y7Iu4o5A4Ak
psoPGAAPgY51X+xgxCPOOTpU98RvyI+L9XDRbuvvbnjxt9guBuqB6JPvfpmR8RlV
N2xbzdm/P4TFgZNrbtyukKq8zKE2Iyg23cLc4nuTEQJjzEUb9FJoBW9/JzqrCfQf
rKQavjLgiAYR+WHL1K1BLf3RRrh2S2y6AF+r35ViCmuPR6fnTGN+8MfETVLhgnC+
AYdMJKXWk7DU9/3Zgv8qmu3WUPTqN5PxsqZ4Hpe9mKFW9B1b5yh0U6ImwVlR7fxq
q6vw83nXkxKb4SkABfeHpbLX5xa/tdSIMlJ91FqNt+JjMpnZQObJx/aiOB4Rk+JS
WJuniH5W3r7X+7O6Ba16IYPfLCngV27SIam41Czj5vdj4a6iHXwcOHSBaqklBIyZ
jarVeJAuFc4H+cTj1wF01SNcE3/oTCiiYtpOpAMInRnB3c8mXBN42RN3rqzKTwdM
7wCYspf7qZ0oIRJDLusPZLxC7H72xuiiydfUX9v8r6vkmGNjYRyBEgQkLTAyw+aS
B1SVk9VX7QXu04Oo/WLJkqVEOn7zm1WsiVuGtqX4i2uG3/1bjrWyOJSN+LIHbqTV
NeE5ee2h7cbz1YFuirrp0r3ZPOu987nLb0VdKVpsoZkh1N+h7PHjROOrdeGdBQIs
wAJAP5dpwo60PZ8YxKANEh1lEvPYjmAIxWhJjJrtdUZE4TBlgBaWNnL9Z4G+9KGM
Zp/5x7t/7SGASPvV5bOugeI4ZmBVYmPWOqtTTIF78KfVVSbwGJ76m9yFXQ3geawn
eFGKolDVOsVE7rI2P1+iL7R6oNTp84MAAHA9LahC7HvLA6bUE+4GQNreaLX1s3DN
ZBWPTxnCIQXGs8lTS37NYCbu8Esrz8kJpuOAHTKinFhLO1eT2eUN0tHZPs2rocis
IREn3u/2BQhQBMRrxs+MJFgclB4wux8FIJMC2cx4OhqpTtTQCP3cQUly10c28ThL
`protect END_PROTECTED
