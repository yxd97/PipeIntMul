`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbXpA3B7NPylUfwdC6+MchXN0vdhp5IahhnIcCiSBJj5B6RlqhlAMLXS8s332G5G
hKbmHXbtbTDwiTagRSgs9GpNLYiPb8oGQ/0fAnU713VY21bmiJ1dMO10Z77RV1A9
NWq1GfpG+2gqJ0q78V/70XfMA+mPjbNubr6ZCkITtKHGasoyPlQw31L4Jncqp7ml
dgO3h2WjFkJ/gUJk4hvTXF/IgK1tSvspwr5TnbDkmIXssxplX+URI1pbePgdyG4t
NKNiDrEfzklfJIk2RDU7y0gl4KrL5InVjF/4RM1jwOTWNIDhmwL8emm/R0pNMqvg
Cz73i16hcFWs8nB+dDHKL97jgM1vj7HZ/6odUbSQApgzpqYl5tE5X0mV4Pl+Kz4E
hgk5YxpnFzWeVo0oZLArmhOH32m0nUf4NtKMCfvIBBYyFrXiFN/gsPcZXjGtRzpI
cTQ5m0gJDACoY62mZS+0dArOXJQ4pKoPDmBNy39xXgHyQVvqDo1fXOBO++7nbkG9
ZCZxh860W9TdO+av5W4FaAsFvlLCqbYtcVEgXJju1Eszhw7xxoD/Nfm/qxjtNt89
FR5H25KNmHRxT97TF/r1BmOe9o3lt4S0z5EQ5DmGjcmg8DkL9r2osDbwjdiA2JWJ
FkL+DQh7eXbgm+qCj36of85ffIcfDG1VoCZOk2FNyuLpjgYK3c3cOM7DpVAAErMb
MDIopxmtO1GUkHQEO1rXguaEkpLs9f/Y8LC4TFNTWT2VttOLn6PkBBirIaprwfgn
H+Oupwx3/kYqWfGOAmC8iGOz+uYQl9iAdt42dZJPFT/wx4QV0rtWZndczC02DTak
7r2LZUJf2q6XOLTCungwTRhp0ldhPamVrtqkpNhw0fc=
`protect END_PROTECTED
