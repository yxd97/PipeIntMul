`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P+dl6vQeBgpcKpeLnz66Ym/U8jGXP/tFXq1yGE0LDB7k0vYH4agjgY63m7RN1zB2
4k02GYEGYAGemv/JmhsHIWD1QF/PacI27Ehp1Cl/RPICFfjiHp6jGkRTTmqVDEUP
swEjBa/DPPk7yqBrDr2LbgmCcGE2aZ/yY4FPKpHPKbyNYiDps+Ou/tyCCloOs1M9
IDL8lSHLWm4xkxWTq/XQq3jpf12Sa813LjMFrI85f3INtbggCbfZqPIIwdXD2No4
E8MGe4py43MS7WpEE42+jd7OwAb9JTD7WFssxGCxp4Gsf283v+5H9jUFVIMoYUzy
VqpzkDDl9raa3nVRxJW8BhUFxv6mDHp0XWL5hhc31kJU+VxZAouIF6CdLc2HGjh4
KI/HHUcGeKk3zb0DyHx0f/Zvp02DXfPqLe+1dTP6p0viR9doIxElSUN4OgcXhz1p
dYHZJckHEfBv6+r0c+I4sskCk4m5VJO92wSlOaB3oYG2qcbAUE1e2FyJoN0RKKez
`protect END_PROTECTED
