`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aJr7uK7puu0YjPDASMqgFGuk8x+PqWbdjAFHoLDmAtIHava40L9ZBujc7G1Sa0LU
nQofhisLcVIY3H1tCgWf203bZYFd1JiQH9x+wnTFVjjAgJx4ma4B1gpzb9LvtWh2
zM0c7+dOFdtJKbX4DwvcsVlPuu08X+wRJeQVTNekXkgif1Pd3S/myDaqbFavTkq1
mAXc11v7IT8MbHXZaY+wk/jcgojpaPXBAbZR4KrRpkSh1XIm+zcuLpqe7WwI52FD
dKtNLQbuiJTHWBVee5FBWWJDIHSg0JonQAkLjKTJz0W1V9B359wrTnvc9EK7Ij0s
/kLTtBMg46q71lolDHrH/swIsieQW0BbdZu8TnOCtj3g1KLULoyTmXCTxU8kkhk/
7jSbjlLpfKIN0SzpWj9b7TkGBi4/jzebmmkNbiVVVrqC/mlQeRiX0mgM74aGnhzH
CY/ChrZIOOc3pzHBn2OhGGcM31tLFnqZrK7Vi87Kkes=
`protect END_PROTECTED
