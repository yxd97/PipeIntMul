`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VctgjdHpAiJ3RU2KfXv/Rko1/G3hhelZuRPGEupPxFx8cIvsY8UAxbV0lJ6t0fax
nm4kep8Ztx4972ldvZJJdfeY91YITAhxhrtdMT7HMxros1iZfG8UI95WXdGBGSgy
muc5J5u+iIsRmBW4oDYxvG56S3QW7D7OZQihImHmHtymLqb0nTY/a581wV/md5Qh
AZpgWpSyYxSDyD75Js5ZomflN208ILjGw3ZVj5RhgZ/JCKPGFX9vWFjagvNRKUgV
Z9L4S5yaDW7nds4EIDFeeL8wCxsC8WgYe5hdPZUKcOeO2Vqmh4/SBdGAbEyFs3gd
qIbVdKgX6lZwVriFQmBwB15qrQ1GygDjUfaNiODjgHsMjulQ37QTUpoXxYrydWaQ
3MxIYA91A+G4anPv0yZKauk02vzhTsu9c6UVgvzzXRwGWQxaWeBUtAmu3GsGquRm
HG4fiV/jJBjuSHl1MQx7NJcJ0NFoO3oBwVRBsD0JXO6MurPuTMV6w3rB3Lsi0Hcv
UWL2YVYsAFReWMI/f1lwFlEy2NqpdT41S4KB2ri2/C5AxzmT+XHmWe78FIFxSEW1
Ou8Gt6eDoTYOwyNcVBPs2oUXhKsTbyBXjM4BlJ8//XA4GvgPYqojenofPL5fyk21
TCkzZuk4j1lAQxBdJ+weeXQwtHszOaTENy+0trhULGa+nUcCCqjM8kMcF8f6PxLt
EbnUZokCBfWrJSerpTG3DA6nXj90jAUa3H8c4TPjHuxv5QeOqFj4vCM/fXffGJbY
1MzYekTKiGNHgPFm1R+IaSjd98+RDawycIN8VV7Bm+prNtK6n5RxCYm9wgDAiwfY
I0cjOhm8oRMI0t/LTySfkybr87Heos5ptwq0JcLaiyWwYA5WPpni9cl93CRJeoTm
pgH25vZETCkZ8zfsFLXy6/WOgVAOxqK4YUgVxoEWYz0wIl0MOUATQi7IX+KUpNXo
1xloWUW1dtBh2JD0zjnzWQ==
`protect END_PROTECTED
