`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PvfBFLAOohsURkIWv61dxz26Hw0IHkzIUIXqtn7anU2L6RpiJNW5SLZupJxsWpY
C6I8LHD1lKijsKZOMvOJGRPAaA5q+L7VzAU4xnSNU2kRMOBlwK6wP3ebydmS2ODd
iXEE62rzbKzDO612gx2JmYX1svmPpl88JNpK3w5UikKXxcPGZyCloVeIiUYI7nEp
C/17NYYZ0cJNgdsuyukwer2TZNM/ZAo2kVWVMCy5GzvDP95LZlrkRU/nbXzOwV0M
6G+ZL9jCGLxW0zWyiFgjUs7CPQ1WxvfuWz9Omux1LOEYFnD6HdUYD5Dzji5f8Wma
6IbsAwpwsnhUdXyOFVHh/6ehF0c2PAa2/Utb6RcypJnJ+mP9GXzBoEEpXoPh4irg
DwSEAhrWKpojqtmNjC7NdA==
`protect END_PROTECTED
