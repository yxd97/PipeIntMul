`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lGWYD9d9mVgosyo2AtRYrgde3Ga/3XhKBs0iJKPsQVRQsqj+ZTsUKL1kc1WjVPl3
qiaIfnf9hQpebF+PXR5V2hMF86STFkzRIPqDsfmva2KdcZFTMSJhIIEaTzNwYx9H
/JR8YDayt6vLkFQSAK5fes/PHUHTXnODlz2TVIQ0v9pNC0v7+gyFJB40T+V8qpjN
JzVW6ktJg9XTTIgDsXV9MAvisnKja4asPHwl4pf1tRsfJlGrM9+VHueKZpyKHh79
AS0ZFCQ3xj073Zj5lqcXI3iD+VCkgJ2tTRxrAURAEz6xB0XSdGnsY7w7/75nS2/L
i2MMV3S+piuikasLOTVuwUl8syzkH5+TDZFY3ngt7VvAkHQIMKvA5ok8B4R3RcQS
9kkWgBnLfhphtpmTtt9t79cdaraLIIHmZ8sfj8/AHNjtKLU1OEuxIcic/A5E/ipW
216PUAluVwha3PYsreWTj+QLSrgIxeEjbisHmMVwTUc=
`protect END_PROTECTED
