`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1m87PYj9d+kHoMlm5pzZYF+WdeWXO5JXvDK9pkz+KpJpjB6l+xpKZtNm1qRN1D2e
aimQhTxEHpWsxhLdBYtglFCvG8AQR5YyM/ELita/tZ69v1MthuenJhxCfsc8UjiQ
3W1IktmuYRIn8Q50jS3wBz6h/Sytu9EJZ7GohQkT2q7pJsQvDjarEl3AGWYZvqxu
n8mWb9kSHvoIf8rI/n7s9mwiKUYef+8RjbrFgzFMPdTfTY856IZeTOMm4J6IfJYq
1Qy8834rWsk+80PGsdAE8xwu2m6i6Jgq8MEHG6PYpTqtKAMtB9zxivOU62FTm0Lk
CTsDMFZD9yEJVhl5HkBOLMTC0GkbyTqGspf7Lh15/i0bsxVCwNT2NGKTZ+4K2+Yh
`protect END_PROTECTED
