`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o5wbsXXlLwm6+pjpBpYfgm+VoHJFKk9EU58JEf2ScqW/GYIYw+vdWVjMKhCPkHL4
1rYGunkRkFKQBfF+yuIvMK2vxZ0nHbG6wBnkhl84nTTM8n6dPl0IkUOLBwfdCecx
WeUx4HwWCFxHCxTZPjJgVnjcNpyy+4CA6RokpQtuYxigr8yfR+3Hl51CuQkb2OAW
CdW4ttZ7mq6C8KAqg6H+Act/S+LS7voTcCYDjDhYZCkjD4cN5pQg8XgP3tQF5ihk
b60lVGbcBMH55kS83wJZe6DOQXCzb4d66neNf2ecK5zs3JA0hF9q0vmdXWZeVqUA
8UnHQICl7RBLO5/kfdRehPj0b19piVu1nkUC9ymeJZXkZzbHicIoQVNOyevwU9+K
4yj87kyIvy/v3j1bBjkm9kW1vU75JL1t7CfS7KjLa9U=
`protect END_PROTECTED
