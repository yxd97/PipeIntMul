`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgnAdgAdFzAdwNbUK5gNe0Iqgq/B1T+TKfbRhWNUhqdM1TyJAew0jy5HQNoPVHJa
y+7KG52HGuDOA4Br4XpPspq2yLLzciDEwqoYhwSG/U+lqukd8UN2sh7rtbQT7Se1
8j6vhKvmBwvQnNdZTUcECU5ddEdco80QQVfGKf1XoddKNdi1Vz2sLAe5V7A4DLsA
F8Kyu1N4LgbduzTeOqa/RlzFvFlhiwzlhgcqVy3AgKC1/l7Nu5Ik4jFlY7pohOcZ
eRmR04FLheW65NZmMO1K1PoY4ebIceB5qa/RXEZ4t3WhWlG8ssUWQL4f6W/7yLsN
wVfCqzWJ5yQV1Bqzvqfa4tWQs9+heq2zAPi/onPAJ9Pc8VntZ3f4v0SBrkD5bC3F
8IxvWCKUEt7zz9xSD7MrZRSMyneANiarLkophO3tOwKPUPhWxnZJeElOrR+ivEpC
j+oWyI4DTZNIr2ThnBt7ZxRIN4HQpXEpOfFQB1AeJeKWGQpeVhPkV9DbT39VKuMF
BysunfAB+iIfxlI8Od+vnYtHmfKcqfd0tDt61UGV1bFUQigK/QT+iXSdzuVVcnwe
g+mBeJBIhPDd/Cc9aP4xZmkKuVe7G6E4uc5FzheZ86xuywMVKUfka18N+aqCEZST
V/+r77ZHKMXnQX25q3yDjbyjJbNw2o0AFLmMJAoK1DsLepkh5Ub1/W3w1Bjpt6e/
sDXrJ9Ns+vTW/caK9AthbG8akiJVhk2PRxzyR6aRC+nxF/XJiZYmv/S6vndE/RI0
3h83UTGSSNr+DZnvnjVWC7WxJzC7EW8qghAC3X2z6C7CQj/niZQL+OplLa21e4Ft
0Aj5MitU+ZhQ8VaXv9DNRBizw8SPGnhBD1QYIYGm5L5ZO9aG+BHn+L6cJ4oZpLsB
oMQQyRbITbePsDIO7bfmKHL5nJE3FSmsHw4o9rklJIdNoT8/yV9UIXcjjIrSbB0s
9eh8na7aspryZJ7DuYcYJE78p2ASlSz+0ATmkwF9GBWWOoMMMKEISvjOr8m3IlTq
O7WartUkbH9Wh6A4XfeJBngvKy0l7oreS+Yz5QqW9CTNvD3Apsc4TnpEwatOnXna
`protect END_PROTECTED
