`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RKjxH34jWCWvU0GmNOgkdGmjaq7YtYuCNQI6I1wTk8e/Q90MpykkqE25ChsWpnWN
sCqwKsDI3mLn8cf75XLIVXyN+5lx01/HJc1sk4/vOJXjFB1xZmgMN8ekfNePmfzX
cVUmppxUtB2YTopWZmlOVrnlc/dOi0bi4jvampM3yI/KpAalNBar9m5XlWHdiQs+
qKmNLvB3Rd+QgmMKvVrc0+7SzOBV+TWNDSCCqTk8s/BxDlALwM1xYHrgG0VhfgTw
wCJBldB+654cL163OTKhM4XOhjtwdgRHiDMkJZmdzR4vQ1qncB9XSB73fDzGp3v/
5ZxozNHmpqCa45uMboTLuAVunYoj/NsO5m/7dph025zz+7pWlegbAlk/9NrgHCqq
QinZLpHzVZce7iK4PHJTzeqH98xNcQlK3ziUsoI4IQ26uQNO/xveexm4v64hUEaM
JBjSb9aK9vKzUzZPo8JwA5TDAzap0IsdpsMEcLz+QlzT7hv2vSUDJ8vxZGp3MonJ
+KCcXDdVvJ+pJaj8yG7i56wFDEXWv7QoC+uIm55pa2qfB35ynhHPVAfzHSEeT5M6
A9XLAYPPu4w4WJBH4/O8sFDfEsZFAMoEhfJwax+CSX1GpBW+yFQxCiEDCWb7XoOL
5SF6bXCP+Nd55CnBxUZqGOZaxoz5Lkxu+6GH0nMpXVALSEcNRkcKCVPpeYFx0tjq
KefBxAzv0dPANb33a/FtSVV3gUM7rLCK4IT2rCBzpOWMLqw0EHsH40U4YVOr/VSZ
iwkRA5NctlCiJpiX+RbFRJevQygKdNTV0ZKSkreNUrWOyy2izCbJgMiCjAFIf8vi
MccmyFIIz+COExJY9sVXSToVDxpmQSmKPu3Q7pc4h/ED/6BCADX+MJqLwttWRgWE
PjCDNIVxBhEXQDFXKdarapVJ2UzjUU0Y3nPxOWKDNHApZOmF8o+78/a8Mma/E2KO
51+h3kQCTLu9nD8Nfd6qHaW2uxZs7sWEfRr+xPn8QA7oLJCpJx8R1Ffy4uk/W/jN
ijGIz8nUaoJ1zM21NIdj/yJULBDc1p4f7aHhX3YWggnBOlHh7qt//nDVlfU1bdAr
bopVJ1Is3MsHRURAMXS/xKwJ+hiAIyZ9K9XAMzZQmq0wxZsPjUz6jYa4FFFzsyhp
blh3r30suFOqNgpNqlN8pikQtuGUEJwXur8ek1GkCSemP+B8RCnBkFrz1Hhe5ccv
cxelS3X1w6wv6ZUsB1E+y6QPpKttc6yM+girYMD7jEADAWEfvETylaVBSS/bdOsI
XWC7ML4K1mA3v2kX5Hxq9nSbSzED4HEnzTiegBbR1ZLXOKZo3QQzsKtdvAoeANQ6
mjtYJNbAI3+N5wDfCwSNRk5JihFTd40XaWYIc5kMep2y9zBi8rxpoN423JTH1eGI
rTBkhbu+ryGQN257gTjK7ZdO0khM7IYPgPiPBkI7qThy5WFemTRqbnSsI1DDd1Hd
qiFZXsYD9OQdMgNV2ExYxN8nu/UzMBFfkXvQukPwpPINL+E9g8eZu0YEJ9pxB23v
FsRoudyVPc+adhiRHHG2kkyDNFe3BZowx/3yjOMCUtFEn426O/CHkaS5V/IW8iZ+
W35QjAyuDnwowimiPngbBSM5Ri6Bs3/kynCoFLPIeDbq8j8vJL+2p4ccdOPxgXQP
xOYYIIE828YzSJM+9RWYjt4S1y3f7Ex3eX/GkAiUba3RxY1FAFOqW2RaY1CpXLRm
XieTwK/cYXkXiMTbnMqL19o+i9qUJ4MXtUzrkIp6bGBqIr4gDVFf9wFcxfoP1SqQ
DawwnLtW5Zvzu6F3g96W8op0w4dNZZVZK+icvhiNNLo4JQl78KZ6GnutYzkjajLO
8LCT1W1w139lWSCGqzuJTpq46JXXAX57XVGxTNCcm4JDyafRvB3yHzSpyMjw2TQF
boGTWJsmxm0wR8f457Dru9dnIFgadJMr5tcvv/MXTrrY2iv+tW3ufusEuUOA7d9b
H3sRUxkTONKXuSPnVjLua55kgTrVb9JJItSS1LwZTibeyksSom9S1PAQ1Co87T9M
gRCLgf8umCn5r29aZdsdWZzAYDbrl1Bv+X8wvu+qlT9CrqvEQ0fEKWPonk+zTnfJ
YlGHFHXC8bk//ZZcRQa0tT5i5RmV9KE7oorgLisWhTdsnGBYjiH9LRsIBKXrdvCp
3AzzK9DtXpp+g2haQdrnozOWzgToaLrNWPdz2tvv9PkB7MmetKABa47BDYI9Y9Gf
BgMqbrSQ8zNINFcXcatG+tvP5l9E8ZSwCCHshUoWi0nN3RcTzs9qdczHJyEzozUh
0om+lrITOS/Cgultimw0Ii+nDDmT5sTasKC4zycaxqOm3BwOeGuSGPt4ZEhXu1kM
JGPWQ2XFdNE/yN4oQ2ljY9dUQO/T9MPE1Os5P59VjeH+9yz0pFXog2unqlj8Z42r
qbexeZsY0RoA6OFfS7jCcoMKQ7yYjWp8k/CI1VVp++6xoFxIs836d9ejxoQAh3Oq
lgEzp0hBjbPgdU9j9ChkaRJCLDtz7tQ0ppDH+yRlzCMO2vHMMaJXNHuz7N4e9lDo
4xEhuGDwGDJY1IohxulFSaIYib8QaSdfEhQ2dODEepq9aNRO9RbeitIHA5MXEg4r
qYT/p5dTxFQFJH3K873uZCgXhTsiPzwYQ9UBSGlcNHKm8ojKsISiXNDnkq2ob4FK
7iEtqpj7rRa7z4aBVz0YvU9Gcn9ARBL5LI6D7mGd73yGUJsFHC1Hzx1Ktv7dQ/iF
S/hGkXnsLxHrHP9hJGEhGnxR7h6TGem5xDVCvEVjcgg/kzVRjoP4UeyUceTVBDyi
I/Xy0vPKR0ZU9kQUYCfSXhg/E0ORDdA4VfknC53v0KVnqJtj9b1u66W5MqzQJMpv
wwnZr3maTy0sGU7Zy8ERtqNjLStZkExl7DSorehR+FYeGnamOPK9cAgBRwfnDqyK
kkQcPu4DreT+Pr1AzxTOBkKxuRJo/CIaxTXk1JMrOoo6ezo7hC4Wbyqu4KFpsWb3
ncZCA4fOT7Z6SwXq6A1LFA7P+3qnCDZJfslTH6Hh0+z4+Z5LFLDsI5SfMfEzYEtu
DF55sKNNWojGtPCNZttWjoH5nbL8fytV2iBmcgfuvva+GYI+wm7kHY8xKWpAg0rX
JUUXtiX7/+ShhuehrpoeGUofv7PKUIHaYYCVVYP3Iy8O9O6oPysS4B79GPgdC1Jf
KAuvS7TH8mkPLkkhGc5nuuaDq11OraSNHRakqFHhWPxLM1IHrRku04YxHAWwd+1i
xw0iq2rGVXVkvEaV9jH4WZnCHW1UA4O+A4kT4+7V54jl5AveQDUY7WDhFOopMhdH
m9x0AklgF6f78eVGG9FJ2oJVq2T64cUswTZRqQ/CX++S1NCBD16qP1/JgV16/PQ+
jP5iJsfZaiCK8fFGrnMLxWN1i0k2fPNglxm18SQYzDrHq0MFnrPJCCvlGJoQoYD3
XDIslsYwleG64ne+8bRwgK28TdQmmSEnm4mS3+ql5N5FaqpAxFu/QUF5UuhkFu8y
AqZxHp+5MI+aLTci30GCGxnnMwVPnJ03BOYdqkGCNaw2oKKLSfA1a7yrZqf3Yv8u
FUez6bqnEqnHjcZzNPSJPT5KocBoWukHbopsozg+l/J0zJavuFstb4xQOVobIa6h
XRn/hwXJVe9NUiAcIioINGPBY2uCS7nlqZqZ9Ps/x/bTONqM0oE7k60R9hbR2W/D
1fAErDdilsIyAbOEgS/rGkOKSSAtlvqnK3TU0BPNkciD/qcHZEAU8ERPsRvirh26
5HwjnkPaM9w9AknBQ83DI4W7bqUl6yQqUp0PnaNChqEYaJ+gsExyD1ldH98f5CWX
yQhJ1P1OmtlAF/cB7sEOo26JgKTflV7KQ/a6bTQRm5eGCx2F0OrVWDEIbd/sK2hE
7qHcSs7w8Syt9nNtVRARzJuItGMblizJXyhU9NInhNjd3NNkbrxdAs1QXWZWrHlQ
Qm6z2GYt6ay39X9lBhTCTLTrj7HSO7BpwbYK4y2lSf4VTFl2jHL0PS2TeNq4YmRE
y4JE+3aCWWjBrGXCiZCN/S3FBvMHS5PjckvO17qBmfcC+bTxPgp4l+4tAmKFyFK7
peoEJ+npez0jfbJK3mPaCLLiQA3xapDdOfjj9dy+QdII/UuuiprMm2zVQpCOMdYF
MG1mHEmQHf9dMmb3wjNa+hjS3FMLgOzmD18esKYafG+hS6aHrZYteFSvio5P0Ys1
o2hRmLVWU8e8Oe9BQ+RlWma1g8rOhWnzM7lIsgGjBe/rRBzbpBSbcP8kQdZ5bWDp
sXtb+yAdfaXqdjs2IniVEMktl64r9vfP0AEgoDr7Jr0aouJyVMdC7KuebkFzHUYH
wSYqi0YqIKombBe1beR1rSKrmjJ4KWjM8UV0sp8z/Esy7skaFA/0jZ12qkriUCgr
o1Db2y12+mXR41ykgD0QjCXzshJecFZ18hwnukthl2sO9GxQ8KznHQ2qFvADasW/
GV2JEcDpylLizWesNP932pVQauzKyiiF6TK+aI6o5/3p+3mJtXlhihGP2L9TKVaV
+azFaEnETqwGfV2+r65N0kIL9lwIpgJVN5FJHk3qUXjXiQXEH9alCje5sEY3hpBA
Q42pDMU3U4We08ZBpCZngUZwAVH+t4y3uMIZLqJlN6FrIFuMxsK40jUhm4FFgde/
5T/170IFo/wojequon2eX7sZ4jmiJLUIDLtwXBTgtRMg+JaS3J4ysrgZIfxbzWOV
4+B0Rk55892e+a5d054CIS+LH1ajwzcoVjXRW0rH5CdEaLhlP6bx78MGm/Dx83xR
UBWJ+/RDOgYKDx5CjP632WrnIVi0jHnoAt2JMfvnooXDvbioIlWB0UdMUEH1qzsX
+ZyJbckFmjQFykqIOirFSHMnV7rxJw9K9EVKsHe060bQAMPwiuEWWatcB/CBJohG
DyJCOzJjkgGG5lkJNxNbtP8DowhT/TKeFooXn95eqIABbhXfN4sSo65JvVBcYubf
qZ8LVgeD8HVGnH/9k+/wekEj6vAw1qkZE9cLYijbiqsDTer6CilBjyhrO40JWiCy
a0UuxXfr4Ijo4E4fCVAMOZBxtg997GqlZy4j8jD9fMcRHZAdvsZoVa0QO+2CulD3
LybtPUPdx07VPKMThZ8bk3fqr5rvp+qfznoSp/eq9K4v2ePrWnV6gj+s3fbf+AJP
Z+B7dOSXQHOb8izpm8ChwgIiO8VI2FwQbbwLi0uvJJlYrosQffoQJuckhtIJhZKs
f/nlINQ4G8DX3jNlfSeDZFIIEPF7SJLRpoYebLhWM57NzQVWWE036KfUvVF8pCXs
OuhN/te0eBtkMORGxpQ4DX+lfuLOGTlnrvGuOUcKU0E/1ZSBF2pG36OI81LW71Ib
tyOrvaayfIqL3dCVF7PmSWiS39tHxrBLlOQeuhCqcSKixe8ZvfuNFltK4Sac1IN4
bO1V6IoFzcTTBhY2Vp1h6/FM+Mb1nprWRPC87Zm0gEvvK92RB12JlKu9W/zYR4yG
zlw8RXGX/3g5bK4VnV7fJIBqhJNaJjIDgPeUq9yW4GA41wNbxkscsi46UV1otjYT
DgB4Hhpi6NtP/KEU17LCEon965jl/5ax1OnVdDtrTZXci7xwY0qNfJ7G6lXz7b17
0HDyCBKUS7suKxEYZl+NIT4fKgGaC27isecBF2mBcPjeetWEn3J/dPHUqwI37IGR
Wpk9UQd9oDxMqWR7qjjcaDXTEhUYqXX8t/VErzrupwQ+ym9wLHgz2VSg5W/SbSop
quZ6Hh6OcABpNT5KPmILDGpxrqXqeJ01xxYAATweHLrZMzNmPPN73ZLlPVjCWskP
hG5pWq3jz13S5j/l671B/WNMGfZ26Pp3vg798GURc8KMOd7doa3Ml0ejovc9ShsG
CBFJFX071NCMoKl5DMIhAzSPe+6NY9eU0Ayq5RlwMsbaF4cso6bO4w+sWFeshyDF
HmYWW/LoboNoBhFCUtnlRo7jGZA257sUq1SNfPRyrEaDBEYgVyx5r38p0iQt1Yfg
Hby5dWOJykQwQnTt6+8GY0dwU+05U/8Vt7cJgVEmb0NeK7Zn+M6v4nC+GBUX0GVH
NDLWuIVTND7dL4m/hboGHBZP1bE0hkrxj1HF4S2YBF6GxzuzWiHW/SyrEi4sG80o
iGCft+a011QEVgDN1cfrtD2t3bv8Wmir7dGExhcCVQLaNbtlHd+7EODin1/hitCT
y2kFJ8o7nh/FS7tj/HNLovORkbbcSR0ORBVGTFl7HUgj/lvVoRBmqGzQ3NmTSfQc
D8f8QpGTSsEaTO1pV4Vbzfxw7snzA3aVrg7jqogaCEJQd9AQ1xlcPZF8IzwQ6JR0
FsqD5YEjcfPI1N/5g++gmSSKTdOcgHz6glCmjpg9mlZNGXJUSkcQ/8g79uePjNmn
xic/n7rCUo6zMWVWUvipDVlhZLE2Y1+SlelnJHZz7vziYo+hvqNE8vq6Sho0/eOX
WDlsbskEZTFzh3tMCGw09w8ZSaausVAycX1caWkX/jcKO3kp56Zz2iL16UUVtRgI
jjb4wkjsxDQ+NCrTWmycxvicR6bMh/4OJZPdCryl2TMB8jHm7nP8Woj6NzzhoiTU
5Jl/lcGeOa2uFYhjzaBtEcBGZQFDDkcKqUKL5L0EI+u2AfIl3T/6htWxoxgJFG9p
IO2V4sha9Nct11Wf5l7h7DwiI4pVtp1hBQNX/JaP80gzrEH1SUufJB0UILoLZs2i
1OiP3KvNkCLvsn65Pe9I24+wQrRXRfzHE1wb2cydPuskMK0Y4gRXYUGuVn1vRWe2
TZ+ZIJF8b+4SX6YHxWBQKugvjAIeQLp3J1nhMb1JOjGaYpzXEYlNREKFr/U9Tb+p
WkQxdazyNcmDgUMz13DMV7siEGBj1JqsOd87EFsGb0gsoaSe4xo+rFdw5/A1AdVG
p4Qa6WCX9kyTfiGdihFhbOhMcJ95qRX9dBLEkMHEyJVvnRR4leumpl55hMkqoRPp
QBPsRWCPOdG2+s9g/493ENQ553/qyp9B1kh2b9lYoCjcfDAW7l21XqaNMjIFKaOE
T8o33Xs5xIczo6CTfNLjb+zml2kPO84klbb/Y9DOX/xPejosL9ZPMqTVZz1y02Gy
PV9SrkfvuVt0cLX8RczHSgufIwx2Gn/JD2H0H2gO6p6tgiOBDjINK+1e2Jt/X5xi
tuwqsrPwgWVV2adVy/hc8+tcRaCEcbmIlkpL4imA0+B4QtbqsacAHnWPt1ztAp2i
/L2rmMTd1Hn5nuHkFzr7zw49M+SvRjSpW6uXaLAW5s1e5fNNl5TV9G6jNNj6B44z
5Q8X405rRxmxXvdwD01HEXea1P9iyKEE4AJmKJU7nvtNWpqtjNGmTXbzMCsgXHpO
69FHyumDZFy2FfdCyM7f3fgXIiGF20XsLb1xI5ittjWJW+Zh2786kkzopGtFb3QP
rPmvwYIJXkGMh62h1pnmXppIXjZ8RLGsbgDveHG5hbW2M7835d2go1Vm0kgRRUhD
FUO78qPYpuoaHiWdbvHw3zN7XTbRK2M7mIN9fQohcb/XPyDMYECWQofWtQd7E54/
dSgG1jTECQk33gUlYGxQr7LUOS5vOuHbG1vxDnxErcRtjpNrnfnePamWuFGaK9mU
sQHQZzrHZt1CVK7AdAHlbHKS45cSMxHUOLB4rWAE6+vOFuGGhwPc9hGSDd4Ik1ks
Nnzr5rcC6eBVWjC26hyZZVo3338rP/RHvlHJ/taneS5M7E3ham9VDG5T9uojkbe3
KXZXVIvdrpTFu5Ou1ZyfuTVAEUjMJV4A4PpFmy9y022bd0+p5bGTtXsfCtTUUSft
DqFfyvdsbl5yhGQj8V904Q==
`protect END_PROTECTED
