`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VY7vHHP+115t+ud1DSmJGkG6Gy1uj3HJZzdI1O7WptqoIhho8yWD+SWzcjzgTmT
LmSsJJCxFgfUp2pSrC04GYkzEtvjOlBIwYPZaYkBggX7DWu8TrQCl/7/O2HyvXj9
KgC4r8kuwj39Knt6TPhvrE/v2++sgYImaJp1QGds55HdZSS/mJCZvU9TNCxR1JRh
FDbHdDEFOT9W7HKLB5VwPTsQnCI4jgDiF210l+1K/FbQR1tZ5FRWTLeQr7wOBgaD
Eldt7Rmiw3YmK04010SDEVaHAJkIXmybGDkjqDaAgaixs4k2WZuIJaP1lmhYCIlY
KTeUu8M9z0xvtRDs7ZVKDgxyL2NwY5ky70C4k0/1bwvUr65ASRfbahZWBKUUse+c
+bOjXj17T2Rpq6s9dUYFxmPYgvejWVsVho04Aq3j+8u4Lr9+EDLwFD9JzV0srPAM
CErVDUS14o2Sm20OEfiyWl88fDVNaWCONtQOOqXpm2oEqJX4K4Bcl4doEpIv1G96
ZHyO7dRLzxHkXFGgORPlnKpsYmEdDG5YmZYJtXZFkXThkLECjmV+ZS5QfNwifGyq
WowNaaRYsyXjC2qq+zc5NJ3FpuvCQbzJEvAi0VEBOApuHG8OoHr0vVs4fGMoS3uu
CL2YLI31QsA4i0vrZCjfe8VlNqfYbed+ltEYGz1rjpn9iPsIIyA8WLxSxkbmYm0Z
FZSmYXqUCaWjxlOWjzV/80uDNFE8OU/GpOkz7HOjR5hPY5OJ1J0boXM5CmxenIdQ
fdxbuQvtmfeiIrIaHRnxFsMzN01rkKI/uIwxaYbEd3BmvmtNss7KBYjaz03laOC7
qOVb8N93ly/C6GKwBLrOeLBq02I31yiQx6xGnmIYrbp+39KLfzEqiBNqUvxjwwfV
xZ632gMPnrZS6fK/3Ntc1WBCuJUvLXnm3ezj3tqKtK5c8vBzBwNI7gSQGm0R8zwY
Qi2i//8wUfo6Ez87ejzBhhEp//Nfng5Up0UGfu/sFMl8j8pK5DCJy209+jR6prtQ
DsstPYVEa1cO6W5zj0f7fhjn/qzsN3DBe7UEQUvgnyA+XxbAOZoeObVgE4Zbhekd
AtKws0b942rE+It3GXMltlMlvmHXd7xrBZJbDy2uuzOt4XxH9FHK2Y/myofiNje2
kL4/SIoJHujQUiFPGuOGft8lRCBvrzisUa5jnE51RIEDnqvTUlFHxFcNBsjwcWgw
zfLVRAmTyEK/HSKZfobFqtbvPhDFlj9F0GwWkwyi+Zn7u2D1eOZlNL/Bjpxa4EpF
IVdZpgdlL3om1MRLU1l/Nr/vcmKk0A1pUjc3Ecfsc+E95xmJ78t7fRnvV8SkT1Fi
zGL5SPnbCX+1FIKwi0AZTFxIQmyFnJt2/vFq2q4rklpOtjks7+szFKiNShTmkB3p
FdkhKqIRn0QZBiecxQV9Ivinay+lcsWSHAnAh6FRMpVZDQuBYW9rtijMNJSKu3al
bHiXLSGxZ/HMGvzmv2dQ8JTjLnji4AK4ZCImjSriQI+pp7aciSzBAtZ/0ur2W7wO
+HreA/EGcHRPuRERpANl0VzhlcpmliMkV5TAbfTzNDqsd0/gPUDG2w6qzITI7r5M
yBJn0Yf431mF3EgndEX+KqBFI8gJK2VaF/GFEDCr5QLjqLyg8b1f5om6Pnxbi7Fx
nbj2eY0OMQBuN/bS41Zx/+8R1JKRaskvlQ6riyT7omzzx3q0SIJaOeqbvUwwpd0S
FTAx7wPouAdxwNmbOy8AnVkdfsSG2v6t/TM8O6RJqGU1loecinZcxYd4jzyeEggF
rXlRw/FFokHp7kO3aZpEoJoIom7HBSuY0TjQXDXr4xC9nLBB9RJuYxn+RVklzMfq
ignItXftSkt8mUM3DZ1bB0UGBQ5ysU5105Fka3SDul9A+JVp/5mkfI+B1keO0aKR
mRUNA3guunU+ZqZialX9VbBnbkVtLBw3w3unLh9BWNLrRIYaBnlnI8M3wK16LhqM
ea7WDzVj0k1LF2HHtw9MVULaq+KFcwHJqif0+fRhpUzweScQ3ByYF0JjaqC8mZMX
P11D6mLgd15Bst2Gd/Uc3Y/N/sBfEUB0HTk8tiDKTbFowSy7wTdn//HTk/IHXs6s
lIbAJeRZVSCT/vDT7ow+4Wh4MKlyM6xHr+cFcTAqfHVye/NaXK5aPOYxJpocFvOP
PmRkCdwqesQOw6pC8RuRhZDbo/A/x/XnK5Dmg56i+vOiV4GUngPZqyOzu23EUboo
l1lU1QZOBIlKvBicr0UZRZayaTmFSi1sQVSwzUisi/F/LDUSPOwIsqUGU0Xl3gnr
Et1Wmbzl1XGca9gsV7zSUNAjOjiqzIjiGnG8nOW22IOMCIg4ol58T1nD4O1ClBem
`protect END_PROTECTED
