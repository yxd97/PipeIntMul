`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Eb9bk8w9JSSJV5NQGGtSfhYzMoo5lmCUbeyzTALtEQkWNf2g5he49dmwnm2UCB4M
8kMSJ6nnYaIPwVO5HQWGb9Ne6uuJZei94xorRQI1yYfIRwvX6ToKEHqLuahFrPr2
PSBrZv7orM/tNvTkGjemvAXUwc+nFsYQAqNAXpwTDSEbKHweMBVUPwtUBmEMWZ0p
1P96fcIth6qlqf4tdmYgWY52qOGHPZr8PXX5H1jcBBFKG5rdgzyGMkiTHMC3OqYT
058zexcL0Xd4Zz23ms9PR8G8T+8ZmlMIhFQvhveIIDDv/DEQEUmaYDO7tNNzQqOJ
DKRtK6JNiNy1le65Rhm9ZtW7oUoRpHZG0z0rTSLp0EYpvFFnYXoSQK3K+1oC49vU
l1Wuh1n2KL2I3lvatNEOMA==
`protect END_PROTECTED
