`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xr5cFYLj07yPh0608iFznmWIi8v5GwFGcB9Ldid1/HX0FjKKGa+ZMx7DYjJ+3C0Y
/KkR13L+jD2UWB7CJMK9CN1WxmMuyLTrE2hdBLNeMTbA2S9ABQkF+slJzayP5mLa
i/pkKIZ3FcE+p94EXbaOgJ6tqQzHud67+xFcvHSKpti/82EN7hRFHmFTqLoSAeHT
P0gocCJ0OheOkp3PGowjyxg20qp5wFhKB4W3gXme9InQJ23p7hX9rg4vFZIX471V
Km3wuOvLtFbMTszc9xicyeR0tJ9PIDX1Vgjis9VbjzaBrHgzfgRGpce6ifkMgLJO
tAN0yQqvC0lWNi6PITmNWLjQS0VVFZmY/6GwVzTv5YxZaHJq6zwptIxBI+X6IwI+
`protect END_PROTECTED
