`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFNXbhLX8N1UOutSwL/uN+ESQuOJ6QI93DwyklM2VSThWb6w2IsCMYIQKqEGSzvk
QwrCagym4yU1V5EHU5Cf6CCG6u4/N3L9QfXMtg63slO4S9s1NxpahHEMk+4p3dro
WPvAOHQP6b/scCR2Jc0av3ZUTDeDUN7ilEYuwweqbbUNAdHgY/Bbo4HPdkc1TGDy
5M/zd3/aMeLQxJxNoWQLwJWf8ZhVWSi3WpDDrB/GHKsBgeOCVNMephy7idRKaZ7R
Jd2Z603p4YqTi9IyNPjYRP0Chz0eMGKP0zedFiU6mZo=
`protect END_PROTECTED
