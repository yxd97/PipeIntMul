`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q+NrgJ9CLujBB3hRfAAGcdtFnb42lIKtZU5nM45YHFAfEt8rC3GJzuXgghikBu8v
vMwrvmBSZOYIcWQw+lSkFQdNly50rJzDjJm83YRTWCt2/JTB7sJlKXtpSnsxR9+Q
VUdYM0UwmzxMmhAjez7cKCiSotAXdjqUb8mRASuXLNTa380jnwhVapzIG3W+gnj4
ucjtgJToPyW1/yVGcH6eyYgkK271Fdm2rcK9R1Q5/zacReGCn5l7NR2RjKtFFbF8
84bEBrS4FuRbZOT0jZtW2zzMvYieexv6qeyxX3Vn2xs8KHS1UrcqTkyIadqkKVLt
pCjII/oHaIlI6qr1uAqmhJIgp19gRU9/f447orzS992XXeLFipC6jJBABDMlaBVG
Lniz1JMEVOIPz1vz+irGUKxeX0tgOWtef6LT0hwH2GeG220dS+POsp6JN9F68/kg
f2xzFmqeS1bDHR7EdY+3DbCGX+CVmUlN+ZcB9HQsPw3wkILNe5KclxNqtEnDF+6e
cSbO+rgT5IDiy5daWga9ts4ahDcDzKCpisG4wDW6b4FX6o0Tzt05tVD9k4YEUAFn
NgffY0tl5WTtafK02Z0rw7ib7RRuiZE59ZxO1519VSMrUkxpUDx9t/JxJd6MYyIl
ZMBi725HYR6WgtyUPgJYt0QwGu+Ve2SkIGkgfYQlMLbZBd4Jo352swiJPGwrUGtD
7MYMCWaWIpq+GhcKotBdihfC0Sqwqy487OFbvqi3ixYnXiP7H0s/U5bpBCtfHDrL
/rz39BhdELT1p6qhbjT54/IodiBOxEoTkwmXEgt8blg=
`protect END_PROTECTED
