`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dcpgKdx6gsel0NRedBTwudYImhdWsl1aN4FZ8RHGvRG54d4Ti1xqgehi8sYjcpAE
guNpET/yb10gk0ZVcAoPUwXGLyUKqP7/pPiwXBVpU+4cinabRVZ7y2tfybwi1BM/
SjPLtryBpNshSpCcB1AujgBnT/8ql8sfvPXdaspJyZE+0HXvWkYwnNlSs1+a1+CI
o35rmAUi6hDHldQbKc3CNfLY7u5+77l2NupKra0/L6s0hRCkvODGgZj46Q0F3AQS
4fCdbL1L37gYD5QNoiuiYJCKfrZifawLlR403tHjKbynHS0BO9jsNlYG+GurMKi+
K5a0d2d7FEj0oB9CRt+NQSBRG1Zkz3y/xeE9O56nTkRzly/egUB1uClYIfGc2jw9
FBj8YQXuEJQaYDy+2nOfxKqQ9t1WuLUnCiU4qyCa/sdOhg3I1NuME2q7C8kLGYq6
4ZCwvOExkkae/ny92Hb9yqTHTRAgo7JN3k/9JkQ288uUndFdzKODYY91aM5G9rz+
h2NWtg0WaN5sPOboi8pYju1vB/rPnxdzXA1WsalPKjO2sfDHOqNjf2RyS2RRZ+u5
vjewNKe3GEDQc2hGLh4TEoyxHq2JdO24XMpTBG8+xTATw8j9UBTIkMpfYkifR0mJ
mQn83II3MXx5d5IGky+5LhEeJNUvruU41sPxOS6Kd0Y5OfhH+4LXSUBYs0S4nWHt
1vXW3S7itrr0oeXwrjDGGoeHxnXQzY+gQPA4jzvVbxRjhOrvrx7/aKU6c9cFm735
XKgEcnVYRLisDSRwnzIB+CFY1AP4j8N5C8EpvRvaq2w7CKXMHey/D806lNGCGffW
nFIjrvMj+c+MbQb+hovUU5TzgHaz2DSDIm7iI3RfMtgFYAg9ecgrznwbkNoQpndU
A6H2JO/SREZKDEUIgSTf5kqzQywM01ydNnohLLjjul0ezfDguhEz0vutkGweGVt5
U6pKXOroiyKR4//qC6Yux4Mtu7uHUiLs7CpLnNNoBUKSHWz3nCuBEY/Robillacu
UJqGLzjwS+sWEh2casqa5BnunPNIhNnTxKkdqN0pJNEd+uUEQQ69LLhG4RS8cukr
ajWCSfchlwlvqe4T5yTGYlf/TZnAM72aoYl55GmnnWka3QppqKdkerIeRYtwDafr
tpDEMbTom/GDe58rmDOHrusBI1BOQA4bav+QVABRyFAZCj+ZPaXgpJ597k0Rq5oA
bMg8Ok8TaspQJ62chZOs0QRNT5WGTks06k4oCe9k2U9B5Awa6pzZTYbAO0iGyejw
i+ABdJYfnk6iixW+xe/TnE7vcjTd+ckAZvkUlArZei/Nb/j4OKWdhfB26K0dtPlx
iCfNSNlf0hMYYy3MkSYmpyGZ1p0LRxeD/VVGVayoDGom6rL8rLWxUjx2pmDgL/p9
k6X79YIpQ7Eujo+J8Zac84WvT2UKuOIMu6vcyyH0AvEJmqEVnAlcU64oBX403U5J
Yth7cF03CE/jaHucB4O5XFE08GEDvy04gFa98t1Ejm3p/G0Sr3x79E5TOJaK9m6a
WlrcgOVEmq8dqLIw6nQXKxFR/yS7Qy7QLv6egS+M04j/Ij2s7mCyuU53tp+0BoEW
+1mUTNI5/NJuyf/BEcpq6EU7i8WcTKfK8srqQzB67NGaN25Gq1J3KdFcKxIjKqbx
MN8g8uks0ZbMiLb5yaQlG1jZogmCTNmX3aOmeH5i3oQByURFBbCz3ljOn6BDux2x
7s0s943khWx321eGFCOQtPtC1TJaL4VbFhTVMDlyWLBz4Tc3rGwSS93eE64gp7j0
fcFViTlRWbah1QjnN83okkwFEzQGA7Y+ZVU+J75dv35E4N7FKPnILiffYKF/TYOZ
BgGy7g/Enlp7N38FoxQt8o1s0lbHzMWAvyXdtrRu5ZVCmrREfP0DIRzxvr+kjbVJ
L6gA/D/TlkW7MyTwJJrKYpPe7yS3mRK4xnVWxG5gPLxv4Gyoy+nS0Cm6gbAKcVAr
8UbwBsn+5bq+20bDQWZMG8R/CJT1EtZen0s9mJHwY89gOIY1mtv8xnNqgC3oW76u
pEW3VgJ70KN24F+xWyELgSPWkj0lFPimFts/9HAdFTp5vxIxX0wbRN1SzwQBywZS
0scfz7GPaZO6bYr0Mfp1RNGP0a2vxJOCpIIB4PnYywoDUmCdy/YGWAcgFjB7fiW9
f3dpq0KXySYjVW0cyqKrEldUmYeInfsbLOtCwyRKUtP84s7BSX6JIHPyqKw3Uq4v
8p5V5yTD189gcbndC2CvIbzlngap47x5xVNSCBfvA8wNKffIhrZYVypz8xY91zUZ
qYaymScLO+F9YCpsG+H8EubkYFSNVksTP8J3eLbUb6z0eQv3ZpIz4MwqDvKBBDA4
qQSUm9GS6XWhvKupaOKN4bYuFcfjgmodMuSMx1t1vWUVUZWfGalKqXhjwJaX+Oi8
LlZqhImrOQqcPR20XQ2xAodCSPDdmIghssB8fImC0cKZU5GXVqmOyW+qo5vEKXeK
maGgsqO4LLICAXJyjAphfBZ03X3o3RDgwMz7wa2uE8mpac1a8DqYaLEVIk6UrXYU
sw4W2iceOP1CvmHa0BDk018ZMd5eo98Q4OsemEYVs6yf0sIqwY/XwYO2ArSU/m3h
wuLv7AABY5/oeoqgycrFU05KN1F6QirqYkcJvQVBMpLaJv0pD6VtDSg4PwRJStpS
YKz1eAXIIkoNT17xF4a+Df8R/3Cj+dWK088LDjE6cN7yqgUeieNAt8i1SJbVUvVM
uDB2Lp2k032Gd/Q/+e2VFh9zGsulP8hCV25M7pTB8/EQpplxycbWlgK4EpbCxVfJ
WPJ4WZ3+Zn5v2btvdzj3YchxYleWO2bfhzlBcHHuTt9rv+r4o5TgJiCUnVE/2f2M
pT6XQfI/eT2Ur9wIAz3u32MHQlUuRG93hllC0AC4ErwnrfB3M2GK/3inmu9VDkMp
iV23tjyCFqCPbmPgM2sj0Iq9EbIRbBmN2gqEWSMizQwMmRG2NwN522oX/VIBlZvW
ReAtjH91QZRtlpv8DY8XSdYienkstLj0wMkLdyQB0nxNNoHbfbzOxuzB5W05L97i
+C3StIj6CZqZ4V51o51r8YlXK+dkKkg8bRekrN1B+H6d5dV5fsR3NG1JhVEI8YRh
X/UinMJk3C43SaXeaGV7MhSlwQAKYUu0mfckhg50lAmQZ08pxo1y0AaqRauKlhoC
bOXmH8iTB6Rj/P9J6rP19HPVlUkKojyHNiVQdRwlfulEOvk0J7PVXJdVUKcHxsAT
ZcGX/X/RAgqIE/tleZcMzSOHoSyDIFjhAl0dpS4o7r8GgSpkSBrXnill9EdQL64d
79V0+CzHuN5B/5CQU1r+4WfYi4Abft06RQdeBGAYndfrg9DqnGy2mj49yiFNhy+/
6Zk5rHiydRB3uF5EWcf2IutYD0LVNoZ5BhNFn5WwdSbE655SR8JtPx05RuHVU6zw
mQqGVh0N4gt2bIOxRHrNVXBwr1wsBucvuXlJ17lOnup4o8IxgRsoRJlH8UMMw6yf
kHJr6Vh/z4mZ2ENU/m6cnY0gZqVlTKo4rX+R6f+qvtsam5obdb56d8u9zbQJ1JW7
JLdoP8XPCQMQKdoJZynYnyDnxv5Im5GhBUL4t2Pxrpk8UsEI+BeyoNcy6g9y6DRP
X9W6/NLSUO5uFgmhXcdB+zxT0FciT/x4+3a9Obxy3OaDODh6420xVELm+qLwptsB
kiVY0Us0bnH1TD0Ybnhi2VgteC4FoON1jUPyCSudkpw+UQeeCCYPcpS8H05AHOUL
sYbk9esAMz4J8NWkRXAZQhsFXF3irAyPRF42sJPI0Cx17nNC0lKEFxsLKWav5aah
UqQdDfCyuUR/PauL/oS2UZtAc6TScUnSkqM0NH+HQl9EpiFYNYV50MTJXfxizbDH
97dTJDtL2vrFYfT701qhdxYXQmC7AGm0J7nL5v6y2SeQuwZULm1B0QeRV9N+xAgo
PSxF8lasFG5pezLTzRszGZ+jW0rW1uS5OwQhNAaA6qrd09Rpz8/ypOfXfZYHaZoi
4YmibDvTIwjU2AuLfhiHb6ZhAV9Sec3Kk2ao4LXP5xqeYPdEJBVOVaTJinRXDy3a
5zml63T9g8y8jgU2nfkb9yikqQQ85PqSSl7pv0KRoDWM2j+omsqwkemVqdKI4aLi
+OtpRagtLGQxGs+pU8tXsIdzJeV7FwEpcaxIpz69s3xWV/87v3FCfzF1pImZ5Don
8HctcFNUOIKhAdQkB9Wpdcqr3yZLFtX5LV/NNdorVkjJ5oO2iCW4h3yFSGxGr+YU
olm/hbcTpipKskK0XtbuG69OlHRwSw0OCzafDNotvc9D2/Wtfc7EDcjViND0tmOP
pP1BggSZOA2eYKPIiJsdbg==
`protect END_PROTECTED
