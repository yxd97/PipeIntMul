`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hSlYdGDjdzD8R8r54moA8w+jbGhKBMHQl5EHf5vLuzFO9t2o6IuM7ibTa850yOK1
6b5v+YPHH6akd/61u0IWmxjR3eKlSiNzsLnWvhUIWPySj7cAk7jMHoqZ0UufvvNw
0Wja5IrpJ7sintq7bpNLvo1oEY9R9EZIjw3RpvqczUaGObRshknpL7BfEUZWAkIN
5z/6IkgCpkSeuhftryVe4ziq3XhrSHDAElw6sLkYKAKYWf/SeSRwHp+UH6jzZR+9
LfhuudMXMub9gq6KgToLRYHZx5TXNmLICmcpI9XovQFPU2K3Le282091sDiF5/lJ
gQHPtrrN1zLUuXkfyHfYEIbW1Sgx2lXIAgv74t+EXIhUqlHGvHKIttWHIFVOsHgw
BsRVlHVG+wBLAxZwpBFYjYGq2avrzbHeOveEKtRv39ijnhuSmjZBvgGe3EK1RpW4
xPJGUMRuUmXgoij5QfPULjLquany4lfYNbsQnfxYPP43mxGlaqS41AeJhm7oTT2U
kwr0w1L2Lh0kbHjMzkxWYjVn6grAIHVFI8CY7AM7qkgUSF89CadYWP6jNuGmr5ze
uLTng94HoCOpPBdKGIxEByxamU6vnnZWSE41gEUrenrZkitWLaXakjFSzlaF1MiK
TXPOgaHw4f072K3Zvz9YqPANQKPTp2L/lm/joB9Poi8=
`protect END_PROTECTED
