`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QgJUztkg+bi+bnPL6nt4mZdtIh8/CNQiblkF5ZzlSYvjnoG2G4e34PszeyyyaHOJ
5uxZaljmWwldsOXCiekSCM7xIV37kUu3R7KBN2+wkq18UbZF+YiB00hAQbzvFC1c
J1yVwrNGH4MMm1t+a+xr8PgGcWJzET0fkUVvF+O8pLWB26VTcReEouytXBbtWCkx
77/pvrisD7xf/0c1t87GDYP6slC6tH+vPWzANNcaI0FFaa1p5CMB5nqAEJvX0kxz
hghwyHcmwgXcuFgUoXDvSZv7vNkQZPcyen6e5Bj9H5onYicx4TE92xNVkFdhjy1D
oOfx9azfw29KQ+jucUi4NKbDQQODKjCcjjl1+qDZd0ungHrmCvWREEn5/WH8vih0
7U38KCKWEfSxpiebNOgzNibaWAzkpc9PJb90e3P07R4TcFGZyk4H1SKaKGqtYf4Y
r7kCLm1KUEA2kvEVd+//WOQw6YtLY/yzTAXWogRuqhSnzQfxlMCzulqbp5LzZPXG
WStOpONmoGhEbFzpcw52ew5LtULAgq2KYo+aSZ4YBLJZwLjF3oS0OloE63ENBqQO
h1GUcstx0Mk65TVkLBYCMl6K3isRIGo1g6cNlN/50Lt9c8Q1XzEP3eyNPIhuM0YE
FE5Lv9I00/Vv3wgPrUPoQI3go4MKLTNWWTB4R44CGNNYeHH7gamzP160iJhcU9C7
NrnYxuH27525KhLP8pxZ3Y2CUXlL0UV5tocBQRRJ591u6NNFxjECafs4el9ApE/L
zK2Zwpd8gb3Dp0PgjH3GODzfraxzUeAsRWNeHEV2DMwt1NB7j8bUBevMAtDQyGO5
nprIQF1fGHtxIaAEfomxlg==
`protect END_PROTECTED
