`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qzyTZsqfORoCzG1AFku8FvX8B8s0sQx4jCnk3qnzWMdQRu7V0zIPbF1UE2hWP6U
NcIOCMhE2NAwephYtEnqqDssHMufCAFy6LEJLjsJbrFKqaz46jneAOwCYLAI1uQg
/8mxu2RDLWI53L3pjiElL4/B/YGbKARgmisLtCBI28oZnt+RIX+rDv6lRu2go39T
0JPpH0EGNOwSO621yXvncw3G/tsQkbQA05B4bhcMGol1ZXRPoAjE2zkA1EHDpG81
OLc37P9nPTLaRv+w5SNcDGGtuLfsCJ6+79VEDSVxLwZFtycsX/DJHbEZ9bJq9rD4
zMIvkTw2tP8gyXfDaXf/xSQRP+jnTMfL8o5KWiYvJrkvDtyTQ9/riNCcQOJQhUeZ
Rm73BzQaEM+9iLa0+f3t+q8wzAt+ooOJzhXKGNQMyxpP8conDt7afAD9OC2P7tKq
OYL2xBDrnqpv/+vOBQAV60ExyaPnhFfQ86IU3tE4CdXCg707O2tf7kHhnw/jc+eG
dtuJQ05yyuerXa6zRchBbXrJai60OM243zRZpNYRYm/ReUWYRx7CIrMEW2s+X1lS
PWg8gqJjJnI03w2BJhTqkAoYde5GrkvbjaYM+wrNRI2N0DaMb1E0n1qEBeTIB/6C
7b4DL2WmWQT/TG5dPB5pr2BMk8M0HyNSA8CGlTiNEnFJumWMwtmIjQocTQKpQUkA
u2LQFw127mdN2I7WUy1VXcY4duBmszj3XNlAxUyqPYztFx8iWCZSdeXmTFUHUdA6
nUqYTU8epOGjnKequM97hgWFzcgl239tOXpNtykGToLomMteu5eAj2hq7PDcEX7o
7cU2O/KgsMKIMX3bjFGgNKklF5Dz6s1ydhIJD0+scgElClNSRWTTa9aqlbLafXE/
Cd7iD0yvU+rKOAxd5bPj1o701htPK5tuhsSK48F2W282xEHU69+wdj2sKf2rs3Qm
Ry/lMAsb7WfxL2EMb8FrMVjlQZLw8guZsoG4ZOG/T6Qo6kIskuYBxHJENtrhNJkV
Zz63nTMgbw+Wjz5o1F/e4kDtXukYnZVx5M3Aziw42krsKMghKIJaityX0enJLZfo
WrYWBrJAipoAYYsavPX0qps3UqynS2NdCka5Tqr2XPoKRuuyq0pOfTTJxcMw80yh
c+BeEiFQjCs9TA4D3qMowFAGgw0A1zI0tWyZOrdu0ZlZrEt3EVS0pI/amZawsB3e
Nt9dd6NJBJD2ZiiEDawIFxuu4bgNiRUy1ia1wSO6C1xyVb5UDLYG9Fp5dHeEqZhB
+LVFmgnrlRpjFahOTupIl5C/0MpfMHwRcaI0T+VDddhg85158eAAZ1l/mCiVPjrR
NX8F98OQKgxYRWaBPf1hiZm3BPQ7+lHohMTiNE9QxTI=
`protect END_PROTECTED
