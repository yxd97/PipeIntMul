`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiPhY8PiFVda9Zf+nOJQYF9kcYCJt7jgot9s2aelWhsEG/cg9ghWZ9/pyKaDgrjM
oDGbv5/c4y5+U6p/kLpwRckganMq/B7Z5bfpIWTeovPEqXbip3NzXS0uuxX++eQp
T6o4ZCWMijZVTPJKIa6XXpdvV+ruwrCdOieiGh18nZ+480tCE+1MIJgyx/1I3pGt
bIxMJTsKEzNdAFT2lEsw60DpIr+CXdcbAT6ZeTEA6KFM/Qmwqyveiv6BqQK+keuS
LNdjpjID5pYWPKRBZy8DQejUVtEYA0JlvDYF4iqHxXqMFMZwsmwGUr+t44RMzoVI
1NtuuiajtZv5RBMWrwgoYyReocUpatANveNAlnakD0WgBWE0k9++9PdVedDAxwT6
7Ns+Yg9om8LMKlphhlZ4Sal5W/lwicrQqKizPBq3qvf9WZePNxvfbfQG8p0D3Wtk
IOHDapunVO5ey8SX1TD0EQ3UK/oTCi2sLPZibuULjDj5LrRnzLZ9jbj53va+FSBy
1tNA6PLK7JdhrnPaO4W7ntJ+g8Pk9llYKGE6yxb3zpXtuTJm8jqSmuM5ncKsNAWi
`protect END_PROTECTED
