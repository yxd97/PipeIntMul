`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
10XR4aZ2KMSOL3QPBuJF8k2ZCQY3oX0QNZVZXd9cAG7bfcrDKepi8xtyzB/PFG6K
PZhCu16yYbdLo2rZnkKew2oCTwEVh0RlsGT6i7JUmQKUMjAyXhAYOQn8B6mBhm5Y
Tn8iNO0FT7jHVigelOB6Uy5CLuIwkSkkw/jD+aUH0yNP4CMMaDg7l72ztuZn78FL
VEWABbAiJjr6CuWsk511DcObMtQZZes9Urf7+ET4hPUeo6BjOB6pDyuFTftUF/5D
mDKRdKR5lcfv5e4NFs5BMdOem6RmBEeUve0z/Khr+vxdxeTvFOo/lg5ytseF3vno
mcY+S0EAGSnuA+JoocyR1xKisdvMBABiEH3CPz22WCWT44y6LUNpYIlvth0nTrjs
zWG2uhhevdcJ6sjfk+UILQ==
`protect END_PROTECTED
