`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ULOR8r824jlzcTB4MP1KbKCwpNQvlXUjvaocD+NSdDrFidrib6lYB1hIMvPpoN2
wKYi901lbSirSvGVLCxKo6oZIQ8sTyqg/Kw7wxWU0atYA05EOB82cChUj0qI6nz9
vM1kxQqPCeUmAa7nqp676hHVsFCVxrnfduyCAphilyaFY8fJogGMK0BF3KLZIm4T
mFMNqx7EaDBRsJLABOOOLvjX78k4wxxyfNaNQj0EwqA+2kK1QBRj6Pu35696dum0
`protect END_PROTECTED
