`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UoHu9j9Vu5SH+nWGOiYZe2BJcwZ0SrIlX7WXoBE1rdUTEqDDbUnVBPemYpCaV+Bo
NNEM6UpcSKar1JsZbDuFbGFBzPJkL0j6CbAuMDu3Xlw6HDAdq8KGB0KkAv3G2pzi
7QO7cLxwAHXacHPsCJpZ80igcVRv3IxY+oXhbol7cGq0ljjCIWeNR5eWo0JCR6zO
Wy7+QHUpt3jdIpN9J3sSpjnrzDkS4PhQR4zjGngttmO7ya5IhTmX5KgcEireKkw5
rgdpoDPw8M6mPlstyQJB+wBZF7Vqe4X0NYfGwJqP1/Og83uHAx51wPhD8jz3uRSs
er1rLZOZ8dzAA03hdYBATA==
`protect END_PROTECTED
