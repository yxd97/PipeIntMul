`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SxI8+dTcH3JVIW9JjKoRzmpav4RjjNER2z1mBb1YSTrMZFNwXhXofkJiUpymLppX
XyAWFb95rs8Hnl4uWgm5QNzChI/WSJaKo97bLmUnS3+SXn5612DSCcuZql4E6yhW
m1b98XJVfNGzWeNTxhNIigacrlKha77C/FCq7M2WuMquInXjU6WUZ37vkuS71gPv
VFccey1D8fuaMm7p3yaUovZ94T46tN1Rbov2B4RcQW0e1E4SuIL1geyFQcFHL/Jc
hyWldQVj672XFqVpLq9vULzxseG3iFly1YjMmYPbmqLhtnRoDjcXKCrAiaIxznBO
eBuNxKxJhYhz6t4fIfST9XNngSr9W74q3GuWCYNwcBvopFG6uvhL19bs7qVQcyzl
Ux0eXTKog00vmQCxxkFNB7ktuJCOc/bskd3glWnJG3AcplavVvGrhGRazoNEoolT
xEEky+nlSppWRLyII1iiKZUfpwBy5ikvjDTBt1hfKHIW/vRBYePHxEfbTjIaKIFV
BjNr7Wwx8Hkf9XwbFMEDn+TrL5WZeGUpZFI+iPVMxxdwxo2BnDozrVXqPSRTpoJL
pF9SZ2o7lNV30BE+ISPavZgM9lWKa09yKwIFph/ovhEXYKTsKE+FOFEazMxw8HQw
gnhvKqpQbDxMdpJ3ZJQFUouK8HzJRmuRxR5ZuiliIE1CsLmnfCY0TlHN90uuygPE
t0F0V69Mx5tu4rMiFSkLofypuleWwgiBTY8116rSy44QyMHAEBD0HC1iesgQ29oS
y1gjN0JoY5ieXjykltpcxqzfZHNqt+9le76mxx89uBlvTAwUYK8YUFbLXATB2rFd
NctPRo2Qfaroo6v3EpwFjAYwUR+0nXPIc5l+vAz9hbE3DQdzNa5oQOSe9VZyGbyQ
raKMjvAMoPHxWeIYuFcSkNLN1FKywBfKO9mQEA85wTu4v6dVvf+Z1aAF5L5XWKZc
lAGeVAqp3Qc4iPcWOGDDPEZo5mJFKFaPhSp6H14CKo3yZgVSnXMEa04ZwWcqH6g0
oXmp/OUkqo6pZYQwC9DKuVUqdxihFkplXh4JIsBLh5GBaZNqaSltlp+vvBScCWB2
2hu0wVv6gXGL3lUp9DejafFRR5U1AvKcQwVFXf+J6N7hFwc09SDe1y6rGUm93/kM
tgHH4IvzOMrT463oRGHwpQojm7tSep7U4OhYnFYIa2CkCLKRh4Ta64zsdugaFdTn
posVrQkcH9m9mWeOOfDexmuQat+FlwzRuxZP9pl8VGKQzfpJhw8Ly6LJIQD4cck4
L+au9OJfj2rr7RmB0Jq3PRgokyevqg6Rew+1IrekKAU=
`protect END_PROTECTED
