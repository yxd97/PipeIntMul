`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pdARrpnSHXRYKrL9jWeKtx3eY/3iL/hMLv1K3QVJmkCh51gXCVVkAX7FFKE6AXj
2YTfrquWH+scdhu2D+P7jPDyMAsUHIWTaifCCNhWq/opdgjgOnD5tihltrVzDGVi
4oiNiorolSWw3s1jFZF1G7ebPyw4OWn2ixUw6CWqdLEl6ZSzjm7iiWzcjAW1C1/u
e/Z6I+Wl43YNB/Pk2Xt0tIBTb7Am3dvL5+G+Xw/qQaWw8gcMS2AohK7Gr/ZfYkpk
0fcnZFCgp69Nioony4bzqnVbc2/2DMCs0mkiuImyeZI=
`protect END_PROTECTED
