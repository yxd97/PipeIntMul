`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uF3RtBJxtrb0WYK4rTZKdqojnvg9/UlGhG/weGy1WUNJ/PY2dFF19WrdIjO43+LC
1A3JvrS3lSJSLsel7Obqe+dPvrToE11ekfF2yB2oqop9FXzF8y3BkzS9jSs1Nr7S
+ANxF+DHxd1EGGlwHGATkTJOwrQV4ImIGzXzlYIlMsLRGSsCTUqRTqgzl0Sh3xtX
6P3uIZ7WemqrWBD0ZZZRQqG/WdjwXWDjbL+LDV4Uu8yV1zrHbQEJVEVORVWetc+w
TWheeJeQ0V1fAp5bLP3mYhzlq1ekLprJrheAvEomN56A2b7YI0gJxPpCIirMOtM1
VzV6P5Fk7TrMrrvh3HmjKEk65Rik9JGSF5HmBFwnLj12S4JH5NKG7W+uiZzai+bC
er5vNf4k+myjdT/UPWkXFTLcSm1S09qiNEXuTybypc8/HQnEzmzqQo9//LGTc0Vo
9IOSEIkiFgB8V132P97CS59M6+HYeqDSOS6m0mNIlgfMJ9a4D1VHq2Glm0+NsOwn
`protect END_PROTECTED
