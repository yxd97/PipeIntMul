`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
trGafu0Z5wGAfqizsgm3o7DbzOt/kJKEjw5kam+6fpsT+43Aa5ptQ3S5sHVhANn7
gt8XDJ+VCxGOl4XKCIpLq6D0ZZV3FTqZGt97DmkET6y7szys24SyRh9T9NJj9EGm
mk98WlqxOp/eBSD24gc+9dEyIn+QvmhdHcEPY484FPMNAk9clD6wQ/bR0cmHnHFz
md1FQmMps/e1nk0wid18DdRbN8YUcMku7a2eBiCa/Lgwmijo6GCSZgyO92R1wirP
/Uanj19TT+u0Mb5Pt9IFZUsDVAZ0F7KkJd938qgS5OeDo+xkALiTfmuWSHblYJP4
FlE05Sif2hacE6Qd8ICFaKMKc/sD+IodHn5O95FI2SDl/ifW05WSIbcRXX5zPs4r
98DSpeM1k4BAF6xJG3AAUtGGhYKD2IdRQi/pR575neWQMjKskHnSO3H2qFu99dni
4ZnoNHEwR7wbQrKVtcVkelK16FwBWKSvk02IvJ6uCA54aNUNiQLmFwhWXLu1V4hz
hT+uHgcUEhsSEg8KTRVzCujovRYZOGBpGooilCxkr+n+ZJKmrIuSjeKi0mHPvLMd
sCP//IbEmEqMOdYK0qd/F3TDG9/y/KrV4ii+smBjv/3NrQBWqHtZ+/SdGQgew9dZ
kj4ZhNOEJ0xDw8X3wDIm1PcanZc/rS4b1adpXV8pf7aGm46KD1z5pY0lEEsgzFH5
ekvlpWM//JeBixgEa4gOP5Ko5XcufULXDcKBJhjbxSMNw4mU91Dd8YLaqv5mZ54c
RfWOI9hN+Vc2A6Sh1kP0lBm0WRx/x42ah/ZlUGuRwQHiNNwsRfKkYLBW022AbR9V
lsqLPWa3SSIAqs20Vd3/hwgAHuH9iBFzpHRkHJ8cqkq+0HQ5kfB1nk8FTYe9Bdjf
T4stsvMOBSNmhsMx4oUxq4nxPNU2gd5OaydadUhhS234Vz3jf0muPB9PmsVWO/mu
iESmsdL9E05RydvCkhtWjmWpkdCURgFrK8RgOFIgkF12p5K1ay7mLzUDMJMvcXrO
m00Edwdjw61qWTeJUzietHSvHiILqiG4xvoBnOJXdMFFIeRyFc0AIvdY98MhBp9T
PO23ciUG2/j6+Udppp26wejzrr7O7u+WvSq2uUG3wkAA+2vUYDy0f9AR0tS7oFT5
Ubjt1uqBV95lLK8UIexL4DJFeYZWmnjHbhzoxgg1Gx7FxrmlpqoEqzCmRLSK5SvX
W5m0kQJ8AKxb7cnZiDDwSMC7tfhz/DSa9wF20MRulauPKv/3+VU03OTwkJOLMe/I
7RSORmQ0WI/aiSKdfkBMrKteBRaQDqGsodUCBXy+GAs=
`protect END_PROTECTED
