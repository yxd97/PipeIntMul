`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35UpR1PIKn4xso4mzgjI7ImxdjwsUHtpQpt09+KZVI9///+A3H4Da6GFGmollB/3
nf/aTulwgkRFrWJ8O6xXufhh4qyEKWONYvs4bRIT65Yja9Yv5M3mPa9AxYqqigfe
v0sby9E5F/l6LGdy1x0vj6XNxSiJbqCCa9iwFb48rSW3UAZlUS/85aK++ayHjSTx
oUr/E1i3DRwdjXXVtgoChA==
`protect END_PROTECTED
