`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AImL18fPySLWGBfXqKkEB6E26vDdUAMo3fz1PRTsdwACKFtFl1/vAowR+DHRmIWZ
iLLoNya/nluRJjuxq7/XdtFTVGQUKtw3tBg3130OCYAG4biBjqp4RRJcg/DYMfyu
jv6K9nU1W33Ev5a5XD66KPBT7vS34jlQNicXMd8OTNGGwBTWwhcyNnPzJYSYjlpJ
wbiMMg2GjQi0e+Fsvl6yZQUVKMAyPh680Ki6AOpCKmpl/bq3zdvtO7zZ+LLeC8vW
0F1x0momq+qx0xqxQIeHz/AkxTXbnskXPhTmBoIBGQfPgtWP2lAFywF4mWH2Ayfy
kB6m/5UQ/i4qocfbX68WZ+loaYbxr/bVPmSi3bjWNkNRzOjMvV+HOxxVFXu/+HAb
WFOkp7cmLw5i7nWN2TSnWlZLeVDT0xm+WyLgRaD0pkPd/li/d3gvnrc9jjJq2P2k
syZKYW92y8cIC36OXdonYa7aDrmgmMxqK+M0S57PpCIUKfQ+e8O8spoLrdtb4Utm
RnlRJ8kKgWvUDqJmqcb5No7cTyoWJmrIWm+q9GEs13U=
`protect END_PROTECTED
