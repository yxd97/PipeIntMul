`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4kuJODfhqJ0wx0MQGQNXTfJXLABwiaOggRGSyCF0nMO/YHcR/3KmJfLJNpx+wVkF
vm85OgSBIdWlVvsa+6RfavlYKLgLDmJcVFw+h6c0VyDvLDgiyebqPs9JEl/3YKYQ
1u37NZwGcgUMr1Duz4URdyX69zS+3clwjp8W+o3cnwhpLDesJ+N4uECDRkgxRFeo
g163ECEr6C6pzuyGoYIeKMkTVGbfMSDWXnNppt9MhyOrQp71OZ0cxwp2HKXZ3kyX
ywU98i26IzDtkUyZ/xdkKQUt3ulB6hAX9dLFGbsBc7vjQZIYMVmBSHMs1SzCdYm+
rgYUEB9hB4dwg8gw3FogVE7ioejHdTuNy1eJSKyqLb1Y0yP0/vF3eVNvLxHmY6sQ
MNIGF4/2s7wtKk0fcO8UHxn32Pc4xsWqpYFGc9pGEMwwo6/+Boz+LZQaKAisOR6t
`protect END_PROTECTED
