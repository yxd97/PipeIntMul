`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KV+1rQGnsXhnh12QKik0D5Yam97bOv7C05LL5EQWf6nzdr/1Lx9kSr6R3YX1kHiS
oe/FEeiwSUKOfC3qmUI6ZA1eubY+ulLzipwpt/8ohJFCwQMvpyKnTFMSV3r2Xnz6
Cjy5rTx0xHtnzafXbC3nQKhcaB0uwOw4Eh8LrwMUtgCYZW/qybufjkRNvAas38Ko
e+taKFKTOnmoG2h6vlEEY2pxVHbUPAJVelwH2XIVTL/1j+SSNWudWyHAXPBsof8I
XbvqiYkxUEQllvk6CTq3Hg==
`protect END_PROTECTED
