`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WGLdbeXc7L+FL14z1PqAyJBrlCiTzUftRTo5+33Bpr8OZMCr25lPaEcTEk6G7JhS
3brQQ1BuEowuKywbVec9Y1K6k+JydXswlghetvwsJz1AGI9U1dgUWwRfn0g2Afg9
EvpbPhp0rkwEWOnpUYwVuvrYrdOp67HsrCOG7oR1a7q5y3KB/Y2SHSqT4wCgkIYq
ggLhOMfIRUwo9sMxqTYUhJq+byrHAOCAzOCayj+OqOUkN6ilmfW9V7Y97EyFv1Tn
N9aGYhi/4W8VNl9TDLktMeAfJQiL83h3W3i2hDlCwk3aO80rF75YOfIu53daEdfy
6tGyj+KAHwY6+gmS0jM7A+T4xOvuVYc1frKLIHeyOIWutVB2DGDDZ5DHxF6B/fvv
UcQ8NYmTRo4ykZqIhi3bGprm/jzrCQqoI+b5fJvebM/KMgWHdSlf5xpXA4hSH+aj
sQoUHzPEaoDfwzyD/Mxw4u1hviklXQ5oWJ8lZedjs6HADSyqzQZLyEj+V75O20OP
85Ynrjjrgf6RyWgejCUDK083XsKx2B173IWCINLE7LASZ6HBN+B1Za5vbM3AMFWF
v18zNEm4KpbZiHMQR8hytwxnq28i4daCaKNsKxZUDygPbmMLAzvPSlg4ZY9crMYk
LbGYRSGMe41KvrESraGQlPBiEpg0o03qYiyK8x9Ncf5iuwdyOiqanY7I+mSFf6a/
dvLEghX2JHAiiC/X32rIqg==
`protect END_PROTECTED
