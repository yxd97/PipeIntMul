`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5JQ7aHl5w2G7B3ov2BeMyJPy3Q4WUDAtqfLP1a/96Wxh7nD8T8/tcv6buheMAOsx
+95+BpXkMtALN2XeER/aPzrHaePWwt9d9vTzxDfDIkyzC0+VTHdE6rEtuMo+nEka
XbpG2CvOGIPmcpFdBBio4WBdaZY05yPT+4IyaxX8S/9LeCNNSb2Q0h/belb5Qn6F
mbmahuP1jNIC7lGL/cF+dDW0PyrcyTArFR0z64fdG3lSXX3DsIQGMnISEox14T8O
2ZQq/4CdWfeAddTScUnFdRz1m9SifrGzN1EICfcTENplXP/VEvVh1BA1rxYZ8VEX
zJufYVpbct1Juoaqcjhrxr7ajSgQqzj8wIzYMWKvQ7YtOL2e3kqT7tigK/4B1Kcb
sxHScjq9Rg4xlk04y9Z4BZLl6oXU0O64uUFkrIekC55+Ld4dafwqA/Ko8LIKOWvA
m2MyU/XOQ+SGaV6FR93DUzDDgk27kGi9+PKtIEiafn9ZX0phTsqxBwVjN3AdXOzH
Kyq4rbg1yH40Zt6OdO46HPwgq6IbOwKfiHFZkQaC18H/LuUKL6vziu2pMSf4zTU0
D4p0HS9Ql5KrkmV3bFVvihYNSniAB+Su6oNcb3tfb752HTVywOitRjcyETHfikwq
06uemrFSgfBRxIFfDQY5CRhMCRbjm0i6ScbHbWGWxizo/l436PamahLHfZ/Xmw0y
dGayo9JTbbdn9j6w5NDtbwOZyHGD7ji8uCqllAzrbrzdUeTvx0bVrPVjZJwa3EBl
3opvKQzL7wndQYjznQU/PkkKsKc9Y5bafNPNKXrpGlfNlRu/pW9mwyBj4FcD/HN8
YP06uU8euuGN4mHPnQVET+rZvLpbOKcAI24YasnIO9FVouc1fkIIeGGAoq46ksD5
N4V2BMMb90Eqnmuuw3Jk/w==
`protect END_PROTECTED
