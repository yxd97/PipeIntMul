`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
el1QgEZ0CPUewlqvdQ55O+8B85/xQJ4bEro8AGD07Uo9fUOyJw45QOZurgNctwAi
zGvaB17lJXqp8Klsj6GEZOipsS6zkV1egb37Wep5PZfatJIcGJYnVjT8MUT8z08r
j3VfJ9Q7zmDdJV6+SLnWx7IBuv0mpB9fEnyGc2pmtVT9HePMytAsv25NGJopy3kR
ZLoAk2FAHKudusyhkM0ljaIjNI9muu2HPqloM0tTFnYGmExXVInYSh1BmOU12yyb
ey1L95Dt+Y/cj+9c4SHg2/kNwA4696B1KLKx+0KzIpW4ZTTbm8hbWw3kTPUuaWi0
AkYyDAkF+ETT2avEard+E5cV+LhU7XApU8O0adzAvHu/Owi9oYVnHvh3m5kUgypL
k8er31bNT3F7OB0m7wl3skCe+/Ef9eiAllDdtv6XFfWUb+n0JNyn3yZVaE3kcpC7
`protect END_PROTECTED
