`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BJctN1uk3Y0voVEaocu4bGdFUJdt3U5a/YSp/ynFzJooszxCYHpwBV7M8NgTaMW
5mCxIBhTfm+RaKO83J0wkImIMSz77qunyn4BkIg4L+Gj/kcvOb0MN6XJFORrHBBD
x5lI/ER7VsmVbACbuAQlJ4qpHmdqyQ3Qeg0p5yJXFeh7QbnuNZFVY7pqwqMlubX6
mG0hWDCCyjqbW4i3FFevRqzvgi3mTBCpqkaFur0dMReRAX/lJgZounZWmu89AaIw
TaS1L1ifVEG0x5ybtvYoPyZ88apmOLSL6A57xnGdrTy+ywgxydxBEDOd8Z6XLvHL
PgGZ/UCdERS1kn/U4rmONcBuycmFz7kJ/cDTsmk6gTB55H0N4ow5bmQCCIcvP8GM
IKn4WApiGwNJvNNZ4emtt4/rhPieZgnarB8p6o0RFRtWPCvtk5MwQKg1HeIlx263
Po0I8vI3jSQC3MZ1UDhU0oTWPBkHHxxsITANa5AuyCmTZScgzSgo+L7rw9sw6ErR
ZEuCzkp69GhAJEWXkcyzJpDne8xFlbiQHjQFxEQJvOxGL/cqVMeV45gg1iq1Csgo
r8BE3iXJOnWBOxfBnFkvSfJo+WkeqKHuSsHyBJespp5FZHr3w2uers6ByFJuyoGM
wAPrm3r2kF64yv4stUdHzFT9O6yWhgbiBIGdCKJt/CuEtWQaL1+n6jexGGF3ENyx
dL1q9wIthFRNKO+Rzz2zPneiUJ76DVzxwlWVeRVDgHcsZ/FUNDilSsSSUGndADj7
qCX+MVlHB0tlyMzeA77ypyaR89gu2ZpnSR4PFLoidN/We2kJ7FuZEkKgDYspF5Dj
oPsYwbaYO9X3z173xhY0L36TJ8euCCwlbRWW4dwXODZFTT3Aicq1JVEq3wkzcVQd
geh/1hLRHfQzrnyR0hO7wldAhJSbY9ne1XWvB0ukHQQsrH+lHwopWG3+wdFxDjaN
KtZ7Rkl953CCOivIA2odI9+cewZWX+DJw/K8PsB7AYfnKk8019trIq9r4RE5I8qF
5H4amKUucMmb16DZmn779XGs1+QnxBDG8B3zVsgNVKRSY/VrIEMUIzOiwBnTFgck
1y7BFMhryBhY93Gt4hjHGHvH02AHaGrgOWge2slqRm+0f3z+g1VrdB/BhzYuEXfP
4xxnK9V+5U6j9/FOXW616yFDyp237nndXWKgMhSesT+RjSfi7InLLqCeJ7DRYJMW
d68qhVWS5Lr1E4yQZP+eLF9Gzl73IOmj3kUOUJdunc+tiWX5oFTIUR9dKGA5DHk5
UnHHNktShm03adqnhfEnTeQKXSWk9AQQdNfJ8fsK0hbXJEMKhJ1KvJeBagJ3xJ6r
YZShAbDjxN5rexlv3ZqKwVPv/UqCLAlvn4lCO+8sWcmedOZkwHH1BX0bKq1at0iC
1XCnlC624zJlL22/WfkLMe0iNUGxMszqO5PFnzVToNlaVWef2ypU3egSCmmMmYJt
p7AJimy+/5TtgoWPHeZXzw==
`protect END_PROTECTED
