`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSTb/0iz7saeb/J5GNGZgsgWwEuLmdioGUX4n5/R6aiC1wtG1gBYzIUZTlnPqFpW
lWbulUuVwRgEPfDrMAsDtEuAniPFQwb+Lpyjp1CDhsVz6iVkqP08BNbmc3J5/Zvo
mVe/cA8TGMEthl0gg9siwR/9zGOLL9YgF7lz1djxXzIIzSUhnhBzi98GC3jAEGxW
PdZhQXqdnPLWR4CrLZn1HLrtmGL1tAaUHOLDePTC7d3bQVAna97cfAJQBKCFe7ML
eajPpzsYaIxACMpYrrRTWktTL5Y+Se8QGO1Fo5aKidprWywI6F6+rXTe7TpsIMF4
/gE7TdiYh+ndnN6RkjDLE6CvdzQ+UqFYR/3pZkC0Nd5JBFUe2ptBOXk6B7KZYhO5
gEhKkTV+IFqHnOFkOvuL7A7NZx2R3NGOv4xsRGDx8LU7fEhA3Wpl/y2e+iwi4X+X
5JPkstWGMf/vkZXMr6CY+QskkaDDmSBaA1baVT2jF4w=
`protect END_PROTECTED
