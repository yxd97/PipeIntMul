`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kAdvrINt6f4QGKHLS6nMyC5dScuHdkZ3VVd1kzrkfpzImTKlL2ODNFjHdu3vJ90s
EJ5U/wQ0G4WViGUxh6ABH3iejw4E3l4feJ5ZRGMcDVZOONjKicLeIfvD6v02eM9l
voeB1iTBA0LcATvC6Cb/8XZSXnvTQFqpPyZMEMfSFJBQMlUsUoIqcVZpob337N3+
BHeahxokQuVZlDjVw7NrjIOtSbKGfZeBDzacNNgM+O8pacBZGqFhFrenzbrWdq07
Snv3dquIgZHlqQxM2MKWRbW6lYaI4dHFWgxRlWceT6k5lgRADooMkt8XPRa5X/CX
9hhbteyiQS6mCcvwfQjikKLUC/xjYCnpwICdpJFmHB8JqqJTpovggFBtv6sDgl/O
Jw5S9zUnuJvVZEn6oyCI6OX/9GWVQjTivj4UZxMVUKhNO8jBClu0OIUjo0ZT+7jd
FeAeVcfjwQdp8r/aMsyCKnvLxf7qRGjI4BWB6kh12/oG/Apx0hWqCKJqpecsF1WQ
0C51G/Co4lQ2SrbKTaOrYEBAifzaYWw/PouxjaiCkVaTLdzB0Cw0exzWhbZHtb/u
hdtG/6iytd4/Yr9Cfckt0LBBunid5iHsG286oORCg2EPmh80JaJHNdNg9hzfIVMu
1JX8jBbd02GhedKZtVEiNZUKWsDa3eP+zdDaapudAsnxVlArkfR+dCjHuzwuDiOK
8BBlULi3kMhXevvaDRKMs6DRK7Nq6cRVqsEOonS0MhzAyFezqMgO4m2OAO897/ZZ
edCK2URrdD5DpJQqFHrM0nLhB8H0FFF9/aU4NrxBoSqoHgJVeBwwJUkgB03ty4D8
xPrZlCzRLY5saQR0ad5+sLPJuXOL5z4LMuJf6ECRntCMWXL4RlaNo8e7yB6CSLRV
EHMk3zOufSVFCuKLTxO8peN5SaKHQDkSmtD47te/EOyhENVAVGxQvSoRrK2GtN/M
aJWe0lYyTMpZy61noBhgs0wjklvB599luS6lz9omiLTisSz+PUDfE6pfCsr8DDBw
uoqIuyAJM+SgidaCHeLVI7eFFre0QPYBCan36D/Nd+HIvS38SqBBgZ54bJKLv0zG
5Xg/vFuIYe6ZCL7SW6nVpThX+cAh0YfqhNKzxSE19/bkngcl+TEWhVPTLrgOtjUq
B144usCYp05s2j+55mC4L6Pn10ZQpEvM2X567xVPc343/dXtxhZgY2N0ERIsupD8
L+Fi21xT3MU83f8L7e6HtrKgbP7VWswtDj7NgvyldxBRhQjDaUy4MlOKMYKEyDfM
qEPG9R4N4BJMB7UsaqZeueJHcTje/FGQ9Dmc6QioV3cKcBVUkt8VPwp6gsl0+bDf
wErC8y2epxBQZCqTT4wyLOY3xOEw7zP3Ae45+genzCzemaUhKj9t0Cgpy3uV4hVy
mi4IZTs+B43oidFLKgV4mAHmRwh0cIdX2RZaI0y2GomC/BG92QJHwrdNNHt9C3No
mgFO1eznRoI3Vc6QRrtcaFe1W21OKRirkxBuQywTXaM9EPY6F6y4AItBaaBgFq5m
a7ZfrIu9tmOKBvrOSGp2MkJHo/QT5IZBkaZn7wHWksRcFnC5JMhwE3zkO1uWSSPv
KGsKCbxUCAEQAaTOo+/GK3wt//KwgiZq7zRT4+04cqAQPkRv7PBtaFGlfL3AyBUJ
B1g+5J5QMtG80WbGg7zhVEHiKYOpvq27sQ8qFGs2mBdLVDNbb4Yxk0x9Gc88Ro5D
`protect END_PROTECTED
