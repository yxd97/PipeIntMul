`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoBoRoDZfbCAfkGCvkMQ1GUTR/TccHAqVNog2rt+c8ea0BDcD0hZO7fivtoEEa1j
6hLixReLSicLSPgzNmEVppfJL0+AGuSKGhzEP0xjL1/1N/rgrgPBQ3QqrpyR1sFK
eqMpCo+MuXqy8dSNTJ2HPeCVsd3bWdvBQykSwRhT6+CwaUB4Vk9Jo8+kXtaVwY3t
4zJdwYtgeTJMpw3GJEqxQ+geZAtyv9IaRqQktGge87dtuuX59RKB8uKPGEx04KR7
Bvtmm9ylOIcxe6ifEN8tdI9VXG1PWiKX2G9c7xmrls/Jgdqn0cM70oswoftHMt+l
Snknl/NLHEKjieUc5gCPZygOEyRi2zD1HZ4Bj6LY+mbVDJqhZVsQvNARlBJSi6l7
9Z0R4B9VF06BS/uSZe1O9kVEjQ7oc7mKxKbGq5/fNE3NXg2enK4hth3zuRkU0hwX
`protect END_PROTECTED
