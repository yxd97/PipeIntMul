`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbKaWhneppykAxhnmAGRTPM2cjYxPOBbLSyfIV0+Q1fOFT8OsLknILYI5XCzofAO
N+x/8DAr/leEr7QFKrQi1rzXQAbviXK7ZmUmMjpj3hRCkJn9jhr6CnzcYs+ZOlA6
WRe2+Q1uf0VA6UxnUwic44jZzRop3WY1cBMddoDyF+0qoVXZ0yk9PbZPyHkEZOpc
XHjsmbvWuULXk4aLKMnQ6QQv4JeCVrrhiMvloqOjOs1lJTOkSc+nQ/remV5a6zQZ
fYp09/JwrsZggHijK7kjpmrEZi+xLWRWFIWr4NPI9slNikTtZcQJYiD32UBo8klY
3rxP4zrYpQys9JTX+70lvtRvcryf++j5rdQwSrJ5AGWmxUaxhEY3S+JpXXVY2+tb
7fV4v+9TKtZs7ZJXFPj7jLDKag4TlLS+N5aicoU6K8o=
`protect END_PROTECTED
