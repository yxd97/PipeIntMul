`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZfYnShHrNHE2ON1WWLZzqCjejqiELxDh2d9BvRqH/lYOVJ9aZ/On/LEcGvr6TRNr
Uua7aTg90FkhIimXZUSC6njzyCW6nDzCSCPi2FPgygxNiWZdCC9WLCVlozhKuIYf
sw5+tOIN8hmh5QpKMn7ECrlMAxf2LX8yK9coTZeMOuyemTMjvCPjb7Wu51pRzI29
24++eMmsoDELibJFWOaupNrR1RbYxRMTXfVoM6XYqiZ7+osGKV6sHgHdDH9rdq4W
d9lwQOSlhIznSCUgU2cutj2uXJv4P16nqJTE3MLt7SQMP14AwlSAKPIxQ8VUvrtR
6TiSsvE31vQEWgFkxlzZKC1JbuIlYep126OuiFHwDwHNvNswU9JV6JBeRYhtjDpN
LvbcyCNnDO3ZkK4rjxg/ya0If5VCDD44hJCZfJ9pty/aP7YSoZ2lrp4u5rRRShbG
/fEhvYcL3gyCCEeAqB4cXvu+O14/J4pnyIzwnFENGs3piHKmvVmjGRyhznwFnnCl
6hTLdctjrEkSgvw2lJXBuNxTeASgdu6Dsx55iQmL7PbaKqh+P3L1/gX2HRJ2Kmzu
kaCJh2vp+kFhPcNudw7lOovO5e4jJJxopymlpS1gfc/h3xXrVxPFtyWVIrIXimVg
kXcFCwo294ABVa4foRmWIqEAXm+DDuP0rDLtH3O7KMoY9GM5awYO9lONFM2n4nWT
ibwqBParqLszf40xAr6zvjIJywfMUunuAwboCJ+O9qtt01xh7BOUhCT097fnDjPK
Uo2OuT74eSz4hZ1LcRJppQ==
`protect END_PROTECTED
