`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NqvEFGlkugVcO4SnHsootOfxZzrTKELKa1lnCEWZhM0t+AQQbdAE+KNGg6wnzaxr
b6HsF6l5vxHLbVkuoPS6/0LoILugHWW1QwIwa07fx0Ni2Gxh0K7IR00I2oBpByJK
1g6qtPnNPI9Gkz2xgVYhxb2Jklm8sjN17itweCWHTtBZyJ+CZtYEhnQ0ZSh3cOke
zY/UCNxMG3wZa6bNRL/4s64parRt4lbQTx/CQoyhcA3k7TybnQPjmPpxsg0WZZwz
LUglY6mkFhi/sC+Hct0yRc+u76beKC2g6/S6WKrBG77IrtFoaIDvqyRNvdCxxlgV
HOQhk8BGz3eqM50oGqdQf5wTA/XanQaTFRp5p9hlHJH/XBjFN1yHS2UY0pA3Lian
5WNhpupXH5EmvQprQJYtZAluTpFDe/Atr3kzuqub8Ve1CwNlKKVskggtsaX2Ncju
cGdMBAr2r8EJWj1DL1aJH4bvzmLdmUYwM99cvykPWuzO++0aHDN85CNAL5ux1viV
7NA/8+UxvUM6L1vn/4+xdLkkwOsQh+2RWUEnckXcRZdC3BevwVj4E3ul3DXu02HU
0coKzIVXwhzoXG2pNYy2jSF70ARlBemcIySl+6AXodDImJic88y5sXD8xPWOgTrB
eZ0jDWX7kWNdRIZOhbWYbTc8SjNYNDRUX8Ud6FXgufBOsTz/2eXr8/wtjLy58dR8
HWKtIxucN6kFqOFaWd5M1CxaTdNjn6Rj2du5I1cyFfkomJOpsa/Y9viiYgCsP9Qk
pjouJc3bLb08M5dGF1W769qJ3Gn+2uG32ZMERPaVKhd1mbSFAGtP1Se/bwWSQ6p3
NwnauubYYZnzpr2esQH+jCRzEges+TLHVkyMnYgYbhNEU7DEcWQDv2kpKd9zoYjp
JHc//7XPXQdksU443YBc6/pkTa0qI9QSOpQvEwfrrK7IuMXpxB3HIFQvUx8z9kIw
csaMxFFVHtRQN6Y13dil8tYF9zE9Q4r9srCNd+CHso9dsgLgc4MZK39pkcf1B9Df
TsZp8c589OZ6DyZQ/PqPfy+WI4Ozs7psCYBWcAbQ0CBYqwbeiTxlgs7FDDwAZZbL
g4UHiGJSp+LrkNwoSho+tg2dsG4fzO8GRgFPnzZ3RaADLZO2zlDx7PODHiOP+RFd
Z0UXaJTEEy5h6x6EMANQD6nWF4lKBO8OVnM/YVqjREp0h8Qucp+qMOZokXlv1sOo
OEAfwMn9OcDRTqS6TvjZeH4Fyuzu2SJG+Q6wOxhHsAXR92AzCjqWMfbZiryFXFFf
5RPXS8D+FGECXq/XlXSy61JS5ywWJ9iLGhDzeT2UPq8T6uwocPCDBYmSbKC1NRTF
58Jw/rHf4PrdeYu5Ahy5XaS7WXaieGpalEIcnEQHgGBRe/XK9Jh40ObsaRmJiBWg
4f0r7Htw6p514V26wdW9kHLEGPV9p/KWpIcqLB3+p659TZDWxQG5ikpMWkwnP/Vo
0uYYavfQJce/kLpi+yt0uxMLo6vV5/OpQFvJZCkl4eQgreD9PnYWltLCxxzMWpB0
LRkJuAVy/dfx3bszRzZ/ytFjTNjP/ZO9td1YcY2nqgxD/1UX12OmL3tfDmDPGEfF
2Mr1QFg82XWUYDTnJXhv/09SV5Tqd6LD6QKceO8ngPy8atu9nPQoZuITcpvy0qTo
7S35zfWU8dhRY3kDvMBL7A==
`protect END_PROTECTED
