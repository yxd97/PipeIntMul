`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3J4J/dFSsUzysVWg2NqF1ZF/qwNuG7vmV+/qG/4Iklukps73Ly0LQN/CXCtUKMJr
cB0f05fc7BEzIlen7MgHsYFm0TVatq798cMdl7f1x6TS5VizEMDVO2NbXYFuqTCZ
5TbZqUwuXi8cH5HXT3QyxU1We+83gM9GTu9y7evWP8eRA40zriep5gv7oBZersql
fL7uYjdm/LMI7Ge85bgL1/TzFaU7+7rTOJDQrEG4NRXTBR3IuztBaNVc8TylUezq
3Z8R1tCCJMi0ZFg1di/7PqCYT0Oy3UOguEvNUoRKMHHCFdaSpQbyBPVZrYdkSi+d
U/YKrcqc84Ylpjc3oRJJrveTHSuyJhKQ/b/Isw24GujGOUUcjFs8AB2nEc0hJgeN
bGMGaOhtVwyxuP4YLFzFC3YorOyShZdINiY2o2O3OvWsNwQuEmQxeoeND38W6CgU
+uebuXOxAreqvnSM/oYbZKAuWUK5PMnd1cv3ezuOUzGZSnuft/bfp1rsGMdKOKBf
cYK3+a0FIIgGj5E9luh2OiGuMmv3eZZxfFK6adMjj/+SV6b9aym3zG7nmXBK3q72
J9VlkMBqcEAx8Gc1FXITxfbuUF4O7JZzHjCocLyH20inop+ozY/LcUAeZY2WYaWu
x1r04gpa56CYPumA2lJsRG2YY5AYZjlPFUOmBQNh181Ol9EHl7wjDYPQcJXRIX+s
CAVWtNHUIVwmH2Rku/jRL/7PlelxFZL6XvQPgboz2PmmnZvx9MX3Vo5OuiYRNcA5
t6udyTRXKFXNdpyCbtxw66BY4YWZyHfc0ICAgxnPM26flAs/G1ynLyXe6/5jfALk
Y1Cpf/xoWdPfKIC0RHnwHSeCPztUKbvHUc1dDxihmuNb0NFpx15pTSEfWGJ8r80b
lZAB71+LyCB1dlZD+y9S0Oo/BQ7EDNa8eyoZCQ1daRM1ciSvsS8CnLZsXFrz7txB
ZZ5aUrQMBkcFvhk6er0zJDVku/NfTG/QTb3X5+hXSgzIy+oxYOp6TORmgMRRCcJw
VrHw3/hrLmqTCcd5EqDdzGPeMlPXoRq1xZnE2faa65CfPpf1LX0Gwg7I0f33Mbvb
kxvimipAvQhU+o7YMPF1GQV0Ug1aiTXEH1cFYW30h6pK8Vsoc+Z0JePzpU/7D5SE
mY++oTaYeNFqjZzcABKPKM4Z+uvb60E7OnlyjpCW8FNpzp4zroEdIXUQxF4p19UY
zZKW4iVM9Oa6hlrSUbehPv5W/w8tLh9MbY790CrbKnZ1VILIvhjhMLagr+o2OZ47
uKUWTT5svUv3O3PCghevzP0P8dmglar0+ilK/uqGdCBhDpUJ3Fdk5EIBm90sANf2
UOYmMWN2TsfVmCfGOFwNCguhX0pihRS7RXmWhnVYcdU1KpJB1urdNroLh/J3VOwG
Pe39gUVz18JKm3wXgt8GaEjuvYf+z4hFe5g9hF/cRiY/MLcV0n5KDaraWq9hwdMw
NQwotCAtJnYmaQoiWscysFxR5LI885tUMyrOMFoShluuy2Ml2S1LB1ZRcHllvMBK
X9GVxkCQqoAuIhyfF1T0/9wCUEAU8pb0oE2ColGdROc9GAfTGcqwn66ai5TaOOe3
NGFP0xl04yWeKef8RbJO1NoGpy43oO2bHXmXHOheDiKm2QFYHQ9A8pu67NBTSodV
e/8LOJEI5TfYsja+cOVVGLn42qUrfHUPSaAsNeK3L27lcHo5PjIOEcAqG+8RjlXg
GQaZWCSOHznvZJS4TgILlAZb2njtDanI1/JmzUfcbqTUaNm5dsCI6tzcCIPB4pDa
d9Zbpiy2GtIV2DueWBAw3wTdUkQBcNvjeg3u1svgQJngwc0D3DqudtQ2eL6f+mEV
tUKvO7ht/GpLCyIjZ4IrPB3vA2OR3/QfYvqoNAmViSRwsDzyoJnmcBaqID+CdDV3
N49BWpYrlAAS8hqMuH7295+SsTr16r6051PsUIN6Jn1ihulHNNCW1J0RdJvKd+KI
rD6v+1VtYMMaZKMcsNH4nEjDE+K89b9vhZONib0FJqiNeV/grVpH8o+Qcno6lgLW
r/JCL10Sh8GLwzXSVRWHmt74YsErmUdYHyyL7Ltaax8JmHSahOlTSz+nfEiRaa3d
aWTgW939tSE3AjywV7rXmYVHmbjmTAtdkNpexGn7hG/FwXj7embxnmOoqXURaIJV
3G+M8koKHwYg05VXehe5AYeaTaE3K8G08hbFyqrdX+ozHHEvUEDxZ6kZgsA5j6rx
51jaAzckECu8GW+f+PVuyUcKUfTGBKyAGvIZoRdf2Z7pGCZNUJMOnQIqjyHZ1Xyr
7yOfM9ndwTR3P5R0BqGmvfDD33kTtNK8wf+gdKPlv6EfG2cwFB7PZYa2aE+ci89y
h4mi5M8boxLxR7/5FY3SWBSZLIgIQ0/6zwpIRDe/Puy7KG5WBk4JHJ/dsNIHSch8
tJPdCkJnTWYetJ4cAP9C9bVjPmpjjzpyl58NqLWSpc/AGVA0q2ZWUaykSh5mSVRm
2FVMBYF3+wewP/ZDyCyuhe5ecLgjswJC9alAmT/QGwCPDxXnk/EZCMJgsSUg5nZD
6fdQoBWijjkrlxmUy7oRouMLM5LySXHZE2qekuQ3pOSpwp0fzEzSp4J4PegtZEcD
fnl6kAsaMvfMJAk3mbeemRCLZKnW162GwwU2iAnZfU5zDh18cOG6++QQV1pcJ9kX
xiyh11ywg1NjYfoFq5OAJE94quZ0CYjbFeW4Om9+NAzKhiffTF6ZUn7LczeJ5lTm
YisBbk/GXuQ1pwfMXch4tA3ivW1WA8OGt2mKMcdia42WWk+80IhYEiNdS80l8f5O
yfDqpEkBEXmRZAD4rZZ7Pbwf1s1sc6p6V4ntw+8KCGBdziBpXAUj571wttoiB9KF
u5hsrLAymAfTa75L5YRaEWqBWQHEZcBkFhNl9TAAZnKF16vD52oTxi7sHOJCv2JD
QGw2RLmLPBnJqzXx8FF5VzIWhcZ0dKNG2ee1VR0x+Ffj61CX7FlEsLqLN/TRX9MD
Y4nFu1qDcTI2hwUtpGUvawZYB/GjFp/laB32hAAia0hxxnSN3S68v+klXJyZcl0U
eSuVnbzdlylDKH01FAL9XUt0tcUZN71e9Ci0F9OyLbgU8jAh4WCVFgBsqGHSC8c4
3/1gBfaMZzzs9lBXqZ0JH/bfopsobEtllvb3NoBFlIWwDNEk+aGB7oqYRKiopE4Z
BCqVwL7JhO3MEOLwXZlfurB/nHTohf0iE/k2VAdnYQqftvauvIfaEk65NNK5thkg
88GjuI82cd4kX3vNLKKYCl2ex3VuPAAKYYgXfir8mIJb40yZ+HSXm5m4dc7jurY+
aIoqU3j6VyJvUrpbOx+/ogAzojMl8Cr3XCsiE9oN0jx2y8jurpi88KpsGJsQl1WZ
wDT9iENJgXPW0CgEJBis3qqwRbUMh0bKtk/R2wGGEh14oSVG11Y7xQV0Yysy42Rx
5HATQCnKD1GQSVzwfbhG9dwewKJrDI8BsEGKFnWcfT1GjrHU4eW141h0KYsbvGu1
ZYtV60ClpnKlnW+rUUup/hPZGeN3Hqpvoo7OZcadMvFgwy3W7/3bnLbF4Xi0ENjl
QVKGVRIwzIMc2iwFO+2T3fjFJ3eJ/jy5+V3b3tqXzHLc4oU/zI0Jdv56W7PpyTh5
RqWQT/OB6uEPvvOFpoArauatRLjmMNX9S+EwJXRtyBNLy0SURo2H20hjBOkG1B38
GCH8us8wQyCpYiYwIcUWHWrBCOOMJwV8jXcMWqXsI/3/W5vbTNP6Xz8jzVktbFuc
magJ2rLfa07LWD/uKApuU/ZHRUnR0kUmeiQ76dJLyUPpuZBH2VOCvdqOcrk7BNbz
T/jOltcdajvfb35ddGZC+8Kjg3kbvnPegjNyOL/DebznVxXbZpwslUukxE1uhsYb
j7KBD13tV1TvxGnetmbEbQlns/6M7JgJ88jgXB9oJs22jYIwRFGK/nxIgZqFZHr0
SPp8w8ONVyd6DIt73UNBUyhEzvufGCibCfyQoA6NGK0DVQ8DlnHsvnmRY3DlDe8f
7x4jI2FvCugGww4TKKeHwFBTcJt9MQvlNK/8wZkL3XetHacriPUyvj+lNY5iT9Pr
8N4hITwFCh2GgY707e3yZO9uSwohVIy8htWkQ3IbTHPokHuQNzytqzWVSRqrtx0j
lsPhb5gt6FdGvyhcNTS3HSjWSzgSgUR64Ppk1AMlOESzZpZ4wX5FWO3Is6dYnvnf
wWiSrqWJ5/vtB7ikwPiJj5dcR7p7t9EmeiaPK8xOIbK6Or8M0hH5UVH+8s/+wJmr
6XIhJWHmnLChTl3pofM7B43orbDi5TIlernINHt/0yLBUxuFVybdO/O5uPCrx/Zq
rnLYkIcMHn8cN1Z5+lfK5oqdQJwL4msWbUwv7RMaR/GXhLCRw+Tx/41kGTtkIXjH
OAxLl3PrJo/PRcyJxAE28zsNnyjHi34G0RwPb9JFO2KIAYUPEX3aPNqB8BE1KXmM
IELTHbDvdOoo+xRJDmQSNiIqSx2zQ389sUvAkYTILskwscFfML5zpmNmPkahex64
8mHJtoNlds0YuezSrsq4VInAQyiiwJNRYqReCOwoQLHRE6kcVv9P0fhpBqMXl1m7
2Ytfb4H7/88lxI2rXUezXnZzFtPxep44StaB2cNwJCJgdqn96qIgChTVxFCNcpiA
iVz6kT80kbhkSEkbil+uWPBg96uUCPs1GdzsJdKC7lg7YUuOVW3uTU8aiL25Rpmu
a3c//ZOBJI7035e1YHzFmy4kV/FJ9h9SckA1dGt/VahbULa6Vg1wOH3hgiHBYAe7
BJ2Cklbvd0W1bffBouAhoiOdgmDXEtiLcQ6fIDh4z3vgSUpmeL89IKVZhpej+4vt
b+p/NH2KmBYRt2PyhCqBRDKouehic55MWIGU6IK5t3al81RHgRdAmwbv4waBPnnr
7VyuOEBm0VpkYURjPBBaYHT/QGpGOxdCUMvFCe8eYfa420LtzgaQsbfAFt591k3I
jDIkHe14Lb4VaSKqnwIkI4GFez6W5fmlbvNV+X8J9PgaYciOBvgnUWeLvoOeT7O7
uReohuAPa/C+KF95m4hhdpE3RT+QQIId53cVP4siyuQmxZua9pcGgivHfj6ZwxJS
eOZdcTU00yEgCv4/bqp336xWIZrVoMzzwXclSgLInUNMQizo8dR6sATG2bt5FrGP
se3B66cXmZ97x97kwISpC5JDzNLBBEpR5FQi6BiyMxlGUswq6rLs3D/vd9j/b6+8
x8uOi25x2YLHfmboVjY+j6asyLt1zFw+6YKuZwwZJ33IUybwc0UKQi1eLteP+q0D
09NX+Y4AS5GM83gbP5i64slUNsO0kRjsJz2Gy/iByBxg4XfOTNsqOqtStWWTvl6l
RiAYp44HD1O0lrnBKDjKeAOuBAYixs/Q3lfmKrFp4/gEcWTS2n9gjWcWp+M8j0C/
y0+6cvFsCdZFGqxk/c3QeckiX37iEAXs4IR4Vz9w2XcRo1rett5+YZLams66/+Un
xvGI6Xfu7KkhXG5m7aClhtZ2BYEfe1gQ+yPWw5AVCcpJjuQOQHRvkNCFhit/gjrI
T64hopZbyOZ9mJYVN0WCSrZAn6YyhaZgJoxyHYgFu1HOhyyTx4S6Pi8+9T22GF4v
FvKwy1N4RGrWTlKGLiQeKOv6XHHo8uJcpJ9PxagvcpNGymUvK868mktGi5bgMlhx
p5a+rRN+uMaiE9kGofPUhsZTvw1C4B7IWGsoK31dBglq3S8I4AknwTRhD3jHP4q7
lQovOefyJdK7BRUtBhQSGKDbuLks1TBVmc1uDZS018winJi/C05YGxSgy/SfcI+C
M5ozuJL994WuWIb1sQF3GPGkGxFWNrhS7ioi5ogavOuA1WTM4MG3ZimQhYbwuW3j
46yLMH/K5Nn7zzRGOUhWE9phlHpqOdm8sr0bQQywejJuzixPtID+Go7NbLkbRyGe
yD+lbjO6d7ANWTEE9sUerB6n+QuXbZ0rEwskrd8FsA0jFTXE2RyCsUT/fJ6miVmn
wDAS2erDx6sKjj7BBwi9z5UfaiLaPmBskclsrifSAeJR2tkyWi3J/QAimyXPzorb
ELnFC5moMM9BV+iiEbSATNj7ycZVKQlwbLfbBfOMWSJk/XjW+BS4eRtWb3YXG/kK
SotmDFfUHGX3vqwCkW7vEzW9yDk6239Om+1OmbUE3TyMo6Txuf6zERd+4vDIpBB/
caVh3QZBfpxxSE6das108JArdWVDFhRftPu0qpJXMgRa+V9m/dAzkHoeRLapRxQo
Hx0wsr+HGXZMoBwIaJlKFugZlr3enfCdgrQuzk8pQNdW1b70Jfa4i5pSD8wK6lcf
H2pLzKO6idDQT2S6lImIJ58N9it9FU+7OJ9Ia/blaNJPqN6X8SZixVs7l0LpSQFO
mOcLP8k6DYVbk255uj0M0tzh6DTftM4otiMxTfPBLCi23KE3Wke8uh4XwxKXv1Hv
i2i7Aqlipj1nFRI5F5OFABfmLYyD8bvdzsM3Y60Y4u+RbGuJl+krxyKAl2x7DuHv
vLvASXM1wJ0BSnJmDe1/TNlR9zUNbkr+KpyA31RBNC7pl0FaO/jfyvgijb7QcqsB
K8ePohr51W8CgbjP0H76TeJ6p6arAhLcc/J4F/dq8a/wBVOnryxCcR/9xQSX6HZM
lk9X+HYw7cP1Q/LF+JfpbPxLUrs8ulQHH0386s5htaOxiYyUVarP52p/OVs8aLJW
zpXDz9QlK/T6CVnpMQDpB6S5bz0lUdN+5ptZHMu0PXCONX25q4By1Y3xmyMPfCwa
THVM6PftflXPSa1BaFbr+hmV8MnJHlxx7X1CSdBE3nLG+HHFdakg77bPleSUzn19
y9MrB6Cn6z8GExoA8M5BBDIFMwQidG+ngXz9Rs10hc4tM61VE/cPUyM1zkmDtAa+
1DP2zXBjy48aLsg2oxss7GMc8sIQ03inUe6tAgVKi47PhTUCoaGpKiE0qDAZZ6gV
Fef8AsmqaOl0PWlLhKfk0cP76k4WIw4820S8JqMSMNQtAJNOtA1ZOOlr1gH8ITDg
4re0HrXRs2Q6eCvHlruApBZ5MKrRoJAkVLfa6hkOH2TactQ4lZ70pbR76N+WJo7e
R+Jznb0yyQcfVIXxk2mL+Rd5g1KzKi2PQoB1yuJrdio1nXQKzryyZ12xTxQ60rAf
xB554K8LmjsFLOdCneCIoUi1mju3qgk8kTAFFyhfp/9uHXj2ANFE21DvprWUE2uG
Pu6oMIYPQ4BAmF6rnePy48n+BF8dSpE+hvGxSGZwJmDFPe8TZ1WhAmGml8Vhjz5e
JSCTtmGMVY/ERvIFALGUdMerViGaZ01dunsUUiJmVMQ5mVcHguAKpNw/mLBGaqsJ
5wlspMLocsPWep816FIg7lDryGAjsmQUCLNXkGic4Sja7nTY0sb1dSv0xr6xbe2v
DYWIWX8qHAw5B7622VgXoRaJyomZje33WDZ9GQ/u3R7KvDMypDYPJIGSXTI7pilX
Vu9L+hTYCzACw2OCgW8hC0uuRrEMAiFMYF7ktFB33b7BHEK58keOY1HGkbgJAv2u
Z6aeE9BFS27j7OvGAqCbeTRSwRV2v9ZexzguXuYoR3FB85Mk2zP3+Wqiuc0FRU8n
Easu+5Yq8n541RDAzKwDZgEL8z3NbEs/cPdKMyuSZJ18IRuh4vgd7eMpofOD++aq
YGSmERjd5Ng2H3a2uiqGpsmb54bgwzNLwI8rzdrtozooaYrXZwGCFwxjjwuhhSns
A0tAzwWjZ8wI3B+cv/++Nbbi76AA+HwEyqwsOlY/uMzodNvcA0MEXUpvjfIVn8DM
paA05FRH6tg/WBWFulz4pH4xAlt2p7T4pQnQ1ZzHIPadYVpnUUFcSRgYJNvipBbx
CT2sAQy2Qsr31mEQIE4C0kDzy0NCVMeEQfU5V2kWhzSqxPd6dQAf4arCBKDsfNhW
6mioWLqvqC8VDLJw8DtH+iBCaFZO2I0MbMM8gg/DxY5EvPp7TUwz/Lr3tsKHOswz
NVFEUEY9sbJxtCWqBkyOpMhRSHcbP5fr/1rRf/3ZCxaqNReCe57uCR9PNBIE9uPn
6lVNAkTdqguphdUWyvUNf63THLqdAdPArn3F3N+3gXoyIyVSNYS3z5QHV7FMnODr
3p469d6v5igNScWYm2afNURyFR3VfH+2eKneh8RU8vJSSmgLqSNXVeVDL+RloEes
yoQTO8mf2cyU4sqSkJysW0QdIsG0to3wVqarK08AcS8WOrvCoIyFYmrKjVaY5Lei
ZI/EiQyhbIJdasVKwafEZ8sRCdgU7ESM93c+mw57+kGz2pmtlcL4whoNETNrXWSG
yj7/5/OSlEqRFLlLPPiVMuSDnQx5wbS6tC5KH6+Ow5ZZYEPojun1rJogi/3Y2Bx6
VXW0pIu65Hdv4vZ6KUrJWUrTmMVRiiKmS7LJFH1X6JYMJN8bXqlxOBg9mhwvMqAn
+idujIsstWc5GXiODm0aJdoWUmMYxrjPP0/FUT5Ex+DjDao/Z4jccOtkskDF7IpK
/runJtYoOrm1jTKis9pejnSpLXQCbC/xMlcCnTL6DcfayYUfN8RQpe7h5gI1oRKR
cCP+Xay1XxDv7IalwqGd0H1PtC5xUw20yBUjtNdRUBwlYsOFPCDgGI+ZwXeglP+2
gG51NZuJqYDsz03my5FCbFdRZMWC82+0zU+NKyKDOLCapJCSiVYFCOb9PrWgLN0A
tV6K4QhtB1YYc+E1KpXCBHeotMbY6PWVB3VuP0DLaLyWWaAXRuPbJilVOKoAF5EH
mkxjYUj7QPSiA0N5wqI1qeYZWp/kJT6P2j70pbhzrcTkXeSz7vxYj+Ml105qAIfH
qF6r8RCUzm+ad164CZ6JX8WdzAilJ9QyJqoFT9sfe87IC6wOjN8+ercJv37vS7gU
KBmfIBr7yWMWpNb7YTBa8i0NAEcFwjk5UJPxXgo2idNuFc8hMj3ksuvNj4fum1t+
MmjFVQ/lprO9+Rmzl3RoIASOvi2AmGaqkFqQazxpuNwLoisyTYw+iOuxYJ8fbx76
3YbHHUqkow7laiEr6GZbR1lu8YNJPsZmwzCXPNe/F9l5BCnDBd1pblQhLvH3lfS+
sNTCWTkW5fk1yv4Jz4gkWisr+SYQB1COaZ99/clWdH6RA991jG7R955W1bpgttRi
wMIO6uvLy38HPgZz1D8+Sw3W+77HRZG0Vr5XNVNxBo7GKv6bvXXF3+vgLshCQb59
b/F+7LV3pALqK0sgRVSoIVSc3haKj0/THL3mQWtud4EmUB4bh//Te6aklmloO+sQ
c8rEx3/Fm+kMJ/z3/FiG6kTJyvDU+g/OSkfsoEypoY5W17leEjEaBaL+gTfnHlyc
OBdlA8eqERFTyADHWePFgjBDSFEf0JL3vxV2zzYKflQITTMhiaHZYerdUiSPr/0C
r3S+f0YXLe3HeGxrlRGANR0IPlPmWRAFLPLzRRbtdF2AMLQ6jrV+xWBsWGvUXphc
ZwvGZtCykowdqeDiyBUKQQlcMSHyC3ZdQ849nLzYairI2e2QPODgclChGU4yuF66
rjUP0abATDxLzKVCI5KU1NJwutLgO2E/jkzFEWM0zXb5GT+8dDemyuMZkN7l1rrW
Acgi/i+gC0yrlGSaH7QY4sIx1DW5PP4m2/5g+OgDysOFOtpMDA8dXVlYzYNIUGyh
z2fiH3oVMKJagEyM2Ax6XdJKhH4Qsik3XRF3rQSsEV+K6whbq7Fo0fLt3onhA63S
rVPHkMerhN26HemAUVhaMbVfnZCeM0sxbdcAiFCiZyGIP3KoZnSd+APsaY5Z6FE+
ua8uvIOaoytoMfKE2IHKdqNj/HeRe1Wl27BF6aeAc7plQzp+LO6RaN4pHwYNRD+3
kEITIFn1CMhED+bt3IhJsqigumyoZ8ibFLXI4LpYDxxcTJr4Gn/wXBQurbGF+tq9
Syo2TFDTQGScP2I7Fi13EFiyPeobumAbg5EbDsMjZTel9Uyu44JG58F6c5Z1wWPN
V6J3f1l6v60Q842aFVS9Rfj4Bb8bJO378LtF4y2V759E26iscCsqQ7K/0WCKWxTu
oqv97hdFKfa0P8IW5fa4mFgeJdDapvogqb6cweE5G90p4dVwGYbJty76f/W7ZWme
W9VGdkbqjJDUioQNBZf3OwRl+1MpbOeIryW3kQ5lUpRCpKfdvkANAK71BoMmX92Q
XrJs1vp8RLCYW+63pplm26SePZuTdHq/G8kJARWqWq04k1HXewwc51twZHpJIh9u
8GNoCGOoZ/1UVwnMCgT8HW00jpgEOACXATE1yRbCzqQGBFHver3tlO4LB0zDM4J8
F86ghvcCu7OsnFg83agidc/PDpdCR2H0l+HA9xKDsr7W9OjS6c3NQ6GbxCBdjwXL
3XuC5iBPg9daq3pAadLup8qjdgSCI4SiPGQD3BWWWBWzvtbPrP1mHxvzrHdW/yj6
AXH7K7k1DIgMwVqREpXB+KxXHkJrfIYyUBPPJ9R94HhiCo0A2hJIpZVUInoHVwAY
LMVgRX5opMcg22rd4ssvSplNJjEfD8SPJBFVOxhEwPG5oZcouJTKkFWLAq4VVkbN
gJUg7PdEJPpQpFz9SEgCvvI7tEh7MvPiXKp/e5dwUlODDxWv0C80Csqn7Qii0Gg+
TK01vlNZeFicyMrPD+2SFrSSjqHoExkxZQ+iBBZN3YRxDawaxzwsXnKNWrvoaQ/9
TcDZEh2bPnL6/sl3AS8qTBYls0TC362DWBwNGShnuzOPgx3i1+7d2QcegXNteD9s
BBdE+UrKe1hAlXFQhHvmmY/AaYvEb2knjkFg3pavR1mEinMiLs6yWYqC9i0Thgbh
wFRciop4F5x/wHBMJrJaWklEE38JoxIw/0AKy57HJ3asv11arUp/xzPfzEmOldzO
a3DhHWFJ36OkskKiykBmkbf/qhjnDj0ATQ1GUcz4m806ayHHCBZ/bADFTBCcitIm
nuQ/HcMps5oF8oVVelIF8Tw0ABAQYil7jSbOOuwCI3/0FVJGMzt5nSmKo1IKjElD
6g73jKNjZ/9V/edBPXcNiZvOt9LY1zdP/WSS7KEreAwTgtn9t0ULXpdemWmYB6wN
KaVEyPxsG5P3BW/Uv8FHxB0hTG2dhsDVb1ms+/mAPqF5yP6fZc3zxIbOmY4n/UTI
lL3eW1uorETI9ONeV6K0mq1gACuqhSscV3Q5WbUk1P90X6a1WdsbyPHHLQqo3pDX
gBumKqjQflTLiAxvv7Bzk6UkUpM/gLbScw3LIHWNtjQUqxBxqPbMg+jtSQQtiSDJ
/QyTi1r566c1x+8Df/2nDYlyJuKXE2xKT9PogqXLVnT8F29GUuUcT75dB9OzSuYH
1QKWTi2hQt20bXS9joqTVjfAQTcw2J9ISYtSrTG0VLUixOM/73D6vqkWL5PD3mmu
Lo94/O68igMSu/EAkKskIEGg9n2A2rj/AxTKfN4gR5nnF5BdCbKVJhnRVtuNdij1
FISfz1S21DNMbh9AHZrbxIOqgXs0+t02tI2UA1PrWNddlYuKwDlRGTZ54VH/WzhZ
xJcnkOyGxvGUB9X7il1OZdc8XNQYMrOtcYGMwDJKfXF7g1T4R3+B16uVqOdsix2i
eawCJytcchg/lZL9Irf73qpdDK9/XcTtgBgzenz4aQDpX2fqFZWCMoGSMVI5kf8d
H+sTTCbxWqAm4OBi8AfSybA++aa0lrmncaNPAznMi5T4bwYskIE71Qdui/0WFdYK
R0TWFYgHDWQmbmqnPEsCbol8vUv72wDAb2+Kt6j7VBeyx7yj4g/FgZ0tJgpgPE5O
EU6FbJH+PGsgysKVl+oUBd/ojG4jZgtwJPX9QvHIKCTIWqPp+THusUKJkYmdFh1t
lj4L2EOtopOwgmVflDyip9lI9NA7jFYVAC+GLDgxq2KLq+B7d1hKaSWdM4vnuyXf
suA9U4/5IQLeN68RCmBxKeyIOCufEeQ031FA58r2+aawRjjTj3c0/hss+Jk0h37E
uyrmyeOE/xZYOS5z2847DcH0LHWkCTnl/913St5GG1WPdo9ymDPtczGK/abtjHNN
lYWN1UTFTfd4ZsMMkYDWH5KXzOOyvoeBCri59s37WEqrY6G8pyOuE3cRhzTC+4uG
T6CzFaSIHOnyZH9gZJK4Re9gQt4tsubB421J35tV92n7F96Njh1Kl4FiWnzeaNFw
nsqa2n9dTqccbqn1ZkJXcDo2n6IaaGMmHobIw1jYTGX5MGKOQuVCOVke5GcE/bj2
Lp7AwvhrJQUYC+yugrTbp4tXsuex6hMKHSwBiIZtDjG7jOOHZ9GAKPIX3sJzI1FY
TDlfFpTIUrcVcXBiMF71r4V9ImopB2Tlp9nMD6Ndd/a2cjZjtu1r8PEh92lFKlXA
q5KuhP6+UkLZH39Ry9iZFrDyO6bpR47AFtz/tZW44J3kTLwj6qMWhov+PE0mPP70
8gUV/Gdku4qv5CNMeOvboZWJSA6iAfOTsTduR66Xil5qhachrN+J55sp2fnbnB7x
kuHBjUtbiGEIhBUYB61YBKSByUEYuy78ra9VRm1L7opvjG90CLSXkhUpPWNcpU/Q
YR+8aG6hEOsgf4xBTha2C2rWnEwZmj14SdJKrRvVYKy4KolJZfsZ6e7BK//I62W/
pT3MzgNZROMSxTdQJ6HdODCWdZYcTK2tvTvbO7kR1+2wbTI9FFStdFm4Jo3YPSPm
pBQrfU36lA5FSAJFnT0xYC4Lw1PvEYy49DSgNuCvbFJA6EQWt2JftfZXjHlTcCsq
LzxjQSKz1q75sCbRlpjc1ROkdhqYrA4yvKbRZZR/S6JSg3pfgm1GUTjocTM2Thtx
OezpOQq1SvkF2Ph9DAgO5td9+HuhbdnYfqIA+vTSPgNJKYaC/36hatDDk4ICVr30
k6eCZRUR25jMitgrIqwDtL4EA3p3cBVfbUksIQDnDaNrgCq7gL5JW8ncYM/Vm3Vo
UZMm/ujGYer6x/iC+BWQn7yHWujx23G27YsmsXKoUefa3eOXfObIcoeu0DhNOIrE
YPl6HWR0k4bx4wBNn86eStr0Z9tH+Nt93tl8irEpifaUoNscrNp0Mdb0LRd3ruGJ
tJJrDtu/+wdUttZBqCOZzFeG2gu5LsXLMWUr/Lekrt1DjzhM4QvK2lk56bNl9vMz
Uu7ZuPTqO+arAwSseKuJ/VWlaSkeZmEinQz4doM9b+jfig0HtpWw5ECEePMw1I1M
2fwavnqBWv0Y1oF0tR27vaX96X4JZQs69vhrNfScF6BHcwIbI2Wo8ie6hc3qtOJg
ofkzaG70CM/xjzf6tUu5nC34IZ4ji+cGPvSOFgrxTyPUl/ezofG0Cv4opm6KGvhS
RXzR7V+qF7paQ/1yY90srbTl3BFiHhYzC4gK9wzwlB5cS0tGZk1yyQAnpwD2EdZs
qU4bU+GA5PaI1wqg3824NsSJ70QMpO5eKtfK18+1ccva3zdkR5ugpfZxVdwrMHEA
LZaKn+uH0efEBasdVmnCKaVvJG2GgzHfN3KXO7IZ9e7H9Wp6xVQUH8qxDB600gXO
3IpRr5SXxDn0eFg/bd86FELNMB9XnmGiMJpfi0JbmsGCaEWEDzODj1IMvDnmXnRj
fAg5j2XnfvteqGtXHOI9qIyBRxXJf0Qh7/dJzSZ/xA7YBB46s9CqFhTMaA8ljxhm
42zKcPY/nOz6a3frlDakWTm3kbtoJ3j907Q3lNVsiNOOFT4jdmNllDBwYNZSSPOb
qdv0GK0AXVrQyPFVqcUzg59Nw4EemsW8i+5aT1epod89DUvUofK9jO69IxojLBMa
JvddUEvrX1n+wpx1VXbUMlpE6e5XjRdZ1COf1Va247Rt5NG5w7mzu6Zyd9nkXIub
GhmismKq0vpYErGl2UHXY/KURys26CfQeVu/vrqw5vDehG87fomwF8UTdI1Ti4Fj
zPvW/0rQrmpCzG1Ttrc+OUKkT6Njq6ccYkoY6AIxlOmejRRweHRfksxo9YSHONoQ
Cu3ZZoslDDo4HGDnml4+MNYTpzg5dRea1fWocmHwi9V96iJWz850xGcgejrQpqS0
w/6DOKubT7XSWdQmWyXxewFIxBGTm7MJ7B+/d1khCChEWu0480XL54otaFOlRWNN
uJBta7Nj167MbqerGpvcJoGXoSB/0lya+MZaoJfGYORH2uCi2cK/a1dCb7LmNOiD
C/4J6Y0aRNRj5z4TGRvzDWY4iz3AAZ55qRrqfLrRAMc4D/1KIuuEAhlKq1oSGjRV
1wDa5rDOLMcfLiJNZM1LGB+jPncBCzKQ6oASRt/5DGJvoWaq42Sjc/7/dY4+Vzlk
WwH9+MHmgAvT1e0rdUyroYxN95JG7dzVTULcypKsAk51wFCrQa7i/UpIeo3Xs53X
3nTZacCS3zYXYMU6SYS09IhxnvtCsWDiwm92PO59JYghtX6yGB4QtGzoo5x1T4jU
Rc7tA3ufipa2ZGpE7/jSFEA8t9KOWbo3Qy9oQzZ1r0g85C+0dOqOaIUnDOEf8bg4
zjdxiBVJzj884fm05FR7E1mGMcYQ6DA0AidHzfMfwqhA6jUcN2YcWLlIedo0FbRw
63EjdfqUlO42q+flFYepOeZ42RDNcO9JULa+ZBLB+mUytVL0YsZ8GXvFlv72mwN+
srpDGdCvR1U10EtvZIljx+wICGW0Ys0OURAJ32HruMabDfQy0uc6rpQvqcIuz2JB
4xtQbSmsZquDWSlGrgElVCd+3nZ7MpF+806pM2YdX44n8dg0tA3C7rien2Vzc/Zi
y3F2Ew4X876YMuDA7MVw9XEiaGY86OHilGozA8xdayAF8kMsutlpDfOUIVjbWdrG
Q6U55lF5n3FJwsJqY5algrH8ewixJfrAdrFeVEDbWJ0JKeRHBwoa9eSX+fxK0gGF
807KzRQ8i+v5cG4k0GOL6Z852iyqs2CLh7jac/XU5RxbQppOceD6TNChguf5agiz
s7J/Y5lqDPW/yHQePPahgnGrrKTZLUFm8p0S6mhmXJR75OxCX3tDqNJUKAVlTxnC
zCDecv23IPBcg08558cjZr/r1DmPn/J9Ad3HOydQqS5PbB/9m54HaUWaWinUQccJ
UnuN+Rxo40ZGKJSRgCHkPE+c3fWWx1p2M3suzbBooaUmc9B8xzh6u4yzMSMRH6xa
D9jXaywkDz50tOxfalh4xrSqbtAUCd7+d+8BsmbP50PagDO/u16rgfBHajbDsGjA
MHx8O9u/QgzUbiJUx4KTYb2l2U5vm6vJAxVkKIKSDvah5ZryEFEXorp1tKoKM6dC
kyGJNr8jg71HOw0IsLknihzx38qpKLQ8FjoTwYz+gNLdz+jZ0LAs3tGxqG/cGqKX
Q5Tbb05gqNZf1oUvC9WyuVqqahw7V4j3B21gRJzzx0+ujP6e24jYwc69PMqDgOXc
wakxuMwqY0lxc71O7/GLyop6MYPPyU71+HReso7Io3htdX1OS9h3gH6FGYnf6seC
GP4piiYV6iysGG2AgMlEgrZ0DCPuYlRd3HK3l0kMcPXNYp+T21gZUp1kjRFfAiHa
eFZmdEqmklsh0BzqQ3O2UzywXJQuQfVbVH2+dTNKc9We2wOfVQ43131PQ2dEZtL1
le0Ez92gCNGuXte3u6rSqssdrWO3zkGUu6wdgIoCK4Yo8cAhmas9BPHy2ICb9t1i
aSFbcsQwHxPdJe8qEAHYmwWCXl7ZPbxKGZCqrCYdKmhMGkR4re+26i78gXLO9rPL
QyhW4b0glU98zmWhN97DYua3EmEweLXmB5cYh1vAd1NIMfwvGS+by/rO3MhNBEFw
mPIisBXl4pQSe1Z4rIaHzJLAtoDBFfFPtANdREF9j/v1mLgSx8XnY95pFxXZYl4e
n5QbvrbugcESrqwLR7XiqllMU54CtpE9F1Oo6YGRdwOTXRRz3hnzezDC4UkchqC2
dPwpq3mlwyhcz32V+hbjtu9mbnM4SaB/B0VC4MBinu1Ga+wsoBxSNijqO2Sc+RKb
elX5FizjkcU8eWT6IyLvAOYLZaHj6NDrrxcmpnAsiVNDo97JVwKkxLFm3GK5X853
4zB9O1vtKC1kRGxHr5AGYWjK/5IcRwGVzOzlcUBUjKpHMbhZ9CXKz6hcosRyN+EY
i8iyfXyWmWWoHD5VkQJUFqxA5owuNFXcmOsVf2/+RIR60C40nLzBEDvjvVhPq/s/
CAE3/VxAPS6GJQjHckHK1QNtn+y2NHeBKSJqb9U7Sy5KF16FIqkcEXvBmiRmijGg
wpgpRz/MAe3+W7GD5wyMjrVRD79dzrWpZlxxvOymPM3p4djitLE05nEfZI6tYWiq
K2cf1EC8PFI0MXzM7GOq00KBah2Da8kagOwG8wgG4KyhIYXX/Da7tdPptGDIfx3+
NKmItLL0V2ecPd3KZ04RX9bqF8ODwHQga8Aw+nIS9aS5qMa9qHGdT4soEGp7UPTx
aDh8eOwh/pWm0rzQAFHbeQu24avJduqO90lkaJAiHlMHtf+Uto4g+9a/NfJP+Y6C
9RpyPqmSmtni0ySWtxI99e5q4usEfzFXOTinr5G1HWfvEjQ6jDobmi5b6vH8WOae
cgPaKKHWtFd05go4tyruLHwrbgdisDmAm9Uc6TPebcuzEzA807t2C2pJD2jKYuRh
ohpgHKv5IghnE3ZcgQ5hErKHLBZ+tuG27hcuqtET07YTbruBnXOrPXH+CcWu9ph6
haZHMldQATpivq9U9n1N+k4MW+mzoHIDQHpS2Xs8MMUQnr7zvSmt/7jdERqmFA7P
4dCKPw79kPRr1oOBSr1iEwW6SKg7hUXs/wPmt5juiFBkofS/U3Vs/ldGdXS2MGYP
m/baSzIfSkMyHLU4Sw3eVEywC8QxzAD0CZySJqR/fsrjzppy1TXw+esg8fJbvLI4
3+ytbYCM4on1MbO+JhK1XxKp0XWBOrRnnedWJgc0ZkYDhxAUuV6HxggirRYz3GCs
wBf6dO39aOjV6eq+hJ9BzN417zr5Z58W/wtrTOtGtVMSfDJxl268hibTRM7oLY1s
uishbV4dxFIXDN2oTsE4cRmohFM1v3vBq2Sm1M3xFaO05lLyClIvHubPKtMpfjTc
/WuEU5Ws1FNOUtTT2p3nPRrM0w5HCgQCf1HVAEyfFKSd2Nr/ljD4vDoYGcm/MIya
ktF07xOR6zsiFvA8zEghWlYvqajcUccnllnGDZfHwuxrhMxdAl2aM8oBEo2FbKPS
uwY+AqI02zw7vcXjr0BK+flFjc+9bkYpLTnaz2esjNpBaHGHB1c9DJ3rKWZz6GjO
aqwzTJumFSGI41cPoS8v6PxsPsfRsqaegnqNFZe59AWUjNulQjQOtNKxfNwkdu0u
No8oyfvYHOJXo7xQvnewxBoPPDi5r4+rxQvKeJwX0sybpdqoyKglOLf8RI4eDBEF
jr/+YtlC6Idv3zsfi/24iYGDhO8lFG7zzEl8sTKOoenwoO5VnWK5tHnNyVaneCRw
d8RdqO9wz6CMYcTHQ286T/z3Y2IxcnoKdFtuzg1xmqIytAx/8vyUzWbJ9bo8ng5+
JihxVkHZQ5JL/xi6Z2LnDYnuA7k8E2nOlHg3W6twOpiidVF037TicKYPGmpqnoFz
600H3jQ7sQOJ43hvpnvPZu8y2JZphYG8hJF4NgnJHTFOTRXL6dv7GcPyXHdwP6Ij
0hheLquDc8HHSk/fo98LmDQCNoQyx3+9pYbyeirYXm48gD5tvOIOT+nvyj4shaii
LB3IagkLIdFgPUbdIPY+JcWf8bKufX0AQMN0dM+agcMCffDn3QKBN6ZTC+YNKG3t
yFFjt9a5oxuIzJnpv/cwnTcwKifT/hx1+rv4S/Q+zEKrkmp3fimtxQNYdW3UFdBY
rnazfa78CyZF/m0oxPj/ttV5NoCAOa2a/cyce/9dhvHJWVSCgS1A29Y5s+g0hZge
vekVJiUEs7Utho88YdL3re0d9q2XCUsNkrjsaXwA+5J649Qmb8O4BR30RjOz6toX
EZLJ0j4HJewJmRqGysVMtBYtzFOmCD/+bXCysXkrcsi+b9TGYWwtCmWUChpgYKe+
xdmwFYhPSm2m+u8qcBLtte3zl9w1bNkuUqxXlHd/5ebCihc44hVgfJJq6pjoJtbs
uA6oEInPjfOqItW2PhwoAhI3MnwVZSdtd9fPcS4iT4vvqH0PHqyJv68m3/tNW+bB
U/NoRw4dL+/MblByogREekVOofHGM8/GJGaEbqzZFwyybXyDnnJoiiO5H0bkvyU6
GCuw/dPtXVVYN//+RQM81t3lfXL7iwk1kTKCiAcYxM76/tBSerSsQR6NeINlmWdK
icbpH4bN0eZiqlgutO3OoQoMx4NOz0C+EeSyj5x3P4l/xLZZH8lFyqR0i5U1LtJC
KgtRZurZ3/iEPL5kEGjI3pE4MqcblV73txIgab8Bew0+z2WNsJa62ru87TA9jThr
OpSneSc0tbZqWRzAOw7TdKhHWFyss0UyYwNS8xTzF5ddCZRLfQFHr5/st31hxEUd
aMyuiHHsk0sSGkx2Og3NKrrz4EXqNhVoTCTitApi6khybW0UCRvIwYatTIQfeuJ8
l1Ihul/4IqgWHcXTJC4T1AJTTMFhg5NwDt5ZuqeKHB6+Go5hfVwvPBWmijoKOZ7f
omiTk0quqJRkyqhaVps7+eNMn72Wqjcf1IOMAwQQEHi9IDnk+yk3bZTnsWPwUIog
u+70dBmkoaLKuCBNNG5ORYDyoOD6QROTUqUblIsCGfBAJvVkHuyEb0uywzkiHWr9
kyBg0zKpstX+3TrJUnW8VDRSGpDXAskG4frNW9l3YjQzEZ8yXWYJfgiQ8MInD9+M
x0tNcKwoKKuFRKkmqT/mlzzecRGDO8582s52ReO3ALRPXQltTmCQznycnZ9jw5cP
3n/I/J2lt7M6dHVlkG8Q/arJHXlU7wwDBWxL+1eiwRtvpRWLMv6/k5jL3xeafQOj
PEdikVfP14SR8/uk1mNAnlSQ/+xXjFYyQh9P8SFEOofRXBzTvZJ88PnpGp5Kmm5v
UDiDrn+WzwSzh6dxsha8uW9rDgVUIP6/SXntlM8L6KFF23WRbfzCz1XuPRZbSciv
OaGKc0CnlaDYCMMpoQnOi5z6Y7+/mCxei9wN9/keOnOGM45ovLTFEqnfUphHTkLF
HhDq3DzVhTYpxSrTebdAgL/YLtD4Ph3gke7QsR6THbYxp3/L7ES7Q0wgFotlWS8g
mgzZGFYtbCzoSlYK9avpRYFRu9f2ioM+lKNLzoAEiZnHssvYVisLJ5SGlou+sXP9
KiuCADT/uWGGu5axrkqVy1ZnB0nOdJtK0NG6l6PcnSEYv8aLL/7bp9ktoD6UQL3E
AfxSziLmQp44aeqPhp/3l5PzuD7YZuAUVzSKQSFuCrL5MrUT9F5Zwtg/eh989ruD
vjkkdvlX+s0qNLuoTcDjicYKx0PCItCbebEM1zWm0SSGGi/TJ/2EIwkkO3cbws00
gzeppbdeD6woKrUpXZQxUHqppOTyl6LWeL1FrTiaEDOriA8B+Xi1q9ZrEw/hHQx+
gLGknpdPWzEI96jTLdMdcpZ8ENZfkBCgPn7xuxMFQtyVf6CwS+uiTPaeEMkqgqZz
/L0E6PtF2qs/sVfCYc2ilEBxY8WS1oB8CM0VALzVf/cDnFlSGz9hU0hSzJ852EiT
EBrFA2Fw/cdRh4HFP1dZcYftgKeoqVFOvbtfc5XPkTUg1G306hcK9Rzvrdo8ZW9G
fToLwSYqKbwDS2qgksqGZaxyNHvgy+bH0lq6TwmTnNQdWsd9IyePy/+FWBl6mDgJ
qCIvIQhdenmL+r42eELxLP+Dt30d0/N1U/mpGNFjpEMUhrvbFU6Kwh7P9wbdQ7eU
kSNIc0In6mmryeioVWk/E5YzePCPU0IoXyDeoc1KihAan2clSf2U9ktjXUnzdimi
c/9mi4K/yEhvHdDh4MgjRjogy8RBSYZik7u3Mt4FTx07WqHD/TYeaaIczwLLKZNI
IXAHh1q7GyP0SRJALh+312inXXqusP0fN2G/3eT7zlVTHcXVtfDmlirT3WdMYuO7
4HQ5fbR6i4GkV7xoi2Ms3dUB72W5QU1So1iHC8tajSwzJTEAzZV9yTSOseooZIO5
RvfdL+B8s6fPWn73qHeF1ZpsOL3YNX59OF8V3TR0Y6LzbGzkae0suhKA82Tm7QnM
Kz/P1+KGHuRozCWOI9vQUQRYUivmIDLL4j8dj6irIpqqV+GhyxNnkZXjKJCVpPeb
u6NJ46jpxLMCn30VJ9TWpU2suMRFK9Qbgf/24PEEEyZ7maVD8gc3SdW31qZ2nK9R
OnnYgaJvySK3HcPK4vfQ/Qo8QItOJqwZ8iIfRm2Rojh4+rgdhxgFsBE4j+X8MqNc
qbLwqKUmqmnqfNuUlOOYnp3n9z6jsilyc3fPep3UR3aWXTSQB4gS24i+KZHqNnaZ
8HjgzMtg3j/WPn+Zen1S7OwYstfsoceEy7vmgJZ7Shpqk7KodCnTgfm00Hb/cUGg
pDOAoZ7m9IXWdwnHB56NwniBSrLyoPOGBCptNex9T/QpO7coHz2x+Jw8faY64P5j
mOUn6BPchgUX4IxNiDlxq6T7Lcxnu6ch6v5qS+PBp1SFwUNhRfvlTFITOmS+zLWX
aJ5aNdIVzIygpDmYJu1JjhApl6ql+fgChKAqcIZV52pDfW54KMPwH5fO9eXbc4V6
MAUEAmXbstnyQmMonllKYExt3f4Bws/hLXQBjDtLCAMH+9Yocqy/LEeHxXJA+OkX
lnHAKX0VhOwCOGTlX81jmzFqwhOFN3m9HKW9RBFCDwymHIRmj/2TlodDFqaaA2Pz
suBJwqHsnePW4czr739GgkeBorXDx7Zg3UBi4VImAWetWTTH58cyY0/BhJVs4eoa
YzxP+zKZB+2jmF5GNszLJq8xKnP9YlTW7nTD+xD7K+txSRBfdyKahlzUtJpcQj3U
ddAE6dZ/ojOacNPxhQYv5KWQR/EWIfCGFo/mte5Q1HpmanYgrEB6CvemytZbrz8j
SI85Id8n8dz2ApStAXsaPbipGXDNQMKn6kTEIPuy3sr9x9fHVRD22MEDAmrdGKEj
zTOQSp+AOyX58YkB1piUgwVYgOx9Uwp4DTP/2ZLsd5iLgHju2i7LwAPSvs+no66v
BT8whPgOZRbkX1/FFKY2cq7QehasTkiJZ0jkwIvqzcCYR7HNlqtl1gZ9lZiluOGW
lCeHcz1jLIB9o2RYbGnF5PjxBtYFQoyARsrJEr7jM87VRW0E0kXsoi8Z7MqfNlP+
jbryHO62XVKQu9SE0m+HcwsBXJc9XY8gN6b2v9s6X/JAIM2YILH8gB9PEZjvxSzW
q6uhqjAFPWwxCk4uEUzT3HTdhO4mhPFkvVIyKAxsYT24l5CkUuwoX3rxCQPo/mEY
uIjmZmRDhBFNmzcb86cZLYbDmqfSmEhyMGs0xSsEHQmyVmUMHbncuUdp0pSX0mMn
LZmqYI5A0JZZa7HGmcGaioXdEYD4hCFs6AEjB0+dKLBPimN5fjzD74tJfM/yRZUj
A60pQ8jih8Ep9FSIoadmzkLfhBoGE5kvN02uV7ooZ48sfesHQHMVu52r6UnGpoIg
DSYt7MEdFMg5ppMmVhCv50MZtAUwXITeaQws2iEfp+TlrYsAzrn4YkgspCEKJ0fA
IwrG5Sr9+ejHqsU2AdXhAaC5woV9/jlfHeWySzLt4V9u26YHGBHykWVGMjM2s/M4
1AVcH4T240XC+KpK400E98akA+crcF2h/reX0g9frAsBbFcAm48VlIBvbNSJqnMG
DzBSbuTizQal/i0DDExE/ZbxLqYgrZAnlMqjZcqh0gZyMLGK/YeJV16+LAvxtpzT
y+k6M2lSKXdE7w7Bd0HV1pQj4o5lj0U44p3pCV3FzC+iUbpHVoq7oBvH0Ur90Qmu
xgl5smpt2QBuG0nf0wcu6KZ4VlYn66Y44gH+UoqLPyWQSdmztCUnhOPyqEPOdXl5
reF6x8WXHduC3wpvYVXQB8ORLZ1FdZwSOBN6oA7Ou3cKVGVt5WsUAyex4F96tgOB
/TqIS6AwCSKnEx5HYsxCL91WSUtbJMuVNu0p02Ju5z5PZZo875hx/hrPOcRCMA29
iIFVxgiTYc9TMe35ynzcNcXIw6d3LWd+JZo5AxpVVtY/jUCwJ6FeZpjU3kRQrsLm
LgZtSTg/9+OOBID15DSGFQSTKWrkXmNz0IOV6/xZQ/TT6ExKPVMeDTmjZNO5LNKw
uoSLE2jYlFr8ROYgBXvpPX8pcBa8HCBRMkJjSOsOs/50ovaCjpmqkWHAnOwoAvPH
hDMEcb3K9Zy70rbVIBFPpHBPBJ/UdAzFZsRr2hS6AL5eefLGyItNwarlXE8RHlIP
TtVB2m8UHo/mjpVlqyseCuuhl0ECbKZKUYnwSyQT/A2SVTKKOytRfvfoDlyHU8b/
4CYVm/EZkc99qWpFfJOwRvo3rRmrGT40q34dmG5GD5MvCGVHS4xdGh0Huk7B7JDy
DlDj1G9Cf38ojNTwgIwURQ8paf24VjxJCT2HJtJktxgCNIHZpklRlp8vqE+HwzYu
sU8mmIII1QqwxXTd6OYFxI8ydNzTgLhn5cDaO8RBO+UV9acIeDmkNRay+IGEB0K5
/CRDzu5hhjHVxGvTBeXdyXHX6RokHOtJHVbbRdfoNlKkAWPUI26a/6sMBqacoXM7
2iC1unL9SlsCbFz2dkFWH2UXF6uMDjseb/sgwKNTTq7Dn7wMhLtS456+uZzTZuSn
SYoDNIHqckHBVEJu0HEzXED2aRgECScj+0fmpvuYNfv3ffBIVlUTISBQAmUwjTb6
+d6TtM2H04EGumj6v86p324OWZVQ6DsH+pQVWG/6ObldztAlc3wRdqlrho8SJwDz
2kuyxvk1AuZ99MSs8DtBm2ur7s6Rc5AHpgQNkJRiRcDhraCT1VvPrzvEcFvcyIiR
7sCdnbwbcnkMCdFWPAAbGYZo9yXpsIu581uCreMdxhBHaqdQlfjFv6CYcdVo+zvo
rW+B3GF7zzLhoeC4xig86P7zIiNTS0o/BnVjGSj1VOB8UTpP/+cpCZVp5MeliwvD
w40NItzcpZvLYgtg2gb6qlZXw07C16jgLKNzFsGPLAzbT/73YbaIvSOM8CP6x2zf
QPZnQWV/m+vUqboKylxskygJPPRbze4iXobvJ52cCh587SkTAihnEu8Geu+U4ErW
sYqJ/LlsbTKojNDH/lTkikr8lkFlKRBkV4nHg8R7nAzjzFdFI8Ft+WoR63GQs+RY
gJwYS9nMnU45K1+hrjcuzZ1UI9C6kPjyYurYSF3Hm0CO3Tndu9etdo0tCLb146Pa
3Eq/rwculJKxCAhEqan/22UgGV8BcB9/2tFJMwObvFjOlYSoUflW9n5P7E5RZWru
Sr8LpKnNU87NJy9wTKvG6cpR/K+e+4ayWqGnr2oLyWQp00Nr/lkECCug3m9RHfnL
Fz0HRcw4v9dKh9EyBuOATKaH01m0g6SZVD26ObMKm5nJYN5vNcFk7K5DzhBnOWNF
PdUAVvnpbjO+HHRI04VlXjbGffZ1qf9czSIPT7LA6nAYAejKeQyNjz3PGjx8x7r9
i0EH7hi/EQlJtQg38HDJfmpzbUqovUfzqCLBXVf6tKX55zSda8CgTi+hQXqzI5gD
KbAM0HFOsG+4j/OshXePm2GHQPGOMf83u3HGfPqxNlfNTDYcz1geU2TFzfTAQOMb
rXhBsQ88mp0naGQnTrC4NjJFOacfZhVUeuPsMETsnGvymADS+y1vgu3STHfqfP4e
fJJyLjVzEV7hZbpyBLoHXSzvO7ZSHoAeObbSOG4AaJrP2PxYYqDBXbuux+Ttw6GK
WwGFBf/OxG+4oOFXguRwCPQP/BzC8J6vC/OKg7sYVg4QwUipBQ+YX7q3YkORNe6c
ST8T/4Z5wTwHTFFtPczALrsfueeWp2legCNcXMN5rQiO22D2JEEqRUkBvE1R855i
C4jAyPHe+TsVLc8ZO/dPAB8c4bgNVpXo0p22HwXeT0R9/bCBLobXIZYxsvJtOCIP
+ly8VqCHfbFLNlTMZGSDI144Cu2NIUQrrBnAlRV8VESCqSA3hFc0zsaGHm+wbHR9
2viapdey+KSigbV2Uqjf9Y/p3yW0svVeOfziF39vbGkN3KbMia8Mq7y1HlKpb7r2
WaAkg4Hn/rjbInuixJLdxnzcjZlAsdW6v2CAEdHC/+R7icHTpokHU/MaxwAkgOKR
AgEvyJRQxvrH3kgPZZ0LSY5yvKWLGDBC+BE9C58Gq4LuCkP6VFnU3gf+R2dLlOKM
OG0cOLIOFh7QFMu8C0TOOtB+hxW22+mH2RzEWVRFz07mqYv7rdnzqIDOiCtab+dz
qm0ycG21jmKNcOTNwqntawIUlD9Yx65xzQ4QNJz6drzMd5eXCSZmVK1KWI/cCbos
iUSuyCPD8o3E5dTBLD6fs5TXpBXfslHeJkern+4lZXDQsG4JjoyBnP3ahhJWCF8T
qtATxLddbURSuYxZXHIDlJwY2Z3ggsIgyB74QYbGXsRj+DaKKIU1L1h9y13SYyQa
Jcq0Z84ETxUtFscPjdqCAmh5knwXl6kFc5AYMgscvKQZvveqVdst2jBbnVdnII+C
M4hx+uHx0ZLZ4Pvwiun6k7zsGFVoQvgoI7SBXdtHPdYWh5qg+NdcZeCIAlMSkFQK
Xl/wGTMbdIIlGicCCUSCGTGUXJ+x7Sc9zdtsBCAVsnF46TKfqBNYddgxMebWAIM2
ui8gHKlf4lGKCyoAj1dyJBYjsTnRGbHcNHhjykFi7eyXq/bQyScpQC4PS3w2DxEc
VTCpT1NVzZbLyLU5XclaHk0Hic4aYhvzuRZ9+jDVtg7IgKbX/8CRENQUaYsatbQM
U1ry+ZW45YvW1lkYJwCx8MHaC6SbnG8kqGfLYbT2u28ycuVYqeKoarbYni9n9P8/
DaQU0fRd5/or2sAFHq+WMcFGWbP1VqsB+9D1Au82Jsv+uFl9vin8er+Gkj4URnx2
SIHbjpRWBSMipC9h163wGsoaKCV4xDXL2GPqd0U+Xt8PDvKG86W6Rz779MjJLrup
pvuXg9NVdr+HUg7j6hLrf/lQXQMDqONptaXvStOSLZH63w9KMTOqqaBlEeU5f6ib
8puko0CGQsPPYG5/mZthKUHVSrzG7Gxw89nN0ilTNFYCyAqmvQBgIOkdRsxxTXYJ
QwAjl0bVLKRgfAcjky7mJ1DYWF6M3Gb/5GGE0jlVYQfls0MSvNYAP5/Ey4NQIsXt
OAeAScgloMN6OFfM45ZjsNhAyTP5BqjhOFKxilehv1yTnqW+2T4GdQQF0J1B2fZc
jIJvXdaKdYXgSSnvwojFAvZxcDlRP0Yvn7Xhp2KizIiBbAuneTVd+N1qn/cCUgNx
VmU5ckV5fq1DEEcAN1hY/9QefEXWifo6SLArBHf79agdRZkKSwwLoogNFLzpXNFc
EcMfBh1et8iaYMUnY9OaBcfCKeEuRPnc5zQXb7MQc8RApLHZt/63gabxUY6guThS
1uZpukLQcDth4nygB0nj0uX58h3NPgb2Vc9C8ZO1MQ+iT6ygiCTpNamKqQL6JF8Z
TJ9Sy8UjDU2+wIOaFsTCEykq1ZvJ2IscY1UBztGc/upMRvJMYc+5A8hOHTBnhlWV
Vq24oD60+oIdJc5UTqLA7dmcROa8cDz8cYNGmEVZrqvwyFPh4eJVnCgK7QLiXzXe
lVRAaksGAk1Q0Di9/1mzU+UB9j4D4dIP9lWoTY7Z08NguDxh3LXIm7LOoy3PVe82
Mxed7UzTe91N3+DSxSHXG3qKqZ895/XEBujkEprBpIPZ98v7K1UShvstuwEbi840
1uVkBSNvBiFSeQAAfNfDNIycKlxfr7TYllODLW/H1H7Gg53iPM7ysi46ClLIW81h
LHQoiFDXLYrTqlUN+iPfL3/0r5QUbO+M75YQWa8c8NoF/0tRUOWyQz1BAMYsJzdX
ea+k/QIKOsib/5VjzHrDD1VCfVddQ8rJ7zhdvCgXwxI4aiiCHSt7Vck3fePkVw3p
Swq04iSfkv655mTzGcs+kYGbarJed6t4/NsKn9CrPMxT7yiVh+2fEYfAqXr0Fgg+
lW7DPk/SFjpYoZ2jRnv5V9yO5U7ciCZHnY9Qh8ZSw9s1hhpztOG+g+9Vhz6xm1f1
9sBUa2aonwZO4xkj8Ki1MJKYJNTv2vWmvpN1msJoZU3AjeCkGDxpd39QMUaSqjtZ
+mVRvpiXzQX6TpW5ly5B4brMH4jSo1EJBHt5fPMd+La62uwOfdaebPyIak6EQbzq
+Kl1sp1ZfxTUIaxtqAtUDZEwF8U8S9fctKjA4ro6BH0Fo0UjkaQxXLwu3zQml0G0
KQZeDKsEXnZd1kicVqmk/KdZW4v3NbnYprx/1pXB+/nivbzgoP1/h/vKjxiGYlXz
OSvN0qliT4++IHuN/gCOpDefwv+x2F00b9xR7XK+YCM7Iq0LgYhsPTmXvo0ihVFk
/rxRoP3I3LJWvqckdzn1Ewd70scW7zmZpfT8uOvBRlvQLv0/UByebb/NH8BH13tM
qjh7SV/tELsjWh9WRlV+rQwlfdctmLhtUH7GjsKUzceGhZf4sunCdvTYw1G5XLR4
oXUvni5SaiGHHh5SmlEJYmbsJZVPqqVVGeAHaWK1S5JIqAt8DBue+yjK2nD11KXo
CmqVRYHKHgh4IDHl1pmgveWzHs/STwWeHoxWqgyCSR/4R79YrGWqWDDlWsUFUcB1
+PZOffX3L4beludq5Fd/V4nh8VYcC/ksIff1saYjTA5oIsodRWss2tZR6hOiyHv7
coCd2rTyp67PDyE7mPiAB59BZugdjP3dKcJvd5O/kKY4ffmIMipPr0YTbv372O8i
occ2fYoVRvWgfwel9elroPBlTuDkk0xotcVHZRXJDVNfYBiBU7VSHx9iqtWeiLJg
8Xqrv+Sin7gcMTIuWUD7TEw2+dZeH9FOsitBPvJ7SxImzB4H/E67n4drM8MNL3Ck
YHpUt9D6xDBlE+qZa6AKA6TEAMQ9HGXZV0JdfA1gC5g4HdCrYivRuhr4wlElhhnC
TGZzednRqneZWqFhkJmVoajr39nxSGBUG8OyFekcjHN0E3DyELohdTYeefedxMWA
JVcTgswUPTrrVG1/IaOxTEr6QoR9p9gXxUBs4gmjHOgbxZ4VNjaaPQiPoDOHw2I6
jI6lg3e+X1IGOpcl3AVJyvfETdD7s7lJl/4pSRKqR8/SG5sNvF9/BVNW8SGvcHxw
DdA8XEj4d44AAD3s70WwzmesbZGsK2a+Kd9LNUMhzr/WzOeMIy96mf7GRWWmdl3d
+LMz8wIb/MnnyMRSjbKB9RHKy4vMDXXiV6v0cRyZJirPfrGhPKPHJzL+R/X8pAri
JeBfnqV34yG8pYyYiVtDsd2+wf6k6tf0BiRaqayR6JycRN0VWdPSPl6aXoTtiEeo
rXz5ZX8fTAu0zwPQkbSGERRGDIAebuP90/xnm/aj7hy6lwex5BduJglLiOGiAoDi
OV8lLAtebJeV1dSpfJQSgf/HYRHac5wF/G2CfIer9swnYB0TLWdwgUMO4mAUeRUi
DRaBsIUBQBe8qhlOxJZp2YH4y9H6ABwaDy6klW+BaKi+Sh6LCnAEY2fmtw1ScalU
IBcp6Y0VgKUl75+fTtZMJJPD2LAY24JDsxUjwZ+NZvcyk+Ukh+U1I2f+6S+HYPP1
yclJnTVIsErOsYzhbomNNe9vuYwDQCeAe8h8EZmKCod0b4TShzrWP3RdULdqwxEs
g6TIEmjqS0wJYB65RjcTwy0ILG0OMFiReJ2RYAv4tIw0eqyODqz4QhPs1Fh0oY30
8duTqtF1sxHpjttuxOcawpgAQolHpBK1LhDKSDXhCGQXWYBhCLM9jKlDNIXx7FqX
mzQcJsff5ikqNLjfIO1sc5kteiT5dkK7aim2o8N6bGrSbfOeb5TjrcMe07+IWWXx
gvxz3sHzR9BkiE/OVyqK4q+hA/i5EcwKLdprSaDA17q6yYFcdN4Ii3/SN2v8VvDC
jHDOtDFmAt8bynyVpEslsMSj6W4eAvpoDsnJecVHzz+Ie2CruhbrSyfKY6ffFRA8
t6fnTLn1YXM/SHX549y0A45CeL0tW9GKwYHMHtJGzaAE6Q8q3e2FNt2oopNRb5Oz
l9yQn+uIDdeSLhcmPhw4nyu5KANOnmgmv0yMarkWUhTUtWeARkwZv3wyOb3qkYIc
aUPvU5mIApSOWHwF5Pbas8U1sevMYuIwXxzITb1DkjEOYZbokSb6Km0q+M+dPbEw
hv2WyQuibdFi8COB2bl63fApSPRHAhFysHUV3otFtXNyOwLJzcRC99U/BiYOG7IB
ZliCXPBuA0HZLzKXAiL9OU1+TOI+M3hwCcRhGoRdRbUxDtkaFhVoM/FM9KSl/5Id
L3CjFz9WGbjN97OuLCHrktUzam8Nwe1CAkYgbfWH9wVNyzVr/qvsmc+8UTxcSUqk
CWArnwWfba8k08wb8VbAwfYTEviCoU0c6j66DjVvQ4ETgrzgw+/UT+7lX/+tVf5N
NaW8168GWj9ZIgHXLTYCa3/k+WuWtiupWYuGrxFQiocS+0zCujjaXGODNROv/6Ot
ovW1bNtAr/BffgbpRUyWbkleyJkuWyGn+5HxIFscMnc8nnTaJaH9jK4xIKIHH/MN
UO48ItqJj8iw43x60L5AbxbONB4G924GOb1OMPDrIJhzHU8IW2t9L2t3XsUFJGjh
FE4cfSIawdnPO9+A8BxMZnUj7CMIdFn3WSC9GGf2P3n+9MiKBcz35mdKxn0gkTXy
PLPf1M5dpHkXd74/1ASOwEZ7hm/UKpBV+79FlvZPTWDljAsrtWPp90Q83UErpEtA
Dnh2c//9NdYSUf08f114hRE+BlxDcjiggoswcfQ4ZKJrwYEM7zgkO4uDBEVVEIhl
jPyi7MdSzKTe6LhREXN0RszCh1x8TYfJGJE63Is7YpIN6nxsUSPNx0M3QtcM/N4x
DBDvf86DmPDOlw2cxviSQwKrso5vfbGKy+xd8jpB3B52icOr7d0wAXzaqPoK26TU
5WfoDBi7Q9vUUtDGXeNch1KI+1W8GkcoOy7ceXL0uo2srI+cMz8o1UzHPHyXvAXm
2AySaxln5dAnLXk85aaOXPcNNKDXGI/lOvXhfvOMpNMBvpscs3Jlwxw/Z/jx5A9z
j08Q9yNhp+d8Z76a9c96wMuesKI0hcHO4183VTwxxugqlfBmheSGSVkMP8d5eeXt
cGx0ITJfWiz2M2vhsSmlGW2HJQ0YM4exY5Ia64sk1MtvgCUH6YQo9I76YB6/49eB
lwNRZIiWlS3JTodLp99F4eWnlRdd8Xsyi7Ln33zKO6wlnhBwE6moC6WhhS5mEg6q
fJOZjwEsJ0J9ZnLZ3vYQLtUUcKhg2/bBUXw4LAmDd7cGCMEe0+wxTuacouLvRIBc
5aBaeiexETEvem5xGBfuM5W9Yn6+VJhnD4iTO60GhilrCrsog+gViA5+KrQ/DLES
nRw7Ylh1zh+r5Hg0sbRhR3vAypnC/51nfejgmbA+9gRzAuAlhsjrjCl7pIXuZagA
+I1/s3zWZN6X9UhVWy/rLlTkAgLD436e6sR0brxXlLGHyAWy10zLtTzoc1z4o4Yx
0gwDSlNkHNH1TiHgNtMy6gMCDMZnQPPrzoeTT7AsK9TnBboULBkofSwx+W6zyoMQ
ALilVoRt8boW8zORmt7dvSGbD/0FR1wgHX0k3yv4hygme3qeXQgX7iu8j7CLOTvn
XIqaMfEEu+PCnjUsy4T0d2ufZivE7t7wyE9hZIzMKt3hGmiSfjAiGCu/ci4fmjOB
ZN2Lk6xyv1k6uP++v3ZMtM6mAbUoD7N1fww3L+IjE83ao8nbVOKOsMY/9R5M28RI
LM/MkW+aL5qx47c2qwJldiweH9uXTlkx53oTyS8m5kC/3/27qeAMwmSYX55U2Q/2
Rc6vWf7Tw6s7Qd1V8/trL3uwRE3gjTi4P/i9tMB+joEn2KYcdRDeJ9Jix1H6Cd0q
mQC9WkYbzt5EDGId2UneGhAccfpyjZNaenPhzMED4HAJCaC/xG5nxY0Wqc5dg7xk
kwYPaAK5wa4Kqw/5bzgsuyoVPhDleFiv98QWlEAKHZ/0zf9sGV6KAARagAmT8SY6
b21YsW0YYfKTlqwGy/XTvUMXPX9ajgZ2eGsw4FQraaGsjoxjE+nuabYDkNwyX357
mm+ZTCE8XwtO4ACzxhxWJS7wGu0snhoLgPPOpalvCNj4E2m1+Xn1K0zTUBWLPHYU
aHks864/QjoPzHHEoDMQhZEcLZZkMsDqk76MYSiDoYffAhjoynNjHaOJxWe76FUk
rZ9bqC70ThSIgZBuycNfMj+4vIjbDD5AA1IQVzj5GVRzmTHhMzsa0rPb39jIQIss
2CCKAuZXfA1dih5ma/jEbY35vVZbLNs+59JPNE1L6AVW9BzraVHdQcAC73MwObm5
bYG+lBKgEwtTT7lEAFFwS2pXdTES2PFE770JbCvLP3Arxge4X5YCiBnvFjszRaOW
yNZo4Mol6QM498MPbXqnuzCMCVeAN/OQfrNnTzTLcPUs0ytU5bWusRIxSQZWwBb6
GRue+62SAmRsisaGP9qwbIVskE6i3AZImbHhvPE5CxzwuPF8t9dZZYeC/QmI/5sP
VbeiKEp8jINdT7qZMeqggIfPMl7JpozzosJhVzia0AOsQxaz91zAa+C3VxgSY1Xv
sk+LcJ1KM4mIZexLJVyCqZTWp+bCY9tEP0mf2t5VPuBqbRcnA9Hplwddjq8OM6xU
wgblAobiNvlMK3aPCyTXZG9sJE1YPJwjjHUwUShDPs2k0xefhE6ET+KyuQuait/O
OO6azKyAw2Dr/KU/J1jyK6VWfkOi9sa79xVGzeh1clfAs+XkiafiVxr04wMUVtSw
9AAzryn5MBpA3CxO8S1EChV80Nx0AgJI7SMAkTXeiTicIheakJSGWtq1qXUnUmHw
ify9EBPB/5djwRpYFVmzBK7PuTarpGcikrSaNqb/tvyqr2El2CrrIG7w0jCH62Rz
5gPjWb/Klr05GC/qskY/puPJJF9sid5Ri+bH3JbNzHaDxcR78P8GEyWtVvfFwqtj
sogponuHvGRcK+qH4FJQk4HdWlN/bVQFQ8BRsxDIDhbCgLIDjozW7tzf5Ce/jnuf
T7eiWAAg2HAmPubWzyEwdDKHtCwlPr0BCFpRvMTBmYr0EFgh3beM6tbLDZPgchmk
5+LDFhxr4AXyXrIJnXWrhwn0ra4iJblb6ncmIBfAmuxSdRNz32u+8cxZGFVJ0AW9
S97+KF8Zapud5qhut3n9Mko7ytIFqnu9pYpMMYTG9kUtnbsSUQZtDAoajHbPzvEi
a25aBn5JpPAWy0aq6IcT5IFTBl4q+C7Vq7dM7NUM+W2Ux6JLLMDTtSDBmMOK2Qco
qv+LtN5VMam2j1l4UniuuXpgiNtBQbx1/AfNEnapSuzx26kEeXXAgnWXDebPhN6w
ncN0PPLyQjZj0Uoqzq7znmko/eTIqn8hk9Kfp2GC0L4tU1oUYyaZTn0PTPAqU4Wf
lywLFoh2yXUJkYhVljme0xh7FcVJNZFQfHlkbk+r3AlLfehILt4SXXkmc2kMRgxD
3z4/grTW+Kvzhz99tqmqsb+hbt4nMxPx6P/U47+HxsK0iZI3mnEJ61bWoewaR7Tv
fGV1ggiXmHRBO4l+wrsZf8cSajA0qH6tp7detVeksAp6XV4yibjItZXOgW6o94ry
12l2ZggAzK5A1+wM/vPYPQNlHK1X/Kk2spAMGqbUfpRsaSlIQWTERfKhW7sQuBt9
XCcqCP3NUAnVjsTKCXFDGl1I/x5+5HpEFGe+7hXl/RQOJsx0vWorW5s7BI4IXc0z
tWEjYKP7rjxAXWByN9KsKa68fs13rpGeKgTvlSydEeCm5KWxeuvnBngTuJBl9lUk
TdUyXhUU32mfDiBjf740diK85VqH3fDdXLWYX29uIJxcgQQuFyJAbibhG4bKferm
av5QIIL2HHH1+XONTTj9L3J3FUY5NeQBKBsC2P2eBmzv5ddV0fMXeRAFJll428+2
f6pBdt9UH05rSQVVToURMhzxe30U3wD5d8A8qPjjlAYGL+PnzPGgQERvrj8aqnj2
XMONFKs8yD0UhgiTesBKlgPHPgHsL45MhS3W3A3Al+QTuje8kKoFb0me/Q+q8buw
NPXTJS4mojIpsvIsOyXKOdqRKphvDFN9l7/8h3RicvNETwYCuIz8lFHE79O3nCew
nbIbC4oHpCrYnNFxD7r1MxS+eunBfA5c9z+aGxgHwnY8jtjhR0itgYPpx0pxui/d
/dK2FD9VkeL6HDNfLQKx9mq8EeZojoAi6Ap4ue+wVQXbsooEEUiaYe2JArYj+cKj
Q22X4fh30rSSRDcqBZvSlAQYNXN2YgdA9Tjdsr5RQTbMW2nrrBCk8VM02uaA0Oe4
EHKAKZ+3ccKIjGUcyxmRsPUIDvlE5KpplQ4CPYeTXiZ0OpFVxj2uQOK6fTbD8mAc
PCyMNm5cuq+U+0+dPBAseIcQ5Rn1SZFl3pZGl6ARNWWcmTAWfk8ubGpAfQ+EcGJP
AhDaj+39gUA0oPPNbwCSc5ZQXi2HwfOwXgut/LxQWjX58QPzQCEPoaXI2+J6SkhR
SRpTD7TK71c4l4lC2irUMAQRJm1oE5y2c1BB6XlW/rieKPPdhq65/0L5aCaVA294
b7clRSobYLi/zFsjpPpoP3VBVu/w+mpwS5LiZMiwjIA8PBNHhgpjTXdPBhCilNSf
7XDto32hXXVbwTZZBa9IQ4rM5TnLh+UclyB/W6NczC/j//wjbn7C7f2pUk/pnkOU
eRyktTNWB0xTMHwy6NllelIGv1oWZnCu3wAbp03ddjtDV2WLl3Lx03h4bGMJC8sN
QSqaOSkhrnVbdDJhmyya1J4o5veI+G1oyZaLD8gOruyPkrHck974eTDe/eFDIpP9
/67wqPFN1s3mKXwbnGwvn+qRqX1DRUj8k6MuIBVX/oOrneRexC1QCbRoG24n7J62
N/CiZwMJqNO2K0sAQdfiMzVsg0zzq3QtCeaUfkKb/57UBl/Ulr7jaza6/LZNywBi
nifspTxrbo83XVZfXTri1b9y2cnHxfOAWFC6jrH9bb9foG8u9CC+nmFowb4HiYPy
kQY6GevKS8E6lzUITYSyk3S5ldu5qYRQzj7Xe3JycEur9VyKXTPGxKRUL8olNq4Q
hEdS62pootLeCNg3kgQpZwdW1xjh5iFQ/WihNcYjyD8JUUREJSovgU3Ts5YlhCJu
lgQAFquPhDnrqyJ3E55c30zun5hVc657XUIHhf0dqyYaIEOiLUR4Xq6TOL7ztZ8L
l85FSmagvuI1zWBLw2Kp95zaNZvOfcccvTCywAMt+B5YJfsXDaE7yFJEM1YOmsZ0
YGikzXe2WE12V95mrsHpadOT2rvIbeH40mCrzs+N3wMgKd2zpWGrNAY9NzPFzJKo
Tqwq29bXZjhlgbwTpa1PavmqSCYHdck7fCom6ApUUoP7WBcMlV/ueGkeQaOa3XIc
zPD9TgLaVqDxd2+d1mxlk/B5vGZV+QYF91mhPIL8dwxFHVeU75Ta1OfJsvc2LHUV
Jh9mnlfss/Nue285JwAaASb4CHbXBo+2G0DEJovyN0BgjFsoT+u8HngcqyzDajcF
6RdAENkjGf56zYZmQCogVoRNhQnXwu2V3NEOoeirWfqrPVMJ91pGxa2XC4FpikqD
ilOd/ohaEWItPsJ/3cEkhFjHvkLO3Xzl1A9leyk0/p3gU30kLbOrxox3lbsD781L
aD8L/8MjDAPV0VEosJEX5nbwOSpXQm9kkpn4hFzO8FQluld4MPlVbigPrgzXV3g2
VB03pgK2oh7yS9k5uLR3tZbnCATg41tPPs2BZE5cNUJUKXoTmD3qY/fajz71WQ8W
qOQ8G2zRpz0fzTNijRR5Fmp44t9JgHhVeSBrdvsnXMHTdGilotHff5ow1NFN8N29
AbKZ9Zy4CLFgrmqtCfzdTJYxDtBt59gLw4GNF+H5MNKSKMziC6sqhtOHZm1ZcK2Y
AMs+5iYH/etfxQ5K0WvgUpso1GWGZrzzohnRA48AjsB1fqbH6qbhBnILSPGU+5HO
lB9JrKGQrRdawBwSeWwewwiFpknkbwJT0hpUES2zJrrVoEoI5iOl72QObueaMW5R
dvnGOC98s7SXW/Vxg+RonK13vug0YyAvBD5LxBcGMUzCHY+GYDFC5BWbW2PcDACs
3eKMx5t16Sb9x/oPtat/fAsQGLDjtFn0VOBvKl+UzmVXgkJmxvyIWhEOj4ZSqjZz
6NCwqTwN8IsQe7z+nFMNrAtI2ubUk4H8Ivcarft6UKc5siG04srZZtAtD2zGZ25n
s+UBqi5ZSCMRqnrSLPUy2HPcxTytTOqvPL+iwyKB3MTP2lRDdte6xCudOAPwBXpd
qo13lRS8rLAa+zVMqSPYBsTZKlib6/5YYcn7VevLJ5ltVrGbbkok90ZXQ66f3wid
Ms3ns4zoM+hatH8ahjTNmXBN8mbNmTBFz1DZT33TXJ3+QqYlw5OCZ6DH2W5sP3ab
GhQcdyJ+5d1h6/ct9w1NjrPqRmEL0d0TOFbWhJ8PmMuig1TtN+rtuoT8FJpsLKMe
mJJF6jwolmZBMegkm+8Bc/NquC+7Te6GPSjTupLi6VLLZ0GdDw/VgSOgj7nPba/o
pqMxNGcCweD6bdWFLFFHqeeJeUuUby9JBKJV0rfnOamnp/hHn39TzGylbZaBF66y
2IGOnBX95ayatXQRmh+qo+uwPooaptZ9CoQnsRy2KcKu9PkmQtIlCrzFw214aciM
wsjYvwz8l7mue5ck4NGCzmjKtlmJ6Ls/GEVgQY1C8n6SXzwOONa04r8FSA9q7yZD
r9M2UTCfNAmXqomhD8wTFWokB0Lad2T8uG14WoM3lsx5v4rUzYVssUtuPrO9rDAV
rxVAT+/lkIS3ZIFK2ErRKdqe2zkTpZLsAk71kH4+OYpvUkandHOe9mYNSUZOKuen
H5QePu1VlrCkY5ruKxdIzFbgpUXAKwWL9yTD/giQ7MOG+vN++u94NqqJbNxqx270
6Xb8vCwaqaW2XmMA47khV8XhXoyJg5ehBcw29IhPSt0FRPgz/h+Q4l6apkaCCjUN
vlKlLN78HAgIGAeRrxYNvbuI8Nkb61mbSBh3kvqo5EpqhM/rghnxpPFDaOPeFz/w
9ud1lNVxNQgtrDQb3ADJIVMuBKsrvgFwUQ6PJHKrw7EFiHNyedQTur/ll88CPQjV
O4A+0r6AVITilcD7WTNac1mISmSE/ibWDb3UfSqos7IY/HX5saQJ1vtJG7ESLXEI
3WpPDJZyNtd/ea9bhDEsZa9747xLyftnuFqhcDyh7tO1m8hBs92Royh2czODDGwG
1QUocuLtAnCOKnbOO81XXDeDIKFinOuyzziFEZtwAyUHbxv5P/wUO6lThaHB0Tbw
f9KKzuQdBXtU7ORiIt/YJNSTcSTWJCy/a3ZvQ8plHR9Fxsm5QIoCRT/DxxRKICCr
9HPH3XqPcBvO5opCOw5pVTigJqXpCDx1aW6Hw5o8JZjMUt/Ikhw7Uk1F/Wet1QwJ
q9kJajZAD9EkLkoGqxIYxg2Ek3TVnmxRpPUIcTUYIOaGpESOxbvAJhnv87Fm78Ct
mRvBvNVISseOy/NGxPmx7SrwFMLeOqGN3QFQpqEM7Tiz2gKGc35+R9UHIL5Es6Ht
c920p5+eqEmSYL3FOjlXeBpdNj/VSlt/+l7t7aKSMeUdcjbuNkfjfxvGbOxOb/ZH
cQDkbZ1nU1f9pd3bM9/tuaOBBF0MTMgFACWeLQriTUWGWG/9LpSE5gkG4JRej1cp
pCzvQSybmBz0VaLa7//hFGk479PnrahHva9BPRLO0+PxXQAGEAfi5FsVSS+vjSd8
iens6wysR+8p/AEdryDsW94t+ryhsrBsJfhHleXwqy7yLpuj69oP6i+HlNkDmKE1
f0lRvtwiM8AupD0LWgv34oFlhpEhBUib9ftAjMi75VdGQybjLwaTbKQE1clUCC+d
cJXKT2tiYL8SHYWAhn2A0RmzKMdK1l8huTax6v5NAPsImHl7ltdR9qrH0dZUXVfW
fahlIa0+/HqKAudNaKBHJefZIPpXpsa5qyhu2tgv21s+5oVDVdgp4lsgAh1klk6z
xHDCbUFtb6XPj+djNWAdUXjnkzm+wfHQJ4ul4u2RPI+JxOcONIXt2zZgVEmes+Bm
/eljZztKwUrDWhDgomM0Hr6jEPuP/sJxat6abgpTGRrbspuXvmAJbkfVAp7oJSFb
i7albAK3gShzxLuI1NyaGcysKuyZ6TRKXVzkJONSauDbjznqsGCznzV/IidDCN7O
4lIJWkuXaFL0WHjd4q8k2ucvDCOoaufHHG5sWvFxKJFcviUcfS/lwlydgk0/ffB3
Ac9w3BN/KHEsQAbrQQ8NSgbN8olsZ9obsqhZ5kY6rIYA84xf5J/u2BMXFbWohAmz
m3fqmLRHyr5wAcq3JBAzRMSYsGZl+XIFMfAr6jU3KgFHwTvnKlZNPfkfI45ittpI
oH9kgpwHPRzj5XBBFr02UkMdjcZ4CSk0lLkwgtC/RhlSYj3ka2UWhUI5RIfwFowg
Msiqm9gLkE9JfKyFwt/JkZ/OII5s4lLxPEVhYNJpWH8wQUkapxDyyQ4LVh3a4jC6
QNGZzIF9IjEGd0pssxMRV8nV4VwkwozthmbHe+b4XQkgDvzcaiB3qv4CsrbGAAGO
rI9sWM77jTR6St5fa4Cqq209UqiHz3cnoy6CeQH0JqLSa6/RLudt28y2GVkB8su2
wNUBh4LUoL5xC0gGdQWprx9O5yCIJBj31n3mB0XROUOOyBdyEsJ9ogfbBqEeW4+3
sS70PzGD5ems3BEOB0Y3WqnFyZZ1bzAqVcGX8b1blqeg8krS9g1AmupOF6NsjfC5
Wclzy8NHz5Mnxeq6Kxepa1V0ILK8z8puvO/ZaZDSYbzXjY87vTcRhX4ppUzWHtp4
7oaJL5bC/y0bOemew38SzlOAGYs50eGVfF5OpfF5lg5LkJEK//niEB/nPhLZHiG4
2/xIPYiClHl4Kcys1fQD1UM+KnRV44q24WtU/oWb5GYmGUBapSwCmqXHWXj/QHnd
5/Y3cRwSXP6/xooCEE3ibH1j8G+2aZgmUzC3bdDh2QwoamI9XyLMFx/jUnSio4iN
DiZYye/Sq1WBj8VhIpRLgZmV0AC0/fgUSY/CNz9LMWXwrRwufyebRicL1mqay2LS
WVBQ1CoiKDKUC5YLgZcyNIlry1DFW1BSU/MTmNJbWbLxdJjq5GANSPh0Ikk8f2Qz
hAMZauQntYDtUKZYf4XEEG/kz+q7TCf4ZmOYsb8AFY3f4THgY4dU956qiOdCs9qL
+2Loiu33Yqdu+VhdZ76Jz82yFwYgTWjzvilvmUTlNBtzUEZMBGR3Qc3EfQKI1Z+7
EVMF+eM/a4sgRPqBWUoVztENh9PXOZtfcTcGS64jG/caQ8dg62qHwxZPzI8Oa8gJ
yWlWs2RHqOOtL3tSho46k6hQ7fisUc/dmZEapwGCKTCHkdVvuYMHL6pWBqiQ6gnR
IrdukUgYr61gEhnwL0LvDy/YHsYMIdXT/SapLze8H+lF1IOpsjV381OEjFkou0aC
sOUyJwN6hLksqtF8pmJyUkqzXS6bMAmf9PQfXMEQ5fH3MA3ScZVaEjQG/8YynEa/
ujQmx7/SGx2Nj5AZiU9xH9S/osOU1jJWM8a2vkJtuo0lI/TL47j4kgSIHv48nJps
QssvWseejKansznGnD6AL5Xx1fVhobw09yT6dHJCXmrmc+6r0UYNzSkXc29iKw7U
fUR5GWP/6PQxD97lhapwAw1VD6Vi9EHv7wedX5EO2OYV3f7OnYSi/K9z4rW0x5nH
r7EtAcKArrOAJcG4TdAz95ks+NUsev9ChLMpi8Rzuf6W7ggWJ5bQrQ34YPcDtPNL
jTS7xy9uoKs61yjJIACAjgAbz3Ic8kQq+y39rJyxeWamB43z5z1cFiNJARdESaiG
ad9Oh0laH45zxrRbS84dy62FtF3jYCVqeTPG9h6MRRZHLdPrkM5OrjmwLHyGKNAM
P3kCDbmoDv7ysiOnn7f+RRm/uKgoIlqoRKKOs7HeJbNNRYhvkMcrBH37ZAWPKGVR
1wa8J0L83+tFYZvdQN7XtvNF15qNVzfyN6O2efhZiIH0IA0JDq9n9A2in3olKw/K
+MIrT+owSMAuTkPhyJtQ0Rjg9XgniKG1JgadJmjgII48y590WscW+pQmjXPnhpMj
wqnKRsrveqbKIjgZQjkdvjcbQ5XxfOkNXm04JQFIngc/RI8Xgvvnpt/z9OJUQ+WU
DesfoWgW24kxaY13xYGbqn052zNzjzLRbAukbGpQsqQsds1vg/zSp5MeXxdeBu/H
c1uEKXKwpe7KY2DgF7bE3wAbvT9jiK8ZGO2VuENlMRMzWlX22EV2MmbJH7GYxR50
/n+WkHurnm+Sa9z10gvpDLv6TIAzZPlj5Fi0udQpQmFxMIc4sNeQM8DX1ijopbrf
YjTPwFgmVN/sMNFbaUEOBAwPPJeCIgCmrZGOSSibUMkMhlc7L7uD0tkqXUoccn3D
fHxzpKV71nTe7MZjjgy+xzfclGT+gNG7M/D56vQaCJa8BCjNlyextoK/r77BYs9f
YqxeWozN42FN8YXiTY3V6oOD4PGAVRfcJIASJsHhPA3bZ/6Ebb3weQJ9olJg52uX
o5inaR8pH7HtV98bEcOI5DWVrfwFAcz7AOBvboXqLydTcLzmmv4m1sD9Ol6tFWx2
XvhgRmhotlCTX7rKd5m7WZWEdPY7Spyc7PjhhjAJ+phduvEQvLgG1UVC020L5/9B
RO3Y3B1V5G9g/OYTvGIWX9O0aUCplc4RQqwlquQNOC8M+ub1P5QQqExHhadbxsQx
3ZMzK1jbFh/iZpT1iDpPz9nIA5+MajoUCIERB+/oKDg0chJx3+ogrPozc4vZhkYJ
Vy9R6QUleCp4WkA6Dl2UdZQ1fpiqHJ02K3sytyrtItvMunIL5OissBxUkdxx3mxe
r4X/UhYSCqW1uVQ0aHwWBBmhlzXhFDUGxXAeH1c0Hi9GzPcEJAPeMy/tcZjV9KMx
2rVNrKSwVWncNPrxkG5hdqjjV1zeshGf8XmSJnKSGh06otA6T/1a/M1hhz+N8gtO
R+4WNTVc8BFwvUnLuZ/L9eNeaiQj6mvfBDQkIZveLJHC8yjbIPMtjJnaSXfNsSQD
gOmG4g4s8sV8syRR1Plpu52HVANSjDhR73uGKomo7xxZmOCO2m6db/aqPV8jZVcj
+DRlZHOekpbcBf0yTBI4CK/HIsnSd/pU89aFCSZV/laukNgvCW3vcS1G4QMWf899
G34xWaS1JVeOYmx54ob5yR+1VtXevz4AA6f+6pk/Puw/evGajG5cxQBceTgxFSpe
VZIyC5jWL8FAFJdnAJ+qvvFZqFfWGn/5EENrQQXt/kMPsu9hH2kUCftjEWpyiPlT
Zr0D709yRxYC9BqqK+QDr+Cw6+JI5vzP1lQi42Jh2hCFHIVEkdVilOxgknPsnrml
8f80OHeRroIUBQ/af71icSXG+jDsq/Kq+ruLX97Ejjf6MEcSmjIehxU6Sexw04Bl
0exB7kOsBgo965Y8ZtuXaHqYncoCIooRb9TXiWoDYRF4yliZhE4Wcfh9TfCcymGx
g9NjhFN6xdpOpxniU+KAUHW+uANWwoFHyGatoylEi3rBnwhBjYWaK2wF65DOR7O7
CEkKZZ6XNIhx78iEkOOFmI/YGqcwvudQPazJWzARkziHVkIWGxY7O5hm7O8tG+uG
3AmRtGedIEUB353tRcnLp9TQjVGNKDirfVcaVZEzcaA9LRplQ0wHuf66wblaiuwl
G0NwzJQukgqaaTqYkvaayFbtiu5S+3uL0zXztSy8RZirXa6ayoU8B5KR0yi7iCVt
l5bEUYx5asiRSzYZ/p9FdaxGtjZZgUxa5gU1l5aT7fN1cJZ7ObL3EVQkfvOzC64Z
p+Ij1jKf4fuP6FrOWZGzabqqLcKJl84uRyH67ioV7wPrF1B09AmGQwTvQq9PB9en
fsZrIUOLH9UTWN5+tPNNj+L9/hQKFo9kW8CMLBZwG0I0rFg4kQPNt2Nzgjvghwho
XGMHlSdlH2ZT1ky862vizTCde0IXqqaNQLfz8I8vOJSdkKsjTM/DwkBn2cM/I0J9
07K/gv0BCyZY9XrvDlkBagVTOY6Hk8YtXZzQTN2KoTPxaNBQE3F0lSanfLcXb3pf
iqv0xtOuym5oCiXVosPbuZQkJC4el6gfdMZmSinD6RkPzvGFEO3ZfZk7uRpfB/Bd
3qI47de7OQrMEjB9KCqiLzEGfE486TpV2J+fnoNlhBGmQbFhELW5+Lswsplm8HyI
NtgD+YKLyZ5CM/afhIMJ38YjRN/UM8QRKxuvpzSvf+VRMZVuh0hhb9zXkdfg2/h0
/Js5HqfdnVn3Uuuy1RYbqo92oxTJYKMp4R2sIGXChYI9oabtUVR/Qo/E2bVCodwR
O6rF2I91RZ5Basd8HdBj1eo66Dt9W+fS4h/UCSfIVGx3C/YmsgRvYp8shu6WcJge
ZNTr2o1FQ4GFcnvreZzY0qoXChT028QnacI3mx1lj9/rtlFYWh5Da6U1/qV6UjCr
xR0CRXu9LMuK7SA4wXGC15uJhy3NjAfRH16oidz13xtC4w+xyFVlzomksBjZylF4
YiC17G7oDDm9v2zn75QUn+9SxZEigDpZCxXRjCYfxZv792h58UFtFRZ6fLMMFh3t
+HfYH14OhEC71yKSGKFuuNB6dGJEzByDG2SFMOnYyFlCH9LxH2a31atqxpn0xBeq
Q/4KSCwJ6VlXt7du+GjtIIhCgUCrI/OVs1g9jD0HNnZSzz+U26NXGcXvP53XsgjS
+HAAVsku4JmrZVhGOEFgy/vp2IjvtCtgxLSfRZmTyn1FCHNyv6egaX2fYqBuKbuZ
R855sqnOCzJmKpOmkCzqnxikSkTAB69uh4cl2amDHc6z7J2S5SBvtZigyocb547b
gLaBG144csU13vimBT+rfF2BtqNjCga8zDiUCt/JAsbHZjyQp0WbM7/1ONgprqTL
gekGlcQbyjx45hYCRPdvvuCaEPvtVZa9U8rMAeuCUhMY1auLxuH4hpyQw9+/Ia8q
iXOVX75KCg1WIi9htF2NyK4e0+ADvIT/69n2Ndd5mdCyWoPUz6zZBsKUB+jpP8t+
LjR7FMgtEqLvBsRkTAUg6NzgKShrTFrQhDttfh+jla1LokQxJGkP7508ewsjAHz7
njeDZI98R6Rxpa5DtKgd8qVijT0etG+6RRvN7tRgBiE1lAraF3cLx7w8YxBzByjI
nN6aoxW54Wn+sImYS3J/eb2i4IV4rERt9PLblKHjsM0C6NJBK306gZWwFcgZ/WJH
PSPMCya+NQe8WnxQSfw4LcLo3S7LiCdev7Do4xfUKv40FWtW4EOmNuJ4hXAIPXaY
DpkSnyJHwH33G3a6B1Gdn7fYz950fJH60rbB70rLzFr4cg/8Jrh7U53CiBYAO7jg
8WYr1DGMx5RXIr0RvO9l+QRD6ufbxU9lWVLKe1QLn5abRS3JdAqqM68uys4xihmP
RULMClbxTeoixJMSCFI6sOim7rV5W+u/KmcI4yWVVkG6+jQBN2N43wJzbDynvjmi
nTu0S/93HscOisUao25cNaKIwhUAeRQkc38Cg3IwOL1Jk6ynXlE/wSebTbBloPNO
jb4cBnKopFdG31+3R+QAMZFCVnFt2bfkpCmMgcpvO0IIp7nBLTHc3/5NMSV5AudD
OVyl4wPH2WXRQLBdP/GJ0LUUorjkt2zcB2W4uotTf1+QAhqAs/9B2nUwGQ6KhWOE
cG5Opg0KUhtm6Udt9ZBHdAgATIiGF42aMAteDyKtoCw+gkjE8c7SqWXFciZG3k4N
BGadyHvoBKqDZbzyp9S1rkeUrz2MpXndmRCD8/LD8iDjIYaO7QcnFj+SNYwYDFAg
kAXaZ2z22BGAZ5bFIM9bKQ/uPOQZUBIN3OWbD2zA/weKM0wnyz5VrKEfCHyVB47+
CHwIMxW7Bz1yq1BNndXS8BnuDvz42qnD2ne4grIriW5st0Zsm+osUAMygmtZvsdc
/LCYFUFHJIKKpvfAAC0eMOlfhHQTa1HJA8gWVAAXBV0LE+xQ8k7z/yrx0S3N6Wj5
eBTa/WxmblhCYBvNGq6VWWIlzwrSl9UcPZ9Uah68+lTYl8pUI1+o9GSNeB7l7+L/
rkz6i8GavG6YH+pAOMblog2CgdYQSwL0IJnwG5zz4XYIZ/DpbbxIh/Na5vLC3V3L
U6eF28cOhMG0NOnOQ0FtCEllbfuBH23E69LI+CfZ2a0VehAzWxDMTa6wwHAzdbZU
o2+GHMTHaZviGeeZWPC51apjps8CGOQjP0VKZkQ4MRKuIlp9qD47Rf+fcfYg/jDw
cSMgWpsTYqj4PSrbxK4At2YqlDXPpEG98Vqib0dUcoVOuHW84nSVyANqmk0Fbo8H
tgTWFhkYkmxDpGs3t/4LeKdiWRmafh4t3ZHfIfSSsYNIMRAlJjMZ/fmjI1cUUkJy
3zKpFxlAXzkVMbR5n+qMOWw897Fe1etDEg+OCE/WlaIpBV2aam0nIb+lJll9j71O
6gHr8+HezJ78tAKe2cBSBXQMJUymHCqobpd6qegFForU9FUaitaL6mTH+dV4M02n
6Ca25XlXUX3oevJF/dZdKjjO+MrsyqLlVPPRqZw3YUb6eEXJO1wgahCpD/G6oCfp
EeOKHfjdgeznqTnJlQbaZagZcO0ZDDsEYJkDxBOcXLag81r7XV/VEGUIAwKB9t9E
D4j6gbZtB8yHkfIeRjVMtbg9Td72sFIlWlea+nYElnc89wyEztpNC+PNZr7KEByM
NUl424RMauxPmJWFd4j6DgtPDnxiUsgz/NorsgfgR4vzZt5Vc8OhF287VchZSXFQ
zHKBxfspyavUdSMWHc9vgrwKiBxdbieHoXiyEA1ErH88cVBQHWWzGJ8KB8uLjm2D
GoPY8W+bDeHD4zgTyYlV9V4B6AfV9WCAisqv3g2b7QScgsAQ0vlA1BmckAYRs30e
Xilj8D1VXlomzGYVUoFmYTYCWkHKg+PHu/8COC3fNKO/ksrgJuLme08ouMjMUuNB
sMZKMmKFN/NPYrqf6Nm2Uu0QAJ77nMjknCyQAoFlI8tRomNXT1w1rP3a6NSz0Gym
vGkYVyqUWy/F1zVKPQxFwNcmtfLMcsHfJtMf6cxAC/ukO74m5X7T1KkqeB78U6TS
VQao7iXGZqK8U7HTB0Mb9VXf7KKJ+8UsMsNSRPmmoFae7bIMGVjxuAawgB2tBD0L
kgzX4wmbOpaoVL15NiVJOJSRMIPAjX6BbzXamoY20u6t/i934i6F7Y5849/M9FvO
MGDlk2o7Bu5r+HhmLkJks9yFZnMEbtbNjgMGi1nhl5F/CvgshkunMqL5xC883kzm
nsoOC6w9uaSRF4OFrvNtmyFL7G9CCYAtO6tge+aGTW3LB2T/hk4QZqtRGqlXMdtb
p2EQaDwYe0yHOras/bZGEQ6em1cDWAclo22DxikymYRynUl3sytRJHDOzOr7vaLa
TytAv62Tbw3N6VeXlvINoH378EijYv90R9MIVwe0a5JrE2XwuLeBf7x7PonWvcYw
A4e/Y4sQiunqd+Ox9F4BQtOkcF8Dbw567blSlMQUJRttLWC1F76O3Z9HBDGRevVE
cArkxZV03IWAgixUnWuL1JeSXun/xg+z/Ol2Gh1UrxzLKFtU7qnNAo8PaysvReUn
NacmjaizQvNYAk4WqiOy9T9t9gbZOAMUAkh8PnlFTu6ErZ/x8riQ9q5OMiaFuO8Z
VHrMGwI7lY34j1FfSlfU1A1Rn8uGcVLc61yaJAA+gl9CCi4tEKOS/zxHsYWOwe48
HB1gaK47e3BfT0oSsOsQj9C6FtYMLVQSxCjzrIxRlZgasUlsrgk4HbSUqPBqudv6
eniJhk+fFxbabzhxwP6vMuHoa0dWcEEnPwxROhjn3Us0eRLcqVpj/XIxQj6789yx
URKQJZtc67BgRkNUHreSMel5susg5cnVFfPa75XPuFUilZjojsRgTmKykHsDQDpC
RpTiPalqwLyCbcmO0E0Zit9DnzUPKJ8aL87Q61PEeNTSe3M92D3/rfHUWEgmQJ01
U1jylcQChZJ0O19ZCiYA9myPJrImpcPygvG98rajPxVU0/X8GzED787aa3j9zS1N
eXYf3BUlKcnUrEwgiP5C9P3WmaRL/hktIwJfx/qkCqdjw+atlJ6GKptT+2DVxSho
qj6LKrqGnpOr2hhUCUDl+VD9kNG09NXaliXjowXhQObDJQQI9gMr/QwdMkMKU9Yf
LJa8oQmZ2PYYL9XrSVq1KzdPWKYud/93o46PgmVKIUDQswzPRuOrWhrz/65ezPWW
HInAbQUHYYwRT3l9g1nSOYVf8t8hNw+NfEr/AZSEUcHxgl4jGmFFqcdSGt8EGTRW
VRxBoLJuqGU62mu+Ndbh25fNtzzQauSXDETRCPcxuk/sGitTN9c2zEvQ2TGUCl6m
OGiHNyd7vlFiUALjNWV1DYgDEmmfH+awvDw2DU9gHMpVmmnn9Fzq0H8kIpb6Qrvg
v//OEqnJ7ef3iSohwu2pfaPmAsPtKjtJCg5Cp9LDnWxNLptt8cv5XWq6t7vfW+3g
x5KNNf20e3R+jmt7bjhdY6INzbzuNASVXvV2Md4GNJgpw5TPB8Gb0zHIHf+/9eGn
/2/v37K/H7n/YLd6zkTberfMLSdfDMjT9PmStVshnl5jEvxYVBd2WzZsfQi2ycqi
6Ih6YEJocULAS7XOSZDIjNZ+gwisfBe6qUhJv1pzTJwFOVFFicEojOQnfAvrkQsW
vufBvzOvJcdaToNFtSBkw+KGwgln3/EAJHo9cZc9U/KIfEAtW1oXdUDKBAEjfVy4
bWHsmk2JLnP9Gml88o5eYN/QJydy3S8REBC/yuO+/OlW7XrYnOE9T2gRpwgXrxaU
I0kysnkvuQio9cjnJJwif2YaM9JuvZfuduWFxNaPHzWpYGFjHpPJJ5ojcqoMroLR
MFgOb9mQGJ4bL/I0amkktQDfq6P6IBGwpgkgovQg/JU3RQPkN8x4HGzypMKCtpiZ
7BL1UkcKkwCzQDQRR9MADIpQWCbJWrm9VXBcy0tngbHrTXfhWxH481AUJuzpJeFl
QGeWPuJhadXDFRmAjDJwf+pxZOaqdftDfjO54lyY9bIMhkdjYsE+y3oLebezArQq
mJ7faNgvgx/AQML9xNWwfFKiTZBEZaJwc/rv7hc+ppTN4xu1rZPmVZD+Qfi5dLzu
W8PkJI4BUtSs39NqhTMfv8oos8FVC49tY+CyDm24Au9+S5+Qa2aoRx31diUDT6Im
k3eALZQG+YVLSeIRRZXRK4DmiRFvl7H7Sa6jKUKDJ5KIFucBVSK2iKIr5sr8lMkN
NYW9vL/YbJx4Tle1Q/2MqiBFWsT3BVHyet4134GHFrhHjah3g2tdZvc1ftyvTIMo
YPzETsVXwtGYnpscFIQJtyfqDRswuAkKs7EzlAZ1+WELdaL18XEznrNdRR46EhIr
GYWESrqn2slv/CuaoIEU/C8a6PlABSdDjL3wm2Nui109Kl5gvRTXNszs8brNsr2D
6LHyC7drZzhTJ/41PIG/JGR6uAUKkxEoEVEpBosE0t/nZqwHkI9fdPtOQ6GYNWbD
sajVwH8w701zu6FjmkL6aM3yPSXdiXTg0X+BhT4//ZAH54MS/FqO21Fb0o7y+xmz
n8bKCw9YAy3Mvw4uH0V05npJddQymlxIeY7yefTjNGvTaqy8Pgczfln4gU27ZHeS
HSFhDRyxHx/25qA6yqVZSCYcLzI+icF9Kwas1yhRu2qp5X7tBa9vXwQ0PEoaoQPG
mWisk99TXrv8J5OC6kzkEQxGQBMA9CBQSa7tfmDSj4pTrsPCGJfrA6YEO61naRqQ
QPFBZmwP7/LPbTY+eC0b6E8nvmrxMJ6dl3hK90OYpWWWVydCB3xfjCAVeJan6ciG
l6OgRtgUFAGQlfd8YuqBHoDIZRx9gMz+Bdo1rwrCMl/ov3wn1By1QmYIFwfdMjFy
IEDltfRQT3ZVshz3gZ96ONsL41OVdzfuYTutk6VLuGT2H86lDvl8izIz/U6WpOuw
Gerz4Hc2xNn975rQMqezd4M0zv6J8w37iISAzy27MUaIm5biFTkk8smg5EOCzqzW
HynNgK8dt9F4I6J+GbmhJhJmIrAjlx2AP1YQkZiyGqpzTuTqyKFnQmSaWOSq/Inm
ZxGeGk8enUHZaZoa4RocZnC9hkWbf+/LH2rmHPskQrGxv6M5VkZ9B/u9//Vc+uyz
dbav6WECZhNNhTQfItA/aByi/SVqDhQvoFdKtLVARsHHKAJW67DI++az3djO2zbU
4uQYv2LsjNALNnlwieC2sqpWbSZ3fL8y1CqUwYSnEkOM55OeNZJas5ePwBf2SAAF
mZOaShM7UXDTsxANKX9SbTvbqijPK4foVcbpgaUrw0ySpj1pUJzN+libQVLw8eQr
gIGI2D7py2mWiKCjm92K3oiwJmXwYpDocx1YmgGJ9QVqchH3pu3EfUQPJs5oyyDk
bBdJK7SpBVz61GxX1kfaqzNv+m9qiy1g+d6sqoEnFn8sePr4P8YpWccCix8XImjh
7l1Fu+rwsGo4mZd26En8/kfix41i8ELNM4Tz1GZ5J9t4GapOfQv90CArSMEHrcjM
snnlzi9TASZP9vIPPhfefcGtbG7a7WFmZeHjU+rObuA50ZhzS+i5f2o8YOu3FXHX
LI8cv7fGviGD78OyFxRsHMOhvVNG2Ne8Xp45+t+t61qHaaon8XgDmLmrwQEr8RHT
4B4en/x7T8+riOOR4FgpuGvsuzaK2Fp5IifuEGxbO094jWe0PcnIgKPHyN/t5st3
pVgQpbeIwyZ49DzOzizOJq4EmpxNKfn6+39n1hM4Y8EW51tQjm4a0J/bPVjb1DRm
j8WVrk+siY+8bU/iDtKMRqGO1g8UBh/7zwx3dgJ+eI+XMKaG6bVnH5eZJCrKWu6Q
XXfc0QRKO6V7Peutpha6pYkYTQMTtxxM+NzwKny1ytIEg/wA1iFnV6nXfhB/if4z
FJEJiJ/YVHQH9PhKb9INIQNHw0d9MiJ/jfHQcO9cMDEl8L6JPBCrzlRgeHS/GVQJ
/yADbyQOErthmuTK+Qan9JbZ7slkvi5TCwt4rJyY7OWOP2Cz9RMD8Py+Sy5tA6Vr
aW1RJuj7gvD6PhQQZjGasxsY5LANi7syYTIA2A+yp0fbPbudhPImflZszU8aMcBn
1QbjjSpccj2Fc2t3MqaPnc+wLMTgVmProIEi/ZYtAUzTYrkw/hMPPAs7LTvZYQeA
hEqYuNDGbjQtFk71CQAO3DgtWN1NaQbz1iC5LaGQnUPfJdRiIIxJmftiXS0TDm8m
1B+PUvcLtK3UGTbNCQEt8wK/On4D/w8ZVOLYi9ZCz6uuNTDbLdO0fHOMO///PmIb
cDl9r9UCOxS0fHnPDoSF7RGMrlXf+UHi8ckttpa1dgEbHxzcd1Wf0HSyBhbTt1QK
gYJRVJSe4citr84LoRVW5kHvWterHoWhxXVVyZeLdfzuJx8v9Pa8aWmkQNStsPVp
BLU7bSTCcfQKsNzwVfeFGL0kmOjsOfuEATgM0e23Ck9rm85RrN+pS0/rMmBARbKu
SNuu//hYpHP7QOgB8dIS2NtinAlVlt87IOQ8uirwErmP+GSE4bzHPZmf12mKQbYs
5Br+IWexLsy9nJIXmOMTJav5kv3whvrDAYB2Lql/IVPFuPhETQ56z/fMee3aXz8h
yG8fi67SB1FPIVOq/hXoPhbaHOM9RqhBPfvuBLfqtNwfqH1mtWqPral+pYmKrB33
7jQ/a8MI3b5vTtMHJRAyG6cLFJt5TCDtOPF3FUI4RrieEjGyatpB8GfSlOuCMiyn
miuHicFFeyR+VrSaxNONWiMGLEslvr4Uf2wTPRa1jsMq+RYc08kG7FHa1ZNiOKzi
LBDipkDz9ynclFPhmdgxsWuwMkSKf2dSu5kjzON1lABBCEtwoWlrTaREICPrg3YM
l/8qbcox9qJYXTYOQ0LNX3he/pxVF5JY7FUmNKf868j/4j5GgRfv+OCTG7F9iyku
8FpVTQaGFxx8+M5U8fRQFVjKlT42dY/2ss6ObUnZxZnKGMlcUBeCuvJTJZfyNQCx
aFpFBzdrfXMmnRUUN5YvA1AVd8tDLr9B872ptYCWz+2DDAHqn/BrHUIECUq9g2+n
p3Sq3efIUPOo19H3AL9UDn5KoBsU95QTc0PKuwT1uPRgIO8pCA+1yDu8fmbRLMuo
BeE0lO+sxE0r/8WoQXhaJMBzWznlBF9Gj3EO4Fw1v4d9hCbBgoloj15st64WMcwh
h30kUnwsZeT0CYN6KTP0tfUcJZRvvo+D6OGdrhByITYSuPBj1j81AtCg24SVpS8D
QaZJBJhNurvaSEDvXxFl9hEyB3Wc2BgK684l3KZor5hkJKdXaqOr/lVxFEoaAwuA
qDnCUFbsOcc3sFfsu+CyWWds3GY6R87ic12mfzGNXPTms0JGhmZ5rwA5XAMDFieS
7bToQgxlslCqKfEmXFm2aS82NMuTbq1GrMA1xLq435MLRc65X7O71iILCRdyR5UA
TdtehNkao6JYzIIuNhFVhtjZlfI6fAF2RPEVrT8HZ1knDRpsu+EBY2dCQ4D/ZuNu
VL1jN/yKRK5RNop0Va6Px28u1XoTfV2pLjFFX0DY/Q5QSXT7uuIzanful4+B7uGe
4J+gw7/UW/oe/ThScbClTVesf116Ul2eesmoujVosMSQ8KXgcIqsekl4Jc7vL8GC
HYPPDg6K2JIeRNu0rksSEC1/d8piRFSJbIwfgnPH4kflZXCwzermlwtuh4deJlTD
dMaH1AnFSd9Ki5tDqBkDeehJ6oI2QfsO4sSZMp+NnFUd65i6DhoGovj1wcvP/Pq6
5Q+LBCyK2M24H1YCa15gj/9boj6rBW0KIvLYTxzL7VF0SN2us9UgwuwNrZLhMNBQ
/UluYFvrVDdhDswHhDu0HTH5OkehR68x+IzDRVjch2gs7SLkZuQIkrVfKHplQUdq
gcMi+P+OEDKuyD0cWzdqCGJ4gd8wXndXZpyxrvNaBBa5PAnrBiE8JdSGeeLNZZAD
klRBcKw8UsXXClB6g6CxpLVMrCvLbuoa7pvDMqfIP/2V3PT29oXDd2Z5B+XubFOm
UjYXps2m+A4x0m8FfnSlag==
`protect END_PROTECTED
