`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V648Qsbt6jk7VL5lPZrtP/RaZC2yMNEhsN1mTRHi+ZdRLGgPKI09zd3T24hQho6A
p/LGUgayqzKYnLDZ8pCJR5T3HD4492OFi7e5gRbHNHPcE9CY2LHMYznu4QmGCdbr
3fr54sFtJBZCmhMgArofpc+hw6MKpV6ccRAFPk5MAUHHkJ/D1D1/fXHMZARG7vVn
+X2ONyKaM84WANrBeJwYee0F3aFuigO3bylhwYePnIzIySP5kos4qv3sT/CZ5Hvu
h46lhwDig1DB51MJNtropjqe5JoubADX5GNXW7Vz7+b+nNiYxOqoqpWdlopx76rM
DM/O2ybZKe3hYhhk2fz2/AH3veFM/WK4Ynx+jxsMPcMdunTYwGV/Z0FxtQ8tXIB7
U2F4RpWq4IpzrTFWieucBYxlTWVbCNDXe6ltmCzWKkKpno7zIjAeayCBuuxdLHK9
MmZgoACRT+C0F4wzyVqOeVdmgwIiQRL1YeqGLpobJHJ8RlJayqUD6p7sGPiBygyj
25WDWopLFgDR3RELoNmNXWh7/wuOAlxDhblRg7K+MA+JtZ9XuXdATijTYMn4s/7f
Ita/bC+PzcYy6UasqXritgr52oOe2GFS4JXLzrXVIWS6KW0gKe+Er0PpR67/rjQO
tADap5bYrZfe6orsuuwSPH+9+TnmmhkFOd0UTw738us4CaA5ppgxGoINvC8LxC5O
yWQzCF21JDxPZ4VBRjkJYaHbNi2kjFiwPCtCjoeuOjo=
`protect END_PROTECTED
