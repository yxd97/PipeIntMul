`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h9rjmfa6BSVUr4lqghQZ1MrBm22VqqE0J073di2moJiopUjwK773mIECXENGHeEK
+WOz7Lr37YNt8tgW/wFT608q7hY4cM2K9pv5Xz32M5Jfac0+dvPRAzFRpVLFHIh9
1p1hycIGvTH8HbgVzxGNlkIUYUsKQG+mOdT12bu/WhnFZFJlwfWG+tH7FmzYrzSw
HwbAz0HoHEkIwCS1N0IXXvrRs9Cb9yNGXJEItF8vnp7sYSu4deYBg6kHfSxjuym+
stxpbQt+rSBlYhcZDqp4UWlH/oTzoLb6EGFSX5NH1bIn4ki07ULoXxP8Ba/9NY94
q4ZUqlZGd9W26YRmLfMoFS97kQeZAmiDpF/3Mux+CiisaVjiYbk+XnA/UQyBh1S2
3KltP8quSaxAFo98hRd6j8ulh4CwfBb3zVJTyHQl0tGWJVw6UoqJUmU9Z2BgBBpn
uiT9zpEVR57cyi9sAwEG3xU5kEXkUvOwjD+Hw07Yyt7izO19ccpFLRN35wGruzCD
hCKtUwNyfEkpTZ7plKpVkWo+SiRYo+RUwkbe2WUfb4UVsThnD8FCMlcAEXWSjzK/
SJS+HHHySCkCj4gx0Fi2kWhadCGvBz88QS2K8FLiHzHOTlc5/WJJwXyOvufCDOc4
he/mfvLv2WPfFlLVehhVtBVST4t8VNS5zGxNhrLQq2md2/fZUjyel46KcwZLSN9+
hR4NsA+/GywxooikoAgDOQgGmSd9QZmm4iz9Xs5t7sx6R4Up7RW6w8t59PH2acGc
WPEr8OxyPAv0q8kIFriykxWuNVT4QybdXax7LhmmZ6ymWUamxS2HySHVyhkjByrT
KUaxw0BZGoleUOkNWsCDKILfMF6MlkxDsESnDAY04m6oUtY/1AGMwNSZ9cle20b1
NxMkIiE++RHMJUGVsamlBlOHwoEA5Xc0Fn1+bQ8jTrM30t3Jqygat/nI80ESceg3
pWFQo0gwoiCBaNosSMyQSlPKyG715aAcgorX3AM7Xvwksx4O1oyjg1hVmK4yNAKp
QFj/ce20uJnZLPv7JuhrTn+0r+TrybM5YSIklQFtfsIyFxVChxir3tks4OJGNYIc
h9zQgWy48vJ6+25eY9ZkuS6pIfXfvuK63oAFfy+7gSj1eoejGmxVsaJ9Cik0kySc
Bk9QZwkxauvL/eh5rD1ff6y3xs/tZIbo9DQF4N6/ihMrRe8V2j5DSsus4KPB6n8h
vBJ8LUVNyL1DeGropU2rp+QiQRzkLAcSIP7ASwu1VX4QpUUuXjDZuTHVAvthf8YW
iAVSLEwd1s3Oga4NaZshX3xgkhTS46kPjFZj6iWXHn3bslz4H2WoP4ZcweqovipT
FBqGNVrEB9yJe89ds5XeN0L8r5Y7GtK7ih5/1108wWWrj3J8NYEvAC9T34MEYdAQ
8aCnISGRgfw6HVTjiYby6wqwPZqI0gfac/D+80O7IhRq86KE8cZQoAJ8rhOmkYpB
iPwkmjfvbgIDPCjSelQwjQPNO+zS8yl59GQtiejOPGzmBG7rn6RNqI8+9ubiifXd
59wWER/7MS97Vl42alXJdNpLblc66TlNzGUcn2cvOn/g+EOdimXuZvM92UCPEmN8
ozY1vvtHPY/Z4Rno2F6bUdyWB3WyzRKrCiINCmCr8QhmnaZXXhU5cPc0fbWU6mZM
B89OKh3qXawvAkRLx468wR742IihRcqBBZWL4S6ctjZaI0bu1V0nFNtTYfL70jmz
Ldp5pRfa2ataIe8WnIdVAmURPh9fHOwrEq8iuPUQmJcXigzEYu2gWMUGi9tWAsY1
766vcCvpsnpOwD1sMI/q9pD4rQ1wp5uYSrokU+hNED9ZZ8MfIpVH0Xp3QvCvHALD
AnzaBdNPl0AZeRvxYhHCXURFfwvtQ+WJQc784Gj0XAlfi2MISu92UZVrapaGXx3y
RfkwEckJkgy32V/Zfxg9OnkCFtrhUotChSDmu29FQ1A9Cn5xmzAxAe4fqgMPUi7L
J2htsmluZ1Qi6lzxF2Aen4hmiKe2RyGL7p9XSeRH3w6YcwzVBzBNzwBvUbsPmfhD
8SvvrporUcjgYycS75JLZ+963B5C5ZDV5WMvJ+2NkE5pfGwFWOoUYj/UfqRBozMT
8AL3VV1/ZHbuEN2dquwEVbeacncKE/Geyrqjcr0Sj0/KTmysDg86dC5StdE+a4Yp
1h41smiBWR7/AHWzl7hDAIMQkWQbC32nHeEvk/NB9UCrpbDjnXvinbfQP7i4KNe4
wtXs7zFx0fmrCyDUucNnU4s8zrgE/9TxPeKBaZFwnVyVrpk2VCpNLQdD1tHhv20e
Cu9qUOxK9lLqPV9FxG0BRp0tVe6jiG0tAtCnXZ6ewH3OJPtrvYEYhrU3ccpJDQIC
pH6h+ktbAo6XOWBmuvhL3FVgB3rA+p8VsJ4H4jTrO2b7+S0iRhqlpL6ExaoQMxnz
CSrNztUUy37LSSXXa/LugCm5BbKMfVsH/2vLzbPdLm5Cp0DzeahNuF3kotufTSn+
evgco3up1oRZAjCvQjAawpPeK17KH48UNV6QoZq12z08L8+G4VR8bJ9XTBmHNZbY
3/3a/b0naC9lumXDKrd1882GrYSXDr3kq1ehMDSAngaFAWLFlhUWAjJV8A6Rr8ZR
IJ/vmS3eiArj3Is1hd7iYl803aNV9qEguq/7nRu55i4mDuQ4bacr2OKvNanVXL9n
bpS06XA4hc/SFoJ003btZDhoy/asMbLFJEz1nUydcdtTeoJmOn79tzs4Oojduxfh
Uyxs5/j9OLOHbNuBGKGxZbtsHhXyLtfOAoaBSIL6/gHjm91m/PLBZmSVlSbBk8GH
+M5Q2+9w12FuPqaDjN1dJ1kcvADNig5avY6BbyECb6vTjZZjHeycQMaiaf+miP4X
5zXDU8kLGz84+oEE4b4bm84Kig3JmTkBZWGdiRVCAoiE271W1cC8FPfWQf7JKyjp
pmxK/NTAND0wz5Eu06aA5dMC1HdtXA7rKB+1eERb8QBb87we6/u1dUe3d9X2UC5C
yJtVTuKefLPpK3vHzsJ12alaFZyWhuBFHbRC57Q2ujtSdN7BaLP/L4qxVwKwRbf5
zRaNrDulkQ1hCH0L256NGwJJMUFelHIuQk4ih/aqHjbH54hoiElAyuBaE0vdlS8U
tUx9uu0/56tmcuagsvbqRODWaan9w/ubfxerLYCMq/AKJm5rTwYSe4PAF49Ys+mz
Cg2Vgr83W3N/AfW2p1vC7AfDTF/5TgJ3OQfWvju9bOAgBPom5iBC0+5lqJMzrgb6
VaEPI7i0F4g46a4t90pU7jDoTXnqhva6OEmkBNePeYuHmSv/QtjWKz92WBEINpu3
fE1xF8lv5Zzh8H5LCJmmEt0STfiwGsofV55XeQNZRmEiWClIdOJz+wKs52A5gZZk
sR5VLXFYLt7ECfb13hTHCrvwhviNV3B5TQGISHWlHnIwav0OVgjFKNKHzJsLjXEv
K9iXkE1pHoQWPNYbAHM88K8Fd5OXQ6JjSqMTSQavCDmJBJjWSZ/2gVCQeXQfKurS
+AFueCcqABoLfiTdFCaNUKcDmLNurgGyQyd9w6jhyLkVr8fVUXm8CYq8K13TqiP5
aDhF7z59ur9QvWz3orA7OyRwLKTCdSU+xl7KPIltyURu16Xwh/MO/bnR1NnAA+HZ
hmd+vcvvTk2jJ3OJGmOdKtM6tftprdqD8fAoJMgf2rjfD7zb6rISVHtyWtz34bWq
HdVi7IW58/oBCXh+/W9OK1bwXemxz7U+lt4zDC6AqVLgF6mMv1DIFzJWmA4TjDoX
Jlos+cMo04tTIAOD71ks3ZIUVbrrtknXgwnfKklYUD0dEKnuakZmlfJA2l/s1n31
gtsLECFSU7IR+2ekAOzpA3bE79+JYmo72xJBqQY6KhgQM1tNzL9AkrnJen1IEKUl
TsBps+gQEVr9dw8WMisjCMZFTuppS5fs9zYzSKYp4eZFCod0nDYqvrX9WQkj4q5U
hrmEL8s3ZPUb/dzXiUtoLt+jgyApSnBnAtagww9dBHfq4wmHlpxHfMHX8knmRqRg
76n4X7dBPXanii0PILHmnzKaGnzdRuJJokBgEX9jUblJMd23ugnR6GJfsOZacMQk
/pJAYvHDxIegl3g9KJfDLxzpMThRC+bms8MuJZ9bQnAIc3NkHANHwarURyeiCQ5Z
CfxpnE94c9Kdwbjv8WS5f8cWRZdDxfemOVqcsxOLy9gyXuhIrQXH//5cjNS9PiOm
2GBJTZCdGUo62yFimz85JvjGWoB9hQi/LvyXUibnJLR4+c6jxgm6HBU7UUWDbncD
4xuzNDk2NxGOuhFWUBO0W1jDjTqxQhdBRFZcbJv4wAbuzbK/vHPHsRfTikW19eDX
I635ndHAnme0JzSHMI+mYo7UK8CaLCZVnQ/Z1jZUNByjnkbqBBA3ReTT2ktnPVVx
zIgoA9HLJ31YKmx9y8IuIh6QjX3ZJ9AXdELyTvshvRsMLjRf1bMDktLO2p9MFcRX
BCLDClxMjRMlxPk3AB//pQQ8GfmXU1LOJUYEGdJUfVx5uojZBbgwtnIBHrPHtCS1
02SSU45L4fPFZE16NoL63mIXcxbVMZVKOZL3eKY+0WhCnucDKDxG2xp7dBcc4bV9
DQO3k36H8qSzz8NRoKx9DkXQ+pq/GFIF3xrgYfi4w2Gr6kYfH/NASbfERFChSsYc
IlUUoHBpdZmGMfpR9ubUPr4LU25WtGuYpKmGk8sMuJwO+mpS9gPbDCahp7FIAsGL
nbueoK/qJIfmiAm5HsCDRvQdabi+j6wl2Je3YIrDZEIfsqZLJbhGOP/Irg0MzhzV
qW5GbhhLM5ipbJWY4Z47pHQjrB2Alqt3s3xae25T5RJzcbJXcXFZ8dY0kNUNqkTs
iBHWEhra2irvWJf+BMPyPTW79U53IEr9ibl3Z9vNVBA1dXnzU9sfq/k6SV5txsGF
W/290wUa8i2BEcTYPqfgtFq4Fs1p5IO29EV68zXYm2qcWIaUcl+HaDqDpZpLHfQN
ZpV6mCjB7IMkU/ZA07g4xpdVMTGbSG22giq98c8cAr6icwtxLjqMcKThLcW9H2jV
Tw/CshqEi+PVj+srN9IIaiY3OODD74JyZGSQbtb5ppqm72V3ssBWSuHLoJ49mPPt
DsgQqv2Uxu4ok+zlCyR2vW1jCX3FV7BJdy2ebL0rmjBTxXas6aERXA2dUOoLZ8c4
6vPHInDSMqMhspG/GIL87xM7RIvC3S3NpLPiR2K/310sFm+iv0XR4aJlvALbJlk/
d77o77Kuvo6dNj9iLFRPiRJgvyZEfXyIKp2FTf8+rP0wHokxRxM4uw5p++mNBytS
h8e/EqPMZV4XIu1clTkHQcSFhPHJkISVDqpfcrUDndNu3r6NFbBCkCB16xsEBWtE
SKxIPsfrJD8pUOtciDYzOPcJhn/6ME0ciFKu20zILpThfwrP6kWk8UaOGfjTNNDB
EWaXAD4iYnUXPoqzsx2jBIr1GBC70kAQHjRNP+U9CZJqXQFygXp/O4+9KR6/F1bD
Z2296JdyaFfQiHOuZbZqe1pKiBieRoBEs++SqhEJ7plSr5DOcYUXUWB9Iq09zgcs
8IsjzbbhGT0Fgl7jOYTURP8VNXm8YyQwMDkfgFUVfDSNaWoIF7DreaET9hb58/Lg
HxgDx/zqQ9i8ctDXDdolJQB9vWYNGsmqvAR8eiXHjlovtkuPzjUe/80U8pPp4qYw
FuXkeKBsJoxXz1e77IQxDbQA/x45+C04tccDHLmqaioShxMBDqi7wbUY7SjOqBMa
YYkVRqCSAfM95HtuuAix11jd9C8aajTjf9zAkURpeafNRxhdO0qw3vhRHYpZWTrC
FVi7XPeMVwjROFLJYoQaRqtbyq6yNprpJRBaravgKYMi2gkRA8PzGCyxUivJx9gg
3xD4vCJ3KltN3H6MO3gi/3cB3E2QUjowU3ez+cmM9ciZKup+ykz5E+PL3fUGfkMf
62EvAgFTqIHGji5x8USQ0hH4MZF6QaX90Ck1QaCSIX32E8VeZL9DNE8gn6VZFghd
hVsdXS6FPq30B9BL0TY3L61wYYsqce44bc6PA7ROSeHNtL1Sik/ryLkjPLl+oC/T
kGq8yOoFxc7xNiwBl/7S7DMmOBgpFfMPRbG6X1qUKftqVArQAdKV1ucxK5zUFPAU
aM1AM+3usIDHlabdcEXw8nxIix2Ij3/d3WPIh3PqHoY9CEDTTRO4Uhs0rsoYhsbW
HZ7N5NFNAlks/a+EV+EvhaumYxmq9tfkzxqboFG+pdO8znqWqwzTu9DCBDLio6n+
rCwIRHyfRO3aMm+QTgN77dEkSnsaBXi7rkHwZ68lcCwyCfwqQVP2gFgAD9cckol8
oxAdQ9AhH4u2UJYSVMYL51DNppqhygH3CUIa6yyKA+ptzl/bHaR4O86oArIEpVsR
2OXzB1t7FXxzIWXi2wRw5wPZmxEnH7nV6JB3/l40m/2Tv3+z13/0HGBD3auV+jvA
Fk3NW49dDH13/b06WwmlzT4Ldn/ErA1132IvjpHyEq7n7hkJoZiI0BizYKq45atd
AdFSx1JZ7Wsmo6DJAzFc7tBh8gI39EqAePQZgS3p9/1PwB0OvafvBxccLZxpSxOm
VjYBlggm8Vbeosh+Hs3zo9t1HYB4ZY635xut7ziXZPUraRiJkjl2pN3C83Evcrb0
AbtIRZrA9AEFaq+XGOnOKysf/EedjxTX/k5IYISYKCsfEmgWyO6YZZzy/QjTMOq/
+44VKfzbrUrbgWj6RTtDnY05jRlONZT4WpvFMeQp6J8P9AXIWxENWNszWlVc1JXg
ojnQ+vP0jUrL25hp0QUEtDV7lW8LMAOPcv795G5pRhmwN+LJ4JQ/etWVEvYSy9cD
KDgU9qGYvGoW32hJH3OeA46bxMBK7yYjQL5IzVS1r+fisi/7YfYK0iUkK0yKWPil
/zdO0a8Sq/tIUIySCskcHvwld/6KSRwl2HUFvSThUlHPdBuUZEEuzaUIKo4dosOG
mWuOujO0AgHyDzU3VcKfNuFvA2J0WYQIAGBzGxq7/9v7pUR4MjmMY6a/12q2dBdw
ukNhkhxY8kL3NZ1FWeqO/pg4ThEESanLcqP92H4cmUlOxghuAHdtQOiDfObF6IbC
FsA0p3GFJ0ohqUta5Ds1NNZA2kIL1HIC0TcLPmW5jj3w82hoIXxw2f+ch8v8rT+9
fb3Jz+VzFA22Bde9amTWTbstMqv0IVbsQWwRWrR8rwjp7LUICFBGTyf0RaLr/moF
31BcRC9G6yBNi9/xawl6Y1Pc4iiP5Fr3B2q2kbsGzSk+t/M/JtG3rx7A4hoqHUrs
fLVIyuwGHxxlpCYV/qdtzTHFiQHFSbR5N7SSVzeTLOWK6vuaknF4KxlPvM/qq50Z
LV++eJmOwP74J2uODj7kkj18BpofhxGlh1JMsVMmMFpn7260YYv5S4TcrqHnAxcE
NCz3h+YzQDUuEE5ty1aNGpoXSYxieA5WETynkfP3/w5G//W5SWfYFtAX9kklASwT
dRvUDitzX7ezzAnLH6xiZycnhN4tiPvsmRQn9ZVJnAP5ZFWZgEw8gqE5+wZ1IKNb
MNu4EWlgzXGC+FEkyZSfqduPNSBedihIsO5sdC4eohlCRcr3D21+vv/lCyt4/ShR
UeucCYqFyNYMeJbNRhrtNscSCNM8aE9UBAvsNVuy3wfScMMhAzLCUlm62jCHIhZI
Ql8F2u6SMVbIUr9Fnx5s1vl/QAjVDWE/iZCLCfJ4G2+JeF2iug/b6YRTNum1M7cw
H5nCGnX/OCxYIffYhn1mVrkCcjZs9K9AunhT9ooy8vGEhl1H9Vi0feKDNYaf0iX3
w/6oHEyw4eiJisaZxieggkwKGktkVUK9XjGKv5AhxWPmrQ/C0jCCwcgeVFKyv/Cf
J8ajPKmk7wqxFdZ3cjUc+AqI+FmxD0JMLDgX5tNcktm6u2f++MK5dIaE3HEcIHxt
GgUgsJTaL/vJGvdahJc3AjRpUVoqGkSYqojMhiq0zrpFqcMLiKhsP8nEnLpv3kh3
i+nCRhY6ML/u2xIYpSMexb4atHdW++SX6KzJVOiEpw8ainCRCLLRkCUMUJ1Vd4ys
uSKZPi1WPFyiLJW+4Lz2Q5cFheDtpz2t9vhJ+cg0WlA9aICijTwoSOZVr+QcNpIK
Wsj4tMLFV/4rFtHJVksAa90wr4yDo9GElPpBlNROOoZCtCTMdFjPRR0UXWiN60uo
ll8gXhFcKHp88bbasInUx+RiaBCzPoS67ojwn3svkFxE7FfuDBeZwKc+VtuFYVYa
USQYDoO9HY6cNRP/oNEj/Elm6u7rlzqGnIj0BBp01H2OtNqAWVWDiiYJe4nk/YcU
g/yxPl0OLhAEGm48uSDNUcSvQHHQqrE511ErIxA2W+V087c+L6UmLu/7qVQEDJZH
NuVlS6ldfNazLyHrnvv7kSfUyIgj34zpu7OwCADGq0vq0/S6S1yU8GJvMrO2h9ln
MCB4ZTRIANZsj1yWazA1FgaOHmlXyK8JEzScoNjwxyxFrQ2Et2JcwICnszetKdP7
WW/tK/SxheYZ6iFTPPJEemtATJqEbpxgOHUJdp7JXEQmOgknH63OjXqgYlDxKotG
IErOxdFycdFrfoEq3tbICX/DEjwjEs+OUger5hIpfB5N6ANZG9yqSkeR5U4NNU0r
RBNGGsVzVt5k2SnAnKL6LveCNtZlz9L1J4iSWxrOm+pouInCHHBvrZaQfUbJC3t1
K9smHsLf7LxnMuheJSOk4xDJQOZQzHZNvAcOhShQIcWY/jZ0Y8M6L3Xc6UVM3vNd
9RABYD2QgmLOCUNmHkMc7khA9YQSJ09YdOtcB4iPcHv/bXZ4duQzFYkWeOz1PkwH
yxWCBjMpSFq6F4Jd0DoSK/giEGaOtYd6R4oojaC2RmkKXLOTNDV5qAIwb4/IMoVh
THb0bFQSFi7UWD3dfA+j3MpryPyv6m8aOGzPtN6dWigV+vrfXBQgMA9fHa6RuHuJ
ZiI0fLIz04+3NyGbh9BPs/nJjRbTcN4SQewgK0xhFfkswptpak7z8evgubzQJ9uk
8x1rHNa9b4OsRJIEV82z6U+Qn5Bme5IC91oNRd6MusgnXuxnDj3ajgLPLXrR+kYy
rMlP7rl4C7ZawiaJ0bRlWTWSBSqNZZrBJ0cxgoEvDjeszlcjyWHB8W2YdJIiU1yY
feGMbdz+IQ1ZewiGTKw92vxaNMuO+Mhg5qWNJzbB6X1aYb1gExF1lE5l4meY1wiJ
Bk0vSqgLB/MgTwtQq4fMimrYS5pXLqvEMrXCPDEIqacIcXwitTg2cGrpzpKMEmQ5
vTztdiPLe2jWXgwRSf+U5KjKelRjdujwy7dV9go+Ptl/lickOde9qzUCRQtZDhQM
b5DUCaanIBX5Onzzymi8m8uO1eZv+Z4j47VHoBm5LE239J26AQPNUusJWPMDvSvw
j1ToesW43oxjuoqdlg+mmBc4Q+sU3MzjHCcPnb8PHVMWcob6B5ZZs3/ByNBy4tBb
2Sr1rhmoo8eVMbsUqSRI62RxMkt1oND98XrNCMrnEjONK4dmEk2D7wiZ7tgHCQqp
V3ZBXRLkwHMTiKna2mTdhVHeEz9KNmQ4hiMp6TA5xsR9zmi4u+TNm1cy/6f66c1k
WllpyKXDitCw8yRth4w4fVcRWGR2Lr7PUhaT8cTnhJmOLZniFqsWPU6x3Ao3Aa72
epgZSWSPq7uP1POBiyug7DZmU3FWjPXdTpL/4V6tiM5jEuCW1d8OQ13YLBp8rpVU
qjSt8Z4tDPFKqMf8IE57sgRf7E0H+XdCiGrQRJH1pKJrkSwKnxOJXchBPW9PXvn3
sbqffbPmOAkMVzMGrA+1QzSv2kOHk/KtD33VhzioNmxVXZ5ZgHGcEcBe1X/Guy3p
3D8wdAPqODstL481lKcfDDXCGdSfn1pecmQoRYR2IDmlxZDD8IOtj+6HCqPHW/qB
G2CpWXaqwdDoEqs422wO82mzCqPtwSHsrv+T4vba6bnOy0aer2iSNuZM5yrO4aDE
8LL7vAjtib7V9L8SNKzmHqDplQz4+yW3s4aNN+RIR6sD92SqIsTyvo6ZlbinBdcE
2pIZ9/n4xvkeFI00Zbmf7nw5OZwMIHESqKpwoJuR4NYo0w5+pSMmSaBLRSSdkiki
xiS8897ZBI2Uju3xYyNeB+iSi7BQCTwkhRxMeMUsMVDpgQu5AdKRQu/j31Dd7fxZ
crI6SwIgIgZV+gQzwi4BDoi4baOTErW4zDUMhKN2m4PqlXQfM7kau1CtFULbXrqi
eqRtyj14HFnahu/yhGlGdL2pq9kRVAi79qsDlGk3sPozYWnYQ6YsVujEMEy7qgpa
GdiV/KUOp0Z31awjAe6DvGXlmvRL8hF5Rtq2mMHU7DHG+EotHHAYsLlvyS4gjrHD
xLKft5Ce4ViX/3UkPZHHg2nKJ9HWQ4GAFhUvgL3uxpRx3UpSPKOcB5zY1jXUm0jM
SCKuDSo/JejHplLOpwJTZYnAWzbXylOIJN71YGpj91O7iyhekTFTDhbcsCJ7+ZzE
Q3GIQfLjaQVnWdOMz5jA9N+itUCgOoKYGn5XUsMR+aivcTT8gXwQdryZfVka7Nrt
2Jj9xsaCpE7iN01UFt37wZY52CNPmQRQbXW8L+ULOt94JpNaw15AYeNN147lUiJ5
Nl3WUnn5GWljXAdDGfg1Pix3qu0k9jN/YZklbTcxNHdb1UVIm0EHW+SM+i+2QHDR
J3YLHM8eNgevd4KLvBK7DrreneadtdF4S4HHr6XYhwKEdhtPmuVDey82/1H+X6SK
RUNzye5UhNxuv32idflQa8ALoaNW9NZVGPrC98W8NbeQCQAmmY0WnTPmmbvOAZLE
uRrfG3vpG6l46HF21mMVGnSwAkf7HUE40povxOc3v9hzR9GhqBBfPZ1O1qf6QDip
1CxTzK5lMzwusGTEIGgTVr3oB3b7SMvqV98JHNB2yZo9BtC+iH1wxA9LjPZ3RN57
2vzLwbhK8CAl4tebPYOfy50fLN7/Rx1CczPF7BGfcMVOJlhbdhUToWZLkHTnVkIQ
ulSFKFAF5ZzI2nTvae+4b4AKcPInZeSxOXgYvnf/CYcKnGV6NsKJECJGbkeNIe/w
ChfBgOLnFECCPbFuRxUE3sJiNtXux9y8hlct5jCqRIxbDJt5F4pjPdevv8eHSLz4
GgWjO6TK6+WsVqweZ/FesqNS/Vz2H3KliTbp/RweiKP1/9EUsXb4XZe4EBg5SE6u
VkWOfl/l7IiUz/tDOYtOofrPUV4p9lIxSMcZ8CWZKxk7FmpOGWwK9SiBTjSuF9qC
oD7pqGGDz1oXFCImaH51warWpEAztDsscNt5XlmnsqPPZ+/ZF2hGs6Cukyx6AqRl
qCkRbwqR02r5uw7WQcqdbVCVFKmsDmi9mS40Gvgoq0mEZbQiZ226s/d7rLj2E59l
ecsGmBaVS+VAoAi9Nmc1NUGGh13W1CCpEcLvXh3qVuBk7BtsZy/ifiaNUohkDbbU
tmu/CotLDGdo6+Ty4YkJ3sVttJHgXvdG1/E57KJM8SLFEEztrRwqy/7ZT3KtIuAc
9TPV2wWbEGIR5grSbjwoe4SNJIP8CSFswA9T9iWTmRBCZWXPutBLIjd8SOVGlD38
d2GJ3catz+h+VYf0bXxbKrAsJueA0EdR2RcBui/hhmF9DCs1GBO61fDizxXZwALK
RqxI+BrMF/LzlCtP9AgnwoshMoqO9DicckLfws+SbsmOZlP8ip+hFx3qRpRtiNyU
RYB2vnMvJNyD9qxRhHHIH70iLB0lVgaRQLsKUnEgQsAqQ3nazbycEPnm4aEI+PGk
R5M1nPbQdox1ckjbYG8rhTgAF+WFxfsYis/Few8ROw3cl/qFHPUBay9KSSe2IYy2
2kVp3U0X80wspDZyVOUItXJ9SgjYF2WEgmdqTIATmxos7gfTYMFiCDTzWKanMW0C
rQaCVh0GmvgUwL0bGIs+AWISd9m712st+D6Qad9DO29XZQZp9NBnn0pSu4H4QVVI
TimCyLo4oFcZ+AuTdjW60+BIAB8BQ4gmtvktP6UPQR8cIOokNwACNN7HQKjI327H
91QwkA54bruk4lIyK1Af0k5HNrhyls4fQXM/Wkke2ORZRaMgGk8RorMnh15hpP7x
kTN4P9T7VlljW0v3RMOQLJbCvk95wrPUJIMU5pgROpTMbVwbyglkADgI0TT/xs4y
xZTCufptbB+SrOCoiTPumQ9Nie62r2VB7bpbs927A5sjoAbOnQ0bDqw0oDRZE5Il
ishNS16czd2C98DBNVAGXycp4jmQCNjNejARHgrQiDhlBFd+lU+Z8R4UyNc3OG2h
oam90KJgDFC/SwihRqu2TjxD/yu9vmplOTYTKs/4sI7JJAKVeZ6N8kB3B9inm47u
GeOEF2ftqJ/b0yjyGGxT6Ww/NUYhjxPWX7obSvAVoYxmRE8DtzJ2syBcx2P4Sn0L
V+cKbvO/R/N+4dcUpEsYGqLD/JjHz6IR1riRJ+XWnEtc1r142b6zhjs4Q3tqv/Kw
j6uSWEHGzE8t0vdRFTDR22BI482RRw8BmsDMKDcFEGo6P4AHL8Ef1uYMbPBcy3pf
YBEyZ3jw0tpQjcLwPpmKObnpOWpzORouvfiQMyRfzB/IOw8jR2ocvGeR6lQlDS5v
SntWK9zvMqTVOL4e05TtsgUH1fkjFxZtbBr3C71JKe6brlSeJR3Hm+DeCBQXFZOS
VgcoYOnoNz/kC8EgNeIPGP9hOLMclFMqF1C2vGU5UX61qJUY0hDkcMj+qjI8Egl3
V4xv0y/iyDm13gab7AJU1Fc7JslnzNWAGJjVy/9sU23kYEClRkn1TQYwxS3EaW0j
Zr+cVEHKRdiDDv8CmQjOy9tFPMPtJPC21GxFL9D5hWnJ4vU0CVTiLl5Fz96VoQ5j
YjlKQKimkduxfAuCzkSRH8aa+INMk2VgKJSaYv/PtD+nA6R1se4pRijimZ4TeaIt
G7y1fSc2JY3NH8+GR5cHjQraTlFN1NJ0Uos9ehwgMbZeVwZ9O1vRrIDU9OBfX3rp
FBjezBKGfnQqY0FCP06sl5dDyAzV7ZEXI4KIRLJEVszv9Rh65Ay6OPSp4qUtn9Si
BekXJ1/3yrKfB1hZ9feQpMpxvalLESQrGfJNOHA5zz4gHBno6q3YdwXZfZFoagKJ
gfwB/3QSN/uBL0+pPZi+tT8CsAcncHCGK93ybMJlI79hnXfbt9tGJgWp9d9ksD2l
mucK5EnNl7K0yUX7WRocwihi3GMqZh0PNwwpWtYYpW/xGGwlV1LuwvLAh5xodE++
f66wY74OVtXAkYxKvAY9lM+ff1jKCtHG2PwOOtU0/vw7TZ2vEG+ypzYHFrBO9/Nw
TVBrzBgJiXY1zjtVzx4gBco8v0fxL2A09ImEXNb90O6jL7+gbbZkH+IRbmCk+8Ms
yJIga9n1U9lfSv5XC9mULTCpMKW0kbsTYhh7RYpo2eYxzMSZuqURgyFeNGDRS3GZ
GZ4DtJPbnMl/xSSTS6F8DE585AwzUm5VE6nlgp1eclnyMBrLi7HcshNhiqEcfpit
ynVaL97MqPVjb57OUK3q5O/+ly/dpxRI+ojh95Rw+/Chjr+ECURi31ssgfq7/val
zFGQf5OtBGVefAk3melqKoY69fsODe0/qeIS5RV4qx9YsfAoZHOVs8C4dMx/4l3J
YC0brlercymljoJTwI2kRqmyXbs7QC5XsarTy8ei35H/YhBCTJkcGWF46VUTc3Zr
YWto9vPD6jOzojgtfMUYcRMN3JuNMVuFQyKK6j9som1cGfylE65bkCaV46YL4LU1
6Dm9edcdzOUoDfhDXL4a4XbL/rR+FykJZzOFAM4fntK27VNPlrZkLlZzygAUrHfd
/C7oU3yjrQjv1Afb0C8IcffZquFcRi/4imf7tbj1aL5PcOtMDuWhguDsk43sGGfH
sgA+U7Cm1Rttz+JAARGD88bPmkqO9gOzWYSYYm1U67TM3wXTH4tS9n119vLROkhy
Lp9IyHf7Ca71QROb7ofX7CmrvUHZbU4rF9FnDbDq43J3F0R7BzzQVpyZsM5csbb7
yskmNmi16/qJ8fuxrCY1cBqLVEECBJCA4cqEQ136tHng5g6lezzXqHsoSqyjNWOD
P1lnKYZ0k8j8BaKfcwJ4DHeTB7oaJRekfDbZypDGInA465hYaqV/OhEDzyzxD1zu
uPOAKsEwDbtViqOLHdvL6nrJk2kv3AZZharHYJ9UqL9h5shKt8DJAl2uUT16uTpB
Yr5u4/7HJU+5qmOPdteRcokBeh9vW+jmJzLVbfJ6fM7KUaFkN6bHH4jHkc0gWHCj
q7ErdF9iYNIcarBZRc6Po+C12KbDgd3WXLr2jCE5C84lkCeZrNVS7mydmDzwUsfa
ZT5uj6vMHowzpL6NnG7XBR/EK0y2VGljZ1eoWq5I9HEpsjHHzF5uW3tHCH4zZCGz
gyzg0xs6bhgfkkIfAN8r/idV9yeaxS4xXLrnSbdYejAS44k62yYbzDJojtNWbmZN
062aYK5mUCQG+76P4bPR1JrK9QAC1UTyxmiQzrqpdnKEBCc446cQbN6fCHHrAa5P
ZBnHyuzDAcF1SYoHy5ysGUkSba6DcYxqzBNIQuFPrZKxiUvFjWoP+/Ww2qSRB5aT
9AXHHilWBWlLB9tiZykG43nr3O+Bk+TjMV4qX2yvHMl5eG2Q7GmWi99P6nBOMtFG
fpsRb1UKFxauFUChsEIJzJedhTZss994OoRbKfqzc4R0hWJSrYBLVZC97AC/Ni2p
jv4Iyqb0dE+y48W/f/7eBXAbnfRD2lI4eXuZGU9bYTJv/JFawdbCPlN7babRHdlj
K1VB7TCt6iPLQ3R5GbPbDOVwqGSxPdSls54cvIXXSnMKdIDT0c/oHuyfUeVcDPsB
nEveqxcbqnHZLwEzeT/nd/QH8kcrsz3jquHHEHZ7D5bKyn++h+KPE6h1dHbfXGn2
fE52atzcAXCCvkSCZlIc7dkQ/YZdkiOGF5DazeQoBckZakwUuEXK6itzrTuHJbo1
cSMIRqaDCJIrrCwP7wmlUp5ix0dVU8yIsHJMwaEH+ZO8AlWWYdTUdeQ7FGPW43Pn
lBjUS529qF8FaI61ULJmNEqCq/QzypfFGeRnTPfaSE/45fn55vGhVzc36Cx634d4
JzKgOGjBKcuVrqaJyB55h3v3M9TY3YF1d3XHk6tFxmGaO5T5SYf9IrZE7E8f6gth
9YaEe1TBWP9PqjeSvx8EQJ7j8HOldXYV/fDVx44DEoY+nwGSlHkrvTxlI4/bbds7
nc0HOaRtJmATnxFyOm9CTbuNHJrEpRP/FigXaFvKvp/9IOQkvjfJrlsRHyyeLQML
X9ToQxPLuxlIj+e3uXCX+gI4mwS3SsCT0pspG0NnWDMqD0oVMsZm/U2DnqcKVlpH
NYPBW03clxdH/fvQ+TXV6Bt8QawWsg4dR+zCdL0xEhpbowDzmZlO4spT2WlHKWoS
oj4zT1ZC77nrc42RB04NKjuq2/R/YTrYquTa6trUpsCZQdtd+WT/i63MmkVgck/V
/hamCOe3/H7BQiZxDhewdMVbO1fUTj6VtRiJfhefXCWI/ikxHviGX5Vt6wZZbKe9
OXRsfqVz42jlanypheuN9PhZs8iv8w0o4NQFGf9JLf11nE0iVYEfikBlG27E21pq
PkwhmMi5VRIIXbTW6OIy+34NMM/jxhawdQXmJ4bqk4+A+xg4wNn+LSY+7wWPSnKD
9pn0+/Km5In68StGnMaWVj++e8dPlatPfB9Kqd9DjEGkwbkZibN03Hy42E6PDtiJ
xQw4vhHZY7IInBfQIt/70PdP/OXxbRLSnHnxgC0dVzIlaBzSAud2/AjHqYCu33sK
Hb/c6u3Ut1wqIarSJLnVRYtFQwOECZ9s7+030kIKtIMGtJBS+Rn2+xGi4rs1mikL
0HQeI4tD2NdS49iv1J9tc8fj2L7fenA1LbcJDh+lud/0NMH4/WRCB/yKwsIkJ2Vd
mcWWjEqYHeGDXPWR3oeS2Uqg+M/7NfIq//JIybKIm8at9BbF2a3FS1kqw/eMqrAO
Vh+Pj/2Abt5ezVJjsQxHV4IpnXFLXe3wmJhWnwCTwHkELM2FgghF8awQJbqW1Y8b
pBtGhkq7JZA0uqWm2zGRMZfR7+8oKGmHtnGeCwj7YzQz3h/Icgs0pzm69dHYE6b1
xhsD5MxCzLzT6a2htMS5taEaj7XJy41vtCcmyEzDD1CK4DkMm38+FRZ3YeixKiAr
KxgJwju/qxOA6M2iD0T4SV/HJkn+geB9bvf4Rt+L/HPO7twFrDUR7DnpKjbFCZvi
xY7zOvrajcNxvjLR6ybOGk5voXjECl2svKG6rDQ0E/dV1sEMPrEJI+6ZlbJSF7V8
SK7vt3VMkAaXPQLOCDAGIyfp0ZSUNGfVNPJmHTwo3ApDWqE4zh5rzVlNOq7s87ud
QJNIII8qaO6Sbb8vhqjehowIQugsxCdykESNteS8cb9V2f1n4NDtvdGbGJ+nmDhE
J218f1pdk6+cN9KkzZJ6YN6u2w0XFLtbCH7L/lAfZ1AJtL60FOkP+v0eIDrav62F
U4lbauKyR30k91MywWI0syyisvqdaFtfSWmeneRItNmkKnmYexq9PtNhTU3TYYoR
QFUd61ob1JUNiZWFFzFua16Hv9LJhw15/Ua9fNHJZd+KbLPyqn0nWpdHmzEvJMda
f65J0RVnwerxCF2VRGb872wPrEnbW+ouWdDoY4peTZF8oYxK0h0nF93zP0h7wyUt
LMzMjNq9TNu/PQ12G0etdqMv1CD+9R66K64xZa9YWas5axNfhxaAwzfzrDjnnw03
Ic0EGrkYy9OvdiI6u6cFLLzpPxM5/sQzBrktr75KFewm7+WPM8vauQuvE3cqBXoE
5fsXAOyz+eMneGz8gr2tdQSOEE2bUo/9wnZIpFwTwoHMkkdtpb2D2bIjJASuO7Fq
GMbz9nF/ChgzRzucHp0nIc1alnPWNd50hGJ6RdoIgU8bm+zT+9kUASGEPh7v7HO0
1HGSxyZEYJLyPti1wOjcPDL8KT79faF0JnTy35X4atu7n5J0/UUqM3yJtfJQTJBc
kvHZbUNizNXKFM2yOliPsAFxmoO61dR8aoXg0QYmjKwjV34GreNEIQg6r6LBlQI4
cJJndXEi5rE6J4r/80/CskiYk9U3P9F/dAPLOQHlWw08AA8rS3QA6qaEQoEaXhvP
9YCLJ6AHyj9i1owVTVBL/zVcZ+LMAr7dt/7LJ9KLZxgL+Og6ILYlb1CDPWGPXsTQ
aSJf+EjI0XcoBWlSMYWIU0JsK9pqnXcfxy8//jYP1rGQ6t4zOkBXmETnYp0yo6VH
p7VIkNff63biuK9kL6R4jqAvvYtpzvdHO4qNRIUpKzhCyUFxUroJ4Ai4DsNiubVP
26exnaZqIRJLNh6sGgjOgBFDKCOHbnFr0W/1lKNHPxvySI+fJZ9FQ8SRh99Vq1cB
wNq7hMLD1LdD8Dhya0zail8qO88i8rf5o64NO/tkgJcahFBoqv0aR15wK8GqfFYX
T+LtYkvjDt3/LegtTWP0QXmmkeYmjs3OvNNPsgWJ2YQdce/2xGFn69GcGvCfCaq0
8qHGoPqal0d7x111p6fWwtTA/UO/VtlKofTaA4vDIUP0LILBWTrONMNEC7OhPSUP
hf38OEOOMP1nwMfs5X9o9ceEf6pJVMhISkeh4gYrM1+b4X9vZnpfdL6IilTeC4lg
eRYdrbEWu6AWqLvnWsk5W0WgOIwUWQhF7Nb0ecw8qdNhpWhJ9XXPfa04CdM1eKjT
9RtqtGzKuS/fkt0wF1Wr6+n8BrSfEsulKi2BPlVzS8Nee9SzJgXo+H01bhqjZgrq
K52g4UgLfLoGnsAoD47OkH1DpAw1bIL89aMNPtYWYxWGmmwCSU9g/FuLoZAvWSVE
T0W+cgWJXAnRnxigHUECS6VaUG19VEoFdgIUGvBjAH/Vm4ftMXfIJC+PzDREYXKw
q+x1/nY/mOOho47McQP/J3Ct2oFpfv8mVlQ7v9shbtYJBRAgmnYIUCiO6EOwxVMQ
xEoPNw34hfgpe9Bei+0NVgS6dM4r44S03WsvxCL+8l9lROj54gxfJZf1nK1cTxGr
ZbBcah/ju6lnrtRPj8d4zVwyopnmq5XEaRv5Eymd7sDjzUrVv2jdjlxI9EMM401l
0PjWcuEkyy386eaJirUQiAQdfz3R81B5MhtRx74w8mlGoZ+IGhMCAT2mJCLq2rLj
sqO/A5/GlIB6UkqMEbChngbJi/9OQOu4tZ7YINTIcz/tfVsG78LmfyPVVKxyUUid
/RQ/BchEHvRwdSpbUFSeD/YaO4SpGt68j7XtyPB1HzqMQPfgISzB8EJ6qgoJvEL3
Ewdgm875sokpQhMb6sSAFxuS/wQ8Mbbmp94v8NClUaYVT5TRIF12CQ6ZFPwOOZhK
+sZU8ot/FWboyuXhK7yBhWI5QEM4VBcI6377ZuwA9RtxoyMYuBah/uLxjWuhk5u3
hub15iATqkrAPvzr5Jq2ob1FGTovlWO216wiY45zbiZcMhExLo3F8NkqzD/2g07q
Wu/J3gnjvQBdHJPQiv7DTLmknWK1JlZnkF29pJpjPgL9Nwuz0s+CxmZCy3ogrI26
muE20O+jHIksgCPMDTiFhXusXAwPmM2YwKt2KFuaLZIeOSfYQ0EyMOFIQS9kTuH/
jytyYPmTmNz8k9SLB7nMmPpCl9H2q3qVxSguqDm+jRj2QmTUOZv71ubl9d4lbH33
DuJBo6vS9DuFaAN7MI5+KLSzrJYeQqbsXpgoJzRhWKQEO9gEJ8xg9MTcyJxwg0FD
gV2L0wlB6R2WzM0T6LtoHop5m6HPD5ikE7CnyLPKCwopJ22HhiaBeSJ+KkG/WrBi
HPamYYwXjYymbGXtIVPK/eSZ3UHOb3Gl16rWW47f7IIyOF7ybA854ZMx3IFk6Ut9
y+6mM/fQ+qx77x5qtngXRgFeajQtvk39HFtp5szI0rGB3n1sWCkhIWa1gvrOZMKQ
dDMC0awaX5VuayPheiwIuWNyl54gR1aijB+joDvwuIyFgzlVylp5H/Wcz05gdBNm
hBsFqQtVTzitZHh4daedEm/PuZN/BPm9/dvcyfHzEs4OEOrkhaaEcOEAUwRkpl8y
c+AiEswZkq4jgL8WHUjOV+IbKit9SVrpl8rqyTKRT9S6+y0a7ZlPj9q+fTaYLqIf
t29NkFybqhoKzb1lkSo+HhdMqFipAbd+uR8+Kh1q3Ejbe7hWU84jZ8REW7jieseG
NWXV3uGnE7wuFfhEXM27ZtFbR/f6Qv7Meqw8c+kOguJmNnDpboJh/Y9KC65XLahe
FNSwkuZJSZGQhsoOZmvKmX9/VV5Jt4ViDJRsans7wwAv2cTSz/Q9Y/iagOTGtIuH
6dsZJL++wwRKa3Uz1l53wqc4FsZkMmECGrKwJL10jgQD/O9lQr6T1GVqE/2w8eDh
NiHaMT13ILAhh9ljFojFOO3dRovztdLgiHJTaOpAtGej/K3F2KzFzafDtx73EhFn
kh5bjKO4e69718ieW9nfd1nPy43VPIeSwkjqcbAWZmaCJDnDUlStvY3UlzFxKcUz
DVbABix/SNwAHL4OPqtKMatQxhbtfV/S2CVqHqr21RSdGHj+1YYJdhCjp9QD5mp3
z7TcwqwA4bvug6vkpZ6BXQG7yfG6AeKL7rTmObDSqgLxWbsMp70M7RPXs/6z4gp9
r4uI/wkP8UvgT3sWyv2VRrg8EpuzGOteqAP5KV51jmqU4CHTRgdsbHPWmMdCPTTs
tiOr2PaoDpeCnw+Mx5tSmONrcCJGJsC/tNkqKeNEqotZtdSdVbFS5D74T3KHtMyk
w+YpA/4HM2UM89JzzDInFD4KPNnq3kS6/vacw/+kpjqqr9vcnQ7Q6iMWd+sdjbO1
Y+b59lUCTp1kBMHvU4k/jYb5V0rdkK7yogSOC8XkKs75/QZmPyztaq1G0xLPIsvn
12tbl6aJ3AlFKO0l6mRvVQvbCAcmt4OtgXh7p3Fuj+fbGTnrHzxgH779LfPVQEyx
/JfnevT/USo/5Lit6KGvMNVMfELWmbdeAX/LF4/ronPsSgXr79ifGDXy6Pj3k11j
KlrMgI8HqBS2kbMGZ5Cna44Jzgdh+rXZQHOAnVeXtd8J+xJw2qntzCWmx7kXDdiA
6Habq0M9V3RaPYjYSllco14GuaY7GzNKR/rVGPU997gLR1Qkknrp4n1DmM/C+cvv
ixyIFOs3EmUszNZCUVbkIr+Bn/uWwuUsQrb5da4goKVnOb/3NXDZIlAbpYVIzJkY
Ej6YjswE3vp2d5qmtdwC2rtAmcV1GG1Yd+2W1QWPrHRYvpH/zURxUbqdf+57ggep
nUzeKXls0rWZySN8neljJ3h0YmVOiqDCoBaOXOXDJgGyGLZIWFzLpXhz3g7PF9u1
8rM6qJKUrjO9n+KIS2wG4CnLrNUxYeTmtOZ1DieulwibSw2U+rDrrlPBNke8Qv4s
Ivd/T9ga6b6iDSfb7Ad45VBjfQ1c+zSYDVRifK0q+m5xczIuMk1Wdop/y9XyOfTG
oNkxzlizI8uT9WOgKMuobycNEv40zbby4tZDBIpR9ho+i8cKzW9zcfAHeQWVxBUV
Pz2tH+ysG+XOg3VezWVAYg7UjlQGht9suEXh19uMBZb2BA/+T9WvJJUEwh2Wnwph
U1uKx2CsPnU9Spqz0wBA5ZawQrFm/U8aeQJPls+v6lt65IpUidwfJP3XvFEwUmHJ
ZkeegHEnA+3rOWeha9cg+GASgteXNg5UiuHQd6nkdWQ/1RNP7uz/NyEYb2yuMh6t
1vgMjwUKMgt10IV6XlzE4dzslfTICNwJ5B1FWAa6q+ur1wCSZBLUj5dvZ/zhvEyU
FBBeLZoAUac7W6vVTLgto5tqkRZvJvwUUAOVkF97gJp9lSdq369HqONXDCkMlTen
HQ0X3R4742QczKhX2JnVonVM3QKmfzwLx2cEHnz3t4pElRL/GPfpvxl/QdFMNJeF
trIKC1bYeHN+rbCrbPTfncX/eeXjN6Fipu7orAH/NQbDf1BG3l5v7eL11DWH+ech
raMxu8vvyV8d3HmlmJLN683PtPa+JEvMQ4eQlG8rEjbAV/ZOoOS7I6puGYFWqOxP
4svaWQ+XjpbrGlaqgiv/5Q7XXrhLP2jq5nOWQuGw1cFx4R7gejqj5sraM0oQ2Gg8
2TeVUloAsBFakHLVMa/HtSmRQC7ac7WmfJCJD0RWjq3VSC2OCxN8fPjPnKQQglL4
p7sfOGHNWpi8yOv68VBVZzVxgRQ8J/ABjoliLJDg8zftMYnnUQi/lvAadqa7htU3
3NtDCK1HQE/1qzp1kRrKSkyaW6eiJ2nI58NsrDhUBl5tLhOU4kjHxkKd/lfR2fpa
xXY9DXiT5M5pxpWzjcJZSsmqnFEnw3Q31xb0BCHrAdMd0+I7lgl9OZfEm5Nh5m4D
lHYv1W5TRnvXQ7fGaQLDT7wguJW24SWr+TM99jkqLRW8JiSMT3hZD/Sp9k85l7Ww
KU4NGPb8m7PVbpohGXD1zDRG3yEx89Koaq+TACXkV6VIHyt6tKdh5SJRS9jRrTPz
7Y/eHwEqyVukHoBxTVip0NqIFwohd2xMurfl5NitZ0moOEZwJKJLrkGIbSLxTZuu
Y1tj+urfY1X7U2gc53MlW4jbjU+PLKBQEG9wOwWoOQUbD+HkmQlOHA2vsUxt52sR
v+AjxgOduN2YyG5jiRLo76Apy9pyT0A52Gq7p7G2ms6uN/jby8H2ZVt/MIBcuE66
touSKCvbGQowS2ZZaZLf0KChrbKG+DMc+ns2pl0tNdHQUuBId6HQaywbzVWVnlbg
KihsVIoydb49AEY7Q/DOFlcAxTxN0Q4SmYA4rqWOVzssopxrpgV63Zzk6/AhBjrR
PzDc7noFauMyWF/mi8X8T/bEXJe6NUCOBUHP6CpRXerV9plmhcNXQo64YymUdlug
cRc+bpp1Efe89XRM8yGdwZfvqUSYiJw0j/9etdNt4npsA8Dk4h8K3kWi/LkZYvA2
V4056GIJiYu7ZauWCIOPFnWS0RgZc1ehc3KgkVqSH39t7Nmd4ckxa+xRqHp/LeXM
EMlQu/fFpUuGNbIpoZJheBVtTJvI9p5nFx6AzoxzTLqC8cd5M+p2J8YHB3on6XB9
rVfQoBbs/90w58xylqgUe3T+yZXp/gDWWxzkUjjWOEY6KdlbCopkZeUmCyg/sDy+
+niToZbb4+2chKCZ5RIr+ZMWIHS3JE+5B4qH4P6s6P8hcIp34mlvOykpUZ7oCCpa
CS/kwgmTo8wYK9tKo6htAiIFVirvbB4iEuOuq6VrVsKlTFGdkAcd+/lJcUoT18hS
2uYxWiuZUKVBPZWy3hRPzAjJPaUAIf/xDFxfEFfQBLavmpJhwXhSGDxPBZeiU6/K
8lQtKZIhobRoEZutppATHgqmFQDW1Ezps5moI6hjl4XQB4esICx2cJVjnCNClNzc
YWXeAoTDUGkXjTK20QrFymwOkmUzO7sYIjv8nj4CcAmRvTKIOxGCww/fiA5at7m8
mYsbWFQguKkJgbi8eAYf8J9bfzcH2jWN9JSwJmDF9Hv87HAAlrFZVrzttd7pFboc
7pMrtxSvKWGFWXf2/rkx/5BslKXmPB2FQFTcFGuZju0hW5wg+bOKXbNeeefvKWmN
NrK2VTdfEX9mAva9RgE7DJl3+wUksVm0yVdk8G1OOrVNjUzMICEukEgOIz9Ogcr+
AjabFOzViIzdJtgBOPkc/rf89YN+AyLcXhWPhhJUfRS6I8/gpXwazqRRbXwkvyMq
qGQZ+hyBP7Cf/coy7+rZ8s5oZLkA8ryvoCiT/kuuf170JUTB3cCIxlHNU6t495xj
TEwsFlzR2ZGbiUZqiwj6Sc+Ex/szhOAvTAHS9LNAy8WeSjE4OJFbjsZv2hpmAxgD
Mwx55VHDU4rF31yyFxAVF645UmSY0Fsq7VvbgM7HUTymKhmi9NIV3aRh2bps715O
zV1wnwPBcvcG29irlYXs/2RuTP6Ldfy3aVJqdLVUzx3RCevftTehUui/vI5OlVod
5HDe+0zHPw7a5a6114gaV3z50mRez+DNSLINgnLFbQihNNIszoqQQo4/KPAAc5NE
eaKdCLV3SunLFY+m6ahn66OyyR3RRHp6nqgRWaeXn1+YBr1fNBojXc3SQszTwwI3
CJV8G8nZySg/jZt0aphvw/T9noox25LpcgaVtz7fJMlLKuSxIk/ASHBoraNTRAKi
1X24rC24pSeyE+FzYdXHVACohc+W4YRSdod7uJisKgGMbF/wr6/Lg1bQfLcWwu29
0dYbqeEccKX24gMavu/ITmmCbDdnQxhz3MYIeu5ujgVl20+8Jjp5Z6k1DCvXGmTC
dAWbAaXgo+MEJp/B3YV36u0kDQu0CqEThqlutCg5kWZQoi9LaNm7+4YTOKXUntW9
HO375dYHs+B4+tytFq8Z702BkktqroP4j2ElzO+/6LW0Ek84eCIy3zZDjnfgCFBm
cF+piaz8ra8sWfU7MfYLRNH0cpPqsP7uexrIFgbRQKKsH6E4VCrrkTbgfUt30dqP
FSGpHBK8QkbBt2duXqSTsv8/GOI5blw4xeppsrfpuZuzH+S89OzqOQ4pXUnUBa3Z
7vTwe8ZnBDrtqhb4MDb3Gp+N9MbNhKtsCM/gGLmHXlQSsFUCfdcO28j7Kw2Fnstq
03CxgIzOzFO/7qnHKuz7Ox6a4pcDpysYr6V0v89YtZoka5nHrAe+EOxI+UEk0nzB
n4954OtywAOn0Ys9WUdUa3jqRx7k8ydWMs56q2nfCDrdzefGRypn0ZW0XoprQrl9
ZfbI7Ly8IV1OGOIF2xlYtt/LmpopqYUAtr6uI30utoCFTtFM31hf/vfi5spZTxZy
vMu24WZskRxXChL0Ul476Z/HSscbr/HhctFbtigdDbp1tygreEzt9Uaa0A6JF+cb
2uaq3iFrk6WAH9QP8MoP6pXqtEZfY+ZNCiXbVELTJB1Kfv8/k/4PF2biP5toZY4a
QlCwaT/Jb+XiBmavhWBOdqNmHOmKy+ri8VRyaaXLHrvHwx5Xc8Xru5NxA0rNPbiD
3MHQqCJuxOnjOuur/ISEpT5DQJdsUdHeGy5ZHfOHLcKdxL1X/zCFuL0Qp2I7UQee
U/p5SaHVcoxLD3E9s7xeFfNmfYPWOTusi0WwIt+GHqM7rs2PY5xYQlimNdxbPfQz
jdjnOoUo18los5D4hfGHVEoXYHD8EcVtlRMjmUTs8nyYLwBJi0qL6PmbK8fMD8BE
Hc9Df4u2UzrNim0wivlTIv/TJB+IBOMeYyGo7exzRd/BtpGY57N7fp6NWAAtEIag
KnrZcCQWs8PRSARxuopO8I0n4KUt3y/qAhiXIQ58lKTOZwnm6SdGueRBAH7e5iTJ
FafSaRGczZ4a6N6RehKwHtNcUy27TVzLOqYVOsQbDQ4YIUyJKckeTBVnGRi0z6HX
kG/d/vUogc9ESRh1kdIZYATKdxxMy95shIhCVHP7FCMzKOKpg4x3klovmMHGOXhZ
aoV3LMJ7swoPW4yGKZD2Ym9Q+yAOJ9ZKlXeGcFtKsRcE5S305yvy4x4A2PZ4sEL7
hTDXmqghjbgao/6c1mJKSfj+onBpa+ZP8j4+okTD4fRQVjI7PJ6Wql2870NT5E3/
ZgvX1VftS2Dfdy2kPUb4JT6rQLPiPoEYFriG5ALcw1ZlooI7nchBB8IiH1q9ILdM
zK0NuDKK0r+7PHVCfpl23ts85WZYsnhZUboN1QOWxM7Tcl378bsy9mMEZtvuz93T
ttdiMljOTsPfpbHCIJ5hIBvXWBAY8nc1wq1jgyuGc+Vsgt56IZ6jZebARR3qktux
TqYQrZ5yQenzN0mwIBDCiQ4VWfxXdfo670loYOv1FbqzKRORD92ZO9XC2ygmlF0e
6OR9IluEMpwVXPHWrrqNVKficVk4fHS1lAxz9V2v5JE2+E0cwkrX1zO7oG1z0iUp
7xlTjt6QbWcxLdI7gRCtAky4ZHGWz0gDVkr6azNo79zXWGhkNGvyc4kvy2ikA32i
fS/nE164yaSTRtq81Pef+MtIfmJbyeuZnKnm1zKuyqRnD3Sdg9b8wJnX9pOO/w1n
6ptRcxY6qA+5m+RcXZd4TXHGYfDzbFsnyWrA8q95dCJwz5PW3s7a2KwHCDyDjZYv
DZUwpM68JSGZ91GXMYtG7lt/2jeNmAsnTYPzfI3zv96Yg5sZhUb8XzGgvljPCUlj
IMSlPjrN1RaLBXSo/6NNENMCp/2arcBYCNJeyEAM/bj06JTUTg5VGYpQzy0uIRCY
HV6Oom0IS4smZfcmbNkXb+X8NhvYMGlsdGovkotVgUROrn9Y1St01y08bFfzWhOX
WL3FnL40HiscQ1cTWioZoenYJCf+6cTGD2eiTUhW+rwJg3NAE3cqX5Q1VAt6Iqhs
acYjH2/74JJnA5CZ4h59+RMHvxetA++RhSU/1mQi/Pmcj6EjrpN4gag+zSu0+ITF
C1UikegV+5eVa0UdeuU5xdjUNkf7fD0ZuJf3J0zdBtiCnEw47JZXuMvOjcELQ1Hu
RyOtEXpgcMWSx1VcMvi9ebh6IQuJhyFNQHDpWABgP3Rz4MwJ1zPcDf96Hve+Tti7
hrfzRvSFF/KNzq17SkuZX8c3r9r5CqoLfoQx1NuoATwihYDhrzrsyG8OpXsZiPki
YaToV01aJvNrtuDiqrzwI+Ddz6bUNcJrXB8YGhQIOahqEppG+/RqiK0fGkqSZnKG
+6po+NaaqdhRmklvLo059GV8Dmz9IOO96bBUgFCCzcAZY0htve34kRwtMJvuHt0v
l/xSEQLubs2X4F+FMimmncdQcoAb+Fm8OSv2J/an7gIfMITcHGDJLtW/1BscsF61
JKbzY7bAG5qWYqkCu9OsYjj0bwl47Pt1mlibOUOJanDv6AAAA1cQ33QiQWypS+0P
ISSDgTxTXPza79Fhl2Y/Nxnl1sHUP6O62trtkbma4NxOdPbUecuw5GF0DLcyf8DL
rvhY8eDqlvetqO4rYgx/PbQh6AMbgwwnIdnVTI6b1zLrYpomFEbgu7C7PUgTZ9l/
RqBRe1mNAxl5PgI+iVH9fXPAbGJHE/Othvn+CzIXSfrpLKOWLfJ1pH372BjWVBRz
o0hFDUWasQDpZZzN+Fdcqq4cfwbogc1pFYu+ao54ob94zf2EsizznlbdEh+i/Fmr
FN6mjJBRaDH+Fq+rLqQQe9eRoiiSYx3EJnICX7qmh691nX6wgTO8C5En+U3jim3j
1AXqhaBi6DCx9/8p0wh1lMg0Pl7LMu6knOG2WKY6hAXE0d/9lyc2VjQ5rXuXLVJB
Mm107I/cBVSoFX4GkPkbFVLCyyzc1Ti6ndX+CXufTwCPiXhAAuSxstRP0mHEErdX
vDSAM1U9pDitrasIdHhRz/Y5Ji538YuPt4ORLbsP5RI5R2D70d7QahUT+3JBP9eZ
AWi7rgF7tWutcTGLfIJAQt4uxYwHAmN89/jd1RaB2plSNDKl8b61oVw0Rmkhxpuo
v1x9yzBJUtbeHwlFB/W/rcUe8lOU8AfAHxr+wG0XFi8+ccku9v1OW1Z3HG9eGNin
XVhpuhYzCCUPwplVkpcM7OpruMcRIztnTEOLRp95s/lgt7fza8L7L1zxGbVGe4G1
d1FOrE8dHlKooM9JKBGIdrErZZCN3Iz4K7o8+xhl5qzNFMejGTjpix659TqNOlOx
8HvCGMVfCSgNqp1lHvaHtRUoWGQHL0Dfs+PyLBAYvpg42F6D8GXcKHFsND2d7atn
k85/nP7uCgRV+BYIRtAVzdtW8wv8WfsfkTp+TEEYCCwoPvFVDPTSf+9bZeC8oYcO
56r0OfMSbFSYxFkIIno4yxDCFrYFfkl7OLB+IopBwE1S6Bw6UqvXgvQvnh4Tt4IN
GMW91lCpY5awRNOPstOez6I4RcV2NWXes8JS/x4xvRQ081iwsmm59rG2GbZH2gy+
bxuZ95zlZ3EmVyIhiTq+PkQCONhl2ETMoJ3V5r5Nr9WK7HcjS07gFJRHCL63MD23
O9sXKRJmzAOEg3+PPvrtqAUv9uh7uioFNEu/zYKOg+vmDuFIUGxfkDK/en6Bgv4T
t93fpuP7gpz5cEO6fc/qAFEpcMOoo/I1JZ0CGo/5eD++3FUvB41mnkIcuCe2wBh0
Pf7jerBTGzFsMADtu/Q6e1nZAU/qON5MnxjxPztptkFonJlfTrUZO064xhKQwRH0
kiug/hZ8uShon34r5WUi3a/zzcvyrsCRzBudWUgFpadXif730ink6CMV2T+z7A3i
99Bq4mBo2PWBrVLEz/E/Ef+kvJf936d0lfhqNFsnJ1J2OblPGvfgFZm8TkxkB24D
59v7ASlAVo+0h/YBTXKCSEQ3BWu1vwGO5lRMVpm5ysz7X5IlvNybpJ8W09k7L37g
WrwhLKsbPXX1E8/gCuZs3HGylAOy/RN8oN5am3Q2z+t4aiGX9f4bJjDbY2M6BMOL
GksrWyqJ18rLV/PDj1+C04QQHkgA5CGLzNnUBEYNBQK8gPnB/yB7jVcVZ20oS+HM
q1Wphq74+/aeRdhqu8QwYhFrG0B40WsJBEtCCxvIwSEzbxJRgLXJiE1/zSrWtMK3
7/vvxIvfz883DlOe2YZPT0hbO9/ZjIbue+bXHhoc2gLjLv21LtdGWEWExyDm6sqk
70ltALhxwTPIaeevxhmzq/LYUuyKcTHxQqtIZVzSuD0wxl2+pjeTpGt+mrkBP2U9
W2Y0UVuiGcf0nGI4ra64cBWmzmgucQ6IRdAiMv6SiXkglk9ekEygyxCotjMj+BCB
ZHZMnfcbrjA4J7S0SsAXelv1guJshTMPYe0LsKTYofni1maubEllP91BtYzE1ka3
s9p685wQFWqIFrGCO32CYTOCT/TtRAA1tSwAoEqTLMaVHxyjplVyrC0fcyJq+33i
AzLQLkzWB50+ZjhufVCFWbQFcGuH1490u1023muu2ftflu36FAO1BZu+tx0BM3dP
ddUAE5xKMFAegJViJI6UvFgnVJn+Pcr1OyuwQ2IEj1lfOYTBG9TaTsLoG2b9j9sK
lQ/1RYoMw0+9romJvPUEgsaBt2VXMGDqSiRvjfHDg9YMhHQ1NbNrM0z3TJnHuuLl
v7RI5KPH2p37d86sEVW3NhxToDo3yFZqfKBa3sGB5Aa3QB3BM+eto+rZPEPqMf3e
jUuOQeFIoWQ9mYpGfcoIU77alXpiXyKoouVzHKAxxgIV02qImheWZoK9N66EUJ9y
OtKrrONu7MTR5CT5VCCaEQibmd3v6Ymsn5fmg135qqBpRwHAZ/MUypWmFwrSvsmo
MGJEMP9zYNT+neLFwVVaeTkxpPq7MtBxB7uVt7zYb63VNWsI+1MylbaC042cxUy5
tyjDYdbJkcj6iAj6eXjw4dzlZqXFLU2BPgKziT7WCzmfRpa9fsSH+OsVo9I+QY8x
fZH3ku8/8ElRay7nOk7PpvHRie70W2kB6aPmPF7+s3ypurrsboWlXq/JFJKO5xBo
QfMx2uya2/b4kuu3+R71fSeMyesZUuXAEqemJBtxLnmqv0GPsSsyhic78qKcIOM0
QjBGsZLo5tA4aEOaSEHb30TGepsrsIi5KCPBiZ0o6WROtee2u3iUT/uYpYFZZ4TB
rNJvm4j8qR9prD8ZTN5I6SZxLdQChI/Rb3KEGK9Ck70jSIWfOyNltt/cPDci2+gA
6oVhCm4PT3PlSAvl91trJoiBzLPVX0YReYZJ06k8LLgub/bJw5WDs7H/g7pGuvTz
CroR+dLfCEzTLEqqHByncAkTwKeEWAxtMf/qCZ0eINdtc8S8NNEYCUGGaDzZP58X
sWOkGTAkdrwg+B1ehhd7AeJgEihsmfg9A2PWmdo4cuNY5Jx+CKLZlC/NDmygDxKl
3Geq9eZd1DFsdOWDCTYKWrYZHJLQcA+4UiW2TZjXuRl6D3MdcU1l7qph6WJeOVRj
m2qzXP7ZRZ32FcvLKCuOL2Y5AqAUtPzJM4vGY/SoK73U/do+bVVlJTBp6iCG6RWI
QH70QpsfVArJvSZ9/12S4JJaZQ2EVmS9RZzk8XBnPBZjS86KObd9RqlYy0Ag9XdH
Th9aYRk67NwTs9BGJF2Gg7STrigCR/cyCwsoiXyV3GD2NQNLUIcEYyna1FUCuLtY
rFqbJxSdhwSorZ2KisPBLdwFyoRAzgMA8HIbvrUgvlglmhDQORZORldmjN2Pg6wK
+NuGvO3fSuVphLOmYwrbUv8SVT5xQIdKyjpIhGA4pGFhEBGwkUC5WqTjaKTjAnUN
LSN1fgFkZDOZitN1GB8DF82c1LXjgIbXhm7unjJxYBtYgcZgMIvhmymi0zWe6Hk2
aHtuRNtz2NpHuM03uHRZqxKzwOELaLZ/rnjA4SwR/JPcYMQxCEHjFSGMnGbu+3zm
0ZJcb7jOIZ58baMvuey6M/o5iIYhm30WcJLMYX+wB8YeFLG6e+uPTEPfO38gZKTj
75mRo/FdCHFGNxt330ULafDUu8DcsfI4cEMr5A6KOXF0s0TeCpmVYtEn++l+kTj+
MNQjavlQDcMYK9wJ6uqkk4QYqf+HWhj9mmhVixZ29lJ6UvY0Z19Br/wIsdV3YwhU
BMao02mERfAPDq87rs47SO2CVPpSyTVfnbSR547dzvMU/5oWlzFffXdd1HeEPmYm
/QBuei/yGK/jxbMY7atuTxtiM039ztKKIEfXWNxbwn5As+LV1ai1+EczsMwz26W2
1M2zTH/Olt4fWgJZqNUUfDOwQEvJu1tA0IpDdiHBjfSLEy4stUXm8so7UQ+xDzQo
Rq45lmg+5/0PfpBsuNUoAPEoZqmrQaV1B3k4ENWsuQvgocuzYuYqrgu5NnP0uehi
FNxzFMNvTGW5ew8plxBa/4W0WopoF9Jrw8LyEEOFqPDLfQpNCAQsl1OtI4UNw7Hb
OYo5cbZFrkVPnf/GJLQ+eAvFJgySgHeKOX8W9t8GIWmmYuxSuLpuBjIc78F78fPu
vSb2vnL72ohEkocNk0EWGAHaQXMf4u68S2RFoYpAdWCN4B35eWbOeBdv/sRGfVGu
aU9bKBkoId3pnX3WvUQBcRBchr1wVe00T8aDSf2izSIhvItTMn7Y9FwHNAt9B+EI
DxLRGabRbcGs87me/DKPgkVqf0WfOVC1U/a7dYxJ+JZkT+ijgiFdDi6WGcCgeNQB
DNCb8kt++S9mnKevON8MY6vPjVfUIL696u+xiT8Swg5HtSNEt+QoVTGMl6HrO9Av
hcf6we7Jo/aHvseabbUMIfJwpBoP74sApzSZjnHCGUW9fIcqGhtrd9PipJjDwNQU
GK9dZVxqPYRDsVFkakWCXZvJqXedqvA3nlCc+BR7sHDoxx1HiSTtTp9W/zwP6Zzc
DpgvDtUV+G6ozQ3y+v3d5KTx4152tkPrqt9MJu4hMu8XXlrTbHYwToO0EWQ/UOns
oyBY7DjXXviA7kPXWrI9DyY/OF1QwELNhfTbMj1ApT+sKr24GxXCCd5S9gHA6RTv
SWaB+UPZ5AQQaZiMInkWRf200i++jQmfyMaT/TyhnWOLdjUA+9Fe/tsT4wjMWWWj
iKnpVS3Jp89kZ1wdct2umXoEo93ppiwerLOq6+ry6+3dOt6rkgglXFnuuT1EVk8j
u1rizTxTVxsG3VDlnM7CIjEIem0awad6f6SNvIaFhbkSarx1Aauxf7q5oVuAOfic
bfzUEqxxjugz9ejiDTCw1+cRlsDFiuJ0aquqQ72KJSLbmTs2pnO01lbY4ircZ4DR
OyB44l1D6byYUxlP5lUmiJ0Z3raAwMXJX4gSwaBetGx6SFtIiNkBp29YM0gNf56o
SizK5hZgC91SXWNKJyVpWOK+4gf1pwAwtOuwPQgHN4e0iqEEmU8Iay7uT3bnuBoP
SqGqKp5FL/OLs4vxfgTqqVN3Z0B3sEOxZWtX4FSRO1cRmad8/cH4+SxppW5mpvDl
YOnkN20GaWa0cwjZu1RLxwctyaut7o3ntc7iqDj1fjboCSzLABANOB4FBc83qjlT
xVVSsKNczMtL8XAKTkI5h3Lc6rbU13F9kQHB/gkGA3VEIjOPfET1tYWyMbUvfWF2
6yrdtt9J8BAGbYh9J78qmIuXV9vOY3R6SsfrWVYSheOyR7difeNe8KCby6pA/qju
CoBkS5h3rSLlO2kepEIRYbPhEMMRSFZ2EqE16CdEhCnGV/g217V5fGyHuXNtDN2+
ReeU3EAfa4LJ0QK+kH3pA5sqlVgbQxhoDk6cVB+AZ47RgStYEqf5QM/uqysisxo2
6kXCDUuhUZySHisdrhCQ2Oi+lg8cXZzAQUXXqujTW9V2tzekTMcEJjqFoqfd2cf2
DIbI+AfNoztoVH5lWnJ9YyKwK8MhC8Z9hxTNuUhi8McAjLrk2L1NwsYFRHtGsedK
gi4oy4r2G6/O8BkllzA3nzPX/EFyaGvAxRzsjv0Lw7w77BefqiWvUfyRO/3sD5cC
xMcTDHgvo49XlHBnnNwUKszO6DcGQO6TY5oPQGrOXL0/gL4KDmmG/04rjIzonLKK
ERaLFdDELPlHXNrJsx1jvcKGXGMFjLyqNYczohyvbTtWVyO5FpbsKPqkxEFqpeD2
AJFlGuLWSenEW690kT1DTla2o2Qww8D55LVb6t7rmXbZIIVXXm5eSKUcXC3Vjf5h
0k7gw9dh5pEY5kONw7B5t5HvCn5gD2rMbQpAAv+fJ7KbwuVEsDrUNlAFysGH8Ytm
IM6YQg9Vg45xiuTIeg9aHBz0yxuicndyWm5joGqjihUJapT3nN4tBFDnRx3Ppy/a
Vs4p5g4mo3QYJKYu4UdNxToJeJkhzIWUhFZDGBmkTmIcyQRNrf22W0OCP7wbII4h
0luWM/oxDF2TmbqQ/zIfdR8AEY1IpduhPBKeq/oga4tULPn089NZB/JNTW6SdA8F
zSSrT368AY5BA+dubgfoE7nnVZZTKrP2aUnojRQFwryT306vcE4DsSKQ6NvCshF/
TEW2ZmjpXip2PwCR4wQKe4Q85gOaCwCxnAhkxTgI78FoRrXjGKzGeWw1sIjY7lSn
Sc6OEa28AXbgzpDIJmxUegTDey5Jdi11P7T5MFwvo7MEpDcs9Xxb6yDQw8armcIN
guSm8c4O0L7Qq9S3NDLZzhBrH+epXteP32r41qMO2rukDl3XQ+GTvb/9jUdz43hM
V+LSkTsJBC9fM0/saQUHqicxgPWuU0ybYHw4qimAf2PlenS6CHUrQHX3mBmYTwt1
u+mXHQmXd88um1WQvcYr2aF0gU5MByPCv0gIXXfR+kCN3wyiWwkI40CmRtt/TEmp
2jG7rBomp3RwUz+ktVKbgb+V01/w2ZTxIX4SEWNwHJQ6viYfNYdrqKEIDeRrWqWu
9Cyr8uN6hdcV4T6B3SvE1IbxUR6+WsUBfjCcbBMymyCOBhZmwv7uJrXuGwUMP/pp
0ycOlBO8raySSPu4JwcQS/+JfpOQzdC4eK/FcMCe8JGMKmDYg3ZBdlTCJB2jvNos
jk9Py0w8RHEPd67SOu1y9CtKdw+NRrtRUd95jPwXqYm5prus/clcqlp7qpdWMK2s
ZGSOtZ+H0KwpeELs3poieHTonc2a1DtuoyGth4EMWgfOK7a7pnq9dYGUkAJ6WQep
iJ7TcQUwRj2wRF43vvz7tYsbvIodfx5TRJj1qBT7w7pTkgKTMGJgb9fb96eKEm2M
H6UkPheAhZ2CYsEOdEmKIUzrMDVJOV7G6pnqkls29nVNErvzdjQs3DDdSHvJnm51
JoG4esw3Z/2VUC6NPwYzytKs13CW3Q7fnUhiIwStMgn7NmH5oZet1bbtJJbaYNf2
GF/0nPl/Y0ak/dQ5a2vrk6+Ic23n4utL0pE28rIPRpT6FM8zbUi6h8ISmvE3bWAh
PSdgi+gYjLNA7xhIyjlAsS3LN1ZkVus0lQff4jILkFqclQfJeLEGQhn2dCCqb9PS
5/DO6KWUa7mxDSe/h/1GyChp0InuMBsU8gU52Btx8EzPtFskgaHhdNszqmDkqD81
U483nl/HfjIPS2JkHa4NYgdk0MTqhS2+inYqIZhzyigq83rA2xZK/W/pGb6ziZ3b
z3B9JlHxjMjPRWrcDRQFYSqndnpAUrZsrPTClMm39Z1+cBNGJvwSxmnIQcWgsz4F
pY5nR/rqMNVgNQsLJW77L8/Hj9jXyhPRnqokgq5b+DlwYK3YLVxh+gU0gsgFr2K8
nTb5IWF+B4HTVoLg2qoWeXNzshKkTJ9IpOIu4mCcCOwx/Naqzi5Ea2QxabkihGAJ
jR7yxXAlwZ1PGbwuaMbiN+J+hHridNk0LedislMa28m2E5O/+ED1XqmntT+obEjk
nq0Ia0PyaXd2Tmv3hSf5eBO3wKxJ6l1hdcDajZuch/eqYCByPllNiudM9/SrJHpq
xPeTmkEUv+Ge4wJZb9tEAM2T5p0vyaaQjZO45kHaf7Gti/eMzQDEbV1mPg2WGAeH
d8dh/j3NMYBo48B7iywuVRLZJ/DuGFkBEh9dp0DbS3eyO16VP6eQ9ul6qgnfr2v8
F4wdLmeAfs7wnPwHtJ6sqx7/i0Xth92Xkwa2eIpUWT5LJk0Zej+5Wt8icRE0DPc7
qniY+r/dO7rxF1V1Fva7KZnbOJFbsH4Xzc5u0kWU6EwmsyFmo21sJUsK5kKn6T5I
NzBRanaW+kj+AYFNQKhcTMr9WrVj4YuW2s6PJCH7pramxa8SwzEXtxGF7G966bZ8
Mtx1KFoSdMR947U0xO5UQfKgEC6QPnSf8rS5P4NjndeHdxXf+75/cyqTaz7xzi7L
cYySJSKH7dxcDlC0IAYdZY7BsFkfFOMs8h6e1Xp3FxWWwWdrDQBBNthnrbbW3rWR
dwiS2vDG/92eKwPecgQKNR7ruxuoXt/dmzXa6ucwWpP3iApBAlh7QA0Xab4dXoVv
4Bk3RsSBuZS37znmrbNxw7Y614PRfSURlnOOA1JSB/Zq5eM7ZfvSZJK4v9BZQ6n6
ZtFUtgChZ0v4yXVsT5vdoJEsmOpJf0j7qu3z4npjUuBrxI/BtOCCCWnWPQoyJ0yp
nW9MkHL4BsMucCq2b85wDl3k3gloY/AoBWOn7gm6XAz4X2Fx3NOcvHGImeHbgSjM
GfLOxguVjCVJLuVR3U3eADKsb3uungJde5YyjBg/W284DTEDcMrTA4VvVYvG3F3p
ElS57ibxdH5BR73FEkr7C5Hpm+5BsyvrRi1c+ts3g97h1GJvawEWzhrYWVPQOxYS
PCBai4A/X+/BGAFIc3mmw3Hb1TUJXwT/JOj4iF5Lj/wrXpg78fKptvsp8PyKwAYL
9mRA/JQ8dulleIIZ7hz0A3Wwg9e/+BORDAyACGhpg7kBUpghR3L6h3DYKo6SSYnQ
98Xo6Ik+g3sAmFwo3mbyWMCO+G62IqHnwvE1FidmBNZiusorbQ1oCOZof8ioHqvy
t+oFi2eoLrR8pNw5qZ2scF/XgtLalXj3tyswVkXYKPuPp+8O19krfWVKKaND2rYo
yLEi9u170RDfo2OCGkIZ87bKdwKRPiVhWWmuJDaFuRqPgChr5zYflViDikEsIDw1
3LyYTLadC2FXkutU1AGo5sojo5lIlfxt39ESdfJTfYbgQ9zpvASEeK8a5kse1KP+
KKt2ASAhCf0Ev09KqF/RVnP0GuU1OumHRuOLoEvnNySrl7m9eqFRwYGw758OmxJD
2bCEXlv9mDyE3T0k9wBx12Wa3a1RGyXjisoYcRDfQmk20OSgSsE3Qtzxi17oniED
89dcJtibAuOEgg1oLlna5eK7myAx2WloMjaeX3v89v+6HRNedPDkHIrAP7KWugtP
9nT+xvBTPHEiOEaQ99wWFp86HtmGY5Gr9VCvswG5qNgXtRErrjW6CPP2iSmzp+Xh
asRM5+Mpz6NSryl54vvJwgezdaMmBU+ZYKQffZLx0zWJq1GEACJtQqm8OCntfGgQ
+st9M7GhikbNd/NTX1rXUUFU4RLO6zckEMH/GvnoomXNk2Rk9i107VwklUQqvBy5
sZI92SHd8Pkr2Elvtk96NWGHzS255gP9UZAMknvHIBD6cUdSNvxhis4H5MmpDbwA
rGd311Go8r+LZ8wLaON0AIijc0b7WL1h5DRBK5j7484+dLCt+mSe3gcKYYmJ8e6V
d9peOKmEU5lwwVV0k/zpq1SCvZGkXEVSvtULYUqEu2EOn/kark/Nxncc7sv/CGMW
ZSvdmKnzrByKbb4HVIKiEnBPDZ0roCm1z200p8wubi0xkEVyckZU8p/3HshXhGxT
Iaf8hOj3+b/+WJ5y6cFUw9mLzeiWpW91JujH9r7XK7cgY0Cv+KgeSdHhCFsbv5NP
Atur6XG7uaYVFfkG9cD1fcxi43oDM/tJGy7PVAwLAMh+IrGD0J+GQXnqTkn9pKSe
wunu9298A5aV0jMklubnSA2EqXk8wF4E28jKjLlm5JlEyy3iFPXrrLC8RSpYJ2N/
GvGc/ZXa3OqifjZj8tKtMAR6Gfm9DnSZ+NaDWWJK2lnAnSGRn7b9X5yBhF009co8
XcBB8fv9HkKDPMDmpQxZXAKpWgD/a1ndVMR01ucV2CxkEOJYSlT0XN+IAi8a10B7
qmdn7hz42OA9+L5yPSgUD0YWEsqaAK+u8tF5cMyYedCnEXZZZ1R5VViGfYmhW2Sn
R+59UliP7e48/Tzu/xCJLWkM/HdVygj2Gze7lveudxv9z48FrtSmtEzBrnN2dvmI
/A8RK8ok7Q76/HoBop/1pRD1M60zxp2HNGjpcoKc046pgjntoQN2lNStKsA9jauI
QWRP5Ganb6GNsdgCarheI0b2XTeoVqnb3tP1W6zSy77k586SyLgEdy53OjsGhfCH
gPryLMNhZ3Kdc0MSmxrhfHR27jvcaP0+PwOn2TZ9jUjx824a5tQnc0kx5KgBvXLO
olRUvvEl7aTBugMTELNCZ9kxc9IPJQENhovSKJnVP7jzh336p3K48Chb5QQCTLe+
yN+z+vTKa07kyGqBGMGnXrtnTHFinhPfREfJIed3U0PKAzJcaWGntHQiUjJ6FFvh
JtvLtzI/2kXqRyqYCaBIdTYBvU3T0ggp5Qp21+oz35n9kCPnDTHEq+qhLXwggCJ5
tJhl6JC190xZ+9UnmZUk0j3whcF85ZHPfAuZDKQiRXvplhQvHkKzULTxgyQ39xon
k4Qxjx9ViPrOqQ4NupTpF6o2cYC+wZ9WCdxkNH9hxYSDjb4Z3Jmmyrk2lEqdkPY3
5Rj6/ByZn2mD10Lbs5wPJ54iEAS0rmwahGqxKh6Qd4E2ayIKdomf3mlMLY2MCMYS
lTUOXF1sM00rhbgaxT7GgcscLlXQ0FlqlLignYdXweurvLwvUxTtQ/yqNXWlJFP0
LLX3KOhYu9PZ9M9iI+4Gf78OzZcPkzqrOVEQoHHobbg6vMKcAAxdrU9PiiK/lXFP
SiTYGNsF60pgC/vwggdlCwdstTMAf28WChjpiJ5gxk+NmrWXhv3TcatXX2kfo0B1
0gqLGFl48FNwn7LpkF80kOtnCtcrfwmklKLAWSM1MazDUcQmZFUobVElxX+ni6B7
zwu21US9nKFDhjqjT4/aa4VwVVHKF+AXxumP3A2JYvk7vVqwj2oiCbKIutVHFdWv
/y1VdiP4kkcpS3tieM+ekQvmqcYIgMogklgcvTQzcC5sjMb5VPFnBNFGoEmHs4OH
WmhyXBD+ReZI/TSza2ruuOU8OIvK1bcSL1S05m79l4E/68ps7YTBWaZtLSc7eMRC
V9PJRTum/01lENFv12x04u6Oz0VFm9muGkt0c7n/yjCzO1jTlzVVS5sOV4xAkG9Y
QKUVXbfrS3CYsl2GWD5QvjDDndBMEUo9idyafhQVEQ+9nLqade1PjiwcbOtzlTNw
AftfQlzunxrMsO/oJDBdtffFUbG5kQk9W1mnJoICAyDLnfsAL/XnSq+j144LeAEp
yV2lnGXyMrNtHvg+wv8t7M3hfN4VGVmjME7I4IqFBHHAu3kVVCbxo7cD6KfEuFCS
nhzY3nkECwazeIu6hIWHV+/Ty10EGK+KtpfwcOMYOrTP/GQAG/1Bl1hgYkQu/Jlh
NqwhB3h72KUiAhhFLATwKArcUzemAjJMrlI7Zeyf/E6uLZxPsDUX7eP9VDyP+iYx
B9lfzU1XyDMYNxikW2tkHC92lIC/gQSAb5LCAOFcrOWM1XbLEmEwabCdk87hm2tl
Gl9QNmiQJkfPNszLIClqNXLA7ZMx/LlZJguCk8yPVplExh/kNNP4zDHvQMkU+cek
rvJ8546hbT7zKd2NzmNIbjJK8SGUsCd2Nu3yf7JaQhqxL+yNG8Yu0ssH5bNDe06s
HSEVnQ2XlFfgYOAc07JUXRjv1CB7fRcmNJSHQHLLU0zv4e8VlyNk9gUaJSvPhaHd
0TobWM6C4Z98oh1YQYEZ9BPIFcms6lODDlVyoPxfUdNqUHa3K2vI7uhcQhbEO1NU
LEpOXuDnMt/pDXQB4mceJFzvIwaDJY/GljYKFbjgOn+JJR7mI3hMVkZNfbKAcrsc
JklHnxn3q9V7dQd8UuD2Ns/volfCOlpaMKA/j1zyY8x8mLnTufRymeVedS7EVrCF
CqqaWP5JAvvAzsrq+mwo2Ztw4sEuikU5CCz8fRncpuNV7684U4ySU4R87yRlTp9X
Ogu1mt8VXX4zzqvYQ1qmWYs7+aCVaoqSH7oWdI1t6B/1YmlBpvA9B5ONr0LqJnGe
T7rzwbJmoVJeleQ51cVD9u3nqALBDpcrW6fozivS8m67v0/IKyz3uy74h29kToCJ
CUrklPPubc6XSW9hN7U8FnOJODgC4XiVe0DEmFKqZRHnsZpt0yFrfU7pnmbQqJ0/
g9juZlqRKxp9Zgv5JL8r9taxiHlPYVrO6pVFnLEsHbX3tKikhoq7tr47Z2svMcv1
2TBnFufrveUgwDrqkTg2+twlIu6AzXnMhjiIDoUjAOtgIXAQK9NYdfslDiRX19cq
ni8/+3uAsC+3GRaSj7ij9OH/fd1GqpOPgcPf7bleA9R0o5nzKJgZJ3VmEr5QImt6
viNo1zRF4lxRGXD7dudaDltN+/cyQE/ktCsUoEki8nksSxkExvVt6nA26DISm+bW
Chc9BnA5p8n8EVCSquqaE35O+Cm7b2gh0v/ZNxDe1AgSEQHQVoE8YB3Ze6BJ6bf3
IDEQ1j1e5p12f5QcNRElo/fBwzFfhSDmIXaKjel+0+zFR1HEVFfBg4cbrItMrPh1
rSg8M8KlEZfNa9kg+1Td+fBxWLF4Ig6Qw9dg1Qlwke54An/MzkBCzxEoLaTArYEe
8LIrgzIs5ky0oLw9Ku53qsFbGu+mAMuGp9HS5AMJ1sDBX2bXYkK1dP2qhTgAOkmo
f4DXtOaQbvEtA4LWna1n0MXyBfwjPA0MhWmhxKgP7wAIMY1IbJ57gG9aQtDWdJJ5
Gfrtr0Y/rqAUpIh8J/Tuxn9IT61lUDGKNS0MHy6PCt8d1YKvbzhqhefgtHzpnw/M
E8vbQbUCJ5HtEGUFJJEU8btLl1MYWgoC2O1NlLa67JR1Xev85r+MYasVZB+n/2RQ
CDsK1OdAu05GZQpj1uBntyEJClU+YazD2vycgbKqvBlZBHIDripS+LuyB9W3GhTh
nK4yDqP+jyFwyLpvHuBFogcel6Yc8mpZ1TEIEAzcR7B1YeYlTxshxWcPlG4POKBY
JNoJT/5uCZYo5GeeaTFaUN8W0cWggxf3Fx/Cw4WBKIhw85cAfbFDBrf/PaUB5N3U
cQ9nv5qlBI7vMTjyOK5SsiNlGYsxhPuwmGI/PaG51On6SQEEE/UenfbGYK2V0e/T
bQAz6lwZu4AdBFPQykgpPu5h+/hM56odMCFDGdLRvfyuXAl8oifMdbPkrNm5+ZvZ
2LSSyMwf40Izskw7NPnkw2H15Vc+Gpe7yau4B7/esmTIOUbzPrYhixnwiTQBYw1M
zPR6OCvJBL9YPLXl/foiGTOPsV34KcNdDddRmq7y99e3jjg1Eo9taprqML8tIjKO
0dH99uDzIRQjRqMVOW+IvRDWGv3SqlHdttPA43MlAtWqyXqpIN1XELNJ0GFXixQ2
9SRIpwzRLhUGBJ7Ke2pMZE0KPbQA1C2Yno+HBWx7QpDV7Z4i9khe745LJoO/2Bpi
N7/CIsexcMXeoz+XTPxeR2KGtCwQA9vBHaokhNzD4yz6GDpIKh04SVHX5KlxQ6KE
r/NC86u7FXTRjzdEFGUi1M9bPE54whgDyqv3FT6rGkBbXM1ihiGa+uFBrdC1g1H7
ajYjvw5ah7T3gCPWC2R9UjwciagLYXHn4DCCr3ax1xhWbWpoJC4fzi4UTao/jzNi
52EUX3V+Z+PaeHKUWU+D3Qnsx3WLHnnzPFIICAlLpX7g8JuUJhn+l7TBH6KTBqnV
9Iu56uhpXT8J8MB/kRL9I0GY40GO2zq3EgpujTkB/uuTeSqDqc+k6NzwsmdLtU1A
WnWODZ/TEdUoWiRt4khmHqEGQQTea4dEOumY2cJVJmzr8sZok2mvXrQAIE2YaOeY
zk4w1fcjqR0hovo+7N54yVSeQGd7r2tsc4ASDnpZlUUZc+RDTogd7PyZQSGn1axy
0raSs39AflUtvkCVuy0C5Xi3Vrl4Gz9KvS3TBuksXe4v94bVLYKOVCtrY3OxctZx
EYzgNlW25Oo3jDQrPPT99Sbo1RfNx7AUu7jtrjStsGqFyndJh+Z0z5LQrrI2QGwV
5DsgLDFk1UT3Yb6QZi+CmVhT92OuotXCW5CYkqVTUugKdd0Gsuy/qvbQB0aIDHU/
2ubKs+nWC9rtmMDt4qtqhvFzSsfFqtbGydps/qwQ2KjHu8TjQRs1SSCBYVDSyqtG
dupOzEYllJeL8NDaB1hp0B9xg7H4AlrZBbCoFvV8f67V3rl7uhYuhQBk3fWM0R62
ntkRgJo+kEnYfOtboLLIlDK3m6Oo2WVj517nZvV3YOwcrjBPix99Okna8GTYdDTw
MQim9OMjfIPG0ALy9uWxNG5V1I23Wv1A2q5vDgFQgLw7pjhEN7ncuZZe+n/ITxaj
OAlXSKwbKfOSfA0lNReCF3V+X7ooTU3rrPrP9n34NRH8qpq1tQrYoi92t5AEc1Pu
nm9uOBDbRqWzP1SyBvhkS1iQDZso7oyV+etr3TIOwNE9UMQPOONlEqtYDP9xYj8J
OBhRgjlDDCjRtX0HfwavyAzyv3wK31FsshBoq0+9AK8Cc71bhRRsu8lVTsz8QGyJ
qdyWZf48BFUic7UMR4QLH190AALQywlaspuRA/MBnAMuimRcESXErAMWAh/FSf50
pOjsEDiCL/aaF7exPtMllEzOPSGiCbY5WKFvebVbNe0q/OvGkZWpl/cYOwC7N5vf
LBEocn171pyHPApkH72I2ieZYR8VyujZgywqdh+K8f5VuYfnUnaZ/k2L6RVbw7g+
E/PS6tnsKHgzPWGFrKDhLN8YHbxDB5eVCx8ZlYObrS2uqCERzDLhapaQsSgRCgCr
1Dffj/JZsz4g3qQR5XNxCWk4gD9n/DVupadDFs1W3jW6d28Gndm/ZVKATIzmf2iK
Thn8enEsBkYs1Rx1zWfGCozoKnF/wGTeytL6XjmGyzT3qEkK7+TE3UNXytXj16gO
1ZG9pjIHEteUIhpVlzFwlLFAwSH+LaPpmApi71rUkm9B9WxZDCWPYO/cWbHL8iFz
YAdZKQdq8RjCIwJwLgIJyirVinDc/QVXowk8b85EGo76wcpuVjpxFWI5vNdO678M
Z4p2ix3gk2ofPg+tS1Cnn8sHkaXDteSHYjTJZmU5pTSKPfOtGBR0HjP0GIMM1JKQ
ixoApQOuHrilDM2l8MWFqdQzgLL4oO7Rm7/bwV6YIWPNFbqpskQzbYpDKHjpAw5N
/r9DK4hVKNL6RljrhuUGT8qPOrotH+LfokvVqlCW0Y1wawMpuAxwDxpufqRSZ+nC
jWwHk4DQX7AX4M6KkSXy9cwBazHhKk0ig5D2mIVzqHTy/6cQiPEIU57doMaExE3C
77IQkJp/zeLhbslU+9kebj/4QAADhPEXdJaSVqzXCoSNz7u+aAp0hSzzLKucnqKL
W9LBKZwfT1My4btH8MQpkCg8Iqu9VLCV1URysyij40FuDZbRK4nuKbXbAa8INHTz
8zyk9B9LJXfiIUk84qzm0tzhYjy43zLSE/qyLBD4N4e4ZCr4Kmcd9azkf/rVql5X
8vhVHE+BJcRst2ELE41MFtUbviNMlvS9IYSnpuFUzmAWCe17o8qjkexw6RuhD/nq
1ReyIrkQfpVXo0wF7IuaoW7tW2qodWndxUC9870S3kujTzkSRCjKRRk7dv5GUF06
rwPQR2DES8UjUwkA/vqGqOT6soygXAWc0Y6D4uYy6FzUtWmfDmeh0Lp764L63ohB
ZwGJibN64Di5O4ocLU2pDnctww2ZYexa8F9i9R8Dg5XxDQ6oeqgenQAxeTNsiFgH
YrELdHP09lfoOTusEpDmMNF36RSPY1hqhRHy+Krslc7bS3BNU/91PBTt9xeEa6cO
KKp0MEocyanOdxLv+y8eMwMr8aEUTYfhdvsJcfIXO8d94xdLg5y3QW55J3TLJwW7
RpUbGIACNdubA5qTW7h6dbZ5/cKfiiLobEniVLClvRsbnO7zSPvAFg17hCKwjeez
k8nGEIfvroE3rEue7l6GyTjlzZc5bTNir7d78e2fQxAvzwHMoYxz86zJBZC+zyFt
9G0Sc2Ufo6fle0gWCTWOX5OobVnZqAj/sLKXA7whIwxqvcH8Jyu3x4iLh/FuLujE
AwzeablHOms6Uq1mOykq/iVPjMRL1BP36sehROlOOcOsbyDq+sWO5VJlB8TW60EG
ySIzmjeNKWua1VmV+IVB50ljemb/WQy3/Ch4xJMQfjfPfjUCInsECMfzDuqaUTS4
nMNjYmaAsaJdujGtYjcRc04TRc54yxqs7J035jg7dLQrS1ob95v5mHbnU3pRHyiX
3/759di01aLnYYQ3Bcx3StG7tai0IKAYq56FaAShJBIRCdUxqLKZ5+NJxtdXikW3
rSncOGjjCZwcUDm0JLviSWaiWEpm01YzM4s+FGCjBlX556iVlzdxNbhlRhiu6o27
8coXFLTH3gai7/9Ljq7U/RHQqo2mHWqvQWyh41SAzHUwFZZmsgAevNT+b0FAX/aG
dYDUqGHQ7KbRlhHTncWYD++PUdJiYanIYsvNC8b9y3j9l/nVsCCKOiER2vTzwZPP
UTya5vhwELPrvGIu8AkbQ3533QQP1d8VKwFP6Z28Afm5Ve06AT21L1DhEo1epgfa
wLDmy77QnBPjeZE0DGuursYLjtLnLM38oYhuMxUkY76TSReIEI8l5YF59wSktlCx
T7r5PBFdmga5uI9oFj+xypObXQz5oIF3o5/GAnSy1XL96WIk0plxpleLIJPe6/Yf
JA9ym0ZuqLkIAOxTA19IyLrPOGelL58odM13GTIDbS0c3dnJkKQB4XYnwwvwhoyJ
zcCSMQxjxHaXOUoCYmXUcxvLVbmZwKknTJ0lraBYxbv63V9jpbjUXF31QzAY/oNF
tzTRREKSp3gKn8zJirEQz5LHpP9bL7dagxErTXvY5475CpfHp1v+9uU0ulqXjakU
qy4XDoD1e74jItUppjB74R1O7aM3C7B6X3gKbdR0J+s0dJKUuwGcXpQ3SAOIl/cH
WYmcmrOeUTrujwm1DwFR/SyaVGMG1TnpxKU4whJyM4JZ2BHEwmNownW14dY1oTvq
zZLPrrblOpjLBW/vLMZiuVqZff688m7DK3hP6EouK5rGNO9OB735IX7bWmyXAMfv
0/zGxc4Mg/VBDiu26rNFmZ5ui4v17cfyrhME2ZJptRhRQqnWThmTiOmHJPjRrRVc
wT/n5jP3f/x+8xotG+47toyJmi/zvkeWp/VaH5FUvMoweAyTxXnIcQ4bVa28atnV
Hoi/ZE381IxPg4kjgoX7vBfmQmjk7ebzY1ldewtx86rBIZTGpEOWS4K4JiSDr3Lk
jQJ5PZQDljean5miuARvaTSHob+KEoFZUch9Yj2nh4WN6ct+EiJnznblXel4Niud
s06xh4EH++fYoSIUvBh8BI6pwtqQifg4Nm4S9t0vcL3+8JdABU0fyQHJJhXOAiT/
lRZYq7CsS6yfVs7FEJwmW4ZcIRiqRRCPO8cByhIFgrjskG7WllWNTVQKxoka3IUB
H/R6IuK6+Ix+RatECgfULNzC6t0iSTBsgmL3EHVsKnnd27DllmjY4ZORZPvnB8V8
3FuX8nlGoB5AmG9IkIOeJSTrt+uSBIrQLB4ulJkPhkGf/BmyegJ/aoNa/i9jxnCM
OY2y5O7Awx0m+bgp0vjRJZ40yN0WVCqgRDDM2QTy/YqsCnPonYtBjrJKSPb1t2bs
uki4kYAN/sSzEjODB82x7Z8lbdRZYY8qk+OXva7xbIyjRc6SrQX7/Iriy/XN3YLn
ygZbC710CrSaddVnplsvXOewNBojPNjAtWY3nILTxccHHDcrB3ieS6iZkQ6knJo6
YB+rGJekdvPRowVuDX2dok8Je8VTlfz+eHshHzg8XiTMElayCYsdWO98HUPzetjF
HztugmN3b3XdNqT5Ecx5cVYw6gwihwXXt1rDkoDBlGtYZcPOuYB2P0DHJkxF3j+Z
MjMRhNLnCceMdpyQwi/ReXCruAj3nOFQ/z88MJN5+m4HjJEF+X+JBHrsR196r4pk
VGCGZjoofEB2u//j2s9SZEzCrjOJgvYjZNi+nh2jc3PLMh+SwZg6XzCwoZo7zvju
EPALgV5MhK1MqSD7cr+uZ1doUh+l4gbMFwhSr7cBqCeHF88Qqau4YOY6nyWdpUqA
SLFXrFqsGtJz3C/7JAiFaeAPLa33KNCfdyqtFYs1C1LQ+fGdDU9/xlvNXnSJmt9G
F53So0oIquGoOp0u0DCSWTj9MvfpxRujSM2UQOb6UnWb1h7vbGJM9T6C+4Wpj3cW
HgoBnbm06Fqvv9w0IIkmJp6De2A4geSurfg49TBZSuyldPRBWps2ePGtwWM/kJKG
ANenFKrSFab9EZeidBZvneBC8heEaaLhssNn0rraoWVIO+KdZSyC0MRfCckWWN56
Yn9CiLD+Sn8mT/P+noy1o99alEEveWvib6UjB9/SspuAECTpQuHCxUMEr8RKXh0t
Bi4YrcN4hEUszOuBwfbMbG1o3ax+Kscs81qphZCUXThFE3rVXKPGFjBVJu2KDN+L
/Xri/SSPZ+aoAuEa+oHxwKO9zJywFchSzUcB1CcuH9+k8bJd096/iJ1xChdUw0aM
3DlOH7CJmvt2eUVlbQvLAYmZAISNYiibxCyXsNXW905j5mGTvNJcIii0WHghdmkq
59/qcSJPRYgD8QjdKfKoAG9KmwG/JeyMnM7YAuFPQ42v4PYQWUnXPM8QSu3C7bPU
6cgRRAyePF/hwN7thdcAyqqCjRtcSGv/R17HR9yTNMh188jWiOnE9ZwE6paNPpwD
7F33TVrH1zOYCuHzAGgX1WOGUa+A15tWHe5/1kUVJwDhtgNjgCAMwVah3OOPQ96+
wx7NMf/WTTOCDcTHSE3p0xtg0kkQJf9CHzoOOS6tGSnTAM2RtSKSIyMiS7eacrTr
D8s9kSFaO9DDQfvk1mPorBJrY0AoMdOLZnthM/d5a6sM0saOe5eq2B3IacBIncyS
XD9n+xBz+PEUTN1RcPwao9g9SLHPa3norIjC97W92nOrSSKxEDQwaLNtyabWGpSb
dhJRACHoT6gMA+VVZ1hIJsvs4Clv2LkxAD1EKEwT9+uTNoYMXV8aljFeam+RdlMk
w/jeCHUetJpUMnm0Ovhjo3RgVDPhdTgYHg69YxExkHENB0iWlp/ToExdaXirPoOz
sm/FtmUp8QEUAtZ4L5w63eXmoVh+n+iwQlkk9TGyp5QfCh+lvm/aJQ8VM0DxIKDi
48wQrKBQBbAQy1Q43kXMPhp1OfQYSYubL3Wt3hBlWVpWqseiUwUenmTT3XVi3Vk3
AnFg3gWV+97ZhwgOTOyKYeiE+b/BixOcCmDHfEQrJM0oNxOM759kzpwm9wd8pzXE
0uiE1lddaStUCSf6QxItjrAo7bhbWL+eRMyyPQxD1A+FlZTZ1hSbKAykx7oS4oag
z9kYX8mAQk8wrBQliEM1w5F57v2lWIBW/ABd05xfTzI4cIOCvoaA/4lmYeGRe1Ef
ernLGdEhbjc/mSKdbiHN8DB4hvJJhNYgRxKGuzHk2t+nfzKvrzASBHkJ/riedR2i
S5S67WJLSqE22ra7WqMSUcreS2U8qggpCQMlrcaecxJW+N1jBykZ+NEFFP1AJy4l
/k9jbp5MAJ1gkyqcx7VGvXFUOVPv8s6+1HO0+5bWq++E1v+msTZU7DZFSQ0Pmlb/
6aaof5Um8F/PuIciEBjwIFXEf3MjPaGUrJv0gq4iQein+U04qtyzaRhEuMnZi6ms
8TYWVPvOVRCdl4CYCFtzvx/h3eaapf00iNp9UGAxFfpzFL3bQ2zpx1vshbDJZLZe
OObN/N8t+m14H1gEy6ykSxgoLcSNCzdep2tEJhbcSBDXQvF3FwcrEstq82N7wpl/
XuJI+SPtmL/Ql2fkZI5UbOPVZhbXZlMXMGOvlBswUYRSN0/cnqOQOK0405Nx0K/K
CTpjoaR0irxqYz/5TVEfhvbI4kUaBB/Hk9IKOQnwO+Hoxe+QyynM0zeuyBjtkoNW
48DZ5v2uo0bInbD1T02M6bpwLSpVtmBvehGMErMqtVYHWoZwJrdJAKRjawImw6hQ
gD8fTjV1TzKJOqzX00PlU8Pqt93JZq59a3AbkxyIo1D2lhcH8JXW/tlf0moDFMCc
NrsyTw9CfAGKKtzUXhIWyr8llzKO1xxhHW26wkgkmhjX4e5NNNwgr31Pra0pABTh
DZ2hDYgI6DsTvoy3Ca/OiJXS0XdI6JkJbuhSH6PeTvHZvJ/O1iMe/ADS9HGbs23n
/Nhi1UuGs+MgbF67Kvaw6pTa2LoEChy1UnNE42G4/r4cRDZU+OfP2RX9u6NP/9lj
B1Ar7PB84tWB6Ty58hARoyDmEQHlD887s9P3LBuWCPCcwXcvRSPDjoVfFHKqJNIf
lyoLhOKwMHTl5SJfOOPPQXOgIDLsFWTALHe39eVlluAwk59XZtBxKVBgTmd1JE/C
crI6+d/WIt0SF6Enn0vu9+PYLFeGlWS2gIdUCQR/eBjKeEEqOJvpGaqh/90TeHmy
Osf7YUdKrErFzp2f3gNqPAWPw7P2CAZ0Tglg7zJdZfwzjqHZZOJRS4+TssQlskD4
+ABD9x7CzC6WnHWMLMeTvI0ZaVWoQmz9jZwIRcNwYOfskkxmB2uA6KWEaXFyxsAN
liZ0tDxVAms4NEi4yDfNE4VTnX7gUrBiesDKhjgI6ZyOa6gIerARSH87A/Iaddn3
oDKYrZwN9AVWUUwaSsut7Ai3dStj0wVC4CEJrfU83rkZrMu9VOVSYWKsEUdAWcpH
rnrMCuTJA2QZSR3baX1gNbk1BC0bATL0Alu0Jl5Y1B8/Fj6wFCUbg77mb9/IzULi
6abFiVRagkbgT6iEGXZ1fpa/LbMG2pF8tKxeJdTXNgzYcsMqIG4AIoZpcq5QSbgk
BC4HdmpBXXknmcXYyOtyB9CxpZHrgFSuGcNUxuCQnDNRDswZPiFeUd8cvnIxRFHB
1NN5IcYL98sAOilbXj2g/Z3wPPKZ9EeGbJnKBjMo/gtlmXx7pNySL2Qu69cfZ91b
6g11O45TYAr/dh1e+Dcbut/UL3n2uC6qNwJZDOMfGMrXDG3lqW+cAlD8botzalO4
qM+tJxl6YESIE2CoReqZLQ04Xo48Dnqf5u5X1IupFUet9i0RRsomrVPZXNCZT3AC
vv6V+7wWqecQcJgDpWoa+ycp5aBqL4nLHsqtAMw+4QX8C0ARPUtnTOHD2IrBli+u
j7WYLJ3w2k4lunbXGafvLi7P5YJU5akPkg621yv/vL6VegLyshWfKG2o0aLqMAwO
y6Zdj+IO+jTryOCgAuY6cv2QMXV9+xF8QtJVBOmOpRodX9hbLt5EREeDRCjfe1Nk
9OvWxgVYXSdr9HNNzInpLg6QWVSPqSBDVLjbyMHQeUmoyc1nqm6iyQSa9D5KRjST
L926VfQS99/H9G2rx1hTOhZKZTG6ugQhxSu0Cet+McftCG0tNpkNt/h06Acvt96g
VprBjplvOLCMiMHI6/KSG07UjeBN5bl0XULaNf5npTN2h33jqfbBs4fcNnANRFk2
8CMSzSIgBmMRmLaLiS2YlbJtizluRaZftQ5DZqdNRIQc82o4A4f0QyQ3I8yUu9Mt
LmjecGVDBwCpUwx2zVNIVCLcqVddbNz7/JRmrZelaYVDfUQIU0MDFMArFKS7Jffh
HHsTUXJRERDKGxHx2QlsLI28lvUP0UQtMeWvrkZI8y4cgURStQzpVSm5ikYFbVGt
YpxOu9nT9wCGxOnJnS3pK4rPM/W7iPQuXGuYcBVapCwXlIZ4TXjLP/lyGlK7bXme
kV2D6kYMqRC0YogBvuQVm1cPWOp+oQJElogArB96RV6Jm4QKvRfbY8AgIX2KSkrg
g503FCPnwQv3D0JyhwV/Kc/T8U8nozUgd3ww9ou9FRNjBYhQ+GzG92k1v/8ac31z
cVqakvVOl+eOtXWFdtZrzMZYaIg0GNT2k8zM2QnBQ9N5tsWkWxyIOkdJNgADNUO7
LCIy9bG4nhGQk8r+k2LDY+Hy9y7w2rM9JnEPzOYCwmg2bxZKq1ryTh14Bk4Q+GXs
18ML0Wq/DY/st3GLmF5RuhbkVGl3b6lqIlQbiJJ9QxqZkJHZRzR8GPR8qx0vCH6Q
yZRaAsFvX4ZEmQmX7KsytCBUDZbq4MCyhOCp6QQm1O5dYIzXT9yrtFaU43uD81pI
ATpmaaZWxc80cGyRdGUWH+916h1WESzrGFEfFxGhlwwApzIJD1+09+CyHps5x0x2
fKiSRxMFvNdlhFBXA/14bkLT2NtddlDAHpo/dJkjEAIC9m0ZiD9laE8cB6MJqjKw
iow+U7oPE5u3akPGu3KloYMXmhb/gH0WQL2mdFm3gaaFZ3Pm+Bjm578P9mqoORTd
0YDLqXsyWZIZTsDVDJ5Cn7d1gkPs2ISH1jCBdvxIlx+qt+gNZZuwNEp+522JDyb+
32v/YrgrELccWfPlpFI8ivg3uSrx/E7MWzlNO2TYRPF06iFTB/5P6+2nNuOYzSQq
YRPJHE7VmJL0+yS4tRdGxkjwAYsUVnR3ywX/16EN+dbFYThYfRrGFV3pkXGJTdCe
84IVkK7gek070bpGaytqNutuX+zCHY1duF4MYpVVgmVzI7b61DTI9H7kaGSkDQ9l
NhnGhX1a505H/o3bxHUL8dGG89+2jBXDivxQgyb0q/bZug4Q3itSEBTKHD4EPGpP
6jysKpXwsBtrR8e5xFMNuhacZTWOpwYEhicR3iwobPcOiW1wyeBciIMu966lo4uh
gIwQJ9DOE+6R8oR57tVJr1rcst/dRwdTzpd/2x5UpXihRAFXrJM8+R325+4KnVd4
FKEnGAP69qFjGYjY50sN08XM2U392Aa50ZMROg+vc/Je/yTkb9wOde35rMrXg0zp
lUFN9oBBYDfXKvAz+ApB12d0daAcUQ0nUNK/ijWHnEC7n//YbbKTRKtscnbqqiv0
p2fb0GkcB0B/dSEaDID31G690S2+OSOhkGpgVrHtcQybHKtm63sc/9cPmrB97MMk
hRhENa27Y/+a24ytrS5WoRZ+v0zb8LAbspKR0ZC4+CkmPm/X68vEdQXxgPmrFzul
ZQLyf5V8FYHTb0YxeQMywV8RKhPi1A5Q4F/vJNQyiFeQls3I7KXlVWuSZVjhaNpE
RnLTbSX0N5boYiGZuZwK0MDWR+2jXnftiis6P/pqhp+Gtp/4EtI11m+VVDGPU2vM
FqqeeysLEkD1T/OUDGX5SMAalx+55jlIeDMpi4qB5BXubCrFrbL2n9HQ5x1N8+ya
+aYgTEPoCKGbhAZMI3zDAkhYJyl2psdIMi46jTWVIV44Ct6hvsWefrnNR2wY9un4
AzWyP3MQnSzFGN4pAn1lj+CPxaNqe/6uB5D4TVcwNOmX5MIg+51VpclSELq5EtKJ
sbAipMj/wDq0zW97KM2d62PCxZnCWIJjSD3ctKkZJuQmWOz1xTdhrJr1RpHqTWXz
5y72lzT8srHWJv5+m3mT0PRa2zzHEiGjRIs47Zj9fFrcCY79+yAPtlyN1z5xnPCM
g5zi6CIO9jjMkrjfUBHqtzTW9eRaz3NBFvMHojA8unNbRgYvVswFkanRSrKdKDED
Cz2C6lpT+ntkW7P1vIGDwebD+4fnp0+2AsmJGFdEiAc6UyfL6EAQJpLQD8AqzqjT
KCrofY0RpG3mOM2RXAnSpLGphak1Tv844cY0pN+142pNz06RibeyzhP7sZvedQ7K
f9rF5F0flHNvsPd3BHGqoeI/8+xXE1iby0+yrMm5AuhstulFjiRsCVdf3T5DYCpp
9sbF7vj8btt7SaCmkQNSLiaKnZNANuxQWLzvSTCIchRZlz6ChDG/SaGJDJcwPSe/
6j4+VwhC0iu+eFDx+NXi9vavWECCDra1gSDrWk0xZp0kI8wK++fKGXbtzsm/XD28
FcVesypkg6Xo4NEqmws+W5TLS/i3bKIdHaroWUMKlXT9nY9ZXaIs1a0muaIHPVt+
ZdR3aiFHkGs+EJXKnRnkwIX6kOv4D+cyWWRw/+vkFe69PFEpTaXf8+hkXeeAnB2M
e8U/xbiCp/b49wb8HVzQmqWevd1OIqeJxlYPyigTit2mYrR/GjoWly/f2cgfNVt5
aldZUIr6cH4XVptXAfYBWh2A+mAOsJ7PV27Nly1Zv2TfFC+w1zmBygim62LmXdDk
pmiN6t+4ZhXvrqR98k9IydgMBv1feWojnvgwBIMc5+2L37HzRnpdNb2FULEt5cPZ
2ffrTz49htwBZRu1BdfJm8nH0SkhoEveEP+x1cBBtRznPiLY3sWbsR5tM3R/aIQG
TQwcvCVED3neItqdrB3RMflEY4k9qXPkBupfYi/I/E0AhdRtXzOBWHOFqDvouryS
wxTTy32/j5lb5RjqKURUQ2rd7FfRPUqdDc67aKLx4KyPZ5KPzBdCjWkvIRlEd/ys
9a8J6vClvQOBwQjn2+INp7P7k8VMKSjbI1IRge//SJqrHJvNxbaDgJcWNzjsG+GP
5FyzXT/qG8DhyYKHUogKklyhFd0xMg9Le/8a8wCudiSXWOjMeCcQlCKQ2ZolPxiH
qbfs6Sfd2hhPIF8VKNJ2Jd5qWM0SCFEap8L1nakYFu262RhPUiW3bo2ver3Yumuw
XuoOdOPrUA/rZAwuGCqUT3oV8y3yRDHTAdfzDh+93TTKaT/Lu7N7nf84Lbbn0Dyg
lC3CqaE+Ot+xXxE8Dg/wrOEfjGxD8L+NL1BTBjrzepo5wRkBHrEvPTzgYjd9mLcf
VN/fl4wTZ68zRjKgLcrTTBBtkr6Fim5QyFREWO585TsFmPWohk69f6MePnoUH9hj
vCbk1mPtmWiHqJFcY4l6/HsBXTBaa5FCBu6IB+rdOgU5qlDAfEcnVXUR4VO1/kKp
Zw6H2D+gDNCCTovJZ9dunVWkRrja41lj+gsANr3EsQP4Qgf+Qo1V3orVJdqHxq3L
CHt7d5FP5dlfxO9JeaOSUvD5k00ZDmpEHO0v4WDPVot5zMFAfz1QThVPsZt75Ovq
OLwNG7tCoEl7vH7WNkJGpWMfwh6u0hVcTZvHfz/Xh8eHNMul3f+RAKEJ6nvc3tDb
stL8SLgTIW9KXZl3K83/XwmP5CHDSKhT2MR82yc5sXv/XINaYhgmHPKqx8zPXdOB
tEJEaB1pjv+uuiUpvcnKFqeu/N8uvT+sckCech7MBw5t4c7N3iGPz8kSUOXq0LZi
PMiSww5bw67+8LR2+MzVtoJ7Rt0XyHjy+yAQQbbVZl9Znr74s3qN+iXQwiOmvuEQ
0ogO0sA9wetBnNG+idoXdAhFlWJLPVH0gcgpa7Im2L9aj2WUAdGQmyqvBldvaNdH
dzaLvR4Pvh7+Qzwi9dGRiLeGdvW3RJPTbxz1kOACVI1venLrp/xsTVGceuCgknaT
DcI6Z82LpDvNW1gc/35ccbxlBjrLFbnk8MEG4KcPUUqd7BqF3vy9vmrPRufR+PlW
2ggc3vX/4fgClZsvbHoH75wZfNm25d+Te1CcnHsMP9AyFm8bE5kfGXXeUBQ99yZP
RcmQRfrwlyY8G0cUPH3V2sTEGJLB9QfZuNTAl/MjzwulBuOnMuyJ3iMuW2THPqYF
KpqKp1lH5bvjf26zLPcmhSprkQ9t7l+4uJ6cF8AG11HxdqXQtvrC3ZSSvlVAag4R
D70cSaCwJWzjLWm1pdNa1SgYN26Xg/PQB0dI9/7wLj9gqXAINKMYXUQp3KmvSmd7
JC+z19F1BoqXsfP4iNPQgqYfoIGLavDxDVaNxfjHVmwjuih5uNbVUZAxqNmmmNl9
qe2C/pGVabkawip7jKpR+KV5al7X3VBm3XsEksggKhAWq8NgsCzpuW8HZarKMoeo
Ai3lUVWnrFv0brhix+cpjP9MTvY6zb8t6HYLtBM4F18pZazds6SnnSySrIDJQZ/y
735SfhdP5P1I61olQGyTxFcmC31oXU2ct+f2fIsTsEstLKqwUYQ4eDCoD5yJObB5
4JFFkhe++YiybriHQuryH23dyy6IFOZDnjWzhZZON2ILVp4s3xvgQ537jm95Tg1b
l/Fz7sikINbxm2x+tHrzgXeYTsOSwA6zD4D2UjP3MsDRQyWkOnxZLUXkeMNDVtqV
7fy7nWDsw0v2kXbAUH0najaVgim0UJPOXzuisFdbnLASN/edhCarJoo3Vaj6QNSQ
UYMUKbUrH8dH94MP4paLQoBat0XcLtHQv9+aMHybAZIE3+KL06Jxlug0xB4iLzc9
KluR2TS9G0YpUfvpzXUOSg+4lp2B6/vfxpz0To2dkUj3AJvlrEtczlhNlBe1JKxP
0tGAotnmoJXJUyCxgINK/p94ee/OuQRw4MoCfsvSoPNEVdnb3JH/y/fnRsh/wPK+
bUtX1dAhkimrElAfkjGkqPNR/EVnxiNujVesrO4QiA/t215lAdWWZWs6TGHVA3ln
/+yvIJOV3+EoJE1eBdeykxpUnK/ZEP/452KKIZr7+um8v5axR43AfiNmFlGUcyST
t+wJSi7r7pDGapuWXxdH8Cy6aE712syCypzPbDzrVxj4BaxSppEvc8Cirvzm4+SJ
yyV7mLbo+bPJwbFC5CuF5EoslZ+XKJQUfmEdUYvCghdPRDqchNyVVWxIhIJePDYS
M7CKWa2+l+19Tnk1kGVTivFsUiQ8Tx9B2PLLBvWWkOWiLML0AjSOJ0kDHAfdkZKq
ERo6Hu0k22/rOsdlLKvLerbbXctLctO3FsmNdZcv3nc33/J5JzK7mW/gFHJtgCLd
Xht0m9SLrqcvJu6PMiQm0DwmV4FDh99tjwiw0pDsU5zz4LANcdzi1TsWRJ2/nVI5
x8LYrswZW9CTgsuobIw8Jb6n616NUEOutsXT1M8xPZWU6parVT/BxP3U3f9LICoI
S9pTyCh//KxWhs0IH6kH13yFOBHnJgeQPmmfzkid7Gn9J3+MPOS2TOJGmRzOJMvK
sftt9k5zEehelC4+5nErm1qOGi7HRYisxbJnEokWW3uE7QkNL035NBZpa4RhZ39B
HPofRwTJlo4B7+/ZNSJ8PUtsAeW37a2oOem3IopCik7QhvG2f4Wieha7jicTb2eB
r8K93DrQt0YlBI+bDVTHggkY1heGtmvcj/XkC+/IW98VBHJzrJubOiNGVwmbWTMg
CkKPHtWWe69ah/um6r4gsBJtQsvC65YxFz20gezfFru/DAikkAaf2Ncljp19UowC
ywzHIdRg6uug8HR5fZAV8HQ92g5XSVkOhlUDmXMiC1g9ITcgdNRrEF6hvz7Aa4yJ
fim4Vpb3ka4KWehooXO59qOqS5y/3zWqbZif9ge+Y53YLEOu6QMyUcoFx0SD4Zyo
LiwwwjsfiH84KHkco6Slk0hvBVB0zP+vyp7QfjmFOJqF6Oa4yAh3a7kyTF0T1m2j
clPBH34lMRz9Hx5lw99/lVKI8VhXPyXn5g0k4/PmapdfuYTP6M6m+sITp7b92Wyc
MZsTP69o1mzk3WgMhoc26zSng3AuVz1smAgj6nakGTdmGflnc5kCGR8DoNP08k7d
8DcXbK66ntJ4SLMo4/+rH/tUEJ7fz+m0ByGk/i9mGtvGpKxZYYo0aQLZhYTAFwds
cBYPuPi/jmYyK9lu7L97LNL4yp2qg/OqgteC3mnB2TebPJwOn5cd4KkFH431iUWn
qdqpHzPUJRe4kCLvggwsdG4u4UGbuo2otLChoFzADpaAalVbTDrKzc+56oq1FFuX
7DDQCIbX3GtejRf8rS4jYF5/vHnQLcT9X2n+YezvuKcFORPTcdTPvLhDRClc7lqn
w8iu7Uoa7SoT8vQdnIQ8rIcW0T/QuwucNEooUx97KrQi28KaRw9QSwOZWBL4xNXX
g0du0+AOWIfDDquub1BxFziIRw1JO+mmz6qfHmxUP1M0JyA+1NQOxJvlfXZYog2U
mLmLCIHoKdtSgHyZVvib2OZoaL+j663Nyt2pgiWob16NxBemEQie1nFX5LhWwzqv
uEmfkh5a9+OTV6BgVCpn5Fgncqv9KHq9FbR+QfL18v5uw5rjOKV+xvkLz/gsdQV5
8gFw5N8EFGY4ogFLc1dYvBn+KMqDosvUGp5l0B1B9dfaT+rCd8szKPag2XtQu0Ze
LJmE7kea++x0RorkyAXp2ekr7/xJFo8mqMVNBElaaIteBwdyeybteryBJ8jQLrAm
giJd+UPWkb03d7BfZIZUYRCehh2JsW1hDmTSntmJ+eWw4vHh7LmFH62471RLDjlq
c5FeT4H5+33g2DCV1R9yw3yFCTyc+zX0mtjudEgeSQL8/tKtYTJLt3uYKD5+5laK
DGdpTF8f9paLCWTb/ZAreVVpNrZ1qV96UbSeJQWxiv+XzJ7nYRia1feOmcLrBAQ7
AnFDcDOw1alzmJGcnXCSIOMNwE35EahNUhE9IXCAW6OxpQX69GQ/hrY1vp5W+YWV
CMU0734aCZg1Tok+3Fm1GUZTYmdNlcF5WheVPCdQ7k4F3etEksvAe+UtVmPTl3jb
gdNf+fBi0luKbDyISw6mWHyziZcMJvi3Jh/SUQoVfz5JHZqVFJ80BP8nh7orvgPx
S/k2nTKhr9hNXSIqqIBIXNwmpLQT41+K2sX1BuaYX2mX9bTlobfRjds7Za4qNhqo
6ncgBOYd9/osCb/myQR7I8GlUKWzjcZXme3vDh7KLtj1QDmaQPjRombt7OhPFgdZ
h0LpB4bfZb8+q2O2DvHn33HBYaMfvDGl2X1wq3PvcQ+LmKbkFTuEsibeEXnlFQpK
ukLC6c/kYE71zATC9dAviUcqColnHotoYOWy/XjnpTlHhBgxkJ2iSFrR7UtGM/2T
1fDyH+Wo+HjeuF3e/9epko2o0axoqQm6YA5cIh4Vfgx1JeAuO1WkfucssOorIAle
ZBQGksOxl/ZDBBQQ2mmLn4FIztEEQ4K+f74APmVbXhp8AoPLOD6DyiZ4RwO7jlLw
uUIfI2BCeRESE7XN0T2orpIQq3bfJxGFt1J23VRqRM+jxrDqIfrWtU8l5by6Nw+0
Bc609X38CGXNPOrXHPnd1w2H6uKSBySWtEEt/90CXj4LqyYCBmN5uGvv0N1n2bEG
sPlpl5uZAsKW7fU0S+PViATY2l6HAe3JGu3ih+HGPv0QltD+MM2N4OdPIADDIN/s
7JvlvhgR6ZzRPYu2Ki25Hjl1GZxiGUEh2jEJv9kpXsKjbAIyRSfYlTtPPamP77rK
mMc1/bIqw1qQ2w19NkL4n/FRt6tgWaz3CtnxhYZl4s8SiUlHRFzRlzgv7YAnZir2
5dFLFZ12zg8GOGrSX61f/H4aTvsTeqciSUSeKqd1k4G70nUYmAIqEriTqN/nuJXq
S+5Qc0864QQvL0+PeGbsCeqJhs8ms5r9KQrl49hatJ01A0PKClCQ5mik8ZnX6Yan
YIe0yYvKAXgN8NZ747bo8GE3sjxCVxxGScLJFcfpnUsn+zCFk4tyutCUnBVtlg8X
DVYsYFt7+w0ouILeGBzT80ra/ujT59jYyWtz7deJGbxMd6J4ytHPVvCDZu7UW1+5
n1F6vZhB/E1P7QEJAuwG0nCNHwFc1CR77B3ic1bRBLtupCj0wRs22nJf4h1Etlhx
Mmaxw6DzxRigYIqIM+9+6Yn6LFTHr+SN3ZMtiHezGYZlL+BPYhd5VpgTgCIGYQkY
4ZFpkYSGnCD2ljBovN1yIWSNjt7NWhzZyxrUskovEDGBwoofoDmb4mmHwsViDIO/
RXI8e/ROm3dRUBWoCI5YVi+AzzbSDDEmyKzuMYpTR1PtzzSK1XgcT74JbFmTXSwZ
jcjvwpNG1YqC72eYAQYdw5pAoFNddraOJ0zldGrTX8NXwPN3TnfzzEBSVQwkAroe
NtouWb2CsJKRTGTLQ+cw+A2NS2IY95FYbVmxrK8XxVCluUCS8eL5AytVoG6LRoHR
neq6VWZC6CPpAsv9RyGO6CkolIQEHnFxEKleVdGmsFXx5c3EQWAaBXQL7AIzUB8V
yTGp8hgKKNPam9rc1GIhzFzDzEdj/Sl2CgFDN5AgYIY5UkdK2hAtbOXxG7URn67i
rnP7NyrfIzCPrhdeJ5otRE9ubYkuQbES4iUccikAlwxWPgw4DQUYyZIzTvj2z93d
aLtgRQKkOvyzsLeR4v5dSA2ZXhbkHXa+hlhmES9UYqUsaMpaF3eh8Ep3j7nEdCoy
lX9PFMughaBvm5ujOqQq2S2Kuls86HBGpo3WfrCuL8B49fjwU6cLE3xLmTW7sU/m
i3rpdSppu3aOhAe/bbog91l11g3tYwCF5sqYc0Knk1zuJH2NSbbiFkdAxq7CGJkD
IVpqOrj6R4sA6A//C2KuU1iMlEk8ew/U84CI3dh5iyRk0Gy4a0ZVX6BCE9iloP6k
7NmgGUIVyRzQU3M9J73P79ZaR4MvtRa9jerYQUdhaF8tfEVShUn0ijjUq46TXw8F
0JdI9O8r381Qk3HDXqQAEaCB1R5s/BJJOykUTvAgxnVio6QX62NPnLe3SWXtgImH
eC94aTAaNmSY7/hrCSi6udGrA5x95ihgIBHOjJdn69NuJyo1fOVFjnBE4psUrVwO
wjdxiwNqa4wWYG1+tQTC64ukXSYUd95DAzhy039dr1I5GlM+/evcAhsjqtNdXq/7
2dcU9i5tdazKu8CpFx39k9rE80u5x/6MmioXtw22ZtOqDEMDjmRAfxMsLNqEuGyk
G6O+nO1l7AonPdzZUYGMrO+foujvJ2bucziEZJ6sIE3y5HY9AXfRRSHjlBzRc0+K
/mpV1hVic//apd2s72b2/L+aBmvoFjVQG2D2TKUWIJ+cmaxQFIDJKcQx/ugU3p9v
y6XL1H6ij4ukEFHfQ9ny3saODnEFzeen3TfJbNha+3pQ9SkCEZj/XOVOB+qfqYZQ
i87Kw73ODIfZf9XeeAoCyLztao+QQRqPQvU1oo7RcdHxn3kbBYdB8lttmIucS/ak
LwkKVw8dVFdvXNcuQ0prDDb5e+A8UCHkkbQfiyF7SGYlOwEehMS5tOvmN02dU0T8
qgFMRoY1hUbXTsMAHtiFVijMfXalWhArKxfkNY5hY/gR8N5G3Y34L3d8tTxoePgs
GGFgKY8tS4zLWqwytiTXWDTWrRrgUvM2KJmTAkWANr4bNYcHpyNHA2uoaWZm3LhU
IO3dnCyDpGiBTz2FNoo9EAzw44a0ulgPo5KyXzYVmN2cqefcHIPAhX3lliwJp/mw
bKpBT75mvZhZxiR637hE0EQUDs5vwwxyjOToebK0p233LSYqK2OLY8KmDaOiWDdB
HPmrfIycHwREHzfV4xRAc7morZEwbfiiPHquV2yOuIP1DAYLOiwzXaJaMNbGduJm
CtWUu+oGcDCjtbtp7iO02ly0HuVDfbgxEbiFoDJj62l4vW6/8Pq7xXC9VP0CutLO
GY6cFaZB76zuXqLrA2oW3/P07ErHoaBlk2jafzfAGve4OCnyBJKww6Xt1vL9NxS6
6I+0UqxDe5pO3dgqHzzSjd7n2yuGVDQ0aogfbYUcEz1IQx+s2KBeUTWUz8KXJsOB
vFmE59bjdmrOhMNVJCg8Z+BQtcyI89j2nuAk09+zVUR/zNqtBbq9mzqb8AO89dGV
kmKghgb4YYH1l/6DLjwmZigqNec/L3u+LmLqEf0gj0u1uk6Q8PELIknQtv7i9enk
ZJl2aKNhlq6Od11mUt5ZI5lUYRYFKWdiLNqBXih25HFLGOddvthgCSNkXqbVKiuf
S9fHmQjTP8gtIEfmTNEq2EDaP61bctY7Cx0OfTQGHBwshpK2vq1ZUexdfvxFdrnj
zprLNOgEsf6qcE3Q0U/5OAZcjWDotM4tIrIL7KFLYx0qAfzBWlLcTkDPV+e9WZAA
e/KiIu/u+xZuR9l6L9tslah3WWIbmCaMRBJE7shfsfObTuH/sxRNi36+xaZOPp6e
ivN/Nb7ThHgLyuiCn85vljtemb9aMAfu9E2STMXmcrz/i6tTmB0lY6KxumD6vAzX
uPK3/ETCkY/BShcn8xdT0OcnQNAsnqrjpsawNhw7XZLLe1dviGrN6dlRZoYSpgoi
U5ma/39nDdQ0+MRR3UCsjoxJuOP+FfQMu5mxRUCpMEhPari0sPm1/KJTO0ifOXL0
eizG0jGk88AldX70Ch3IakQQKixl7RHqboG247vUybK08YQ0NJ4diWFFGilD9OoE
SSs7xMHMHX1lrmDJoGPkyjpEYEt3MQDotkIHbVUnwon4V0E5xVyMf62NEII0iHpO
atKBvO7YjfPCmm17/mDmxmDUrz879nbEEizddwJwvFd7gVjtnQnHTorphcLxLgrp
dXlJooKdDXjliyHrai7cpCyHzdSd4VoHilz8esvPUV9izB5J4EjS9xS00XvcnYXQ
PsohhnGcs3R0zFzxLuHz0aNdsATl4RMOaU8QU1EBSmqPDG3xjGMZKYKhgcOsTvDh
2yjL5jYJP+9cuIZS4CiBWCwwjwibouiUa912xhYEXWD+U8r7eWeREnuseY/Bmax3
Uq8T8DO65tUrZPr6AE+OgyHfFNTFX7CXCTrTZPUBA2hlYoWlNCaz8U0slEGGxCEP
FwbbazJfgza1U5BgqyRn7jBn3+XsgqG3jeJoyx3NA+R4P3RJCP8MVBhIYjYsoSgA
+x6q3KFIoOmIm4ozrsEZYxsT3fvZRxEVXJSdQ6QSDn/ZYLspFHVIwSsL0nHjVCpp
8BdjeHyOeJ5ZIk7xVd1/lzJ58dPgSLhZrr80SwKBqOdwSoJ9O4/vh3LfjN8JYAtQ
wIwJb5owptlLDgtNZCfvJv1pi1Jbrh++CPM+9lZ68T9r6sGoGu8X6RCIzY+MwhXv
MSvbqHMDtG2r+gbTzGHLwHyR55VZ10KFfugTNi5z7Bd2UWSLyqhk2EgGEwx43ojQ
iYKo1qVjlxWK/36in76UN2N2+ADALWZjEhv4Ig8bNoIvuEABqYZ+3/FccMUhEghi
oKlaClMqfOBywzjzduHWNPjavVj91Chn34HnStrzmngahab8xmzJ/NFw1a3hBRhj
JTKyUHZbF+flJ47diPGjNU73i+Isd5lUGCbZZ3hguqQFasWngL1S0dM0L8V1qvWh
+Cy1jKAd3Lbqnl7envmpuxvflPgeo6l6pUtet0o21nYsSsy/c+dFYFlfWNS85o+w
gy+Jberom1jydsDoG8DWkHBQQ3NYSUnJE0cPSf8A9nOEL0xEiseNJda9CFu7cI8M
poCcWptbQuS/UseVLGjHIMYVaw+VB5SRzI0xZyjS+BDdWeFIDuOsJTCj81b8VZti
Sso1FgSW07Gre/OpoNhIBc7+W/ZlYzBROAxjq1pRQJ7VOc0LK3cQOcxq+ZkZsj1I
wn2xewCJgh081hMtGfx1zFyg3D3XA/voYkhoD6PBqvtsshPiZ4OEo9ZnstweRxBD
hZ0So+F5xcvLu+ryngxLqPCcz9wq24YjRFnvHAlBTxOJU9s4382anVaKz/lU7faG
aWEmWEsnP2/LHCIPZ2MpB4RQs1ltOe9ZcBfVZWGd5ZKFMjBBr/TSQanuIh2OzPA/
dNg18AJZEEwgZ9quM1C7OT+ocxTDjFzC1lEvH9GtYOhxuLNtypCy0Mw1h0gPYDpT
LNUC/KtreikN3ytHZ3HZLsqG1fZl6TWSG47Y9k7b2kYHegdQN8C70iJ/iVlhMkGC
3aLorv6J8jjUzjc66lc/t5Poox2YhPC0qyRYKp6D5ojRz62D3/3CEgEHRAMPRmyY
EfceYp8lPXPr5+wfvR/FtIhGLzC+etok5qD++Gy5I3HXmiZzZS8w9RYqcbmujFql
zQbvlTxovzKyuVmAc8rg0T/ApIuMnaW7u6T0fvAX9DUpT2g7P2FJGBjuioEv5jNO
HABYWcCYDsMGSdY1hcL2OcIqWa3ehNXLdpcTL7MMSc6kKOr37Bre/HjZuSu9F7Ke
+ETpWGoQ6cwJBle5fcYy+ZXpbiRi8jLsAF1L4JwbYtqirot372bgDhjOzD28nAgk
2GfWv8YQ5xbJ6ue7YNeeuucGrBEiqhK/qncg2d7uJezcYLUB0XFkoERjiyA0bwE2
G9WApj+vgE2K7PFIbi14zClRiBwG8JAqFuRrwth0KKSPVzIkIZA3n1GssPvmF3Xq
jhZTNvL+vl0BB6l00vT9Ekh+IGO1ry6E+Jmk0s4/mAlwGxK/GpmfUQLfK5epsC4B
JzFl3olcSuveowEvfrz5j0RS9+X5xD46kSYfYZb2Inunvy7YmJyUQ5OrQ/WJvWHT
IIvpUDy60P7xsUBplknvsGrW6ZHhOwgu8IrKKRi1yqxdRMOq1OMxiby+bXN/bvwF
6/VOjbj+Ja56et+rcTgeYJBbr3TKkP9Cw9m+Lyu8l8jMaOx/gHYWHxq/9olua0aZ
80UDmkFPEqH/RMAHXO2yWSR2zffkxmk/WJFZhNESnBr50na64eF7uvt8T8V/rNFQ
IqAP4KVOKuQj8GH91uZBb1tk5nqZQlnPPfuqMfrRUoszfq21+7BCveHD5ZgRMcTC
Z/xswJki1PTzUIeGiK5oehnjMCmtJ8ZHpRG5bpJ+1CMJo2whYhaMV3r4z/ftV9jy
R3Iq2+bRmG6LB/yTWZIr6gOs2XBUoWjFoqFo2cQWteTlT7NbGjwCzWudBxakvrQR
UVwoMNncNbx9pGBTVwztGh2/+SV/CKpz6wuzZQ8HjQRVO8icRX0mME8p5PxxMFdL
fpftvj9/XnEIqRLxZp+6PM7qCNNvRiAhlUxS9tIaSkL9K3XDEJtSf7yFwT8+5pRZ
w5wxqQv18/hAvuSAvldJRAkMmPY9IMGR5tYH86zbGSJLPBwEClGe/dAuxzfiqBtw
OlnliHvnzU0QJdwzD+ny9vo27nkRaSJFtKCJ4kdcp8i893krG3HJIJrCKgcnOA+s
82UueWY/WG5adJsthl7ZcJDp69qp0NgtGhiAWDdESMirde8p1gAlqaAN22TO6FRH
fbWlylbi/fS+09W78YPQU4eIbUN37ONnOqlxrWhop/koWPUPUnxxEJ1nxK0i5Jeu
TkLYaB4uL/lg3tVX4A232QMiGFsb4PFammlDlAwfLVkGnEvjwWI7KuQ8AyeeTgs3
7cbkjXNdHzmN7tvcuKiv/g0yUVu7me6SqbZDnJps9XjhBeVYIWLs1be9p7RtJpEp
bN8L1rWJOdKQ0l2Z6i4Lu71gSd5aF4/e6W5ux3FqGPQfQP8rZB1PcNqXx/j/4Nhq
CsmuYcHKjWR69hIAK7F88vTVrSpM978M02LkxZ566c6ZsMq9mdfZDhwzneq5N8sx
d9NYq332iqP0dyeX1LNqDInYr5mi9tY2SvZJez9FbQo1RItrkH0SxinJ9Dfijf0U
db7wtzH1MzsEezsw29++E+W8E2rPmm0UPeLacd7YdeYC810yScdnRJsai2MHLMmf
NcM7nHU5ulWV4dKL62kle1iiY9viPUKCb/6/FC6hk4Mzkg6stc3K7lgEZ7DU6PZ6
0Y+4cgJ8E5AzBa58rMGC0DjdTPQzhz7jT3mCrmXDXZCrwdzi5tA3vu13HWWVRk+j
R2YqH3dIuJQbdTQi1+2AcNKFd5heQuYj+69kfr4lhKiL8lppE9ml/dIGveEdl4GS
Zhc0CKtXE3rt4Y3HH10ouJ6jTeyE9HO1iRbe4LGIA4vB9mwL+9q0FOGpwvMnUWM5
MINEmS8ODNRIjYHBls7c/kN4Md9n9DENIULYr4SCkAg3zi/MCYV2M8M8rm0BOAN+
a5Wg7nwdsFf0l8ErtWIkZNAIBIrZXH/HkxK6VIVnS5JY9QXrv7i8Q/r66BcrhzId
YHV5iYt6qR+SzOMDBM0T5ng9bLUIhYnymqpdeJdeslUJi+dvYN2j3rIUhi4/l8qV
FwhUPaJvdEI1F1bYuerHBZwsFDMOqd4cSXgw7kFG2+LILEF9hg4LbyGnehV7wtT0
4Jp10Ywno62pVmD3wprOKRlyj5FUO8VbLs8Ag3rn9Fx3VeVdU2qidT0EFcazuLQ9
FZ7XRY9FpOnuHXvdG99kDFpK19Za6dkPvausZv8AKghz68lvLUhfAz4v214uXpHf
B/wzOuJG7HFZD2cej9ZWDROCvJk1LuTvFZ5Nc6S4rA2fPE3FeyrL3/OhZwMdjoC+
pmt9CxA8rH9tf4x9YoMy9tK5U/p3DJiqXWsQSldnxE2anEM5P3UmSyGYxS27mqTc
MWaxwzwZFhCrykEccRkjxOV7yEbPWH2053VvGRvJVuutsPqdIcFZkJCxU7b6qVG5
eONu3hnFEQqjcq4aGAlFvioRUSGBo2VHkRabJa+SlF7QFJDjc7rJDb49Uynf76yM
SUpGDXz+vvuBQOjq2gDI5iYf4h88IsyFkOk7qaQxrIKdu4DLQWXv6Lszcf1UGBr2
q7p+TBGMsNM+VcRgk1Skv5XyHueG6TnF44E+OSMdwwGjUY+qzuqavbVT8X6TLiPF
OxCjlZZqBGYVOSdfZ7PthsxZA6TmKi0/XxrK1CcOSYm4CPgQmIUCIcS5qf4P39Rh
iii60N55J8dlLoqQJi0FaWLBAOP0XYGUMra0K8mbASwn9NrzQTu1vcZ/IyNEUlHq
6uYdyWznyCzUVeZfFEj1U5IImpwLWfrG+kiUCLKfrSyaNyKc9MRvViyEMf30hBH7
5mmQCaf5ZpT2z5yVkZndarIo79rRmfUOZyeWDOdBdpqvbFxe783IHUF3WmxIhxG1
3v2Kzh2XN3fYUFCBkcaQgH+GOhaMTgraZpDTix72sV02luAhpYPp963+rqWxmJRR
JkE8Am3w83iqe/a4s/l3bsoF+dP+UkpOKlN9kOMEVmIdVQw6y7vsp/0iPV2NNEwr
fWaDYywWH36cf0nlGCv18+FMJ/p1wsJSATuV8czN0xAnCyYbZCsTvW52hIp8A/dy
wnM0Slnamp4K2PyUXzKz+bZ+zMMsD9887p04FWlh/mJ6eI4MyAy8kbHSGbp5/a5l
dOFUeTKr2JTpvBf/xepqNeKtp+07dcAVN37Iv0I0jR9QJnl5QyP6iw21OJ5z46tG
9zqUUiWBTFlf0QCCoHHwa5lphosoX4XHzzkf9n3nNN0eyU9iwKiZyajy3UOa/6pa
45gwttClWv+r337FFDVGyhistjJlHYxm5ZBMi1eWEN10CsTpSSLIpQsotD0GIZ/x
sJhSHJXzGX+pE+ZBNw1S6v8mxElH7VHi6075AcHh1G40aH6tmM6OEee1jndD9B3F
rcPy5XWBVu0KR3qlcrVzG5vjsvtnbg/tnzzCv3H1oxtWqDQ5N3BTxlA3ioBW/vQU
sCABnh5g/SNRGghkJNZys6cXalYLud5RUCylD1xjL13lMq0KE1sPNH1wDp1uyD47
2B/l56pS+4DxF72LR3u4g0GLwMz6HR5Sg/7caPSgE9mBr34B59RZUEkY3zp5imZb
sIBbh3VEAPm0f9yWUWFBnwonEJtcocB/rhMup4tfGSMRuIHLzC5xfzgDpy9/nlqu
m3OvCZ5isTkJEsXBCj1oj267iBdAeCffPc1QBdrOyl2V48/OmAQG8iyVCyEQWiOB
4E7z/Ei3NPA2BkZ95e8lSzMpVP8vvCQ0xmeChyj++y2qxdTOOVGLo9MRj4nnLDLV
IkwJ/sBHIi9fdet9tEKFYipOHsOPnZxC9NPHT4Cl6Z/m722COlX7VW9t7sGjbo93
f6ZTtghfIPjdA+bCcUdIL0tlmNBZz6XHs4WMCMbRtORjakEr4M9nz/yvGZ9tq7qL
EggKj2xh9rBCz97+/1ycoWmE2Q7HhXGOYLiMfNXDElouuoJ3SUsft4gFgmoUWx5k
OYId03lkXOGAwN0rhuW7whcG6GolK5VCMNaHq74dSu7jz5ycV1gT3e0h4ZxncsQ8
uzQoPTkqeHv3K3TY2NexDm6VhBom6Z8Fxn/UcF0r9yaA28dtGz1KaRAoGrGv3qPY
8vrzIrFpi2Gp55hu1RRUzyjz8YkFwtv2we2hSTRaT32tJKgHjVN4/xUUNnuPh3wl
xQrehO+NDMFE/Gq1oyEi/OaaJvLYBRLMU2sD3nPIe840d1P/d8xRvosMpuXoXuY1
BgapVOnfMTdsP15LeoIdAz+LRUs/CleSh/4c0usms9HER1HYV8RiOsbaycesdxQn
7d3Xpqu3z5wkGo0EYWajLBDYQWV0S4gIVB7RoEPLKTRTdLIMKVcTpXrJjr37kCxQ
qihRrO2ZU/bWUJCbPdPsSQvebPydm06DxMUlm/XuNPRILbpkE/wvFU+NVDD+X9cf
5O//Cv7OakbTcdN45zIRXAjnHYYPJkxE1IweHDMlyexwU4iq72vCKj4Q5MydyBzc
819C3ShFdfKTeuPmjb5FOZJWqt701LWZQiqzgEmyG1TBBmDf+PBE03ynmQQM0jjK
qOvQ3A4CE4poqE2to/FA39RrSqmMpTtXzN1Y+wLaLc2MY0DZ3CfETPjSXF33OUn/
SZPLhJx5jgSqO0tv+PUDwOIrsHKJYFLyfeXIR3Pn4mmuKnhFg4bpjPXdovnkR+R/
ixiCurjSuQYQ2YQ9ZeggV/fCDdjbwSe6T0XgJ6buOJsPMOW9naNngbUWNWGXlbMp
J7ksMvQ5b6wgYtwNUadCxNN5RE4vbolFN6woy7pkQY7n3/XzAowS6Szpyj/HvgsH
b/8rOFs6QbSVeFESaMhF5kF5whFk7XqHe9Q9QTetjJzrX4kAzR7dNInlFrxPeK4B
634hqFYF4iguC9sUrnC95tgDN0v4A1wZAmglDX5KafV7n7dXghVUtBUkCMuv2iF3
AKdA64WXgi9YfxiJjjByulzFctRVQYnNhrXgiSMeKZaqvXR1QTB916XIgeooupy3
WUJUrs0aF5V58//uGfXxKASXf/tKx42hjImVsSgcAqCZ9sPM44+FdaUfiwYeieaZ
mHfKlzjRuVxzZEkAZlDyh0qog1EAt7bMQfnXpMFz/QIHAZnGa1KGiozB++syjLZ4
J+QLoqg5ovJi1eyHwH49nhzSuKhIFGI+yho7PkAhC/X3ay91Ru0yQEOK781lSGiD
Rkq3sgDj53FLvlUc8mxsbztgh7wZTSnGx09SC98RIUMp3qxT6q77d856q6OMipST
rwVlkwxGGO0K7VfbodSFvUhBl85dnGo0X84y14WVqLMzy8/0YIQCpphX+D/2LA75
mTa9K+WhWGezjzMH6RkTpjKrrAXNMHxc9yTDym6FYAxxpdTL1YiEyqJY9bRZKvdd
8rhTmFqicoQ97/wZ0XJcDkoD8myLep62CRzUM8vyPPMhFQvJO9ackWUmXpzf6hMj
4RcAjvPzbZby4VFcn8ThYaEk0HNowebjspzX0G7C4v2X+x6qbRfeMud3wM21NLJV
kM+fyMpTwtMMt0FcE5ak1Ubf7/tgW2cYbzlBYJCum7GE05ONT1EIfYFGiV7uTbiX
IfHTPCFFCgK9uqrfmDNmkK0nOllRCsZc4qkWOZEHi2QbiMJ3QxdjKk9vT6K+m0Z6
Ffydpj0T1sXcbdNqHSw15sUfHagi4dTIFuB94ICXaBIRBZh9hCkat1qpp9+hrprQ
eUQvhd8pQMk6CVSwP2c+H7ZJLo6MxcRWEoHDQUkOH5KC1fu+QdcRhOuvCOYSLVJn
2Ul9iROWxyDID8Ce/eqh7vhs9WtvjE+3OU65W1Kcz57kU085peC8vY5xp+uJEzMq
3Ual4/snptTsB50aEs1N1oEA1aEBaJW6b58T+qFqmmiLIIe4qH/N4XgQbDlrrH+Y
Je0XpNE35YaRy++wPqvMNdm0ZBxTJM09oFs7BHBypupD1mW5dpipY+/+u88Ktzw5
QT7uout65jKNIi24iZGqTLWMM75vgnOskqQXOWlWxAkJQCmV/pWqVM05lixB0WW5
uyIGk2Hzu874WuPUTPyB1kDE/rzaQ3wbP1BPrGy19A8WS4W8inz2PBLUbGOALne0
T8K06tXDLhrfIM8g4lVnyX2P2dBIfcEJwh0dQs+QefA/8WyodfBj5XjieyxVSxME
HPc1+8O4+cQeb/XbyVXhp998GOk16iHPIdpSFkoH+JAnZyBcgSUE7fwJoUTOH3l0
sDmeK00RbPMFpubEBzLYRNfVkLoDXa0VnV0t7/9OZtgDskgU/RR6swXgStJuBfSD
s6vDZByQ28KZeBrVYX6C2KlwT9xk+kY56Ca87xXSOEz1Wm8QtP8481K8iQZkVuql
ZEGG5Q8VQfJQYbvNYGEc2CFHbXUuSZ/pmN3Ykn/WJlS6U1LvkQgs5CZbYjRg5JN8
R7f9OOnKL+xBWUdllYnoDsklBRKLwT7eg6Xt5SYLs4C+reizkU5th0YYqPuK58DB
Rm4wUU0JR18vZG8I1kuNavWZ+DwgkSpclCHdvnaQBT/xEocAr2x7EYFvYQf3Ka/j
FYGefxMh38BNfclar2k0rVdGEe18ZCHJTjvQtL1E5fWj3jiRF6NCoa++HHLS1U2i
u320X7zyRNV2I5aKrJ6QLoppjfo8JX+hl4KSfHkuzgXXflEcdkCpbhCdvonAt6f+
yihtbnirBBRAtAQ3TywDlWvbPDrVKZewfyBaBftedW/BOewxK374oLjyoTh+MTDa
77SFStxRjimC44DMHwhR8BRShodGQfLNm3tF96lQ983j+wg85FWYHMxQWS7Kz5RH
g2SPimDqTlVcbV6gyWpz2qy+319mUIWaDLAXthf/WeWUolB9aM63TI8YQ8kCa0Ie
V9C1niiafLXkf8IHQMu3Hmzg997cM0XC4XbUAw4nJQgXGEDah+bWdst9Svvskxo5
AEpEzgtT3DpaRtnhhTs1sO3c6ogDLEK3uug+7bXHRZd5h5mcOJ64dU52LsXnZ0fD
TvAoiKHfN2V86zzi3tRTZMF451LLOaMUkt3KpgH4l0KJsraWJbXr1XJntw494xNg
I5stPIQQ+eprjhbYHrjjadukE8UWL3UU3YhFgU9WrH4A0pgFWIiXRjK5hxIIfGf1
sT+6g+WD9t0Qaz4SzYshBWBzMovzyWDnqUEyEO5IJQ5KhbQv/93d79XJSSEHZZZg
/Bn1kGxrKHIf0BixGtLR3d+/LIUf1tZZYiUYDaBi3c4z4XSdkakU3Z90Cb5ycxME
9327mJRbapyKOxlbllqSmFM+2puR14Vjax8Bnr6hL4JLfO0aGRBqOZuqV6B0IqMh
NUe3EXZ32o+ZBkPP908ODfoju39OMrPqSaKIC6Ww59y13vaGnR1lSzF0RCjtW35J
L/4vXDP4CvfFZ/awXhpcdRFmW/WLLSALGWmTzhhB2qIQG1ecb8tloQpxIbqXflIx
umO7PKWIJEjwaq0edLsnBdI4hlYzTVf3g/ZP/N+HWO8QbqlRtfi0b9Wz09WgmoDy
9L3PBHvkiT1oUrwo9Q25pegyfSsMnPTmI+xWUrqSqgrBZrZhhxVJ7E1cSqGzHUCD
Ni2jXFKveS1c+euKyn/WqysQmV1d98hGAwtsLASjAZZHl3TKUcHB5h/BMk2Jl9sh
L7lTbVMxhUrowFGbY4pO88bisZ4og0hrmqhx2YAJTjjTSj+y26McxDjvt9lvvx+B
WE4beKW+D3zXeVnwTS71RF/W55k46X4Pcb2LEpY/c5tCM+ga7/zZpAPnZdGgunYL
hBZ6EVe+zmNcv9rJy3MJcz/NwrT2H+c2VNeCzNM82b+PbW3FeV6w5tEf9zvOVWHP
8hPhYhHS+0C6w7DNUwyTxuSlq3zzSAOgH4lPySwc6PmK8LMPyUZp74AFV3C+HC1d
Wq7VUT5mT/IX5dsNIdGKNM4NZ1RaCf9Fu1gTpQOehP/FZ1mKGIsMUo9f4YpjRVrp
Y6qwcgUt8tKgHGMxEX1Ozo838Rx4GN4fM9iWMZblEy16Fwc2lOmJnHrJn3ULV9Zy
NThMT6GwuqudMu0NjzSZU0qpkJgxjaWQSBbysgaQKo/a6N1ZIz26Ie4b7eX+w83B
XUR/o9LLfOxc5/D4hEqr93n8j+4XJPaBKttmOCw79xm52OgzPYfjQbSGvy5BVMAu
Rtl5ONPabrf8drQmfXFU3L9XoxjQJoWV3n/nyGMmUlsoHAxhx+jsqZ07Iu48iX4+
IOm7TmFJTR0tx7qv2tYtoLWsjWbH/Tt67Nhd42UCQiYbJyrJYTiqv5HRQefVj36s
CAvLOPE1Py1VVMQsaiHwFvPUhH8vl8Q/yy9TOi3CtDALQ5BrzlMCVhuIx+N7zAay
lTgdInDnLm2vYBetUM8B9/tpl1/v22JHegnv/Z57qssED/PbH4fzjpZS2Zx62sMo
lCDIoea2//0BbVvB2aOjcBTf4YhMpZsd5+4eAItiDOEuH0pSrMy8hWtvOh5G3WRQ
63N7Ey5lejGtnht5qrUld7Edf8xkE4EU+y4WETeMmjSZoXAXc1gY0BdpNMPIKfWT
mrK/Aujx7gciyRVbaPLFa3vSNaPYNpXNlz05qKrOfJau7wH80HhXCf/Op0HZAu4W
+MA4JjLIsEAoXClBKM2O+b70hcMnG7vLIzEl9EQJgj7Pi4goJtVOnkd1xNyG1xCI
x0MPna4yQjCWUZ53rSGMFYyLqrAw5JvKk1DsnYhf6syUYqn0z6xvIY3srWpUPg+T
QV01b1maYGcPJ09UtKreqcXQ+2yX+i2dF60/KeB2DU92IHZYv40oSJChEyzCdxpC
dQlBKRHYTLri3qf7xcmWE9PJU4n10Aj/wIPIMNnLkUHr944Lw32bZdeybDbH8i9A
eSju58/w3k0IK8swDIwpmE3M4b3d/0TywQO7kL07sH190bfsGXqzN5bqOIt28vEk
27f3dmu6M/46PxicnEUEkJYaT9lGWar/A3Pf2m3QTJGRfio7D+ObZgTZV66Y62eJ
bcbGMp5NJSl4+wwM8ubrRFGIghCczhRWm2/P7vR8sptHuWQmuAOEJSCN98q5ctFk
GiCYyeinI3AfexaUDK6u7F2UxkDUGr4PijIsFCeHJUro/qqZl0qS1S9Mj8c/UKSl
97Uxn1RnXPJLGLp3L3EnbAx3JlerVRLKYtnPVd1H8MAIND9VNKVX+DSdTLMVDYzG
+IR+D3NG8WxMxAwhtDpIJ/XIiuMjcZEYpWJVWE2tIK2QE98iw2p46om/Q1QNQg5V
88DFDaw6VNersHGAN5HTjG8sCH6wO9grImhdXpQWGzL1jVqTT/Vv8x+ttpDNJeTl
Fi3guM0IWWjxXJDIPyasPD4DceBmLBoSJQ/gz/+KtlbZyzniA3aE4NJnX0xCkPLi
VIUZkWvzP0TMeHQvLX5mVU2XloB/CyKFAImbwlIWiqGv4qqZlt3iU2VLIqoVCov9
bdy71vPR+gucaUc42rK7tHFONn1YoT7UWFdtJtSaxcDzETFoF6yaI+Ow+NKo7hQh
wRfgjnbG9hQn1lbT+/yGEVTJ1Y7g2Mh1OJ3osm9u32zhFL1INn5XU/mBt9oUT8N+
lDIOv1gAist4HKVUDthgGl3xdOXi8OTeVobTkVWmDdX0UX6HVhdamDjSebySbU08
hCxKFcuzx4BZfxiXCaaW7SIa23UWgrnlnN795rZPi14Ov9Boaq6Y0blx4NNyqmcu
N+cFIdvSGIECcRsaRPwpstM/J09L33d7v2BptTW0rZyCWYjambU5LS7+9/Pp3l7k
R+XJvrzbBVI0qJ+zhp6Nlt+Jvcu2i2smfl0L4xBc+a8VblwT7qW6LG7tLE3SXVpy
O7knrswRMJwMlZaC0VCh6Lfx+9NMAiJrkY6DT8qmismRY7PjfOCgxeXgtbJYh6Tb
dFiWOJA6KW+I/KX1QEA99a78Avn3mS62XGlbc5dyZsFFqhCjkqZpMWaQsg3yLyTC
xszR2ySJdJItwhNvokI05aLMujMEGlBAhx2DElsEeV9UzH2udebvkPbhA8t8gImv
6s2jSwCGDK2PSFaufkIwBgIP5u9Aa91a7FZAKUpPgF9h7elmxAc9sloqPHGkm2rC
Cyq3iSZE4d8H023BHftMjVph469NuLc18aT/UJ+RzpFOdIvSP/Acd33si+N9bkox
UWrI5TZnTPsOH9h24EfeuyO+AoC1PEi4Uk4TvOv6oM/mhsUMULr93EIXek4vCqtt
fXuUl1/WksIUFxcsWCazN/h+huFvXIDObHWw5TI/kswBmYJsAFaV8KG1q9qkzUvM
OxaQQczRPTIFgg2Qu7AEOJ2Ar39zyt8c3VATz1Sjq53j9LuASVKJuW4Ecr0zlvZ4
FEuCInGDkxehOz+txw78pA9QNMPkQswQKQYWj9nveP30/0sS6H3SkmSLO20uwvEa
tkEPMZNWe5g67SltTNCjuC30Tru/HhgoCn1Of2+fph3PyKQ4339CiRdhhob2PFEv
xFNH1oAJ/d8HP5mBSBl5cmLgUdko1lRzvad/Ts3XYW4CJcjwGXz1tjR3jD2igfBW
nWD21SbHDXBpF6N0RiClxXTpHmKP7AhDPkf92Vm9J8mYkhvQxANXYw5um0w7nsUM
qiIEika6JCCg39QIfWS/+SD8stdgdDr7VZOOOuXaoJCSpoNsd8riLhvXf3JpGyl7
Wf3H3AX1nQqzZgm4NknVMlDkhaj6GuAuXG7EL7TovqGvtkyE2sv+W0s4FrkZMsNz
ZzniW6PAdRCZi7eUt1xMbumbw3mmNHk3ggrERP2juLgVJDmTm+GnLVyIoqE/bhXo
WYkbyWNVN78hWf3BuMe8f4gI/ILLmuLoJCzVYopYtRSBvRF73aK6kBpo9/dfCFAQ
YLEtxsa+1TdjHIUNqhcmw3Mf59syYeVxpcYKdnmERuvz+IIaTgUcO+5CG30MZYMe
3Qcu33pYRFKqZRHzu/Hd+zPSbPjtbNj2/xhJQduvLSe2ri5XNPlsdbmbHSgI3S7a
ZEdL9mhuAeYU6nZ3euLQqOs/mbtZ+vOV8ACt8jxTqofQVCwpl6gODuSB1BNUF4NU
Fk7Yz/2pFOA9iG+ItGLekaKuYrCkSN5b1wI2Sg5TNkAFIlw1glPwdHcNT5EU0izp
pLt8LP0Cxb0JjE4wnp6qGXIMIRpuQIqKE73/vJUrSvXyCS6nxKovMoUpb5Rp51VU
JzE2xY0tXIxqXBl64wLm4GTmOh+hYkUY18y/yJuJ9GjkDCYVp1BxguZtp3yIao0y
a4CcH0JXa7OYV41x0vMo1fbL+GXtAJctPSLe8Yh/YPgZE57Tprj9/yEPYwjSDwK/
dBCgzJVa9GBVPVbynNAJbV3chMCgmMBpnVEQkt4sOkXXmOBtNdJTs5JF/nectASU
kBcPz8/rxDzaZ+/COr9GSHfjoNDT82du/qBxtKA99WBChUgnGmbv1LcwX4NbEbZv
5cP9KcFzJ/dNXPsaTBSapTd9zO2bKQ2JSdrdsvJyCcXI+JOJ6VspQuFGJ1Pa23OY
3+6xkOzvq3EKACFU0KPmld/DmGnXn8O/UkyLlm1NE4p1m8IgBwuAt+mzmiLqY3JL
SJRKDPqJHHKUL3U+2to8I9WQlRQZq98dVP4JsxjL/z2h1MjK01CNuuYCs20fwJ98
NJbY7OJzRzS6X+jcvKUO2Bml+u32Ya2iY9CyTajMp/k4mbKm4efN9w21V//fk9KL
P9ToqMQ30HwLrpIf3upReuBAqh920X9bzmthU5bFz3eoCM+ZtVPC9q9wbJqmiSLz
dvyErUxo+5BQrUmu9pUbKASNytMvzWQHi6lAzBL7gWo31Wg01RGxRZ6WQlEM9K1B
0OA6w+rdvYElHZeXl8INLo9cFDRnSGbT2+yOu6Zv8LPtLBd91me3yunC2KiqzgLI
s+yOaolBWyRcH2TCAiDeK5KMlEKeVvi/so47nT3kF0UQK6/VvOaFSam1MJ62S1yF
SWaUn29BKd3NTCQ3mlMVx94tS2eG2iuxHiAbDvuP3dE6MIOFi3QnDrswb+BW39ps
wHK0EOljWnf0Dj6laquxhprHSIWjK8pIYjuQncZBu2pHbhML7+wQaWmUclNAb0uV
XO/VWksfNWoG923NeWFEYleB8VLovMHzEa6fNzSZnWN2YgJdLSOIlzEml6bZiJEU
TRK6YMKMFAuJa49NjlJE3MMMisncR/iWe1/kXZL99/wspPqz2qMgDANLX576gOys
GXvXAh2llD4cP5DPlaHKBurTYSuTV6siLjBqtNxDwqbuSRsq1UBJiVJPclmv80K4
ylXUn1g0NfTl8nq4kkN5rBDAJUbxMIYD/cmJSZSTq6EhhdvlREJ75TninE/2GpWq
NmMGrC2Kc4RL1Klsw/3WQ4dnShKGg5JYOc/wUKPF2rhtTWPztUZOceQgWiSN00ZP
GDGgOXRoj3yij8tPqftJwqWtblJyv/DOHTkxb/ixm2j93lUGyuLSwY0qIR2OJWDA
UkTX293O3ZBdkcb6IsloDg23Kfl7be8pTFwNU6tOYh8/pXa8r9l3zBnlxkeUJDFS
fp3sqXpAZcc0zxDuGCY9rJ/COJNRscnJnj5PBpDh120vcXau7UwKdkexDzqKnas6
ZETCEXmkFrugQtxh6+LC8n1Oe2IOQjjOdmm3WNYB3OryeOskLCzT7zhhEgtFfXMH
vNqA54uT5dWU3zKr+Q2/GKjFgleTuiHnxfXTXy6Yn5ieAVTsLL6d1I47yzf7t+M0
L1w+IFxLwKjy4+0aiQOikHEGG/6iPyYaRZJnFjQOnSttXPmNTdEpjeM8ieu0m9Vk
les7I/dN4Y+SRgO3O7YR7SOVAyA0Im0MNEYEGJAaxOTN3F7ow+sS47eGFsNO1zwT
2KVLGqCW851v2GMapZcU6i//sCxMA6DKuV+hBw3bYavmqGZKNsQmYwuz16hzOpF0
W7zTOBc5oc+nmaDTOHeaza/iMdbl2sK/2Fh4KzPb8eIHZ0onrtLhD+Hm/i+GaC1K
Dca9zZKq/bZqmUmuiZWOAwXT3NfeZV/kCCpN1Qq+0D0aLcOniDEPzGHnUIGx9eQ/
eeMm3T/VikTYqmzO464a11iX+Z3qHa9kmR7ZqldUBPuafswWAc6eRPrCQA4leqQC
WnxU6fTu8zopkt+X40O1mj/mL10/g7KVdn5Njps6KkFkmpVd6CkbyfjfJ0dCFQhc
3iZggIFzwqbT9FBDQkT8ZAuGywilCG/epxHM09MXOcOVVHrccjtXYzQCh8eRISm+
cauua72JN8NmV6Z22uEKPlk/sWAEAioAIzhdn2nxaQNaE+kpuhCdQsZt2p+rOBV1
lsSHL/W3ueBggLRB+Ax28QJZQHTeMlOIA1IqQxjiYjAkhW1FEZmbLFmfBETW8r63
pC1tAM6SE/24XxzsecC6/n/2XpDIKyVnnnjhGYt1QCAODXIPYRjB05SUxU3M8Tm5
pswSzjPZ5VcMr0cCJItmS28rI01dpWf97tng/zBXO39AhoylQg+31yZQ536p97Bo
QV5naUaboNgs8G59ilMeTlufm+OGE+NnZtF/8uiqkrX90D6HlQWi/mAwZWvcu47f
pCgNHHJGLiR8glqCRj8FxqUedhZRVQvZI9ehCrhr5/H4HtkdQ3Ngpd3L09zp8WCP
Q3OZrVbCfeP4VvMZpm1O/Vlr9gr4VHLia557UqKRxzJdH0q2/T1E2ShunwFQjeKV
4M7twL1KK1ZcKYSZwiEbcE7a1vsRlG6uTUr+uE4MxeXf/w9BIyKVGVnb6620Ssyq
vXkp3D9ipze/GhTMKI/S3j/P8UIR/yWQiqMTSXjr7sZtGDu8nCCviJv+iya7wI9M
Fgc9O4ILGVx83B9gG/gFItrStiCulg7nHJcCNMmK4jjj+0J4o9U9KDopZQ0J4oOs
iuI+SJgMOCvPqYoqwAfMrv/uWvscVWVv1kImkhBIZKdhRWoDl+c0NY1GjCuE1Z9/
tSEZ8sczaMMyPeje7evpMKeqosnvBD3LeILnpM5ojOuVdvdM8wGcgRWqyyaDKB/5
wbs/EC7KiFl+VA89yLzZOPVgOPNpRejnI5JSuM8Qb1wUxCtWmAbLgmur5Rikb2x0
Wac+IAsXP3reO+cy4l7U4uOs8Dh3Sm30I3TWdi3gU9yRChI1s8DOVf/9IiBDLeFq
gjTvkfCMzu83yPoz8l4Xwy8yIFlmfMSz4ngwhzJ6gKfdxxBvZqAndt+ycEdE+g80
rTL/Lfg6qvQ5vN08/7wi5ubY2jn5IgXUJPa+cZ6F7A/r7wCF2mdRvaT1t5M9ulJi
6l8dipecShuhtIO5cRtEXXxA9EyKW5bWgGzAkoeT5MpJURqGh8CwwijyBJr+iNHH
PIictnw4X/btgamc/sUdC3FahUP8SMKDuNOG7/ZXdxyJJ0RGxenIRB9hZIMAP3qP
KorlFg3olP2ONGVA9RuiRmywwCDm24OGuxhwisdGFXxWKyVGe+MLigmpatCyJQ8h
Wiy4WdM9dkOv9NB7p4spBn7fiQcU2c3qdGvkQI/pWUuSXMnKuZ4bKQPvH3XjOqqQ
0SkCUBsz/PUcogRd6p7bdo52/rJW6XIQ95f67qw/AVjQBkuByO4h4MKR7tQ875+C
D34GP7tEgjSpt11zk7EQmJnq9ur999tPrJoDFZlzUzoAr0sB+I15gkom0a0bJbAY
iCqUro3PRMh3MRXYPk3kXPvjaOoYDARE7pv7rY8uUSmO5K65I+DAqj/GHhwauREn
J0EoZQ9IxQe3pW9YKRg6tDyDalAwnK/HxysRTZJAjHWfk8TG+WGSL77XEKj0uIPZ
mgfK6aJFkZUM+dvuUVx+j0Qut7FnLTtpxOqIna5Jn4Co6kjGC6ABCGwY/MM2F5ZO
NFlwl2NSfhjhtry7yHAMMCeyrKZStUYmUu0WEgbrL2utIJtd2odr2khCsYH2edkS
jBRlvCItqDK4kc1zZA9pHg/swe5lRXXcmfBEb+WvQf7zgxUq2fqutUAj4YcXCJwV
4BLljUG251WN+DJpvgmI7fjj84gjPf3yypFXWJ/i/ic2URYvikQ97Fr59QW9wizZ
SMsXlb9lMami5qvFriC4JwvMDfeS63F1IPiQgY0ylvN504RC7nOjh4Fz931EqgcC
z6QkjxITj53law7e/Lh6r+PINxkGUnz4NyrJZt+TDFJBPBZZ4mRe7i36fbw5X3T6
AXDNbN/wgZNwQpzATiMopBfw5/9TcivIZ4v/ST1Yg2OrLyJD0BgfyAW4826b7PiN
UTZfYnmV/FnreKwfHw8tiq99zhu9we9P1PImZ/oV+cEjcXbn3zwv0Os8MGGzMdhf
eHPR18LNEs1xrAjiD/j/p3eMtTxmS/kQIM/4JfJv9G0j8wRwGanO6FKI9st3x3L4
VoX53uSXBNKVKRrYK6wCVseMA3UpVUWG4bZAvTqHbU45ROhv5+UX+zn/+n6Tk9jy
JHYzV+vShN3d8ShrFMlBK3rDncO3KxL1v23Gzf2HQbmqJF1sIMOkPh3Kh0D92iOI
aOP0NdFFffwgZ9bKZpv7WBM9qHq/KSpN/WisE+khOO7HALGvgbIj10Uge5CEK1FU
U9K8mgXk0rlHvFRMbupbc2eOfZjM1fHJdfAmWtbfQeXjxtU8w3Ex/tpCBlaQ9+hT
pAKA5StE0k5VE2e7IvO9CFKiwoWv7aqEqTtixuNXff1Q1zr4Q3jP3JR9JOOGHK1C
GWFI9FYBmp3eZV+Y6OFyADOzbNAn2bhL54blJ8kqVjXI+OEyh4NRt9yZ2HTGuPz5
R9HdaXW5zULDbBT1/dWeIt4H8vpgDPz02qqHkzxSrkGPkG3SNJp4Vp/2rbtnbgBx
FkAPPWyj2xwdICB5R1wrvZIGNgEL6Dj5L/s9U25bixOj8N2dZdwRCM1FodxdwNYj
fWc5yvG5bzIC0XkRvytDmVdgSKR0NCoEFo48HIZSiprcy1Bx70VP9eDkH7NbQKC9
FyvvTf5tL9NRVmXXPB9/ZjPURQuwohHPxmDP0HB8laN3ilWuoHjd/HKEsY4rvNma
8Fi2d9n8Dilw08yEzdTqrICryzc/YAcFPZShhTzIHBqy95XN1+7+ajNUH+wUKtOS
DNSQFj+qOJnoOMS8WxoCNvEgEwtnuS+dkN48PRlwD9kTeZ8OFjbNUDZ1Fr1edqqr
dBuVmrdnA/tNoNJxtjZebukJdJ4j2cWud81Q2H7E9VQ6/7JqkPdvoY+R4lm9SxQq
JcdbyrsbMf6fQQHyoE/MdruOnQIXCniAqoSFAXpP/OIodPj0rpzDR0e/hPup1o+P
r/DGNGnv0/Xws1LD+FfKxUuyRJSBWxa/aeN87+OoOUKad3l6hW8xb58QSv+3YBp5
WSZuc7fLeq0IVBnOwU88DSivVJQ7pJiI3ODCUnAU+33Iip5/UKCFVg8lLoQ5iVMu
iaGqA0K4arOcpIzWoV8F3EPhO1j6yMcAYas6lEOW/GjX6c+ZG73pi5q1U5gtptnf
7e2IX+tLfytjjzNnvTBv4J8qXDxaVdPF/jK3Q1PG35LaV4p+kAQnLCQaQpKV6e5E
BP7eMLNqp3zqXQexRrm5VOsQW7OipHGAwYz3fIO0GPcDB52pxh/ykVOyvh58hfDN
LhLYzjJP07n3SvUhBHRbwpD2QNOqYVahOPot8Fsp3LKeIAuCiCnDybDAs25YdWlT
GhdSBNdW5XwK4ZiNiqUkdP0w5ZUpZV0gcNQd7AetMDEALTj887GLtSPEMMSLhjUG
28HlWohZdZ1O66Gu3/q+3ZYQt3Toq+OMSrvXpXTwJFQzSfLr+Ws8Lziy4RsB0Yvx
9xCQu/EKNJd1NddstrGL3Un0yFsusHa11R3MiTTSWkfxbXpJgPt8ni1sk3VBegPS
F3/q3nj2IxjAUttNlBtMV0O02vxYNK0R8gCbOT/gRmaBVMC8NBz5JNFZs+XtcwOv
CzviFCrwnw/PS9UdSQMBlBrbacR7gGpPVySmID5XlyAFB6L6oHyXKQcgLwa7YKQw
Trb7JsxsVA0IYsKAF8nGlHdeVAo22uOTEt429e3+lKy4rcVgv621vK9NOlMgA4Ue
MHMXXWXxhbSatpCqK/xZ8t8/g553JLzk8uAmH5lZs9Odhmw6if7A7ho+8Bo5w+GK
Cw3HeJ6vMXs8rTcTc5eDVLe1Qi2ZPRKDaEK6MAXfFkhZyznvOA/9UuEc41yapn2B
gvQfC+eygLpbgpMZRcV19V3pTY+U5WY4dCrS/nCBB4jlUfgGIHp/G128Zp9LN8d8
d8zdxjcS1aVDfUYOxat9LPvwK18hebyO4RTZdgeRmzfWeUdWF2JiusoEZPGQmjjB
m5Rc31s8G7rsfButcI2gCG0saK+SgLwndyhEAq3Z2GBdIcynJMtLIko45gIzcZa8
HGLPeKX5sDvKWFgIOdLgO2WMUwMiS+Ca87xsdEuF5az5FUy3xTqEr3tedPp81yP5
JNc345RqJvbj7ZohrMko8jDCS5FtdUdm0w5jm7GvJRbDLUnkTNmw7GKtBxqLrxy6
06JWL8fFvtBvOVV12K0ZFbbH1KaqJBhA4pnkJH0O2DkXViHLsrwLjrKDlUt5g6cf
YcREr3/GmxzHKP9E3WKUeXuaBvMK5oXGyglrlvt8IPebmHR9xdqH8iAZ8OIX9xcX
Ft2eTz+v8eMJ4ZwZL4XQO2IHsbNSQDzPiivYLeZjuaYOMH2lC+dWL170wfbNvszl
cRnSdpRfDWW3yWWoYFsprzww7wv4j5XVirfxwv4NodpbgZrBpfPHafNGkI9nrhMe
WhPwxjv7WdnrkrMsU5vIsMoLKnMiqbfz/mALLslRThaAc+sBt+cr07vrW+jnRtHo
tb5Y2vMYN4rnuaJmKGYvwBIP60VW/HjitbQqskK6jwhEdL61w+eNd0T4r9n9RYEz
iRLTxN+oZJgjw6j8FBFX5VAiqTPp5V69YteaXlMTvrB5OGiJVmxW2eGlvWOYLMyz
q9ZXybfXRs71jQS62seRmDrP73bKW0Z5P4gzcv7Rgo15s1J40ijH29BaOETcvAdX
I2rCpa0iwHb8UI2jMEsRZDq3VVUuIYUlJQHA9nIk14qb6/9v6eXYW/ZOWd5STZ2v
0Fpid6T3NKlrqY/eSGYdP8J05o/Lm77LW+Jn+ldxj22G8Ebf6UOTTgpPrpsFUsFv
cG88VqlSJ6ZNaiFhqggdbf3k8VR/h3T1P4uJ0MawfnE8nLgKmJmcNU1TcDxiuH0b
L4knJkjTM/FjmmW/WawTw+nRRNw3FAaCG/mgVflWxj24xoTm25VXcPEu4pqzbCqn
5Iin15r6tMwR+jLdXofTuHvDEhqJ2/ombMBGJZ49/TgVnzvi/8jS9t4jQ0GxNZbO
0ljOjak1gdxD6Sez8fD7m4PG/WtjOvv9C8RyKdrQuMBz9UeZXuXKlbingXqHntYI
OuFv2PVr51YmNIdhf5HKSSgXrXKYRqfKF37Xx5nD8XqshhBWtDg1rhG02CxZFu+T
5rS7lFj789/JopljLhuyamio2/e+BTh9n+7ULRkArl6EXDDF43LYT0Lldl9YUC+w
/oszxQijujVYeOTpyyLkH/Q9yyA95N+1ur1RdL4sK2JkszM8M0CkCOUYcVJJMsrt
pcEZUsnX7N2PfguBqW3IUKwpqYDfIRXlcDHvI7AS0VrJaVcmRhoEZUmro7lQJe/y
OKe/jmKX05cM/C0/QAMLJNuSpqR6GObY3Q1ocZ54tgR2CLysEDQwL9ZpWjb8hqJs
CMapnZd1Rue5shpK6OMR0R3a7hoAgfiTLi27867fUVS8NBQvth3Du3h3Ouiiutbp
W8lIRELbn8YWRqRdz3XTYuRwFLSIUDXLJB4wlfHnP1KkRqh1Aze15FgOCYSjkqPl
w8/BPeVTsUfQc8XuJl312peE5YJ6wUWIpOaAN/uoHZZtNrP/yh9vwqJheSPtMXV7
R1kTxHLzOjXRA818Yolb2PUAEv2LqBPZFlkkeVDVJMnKIHgoZzr3ZMMNjDwkGx/d
Pbmi82lzTLhIbTm3MXhbu537CkMGGmLmPG1N81slsG5aoOT9d3/KG2yZQQDJ1d3r
jx2xYQeXT3XTr8i8ztCHeDvqdWpKTh1Kz7iRLlrCjT1E+n9pIztP46NON1MV35Td
ttUuACO7wnOM7fsa9r8EY9DJgA02H/1rJg8pke0J3PUTMi02Y/Vfg6fRLkzZRCPs
SkL3aoTpGs5lpnHsOczJMRiPVEbi6ltDENjLGJfX382dKU456MdijJbaVxOLBF4t
PYiln3tc0mnwDmK6SwzoncPB98wBcisQOTwOgbeUCijjTtjTt/reiXEOAp8V1hlU
+wbYq9SaCdBeH4RxuS/j4nIhd4xdtI73H9hnm8H2griadbDU8VxQb07Q1LWaauKH
vlaVcyTc8ctomZTQ1kHpx9yb/ox9l1pIm22ODz9sUR5HyZBoSMrxl19ETpQMkgl8
lDPLdZ6W3R2CrQnc2Gp39aOfB+ZKxtk2BXxTAkbz4vGSLRrYhXJkiCLPpUXmiZ7E
AHPL7wJXrbGo/spddj6Gd/G6VC7y1pCgAL/u5Y9C/8CdiPelUhcmR8C3ZUhBaesZ
FkN63UW99XuYDmje3whc7k3pbDKtapzEz4G+o0EBoCyV6cnGXnVfvwHudgvzcnor
sye7Klqzwu0iE6QMW4hfi8E1p2SHfKfFY7cE6WSAwbXjpsSEGSO32J/rfcoqgjAy
cJdP85ieIIRx9JXXFvvsatfCmzIaFVs/hDl8dz7PsVuhKn+8eVKYS5T+MVxcBxeG
0h4sw0KmkIoqkgmgjI26UDXEhGpC4l7SwX8nmHHkYCc6WttsT0K0Ky2clt3JF4wb
iXo29MJYe9rN9czj1/zp1XH09W4smPQsEKwl42v/KYEnplAcVk8lpJNg8ejFbSZM
IGYERuUd/NvNIVaC8ZbCG6WvtJ/K8rzL78SW53ezaL3Q08PQR0h9qwfsxeSNR/tX
8x6IFyCIuIThYXDPHKKrL0WdoGEqN5ImxgzK4mVBiVnqkp4noha2VRY0TTPKLOSO
J8oyq5EM3OC0jcYSwWFwyIqMkv16W1OBH2NtEleoddSR45TUXOsKzbxeN0vAAXsH
NaFrM/Cay7wXGrLu+E5gmpvK5A6HB0qJRvmCoi1sSQKGhAED9xcAnz2VfILQVHnx
2IxGs6Cz1XpDYWCVURoAlbt6QwdZMxv1HqmqfFXq1zxp2Ht3oG6LdzQr1+vkWJhQ
2ReZOG431VQ9WdM9IJyw1+zt80hofiBDz0iZNppCaQnccz2n98G6MRQj90w6UZ3w
QujsL8XMpWJn1NhdEcUgz7grYZP2c3GnRRIBeZ0mRtMheLyGPkjFIX52zgkImj9F
llZacVWTnSKd+raUwOnV3iCro5MPlReG7y6rRJ9skWef50aHge8ESA9KTbrAWgnG
7umjC2LzpxpMTBKErQoT3oP8BXmhMTO/W0BRVZ00nwaZ89/AeWT4RAeXIGWgDKC3
sBxLkvI+vWjZpjp2hKumVrFjvT+ThHtNFrAHc4nnb6snfXuwQmdcbXzeKqrX6/va
Z+c3aR5etQY2uMoRA7/jEtPX9OiSERGZjgX7OzZCSJQ0XF6iemlGZw00LUdX5NCr
cv4EtdMlgZBR+kp0MwzxnBvdrsdgimhBE5KcQbgCufYMZuwcix8pCk/T9Zp1DgCH
XwI6eaHiDxsHQjgB8acLJ0NP7yDDWJf9jy83C5NxgmZcc+NrdfTZUKMAZr23jXme
L64pErwBcJkj7V/vapvwkJ/5wdyQBFm2R2oNzAiPz81MWU4D65qVU/N/A2bmKGvF
/hyPv2epL5AUNBtSZt9J5mkvxm5teU8IkRkpsoGV1tTMyKoT9YR6/bXlz65ZIi20
4b5HikERuvCnIaGjzqVdHLeVPaTrSPkm+pDtjRyf4f02ircG+PBWYURWkjc+mnrd
pr90AGmiDcKXhrw2QFxDtvzT7rnSpxRuak9p+ky05yCvWuGkgnjOBTevFlmIMzLO
CChHssh5l02APs0yZ0ukSM9aP1IGZi51CSzLBKS/tVm2Ekc4X1rH3xY2Uhu9Ttcp
f7Trzvt6Y7NHWZBRd262hj977aRHRwW6QfvXmRh+ZpgswtR48ld+YIVH8ey9XwXU
xmQVjZluHELtJ2jN0mDaFrc3W2+I+XJOMrkuMpBaVHrLMkxbFyAM6Q9fspoxrxRJ
yRm1PFEyoqs/0lYxJTYX4fghBOh7nsfI/xNbpvJ5p2FFY9WafU1TOmtyrIsdA9F6
+4nIIrC5DqQU7V1feq1m4J6dKByzDSiWoBfZoGCKPWw2CaMwybEmLYshzhCT/ipY
IH1pHmV9OqEdVBcwH+Xl+BFoHvTcnk3pacF4u2IAtKlTMfs+EY7SVDDpo+NYy2Co
WYdcw2FURtIWgBGe1bCe2pkqBhDx3zEDsdCwpbpPjHwVOG5PtUjHnq+7H9TRp53c
vTmeOoW3DiINjDI0DSo/oZ9TUl7CGrZjyJzR0Dz/PDP4q1IzO6D2rdYspMSnu/yj
WTNpRoGA5SO49oMVSdUsZUhMmho7FeS3Xj8HEzR47g9ds+xNNxvw+i+798nC4302
8rXMWJbjR12N5te0LLGS9IDl6QA2ZDnrYk53nkv1PG6ho9w2b7FySJLgj/QtXL5I
mwFaaD2B6gaSA4FxYkFI0LCwZPZl9/8Wn5TwbCri8jpgeOhr6dpO2tJ+yoyqktE6
WL4glpGmn9MFZCbfCdMbriL0NdQRGh+mfijyKoC/ppewcmW8R7HMncUsjdUunLjF
UhBGPdUp9mm7HpjmPNoA6dEbs8o6VKld9CNJyEMmaD9b+CGtOUmFbb9yL+yS0LuX
G3HY3f+jBkX1zg8+w7rWEmd1KhWeHNwoaYIBLODFd2aq2j0LtUIOprBHkZxlDS2H
1c/RTjCdUMhQjoLBOFMM/WGXDcCpXuUyQZf48w9NIzVgF8ToD3rbiQH1hjb6rpZ/
GpBJfJvLlwRO+D6Lj8uEmp0PvZ+aA0JYkMNJeOz0tM4R0jtjEf5K6AnQuNv7hdGC
k32tOdLDKc5O11e7Ee8tSfCCE/Eocoz6nCoZEHydXWtWJ+gYrg6sZ2ByzLHN9n9O
XIletS38FuEw9LyltyK9kB0AaeaVJ+np8OJOHX0lguuGrcdXP3UixKuooIqUJi4Q
exNJHVXlblqMzHBT3J87qqxF/qRxEK91jRJrIsr12JpyaUbz5vmTKw8/iJ04mpwx
AXL4PErzKiv3nELyGOTnJmVTlcCuURN2GSh0BZguaxRQ29Qsorypf84QTYgpacbV
MjxCUfQn3sr2CTNZCL0zATS3IKmSURwBjp+dMT/0l0r6j9yOdYUXvslDvAl2Y8Xi
bPDlpZ8oY7fwGaz1wv11b1EOZFy8EEf1Tzq9oVzetK21KyjnoKWhHqSOwYvoACdK
yhaAzLddGXmXLUYsQ+yhFjKxJ4yVRcfyT9eDPoBWJ8t6Rtdxy0vkpfOemXraDvvZ
x/moizyJUNCOetLPJU61kYAuRH+plSyhQ2GktXWUSVXfR6XYRPNQGo60SNhLOLct
ln0REj/xhKRPbkdhc98Iu7r6Kl5Der8WFj8wMaIRu8NlWBdNnrL7nE0IXWHnZvDR
tT0XHv3Uz/R6M7mYQTb4LDmkKz3l2qSw+R00G2hUUJLmkx2MVqfo3jDdWtckBisn
1+Qihus3TkyuFNENdgjZCMxgOhDyKvW6Oa0xmk0FgqxX0Na2naMM5oBCSX5/LzOt
xxDxbFfya8g5BpbDh0brvthWv6oGOQGasA42ubtaf6m1jPObI+i5U/UgsDHwLP0O
7DEUVDNwmJhrJe4KHuKz5KE57duPRaFGx/Rn6FA5nV2ev9sG9OhIgxvwP6u8npyD
j/t5Jtu+REapthQUA29NeMvUpzt5cqW0vhCw0yFdXdjtjt2Wwm8r7Dom28BixEQz
Yn3q3uVg24or205usYGVxZ0jX4Q26xShPi8SDOl6yJLPWMTSNF+qg1HbeNqiN+u4
3/X+9JRzF5OqFEzGHmpVPCqE20pQPA69BOfDLqN4E9riD3P1WBFQswjmiQY9Mm9m
FU1PhI5RV04O5hEQbWK6g77xOhfp224/nZtP5ecLTO3x9CRB+vCPanWgtXxQZmv8
VIt22WaSw9JUOpou7fmq06lXThsD3hrjUNVphvEG2hvMTSRXSFczNTDXk+FPA+O9
Q1jKG6JaGpi43yKdXM46r1f7tJODyFlBYu8lQ5s2/R8lEGhbCgwBnH4a/Mx+Bme0
HAjqmyao/nJeDB14aidz2SZNovdiyf7fJDiZtzdN4HqkkbbbGCNRgvC3m2TvBgRC
VdTFImySkmjPkysV5dwK7icPAnSm1aMSaYkKehcf0zYu3PoKIIi7RATgsV5Jhdr6
SOSQABZ7HC9k38rKf7DaLVIH4wBS1UPgDe/Rwv+qUe727Zax0tjjSvDK5YFMaAZm
y6xnTJ1+7wLbujR0xKnyhXMI8cLLQdi6MXufKEkn90vgeEVvb77lUbC7HgK+GO0I
vAe85ZrHKmmAWYIFSqCehMfbjyX5Y3l+VCrFCk7eW3ZX2WDf/0lMTpAlgt1BUDXK
Ex3VYINdHL/01lTFMANMX8NQMwlAcqHp8s9pfRE3xMEQNd1saxXrAympCbyqPMD0
fcJ9y7lngIj0q+71B6l0TzGwo42Xgn/tfbrncXSwZQMAMmMDw6wOcRl0m57u0N1o
0RnFGGPQF+D9xhex6u69BLLhQcwuD8df/HDZjLAQleBLwB243MLi8JpLbngLuJFk
gehk4r2dH2XIBKhh7Tb6WzKju6XdqLEpLZv1EThzDcS837cV25ftE8ChYHqfkP87
X4zvai7t+99esZxgYDqacTTbrEid5wdNNnMlZ+EpjKPWPObmeAM+QNhiE25GTkl7
CIK2Pa86lEYhhXsdpcW6IKcYPxwT+NCWy6hSET8ebpOa8u0b3q5QBI5azWDtZyHc
8QkVaDEXC0sadncagnqHjethmgmlKZDTthqSgPVyKf0yjXBOKxP4BZVSo0AYpoHW
VQKa/hyZYv0kYUB3kcpRcxyTdJeB8uJOM1YkHJbWMfVWRqndXPOc2HOoyA/SiUwZ
BFCD6wqU+O/ofcns7rvY5nNZURDv9Ya2N5Gz3Q6YlN9JojrmNr3SCIZpNL5CLnyz
v6Nj0TttfQ6nlx2JuFGUmArUTFzJF2VcFXYnbQ1M93osarEZPHHh+YKeGtXwmcEX
4rQDnhWYH80WF1KteiGUtQXy+2rhqjBZPeiwifcP9DKxq/bN9LM+JSsUkv0bKCgW
sAjuhImI9bAC630aGZP9onRpPwRJV8A9RsCWk5v2HLsmSk/c1ECQ4bTCyQxcd1U7
ePIJCpoCEMlskVqkpMU3MvsX0jPyWQ0VEadd+sb7uyhGn906ZlkS4Hxf7KmbpOya
4jSOOB/sT/Qe5ljI/p9/l5cv7vXric/sDSt3vpfnYhOwuG7hVydKeBsFcgGmwc32
CHMUPrr/YCLCy2r41lBwd+CwhVlBKWsol2EdX7YPSPsSMZq5MkOFoZzHoUGz/ESS
Pqwz+cE/gjdfatJoOkrnILdhYnvQYrlLOkdlQ/W+UKl8+ZGA6NYmdrKiVphFegPt
oU53aXZX+l5VfC5ACx1JdoRDEHOCNsgEQRchgsAT6idPzCgA3CWjVx2ygtncdD36
k1NY4fDdQrmLNOiINlzs63TD53BfZz1YvjaKAFZQvkUVLUt7iKCOa8oIOFi6A39s
MGRtMZGfLtUXBqIaA0UgtpWj2HTsC2Ch5oq3BhqTREi27I6NEv2Rjkr13rZtkPXS
q9d8uX9K/Ogj3QjSDS0LLb3lcV01IBTNeJJFry0bX+sURHWR0rYKTatiyVWdaXrK
L7+4/+l0yc58E1g8s4+qSAr6YRAJ8ijj55bt93jbYT78VZDWEpqD0jpSEuwheaFE
7eHr3ctm++3sBz6aFh+U9Qhj3nfWN9D4pXOX+0MDp7CcMXCse+oMd5xVeGsFD7BJ
pqo2zUKoHo0nf4BPnuwRTqOymrrQcbUg+XZWpKAhI3Yr0XfWYR5vgDil3m/mv9iA
xePllR85SuBH6xqy62dTW7eHvAdPjeudkvScdg5zYGjLfSKIZc5U4OiF1j08UxeM
Ky9uKiGV+kYFr78+CgiWah3IxYqDOAh7GYOuibXScFjLH2zH+76/gczOBps7a6SV
2jfZ4TcOUcacwmfBr5zcZjBKpCdZWUTE80uJ9ZPsqW7MV0tyoW+TDvlL1G/f+lay
rjjD8krYDMuukB/BTIv2J0zvKYmm9BBgeTCGaSAk9ExLdu4rpke5bnZZlhtASXdQ
8V+UcoKknI/ZfddgiY0lkIniFnYk+kucIcLs19ANS0FAfTA5Xfa74RdCglwv0DXi
/0xQWSbelD2Kq0PdupyESOpTO3KbL42knvRBveMycUnwIySuCTdOfO0FFue7xjqV
UIou3ATdBVtw7KqI1MqAHGOZegc+dTYfOt+aotFyOCkv2LeUliVzISnoCkqnQRZA
9ThDik/IA7nt2SCDVkIpFpk0LjjzYWfNFAhBJeNEAlt4VTd13j3qCsn077NRrz3H
6oSawqLcfe3CHeyphCDC7EXBGzJGpBgRVjsGCIflhdLQNtKLVpo6rMTW59mzasSM
bpW5s6gO488j4Tm0FDjqKM6BblvitI2/FkJiS6xYuKT20Qy7vq/oHgMTnBla9a8z
WpsJ/+fo29IV247OqnE5sXo1ZTt+m3gBwuB/R5GaJ8olw/gKP1hX0mo/duaCZ4Kg
GpZ0tK+M5fRLbbClLE8053MhCyb4sVWhnoLQBUDAL5XJQP/oX64o59DBcq/yHMdL
UoTDXfgGVSS/1rbbsvJY2zaeDlxOroYd6QVoWn+F0XB6SLSf7uDBXoL3vHtGsjKb
KYMsDdEYPFvU5AV8Z+zSuhvoKMuNocC0ZyJWptd4YDruIYu/m6uQQxaSHsxRTvIn
bRd8XFmlct0v1lrpHrNOxz4g/mU98pAfx/RNQXLAvp7PagZoR8wrCKdeIkW5Ecpz
izt94BMD5eAxZ0C7gO4y/UIlMojumhBQIyqPYeWba6vAaG2KJDnVGQfGFyn1FKRf
LW0bK/ZU9To77v83I42N9V6VmUwDTB1LOO/pFkJLw2mPytf1GRSwwK91IRLtAtr6
Q/CnpgCZHLYCo8ac4upB0dcMcixfEHKSHdtZgxS8GM1nGlJmGvC0GJvNnPM19KoU
hx1LGc7klJOKnp3+VHcLhqeaaWv0/erQUGEU61CzBt9pOqx150Zq8FTOqYNgrOvP
QdlPBrKHdfFGpGXzvkT3OutMlYdGcSi0+jg2biOatFT2mIHF06hlknEbT9a8PpJ5
WhsRimNWrYRIqF8ef8TjAv6lc8VwHnEneXh5brpRq2yLwdWjDCQDrC4GDAzwMNOy
6v9HQUZ2GlWaqOejaFXZMSwIZlJln3iuAy1nqSxtQrjmgTv1fbM/GVSmTImxuxXB
QvH5SctG3L3MVLJQIjuh0n1zA9F3KkQabioG28zNq/MVGqBFxdMYAMFHEJ8OgINX
iuR9OsoftrmiCv5H4xcRS2H+wVihg/WT5Yi1bQyxpVj7hyAwV9+88fviBqQad1j+
n27wBceUyXapXk+ZcqM9E+lThBGXGKwT4LNK9c6Wrh+lJNeWA+1qONBVuGdMirTZ
Ag39A0pC8yJsdPmC3EDvnsJuJ08wRBC+kDEn7y51rP+FC2RlZNpuagS20hTxTOZB
kE0sTaL+TFwBoHDaduLHXkgo+n/84jU8nYsnXIqBz5HWDK6+6z1lYX8AwWxDibiI
ygEM+Hp98LZjODdMETiO70q3k7sm/lK8YVEPX49RUb+3K1O7PIovP0ERbajzDZMt
qr0YBOB1sQ4wrR27YU2+S07AASEMXcTYtWhkZy0BpxfkzahnHVm8CxpuvSDWWDKZ
SSU/zNJ64fuxtu1oCsl88GOUge0uHLxEVs0HxoSGAEOTmMMHaZXQtFDFfgNEdIxB
p3LxDJew+GW38tZePEdfpHZdufaIWQzLefyY0yz0y4hFQdPQwAxoDioaONusCPhN
y3HtRcWW7iprcyWczwZRG72YxAButiCONuXLCsLbSZDqP0huK/Nrd+GKaE3gWlme
EVT6DmWGmvjV4D4BmtPnxrCUNfFRb4EQ6Bn7WrJ/Js2H4sr5onDgiwCDohtWjoEs
6WtXPxcfmO1ieCkOLOraoY7bOv6FPXgdmqxVoxlIIBcP+gv+pnkpcEAA5ZYIxH8V
Atr8b0yL4qwgPvpq+Q9DJMV6fMm02s9OqeLYZwkAKhIGXGjgfZ/PT9VhQlzkwWSa
t+XhTM8DaK1arWPwwbQi7V61d6wgDzqzvZ0DIOiaaXxwoj7XynXN6A+JSxF0WxMc
pGolIohlCP+8eYVCUl/UrBrDGvwvcTR8QW7cg41S3cvdZr5kzsW1ZM/cU/2yEsIu
WVwE1F3sJCaM1GZ8lD/lm9BSsnXZbFoJS4V+UxQEsSuO48TFFhKyu29rnc/3R0Rk
C865FL4y1WD34LCi+x4aMp2iIDMefTTGFQLYX0XAdX7RkDXppOcxUQNZqwWBQ8Bz
YUhdhV2P9z/rspRUBWkMMjRIMAyBuEaFwAiLi+5wpEUDfaDCWX8rzwNLo46TW9eY
1ZdPxyLbmyzj8PRUIjCcHtKr4ru5y3/pymOrhQHW/CnFMBv2QSFdTXEhpDHkWQKf
KlAXpsIZY5QrpIfuube6NSw78lsfZvHGtFqj7cSFamfXDGJr8nlHH/glCRwPYDvM
DEzDBcms1YC4QFCmzVd4ywl8+kgZJ/fBKRujPinVArrd4bLqm3Fi5RDnzW+cHcek
OiALwDQMlxSNphhmtPt9K5OZOQShwRrIrq4WXWZ3fcKxLmVTv6YjrGpSJGIvkFMn
nJi1AZHA7hDe10U50rYVf8FaGuxht4eU2bwzGNXqW6z/0JKJhReK2qjPrZ4clQDy
vQaVbmy84YBrSC+k8eu+J6KdvWP2EEtZ89UZEelxtglSALXfIpC/eVqAZhwDVJJj
JTUU9jZR46xmJWy1ojXsxXRtRnf6QIhDxq+TUXhuqG5WhMnSyJ8ArR8Wdd2IwATV
cB2aXQdLRhbNIGQZpetcyGy+eAHycILZg3xGFVkIXwVEpnEGNm3EVw9ku+8dzxUI
eiiztUwdGXRr7mPp1djqjeJ9x6I0GsS10Y/b2Xxdex1BDZdoeA5Rw4dR7af/4qAE
VAi7HiJsAL6V7mPjbPmqSWcnioNg+uex3uLJC+5xahhS/wA2HjMiE6Um7ZW8fgWu
6B1GL3XotORSkBgOMvIFV1WSVrFBX8VEBLAIQ+h+E1e0vyzP/qr6Jcr48VpUQ81U
aZFkYCOJZvyEs8nZUIz9egiBL/S6qAOw4RfV5qfQz+TTpSTKFu0+vlmf9WlWRs8z
Q1HO4gi871MHWN88FqJ7YLaLH8rWD1oIxkiXlf7qsxTL9GJ49rn8IMMxwHdMtM89
8KFoEVsmy1STZGdVMUVU5TNLvbvczostUBcyl/Dc1+lZc6xnEsimQo1CLX9dyK15
Z7PAngOSXQZu5UZRt6ff8rWOQESi1VbiH0ix/k4mHVOGjmlipLxfj34vxXB6tGdd
AdMM6zEaeIkILqLgmGV/9Q+VAOq72MNBdlOsyY7V/biJJKvfMfd26IZ3GJL5Cq/q
HEwHHlqWOVImY6dI53HzIv87B51fYTYllm0iJzGWw7U83YK02G27eygws80aadcX
6N5GvIM2CNPeqh80K5LDQ8b0oK9E9qd0/Bi8k6W/3xwQ2aSAKDyNbHE4bl5NryBz
nKahfXUHgNAtM6OdvreURSZqjfvtR1xp46rDOyaq3f4t9ST7ziZQIrfqjWaum5PG
HF0w1lZIP2AATkD1SSaMYgZNeajI7yUUDdKY9UMdMJxrq5HBIdgfi6aTEjghdzCV
7GBW8/DaHKQtYu2sveMsfViXMZGss5aI7zQiw76Onv48XnRltFwFKjs7KXEGvDau
gy8i2qWYZoET5tO8SgvBNlsEyton+buPPdSehLrSbmfGXZxD0dgAUi4AU8no0qb2
ihAMZZh3lI9WOPvKuQ/AGfm0LkeIKxA1/moQjknT5ac63NbhbofTH7EQ+tfKSnGN
LWoIW4sy/kjG+RnUiCK/QnxwTgasCCrzkltp4hB1ZCT8W2be7paR4VRtOuUBiCpK
nP2KS6KNIjLf11+bpz1DWtuVFZNFY0cFlOPuukWJi/plL6v9Iav0hbErCDFF+fZL
Fpiw/1ALzQfMQTgQs9GoiR/W8YFiQd0ZlPobtK8kny4OQCXom6WBcZj1ghjoeNoh
w4RW0eSkQNKvwHJIIsEf/Q1HCDOIh3plelXjYZX/y8IM99ass7lERWsnqCpTJ5Mf
gWXVzNVhYLlR/sWTISitaAie6dHhloz2gizeV/3JdAICA8zVue7zZqSQh/cxUM3y
u+YIcPNRSYGQoeoxmyw33iAnL5i69LCT5q/cMjrXgTf74tMmQlbYvRCYthMyiFbv
eh7JZAqO0qWAMatwqqFxRyFcy8/gZRAWHIqE0i1kkVTRK8S4fkaL6+mK9B/Pbpmc
zEjayTy6jj1O9F09/q3UCUo71KBL0uL9TEtjiFCZVbKuALdiudV0+t57Eo5LMR+i
kuLM0C5rEajGCt3XLdzIf+h4dpeL/DT9BEskbhzg9kp+EbnQZu/ZowtnqkQOhlGP
8L4KIc/8/JtSk1yHgSb6HTfs6rw3ULhie6JF8uCM2zLOVInDkaIn342uR0vKCN/P
rT4Ycoh1apGfeJQ9SZ6J5mgbuBviWjlskw8VBJg7dKaGDGKotTyS2bEanLlKKOin
bSFp6XSX66/wfs5u8wmKnMJ3GACo4SY487DYtOdFYjrZKl1cTT2bzvjKASZF26oV
bKabQnETzbnXLm9C0yoviMxU27ZhC+2evn3ZZ8KDcIYrzRHn1rvKl3iXhSst863U
4ReAcl3OfcFs/x/KRSaTg+sdS3+z4ha2KYo98LApOTJMUp7M132zu9n+OW3yDdRt
HO/K9t1l3fpSZAaGrydvkycshsxPcrp2leTdoA3tV/ywDXUjfrP0xWdhrTNYJHzR
G8vnngsNFCrv7+0idGLab1oOdjkNQWl2RT/moJhFvqLMa3vr80f4bRkQxjVJhaTJ
Yqg5pxSgglbj77j3nnWTYUnugON2UD6NFiSKtHGnoh04v4/pNNB7ItcO1nt4XFwg
3cYJ6pskfYazjgWwjoaUOtOs5sZCPzyOr0HYvGoptXdNDvyotR2/lJXa7MSv+jKe
NXESMbKM3FYe7Pxic+OGmxFQC/+cJyYjgkah3DeKjBCR7muUfMFmA0L5/pOg86Zy
+0q3/jSQWKDCH583nTd6fMHJmh5WjSL3VvhpinMn0KMonSuBIi1H99b6VEZbJEFx
9/D5TDYyR1t6FofbYkpbzUCsjbXCSz4WAPtFiJnsxnQWoIo00IIw0/DJ6ZXgYQaT
/aMPPWvMBP2m2gX1YIEdibbhdumXMZ8pI9fIntY6hGFefOGD28EZlXuV08uNp8SU
7tQh0DWRWea7lxjapyM6NSPfvHio/ZtpiFumjOVZZbU9RxtGAfLAo5URMFy075oH
XYcYW+A6k8dESnPkNJINQ3SsDFenrY9wexqOoEVFs+84KQt+prAcuy0ctYuW2KAp
c+lWvcUrN9LSHI6hZsV7nMOhHQEtgqb1r/WRaoxYCpLO+4AgCKZWVoBdHf0UoBsD
JnHWQnVSYQDgqZLgY2+gsNqKOh3jbkg2vKuKTdxjoACXtJJtDcwHpdCd1z79U6d+
hVCoBOygWDrYHH3M8o6JMMzmonWYfMsNmzWWJZr5Axln2+BO3sf9m3yYN9fXtfKd
1yIc9pfOOJsZclKSCEO3CrvH8rOhkRAMVArWtDMs2Uj10qdiHQFv/wAwR8GggaO8
2R0eLvg8SiI7NlKfHTrecqML/y4bHggf4dinzSuQvlN1T69o6QDkBRBosrb2KNgI
fSbYEZoJOTOgCWuE2WwrECq2ezjoBJM3/dt/pTP8rp41j6T/K3/Fiul/9bMjC8Ae
gY8TNsWtvEw4wbCAtvQyYK7Q7Dx33+0EjkL0E4gVbmiREOYqn+HFJP+FZjWLSvDM
z4Ys9Yw96mvswYX1Yn0fBa3pICY5ic1L2zHD9Z/ivsPAOEWza/FyCRQvspPtWEQk
nFdfAOhWfhtGbQJGu0LaSggDyOs+Oyd/uXqNi4z4qge7x3wF7H2uFJ+DuKcaTf9b
TPuy/Z4XFqjcS0J9JvHs8HcxEJKba+UYbfG7kQOozk4D80qRL0FLwfdVCm6kDh0D
xtcnDgQZcHJrNYYRsqIDAKsnHuaC8M7pU10xSpwuvn9WHwyexdo9LcU/FIsrCRhn
eNp/6oLfkDZrKNNrMJwcyd2aWqfV+RgkXCXBACBO5UsfXHWqFVGoCPblt1EJJLG4
KDsI8fCgjOkvIAMXchhUtBKDFYGFH5uhq9Jvnl3IUZRCTHvb/zZO24/iBBafYdiw
wifgEnU4v5ByXEn17J7dmRNOg1bk1yFE5/QDPLVJ0eGr69PVK+rgveRUZmnxpG8c
jraVrQkpj27AkrrLfYibQt1Rjcr/SzTCB3clDwfm/5huF9A5wYrt6DktzOFr4s6k
xQ0AMpUtlZQjuncAphJqbjwZJlSJdf1dIf+m70Al/LwtOIeM9GdfiRANEIvZt8zd
Is2KgunETAtbADRBP85LCrkiZf1I+dvSp+4+KY5IOxuhf01A+wCxjwJxGumbtj2l
tzask3noyt88QmdmHmzKDriyVYEnZVtLBWF+P/esp8GRi5bOTymoAPUI0ZCFqi80
UOZbH4VnmEBpV84DQLC6bhBiMvWHzJZA5VHkA2qjz+LHzQQKVCG8tbET0H0QJQqc
zH+G27a40uIZngh7UELh2f7XB42m3f6NQY1GfcCYo1AfKNol5lrYS/KEQ1Ph2mqI
/0+gn5wbOccfhXvpNhgl//JdO2ZhtQyu4kEJ2wXDrMoAAK0G85Cr7CnAnsEyxxGr
UmiFTXnCZkrRct2GTgCWtpG6DIKqV7z3Hq9bZoxOprk21sK0u8gUpy2oNJlROfUa
IrkFpi65TOJn+KqLNRxGU+LTfE0pQexa6P03M8P1wm5IDWF5qH8IVt131gOJdof+
IWLEAZCSEmMFdTiOA5YptsLuZwI4PX5L4WiLAePjYN3ExLcfeTbYNCSqmOE5qjKJ
VqaF0nAgI1MwatF8KYCRoVuWCczPKzUAcDaGDmVx2ZwEN+DPBhbxb8uFla15rplv
7jttIBc00igG9WLHifblj44eSHuzToKv749PFtkiBspwLpn1dNik04dMAKJUxRXo
pD0CJmJTWMQ7B6oNroWUP+hueqHTtCOvCDYiaKOmKH8Hsy5DjfaGnJxRrvav/qvw
YSnuCiRByyeDWSOvfzsj64PCWh0uCSVLniByVJe3KBZCAQCKNjmDlSrIXZlJZGOq
WJ+XIxtOMovwiJ9wuLG5b+lru7oBuxbfkNxw9FU0+3gez8zFFV+t3GnO+YrkFLku
QhkHIWrhZ4mtveUqvOxlB6gHnSX1q/oivlcDTf6NI6CSx54vsogqPrCfIKhjW2Ts
Fwj4yL68qxFzmVdTwDU2P8bT/tYS2xgY4gl7gwXhWG8NnJ9zRkvkbIzEiXmJyDll
j/0D94KteZ2VUOCEaqTS8Yb2RUrmUIz0Ymieb5y7c7WX+CMRr4RpGOVPvu/vRbEz
3OgoBcpOn5RQ7wNAH67IiggHWS51D0HIsnzRrbSUwe0BrXFm4zENE2qPm5gYNE4Q
QdfdLnz21PeqkNXsXRbYBjcjjOTeflUeWGENWldQKm/UXLR1wa/fqDg11Tn+YEFv
HHwYrg0kcIzU/3/GNiqx3jHvjpmsKHuGlN3FLwWseuoUcyjvTf8d+551g46bdyE3
6pXcwjElwtrgog8ExjjmVUBsN7QgzTTFchNBaevWjDwaINIj1Lhp8yeZ/tsMKOxJ
Yr610kC2XN6l6A4Z2ARjNiYOMQTT2X4CJQTXarU+74Pjy+HPOdQ5J2ssdMpKMm3x
G+z0tZDJPPsv73qpaauCkWWwHWwendE1ukzo+BlC/sE3IGwtVgiiWXgENBLwjrT7
QAjfdn8yktnxenYeWIHkUBKXRNTVw7LN00rCYJUjQpfetn71X7k9ZKWaPKm1wd3z
acTI8LPQE39wMY2ILEdJ7x587ny6hryBnvnmP9QddjLDiA8f593NvXGF2oEM0Jb5
0I0ZPCZQlmMYvr8/X+QaphF6kT4e++qlBsDL8eEkNDkQq6KesoFcLLtdAbpskpq0
mstl05QpdeGfOs51fLWoR+CliTUq0ObJzBsqwXn2PeqYR2qDk3mEFb4gKlzRooWY
xGnhIcpTMBlLkXn7ljHwBhWAl3TEAyjbr+tAiVYcXv8skKGyGQUBKxbTwe3eqcod
YUxRNjoMDZF0vbgZVts2SyDQtnXW5LNRLi9Y50bSnDU6wVjlpEIa57yfyBnShU9X
HhOXihHzJbrKY7LDLhzC1QSJmMdokF7OXkuU6xi4b9SCPnzkzyX7D57qkzlQZ/iq
3SgbiqUlnAZxOFRGlXrr/Nj+Cj+1o3GCsbC/8carC0f7+v8BRD3Dt6j2F1lhAIP0
rcUuCMO4GtTYn+MuaNDCkFvl1UVYZNod4ET8bF7upfboZnW+lZXAzgh2lpPasttE
OqXuYR6N+dikp7BMMsOdZUB9Dw7UMh+vNZL1IdrOGS3Zo6+efAg+ig+zE9hsiyXP
vTVbqpYDJptM8SmTu/quTQcoixZ761sReDanNhvm9R58ztQGRpk2WNDWe5eLmey3
rjufj5Y6TbHaZWzKG3894dzMSQZZ4a31pyC5LQ58XEPv61RPCZVIXpoAH9N+Fyvr
rjyqi5gxvAqLTBlQygey1w1AzdQKSMP1mNUZpJ2ba+DyeDDK2oNc7e85mYX5zXL/
mWpof1kNDAan8fVFnhBNw60/8F2/yXC0Er7jUzl/ai74uECbfxqwM3DOwS6xZwVl
0C+c+h8/ZFZxavyyArTI5ro19dR8dzGOWxLFv+8IXtzPjdFSrqxk9I1WdIzgKWqe
Iwk6Logj5c5JjT+u1EQ2rtTKEUsBgPTXnIpuIqu/ruoVXhA8zBBmhrtkDfA68PGd
IbTWYl7W+hTsA23SS9aZtjvWgNTNQZ2lfhtRQwu5mVO8SjrGOP+SiObnAWNE/x7v
gvfjHuNJyBTJS9L6bH7VkhJcCqdeK/9XCiHoDgdWPN9uS3K0BpO6vnkKKF1Aj73s
d3TnU7DgbJuXPj0U1G5U2xHCigfDJDdo14WeJ9KxKCSgNU7jS0i2pewBbLjUBvln
d5WJ19TdWW0BVZFHrNB6Pc8+ssuyjIXioaECu28nlRvvH6g3SWHpZ0dFKi2eWwv/
6C+7rKYKv0dL234cHPtIZgqQUlSltDlPfZFiYdTxdTRg3NKrJAQ1hEgv8pOkGpVF
BompqdLjHm7rC3a3LFZ75x02ejZFWzeksuDLOlpNmj3VOiZSyWWeA8/V6jAxXVeo
hGHiEE/HrXVB4NU8uA/MOOB7ervhVtypr8TshyE0GPXEBl9/d6kJZtsrxbJKX9Gm
UGf3h3wWnS7p7czyS2RykNbceIerv6oM4H9vAaan//BNw+V92z0We33USa8fi2oN
2/McQC4Zl0ibgvIXzhYeXKbagqeDVT0aBiSNxyKRsA0YoZSDs99kXv3VQ0rhyvfJ
shmn9kmgWS+fE8bslC0UPJPm1ahnJi133skzu9lE+oQp7qOU640zA63GRf0aPVo6
hOVWccZ/e1G9q5qqRkavkb8oZQZV794TV/ZRtVLCG2C3xgys2WhN+n8EA0M4D8p+
CWaDXTO1PTH76lqu3mt522zNNIDen0Wt9cYZM2MX1656xPgtqwYQYB/qI2jOaNkK
oxpBwZCATX1Pdhh55NEXWT0n+A0S94KFxDLq61leaUmI0ysGQwSjzoe2QEzhrJeE
rNUyhHh4REtce9KOOZnbBkx97LJhsy0SdLEX8mqxA8v0wT2PV9rxujmbSQSgcpJL
ynDd8hNrUdt2fGlgBWvxUzwIjvH48PNSgwg5HbQPrx/GoPR6PoIH/fxyxsR1g6Lh
g1IVSuw17TsHk7pUZHp3LOPJxEKC4kSwXmyC5Xplo7eneQfstpUB+733gBLksBzk
6XAAo2cP9Y575bdAguvQgc68xgDhiY3IRSeTrpEx+PZBqb6Qp2sByomY39tWByS0
uLVw6dKMH/iVdguboGr1kK8Kcu1GcfO2/nobF30J5SvYutR2jKulB57mImuXjI4K
h/cAhFOGbqvsbrq+whYzZ6KQU3BVqmHJlRTStNPhjDj5C7h+R+3vc7Yy5WSE6ev9
vUFflZuIhClpVAVdhfxFJjS+khBqTUUU2pdFZZEVnNC6v2xgo/cllaeO2YXB+TmN
UVZacQrCIKGKmHeVbBEGjGH4/N3i0gHKqruTXAJoLdwMSFUliHUxfuFKxyrX4pj/
6PnYE4Dd76FY67Iz4KHnvulZZFkoZ0iP8hohx0A16qsI2PgJWbhN0i7Jw7JM80O/
qOjrrYrFAjCZU2g+1xaazeU03FF+NTDt+7ukzFdlH3YB3dZb0eD4JjhU/irMhbhw
0P3iBCR5BZM3nN3WAYzo84f09IcXz9DY+f23N5YuA8E1BILYUm8gMTIww4JdvQr4
84tOaVWkeE6efkxW/MUeXr/5ajSs2wBEz8irGQWSW9CgUpsmZQcPUsMxI5dcEF3m
2UsIpf5iIssDpxMfmirWOLmLgdl0OEH+ErjnGKzCqu7F0Nt5f6PkL3TtSr8VwBwq
0DCi/ihroLh/OFDGO53Gbw095nqqCJxb8W3lx9N3dn0sporUd9/jarhfdX7RmzZW
cwQXYdj8fZwdr6zVDKrlv+ZegBTbui0l7wphfYWiUorXHsmH8Pa1y5zQbbpG50xA
F6SkMnCLl0NSPWTjw5+A6uGqxxx6nqOEcXXbT9ElpJHnP9hc+FrpW7as7stKT1GJ
Bt14182JsAigCIAmsLrz7JF9hmk1er8uNsj//B7u5/qJM4Omhq//SRaDsG7omGhi
x/W9/VQPTXXuatVBJSM918zUFFJytoiEh85xzLrLiK/z8cI6Pvjuu+oCVisq8lrB
xNcyv3cwLAUE1jc2RWOTnHExZjM+MjYdfufurkg8AVyWT52kkv3FDk0WbEoYJ9I1
hUm1suXOtSJMzJzfw1KizsekVmQJuVU1fxvEu7BPsoCea6AROG50Ayta3idbGtKC
s8ZZS8SGNvagJeHeOhSJyGG6uMiXqwaCy9Wjy/QrlbvsFjwvCgo8t7Px0bCbMfwe
bxcLEz//839PfjbEnEtx2bUOmtJX3wJMnAcdAmtIed1Nu9vcuvDWdroKZ7hzmyQp
yHHL0crB8SFYg3tMz6PKgLR1anspu2ORsVUJCGXbtbgIsMAJYVzXkbvjGPozFYYl
9GpCej1XN0hgyxHiyon8ZwfY6TiMVumhxzrd6QyHACqlU9gvXe9C5h1o5A12mpFu
nGkJdazdBRC8VR4tUT4vm3snZh3pMFY3qE/dPLnmEDXsOs5HnLlh2hkeSpbaOz8g
5nXwhSC9Ont+qmd1pytMJukqU1mRArE1Gdf8SucwlyQ3rvFqtYZlvsXN9225CgQ3
rXhTVrpz52q+syME0wAtJNB1WKBYS1Sx1xH1M5jqQXNmomQ5+tgUAOTVzOLOOjo9
pD55jT0jWYykl90rc4Ep2nPOjnR/sAquITMScngvnmvGrGCcsKS/8TsXnPcedlhp
ipskcOTTEvlEmZVUP6gJypLy+hNecgoPIBjfYnzG58bmSsmD0gzUDrkQ4dbMjGBq
H3jpwjfkLmUfYukqeEChc5Zrvv819JulEyirt1qbp03n1mKhlnIFZUFUwOPIBUCd
fiKqQOS5gyswJ5RvLN0EEBn2YloBVxDfRv/37KihFt0FLOtMnDRHfzIjmQlLyflo
K1kKCjXx23jMaFC3nElT9TDqqX9xFOGcSf46G318Mikz77K4UyO8Z/VoQRtMaH3A
9AT62YKQXH7ZdZ2bEVhDVuoMW2zP0eNYLIoTZEEQNDcrzis22zIIbYyNu2Bw+ZpY
ySmTMkBUylrXBy+hK3g1iEeynQtqrMGBC/M9G9WWblPRg2LTbzVUgpiTFLerdC8x
c5VC8Vb2okbFJQ2G7MJ6sAhfZOxEyjEyy8WZDehGUsomWQ/wm3opDm129dCL/Tyx
1i6bZpDtvqgCKVXUTB55j7JDMKYzDfsj8yFg1rLIDAcki7PjP7aQH6p/eusGvuD5
kqDFwIV417ScsmxSckt+zD8vy+LKXCeC+oFgl/DjKi+JbURRi6wHpjBcisJH6/to
MNd+yj4mGFMCND2gsUAiJaiyLAiCRQ6xX2Qwohg62D4AHoG7S+LdJXthTJfoPIjV
/KvzqMcWbsRXlHtwbu36vD6y1YH0eAGGNW86kElbN23jj5FhcpOZsrTJjMt3oFg6
fheIFIPBBpa8jrvpiNEc4a2oV+pNI1E2tnitUPe9SQxK9QqkTbH5pRYHkGKpipKr
KoJZRm2iO8n/ixy6iJszq8F5mQIx3p31r7jUKMFiZQDnk416zqSEdsGXzndwtPce
qxFGBAGhC0XarPGSfqci0cJTFylrzC1dk1vvJNxHR2MSHO2cxCIec+tqe7ZshG/p
6U8v3Kp6zsU8y7WwqKAZTPaMgf9ARtTL/uFdhkCIX7HYjooJAUdDWTvD0/sn/Vex
AM8rjtginTm0L2xvQuDEcI1DGQVYCtmOAg5F+lPn1btadI4ojG9XPVaIc4wKk26E
DKZiF2ZmT++RY14gUwmZSff+2vl4XwHGB/r+gWefHuBAbHeerOPex6PQxzNxQjlu
s2FYDr7u66lhcubUwDVQWohytxTAUPIdChRooJEzGTctvoSGlpzsO2AdZyrNTGOt
DAir527aCxM3tQdiRTrKIsvxF5P+2tCSFG5KJAtqwkivNnPjZdTbtmHagIDp4JEv
goF81gicARu73j2eqSuKI9Lg4jocz8txtpJnNZauKUEKi8F/NjoNar2V/NNWQ6RJ
GUH9/mwk8UZES8nsG1IA4snoGVxx2+6ex5pY4+5pHBxnjwV6DxxpsBhTVoQmqOyG
0JzAs6wKcHzhZ5Wz98Yydo8LkgtfpjK/7fR5nDMX5mPuVPBVf1VnnrlM5+FU9oV3
rhuOFx8kV3liamg2EVLZ/qi1hozjXEJiqAg+mrftW6GqD9BYLrDDMB/oYxAPK1ws
c2HBXR1RFQYgUdaOpTC1g9Qe7ACJCSwSqrNB49pDAhpC8W1mJGpeLEvpyKqZmyd4
rccOexgeW1fVWZHlUn6Z8FU9xSmDdLQZSSbXx7JWlWRC6/nJuJ7I73YGVpMY4x9h
oYzbpgLWc/kkYzP++ZfxFhPXovw6Rt1py636/jZ/DPEpqz/73gLwugd/BnLNqwtt
JxvS+BThecz4qIXmDRhvPpgBlewgglNDHA2YifuOJBtIeSy9nd3phI72rS3/oplq
6rPPw6NS63U+geYaXC30pqiKqNvc5jG6USd+v370C0l9DTszwG+KWZ2LfQU5Eipk
GnDzdgMQ9z9/22F6qodbiMKtJnK09za2iJvEP4AUI4QvcriQdBXWI6h09WwCNsd3
RSt8p6R6LxPIlheB/xqG//6oxv2unON9MTNT+VIhboydXvDgVVIKqu8Umz1ZUYdQ
yZ8zvkHxHjP+L57+CIMdA3SM6GAIU3C9mrBgDg+QtQAvCoaWLRQg1uiPvSXDBHr7
gthfHoTMELi/HzmKGrdBQPX4lDSUfyG5KUaR+s4k0Oi7Z3yoVVlVdQBwSrUjoe/4
vTi8Ay/p6VxwReRhn4zIH6yCeSnaQkMgGfIzVB3F1rMwR0OnOuWyI2cER8qs/wPe
b+OzxVJBXNuxz5F7r3DtZUMxAq7Pe9wWne0S5W2BvmPlRfnN71oQp26SQqbt8YFf
mJU+VycQC9kZzj5QX/ME05vzyd25P1szYZq+NxEjiCPQeyWoV+aaP10g8nLuwsAG
Ih1AXmAdxUKUy9cKqCO7+aDsMtaldvQbLpE0vptixZpjhh4Iab9Wr/uk94EVon+a
CVDNSn6EcbtlgAvnUa3dPabKPsFmIZEiXD0mKGCDwxkcXXWXm8Pn5lOdNkZD4mxZ
2tJxRrqwtRQ45i7QUKRZcxz8B4XUNkuVb9dibxGpYSogsDqpY/KnvjXRjKnZQlNi
CPCIparRtpy7WIfyG5srM10wKpxtbU0BZ5Q6RijzrhhWI6mSKAedWM9Es0Zdl0Gg
jPQyzaP8cZgxvT2n4zwpPnm+hdHsMkVScU8QyI0G48xQUVvv0o6bSILO0cuCthJ2
FiIdW7kXj/FPYxRNDJqM1r2G0+PPLoRMyUlaq96qS13TauUpgz2HcgqY6hC6blql
ySPB6RHEh78nQf8BxzP5t4fr0B0GLqkYYRm3/6lA8pmbdispU3/EZAfXW+dWAf6O
awxaIaPGsR7rC9911UlURU8PaC76+XVpVBdYGTNAaAQsW/nuTbElCtQ+Zo59ht4w
WG7QZZW1LDRmxDUOFBeuHV6V0IIRfUpDGf0nDWz/7/g2I62xZc9jU79eGHX/ZmU0
EVhUo1R6MnOXjtQ1a7hvkjtiGnJO5Cx1Qd5cHHiA+2DCOILrDxCrqTT3l9Kw4AEY
QmX/4RK72ob7VJ9BjpXkqucdRLrGEKjJTGsAxt3XEePkkqd91B82LF3c5mB287ZO
ExwpZjHaOFLIHnGmPDCdQvYHm41YXJN+BOHF06CueM1lbJ9z2KskyX/ieCyKFlnN
rDC4t33fqQKxKvSO4x7moDv2q6LO1ePddpmWKHASxLATTBhN5/7pDN/8uXyLm9tR
wJO2NznaLWWPGXENZ+GlQUUSMJ8DMPx2AU1TlJfTQurpfvmoWzkbQS7rjHKCUAPk
sCbLpQB7iXi7r5bXFfOAWVzmsqkQd8OADI27MaCnZOnGdXDDDNhBtBLpojXeLYSW
zWpskYiBnvVXIvR9zEuCjnBDlfIminBr0BpuWFi0JsLkl1dOGh4XoWTk4e3rxQYZ
bNDcEu9MKT6gUVrgujRngfWMjCegfA24Tdc6vGX1inTzSyPOHC2p48JGAzjb8iAG
WZs7u4w+aDyQJFVxdPAe2BfLL57choixRFWUgkRmrHgI5N2N/jA1XL6n9bmkH9hk
C9+vokbM0zM7dMcG6o1C9XEzQjCPR/nrghQ0GiHRvocqMcE7Qhg2ObJJU2MV0o+R
4Lw4VDzPWM30tMv2+HVlQp1rVSVoKFDSBYt9oEFGvH+C/eCy40gfxSvb42ZeKoZH
lOCTnl4WcxYcbxpbfNXR3zORdkIL34E2+kcLR6mGJ2s7UVX0uxyJaLL9iu/PvnI5
2fO3UHKFAzQXpLH9qX3orvIsnQ8a5C0eJF8/jq7FKzKE/krkFFpLvyCtV4LmVEpG
3/bBcHt59wY9QKpEuGDfHQJTc8SxTe/wdBeaS3bVdubkHLGx/2wX2N68vgaUXfeB
S4okMUX9sWfKBcZ1aZPiuBkRg+PtE7k2TAkK5Cbwlxbvwa2D9BVAIz9wPfYGlILq
9u8tGpqIGEtIV2HO6Y32VhN/5bSkbdgAFN1GXd39uuHd5WlnA+BU/i2o0eplR3cf
fIIvUIacZwM3lyYTF1EaagaJ/aKzXFxpDQakFJFEuCgLjkzxd7a0TMOcdiCuqnKD
WsAgSosk6mzdviKIQL+LIrwsKGACGcszPzku/Y7lBDFUi15nYV19Jh7BHjW+Cesw
FlvOcSnhuGqvNbZ+ZUBGPRnHSFE2o+h85xuLKgu+a7R9Igq8E4WSlQqs8EK1saJN
+7uhyM4LhGX1rrVXIicLZ6WU2ZH6V0J3EYINFsqsqedkyRClVxWzv2KWZpberWme
cQhpkEeRvbQ7cNxdpG0lWu/IHwMSubL120p/N28KVq1Y5S57LvSPydWwtEKdOlen
/ElKZHGMwMx6OaHcv+zq0iQ8I/vdyINagw6aTO+yyedHZs6lwfSuJxaeTwXeyPgc
TQS8SgGTwUNqIOABYFUYc1YSHh5GSDGSoK2J1vbigANRXUnCuRjkVDfDNVtCw0Zp
SOmElY5v3wOUp9yPOs2aijMCnJb1OsmL2+ghCghUmJQrHSopwq4FSe8ZczHPSRJZ
7UnBjTYyltdNCNgyGqmXQn08IeZIw0SkRAIxPDvJ4UR8tOVGQ0EKga3STtMkzG0o
9uGs+C+G+qWkBXYWTnr3drUlne8mhS5ZxwlPpierY0sfl6d3akvUX+yA+PlkLoOQ
QaBiVmTsjG2898O1l+3RlcEUStS6Xq2WqEzCGhGhjy4VmgzonUFI56MRwBdayl+d
TuT9pX2uSS7LLlkVu29EOnwaKg9KfaR62yK+/fqWvx4rd5PTu6Lq2z0FuVGlpkME
IBF7yqzhmFhFqAqOmtUpTXHbg8Slu1j292Iy2DZoGV80YBGeOo7AsjdRdHrKgdf0
hJx9TLzF4goskEFop0eIAV4IBh7YCUsm6t3QDE3Wlk3bOLDOq/TAP/XQKlFwIr+a
qdu0RCVDm340aadXtp8V7IcrqxHYtaTYZyLSfVBGw/EpeencPQm8dKTH2bEa2WXV
PvfFVWBK7JuCCKAf91rP1OBZbeIzgSa8QYz02BWqJnKOwOAM5rb6o8WhCWjaEh4E
vfiucs8vbxFWJ8HADyZgt9YsSo90clEco+M/XsNn6KcuWCv3gZFusWKM0NiRP40b
uC4N+j49h+X9IfaAxPjGWJuTGzlvraWSpFrNsO41+rwHkVIX5jxD4MEU2HsxV5GY
qzJiCT5V/NPf6sIsY3ktZbY4bVl0V0bqUUz79CKnFpHfupb/75ayczDMsQb+nFpW
Mgog1QhHBpKxm/twuB/p80nbV+TChltxW4SzvywdTXO630mgppGYkezg371f9k04
5KexfzIes2NlhiSlMJlN+jtkURF0J4CRVKzUjUFfR0okFBFc3NjorhPNAQD8wvWZ
zbvNCy3U43XCDcjyOw/3ndHdXOMUP3fYRrclwJK3XP3UwA6pHwMP7xtoAymbN8Vs
Nov4ez9J1d7OciALzkqW+YwWwHlZFQs//F5htruZ0UN8jyArZllGQyilKH8Cl3tM
CW/5kwib8hh+k4CUBOAe0EqC4yHQY5HB/zMiY3VK3pFpm3kaEc1xXVBkeZJCHdkI
Ntpb3uZR1vjrCXkuxtzidb1gvDoK/OTvYPKqyRJW/iuRnjAYu/HyeNVQmYQrI93L
EgpB5KeXs0Y3qOfdaR3MQL1h1s3p4PlQK3o+0RinEpdfwzUGUKnaaeFOZF8cTW04
sOg2FnBEdGFS/DX9N5guXkeVO2UkcAXmEFgVyf3bDVcSC0T4qyeMExTQe93PUMfO
WtbKAf1WDIUd8y6em29/ulU0q8gHMzKD0DlTu7MaoKLBe6+t22X2aANA1Mb0boSK
ts4NN1OLMq3+N//5wICyOpuWiLl0ocN5eB9BErqqeZvcqLiEw81ihonGurD6K1qX
prxA//efGYOxgj2zZ7JG/cGbPKcgYRyIQXqeidDCVrNRfTgyXoZmAxjeirrlJKVP
7lewuEqlrzucq1zL9AqhPVyTjRMN05A4T1f5Ia0CE4AtHvizBFPnuG+SwSFyiblN
xUhxYWWabB7CdrIl4RZGFYaMNZ2oTgKZgipYtr0IklycQEHiUxYPU4VkCpQPng4A
m8rJ4CHWZ4gg5PiDPfILAIuxJIwgrG+ZhCIxQCH8TKIxGIzTKbMJCKrGAhrgTOB7
7j/cjmayB1ET72GvOIOqEPqvNiALTBsod++UAMQSE2pPM6rLjX2c8S4+1Z21NeG0
06qV8zOHEIuz5Pa9ft6H9/hdYMkOo0AMX5QAs9cpNsaMc1alAs7ywIONrox66ygx
bh5xccWOp8w8Kse8MPsdG+KDZwR6nutIC5N78LBcVyc33yTPfvCh2Av6VCYVSApf
f/LIROj21KvYswE+b9SArcZ35Bi0HxvD8o75bKLlZSaGoRIckcRutX0Jhp82zHRM
N2Hse3N1sJACS3J+Jk/G8nLp2uL4yxY1ZFeuHfb81uyg4BYVu+iinBm98W/DlPxI
IIlHGgZF/XI/DkaEu+OYkpMDZcMlk5hLyXJF0sKYVgPDax4UIfRzNQ7uqDlHnENl
VZ44G3T3vWEaAm+7n3f5CrX2qlbXX2Zc5oTxxQ81z8Ngq6sqtVs5hKew3e6/pu9X
zSaCdovhAvfWRAMLgSbY98seTEOVFVCjgKZLgrxysywxcWwQGXC29p7YFCIyQegJ
EA3f7HgTg+bdU7X+f0PChuHcFvTK9W4FENolMDrOo1Hwnc8sjLlDEBNekGT3kaT7
+K+FA7VSeOcSzQEJcfVmawwqQNMjSZGrh5SixpEXjefhIBQGgAM9bmrfF+wjEctc
3NH6hagYs8VSujYKUzUQYtK3ikMsdBOR7mjdrS40nRm+8DpWl8WKUDgPNEADIfoj
Y6kGD+t8Mzy/OANflxco/OmR6cFtWDQjL51VfujLkoa5bJhBGgiGwOjKuGkMMuON
DYhUKOugbEgJLOuAwKiO+bEbxT/jkq6sTmFORMQVnWKoyZou71FlOJErhof/1Qcq
bLWi7P6O4dZ69ZJ34wBuJdaNrZNwSKTo8hmtUyVzI/PjrvNKxUiItSdhX+abkdGR
0jNUYb9NW0CA1LVTX8hMS0gp8kfzjs0LS3CQJ9AQjXLSi/bwX1cKFGHGc8Rk/S2A
+g2aqEPyF8ZIDkhUIfKaOH1eHUHi1JpRLHbJmO8c6Rue7qJZjRDWbwCcS4e4ut3J
t8L/TlMgqZ21EHARSyszsuxp+5onfYs5Y4XEpMHfkj9lK6StSjYBfQQKaAGxA53W
1TN+3lzeqwKFLPg1bNLQt1b0CcJ2R9PSpUwaB/vUXH2Tn0zhiSiMUptx3ipPPjgy
2Qv8pVpQeYRiRJbe849MXotL649Lv9E5pEOTRiyqRbnTQOAcN9CjlFkBmAyw6M/b
McSx+3n0FGZ5id111yNR6SiH62enYwGRc6yWMr8SPDkC/AaCx0OF8cPp9PZLrD/n
Ew66tplQ5jtMrZpoi4a45FIwciPj3dFAWlN5iRXG3ax3OBm67AGsaNO2ZXUHVcnV
r0VCeZl3Z+RDRfrugcrH9pTQ0lcYJHsJxExFDBnsXXJ37GU0vJUYT9s+3akhnoZJ
KoTQJxszbrYEqujXkCaOWUA03MV1Xuk29QWKKo7JLMrqmCFfdyuQHJwukeV5TaQt
PTOkzdjOuhbOqzQ+ehaKmyb2uiiVlUH1UaTRrPcjcaDsMMHonMw0QlZ8D15VdlcE
JwrRmOTLNVAR+o5+gp5Tf6uf4WYytnYJoWVbVuxjINjcaCC1EJFmTQuDU54drowp
ClwMMHADQRUaGRUHzftB9P2ZeGu/z4HoK9m29isiJ9RQOcq7cRxeEEujbVKirJ6R
DWu/S1i+OCIHEgSo49cEhMm0U/W1J3TPYauczdZDiGwWKv41M0qVmLHwE9QRbbqQ
K5uee5UTE15zl2EC8aA3dILfjgxKQTUt927XUhyTOlzd/QEuo1WkRVdH5dcsdRRG
2IYbs2C3ocNtWaGt+4YI0GZ7/B/BHxDOTtEkOuvbsitc4KIR316X8c0C+jIMppC5
+wsWPLY+6K3YR0eni7Jl87bVA7YPnd9oIv8ahVb+t1CBgMPl03+4rBV1vNjfi0XU
yvlMHINcDnOyxuupwffG1J8GPrX1n4/s8oVFQ/cSOhtrVlVAmLy51XyXBJJz4vSi
6sBBDb0U0rps27kfvxNqtsSEu7jLuTXXTi1h9Tm591icoor7KhLtggysvWKaFydP
Ub/1acgty/OFhISrtaGrK9WkUheKhKmcmtNQ5FMnTF7O44tXAP+xZ9DhDGIfjUH3
220ec4PNIzmxtdWQDCoak6FrvDbtyB5IyTIZPU54pCVqKmbGvGhxxoGHUej4hO/L
xre0BqejZtshSuAzxuvcS2Q1lza8DMG8pBhmVcvwtB5zr+tdANJReHSlvYLgjpm2
YuaK42quzVEutIQk7gUtdXMW4S44+qEukAWJVnP6cbdyPAJOdINXEXz8N8tMIcrq
Ms3CqmWyuFFuzlWbIFKoU1likWiCk0A7ClWwq86McpTVxDW/C9qLrbRa70lA/o/j
pfbFwvilubs/SzTv4/BQ9/dZwFre4yQGHzypDGIH58bd95pYUBXEpekgg69UXwwM
g02zKuI1TEqybCh9QvSgX+2WYgnt0qbz0aUOHOTxbNQzOY2nGDKX7mvzBDw+ZOX5
3jcae1omd28oZgvZXHXvvKynet18715LkNAGshaxZEBzKCyjpvipTro/3srE9NpA
Q84u7ILX1gpmoZkEM2I6Cb/YkJbYLhHCZSYjmAQsk3nKrJqpwVcwADojUiPmcPJt
twx+omWRFB9zBzJ0ykk+EeUXzQX1mghapMGbBaDYfhGGeC/gxMDzcKzyhzK5/s6G
ecq+diPpRT4fdWeyhNEIHSas5MfoFHP2Y+rqZ8HHnps5Of8NlYrut8/QGkNwYiE3
lKAy/jRN3oKfNql3F6w9MoUScPtZRfH5KX6tXl4rmhsDYryLV3iNZlUR/aKrzM7G
oxAtY0MJFBstdxSN1oOcKfx9FKKf/uDOgr1EgCLFSzXke4UQVdfnQKhAi6ucM3JT
USg+ihDuIzgaFQWZxRIQc/sKbysfW03B7IUKVug3fo/NVV4BbHkx3v4VP7YSysG+
Uqurma/DtrJJ4LDbghX0ozMEgZLhszCrXjZ6DnwgnRrFlP/ExrnXpbqWWZljUpHn
ZrlVhtzBe+7jnX19kuXHvlNS+0G/vVfvujogEwXO6Bxmt8ZQNW/nx+cijz9Xn3g4
ubKJsGpXTEHbfmvlxn9T8G1+PVfj1xVk34yEg0Sm8IzZ+jonVYo2Ple+6Dh7JmR5
gUQ9Sy/m/q3a8tLfccLVLeoDheb2ZVKor9WvzcjY3V9SrIpVtBoQv2Dk/fVwd01e
zEHIZyxT3/XGLJtsyqKi/eFrRxLR6A4i8W/ZY23qfxJUCcjXOMG3Bt9kZZAwKl6i
EJveRd9lts1Bk4lHe5Ui5Bp8pAw8unXYIfzYTwdJa2yNwCirk2eKPla4sdMdTweq
3w0eJ2tqjnNcRwXXXZBqonZNeRv22hObnQ6x/meDNByB9wgd9FvZ4hLO6FS4Jlgf
URVGSrtjMJkjf8q88gOq4SxDmrhDJwLV3mQ7lLUemURKNTTN41XbjMtPpnPhdZ0I
f41nf17nUe11Vn59vpX4LS4qEUvW1xmX86HzTvZEMdSMAP5mRWzhJRyQf6gSaSk1
877MwSPbXfnfkPMm1jxs/g/ZDfV3tGMw8Tshl0Ax6VeWbkJrEq86+4SQcE+++HRH
H3//zeFFvQTxxZXIlp+tg9Q2cxoZCB8d2cRuRAv3YjNdixQUROvdyLXaP/BrMMOB
uR6w6f2Fx582YJxLJJ1J5O9q4stdwCxM6+Nb8yT4SixdHddlQ2AYn1GpX2cUcuAr
+T+qXP8LxY8ksPzf0lYsyLaRjnwUFI0bLTOTF/pcBI0skgKvTKe348mo2l/yANzA
wEeANcgRFV6MqU3Qbn5w/RlkmnmuiDpYGCkQlxNkB9ztZT7/5rOywVg9wFKdvRq1
W0JfjiyQ/BiPZM2QBHYcYCiVo6d3vHM+tRg3UNDuOrX30HcHGsFwi4DM+UfXcnrR
YyQ9FB9OcPYR5wrFhqzdPS1PLHN64iWOKMm4HSTdOZ2HGpTkeH+Iml0dFbMtaYP9
TfQ5V0Mgjyl1Z9FuL8N5MUfjwTexkHCcyELzy0/jkNtzpawINN1TOJlK2TDLMRwC
M/SF9K03uziA+ao2dy89XPOPE5Xs0rbrRTpciPYrD3uLHTpTIVTuVTu5LlhrbPQJ
4B5ONMUuWcavpETu3/wbyc98ZNnijzNftaxUC7vZ8hFK7zW/Z01mXA8aYPihLiBo
JwcmdgJAkzcmnv8UtFBl37++V968YnzZ8RKo15XrLlJdU36cVPtVssmWONjTAWQ+
rZ4cFVQmBczb4Yel+LMKEwzv99L4Wp/ojjH2BIU1IZeXKdk3Q88+dP5Xy3LgsO2N
cvkBpZmL5F9hl2VBO4WLgqiWconbnlYHVaAhz3GGQHuIAESBRyaVcPBYK1s6x4yO
n8i2lm0ShGO9qlLDheH9BkVAWY4O4VO7kU5oBuGkCcU/RG60tBmM/nUDRVmbDsqt
EDN6V0vOlIJvdWFvp/M0lZbU3HCY+hoHHliOMtnAGzwNafpQtxgM5uVdcSxX7jWl
hT48H2+LtPoBmeofjm51QB5dsZrEBbIHNQcPPqkm4uv5Y5rFyG+c8Z0ogB5pVQU3
7XDiP+gwh/UyIP26naE9PbgM65xwNSZgHfMbspCIrzf3u+vAfzBXMPbS1rYbHZd3
/Uwm9ad+ASH6OEdsXdoZX5v0M2ibOloOOwa9IWFJxQv+dT+WGoVwNJ+jpuMlpLse
yuB8FrCYvMztSRMNSxXbU1yshfKpgR98D1V3PTyjYx3st8LOPZLgI/kOU7FTnQwr
1X+ArVtLnPXfde93rKnIIBc+MLXdvlX/7M2TzndCBqZTaVmxzQpOxSqBmRny/Siq
p8vSHy0B6LAchsbufXSQL6qtFyeHFC5YEhBOoYWsr3e7pYqxYRw9fP5QLLYLdUtG
vW2ng3+j8Quv2cjtpTGswb76UzgO1HUH1zEsVXJxr02NAvDESCR6tCW9o3GpSMdI
AxLLOtpQBVOC0jGbBTMCT50ExNXEAfE9XqgNqPjurZMEZF7wC1/GniHAxDqHhNdg
/PeHVTivwufCe4o+MsY/614eL4VOQlfSfl9Kt/wiqJs85VbXiLDh8TyPETe2vn8V
h/xdQWMMSpvnnfZen8IEjd+3rN8rHXIJId6KcLLgLDdfcabZLVv4blQ86vcsVDmk
FPxij0G6Z1Cr65Te/JFWfdEAjE11ZmI326kbHbTsFgu7DVFS2FL5ZLtpsWwwYKxS
I/+0qzhrUfcrnBQxCqZ7Gt/BoSsG6Uz0OSkZ2sZ3Gtb/VGcxsFWUhg4Us7gpJl/U
y+L+COKHQD3MiwHxVPn4/VCuzywJg4lIM27aGImahe6EqeeEinZl+FAdLoPjcMoc
h9DxVhkHHsevJIgWTEzBzKx0jVEDiUgWUvQEPWDLmWiPb2btfmEdzCf5hcFqOT15
b0ZoyuBKrRHUl/Wt56BxGox8QsQerd4x1BnBX04p1nEVxNduLOwoAv404lwV6puM
dQFgFrj/evxkDkEUfkFD83GRc/z8aX7e9fJ/5v9fvMUOImoA+7cFoTySogvSVEOx
iW16+6fTw/hr/Ic+qUYYPS5ZUbOjP5pf0AOijVEXLxd25t1/YvA1kyVFyLxOkGEq
wXV4CBE/Us6LxglhDvKm+7Xz8q9ubqIryiNlDCvTXRUSKWCz1feXJCJ+1cjzgmGq
XTm4tPAQyC0txuDdW+jAp4+gJIgVhcPbamXpgdqljPSpzI0OtWt2HqqvccDG6qdM
RZXuOE3VAFtDtihg73Jkh9vAndvikuv1tadXIb9CRY2GagWVb46q2igM3xm7YbAo
zunyh+t6s/BYcLlS3hKiexamtLL3N00Dipp0cR4vtMjLc7/H9wL0REE3pgIkENmL
iKZaI+MP7Mi9Yrdu23r9laeMlO19m0ToDQF6czaVpmkvXFfheMbRCkVnYtU966C/
O0xujpgoT1+YyRg9R+WBFEMJdP1tR6p17S9dhmdDKl3z+T92PqIUujOgmDw2RUyb
0BCNQoEct0qjyXl/mqJVTKJwAiQWzwCJHSXqUCYL96Ihwy12RRFiJrMlI1hXXZBD
8t6Jz78f1ww7OufFco9osbEwuUUjxhd8sjHjz93jbhsn0Hzs0kJF9r4qLYhq/3WA
uMcZQv0ASLxfNRZMGEetHax06QkuRS7jjronebCpr8niLTdoFVEQH+gO9oad1fEj
AX9+CMDnKzqKEA4N7Vypssn8YuSRsKQ1x/c/igjieJ6o1PA+15Fhv9JbsTx9yQt9
QcJ0j2vtl3GmSiH7HOwXcDH6yXuFBX8ZE/x4f8e4NQ4kQIUjaXtrcXRrsgNd+ZSi
O7CubEu3INAepIgc+1RRd8PTaQ3oJCxYGyZsZVmBd20uR8EoQfntZwapG17BCfIG
jifwgIuZsMQ1hhd5sP8GWQ0RdUXzF02HYTXPJV6jmUQuxzSVgHACT4H+pgNhCVoP
d9lCzmo01EP8OSZ2DtDc4/p0oL8uoiysmVTFd1Oqm8KKZ5arcA9Q/Y4jeVoHwPMF
FnsK74gfyZJreLJdSefbkplXtAGwl+xUmUUy1inyoDWA6UCa2PaVdwmz/nIp5oAU
WnoojYTjCcDDaeU2vHAAfXjbraKlH5neV6GagU3LpOZT0wFtYsIVNfWqnYQDh4qr
Zg2jdWJGJbFXurFaY3/HUetKfJm/YFRRtZrAvY6YIXH8393z8tp/5teQhBVQyby2
6707L7mOU3KaCirV18h2krm5ASt7bMVRO6y2qzO40/MoMwXPsD7p4mrnzIDGjwbx
1mtvNytxW90kX8TSHjtBYJQ1dT6W36gIa8ELDTkYl8CS7LiDkF2u0xAm6NwxdU64
SoTxVSYNICZVA9PxUbbBYz4cS4YW0PGMaBKR1H3b0LvaFn95Zn/GNxLuzVlxWhTm
Io2xxkV6KxxBo+utwhfFRiexzPkGVr4wmEduSpBb18G4NgC1tJjrJ/ccZ72ZIgik
gY6E57SLmox7StKlCO9pzh4cvbN0xRbbN2vErCmRNoZ4KVk2JZshfI86W27UU4J3
H5Ot48ELznBVRM92M9QZIdG+XnfivTyATsBc+qAjF7Ev1HPX8XKN5pgf8ktJSqyO
gPf++zwIxDWOdySPac8mIinp4X2nMzav1fIovyVgHhrUzfOeXOLduNTDNblKnQHx
EHp60uFJLP1ZOrUqCCJLpgpzdfEmL0b9dSzvJxYAOgX3QJ4CSIentma/2S+kNMdF
xml7XrUX1Yu+3tPv2FEAqp7VgPu1jFmABptMViTFKmxXoxYJOouSdLAGvcdjjZEh
xLpNDigIoJc6K+ngNf1PZuhOaPmmTRiJUV8vJD3XeVMX2eG0BZ0CIdo+g25gQQYj
shimlvQkmmzZpws7AZwGarx+i5G0CVsDA1H85UmNR5HZI6mQOqPKC+i1bcn7R1h8
1pXnc8EmrZZ1HzXpMVmXZQtxXDG1TeHDE/Alm+KMTGP9HWQPq88/cgoiw3/wi7C0
J7JZ6LE9nzUNHfdWXk7BrvzO19J8VT+xFWaF9F+aOw6e5EF3IXtz/HsMIqtCT/SM
k5MM5XifLRYzqaqCEoajdmse15KmBJFkvrPnVqKBFGGLPGEhieCVbkRHtlFCD/ma
Gis5CxFK9Vtk1jn2H5U0aRDyBG38uMzdwQoZNnsF/uzBrDJM0JdXiQqORa4zkwT0
CdnxmjkHNGew+dgbH2rmlgQ9x8H6LXgQPAQuzw8ZHVCyUXBZ2bPM7pAmj3EB2eVr
YWhY3pB8SdqO8px6DS3fU0mZ8uZPScZh5yOUhX478ilRXjC0TtoEP0O5vhcbfFHY
/vgn59pdkO7zPUYDsKoe6xjsgfQDLkpjrN5Z1F82apO0g6+O0OzaOBL3YmolpiHp
FG647cmu8I/eF5f9ia3/fGynPSFe9IFlFNO0bUBXyn/8wM/aawWrtlU/zn+CjUSm
spAilPgemPx6vHCpvwMAyDKR9fHO/GKUun5ftId7ZD/gEmbWSkBk8z36jwXM45LO
CmUElGcHqTRzGZSHLbwGcUXZqfqgZD7CrjRahQfOcAvlQMlFGz2Gta9hhs4dgsyg
BtiDge8vVW0xn74Cr1rBmzA6icdX0Jl61PdkCp0RVS67WfLdNZ/XifU1GWLnxyFT
lR+ra8pG5r3SaoAxQPaG3NOpnJe1SNQlD3sfwrgSdQZKiOH7/QqqwHt6ljZ5xNth
fx0y2qVMu60WDDgvMYczJ7zYOLmsRNSYxEv1yQVX/k80kO9DoSaMAe/wHZqe+TQ+
DNSaTZ3v5H4Ma3ViBlLBo5sClkyfhpg5nhb1JkPdIKaKJ0xwd5MN+QAfFNqU5L9W
ZDzLqTSZPqCb0/EhfBJ+X+aZGijzr+edyTZGV8Nwh882ySxbbS9z3jpM498rwB6q
tb2et3DyAuzOXcrSCplJncOTDf12A/g0CLkloJ6BF7abg3bukOGnDUXLuWRogn/Q
RXuelwuJZpVt9XiVWHh2LIGslWptj+SUUjCuQEv6KCs1Rl5/wTPoG5Sz4kV+6+WA
P6N5+womNzvhryK8zjCXGpUwIslE/v1GH4eIA7c8uckHxWH58fOCDp0S5YXHwq9n
raBPpnQTqp6HVe9icY6DFl4ryuCNXU1qe3+1/Cn2hD5CN3ofXU+zvI1lODywpFWO
F3wOED8Y2e7OFZfAQjnBqTCWNyLMKER5B/ydAAfaddGQ1lKG54bA8MCZtsj3gnqP
Mwo9gz7vtwMRL44Wx+3x+luSgJlVG4pedoAZIvVoCFkWpAlNHsAwvwYH5Fimy0V9
fpLWsZOLtEQWLJhTb9iDOxHETO/tGqg0qlEB2Y653SQIZ7fWLth9t3XkB24O4fXA
hQ+sNC3cJlw52ESaKtNhkLeoUxE782iUi9C1g/IYplS3iqwkG2KZXTli/qQMuVs7
IrOwq3tP55PivkrbehuwA1o3s8bQaY36/pIAWozx+MmVuaeCSzs0QL7c3N9Czris
HqtKFhZGTVy6v7yZO8cDZHTmUBPH1fv284fYvQp0xMsaR0p7kEuGA1KihKQDWMns
Al3bxDW4DyIcPYYElvlHpLIc8ZllY6IqYbOSVevttXAzwK0LI4pxVDGgXVKzD9KF
xGcg+Z5DP5bABmO1fJM9/3TdmwEufHCYbiguPJ15vambVGnJl2FRkEIOYLMK/MdO
TOs38YZ43SFpoloKvgVrmKF7FkAvDkT0i1u8kAo/5E+3NPoL9MbAkrclSwF2Xs94
M1yDWsB8c10BNdFH1BxF/V6S6W8yCmmrChZpQNQbnwzAxeCNL7HDxpfhZM+nYMOO
8jdd27QFfqNFiBV0cHRc8eDOadKJDisWRElVrpJOE1+m55xw/sqJMfCXq4rlhx8n
0Q8H1zN8eGrqTBb+dM92TifoYGoIujMbRX1qAzZXlAQby1bNEmrGmqw8W0ijAEIK
SxrrYL3H6NJX3XQFaxS1c1bwQhYH7hfhNsc3PzW3A9+Lvtb3Yg2l4rPgYZqgAU82
GriW7CZLUVrFk87252cHFRED4AM7ChBtJ1GrgUnZErkLdWoJwEBgwmJ2imn4TLWr
ooKQhTmWapPSpsacc5Ns6/r5mQhlKQ4O3hyDBnVlx4vc9ZUrqQPJGTqJ4oOvEJt0
7rcAmSCbMFGU5iOlEFs3cNk4HPdZujs1dO0XBA73mIImd3JAo1Oj2Axiy/3/qVDN
48e5ykYO4GSGigXrJP26glNm6YoCZvbyHble1YiGnfaci7ID7WdlPKRBgIMjV5FQ
YT3rBKwInBuiv61t90VG+t5ESEHM5Y9TkBYc673rv3+ZhSSAYw2vGV4seLrjYCSc
6bufgFqXjFbMTBeRa0eAdKM624rnvNqvYRu2YI1pgz2RijwRnW4Vibusd07Ago9U
OKOZqToj8HKeR2Adt5oEUAdu4a7zKpjhkqs9a2Dnws7QBHRb4eoi4mqv7FVFqjHR
DGXG+4UeZG4PyR//pvD8Xo3JunmzpT6cXr0wvGKuu0dspGXcxscXzQ0ZII3qrJDK
eD9QjB4HwLVH0lGY9oATbb5mF2O/sYKy1nlynW2X5DdfB87VOf4k624S7vjSKYRh
XAoZnKXgzMqs/AJ1ZljNX14XQENdHS3G8njoCfXjuzywUS9Ac+e5qrUqy8Y9y/J4
67EFjBH897TIEQwQ1lvWLhIfcwNpGOAxwyNb/770jFxfhDCm4yNozGRGOdI3yWfP
V/M19vwvw1x4rCgpnfXaH2xcYxzCLD2dyATPCn8ctN2yjdksnCaHfxtI3C2zZ6xw
pZ7bmLHOgpWphrCUAB9Bk2hMF1GMJxZJANFhZLGtRKQYEQlRUTWvFOQiksgcLSif
fHpkcxW+SfUHxwfTkkAhsJv70Rma3XjFN8RllJEZpOWlw0zcj+Cy4c1KVxNLidQG
Xz28SpCkoxezkJ6erqcIQyIiyUlXkuJQzqBT3GBTuGPEn7eOSHKexeeixjWZPwaZ
FqJDgXa6pqxvPA+aHi9QTFItsckUf7G0nc1YceE2SSVmm+A2cDPZUV4/nn+X+Ai8
v7CyB9GiHEZiweFvh8GXuFxoUkotGGmKmPpb3zKaxDuU8X9SKhu8mW9c/BHuXHxq
Y/pNZzcEaehUgIyfqgOxEejTGCSG+ZSZn3axIXVEZtvzp8/FecNj4bkjd8rTwuxB
fQSZZoeQ9EwnLHwrWk4n61MEa91OnqZuokaPs6lMd49lrI5poi+76cJMjmR1ibkd
E48yT1VEX/pKieOxZaHb9Z4LMkFbRkf0d/DZZa/IsJKMBe6zXmrVqkUMbcyq8z8F
gMxmXx8nCM8ikH2ELaKVuWPnwvITLZr9bX3Mb1W6eo/muu1s2X18KJYHoDhZP/FU
13ApyOsNRoRe49HGdjBfYnCcoAWGsO58hyD7uxIKMvbVJq6vSqvey5vdWjlzq8HG
ic7ktHoNvqDGFoVcMDdQs7DxWQHDQwUoXd/GtiTRUUmPTUNXaqTGqEubFYoqS+U4
ht5XAm5rQqKTRyyIrjwJlFTFLgYBM+1NDwFh91SmgKybMrviU43nntA9QdB9EQH8
ZARZQQTFwwan05htOSlMoEKPuULGx6CKygUwFB337l5LL5fIgwwBKeToaapfiSgz
3R3bxCM4qBk2K/coMsv8JXDNa27CyQxi6U9j8ecjtZup+JZ0EjT9Td0cZbb+fcA2
o59qLpzoI4CxPtDQ7CVYhcS9XCAHDEQhwyINmDEABV7OTWred0qaRhTKAQIALLLM
030Yi/BbMH810/1Mp9+47x4K7+EXkHJfLXP6gwLsRwjD9L5Ojy+0499Bzl+E7Kk9
kbPHdiFWI1wNbdUxuXgvOb2Qr2RIq9hzD+bQbhJ3hKyj5zk0ZnwPtpIsHUBb2oCo
26DZuIXUaETq6mp4vvGZYFgYEj/oTZ8gl7lQCV7B4b3ji7cyIGR13GKe5unGINmK
0dqAj9ck1BjbvdDEK3gWc1/W0OtQydQcakjsC/XVpiURmbhyWlVGKA15h6oqQHe9
QsItS7Y8LYrjf7GsliurFH3tz7O6Bs2R+Snar6C2tB39GiOGLFFyaCPg6O4stoCd
gE/t1nDNDfk0kyfGZpFtS/D4RH8u0hrKAkPOhyLjgOimm0BVkvvN4RmsQ4dOJM1z
3np38wgQUqucpThtEVpbH8sMLweve+QCXb3jbh20U1PJZ7dBvu2oSkXmyqkHaIDP
Vbac5wQuIy8tw0E2UoyhxbFuWEKjLs2SDF702+hc5cPkF5E/buj4H2U6daeLMep5
J2CPfxuY9LaJzm1ensL/hEUlDRPNyiQF17LO9cZ76EmbpvN5RsFQFFOQRKwOuZO4
0j4mlmpwgfbnfECOMKbNbO/JbuRaAUv+ELwKmJnVR5dg7lBsYar8DuWDj0iJWwtg
Bpi1skdZB2u0bBvvv/rMB2bkfjDuxMYZp3+cmhGEPwVCKfl88QDfLU3Zy9MDU54C
S9FfUqvW9TKAyxNb9NUFUga6i6stBH+TA5iy51ObofMxi95T/DNm1o4LTF9t72D0
hEpYTI+8xHpKjrWwj7u6vzAUCS6Z0QzE0RPhJFntgKhd2Ne6dbJYima6ftL+8+e3
VBN2pH74JlbFQ+VT874djjra772hPAGBxcOiKTKQ3xmGXehKiHMtKUQ0ZiVr9OcY
DIiXOIR56VdQnGuQLtpHlqvCGH3n02k3R/+aFuOqaYVZFCNuW9Rc2QlKjia+SD/3
gP+n8AZ55GYuxMFGvKrRxAFgQ30xkAxi+jIsaQ4GMdG0HNPhj7wmilSn8gOzfiJR
8Wiq0pdG0jOYDkjw/Q7Jy1DNdbV0IHgGQ0R3Cf0gMjVCYBLtFcboj3M4Kw554tUY
CChUs0U7eA3DHxc/m615he363cyjKIsiKGzsPtHc4LJoVcAoW1A+mb3wyRiKJxzp
IENDQ7iXwbFJguERSCmwCucFAaLYWaepBJLAU6lQrFZ6cNP/CHCb7hlc1kGBroRY
Fl+gsL8RPTGVP3jMAFWalIhrL5ia85e/f9WRjA6i3DOyR0x50/clLTHmcobY4+0L
5tqdC6roo+gKTdS8wiAAQkRlCfbCFQNEgMbJpAvo6RvcLErbp5JWxykyCdvhxpH8
DcWQAkvXNMPrti89VOmXm88IXWTtd5CWJqs1izV4TUvx/KmTCfgzShGAktRxiHHP
RulwqKEQWW17Wq/biDvomYDx5rKBAjjOJ4SDclOASBISTp3ADEe+IScqpaCl8iKb
nTDEY8PodfQEKCF5lv7U5ZqVYcsRlg3yOJ2ziWf7QmtKHHLKpljO7/o6hhD2T4Ud
VLKAoGRPiZXPYnzH2k2ttrbrSSqhpVF35U4yZa72d0bnC9alBdw+pCErcl4ulnbH
zuVLt/jWkBeq+cpTCdsmFoblW8Y3P80rKFDI0X0zAqpgo/Rq9sWCSOQXkzIq8bbD
d2AkzvFYOpaYM/B7Jh67bZxglJVrwvQqKUbtOzK4ra4ATZuOwfU31HTCn8IL0USy
5n7LhGCEx17CmM/1cIqmgDXG9eh0Z/tQfuYq7b0upaCLdeL6DPZHi+OmiowUPyMO
BRpXSly9zWKATctxECO7SrnPVTir+WYRlhKQbTI/r0sSnH02EdSe505Uss/H8dBt
8OHRDbGNDCGTCiOn4T8Gcj8Y91ybQv1nEmk5n+nJgXVbSTdGHhCthpDK91SjdUOp
Eg6HRBntsIPRh03z8kbAaEUInWeUOZBFiy+yZGdC6qcOSDwEX9TikrOUORzxtmpy
fA5Ep3npfybU3vIaOY1JSDiPAvGyZlm9Tu014uuxm+qGtFqJ1its/Pwa3qmcd58o
c2L0iuHBexxK7+0KNDMMV2NqQzhAzY9cDe5jy8hA5I3E2ajrI4LZjJC+Ex+WYA3m
xxZnIzg19YdAt8hVgjWqEXwQkMbFEkBNdIzzZVuCcITRs78FdOSzucM1veC+pKsF
uZTrilYb5dycIkWW/CsAKSyIYGkDfD98KfkohCscOJwcxmtzOB9Nz6rsZ0J6rCMk
I5UopI4euUyzstWQG5uSX2GCmMGJ7CdLHC370GU+7OdIgFP6qBD1jgc35tTgeTO9
R4SfyOg7sFyeclFCpXpCRjRshB3YsmdiSMNmtbUqi8PwAqKwb9NjLCRMJntVZw8d
f3JSB6Gha/RSS+D/Ex1wY24fJ5tfUyXOQeGRskaI2BNvfFJo4bV8/ViBxQR3ONvf
9k+RkwXsa691pJIZOMT6NmsrWAfT+qZlierh/i2tri0asbqwwmaa9303UTL0Tz5x
qxiS5BbltM+xLfXzbB+iQM47b8g9PIgAHURl9I1YeNRmouhyc43tBOJTDtMDybkz
amoZljITAnMRUbzyAoBTdujEgzfRfQWCTFcP759J7A2JBwtE3D8PGKXTiHn3mqlK
ZrVojIBNJ3bhIAJczX6CpBnaUqYcM997hDmCvJ9FBS5llgoePVtwICqLn1yTnq3v
YFptRgfgi43OV7MrHeZpfMf6zrKipTmF+Yu+izYTVZ3WZlLUgCQlZgxeSWEUiMN7
pxvQswEgNVM2NewJXmGya3wkGGbveRsjvog0Sp4OC/Joh3ozaalUxNrFXccTpJzu
2aHVMIGBTl8IgYZlvLyVWa1/nDl0vp9BG5+pvpVaT1x0KF0jgqinGna9sIPVwfPK
akduEQUkkbyxtOhYp/ErblYP25epsiIvu569WkWXx+ikDawATsxXM8Y8YsvgVyu7
9kiU/5fuk8TaAG+xfcf2rt79UgleYSa3d/2WO2K1FxQfJpYyCnRN9NrqChHOGfqz
Jz2QxL+cNiOFetcG2yOtQMVCk4m00yLGkefscZub0DI016v8iE76sFABAPVGd7U+
S/wxuIvlaIMZuMs9Ar7np2GEUZli4PMAYj2KxO4oXarFYbc0u6kQrellpGv7aLph
C/oKXWTzlSnRiU/wR1Khkyi3Om28yR51Hy+XHPCT4dMNOWKItyq9VOgk0Zp0vI7q
G9JL0KzqnwBRqo4D1hHvsQFOHJQRWzEQA9y6eJWIJXC1U0qUc5+P7o5N/zw6A7Ru
Ub0V5dMlEtY1dgbkdtEySru1G9gcO75MQeIxxXPdKLgM1bwRV5AntGVPRdMxZwoW
dZ13flxaQ09kIeStNsQABcAeVP3If8oKDBFCtK0Bk1ATizwhv5EooBSka7M6OUMq
TjV5pingdLHcL4KrY/IH8PCAde1JjrKC0tq1uBz+IL88TWVGXvqnljONjJWYc7cr
wDKjbSkmDyDip/cvR968mtiQdzaJZTDCjMpwzbvLWHYK/Rog5PR6p9tl3BU1MtfI
32OxPNF+FQRnVxHgjPC29CtLBpy2xcNfHDUnk8rWnOWNUQzxAjjjQb4YpaPZ5AVu
00d95w7SXy9PRyVYYAdWY+MJgM51u1sBJ/kQ8xEFUhXGxQ+RStPm6Lem46vChaBo
gcGPyPIHtKZihRzBld50plftX3bknrAyWDKtAYZ+l1IG61o43YYSS1wcCTJM6Kbx
ZFmS3tI8HXLqSrzdUMeF+mDetbpx0DVNwWkvnaoKZyZhFFOpUTo9FWVtFf03g/MK
9GTP6d00vMORW0PzHqydCJAKxvbtsGfSN4E9uW4o2maJJ5khnWJ13omBzzB91m4d
3w7WJVHVxPeT887PrnhxLtK7/EbpPwEDazWpVSbaVee6TvlXULFJWx9oPpbV7Jja
5hOLpASsfoVNiADH9PAWtotEF7pXCPVzL5ajKUfAckFRZ9lf6/o/k9Qlv3kQ378t
TTo/bQFQErGglmVxxsqyYYwS+d1ELwigT/GhmWSD2p3KbKOFFHZpsJShstilIX5b
eyZjTaJnc+kx9LJ+hyGQIx4WfXvVtXo4mkgwMBMmTOjQ07bDh3Dx4DGIlcXdfFbW
HIHZ+YHpWDtwfNkk8E41EXjdyYAznp5NgedtVMbRsX4PdQaZPYKZ/BuhsrJfeUdL
FY7obgtl7JvW8HoKduxXMq3YAXk3LbGZ5X0rnlFxNPoJaYqyUgfDkNqprRBi7ySP
VMwE8ibX1TsQw0MKV+WG+ZMFSUPxoSBSnSUVZjnpGsuKyw0lLpswm37KBah/WQHY
9IS8DGz7oTbMBhHidAJN7EPIPWi5sL94ZFZUUAsRLsrMQVzytn8iTZG1iGVc+ZpR
en9MUGLOMlKOPX9U0XEOCpMEVDAa/WE3S6SBOuBTLvWqtKL7BQ7BUBV2wO1qnxfY
E/me+kRaKhBUzEYg7NiFWqoX0luUsdw39cLrlwm2EjUf1MQSx6sfS8p3+Owfr2sw
C4IJA/77iBO1aHd44Bx2bYAeiL2Co7NRF/jprKkC2c7JGnxsV1/UNAHL7pJJicXE
u72kU/XLQgSgmb5FIOCQfGuk5s6FTB3VekFIh7QjcfS3m7uOiP69cZyYlwMOQIQN
AOA2AGp1GN7eSuOXukDuOKEJTJRmlsN3JWjlm8NjTLVC6goPQNS+HKMpf/nJOJSf
PJoy2p/5y134cei9VVIOIZaeYWo8nUrPbPlRLKl4cU/iEMD8qNIKLfF7KH0Y84El
Q6MJ4lR36xWDXVXcYKjarqO9vlBldyu4pH8jWYGBYBd1uxLNHhbKAEqoiTGgU9+T
CGg00dv3pArNEXEdT/MocFELqBM45ZYnjWcBB5Yu5OfgLTMURgGgaRV/mIBwBxqj
vL5Eeg/XNS5Fwn+XNEsiSYtGMkTsYvNVygnAB2PwjzBE0fyQ4EXlYEhEhUlhCj+P
xyg7IIo+b5cy84bsLGoetpHgwu2Hw3RMoaDBCVwi/w5x7G4CPLMXcQKj8Ni07lIQ
YKk2eOvr8G6sieHJ3ZPxm+3CaGr9rU0gXcn+976i96MKz5k1y+oUoT95lAmS4J29
sPcD77yhjJKUptrYXfW3h1q2Wt/0wiz0GWE3NDUk8ouDxDNalmoXvxq7dkR7PFrX
O1J8O7BJxNoiLlttHonAodsRRXRSiq8n4c42UWR4cguyIiI/PBHWLEq/+VPKXqdw
vjLgb5aJ61UPacz585PhC4rLSS4OReS0pkiy47ZmArzF0z77gdepiHGy9O8tamvh
lmXI0nVAN1m28CVS5UHKOFBWADpH8JXvLUF9vUu+ce3uMEjfHS7tr6qluGGzIrhN
hxZwc8/GGe9h395Qkk6AfutMXStyKIaV8Qp4MF4qwn7j+TNmIOAKnKeQqhiGRyE+
fkWGZG1O79OdgyBvhg9WqvUkCeldwjYyCbyL2WpN/oPXgmv4HZiUgV7XlxkmVLdT
MYgt9DaiHhScSoa7ta8/LBDZ6DQafulCephThxcR45ReBHH2+MsgTMWT6u1zBwkf
4kxxYOMf3fTph/2G9QNwf8sqO/88nb2aNo2IDOU67APqGt2nMXbzDylG3WAijnSq
TWtaNoVr584FwbkJCuiKsZ4c6Zzl9Dcarls+9X4wgG/6Fe8BbvsYh1EKEH/lww93
VjvODny6SZAwmUlZr3aqPcX3EijEDl14WTJ91/SXkneqrAcb+zzUhbOyk8/aJVmi
PsYX1NHAToAxu2iLzXELD6cTQmfAct1+P9w9/RXpVsrnQiSS9cdsjckVTekQucrW
tiKvUnt7Md9avJP8g1tQ0brFRQtbbmlqHQzR/lxkQilXt42gnTBwBX6lmu+iiP4m
1waYrtjMvfi/JNrk/8XxvE6r4s1d3/tg/cYw/HbglHnnUCskLqPGIpgiEiJvHIte
pzkLsRCX9PtW86NZWlrWxbAyq1fdFNqCgwdiDeP49CUbhJDVkBRM+VIalMG+cP8G
bMZVZ86kUt6Qrl6pP307V8GzB6aX0MbYyn5lnEZUr8wvcVzJ3XK7dMB/SEln08iz
C3jhhNFukv5hgmXNPK1VrUtMlv65OGz19LOWvWYjslgtfvjpnbAv0wjDGvhOI8RP
nmCkyGiMnpGT6dftoKxijMGDvjhLH5+4b79YZXPuhCwYdJaSbq2rE8wFxo62DCI7
l6XxGahV4gop2efCSBVpitIqEzxCZrg54PRHZU7jTMdp8YVPWbqDpgBl9jZqTVtW
esMo0dftX4mr4yMXNW6mjy4uAGI3Nrxo+r29N8xpk+PFUmLEOryaap0SQ2GQBpNX
7pCTV8lVMX94muzHnvmZU3+z5WRm9SriZU5DQ43usKx0Icxyv3h8pX6ULO86BAuU
Fx0wopDxVR/OZys+75Z6KXGvXLRnK7Humm2j98TmbH/MjceladI5D+axs+aHW2mL
h7PpL8zJQBxwmiRPaucYOKGxKGqhRkDZk7c/trSVB6qwJ2XEjNqVEONhFmOLvkdt
PaIWsh/S1p/zfo3v5cXn4lHFfTnVJYjPyqK7dQ3tuwLnXbzrkuubgp6QHPa9JIbI
nEwVUX19huJNHXP5U2Ve1bWwABVv0X7z54Hc/bMGW5fDWjRlFptPPiihGys3lZij
yCzezQ2B+A6u7SuvMpsTXSyhw5Cg8JjT4TTMLM0S6JYIHF0t+RFr/SbbpBnLcdWQ
9Rll34w4weh04duzoPvmKW/76xc43GMTun7cVnHgeyQOvSXEd2LWoXpyuDoDKrvp
8q1UBLrlvdToHs4j5UxmLZc9gIg5sTpl9xQZgNy+/5TNTjACybpIUDCI3jNpsaie
skwCqNuKm+0HgzUJKcwbRDtO+yjyJrvXoBAsoLCLD8lR3aHG/SIFupvcnb8rExrx
bEAU+ePK3T6BrpKooaYnpjCwWGovOgqLYxrR4asPz0ST3P7q2GMJBBzagUeaP0CI
zN1Ui1TkqaA++yI9V4QopjPfhoakzPMYulRFJG42bcj8WfGOWo3iyRqig+BXseyK
l5TLj34O1L1bNzcJixRBygNjpYwy5xHi13nUEPNtpUNM4PYOV4bQUUkNEwVAvovR
AKafB6dkcKCjBpI1dXFKEh7Cs2cdoOjQ0v5qtblzl+1KZi5cVY2A8f0IsZhwfj9F
NjoTzC5kYHyFE12oQBciZPXvqrlR/ZsjdvHCdYQhkDaJasPRCyLR4pMhmUcUGV2K
cztj4XFYerM7hVGbJRIbm0LvXt9F0CBpJksIbhBqTk75Ewnvzu+dLkSfSrmNI2vK
8jdvJf0Y8JC6Ep7D/11ElIgrl3bWiuxRb43UiFNDJmKjvvBhGI9AfHXCU3fCPPGl
n93Cf4wlCvO/Zmp/F2Ohhi/dMC7JT5aHhxmLgI0d55D4jXIsZAIsTBN7h/l8pDNh
g49J+uIallFWm4ZLNsWvHthCaCjmxYUvUIVjCJrZG9GL8oXx74MJoKzucPc5nytk
18H/mV9IXxfRhc1BwZ53orc62N2sSNzV/CdodvoOy6ncpgDX2CVRrjDDbZkysjAw
//xbE5RcDSJpsWnvUFWm/5kbiNeSsoIaGXclEpG8fZntTIrLGNeNcqf0CNmZSz9i
jEe/yw3rfVPkykiIlMDBuP95n7c5RuA32GXc4rcq7eNaUJAhrbuaiDRplWqKNRAe
WTjGh1HHrAG9Wb8IOoAT+VmoFN3w6RDg8Kt9KU8ZAc2xEpFAJn992dZKj/NGX6Wg
aV0SbFjLdXpFf741T1d6KraPnRs6jDgACSnIXBaG/FXGlIAOuqGpfuz/aOZqISFK
gGa0re4wa+95ZBXzdhvCq6mlFA6GuYVBftJCBTxqxSuUiLHw+qWe4sPSCIbJoYT6
9/gzsqrAdUelFzbNGNuvX5lUJkFbJSalnHbFN8pdlgSN23KQXlj4B7FrhRHzN8NB
zTWfmGkfEkEj4ZrLEu/swBNWrMS9KPI4yD2GiAVwu9n+2F9MfIXTVH3UCX9G3yyH
DVqoXeGxfEyvR+AeIjlXimRBUfVGJ48qly7VPHtMz5IoJKOOE43xLDrPkMlE4dDV
gx8wn5jOb41QI/NTQoAIoUuUeuJbLfYNzgRP3fo9QJ8hUKpOV3kDysOeMtXv8FpD
NcVDcLcLumv3+8ws2p6JOfDrIJdg8LrsUocRRfifJshx6DkkvVvpOktK9YcUmST+
VJA2B60egF1EwhKP3xiO8DaxWTmnT+U+5E/g+T1eQH2P01DuDVkTYE29BfM1sALD
+p9N1AObXI5RImDb1t4VXGZDIKWsARi9+DCUvcrdRkj28D2Z8kt54SypzJvFmzCL
gS0lxktkVIoTheXhBFJ0bBAUGTCNy0LhNgm/9fS7RQPoZJmj0tTKZd/D2oaM9Tct
j/KX8h1ULBLkaBIpzDBd1qfgdSYkgGoiSB6e9sA2FjAn8xRBMbW22ws5y6nDJsLI
rpOdEZ1NocLB4hh3w6cI4XvtAqOWArvjUS4YaHa7pVEWkFNeK70e6HXX+fVdrLTK
iWJDmUejA9ux65ki2tjQ0YhqbI0vl4+Xbm2UXFkZoP8yKwVDsUVXt78OWYfS5+eX
1IKHZAuxaGW8qyMXovvJpVhKR0oBPNWwYbdiAC6H+wq8m3qiIN77N0303PYjLscL
Q8HUvZ9HHzTXVfsM4fMuj73r4kx8FIsw4EZKR8lz1B0fRCYUuCJbFZ1VLsweg4pV
2BVyvb10VnRJhGx0PRk/xi+uuhJrdXmnFnXrCKi83iqnaaqtGDDvW5JeaNI0iX1o
RhxNxPbVY+I8JDeoKidW+3ZMyOo+TEBdS7C/34YGRAM/KylnLhPqosbRmg/SZ/ld
5zTxDHnf8vtKCoBqJAE3DnF5LJm7KvtyX40UFXabGSZrzsxQw+g2SmeQ8kqR18Gj
DihPoL5ZHGkiYqZk9KdwmbN9VgcIKOd91/GJ78edYi2Z2s3YMYIWakuRbS2el20a
SrqJZS2mahIOo3FQtEGmZGIfYpchGeyKELOJB5JxvL60zjTfA7pmrWv82TpCJJtz
RaIa4JEcOJPTQZ9TolNUSGbUzw8jJlGaRfAfecf8gLbHBSrM2dqwsLyGsx0KWwlI
HhltP2Pum3hGxSiLk+PCrZeNDPEItZXwYv0lkauRy/xzVDt2TN/CGCi3d8kCn+nf
/M5+DbNDkWiSV1J21KmIYyQ8diI5RLxBO8qEijPpjZNIX347+YowCR9M1aD/tKgW
w8Eec9mveHVgZLNXiStNFKVVOFdhbFwX7eENMCV4C8jvfeq864o9ndSoI0Y8zQEr
G9oUI9uOPlOCzj8uuk0DZSEkF0Pk8cPTeW1Dzrt4ryfWy5W/yyAiJLTXvGxiqKpO
sq4aleVFY9az7rOpWjlC9mnHK/CFIgZJYQ49bOZDPpPYrJF2K50vTpW9BRpwb9BG
S77M6byR6Ooa90864m6KoYDJveEJ5jF7f6rAmNhV7lYDDP/fkpZlevB2qxzK4rzi
n4LImigLDm31qUjBZaXJtuioLg9Um0cX5dJPH7DXbRXa1W+BxGwTCcNOmgNqQBcK
blvY2J5QlDIWHgAhqkCmsC+rgePukMHdson0333/EvPsOGo/NV3b/XwpB+/jMoSk
KA7slS6ozC9j1GtYJ41XYcUDDAimq8jkhWFKStp5kTQv5NRmaz1YDQCDQD66q1LF
hDjQhOYEjlZo4GgfBiGgR3IoTDWZspcn9gfRhL7TcyoeEy5ee0T7FpeeGvj0j/T9
nxb2Nm4KwYbW5UcdQmdXz2Zhrwsj/Gam+OeEBOcDvReLCltVqllQ0mKiPvu233N2
6hL2VXmfUoJOYj3/o5AoCmRCxFFweKMIltGK8r8ReKvWAj1JIJc7YdOIjEYFbFIP
oTvFgwYXn08lL12kqJo0N0lt3qXstaGu6Q2iuJnAGaVspV9XTjeGTSj9fvZLUdT3
5N10uTvfI0OEMstUfyR33y7Kp8BCpdZ4cds+gTBuXp3kpinNO2lv+U8qWyesqo1V
uc7J/64qoRo9loqHzOkzZB9di00e9icrlo1r4YcNt8nfySftuWvim2K2BORyN6/W
Vbuibclt88Aro7AqnEMtO7LzUfkdSjWLVvtxZurdtgo9ZnWT6raubkmgAragPu2V
SZsF8aBvdeIn5YhzxS7leOR3/o30Y4ni12D9yH1v9Ne/zg4WwsyxxRgEhkxZZTxW
ABUUsnXBytPcrKxUWzlZTZ2MA2UwFBBGWqyK8c+lRlSD5yT7qdzkLxhQCodC3v6D
DGphDMQ5Xh63YD2+Cy3GT6H7jiSV8A8W2LKo0YAPYPxfr8M1+isQGvh1fMSfm0fJ
3kvl9ZnRDEblEnE1VgFjAmpGuq6NY71acbnUmnrsbDku7i+Fa+gTtNKX7BoQ31Nu
+csAjNO8MsttkIN9Ir/7Di5gtKNDMTwMGt3zNQ2kg1+Ohb1Gpevl8kCOaKU4fj8k
pQczYzhcgN5scCz35aLQwh8jPuZ0ynQd0broQfhkSTykOUEsBKNeJVAE5KXI4rl9
dQLhKVwbnIhtx6TaOnRI4pcdi0gPax/5MeBD225bq/phnW6KFydyQUlmOdRa5UFP
JZuURaF0aJ8qWWGtZrGaSIiWMSjcMVsCAgDR7PboLp5tEBAE0dyaZuIJS8s3c6gX
quXyp9Zq3rWDKfNDC7fgE6MXSc8FR+mFhIuxs/USQ1Hiu5KaLVe+fmyFRcILLMGF
ewC4vF9sv0gpJvkRzIcI/TYj1+Vue2bAEHqIUx7dL3M6ZvhDJXKf2yWWDj+jmx3u
NGGatyi3GFjueoq5IdwvnjbweBk/GypHtZ9H10j801l1L7DrIKxYnTxB0Jdivoaj
QDnZbNTQ6Dt3eoh2lhrDOR7dL8SGAIYQaenb2ur1g95MOpt33GH0NDU9QmCxjnbq
AvioqLqBEDjnq+bmc70TYkVBEn4//7PB0HHBn/P2vQRor6tEZabUVEenZmv7Mud6
GRKPTf9Fi1TINoDyuJheHATRxnI5N8xQxzSUL6sYMXIft75U2ApMz/rq3zWJsbWQ
f/aUovkDBaoxN5uF3FQiFi7JqkwRYrqKLGEEf8QKlpsJwenGhBudG2KZh8EQ9hAx
fG1xFi8jd1h/c7Zwf/rVv9W7WijWQo2zphvFx7XLhYOocp1/RLWt+oNVsxedUP6K
svoxtrk3zVYjxDk9MrEsGVTjCH8+BLoFn5gUukn3c698VJbHe0HlKr/fOwJ9iNIE
1+Rqbiuu97aWGrD/lPLXAMaWHDFT6lKgN5aIcm0V+u8ls2UGWMULV5K/5TInYPhN
CiOdGiuWAI9CG8Rg1adR7XM6vDafQMToeFzqs8MGTIQiW06UFCGHaEnK+OSYo6jT
eSVbIb7ioq3jxVKXQYPIh9umzH+xq3lP0GVddbfepLeZeSwlQGOjsHLeCDfDmsZs
epO7Rad13XQQ8Tf6Km55+Kps3GjzV+aSS+LwWxYBoxPhXFgSRvbKj8P/p9wyEocj
V2DNM44uJQJ7vYoUyTzxV1wgerKjuuWXUlytNBoV/DCDN1kXNRUMU+6umMV5vZX/
fVR1GT7oyc5X9NvalNm6Gy0sOKOOcUB5bzbG5lCPlTHiceg/n+imSOXld0sXyGOx
T9oS0Zo/uhm/zajehaOP5p2ev2rvzS1/OKVnerf1b7aC0YovTE8ZmXYsDFG9kRk1
c1WyO0dZQBj8K5EFUAqoYjgmZiV9jkd05iDx4WJRiMsqKGpJY4PLGV2A4wGQNLDO
+ERlYYS5YQ7+Me5Jtcy+TqSG96jfypnm3/8Vci1h2zmt9rh4YoZCp70CvTgrZJOM
PbpDjA+zzD8muS/S0kdqyPXZpdHwou4yN6vQvFnSH7p4hiL5WShmSisyF6FVlCTL
35IaJKVRNk9oYmBD1Iv+cZ+jaIOup4OGQgDaRrRpBST1eWFjfDUzxlTHrMBAI1Cb
tCdgP4Phy2bMLOYMIME3oPNZCGrTO8sdt3XW5iCrKpmy6fvhXj1XFKRraeNcljKJ
CFUC4QL/Vd3TtzxqDP8Ql+wQBPESkRVH0OIFcQ7da13jff1zuqXNM18ekkEtXTbi
2/A2RpytYHNOuKzsWXONvIMErYtoOlzsNg+XXuUhPih6wobI3LH2UKVIb5iNstQ6
nw+o9/+5KYfjaSZh4wFy6/GX3T86tIPpLmeI2QACe37T9oAwmLF0055/HxklHlHA
O74Z93lpwZcJjSI5oqkFu09V3VceWiJ7R4ZT7hiGHnB5NMD9nD65FgVRqwuI3UTx
xSxXMVd/Ai2FD3dupawwUCGwbhi/AoOGW3hKM4ZiK2tPIk6VIV0yH6fLZRKPuI0m
Mwks+fOo6cNcJZG4GG/lV5Ny2CDw/19wzjuYrN8ocX7TZVt1/KL/NvVzIYu92eqo
k6CcHJXSPnys/+oF8dki7NbZGA346t6PkuzJO7/g/xHXNnkAwy2/e0lxH3V9tB8X
v0PwZPPx3mo1pIqC+EbTGQf+SHXx6E4JPqAc+9xPkLazJT+JVX2j/6do4i1E5r4N
3PH3wKes/EhUPoZKzgCnyuRhPtwABqAHCeO7UHXvzc49cUFYEObn0pRcDTFWeF+d
0rSyV0G1mI0En1zwZX4p2Cv6Cee3LlrEvZqXmvtyvdOliD0a0cnfeMVuIns9GMGW
/khVIlWSAFQdMuft/omSzLk7M3zfiVxDU2c6WGtd0djgn4mh1sqFvvhcHmTTx310
n5Zgxh2o7tehHNbRna4gKNliYEdHgBRBQbuKUFcodtnnVEqMG+tYJCHwzXzWari8
UAroq2m/DnQuWVv6agpQsaBuJI8ubRoqXpxC61MCtX5zC4nrXLFbw2FKXvAhhdh8
D6p4QIvpTYP7+KzzshlvJzBU7sTmqm6/sQ5PboXFM3ehYCS1vo6M7vWvJyXHcyip
uEFDtbtJggT+CB0U2lTRDKuJhEn5/UbxapuYYJEfQSVerVjwjDZvCMacdcUTZas+
GQNFO9x8n9MWlI5BWVgqNb/FP3cq5ViuN9UYq3cUOg549l5231FnW85JZ2oMx+Yt
aRayS2lTgE4gI1QcbELLL705WTMcDu3VlC7cN8Otrl8l3FbcAAMI2V2GCbADnaMm
1k3llAzc2O0hD0ip8J40l6E3dgL22oBR0ZCkuQ6UpDkBeMSZz59QlI+iMYhjca6A
CuwsmojsWrDeoBlhwcj7glou8GQdn2E0YyZ3lD3ZuNtdoxeC9eEqiHT5eN0E21Km
qf+69NVCXyJAR/6RcYmVAyY9NEetYicxp4+HfDc1OZ2Z+zIW3v7AOSfEAudCBNth
nRMS9UEFTLmbOeNLtX0+hHwiZgy+xJUSZt0KoZuSf8szG7h3dPt/txGPyYSOmr1a
5OQtprSTt11FMkDn6mFO6z3l2ZWGvz+ywCjm4ZdbhwIvj22HXoGUnpkA4XIMDkbS
mETcJ7TYaS/9myUD1UYQpl4L5baFId0+QBNXpTOv9O9J6yBb0/CoTKGJhnXbIg17
9HYSAOlTDRbULbLKde8om6LBhYCtLr+te/2IQDv9BwP7UaP5FLQMtvtYuOIoIkUu
l2WP16/0rwNO5phdjB2B8C1VzmuOF6fmu+ryVCPWVaKMlyfstcoKLojV/fb++F+s
+LFKRNO+HcP94vMeBzAULlOze9veuMx02Zmrle8WOQSTFy91lf7THl+iB9vP7WAp
aOyXO9j226HztoaPTOO8TIEvTRSxmvswbB+M+nRhsGnrFqw4A+Py1RYG4JO6ctIQ
m8Ra3ZFFs4Bvn+P/7oBgeprt5XcXHpCXXXAofWuYmJ8h/wXS6tJPaxLoICxSxQ6P
lFyq7A59Px4rG9qj/Mg54DBvZy7vdLl83Jy5ChFZ78QqC9z9o9SPVMPuc6++lhgc
upRIqvF2OEqO1RgyIpBL8Ipc/LvUSak/H5H/p5JtMznw9FsrBHceKpii+1UNpGbV
QTLFeKbifYYc85twlyeyuxXJIN/EJNoQLg1OVA4Lwbq4JtB4rgrxxoy+QVzoHG0o
tPM5tHGbkKLH/CRIyoRJq2JF6zzthWVbSRF1JyTNFNi/RPE0n/sMcqMCto66FfAo
2gT/ssAefgHgypvBX5xPo6ZpSyM5rlO8scqBVbU8fL5JI2zU2BXVOohfry0uLV1x
lypgguRynybY2q7gDv5kWc2ATOYfSCnkvAJgUfDO/Rt8qmHH8UlaU93ZMVZ2KqSk
xRQk3G0DFZ1eFASxcCCYfVkVeCrp8/3JXjwNok5nhvVD1zpogFkcHzXB9xCYQosa
5YKeuyYoxV6qqo49epFgS7ifc6Wsnl1Jy6asO73VO1ZiaNNlGUfTKieh043Aql4s
ZMv/k1/UZRFXh0+SOrkmlFHFBYFJPoPKyTTlIbxVCiMVIzv12dr9EznyTeXfCLdN
IWDpupIT+TFBMCLv3WOI60PqgiybtqukIPyRHPVJAeyYaYOW5UYQBmQwenZcI8Pm
UXP9N4dZvuiYMYwmTcCXwAOdcLtr/2tmg6OmnZ25mnyXyO386eNuSVq1ThsPW0w5
cNKM+hgKQPd7Za6xhE4XeTiIfbKewvqcQWAGYk2bwMUUeEMyISTIBbO5rSoP2UmZ
q3V8NCGsmAQSPhoO43P+Ev6JdDTVrcjWm8HmaEYDi8eUgFiqoBYlPXyI0WMDOGyC
VLLZLTc4DgqrBWNRTtrP6krvZxtW8/W89gGgEpxMAel6OWfXnwy9GChdnAgv4WQG
v42lgkBvPxG26MXRmZSX53hHGF6OMRV+mrOadxgytONHRTJ8ljVx5XtGW0+cECHZ
ALu7EMp0pmvNO79dCYQIT4WGhZ9Q87Jx4J7VijbEarzalwvRhCnpzhBJeJZm1RoI
a+B7MC2KzfnRfkbS72htkvYldd+z1MEUJV07gyKTu+kNkRrOfiGbhvLTc/nqvwRJ
v25ww8ZcMMiLlDMjnkPXKtHC5EgYYtBTKrDZ7q2pn539m9qQgV/w33f8iQNKsc2N
b9PY0oxBwPk3wwp2sm4mDusq5MN0iXyujla2r8L5bgADNpLes6zxdnSnXaoVUtRd
qNvnPntECWoRIGVotTYnGpCgqrum2veoUlyz+cs88mht7mrNr//KSd010qlNsngo
Bp2hcxkiAAhLBZNa+9+z96XZ4HK/9HaGWyrS5F6w0422nwvHoRZhdaE3dsnJ40s2
ASjL3zJrOqZxMjKv5i4VF+Ii693ey4y5WtGPGF2bs6/5wgGvM/dBoSgZDPfJ6Z7r
moyPZjm9vtryDmpeAoXNwSQhw9c6ve0Ka8N7WvB/N9eldpYrfShvKsEhSNLUNvgZ
n2YgSVakUUqIpqEKCR3qtLbjO/uvCETjc1V1vEpNW6ferHKm1PAQ+UqklTW10UvQ
XPfVwF8Ay7fbsELaGWywIyRhtnqQso9iK0RGL1mYyC6VOAzBDQQLSHlNATZ6Gh1q
Aog6xQJiHnb96XKVOFRJdTGSxCkT9OpHUlFRTFfnDTu0KvRDlgV0FB3gyJIciWkQ
5D7ByW+lBZjQTgEwuLOErZ1aFlv3zbyt5xjPmOnKxsngyGQi2cniGN1+C9YluIym
Ehdo7yliPPU1AsWJJcrDV6VsNXlhAmzD00FAGdGzDV92aLB7QsNMylcbtgvxj2xB
Ucg42rx1mihcxcWk1xMCsy6gVpwM3NJq/DbLuxgh5b7LqFpleU71taUODQv4aMsT
gjQqLGu5L7r3jRwqvcCDM+09PwcxJlT/ayHd8TnDUcEF8+hBfv1cZ/w2gcAKLV6b
vtgoKTM2iUTV3M6zeRw+AYFtyZsokQVysCbJDnlqB8O9J/FazMbGK10uV6Uzh9/m
XRsyx5xednsN/V9AthN7JXs8fcKtqeJAROpSRC84P/fr+Ph54onQBaYJmndN+g4b
LRlAp2wiLX96Pyd6HBPMs5oj68mjoEfdE/2wb5hVumV8D/jLY65stMuFwQ6P9B8m
YEJisl0YK0YpmPeuiJT0vX2PMzWW1ETUD39xM6rUGqwToXwkSjzVEsyyitZFL+5v
IoMBGfV+N2/IsQZ6wCVgyf1od/gKAYCU7jIToEYWEbPonJhS+M3FOI1vEQc6gm9L
bFlB4/JgTXkYLeR7jNJWoi4whdOMIwhsYq8h2/SE4WlYTQXC7mL25SAjMu45IRIo
c/sDhSgMi2p8H5VZYKp3DvEZPVWMovTFryyrPnsIqMt5RPAfgpsNVx7GVzHwQ2Uv
LW7zNHMByPUdmKElFfux5JgLd5N+4EpiTJA45LzxDzIdHP6p9tybRarCJxJG9GwG
mnHt3Ypu7fairwx27mfM4WSfN31yySxn7lapCdxaDnDawtCJwZcKflsNdONNXLnE
H2+FDk8FFbxo7K/od1+JJSUc5aXCCff+22O9uxVlXO3ZB45BYukVyvbBTq0ZnO+R
TsiF5A35XQVgr9wTN8isj3LMF3vHWVf7BuxihKjYd8RfD+2/7KkhfQwOCK2NEIdm
LM0T+osQTH6mnmph5V6qLy6iuQiSbld3hcbLf611fiOlFgFk83diePqZlA6WnvWI
NZvjSCZAR3Rr7HcOZ8AmyyNR5pjOngLd11uYkYSQ8D9WLuagpnj6dmnNz0+sKCWC
qbEcE1ppHGULdhPTfpfO5pyunQXDC6kAxjR0rzeO+2wqDpBgvu1EZ20c9FcjOQVR
OFxDU2q9b6UQkCxEWtjud2hRDZM5ikYWZA2Tnm8rtSd8NOMArKSDX8Ee4YUFcwQX
MBos6J5qnZo0L5Hi5Tfz1PrYPJxxmOGxDkOCtuI/KCKkPO4S0hmdy7S3lm5syd/8
JExbYVr1Aq3jzOtta1KBjiBBlsshsr/mcvdP0Ny1sbXfnOo0FHUGnA/J21q00YLS
p2dLusDk3gK4NCbICBFBBWMuf120bPrV75HngPXyTai/yTORsXw9pUPp72z9tFVg
g7HJObDy+RBwc62BZ6q3/XWo9LOwrqG50zXweG82kJoOgwpEwbrEVN/9lfEuGucw
p4CQuv62XxNhj0MdFfJV8VFEn1eVWy5KMjokbFgheDulYlZakVeaC1WMMhOMHiDs
dCysTiLfx5CcyH+jBqs0k97n0AvIa89ewNHdKYKjhn12V46eqKNCwW3H0nhJAAgX
VauupiB9wuynGpDUbJndfWG1PTPbJ6/2JmDF4WMesZJJiYoAECBf0KSFNS2Y2MPk
pcgdcNiwxAPVYKhXIARew92KRTkleYu7IOiGFokLyalGZvjRZ5YUpBNKVz97vB6t
8rkq0YRq4fiEET0z3YlveQnNl6cQVg0yqsrRDrvRv5ZKOd9mhosLXUIdHnr3+fkk
MF7BnWVpw5omZENz0giPtAYKeNA5d8CVXzBt+BY4jzTK3SJ5YTuyUL2vL7jTgdjU
hcLmJZAUKUzvS9dAguhiFp0FbLY3esuc9vHCg9NI7t2meR/3vkrN6kWbMxCIuIQZ
ngXbbFwXYrZ060AVtMLJSlZQBxTvutjlP/GiCx7s5qFQ7H2/LssCLOC0p66aXJS1
U9Vjn+qBxVoBuqFBmv3PPBVfViyQhJUKTMZx4EyzcRSuW0NOZzJISopfK9OQxwqe
Xsf93VKvnLXSkVTDONyIyLBnL883F+YoWkZPW84Gpcn6eKFP1BJG3Qj+cV8j3czZ
xmQjQSIJkSYvRJ4H24hRb1TLW5g8aO0Vo5WhSi5NY20dVxAz/HayCARdF3HJ0avK
A1wtNpb8jOwIWx+FqOL/ykkyLjeNhQ6iSx6EmUnfQA7bqJYmlkkiVzDUbMAVQSKV
zrTiPKoJhQtKJACXHMlCq5O4aRwY+rfau9z0Qp3LbTrS457vjJ6y/7YEa4Q37dDp
yWsOtwa2BdVuxCnXf6dJGH4lNBrKtBeR80V4HHqCmLTJT6kOfmJ8Uu3hedqtQM6A
85y+CLbKAP9OoBgQfz+wZFJvDueVeTzaQL3H3xRKr3y9AwXKqwfqHBGC3hzUrjFV
VFUUHKa7BgZ/9UULvT2SgySB6+xHrj5zQ+JDn7TvhrSLxOseAhL7XwkCEEs3u+Vf
F0PNhLtq3Op+M0NzzYwKgP/byQL46h5NxTUCuUUXV1pAeGYELuFkOUAk6qO929aw
FCCEKL23WMGvuKyvvwg0LvDo8UHfRRpca7KTO9YB5s3sOO9Q8xOGkFhD6+F3StCu
8W++CUjxgxBCo9vxfzj0Mmto/uXP+uJpDMd9+8fYKYLZj/BwJDfz9hyVyZuvur7c
Gcy2hiasf1RtzxehXFs8mqxppebZq7nkCKsqXW5Bp7SNsHRis94skG46N8rKpiXn
Sv5v+jfgUTkEaEf1de/oPmvnIKnmyW3t29lCQJ9yXgNLJ73ECTogj1K1rtvbvXFp
sQnJk5c1dB0HBERrpOcOR9c2AzMKXZINdpZVDEeDJMr5AjhIcfmWjbxYUfAbFb6+
+7QslSVjrR7BerLh71EXWclaJXtgPX5ZgpWdi2SWJuiMmq90n4rKflaoCXhrJjOl
NFkfM2n75ADUMh85UDVhBjHvlnWah1O2LK+4P2MI45c+5EN/IgS/8FCnWKq7D5/Y
4WzvLPSn0Jgf+YLjSd9yHzptyEyoh5w/ZPy1DWxUTO0Se/PYwMzSS53ZD7B4YCyp
o/1WvlEdk9nQw4954+njF5pFkQzweQcvqrAXagpgVyyVGXA3SXYd3TfC7wVcD3jH
q6HDsI4zxEe4L7OKnNgQZxNozElMbeGmA4FL95vf8aMAj42KIw+/qQvg//txxjNT
aPu6wqSc+EQfdPSgqgRKdtIv2JQwAp0uaQmyy3C59/N+hptYRetITZhVyBQ3AnNv
lc0mkdXAlf5Gz8U7TKVUuR6iXf1dYhUd/KN5AO6/eaON0k/X5UIy/Vt/1EHdb/2P
WQORcUAbfa1LOI/1cB6ULiLBVUPmUYSztPwBs4Lqs1CLsQlfhSfrCIezHpBAaesG
YyA952P7ua1JoYvlyYnznm5He2tt2oBGSqSJhTtagh6Iw0/c3gJO0BZzE2DuiWSx
V6LGVVgnEMWFeEtO57uATAZohrKhJSheMcOC94lpFK4XLZlBUjLa2SRZVQHmXAeV
V0RtqUrnQq/4+P+R5OZkakz0FwT7h9N017u6faHszjuroWpoBJQKhkj/unw7r9Fw
O4z4GAcWHdc7LmNzR9WlSZPu5DftQBNl3u5kq6MyXRsdVG4mCc4PxxydyomY3qCB
x5MCWCNpuGSdkbFGmnYL9JvM9HrfZ5lmjsIqeF/l1juODdkuKQxDe6KXmbwfJTl5
faEhaKp7iDfWnYJpUivAIDUYgXPVfrieI/sNmLKMaKL+OGYtcrXVkZ8dT4Ftqhrn
Nz4nFAfl5gDTpkmOhKIdRGMyYYqKkxHezkVeouDePLfpsbnNnvo8xXMqSBGLhppF
FOx2M1MDKClcQdBZaGYcmHs7MbYwTpf2/p3sGXv3FRCbyLgcfA9mSCLXlW4sicq0
3it6rqcIEf4m3kly7WAcrppNKr0Av0X5x36Nxz9jufgn6LUjoCUPV5gA6CRVbuCq
pRDTRFKaU60cSAY9xG76Rtej6YQaSlS+vuD0uyNLQk5QDw0mKOnam+zoQdjYIEIX
/G5kVkGeVklmgX09T2RY9E82kcXuCz0GUhu80QNA5SylvN3mordP3ZAoYpyvgr7I
JDEgY6iTW8ZZzfNLCh2iboGEiUE8HRlZwvdtUbFCibIq0RrvwEusgbGfkup62j/E
xlD5E/MsdTTLd22o42vz8RhqZGgrEV9f78EmkSvKyPafXNccdB8nbIAONu7NQUWW
DU+RGovnzQbH7ey3oUi4I+UIsCjyujvOh36VtinnuiIb0+apW1eJLpCRh/Hm2zyn
F0DibX6RC8RhNAjHcHoBybeMvQI7fv148GNNc0l2jkoWW4N+Pb0YjP7L6r6IH7Hn
K6bYGEwSuxhe1pEIEsTARnZPckHoZFEZtoYBwRfso/XQ8YIMH0oFIsIdQ7KqUZEp
Ma6c/R9LiTIk2bFHyITfWDnIIDxcD0xN+0f9HA2hmXN5AF9VpMlgAkmXd4nkzHiS
tfHv1Poc8t4Jhs0zyuUN0pOjCvXXFVqv2cJkDfFxlAJ/NScBWtqVPq9saIYiLKlu
eD4umnTpiTIfTR8lUkUAWZDIwdjOmlI6+JiOjAZIUyyq11BgkqenrNZdJFnGxR1+
PqfjkRmt0cWFlMdD/mF8a2txDZO6980tB6BEY580S/6LQVtnK4/mUIUUkfrYkTwZ
m+C92oykGOlFvzLWSzhL8GED/4Znqhqf7cjd6ZrJpBbPaBJLbMjBPLygJhTyLXY0
Iz9wFQHiJsjr9XRVkupkoVZ2NLSZBuCLM20vh/5HApRK+ax9MXEvt7q3rCslh18r
tJITMWlSL2bpOH3Spo4KUwMZSq7NmQUogDVZg8sA7zAafAVnOOrisdAtfVtuHrTi
VDUe5odhmqGb7l5ToTVNO7R+FuUXtG6cN2nUfH73U0DNwfPGlH5B9Trsjdj06M+I
M8QbyokxPi/v6uxw/iIUomQ9eA5Di9b2bMyVLukpJGIxK1IVkQXgJCuGlqjuOTJv
lQapFZ8Kw+amG+LJKEJi59bVCVQNbFuXbPnN8Mm3I4jPT5cyTcUQeL9VneVM3L1t
T+K0DEu5zoAESJQVnCcuHFvf9+wY+PiKwBBWFqxS01belzshyWVPz6/Zl+f37ulI
FKN/ZOFdeSoOQEEFHzc8bAT/EWYzJPElxU8S1I15f8Sl7KORVeCnTN38det6h9xg
zt27Q0p5jPrIq6h+lxwREJJ2edPw/5E4Igfnj+jrwkdVvW/zovEYL9TD3+lqiFDB
Ph+EXoDKuimOEdkphBfehEBHbwP0j1jqbLu6k/MKr0k1XlLf4r3ql48lFTyzPbj1
bX3CWlEms+r1eUTYINdrhTfiu9b0kglXRapoVVTDM3amWhTgvjpyX3XDU2/TSxX1
pVOblcuPqRBD7n0XkZLgadWQvTiY3nmrsvLVjd2jxABNjiNgTeqTNowjUyhd12Sp
47J7iT3v5NqjjE8oxeZMV4eh8pyzXF/v+4hUN0as+pmUE5gSuNHYUiKo+0Mrdqvp
`protect END_PROTECTED
