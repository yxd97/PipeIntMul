`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2h242zF8plvrRE+nBgShHrWtY7MJAozS9tZGeQorU5B41fEVpseX737VnxJzpopF
De8orvTK7ud8/zYQC+PEC5IWGz8Bx8jgoQ+8WiHLCBLxFtwfof+WFikAG+QQZ3gc
U7tSiUDIWVDG3h2fKswpaNN5O77iZtGDA7wsDl8mycSzNPPDUGq6/sA8hez9Md6M
oqtEgFwTiOlkqahzyRlQ5XdhUlryDJLMI2LbNKIN1FiuizH4qFxLTW60DJ054eDX
76Wb7Fo17FWfAkyuQ8e9iTrRFYbCzCeZ83MdGnl47xXQCiZG14zkzHUrdeM66v4t
`protect END_PROTECTED
