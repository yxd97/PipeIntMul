`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RkR5Mu4C8F3aRzCv1aHKwiTn5j95dwPsPZ1GJx5IrICOShJRHHHFsCnVyu0IoacY
zf47eQeOwhqK/+Z5Z3+NQiO8VA5Fb+jRBn8thO3jUbKMOyihvdAitEanVZ0Av2Ci
iPaVnoUyWkbYT7Fkf7s/qbj7EAxGtwN8r4Ppsoe3da5E9kAxEDP/b+djHkI/kKCp
O5dZPbvXWd0CwZHpfauWwWgFhCGo/blMbbvboRvHmJR3tqKZkKcMKSQQftRvJbbJ
xYNPkRnzDR46IzCkUOiz5lFLRfr4IgI5kO1TaKkhaWgulgzH3aOcEMyw4niMwvoo
H5zFPVnLd1tYXFfI+0llGQ5zatJt9VKjU10WDVLByyxuKNNE+CaJu8NhN+lmZMdU
qpQtIjs96T6cVTJkIb9GfjwryNB2QS++khqciPopHOi/Zel7akCYtUFcv0qsitsw
2WcDck8JvPSPOflZqsHHIdTCzTLL27eoWT5XrElhJHo=
`protect END_PROTECTED
