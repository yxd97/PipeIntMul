`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kr4joS7/inN6slk9WFakdyjxpn9/DIQECpi8zKqN4x2aVW9NLVAMrsPIK5XPk3zC
vxfe4HwteNTqNxHwOoNBUO4RPoBg6CIzVbjTPa/nDH/D115q/CWhac3O4fOE9z36
H7woZR3TAto3xeiB0iJ3F4BT9ntntJwfSmW+grC7hfNnEMr1LS4b7bFM+ndb8wyT
dy4vsmQaZQ3A23h+T9X2jDO55Mtvjj7wM7xt2GsAk+ckxdNXwYQMTHHHsB0JQ0Di
4sScm/sG5h18QbyWh2cSz9mEs6XHvQ7uPnA6rYaK5rQH0+LjXeej+JZFymu1LSv7
c9fuTYQ2nSJx01w9Zoe+A4N4cBtBCUSjTBrj8l8vtJVmooCHrUozk0S1vjEuq/vY
KQXj/8vBC8YJ1fuYHdFUVnR4e9ucxhgqfIDRTM/3MipzqKqfyyLtbdFq+dQm3gY5
u/39EOA8JSX4lT7T82iYj3ApNiqpUgnzUZJs6dUw3R7voAlYA1+nLIslHiRWLDKC
eIPJSB51IZE8smYrwWetq4QKd2usEzr7+hqegfLW2V6D7vpYRumes3fvKeBDboup
0beVEipiTX816lkuJnKN0JTJcQddJKyHjtX0YzdpvMhxIBWqM3PxALutaAf+C3uw
GnZLQ2zdZw789A2xbgM/8bhLUromqaJtBzVHlpD0u6MxpBzoEJkZC4AQzaoE1e74
O8pAP6KQzqd/zl1FcLCHsVkqynDKpOJqiO4T2K6OTok1POnl46QjklcGOsvW+TiB
cYD9Igj8PJyYMx1C7p4IE0zMUzx25/wyH0ex0xYZ5UcGBHCAmv6KPUUoPhDx7vdA
KVb96bkRPRKMCy7GQ1z2mbZSP1oemAwNTw/stmav03vYY/uXEDQnpxkQyJURhPu+
1eaok0uBVcNUL/j2W1ktLAmURmhJJyuHUfidkGJb+RPrQF9IqF1wb7SeL+fX7M7T
xN9i4UHR92NwCZHX1XszCMIUxmkUP7E02hWaEo+vXbE8uV/xR8AlQn/bZPWcVHVo
FZoh+863m3+KoFIX4hDehYXcqQllwI46rvGV8jPCwO440CSm9dl3qtu/7BhiMJtC
qqY1J43Bca6rsGJpRkpss+nwO3CUH5pLk6TBhghJx7KMaeYfljFhNMAkOEo7j3zH
Inu+/l/fGVHj8r2hYEFCpglue8wgdDsxmpEuNjFA+ITJY9H0XD1vGKhF/Uoaiquj
euNFO2zULyTCl7lqIr1MLYLlU4oSLaAsUhAvbqeg5PVPL5no6lXMc40YBF4qHKNi
8fzrAPTS2zYX613SpngxH3T3HmxRHVrxOl1k/bzcjv7jaLClcPfVsi4JRuEr2RsS
6mV6WUhz8PhRkFGHl6I5ye3XF5hXUGTvqMsZzsKWJ1VRoisZ55zR+5ITpkViNGua
RFcdjA6VGLix2thpwbqLZ9ksMUo0tzBEnszbXRlKer7nxijXjDXnIzpGPQvPFKFF
PIAVlSKicK5qG0TgAIxdBfHmmTWqn0l8Wa25Mofldu2mOWOxA0elEF6rAToEDw2e
GkySlAgTX1GDql4zv+wGY9TcZ4YLrYRjW8bL6KULClMwJPvN7D3KplcqhxG+wOgA
f+HLNDFKCHErg+rA9tf/4QCb6FkfP/ow7svBuDaVtQU6Hhwitxo8L9Q32uCXQz/O
uXOKbGnjGovEVt27jMci/Y4Y5CwBoq+V42YqVvbXQVLHIkkLotnB4RV6xiul3nxT
2TrvC2b14AVeDTrU0qwpY2GX8/4UmI4VelBKPc53EFp0bDEMKpMMCR5ebTRqJ7Ao
piWIRIV1F/OgmNs/FfDWflvY/7hVg5KzZUcz3y1G190=
`protect END_PROTECTED
