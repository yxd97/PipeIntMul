`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqavNF5aoSFS/kWq38hsWav7K2zIt48It7KLdNvFWfbcQo4V9WQcCrEvEXW8BWBn
J0pBN/2JZCCMy6R3JKZPeaKJcH384FxxhEIPt5wJLemyOXLFEJHRHcsjeTxZVcSX
4ldUiXsnSW9vB9nE/Ty8e0wZi3IJ3PrUrr2bxJHxUauOQYF4DUHeA+amYnsgJ5jr
RmsJZiru2YGrpvkPQqF60mx4uOejlqUkmfzJXE+C+TAy0ARe4kjLXWGLT+uSTmVw
rCdK4s3x6HUu6euAkdawxZ9fDGDthKygVKrjlSrf9kcg4kqfCN2nLZoUl+AtHlnl
JhvugwDvCKTW/vnG6xaV+ZvHrXdmeFLYVgZtsxmIOug+kCENEg8vdZ9xLULZ5Er5
X2YeeyQGwEBoaYbNMnituKURTT+MHLSrRMotP/W1b5LBk7lSx33ibP/QlXaf4zYu
flFDkPwXIh8AXRWhj7Lrp6SzuYQgv27kNnJ3TP5LemAL755gCaF+VYCa3U9gzt9a
ccv0WkA03lWBiEEJmdjIAdgNXnQubTZa91oAAfY2eYKAVw7ApEgeIIZz1C5wRKfV
Km7ToHsPrgSP///wWR9dMiDsyFZHyLq853jpRz4UTtt6jRxHQUkJCI2u77BTC7BU
4uCJRwO422ydb5MASC/BqfCOTMNTJ8xeVbpneThR+Wm1+HszgLniJGgB1zLFGBf6
0UDWJu0XjZXKnjYzIjT7Z2eYc6QDa3JAcrmXUhPMOO2vh4+n+LdJwzMhNp6M8EeG
rAeC+jYDnAtVGc9EZGtezw==
`protect END_PROTECTED
