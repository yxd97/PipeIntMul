`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twMRMozV7X5x+2en3NEmUCuyd5AF7og7J5Q/dq8kGUVI+P9+CN3NNA5baFU9DDUS
w1uhpEjYi5d1t1KrceiL/E+zboEzXMlsI/DgB9uxz66BpOdcpKPvS3vnVyRVYMuy
zclhvMRUGVFR/Yo071Jmcl8XDBMfGhnlwV3CLxfzqub9J39Py0oY033gV3TJcwjX
ODJg69tgMlrhoWUEPA9H1nxfdJ2udCp4TS/gqfwisdyoRQbgOiiT8y77sj6DNv3e
j+lU1hDAr5jxZJ104VJf9RuKC2ProB2bejw7PJKgJgtLuX99OZSiSCAlaF+uCuG2
bipph8Oxx1OH4Y4fdwsCIHkypD1TgVdz+sbUJK+yWRx09ygILrNLHo2/0WfSvAzh
cbyW3s0Px5wHshYvDOL50XwCtIfIFu0CvOGbF/GV1MPt6gmCfDnWcgBSNMfdyeCd
iSBK7klJDlCGnOl0xEaUcIb5w3L0U9j6UHVMuZTvofSm1IHwK6FL2y+BjCFOVV+S
zu3EnJ/J3ll+umE9+Tr85pD4UMcLqvP6kICApgIXGhmsJQJ66TKncSXETAtC/Qj0
c6YRpKQ4PWInhprybwVvAMrRC1KHkm+NnhWEgn2yJDs5g3OqDC8mmUizLBcI42Qh
OaaMmCTkwrQye3SWKpZ8mCKNGMMEVuoprkwMwPbzeBuuAZQmZnyr6ggwoHGPJYXI
1Ct+E7Owu5gWX3xjebv1VK269Z3atYxg398J5iVu+9hRO688ej/m9w/p9CbPZw1b
te8HXU7tLQXT5OPNWyROEqgNP7P7Xpgdf1BeNqwoN9FtWZ+9XTGHNWqSqaxalxYM
NUU7dYtCCs9OtoHrJ2xDmYzm52xthKhiDOprF1P+yEs5ysLdb8VcqZljqVjEEcsX
0KB2u6o4QZ5XvBZ6TfS1VhD7V9inP5yfDXB/IqGLn8u02zzd8jFJBi2AHWupyjnk
`protect END_PROTECTED
