`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SE5MZq3Hlteqtmz5IniObIJvXDSX744WFloXQHyuNSxOSsiYcV6XNRyGRQ3QDVxS
E0vAzpIIheeiIRe56+gTnhiZGto3IyjhD1CnaTiMADHJ+48b3TvqDf1VQ7ilHFJe
1DIcfyg6u/jQDlMg929+fvsg3TQYhiw41UqEHrb0RN1/QK0wAbGfp5mODhoHlV75
8GypvvaT0f0ctCTPD3+GXz7Gx3Esurfh2cUfpjPSz1GL0GN1WXkBenmZTfyI+Y0q
E4qfvzCyzhgD3IzixZgj97IvoAYhrzWDwDEbk/Y2j1UzDkhy3yYy64tXFOs/ua8X
mYOimenq17lZF2beBV8F5g073kDRJ+T3796BzBtk0pLv9AW/MWEsyLfptqOP8THv
RB484RwNinzAv51emQD3H8PP5NgWqsukqchhDuTPDgw=
`protect END_PROTECTED
