`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EIgE48cNLcl8547dlm+/hfCyOUpXthuJ0uPfztXp6Xs4FwU4/v1o1gg5iiArib9a
kRLyjMoHCdg/6I8knsFbnAsVTpUExUbgdUAQGxEDoOc+VYzxdmLegt2Wp6db9GJf
8UFrmoFYl+q9cK7Mu/TOnmM1RxSOEEtd8i2GlF/FWaS5FqB1oEBdqOVaOBD+N0EU
+/rhVmba1aMbQwP3dedslRCLU5Z7ecn6/5bBYKcsofz4WSK5SpT4QqKZAi+MTGBo
tOY5krRz+gbF3ve9LbuxZhzvwP8+qoQt93cj942GqjhfZzpfhcPXwWh6WUI0LHyp
m4jjJIaOFpDvGlKTMF5VBzWpouEjMAB+Q9KL3PrDZoJumarsM7pYv6jCnYBa0LDe
9lre3MI2RGjcprHGHXoR/jqglg9w6q/49g5w7HxlsaffukB5OPFRinySffa+z/jc
WiBBRHDUGLyLxwTfe1Tiu1nZ2TCGTgKp/9fb971+/BpS+sZu9o7njkn1LuzAfg0J
0dFuzo6nGGIImWk4HxJj9TabeUgsML1BVrRbDochxIccwjFSjiPh8IoaxkAB0dVM
/uNR4m+oReVkmOlrqnqAd16717cwmqE2oNUSR8S/S6LDBHImxrXuOJ7R2sclpw2M
+nFhRUzJZ/DlNHYYmVjIxT4ww2puL6m8HrXgKxtoin3qecD9DVVZPoGA4EKHwQUo
EJRl6gJYut7+de9gC8z1psqx2IfajguIRtoxHTukdC2EIPONJerI8DQ6z6o5Obn4
RLPE87DpTosav70YA/pz3M9q01TvKZWhvm5Q9v3YFa4wc4qVPv7LN/L3wZ2bL+xI
eu3a9WCAWumYpcbpnw7LG4i6RPLE1ccx0xYv/EOQTUX+cw2KNvrF6Qo1gkid2hc2
SSbhDzw4l+2c7LD18KGj1AEN6xuZ1qHk8VCD5ePlnv7xNhSWlMdjRtEiU1lhevJk
g8j+8NKHStm2UcFStowclvxpSnrgSHoJEdC0lsuCG0ySeO+Hh6G9bYRh7hz+ik3B
pajNg0e/pSIj1fLiL36dAzHRRhzDaMsIMRZ06OWyeAV0n84UncWHVf1Pg1RA2oZS
aXKMSWA1ityLPV2WyL0DSLt+bdE7ikZ5xdC+Itsp9so2UL2jOdJrfwAe7MP1DSQN
mNaqScEiOTsNW0X9oGfmz4X+o1Hes2VWn4YgFQ5JjY0=
`protect END_PROTECTED
