`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2luE4kwp3HADXoEsMMUbQqDVsLOcw3fuijU2v0Ix+UyPV+4Yn7AT41ldv1f9Qmp
veWX/sT1LFvNWdOF7yALaeub36HhfBFSllakX4dc8U7C3/xlWuq6f3tZYna3d+E8
72obKYSZ0CZOgHwzHAEcuX4JEgVV/aLgY1kgxSLdtBI+RHxlnag1gyIqLcP9SrIz
arDNjAVKmfkXVaCJchwMK25Ku+WNYpYYRpNBrAwsgL9qPTmYrw8CxsZ72nZEJjvh
`protect END_PROTECTED
