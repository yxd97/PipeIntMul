`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LoA30tdWSgWmLVTlSkVVWrFIk6FbLFesC4HJ6aHT7LI9tQ0K4C0kf8YxA99SfXSm
vzeUyJ1BG0sb4ADONCT8deZN0FW5C/STmKT45w49wcASjU6IoLYCuACZSRfZ13CQ
sX2g3AAcjAgoWDCWVxjKRP5P95scB655mIXoRVgVSo2Rj0t9Fg2SpeqJ3J97q9Ve
5vRQTE9glwuWUser7wa5SuiPKJAVSJ1f3XALOgRviIGK7OmlCR+0WY/no0mBnAkX
DQa8bdHuKPL2VSeh/bj1QSO5PoVb09lr+VEfD2iXd3O1nkPf9ryC9mfsr7a4zqRn
u5ntIbiRbHjQ0HHsJLm6dqvBdQZKo7U6EsnxGlKJBhv2AjoRqW/LS0zkqBLejT8Q
ptMOcWitVPJkKbFVxI8aTreBfWQa7WV2PxBnh9Uc0Vc=
`protect END_PROTECTED
