`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kpNYu/Br87pO6wi9D1VrciIo4ly//mRDM5v+NL0wv8fFx0l1IsltHy0QPN9e1Nb
vQATca3/CebJ35fzrsPgQTmAPNoPxIMTOK2GVszsu2RfRI64QuplofVukany1qLk
wfzj4O+5QdopfKzO8AxDBYKxl2ykIAw+APENhFlkL+BfMp737cRi6v302tjasqHE
+ox2jVc0K5Hr7USwXhCEigY5UchbMWb/Ic9wqx9sEuPQbMA4kIAHnGppcz633KVa
C9ed+2cqohjUyWptkzbkakhH4rOrZcV04O+Ow6czKnVsmjka7WUhFFdJ2+itJ0V2
2RmHM3bQAsBLfWZgeNAlgiTBmL5YMZqsoWxuYc/3ZMtJwTCxBRmzfhwyPCtS2sqM
PdyUDz1UT5ojOMA7edgDVw==
`protect END_PROTECTED
