`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6y/q9qo+vDi8qZtyj8XoyfUFPygq/Rzfy8Tr8voXFaB9FUzteOhRUagkhgDrJze/
V7ZtBDdyJgBpCPujDQI6+iL/ps8EtBRUHCbpSwdlNT9qYiroLiFUDCP1a4cfFC/e
uwerBHQulImx4AhvMAmXx9lYDBj5SuP8pvtqnn7ZrYgyA1knq3a6S5pzUjpeSJaq
BUPcZuoFUSrShKONRNVmfvGYs/CpWQgj6sEDTUClGUvHKb/IOhjVO7M4c8bF29fN
`protect END_PROTECTED
