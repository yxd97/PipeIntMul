`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KnQq4ZP5qaSlfN0FWkCcaReElIJvtnO6nvdjhhnjdijp31NOZSC8wUcFF3Wmf23X
BtYURM4Sl0RuRaILbfUcJe3eWZGJsOb+69H80KvPDHJ4zgWcHy9N4vnfSZPRtL+1
GnjBzfooBKg8+24OzYgFOKTz0ky8dTy+978OiDHF9Z7qkEmaYsJ3oggTIDUVvPK0
lA97D7eVohXmnOeUranL4yLUU0yiuVKJXVbxTTlDbqBM8GxvMhZOJWCI/jsMkrvo
BKHAsOJeHiWweu1Mj8qVsX0sfASnSqehALPm0Ph3TNgfepKpK7GBqd5E827nWBNm
h7n2rMzwwnXZNktGEUL4uzcftw7FH/FeGv7KBH0EPj6cnfWS5Xb+W4l1tGQyvxyB
4ztmVgKrzRxjtajo+DhpsS+nThVnLWYLG/XCJjqxMEdXIjbvZeMAaVhfIzePCmrL
mstDP7+0wiE1NYUlg3Z1zeNWBe+zKsVSBprJ1EMCMRa0v0KbpvVYTIC4hiRH3/cb
C6zdu+CBuLSk7+dSBdaqnUzrDN3eZX+rx0xbgZfmQMU=
`protect END_PROTECTED
