`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LFtRpn/KNynyxbLoNCxUWUb3nE6udNPMwtg8F6F69/C1B+U2kT3fc4wv91HGeB/W
JT+QAgxhQVnkLvW1j+/dz7p/ItdjMdK/pLLI8eNHyHkCeXo9bozgid7UK4wcecTD
uIUpBnKZ9I8c4lx9G+SCb0oK8G+U+ngRaybXDsqmbPAz77PRBTdHU66E7zaZ9zvd
3WmQ6Yhi6GyHwq1lL26pSZ2fzICe9VNzoXb4/kOu8BqyMlxqHnS8/UiTSfsIh/fO
4T90yn2/zxqk7A4AmBvBq55Ay8II+JMs7zR4ONov0U6yg3g8GTbjfCRWADs3BMdP
Ypay3h/p8hW/w2/YgGgG1XGZhKmlQmsVUxrB0I0LKdDi+1EWyFUEYIxwn7qixWcb
ikgOJK8AESt5gjnw0AstBQ==
`protect END_PROTECTED
