`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wMULeNKvkF3sVBzytDXUy/wD+v2zSfEZCj7ugw9/MdxYwaUsHApiPGObN5EaUykw
frMUq3FeyRz7uqB7UAf8EiuNTcTDXHVEXLrFW+tWbj6rI2xqPUoMq5i6LLvTHu94
V1puZv+mXSWagcHNjx8eKTmQr3L9538ZJbODe6N8zTWRm5revvbyXoUnjFmJ57Wu
2ve4WkFoE8qh5o3ZGp7M5GOrl5uLeTgwMoP2uzYnu2rHmSTEsZq8EteIt6VJNN97
KOTEqQ3+dg4Zq2uvpkx1BbTnuBak77bFyIHHYw9ZF8k83h2lWZKI+sk2uOL55REy
ZcRGS9EmrT6m1n6F3g8WqD5DjVorGIv8sfL9/MQDV1PcOvSdETx9CIl9KwbXg+nW
UasbD8dk++vB7VFGbUQBdXG/t7EYO9ACfV6qilto01VlA6mojdfLCuzKNq8lVYR1
Dv16ZgN1/6WC+dPLI54yA8c2EZf/+0Hmh0MhsJbrpW3NngwfDBQS4spKxE3LNx+U
TX+MYUfYflauZ521UR615RpZavNiW0B/ks17Rn/fBwcEaCILkGTsJhkDhGnpCLh6
gx3wPagWPeze9Z+F3Mjpkaf9d1wsmT8Euq3wadaEr2QqEQf4NFwrhUsiNkxaelZr
Xl38hho9ayqNO0+YT2A6hBHymiR+82SLBfFzgOOhVUNng6dEF5FexkUbFbAKnYhy
7r3dOkyuZNpFClOU00b6TKVqaSWv+RPyq3CjV5sd4mAuTPCQwi08rw/1Rctc3p1x
4iiVwJEXZoTbsCNS8DjOy62M0SeFtaiTlJLqqAz/356xlFuMNWvAoV/oH4Nz74Jt
amDimozbO5hmgH2JrLEAavvFc5/dz85l37EYoepoY+8AF7eNjknwy3GVwZgmTP2A
BJIBwHuG3i94/X7qYLcajzZ/VC8/+ItJjN7tXAf3pCJOLryiaMZ1FH+IwwkiG7wk
IdBBALNaPQWTrHUMsKCSKUwnxdFcIC6RKc66NBfyLOP31wpQbXJp+diLIQlTy8pq
EGRsnnK9pevtJuboPfupPeKPMgahaZ5YslzPuvzFsLVhP1Y1n1i3ppSmMZHU+Vqr
CdVOOXPQ8SF/bVQDM2LME9fpNSNFS3NLpszlyHNXyIEq9KSVRRWOKByAYQ2FEImz
v1sNsGI9lP86nx7MBfX1tcZfN5NfZU9QqJA/O+4K673vKFVfF9plGU7XXY4YWqI8
ESYe5V+4o7NOR8cl3dB4xUmr73jAMEOuWGWvEi/7Q9E009fAAygYiQ815f4WDoqS
DA9+p/tef8/ptSwHwwuvRtYN1fiNSkYDgLXQL6GUaYIA1UBaLVYLyYKb7PVoN9Pm
V5J/FpfQhj0aiZ07u2Orcg==
`protect END_PROTECTED
