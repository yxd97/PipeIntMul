`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m9/ct75+hzfwjIBmHDPUKmG3WYnDDM9x/Whe4Gc2tVZd9E/5X4mYsz99VO1xMluj
GjGzmB88ydby1hfIQJihJjCglflFCuoxZfQQxbtFHLBWwipZMc7AW+c6eHNFeBmv
HIwMQqQ2M+YHS2bwteKWkuscoA4f11P9m+/Gd0XeX+8KtQ1GicY7C6BrbupGQ6CF
HKkkDJTtrdD39tk8iH1o7Vc9QjIqK7Jm/qd7hC5wgtSWy+pmdm6kzVjXGrAtTrUH
SoBp2fenDvJ7IxADDkznFw==
`protect END_PROTECTED
