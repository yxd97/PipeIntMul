`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6t9CXnEgqYjnt1NT3Db7N5EYufq1pD1yCzZGAtl6baQJ9MTbOGpDERV9af0Q18kt
ygeMNuCKd/o255+s/T24HqThb8Fo//FvWYcTJ5YaBm+HfzeH89cCJhXU/LIO7nUv
6NVp90ohMyrAlK880UgEKpkx0GqYHQ637ZYMq0al8vYxq2BNO/ZldWKa8PitJ8yl
74omRuHQO6xacPx7H0JMCPPa/zdFKcVuvI2+jEuenDJpuU/3P4oA15lWDcImNMPw
3YFjju5/sK0c/jt+Pp/MlGJqSk3UffolLm1TgJUTWffG5lN4plWTkrGYLBwIw7mK
or2u8Cod8BeeAzupbJU13SQmxrpuHxNikKmlRyJRLM9FFTFM/1fXNiZHQtD9COS5
prq66WmEhee+AVX864D3UbxbGinZuEnPU61Zspj1Mc/5GLqxbX7GaWKsvdj6K6wy
vVju0qbx9Dbmd+itpovj97dNpBhJFGrDFk5KvGTN6aWU2J+I5EC3FGnndQtspbXa
`protect END_PROTECTED
