`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2CCTMUbgVHDPkAlRGBwUjeGW3oMQjjOy7thCYO2L0rkRuPwtaIje7x3cJDmHvxfS
paLWeXW040IysdrhPK8Nf2ZdAoLEs1XlDGVltSkLwSDsfMnlSo9oj6juFP8cTePv
2msiaxE4LyNGjAbKfHlWlw+WpaxtaB8CqjpfWscMRUm0o4WYRVnH2joQ1ko5Cjf+
JqrNpK9csEWDb8AK/sVAAsApIl5pjh63/rgMHoUuydmt0+wn/FrxNXMF7lm13Akd
zC0SRODkQKOzNnYKFya2kVQMzoVD34QZ0jAwWLIe6MPGHtlX/1z5Z+RYxYVJYfXy
1scJqc9zOAJ7Q++Ni/AXqImzEhUGIhzkmt+lsyD+cWoJJA5jg4eNyPWjwqFguSHc
EdqidRpApGELUJTgih6MBQ==
`protect END_PROTECTED
