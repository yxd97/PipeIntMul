`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KP/TdjYvi1LJD3kJqcidwg9q7OBOKyD3Vx76rCyHeKDPhc0L++AHA/yyuqhYFIFO
+nVEK5D3rleBPeeIxOnfcmnvIapbfJbF3ae5cvFKFAW0l+Il0FqBKD4cBDY4y9NQ
b4RqAmiuskhAjuvjC6UIdnaOxmQg55U9TYualq9eLNNTcMea4cTI6G3XK8hUgbd3
6zhvkgeOvYJ5nsDwKWINPVXwVmwhUqRAkWRyFd88bEtGCY/sefHYcz+pB+Ik+cFt
70C3t+FvJ77NJw3VhETKAWPNaK8SFp9B4FU5t3jJgcHRnW7/oeDdPFVgi2IGQJIa
Gud819AQQX7ZcrHkg7XMeIoEBoEOGMPRq3sdAp3hokkFk7MSa0zbkcbKel7TzNvX
t1P1q+SV/vow04kaKdwuPPAFOmTkOprIhff8qPlDoPxtOKa0z8R5MJkY/jPs4DRQ
FGrJaxVHvvnfEWYYk4njktOq6F+Ou5uajIqcfhYgj8ibcwm5LDG9M+ULpfnnm53i
6EQS+pQ2o7DkddCYlu6WglWODnNB7HARoDZlEo4ZlEKv7GcptJZob6jVmzrRCJD0
CHB9Cshpt71O6h/kHhgYQxs3Nyyfw8DG8/4eKQIJPE0ZcQVthN+5nnvfcQ4uQZi+
7IMBlMGA8xjoQSXgMJDvE9OtrEGxMEZR0TBG0nrZqb4y1yxW2+9b3Y4oiw0rrpMe
PSMIj0LXDqVDVzCmezuRgb30v9Mco2pDlqk8pawdUBZvwRqis+oySBupb+CZXsmf
IqyoH4B+ONaWmvsEnKRtsQrfD51silIZaHvELF7nA38=
`protect END_PROTECTED
