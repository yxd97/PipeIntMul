`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8mJ0Fcra1D7UoD6AEuMU29k63pgh/rRE//fIlcbZPR2aIVVzVQbOS19noPcoHS6
TlpfzGUuTLI0igJlDuEoSVo8/uT1K+mCO6vf8ja3nJkgaEjWaIvrrM1SI+inb8UY
5/wuXRFO1iQB+CwLDtA9XY0XWy6wd5nVPAiuVL2SCCqpxanGgplniL8MK9RqYO4E
w3d1uiL2/hHOBrIsTf9MzuS9CwNX0i5AE0kfaDv7TmkVS/VC9O3d4Di441WocjDN
FRc9zIoRxVGbrhCUzbmCkLhL55k5x0CKA4FxHhIcfIKLbj+QoSHMgDpOoLQ1vFdY
Kw5vjywpcPIzRMM1AP9zNw==
`protect END_PROTECTED
