`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NH+2V3ocH7mrgP8uPjhmEestojzZ47tc5vjnaxco6krOthb77Sdzy9UviM46MHWt
nPJBnXoSTibYEea4Z42nevZoBA+5jhsy7HHDc1mKwJJ57JajF6ouMxtnaOz8I/Pt
wYhCoIwIIfkhr3aVoZCKfU20XXqtYTP7aDr0in0HDFMR2UIMQhh7tjI7m/U3RAtk
qfw+jQapCuy8W///TY2QUY4fDOyd8SzK4oy2UyoyLHKz9QWUNR1Sr4RzeiuRvc6l
kQ319iylipocDthaL7ORI0tLH8j699z2142ZLkO0aMNa9jsQq7O3Hl2eFZ/lnbuO
+mXBDygeXcLPdNzhKOWSjhuRxYguGB3AYp+EQwWX0UvKKQ0WiSSWWuprQk6FzASI
9Gu3jPQOjXHKwR2XGLP67rAiOlb1fYmz9aBHg67meuw=
`protect END_PROTECTED
