`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Js3r/pgtpOx6B+nvyMKLb6v01lB6UqpSDV1gVSpTOK+kqXBz3uvuw90KwL1O/WgZ
S7WuCL9/Hl5zcrONct67uL7RIXFhoG8TyOO7J5DOFsyMhHZ06ipC8F8AbizheCAd
EzS35k4sjXgYRhlBcJRkukmrLcyknUl1qz/IuCg56FkvzkhsHH/8KU2D03dZFE5K
Nzken7hhUkh32C0ZF8bI2aw5MKlSZ4n3sb6eMZcvxzCMZiA6G5tmdR/A4hzXXZiZ
niDK5ez3f2gu+aS6yz2Q4EaOkZPo4kglmHVWZPjhgoT5RkQDeJ+c7kPGca6S4AnP
cCb++phFUNOM3OLIhfLctIqNdY75/p82obaa4a+uOn6OG6H3VRxaWF1buvJbuLcS
Qjd7ERdNECYvQ9IqhmDp7B4h3ULFFvZS1CDF6+ml3PYgfAXWwbcdwgEeD+uF0spL
yXcxh0EQFhEl7D3y5714jLdDUh4p+L0+XgCD/5qHlrmLB9X7luF1pCZXhSe687Av
scuaaB3XDa8IVzkf/MDLBKkeIW0zKi0x1XenvmLvzaKp8wK38t/r4DTUoGeyEPM9
KHooUo2bgq8Daky/fvBlzwldLRInHzOtyMYaFLlXIqrXVvlHh9uHf5deIKQxqa5R
lW6qEooipjS40LTSuAZW7GghobbMAyY2xcvsu9Vud+UzKbTCqKpnhpJ4zSgWMrn9
vkfI4Q+Qcg60dC0X0uEnYlhPBottY8D0fBqaUceAnOKr6h2WNsDY8BdHLBmGjbTx
WI1/JtHQMV1EfsZ+97u3Q3V2r0YJKN1kEFi2fVYcHTRa32Wgdl4hW+hNpBlNa65L
sj7ySxJFB6Oo0yL2SpA2ztk78EkqjGr+doPoDyoZXDLOGcDrZf7LcIoPU2cdkx5q
0XLID9Ub23qFy0uViQ2VzUAdsMr9Dxej+g6AEagLZI8jXN2i3CqcH2WPspkOW5i5
UsT0u2tdPkGDTESntLZn5RRVeHuXBRh+HUxcP3SYMMGK4LkDpsDztm1apPcZ3Ivs
JUuenlKgznZ88IFeood8TZgdlU1XcoRs57S11seYtZYNlonDJirSfMa+/li12oqJ
HsB0o9uIw8V62LJRqJO232M2gJPY9KedTDJ9IXJD9ILS/t02kx+PVBOT23bQpdzS
48q3JoctZt1k68xENDOVctjWJYdqRX5pATVYFc0sQyuKWpygX6JXH/wlteflFOsu
kCyL7Ac4324GaExq79c8g2kGkslkGm50y+zsL1sb5vfe3XNAGYAzlx+6TpdKPUvd
gLbITbf/ZnfTV5xE0lK1wbnXU1Yl89SmSs9e7bai1An4UoVG3crs2e7Rc6NGeq3f
Un92Ix4WcTAdhDJLOZDota9bW0esRxclFKBrj0z7eNyXngicmwoafXZcK+1ReQan
1bLDhzzxq3sdHiCc1jtuO5OT2KakYtGS/XDo3Jd/8xLcSL9rgux4m5bE+15n8HiD
WxLV4vnpH9AFClleGCdfW6Hv3NQWRZezDn5MRVWiALCM5DwHbBeQKQluAQLd4nEF
XJMQByPNsGPZ3AlyGVPOD+hf6DkEUHOnSuOBEYJuFH+6WQ44/Tzj7zxYR8lSE9N7
VK5wC0jzqmMqZqH/W00qIUn/GCIhxj39IUj1tjQZZkaPP6COj3rz3654LpPNkBxX
wgAVSuJeBWiHtfRSeqfrBpSEe+tQq5Y0KaNCM3QW9I5xdm+b7mo16pnLex0PKRT0
TNTmBeEfUDlMgMYNYtQWHhHVnosryr31E8LX39sZ42U4gB2lX7TZk7X37nEwTyz/
0DCCoJcIrQhUlcL/IKgkGJg+qOlPP8Bgc+n0RkYyKHNR1skbBL+DxCSjvDM3spQO
o6p2/hlD2ufNcRbx9Y2DrF8EbBZpGSy6UvRiq3p5mcXYC0wlmA5vUArfDoiGMobb
n1GmKGcCOsF5pCA9sUpZsQJuAQqlAjQAgb5QVrlGSp9kBbB3GEZ90EalrXSDykkh
cow09OuvELrnJn1gYUhaB+FSwKiGeoGCHlybQvi4qEwh0LxhOpFb9mYjF6ER5tQ8
/Ef80dHIk76wM2qxsphH2pjeXM1YCP3AdS4iN3nS5LV4S8hWpMg73u4TRYR7M76b
kFaOV8Zu1uFPFEHA4eHLf2oio+peNH/JVnsjNMl9+OsvUquWQvdENw7oUCyTxLUW
+iUfI4/8LFJUV5fcJMdn5ewd6Fb8UmXo1jkP+W9uM7AWmV70EYha3gUj/qsHApP8
gcWnUewNJX/Mou6Qv8XAVuJxie5jL32BqE61Jefn4/9mFwlJSUhsFT6Iu1vycO+C
l+kdR/S+saFEr62XEc2eVtF0QROVDW8RIOgABOEQe+KqMdgVT7bCVXnXQtSaWVyo
OuAFu4iKbdEtfKu+4blHXC4mhX2ieAg5+pA3W9Zo27B5d9j8om8aDgmpfqHXCxiU
nelICg32Nkceo368mELinyZ93cidSSzvgtjMI6E54m69GrtlTkUJV1h9PbGVvd7a
kztvr8uqE44ds1bI205KUlneDajjR6h7cEFbpQzFgNkSrXW4Q2t1CQ1wg2+wDZqn
vYPwMI0jIxj79J4tNyDTQeugyKi1tGtqa4Eq7tKXKOq4HHxG1c4VWJvYDNpzXlRS
q0WM3D7vuIFUTsbtKNJjlTSHo4Dda2PiNCbX0S1Z3eUWh0TKbIUWKfUDDRi6MZMJ
iLPxuRYWpd/kBx7GwV/f9IxZgTEuQGdu7eug3QCQen6aJqsNO15KaV+Dk6GZ3Y+o
6S+Q8p9cN3fFhO6kqqZN8wIC868sJBTp8i+JrEPTg4Lga9JiCQE0zWPqDZddjlqx
A0k5NlCUvgaSu071rmPR/jmiE4YrywG2P/VE3aIWUa5Smugsonqdds79EAhamzQy
gVHrG6mLWdNMDmepkNO6I1KvsyNf1Qru++pZp8MBEC5VPjMgGRvDZY9slun0xiE4
/6wH6FjtYt8T9mWBThnrhtgqlk3ZnlegT8LfPfdwgf7K5C0bQWH0OUYk9ZVNqbOx
7+Vzyu+hN1+x8RfKoL0xEN8MsFE18M9rOPXubRUER5b0jI+dhHOLhuibfsW3gkRV
xND96mPno+uhtfI+DjYp8cq4P707Gb1VE20qrQHuXdHO2r3jqTcfMddCXE1tDOAS
/cDLsjSF16SB1bVh3nEDZw==
`protect END_PROTECTED
