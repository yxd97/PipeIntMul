`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSuAw8O4Jqk1N+3W48KO26QSr1Trfnu9vBhLz/zsh8tR9sXQ2Q9lwtqryGKb9+aC
qgb1RRLdgly1AtF6zjUhEKDXYnRwHIZ8gvO6OITrHS6xsQtVtZNm9+P807fJBcKw
jWtDtHsLVvmtq5zd8Y+Ik2BbK5/QXYv9TJHzLdXf6czPZsAIZZqy57BYzy8++TTS
F4gFt28iL9j3DPGCXqlGfkDClqFyP4ShmSFONRepgWmXJoluf59twq2J3tnjC/TE
ZX0dgknq/z2ER+oWz+3E4yS8p5aIgdaG8e7/sHpb/Su6OVEIMa1Vu5bbwcZyPhAy
Rh5zPfmWuKZ2sfX+/PUh9KpelpdK6TF0fn4VxD5qOijkdcEIOy+LFLBAcxbGKXAw
dQdhCHfznGtWgo2aOiMUTNbB/sL27z3SfK4zaAqoMN15b6CPEU9u8xphHJh4z73E
9Z205pJ9Qrx9oATmUN9J3/2KvW30c2aDpj7WxHwj2L7Y2g2rbjpWwemWz5vwakau
iAZuRDxmpn7voznfrv4O/o8EPybPUrGCk5IFwtjF/SlsilYEbxtAQxOgkVJgQxSA
ct5MMvfeMl1BUAy6ArqOzW40/lnnRIrcP8ktsqC+VFAuW58gW2ggIgyx5PhVMAH8
dDAMJZ6JeACbibyNVeHoQlSPMkTP9sPuv+Hb9ygridGeBqh9ewPGRabMMfgX2msp
4A4PkYfs5Iq43PBItU2ka78c5vqx7xGcLCxVZjUMXffqPwDJTgjDktaRCyefjCl0
4WGX4PYN9c1gAZvyBm/utTZdY0++jvBWAeVdH/+WXA64TVvKgll6rLutkMHtIDg1
Y+OMqwfUtUuwI+KJMKh+p2fgJLO3/fBDx7NayxVT7tYxoGApA8f5oHmn2pL9Xr2Q
y6Of2gJAEhc3NG1CnulCav24c/47Upgacy8es+dWYiC0+LMprEUBE1n4H2Y9RQZI
R9wX9LBeC3GKd6Ohv6PlVF2xhSAqHwqyJOfZrMQkKq6fx8R9Jkmw2GpQR3fJxXMq
FLohnSrNeJdE0g7RhkfTiK29V03M6wLp2+dhX8J2TLMRV6roXxTaLVcLdgNDCQy8
z9s6FXk7DZ4xZPAr+gAPU0uSgZfsEWA1auCNtbB+660dh41ccWLtPvpiD5T3gCEN
`protect END_PROTECTED
