`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rblGuBIkUzejOZfueQTnfCb7+jlgDbnfUO1tANSDIxC31RmvAi3mWzHvF5oI/3M7
Ap2mM6fqV7Cmk/bJjkbKosLF7dKyT/soJEpbkt3yW6nY0oJY7fquZzthSRhAwOvt
pzb4N5ZdjLnABuA8RkYo263twWiGC6+DBct+lNB7vrKJ16tnhVbUZYOp3KByFdYO
wXI4Vt4msiR/QJmQQ4BeCNi1NrQQ9CvqFcql30vVuscdPKMeXheBTprcKm1JYR67
QA7MbP0hQSsQ4tXb2Uf2LvydmTXrDuDQx/XD5wwT3xe7QQIW5HFn++SZZlcmYLg/
Rdoy4KJ/J4FlUFXi9weuFmBAWm7jF5M0jQJnqK44jKJYaEL3+t8D4hcc1Z7k4JxO
Mdfak+Ehqv0ln0BzoxdH9DrWi2fKsX3hIPlpKSeo5yk=
`protect END_PROTECTED
