`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WCQjzdPMUZQM5m2/XU48jdLWGONk9sZS1g+2OntQHi5YMty/NwiD/iBrh5VGobG2
4QNh51XZuSiHfKzmmXAnejXhZmGgMjONok/4W5x2VuTv/w1Bk3SicBMGcR/cRPvx
O1gXLh6pHlEfkOSzsGnwyo1m/rKynDJPvnUCzK5TgNoBdA3WlpedazKfo72YCtoU
OvaXXal80B50w/0HK7lUzf6cSrnoqfdCjYMHKYgg0i1xdsO+dkOGdv180YjHGJPm
RLT6V9ID0EkSC/rvJtntBuKLd0JpsjnU6aQkisxV+Bv/NWNYza5faVGfgSw01Q7M
MPnjDf74oJEEHX84x5S43pvnWo9Cet0UgNq9i+TVBwk=
`protect END_PROTECTED
