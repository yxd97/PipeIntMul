`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AMzcgDz13SI4l6S5IPak/R+Trf2Y14QIQVNbrykMgDdDJVAqijMzr4deIIbFPyr+
0Ro/RtXwg16eiBn7Wy5A5WvtyrY60IWHFflbai4EHzFzIXy8vBYSPEsbscMOqAim
u2/UNbP9H/j6JRN/0iQslUVFeqK+xBIidAbm/3xEtZtnSu08xrlF8Csddg/7zVF9
v1AAh2hYKIEnlqkWdFspjiJrZUcIAT4mDGBBhH/4HgFRuBH5URjy9SXAE/BnedU5
5W2xhny1U4oq2mO65pijCuqEw6MH/ef8Ika2vuq4AVpt+hlO39fHt1/a9QbPsZsV
/gBjE32sVuoUuCFyTSfAMw==
`protect END_PROTECTED
