`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bqoiY5M+eEouKz651TmWCSqXFDvetgFSfuPRMUL12BQoJhRY3b0kz6ugxNobn49l
AsOxzNnFSVX+yupqu6/INAM+4hGcuDxxYf0s98v1YWsNNBxbqWXcwYx9M/nnb8tl
cZmHU4Cy0wWkpcDhuu7i/fHDbZq6JvwFvl2DUx77hrio0H/3SfvTVdgyPX6i/gxV
QWBG6Nxnl3zhZQ8crvvJ4MgQ29WUXBd5LRMtgedG56DdBaOOz7sqOZb99jzoFAac
uW57fpt+q0H2Cz5UeP911lFnqhD1MIFUyMC3Q/wQla+6qS+KUYGuvm3Wz2nZSuZ8
Ho23qkU4p3wq4Ad+xDfYrqNsvXuzM/c3yMmn1I4PSYr5ROMt+CM+FWrDatAoqS57
xdwjtu+x/q9Hu/mHXwBY6kuFMXsUYCx3VQX6IuFjZMh9+PkmvG+zvl/DSBdZY+Sf
gosvsNkNZwygUGPsNBgxDBYgH2gPbnM+OCB4tq/O1YpPq1FB8vewbC9laSuz9wlL
YsWxomhyltbtHoNyZ+4httnGXPaaQ/3AG7+i/Z322dkgkRoMYFDVm7lep+kDbRtr
D2ah0+K00qvbwFPebJa9blBks78ga+VgXxC/wttA4BR2ebxxmBt77YSfCDSuMpPs
r4ePC/+nVSxPxZBp/S/xGEjc2Gk5dHW49ZNob1uoKnejqHAalOPpj5pp5FE/9/C6
lXdfJXiEt1h0r/ATIkyGzzSlKbzK++wCO5VglMuSOhqsqem81iuKRsP4Tihjw7xj
uADdPXsvihQ14g6t0ucpwmXUAxhww24sAsOsiPiFSFETSY9gQP3q6LP1hxAKuymM
YbrQyTJ8R8Yu0b7H0SGUgabGJCjYTR2c0qZ2i/+4cMY=
`protect END_PROTECTED
