`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LBP7hpp9fivmX9MyF4pwRq1BA9DjbN0Q3g+e/8XGRW8ZMP8mM6leDgWbSQaw2GoP
6VuWsAXS4fq9+WfSSv/CzoLvEKgWNbquLzIuC4jSR3q66vGvycM4FyG/fGDH4aWI
kDc3RdMm2lA+TUVRcVu+i2KZ3bZXpxwCwEq22d6+WY/2RwddldSgw84r4bv7arFg
q8jr7Ti0++3HTWKit9EUJiq6/NG1hOc3jrbFb5NcntlLoMol/DbbSYJTjZ/xKhlQ
xmpPH09f5pPxvpzZOEG8xw==
`protect END_PROTECTED
