`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIuOkwSqPYdw1U184wwKhMPmAZHa9TZzlmEZMbG2SkgM7U1o2vSib0wbHIACdwSp
td3M88WiMgnLpoc2g1ZHJOvzttbtQZ4KefRc/nPFXztijzSPcVfwbhgON6QiIRp9
2ANH5u/pXZ6a7Uuk/hDMmEVk7cJ7FTM/9WCXlsa4u2sdNF3yJ7v8sB7AEq47/q9/
w6ewDVg76Vn9MivPvBlBgGpL7TmV2yYamAR8j96qV2LTDmNEE+lNGtk9OOFHQxZJ
EhJw4jCcuMTICV1tV61lvG7EAHfaq2RLfX+wcYyk1SdxhFQO/nR6ujq0gjtouI43
wGOcUb6dCH83pEBVa/doH/4FPsabkZYK6wtAm5LTa2H2f42NPgi8uzVP+ymVdDYz
60CLqJLIUXFJHLBiyAoUcD7Q/M6OnK/H/rxq8FAU/Ug=
`protect END_PROTECTED
