`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjgSg5gjNyp0opcMaNs2MjYQ+d1AGzto7amWxh57a3OBBk1KriAlgWRS490tWYcJ
5VfbBaT8k8XnVXeSbfY2Q0AN12LnnHP8bnj1xJqDzriFZ/4+inRLJ9DD/GFru7tO
W/ZvLXjHpLvN9AT0GkfE1SC95fujSCet3pPXpUSmxAjQ/qwINmclGVkIElCLp8zz
HvM7GCS43HKLPzW0jSJ9Uf40QdOnW+g0NjxOm95aHn3QpyUXuehv6ySPEJnchDQT
/n7FpAI7uQHgCM9yrlJq/JSvZJrTE4VtTrkdt332cFqzrpREuHFz9bYnYsNk5wAO
upcUCw7KPemZRXdyKqSiJ3BRn1WxldwjWkCmC3Ejpv2ybrtC1S++gKGrUEsukO/7
lu0OBXrmViYuRpEFo4OKwuIUluH30JrmDRbyujV8ESQQlUXhHhgBCco4rQm6ZYlh
hVpayMC/orIQOv4XphPbrJumW/URb3DPEXMlj4Yj8IGLVCzut1ybLHi8rPNOiS7j
ouH2B7V8pl5NCZTPQaiFbpYccKhjZFDIDpEvvh4qufptGEj6xlFf3sccTGt9JNnv
HsftYgoel+27aq5tdhrWpTQDtAJgHP/0GGyJEaMOf+kacjdS+majoOSECv+qGCtA
DaRW2HWyebu6YW1K8eVzl3IP8aA6tGM5kQWlwrE5TSTtlLWksXdiOtI3rfPIr6nG
xWsS8aY/iwPmtzIPAQlZojr61eCe3rHCMESiISNNsOuULOmGSf1JnKFu+T2vhIKv
XejRgPVaSw+d7t47SaZo9wm/o+lZjDoJo2dLrxWjL7ycAaS+q6/fyiYw6LP2Ti1P
WFLdy9NKbA6JOEPyVUgf3JRw8ydQJlwuLsiTzANRXfpUKijzwrxmm8z7jAvd+jWh
M79GOzZGEB7BBtEzmn8RN98SM4TUeOPL6v+M+KsYlzj2m3HFnVodWfE1wctTJbxQ
n5ofR+oB4xgD9ZSgdp9CvWYMTL6fsNqAqPhUoawPr4QxKKO+3Nma8o9UnNa9CHsF
B2hTUYU3gM3Mlwr23bzC0U89gJ3jTzkCkuuwpheVKEvTzWJ6vO0tARCXfxnm2J9k
gGBiVky1OGe4UkpD/e1gUypC0zLQOfj9eufnO4NDB4UnvF6aeoJGyHEUDrOpYz42
4pYukyq7zt/Y1gdSwohceOdkM364c5yrL2QuhkjkuOrGEC3wklBmvU994fX0J/oR
yPSBTdgpjB+WW5lG+9E9zA==
`protect END_PROTECTED
