`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Os/VMKq0zVI0kGwTwO2U7l2m5X/Vt45CWB2xYLZywFaZJrwYwt12SCvOMUdZSOg
QyXsmMt916Ce4bllS353ftKk3hX3CTwNyqdLUpok0a82sxRMbGlVauhVCaId4UW7
+y0Y/1Ep+8Hrb3wFz/uFb0MBuOLuVM5CG+xVHJxdDA1fTyEpIuif5H+3ZEUgGfG3
Z60I9Uelo7TqOeNkl6pGLYHz4fIFoXVWK2VXeVTr1EKek/bZ8nnIfaGvK8Bk0tpt
Jw6E4yI9TbL9sr2Y1C6uwQoNvIyNxaVxDVrGak8NsE9QvW9qCzmh/UG5wla+rs4h
RJ3SilG0pHB//fb9faFTyABr1n1Ml9t2AgYLJHBKduiWeOHkpXv+Uop4b9ixJBfB
F0ZpPqC4z2HVC7dTbCZq+Yr2mXVKh7RO7RVst8N+X65ZObfcpD1aLPXNir7tfkAN
1m8Z0qBpKGI24BT/GPn8uPvVeKOxYuPSQbtAtpAx+wrrGE58sCUNwlg0UNnSr7Cc
4rp9sXaTgTdlG5i5A/ipwpJEtv9Gt5L44t1n4tmTQGrJQa6pMhidumPqolt/G1H0
`protect END_PROTECTED
