`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5n7yPqXbrhwPpT+dgAFR9m7FMnf3DXxd4Stvvr4sFgOhMPmQBUwwhmUl79FV8vzd
IExrn7hpy2X/QgFOvh4+gZCoI/Ij+M63n6CF2HGs7hJumNrS6C6daYus2Rjdtjd5
Qh+zw8gRDYnVRyX98excVuRigD8zqbRitDKFpIUtrn/sQVBNhsaLxSK8zwzt1HNy
vlSr7goPYGNr6LG5R6ygpElavxhzCuWORawYJofAJBGivIhUL9PQ9ZzHlPv/5rbZ
hM0vIg6hbqhYcfMc9oxBN2CZ2pn17vD49xPzcMWsNXYExryxwl35rDdrxCSKEmd6
KLwCoAtnB3u90Ng7ckHSO96wLkkoXnso+jjNs+ZAkSklH5ScsenuYict7lrKO0NT
xqOAju3T56ukuDbwNjBFal86QQwRLoHfVvmIzhgFv2uqh0Z1drttN+d4tnwmPx81
5uApr/oC+vucxZ5KEc7kRx2/mmxLbrBj29w+Sj3Nbdub9Nb+zgMGFfPZJlJO3+a7
kxsXQH4mTngd3ZWTv7TBiEgG3YujUQ8dF05tNeVDpBKHqEctaPCCydyzvLJCK9dK
vskEK1D/iQ4OJpCVmF427HRAVmDWmiI0yUBeXLgb/64NZNFImVRfSSUi/Udl5D1i
dI3alyqprjA2Xg7O/kBXlw/c8zt8Im0fT5TSc6hYZxxSVD9qc+wecNUOj4QXAgHx
SSyjikS6DArPWLF0AZvo9M4rF5adrcSpIQk4xqvz+h+QI0Gp3Z1bDcaVf/D+eGHY
P7jYSgKdboIxHt+wjwyeK9XuNOEiCpOOynPKhozv1LjDHWXdD5nfRNxs4A4l0FeY
ubUj9RAprLzzk77pGJK0D6rk/ADHTu1Mgw6cdnA+9pxOcZO0FDx1EXMbHsMSh7ea
`protect END_PROTECTED
