`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uKKO8riFxMo+Hp7mxOokUpeyJEzEgEIi4u4wZgeT1MbN7UnxeEAH38ddwma+8dbF
Uv88T2O/Rcyojn0j1cSVq/gEdaCabgHsfsWwI6JTiGdO7hlex8yJ8LMLrlQkzhsn
Sev45kCx0w8RdOt91JqO8ZdiBQdWRupP/ZqiIe/Y3v7o+UwtBxXepxIwshFQfzJz
AY9racYKEZnJO04wQHQwCLiBxFYlUKZEYiegfrZmW0dOBgn4jgc9DHr8p61EIBQq
Rd18JYnn1/pOGtFtAacUZBh8VO+KJhYXLY/xNB9RjE89qMtfo/Q3x2YN8IRfHkFv
xTMtJVMY2FsxASHli5hdgIPY/SlJFhyvDBIeOjfneixzSxH0mHL/L0bb/b4rynjo
ch00Auy9f0IJJ0UlOR6yrmbiAkVFxlfCu/YJ1JNxWOTHICYXpkPYqFh8h6d23o8W
`protect END_PROTECTED
