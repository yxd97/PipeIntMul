`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6Qoq8ahO1PL6Uqf91Seo1nDlvOvwduyKAj+Sc6NNoxF/zPqN4b3LxdHLaxtO7vdP
9RPqdVhDk8S9QiQn7keM3Y7W3YbAth4KJJnPGES5XqVdTBOv+45PLx1+iR63QNlH
C5g3LSn6vyrvuec0MSS/ECE9jIcHbWfR8WIavio754hufljiedxH3KGwo0zpo2Y6
tmCGq7VGsakqeqeHBs11KW74hME1nE0jAmkAiEBMyKIjWOZffXD336AseRhjCVXR
VjRxMRLwep8yaAlc4hYMTgndkwMYwpjG6jvDwCKf6ajVW/AjWUQI+pGBwmUeZAyI
IUlLb/YkgsPVXFqLoC7Q7h+wz00dMqECakks+q3lZ7Lqs15xMz2Vn9XwqXo02t3f
8xxURIAWVGzm79CC7qfEOmUtGWVrDFmvAu9m5QpIELd8yOZpmHKNl3UUJgpj/z+x
f2TlSdyiidzA9ucrdaG9enp7QFNYvJjPvPNzGnkdpnpHtqTWeFxIEFXfpAgy/Ujk
`protect END_PROTECTED
