`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e10I/5PuQ9QJ3hExSvd3bp8rb3w9M9g9es8q/1qPtki7PCaKL8CIMCjfpvjQFSJt
Hes62oWhVPeOjGpw8MzzTF6TgbVSP6Xe4ibxljoA81RfEwNuNP7Er56f6wtwSEjw
J0NgnuzoLg4ujheFRf8CwGjwU/O+fPQ/LmNTOoOcQNunYdLBp8jnwSsLBMxkAYo0
XPoNdqLwPkOGxAgf73Ik/2HKneqskLrXe4nlG7YkTU8dwN8ytRwGfjmhkFXkmRo6
7bcqIY3XyHcDYN3oDE+6/A==
`protect END_PROTECTED
