`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cJdghnLQtROdKupE1znLry7EhBGsShvp+Ku9OV+TrFvjENsKNLGlLhlB42cwvyq5
+tDDxzOtl+mM7xmZHkqcguU1XBhgZL/JKv5HwAI/Xj4OtJlu5dMqa1K2NVRIn8Od
loWFieTRx0uUJGdJMgCR8CFDUm0wyUeKGFI4d9SsHr0wx+vENI+/ARLrkwDK0Mx6
5+tTC4y5VQ2h4uH7A7pdACsxb+gynF/VccMg8nO+sT5Yk5g8jP+9xiotDApos2OL
l870ayaH+8RLq6ukysdo1SlacdF0Qo/V8aveFUsBwJJU+/5lSbYM2PyLCUf7zwTI
z8oU7BxWjtFrZXcTqInE7ajwT5BcL7+B2p1z4tra66WScZFPVJw8K088Vkl8kSf7
`protect END_PROTECTED
