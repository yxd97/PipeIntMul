`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pRsM/dThx8sNMnXbiyeIW4ltci69E39JEuqF/0xGp3db4e0doEPXI1pP8HzGXu0V
Lbi6zg61fMJCIvR0HIOAmrpV7DoCxOYxl2nhEqP9r7caIdmuCsVPNQ0Q4RBwn3JW
hhIHWx6KopcTNhlpGKjDzrVI5iFlSJvdPN2ZANN1P+aiTkfsZxeU7UPGFei87Mnb
YHqzOZy2+G3wS89Dlby8PoEnl3Tu/fw+pU4+mWdxhN7Thwb77fyoh7+OmCW4k8AO
9notbh36ywoy2TbVIcBR6JPKZn4mZmEhyhmFeKcIFWGEFtQk7/R+dqUNL20JNIrz
LegJIw3QGr+S5YzMQay0DO4oivvdrDvbMtfHQz7dt33lCffJvEIpd59cXgZa0C+p
SKWtGlrEbH0Gg59WJxS1kHMe16lotE/cqRSuCBn4cic=
`protect END_PROTECTED
