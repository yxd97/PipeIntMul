library verilog;
use verilog.vl_types.all;
entity IBUFG_LVDCI_DV2_18 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUFG_LVDCI_DV2_18;
