`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vSpTwTNhrLSeDMF5PxvQCLWw/uWEmf4GchpE9M1ZTjk7VVbgE7HNwfmm13rJ0127
VUZO3L4Bc12M2U2C28egjMmxGfkOen9+TVB2N6uVHK+5IvpTd57PgtgnivE9VSs/
HDBQtJ4vO/Opz0pWUaAGoAUN2gNZ9rSGWyL0UwuEAAYqdoSkVyol23qZQjZDQLzL
3aUoLCUUjyE7lenMxwQOcLdanf/8DpOP4BPeCeKWqYbWfEZx2g1xm5dc4WGa1QcO
prDmf9C7Gyuh83ZiTz0saQ==
`protect END_PROTECTED
