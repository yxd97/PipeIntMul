`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iznePa2RXy2Y38K+PEFwFuGt1VxmYE3NKqJxe1s3LDAqZeVxoVQCWrFT40rfoxbt
VFGPrbb6Tl965E8lVCt6Xb1PM9eTMzp8uMacmqucJ3eHRmX60YmpSiyEtJlv1h5g
3pRNNYbNwte04IhREOEgq2gmWgDPt7t0MUp9Q0O/3ITF5Q7X3fMLQkqAyAtTZRLk
dTo32kl09b3cahSfYezMzuPAaa4w5PxC4UBMvFtV0hLTCkEiPUQKbsJ5zVbUELs2
k0RCk5xcAG5YGaIgi1F9uZ2wEHfJ3hT67YmC1G9c8YeRdyU95CANAjcgNVHBiPJf
6vuQm53WS6pnm+gKsxLstXqSQ/00fY+gVquSHhWXqEdloMhrJOfHN8po1sFFPCMI
9Uo//iN1QGbEPU1OZ1KtzcBvjElYKBYZdVT07b23lY43DU/wOKov2CLupGN/JkrS
tey6OOYuMSVosrNTe+BzFZmuUnkg94e1Bx5qpB0J88cVCwM2anpvFay7zcnHUSh/
0OR6K2zK1f8Clhu5PvCHJ2y3aNS2zC6R9+oBWHY/zMzDl2gP2LIdimvdAaUM8eu9
TOJZw5g86w7uNXoU9v8K/bzGG6C/+vubBYpfonpuWdI=
`protect END_PROTECTED
