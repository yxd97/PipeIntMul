`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CmAya1Y9ZHqDENLzT3gORz+6dJ23UvgBEB8/CNbQpd7VO7cOaLu6wohM87xibv4I
yJ34efm7Eo7qk2UA4yc7GsGZ6spKkMjAvcIoOEV1I5X4hl3wVJ0bBFnOWKnDgROP
ver0QibvRaosOiS9M8gtrdyywEAjd5eNiRGlSUzQgnqy2WTLqs3dpGgA9Ez08a8E
1aE/9EMWDotNtG1eOJVsgYY8gw/4qkQzllHZFII+SMINPH2lmcBcjzBoOnydITBU
Hrm8e47UgT6YR07/PRyIVXjis3bAhxBVnoN5AhymjsurCBf5rwamW9BVW3WTxXmk
xu0iMKDJP8OzNNE0gZ3ekxXMIdxaMPP7Qs5CcTPsD8E+d9TZum2ygLZMr8DKi3aE
vSsK93juuKy2QxbY2ZhLgtlXLIVPO6vLIomHOxmb5+FVrra7wqRdIOoNOztB7y25
2MLNdXx5WseSka1+yJNlGv/3MDKvRuzyNESg3iAPEUeOPzdBl8IriWMN9hR/9ssK
iscacxeguK7Oq5oq3l/KVDFZPmn0tOfWLdSNTpruskl32KSzryZmArTwxqAngGvb
16t6For4q571v3q7783qrSHqVmZFAkVqGxWTI8ZCxEuSxH9OEYMKMUHNmzH4AM7J
SlIo8017z4qgjxDoKyxSPBGcT0fpQWTE7gIJp4j3tjWqYj0VQe/HLdsMBw2ZF757
Wf/7dYwbXnG8fWuVsz0cYxW16+m4A69IaSmQQI0VhZM4THcdJATdyir/2djcsQOz
dhsKYECBqDVHIxdWvwYnrbRs1zB8f31MtMTi4kjlt4nGi5Kb5lTPZQwnpl2cIxoB
oaLUrWjZOtrHle5G0JrUx8bzXrznsAUWuPtJZ6xE6Cbduv22sVQ8NEV7GzGeyGfj
p00Ir+HPqVxkUg/j8G5VW504kcaN0Q2MxCjQLpgbIphGiWzdr85IdcEVMOKxePQa
1Y3wmdcPObpXVwdtzydDGfsyhIMn84nvWZ+y24Na1mM=
`protect END_PROTECTED
