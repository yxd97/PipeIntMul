`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PoXIQnyRJXXGf0FIRr07JRojivvB932fDix+CKsnQAZl0Vq5zSrgLAuo8YOcf9ls
AyrA0dt9g0nWISrDL7yQ9yaaziqJKymg4nuJfWWloHYs8dUegylb0MLmQSmK0JKt
4YRn35D7zc8Zv9O7fGcSbe6W3KQ04596r1C4bjaBWM4+hIFnc05Ix0WiG2yyNO/4
i2TYurUOivT6sgIyuVAQNXR3jCSEaP49BoMcNbpLwLXgce7+7dCdFdBgC23gBIWE
avBteL03GZXFu2qUidMZD2ldh2QJ2qr3SyGqExK/NMYQdG/knBmSKoPRrKp7S6FW
BEDC9NYPWTXrbPOFPszI3WUx1wgfk4QPcbvUd0MK+IA=
`protect END_PROTECTED
