`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Av2AKPPDS+6ujLAf7CQfixEI4kaP4KSKUHVhADniDVP5evKlU1U1YzUkHbtMROiK
nxtJO3tUrqqazPtdYCeBudjdA+3V/mVZs5HwdpodRWg2eWjp+HnXjJLMiXKR5pSz
xiqXjtqiVJ9F+0cJr4XPOQvJmeUxBTdnz7ktjk7fddXQpswxVJRSC7AlkIc4+x5P
Yj7zlARQz/85BOFdLMLP6ZrS2K7K5NZ1JnWE+z772vDtHCncH9TJxUXVM56wAC2l
oHMeEqxDlhuqVtyMeL+c21UDh7g4lg1486wewU71aYRw2LjGSr1+xGIYdrL+dkau
ugiwhCYhTF4mmLiRRmlxv5loF4F3+tW9jYUAPRw7G6h+5+GJNNggUiSAzg+vfwrl
ZbDj/ApAf+MQ486XQRQ6yIIPEkdwrya7s8ljOo8+hkTvutE67HpoW5NoJcdO6dJn
HPssbOK0jviqki1oT/FGPOYgC136OV3bZYM4ekeoOdzukCHx0f032LgCsh7isqxF
Gpo8PKny3/0O/vVWZDq8qDXuTjstnCe9NxioZ368fb7HFJVMJpJJgcTFAdDWIF9L
1TcfyJF+PjmVUySlw7eFF+6d4znL4U863LrdjIL/TxILz915M6DhDkTQ1EE/8rHH
dZrqWhWISsOqbogwoCqSB5OU1wBtiTLZVGHw1DTeTne9JFMK0ID1QcpSScq8YNaW
GFrhwr1GE6evd7qX0PQ+O7SMuKq7nh38vvpSIgulMd839pRV9iG7hHgppBVt2H7J
ZXaE0Z5c8lyc9eZEYZrT3W1iQmizWl4T40X79o47JiKIkRsXo+z2geZa0xtbQO/y
`protect END_PROTECTED
