`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3lQDksAeP1en9QZ3532LMqmVpNVX+QWGFJ42fQaxDNcJjoByhjyL2+shVJMYMSr
f+n7DwbK5YmIOPWgtwLPeFHYV/YjaqRTjLTLv+DIL/IlDiSnXZk18nQBfFwknDP4
kDL0C0PVF4SpoltO8eLFay+502Y47zWj98H5/cSn7xz9JLFGgTSqi7VfFj+YEZJi
CmLi6oVXcXzeBygKmyjwruxxRCO6miF1PkscRD0LgDg557lewAAjRF+53BNLHuhS
ywl4EDE5/rY4vthhiONoiYwzz9fnkF0N6aE/G35dK+CfW9gB5Diw50lNJMi05h2o
uhELI6I1U7ye3zrSTvLH3Q==
`protect END_PROTECTED
