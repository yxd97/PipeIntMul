`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Uhn0hwGXohQHakqPYOeIZ047ZWv+2ueApxTzT+52LWOJ28iIsshPfSaya3KKD63W
iYf6atPvf3FLHf57iZ9icKiO1ZUwtsAX/PxY3yda2t37d+MSqnfEuFx8vNuNyM6t
yExpyfWnGprdsrrW0kf6Urgkw+ef6B8erNVqb2siVTAuUALn/4BYJu/uGkw9LBF9
SZ7Y1BAJX2+rGl5rkTLCPmjF+mAoyO47myT9isa7NTcLFVFuxHgXfkSva/eou3YW
9SwT2NCbo57cprR7okBKYCGsccdO458sD0tmEKq9xh3upCu1rXFSy1Dgwkg6NWrX
rA1tROcxZIFMIJmoGeOk+SAj+jm1ktnZnwDN8prMfC6DnhbdAXde9lLB0TvQ0735
frjzzXUd9MI5rKIFiGYmpeDSI3BlC1iP8RwRkbqBZc8SizCGVZb2LNINMsFa8nUq
Tzdny4uhyH2x0PMpz05lA9t4L/z1GjBabo0eXxNVc3tYOMsKBjJiy/T1GiC0Rcqu
LbI/DIwwuHFCFdHjCSCMkBfTvObkARA9vJr/QczqMP9FSJ5I8Gm+AW529mS7Wh3u
vMC8nwujLgkPbtw7ccATnDoeeiQx/bviB0WjOryImWHn0diVgPIKUpG4H3KdVD5/
iAz5WNUOKE3cwjZGU4Ae1j8c+se2xPh5TWma13wj/dVmD1+ujflK+TBO13U4x0zu
q2BZsEBPRUr0YE23SrOz0Op6S9lTLTtZaxJR9+vGPQPGvR7FGOMoamuyhsig/eOW
8xUCIVTeaT9MyHj6l+TmQUVmq1zUbgMSHg+MJNzZGGXNTuQRmepYnDNfRXuVh94Q
rBkacxsU91tVW8C15f+nQuRKa4SbLPh/6HjnGfEws6V2y+4PzPJg8QgbBnT6diKf
gRF0gyJCRgWubYoPAldnnhP4c+Yly8p/MUvt4nDz9OdKcf5WtzU+CZ1pb/RtjkXA
4im3tDc36k8fvXCJ3DapvQQFuBqn1pRdGkDGGw7QOwWIs92rOevY/jawCpq8u/un
OUycyCb12ZkVQ2dkxkUECubdCg+XA+5NoOsYrg9Hwfk=
`protect END_PROTECTED
