`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A1N4I1oEjImh3Hegkf3+7SibHp4qnWkVbLBlzZZJ0/G1ujAeGNvBRMeELRETq7oe
d3tTRLEarT0oegsUgDwG5tlddnqk3BHKoRjdYVvvZz+1PuKWd/HF2DqZIKDw5t0V
UdFDckeB51CKIn9AyfixIYjvJ1XWtIEseWBSxTaswwVcCCvdd2NDbYQJ9luTUYHl
x+cEKlF4BOXuAjKQKnR4SD9gSX9HvaetKjKbfnzyD34yF1VWXOErDnaJBSPBH0Wb
KZC0TKB62yUNGp2MVtdn2YomFyJVRkx3OsbzjWoZvKTz+BL07MHQz3f1acPIwWgV
OlSpXXuRThGaTgiDjLviE5sUs9CyzwAAiUl1bg1TuCgbqpkodTEi4nBL6B+8jf4v
IP4arJaqk6pR1DeqNo6694PvHvHEE/G9ZBY6DyZKUi8=
`protect END_PROTECTED
