`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sxzdL0rFNtmXU/THGdNM6CqbqlkE7oJdn+iCv21o6t4Yg0CejVc4Cr+eBoYD0lao
sDctIpD6IKnawJ7NE4X3HS7nEvEg+YT6gPj+WAzQvbXPz867QY13j+6n6rkZkldd
i0LSa2tRCCdgESeAcZ3BlrZ4o4nfaHdvjekbOXdJ4NfOhrfpln4YaXf+Jf0DQ2aN
vlwunTryB+Z1HAv9Uf0vIJ6nAKNIbdyH3NLZl0O3SHZaZXpcII8YJ/bDmaPAb0Hv
VJq4eHh1sF5Lt0ezGcyOp8Fxic4FsNRc+B+XQRNwYoTTXcei4lIGr+uI6ly89Qz0
r9Hf7mMPRPPVQ+rDhLsGGcU17TE4l3Q1dEV4wHHcGPaIhkJF5b/AQ6sa6CeHhLUR
kvPqI9w+SMgrHsJ3tpJl2i837HKiATBg0MaXpdsXzcL53lz7OKNXnXfmniAW9Yfh
RsyWTFJ2uBEkR+MHI/VW4+iqCAmaZUTLDXEYZrF9w1XpiA9cbsRDldgDskuenOFE
GmSLwC4vaDbIhjR5+8U7UcROv3NEV4cXxUWG8xcj0aDzSYpeP+Blc4JkpayGa/x8
8I3Mb/7iePhvUkXKuJAxStzV/x6NZR1W1jvsx1scNaY5Cgid7QWV6qWASt4T5NT5
dIlkg2s3o8rsYfe2nMEqknBXnP9PmCh5WVCLnHpDQxPcvyAXjCHn7L2Jqs859X/2
gqjwi00l7CjuhNKqWxiMfEE3Ualx8cQEj8vQX+NinMEIrw5oAbVCE0jnh5onE8Y7
Orx2M1ek/maF5J4veGtAtc4ueyW4bkelxdJAn50AhRVtnsTjfrjwGDbNeJIj+odf
/910DGl2/Kn/Y1HHzaxZNxNokeICEy1hLNvFD74yLNXvF7NLH0snsIRPQUke5qkF
1wig6afH+J87FjhFCiNsbCERX4T6ZanwWry2uajJ5Q/GnguD0LekghHSyKiuXTxC
ZgwUf/AO4gd7K/vAimSDgNujq2IjxDLhflbRE7wVY1XhgU80Z3JeCxGEu8Sw0RHj
cxyn79s3XGM+YvT5X6d33Fz8UtL7JRRC2FczY8BiKsDr8yUVLQLdW7fueBbj1uvt
z9OXeyA8oz2NACy6VUUueRB3eI4o4PTNE5/N5lD8bKbJ1t7WCHZKYwdbDI15gQre
kUQrn9qd66/GpIoF4R15DDs8yb/PvY7pTJlM1M29bYM0HAhJxBhC/ge5sBAH8+F5
eRz4HuqxQSwNkIe1QHk1OFdRJOrDkx+W8PStU4Y/rX8SyOK7+gDiS4zepjgr/da5
2AmVg5vqh/QJdrsOKzwm0ae7K9N3731wa4DLdpRv7RmZbHclxgF0tx7X3sqzBRdr
XQIuy5/xc9/TDfuYB0gv2L3XC9WaIVoXYnUC+yWaZPqRegh7eM6QA4AEvvaZANu4
R//1cxsBcgWBWRo10/t8ULD2HXBGIeaNFlwlqIHDJ41gz41o3cmmD/F++yoK1DPe
A6n6UGf4lkp923I/NUNyDmSnjiDKqG26WwuQAkCB9GS3eRpVeORwea1+cPlvhj8A
PDcZPUC3sPEG375ZlOibN8botMby+bi/hmW9M6N+QuOYYyEtDrzy0PjEZR6sHd23
LCyrtYeCjhpednoAHboHXWZ01V20pq2OXPBpS1nNCijk6z7dlsiXmj7IyFYXQnw8
RtdEndXXqIMhvMYlfP8SNcTk4jrvfvne41swRPwo6/f8AaLGezHBy2+yRSdhvJst
nfPldPk36a5tXvThIY84kBm7cAA32HWfDmTJNYCAkdVRjoWnHVo9Trh/nMCn6mHK
aQOEub9vAz6Mr1iNU2hFOodEhTqu3d+cBQRpL60ZqYTU81YvGCsyzxSSF9F4VXvC
QfteMSUXVnVDBECcYDRz80lz2EWLGEavn0fqyfxO5/ykTqTxA0xgYWJZpPLaDRho
lYn8aUgUx+vuYJ0wwXuAZE62YOLTygJ+s+rNwwUg20MBK6HryG+U8rdl07Tl7BJd
vLFMwDdgsmmtlxhA1VfZ2S0owAw3wL9cMzYgVbvAP11AmmZwZKe3rXSa5flXV1Mp
OujtF2ru71ptpKK+ThVRrAx+kXPu4rTCU7JCUw5afbDeq/A0a4RPcKgC45D/o+w2
PM6o+1dgLnu9EAllxkZP4ol2gEst/ldXXOhpc8Ddds7thrEtIEdnZlSWk0Vn4Z3l
Pv+cPUjMIWwU6HhqsXjDjo5FOL1yOBShPNafQa3umGD9vtBB5bW6s0+Jzq0BkDea
fVefYw8Zi1DytS4SgsiZWGzalOLTMk1l2FZmIfNCbeRy4+UBOxM4ImgWFbokp2EG
g+Rvnv0yw26Jgd6aNpVdZZ4xXkt37skdicplsUD564ylOfLChAHGUYEHd/apUd5d
f7zTzjAFU/Cfn6wSbI2k71DMZx8+8+kAm6RlJzT3otG9uacKXFD64qI3TxqsOCL3
HDib+E8TIIZqt6cEpj2WbqtYpRHS81lTdtqmrxneEHkazgEkauXk7hjmlR48TI7X
/L7UaQCLbTNfsNLvanSoioOdrOO/x/ykNswL8siQpMseovfJCygnSotd04Xsya1b
uoekOee2CLclbXIYUsGn1tfBJiprDPGNEqjzrF+k0HHyD+KpF7ZCz01cPG3w76RN
2DbYgUQGNO/EpkQ3FD0Nl0Y68NG2bo4IFYdc8tuS6U6Ub1CuqHi82FewsvUkPCtr
o8mcUf3YO0qki60kGE+yzGD1QcYcdadJZ0kHvDMTzTlxmFJvx96FERQou46ZP5tO
T1nrj96m2DgaLFbwzlqpARgdGYYkT/8zY5KLS2kMSp/oB0iwLNji68rIZysSov9o
YUs1k0cr44gp1o0NvvkyL6O+tUr+9+pUQHub8bfUGMBmwWEREgiSqC6qaJH+PmVE
o4e/VDhSkvVTpNFZw+83qRAYUTQxMxdFFYiWJ/HU7ndShBfaQL9HeYRLe6mHPaZa
0STPM3WHdRaWgIgxfmkjpk6Kpog1Mgf4Y+z+rw1liK9Nni0bxHPpfHhIafA/GhGt
VkzgOm4lMRlP9kGfcMdGdyvCtttF69VIrdEWEh8nNY+wu+BfVHUhZR+zyy7izVXq
Mgw7EuzPGfOiQLUWDAgDvM4O3dhZ/+Yo2BUpT1iKXmSQ99UJxzsQgpJ2M9ieko+R
ilXvPzEBfws0h4YKpJxqY+IQHVVE0SVp9sysQAMH0G0NSJiUUhpBK3aKaNOD6AxY
QyLOtPIm6N7DRXZX/ItaMdIB0P4gcQUoE5bIebqSA6SA3PJCECuno1wg+EZID6Lj
cWsMg4K43B5I/5MR4l2z6od9arkJIvH+GuysNSz4iwTZQqG79hjAsomDGCr0howb
BFPIEDBWIwL4cnJQ1UvcvXDXgL0asX+12UcYEo+knDG4EjKiuB7NFjxTJroA33k6
MPu4CoL+8/U8HUaqYx/6H+YoQMJXUotqYq3Vq40hsJScejleD6N4Hh5pwmgKzZ6C
RjB8sVHJjie46RKBmeNDfmYvZkxOZ6GbHtQkSuCsXPaqWZWI4VJpD9qpUl77ChoD
rTjXst+YVr+2/x3QdQnB3Uy4B8rW1zZuHb6H7yPYNy5naUhYen3XDsCHLD0c2bHb
cUmtwzRXy6dc7G45Sz/cBovRgJcdMrybFtKhE5ZMOJJKZL0lWyV11Lb7IwFLKF3O
L3TcjZ790GyOca6vfPjvP58o0n8wb9lA/uqSkValeqwDsUQkjnQtHz4nXzENSTsv
De2lYFNxtwnJB5TTzMOdUO7mqproGRoKFTHLblp29PM1fQeNf+njS52W3tXs7ldj
aXth/E4MoX2SFsCZIabxLGqsMZ6eQypaiScGMX8laSSMjuWnQiXPlKy3iOCazm7x
gCXjhnRGZU48Zo2bzZ1zrBLISIk6ehCmlqcQRdbxIPoq24K4NtmTA6JbNwQCiFKQ
xOLSMMQ9CSKpCPMk2ZKjlzPQJGzdtt9ZYy5okDvN0WPpxjbXNPVsHFOmmcVTGmyE
0rNhRAO1pMLu0DPyCRcV++oJByJrP6+Hiz0XdJJRJBdpmtyCWQ3qcgVhyicxE4uX
7YSmuIexBu0WsStQZ9dr7XzEFLkzo+gCuIC4SEVJD36kHHa0xxiFQ7fTJu5VQVo1
zIk7Gfcl8wlL3rR7F+G/OdrzXiO/Ia+cOjbp+rFS+93szanmVZ6xbxYvWO3hklo3
Y5bCBjy4ZmpLI+lvo+RI8kcHTBlZ4P2UnuLKo2lhj67v6YMkEKlbiL5ODt0Tj+Xb
vqOOfRSCpr65OWPgEHq4epoB69keRH+2eTXPo2sc0OiUmIbT00HPXaUmaFoEp+tZ
hsX5AvAqd+0bIfNC2RGtNM1yK4sYSxzowBpLxXgMqHnW8gmyOUkdhCr3EXW1lMjH
evmyZ1JEfmmjqJG7ds9fRpS7KEf+l7EZARDAZ4VMU4vy8EeQuNRFUX6npwJ74VB9
uBQ0Xnc4l6tURFC595b0PG1PUEjR5+3al146a1eiJfIsPKhrsnfZ5TGybEwlH2l1
ftoYLHTPp9pJEIDl2bS6ofgVZLi/k0eIOVn2+eIs+X3saCIavv/fWZM65RHFbhi0
qPPkBg4m6PHdUlyIMomoJkI2yYHNWk4x8okBkwmG+Q8DX9YbXG9dwva161XIMBkU
/Kbx2W0PYYiaQa8y8BBtCCJDsWUobbeRXb0NS0uj7lHya8xX0ghNa+WryQ36BGqo
+Klal/9fYgGlCyA1Fs6PddpqYIiKMFs5Hz8dyLQBbdgAYpg1fGNu0pGR9NgeYRWb
ok50+gckZAZpuyxbCEXQvfNi7raxm6Mx7g0UILCbF5O3HyHZqYX2TMuFveOjICC6
bG3AYclyay9hSW8xY0ZDWMJCEs1OdLuQnQ9ezhw2D1WH7xkHNod0GMBBlPzXKU40
OLFI06TBdgAtkXJ5EEE8DdSyi28nVBa3+WX1IiEF0cZOiSBFKynB5oZLiHAfwdMO
4dtPV0KRQ5U+v4RY9lsFd45uJ2FEX26L3jiCF6H+uxj8mDqnNQ3LyMtRh2IAuo1C
DBhQdmhiKXm+o+6xTU9U9Z9Qt98ZpBC1Zo6Aoo6pTrOuvewn75wf3/PAfDtR5CqP
86ENyZZROufOChvTR6Wd3nKOUBkKChGLWwVwRNsv80IIRdNUoqLVPwgRF5XQbWqj
MkuGzfHkdm0k3YnSjqdT+yTG2h8k3XjECQHjR9K2I6u3SrHuJqhXaiKiTlulJvmJ
IgvriHFQBPEgh9PmERJLfiRA1cfbSR/+IrgKZ50bN5jquKJiNlOxftd29Nj4vaVT
5PFwOei5Ai5SXvk6GRZCJu3Ef7NT3J3OmNwA4hpl2pBW26UkKvJ+lCIQHFnTLp6p
hBetmIEV/k94nM2IghrL04ZIUFGKVymY1ZX1XE85BxIBTvXZTJqgsLGjYDuHLY8m
UF8DARSy5s2oDd7vaJUncFxcS+xAY2xLi5/0isoG/Q+KEmgmsHaognZa0MkwISVW
aZBu+sNs0vLQIylCCz1YynUxBjS6/x92rqN+OstqwH8=
`protect END_PROTECTED
