`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6QB3H6zHVr9k0ydrZ7rT7FRYTYB4LwFqa/oJC7AeEYjO+0E3+qpsKorgRbf9NDbN
GNZicHnEbW8p0vpzPwgZ1MKlNpHoXYEBWX8t+1rmOt6DTsaiskv7qsZWbzMaMzC6
AhrLsEncpP3FgAowfI2v4q6tJY8QTKOKPSEfaZJckas5pn52JMKOiwATcecy7kW2
dp8OyflJet99RWxizG8WXhBKsl0HRupDgY3qgxaVBmEYysPlITL8NM/bnDOFdglP
eVRv0hSrZ/HBLmib6nGoIeYp81IR25xXes8EsgYjGZeFHq93QIbTS51mKIQMyHuX
lzRSpjDRJnMDh9GzWpnPdjMU/VI/AT3vv89nhA6QYNVyvu+dfximEJxfx4hCrmnJ
XZErfqq0brrr5dsFl6wLgMzkEYQi5zal5QnDtN7XvbX5fUWLHbEq0LxB+4275Kfw
XB5t3V55jEc1QaK5EqkEigSuoRcG/KZ7bE1lRVc2lSjyzgEAwLMWYNM/77MT5ZWQ
6WHQdREYca0jesfRhgPHzLIuIC5HfJD/koRu3bEvPZUN6aZkh8KbR+BRwQyQVkF/
P6+no3ApSSq9USTlWBmZ9dCFUBg6XRufZ0uFvJ2NKNNfvv5kEjywWopwoIi1oQpA
BZ3zm2VAno2ghO76cnx9exabIz8JxWibOkQ2GKXZXmeZrKJnbq2LrLitG30/U0DU
8eMIMOG1t+RT8z9nuSyd/X66zJS08ToyWf/MsiX0FncCJkNE+cjI2S4aG0WiHRF4
iTQFqVYxbPFnFAKugIOlGgC/oWjO3JoBftJ10nY7LKGPhrpUz8P7GQz+lEOgmxEw
y5stIwshiAwAN9bB7+rzIKcjJixSCHxrckYMr4XfNnkeZzRiAyntbTzt346pq6QJ
a0fJNrQHcoFqDEYxOo9QYRlwRdZDnSQ3Q7eQHUU8IeP6mRYVcfJf4gIxdc1y017+
wMcf0mzeyGVzJhtp+aEjNiipjr+m1bgaflnAKC543UGiXJh+wfG+y/DlxVtZuMDz
fjQ6/0hHNLuVHOvDO5H9PlNrGPOxOj/fJXoYB0eb1Ewu/SjSmnklb6ATOrOA6YH/
mN3KbkuBWR8QL+yqz1HWaSy4MzZqbqt9nwiaDv/s9zuStoKzIyFnYXLYQZjd7GaW
5+Aeudf/12FLbT93zOFbKSKsH5sI8ySFLEMhZFBkE4j5rAAD+hGKBhMqM0KtWoDS
J9UwtrqmMS3LwDAyimPX1UpVYLdF343CtU4YZNQ9DtgEUYhYn+z6ExSyOCfr2vID
n8SitBiqxj1uLm8OsFqVZ6ApVY3WnzhB7x/rNPQgMbu00SIufWeORZVUi/uOGUM5
jSHBiISpU8Qd/YczXcsGRysCFAbW61VNavGZbloNrU4hoIziPAZ0AItHJXu7WZj4
DBTs0K0CUzBczAHFgfRco3qfWhPp8QLGsnZRV10CinAcP4JA/dixz6YU+J3Sq8Ij
xOE7HAwjbychdUEuGCxWcH6Lm20HdFRf4/+VP6GzEbMCO3N99PtJZ9/Uhn/ONB1u
0tbUFgbRR9iBxjIvoyOIeqmS/EHQ3Hkztv06ImtV9zj+Og7mVVTQtGw83sh0ivdo
C27HnLaE0LOGsqg00RHkXPoxY7RA5p3voDCuoegNFIdyJb83xRYrzZZiQG0iFA/9
MIN8j3haq6F1vB9IbJvouxQ3ZfBtXhPeXeryITQXZEt453besHhkD0oa3qjPHrWa
dNYQTfxMzHaI+NYMlQCJALCRj52KWAi8myNeInjJNg9EtZEnT8Ht1eiGzoFn8Dls
8l5YwwOR3o45405+d9YqlNedwbkeIWNQukRLTdqJHIzy5yYhJ7Plk5F8wd0qlon3
hMrEx5NgFK8C7qmJUKmetw==
`protect END_PROTECTED
