`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rmeogzG2HMhlRwZa6VHKvAZi7txCQr1jowvfZu+NIIOwjGSuO+qSjjGI7ppknUJf
30JXV7ETFiJvSJ32aFtJ/hzT6phFJA5MYwQOZbuqy/e4+bCSEjoosp+7eLr4vevx
qRR+6Pk4EQgXNQimTV6qP5yLHm1qechOppmlJXcfmekOvh0IjHAkt/69ceIH3/ik
HmrPdGMFS8xfwmPHi6vKYCU3EmAqJIk88tI+1mLN7hOQax6haZqjR2zOH2gY0DI2
K65CQtKuPi/IG6buimvL7mbE3I4NTXKfoCegcwhrsVV5f7DcmQ3XdkDQGI+g64nA
`protect END_PROTECTED
