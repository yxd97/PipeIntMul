`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4bmXhnwa6ATL2YQbtwGb9RY9mwGAH6CtNKdxCaUWfl8MsdHnl5RDhX3H1ijgmRn
VW7wV+W9Usk1C3xpgLJTH3A6MXOeMBjiqFjUAswtbvnxa1eL0ZZBaQ4xUoKfaqFF
llG3JK9+xdlzy48LQXmQRrn50pRKmAqp/GdN7VT2wcAAZIH8o99JCoxGCNWcPsxn
O1cS1JHsBorCluB1Am0JI2EZq4oczWLy8KKXVcTSkiqD/n4WthkmTMObKLreQDD/
8ffndbYJbe8FbMC5aawO8P6srFsxVUWUOOoPJrw/qK/nsfm9u7ocEjWBkHI0r+JG
FYzDGCto5ghLL/XFdVrF4w2yKU03aTF4sQfOgDBN4CWWqQwuzazRC0p8Z4E61hFG
`protect END_PROTECTED
