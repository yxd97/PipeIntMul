`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCc+mB012ltOqz59Caz48wVoXlARA0JIooHcfhefqJHO47TKiFEazn5LeQUE+mmQ
XB2CZsJYQI9N7E5KTf/e6QOrx4L59O7jCxeSbkUN0N5aO5Qn1TBnFpWH5EK5WoUH
jzIbcJhVjS7bzrWRWUFpWhg4CAiXsQj8oXcBPbegwiBQdqkip4InSEv4Jd67EB/6
IEfusFsl1m/O84dZu93ADvp/i04izHDyMydhkPRXL5ko6Scyze9YNmR/67NR6ytw
bLun5e/hl1vT+p3svktrBRU12GpO3RKb5/F52Yjmkjvw/1aL2GlbSVtDj7vTb9xv
wBOWapH7Ob0L360zWfYtzPSXM7/JXDKv1lm6vFS2HFBhIfVDQir/bwPVKDk2UTqi
e4+CM1tPDefZGmeh89tbBDzUl5o+q0Yk+JP3XQEH/UPTt66dSpukyfcGtoW2yg5W
2bGUJ6udsGtumQIp/5dEXUnJyliK9Chw/JcgiWGqMOB8OVqq/ZFNJ+scQZmfQhTP
cOVAkfobORxLRKVCJJDaurGH68dTrQxoVBqQ+gJlsiM=
`protect END_PROTECTED
