`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bF1bjat6l0ia8LuzulpdQ+YYjyNjYy9gy3pIioysQHUG4YhrzpiKAQYa5usJ4w5q
LozPJt/rcWlkZsnjhOG0sFH2PbVrz/NcJPL7NoB6KFdDQyhN4cAgmAA2pFMhrVLB
shZgArHukAtIV4GSDpuFu9VY+1lAG0gX6/DYDuzUtFJ8FkYX24W058pJaUUN4X4+
sFo3TdleWi5KyVWmJrx6DvdByYPhN2TiI96+Rljmq+el1ADUzjKEaofGyTriINWN
947YuCKPA/jUq5GKd0Gv8w0Ab11iXRO3/7UM5qI+8/U/2Vu2TpQVMWgyH9OT2Zlh
IQIcnZDDR7bFUZllVa7bIMFha/25GyLJQk+QnWJAQMnNlQACUXXNs5UFvjYj5XJx
VQrzOgBXtEFwR9yEv9hIYt3WSMO22rQOJM03M4eVJkCU/s4Jpl1DOPl9xELuC/4/
vbTLNB2q5V9iu8glouNR7cPKt6Oa+9Ws0xZy07Ml/mE1N7T5oD9Ikq968inObRZh
rb2UoNxtReephyWRsO8N/KjMNBjXxl6Y7cVd8ZfFpPjd8eK9I0IQ5hFOlp7MLeW5
DA6xiRJO85+RabkMpVO0e7uu8gwGCf+Nm23C+sr4FBQVm+RYVSoCVHu7eoywqaqC
`protect END_PROTECTED
