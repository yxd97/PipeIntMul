`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
86POTGkVMl7MUSPGa4J78Qki/YY50tH8xyKh4H3e9mXvpNuYbRHe3vnUJAfmzyr3
49H9Jta37MFkZMZk+Kvi0ZFkJc4W6wLzYufZY3exuLJIwZcMwazrWz44ITxE/3k1
1jN5g9R/4VZIgMxt74UaDnPuP3gD6QBd7nxVjxg6yoFEK+FRk+yd5DYVKWtgCZp2
63h7bLjpi5EiBKI3EtOHM0OGVYrfbMWw0bi6l65E7Tmb/34NY7zfhlQGFxRmyWiD
JimyPUcGnX40lRvxiU7pcVZEzlTT2i0Di4LO1hV0hOK9aTxxgmTpR/9m2Md8mUrV
lKzHXllllVMXSK+VGuk75jFY9HlOrSNQaXZfFwGbYIJSOkefPm7fOKPSDxfCVvUv
`protect END_PROTECTED
