`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLaDC8xwl0MErDKtUMrc3fmyE/TuySLbs2WkBMN1SFV0rtamHWmqhBCvZ/nVLrti
SxGUxCLE9dTd295Rl3Ib84Z8D0o13UEB3ejFyiupwpzVVs3uxE8OoH8KpSmWVVUW
bk4FUJ7450ROzRHVeVzrePgRCgupNjifL2NQnqbvE/SNtosYbyFIKWDIaDjvghlx
Hg/Nuc23AdRCmu/SlZ/nVaCjVI2ARJMbu4F1+CBuiHS2u8j1g5VtZtULNeXDTvhZ
`protect END_PROTECTED
