`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TO3vk0cQxmEJx3TOHdo41/9e2iDGFbRq9X4CtLroxDVhL9J0y/bnPAzGsaEGg8pB
uiDnS9aay4SdH7XElqNXamZZrvflfBGirLv6uAXxzlWjig7MA5bhVO0xUBWA8Ty2
GEGZ/v/nAjUR3o9L4vVzgCHlFl5lhasZEoeDaCUGjbpMundb5DPqunaIPeKM+Ba/
Ah5SfTrZfzWIep7rtg9W3ag9bcXgyuMybYyhp0eEGZfhfkDL+Qt3/hXB3VlA7qRP
8dp4ntFti35TqakzztwozUcaGhkwz8lnE1X+rPWzRW8Xp/wGkYKbzd2xq1BrYlY7
DjxqZ7Br8wq1oQ/A+bVpe+7CkhTQqoO0Wmw9OZ6SrLlLKJ14bitCfzoQxA83mUou
/qrJ834n6W5gQZBXfx+itfnMtEWyne7qTrkIe9VajMwRetOjzuP8cpvCPjBC8Tav
iIcz6987l8TNKMMXU9afiuioZ7KKAsrxz8RG7fxuvmN02QUz8Qhl/pjjFkz7LA0t
fibDWJWX8Pi7aVbf6dpBjXrklvfkydbG2YkO5JIjDR5Gt72yegaRhankmexagf7U
ZwKfN6uhjh31YEAyfUko4SsAB6j3coNEOOZWTxel5ec43q/wIjswS1J1FM0GjBoe
ePxqwErFsMqMzTdZds5cZKbvkBPOSmmi9OUbk0+MVcZOfqwqwyJoWibMXhjHr+xF
EQACbUabsg9k0uDi7qviWUL1IVdiQPE9lRbzQlO+pd9omLHArWi7eaZmC0d1WL0g
wdm8oBpflmvJR103hT/YdBBi2ktltKCvTzrbx4Zh96na/se7wIymEJO6Ybm5KxQ8
`protect END_PROTECTED
