`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHTWdQT7+7pvzq4vRvjVLFEb4KBY0yWy/17P56KJmAscfIST17t335wrKXBD2bFP
JbLvNUt4MLuqB+mkOCVKl6vftB+tP545z0RVb9n53oImUfuT4MCXtGdq5P3kYuZL
XQpLIhwFQ0qV4YMVrWrcCCAYZA+5AIr/5B/InFSeaXt0DNmVJQzv0upMZ9VIrwJv
Hi2rsYpDCjdRzIjGaotT1MTuT53dZWuk2tll2djvXj8gio8YYGtUd/VOnJikmfDk
pJcpBrd70t35QTTB+PAsOhJ62eo+7ae83OgLgpowkASgsgD2PNulj3HteM9PZKuw
VBgTk6y3TrvwB+ejTULUSdpCttBm+viotvmK9nSRrUL+McDNeVfd9jIgSx2i0pOZ
zlfgxA9cRw+vrIWctTE6+wL3UJ+BodtVUeuaIb/VnrwlzdjZYMdtuEIKKdKSSD62
I50+CAhlIJDSdHAgWh56ln2puqWMoLYziMs31RFSLhr4PdfDOvBeD9ez3nYyV+RW
Mayvi3smwn0OqHZXYClX2XnQCUkL7e8yrBHsdaLMG6p2zQFzkEwTlh0Wm122MyE2
UmXFADlDXTSBcQWxSRqi4HykKVj7C3vgMniJMeo2605gpoE//ivYpH0aATTKj9ND
9zkzw+czOh/x/mGaXYYadJ9ec8Yq5Rk3QocW8RsaUWSN6v5gdB7ryw5B1g0Tc2Xc
ActoWiOL8emHPx/cbAE2vaxZkmo3EMVCJXnCCj5ukZuM5rnjEThBo74ZuIifCb0p
MwIxl2Gemx3os1aVJmTPTrMPSDo/qTRHiPsSo6ZCi1vLRY4LvRHE1+J6qX7kb4ek
3TvD7sPlz8wT7Fmhf9QBwZfRJe5fnC4HYfKis/Mv+F3fKFjW4t5LuRv2Nd0nBrik
LBmE8D5eCdtXdYq/bJzupKKxfLCVuKO1b8eru6WbmhO1oKSRZJ3H9sbofrh2xF35
43k5UAKjii0oj1b7rbl0Irf5gzmAJnFsaogJEWx7pELkBDFlKSx7ZUKKh/B4eGRR
S+xdBAwy4JM8G8UWBDb4vlDIrSSBjFDCGGA4wkEance0RygUZAMRwmF7tH7ePc1h
KmIsJT6jyhRa+Un9UmyowgPIVPN/XaMAMYnOsbkOT7olK8ax2ShFWBZ5xOr5lF9+
pOlxj11I6VN0zuieEICLHnR9IUlWEtQ721qKlA2O9fPvkpL1Hx5unU7lEssNcoNV
giKdpGSL6ujMcK4+CHOuHp1cY+SiNhYt1GFYbEIbm822HXb1CUP5rI2ZRG94Aha4
TwA1T66QXHNxT4KTuwE3tLvrT5/qRjzFiJ55+kFs+i/EJIdfOFDHdNyS+ProKjsA
vfl1zRK0uUNcsMsmQNDSUCN0EWcwaPQFPWtr9DPpI0IvwML+Z+b+oL54gfO1lDpw
xD9rleRADjYz+5qTX8Vk85QVn+TjXg7xgIHx80wn05MWlPzWj7ZrBQp53ZSartRa
N8b0sEsiFNupHK1A/hlee0VYv2pN9d2SGWAsEtUjKzeAbgdmaBgmJVGczrYCqZtX
Au+V9Pk/2whf3bZDhrLVobHrU8wOAjVuzbeNp0f3WGkhBGdVlD5rr3GCN7Cg+M93
pVI0RxabWHS5uY+JFLkyhhm7ucn3mkQvtCbxBmTC+BV+SfT6+MUAH0J+CcIrAfCe
sLt94UT2yqfM/Jl7lK6JvKvncKHAdzg5AAddIN14DnvlUOF82+XVbfp9pczA4cuo
ruN3+E5ET4Tb02vGTznz0uTDQXsY1EM3bwoLzJHC4oM0rfizSLyotK+F3++zYoX5
V58AEEvO+aFD4aDXfF0hAncZgjTvM8Np67JVFxQ+gQ0fRjPkuJzpw8Vol3owcstf
g4umoxir2zh/AmX5chZjThnIhSyu9qzFyEXglfYsD4zOl/4Pefx1mUFbL3ihSurG
ozq61SrF31V6L6GI+GsU6008NHtyArCa6wC1vGmiyBaFQQqFxEwqGvFZfvCKLHGZ
SAvbGPEzmCy5UeWKG49uqU4/50H62JljVS79tFDrycuyZXCtPl5NOLYmnBuqt2zy
lJa79GyUTCrHqnFruA34pAm7RMvyXFk5CX0PFjqFfYMdMKeHtyrH+lrx7Nc3D32w
eEBkCgt+bLhND5SBgBsrzD8+2M5Jk/vZ6x1z7PdCV8UkwAI19fqNWR+I7O0Cn450
bufuNv87VmzRh9ZVdW7y5Bm8wO7juiusg2kCGNVHDbXusZphu/wf5pUyZ8ODsI+7
xokUGz+u8yCf02jqyWOc+4Z6ZdAO+DOMAPzYt6bctNjlQ48woIBAiHM22iOMIbfX
jddWn+BXKkL0TP146ojoQyCOQw+48ZF/eJ061M05cb0TyPIpiUo2W3s2lGycFlHd
ZzqmRSbD3DgbJPvG5Oiw3AX8vVa+yLwtCtXNEpD+hFZesX7XZcQua+2wdordJfTe
2fUGLy//U/qWh5y2+5ccakhHSeRbvpr/OwB2s3hDK+iLAQYHznP73uNfo5SDueNu
dSDniltfFQLu/ygTKppCHgFB8U1k8xx5oEVnPAxxKIFEfoamrJYg3zFSXorCJE/K
3PXzdJwMidCdF+xDaPJWpLWFOOuTZmYEghCPACmcwZM2ZAW/cPTKuCmopaHU8I7b
`protect END_PROTECTED
