`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EDKJT4HQOgbz+wve10hi5R0yGqP3odvlsWi4qqfuebDt8JXupzdfzAgDqASnsjdh
iv6PgTvgwGi8RdWkeaJvR4zkUl7ZPMwFQYGWCoyOmElH+2xvAEhkul2V/di4RLQ0
sFXMgxbe4QYgovgPlrPfKjvE6PqLrAkjDHBE46p4fBRAHxFiEU5geRzfsQl9IoCo
mBW1NvqtKFHmvyzfLUBSTwQo1irgi0gLsOB87DyMkevZLFhkKr8RSI66p+6RcTeK
LL5/Ev/sN7CdPwqufhkqKGDGqU3XkcZiwofQO50488D190BZwUwWBkdPhzhvs5yi
OaRp/jsxSR67q6Q3ru2dVRNvi6Ex2Fbk7IckgDo3eOJxgNnMVr+l1CIk7JaANFW9
G6lexs7uufSlgTEp7HxRIUDz673cPc1Q3MvF+WhPlh/dk3OXW3EcP8E5x3GrIufJ
LrHAhfWWLaSCwWy/b6PQx9RuhMsWnR2uH40dAu3KVRKJueR0GgQzJjnEX2mHBqmR
Vl10otTl1o/hcORgv3PHHAlZDS4uWVUnbOgcIceeZhMkVwMGZbCDVQ+zsGk2nbRu
V/9x1xPJDCRCwANM+TP1Ow3KhNxqD1Evcd//A3p+0c4gVwbKMpD5v+c2vP5ixyhd
v+uEhg0D8bBZNxBITuWSmfbvBWlnVoW5pwt+lo7Peb4fzEW9ak5HzHcHHSWuGnyx
rcHqpywx3z2A8pIKigWo4CeYu9jMC4QW6jxdc+aXy1oxwkFE5dSWb2tGyYVpPTez
ZL9h24PNkIDziiQqcXrDSpLXqBGfWyaVj0gZzBBRv0wTeUZMUP2LUPZTF3rxdDGA
DQTC4aNkOS+vz9Am5p1pBAs/j12RcSXoqJmiYpXdD9pUUPn9u0lSrkp1V4vijsix
DvE+uE2zMhbxMQrVKU81MTN3cVxBRTVbW2BuN6Vc4EjnDfjHviHRfB2UvIzZpdCx
x64rhykLi7YHBQxfg5sAqZaknYYR5DG0d3iy5dzBBUtLZ8V4PFQltfeJqSwhTGyB
L7fCjcSnrgRYD26YVpSJv283PqAn/sh/aIu8VmZWuZXnhu/dVe7ajAiEuIJXZhPZ
c8awqIplsAVhEGFPnM8Edw==
`protect END_PROTECTED
