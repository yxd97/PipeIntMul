`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YsmcfGBlfOE7uHOBPaD7ZxelEbZv3Od2+CmWhCogJF5eJP9FT7MM+v5INoUidctg
5cI3+WkAZOO4Lx6DQfUQM71lG2K6DACMA71dtwfhmwg/Z5MU5CwFVWJWfYqjeBJ/
vtzDAX3XPQkADvBN+rHKAeR7tAHjEHIrTEQxLXyN9MHzcf877mB1XOrsnpfRr6oX
lA4In+ot/gOlbFBeikfLkIuwFAbfSGHZVTfJgycOVEt94YnYOZlmpHJMju8DuHAR
EpKBAxBeILYnp75aDevXagFacwebx1taY7NyaLwnXeq7fES5rBBrG9U7rFpqRizQ
r5Hhsn6lh2y1xsmfpDZVdP2DpsPGDeLr7o7As4I3DnkTAz1u4S0mzgrDbIOnerVo
uiuG1wlAxERsQ0DkFVeVZRfDXWvkZgp3fBZPDzT+QbSRg+mpN0zKLIsK3iYIIo/7
DfqRFK8pBMv47X6IW3hMFgM99B2jx1mcXzpSSJXlUNr5uW/eT6M4701biOkLB6Gx
ajHpCRwvZNBmMmZiZs3d2NeyOp8QAm+K1s5l46nzRi8Rua+FMAcR1CiP+Ok53O9s
FyUNIgEiaA29SGvc+HbTMpYhB7FzHtc5Tmv8vXq8weWDqux2dMg2nGRZEDg3HDQX
9/0H9RSMSHelrpwLlFL0nIoqA7zPrXksF+S0kA4ArQHDQzjojvdSSQk4omfS0xZv
XwzgUjlpCtSMx7Gxg/8P+FgpZxwXwhNJB8qJ6npL2+ykGw9Z3wySkNEmUKFzP/WM
c8uOMD/8ppcmbCEyktb8KFLDByUQn1ysIL3sMIgDbll4/yQCB3rI2l+YL5K2S4n6
RCBlIgBp6iRk6sssAo5zxCZ+yL5xf+rVOnuQKOPGGCUzSohagMB0SswvaB5KGEHN
k4WeucNwOl+28RJpEFS76p4UG9EjrGgjfG+4qHSWd6FIayKdoOuirsGFEGopMOsV
Wg7XELSLWZKuEbOvLh3QWktoLfVweCvt4je7tzM0yg28ik/whPRImg7vrkEf7+yP
tEPZnxo0Xqf9DemXyYnWIAi2Vj5wZ92rSt/c/qiDn6gdJwI/j9d6tu3x6ZmBnkxZ
VkIZlPTj6QeuCCdbakPAMqgQfAmiT58vsjD5O69yEe8A0xpz8aGakyhGbeQIWc3Z
It6Y0YKYcg3gF50QBE8OYFHccLgQSM5gzAUaoUC1gIdPkksLhrz4nrGYtnoWEMw5
HUWPJDl22sv6UxXybmwaPvNOKx2LP/yWh0hSAdfwXZNGJKybV7y4c/kTcCBzNZd6
R+vXJeyJW2hoGV5yaO8ByqBSg75vWkr9qs6zjtLacahWs87LE73dB5qvfsYiezC2
GneZusd5oMvXIFMh8Dhh6tJdgqhTSzqYc8wiSq7ARo7wKrs+NFgNkcQkj0qLvp0C
tbTjSei1kaqF4C97PySWpJlV5kCpkLxyE+T3o+IIaizFKzrAvWXg86hZUTEfAuNy
VHbx16QdXGyeoDhv96bOyxCmxieMF8utpscNTYv96jLHYzIdOzrFb1kCjAXZMsg2
0y4FNMvxC9lcLXb/aUroP5OknMnE+hevW45MIVwrF2eJcH8JAjzrCmpllofDiZ1A
raUuBYtFzNvr741B+pS2gQVO6ZqwPrEK8oQjmBPduV/M0XRYYbO3IVbdP8lfJ5g/
V/TBNcVAnp4yCve85Njj/hwJvj+x8qc2FKzVPzAjon6qYW9Xy8AisbKj6YBTzeHu
6sjSzEAWF8Y5C68s1rf5Woyd/gHt7NUXYbp1ZVcT50yyjcts2l4BUhamgqorITwD
8VUHXIYr7MpB4eaJ51Nqyd0n+nuX9H3h9vn2e80PDakAQsEw0FgiF442ZJZLkJQM
o4k9JhBWm61fLQzThGTUevf2G51pF9b7oTLVz14FNy/OSn9BhkZXdU4I74JxhoLu
lhHAk2lSx8e19p42E8NLrpBlhn1fHcKJf5yFq8vIDBZ2Cbr52/8ii1TT8V33TTIb
u1jYfCkSfS0NT6BKnv6UnAjOYJOPsdcyHGnUJC9R4287Oc9k5V845DeeExJP1svX
UDBs1PWSpuo41kkTcBKIODprTvL3MfI8GIioUKHtP9gG7kWGS3g9MDnqv+zqOQ37
cGreZOKwcRNaqS2BWheOFR8MMrz6pzuvfnlNh6SF+ciSlUUolPWP4NZ81EU6NHb4
VX8GYJfKJqr86mmfFQIsihashSn1BTq5NR6vJNNfeHaYebTo7voq7mR8Mac0SFY8
v1rufxTcK/ganAqlY/u2bYsPWdk+ezOkeUBQ4bhR47SFC6NWOkh9fee1i94ZjXMC
JfaA4qJogjgo+3yHTgFuJPkIuFaR9cu5tffHN/VhdOsoLPqX6uFrWwcO+dkejdlh
WMSY//TkVK0LAjmH1pW5HfKCI8e3e/07o3qm1nr6mRu1UnOQfqNgbC19+6DMcLcn
TLkp/mewvvcf3Rd2+9gyCdjcA2uFKbbgjf4sbMrlDXSFE7UZjHPhRO3kFs0QO5tu
WffHmGEjeb4vzzc1n8De/LzQCf6sWYY316r5dwHx4clkMFtq0s42FyEG4+QTbjj1
qIdt2ZsWZ1CxODnH5AzDaoweEgYNfCjn+3dJ2kO122BVdq1gqdE1ZdVm6/ZZ3WcW
ZgMxvKKUCQEoekwrYWOK9aruPpmZo3lDZHyph0cGQU2bzByPoHenxUz9E0QolrQb
pijHoEVErQBlWd7SLo70eNM+QRWEetO3Wtfi68x48M6UmsMK4XI1QbVOS79kabG/
uwvVz4cntWcTRJKh4VI3AGaKAeTxqOJKiqJkVFelkFh9xjJZI6nsUSWJ7BXPIcTg
7wXatvv/7xEacmFnb3MOWoBaQGA/mSrNxLdbx21A+gldaErJ8Fngu4HzZGnO/Wtn
AuUiBAdj0ASTM34KhXHSJlkgrGwIIwmjgCPxanRzLF89YBoKJwpO7K8WM98wUybZ
9sufGLRW6sybAnkOuyU5itzoJKFoaCKI2QH4cowXFNv++GayETkMrjFeetR7yOhG
85vOSUrWuycq+KvH16oZRsy3aj0+EIuENfgBfIizSgPkDBZGUTtKtmGTsKHi3b+N
ofQTWFeSiAsXJA6C6BLyXx44EGh9InzdJ4Zm1J6xYiAhsRXdpiAzOjG7AGnTdPNU
Rzl7tcM/uIJrPtI5nRNVf3uU9rzQe8B5Po3qBw9tyOG5wHh98ncsGy9cg79hx5sE
aulQpI9t005sVbPv8psg7QwSS9lMSIUb7tZWHbwO8LgxuMuqNSbF9rC5OBzr/ijo
SwaRr5OdflbYK6MdLnjnNEHZW7/TtPGvyx60vrVB8tmc2TwviK32byEReg+EmcI4
T3V73wRURUtKo8TQGs/NETImUHTfDLuidLFDAHqLX0rhw0BfolHT0FrPl95+GA6T
LatiBoQguukZXm/dsqK+pRjLqxmLPss4V2+kb5jqqyRrfgQoZpz8qyyrgFsyuibs
c1uL4i3k2wDcstjbcC6ODfG1DyxnCCyS24snxCjj4acUUzZnpCOzWavaqoC+8qhH
TGT6UxXSSk732jbUSyLpaMLlkqCCyl2mXSaoVwzZ4wSTVQ1lTxSs2n0hkDyRYKQE
G6ZfbwWIrsZFC3sHH5AzxY9pIs0PCiX5asf0T0/4x9HwD1jIkaM9IW+sCIURr1U9
N2rPJTtYSsyTv2g/HOzQvEXQjophtaL9u/B6+1/8bm1xIF88CUM3lQ22uewWiDl7
YJq6GHsPIB2u4zGBByLf7NSPQHeJOj63F5AYGMUYE/1g+D3GfgEnSZa3jyU9NF3t
F/G7E/4hy95HIOzU4FcFMHxnHIxw64Iif1Sfmv1mw/dccgUJeJossMoCG6J/SvTA
RLGVm+Mu5ajjX45HjMH6x68knyQq6yH1GZgFc6FMQvcMG+xgTfI1YMw+xJH7OS3o
rrrlsKATAlxsiGKTJv6woTanLIySUVQOH6mVeJ9sB+4Uskbi3INT3sFNz/x3C40J
J3OUvmL92Qrm9MGRY/CiBdzowkYt6fVHmhX9GLXa23HpyVr9uK90kbGl4qpIifGK
W0rvgoP9oZt7/aqZCM0pDDz4aq8tnceYkT4oeJcJ7DCCZLq6gb8cSzskv7F9S2kg
mzJDFwktleaOqomRCvFApJnU1Tuq54RD9UFHGcGQALD0w7eyqfrWj2+Oq6/MWkNq
cVkTFJPGSd0yTV3OA+k+M+WQHK7XRJlbKxHm6fQ9FftUitabWuKauSW7f0H15VVa
8bl/W9WXbV5dDtRqRvWxDj5dF1dZR9KiuSnhkMXfECLeEJfTA6zgflDGL0nIocaK
ZPrLl6OmqCyQWzvDh9fHEkGc6Io3ACcmJsHzYi1Yhqp6nLbUnUNmGsoVR6Qvt0hm
7iYG22zOpoTohzZF/7mEIgsS8I8EKPZajCiEkYopwQcN0a8/XRtbOfFYUhRoMMqf
/5003D6P14lPz8brbs7IGX56yoTkfL8+30LZUAIXxg0UdkSpAD7LD9uqDLU8Box2
HEkzH0AaGAOMJAhpYW2/+EiOnSEJKjKuTWDrBDcnsKD40o0xRSR7XEPuGwTeGn8C
f0Lz2z8HLhTeEQ6oYrmO4fbz5DKwPNQr/x55qNEy2VuFlryPZr1/UdXmaFyfoIFu
qrZ54Be/5bjS87Y9BFgnYEDT7PVJbKUSA42T+OMnbA4qmUYmPnTVR4YX6mRVZcxu
P9BrEOQIYlcfe0kfnlQz6JqDJOMe/4fXkKeSdpmiK6ZGZ0lz580uyrPRIm+PMpp3
+wgzbBBvPx0+QGBdBAetgi+TyU62KjVaKej0YjlSQYoYq2q+m6n1ewhUMsOcKx/o
nPji8gyFhR0iLbhmT+ViNvXwkUXEwFogRMQKvos2C+KXZB1UW45P00nAV5y+9VCu
nwiqqSOHLXppaebM1//VJDKb4xLgscUehAjZ8wVXyeBHbbxVbU0ADhs5Kqw60c2z
+hCHqH/JIFWZqDfe2bpklpewhuAJ8XrkHH4GlaaIPJqBOkcp7VKfsGfiTwf2rFpn
YV/8ssYdAcUdPrpQ9kzgPY7xt5QwTBGdH9wcLmDhrWR+y89gmndbVdo8lWu5tlms
wPR8OZ7y+roMd6kSHut9SCuu/tz97jj7ib3clMnR4U2fIVTrmdrM69jPFFCIKehG
T5V/4rCjSK98v9EORx0urwUqgCFXWU+yGz830x1VaEh0i3hTnJ3k38F2csIqDgIS
3fUvU+d4UozDT6I4NZ1n4+JNKq6AO2+LEGntGddUyP0LXDhCazgetoh8NnDcyPg2
s+GZW7MM37eMTLtrhz48xoSn+bSH+0aRCfoU4aWtBn3vLRO3nwIFjBlcVGgOLY3j
HBedwkfOuYdUr7m9fRKBlgbqJ12i9hDgZ/UPh3dpX/97KnmU6D7/Br81KImn6MZf
iormGwlCVKa95xQqWte4Y7XUYBgcKcnK7l2FQC8EMbRuE7IJE17Y/dktpPeruhsj
zJtE29F92dFmt3w8QkOzlX2nHgifxkfByHdbMOH/rEffLcPNYJBTpKzNxWbS2nfA
j5tyG9SchQcYbI87CDsustZIO0/vNSRRRaEu1BDmPcrJbdZW1I+/CpGusdUH5i5P
7Fc9wL4bry/JMYR7f0lQuMpmPIh1DJPCLzyS89gP7dwJvzErQvuTl6rJtFbCcyC3
zW4wpaUcpeuQnq60Rmgv/6OYetCmMtigsprx3undW+mYqloC7r3XMEOLPEceoBfZ
6v2ewKmh/lKBEhZB4rNi5n4/R5pE8LWFqnPapAgggKmuOipvLVFgcOnCaCamVb9V
HzHPHBNX0oTPqEE7+G2IMglL2S6gLxxojEQYudnyX1Rb1LU5p1Eex3u5AgmYutA/
GR0VhODTvj8sty4qk1vO0u9MF8jUPATkk0k5VI4/S3yCRsnN6dc/h9zfkwAwgvP7
jNARL38Id5UUIPhmr+lbFfe4TTK8k0xXjRbBwoRWxYAAMYqdLc+keD5uMIAULf9t
XACoE0T0xGLEk2aJU59HOoGIYsDESvh+BKUnaKQbdT5fOQtkxjGXsXvB9TnofSK0
Dcuysqc+j06aB2PMyIn5PrjfbydNQMWsHPXIO5s9S0/5y/CPTs0xek3AGmYc5rym
rbVV6ug6juR2MfJB6GvCk78Qa1g8gtB97YCKRs9fqJtMbUkSXnU9FT1ZSWYJ4K7j
bFhYqjoJ18iyZnULm43Kyuh4enhXKfY4pe8qdAQIKOIXzqYOt/T5HucXnll/koMn
2UptBqlmE3QJOao+tcTm9XnFKKV94tvKCkKEUeOJ/8ZDrOJuOUh8ndMp49W5kgSC
rcVHg/iYcJThp+hIn3RXTICffRMMMDs7+qVYRhwLbXOapTnM1r2s5ZqDWP4IUTF+
x7KirGTEyf90va3a+1M3ppsoIRUKo7CGqEX4u7M17yVs+U7s9Nhxm3re67+mIxr3
g6vPJivpvIPNC+nBbCPW+MC3REOLcrG/16nODMWhqfVdfJVzuHSgOxHVOA/gfK0L
7cr6gFwWyWf5cVnaAPkUjDW4vDGf53CotKdPW0WPFzvPGyWvdBVG6dH8fX8R5DA2
zPY44aZ7BNzKQwQ8X6okdYWD/5r2dsrBsGj5tqhW6oEzBGsgs2NTD3MKbtcy6fiM
7vZ4AxtsVCYoR9t2McHsP7lg7MugMgkp8kKVMuP02z0TKSeMCsn+GQYzUvx7v5VS
KIMmbvK4E0ykljK0ORbojDL35s4gdwAOVjIHeQjsXnkb9X/SgEUiJthLM6+vq4+q
N6eow4CPdaspBp0NXbuovj8ADIPxLZE/Ci2Im9M5HuYoRD+ZpjDsVJxE6LVFl39n
wDO2s2AqjUc4+XsWx7UTwHmbRz+s+71iEwWmrVddCaSdsQ4sgR2DFlLt8BjBbHMD
C8LAd0mUlT/5njkQtIm3OFUMqLia7PnR0L/761Mi7jEUB2faJUlAfjOB1YKaN9IF
gv9DnPv05+JaBDxKPyDYQWdubzWLFEjqnutFyQNYcpBLM6U++efBcc4v9HwZ9njI
KLeVoS13iP9Qsnmx9QjABuAPyeOvdrqlcFa5Sx50aW0xyR7gJQU/XwrdvYss6AI0
1siHtlLElAQkyO2qyNtnLtcQ3epEfQRH9Sw9OF33lud2ultG/W50Q3gCpWXpL0O9
ocj6ntAgNzqoQSzZGi7XVafwEwva5aFpsQ8GkMakI49iW+fPguVh15IGh4bMNWKP
lO+BtvU2QbM2EQU+fcSAHMfdnMhPqQRHp9ATIkbRuf1NLLPAEWDA6c+z7WcErG0I
0IklvDVK91cW4SDhLCavGCRm0BqQ4ufw+OmptNMXRk0MHGgIruBExy8kAT+ppURM
SbBlPAzYafGzSh9bsEmo1wI60w0L0bf9bfOh0zyUbTiu+x4goyL2fvzOGGNDDmwx
X7kYBNp4pQ8SY0CqQCRH7yB7VJJsGKAn5eheOX3M6h7+Y6LGe2szkeQIY4KNPvvn
jOrp0ZkKC2DUJEHUgesTrHAJsTbsP4QAorLJbE2qcZhxK6a/L5oLIjWMZ7/3UbKL
hMltMfwyE/bOhI0PBAZ1qMB/fwWNt9psgkkO7dj7PAL+3sLn7xRA4AQ2sJ22HULR
vjrbGtKTSQrzgWWWCY5RS3Y/kGjXnchSGAVGSR5POQQbDdIWZ5w6SoMkLHnr2BtJ
C3QwIqfz3qzaEMW7CBsT0EmxF1BX+qd5z87lDoPxGbnw2zPCFbKFQVPcDTO2WweJ
if96QrN3Mlif39I3AZ7eRiQga9q3qctRQtjimwbxXq9WsaOCqk0cyOb5MEaNWQSa
S1EAaG3gh8rbWFSXOtjbrE9GpNN3yOwA8kBbi8jMAWQbdzQtVKPUwZ3Y/hnuEm+6
/Tgh9huueyksfjpH6A/Ys3yrez7ogdiFNm65wZWc2F4Ts7flq+DqvP1bEetBnZ8t
WeF8eMrQ7XJrWZv1bPnIGilGKNAyFMMpSf60fmSs4fwHHG7USWfxPQKtfcyMhlHf
gAeXc86AHQkuiLbZxgiybxDOZHUZnDaPcrkwrwAW7wGBdBcR8Fuv0UKk9H8l5h87
VxNfa0qOLEah+/QL654Ar+r49HYJifQ/i0DZ+VuigF7yq/qKHiLmyZoQWKGHiCq6
GkHJKcrrVMsvrs4EnzGrtZFPpoZHuvD9jMFevBx+sQKnDPyjx4hxklbKgiIkG1IM
7TIY/A34PCfLpb6Ksg0e/ie6yQCuyG7kydtajmNPt32a/aJZ5+HXJLbKUfXD7EwG
wysgHPFUebtxdfhzN5uOAEV1Ey/FYpqrD7KX1cDDq9lL9frSeRj1XrENyA8fwmAf
3fQvGku+LtbinFAKVkYbo76aPrpc4ccjhQLerZJFivUO6F/fWE+tXJ2b7eECUT97
2u94hbh7BO6Gptkv9o7o7Mpf4WTzzNG173DNLItyfL5j8fLz0/ZrB6vq2Lpxwmmj
jX2xExww7e3DBLvTzDTzLk+/lokkptmuHdAD2sFnynaKz2jd8MME0SDr91IS6lWT
toKU357HpEZ+GF7RlgAfbOapnFttMpPTW71QAG4Oxfq4SpAzrD82kiXtqdwhgEmB
HosCY30pnQMXqPDoOlYH6wKgC68IWF/tmtZhk1hg0bWlg/iBNLtS0j+iphnZjptf
FJ8ecnv4uID1Oz0wWlrKu8R2VymN1bfwBVZ42RARidoEHKkf+1GIoxmbiLiGduub
uj20TxgCq/TKEwBhGtRRoYAwaHpC7N+ykF5NRyUcF2VuK9r7ugBdRiZb4zKibcYv
s0kFGrLO2W03pgBQqhyqE0d4NowTbvm54prhnPQJJmep4a1R18aCUk3mKInqewFu
1+tV26jpswTKVyNdlUwtekHEZshwYmVKndozTRoVX8VdIJtGOILoc5ReR8zQqBRs
Dk2VGyGIukI1x4AVWUfM7aWrbgbgjTbxPdvdupxmsFB/EHfKdKqirRjE8WtOvJ6w
6SrLwdnHH0eM3urpaDNXCvU7GX6hXjGQcb+NXbGcXyPDyxHKJiL31KZ6YvZx0Wv8
/8RdAj3GYM/2QcCMNAeW5heZZzwdT2rIVq7+qJCFCFNcRTVxEaoLGv3iLVpd/jDt
WiAWfNLDLcOH7A4vO+Ttv3mrTpolg7W9MIpRE/D7G/ec4cEsb8BDjULXIUizgoGS
C6HbxStOgwR0TrpjivvqR0MNvcjVAvleP+TiHbLRyWoETElOcSdBzfNFJx54n/r2
ufSHYlqCl4b6BlcDVlKt7MJQUP6c3YpXkEJbd8JMYV1F9mSsdqOHcRXsjQn2WQSx
Wbxwdx0bKKRMxj7ZQAZS/oHTEWFns4Usz9bNHZ//YYC8iQO1DAryAMHj7KxILHi+
V2oipG61kQ4PXLhoekwJX/l+BlWc3xz0sMDvYVrdpdEFb55onJxhKmd/TqoN2aPf
2vm5Ju4YEfcwYCn9mQHqUzhCtB0p1Boemr+m8QqgzKmcXCWUCA7uyrZFFboO2jZE
1w7l0KiNj+fhhp0mKFZixlSaGKDnoVK53rHGme2sUsJAOlpACXAsibXTTq9M6lpL
7YuBxZH+y+QVQvJ+crahDwNeo5pLXOEOQzmogB1VDUJP0snK6Avfy3rLeIF0055p
hGECr7OE6eWeFZO4J/kjN8O3JeSd/OaOt7hhKswv+lcJCNZz0EZbcGvqR8Zmi8i5
qI17RQf0jN2i3itm7r9bJYxSUJiHUkRBU8g/wbiEPoBStvFMxDAdaU5okN/+/n4G
lXEMZYIyyUTLFxZsrCKIrPEAGsBbQlS4BD2YqyBVdqkhwF+Zv3oEWj/p2AApBXNY
Tveru76OPjgVmpz8lukjEE4zs85w/+WAD+kQhcr1LtReVd6ACUITvUF7brlb/eRU
5HrSfyno9/2X2pT0aGu3lUaC5aJ0l9z35a/If8C3slCTs3wYnDgSb7GmgfLwGOyV
gWLCvVaamklFeQFMU9zTryIhOnH6kBSoIxnmuvfs5Bv5ImG9eUqwxmE/pvYKztRl
xIGvAGOw80Bt/AgcMlQJ4fMDbEJNO/VOqDiUa8h1oFcnW56+KjE9Mq58g4SsTVi6
ZuIcrNIu7oTC7eJpWdPQJbd+lBk1OHnop/0G+3FQvS4mTcGfLnPYxvPxoghIxGuu
tRVL4fdEgw5Q0h4AP270LoMVdL68+vOJSpf8rzdGz72W2XZZf2oAmC0od7mcNrZy
s3qoXuyvHxnZuQvQ7bwXrQ==
`protect END_PROTECTED
