`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pXFWxpjGKS8i8EKiJj6p4lXQNOVMVX/CKEBUyYcyJBcRC68deK7xPizCla/NSMw
AfucUiGRCHh58DehWww2z+Q96zBaKpyNAtYljcy/zWLxcgfJQH+ChiLt6Rr4KCDq
U0e+7AWP6xlu86mGA3RHEilGH/q6FQDQYM4sPUuIqRO9aZebBAoXP9DLHoiGdRT0
vok6FT5dk7L6s0ip92k3FxLWUzyabFSkp1MGisOIovg+E+V4QzFZNbb0W8NkbyPm
fYJryO4H0OXgjfPmaaPES821R1Q+4SfCg39C+0CQo7e+IF0zeDI2FoDruMuznjzE
FZfBSPWnQIl5zlub1qvzZxwrN0odxDtYqzxpFMRRQ67BU6YszyKwLr17C1w4tAlk
G3IQwGtScWBCJscfjNETWvMrf4uIR6l7tJVNL/9f6NVrcEL1ZylxycUqzjctck4X
23NG1I0VX05l+y7Q5BERksdNzzroJVIym83Rz5FVIbUB5iV9WIujU7VNfRwO6FId
F+C0LLDEE3Rb3j1Wy/mDa6JVnqB2ITo/KoIq0uMPc+h4ilgQnMC/1bOcPVeSOxGB
cMxde1WH2NymBvq7+rc315RpIVInBVRy9TJIF/0Ri7UD+n8TcfzNSZrjUJnMb4+e
DpZ4nWCOcovNiO90rLX4olVKjUsLmGw1zkLqvWmaI5H1lf4vRzBLkK+29rH2OKko
Uq0gR9CfLdYInXmtEgyeSGhHIZN+k0mZGH8vQMniUE51wArKmu3JmmWHA+pCZh3Z
yM/UzaHjPJps66myKC7FUoq5KmqlRY3ouObLkKOuLaUf3Csq6gm7CcETXd+Q7QKk
zuL9tvs4/fZmNLQ1GIjQxM3C+TLEJRXgg08Y1ankXVz67dTNxBeNwjsTBgsedivK
vMkc2/OMsTcaS7mJedjyEYj/jxGncTMy+Yt6asQ2PUnF0cR4qTGz3zgNIXV2HhJ4
M9yjGiKZ4s2oOkAVY+qJRanv1KqL/vY0Wp7bKrRk1W+Lx0HzKn8iVOz5Mz9+xnmU
jsuv3cReoaQ8xDjSMMuDxG+hGLyS9ok3pQqyHih+TlTsmKHxdhVNQt6Ws+FZy6am
17KjVS0k4ZhK2Q5c52ygX/qFFJo4/Jf95PIhhzJe7Wg7X6hezEShzvvFQAxUtuuu
0TypwhkDEyWdn6k3R+L7YGeW1kZ8/Wv3y86th5TukTUU1WU4IZufBiECGFhpII5t
LdQ6INwk93BLGfSei4yiQ3CrQiesNOaAqI/18N298LAskbnhSJB1a6QScY6ZJKdD
md+GTigwrorVMJKNPdGURoRONZkjAYET08OWgJcaC50eD9AGNCUSRylevSn5CZe2
OYyZ4+iaJDtkXX3S1s/XAN9LrzdF7OUc7KsD4yWlA7hJqZIT0WZHm79LRCqthQF9
asdhXH+2/BlJkMWYrjcTA1iA+iFCmClbOKV7/CNi90ztxY1CZwOiPgEbJJKnlU+o
9dAqCg/EpVG8y/eNr8zVI4s/9M9ASixwatYZU+2HJSyKHGLbkfaFkUGV0Jvn0lFc
iA9FQkYuxRfch1dhR8CYCcTugz2IssufRX62QTj4cExTkuR6nSF1+/QiCPoZWva5
OIcLr3u/YWrPWOzWem8z3MEp9Nv3zO21FtBNLNKICONeQ9nm7/s2KBhbgW4uyEas
QJf1GZ5q+rTKY2vBuCs2oiKLDM5B7/UkVe32Dzgqaf+9wqW6vbg39+8irKM5Gn1n
QFuLVEwO6PR82RwDMc3af6vx1JJlBgNaQ/2RbfN+/7jfEahZDuFf8kRc0O+N3ndw
/3YfCp7TG0YFGssBIOosDXPnx0OvOUTmV8M+68XR3tyxQfl3Iqs8/iHESIWawfKR
9C23U318DJ9fc6in6TiYkpr1xs8mDcaf73y7B+Vx1Dc=
`protect END_PROTECTED
