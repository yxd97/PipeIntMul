`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xDn4AcBNKsRwtokCifzN9OdrL1Z1t22MJFnQ2mv5wsoopS+g6bMr54815xwlObgV
2V1FVePbk1tUUs9VHszC1Y9+Xnz8Sws+5/gyny0VwGJp4SO46eu1iO5kxuFVMDhu
UeFTBGtbb6F+q+Ly5yaO45koDDtCSt4B6M+vuKQgxt2M2zxr1CJLPSo9qR2POA0K
8Y+j6kdO7J2yY/epdpVhqFt99Ily1k+TISD9oDRhd8+tqhZh07oNSwCHwc/5MPX/
raLxPfoY4tXW2/fcBUZknPfubRmCp7FnvHDLokjZl7pCdUaUm1HEc8c2mcJKKUZ6
V7krgeUOKpol7tTON81scjn15Ff2ErQynm/9AvCHMEgIXyTw/hoQonNjXXFpae02
ZWGYn1YqK6qYifGUAn+7dT+Puy9smt2EdIvmc4zfw/wZ32JDWA+E/ZWnbkX1OQJE
vQHpOBQEMXbyuKQX2YDpO5K+c3biqR50rpALDMCUjn1sxLbgmX+t2vTOeLylBxEP
mkTbGHkcOQXHG6Xk3JOntkWsz0pUx1sVclwp2KXVPE9wKFvHUTQ2+GhcoKO92q/D
FiGDkmKuaTdJgGwr02f0xX4PaRkrCmB1y+Gj+O8OkJjDn8TsJvXzlCRYmld7ooaN
Vk31lf7E+9KH8F0cBX1oUWxvyCXbK6o5ZGta+B4cvXNMsrh/pGf68hS8f+hMQ+Z0
iqnLUJWYdBQRsywNJutprvkpt16lJyROf9JSkylh/Tz1DN6Pq6AheipIkXeOxj2V
LYLZYsGCKOOla8kUCIUsVVEkKcJfhFO7yAmLkxSlGCvHeEJF1EtnIENWEyN+PwBx
jZkSF9bVYqocpgZ3noTsmxSQntOA+gGAdd+8APNrmqr6OHoC+iF1p8+qysGJFELY
hxeK2NcpnOy4+RAwKNb7TP/3fGXVHWy2MMjfsARaUcXQRih45lMhVPnanMZAjz1P
cETfIRqO1dxUVq/KH/5R5tV6MHKzur+mpaaXE7Hx0i5wBK7F3iJeE227rS7iNfmj
/vcOqA9jcAGaCRWQ7uop3pG+lMih1Y9iQfSvbUOnJ5F2pzBrj9+7qcgWNNB6khs+
JGhmV+aV1fHMB7rEQjjDcfSJ1XS+Co0V5Sw7SYdRYtBhZV1ptwfSL5uz+a1eG70n
`protect END_PROTECTED
