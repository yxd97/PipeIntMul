`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l+nepVbjR3hX+KSBNiNzT7FEWNJcBdi4vv8uvWRrj7UsHP+72nSCqzXAsLr2eMoS
NwJA1pJf8js9ymTkjEMGVBBKZ6bYLCdzzcy8hf55UUfHCwD8vAbAHkHOfeUZ0J9A
w8aS8eeMLRH/PpB7A3rIwpjFpjx0UoBbse/2FDHj2ZPRTltijKF8RJWocQEk2XMa
/ubWMAiNrqgydE0c5tXyddbJV/XWznE48tOCqqMZRiPpJfUTcYtNQMeMrmGgcTw5
1q1yXKC2aVsyLa319fDPtgtt5+DH+NVFfjE0gmwJPiPU7/6Vap5uZ0hYA5xFhU+5
C9xAXMMBFBQuhuD8Up9RgUG8sTAQ/nGxfngNyxJ3xvPfnkUOBZ8UKbpcXMQo87/p
zraog2OyGcchCcuKhULcr5AxpB/8x76RJsA6P8Jb69kqZ87zHyRAZtGySfkEHH4V
jSwCM7r+iEn12b6tVSB65reCmNgaBaRpy3VQPA0kd/8=
`protect END_PROTECTED
