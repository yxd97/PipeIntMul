`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1KusdifgE+rBeY7jGnWjxUUxwUJXYh+t2awtb3S02iMfZ/IyY2Y7YdxM6c86mlxL
Ay2waCYLR02QOvo1sFZhy1cQrPoCBH+Vz/Mk0aWvj4mYWJyeQjmH7vQsOhUyZHhr
p8RTSkVUJsAchbCL4878DM0nUGRGZCTgVTaLY6xFIfhDv+iJaZN5W5u94cYuSqDb
GtA+jTz6BFyJ0MHqzxvk4H/ZHMR9dnRVL9uCesMEKcfEzgoC0sQKFcsLgOlnm07g
OWxB0M1ZV0RR+CXzg6g5m4+3CFIVUdDnPGHR6ufrZ2X3HcadjfQ9iApNCceKEBnv
q38OFh/hUb+ovcbqaEms6g==
`protect END_PROTECTED
