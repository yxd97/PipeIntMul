`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9fmd9DrB6AW6ypbk4RjUatx+HXe4FE5JqhH2fNQxBZXkfzvyMyYxo0Ri0nz5eSf
HHMTNqcEh1U3426vH8o1ia25uXUnRQBJApcgQcsEAL5KvroAu+nebkd0w4Tv0Rtq
0fKRD+fjO3FjkE9Q00ghO34iJJSeuYT6aOWsSD3MleqDz0FotOu2qCUq5PMS0Sjg
VmQsgzEtCSqDkYooEt4+HTGCjRjO6W5Eb6pMlaPoQXeaTjmRpwGzqxjjBsv0zfK0
viA3DEo/fm30uoDgfj08lrCB/7os1OoeZFlPcruKbL9k5RvPEAD2+b/tSZhNO9p6
XzN2OJXzvCD2QHdF6gWex2VI1S7U/MVwhgO2L/+ZBr9TVdlBbWmQeULOyyDjpzm/
JHj/BhQwitdVfCMM65LTpLMwnXivgwiaGCSOO41HtivUqwEBT+S1WkN3vNgREbY/
yEER7/mKf9egH7wNkxUqFyWsD+1pjIifGCLieQ9M7o26Rf9ID7Zm8KrpXY1Kc2yN
aWqTpstBdm5NcOOJrpZlSzFK8I3sIju60uuuMUQZwmO8ckRawsZIcL4Hfn5JCIJq
obve4nNKV0Eqs9ezaUYJ7U2jvB/OZz1USDlAH/4w6RX59Y5YzGmEdw66R+LedSDU
vufDZTnBCifamxEVjhWsBuRmqgSdxEurIFkbWiirSSdtoPDboZTPcx76ArsAndJ/
9oyCATGl0Thu/CTPxf5hRk2Y/XjdGE31NdmFxAgryjajl+L6iz2lHcQQ7fEXBmUp
CzQ3pHXbPT2dOQ0ISIO7eomSES2LGXE8iqa5i3jyau6pX86d19pUDG+RMqJwEfPL
NmHrq7m/np/7mcK2GBmGUkZLJ3VQ3qdAmx+n9KdPAdp++wAicoinnX39CXlyszSl
RhXdjYIV9ye3CboC39sIkC6GEBCqvqrUbmd5mqTxQMOUdAZgmp4R3d0Q1ceCBVKQ
BJDoh2/eSvS7zElcCOAilE1a3gn758GV7yvhJwrYEqb6dpFC0DTGQEGIZgDnWbSm
5rao8nCja8Ky1CQKc0oS+p4e/0R0RDZZ31Xaz0IXvUcjVrOKibHQl6eEeoO99bHh
zjbuzWPPvvZ184/4rmeB07zZ+k8xlGhcH8yUhKTojal5xMn/Xdc9TZxL2TjHlsBe
/Fdo/0Uep8MQPe87eJ+tVMe0TDtxou5UaKMYJluQKpdlX9d1zcpi/nWY7TWxycgM
PJcH1Hb5v+UROWn2kANYU/zW2c5tjaGPxDweJRUmCHkoidRwtURvGNv6Kz9hDbcM
ODklKaWWGk5MR9ODCnu3R1IMSJWPX06TQKgUIJ/SVs0klDiaezqoceYaor/JHW4i
5h8keaJzLuF8DS9cAFaLmLFwlFExM9At/isefweXAhOlCm0WGhHZ4HJVY7NVzfev
P2xe4vKUqfV/k7gXC/hS2hi5+aUUeVMV9qcpS6ZF6JRcAaYlWv7D6+e90PaeU9zC
PGdea4rXlP7JDqkjuItJYaCd4Xny6nuKlVdW8q7p/K7KYvNK4djNOYrAVxIXVl1J
vooqsXrGJvnDF269/tPqyMU9klo+Az/aOwywam29Ofxj34NdDnQ+b3ZPnC4hT0Kv
zCn8YGmWqFI1ABYASk86ecksbQ69OOzvMlxedDFfE5uvUQvhc17hEYDskgbNoKCZ
`protect END_PROTECTED
