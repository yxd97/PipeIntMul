`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rduLMDKcuM5B81G1IeABDRccepKry/F16g3U1LrQw78MHXkxfvtCSK8S/cDWugoH
+Zo214yofvkdyxBIrNHjmj2nKQzkWUj7yoRztrcpquEXDvELu+l80Q67HHqucnIS
njZE0P4eobmoqkAR2OohZFoSGTe8EzophILGOgiPLEGCShQUVcS55lN4p/VgwMNF
LVb/nsuc+WvSmvmqp7aVlHKzRg44rPQ2054a1/NJccHDHzwPO5lxWyQ/osKfuK3E
YaNL82Qi+ZQ6Qrf29susUCC+d8TplIC57n8kOts2qLfajjkiD4YZd9AddsnOTIJA
xmnhl5FxnsMO86N2QBW+Vg==
`protect END_PROTECTED
