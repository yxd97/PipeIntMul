`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1NJSEn78DPHzZgkrN4BVV/UIb08IIZ1GVa21v1/Zub/qOnvo7AeZjGkwBeSR7GE
axK9i4K0QDbspchfcH1sfYMzlU3XC75stv6lUdc413UKyVK8bkouirIBaPIBx7o9
EkuZeH6i9ikny2HRM0vd31aPW7mEbsgnYddCSB/T4lDjFUxKgGVNes3HuefnQB5+
3kwJFKMLh3r+dhdTyH/0B9ExC5EDGOuQkarg3etKsN/5bSnEKbvEaUMy++XsxzTw
wqzpHWzHGuMGzFuIKOSIq+bMXgYjFscp1FxYR1jmzzykg/fop6Ms8kFQblObGLKR
NV+2y1jqsp7x9HIi6TLnh2YaJqW6qo7P8cI1tj8BwtiDttjgmoyaaVvEcosE6Y1M
TjwRR43l+uScBogFwmnkJSMDhv3tOdF+MW0pETXMclBYYTunNq8mHvD23oFpk4xm
S7c62X+OyNrSGTEfU4vV7hLshzCodLZiCHfq8sD8dTS12jFprp3pG37Bd6qGuXFd
h16f6aBBwuYY1YyXM1GpweKSPzPcMB+qmQy9IdnKG6DcA7je5AWOMcEEGfhU9FJw
7R06RQfR7IuVN9qORCeZEku3YY5iB2brT6PGIl2V+9OKLEdCpIuJdlsSoWS0Xcf7
IMpZjHgOsVCGE0Z5ZltCgcmovnekVXjucjDDzXTSh0/0KVkqiw8R2fH6Qwpb8MnE
z0FBy7Jyvgj+79WXp5Y4O1OOQMiqx/iibl694TeiGceJq4KnP1M/gHEciPOwZQON
hUUcap/dPf91KoUnN6RJ4ArexGzwBpMciRKbUAbzdOkRwOb6CqSMsK/rLBx3EBnc
qdAZl6F3cJe0aNYbtGPT7gX4sBTh3CMhzmUBe8CRjOYNVpqYlaysuC6tAigviSBm
10k1gaCOdWd50WieVFQTeCAcvT2OcPj4jfu4ZFWLtFvjQEQDxk8EOJ3l7GbCK98/
VuJByBeNsnWsYmXp/S98dO0413GcX8hmGJ6DilzFycT9uw5qAp/AduQOgrFVzEl1
vThxcsggqm/E1DfTervoNepfQg7ru/7PyZSYz/U6JK1/Dn89mkYgZKXF/r4k49bV
l5qHHl+WUaRpsbQcb2jOqfeMW1f2hWkxf6TVG77LfXiz7WNuk/0ZQOKeOi0wWroc
XiEcysl4G4fuYTkVnEiu0kz3y94P2A8wmG1ce0P17wcom/Q7bACBb0ig1XeOaKEm
vY1SfpzB+qFv6BFKGDdtxb60lMwxrhja5A17GxQu7YkSwFEqG8SEGIh0KeW4tRFN
XDPPurawYQjTb55f/XikuhPgDftBOonCbdwXXoKcMi38i6gPevh4SHAJ/0ZyDmN8
3mZ0GpmNWWGSSN4QFW2Xh8tAVTYE/E7MwrjX1PKKZsgqGI5T1RBJKQ0hDllAuMmE
CfHwYBLws/1uow/sx40w2YMhpVMj/EC2XsWgWC5gDDhXrPi7XTz87EEqo2HZQiTn
CQ5iVmdkvqgrsQbwgxQDGHD6bNiqHztPPRgqb9slJLyWuaVYFi0QOrJGKEENhnmv
Mp6nXrcgUy4qysyWnJqONNN2H+ZlusJOJFzBdHIMa7suqhJsqLkW42oVIkqzvqbr
NdJ01O6NTzbIMA3F37F7NKnRlrN2y6pLeOGuRKwbMoIFQgjLVSo8E1cZFxDfE3bi
CAOUwSgAYxbCaAD/jMSWY8ErPfT4J89uMf3/4WL6MR4OizNmDxkINYyryWJu4qkt
CSUlUjlIStZCr9Q2EdeuamhA/MnLLLuYXVDptBQZk8OkTA6waBoYI6KJRRa2FacV
DuYHe7G68EUo5fwmFtP/9lh/vIXdVvyawH5J3ybkYg4kUs1jAWEfeMVRHyFGz3kY
XxQPiYhW22jHYblmPPTBGZvlUyS6GZMynEiREHUr0RwZhOafhFDyiWQNkNFmql4u
fU3XLmkQd0RaTZiHeNKziRG+5QK0Esg/x9VhYzJejFOf8DgwQPuFMpKBreV4JDNV
ezDMoVQsuqb/pSV22+SnXebhAeK4E8SNiMypRJMjzj8biPwH5c9hCHekBFGNyllH
7hIoTIIUPTRmBFe/tb94ya+aWA6WKZHTMFWN5k8Hxg8IXRRDa60uJk3XcFx6WYUv
5aY3mLyRzMggMLzymN5ta/4fR8n912G9sJlTzYQLF2+qt9Lv4UctdsQ9S1TLbvAI
QF98cAgJe+qiVRfDEam8z4pd4mGhDkDfT3Egz7zuGClu1bxFqaNV3IaJwSBU4vLU
E1XV8nTPlL28UCpgwhkWF/Hd7xj9r0HvMD5Dlxg4P47rfr2yY/RG2QkCvxCDnlg3
AQTyl6LFoKMkS6OES033652G5US49R/IK3OZXPe49KsJrsK5M3CnrbpWDpopdYFE
p0csYVh0ceeCMXbiK8VhPMWm8wEauVQuFzT9vcEOobFpbNkP1RP2L79xvaFnUCuG
zabBM7MAS1HAgvEtw18iuoU9hS/o6XYhSalr7vJwfHoPHQsSCY+q9DPvFJq6vmHI
+wRiCFgpfPtSLBnHylf0qeh1GWCMmi0Hm86veU8gkkYN7APJ8YJvotdv2k3gEAA7
pCehQ7qX4snJVTq0CkMkF1LqDhrERyIPAhyyKUGTnzxNxqJFMZZHLRnZc12Jwnh1
FhQ0LiiL9AvPX95Ke6GP0p1HjNhAfyqcp3wgdU1zx53Nl6iFHpMEUCC/LvmJEwFw
Vlq+GJ549iTrCBUbqZf2+nk2uU38Wv4s0ynKimXb2/+BZClkyI5nUm2YIpJJ+lAz
1w4/fn+MoZhzMwZEUKQW7yJ4oPIfNcbEmn1mfk0x1RkBVEWuWRw37FpviDtTwYbb
jHhTyWyhJ0khCTclvxsKkinxfTsqpQu1pVYNe2l5cOOa+25VT8rDS6QfiIGEGwOr
39rDJ/yOYFi50/r7xS2XwiHMYDxPuBOikjmSd1ic9MC/zFqUligk7EctlT68Crwz
tWKEmiErAmNoouWGTzGRS+4rJqjBLSaf2UOj9VNhk4WnWn+zP59HPEeqKxqoGTlV
/tI5Ti+a1Duu9QTh1Ig0ajejih3reckZp2KSBcfQ7hE9v+uvCcSRnM7/xlf2l76Z
ECcw2vvwHQwjZTpajPC5Lg==
`protect END_PROTECTED
