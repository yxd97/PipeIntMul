`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oexVrj5hWAsmdDXmJGzIxyNBQYjuyMN9eXyowF4qfhTNXSNWJRKs88Vjn8cBnrcN
mIwySuq16RgI52MQksIhvw6kW+ZOlJXnPSQc2xAoZu8k3Awbv7ATagTtCKg3OEvU
QX8sAGkvFSbTf9Q1Yuwe0jaF5cyRpXqqtgm2onBK75AC4+MBzcKCng1MTrHUpSQm
/KVPAsrGhch32I8sSRNpd0tuhtxErnvWBCOk9vfc0XWEth0P+p5FkBE5llpbi3Sj
HbreMbEXMbX64WEOylm5hAMQHwFBJIVMm8caeh4E287XePcNL3AFtLVLivGG7nJI
K2BM9cOpKZ1coeL7tOHVdlc2C3Cjah8RuZlnxknGRwsmBsRAq4vq3t6qfqPAQa5V
owSV9LUVeTzamXQPiEh+vwkXzQMCHCwRs6xDveR7VVc=
`protect END_PROTECTED
