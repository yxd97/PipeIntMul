`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yP7cvcQLQuxO2UdcLOwjShRLgnHemT/MAVnbL6Eu+uHDC2JmZ+V6huTi5aoP9Qlu
4W5D39PAjnl9JiUDRpASJQRHDLUdZklAJWnsykcFOWZVwDZGvpQu6rgVVgA98PBh
aOkhe8UigcqL3WGGMWq6HXXDuc+l4TrEyLe+9fc0MH6sKwL27X9xQwBU/uwR0jsB
OWzWoU/fOhBrjPJw5neArR/JhftqUBxGHcsn7R5wRT5ehEn13O1Hos6w4vWcKhiq
ZAqnvUmJGKCqP23DzIlipo3BpFNMfgrDBf8MllVcb70x2BQNkVN2vlMIir9/2BKA
iEZLzu20FW/7kBLvJhIx753cGQTKwLoo03YAGECJibkPw/ZKVwQDTQXlPDiS3WkT
otasLjgni6/LsZDLohg2r+UTjYK73vDnJKZ3WpcSbs4Q36Of8G5qPQX6SpHUBqEY
/2bikIvn0dJ4ki0O6Qd9WKUIVSEaWzEfpxWQYnYBp64P0Sk74wwj20jCLL+x3f0b
B17XMD7tkSk/rXXixAE9quu6tSFKaJTjlUpBFAuSJDyprPOMBRKzZMQMSe1vZFuc
hJG0FDbpRLlqvpDQAueOMI4+7VyHKUrnu8b42hTVAjCmi5BmeYdeGPH06WCs2oKg
WVu+NhEaTSS7UQbKLUCNVa8ff0RV1t3DBbt859mQ8wlh55UknlL7gTdCmV7vY1lQ
Mp5BLSEmebgfQLnqXjaY7o7gwZQZqwfRJD70jvdPhBIAdZRxK6IdaWsIPKXWv4Ah
BgHNpZJUWHdn5ImyEeCBgUi3U3V8sG5zSkXV/7fdgOZ1HFZolHOLF6hRwtR+I2vP
Z5D8VsECcEVuvt9UQD6vh+ZXkEVkW+E8BL0VqaazwsLiugEpi3uczOT1hwzj5pWQ
gvUo22OV6m8T6Z5zASk9bsSOt0oor39YTj15ddUVg8wNoYxmNOUrDr80zPjV2wfH
zgvCr4BAHHLbaN0KwLFgoTs1AH4yrEV9gr3+J3H1bPwwDsGEE3XU5iY2rX+31zjF
N6Gv0SJupRPompBkzLm9X/mQrMe8RWC54RDFPgtTrHQ=
`protect END_PROTECTED
