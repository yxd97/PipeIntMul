`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UlSrf0yjzgc63/vpEKf0WxTzPkzl2fe4T936DUG3MGesI2h8VpCijqb1JwBtCtKj
Ddyqh8LAyw0n17z1vYz69B5EJT+q5X3U0ZK78+lldeph1iRYO2P7o6KeXCtIVJxm
a3k63aFOK6Km3/HoOjJ69NF5b7nFYvQdT62lWDIAtho2Vwn8W9YHWOyp0LykoLXy
E4hrUFIcblxLSmSS/JPzR9ouFDZ8VPKRD7qhbC24me2jSU6xoNO2U1THKb97ZSvf
JvzDD9TQmf4IZbeXq6DLc64/CCmPIAeGHOjgAsKO9RKMg/dr4LksRewvX0/eMJCn
pCfbs9buzL33fEpCY/oL9hn1qWHuubKCLPARAbuoN6ti/YldY2JylEOqhmx6LIfk
tj2O+xZAboloiLKnPtA4E6UaaUf2HWNIFWpji3TVpaZKYaT2b1Wmq0mH3QQmuaPx
tIt/A2g5gAYhH1ChgVXKkreSPoiW84p2Z6VnjvbC6ZzgxFRjh5hb+aCpj1laZxSG
QrzPX+KdAEndzWnRKUo0Xg==
`protect END_PROTECTED
