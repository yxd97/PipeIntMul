`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DD9qI4y0LdZNnU5VRekwA40OP9sQgFmdSyPJEcrfLQl/u0xVU8/AVdK7deG13XSr
JLjXgooCLgF7UYincjKOrviCqTMvIXksOdTaxASFheRbEoXWWkXY/MFcSY5H7FBz
4kNBcuk7E0ePtJronLQJgvu3kFrSM3NQnzhoKouVorQpRcGWEnmqNSTfWLhcwDv9
ibo9ouq73jdwSBDA3XNd19EOqklN5GzHrydapnqxGUiCOH4AAmu7LXHLrysHG6fe
6jSMAfUDDIa4xePOWkRWSCXtmQn3l+qERggR/4a+3/gBFcBBxtxv4KkOrP2Vroe3
cNamVnN2nsEpjSvrEK2K9vsTlSxwzPlWRKE/OkUQjMM6kdC7tQqJv1SwfOsVds9d
DmMKHd/TPcYCS1yfA6z6dwmJngKZgaNFIhoZMVa5Rkij141RBooIW+Jn7ZQLEZ+z
xRqL2+XjsTzMVdy3H6XSNHk9xeNr/DzKbS/DVmBm2jI=
`protect END_PROTECTED
