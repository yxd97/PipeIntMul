`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K4wNP8fSDVKUns+y9mQ2RVyt35ewimCvRj34cgFBioZxaaTK4Sku9ueSCJv6nU18
JIjQpvX4rjUwYTd55OAj27D8gMA6MwxVHny2/93LLkK+ktbZ5AT1yJku09HgwcIx
HdSWkMpOT8YvC7WALUQLOegA6buH/8776YZoo1QiqhqNMSPQoNw3nS3+riKtK4WP
dw8xpYmWazy1MA2A51IKYpnbwvC5PNovxRLb7iioYiAK0C3CW5sPWKMiWYr9G6j7
kG8qe0EKiC+YHfSf4Vrf6NxY+7CsN4JbZLfNxShlpDaH46N1e39UTI8Rx/j8B3G1
o+pBiQiLRipu7QwuzwLldw+jJv8vcnFl3m5i8+owWin+GGUNYboJTFlI0da7sDxa
JYyj8wYqkCPpKTzUtTzXrHaGzHKVeDrKjyZLNOoVxFrQ03HQRqhL7aCnjnpB8GNZ
BXTE6oLncvAl/32gqk+cBqhZDDSr75uVcX7WCfy+nJYtduKZ+7qJGiTWVr0HTerC
yCOm0TyLnv1sbITWZMFS4XgSBJkInhjj+9QQBWgb7EA3yj1u00oQTphNAMX3SoHE
TXznRN2a3dUlDdBHg65wGo8Jbl+2e/dRIRboFIll47b4iGMcwIe/8IrPq1rve4yO
BfWuqcYa/aRkWQ+lLPUvCUm9m5H9HTztBWXRAO9GGb/r8FEOeQW4pcinwB3KYuvU
ly1mWm+WDDq0Wfe9wgZAt7IFY537KJSP0BQ8/aBWxls/UuwCDFKqjtdUM2omKCb0
Pv7NwxN9EFMXcc+k0eSlCAb0z8ivFyDw1Eu8Q/ALaR3+pVzPpRGyvdg4R3rID3l0
feEI3wvGF+uKEPwln7nVFYWhSSnzIEY5Pz8/K6b42st5Qmmk45YmXmso0ToZl+13
QF95OdC7QaA8qOHCAfsLAQ==
`protect END_PROTECTED
