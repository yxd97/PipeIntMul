`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iaaJSlWkjTOX7mCs/yPdCL0fFknh8jm4NCGs+ihoEfbJbTrF13SgZmgdxPlPKSpV
egGZMMqprEvI2wuR/uIZCpA1zVHLy/9dxV3L4FxhSHqb9+0JO5RQBMO10DUfGtKr
DQfCZEaHGhOQq+MvTmGSpGEn8IEDJM+Rp2AZvjgnfuGgIrxJfoYLTQkrJm96z3eS
2zNF/TBD1/q8tgE7U5hN7+4fK9c7MEVn63Ype4uwhoMm81QoK+qNschbjWr+pn6H
A3mjNnrZgx0IE1DeADb3rmB4gircGN3p+MNjQyvmfwMVKiX3sYMKvwzdYd2BWzBW
j1KIclZ/K74tLWTLQhfPo9wv4kebs+CD2FtlJPLSLkKs/Papo7k751GejoZArfj3
efg08Pgo3kT8eeKmGnIqrqBUiHqiHyz7oPe7LimgNffukpZUaPYekzIedFaVRHWX
cIpnUz1ABH3rAHvaN+baTXObNUO/WEc+3PuRtHjLABxtgDrWw6YScYeil5Qrl2de
kSn3NGd0tCkVI550nwXhfzV92yN9WqbiqrDK7hANyFqkBw262FC3HERgfrop2y2W
2b7DiEGjuyETo7oSkYt7TfMZCWVCw2SkMq44mzMzpolXK31/mPPIchnnngYK3dkx
I1ihYBaqFFPZx6OLYWQ7Ir0k5BHcihHBwdGTueTkeIOooeNBxnBWGEblAyVrUPod
MIH0rLGX5XllKZzV9/De0bmdDaEM2Qv9lhGRqFiCLAiENT8nsw3v9aUnfmBtLH45
PECTev8pMzy45ptHg53F6015vHEKzzcx8N3+i2eoHBy57bYnirQiBg2NIYuB3G/C
TTgCUUHYU2U6aL1oRS0RyWb3Tx/TuUYwYfiRD94Dgfoux0UBE1oBANS9TSAS4TkD
BZQMnwTLtGY72zNYx7p1fQ==
`protect END_PROTECTED
