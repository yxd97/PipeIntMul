`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQ2oSgyX0vt/55ryI/zRBUbB6yOn/PLbfAPYbRvlJtl5fAR+gmnRw9Uowxfyh+M+
2xOqWJ3vnRa1E90EDFHDRjXpgPkPxYKXOtYuaz0NfGHegqJ+PnEHcehzEARFIRu4
ZGJ7FhZD+cUF4XiSiJjQGgppyv/6Ym5wVNc7EJcO1ONRVWRPi1adSAVDFMAnyCEy
rYmQWyx5ohHtts1NvHy2ABzkOeGIlATs29eCXTR1se39vDIj8LGa2xuOxZ8rz6AZ
pt5aFhe3pcdvH49sH0Wu1A9mbs+PheAvnhmasMUt38f+yS/XOioOunoO9MsIOsmX
9K2rIaZNmvz+OUippEZ7t9fAoQYyuZcf5ANF0G5f2SDTvoq8lhLpHW6SIe8v0Dbw
36ueKxDJ3cdTuny7pXwZKlA9cw9+UoHufdI2taif1Gg=
`protect END_PROTECTED
