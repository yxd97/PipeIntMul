`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9pkFSRvYUCzI58ANMgreTJzoCMH+D56Pw8/W89b9hmjTkmUVaCtVTpV1WVv+WcRX
HJ42AWoLmJXtCpwjLadlz2WT+xu6wy237P5wmOdU28PB74S1wjf053Cd6WOo4O8G
dPXZ8WUO1Ni5MgJ+K4uJz0UZUfuOsXswuM7v4ksYTdbeVyLyyxDumPWSEPeskc3H
W1wxPtwEuEe9pYdGedhgAioA0ru37q0Aszc6p2EnyaPpX7GjK2usGZEMrItozAzR
pkYJV0lQLzmCNlYOxxv+E0Y77VKcaJcXFe+5avpoi3V6v9QmU0rUZn2GfdS1B5bk
iR7mC3gg86+hwceGFfQ2HfGEm8jtrQDNVk3Ca1BimnvnBw/HOOt7datdoAUBjh2J
xbh3Irk0gJgpNPBEhOTeFyNtT6B+8tUPuDixayFhlasRSOGbJ1/PBrtqJE0iw/WZ
ysgCQEL1f6uO6L87XhRs9zbjbgtNY8BcZDytvkoKaueWQ6A8JtvppFOWZZh80agq
`protect END_PROTECTED
