`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Rwwud9dZ+tku/9Uvy/elDJDozJz4pnjy32fFORDmStA/E/eu93lJgUtcJ3QPLMn
JSxuB2KNqOLT9SvIb5Tm8tFgei4Karry1TBcn3vUqCsjFjETzC4ieJsA5Dq07OG8
TBjAOdB90C8Fv/JWsgBHAYhSec8mhSaDGL/mGdHbtRmSVYd4JuQjITzzHDDUcdxp
28h7J/2Mdg0aiYXXFWH2bUmR+QRQHpRJ9Z/xRLcXswrrZ5HH40ojWIawVVSO1ICO
ZqWkN3Z8gUfTlcNBFqXSGjVrFq9ED2hHSJWMmFfE1tzjY7HRHdFNBXyumObcuJZM
EfKGcSdyqYAPGHlqTN4FKpPmeh2sPQVo1vUdAi9TYxEXCqLWT73ikradGAGJF7tN
6Y+C3NR6h1o7uf1sGVKsYOXHW6shQXu4FhTfWvt9wFhu2/mRommVXoPh+FJ2/a7t
P0bwNQVUYVM+bWuTGhabUlOlusoHXRocW/r+oEHdXdp/xkP8vHlkg/q6PPmVatg9
ufewhwb6jCtxhqApZzzZOs0heMG5bfrhi/1wKzjUv4DYlb0cne79lre7/rPhiuO3
MLmPvEWPJE3joR/TrArvmtgiGqmzO5+PMWd2QYVkO3o8sAf4CLRTj+XVFTWsAiCl
erzBUG9V3ozsjHvawbZI7A==
`protect END_PROTECTED
