`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YFLHIWcsIU1R0Sc9NBx27L52DTBtumgOCrJoOB7VxpVqF8/AQHATkFMJrBmeQKUC
YmtT3i/zmjh1gHAkGWg5ep9YcENzV64u08ri7JBFMbp7KiF3uqaX4lKv+0mEtXw+
t8b5QART3ygTMW4LdfPFdhp50IXLSq5LKW68Ngouh49slD8shEDC7aSZG2zEg3uN
tOs2pFGIYr6YB8MWcXSgJ7MhCEa0nDdAMDkBj0mIIbLWtf2LQTttJxAWYOSSVnso
/+3C0QdSU2o+fviDzeCWclIECnoeH9pYD6eO2VL7ajM=
`protect END_PROTECTED
