`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
scdUVlci2XkRQ5dR56ild9K/XNfi0OQgTEbnDAFwUtXOwewo7DMLoy8ZjYn5o1RT
3YQksLD9x6Eee4QzL5AaEZzpGEUOehNcNGjj44ckJpCc+41CerpYrSiJHb6BTm4g
Avstq2f6UUnFtUmpCRoXMY1nzmPOXDmLeJR57A1HXM/pCsqjmLIVCLyCO4ixpnsE
hY3N7PnBtLgUaYlhBJl24VB4I7p6EuDZleV4p4zf4NEY2jobWhm3gFaZK9pwgCgz
Q3MS+4y3BTFCG50l+E33RG1lm18cS7hnA+xTIi4QFdkepCVD9Weh1TX3aqjAiEAz
Q4j2Tqkm0jY49fmX3Xz1cWDfzhnvujG2JdY7+G+IxIDQ3f1tf4LhtsWS5KF0J7z0
PkE50n5zlnlbx69fKpgMfOcWk+9OgmQJcPyEnGsQgvK2Azvk0jOv96Rgav4BTdzW
rnNpaEdKRx+ecXfoiKZlRV4fP8nRxlxGHvleeu2mPNF0CNDIHRQQwbKXDFzFqbdR
hXZbDO3GV1NEcskTFQRKpAQGZVA5k+luTe6YiRR7HBxR4L3EbAwdrETHUsZ/5SFd
H3GcMLk1mqZYXbagejrsijYVK+GI/THVh83i9BOg2JjkRI+655rt1eArhuoQF8JV
QpgK+XphRm++ZObfmnPRDA==
`protect END_PROTECTED
