`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dF5Btoi7iL72WT+CsEDQP1rj8NDO7r0H7TeUFsFAdS+4gNXHqBQ7o4gfX2ZGttpg
JgS9l92sXZwjShCzapCfsywhDuQkuvIhvHlBbX7R7+RlYRPjErI2OtGb+exioWKH
HByHtITBMkSOcseuDBie0elA7hpMaJmLPVKb8t05Y7Dok0rniWjyRnUVdmQ725SK
0a74Mx1jTotwSUSaw7Bf9HOYuhJaRFy4OzICKtI76vkNak8Cn6twMuB4Ed+c6qUX
DAdOL7OiwkguEpiY2UAUrXEj4ssOZejj4ooZbKqybl8Loo34LUf96S/a5a4aMall
AcQrEUeIMmNfSYS2XB/N/xU2b5VjtYksdwDPwUl6zqxJYk3ukzNCRcAWipeCFY5Y
s22SfsYBoS7PlVadf58yu4WtakSl/QEjy0ifA9iBqgZcDVQDC5sEWgefeAthm2S0
sWGwQ0BE8KpFpuaxUDkr60mchFO85dA83DyIs5Obrk/FDQ7W8ErPV9wAumYInUDx
Alr6QV6pz7yL9C1i+r3sVoFYrW0vajxSZZS22zIvAXRhZcBc8VinWvHghti8rJU1
q47ps3/Nwc/vD+ZxLimMMwD8bV1vl8faj06BAvQLWnR1aBI+NjRz6Api32ZFlt3V
zyQx2EznRveLE/8tTex3c4bu0Th8oPubnx2m0ecJFsPCpiL57Lgk5gLPvcvgdg/c
CgESh2obACqc2gfUmhvgwhwK9IGr1tOx4mUQ6ReIpNAEPfwxiQd4lZgNZZ87/soB
9/3rGomZKgTCNScJn+zBilugC03zNVsgGxWIBOI+9wNudLLOyHWXYOiINymo+I3c
NYNAwNPSyqoUNnP/TxXY9HfEkEf3gE5pt97iQPyyYpIIOnuRAB81IDAHOszUrLHe
hh+DPgOHObTDZ7qAW703R5pMV8LECBlOfM8KuLMNowuscmSE0EtpRA5x5YRDl19x
Yof9yAx1c76ImKF96J1+n+PBEO9i3PVu/Ls1oospBFbLixkf5u1m097eFI+YqJw0
/FRHVR9oQBXQBazDVoTwP5fOlJaIN5n4w1VG4A5BSG9ksz/d56V4YNUOwYOkbCpS
TXTomzOIs6Bi0lb8BoLRCnS6E4GdepT6qBZnWKtcrFckX+4pY3WMvn3M3dqnqTsm
WFeJ544WpTmRhU6UEyWf42n81mlBDLmIqLJFIzIWYhqpcNYsLd+ieAPyPX5qQp3g
qllL16oSsEqqhHuWqrd9pE60+AZQIocgenVFCjAmDq14PVRav7mirTr1Fft1bTrP
d3OL4HSJKlwq8Ka+DO0lDCEwXMrJYuoCjh4nhsiRxW3oHA25eG+my5vSj0NccbQH
T7w4A8DiKjXZTigk6wtBhllwNg1tXT58ITZPwM+uD/k9u0Nho4jHvNca6Uys2wuF
ehBzfT6fCyyHbuoWw/vq8fZJjbvzul6O6vlARt4jvTXyYizTgP5/UNDggfvFg5Xa
m389Tyu37s7y+0mLIwIwmSfl9rHmEEHMFE5ddSFaWxu4Bt9TALuYUE21sTB5yogL
0Ze4GUsi4I7lex1ApcXuy6NElu5x6qjIu/cjGdk0Syd8VcphZfCFZSPkmMuz/B2w
IYGONW7nwM+0FqSDGdQeqUGmYvAxk1nyxjFCcvd8IyxhTzKaTqM3AQy/ETsPqrO8
jUVyLo6uUP1yNKm1GoHYncdIMr4QrIOZte2GRAf1G3wQB7SX8O+8/yr5oJ1xi7Gl
bfXtvwmKmfg4OmsmY/YZniEBh/emVIsgoMO49BAdwnRN0qm7/8dgBoSKuNEW6QTa
LazsL1l1oPpQnXI0K9T7UJwAUCYR6619PczxMIS9A+Fe6rNKx9XuTwTAlbD73LQC
vhUTjfFuPVJl7eMPQTixiXYNUFt25P+8xURsZ3DKRzAxWKRoHcgDlB2pdDj4/Sw3
Go2ZfdjnS9t8SwVJyFqo6z+pDVdPrrV+F5s4kX5L6X6uQAF5MCSktblW4y4rhNc7
1IbfNEMZItxD0ron7dxFdQ7JkNGpRz099zb1PXVwX5FRpUGIyAnj3rmrHPEFtfx8
dSedYKfjbVPbzxv+xFC2PVV3950+B9OBKH12u/SsI7HbAa8V9lv+kNa4dn/8N3EF
rJD4BakRB773aWLPgC8HuQ6ConLxfPObwF8A13Tucrusf8DLO64tUsc4x00NqwuZ
uwlwL+homcVhg97SecWKtsfg3x373rKNVUmlMzj5MsIyCHnIHcxVhHf5UESqWyz+
87T4A7G1MgntJcPkDbA2/gSMgdFdFErxZBK/GxH8qJjIl2G7pySSQm2sxiMzKcwA
6Nu9CbVVXA8KPzXVt4AX0/Wb8pk/OUn6/YmZnvB2xXEioMS/XaDrcNZQi+zi0edk
POxEKyMWeIw9T5IbGoUsoMDt/8qUhYGnUaDS9GNwnDcwKcI0wt4zYUnKKJUk7m2t
SXJVKfsDhi87+FuUwrTpZomcuF8xiUjLTKbxZM+VkViYgGdZE1vOu1kBOYOooO1U
w6dUE75+Ul+8aYIEpUHAp5F8NhHeMxAdqXR4v2/dUSKmTFDjTnbBH+Pyofvtnp8Q
BU4vzv463ou1qE30Jbqg3wNZwd2e1Z0eaQNRM6Y6hV9FG6VyParqhxGDlc7m9cZk
lhjUl3W1wDccF1xVn4eKqJPxpVBtIg+OoBJJ608xLK6ov3BSV4avcchRWMuxx8XM
hLg0YgKuTb+rXHCuBPbI/2UmBu2IJG/St3aWEJwgQoTS01ODzjZouW2DbUC7y2ba
mOgcZzlnR93Q2yAw4olFWr7XAEf405xDXlzjB/ed+3jdDLniF+q3t/tHbG696GfL
LCoSQG0eFIR/KRSuMD6moSGsg94GoKKgq+uRLWbqTKNyHnYWQuZVHity4GQDxV1c
fMOiltGz+27FytuKK70dD0D+y5C0sjYROHMmgivSGF4E3W6RmXW2bpKItLt9Tcvo
NHVP2ViQ72EYcJ8DuB4r/oeNJeURE60n4gkQLqnQpKGtd78XhE8uCQaXi2LEMbnB
X0CKftKVNa64lbYmIXfyr+kbTIPIvc+XEzUu2Ut5tVMa+fW5vhoHPpybO/rfkWmE
ilsSciu2cCgpyBBn5Zw9x6SxsvhSgVFrjBrrmim9d1TpTi1eJvCPcnEDNaRd+5uI
M2Rsi2udeYmjE+WprfBnoBWBn5qH+cbsrIvDBK2LSk1kFP+60E83wdpMcMtgZTvK
7N7c4rYNU4vP2Wj//biVAqce5u8fzLBWK0YwU0XPb7mgqOzNPFvz44J3qCH/3Pix
xrFo72Odmm1rbWsRGf7r3+ghJaBYiVt/aBdnI9trZR7eN8ohS/lYP2DPw7/CTHP8
f+fNVynFRHodJoqeNMT2wg==
`protect END_PROTECTED
