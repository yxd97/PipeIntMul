`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RfLKOcjfR/LacTXBlEt5CjOcxeYfwiM1dObvnMPGRx3Xkt+/0COOKMyNpmP8YLUH
chM9B0lwNUq+k2CpL8fsbdBB2Ry6aQskeMYZhCoHTjm/4yD3cnW9/hm79tLRN5jx
KfPa2mqJ4hMKR+E23JNZHVafBoIwpkwgJw5RdQxKOL0NBNi4NrcVT67GNiXpA7YW
OMvwI5sRAqlx91zGC8PnZ4dxqmdH2+8Qqxz8zcOyY92xynGiS2JfzQUEBftfn/os
KApA4uLAyaPV/z2MYbziUQ==
`protect END_PROTECTED
