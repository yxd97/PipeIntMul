`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8EET2jLKKG78a5gZehZLB3UaLvmgmC1FwqxIJN+2ptouENhuRT2pHB+84PX8C/6
owTHckPpXRMdcv/iVvqRIaJ3Y8RCqWWO8ovtuP2vROvLZCUBOlnoZgrRivWY0NHv
ASLBROMDs7u8eMq0/MSsvfRlVIKWF1hc/juUky6M0AFmnlTmmRTwKhuBABj83XJH
MoqJu6bSogCquNR2bn0E8RdjN9ZiVggECubn4pd7ksrpS7HL6LChYpcJpGPdWRTd
otiGFdk23gv04cIgHYdk9ME85F5KiIAga9uPy9GTdK0WG5ktfJRlf0bURbgw+XGr
Id61cLflLfm1Q1Ha8nBiZbLelTr9Qj3ky50d/XJF24yARqtxh/xvmaFRm2aHBxkw
1W6MosjtjZIxuKHu2TGv9GB08c3AIhT7jyJ8DjhcjC/SxNQnsnJP9PRPwiWdyuGh
AmFiC7Qd3YroTQB6H2GngbhuwcbGVCLhb98J3u1Sv4b4FY+an067T/jehLGDG4U1
S+/QTnzonX7aFifpIGcMu/UPcnvd3m3bHqyH0wKekmitnmz8WAFSuL6gZ4fhJoGe
uQB5tXitJ6zyjuKpBBDZvN9g5Tz04F5nix8GffmhODuuhMZgGrW5pkc+jML09VeG
Ad0KNWCtSwCJJnT7Iz4qothzicKN/CglGvhLzjNbHoylbOMNjOESDfPN3diUvvfc
4FpH/+OPVC14zjJA41lpI3tFLfKDrggSqvOdH6DIUCtD5S4ZnnYnzPzMwI+Ri6ZR
Ia2NS81DcZZpSDkDXMkbwEdgr91jpTeyLxQuHCuVgMYNk/EwVxiRd/yiM+AX4mFp
YaCF/fLWERj2caYvlJE9EeiSIlfds/zGECYhqe1Z42OjTzbzfoXbF9xYkdbEAXOz
hSg56JT+/PRNxH+xTlNJEZVevEa+FukmsdmB1xyL6MOtXF6eC4t6e8EV6Gj+0vxH
Y5sAl+LGg+9Eo64FjjewB18SOUitbargVPjJw4pfLYfCG2SC9HaSX9XtXBnvXkO0
6VNbv+QIyDIXBRV12iwcvW03KscogaaYvValQdSQtiGHhLmU9PQtDOwsPKC6feS5
LjJqUGllxjcMqze62mePAPVhhrg/raZ8Q32+b250+bUdfYxKtAEc3TBH6kluta4b
I4rWhYR4T2AigdSQ+e2OjWzsWpACh8gqk6UDFbNi26Y+ghdLHoX2b52mCQ0PkgNE
0296O1etBTh64cVeEQTl0IaJ0SEbuGLc4P4VlFd6wDu4QA3ia00xUCWicUyGEhAQ
H4LyDzysPFb9em6ccX/hIj7SpxUpEo+fc/XJXGezR212t4Tx4RKn4j81UDV+71yG
qxxGNF135CrZkjIrda+NJg==
`protect END_PROTECTED
