`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
twQoUNZY4exPannM5uEJ1kKU1QoyBkzumMNznvkt7Ep3Orurd5y6owNAU+0dNcpU
ePNNYGgH5LLa//3LVMJ7mRiTzDBivly9a+NzqkWIFj+916wH7iVkNuT+v4/K1JYG
Yh4yolxzaknRWPD457FNEnEUPwzWT5dxlpE70TyRMcUR5tOC5ZtgAMH19xVMZh9a
5X+4fqRVZYCYNkmIZtUodrzltFntBo3rqXCFTWI2Xe97IFCALAUtDDL0VCa9UzEt
hjHwsgi3lY+C7aG51odoRAOUcnx1zpIyb9AAUZf4//LEGMQgOdukbZaMej29eucq
aGOifGvKqUmBgKx4sjDQS7hu9FW2b+ro31gVsMvI582Pw2y7Ck1A1yTy2TXC++Bf
Ra2zmuTZrKRM9Xm0045T5/lYQdf3tqGqZVYckrqeOLWDSzWwyOGzYGzL62Plv/8v
yUvarMhdX9Eofcl4SZfYsB+72n302yXqhPHsTs5klwcNsQ/n6Z7BBe9z6VaQtx8K
v4byhKjMuEC4evCNBx+GPg==
`protect END_PROTECTED
