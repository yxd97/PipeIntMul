`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ggdXWgnnBzB+7bwMH9lYNv9g7s0rLLwU6DMZOZrzbPerxhB6hkygsG8UPqX4DFzz
I1Mv15f57kXZB9cpO5uhUfj62LYYNADfg5XML2qY6+9vnpcWCksQucTlroMOEv7Y
N/JNy4Dn1JUvchxnEcWC5r3QhrsfaHiCgOZR0r9Ffk5dQSj4Zfc1h3LSRphKQGZE
fD+dAYo1701xdrfeKMr/ixcD/hG4kctOPiK4O6pSrjGGvuNEs2ayHOGAEkdJL+5S
watLm3jCfmg8ib70uDolWTNHaRfpQ+h459mFx+FBj+MGlgg5dfwGVlwDF9uTDS2o
M4KUaFYS4MGNUTSdh61Nnj+o/Xf/o5KOQTvs1JR14r2sXmD8FEQZ5TvZlBqAoWmm
gHXNVtMZnftl9Heu8rmv8VD06Gu0amlt1eYR7b4S3xTQv5AW+iTcUmgGQUkg0P7n
GkPUqnFTmMyPa+hbC+ox8DyJVE3Dm/BK925F92KzsZ07wyl0YmteUXzi+/zsBk7X
nTlgfBlbZepdQ1eLllHda4QWkr0M6YCjo6azWpIUa1cMGzaZW8/fcsUybGuUnFAY
oWS4UxFRvlCxVqAxc9gEZkHbhj39ie7F1Re1cnPHq1MxVWAK4/aJHWKX1k9Gon5Z
zkQWnFMePzwmOr/zmZHoxxDnvAL3UbV+4n7NcLBF0rDz9ga788fBOEDpb5GdeB4f
QyJaB71ckfaqDfwr1fawnCdW1NttHRX6lCGOhZxiLyjSpnOVDgflZls0vTeoXKen
K+DujJQBDB7Mwp19TMvx/9w2DVhuR89BECXjYl/+tuUeqJclfZZ09DXNh1jmsI5q
E2WfCjyyiUVertkyN/6v0A3j0ifjXKkdjwo4SQPKShq4LpyVEXIAAj6OI2ZT/SDY
/wIsQA/zFTg8Ozp4eL/xhrbYbZ6d20wWIsLrbwIrBUmn00n2VG870QHFzlZgl9Ez
cw+UA6FIdMMoSBenx7X7vQ74NwL/qclBoEKabbPpV6zLu0OyioJPT4qhc+6iFi2p
rWImyrUYW8HEEU/5Yr8ZuW7Nk4WUKfqrHqcekotmIRIhoeH9YXs4r6wt3aThtQku
GriZZ+VGnjlhEMuA0B887oKkHkUcBEebM63LN1U5erJp2GkBey9k6rYbCwgSDCVD
8Im6GIrPLyApyb3RLukjdMDIrCj/OqXG0iFCYwBeeUVZRZwegbFq5WHMJz6tCIbc
zD6dm3Bp0U9/pd+NA74RhdZARVcfQJGzCvsPLoeBALw965yh0Py2/fj9oplCX3Fu
x+hwxezvDVUGKC+wor4YSzU0qsqtE8Q396eu1CzNyEpI4TY4MNwAfe0M5fwkMfIA
rBmcFx4ZVwCt1SIujIu7zZSyAYMZlJOZdV4ws7TlTD8QFJNOMCtmErHMAjIiyX9o
Pn2YLvuatKvxOkiM8TpVwxSwh9b+ol+4623gAJR1bbfYeBV0BB9iC4+CRTuylGW2
D8M1xCSfubPczfRxp84wq/opeLSUXxmsM6Z+uR6B7uxxIPY5C/mZwcWTNeu4M9Lo
ovkQMdrnLuO36WofZtI1SxGfImjGSjzMrymKRurwFIKH5mWSWbpRHMhoyWyBFDo8
omsOrPJMVho18Y0GkQ6XfCxa5bX+54BimBdKoiQs6ulOZ3HaCTJLKXMl8IU9THhN
nR9XbiBTyzgE0JzyixcQJY9wNOurmYdW6Q5/m04Pd+W+B5m4KPWqLVC0suelDjZk
gbBU8pbn2+NcOXCrTQHo+ZmbJy0k554vUJ6F8Jk/3P7QWJHcKThc2y7ThxiEbrbY
mMZxt3jQZHxOTcXxgM4kvBHjcHbQUOeGhH4uKCMQIG+nj+GGj/+R8u0HSeGK9MBT
Ivr8abK+Dz+1rD1vjy7IW5l5X/D0ZWuN1yHGz7EY/Rmg+JeefUbFwee6WstglujR
/eTL8XYXBkGpGPNN9NuR7+YZZy/VxafNSGEfGCQWZtYFDO2X6BuSqMSIvW9edvNS
sttMG0zkgPImT3X7rzqN7Rw1ppzZEmY+vTSYLsEFaiwbUp+w7olDGsyAmIr9RfOx
nGufU33faBQfKcQPXVmbzp2Ixn15oE6ut4fXoVVpjWLfJH/tJsYHJnqDGTYPg4hm
ulI0fTfjBmZ89QLxdqEfXjQssP/Yoa6kZkMfQ+GKKFK2WiP04Ojd03K8c+1PDdoH
TN2ZJ3qjYmVsQfPqcbtlZeug2RFGqvKTB9UGW8omRcEXZ4G/zwC656G9kvVYwkVK
D0ox4sb4PpjLuzyqKZ2a26ly4ZTkomgsCAa6UKtshaPCB4FsjgIzaLT5QRtG9R35
QQmfvxKb2ydhBEra6N0DXQ4ndLvc6f3PTTJkylZwg5cjFyFdBGFgk4KyuFFhiWmx
8f6lCDQZCM3MG5bvEFp/n56z/ehkQ0nQ2MEfoa8tCv5sPkgJQs3xy5ufmjXtnVE0
jYxjh72Lu3kcFINFDU/5uwoq/FLqrfqK9dSPdG85Bb371bh/6eyfhHZxOg/fUFxa
L1lIgR0u6THF4TSEVVlBe5mZP5M5fp5bxncvGQmHPWwBMF/yFWriuq+w5C5x+4wk
drKLVPsKcoVhFgKk25CW+WbIyn5cYnSj16/widCWRSJtLm4G5XAtcxb4tOz8qah/
gwb/rmNsxngP88HYrNFNuzgf16x8yyHnK0SVPq1v73TfjyLZbvC3wLgKyGsSUClE
C0lbaoFFbd6PEuIEdm/9+vDTpe7v95VeNby4KFWyqHVizMiW+Z/KrmD7ggK7zSL2
GO84loXp2T1UlkxnsNbunpVZFz0RDgisGvaCciOszuF+W0GYRbDpa3yhm8c2gkTI
Qs0O2VDiRLQp5+M4mKdIHg4IcTB2fWFl8A7I09IS4T/KrcTqyDZSbWfrBSd/soPc
5GcGgmgvGiitr2kgDAcROqDS4KJiXMGyxg1L2WRQqL1Rk89t7eP510PViAMAYgUy
EZb171Ta7HMWcJAckjTdl5gHT1SoC+NNJeJ5DL+G55kSKkomL9Zcn0+iDNIkJh1L
z4ANckMWVBNmejmnD/PtemRumM+m11az/pn99rmW0y7CGrtpHyYJKVFj2FNNKVhU
Qp/zTTCi350jvkuqG+++G5/mTFZ7oGwGRgv5b4SIVcjDuIrhmi57G5kHxqjOYjbT
fIUlhcPFT/+MUKC4MSfPZHm7Br3JCdgxA6fH1a7miK4twffmPxzbw8/f6lPNO7qr
kuJsjDFvGL9h7acOcnEZ+tYQJ3oQcAHhBnV3Bc9gLrTRb1Vz4qOZ7VlWMDaJjFpJ
MsVysbN6N9VXUFkV2MWunAyQvQojQdgm/aZy1RS8dIYGZTUdAvfe3NlTloudRG1Q
VYNet831riyRUVRUNTjN1qmJ9IdgXVIgkd6spQlPbvFmuZjmz6DSG5yHQ6LPZJQS
1Cj4elT5vPFVJviFYHSCo1Qn/qXgTIA/2C162RPHzzKpJfeqH4mAdKdIuMWioTmP
ursRgnfKau18IRnV4CBrUFY8D4xij7lK7vIUeltAQLWWk7h/YW2aAkUDViPHJZnV
wNjPnNFiokU2hVbR0Tc29MuTNELa2AzcUB/MsAy1Lmhi2ndwNXtkNX2m3qgk/nQB
OCsxYk8NHKacctZUC8xhNi1zu4DlJrBX7zoLXS5vzesLd9Idx5JRt5d6IkH4xQV/
KJsmHzGVARqdMyci3Q1MbsBCox3gwbqNptwhrn562SIe0k8bIxIhA5qEPd6N7bzH
gf02QarUagNke75w1Bl2aPzKe5KzxF82awT8xxjd088RIzYg1tvQ9tpz8dZSdUtv
qnci5BgQOs3VlML2n8WqwKQdJSm0TjfPBFRnupy52aobMsA82lIzzFFkeuip0GQK
awYJPodm8SxonW23WNPZOmd8EGZur/yUh9EpPaAVSJ5zbUzjIwnPQAwlttHOrUMr
yWCR9EfDoGvCV10t2bdJjnyF0WJ1pTAhkzpXffdldR3PXZQPKzXaFILlsmoZ/p5X
BvviGowYffOW0VWSFN1lZQV32na+JMXTaNsZGNFOaYSzzt0YKtXgK42W9wSfe9xB
oWhu7lnglMzq+qsCDdI3FD9sk90YodA3Mrkj/ruIXdSdKtR09HNF6UT+nPZsQohw
Va300w6Y+Lj/iPMat+s+3T/d06Vp3SlmVoioLHTBDINsHU56U2G4gEDTBgYNg4IQ
1hnjnCc3Nez2NaRPhs7q1WCHWEIv6aL3wQnAI2vub1Oyjd0nISUoq+dv1HsuLKq7
VYzk6dhz7JjfWoSZpsAM/htQWJ/yVHkl/oEcl55PyM2CELStPOLYY7HHFHQ9dFIE
1gyU/vzhsma88isGi5CVk/igPDE+9QzAXKyKX3vPulZKfV7jyQl8Kyx+WLvXyaKZ
uZ0bbTXpY2sULxsDkrDfy90ajNtFZNeQVeWjnd6lIDUqJ90wkRKi2tCEHFJRqV+V
gnKQRDSa3pGxtpmLe7MLKi8A3mVxkd9RqCDU9eFpXpZU6K/+B6Lq7/m1LSuiCV/C
ObZtv69xbe7nuTy6x7LjQ3IVBbFIYfWB9ndOih6xz/A1DO3afZxAjFTYRZ2RpMxs
fYEB+ZgeMcV5hu7U/IlRoKRxnE8RIw7gB5kSsMbjSs03p5MhP81HWxkjFz+76mLL
/KyVrt7fwh8MzENYk7yOEN/KpR+SLrXcQEN3KVLdCLeYIH0Ix9/U8HM5HHW7LORw
WNT73FVKUoP8WTZqxDbJCraY5rLKlggh+USzs/k+FuTK436Lb01bkV93Ef0RhFB4
YpjL0xmSqjfdW9fWYS2ZwDZO7T0TVXIuNwYLpB+9j77GR+c1dvErpemz84nhXcj9
lZFUVTU7VBIsRCEaK9b0xqfPifACEmJ5UvGHqpUsjkPy55qknCWPoDt0A5liwkLx
TS2BEmsggZ1khGXl9bApFeLk/6FLa+vxWCZOoqvnAXftU68ptSPcufM2WY/vPoyJ
4Eb0ARUKdJUJ2tQy23QD9KSDsZQwggsHYzQivgyjDYuPeVU5a3vCAlAOv2uB4ggg
p7+utBLv9nAIi9ld9N4PVdz3gZYHpBaf2gUKItNccZ8+6NM77eEqFQQYs1JlgyLn
/6XEu6LfxmNFmDDdfRGVuFP1aPObI6gceRyPXxbWBSy6azBjIOhnkzggxlQsaGoK
pJWYmbsQ1P0aPqMtXpvWYS7d/VPMDemitmIZaVbxxTzXcccAYL/otdGRDJo1xba7
kEBTsneBb8Dulvahu5diFOXJtilAXMzUwPJ0aLHjuju+n1H9Ko4Ij8SpfyhuAD18
SQHt6NYTGK+dpRH4Q3xumFtMfoZnIIdZmXAK1IeuCi79agvvacj03Jz/r7TvxZ2u
cQ1ItnnuAiYk9n4alDzmBY660HOFP6WfHSGLbGRWtG1i/mxQ9UEeJ86O0DVBSAKu
FTBwsVJvhB4PWEnizYcu097fctQlsbO3wDCthu7si+0nbqidMX/dTE1plw4j5hLq
T15gMQimr+VyjWB0H7Mh4VhlsuOWy7hxL0oqGuSEtI7ZBT/a4868uN62JqR5KCYf
6A7PfpBGZjwTiAFDCfKc18fluYoqyImIaJH0/c8dbttZXS+coFp6I19O64ZZwMe+
vDwGkuUNV5aD+vDUgqq3G84XLQpTDDoloSgmeMZYZutwwshKSbVh0DyE1FubnNfP
Kj0l1URFt3kvvWLMDq2F2dXu5+m8bRCllFe0fNRTxcGhGpfdCh6ahuCIl6sTP8l5
0nMX1e7zuwrtkLLxoeXEiof+/jShgHtGFcxdfAjz5/KFGtmRXQT8JUqCHlLnHelV
W0lFMhQea68PLGgXV4E5lh3kO703jB9nHkMBTo5CCzaYm8z278dKDPUZOVYT8CR7
pCUypI3738xs6EgC/DGgsHA+Cxl2GWYL1wcMUBqNZZ0gPB6jxOgbznkBgwZJa+WB
/Em3isMqXRoWeqWj7N5p+zreypNNYKHbF7+1ix7XGSdxvNSxZy27zGjoxr46sQ9V
`protect END_PROTECTED
