`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRB0oyW2+bO3PCVS9NcdFapiyZ/MRdK4jzn1eiH7GyDbVXi7wbJU+Ohoqt7HOY9s
KPcMrZHGGrGAxJsyiQEGephXn6rnE7GC8rAqRAE49UTPecAxFxmfxOwqa50/8LGs
uS/kF59o6/U+IU1vSeH4HSTRp3p2gw+16Bk2omaqySoTL+oB46oze1lu+CqNUpej
h5uq40f7mjxQ1LC3zljomcXQLK+n8hhYhUR9arumbA4d/ekuX5Z5oIr5rEEv3veb
l5F73i4C70jqYmpStBDtiBqFWp5E+og57TSGf663HShhKLPzCOnWxQfGIxGPGDyK
0b62bkerWbRg51wDZfDfEKHS+mG1h1zwnVF1mJvaCZnGzw177WNr8gjnOzKKe8Gt
aQF7XBhghNDCkerceEl0EHn4N2nHwifqHIyape+JbpY6zwqfJCCLXCXhEXkVKZkJ
B1M5601yByR6ZX7eKjb6Z4IM/u4dCNgz9oc7FI4HtQHnO8lRihTSgyxbifzPRA6O
Nd6cfZAF5hPD4YIANFXqggSxPwk2dDdFdJMQCmC3Ge9N5KbSI//oH6/Z8wXgMTli
xGb0GOgDhHQKSX0F2kzJfnknvWphQmvKwxIdZgovvcFLNwhT/chivWzTb2S5Op26
/jZgLjZaAu2ML3aMwrgOgEYO+uYH4EOTy7JoAs6jAqij5sasCi3en/keFNh5y1Cm
7PP2fK+DENkDlP8vLwRG6GbP53fqUQ5RI4lLEQ9VT6DgnwFeFMxhgmN+PQWRWpsk
PZZ85pDDpo8ztHzEqhgc4XcYo1ndQpk1PYqFPXMekzs22dMPE6XAtVUcMW+hq/Ad
qya5/T+V7ZNWTiZTNrWNAw==
`protect END_PROTECTED
