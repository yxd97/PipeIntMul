`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rFBqX3EZiOpgA0ZffjOcXYBZxroxy+WSgdPyzc1I1HGLb1EELzc8BzGbQJ23rDDO
HvQy5OZdm9t9OnIWjciQzM+H2UkTUlhYVjSsM/azuhIZifIm71Bz2xZYjyYWPC0z
zAydjV+2GC+tW06us69CA0BjpkOScVVQtiscU0ZrpeQMdP/WkDvtzsCaH/ZC5Vs8
S8dp4vcacXA6W+rfgzP1v15GCtEFpxk1YMeGXrSn3ch4vfSYdhKYEm5oSIT7igYc
qOXmignRFxT97iElSJEf5+ojnd9TMy1KCbTA/WIwBg/bKIH6KaMsdA8+No9FqTQt
lVc8xeOS4XdbSxqMQv/7zJMOVSEHf8PCA8q1bEvLiWmCFa9EfJelSW+mNgGydy6u
tPHaa7v08MFu1xo2X9ydbHfURnwir6DyK1dqZsM3F3IanQeHoVdIKw4VByNeHq1I
YgdK3DAXcd9f8U/ygThcH/aUhtnxvCnhmjhImZ851lfA1kgIYFX4uyPF9UWr7EWY
WZYoiqt1/GaYQr7Uz+o/4gUfaU5o8W6ddS2wBPgLKl9gT7m16nkLCkEnC3ouckus
O+jX+jFtdp8sDGutU4qdP3JNii+2aFbVII0Kb+5ZUpo=
`protect END_PROTECTED
