`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qe7hkLe0loiCsRG0Zfzlj0INAGWTLjwGDjyI8/zM9A8I6yzMqvYxhPGgmZPVwy5G
dYGGVM6DL7uczd0fXTERkv3Cn2uXDeSgF410p4sG3aeiCYJ7rthLSM95+KOYSIlY
rMyDrlmvIk98ESEoiCwRGVJsvBYrAr0fINfwS2zpstIV+0EYLW/lmPIg+ib17GLw
J0wDPLP5t7LWB6XTHvrUhunSQcM6MUHCtdWJhOxLKjV7pX5fzdT9ms3QxYO2r1gu
S+RmsfyURQVv/qJoslH+gY7N29tyN0EtWwpSHymVyw86DyOiTptF+nRSMXkwO027
F9IhOL4dWtWvlpcCRDajLl6/VPEW/Kaxx8t7G57eg1ZaENLA1F7TdFsYxHdF5VWJ
0R/bd/3opxRyLjwJnMi7ywwqDysYZZt10pMYgWWeTJhK9ALbiG+2vEQ9LydWaEhk
29VzntQo2UmBgShGncziUl7QOgeShY9kmwOaVN2gVo8wRyEPPAOEZiWPM5sO8pE0
mWszRpoY/sXpdh8bF6yfFcRiSZ9beFCpUjFSte4dV0+KUWy8aIodCLvCjw0/IfN/
KPeyB6eciIE5WbpiP7Hj7JYA5ca7eonyuzWOfioC1herqfZuQ4KLlC2p7wfr8Ice
Z6SskZx4hptNwzDIL97fJt3eLWArtvvUwkK5RzFIR2wmCZznho4NWiH4dw/35HO4
ha7g950+3ipVZA6qb+FDTUYvXcgkZ8R1DgTB6LIt17bRs9YmCyEyyOZsTao5srUJ
+lAPPeQeaEHokBSmbH+EuNUJa6M5vwmZ5G9aYOQqBPUgK6QplFUP3xxytj2sNFAn
vdQ6al9X4dZsR5yFTNNFYkWTs3YBHeLR4tyGf4piYlpr4eYFI2qqf9p51425e40C
QIymlPQg5JH59U3b4tHFcye9UPVLyz8F5rBX0zqY0jjGb7UGLwqSZs9ZUuzr4fbD
JtZW8WVgo918meOoSvyMAsiZoCuNKqLM1fwVEr7CiaVaGa65UEiVFk2X24Hrlpq/
r8zkVlwNpczuA2ZalcUWb7P1j0LLjABhySSVDame9cXDAsZGpq+eSYUqNfN89z8l
HVVdlslnp5IWmE8yJyjCgTHOCMLoRWX3yxdr1mRGe3Dj24VqqvhIzjBqD/gOOlrw
XqlHD8m4e0oTaE1rD+dVTcdaV7cLd7moJ4Ak2Ab7b9e5ptsaCn6WLBqBwMMRFWXb
f6EZPKx6eMw9zjIHCqFH/9wCLVc+TmTGtDj4uXNx9MqJ+3ML+NQ/2gGU7qFfBFeE
F8Ktwu7YcygdPjWRRuYfoyId0tBBA8JQlXvhey37vnUAVtBd2Rda4dHlqWbs150e
qCR5sB20k02uayxtdxSfeqG8IPGGkvLdHun1uatkC/pBmNfs3oETIuek1PTdnJvo
uWi8NZu+0Op7+Ve3zNmmBqYxinoAn7vw99/hjusSgioSsMcR2twuD8NCCa56T9DL
QyrfsMadH3ZPyi9DC+Zm4s2euPvwHpnEWFV5XfPtugrgFGBWM5tL3tNvUbbiPmpF
o30fgXDwwkt5CS4QAOeWTAFVSOQEsb7Io+rLINtIGnvLicFUMf6CKOlxhC2F1qFz
7AbEeDlarOZC1PNGRQOFAPQ1qyWoTafAej6Ky5qTHy4ChV9i7iO6XlDNAMUJSCgr
8wHV1C18YERDhTBmMPb8ej8dbXOcG5skzPxD+8uS5B6jV3PuMM7kXKitYFiND6fR
u/CXFEfxZsoyRc+UknKMf+SyWAuHzdo8GzjBMMIa/u+Smri4C5UdeXa7qwvaY0FA
PO0+T/KD/vF70r6njgWHsLWtGAAiNUlZjcuX8SKiIlYioBKBODkJwg05OcopCe10
y59Qceg1+S9lUWMjWXZgoARJcpr1fQbNc2dRixzZlv8ht0VP3gfR7LdOzPFLeKBs
u94izQq50EW/lA/lL03TH+6WYq1wysOv9//D1HeNUfnA7pd6s8mV4zbSttdzWxdj
Oquyk9OtGLFCwl5Ttc64mHoQYhK4xbLSykoEhZ0VajmZLV9ca2e5HyJuT/KQiGko
3tTR9oXn3H8t96ma1GXH8zsKuQ8AB7cYvUPZdepqrvc=
`protect END_PROTECTED
