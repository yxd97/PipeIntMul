`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aj26FiO+hy86e8loyFqCLBIXuiChgop9AEkQVogSKSGcrGPOE0OWJWSZz/IGyLc3
t+GrNmlGgqLDsAPPjoulIBi7xuIF/EHcbEQ0/djCtVtdhdSvq+Nce8HQDWwAzjfk
BiyqA06dftoRPwUzr9QlDgn6pLr9hlVNUP9p+KeZUoFDQtkKq0pqCtqbyYQu71pe
TvR7oeowg5b1OvzBsSNmxZo5R2SB/LnpA2A/caDz0+f7H8MSr1q09ZG0VW321nqo
UoKu8wHVkhhebFlC+L0QQJ6clNZGoPERQ9gUffJNomlc/nqHTdoDn5oTCffqRmTl
zbi6VZDLCiYeFBZPdiaiEg==
`protect END_PROTECTED
