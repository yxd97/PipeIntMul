`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vNYkKiRNgaNJDoHQBF0b2xpisAI0b/e7Be366xdy8LsIOUREDtsmv/gCurMrY6pU
msYgC+yzMjYzxzXc6SBz5l9QBGLmkH7Ye9Z93molEoFBQVIK9gFr8gzDjO1M/4PB
Oj4pe+LoFuSdXCB6myn5fpKbsEZFZebPe9e5UbKkF+47IyCikeuGkJePWnRZw9ZE
4qGrErfm2Cia+5N0dfSrnDg0SGELj56oH0wpaVrn35xXk8iBIT0I5rTFsIsr1XIk
BusuVD7izjGXCwAKrViEHHb7I0m0Zr/irbs6RzQVFSmqAJnuwblw5xg70oUWs4UE
X8oxi2SgJ647Kfnn+e+9RAU/NGJdc2xrbVwXo3vl1tReOb7iLA9u/G9k5zFmoO9L
tbOaxU/LkHuPKBZNxvc8L0BCUIv/h9Gb6GRC13DRi+++s3GgLEM/tpU5+Tnr6rh1
DxsSoRoUAe56hksme9vlpDbVsGm1WujotJuL5A7991Yn943GnqRkd0dqTxQYfVso
JdH5HEmZbzegppbkA5LXTTTwaeAVJ+22DEQmv9Os36JpyP+hReFuspT1v9n+Dh9h
VlmpvbtfrfVVGEWTdmW6bctla4ev9qs0otvm/oH0sbr95aZRPqvW3knZVp3T02FJ
kQZUvIwygW2qaoYPGXwArsuiY5/jzwgQ5TD5bcyT6b5d5eZWD41NE/UET7/BqhnN
7Gms8Y59wVac6WJ7HPXA6X2eRTF/6PISaCjvnxR3gS4QCF4GguvZTjXNqjGoSjuK
OQnyDIcZNXkyI8EfEmbzfIKxh69Td3V6haRqlNiRicKLBS1Xw4KDqw9Xqbhk3hBM
GBXH2sNBenJ/cBH0jQCurA==
`protect END_PROTECTED
