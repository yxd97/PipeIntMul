`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9vltT5qT0xM0u76wInzvuUiPmw75ZB8w6nWSjAyN/HbIjcSGKnsWV94nVgG/iar
8D6vD/AG/MQQYcNxEf7MvCbjja5nLhPXtrMf3CstnoOSL5eZbpZQOlXwUULne4/A
mgTccex83qbufSPY1XmNMoaqRFxo5PFCrzE1PsIJrMYrao+ePhyfm9ZaFrDL3vsW
unWuauDb0vw5Ge/XQLsuALBKcuLjuK1ST3TgKSdyPX1QAr6Nmun2JWaLvutbsO+E
SQjd0vP+Y/UYQJXRP4Ljmlr3CkFsdi1FOdAJdgCqBmFw+i9I8nD8WbAy3c3MOR4M
pMcIpMH3pd55VpBhzd6loZYZ3lY9tg+zeVTaKWUxRlU9MLtfNRSn89Feh/LWDZRq
`protect END_PROTECTED
