`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oe6/BduGjA0Kp7XY8QTbxekJ/dQHQB/zFp25FG7Pp6w/bFqoOeN8kxlZkrld79Z+
q3PAahFy7/oXC7U/CC/2wzFUKNSBoW75OMDfiabN1MLKWPTief0oTUXXH2glHo1p
yQMuUzADITZt9k2kAXYvt/xTHsLYQRZMq3+/Tt9YJYpgwGmQnJTIrCOUjDTSP4Pp
GVxqPDSPGRpPkKoDiArYoKLQuDoXow+6hj4ZZF3x/nGEMp4F+/o2aFw3kR9zp0Cm
S8WtKHGjj6L8Nh9vHssokdgqdjdFZKefCfMSwoQoLU3W4eh/vqhYXsaLRCAwLUv0
9oglffFhjfixCc0s0PVqgQ==
`protect END_PROTECTED
