`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TwQXWjb+ly+KU699pqvCUSulSh1otwiQGVsHptS62o/KTVJVs6xUIUpxsmdJCUez
sMvRuJp+roZqceHmXQd4VsQxcmEMlVm5BHPVVrmiQMJZt+4wtx+Bl2v9Di+Ftz1y
y/QSd7HLBtV5DyrMauNZ2MJIrFpmIMmHspi7hAEoW6y6vxeFS3EoJQu0JayMQAkX
0PyUSO5k2lmJIIh0JGCmuLhIuQKx6m26ZGp5YhssdoVtyiTDy0xMhIfMY0OuyHoC
2GVYQ8bnm7gMAT+MLAnzB+mtynb4JCBl1338uGGgxfrZzYoAgaGF4Wks2Rw2CzQG
ek4PpVMoxJDgL1Np45BR/+r4Ln2MMCpt4id/mEBzNAw=
`protect END_PROTECTED
