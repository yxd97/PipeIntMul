`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
beuqMe0sEyjEwqOKt9HhlvBh0cD4WbXocCh8QGqiTohbTlaRiPiKy0KrwkwZPtLX
xrdqN12C8HnpTehObPFzGMZdy8nks6YqNbfRE6teeg4zjhbbh7J9YFawXs04eJYZ
47C0TRg2RdMIM4yRzrAQhFoE0d0zGqkvoVuNEFG7xLot+/in5HB2iNh519wr4a6h
sEgvK4L+qJggZubbOLu4mtViJfC38DvUnLEFKcWobDbU/dbh83DvM7fkBZpQDRYA
/7gd8rvdM40SKKGgxSMN/7EJzycV4IVGFtowFGpm4XZRI1N1svQ3EzWfjVKEcuZJ
0TfashAciFIJ+QM7ebsaYWUIuIqtSabVzTHXWUv94AQjnhsp9/yP8oBzq73+l11P
Lhl3EpUWqIgrsanteXNE1g+E6U/hdP6/NlhmdbjSTkVBVZdo9b06ojbsBgrfOj4p
4dJGHVgzDarvleUyP3vjfr2aL2mrSOeiLFHCC0LZunI=
`protect END_PROTECTED
