`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
//hUUOTq96Pbf+VHobsg5eskXYkrVyIqNVQ9PTNMXXcLXp9XaiIZLLwmBUjPbUL6
EFZfYvlQOP5jj0ArbDndEEZXf+2UeP9bNI3v9xAs/l1l6vaE7FJMB3/BDn8GjB1c
8r8V0rnqFwwhDH6V6zCeabv68fI+13gGMfcr+iskuKMsc8CLkJj/KkNE+ikIrXf/
6qFiYhlqRfGdgflRH92bLrCBOib/l5ohK350Qr9Bh2kyQ7iRY+7cYrWgXUPdk1Py
FyePfD5Ksh9If6A1tDTfBW70ez5aa/n9RKXNOF0gv5O0OwK5ZP9PU+WTDaFbZ3Ef
EZsGs52ijO7Q7c5oj9MprC5AK8TQjhaKh984SZvouwo=
`protect END_PROTECTED
