`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3qsiQM+iJnzvs3FXnXvB94EDtmHWsZgsnFXaRCLUUXBaILMDnLw0RxPmfXhrrq+6
wpCrqvIfZgNqbpEq4cdkntacf12Gd0iroYpJPBlAqb1BZmdY5Ygx0MFh8GUx40Ss
x6MjcjaoMNshhE0ftdUivy0eFUuJSXyDyUHoHbBsuRk89qfMNEXDGfUcckHyuLW1
6ICuKfXihDx8ruEdJVGjsOvPTibGWSdIpevR1+7LzLKUJvd1XbDPErVK3iW0pL4H
6PHgRSU0H3BjkymIzB4fiyeixt2LVT+aAiBRBIPbR4Bpy+cQXppmb/3v2MiTeRmj
B4LhQKxC7Ai+kHFna2Hy4A==
`protect END_PROTECTED
