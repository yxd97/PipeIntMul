`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7CE3PfS5B1+RsR6hNkfK3ajI6DljJ4hj4L1Og1dOFtpy/uqSzjsdrHwK6Db/1/1
lthZKqRQIDzozi0GeJeBm3eeAwk7qpRu4LflzrIEHJY0Gfc4hEKZnGXQNawIFrqX
F964SwxhxuXPH1RFFl8dIr5RfYgXV3e7w6+TdSoPMA2NCvY4MIBWx4Z6s3rK3hO/
Y5jah94nM8A+zmkNFvMUvn1Q40iVn1lJXvayX3J4fsbkpANhkc70M6mhVKuq/AYS
Sv/QiwG4wdiC93O//zJRuz6i1mYdKZc4nMsHGozbb+2uVFAh+LRqJuw8J8OoUmfk
ciKsdvMB7s9+mdSudwca3JVQL5pgbLh4pJm90/dCIiwUegkumiqmfUUNQM7mvsvD
LxAzynAsmif+WGakDP0RYJGQcEY+eOof6Z3lC8DqyzTPJOgB46S+5VgC0/xBMty1
cj/q/f+0bMyo8JWeFdY1ZIYiJ9Hrzb+W+OP1RaxIb2I=
`protect END_PROTECTED
