`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0utIh9CVuGSH0Jxwh8osVrvQLfJ1WQA1WhDXjusyJGddEUT9RMrdBUd8+bSXHPDI
DI+oF+NqpeBg3u8PuRV8CKwQ/Ra2CS+tGkgDZ9YkG4SnkJnrl8geuB/kkNrHb9nX
hkfPoII+uyr2y6a2CMzNOH41OVr6/V1pn9Nejks838BErbxbM45qSDoEKjVguXfd
UGNDesUf31mDyI7zLNUBZq+TYTow+/0dC8TJgvhsIJkeDsojcxuFZqLmR+10qvrR
1Im0T88MbyQ2284DFhRBkExfNw4dOlF12W57yVerfWvZ5BUiTbFAc3Vaeg6cB7Hs
OwgrmgUM1GnoyDhQVgkXlygJbXEdzJKzj0mu8rnw/Rr3ARf6dELQwhqtZMMaUmLm
x94ilwD3Enl9oSYFBfr/O+OG4epB/SsXIrmLEIt4m0UvtmOq0rTOnH51UdeNQngx
4Dw4BKPkpaiKZ2sZMTrlMR6mLIAYQY7pDi9sUOGHlpQKnr/RFrafrUdmPJG1J0P/
HqA484yqL1sU0LzU8zlzt3FJ6st6VWwZuHgmbsHz0m/H3vh8Au9ipSQFkLvkoDyS
Pp2RmOnPzuZ1gQLEJnBGbN6Le5dJ2hKL1d9Y52C7zEo=
`protect END_PROTECTED
