`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fCqSbWl1t4lotQwmMKh5YqhOzio5n819+0+Xq/IH6EcQBXOiXRLiOXwa2TY733bd
KdNik4FjqaCUktSpJqs9yWFN2nLHYnxonDVGGWrbpMWxfRZJIDKr0hriHf1/AzB6
Z65PDAk1CUbzklMVzhSigJBcUc7sStiEs1lrijHXOPX7/VEYK/Rs1TfDx0h6GOEa
zGufKw4VnvljLT7x1XRDLFi+S/8gkZSfVxhIlvdYWEX4eFgRP9CDqHtowxe93IJS
6qj/RmGHP6AXcUX3GTY1qR+iBkPsvwhDh5gc6iA2Ass026niEQtvA4dT/JrEUg4D
YwB7cmZtT59XblFtJp/Y4pugL/81ht/LEU3WwMUfURhdOgLpsUSQVbcUwjGDBteJ
`protect END_PROTECTED
