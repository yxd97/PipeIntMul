`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T73QLQgpG4BsDAGEz7g7zBjKI9hfSBp3e7QO0ufMbsWOMjjpOrTAB93R+Q6uEsMl
TJokqSLqxx1I3g5Zp2nJ/yKLrJ/MRzTttyN745xSuD7OSCMXYfKiz7jvJn9PnTCi
lr3haBw19wiYHy1v52faoikbwXvRTlmkQ4Z59cv1QgKq8KMDvvudvibRzXPlq5YS
I816n9WlfJMkkQQkneYzzqa6PstgMJq9w/JYbMAB3OfVNiimtUYm/QM05ma+ORtB
n3nHvcgK4/Y/hKgjOXD/a1ghc4H02agkEiFIBiKvA+0inSKkZP08auoZoLvnuhZb
BK2YAszh6yWNtUwYz/RcgVeDTTD4F1X+NHi02lhN/PrNjsbE4aBE3eMi3HvxEcW/
BwKwZQm/0s41CSKcQaxbUPI7qh8QBXveyRQw+SDO/onSTPquw37BW94ivKOOclBe
pTokosPXOUbNDsEA/Z17WI1fNFj3QsPAQoRaTTUq3IiJomABs1g+7XJXbtI+RwKh
ynsxLAgfZ0y6KsZ9DJkmxv0lRTwDl2e4Y08OLEX7x4EnqYWW40Vpdg+83+506f9B
TquqD6cqyiNa8yEPcZq15Fj+Ug+MZ8eK2BsXEoXHCLGKH0jTSqeKgbnwXcqmvw0k
`protect END_PROTECTED
