`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqiVGPNWlOP3hlVmXYWZ2VlC4iGT/NHOjgv3JMoZj2QuB+leK8oMdqekT6TUdl3j
+IodicLf5/a2P5GtmrYdlwYYritP+YipEfGbVeOewWc3bwjOFSX1ifmPEl98I/5V
al3ZSbrTbVmjv00hoxj1S50Uxk+BY+RP4N3SmXa2oad3R4gx8Yzm2xXZwFMXPnoY
ypsBDMBZzoHJwzKwA7YyV+THy8nwq7I4C4wMjl3bFOQHiqVa06kC+Sf5YLL+7LZ6
SD1QEsvie/ghFNycrnvA0BDfYl824cZRkpzLcKUcFXC+rHFUIU0wwatHmROVnM4M
AGAlbAqZC1daiUpixc63WADB4BQY37MCM8hDP1BBQAyAFMQL9XvLx7e0M6WcIvX2
U27qRiWvuDAVCRAww3RBSyXllo8M4fnYOGg60BziEsG1tI5pKGbmmc/s/rNQaEqv
`protect END_PROTECTED
