`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8a1noCbPAeV30GeovXhTKzD9NIXYXebqqNMYmPGCquyPx0o0xci6Lef+YiuSlibw
8mme9JY/Znb4CzWLTzeQ9DsQMmnP1rutRZCqBSJ4xBkywFq3HCkuLRRE/tWf5e/j
2ear4ORiDp7e/SFJIBkIxp1UGWtqHuHH/KfkoFqc5rGBM1GMFM+rJb+KUOW89DXP
bW/wLvBNst2VwbDU7xxP/oT5vnSswlEumHAQQScB3R3BD4mgf835o2xSOz6ueoqC
FcNrjjbra+DoG42AMmiUY2NIYwhM8yIwptOoayZ2i3666YJwFnMXLcVfW0/Ht+/c
1i1QpD6GIDoQToWZmCuSPdNk2Q/0lrFZaV1uJgYD3Krj77CY2nxO4Fn4VtESnvg7
7597oPIhcpPFRs9jPlOnJKQg0kXHPZfEItW3ij4OLASEs+oBVnuxVz5fBhun9ztl
`protect END_PROTECTED
