`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
srmnF4AFZ41XnUCTXnUX8TYIDmsduG6sVyjRuEV/bNCqsf7NbRzPRbw8MKZ+NYX1
eHp5Sm2k3iqe1AgA6cbe/IA7InJdmVoIcNiYAMFIwxenAOStC5O6P8HOqfbEwE7K
0gOwiDkX56xWcjhWKYKQAKtBOuwA+HRNyIMz+hT3BaqmB85i4a/avuMDUXIUj7hd
yUsCHKXNfWeHf2JnAYBjhoYn9O/r/MD5vrO6wISA0lmCA0qNuTfGrVzkZoQWK3T/
hqXABgElb6wKXFqvJCBP4nAKHjV27UnLqNpuUXTCThCdEszTOSN/ws6GDGaquLyq
lD3LGmWGYdH2PTXgafpoghFRLM3sGnyaJOs2RMV9Rs41TQkunvg2fWllNjCDsghJ
qA3JwODA2/Sfv/taQZAch0fYSuKCIuyiX+HHdh+9qtLEchk+ODw5Ovjg5CESQXKW
WEuGZBbNvFvgjVDoy9FtkOa3J32O3KJeYVxaCNkLkasX4QIknrojuUxsUoS0R7Jv
YpXalF4mukShtUK82gVM3fFWLLPpPR4aPflVxNjuWAHx/SrwrnCq7NgrchcLZ7rs
cqpCvuPkLxTeyvVLRP2vVBgFlH4vQZ/2/m4f0E0bC8R+L5Ejzh16azyNw8mkbJr8
62zKo3Ah6SO49dqrVT5qTA==
`protect END_PROTECTED
