`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkBafVoeTkLMEOQbI7WsoCkpbu+AQUulPJ4x0rVPElLKKGQXclH2YZ2p/Kfw/DGR
KwSxFzLUwoRD9L/SQkBnkzfDpvOwFDIGuF+oeTrYcDDy5sm7EXEY7WatkmRpIKid
oaAQvU1i1nhqHYx6CTj7cGh0/81JiSCnizV+hqylUyt5+UBnH9ECXGLXO91yKNZf
0wps3+LqBvWTslNfBgn6MTJ/uhdsHld31WFa4c9rhXB+Elzt5ed0QwW7xroS32NL
18j/IBDGfIJBVcIhZxpYHvK4XRGRpkV98F73MS81o/JjD+VMsldfrlP1aKUajbKr
2NkmL9I8OrFFcjM98QXwfZAPRhNAWDbunIKCW4122j2cPsoKtUSo+Mc4OkFUyzf1
zW41+9ySV0n/APpSeugGTuOGBtfhWd2zHI7fkgo5G//Yi0mRahcmbTQi0/HxjFK5
utwhCUG96dunXDU53nVzKzAYd2Coir2G4Mc4RjsqNEZWDRErtICdNZbfmD49u5BE
ZlqCuDlmk/Nglb2vbgMZDDPbGeHpg/evvojA381xbN9Syv+WjA9DHLbubaFwvgNh
cffpGzsfwDGAg2PhQ8Ysirvr9H1ZCoSxV83WpWlnlcYqUhQMZGPf0vDIgYJIuIiI
zW70z5/KZEgsjqomrNJQnmygOGFkMsCYtFpxFfDT8FM=
`protect END_PROTECTED
