`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFFiZNVw7AV0ZcVcrAaFBxmaA4mc9rF04w1fqWusoOmoJYxlqQ6NL5Lj8z7AqSmT
B1ivyApjEt+GokFNObrXjGth9HnmWy7PXRx5NhVe9CZIr4R4MuYg7Gyl2jAZX4Br
C43W2gzQ2nxRyZZVCBhf5nrl4gQG0Rzy1wlUSPIVzp6PRmeAbe7wFiUrnV5AG4PQ
h8eVhl3zeq0Jm1dDgrMseuOyi6MY6YHmc9Ff6Vj3gF1ejgA3koUdU0BR2fhlPXlW
n2LcmaHP+SV/anpUOO568BUg6Y8mAANbpGwgD6IyYHzokjSaQ2KzwHSilAprTftA
mCGCeLSQgapsNGPhTm0oW23SirbgMPbGmROtliKtWzUZjd8rH9v4v3LaVvIxqq4v
Ht3f16ZIX3cTX9EV5xfnqiVoGcnQxqERhhn88JTAgQZoADvDtP+MqTG0vA460Seg
5uHtH8dMUw/CJtod29dPRvgT4+GS8bCEeTS9oZbym2y0iWLztE4YbZ+mFo5xqyfa
LfukxHPKtHiRmF7R/ZMSBzAh2phoWxjoyaG6F/2J3njjhn/0x+P4FF0vjuK0EyPY
rNE8e5NnLMWenF9CQRrpufbCbOJcjrbSX7SyEsAlwfHIkBT//LtazccUR8Y/cnBL
H32tcZl9I6pmNfl+UtmRzWVGTcazQ39bu5wBhV0CGfsB7+ynXEvTm/Nl08YLl2xS
XZ7HAR+DQ22z2R/z/rZ6SBIpuPi2L75icYJe474LLBT9RNiOXsolMGabNPmrdf3v
2HjWWlyrPJavT7Pbq06j/LjQH5oC0gpopLo37N5dvyjDCSq+KKyUpugb3MGs2KHg
i0yQkT6FU6qlcF/YnIUQm2DNn4qzrgL+UXkN3UtcPBsnHLdl7MVD6g4yjiGcFlUK
wNIEx2tUNMlIl/efYxhYklH4B+KmDjJWEyXWa/hfQAYEn5v0CatrOH2k71jyLem0
hgUh/TkiEAFlWvrOvb/Fkg67qMfiS8mcvUwugCsXrnpCgqDfD8d3RGc0VofGQitN
Sj+YM/ZnohG7QQRzFYsX6pCBhooEbA1WahFPdESq2LQEbczlanVoPF5zXLu76pEu
sosjprfTQlesie/bTDH1CZD/JZHrFO26VuvHoItNuwD1G1W5/I4DvYhN15r/pLw1
f4WvV2C1LxwzhZIEVFxg1NzWXEPQI36LX4kQi3nIWJg1+xNECcqgTqyFq6Xb9qUp
WgX7EB5AAMgvQ625PDpuYFnOMe7noRxAYkfIiabV9zozdPSt2lhpfD4bajj7PJq4
4FniNzWUFAIqF82Ft4+XRLx7MIxMQhRmNhPKvTwP6I2I+ufeLNtsTFNSbn8JyJf+
VvGfIHfsZbslvi9gX31O9Cnn222RYjfIsUDXZgRnZo0oaG9qiT/7Rbjfc0aL19Cr
b9s8TpwBWFUyQQv1E5LH2JCqGZwLU7FzHkA1/tq+0E/oorzeie602vRVR3m1fTZu
01NlOTI1vGBJmch+ybPPXWEkpqzwaoXVimLkVBtRgk0Kv1dkhhrRpDNLd59pNLTQ
DLjJsoXa6/PbmJ7RgPSBqavqLHbiAU1RjKZRzjimIK+8jsuRCan++pEgEiOHzZHe
0Bg75BKYwCMNgbXreluW4g==
`protect END_PROTECTED
