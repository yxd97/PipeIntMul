`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uAGw6GzSvY+MaX1ggVti6QUlPpXRpfwY4EXcg38rFhz+X10MWcbVRAaz5aFi6DmT
2QzQaESGhregWGmaA/0jahu6iIYhOS4/IpHbISU+nolQioaBdjPAaD1HmsX3wxRi
MzzxsJ9ogwPZ8X5izEL7EhW+Qku+GSTNj/iLmBy+rDB3KaeLnkXN8QklO9vZJjmA
/s+0uLnp//wqsYtmygc7EAsqeVHPx9MbqhN0xsXQ5EYkMNcB4XryO2hyG2fd+ClX
42GNOATtrIzEj6P6TkOBubDF6ct7jN6CXH7Ls4Lxi+Tv4t6D2cTYdKVR9nJDkhCh
9oXbt9CPxwswInC7wBnT1ANog70EF8AYEhKruVOLvGzMee/47823p7c6KfzYXSJM
vecx8KjO48sX6HeHZLSbFgg8q1cc0N1LG7HVbEYP6fiJ+dpnweqjg9NYkPkzEa8v
t3yU/pQak1arWQEyre0swgVaPemsdEeEktJtR1Rp7VZPXTZj1qiOT9FpRxhoPHpe
Feblqi1Y9uqOk0UFL7+wBhUDZ/20ANRBchHBD0nX4hP0zxnuyO4idhLb2EN8BVa2
FpAXrCvV8FbUxeVOgdvBPrC+UN49TrFVS88EMnnEPseeehCRCO7pEraKuGBjCq5h
CF/PWvfYU/CgZsByUEiWgVb5RRCLgS5nIEX6WTPo4xhH23GLutD0Xrl636xJm8eM
2A8L4UvTCmtKcO0eql5Cqg1Ebqx4IuTkhCOOahtOQTz4WhENeRC7jn1MT3tbe9uX
TZovLg37kewu4C7u3W2ezG9XTpaSCQHfPVAjME2MVHyD1qXPebGnQzyX13hht4Cd
Wvx8Xbmw7bUcaeJZvKR/twqa60pjLgDf2W+SnTgd1G3pweruhGD+XhY0gppeo4Yj
gRa3FaDKyLPGSre0ufSzjQwyMxohA6IZJMM5Z0Mdu+J3iBBr6vqf8zUPgHhTCyAU
mFyANrT69jS7JeheEClETCuiprfrTJJvgvRQYYVGroydFod/DyQTJHcBCoqB8jhG
Zb1l/iq2Hj3fyR/szm1O7OuOIbXgoruiHXfw8Gv4XxzXtpE7obeF6i2HJXLM4i+w
6ZbPQ+9jfNOgTrYjfZaJrtSpBnuSA0jbfxskFOeLw8yxC97+zbhr7X1LxHw7X/LW
uU+l605dQGid7J4Jc3khUAbjEXm4WVLsDzFBbR6NIlA0CZmkVsecxJiwO7iOQ9V9
oePmoLupNpcqCDByvvP17y+pc2LD1uR/uK4b1JHBcENK+rexM3dwONKqpcbtojNd
Wf+fKWpylj/MYEluch63g8M5wWWM3KYwunlCrfn9mHPNZjwABEtCA19cyeRnDQ62
ZJj/pwAmb5E120Aoz+nT7jdRZ0BKULtZZHLtwwBjNlhTa6LFExBjrUeSi0Kc+5IC
mvJAMp/0dsLYWRhZjwc4Apt9NkqSLNNUof1uPbxqsyfnW6nEXz4cPWHiPm9cFjV0
V5g42ri8rCDcwDj+wtlqeSCX1vsz/LxaoDvC4+FH0B6iHNiJ0WqrLSZ2pEc6VoSZ
cE+x8R3qGXeVOqWQbR7xFubqR0RJReOQlD6ADAAXqnPa+JW0JCzfyGOnQ/O06Y3o
9uCBsutEAiRrxD1SYjZAE3rbPf5NN244wK59RzbeMDRjuh++Np3bsWYzda9kvAJ3
Q6EqO5EL8NQTo14DgMtDT0UH+XBlJc55LaXJQds2rzW/7j2PSUysq0GVTvEZlN+k
FEfk1qhG8esM4KqnNgeZGbg86hT5lIjja9dtIx+ndtewcOM8zakoid/yvupovdJB
lSKiv80xyk5PaUc0akS2c7AMBYaNtyS34rBA7wzA9twA71POImrv8WhaRmHhGMf+
5nAsObUaOuH1t3tZF3WX3zKuksi/EJX7sfv42Y6+NAph1zagCAma1FTq7qAjx1oT
Eitnc+pBJ6cK9dOUeSmJcA==
`protect END_PROTECTED
