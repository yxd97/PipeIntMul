`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyAhTKxJykEayKz13jiZrPGXBzqImr1uxhNg2qCvExgqw3GTJgWUjE8Hp+EDOITt
CHL5JaQxZ+NqNH7pDih+j+nfgVLz4SgkT8LSXN9XiyGnOI19G29115MwAre4GT5w
KS4Bucgfl5fpXNV+S9ETPGzmRscjef2vRCjEQzbmBfr7rD3/oWVpASgjA5BXm6X6
VRmSs47K8o0rrnwqF/5rAyMUluRKtlcLF0Hsl4cUryWvXlZkTbBsyQFkQ4DHOZNY
PcauhSyEhJHHjf0nNaX323GUUXIDGHQJHjP4v59rY0o8z2CObWGuLQASKWHssVb0
Ry1zbk2iEgI524xbFFR8f+8H6TKXrrhK7v5BUOuhCDeBkbYcFd0eo6IWjUVndQKc
zgX1DhELBoaT/78yLdcInnnAE7xSaJ/wLv5qX3ZdmXzopL8iKFa9ak7vVDwXw1Fi
Td+pQkHVbnn/jaE2+LLHCg==
`protect END_PROTECTED
