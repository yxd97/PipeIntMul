`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VIej8p+OGXz2RO0IiM1OhRUHueT+DzxbUU8F2QFOmQU5mU8CpifhWRkd9DNVARnh
nbBLOfQuGQ5zD6v9xKk1f0OQz2zEaw0phniLeYAPorLErAiBGkfM6kEh7tfHTk3e
ehoWMxTLAX9zc/VNxRUtnBhOXBrQSr6aHcZZQPptv5a0swxlylqUoeJ5Ycl3792t
hYAPBB1U8MzdIXqVJ95tczY/tBEba+uNQ8sDJyfc0di2itOmGpXlzFM4e8UcFCN+
BgjH/7Sepm9ApZ+wTsTNQF8GgdcdjobaqrAuOMiIRvRjfwrIs6UShlLeSUFk0prS
ZBrVqxIMlQGXEZk31c1osLirnrev1ufau7xgyhJm7KriYjJZKuuXmS2anNHFzSEi
uvxhkTmqomtPIslE1sWJJTlefFyc+b4Nkp2F0aaCO3sQiHQqx1WJ5gpCmA4nutWH
vM+tyy/14i8yH/92AtV+1c3DnGCLCd2TVcEg3rSjUmdbI8SG9JXVU+LjcuLkB9sE
JTY+7Qmf4/6pjm5Z5nxIale+atrAIHCJVH7HLI315vCgMUB5kL5cArbN0cZ5Tvga
T9AiEUdoUzYUzy/B6Q00xerCjffaXg0dBHJW4H27FMcYmNWmBVQSnLGjILKXUMBK
`protect END_PROTECTED
