`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L0IWJSZ0o4wD0VSml6oz80wYIrUIOXO1XEjD49MJqIGQzp9EvbxljcGidBOgF3mn
QTookop+RXk7u5JT/v4aqD1JJePE4sch0nkXdpb56XmX+/TEfFO8Vqtvp6sJYhJN
Xqmy74GNGGuLJL0jjITjNJgfkpAiwy4fpL2+2Df8xfqDodlBCkuLksgqgMoy3ki/
efMz/NoDICvff4BqlST7Jz3zlm/j9uCErop7ydM54dogBo9QD6WMxjg4MafcvByD
im37Od/qEqRkZDbFjUBEbSXkSI4h13Kid7c4ZBx3cjxGtLbd9JJe6ofX4Q5iK9aN
WTqDqFmY0A9L9xsbGxfd9pGo5hbp0QvaVHLgOaxBSRM2+uIZuxtSoGqx8Gw+rqHq
McFPCK+hI+PW+nhhihTOig==
`protect END_PROTECTED
