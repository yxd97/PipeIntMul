`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bkEbjYVHb5Zftl+/ZRBit3SimuQUyAueAzA6HxKrrr1+OfH7hicztansid0HHbF
5iAYRA+AyRmvrRUw012OA4ubI6jh3v7pU0V0QZX/pX9dpy11yi6OW9jySrxDLa0p
TRrjFvUnw6UDitOKyIMVs/oqsi34WWY4Ip506o3qQ4jVi6Yhnxo4iIF/qZbhR2kZ
upfaoPCwO5qt0sQ2KLC3G2ZG/FZq1rO5gTQ55ZSnXUV/tYS62KFTRFXX+GfFycpl
TqGvTsAqICWc2K6pGWds7Ca7NYJck43jDrhIvAvb4NNU8ofCXWrmZ2BPCVXXe7GJ
FTVtlTOuE/5exXtWVrBsUrXTsmSh70QDtqmDo1Tf7HWX1VSnJVZBwsTSmhnUw/n4
Irxq7XnSxAsDdPZe4OxznCoPccmv10xJkboWccZEXCL4x3nKI664uZWlCYi1CKVK
`protect END_PROTECTED
