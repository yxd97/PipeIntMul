`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jCKPNQsjF/Jr/Hh4TLFz9iYROJ/68MnvjQ6ZqDBBnB8H5RcOCDR7Jkd+spHx2sov
GjRTXq6o6l5lY23M+CIeOD+fDQKkxkWJZclEQTuG9E2qUvLEaBGnADLaspjblTNB
DDusj7HWW+ZbHBmT68uIfjF4LwjaXE97zNwVOvBp1FeDwM/jb1bM6uCJUW+aeuQd
h/9D6a4Ghyo58u6nQcPJ7zGFQskeYozClGU1eQkqpeZGEz9oxJaifGcX6wN5bxzz
eEQUm37zR7CVzypBegM0EssoVch164SWLOeS6eOKvreADnLpxrjA/9yaIm+IaK96
l3k7pCfA6v8bAhqAEcPvUOXNXrVoq1CHRPW1Ansiq4DeZvVgT1hVRnmzDzdSp6eG
SkwaLU49p49TM4EL04txU4+cUpnq/5/wXAbHdtmxqAC9V1RRHCaAhdqs4v4Yotts
dPqRd0jLO3Gxa8t6KFR4dTRkEx2A5W8dc1Tyj1I4vYh8Jap0BrwiJxrQK1wNStlI
xkyujkKnnPvp6eaVEPtBrH3eNhu0nXT720IhK448kXCRTu3oeynuxy0nI08Qp/nn
f9/IzGEaaiEKMSXG1oSAr0z2bwEko8VrwQdd/g3O/ntynWPczz12mBurcz2CmWkj
zvD3oseF4Z/WibtZ46Pp99uY4b0YoAqr1NSgMzIUSZc33TGLRKvukNhaIgFSzwhZ
w7AY+XZHKd2pAdL40+ktMPKDy3/3XVFiPTp1Ue+iEmakwzY5cxEisA8dMWszLMAp
gIKVCU67gdr+42YIkvPZNc3vXFisvnEy2kwr6notHScOZWWDaKyjpaJP+r22DhlY
A+dit7F7+ofcEthAoxDRLVPIvutTDcKAJ6CeK2fc2+BV1jFCzW/Wpz45aFUcOn85
ug+JGE+8JTLLPrmEC6yVksQSxkJ6dEpwaNGYNB3lxzI2qrzbSO42SCx5etCU3x0S
eusPecyZ5c0lpaT9yY7S1Cabnmf7xHCIojvXMhaYYGd3GNF1+rcC21Ynfs3cXyeU
33rKUz6OE7RG92I3HzAz7nB6mVmGlhTEEvl0jeEgKUj4Gn5GSp/ssEP5q9DTGua7
VuIRnGBMrqqMR6va12pma4k7AYS/2BNNo+jKuOkWgGDKvcNj72MymsRtADEmUutB
LbRH+lVISAalOB3EAv9aqV+XRTMcyi4/OLGx/UxIyPcl1sydPba8UOhIcm98jPx8
h5pYEZSW3Y4M1kwlGl7UrNRN+eac6a9vGaEeecmEIfVoq+7VjDxDQOgm2odWBU55
RD+UE4R3DFi/ccgVczPdZQJVKFc6ADaCVNd9F4VBqDer/4LmVwYaDLeW/4crGGoG
A/+OfJ7MTGalHTZ0Rh3nO21TslrZkErAQ4E33YYin9rO65t+ZxpDYHdFlvxYBttX
lBvMkdg3ge4R0Sug+E1NldtGt+f8VYlh643Fry8kxMmBJrQjWwEmOyLU+E+VJuAg
3KGO6r8XtqkQ8Ki0mrFZUxj6ex9Vrs49Nkj/sWtKPnyEGo/BP8ENx7m7zbxRDll6
IXADktbYKQuI34eLtK9vlxrO76MiYEbC+MkrDHs2KfWd7LcHqRo8m2BSYN7mySVg
RZNZfxksjIIxHuYObEavzZAcBSapGjGFskodd+6s81kgRgDDkpGUOUFf5z0+iXpE
aj6HgQBlzBsM8ozwE/rSHas/KyMIdkfEwQ+Z/3Tu2x6foBSZsGkOnJJfdq8+hrEH
6CCnkkif75BZZkUROtLbOw1pXooakC9YmvWKBcpwE8Cl3uyPm22bjmh3mG+811t5
kfNVsVq8OlPNEY5QO8OE3uaDlsFw48EINE8gmtGbUdSx3d1PMw4hAo/EmQI2cxtT
Q/5ohhDmsZruYsGubHjDLaEifOgclquTmG9YdUhezl5I/igtadMm2wlVN+AMFVJp
Umu2lOCq8WPHu62CM6PDqKx0AFliIWAm7G8lrqdD997QBcqS/jldjgd92CM5NauS
oAhOwVaDvh3IbQ+q6rRPBjg5WLE9ofsBkltx1w2TTiN/K6SoiqGs3+tUB17B20GI
ASMSuGNxfTrk4nl18o5wUf+K5hTFK3LTeAsHUPShbudW4vpVfwDIPMBeO5QNpM+U
02E4orNPBm8LO9SqUe4MbuHK66G8CA0Z6r4sj31xHjpj/U+EThFi5gi3bXk6OEhv
3UQMC7hYWoLRMULFX2fB0y8fS+Ig5fw8KPfBdM/6ysgwcJj4OO0rWxBeYkAvi5dp
c2wnHyCMu1qDJOAtiZ5Qj2db2c3rXpOiKBwiEfpTNJmBvnbqXff+x85y3GlYI4ut
TfBzUsXbklUJUgvWnq3THGq7ANhjfdD1DiDS9uYGz3onQhD57xk9hB8afoTpkN3O
tPbQGTu2j/QlooCev/6jxVxnjGca6XKjvfoxMmwnohWjDHPg5CYUAp6sEDNyuDMO
hfsT9EOsC2htdm4QtT+p3mSlhHjqicXNx0uAUbEPC0O3lQTN8yBaQ8xbLV32fS1/
pgIeHFFmb+NyfpvzRNecCRMgeDWG+0hRYa/9AcIX+G+y/7oQRoMj7WiDEe76qVMo
UlxqMTULLl0iPPasFZmAPlsUNRH1o9QA3101a55dSbhCj0oJpS5a9DDRI9buiDak
fnCAAqf6FNM6VVPh7fKCMB/kW5gCLG1f7o5zT/Du11e/bRJ1/F+RTVAS082u3hvg
dyvUC6TB+6fm2jSBNDU8hkzCL4sfKR+MHv0NOkIwlskKyKEZXURr9rT6+YmEEUrz
5MfzvBOAv4gyfNMPqzhQLEmfgNJz07TeO/PiZRJsbxbGyABZSTW7HKA4W5s9jGeU
ZwRw4g8pBie2ZTAV3G5DlP7Ap/jioGrElU7nRTsTjhvKijmlQeyjS2Y/Aon/myYP
hJB+yHP1+5ovbPC6xHnFfkREzKvv4H1l8l8/EmsUFbvWX0WMxsksVZW2bfaziFmp
MMEHeMHpBppr7MEHuUuEAz8XExE99IuLKWCk8HfTbNcFq+gqJh6eEmRwb23RQdhm
M5mXre7VZ11Ed86V5BchiZ1EgpHmFZ+iocUrMW623bnO3eLNaMHEbb19Ec/ynt7E
M3ifQ4X4Wi1OOTDe1j4ljzir1vyngpcpwstYpEvVaVlMy58T72oyajstweFJX7h/
KG/biKC2u7wihfbsbIyYVXvg6lSPQiku97tRJ5VEmZStgevMwOHAOdaApc8OJMe8
QpK/8zp63DGKuO+wcpwulNYYJ2zHQgoLRuiITEeuV1dyADrG4JydGoYdf3gPgig1
HUmqZeD3SC22RShFKdl0/lArMzfs1xi4C8gQ6rnhwXRy3bVYXbmk3VNDDZeJ9C3C
raI1ljJI+qtk5zWcSqzk6N0O+i3lEMCeLazGMca6NhthND91qyyqxWspd0uZd2xD
nQ19Vvas28iefJ4Cs5/xMFQQASyoyA+7HsRv+Y8DPsedmLbUOu9BgqCEtuKwDbYc
+7MMyQnAzlBTLIHojSupGX0aXOStKrZ1AZwbd+sUtnA6w159gI2URFxZtyROat31
Oqk3VbS0YgEB0UcMynq9qtt6Ru2m6xnLjIUYdOWtPEUdtnAVPDfmXWMoRk1w0SZA
wx22AfhnmUAnoeoMCo91GZq3m8joQRK6r+biZsH44guvTZvSBgrWseS1noZvsoTL
/af53zV1pcEdTtCo3qd7vsTNOu1V83f3rZZRqhaW1TYCRQx+7q22th9YCYCdBBUe
W6cwlob7MLnPTHbtVDchR1K8WKW2iKAVkyAAqR6tXjC45B2RCpNxkKTdP/IwA8WI
7GSRXu1iRy8VOdS0Nyq/5FNfxH/oQuU5KpOlAVXjX4jYF546DHESQVWcEZt2j78N
9fokf2wo9sRf556Nowb2LWKuvJcT5fmOVAF2MSGlDRj+utNbHv+HNM3qXaLMqV2x
uYOv+GNs9XPWiC+W6gbNvBGIL+FaEsv/Q6xdh8RAXOxFHA0smHfdZudp/LlTszHA
I23fdjcbEDpDkgpee6KiTvAUggmTnX7BmBtEOg7pHqT9IoZgCiqWFkhaH5ToIjtH
S3J6N+gHwoAbw09KhRTumIa20PQpagV2xI1ihbNY+Wdfy4/QU3xIBQOf0vQTZpD8
Z8yHWtT9lac64QESKVVM6XfY1Q3YXb1Rfdr23xyRRhNU1wCXqo2NcfUmmPVpYkJx
6gRBkoI3+NmhIbfRPXZlu8IG3MhLBPFtfYaYKBtfnPjuqINoHwunykCEsLyrP/hr
cDFZVWImOhkNQ5AWvLaq9uTeuwAcKTgaVbrlkR/zPrxEfUswf1oe0b1crPwCKqEZ
vZT79ZgbCYErU0c3YqyVgQ==
`protect END_PROTECTED
