`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l8M1RIzb2gfk1Um+zFxAWa3Qn2r7LDA5bWmwYwvUcuSTJehFuBU7BAXVtp/ZRlIO
t3mFPeEuGGOG1cnh+5pmaf6ciTtyGHChyeve1RLvTfUW3hZ5VkyAY+XmyxG1Th0j
Pt92fmxsTwE/xcYJAIBEbWOGXNqMKcASRoU+8yxfJPVinc+u6riDZesxLTvlMmR6
U+TVWCjTULAoJx/9dhs56SvVATH92+bohz0BrK7U7brT+4lz3DW233EHOZFG0xiO
Vkh24tF/LwJSe9HWk9lwd6+CJGBHad8bia9QupZAuxH2gKwlqXuqrSeIHOixrCGN
s+ztgoE0qyhNf8lFBvAZnT5byeyXRwOI1mvVeVezZLsNOPH6cjaJLzWkxj4oCunz
7epgCpN9BPlO1IBOxHuiyq3VQWFB98nb+5rlXdqlRdgjfofQ4JzRpvyhzbJDsB6T
QtAWMSajrcfO3WpM94e7PKmWAceQy8bVn9AbQ+wGrHaWsmmeyzoaHJz9V5xJHED6
DMPTIi6yAy2+319TSqlM2IPq5bXUKRwZ+t5otAsmyq2lzQr29VI8F/hdI0S/CUoz
HFBdSA3e5Ffjw8LckSmFaKFkqHouoW/Zw+fzMqD2oazTJAlScXERZZ4uNH6AmEaL
RjpCpWu7g4KzZ2xefYpe5gdE0voAROXGOIlkpGA5ggFV9kEdjtyVIrz9TAB4QFag
2n162RXp7xD4jRLJPnBS2cJLiybZDlhM3xk5ggeLdSxYwfjvjm4V01VcQs0/Hlam
dPR3UV0N6ygOH0jNuQHXvyXSd9NwaX3nDJiCqyyLbkj18ys6Oxmw0TqDCwkTbA4u
PGeZKgKUuTao9PFUg2/9pal33mt+cNkiZ+unGa5l4bHqvjPes0qqtLKcjQdW5fh0
XsHog4VQSQR0TlNexfNStHn4vlci77IjXbgjjzqY0PP4jy8SPjfrKtAXkl+LxDga
gKf4SRklIsN7X0AmMs/4tY6hllW8to5ew87+OE9V30pLTx4i8Sx7gnaUax6Pr7M4
aQyVMgZ44qQFt1iSiEMRlakdNXXFsFNLzChIz+Y/mbIKQKRNPaRPBJf3BjTM4fgI
gSDBJDqNFjxmhWOcK4l1g6IkFphYjJrWwzCEmyk167s=
`protect END_PROTECTED
