`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcfG+rcg7AUyCF3Na1k9olr9tjYRBagUDOs4QfX1RSgiOjkBMLryyKrfoeJCp/Jh
c9zAYL9NRfhKh0PHtG6Km3oehEmOOw/T0PY8My0wlSZJntnoILKgn1zVRgE69wfl
rQf73F40jyKrJ3OGA0n1dDCDFMd2ceEiAEzFBKKX96o0fue+WWnusbNt4iAiZpQY
66hJuFwbO1mkdoDs1tj9IYArP9/znXdywgAZ+ookF5Z/ctk8CGWDmaBNL/9CpCdv
Kf/2konkCITd38KVLR2AIh2NXpKXFDQBs/oqgyUzn4lRor6pBTvQrTC+iH1Tb7Qi
Ze6l0PhDLEgr71wr/OBnmgS9myWNfnVZ07bHtsrDwqzre8BEBo9VNDHuJ7+09qAU
uGr72xsSqztVYa33+w3moL5eA998pe4ol+wj+vb2dc3zDCJinWQatcQo/MWzK9Ch
yl/OMRCwLSOH5CgM9iOQ0txv0KalOde35G73IGo+mAvysC8n/XoBOVjCZ1GKnrM/
YY5gjjRBG8G4tDUcUbCbyz51gARz7bZ6wXlNcVCmrPmhaJ/AHfKb7RBL4wcFgrjf
+Cu0wnwKcvqXQfC6mO23zA==
`protect END_PROTECTED
