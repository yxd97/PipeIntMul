`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y+mP4NQL7AiIQu1V6Dc5BVnfkMi3eD4dDscdGUtNv0hMGulE6bEaEjgY39Iv/9sV
BJFRoIKyu38W3zHL838AfWU8wW26KtYjfYPZznOzLEjPGd5pKoWoBx/HY1o55w0N
fCtWjRWfnT2PtvLPmtzYbOZC6Js1FK6zvhe9joOF/jyfKtqVBmcTW+uA3LVkRYsE
y2mTs86j4X0/IHPord3NxrqKEpykWnr6RQLKbrlIMnd+CRV33wgq6L93H/cFPgLL
w9V60z5KdKEFU41Utqx0BbJCCrAADFt+eVhLTw0W93EBfeL9RQce7Dit/0zvgay/
DOZWYLBSSCtXQAgiU/ux14dxUon02lFz2vU9UqOOUyc+K6w6K9DDMTs0JfjTYbFc
GcHUdmGyLRugMQBs7qjV6lGa5Gsl1n1sAq/Q2afG66+xezDQHl++5IIfQWZXhmhg
8WJNfdNZFiH/l6yP+BjVyhD9H2hgHpR6I/53AZQ7CkG+Hl6susNqXZF9Vn0vZ50K
Z3r6ELcyslsf4/ImQ/iy1aMbxtzXiR2CQzxsfNh4cW56dI2P6ge0n9ZfkF5d3KIl
WYxRgl9Je4wDHmE0ipjl4lbw1OjrPga1bYkGqMDm7lU=
`protect END_PROTECTED
