`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZTHdomlK5YtsIiBlO5zduX2bpkYrsw2cty/ezO0UXVeJ/+8DuCPPgdLTfIO1jrS
x69THtyWsj0IqIWe29HOI5ahLT9BEdynI1nljQhM2Ja/DflbTMJHXLfbTBU6R2Pj
IwwjuwErRpvcfibcInaRD3J0sW/ppp84ZFxXpZ3emGF7RDn/bRPKbMnuwVz6RHy6
+Vb7uD4QsUeZgMrasghdYKld5+siUZwmYLXCvQvmlmJHTPuF5CK4tMtM17bxe5lM
7ckDWf0mEjxRJ1K7fM4L9JDcFAXP18aLfR6kp2xf0xUoNgUh6CnsLywmE4YgMChx
1JvS25tWJ03xER/PTBbM0Mys7VpxnkQcnFgpJ0N5bX1kiqrPCaWB6at4ya+VxhyS
cDOBFqv3QJ51YRSJt2for34mplb0dfwLcz1zpZU1uk07UKCdy+gLIaWd4Jhu/mIu
aDukS3jpDRVTJeUGF/kldnLzIokjQkozyx+Kgcuz/qSH6lBf8YJQZleV8BtSamhc
7krxFGSb5GlSQ6pXn8oiyWeHq+bnlWIPt6Aoxf+WWIXoG9NHwC6LHUFMOCWAsTsF
MBQIn8slka8strVXs6JJMw==
`protect END_PROTECTED
