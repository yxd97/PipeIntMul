`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gq9kbbEMXnZwoFl5AxJXdum2JYnffHva5Kvgl7RglRLIpnqRSDJVfr1GHUk2Sogl
Gjt5V/PLA1cC3BrUfidUvwfjlRub6NcDxSgD9CRzVIfls/XPW0l2SC610Jq+SLtw
wRsrt2hGzypbIRNLZXybw5O/kT/3M4R3yTZXoc2bzrh0dL9N0hRxoL3uNj5ECraG
ziQFc6o+ibMEKvSecnpI/jsYHlIs2qiBF1iGkRN0xqLVAQKsUCQuNitzH10tm33g
TxPcZha7UCkYoEn70iq0wQlWhwjGqZJ8j6V7fD0ZYgF3hengKsgZ2Id3Dc0s6MQ0
4IyK4UYZ78dEmJM0+GGxpYU+xy4A9HR+Uki7V5ALoTuXsFazow5V9OpA0QF9PHqo
lX4KDDCrxS8T0/dETHRyui8OCiiRSS0wr8GXk75YPQa8ivQkCo5e/ZC04JqLhBAh
eMhX8wgRa6PfbmPKAi0OdIUOGZIkHc7aBCI3n/GEBEI=
`protect END_PROTECTED
