`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cTXZFrVK4YQLl56Z61FLDMFEIMzyLZpkn9hdiKCY6Amz9JilyrESo2zGXauCkyNT
ZTwimfwHn0AZfPj+6UoAbXncWKzYitnSDT8v2TOSOyOk07a2MygMXkbgzCXztEH5
EIMQiBg8A11zDAbvlLbWytLL1ZKgoRF5b7q+GZ+4iu5ukhK9+4DXQqh01jWSZXBt
eJR5AREsE3e4wpLdmbwPqZC3MGMxjAUvRqaw4sy3Y/snKc+diJnYjINjvo7Q4gES
/yUtH8QggbsWeMsoAPqqKiRqTDXJz37psOboE7f+c3mAA9Ze4Su3ii26/sIleDtK
B5RN79qYandWyWlfNX9gqMIHw7AbIjWu7N53OId4I7JWzfBWprNPWrkWt4jxek2J
z/TXDWwIouoL4nOzn98K4S6wzsXIpHApJ28DQ4tyKIJNI1qwNuYin1ugKr3KZFMO
Gf5nqMcVkjGWD/Y4OgIjy0ld9xBHvVnJnT7NhInm/PuBvW8F96gfIgkH3cC7Wch/
l5BaKjeJJpcQcEegBYp7NOp/kxNyf2BqnzZd14zUv4K1PX5mnRrr2cFfUt8ySwbz
liVK8+pRAJh4mRLm7wmZG0iCCBLIw4R9tclJx1z5CBl2hQtu4IqfcwYiRwoDis3U
/9HL/NrL2fBIGIkE8lnZKEwSflxyCMsuGUolqfQkkwmaaPboNOgJ3Do1/S8lEZqY
l0vfg+3fKIojyD+/2CcaprxgetGwJWxMxdzvBnUTA0iMVYPk/zb6MwthRSGYIIjy
IvG+DAF8UdVCkC0JSQPyUX2rmpCp8M/s68LmWdImWslS1A9qGoDgs9jiGLH6AcAN
5wAA7gt/VuzmFQcR9J6c9uDK8Hc95j/OjnQ09zH16u/QRpDyI1J6Tr6BQTIl+2/F
7eBoCW8PX+OV4oEcZPcTN+KmsaYpJAao9wtPYFiWRcF9P/iVeHTQTD0d94A+gAWI
KDDhLHyLhU7aeLGhkSmozBE5MEMV717WSOaSC1hr+nwoDMtT3hqs3JTQnQDvTtsZ
/gjuuUKh63QhwrZzD1hyIu7CgcCgU9VsVag5AFrLfpv1Vun+IXeRkTOtbSjR6dXB
GMqDZGZ+KMBEDCXdJcV5+HkP6D4rqVhBg2hNDM5pTWDN2mqfWH9wPS21h8Z4UnZS
yvRoxZ/ZUijMPU5HJdKSPEIC71IxOVHgTPBBmJwpr2o=
`protect END_PROTECTED
