`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9pESrlUdTcryv6lIo5zTBUA5xd0ZNH8Fx7+hVWWwksWgSJroHCLegjQtgMQfr71
w1P3/T7cfubZhwC+YrSr3emqeLBFDaoNv971N0p05m8wcK/duRBqnIqLiKl7kwuO
hwM5FE8CX46ZZvXYpDcEXPNK9gKeDxNFFcHVF22+yKFibvpkimMEYZwVKYYVeP/n
HBtOkwUoC1whMBl/ojFfJYFb65N48XZucyj7h+tjJNKXuH6wWzrMNeVk0Q425AQR
Z0YkW57MSX1PJdmA7K9FtEO/PxomuOnl9skAYrOUPgRHQ7MOMkVMRc5rhs3CqWHW
SR7+7abjUuVdRZl5FrPieeFfkr+3bVzCjq7yE/ayETBA57rQUbWRiDS0tNQ7n3Hm
EHJGqUrZwqvMbw6wIIqQm5zbdyIv+zWufNtMsr25hQxYbJl/fIkLTGwARLVOOH4m
ZZpY0RMBivQx1V6OOV4sFshfbwUOghAV66FAvpg8ZJ2EGbhddWBWymm9WcpOMVes
WGhLbzJrCypeUdQQVzXAOOgZTu/8H/vdaBvkdI/6NsY1K3xMmZZUygDyOJzUHZ2Q
oKmQ5t9hDczEM7mLuZmdIV4uZYXI+DAAKrYoS9rnDTmLLO8nqhO/w9Qykbafe7LC
BhSCeh7lhoCD2DrGCjtN4gYgidHkEX/hj8P6iJihVi6GkKnS01KqIK2dYUN7F6WU
LLtq9VV778PT5opzKjwGuXrhySASzTi0yw9A6FWteDFrAzoe6HtsDAhM+Q67fk2w
yvgePPoTh/IxA/bw6ZHc3FSa2h7nIzXa/ZkfFqWmCVBhZwXgQLyazf/iSyo3w+cv
G4PO8UuT2KzPnE2tb1cQWLwmqW8ivMeXBv4pOGVKWXCvDHRfIjlsH+8E/kazicyO
PsMRNt91UevnfHosh0XOqASao7cWRh/tlLEMPJTc/qCB7iR6CeFvN5UoLpq24p1g
88b9bc6rnLg/CtPR6w3LrMrRZdq6rF6UOFM+rVlF/oU=
`protect END_PROTECTED
