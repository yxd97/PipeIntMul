`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XhebXJbvv3Fn/Jb/q9G8Zv7XDRdbp9nSZe4vBM8dOkTH40yqhe1nBD1yWGh7WHDp
u9kYQei79iHzb1SGKCC2tlCQwG5qFgXNVc7Y67Xk6WMBttLNBHrhVSMEqFLrKZce
GA9z1X6eCD/UZHxeo6en9W3edIZcb+McTtQYJ6w1lJGxjpnV+oV4SUY6eMQCQjKP
EgXBRGFg4PRfSPzsa0QBXjI39a1+xO4ySrS0Ve2yljJ+d3VHMsHKVL8W0Rt3zFPA
2a0IBcUjEu9Ht6jQYkERRrjkAGqKRapu99O7RvFpafosb4xsb81Si5iH7hCxJWEe
m2U4+9MQUQWHW8nTjqyYIt0pcIbY7URmqzB6pUpX9krZxMFaQP4M9QGuc21sSVL8
Hl1TqT04LODqxQ5CFAKJEmddKn0L43+Xl7VpYNJtt9M=
`protect END_PROTECTED
