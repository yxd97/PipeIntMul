`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UmqORsQD37pjeh3tKd7wCG3ZZkD9Fl457fR8qOkDxrEn6OUK0OJRFNuDPyHXXZ5R
bDwMgNp1c/oOfp8QpCy60zrC8uNPjfGEWN1089MhXx33U3fKDK/IXKRboPRFk4I8
XXHWoHu9QBg4fRnOVzkHEh5rQ2in6lcK5uSZi78spG6NrwJCwuKys4vEWYTkZwP/
T7vNG3VMf0C0hshN0XM5IMXzRrOxKIUmGnfCYkZJyICryW/3jFuuavVSiiOBRl3q
JFWGS7NLvpWtrcKliQBdoLoGZfD0HllzobCQz5YhsezOlF5vu261UAUGHow1OQ1H
RKqSi8O5KxCcD6XzBMq0g92D8UaviCvH32ROyHeGhlpyU7GzL9ESzTrcSFv2cQmr
qK58OzhRwXEowjI1CaAPPYLa13lPNKnBUR66RxTPgaLd7nmxYc6ArdwEJZdzt3+B
2jU4dkCVkliW3qc8hVPmpVSwgKhkl7pVvqZPFc58Ij6OnQ/S25w+z0S2wQhdsvwA
icNpQnaooiJIfXcMwImNuYot/im5Cs6Upa9eVja7GkI=
`protect END_PROTECTED
