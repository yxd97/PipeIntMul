`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fAzSwTiOhbOASZ/H0neF8qZc7ElEPRZeeC0iQdEc7h/PRezSkw/XXnebcbF4aWkK
YlqwdeRgDJmNXETMXb28sG3Vg39xkAviGvWixBpchdfvxvq1TwDyU+8R3yd6S3D0
xQHaHc51VJznO3l7J3GAREd+CTQggBY/s179ViY2jtA9rAg6xemb+Jp6vkivjOs1
rgqiSg+LzcYsxEVbWf4Zwu+ldUdR+Pem7uIwOFe+9e0eymjtjI4+ixz+YkWzBp8l
aNWr7s2G7N3pFxrAQOz1OQhIy3xV2RP2sPER6an8GoFT5+CZC4Y063O+23Bzl55n
WPx/FEmqj7aJ6Vvl6Wpsera4RLp7A/q8TNGeNvvoRyeq4tfUQW0nayvsOsjiVYm1
j3fifwI+L2aKXXX3PTFxt4mB4Eih2H631UQdRsIMAJ41omh4A/hDFTdIjcv2hAhf
Nt6H372Unaxl+sSJH8HAcD8u/HcVWiOGiBi+d6ynwsxluU2xnz2sAOAcAJ8x6uIy
pBg4urpOsnPt5aIP4e//7X6GoMo8gKi90TDr+eg4ayN4Bze5RbQdWVSnzDRg/54R
6Gjm0r3Kt8X6iryz40pcu3ZF68OAsYYm6eMLJmH9ukejLyieVAO6KhTh7xF3g76H
HakNW7wpVIct9YR4CkSR7ELlGwI4JaBuS92X4cklfACfjAyRCsF9+//57i6oI/Eh
WEqv15oDZhEwBLi2LZ9dPLlBDE5lZZNbkflsPt9CtcrJsNMk4MGQ0NapNnANkPNC
6lvOpQOniDY1338fGENaa3Jkq+7WyBEQjecNXqhdSKlXEiauHXEZHEJ8+WSmDVp4
P3ADfXDDkKtNSLTnBWCZ/mJ7yTg7wd251FLLeE3T4FwMik0iP1MV64aljyKYRb0k
EPOGyHQKii6CxeMkZT1DSETuHzjqHnpV3rt5nvkFl2UZbNyEe3Fy3CrkavQQOeaO
xFGUPTrnFIVKmvvWrfqCWzje0FkQ2Hrh9LHxan3HDESL0r8FzXYtSz9Y+DhLQiZm
CiGV4+juSOEyBGOgEvXGY/z2+9GnHiDye3FByWfmizceUsYUyNEFlbs0bYR0A+C+
DFR/MsqNIPBwIeeLeIPBy49ptebON98FaDasE5bXlKYQQhdUjFWrHDeLhYia0Pgz
2xuWRmqyQ0ZP0S8LDoR7M9aLXBhB2O7dteZ5TOo/B3FGMI2Rl4Zse8/O8sNLWZOq
TGvV7AWtaGQantAv80anydRt7Ycijcfs45/+sMb0q2YPBJKh1+Oes6YiEjqa7zZv
8X3oFeBeWqpJP1BqReJCIc4d0BzyOMWayY1TZvLpnKW4GIMQTS96h5XMU5bNfoDn
FEa3foim54zc1b7jdLcymeDN83x0H0ldgMnkNnEYN5GiZ1suT8fXh5Bj+jxUA8vZ
qEfNKQuIrxeNnQK/ZuyZ/MC0pr8dxrF25zDM1THmS08jq/a7zol/FS+ugIbND9tH
cwlwwXfN4K+bq+ryY4bh2r5Yn9yAHeS2aCZwmsjkVr0NFPFcNRYd6N+NxG83QM2W
jkTRmDtuELB5xQpum2yAsp3e1N3bru3zi0facIAKKNvXxWbi4rfPaQWDIMK0W2ox
NIF/XTzmbkHS114cM2/DWXQhKmH9diazEAO4qoJnJoX0fcqQNnQIDMfADV8H7GIS
I5tQUt7asNr///TGWcrnDL+StrxKmgC3NZ5MfjQcK1zpk7TY30YxQJ403iBdUL96
r55fyzM8hckzrdPcJzPEGdqbimTtypYrSDNwjCfAwqu1enyXqZnR69DDsEeZIy8J
hNSBfiASKQDQy3TFd0GrYXY2hRpj1she+NXyOjebAua+g0k+qaUUvi/pSjmbrm9s
t7/Vb+j6GaUkDSXxkk+8/lDs1rSp6v69OjJocYpJVkxPoteiBkYCxrsDRFqss4Sd
83eJz6KmjlOI1Nzo3eVEvUcpdSJnvB7FaiVz4e/eXtADQt5c7K6pYnKX6gtj4vV7
ZhGJ+asEChk60aRS2I8Qy7Vuxr1EO7AfwR/J7bvdg3pS6S9rumlC3RwYXrpf43KE
/5jlj5zthokzQwz/0SEM5qAENwnLCBthTBFBlXueiidSH0S8xMEqPRrmepEfmsCr
zfIsiZwCLFAUauSbf/17iAvXEH50S7kGtjLk8Z1zw2rMDOsl8Lk9qGHAh3FJj3dk
X9yg0Tk5xSVyVfivHFHvFxU53MDNWgofx4jUE/noVBpSb1a/O0vzd32jlikDu3q3
F+h3bGb2nfZ4FJTOepTC4rvlGv/XmHQp15vHUdLP438KNrqJl3yheG5ybsvGsx3j
JO13plE+YMrDM2Lp6g1kEx0yhdr1tfmxkl+uftCQH1fdz+9giHsRvo6491MBzq0H
K01VL7kW9otu2Q2s0KylO3odGtGlnYJw2ziiAEoGqgAg4ETCwqX9nD2MCspM0U3M
23i2DNz3pjgW6hqBh7tOP8igCHkrm3jE6odLCA7X1sVmgV11dEmpZwbS9Ih6J7vd
l5P5PZonwreVxsAMGn4gKbpPig312X9umazVkMZL+OXqmrWm4/6FpNSYVORTeDaV
oNVbHqr72ojrn/kbJQjvvXPRcGpbsBvTjxC+RKYoHYGKL0OT5GdRCCih6kHCAbP+
SSQNfxzIj8YaqxCVfNw8wnigVlnaeuC8rcqGRhmO6ZAgr4/obhurychfQotcocwW
SJ94zIyKHNESS9YusBvU/3lxHk/bnPXXVF8pJd8OyTEaU3zrBA2sMl0uZ1XhV9CW
SraQ8UbLKRKbHD9G2KnUp5p73W5f+YuSHG+Wg11m03DzMYrg8ycJvn/A3YvXhGMU
KwCsTqb8z51G2+S3pbN4uxHia/Ab+mfmkzJtxEHR9s/tmRKTWN1cHNu+GqgC584t
hzXP0zHdckX9f6cnbwMR+O4p2H+ywIXLtHAYzKnR0Y9ny41elv+oN6Ci/Mjxvj57
Or3F6/fjKyCWQD/lj2gnUy4XNzWnw4oqWwYoRzgB9upeYa07amshHootcGWSn0F2
FYytXJ/XqQnqtGGMpPVTuUT3Odb8LxflcxjNJWPCPdEo0ET2itYESF28MbSvsY3k
AnaUMevlXniQYUMl7QwroHeKTBGoA70t+vDKnsGdGBy8am0NTrGIviYokjmDBcdG
pD6EiLHcxtcqQMGkr7WaOx8yanVuaH5Qn0SYIOhGJDLGd9lPDqz4vnC3LnDMhERE
VP8BjYmnsslPgv+iFIYAPqrXx/5TmzRS91xOzKDw0ZG8bmoJVoPkOOp2k6Qz+whn
V+i6zFhXBHjpBQEFFb0qFX3D4vLAaoa+5iOEQ7SSjNuJ5ezN7WJ1LN0vvyhcWMg/
wa2IUgia3n1EEEAHJgBrwdbUeRMjytYNia/m6Nn4C+ogJC+4bqQYo8SsH6h9cDG0
LUeKV8QX9fbDKN4FMMpftycSiIl2S7YzmMVA+2y56PH6f3UHbJFROHFT8hU0J7JY
xrr98Vydj74dBIMdXIZYdpGiLFi0MOB+24fZrfhGjw9IUZI0m+l8JsVh0T0nlgc/
Kfsl0I0us7fDJm/MUlOUcTCUlw37ctKitmoNWp0GWUwau+3Cq5o4R/fSY0RdD40k
wLvW9rQyuhBvK1UDE81mOJwpg9Y4MszSQvs4BuzlAxeK4R8rFmDmAsBQ6UU1pmsL
uKhQkHlko7vd79lxSOADoobiqlkMHuYHF39oMDyCsQ02Foww4s+EEDjmsCl0C12R
GxfxrjIuuMZ1R52kNRG4oAHYZ1sew13G56t/DHSBaC0NsnP8IU/cuBQzCwfntQaj
mGCVOblvbWkmNQpclN7/oBS/6pgMkIzgd7A8irqBoqAMUKF3NilRZ6+EGXC6zrzJ
sYJlIDH4rICyff9ob2m7SNTd+8hm2QZHVOz4o+XEQtVXPLT7imLfTpDAK5/exvQR
pRnnyaCDeoQzZATG/Wld8pZKtawni+Sm53k8yMJx3UMHbN4w4psvRFZWkn/CVuYW
uUf7cUxlqtbvhglkQDBs5Oecj5RUaPh9JFe9ao0BhAtSiuIGUacaBnAldbMyjgdb
ZPDeeVt4n9Ue7YEff/LkT66ez+Et5cBOOyyqlFUSdy70OcIAtK4t/SzJ4IKvNNuy
FUDV2B0G+uODwROpAqOR1mgQ7KFmItqqXeJ4hfrT8/iJtie8zXOrmx3uxKMBGGLk
+93UiX+cdImeW67XsH63CZH0PFMKjGy+6j7aPtemVH1Hcshz9l932NlvFWls+UOE
RXnWi36zL6lrHWSGCstEji+3Vicr3gnQKNDbOhycC2hQweR3BqaUUiOg7XlweTfB
O8K86rIgui2dm3sOCap1dU4R/ApHeGHQYL8e2zlUfgIAhrLn2RBcskXlLbPLvp/n
F1y67pDAbeonfYOfGoZIsZN4t6xZeBsOAPbHrlzNES0dsM/WLBisR98KvFqW7Eyo
7dH0JVHW04qxjfgLrX8xvyO6DzDT9mbbiqP631RrE1guozthrnpzS2QIXV67NgCk
1e8P5x5ebC0OuRuk6jeMg9SCYuUQKBChbwxvMEcfLmzKB1llsmoRKFPIkFVGWyzi
1uL0nnxaET8/8TVzWnbFvtiBAlac2HsLiUbpozhsOCDqlUgUjBREMmy6oY6vzGo7
RB9rFhLn7H9ukLp6k1zsb5UHa2uGshk0RSd+GGfzjkN8yxIbf7/7B47M0C6JvIDN
3TYbZ3wzr1ZyNGisthVCtJn6OC5jCD8za+t/htZELn1cyEKNXVkExyNaz3cQPNZc
3Qv9Oh7swsSRDqXwDVO7w6X0SAPR2+g+eg6AbKVi6PK+YLCjPSiCrW38nUjAyz1u
o8iyQvNpZmZlcaehpqR91GDSej6i7oLGpsuhX7cKy62NKeN8TeW1Uy2xHCocsCl5
X3ZNT1RPcCrz2WiHB+QwFow9iB59qw+s2JpsNTwg3p/0CCctrtcff0LGRdPnaLjU
vkAxmtwE0vRzvgb6nVRPmmeDZnCI83260unhceBfsKihWeglurjjUQzX9sCn9ASR
r3SunubilYOcJ4NgTgPLexnz1yeMfcIxWZp8iAJ6rMMThSu3gMpMseFnB449m7S3
7pyWaBnidgcLOVasJ4xIqRm2P5vx+77N41Q790Y58fAL6T3uUI1HZLC4uNi0fzWa
pExwCAIVSQrfNFY98Mkva73vGTNFOzperKxiPLCZOKeFkFFFI+GsPMKVQkDOsgHR
p7DxVoX0yg9iy8DQjMAY8k7OoDAzIn5ef8XEsh7c795fQtXrpVmhg+vbBjas/TSV
vSibAVjPTBBdFrSS4LzAygs63HtSSmp+/BUgRG/wnhaHYs4x1QVUCg8Vml9r6QO8
KKSlRdzMihHo22SR/sxdQ2DKjWN+9MTGgt/m+p2I3OB2aBWxx9zwrim7u/7qzuDP
BuOxwqh4mUAN2Gs56+dDX73EOHdhrPt7sfQc6X01nNuNIIXjKi7yXGqKsflTRg+T
wdK5ymL3Xkq7x/r3Al8d0Ndp7wDxCtI+BvniWlbal/jDJslAbqfb1MdMZ/89nO1U
dChh7PWeYoDFAjxbMFesz2aO97InqvhPaxVFMumhSbeJ1LgxECIYMxp6bADqGFEx
bQlKsFeqbSzsXfNPCd8hrQxoIamtFSWampGgCkDhHVgsAfXSGGw/SGQbpj/XkCf1
P2QxVuJZQ4ivlLiHhGW8zlP92HPnyfXFyyA+rXSYXSo0L2TzrHVp6DlJsltZuOaX
gN1p0SagYtLQRYskI1xlI8Eiie/uqC7RHzaC7cXsqVsfL5TIRRCpAdDWmsXxjmeX
ucFVK+9zSHWvdR2+Js4a0sXOLtP6x6oRvq2sTpB0Nn61TL2Vy2xMorPuZkcJ5JMe
SYyEJJduzwwHxzSi3c/YFh+JCnjQui7DYSiCa4ZZmOI2CryaWpSa4quc5gmEP0+b
wJQMbUevoVFFH1Ny/+xRsgUCjjAwS6Q+5Bleup6m6Hyi3v8yE5CTPoyPfkJTnwYA
1NLwLaOMRJyNAaRMyO7loaJm7VcCOYv5e8EA4A7MA+I0cYL71+TDAFdrUBOEO+0X
jTEPUdyU92h1blXieozOU86R9qJwJuIowzd9mNcW+JpkuJOk33R41ho0q+K0zZ8/
YUnR0XX1lWCF6V+q76CsQNiXowmh4poCOHLiywFT7RW88UgwanhYpnenL54mfhLp
oOZOafBTdLTMcjI5acufIHtrXS5rXXORV+Asm7KLkghO9xE/IThf/SkMWRZFQJYx
C7VHfPnS8LKgaL8PYA5PTLT7z5k6BSBKyQdPPWN7aUQZFRnAQsALH36YQo3SQC1Q
+dM/8WgBp8nTD/FjIR8WY+BuH5ljE6U5UVBEhDcZ+8SrUIiMcNVFP6LZC9Sr4/70
4co0Lg47Bb4mAtDeTCjIkedtP+nZFfhWX5BEiat3cwE69rOnaqDLuilqaCKJVwn5
/z2XhCt8VkuFDkrZBP/Ow7FaASbz4a/QnVJWtRGtGKwHt6fJ1nApbN6Mq0aNxtu9
0nrcsngHA+HXldUqH7/M0qqyHzohYE+GHD+7kKIJ5RRunPaQFvT9D8c3Y5OE1d34
dIPUrUnHFgn+Sp9Ala8Q7px7Oh3NGSYLRyguagmzy7an4pRkeRLtBD4LjoD3A4d1
mIMhUCwvSnYmY5p83kKPKp67793NOCH+wyJtv5YYWepq/lR0s+cxAzekPKexv987
T/IvXM5WaLHoYxjH/8Y4znJPNX2JMUD6qVIw94Y+j45qPh1JzFsOlty9EseAN7I4
YwJbvZ1I3G5jhtfXBayO5HllZqmTMgZwRg4qKOy1AJbJdirP7T55OaQpjfQve4gb
giiL/MwM2qOWKbtUhsxuaHDLHi+p4qPPUfClT4l1+SfCfwOTCNqizTyByF+GVoot
BaQyZ48NisTBk3HBlRZvYlx3jv/f4juFTyLVkyEHKWJwe0QDoIUHS1bSRlwhdoDh
r4lPJsOZfmL60Qo1acRaOYgkO4ZF9AL/s9MB5mJGcnK9JWePCDETF/ixHs2eVOai
cqiCNom8A2K7/INeSE12HtQYzahgl6bQT2a8sofIy9+VQuIxywj9iIVqC69yFjWH
kC2lwBkbK4YCqeq7LvNtUt4XPLd1QSViGTu7hWk3DMGXiqPJVuy/p/7FKznFrmmm
+Oqrn7vuZOVzWzKTiMP0pg6pVQgHFmYN+uGmpAy2piUBlurv7C+/q+/eiTbBJbhj
NmfUqlbjDA1Z2UlRV/9EYl0YJMQrX5QV5ZoZ3I8txM2T2ksYtUgkZtvCrqFr+LIx
UZS1KsYa/B9o2tbCFafNYJ3+l0cuiWnqT2/M3kTB4mQ166voWQnLagpJmy8Ee5Xn
yO7kKk/2KO2D03NqkQDha+lWt9wojVITMX8ZUaKgtuHyB4txqU5cs+i1dd2E+/Vi
7euQYc0D6Uh9UWBrHiuW3nd/DMSHqcFhZP0p5BDK5jyAWfAjazRocH9SODHvtI4+
zgyIrH/5hvdkuaY05BMuW9AfdmKJZROFHIoUNe965O9UcT8W8ixFWtdntBHSmCzI
Q/vAbtZijF122Q9FmjJ7kUP+eHOWGKO2f0/ieXPK2BKKFl9a+1ywF6PGkj3ngAHK
IViGMg7LNZQFiWoI4OaCmqbOnru8PX8AkEootfOQ/kh2MWfGFHbwqk4qkKA5ugzF
zXQA9WSMBqtXIW0g1r1k7QWmoSzJtPyQ5Ya+YPlJTaQE6CQILp9nKD9VUjZxwu0A
xglaa9VPtfUpz73R47zG9/pV7u8Z+rEjuoM8CId1/aTm7Q5Y5d3UUkq7K0YTPAYy
xKwZS0VRW0+La+YBcqTaO0J91/0/ggidZe40c+crn07DRPLif3tV6gPk/ujt3gmb
KdOvq1z5jhJd8JqxKx+ZGitF+Bg3P2a5/6GpUwSK5MqYWloyHtn+GSO8LpOEziov
yaKjYoWqIabdR0OGvY2oI/kbcNdu0q+t0iDRzmv7JvIvTf+h3HJ8stc/gH1t8dBt
NY+1N6ZguJr8DyYGvKh4sDlXaKtVobzMO56Odu7LyG6JdwQ2J/GeML/Kau23EaKf
Y3GWETmMrLeCB4twZaY4z21+phjfGqxONSl+1dsxh7ykFGG4dMZU68gCltJfrqzt
nB9RUH53DSygvjoAu8u7pZScblJNQ+mMrtuD+j5ozOdbH24ok7G2htjAhud1cRmJ
deBKTd7pKqNsFmx05pBb0I8Zj0y7XGOfeJ2oGeP0IP6PNQ0ujbbnIxwru4U6CoMv
UHWweAQDWdLQAn8a4upE65lNhCtrYSdurR1FV1VkeJ3XfEX13ETSwKrhCFaejXR5
e99yrgd4FUC2N4GzF2VLpxKHDKtffUnuBz9OgwQPDZw/oQ1TeXKTQNHCW+URI0NZ
k1VIk6Vw1Txg3JfE4zCKuWfJzsHHkMYbSLCK/UMNths6w241hN7wBjM9Eba7FZMJ
69E5WIvt8cgAYx/so02lCbKkDDQUjRPnqKK8jtetk0BKl6Kj/91vQGCe20kQ8IZ3
yw2KpuYIL8LHLDHU9wlSAQUqMy8ylh0Yg/6k/aUjQMhvGWIhYMpS9o/Mf/CjBU4E
z5Lo4i9Fd1cmSWkr4GSKiCMDxETKueNZjO6+4J6ydvm1UrGVAP8qYXTIKytpf3k5
Pk9IvTAqdpKVirM7wvgEpsGiPyKmajqlQD+xpzsGVr2L7+5PM960b01Sndlq17wB
OdozDi5tVVALzkokLcAcko/2KOLj7eFczGk8lQSn9cr8dYCF9C1U7Iar72gVTskk
sMDRGptbCvvrW+cEtAU7ePjZmJ+ceMy9ZqhmU56rR7T/1NkjfvXR0IYu/S0W5A4V
0BqVeoTqj9qIxkDxBMEmp3FDbHoXVBI6Kq6Xy7bj4iua/KRbSCfoU09tC7FcBRxn
KTD2Xe0aTK1I3YvwC2evRiw8Mw6e4T2N26rZzxBUVaAafnpaHYOLg/SbZ/u22JZJ
87DyZf7DsMYzGb5Nl7jyRSv8ckx9+yL92SbgC/pdYlqiDd1gzBd+1xVaeOD8vaFm
tloZp7s/nqCx1QyC4y8Yw/ren5mkhzQJp/c9GOWybrxCanNYofPJ2EHNf6hfXAMr
8WFzN9T2w7vHkStFgwRt1at+hyP1koZV18geSRG42sPYsyg58i8BUWhQYZ1zYGvK
gJLFG4SGk4Po55Qo4aUwbbmMmLiWYv0X9y8sJqZcBN5eMI+Up5ruVEpvz3x4VwpN
l2k4Tuw80ACO1KiIK3EfWnIdMcjlNDsWWF5bJrCy/yB6iPQ6OhIcZNLJ1FtENyND
nryd2xclkrXVXleqxjdFKEuoCYfCqwk6CF2GFHq5JbpJpSs5ewUukwX4szOVGueK
r4V3IMjp0Q8dRwH0UJWEvnI8T9odvpDc2GvmYTdgR4p6BA3xjeNmmoSo1ILm/Shj
rvN9oajIcD3WNvCd8M9AiCmZlUVy+I/mWm0Pr5RY+T4DeVW8p/QS7lC9PltEqGZh
412878sV5KmFIKeKfn2NUKFJWN92P+VLzbuLRjwdQty60o057lRZAgjmDAFjGIjJ
Gj+UWRv/33nmY/NAQkC6STdCXddnf3zpbXkHWe98evKfu7H1Cn5VmvXhLcw2GLXu
cYhW7+e8XIZrvtT4YyGla+fzgqvWPMeZijlsqaLIN+gah92IaPbrH1Imo8QNVwtL
qqRO6tCsvqiVi0NAhFA344zprkiPQnFOk78EyXuRncRq/JfdU/nb/jHDY/byE35B
ih7EC9CfLnOq5kAekbe3LpnyRWZ+NOrJMERyTO0IfMxCxrOhYE6xObuqn/Y65zBp
zGifsdi7LMPK0mjtQRqjDK49BztC4ROqt4BIqvTS+IIyuTWd6K29j8Eat16omlGE
pifD6TH8M+g6xZ5+ZebvRWb/U8/3GmmfcsoQ5ERR6s5qqK8BIVVE+0WLJwo95KUE
3lG5d7sDJOiJDoOr9b4wMZwZVQY6AQT5kfAv/0nDxH7L28lF1BtYuzXQJoKeRexj
7wf7Z8bOxzc7MAU/hK77LdfnxE5PQJ0bXiujitXdDE2XbIxV644QU+7qDz3eCa15
PUZY76m8Surln5/sPXord4S25ky0VmSRcQppkgsfjC9ug2oOLWefbx7kA9+w2NdC
qwT0TX8UQFsNjPtav3drbE9sYiw7um5WAbd5xW5GR6KI3NSvC4IcQQFUPqA6MIFU
28bQino6ellYlEc4fSSSD7088qjCKaQT6+o6+Xorv6yDT05yr7aeMe3DB1b/NRio
oJfE5oLE5suYFq44GLyF/CwgObmGHbMC+ICr+ptGMpxbCVHpYnH3D3W207JWiqO8
IbOKfmpuElqFeQLfS8wG7yfR4tZaezzNcFwjJ8IBpOht+b+28asq376CWTcU0uw+
d5HFw/E5HmTFhSLAxxnidp9Zvd03+pJ75DOo3Xuw+27nmYrcrXuCFs2zjF1DByoK
NFCzPVsGRMfJ71oGeZKC2tOxv1HPOl6to0wY0dJsdkW/jfvHb33H9O8nOlZISF6G
MQ8pNuwddiGIKRS5QpncjB1eJagTpsSCxmX7GkioJwypSSrmduQNDDAlxKYihcDI
MBpbthichsl1btoR9WhLR1obA86w6NdS27B2YjZrYY5sKjlb27P21CdrziC2h85M
77V0VLq3cbby82htV6mKCvKWIQZaIEdQZoid+RL9HY5BikdPAb5xMVQ2WUoM8u2x
o8uBRLE5rRio2b1aKHY0EN8sHaCbQQQBRC6ISsBnMnV5doZ8anX3fp1g6HtkUOL5
U7mx7/dy4QII87leAxquTdgLjNOISWDJg2qubK8bK9O3Q07lQLcqMVNURMqn8qyZ
g3REu5BREho1ZgJe2TIJwQvCh1xCn7awFF/Ze4HBQyIT5IIL9RwUT3xiHRD4icJD
vyyFvWCRJjjjldrtXr6Npu2SQpRYbaGRaHFmMv2jCp14HmJIap32A6WNCz0I3loY
oTheVuNF/T/PFDhz3y88rVVcaWHPI90qp7aH9VokFmc9TtcMfsV9s4R6C2iy4uql
S4HMAgw7aKoRGr/gWLoHHYbQFwuGHoUyOIuATk8DVU04fcdrhBrF0OWEIwNhycFH
Ly8vQDLQp49fhxsA2bxW4UcD1xlDnpE5xDv1U3amIddP1G/T60DyFMlbll8xayto
LZs9jbIPBRJmpLzmNvifTx5AtKCCSw5snFfeXAPk00jYBtzLkGVWq0gm5yjVjGyq
C43EP4pluMczcyJA0ceWjzZotvprUqK8toGdNZKu34X1VOCe+AmUT269y9io9xTU
23Y5Q7RM5cAoBJkUu02itvwL/p13WnHY5xwatU4LcEfvg6XfegTN7Vb0lXrlEwW1
kGib8zbKJNR5WsH6wKEAOxvdUNyl8d020h1bRFEyAFJadFEPLKyj16gC2QV75iy1
kJ4IJpTgHbhEvJPBF51AJd79qpIYWjFxvdVc0QOHlAsqg5zZtafWSG4PmxCQPZp1
CwZmJnmxS3wyIeZGBLZn9Y/dLLFuaEM5ukFBCfT2I8LB3FynA6gYr4LAe6t3BSwE
b+DfninnC5Ip2qJD5q1ynvx07m18hj6wvlL6unTYTJ5yDwDwDGVrqqbaahs/gLvz
FOPFbNThZkTIrDgLPcsC1mPW3sNaGqBA/9+XT6NmVxJjHQGb7NahKzYWXNQ4iNIS
U6VkFp9hn+2iFFKp+vLFVpLqBpJf4zEqpPHuUijBEUnaffZY4qy+6hH124dtpisX
/nG2HSUiQelBh6Ch4bllYrG1fcbQFVl/cVzLv5Lwhzmgvz5G+gADNj2MBfTxewQf
J8g4uOKAK6CiJIUMPoetSY4d7O60dEzpwJ+mc0oFRVaB76+rY17IP2Gw5Y/bx+9a
GlL+5ZGilIFzfQsUD/pgwSDuTtNToKlsDRtbowWdgpAeqmGbUtsikTd5/dVDzG5h
0CgWDHhhfHm+XH/ftTQPZEeHuHxXuItBoixntCGLUGzXDmif6oB8svJn3QcVdE08
tC9lcOz2Qz2Y24KVyDYmd7Hg4l8+rrbt6g0Pi3J6NNnX7LaZYMXE6nIfJnTLJ0A+
go9U5jSRk0teAgjCrqRxdsB0042fvxvomV3MgUyA6QjSftx13hoviH0L/TMoA9Mw
DStz9xRULBMr1EZ+ZsktXRxuCQR9zIRsQZrevrtj6F0gcrXnCzq5Uc6ybFeYvpAm
n0W0X+wyXqbFLeNRaZ4Xmca/fbKDUkPQbgTVAtnGocruWg0yH6WNh33H7jIWgLXR
5NK1zPSo3oYCLryl9n5V1tBNM9wYs87+PCeJQNkdnneaUk9capcV3dbqG7pkizSy
5yNzInN9eIOdxSkd7YYMIDdk6TFOq+DU+1pHwLOQmIXc5ncTFWxL8R7tidLrgzD/
nLUb47WEOHSreKkVhQ7DfW0EmaaKHJTjOj/SYZllzljdOlm+e5YxdWA5Mx2c1YJ8
cL5aNGHAd8urdLEKwHfbf0EDyl6/Qi2kz+/IBfQXVBdaCOYiofUBVduwddbegUSU
GibKM24Hxt8Loqn/bCzx/UalJ1s4wXfGYGMMRbOmB1cJyfcrTHuVvpJDNavtv7hB
O3wwZ4+FcELTS2/az67E9UF3f0fHrZw8LE+UphfpSGsymgH3uL3zNO61Ma7YZWxS
9EFeysVDr/5J2foba78bhf1/16qV0ujAtUJl8mPtpSyY5JhuIWBzoYj3Whx2CU1Z
MgGYEfd02jbHMBU70wxtDVYO9njNN8imUNu/ljwbLvJCIyDYoCgAX7+5PlFcskn4
Mgv/8sxCPtOew8jwVIvAikpdpqMyF6ezRHEcjra5ojPjQK39QA7c+mH04vGjM/rS
5p4TIcrFRZWGDf4ly55REC/YH3wurABhDXo2ntQ0HIsJktPTLF5F286uU+lJbCxn
HwOCxmO1lf8DenK7Xyh+U2UO1I8F1SaFtNdUbGCT7DanpnDMg/5N2N7qZWQ7FDkf
lgyqSPZrmiuDNvS7e83sfLds59rND4ErrzbdQ4DFqD43yAwTysUzZ/Emc3cSHZQL
mdmMmExGRetSb64BgXwB916tvwQLRDGiQS7fDAp8xtbj1mou0I+axkKixdCqweqa
A/g7lnBmvPiXCVB6HaxqrCcDVOwSsDzS/9UB6KezE1P+C6kxycOxJAXWBBgAVgVe
6R8fJ2JJEVXB3a9FFSg3PB6rC6xR+euIGuHaAN2ZSU9K0wDXgDll5RZJkqsEtK4b
AGrC61U0JNWS6L0Zz4oU12anPcjyOR2XTIa6rs01oBLpAQ/9dq68/s1V8PpTMWdm
H/zhWsZ7fuAQ3S9rLPvjTGrYlIDc/lAGKragWVq4y9ZhLA+hSXj3evZQ2s+wyWsX
KpFt0gJX9ZpvQl1Z7hRrEjMZISpdW9kn2tqe3yxwBEfLLw+PK7tBL/AHs8RCVam4
pOYAHtwsZSzii26mILOeHDNiKvwVIPcyVrZD3kK3SrHFq8ZAzCqr24tQCLrenZU4
HJzlYzI6exgWWYJD9aJ5Rlt77BMBvmSapsrUdFR8IL3bYRjmKmfw1ixH+zW5aAQl
3WAU3nUcozEP7OF0E609xeV0iWexgBTCAKFtkzzz7F+3DoJSDR+0WTJINb9SeI9f
zKiKoKdXOXgTZzCkmQpAoxUTukv4wtsjKQZvQn56BxQZzzvd0UfSa/7TilAvuocj
Xohe6/OlMYCVtETALA6aJzhaTLArUcCwkFDf8aTH2NDN5O1DJaEjTNpxKO+69Z60
UKoG1uqcPLX4GRGOiSltzmdETX7pNYT5KdPXpgC9dtJ5uI6vO00rl3p8h60jTCXa
tMQa4nvUAuNk+EhkrpP3wuz2JCc48vTSyH++CN5oRIlzklv6XaVb3rBqOcbKvw42
f2zURjgScyZsUYG3Mk2fYRTAIgj9fNea6cCafuKVqYSaQfq9Zrne+kpjTR9Xz0v4
5SOKroIW9e1UUE+90uIVJZ2vx7JJKxiZ3XiNjaDe4a2Q2heZLxzNL//HO8MA7VPr
VKUk4KBTrzer5yWqBvv9yrAD2Jv87V6Pfciugvext+vlduoV3/jTWxoj5drqDQZF
BMbkf3u1z/LOEzWogUWUNQCLbrFB7HmEnPRCRXWGA2jtysvHTYSlkdQaQGq1kSKB
i3xPxiejSQj0TjT4Zf1CIAucwok+tEj+2IPA/2etbFo8TC9K94J7l0EexucgCWpH
ZYeCMQSmSCfC/RmjtK3EJi17gRZVh9O+SXu3JL0ATRoQBKrfq6yX7KlSW2wBBbkP
SHllJpwQdmoylpWe8otdxEcmJ6h9s2FJUZDX+qfgX9eC1EREwJP8BfgoBrjHRTfW
/lYmx3z3AFhtdDooD6/6Y9UgL8Bg29AuMIthLSS0qg2Q25+PteFwMAdyTSC0CkCV
X6rZq3w804K7NupzOkQdKme1LvYu+bKBTslD9lKsrfiW+91GhWPdcwuhKUDtmbCg
r0rNLbFoWhEFOpesvqFThNcVRcRycQlrST5bsE3UcyayyowaWisB0n5LuA8J1mOz
goGmZuaozpjKBbDTGqD2hZrNJB5G4Vu3oGFX1wuEH99eteX+SYTpkC1VVfpyISwa
BIbGiJzYByjSGxRJmAUk5D0ebpfQm/fVEM+SQqGdyElj7dfmDQzr9NvcRl8DO4ya
5NAxbNNil8zmEGxZvLesiuo2aTAc+K/wXVmljSieNDBjtst2hUnFiCW3cu4yLA/n
agHw1EzfkotY/2JXTOdPCbEnR7QTqmdvsL+XS69EJA94O17fceS6da6gGA0tJQjQ
Gh2Bh7ffvCzfa5H1MlP/xdWIo8MeRiv0J5FIHnAQq7BByvETSY55Lm5J46UmCzMG
OVHTw4Cnxbzt7TmF7Huo6tNandbkiTd7XTQ3dgwgJzpeuN6pm9s3lKDx3Dgu0VSd
6zHENwIsEj+ISn227lKbYpUOV7DEkQeTLm4ckrael+F+jlAxfv1STVrA3UjL7Kh8
wrnRXMK23dCDE2JvzHWlZ3S9+SD3XxhXeNNsf0B9FpO4MpOS6/mpH1Hh8WsX0EZO
rRjpJF8jJbyDjhmwCkvgf+WCAzwypyIHVu4ToU3nAfJ6/8wFZxxywxpeO1Txdxv0
tAdYQKRIUaD3ITEsmlIEGtZ13rj1a7DI4tgT/BHIWi0Z3fah8MBOFHLfzg6VVg/E
S2r9+Ji+FQFU0RuG74EDG3oyHstaq4e0B61CzywUj4Y8Hrhy7DuPgoF1AAXDzc4k
JTUbU3SBfHbwW8KevHckCE78ZjzWbju/hRn2TgxE5N0Nrg/MlZP4VJ0zphANcwip
bKKh1gzQt9qFRiZV98KBoH6bMtKW2bvmry8uHmfAeLBQE/0luEdjKUuDnACSJMiZ
vzF3NiBmp2j/yOxNVbCFkHbVAMnDCh+Ts6WpVk4AUyaTXEnwYVe2s3zvmNBAL5O6
W10zt5Q1h97nhhNO+mWzRn/m6cab5gXPuBzorWHvu0h3M3lWjB/cM+71NqMnv2OC
ld6tOAJ3NjGDfmONLrAfI9HBOROg+vC9ncX1+boa91FazSMQWB6mOnZKSl3Rl+a7
18TRn57ECW/EYCpHhN55Ie/7+v2BX+ydIpSz2hA/pn+JNUvvG9Cd4JUj092VapRA
bi4gta8yrzxfS+Op0OQM2LyEmikDMW1ry+9vPkVWzBbGfkAJYE80yDTYo/k7XlOb
OuithVfWkrUJuVPWkrhsZRqb72KYz+d//dqMtcDWxTirRTdzzEAll94N2XpEkonX
aElFWb7yaVpnZfCsVUZHhW+Nl4ZE+BG+3CRwf7S3oYJqrrCufl0SQ5YP7v/uM8Fy
SSRoTOge4XOqcHGmDds0wok4HBti9qah2Ju5kaENfj2x8Z3HmKOvX/TjPYH4j4iO
G3eswU6LTZdcP+GxWIFGUJ+K9YI6nvBh1p6pIaHmvw5F2AuhNxOVusvekE4UGrpR
Op9whg69sfzhslsfcSkX/vyj5YHdu45mjERpOtaEaw0vBzIsVUhaMlan5UIxZhtk
b47FfrGbFS3xzVQ90CB08d51jz/7MxkgA3ypPh4ToO4ZVbKzU7a+Qr0Rq3Ra27pL
KzSyrgX1bkNShHf4I3KyswalJHx8n6/ITV4dGjGBcuVebTu7edRvwJhKsFNeuwQ/
Aqw6Qgm2YxllPnKGQXxGYuCcPh1PRp8tzQs0nqXt/+PAr9Xa2PFjlZ+TLwQmBOef
EOagUip0WDAP3vG5sVnf2fym7GK9J1L0DxdnlJZ/mT6C8a5xbhb23NAHDFR48OkE
vSV6VZ5ehkgx8Oy+KnkvenWLlKILtDZDHo3ThtY3iORGhTKXH7ssfr8StGDd1X7Y
KecVcH/sk0prN1YOQq+5CEq9i7upx4xkEMKqOcER2qLhN+HvOCPL8HkWB3tykzGW
sTgKGzxV+Xir7sp+cUTx2Hy61vlEPbmna2kWoKbbcPxQsJrgfLLdtYMO9xwrEXFM
fwre/Ddw331QF4y5uzjwbKRd7xrlXmJBaVCMqGTASr/gsegm3ByD7XNSCnCzzzbS
G5nx7HPsYy1W+gBJOe4WKpHejyC7NhC73TuuoyWjYn9TEYdX1p2516z888Nm6b1c
nOJzBeYg13yYKOlSFoWc5wn0tIMkNtRQ55tMVRb3UlUte71YwXH/hrgtInt94XXR
KSijJrmwPvgiO1kdrle6jSpVHDUHN2dl9YS2vrsOMeGEGY7BhycWslcKQ2alZWAS
TKcYtzbhjcRuFBd9FFU4nKLUdRbJG0rqV16v/dN2R+ZNkAkWcgxdmKcBkzazqpV8
k+SzPGgpq0vG180jHM11+HvvCV7R+VjvqaL6IfNkEdis64stVzPmQqeM65tFJcnB
zK1VOqVC7vEeRKASbgkl/y5PSFFDKnRcreqXp/M2uEt5tUCRa3mV2XQVA+DJjYq6
O2AWWpslUGjxUDqW4Ec4hndsiJ0bcFexzDGiT0lTFaZE1gu71A8X9XTiEDWAjqxp
YS4mFmsBcmMAovNih9JkAlVN5cau/oqrggqiJmFWgH21Bj2x3FUe5+KZAilzHSuE
q1ykWWWmj5uEceNkotF6WQd+Fnm3QckXDAj34FLGftKIb/bRNNeblGaNqL5neH8t
bho/Bgx4NXGr9rRS6DLoigOJyELte8HjrrurR3D/u4FtjdwVCd/fSR8A7PVsGpS7
8VYNlMWdug9TZyahD9NxNTD1GGwdYRtGKc93+bB6/XhfiRD9yJlvjuK4bbyLVOug
LOdo+gp9N0rqCAaiOPy9c7BRvFT5BFGIshcVuJLs5KohPYols8zW0e4J+GD0dn5u
nFciRkta6BXlGy0dp1l8RG7xQqVTkHvL4+6akk6IiF3eEaDCxeHp2iCv5hIq0C62
I+89VjsfHBdVSa3FdlWDn14qoYenj/ccKjVs8EfGMF4+CPTBFEFl6V4iCuRPlaMr
Smdv2OCnnR6Gi3g+pPMh0DIqxsOPK/xlvljD30ybxbPYqWEAkFN8es/Uu0VD5Tvf
nLvVp2qW+snX8kHI+E+r0VokUqJ0Fmrvgn0c/4uQLh16dpkKO7Sy07yII/VdS9RX
2D80hK/sc9BY36Mmuj5yNWtzBVjHOFHWHVD9b5ZWYHsuAsn4Jzq/QsJpbffmh3bm
Mf+/VNTvZ+Y69lIgNAKN7uW5yKnoTN1MD8aGAgHH8U9tvXEHy6bFZS3CTa0NsPuj
JmnIxTPoB+yrgc01WJaynYt87psVZBUcBRaLdWqdBgzNYMHYNfH0wN/qOg7gyvRH
qWHCNEOhRh5LRCoRMxPFef9U4Jal6svQme3p5KmUckglwS2WtK/xQxRWHZKV6nRz
6tH2B2AfV/HCc9thr6RKUzdFbrwF0Ys1d+gB24gpOxL/31Xmot9KvUDsnq+37i82
LtFFgw7RJDST2fZ15c4bSBdeeevYoQEsnIc8J8QdQlsNrRqpQCrYd4BYNn0ShTUe
gs3xZ5GgPhK0Itqm9X32CWtHo7JqEPAYBQ+mSzyCFBx+dOq6/vJMrv9qdhXFsRQK
7qoRDf8IeJfw+wx1vFuEAZr9vYKSq87WEsncesb8FBcvZVGDvh2tLVnEt0sqn+nZ
xt2NqMNpU3Kv9cJ3Us/Sw4OS5vnBCZi75oeV2C3LFxvD17m8wo2Skg2esmk0NbFt
u4ilxhzMAp3L6x/5bD+Om6sHQ9QrLKHDKBdmXat+1g2ZcGOhT0R3braUeri+WlHV
f9uTP00SsVS89gbC4xX6/RJAG6OPkBYe3NrsAYfT7WmXZLNBUqeeIaUmRB7/QvWt
kO70y20uoj+OOUsh/4Nul7zzNpzg/UoFgEXhyghldHG+XED09Ilzj0OnZkE/EF/9
61+7pgR3zYxLqbZU94l+HWC/6WTqTyIYnwlyuxFry2ZInCYHwoRc0ziBVGwKcmpP
UyEl6QdR4DWNMeuyHEhCbTMTUMQZWuHIHeA8tZGXEUvtRaOL+Gm2L3yKsAwIgzUB
MNWme36FOyf6IXjP6HRENWJ2nLqUvnjBUDlPCTVNhwuCiJuMH8PydviXeMmRnm4r
zKzcLgt5eXvLcZwliIrPTugkErCSOIalwYdUI66ztQFDJ0oTK0/8edpV1wlNi5sU
HpY24DhyLXqu7S9Q1OHuaFtpPVxfEMVXUDN1r1n6MSJ4+HcXlF35bbkohKUoBHZV
5U/Ch6zsjgoUGVU6Ud92rM3zMgUmrwcv1AWOz3tHrw6Qu7SM6TusTs7ub3o6DBCD
oh8NekGzv50q1EEnnOSf8VRc/kycNZ3Ztu63FD7hoLZ6NoM2JanmAgw0LZi9/I6S
aQmvjtzqYHyyGfTLzk/xwIi5lkUNdoCXZ1JMAnyeAEMk85dgWm73OEzwKCD1t9fl
WfDRdUyGkI1iJQOrv72mbJGdBIEVmxZSxfj+jcvB5dpJj0H3WI9bMq9wvsI5bFPq
HucmU0bjT/WKOWXdPbPvPm1PO3IEBnHgN1Hjn7z7evtAV/MnLnQMY5COyDnesc7g
n7Riq9urfQ9j+GqZB5BsPZIDBp/Ap4jgWUHGsn0wfipO8Rohh0UXsDhfYq7XHLe+
yb8Z6M7HOfzN2/x7xiu6EGkrBsfzDFZsdfRIhCxDj7zs1/2NhJUktwnqbcpU6DCn
HFyTGVtfLHdEgy7/SQF1u6ef5exhtnkOXX3iOMxwFQeY5qRix5RUjeRlB3WPzIRy
lLY8kSSwzyBmM06jOhkdFn52MQ5pu+3Lf/qksEGLxQspIeRMCO9R3mPaFMSoC7rn
Q86BptmIz8BBScJsCMulp/cjNVvcj3YeEVKh9yJVrwQY/p3it93J9aum5QBf75Uv
s+tucjULGPN9vHJbhCDG154SSSk1qKy312A98APXR/PHpByFz5hCFur9iUM602T5
SbnN5/RJJ3MwiUBjWV9t1N5d6vwjV8X7FGgnLx1AgSoIGmN/z9s2qPsWZtTuw2x4
hxStxgxyKJ9X61C1IBinvBQdaYw/weqI+Npap1RUspt7y/YDPvWUfGyI0HFjjVfi
5m7QbLDQiZZSsdnmiI8zDG1siXf0ZoiIabzkQdVfCXwnIppMPczRSywMFie90qfa
xCegkugrxc57bBF2jaadKyWXtRbDT/RQtKj7zyF6+Lo6V4+XcG1XfhpghmB6GEjt
jRvsrFwd711e9xOCYJze6ZdIF5NUfLHeU0pHJh4cMnGYSbz3MlKt8rZw5EREz4e6
885LQZoqj65P46djhRzrUc3T/tkQtvHP2mJKw7OqUvs3RCf5ApB7afCfSDu8bWid
8Ndz87nlElmMDVGnM781YUn/49tO1O3zo19ZPj6M+oa+RE6FIYYeo8EwlqMUX/87
fRiZhvI6kYZIUasqAXqmopEfKDM+bC92j5j++19WCfS9B8ZIVDEhEaTCLL6ExlPu
qXHJ9EaFTunLkrp7U/cMovnZUki3yM+Cvt5COnUIwqw0157dBKswHHRYRK9fTIB1
ptWoJ9N5P1LwRRv/X7AcVBtNjEXuKi1kX9gP0QKD/dgAXHtYBYhN4GHvardfdp8R
ZHsSjwEGbc1IgxYH2jFeBnsIXY713n08ZSsltwxu32iQRpePdYBzGMfLEgvEQ8SY
J0xwAjxbNxtQJWlzaz9ihEYhUeGyU8vVcLm5zXvAhTB/UScpvZHLvydZEogm52hS
Q967cO8n0tB7hHWKdb8eqlqludenyA3FVoFyNjizb+oX2352QrzgEXzmf+dhc/MM
+t8egsdQzsu3NZ1koXomuKL716U8boFaPEvIP8HBs4hGykjc5/5crsC4E3RwL3Zv
985ldXNH5B/VArPv/+UpdOZUK+HvsZbtdungoNWgj+rDp5RMpmRE+iThkMI9ijhd
QpKnYd97jub1pf/eLkNoPxleo6pQE61d0/YF38vL/a9NNmtuvIS0Yd5M2BourGgY
G9mA5y3noA7jc+XCJviaYmYy0RD/pts1MmJk3aRX/QR8Sgu8jxwR6Jg+XL8/9Oh2
RC59/b7G5s1qkHhhNmeQK3DgwOPBZ7PVMhE+ZbrVhv4muhaHOt9QwOw8yN3VaBrx
pOZcLdeTjRObAZfmFDTQInqwXg8byeNSnkXTpMcQPkb+S3rEF5887e069Uhymm4Y
sCIeoxLgubk5HhlOwr+KB2g+kSXb502FaetGA7k8ozTVuGAPnaWL9BhHP7pXdYY1
71+DnAdYY/fsP4oinXVLBzv6Jmd3evF+QKUmV+vCZwkW8bVmVA3uqmGyRQQBqcV7
sk3r8+7764tVwDMCMsEXSJ1ug0YH4g7cf9rOxLkboz7OQrDbXM7JnZJKHkGLdO5i
QFvvyOFok3s3H2FW9QP1ZwzIzsrDu1mICOYtoGQq9ufznfNNl18ZVcDu0ae640yo
V5t3Jm8ekr9r4SgEusaYjn4HazpkpNlhTAqiCPFtjq8xLm6sI23X9vAutnOK6KcZ
9ItcmOa6fd/FgBwE9yyXDPHIb66+JPjcfHUrwZ1Srfzt1yrFmee86qn6yKBprbcj
779C9mEdmvdhbGtvdze0XlUmOGFlqTanf+b8owPjejDv9IuEG07drQue7JMccXNR
k+tcuEUm6bmWhr2l9/LFzIN+1Kfqajtvr4KtD1t34ovSmTER/AFqbtFX+QVcncLa
1cP9GA2Vp8DWf9pugOJ/VIgqOWNJO3omOS9jHvDahYRVOWdan50UtBV4Yq3vPMMc
9We5yr1/5P/LntuV58fx+nP1wbpb+3uCH0F65ITmz07pAUHZaIMLnVJCzUbBQBId
JYK+tbFTCWRFDSaO2koOR1qsRska1J+UlhWJnzdmlzeBc57G1K0EEGvQXTaT7uHH
saXqHAaFrCoZfxWmnfXGQ6V8RBIoqsMScKkB7aFMy2oLgBpjOgdR7xElMl/BkFKl
Yu1AAB/WwcvL29/JClNAR8i5OmJHhQ5B6nR/PbODbIoF5cmSs21aFR/ii3ni8Q+I
bkamge7EKELpgOw5tAQhZ3Eqdff59/ZvlabPMs0wYZL+rvrXBEEcEgvRKgrMqlQC
sOZTPQSei1OUJSDVjrXwDVUNvDMY3UcR/8w/ejTK55cdCP0dg1/x1ZGmQglK48Rb
IfSgjh23U7BS1XzOeFAYOWOei7HKmiOgK/7J4J6FcCjL0RJgA8eVuI7tJqx16a6R
/5bhx2L1qUmafkYnIssk0DrhlRPi3dYYD5eIk2GwNyuTOfETKGHjA9a7ifDFcWFd
Z9VOTPj6uowE2+B33cVK5N5GFOmPJj2CDfOxXUtILPgyHvRgj8FhhBfP+7bkEwf5
vuEryilpNFpVjhSEvWmFrWKlspqIaB2NrihTrzP0Ec4A2pW+Vedwl5Lb5lY9OBo3
ZxZsgUTbRGMtDG1vNK1SmWEyCsMepoZD5w7QF3mEM9qO3PB6hR+cJ5FR1dt/03Eb
b/rrLvPzSxQAgQgS08V4MOaa1JH9YTlyPjqyOh6V2mzSVjHHJASjkcqqKMpRd3mL
JC3yqfK2TaGg+nmzryBDn9wiL7pMmpTFAGey+KnojJ/8qfTmjrukei8jg3I9MaGJ
Jtjx8fWIzomrdmfw6wQWQMx9FEIiUvAr+Z14c+xfWD0rULXEYSBOUrviw+dg868w
RC6iWMpHOAFgJA4dM0ITDacwvf0jglqgDs1VoqxOy2it6jDclfN5HrvgqVEu1Cox
MSMNpcI2b2KtpRlDL3N6791mBGuu+EAcI7SVPdwleWvlWiJn2QPDVcq764syKLV7
4ATcF1KLsyZtme2OQcnm/+DRxdBzdBdWesxRC7rAa3mhUKfC12BvBzd+2qqTzWaV
gjNC9zSjbUASpJ18xGpWGupvCxqMaHlVUAbD4L3juoO3pyln11nME01dO7UizcRu
zG1BGkcZUQbgYaMxFYPcuqQxnoST8wty3BDiD1KPk4Wzs5Tdf5Ih9/xBBrOnY40r
68p8xbqBJYwulmn8iAHT48y2I78IqNFGbqZtlkdrJWVmxarmD41VAE5G3eISoepb
umoC7Q57OunkkY8igOjgMh0RlBolG9wOjD4jwb9VJQpEzvQvePAJy+kMvjy/9m9j
K71sfEmGgucyRm7nyArDbX3as1FFC6H3Zet/JvNzR2+ebi3hlf+suoZ4kDpQ1pyA
6oD08rgGBD06v2oa5Abaw+0ncCWrNQmkf3EUFiPEL5rLEdyDoAjF5ymLr1mdYS/q
TPWDQk21q2kiW/k0e3TisddY+1xQvCTgbtRvO4i3dTWDIlztrYrSw6zNeM6QjSzs
1dgYLNK5UxHlsMQFwRNQg5tB5qdRO9Ra15we2a9dnSv/M874koPG+WEr8WAqRc/y
3Ne/y8NfuoFYch7zwW8bDrdgA/+G19ES7c5EHkHysvVTYpb3BSIzNHQDcBIM6YKx
2bYBK18s7cLfve44Wu5xQSD9ghMlVyqjMaqPmLN/r947kNhcXGLz5qsEG63jA122
2EpKZGtv9WtlMpV2sX/+RPaXXd0Y1Ou/bJc/sumq5BikcHWCK649dHUj/Z9NVb+e
NgDZyck6smqqhuWKHDWC9UiX01Oz6fQ7atYh6GTJ8HhOmLNB4jkPiFgFGBty1y0P
0l6i3pYRe0UyULS5ZhMy2zZxXoEan2wByAXnOj8y9FOMxTs/blPv6OVu2/wSXWdF
nHnfE/HQvrsdDt1KSghEAm/yXNsDNKRkku59ld/mZiCaz4VLWZcAHWudyFoTWeB4
vc/3b/pk9Vfe6YtwuzGeO2gbZrdW70LH82Y2GQxRadq3CjOwMVgYYNxK0tCGvqrG
L04/pN8tpCP0ShPgGrlv0pscmi6r4DXDvSoEr3uXFmmHa/cA8jHgMSIeXjvr7Ym3
5YlmTj7bxVojWHP27iO9R93hI2dbseU4fK4cqdhfxc2DLiWQQJdgN7v0ff4+o9Rf
PduNw74+qE/t+xFJtNL2WxseMZNzs8HamCj77xJHyKpYG2vnUMAmfPH+SOS28dZ3
K1kLjbrSmQBKvmhmnjEwK/HOFmdMS1f93Lo1Qi1v0XptcJdB/kbgGqV9pXUy/uAe
BjPfDrLaZygeROtmyPi515kgYQq8oMjEJPQ9Suubt/ervlKXDW59Um5Hbc2Pe3iR
472QozlQMoiwU3TmlQEfxnQ6gFrjHzSW3ffyXcJJRflJtiZA3RamXR1XSIJ7As2T
HeZYsJLulwSIW0T64QHeMer+XAKHzQxe0o6YKTB2TL0tiRhQZ45gqZCGgmRosI1I
Z9AwR8tHz9yxGipA24XQtU93Cln+olpKvNZiV7ayquPv6x4MJHxmTghDqucwsUc5
POdNAbQyoV/WmwoAJxXRwbAE8H2seU8GYVk3cpYWJ+tbMQwXHEcL55DtJz++zGJ8
SSCyMWdd3ShXLEVgot35dycgb6quQXyxcJS0pqeCGD9/uxU4RJv0NW9gfYdjJAu4
QudH+cWEbkGcvlUKkOq3Clxv/mW94g9UbQvao99QwkscPkG/JAHY04FhQYdXx7Np
tdAq0SI0jwL4bBaw7U6J/xacKJs/pHkUEiPeCYnfGa3R9KbjY1Q7zyX6eW+31/3W
BdjcZ0c8oewYEPhlkOK+7asHtlunQBJBAXZ9UBoy02HRMCYWYAuz4RkmlHCA7fHA
2H+liContvdFb1guFLP4pqT+X96Kdy3FZG4udzp6PquJGSGKgtJK4NjNgXIf47SM
apDy5e6gQSrvc6EJlH37iagZIbyOBn7TO9ujARzWwg6O2yTNXxCoMn9SQ1pR9kyW
Stw7K+5YQEd92R9/LWBGESuZZbgP/+gHOoq8LlbxfYL8+p6WK2YPmyyXjffH2BEB
ZHhJOXcjN9Teersr4VIWlSZ0lWBvh+tsZ/qs8x/hNQthQiu9fKzDQRbSAjGD6ehG
NkqhNG0FWa4DVDt+1rS2JmnyU+VsKOIDn/Y9/I8UPWMe5DmWkBR0jet5dg2iFxlH
ZeatVXAXRuBFg9aAizOUWAkIdzQ8q5ydj9nesoZkSlSFCqKXhvRRubY5X2+6++6q
/K7TkFCAXADKBIhQSlDE9lM9i6cSQbFFMU23FWsvYuxuycrJ9J/GBaEfPH6f3tbg
iOD1vkMDjWJPp1trs3niTxpm3WZghSLk21O2WKwra9+8Ua00CH6sh+2T1BBGUs4o
N75um/yVg8ZvqPwSYA6VeIQNY6air6wgBXhjONUEvIJPArlvZsdg3AhW1dpQl4Kc
QmyH88YBoT0RUTXKgGwmwr4Th3sT8shcAW9zRBJduEm0Vb3QZan/IrG8pvd42KKX
4Ln29jGm73S+kPRfRoLVIzuhuAWZz1Jty4yjd4b5AgWR3lJXsBAs2XEkd+c/yHSd
ze0yBFyT9XvMvrmzK/Jj4Y+Ur7+uas8/yfwa2FxynXB4q5XFXALSXjzHw6HPvKkN
omqLDvkuPvF57EpQmu6uOUesXDf05xA6PEg85ZmIKh1fflbxLpcgBVy8kDvOKJ87
4TrHMzr8QcYq8xhXcHtEhJCw/Bo2C0KHAFRraqUAcL5kY7ktHIAumVFIBibNXfdM
zXrC2XtV9v5YKYVe5Hl8bipJZSwJfvi6CeTHw8HEKbvjr/HXnWgKnngWI62KNM+Q
/kMs9gJ1VHj0LyADHExPpyAiAXroNdogsriZ7teJqQWLAWsFYqbBJKcjLl+cx+H6
Ekx0j3YXsgBpG2vdrCfTbWLyzkXErJSMr6ugdk20b0rgLOlTbuAOkHJelyKSeQ0b
+p8WcTmgbeMRT4rBkaLR57XIhmPrUzopwYcoQKJuMOXIY+hqCz/gFpNedwVk6gY2
KmSJntOLfcaFMLuE+x0QMC8VVCpnCILWfzCLIAy6c2YPi1Qw+UNKgx505ViMnKRE
2a/qSPwqMr5gJzJ2YF8oS6EZ2RFEYX02llWlIhq3Y35I6Cxcp+peAOtil5A4n2op
I2ozEStds4ASRRQqBig89oIrr3i9ChI/EB67y6yE4geBamNHn9P/knPaHePIJHs5
iCmZ+Fr6YcNFS1YXk6WSwGrKhh+BqEgXR4J2F1HgFPL6iw3y3WOf0r2NaN4Ao5Ov
MrNBRiUXxAOEGq/A6uG4Bi91cL1gIHOfMSmKrI55XW+rt+mKfgwSLMpWQWJm6fXy
yDUf58GTtHXUNl4nSH4AeEfATL+Y3yd1ms3OQH1GgDJ987w0Zz1DWVGivXXEEGZA
feY2OYdk4W9e74Rc9k7ZDWvcWuMD6wP5JnoDxPLEC0CEYwPXxTQU/Y4HhIh0ewyr
So/VEE2tRKk0kuTTo5CMpWX+YKDfHNNro48oPr+ES5pvR6x+D/+d+fLwZzto+F+s
4CycMvlKW2FStAdWfAQHp0v2rBoUBgfzVRSDI+jAqs6jhrO5QBYbdgWQoCfeWr8X
rVyu7U0XbmibWjoWG0a3iMQ5YREVuE0YFK08zFSvBjDKManmjQIeOpSngbqvliAs
StEsQaenJ1Qio5gEyn/6ugNoPYheDp4GqQD7WPUYfMgBzFRKrM7YfGWfhyIAxxIv
BQg/ZaOkevMmPuNK6M3K26KASqx7baKkqc6lyJdbyCZXHKesd3CD9lZvtqOtzsTR
8uWCd1k14aHmfWooCs+TwFLwu1cwrFqNwRN/b6+xVfcvXuXdkLFrmHS0AvCdM8zE
75pgUaaHAkVKXBte1yZUhf3fYHoccfxyK6xUHz9drtsZFgLjlq7aIgLAodFfCfx6
3kkjNnvvsLg1PAk0Mmr7qOdPcgkiy62Be/yonorAOgXJNLNcPUOaBPwsW3vT+B2d
sF20HBuXwiViPFm9ysCyAXFqUasPVz0UxFH1S4KoI9FzLb21X8xXEy3Ly7jwesRm
e1DioCnOzKF92g/L4FWowJECvqjeG2PlbaRvCyqUJdee4foj2YMrgFv6STTqkc1d
tfuh2jWXmY34mb32ZRFA6pyBiLZ8dHjWoGzDc/FAkmsY+L5cPjDJ8/JVns3H+GWl
eSg9yOWhEe0Ix9cAgghV2u03+xrFEOzhGyZgSQ0rhh8oLVlhFjmfvGmkdSYlzAt8
eU23LLUgni+/oteIAnGiMXTREvgvgvOd+u4vJCB3iOJRZv7hjSkUOYvOlkgc5LMv
6Yuar5oBaouNJ9D92ylwSAhLc1ovBMN05D7rsJUkj+IvCuA+u6AAEzC1Rqj9mSr3
F67DaCLKrUX6m/HQfmlyPuz/EOAYccJsilV+a9IjKOsK53UXbO5K6+GShwtN/uE3
nv1gj9XXPHNgoWPU2CF6uKe+btJo91TL7OCvzM4RY7Zl9TPT+U1ROnNlUsvzCyoh
dzboXPz+TgTlz+rT8s3aPYI6c4BeCKtrPNQ8CaAmi46j8kOGjES20YDiKlOq8QR5
gFEpnvaPGFiC+kqOlLOcj2vilvtg4jnkuyyOdmZR2lZQThhtI7GVpA79lJXTZX0/
4/u3H2fawwIbgpa4aD7HGaA8EP7DCGwgg9BDn4AX96DaMmGapoLQvEiGICydOdMT
R6GE8fEFMdzxXTVnwQ0uIHPdQ+sPEPi7HT+6ujqW1uFM2l41Y/sBQzhXt6nHfEyz
BtPXqYqEJJZyWyPT4bgibtoFqg79OxvQe8ILq1Kb5aONkqozQn5/id1A0/CDgll2
qTI6eh6IsQGum+ABL18Ie3MXGDD+6JsVxPJim5ygraLZMK8KV/plUUIHSgH+L56s
GzaicDtjIrVcphAtHZSNWvubPg+W82MJZVMg9EaPBFWBrLap2QKZ/+0hWsFNL3L1
MigvmivIHQu1kxHKCLuE8Wm3SAYngrfCGGxo7ikaGKQb2u6dFUofPh8h4N/5vI2C
oTYx7IW5fcLUN+VeWyWKE3sHTd6stXcon8PQ+c1ri0aKCtbJm4AYGltcZLl5K9xw
N1Y9fSO9HnoTBX5V3K7ymWYYY/YKAL9wH1+kBnVzdpehYijUivXCTjBjpSZaR4+v
APud3ZKRf/g+MpSHgCI2EqIUNPf9vrDs4uKj+/0iZHm06G2vcOo80vEmnDfhOoTD
yC+Dbe0DX5AVMeI3fTwhKc+YYXgr3OvSIV/UlPVNncIIqfryPWc3NJviBBkLvUne
Ls9qKV3E14kNvriYxt+5gSZtydn1t7xxaYMWC86TuisCZZvnEeKEN5FliX2teT/l
X//xcr5p8vl2h4/w0BrTn00IVSvJ0O7PaIp1koUgrvLEevPXUoY25qHIInhbr3/I
8o/lJnReZoifgg26k3mkMNAInOAnGNOh9N0RC1Mt8FhPJ22EDVkocZfk1Lg81+r9
EfNWglPLx2U8XsNNxnD2V8p8MLlh4EJxvc3N7yjRIabIZqHgDD9HhdXSqqGTIKFz
w8yDmYne6bGKiwtteLkOVMCRsWiTnaAXQ555OLiUHtRVdSnWXhjAJJ/NPKGc3Si/
nGXKZly8W0dxIC8bu14FkBy1hCGCEu/dJfjGJEkDv85qnLYBIGr5i3lnamlDBHJS
jdqDfeegb6tV/ST+ORGIhEMVymX2MOR7gtoBcfpyXKBpWhAY1DWtRBZwie6EHXTT
S6nXGj9IR4SNT62JueIBQXZ3mrllT0gIl4+89HLilAGDu28iQJsnNPOT6jCACfO9
ACVNrC4bcl6oAoaOmBv/D2AvXHCytBN6WC9qma/6EAAAzQwrF3ONrDBlkHM6WxFw
HMRLZe/5BSEGP6MOPLrPw9XMMMW7O2V5pXtML/Qfas4YvazIK0mMxR0TI/mEdUYn
LlmvBpVS94SmSOq0Fk7uBLnJ3KMm1yyyzgsXFvIajtKy6TeQDZVLreXXTZ8aVyFO
nM/rEvLlHgBidBUIkHG/njkDBN7gEsfVUNTCglC+Kd/XKMY50GhQ0wZ+eK6yfND1
rLjXorz9bhyCt1YGWnmK5SXl0hdVxRZgeyMiUrMqjyjlnc499GC1vEIHQcGZVdSQ
R+GQbQTyeI7IRN0gE/xfmlvGHJ89kPJyNCEMG0KaZwfpk3BRMWpJ2lTaYGiHk3/O
p2za/rER2lvPLEvNdb432YhMQcyiaX152Cp/Ss7Nbd1/wCLHBS7FMyb2YDCKwy3c
Ti7aSsZLf70pY7//atgLRnrX5TdJwfcSKPFgB0vBL1c2taeFenuF9yV33Rz1+oyc
vmM+xe7tar5Rq6g1a+MsylT4Yj1gFjYErnpcUdVdVc6E+Ll+blf8OrBRHzX9bzJj
y6EjCe+Z1XXP6wEuHhiGGgrxcCgKmDmC6RVcmezpB7caVlluajPMbnEojNNXTelI
cVeU7GH6DdzbWou4lZBuJY/b625k+pvT/jagis5hXeHWIpYnLgZCT4E+nqE5BuQV
JqOgboG770Vx1fnTEsA1gXqxoCYdIGOKfHljyiJyLEEA9+YBAlz4Oajzyz/f0x0W
SVMUz42F7tLNB5t8denGxphCh/YTvjKRGisRUmwxvxB59WpMUYoCM3ffGXndMBsX
xxJ4+JCBl9QWhMtvXW3mzLTRBCjSwWt3x4Q9+ISY7EH4yUuYfzWqdukvZiSJDif0
yPIZns5kW7+6H2pb0pcnuvh3rhqLkVx1P4Il72FJzHsqr8jwPojllCLH0lzUWChH
do9fk4DWd/iF40TVECO4Q6OPyUsRPVCpruDyCvlMLoPKWNUjZXnwQox2cEYoTBnJ
lQKGIon44uk40Yu5bgBzTL3CZ22OoIBcHRBrSVqPAGoJnUHuq/uJlf0OQkAw0slh
Lo48es6w8g97VwebPeD0I7uc+qw+cg80hPf2M8To5xFcwkArafcQsAIhfHBnpUNn
FnRkoC/N5fhMdaHqY1zQCSvQCfAfCM6KVZDcyrkS15Hxy5YHXJkof6uFdgAHaFrR
/QpVngqRdBjGhPxDDy+GKG9Phpbqdru4Xx0B8piaF0jthzaclOs0wzKAsNW40gFz
bmXEiP2DcEZjk9Rvl/HacLu4TX9t+z+c6mPBIB7gjt0oIltDlfE5tXF7zvy6lv6V
lYou69ISGF2bcYNoIpTxgZI4i86lLN5WLps9Yc3SzR/QsvHvqQ5XNG2r00kjaNR7
qi8K0J0s86sPhBVezmSVXbRfQYKacncS++PwsC21IImSgfaIk6pzydH9uuLUmuzM
A1iiseWb/B4RsWIptTxj/sj8vt3HO+VcRhVxPFm1XpavMrONvjyRso2VlnAlfO23
22Qephv+bfdKZXhfP1Z+w/B8LhI2YzYHovlA//MEkNUzP5BJQ9a0PW3hbHFc+BbF
9XSsb0YBReOCwwmVuyKO2BVVB3D8YCIxxhcD+UJUZCGlq8D1VDFWWQUJXF3RaEg9
zE2ak63nAv9DLK6bpL9rhynsIQQhf3dPN4e5NQc7/NyczjJC9q4hsMpsAB2tRT3Q
DT//CQZXT/6AyFYzOWwMtGytoxPa74PBlryHyphm0uJ9eYPdK8L9BBlHI4cnG7Rw
ePYSrWIx8Khig93GjYBN1dBSUbhwrLaZvlqm6NYtnVbk/GarU4FSbT24TTYc3b8G
unP2bA9IlgvwpreSUuEkzOo7N/jt4svlwI8RkUq0Dxu2sAb+CCigkP/UzFfo2tAW
euXgSP3weWsz5NoLWJ1soRHzQmrgBDMw13Vryt5scFYgcQOlAKVr9DRISy74Q8+6
JKtSQc3eNDp6/v6qIUEeb3C4Kep0TDVkmOUpWzNigUsxKiUPivLaqirifhiV/D5O
ppIagmXBEaCi8F+/lSYWi6PQxXjEZ1kKZTFXYAY73lri9jm6LC+6+Cc3X7olN0a8
FRl/G0TACMsAwUSNMDK2aaYBBo7+J0Je/SdLQI1rg5tMr4Ee+DzWxVy2nXd80K3R
15FQeA9/CuLMYJSwqkL+hB6eNejKt3bBJ04FbAtAarN03eqaBSZfoZXGwZpWEP4z
VqADYDjl2yFWnNOVAFXHi4mPyYUUNO3AwN8v/QrAMvRYN8o9scZVH93mIJphKK8x
vUH7MTkhGydNZ4HHY2AQ2Q3ZOSI5goa8Cmaa9Dr9lYkLX0tPlDjwq/ndoxIc1ezI
4jxgJXi6EBSgnnYGpTwKCZqFptbUWOyh4qEmbmjwd08ZH0pEjGWI6XPj5DRJM1Xk
JAvXwJuZjdwKzCmO4nE8jkvpBLZvr4xTSdzuIDeCuldXczr5rekHBTJZyiBFcbfg
H5l8epoi3PWVdbMV0E93Tor24ZY51ILBP12S/iiiCYaaS6b1R4nHj1wu4Js0X1Pl
TMhqEYql0q46vMWpXp3yxPWyG8sni0uUjGmGOYWYRU9XWwsWPSTQEYAHxMd9ENl9
kuHcLhZl34l/q6ugNOUiJ9dxJKmK7Z8tyqdzQACnPZOjQxA/3wG7gkU7p5zlzrp8
28P0/+Hjd+I9MDpLH1lbVWWeeptqCCZdNYuR5MZHpEhY+T338yhoOlKkKmSBDm5F
IhO2Ymc50hwtWzVpiwoO7MFGycj05Jmz+7cFqeYiXO+HNxQioWUJ2yhMtA6jfVV1
CI1tm2KybaZ0uDZBrxTwiFkHBmuqCfgNxvNCOuKBVHi3uB6wGWNg4KaecvBS1zpG
QdxfPM+4yq/DYfJz/xkBInuCafYA0LvfwIIkUmTwQYZ1pATftT8oPnc9uICcdke9
sERfAIkov+5v4NeQfl46RlaL25FnrWyHXvBmVW+e5eWCDMFotddKD0gtHDcsiA+7
rnWd3+XnIUursi8Xqicd4BJIe1XMI9mru4VPLquvcRNrl8LSXoMuihtAddootrTo
BOJGzysVeEV0nlOMGhotRD53WJHC+FZFRXFFS4px1v4S7jS5YWcQZW0Jkg9s3180
cWhIeI9aHwiePtuXGjQRxZoNMEf+JFZVNdgoolOhOgKCxYziASGpilASEFrbhf2h
xhiX89F/gTPQdS4tLf9OqLAmORTiQLJhi+DJsKWcw7DPvIXMGpXMG37o3Lk1bh0H
sQieGIZmJuGSrFz8mQldmuxq90CqaNgetajmIaOspZCfJHhbrq+2xXczifWm8yDb
T6GQqqRKPiHDNkiSePzgPFborzrh+tWq2wBwbNu2Gm3jA4XIOVyoqIhAg/3KScCC
WiL9IbLlRhb/pf6/NNHDwL9Xd0GDOXlkky41m3yrcYps9GaQ/ZJLV2PfHLNSS12a
sEGmZb/KV2+LmQQQkZZ74/KR6VTmJpLRa+3kOLymFK0Y14+Bxedoawy+lZLLyucV
8NyMvb5UC5al7IQQDNdJlncPikP58oLK+P4a+yb20PLCk1kLVY4rFw1xTqalyO9I
c+nyZfXifRm/hnaVVwnvY6TqmEhQkGhibN5fh0dNCRGhnIZrD/HR8/yBKS42zxWk
paeiuC5rTs6c6qGopX0/PJvr06ljvOhyx63061h4ilo2c5F1CiXZJbyYD//C/2q2
nKWFNW8ypNt23tcHoAKwRfZF8g+rZQDh11fCWfhmhfk4TIIaO9LlZ+ZqMpXlvx1U
GBCr0opr9TceOolSdhWuBZn5EvqepYzLmkcQyf645EFa2+SM/EVNNO5biETCmWBZ
rLZdrCm+iKjo7heQnf+Kv9y9RgtCg9ABoUXGHBD/0LQHKpqQ8MWVp/ivSjKIiPkU
mD5UbTxXg26QOgQgS+2wMwHmUjf7Aqf8NVdmYYKiWWYuaWz9EoOF4N3bv2bIZOob
5jmvjMoqW1uQp/PW3x09WnfA28VYyPHILbsRR4xMhW6RvUXM9t/9rYzvXcwFRpqr
L2T0HjYCnm6lXZmgEfYDkLxs1vbvqP+brSBNrjNsVaf7r+dlUZoR8HKo2FNwT2MQ
KOFgB8M5KgIoq7bZYEFdSMpRbRIH6Va7RBEQIj92fALLeMLRJWQPq2bvAvzQnPeO
ITAeO9H0tKoDgtjKNqAF0pBMHERsPq1pkRTBnc5aTRy4TRuSUr8CjMHLprc3DLly
up5mjzgY6vofTbZ19BZHpCcC4VzbfWeczPF+AwXZtwYm8R+Lr0YHnoH5La2CL85g
4UwMCGOHEJHdzpV8PlK7mC3z9gYZWSaPaKRj3Cz0KFUycHMxg4rapehpi8t/1eVQ
xMm2MFMxmZ9zbdnpqIxzlJu/LiOL86XKokclJCf66G4EhsLmNR/KHMbhD11PBGug
4h+QrweDOKgWp+8xAHKvZOhTSBa9/65qAlWy48seecACqnIEv57nAIjQAYxtQcWZ
eqWGqSQTB1Gy8eXmKYHw17NbRsSBPm4rtnXbGbjZuwLeisC2x8IweKiP3j7pQs7c
K21jyficaeRHrCBB5JEEis+BP9RbpXVUbUQ9K4fFLKtG3ql+WpUUFXrTYLUdNqE4
WpZBqjDo0RNqjl3J6Ew5u0z5bu+7y2GFQFVnl908ny5kME8rjtrufMS44Z7s/PEI
YyZynYjMrdKmVOpylKpnqSzcyQ1PRm6rWVfCiNYtTH/tP+RKcactICVMecBp50tZ
EAVKJD5mYzqYVERnW0A1Drm0YEUZdHxrBGNPDRg75BBIZmrvkyBaRsnq8Nc3ATb0
5Wdzzu/qpOKolAFHkgkQjFcpuUbsE32QE+Wm2og/XnYJL4TvNFxc0SnH05ixQGoh
Kf17RRtEm1BbC/4ZbBBZkfscIGTQopHDoPe/Zj9b7ry2cbn+S/7Ac9HPVcBbDCWc
FQxBPkZ/SQZAPvrjNAUIzS20uk1dkulp0tSlIMEU60PxMpQqOErbpYFMIySFgU8s
oMeKo/zIbYLP2GZBLiBvYvXtEB2UIM1+HiTYAQdpP2r2xWXhE4r1HraHVI9qIIYv
fANJ8wLBU00HMLU6TknDdFHabNs2miKJIIA/m+WlLkrBmQKX9Gqk5WZ7XohXP1m5
wakl9KgdzB6DBVdfB+z+pG7ZeBOK3q2mGOuCUUznKftSlPN8NezVgch605F1UJGd
yt2nHGrwroIOSMnLvTcO4ds8IkcRCtGUP5qeiptpACXNzZ1WncRTtiOyBDjSI4t8
PO1ICVOu5xvAQkAzNPS3L0Vu27oCgS/hcnZI8W+/iyX/gga2KiOvaiPDBrkjLW1a
gFov6iLrqWobm5gd8gQjh+PL/8w4FNbND8PWw1KwsM47z0dwB6aBNhC+WtPzzLZd
7l6XfT+T3JITnRflcVuycI1xBOBUra677x3gClG5V5rw1hDJ1Fd0UWY83CjQqZZ4
dsWDv8m6RTDDAGwA78psnVjxZTMO9/zk3AAHXeha18nqezfj0dBILQ14J27pAQIu
tI/3SsY14gS4zb9aup+EoY9jWBKSTzmEQY87N51S7XoVdFHzFwNgXz342ONQGgPX
q/PBw6g9QZQnTxzDRXa6dHRTkiCruKKaoZ+NZtUF4incalbOI24PTq6PlL1PwGQl
A/7W2GKN5YjKlsKIGYfK1E/Kup1erAml7MpygaFvFlxczAaRmQGppJhuiosaRv3Y
jAgW0XdRCYE6lcOpOWQco3OZ8Jk1TDtq79mRLFscdTm3Q+5/t73KlQ673yC3gk5l
dDTyh6R8N+9ht+xqWxxVjuKqSVfN6m89bYEd84plrfV8lZl86BFgwiiyd8H9PjqN
Bw/CLg19MQjId8r7Ct9TFRFP5tUq9Kah74lsX8nEUmj8QeEqrHAyYztXeaD2HGir
ZFJz6mMj7obnC3vnA2bxFnUG7hwPaI9kIjfAR1QrfslEjd1iuFeh4fY2GgrYtt1O
ZjnUPlS7oBFTl6r1pwTpXAm9H2/8O4B/jqGqcfsWhZw/dUkjR1ZF5h5UsfgnFvc5
Uh5tnVt5jb1Uo3gVD2LVRxrXmtTcBCbC+wfEd8RxHRykaABToMTQrxpmGXnfUFPS
5o6J6fG/taxZuu9tOUC8ozGrC6WDvOAWcNWaKUtGQgKkfWGsGPQJu1ocg/iBOqzO
FPsFJBV//gYmwD3RuatdGxz79VtG50L7lyjFnP3mfvIhfA592bpUf7EJVddX/BJS
6nNJytg+i6eN1/GoOoi4qZVh+pHKORZWDpJ/bpkY39KOjp4chywLEhoUEArOtid0
X9A7ri4TSYbFKxS8fi8am1cT1Z9WBbjb5yb1FmHyCEbc2v4GPYsu4+1GtFKlUei9
cB/KgzQcxHLxl3bnKdsqB0PxB3Ht6dBjoYQUCq3vo4ZpmdsJEQ4YgekYXoqhhlhE
fk53IJMmg3XM2A4XOzN1nKldG6+XEHFvle5wrriOyCgyHP6G745kF+oIsUXeeeaf
w3U5hpCXN0wTsTk+9EU+Ab/UBuotYpEWtsAcOtV4pqzrQv75UX8WxZjuDDhOzI9r
L0FZLeOOtkv+46F+48h8dCbyUu650DEnTR7uK+0y/m2dfjmmKRy96kc5AVtQpULQ
i2pBqdTVi3avEZCHVeM0qB6+0HqxP4rAge/rFXPcnbD8fJnY5XaEAfbgu8KwYXDa
8hOLYNqH9gqMUhsljtI5sGRGPVeOK+ri4uxX/K1edPn1Na+VzCqVFTISxt+J16r2
AUV93NIr75puERB5H0zko+xi16KiFzrM5z+EFviCkmA6JtQ6TJR+qe/Zn1aAmNyR
Xm9k5NJc9cTZyICfxq+o4I0X2LMil9wkjnwvkkklvm9g9F/aDkFgVSksKhYTd33p
6C7tmD4mTyK2eyjPsMtrB62GTJzscrM+erueuGPp1Y/PuF33at5gPl5Uff0BJ0xZ
mYZfzb+J7JRk7Ader4Ir5f5SJXV0S8bDrey34E8Xhvpf3Dt4aqVkRaYrdIs/orPa
R+MAZh8TYncJ6+kXqxCIZzctP6BdJkacaKaubp/99FThelmvOjrIgD1tN0wzT7ey
d7sv8Dvg+awK6K7qK2rFBq5V7cEwiKBS9AVqt3JpM/20K+hPiNYPGFL+usxUVzul
Z+skCidXJvY5Lw6BrsuILH4a62E8BgUGAM25B0/vO2+YfzBe/vprVcjPpy50Cnw7
HzTe8OPBpRwRFesUmS2bc1JSEnMXhr326ppY7xJIya1L2TVL8XTcbaUIsnPopBU3
IRpEKJp4NDVC3r/1k1PEwRSLsCM32zIScnX20K46iFcH0YW0gO/oN+UL6qBjEIcq
tMOxinyDn+A0RD1qoOQvGA+VMcZ43mDqYQomefYRR8FjvrqqKnmrsk07oC1NTN/3
9MCWhP7yL7LiWq23kMbHLlr/UFkpslTyW58LaNBUgnECsxZOhhSUpdYGVY2O+842
GXjm12VtIabhsmvyM7Yvn1kSZwvt+w3nv/HbA+218EVXpvkOApJO9Pgb7Soxj0YD
umEQd/QXusNruG/gPhknXUwQuWxnO7oe5rNX6o+Udn+iBvzGMItS7yV0GJIDZyCK
aVx0OX8Z6uP/sdbMz9r/taTaHNQg8TsAEwqJgDvD/elchJkpzvruS6xQOnd5zSPc
GuRLBWAk454m6XOCGeV6mFkDLXSYii3iyKpPnmrFTZSe54mX/sT9rl8wuwNdYtiV
kbqpUFYtjLB/Vr4tMdbF1qLulYMmofZeI8pECeX/8vxk9R49jiwAxxHNBBIQYoNO
b+DsmOJSewMq2t+6Wotb2zuVz9yWG9wQ/+HSovdkRg0gUx0Vzh0xs4bxpJDL2v99
KrxjwzeUPdczYcDJkjG3Z1gYwivjunYivL8F42deF/mQeZmi3irau4jvNMd+07T8
VlQARBXHIqDhRB9p243eHXvqCb6GMCahfkJ8ct+ciyU+sQoUp1zxGQcjfEhPU8Fe
u2s5ja4XfQEr8wRGiumbeAlNXkysmmFln6soy320+Ygtl6xoLAYnJ98VcY/g7tFu
IB3/cajTp+tQSftGxvbKSmR6I9jphKi5a6CKcg9JH1pczzvlAbNlBJ42vPHLosUA
K3T7cNOXUzn/roLimg6ujsWFEcTHczj+uCEIkWb14/naXfSbiB5OeE0AMzYuyw1O
yaorTWxqpcsnLSbOiUk0Z28EfZdhhWyRQSr/4B1libp/EnHV4Zif9QdJEKEXvs8k
EiNqyM0cZxfx2YocJ1VKjhiwb4boUKMGh7ZAsyQEbLpFqzcaqISAFFwsGxllP6bP
cb7b/kuYx9TeEsUqF+TeY3y14Vedcl7OYSIFF0LW8khr+GtZSrMXJdqLq7TiExN8
lCTK3gvAlvKQWQho9iNdiIDw87C4c87AluGULcoOxaCY0ow0+N3fJzRraKHaVq6h
rxtVrzOeVivh4t8jJ7DrF561fvtxlbAT9SUnPjt8prbAu+IclHKgTr52WDhCA0ng
PumKI358SfwMxywU7bRWm0q4ox+Ly5GfK6ngevwsCOepuSwr4uEAxj1rNJB+cGEc
8XTg4ZM4eVpIzwApF7BVY9N+nqHuLUJD463Yd3H534ZgJwAKCw4UWjEDERHtT++J
9i3lEIqaQ5wThRI6rkhCXFy0IvWOU2F6k/w3Nlt1XstPsKIUwbnvIDRz+So/pLSp
f/ehcpULpXvMtquI9MvWvWaAqz5hJ3iPTOZ914XxOhHSM0su83+LWBcY4l1l9jaX
bK/SheFWggFAY3TtHo1YkzN2XQgyYa4x+31EKf9F/joYz27nuMfJpqFIvwQclXj0
AoIJMFqdLwIPrdYL+Mum7Jn4OClD5cxCFu71h5lVHvqmeXrsw+cuHupJf3E/82nC
pOUIl88quSIHMgaI7C9uH9VJamlP6qLA+rrgSyjEcH/hGhsKZ6nizPO6lIfG0dfl
FzRjKlX8NAnX7fmb5bA7WnlA8IH8YMVbZabdnV2eeFWj2zvmy64XJVt9zwu3C938
8Z1QBVhKMn3lFbPr86LvzgGE4+zqWmuXHj3hOLXHU7bMyvD3wZ5RpbSajllQ/K0m
P9iCthfR6Q0+qQGPF8/ijHTz9Wefyfpt3rZwqK5l9IcjjpQcRAxrvihyWDo+NGXl
4eIl3MI0rgnX4mM4LUgkwNxDn5FsW/8hg1kg4rFxWBquOlaqXFNtZXoM07flgveO
6T1akn81ZC607323RTGz2WRwv039wZcJEHfEXHBSwqfb3qoN4eI6w+EdAolrN/Am
bSRMLcCYVDzjpG8onu5CfiQvvVUtn0lZZwKAG7STbvGPP+Qsf21WRPJZBwqKqNwf
p+vvSo9Agf/6KedZ/RztPCC8U0GoYpyGosp2BAzc2UXkzmlt9f6jaVLQPNfxoX3X
HoKe1OFxiDxwY2MybNCvA06aa7ZykRmsxpiKelErz4aScFUmK20uUrxFzi4Mmhc/
WdTsC6m8HiMxh1s0SvRAC0r7H2o7g44fblHCvRAJGIoM+aotfuUGQ8YXEqDuvDnf
b9xakmzNCiWv5eZZh79f9okJ9EhtcRbo++ngK3gtB8wFeFNwBIQtG2jwdCZA8Ocn
B7VT76ujf84NA41VwABj1/OX8BVh4luNuyXBd47KbBA8iojnVjRi/nwdPQ5VQPhx
LopAeHodpCErB6PZGROfrNMuBqP9ZyZfXzQWYRQK08ZfyVElp/ob7UJNuEkJ7+ha
+rgjv4j/ekPIhOLthS0Ure482WV3WTNG0jRxjgL1WuTo7wMhE2aMBih6Y1dWVij8
eu36FNrJ3qHYnf5lcfb9zTZMAnK/YtY21ndPOckjcN/xL6/Mau78Esc4+W8jD9zX
RyIGOMu2hCBfDFwwfB08YYSTI/KptTa/74du4LsRk5gPFebPutNvsszaQUIdNbyd
r2W0YhSJcMITdcaNjtq0P2aSK2gGfPBtbEDGwt55ncqZkxA6NApXiOROXZ7siABr
ySOIdGAlVb23iq8fBZNF5L1witJ2ldimx9AboN1S5ss41kSE3j9vXQy50CkZKV4x
eVTnnq1YRzFxqwecPmvGEvZAqAvwvCAW2VqVBuzE3MjQDzJxg2EW72Myy0ZIGqc5
VaMWDEYz2sysrTwXTuysSqXwOL+vpfsVEEJUGJk6qAqmEQS53EoBsRg4O9CCv1L/
psSsTvV4bRnmj0vFCy7zSGEhms4mNFo8NpYGrZwKW1F29zuhz3KJzBqJ/qxMxUeA
sfCeCgN/9jcYr7/8o8MvcJOhGPy/N8Wj+0iTNP2WhVJNks3/NgO5jKGEuvC0WWTT
m6NpUbnVmhOEre94ZmPM+wQSFnpyUOzp4jYRgwVuBK5zX6FrTax7/JF9qDiJKw0K
aNWQCi2T9A5oMqZ/jADJ6jByrYTMnutu1N8zeidy1uLFoks4onomC6zUDv1n/NY6
645jpt0qh2u+HI405a9ypvKuPwlecg+AxlsQs8W++OJdDBklgFN5JcZP/21JpoQp
QsPxumHiUTAsNjzniBI4g4SBzpOc3Y9ZPDWzDar97COOPv6i++zhxrpWsyFa43pc
WJqthhIxYA8JrdapULw0nQvWxa67LZPzTkbWask7BT0luta0xLwgfjeZZ3hM2Lzb
s0D2zi12kn+cHLJjAqxYIsDryMae7cpaybfW1uC5pazG/EQ4Jg0JSYE7Rt/w/5nE
uiojASAE+sR27Bx0eRhKjhvVVdYtCk4Q8Zf+A1wXO2cHcn7QHFmIWB8zW288F4Q4
dhxxkTH9jhaXt0YoArtymV5AWQ7uIK5QTPVmMQcRHNoLaTLtQaFlfdQDCv5OnLPf
SvgrsiaFDlIO/dDONbtGcZWmePsm/0nSXfOzwCl8ZtJvUeAAI3oDXsdJRtQ0kgI8
Qa8yei4zfiUdBkj9cQLSev0fMz+QmMrZNX2/SOv6ca/eeq85wqVNhc9tmlzewaKx
jBgfYzo3TR/pN1h0NtqUfhUfS3wK85ZjDFDDJaG8vnPVH2WB10HHBFrsAgZhXelM
yog0I112If7XNdBiohEjqHUVJ2Io/PP4KyUNFCLjNx5EZzSiiL+LUjLfcCQQVbjG
hi+aWEOrJP0MZoOd38MqWSB+xez88BQpCss1d1wSzqce8dhhMN9oEQnJ4g0kJF7S
r6RW1WQEj3JpAbvGmi/rWHxZ/ZH75/qTJml6yQhzY2dTs/NIOptVHwmqLI1MIMiq
YxwAoqkBeprEfViZoPAUiRtWifHW5OPGngZf7JgrnFuRE7x0CNjjNQDR6M8DyeRe
u+pdHDNOSzBhM8TkYHsvlUXSY/iTKa5P2nEuAIynJFIVfbyfme1EPGh5kkeoNKb8
XcD1H4VTdtlDyQ7LJgSCHlrd7o5ByZm0f37cGLUnhNLfQ+hcRAI02V2mMZojnxuj
vk8rpAlyZuT5peiTMmMbc4s6CFgSlWh6VlUVmw23vf43YKfxE6QGsIPbPySN7n6M
hPMQyidpaJTLiqjF0w+na8UuFDMkDLBKQ1WN+ZlqxGiwuobNvPJUSmLtBP6pLCzh
9gr6A9rzx4Cc8oeGk1PcW8UdpLdtFv5Nod7YgdfUpeJ7ECO9Rty5zSdyBo9i8GpQ
a2P1y9wArE2ws8oYZfhUjOBBhhNFN+SnME9qmeDu5yXbyAlbw2Sp6cuFOZrxi/Tz
JArh8ErQE8yCPflUrDdpLTvVgUFQYmuuL6PyChM1JAr3MjeA+1xQv1QIbXZUv6lw
1jIiDC5aYKzQRYafLxkvWRWiyjhZJmTFylhjl892ORLlDYENbtINj1H4gKqgZ1AG
ZkoQBubsM+EWlQP6+XeOpH9WTAM8910tG/ayHirGKV555F01pCG+tk26MjCfK8SK
oXlbtEYOPH6OTfe/qryZSU8HQC7lNf3nHTaeZ2hhfREO4ONAp8P/98k4nUO4F4nF
FCEQw7AB1cl6MzB73V83dPMBS5Sxl9tMPyB7p8canTAenPzbIUr7dUPXcRoPVDHH
y3Dh4nqk/diLpWyB5Fxu7tsJHrshBWO2qOMrfcH6dI3ZQTfw49DSt+Q+Dwq20Muz
Fm8xdncc+iDjfQzDUIIsDZxwlzkHwDLa/KVQHp1kx0kHVG8x005zxsZq7DyqWVrT
TAKTb/pnKWRIKXOGB2DODPWmfADKBQN8LEKpiY6lIy9GihgYThOfhvogBkFRlEKI
9T7OqseRBa1LwtQ9myg3zjU6QqLBzlt+bwSpzlZgV//qqW47VJbixRx/VLHyRhWq
1wsMKAEjhl2SPqPi2UKQy7afJF7fIP1KR6kNEfOhwCYtSsPjX+IJG1hSiuOR6mL2
Gd5XGNtyq2SrD4CLO28jQBINpM0JjRqe/WfbzZI0VU3DiRfRAi1BgVamIXMiI/np
SU6cA9LJ5Uwmftyyuk71rH7K7V4x+2Pf9o4AScwhcMzHXqXzBFSOpSTf0LfuKHjI
ExDwIMDJSnE2DZ3STcwb67ast581nDDOeCngsSK0Ph3FzbFOs7iz08SwrBJnYk3/
wtBKAjf93V7U5GrczOGgRGveryr9ilsQpJiAaQY3CM0dVEojebg5gQERVEmRUZgS
h9yF9R76lXeG9xrAVdj6c1FLE9HOfMoRnr2LDA4QoG5Env3FNVa8DKUCTuGQFVSQ
jvzcrvrDF9DYY0Baf6VAQd6ne3W9aMx9MAIquA9GQqg2/j7iIekfHyziDYyRuPoX
uLF+m6ThsX8Gx4io9h4uAkQNtWG/VsXitw76PJX7HITvV1Pi+iuQnx4/EbAgMED3
vz65RpfOEr9Uw2k8AKazyPsDOEozYI35hKnBXHm++UhUlEyw0shyxj3usfZ7hPD9
eJdc5L4xkCxEKmBfN/Z9ZILB2E3TiFWYGBOIr8xpbl5zhudSFnoifhKbOLRWktxk
uVBsMPfrRemRrhOy6ucrOHnhE5+ZCkKpt77AYuwqA7fhdzasntuq9ivUYjrKnPAz
jO68M4h8fO7zXQ3bqLKCkoS2g3eO27yDMwpXk3l+xDb6aLanlGkJW69XUgesKI6b
1wWwZzhIrCINQ9XjEb9D8MzF2qk/55Xo17JoyhjXnsHCycKhaHnoJ+S4kOtPxym1
SutjJ3c+EofLc6oH573TU5izoLR7S9Ig/EOSWNfSjZQZh+YFYhsPRflDSJvd22ME
3IbrZJL8UIacRPPenSdMUgPn1tZLe9Jy1tspL2PpeqtnLVNOilNzGRrNIR2G8Atq
Imvnk6VkST/39uLIoAzXdCA7BytNjqtCBTaXujH6RURCtPJUZCYsUpqgOBdd1VjK
CgDQ34Z9GMP8AeKwSkgoCM5FBEwo5Iw+bxSpKkMYDTugR6QHgyag8NMV/uGU+mcZ
7l8mJf9T2oFVKuFkuIczFEeYzC4uQCMvwMr02UM09Xnl5SXXOqerHw9tVZOCYLrc
n+AMdfo+YmOYbnC8mYzIexGOlJvSPvShb0O6etrn6PzzbqMWyDC3D7lafTkItxUN
NPE5tCGTIvTf5rFL4hrOmWTm2h2e6fu7pw3XJQcVMlwDvvo+JbgbNa8nkhzgPJ4U
KVnrlU9gNULJCc9EawRrP64wBR8DW2Gu+WrDOwUi882giUWkzELiLRYgrduLZHar
6CW6wtYYbUQp8JalglqUNJ9+o511jMUsV4O1K5JiFl0VpJ2yuuNDtqr/XEsC98lw
R0gs7Y05Uh0YMNLVVxRu9rFh9qgGKF7eMxESGkBLQhi+RaVZ76Zzk3/9YK6tQDx1
h3rZA2cAooNKf+KiZz+U5NHIz/XyiUHE3vpG2Y3xBfF5U3wOBUBJpboADF3Ke1pX
KqHm0zlTcwT7JZ4y72P8qQWi6uA5H21vAdherlRpEIkHQdecTl7lgPMmknYX4i02
pzUmYqozivYEblDSJdudeEgDobQvk7ucBXyQi4WFpe7Sw7mG76tb1hFOPnaxgLKv
k+GACiluFklrdSYfSJEH3+p3FOLha2vxEL6ro0deszxDqShWBWlXuoALhz/OeSPB
rUbz6S46b9zmO2d3d+vtMSls7Au4rxasZ7CtE979NjFpJgcjfMoynQxWm8+wbfBP
9h09Bd0PQT0SzqZOwzmn+Em9LgJQpt+t23X16rdCHP199hTwWIInrwEkLsdRlE2H
UYZKOarNmKtUD8RunZjrxAqnN4h4AN+yfctId8gRzfp2S+6guIjLi/8i2XYksDj9
Mw1exJQvI1Dnw/YAZOJCdYMA7wfX0a0xwVfvCbDVTILau8/ehhPEcQZB7ahxslOr
86xYUaDTh2pZY8wdmoHhrNXQ43y1SyN/npYGcGvtc/CnZPPiBv2ElFEJ/TUQwHSI
aUVGBniVuAFXQ9bMxSGZVL7jAC8DS0rzxzzOQl8oiURBxLVpa5ZwXpT2Ez1yWoLr
Dwe97rWciboWqOuX+wT1SSR1nbsxPeBbape9rA8Ob9H6YJ7g5eYZe8NiOyFEftaH
14sI/DePan4KY1Vvoe3OrR09/J5AjMWYO6vzo9SAEt0GMo9+WSDROvmDSl662V10
MSOWqnuDUODRuNtlmBUFeVMjHCsIBrGewXdoEHvV+pRS0VoMcpzyayVSX2KsSLYa
BBjqpdj31ubJOmRroYzBlChJHXfIyc0OGXna+ZKh4ZoYxkpbitfVhKsL++YB5Pwh
sL/Mgu2jR5uWvipVXUUXG7ZpqUR0x1VQb76xqtnsck4GwwdlOKd+UHPvFy+L7ycu
dBRSqFR/gKSDWmHTPCbbnYMkFuQ0kbmmebYUgWcOZyghQzgpdeBf3zUetOV3iKVs
uauBCx1A9fzvvlVCJA8vviuH1X1//EYWg8gwrLFlrUO3pfnvMqOwfSds1NpX1VU6
Z6R2ZRaSJBeKF8D+0pGnDE+cUyMdzU4tZmcdAIR01kT9c56SpGBHO3h2aTPL6GMB
Xx5+LNDIxXkR4mOagVxw93tuzzB1gyFYu9O23resBZpuCY/DMPXDM2keurOyZPVa
rqGI2CLg53ZObk/YwKlXmOFypjypPrcAvrOUUACMPbQF7CCwN0xrH5loJavLclZU
VFfWFvUgrtcSLlPhRe2xbwigMu+j014FCmnNujBh7htVzqeE00+YLP7fJwlEF5oU
XywgH/xU9TaK7WJFMfqGU5whcTtObslutJOPQfczsXT7AFS9HSmypqq20ntl4cQZ
to6xcz+cDRR/3vNiZmxhenpg/690GilAvetoEC+FSM+bNDgUPLqkosFHNQX2z8G7
kXa9x9RR3qJpGYF/e/pKsqQqgQv4g4yG0z8S2e94E2pUmERPS9t9gzGxqPiKLLT9
Oy+7eblKYl3UHF9nIakFPJNaUAholLk8pTTOvzzJSQQWXm95dZ3a+Z0SfYEaycW0
yk2hYeBdcLmf6gYwwoa1N4APodaZHur1xvHU2VLF5OJ4v710BWt82GVxy+3DxtYa
mFjC4tQyqHplQNtdyayn4F2Dkv0yIfEspnErbPPS8Doa+D4xCLKr3ImqhZ+dSMSY
RyEy7lHkow2CLkVbmbX8QZfsmtcg6iPw1J/7R0L81sk0j2cO2lX8Tf9ZAw5Xiws4
dhqtfkUiaFI8Kb+kjDeFNQm4omPNcFv+wgM9Z6ZY2sBi373d5L4EUvJbknqG9Nrm
1T9apPHy7ppztxkkzPN4tT07ckTmNT75dggPUKNde4tnT+tNtMNvXoS8qVnXt4ct
fyyBnfWvpyY+7aaa6nTn4f/mBx0xw5I/AWxjSzZax8/AGM6UnUXDmTl53quu9DSV
qb7S3gUlTfayke6sLVMb0n2gZYipnaACDB5/GKVAdqvwcKtrOUMEbqumgEy0zoNU
BvHPd+jB9F8ZQeQOAu7MyjElSANd0+yFmwctmTV3LSJHza4Xu7pjsMzAlE9hai4P
mc2YazrxmkM6iIt278vSOGuodaLf97Y9s6F7vIzS+I1PmRf6OjnsBqavU+7zG2kn
WH3XE/k/KHq5vr1pxRAm7UjJW04f48pkHTwdl/Nr7i9XIOhxa4ngt7Hhp0scHwfS
DpmT7C9edq141KAeUOXypW++bzmkPnGVkLLHpxsySLREyvaKAqFBHYdKjki2jxOW
od74D7jx2EJ7xEOzHtRns/jr41Hw8OhKhQ8tBeKZFD/OoEeXivuWLu1un9NY9p6U
VOqe2ZGTjD0wAf2lxoIe5ChK1rYKcQrm4tbg5KQ0AHTFpD3TbnJ7U6lRutoihx5U
z2hUvzJvjtVXr7R3HTO3NAybFRzAwS9US33Yi889jiJ6EOGoUVeN12BinDvHVem4
uQ5+kRuyiV9ndeGnDZabB2GLcPZpwSs7YEjoHIiAjaGw+mku9derBITpZMLFiEhW
+E9L6yuCMcqr8YIPAnVDvqhYdRfwac/wwY1XkHYZhfUN8G6T/QVu1gsAF5+AhAfR
b5dl+Buohnae4ah1sE3ZjlkWXvNekEI6Xh67Lc0G8Pm2AldhL7JNtU79qtjfmBwh
s7KpL4/xJbxZvlaeGCF+lp/lc81lVuLIGqEXzPTryrJynl5nG7CavEvu8cJfoOIe
aG+aSKKzUKt7JA2JuBDOa9zlXTBvIS/ExRTzSOsVps7LTzWW/rlk8utgIYjtEr9x
p9HG+dJWvthldKQQxQyA4ZkZPEal0fxnmHjo7+N/X9rLMIZzSIVTkkh698lB+z8e
C10A/mDcB4xtVxwUrUPj2++RIJVvdofr3YvaSqvCnW6MF71aO7PBXdOXXuXYgjkt
fSuICmN8HdCxJq2N4wONGeZPHVAQema+RaD1u541n3EFBLpizXM1JFX6y/J3yCST
/79u/HdS7r6l6yvgCqzvu8GTZDl3/i+oHqeoyzQ7Xa1MsvUYrwEcOqbP2PJP+6oK
sN4SeHpfhPb2noMoUgNYjmLQ/1/gXi6XrT3dhwfJC9X4oh8UpQZSr/arNsteDCHq
GqcyQRb3vLjZ9QUm1Y9oGKhgPWEdXnJlJVrLOX9WSw/R+ErKEbDNtg9e6DXvTenK
SzcfWUkR28eJqRFpmDGA9VT4Znxd52zKZRyd4rrop5MShsRCrBbVUhy9iz5mASPQ
9vu48va9hBXKhg3u2Vo2elNBfctexPAypAfL6VZZVlGv5d233Q+QcoDcTvgD2qji
qYJ7zgY+5StcN6cV8MptuXb0TVe/35uR6SyHCl1U+BASOhf6lBB4SYIDFLLZW1Zl
frnjPwNIgCHwtVGDSkJXvVCoO+4rUuOsPzo0u8uxDrTQ0RKwcx5txdwkn8nxt19s
zZXuUbLpnj1bZhsTuMixPisWnheAL6tjKfFK1/2pIGatG/fyIQwE95V67ioQ9C1P
OCzetdUGGUzs8v08x+tWMbxyoS1GcfD8iNSDiqrd/HyREbF3rCct47Bhn98h7/8q
FKUEXx1dYPsNQVEivzy4Hlm0j5NVvG6f42cW3hv+PVuJF22YA8dls1l6Anv0uF5o
BjoJ2HUljbu8LZvHI2nilK8fLIyqOg/hW6P8xjJDHnqdH6bc7tvvxa5d/2cYiWKc
QC9vcvdMfumB1+lICwZ8Nl/ZJLOANOcWl7Fj1xt1J9CiWAe8unUFTo+qjhq0LwQE
BZUAOt5g445NT5cPbXCu7IjoNsXu0znQshI/wh+y6rwr+Xndqtv0OOPSce3I52d7
MadPj5E8vYoO0V80IE5WsZ69A2BfUytptpjMqYSI8Yf1R/YCufWs0+bitRh5xIgw
JlJKIJ3Vh86027/xosL3AXuXwGosvx7jmhXgEv6GvgnIrSE3r8u9jdchAt75vVGl
y6LNow+ac3CKWFrKFA46aOjIFNtNY9db8XfXYdcVLwt7ghxuotORzWyuXtuUV4cn
IKv9I+QaRt0MPlDdopuAD9te+MsAHfVrNTchNDqjEdY/8qcL52K/gfuUnc5igVtq
/NCwLWdl1Of7FWscJC+l0kKL1hJ2c26NKhmQOnBfSTJ8R/HdjA3UwZkP/YKWR8EZ
dzpsezErvtwCZa/6bQcWDmegYsCy/WGfp887+hbd9dt4EQEhND43Wi4gDhTB6Emz
VHNAJXrU9UEKQeRgEMUb1gnWaPpkQQHhl9oKZG0st/IK3MZrMhKSb/V+GJrh5AFe
UJJA1sduO1MctG47qForwF1QIubuD5wpDWVOyLBtaIqo9PhHY+VZPuVN0Sc5W6ZM
0kiQ7rJSDor0VuO3BgJr70IzCJW558faW96vyrvKzaWOwAMEvYgOlX01o9lOnnXL
u+0+t8jwOg+0v02ceSsuGrTp4/++N1UqGy7/DiB8FlHIOTsJft6prYNcVVWSWpKM
ljfooQ8pmWQDzNNfLvb+5wkAQ9srPmyBCZFPANwkw/giidk2dcPjLUAUQJiJfFeI
Oxg0mC0A4ICW2z2+HhapxLcv+85n+ZHmw31I52/MlgxS8gJnp8bMEHhzgDRsQWTz
l4coYjKODwoErlIDnlB/HJHLw85skYd+vk+EWyecwGzi+XqKjdYH8wM6LpDKJ0U4
DyXQUG3Wi20ITLsTNVHfahBeGrdnAQCmBWGjNesKHXhblZXpBT47doy5VEWtYXwT
4tye+Ts15qUq1tNNO9UWR3gfD8F7HCEcwgnuS0UcXq45GiiW0V5dsnTfzl03kerW
wILq5/QvnMIRslsM5S9PE37F2NQuUXJ+E9TXVijNTeTdQ2EaabBTiYYOzlnUVEwi
XiFVlytwsDTU3V2n2T2R3rL/FISfPUdo37Glana0F9Fg8PY6SQ0A5omdRfxekDO5
Rn4i7aWCnzAicWEuewdIbTer5yjlKCSMWqAsi1kxSb+yO9/aBHweG8iHMba8cmg6
LYl9fVC5LK/00uKFgwTwGK/SWYkR4YjXuDmNQ5b5EceXjLE0eqLDwhiKOQmvq0vG
p4GxK0FVWI9zFmAlLFXWP+0QRC7Gm5peL9gCDkYjn/XXDcHQ4PcmNiGzOilKeZJF
zu3Ay6I7bsmm3QjN0Qe1c7ZKFbPqV2+n3sAiy2pIeDFgWspqK1kAWUP9iaqA2E+e
7KwC/5YkzEbz29VGQXMqXwkKV0x/A1Bry+g+GJFoZluDkr4lRqRnP8/bF40hXlMz
+OGuzonna/nlkVPkNTbjuyJ2uWGdkfF1omI/P8bPKKWkQzVy5fOQnJuOE0uW40Tk
1qPyMfFxgpR5iQ+uHM0v6Km+w1mXY8l8lHBPx0Grmj0wDF4XizuLYY0OYYi1t7Ct
xMDxFDgbxeSQnTiWZQyW+i3PM3aYJe2kgSXOg1Tmt/8kpeqf9cdWpUVD2shBvDJA
gNBMNHUSQamRFSa6zj0vGQC141xTkewLbp/cHt+Qgn4fJbV3JwHVMxBIPMwAywDm
UmzWPXxTG48MBhWFDl5f3ImZiLeFTT1cXiGBkgfpKFCLoMMjU4usuMfivisvrF29
+7LmwVPU3rd7UEqLVxJ7pGOw+L8+C39Q+5ruvwxEM1HDND3lczVTseHRzs0M1iyx
zxzinsO/jOMmVER645pcYksQjPS0xotDm2d1BCbAvPwc/V/B2JKm73fWDO//enlw
6fedpI/oEqKabbbtiCnCf+2pBDwlsCYzKyCM4W7a/RUX0inZbAEOF0Z8TfQ7+/Dx
SzG3PMTXsXB5sN6eDZ815PQuxnxhOO/lGJEEDwf4SK4e3d7OFaS/ubMqEcVGe99v
vuylTq9e72He5YOEdgkFlYtONFTegimGmJk5G30JTAeXJmTPIF2dX/8F8eQBpFb/
4TeqKCqTeKuK1W6fCwECkaRSHsEOm9DqDyWrGaoQUhOb06U4zi5G6yQTDJg0Oaz+
GN6o7oZznDXmaXWaWltc9qdp8gr25ejdWmFvE5LteqPyfm73fSEpmOf/x/ib120f
hWAOFAWySWPSvlq3mMr8PtK0OMAMtNURusWFgps3a0lj0CElKoHCt/oFGC+LBOgs
IjDNTwyZStQJ/xH1XdAsJ4/AWODtZ+HZSgEPWzcZcs+rtam0LMJJKlaiBQZAhDmn
VGbv8zeHfO0xHIEyuJv3nLh5177V5jePxB3iE31EhQcOiidwKGBrTZe72QghsQmm
MG7TezRSK0331A8U3M/JI8G1OZDllGoBnGj8+QIHYLRgx3Hw+Imuo5ffm7A8YmMR
QQnf9z5dvVF+6dq7O57WEE5RwZPmHK5o/MWI+9r12OzUgtK3fasyZAtq2HP8my7f
8Do09wyYeKn0OWJ1+YEoU+e2IqaP3/0OO+xJb2q5D3s56r4hNvgl8Oq6k6WKnUNc
zPMenoxixD8x3CB64AlU5zBSU4nDpbLiEXrccgllU8iYJnxVENvxfH1hd7Ro0iw4
zMiVki9eN0Te27L9DA507vozt6GDnegymVxcP54gEZMPjpCCKcwYyS2yNv7Umked
uU6X9MxSVhwGoc+uq5ktRkzrx7td8OwEXizkhwOAyEn75818OM2Rj4cAOxVr1/uR
muknXpK3dvx5t/zxPtMufXtsF5pF4OeWtrEdzm5fQ/voEn9epYp5Zp3ddIpCFOdx
StjmoOPJ1vnagrqyvHqB3lZ+bQ6vsx++lJOSF8omFgGznIA3/Agx499ouUFGkhOR
OjFGVRBUHmCcYPtFqsTuiafr2vMda3+0tVWXc3iKLzOQsbYyPXIBYNlIK6xy2hs8
SzpZJ+vfr2D9raV4Xe/tmXqKxrRfViC10WvLwzGv277PuI0oirJOB6qIC4kV6CRy
atxVK4tAUue+Pb+gJfOMal8tYpAJBZ++1DEUdeqZS01Hwll8wG1GT1F1x07aa96U
tKawvak7tNso/ZjxTyzBU0l44yz7hLI6ed4SQk1KFE61p0/ZSPThrZ6sBQUd9hh/
oatMcGbX/sBdQMj/DYqEmdzOlX7QPOPmUKoDUrvlC0hxOUBeps6SjIIAVvudcfUo
ttaVYqzeHqlv7z5kW4Xc6BHkO+P2OnQnUiEhW9EIjpHai56arxlpnjm/J1BDjyz+
AbhuMwLiUqw5fJ+H0ysr1jMTLJDe4ZvyrYtJOnKu/0noR4QgvywXKknxmztzX8BZ
q2YI3DcvOL7vm/WlqO1nDKddtrYA98iiIZTgmh8olu1bVY9wCv08Xurf5PddjXBh
kkPKWYC6/0plXYPIb1bwMNgW3NEcHdX6xHnh1nZfVVHMiqGxCs7BL+8vYW5oWvYv
JtjYGKV3AqVrsXlHcaEN72eOlRQSt0qKq9ySovYxidQXTGPZLWzSvTfJXTTmfSjJ
d9Jk4ajsK3Wh7FID75/h+ou9dgrkzQORT+STyOQewHRBZN44xbuYV8nbZDBSlqUe
tfDMp001Wq7SJwvNkmGeB6Vl7asmT6eCWrzOH5duhDAItKCRaT8XQxjUJV0RIj7/
lMSFqFxfZIY6puJWmxVd/TmObsYbNzK2ZTsg8y+EHymxNPP71Xbu2qSm/v1YkTBO
M1+rgu+/xWzrbR+yCfjJlidQZsVrsPqFEpEwpyV708li6O3XH/0clqGP0IdQyVrq
SJ5KSgcsFni4qA384ldFHkwE4Zvf+qgqqA8fQBDKRk914ktwFnT1dNcLIq+/9D64
qVuKMFc3Px0Gja61N0rmvQM341vutqWuKQhBjfxp4pUAFF9oGZHObxrI/2AumrEJ
DXw5zxFuRi/7Tr+0Ln17dH+qzWyTaI95obXCzzRkdNp1VN0jub+PodWPFcle0qy+
/iwRBdgnOJYPzQ6PE7zH3hja2uGJDljqvDZClogo5RIOqVgJJZWK89XBQpnLQ57L
wV7ANsm7qtH9KzXoyH9WhL9mwdxYBOuDYx8qaT3dLxsIeJoDyOYHO1D6M5sO6k8g
hiSf4KUi+QOUa7+gOM5CtLWmQE7Sm/0hiIfg5Y0wAzepPkxU255Hjjz02ULXf1Gf
CKiIdTrMFlSb5b8yCW2MvUQlQa2VndQOYnrjuHZaH8L70c6U/90SnfVrIq+EFtTF
l8PYAJhwvuc+Ujpir9skQ2KNP8jhoBkWEqaTuZbbG3rCsryf6+37hkQzQAbnLa66
+wE5R4oMegUVzEpuOcKz8Gezx13hxIk+xwCSX2jBWbZp4kWOlpVcS8p5TftNpBTf
eNRnt4WKOWbz/eiHWrQfbQkd28KOHcDmd/D3HCEnLH7RCFnz8J0WsUZnUx/Reg96
9QOiU/jeLs/Un8NYwZKPrmQHeXu8lJaBQzM5oSFzoNC9UOa5+TeFXdqSmTeDXWLD
vh6cKk+uDlse7mKHh5T8scSlrnsebzc4KcdWl238GixpOaYJnCVyqTI6m4pQWZ8T
rorffOaNoUyR/ommMRR/KF58c88teLX7VIG3VTJ3f4iceZ3ewTPEvgry8SHYSFzq
OPH84BUZxoTG+EqTMHij+8Z6iDWnr8o9Or3KPFbq6e17vKT9sE4hTyOz0xnmj9cz
87+5qcXKhesyTW/XkgiV1C1W2kGZgqJpvSMJaoMc4W507XCKhJ/S/L6u7NmLAhwC
SBK4jXVlLXM9BKDmFO9VbiN0YGm1BJD9GmyqbbUKOENjudNmNYLlMU4NG63d4y4E
yYw6mwem3oi/1XTEyWJZBfon8/bgCKr4hhTkP4Qv1rxZq4vjmxD5u2RNKKPqavIM
pzJe8ikMKAjU9XZ+vAadhQx2qitiuaE5SJA2qMiN0T4Lkup+pGcYzX9uf2liU2R7
yR/IErCFehARZvnobkRBjxvl6OPUAXLnIX/2fvfqWmA7CUxS6YHj+vrO3RQ9i3A/
8jPprUq5T85CahqDzfV5rY7l8mvDabYe4u4i+8lXS+lgcTZV7FckYu5p+hXfMAYx
1YF7Qf29/INoXvQY/YhenAaxisEYRQIRd8B+v4Wwr0wjuCNENNub8LIX+bBUrwxR
IJPtdnDtlubxATkUYrFYXeNIa6T8LkNMRCtc1kC90v7D9YYYWdoeg6h/rDPO0w/D
d0i7SdSbnjfvTbhqRFPbjj8/Pfqu7vG9k/L8SnTWpZLRfWzznh5Qoz4fZSsraVDI
RXRT+lspJj0rk8fwkaYT+8vMY/j8Xe7yTOQ5TqOhHJAM1Lv4K7/Pw/NaTg5+7iIi
vYYkbRXrztT+FQ0tPgJ4ajrdyfm0oQo5zbzm9Vp/JzE6MaVtS5n72UYeI/2v3+8j
fQ/yO/LEv9yt5I2eDVjAG4QwHiPaSZSYlTceuWFo3YZ8tTHx/SHaGqqtbQYP+WbJ
IZHh9Hyev2e6+UZgmEGW5M+1E67IByy22IXPNnlXySz1JeMmBEfLhCW8H7X7yNpq
1S5WmBlMUIDOhPEiXMMsmm26CChLDZ5EcFciMOcGX9/k2FBViXaxVafPCW4Z+zv5
ptjHREV2CHpCTHRzWjUWRY/xsji6xNztj0EAdgbswYUA5p/0uSX4b7FcODloiiK1
dP/AaTZeTdjNSrEFwhVY0Di96QYqc5aH6K+V+KcV9Dp71N49SOrSDeZD15/ePtHO
T4ONJmRtWNISKFjrFNSM7MI6FE32rmuEyG2ykaC56YNvccqCr1vnBtBtIBlo6rZy
fOqy1bXZTaRx4XtQh5xJRyUrjpaUPp1N68gcPzqOkwbfJS/4MzlPSUAl1ux7vCD3
igwI5EBIWCd1oaPK/CzAbgr00XYNeRiuCxXWYaaVQWQbdi67stzXY41lAU+zyukr
c1uOz/Csx7GQKcuHrwvJNv6xFiNeh6dBlVAYmnJ4OYGeKpPSgD9IMkPKheRi84m/
iIvjXRib6TpfPFj69yPHR2+ZrXYpCl8l8uGrVpH0yBFdeWAk/dUySPodj9KOyv3L
gPZweKRctxdvabX3eHX5UUIG2jknoF0C3b/9wrpwFX2pfr2olaZfC0Kda43DULTS
BqrLbv4oZEhshd6qHuugJ+MyUDNlbSrc6WrHUGQmVFcVLpTajSh4xUPZITKDSiqQ
vWifOyYmi18X1O59+0+2TNhxC9vga9FDVxsiZOrC06MwsckGMd96EA3/vMyk4ODv
WN95h8l0iG2s6DezGoE7VZ8OB33q4Kg7N3K6Gjbk45u2CsCdeRddbgk6BxaAwZfZ
QZRvrRP4cJee4/Ph7J3chgw7/73Dq7n01de/RXwM1tUSEMX+ov3881l3H/bmkOAO
5bZVu9ZjkYB1pGhr9pwenXAecGUNS0XuRpNFbu7X/Aeg9f7mJqYKuE4EHP5LrR97
xocXkaf91kpJSbS/I4JkP+IzTtDA7MnB8a+47uHI3yoW3anyPyvcX6XoA5q4pxLB
h+PFP4uZ8j3ywBuZ2Kps5bTNME4b3uQNJzNBVtGCRqKj1DqVr7GM+g+A3NpR82h8
1hXojZ4lXD6BPsGFV7NaM+GqYnfrX2NhjiGz38kErelwqaXn/zQvXofrAqYdJpW9
is79miq4dJJWnTxMoT61N07bGK7W7AKEE/ezUD8f+xjtkvNmhIMMGQMX2WKrs735
bY3vkIyChSBhzvwTRYeZoqLXE8+5sLlSt8hpQ2JTP1D22J3Mx6GiD4ir1Hafg/cs
CBdpvNreARGlFpQEqQjG7iMXGsz/6Eyqidbi7i8H95s/smU6quvqvbK7ONRZC/QF
YAGUSpJHJCP+1Ndj8rE6XkTD8hPVh/rvJknBdVwG3WWQrnlHcH5BVaM3Q/K5KN1B
0FW/MWR94gJD3ihCkoXwJ3xVh+qUQmAGUoql1e0q4dlHxLbT5XRCeSzmdzB9ojm+
EjJVM5Krm3SnG3eCwU2hWz+NFvO7nLPH809q3tl0BpNU2OCkB6CfRtTmgieXxlce
3RxQbM/oXeifCTQWWKeWxCGyN5+kIWomR0wqMKQ5kWqZIKXTyzZq8/AtFXEBHmhz
y32WZ+BYtFm7jty9kosyE4Bwgd25eHNlVYrTg/lKQydpoBvUQpjjTCIeM5fmZboQ
cmwjFLxUSh2GS6by9zA33uy1Rhlb3AUD7gzw/uUVODZETFOcHzwjfY2L1cJzofmz
JieE8ZCgLLnfy8qScwQ9wLKlx4zP2LuHcAOgMsWnrJT/ptfJsfvbZc1G03i9L2qj
ZXSVEwZkvAT/NNO/vkWdzZ+8n1MwLR735klQ5RWJtt8RxZfH7eTTpMNHGVFqoyKn
oZohO30VjlJ5xCKwBw/ELc1LdsARy4wi/bGwwVYxFkfwPxLFMmFXIV8aRQvHyPQp
0ubYDRUg+qvHg6jAtGk0bhHM/52zIh86tKy49/3AQ2C/7y2d/YsNFWcJQFq+BtS6
U3q8jG7bsMsy592g/lhvEzh0TCVGB0INsqGyd/uK9fA9gvyn08zXq4r+FDEU0J0J
gjAjKTBAntNwgG/9fUPYPib9Y7+ZdJ+9qM5599JWYKtliHXKJXDzTMgWw5qadlSC
qMT1TRVd9t676SMoIfnaNYNKPoTLZNG5KcE6Xdfx5TxVtbjqTLje1WFVOIUESGYg
7ESQWP7wocKp9SpZ6Zkw3W0Z3k0qq1ZlRj2u4mwN34MjT9r3U/xUp0ZxDBCFFsmv
SOwAMofcWXRW0ctF7xX7Zl59x0suiLUUs5/8hAMIPms3IEz/jP771YD3l5g97WiP
rALdk3OIlnElxRNbjp98U3fXDEWmnosom/IMiXac4MuaoTmlCgPc8rRfwXCFIKyE
31KcYNGXMqZDr5aRTCO4AquD0iKfoX5OjI3aMu+a3CzHd6BzEc/IJEOTO6eGyCHD
f1/9eOFvqRWNE5yoaa+xbyhejy5KAsDhVud7TL10ItVownfhlro7DK7SIoG0xHdl
h7T+cdZVesQ3+XerQnfZUx9SW1SFq/TL89c/Do7wPPanF/Y+VvxRBOWw09o6CJ/8
VM8OBx3w1MZQQdo4Ar5sAdtxaPwpiDOQJgNYkVNesnw+GZXXpRbBzJR6LzkTPGyp
Efgf39u9rJCIcd1CqIFF1+dWDrQrHqyUw/ZHidlISQr2m6ESMmlhLcvZtnhQqbQg
OTBmPMIYXNCcfKvigUvu1Edqb06ptINkquBdvxoGV0fOfbDzTnhduTlFHJJtTACS
K4hDkQu/Ny+GO0SA4ScPk25KV1fKNWnNrKRQ9VFyz/8/L6oYtfUzoM9K5aeJUHOX
F9idMXy3aTNwYX/DViHOEqEHNOaq9Gtn3IOUWYhtD3SI1H+Wj3OFgfdQjep/iNv/
cLESQIzaMvuEeBxfyn9Zr4HoZ0dqtJvue3Oeg5ILKuG/oqBco3GypRI9yRT7IEKj
EXayWB8qBIN6TrEGBaEloslFjOp7OyRqbm6wkvALBnifqpw2IuZbmSh2MPw/TeOv
FWgnsj5okn3AthzK5uwh4j8uIezaFpiopqOiPIEEjGIwKIMJtxx9WT+d+EcfJMPP
hmD5rA5bjVmVWWed5Yko+Zi1k5HBw/zYJTq49Mvtr3Sj13zZo6vPVHFKY/+J5RGS
1Yn6JdHjH7wmKvFnSdXwONc8a8vPxfYio1+JrJ//8YrQrJl1X8qmwLMHHiuqU49O
RDm+I4KA26fudWIew49NnXwiTo0Z2NxEkH2GaMOSxDcV7HuikDroxfddVOEQbE1M
QkwbWjP/rpIfG00oTywW6YkmmH6nHiLQJohY7NM4Lq6xNpQ6UXyTvvmLNqUqSxwL
uhlqLp340kr7mwNOyJn16De5JJW5GVgZVgqNj6ElauoJgLdoBUmnFFCkF3fkL78j
CL3fsYOKax6V3J7qnVar0n1G7mvpCzGplvclr6+XYVYkA/xV6UcZmCuyTIOFkPYP
gn8MtaULoV4JkZfr7IOzRuvQGWX4lstdTvhl+ru2Xxukrz5DGNYwTao32im82Rg7
RujQEJQfFBRvZi2w2duso3ay+ECXAXhd4ByS5FOyR0/mlgImLNszgF15umyBNWyP
D42OTNqwapx/IjrgCYLulUyG4Fq/ydOBuBGM4ksudeYJqazxOx2sv0Zi7yTlheQK
POws8FavwtfoIvlAnWqOsO8a8fkH90fQVQywdxFtBWpXXOUbEXtlvw5oNakVbFud
F0yrkEPXaukI1eeaZdwt8hP7vBJvaMoJE9BkGUIBi26OswPkeoagzcUIC0XcJ9m+
x93FK3ACyXj47H6ZPJ1NoG7jigV/UWrClYaHizLZCFl/6eEDIvuOkbiRbA/Xdg/8
aLbObehLjEnQAWruqWABMpDQnsnhQxIyd5069S/SVN8hF6KVcJtruXiVUE2HzD8z
wafxteIb2diBtOHECIgHa7OuQKiJ4V6Zpac/8yrD8txA7+NnMr3jSezrwX1ctYao
4QUJGf5eyZfRdxGBc/rHUr3IPRJnYJ4nOGTNLUuevPP7URgRdcPtUKB90JSdnZvB
pMhguiO14icM6At91z+YpeF8xa0QKLxLc/Vrpr6XAPPuYaZXXggsUQiTv81ORjBC
yOj5zpghDi47ItP23Vf0ZzlHOaSaTaewmzVp4q5gxfPwfbEk1c7vrcZMCF3j+bWI
OLsSUdU/aqUD+nDfT2ET9gF59fWAd77HbG6Am6hgopKDWn8u4F8/da5hoZ7YnOyx
W45Ix6L6QEQ7VLYnppM2aSvE8g4caL3E9IBit4jTpk8u6fy8eHn6JcEcGnR5539X
W8bG1zt4OydSWLczUotdTScGIZ3zMaqCrNBUe6gM/SBscUmqWpvPofT5EySs0pzL
+8wr1ySZv/G0PqcuwmAx5RK9/zzNoQU7kZqE3wnkPl/Fq0QsuebwfYC7Aum4VHms
5ZLyizkUNydq1tVkaFfkVbQVzSRUrWzrBQTjoeozdUasTpeoA3XedOcr34lAf5+d
aXo4f9G/JKyaAHTYDHTIvGbdI5XGsoKCINyL4RiNsOLWI49nHP6O96HMBb3gwFii
9USUr7I111DUuuW6qZtO+KuA7jPEzxFatF5/Qgz4rVG5bg6udJh+GVza0pEBvjM6
+awkngIsSrxRIYKU9ByVtKlVCHMIZ68B6ZtvZwfGSATvhoZCstcS751xwEn8NEWe
0PDzeyGZ/xAguVoWk9im/AKtTAzjLqohAyIFh4lnd2ZIDN/Dx2TV01/GsYv0QNkj
eeiHgy15vAqhjkDb2lF8dlJjRDLjLDad629PfQrcL4FQdpP3RrVipd6Hc/m2HYNA
gCYEdX/RmoGlGktuCZmN0FcLjIkgc5U88hg1TgkPP/PZjj8iNG1UzFY/nYgMDVym
bkCIjpUFKe1GLOy5XmBBv7xJmVb2Bp6qe/T7tEXDMQ5MZ3Pm2R/7P+sVNy7wntyy
ResumKd3xhGp811ZnAolap5zZCB0HsWBLma5SgXL0qIGYK+k1AmqRuhOZ6Afs+Ql
gAZnkr0FebKTb9zjC89CRnn7AJO26MZwcbJviJr+5dCd4CiTMfSSay2IE279DBvK
XGAEB8lnu2apFEc2nrfRlHsP2a8PUmqDFFO8cNbkCyYyDgWUGWTbUUG5Z/eMVExe
/NsaiD/+AEtC49CyBKS8Mp9tFgqkeNZsM0YMEMDhDHHvBmAIWt7unrydq8HgbchT
iNUaxh/hbHsOaNKzMkfJKVbMA5QzQNJ2N1a3mk/FW1CtocpbeYnGeeK8cy0dwhma
SBM+vpGiYKVb6AF8W4wOuYrhf5IELUnvdcKONUd23kL31UxesGtq3b3ib46I7Gyn
Zu3s8HcGE5Rd1iMn1XEIXWSPZnyB9Hj8wu2nXPLvndFCWcikwjfOYbqmE9ffWtGi
Oql0HrAJdzJM0dAbi6E9gU/npPq2VC+81eYsegWr9/S36L9ES18R8rBu4wJp1HNz
i164wlfCd5SlxWHzWcSeuAEKfyCUMUqlnj1tRdDZur/S7M1YvJ86TKIzD+4d/ydl
n/IDSbuqcnQqU7d4oQLZ4Sfs87DNR7e8AWcsCI2S7XklUuy4jDs1wOaVgRoeSbzL
5oHe8BukVEV3oE3hNBZWlsT2UW2RRe5s10XdCi96/W2kDwZbzyMrYokVr1Apbw9O
RtP9ymoTjsHmDMUQXcLP59WV8zqoMJslty31rctEKHhEF9lRgIMXrV0DUFkMMmxw
HvofbZ5Fss65L4zVo86Z4DNv1URmEK+roV28d8HMzskb6nmKRARGhPH8v4qtJinY
t3UJ8Ydu+1cooDgi3CLg85rRyZiTRh8S3kLz57/OrxG3nqEXSXevzyORtaTgDTBA
ci0d0eg1mfQgHhjn7jiHS4LiQqlMHp18XlSgjiJVVhCwF+ohvY/5c5K3TVgMc8lb
84Im5rtWC+1IdDMaC3RxhU9rQZAX+EN5gHuAj9dTD/vyxe8d88KsziOBkqNJiYrv
GbOVzR/1E97ExirQOY8T8E4QThLXJAUs23pjtv3gxdVK2YSUFsiG9/M9YfRcbUqv
Clpwt5ilXKsCHoPK6YywQyecUO3mB6YryJJOmMP/LwACmRRXykegK5ugrexqA0FT
bXhTbvB7pkMH97a22K3k+fIj7ZLmPAwdFmWmXXZ/fmdkZuPsoJI0nU8qAM+GrAJT
89CsMgJwv+R9zZ39gZIwLkZ2G0FLq/HUwtvJE968OlVr8h+/SKL+wdqNhVXL2eXB
6D5IrMzm6nZy/eSnQx2Ktg4ONvbax6pwTRGz5m+lM+kdJArwWUuBFVc+Yv8ZkGwL
jVFUqwYYwOOk0v4C0xMYzHEmI2d0F/K0sL27p932azMtMAZlN+4uKNL8fZwI94WV
l6zbjbNaYFmHUy3uVIJb8J38GfgLmhPk7pjizJy9NKFvQkWEfiQ9Nk/X7nULxUu4
AjgHNNufnnI4wQosxHuE8TEBsUIrYiSCLh1SOKbLHDMgxyuRL4ooKb8sWrvFKhq8
Fi8tlcK96CipQQN9nQVl3d4fKu3suJNWE+fBlXvUV+4v1jxAUmfPxrbPwY0qs640
+6JfQqnkPIRzybbvvNTkHRGDsaao+In4RV60F1v2qhM6aVk1D+XkDVkndoeiKj5b
RRW6cGiEOHDzceTdxgVTCx80yJWpFi4qY75lupUvehtBXgbd2aaTDi5T80c0RrLO
s22pfRn+AG+ISghIEUGNWodbRwv/9yuiHQu8W+r6Z9cGaaXJQq/AVjTyxr++dLmN
jmh1kiWGNUt+Y2IQZJztm+c1Tv4vC2QD961Qn7vPw9dd+tXcixvEMagQ3Ryq6tYK
P1flSiSQ/lWnCKRpVSmmFetfDqtu81mj2TLl5iQpVq47T2RXmE+0jWIaq7N5t/GH
CbZNiHI5JPFAZvxTxEaK6Z21qDA1rIrpCjaIACDIz20BadlHiLc0SkRAy+KDykGg
l1j/5Pr6TPe8Rtvm9IN4sWgF3j285r+7t5dIfF4MmoZufsE2kaj6xyk1mU8dw7kg
5B5lV2v7bl6fxm2+NPKlyhYhr70C1TNd+YVk7K/E16p8kYfE/5Wkzu+C8cX+1Uns
AQxSQ/eTtfUY/gGN6Tg25hXMTfnhmTzI13pctnIgBW7k9KNHLVm4EzaOZfFBvw3G
VJP5piWOQbtQMioCmm5HPtrjbPedTRUb4HdRp5PdWo223EHAbNPPfbGjS6558KFi
yqbDidDe67IGnEIPZBjyek9GxBjGzmSZ5uIAy3a0krHBVpztvmAvfGG7CsSrb60n
wgOYXjIcyF+fScTxtedqV2/InG/sG9dkoLjbTHTYLGjbJglzFzoen8WRmGN06dfo
ZeP9kZNxJA9AH4o/J+p4amx0r8XguLqGTlBwtJ6GKKmprksSZYjEkA+CA5fkpIoz
Yy/IH5/NMqtpwxbjIK7TAHF7RTOw613KIozyvgtBMEsujE5UmYoH8MyPw6qBc/e9
Jt5epH5u4iKrCoT0KFEFS/5gf0WvDfAfM5DkJWbjbR7MpYFECj+moamRtFPc4Y1/
5YZ2vjutW0nVrKojfe4CEYw5JcGHj2+UrINubT7psF1EwyhDDZg1HyTif3OOpfUX
kL8q7LRhQ0V05c3gQuwqbmJZG5SEUbSjCwPseus3RCgqek+urJqUizAAMnQycmst
xTrGK9xRmy0/R7SxquHRrwjbMl6T2ecaV0pO3HPNH2mWl+VBTdMuNZfUw5FAuwD2
WsJ06td+WlGod1ByK3TW27TuPNxMbHtGJ/bNKHkj+k8F1ByvVTxl52aQBbQP26ov
d0LxTeSCACrqgLg2rdpPgn7KG5uZ13wCGUITawOjbZHbFisTKbsOYsrh9xqT+HqZ
0R1V/pviGNIqI4r/e22XI5qDgSrGnGmm3Og7JgDdLhlNlbGktt/EbH6lgpGL3U2r
MPybzkK+vy1tsdTefjXurUIoSIa+uZoMEf0McFMOZhy9A5dR1LVW23AJdxpj/alB
eG873TaYUyFJs9A7gCc9bAdTLmNbVZmd2NdqidLZQihWlx18As74ukfdzWU7MRhP
WxpO2u+Q5m0WfonJnfLkJGlk+WmbedR4tcvwzy8bdGxLblk/LijUarL2a9qPeac0
O4LlJ718YQP5EiA0WKlq6g2gGAvJ26b3S9dAgA1yfkXRcO9tHwLEwSbKEO4MS1xm
N5FWSBzayNAMzDe+cAQEGbw7KjzfXDo6+fcudtzBQInU7HY8Cm/Xb7s0yvd4Zqmt
VWtT6a0IZW82nwnRcuyoCDVtNKjxB7FJw6RKMUQOmZWnIg/U2AbJdMHGSQpbS0ZZ
DPZ0SOxM2mng5Q+Z53RS6gJWs0FNuL6w+hjbU5zBrV86WOH6b00/DUePahIt2Ri2
3E3RaLGqxx1j4xrvM8V3O9cEhWYAxR1ZgCH+6HttlD5myjhDVnHNRG5vhYbC9gPK
jyRs6SNG03qvSCSqxZTJamWScvanW2l/co8aC/QUvn43ogcb/sfPH3/yC6SmIp3C
EZrZT89tuOgpeY3XsbVJu8MZEhdFt0UwShcaV9Qn8XrJ0lu/+D2CKrTyIc/lsNUM
jDC0Hh4HslKWmmC8EYy9kZ6oK4OwKvsTF/SbdplIJbpXUtFwhU8nH0aSMqXiy2JE
jAGIlzg+LvBgnCPZRXGKwW5n3Ykri8liKEEw64HyIL+7wRE/nAQ7a0vZQ8s7BQg/
ceko+RlR0q0tKt4F2nquZ5NSiltgDzCXtm60HY1gZVLpm2az7WI5OXWWNdpcTgwv
FzHSCyBHwQ5RAxD+mOun4fM1uIU4W4sJIHxD+lC4i+OEMwGszneBIa7cFXPwi6RI
/E7INPaqnSZumWmKucr4JWsW6NHMPnOpNwwkYmSsMxZ0I2RcHWpsl3+rHO8/JH/y
KiJx7yzhatP6kUWDWvxvoB9Aqnpl67pGwHuKD1XzmoSO4lbkW2g5IMoXsfKigNN6
NWhpeK2Othp+JTka5EiamvZRARTEGdrCXK8ERLdquM11ESDDFneHSHcrJGN/30AN
9dUqge+gcwRhLKQ8B3kGG1EB2ojMr/a3rQFouR+ZBYy64KkyXvBjAV0LN5/HEUSL
g7f4NzjemhKVqiHkt8R53dE/eC+AbS/1k8AoKqCd6uL0+Mh4ZDBZ+5zvrTiFj9E3
1xx3ijx/6+x6ybcPLGYuIxIMN6JYaFTWPsLlvmB+ZP9zDXKrPL25cLWp0rhFbxwY
hU8+4B7iwCCNv+a5GDsNGNUX76yuLaT/17M5X7QjOwQ+N8fOwDZdo7w+fyOgz/pv
kYNKCfbYDEGCvUWtzg4uR1S4GAk+6D/o3l6/krsXtTobyWDvoQ/LH4t4DUUQpd1E
6I9k2YhMVNTZ3uEwPhH1MfPrQizkj2cueI24WeJBKqwl7f5q9AYmWEQ143/YrkTQ
xf4FOo2M8+HbJkKuFgAIigyQHBmy4hInNupS/QecpjZNhLNtCaYOTXpY2ODZ0SXK
jmNGvGXXVm8yrUdtUyVRzrCploYSTBCiF87HDR+YfTnmHzkX3sjEwKheARtrO2pY
Qey/dplFMsRV4RJlJJ8hPS29jCEh8zO4SzQa5rQq+BnVB3uh6jIHogaoDjXRkOy5
ixpL8Xgv4lFCYalAP30ZHUFnNuswgPyTMS0Y4ImgYMnMMY9XcaD0ee8eAdL506sK
OotAMx9OFFCfpkAYKo03OMwUvwV0mjc0Y1XC/TTmQ0GplwNq06h6AnkSqXskMbcJ
fUJi/y4l0R+d9ZhpKpugjmxFpLUWhkVkzh5RTKSWEl3zt0lGVVazJpwlSgzMpOWO
WIYdl9rvAKNFyGQSwS0CHED1GhaOuXsvtsr3zsj+gKnT35qp/5/XsLMwk56QNmHN
YP9wKQNbimfrQ+JTjA340JAt7hIDw5YzKG4D1o621a2QAiheJvlceWtK2i4yZLVV
krRoXKm+f3NCvUa1EvfhtIutFBVDyVHhnz1L4CaArhCQ0KLawCQMENkyA7zJ7+iX
3nB61gMGgA4h/rkZR+uKvMsy0DabdHOZeuNQ2NaMzOw3aXaXK/YQle0dLLo0qmwe
tXGmroiN21kJZM6/ua7OD+/l7DzKU1DsMY1rVBhOSGaNlrbt29VX3TXpKgVH3fTW
tXT9ylEHMWChuL87UCb8Of+sBkGFquO8XYChIOehKRgux0FZgN9z1EmXMg2yRP9V
7WZwkIpjFFLVNO0fp4/uW/xBoFcCm0c1cDbYQ3Fb171+p/5Evl5fu2YGVOEZ5DdD
ec8yHxDcB0RhfdNf2lP0x4iPB3x9IQf55LKGnfA0j3clZdeb6V4JeR5COkaE/Pqo
5pYzRHgBDL2zaiemPrhcd9M9YjRJMGTp6GO3YQfxJXHNL+615MCPUHSWyksUOQaH
EFpGCYUmgxUN/8hqdsihJBepnuegb5lCxBTkAYE9HoNmvewsvEQAKsDvz66IuqJm
wjDom4AGEGRs1I5ShCj7WGkKKr0veH3XtIN6D3l3jIQ2ul0EgFudJTuQAoAseUMb
cjMsYXfz4iybCfA9AFyHsxY6NX2zgrrg1srR8f27K70oI/nF3Y6MOwa62U4gXa7c
2Y77h+ivabQl7nAj1ql8tPN5rYiKQmh3fmcF4Y96oUm7i9ubmZkEizM3fY7+uI7t
BgIBVB0qLhVusqwCHZpSM1eG6ORQKhwy++nixeFnTVGL2HpwcY3XwfkLmrtN2zWT
Gyjg0Oq8JwDbTQa+xjsE2sCIjymbZLRGhrGkS3R7ws5pX1MpSQQoDyl4cplfRWpm
DoIws/t+Z+7c7+HRxJ4MYasAv0XsbEh3TvDUKibJ09xsLak06mzeRsvFsSUReWOT
Syl0+Aw0uP40MU0JceozI0zyASIUPlU0fjB0L7JgYtk9VBe15ZvHAk7U9R384gi3
sohvr4nrMJAncatOpt5IW49G2jEPX4ZqR0vOW/vBPxiW8OoGYJix7bMXxEic8TIw
WR2mtgdo36x2+GIdtRpdrEk2pGjxjMF7HZf4ZzufqwIfB34laXGfP3HQsQDMD1sY
2vyP8BnzNpDe7HrvJE7ZE4vNM0iBdEXVE1fvXKQ6/Qs0UlbhsjsA9sHPYjSi9AaG
2iuMx58l97ytJgpK99c7EBDsHkTakIjKw9kEYoeE6c/nIep/Rsq+sGw9Xe978rn0
uqZ/315sSF7i9EOeqYaXIgKFEOabsRESJ+1CwegQvTtGU9EK+3d+TECDY9vg0h1X
zxG6Qh36K4pAt5LLTUwxU4Zw+Rj/D5/UyyZnWPL76fYEvBDSXbxBUfpGRuq/rgx/
vqI8CDD6l9YDcvhFSRd01hRdIdQGSpxrqgYNwMuCI0rv8uncaQoDMEV33xqTLw9s
u1fP1tmk7fu8rCn54p4xVSlPSTieJ/d6U4E7nPe/N8WyTYxjWSbCyy738Stbz+8J
4Dyvln1w/7RR02pgsi09GLUTEZ9CP1budLxtT6RKOfB49CvLABsb6EBcHuD1BKNJ
q1DMb67KT4BbhG3P5oR4UZHSemjWE38yV5xfG2if2qmJHpeVCiAtnNxOXP2lcLsl
h06+q1mKB3VkdWDcNw+FJvavH3C9Pc7M+diy/zgraXEfCPucnHfzpSs0SikODIlK
mbpBbpQ/7NDhIwCOlMy301R2B11koEfXDFIzHK+ORF9EMI7LM+wblD/yVrDB2q47
LfTy9sPNyBWiAv1/V8GplNWL+QdYw0Cxa7SrGkH6ctyMlgVvSvfoNTsZA5ZlKZAU
fo5HcElabqRkoloaTeS/bScBHL/KaaORDhfBu30CGMN+NenZzSLzebMGYXrH52M5
g65yPwdonBaaWykTrVPmI6pbavEBEIuFe78xDxXkxA2A5rSOfjElVg35BzthUD8x
0HNB4ZHiWLRA22axZC8cM0s9LrhRo7eKteRxovR5eHhO6Bo6RYnzgCR5or70TmDm
mVhCy4X4xlyOyj7K3kEFcjIuyJpu4+SMkk8aRGSO1lIuuvbEu7tA9RebnvnLU+Gy
pIMG0c96QRfipDOrqmm4c8RJZS7IBUMkl7xXJch20/ldYugt+qHQOVUQ0IGPJQng
yQq9+1TNLnnbWWW2oGYDhG4ktZfW4jtTAnMfpKmdGH1rgXcXuzT35BBY9e27wm8q
1b0rIVHDOyA1KxQiiJdp/tuI/cAQsAGotFL5XOtDnNqkhqXiHU04zMfz2tTRGMZ1
Ts3zF5j/5x+LajZ2hrxoBzGDLVMho/3VoythiqzqPmCRAm43JLJfLSaHre559vgX
W/u7mlNtkqT28YgB6iWmhu6zj6AT4OfRukOCtDKFRn0ToLZqnSB1elv6h1y5W9RT
3bnsxJAmzPU3PJMpzZamgVuY40jYCHb+FCoBwOmVpDbxFdirESjX99QZ7XP0d6b3
pIUW/KwYIS/hnY5j8cm1C1daHZHsScXO8OeZyBjqyGoHg8YCl6jDGEMQfvSCw6tB
ClKyRch0q7C1U2IA6GAVenl9iZ/UGrpg8i+ic5+zkA/ZSLuqKalDgk7AQoNJ+BQg
auTPQhHlKfrxHLijP0C+NmhMbmDgc5GixP0Zq2Arp1/N1vAnrS7hKK2mIa8acQUA
XEY6mqNqHqRcu8eHRWRxTMSmvXhRrenycG/AgUmEMd2Ri2eyC+L2OugW2Fbf+Jye
KT2T9pZpBrmeFZhzy99w8t/b6Bi5wbwAMp5Y9xezK+AVLd2OV9/hUKsIXd0PbALN
9U1jjzdDePe0g2IM7CCNw9q6/r9f8+kYzoZAH/eYv7aHjtj4MD7bx2x9+rVui0Gx
FANcb7lTmYsAYHzfWpj//Nr6kHUmWpzJPyHcLa+jTCh18MxexHIiodVjJvaSA+u8
QjbDGvGtIoGoPsLmKxSHmCdXdxr0noEgIJCbDCTs7dH7HxgGMULDFbBQQbOi9fl6
o1gj+0mGVlB2/Jn8vFXFuq1/H4wnq2x3YEq0EtTH7rzcmCuhZm/HasC3eaEIw54Q
qKSSFxbnRQWjXePlN8eXjOC/MijwX79yDiKNF37JnWAYmJNC/1Fgp3C6d0PWdHox
OnJPaovYHMyU9V7n9rA6qoCLJr322kPRIzvjPWnHnLMG59d+8S9mLLa23eThLSv2
oymkD7AFbS57RyvvqMBJI142y//WpQcyr3Cl/4NVHFLA4SW1CWtybZQ4wHtIEE8i
iAJerflUz5RVclVBLi5gFv2rbJmpH+5paAMY73rHlCHGcUcvze+3rJ+51qqDmWrM
wqlfJVgpRDorbqspWNlYBnRJ6Xec0Gd6YKt4JqFC1BLPL9yi6Zjnzu/KvUkAUewi
GBKGrFdwDCLZrOW6pcTxkGO8EnP490gLU/N6rUOMb0nYvD7NGeLhSVC1+4q8Luas
cnqny52naY9bxC5imjCNYKfdfpnaWjHra0b5OFr6xsgDq+Zu4JNUuLOLwdrGnSUC
OBMirNXqsnA0Q4xHeAO2E/9OAbWKhzYnrs3tIwGD4qJOtTOceMbRdyFncYa0yzto
I8DKtwLbzr+RMNGfPfddezU1F+K1CQU2Jdxr+EyDCAX34zKPO3TRjLjcsFiMfpmJ
sPH5zAVxf6kCR/mHOReOZyxAmGKXZVVfMSLuHL/X40ou/X+IJj5N+LlTVzEzQGpn
YW5fSzQu6JnC8Rmlm64YXHqbARDYQsbRXkMoLZKMHvZz+COFm3qFu1khe26l0a2Y
UsLV6BYjZRy7vlv0qNKV2GKepW95bOFDc1Wh/RxuDCX7Fp6oOueqD7GTkAHvVdKq
hneHPC1e0tr8oO6MVVWskWwbgpEbuWs+IeonrhS9BoY2o+nmCDlFQePDzjF1AZZ5
em7niMGgpUD+aUD5sr8Y9lCkJs+jBQs/2PN4KtZDHvAeUHuUBfBp6dllvFstOB6L
jfQ686zWfRIJPzUGvvmHmYVIn0ESIesh/xG7FFxhxutOM4hqtl5PkZ+47/tMSj13
o0L/dv7zlHyTdLMWiJqHOiDPEGGk1uGGwGLF1h7os5uWXlGy6XjQl3TUjUww7uJ4
I3IZtxddBeVFIdMvO1f0JlHd8BdGckfoYw+/QIGRmVUPfWN21xbsgkXyWDZNtVHw
t3tkOvCTDX+tYno2LweaZj51dNRDW0Vyhjft1Hdd9FfXI09FBdkUg+GwZI4NXiNk
5DRANvmOe4cWxfxmlio9dyHlKIUMzV03u9WxJwAX+L7zv7avp6NEGaq2lKCsZgPT
aaHsS+6WZRcV86S0kc8X77RgwFS6cMtj+fNnIxZV/SkkYQhuOzsx8+FfK5OIenyQ
piHJf5dxc5OyYox2ImUEDZvhBfuXUyo4MXHsu6lsE7eztwKXliw5Jul0YThGeqno
8biQM2jhOnrUfOFFX6+B46J9R+JsV2yz2+DqOv5urwtOGCHtHTyOxrbAx04ljDRZ
xleNQB3/3EqPYDE0B3YfOEf1PDEpPD60S1fILIHnKicgyMkZDjksQwh0rFiQBIlX
RF8e7Ga930zDHbjw1tq1Qm+TfDQvrKG+LnliBWe8AK1aJPcgN+1FAQjFFJVNg9Wa
1Fcuf6gRGmqV6p2XdQ58/FjCNJZZDZhQ1wyZxVqxMbuKVaANB1bLiLCYW0RpqE+q
hY2bqK3aoSc0m2hLOoln+8mcoZNytdxkOyqtO9JGEEsO4qHUhXi7TsMKeom3nFG/
dRzNTEKjQTngZSaiXz0r7A/8OTxzshQx9h1FfMaqJ+aXH+Rzw7Wx139aWtRRmZHL
8xE+xaIyx8uH5xVIIQngPfCzXXVSSIXc4LaaDo7S7ORYiYsXq/vKMQfyWuXdPE1p
h6mT7ScS2eHP0+Kj5W4HSyOSo2fhMjDb9hPrqV0s2X9qStaYaBAKTcGtjCrhyDQd
YkbfV0tkPc8xnvdB5ZscTePH/3n/BKyXYKc6t3ONeZtqr8B+QrCRELBpxvaLK0Of
1kcBmmhrDgvf/2odgEzwpqGwOwKMh9qPDWkYXQicFbYiz7wr02+snzQuLBIUGjs6
uWL231ZE6omuuTQ3y89bTKL3yfVlKQVped+g3WmXFie9XuoDg+U1vIAKn4+YBrhI
ctOM1+cK84J6nPvccJV2f/bR/65pv5O7tYV1bO1X63p2ihe6XXtsH9015KTgeAX+
Wu10UMpeNQHMRoHY44xLY4QTVq6BKjFvmLqJf9Sxw6sMR3nxxeWRfoLXXlOQBqC9
P9dbav8R4hKxEvNHm5p7kZGLxo1drx4WG1RdUHnXJxnBbo3CgclkulxcCgv+Dhhd
40+u/cai9wxj2U5BecvHiW1gswMpZisPJxIUNlvTcy8Q1idLlgYRg7m6G+cANeCc
mYFlGTvYaVbqzxlgohpy2Pscs8Egs6M9WbIDzZsIorOzYzSF3ff6TbAhJCFO8s0X
0+tQFkCkspE6Pbvkf/CnDSVWJ2ooyG3rVK1m6rXMOdhXsMEFBNrhTNXYcLADw5xM
A1w4Pxmc/6ngJeQJQl8qNaaUrEwhu+JB62VpGKBkjhpjAELjaSnXjjXWYAEJNxi2
zk81NsCJW5y6IxeMWQgCHV8f5/GKThEMcVB1Hc0OG9OPQ32DZlEmzU20M23AF1lN
1tZWW9dN4um5T8TSVpigByye5j0idmaPtD6I2/qfDVkaER8vEkQ8P+/bTel2+TM6
ZdvM9DP/TCvqJM4wA2E+aleOX3/MQOwLJYcmXw1RCshR83bwgHcSIDEpzEsx0QSC
F99A5cosRy17yORhhLU5BDnazW/ntO9b2hi0hgZJ4B7KNwe5i3hRPuKWfgerI2m8
OoVHyY90bLRQe4oLTLvvCB2h6J/O4SxKa87RZ6FBajZx1+pKBXwZBxL1o7EO/15v
e0lpuSWyc0d2f+e6G3gbRmp1o33l2W8lY1oiqs8eE9tAafWBgyHpuyr1I4aAKqyy
gIlumP7/YO3ABRbANOte4XV2Bq4GU5jJ1uH6KsB3D0VJqcBQDUUbiv0BEbHFuKdo
DXWnnKXu3dDVrUU3KAh8HyDLUVxw0QvY97KU6BjvfaGY3CIXp9NyZx4VNvTRH0e5
GaPIEISe5dSfzRhQLtkYZPCExQXVOfofjM3MdXMkbUwfVE7ttYuGSUvn0E7jowkC
/eR3PRX71jdjcL9lP/7NhrP6pwmCSM2K8M5rEnyiKdjBZFJWzwy12E+1E6Rq53XO
yhXvQoPrlxniK8ljOIbj1897VD4PHQAvgQYrUcV4q6A9tswIC0jqUdC8Gbpou5kf
vUYvJ96QLks2zME7VICK/5SISQT8UyhognzdzLn8hwJefoAZy6ALEyNf5q3/xVq2
cmxl9R2tCaelBQGT3ZQfHICZJSHkZ6BbmHZH1K3jvlAso7b1vpujaXsJN/tLkLIp
sJ7XCCK4jUTXSz9x2uRoZ9wVwwZfu6zRWmrtXm0mc/D2EGc+yZtw1jrW4WS4vc0F
rDUFRZbEYvsAPYigVmqAe2JtG8yqY7/RJimGBBnWnsmv9nfD+d4z6dgKrgcPcYeL
3x9PdxmcGKeEw0rMAfPINOSndRJd4hu6jBeuHdIAJBsJu0mjQ6zCq8LaxDliOyqx
3bMbun3LUw60xOG4rVYRe9OcJKeWc9BSC3kptLi2uar7pXiUoSoLC5lienAN/K9t
/UpN47wO6wC2aYgXcu9xDReulaT1tWr6qpA6RtgUXEvD2f96FYZ42XwDNJWSpReu
l90xYzU1kSMqmfHaGSNa0MTQYBi332iL0VGnNXYWeGiYq9ZhX0lHYlIev94cZAbF
Pi4vkaoN4hfEjZ1J0eZ2Iubk2J7AsW9uVJE4ckq95XtskrmZZ6NlSKBnQudbrc5e
AHW6G1Y7wHsGJ8iJSqyqsM3l5bWi8QKxEIOIBVv5voEVPr/ezng44UMXRS6uCXRc
HIG5v/05eyu5YmMfN9ILtLmsp4nIjpw/yUE84s/Fp2fSLAXAExE9jKIYy7FlLEnY
UATIrEUr+TiGc+Q5KS48s4/SisZ0Wq7nM+JiuZBr2E5WSt5fOSYtZ4L+RjgT/OJw
g0qwDz6o5XS0kQjzEEOoL1B/ASLHkWNJIvAj63mCjOlIEqMbsmJUXo4zmlW9ZnYB
kVaA8m1l8G2RmcSlgNMyrvxYO5QFx4apEFJWxIta7YD+dAmyiSu/x/Tci2sP+cjS
2SUBQa+hxzam9delLG8wN40R0j2ogYL+VYD7uFtR578EwEzBA77AH/dRvIbWCsds
RRv8IpyqpBlbkJDwA8ME1d6Ho2ZUPOp6mO7xdOidq+oEGO+OlwMiFLztqbwcXbq1
/5OiZ3ESZoBCJiqrxa0A95zCx/Bl8aUAdFtir3OMZwrs6nRfc4CbPP4q7LPv+CzM
PXftudL0ok7mh/46d06m2JdImt4uYmayiRpbUo9ABQFfNlxooG6/a5kUkCz231Xn
9i8+8QMsrU0FcnO/gb+rTfEq+Rd1q2v3wip8rQa4fQq9CYn+0QCz44XwDQNP5afQ
ioq4uRkUzW2KeLGE/S+QQJpXUAw7FbtBArWpc2EdiDuZM8El28r2Wf4DsvQMzhUL
QDOZfkkNPhoaAoJa46pJwRsQbH8u8dKL2Hj4IxghOyYc3kj8C3xSDA9b1/YiSTAy
5vUgIZGR7AFMYZVkDJVaQ5oEnb4D4BQjwwVAwuA8qbCM8LkGsS9RpVokB+gvBl0m
xB1cPYPekmYBjjh3sTrXUWlilwy2aLPGaHHyrtlv1alELVI8sU11y/ZXW40a8b+8
7k5mNWS/4iok3WjaIcSt/4xko1csRypsaOg0jLNMjSiBmxn7xs5kyM/YpRcJ50Fo
ZV8VgJq3NZ2aska9MJLVA8aqUolMu5/oT+qFxKEFY266sZyvS4xmovwZTethUhOV
WScvwPoy0SAsRAgcmoAeW0pOlXlUSz3mzDS+K9lXcusw4KWQdYraBEcjR5sDMlj+
dNLOruerYPtt/aQgEMuz9mnf7yhg4ajyeCOY8Nfv62gO427cJ1AiC+cDaA3kh/Wc
OuyoV7xsaaeUJddsWLWLoRlKXr3EYjkNlYuq4CM1y7hCHkrS5q6oB5jrs31P4uUV
g8sgK2zz2jDg1XIyyqw1J3i7Y8ktl5yS6puYit6tHOR7CeXeSnIcyS+mspMHwxVy
OC/JC3yYe8N0LqVu5pNfN0r+7QsFVUXZqw2PKDlMyyxcejzn7TBj9ghX4mh+VWpc
2uayPziBeFgQvo9g4UkCNNU5o1pC0DjAE8yzfQQdfXJse/SRkCwyLdAmHP7MChjh
W43QLTQAisQ9ddyZdamodugjjZaai3QL1M1EfVOnkP3MU52jElhtoD95CM7ORP6I
LLe1MqnDEKo5ouGiF8TS9VrD+d6WoAn6yUSYnhtEFzZjAb9sfjNPRaYbkcw947Q+
bnWVNofafasMrSm4+WXFaqrPhSLAah0vNi1FuR2f1Zb3pKR3OArQhk56NkGSs36O
r1uY1TjXpYWj5Nx/k5XdMepi/10vX2Jtiwh9kyzE4oaJ5ScM2EixLQklh+Yq87JS
rP0CEEdA5R4CLD2KiFprTzDDkitAi5sWOzM7PRNf4uB/Yw8sATPVovYHyEti/NE8
tBD1McUNZPZKv46/Sa8Aw4UwLhxWE1JGnTPd2jwKDlUBA7Po/iCrM99A565Ro1jx
LanuZR0ycLVv+lpg74yGs12hLp86wA312e78Et4wjN92Z6NxkawTeUDSOiDuuc3t
Rl63KAMfjp/8D2zo+QjQFEmzu8eeeq0dN62TN2b5Iaz5v0y1bKskGOZj/0u3wKZR
84IRaxjskkz8pLfAI7EmyJcrXKRHPZLX+EgMhVfS4Rr2qb+8wnDItUgcgZWnBB2+
ep9Lu7GXeNbX7OHPjf3CM9OdcjOmkSGRjlTICdGuq4yKQ4Dj8s1YmWMtl9w/Jvbn
tF7oPNdbD+xklNeC5Zqu8bR6NXG0Kemi1fWtXm3BOsRJuFv2fHjg9hATou0tqXwU
rQcxH/KdlUYu+QR/9+ZaJcHRSimxvwjiSKwd401Hox93JuzO88sDWOAV1iQdDZpK
oT7UL2jWZhYpolfk6tcs/hO85FDoYQqIOxUvRg5fO5xZDoxg2WzZS9EZRHahNmml
H+Z1qp9xpVYjzORjYIyHUQCtuhgCJCDULBbak5yCH/k/ivHLN7x5tgrYCap/qv9P
xckLp1+TYsARpkYrPKiXCRmajNBByfnn9Zjz1h2b5Sjk5Xu6ZsDNdO/YmWf/WBn+
P/MUJogSgrGRa4CkUYP+Yw9M+WhkkBJJaAbAC0iasARLQ8AojB9C8qZEHHjxOS1D
N/ktuLbAyC8205lFt6aZi/1pVrhgO6KQJanNZfgtSm92MY2NwDseI+Gd05Fw9zBu
/t7XOzDAJkicYC/LvRvUme5FHImishRoBeusJG3xhZM4k/2OdEah8FLJokI2xteB
E0KNB/U81vnLaxxADVpjKOibsSQ+2+YdlKZ9OoonZOPalWfb8+qL8gm7Th/SNWnn
hnHzY5uzyoi2w11F9Gl40Ij06KpPnrHsSzJskGyn6megMJPlJz9lCjcYe51OyoGR
Ocwk4hn9a8gUXFT+izWKBw4Mr7JFHzKfQy2GMzurxId9564OenZK9sVeCT6AGb70
SEODeV3mrzeOeY3apTGga3etcRvpvwdeRdUFC3lq+FOmfiS8fekfBWgYexq7N8nF
uM90UvBq1jWvsjoBOUzSiBHGyyX2rHGz1blsvaLzDtUVovqK2J1ZnvGScYvVmbHF
MzD+fkCwU79wA3CVpwfZ7qqcfqtVBcL3O7l7JJZ+UIjY2di4b2EDvOjPnJL2nBN8
xxRynq2Oqr4czBBHXBSGCHxZ4IiXlNWZkSsnZVEioXNW3JGv/67ElZuR8NLr5B9Z
LqDyc4xC0dgIEUq/rOZpakG5osX7dTF2rQiz2XtREu8tionfaLxUaez4k7hMpQfl
MeZ2RTFZwCR028tjBXPzzOz/gND2wcJuJNCcCIEZmE8wIml7xekR0Kk+n16tao9F
kA5Tdu1Nco4XIbT6TXpvbNnj4PUHarxC/z94skRJ+RX/CBLk9R5QgxrcxHcRLrEa
riRLHEnVa88MAC7Gju8WX+4Eei4gXqaoTzEvx3z1EqzVJQTx6c+wEqkuFXT0qT5o
i4+9Jyv01eUB79T2nGoQtJmO0bNp9MFGWbcfNDUBx1D++o/kmdOHbgbo4MREAXj8
Y3yqBf8MJEAbrFGbqpymxn2XjS0eB5mwlx9e89+iYwFjZIfz8ctnQxHk2iJlAD20
Objhkv03mIw2tgZ+xLVlauXfLxO/R5603yfSIizOTBm3F59UJhZCtlY/GxpItaRn
renGHWzv8NjbZYHKRrtU+fTeUzQIJnw+kYhvlnt15RXCZvyYsi+6lMoDw3F3mWWu
r40Yo3R/DFyILHApKRFmWSHMzfplrfqQ/+ZNFNb+FBZBejeSbW7JI3uVtO0tzw71
afNkfVUqWx7zcS/0H103GmU1ZEr91EJRD+raG79TkcbRyVi4iPS2C0qtrPNznJSZ
kkK4Mvaku2MWrjs7JZ0aoALOYs0c6ouEipGagtAsktr85dq8y1lBlfV4fP27sLRq
Iw3Frl0cWwITz4UCJgDfY4ykwx+pQ25mbTb3kAAJ+g9Ntej1j9UhSSxlBM5ldDKi
5j7rguslZvnwuwK9YVlq2q2/zJMiwHFizxrQ5QVPAf2PABjrQ3RplRDTXxDlqbFv
87zA7bQIcFye/voUfbaSjglfIYZ7kqFc5T0BvAas+D2T4exgPY9L6uHjOOetJ9XB
g7O+Hmy9kNZ2SwNG6g10paAjAe/sL2Z2N2T3oMRWcMO1b3LPM7EXCoT3iOGvcBVw
TvUvlx4v1wZLdRigp0TLNsWr4+YyUlJ+BthoDcADoGE3Pg+yPPQ6OlikKzG2wRnh
N/sjI+jH3qR54O+q+ar4SE7E7DWn0OUcgpwAG+tEv5EoFEjir5NFHFR6thl/Sqn2
hj14VSA+AQIsO77J4j2u5VHNtvLTfIwOKcA1NwgRo5hoxeqZFibZEQkrZtwtkFqQ
SZBRmdBkWPJWqitJZ+EG/5IBQgQNcKyXg8pBZhHLk8C71AJG/pKV0NYjvoc0b+Nu
MkDVuBQe4Ksi3NSd2J1viMXtHWSqvKgLbU/4U+OLTK9mmRDQhKdVkaTn9uwL08e8
Y4XqCH+L2QPKNpqYNO5Z3IP55RenIB10l9lQwhffGIQzswz6nXwuWLdar6xfkJqV
73q8Z8b5H0Yh4xKmXzi2BowsExDuSy0Bq7+wjwOkewpZ1VRcQUSpZEEG6+XtH+N0
YK/h/XjSMiQnb8K3nMkx3k5/U4q+oQy4F8PVTHXD6fU2G1OaVvR5ZRG1Go4h3+mq
zirj8QiP8KgtgILUwUT/6LMQD3lEHI4OeLFeWyt00l6zD7W7pMiSkRlkjDy/1yO8
6ArxwZODh+B/0yfUCkv2opFHj/6+G6WzEExzYedVrqUJAwRDoOZmaZIjTWP4gTcQ
kWCscui3g5M7OiGlmBTr9CHjzcrfdh1ud8qzI2uI22uBH1IiUY6bI3i1V0UYfWF5
NHipajezpWGIsUBmtr2eQVRqY5ZyIpGdYmayFCjWuIPE9pTFECYwjepwplhcK3Fh
Q4591ZYSR2CZghdMFfEG2uHxMosUm56U/iSiSpzoy9UUd2IoTnX3v/v/RXDCudHh
BFgjtv7RCbOVtIQJ9HbHBPIUuSXVcJzT7Q4lMioggRgEPhnB1o2oMpB82sGhhuk/
ZRimfaS5ylLow8Wv2jntr7s38I/gziOnQU0lTD0nfteMuEXhBhsunpeiED5xWTO6
VGKCbguGY1oZPEe9xDkJdCwuLTa3sBKCa0paHzUk+oV5h51ePhtpZpOfUm8dIXEt
hj8pzz1mmi+NFz3tGDEWGBIkkJ6R+zmIoQbxLF7J8q3zHOdDVASq1nCVWnKFmssp
TdnJ2bzX6wIGSvEi3hDOzC3fnaM1IXvBjRx5A4q9GXngwmwvfwH57UF7fB45Fgz2
qjYX8xEeMLFKgmRr2mDNnXSmObqpLacSWJXhhTnvgYwoFIpfNmnEy2NHZltFSbr1
U2bNa66HMRIaLvEsjylTkXSG9VwMj544Z1/qISPt47lG1s15YCIRpMsBCM0J0pCe
7AxeyqhtCfdgzWWCUrOidC6NWXTdsIF9OudIYl3lHBcEE4VvlMF3PQJ4BuNjzmUi
rSIegvJJtw1ma9S4Lpr4ssFI7SreUOrPDnX4Wiqz+KAS6XWkm4toAHK/2CxuqSFI
3seTJ+MifvrkvPm2PoiGIXkyypK6vdT+i9EtV8/VnYmcrEIr9G5WzBrbdE/IZKAf
UiZsKiSi7LX2s1acdBeX+4T1p7y6KDiVOt5baYvWHbwRG/L3XGgaLivng4uer+wp
K3RhFmiwrVvF+8cJKlrJ/kpp/ZtQcyek250BLWdMk8ZLtDubdVxPys50qYBSaySi
7Ig0TxT9SA0KLSXoK+64/o7CaoYq61TiSanY8WOBXvny7vtsZMixaultv6hqdDkU
havyEKyoZMDNzuvq0yHt0KQ35mS157KBK4euf/d79n+9jbyI/9STACzB2tFXbwxz
EEHd9k4F3nHHLu0/vWRvKGp082Nasfe6pe1lG3WelD3CCRJusXAbN50aIa+hVXQi
8qfN80cQhv1kP3BT6VnOx31OGUTNElr568qprwyt8ks6mo+mElNWLebEm/SBeH/B
WsOaO33ger9dNN+e26K1XdarIxez7lh9ceaWQ5EZEP+IS/E0IjDufhsHhBWisr2M
pyS8X9YkC9i5INypEcijTer62EtXTyZtBFA0+qk1VTotWJRUk6RDl2S5HaRbEFCQ
lrTpEeJfW/HfDZPv9h+l6Nr89qzcwRzuMAfQZ4jcFJqfioT8F/1cuCpIUVFkirap
u1fgLh9Dbnjeqw7TBZp1Wq48Aog4U7J/kqFNxQzbhXGbIrACpyKy6LcHfTfbXDsb
50bqqkW3Z8IJEuvYcq8ToKHCYbda3gYzsZHISUVtRPazqj2dyVPiWmS67k8Tw6K9
Gt4iO8BJWkKFBg0n0jkPjh6QvMcUHXtAsqC+DOMRXfcPSnkyG6FSA6ZeVc1Qq2L6
k+rjUwY9JV+tTZhn01D/nvRWiJW/x21aUBQYBGdwUO0QlerTL/oQABDezQmkkvtw
kqnKyPEkZ34df63td80EhcHQjEEu1RO9KyXjAQw+Tcs2sfDNIYpbm5U9xsKTLQig
EBsMdKpN9WUluYkmaef9nsTgzhxBwXWgK0GR5ZUwlbEE5K+QbX5w2J5zWo82xMlG
+xafK9vPY0jUFcCHSK5VHzAYx4wPwBfa8kjUGSl6ECq9HiD5NW4peXpDqQOm6vhN
MyPWLSLvO2cjsuPaP53AgC2psY4pmRDF5KTjD2SAleRfxs7JdXe/jVnS+WgaJTe1
PSUftU8O5Z6+xJkbttzkR8AY1XwAz/bNKKrlc0pl+NOD5NWxhpADYAuHTvol+pXC
lXLBZQ+3QXil2Uby9dKH6z4GdcJ+JBhZYM2rYlEs4OvGUbVygoSMD6IdkzraBjsc
wELZ8GcqIHjaRwuy4Q0RsRhj6Gvvpdxni2n5xKLs/xv1k7Od/PitGaqYbiHabNGl
8xQszc60/VKYVSoBBWkRH0+cgMbgUw190KJnHgVOK+/jIZmITBPv+AurTkvE0foZ
KZiHT1j32rmv6qN7b9k2tjgK5Gcc6B4unfFJ7H27OVXsRCgh6VGXn31kdeAooMgl
OinmxgfNeofVQ4HK9y0h1hJDLNZXqCFfpkHWFiIkFKZFm9Qx8dtwEJVmd1GYF9mN
GvHOzy8jgKw/b+ZCP1NnBfZI8+fM58d2aiDiVMj/gxq9x1LykVTi9tyFpoFYGj03
R8b+mI8UnCtVu03QiLEpTX8nIsCIGbak0RAO/w8nRTEUh9ZybZma4MbvxGyy+X6K
d5w22PA3/9QXNf9N744OsvghqulN3j+CfwH47j5OHTBMeRSu4BH9kVPGMoBiqrx+
31QiDFDIV/v3AbORbplvSEs4jrFgXyTZsrYspXdy2YBh+xaxQb65P/Fx9ZzJrowP
/7x8vcFDA1bF+CLhnsOsKcVs9zo5Ym9pAqfW24rTa3f3DkwEvSlyhY4Rd3mrvy+u
tZYg3vUjVKZkG3xf/fT1MWqPcP6477xjOPqimanfe460Vwb/k87Q5j3gtKlgrDAs
4ySRmHihZR6fw3zRzV38bhtFTgAj9Yji1dvw+YnBrdw3wffcxzoa7hxX7E4WVLym
aS4yYg1i8uzvut6K+LaXiT6IVxNdhPDqvnORdm//V8Ie/5Iyy4RoAYNUoaztJctG
PFxY5LMokfaBLOMF7nq2eS/VdVv0nIKnVHxidqImdV56pJ4YY/bSa94y0JPsWL2V
lEDTYzgNAuFS1Icrda6bvATyd6puM0xapowP8kyWJRovfM4ImOpAkYluVxAKBBvX
1H80A/hFBlwGhPR8D+KIIlPFC36zXK/Zy0rSg7NeYlqKW+vr2Ip/KM5qLCREA0LC
XEsd7PyznS9suJFwOgRbHHNcN+/QbceLtTyelNyOg9xiNnWW/f97TtfyCx6GOyf4
kNyTKnjyEyGx7Se193o8Vf7IrlpC37VSwLXzkgK42M7qi71E+wDP4sOA+1ZTujr1
E40MhMzVNjTN/YoqnZelVROQDAGut7Kd3zb0B5xjkLJZ/hu/AP/VPZvJVEZEdwV8
PmG1rpAyZJpoKblBjQN/1e2N/ixBS8864GC9WOWCg849bB+EYCCq/hOzlSSQs35S
wzvikfKr/XUoRG++d6S7Nl3P1gYlddTyHOu4axbc8au8CkqW7nVhGtXLA/ustXvb
zNdcnFztYrxf1mbpII7TTKYOZvpETybwDw2Xg3sGNCaS7+VSkCpI5MZbOwNjDvv9
PDa/eyfs1yYLcaLMqzU30UPvMGbfanR8OwpzpithhqlEYqpgffpUt4Cb+gMDK4JH
hMTo8Qgr/Squqf04gOTK1tpra45EemI2ioJilXsxkJzq9gN8uzQNBG7Iul29g91P
UrY04i8vE4p0YpUEpRkO2DgKtKjSIIkMgBZEM6YAiYdL6SYtwpVyqeAYEnu3bbbA
tr0ZITMD9GPXYxoHHSlR/AiANI3Gb7rahICqM7Rq0BJTS4wIKBp2alRtplIBloM4
imDZxT0M6XFHU5Cwf9XXlEqECRKq9TgCSOvPUeL/rE5gipGl1Y3phuNoiF0KwYr4
ONkmrI8fPkjka5f11kCEUKD3Vyrd9JLUOtl03q2M+yurzUt7d0QRYHRDwwOu7brB
mL/6214WOqp1MbNBvoPVzxJyO8Y17Sv7HUSGQAt0DZf202jOLcgBGVHz6KUtmkYH
N9I5A27E8BpmsL6mRlW4ViTltv5mLl1bqjW8WT0Y+EL0tR5b2uYyUsmhQn8Trpkp
3QlOM05J7UBFG2uj5EfsPXy0ZUmZJ8B69VPuXeDIjVd/bs5xBOsH7XXVL8Q7Bl2v
qtamVnN9dZ+qw4KLyxJUFJIg/yzeo6yUqk7LBHmI8Gxl+RAYBv+JsOSO+6atrJzM
y81fcU5Lhi6YNHp0UHJgDo3M4PTEWbgk7gWN9zdvoaYMg7e9nhU3UkYzLDnBHURk
S3SmfmeY6pC1P29cQvskn7JNGkQrU7F/nflLk6b81CM5TzHYtubiJoLyg9pPnkHG
rZZ9DaBpXxcIaofxE2yxSH8AwZHLzvD3rz1FDmzzyeExx6seqgkvLlnBwLPvd2BO
bBl2y8UyTUV8tbSJbiJrNNJnVhdDmBAA7nKClewzd3Ycp5qk5JwiUR1gsjUvV4TI
VTIAwGvGZ+jFVazkpsC0d7z2wiaPjoDtlWYIeWNMpzyfc2HjxZK6Y/eaSYgej94J
VJK/ztyvET6tokK66DvL9UGp/VYYlEUP1ErPu2D0mojXbekNTR/fU3AJAL43wycM
11MwxiGxwvsIu87a3dtr3pNlxe0pfTSn+X8o2UWC9kJXil4Dojl82jLljJKnTHSe
I6T46p/HUtmhLtugrnrT9wmmVnhY1DV3UDXcvHA/gIwS2hCp19Ht8b/gwa6QXVLa
+gncXzX+Pvn/yr7TJ+cw9SRG80PAFfgk/syiveJq5pUGPiQrjvVKGP9rcn/r/R+N
fl2ZzHYv6Ul14Y0VQ2JkwO2gJZgqxPG2vAWuf62iUzSO4mVQtf4yu1T6lsAGWSg/
LYIBVMnkMj9acAho8gPnh7PPFiN/ChhoXw9GSur9WtXET3+Q75SECvV3XCSZkfJx
aQpAKxr8gX/Mvyq+aaIm1LkVFGrrLNHviFJCBlouUHY9j4GZ0FpXbQrVLFEE8Jx3
bQtBphUaYMDnpTDavsi596TOW9NuDt8O4yUYWwLPxswHxp0NtVX3131xo+gsARjR
35hJzRCj9oSc9u0jOrwhjlx7wv/dXJEem3zWQ2WBQwWlQDTuoD2HHJefwkShS3ge
VWSSxv6jCBhJSorsTSTTmGwyouQw4LIdihLXmXuH7118xDVEc5/lm9WKq1ooXdIJ
GBqzOuA+Q9d0yRPUB5e1lift42NbYuv/qW5hP7b8q99N4mhmVvU41bGHj3AiLkmr
VPr3sH99/hon2VRlpvOUPHbi1Gj68NXfimlhe9wUG2liSWC0CvLiOqjU3HBZqiZZ
q71gaAepc36Tm9r9ISJ3DstGZl2gbyBihFg5C6mJgH8vLfzekhTqfGfPWf9eWA2y
ziHBq1E7aYtFUMbOtRC89L3J7RDZwqY6NMAF016NP5F5boi4lzhtRDEBaInJzse3
A9/7G2zee6dAvAyQH0qJpsZVsdB+E8H7QrSQ7HPQ1dmcgBXGT+ZFyKpFQe257HOR
Q3VKqp21QdxZw+myCf+nTemq5R4Lm03pk290Btebrw+ym5qKwRTm7FhbWvYkvoVa
kGk9+sHrxBNcIkkTX2sZV4w8d9RPePkvoSOVSrK9N8X4IVaDHm1ZSDWOgEZXESRN
K6Ue3qbM3UtWARF/6G/xVTx4UyDEg55HWL604qF2cod44LWg3xkIBmR2eA4gVNY8
4vLCHTPa3J0yO6jaM0y1vTDYZjD1O3bFq7nKnCdjvNAC9fvN4IkoDdeoYJzS+MWB
dhd3Fuy33CliC7ENcybDQBTMRAOqQICaaZtpjOwTSawEalo+5vqJqqQiRKQ8qeEs
+LWhWUCmvRZdtJe+wx8KBOFY8PsUefw328q3bH4SZSMcPU/MWdgz1Pp408X4RDxf
Fl23m/VkmDvx6vuGoS1KxyUhpN25bpZjhSMAMHPU2Xy65Y2YAWkuA9JTBqWl+ztz
UZ2z0lIK7euemMrtve5RiYMoQwhGUlhB/B4G8cYv+SSJblT7HFfuIpZzDSxr0pTE
qtqX+QWBXDjRjgjBrPqPvGGcx2lMtqaoseE822XdMjpnN6uBwXGKLogI0VtSoHqK
A+LxZYiofK9V+sO8YklpJzS2nTNMw2ndaI5vrFOaFioO4lauWjKpihEcz5pXKEsN
KR68zGxRoy17rOxuEIh/qqJlrJ8JSQ/D2P3gl2129zxnpPTq7u2yapi3ObWEpO1e
8RWYlgwUilDGewNjgfU/4gsfZL1VtiPzErBg9X3EOL6zwGuX5SZKYOzWK8Qs46GA
p7cNAKPBsNrfaxjEyiiUAxt2fWdAi0X4s0pujd8N9/TlMdJRYZXaJdTaygp9idYN
+1x0WfY/C7vA1fj5ZVfw/+82GXqxN9UogTaDIaq4FhumnkDsgFLRSWC0ur5vzEG8
4gxZAFTBTchtYLC6UiF0SBqZhkgUtFLLkpogi0uv4zcvPlMEPnHqrVAXNXiV4DBC
2EUXbD752ZADIGSusdzdb7+55D1MgCAIjJIL506XEXVHGZTCUMFtKi6p88UbVsU1
RWkwXwtovZ3aEZPTrtVv0mMLN5a0Z5WEfg/9sncKW3gMTM60tQWhoBiKWHUOi8KC
4AZzg3ToVP/PD8CDEL6JaxAlrRQ/VlYIV6FyKJEhysilM7UUhJSxe7DLUV87L82s
I6DaiM4NJvbILggFt79y2+bMGzw9aPTy3zGtLoDnW0IypzNwqQSP2P99UsumfMV/
ulH6ERy5s1zkznvatjIOW8FIX5Y77DS00VarKGMCkt15He3rVP6+T9TXFgwf/H2b
X15F634Jhb5puFBuBuRfFa4dojwbct9pYYWoMMcSJQx7WfkbYfYm4ZgNQNFQIdTr
o85OMSoBHj+R2401nX0BNS9oKaJFHwcgZD4L1JCP0F+C15lLfvHOFZo4Bpxcz8KB
onlHXEO+7S3G9206bjl5jdpr1+Ddk73DZpQT4HMLODIBPrGsaoUjeEI8hxx6vZrq
hv2UP1zTf9gkLxIuulGxYS2fcUnoptOY9w2lrJ1OPLNBn3+iPuIKRHOx9Iwuyh2h
OoFq7QDSJ1RMfmTPAneDI3geH6KoPsq77jm6/DzzFcsw4PHIgL/fLRlJ1D5PxMZN
aKrHnQ2B1eM3pHdWbxH3IKWGgni73RZ+UwcrAtPm1+V/Dyr9cjwvFapfZcZtiSru
yt4Dv3O4xsXq6g+ruknfIWzO7BTHQXp6jJmtXsnxWhUM9VMu6JNHg+AyMd2ygeRM
Rht/s56nw39tZUtCZDJ4BDaJZk81oNYd0pxUR9hFBVIiw68KbFtZMtj9ufjgGk91
bEU4eSnYOuXCVgeV51ILgw8//ZE60arIDY3uzr0B/qiH4AJT0p0E3pHP4w/JDgHX
k744/BGcCs0uJPWWtfIbDa/bIGGO3OtXDaQnhsfybF8w7qkOfzaaMRCUW9UOPsZ3
4gBFsgysEicj/9wY9JSOlK1AJS9PSUO47YecR/JfaDDcPKUoeLa+FlIZxY0LFg1t
OduF2XGZFWAkEaPGSweBXpK7DCJtkUgCr1Zd7WW2CjGGlIop4Gz7nDh8ZNuCUjgw
PldlpfFVp5bOAxSkyHwxd5WQPv4Tz8/ChiD9Van609aP46sFKP5Y3nzbj3EDtjxn
6Jc+KW5p/i8SCYAN4jzpDcnl2NE9udLnYblkmXBG4sNVom9tNont2fPqfiE9Bkl9
sF9DaVtMQzqgC4SqZGSiEkD11fyh6Ynx1mWY52IOmtwy0KxBVWqRfYWKcWIrct06
PSRERd39onlmq14QqT+7Xc5Jl0f81sMpouvem4OyKNwfC/bLnfT0tFzVzXwZ0hct
7xW9RJ+IP3L1juYLWTHodEz3j9zAhyuSsm9vRDTlBpzz8ADcuF+TXDMfzGdfKNmF
Yr8g0YVrRMgIY4JqAEzHHCAIUkY3I34Ph4LX4tDit/fv3oFDTEoXUQn/MYgy3IB8
bU7hVE6X2ByE4FJoJIB2SAj9ULARlyjZE91klYAbIbj8cLshrpeoO+hL3VmY++Il
MxXWIu+vuXHa1JlDG6knlX7PCgDNgwNcIaHz3hyZKcyymyZ0LznrhCFTnUp6z4v2
kYe13aUOOWu23fN1bwm07kQpWFub0N7vhMOFA8WpQYpsWx0VqiFpymWgaWofI9Vy
qhgbFrUbH4vV1CFqSZQjpOjVCkhkVCSwzr31+VfPeHJyYHjFlY4crUF//IKRmbpy
Dkhqs6HATKWXzLv0mWGtZM8f+K9oOq1nvWG4o1RY+hRcWOabmkhfZSy5QjcEtrsO
r/KRMTZ0gom1TlufrkATiVBFvij/Gi5rO+QgcjqM8I82EvDNkymQylW34kHUSQXC
8m6m8LNcQqZwXH1rRFjcwbYEXFxCFnlk3bzfXveuifNqXVsJ3p5ZyB3wvjsNGzpk
6qseLf4/uNjf73L6GS5wxRWZPlbYJdQrVCX9pQIOvI2ZhGLjTuzIO3OYaDZsDcWi
iVunYWPMnmLA3GiUxP5m7WyLJHumys6mFF3+HURgBk/0UHnBf9zx4luq16BNQ4pd
iIyErU9sRFvRnb0OBBl6wehNIUa7YqsEWYT28JGEdzBMA0w6ZZ4V+AGIymktlPqG
yMxfro76bA4KzOTEOkJUlQ/yeLBjttWeUFq92gDlj+90i4wuaIW3g/dHNgLzXyXS
eRhe8MaAOALUr5K5sAQA5tMKGgoZ9Ya6CGNEOt0BW71cHgVu8MxbFoe14WDywMav
/4RstedV8eJxSdcW+EZ9986wyTSSFTSkMpeCsWzcSD1RAHGVWH52AamTZhQnIH92
m0EeHQJ5+WFs/MRriSEOBCFIyYub4HUAa1YS32SbsS4sMqs8z0D8ZhbaNG9Gk65F
sG5idh7KKfmSrSogK0WU0y37fdEMTOvjgOkwXTVXf+4HfdIOAAvUIepysdO/qI+c
7iUBLMToQmWL84cosQtCQDyrmxIBvwmWW7iwiGIJio1rEJmfx6xbEtLOqDyMeOKt
OWLzcoxtmLa+dYDl7/+QgAjhaENjqFTanrNYDfQlFgxOgIyFZL3AbzkkMkVMUYno
28zQPlnKPf0aKDBWz6cS62TqJmfSGYXM6EwSHVSf6Hlwz1cyr82vhyjdcLJQQ67+
xDtQltFfo+UvrkF/KmrUDp7VtUspLJTIz3ANlyRaY51HW9E68Pl7f4HE6yBZhMg6
qHRlxX0HCq6SCscjOHKGEpbZsSlaquWcbCuvaejtr5FVwrZAZDjs5MJPA2BtURaq
mSVZowIqKd5ab1cRimffztimR/21fR/O1QVEso1EeZTI2hMIc9IKHcp8MvmT+t7d
UGNtaBf5sfHkCqcsmDKqwIJl0YlQFP8Gzvr+v/zkpSpZ5KZlT8aYd+mf2qjID6m1
EeisGp2kELwcDza/kYZFgsTogonz2ybDtJoGg1nA5Z5H+exFUsCbYLF/+y+FhcNw
dqd6Mw5a69nL8XKMdPWAZrZnzhPlL3Zj8PDJ3zRkT/a5GB0EyCTcClQeNVmemsPG
xsP0Rp5jz8s2+N0dS8JxmvcMTSFqJTh7V1BxBjp2qyVdL96b7fRGYmrZpYnkOs83
YoQG8BRG7vfH1BfOcwfImKzz3vK3guNgLputzHzuOY24AzTus9zGtV/5RD4f4RAw
SIreLRo58oAtNhoyoAAnzzVg9kpjPPPMTOtJT5RZr0yrZPIWiHiFC+gmmshoxnhA
0nba5Dt4WXiATnc/IuauF78vurM8A3dA/nbxZztrDg3sclzfNSNMHtsD4v8DfGWJ
DmVcXwU6Pnz/og1UWP3Bw0VIyph4DTQT4mJdrqAazRBCZDL5WPzMxQkgHHezkVAm
hqc6+DYwrOm0fuqso+rNQjmRRomc5WOEwllaQQrIR6pKM2zFcUXW4QtB8+DFkW+K
/mZ0NyRihriepoze7scD6Wx7R/SZGmSuPCPcLShazptUA+b6zXDznq2ijk71mJi1
ktcJsod2VomSq2QmP+mjMGD81Tbkf9c7xZcUmofDZSPAod/cdNiJ8EL3W1PJIeX8
EO5zIbqtYK/tUb3LyBaeDaxQT6Gq72RSSf5oesSo4QeV+4/oOBZLPDZHeWbUwxoa
qS5Ixz7AUIhh6PFi/WeFrk2RInBLDHcxyMdEivRCc8uuATQ8zpdDSTyxZY5CUb34
o7oEjtOIuMXtBz6J+l/4rbmHmacj9vyMCbD9JfCRuVIsZ/1tyOp5wb7fHksZJsGV
leUOEwU+nHJPapGH/rYZ4KWPyXvEVGNtfXmIrZXaE6eXf0YM9kfGGBB7i16EIUOm
b2lc/AJbet+1l7ykcDc33EFc37q+MSFsTIAPlazDLUOkbKIUkmEZn0Z1K4VaYXvQ
Bpp9NlviqqXOnqBOlLxOFDPmQ2NaoBtSxeG2sHQaCiDjm4DpUW+le2XzfYGJVmgS
9u1Yjj2uremxGNUfMxnFPF/wNYe+fTOaWn7mnQbHccSNsn591bRCo9H24juY6dB5
p1ncIqdv+vaf7+3Ci8hN0nhWdyN+OcsS8fXTIgOR3tq3RSfISUG20yalUf77xyum
R7/Y3qg0pK1zvRwDl/PhsIcAD7ZufzvvrB79QtZrhQcmhcQTQYOaNEyDUmgJbIHu
JjnHo7y2K/31WzU4qv6CzXCQVh+qqG7DrPdWh44Ha8I4+w8u4Vu2J6hNbm8z1gQy
8CCStk2cFpiCa48ZxGS0ViWRa1AMXrg7NOwDd9XCheD0S+UEtlwOllomGeCWPMML
WXicIKsNc+xgn6MadL9s6DGTdGWg4OKLCHzPSpV5dbNJpfQ8WmqrQRU34iQxsAXg
fOm2H/lxmiPZGQvdalHhjPV+7/aIewbBOr4BrPb3S/4iQIhnwgNw3dZu2Z1DYufR
fpjvVHCmUOMkGNZczBK+RmV7Qx4SSXJ04AGtp36lB3s4zbuk8ZNQrx8YoGhwyJYJ
l77b8ZDgFS526hIqu8qxlNWAWKg4AJXlFrcDi7qxffmz2perLr5oxhoYxCGreSWt
om5GWbeH2qQq8VOlvS8N18S3BuFAIe4GyRw5qmp5Ur5YNR+UrtEdbE16uO7ScUir
9XinW25mcmhwoHra/YLe93SR0smeiY3TorvLf5V/VTIxa9TZQp5+jGwsePTFfXD3
59ZY/fmXDM6b5a04KHFmM1KX8dKJcAPHBsnMsUc4G9FXhSdu3LgxNqRSyMfFq9ob
O8hfg+XuTdb+B26/V1tAEz3b7banWf8AWtCvs3tbGxtPVzsMmSclIIM+2atBWABF
tFfPtpqxgasn4kzgQUXvPoDOpFhS3wGHB+s9SuPOKcLKES/1OiZqi/LBLR/vPUXP
GvU+ZJOS0VyFkr041LbYizl68glq51ZEXNU98Y0UmJ9tRHblmKXYIib5lxGUUrs+
GB8g/moodAuDgtrM/l/ZXJUUYP/XGWbC6Ds2fOTKMui3wj0iRkmPJoqjcWwWTC5T
BBZSUTIMp1zRNxM+p5i7qkD3xHy1TlMgbRdEJ3IczsiFXKbAQ1ftHOHQlILGw1CS
g00VdWqK3pd/7bXTyUTkXwcLfeNM4/SbSJBsu+AKs4fxMAvsDc1bT03wh6bXGJ5f
EGN9YFNOo9sk1lVQqeC4mqwBdK41vHsnf8DpjSuBQr6dMgFFm6y0RIS3K2ZECE9n
KJQB+vA+bS5G3S8+ozEuV7YejKSdoTH7rHIPSBvmbZs19yFXJoti9ntplalx/f8J
/zsxBGVgw7/YxdZf7dwHKE2Fwx1iw7pA0TXlMznIrXqRRiteYELMfVldpvmNDHnM
wshdOVxSnC2hHjxhGFN/+SUu0EuFOg0pWjD5RsW+/3Wx+J71TPlvKhutCTro/mmi
8ViBGIJej9wIIYUsptlAO2oLvtlJiC+GoBIVmdr3Ylc2S/v4JEZJdwLc1wDErEkX
+ccKVFzswpGB9vtziEQm7BMKblI/nycSCzH17XeaKchEd5qpvLC++Mf76Zz3ESa8
QJuTjoD0wOG+NaGy/E4EFls31dsatgjxWSngdPCX5D73V/yy6elfbOIph9fx5TUw
l6NQyRiTRlgRF1xuMKwFOth+MR0uJwjlNF3YNMt+CXNeinUOiv7EQbudb+p1Lo16
rCT31KQZpEwHxiAYIPu85BdUArs49dOBR6j7OvtzS+oP6qJSzc2rk7y5nVrO2H4b
zHPQknpi62uH9P5Z/D+WyGrpq2OdIPbjmt/HZRK6bASwlTryjc9CtXblfEMBAW3A
f7rHGVV+Z6OZgzL/KJ9oPPniYa9WEp5f/06BkSxu533URsk4lsVgOr234LSaVnlr
p770oZfoc9Ru5L/t9hJckLERU5EZCcGWGWOYJRDOwYxoN8HmboDXv1mmIcag0fkK
2ocgOPbDyOumJYDw2s2KGqPyzpudURGiHdqVG5DeZxsrmvE/mRZYOssU05KxUZOI
24P5fyYP0R0XQ0tIlcDXJnTLlRS0lhV2GdJISc+FdpR7sRlTbzIkI5uFLsm4Q+r9
wY2GD5WifHbSk6ET7U/OOXRcdcMCprSJQ8dnyY4TCmUaCaQXppUqaftwKVyVSzPc
CftKdarBGu44xxJ2O8r/sZyh8OsnhHSPhF79HWjGMmGm9Rj9adASfdleth5XpCzE
NBzjj2dIbXcS/C/j2Mz2Ume1KnU9hlbl3HYwD075xbZT89I+pNAWSID7BCtrjU7H
PgIK7B4SK2DnMS0ujPUcHcnD9VRYQPdQWvyHVnwI8AlgAOKYpLhrnk+DKxwDAxBR
y1eP625KIWEjkNFyIbBhnPGhMbfAw3X+aUQ9gxZvFcfI2VM5GYZcaO9e6ju2I7ko
87BhHokyOYxpFYT2VlTOve2OAbQG9g2hliFa6qyHfGnF8WOcdSaZHBCuBKhn+/zD
+b/THMlAsIfQ33tYwRZ9LFD4HGL2Ys7QJ50HeqeITnXdq6QOmHjj+e4LHVqJoHv8
/6WJULfn4B0UyLd+PeDHO+vx4XwtqkiGUE+eB1nI4qho4mKizztYG4VyuJ9OD87Q
8db8pyX4oZnv7qy2mKUozB21pWgUrZnQQmZDUrEKy7yRQ6iQYa9Y/Z8QdM0b3JW6
H0GQCJn9lDtfiN1fOIaQLZDUieEt43u510QipfCclE3NaejZ6shp1sCYlWmeCON0
7xjIEMoUcrK+8PkqJSjVkafcAPt1GW8RJXZZXjkR9FbOoJWoAUCkPELZ07NJtbxc
zj3qsMrSTb5Q13VzJ8heAXi+2D3nQJMTYpqaCZtUAudxoI/h9WdKEKLrGFCAQBaz
RuU6A9xr+V/xj5mFe82FChG50F93tTBlVdYd9tkcnlMGg0kpT4xDykG5x9xvgrIS
Qwbb8OFAFI/04WZ+GVBTV8IeGzAGjhVQP5Mk+FGiG/igllzauUy3jhhsArePqKr5
NqdnNz3LeH2DixGjcMMV7O+F+OZ0MF0exqrHK3Rl2bnIbFKCznEqAEO9LlXf1f7e
W7IpBDPo+9+IH2EaglNAgQr6wL6+rUgUiT3hV7DZrpCSiTo7d0vbzaGvBRTJLlL1
kBZl72MtVSujYcpMPbEHmUEN3LOSCbel0NjsynzW0bjiPCqU8Hd98iy6qOTZYFEZ
YTCJfe5NZggMi8+5Wjm73LByciKpEm+MzhfJYGg/Q03lsuWLL1GoECYLLcIsigg3
jUZvzBB9YVBRQCsBvmq/x6O4Kjz51qzW1f7/KBpnNEyoEnzSh1ePu/zbGH+bp2ao
r9ePPgMCjz3ve8bdyPcUW9iimDeZeS9oBzH9/2i3PiFtniU62htExVu4tjc+IdDT
v9pyRzyXOzyvuE0fKESVz6sQyVBpGDveUYZrDECeA9/oNpTw0LDbSVoR5x7FyoTv
QzW2xPUpy+nv0LcAYcmfUjaXZu0ikeHtTCfa5JLrJsR1RkrYxF/G7YjVplB7c0nH
s9fw+LU2f2D1y8WfmK3mm9oRY5vkMT7j5VtZxE7T4GAMnpEuSYrULJ5agGInZvn0
x2a7/CJJ8UI6MbHqmjZmrnma4rqBw0KcApvXyT70xbIuSMnGnqsg2l4/Myi4dMZc
jJk7RxyOzvCbdb17GoE5RYVgik/u6ZJepYxHUy59QXYwM/dd3TE2PKM1lfNENbX0
R/Dn9sUfHm3yXZBMXZmm4GOzyDEVbsnA9vsISWN0z1rcgMkEx2oLSEvwTU4ONEB3
KR76qdx2wB7oIZHHPUT40cHLJNTccPr3m58banULLFktTCvu4GACChzNw3xKwiWq
BBrQvJlrsHMy/5M/MmduNm3ivhL98VXpwzT00+MSRu7/O0UAZSu5fhmzgTIXOpuu
f/0YFNssQnx3BGms3RvnDtoo1f1yO6HAbZymWfsFuCT7H7vN2alNVXeGkRq6jnco
X191Tr7FT5QgKFOSIqPBxlXS/GA9cgsCyLbK5RQQzqnZg0DlJ3zumIwnj2CWOCXn
7RPQo/R2rIJUEPX3uoF80d6byOfR9f65SZp0Wd7DMX3Z8sKRp6F60SJ/+cnNIdbY
eJIOiPhAkek0MK6BcT2IajhSUOUB3CHnbQnuU8CrUVrqZ4Cr8ifB/P/U8nlY6fxc
8QHBXUuLFwH3MQxeKSRop8J7La9biL3ygU+j5uwJCAL6hHnjYv9XS7qqo2s+ZKUf
QbtB+kQEv9vzspQjzF+cSDraOz/GHPbnEllqBXIKeHsMJbx9eZoiQkvoTjzw94XU
7a526pw7N3P8lXdp9IhQlYetjYjX/FOEhxS154BOUWk3yfHakwY43GqIyr9Xsf/8
a+sCqxuTH3QPJ9PpepnHOaM/71tqx3/5eo7RK3Q6h5QAIcyNaqknlLMtvKyeetE2
alNSOnCz+zBhNSYho7AQdkQxXt+kj0Kfnp3HZU+lRBYpP7Y6aUohbl87k9Ua3/Cl
g9bkb0E09B32TPlwK4zgSNQ7XUF1/WX/OW9lHfZM78zexk20pRNfAEU7fjDUDeTr
eRo7Al/mybtrrac7SHtqj43ZXTjp4/vcQIvzNBci2G72CbvZ2K16T/6mCAWtQS+H
0PlTJ7Is0QEsI/vz8mI6HDtUmt98odmLS+dcjwbVQkg6zi+0jd8koZ+/VAMBMwrM
JJN4mM/s5K+go+UuXA/nK7OSYtftbpt1qM7QBnb85P9vHQQoxGkqrpHq/P5po6l4
jl0A3vVyg2wMX+SBcy/2ZUIHqxTaIueEmVl2AYWD3m37lnGUZQRXGO3fH51knP7c
VIvnbJk9SETq56QRj80nEP0kKP6Eze9tOBJ39AgfjC09CrtY+WoNKcAdIDUO2IiT
ZtFr7fPEXoKE4wiqYXj1BQM8i9EIXnRZt3r35xN+EqIoiIb9nP2sC9q8wsbaEUxP
7l4ZTthqfK/xVsU3uNkR3JukSTh+wN/lp5+ma/cNTEWj0CsaeuEWdNtmFYtpVQnj
4MXnkgjJOvHwbYvD8hOcpur0Fu+AsqIzcMq1TYLqY1T8kmDNq4cu+kpviZ08vqKp
eOz4YhFhE9usrDNyly5EtIDeErgxkrN1K3W1EkWXt3kDS6yOn22TvWL2j48Ma6Cq
jH8L0f0mTwLr1aYCQikBEpfMzqb0AwdEaIrKx1d0DoDN7+eH6zY6YHIKJ13YFtBG
p9xCbpoSDwkc4tVTA35Y842csqjDQcUaraZqy6TXflquN9byhi1bsfaLXVCxwXCp
cgMT2IKU4822ekhCSiJQ2hCMv45I6EtJqVy1vzz5b7JT0stusBttNVjV6s3/tgpe
22lx9ryr+ahO9CBFko4dKqqKeeuBd7jOK7CRmhTEO4DanBDbX5B+4qbcTHRsIhbl
ANBPOOUCiz6rbLN9UDzn70epIQLcYOwu2wO5rz7Dr1ASTrEqzzCRODt4nWKc30GG
ex41seuqVYx4dy6iDiV2d8/Zk6EIDSmfVuuJUXik2B2pcUYl5e38+F3QQrckeSTN
RAB2Egtp/UbacwY2IWVpI0suMtr46RHnai6HinbFiysPS/HRR8QeNBTUl/A7xoDQ
4x+cCWvGdSuHFSTvyW/q1VxcF0CI6cXW4NSep287MOdlzeFGtSwq+WrE/IiJRj9s
QqMwFUxkRXS/56akTzojpG/PrKHgsXaHPKBfaRDJk42vrIlA9Tkj1ELwi8uFlzyR
iIliBNY83VBcKJUIZVVRB3chZiUNxd6btdc4IUrAh76XyFQNye2kxmurFii6m9fp
uMGlM8+fh1c4/F/UWJTQIoWo8gWQWF+NxVaLvFc+rGOAiYNWnKhl2B8+JqdLt35s
pvPA0+k29FSUYnEYexOb1d++u8k9E+L5s08AfmwNGUtD8WnGqfawX+4Te8piwMsO
SpuSOqd1nFhiT8aSvR0DwVHJYZxH7CDtv/h2kXRTzTd+e+9vOT6usCrELjv6oXbS
M70JGNviVaN5yV5g1x0e8uOOyNlhciKJr3IizTFB1oof6aYhiH2Nm7jwGCO5R4j4
qeZlo9FcuCXOmtQ3LuVTKP/dBfQqEnvmxnUvpu5g+rPalQNc59UKMZYZ6rpfZYZN
QeXNGSzN1xzFXqhmk6guydln8hb9JV8d/UB5WK33f1LToyfdRA9yjK++gACuTaM8
K68Dz8f+wB/174RijoiXzxz8CZCNymO0Gyn9O076aMxwvVitFmDho1JROtzCGnxL
x7HpsEKobSq778QBK+ak7TMG9z/S9j8LrTbeaZi3giEYDMivjrEL4n68EdHnPMpX
ycNRViSGaVjZWNo19SHaWlgVIFZ0KHF+eY+w/yDkPE6lkRifTq0/0W4Y7zzJdreh
8gy0oTqbPXEYBsDZSrQ20ZWrrGe2INO7+3S8VnmLxYf1MHkbavYH+ADu5kq3eRJX
u6/vpyBDx0NtA9t8HeJev9zRGCcvWMJ4zlFARiqsllsImOlAZjDpdsq/SaJO6MPX
kmyZYnWiMSAUJe8ZUzeSj7uUvVUe9IgV6kN4XxA2BW68lP/4RXKfxbFva04/+5J+
PdO9UdcSrgg+sUdwjz47Z39jX9RKccHlrJVtlN233hElUsJrccd1rRAivgY58VEp
i6+SBz3EBzxF/4DHwpokvPs6UwFVohvbAH3nCFZIzhzD1tD9y7RcCID9Ns+FdfIt
//As4cne2JoTGQIGUK7Mxn1FxfrtCRTkX/AzqAklXHDQsEAHj1+kvTSDbwR+2ZJK
hy0Gp1K6qSE+4CcVtIiggSC3TCyfbnMN2vYmEtbRCy63BZLAKCaEpwUZ6APbf72R
qWAV1+4TDaVy/pnKvNoqVu4djE4uGDlhDmY/jDd3A85APXlrtG+Z8BD5H6KJSK12
veOUHagAaIyC281d7uRcycbtSfbSCrbugd/eOhf1Gxr3xQ8vpiQk3wygdTBFmaK5
wh1rzOjcyN72bVkijQhLQvcIutCT0Hec3/IDEvT3/ehcXz+4vPoRvjP8Z3SOcRyQ
FltM8gBtbHpwGXWRw2+reThsfSHlzpInt0E5RTYWM1vwkaXZaBLZ6ur7cRg66pUO
Gl9ViMWj10eWIbNpOhEWLU8U0YsQvjxTt8mumL356FPEpkcJ9NwbpW5Z9tR11vQB
JfNzUM4EfyIZclq9E3LQFM5ig/vAdGVrgg/QrPeRJlQ+lxjOxWxxatjSOZhPdCwA
hAP9B2wPxLwfrkOo6dc1DHgyETYvGD0Nvwa/TqjkRsBmd0gblNftbtTwzYouVjCg
/wfvWTxHPx/l00YAp8vOnIFavqpVxdlimJqCgrSAaoALmXR2qgarlsEmBYPQLCSQ
0xRJyEqH/9aVRBHnSTjMZuHvHGcBupJOKgAslpyIm4ooI/SNiQsoDGChl75Cc1Yk
2kjqR88kfIlqkG7Enazzkr2lUBhudRTbsGSdSypa1jTe1YrbFPZxnChMfesRX5cN
/c21f0TbSsignwKdpR6oce6mVzywl+aEGOhZ/kkLa9gHpzn/8mbZU34ES0FQVcJQ
aamj2mXl3C877aIk9vSF6oS+PE5u5HH+L46ywUxfTrhMN7tfZlfi45vemp5Vy89W
NIskMH84qnayiVNSIc7RlplkhQKG2IO3NFbLOtFWOrpoBNgLyioSXGwxepTnwXCx
wIE7QCBFAjid2udF+ijo63h0e9jvni2JFME5YuOGhyThRQVLA2irxQqGXp5OqxDS
7sauT4bzz7TL6UoMJC8biMH570ble/U3fH8BrPqCBDdaMRR4t4KIK0z7zVffz3lY
n1LPyyP03ZXNPQq5Op5huj6gqJeq5I5a93sZVcyM3lbmb0fnXDteOqfdXAQgl3wy
jfjGpUTKqVeIvQXultZ90C0SdV96F5d3UpLH+t32L/8MCP+RnyyNN3H4t+KaFdZS
P6csjhN+vg4a1EGZK8wj9LonKcJEqxO+BeuD0SuIJ30Mxkzin0OUZEGmTITmkLR8
9roGuFtQhuTHwaq9+cHQNcsz3xCt/BH7/Ngo/LZqO4b2bVlqCXYmUNYAUdwJtxvs
I3hpIkyIDPuE992y2HHAr3RnGNmlTWKOtGgBMQOF2Y0HPKGV5IakrdfOdrNUmp6N
hSbbIO6AQ+Vp2baka7Yn0/RzbWzqrTXQsShHikp/o3HuPjhb7yma/HquJM/q0x1/
Qi9OnejO2GOMwVJqajZdUGNaUjXO3v/R3BHAjZPd6i9VrEG5T92Kllj9h+x/FlQj
AS07cizHL9ieGHZclujpZERx/hE6qOZu+l//U4Npv+P/1FD2Xac5eRqVxD1EkvEu
SZezyySGZ+4yIkzVPmLPaMXeTToJlZ+YmmKzr/GcrrYdGZtZNVP44kMUugwhj0s+
uGlityyjkCTBg9XCWSgajvWNmQPDf+anEU8nv7fx1nRiKd9Xb09+6pYPTW2x3HRc
pDAc4A3WHozGAMxvJg73shNVGU7wbErtHc803TpTRrF8OwIIqvAs0P8LIm0ypIx4
NtwNKjVOuMAuLTQyAWpYwtVekfPG5FyLRSnxkxHSH8zI9qN5YtFcp6w5Or7bNX47
osIi0Np8N8CUu6BOw7wHqAQ3nIembu0/u4BS4R+VuanDoonjHeMgzbbomRCsRaCy
/un9ZdPgaZcwdeSZnUf66TLxt8C93Uiw2UYzLptw2AW9JXlFBeAuzxFNUK5iXkRz
cqSd1jNSVvMP8L1duVgnnNp/HqMGLfl8Bmd2DAbsiDwbMHqqhKsLkrMyDnfa6c3d
iZ4nne8UMsEk5lJRryoVcjdwilGKnO8O1nDBQah753qZvB6ZMfK8xCqeqdD72Ige
1YwoJg6+1Sxmimu728D93v8ZJVKG3V4hcXC1dQZ2oDwLP6PL3sbJlEqxQquvdpMO
Udz/hyyE6PQuu1VrUTtd+WqKHywuZMuf7JoD5IW9kkwN/6QxAjkuLc+AJF5vi/0m
xmCpdYB4lpsWVXjThGS+zP5D4n7tUANRLRUusTlJAn4YOxEVUlAuKPMOA7J0BFT+
Kw++fLcDYeymReysVICTNKcwauBJKrEi7+keqK1uAE2C2Ls3Ceo/PVEhf+390cKY
zkmpZwFTrLJI46DB1J+AynGtF92ymmbM5hu2ur3c+SMn2PSJ9h6nX1FPm5mU+SmG
CjUEhUzSW2DDoO0IMgvNC3rK28H3BfVWqkL5DA4MRuEtwqY07GOz4qAYsGFQ9kGn
aiO5SJfCL7fH5B9nRaMOsGBIHXc8G7sSUEokGjuWdL9uMFm6eMMRRrzsOonlas1W
ktfM1xJuJk43teBycI/os1m9j6y1o92NBnnqa6P2OPel7d6bwjqkII1b2OnhQeMG
7H75zWf3y0AIqsWsNfw4YJUtYMumHVd1khNDIOiLWKkhaWUA+DfBzU1K+ep02G9r
6mHguz21pagLyggyC31nj3gz7uXCqM3l/IG0Gh+C4BbfkcCmlxNiMqk6nHTPqZPp
FzbQOkSjRfgtsVkrm2UYqtOwKvLYnI0TH7Ib6/YoCPdCbyPSQqTD3Crf1WyDxJ12
w4Uw0sUa5opw6mEdDlQIxofNQ75n/1/gGj7xiD8UGv17BqBHhCFc7fsZl0UfxDfb
unDi6Lzfu5RtqxSGrS66SSO17g4wZknGys7iXrjlnW0GmmHE3r9EXG1MZFEXRWG9
MhuIn1y6105eAwZ1T9y3MEnPV5vVsiLSlhQ7rzZcoYSDsadVnu0U++sYHoXS6znR
Q9NBta267nS7MTIdxIeGj7FObeQbO3yTX16RlY+0onEm56YU3YQVleKE0Y7UmURq
9HSsf4+epBqEE75wTC6NAwiE8EjxyZ7211FZatAzL+KUechBspk+A01aW25sm44V
lGZUXmkOBytZ8PTbOM85hkUpqxHvdb7bBJF0oVS7VxUOHXVD6MWgRqA2mxoFhXze
a8gtJALLXMZliTacKTVaM4b56LY6ZodTabXPUI00iZblSvTzoH2j/yn63ghskzu8
fJ0WCS/q9U/4wTf+zMSU3DJbFKv5h0Ex/yyRdv0tuCNdejH6qW8JORK8Mkdqle2x
EgZ8EqhoE0RzR5aqf/iAfrcuqgr1aMyZFpaDOFcZGGCx4gYrOztuEZioECxM5TRK
GOnrSSkS8LpgPtrwwh7GRGWMoxEcNM+H9hC6cb4yuWCgdQMrQzryCzGvufDJm4w3
WZZA06ZXGvy49TNsrMZ9dGWOVPMiFVzIt/xKUcd3b6nS2bXe4d0b6DOEUSTvSZzL
5wSZc479ELvDww9TJgd4fJX7pgP3LnYet7Wk4KgyO41eunM2x4yqUJfAWR9INZF1
k7CvCCKSzUMYP7gV75wGTHs2TTcNlzTPt1akJvBCRXPot23v3X0lLLsgkydwJAIZ
m4fllPlVpfAN9HcjnZ2vlVB+v1lCEBUga199olFqbb5tbSN+NNxENmtuOSTYqQg8
OHvD629v7JaZNsta/oZM17b8Rqw47oi8pQSdMinYhWo9BdTCIkcVUeqXtV7YtLD3
4G28MsWhA+wTADNpX6O3MqS6eS3qJG9iq+rWkTwIkGaRa7RdpjDyFKvFCrghe2Ge
qk35AOlb+KKxiIKtBjPIDNuGbL+YGi5ZPn8yiWy9OBo86dfE0UOh8jxocoHKxYkp
1/2TstUBFrbCmhRUrfiUqeesbUVbfO0zEoTT2kWdXMqfYeGh8c5lGSO6eVs/29Al
LY4vegXtBm99nMPeQY9/Rq0uhetXM/7AkeT7YdHwSExPLkOA4MOOooeYhF7BeRTK
D37PSN3Ztu+oLx/OMRhAFCPUP4SKQITsjZSfzNbFfj5P50g2f8pdEfE0ngOyQKWB
mPnplBpa5ich+GoQYHTz8rR5ZGsqaoofaqQc4veTMSpQYjNfSG2q+mo/bk2IFziY
ZoyKrnC4sVnubsLhJ3pcDKx31LG+AzD09+Axt6ea2VRgSV1tMKtUf4fttuD1uiGd
Nr0Xva/f2GgeA/v2+eu4BsR2WpykP+O7UuPcHL7qZFBbAwA+j3DAiiU5E3VjMBLe
WuEjVJwCpNKfaxUmQ9Hpdg+CBPWjQ2jPhu5GkuLtz6yX4i5Q3BbbSu703Q9IeJeO
W2E1MYlbRyRtIJGqE3BxiaeRZ4U8jZU9Cz2Kcu6w+JHXJuMA730deHUpogvN9dlA
Dih43F+/X6vFQL/Rx9G+casI4VoD6ZQmiAVjGfNWS0AvNJ337SI8dKeBBw5ZPv8Z
U8GeHl964O2Rgka7+4ulVuG6iSzO7Oo4xuraL1h1PO0OQiA/VF9Ld9AR2beyMpom
TO+7tnhJLuazYR+VBYSdYqkk2TY6g2N1D68e7DPzwHuyEB1NC/kALk2omlnNuuyc
kQDYI5CYiZyq60CflOe/j5rzsUwJBZYlTB1WESGQI7s5ZLc8Ojs4c9ARmNuPhz27
NR3ZIUZ/72IGVreYDprNJKY+IBNkfP5mcq2ktSMDi1HlRaVWDa/+WOXsiId11LBe
aCSeItIVGC+r0HldDRXQNDFz78sjFoC5CsNtxu5SXR2glfV8fuasEJdDoa758E3Y
SxqOeoHc4I5ErdlDi3pIGhI+31WHSMFRlHNZ1aq+TP+ZnoCNU0e7UV38YwlcjpQ7
IYLjFJW9BSctku3QbE4NeKkgIbd9+pdYhW5jMkczQ9VJwyJzg9OcjgzX1N2LaTzX
1Inc8794QlRkG44P1qSelfVBgpG38MPB0mklDDC3cHeITJY6vZpsxGXgt93id7OD
xGnpVR5ZC5/2CNiZnFW7SVWAe6GS8AuKePuYvsmiR3PRH3gXJ4ZswSydLrDjZzGB
TvG0KDhcJ2z4cKcL/vI1fDFNWYQQwSuhW8bwTQLO+g7Q0hKin5JgkRO8kvX/6eY6
BG5vMYEgz7fBHH7/oua7lFDIq0UW666Hv3CbWd2IO8AHtZn+FoPEpzqE4VWKQ++q
rtXIp6DhaI84/WnpqeUUK8K8ixXK94HyFVSwqzrxpDn1PPptUDiSDoyqW+OXFEcj
302VKykeVvxh8LRRhvd/Iymo7FiUVp0d+eLCY1YNS7ZBHqY7QUhAje/Vq2HlyCB8
UjqIdSluwvARMpVQ+Ri0LpdvstBhpf2B/v7K31hil5jbG5ZDpkhWkZRN2JcregSj
akUBHJsBVkWSd33sYiZFjP60FWa2+00b9bx3UH4pj2Yn+HK/HQpUATEC8zWKmDWw
BPAd+e6s4jXz+PBxJzApnZ2AM3ZqBNBe82D/BcuZ7xyiVKrsOYyDbQwu8IjPuMuB
KJyMVTEAygOQtomnLNZeb6TgQAWe7JyuUg90WH5f8HN9xGdj3b/5/I8RxbexkRIJ
vcYMYd43i+R4oP4AE3pBfxQOP1FS1/lK5snFyPR85oh57I2hffv1U1eX3BbxqaZC
JyFdF+dX5J6WcKtUTzBcrg+lZdRwqXX7PTkaPEss6LZFlxMtggYiytYq8dnQ2hgt
92k8XjK6qMvcrp5AkwwaNHe+SkutvjxAZWKvLl10peNQHNqFaPTweK9JWXewIISf
mmn7VN+2YQ5w/BFSZKT6ue8XuL8gQZZrZX2TyJBxdwkScenwa4YnrnPziU2vowbE
mYSaLibo3RrmquaA3X8RgTpLZEU0DV2LrHAxgEQ7y6zHueRqTq7b2IVWVLpcF2w4
Pd2ewXPiFykn4+Mse71/8w/WV+S2Vgi7SMB0jWOvy1WiQd7MxLZIZQHc/EWkXHiS
xuRSBtsYUZKax9OpgiWW/vM05nLNMpfx/CQz5+sLJBDibXf+8SjVmC3YciX/mbW3
Khd+S52jKgb+Enmsw/ExYX3qC0KsXeX4jXPjZ8i+aE3hrU2TvO0TToyhTqf5eaum
yO74Lo5u6X28hSdPLDIEsHubX85AnUD/amLMJ5cjCa9ND0XU+RjyYNAxQCffIhlZ
SK/Y9Wr0nZdQqniZa809Hxrsa5XiMQfVIwZ/VHU9EakfyqGlQIkTfugSO4lJ6Rzg
BffMVz/oBKufdIjSJ7x+V4s4ZYskoZYVDEs7jbsxT+dxpZU2kfdptOuhHrcUs7Cd
v6wjgS8C7b/4G5KVuI0VStuKQtDmKRprTuTonkgdUQ1Alz45KULXaSz1VCqXXWAb
SCRiZQUy8ZcS73PoccyEmEo2lHM8KX9EgzY5D1ddLeOo4Sk+EmU86SLrhKOZCqw1
lCDRzHJLFdI+xltO/imbIDI4vLoINJVgisvs9XBQgWN0WAf2+bLPiStGSfOis2Yo
jwBKIVd6PDsOhHJdgQzjg63dYlytyCAqk+GP/MWzfjmbqdTsDAFcDqAWS0VcHDXk
63aMhaagBYTIrDDtjYtukRG37+f6xgHGvTmW9rUZ2brHBl+c92uUdKN0h2HLEluK
0ovpbRrqaSw48YzkjiW4SZs+Y0UUwExRcNE6tIV54wn2PKlo7Y/JahHm9msIvBAB
8NQenNo7rI1c2/9Dk2D7t3hyWk/bZ4Iz1WJVrnisJ8bDThzmjN5+ZH2xqJ5DSB9K
X/eE4oRmCV86I3Tkz6Jy+KClEClmhnquQVLgyUEFV0i9Nom7KZZ1h9n0abf0vHFW
qHWxiN7rWyEjGbeoafunYTqTpdUNJgYIQCE8gHFAQNLSGYXjVKUegoL0Rbp+z1YJ
ygQ7s4JyK7bLuptf+LTSyiCz8GdaR2Ln0b046y7Hg0oIylxNYNNtsKwMZOjV4/RA
LWkxi43ewUJxRev9V7vwCK3THC/p5/zAqfVBNBizJYRVPIgWiDd4I3pSKavg4InY
2TMZkJrvdpaNeS7OgGoNzluqEhmgkLhZVSqcYD7BqMb2H4r3/4eSezBUtfLtNjyX
ChYocX4wV1veMvcF5twQVzJW2s5kETcJG38ir9Vb7hQINDkfxRbgYl5HvPZcIAQ2
rgYjEsFnNB/dTfqeebw0otcT/mziRDnp02flHq6tBLWCdD+Z4OE/27/zpaBTHzKd
MOnp2I0qQu+Cx8+aXA/DYcJ9RM4+JJCO+i+NPvohjkMEavNGG5Zrlk+k32Jz1se6
sQbXEa3vKrU9ojaGnRr6Kq4Bx01hC2A5hdAO+V6JweikP0k7/alysBmBvcAhLVal
xpp6PZZHFdytpIIF8z2EeY+cBQvWgcz8YJ0U5IEq/XH1Yuy7Eez5ZZLqWbKts0vh
8qv/6cchRSSUL8br1PWqIAmLv8xAeRzK4mS0iOp1sG2qJ9B0Cd4gWCRYFAYfPjcE
RaqOLqf6Ez0JYu9pfGqpoO42eO5Mx2USyPDmEgz8aZ4YIQXtUKSPKCInI3J8xn9r
OB/EKckI1YDS9M0JXt22izh80+o+YypmOo6jaTHGrSMFppy26zzYqZvYWBEmj+QL
5M8GF01Iz1J1j5Kq4H1PvGWBaxO3iZ5Vl1D0mvPJbhfhZbVlv2/uDOi0tDPAd2ab
tiaxpwYc9sbnuLpTKBPUEXMvZRDG96NfGvWMYtYUcV+Cpfxr9LvNSXVhfRyszxYw
bcKQw3SgJnkn1z2wy9VpHPCpdmQcbUOThgJQQ1HiaUQmZRI/SThot0vcMZGGWHJb
xMbCrZBmnoIJjDDhlwKCN0OHhMloHKhP8JAvor4xr6P5usBNcdxTji5khHeXlEun
aTiAvrrZ7qZ35DrjShbYi2irgIf/CcUIkukK6sCBZdxZ2CbmHadXArBZXGYhPJt3
dkEh1EL8VZFfUyBepWHYC7TJso5kIE2lIaq5seVzNw64UgR1RyJnekG0eZ7p3BKS
5MJrNyrzwSVxQNdBaeh8308lVMo5g7Rdl6FCaH1XC9If8n3jhHD7a8ZSV+AFWfqd
MeZUTb+52+FfKhACv4P4i4AuM34AW2yNlUg+JuQgB+sbuPTZY1C25MeZEd7KZqel
FeESxQQpaII3ZxYM2BM69JvlO9rGO64ah+B9cYQSaEx/bqIt/X5SzNQTX6I1H0/8
rbITdeRZ+Z3nPwdY2j+AUyTYPQgp0ru/dNC2+9MxFw92ujuRrqVSGlX2bsDsNkJS
0baLG3d0ymBGPnRsWj/pvqAc82Css1/JOqOL/uKyW716Hjlq+QmpcMRtEXagkrrU
CuNK8IseVslGR0P2YNynwQ8ngAN2Fdr8uzv/HJ3OXD8QhuUcM7kSX/qi5G2ak1TY
/zLZBmkbFU5OUOQnAABrutU1qL6Py56GlLABMd7gCuIbqwd7EBpA00kwTUc7cP42
MCFmIC8Aw/OWlPWu+gOBXDfIzrOFDQR/orfC4BVU8pdYykacYB1PwHN2SQRoUmjD
Wjqh1rtBO5DlXIZEoGBCfshoy7iH+2PK6pLvLTxgoPkJCexuOpn+4ahhXlaPRRdM
6xfbwwd3sdyesPQ+wHTJo41QwZV2IO9sBEupwfdPOcVDK/n+P4u/jkIl7zCX/L/R
Xi8/yWNVpwXTztn/p3WR87aSy4EC8D06rnvUoj2X08ID5zXqkx4dhSjB4yEWJMGR
1pcIDoYjqnb5IU62CproLV/9B7jejZwDojXlJFS2d6wrqA55hX2pn/QvMwLDheuQ
uYP+8ydSQjmGiI2XAE+b/x+UQyFKNW2MQgfJV+jkpSK1wWHW3gbAtC7efJkDsYNQ
bamol0C7fUT/1oVxe/zGxTLazevlJvPyc5En8ik0IdI5zh5SVtficZrhEdlEjLYd
JA8GnZGNh1/P+SR2zfVx+8TuMdXcq4EiCXz4V1OjVIUCM4EOoj7FS3+caHj/Ys6J
SBMtuYRKzpZ+mjTeQY6cxsxqYblZMFjV1uOmYZtoMSJsfggfnNoOYsDRPOE2SolH
7ylETWHpYqLsIqnBQek6SIHw56WyKOv1MnM44YgX3hbhBW/UifyiFJTZZyFy7PPf
7j8T/FzHu4V2eoOratGXW0dcjJ298osWZ3DB7qv+fqymzd/5o4bH/6Ddn3jrjOx1
IxRhaF6HfUVb8fG4f4ElkhuorChf7wBRw4SNrK0WEpfRZaKimeJszfDWaaNKTe9X
vkRp+QtoEinfeZkCy2jF3SkiYXL6+18CqcEROflXj1Qi4ufteqIfAD/RGifg966O
ScJJGhBF27iKZnqBqmCaxbmUXHkdOq/N4b1FzmPy1CuSX9hYLoUvk2BWLxDLYvI6
WVPJsu+jVGVHLEQZbLgHjeKtWoeFEaf6+c880ejVoIPY9rpI/PYsxWi2DF/lUnVE
kPxEdWshCqe1bd/M1u0VP3tLwfjTp3hakjG5XxerVeaBY0udM/3iK9++gNvFkwRh
2w3H1JnsXH7QYp7xxGON5lZe6zH4U3yPlZNCUg12kymW/wgBWFjbKV4OezQGb3kl
tLdzKCEytvfEsJMoRcX7gOj8Pyt8pOQjcc9Hq3L4dp8ZYGYUsFqfwUkqeuWcZf+D
vm5WqK2naAzb5sLJSmpAqhnd6HSVE8qjSpbuRIIrF7PKlFki1CwOhWypoZ8WzZi0
hGiXEtrGAry3GTcVHGFtJLaxkKBV2u5owq4GcsyqZJhGXIrdHQnYEFZ86UVwS3Df
QAYGsuvyAunRQLtm4ITpa/KVtEU3uJET635Yf72WiqMbis1AzcmGTw8erB4vbNQ5
RKIw0oebqlu35/ua6MISMFeLvUs6Vw8TMpQ2Qbp3Gssgquk1+T5ayL941T3jEH9R
sSSqjSmUjgTLS2TQ/2lKFC3YiSpxG/w1XnMWbzGwSIJtw7wv5LCxSQWSfCwSRuoz
l97Y3NZLXYp6aLIfdwFPkV4KhGmrHaCneCzK/PNG/YWh61KN+SrQ3lvl51oH95il
I1R10ewDGkbBxyuE9AedKwFmuvyxmkuwpvZLxDhP0qcFme65c9OWukuUFZ/bQond
v///Mq7C2ROlX6/KP6m2GHwW1V6QB4kbBcz6ahhbu83U6ut+SS4T9wA9ZUiuc26p
E94RCWfMbWIypRn25oGSAZtFh16PxDCZDVERIOqfTycFrHM864A66b7NLEZl14Ty
o3Iv0455GTe4ddB7WUzQGyBqPb0TftG1onIX5wCAqZxyI3J+RZ61kJIMmiS2/qaK
ZkDJqiXX2HGPUo1pJGcdbYanejoW2jX30AfKJcJOiickXJ8k6qB7DZjwnrmANZk7
yOGAfcylYW+A5FngbLQfidG+9cEukq9eI9pzQQTxXB+f0W52o69eAV9fYROBLZDC
CP25Ahji/zZzIjbASc2JmmworoHqLMmfd5++hZcSnAYUsDGC0yegasTpg0zKIBpb
o6+f/D1CcKgBfUKF/hzi5HyOMYSSujY2469sXDJVJEtpH6APlokwAVMh3PSYKANv
7+QXqgwUmBEbBJmpw1Ce808wIWr+L4AqB8Nojsv9EUn1xqxqlQ+oJ+4CHNYkyWXf
qKp7njQuUpBUl/z6cGjT1tM4aSj86BXsqq3W80jafPdTVdb85nyx5wV4FutI6R9V
OOLGCkCf1Z/ehJUb8kRFnf8jqbMRW9wIyfXuiKGrQU4Q2+b87bZZICwGt1n1kQ7r
dVDFZ0BsIabd4+HH3uyn8LgS5/gtMVDP7M4zY/8T+Fz3s/jQPs7DuHA2SEbikSFo
Bj9xstOqBcejJdQC04/+SejDE4oh9EjvGgO68vbIAlmU6UgmWn9jGDNm7BznSjJo
GPQSQvJJVOE0PEZlrZalupIQPs8YuLFDw2/Y/Lf/smHFO54I3/kDFW4xQ2Pbf87v
oSjIgsYrsxydSyL8RsjJWUE5kB8qxYXbdfTMj9kukuqMKGrpDfO2Gz02//wUTvRu
e9Xa2jntZfJcP8X2FYTUze6XAnEk5E3tMtmovyEeqIvmVInjpPdv2cNYW6Z54Wkw
+o2GqK9Nr3bx/rOHue6S2yqMZ1SYQ3mAsN/rn6GEiiudPUliDHSmS2UevuVv5sRj
NaSO0w/QwV1vXZbf8vIcGzkIBZaZhnXhoE35CUZ8DZhSeQROPXPLXFl0eqPpB0cn
///Kj7U32zfK0RVlm5pVdgzQsyGLihDqxN0AKduU4LdMu9qHpJQxuDcdDeKgygRs
AetCVvzpWOC77BjTP9P5P9ag8Zox9c97xZ4AE+/11uNI/k3GSUPk5RDdbFx5D/om
4RH9e2SYTLs9BxwbgDW8meCqqC6d0k017Gux+1Rv76j0QmXEuf5+Y4bVvNITI55h
yDA/MwaJpwdKxb7YHtKqVZAlXwnyeZAt+RaldSFNv1Qk7oxUiRezDqD045Jy1iYk
pHFXisBFRuBupIJFz+2BFXdTWxP4aEvwVv7xjWFxHZm+1vcT5uNdnNUQLkLugIZa
8pW8AznwPdeHSdTkx2Hejja+5t7mJuGDp3VEjPvood6XW1oqsnSlqxHe1vF7jJE/
Jfq8ThWzL9UJY8rjT8AkOdAdXL2dfPSphuSmuqrh4ckI/ry/iwgYKcCF1pAKOuq6
Q7AAY1UP62ZR3UY2/fkqaCbPOBbOYLMcxLr5Rs+TuPCmc0F9vado/NbmWXXhQWaf
YObbWPeOADXT3lT3CKApcuLtH34j9UnDwhgjC73BIvYcyqFNY7aEp6Qph8wnHc8W
FBMIoWdcH+Aj5YbOmDsi1rwA2hR8ije4/0k9GcE0ul8NQ9Mu9Mal6hPJaLFVaIAX
URC5h8WQgCdAyyZIzyxjtWrkrN4HOKZQusg+r6yRzkn+yQxIZedT4MKT2SbXxMMK
fobpW8LaiqmE4nVuVfYgC4mLbDSNLhERwGgpTsHEktL0+TmWdp6gPZqWn5bBsxHa
DXcBRBHJKselUmeFWyEND36gEjmY8BO/xhC8Br28vf23ef/jy6yU57Z1GysouGR0
7bBpL5CwChm4Zj4yr4XXdUzLkGypQn1/kxznKU+YiTtLxXHH6THkM6BbCyqHGw90
mzjXAdkHuPBcbP7uADs0bIScBsxg9LYYGjPRIQtrg9FbDaeTD7Virft2D9VNFxu7
aBeS+DCJ4ES4fBJgJtV8q74nZFGfoJE/FJlnUdkurs6LBS++cZQ8DpbA5tBSCNeQ
E3iBq3Vsv2pkR2WDH5eOxKKVG7CYvAOrPhmQae88p2Q5Njc1HstEC3S5NQt2OQnA
vpoBHEKc7p8LXqDf6UzFxxALfxJZEnOLgqrp1hohTlvFS5peKMlvpBjDhDRUOhxC
8ptdoBhfLPXWsimRICieq/mBnR8ww2R8iG/pBJNPZtkfbA8De/6a8aNzph3zAY7s
d98TvtnR9ZPeHgxR4yZ5jI/mEI5UOVv2IdnP6P4aOToLLhpJ/KbX7Fa4PKSRwbTU
VycdxchClTlces+aMfULtqccW7gADjF5B5Xcs8Qs6haV7nDsudroHeUZUk4rqr/+
TUBIliIizcGWEDWDRb/vJ9nq2Hzmz9KYGRhrvFF3KTp6TLrGfD+FXCAKyZoBcf+E
eSWQTHHFAd5cZubsGRWE02/4Ne9/m24+kSdjx0YXs2jj1YhmnLC0dK8FujFHHz77
Ca+0769K3800pf4U799GOkh1SQh4Vi/Bp0PUprOFLmLFQGuRYEjBgkPjjfkLnp5Y
9VQxFXmzJVpJotNmg+HaDRuvowRIWcnkhH35aEQPXuMyUyxwT1cuAgO9o/Ct8AvY
7HmLUEh+Mtmr9CXOkmUM6Obzgq2inbQ1pLJRWaqN5SNPoV1hK9btWqb6+w/CFF+p
1h4ejU/9oos9NKgv2JGLgRhvb+MJla0czE5fpaMVyvTxCTO5q0byDx+zCd3Qy71h
Lx1+d/zEAf6JuispRvVZQcmvhuPOE4Rf8o4/iVjkZqU0Jdspu+afVV/eIBkJpm1y
BSXtG4buE1jzlLQSNJ8xj4/mzxMZ97OAHZf/HSJy8f1hWDcl093R5p6HSSQGZQ8C
o4c+eTxOWCeRwp1Xgp0Z7zMANFOq9Cst/TXozlBjivTksXG1fWvBbAOeM+T9SeXN
2v6kZndKH8ae9QpCIsd0vEtseRSGF8f9qChp1FhaBZo4cRSagpL/TQlvC7h9iosG
E8qcE0KixlN0a8qLLNpRTWR4bEffV87eRKZiO2b0wcaxg1JezwEnGfejB1zIjuto
xjQwFNwmxXeC/j0FbBlHL4ovqXtfd1m1Jya/8PUN8jKC0rTWG0DTSWBYzphBT2xg
af4j46uN40IRPGMFQ+vya/ucNLmw+rI+k+mmOVhjYHs0WhqYRtUZhSpgyNAD2iJR
ltuKuvEB5vbTilCRQlOEw/FyChbxLp0bzvr1yk7xnDjCJVoNxkt6v1WlIiDI1Xs6
D9jEuj4ApGFa89IlcguJv3I40EvTHBLJM4J+d8WZOUzV+D6GW1eXQE2clutIlXc3
8Gmb29qvLiM0LdfRZ0roopEzaXjNpybZlcCL0tyHHrzf0gfDb/OdsAEKuE7X9sws
0K7iz0TmPVwXPPxvsI+tZ9moiWypLAkU3M0diVyIWN37AYSst6DE5dDU4W/L5oAI
7ORU1mgGutRaqM+5qnLeqvVDT4Vv3tpMzmWFXW5uivux5NLtF75v2rCv4ZDAiSOL
jlYeEtjLl0acGFOfXKUzS8pglgLcEs1OdTPC0b9VmWjuaHbKkE/No+diVZqJ5yad
nb5FsZMa+eV71FwkKKUCqTQWAi3sWr/b42aCGNO2ep+sldvy/PYL0AhZwLIdR/bJ
WBt98+vV21NCrbUb85Na2NeVulLeSEWEruJDMmQ+0H2p6D/jS4wdW60Awk1n4q/1
FcLKF+DC/pV8VbM0ZXw+qIUW6zRuWitq8ymot6+VexXu7Gr0Bj8INYf7UOMlwNsA
wI2r9FHC5pFBbg2TMjLnQyrR0Ca3/0toTzc6utSUK0uXKdHPiKuGHfGdI0ZwRJxC
VDdhW3u2+QGKCG1FMqtJVyep+MY2O4seM3oU8ECH0DMN3SSsGiczX9pd72ScLMu4
QzJUSb3jHh0TOi6nQ+qNwny6MCrktzPsfMrYoFHSQW/tTbvig3jYwaMSXtPokPmC
RWTGb8J5jTkZxO+T7YKSXFC95BOnLd70HpS9Z+L1bQkEnYGK+UGSebXypO2r33m8
qEI/w6c8IfDmhCxRY1aA+zNooD2+5JEgFYgQRLr+SpBE5bZpmOP8GMdEJcW3iPlx
CSbDTd6nPriKA9jPeYoPlHKPPCG0517/5c003n5I2DJ5Y728HiHQhxFs+U3mCbO4
xgvkXnqTKigWcausCT7kaHDsAZNF166pKMvvETMZz8RztVbs/AitsazgYlNoqmnU
zWSLH/u3/XABEvIaZq1ejWjEe2xViygK0oN5VfStKAqQ4wKtWuStWwCmGpkaN1kK
gT/3eDAopnpNJ0MDDIp/gM8OMi+0byjkQNOKBM3rBd2OvzNhcgW20HipBeNjjXmA
9eKXibadkXQhHITrI2i6Jr0xsipICyW9cvIxtI7pyQBKPoLYOx3AokSsmGG1/Apg
nDMBOoNBhFiwn6l1PH5nOWQ9b2N7cS/Xs6YcgtcdiKyPp6TM7g6SsVkpWjQb+jyB
AeGUthmWEH3Zw51I0yyF9coPTkvZiehX5TwZRh+pKX4ckeVfpyx1yXkrJ6GADux6
TDP1HVF2Clue0ZHmCJ1BgBYesBykyyttRvtiyPudyKfi5xKjJF04aizQj6TBdWRP
UC0wZ6C0vFninFKuQ5Oljr+gA6N2XKqB1N4BWNa4oNGq5lWuzGA4EhVOn48a02xR
fEgVcY+fOhyC4AHt40WbMN0jBbZguG0HbEoqpVqacfFdQrUiXyIGMQehAW8m8ysi
bpBUb5PMb17Q3jXvNxwcWQv3ZS1n7FpWKRbLZYVRjQoV2Zk/ZCS7+fl5KXemqChk
h6gt2rZl1X1oKsCtZRXlyX75lIauLcmlJvkTpfTA/t66/7FYHnTgL/8ghX6O4+sM
iDe4YLjUlYDyaZINZaGAYl0MTYWukSzRa2mQ4q/pAzWqt2rHALcQaaE3CZwFoNv0
MYDDxBKkrI6dXCpK8RZseO1RGuz76CwNkNT/zz44VrIBBugVxL5qHwfpx1O0BUW6
Ty1YVp69GSkSHwJFGuXrrF09REx4LU0IeeciGLt2VzWn63xIDwcD8GcvL/EcelLT
mQaZQnPrp2m5HPs3+yMx6+TXWl5Gol4/Ob6t8LfRG0D/0oz/zQYGo3SKgihiY+fO
zMBekUhA//wge/Lfv8WBwiBIiAImYXNbj5zEwgwCGgVvIrvJfT9/xNONBBCreulp
xkR2IKz7BFVUxWs1aAb5T9ZE0047NEyN/24qyjSyZ0/m0xRdB6Exmf9rjEb8XFQc
Ov2D5C677+oT8eXreOkBXUku6vl+bgV6BcusNWCeRSByskDnYoIrX73E+0IlN1Aa
6zVu8UHdapUyru6oq/LM6MSNVJZmlfJ1zPeVcp2xBhmaRQ9kQjPCuVlhEXptq9Pz
/j+aSn97VPxvfkLBnCLaK9FRWbAU0vtGAMZFooqez1H5DWYsyhI5shrRHVBQw+Tz
xWsqPdXUWBWW/huiNgVrsxniRGVf7XD8Ha0yP+GxA4A5O4I+UKDaY1O+HboQvpVu
FQh96iq8NFG/Eo97nPUNRvY8iibo0yEEtS6Ee01u0rwlKbrzA+ghfgitDpCvTHKh
Qq/r0YgKypTa50M9avXicC9TJaKdoUcRqcN2mmPtUAMB4OCC82nAczmKhv9BSu2G
eEBdO+ATsU468IdtoT6Y+dxghlINAybnvaY/sWw7ZAyyg+VdqV8gtQie6qUEmlAs
CDm3KOSVFsGKxtj0v7mUNQt6iLcVwWwAb2PaS/LFCVKje8LeUcsq5r7YZzvE80gP
xiDLIdbN103Oj4pKZzPTUu49X3XsA4O9VF1Mmlmc6zdQEN2v5MVxI7cAtWDhNzAF
REX7i+dnuGHk2jv2q4TpuQ2rLL+05mPzeCAB2C/sOG2cGQ5CJZf4/qCuo1OcuWvl
z+WRoscXwroaCYAHqDzz/4BRr+vRTSw11olUW9OPR8JrTYeMnqu02JBwh4sdWU44
XEJ0dbBsINx92S7IrmWjO7P9lE3z+oNn05mBi2hU1HmaICst2mHFS7U9j5h1XwYi
Z7WA+t6apoeIC5YrfqlDNAXknhkC0eA0bv4MisTCbWsicna5yuTxZlrx8BjDH/Sn
t1bmRz6IxmUADRjczzFwhjNfXohkyh+y7K4bHYoDoqfTtP9qVzCldTYQWLUoY/EL
Gkg2do9iE1HpTIcZvS+sv3NyfeJ5tS0IKTl/FPINxQthoW0LnJRVgYijK9aptPx4
cj9bmb5pWGPIcg+y82PX4Ih7iKVr1p96cy8U5aY5Ja3vFkG3hkZPhIIauysuJFTP
ZqZcK/aZhjaTVl+VdDPIJwGMPUrxm+nJMnsYcoghTY19NA8ZtIrTyW5c23peySH4
1HfE5VOorV0EPGxzbkl0AjfmvYtw95tkvtSI6qy+wqRUbXQDm9c46zaL3XBSoveA
hIs7X4klVxKuD9WdM3xR3DzdrqYga8iAe2XZfqW4N8osIl3sKqnhYo4b/ZLV3mst
gMR2kdVLfqIMVyUFUjInSIzFPnLh4fjjkCelgjvdbDpyoUJXW7ZYXDPjOoXhpYjO
hX6gFU3dMYIaVsYJUe8SD9BYyjHT8LxC21gYzOmsws94ZDq4VVuElBnQpdRYwGQl
P2y8mhtiX8B7lrgFZmTdkhOTBFPh9I1ByJ66OoK2Ahq3DKLUyFSNXkqqKGdWGJN9
yKNCM7MUuHBya3AU5hXMsJs3U/KenW3Y24bH9S8sn+Oz/mvFc0royi03W63YBgHi
5nhOoZGkOyz+GSSmxuAoJO3zbo9TU7Wg3ci7K6S8AOxD33QmGAUJ5Z6cHpofG3bm
7Mt5WdRBuzudsQUiz2MBUyYvpqOZWvfo2o3HS2aogxo2BD5h8YY7p+zcMYy23YMg
TSn1s80rgNVhWMErday+OwHsnHbeL2PvtzJjJ98v9s7PQdfJlIgmLNgJXAUyhG0k
w5w6JaovlRi5hxB9OpIGFDkwF71EiSdFZ8hI/j6TQeNPM8cULoP3qNPJD/vrWBQO
uCqgOxz5NYYs7/i3VBKNE737/x8huE6mvINxFu/POCrA4CsC2SRQB6D88lEIchFP
3w464ULcHPlp0A89pZmMZmYnUwS8gcy/OlbRZnddpVyhNAGsZNPvZ8xyiaV7+SIJ
m6bNiIKhJsi1qDzLEa90jasTtSWmDQGqCYvEZVmJMf+64Kwyh/Hq38fniUpXox0P
/KW0Pmm8GknWM9xmcKxObpvv4F7+q83eIshy7hWMMXielbXwEqi5GCOuQ9AdHzOo
uD22TEv6wKqHkEXFFOYzNg6EpGf4vtvsSUc53Tinra0FESXAPaVPN3nrZyR/Vnq0
A9PCbaUTEoYg/ku9ln+H0AXY3eDmKo4sZ7+/6GlDXuCsbg2GRQLVaOwkubCzn8Ca
vNH9t6RfPFvgBEhbLj4f0hLmC9fVqwZGEZryPDKPSdWrBcwoCYazS6/RZWKXKSYF
ZJA9h18242FEDvzmYTb9QTkvtYe03aY+jAfGgpr/SUkHl5OJEUO+syuUFnoBHKOc
iepcALdKfwchSLzw0UlEvxUuVt1Q+CN/U6D9vbDG+0/Hf4DCZsDyyvszlHgoEPbx
q0a2obyG8S4LqbCW4Rq84EJ6qZWn/Rlldf1Av9HfVBlrPTYUFxkSTHY87fKlkanU
xij7c28Z6+T+IKesOmogC43Kv63VCbjWitqw7Ut33ixWvsKPYh+9eGBCqFpftLV5
hKSy5+8/tx+ScjHvxJMTXLmpiBju9PHds/TuE2QbrcbadtojB0UiUPyanPqUNwpX
igUEmyb3ZPQ7z8Pl+mQdu1jPkVGQqJVIzCmO4FYrM6AGNUeqtSmfDjPYOVE40J/z
2424EiNX7ycviHJwb8MEmB+GirU8RYOpk6NAqTkHLIyMBTLP0RY9oOYAnN/C1XY0
cgMvEjHOn+vZw6Cur/jW8iR4sat5eEmRPchmWqtFB0R4PfdQonjls3z6w3DgzsXZ
V7tWFhXnJjHeoWe9lP11C0VwHO4X493Bp5xRQcxT4E/pTkcyh9wYi840yZ4vppD/
ZCRpaQrXqRDF4VId0ClTwsynKZBzT5QEOWAPFgCp6kWl6TimDDxRtJuFO5dtdR+6
dsKN27MbtE2gDm6lt0B/jwb7e3S1Ra1ERH6WAynpQ41s1JyncXNq3T+5L5+PmzeP
9L7ACBj8JC50ZqD4OSyTWCERQ+tF4E81Rilxd3z9hbIgwBk4Y8EPQtoZjB7Igngf
u7b4gzO/LBrKSza3N+CPrC5+cJYehy7m7xJwrhfgCunIoNa6e92ZY2K36j1rXLiN
RiubcHUuSqqCz2+83D+RLknZ3lD9YK6EsWfVHVt6oBa7CW8GZEVsbeauxhyeiJ2l
cwzYsvFYCNioOlLi0V5/Ri3zxCL+wXHE0pD0Wa1+YTdOcXjfiTm7WqfTgWHSXl4A
AcMZch6+Oz6O6lJgR4txhgU5syhJVPWDa384JGv5216V/CQUL4sp6J1iQMgHUOlz
5rtZdA4I+wo6YB/zWHTGnd8mMDrmoSfav/3hSzmuksRC5iXZlRqBAXvzJM6O7DfF
PEwbW3jdQu7+bqghwtB2Bl7xJuQ0D+ctX7O7ODmgyCuGeI6EnQCHxECqPiDWrpvA
ORMzGkeENS7Vwx7jTQhfNGKfW2Yg2fbmncEk8g6Xsz34JbRzz7EkLkmxebiiy/g1
JnaWSpeAusC21WlmDb7EUkekbaWM+aqInvcCla/2m63gUCQbggHEcK+BHiA1ykbL
5aQogqrTVUNnApHuqQVyg+1lUOIJFRwCfVrU86NOtz9Ef4zDyzP1LDYkWnypGImE
Koyyqw9y9bJv5TngMR811Ixz4WumRytBNN/uKSf6evXlzzH0g2X8XoLa0mGd49tm
hhn6onuM/EUMO52nN1gTu62cl66H8gWbMOfijvEMtZAdemuahcmoI9Q+AcaQny9h
BZc4rm3vIlvO78tVP55U55s/pJNDlLmcdYnODWTawR90G3mhvFcE2hPMZqgTHkhg
VIg7YnavDVrqXMQz2FYnutuwEnmybpjMsJSWc+mZOuhnpZ8kbfFhfmz6+QpZfyDt
lQ9gPA7rrnaD+Fq9KuzeLUijjPwvMrbpfmP3+oUYwYF5Y++RQVAYmp6KR/rdobbt
M1lHZhqiblc5R05AO5Q//upfyj2KOvize5mRqgk+mTahy1ubPM+AU02rC5vTGRIO
3ENEKzJzPDxYWP14iuuK01cApZfzo4kJ+3Xj2CT4+NnUrKPB2w8JxU/s/OcJCK7v
0CZCrRGPnyvBK3Av8gIw5kKLjj/XsZzPdF1upsVXuGA2GXPbytdlQcVq2VtF10u6
OttE6MD5B5NFIWueHYyIXZRX4wPyWerlnwx5vSdaylWfp9/1vBjsWbrdDx1gb6gJ
DIgQY4IfToNK6rDZ74/O5HIdJXM9WJIPioiJuvT6WAO8wByaimLk+BJH3GMikfUg
cvlJil5szkIpZtlAUWrye8KCVj9DwfkTMv6Ynfaz8ZSHfj3tq76hJCaWCULpb2ig
cyHafLP1KGank/bQ8m2PwGIDU57SZKZFklTycMitkiFitLARJ28oaNnY0tWqJkeq
stDW8CCGwXr0lYIt3nI2bDLgcrJamvKBRDufeHq23yRVc0rSTm5UTNX9uRau5JYZ
JHZWseYVZ5cFZn7rVJcLKnPU5NVD7Euel/fpyb4WyB5ahucawy1HCemJDQ7kdXjt
NdMx/3+x7GW1J+t1MtkLnYNVUNzu0jCPgPZsFpWObL76RbX/LN5ee9dBhqQyAPi5
+uSa3VAm6YoS1Gn/tueHcUVg2N7iyqoXMkz7mK9n3TcHOc0hV6Au3UHni0w0c/wG
KUu9+bs9KE4QzV8wVZpLZpyaJk6RdZRXVyQcNqOVQ8/ZbAVmIIjSzRgUC9C+9LtJ
pOBNfldeMucG72vrwQr4bRuZvmxwISC3v3cLlN4KWLiM75gJE/jskPNzwpoO9i+Z
LlRJ9ixNseZrCzrUT98TXUQIcjps4xvN33tCslm5RMFKy3fvBfZCCVAvOvTPd9xI
0j6/nyNVJ8CiOa+KLIm9fxD6a4guOZTNXhR7Ax8xUgUxSL/Dv7wZZHDVz/Gi42KZ
CPmxi935C8/ZQuwB+QzLlW37CFvBfeTdodXCassFCR8VoWXveKnGLdqATqbzFpZe
ka8KIS7RizVZARvlS0TovU3DJFSWWcEtkSilZsCPt9+GsE2RlWsNZ6JTCyHUIDxo
m341wDO0bLdZWvkxJTaADr8+a0zILvH1LDBSjprkrQ7CdhTBC4lbf88pozecb+xE
1d/S3ahpUJ0CG9X+R3+6MWHuoV3YhZHvS34GwGuFjkVnsfRiLhOYcPtowCeKmBQs
jVw/7Wi/EnAn4oLIJp8hMTBjFNx/00jf0ELa8gmJKxkqgXxTKTpn7QRtHkj139CK
Hbl4gl+8CLCoKCuMuNdQA/57ELDkCY0c7jzy5SVQtnrmC9uVvnfLOPj2df+LyTyE
ISNNrR3mC4kwSJgELV2buv2R28Nkoh4IxaWAOL6Nrb0oub6ghOgDeh7YB002e2DJ
LvPJYYnqGIBW4b38dg5vEvFv8VSB4FIIJQyhxSpUfICp+tsc5IWWTpJVaMKVJbqQ
eharbMeiSKsaUNYR4oTS7dd4t5S/6Xjncqppa6vT4VV3E4eHeCPZgIXZSxaJ2Jow
hOdMyS9kRKox0k4SXKUIVj65r08i+mjf/qMv1rQcenY1niRH82dsg6G+gzWY2Kip
3Of7CG1OkkREGnC0PiD7fQD59TmTALs8p7d2tr+5hBnmskGYjTixvkUSqNsaCHII
1+M4p+t8/Id6bWhGSvD0Gn5S0fwPF19uBY8gr4WCb+Tiw/3uUB1e3nJIdCtggRm/
7829pv2At8+CV/OV7JYlr8F1jh+Z7vPPdX9PK+Fd/k6x7obwIqZJZhMVT4SwkZQq
t0HqMZs7NJ8pSpt1xm2e1bMLKhZuPeRm7uaGs1d92NKu/zPbJTjyeCprd0VLrOGi
+ptitvxr9yZJY6pT2i1hlHuY/WpC6Zoo/BdnAAhnwU9pawEM7uco+K4vvIQXhRp2
rmXsvt+c4h/3LIy/ZbHcUa6lBlE715vbgKWMtofSnm7KeVgzxdMM6ZOwqLFfMAY9
dWPQG/JD0gD6jJRRJHdp5Wz7hmZQC8EPPtxMo7uz8/q/RgJ24Z5nt6ROeN1lqbsk
yMxXAvIrvq8HliLIz42z8A0lYklGfV+tdBOnmOHHcwz2cXlluUH90qnJhJUOvqKd
qKO6QAOSKnPkUP7TAo+PSrAWRpVgM+w/Thhub4OzfYsT1wHHHeZg1eMSnQ35fnZg
vET5nUfIAh9K53aB0Xe4mqm4RKEFWNsj00GsqxxGHc2ebiDNXPyJW2NDAKsRadF8
WM2qPnRvgBEOC0xoat/yZXIIOoGqsVxmQ3CloxEwcgnGNg41mfVJzGgNb633S3Jd
uPP58V9MWeer7fGmu0l6HMQ2igCMyJZydkjthDDg20fxrr/z/ttBnpeI4oG06QBP
FDjq/WIV/2xOM9eb3NDnO4xaJlT1siXtzVK6LpW/glLOjkFiUFH5IOHMnYcVIl/D
Qlkxlkc3UXWkTkxVftcoMRuF0oiI4wt9jhSYMRGjagtgiGY85Ig85++KSGExLXGN
+mykhHtFfwzHJ8le3w/4Jv/0BT274DpiOS+RaRsz0fdCTXr/t4fP3TS5SXlD1blu
rigsYou6Ej8avrrE6qHMuLLqZ/+S3vHG9obbX3JJdODYk+WnVwyORuHhWow7uBeb
SV/LyhPgi90YzS7Wq9UxVyFU6hooCR0JwfUHbxQvAZ+x6QZqH4aVeQwnv2BPo6Cg
PGoTs3Re4YvcR9/17w3Q6c8e7ar6FCjGr7xdZxaIDbF+ljf5MXHPWZ7Ha7E1+HPS
h1a2c+caY5+cHka6/5jfp9YZ2qo7+bdMSG/Cwqd2PDXbLigFHg4TxwBzTE1pgHjY
aQQbjJolAB0cRQpWNUzNdeU5CD/qv26sagqQ14jvOt/rEfIDuuEQVqNFNuHDBB+P
fHUB0r50qyIaaTK6KkzhTEUlujNaEG2kcNBlR4NXTPbTr/wID1F1x+Lg0csxupTR
b3zQTSrX/LsjIUlRKsbsZNs4TDPxavXkIptrknf9CKxN8n2HOarTq/m206SJ1bR0
q5bnI4R31S0B7QmRLoYRbQ+A7qBMdk+4P4MnNZQEHGRjG6bkhiIHJZY26eOMeio0
TPiTuEvHxYsWVWKb4fFic6QkfrpMw2/0yoSD+V68h0cG0JO/uBLddiuUNF/62H3l
XLUhPiCd7PMniw39hUu6AuUU64ts7mhHxDzCdnf2LkpFMkTWOZ5QcU2mrzw7B50a
tb3a+pSEMPEY0rXa2qKNe1X0EGo+PGJ3R5WVisODF+JqXcTt1zGNrRAUxF5KLGof
9RCm2lwbhDt0UUBkuIAtDgAG872dB5x8SKGDyNA+xbQBHoLERohXNp2hhIclg+Ht
4FZTAXuMrI3a6mjGNdXrTKps7lnmkwwe0uEqVXErwB9jzHuUUkztmuwxlbUGB+FO
lycWzD+Azbs3gODFCByK9PWVFXG4gTTcCji7Hkac2W1kKyixOeGcI3RQta3GPRou
uJ/21hg8uvXxxrTv9C0+gblOaWweyDUzZEKPygtsVnzSBxfZT+JnI7vJQSKn15V9
hG6lm2wqIzvFuU3Vhw3ArO2HjleDOVMV/+AuxsBiWaGTqiNyajFNG3+8WwV3dqsm
FQau5MWT8+6286gsadWBTW1qzfQ+haOKt/n++dEkDCR2T6lqThNiQwA67HFf9uix
nEf3+FEEq+cErADPwWC/F7fg+hkhdAWvOmq92jHLJrs+s7HlJfi2s6mTQX3o0mnH
2u+ru/Aox7tYii3t7Fojvqtr61G9fliF3tev1xW1+XqI+mNErLn3X/rGKT6XOwnl
G3mzoLNDR4gtSltDgYVS+YPOMDTVAEQZNQiSPFnc7QUcgN/ylqK72FMP5zQbkRq6
DrX6ERrfFJeCoyqKH5d5YxMAZEgrEa2/WWCMTvSw5ajEYv7aGiBkkp5PTTxC8dpX
NdP6GDIO8IfG2vcYwphDr4tI+tYc6OJWclBrdMBazYuAoMBzjmzyUosCsOqsDrpg
boixHRJWHJrOXtJ48rKU3lECXH+j22JwqzVoQ/MJy/IrX/4Ac5m4DKAIvOX/f6sQ
5lzsOJStlznZ9GVnhSDjjJDQi1YUehpOfMa2Y+HUnFUAb/XuUH9JKjpXtf9cwKpp
aPftmS1EoPBJybsRr6Hz/he1eiA4nzW9rHkcUt0mMV5jsmxs5/bSl+0s9rqh5IJ6
C+062HCa++QINkUy0PByvWc7gYR61sraJZtTfJw1B1QRkqNriYLULHFUr6jUj8FG
ulKKv5M7m/J35LF+wps4gOcHsZTFeBOfQj9cZKOOsdBEaXB018cso5GdZZrj0/6R
pLAeHE1lLSMRmeRKK1lnc6CWZdPdDGGFunf/Z0O7G2HIvITgKV8SfplwoA4JaLZV
ko4FX2dlQty5qvGAHcAvh7+yArmTu1UZIdlIhruAOeluV+jupLDujQQTjBzjq0H4
C+W+nV3xenUCJgVnIlFbvjOyHouGHZMsnUVxsDmWrH94IB5NL6E3Lzi8o2HKFJiQ
n+q9k0huRCYw4R3dHLPNSHyhx292GBRm6j85Y6tcjPyIISE0VQwQDdl5iZHwRGMw
PUQoW03jmvZKDVTIhUl2lWE63bXwrzqqFj7QXH6ZF9zhD1+TUMSY5aylt/C3sS9v
VCFlpzaA/oj7Dwrm8GdwUgfctSw4w8M8TWhT0WT5bA/G0Kla83unG6KVnWDNYWmZ
VxinimcXJBtqg7K5iPWc8LZiteZwkJzfuW9LX2eOu4hbnMbapmkU+15Ty3dOd/Wu
RGujOZJV41WrLNg50VKAaBteHyoMRrl4sHAX2UFNAoJNmS2aGg0x4eiTVMX3iUHE
zG+UdukN/vL0hkif55ets8o9D8EHR6P9X+9ki3bQ8tVGIoB/MYFsG5Pks6t4LtyO
634eGLiiUbv1PlurES6YwmoaiVasC02rtRiUoyvaZiH9oNtIf9+EsXiC1MpOMOiE
/izcLRNfQyCUrBbemW//epjpb8Kg+mD5hIeeM98ULbIiLJDRVWdz/p00aBVZW/6x
d3FgY/oNIxT55BtG2u4+oraTB6f+2r3IuVE3fYmjKQClhwr07b05wxJkazS3LYeO
37bLK274sk+402NkdozVwx9J8XiFfd602YBR6fpCcSyKmsO5+8yqBjJIcALHpiQ/
qwj9UVBrxceIgPDUaaXAV0fzLM085eceTXzLp4ktUMZa+h4W1RBzyw/zSPl088ZK
9lF0zgg3EjClZBzHyfSwL/7V1Svfk0UFDRsUlbzgmvlMqIwTQ7VQW+5dTVSZcjyy
mFKX6X1NmR/IjyUSqywQG7/7GdDXjIfJJzdPwq/rPoExmIzMB2xxFFOmAcDeprF3
9db0PJGcRoNBLQ3nKI1JP7EW03vDb2yUeSFfGetWXzT62YWW7sxo9KVC7aAa0Ut5
tXB/3s449/YZroCqjzYMAGFLPDVyqLzoztBqR6yUpy0oUokslqnYGkvmtfjulgxC
dKTrVXLDXnbo8oIP4XxSrCsdKNCfr3jcsHDqjzj3RlSWDJJ7DCrgQIHaB5pafNop
pcLDhD4TzZXp3eRieXpx1GN/oji+ZQInzfmnR+Hd1WKyW2d2L+0gr75rgmCVO2YL
6hO6EodsD6v3FwTFJfBx+x9rJM8NHi+fN9y+Lbf77GHlXYBdBgNEfNEy9igR7QLh
kiP/tREO6nVwWdM6ZPQu/6VtMia5IPzAQtZeKNgwLvNFrIyYMyxHCuwThAqkSTvn
R0QaHzkPAMP7pmDDrYZnyF3Bh2RUDD30dsx4GzYqX8+ThtyZy5QLDZncZOIAvzRo
PePcMBfLi8dwdehar4D4t9RIXGgCFBYmkH/yCh4UfMUNBk+FWueHtd4zrl2O5Oo2
rEelzt3/2yUcmLA9XxbyqW7wbNjCNMxVLIUcdHO6QEHjJ+KgL63c586HAOV3fxMb
ch5bj51sgJux4loPRrh5rhfzVjx8mgsEC70ANoAIDTs1Vc/eGhoekYef0ZYODiPD
lCZ6qeRWoOt6lIgjg39Ms/oAsE97qorkXjBmcFkArHfkjOmNKe0Mv1ObbAkqn3Ra
VcnG3gPItj9ecCilEm6nU7aYyjySfMuuGKDo6zbbmZBDgN2HqeYeL0lM+0pPThuK
v9090vAc8fPN1YefP+ad2w+IfDuK946ydL4W2hdRNhQv70Hzx+U1m7fbAFChOHsK
eawTw4Z/3CrU1r4hKABx7UGO52sE0WthrMql4bGX96+0YEzyqLs3kuEpfVUKvH2S
Jo7CABOGcLf7VKNhQCDSetugpiJa33N5BuHAs5dQWAE1rhFgUxuiDLOfK2HrZ0pa
jip9qEcwqOHAyOEHwh/HxvIXa0Vgj2XxpigBGzxEyxEgM8k2POG7c6m/JOKp5pr5
CH5tGte1BzEeXbdYkhgzklh3bgVc/fb2vGLwYRx9lBsOUvTcU2HjtTHXdExwG+n9
YB3ivniGvAwjgoO2bftDjINacdEpV2QfkDYSaoUOcYJZya/D/3wqccVvEm/vGqpv
7F2ncweNoDEUaLuIxdpu8pRvt18y+/jhByny/cOSR/3Br2Z6GLwJK4Nycj5kKIU3
duHyx3jPx9pwSTIcf7GfuTGgvx2iiKKy2jXYUjrjm2Gq6/9926bL/YrwbDJdVs5E
iDvhDI8KmGn9xf9fLz42pygsTtEQSHOvS+40OtRwGEp+tCrDxQmrZZcQg11QWlaW
N5cXPoI5xsC3j0nRmki6nDUC9ALoQDT75x+anj37Fc/RZjF/p6BtBnWSxLSSg5hL
WAQQXklFAxt6jPVNtm1i3pp/CTvqj1qyK+Xm4vupNwE7aA9C4N+kOJ8PD/MRnqwr
xuSU7F0Q2e7kXK9eN5MDaZFCvT0vipyKsh0FkMg+3dp7VYrzfNSGathQCgLLzd7R
EzusKkjmlEEuduGbOn96DW0WYlY7LVszRmn5MIhyrk6WSXB20JAFO2qIk+lR1oVL
P0Cg2NIPcVo6KZHr5j38MOk4bZEgpg9ugvbQF5cniuvVnbNEPQo5+UMb0O+zWnDP
mxffJi8TlcT5ZHa9YtgTV44849JO4C4kc0QHzO6cf9Pgdv9/5A3ju6IaGHXujKdy
GOlbNz85+9HuQ8ULIsjKCpAk7D8wP4bvQqc/tumhpkFtPJBzdDeCfgmP/XL2r5sz
OunOJdiQWt7RK+ozd+V7y+GJ5BZjIMQ4tyWW1w6k/9MaDqze9AxJIvGohVyj1p3y
uAqElFBByfLDwv4hTCxAKKWllVuFkxMCfIC3Thjxk2eSVBkMQuDUL3JXxO5KtyQH
WQB/pW+ZVfBX3+Cy/V82RyqaQ4A0eiplTW4bXXYhycbhcQn7AaXFX50ih/Ch+11N
zPHTSFPh1X5hPrKWutEyEyAu/+aHxLiWgQKIJOyVB70dFvTdn1CTwSZs2UYaf55r
2vJWxNy/X7wc7pAd9w20otAMxenarHydbVr0Lco7SeRHqkDDg1GJvELDjLuihiWY
/BSaru0iUNrJVVsNsjZRgWNA6euGHU43oZL2T+/H5BbePfnFy8BYyTveGGCVA3i9
6nTMi0KFKo3VHAYBum5lbyq2Ssm7x8E9euza5UZBx3zIQ/y7VR/UOC5Dx7QU+aXK
pv00AS0I8v1TTi740nEUiItg3BXtfqOitH5WUXps4LJ/wCCTMNXtK7eW+SPX1tbl
3zxSqHVZSjNQP0FqkOZ2BJ1CLs0zHXFGbdw375R/u0Ly66qBOFmIlil6Ozho+blK
T2wO0z3W1y5z0kIH9e6R/yDZCVCt/ix+HPlRGh1PWJcXnSc4u4lQLYBPQREAcCFp
0IRyhmx4VKMFeROse3CrnSep6vEDBkJPA8638kmTT090bCLIJE6xOvXdC6PCjf40
iOX6hiQsvm2wyCbm1HZIbqgOddvEuB1W3wIP80+QxQhQ6IbVX+Af3eztyIp4Qswg
1RJ0Rkw/mJ2B0YomDp7ja4XfKeEEdYhyVveDa0uZ9iTZe36GK2pWttoYW1LjDLvy
UgthEb4JJmrh6SZjbcH3SBnvwzB20oR01HB3ejnDBQEeU9dJy4rugoVNbvhNIXH+
CcXqMuEoayS4zz2XfCgo9Hw+V8bdj46mGo4WGtCjQShcKgBwqOnD8NYXa3JjZJsM
8kb5kofvBKLJDadLibq/PCy1XGPKjVK9ZOr7XCJMV+8zecAazEazKMuhR2RDf2vL
35IoeryJCDmRUjjm1bvmQfSFoQjs0S+P02bCHbOxwaYI6IR3mPnA9yjzJ+AaJG5B
4V+Dw21e3BTppiDu/FtrHZw3o7rJ9Qa0JcOV6KYuQ4UEAlqhRzzfU/WsD4f/+6eC
+KyS1hW9TTrN4bVYGlAi/wN9PRGCIN3Ae/tgHwqHjdIFxGQZE5aBsYqj2iiQVNYY
umTfqOlOQg4XhpUJsSbPIiWktLB83RbxkYRhnNF8Zg/e5SFKt3TtHIbUxF9MseNb
A23AfKygrdmJdVeUQqq9r3uDBOJl1OBZU25jDANZidCod2z+nT8Yrh8e48CBYSGy
uzikV1UQhjZbQCs+iMWqEAkrCDiIrOQy5eBfBcoiWWlxjoJq/khkyGbgwsayXfbi
iS2H6nbLzPNUDHv4sgh+RQLJFWDofxAuL0lD8doFEeTKDt4rrM/h+lDYtrriVeqg
TzuMFT6Tnc4MGvO///fMIagPiXJpdEB5YdYsB8RUWS4KZDLcyPQZlvre2UtKpqnx
KB2+z/0kJ3Lc/tHszXpQCmZpNilZ3/4OqSsAuLvPnvHjbv8wgZP0FKYSTF4Ludrv
Qo2JWKCUvKvSCTWwo+rR7uLRoVX1VAqZxyQURQElTjgK89Ff8FqYxvn0AdxR8g/A
Bheu/ke8SlZGgt3v3VncXNT1chIppwox0DE+gNc5xlqlLix/cgGeXTammBOh0jon
1ZvVg3kXDxoZHdC04pdC4D1qBxk0oy4lTpsKlR9Tca7idnS/LOjcFBTB7Mko/oF+
00Z/hdg8T1ohicvtpwYQO3kOSWxYH8Aryi13Nmi6tnNqUqWLpuKX9IZXM2hH2ksm
LfwuknfjSyaJTA7Zw/OwYS7fYZ+PivJI1AA1PTTRbXgvornyH1+eYrv9M/nwUf6K
iRfBNZGZIiIguqIOWBnoj7VGg1Wf/ypD1tz0JZYV9B22JMuLu83n+83Z4CNiMOXm
jJJthiUKDafdlkjQArSf22Ih1utprWtzUHtbxUUZAKm5XDvlOwKvymlrc/bTyt+u
motw6/XsqjYHlXT+IHxRlfi+Kk9EZs6m4tIVx+ZBVAwFMYFNgmNZILJ8HaT0F1FM
f9MgtOdpSo7lyEw7CdUZrBbEyNgy7jbqoX24HBWVO3OCTAu7WUVOYxoc6nnBxXal
droWnIsM96RK+G/GRxOQofhd7ZxzkjYnLxgzq0Ki44mNoHqycPPb0NpBcaXHX+HB
Mn4GkhTQY6HDgy6AcuyC1HjeDBQdpWvvCXSlEGxbFpUToDxPBwuU0puv3MLka1TA
fZItk2Too/dhnAw4NOUZYHPZbpLH8/117YrLOnr8Rnieb9svtX/6kKeCC/OymEHb
QALjKhYQvUV9xW9Otr+VLGICqTfYK+Bgo8Wb/WfqVXp2gz+UWosF2A0+K/rs0kuN
dYReNM/jh+6JmpfNajyRUYU7GxqwV/mPscj1/+W87tcAxehz497zuaDR1XbHcbJA
UPYyaYeVGyFZurX33iaBslxsndxUqMRA5yjBjoT93Pmwh+WIIV7q5sBrugtfYjUp
gKdkyWnttVSeiKroSo76x67s6PwzxAaYqfSLOMt074OyXKtm2+WK1x5n5Qiqx5Q8
Ro+cMPLYltDcAV2KQd1PP15sBEuoiqYFy1D51PZx0lL84i+a54qVZ5+XSUuo8Cne
ATw3iMf1sO389cizRT/c8EwTahQLu+WZzUhLt12+gw0p9smacEPLCJNutxb5zN1j
pJBXQ/iXcTj0mNc9nXx7V2Ar3T+Nozx6OsJeesGW2znRfxECMZaxjixb9rbaa9QK
Od5le+0NIwiowg9xYSQngfAYR72uxiAQl4ccROiEPz5gMjp/CEWU7wYcfR4bEH25
OlcMKgE478vZPr4JvMJmnX3vfoDK8Mh17Yl3Qu1rAT2HG5jufB8rY8+mESxMitE5
gkB9AA9qTt+7Ebf0cqZiip+FJ1piflKMgMuMFtS78V+29GpeGnGdmwHB2vd6+abj
uUQILZKvhtOFSXRUJf2wNYq3kx0gm+12enb6xY3/OzeJn+SL9fW5YNZKvCz9XLiQ
Gmw9rFVvJFfVnXGBlrw63IMozF/nvTYWLpcAJEJFD04wZ7V8obBfT0l1WlAqz1Bi
eBDS7AOXv9sDZ/Xg8Gq+rHOzswONpEtkOALU70WhK/sinE5eeNvvVIGUSZ9HhS8p
dr3+24HujW4Pl15h50myoCyU302mwrUw0g3r7SOUJnRwMtjQAwIITUZKHF6i9wtn
lGf8KgB8lnxyT1bX3ywAtANGYx0frXGGmUSsxXWdt30JUzXT5+rj6B7GvbKOv1vl
HOr1LGgoYJ+XxKBVrnWPiwPabUhfmYuQu7NSY7cQPuVf+E72ZWqfzGIGxZusoJCc
qRKJSMxy64TIYYlAqhWIZh74++caqURuVa3WC9TuGmjEow5HcoOs19rCoBDYd/Qw
E+TzxChItFr9iiK+VVBkknrj2ZBv7+baNdkpGxHTgTB7B+5eV+dZtdPoam7PzAJn
fRMHlgl1CjMRIiiHqZ6fE1LA52MOipA8DZWx4U7wR14CK27pytHL8M2w1TZ6V7XC
M8Y8JKaOXguB0Mn+PDKsN2JLdhtAeNk/X9tTRlcrrA5eRFUKpS38lv/SR8mkJG8C
z0CTVT9AHj0hP1ReQf91ubCR0Gt4N1NaqBl9w/LzYwfhpJuwAoLcpBBXca2gYS+m
657F7Rc+qxfdmiPTt5Nox8y+KAKWIn3e+zso6Vnivhf7IpXoSzJz9Zy4ZDvbdobK
WzHg8lq717MgPeL+RDYgouyzptRoPKTcx6k5uPUPaxfMtwdGOiiynJXOPr275fXY
5bzvFMItyMnN4n+Eyk/F28Ent/n1siSMNOyXkJaQ36pEd8ubrlCdN+WEzsVE9g9w
SmEQLiHZCK98qjmsa12W4uaztChL3MPVnUAr2sSfEVXN0jC6TTqZhIwn/0f87egR
K0NMImKjhMOQc+Vi2GVaw5PIBWhE0qGgXoOpNit5bYXcGEONOb1uOoQp91apKdof
0y9onutpA0MWkGYRf5jY+G6BJwzKzJ9Dq4yZpyAo8mf0T4Y80oQSs6mLpr5zEWZQ
KAr9GkwNXGWrLP3AMBaqOTh06qEuNeqoY5AiEadne+SLHmrgX5q/TUJbBzRuZGuE
qIv0FsfhxVMR9ep39HQM2iz+S67JSBz/TP04bOv3BB97QH2TtrIDxOoAe5p9tJzS
qq4TQfihWVA+VI5uxFSU/HEDZkBIurrn0LQ8JnFOj+6bygSlQJRrWBOBjFQRoljf
gtuaIMoUTCe6fEt6uZOMWvm9NjJzXULhKbfH5II/97WB2oFp2xLzh7/nY08ssDe5
pGCs7ZMCkpBUSlnkdeQMldAYEY8MjvF76fddcQK45P74iyQlFQyWiGaL93s0Xf+Q
8wJQYHr4d/eWuCkZcm2bL+3ClHOQnSP4Ji73773AEiXO7/jKiZ6YfNv5MXtJOjYi
xJvVISrh/GtQN8l/TuEwOJiKh/FH9/iDGYJQ6JrztSaGIjgOU+/+DWHDp8cZhYb7
HMuAX8rNYegZXAVd0bUUcnFvw8bnw44bY9HMsdLvJdTSRUGhGV+0x4o0Au2/S74o
XrDl3vhKTdeiYAvpt8raH0qMWp8k7X7QkqC+v7O8YXKYlq6k4eYjjq9p5pzQ3qN4
2WMr/ivBmgcu+DTXqOoEhLPlEDVST5HAMM+7z9Kme3h4N/BZrpsBSXosCULhAFix
jkJ7KomfoITKqPWM9Ya/RSQAj3rZlnDe0VTbNqpDrpju/TQqxk9fFLvM6d/A7fua
sZYZ8FS6rE3hA0epdoKbVaLQxL5onAghGx2cZMrvWnQPCbfv1iNf1jHeJnk3UPC8
xL7sFpWMLdJGJ1doVW6vACLh22XWacFIAvAtoAGlDgTvbsi5bm1rQWDGAaMASZB0
M2LTFPSKwyHhPtl0dinPccYV2gvv0lTiY/0ophm103KV4ExngBz2pD/PMZ0n+2H4
38TPOKFp1pqx3lMFQLpCeKerRXsjTmUoT5udhbrs8AGHV3Vv1+2AZiRuQDF0ZZeL
bzDg34chhQ/Ur3YO0m8NIw5hSLW43QYk7Br3g70ygov31tmaTCmDEoXj9HWjOt+z
e1raiYPrku36TfJFAj6UIfNT1CJfv7XQ5ZIeTV6RiBV0DZ878zvFja4sBBMBas5s
JpG5OfNNfb7LXUiQjsl7kw5RedYSJS6J4dQv7hBRyi+3a8L0stxwDGqFuJkQJEtt
v/S2MQL9pCBhvOoui3k+xhSr7KPP8+16b5S3LJIojfzK7zNogShio+886/3WeoaQ
wsC8Klk62Y48Es5JZe51abmYwFo4UyqA3pVU1SfOBxGwWTzJPhou9fV+dZtsi1Ru
b1tPVv2vrWpz4WP31wwP0inAknuSdSRKateBH+hfmTTsyMc5yP6tn+sdXVIlg/iS
pjtMnB5pOFDrDirvs7wC3KYLjRYnhfecDxY8MS52d/2DhGPbCGNursnsoJbNAZFS
1vMj93qGT9C2IyYJE/LQ34YlQcGDCfRGnhbPPSq50yK52s+gNEBRo8iTnZY0IPXQ
s34wL4Oagzu7MtdIEJ2syn820tCkFv7a+Jl3fgJeLKyRqcdSXqRz+lOGK8UwO4LB
quwd3aSvqdp0Va77S7jKhI3i9Lfg+6v+E1zzdeswsBvS5L1xKprvSLEuCiUkxY9V
XhdRC1WxIFLULTt3ZdW385zBnUc1lP5tbSqFS/pL8WciNf7SfM3g6TZk+Iw+RUB8
F6ZCkQj/JDawKkTUHrObyzdRR5BvF73A+lnRZsOC/qV26Qjc9X/e0LL/0obKGPJk
I1kN6MbewrKFQmAeE6Uye8QU/cFIrQ1Y7UW89j5WfSjtxYz67vsi4CXuLYgDxZgy
csGnD3U1tL7faw92aKOC++RFNgTTpAN8PezfR7v3MSGqLDcER8nQcaIHynUH7XCj
9t1WDCdtCX66Oltdr54cZIvFR0WsaSaDfFDbtb2Sujl/mVVm+xgWy9Dle0Fy6fJT
kbFhDPrlmKtVOQCxefSd4Y0qGx16Wc+b/4EtCF5q3qi96o+xLoSHczjUdYEqMn2V
LiyJ6WFtthZx+RXhHrkd0KUYlezYmqJdcaEqTmEDuTzQblMAqvwmNIe70HiHGCNB
VUWY+gn2+0gLthws+zn8h4rjy7fHmzYTMBYWZYUJA7LWumDiC5sC+0+NqAhXL77f
WtpMIkT75rLdbqvr+ocmM2dI2rXDkjB+sWupjcH+oTxGJsv+uHcZRavTyN3iXLt3
SllknlwL/vUztNbXkBcy0wG0A1rlGh/MGpAOWwxDDgpby6oqv4NdPQbDVae5IUYS
FF42Asr8uqlDPg10wOt21+R9jHs230pjConyMcRQyP7iHUu7rQXdqLQIKeET/qoE
Kbl/vf5MNMAI2N449bqPabQ7+fs/9wJqf1GT7sHUc93V+uqTEOtgc/gn5mdlmm3N
FDXdN6VLEBGy8gR/xHGsWuDhnKGaZZwETdlhfMNJklcGOm+3oTkZylmeh6nESpKH
hYJqwJLKSTE4EBdpO0pg7MHZCXXKLxKS+iv3IogAnwjmiZcBfC73RIlUcn4EyAxl
D5Hx688ZCN52d4v95gIiRSU5eI+eYKscU8D6lElNOxP+cEr02R+aXze5M8itveY0
P5fGdnJvwpBJhfYwKv0Ikh6AwW6l+lZH9yRxbYLFK+N4vjLxTfPQ/dtt8wVa6G24
osTiv0LDL5ywUzM8cOk4adCljdzmwcbt1eWVUJNEA3w1apUN+B/agMmLFgw9mceH
0HUUF0nxWYXcAWGYEbphF5sZEkZ1kiEHPL5W/xhOF6J0Wg6bouz6m73+YBeWnxYr
dpRQBHK9nDKZYF+q0qeT7URfLyx8FVy0GH13LWO2b21EDum+TFXxTlb1sJ3U/GC7
HVK0QDsOeuoQKGrehCZWEcu5tsCOUoyscEhZAuV1xTRpxBt312b6n7HXG1HtFqjE
Vsahv9Z533EyMRYYT9lQW0Bj9VrmvmPaw8881kbQdEnRSJEtXOT565aAyM7PyzZy
gCFdkgVIul65cBZRm1E/+UYfQ6FPyFVOmGyEyfMj0RH/6CtlgKMe+J3Cic317EBu
VrrS4W4YIBbNzHV+bz+W1wjj5FKZ7BTh3TAU1PfGh1kgE7T59Tz9X2fc3AhYIgxL
Tx3AEDetFk5LAucEt1JpZtAKtrdbcmxcHzAFgwje+j5CXQCuoqpAS4lTe/PzEy3G
hPxENqBEZkvXYrXeFkuSTcvw3eKHPwNrDRn7qjmpju6edjKIKhotnvfWX2kuzDVB
eJWBUOyg2dvWNVwYcotZCtU5N+Byg4v12AKxp8c3HYvZveRk091zLmnmwJXSvWHu
jEYJIRSOe/oF358dNpoGm2cI++7ktPKhgaCU1a3jIcfUJBDfCbBVUmwy6RG73fKI
NOWJQLzQoKxS4Y82HM2Qhv4dqqmLM53O+5J5bKtBo+rQOSZpzlrDXr3tEZNxo9cs
Rjo6xtS2Y0176pS9z/rcg043nSLty2uV3YJG1+MPBktfuDh1+3u7qBtlwElufQ5x
kBYCrGs5WaHdNUpkjcsJbXqD67SWN4d2l3FUVBuw2ND0c0QfXw3QISziICAjc1hW
/zDDM9dSaK08n5KMSt4a6Z+vlDhT5oO9r8Wz8JqjJIFfeUP6H4AQM1QIQ/y5k1il
XjIwPfy+gzom4AFLx6XzdCPmAxroRUM0r6VHT7Ae1gsRkNBmjK1VbIt9SO0OKdRJ
wBz/vjNicq040VUuQKKT1ds/luX2ZgyQ9k5hXCGUmoREeiF29DkMTIMyb+fZaaVT
J67XxwWSP2E7msiBjme5E+I7mMVDPtKQFmoT8s0MrRHY2dw3KH3zLyPICSbhu4YK
vvN4prNkvV+tAPKgslbu/JVoeYRz/LyhxQtcwviqDP7Qg8T69sPUcaFquWPz4uwO
FWLpXRPq208Kw0T5kXYw8ha2ODAkHuhAqS+ATO7d3SOZtTrf3+H5FYw5OQZTSMlL
KxLH3h8Dbqna4sYcEK59s2Zmqea18X49xtfci8WuNi1kCKiA447lhZOjlbzEKdfR
dUj11uh+nA0yiZODODB20fpm2edOSgzdEQWHNBPXB/OgrCy7PEnJWkxXwnzc/AL3
NPJRHb0IDeqX8ON7Ihlx3JNHtelzajAmpkroOj8/j82gpyn2VF8u0nbrIXtZUUAh
wE2JClTx5/OiDGGRV46qwAP6CQMx0620XqozXCWBGMFRYg/nwavMy/zhAtA8PsZc
NCbX73DcKJAybQFP7PEFSBlcNVunr1AjdNQsbfT6BfRVU+iujTokKPhvEbJRQ0vy
r5OZIma0xwOmKQy4NkdsLGuhJMpRN0jOrqfm0+E3O4elYkRre56+fu7osQpF9P0K
yLXIOd+aMXRg16uwWurHbl/+XKycm7ZmKWH7HYqB51twBpnw1jbokwmbVV8uTlcg
IgU5WrvOrnzOhhScjrFdggPcmNaoXn5Qa4VIGxtrGJh0SbAD78glx1ut/3j8M5Lz
ksaJCx9McBshvbwwVJ9g7NcKqkHJmy2gUuePgTRItp2vrramDYD13eO6y/d6E6q/
34ydLXHbqzOpylNRzKbbmOndx+Y1p1FGmN4OiLI6eb//c2tU2GUXI1Kt6RbfLAN1
5A7YoB6/DKIvJ6cSbGJRAGeA4UoRximqEbgtU5q9SAQ9+jtimdKumSRSzz3ZxBba
JtiM7AtrejfBy5/vLkZg/UTUhzLbFxRHePyMHDULJ5daBj0J03/wGp9gMiMNXA1H
ptLbuSCeJ38sKVRN0i9OihWqSa1mhNahHN6AHnhfPcx+mKNYpDOdJ1rlyJdgEOru
RQRp8/nJ3JR+d9sMVg1nsIO1ZnPTuVkcTbhBC/e/6NeOagkXvr1kd/vez4xvUiu7
jgKaDb1tP6gNUEcR+tqX+mrU7RoSgn19b1rWCrdu3l24eWFIqW7Oc1zIGNxO4IhO
54oy4Zn7ftjBN636OND+7vVP20gqq1ne7jNPr50HnQaD4Yt7oDG6HYFGB96a0Wab
xbwpcq6TAscu5LsgOFRnfikRM8jV3FFUV6lrP2RR23skEJJBS/uPsdo0LLOkagT+
KLdt/Ay82URPM3g5hlcX7kZ1kbNuLgwqOPVSSTT1Ayh9sNj1G/ZN+84YgHhkifZj
5wKwaOIB4wTe5Q7jvmwx9+jCMRRZoQ+yphI/Mo7gCVRbvJoRntvsOv9V+gYIXe0e
1wlPWZMnz1dXjmc5kgXpzuyRZo0h4Vb53LBx/g9oDG5xZKOj47pJWBKWXfv+ibPN
6Sd8TVmmwrAtWylsWH/LmqyfghyhHMvZ3y1CQOfifjdhyHBoAN2mpWxfLhNOtSIw
EbukJNmTdQ8ocEkjBXLRUUdYQQQGCzbbFyJ/YOjc9DwfKuaeGHlJtosH9YxI7/8L
yVVUvWp7ORyCS63wivMrj3TxFrHyqGxYwgP/ZlJCb8k5+CLQvWeLjt8csv98jtpU
xxRcGrLdv1awUs1H2eQYsMshBedqLVFZYYIZtmRbWlbMvZ2EJJ8f54v5Y8DtbSvv
OMBMWwY0yrXmOrnLZKhUKiDZx/1SytD9SLX/33O7ijYEhN23b1XrJD8VBa6fdzM0
kfoShHGvrs9WPD6XCawcJG6/iNiHEteex+SBCMQ5XCygRmSQ9RuJxb6iU1F/Y9Eu
Tsmi3cA42m4kIJXe/CTPAr9R5hK1qqWWkZUidVe89zBjjo7609ng6ufCM55sC3+f
6+8OG+2ROyJoamsK5c4RQhchpcFnJ6+QyNosunEi4hK/5xUC4U/4XZXaBTUW4OpZ
Se/ArnC8bNr6+h6CQq9+IzA0PJjabbBOT3fhgoE0KGYMnBlLNOn/gos9UjsxcbaD
V+cXPX2aI5DWEndSimv2GuBJlO9GK+/bQOtaI5lBUTZJxxqEtCNp8+u9P4lHK9aO
Ujrw4elxs2jlywRINhaP85AhV8Sqw5eDIagEUAKqMwiQohqqGFdno0Eg9vUgopkk
huBqU2hi6hqfjN9q3iP16t/qbK4uO8lYfB9TgIBA34kSfP5ef1j0aQGQxbMpP6XR
a2Nw6Wr8C2Epd86Hb66Tl8H3BAxd/JnqQNHF0QLuGj8mh5CmkwX8eKmSn8Mr3GHx
MFB/Ov3f94YeasW4s2Z1iglSXUxTlMpDT9B8Tt0GrqNRvKBJMVwJqAMyZgMepmcc
97nDom+9yXKbh9uBq+Rc9qP7rAR1HbntDLB0eUm4/EYsfMe4cu/wpsk9oceOh1mo
tqFeMBK+z8CXMnyEHNzjgiOg1XdCbB2PKyVg9OYRlNGOrCb9fZyGOdVaO+p41z5m
fXtmUk46WJbpNuhGQ9n3EQ2cVbPvsi4BOFgZqx+I5hwVOKdp4lAbiX5SzosDPX23
CCMGIHbyR+1Py2uya+IrQQKoKb/7ZEbhRYWomsY5lr+ytUxyFgpcK/2jTdBTmXLz
mZnEuDYsZQAk0Z9eIw0MUcT2S9YrIu3yHGULNTwEN6ZOI9x4F1JRxvef2UeYSxkS
Dt+sUAy6YISFMkPLhFzYXPqdke3Gyx/+BO5YCgaxCTldoOczTxxLZj70iwZHQr/F
b1MJXv8YLywb/MlCalfPSeE2yeC3A/rM10CqtjDPJED7nIBFGJ4wCxtOUbdwDjoB
+PbnVgbYIsyQgliQrDTREMjOh6LCBmAUOg4K/3j/Kt/G8Qc09KqCpVUAXI1YKAQ+
WuskBEBrnlMuKVMXoJlyKtegFjHaEkZhHv8TlhK7uN+E5AOCXuv7vPTBszV03hwh
P8dRr4vIRyQq7M2KYQWJDbzX3D6mFBq1Aj55l0jMbeqEKt97zdAfMwurjysygQRm
hygACgw5BBFc4d/osigDZT+WBKshiGwHfZ3jPGMR8i0LAR4JOg/nvjnIrBB5LueJ
ZtAmUGnXNUAKj2oic8JUbN6LyDfhzzDwmJ/8rNRucZYXeD/YLt3SLcchlyPcD2mo
sFVhd3W89+nlEa/43zIS55TpFu82DOqslrDTnS8U3K8GITt/BcP2ER5fV86JE1rI
AILoN6O/8qaXp8tJBnYy2/roP48PknjOznOmx6cB0cFQ+0QQLHqZ2BhpzQaHxYpf
lWRFxzK1XEmPqz4XrGZIVqDp3mv7z0gnHkqMQjEuj7PZtKvy9Tl+AurMMVYDsWo1
G9vbKcqzXrwezaC0N3MsRzeFdeXI/tXv4u2BAD+ESpnZl0jZFoJy8VHi9esUXUZg
hoy62D38Zm2RqvUjq/BX+NSV4dzikO/uvoO3eLNMOhON0CW8YH5NntSrD2j3hHsk
kI8/S4I4qb0AyM4r5KpryHhHWX1htx1kgdaPqtKpykzlpuMawP3CvLqsVDQInM2l
kw1n2rpiuNzV48zbTpUFBXW55e4+17+4HwePt7bWf9TiGlJaIHAg5X5keY8k3f20
zSxarUCqYHVEQsWG2+IIoCuFjoU5QE8lNd/kMwT4kDfv418wlZmJcC3OdgGqzAJV
MZgbGDtbLYygmr0XszMl3IWycI4Gzla3R5qRPgOeLHFyISNVR/9SV5K1x6+Da2oW
sz9DWmNZOBfnuTwa41Ys3Xg94ov0guhPoHdhkAdbQnsplTXy4fs2IF9z3+FRa7AD
xagm0xs+rSdHYg5C7c5UlupvAzauyzLIazG//blXFMwBW1uau51h5uMp3Rw2gSnO
+VmyRxzq7iXuqP2RcfVrw9IYk674ARvhvmSkfPIm3BkYhkyY7tlUL0NsDOQxKe2M
BAZN+wcYZfdzDTBLXg2tLgjRp4GOmFnRD75tXUFMj2Jv8nnf1az5GrnQskr+mTWw
Qs0VRn69FaAlZUpwGoEoWZZM+UNzTjgA+tm0MCx4Ty5K7mmVd1WqZjy5JL7TB7v3
xidmseUWip7J7Z/tpfb+4Nafuk0VE+lf8Ll0enFzBQZMzLZ6slTCGo0mQbekNGep
09Xpb41RLPw+SC358x3nKvgnN7xB2idNwDAS6Fx1YfgwjYorFFPsEE9+QN+XWAwG
9i4ntUI4bbY3ar1/yfIpHMfBawUkxwUcYZk+ep2l73oo2/idhu6BsK6Nz2uMt/0u
5U89cDgFjsUsE2Hve06R/lpiXeFAtqJPrzuGFAr6tyORBM3Rh5TUuMMk7H+/yjkM
EVxlrLkXbhS4D3fJEFd3ByRp+nCErLB/uL92/tnmBY1CDdxu+Xl2Y06UTSbg6owM
2CtAlGNlg/ArI8UeqB17Q5KFbrKlQFXGB2aEaEXl6cEPM9TZC7R1SJLoZb7JDdVy
EGgliRWH8mZM93b8AbPr5hFxOAdRvjtDKyyWH6bIwFqzC7X8SNLkkWueuaaC5jjF
tMkT1ZTk89dsHigycg3gC9vdIxtgfz8DT7564PQebXsjGTUSlplUARy5FCvhjzsk
SWMSJ+fGcDrnEIB8/oxr7p8CnpYetVuXNZFkLKwIcyUxNWwuM3CJmWHukwejAxyI
JKXUbHyXxeCXp5q06qBO0yaud7hM7VWrL97t46mcs3rYR2zFSD9QSlPi/xH5Y/cA
bXB8CyRv1NKklbK582wi0JFYyy3VuRbldCjyVOcdWrQpvUvb/DJQlhvqTP/VCznG
0OJsx4kHfa6hgVJ2a86/HehW7O1xr9xb9my83zT9uNfyW92QvJccbfe9DExzd4xv
U6eR8eXMA785auw6Oehr5mNMrmfsRyfcZqHaA/XrjZTEPbTAOqXN1f3PgBGlS0+5
b/PADqSD9zNZccmfjl+epygf+CmIGmWUlUJmLhf03lpdRlnQOvncZ49ccRgfeuar
XvyFzGlzJPmHCrUfu/0JVJvgYwXWfsZ0X62eyOLufIWAnyQJQvbgL5Wj2v7ggpxT
Qp5EqFQEc9oVnSQdxoA3MDdvVuIYzPjNMozZaepGsnoLclfxLZQ2ZdgrLQp/gJzY
7bZZyAMTdoEWQvb3yhIkOpiOyjpCV7Zv2qnTDQXKAeiQfCCP1eW3YmWQEXKhwvre
Bul32oCmlL11Z07k4nVJnF9S2ujHyheiSDeZPIZoWpc858sYs9R6eqGQ9+s4yUED
61ob35EhH2Yj0xXFDh3+qGCLWuhK7iD8TV7IV6quClQ3yb7CgfYeLBKONEAp9EOu
O/j/UyWaAWumnFYR3OUEKbcHXtZ6wv/vLxm+nEZPeIjG/U8tQ2jInqmF3fTFTUZW
DDNUlcV1hgAoKcY6EccrEobUxucQSxQLeyVlJt7weUUNgk+hTvPGOUeC//L80YGG
gvDSmP4Fg2o2u9AGDW3uJEOJyCjsCgkY2Lc9LVI0k/xgvMRgic9aGLYehcjx2yjS
vHyuveQRSP8ySJNLyDG/1JoAAopdzqbHo0JY7VfJJK7+Q7mfVLnkNQ9O88t9H1QX
TFZJqCk9/hCngSt8W2jk4ocTk194bjTwOn7BIagvRtJ++kdGd6/RRDsiCDiZNrLk
zSlr8BsGdfz/PPvYey1n7A2FRbsWyII5Wi4QYYYipWFzQOWGNKLeZ8Z+KscYjxSY
HNzxdPaHXb2K7pNy3SOmBJfqeeBV1XjASMqwyTci3l8/Ov96g4MvgpWi1VIZyLdm
NRman9v4hAZm/M0McsaokjBaCRp7iggCoRboXYFgd5Hc3Uo+RrTFygEgGlV064/o
CkhPkBXeSgseMYmCR09O/BraRDfLcLwOcEJAG/zsk/CA/xUpFYMMStThqAgsL6cI
+EW58q3M07j3oIXn35Z76Gq5KJFR0sdRej+8Z8xfM4pPd3hQEi46bOHOK6XHEE0Q
QP2vxQt1E5JrZbTfk4lLOz2Xgb3sTH8z73spy7YInSStMBPxgk6+Tx+pJW1WAKvH
Kfza8gipK8ZUEpqdOvDpRmZ22dvLWCHLvDI7kMLoOYqc0aAaucr6IwRVBOdnSPf/
s6jROV7CmgPN1mn8enLXjCaaKH1LSGRio+KDRRChOEq7gxQbdkkl4ss3ptob274k
HSpYwYyOh3FLaeSG+ET31EIW1NwD8mB/5H1mH10rEKYjGmj24CRLRy8A9PNaVITV
R3cjAT+a0uR1K3g6WZv9hjpWLDgKW8vt4wG97M7BH+40/X59Ue9vZBFEUQed3vua
lSYWttxZE2FHgzcq47J5GRfsgWrBcnSxMEN9Fijovg+O0CR/lG1lcvxlnBkpesu3
ExcNmM8kuOHut0MpuoIMtVr6qG/YOh96Kr/cqlb8meS7DKRrSnNe+qPMYteNdaRS
95iOoh3WGdiiovCSAOr/M8ARMSpQeJpPXMm/oEjwsUfTvgghYva0rvhcGyCDc5i5
gtWp75lerFS4WS0KmeLbnhwwJYSUX0FmXA/XJUpSXeMOz9kbgtng/E+cdPBHBe0O
Ja5r/uP1AUZyxAFkO7Nm/2cB4v7lex1jm4idNv9QbNIu/jcMt8A2CYQczFrfnvZC
MavgAyrTbRpH5LJvTNMv3IB/3KbNTb0z8HSOJNC8J/LVMv+IWjukNB/Q1RnSIKF0
KehlQ5ssQSLtxRmXaM5k6Fps7mgKCQxWZA6blsuFxTKSYHR2+nx8htvCt3yt5Cw5
vdSYTr3OoQxUXJxzj6pQn2jLwhOikILBbN0aO3ZhXxerSjxageCk3KoMNGGhsAMM
bzAEfnOiAJvIc3/itI4Wp4+8Qdzx3YjElu4aeMaNtMY2gDFUr0Tp64Zca1inBq11
tjcXO1CKF3LZYDYYYOvGmhQEwFUMGKNE0sih8bOGb/fpKYlXvFUMiWDSk4udhW3W
f0KXQ4LerNdcAn0eVUWQ4djVi9SN4A3fZFgbNewtcsZ84BkkiZib42jxSa32waDt
p3vJgl15plumEOSdMoZjbJFD9Gsvif5f+HqZH9YEpxxhqH+y2n8AqWpNWRMNk9yW
2uh6/pDtFGcFTkUcMDZuj2eqfeBTmzXf/iBbXp3+HLOtJsuauPeSSCWggW3bORXd
e8tm56WpZMdhEeYpe7iYsUo/9SfMrY3a/I24ZaMG/UrjzgATl2tQ6BBjmmuaVHxw
uWFTnLFsThqkuVEF8hUYXKa+G40+Xl6QTZ061ZzWvkBBXmXmhvwNg8mERb06vSTf
ZCww/6/equx0voCYQcOjNuxHwcMnQ8S1O2ALZVMy3lHt4Wni100FxtTJdZHwAHlQ
e60i314YVuot3a3q9tnrzbtCm555o8PGgZwbMJMarNOuYYhlPUKG24kIHLr6K8hc
GELj8i4bQszq+OU80BTM0sH+iuXuveNAwlrxQ5b5SWPAPPzCqumVQDHkfGM0qN4v
1uPA4wdue61OFgPIMJfyxg3qQiQL45XLYVH44r+1kaMvnVUoghreGgI++CTfhhnM
zu1iGdF2PreHYt1KozPSJYVi2GpMYhQV8x/Ub+rPfFKpRmizlZsqSDQj/HaZ0i+o
mEbESRb8g6ThDC1hsVXhHI04ty6rl7zmur9gPSj84uajsNQcDzXjEa9e7qhbSOPp
1e6q20K0oaZyAwueZ60DYeFmcO19SzdArmMrBhuZt08fJst57QesucsUry93OY2d
Kdr3F4BkmO4WrEX13g02yhM6isfFLeYWS7V44UjDiTlQTd9wwB1wZL/ZouoA89Sb
MkJuxPFQHd757Fmz+m5YKJsA7eK3xJ0NF2NnzSRax4CuApnlrRYYHwi3TWMm7o0T
KR/+P//stVrACZfzhh64Vh4PR60wzszod5j8EpFOOhpUlgs/2jniOS9WxVVZvwpN
pGEhTC+VAPzzlYrBLeZBCwsa9bqZm9R614cSd9EX8J9YOqFnISvgL0j52vLIUIpu
JfqnPsh+xZYBwDKdi5iderBLgR8C+EsHpYX73ie63cQSFt4lAe2fSuZ4GWPfKIum
O1gbrJ8buZjNrXSAAc3oN9SuD3LNZmmH6O9MD9l4FagOVFCdaqPuUqTysAmcxWBk
opm42OL7ZNR/TfnxHuME5YoMBgdHPbfvsVm+zSUlk94aNpB4yjSMOnuiTZUOq6nE
DLb3GgfIKipJ9dt1jnVobPjnWPYZ/IGH99kQsR8EbiGAirJeSUCQM9N/43PKAIPM
43uuMhDtPhAe0y+4HtymL/T5jAXSwA3J39YYjH+oJdIbJ9ebwIgA1WdNRWxSSUWv
auARSoVODtlf828fPZIe0XLYddxPNfL6ArX2NTqfzLAU1KT6uEyTHa0IAGbBVlC8
5pBYAHk0zia9RYn8aY5UJnLeo22QZ603QJzYXji1u3gzbj97aOxR5226K9/UpaXV
mRMqXyFyFbQt0s2Np9PrCuj8vxDqxiLy4YQxFIhxVBefIefjV4XVfgh23EU7S3W6
Hj2fTutRyvp0qmaDkmbSfKBXbKmk3wLwZjjNXY9mAWCj6pEeUcIfJU0WGIstjDLn
vUTr0HtS3D3f3e0gDh7DwVPh0/7sS3vJsYLI6A7S8B1/IYzTulhz8PmG8hpkKAPY
crJXDfV2ccarDRE1PLQA9UjL7+8GeZmryWl4Wm1Ay46SE5zGI8+q5D8c4/9NYcQm
qS9nXdWj/5YNF7V0f3hzyVgSJXQpBW4mfvjS4eHFklAeXwY2Ru2sLKOf218NHNWC
p6o78phHp7reefkG9/l0coVh5NC46kG2ppdnRlP7u2+3JZjGn5gO+0R61njAA6xv
MIvn2bd54MWd/EDeopGgWcRDjMaC/8IHjwJ9IbE16d5T7gh7CqQW4CH3mdd5Osr9
x4xc3ZP6/HWx37MeoVJgrMtVnleu7oYsYjD6WTV+XeHRCm+DfmI8NCzKzRWw5jV8
kMfHI4XJJ/CJa8X86wn3sMVje0BTfy39YmmQLl1Mo7uIeySFlnWnK5NGlg+r3gEG
ap4rl4opA+6lccQHxcsMf3BwS7j8D7bXNpeP3C/v52ucFVrGiQMaIhnQrus1b/9W
PZSQbqrX6yi+Q0xFFmp2gRYC2gZCJI2jJxNuDl+RF0vuFMVRtO0KtOpAezp1TYlw
D/1EoEBIGXMYdvHz4VmODlaLSd/kkzuoA8wKM8RSHVzTYLayZZjSGYHmCB0DLyGY
B4y7OAbJRjiKv7/1NFad1TEhYGo35B+O0JSTUmsUZM5E4nby8EhchMSTUmeO0X0I
11vZi2YFMizLwV7dM2l3rAjoGz4NmuE9HggPerT1XUeCvALxjAqlT03p0tpUCY2Z
jb8LeWVFtEmKX+OgdRHoCGesi0QODDxcZ6WOjAENKhnBinqsJ7Ta/fW/mor/GTSQ
f3GcKE7AFaypEpTOzemv5mtOVPwa2wi4TdmsG0ozA3a60xFNRSjEi+x5ZShe4fzj
Luxx3AOOVJ+Vt/fKeG/T2qfAyB3AlXdjnzKSK8XqNCdU2hWInG+7i9TA139vO1Z1
GvkeASFRke40tqfJxQI8DtkYpGhpNdoHF725xMLcDamkfKGp838ExQcVpqvzk+fD
tZ1iJg2pbjohnyPLTRHOUKBpHL6d1egwgjyLz9PXB1F4BbjC1HPFxm0iLjQhVbaR
urYj0cysS1/gBcxdBLNqB62eG/J4Zq0ty+PYWW9ZuoSJhMgUZxm0LLAMDgTnvAm7
hrnFdTOY7wH42AMGN6Wwd7wVjteJBGReKYX3vQKWbUXPmj80IGcL/+9WetF26OgX
P7XL6ahKFiieFBBLt76acQqSQXiSE1rREvjKVPOus20l4l12Vr/fr/6G/scPav7v
7xwgu5EjBhFOiAIe0H7qfQjrhkf1X1HhISG3sp1KIE8ODgnk7Gcq25YSKIc1h//W
H0lVYDXPJu8E2MKlaoaDQK0RYgJTcyhSp3hU9++jr8rHnZxwHLVZtLmKPvJb74Tu
G2tGQOJRJjKtbFNCsLG+Nuqcf+fSrX0PioUEPrHAme56nfJ1V67efPnV28SexNtc
7Gg9u0T895fGq2v7CM6b49Ofe/oeIUT9gKj76QF8Pv+LZ+s79zKxAJvrNo07+J6s
otns6OgOdF9nPwUJdE/OPinUZ6W03svp/MnGvDtA8ClV50mC6nhDyUkYnFZJMtVx
l4h7HvUvw4YIVFRddBMT/JZLhJ2sMy57vHf3zuzVvS1Psim9/ru5MCGrHYPet025
94scyfovNvfdJaaI2AqTWHpcPfDRcScqRTb96TeijhCO/FO2XbHLrENqIpQ9Cuxr
tAdmWqvKdV2b1OzYaTclLvSjfW6PaAKn49PzpG7acJ/kpHDjb+5WMv9LiTxjJMCz
kCZKxrsar8W0e4rYHXo/RhACp740YObQVl71WJOWR7T+28sWV6ecomsq+bLTQM2o
q27j7KUIlpaWwZ0RHk1Wk3OT5ATDBmXeNI/uBBk4Ev5BSzouiUttePGw514ucrhF
rCoT38tebA0ntvezH/DGHO1kpbbBx6OKDHiDRuJfWIFxOpy4QDagUBe5aRA3TScT
GeY6+OI84VqeDJOAqPcNKD6BhNtE1WtmBTNrCNqpZ1fVvgLo3PsJZiqzn/JhL8BV
EDGsAD4DQ09VAwfliZ642V0W4N8SiNN9wP2iXwo2ug/7fHtLUNdeoWCQKnzTrJ7h
3R+SlvSfguJQHSwAlmHCdtvq9xQJ73cPlN+/Af5+nNTgehQURSWQZGxcwANiKKrB
wp3CRbqHxdpAmHrjpm7s38W7DWpU+HZ1O/iQU5tY45BRVpvav5uuESkY9iGXb1iL
tt2CdbZBkGmgXalfa+KJdV+gYi2lIXS64N5IlkRGoJL0/OmaIXcXwSz0ngo4JYX+
y/SUrYI2FDwK4nO9v5q1Q5njHkUvs2OAsmPQ7faepiFOQ1VeyjJO0jGS8pJ3owuY
n14lnJaEF/74khAm7mqDgKKG5S8NjjMhQY6rTeN9DQ6qunNfcY0R1bGXzVgSUZ5/
qh7VA5puIqHleE6XzF0S9mGbpp4+rGdDxpczXVCxKMFRaWsPabGDeyzhUI+yaTrD
tsOXhVHadhLyNDAnxkYrbl/b2ggo88GPScN4PYxa/bU+i4VUqxfRG4MODXJjHTKP
gKo6QOo3ghpkasDSadxGmwOP9CKsANIa/Aj/Qwqr5Nb755LT0gk2uCyJq8zpwo1k
D+vaciWrLct3dp39nCOOQJ/zDtXl1p7sS7Zk2KFWs3hmY1RJcXB8zYnXeYRfqKGO
B9YVShFGFbN341yIxHvOooashnWHBxnBk7n4fo1RRBc02FqD2sdZMneupR5qqGQt
InO23rwsIyLmTLcWvpMDltFovZ3IydTaTyEu3G6GOjAflX6yWVsHf8LSJAlJPRvC
vvGjxnWNGs4g1q6UrDtPFlqs6UXR05Nlm2iCtGb3oMaY9yViJ+JB3Wp6/ZmT9/eA
L522YbNiDo2QOo9/cSHk23TjKTq79G/A2zs8y6Oml+ixDaSPfp8Q0ss3AxBNf1dU
b5v8dq1UMtoXGwbXDULlLst0lX1GMS3LS+iQVqG+PV55Y69RWn4p5WpcD/kKCF6q
Cz+NzCsCwHLoqEtAsThA4xcFdPQx50XuL1gcQmS8oeskRSBFJuaatZlQ4gA1JolB
Ng6QPwSK/BO4APMXmEz8Tyr1wrWU+vZ2k+S23JW1geaWrQIsV/Udypp8myruZUKA
g90RHHsSgC1QAPCNb3U20+1xeMKzeqcIxrBpzjMiTtEzEBvKfXnSPNTKGEALyvgG
zo6vJlTpr73RS+N9qRu1ZTEgGpVGVw0lVLOzMT5uy0QTxjoGr16sKo48tXOE21Hp
sueqgtw7KaEV+uwi2Rb6QSoOTm8LIoWK/1OpYRaEzPkJeLpQuhPRtqyDPEGY1H71
gY4J4Q32F0taJ8g2ZxS8rcUv50ztKuU492FUs+c18+ijnkfqc6nzMnlBoYWXCaBO
vjBVaVL5Rw9JJqUVUlv6j3J6e9qaz3/sArzn49m7ZOhkKttVn1p91GwklJlLHocQ
N1u0s9us5zHccMnKG2PmTxPvNWNBp5mQdTr2sKXDAAQPTUHfqPNCPaUfH6oOy2y2
TU3oar5IcvaZ8PKX38NJkNdcKTofR/8u8t+6St6/sTjzFYGleR1RifoHsUVyzjqA
fHLKrNnXdxq4b1AJPEQRwsQWClqRbZa/FuUttcbIbSl7WM6oGtK0flRVJIHjp62J
Qi+L7MgtUtoldLdgpnOhuQb3sQm30m/3xTneIpAvaPrNX62q+ivCFPQA9jn5nThd
hdj/XF+DC/f3tKq/IbwAPR3U9DulAIfxuNcmUEgb96wPBITkqSKOUN5V5OyJGKAi
ns6xsI8npOJIOeVSiyg02ueIcPsRLiWNEpysZp5Na7Vv6ewsfm7Gj1lnBNZkSZaJ
vs9J4piLYgY/Lr8Pbn0bcXwJglzQn+oA6axDXSMh3gM2Wwt28h8RsRRyHi79GpTA
DSb9QgMFv35LdPCwpzaeljbdW/L8Jv0yn0yrqCtkCosyUdAa+9Wvo+FabFQlpT0l
RyyiyuqWMGmvFyv4u+0eRsCvzujnKw1oEvJClyGE8mjcvqF1q6+Yt2wyNgvmQxvH
/54eaDpfYqwe1232gWu0oy9EDVMS9JldU+xj6Gu3vV5cb78MUIDoLgQrDdbRxj1K
SCCkCJqCfxgUjR0am4MgHtX74367BCpdXfV5+ABvFiRGnLicCpfUzp1sdIRqbmoD
9HrVimYMZCep+PNFdBapl6TqIdVJDZ7nsfAdzbdmIObShLP5mWSVnz7pmmE3XmCc
zb+LVSkARra2EOxSJhyahb10MZ1Vc2Ez6YD53g0pTiFtK9Wx7zJWz9qFTbyv3IP6
7hbFzfpDIaCpk92cbIQCeYekAOz6MUbpkZAmc7WzRXWtcGZVzYRNIADb4nJT9/6C
yu5vxeuBxHWeh2d5u1vvl/8EvqNVRY6F45BmC2G5StxdZI/RJC+jw+8BKVn4w+5b
7GVJxhWcCDjnghrvNsIDwl6x9P/pqxcUi/TBlFLFZ1DmZabAJ/tua6Ko+GT+TuEb
vXS/1rVGOz6pidpS/oCKA7KEUuoVMoKQqH1L4R3ErGvtZsbmKC5SKFUZepOqdEtP
LYEVrYOSqe8IviZkG2VRKPfJ7tO6X9j0aEurKaygMxqBnoz72S04u1+Ko96f1Lyx
qJYDFksNo4drlGOhEfgoaA4C2xyAI1YCDFkM8ZBsockXc4rQOscCVu5AuGEZm4GS
x99/i4QFxEjtwUyIEOfgVPeqFrhX50pZnsHpTsGi63oMywYkq2n7/pspVHL+sOhv
I7sOTWe7f5/Zk+uUesnI5aJCpbGLjbSEp30f63G1d5p2pcH1tb2lQYUfEl3m6hfv
685mlD7Q6lZrm08I9CByQkdo1bV1tooGDJjIVSPVHn5GGKqVNLtbJuXAWUswSczl
u7NHPbd14zdHco72uLOocNXa7EOv8LMsyk2IdPV3qJ2VJfi0MzKB6hGbxkaP8ky+
s4j5v4GPAMCt6eZhcLV8pSE2IyV03Qm/SddCOZr/pEkBd/pKof7TDEJli9nl5LwY
cwEkd9Hu1stfzXsCnfGN14eOl+SWnWmgBo1k+4SH7WnXKtgpWM9t37M94LutJhWp
9ek7qx5YLO57S24PS8Jn1pINF1JyDHajNAh+Evkg72RZ2c0Tq+wdT//qd+RZfl5l
rZ3zmSHbnJszIPuCPBD3131lltNR3uHi/ScaMcgo6vCD5Hfcc8B5p36DN3ufrin7
SgYgdpd4zB88IP3iZtLvtunitSv9slok4uJuXA51bLK3WZ73H+O6i+PszXBS2Cao
X+raO+nfkhCnhG8sUVZLpOFQ+IEUkGe/ZPqB106UKL0tMlMo3bfpRI9nHtjN6PBo
Lv4m91ZHZ6if2PLpfd4LnL7k0eiSB0FyIod4YalQA68pmYOh4VqKz9dmYcdbuxGU
J/3EnR7rrR1oLyZrtzxqrN30npf2eI5MEul5CVl6nLChY5qcH6sgpvQ1UShHN0RW
cam80vE3f3nFo+cx0Vd4/wRCJizvuukGP8ErakPGbvXrP+Ig8Nm5RbORLM0gP/Fn
Kz5+vQ0Q4JZCgbKGtJ07ZrRpp5xYx9fKxd8zABJCsx4ewE2dPlBLi6gxzPj1Ce8R
0ZRfOO9UKtyg7VDbznXLktf9Yxo/bw/VPm3PPCRvjVqjKVrYsxSulhQPti0yNeuj
cz3jT3TPbPeQ7wbENvdMmAFvT2hhR7hxNCVOyTNXqa3ykBx80cXNQ5qXIBjyusrh
Lns0fA+3Hl1q7K84L/9/ej/PgNNYw0164rrjoBHCRVfqx5JdGwtltnOGuJRGbUz4
qUc5+a9LP3FHzY9ip5l3q7Vl/p05WQc4NJSHWsozstENULDaTuRuQDA65gcBMmDd
u3zq1wDDj0DrCRctXONnniPf4SCnqz5BXR4JWbc/PZFCJBPuRA7hL9PP7S58tkyM
BO3ok15QHuhWW5n6qZ5x6mp2my7YEVv8KLGBsEeLPMZlByQTxYJzboN2aRzvygJF
mkxdJmn3HEkMtES7efjAXPGbBky5sstDuE+8rvD2jHyq2G6VlcFj1VgHeQifO4T2
iyfcMb/g+yrqQXnyTHFxm5+pcUjDQ/FVQdRmROEtsaC8txnqCs2HQw1qPln2OA4b
oVEEuAHvMohwq1Y/i6tebmC2FC+kokOHZL5bPY35/YGOaWmvJLrP3owX0nHBtTP/
bBq7iGpqgh7ZkOEt0sG/1R8GtFZWNIvEFeSvpYLUqnO59CFL+ae8Ugjxg+QXF/wP
2omChDbZfK0t7FuOYAVBQYNQJ9X5i9hdG23Le6Og/Wmta/tWiJit2p6htxHUSbyu
cxCuM0FXzPy4t1A4npDAlK/a3/ajYzmXX2wIVraUBfH0fN3SxTxK5ulZEp4z1Ac+
OLnNgfHwWt/k6/YMT1hZ691BrX3KMOdKAwWNw67lJmvkqrN4OS8suLM5VUqFuqNW
2skpsAonv3eSD0t+r3RrtY1d/1EQDdKUbUOgZHiQGykfj8VE16RHmagrpr2r7gkK
mY5xpGmAjKYb7Y+mggyCMxsrba4a+i+QT+9E3aCjCplsbjspmqNx2b/hnhqQRWk5
hXFdF5qsCPfPxgosumW44mPGn/67yqrrfwMhDOZlcSaRREieRVa+pmEHod0KAac5
9N52M42kyJNLGB4tQP1itfrZ4EekD56N7SWLERQYmTsPYEoosAUUiXHKL95ec0iw
LUmWp7AjDx+I4JM4IQSlEDLhSrI23RQQqMlI49KqjsGbphXqltNbqAbeQR87L59k
c+ngXco91nzddvj2yJ0IWxa7TxGhBQ9qd+4cCLtFnmPCa8o0E9wssY+4i7V/JKA+
KI/AaQS3cCFA9js2Joy1m7yfgqLhfrlxuPFBpIeG1MiJDbvKuf4MAAvkYRTK2xdq
A62vOne0ofx2M1DsVp8DYGPy9gLdGi0w3Zkw+IAjBKJ3NhvJltwkeVU122iJRRAZ
VEwp+tVRg9r7cSKEBtJV2U/I3Gbi0Huo2BN7Hcvo8ppp9rzSlTsLrScybUm8mL97
d/UM6CMjFRMbEwXNtTjM53jE4bttFgnUwOJEJnaUfsmWoVpCy+XYbyL0fv/mREhP
r9vdSIfXEXnOgMR1YnJcb2o7V0b2opeJx3FCEwt+WxupcvgOMzIQNNIeU1aO5LKq
Hi5OrAypYuLe7fGzvu5U5sZ/aq20ZyEVjAW/0SIJA6B/cu8xGOiTH4LQ+boghwoI
c42lUnKVI8lCQwPCN15hRReSDUH2CywdT6tm90I0W9/ll3o5r7+opBF1K5ySyp65
mrxAeNM0Pf2MyS1wpmGULUcrvyKvMpkDjRtRti8zCVW8w5Ji95Y1Z4vzj5keIM5B
LLIQj4/slMkTuYI66xblE0S30CaCaWQypZ7QtLfkjUi35vvKXuiwU4PSQmixQ2mA
ATFK6nHoP6WYcVJkPfWHOaTv3H0l1PhMN/2pEDcZwT22keWTOKsxJa/YfoJRg1Vn
uze1JzGCKmev9ZqjiqvKdt5PEIZAdZ0Hm/CFiu/XYNRCkoaZEhQjM9zZsblPO8ln
+/Wrq+7e/ap12zRZJQyacGFrRz+m2FV8NBYMukY0k6UD0tbCHAm/LtmoCliHIA3R
BrzL5FUzoqjh/Zw+YK0q9BqQLpNTWpLD29l66Tz5IfcOoBYHuTHChNAt69MErFjE
2DdErCg+JgbEpN9y5tmY6//0jdjHjTzItew6kGITYmXvhnjXg5r/oiz7YvPvJp6x
81FUZwEguzE518nSxX9lB6Vpd5HUJR+N7rflIL5ivVU6ZUeWBOCirTa4OzvCuzy1
MogAmge8BwZIeiXuXmm5wrxTd6RgG8n+UDATVaJsEknuJ2RBvWv1PS8Qt56TIetg
ES2Q6NqNifP4BdXhTWmjhYeG6EDqftSbz+kN6d8HgUvMyc0aUsbo9JF2o36rgRTB
OpCHlLVmLXoKYPrb6lBpsQz8+1wY0vkmPod6iMS/GPCaoH5dpvs9NjNYqXNft+v1
g/vEad5hgOjZNCmtYfob56A98nUZTSRRc6VBfdfnS1lY6U5mBp2ZB/G5C/rFdaeA
zaMcuSAcOf8PCyvMUx99TG1hDRlpBGFh6NYrxo0Yiery6TeFnhODHa/9jC0m6Tcn
fRS3lfrb0QK7EXf04QnCWyyrSjI4gKOV2yQtWJpC29sYWmW9gVikLRRs7M41pQLJ
xWqE/5Sz85pG373oc52jGU6GK2js9sqVLGsC0QbauEebyl9P82umuRtQMlJnY69o
w/BuzvSMz9nyokisKgXQkmTHmEkAqF02Usk+dqq9KlUZn5JMgJXcYoQoRigPCx+u
CLfXUBPgRnsaY7dJUWsYmZQdGaUxd5G5K71ghdonMbkLiASrBKzOCxhtevJa9N7w
nJbuDtW7n1DcDI05nZK9Jigm8n8pv2+0dPFe6zYxleIa2B/QCBcMGOlAhtzi+jdV
c3LGwvslOMoMZByivzHGBWEZ5dte3dw4lI6maLzU6l7BnisPnpgv301E3Tw3yZ3P
BQPhYHbJXVRSds38ZYqOnLzRDJrO6bktCwlV8tsdB5oqpAbVV5HFMC7KaEWQRDpN
huKcJIr59Sx+dMxBBFIEi2Zyd3hIiq0D65njK2epqFgb2Ve3BEw3kK2jGYFjLJ3+
P0JLdm/D4ALJujJLSa4RzILtnfCIVPnI8nL8YtXbA9JoTVKTji9QIGuzgEZjMBEh
IY4EKtAhMS1MWMogKAFNhjD2fwJ8UZrJvjvgTy5gSjA/6qxxJ904NjSuHAsgV/tA
fMjrEpfjrgRR2LYaIfKC9NnIOuUETN+BDtMJI0WrIuyaLAAb77z7t9jCHkDLLsFN
i83T6nXvFU5NYWObmCGh9hRpMFeJVjg9QsRm2BTV09wVHxOaz93rUjluB50ofteW
nhoo0QLytVpelAbZPA5Acu9bG6SQR3O0pA9mpYtSB153MHIRkBLCpr9xLbbth0MH
sLMmaIYMrfKdl8MyQSK+PGNb0zfcCPj/HsOYn92XHBdLRHVwMZQnuKzobOq9XOk/
h/LAHmB/dQD3V46JCikOfrnwuCjMdyoRzySjcuXplIJjkNySC4KWyjgDjZsx266j
l8pN22hM4WKRoB2wkuqrgre1/diDko6Jf39wTbqWTjTR1Z5EYmajQoJZBZHyL9bX
QrVCrq9z93Gjurstq0jBYKNSKPJPs/dw+wweC9t7LnijSMQsbMts0u/4A8PWoVTN
XgQEelECe5J3CS0/IH7Zpa/tt+5aBSHb1MFLHZPViKBWjfv/zD77Y4cMh8Gm7Tkt
iHODJoaRFH+JQfmMKn7yWnNeyxfcvN0IuineDrhqJtjCh8j8EaLJAVTJKH5S4aTY
bViOzssnRLdbbTTZcXzTKuIWPnJfEgxytwiqXtdOUvRBOKesoxL0XjAhaBM7C2o+
CAsai96xOat1U2c22yfzmy9h7EqnyiqTjjwtlC6qqprNZLFw2FLOTKGR8Cb1sVQ6
LZ5nwDocCVnDy9DqwblEIDSQwectU9271cfafoi0AckX92Ob8ChZLhNAPFZyvcHm
sEnYopZxp13wuTONF4v3beC0MJF5cRMOyxGw7NOQNh+nAHhqvSBqNHumCJwM7F85
OIU4sHr+UhvHcxwldmQ4iphsV6gxGmAfDZoO9jNGfgbQJ+YMcSHmQrgHWHDaYdgJ
EDdYzHBZD8v9ZIwnpd1ZHqsXOGshhGKhqY0g8CM/Qx+GHZP+EwCGND3t8x5oijnz
cd31viRApFYG9zH4CaLOlquHyeAju8ne01JNPJf90l0TdrV2k9k29OvfubVHcjyl
k1MrVKBGJSGCKxkNn/Up30I4vzhWkJHwUJJJsK5Me7W0KMTcMcOIcBxg+N0UBAyd
L78r0224z8t7cgt2l2ycQTKv9aCRMbyfOWtS6gqmi9nPFhnIHoqVDWcpZk+8EQr4
SLdZlK0i6kLH3e0IPsu4Zg+YdrWL+PWcJ849zdocjL0OrAMENrOdZj+//l0+nhAD
v/TJU/smlGdgsBldhOwLmdBgy+7RGFsMpSQoighJspKXyeEpRhnw9aIjjGSM/4fg
yqNYMt6y8EFGUctG26LxLR3VBCmM+vnnNTYXqYGrsaDL4ClPu2t7vRkZJMQQzb86
FCIWji7BcU/42+c/grglhOlNW7oOGiwKMFQuDaxRdLguzIKsY6bUNGVYJ+T6/jC6
Gif1ktAuVoilwEi+ONkYWa0sIG65Kfqt1FSwgdtCAKMLKxPUzvdY4oMKciNci8oz
WGQtKPumsAwPrXoozYt+dkyc6Zkr1QsiLM8c1VEnrciIIVhyeRTz+hni5iqqB5ET
4IUZ+J2yXN8z0riykBIQ/z6lI4nT2sM+erGaP0NeVHaGUdZJOCn6GK4HDeoCl646
/KbhV/DfqDzV4+wL5sOBPCj0sijxqfk4Q1W+UhJbCBHlnKVo3HY6tCLRVk7HaQnj
DZUeFkPh6Ug6Zj+w1bABhRAtOo/A+Q4hOkAuzntazwx2Yz5qTkQ0AnY4lADrB/e4
Z4gyiNv+pBGpXDMla4rV2Z8tfIVJCTJRNODuqc186+Lwyh+DTwLCQMTO4L69O/1d
0uuaAOWKb1Uzj4ccoNMgxEnN7BdZk9vyITT+mS3BsLm5nPtsbO03+rFO1hz8rbLi
Pli8jv1ap7rkQQWU6cYCsZSu651EDGKa91TX023YjgNY/RPr2cFbA6ponph5zhT8
F8SXUqHH6eafpCiyLz2/MCyL2KV85GqE/mc45HaEPjjXeD1O9W1Sgv4W4h2QjbiO
zSKSBrJqpM2PtQQB6La8ayPm6L3ujdK7b61WODjJwAwNr4vNCQ06rCtq4V1icPfY
W3uCHzBWDScsz6SiWQvGt0fVon45WMS856xMA0QdC8spI+AWkPdwVjN982CQBBT0
kaPbVCZuGBQ2NPj1f18QqEx5zHhvgt3Ec8ROxLhr1SVVAx5fcQPmjf3CErLk5Eeh
lDjDhYA7mKWJbaz6HBBd+RsDvsYpsrswsMatfgS0bDWFj0kInE0yDJl69uNaZtsE
Gl/Hb5I9E0lLev4SmBR2ODvPDMyDK3ZAYzA1XTQ8X96WVZcO+gYhDLYubmbDR9Tz
pU9XuFGMoDpHSMx3JUbhU0XvypBWmsAJ2iDKG1WUF65EUVcL+4pzRCU7P5WSSPO6
mkkf0QB/VVmavVvZT0x+eml0iV7mo/1XLMxJGujJ+GdUVFdzUyHY+rHQ1L51BhB2
fHsTuQtvNofibsLCOtN7aUbgyyPpTyQfekTV9sKKusN+ofqvkrEdolv4Ln6IliHI
N7scjrWlBN9gT0N64NCNQzxkVQqzOxPbbI4GGUZnh8Ytg1YU9hBFO+Jb4mLqoj57
Mu73bN48ZIWZzmxuXtQUrbO5ewPD622ddD4kIHP5XcWWtj+VOTvFqIZZl6fk63vN
p8UNDyMH8A6bzVoc8IRROGzoEXdIiEuJYbKMIzKZMHJbPYXrjExuCi4anl0/no7a
0eLPRufrC+qzgqL91X+yFIelMuhDChF4CUeDdG1q8SqhEDit1MsI9oowXBCbwOGc
wCvnxtkTgTxYwETsccKG43LX0OwcrJ8WWhUCBJJ72m0YEeQmIlvdCLFBoq8+bOfr
vPTMnf6OvdR8Dv9qtlerSDEWix1WkBHtVf5Ma3f53nDXaN79FPcLiUFxPusraYlK
eyWKbXDRCQdPFhYExFS3cQqCDZny0CmqD9L4hjbt4USQdWxYBWaS4lo1ajFWHVvd
ryMfXxxGCj3QynucMzkBu+pe4oCCuEGjhLTj0pz0vZWDjew3c37PEhrknGCk8WQR
NoPYisbM/X0Oj+MolpmJktVloDHBWVRRpCmuvuiiTgM3vmK8mDv6fQlIMNX11K3G
xXjWwHhImtt/A8ycyLJHncgkOnIz8TknfhNHp2Ed81A/PQHJd6i+1YFBHvba9Ont
ozwhc03eMXF2DEhPlTsTFJu6t9wTIy3KF39LEigG+eDi+P/JZa/r3cbyodWlGc1c
vORHsF7QrbBuwplkNkQnDAB8FaduKvHwv5g/vT2PK1PjkF4zix7g4v/O7miiK865
pBEb4iUI18ndMkYquyNpdVmsKFISuC9w1EtVWZr+5POhzqlLzl1s6r3aeFahH1Xa
XOrMEB/8M9o9q1j+BeDSJd1dtYODhlbhfz6X73b81QsPrrF/pdKO5n1nsYvzemXI
P33Lzyp344x35OS3kPG/EAesIC1dcBDrOwGfZeEWF80hS6crm7Zd81i5uAGCyQJt
GE2gMAf86XtoAi/ta2JPDzq0azIsnsAeZ9bZwspQLDrvupPXoe7xs9/OjCrqyqVF
KUYUGeZr9A/2HQE3et+VY8JB0PnKUzNCZbHNK6DkaKLU8BGDku5m2ClkqMImYKaB
JYSfPkhUZ2ovRsp8vufY2j/k06ArsZtz9DbruQ87jbg84+gZOuEujM/zu4/A9+cw
FiElf1ExwpZxbb0CXGGQoWcKV2MnwalhtMJy4Wgx3HJ+B/iDAJstN1B0g3Ocnapl
l38fK5HnKWcrXkO15IBpBjwh4YZy8Zlin5OQf2lOkM/8sskl5ShgpUPgpzCv7erY
kMILO+s8Ahs8AZCZ6TcrkHszykDNm17HfwTeP3WZqcELpkK+uMWqo1mdB32kz/kX
z6ToxR0X7Fo2ugFlqZDk00QUwOgkPTknvFjeaf4amvw84Hv9H9++gN1aXIsrJLmE
TDO/EZiY80yU2G8TmcLliVOeY2El+0pgkTSbC5EhuMTSMMXTaNYOV6uQFGKst066
J0ZIzA6KFSxo4y0XR5eAs4BEkMZn/ZZlvhyiIZzI006o/bCEznJZvmUNSjOIH4nR
eK1sWo2NdltE91ojU+5eWq4ya7UUf3uOu6oPtJBKXNLaUtcwHIMnWzldO2nokdFS
VUGQzyZZQtBHcbBUMx1d7+5qdUh8oZC/cVM13vKpTqUkYOA1Vo+/uCMrpvwe2obk
97mpoqMXYf/ESVVpIAQXsce5KosGMINbH6i6Ejxg310v1syde1q+v0CxpLqHPozD
bHy/XUUx/QYGlArkowa3xQYlZtXrNpbnbDyNPzArI40BKU6+F+48Os1hwO2U1AgP
t9CYbEUMtTC4fjixsH8u4EglGMa/MVSHDNTqzfAoOBL3aIk4DAbAFT9fP+R4uENk
UPd8l9usL3SNExmwHDRmES4qZ9fh/zApn1X6P3W34L+Pp/Npl0RQ2cOmej7xpwv5
sIXQmgbSDuRVA0pSQExVLQLibSaaFUlDhXPgOyb5IBg8aVR831ax3MmN+VpxMspR
qNF9QC13oXZUgHZCN01VpTeqgsNbr273PgUjsFATV7lPA6d13wWsd+gswun4TrIs
1jrqyjLvepmV60WxbxIMcHHdw/ELHvNz6lM5L3hQQhWKbYh/LbIW8i17BWqvWqEY
7oSsNpqdaq6CEhD2DTLN7MNPkKPHBFXxoL1LfL32sYR/pXGZIILno8jQkKVmWuXY
P7Fm/POv+Aya0TzIanoMFIdRoAQ72xVzIoZSan1RQaYy//DC/jlGxg8ZFaYnA5Iq
VeR6zIZkCA56LpjUAjum/tiRev2WaMDyGIJ+qY64KghZ5BpSCx7R9eZ65sxlIsSJ
hlgsudF4IrPRzFnRNtClLg1v40lbGF+SnvD+Vj/oy1e4pJkk9rWbydjk7A6daYG5
1BYw3XKFg9xqz8h0kIm8nGF1bp7ztPHhTg3JqyXsNMQx/PAoOLLHvoxjtP6XI13O
vmXkjaGOiQ5b1yCHlgikHilRktFiaHtqbDZRPJijhgVvcTeSQK6iTFy3PIFheSRW
oi3MvlUuGqlNrkSK6RI+/iOa3w/6VsFeN8TrYT6gtTOTvsGXvEv9g0UYP1o8Jz8B
XjLfP76UbF1mDdxZTqNlklhkIEUOb7yQ+eLvnvd4X06CtuMofZadigEKKVog4TY8
0X7kXbvJFHRxtJq73nI1NUMebK99+bcOT8WmpntguSTn2lkYv+Nl2AehDQThSru2
WjdoF4cg0LdzdrPgWvlbM7ipDnR1BOebSb7QHFe1M2Wa+GplxndEI2SbLkTlW2j2
jikD4bXhOmnJDmhcCCZQmTZa8q3fD+DBB/lTEI6kJTzAem2DS9BGykZTNDqM01Ss
DCX+ahirwVuXs047dQVowLRIVwOIe3tYaU9Xf39uqaDiWRRtvuB1yxcv0yYVd8nQ
dT8I8H4kHqNJ3G30y3k5AWo7SARmPSyUchfcabsyRH9r8EJynWdgPnhMLzdSAjjd
cl6JJeX9D0BUnb5XzvmBA83ppTnCfVKLNwjmrYhx6IvYH0ewTWMn6Y/WAgoyVY0o
nRpwYmjf+B2MTq1i764CJkYtfu3MdTWCnGd95rVV5Y0OtG5VmYwD7gm7KRI9Vpv3
cQgCkaFy24hekLykHai3u/olQBsklS6j9DAClQcQoZBafHKC3Iyo6o7EGgM6Y3R8
hcrT0RnQChr8EKeoPNDuTVQ68ycqDjQMQbR37ZJNJAuiYTa9Wv8CQq0tyUZE9EDi
ETi1R79Uc8NpPjfDnZNQS21fyDezAwvc9meV30eWYKZGVwMBYSeaZAvgBfRcw854
hrt8WwciWkZcaeVlsDF9U39yK6Br1dbn2kiTLO7l49pHRIsxXAjacpX8Anb9ikGC
w38pcl5Gr6OXh/G3K2ptmi3/fUTAAXpJFTSm9b9HmrZp2vcFA/8ycjBrsbmYWkMu
32nZncy7d94yiZdhiSRssCl4wSH8kx6nNB6E8bPeyx2R5fuRMbcLGBf81iHlHW5G
67I/mL8G6eJHga9Rspgrr30qgxnyhTqGZjuGcZAYRH3gumkfWXZTCVUweOyhBElX
ckruJuaoFqrBc7V+cJqdqnA6WecPHked7v+gHDNJZJYz2ZVO7aH/z5jQEjOYMvsT
MvhWKCEHkqXpqN1daNUZVBURheV8WgEjBkizr+ZTQeAcf7oDougSzce/WqFF+Zqg
diDgW+SbZtTV7i7sVy7Ap/6rUDBa89LTnDlEHVgGUNmXVpAGY3GbCJGTreOYZucI
ak4h8D/RGrzvtISoAZJg4eg7YSEO28hkwm6E5Ap6UXnFPjrI8bmj/cc5cGvbxH43
gu9Pl51TCctGUXSc1lv0qt6e4UIXOn0q2wOJkOoWvdrhSltpr3SOWZTVIBL8iPMz
bFIVOIoL0T1fDp23SRiRCYgA6TxCeJN1BMOoAaCv0wWegUhfPG2cRblb0hbMxXCa
YeIuID+RGp2gf027RDHbDn5pnQND1FvAroilraDKP0o5X02YVkKpPMzUgIY4Q0p0
BeyfWBZzItivT+LxbvxvXLNgl3TCag9FQidfT9CaPpr06wAFNOe8Bb8hdFb8wukA
64CYCrD+bVOlI3YdBKNgAWMlfHCU1jt74eEj7nyKsfpf9VFyVmBfMM6pXTSXuwE4
rPcqlTTYz36CZWO3TmwavKD3Sy8354ZB0vqwbMJgszTRs9ZcFfHohiv/kv8Qj8SV
uXcAtPtb2xJuD4lPZfnartYKwN7NgLkCWNojbQqvOvXTXlYfnklX1DGxHA1Oj+br
RsO3eZ9stBgoWZnuJtxOv+9W8ucG/G5/+lKk3De5AZgRnqFuviBRC5CMpJSTlZeq
xOL15s2tS1bgAJuX3DV9OhNrueYaCEF8CVZLZwt7kFF2fP41cHusCb5yhifzUYis
OKvrzi/7xUhGsUpGY28GV9V1WND4vJ781wHAFvXi67BMDdqy1tgcD9O7GnP3txfy
tFe5P/8vQsNe9aaAw4FXeLSC3uAgqV5gs5mR5Qn6Je5gpL9rDdty/YW7xPnigbh2
ZRTJG0UK95awsxwinf0EZdi6cq2Rnija4YLc/q6RnEYH1SRSG5vkngefqbKTk70F
6E332RjC/xHRdaRQ7dqM6sTGaWZok2YznSD0UmgM6rcnDAi3PjEExM80Et+PfQ04
Fdal7l7bgUp+Q577x682rTGgLiHjDSIlHLprLZHxuucj1pfGEaYP7kkrI9fyUhd1
Pj+jMNyKTTgZ59XLTPCOFUhhR0Znp0pQ8zs/3MybwyO+uO9mQjm7kdyfyWRUC9uT
BOPFR4YF84RWLiCyZoM5RMHgDAZVAfPD4w3nynejC/hnge55XgT9SZTO03oNDwhJ
TP95QeC5XR/TyfviVyaqEIFOIv7w506KSNd4OcN6C9gAmjRTZjB1gTCM5TQT2FWx
n01esvSmxNPhCATOx1naS4+C0hD3WfnFjq/Ca+BCaDmPfbixNNTpi9xZgbpIXvxX
+aqjX3Cb/9i6We5QcmwUqRDGMIEo6g1qfsWWJ4BGIw0l7/dW7IIcLoHUyXvNoJGs
WkcDHvrJaXq9kmqGoVjnurNUd5f3iAqHRsWUfRmg/ZxlRJEV/f/OCFIHALy0SFF+
aZn9+xwGWXbzsZB5fG+/Sz2ct9+o/O78p7C2LbuFijawZs+yTlpeda5YedGwER34
9zbpcP29vdXcbb4udkA1/T5ZywEdmPL6/FDA/lkZgQkesqogTsdQiRSXtiaRRPKx
e/GWmWQcF2U+6rowaqNmuoZ7i9GdAkZ0NosD/SxZ3VTaQF1ppyeLYmIjM6P8oiNj
hhnWT1rS3cVcGMXeFcjlVtirTQ2YVOCD/dcc3++5Sr1MnkmsYGMAmLrWcJ/4Meif
4MicSdW0g/kKOVY0z6OBh1FMK8vtKm0ZGCAyYElTtaAdqNqY8HCNB5Ra61mIc1HS
IEs2Mj7Ja696RJY6mdEABdk4vop8U84SE50+d84XaNYnZ5vI9xLcfiZxnvpPZ/Y8
TOqAD1ssxeAPhtb3wHQotNSNxll/jakykH1/JLt3XBjP4hVfdtPYDMiginJPEieS
xKbVrHwQ+md2N+2ssUYKA6E05Ib4TwK5GuL60msnTHmDtSUdDCjy4cYcoYXZnpPT
+LCAI960gDOfpu6aB5NVtZt/8R9iik63hqTEq/uePbOvvzi16mX5ESieUQaKFeT5
iv7tERYFobtfNxsL0yAv8POhPU+tl5gkGO5wiFfyBn2tSnzdVK1yervTnRyXJHcH
VSoDCcGtRl8nCwNIJuc3YX4ZEPcEtTNIJguWJK5eZkjwiw4W/jqS2Kzy7tfg8DuR
fEn7V+G8TRCXPNarCMpUFXaej3CFJGJA4fxrQgur8nuiaEVwTrAFDMUh1APK5IbV
ephrIrH0yfQ1b5Vu5KXpIN8iMaEvj1VFMumLIYyh3B0KoVgs0iJQKe0N/fhgcvpr
BzFMn+e03bmBsehLwF6vH9o2b0Kx/aSD/PHz0v+9sZNU2Xyj7bF6Q6aVOGX6TlSx
Nmfr9VIZZivLxHe8ODjg0WQ3AZv3szA0TkRrpupUE66ccDXm7sXWp9C2H/Ggl4H7
vqP23/crYMJ+KOhcsm+BtZuJ1rrrSlgUVCaOcvq715fowNrzae+H2uL8JQUZjhVd
yXixnvYKiO9A2gpJhQ00FvRKeVwVCIVa4yoXyyf+lmB/s2hcrtGVyA+5cID7Nmbk
TuVmPC+jWdgxW/9yiEIuPZXK8+g3ZQGktp93FCDCOGOm6B2yjo+2t3s9CjPHipY3
g14QaVY4DnyZbC7A+/Zwppa3xvcuDbIPNYWuJx8e2OHMus/3oVmpeB3WZTH0L7RW
fz0cR0rtUNZp+Zpdc0CRlamS/dvfmym9pxyF9H4rjt3XL/THfIL5rQqxNxlr0Owh
o/jyGuPTy2UXvw7xGtQgdN4YVqYf3nPOzYBAz6lesQzQ1sEUlycvIETwo9qKOfrS
ZItpjHhSOndrjgXOvg3sLUeTxBz1Yc4c1FnjcQNNH/5yizS1aObAyqlLICbf6d2T
rVDy8Z9XtB1YBIclfCSNKpUoeHPtM8PNTQdsHsiNde34ohx8Oe6IbqEwz/34/Cfr
tUz3qemqtSvb901uBpbswxLuQ/t+L07b8lqUIRhkU/gcVaGkREwmLlygpWIQF63q
prVWRBZondDz3QHDNo09Yxi/KVKMqNht9hSicMKkZ3hMc7S/waVjV4GQ2Of2fXO8
ecCYB/fpU3vd4DXrtIXVdPs8ygnKv5R/clmjWCMcb2yjK5Owyl6YAouzaPNObGGg
7TsGP29K2D4A9kmZfJgGOpcfYDhjgqVudhGzbNJtI32BnQnaQaU3tvFUgmC3pGHe
bnb7ZaR/a9WBUPTce363W+9KJ9Cc0+B6bhDqP7NHmIWX34jtM/6THquWaxxVj5Sb
vDTa/qdLgO5g0hqJaYkkRGbcs0cVwaLBWs8VmKQ2f/Q0mqFSImKpM/v99BWCVs7F
wtwlAaNKL3sRfB7CP/JF1CCRaBqOAw3AtMScSvUTcfkuytxr8XuLPcP50szY84LM
qThGAN+DqgW/5Hgk9WTVCyBWsgY/FVsNQ3RkTRFj8vicOUtDuAK5WvnlhoMhhspc
rJtzzfxZTxtcIT30T7xgrMtEy80SFUoIelb+hLV94MFiGiPaQPmKKItoI8FkflVO
tWUaq2Vi2h8ZFqX+FjfwiMtfPIsbd+KPVRdKeF826uRdf1yYpBPdrm+0Xm4JslyF
Hk/ecJlm4PYwXKFcXy6tcahNP+lpHakZQgHPWLF/p0GGhGPb/59b0JJE7AHt/25D
gEtfrFyrxxbHsa6VEzhDhWSVf2wnbRB/fwbqUbI+Bwa5Gsm2DdS0jeNvWf8Kar42
QHw1z3DaMI6HWO9ANsZ1UGpEcTpPnIVHH6SiOBU3MuLh+XzuagfekEyeqL7S52Bf
6mftPwyN6dxgUKXwx/TbGouUF1CqeA7EfVXeXQl40VUXfz8z6N9dCewGu6VXaCeY
06F4WDPt+ek/TOCqXMUJQvNZalWHw99oTMVrgwyOvqwXPmimlwN3EhJzd4afb99o
QFI3MJbsTO7XnLIitz9MAeSet67BQNe5Kf5SMR7RGksHlPMsibPWPobd4O1MyGQX
4cOrvk8rpO9HQ+C5M6f/Kt4KC8vOGXYm7asKlTGVyJ6lWl7OAZrQNn2f9MOlvGri
4gN9qXw4fNvkCfQ07r+ka1wEN7bLR58sws1M/P2+YUqSewffRjUqh33bK1M8qUC4
SzEfFwIpXvDltn7pDpRGAuKApqLT9tZ7yhdQ6CAzLgrSlWRUhA9qc7PcN0NitdfD
fbfb5rQoPiEqi8msH/eK0aqYPgpTPlRVHfTDwjyWyOeniiRgFKSOBSpBL6sIyvX4
KSIdUOn5kRDpPeAN0Ctf7IsRyGE9s/WOtkSQcar/CaRyEawzzzuNTIpIQFpH61Gg
/YnY9FJBr1dPd8N3GprqLEf9iQ3CgNHImH/CkUdFhZkApMqPdDJ3CDizmGUykVz3
3W2bvgpwoHzyvFccwmojvfhHpBEJN8EbKuL5HPZH67/qy7AAFHRoGgrULeUxWn+2
RPDSlXI13jFvZ8eBpuk/el0VW9Q0PdWOgAOvp7YA1Bl3r5uf16Me8YjCWrmPKfAc
4Hi63DvCTGlxeBVdSZSALkpXGEeddtwCT505VZnD20peS6wWCZdaYi/mM+C4KjGr
pzdFsU4evqrUMeE1p4fku5uqnHE/ifRDwidc/lW+9uohrEfV5C095rAdqokw45qZ
U4LXAfGR2W/nfOm7PS/l0IblsDKElP16OdxaMOSHdUUUV47xdv6IVyLZGmArEvqE
VkUCwpdu+ZI00IFcJl/6JAhQN3qUFVnJ6tqv09p+qa7tCGNoh3pCBJUkf0tXgMdP
7iz8GLvhDN9XRBxXvb2rxAwAc3hOuKcv2IpdvWT5cyCvsNFwZ8C6P+9FLI8QbojE
gXnEzk2Y3ZHiEh267N5LT0r48YbNOxWT+ovcklYL/adh5R96v+CIqSnbhjgAOESJ
Je1Jt3J6CHZs2zAZjbpt2fRWVaZZ389KspOaCtHunDKlNSiZ5Am+ulzi3BntWoeG
D1xYtWhKvYfFRP3rjPxH+sbVnPD/ooJzSZ1L/U2jYzwBJ16aBRkFztVb+BGRQ6xV
AVDCJMagiLzpK9dewp4upK+NxqHeQ496tI/sAOdlp9TIP0K0yprmG078HBPGZqlr
GiF0e2/uBD5JrjYhtGqwK3q9QKFWUG9c087vF1nvmP3DmKVRbnKuChNtB+ZwpLSQ
FLhmO/1Ygmzc2COiC9qxdRephVUveRZGCFsgh7GBY0hLBGaAmIVG2Twb7Ny8SkLp
Nim2K0mb6I3j3fVhZaRuGXZD3w20fAH7y3jRoR+TNDWH+g63fJUgHzb3j+XpccTr
29W9iYDyK9zfF8CWUnlVEryrA8KccUQJ3fGzkUzl29th2ZJOoUK96JcL+NsFk0ck
bsS62nwcbN65Dxf7FmAbUZlTDd7LdSv+BFX1rgeGeP1+qV8bBAzN8SUkHdvDAhd+
ExZPPYmIGWvJcfYNjYUMgTLCS97LI4ROtLvYYck9SvLhzut5Tv23F6lsdQx/voqf
cPGdNElFf5Qm3IHqMgLNy/K0vhvpLgziNBmlLrw2xnY7xuulIPv5s9GZIPLdxpCP
wX1Lh5QgrC3UwFDl4drVwDbJM0sU0vAF2nV3IfcXRwxrxLt652M+UY970LR8aGCK
kXys/vnEKzde+MzjxugE3sL0HFtJGCmy/Af4OCFPkP1A3MgoPL+6/vickfzFEMzm
nktLJWpRhID3JiaAFh+cYO4PhE+pt9rqNDHa0cfJ54R2RPNOoLKUZ0ub/7yGJUsJ
ROM+ShjFyhBqiw0cvHfzgk4fHxm0fi7Un1w9ZhhljBeVTABgn+msfYEhUPw5fDkr
Tq4T5KK0OmhKSKRLf+CpwtLyVYCtDncfYapz5s94iNEzNCiwbIWkIhd7BISFde16
06SDvqiqyt1AB0TpxStyrQE3xrPh7Jjzwl4CmhIl3agUNkUUqxDPf2BqBUlyFZ1f
/nF5G/4ul7q0pIAg3ggiTLFDFOoGrYNvbuItmV1/9hXwSpmcY1vmQUCczqEJpAgK
KVfmn4yWpBCX+ektHJRcCsYvq5WBQxOuPIdsZHnhP07wY0o2vAoF9Aaps55XE2JT
Bwzealb/7PkNQD31OZ8FiiKC6/M2N8T3mtliqoAWqCFPZHmXMx096OxCOaLJBX5Q
lzZlvsOh1mPTQUpTFpbUvmRDa9CqGiisfNgCl6CfCXiBwtwENLfL4JYrcQDfi4Ep
xhZvfvnhp/XauPl0axAuUZft8W0hgcgdF2IsruTatD1vEN/La1HGTpy4YVgjnOfR
gRpmKE7bAhmmzCP57A17iSKZ1Yu98Ul3Ud0dTd4IGlTywRh9ZvJcZPu0TkUbDs8q
/AbE9FD+CieMTtHQG8WjGBx83+0n4EcMAE+ONtihiN7RNbWQXtVxlfShxKDQmiGb
Wl3Q8nIr5LmqrBsgw2XiFJwHtc9+rfzqaaT/LO6hY1X2OMho0fVWYU9m8Mxx9UjD
TSlq+0iAj7PM1f//O8hSVSWoioNJe4yx1oQfZwK+PSmkBqbZSgEiv5soMFDG/oTn
h6/5sB8SVxtNCU+a6K9rhaMRniPzS5BLYnP6jOjGti2NON3LjMzIaen05HuT3RVw
AnXof9YALXjAmW4ais9LAceW9sQcxDApRnAhhml4f96dWRmQDdbuAKBzEmnZsJEy
Jip3R/oR7GqK+Q7mUQ9G2c3yawqNXLcvvJqF0e3Fc2vLN9Tg3Utmyp6SObTLvcb5
CYnQRNZQioTl6gU8Pm/zpVoDJQrFBkvPZ0s2OwqJxCUU7+4iFAXy7ljAQJM40dKI
5GZpq4GnNRluAIRs5UF02GFlTStYkfJ47rHpmny1+kcBngn77C3a223jI6hs9yAm
O97gVVIOshNncytHHfFmJDC5j6GG7oHhI7lVJrp2rZ6uxwcCGliuQY1bBlfVwQBJ
ZsDPfMm3cA/zOlCnagFSXtfXzX+1gIvU1hynrwX35voJB/cDCcN6fkuOdUqFNRCq
CBqEB+wggknvOEmcqq6N+vFqFiOnCW/zbxdI7yThI4HrWINDVw/MtE5Ohv8rZvch
5+214EOBCOPixKJHIgVI0psSzz6Zl2+0Svq5ASFOG/59ntb/n1RM0Y1vcdChW3t5
27CiKUZiHsEObvrYC2M9osW7kjF1X3CbHu0XIN1U3gGW4NwlKAt90DvOpIYqpAuW
ARUVPLE0Bzd1OQLajhNRZ/aMi5XsEf9TNTS2kUbEFd1EKVDvA+R1NaNn0vDLl2hH
HBRHlAfydKizKEQyKORF2hW+7iK0V0qp/rjjofYz4AWfVz1Rn5gfX02euPCgPKyG
f7zXdoSfRLQ/HXnLb2/CFdw2HhiG7hWurdXktcmtbe18PJqHe/+7MxA3j70xi58t
wP9+44C9+AabizMurq5QULDcyQRU1/4lqPvBocs9u1m7T5YVNcWmJVy6MbS7IWTu
j9BlURynFRwQ9Mw7045n4JcMdzYLatjfCPaaB8gDvnfxnQT6cAzo5MFjk1y3fe0n
AiPs5q9gwgYZjq7an4Ua6G7V7W8lNIgAAcR0ym0MB/TwJtTQJmaK1N2V1w6+XdJj
ib64nsSq595oUSUMjaWsFvC3hvUK1p92zy5mKje9fyBVKmeF7vJ/ToBay5GRzq16
BNeAWjQI6cW6Ca/y7T/v7bp4/JWcr5J3vV+xh9ARfzqE7a14VLbkFgsf38jgUgPW
NROgsWSyx3f6ZUoA/TWnY59bLQGaP9ck8WOIL9aBCP/gxkghs1RTR0ejmfTXMNSy
kjIIDjagjDgZruBQ8H1bdgiyBIsHZS51ppVvlvGRObI+QMIWVppjcvs0T91uVELB
FGqfnmnEd4BxKfjLEcnWAcMcXtDMVuB9OwZ31ipiXmvwDIpiuQHuOLPTzB+J8Nrg
ke2GQr+2vMQ3LMKDWjcKAmkpdC2KdHSgvLwViYODuhco/+dTBYwGcxnU0iYFbBpy
Ls1BqhfedRw/UUWe5fbkaXZ9RsmjWiwvhKUT6lTWQn0Lt/Y5BqQaQhkDSVd49HNk
G19nP8b96T0mEgdlmY+FTHDV8vot43auw9a7N4TDnqRXnX4fofrq4OckZcJ5IUO5
dRXMlSlwjo8FsE8UYqTZPxdCkm5ISub6wTFt2d9VeuvFecWftX5PqLx63+Bmbx8k
jZKE5dEk2zYCWMn0CulLeoPTiSK+V3I7woKA3juQhoonZ4pTJmd8/oKroV7EUzUS
s8LIylAquLVhB+kKyl7c9vepHzvjK4xit56T90mtM0s/gqU2xDjlu0MVTjGah3GB
hAq6VRZ9KEx6IsGjd4JD3BhnZMetF7u/z17AMv9OMM33zdEqkQ9le+c//60UEoSg
sCk0+gC6LthxuuKefNHoUxD6gSQkDzXy6R5ZRaclBmf5npPiyNrpV55hvDM4L1bJ
CjhiapUeyFRw+n1o6ndJXCx1GHlizjuljGuLPTqOA+6CL+NK056aoXf2E0qml2pD
W/ufmjpki92X1pdF2mAWkbcXrFEwRMiQpbtQYyH4pWpOlv9wpjlg+KuwN3M5UYft
9hygzq3s20KRCapSFQpkOMasxdK9QAz+vkNQ9n0kw4XQmegZR3wyf39MYkP/Ya7f
KwA4ShBGYIgOW11BLdXeiWKcVdDBt+6Ps8ZjkuMXxML7YEpcsLBa/fdGMl4BSI6h
5J8kAyi5G469patYDoVi5xq2A1zKpDFs9v8ZGCZfuPRzbwJWjPlykJJaQ8R0kiGD
Y6KU4xhQaVBrl5EGOn4CLSZ2EyVMhdJbHEjt9U+Y9q1/90wS8HxHjPfXnVrP9Qup
imAwBNJQBKu+74VBA0gLmlmxuCMJ9u+5prT8rsg0isMULn7OFORQp+UOOlmX1Sig
mFqksYsnR6om2iRn5Y6XG95ep2+w7L/3/WvCrVY6vj8j2u2zuXmXjexQfqFpqZpM
p+HBiv5z7XD/6ZNSgWxQGfbnBQGA5YTHuvA0c5kkbaw/+6kG1sNb8+Keo7KlomX1
7AU1MbveeKvEWBWPRRQDUquD/TmbzyhBgx4k5cT1sJx9sKpQsJBAW06Sn4xnIyd9
OtWHkn6YiWHL9NDT8bV0GzK/iGFg0Jn4C5gaCyuuyBpZAzSBtWCDbTEdJ3RmZWVu
Gz/I80JSzuyiIPgTEsuDifhY0nhkT/gyWiavAejT0Uw5pKD0GL4s2qXpbT95mcby
yHe8KQT1mad1NUAVXJC9arVmTWx685eUUtpQD3uI+pl0RaoY+8YbDSx26lx0dNWD
AVPVnTmrDw2c7tk0Is6WUfbTH/wew8U/GGbyPKeKE3irYG/mgPPVHO/V2Ld0RunT
G+x3vCqMIt3HckoDU+XF/cIfZe3jhs7dKqVKkwjEFjWHd/kSVMLEA5KN4t/3bRfg
brItzwQFBYtjIOnxTgqEQXKlSWXZLPnKDumT6JZytfufHYNRXeNjEWsP9S6RzZOa
dbu9X/9QZ9QtNPRCrGVExtzpDBo0JzT472NqoLhwCSPNh3XKtUN1N24SGObcRvQm
X/Dw7CgurHxlTl4pfabNbFPi1dn5MD15ByRtF9yGCsGo0vYkIQU8CWH92+RvO7rt
xkOjLXtEMLN6pJFDIEDFGs3LaSsgtCxkJl93L2PsH4sK//8n5LBE6essi+J9b3g3
CFWiN/1Z6bP4BHX2n/iCWdZvYaI3L2SUHGkK9HHy1vQDZS3qiFt66C/n8FAwdE7g
6jziJyIsEqKdoMvGUMNVhv5Gxu7QpWjFAanFFZTvH3ZGvLi5K2PV7EIM+gZF09yO
L1TOkHgbDmIhmVlfvbxQl4LbdnCzReElP9IHAgrA4MDTeFtJF39xnUE++NXtbGqW
hg5kdW2imKoQfYEOsMFG0EOKjsOhWiq7SZCFOxCyss6TVRWSz9F3ydjgGKKb/kKe
9mVeu+yN8cy306mbK1Q5wnefoCCjaD0L/orLwFm31CFEIS93CxcwdGXczXXXYbcq
eCqGDiigliiTAWIB0GIhtyzEXIrPGvYeJZItB9SDr6GFZThMTl/8KGiGlUgT3RgI
A35HBM7+KRLOy5cqbV4EdfHtbSbzCDnb2vNAhh5CPExIucz8DE7g3ANaZLMAdYWP
l12CoULa2fWp2FwfQV2uUf0Q2VL664slj+lPkpU6vwq0/cANdZueYtsYRHjYuNpm
tj4z6IiVtdjwM9UayB6Qfs8eDeS0W2A2NcGPWmTtL0AJvAIdHEipTQe5s4Rb+rlH
EV5EWzGftPuerxgTVerwvE/8UbfFpjaelPMCTJnEXbSZUVTMoTtcFvT/B1aa6uGN
BwKQlAuswcMNKoc73q1il45vWL3YGBc4P/jLNbeDvqtS5pYxJOj6j3RkjbnOtn46
GCfTpcNJcnTopqZyb8jXipSZe/U/Rz/Dc2Xl9rp+7RbcCAY/Wv+8+kvxCU2I02R8
CKttpFTHKcL1jApnIIFR2ta1A87WNinw3X/lug4Zm8GG7iw7hgWGFsSJWXN6apIe
g6jN0tBvTszvob4OfJSsrFMJl50qrOEOrs45aMD2KgNsQFBHYPCgmwEcdLMuLsYK
RXKInDj99ZWREkykzep+QJpueizWCh/DoPg0UfdnVsnfarDwj+2UupTQxcrGMZAa
Cr97J6KET8cKzuOf6A4frTE92+ztnkH16L+QfH2T50VTaP7cBY3eMchOA3npZU8/
l2fla9UWR8h5+Hk31KGkdc5ZMtme1Vmbbu03KYLHsCQxIxcnjHLhHcAvIvCIEkDr
A6BP/pADyAYnO2l2MqlCP3dP1f/XWdph+e6zksBeQ80Nxvs9j56Xov9OrG0iJoRk
F4/NVbzt7hBnwgLiKXhoNYoB2aLiRAncewgblIm+UcC4SlZfiwOQ6eres9ssgFsI
BU3LZAeuExcoyPgo/LcRsRfzPHd5/dcY8N6+N4JOFSzewuXLUIpQY+fg/uAF6UcN
7r/eNvbxJ/GRd2ZPGD3EqTv3cF7hYBPD9MbF7DpIUSe+m7iRFlJPiDJFwqeDBd4W
I8+6vtKPyM9NjdaWD1E3eoRkedV7aGY/HXnd1CK2qmpBAzUyfHLTb9B4g6rGEkD7
eQrkdu2Z7FrCljiGGYVQvRlFX2rItySOmrqfU5mjFYQE/HPV1+XUGsHP4frODHS8
p3LdCDVQsMM9o63Te9a0UKMsRQLeoKqmALZefjMXtgllLV6YIMrloZMCbQGXSffK
+2oF3XQ0+OvofG2Wdo8zu0obNGDri4814gLujo1BlDpS5219UVC36wxTHCdn+HP4
9Uq1sdyM3s49L77uhExarvbFONWJ3wOAb0TGriDvmmPWpYCizqm6Cly+N3+OKMh4
wcBycdCssMZFAVrdwezpo/LRAW6OewomSNElM5jYa2CWwj0gt+S4u4CjJxuQAaFX
hB1Jc37wv/XRfg+PoIKpHypOElusHW1ThzvkagokKYwUCoCaAr0jxka1tfpVzr1n
N1LHpJxu22f0EKIkIB+XzKbyPkFvXwYlGQnZXBPC06yoajgmhDH7wTmGyeak+F7o
Mc7KOTKpxTm+7qrB7Y/ygbRRFkKLJs4sTI5uXS8bAmvdjJsHuDkduDDeBHYklgC2
AZ63rv/jZX5Jgg3b47Z6ztZ6JeypAItNsKqavOu5qaNo3wKXLiJ3RcO2Qv7kQF4p
Aiz8Hr4BnoQS9lWUIavxJ7gaYREH8EcvTLT3uDnEfmrENcU59Htdu7by/ruF66L3
4ttvvhnXva0pX4VnSBskEI+JwcCqI3iiYNeTHkPMW2Ho7aoYv2VnAOeb3j6HrOAQ
M8J6IhKYNlQdlhqpPwD7AoW3y5mx3dSRUu7w8nX5lPO5hz+UFexEG3+Vs/yOUpKF
8PTIwwW1wLT9rtCg1Iy3XcOqoxGd7XuMIGv43sW9rnVHWb/Rewxz0og3Bu4caDD9
0LrSzxv39y82Tn/bKp11IAPNms8cbG4+Y66AF5dSrOq3fT5IqsogDs161RRZmiQy
+fqg04zIw60wDHARAox74OHewO0mmMWnPPgeFsHCGm6UIsgE8yvu0hshYS9L9OoH
Hg4aGUgQ3+TOS2miGVNIeMykP22bNxkZ2w0hSgNzsJ3DQhO5/TVTBvY4dVLDPtJT
s71ahfYjQHKBL5RHz0CcQvrybbkIbzeS2b0WaMRuvyDnZATs1jojkUFH7ioM9lnT
aAgzcGvMZ5EAflI6Sp5ySG0aau8vJL2JVY0tHh1Lxnuw/YNoA3NZAyN2Bkk8htuu
oeVaIbeLoeGBH2MMLfmyq8xn1CiQRCtn0aHzrCmGgWSMN65xgSKxPrgTEPvYo97o
LuHdohGoN+/gqgND+avZpOe8r/DgGHF13OwR1HJiAXhhBU7EZme+Elc7bRAehR7p
M2LmBPv5UAE2CNE/pc8fmW4RtmNTJCmtAuHUfkOwDgjm5VWZswH4r+tBrK57Tu4T
0F8hEY/6vuSbSYbHf+Tl0iIG/6NkEv0TjBkozKGTmNvbaTA2kaY/kPTLNJEdzc5k
yCVQeLzIInTUp9hBF6v0dgE2kTWZcxeFeKOrdBq63BjExLenreMCP+J/wnlG4OyU
54ppeMgQlUR5zCrbJbaMEw+F6tFDHSAzf6HAZosU+aWFitl9GWaSRoscQfj4H10f
FY0gX7LnBoBrPfpTQKd4NRPgy+wck8rrKoVu7pl13Vmd78v8TNc+WKRA2NcYpt8b
wZN2bGL+8o8KoYTdFKt6Q+bcVz1JGH63O+dQGjrTBBaN5TJWKhFUu8tYmJza5GTn
jd6RQ+d11inkilh0HV57Wb4c0YiBFSbSWhAkCpNXBBVNPRCwTRW2PxfqQDIYHOhQ
PVo/08TDy+WaZg6z+/xIeZomx7wXrl4xngofEhWOrW1y5pUH4lunkGJlfHW88NuF
PhvZpvMpjq4F+MhlusSA+0Zj8zFTvHUmNbK3RErhrtxMdT5tAll8EQpMb6nxhvo+
snFiuzKp2MVdlrfewjgIb+0VDZGh3CHiTEH2WUhmt6Z4Lnk473zvlu/mH7WaPCPz
vJqbnD9/j5Xfk0ccKEGrWWZrQsHm68JVWC5IUQyP2xhZVTx1K0e8yvkFtpo789eo
PiNN1s+f/75kDINOFBNjR0z3ndRI9hN/B/V/eL2tmCusybTtt0y/rU3DfTCmuOmo
YIf507T3xKttcD1g9BzMjbOWgfu1GngDmnFObacx4SdgV4A7zgwPP/qd+Fnp/iCJ
F5ccc5zmKeLzW96RrBqQIgW+GvQNAnl3bfIjkDBn163nbXZjGGw16G5OpO4taLLI
reoDnckFQIAS5Iv5IMWtcgppb0ZTRIw4RnS24SLdWtJHjeta1nxHFZNOw+tmseu7
IOKzP46HfASn3nEFSOqePoHV3LtH4wShNM6HNfb22yd/n5bFsP/mVhqsKR4QjNak
PGrRmM+NO7jSt2cmcoVBvV2TkdfcXDrh0iuiV5Y1HzEeAoOJmTE6j0+JevC+GPvw
dMLuXPcc4zkGTzsrsxgOl1OWXkdjBrWN3yzRF7Vr5joBfDSXIRf1EEW5itxam1Up
j7LRbTLKfYbPeyYotwIDNlB+21987YMvoUbbdc0cCjCrLqiH3CmQlaCAt7NZqj/Q
vEXAgz1U606tlG+CLvgtkuW8wp8GzeiWLw26P1ZeffVBIU0k00Z2Ho8qKFQpNzJl
wkkyxmZydPMh8diTp++JOv9C0dJUMdd1mGwJwq1vFuFq7Hx6mlZ4NSbUFho7WHlc
PO+lBtvPokPcygmpKpz3IwgIIRYsQiaajtEML/sJOFLxyEIgMs23UkXhzh5rJunw
Sw4Vm2Q5W/k1U1lw37wFtYtFE5l8xpnDlTiG6YgSe6NJ8PgyuvBbBvKZb7UZdvvN
akiAElCDcvOZ6WPKQRQuefHxQX/sqrKp53qd/0j/wvC2xlBHYn0BCw4WyOIbLrOd
vEZGPUi29LFV8Z3axcsq6m2J3axHRd+XA6LlNTjP2A5610Mb1o+tZOpY9JlzCpFY
YmKsNx5uf2Bvdqs6s7MZxHra/lJwuBl2Yl1wZ2Xy48+ByIgCuQvJSRMtTmelzpSu
nDgjiSqJ09W1Ts1+PuO0CzRzxj/BbzZYDzOk/c826eGLsR5xw1qS6c9XJtueC9tg
aeLOz8omHiu9U287tNFI+1F2nNZ4CFEMr40QOPEGhvUiEGFGTIPMD9V4wJQ+mwtk
lrcXEA1vV3BUEF2bZFnNDbT9HnUVAYtlSxfG33KLmpyzESofftXOwZgjvhW7N6y+
2Y+OksLPhvX6WkOrm5T+r9bv6y+mHJtMiev3v3TyEnRz9lQyWxVnR9snw9O+81WY
cMCWeUAT+H+vzfstyK5S/7zXl2mDmuM5zruKwI2agkbdU/O5MCnfMhcuA5MP6b+m
E6G1ioMxlgy06E5UKdTPv21/KFMMvQ43eweDr6SojZDWG1BnX1YaVIvd1wvYWVom
wxtc2+8Q1BqDHv8en55vcLzFnHMjHyRIZJ0+Pv/gK9qoVRlbaoNb3cs/fH9RmSi0
ZNQUxteQrdtTT/WFOUzNGhd2exmyrz/hjEEiASfQFi4f/HBu1iud1XDYQCvr5V8N
oaJIfnirgBhSBi5bzxCzD0LvTzomN1rth2V1HAgkdumvsam/S3/H4fKlmxV5m/uO
4u2UOBcJE/8KMAgFlE/WcaHCeKhA9rLNNpA9zpBQdpfdY3rlyCEHyxbNh+Pk3aDk
ejvgtYE9/gpBbmXGfQHno6TGYiXxBjk9PypS0gJAizlF9vGktNV/HaHLwdez1eUB
Yrz57AwJUmBf5k6NXtl6L4dz+hTMLemI4N4HkXIC6VzHmuLC6E/fh+MuKKAkIW6D
f6H7QFiZDkycSHW2V5HOpHSA4RemoTWKon1+dFBURYFTCU8hmTp6cwlltNmpzMeU
+tSqT04ivQMmJSkGR4s5NHw2yYokG2MofOJKHWq16yM51RdPYAIjVMEkU7aQQR7r
0bqpsYdPOwkoxthcdObJZGo5NsySQnAaVDiZCHVNwyjB6dOQvPRYgfkqPSMH0pb1
IOV5MPIenp8ZixAJCf3D4dfVJ0qk/cuCxWBvGFdVq1VrJdvBzg1J1aQFvPKNab+I
Eq8mSCo+kTBEoXZ0qGRcu6As+TXV36nuVz3HrGzqEsIcHenSWJjydY+unlL5oRkp
X+qPavbZB9/VywGfXzCNoScZvG5WzWzcfnP5pU3QyKqvOaERbF5JYkAn+3+tiTlb
z4kXRcMz6NjRNJUPb48SCZIR50NhR8evgE9e9HWTEHwTWV964DZOi5MGdZcOS3NI
eJw0Sy6k4VC4oJLxuyc8HKkcQeOeHJ2Vk4vbIvV2KPck09iN0cXqXvS0qRARAAN2
snPvPITuTusfzQTbQu7DylSUiyDiBveKpY1sHU+IXokABYBx7Qo/oEItM47pC5dq
Zfa5093WQEV8WcKRkR0sokdJ1/V5XKBDHlixmWDlIzaoo4KrHffSfKZdSxs3zgQO
YV+g2qfKa6THJAPTvx4zrbkccx5t13X7PbxD0SEQbN0kE7aGaDZRfPIudVUBVFDj
7N7TCfZG7V+hwItcljpssUJ8NoPS68Hri3hIRQ1v9VN0h3k96KUqiWq9+TCpkWA9
+rzQom+TcemuqTjJiTFEupGlb3zb9s3oN9LH2xqx2sTgZiyuS7Z2uf3WWz6KMucv
mwSdXleeuy+Dv/38/f0/cFvERgZmknXXJvcmK64JbCoGYsxxPy/vooWF0orJfKcZ
6aCuVshA/fDVFj/h7td3I4l7FX2/56A3A3EDA+3nCNcBpNp9LGHD+cWGJ+/ZExg4
jShIsUxMR7y0FG20i9Ki5527YyP0/mlPazgQ5s9fmZ+ymTpWmz91qeSgElq/DbIb
OW3wnQ4O2jPg1ZDocN9oEcNh7KvYQViC/EUP6J7cV3sue8L5fjW+1eL7yAhpnjmZ
PkOVJpk+Y8COWaZJtCQg3hNXUV5YWy2P6L8NzMFwH8Yq8+hEYCoySkX5buDYE05R
NhiAQsWyV3NC+ykPc5smGPSXod2E+VnxDihDEM4atZgVTXoMwOhWw6zr2gO7ulOI
TgpcowyOxFp6k1DHI5rUoZYgFKCa4sX6DMtqxSIwtlADPz1cYQt47BLY8ub3rIN7
9fdo01Sja/xerckzExO8Y3Z6czwlIiDutEvCmiJZOB+RSW3ljAx33py6sC7b0FHw
HsA185G86zSpGS82rPo8lPAHI8rtHBWTpJVyS/4pqw1flc+/K8siMOYY0WBcow8m
pyopoKF19S4+/H4qAguM4K0Xm834LleBlEcqrDDNrxh2NzxpKmbOovMD0n6R9mhm
gUWGNFDuyIZvHHV06+rC7bQcGwRvbtgsBcL1qfi8ZM58tnHvW+4HlMpMucfdEmK2
wPuh9c2GdGMe/Row98VZSHBTHC+VKZAj4jC+Eufsa80643ZFBDoxinuTQhZmFg/p
4w/3nrEeXKOPP68+X2EaSYeJJId/DgnQo5vRL1U11GtV4JcgUU5gwvrlhMx3Vebv
0IFNDLKcX5/eJtaSXflBNpyoAmJURIw7vEtXnEjzZMGHd3XXsY1SRPPCwQHrZeu+
+5YFXiCAS7Npk01dxLO37Ti/pBPpuVA1RrL9l/tX569d7sJgKFJiX2eYhFySLLQO
OX/Eisw/p6ZBHsV6rJrylF/E8ACECQfuVgL30azANXn7bV4e+0v8EZSSTpaox54C
tLcCMd3vUS8wjizujiyWGUSDIWnUVYy+xm0gArTZFG6VTSfJAw9xD0SOGfKuzT7y
8+MS0b7PjYIdIbzFpWT4E0wD2yxqKG2N5Kupxa/7z1h5S74l+0nAEVdIFokPe42l
E87xGAHcOHN2E8r8qjgKrILYlh35U1vJNc+Q0hq830KnUZnDBZoe4E/UEZuvhbtT
l3C3iTep/NtrBLWgLLI61egv+5j1nRXpnit+z9WlrqBPokVuDROKzNCHSK8kk5qc
fAvtdQwbcnHTIBEhZU/2qntYe2MyHrJ1zwNBmWGKN9/XLuHl4yhfAjJo3e0tZCKD
8zW18p0axgFRedMtZnPz+btjjeeD7ygakh9SRoI0MI5gXPKKLpT9SK63thyhcPbx
mDue1BO9ydiGkwWJpFaPLVTIcRvqjL3CaPh8m/JWa3DZc0RORdEQegYnEdOPpFP4
2QPQtbL0O9UiJpU8PHXuQeeaS7dSmbLIWmEASxhcSQYjQmZN+jqZIAWmiJGyLQKH
/UX6CpxuUU4yG70f3QdJZ6BMfVE1E0EtRLli63y8Uiy8uCGJjRsgYZGXEG0SzDDZ
e+xFWxeLP9offSCWeJtbAZt0KahDKKB+bxG153SX+pDldh/0Qa4lEFcgBO5Fgotd
7PmNIZYftoC5kjsDf0gw3TZvyd+CCp8+Om81IAo0XR++IdQMPIjxcSOkk3n0bUt8
GiYpRP13Mea1jCYdDEv3Q3JQGVgP9C5ZGxyyVqFSa1z5X44+EjobQcRJt+zhM/FT
POuO9cJioCCMbNFWZNYHVheFKRFV/7M18gEsPXDi6fBM1URUdqUAHc800Ms1hPHS
zaPGF3NEQzLdyFSxxhKNrlJkN1VUfDTyRrNQrFms2rt7mj4/mOwZG7UFudpompD5
2tIM454vTslqpP+8jSKv8C7P8HSVEeXttRPrpvVfwOCENhOtdX0JEONOfvUCP/Px
07bDY9RYf+9cyiPNym6L2uRwCEdcf6ooRnATRnokak68Ryx0qUGlgl1jSLLg2Duf
oNDih4x/S2fpRfHn1MBQtY5LqX+vRQQLGd2TWPxQEOtQHVAccXvBo/z0MtENuzxx
OiUZuC9ZZ73Z2ITYU82ADkQFfvERRK5emehdGJiJtPNtOQ5P6YgWO760PwhPs79/
Ain54VdeiqwUQfXBVdGyHCll2APpnXEIkAvt9k256ybmJAjYpFUHoQUCWBEeL9zC
nm3ohLZ3S1lvtgnvMEEXwVabVvwd57tT+luyy3IWXMMmakucFU2449ZfL3Lg2Mj+
bQKZSukQjGXxvubZx8s7QEdDHg0XSZ94BSKmgJLC3vQh8gZMjHSgVoMe9G4KepAp
vAllCLT/g4qRZxcWfaueY90zqM5ZijaIlifO2FwTYEKpH61LmzHdhhFFhQafiUd/
t5JifptA8B2KKayCNRtCO9H+n7eWpnXhMF/dp0ltlu7finJxmqbtIX6BTTQZebFi
aF8dbnMVJ3N+9cdL852miHE19PzapahslQQ/cMAlm6zjbz9wv9LbESpaRI3/2RJk
H7zsghXHp3tXphjz6E8HLnqVCzV6QfEVfBzIq6fEH8LzKJjNfQexu/qE+1tMWrlF
Ma6HNROKzIbr5S2ZGZHmkldYB2OYJcEggADc5NdB6zdwosLHcN6vpl/Ok4T4Mu00
OXh9b0x5vPxKi7uA7p+yXbBIx7vBvi3993+yncVuIYmUh0LuzviVUCQ6kfVbtog3
5nQX5sTePjdHtryjepJEjDKwY1TdBu3atoGPwVlN9hl26xKMaEa3IgLptMvDm35c
npRJvJGGJ/2ncCK8ghWUAp1aLwkApM38aVtl82SaCJPUIGX7yLd2oAlPdTs0odyW
uLGVu21jrwLgwRSiyL6G6+EmhNUU9QwNJ0uqxYy7+HvBo15bWKvRH6w2carBzNnf
vEWI4oU1FcwVwu1SNueaHtnDW9Y0qXbs7jAB9GuBE8JuZ26QobmSPtDbEvX2JKra
rIlSWVeCsOL9EEveAOyjVMQLVNC8Vp4gg/X+tiajRHWkcldExg+caa/CpcoTVyf3
4zzUvhAr49RZd6dtK+uCSi7wcs002pL++X0/cN8W1Qa4QmOAlEzvKSil7Zk537zm
QtnNcTEf6BDfus4a1VOpTqS5TCBRQatwR73RHKbRVSmFf8bbm9Nvly372TyClegY
L8C/Li1dr7tpNnHUOgeriAZ/jwuezqC9YOPHKUj8gdHJyb9inEEqESJET6skCdIR
ztnin9Z058T1DESRVoqMKTYx7QhZhAn2Cayi1XaTziVBPS+II6eW/JR7B58puC59
+gnOdTcW2fO9HxvRzhdObAkc11SNnug92tj+Tof/wSwD2X5AhYSELtroyBZ8U/rg
pEWH29fGz57/0ATWZy0LUJQ6SlZi+/XN/STtnOSpO1kxrjllxebQI7cgJQgOBrlt
OZqnqchXwrWh1Ro4B2nyBJnXm7cf3NPuyadgGn0gw/ImwBoFqNvraatQ1ls90LNq
MzdO5/H5leOw9BbeZhz9nmz9KGh3NEq3icgnZSRYb4rKzzcggNp5fUzwg3jNrP0Z
fPY72cyLQxAgtO7cvd00Oj4uQ5J4++5V3QqUpYK9ODyJVjaPJVSc+JEfk3JjXjfB
9HKu1KORZzF/uY/MY2kZ0NAqiaWr8KfT/qEwLl+EzfmS02l12NTgPkcJjj5LJ25Q
wZwDSsjfLIA2HKgYP2tKirThByZSbU+cSaxr+8oAfYgOTR/GZqbCCErK6KMBJr+C
bBcklYfLe9wxXvzYjjtbgWG/nbJvgds5FEteZnvuSd56ydcsL7upd0wb+XYGhbau
lhbtpMMe8b1zsmdAMZGqwiJJar4indXG18y0oVrm63TJn8pHMf6eKCfbsmJwYM+O
X+M9QNUwVOwKjPEiYPZG4OrLe4uufJplRW/JjNb0mU8+EFhaVKVHkML5e8DjmByS
CKnC86T4VRJKmi61fYvNatXTOl7szCq7jnzlKHptdBPOjucxbPYZLR5ydT5+BeT6
aGMRjB2o62pjP8aJVKTkmEng7buHSxpif+EfBQ5kKo/rAmpjaCWzzoanhb9ddUDp
MgbgpvRLrDSTieuW37B9GKdj8zWa/7kvMZmbt+YtRSE77AcieDfMoHlfCQtSd+iW
HSqJ9rGQelAbYPNoha1tCKRTzix22/eAks3okD+PxImfF0wKA6BoJm5HKBSCymiL
0LDaAggqXu7XuoSzb0XvVyMqi5JDYVobUeX61D60lDERs9fvKjT1/tHgzpyPwINv
+ZguZreFSyz4kCIXHDRlENsiCufE2w9ck11xromi1X6CSeFryyj6xu5XHT9SrHDL
PDJjMGitSdRqIm3TbGAJw8jHLcFEgRtQQHdqr+OKspTYZhbyPBdDEoLIrafKI8cb
iLKpSEJ6sYs9oGZcjkgDcZ5CYy/kG1A14mVHJi9+dWD6O/0VpBlK51h8xube2cE9
tiEzWnkM71zyZ9sgBPzlgJS3QVtRnANfyzHOluWIw06cC01k6g41sX+jo9IXu36Z
WQI20GX8O8hEAGQTAL4DrzzbaAz9EhqpIO7WCSZMSUOSMWCva0mGmZzbPeLCtmDh
uEKcT6JenTn14kD7F/mTINTTKflyJM7q32bGb+VnrmTzpKMnUZIrWiEzMWpf3hNO
umkQnhf7XononL9rwg+64WptAIXDXaC3dWYIT3koUTig9lDHxDJkfItdcf9Un1Aj
2EJheCvaoPQTlyNGpbkguEwEFxcwV3wJVTSFdh/Wk6RkIxPH+GsYCPfhBGfzaBt5
JF+bsC9LIMxI1zamA7SB7ahbNOH6oJhuUKRQcKo2joUVxGPDKeN/MdZAXZRUyOdA
ghqVdPA9YLZBIDIKmGbjEdrpk6lp01gOJrsgnReu1EUb4b4pV9cRnktiRS/rAq9O
viOYwPs3vQnJvn+S9nH+7yWmsmUVym65DVET8UYQjRBEMaqC+/cLS48+OTYq/E0+
adQBT8re35gRV7XVGzAP2FiBhL34TAAprm9H5qViRekeWuNZU2pATuL787TcfedD
l9mXQ+KH3Ov3a0ImWD0Bf7l8XBE6kyKFvz0uRmnYfMj0f7IMfL7roDYJlgPy1Mzs
YCzRbvth/LydovFCbPTNOj1tFsTaIvaBHJEuK5XkqohC45QBiMzEFx43IMmbrcjD
zyrvJ8V+MohwKJ3VAMCBxl1ChIdlBtzHIhGkhYSnRsrJLqN5unjG2j+tbKHfGZVw
ey/U3QWMcz4jzkOjqj6DORdxGfhv+b7msXSib2EauA/5lStZKj0C4COwk301yUyz
vHf8oanE5GeXLVo9DLkn/cWQC5mutjotvEG2UUG9yuwFasT1DcZOw4sLAvnBJLtC
JHuPeTOjbkJaHWxg27IJAEj33Y8WccJVFeMj9vYCVJr66J6kqoixTM8N1GQeVMD1
B/hMhsmZN313ZMHX1ONYUk8VOrafpMMsG/A5Sm+DH1HTU78rEhpOOSO7ZfUFZRd1
Cl7++qny1n3PyOteSmx8gJm7xIOwxMSQRroYQfNlZPLq7lphJm73K820kpkZTlei
k88W1RdYJDYS4Rp9CZhGlTR81lH6ULbATPxX7IHRjfbBDReLdW33jntMRGIlW2lP
ulpaeIle5rTke55MW6xOvzbr52hogHt/rivclLZJraeO4hO7LvB+noA+RvFCobpv
9aCUKEo1KcJmzqlzhXIHpfCBkWxaaxcj9nfVq1hdk7F2U/PhfwXbySBIvBlAk7zv
h0+JfNzHZAd6mJb8ZW77G4nYEoeajVVOXBBbHwss3igVE0LlNl5uGlpWUXcx/t4d
WaKbkK7jCg9TEYyADDsL1MOagiAQFqVqYtbIS36mqG0enldkM30IH8gf+mfwdx9u
bjVWHxZjDYMhE2D9cr/Ng3H4cFKSctQ1JzvMl5LJdA17qD4ekzK5CIZISa+QZjPI
8/Jmz/P0FuGbVAPA6Iyn8/+I15IOQ03KuHfQs8a9auwb4DybB1incvfciQZR76b4
W63/sywq/tieJ16FFvJEqgvd2xZiyt+r23r39N3T0HRY7pE9is+hwdFyHiMWKugV
mBUmvqBZRZa1mbzU9Z1NUE2suT7dQZ9HQ7XbSir9qiv5Oth618EuMO3OuhNLGgkb
dYnf2OwfK6NeEXL/cE6nfrdMV/MAa1iiHjfb+aMTCUVjF1d5MDA0oO0FsxVg+fo6
eHqsIl3posk7N5zhjo9RC8e5Xh1/yGGVud7FH3T609HFmK0pAdKACkqwvcCr1Y8q
zVgUfsG+60eUcSrq67B+OG2ZwuD/hTr8DkUM7Pv9PnYOCIHaFGtM40mLzY36WgSY
ZQk88Tiea+yJPj1hyAOiERlQeYhTBJjOr5AdFVvI+BMOr0ZyJvCdtQ/V8zCQpkSG
yYxagC+P5rYBc2V3KJ+DxXUyzFadrxiNX5IY9GLfuanjjWZBJTI/+g9ycnBrgW9G
WLbD2H4Qv8k7VmDu8mPOr2nEkEjbNchWjB9P2FIF0/CX8PYBdkthdYmabCQ3C3WY
V9hyG9/zjpqYy9mccaKkv+GEyMWjZCrzrR3CooqFFdrV8bNH4xRvFRPxLIcsYwnt
40PammBLzC8xSPOGNRF8W3FZpv1ubV2ItoILEDvXNi6ZdEw1TSwu5EOgQ+7KkoKo
mxqmf9IBG2q3JjAfRsvmw1C71NZGrBQhllovtw/DruiDC89xrakUnR2EG+zvlb8m
UxYTdUsYOOPsvVRbh2he2TQYnTe3luX5s3Iq+FfKut5+d0BTJdykFci7vybQ1H4s
vVAy4+SBrd5B5UdCw03IxvrjTKkZWQo8YR8V9CUs+TtldBevLr+mthompIH0I7Gm
Og651M10f+m6qmJo06gsikzXzS0yX+hdIjusgmxiCklVX9/HbrtqP9H0ngSbkP3o
e+hkFyaNjE/yKo4gcLkTLnvBM4nFKMVuqYNVBgaLfrumbpJ/5eY/OG1X+SGM+2G/
hZ0dig6HWGEkc26lvA87kQ0OthhJJ5JPZWn/SHCuv7ZFZkA+w0+Ap+a/VakEMdC1
zDAlzwYrlgwnhgJww4FtGxVR/+L90R0Q77FmeyhermKC8whPkRtBAJrSPq7OTYOF
cB/CwzPi8wnmze5dYRVTkHhF/bkdjcrV+2i9iSO2Qg9WcIfBAGIpfAFTW14I3F2x
/xnGlOUt1DWdLURSZ/DC8nJCnX0JrVTKkWyyf3U1O03WBEuMfBTkkJ/IYuUYQczP
bh5cnqJfGrB/Q4sQgmAg071EWk2+rk555F0rZTfZ2fYhcF3882czQb21VwZnrm00
AtxtUs5Zz5Zwo8BK+r1xtdYqi2z9cLnPaTlTr1dVL3DEspW3NTRVNs2movTM2xAI
RrnOoawZr40DatFgb3VlT6shCs4FWG94PCe0hF3TXxr8ABOSdGONXMsAZBk1FhDD
cXXFMtMqOO+rt07ldtVDIImSfwXyQkqUzWD7YyDBRufaUlnIdtewL37+jlEBeog7
mVTcnnIEYwPDUXlqB6AxWvL8O/8j3gTpr/F8BJFTuxsvQRCWqbR77dxiEEBRUJrk
5CH9MikzXuu/lYylf3qPRbin89/1zvpKo4Xs2hdqWPmlPcieHwKrHn4rQmw+1uL/
RNZoBz1XE4gTR93Uom16452OOe3Kq8l8/82tcbARgbTDBWmtQ7u/hLwxub3l6vX5
X6uw8kYVCPvBa50ySRMeYuFMT2Q19DxRE+okJI+uPMVXST11hnBpmVgM2Ogu7GWu
B7r7TrILR2CAj/UEdvQs0l4FKt68zkT+OJfXA3k3AQ68Y2RvTuA5qSKZ0D4pVOPb
0s6YC1NnHqTm0BLEXWqZNaaCyaSM3yigRh0QvpvG7bX2H2vdXeorUs2jN6H7oi82
kZn83O5TugbDzc82VU95AeBNZXHgMdvDQMyrmT42FdI5srhw1xmA7GnXAQ76I6cj
Ia7+lkzuxWpdQVdmgN5bMHb6Vn3AYVWFzdejPGVVhygR/tereUhwmwEIrpcIepOB
YNYIIW2HkpqXxdBbZ4LVAwrPupozdW1zbMlrZV6xbffCEw47hin6LMnhfJpB8CEl
ce7aLv2p/Xh9g65W7IegUf6S7u3RePtPk3eumdxDaSmrdZVLxEjstPwDqw+w2cjB
lWRS7lcHTBBwtciE/zw5xyOZJpbDQHeFiwUp/CflDyuzsDe/MqO587ZDWEM9aqLr
An7XeLoKbNsv6+3k68gtCiUzOV5TMj/3L2hk06CsnbsEW0s5S9XFWeLujofJTIeS
8XvuAhAgqVRzMXJF5yjYx/FqXbeU9pmhoDko9F/LiiGRCFmrkj1e8Nrjl4qhxHZb
NNynKkI8w9hCGFA7vUD+KymcytMquieQSUz32nJ6+APNbv5SBe+lZQBEF6g+bZVW
0ixhR9IB+cCywsy/T2CFoQkVoKSzXHE95N2t0sMu9+M1X3iUVsh+aro4rcIQLViQ
v3TmFekX0hSbJcHGdeNbru/OpiL0EIOnBJqQNoFv/s1dZ3GpFYkQcF6n/TQ1T7dW
fGvEMHV0ZUsXkZetQrJ5O+c/y4jmRAS5Jqlp/xFcJwOZhfdfEFXO5hTFwUEX4SSV
I4ey6aiq27xWgdJze1eraQ7vCcRHU8x2ZFHubpAYy1+qDFa2SkFkV4f5QyM0/jzW
AF3kPAYPEcO96OCWLSRtXMOcGgDnX8KNMcv+tNnWkSz8ep9zryYpQAHumrpzazXX
DAeSLQgnChpmOaFxdh2MtIngtvSR/+eiY7sAX8tw84yDfNS8NFx1Nn1MYiWoLwpv
+BcAy2toxElwrdxR9gRjAq0OM2/rOLQZgntMU8tnlrMpp7vbtENaJrztDqJw+AJb
fgpMzJcJzqsxt3NATYt9uzpqty/64Alh/2Z0RJvsrDmzLWrGTi6mNiXgPtJYJs18
TkMVcvLJ5l31/ioXGoI5fQNAB7lENamDMN2WmfwCr/WIoWaQTTF/NsoPJyb8LGRD
LGDxuHV2ZWkA+bPyohj+IugtDPe8mg4BEk8MXFSILpHdjz1p/8psvEmH5+js3V31
wknJx8xutxhTzCMHzXPEcLoHiJRLOdqH0bYfFLzGSGyVYXlO0coS5/6RzLEtzlwJ
+yORFjrCV+FL9Xj/GSzqZ2qGwEz6JqrZZ94dP+nnbKKpxpNL9E3pBPhyvM7IXEwJ
dyLkoIIayN3gaKmCdwwPsrtnZeRpP7ecXCLmGnd6J9DOlbDQbY6+qSWv/rJ4TZNg
EvcAYr93EsbC8EMwDgWQcBqdeabolifAsEm2H2+dwWY12ccHSzA6p7KG/zQnFRwx
HXtepeIhr4rbhmUZZ4slAy9jOww/l+LW3HEUtlps/7nJaR9Iqf3OJBhTlyKtHMpR
+E4YppVupYIa8qH/QynDfjemz3Jkmf7BaPihRCBSWylZ2ZGiTOwlIA0gMKsf2CKC
H2B2jmMRioiglSmT8r9+4uaFv8wy4H99emL+OrJOBWR/6myGHTTu31+IGDNikTC/
z+VNpEuGQoCgr6NLcVK5h4EzUQWK/ter9v0epVAJrduCz4TIOyjaclcc95jGtKmV
gLieVBPLDimg3rR98f5t1aUOiQN+xdUlTY5cfX/3BL2uWTXRmZ0AYc/EE428olER
PkG5R9yRrqNaNYynXnDeqoC8yXgr0DrfHZVpN1upAqri6LZC3M27WsKFZBg59Qs7
Vys6gSkl8S/5CHAPo8ixqAmOvf9l5wUlqEKDxfuQDMYCnZHBBu5Oe6zy8mFAcWyk
wtfwzBsKAK3KAysam6dzZt2SGwdR1PxyAbtidsPfWvfWZOB0f1WtmcLHn/40wHye
rdyyXnNMxwhVPCexTpKeC30d2h9Rlw9FYpRaj0GfIVV886TShP5JyS+NNGynDUxU
XV+4PdoB5oU8d9WK/lOgZ62q4NZeCGKzAvjRTz7zsv5LAblpBCdY3+34Jx6YU3kg
OMXn+0NrDN92FaFJHDN5vNohhUT2ogDmdH+ej7GSyjcnQTLYLX3Gxy5k+rkVtIZG
WuI+Gil8DJRSTwkpcPQxctH0RbRN1IuOdPiyikI9L2+Ry7S3SpXDQqQt5On1EV0+
Sk+/GtSuGKZvDbpyT8PQ7DBIcVDd/OFbGJA5ew1shYAqJ+CvJEme7Zq/OmK0EUdU
z5GVfQ6ddcX5+vjDPYILqMcdhJ6iJ8MvXolm40B9TmN/shnWY9YP2NE4+Azh2RiT
xl+t0fzwi4E2oBRuWsCro7Dcih8R8PaURO+ouAwBL/R6XE7qMgH2OY30zk/Rk2yj
Loj5vGAYUva2UyOmCAjayfR2Swnm9B6iIN2m7WeUgvbr+y9Tu98PZZTa8FSa1kk4
o3UwJ7cQ9l+StDaKeknYmfigA9DqAatpz6QoApa+Jv6XM4JGkuKscy+3axJiVNxC
qnjwVl4AGmcG7+lLwPHEptII7iCgbaTKoMIbeEGFVuh8Ct4p0/d424UoEaBwssOh
QsQ/OwrBs4tfQak/8zDLGhSN28NZNxu1M7XRUxQ5o5G3DQ2chXVSaEPs/q8zp2wb
FnChjsHPY52L/nrx5qAjTazLr/Q52aJn8GCUOSu/h4p4ewyFBiStTcLHod3eLV9v
87sE2zGyT/lP1mvM77cBGTWy7SAgrn+hOX4zLClGNwYnmMrkt3hAKavdmcrCewus
EXCQy9K0PScuUbJFKGNVtoNEtP4j0pi3nBSjQ4gsjCCKU/HXahYaCcB6wOPkYFqJ
oz9sCWl47bos6e1iOUt9fBhYuzJ44YchUXQVkEj/fdcmaAHF41V98zkrEQUFR1Xc
HxJ6HhzyFRh1qEO3VjZ/KGK+iAvTLgxPt7d5ky1IXdTkRjQXtkp/UNBNrJGVj11J
aca3fr+JUzaZp2x11W58AvylFq+IEMrWZwa2fn+1xLQAv8GB6eKAG9k2XcQii3we
w5zMaHFoen4gSeu5C+jlkaAY+NKFd/W5+mU3V8IRT2VjD6f4E8fy3vm5Ma8QfzN0
hTn0yu0y3qZ56xDNUyYzXm5rLI/TUas+nw3MqV0kAvjQNfEHTQcpaeSCyZXdq/R3
UqMEkS1Tq4kB6cIebspmuvdUy3hE3z+RGq6jAZKDxe1tdpu8/2YNp0VZwMqTcRcl
vLzooictwVzcBHY7wnVly1h5FQuptARl2Mc/UgBQ4X4/U1E8ko0cH0+SlOLDOPjZ
rz3o7YVMciyHCmFn2QFpC4+sGZuDJSqGztskojRk9vGIvlANHWJn8Ei1TvKqrDkE
PHT16PVP3yId+xZ882hc5mGMyRks8KziUbEuiSyIWXdhhzy4j1X3kCtDOHLOTgjh
aV/1ctRRUZ1CHM0TOJiQ7lx5acdcg8fw4A5AYg87Aq9vw8cCkrlmVOL79D09wRNx
ruH/qIlaenNXfez3C01eBF6Qmdf4whwCIfyp5v7kaZ3ZtsBrt6/XUIs5Q9OUfbWf
31n+06BjPHMgBxC++dKcBS/wqVqsOAcBhXgGeMxm48z7eOf7WEpMsT8Fyg6BgPaw
bMWIP0sVsLtmvxGKx9fj8Oqc+vRCwNfiW8aPSCUmtn7Z3A+a1xld/wp+BtrZTAUA
Gek8wMeKGyuqdlukzxzZPpb4HMvHk+lqQnU7S65GhXuAtvapGGNBxn149yI+EG2H
kvwBbSCwIH9RG4B3++3S4Mm81yIzByu2UO6xms0s7TH6isReMFQ8jOyz0dASdV+q
6RwN+Rdo+2Pc68zoJ2K9thrmhx3xkveRM4jsI7J5y8Gq2YEc2+1YKE2//dxxNF5F
HxMkJyR6CeBGTVCYFMAqUR5ZKzaLD77YC4SbnOP/UhDOBfsEW+NlaexJHD+67+j1
KonW9qldP/tPquU1I3LOAbe2FJ+x0OcbbK/E2K4dVEO7gv97oifQMW4N5eBrfbvl
sWNwmC4ZerqdHsIajJX04LYci89kDtkPrz5u/QpwNBc8OU/+zH0Pz3f+gdW7EerO
OFhPpolXprMyqpmBOLtE7s/yBGdqK7W+jxggt7INbh5fPRX9vGOpoDBiiQQjVoae
+9XabSRjWLFlwmBZzqPSryttF40Vt5GtLvQxZqbjcSZLjojXwoPSYAx+2GgiyoLb
qIZngkv0U/iSPwz6cvBemvQ8VYz0lnixZ0E3IF7Aqbz+o6vEw5Ny1ud9vyIkQhJ8
fgeK5M9mc+CFGe8r1bQatH0PpC5eiLVkPlAa40B0BRNsI6xaKweh0DNH7D2eohES
Po5BuRYSB5BwyEFN5jydkWHu2QT7p7EeRluvX485X8vaUyWtgeZdc2bqeJCybCi2
vzSeN+0U0CNMG3yN0dQ1+XfExhO0EJYKSpLykWegRiwp99CUYCAsSHRDcKcptlNc
oMFrX6aAmqz0Bvu2eKa2hF8gC7+qgOmDuUkSMiWQdx0xvSchgbCl+p/iKiet006l
0j71ozjcJomaRfqFIPiBJ7veE72sKXlXAuxcBT4VaMDPVgGLz+DnYwi/J1eu2V7k
KkWoZd4Ya0vV8cmaIoSuWur0vQUJ3X0WKECckevjqnI0LDgkg5gBY/oG853X2EDZ
hjEPFmnx887i/gusCpTk1EvyFb/4yMZdPcHDijapNrMCp+YNjLYG5J6KQ/YtImEg
zJmiUq2wQXyyvsrlUpFKVhNrPfYydMk7bY8huH3jrcNwTo7eSkpF26sVyq9n0QOC
Rzcewlo/Bhumm+/G+3obJP5hCtCmfcV6s/WxEp/oFGszGXOtGKpk62ZfTBNxcPfh
d+BDlW+v1tshE0J1hkmjyzxsjmp3snmnL5c7rikgzcKoJfPm1o3naugf7X45Rw17
oyoPlRsig9DWZNyWl3t1cexHGNFmDeHhTIcYVw3GphVVQelw3Aj3JPgdMzS5gnsD
69Ud+tsUdRjjwZcdSEbSZ4op6kz1ePmme+RZJSCIZAtv2nBh0NLid5yNI8qPUxzc
skBITeFS2lxIKAffF3yCIk7amn/BFsB+/H2wS8dTJpyclsr8bTh5XrjuoOIqmfuB
j7U2/mNgMxbkpUmXA/c9ZNEGDsUy1uy1AIXffiDFEhndp0Nmc/GxaktKYsLtJXF3
g+M2OZgALWxMT1DDmcPOUKJoDNKGzQgZfbWuxezETxnGGvQCPUhxllUfF4B8ic0Q
8yiMVglb6oyIhbWSw1tjF27nc5lc+aLwL0RhMiC/h43+iZWRfHFzJfyvPl/x5rlA
Fgi44tEbZS8veQBBeRSfnwr4+MYpEbEnB37aZiOjDpC/CrFnIBlFDWD6jINGz0Yx
fHrAg/lgXc3e0hye3skNN0lDfRY8i6q37cack+CdbWL9pTsPA1hJ3Qxs3nxAwgR3
MOsHNgytEGw+3nXeeET6cq50q13JsYwUCqQ6vrBkqcCmqHqdP1n5iL3Z61hIREmG
S0glsAl1jpCTmP37aD6rl+l+/aDFLEZ+1R3yUiWNblseq8TblYDJGySh9M3OTvR+
/KWjRCwlfAbrckSccbce07iU6oBxI2lgKPMlxYFjqdsMC10r/WTUb4zyb/l1BemC
qAxPzsyK2iX1Cb+yjnjxfR8d4wSHD8bqMgEhWbdzDS9AFBZZdaiRD70BxhYo2IiK
VEf4aQs+DTAuQhpK4dh/nsM5mQ7eySmp4FHCSMqgBnHMzPGCegbVZcH33TB593Qw
2vvBKhPqevhq1tGDNPpyM3TnuG6G9GiM/7Ovk6+1sLH66liywZQsXRi0Z0JA5RRi
L6t0BsBWZjf+o9pcnJ7SOPMRY6LJkJGizDmnTnKr/Eh3n2vAv6PxcEXW156fBQLg
944XSt9mDX5lvyKUsufEppUAMOSo1qLcR2YRsyje0rjWdnc1U5ZX/OBMqzmX4Qzw
sfkKoOL4elD5S3y2u4tQzrgk4TuAebKaS5AEVBRBd38/MKHkPCJBLedk1yOu5DHj
+vRcIIDniOnvX486wNp0GJ7DcEOE7RqcaYVKG+9Bq/dNWywk5Bm55BiE34Rlzl6C
snh21eISuurEFcrAGKodIXD1Sg9BxuATrtLVIBjoh5uWxbK0dxfiJEkhp9vSU8+B
VmMLVqqjspkuoOrehxoghul2XYS7G8T0oyt8h2SLSKvyACeNbvZUuc4LVIIx/t7P
ZatQKS2owudsFPORyE+ZCnY4/UnI805QUvWwqxpGCsIoM0SCcNmcmbjgCLjIajcP
Y2uSAr9nooFKPkCSR92kkOkejrLJBkXp8k+lfM/dT+hiHEhgMX+4VP37+8g8msf7
Fc0uojK8XEGN17/4raBVafBQKAs5OB3JyC2m3LUtngH2DvH+OegJ9zmCD4xZ1geJ
yf6GkAnWhYvg7opZ8Qft8uT1YuxRmMuyQdt4FOLeCaSm71qT7nQFMA5bXwGMhdbY
KdpMO1q01T2meDdGMVmVOWf++ZpLPmmKCs3nwFs63BYZy01vOWlM33chYgqRicB0
x8iyHmJ+/PmO7qzFsL7oJYWu2VJV9imDux3zBCDnDIHrubwF34FMK4SOJPIklDoz
0fZTDZPlKdFNsONcR5F4JcJS10CRnVlIctDhSSUBAL5Ab8X+GNb3iUSjh0ayq4vr
sBc3qt9rI3c1Yu5gy4KRyp5EvpcczMOv6KLPQXKT5LsR0Ge+VTcYbvb5yDhe6k2W
TsAhK7BLDwErWWIEM0eH6TgOmMA3vvZL+BfHIAfCd/eIOgeMTP8paTbz2QrW9eq2
SGIoP+Yn9JLIwlYeI+BT2TwMgajxjIZ1QCnTenEwgYBbwev+W43ous5x28gsSY2+
w5T3SW9cZFeSgP3roa/Qd7/NtagUB803QoilNfAb8ehz3p39L5vHOka1KVjRMD8D
fztej5UjgdtyVoXYYc5Y1IV6UxMY0AtjyBKkSkSGJwVsg1+ncKZRpN7mxXV7hJmH
wwxRR1Ufj9bwFEIWht1qiIWf84kJ9Ib9rSPexfEYTCS6Q9prvEQ8dkIx3XaJ2CNw
oHkinzaN0rwl/iZvttdiu0geP1DdFrwNC628DK6ayol3T2pUUgttHwldOLOFsX5g
qADPFZDfQ3FyE549AJIS4JEislLDmGo6yf1NgmI57Plt65h/gj8/MCcMTwHofck0
EvO2aWiXFNBxNqflCqFkU5/LXJAhdLTGXuJGHmoO++MQc60TFMP1BLYdBj6zo4Rf
N8B2M4PePSGzfhsggOSngnDonJTadmyfljiatNccGH9zcxKkBh4WoWJS2FHHK2tf
Yqll+CHkv1ONvsRrS7Gh/g4nGqshoIbJnzCwkyvKsqMktuo236yy9LwEkQB1xTxB
DL08ytqFx+bLZUinP5fYJaOHmU7Bxkv6QZ0gH1qAzeoRJlIvNMprNyWa+V5MuW1M
ZFSDXs9MEjXtbdccm1vASr8DPtzxC9yLAIzkqr5BR6K08VNPSZg/ELDCLJ2DIc1E
9eOzqzLuQzpGijE4dJO1yl7P5aZi5UTMlhHS7JT45DLq8QuRWY27tB8bGMaPvxmY
ETUv6rQ1tT95TIEyZNvaSVGYX3wqQpDELLcjYA27B5LCdlkdoQlrvtrUg0WBpGMN
cvAX++r35u+TeuQNEY2Q716D17pj2jF0bnzpV8+VATXujdl6aljzb1L/XpoJkXx4
urS6Lw9KBmn2LIR2pI0jNV/UJ2NcKFdjbshUZoOege0RGzGcCNMZpqiKisPU1uaj
9s63VezMTWvk/Whd9lm9oH54pHB2/jGav/KLVxY+TSRxAsbWVDZSKVwokxAjP5u3
u8Z47e8MYsSHD/nzf2SjdT86PbXB1zYFZHQXvOnImELZ00by21/kv0CmTh6Huc0Y
/hY2AqJiwrPJ3HVhXTdV+Xzra9tbBR1qQ0YLk4rSLsK1Np1Kg55o+0rz5oC5bHLz
bqUibh5swJagfRUaIv0Tnx54l+byPwNbLCp9BQ13kZRGC/7pWIHyIk5osp7MoxDm
DOS5Rk9FiMxz6c2KzdAL4vMFi8PEWpriWk1iij1xC7nGbd0MslfBPTRSQuSnvcui
wkrFjcQiNkvQ4Pw0JAVyQQ9twCwdGBP+y9Ll/GouHcnSxRqB1wkVH3T7FomVlmNu
6Fgv3h9bXEB2z5e6vHGk8784TDajOPdj4amkVEwypmRKDAIg28ivIZqB8pmlQ3Xf
lV5AVmkDbsPfr/6oo8k8Ij+Ll3prH3msWOQQJUxSz1icrPiyTTPyRLPjTVUIcyu2
SsDOkcVwlCYfV3InHz4tZKRs9xiSjSC7aINMJY5da3dunbplSeYbOd8y3HUQ4ixO
2ImUCpue4jB4GSfIzFkrww2hoSXQxIXEEiPuuUVfxz/CXdOkthIkR3NBi39UGeeP
M5Ct773qJLjar1XSMQDudVKkLO00k7C6k5qqHOnWVmOTAgBbHmgdLEYK3XlkzAXt
RuXdlazLRR7R6lQgl6saWT2Mzkp9Oh0lkhy4TXvFQCjL88CQFXTrF7TIwVPuvCMQ
TZ/ujekBj/PaMzhq/W9veVC5UbcJ+A4nxBytJcr4IpfRrj7CfyVs0S4pzYUXa+Ha
bfC2nnFiwqJXbHXmUG2ttO+2fyzs9Adcq7zQ38F6cOntxcbCNb1VIWiVqttEjv82
fVNyWOFJk5Sk9BQ0SK95LjmlQgwig0p7OU1bX+6zeJ9Tjr25QDZKADIR/5U9VWLd
p2u/RiO8wOIXSPYFqCDTzAaO5kwfjgqmZrksZInemgqNRCU8AFaFqgfyAe37maUR
OsR+tjkW2PvBPIoOOmQ0nKtq1vVFyyb2q4krZPOBC+ekMn8AB3dZAWSupcWy2Kht
qQl6o/1Hez5hlGt1cD36MCX/oaMGiKXo+4GezqHKF4G01MAXR4YOix3ouedzxIDI
GIGVKt7pKr3qfNf3II3/kglJRBOe0sgQ5UdLjUqp290RWNLy0MUiSDtZX1GruQuV
v9y6jUUVnvc+MqQ+O125mQ3oppwu1P+7KiWeR+ZerrCV7LfpiP//MqQYpZ+CWvs5
cU2JwqyNyJnczXTQNWTrvw5u8Qo6pljeLZue+ZGIOiAaIplyyX4TyWBx87fgn8WK
Wi/PAR2HNPvG2HhnlvCbDBTGmqFb4h6kOEzGaBsQOfKb8G5kDAOKjNTuWIXPcEak
aBLbGGy7amUmBs69ZW4RosaDA/SkOZOcHBd0gNR/rQ/nR8TdfyDwndyRphEJHDka
N8E9g4tcLu4tGg+4iiqdJB7Fr451zxnm7KPmYJx7tar+5G9iS+IJW8Ye1ocACcZa
ttCf5h5WzHkF37ufItbt4rCZfXmlPQCvIPvamv11e3moICHZAJG8isIO7/Ed14kA
JH52vcqvfPYleDH1qn03O8ynzDDj6xdMYDmq+tE2+T2DfKLPEKzZffFLxCBF43KD
IG0LG47BG6A+izYbgd9vDxaTkXW9uMkyWFVNxazriX5LJL3k+V3bHhiwtGqOlkbS
9qjKuRnhHDXj0J1A9VcWt91WA7dTGtIJImXx1dcgWlu1q3IyU7UZcA1dOELqWJC6
cxhR7QSDjmMvDd6TDyEilMTffD/Kt45Af41BpiYufTxW/i0J9cc+NI1Tm6uTi8Wf
amrOwLzpV2xCpH3w2F2ClR4cgNFKWr6tvzYzFZ4L0Ey2rOJtAf4TH56dbi4D7UN5
fRIOrrW4d3JoM2pwJPDGkk+4cTPSNMOZAdlOUAJl/ruKyNf1k2wbSpZWRnFcyU1y
aQhehiQadnjGbBtg0SBoUn8ULpmQTTk3H5XK3IAF7nN15IvMpH4oKRJB/UlgDexl
bWZBXBCUwLGbQwuIpoYKogFjKRGwZNcLchd6X9b5bKWGsZKiZJfr61VU1rkuU1wv
cIfj24QSHQkyqhUTF0nGvs11J983KLO3Go9WaySe+CSHawzp1pKAiCBjk/QvkaL7
JzVgcCqa+pSLgLiRyZIuVULqhVZEY/5yBsMlItN/bKvIxT9ThnJpLYhkjiUCGlUD
xlIY0Bbljc5kpxYofzKBq5KL5cqO4tp/eG1X4aEZ4EYMaNMFJCfAK8BQf1OVWjQ7
3Ako39eUr7c3u0P+ORJUZ/qsNy+AdFEHvDWoc99Mp8uRLUsr3s+JhQXuciUmpQGr
/KtqAl31dYtsd5fhCQvpXf44B8cGIH/PYSKbDl0keYNiRpevHvlfIX5VFc8WJDEo
2ZpaWnK0Ne0SCfgExWcRztCerf3OA5a0WtmAcLy03AtYLcNRDWKx0bHlvjue1RdX
1g1b1aAnhfen0tsQn7nDNgeKuGLVsXmvcyFDPmNB+NhwLgxBqS1Hyz3dZwGtzsYX
Xp4dk/qVQ9DzWem9mqWsEFmS+FfR1nqvz6QYhb40L70Bo/Uso+eN+coFOt0UZOWr
+qbgMU++TCm7pCDTZM2mKwojLE92YUpd9SOQ3+DKe+fri/gEHXJ/5Arj9tFdfInH
1ZbMy4Pa/w26FdLPRNjnySaqbijbI6GGz2S09ZVAr0nDiSmifPD20RV2MbbZfTNp
mBbpTJDw0LwBxqeev2DN3nOaUmQ48XPudWHDxnIodNAPKTWK+XHDm5faKRcsQ6dS
tBj3qZP0xuUsQ1xlPqI1JOr5Cxn/hdrECgiiD/3hjL3OMdd1fDsH9w0hq2fh6not
eBvMdA6HtsbTOwzHG7xCyFYwu215nFT8xDH+ioDQAncl+qACYmCvKcHkJnWuq/5O
wsMFwVjCi7M/3Ce36dD8ssw4sDkhYlaVYbkUih5fTOB/iAqudbR1K21mv6QIeY5p
7dV0HTgamL3DCG28auz3wQa+XZSImIO/oqgb33syTBpATgPJFg4AzvhF8MedvCXH
8B30eNyu/ZELT9+GxtWRWZ41qPtc5e7PtjToY2EtErI7/GtIc0k3g5r7dTSE/ChY
tcuY3b45NZlKtrafl/iu6gZga9j2Xh4bMbv5RpM8v/IOD7Dbh7VNsMGwJUSSo/ro
TG7sETP73ojtMH8bCvJ9LAO8r05tH7RSLabutMCKdEHw3gxH/5BGA7w4JrK39atB
J4QzAmrXdVam5vz0AZ4yIQPE2cB9OwJm2Vn+bmroHpyibow09EGS0SvBvjYwgcJX
LVFCFct1L/3MKR/gqUj3gonVOJR3S6Rm+cZMbxkBaZqH5VjXPJW1n3iRDGFip8f/
mhq+xH9JPq13IfKMpRq5Iz+eVRkayfytDLF4n6fXA+cDVn+RjjGwAiKH1ufNL+VV
jC9QT+TgRDSU3JBY0YzG61MLENUn64cwh0sWQAV3UV9HDeCJ5Rxhui0R20Ze1rMT
7NyPn4aoEqIDYj23x/XP99JProN8pylj93z3/Z5AtCs+P/TelJ7f2N8lcxOsmMa0
FRo22XXVum5DqffPkYIj0DVhjNv1QVTKDG5OtLs7tNOJTvX8GN3zeOO8eS5q6q+Y
sISTBUlb0nkDZJU6u/w7dXH9jcOhXWWl6GI35L9WJyAg6ijrC+QCZqT0bFJqwe1Y
VidyZk8Taum1iMpB/95Q4Fz5WxIAW62bpbDk+nuDThlOwKfRzl9LQAuBCmVy8+8J
ZPElvT69KJE94blIvIR1cdEQb9Uriai0oUDN/kdaMmBPSvgWLv1aKDevm7MEpNQK
4QJ17WPqvszbNryuk1JAYoLhdE4L+EMK/4Ayv92OSdq/YV/T4+DXXzp2zg19LoVD
HpJzar99370TvExIiISPS8vEpWGaP/beEBmQBLruj77Ly0Gsv1Q0nGh7ooW/pUdt
pStu+ZBaCY12DL7nQNAVaTC+IiIXkF0HcDv9pvtxZsXjsJ/fvxGdlgQATLuPmrAr
FS29L55EA8QMRkUoc1DSr2SVZlJ0ibFkGfteNcNjaZSwryCPlKciO7lx//mzHpmX
ynNqFxqEutoO8OardsZYaKHeM5rWnQRYvE0qAx0/ahTIR3/X7x7cZwOMhKYNbkn3
gtji/cZQMgLxbE08/fMeJeSuMHs3WZI/zec3pwQbswQxlZJODVI6466fDSy0vJoj
e5b2dqMjaM2XUnDOj2PH9AkvUzXjGPvt649xgHK9dqYXaQrtoGmD0QR7lP+kxstA
f6bLeFiiZyjzX/LYpLz6LNx3o5z6kghX94xJDINoXFt97TCVePI2BA/5g9DHyfjp
TRgaZMQjGysV3CWkmwlyaJ0GE4HJbN0IT3UhqfOsgOqzqAWsKRj8EznW4ORC5DNX
fvksl8/YGRA2orPf3x18crWF1x1/MjFffMpY3Fq+lRVqMBk26r2OjltD/xn1fVZF
/Ma40hxD4dARB7mrjTipsn+iD8SFvvCifz61aNYyIhsrIh364klcmEEJFCXAyeNe
E4H8zgePhZ3+jdiB6KTjjFM93gRPcGkAfr6kTVbCK56Wtmca4JsaT38AJmysj14h
zX8BufBl9facugLOnZ3pADX7xOS1kpf8bI3MQWimrw6tDLJNABdUO3dMT2vo2INF
Fwxz0wrqmBG1/BSB6E7ERDBIOFAoVxxiQZ96B0Fdqxcz/sH6tVjoUS/OWDPfCIIg
ceoLRK/sY1EtD60t4nZKlgDRoQD+afY+V8H/Q+O+xS4RO7bBMDEnKAwthmMKSkCV
PDs9a+sNawPL9vJsdPWE9yZQDyYPP6QZOKjLyRD9hVFdGSnLvVUdb2AE1epx5kfW
Dv9/kaJiS4Ry9+g6G5ywN21OjqzGO5Db5THdo14VMxImdbD7ZbhuXdMWYGjGeve9
pxPf+0A6byA58pfLCS+sQ3E3OJQbCWNkgeWGSVbMpa+nth5Uz3+KEiwMG1Eeg6p9
Huns7mmWa671ZKZpN3Oy7R9H3/lLuSGn30A/Xjse6adhnHXUuZNf+zKckFoiBNu/
2DPlTiOfOHyfGvp6ghE+GCAXadknv03ya5ADAtlhKJT/sI6b9Ufhhf1r8kPeIJku
JsF30IapaQ9QDBJvc++NsBJkA0nHB/xSLky4qf7I6V0V8MYBgbn1/cxu7W8sZDCU
BCIJbsHzgJ8mQp/6XRmpYGdYxv7nXP/3xSwzXt+3ujhYdK31Fvu1WkBCBhf3TLo6
peM8Umiu49U78zjmtnEk8cTB9nc7ltIHsiGXQODdJRXbsjjzdmnwauB92TkbtHrU
+vJ6LQOYGJ3IABP7u2KrdCrQzgDXtkTyGIGOx7OFqprzDCAY37D+xxKJf/YmWXxa
2Kvws1wGT8NkkLZHP5xC42VHIRxGD2qNHgsPV/bNmj0Gk3rpEoRXtgx6StBTWoDb
dIeJPKRCh+RwM9Wdr7vxppsbSQ7aTwMAkF4IgJ3uheArSpkr8JbZCKywo3ZWUG+9
qoh6GkAMLpuYad1v6QvdpjuFJv5CgsfV0wxkuP/lDWUp1za4H8zKU+hBCJ+9eL/T
i9LzS7s0t7pO3CD5m8wm//4uL9gnHX/IdQ85MS2MxCFjZiBU81cMK1vweN6z8LCi
rSKOM/RDZV3TrhUhPZ+yLkyPrCwRm7nuBOKJS1LZB4CJq3OiP7paSmoKbHACsFZr
vMnAgwJ/fGwhdICyJNhxf3Icqh2ZdEdKF/jND9VUc/mbVtMkNw04q9yO0qEOjefa
aQmalc36MWiQimiYzU0RGFaAyk62Pb6wYkBH4iNAEp/56CL2TM3ufn5QWJfVfKRr
CZsmN8a/8ylXchFX1C/wZfWM3Srl9H5Aw+X6Ixw6jUfBEIi+6w5kjBp0KIhHCLHh
3UNVCprYCr0zcsP9Ho9JVHGSZrifiIpvxQIHs7UuVqCTaBnDov9C2fZhYd2rBU/b
df26c9ZjbKQJZr91yESc64Y49hTRSwp5gceiR91qJPLyh5DPtUzggLUY5zQ30Rc9
UvbEVCiRDeOSW+JoQSqAyglkzYNWhcwrVzlZxFoeT8EehnIOK48mw6oA+IKKUH1g
kdzLgl1jWmCrJqoP7wiQXBe/ORXHtJUgceODlmukftF2AyMztCQ3rLuJvAzp9VqX
s39KYsQrnkOBhQYA+yLGvBer92mHkaeYflF6hkuspDsJYa2sAkhZRkQiQpqQQA7U
WnDZlEq3ViJP5DRZHNzvqpx0O6YkPlTxICDoxSfzXIqGs3+MbLcJWbDmRXdZ0u0T
kg1/0Lvsf7VNILE08hOYHwagwY/R7SsKPbD247BlbqlmMtPCCxRq5M8h9hx3XnAi
D/aimF6k3fWa2kZadNhAgsWc13ehZ5kvD+K5lfB038ayR3TISAwEdY5eGR5scDFs
WkzxIDrUz0XRJqO8SLCZ3YChN77GMuBcRx9mEm2eK1r+439YsN/uaqDc8W449miY
29PvpU0ThZcUGJiMQCZXisPywpA6c3g0+CPkKLzJlx8HXGC+rA7V9fgiQ0C1ruKp
pjtdEzQJc1jkPWjDfDXI1wMQU9vPXTl3SDb4rkXaha+qM9n/j7zlhnGUtOCKy3ef
fCptLbkS7jsP9LK3GdzoBDTHtpzOK1AyRaHxHb2nwoHQgvHi+HnAmU2rjMUoBoI0
heQk6oERjtrEApOYYWmPcStjIF1YfPZFtIt02pQJ7ai6i/qrDrqR17XOC+rqTm+O
f93IB34fXCSDSObAbwpAyG1MjZxfhLOb18fdWiM+1Vwh6ba5kupy9ehvNE6xozBu
TO3T2LYV5IQ89dGAiICVztSvRE7CQJiHNTTlmkeu0+bZYTw1zT26WSDnyh1kuasv
kD2CTEE/XoWTa6i8Ww48eve0cnc22I4XcAGPvH6wguc6pZCcbKkElNzerK6YiMRl
Bm2sHlsxjZgOLl2hi86KbP/ybGbRzlyim7ZLUiKiT6ufq7Bk2knCZqF3PW+zOjqp
l0d9KWcmAoGy76Fwf2/wlf7w6fSFebXxmJ/0JWk287fJlbdNuQiJtOd4qvSRzoSk
37TODdkJ7KQ6VSxYTtAIYhoOd0GDQGhzX4ZAxBph1X6CTsJBzzw5/4h6ajAvcME8
RBwDELf0Yu4IBui6/CwIJvcRxx3iXVYQ4x45IjIddGCB9k317camDZArnuvo+rIm
WxOTBHfyrb14gAr74GOlt/IKvjU8LsnjJ9yAeElFiV1lX6fk6W6IhlTkhB+BaAnt
6/15IwPqgnSWrp84adGxhH+FRef4RYP5chgY7Ln4knxK/Qs1l4NLNcIuOl2nsdaK
Rh79kMYEM8H9iCtvbv6KIgQlt41jU8KBoT5zM6xsYCMIUThvxjXuI4+O6+CMiKJO
+hL+SxCYJVbJFNRYad9TfHl8xQhMVs2s6go137dlHFAr1/loFOk/SmhcYHG0G5F5
MVzL+0iJaukig0ndSDdolQrsOS0vI3DAO2REbipBc6nlq/KJsxJ5rejqn7l4ubIZ
1g8K4edm192TKHi2obrBIN6numQJKk6Wf2qkDP/t58TS7TZQ1aGqgFz3uLOim08/
2/teke5F1HbviXjfDaRu/hNAFQxGvynP3UuJhmiG+wV01HfhAVPFH8itoBoY3tph
y8VWu3xOtLWYEbLhNOkYFNAjfiilqd/cB9HN4kxLv1NSy2/eObiCzQdZZJjuBMuV
gwoC0k1AlEWEbhC2B1Z3x3OpmZoI8aPB424Klv+ECdvqPmzfHEs3IzxFOaYthxXr
DzZFy3OUFbaqhDjc5kSHzaQKnh+wSiy1FlgzBVONFq8AK70GVQYG+m1B0XkB3k2s
Uob3gT1ULRHQ+//JEonyfQJFP+KjBy7muNbjgSY3b4neDqdfD4GMJ6gK5sY4Qy7l
HNH6XdB+9z2o/pjvoQ3ThfUdC6SlnMkWTZ+il+qY1RIfUQCPMS2JfjRr/N4938EP
XmrrFpvLsDs+rGY8H3lFoQaBOFVVAeEMHnzOZDwcEjWUQuF/R5O2oLGbuWbe+dmY
Zk1eXxATBNTBB8YYJhZQdKDnjFy5zQ8a7T+92lHVTdF4d3LmIl024d5vUmXs/NmF
bvdw0MVY+Ssb9KKkS1Hn9AyMFDvYcAqNxE5edaSGlwTFngvJEOWOZB2FszJj7iGw
u/6z6jZUTOpvh1vnKySREFlYqp73xztgU0tNIgTDifvLl79K094UDWAnl1mJWcJU
f6ZNczmkM9Xd+k87RBkPvbf1fY7D+oLcQIqVrsTYMos5MK5P9M+/B2lZ5VR4o/2k
jUsC+1Wp8/6JlvLjhQcuGjiVkd3aAt2xdEHOok1lv2VHOR0do2wtzb19e1V92qnk
C5qWMQ1WQPVJySx+xBxDTJ1Z33kXtEZW+zF0bvTUBy9tOiNbz0PWvzPANbzvrADa
CT1sotRHTcGGKLeePB/rH6Keel3AbSqDtHytULPb8+M6qJOXFXIGXqKbe7jmw6m4
yO4qrUh8qgIO0AIsEAgpcTR14TDKpIrT+60DDE9iGGtDTVJ1LZRPKfhcNc9vK6x4
Xg3bpCJisB7FXeJ8yJA0i3/HTdX8IoULQjwcZ4FryWKPExxJFaeHcl762hLHhl5C
XiRnsmD64FlGeVUB7Q8JZwuK10xlF2dnhCQit8casCyTQUbcQeUbwitMMOzOaiea
uFlZGGzcVZwZVBoOWANWDJ8N1d5u3i7D8CWiptptatrz+6oumr98dwNLZFm54FgT
zoCCY9PQ/5HLlm0z+xVjfKxI7VPqPcIf/8s1kBJCOV/GyW/iQMcbCrqcsbmFcea7
1k30VAY/qUgezDFhNMfG1sCr6VMZcnmTf0wR0+cIGHkxLfibcmXKEedH8N4CXpd/
ECZXQ51wbaznMFr6xHNPEE1UTNgV5UQFN9HlYxFm8veVCbk1c5Gy+mfnkQX7vCFx
Z1emLK49mcS03QhHOGwt57Bph+NlxyNDhlht0t98R3tYQiBIFE+YqQHZPrUdkVFR
ynPKNx5zSXIVx51UZ9Y6vTGc19h4fLKuAwWEOpQpLLZMVBNvGEcubzan577jv1/E
8Olt9FQVh+LANXYoP+kwPfv+irf3HHGSPC2FJyaDafoZm2B+PfRd/7DqCJvM0wOM
SmOiILseWREfafM+92X2Dly+rPOWtoCy41EZweqAwDQV0MaBGx+WmowmnSEXMcZM
UpBDFqro4s36VscFKUBTK03oAHtYB76JOEHFRn+lmIDz8MVsjDjcUGTEDUh2oZpl
0aVsEsYiM1YYbvIse0pwC9XistrNZUjLLisb0HvjR+1x5aotNsw5AfW8QZTCUMep
BRy+F2luosuAik6sPNT9oqea1YSrMh8Il7bpELG6/6Z4C426xT4SElSpDMozh0Yf
QnsMmHGMwhF2DuWb8uExGOD6d5A4udbTa/BMJoOXPNCoQBTSC/T292ufFVQ+kfm4
s4b4OYXDc5MmtSdhZlx77YL3ppRoMg+sKUaMmhtGwUk12LfP44eG37tOqSHuZH/Z
aOCtRTdlvA50kvY8pEWJ1rO5YnCms+fvvvzCGwRZgGmwUB+iSm1pWg/lYRezI3mo
7V9L69sA3KLZ4vEcGImAfVanhBfdtKD/4YMw94500FA5W9UHv1+zQVzjeA7+JEBS
pJnQsGNu/SQQw19KvVwYQWZfxL66zb+lBhQ6USsp3aVR0Wo/bmWOzpKxp03pfSLL
4M0UNNprJY5+VUCR74kdAqM6tom6aas6TbJoneLJ2vGUK8q1ui57/bVt4Zr8sAJk
XKfFa5Vaqg9h59xXObSVemHRzSFIJS6QI+pC5w3I+QQL8Z+YTnlfN9j2MNnz0BvX
2hTfv8GXNa/bJOt9k9z/zdIfNIIOygzszEv6FNz6R/nICCaVvjBSATGnBjMByk9I
TlspzF0x2OO4CHkLtjgenIVyNXMoqVSIENeKM+ECcCH90iSvqKC2Okp0+/2Y+U4h
mWMB5xZFPCp7lZT4hVLiLPNTohAI1ieBSqrJzNiPVOVxMvgwwMWW4KL/YCEJZiAL
JXXmBgfSjn8Y2jyP9/HJHscfCvvwCegvupP8NQVEDf6C2zA1nu88xWE5FvX3rrvo
D8huIOpGBM89q3wi8CORg6njZqpqzRnxQbfXqAN4MnkQuD8iIlT4h1QDVaKvQu78
B5fJBhkTXAMwGUu0M1TTKt7dUQcUI5/3GR73rlcn7UbQcgxDcLeRg3Rx8MYqMqua
loBlDYLJfwm8BQ8MCfbx5QRPhfCbhUFyI0GNEij3hbqbaNc3s4mT2OAYLpqOu1Cb
r2ZXyK/ciYnOg5a3LqhCed8NCkZ+jtCQdikePDzScgIu8d9awtibYB5bwPFbvIlI
1V4/2b6ezKOq8rQjSZjTke5ndJm9/Ul+WyTP27YV4y4siciMXiTMUDnc9tpj25hC
5MXgxxxcY/e2ULcbgHTwNxW6euNvXrj4+PwRFMbXG9nUPtq+oPREp7dR5e1Wn0a6
Hs48VfhF9CqhnhHOlLbzFuHsQN5T67gaTOWj+6ivIHyfub8d07tKkI73jOsert5x
9riqeIyxLgpdllfgGzepA4+A26oShCJ6LlBWc3Qe5dQTwSSUpk6E27QUOvZOrsaw
VgKHtxFFlDjzoKuY1Ivk4fjBoNLHH/vHFsgdv/XjKdeRBTlnhzzPW0rx9f5j8wLQ
W9Kw5X0TpUZ0xYzuhP4iKyEiZxmoROrIe53Xp4yo3T6JyGLh4cS0ljwjbz9EsRmL
Y8V19AO0mhi6+RTiXll/xxq2y8xNs8km1D0aFKY3Nsk8D7xmUnGnGl4QyQaMsM7S
VT48TG5OHd/YpJoRhVwiNO26QmN0EkFCN4rYbkEMcF6kXC7bSJgqWXUpRn4m3Nbi
TC9AgGa5mIYYCd/3S6rCxs0ioUB8EbwKnDhOgDcPNezG/6NCxvc05SdRNv5CYs+s
2dhZQq1N6ORl9FKwyyzoaWtl6AcEKW7x/A2jmXooy+7CNO6sUMs1xyN/koJPQrc8
aLXKOugzy3gDhyQOLnRNelBsdr0Vnyd9pQrwS+qL6ZoR07DbfBvBdUI8M3JYHohW
IdabRGYejBDfmxEcDYlAFhAyUgnGiTuQrQtfySSLP8+vZcYMW+gC2aNvIiF7St7A
F+KmC4sRaFAzDtJDNlGQdx8cPO0zkCoqDB3KDNZAkcTk+v4Hdr7n46wLBgqjkDwi
lS1Xns8+eNWmvbRDEAjpO0WYvag8vDCfftq74EjswwhL2H1ueqH+pEs162Y23wXj
MB7KPc8MBJdz9q/Hy56T3g3nD9O2G7xp5qXVvFkkUciWXcmRPDReCet6F0IDoDqE
asOeh8XeIH3cmsCFE8jhqtCN/pfUHaeYGmMgr4vaeBUeQeP9StZV2eDDCMY7G5D0
E6M6oP9uTm4tWeI0+Rev+W2jY7DGE+glvac/TkBh5ftk7d4fSbW4XHlGuZWsrmmB
nT/YFLct2KEVi4POlFO50YHrfQaljZ1tFLdDaXyQIj+TXTJNvDTlPAummynXs9NW
ZZhlibKt1Q6nVR/tVRXMI7CWwOkKd6wCoxw67Ep0EB01e5dEmmanxHn2K+r9HIFa
kim4G2RnhQ8wi0gUN4zonmAcSfE1oiRP+fIbRz3KDI2jheXDIdVNmefhwViWvJsV
gfx2FMobCYXC+QtnNGvlNuquF6f9cZKHe0pj1x4L9GBOzngyb0Vr88z3gex0C4AV
woxdLtB0A2tdqL7ripkrQtxtPDcCwkxKX40XuLK63mKVAvQuH8rpgp5PD38kRufK
xhnxMrTWXTGpE+tG6+vUf6o0eCUecgsP3VI/H+Ulx7Evqvr/u8fikVl5Q8/sR/tE
9Z/bUovq84bMhziuFjzLkWUa3kgYQE6YgioiPjCNUC9z1TfIT8d3ZPGLfq8rtPfU
BSSWzm+mQWAggcnHsO4EyyQfOHUKCE6jPzZ6OKRms0EgXpXdRAe3aDRSgcbV3hPB
+AQ9I6Das5ot1rETZ6tuu8idlATz+iAS9ubO/DC68NXvtGeEiSwtGHXKSTJfbVVq
o2xM6Sh1KTwm+9l0LRXKQCHjGAcoOi5pgZAn2QBi/SEZpSKRLHQt0Dc15ShvZxHq
P0dodT3x6xYLmOMWKbTZaD6UejPtNvzVo5KqNuUouqpwMPizwAO9JCjLxY9/7bzh
kVqNH9vnLmvZRkEQqpNxx7zbs08DZch6XJtYFBS49nB3W/CZVgLOsvXnHbA+FkT1
1CURNeFHg7NI2ClmXUoqYMOf9bC4OLcJQCMup77eUNmjqw1oAog7kM3iSKm/bxil
uH7Q3/jyIl0zO9RkdTvLOGxyv+daVrcG+YN4SI0QPD6iQ4mxRt2i18vZgkEkzyFj
gYVPTEg9Mnzd9woB/2vY03179GZo5cOY25stDRGJJr7yYsypW5XNTHoOa3UGFb0G
OlOnA2XTeKbU/ACMqY/W/TNvoS3+0LSCrSc0AQlk9yDyVw96N3vutxbXitGllmPx
+4z5mlQAVyXeOEs8+Vn7Y2rJT3NrARZ76oSKfjZme53/UnafaJVY1c+E31NQB9O2
ktGLjV0b7yzw/vA3swfL8nbhnYAGQiEmXZnCyJO+8T3ESw1ANT3ZQ6QQUNw3HoRC
pJAVn3Tk49Xd08A3lWYnTqzxdESWWuW/ESiM37i9cg+UoUTU7H+CjYGXHuzgvROa
w7EhZBibrmUb2BaBiUTVKG+GCFv1Y0G06bQusbinZ8en/hov3iLPBqoJIMf7PhfM
os3LFmGP4EyL68qjE3Xbb9WWhd4hYX/IHngLQ672np/f75cj04PhOAoYuTPUSEqa
4SYYlDMDypyN99wgpH49cJG3I54BVtJWzuEM/aFbMGZsmAVncq4t0S7AIhMDMP/f
grYGsqi2zWy3FpmnW8s0PU1fqV0e/7TNtNZceaploQJEFCeVvsaHIRp8pnrpi+UC
/UkuHWyJoNuMY5gd4aBrlcI8vWHkguY+C3eS4x8B7hV7TsbFqx+lBFyKDb2/4Gr3
Rulm/dQof+DKdEh9sajUZ5GLhFq6A9GcKgHZx/vGfVluv9Z6PHN7EmRHmnKZd3SB
172zOInK5CymbGXFk+0+2pqaNAjMzqfKdKCDttLZRBwU7uAuHqg+lV3shWLqmG8a
kKgJ69G0FJUlaQrKGHvTlwVNJVEUVQHB/blwXXw4pfZNkl/fUZwVXyXgfsK56D7T
nz/PdghC/+q2TBAMglISJ4DUbWcD0/jrE083ldFsfzMAvrH0ZFlm7qBJmURHzKD0
2bnRmQLbWd1/q9vhblRqqCm3vSlq2ZaAMGnpe1Eb+zNEprXLjl8LTOOgZY3Ou5kp
JfbOFDO5bt7AzSMpjdQdgq70wdUM9PN5/dFDAmm1YjGpJKBHgTfQh1yRNk1k+17Z
dTwwdCh+nXfbG+f4aE7ZfsrmG2tDlES4ujsh3lSyL8CPR63hughq70cT1FELWm10
Znjf4Ec0ANvVr8S7xb0LGhTYHvWzQwlyyxy86Ga8KXJjCktpjzxcv/C5JkTgbVEz
TovqK8bBF0M7QFq2ZKxyaChxHCQ7/2ou/DwPG1sOTJM+7e27n6+Y/MwRqJIkvG3Y
bPfE+I4JHBTRHY7Uc+b5WpG+MUzFtU27gon+tehXCMV7fnRvn0NIrSyv5Ps6vsz3
ntPrIWrCLlgOQvetUPRQAfFrHy4EpEfp9D4OX+RipNSfXgRXuK0PsmzGphzMLcrc
MwCIXWKJlqsqTgtACQzXVqB44dhdUiPVcSnGM23RKsCzstOT/0dfNKBNBAjYA43f
t5xz2/SjkJKuH443IDOBa4OWlOt1n73XAlu6ocqpRxTobkF3B6S7mWLpOgIPxNd5
TbARMhJts1Izr00K7DSk4dm5H+5mes3ykBbIeKwRbmZhK7mIU5rWRuLrDx87JBVH
vmT6Xrwlg1JI9d5RLRMF+LFazpAUn8essXLEr+vP+UsOv8bHHFwoXD3vb+HsBuQo
RxLoeU290h4mEfU4lMbbyaLm9ERPLEeoyLljfJHdNlOYXpHhVt45jIvGxupRTx+X
Xhk3ih9tn+OwNCH9Hr0MPq96l44c9cppk29Lxm68OeAxZLSpP5UyQA6bGqppvZFN
F9R6CVMlguAbYJH9AukPkgk5W9ivQdiRyq+mUDsuQMNPOAO6Lg6fOTYmYNDrXwl5
0Ir6vHL3xITMCIrxGuECAPUhaEKgY7R09OsRbDt+DrVtdnsFcA6joARn9l6NjUoM
UiqZJGy8Eo4Lt6neuh/p/VSOqIxPqdroWhUVVcQRtnVSr6tjcZoQNnPgJZatgGCI
XZJx/lgZfrk/qCxnXmmYafdQvzwVbhSRm/VoxJbzK/B4rL3kbEZVOJgeMIm6CR3J
T3H41Ud9NEnea5s5jP2PWZclN/WQAUo3KGOsnRwRA+zuFOGyrfIs9Jx8Q8hinL59
R3xJkpszIZmxw5NcN22gJNKYbBnoOXVZx9QJiXpGBDPiDrJiwgN+pr6SFEnbqYne
LSCV5/D4qiVvcu4btTGA6Q4QG2g5qmQg28egJy+YQV+xP57AIriYsbLi8ddhPySB
PoklJMas3XDElfnCuwpVgXh/ZRAstMapUap5XFxhweHd7q+/fAcJs8DRXDH6tz5A
QcFIO/kzvE9UpibC106DlTBDm6GUIfP/6DqzKlM/gHORyYbgA55fUUv7cL5MFRdD
F/e+EcwNmNpJt+F6Zt7vhSGJFvxjDpzYIcgACIwnDo1FsuJF2Kk5Dz0017ZCG97S
7VnF7ZCsQhDeeWS+51QbjbpITZmC45NsLgsqDdhyuU2vvdHJSAlGfKgX9edZu+zY
DvWfuEUf5Ac0W80+YDTeENyHmeAWNszyenzOVjuXnKBgSVZsGFE1F0dJMJt2ySyO
a4V1Z7iEVLA0d4YHWEs56KbPb9ZQ+ScOYQNpytu5nKRFm1JdcE4orPWizLfyu9H2
GvQ9ayaf5u0FxEGrh+UXmN8ZjK+phepreYyk5CD6TKebz5dP5KfNJoBnJH15X9QR
H9ghSvHbHct0oAmyVTQBtLkOj+Q1/FgFHZl6piwcYef0Jb35ZquvypulrQ0E9XXV
rWZ/37oNW/kaolkdbZR01KnCQJeg+8ZmuJTwSR/DOlaDXzlR8QrLWHzMQFj61QKA
CdkltYDuCPn2Ed6N2GzuwXby8qwi7SKniyqOiOJDzjq8gJLiiAowNYLFBIuOpleD
6uhMvvfYBhCIA+1nSzoFwUYebt2E5lPklg9RMPnzB9IkB40BfMti/W9vgtpXjgjz
pqkXokEkDCwivmA0AGtuYhnMxbQD83mNaOXCQx6R7T8DtTAaAlH0UI7JyoY7lQ4D
jJuovXMpvnpWq4HATmVG98aQtnMlW1qGtR/rdzCtLt6aXN8ghEnOwb+4HdYOqrgg
Mg3CdtkwBPPnPy5OHw9S6aflBdFPmoVKTM5emki0w6v0BU5j/oG1RiE3In5Q4Rb+
Bimirx8OgH40hpLhkFuq9cqFKITrw1bagd5B5gCwWKyvCUaqnMBg38ZgYWVQ6gco
TgvZbQH2eWOdO9yk4WRV9AnSj1t0CEolpI/o5jZvzQQ53zsBeZqP5tU1AuOqVnq7
I9pe1MwvzopgeKiDrMpseBlKBVdUDfSvRIocZbuPhpEa0pMjemVKnZQq3fcK5Syc
EWC8P/IDK7W/3M0m8Fn7kW0ex1OBnBBInTPo1Pl6bnS2QO55F7rSGqtJ4z5iMgyS
bCXGi/OMsu6eLmaqhvHomrMhO34IAn0LBu2YoDZ+x/zoQgyyJ8qSRLwBUyMxGIrP
oNBGgtmcQZ7vSWRM9b0bSp3UD3I2wXRQ+Ep+Bp4JZJdcIaCsT/2QIVqpekRto6Du
JhwIT71Fjm9k3vtDEvVyZ8svIjgloVfw8DLNLLG98cRFW5gaehyuClJZ6cq0uIXC
XKeCyWxl9fR7jSroc/Uqs8S89p8IX1oMfJLzQFx8unu1vqMpmNRyuP8C7PdbddJn
UDC0cVVbz2reSMP5PM2EX3ivGmy19wcycMviJfzE3mppxX6KnVYRkgHhQVZNCjRv
OVZqIMsTJNOUHdlvTAm3f4OFeF8GFOtpgGKLbPi0xWcKqh9gvso/kpWnGTWF0/Yp
pRitxGrZIhjtBtUT3apJPWjAMtSQWoXyKmIuU/e7zJedLFooYUZSFfSsdKmFIqzy
s4DbzHocgi1H8F+xMZ5nvTOGR3W1ADPlBTxQWNd8GWB4K6KtKngXEoZgdyFakuz7
1L2B6sLu3wwSjZu/Iu2iWyRQNkcf2Ad1UjcWrdW6pivY3vAI5icrf0ronGWMbJMp
lFtxSXgyHRx2/pOJQubB0UgWTyApxH4WoLRzcOg8h9JfPPzkx83lvWlrbKG7OIE7
tve7gGdCYyF0Xc/m1smTqlUvAY7ernSSrhvklJzRT+kk9AXdQLm1/l0vHGBypWEo
Z3tFggZGhVSDVH/8oiln18KR0MvzHBTomUXn+xwWbFIqklzqhy+6ixAya/pmC0HX
OdfC6oncnMH35nTx9csSY+PRkxtr6DJugCwGaERYlAQYzWYARHZA7GkcBkaQEZZu
I+RBvhMiiGDcwdXV6Ro+Ylt6Hrqa0gy3yQz5m3WKnbBQjP88JsT7F1KolSHkOjuC
WeKEaN+7wcuj5Fz8vg9CCEopTcJTfJ/ManYhUDmvEAUXwAnHathUO/kTAebbFIU+
ZhIEcPmQz3Dj9LyHOyAB+8L1V4Vb0pd2tcLEnKW+m0bspNoNDx7r5FRiS97KMPqm
JavG5Q2dWYNNay5rD2SGbRzxFho5ecBn3ltPUHK3JAiP7iNu2JwzAeozojOWo5ZV
jnNk2lA68Is28nhzWHmUJGZGfMYl6+CIxUN6qWijwKZymceDzuvN+Q6dy2/R6Am6
XHDqaKUthFounVSfFrPHps2KBLymZBoK2Le/Yr0lo64LmmuDZFk7rPX/dFi5+3dQ
0RRqRGf48cyNLWy7cAgSWASPePGsqKlau4wTI+6aarrTxOo/eVMftqcabUrllALw
X+BaDhNzQzm8GFYmmTPBx8i69GUN0f8r2XtwUvl7xZGn9QFw1YdM0HlKSb6U7eCQ
h63pxnyKg+mgR3ty0t6YwX/h1a7UXbivyqDEzoH7UwOlxSTiTPzcFmWfrS4gj1cb
AMVF9sWdqAftiR0OTz6jbMaBG9uyxDKPt5cEuf6wivM4rUNEkHD1uLktudGXZ6Sp
Szu47n2g9GN/3Xrd/ofuWX6y6d9XvZLHEKPsl26JRpOxV9zarbAbhrwVVHj6xjwR
gJFvyYhOn7om53XyHc9oxWRJULSmZ8wIZ8XWqKc8CjLmepFbtHSrYwbbxQ5PV75p
gTtqL15y/1rC51X11ue9CNTmoc1gbpn7cj6T1QdwMdmkoMHUmilUsg+p5YEOXefT
bkTQOQt9yO87g5Z2XPh+D3tYZI+6Pu81lxdIcjAaeWI37SqyuOA6Vwl0npM/3ol7
u6C8pJSCJ0U3y0UEdO2gNKncguBFl0/1Y1tjlPtSb9AHJuKrexbqj8dqPKf5+Doo
cynXY/84jWIJhMlwF4PPRXBKQMoECDvUxvLUr8YfCErv1UL3KqwjqTxpHWnmrW7b
vUc9GnayCmKm/ALWRxI0pNyvpyqLOSXfDcGc81z0b5LIWrcvqmrBQQ+Odx5z970H
+vK9GFJ0tMd7AgpNg/PQm50Bj/5t9JWwuZlz1iPkT0yIsnFHGeuRPkoc/SK5wyQx
riUNDiZpjhNdAzKNHC2RffJAvF39Ze/pbkCIo41kvhA0aUo8snN0Hiy4gLKaaSkP
MrC+pUa1ZDhF9bzWDWEulm7BA9sZeUWLU/xCpsKzzVfijIgTQu3zbqs/RKD1gbL9
4GZsLamoxHCKi74jrE5O98+pRcRWNh/KUzU0/1XYpqNT2GS1xSdQNMsnI6WwXzJC
MpZ5doPAYTKU/VQLLEgYqMrCXKi9vONhF5h6tDfWlF3+T/s7YLakNSjOJSlmixzx
r0OO3PT+DaoohP6k6e4A4OGkR5AGq1cKQaoS1w3YGN45fXzIU2BaGbgwEWxWXo9m
Ze+KrV7TQw+xPE3NmrK5efspNH9LOt2At7gwidNaZMKcOaxRzXITMwkX6dairWro
7sOVEElEUEsEaEI+d9d+pmFVXFzpLe1RXZUPGw5nYhBmcVMXdO9KwK3uL32EuviA
JsOUURY7qjwxwZtsHiChENmY2tDocCBqME9rj8JP0XV5jIL1+kMJ96ISLuz2PwWS
TNxFpZKLHKvdM8/+7AH1vNlPimRkjrYyFLg42OJYZfiLAjfzINtyL/TAdS97wfz3
GgUFyBXh8BaNXIpynqmZEVE0D4l6ZxGvrMoehcuHQnFUwp8Ol7Eyawbjw1bxL/Ad
+O1c3YuAH10BGZKaDpbl6NtGwa3I90IDLHUlmtQB4w9N1Jxsn1YLxG3iuxRT6kLN
J/jf9Kl1iIsl51ms4CFt3wKw+UWOeZztjoYfkVr5nhpzVIUFKlN4mVgi+2jWTCEi
qI+gg1OdOMw1Rq2jB95ueIdc8rkuDNCjgSB7HF/1oD6rPpIfqA3oq/TprxvzA0ox
LeFZRHtZgBdAnchE5ozSP6+upOsNGisPg6np4zUp7ZUfaWIK/eYqCDP1PLd0zPxE
yz91zDAFhk6FmEkhdBY4nM9qC8tKL6gSiSyDlyfcrbrx+/8/seTDl7d8bYLSar+h
EYHji1DAN5tuZf6GelC1WLB9V/0jG0cVQRZAEYe3yFTk7PgukIkNX9EzXA2dq0iK
718nV6qNXul0JdY6lhXBgiRePT4076jLBJklMHfg/b6xep4xohMTfvs1npijHKTD
YCMe3O6qRvvG2XaYCYd7BFOS7FD/8eLuySqB0hGz8SgniMPlMWWOU6m8GHxF9ZVG
ymJm/nNtSc0g99Yu50nXYlMCXezACW9ypIn8DiEZnDnTBGVjZPW8Sil/lppytdY0
NiArYrujD5ogqO3Y41LDKDj00ztHhcQBZatGsekLbOnY2QhAgjYydb5v7Nq8foas
ZNcD266BQMu/syRLaFwVg3BlPFrB3CInS9wHovxRItkA5CaDjtkF7X4hn0V1IOYa
7nO12cEAQZY2HPmTA1EDb3Vtto1+BgbHIxzzG8C4oSAOHOTRnBH2a5y0uVhYjomN
DIX2CY06PgnJ50ctSLoO3/6jOtG6ZfdjXrFCFPMmTKdiSpJ6BDYvBAdtX/RGt/fH
f+IJ0UJWpJFB1otaxM0BZwFHOoYbSq846SNJWXmU/qdy+Fe+F2wBijyCjL3ikB4G
peE1e86ttPImlgJapS0NKQbLdBqfLCA0mMZApHe7FtodQj/hOixIXe8MTXVKn5ip
msYPJ/ranlYHqGGXoU5fgFy1GJbkwmx3m53/v0e8QgGzXYKkpPkE+7mUmprprVqP
Ju3sZK9G/yawkwvUBCTzZxTBu73qlx4297QxCSOOdv66lthJ2WTw5u4IjodshNYf
zNMWos0wO7+l+ELQNVvZhCj4Fjsc3lHmRhDclop6IWGIM1kTuqWrEsi4w6CcCXVu
cNsnmZsZueDu2dP2Z4aSupJEcRjiJsgFdzzpVP/yEjvqalDrqk/OGAcOELgFiLRF
MXItirFFLfMovMFzMGhGmx+nLQeh/8JpY2QH5uFERBcdrU6foBhG7NHGpMGpYdF3
x2IzIoNgESKitEU2NK5YuFlCWUOEznwK0rZXBWTxpGz6ebpsb1RBDpXafimImT9W
WKLhbwbkFcGg2iTpIdTTMUOAlIWcqdGAyw85P9Kc/SW/ZcDT222SfnNRYb4qOL75
rXrjfnttkH8xD4DhyBwafKWNEUxPm8+jybZlZdzoUhnwVUcO+9sh8HWlirEE3gYh
S1myBVmIf+AXHqa4QM/fee4Gg5EI3gj94wY6hRx1EAn6qh+4UR2ORbtRG3wVJx4W
yCI/YwiRdvjjUV9tYIUZuOp9HLOoOe6qJLEebL8expEO0e2W2+o0OvAanc4YjO+u
j3+CiUR4LNHPofekYWtIB8kpZcLUp740xe7e/2LRMOsx3O6xVgQmj0qWoGZ1Pgke
dr/UREeZII85z4W46JofLX8AUuqqQnkVy3L6G6u5m4jc/LKCGWcRBz9UsZRgmY9+
pKs3QjzV5W2P2SJW8kW+K3Jyhf4XzNsgCTfAtEodT+WFdOQASWPdFqfeBdcuI6Wu
1XaDymrm8wRCoDLo8k1dblpXVjYAgHgQw8lUNMkh/CFfEO/RyfrOdStzjqKKLoS3
j7EH9sFzHxrSlBkr9VIOIPbaGEGxJqbho+viPNcErUconogYhwwU1szbiYd1o+5N
r5kd4UQTMwDlMm03iV/+ItFB28bRxyGy6s0+6ufvKC8wkVrSGjInvixfbq3G4Xic
r8XCJl/vRGGXC0wIERlxRpNH9CIw2se3KYekcvzA1VgzAtY+LZVYbUUAbFV2yU6H
L5wTgcJKuiqo0/P3ajaFkcAX/OFwPtMz4+vwir29t7bS0OlpHbxxEDtQVQBrsIXh
tQZxfIITGMm1WziA7wcfn1Y8MdXqh+4oogs7V+0f0613HczW8yluaGJBotojU8zM
XOEC4TF6j7sMnL9MZl8PNimAF5odD6h3b+58w1y5M8+noxOjE3tn5YOASaeuEBHl
uLWazLSCLAgANjlysRI7KyCaLwTzlQWFCV1c3Sf4BLDQOMmfloTo27ih6RIAJLQ/
yAtXDkNpVyrbfjQVJ1WRCWYVmSRbgovoc3y37iX6E4VFap8HaGe3B2goGny6PFxj
2ORMLWcCnTV0YLjQxc9ZYRERUHf3/LHv7w33JsdRPITIMKDUkUozyjLaRkcCIyna
KhMY6p8C1L4sK0lFgZQotoc7AQ0dsez4cUlFgTSO5ne7rLJFQV3n+MaMKdCLNsyI
iOJVlGKZTxtLpTkm5PJXsfHtC5drl+OSnybV+KWB5WNbPxP18wY7bB6IS+oXDLue
AWdeIbjEChVhkohtt/jRErGy3Qax5nbzQ1oCHetNO14DacL3Zmt/4rWZVwbHS9ie
6sObKcYSdwthz0monFEJUBW/y+5FjucehSbw1nLa7UuVz3ixx85bFSLYt8hIMVLu
g//0BsxtW4YiCfCzL/g8YX1kE2Q+cmfobiM+RN/ZU4Q4WFprzjkMEHhsvaNEMS+v
tW5UbvdZ90brVpzFTbV06iO2hnxOA6on3f54tQjQoKARdSfZLdGXCAW3D8icAwaF
c4NHjcSbBqNUjCl7xmAgQgSrw8DKvxDuaxYPa7X3zjyEfTP0X+92Bm1RzcKvOesj
diasIIHeLlu9LfWZw8u4LL2LUPw+jzXpKJKgJx2UeQ+LW9bgL51iSv+hp4Mhz0ne
bjYAVqXc+BO1OeGOUZtBA6R1ZLHoTRGkgOhSv+7iIr7B6oJrVZKhiMwNfWcKeOQ0
MZ0XBkTiXNBZtkjNGQ5MJbL/o0mNmjEuOIBJG/67dBwy8YcI6KXwu9ya116I4rM9
eJCzveRmKoItlhnqLdd+tPPFTuwz13bEJnsjBsgGJsXiwneruqEA7DoIbfy0HxzY
TyeuXOCqdj8T7SJWYyendBdbn9enGmlubDggWe8a9Lk7BrovMfuy5ehoK+JAZBsZ
Q3inxMV/k3vo4nPbQQvqbN+b2s9piRdoEkRqlcI7aGQXzV7Qq/7Ewxhq6Sf/YoJN
8Q1Hy96OxrNn/P4au7E/pBIXW/G/uFEoz8uI5ZZrEysF7G8l4oMgY7t7Rpv7EMwR
FFzn8iSHzH4eWw32pk4ABCYK9D0sDQOhst+ZRyEyAxf+eWM02fybs4E1+NFdb98u
FfKfuLLCw58uspBohMhWR/VzSG8gpGXjQ0xHRYIqt6/PcSaAsSjTvzpKSMKEkkeu
jAJhnQLWNV9qrq+j+2ioQSSiEaeAI709uytdUyEJkb9yyEX6j5Z/aODY1SyIyCBO
piLQ8kLJvbnUkgy9z+epfQrtVMZgy+NUordeGHLLDKsAAGIpqf7lHShsXCaPw27R
RSxLr3hSFA3jhJLfCxWYhUQCfSALBdfkBE65PIaW8Ia+sEZXfw3DFV3KvJjmepvJ
Kpo9PdCJ8V4xmdG9xDy3Re+kAmgJqCvNol1DWzwu/vBWsU8npECOcUw3aAT3GJd3
xwIwc8Tyl31aOebBE3Bk2B37KPjA6oXDB8nJyxDfR2bb4NOiv44bij4s2kf84j+D
EeA0R3hBOgvHx5EEmC063Rmjc9reuRWTNwpJJdpoyl//52bFpNsRgEYO8Ud1gFxg
5ubY/yTUQMXTtQxzD/KGydfCL4zXTHrjtS8HkB2IEXIGw7Y3FCEWu8+iLJtIspz5
jDeoczhPtTc8ZpMb17noy1b9pAIHEwMetHJM9wVtTb6fUwN0MCEXZYU9FZ4qL+G/
bliYHvKEqXZdvwqNd8TUkf9w5v1Kro3xYxs32j9vYdOXrmvNx4RlvAwPXCCx7JSY
2U86fhQNpewF0gU2aeUIUuRlF0NRVp7ydTbz9woufSHkIo6HMvj8MoryY7cKQLSz
ayxpwF//RrS+afSTctMKe1ZKqCtIBuW0k8LO3HCQ9Z5rKaw3kQ0ZOE1Ss/68POjo
KZsdjMf9MW1UjftP/9MZN/EMl3/mRKG/X5eP784Mo1F04ITL4j9Zh46EFcJKnSed
kyEOm3PDMXPDptdV6Zwt3z3pr6i0b6IB70+p9kzjdTODYSjowLATrm0ePEJ0qaCy
FnAxeHVO9vsd0YSW8tQPr5tcsm8tyADZYmOEbGZHvCAsBtWAj70VE6jQ5Zk27Ooo
/X61neoU5NcndgzuH5CJdzQunEuXfT6w7bYFVfcQbSJEXzeXv5YgOA++0b1yztJw
5Ef8qqpjUa9KA0YAT0q3KR+1BbggqDGVu7NPIT6sc/rvR8rTkCSojG1yZEeE/csP
VagMMVjAspz4RLCd15n23efdPX205yGr/970Xtrhih3Rn/mbVXkQeIcDe4agQ1b6
k19IRdD4bMMRqfBrQSa9L0K9kLvdpVGjWTLFvBg8UYxK5xhm0y+csMfsLsK68gTh
vM93+VEsA7jRLrK8pKHKxHCaoD7+0IcC05IhmOiWUcKMC4RGy50jYyb8smeqoKZ/
L2EHtirVxLMMf2Wl0t3hcaOjZeLVCeYDd2oSe0eq2Kp2byMOs6nZUj61Pz/dmpcn
hLfsDB63NT+DXTRa+DxAW5atVf8RwsE/3pkqeAh6XEv3we5QQ9WgyVEEHZw9bAU9
BppPDQIIb3PR+cvTzfxMLowaSUkRWHhKvOD1pvOndO/o9fijmDWcd9Ty4FP3nmfu
qrHxqxEfliizF5JOCswKizh65pHh6V9nTP+GOx5m87QRGDtVTfJA5hS+SWR39sIQ
WVmjh9T44CTQ9yt3m2uVLwNYz4rmlWnhhAhxepvVcO8AIHKmChCKploUCGCCF+W7
nF7pF+Cy5mEUiNOAi/Xqxy3SeXYzCnsfOJGgce+w1sstg+qUF5WNeJautc4ybHTF
Llzr2IHoydKRAdwpqR2l1M8TwVIcZoOiX2pYXe7b/1anTtqZoHShfCuDIoBdSMsE
UFdVUeZ75w5EDqm1MlHXFp9m5AEPv76nxk1NhqUC2KqG5vjSVkwiwjlmOBlXIYh0
v2bGx1u1sA3aYpcALhRViTxlVI3wQL6ZALvbyABS/L5UwZSTd6aWf4T1Uc4cT3g7
fJgMCXfF3NprP6YbCbGkoScQhMzVpRMaIR7XDFZfA/xuhEJtvZWoKcPnM9d5m/b9
PJMbo4o0v23xaDpgmWIAlZ26R5uBMp7jT9zxbBADYBJR6PahnPZ3hHhVqsqZMHJm
fW+rQJgv4zr5d2TgX1dmqSd7hxBr1P7sRgDKrjaE9UUxqPhAY7xq9bwbqOdmJp/8
KRPN4TixCrZObmyqSNHoumD2waWpjh/EhK6G5v7H/4zMQk/0qnEwIQRozI7K/nsK
8lJnxWtInZGCJwSfavEzv/GEuKpXMgVUvVm3P1dGUSWQqq5Jx7CDVOQBfQAZfOi5
502iPSJQ1MOQOse3ZauvehDUOjQcKRrlopN3UaLE9SIoFjiInKB7w/SitsVcMeR1
UM58KIcDUbL2GFvYH5azoFY3RwN0LyesWQ3jdvbNrGisNhwkpQdh6emc7Q/JxsJ+
93cgBFeIWb/k5sb8ClwUIsCe40q+/714kcPorvD8dESdZKICQRgh6N6AFOULCIYi
eNP0WJbPeXFFyIGGZVJdIDECwjZp7yvdSejFhCUhFyGa/QVbVuFjDbDUDt7NOuSE
AoWHSlbpraO3lMpyMMXKyPHwo1dRCfy8wfgB53WFrAuJwS11mZUAARUCQLjY2q62
NSUNUUIc2jhF9FweNmR00JQWbs5C61+66GPSUKKtgz5uR+tyA2AZVa3LtmOXTsWH
nrtfIWd/8ZVKEOwMeY2I9I0HOwbFTfdmxMK4fHTEP9W4mbTEgMtVH0c01U+vL5Wo
JCG/NFrPIwSpF3wyuYNACGQpMvV/OFfuPXaaK2f2mUwWd1mshkHwv8ohVqQst44k
Yg5ElIslUYDD/FCex3A+fvr9DlHRJ6tTQrurqgO/TYXdqt1+aNB4NZviNXa8l/xx
HU8O1M0nDnjse7Eagww5m9viInZn0gWzOrSdtK98GW8xseBCgMi8ZFQBLzKO653D
5lwXYcvDRBRCeZyRxTjAaul3Mlfmqcc584bkbqclpYg+R8sxia/75hI4ZhyqsvfH
1U5momzRnmatnhZTIivUMwUs4QMEOG0NOAapp19iTICkrgA4AxU7EfbAS+wiRUcI
m8ZqPt75ZSp9Nnyw4q6pgUZBxF1RdfpqYBOC3YKEos3ocAfEKBr6rxy5SXESihEL
ERHg1ALfylSxuqvKRt5tyGtKFJ2571ykUcGIwoHL47hiqs82N1enwonbzBTiyP73
ZPGJ98PRhf4qhyGrnzl2MpxTWGxfM8QVHp2emY0kJKG9BIIbHFAjCr9zlfZrOXhF
Y8avFPmJTUXVMFlFF0Ii+llVUnxmtoZKPQskf6Y/kBDHtQ1GPbVt/SwszXLgyETG
51ZaH36WjzW1fT8ptX0bHPnNOGoGvwvnXMYGwybsmEnikcfH5cjUMLFkD7hWCRAk
tKPl4h62N5SA5GCxZyCoMVHGy83q9zuc27oI/jZZnXrYX2g35ER/ceJ7kzGtaxyQ
qF/jmimY79Sas70xFaanYGUk0nhdWaUBmWa5DZszIEH0ZRCDno0QkCjz1GHd3J4j
EXWJq3RUowRf3pcTIc2darh4eYOKIRytsP8/B4sIDEEM/a0W/2Pho3N6WucGtK6k
KWOjY04qbCIueuQvm0iH7FHZnrr3GNXHymCPz8VW7czb0dEzQqAvzFPlqkpeJM81
UspPMie8mm3NptPl9RxAEVzTo0aOwyFIecrs+4wG9hZRPPAq43mdHmSXgVjSli9s
SR92mSaQGTYFjWM9c6SaaPneG3jnya3HXMmTeaQt4uKWJsi2kETGW7122ww/z+qj
a7WUP81//7eyLmh4uJcLrC8bBJYTNh8GFJfIoXLnz7Iavht4fZmGPEslnbRtKY5S
0iz29PwvF0Ijm9ZqZrz2IVdYLNt0keTe9HzPS89DLQ0/pkFTnO96Xo0ooxTqiQND
K+Oqf+mZHyuDvWjxGCOAX0q/NQxKc6PKSKNff6wDfEeBJNmRkCg0wZIPZVTcIa+e
AXrOhiwX0VOStG0trouTDtbMuEMfIdXP92seUmVxD8QAYLYBDN6LPiepkAyn6o1K
dsm631l6OgTLQY6pw+Cyf3AsTpUiAOfKgFkqbgy9h0YRsD0BXXsPIX+dGfq/QEhw
9KyXdoi3ZEaXx3kDMxSfdfC6nZMnEjOCtcrkUPZ+YBcTkR1KBhgSx8WxHb56m1ZJ
8K696jeLq6v2JNK7FSX3tfHIG0HF3sGDQnZ1QdvapMtuvjnBwFokcwLLt4iSA4RE
OMlfNmdmKjYBtIMMoR5RyKMpAagGAVNRN08+UHKqLzYFqpvjfd3LEGSUZdiLj7t7
1CqLbMdYALKmvTLH+Kx3Zgs4c61djr0mtWjT0aPur69DVraIgWVCdskic9sbQgRM
r6C28pI8k1wYqkEn5yed7wRy3PRK8GjWoWtTaxR5wk0OkcNy321pQk58E7VM3GUk
e0BWr9tXeeQBjVpceQucRqnTxf/6tLsHm/hU06G+zEwpMCvP8Lk5ozpKSY++ij1d
hC08rX1St5K2QrTDUQwX4w9G1/tzSJBTFN8H4h2DGqHwMphUJkG7NocZV6GKU13B
Ye7nRYkG2KjA0zl/ytJiCFJy7Vy6LI4IgL4iUbqEASfgIanbfnlt4i2kbAMOi2Kg
d2yz6/EEHxlO7Q7Uj9cADQB5R5KU35m3bBQU4AvjVz2INLziBQ26CaRmPw23toBO
HBYXoJ57En/p3QH8EHbOfV+zjcQpddocdjMFu6NioQ9W737v7tqarQ0x+DelyTzd
hlmVepfsL6L9Yfo1s2b2REoc4YLM6OkF9NrxXgRWARB8fS+IHlF1bMJO2AflWbLf
HAgnfobuEWZlmRkCbfIEaGcAIfPoD8LHTunPe+LizdXySafG8xd5ubyYTL+Qdv+Q
LrCLaFnxWPxTH0E1Ptv2O0q/Dfi+vbid+XySrNd10xEXksm9TkniusSvDtFJpGKK
FbPxIeLD1x/m/ScaZaJx+w/aYDXKkN0ynPwf3YzBOpgbOw1odNx3B2Dp80edR3Wp
W1+u/eddGiznXRm5i9nTkgI+Foso5u+OXYOKHQy9rlquQxKLomaSmKsnWAyHruZI
Jvxc10fcZSBCfyYHYqa4saWphtoXeSHrbB+eEivJ87NCdMCv0x6+rRCOorvd90NJ
JIC6AVqgytgCulModyRyM4ypRYUxAL0KtlUlkNasMkG3jqQCHioyeJEhBZwCc8rH
H2AlZiOW5erhrw8KVm3Qs8H9YZXTPgJIE4h4B+i9vmZ0leorHU69hBHWThTsc5ax
ReNEp+Fnpj/D8j8ZQhMoPw1manExTOytNBSwypyU4C2RXJ8nbIhnf+MNpf43fIB0
8csXsb6cFCxRLSkKKDotrEgDNvIhhecnCPiBCIVC5TOHvxjTqG5uxqbel1mXLhS6
yRokY9zjQimGQKGXdWxB4Xg8Q/GBVjuwhlgpbC0eFgukVYbyK8nIKbF8R0C1nyhj
LaVAHhPR/1bIgqCIdM7xLz2gTirYWlzlCCNz090JB5qcp3zG6I/6FPqHnflXd56P
6P3WL5ghEjPC7X54PHaAsGAuoZOjohluzUWrlusUlSg0gEvB/3xKZb8VCK8nTB+y
Vr0MkrCZNcwfBkfOq5KJWaIGpogMddRemV0oy6DdoYr469XgZeUO13q/MBDP3KzR
de0T+matFFeO4o60SDUwLIIu9UTfYpEde1kwPajrePkgAYJD22ca5CcDrsMmFARX
bf1SVJVwR5ZwS/biJ8Xc2W7ZKUEB5hIfiZx5ASdwAQdHDhEJCWx/XBdR3VLQ1G6x
fwLMOI2u9Sz5VVFW8QqzgtIspRAxwG3ZBDOwKEFVRtju3tdc0hRXXIvhlzfH9AB0
uXKQQW7v0gebXhh014WuKJ4CIoUXtW2MrdX3QvJ8ENlr6zZl3gjCpkMiEIEwYHgp
lhX52sNGDNauTuy3brTrgm9GRRROoc1WmdfEy50UU8cHqLm3h81g7x8+SoYEt+He
d0JJYLpcVboQjOZXO8fBRWd/ZeQMdGS6E13Kamo7mvyIK0rhGyucawx4JKaVh5Op
7b31993skVzYV+Abpfgtgqcjg2p5wLD54LpK1eDNsD2xXtiikDVSuXp0D1qu1bmM
ikUnOE8X4BTGYuU/uV9KuTywI8TT3fidjHEvwcQYtr/1zaFCdu9Y4oc6f0pIBE7r
QtK9XatslnAL2yGY0QmLGeD6T8xUfoIEPcH56AMqJrZnM5+L1PWy3PnNyY2MbQbJ
1n9s10ox9hYrCCxJglWieQMYqULXabzPCYMGGJOercKo79yneg9M6D89nIzVbeCO
lzLpNHr4LzSHAQQRYBj4UaLDmjG036ISi1FwfuPucuV2b+tD9k4Sd4W/NTI9/84H
tUF2UmCDjIGgvr0X3GVf0pEczNonkaxKmSOF8noa54YwORRKoaeu3lRgK5UwVqjL
RFaiaBERMRUk4KH3mJ1RV5mfrvXNNuhuszu6LV8SEKD6lHZm6+xxyrbS1zD8PpxL
kcKRib7fyrfJxU8lsEMZDsvgtPOw+PG8MnNMOcrgVvZe0cD9HVBwXMUxCkWt0xMW
ylZPbCBBTysQIzHcoEio5qMo6ZwpndkReU2m2do7HQqzHxoNGsNfPD0vKd/kY5Nr
kKKw0p5SURRn0J7CiJklcPiiLFi0RwLq9vLC/y2BbqeA9jHNAwTopM1fdKylQ+2I
BxVuD7vesW8Rp0NFPtjZU2U9V4aVIYB/OmILnFHk4I74lgKE/5zs1DjoItFI4zDk
g7ZdsLvvefUnR2hkm59hRhEYbiVg2mFQoEWdy3p2o0GrL6qKAiedb3Prztb7VZz5
Fz3ZlZstpV631PROAtJbMCPnPDda/UuYt6WOYzVcnr4a5kKjwWhHaqKa1VkLoU5v
TCU28GUaB8h0LliTQC74bvho5AuqeLOYS0U6mXCEBy6Xvj+5T4C43QH8micIbgUy
w7NXHvDhV7pu8BcSEsI6vYjCY7ZXKU0TEPs8GwD7ohNRmFLiXtmfo/gK4LGHsyEp
Bc6EiBeQEKNBQnH/UMRFn8IQRrrelpXK1tMLjBz2EkqAjAXAWl7dzZ+8Fs5oYgGy
DHpWPpLg5maM6LzS0n0c+BCk9EWQ/korI1vDvQtdrLFgwWh8xftrncbzopFiXlKq
7bNiIaZsEryedyXP/DVe2QD8igTmBurUs4GJAJqjF8pcPCM7c3mnpkfAKxLJpon9
bjBnBUGqMg9C/nFOPQmCYZdWhXBeJEXs8Bc+zMR/CLXlmca6OFz5maWoJeeiMvb3
gqFb6ULqydcq36by5nCIerTqgoTQm9SfSXe0Ebav7QY/TFlqVLmrICK7tAOayovL
7Y8d4i5eaEFJc7+jaw7dbPJLz99ugasI+Y8ViywW16vVCNrG/2Cmok4pK1NuY45c
1CyuyNcukfvKp/fFsnTwUpeY1dw6tPgs3JlWmJsozPurxWSQ6xu0q0i8dNwIsrwn
udJpvh9Rtecz7813i/a8t9pTMGh13YZWu4ScjqKIWK+20Nx5oRBzAL/7h+XDjvOl
BYw/4DVzrkG2IJHRHC39pRz5YBc3Y4DidQ+8TyTBwelGh/WSKnjWO56b0tjCsuzQ
I96QNPmes+P3+Ddq1Uz1ekdDM6k2R6cTwfk5ObXaP6jSCH8LGkqXSRpObvGz6FFc
6AQcV6lqCq1wu7q+NilxYnPB9aM8OLazWGrohhQGOAukoVB6ZVyvDZRiQ2GxHyBd
n7/rhomQP3IHaicEgqfBqAQP7+vQ7eEER5f+GGZYh+CzEcnNtD0Syb7dX1NQu5O+
KPjj/l29i7yxnp7w3S4FGsE3NraLE9444DpZZQyvUQSyCpmB5C2PAUn6P3rqmn6F
yXV+234dOy0as6hZt6J4nAEJx6NtqGSy5KBg6aB03AQ9pngwXuSpSeqI2X+7GW5j
1xU/3siXtjNYhD4MV7AZGXx8EkEbK+67w6t5ovZzQh7MefIn5mYDjFErfDyjrclK
+QDCYB+lr2Jowjy6F1km8JKrdkdRbnu4ihD7rQ0goORn5YQBK2uUY337AHtJd8Oc
5xgRvBa7oF2e5/X7ov9kedfZ/+1uvh2cdx2XKAE5lWHmBDHEjUJbJ518I+IdUd5A
q4X+wi+Jz+omnIo1TtQ+lC2w8OX/Wpw8FjrpcB2wHoEBdY/+4vDIrdy6H4YUFn45
ZRGdmKWe9Kl9pcF2lVa77PmD+kcqwseDtYDIo8XTSi5OquWUgmneB5TfGI3K/R/3
0YMkP6SfAgoLr8xUYQrUvobg++2jxx3IiqOWyxDv2QTVAZhiK150XNBxEoPIk6zc
H+5fXXWRMu4mj641yzVEYVFj9MEw6sxE2mWOSotbsV4FLo6r0Ar6waRALenw8YN/
yESxKHbsGOKnQi/zcLCeuqOS+569jhzucKMIQNa0gYk42k9gwoaNfJLiBE/gcoll
l7Rw55SkIgLuupnTkS40gIFMQ50wEwTspTimN6A98pEnjDOJbhzuicQlcrVzhaiL
igzU1cHexTQwhGyhNdQIcwGtJcYNxU13pR03H8wdVIKWJXir84Qaab8ADf85w5Wt
JRqGcytYqKQMppeNQ3lplqaas37mz2HhX99azl9YKGn1j9K42o8AdrCnsHSonbfx
h+3tV0rpPBc/1nx399BEIsdejD9wQkTxOhVsGjlNkIetzbHMtSXa15mWmP2AjSu2
k/qUK8HhCO2zKtkOeILgN+NfyPXHwU1sW6C6l8a1e8i7yx3/Bd7TnGB9lFIV6XWa
sOz5Xkb8Tdwr/GwiVjsH5CpuFy3SLpLCpLi5YAZ0ai8sIvjfdE1O4OiplfEn4y+O
tvqEzHLCFJJVeiEAOd7iW+oGQCioPm7THVxrXokBYjaYTPDMFszYYPBMO6gpzZrX
M4RCgZPHltyl86Es7Yqsiban7+V/JAjWi+kjIjKOK+rrn2BDwDQLoyimw69Mylvm
JuoxPxWI6qF6pd2+aKeUbTFDtR0QlGeu/PnHGOuagbcxfzV0KyAbf8N0NJInvkMv
EGWeGQyNJS7r01GnMorbDjGInhGXw/w2w0gw+mg/kjTyV652yxws5omdDDSmxL6g
nG5BnCLQob788mOflstTPc3mAGXpUKWNIN7Tn3t+Cq87fyeqLsY1p69feigW9GXj
fIFR/+ZPG/kEjtYqlaJizrppCpqeYn9UaiCQ+TQN6G8XLOVbZef6RPcvh20mCZCk
lQfxyZWTOjbiyd2pAGEjHAwh6M8fQekuZMZsuhJzTM4fOmzdfim5JOgImQTVtsYx
HHJkUJ8n6NyWx/BIPU+lncwpm7+FNdPg1GRh513dqHiO+RQKU9kVEcZV5cxOUrQX
h3tnbsp+frfDyPfHd1hz9QI7OwxiqqZfQCnlZxyqaoNa2diUO9qZM5bVBMG89ffg
dHckzdw1GhFeYIShpYABrRqmso5hVvEXdQIz96QzanthWGJeos1tF2qCx6aZ6P43
+YxI6A2eDYabk/4kRk2iCqLGzDXvCGnP7BVB6qEncIRRUjr4VIWOOv8pbju9Bjor
M7GD+Ee5/VuLx2minVTRioWKEbiidWyvXSZ2F/eKPb5q+I2EVBP0ZQsHa1U/D1Oc
c0FXPHdpmqEJxoG2EVohELy0C6eDrZHNiw+bltWRLguqcTJ/sgQvObC9tdHh/5dg
xUJ1YfVZYvxX/07hpUSQtw2e7RgfMtrW4xHZJi+RssVKW4+IBTVltrNtYgT8sdQZ
1u0LoHsaHozuBxK2uv0q+AJXh/ra8BTHfGZAI9qVg7ZIeRLTGPZk91VaP2wri1lY
ECNXeWBkQhFt13vZRzBaStZmRNnl9cZ2zs9tqqcBORxtTNRhAs0c6pXhV6DcSecT
B2DkHKcfKbUijqPhm07ax/RDTnvh++zhZmE0tqc7/xIbUqeCaWAw5/x3fLcXf9vo
9zTEI0HKKvaaQBAJAYIxs5xW0rvq+CXCWpmcYnWVSCscLMJ9zT4FacOiaUjATTPC
skXQ4hdY5Skj/3+qrCIkk7VDkwiUmMPyQ8zuRvnhheuruEJs65jhtGpBwIMb41Z8
JZLbRLpHI7BJBMtCrt3g2WNtOBTcPf8nTGh0nWqRC0csKePMuRhbZ50BJf/QFB6h
Vl5Jg+r2MRHg0WEdbk7Efba5Xg7QrIv2zjvGGDcVMG4g97OcTqOg1dYRxfxqYmvL
W6m+2bp8JeeBoXFdda+6YIBrCfH+ZQm+8SIHAsChW/vjZTG63ytPVkDfSs0oapHa
sG4VUL649g1ToUpDmFm975UpGIsyWHiIwyVNAygRC1GvJJorte784SdItuPzID1f
/PUJMWbALAduVlCm0Z6n4U2c1NHZypk3VN21hS2B/vuVByzhLdiI3++Ht50XiJn/
+15UJm3XQr6crmBAQ2rT1EAtKus7LD0SK56Iaq4WXXuRsyd845fpWMkT/cziUZkm
3qsWdv30C1545qm7HCTkiv2RScwW181nWSvwKCTzDuagmOpP4UYiyDvv4Mmq0TyK
jv7LbM4V1Gsj3lXVXMzNlsGhWMvtvbGiNIVXsNlbtbX1Po3pqJiTFs6E8cs+LV+1
is7lKim4tUDid1K9EQo+4RExDWC+FG1gV/lpuBUS81VR7tloPBwvG3SkHX6u35J5
qDjwBeIzzaiiBdJ8VuoOecZiFmE+9xwYht0e5LEG7JgSJ34YtD2nJ+aCdrrxPc13
v7hxB7gc3FPuaWhgzN/fOtwyAbEQRpXqSzmXoG862JTrzfYb8dfoXbBYDu6Tj5cj
xQWoPlsUdSfXplr3FjZ09o5ZrkXEQ7jOwR4qQ9Fs041GhnGKc66urmpPZpqp/XzE
zqXxYG204yn3FZIhUYbHkDMrM273ptyxq2QInrf41CaWag//MhHUbMQCUlLcdEaP
jHwjEmy/ZsyC9gAd6eF2RjaOtpsQIWEiSA+g1wPOv8S9jvZqWbQ21UwTzccUdzIz
7KdI5JVTbpl26HYrfqPtadnz9koqsfFkwxZ2yDR56Hq/e9llLBmsu2jEwPmNXTEt
RKUcTGyhf8FSS9ZGnCbHM87vjgW+XnIGXY5eIYnyYlVHHfTIDwcNq4SWYjSAlXKi
aaPBcEotBHl9Fcnp3QPtSN5KGqacwgsS4pviXYjqJhhFewaKAAIERsJPfOGVNjlC
YOMI51981y/zb1DUfOAqwqIyhxaBp/LyAZ7I4Yg89UvsYFZE2DrTRfd+ZYJgmisf
FvJnX7LwOmklpFVS5UnLjmMIHzC2B04wnvzhRVXTAlNhxJHIryZrITKtkCCbU0EM
9Ykhn84dA73vYXiiCJbgVnBkJLz49j8FEg3GTu+8x2o+/2MsMc9WqC2kIX+EM7/j
kWuyfN0dW71nqKSfpzRwiPj6LzAuYqw1LKp+hO2Dk7iPjL7OEwHMBd2jmOSKJXZ0
IeKRuAgPTHEePdZpr46THl3h6K0PeHer+doMp6z1Z6uMaykYmQNFOMnIcThbUjos
bFqko74c6UrO8suIIpw6D5yVgdsQfFv/SXkKQB3hW2cDc3XhJ9HYB/CXYwLFTrDO
m+7YDHYIxLmcFkBbkOsjAJfDVvH17WXu6YRywqPOYEu4S+Bgfg5H7vtEMoVlB8CG
b8B8hf//GA2caPumPad5e3ekeqJX02Vk0fZm+ygRhRGCaK24Qchu/Xi/bpm2lPgd
PC3UwaWO7NkOdWNra9y/7FJqNi8xm4cXDoYqJ9Lr25B40OyIOne2T5t87PJL57Pg
82WfsqEWOEejGEU/1nWCVfTHqMvI4pyTADXoVyNyQvOrwVH+2yxkdaLMdwlnDQek
g7dRMDwoqkrXPXDW0sQjoZHvK761t9jPr6oFbebydVe7xdBhfw/XljbNMmXGfd+Z
daBHMoH5JP+KBk2VYIDVGjKLMlkBFzV71b1J5cuCckfDL0v4YQ9nnKhKckQzZAiB
Gtn185TbkNwUtB804MXU/I3hisvyof6r7CQccB+p3YCH0gEEVtsb8rrPqgEl44vY
V6Xx9ioLv0mG2DXCFF/Gv1lfTVu8YnX6rT9uCQijKoTkWs5wPbM/OBrA9VrM1Lm7
aPsxh03Nz146Iq1lG5A2METLz6UiKyeH+f5axUPpqC04NqQHYqgguA0asPvjOHW1
yhRbBNHGTwqepIuLznpEJjOmcYr1P1T8Os/rycsFJ2bqvW8pqxttaKgaocYN6TyN
bwEOvcxXdEosHvbcF+xbs0+7JlUMWBUhLBdF9srYMhucsJB+9kaRkp3rOTJEt7jQ
s+dIjUa4280dLlWs5uwT4g1FUsxoY5MdfnOg6tzvl58sYnZK56OttQlcuAAXOIMX
chf2UXABhhR99Hh9/JAUyLzoKOWxui1/e412udA03Gebhdc61OGwathAiaz54tJ9
OLu2TojqXVFjjafXWKRa2rYa0whG1pFLD9GGkjv8zubJ6aJ+BJCRUqxP1kFP7FMe
cZPAn1O+AmIsM/Ya3yi/hQb1yyB/WiFjqXRIhBtQoJuDOMEoi9EU97cHMtI+hz3B
gUVNf6qui689bPu1meK5fSWsK2hCIAcKU2FjhtnMhTA0si9gCbPLuoy1DFaCIJ3r
QmBc9pVjnj13u6duTEwMIP8zuXN49mVPC5+kJWnZzo2xH1iehyifHh7rVgL4W+xD
Si6BIs4IO1htkKTRL3I8CgQsGbTvC755d8eMQmvx7zcRp3Gd024/yOPuqIizSdyG
sJpVr+F2q15zbScd6DOiQSe6QGkd26aeeoMa/DLoGRZIcGtleyEB6ItrrJTSYV+P
yuPQDPW8Cm0sQTABvOKF5mI2llsuyhQi0IKWUFwxq3Cw+u2e5TsbgNrSGBf13zle
DupGvu+1IMexzJKIPu5Drl8gbUknZQ1Bb4xbfba1O5VsGuW/TIjt/nmq4kP3kNf4
OB/K/l9TWo2jf7FBO2v8XUr7q2N5mvI6sM5nW89XR71CtA6BTv6GYTn2wPUMs7qM
M/o41TQvYmoAOSbw72NjQubOcKWPonvPKalIUHyPWVo5Xf32Qi7htB8rFp+mN/Dc
P2qsc2WLxBdShZSO1I4JF6rEZGCbSGGLdua3qFqAAunJ8ufiG6SbvVAZbMLjBj/F
3xH+A1tFD/EN+RlGCvAOWy79yfvOByYDs4hydSzhchSzvf905ZI9vpktV7Tokad1
vVQlzGF4osWR8SZ/hf8ym6Yx/UGIRxcIkA7wRCdxW9veBsD8g+aHZ6gysp6xV5hf
WFz4wzYiH7gbW/q/r7Kl/daxWJNZ5aOFLmX9qIiy/hIieMU9UKCPCznntIdYzStn
od7FjLZ8hJIyLRH4/6k9F0AI6uoCc5zVEs9pBWJsigt8XeMbk+FZgbCosNLONslR
Nc5+2VjuDhRez8+SkGMGjPnlFFpcE4/U1j8hq2XUSqJ3WPj/upBxBi7Nk31bURdI
L7ut7mSRKMWJA4Yxw6445Zy3bR183s2mAPZf12HapYVgk5UX9p8KI35BypV9vmyL
jChDs4Y29m9VQE/FF0ZeNEUVPLZ2VkzdXBlfPztcur06xa/JfKy15qBxEQGFirK9
cLz8qNTfgqelCuzyUvf8Zbr0zktSFWpcc/f7kotN4Ltu6WTWNs7goj6jMm6mQ2uw
inNs+zlGxjJT5Cr+5e0QhcMJEzWwIre720npLcL6pSCIy3Rddb3e9NqpCGl8jKJt
IUHhL0ixWs3zYDYRF5AN0tzUlzKGSGMeMQPtXrv+/jvVWEa+q6OmATqRgnkJyc83
nR3HEJNVKgk7xAnoJ+FJ54Nqi3vGX3fKAEQ4bE/K9H72vUHcNQi3237RX1L7rF/m
cQh5DsFUjfxpvcguNi2kTPTUyjRqVWMlPCwwDheMY6za7V4W93NrfMF43jy6PZUx
CL2cDZp/duGMqa3TcmEUhUvJiotAbZeL2+pGoD13vDOanGCshgGK9VtSn/mKF7Wa
xxWOxq3d45/93soOi/xYT4hcW7bxbO7ownV6lL4gvcwiFa3HUGPopGxojhxvqZXc
ej5eu67zSbqKIG0iXuxSMhgYNUhyItkSYl0SOhX7pLAn5K6PeQeWbLWgWpaHYJYM
1xrW7oFsQFa58YbLDXbZvMmlMrpkDOmOY6N6D9w3s+JcChdJ59Ps2uEbQAxh2GKm
ZbXjVdJvk5K6mGMZhX92u2LFuemdcpzaNxNYPpirWnkJiOBspJDSDmLUtIKfyniP
t0JjXks3Q7bVqA6BN4XGlbFF8zmYJyChmoPmvUKIZRvRtObdZelibWIoJVz/epC4
WAaqqxsRVgQR+ZOIDxzi8KJGiQ73MfxdkWCujgHbiLJ3RnKIVBBHgmFoBsr30kb3
NVQInmOZD+7nxgIzGbaBp7fxnQ0CzQDJ45CE0dqnmcHGzjckuDJ51t/foSTd1scL
hIGyXR5FljDa6zWCCP48LCOp7tX53SgEdW3LRagZNGeKj59iD+hzM83C3lL0oZdW
hDEh+6xxSx3BsGNW7peXd5I97BZTX1x7znJHS8jqfJ9omROWWtdxFy45OCoUybMd
DbAUWzSW63N7xbBCKMNnPsvWxdZq/JijAEa4Lt12QYmV2c50Qmzvmt6cOWBKKLdS
MBJDfD99RLmpxmTuazkFhc9yg0G+SxuugjSxCyy/dcGmrsEpCeio4P1DMZFtO+ZN
14mvJxHgwhSsPgsAnEeh2WhILXFTC2ySjk/r8PRGFrQcEnoS/YeIXVXHT4jmlUck
xIgXVVzcIy8A4zxnfOfXvhtKzyOe8/BjXtN+ODkgeY2ykTSQ7N8u0SZ77gv+PT+K
hcuv4ZSz7RCc8O4zg82muuJfLaMR9JzFKI3d0CbEvm7BLoggSGr54eAaNGnB708L
uoxrOdcB7KgJURZXljoBItHM7GzxykQR0CjPnAcgremIDN2I9O9UNPztytcPbG58
RBeP5oOHei/wvWb6JjAAQ3B0j0IOtjXpLlQtFJJ2B5eEtHzL6NOYCkS3sEcJQcAM
O2JAz5bMdEEiyd+aYImisNNnIojcZOZLVXXNKUYJjps9La4lM//5w8GnQsFf+pKc
VQMSKNbZF4RrVJ+tl0vkWk3VhRJhsH4wGywUmSaQYcw4KC0sKLGszXb6YwUz9QQy
8x44HnDVcrm5xGAo5/O9JMfY9EnLH+TZEuWjltZ+4/xWgsX8mxaUcYDhNRuAfdIC
sUepZR+yiJyWuIM7zitpb9sBu8JRH6lwQ9++6K3f02b2JdAkAKHaeE+okH4+hn5Y
45Fyy49h8ltVBBc+D9qpbFZtm0JzpuU6HSxgubH995lOB4PJHyHBcYTDH+ObrNsn
6GvalNWhZ2AIqc+YX98oYlWqw2lkg4cPXWv1xw++egv0ZMAHJUKXmSlj5+TWnZw6
CtarxudzLQS9Rgb+1kCxRd7yoa6SHh73IlhWspJKZGPwPQpldz5THZssaGzKGSNq
Y4JBGctMt4pfGmpBxSSWmJLrrwXcOYdNBcCf0zNDnlK+HJvWs6ahKAVjb3K567E8
nnndmTkeHRydnqL8RUTvwygjxwCTJ2lb5A5V9yPx2OW+hc1Awfc7xZclbexCipqn
paawrwltJHa8Z9IxK+MFlcXl5v1vtZydk1BlyfDMMafiN3GG+1PLmyluz0WmaSOH
kz1SaLJ/1luJ5ZGfeLp8yMZ38rA3PixBDxTWtJhKhYbCDKzta3hiTsrkAu7bk6ut
4KLbYIIcIGTFTUzfEmPRbb4NQ6MfZmFgWeNfVeFHpChNtvnHLfneaFyLX1RdBlzV
q5GtqyRYWLdQ4aqA4QmMmQkItH1iDZkDR7X4/pgv3G0SeVa+tIAL+O2Y5DJNB5Em
xu9g9DP4DwasrIBZLf3E1UsPELIGFdcfzWYu9AXyFa1mqv2VeT0SE65/mCKWEVD7
NTfx3qqcS4r6fo6Porpd71MxAOfpileyQBZSbfKx8uppZ4f8mOsRk8CpFFSOKHWv
uasjHeJ57lJ8fzeTHvVRIJlS31sL1Y/mcJG5CB11cpfH7uu3fh7xH2vVim0Hz4N/
AoC2Rrh0nfjGjdaLBbuQ9gElb+cqU30Xr9b1dyP0GQbFm/nCuhbtWu+5QkjPzAEL
LBoJu9qBEWr5gXRz7Q4taCaf14OoAR16qGZniUvu7wfjfLRKZEJPy6XOejuKY4K9
nqK/CLfXieCgO2L9oGTHCpxGvM5+L08VGAgzdwtJa778W2EmyKzYX3CvGUlSlbc3
br+J8pUo64paAry+J2IoaEPrGyyOAo0edysi5VFmzSJTr6vN+Ke+oeQWb8/O/a5N
eeJit5WxKQpWLmem13qcsIN0/o4dURvUiJMAgSk3WJCcc/a+8PmE/+erDRBOkAxT
J1DMiu7IoKEGlTbqE+PfABNXRLi+R+9hwzcGHSnvsGW2GYQzEPTks0tOtEWXK0e0
okL+LXl6jbS8KdVRM1MKXMJvP0BTo/NYOu4ZPtPZ+9pQGmfdVCdOHrZpHaaMQDuq
aMIalkDVpk2O5682BngPRUlbXhAASeZgEh6qo4x7ObFJqEj5sLr9yDmq0zok82w8
6Ni6c7JMU3SJOva5DclzfdyfPJ9XGQaa6ZTTznug0pIvta0+qHoTz8lF4KKvCS0+
sgweGOq3zn+3tSPoyV88Cw03CAAG92JXOxJJSv+aJCJ3gYRjFVhTe7NSCLbUbWX+
uds+qlcPNIYJtEv86QCbZeTScStGgghNIAlIcgpX0VzHMe2xKKX+8UJ5pD8eUPaG
D3onZXQ1mwpMuUSRcwBDEq3nglBSwsCNG+uH9czoMvyQ0ev6GIPfGk3Qp8yp9JGC
kvl52mvsC0EgaMZlKtmc+N5B32Ct+G+I8nsYv2luYNsISDCKZ+Lj0wK5ONTkHCB5
BbMAzV28AV4dAp06svx2fQUnK3lyObzshjfTrm62h+7z/m3jzl+BbKAN7QzzhuDp
R70/mAqi3iBPH1FTRkJlhGIYWHHybgNqByuH0Fy1HQLcED/WdPUpgxiUNQJQHC8O
zBCVGhvyVqibRzfSaswO7zJjOf/vd9uX32jgHkbhvgwl7PXEbWcjOFdJPJhmvPVi
xFk2CG2PZRAmd9bPQ5en0QG/aGcY9WKL9plGDhc8ol3u/vECZzJ9+NyeyzmjiPBR
DR8m1JnyGTOhSMdMSBIKuNix/qacbkGKz3bivzPImiynDZfIn1C6tpR1i3w/dE3I
3+NeLAQFd4zqtH9PJYKibUCQGeZZQRY1ptoWUiiPpHKa3EEZvg5wRToz3qVltW8y
tBYX0mqg+SvSctSffa49r8tlZglXN7dWK+ajtD6L51rGZRJdGsDJkxQfvnnLncBF
lVwl2VIWggHYJztnCpxEr+UeTOi26bKwn/uoKFClSduZfj9e97DDnJg3PH2hSqaN
JRjsVs/X4qoDn1DG++eOiccJr38N16VgoTytJZncTtI8B1y4qcXFMnIdiY4K4JxU
ZoJSpZ6dbWX5Tyv4hkV3kWmZ2YtaWMhasZ62NSB54u6q918yw6BTI0g3r5HAOF00
+1VK68A6Io+HWpIk9NWSSuY/UmKEHeKX+a9XvGBxouDRd75CrX+RHWIInlT4vIw9
+UrMwx+MDeAdGxDQ7EjEugOYBRUzJmFBxzIXdK88nybk1pqn5bmLxNbxyBoS/PKo
8wmO971zkCJHHbZ8px2sHcsFqq0JHag94hUhCwbiru7pZwSJqex4hN0Zp7Psur7p
82f8UHL96zT7XCMMVDtmj27Ky5nI4+FyYw+k5UjjKZbpC2nDMW37S6mamsgWOvup
BqWCN9QJvJGj3Yyt6sfmT9IP3DFQWw9vOkjDchAXM1KsgLurFchNqnOuIBr3f/8G
XSqpM3EQlH7ml2gAp04SxEwplEMMFycQxAKmkHL0SVk8ZRRwprTpQR96LbM0QTsu
X6+OWZzeOOj4FaiXG+OrFr3w9A4dPiAC4THwuRvrtB8ZFbnTWwd4+dvdfcCOC4Kx
OPzyQAgg4+5IS3Bplt6/bnLSPNchosxC/IKimF2PnIE4+w6FQawjJX99QfzZLpc7
ldmDIAy5f86eU1qeynunqHCG03+UxR+v18VfPlKlaxCB5KJ0RUtJB6HqnQtkToSj
dJpzspPcTHAQHNgnvdAlYYy2dQoNBKUUBODNj57CBurg2WHAfnmR1x/Fs8VAmAVo
CRxZDjCws+ceyfsbwF4RPrU/p2EPq1lR2oAHfh+61ghIK+Ay0sh0fCmZPOtcSDlx
w11b+HhfEhSNpTcsaGynaFHZNbywdqQMBSW6QfunhNypWUgOzses+9NUvWDLJAtq
3qKoSKJ3H87nhzyIkOnwrv5/QgvRHFsCNbnh/7iHKuOSHIKPy4DneKhUnMRYYMwc
fYsb6UXJIFvRkF4z8N+E8fc3Fu2EqjoUqh9wAjNcV07FIZiLLIvcXmZlbUJDNUej
APoetakKUt3GzSTIC12muCSXk7c/tY87DMj9f3CL4qma+eieE9zE12qc302Fiv4M
+zVjWn7+wc/sm08H3hyGXKkvixz/3uNHg/lZB6uM0fKE8NlSPqL8GVHnsydM2lVi
/mQexJQvDswuyX6tzC9n7w2Qug+bkQeEfy7x8oEZI8r6ASDcE5kddq5coz1XIvKC
USyAWwa0XrrlnhR20GLwcLOZZfyYr1uSOjiFScT95UUa2mzM2VGaYt6uzI6gaZs/
ZVyK/SKEvtYR0SAHUhAscBFUH5ujBs2vpajGpAYmPGK8kp2maKpNt7u7W1iOfE2S
3siLWwYJA8Vz/kDNPbQyoCzzGVWRSksEyrHGnnjZUq29walzwuZtnm80+1nlQHt1
83iWIXuuhJRDa7+0oyS7xIDotiHmXOUcR16e3R4YeQSi7FpXgA+tl1p04suhaS+F
EKEHAYvu0eA2aSAucMhkVQCvfHCDZWxLzMFpp2UACupJ6Lm6fMx6qGSl9BY0+3It
JEdtrFNYarnnrM+cK9NeTBcP9h5VToqjHTriH+TWLvY2WvFKEh4eqxC27L/ZBr1p
1H7eINDq98bcWU4j//wI4HGOxuOohnFdAjQ07+VF0K8FBOy/QVUiX1mkLnks3ECJ
/bHMhfmJ8ObbejIB10EVgjfrpSRfmSquPvrAOaF9YJ73FcprhH3bbznOSvNPJWIJ
IPtFM8hGTo39l2iJgyK43WIdh7xSFe+zyWxodxOKmv0siyP26i52mS966oUtCcUE
TMnhaBHWGgYEvpDYSaiuvRHacNQDMGyAMacti6jQY+sistL9UpYQuO7fqQZlccte
VSLhehNIPhFxsNQ4l2pIf/Ms8y1Ol+YrV/jIhNliGoKUVDJYe24sXJataPLX1IUf
8Dx2NWC3NJSpDHLeRQPxk7iRiz3t2UVSFBQsZiwWJSx+0S01SCv4RC9NC+HMj2i0
EeiVHAO5KlOqbphShs9aWN7eiow+KchY8EzLM5zbVhRDl7d+bDeEr0z/bgwX4AcI
n0Q8oP+siDR1sSAW145361++kIFOfpbieVxLEpPlD4m50K1p81iWOP/wDGQ7XpdP
d7cTamVHwUTQ60a69AF0+ZYAGi8JvzQox9CXKlMAo2ZyrduGuXpPukvMdWZhLjN0
xl/mkrr8ATqASwRLjZiHPQlUA7MuQGpp2D8flj5CmaTFszpesWaXMyuA8p3pz0Yx
tZN1EGPgDMeTY0wFCKBdQhmepx6HfHe3g0/jCQwnEw9GBrwmHjlNEXv/7EoRLtTg
OS8E1/WSEi5KJCaR/DZXJwFhMo6z2YBpzTXPUx8mg7Lj9wr5nmHy1fnfaXl2OmXv
0uTidXDCDZULlEbsZBcMlGm6zc6+jbfl8d3tgkGqnm6fWy5BqdP5H2shBBU5L1fR
Gj/n+qBIJYPtihKgqAy5/UcNo1cXp7pHCWUcPdzXavgCd7pn9b69zYvoJwYI8biv
AfWSfEm42NwErjYq7i3ShUPq4Q74Bd/6s25svDICA9J3P/DqOCqEArKfzquXCQSB
FGH5M5mG2jwtZ4JGjgoW3RgnanjR5MAwHIXGhI8CX0BDnEFNPgwuJWtXUCLTxXfj
ffuWCtOTW4NSPZxqTumjgrJPE43OkX1fpCXXu6sByReQzthudX9+wB3H3erSLXyy
ooo1WiSUf2Z0uGA0EQ1bQAwtWyX72t8ZrMR3Y3Vt5OdbgDauel/ZmzLKROhU8pAs
GH6hhwuk8H6xinuPIr665cPNbVZOgbvnjakWwF8ZHKZYdpo6xQUwN84ZquBwVkj7
QXlCkF67FYGEeASTwgQvwQMstx4KGYClzGa/5SETlfKzJtbOP5y3aZxIe2q2D9rl
Wp9WcPvx+3KOg2LckqlvSxL+kk7nsf1jFvbGym9wyz187Fpzt6+0vf+esNrLCNwz
dSfg/sWT/Yy4aI+8jCI+SAYf/lZHZw7f/2TmidfEAqe2MyENN7MhHJo52JKCXBA3
22wNL/quCSTkvZZzyCJ5JWnwrbQMFagYKmNzCN1ANnQwlpyG52J2MZkA2qmu4syp
aG9ktzpTwFE/0K7SSBq2cxpQL8VnQgs+5RZz7tWP2BFV9EWkcC7C5fhjDE1JofTH
fU4SyH7PFMtYehcAbf5B7BI1qXyZ1O5RX0saWtkVRQxcp1ftRDpCj5yQ2Kk3S0UB
+sXujRmds8IQGcLMNx0uM2xT22HdU73Co0IggAkE6RvgyB5UwRKAhVZM7UzVfxrb
DerTvCmd6CwQ1zcnllUnXEP1AON4C3BHkr3zeJoS+dWeHUllfDRnLnehT1c1fEe7
/1Zou7WedBHlpXakZyn/18VygisKoI59A3gFxmOstwdf8ODqmBUOsBRzYFuBS8zA
r0G3H0jZVlTQ0poXUsiIRHVqVctg7JnBsYKQHGVSSywH1LtIVA+mCNVO6/kvJp1W
D+Tkz9C54A97dikqRt8RCDfRcuFFy30wlqbghkmOfh+EQAfseedrMeMwA2vyf8VJ
0hTSeRWDrokV0J+tlEPA9RCvy7PuFdEK3Aaj2aRZ11k2FrBvfgx1Z/mtzRY+x5Va
frewt9UHDEGgghTgMy2v9Ssvd04JDzQGwTtN4/Uq1TO8rxAVj2hV5k83xB1/BVLx
7/yS7TIbNLYZbB6MQ2+qN7eudK3hXiuh9DnyoD8169mOL2oJsjq6S7UQ2KT1tAPp
pEvQ0HLy3aySpsq8tq40hB4VjWaYEZk7HZxR438WfPw2PqoWZSskDEHi7h0v5syz
OkW6GE9cSV5aQ4dBL9bSMj/ulze+qKMfMwDTLQdiSUQTu6uSBw2FgHnBH1LXz0N2
jdyNaJN7UyvSIiUoc3BA1d7ZwAPb4mgC3pgUuhm5ku0UKqsQOmW9c91fLiRWk8Gn
YxyfeKT6ZNkiN0r66e1Y9KMkDRKSvFYP4ku1qcKL2HDEEeffeyBFrTvs0f9PVjPc
czkiXd/A6rN1dvKyp7EW4waKyDwjX8nyjDp9gKcxeRa1oR/4+CJQSsCF2rl5JmCC
9/zqKWYIvoZ+zViNYJFYfQnOtcip1VbkqBY3xXvSrKnbtd2mKAJPOflBTCtrdJJQ
Y6jvZSX9tkpYynBaNsh/JhblFs8AoboQddOktfX5oyOeU21/yh46nUs+npUPdFnW
vAMBMqs90zcjCQEuyZr1O5LG2UWXVtTBxLeSv9XYHqhoD3j9JzvZEXy8832oKAAj
qBcTa99yuVGwxx9j+HSXj/43PFE2cHREyX6zrrz9uxeOgRCe2sx/7MvhvlgSqPgX
yqfCvxP8e+9/qLxmB+f8EaQn7eycm14lg2VVw85+tfNBf9ftyt8JQ2plnZn8nLCb
MoFTpFBfSNzCb4m40xKpvE+V3OsMcfvTsP5xg96bitz4021iEX4d7T5G+C2IL1DH
vEcRSqTxiMOxSeJwpcEMdWXTixV6w3vrjfHBFdo0L4jOodoydzYjyxV9MkRyxzm7
678MzwjF5oDhA4f04OExAT++/M6SCdjp8m/m65ahqZkUeQ19/g2pYs6Oi/ljLDZ0
dedWfUezIcyIJl6+WXqkWaUjkZWHs6QefCFaoRDVPDXq9HTu3etIXnFSQig/reVN
eAcmMVa4HQcSNLTq/cWGzJBYWL+JUJ+v+Ugrk+5wsmJWP1Z0jvFXYNQ+Qta7Kkow
IR/6RieGELChSqwoH9aBDu4+CCyszmkDDsvvHlbp+GMuopKwNBGy0TAjiI06lw0a
zduHXEHIPN36cFMHWiA2p2DjijGoywggKWyNBrWaFnKCmveqFmO4Dy4w/QtQxPbL
rH5hgXE5L9hC+WNQAacaNzC2kaJxlRU6iHBoRfItc9guQPZoUO2meVhUW63qe3Zn
BfrKI4k6tiUh3BWQihJr9kjrYUfrwwvn2AWp5iHyR2jrxW7a7MTI8y2a/9lbHtAI
+5QiXefJjyohTSapIcvC+pYryoqd83nGyJiQtOb5pGXdgtK7Y8rvmgB+69AyUOD4
ZsExrXNCXGi+Xx8cF8kjPCz2UYWeGw98XnPJInE3g5U0TG9hNpyaSs52VsHHgqCt
3riYc7Puith2rxq9fv4UBsuN82oa5D4/yCTRhG4ZS522qU9jBruGX46ym/19MRvN
LTTfT8VhMHKsZG5mJcLCzR+byA3w9pSAAundC6l5wSKAOoT1NZG+b1Y2yCqMOc/w
sMAb+nUrwwfnDHAQkW042EDe5qr8Jh7W4+ZWv1Bvpsf80Rf5NUy5aEc5sXrW8daa
wfobRppyk6uFpSOA+FIbmh1CaCr6vAXSrzWNhgZ+H4hjeaiFyUp1pilBBWrfBZKT
f1NgvuzJSxtWrLGW0PzlFID1NO3dff/t1BT1brpszvzsf7sL+dtTQf0/jJEyeEAb
5dHpUnaOh+o4d66NQQM5CWVo/rY/S26rDu8f0+aizMa04Wj1dQHwTmsVuqUrtmea
VdvwsCMeumd25RtAj2EnIAkv9VAUkjgimgC/9/dklfeG/z3vQ3lPQYs+SSgZN55a
1r94QXUJX4ssf090Pob17jCiPEhp8v4BTPEtkMkLA3U2lOEwYgzX4klmfe50N0Fs
i1WiRc+7DZcx3FiiO6HtJMP7tSedFb5Gh8i2AW3sVyJ0/TQOv6PcGTlmw1OEYczX
UnWDm0YtfWajeodkH0p1HxPjUkfVEtXcA5fpxFbMzKk6p3vQttC/vRwCXXL2Pl+X
R9/bQmI4Ra6EWbm7ZtTnFWjtvqpAoF974B6SBE3uHQL5y3oPa1EEeAfyKbCJa/5h
GvlxMVaf4C5easWPOQ3O+QoTtWkuImh0QVSmfBvnva5I6wksRdJdNeltJAhUcqXd
sAaS3Lmw30JyXBc7UiRBnVMZnWtYh5/7oOKq2G932rR31QX8Zk6QRCM+wroqa3kw
p4pXT7zkoarQ8oI4EmsdMIRK9QInuaq54RLacrnHzMljGKO3CceCvp2FgdTdS2Qp
/VN2aNlCuHlvCEfBteetxr1Kb2ESZFZXuZG0AeyXS8rL7G89TRpvGbeZz1/5AAfX
yCcqzGvOtjZyOWwrCupdch+bKMj2irWngRAmRCR2ucrMOPhxH74Bp9ECknSe3PJB
vioErSpoca3DTR9hueY6035CZU1c6Nb+9aGIrtlQ3D8EvbWljeNhhSgIHoJtQE/q
HNrFPtUiiFbuLNK9b3Syaqvem2Ih9H6L1a5lBqSpRRejtiUVM+zI7r556Zb19fmN
j5Ehy8ny5i/uYfsgevem6JmQubtqfWpwLlyVdvmxTVA3gBljqkTFhMGsw3YMvOXX
Aydl2Q2xumewRzPASBaj2jBgfjHSyPl4716RbRu9QQopRl1fKZIfSZn9hgdTaG3L
fPgeAYo1VKRZ51UgSua/8BF6wamqcLcG1Ga5++11b2srgf87ov/uh4ZQTJ9/d/NP
y5Pzo7TcEg/hJShH12n1/8PmJ6A6tj0T39+7PnK2bY6+Zh4aJNjYcyI07+rkD0Qm
KJDZLLHp0aJy6FOifFB5MpMP66XU+RFPpEKT0Y0IzTBu6miyUesMto6CQai033MQ
r8qZryNAXQ3Cx4+tyZLveAzMH74Ceem2Rqg0sLxgoAA3IzJBO93AkRtB70E+GLnb
TaV422B6Ir50iWGPQG8XnONWJHNdSKfpv5xlKij7eMoKAgpmKxgFZhLZyHsAVjBX
t4YxAE/N1ycJorLzJgjdz+keNQP9Pv2ypHgq1M5PqdT+yyL3CasHUwthzfiS905i
3UT5yQrgWfVZzIGBeICuSJPJMdOq8h0Px3SOGl9gxSYFHX8gac8DLmXfoSMETuua
kbT7FAKktk4wIxpFoUwtAK6TrPBkcSm1ghSv6f5KM5gta5e8fJA3vld599Ove74M
1rTizvVsbF0xwoAsZNMfMVg/Ycde0BVKRIxO2s8hcImzzEmfmPGWWdxOqAAjaOCS
tyH1GfHdId+2oVEoS9/2IHnRxkndGttfmna3exZfJzOQbxIgmy5r5UEvWnvpjKQe
VUQdLKCFOTW4y/8i4RR7HYdBELBZZgj20PkcCl+HRyKa5x76eXDZCdR/yA/P1B+N
XzrLJLMBx6duYWd7EKg3+khfRpqBdTy1DsM9tWI6wl5//VZA16VtojcD3JfUrZsc
fXj5p9SmUSOpWwUFfNPJFPgSCY9cTy/wQEXn6cSEBDA7sB7ZpqLTbZz55qfUh3T1
7zn23L1hXjVMlmowo5V59cdo1O+nM5r4GB70XfYOQcULUHG4QuTsas/y9Z7BjhB7
F8gF4wyPecVXbNz39lhySeor2A/FyxuV6uRx+aftO0BLDEmjBaDfLlf6bWn37IyH
0ITqbevJBDgNyLtYQ+ifOxoZgxiFTUiUSyhhFBh3O5GICzsSWfjsKbUjlpMqfMKp
XDimlhqCfZqd6W7BMlkfo5arP+5fOuDd6bUMMsQQSq470ERwOPkNpVuVsgFi/Xwh
uKdvc6RVXzhI0oWaaj84gWkny9hQmiCDEG7G7MeNE6ZA65vfjL9ssaYsVNsKasn2
M8ihBLemO2L8sStp+e/0xmwQBqTeWfXVUUHvGMSyQnMln8/JQBjkFKLGYYhfQlZ1
xoxOrM2D/1oG2yVrG68w/Hun92oD/Xcyql5hj/XBUFcOXgL8npFDD7ytykzu3zFM
dHBjV1nu7zzGHCSPuMFmDeYdkWQB10njUQlCkFcDc7M8of8AVkAZKXaeNO1IJcql
ETLWfrpYQa+R6sLc1IewJpyIWOIUptNnvzmiI/c/praeOXr1fNxQbfY2pqMEAha8
NuEKtxwXEoRj07KUBaAoc56OlqwSKn54jOmipMjshozjaZXuq2Y4K0gzHkAPjT81
4CGe7VJwukqAhWF1dJz4oDlJMvqL5x3nigq0dhShz42ylKBmh0i+ImWkgEYqIenJ
M4DAABCEOWb+FPOPVNgFtf7xFkNGMUkcg7kNgijdJ9zhk5cEIRRadHFoUSSsm7gL
J563erplyKq3wNVMWqoUU1j7W330tZ8kd5q5/36AS0JHl6JtitDT4TrzSJSY6rJx
6hWvzXvwGSoEY/G52yP9C6cOkf53Xi4d3zPqroSOrH/cYWT72p17vjg+/04lrDcD
uiKx+CSsDzBSFiDEICoTrQEtuEY6y9f3OnC0o932uvSjTm6t/tHLHjZ3ewv3vZYk
LUkwo4z5cTKVSHCff5YPyuDtDvUhhKiV6YEdz5WvLUbWiPS0Q/VJkKKGNqs4QnfR
L41DTfHDIGa+ICswlhibBqVw0XtTGOhzAp+05Bie9a3G08sT/XNrb6I/g4GuEGTN
3tQEx+YUAb09VCpKivRn/cXRVFJ9udAnnLRfreV4alQf71iB6lSIbGWKziAAJsxp
NhWogqr2rscsNR6NYqm4Ehqny5KPpyY0KiQ3VF0xFobK/eM247K5OrwCWQmaRYPo
Hqos5K/oZ1JoTrmIGeDIUS/zp5PdZ9Gd5X/XtGEsKZM000pS7sJ10Ulau/B+GxXp
3lIjif7BmJrCo1Ebh/o2OeujgLfFJjq1YYRl0Geh+vSfjt0e/4KJkiWWxHTpqQdc
I7kvjoKq3sW+Tz7cK74+OBP5dOyR4CV5B9K9VuOeC/d+/Z7jZ2tbLfaD40E+ebM4
/Q+qdGktp+0bV8VMCwWlmP3umAT1/dwoL8bf8ALoSALooPK64giPXxGW446NSoSF
VZaDF+xcU4H0iYUv8sw5Zol8gnLsQJ0oAb0fu0cUIYwufqagok/ab3VCgOMib56Q
9wCDkiAO7bvKCjhOEcaHHol5fZQ6gR77zu2iX06PSIiF4oJmU/K5qAXaMdjXNw8d
YtFvCFStqJIuc8D4l7xiRCDNxdojTLtJrwgIFgXtDPagi0nrOzCBer4A3PFZwLur
/UDv4g3/ZZaGEG4yybt4af4SaQAgAVLSDMVzv/c3PEPQEOMzr8TXqwJzABniUaVd
DjXJeX5ST0X+b1dibc1Wve9Ak1lESzr/XI7+FioVFsTav9itRLCacSV0iz5561SC
fc0Y6SIkVq9LjB68PVaYQXtIdoQmMB7BayEAKi31gJdKKuJlgEz3yQ9glk0vTq2a
N3qt0PcT8305PiC9xX6ix1jKEBmGJvd/jEYJAKywlhhGTu0UA1QpyAb6ZUPFNBc9
c8gfqcrsvAx5hct65OWDZ2cTOBCZHtev+y864ep9kKqEkQe6pQVlpYk77S/E5Q9i
4iv9b2FYGO9GN+7TSeou03H4Qb1d3iCr0OATNLruHyvkLcURuVRMMFQOAcDAcwR7
kblTQ5bA0C+lE3pV8KVtGUqtShWEgmDcLMpKil61Io1Ex3YCYuOOne74S7dS2uiM
CcR5dsfPi9Re1n/CuG9nJzoH81NXpjZi+tVhx253ZZaTIgfbHbEnCCfjU+h2ZcGE
d6toI9Nw3D/VPppLaUXT9P3jlzKoMc/4iaOrUFtnKFKZpyVAXVR0cFMASI/vlnl5
kp2L/4zaQGUl4SzPiqqtUqYLTP1TosJDRbEvRugCUQkVfl/aXbGkivdxd3OgC8mA
u8eue8O1PTGmPeaszEp4p/F5HP6IIeO5VTrSjyE5mZNVLssADtafP88a6MobVo8j
msIKp51idkklWgOXXaMDXByfOpf5imAsGJSBdEZs88FcUx6oXbOqN6N5H/Bp1ye2
YmDA+24c2gWUO89Ic7qg0TVBmhG044dZnYEsT5K8x30x5ZoT7uKoK2SE0WHf2a1R
Sx/+x9ACDtK8ZZT8DeoIB9X7FJAgZiRDDUlh3yAqyr7c/99JsE4nAVn7JGYOOAwC
V3haul78DEDJM8Tz2CcdZW9sZs+dalmr873BtKZVkCRDlXli2ZHD2qEQNZTSkAs6
tSLeYCqVZFvM/RG1ActpMb47Uw9+LjJXTVXrOyLodwB2DU/cwX3oPo5rL4XdcNUE
cxPWFOVOStUWqnwIYXPINHgl2S9vW9lKc/YTmQ04X7VnDl/FHPh3fkRND0xL9cvX
3ykZkAFNJJpPX0GXFU7SbEjyKpj3AIVIA6LqqMuriiEajKBA6J394w+Jz02iTJoR
AEGCjlr+AWfx5z09nIiq9gkr9gnXiRZ4SSnFKHXoPKd/WiiJJFvOfCYbyNsR7oT6
TS3bxNdhQrBSejROGBv4fAEgda6g4Zknh5nOC2owbxT6q5OoWvxVmsM1mhrYSnWA
c+uYMnIwa4WcQTVz4zJ7EKOkmp/QJJwaNWv5dyD1j07VLLRQVZ4VxbVei9dk1aOM
DeEsnhbhGcYmDx/+4sM51BMSK7QrItMqBdtLZInDa1fC5mkEEKCze8Sm43ZklYmk
fWVwPgFBczxrY/HiHBO1/vgtc+OZv6ZlJjRoK+WnGt6Xd6vzgybvivhZgxrR+Z7I
kEHdr8d4ygrO0vLBM0YmXfadZZRNoOUaNCbzZzIn5ZwG7K8op1DKdQyLWNbbU3fq
ncJy582njlaEyvs7yed9VI2l3guGd1vcNJXzOKSIIwYUb5yzitCOYmMeZFPajRje
EoX6Y2Dk79UsI84xX7n8Io9OnlUutN0fDDxW4CedUuRPxop7Ff3q3Rg9CwWBzTWS
H1RsX7AJMcCtVNDDm47b+zC6kcftvNrw1oQO02hifyI82+RG+Li52AqLEnBy161e
qpE30ajk/wTPj9ZcOiZPn3TXHRtgTNKHGdYQsSE0L1kmMXq4FPfxPB02vhmA4Sr5
LoGSawOeyUeFOr85PsQawAgSJBVknPa4/DCNhzXBqmhH3K/KFpyL7XgS3PHrjFFN
ja15GDW8n20XDUoD8LSBthSXZOQUyPh2ymwBIPSMD3dvm4yQoE0KETyYQ6Tg2kEL
BCTlrQBrvjGpV92H20AXYLLjHScoiOu2Ydmet6CTEyJmro19W9oCpmq8wQ6TihSE
LBf1H92Tc/NFL2JQb/DOK2jto/zTA81Byl8cBSHDTgnrwmtAxGQz5ZKMVoeciCDT
+aEGfahBBEDGTY2TF7W8uWOgq2nDrVK4b8jKJX+WMNbgPj5kWgiLit8oVUAcMb+z
RtcxzewvQemLVXy/ujoZOJoOVdPSHqmO8n5cznpQ/rMp4yGU0h8X7rEtl9qOIHZh
4tmSVwN0ex+aou/9IKSZK2++kGjn03Vfcy4DdHuyebbWcEjGvyw7Qe7QGyveedlp
CeVxmKOg9HV1hgKRBUzKSAv0iEWBvfrXUsDiSzkggFHp4iDpzXtw2ITws9ov1S6L
+SXkMZ20aXefTa3CJ0UAUpOtEQqjJLASWLXpRWQ+lfVoWQFLGRw0+6fsxxAeKatb
b18d5ZNlk5ldvmjW6C3s17DyxNKgw8ZITuSMPd4Ueo1nDM1CXh3mXO7EpqqS4G6H
GsJFBgz1RPuBiZsm5JWZLVJoHNrey/osYCbW+lOUn8TmTuW6zfUuhKXiTzDRZIQ3
ApPi2IyR2d4n26cKiAom6h15Bp4UHc6zv3TFrakL/GEDESQWOPqF4Tr366VsJz1e
xcJAkaVXFLdAmkFdq0YGJuUm0mOlhV07SCrPbc1xGVCeqwY6h/AnnahDOsxL5cGt
wsaRATZDiMltKIDoJaMpGIxy6iQxzrGU9yvAw97AoWDgW6erwMvHTmBJY9LubUmR
rNxiBM2PNWImEL9alc69bJaE46jSW3dgrdpYZ+TSPOFLP+TSdNgLNx4B5rkhIlia
RBkTwK7QXN/P4h8nUqXIOBvUPLJ1p6X3Gfkfke2Tuom60MgPri7kPWDtJBVlsJhM
xS7SgF0prG4KaY1u3tJLEDM/CPWUnk8ofs6HK26H7q2An6JgTKPI/O6rrCl0MYcI
gQX+RVxywiy+Sr2lJ0uutiOLr5Jc0jER8KuTxNgq0brtzbo0AviWFWesSIKvT7eG
NlkNZHYNowjfh5FjnAMxHijhpHnFbpwKjgXITCLN00/GKbe9DWMXdLgweGYaBJbV
mcmkgPG9S9402j108Tguk/PwaZOBfz3ibyRA2cQS0bkrujbzAuC8idJDR+unNEDe
KL1JJiVQisIidEhGTPDJLJHvY3mESPtCHyoaTuYGOm4bNUdeOYCDq+M6bxogHVqU
ptVGc83Bzlodxwp8DEjm3K6jAq66b7ES717wk3S0AqGfy6lvkVXxTAatkkCbDJyX
AexhholT904rgsjF0uB+FmuL7loXKDhoRI387hBmRgS5YbSR3pawkDd59jFt8BiT
A4DiqvkRmlhXWeyWj34l0WYSgA4KELijVnwUZpkBQyy7C9fgPcXkBUiSdN7YRdNT
ap27app9FpNgepY8hKDpd/NCCYP8eIFbWmPBW+9fHTxWn43oRhNlj9cvVIuUWDKK
vpQ79BYcDzysUzwN9cvFZ156BEOnCoT07EtObP1TOb/BNuIXpv+4upZ6zagnc1AC
LMbm70JTasFJZFRDWljsw5Y/UdlcHqf/pq3jKiahlzl5RvcAw49hE4oE/HXgiVJy
Mtx2BnN1SKgXMv7riPHJREv5zaVKZUO5YCCThgvpXDOWSWuPcIOOAcUKpSIryV4K
jWMdDUDiDfnn5qZTVbFsBvaUPN/wvesJU2oWHlmvn/4Vfdft/uR+UZKViQwm6NG9
s0E5e5OozdXhLdg3v2vVMmOz+Z5sHB9j+1RwiZMgPseSevSU8bCVXscNbmSZ5Zu0
AiQg31bxrGphMrrzWwrUHxW/X2uiq2jB8xE8zbAbnFc7ZOTUhrXT1fA6j2wKBSdH
lFuKaNVEZsBtxUoEpoOcnuvSiEbYdBxt9csaKOdaSL9bhUJso71iTN9DiRfmU6LV
OkMJ15fFAEsyQWwfaV33zUF0UJgJwBToAG2hZBKSpa7zoBzyNTAdYUpK87uvhjGT
Bayp2b2QlYTYlWcMrUGfwYkNgPXCMknyOA+/23Pwc4SwF9MG+kSLOFwntMZAUxfr
A9+pb14NovyeN3hoqc5qgo9EmWS14fimK+BgpgfaJue8C9c5ZsP6WgVj3gwHCaBg
IanIO0bfT3BnvBZUC8RKE8VH5pJ0rY+wP4VUayxA2lt8AIGQTNm8Gg2A0BhCSGGC
lTW3ZueUqXbsVxUykEtgDTJ/EGBcEJyG0OKdnGp9Cq1Z6+VwUsHPLnAP/Fs0dEre
+ztgszr2vnRsn3rjfSf6/Ec5RrJNwmRGzTl6uBouhcOekLiS4SZQgpnMsdobFuYR
6SbR4qaPCdddtbp8SQK9Pm8fHNCMiVlIOoBVTsUu0BNkRhuLHAdqIh6m+X9foLXG
4CGwIMqZU/NfV3vxp9SgkPjx1G1yfKEOffTgNQrRKMt5D92eJACwYrnQ4W9+eIlM
ACUO5bcSD0LztA1uwl7LlKe5oOFNEizFltnNmFJoKFRjLZaUV4CRuSnXP2m8sH9G
5vZTgYtYFlqCxd4DiSKkyQA6Q3c11Bzq6paTB0jscJj1pJJGdcaUtr/blXfdJcCE
BvEJ6FzvN6HRXj9SOu+DUtvDmNHNe0k+lP0AJ4dKVOqpECUMfIlFBzwfLZdpFhmu
bMxjtZ08ZTQQvJzlRHnYOPBbcHOshjvItO4iHj3iT367kRYSNAPzstuBS/lf3W68
NRnjcPJS1lRTavAaRka3DrCxjwcbkRei+7gHKus82c5Y0g50/xGDrtW/BVq4HNHb
ifQkgtG3IWT6OobqqpKg9ktDSDKkrze6UNUJ4kNFBcZUQ3uWCxwmNp69lL7yndwe
n8YLZSQebrVg9pF0gixw4Z+/WIykYYFyFpfiJpT5XrD7BNC5kvf9S9yClIR0JYna
oQTG61ifcenvC6+RwsatV4OaNQeRSLWAE17y9fjuivuzRvGHI87RxZTbe9Mfo8dp
NcOo+tXDdfGGSxUnAZhdPoeatSA631fZz4hUMXA/0+3X/zCu+DgXUDa5Xe8S7CCI
c8OeKTe+mHX9XjM6uKK9lbsMdF1uYffhLxERVrTF2u+HAhELBPGUhUmUupYeeZlm
Q9kR0XZowZU9bk4vlyX8simvkEQ5enxIVUPnIBfkOfgTNDMzhSKdgmYWHS8PlsK9
Giu7wxrRWSLnQzR4kjeEVsA2ZESXkygNXzWUsLwpxWIV4bemo8FZK53DrRbMpd2j
tuoB5aGZ+ksh47jVlxNNrbIFkX6F2nki2end+DwFL0PhxpZp9DBtodFLDxT5Nr0Q
kcYc6n1KlpRen/hZMnP8unPXPcwOgvDoQXes7rpDU/merbzT6Ao/xZdUocbhLwsT
XotB/9s+3+zrZv6/MIXV2lOtviJbrxd3eS9Egn5fPFnYmI/EPumW/VBJZhW+18Wa
iLlLRFQayLtV0qRLZefkq9/DZJqYy1GINmYWEXK3r+DPC8uuJOaS3tDmcvnZPqPo
Hh6RYxKdrsGrnEEWKzFFHStTb/ou6AyBY/rOdG2Psd+9Ou3MyLICBKMg0Zloul6O
dH8XstwXw6YwjKU3InNfrTfV2f+zL18GPytJtE12gSL2A7a/TIcsp4B9/I3lhJXL
YceYSRrYmwbqZrqD7aAQnZ7tovNS6Dowyw1HaEDN/KaypCL4VgpEi/lZ0HP8UVao
KpWnH8xu21AIP9y1bdvAX3cbpNAnNceZpA1ZWQr8qUwT5u6h40vuI3jBBXKSiAIz
54TfHQAYgrQ3Maoh7lQmZIMnYIjBMNT1wHecYzuSrxmTqMxgEB1NIdvw5/T2Vy6F
xBDBnMBwf6BBiA9KTPr97OKhg/ojVHC7fRW43idnQ1N57yin/QAh9qP5SJIKXXoV
qPxR9CwhIFzfKeavOMS8lcrDmMgfpVKXZYck3nVb6Z/5CB488I03/AR8JUCbuCOG
/N+kaI4KWQkbJ9mUgVg5A2rFec6m4DWH06be4t04c3z2rmZV1zDBYp3ozQhLWhFH
arf/DmPu4qVKzolujMiLf8WBkN+00SsVz+9SHRriqYAZFPUJKIvegJTO07fYnq/r
A/P78fJOwFv4GE3uAm2TY3ln942BNVXK9qzJ8+m8vj+oWT+y3v+Z57nHrf6EtqUF
p814MzrrzXAFpcN3f8MOyeRqiYbrAEAXxbMZliTa9FCpZhbBOIxessZ5pZf/ebgB
B4EOtVhSvHtTnAg/oPEnJrAho1ASBSuMjAq4F41U6NuhNRHUw4iehsmeQEY9b5md
kBMD6h1cJ3FapQ4MK3RL5LY17tKKc691A/Vn3Rw2RvzecUF2f4Fg03F1Bnj8DHnV
Nxna6BlL99HBXTuq3ygmdIAbPX+KvR2tK01q3j9YUnDuH9vZi62+wrW+GMYSGOF7
+4X7kJSNIcHxSpGbKpMQskn1rtnNrGUd4CKDBwU1BG3nEJ3zC9td5QmL0deEQW2f
BpAc/E1XAHFLIRydjrR83hg9xo2/JDUi00Bshmm6O0jpRiHIdBI23/MMzTM2+55M
S/Ydx5Ht/bn6APUr6g938TeD5fIX+bPrdi2fwBCHwLAZKj//m+JES6/NyCTndXwx
JIlp+5befwbh/yJuqWZI6qEnsw/fblpaRFP1SRwYzYJtE+2Sz48l4iSns6rT2aor
VJlbpIXDwc6F50TNNkjb/Wtb2Uq9Y4OFAUqPNeWsHev+B4pgufjGa1rhUirmMENw
nBQDyHI8a0tMkmAailOwvk92qtecoTTpXURO8cHllaZuHsr6VlXxms26gZEgRNRm
l+EeJ+Gl+GKa5AAwZYuYiet+MmzAF43KnFbivBynN719QhXAbzklMi37Y8MvFtQK
ctev5Yt2Bibw8fwnhZyBqg5syaSEMjeqM/jNDI84qYiMP4Pc62yS/D0ZdrZaP/5J
v9Qk6LPmIbVKaIFdp8gUAWyEPap6xUYqtRh0Pkrn26qsIEH4OEO1pB1bhFLWGMFS
QkI3lOTVafyqtRYGLePiG5jMp+Fq/to//hSouZ37ZVaVmJW+0ODG/dOpV00jmDXX
VaPI7AS2NeKZeNWDvBRDGg8+X057rS6nMXnhzMhMbueyU93QPtgcj0wj1IK0bkR6
56Ld1PE0cP+9aQ+gdFYHVVhLUrlytr9ZUobPHqH8jwQRejdX2eyrOAyRJHsSMUm/
7nXGSDPuCDz6uAQnwz4lBFNpywjDTjpE6RTgK/jJmaxfGNRncMANHYZ0IbDi1F5c
ESnziBVDYgOVYVuSaFVCSFt6uQRLVUwcajtDkxZbvNW8gkuZXJ8M1EIa1Vr80xMV
QXpTxk0SDhb/bWcEJNOaPiwK1Rzx1m6p5tH7b5Eg06Pl2rh6yl2MoCzi6naGl1ii
ZDQ+QBkgIp3NLAyup+lTibC1xANItoRNduc5CFmqPo+mrBN1y0RBPePwQd5MaD2S
BVyM/Z3qx6CuSN4JKfIfPxSo1lHQXp8eD1QnFQpaXY979rJv7ORzc/390kmTW7jC
GR+A7SSoW5rl54q1aOXVUc04E21/WXghe4Hddhu8NU7PAj0e3bG6SGr0nuBSaCSz
1e6/97idyqHTmUTxlyFcq2+C/hrzv5vyKibu/5oEM2MjxGEHOsl+EzMD9bGILT46
gJhDS5az5JbeOmVM8Kveje4gc4t7kHErE+8XO5H+3JNWKxfzO5xl++xzrLHcT0xv
spIVFqJ2Op1Sr0l5hwhJGoL6cUyTgI3qoLOyNo5mDUVswzzni2zdmJts0iswmu3Q
sOuMvNaCBgijevOScxJttieK4ORnakiHrstiG/VsLAOfbL1gDvzM+bEDdLEGCT8V
ZbstOfkLtrr/Fc+Ql/lYB07EF4s5hV1CfmNYxhE7r3VimIUohC177rib0edkkR1y
C2RKnd2Pk2ISa2IuemyWJBxcbi/Z4rb6fi0AHbk4wCd2GRBr76vQjdQzZpZ3bYni
ECcpuiygI9VlrhUc1YSQnZxqsQ0A4vtpB7lgsKLJX31Ghhx+61OmQTA2Z9/gyJku
XYA04968KrqSwykRW7AH1+cbSBp38vM5/Bo/IMDV1sPnFYX+j8+0gUOww/pZSXOA
FcZKHNumhz6kTS11Nl9oCGryLzccPyyMQGB442WRJoU+QUJklyNj1u5fS8awR+pf
AZGfQCf5Li97jBa1rT0XLvIHJEEJ4PWEujRfqKEp3DIOTcKwheZ9b6zqhOhz0+zg
TyZBrxg6Pyha6b8hWK+jUTmvTam732+8VJGb7F+5L6JsrCCCclPLMFI46YmuKyGo
ND3sP7c/lbVQ/9YvJ1ErqVX0mvOZOErcVfzhPMLpp6IzM1AntQ4PvtS2uJbaXP10
dGdiO2xaQ5St6W9gaDctFKgY5dFYCedfB7HsVVhXycPhVRmFJ0FOj5yXY/jy/1Ya
mF0CzHovWB80Lc5x7MZiRSG/oxFApQXAEDwVOv3u4EidVMSnwT0T6efCPravqyt4
DZQnLoDN3BHFtVSJ4/IqA/t8+PVCScVDf48AkIjTJvm7RBScDhCkvTrwaQ9gsdeR
n60U6C+YkdaKBF+sQuX6OEwYjNWc7RYJeReLMo9HFuCQRgSq5TUbejslwphUYjy4
X0lX2/MXyORg8ywBFHTo1rSVAslPSx+3lrNLXzfBLoYVeO5WCzYxaW3BmlDh/Ms/
IPP92K5uUI6HrWRc7bvzfyRqPvM5aqrx82ddC7+/Z/Pojlsc49C972mGAxiQORrZ
3Q+qDr849j+5D2uQb2w/YQR1O6kAq3wUdTSApPvKJ7lqs9WZkwBW7oLZAV83RLov
OPCezidNHejAUOOUvUupXiZwXOXAH06JBx+yeesQAAbJPJsZijF7RwgwgvhlTeO6
5WUUk/vzEuof8XUTtc5alXI/As60QB30f54A2gihrK1GYn+25QidGYZVFshMzXic
ylPeepomEcTMXCLw1Vu4jbxjL638wuNNBFejWQmtnhkPS8+qHbPTxZG7fihKdkYV
b7C6Eov2gYzCM/+IlgQypECa/tCg04uM3p/0YwBmn8WMwKmrDJI/tU5WkIWzZ+3N
lEKgf/IrsLbjDButLfeHy07ux58FhUMXV4RhZrXoQ/MJcTCNi0Yd0wKBC8+ffbn0
Ev4YUhizdP/w4yJLMIHWLqcSUhGddwnNWTQOOyJpZsXFjvY9oDn+rJJU14dOpnuF
kypIuVd3Sts6WUdfzIi7H2L/1nYmkQvWGKQA5W05DAfvhWWWZV8cnyBu2j9f3G+H
7d3bv9WJtwKryqkgKdQqKtaatCW3xd0k5wWd0m/9vovx5RIVEMnWiSkk2SlQ6xLb
5IlagkBNWTX9d8tT3WE554tUIcjww1rLyJD1wHXb6GBwlD6PTpPwLMNRN5abaUw0
ArVGPPBX7DRc80fEkjxQg9aKzY1raZ8eUnPceWSs75RSTjXuJGEMST2hos2YVfAb
ZuAKZ3CEusIN7G3Xe6Ls2hUQMQ+1zsViE91w6yq2pwKvyw7M7sPlG5oOFAKfUA29
PBYbfs6TEbay+DC2Ad7yB7u39hL2nxgG9I5pkGib+bYguPr9qbi7uaUzjFZBFekB
qJmR95IiYnDiCdMOm+jN5o0jLLBSIwTlknnZ2M9t1NSbJ+Ov2+wUwnbPkmU2TZzf
Gb253zfQxD84A2oc8PgzGYCUEBpuMJExzCXkfRXrsJBdVWUACKxbcR1HYMsPQ5F7
swsEubpY3KEmJndiW9FXxHXb7BP1NG4Qy0Fx3lOuLekRPe7NjqNrTNp/9dBV1sfQ
OLNANC3o0aDedkJEBt143IwIc9Csi0WqRuXK1daQWURIo/htgHbrF0ltykygaEXG
OTZE8BkcTBw4CVeGTBksoDGauCeXnF0YC3sfxFfuSuNKAfmucsYoKC516ET5+nam
3rjgnNF7hBCVo5k+uakcLDsRIbfUICM6oT4aOO3J8X/10qgpcaZX5gcieaIruB6i
AxEWRDlp+bEodGdktsO0sgPiPNHptH+vw5a3jla8pdOThxe5yvp34bWpEOqKMr99
1dCjU6y+rWCPAeEp8Fh7vYRCBtg75J7cfTUa1YrQPEUhp0nCB7aUJlh7dEuZnv/q
6sOn7lTMpg8uv8sQlRhZc3lKJXR/NZmR5ULgbz10FYax2XZRxf3eI/ajbS/taYci
PfGM/azMASdCEoXDBDRU9dZqT2B2Px3jVzI82cRRMInwQx7IpYtLJ8mdfFKnwI7x
VSFZUVaSfoW9pOVBNX6olCpJ0fmy54MnfqEItQfK+ACKPJtf81lYrnaCv8Ke0FF7
1TWa62yXwEXaLJzlFPg1SQ1AoEQDQhHL1k1PwqFONvyMHOzlwA7urqykpJUz/ZBl
eI9KafLoKUqeBajkD43zS65RlzCmOHuwEapq16HToPjaOF5sBYKLIkOrbWZecjXP
bqb1CJT8Rn7VAg9FKBhXl33drvvdi9FrU3gBjMfn4KHwx7FAdsv0pTnKgtOUvItY
TfLVdwlkqdgfT82swsDruion8blRqgl+t6583CBO2QIanvNpsSR77Ow1XoHljajd
snu34qg9K5DR5yLtKEcU/Zseq8gb3PO9CeOTAR9Ey6p2fLxATFEZMpEHsEz+Wmwl
Xlsl1zNbWoR6YorYALnGoqQGm/aBO/0rkcOfsyzFDmvEcQAlRhAT9Be32dz788WK
uQqLhQhi8kVImQuI3oh2NKB4o5ybii0CwLQEM567dTO/3sqrOE/CZXNQogr0fpbn
smkhlzhHqsT9bdeyMw4uyfnQO7JeOq/sNPAaBbNJ2mcxPN3dh9wjawZ00VXU+mAd
+08Ssu4qmmM5NadZdwrUHVca2KIo0Hg5akdS6Txp3BFZQD8ITKmrHbanyQ61OgdZ
/3R2L//vMdi2baVn545wL0BXhs5UsZshiYNaVTPHpXeX25BloIhAPWjknWZNUh/W
HswqxcHKkG9qPTCvyFEiI137Rqj4XEGBZOB2wfkaorlyLE60q4BJ7v8vAoJINgpr
JvmB5RrEJmpnfptht+lJRPRpAWFXiXp6X4y9dox6DJ6ec/dMkG3sYiIU2f/g7jcB
Qe4q0Jh7T8aDmHzB68PU9ZnnXDMFqXh46GomQZXEbrJun4on4z3zI84WW8m4WO8m
TaITdkeMIBoyheRWk/jzvptnia4ZQ937aTh6nK+nfEuEY7uK0VhqHtM/QtCeL3BC
IbSs2FncS489f069fUq5UGWjMZpDZ2Sq3cKMQmTDXMjG/VOLPTeRcoKsxMMIeBL8
rKB+xB4PcOMx7wYwhcnX3YPZ0mj1p/0sBnGp/sY7wf+nXaRdobw9Ay6VRfIhigcF
Tr1pKmnFOs9e0BosUgJoR/OXZxe96E0NaFBPXNj33z6VQkJEJA2Kl0vNAHQlupHF
h1g/XZMIM+UkVHzu5OqLRhMLodQF3q/mphrlqvvuhQ46ghsnp0ZNBayqi6y7PwFy
ah0s0kxdQ1CARV7F4koqPKQXyYyJhoIW/UI+Dmpry1JLKz1hORLWXjv/T8wloeKU
Utn2cI/DjVrpTcQ46Xy7LPi61G34jrvRAVbk26WJNYwUGKZY5pMvRbhOe4WxxPNQ
nzcnaBX3jXLQevWPJCJpGFiUjrUS/OP4l/YPzcoO+2FX3kD0TtzpJyMAB9RJG56C
y+KvuZnySw4KvJEg968TIfsQAm2+b99vr6Mv0ulMWx4zz/CeotawnLVbcJWfm7P1
aEDD7x1DNHQhcFRad8G45Sk5TfhTvqowM0tMuYAKnhDORkFtptyrMqbhsSp2fxMo
7oAYem/I9bO4jv4/gJTCusIGb3wLQc5VV5kpn6TKFz+WClKF4OQrpuW30GK3gxIt
Adew2f8pvjxjyncnF/dEbqQuWYueRyaWS+7Go6k6dPyuosGCufOKhIuaPfIEbi1W
nw/v3ZKnRTr7Mxwkx7ABCbYw4DuJxg2houJeRS8ecN7GCAsixpx0HHP5mNH1u/80
5Lryp1Bjxyo5CCO8VYrEYxz8KaxW97Z2su4wJZ4d40SFo9LYe2iU3mHmTMvobDYz
kwdpPS8iPOE2SChHI/KD2bfI3TVSnHqDhwRdsyc/GTyuYZyI38HmrUzymvPdiVQi
zdAXofQ6jUSu/l2as/g+V6PPjD6+JSQTAaoVVPqcOLySV5kPwXv/sxY6UdnO9HbN
4qRiEpKJSD/2itZ8dVV+LYHA5hYlz/qpp0qwQa0mNFYDtxxTTARQFLgpuITTBiiB
Qa7exaGM67dTT0ock0XUh219Plztkv/Vm0a+dUelZau0GvtZ7/LfjeieYVkTIpQd
/+zjlee0Ac4/ZfXbH2Yez34g7bOb4sCo5eeB5mbRQi1Ogs0WwK6TGVj6RpoJfH53
bJhG0sdxnJk8B4fUFuFtk3O4h+CJ7dpVKmm631lW7YppP7oGgnTtJpn0hcd5l3h7
/9LkfO26arliLGQK6TDZojA5OMJY5rVZfx8GjIw/uwRZ1QD3JlEqr0KzNwI5AzBy
QWOJNixjClaeIbqBBdhTrGoANcmUunbK3VUwDExPZOB2DobEmB3ra5L04tp/s0kv
M8KSJkwUDNm8AE9ynWGG/K/MqR4Fi4P3urMKcjR5+lcLkwQVQseERJRRNVD2VqFQ
nvyv2XxwHMASsndVnAM85gCheaR3UIAx8HlgbuVPhCJFi5wqRqtY4M08vubNc9pO
NB9osFfqMt+aZqUbfsSCD+73qB/8zojRrmYJ46PlT1xK8+BEPqfQCfsEE/U45qML
POPbFXPyseanyCcj3Auvj78HFWI59qKQ1OChAYfDmjZsjTI5pflo93XkyXewAPnH
mmpDDdeQie9JBfQuz0wMg651EsdhPuZGnqSGQPKvRsdF/QbTKscgBdZ52U94gP8L
S1IrQstVeIA+7cSMp10fIdaoMdReSVhZ0OTO4gWsc0QJESZ4vP0RKteQhAhm8JDx
uio//aXVXWzI+TOvwkKhehHEMMWCtk/jfmVMOtsG977SFBPEuZ/NcWsjS0gThAp3
EbPSe0vkscDjg92cne1IAWMaEMYer4fzLey0u6U/W5ZyylFzw2pky7m/gMk3P8ZU
C7+FBOwLzzGcJ3qL1LQyuXuvIem7z0lFep/c/YG9luM/y4EbZURoeOYxhrz/hUvP
/VDoxdH/CmkACl38wxlIVWVICp8tADIFIcLOL/il+9cMEwCiaKjsI8kq0w9Kb9Ck
tEeNI6K2CrsuFFJdjAD1j/ax/et918MxKPLBbvsyxLQBiZq29pOauMNDw5hUEu+M
q8rsExuAdBoiid3XJjaSqqsZzMldXd+pURrlN14TcrougNo7yqhx9PTMOxvzCu/p
OZHjQA5gb5qhIn3cVpd0DmzPQDthg9kP0RN1Yx/Q2q4FBLFqOxirgR5jKZI2ED2Z
xQeK6SABN3BloqkhyQAKLKt/Tm5px11fs3DQEHCVOeKkuXI9NwIc4M5nDUWfnixR
GOcZThuRUK2eA01hgt52Zed1x4nD5oKW7mhZAbbv4ye2p7ys0kyjML4fj7YG5kHO
nqYZjK98+b8oLWfsuePm9/LeaKXpqqVUfB3C4f1J/HOpX30StmGAgzUVGgQVnHKc
4n2krC9ppLQJK+MjOmK6R3q6/qcDGUs798cE70Tf42fCdvDqhUeeJPPaJss+zVg0
ahapoBgXWnYa2JEqvDbIVxmION6qdWF8vnZDio30CMot+o4SPGXeFOKa9KGJQkRa
KppNjwed/ppDVVMv5s1XXPeYW9022KPkvDm6n36I+IW/CASjJZ5NwdMAf0AXcCGn
jSz+M+Pl1Seo+SWlYNh3K0jY+e/bThi1djYZ7ngA9SkyOoZGEqk8GCo+EGAL6q1k
Fi1UPzQGaoQtbugmoQzRg8pfSxgSmXF03bdB0lDjTVDl+T88Sa0YuCmMD3Mu+E5P
pOJC3DtztOiG0xELVDVHD366avFTLcnXGFy/ozwfNJdNloyUC+8F5JxxbrZohwzy
sHmhICl44diJenougTNRmLBL5b0kRhLlPsJAYMe0++U+u5emRRuSOrt+rWigYDho
RDt3oPBttCEfm+m2q7FwjZRsx+0Az1RbdNNxTq3UUdjS85xgq0DyByE1kLn8QvL5
Wc/9NgaG7tUwjeSJoCFbFGucWumqm1B65lXXeHnx3PT5JmZcLoKtwMe5W6enaSPp
z15NxmfcJponHJwMH430rc8asEtyvODbr8lW8Dk4iIr+UMR+WlLFKiv/0M55Ab43
bDpor01g5qELFBJ5V+xvQIVhOQ/Zfd90gmpvN/9w8U4U0A5z66GDLQ151E2B6U6A
+vH87xvQzp4JXqQux2ik9N0w6THdsfBd6BRNrVEdQp99RNLyxjOkI6i/cJJ4u4FV
KykCN3tZ+NVfGysuUDer6kHJFYI6MW3PujgRSHTQI5HJT31BpUwprOrs6kSFQFJV
QkAaxGUA0AthXlVWhgvOAOl79wHByZRzU3k5wSF+9C+nQT6mIqoO7o8oAl3ibJl2
6MmksDjcpizYwE5czUKb2KOnY9KfLCNsMQNPJYxuUxD19AQitB0ih86ShnH75Qyx
XdjplTQKXhRsSt4E2DywxK8otPH0AX17h1UBbyZtXIJp8uApAeMZ3DH9ktcDANkz
/4LJt7KAoALodVWzL8CFAfN3d55UYcOcy4KJWzmoGvWeOuZiycRFX40nnWeMkaVK
7XdtuqqwAOrmdySW7lDlJjgksuyCuVBf61v2KUbsRz/t+XDYv6CQ5Nt6sZqZVcu0
uziMywxT1psggh4GOwhOgUHUaNhEWOwhp4jkOVyULGRQoe+yfjFKm5UjxrZxWgVq
YbuqBnGeb9bcfFmcKACSte1pwapf5KbJzhXpYkrqy/ovtoBA/ofLToS8vsa5g6w9
99c5V9FOaMOrlkaZ5BmQajrgR+5R1B9M1RSX9dFFdl0X3Vn4V8LLXQ0kbmsOjxYm
Ffubycqjh+dgCn2nCBmLAERRtfvKcjB8MEi0VZVJYrgp5Pp8KZKpN77luBg+DARm
DIJgVkWZdYO8Yg85zuedjrFgwC1vR8ZggVrDGi70ro0lOxUxglgTQjWicS1pDlrv
0MnLSU3vPHYxPWF5TN8sorbhbgVLo8kgu2tea8Q88wim2QwSVZWzXPT8newk8thH
BA+4kD9KYCyM3hUt+n6h5qcSKYjKr1Cb2nQjXFqf0yV3i8LOV2AE0PjEW4CDJ5SQ
h0mTkGcPc0HBdIm8orGY8ei2IKFxRGmV6umcAN60YOeBSU2mtZYnCJ2ob2+Amivb
9Yido3b2DFVIK/+NsbdBGt7P1qd7VJmeIUeTFzXbXHba3GJLn0gcyNio16erdgyi
l1Muu81BfJ4k3/yhi/MCexvZbY7hEstn2iBlOlKhTt1yPEv2VqMgv+Yt69b1UwuM
qpCJcLs/0+sLqcJolGzu44VQKWhbvAg95Dix2i7wuWUhXxf1egEnGuRWuvdVVZTp
E90A3ntyJFLM73EpW596e1Egc8Ey5UzMMOTUpboCtHqyAKCVgRNw42Kqw365oDAZ
cA/8dZjLIePkOSsm1zLKtCVLH4YPQcQoIR9QPrpV5uGUXUBNG5uycC+hOuA4owZC
2zzYPtmoYFa9A7KvAY8spqbjMOdOp01yJ8vKGuQ854g4prGRDDkfJ9cTgFN1sqB0
R1gw7ft9yWSmhQ1r+BoLD81fSV82TeGBU1qTmMRWejr5IKPCxMPBVdVu7Isn+DMv
57jmTIhOyDPYeNml3IokUMZtNw4L7S/QRKGlMBsibBRPmVMu7mtH8c0TXcilW7jr
sUZWgbD2C4g5Y2sOerG9dDRzkNqj8sBsdF212u/CwOnKEecA4gCbUraxBHoX4Tnz
ztaVzmsvtOOZ/oDU50RW5is5fwtqjwQnSYG1nGRZxxPd3OEqXbbNiMhS8ff+ij05
BvX9fWFHpBsfj6sccD6pvCv4npsHGv8Kdc/coK88tABfI611QM3dmWgGyW1sFNDX
9qogLU775AJvG3BIo9BmbnFhXTzVuAsqjs3q6otf+WlFlV2JZOz5SAyzotHBSGQl
b/3BPR9iZTqcCayo/sJaWj5Saldc4ZyWwxrB0p80VC6BCunDqWYWwIwJM4sb2x2P
iTci+M93FxmeVhk0VMD073KHyPJZ4xtvigMP4ekhW6LlSrJEbXGt8mte/8NK9bUZ
cmk+ZUyAsJa8s6w4Zy9MQ5HaEmL4niQFfkT9x3ZPoxq1lzytP7+rDeMOrwrUoZ8D
dxrLwKRW0iqsgdYlTYdLWw0jxvgIjAPURwK10XPDqv/MIoND29t8UXezefZsif3r
xeomAGjLK0/jNa+DDNzMfMDGzdCfz5wtvbnKsH19+uhU/25C7w0DSiUrgUkdrvJ9
VzFUBwjulkP1fZ687OcHw4bmA6SzGZ1YS8IbxOgKr3OCPMzEAh+dV/pERlXu39Xl
vSiqBEjaXZe3S0rZ2dtzp/cOCNZdfo829YYeBV7wcavFd0MqmlqtzYrT3H10dfbu
uJY5OQDcgmENyou0sZ2OREUkRqMJCfDEfZJwEKa4Mjb1j6XA8tTdBJJ4FTAx9rlO
RWm7VgpeCBIouoICLWrGoPYNv/zYgFyG0N4lgPsqIaS4a1BQ8A7AUKNz/BXugn0b
PaEwy2WAkDC8xlhePPuyRm+IC1BpMZAJB+/aPcZVVuiyADq4740okCRD81BRPQJH
UELnc/ppOhZHbO9Sh92TebuXDc5MrrPPRdhMJafCER+A2ELCI+xsXhgMhxjfS2V6
rgzObHQ+prXQt3WlTQaFR/HBJhlG0uUD4aJ855YGssw7sLAApy8LL1G0YVQyQCPK
MgHHYLzZlfQDSf4n07k12R0oV2yqVfPJKd2VY4DqSe8QMZDuIr+dJGauJN7JNdt/
qEJsdE14kZ2pAJeHGl17+ui3e46CYWP8vU/XJ+xu+DvgV7QKe5RpVAOIyve1Fgxe
WQXr9DpfOwqBRXCfmH6Bm8Y1VLW2+N4bK1XMWahBP8/nG4xHW2UHW/Agp/xUP/2F
5o5EPsUZeVtlrOf9a9R6dR6GADoG/MJGYk/5zdX7q+TijiJUnz7FxP974ahj+Yku
WC/WWvxw50OXKQ4EAGjNMKWkodMo0ItZwi5BJ3U1dPpa8+vTdZ88roWa/cSZ88o3
CxZePC2aWSn/7w9ynU7L9NruPaGd+mbccs95Xj20ll7G/OW79H/UTJpNjbamN7BZ
0EvzuavNFaGt6ZDud5DBd25nTzd24GjAJnF/LCLBGXSDEF07KExfzQ2LyeA335V5
hjUdKPJ2lonLRJ51cnWWXxSNQz4zMSAXFH0pIbnaS+G/J9QjoU5J6MaHc+G3G1lf
8tXHvzBWPCramGJdv4qPFtYlwlIai8P8WmF/LZ6C9KRWRPlMRxW0QWZoL5FkFk1M
XVzmvvyQQ/dJhwsQ8UQwM3T0akXH9llr6Z4ItLJpYUz6+4uwiYUaoeJANizpgNK7
T3EzNoGVkcSbD50Uo6fAIG7lTUTNKRYnGPrBip/jU3jsXY1oUm9xO0H482SAj/yr
NidOdw1k+QKSPlQpYYyv4bOOUCpECH6f8eieLIOZ70dJfuzecsP6qMZMPtFeMnQL
4VVXW5h2Dm8/X5j1y1suus2mIJmbw0nXpgxsS1NvepEycWA2daUF3AgGcMGsf231
tvjv8LOOd3YLbTOAzS0qOpEKglEx725TE5l0GID32I6fpfYj89N+wXYP4IXAo/o3
ZG2Ha81P4fJ6pTVS7DrGYEtIfbdU2P4/lFz40NVpcLxY064ThpZ0clFEdIaAmJU4
EigJ/V1gYE2ALlvpYnXsHVTyaMScK0ShzO6hTUntWtmY18LxJ7sJ+89cJMo0Ulmb
Tye+1sdDfLrJUhAlgLFXrrZuN1WB45IDz+rgSi4fdsGIjRun3ajNzkmViIbEutel
AxhvBLz8ausHt/bHQltkSDF2ktcS80svg5y0lBwcmgZhPgsq9T7DxqaIO+4cFq2q
2b+HBzPLRGromzxMBEG/o8QEhKm9QGQ2hxPmw8oH/kFytK/qIeNOEtIOC012i71D
yqsIflGwhYkrGQFeTVfGZfi8gkoCbDXnFlE8C88BR9xhpakpMNKq0Onm0x6oVhvu
mSXYvg9jfKxFzbuH82yDMmPPU+GO4VazQHhCJd2vuY874vYx/xve6rS4LevflgI/
+TsH/e8l2s1R4kr+6D2OvP/MY3/Y2zlarxUM8u73QUnVkkoLamCK+nk0ZwWEcsWk
lIUOEaIMqQRpqBSFjELttiwoyb7uP1ANPeX/PfOj9RPVHNG9fBir0uTwkIv2kXWl
Ooq0HW1FiznRmHR1UUj68EoCwF0LTEqgWMWSZX1EIB4FS5dNoigUIZuZ5vDXTN9C
UlcMnjo2nDVH8lWmI2WBfgo9L/Ff4UMpFxmaODbPiO6V4b+RptMD5Pozro3eL6nZ
qmgz35uYuIVtZlwocB/XGYqPEoz4QAdQwcJiDBDaTtg5/jVIdhABsPUwn9BZohbh
4o439XPuIDV6KYUqiIXvxXB47QDFTSpckaaa2WfN9+IhmRaLd/PHoIazdFI5C1gm
sO5EzAmhfvaPsmFuW19R9pDY/eDfln1tL/jQ1KfMZhXwqLukjninCZni9NkNb4j2
gCkFN2f8VTfMfSKW14QCPwoW5L5+Dhmy7L9eaHWy0DjJrlucSja8mMhVExzZs6ut
XaZfsWzilS1RYOjVMUb15zz+5F+c6+IDva5DhUNhm1mBYlPypT63zty+b0irbpTe
eQezrwHxDh6ILZkkLD444hoMIR4tXBaXiQf89z/JKsmTA6HUvz22ir/pGF3VAGBe
878v0OULVhs+KQVVsmFWun6cxIVD6st3f7j/wJkEDIu4FAHh2sI8STiml/ScHDY+
oOTuTl7upueMUj9IkohjN+41kbzYc/2os8hK42T8kdbPfV6/Vw9pZ5Z4ggwv3d/d
0zgUHwhqbHn8vGXggP1UQ8wK+AFmSxU4LP1UiFLZNwWfXNRnVH1CoFgtfPRRt4r7
ous2Nh+Vm/IjJ+ERNEFFewORavu3VFOe9wS2rLl4OqT1WEavE+rg4zQdiY4zTBbk
dx+JQt4qOyNPHOOq7tYFrjYligTssUKYxdPoCbxF4TvDGB8FHi/MpmsHT015mKtU
E+QyEj1ddm51xtPqH4yWvCf1g8rRxeUopwlmb+XiPLskI2QWB9HtLNtrlSWp5Omm
59DLgpUx14+1y/9G0+u+y94F1z1q/1TBT/nGkLjBBPA/4NvHCLctSTEtpgNWjTbd
drjihQrmG/wx1+zYyy+B5KPSiiGMpWVzEOf9oy92PhOlH0qrRG3gNo8sNu4O4Umn
V7lCdaluum4ISUbw3H0uTZm0yyrsxYDdxGQ08lgpA4w8KDL4MFqMwN8CP/fkOGIz
JJdY/cLA2SaENM92/mWQOTz8AcvuJkLWaDXngaLF45RI/QlUWBgqqIHNHnaYMHHT
moqymqPGMAIMV8uD2y5u6PAlIqeBs2D2Qgh991oNMGe4Y6ZDmej2nWQfzweE9nCI
BeTDGFtkMrmguJep3GdCbUU5/cOLsBhn12aUU4xd0wLxptIGH7Bm+Awlu/KxUC3V
WyMrOCcuqIvWJcuQoVu7HpLuDwdb6ZBKLAeEuCnWs6Cv+ZnDfGOhtLZ1TeN6wE6K
bEF+z/mGUqfaWMBvVgM8zryB9Ad2cgp/HvPqKAwTj4DBR3AjZjNk/LLPOMQbvvOi
yniyvlhGXS7aAErLI4dWjRCIuf1BqC3rV9FMFwt9Ax/yzvukqp7E1y9Oz5uw1UHH
hGrr+Ug/nMdyM0D93ofb0oTy19ul3ukrN6h6WAVr4KyLrDd1du4/ZRpgKIh4qi2D
sc8HwqmIhdh+aWaa4BaBp1k/e0RuhdO1fWbDmr/cNLf1qMENjaAboavpKkHYpSDd
Y0NkQTKySmGPf+XlhM1pAP6sBR2RW74l4St/wnrIZR8h6wnjFiQPRWfrffnssozm
7NfP1lkP4o7m+2Ue9uFfvK7eHSpCcKnhinVhPUQwhv/yHD8FgcvjSIqjmNBGUHJQ
fu+4g0sbqxU1rKUxAy4Rithypqi0VOwudz1FzlQNcjqaQgLpfsXrM16obdykxhYy
WBKo5FkZw7MGzImrDRodgzLYRzWC7/DQlqa9fYO2yeyzq7oMmr5esNzk7cZBCKKG
wbrOHG7N8WIvxrRM1hA7pOiX3/SIBbIzUiq/FZVs0nHlC/eJL2bJdo2wCptjP/Ca
b265JwcyqI8RamxVF14wq0z2uA/0YVZjQ0PxX5AyD2UaVpOfILnSuLkUp8+9PoaC
TBdFbmFW9QVUgzzD8skkkXoww2o7Da9rcniPde4G0l5u2zWIPgZPwkGN4O1DwfiI
zDPDuiw8BnGihUr1PoykZ0EU1zLE0tAJsCVqa5LQQLu91ScIcnKTFKq3u59kk2R3
Az1R7NSiufrkO4CUtvS63Gm+UYHrP7QZz+AZvI4eupTBYrplMoL0jnMR53IK0Oqr
VEcz2c1JdOzFc/jfOZ4NtXizIPjxo3EPjDlJCJ10jLs2+BcFRXk0miZ3CTpYcV6A
TY7opa/3mWbhfmswFc75p1bq2lUTL174TWEXUQQ0fAf/pSaaVBPaL0nrF2iw+Y8e
vbzTLvK1KBVzbAxW+ozhSELpAEdnUO3hWBC2DqgD2L+1qq7uXJIeR/gOGFeJLuVW
54n0REtUyV+ac6gzGCBHqMMcwpd+KkEuTLEDVHiHmWn6JV8apABsw/Q3hHNKeSIZ
/ETFzoa/MJf/l+g3FSE/AhRDjvdeFV8XU38hABj0ZmhNlDgxc5ZcC2ulROvYjq4p
s3Wqh3QrDgGghPaWKql8xrL3zoL6xSvT/MD+mJKp82amtC/srgBOUAVSuc5bqchm
MAmDCX1T/IrdFD5+9AnvqZZ25QGuPmDcaLs6cLwjL1ap9CrfgFe9vzUC7Oz+wHB+
MuWe9bgTagE99M+/WnRSf57v8+NS7DQfnzGcLvt5kt8zWD50Z0a+XwZbcL0q7Jvc
Yk2U+chPG766lFvOJrXqi2r5PTQRHwIlKb4k/GZ2RXQ7imY+MGcrQZK32kgrER1E
aD4aHhT4FWQO7dlBF2p+jx/2phx0EOfSLv9sndM9M0b4Abmq0a1FGzEwCzZwuWNd
BLD0CECkck/L1SXy+Pf6HhTUC8R7E0aMbPKEX4JdCLy6nuA+KUECIWVGkQEEyGU3
7QaV4h7jr49nEa8AZjxsFqnP7Hq4axMGgj1sBWprQ27IDHBFvc8gAd14Xlie3E7V
KHSA69WUrhJbwWQkYVNgnhYW+7UxRtBvGLBsZQevnGFR9Pu8jQDoHe9WZcNRAh52
q1ZNDXDN2ksJbfXDmlHXXL6d60jn5Dq95DD/Ro/d6yxXQNjwXL/h65v2dQDLV+/y
Ka5phvI+O3CU1DIY9fR+8I9ka/EwEpayIoKCHQHYEKnmKfogZ7qGcDtxzJGmZBEb
ieE/NNvl2afydToYfoxRZiYXBbWZ2lsDraFkT7rDHHTHnXZx61lkRX6IiiRCDgsG
OC/uqrn8pUmvg6STfOLC8CxBqP9XCVTtYGolcujEOS7GxU/6+V4OLh/pFiV9UP8I
yQFCoUlFCgLsJTziyFGiYjWXxyogpwMSTk7g4GeT1vvbvuFb0V5n/CTRZjGnyZAv
ystoxS+Ig7d8Hl4ddEEFfSklrAgTtLZj0Pul280s0O8Zh5UhUKl4sl2XxtXORuW/
jeuJCR9ygAllzgleFh2O8ngkEkl7CpUCu9WS6nvdSpmXoaoFLTJn3bS/0zKph/z/
Ab2w7oDbs1MgMGqLLZWBGGrHp2pTBF6Ze923hSfNzhk49sk/NaVwNlvJS4vaZOQI
7X0bpQNTrz2UzEuTqozIy3/wxHllrb8nWxq7QCeJ5EI4+V+hqWPIqH0lf6xkwFqm
r/0DVPhzXNi3gasqUG03NCd5lHVr6kOMNLBI3mE1VJ2kVe6tXmN5XCqRiDKH5Ii7
ndI01JUGKvrpYxbfyKy17+v4n79nal3CObSiXu2VgtTpD500YrcC9d6OP9sr38u8
l2HlO95sqQqOIt8yFTEvjTEj3U6F/nDJgm/l4i2Ubwqx2nWn+alJSzM9NIGGn4JW
NQoUGhTZ5UeDwaQo0/A34CdlP+wlOBz3i/B/MoOm5lKPzkFqv9xkaeuGvgiGad8v
atY6LVVViHmXfAngu9NnhiyPyKUBfDFNt47d2M3WRypfRBSL7k3AWVIZaYFON5o2
Wc8BmWpUhNuQZVW+XNRn/lFlVYZ2NRE6ecYFvJDptmS1dTYphXlNeKfYWxmFEw6W
0Z7jou6LTYalRckG/gX8PBPkyAR2r3ZRpBXHaGCPX0k5gdanuEOEQIY6f3iy27Mn
KhXSGVNELo8qqu5rlTMaS3q2Cw0KOGKiMbwc5XsiGjF7MBOqRIuFEUZerBl+5Zpd
kH9Ru8Q7LQoupVoRCVTp/zm/jhozvO1lLYeX0jaM/g/JbnUK6OQCeAVrLJXIUhwl
KIrUpM7oFltgRF9oZ5UbYZqHBlVFh5sYiHpfes8iq3sQbgHjglaVmteCbUPR+tTr
ctC946OSmVSUWfjmuCRoZC6jiFL0S3fYNJIoTsbzUBMc8VlJIhbgx+mxxwns1fij
nmlCCUBkxfDXUXZmwcB1F+J9OX4qVZZfinub9xt6qxMM5OHZl6N0YDFdKanbMCjR
e0Eqy4ukuinFLxj4jqxofGTk/pQGYdkJyIBj1b8vcBbaes8opFRCLBjg4TSkib8i
qaN+9JfADU+aOs4QatUkFKgV614U4s+/5EY8E2ZvATegYKfxCrUFxhkf6r9BXPpk
iOHVy8lET64Su8Fk6yQbdkf8gUOSpwqgBanlYHJ7o2qM6kfV+dOfC+2Yi+5MwiRZ
1ZaZMzHdxRVX1T5ZIb5iWJy9oguyk0LNEqTcS4UiS6OyZJwSLSY5cEFOXxrPCHj1
ZfVNNJezdO0uUzcZa3P1BH8hf7mjPVgoFrE8Dtf7YzdgJIDmy2JOYGj5CaU2XIWB
SENM5a78rj3Nyqs4MdkJcmQ05T8mzU1nv8C+e7sGeWYbk0jJSRGIkm28AY2FbC8H
xi2bB/Vizb67+5PSSr0ONIovLlE1piOjTvfgGd0szXGrXfGZ7eVrsCrMof7HDFDi
Drq5YU+tS4SMA2otc+kyIcla+lDREbOc8q57fV7mvAO1gyoAtUWf8tUubcvfO7WT
q4qppoysA4yBWu/Tn2zWBPJ8tHAb027xNAXgPoesp0ovT0Fi9vDNdNDHsh6CtdBr
f8Ua2k5QqehYiD2h48S/hZsT/BJSXeu71S1JoGTx/PCeNhbIOpnNnlKlh+cQVnem
D8zjVX+EKa1+viaY6ktgxbslQs5Ty6lOlfqssD2/fSpOdnRUUZ4jiiGgxDohfZOM
W3oLJqicWLPDp6u3hOxc0QgkpLDtiBTZsOAE8Ipcu13ZYxFmxBLr/MttlXYFOYhd
opWCCJ4qr9u2r0k6NiLk5EEqHeCKm1eKbcWGdB0Faa7NL4jvE50CyDHzbxPiV8cG
t8sL1uh6i+GQhwJY38TehYeEjVV0IloRG1/I9wjYSXXMRtNtQkYrftzlQzK7UN6+
uPrey06GCLvmjJqNYt9wsvUFOd3D+tLn3At/BYnZ2aMXKO6/icqKBMBo5u/wK+db
a7CeBr3QsNgVdEI66bSrDcSdxho23+4V8t+5w+Brab9Tjql4rjBIuXdVZwShsGfE
BhYSbpFG+Ak6PY/sAAfLihpzQ2K2pWUkKLQudCDCPJzZhi0vOcqieAj7IyYhtK1h
TPXQ2p29/P4WD7/OJ1JSHqxc7Ve9fvkRCapojt8rRHDN55Tcn1CIegZUOcHcsyR3
r+JJTsmeSCxJpttFzrK2bCzG3kpDYBPWeQdtztlOi2SKrzdXkHAEHOKQESGYDaOo
th6QDPgEl2ewjFi1QPfhbpNRKPzisIQGw2qHkjgTC+6CJexm+wffWx6akuXb0IyY
g4iM3ZXQODGO1A3Nggsod1haAYC0aqAuu0pJfErGLZjwyU3yMziHAkvDYcogWc+P
ytTI963QhQ9CPEK3P1ovBK+qsSupEkf+6S+wkctnILRl8QgkadnBiFrLsxvLfdcr
rmfJcv+R59DdTuT4ha8v8d5Au9kDG/DB7cvFenWJE6YqO4iIT63lo1pjv1xWIwpH
8HFdMcfA9SBKpY+kDpqaK3FagVY+cGQLf4gFp9be5EJ5/+freT73+6ClHy4NK02w
ZNHNygHk9+Z+RZz3jQWfamgT5BM54HPBcrHzRtQksa4AY/Tmpo+G/s/3phWZz2HW
hHRB5y+gzi48+3splDuSOi0aVsT63BY2V+DuZ8/VaXkxCwJPEOh9QlYsciZ435Oc
0Ou+kHd5zJ8kUx7odpUr3yeZlu3ak5lZ6M5zXRZFuQzhQbEfHezTP/mZecn+OFaA
vzaaMMBrgC0PPCk/X4pvC/aNNZt0VambeLOhvLeTba9wKbqGve9UZyAyx5CMRvB2
hpn9OOUldx4RKvqPO/IEXZLm6zlnPVWarTF4BMFmVaBJScrfTg2DMP7vy7QXRiwq
G5pKCUQv8NJ9pNNeiI+cPEbxNW8HkM7qmmNfviD32CJvhfPF8TXabVQuVLt+n1eP
EgXRukNu4xoP45dK11CbXN6htnX9UhN4QgAEAG2gWDP0VGt+G+F2YRr7mx5oWPDC
jb8x14NDmMqHrwHNjuYWOYA90XBumvf35k/K0RMusRw5j7PBy6D2NSOG7lh1Q+vW
B5Hb9hi/6jSol5imHxeIlnjz5zzzs08btaKexwSHDQeQSnDsD1GPm5fNfpoJHAnq
cgdVzOoErirp3uLrpQ/6JGfbIM2DP9rY0yNgZxcxvCxFBR1+9xnfNQhoRVwzKgk2
25tdrsQ7t+jDWT1I76tDlxf3To0Enf67Rr2dLZ/7ZcA/zuWSeF71SVIB53sq6qCa
TCzK8wBBMliFHJQnshtTSzGmkOBXbMxdc5Y/WxIUoWqD6JN6wTKqhEmpPRYi33h/
40Sgt+oDvbQQ9+sUk4kJo7XiPC/HtvO0Zpsj8bC1Cwg5IGY15rVBRCxhPcBRuJ03
HmHJYtctRAmmPLz/9qVCz98TlvgkLcCnSt/kv2ptGzu3Oa8xLpXsf5XIJaE3NWqx
WTAVnQlax854Api5RPen1M+0oQWha9YKTqNUPB0xgwas9sa7lOKp5pXgAJOW2dSr
I/d6pRIhiX1hJodXlpcn9NIlPqjGRxZD8WEXIukU8ZQKnjR8pVlVEO5fKTquIQN+
X4X34tx258HJ9KoPlPT65sIWK/6T5rA1+scaiXND25gnK2UexDd/VlEmcxR+vE1i
iqpT//Mu9yCNLxGVrILlJpoxWiZM9QSS3QruegCLD41IrrlukFrbWULBs1DblJgD
0HSqHRLg0M+y1C+y7xZghEigTUXxz4X/lCJ6KeZYjn1j9jLJGThmJT+T/6k9F/GP
EAvw/FPTZCPf73MGW1HchD8872sOBwX+GMyjcpKpQbCOT53WkyO1RnSfzs9NLWyO
2bTo9I1uDycbB7cK7tVX4gdGcVbwYO5DvJQZR6/5rJkSCIZCpAR6qvrJqNH6HK4p
7FBf7r8Ktqe8kRdKLGsvijKERcJv2NqKeTFfp8dxv6aMFopGxga0UzvvfYXHAcU1
gAi0LqN3coNS38yqMWTx9stnMtaErQ6QArfFIux7+M7nCOsdjBLMvU197qcxH0f1
y3eniOInYSMSgz86YEqGeLt6IugmYIFqPTkWPtqk0zsBCkoDPd7yoGYCPMZ/+4DC
twbhUWBxCKC0ERSJ50Yc1ocm+nHQpB5dqfeRDixiiojI32Dk5uLrf8qAuLnXEWL9
/VLQorJc0+rr0aYUjgch4bSU3lhFOJDUcjyKICaI6YiwBfTEFvS1PQI3Z65+2xhQ
cbdqpsqd9jGDuXwU+Ohj5YkDcirJN+Lj+RCpgGUNYZ3GbsY/sPdKjiW8Y8mhj1Oh
6xi7xqalJd5UdBKewVGgcQG3Mw1BmHa86+4kv6nuY6RZlrwBZ/96Rnk52gLz+TjM
q2YmABOAWR3bxXwAdlCqouAO8fTBolcOefgjk4VbyblmjXeEeEP6f6ABNYj9fOQd
kATj2s6hVF9DqMPmR6aNbW12eJAzHzA5nXm4kJ64MzTvai0g8ca6ynb2bG+bQPuo
ugp16/T6ih/bFPjc/m+jMtjWXQ8jT9ozd9aR6HZwHgEDzQNyXG5e3blKtVq7AkO1
ySOzTKQ/AmR+zzpa9RiSM6Z6dwv/EoMjnzreYKF6E4/retxHeBacYR+/1mYZKjjj
rQMmj2PKa5bwMZz65j1rpcGef/y0ZKoWPeM6/R2flNksz40MqmQOFg4olIBwOBff
pHWEO3yvbMfs35mE/P38hxWgEj+ifO/p+YphAC8bS74VP2q6ynb0hEvFxhQ9UlCT
/ZslJBL62jwRks8Ymx1zsMSKcQAgUZGbnPJ8u5c3C4Ocmyq757py1EpNhqBm58Q5
XySDshNitXlonDqzXpcyv5POBQ6rnezcoE9qHuEQFTbnzQDW3wKJLdv6bX7l3h01
EnzcX2+IPwIFSLnqxvdaAVBSfdqCX+oUbAeYj13wIF6vVhua6LjP5YO2gqKQbtDf
cgc5Z2RJ3St4mYaQrUXYlF5/2LXzP4gbZraf1rWqMLYrlIX62CCceucmOeSD3cY+
HUJnYBAUHpxydWMyejT12rbzXoW5D3Z8/bzz/f4It75pZCbxqQldHFAK5izgIlc8
sW5aL/11FJG9SCfVleQJeqhEnWUDNX1uv/+35pk5QAJsmymtxdQ1bt9w+GXNd8UO
KN4D/ApMWfnHZyAPU3L+nIQLYUmGQi8DSWyQjDro5pdf/q9K1YPnAZB31HaD6/8S
HEIC+9IlczdEn9ddTt8MVFNJUN0ItGZ33e9Dk1WVePBhRkDJOr/l63cJYAtonkxR
7VX2qk0dotpp//S9iQ42g67Sqg0aJKQThVUG0SjyFzwpoGDdr7hsQUpFp90OkZ2x
pLWAwPIc8T82lD+6Vpxehp3y1oYRwnLjoN81yheihuMXfFuFo85jwjBJhDPgjLCd
EpBcstEUK/5UcwOWeULglbxnFB/xM957qyavaQya8i1GCVbTD47nlHfVql3TNOoo
IHt7I0SSeAv2ohC3hJzCfmBiUSlK6r9yHlYtmSqaiyDRuq6U2GVgleKET3SwnyWN
/Sq1xg69+RH7gpGaGwngjl+HnT5W2r8O45QeNNy3hjXs7qlNbw+UqDRsCBJoJuwL
U0HKpV3rw4ZIuzxG0NCJ0NvfKpA0NpyRRt0d/gi3sc+Du46+1GDTgZmCT1exLqx9
aXP6G7Q8cJ/csx8anhQv2S3ux2rsP9a3flPTXADacnqALgeIYEZpRiMJt5O8WbKR
Zgayf2bB8RRgm9e8/mbeluV2JVnw71vELLCrhdO5MsBkOMKJZV03293bEqjcrYwg
pRaZC7fblYL4tCGZ51REqYZtpZS+gW7/8IXxMuCY9iEYS4RE+Gx0kMpeM05nt2DL
wOIeVWApIIqNf8Z6Xv2kuUSRs8zcLX+ezz1I/MCKREfmmOQms0tPB+CB+m1qoubN
KIk8UAVxDv/PaaLi9XJOGG41XNGCVTUzW6jl3tWayp3wZ2MxVqEtmbOl4UMcJEUt
gPJdmYHgrvoBl9CSk+BL8/7hHwZ9aXvjwYks9/P9a1S3AhkxUDyPZZZFG1ZEJoyZ
vQjAqKmDLaR/IV6JsxeYyiNh0PHqRwdL5AC7P82Wa0/TyZ5dVb+9shDuvVzIeMc0
PBWy9/+I+aSbfgkp4O/nP+mnjgiJO0qPUXyYjoFayEGODLU07R5YhehZZP/foxP+
CXm3hygPLM5LSTYPZc8+C3h6JhtqrvPWMXHUHmq106FLsN/HTUckSP2cyVk9NE3H
IlG+IYQT+lon5FQjyhzM9bqjPRl8bOKFfH8kG6dBDY5hNBQx2VO8jdD6IqIh22kd
9iaHBHr/RFmgfaWnHrqlVPGAeXNnKHuGtC2FvSm5Np8lqj7FFP4F98n/LPkf0J3B
lc6MNm8KL/ftrefuKgK0ukw7yEwi9BsgQZq8qkBBN8ZPA8XYRRvzZe0041/cGebM
186/jTDnaNbXonASk69BZraVl+hS0yLBtXCscqNwJRRyH0H+C248AMUQHKEfJSsg
39YhC8I0hHO5ntyOu1c9t5dzm5B/aTI0JSQxXoraEO3dpg+B7CKmpKVR9zX1d1Hy
0bLcMpH4NovR/VE+AkNdcgOfjGpxP9vCNRHoL0sJ+51v4rrqeayYzV9WUxxT4nwu
gk8OsviR1/RAJXkZYqM2ObKBlZrxkD4wvcl3qa1jYgE3F16gomZcpvZDAD0Z91br
+aVupFof07PRsUgFouSde2KQFZ+APLG1y4day/uBjdqBkomkDwM4Om/cCl9c8mg1
y434Kpb62NAxdttxdXl56RGe2JeOGQaPjpREFJe89VEtkvHR3tWLkIaDfC+LXjqp
0gGCoTWPvoVvxvzvNU083J3SWBUYw19bogC/nCc2QTld5QOao5EByTIGrGK9YZ0C
/wweFkkt+b8P33NH8PCu/R8jP/8CdAvJYsmriSeB1W//qMP9AFzKKHgN74wmUARg
dhsuc/mh4dB2sBfNkxurOuw9wGpnReQ4j5nPcwIcTOmFa27aecdBrnEA32jSQGff
8MJG4ZTCIIRojfqOkZc+9jtRwu5o5ofY4p3SbEqVAN/tqYxqdrfUYjVDwx/sQlu7
EqxUzEPp5HwzFjDIF9mYEeLS4mEWql1SwA/gGlt0Ap6Objyw3Bb7BYjGJHAsjBja
Co/UU1RrQLgnk0WnH3+It8TgGlMOVjoCoD1lRxEhdQY30RpEhH2r0wCD4PH9wgvd
uEF2hApizoe0d13fp5tAU4tq2tKDnTzKP8pJx0ezkEgbMCWfRz8+lkqigD5Q3HWW
5VeDjJN0hrfCsv29+LJJg1tnxhLaVjrLZssXrs5kQYU04SLnGrSLohH5xgV0SRkA
DbPn7jU7jg+bzrKi+QwpPZ4FoHUBMFiKuS8DuQcQD5c7+TnDXzRxf5XQ4UxP7K47
Uz6ynB1uhCYQCOqNjKRKl6sEYTl2Fw7QgdHF+r1o69XHoYFQNzUxp6HEJX7Sh5Xb
uFr24pGgt6ZMOokpjVSBH0IlZhL3dMPwBLcecP7x/cJZ/kbpkbSIF7mkxvWQ5Cww
saarNFp4ypGnpicQeEeTS7qIaTOdqikJPxVenR+C5+6dyC86k2w6Glh8rne3lpJb
Tn1ln0X6Gn0qtLqZWSkCzR9hX8RSdP4a13bXtAkR7+Gz8oOGtJCKKnOjHeV+b2HP
xFAL/fSoO1L3eT/eGxk9ciIfbuC59uOVOzjSaec/APcg1BqV7tFWZF+E5OW7sD/f
/hW7xmg81soIe+5oWUHiijUOZ1KcKrFoBT2F4J39ZgTp+TmJF/KEmmvO9UmKg5bN
1yTq5JL8J5Vx95uhwcedjspi7AB1qutiLGn27DGdZbbVHx+Bg3EN6KlTvadd1tC8
wv3cpKZovQTv4vcQI0j36ItPNhPVKupHhc1wAiOpAPndBnCIh8dA+VqfLp8G61m5
3N1owqfnViaFWmZLa2irGLVDBAllB/iaSQIcQ27qp11W6IfEeRoeUiMl0K4bKdpN
Pf2kEzLyL7jy2TU9joDtbTGxm/aOyJau1GD6AyrgLSL8VpKK8fDcdhJcudLimvW6
TovXxgm1G+GeTFYu0pfH6Tf32skYIjGBHm8NiJ834fBQV5q9dTSpRrvrKhz6Sf+s
+jAjCu1Jbt1gnQEBBCisPW34FU3RsfPzUj0u/F5EU3qsVWKQxcnanhZh0xf6x+1X
z1uYof86TVpXxKCqm7TpomND2KAR+zR5KCtPu0JOTvNuV/lIZRkDTfo06C3OAUDq
5ipJ0QWzMBs+FZKqcxODKwEKrTz5gg+lk+AAVWdBuVw1RgwPXGdwBkmTMJlcvF4z
oyeWhI5UfVUoCYjT7jZ1RWigXTEnDoX1PgstB+EyY62CpRjl5o2+7eOqRnM8rqH1
uxefebI/7s38UdHK0GZvHqONOEClsrSKYoCPx8j6IOHxofWPwcIE9dMC9jsWuprw
pkiPVZmGEe/L3DOzfNuXGQh43vhPudyPuVYdEJnU/cDuuvbWzMuuhCpz9A1gljRV
FHJHk5ACi4ZdQYJURhYO549pltmmZ1aZS91/hxigeG1QNWCUaAyRhlZXXVrvSoFm
0tvda1IgHnOL3WmNmLGmj9dGKlHBnEkFAqIY11aWVYo2Bvph9BX77jE6RRUSpt+W
vvxEUEpXBpZr1M33IrwkDsfW1VQTgBpYsWBVQvzG8Yxa981NPS1KR4xkUtRK+LHE
C2BHyKdlINOoX1Nu5MTKICz+80zRaMq3eOthr7i3WQFzOkS2xNpTwxhVH+1p/Zll
zztcPHKTqg8kxqUtCdqalKxTWgsYX1iOXh0e2TFDJYapB7NVaIaVWOyOJYXv8+lc
f1Yvl9GwjWV9RUozQb6h/FJ7rgvu+k28roPxPszCfKRjjEFu9Hlp3rfl5GpW3hEG
Sfwuk9FoUbBsGW0VOBN0KMqAClOO4SGAW5thIBkeAekAa+a6+gnLHpfE7a0yQ5uv
yqwnpXTX7hAISihf17p1Oei3bz9meZckrfFY/CDoAenxCR2kIPOAtXK6EgEp+Jzv
xTjJ/M7ZZRtZW818aSJvGOmotVd/kwiYT/1Ds2e0WtunkH7IsnzEKSSwWBW5MA5w
EZrL3efDRYmhDUgy65GOTyfHJzJyQgiinGQY79BgA+85DQSrj0qpDYc1fNZK+rXP
5wW+Fos0L0r4sqLN34NRJIhIpRGHY8Ej0KluSHEeeIcSsss5lOUHGLWZO/wz/Vpq
pXnbhlj7xlx/7unOppWHFNIKFBLsFQdiKW0u9sYBe/yHgZk1cxZYuBQTtJpVLhp7
UAgY/H5o0/ABew8zZIs2dBYFI0PYZYtUJG8Djho8aVAe4xZfxuuApQIS3JKe0iLD
tnqipfDuT4NPV0PzEpmSvMHo/+KH9/L6fC81hVcLOv75kgeVrxuMXE10XKx4lQXV
R7tkV1hLq4dOV9uBDvBxU4a9ohcza7UNYOyKDhlwSDrfIIgCVoAjNKoQV/RQUcUI
+kFPm1cP3KRxcs3hkSEfWMLQve8rztu9e/7PxmJe/21yZBqssXRtY/VTfXHW97cy
igw3v32AOQUWKfMm+OaTb9Xjlcs8hcFGpLj3y9/nk97k+qnK8uFeQKeXEt6RRheI
QhzVs4BZSthSvFoDZgX8T8R5JDDvEuBoPk982RqxEdC0R3gs6Sr4JWrd8zDyVJhy
dh81+0/x/1b5IIdvWWp6VeejjOuy/AtjHt7D1zYJhWRUImxHhW5Zf55eCOxN9MM5
xd+euqc/GrAxQQfWb14cKRRs4iC1pxGhkDYNpnWeSHhf0Wb9BR4LG9p2zmCcMoQp
CVVgQ16MhfYmQBlYCfh1H86qQfXjoZa4+mCBaR4ZEiA7zsy4n2nSXzgvol7fwHSu
BABKq2+nOnNW3fstgkQy5OPAdq7PTRGJghdDrUlkw755LvE3HgYe1fDfw4rrHdI4
vyInidxRJnpkiNsQhDsfaVmK5cRq7bh2AbgeWYD7ry3k2xBxtxhXu8Ks1uRZyjVP
Ri9AeJXNNJ1Cm/i0CeVTokwcYSMRIqjlPMQoJca1opsfsV/5wrh1hjY5wWFzlA3B
Vh33lYsy3AJqzQLYauCXbcDeynyYIdhAIgtPSKaKlJdL14Oh+ojVpjPLmjETkIoP
mQat88Itsna/IfYEtW8jQlBcTVNbyiOoUlAu4JvRhb8GFGgBASuSxb09yaCkHmV6
nRHuQU6pJDpN+jQ7c+vxHnfgyJJTi+zl7GwHKvSVMEgstr/CZ7W0iZ9yW4h0ZWM6
42k8FxAqK7D75USOPSZVwrYiCYS8l7VXOOBLSRC2luvN7PY5nnj8AW9oE3Q1LV5C
qnm2B+yDBkXAxhix+KTYxNzv6FYdH4UPOvNHRM2NbANL3e/vzetNHxEUSp/iOJIy
zfbjEOhQoHVU8g6Z+RemkL+koFcXCQxEvt+opLdk1KsG89pyaLS05qs5Fz0UIwsO
RuqZOpmVq8pf12bt143FTRhmISsN33qW10rk1qCm61nJqFJV3MuNYuEs3m4QjBKR
Hkv7UdkDq0Vm+DWrgVsRYUxV9hw3jFhkuiQ6iH/vyK4Q5puD53BB8Q9wOkJCji6w
+yZ3f03suiUCc1JjnBdYakpBA1XLFauzDV1j92XSAf2z4KDf//9P30Be0fgLst1f
FwA9Uo2Xh7NCrtmCT8nCWIXVe+nB2Pejtopj1cSNuu/2W4P9I+EJPqI1TfUrOIbU
H0lVoqKMO5e83tAcmBVtQNNJwCEYSmMNdd0F6LSGkkgU+DUSNj0eDS++Q2plJCqI
Slqk1RRXRzyq43VBh6jMrvBRtnGRsUPWX5M/QVIWjBAP3appnd8bnaw/xpWvqbct
S8GBZhuDuKxf0yr0e9CzM3t9wtkes2bCftOrFhfzwgBSLkurPE2KG28wVYFi5SO0
oYnLMAaB9DkPnTH/TpRVAbZeOrMYv6e972AD3kuOgF+wlF0jwcdus3dTfEVLUupB
1dDWiDy3lN7dtDAbNT7EQHdrgz65qjn6HfSg3LC41u10xeEQDHbGYVdyw5MiD/0m
HzcrExgBMUB9ED4H88k9rm8S7eJGr8tLKbMjV2OaUeTn8izxlDY85Ze45eUy1wCs
GuX22cJ1N1KD2PpB4KXYrxA94bmxRxafNMQpwYPoAlbZWeV9IAT/keWBOAHXlpRQ
+YMHua/RXGFtRou9Q13rhRrepy1dKtZ9oFtAeRR3joagFmcmJ8JIabApn8C5s+2b
Pg5Fb3XX3hNbQGyDFkWF4VAkYGTURpL9UJ5Vc+NS3Svl6ZvuWVXo1tvpQihhIRx6
OREP7qc0G3NZAoDXdWTXH7hsYzo8W+2p+NigFlRav469p0ymlXNw+721B62PS7AW
ZuPrr/tjfdjorG74uCcp28r9hU7O+qNmnGKBWTbPmjRdbjQcOoRRy5G/gjRxNn7s
bi9wXnMAR3e9MbGGWMAOkaHw6GrxwIwdSt7fxV9l4OnCBYFadwarF0t8o7HryXgJ
wPKbHE+RdDw8Xl9Mk58WweJzZkO5TDG+63P/z7uFXhFKCNQ80sryXvbPEBe6+ABa
TOpzKfazNVyhKeT7rDoEq23JHRgSAdg0gg6aUSquGi9RCxpkI270rTBH/sPehnj4
E8hCgiSOWnq3Ywgh8M7WsIzTqHJAfgggybLYuO7y1KgLvIQ6MJ+/enkPpANumU7u
dwBXqwjrSwOomMqX7NPr7B0DdD/EhCCfBj0H+HCydJyvZf3hqDf/g61B38K1PnN5
Wztg+j3/SOgSxcP+dbmcKKIZAOJUO9noT9OfG+ujlWiH/UE4ygFY0d8j09IvvClD
oLXQJCjf2g741Y2lZ1tUNcfzMmdg3YMLhbKf92XXMylKDhUbVr8hm3DU6LC+YIQ/
Eod/VXOg1cxpZKemvFsGz8IvxIkw5isADIhu0eso6t0Jzi9rwFeoKVNsjrUo18Gs
fk22/H6BTyFjMm96INPIlw7rcTYWC5k1F+GyRic7y9m5Dw4Ktdejz62lvpIKTBpC
wK8Df/wy3TFFUpbp+ZxsyHKn91brxjUr9jjVWzbtp2/d5b8u63JAEqy6nzxaBN2D
RkQRuFu5lnByqCSyMre3pcQXpDGg4/tOBRkCIc1qk9qqj38jQ/ye0QIF2/bkT37Y
PCVM/lRTz1LE6g/JqUTokdHofkgAd+3gZrzbYTHnFswYrYA8WkiI0EhBR9LseGYi
mK8OhQ5lCVZ47J/9id1D5MuFqsDm1WHSgcaPo/7qtfD/EZxC8VuxD9SywyE5cyws
MUivN7FqiHeUd/TnQLoTqIxBtVTFfieqhY1kxeTs8Sjs6fbZgDQ8suFpXC+ycA7j
SysLGxEzFa608T9CjqWX2tZ77jU+k2hZhXqJ9X97+weEl+FXGEAsiWcUxTAElcmD
Shmg3aDn67gDaW8Zi6JlDLVIY08YMAf2mN4jFgDm/1Lp+rGZWCHF6QPi0bqR2/wu
xmMCpiApv/6VEx1w3uhjNTwMbasMfsklsyhjqqCo67ioOV0a7BtPql5et6WPU7U4
rZ4hf/8/8/Obb8v7PCm1PM84327u7XEqHocf5HkHoZ3ntxpm/i5bIHuX2WD35RCh
H4aig8NIIS1DRGZYDVHlNnsMAwQFnNjLWtE0aHFJscbJku2NDGqZYZSQKXhE55gp
O/EKiQF9+waXjrurFWNbKIzeBLRqf5giQA9UOsCgNcphrNMLY+oca3i5f89epUIP
gnMNYLfa9ikeWC3WRUkWIOq/Hu7zV/79KIbG9/O/90b+x/W4eO6wZoyWB/Z8vyRj
w3iPA5IBjZzzddq7+DYurIHJ4B/SRqdcc9OPmXb78Nawr3LDtconte3lda86A6GU
JdCcsA3US0ShguznXivtzAJFpN7f8s4b5ZCfat5lqllEnlggcPkXeLbh1yOXDO6K
0VrTMOVxM8H9NDxMp8r+5I16PTJMmvZ3GEy1VC5s32d5ekJMWMtfEzAzHitUNpJW
0SjgT1U3cIOJ1W+Ydmzwkj53e+8Tk8wLtkmY65rymOmQbURMKrdW4QoqF2lVAv8W
2kuLbhYSesRmAni7hIceDbPfxVAizPC1D7SuxQjSZJIgr1vbJFW+YyBHmM3H3KA/
QHqoXRjrC7C0ymG3mLrIu09HmmkYETFkbDjnC/w8320ZvRoeOuRntXACW47y35OT
bp1PLBYMYXa34iMQqRzYtVgFIhvc4pX9KKo285VkwRBnmzt3afIScHk1B9+pYF/9
OM3ptpKYT6oWL+MTR5OtiIDffyWcdMGS/cSBw8SajCmygXkbcoSKZrFIO7L+dx/q
cM+6iWpsOxWQUsYvx2FwereydaGO2w5gknikMCkDbo7xINiC2snSnMbecqER4NsX
PMv3XfkmNGYKOm8/7VRKWqEZkmQ9Lk8Hn/9C7pga7fzmjQUfoF9viVJ8KiTdKYxb
6Np6LEMfmns+fkLZ6q+rLYc6J71R1jViUR6JNUssru8a4v9IZAF4XYkiG1SQFxhv
wyu3I2xCh8qZguDEAKPi3oBC6/lUG7jVgYGg3V7hE7/yU3n6XAZvbyLxanWYRcms
etLFlkQdP46SIBVpjVlPDJ4rqu+i8QnhJaBzz+DlD610fxB04wORCosH6/DOYIaz
Asx9qF8yY6F+ZFJ7a/tkntmKbAdSdpJrTfPPw7HeuVIfFDTx80bXaRRTBF1n6ZJX
UHUoaKP5Bi8W7eAEXfePA6FtB0fAgETECPFQlYX6sRPDKppIEyRqL0TANLfj+58p
IEuJ40V1IH8PoXzticLM0y4sliSKWJ/RTcDvZ9KqVim7uM3rdFpGlpvMQbfys1ZV
uZYNjOjEdI74Z9msTURfcFO9aCtI2npjPix1vIJfT30RbOZBgvpYerJ1AaX0KIeX
Apy4bObCadS0C+NIAgWXQLBPgm6q4OU8ZXH3/Isxe8TPoZsY2IK2hcVXd6nyGQwl
llpnIfD1qF9qDO5bhnanKC6tkY+PS05GUFsZEZi027YAOIlprZ35q6oqLDu+83fN
Vvkgk0hVHXercgAC6alJ+kj5KjuXd47Imv5E+jiU6ByTJuZcxUoBSCb9tDqYhEsQ
N2kJH6sc2XICOhpmAbAN/2itJfl4HbDYDufrOVvYe1LWzzLp01JSqGQm/FQiWe7X
h/vpNbqN7b8g1wb7kZyv+pLvvaByNEO638/bZuw1fa/m6B6QbAHEiWMY5Cj2hKne
SBRCKBRibeGgwHOOMVxYpG/3MvDa/BzneV1Ab4IxYNG45+0yama6aLQCqRAA8eoY
+8J2u+wI+lZEa4Bnk+mbyyrDx9ZYx6Jh/Vkvk/LDf9JR5J9bCWYMcNNRf/u+iPhI
D3jLOQ9AcfaN8XjiqmNRfpRoC2WhTWQA44N25pehRua9EccbE3CnX63u1ZQAydgM
QEVP710oYZCGSStaXieLz4UublMwQav5P/U+r79YAiOzlw7wYiSm1MqkYn/6rqlw
A7yBr6YSn9UMs9T3ebJ9WJ//lAGvmGw+ebdXvqTf6oEu6xPqGJsBn6HZNRixI3q2
qfL9I333ZrgFyqNxiSOD0k83UXjO+Hq1ptueY3sVdGxEZh7+bvQtn4Sv7n0rsUw5
lqY2j6LvyrS034uD4bcU3rDiOVbAGoFpQyv7W4KQFayYI8OtajsdTCINxUg/+IL8
1TtttOLq8LKxvOwVIQpRi8EKvlJS/gjL3wjmgzkhuueMniARpuYPpu6+wqZKlO/v
coIKULPbtpUwNm2haADH0A4O0JHzGAyX8q+tiwpvA20P0lljbvFOefFKiPK/vDna
fLJoWcmw3agPmYfJTmECmAMJ73A+fkIeW7/HAkeyojjmwcWaFcH4NrlAmv2pQ1xu
xUhADEjaUv/YeNgxz2cwHnPhVXdgky1zpRyb1B9Mf3/chJLzcbGlaAg4tio+An7K
/YtCM0xytAuKojA5OQjyE0wnblRaq+yeBI2qxMe2j/zGjSjUEtoNu8jHm6NxTyBL
S/U0rZ9hBjeM22LpZu0C/7B1GtPyJwmLH9dAQEqpiG0oQ5BK/vCB5lP+mCkn3Ykm
zPyrIopazru5Tuvas0Z0c/O9eMI0WtixujNDDtgch+2HRqpAPU4TLkYmk8XaGKNV
fGqU/LAGApH5kYxwM02ei+YwaG7oGTNlKdHIfiXuVlcdpOeELCTMWP/S7ZUD9XGV
MRmdyY72XDbD9lVlRKL9vqCYN6PFax/mot7gzBwsz1CcxSPNWAz9BquNWHZpqmE2
n85xKUSe3nQ2u9YsSap+k9iq1FnxBsnckqaqR0B6BxCEmMwJMOjumyZkSMFX+W/W
W59qDMKyEThu55SElii9MomAHODO0IhjkXlg/Yeht5O25GmaV1pGUIDtNka0maRF
3F3g4Fpq/5s+EFevjke02XD+TMK21v2oY1zHnbiFHCJR3yjHJsJkbsS3lHzS9Ih6
bToCdnNl3Mws1QLN0NTlCAsu3TgAZxTHj4+3s5tQFgVQGLs2EmBjiqbmEkFkjH5M
GKoYjlnBxP2xNc5JSDpI9NOx95FfWY6D2EqGxzElS91HJKh8fBcqs7532CzeQxsX
/8hkqacn9ENFNQS6aYuOu2fSOMEHC+t0Bqnyqu6YH/qCIzvNxofk4REeL901wWYB
XJ3zDWFU7tqN73PuAjZ3ZF9rfm8dydlBQNF8/UBi4PRkKRajdqHpVyEQIzwod3pf
lGnPXewg4Z2PkXNNY1mKEx2XvIE/76XjJ4ekD272fhwiFIAfGapa4SgfAupCzq/J
HFRRnJawh60nay6vIc/EcMtyObnz9QB3W7buMs97hjpSKP05gn/sCQea5Ae5cF0l
bn2D7VabeG5GQWB26aOMM7plHjB/wW4e6plGLMeaANc48CM8fX7ttSue3UUjzWQk
OtDDk0Sz1rrpJMlqXgwN4aZ58DM82wVg670vPGdM/0GCKUERtaq00nKUhx9XtVMU
ddhXB8aRH1r+hirqWtpDSBXqfMQC661zbrjP05RdJEBr8sL8gfsAc0SVjgd7m3US
Ujs3vAaFjn4h0XNLZBc/LiXesoncYs7Eka7Irve+XzdowZrz6T5SZhsSCx5jOjmg
XPHeoazqMThfd7ygbWzyoG77y5aYBUhwxQIRM/tp/B9mBKfeMo7FUQNDuRFogXYp
PeAIM0lHXb64wkrwzht+ZQAA3ikKuO6mlh3Ign+TdUvP0LuGkE+I5TZ3OnFGGPsS
IkdyKSk/VKpXrls+KTeCJQtQ+N07i8L0hm/Au6chK5TjInzy+hpv1cSAZ/vCfagB
acO9lU9FNuJ9ihOVmv0oAV9BSVo2ovvPUNOyk6uRm5sTp+o9YWwAqos0NZTk4fjS
Zf3gmjeHK6mWJZY/IPSXmbjgTe2JupkexybA4YoqLr5yaCjfToJKp7NBBUUx42qD
BPdmzN4fQYviMeXRRC+aNOpxU4IjmS1xaHAcIXrY8y0TO55QA8j4nuH3kDbbqwHf
WvkeMVoW8u2UgLTTcS4J4qPowfgEFcBQvORDpQfKONWUXeytRZlu4+oBk9z5BK4C
dpwKrZ8uvGgFog188ebxbbUX3RB1f8XwLI9CRIyDuxrHBVnk2k8ErlavUhe2V+DS
thqQGHZj4BYtSpEm13EEp1f9ZFrt5H71G3Idw45TS5UkhL39cenRdIXh9pudZdny
LURnLvYvmnyFny5ZohAx3lZMtx0yHAcak5B6OEsEc/XkbXIF3tTbwRByENl/8YIE
SAvveqr0F0IzJynnUSZ6kDXT23uk2UGyXwi8iv2UZ+k2yagcsnJMkFfCHz9iqWOa
TtYL+I/wqJIs/ChE6sFXibe1shTBqNRv42B6WFgmvz7H7rhnjj7BYi+JZSWJkhnr
oR+QZI4xwxXzc6QdG2j3WsEFvkeNytW/WOgSFi89y772Dw5JS7CPMfZjgecRfjaI
SiCd4CS/+E5MKCQA1ps0vyvg7d4Q33NjC0lMblBJ7TPG3+F3pbzqFdLjF/zdiTpf
KqRrQwDf7RY1P6uUyqx6vmJzzXEkwzZEpMIwD1w6omZrVmOstpBkeOoi6V6mkh1y
Xf2FqoL0autGGTW0z0HNxhnGkdbUtSg/Jfh19mUhYfZwweJD1navTXW6/tN19awJ
X2fnQONouUqoomrvf7szz18jBJDR/n3KeGbeJ9lI3zsi7ak1M3VFaS90g/wAoFx6
qIX29XpV1a6xRarX2Hdnl73tU4Q5PpL7u+qqK1NO1JtUVNTkWn2rxD+u34LVk/IH
OeK+Zy3M4h8zh+cKBvObeSZLRkGiCKLlWiKeyQKBaNje5x9wlG/2PbLdxd/MlRtn
wiWzGodPT8dGrMXlOw1p1m09TpqS8JmukNAQR9RAI4GVUFjV+6sSaqawvnoPFRAh
5y7J/Ksu7DKy59f85/7Ef/FL7AnDG2q75GhgPI1IfOmTShK9aovSEChUJ9gTzP7X
H2bLHbk8umJbWdz4f1/UWUNnB2YxZ1S5o92se4/oN+Dyeqf5+pHaXySEZddt9zfN
YUN5S95zZ7YNNhcWei0jvKycVTVlyBY6PTwSf92eO9MIr+FJsyQoqSUTbfM9UqyS
S1x0TNG8VMdg6YiNPQTo3NS+JzxGe1XqYh6UjqS5tlXjgL8FHgkbtGjZebzsLrcr
LZpxIzXskF+omO2egWh3/UJGo0U6AkWXfaLTfIJkyHI2Js3Dre6H2IQfr6GlLLTY
MvKsOJVP6xopBgE/wzlU2UgkNG7vwyiK84Bg32UdmBo40tek9yyXHgtKZtxjwdzG
DXfGuGZcsOwMNKgAh6rDueNKBp9hfUDwNaj5ffEV1N9cW1Uj8IAoWEUg4Z/mgrQc
KQhwM98rYs/WoOW+gByN+oKm5gWvP4xOojAc4rxVStAgJKVMiKCirVPx7fl9O688
PD4c3sekhJq2jBegkvYBLHRkkHq9X4hGvvR8LCI15kO/CuJ4bggrEMhAfy48CiNH
9Xp7REfHtvuzBqdR3dE+S4YxuneCK9CtY3A7PAGaESHutk0J09QTbVyhmCUcCIUb
NwtTeSD/f9uByLectB0DHSo+uE8CKL1BzKVeUKjLuFWLSnZcmVnqZ6WxAYabP3TE
Jp3RAn+RiWbov4xr6G7VDHYx6G1+I4QXUG7WZ1VvqdOIy6pC35G7Naq8XtcTwXkj
5mW2lf2Z9Q0zI0c98xPCgQwzbgOCmC2h3tSKzL4Uy9dXDZjIl8rpgEU7aIJ/MFdm
KZ0ppaM+2b22BVIDB1TDOFe3TUwDBjeHYE0IE0okqHYE8BrmUud7/MN5xzwvQXM7
Lrx+2qEfq+KQ/BgWJ/70BPKqvWVZiS6m/UdLD1Ry7ayqakrpGRcor1HaXpfUfB64
MqtENdgSOINZJeKp2pSYRQhL6UBJfjuPF/AS8JHH+aouL59j3cINzri/hgk3yhTi
ohl7GMPZlbmyAvjTyJix/j3mu4ffg84zQuIl+NP6PTAisrSFCZFilfKlAepwXoLw
Ja0apQ8Z3iFQB8fhXadpPzOb/79Ymd4cPzPyMvmyqdmCye94NkOKLpG+QZzQd/uh
QIcTy5QBaRh9/GpSivEgHnL456HqljnQ8mPZg1aPL7/ew9q36VM1bZHf5JBHUbNO
PlCmGASxBXcxFmZ/8OMVLEctM2F8xOHwPbyqOrLV4nLTeV7Q8hpG/i9mByMT64sr
bqzxlEaoac1sI/AzKecOR0J93ik9t+DLibqaoMDc8CrJhAuRg6Io7jQ73HHrGLxn
xdBHr0G3WYHOYOp7GuONDjOV06GCeVNiVe1IT9xBOg4BGJ+Oq7W3nL9suLCHofBs
DdJceKC+QUmjwz8+r0rt2L5WS5dkfdFirOgTHEsAaFzoqPzUToSgbRFgneChAiSK
NpsSq8unxcXFK6pIHWLCyCAKfa42yPs3lcLg10eiRaD+bPmxGH6UTqRzvdGkWc8C
4FIR3HkkaW4o/s7XHerBK2x1DHbOwoJqOmF9ZpjEkV8adVGUhBL9d65rAElD1rMp
70vL6PuvjZCfl+8ixT7XUiREBqG9rScdEy7UCHFbdLsPGPVFH3NGCEENPFTd7Wuw
s6/Fw1W3IssGYuBLGGSPAWZmwKYlWn6dBlaEkBu2oYdsghYmWMf/F5fFBrdwCv1Z
n7KXr4X2hnXXsy71/cpuE8Gm9wzvRBXjHLPlKT/lZIaVIRenaC16QjRpDWxxYNRu
DbAax9iMfVOqZkJtxveWk9oFnyw+S19GoOYpphg2qwdriC++lKReQ2xGuvoQmgbd
cGiEwVEKmWObMaDo3F8sOqx65plZL7FLnBUsQ/4psxqdKm5HnVgksOncstLFiY+g
huNUKikOW1Gryh4NVZtpcjcyYP1Y2BUickMh5cI22dIVxrStNHcZwakbsDOAALLA
+AlKHUmgbFdKwiJXc+j+mlEFsCVk6wc7TkgdVMVK3KT17Pa9FiIhEaIJMNgLv46i
msmIQg+syAhOqzSZfvOaUPLX5o5yYNc1SUIKJAN1xkT0i5EtSiGAT9seI9xQATjw
uZT/wLqSNyjp7zrrhoEhpqIAcFWc0LPk21N+x68ij1fSCMFCgEFnJcGcLaq+PxSR
vQ3mPgUDs97BpAiNPSuGIHr4R7KICLGZbxtijCGC3mBXt0uU9nEYADjlq0E21UFW
UcTf9y6bK2WhskXIcF/YF/d5RXhzYrGVaKw/bMvLIt0AZuPHC+Z0YA54UWSTBkyH
oq4Mu852BNfgTCuc0bnD+u3MaLl5+hXasSdTfS3ZLL14GeNGD+ZJF5CcVWnDMZik
FdO0gc9UZXXJN40A+pvpghWY8MX/3+IQYRlfNAInX2ZfgQZVOMm5C5hCvo+f6PX+
yDhsuKJy4S7u9gvlGNBu29efQvV6OZD492Fco7yoQK2wBgpoPHD6zxyV3QM1X2pB
TkJ9bRVa2lm3CPQgO7+x+ScTDcHAxSjbzXDC+TFzTmb/dEuF4OBm2vywIcOPdMMu
aRyJ+k8xBMOuH3rlu2KabaZ3WCKCOl/tYj4J2v8kQu7p8b8UfTfSWWH6/W1qIsFc
kgmZQ/Od0YVbXQB55li20mSzYXTwhtP6wv6bTAQTNHQO7fzQYkDODMeaw/H9S6nW
+Yowhx9QZyYmYOqEWJ0NLJlthoNRKesqkHa+a1Tx6dmmpJGuJ7jW43uI7Z36Eyu0
D6dTKmCuphn+yXNTb6cEjskG6ry4FurOAyUKGputBeT25EDm+EdLt8XuAWHOvSRj
xY18oAnz1S5fsnwwmxyqU8j6J6FPq8xJvxAm838A8bhcMkPXjElFZTrlO7si8hxk
mN3IJjlfEKD7s1QxUV8MYs+Hem5aWTDtPBX6UGk6ffbTyblsJ3uoTdj7/CK/eMBe
yQUJHfciRv2wgOZqF3x7x34pWy2ISKtDlPsrcOy+1XuSgrFk+2+T0LzaQc+8G6PR
snI74PuewKP0JXEyvwhr5PO0OW+OnqEwVzOOMS3Zz/r2qgIq0UdLJUs2pHjbitZV
QMhFXBgRtKhvu7r+rUlKLuzXPLvyl/vu/Eu7R+hfjYE7ZSpdT1kb+1W+bV+benGe
FdB0lhc+iFq91DSdrTw/7ox+IUEiYWZx+lgz27IjDkkcuEYa2MEzGCQmVUGM5Fbd
8Jt9skbzecAUMikRNyn2POYAeR/GM78n7jbtD2FA7s8vni2nfjPBmRvA35tUdJuu
NuYPTmAclE+2qI4lORN9GnG+xnSPvPPdAfd9Ft5iYfbRcDzE/SB0k7okSg2RitBB
ICekgvNaGBsqsHoDP63Q4NNuxvjInHwJrn4AUiVNnWp1obgv8K6OOcgsY8J9O8+N
Iq5Kel4kFcIwHN8YvjOMton8k7IaEbUo6FfNWhYCmiI2JqWOTSCfHmDgI79BIq/o
j6lc0T4Z0J7WDznCExatJydFXyp4JeAtiKAqMG3c4/LHMBsU9zkaE8dzMJtQqEp4
PSea6UZVpYVboeQwVeI5IlLTr98wUqlXQfxTbvJBCL9F+riW2j8DyhkXiQyKkoho
/ZU4TvkNh9syAt5VrrxWjR6YcpeAbk8XR/NgkfAmdeWCaJZb5R7/V7cLk8rlU8Yo
ruGmeXCEAX7RNtcyAEV8OjJAGBmyNu4gtLKl5sZS38uIhvnCmi/jZqfIaTDxQhmp
K4LcctdZfdRCnopmT6+Littvd2IiWtaYxnMQz2PkN3/jeMyWiW+og2s9tN+szwha
3o1liEAc1EiRwDjXr0fmfBp4+MPopAbph6liWb7KICiR+UoPjx2jHyoAVHa64csc
ebmv0XlXrwuqFU9gfn87Y443OwS8xmZhaDJchAmiaecedid46ERjsacjXiO2M0A/
kyIWBECI9njRw8zJFUqC9pPQRR4KqJ/K/ufuIdySv7wRsOZ4AeXx8cBtduQ5DYdl
FV/si+el2fIZjcQGjmhQ1alIoe4XexsXtbRVQ1XCKp0cSYSVDdoH7jn0ECsIVtvb
NmZad4GWsYAnOQBxrw/025V9gv6XQHj9VP4UJOQGgI0JQpI/LcJRQkdxyGtZ0ieu
tHiVuXG235yo65XabXL4jjAB+z3vHHAcZoSY1C/sNvxaYeZi1/3uxw2FKRTnikjT
POv+ybU9ecEPFueq1HZyOXRCYmzMLJWabOu9Tvz0Wbo5tDRh8Mh72elYcw27VGXo
7uV5ZX7sSvQQn6cNVo78laGDFS/PJRzuvniIH21R+DQFt9UotgGW9dyp+bKrraKe
vl9X1qwHConTT1tMjzL9S74DWsn2DGZFy0fKz/s9aYEmHS3twbPITXV2W4p7tuc5
ZZoBBcKxwLIWTomzhTWvMA0upHQIQ1tNrMRzBNqXnxFNC64wcT//4Ng4FIs/Q0Cd
lxVkboQijDunk95+Ltvf2Rvvo2oKrdOdcRkfW7F27gYZQME6dJ/QezlIxyO1baW+
RUJ5jLj3zK/aoJrfBsi/m+C1/X07hEzi6hgmEuaRF+eADE8nQ/jtUzorh8ctPn+s
Gzkysr5pIMWOqn2p7lgSakwy3VO1JWAaEG0M7A2+Zus7QPVM1acpvUY+uypmNbI8
f9FzgiamyvJzIDwj6lT+/EB2PIHlRaXLfJGBKakj0+uyx42qBX2mMbEHYY7opcYl
+8XzyY3DhHngKZaZOmGwtCN4hHVlh0+zYL6X6JD+Cn60KM22NIqUG+d7FYYByFy9
pYENNwOhLHy5kiWQUqsBrFYNVcLc4hi8Pej1+XIafgXK4KAXTWdgo6w0tDVEEL7P
o2UwKdLuRiAPY/l3xWhmpzq3u706L5uL7BGY8XkOXgYiL26AmIXRny2mHY0RsNhO
I1DgvMO1Lsbyq2NX3h8qesFj8ZSGNuLT/kYsSQ8UN88L2t9zQ6ngQIMMbRutChZ3
zTGITfYQbFYtVzCgrs2ZhFMqrbWyKZgZFjJO4e8zpI9tDEQfly/L0utkPC6P/v8h
+ykfqrB6zARna0ZT5jCSry0/rGGIprNxGG4KmdyyDB23cbDX1wg7Gf4GqAlYqo7a
yxZhc5uQ8xNBN+kADT4+gVoS9Z6Jbl3TgevY4I8BqIb3hZD0rBae1FFkQOfjLxzm
6Qyh1zU1rr1ml8lDsTof6V2GY8sK9PmX6V6Vw0NFnxKbdAwlRuH7jhnfx6xZ3VsA
ZpBmC0aglVa3Mn2tHggWl2p8RjeKcfnY+qJHFOCPSn2Vag0qJvr9F+4L4kqsqrH8
rSmLS6W362VStODlTUDKClIzwF5L0bLBWk1LYAjV6IqqksEMSrn3Pq08ZojMnphW
nRGK50j0wkfEvvH3Kg77EpOJgwzlhoGOr/tkdEHR2yel/hy3dCfAIJINRC6v2705
fyqja/YI4ReQSrNkQZw9wIKWgyL5f0CHQRDFCiix5hIf+8xOFAHGEejBcyXr7AY5
l+A0hkHYdIrHITQY0Ljpvn4NGtg0CFB5YVtCMtAD8ch8h6NZbFRY1fAxsnV7pkmn
GPRj12SnMnJ6aws55tfGe4aagBWFLvwYcX9A0cJdvicnAf69Hh6BEl4DluEqHS7q
B18oY1ftoAr0cN2p5tzKWmwyg4B9qXR+iHmR0AkHSYXbVEES+Hqv9dyv87iL+mST
wwdZEQ0+5xlxuQiUAK5Kl+x7XTOTVgOb89vWVS800tz5dZSqM6agAIatFbhLw/Fg
CzqffwVxIpnfaFTesHKUpsqFYXE3tE49QqfMORJsCTC6f1LxR4AxCD6R7TccmPr0
LSEqTmhoRbELnTV1TMRAHKBpnWBbrQSZx7X588NbtOD4cM4cDSJKd4JIp5YSJm4m
UDKT9srsHC8FIPcA5Htv6qnuLSXKAn84BijGI5D35Pc+EgjStnMHh1LjaucVLdEf
fjayI/MzYabNHxurtene6RIEdqzDylZBMbo5B3feOBa+IGEFU1mPNr9WA+2hG/kA
UbTHEa3vEZ3DQn92dgscoiU//BcDysf3Qx/0SB+P3MhBrkWV3wJlxv8zZ2i9Syrw
hIH9HDJgR5d6/HslCJ3FDVdrvTLnHZ2pfLLO2VTf+Gae3WLkU6r+hIh/WJEUxJLC
7htI8XNl9XUTRy4xHUYKck6tyACpdan/5JcgD7hqBI51hjwOcO2JzUX9ttjSAp46
y9DAxHCAwi9iJ8XbnIyCW4rdEXcg+n5nA1Gykp/zhUAoY1773UincuADeOGcP65V
2MUHGRbuylYwGJZ0ci6ahkHkQ7Ejf7/+YDTcPDRHXiJV6rzn9wup1EfhNhm83N+5
sXSjoLfUbFzgFz8Cm2wHjnXRBhqIebI+/DOKQNHMxPKjm96ITTRAhh+DJvuZLu10
Y81tyU0tnkCJyqvtHdQ7a++YdjfmLT0eid9aeEM4uz7EQB82Yy79MXD6JLLShRHm
zaar/BGkWVb3m3ul8NPAwbrvD6W6lN5xg4RuWAP9VjdY8mbc1fJj5D9bYixm+Qsl
cP0H1XwK+AXzJICw0Y1Jif6HZcx0JP4zBKyohb6v2oxTzTiWP8SiIVaLrbW/wLOB
geazofhbipZyj4Q6WxV7EtbOho5iwFp0mlXkILww99HxqTZLBi6FrgxpmBr6HZju
P9bhkyk66SvgeZcR2AVRDt4DBrzHJ/MNWvnmlUvm0aFynz0U9T92/fjz/gPmyITD
yzqBuBIxlxjU8LVuGxcvTf7xP1duhVfZ93p9sh28w5013nQIaD9eXYL8opfZPfNf
sEfY3AyICplpQZtBZsH+IfnsoIEuknk8VU1mZj7H7gevxRVWDTPSgFEzvllUs2w1
dysByiCGGu5ZCkCNVWR9fIhNtQwDkbsOnIuykoFCKNI4S1xy/lt1tCmWInLxbibw
8/Ya/F8vtrpbxUWBnNOusTa3fmEqAMuTz5svPrkFM7nq5GwGpvuiD5GpbnyI8jO9
GhlIaoVhqaSKcTMAEAWf/bbCLRIGAowmzLj6r7tONuNLsYApXD4gelVAH1aW2w6u
PgdRCnTwgw6dajECf5+NhI+tGdTHLIDCXVxG02jRxUh6HHFLqAw9hBnVm6OymOW6
6Wuw613XNND+eOlIXWF4BJGqzgDyRBP6FyIi8cF7jAj0+KqUvROJevR4oO7ZUD+H
ZBxzRfUsggu7oL3zgJthfUVW5VG2epiljpHAbFilLaV+ZsU2WHR3FHn7D/42nCD5
4sz8npzNlNTpMpOQkZUfF9JYVVPJmdJgNtQtGH1/gC2x2tfWk/P2bXSSVOAIDtec
fRdwT67PsjhX8MGX7kAMKEbEz3eydnpDZcWOB4ERSV8Oh67lMxICgs3yJ9cHPHro
QNipR+QFsVBFZJaDK8yUoBCnslAbFEypjA0G1YtwR2xHWFJ35IVrrIgML11+zbhs
OFjTEy4Oexs36tVhQzVc67FXKDN+bh4x4Q/eCJisYqkKiw/m4p9z2b1EKMTLIewq
STe4WT6EIKbWE+uYALv7oDdJuIUM3i5E2Jt8fqCa5Cajs2s6vzZ00moy2DAbYPO1
vJ2I+0Tw5Oj5AhT+CHw58/eFrnLkTiFA7mnZXDACtEef1ILYUXFXmu5Jq06ruq3Y
XWXxDAPKsGOe6z2RJzsIVPUO8NZlGI0KG5MZVmMoyQxSP3cCl62rZlDq88YhxTtn
6Nh1R2dyiBAaoe1PI1ldBjgj4kaf/wdW8SzVf9NhACxN4BjkauWYA/7XqWudcKuy
0AyYiBauJfpv5xgS2mW/gjdKeqG1BO99E1I2tRaszSu2H0jSIZ9wqDcCKq9H5gjR
p7zCZHIfBHbCBq+xxtQ3g3lZrSilZA+7VtbhmeglfVknzWd4ejauzB7dCQuqosBm
IlO4OHj+GAGwPMcBKG385aFtApz9YAbyfF4tfEFo65itfV/eARO3euvuwqnGbC/K
G4ylbMjXXxfH68hVxfbIx6tJ1jybK1ggaImapciVqFIkJUP7MUw30TV5ii5ba5LN
SWWcjBCdcCl1I2E2dpXT8iWBl0vsTEzIVsJRDcnpiSq+UbaJHEo7FXW32p5/8gSL
M7rmnCYzDdKZ/+876V8uvpEISqm+atffSDYxHhUN03EJLynYFb1NwCA+6WJQgcTa
s81+xWDgeOhmwT0QAD/8Xwvv8HDANfCQfEuvHC11Hx+LE70j+5rQyq7AWsfAW74M
12fnOFnRGfzxjh8R8wneNnqklw+eYDhPvOnddk73hB4lPDcvskEJGhxvAVEvpT7S
sLxKFgeUnrZeSoWOsIdfGEIr34BSO7YLh1B7NeD5F+ff3WECo2QlHk6k/ugmRZ2x
ympTCFCC7aKCY43Gign0/iuwLjwmPuTbErExS9PD1StjfzkEC3wE6qZ78+AMHFcZ
J+nxbFm6RimH4NGm1b8turtNdcuznti0iQxb9pm6XOuVN04NmonFiO4JfM9Uzil7
PPUsh6Si/3etZ6zUPWrqKsjlleEuUCXwy8+x+E0TM6slK7EOjwB6762EdcThPBWi
xjrV8M8SpTYXy6zidjn9HFaB5m9qYhYM3mZ5V3hrwPXCRFaPGv6MZS2Yog2cHsUJ
kqXaO60cbJhsyb2DUUlQTJo2O0+y3hMVyPKT7SohRqA0ngbBOPf2//uqTLr5cXGu
p+AXxFe2ICHAkEMiGL/t8QUBXMKuDvS2F+X2ruJaTf8s+UDSnUFbNL5RaO4Ea16z
55GhT1WQJLKaUCMiqQzzEUOmiCfwJjGCcJd4H8d1BAvtVHW+Wt9tr+S3I+UUDlJN
hPzceKlhjlvvSt/xKqiYYcuYv7QCv5Qh94hKMFLDpgl7Ktes9zN2xHlrerJf/C1x
HTaQRJ6mWQMGJYTXks6KptcLgLmZhz7ydzkUntN16XryLFxoNAGRK/d2XnXPmTcA
g5mEtaLU7UxS2hwcvcrfZy0Lv4Q7s+Q3QR/Z52+F+ydj1mCZVeM8eL4FrrNQEOdy
Cdw80ZBtCJZ/0OsjrhQTRRl5zyAeioqEG5sBAftoOlQuYOKH1lJYrJYFHCH19bYk
BsR1YaGWKMmCV2f7A1F5FdippekrW/71sTObNl0eNbr/NiC2l0kcTDuHz5tuhs/L
lXBiAZOx7spcQVgqAtpQjDE4CcGdY4IuzkMg2CIe2eJHQRJU87xfWTn5vjb/WlT8
Li90796ZRweLpy7nVva6BqlzALTWxluQSfLf4rEK5L59fe1XU8LmULBCh8Qg7oFu
C/G7P06DNxZziNhqE1sCHprOavJzoSr3et4FBvQq75/1opMQl/Bia2SKF1dbs6aM
Kpiq/ul286BQAQBRnfJDO+o7FjEsaOr5eCH6l10WHnkzR4cxiN3e3WViPpgjrwE/
WtJpQ++0fVPsqnlLpi9JPSkWLa7u1Bpb23xMdgPhNbB6ZP9WE2H4CreGCbVYqkN6
2Wk55z5dAUWhVb/dRwcQrLLoHarl2zWgh0J9hiYsHh40FPeqWY4R9pzNF70abB2/
sprVMybani6IJ1MKB33UIeewysX9UT4ra7Ifu6DONLAbuY6tUaWSkY2EDpq9oDap
QR2nUaOyRJy/AXBF6p5qYyQs5kpSM07pdOhvHTlJEwsBl6Z9svWQj5esrKRzLtWi
VOIiQCOSfjr/qOIeq5JEyLwYjAz7Obdz4Anml9i/E8z4n1LQO0w0URRQJQj4+ks2
Yq1vlnH0Us/DO9U+IOzenA49gREnME5tabF/pxbu4zeF7LLtEg9VSRCzyQk7p8rm
EmqGQiDVboc9H+50hvvoirlZImLWp1k4zqdxyaMXgkn6nu9B3EgJaQWLQib2ItZa
2+9XF+XKjSyPDK979/74g44/lnFQ8iSvMrmOt2kEz3s/O91Hk6Dy8z+AcQOdbFki
YPK8etUQWJmWDtPlG4jYIUyj6ooKUGdqLqtKP6VUsBHsXcLUSwXdExgjdqfqN/qQ
jUHlZjMV1QIXBsKcPn+/1EY6WnFEQ9Wz8DQZBveW8n+mORJuetvVVTcI4tziQYq7
/EwIHO2LzPmhRuj5nPu0RA+5bca1sTg7bLkvEanuEURztQssVmDsJLjwejDKH81f
bymRLBteOiWHtXpeNXmZLQaFFUtpuGkSztIlp1bLqNveNpypkiGaaJ7khdRFMi54
/ZnY0ITst3qo9tEs1T9y9oJRvT0DLNG1BNC9g0LpFEotHglH5SognaLx3KYbg8tp
/6CHB0NGiY+U59inkkWefFfhQNqM59S0r8gh92blJouSoDOvOZGBh1cu98q+D3Sy
TWNzx6EigfuVJ4CFIm829QTlmB9S0FtmBKx+QuNPDGFMh3T73B2BOt4b6lPX1G7d
HcxavJzPVA3AEiBk33ksOWehHQVhFUmKlweI9RBfGaeL8qp4GU8n+nrLCMZw4KCp
VpLLUGBR3MR0SPVuDHJMT6KISCMpdMDoXhtK/CnBxbmZREbnd9GKcRMTK35PSvgk
qAb/3wpVzQtuYyrDtQCsZPc6TjQJ/r8seyvWoPQtXygHRbwq7TWqyrLPOyDsCxe0
O1LZS5Mt9fIAcXgIGNQo0Gce4uyUzoMV/UdSQHXtYPHGsAewJ237eM2db6gOYDm/
6STcHeiE35v4aeSMygOXXtulDFWmscV/5wRkxbJmAlxoPul1iZelC/Bggc2ZtvX3
mIKGcd+H4Cfp/t9eTw+2xvrNti7dDFIFZ0wXTlrWwrcPHs1EwdRZIVBoLXcaLUA9
d+JNZG6fo9sqjz7mXuXHEUov+vkt1U1QUzvchZPyakqQzGMS2RljuaZmpT1pDe5v
HM+AGqukEP2hbm9+1tvtWwPrjbpmWgCJ3eCkNjGeQ7Z3B25G/ALlBn8b8lWGhEsc
bDEgX3VUTaMis62B1nDIWJmKgHcWbg/3WoVasfMlb5/c9WI5gU5ig27DO539j7Gz
M5iXbUn9eCz4Pd4Cf7lVphoQZX6wLq+9dB/oXGRYeUukeX6Wajt/GKZ65VGgSnb+
IqET3fmgOjzcehTigyNVhD3+/4W4//b4qKGDP+AmAe3LyC9BXS3/3RcRdF9Y6qwR
MvUEQGgrMwZt+LLMf3OoxWaTJUjBuEsgsVggFnHtG+ytwIiSsCWDTFaz7Unz/Ak0
U2ji5yUEw9dTB7T7v1bnAsL8qAXx65aSTuVq0LpZlcGZmmdFUJZCmLTA54mCoqff
8Q+NGXoqBwHkh+Se9QHogTs1+orjGMktsqQPkqYF3+3gCNXt4Nc81rIP2sjA3E4T
4XaaR8CUw1+I2xkXnhuDy35q01/puLtGld2xYjRMeTzrani1rSPAfQdxFJlcF4BL
2Xk4PCMeobz0xnHEc6Q7l7QP3KLWx7f++gPTQWq0dst9XPUIy6BG7Z7yCeXe0ILm
sBl+RnwJuiq8OYAw7kf60heNZr7wW3CEq74deVfC6tQXG+65rJPWPyfzr7DAchcM
xt7FANVz/lfeYasVmyev56OXdWBC5TE54PYbVVLphJLjiS6PXo/v+vRVcbc0x/Oa
xRb4cLT4vkmrf16W4shZRq5+LV2O9JJQTooY+F9/WHdiAw+b8LgEOR8MfE073XK+
t+I2YeGCbDdAobcp7cxS5E0X/l1/7zA3O4CFLEn96yvYEdkcbL8efkfQwyN6twUW
dOs4rvXlfCHuSW7U3PKgzqOt+BFY9dltk+/uMnGH3volKeLl7IGVvA+PiFLpkXDX
GjkgDmUAL+DN2MmdO6C4tRZeLxAZnsYZIJ2RJtgN7tDU5JM4jSJtAfApHDJuvQlj
5SRpM8r4WYNgDuaatdYaNN8SHc7qDLKFfD5N3opIT9uwhxEy0tgPFlF2AUnuOw+E
OZC/CxgKaWEMAf2FQ3vkaZU/p6pPQRIoJl9BVPYci0uA40NA6QeLwpq2V+VvXVN+
6Lfo9sNZCmUKx8HCdO+Zn2u2MQh3UkFuf7Ojgz5J1ERXbPSnKLwpWSEi4p9s0ODu
NeijVWXeKg0cRVY5oUYd7Igu0e/PVPW7a3IYQU2d25+iZINvDsMTRG8+XsayYb1f
htY7ILBSPlcX/tNQv2q+gBZQyhmkBbMj+Wxc7zQbZIkXw4WPlevtxtmHpnc8Hcrs
XmsmvtzaleWnILETKnsZLjG/TznCSmJfMZGgUUTl1nLEU1mQeMpJAOLGWOWwwOFl
pacCe9V50HiU8zTFAZ9fbFWo9ojQwzpZwp/dB0WtQtBVhXucjtBVz+MA1BIME3bO
AHCUZVsfj3s7mQBdnYgYYPyhLe/o92Uv9emgX5gnvmtCGjeI/3vk1Qc4rrJNbV47
ZE9wa5ep9OPJ9ChsMlQxTgT7ljM5QZyr8gQvrgP2S9kgx5XDg2KdIvp5UQmmJ1a3
aPM5TdDd2FBmYO6rOzgJWjtnBHAEiKMp3SbAmlybTQP/17iCdEgQM75AsY2CyT2W
nyg4lGSNfmP9JwNzxijfgtCkXZVRE0ElxUW7W6KAJ4e7pBuCj31aYFqPu2Zre82t
B1Ei7ntkEZ7Nzc2obMbE3pWmA0cR9S2e2yibWw1jpMNK4/eY3A4WG7drO3BsJtI5
CdAY5N15w2MFvlrNvvRtEkirPWcVvEDaHHFa7G3hu5UuibJEFPXE8K046o7xr65p
SoLPtNBKWmH8GF1dgijtmzCxgapC5jMY4/SI1u7SUC7FXW3VBNCjt6/sLXij2MY7
jgWgt9rQDAx++NvNIoaPlouw8MEtIxa12KWQMPdv80ZFxNa64SSxyiikKAw/ALD7
PqTbTaB7Uq0xZvk3+y+h4XupRwP9/fxoIfzGPgyXNIE9/o6tPxmYjKl0oh+Hu3F8
OOsMb1HAjp9sEpHLy8mZUtuQ794I4dEfFAHIiVi1oUa5QKLdW/FHo6ifTn5W+W1M
eLQLw8PLFmjL/PWKV77HTixJmczoybC2fB7tAH8BtW/yUTmpSOlu0ww+5mCjINoQ
0d2HrA1W7sUnLJN2Ky/4WLAgEdrJYIyq8Ub7BXME17Y0KGRqyxdaiCXSv/filIMH
nfEm6Lz6ptBgr/WOd9JvTx44ViHLIP2ADUp+8+D6/DrLJACrB0amUwlz2b9xA0NP
mo2tLOo018LQd1Koo3JmxlwEM9BKzXTPdFp8okNwFfDqfjHCjX65jsjEBxFyFlnL
SVSYkSkrltstQAHbnedoWSjDQDQkW76tTT4YuMya/OfZFTypDisf4MsO7EfA8YsZ
xMTZLIE2G9WYFJG5orwnjIbVTIPmavwA5Ntm37DCPgbhS5TxKQSbJ0ivUe6tOLT8
pyiKC3/8HNslRarTDV20f8wnu3MML8A3zEBe2ykcBEk+6p+Tmr/0JTGA/8jUnfkY
fgoqm6bnnJ7hmYtlEsakwCX6E6+/plslljkOwyt2jq6JfEyqxOQgRGlCw90hJjUR
slfQRzuA3e4t5O4UWnbVd31tTx8Yy8TDqGVD2nmRuYUB0b55cyFizSSqEphZLSit
bPpmKV6VZg8VDUjBzUsfe0TC474hIhVNKcWiF650IOFi6CbLjz98x1b1axKbmg4v
YhDNgAxNkUXBDlWdmq+wmYPhV66UR0+HrWrnV3JHUe3ZRS6o9VxBc59uho00BEjU
7hcY1amjRT4147Buu7WQZuygauNyHHSOLjaxCxffDlhKNX4ThAe1k6aqPT6OTL8D
UHthJPoHPSdLBTjvkYj7LHrQ/nMyH+Sp6mqs1uws/NsedfDcfe8es8m6H0/LqW9s
CEH319Z9K2R6+snhQa/QuaS/CjH97ETYjbfVUX3wgHT5cAsGFh97ZUmwfObcV0XQ
kV3/gEnOTfWngnNTxEnYL2x3d4GRAxgpveh8H3u5YbCq01YhF4KoK/9B3iJk+8ZS
SKsMF2yl6DUxH3fWUh/E+HcpGd7wXUOst+RMG6FutZ2MD9I5WD/Othwu2W84On1f
udrwdXvAv5XwfBBbZfTjuMpnZCjI7g1NeClhntfvb2vlNm1OuB44v+WVsgwT5Sou
iLAYcRaEI49XxQILdInp7CpO0T9Iv3tk1eA+fPRndVNj1O2b5r7MsRxTJnyuGvLa
hMi5cHHKTTkym7JUX2f63XDoHRxtjlmpwFut3eDWKdEUu6IPJw52M4joR+EBtv56
heJgYF2HgB5gvE/h0BZZsLdHZuC7A8WT2pvZ2uOna3nqik5JAEDvLTueN7wLwHyn
ZmA82REHrNtUyKFtKIdYQv/7qd1OXxGw4Clra9gDCFg60FmrwNkkPVyP6qArKFXo
mxFEtHQOivlH8bSF5Wc744rWduJwjYqYFnsZy2V3wXTqN/W1sGNqM8GcEh0B/tEy
2EpJM4/AmyJcxNXeEHsUDq7DhkJ4q1ndfMAEU9Az99IvaHDqmqSh2pmHz7JC6AUU
/spV2PEETJAFOKEIO0tzKyFNBZUYS5OdazUOH5/vCoee14hk1vFXrws+ILjX124+
p+EtO8ZEV6Y5mX2t1gBotefwMHble0VQJzA24dQfzyDfykBPOOTXkk00GzweaVnW
pQLBqoBp+b3Qlz3l+Zrf0jew2Ms/kdRkZOmVNyE2Ka6s7OUg+Ge9IgPdiiBqdgxH
rq/Lx7bMllAkMvRyv28BreYqhlHlE06+/fdQUIMHP8y26wmln4JNZIdnqixfE5Bh
V1Rs6M2UsmeCEyI/d5xA59WQQZuPkntPecM7V6peR+H5rfXPrKpLqLznmMQHyCQ+
DP5NpJxTAbPc+cxI/10SSlSiUfxWQGacn5sEnuzCiT5GDSVoiWrq3062EyDoL2aB
jf3c24nX57HlyT0IzXEG4XvpxK03ma1qigTlPtT411IUT4FAje3+wNsYXMlS7VMY
peV1sns04uRyQ9FuPKmUbRr4G8Wk623P6FiH5PUqff5QQ/NXSnbJYmRK+IpgkE6k
bHe7t1FAtdsJoXPGNQQt/QJTXh9xDmaurrP/4jkHnzPXjMfDdT1FkYUWBt5kBGVE
vJtBcj7gfXXx/haxDs6dWmDrCCOnyY4zHeCPliI8EVryv0oNKLaeTuq8r+KYnTbE
OX9tNSINZyVHNEXdrW3AZNHS8T9yiJxTfhWAQIopHQOql95X3Ooc9ERzYebgJGJW
sV0o0xAKQEAkYdUnm/MV59CYuy+M3wtyJu5RzxoJs6hT+oPmJt8xGbn0hu0VlSw4
8GR/n/ne9E8vyUy8rmymNutjLch/PEhDjrpDmG+wLe22+Y2Os48Y4PQkg/GIOdzi
LbsMgkzD4GZc2aXgSn+trL0LkgSTd089BdBnJW+2Tbz/Wv/oiQz0hPYFEKh9nyAB
RPHGtc8ZcFvouu3q+Q5Z9vrsErtanT69QlQEPJPZML2nao3T2c8McMz3Tq29dlPU
d4e7nX6vyuvGbA5vnDxH7XQromUpaJhC+yv+VTDt4Z1kFexCpjWkiNMhGSU20Klw
IHihHbE0Wi0yfGiZewt7HgxNGebcz08WKeLykYtnl6X3JsfxLMR6obgvZCKNxS7q
grc7ZUvnA80AygSNZ8cpZf/9oZggFpTgvbL6mFxJQWLD87TGiCXpNALlL93fuJ5k
AgsPH+y3Xfi3gXsyBjliwUIMuF7aEF7FDwfc+MWQs8S2PtHdO7u1pW33gA4WR7RL
SRMtAIlZgRFy7gs6hUpU6EM+1vIa83195DNRPQQn/fvs+mKtaj/84vOBPOTXT5pE
iCwOfTn2wL8f5BzaJvmSlfdRahu0iZAbGaE8M9KPPaLmX115rHbZSPw7ZygfILAC
bI+MxQNfdaX/2NomhV1Zx7ey43hgduH18l+6tXtyjK4d1IaRGrYWQkZy5EoEiCb5
/3P+S5O7YboLNfjYZzWkxIteqFsDr1/dJxVaERJRS9yNQ/piwHrY0YnWYn74A7kI
oyux7Z2yj3pxjITo1KblZdJklkvvO5DM7U+2CCsZD2SEqh5dRi6HLC7uxwMFNeRW
h0GMyOlzPC0l4QLfkJf719LEmSBG3ccb6TwueKYwmyJBpMBjVPCHBbG8H3sfGPrG
E/4LCZyFPWwwMnYDQDwoJVpJwuDa9SsOzzUBWHPWJ5lop9mxxddgW8Vd2js1Xr5l
W7pT9bbPV0u8VaOfbpYCtglad2Uoz1B3upyEjh6pC0rfwQY42VDkMQQVEedenBnG
EpANfS+qTf9s52LqTSkxLtYlFg+OgDXgCoUilIiU2ASMtrBviFid2uPwaL8h+fHI
9FpAL3uHg2cGfg5r1NkqEmgwLzfjUdZ0tdgtDZPoLluwnXEA6kqtYescd3z2SQDC
+a3/W4bksUGle+AAL0C8UqH+jn4oajkQqNH3pRFmJiThpOJWNyuvpLclxCQfedVD
jWh9EH1LNEvKPr5KlYCKJ14D2BnKzowi/pRjfUZuA/9jfhu5qarJ3A8L+E4ZfO+v
OLxe7bqbc1xOfs7Z5LKuc+En+r0k1WHNIreBxoaATOPD4x1aFtcpVWyQJ8yM+6Pi
sGncoZwn28cfY+TDOBfgy28WLVMmeidIW8J+z6i3QwPRxG5yJpubigMyfUoOXC+b
8Teo8f00uyd6eKugvKTogIoPEP8fNlDGBl+GXo5G924IQ07V0LuS97ox+ifYXh1K
29XHAZ8V4nKaMJ3RFetu7banjfOBN9Sf59NOaVA7l62Hag0FCU0+Ib5o7S9bh3jp
rN4pVrzs/u7Dc7kWpJM5QuK+CHpSR083a5vAI9PZkz2PM0VMMj8p1MVQbjMKmHvI
z5Hb+lsgtlJBroRIenfQUIl6J4v155lHpZ/tHzDuweNYFa0D+LNADgZt+rKPMWfT
xCJPJtucu3Lnqu4CjwxGFd6XLtAd+ucUabycZ1BkAQBGb8eiILx0VvRa+25lbiRN
V3Z3vHyEoVZY3vp5iC1cPl4L24fc/lRuHS6ZU4aIsiJkdmI+nuifiUDnxYGhgNPa
hA9Rg8SaLLCVUSBkFqQjTcwJsMblVZm98tofn+Uu5OUKzEP+GUeF4pmvKdJUTi5C
EJZtQ5QE8La5C2n2RqwCQCeYVkkMSruqddoeMc0bWwzE8ZaxGXUQYRheP1P7dQC7
k6syhyWuv9oc/c5dDw7tPVF1pIma8C7UN6EJNfzrtNS+ywXOZv5QeAXKgZTDlhkU
V2lZs0apgkFeWaDSzTv9XDWct2CDpbmYCIXSdPYLQXWsdtzygca25Dmz5x6KSsTX
hX4U2LmBNzFRIuozJIdfF1ygjKntKP7O6D+dJ1aIqb3+DPNGiiuvSb0zz2x2OgLx
vdRU4mtpussJxAqYO4mX9lhmEW2Y9uFlVbTovJzEIohJIvTMrPoKFtjKWPm/xxma
/iWIRXf5vP2S5iDf4B5lUAuO342rORBLndB9VMD0XU3VNLimpfVig2RRspqTI4gZ
mILWi2pFE9nj5JLTzdNNnHcFIrwICQNa2+gb80zm03svHSkY/BZkqwF/a6CUdQNw
kSwaUYaX0yrXzsVncMwZnhl8wvDDFLRvkdhzte8Pm746/O4hZCCLlzDzSiXEvVSB
2OUH2CXXEinfXVk4XUeJm5wi1EChUaVS2OKPDFHmTopBgE6x30a6cf4W/RcQReln
zudfOioqyoi75V0saPi5qBdhXbdHtakH+mowdbJvTfnmHom27chLZlbz56BwwOMD
m78LNYtEl1/iEqZQkDsXYVwm1N7nmme4HR2AE02mzK+FOzWjCATt9Q7DnJlIi0f3
7tV9VWaPlxeWGJ8Urltng/YR0508P2K23VzwI+XTiw0lfgNoJotbXtwbuwDtUkoK
Jm0NBT+HjDFMyYcrP+NW2AZ6vi/th3Mp2oFWVm29RK7Q9/B2AdRg2twBUzTvu04q
iP/A6ShZR3lpBsPA4eEOOnOvyxDIV8My69xxNeAIHAvz/4tsRvYBHCUg6B8PUFnR
b+z9yLqVB27FlBTebYyDLpqbTawNlqmxQmz4Qu8PDdNGQA+QntnDeo3Fii/RdsDi
aCbfGryu66XWXt57MUumYCuH7ZZ8Lpo75RDsJRYhF0vYrjaad1M1/Fas3QPC4b8Q
MO2Vdboa/DMlJdgExOaMEzkksalaiLrMb2qwEdVjILrPwz8AuG9Zbx6f3jCz6OdR
GON23gIDvoWMDstiAw687iCFFXQT4vt5/Mdh43g3sjF6YuQR2akMJw+amKMIiiKH
BFkqhDjH+z4Ny01YdIWscWcn3XkpJk10EZ0i2mBVWC8mEmNYfzHZ/2954hnoaA3M
9aB/FFtdCrlMKP01ZxYOd1d9QWPVbVmbbp9kOWMG6TFa7cj97bLt9JTqXHSzFXZI
+VRIXIQB17fX1FYF8dBRs/N6rdJFaBQ2geh0cJKORXMbiZizmmUglO9TQZUz9poO
qX1XG/Oyv9TPriEcRk4LqGlRkuYZJ2pzhWqZSCzGQg+ZJAKpLeWZL2Dx+G3MHihC
SUD1uTseeo6ytPujpj5fwGDpjEIMsK6eypf8ms4EPp9Iu/D21xJ79EfIr459eSxj
P+kYB7SHZGkEHmS1ExqTL4ys0gyyv+cmy35QTwY2zrJMXkIbIxrY2bQpKNYISchQ
nSPo8Scws4MpdRKIKj9EL5fCB+YJNzT+IJCqa24eoYL6BWa3+W46QJWUPdH/nJGE
TdBysQRO34Q/MGkAnCeEOeFx7ikS0kDNzY7oOGqH63AKsviqHWYb/CrXuWFfTMAe
jpiY7JKdn8B2Y23vQoTLiUunhWajpB2MAtXFjFSi0DmyNZreInnymzweZIldQ6Ud
zDVUt3CObrLl4Ho2Vu+jxMAr13lNDZn1tuUmttutjQdYAIsWO6OdB8+1L1fQbm7w
N62vOqsRJEztjJ5oGtJXMIxdx7cH+1hi+aOQgdiv5G8zd9Z1BxM+E+vx4bDhImhw
EFHx9DwSgymhyEVcimnQsUszeCDXyS6f61el/aIeAyuSlkCHPlMkz99cxahrjsim
Ix43xJkTHp99p6tx5udd97RQVLQXObhKwzZ6M/zG5JWjEq3UFyh4Vth0v36K7u1D
Pw/zHAoXW7vfPrK6QeQGtGhs3XJ4CBNr/0601NqUorkkb9ERAZzefMdEpZ33zcCu
XK9rOIGkzNgx7BazbvZd3S9QV3J0+2Y2BB2wkX2PJi62j8hxutOPaDaB2F1ymZjn
Hwuy99+6MZLbY3yD8KWeArz+t0/86KpkvQjnQh1sU7XomrO9iJghQVIREhh9F8u5
YCxCzYIIzvmw3/cz3czcAzxl/rCjkgZYWiYGUjlaQWG/g12cXSzNlwzylfssxURd
WcFMTyY6otrjry5lFFAeBtq0tuAQJ2dLSzp/MWhHbt9uY0nIfou1qCP+Qf0FFQcQ
m9NBaqfzSyAoNP72MxowLr9IFJ2W5JXB3gemyJDAfC9hmvhpvIrK9IXJ3Muezml+
tw5MvbsfloiuAVtXhH10mQSkgzgNyGoetbPz+o5Lv8nAyl7rxcxWjyzB8nvUyX7P
5xx3WMiE90ARErK6m3/ax+WT9hbh9uOfIw3qYRQCd+j5TM4s3VLeks14cLBTkF1Z
XK+XSfObBBp+uyUT6nvod25YOU5h5yw+YZv47RD9NQ1J9t5qNuUsNWCE7rrjPPd4
020MVYATMixbtURrqBTccQ5TSnPOQgqHmCEDEnbLaW6KiVeHvt4T8nFqJxSZqj5g
pxMmExUoo8QQ9CiDmL3Qwno1CbP2GqtGIXruhTweWJLiDfDWoVG1J7bkV1uITGM5
tf7SKpA8+xF4O7z/4h0TV4p5rKLGftjg7j6ai3BuIF8ZV2Udu9IFnXfjFri+ZWh/
6UxmN1jIv1ZT092AHjXE+wLs3VvKANjCgc3mbVHFKfYvj00InDigXFj6DJAqluVY
6wzaW+MPdQeNKT0ISAOwtzB4uRpYguc3cAyljhprD7DppiLutmT94aTeDLomk72U
QO3g1cFWfJg1XMqgWGlxbGQh29qxxjcw0Ev7UEk8B5zi68Sk7kd5jkv1IVdOees0
VuP4QkXp/xqcQQ6ijjaaZlS61qAZdZZIvq54btAiyrgJFuLKXjqqv/NoXkozFJBU
0FQC9hCLe48Qf/O1PLZBfMiN5V0zahezGB/n+ww4ebuXuScNldZHTgxuMPOaI/bm
Ww9uGj1qE3ueip+2ANJoTEqh29rjb/2R2njNaADEneBidLE4/Y8O0HrdLDz+G8x+
Ln2KzI0kNNGOZBkUn+0fLPE4JUef/vyLB8O61DT9zrCagdAXTFSqEVHEViWTVCld
jn9ishyTocb303agd/UM5aAxYJq7U0c4k/FbNx77JP2tiBBJcWuXk0skMstCLHAD
fLRQW78h2hNeHlQXyian6NlcLm9VQRu+ElD7nULeeeZzH+3qnJ/sPOesjC0Qd/9/
1Y0ItivDfQBrWdrh+sMjAsgnsAvxD009MvT9i+UqhpP23WSW1tbmUeg5MjvO7h5s
SAnvWagrU6OgGbsLzqjNazEJgVBjug3znTvnKINxHhBOtqEtFk4viIuaxEMWHNlS
kXOZ8GYEtnwwT8Mdb/t0OkYXYdECO486/o1G9SrRC5VwzToBN4gUhtzrM/AZB9AU
1LduNrjIuldbLH+N+bpO00ZLLZFHGXhYQU+Ur6Am7454m8SkoK5nAt4GqYY3VrR/
Q8tjQl6/4SbsVZn3IKcr8QotXlpUfETYVcnT9fpICJahjTvPGdN0yn3EqNFtfiUC
+ju8J1Tr/nwfLEs9twqr5l81d6swdmv1xdx4ouEbVUPn2GWrcJ8qm13amQ6toQr6
vsDqvV4iPVqt0DS5x7sxMTEV0Rii/eKz5QvFxF9sq+Ijlri7Bt0WKjCY5Ko9ylim
LV0640h62qli0E3EaHzqqGQXJnoeRU/cGmPFG4cAvzSdBn9s804VI09PsJJjafRu
m8pVLQvem9f6WNMwuxdEucsMbJsOp4KY6TLyRQWGKeGdaWKXV02aUOAmo3yLZWDo
6jNE8+jbp5AOpX2cS9wFPSn6i6cIhkF0UsP/xITYTkud+HR937hupaglRpqvavdC
GjgmXu4y+m2BO/zxw8u2fbzkWtloK1tStKsgf5E1N2rUV/bRfPbdw+mh9qipSKkX
u0RAT/Hh7vi0UX6L393li2b3r3rixvb+YFHydMGzLVkXRJxjMLN2azwXNq4GVRFC
/4eGVdm9Cv/RRcbSPWc2Y8c5qw+W3i96ffaE82L3uCF242zQyjw/JQCONpRZtqxV
JKVWG3ZPj/zlgHLBEydtGkXIHnkWxs7S6sPcob0lz8TmJ4fBt+ZWDGcYPb+Ty8PW
Nx1sZT1cPhIcjABgZpENrMo9voy0ERQ6hA0JIXD/AMgXUyLplDgJsAld/uJjTjmc
a8xjWifrkBUNzUT60sHCvx0rtCXErfhWUVtLuCg0ywCLuWZWisSostS5Q+cVV1Cs
2DlvTKZ/ph8W3k8rZuNtIlx6AmvoOsuJYvndCjmamM75k+Y/L/gccHtahVlTudF7
Qgqx6OT3WhuupYFJ+Nf6jCgAIesgnqk9A+t2F3M2nYjZzr85FvFBaGPyKh+Afq2q
cSP5JYaDFQYU2kuLebSOX0ZqpOZpRzXY0ITf4OnlJTc3bsKuMsOtz8aM8GKwgaBn
X4g9ld2yaYlg4wPHDHJ17lNc4tUOFbXe5y+BlzlahHnh/6/4V/7hxUzqhAatQyQA
aSioy+jJUGLxXTYgSgEYW8C78psz7Tp/ih72tKzD97yojbSpq5hUDxfMG1Gtmb7N
vTSZ0LIRrs3Cqgn0LASqj9eNiiOHZxfn4pnU6AOJ88w6oyBaJqCh/dHRPOJK0C5l
0T1FZIKpTLNUhQGgmvmEkOEx4bXGTctmi7S0XZ1hxEnYwbB8kX+vm7okWOZDFs5Q
jmgt0LmLJUtmVQaN5VpFkz1Mrj7SsoJs9kCqRyeNXVNgGc1fcAkraPUZPff7tECk
u1mV2vbHHI/d07nLL5H5A1UudPjTTFLXFw1d4TiMzpkLTuXEwNesNIGXbRYpNeB3
TdYmdscAyueZxx3lTCTduowhrm5A6I+jKPZGXFb+TbiN9p/+oHtiEYmazBoYPJO8
qyhDQZKYe8KJE8l6lS5/OUdwm5Q9ROeK22B3Zc6eDplhhkSZyj/aIibttrPCEu3m
7mks/7qnRfJi8ZNnqn6RLABfHC5XDf9YaltA5bpZHUjkNpQ5ZZbguLjjDHMCqM2C
iIMJy+pJ6SzfAch/fT9QSYIXC8OT7j+NtREMXM6zn/Nj5ZI4QBfwcv7NpMB8r8Pz
saCtGYSUIdSSjlZJvClPGOAMPMxQvO7+suZZgMjKzRKdRPXUuk009Vbpi6fSW9LR
1QoCJI/h2HbmWTpeeMYRK7/UYBjSmIjexFmaObJ5ytD9sJ4RBMQVUDXaWJEbYJ90
6YjF4Z0X/lw+rcvhQdwHwuVKmN0FHZkbp30VpdWMrgGDEY27PU+FXdLCBGVXnlq/
s1w6FtklT9yM3zbejlfSoNw8DUnhSLGonR8GlqYUoi1HS+Q51K1wVmIQHAQpe3eX
BhB9vfoNuSqNwaIhjChaH/51HREoYw01qpzpUNu7Ipap/p6iDKE6Kl3grv4kFxq2
DmaPFRZSRPWcmWwegbB0jN+/IEV3pQsSjKYWNQJzpmVnFYVf/4dhdtuUxhu3UUVE
5WGqxMrtZe3GMACEU2pRbe3ZlkqLm+mV45t+Ng0SqM/CkgTN1K9X65GWT576WLj5
EaKpVXjX9o1Hna2SB1ZRTCwIEv8pzQBpM/DjD5p7DrZzzERG1enyAgvobvxEp4eg
NpjdZdXdhE7bMh3y7P1U83C/LCmMlhNonoMliewtDpK6V/HgBUssJGoTzdNzFHvg
POd5dEWKV+JRvJRVOjWA5R6AJUUxCe8Uy6PuKDqhEQw5xOjzsX8bLkMTFFTfUXQH
m7K4KxX6GcoIU944UFs6xez5TDHkXBGNELHcTnwvKsnUVLxRfweoXF2XiSq1q5xn
lPwkH4nwLeo8LFOAgolPMIu+cl6TPTt7HKDzUJFkbCdPgZaScPAynDWK7FlV96mt
hnLQBAlxkh7ydMNdqlmsh4Abce1GU0XbeKJ1iM9Kd1tvpVkL2ch/lwIlR5+C/7QJ
Xg46F4BHGQx/OK2bvQNz2FpyMAz4qr2SpwBYSUOBERwxOnWTdijoibZ8VCqoAoBZ
ddPWyIefTssg8A1c3mH5sUI/LPZbPz4kKTJCRxnkkB0FR4rjKb1KOOf8UG49LR23
95zcoC8HMLjgqIUfEsuSMZO54604/4ZsPxAN1nFfF921Fm/noQeHe4Ju3hVfubJn
Aj6P1ulnKIQSQmDxMdMB4Tw5i56pZwljxgHxY4uccckYGvKLqvK76q1AcQz2ljE3
C18VM0Pc79nzH8ysViTsHao/9jwQVihVBtMge3CPjGaQlIe1IP4kPBXkDS7vnLzL
HII38m00Oyhk8eWDnHRzJaFZYDF4AcnIPvtJUDeOYY1Lv/nAekhg3Iw3Ebmvm9Ju
nWnYYD5yUcaGTZYRmCWUqBGamVl4JeWO6ByY3Jt+nf5H8n/vAFE+NHLCTItxRVve
xrcMYMJCWg6LNzD10Im1rP7ND6TBkmA8mmTHZzug+8GfcXbY1/o11i02q8CgQXRa
H5XzPcQ5ugbHDctfBs91PzUm0oW/mMtfh5AyGaE6CZL61tH6p+m/TPV3Ow+CvZCk
ov7x1wPGp0P9yVs+PFv3MJSDnEyV9td3k9uHWQceoB5dMF4ZuTeMICqIulRb24zo
2EmhjOK8cqR/MPLAVwo+yjSpE/nirkSkGRwtNbjDdLqhhlRjZDHHlN2Zz6yTMKmM
rkYzCO/5HVMNPWlh4/09SlSvzVFXNcDyKEm7EOlDo5a/lEEDTQr6SDkzjN6U7eRD
I1DaHPx+Of94lPaU86AQt7SPHpIItmojH6Wf1692Xes6cBxEEFh0BxpMZi2eA0RC
E4J1jNr/7jnHFrVu59QD9heU9JEJDS435SKkFhGWybUNNCVMt2MR2PXSjQya4u84
ET8qNA/ZwUv/SCLRbgVj3NFLfRzK1LOQtdcQ7gh/+CeawjwOd2dcMOTchQN6O/KV
PhP3ganAyObrzxLqcmdereVx21joIEEk1EEZ7AlMOQ+bJVlcF1e8JmoI5QKRYjxx
ZagQSQwoEnaj6QSDc9fOifEbIbSDEIfOIpK9rbbxGV0BmTesGUD9OJBF3cdLhqJH
jcxlKMUz7LAUzlOrbbR+wCJWStcNqbVS4HtNRn6PBlKK6k+yJVIF6RQhgZT+V2lp
L/n+NsN8paRpmcICiJ8CL9NQbmGZ5nhgC9rtyhpJVo6kX6aTkwidQ4b0fpPiO7tF
DPtMh6whOWOrNqxsSVYWhWsltGh7t5u9M8S3v8Jl4JC3i9t7WyZCJh8xP5kpwiR4
JL2XlkzLY5ie4TX2uOzSCum8x+n7kce581TOHRyG678Oen3SPM3O8973KhQxQ9JX
p3L8veycYFZejE4at6yd+VDTbHU0DIvpFgOy2elxzOtfvYcXeFwJ0tCM6G9vmMyJ
rBq7Zpr0bXy8vXYN41Hl7GX3rS36wG7xHFTIukiyzOWuZ+QRDYMp4Myw2FFwIyfo
EVyD9XGj4HWBme3kWMPYDhx7ux09QmLWH1J4wtEWaiojdWuq08EbqoDOfYVVKBgd
ICl8zt4n38vW8JOGCIePy7X01mQDkFJ9VKEjJaWLgZ2CjNrZUaxx4LVVYvVHzlD9
7c9KBDePRsr8/ZDK6peep6xlvE/UKM/wpq3qAvAQ9qVx7B7Mns+ZBqXhSvw/1oD8
6ZAtyQVCIOSX9VTe4pKSQY6JH7DeE5c/tyU1xeHFDD5aEUncTNu9pvEAGL7NwLWB
s6UchU6+aiqlLz5uOhoduDyUW7kxn2xr1HeI+UT7BfOw5Je7tM7KMTSLmnlglNmi
MhJpmPJOepVwKwAuXEKEALaT2svz/EMcyaSMSAM2iCuZ9Ktw1XB8yP3DEb3itxvQ
CdD9KdUx6DrrKQlgh63v/uLIpYTg/rLzy82YiEuT21BwiX8WTHURXI3FCiE96xID
oCFMlXEl4uHz77LYrbnb0YQPBYXjJVSXBpFnngaW18ra2Z4mFNeL+NO6i+6DbPmC
NEAGM/7WIKZb2uxBbLM2ZmQlZuPt9XkHW8TJEf5FOlar7NdOxdCyB0OcPFmNR8xg
b8IBHMvm9bP7LYoOVIP7MxBnYFVtUJpxwqg3EsznZNKzd1v+PhLgJPpSr9a3LHeC
sKA3zzNZn+yIgj9z1cPVUXgxZLhu5CrrB+Iq7G+idq7RZP9vbVhxHX3dMqvoySw/
1d016+wBPJIcJVkBB/5cWswQL0SY21Zx7t006krtwwtn1PBt3WVbJPrZ+F9VJd65
tOQfAAZ/c/ZopANtEPf+F+dRqgMOKsI63ANPDYZadnccib2PqBAq4tTqQC+Yg8Xm
lWxARnWm1Ny5DCsWLSg9p6pCI2FvZ3yuerMLcwiS0bB7pLynQqu0SaJmN4M4UvNN
rf6nuGKzP8r1n57s/pxoObC/Ldo2AtrcjPJjkMOtBPYIs+W1HSv7/MgmjRUPspwJ
aEgZFb+pdEpYV+fuQJpmk5053y1UTsMIIvsiQSsu/9hnH7Z21vULkUYwW5lP3/ZR
mBd8CZ8gXhHSUnC/yAJb3GfArhM5tK09XqhI2VjmqqKtmMVprN64dSHRt2e8avUB
+GGl9p74e/RgKdr4W/4zY+NYlFtQqy2Il67/mvfS4GbwxjEMRa1q7SN9VXwzRMMx
kW7Ju4B2jHX4sFP9Paw/H2+LFrswgpU0AzcHqf6WWy/vDw+2+QsJuRu2uPOD0A56
ga1VoRhVV+frvzg9OwNs4aAqBQ5EKT7mbThE9Pr2+9PYGQ6CifBzWf6AXPg7xRDh
pgYVlv3r1FI1GabksIfZpyV6ueS/PlYiaLL54XsfqzEV645DH4e1+D/Oj/LwfoEl
wZd+S/FitbKskUVgzoUzmi5yxhm7VS2gNzhtzXPIKLuDgCuGpJ1pLdZ8cQ1OzPSG
KjiyyIdoRT+SJTHc7k/86oJIm/sQJItJ29nQpecl5+vOuuJ6wDBz9318mOpanLBd
6hfLDFeGXhoEMBwWxJ1MIT5s8lX8KlDxuR/Lb88578Kp9E0BfwZJj3hru5rB8BIt
74f6xeB2f/H+WHzKvj/Ojqe8w9jLRFcv8Ymm6azuHkdC487CkcXpgFhFpeWeHear
Bh2xkzZhR9YmmEdckXDqgkrzKlNWBz7/CK5nwnCB0tyBgp4JesiICv0OU/iu0Hlf
R3RtoJUhpLNYdtbGicDTgUWzyNZdi/4dQ1/Fw82QIL1ExWwEfDERdtin0dwSAOYM
yBBDE3N7jw9HrCjfhKVwR3UL7s0BAvvx2iOHuKgNVooBtFCZHGScThdvTpqx/Spw
/GL+vbpZ4/QW1eMV4zorywMW9RJ4WHQhPU+wKrY9YdL8R+NelcXcxo0al3kUZJP5
UOIYPiQ80M5Kob24leyorKB9BbGo6lTXG33HbWEJsoS+xFjQxHhQYfzVUwwDWwV/
L4zodGGbPRJLIgixaaznBYVYXDzkh4ksMI05qhG/MZwTXVkWpRe07uXgjtpdS8AJ
R6q3/WuD3E3r8AM4ZaLccWa/B9pYq4qGlGVE+Txaehp7pYolVDHZ3GHE5kjguVIg
3QMbnNV3ZGu/Kh/T+t/emGNftBQL6BQFxsny6whTySz0U8dTpKdcKw1L/6+OWHYC
dsck8i7Hhf++oJMc14XGaxPLRKOH6OqJs2d6UJ1+vl0SFpgB1tMwYx64OyzEQa21
ylOZcwUWcsw4PC6zQez76erHYxh7TWtDhwTJ2CYPid8c13ZAGJhbTnnN8wVGirJ3
H2Ki1SF5a5afq2Ch2oUN0tEiuYAB/nnpa9vou+1CB2894zopZ3P8TUEfzSfYx/sK
4WZTOjkJSqMZxcBR/5T7nQCtdeRkVY1yPj9GYjxfug7NfaCtLFeQd4PXTYvbVZDJ
cuJfHWCbppLi5JRZA0gxgKY4qXuN3hY8aJm81Rd3XMBSFmT3YNZUyhdoODKYZabs
hxoCsHs/60mEUfJslbuakPAd8XGYREWEASq6bY4SeEu3W9dzMEyr+f53tH5NvVWL
1baqNkBBpWL/0yybxP7Opm69/9KlCIwIfSGRQiLAQC2VW2uE47FAgu5hRnxoSOto
ASIs2iRdqXSc0m7KqqAZWId17hWA8b2I15bkX/Oyi2ODI/jKqz0/a+KtcI+v/m0L
Qr0tNPtNXO7n3avwYsooyige48VrFT4ZU8Uri0ebr9RHmPVI2eSber0w9SVGMUV0
UBv8FUlCZj0RjvcCMR/4Bx6PwQJtJWlzVsvfAN6R3KbCzDyVYsv91ZcyEYXYv4k9
oPXGOL/QET/WrzQda8AHRw/nQnEH2aOiGFsdM3GMIFTzmBmYKAADYVQ33j4L2gox
igU9b3zk02DzH8QMeW1qMTvwJoXs5WwGfoIfB0PwCUkw6Cyp7/2K7RcIbsRkqlUy
3gWGwv1Qy7Gm7TbOrg9xZHUJiF2kcn7NrUkcyZo2hJJHLOaEny+9RnGrtmuviELC
/59ij119ACpY12qfi91G+e5W3hABXgNaUxSBV8KvM/qEP1Gsj/fOeXV/7kdtjcAB
hJl6GXCiY6fe2hZK5Mb+SYb5zf9HikH8MIbX2NQYTfNpJ9rDXjyfATfXYSghssYs
oVwQVHEgT2PzjMkgZLqEyDQVY0fWKl0vMa4Qf0F0Nki5NKcnfQrTb2MLgL+6qM05
hMUHb9P5w5cdvlXXJHy+BsTCLNCvpvsE9tRnQ5cszAdNDL160bxkb1zksmfkEmUg
96yIG5mXv8xaRXV527ziRxswLT8by0SUsU9qynRlVsY/P9fht0Spb5j3lAbyTykS
6bOU2OljpdX4APtl5A3C9ALDoeMoiFptJvwI72x9pCyx/oJ0+QcC8uU55OGKGqJG
ZBCHxLpxeEG6q0GGl15VKYtmug06CWtmutnucAlYQGR/8DJ+LkgVDOeypCI4RxNJ
bu4wIzIGPVdvuaUQ2XY7ar8Bk+4JBhSqKZi6Ag04HclEEiCtnMVFlfh6Fd5aRk4r
UsPtOXRkq4JwJHC1XpjOJc6y0PfXhI/Is5hbH+dFh1YT5BT8n99coMzP6YCe+LQu
IxGRX3pRSW0W1SOtaFCamCSMf3pYGE9ADuqiCcotB1jBVa9ouhbSd3QyGCQXRHHF
9D1s92vHRBROINmpoT+QbREjeZnI6Lad8mT3ETJULa6GPYSLQcZcc+PsWJrI0MgB
VIXOh51Y+zT68qYBm4oM1AFa/cxV3R6yc/tWGOGZkHKI0RDnZrw/WOxrXsnRbQtQ
8NVLdWw7WwEkVojggh8SQFvgTXuMSTyReq++XyyAIbBYsUSb3iqsesrV7MOwoSdD
VKeSrDj0OVU+7Itk6CMX2W6JaVUjCyG0p7svPn+IYKw9W3xy5XcFiQaYJ95iFU65
gcFgk77E7wnYNRD8xcQlhJ0bD58Z/pOu/vBMFnN2P58kyPIVaN0axYS9GtWggB3d
AuQn3U4y5VKfuDJVXNal/PWlDLgQd2PRGMN8BZA18rVVCtZq9YNGFuL4RDdvUQHH
uM3epps0Cat8qg8YNaaV4H0dyPrn6jRFOBWRoMhGjUzF7znlgHp/DIHHcZuiLz91
CYccsESKt7SzDKaud5WpoHXQ3tsoFDz+bRhiXdiKniefsPqDulDTraDLjIlicfHq
XOrOfBxLqES7hBlo6rg63S1cW2/LLp2N0HE2c8lG8rKl1GJF6HskaTheR9bl+CRy
RzmhJkWFgU/q5YXtKnmSX6WPmJt84mMRhK2Y+44Dyh/i3G1TnD/eRtVUPllmBbka
jouE3YRVtkww4LNbzVH8Dmbc0M/rMXENDTSs/dKWRGEUyrtmuEigTFqA9VnTMOq/
n7Uw98LLnM6Srv5f3PivWudsb13kueShGs57RFco6VY70La9UmWgMsxVbw1irC6X
2QaUlTk2oUjW4lWWUA15iHrl9mRrfCcHvVD7M4rlLrWEb8ReD/S8S0wrxsXwGb3h
7olrpyKZtkl2bFoPVUqyZFfxos1gsYZMsy1QRDUviIwNzoKPsKFOrwGgb2wb1HP7
x34McqQfKFIvsXiUuMuwgyY13juA4m9M3M6xLES05mUPAhYBL2X4VH8RSTHypTH8
RIYrGQXD2Dy+T8Zv6YzNbYgW1119NvEblpE5sHjIluK7YJ1oUkwK14t5zFNCBWfj
k0NqCcYC3tY3uQeRjOrNLuG/tfaQUeE+4AiGtmGKaaLu1UNZXCjGYkRrqPD4KWDB
dxudQJlvdHL7SQ5az2p3R2aG3n3OjUSOsUodkdKFRgFLgNI+e3WEcFDOCVq0B0kK
b56rt7DuXvbnxHD+kYdQ537YoclB2h5mwYVUGaqPXGQG8Fm2fMehpIOGFMLZAWP2
2oQ/4u0UwwuyfozRhpa7jytoITUCS+fDyO6lIHX6PsZDtWgtgsglGdSjfQKlZl/U
+n5xoaCg6V4LsTfWwGO2bjsgsM6zuCKnmJTxVQI2T7Td8j7tjmcCMdJIpUM22dcF
7kgUJVyxo8SKFcGgN/0Szn9sT82vYpW3mWaAubRCU4ZwIJmg1220vfewSWsLSbr8
z0NehaB/Yj/YVHi0gOTpypXUNocMKBS/8otv9RelKuc51gZ9qzVGuSbMwLz4axs8
J1wPvNMyioXNCkZF/dEfEG/0VM+RovIJDTzBiNkRYOlMLm4pokF/tzEx+krT964Z
ZnHPVKIqyapP3ENWXNrrr324bP2ZJcWdUFy5A3WV7G1tXccWJw3cGywBqV1m5+Ka
w4qQWVBHifx2Q0+Zth4QajnOD6Dn3SVynH2AgKBkBxXo4xb4ybDD4SbURp9ngBRH
uCT3uvJGnu6vjedClX/meQzTkYdYaiy170IuRZaiKC+QQ4hgfLfCzp/5rsQJa6hY
iZf+tZrCPXdrikVpFjPf8F4Vd3WyhhXoGkHR86HrkIyXeyWQ9I6DoT3A8Fjyu7TK
FZrgVfSouBbxVOevMtcdEOxC355ZiuW2ZuAO43k6PPfzM7mBcBi8u+pikxVThPxP
LxaXcLs0RhEFFzGTSRAoBM/mGyTJcTYREzCSQO9nm3pMtQUU5egjg69Bjv2m2Xk0
ks3ZqLbIk0aXFwROK7anteB3u3QxlRHiFn61Uo9XBG3ZK2MP+L3qEJXjofaSKpbo
efeuyztmUHGVyH//IS9xZGB40JFvaZ5R5FC+pEKdlUFLf8CHlgVyD7axOcjucHJ8
NKtdUydFIyrlK549dBj6ivycP0OVho/WReBNJB8P0uYZ0zzx1jDC1/KjuiHEcxYQ
6HNhSMWkekO3Cp89DDLnPdkk8ECPCPjd0htYVGdcFN1EtkFOlQ4gGx3qTV+Av3At
F9cT5zpgYlwxj/7hCWJzocGG8wbBV/kt2TdI3LplmUrngRRVz8iTUJ+itn+oWTv5
cg7m/hGP/9wjikqxwVv41PA6/yGTXt2PmTGmdVZ85mn76HJTrQIQOV+WoWwzmVK0
/5HgFMmwuR5oRfV/JDdYQ5fhkchgrdT88nR1QCT+FcB9G0cUrFD5vJU5RBXZkveh
Ysc3LSnjUBoXyEXilZMZR7wTea4nKjmeb2Gc1e081kVOJeQZDdCCnQ2K3GEm0tUH
eY+gML/twkNwBNKv7by+0655ITUNrenpADEALBsnU17aBLcBa6eYijoNzJdnfwYi
C4GZN0WpIQDMEfH/xq0WC+c1uZSHkXzcRzpoGZGf03ZFRHEOraJ+ZtHZPIckqcHt
Ht3jAPWnRHSlCxGwIt1aJL2TtzMN4mts+tCF696/pOOLGRCvKsM4jghnPLBbYOQo
BzewJeWxFSrRlkOa+B/Zh/aF4W+L7BGm98azwNTkSngwjfdgxtuZNY5LKxsKkiK0
Q8kJXWw55249B6ao8a8QvhmgKnajsvoGhJRFb2YDxABj6BddqXsEmHjmBKLklLXK
QI5jHtTvnc+PSFXBFVBYPrNNPkZjxc0qLLrnh56Ht1/Umo4GaxHmL8tqwvPSDKHq
k3eQDZxPxlgEXiCVa1XjDSI7YsyfkOeygOvGbrmkvMzihsrBRmwl/L/rW5XLQloV
EYpjiJT+vc8s4LQTJY+NCLkm3/I89fTfeLL4IS4efJoJFM1mMxo8TIMrFg1EHvXS
njt/B41gTEZxJxv8kROfQouOMbpQEcjDz4reTSBZRA88XwXtIxkP9dijeuRxxEPp
ukFt/bPly6Lf5GcNKzps6le4HTZeqJv3EW8Q6QBg7CGNLP0JtOBNpWvK9XETZgpP
x9whaHVF6Bp/pIqvACWJlRUzs4C/ipYDB++x7ys2i+q6rS2YUyR46Ir2fN5tHvsj
8Tt2k3m4lKQmz+JuwLAE8iBsAt6ESnlTgfg10w0N7TDHQj8aJZfLjvjbD5pZBHF5
OMwBIne35bXolsYHnBvd3AcqHgUcoo8+3ZRVGdaOuvbjJEvZBTUPNrFK/AzQhN9j
HCiV1ub4Ve6FtHc3OHFS/AJiAqrIWP+8/fu7my5XTIt4zuJ3dlnMWYc+L7ezRPM4
nHLNY1YY+koFKNr0co41XCs0HAsfic6+zxrAhFblpjOI/jCCxmXvbzu26IWK3LkP
eNSh2k8ymSuRfIRhXTQjsnGiAc7VsX4IQ8zY+l1GoF5Mjc4UVMhD1YloON5xgO0U
mikX0mkFDldbRAdSBeUC7HK8ETsa4IXUlyNR193zGfiLllMnVn4HVd+EUjOFaX8V
WBKleBCcTvjkNwaxs7QnOfwejFCyiV++dkLEXAYJh5vAXK6jt42lhG4LPkGeTbjp
1fiXzG9rmQv+sqggkuxVuy1osqHE8OwDnf8GvGG87FkD0DuNWu7YQ7+4WdW+4+k8
YVwvCwzsARVcJP9lmpqPYCeCnF5hbonca3KMFh6anjWzaarMwAFQkEoVORSxPKJW
AD05+5gs36YQbERslgrQp1TfH6rBBabG+r+n5DRGFWIaT+YBTKhrO6B18qPEJN6/
MDN+POUx0VbbK5oACj84+cHJT7r2TjepmSt3hC7weEGWDtbgmAPT6UpgYFDQkevZ
nyP2aZVDTdLYVP1e4Ki/ItBe2px9Kb+096t/rYw/t2IbQztrJwTjDxK9pl6EiwR5
wTHO9JJdyodpDKLmZDemSXmB7EWVoILM4EN8VzqC/xweFHp030PxAjcjnPUGJSjU
uX8+jlmWof/4H1Ffw+jOWTbcJylVhZszJIXUrDtAdnyPlPohekdToj16VIl27qOR
0YcBE1vIgVB01a41i7tbk5kdX8+Z85e7u//sLnMfkQcvSKuzvVyDdg1AWqycNHqr
4HlZgsP2OVs3++Xym1TOM+1AmN+ZGVunKG4Uj+r01C9q5wd3XC0+E2jYtcY36bGE
2gfANtw/8ujh+IO89Sh5B2LTorC3W1vqlFH5VejhDf2uMjnj9c6M/2550lyKd1KJ
j3/cy6WUjvr8rkwMWv/OHtLAJcazQnp95Njrdf+P8KGB/3aJ9vpyPlG93ULFFY1p
97Jx9SfpVaG0yMsilbdKn30diTwm5p75Q2ULDdzf7R/H2Ei0e4YHIKvG6OML4S3c
KK8QE7pK8RRfUajvrYNRVNrN+gL7nFKxB6boqs/JZ0Hxw43mxZnoRMaXA7Qofg0A
YehEW5GNELiMYogO9gYjnZwFTVU21fuuxp+hYDIzo8WpFoiFYVt/juG9aui8oeQd
YT8Ip/PasSFDedzanVoP/slqeqdBJLlA8vCzs0tpZespeZ8M6fs525X3UkQGXIV/
HBSzNNN0kNa/LsbMATpAcVrrfHbsJHaXyE2yUqOgVyzcDidJ1r2OGFQgO1ttuZBn
zkkgd7+KWD4r5FRQ0GnJbEaO6QZWtK2iN8iUnKXw8oIOz2/LB9r35aJfztL2hbI/
5SrdoM/jYSr6+iRR2xowSpv+Oo1WbfFyWgNGpa1/gvjfxvU+p+ukk6VeG/ptwM9i
l3T5hFMJvzMWYWlsEy/Lkpd2LVHRRc6ikNO7ZcEb/NT2Irr7G8MHN+UVwM6WW5py
yX1kykx0dgVikm+i2k5+ozH/DSSmoDMUnAeQI/3gLh/j3e2PiiM2oCOODcOnwvaZ
Vt8E5MyZ+8hYt1EQe0fTdP3khXY+T0I3sCRhE9tAHBoUjC9uk5VBsFdKPQu/hPuY
X/pu6wZM49cSR1ugu1xfJrCimHAM3887JgPEqp3w05WbtLa+v85gWMDqGUypvjhF
G2/l6+Pp8l4G3pOGhuhYYHgJWVDZu5Oa1bETxR0WvTUMR2wTg8C/2+pMBN5UAStG
LD7JOZ2IziOj9/DtSSqCbz2a8jnGn4wtAHMFSpWoD5hz1WQ6JikYAndUjcqHUcWc
ua7UaYpiCCaBO1dA1pY70ogs7pJbADOG5hay/t+4Z9DtMgk1nw5e6Y3bQVFlVpcD
WjJbgZWIXkeGHSatBAWmkKiBR/x1n6k1ENRuBnw5TUc/TRDEkbp2blqIFqzYGITz
CSR+9uvQRm2gwE105A5xl3jhF2YK3cjX5tjWZgZ/TPexCvpyP5OA9qBOUmrN4/OI
mriBBypwkfLgKzmDrJGqRLIfLgUxSkh+0toAQs6K+S020i4X/SXh5zwqgUpVAb++
K+n2bof7P3IVBfmH3GExmjQjceUoyUQTjkVYfdZgklLnxubBRkXP+FwZLlC0ljOT
HZNFxH8v3+aNMFDCoXvWj4hRwe3M5rbi5UKD52KcE9bMiU5jCuZvxX1qqZdq9ClM
niKz2kQVct9dMM0J+pRqBrGoOEe9qkHZ2n+ojDe20zTQedF6rXDF1QQxP51C3RhE
iLeziU35RnAYRrJKj+TpnX0LtEE/Kq15+kBZYLjrgzNodGbR+w8SQNCa7et5cpux
7+2j7NXLcEE7Pc2eSAr9RS3qmtdToR4udrKBto4eVKFaCXd7IoXFDLNTzzVeqq+4
DXUTvFH9V9XU06ywV3XeEnxlxj4FID09/+iBD/UxFDUmqWA2UI0j8YVKSe3SF3yu
CR6C2ljyrhWo9je3TeD8QTVcW6dZDcOqa8+hyf+0EWpxKSX3uQ4oAB7Imgd533WS
KBZgBYez4Vix1oZdpQ3G+AsZ9JKbdRNZhPycgmFj9izuA5galacJ7DYzdXc6Offd
2Ahso2FgOZ9hJD+CB6gTVR/KG4nZRRTXhW4r5ME5/MBzmMkYbfil2hclstqOFXbq
WNaAFImwWYaPrNM9Go9xvTys5i5MqhxH7rZ0p8/XjTDd1Efo05+f7eWwejQQvITC
vpp8nczCOX1yRYXKUP/VNm+V+H0ouNjeP6ReMlEP+a+1AgVorxrexf71bfo6n3Hi
aUl1MuudtbBB5rUzXfQeCFpFc9mSPchdX0WrZZSck04iBbTmy4lhrHLpmSddOK8V
zsLts8tBKUhKEPJq5AyduQbzyeSDdlz9srAqBbAym2aOUofdDMM4MHiq7t9ZCLXW
74Jx7a8cXftCed/cvJAbowfZRo7egQRIlScBGXBS7zObTYhR9ZZjNizbGxNBmDxT
+mib70EIwL6DT2CV29m1knZ7qMQgqk0dEDY1kXW/2u5JLE1/dDMeg48ebp4WqJR2
2CbQ7dOEKrmmohLmmF2oCmc8waLMZ/7O+gVR9p46Y0TGa3pF592M80OmGuYylU04
qIc9zPjt5G0/pOpXd+mjxHNdol4XlEeR3vi2mtxMYAwvBIUgtW9k4TjGAHdjxpZ3
kMdTTX03c7wFHV0W9ZTsXlC6lpC0fhq2Zk/Q1OJHwEu53h4vdZfvxvY8XcKhhjTe
ujDzYEnYkLO7aJVdAt5vdcFfbfaVmV5z+L5SGCP4qrdOeoVc3rBy06++2AU/3gS4
TezQje4teaIM/43Xfwto9kqHh1082VUMySWAccs//7G7Wkmayywpro8RwQjuIF9E
K9MFLqWQheSl7LsI8+Bcm6lOdIulzT8pH/zk0qgQIWfsJ+uTVe2/qYSWicUMJ1ny
WsLECIZjYT354ezIy6QMNmgWgPv/3lmcaKFfUpdSF/X+yyQ/0xo8cOj60C1/ZJ2r
sxzjkZi7JHAiAuaG3629AcneySAWSCcU3K4rcbpTMOrTYyaLxr765o0AfoJEmITI
58pda4ZThk6nWxySBzbK6+ulgO0bbUOYIhA4ErCaBBppZ1APf/aEXiIVO6YQko68
jciRAwrKEzIZuQIclKy8RNZAkLfoCRcKUpP1hYHoR3S6BI2kMa7/Jyb2HUwQplAY
AlACQgJmQrABw6t4RlZ9/qzhDMKSTjNoCKaFH2AQtt3NHcVmMxAeXQ1eNEcMI1D/
3gC6pWiL/lEHHbqQib6vkflsG5jNnPjSLlMDGQKBTj5tRaVZSGPlYWVCnNYVi2mq
Vqcm9MvmM0Y5QNhM1SYYjY6DFrEjsr9+9vNXM7y2HnmswS4SUGCSCyzEAPPUjYsb
x9qxyDLNWThklBWYd6uXI5jLLxfsy1Gfq5g8PqTclr7VGld/9UrdMWGOTadPuzAI
aIXViiDPITidkz7L9Hd/Tq3Qvey4geNUBO9eztWaI2jljx/gn6qL2hbJTXyjEy/m
pQeCy7UZ33NIxUFHKWUVi41K1c3NzaOj0XFHfn5cq1iamnjzobPRj6srDM8e3iiC
b05SJROAjx83kZmYCOYYb05vTuuEndIbND0hacxG8Fp49Zn43PMl8NJ+UM1wlk5i
f0n9dwwYy6N395JFdzLLrivnWJXozPcpJ+AjTHMFkJXmwDA/TGpEfcua++l0ECC2
3hb15vBmEKALiW7H0gMmH/U8R79IkvMi6g/eGbA2hnpZ/FpxctlSH4rf59AT5Tkv
XA1dpF4A8nJlN1zh4ME2h+5rLVQ46Kq1dvIUN9Y98CRPFn6NzaLWNDCILeUrXt8Y
hfbRWcLG7Lyh0EYuz2JFtdwvvANlop1rRL+u/k4LK/4dBJNyDXBIdEVyMHwYwreW
S2HiNggYOO/ndzrULIejnSphkD6s/cSeq5WrII6LKHLQhXMncch7dR37y1I6Y4JU
ZJF7wy1A9oPIptZOVPEPVlhk++jBJO1pgh9dq3yCX5vgk5DaS9w/1eHmmmw86mhi
OyEu3f0U8K3Z35rJ6s+mmGYoRDnbb/eizxEMeIAgxDaGv8J3+UbSb5J/A80Vb0VE
lYXzt1oFT/qN8NGzR6NkK2U6tsRCutAzgKIzTxGKfIiOfSVBcT4O5YKqn6pTluVQ
hm4dSHbRPudQJimL51gRExpRRpivdJrrKIAbGH3VpvrpkqczPoT/jyrSmaqtOWQp
VGDRpldIdAgY8UAOS5rPWfGngNI6OCOzuQChHVsPW0mSXS24nlGjKhZ0t4J9avO/
9lVKwEY4qmOeSsJ5onGHlUgOglPjU3Q2buY2JOlkKwYZ5MoKLDUiuzKEHlW8XNPa
7Y8qW5Kjj6bwc6+saSWgiW5zFwi20Cli7iepihlWrJja8sbAbPtMtZ6DZXfNqwNL
XnnVFcLR160MAF5sXSDADQFe8XnG5tx0QkK4gbb5UtBl7zJSZFmn5sP1gNRzKD45
bKhJ0NXm1bkjxI0VesBpV8m4fmD8GVVUqzJwq7iDQFUo7jb6uitluCHesUvqvE68
o8m7nW6WlpNtzBPv4o1Zyk/175IEs9k28SYysyi4TX4wOMfhSbaBnbrULeWyylkV
hkwNuWA3LmvxypCNlo1QpWnICIsn6Q+YDwoztWxLzNL9ktM4yPdx/XFWsE0XSIPy
kt9gr+bANtA8FwXpLMHNEKaPLOIjn9h0iDSsa2fi0v2FN6Gusy22dWMbuKs7lB1I
5Vwg6xzBD+8cJuQW+9mC9Qqa+x06brE1eI5HjFzVYysxjaXivgWwqqMONK7Y55OC
TQRYE0aWfYvRYimUFV4ThEWj91zLCMqBSNIYi2je9taqnxsX8yNAU7KBc9JqVk43
ImsDH7lEEyN6MUGdTby5y+Clixd6Z7safmPNX4ZesaPDXA/d+K5yuqaRnaqOnoen
Ed26OMuaKKCtn04oyf1t4Ms18Xd6uA2+6V/l57wAzGk3xJaE7J8zHeeHydwpVPVU
3VvYrdlqjGHim4a+UF0hYVNmJrhcz4V0inYCEYASd2OLtyKiBtU+7KBlqF3TRTjo
yrwDtcqE8+Z3DU5su5Ae4FoMu0PCP65tQCScAX2cu3h+96Co8nU9MGFqZ8aviorN
bpWTi7Kqqfpro+Q5U4fIcEC2JO1j5bkRM9hHZbf+hBoq1OpS03i+Xwn1wkZk76TW
/AW0twO7V5wr8CkuMbsu1bnMAPwlIMzoXr38wRZXJu58uXmpt/+nK3Q4hksTLuro
HbgXt06qkcA0uGMCkcwzRdiBRpkb1Mo1Nv0MCR3LykYrX9zvShlSTUkmrLZTRS5M
XZMZyecfM8A0k/GcXJwNESdI9YjRWH+jh7vQdkT2644+Z4K9nYJwKIlyqNnoW8nV
dCDvhSzN2deWN8tJJ1JZYdZITlyWN1Cg4qYa9SYKgiIoydlYRLv3cnt2zZjQJZhL
KP02HvEc0WOdJ+Zq9mKYshj4W+jZn381UvIGbv3FRA8PcUuJRB/rOwDjGMarPn5o
vuQU3Xuf5QaPPR7MbaWa/SaPqawFFPEdrkFpwLJlo14DQQWAtvKOWaDqY5yPEqxK
jUMBl3A9vAT+9/bHt+U92hfx50SjzKEw4K/3uU5mWAbWkV+fnM/+ag4EdGkTyJ8X
89JeEW98flG4Ypm30MWxcSjTmQKXspZ0KgVT12taOjCHV4zoFVPdzOJPO7JpH5SB
M2NIhUGQTfTk0DugYHALTX2XXcT43RUptQbFhBGR78eGkUfuy/l+ZIP74s6iQiEy
YQe8j7AMTa6dVi6cKl4v0DpET31qpneb6Y/1X0nMIzon46QElBYJHWmlmxCLEFqj
k8dpwOPYEJxGOTWrDA4QQPKaBKDd/bXNDzZrAWf3SzrTuXHe+1838Ka2hgWEpngo
s7Qs60hPsBowXX/LlEyYKVjALZmJhE8G1zPtyvtz80udmAYwFf2WEXfvw81vhUBC
tsY1kIpJCHUsNDe/8fJD6PRNC3txdn1iJ7C/wRwTtbjUm//LS+rcHRqjYbVfXTBH
FftBmFw7OYHU3mQf9ER8p4CNf23TXAieWaFIniM8k4+i4XGz5hiMnM/My9RpOdfu
mFLI9eaRfDllKXIJrjtHOFFtMdAso+ImJJ1TCzS9yNgha4nwNYJ1OXW0yqnoCaFW
PlMOj8gjlbG8mRlgDwwzqcUIhwUTkNuc41ROeEOW3FHYrwF2g1sNMJZM3JQ0+qux
r29baTf6cAdOlpbI6xjOb1Oz06RFMIGDgGP1HzAnYkm/eQb4guqWf6WhGO8P+4Sw
jeyxPERHXzev0bnXKwpaDdLnebFuzLK3lXpdFfSgNgkS9zdemNwOlel/GYyXu9nx
VbrnCvDewG5mEDJJlEdRkdQcRABQgmSF303DBV3K6Mn8JV2jjdRNJzfxyXO+0W1n
jNfeM0DVZnHstutVewt7vguiAchqGaVoJCdqLpZB1Y/rCoOXXUgcLDTFXDCy1Hvo
RjV7PyGnmlJktGRrww5A8dW8QqozwPH8IqOlfZDcvo1G9NBaxrXVIIxiTiZ096Bv
DE27y1Ya4/LEmdxdWqEZvAbZ5hHNijhlGJpkGm2xglujIBiz+bbT+keD79G17zPg
CCOuaY0JEH/w6bbdWw3NIbFx7PK0PsyB3nsUAKwTpPXumpD3xYFrcyAc2CDXl3/Q
msikHSM60VdfzcrF6v/9nu5HJaXn4IN17IRtWs2KUqzppxGB6xy8xxDwLAFejpV/
taoJhwrlT9c4T/HnaHdndbICyTrgiYAQVha3XkwhcwXzS0xnML7R86qK/CLTw5H9
HApQnbvUPHWrvaBmZHCcFLIozNRcyoy4oFQNVEQBipmqi2p+fpsFHZDS/5pgeEoQ
yKWF3W88CvFegupqmdVlTBbpRbtp/oWUkDgW3zmnar7rCzmW69c50NUX4xt/D87W
ZJW2FqG7g/BzSAprzb3rjDIyWaJ9lbpmfstNZxrTGekfhhwDcJ8eFRd75ku6/Q9U
Vz3ay1Im8C0pKXysI4cu75CfckyaBmfj+h+ck+HbfubY2FoAkpaoLVyfXB023Ljh
+26JB7LhNn0xu1FWJQaBz3PdL8GHsCcPEqp1h+If7dI7A22kkblFEwGHEBKXbBEm
X4Tq7U+bklRwVAWya7cUAPeLuaryfk8vfNtt2t4OgbJBEx02Kv1Ysto31XFqhL6Q
OF30dd5S01R4WcpXEJe9cbS2Q43p5/t5K5iqyDUEutBz/I/gKKL6L8Fi6dVMITOB
IDKr7+InkHTykrkcYxCWQLHxRkIGN9rvGygWZNBBoQunX4uTv4wBy0XPZ+eFSoLO
ub6iq56ztQSOlbBfadNhrJw2sy3hLxA/1fUqP/in/5k3fEIWaC9b7po6IpTgNlB4
UBHMYCgVvNl6nC3LndAe0QHUu/vAuSVm9PxaJukzBwUZ5ICutWfJS+AxnNMJ1XA1
flGOQjS2HOqF/ZR9KMPoLnDQM1WNXieHOjQ+dapntuyBijMXsTjW7+KK9J2BEZhb
fl3LkDbFueeg/6WlQVtSQfiaO5hrmYFXwC9Ml9KnzzmuJQ7vB400emKC774IWBTN
LvmGZHJlkdLJGepI6vM5fUt6FJrzq9MRhjzVUhm1sLpNQey6CVsWWgzy0d5UU9C/
uBrMcJpg5mrQ0R3AIoLhGEUx9VzU4Kx7CwyVmQHcT+VRmJP2U7zuMD/tMMu5YQ2b
ja/uwzRuhcDD+JXZoDY2TW+Cu60sGzOKH8jm0e57O3mGJbh0KUitOo47OPmccLuf
AfS+GMp77h355JwwLxMijngCZQLlBdQd8UqzTgwEZ7qTMYKBWpfPEWQsM45u97oK
vY2u4eF6as6JTOwO0mOiCoZ1Uuu54QbfOWXa68NUkCzIXwvK7Z2DhXH6BkB7uV7G
j7JFe3Ut4DgdR5ob1f5ek8mmpAK6tQnVm/3lRqvaaTYxMr9ShV6zjzxlU9MBPH2Y
lcr8TykjPJXmly3YanAJ6jMSsVgLxywQ/RJTgrXGU39hBXFkS87LFCJGwqOlfY0N
YBu7w6EziD5fF/5a9GQIVOARtCk1/p1SRAdE6jJE1axymHwMBwBexyp5v4sf8gqJ
ZSQzQLyIiManEHws3Bls4OHQrQWr6AC4fxDMUzHA911s/FSY3UbIxfdLfVcbfSvs
rW6QwA2jjPxfinrg6YQ11jzn/I7krUSVl3ezYaCVgzfqD+eLcVszTOwvuHptWKRk
5WSpCwlkpV4VrRAVJXsJwh24mcTJrpbM/ugvxzofWAq/GtJ2YYsD8et0oC85sKvh
yIhu4Sgpzusn28Swp/pMhqtGsIVeNfflIDHPk3iNjvaKkv5yk07DetZhCo/wCHWf
GYcUsZ6KxQoKX1cR1fBiQDolpwoKntc+w30UZQlAJ/VqYdLTfvLmA2hiv4x4qIGz
lELEAY0xU/ORFYZa8MJMjaftfi3/FaKxuD3KGPH6/TKbRk0IAc4O8ttXJwrN1o8C
fwaj4Viif9oPV2b7/BqkJ2AMYJAEgWOpaWpwPgrxMY3IF1Kf0j5U7fjxKIMdfh3m
8qYYL9Oxtep7/WAs7Q9HR4mwMYTqZWAvyvnUnLWZOwKpfaxjgI44l5wUtkBa+heJ
JSqbYjhJeUMuPQo5fKX4wyZhq07iGv+cmQ1gN/mWkG8l9dtXTKqoTbQVvS0OW3t9
AJlOBmd2kTL2VUzsVPiljc9/A/3UTmgB9RHEBLAgSm5lLkluoAC0rJZ7oclMhM+r
rwiAcxH3gxG4IdIQ+Umj/P8iE2fsyrIrLzAuyvvb5ZT9PVusel5cN07xZElE/8AY
DXhTBUEwQIH5wmUq/njz87WznAVcPu+iGVRwoh6rA5aCn1uzWVOfFe0+NdHcaDCz
Et9mOER+TyDkPuZ7AT4dRfUElFnXmnf/uEjoY08XA2v3bfbu2cKe9K2Dse227MaC
xK9p43LPU+A48HiIjHlhkwd0RJkdeFvO/FjbctbepcvqojM2Cvx+Mu0W3UqYAaCz
A7oMRz7cV3km2ZgpvFSLPBxFTw+B4+p5l6G6A9eSW23bkvNls5ffa0ZT4NcmFxu0
bWzoBFndMwtaJ2PrdB67WR2dEiskmDtES0zSDxFKpi5FTyh4FIOeIQ5mLWzp/DHq
10Q/ALr1caPNqolMRCXIUp77vrj+lbo+BQo5z5LpAhUppcgqTmANpPBjUkF2whLK
QD5E8MMC0SAOtObRUjbpNRvYqIRB2/b0Zt0GCXkCb11Lf5a3bpcG8cQQdrEK/Fvu
cq8Cv49ySqjUtrQo/k136M1tSm/HkIeA7pbYQuI/bvXN4EOU1EYBUBM+rnr6XlE9
GBM73c+Z9x2ep4EZ8NG/KUFkl3RO7ymyaG4EU4fGHoN01NvJjAHF1DTOpAN4Lh72
VYBDPZDOcWeuDRZV25ctEWJK8LUyYZIzS5+onA8PBclmsLKZlUpRVQQ68KcFGYBN
vzuAQii8FXnsb5pERGEOOv0j7msJX0L/usXv+kWWMZiWt8fTzNv5LWV9/EDwQ13T
6+nOrvsdF/29jpDeaA6EpxPUtg7Vu6tscfAAefmXOCAnfXkjh196oV3cR7aukcSU
Ueb/POSQ+Hgrs4tSfaKjc/9wHoMycETb+dEukPkvH0VVNQy2naoMcW3jFmocP/Zf
jMb/WPYaVnWnxHXZE8TqePLey8tpV0p8/KCvuWn4owVhRtkQRzNvwf8+IjuUL4PV
pRypMq0zEHAdBwqWL6NNJnro+4MTvSF6zoqYSNdqhSJy3g1nHGvuQmXEjIvQh/xt
zrEwypRZDzYqmdNwU8Fo9+yUP8zbIOGHYAEiOCYrjrHeg7+KL7NLHfl9EHXL4GD2
M3Y+0oF21C5uCE/gzV2FO1kbD3YrYjULwzIm8Oje0rREXgRBnwe8ZInNvjJtcagt
TARw14s3+d0RrTfPvp42B3TwtzzRw02zjv7VutDDOXKcd/XRhWPD8+PmQn9KLdSk
vz1aKad8bkcH8qhbZM1Iu2f/KMTUidRwx+IILvRY2VXCTrXMJHN8mKVe478NS62J
LWwQ4TcDtvDDo+T7Unbc0Pl3NcF6nPegYkGf2WHBScYss3Zfh4RIdYpsklNuU4Vw
/qOumqV+hvEQbWOHN0eYrH6sjtBIX5GjIcdS6IxNnDHsKnc5WA1YnNh/1o2oscjF
VgYMVd9J9BngE/autMK8lkmBMfmRvaYKm37i6NpDzYMYwv2ffqtHlJ+011QLXVun
WBqbMSCSTACbhxnPwpPOHW4NveO+Z0B7NDOZIg4IxaA5ez7u3C0Z0PswlF70E7bO
7RpVWAzt5fsJXJcPEip8w+481oYra5qiNDoAko59phaugSmJlyhB6PFZid204lRk
TXFOPAmDk4rNPiYlPIhbXsxdr57/LxgCys+xsneZ/iZ+amjOtLnfGWlwywrcJk6I
v7UXN74FfL7qMJOGTOw0ZVa8wQC8zu1IF1cTVlBVpWQDmrl1n4GhY+vZZkGf7Hq0
stYpTA/mIZi/BMcFnwUEw2/0MkOmmcC5af4dZBgqvLrYLvb7ykk0Xoe4IUbtjugP
ua3eh3+DZzjgYI5e7bG4M93LgknUx76mZyYeSO8xYfTJaKqQfgWPkIEj7v1jdtB1
TveER8IqtkE8e1chnC7m7pscRmqJTpXhw12t1HmNR4sEr9zNYybS1ZxFQo96nGSQ
3aBvUpNpG3bhObTp95qL3Y/19vJnON+8waiy3jkkiPGWD88zj1V9GpkFuvCTpM/W
KkmmJMwT628+fV4Fw3vdbHYBvWQkxygOo18u7N+3X2Hjcx6P88SZZnVjXaAV42sz
l0EV094Rqx8kGQsCJidl/+u2n/q6wupWqVgsqgXkZ3XeLiyPE1+5n82ARJ0rkce1
ZML2uVUuLtEm5s6nISpzu+pl+UAKFaCRy61fZNGKCXaXN4+S94kwOV4cXroHgaOp
DaZyAiaR8floi5geOrhsF+moIj0vNS2ypmABFnQr1qL6+I4eqcyqm2CowBWA876w
nkwk31kayUEQjT4jIiFQZJpHB3pN5eqZcnOJA08vI1AlrH9aiqO8yUNZTCWO6r2f
h/kzSZ/HiEujH0/6mlaRz3+nwiRy4Y8Vdh0edZaXAJUQyvtexO7LFjOx4wyAuHZg
EsWU5+z/Tacl3JWoZOmcPjn8t7NRUZamO0t8PWx3ZyVWKx1TeP80SQxDThQadiEu
JCzsIbPt0LHPRBWl1xXgVGshncGTYJPe5+QNzmEBvWX9/nUUaH2atdDp+qXn2xuR
FQAYZ6wnlCBa+6RTdvYNN2JsXd+qSxdOWLLgXr6ORMIi5zjRMkuE5909vFkwlAjO
5WHE0LzMSGWFeRJQ7YAaPIgDIuovT1SlOE0efQC5YIxg6+RqoVtjqUfmWUZ4QewF
VvowxaksFWKkHiFJZyqkboGMRInHpdKQ6wAJWU6lpYS73x0NHyU9j4F07Nf9Fk+O
Y1KQ1kKXnpIjz5YDTwxy9V3CzfCgqHMqhFFtpPBXLuyE6bF1Y+tRlL8vPylqvW9n
JJIWjwK01jBFbQzk2xG2YJB7IMmPl3BGHJHdXmjMCd+FYm6KW0BGrx+OlOqQYwJn
Ew6aKI2eWmf34artR5gxj7OpBGSudqfn+VIyvZyxqVpkq4WE+WcDKsY/Nxj1148F
8B/sg6TWUm+zrxqRm/k1h3KmlU/axR6qdJnAHEu9b6TiJF+Oeco8DtLuh4WKois8
9PciF4FOuLAQ5uo/YchNupw5aalEWFTcV0kZ2/qYiCZ5KCapI0jTHNNxv4FVNfGm
bRvlGo45MxM+pLNjDL9e4S6xKb+oOnFTSVOnHosmrNur2qn1FbMHpnA2gM6zxGx5
eeAUBj3dvYS+8wiTFO/klID/PPIdpXuJSSKTrIeWguOkF0mtvmUnWpCwoMhSTW9x
SBdXp4EcxD7nIa7xMBZSkr745gs+jvtWznA4IgMdfheYLbJmTZn7pDEoDnNybGN3
M+0U3x+wyA2WBB9XTievdAtwY87BtKrtOBPRFrN8cd8GPk1Nccx6pLfpkkuBSt++
CRtQayMLIoiBqUncUwVjg0+JO9jAw2J6yGmZId1iFybAsGmowA+o11sH8uEme0Tt
ftHNob/zmuSJbrbbr3Gqe8iGmY/+aNdUIZ3uNeulhgd3kzLO/QifWYVyBlmykpUr
Oroie/RebXzd3hWYip18HbwmDgpxTlmk4VgJWN5ZMwf/T1XSUFTdFEx2OHUC/efq
Jy1mJGqSIVUGIPniYFiFNwizR4tIDrL4Qxt0MVUfX8ayg1NIpHmwLuiS0Fe5XFHI
72XazWO8SfNd+yQDYTcng/VvStM5KQssdWHD8Hj3lXzhziRTvXVjsYDIWkEzvxQG
uxVUQub/gYaiMEPxol3ppDLdzVUBhscY4qATceL7AUf+Al+Nh5SCgLPU+g13jhLx
rIehwa/SbwZCW5wKaB74FjzmgZ+QRu8v7Jzu/+cfRrqj1FFS6A1Gw0beTQJ/xSbE
t4vM67eAdMeRGRLg64NS5/WJ/F+ymhGK9cCgVZKa+xl1V6gzeob2tt1kx1uDplFx
u8wphbWKSJeMTpb79vCRCsh3UQ2A0MPeQZ0KWkm/JdbxTsJO6BCrs6yJD4ArdL7z
7UBvwo/7QuVpQo4+jrH5tJ8hpl9j/7Jg/wLT4k0+olCpK86AcVOhrjH7SYqb8gTD
cNkxWePGHZD7L3HU6l6yP6F+W7D640zY8TL5+u7vtFKRB4QyNUNnE8jpPfwP0LDg
xh0XAzz/oHbDTG8deJKlj9f0XCyhAZU73i6uarzmfZ3lAgwhWu2bKqOv2IKmu3eo
Qt4smTlIO4564joMAY1Ys5vUKS10nY3uNCjqSRdt6tNJLg3krtsfkgEx/na2PmpM
pqdMsSoM/Vq190jRDi1029O6nM3UI9/p4bQ7IyvSqNZnZh0j8K2p+h3hw9B4KGPK
4M+nXttyPYoaNcbveQesgvl7stUUpQQLBiJA4gObuC2wxm9sSlniSJ/UO8wbgdPI
/M5ZMYaABug92BWPANP4fko5wzr/f1naN3hBP8GuQsuGldhCHKC0XY7Jg5FxtvXK
A8ntMMzUGLVjDFJEstY4jGIZD+fj1jYWwbsbu+gVTC2uxM2F0L2hJhmlzche00FK
CQT8eiyHYBY5yMC8UkFD9QCMjn4VEP7BP4hVBfc0zGoBjjQnbyGKQuiCo25XHY3T
IrJ4QN0TYZVki46ihC+Nq7xP/TZAkYAvrsYhH/PD9Hwlvq8nYEpx0EiS+fvNrU+c
Ak64fuWkjnqweQbw0JHw2pyxFALwrM4GP9TS521eV50AHxC2VdIljLc6d23gYWOe
zp9SIzk0x4C7mrc8IuNeLcYnpkoEa8mwTuWfEu84hH8U/VX0KW0zn6qf4CxkENbb
JHj0LjuiFBAnnqm38neEgetWKqdjrdp53hngvhqZ6U3quphr2m9ITik+iXmIztKP
s20Ww0CDe1vIbzfuEnFe5zZAPDJ+m5MV8fuT6F9UQhyjssInIjhClmDL0HtZ3UUi
kfYOHoBxUWwgIZdj41bVu8l3t7NSCBN2SHIg4EpLdjCHyx6k/BIQb1Ws7E2HXQZk
XgVLVLDU6i0etzZkFpr4lksvRza8DIelGSmtfazvu0h7K4qkYQ/QtbLHju6+q4Go
xasUmRblBllYyjKN1U449UqWFECVNe36VwmZmXSP/RsRFzP/KWnBikHILFlie0up
BvLFQdZZn8ipW+W6eEjAuROs08eGuSUZyX1tjBeqjUjiJUMFEcKrkZj+uvHjL+5X
KcyhxoD8/5P8HRd51vRm1OxaZBY+C6u0Bt5IgFn/WrqG81EzxHxRh46i0M+hULjf
fUxi97qOlo8EFzc51TFjrJSKcEQgY2KT9pe7tzi59netEK2CpF3NMuF26Rai/dLI
/BbuDdtsa2pfV3fhMNPDux28JApJmaBeavwCRpgE7B5MN8IxHxed6aJJc03DptNX
XOS5KzadjRpgnKkmmmLT7K+graW5Id6ZzndNy/BPf9E61mCJ+TkEg571TQ+vf5mD
D7ppmZCd8A+D5Wk95HtDRBu8EOQ6V00zuRoqqWHWutsD31m6f4K+Soc82hQqtBlB
OAT0gM/E6kTcZjJ5SgtmJUT9Yw+yLs0bFkccw24yCy2frFGPVG9+yXSDZi+H54v9
lAD3JF6VYSqbax/lUutJHZsn3SYJGXEaGskuvEQj5qACenebBYihDgg21c0YNXL9
TkywIaiypRVACpUBswWYHx3f1+o7bOBkrSc/ap2r2R38BPcaqXA0cA/tSyVWQvvQ
225pZvIAPervTDqJBiOYQiIOK6PVIcieekeoMOH68v6U5Cmqa10kR+1KqKLSjLwt
yfhs2KrflvXe8iPjC63aelV52uAiIanqHQjEvjaj/8eNp2kTW/NBTf8nh3iDfkeB
EpeimVu5LPomX53ozwZtvjm7og/07X5W3apqgwXQepG1WQCoVSgVBhsMKOWk8EwK
ClE8Npatw0CBuOWptwvX286wZxdxrts5Zo/khZmKPftH+y3cnLPlSQJfaXLhNjIj
KqRSGMNynHpSYDZIrBvJPUuBS+X7BGaAwgu3puWYkpNrNJ1o+kR7NXYNlP9qk/t9
chfoEBBkVuoohPNkGGRAchM4XSriu23K7Al9vis+LHBVC89rwGsLE9j8ls1DrY3Y
sNtOiL2nHCCHC17Qfs1l4TgJ+RtnyXDvaDUlGNcerKFY0593MoV1q18bgs4wi0we
OgvJpRytZChgMMAP9P40RKk3T6b6B4LjR8XLdjzvvOiNFbI6lThfbSyvD4Uiaq3l
4VXcQjN8CtlnieY7p5HhAq5F7/W9FL4rJ58ecZ6lwdb3g4PmxwFI219CsT/1nFSX
28ic6yPT6dRP22wCrzDG1D/6MozFEcsbcQqvaWDdyO+RVxnfsn1aAXIs1ntkRKpm
RENZmM9Lst1c9cgfITAJNdyFEwZkUotySBO1ltxQ3+WYzCrJSil4majdVngVMSe3
A1eeUK5etKnFybme4OlQe3AoVTTmOa3dyHYC1EsFAotgMOYNyKcTbcgrAJQ3WM7n
FNcaYowj0df4HXvBoLkDG80JNpw2Pv6BuKfKQHy8vG+YTkFZNgYf9wQsQMkoQIgy
1tULcCviULsrYCBmPBZHqwkHTcwTR4Kd8f9RqLQyNIsgzsHIkbvjgmpqYd9O0zOu
5Z/v0/9SJVb9HY/7TtvM+f/8MyQKb1ALoRRpxbSevS8sgUoWGqEfwmtV+MFTAXNF
qLiXmlfqAWVwVWWYYW3FXqDsAe1HyQRpJdBTqIlSFwbWMHoDbUJK+FyVEBZAWna+
3Omke/xF7S9PI8ihwiFwSw3HNWe3bkn/B48F62PzlyeYz37q5XVtWknBHkRAlAnG
7KaqwrWAzFDj1HrVjB7qj4H1CpVql0JAHNSsPlEiPdcQHZzk/em3w2KhArb8wjDm
kkBruYqcIlg3ulkOqS9oojW+Al4Mf+zuuomWGwpFe5c5XcTKWwHuOKvGcJ+2EQDo
dT6QcffOf9qfg/0405UuhE4gaVqEq5WKAf6ke1ZaWf4Ww0QxGz3GOJOEfKk8qrT9
4iRcH14VZh3k7sEgSzcsWrSRAOoXAmw0/yRn3JIrMsvCN/4otQSeHk7uAiq4Pm0M
Zt3nNODuwAfK6yflqWPPECuQmpeAJ0MZOSvGf9NWLnTUsamLul90MrVVlbcHMZYB
slaL26gJV4yyTd1Clh0Q/jTCfkqTplShS+hVhCZpM851bp9zhjApSjPq7BV4xOTP
VPdb25hUsB4wTonl5j4J5dNXM6nIzYpXQ2q+c2+VQb1DiouOOfS5cQn2tZ7B9Wx8
+hUYQDMnqLDnITHKWFXkZSxE3SCcKtjG6nGjWtrf3+4f+3n1rkeGCJPSLggFmHHh
v9fsm7pW0wdLmHO0V0HGBd46AbW4eKPgJYZoKGxYTVWuQOJ5NmU4dLq6+WtOt/8J
BXZ/cDFC5haDJiYntm4XC/AbYLYQHMDh52Lj76NJZlXwpol1ogmQUyHONF++rRO1
WMtxUAg78nCY16KFW0xEt+vIYMjHjSw2HrPusSr3z4cnZv1CYBUuz69VC7/JIWeF
Gvi8ORfidcSInwZk/Sy0PT7x4l/ZdMplZ7tAXdIj+jyViVj/AOSmfiJBl3QvvJAj
pnZGZP/oBhLKmFcUCJ+tMxEt4aKY3Z40nxDcHhV/Ah2yQVrZh/kbFXf7tnI1mlx5
udjhffqQB7gcyTaw5Y+OIJUtaDtk35nZjnTzobgPkjF2rOeJstNTyju76ChPq6dn
PsPLTqvQLvm1Q/WZTyPt/cbLylddHyYiLrJQebLFgqsr0I45z1hFRVSIDweJylDG
IF6WfImLrJ91Qr0+QTyhab+yMNNxlMm6gH2KieexSk+PpapJ3jukk+obr4mpLPXs
2x/lak792MnYU/69eQ6BNADYW9kRR16Cua0ilGZi19ZQ+E2Vs/dsYMrusCYSn8S1
5JVLeiDEa/f22IR42rrtl5Nfn5yPfNd8bPtq7R0pTPVEsHdNacu7TgkFiU+LMm5v
w50try32LQq6zsM7byrG+h4OfS5CPrnql7fj1ygETyh8JuV3cQU9t9SZ4zjFu4a8
a3fOBRJPK2V8hozgJvOD4US4U/SrSOcJGw/VenX6GydH6cwtr4d2SeGvhHhDt/Gu
3i8fuaqVwD2vJw5pPYBF/IX+21cjtu9brwFuS9DVC+3JoN7vW8VHSUjpy2RQIZrn
fjdIlDFqOHA7qRKoQi3WA+PKQzTZ2yLGpRtHqQDBsxK89C5HpId+b+qlnlm5dBhV
6Ml0cA1JC47ewRxFx8oAL67W7b/PwUM4aaye+LYLUIJMhfqDooueSKYVPwTe+a1F
LI5sMX4TrX/ZyNs13wn4Iu0sAalKwxxBPiu71DyYxzw6qUZCmP6fnNzGSo90fefq
gCOlSfYYDrxXRJthGlDJE3/D8Xnsp/ricsmtStAyqe+qKDHyJTiEV+OBIU+087m5
rVnQoHrpa6lvWz7rFHvIcPWsSok3Xoqa8SAl5LNbuHYat7g7dupSjKUpBDnHGtLR
7rbFv5fr0DJHTTU2eRO4ZbD7jR3hu7Yfpv4RLmud7v2ipKdbb6Atjeizm7owXJgK
MIUMF+GHwxpSrQejAqNzQ/R5Hp3l3HjxrDanr16nUeBDwAx1qdeb2exnI52MUnvD
7FgAM+pT5LwK0N4hqjoMvexQ0r2EfBc5o9rYJshql+NYBivyUpD+z/gjYMZQZ1Sy
18RAlN/fbRLtxEftyNr5lBboNgPCay0jzVqHQ4nipJe27s+7sgu0KvAufh/C3MCy
gQhUfVBADWM3l6J2qduPnCDFaA1dbUFrNdak1NntR/MT0uzlN9xhiytfArysinss
iQy9Y8nC3OjE5e4INr0Zb0gmX3ZRlw/z0KVU16eEqKqMfB8MUnfjf44Uof0RIDhQ
io39CDJfVd85NcODb/tCOmTR6/EAosAMUe3JI0l8xcvAxVWPM/UeLEf7jECtMb0V
227Lh3IH6wg1109/2bVe823BTfjThzqKc+IWEDyc6p30X7hjx9uvryiQdw0DCofA
WLLFh/CkOGP96YljjFYsMptGDI9eJILDl+hXCQ4eWZGigfn3SXGPXBs2gz+Vqyfj
ZbF9YU0iltOAKXLCSIX3UK9UXQKmfIOfk55MKpZjkUn7i8sigLxFiwKS9lIzc8xb
J3iZTgaoZ9mzCfjOIAm2kEqU8o0xdhPhIwDsn30ROrCq5fmkC4NT+FB79SKnheTV
qFa8szka304oc23/2dSsU+1mFoxD1kW24SbgHDIzRoeBwOSeJz5lGSja7BKWZ3Hr
23nwcWAtX7+kPdDbeKi9xzr4Tz2uj5xvRjYra+dIlM3009JrU3biv9jbm6inkv8V
l5D4So5eyC1bqVZw/WXQMliNV9nzUtj7szoj/n8jLtwe/kga98k68Zqkxh9yEI51
2mtztUimnV0jSfrTKc2s1l7fYqTyr7vZw4o+32t+Q0OLHfh6MrWUCPADEWwpdlKT
74nTSzbKy13ZrybtZ6z1RhF1nCODfjcY/V79hxC9vU19f9d5JdT+kqlQ6xZb7aNu
TvlXvpCiL/OffUDKequGObF7P0GEGsLAZESTXc4sLyDoswsPh+C7/S6EFzzTTdfC
e09K1TsxPQIak6vW4biDm/bbVanoeJLSH/gZyTID6/iV810T01fqElSiN+Q0D7BX
W8JU4DYQUpkYjCNT8WWzdOteK7rhUp1CEkBwMDBnBuMmXiKV/6w7MnT24cUuXUov
T0kI/IDcN3zIki9agKdcIOz38cFCuzK963BfwYB6RgfLNYVw51vzoYGivj5ax/3v
ukJujXItD03IgwnqrDHnv3Neobwo1ZgdEJCMfhNTmTLy+gf+JthcgYxuIBfkc6X6
4r/ZIScK1xwXKx2hChNdrl+Dn9wHEi6fx4BPhdq2BRrtye2dX5VtyO4YMji2gi2S
+t5p3MrLVFU/1lh31v2MG+OWp+qImwfxallY0dhJU/rgkhCJzXfi9b7SxnemGn/x
O56jv+TYtF7tLlZsSKAnKPRJsCvQ3HvbgKqa33Ln+DOq/h8xn6bbhl4P0W5zYJ8l
T9BQsnxU8HJdrUqZVnQk1gCv6viq4KoaE6yO9w5Mk51+ALWd2LXpblnTs4X8M/L+
rC/+P89wW5EqRMIEDoVqysJAqxR0B4QKTvi++UVi/1CtBLfXmbtCjQm875eCJUsm
n90+ddeUIG9K+fdDBg0mC7JiNl3i4AL+F2LNxtj4e8/ew6Yt9a3lPy1uYIQr66LW
aqyr+wrGoIKHsb97BZixxz7De4ymWjhJp9tkv8uHKW7MAdCJGGborJQ8krAknOSN
JuuoFvBbhb72OxNgTHk1dKwY0Hz7XQt66eNWIQ4E3jESghLVFwfLvzztvFrM9PIP
tnNCq5AK2ZvLV2huQWvGQxCaNQgr3ay0UY2g71B96Wgg33DU4N2yk5S1X1K+n312
lsJ3JSyoroJzT1XWqbT7W+TwnvPeNDkdHk8HdIqa1qVG1fFEC0Q/MLTQiAjf/tL3
pAIYXPT4pBAProWGxOQMRfRfVAtPc+UgNz8QqGpWhHqQVZGo7MAelgksR+DlVFNI
oZgH2fc3ai0dBPS0z7oLk7l9eUMUwITYxq7Hyhizini40em73ORfBFiSUCNwLbDu
vDB73Ly4N4BrH/SczxJCQO+VealF0LP8UL+g+w2hk/aGQRKEaq8iizJ1F1NEU+TX
1jyqvR4Ux53tsNPLfrcxWo8eRIouGr6xvcuqwy2JBi+wdcvgLHEllBvKtGXoKF+K
yos0n4HMJdUe2+NpLzRjTnHsj2EGP9IKX/dBAwN2703Sc12DKHl4L4eQxnD799Sl
ACxrVrdJAzjrEwl7tzd8R/e0Yk48u9h2aBOrszS+wFUUC+UIaJ3q+H4m1ILeI722
KSeU/pf+219122NsbSLZ3OnRq3b661/kTIu+h1Pj5SFSsjg2hzNP8gZ3jCb6lAFB
QJpzoQosmg6lwyVL7AC/VZO1rekl1Xsfl980a0jikxRakG3XPZ4w206xdnoq51Lo
2XxynkAL/L14JkVYRLsTe5esMUmQRYMajplJM9wazCCl/Aqnjcbwe1kYEuGxW/k0
QfH8g5Svn5NOArynnS/mLeudHQc+oKv4aIYIJrN1kJYX1jddeIDlXSzYe5ag1LlJ
OAD3HliXv97vawFS6ykOqlgrwH6Zh/6SkU6bWJpJe/rJ0G1G/5/IlNuf44yY2Y6p
AU0L1wRKUCnvCYSTfe9o8f5HfRdcUBI3K4tCD0uzQ7iD3BoUh8M+Ml+5JeYpakOc
Kvdk/wClKlrxbK+Q0BST6h9O5NPfmRuKt3JuGvcNruN+rSlXBQt8NO9edMbvnjnB
Yq5BJZCG96DcrFvmR2mThbBPcqPi2XRXZLi+qrfa0X0zIycUP+SAzw5DTMseMxbC
pbPBhYhkXYM9Ceo3VyvHKJokjCODhtgqAgE43LzgV09eDgUHRn2zGXg+MMA0lOzZ
Z7fzPDiWjn+sW5975BIyxLe/PamRPFspQpbpLbtys3av1bz+B/Eo4Dn7zEoaZIOg
WlJ+IiIb1QA6LM3+PwA6TAPL6itEjgwJl5VcQKLMCcocZB6ffMZTS0Yp6LIZILfX
ORnB1AAOFkh11QhzWdlNZUlo9hzMnAGKd7MygsRfNftYvAAG+iwxSeo/dNioUwvZ
fir1pJH0wjOXGQC59xlGVEgfeW3ZWjqn1jnYt8LuKTlFF9DpemHwN7vZhAsQ8p+4
OgNuRdz4/tmITCcFOBpOw4aM9ypUsflM/No0xM+HmLSVfltRyaJqzMMYCny9ctuG
6t2pNYzPcoiGjnKFQYL+MjHzSi3bhlseJW+fG9aXkJx9cQW6E3upX/g7WqjuFM24
Pl3V0ocfVdOVWcCmFy3hONTADdkS7opXKmbif/l8UWiM2PkC/1h+0owdW9inZNK0
qC7V5k4Y0jS0cyLGTtBF36dSYpKOuuLStNJjNVc7fNdAS20ROpyAZpAK7f3jTmou
jX7qm2ful63J9Mdm1Gw2X8XsL5wC6oTI7AFzft9X5xWIOtn0DhcdKiMrYU2jzllX
z98TlyEXtKygtvgp83q6CrQyG6QbkftcW3or2vXjHDUBcOJsnZOzkA6KKf6PgJHN
7wjqEfHpWk3NakaJQ7rlhXHwWbSIOr1fPNW20lY0e6uVgg3lIDFArl+6bErrvjCD
9yeV0PHvyPfNEeo3AYhnkG63EmlTjtnGnoKYXgOdgGqSJ7j0dIF5Sns/U4eaFJvQ
umoyfl3LEjWnwdywdzd2iNBRJpTGQ5GJwMFVenFdogt1MrOMA4/ZlZ0F8X2Gf9KE
/HrWp4m1y34uz3PusgE1GuvLVReMqt5xANgAyCgnr0w54OB2rebcomumNOBt65K4
xnN8dgtllNUoS2Qe+LcoFvxXn1Pgb4fexdXlqe4bOr7Yyf3kL4sAmeJiVnzPHBU4
VLOOK29Kb7Qx0+YLm2xuJEU5uoMeW+C88Wh8+sOyPB2DQ7k5b6HREdmcbPelSPkL
Lf8M1jdq6CRraUombWCwnKymd6EceGFZHpZfeTfx7jV8onCMeIl/hrXj/n+EG4Za
tHmCSvJ0TRDxCveymOcCtlMmfM6Y5jgLhxmI07VUsbdd70925Niq8c1KnmnTTMF1
VB0GNWcJXIsaiwbIAEzhA5/JDGUaxxfmvflnjKcdSqNy++1IO4KbWXNhGCvYJCFw
p0R4/ySCSSS4WPfx+kM5eBzFjI0OjMwNZlQQs+woHm3ROuF0uDNx0e4A3tm4dHBV
YRDzZcwVHouZUW4HrVb0DL6o8k2LnSOL6CEgqfKjyTBSua2ZOoGlvBO9kN5uQRpL
enF5DnckOUENxPcx+0J0FBD/kmHZjCA4HqewDH2vyPhjnoNuWeAMoP4Khy8UkN2L
lzhTJyoBqHXsJTQyfH+d6TL7h4K5FIyx9JVm7TO+k3TFVNfdPPRKym6IQUrtSDe6
Tj6kwMYZkX3umBCk7mEJppVfh63xosGev3x1YMPMq/QydV4ax/k8nY7shHQtVF29
ehYNME3KpVfPyCXB6C+axLJawrfOeMgliycYyGt4I4CW0Yq0K0gADBv58k8CJlqV
5M+hmZ7bTiDGIIsPrdY7cYUuXPGzv6RL/dyuy2uxuNFAEia+jsJgf8wXrGHQHa0f
K+hlg45xz+H054t4AZ+nrpAX6oNxZXptTmMeURU2j1WmtYQIpe+3QyERVQHk3zNt
QkwTP49no1Vk5Q14y1Alx+VEAOHeN2wDmGeeQGyp0sENNWkJGlm2TBh6Hix4KiJl
9kDbLcP8U4COgA6L3HSuMzqPr/VaEeau92FPNMWcqTiX2m1Nw5myVf2QMIeY6GYx
kMjNj5P87yamc3peyj5WHu4iGJxmJxIFuQLTwISxogg3qmDWlwKjmE00Z6Zz7gGY
h8BMIZ0WBjePm9pZN8iCWJ69muIXk5WOQaf/IXR0KIdEQ0nmcEE8KBnmdVhulws9
IOhCogbgshrC4+6YytxYeZsBxxp5N/YGbsL4/+r9x3zksMRiOMZIb4PNAS6KMKtK
VVBgr18QOWDK2DiVK4o5tIMxmLgfAOabv/VBW+kZ7XXKc3yZ2wwZ8xseqN8koN5K
hb04iSK2s+Bri4U2cW8turF18YW6Iqv3ocXrxK8okq3E5qAcfRdKXXSNtgLpQFKu
1Twv3NrkMDx1MqxwJBLpfjZVclqUE/zIVO76mIAe7zrM+5JZyrSybyg5g3ZUUOqz
3yr5R62flM/CX4ozwslysA2F9F3Cy1H5ZYVHR4slJQ6OaSxuCy+ujw7ydWhYS9cw
fxQ6gfU2JIPiPnQvWk0IHkOgEVuOkwRu1z+BwscPCNXsXWwck6p79tvHHpG5bZET
ntyoqvIPsyeooYHQTyilWbCT+tWqNzoDIKhZXtRs4vn799+y7NVUCi88EjTbFd1P
T90VaPLMV9Q5mC5snq9z0jPuPgdXqhcdlO5u8uphlgXAe1zQqvJsE6qauY7gyaYT
PZfMuMIICdqcJBC27/OhMmU2xIl7yLOnA0fdRZ51S5/rFl9mAzBVp4XWKezZijSU
SWvq5Z1NpDf3F0K05LB9oCx4mzX+iqNk/HD6r/tL+z/uTvf/GyZxcsJl7HDgW+Ks
qqTnYJvdy61bYT2gRtNLJ0KeUPyi+SJQsGL+lCMnDYXWUUAJyioeyarQTcM2U83T
5Q5bN4lpuvPZl3K6lfdH4rKyZYoAR7jlgONrvUYL7tYuQtrButY5ets4LYea31Vt
VF2BGS7pm4N7HX6UaKj+nvdC7+Tc/5QVqzE8Lbs6PP9fCqvBQm7Y2+t9JesMdsYI
7zH9ZnB62YIcNUBQ3SFfCRsXKGH0Pr17sxrR2O0/exzQ1IqSJs6Tg39KGGFrtIRH
yiy4fzZCvjiJniEMj5z5766grxTc7l5CGBqzd8yj+nGKinW0oWf/SVK1VIRua8v8
ceAUxQHfLn2f9rK9d7/4xipl/Jebh6dN73yD4JATlWXLiKmbgR7GfH6jMTcXLkkm
CsgqfufOPmA+2du9uCe5xLAVRQ6tEC+XCc7ki3eEUSj4EW3t5kLXHKxUgFeO4wZb
6jRD3E5RHRN+I/z0Sv/t5dwzGtL+esEzA39JiZL/rcOm9xl4AM6kg4oi0FmKM+N2
mk/vsfG1XWuwlVD0CVlXNlaXHr+9Z9O0Cxc2+6X4tnOYMfLs49033c6cpIuEj1po
AcwcpWxesvSfD+zD7do9oAXd/qDRqPJI6A5lunA1d4XKnTS5zmPZOpqTKI3PfIXn
tf86JYmdPeLbE+r3Qom24beSnP8d0VDVmXMJRF9f+OCcZLlF2a+JMBLwdTVar2MN
Orj2HYHQHyLqeNq/8CvxMOw/ZQGXg5X5GQeD62MjEMg8SZUfwjenJvTbPE/H1ghS
8dyB2Fgzk/xHhRxTlXsoE5xK4ImRhlW6gOOkV2k5KyFYJiNsofEIjuw8Le8V02kf
jeVhPSav7zBUakPIwDGSQfPat9TeHG+BgXuQR8eZ+vvVXZBg1680sxHOwjhEtNhK
73suVDAVLbMfdANpu2Dc9WH/ghhzu+ww4U4wWMtOolNT1+trZZPCerCN6+C+Zqq4
KxP60V5lhiLED1vJ/DzLlH2ONnKC1pDhBSP2YgCJj467XPi6SraDhHtZBkDO1z8x
jr0evbmmbwLRXqYQ2Cg4oeVSLz1KZKMGO8BCpPhU5tD+m5XwuMfYeq8PWG5+IVsu
xWNXGx2ggksHhUpbmLgrmBy2MIPuK26d0i7k44/gzHNccQT8dRjcoksOBqDg5Hw6
0Ij0uG3IvuhqbY4UOzanD85Nk+rM6G7sQGvoXmFtYSWWZ26AkPuQFfwI2ZwYCbHl
PNFlWbaOa1OgKg5Ra9a9FpV+2S+lIQuMrgII9CXX27Bh2xT3SdtZ/EXnKAZ2SFX7
5Tp15lK3tABLEIM6LN9L8WLSjOh37+azJbPCjlIdlyVabvLdeQXg9xVhFb3P1uol
yFhns8qAqJZ1/pELS0zwqYJYAgA1GxBAKJO2vQmhDAy8PFtVKZfC7MectmcfuW5z
mPBLpujP/Pv5aeUL02T8zZExwvi3bwnXI7bA+ZMIUSlaBRb94PG+45mOMdr9Tevv
O7aZMH1kCABrYs8H21Y0DyboFTZ2mBt/EhJBGufc07mqxJb0PgAfmX1cxCbvxx+o
XDulaUZ7JilfNcO+XQ7goO7miH5/x5yYRbaELMDZMQuDMltjMDrUxPHbrwd38Zj+
awwPv9N3+cwVVeQJnVxwBTx+Bvuk0cg4PkElerX0XM87RqmQYzHNhpB0ES+J+y2V
lm4dfoA3aHdBhnShHRSb2ejlTXpjz/V+IiBbRqasvpFt34SKi6L2zrTwXt1WmI9b
O3kcoeRybQKXbYw1TQyFp/ZMTEzCpDNmFJP4hcrcq3B53RAa1CqIoT9rYukVzXMx
mp7SJWTCQbYQn0X7eoPqfpxyH/Txf+ZLRowrfhpnD2iDtETk4YNVsOlUxTDPBkC8
E8U70G/Hy0IG7fdht9dOCko+RUOeXWPhwrjLIh+COZZUIaJDwLED1bx+0iU6txV7
1gtPhNa0HZSBfPXzOyREOLFzo2Ocov8AxwlyPobWCpDxPA4Ns5TnV/omrLQ5zdLm
0aJt/UfjgsRkVixaDpz2bTt5F2md9N4XxIbofT24P/2xOlsyakCBdJL/+AiU8lfZ
mOnaBWJqOZnq7S86jRc7yv2bIYMvvktfQ9H6oAUj6m0fb5JXiHVB8LOAJPH0QBII
smUqkQCoMboOCDu4y8n80fcVRIJSsgJJGzpXIjP942E65EoRlShv93Fs1kmMa8Oe
Ri9nttSuMQDlnW9NBU9R9AdvMijuTF/rvAcMj5fEYegeOtxklpTJHEVArM5xka2E
EzDmRwGCOLXwmqYmWKfMMDZ9G0ScMCbRAm3OVua3fNmNcOt5YSGb9v9oVHwFdu/a
NBNlo3UDsuQmBG2n6BNhitgqpxAQC8wJ4ejRDU6vvpHRhlyEBxYH26iiIjVAdjDw
LnIdsQYEeQqq5GkQXxqxFo44itIiLHRf821V1NbISC/RlhVx/fF3RmzY8A8M6oCv
FHpPwqzqgBi7XKKjQhzqzpDex62ZNSzKvLcwBOqLRR5mce5/zeeT8bw7Y9sLnV+O
k0Nw46/UouF3110v/iF4AslDPEmo9PSn641gkvzAN7+unKnY6OpzKlJD1sEegJRr
mXshNNc0uIjhJTTyk4vHjLgztOaUwUfbGymMGipAp2cKktV7pPBr/W2/qfcPljxJ
uW3Nj64mZVa+DkwUZQbmTFU5Rz5AYe6HD92W86uB15y15ctJYmKyJX76tKjxoEc2
og++krOTrgdO9775MdfdafZEQP+dL8fxejIkwXNvMwvLhD2h2CqzelD/TRCTYVeK
5QSADftaDdyykzx30SyFievHA1h5wX1GZpvqUFm3+nztHWALRaIaUuT1yLdDlGRE
WxBsHwjVyuNsdyUJRKahdJMDrjkCjwq6EcR6L6vwkDNdhbx0UJfhdqedXLYWW+QY
hslIJB4qYuwEXAg7qrMHcC6ZzZ8jMXF7e2totAFUtA1RU5RGV+i/oWcY8rIvmaFx
XmT43jVeoRnzTsTyrBKJpCEMzbyezwgl6RAL1AH4vsQhW1Fl3oCUErLCTLxKCgq4
qV/SfJCY6WaY4onD2YzYp48iYkh2mZ7Eup2q3NPdH4BM26TC2WcpSDtuZvij3DHC
jH2bBsSbA4gJt1JZV/XGuTrm+NgIGMFqh3RnycBweN3h8KTj/haiBwCoy0pqjT39
K30HGLDbSbyuLsxqdxN4Hlhj/e8A1QsA4RmB7xrh+BXoBdspqaSarp9dha6YKWH0
9eMtXXYqjN46TalHeQWPxemlb81qXryXd+APy4ELEtFPWyrT9cWLfAbTqj96RXeB
tqaWbPBFAPTMbg1esDNlVA9OkzPPPqzICg9IKVFgLmisTzFc8ALMF6Uc4oCjCmGr
3CIfgKfYDgGg1kbIoaCOLj4a7CbRlpAjwZHV47hB1UP05ArgeHKoE6F86JpOGAPS
RJA7Gt6hi727bxBYTVU4L+AImpJ7nOjMNHpDqWzLGvzoczNNY0DZeKRVflsatg1w
Lsu8JgomRM/lqiQe7DANN6HdnWuCRq3FdynfZ9/4Xbh0oVX41RAsyU2LrgijN3QY
6/JkNC3Y2WPdOgxzwTg9derUgjDkLlgXwxnv0g2o0UxTSl6vqj6sOWhKA5EN7LAd
v+ZHt4+H7ZCqJt2wsbwUcErBryZBjyU5skgPWM3OXEcYV8eWIlBH0RXuRkQYf8z1
xiwIWVCjx4vZs03qasVLkLrso/oPvxoYJp1wQPgW9649LsD3HDhDOLgVENq2MGtN
WE/Nt7CuCqHFr/htWKV84TPPHfmHgQlwRrTZq3uEOjDPo364urabr2bHq7xgjjDG
XeLrBZHli4I9A+3sklt9JtsfIQW6PMxcAxsytTDOcuKMtAryH/rr080CEaAKjAbK
/n39Hr6kGkw+Lk2OrdGtD/k5Si6Jm2aK6tzYA8OLZYOtb1F71H5Z3mCdf5wvpQmP
heLUfSdzTSFQNHd5ZdtnnAeSxvfqFVdwWMHUlN+oJf99ynGU6M19TNWcY9XykeE8
cvH5rvYBFUzrMf6TODsIVYNKz65DUuVXV/EM25HOCMJKfaS5sWbMouMINFYYaQj3
dvqdEMliT7IuXxR2dZKDRCaTiLBZPvL1KJQH2C90bkMT+i/xFER7gFGHdT6JUFiW
VvtHVSFNJIvOIknSVl4dVXWZu+rGENUwhJn31osynQQTqu9OKQWvbbroVJZiMl89
ms84rmOXrFwn09c1xnMgt5wUlM9eU+8Mf7wxJPUf09NbXiRGsEt6a6QYxqPACXei
/9EXG987G99ucol4RqgbAsdIvraoyxyL4TV9uY5P6DbU/iygfXyfPe3xcSkmWy7C
9SlFaRl5U3ubWl3Clm19ndXzXPt2gXPNhSTeWaF1gFrZlCs/DeSznb/SZG4i0HWn
gTP2BuPZUdJ74TWvafQqLgnygMTMzxfIc35S5PxHuoAcWB54b4yTlxMXJpNwvBVY
18LsPILGSU3pKGVGSRfWeBjuhzer357lc+KHh9WFJ1ds4Z5kmrVZ5W92pr8LRbdx
xLHBF/Bu3UVG2guS/YrwINBnaAIu3EPQGvHdVlc/Ex45gexHyFKE/mMrp5kVkiSz
G+neqggOu5kjGR046f5p5xDimAKEtT+ODf9SvOLHVQGN778EjayKyqLTlq0Ow81x
7JxYVBa1cpmSqN34cuVBCqStQ+1+mEI8w2jVPn/bd6lsnWvsgu+FvKTznedDFyJ5
zP09Tv6mtz474WcU6ZLeLH4IDTOZ8KS8Eu3/D53F3b+X22DRLS7z8PiQTUvvdVn6
4k6ZkM9C/eX1zyl+AeA07DwHTnYP00udYXJOS6Ymzt1bX99z6zyEcIGaI1uEl4Wr
5M7uSoIRlgMjYquAZZTzN+d+W45w0YBbf9hStthm+OUWC6MKMvqyTvGX5E70UVbg
mD8I6zac2u6xXT8yR2Sv/dkKppOaGbZYir0r394dKdMfbxjk+ktrJX11mHeSdMHM
ufjnnSvbArshjY3B2YmwqtlT+VO9YHMQnQ83EcsMVhwDR0K/O6nTw2uvxNeJ8cIx
3PxWXRcbiawwpJ56uOZ5ogCP6py7DHUtGNHm71MzpuGxSdPPWNiCc09BDjXYWlYM
9E0MSxEaM4m0TYcQ6/4MjdML6ZTxb7rkqrhsHV+b0+X8wiF49U4FoYNxIx+IYapN
AfQi876Ikw9ODmeZ+3x87XIEx+d9/YdONRV3ZGkx5eKaRsUOHjPXHqhYih6t8Tkk
X+m6hE13zuxLAKYnsIP6yC9OhHQsCalzPbn8WK/kvefPLcWRLj+bmDRp26H1tAAf
yBa9QQMeRYizsuaMiHa7kU86jnT+UDrmrp03aiFuIbQ6qc9K7Lf5uhwxFNYf/RfF
oMkNpoUDNgwSc90OtFk714AiD1hYxLsWQmR/tl9cMq7NTDEq8xscKtEAz7SQx17h
nmDmuEvfvJzvYqEFVK5r95+eGkWAI2xmBvFfZPKSjWmTV0/inHDQn5LK15pptQ7Z
b23VU9B5Lk8VTa5gxviE4kW3WH0OMzeKUxotw0QoDDPylnSGD+iIGe3Nzl9Swpz6
7Vf29HLRaoGZhjPvQZFukrCj3l/cegeRQTc4kxPfFbhFZOWSTk+yZrV5dCSqfxAv
BCkneffnuJBKEfa7b9cLQ+69Iy7FuDQAl2iPYcVK+afxsMSCmJlO3PADRGo/Gq/g
gczFTHpV33UzkTCg69reIcYwYh5KXNb2h+dVE7YzU+0kOaZR38cP9BObCwQ2dmS2
tnUOIo9hvNFEUU37T+ssAK1dxrPxcciS5mQAhJs9CxljyHqYdJNZVEhzKuf2hkfJ
heR1Y32p2J4pV8yiKebWBYbjUeb63fiU1h2Yo6Ucyn28J3BTOWvfulthDvNlvOZ1
pEfbV8kWhULJyfM/1X6P7utgNDurBtdg0XCmEt6ceFP/ckPglgG76enIrUusqyfy
KIM1wcCOWFOjXacw8fZqxelseS4NnmjGKOtJljgfD4LP0nltJ1mUvo/dQPKlQov2
hqreyczVA7Mr7pvDkSoXDv/ulNvqxGbkNWPCRubW6d8cZYUMHQ6YqCkV6AwZJY0T
hXXpXMarCw3OuysBHUuc5q2q+G3BtcIBKl6LZFp2J8dJtmkBVLIC7XQsYAiv/gcw
qOQm3IyvtpGHSuWN7ESMn5PgyIzJCMVkHCCWiHrV3LW7NSq3vGsonK4YKlNCQI+e
F8LTWQOuJ0/NM4pDVxZaLCTMB440IRqE9qr9llkOioex557gCpd9kboUTQ8WsHad
rVQLeLBIzEny+ElEdT3UROakk/4HXRbBjeZQLiYLdUFGT22jAnIo3hv3x+pcvJ92
7D7uQTl69p1KULQgxxTMyCbTWD1hEIROhEbue1X2KNFe4S7tQXHUT2ha/4/eEAuz
5/aTuNaZxGtKhUsSd/M9NA4AP/SJRPR01nDa1v7+u2ZiUwJ3XKXTg+JxImv4+JhA
AtjkQhalbxMeV/iEK8TcrKllTs/jXhaAHcLUCvBwy5DjL6pzwKsbtgf2AGHnkjAA
/CJ/PpHsJ7M0pE8WyAXbuIZmAsRBeoA/m7wCKd8qyLtf7OFhxhhu3WEFrK30inHC
oWpidEVJg/iMqfC9oC6cL3n+IGh80xS7j3J4eSGuauIocahroarb+MxL1/6WMyKP
nQkX29FSs3LCXndYjuciUuEBvFQAr2Py1+Ec5Lhyfbu+OubNmiSG/o0nRbmR86jF
quGUpLeCl3VZRs8ywSX/DBwnXvqZh5Vc0+I/5nkQ3G+JMiZD3a55KQAV3g8bc5RK
ozo/5fM1QmJuFi+E/xaUc34tabZWBLMILhY1nrfY0wudH+i8nyAB+sH19BXcHbPM
aUIY2DiykK7eZMX35fgpvPACsdfMPbMmf2wLKeA9nRTlw8GcqszxSQChyUnH6WaR
ox+wtbwFEt5G94UJrl0aCg/JJaE4MncXWrfj089EnkEUJMTA988diqDrbQgbBSLn
U2wOYGKVot//mRTI3BG53sC818RufY99LTtcmL+cvEm5MRj7Y73tOsJodPURJFFN
wvDRInMBdsbqF8XRSkVH4lPcuwfjyRXBdNNGQFiOL0qacmoxbx0Ocyq2wEto7LbV
mT7E4lrwsfuqimX02u2meBW9ocGYi+jnG2akmKeTou0zgy+rPBaXTmiXmgGCjDXH
FKoIY6MLxU0E9ydhQPsZaxGz0Va6Bf2cq6ZGfVWsw6tzLJZIJEhreFZ2AflrbppM
mZi97TRDV9Kp4hsA2uZ47KMayvai9bRYnSDO1WYTAq53KWj1uf2+hs6JGzGb5a60
zDgFumiQmQn+8iFV2ZcHurqlauh+lQyvqBkaeAXNjMSB0NOg9DEPcxeuksDUODNU
UYTo0DB2DxKKVWZWoGiKRVXcK77784SgrB1nf8h2jXuzUMG3Lz3KkS1KDrPTc5KM
jQGBiEsc4cyNjhVicLDffYZU4aimmmFw6ZJG48b9XGiFljERfF3LuOkzJOHc+jkk
sR1+/RNAcnCOxMlS2BVn7Y6aYmQ2TQApq3h+Rb/vz08RiDEQIowbx/IAhK5/Zxs1
eMR6Xpvpm/Vax2k0tgWsEGivlU7THzYLtIoNQu926S6ZIsW+DKIrh4f8oJSPK+0V
fF8ziMWg5XJWMA0oySvlWoBPIHjD64FfJyXJAuRLuGRqe+lwaSdI5m1SVCz3r86H
y4YoDREkEXOisvq7Oniwkxnz/O4Z+7Mcnm0hcclrmVz7cMxnfFE97+u+3aDDDNUL
L9IHh2QMKXD8oyONkx6Mwy5wgvcbhi8FlxG/QMtM0zIKmmss2lyJH7t3o2MpUtZ9
Dez6Gr1qXwVBo6JKcEJ9AcLMIKsyMGAWt3YZYtL+KKLY6cLQH8UibFDhGwauL9RC
TfOC095EcoAuymyYu/EF9nWULtchqR5/EPs4wR3kctNs2Uz43VMk0tCf5UQo1b+l
r9cr608I7T48CmO7YkABiMz5WlotTO91gShACRhuWs7we/MkfebkPfbqkTQIFW1l
yo9QSVwmA3SgXuchzZYVDtJl3E9k+RM36wFn96fxRjHSGOrQRsEZLLIEcUejsZE7
J2tNmbLN/vdnkjSYSoEOXQCLNVamdK4rlb3Ecml+8hA4EEM15qp5ze0upVQVT5U2
5f5nz8ng5smWhLlYXvY6ZGUlSpGpN79ZGyJzNStm4BuGOZFu/fBCNXrr+bNZDlx/
FesoaSrC+QmpJQVNVFi8gWhsnVmMxqibgKd4hC5ZSmp0CcdTOKi9eZYqMmCHH4MX
Ulz4ztQcCmyrmp4ecatoHKF6mRVNG5UwUdSZrYHkYG7N4TS/A06lsdoYXBmqu/k5
1hMTOC/dbfXEYFv2GkcPrkaUwd0HSietn6jAKN/97pIAlAAt8t2p4adTmHZYZ+se
8Pto3GzKIXJa+LtfgYiHjPpgsXpypGv9oqqxzXugfIxSQHlViwD6BdxZQyYHagzk
POUbgWF9Y+k8yU095O9zR+jT8APShVqsWEkXigBxuLKIe5BiaIvLLW3ejFGYQdiX
vTYUH5rE1TMhS2U+8S51u+bmZRxcVLuLlZSpzaDTYKT6lwhsCyHn2kczEO70aAeQ
kQn1JfkGgAyP5VOq7VRgH7VTzOUnKd7K8IlU5uB1rkgQXnD+hHcRb1sK+xATEvCl
jQbhefr8gfxQPayP+MdxZyRCtLOEf8Bw8bG/elfCSTqqdQHVre59Cyj3jGUnVDsA
YiMPRtvfqb/V/DrT8PckEdVYI2G4KV90cI8kVswXMAZzEbCNiwug2qC+0+wwhGDW
DEI6ejs0GSiSCp6Lv9DNSx9a121bww9p0OgfTb9LdWCS/s9rgyug25Nk6uyvmkyW
`protect END_PROTECTED
