`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A4QLvWkIZSlFDCSQIx75gTirRbOn+gqf509jFliZIwrajAaTqcoCEO5NqmJmSF/C
bjzf583FGl56SWW2H3ohKH/49mZdstAvyN29MjGEr91mWGbeKK95m3uv9CQfzfyK
eeyJ+gp7NdsQg6gADbhXwMEuoZCd1oG87USrEb6L033mloZmKJZ1VT/pRizBg6/E
cK/alh19JCMQNAdcagGEsYDliKyYxBpSO2UK1whfJLXDMPYNPP0PtqxPxdGMvshK
AIGdLtEloFyci0IMPK3M0i80x6F4EM2rvIIqV8oS6HAGYEJP7whB4D/3dyhN/SCJ
24JPydzIUrnW7EpV395sDpQGSOUwR1wdj+oqezAl63j6d4/ek6tyqtnAGWNhsj0L
3q7VjV3N9Q3Km4sOhmvAbQnqD9dC9gIrOCQwCY51wKi2/b469SKfY0jzHfgLVnBO
UHUmYukoQuk5uNC3ItNOACx5EJCyH185ptjDsmo10io=
`protect END_PROTECTED
