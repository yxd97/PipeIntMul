`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDJ/Ot8nNFnglkSIDIOXVycGRGE9I/xgKKNNUSgCg5o4d1+yU17tNUCrPqxnC0p2
vHOlAJDK16fnxdmR0JzavZg9cm/YN1vq9v1I49geYJgt3McRQ6+Hz8ozwz8TeqML
o3T0e5hdnXXTBW9GFk2Dj8LcgRDxS17IG9shsbeazsjNgjK0m3GxzypDddSid7uC
CPJ4hLBIpqK1a4SHwlAQhrI/5MJV/yf2VHgNBeDQijTym8InuemuheJGD31IpGMR
58nx8V9lUhF16UU8/UPUURT1UFxagMmpt3SENDYfvJjZ2yFb3pPZ2OKn6t3zLQcM
gEMpD/qxyZ8gTeJ4zIyEBmMs5vRil9WRak5zANNxjpve38K054AyyyG830glCNkC
vufVoD48o2nmHMYBds+KnejdH18pBN2Qjq/2YyPBw2wzp9kwWK6sVl0kgMI2gP9J
2wE/A4SdAWxuERpJqwz1hH3VRvr1nzJ/avgTcikytJ8HYxU0/G3thYSvp/DwYVBk
9Ugt4Vx7UPSyr/9v32IZbykNOclSix7FNg0/CoC+S36zmDxzQZu5jqrXRM/hq/hR
AI6/s5OT+XnRNWrFfa7SqVPRi0WDqF7icKnFID4UVYi6VuKerNFOFHFfCzL9GPWP
eeYGX3CPy4AXXzgq+g3X4bt2muNzbuksttYvbP65Do0=
`protect END_PROTECTED
