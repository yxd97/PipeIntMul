`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wX067b5beLCCOVqNfOJDz7DPLnnXF0n6+lxTrxAbH85uS5XZiNn93mH/oFQmi5bO
opkln3wrioR0RLaFx0aVJzIWdMX2sti6ObyzpjJZ3rnol57SLJgTUW5zPTfqIKAl
1ZnfNkEXmE6h29BUbE9LQemfMqDS5QnvRh7ASQzy4csxeglhHMLdmKhud649nJWk
Cuch0tQdbRuO8B8snEXJiu6NlFktH9uECZTXCyXh/IF9GYnG9G57h1KmMTNHVwNo
k6XRLeEsrrJh0S4eegA3cD5cWDgtOeZzHhIMBusJL1N/fQ3VisLJzdf143AqRfXw
JhoFplkWrxQzRtheJPWr1WdbvkPk7a6JbObRepa0hcPUx1p8pLhawdDO8XsHaDUV
6ATBAPbexPc4eXdPx367ey1MdbP6uGDeZrW4OK8oUQV2mRwmQhAigCWR1IY8A4dh
41ZtQrf+A28iIuYzxczZH8LS5G64zEKoL2gS6gk8MhrHxCGalKZeVXetdn2fwckC
`protect END_PROTECTED
