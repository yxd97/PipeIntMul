`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EyYIucVqVgTZxA7v0zbIMnHn47lAO+VZg7U1+zO9w+Qwa/YSz8zs6MxTlCh3KQMJ
6IZ8dJo2xDgtU00lNzondqMXmhFuvgq22YCYg1AmbTxd+ZtCVLO4LrnCzoQCYLvg
GWeTFmTqgHbiD5ynDmM20sOAZY/47sGIhXZ3btttaK3/oA3TSvLjcJ/ZBR+0l8t6
kZCExvJ95FIOfZRO95iXqsOT3rEPDaHGtAMtNQtVKr621fv8ypBI62o/InpaygHE
OEa8gIqNV2QTQ0Rnd0yV6MHTERV9DJnEMh4wWxLexocRLbKDp8HqMnsDH4jOBtQh
AecAsh7oWtPeExB1kmoJ7A==
`protect END_PROTECTED
