`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rH6I7LJP9XYGT/dVC7JbPOSIVrjDv6w2TdZEpMFWYs9tjeXJ3HAvZ8mq7sS6HO6f
D3T/PlQ57qx1CQMsdvZdJWq/aVy5+TVzmUavwyUmqfymnfl+2GSJlyXAKtb4k+Fo
S1541bj5+PX5lAjQW2HZsUFV5xssuf+cIIxpnKHeA7ET47UZwkXrATeYf2nsVOGm
55gAqLh4MVSRlyW3ERJKpedmG0x//l6azTb7Luo9/hxsiYKdl48g3vMuw+gMUSs9
/xgpOlYUysYHLJpUiGiydwLHz5tRC69pBlVbp2SCfZVtYnTX9To/xnWG/glE7qQo
7QiNKglHbZAVInzU63mGBQ==
`protect END_PROTECTED
