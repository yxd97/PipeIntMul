`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oRQPN8vMCDI7OwWgsHIsKqvXQogu8bqqrxWi2f1AR3Yza0eNVMj82a2IhK/bV41z
JtoforXzbgK3T3lwa1GOWqr4/2KWrCXuLDa8TNHHNhAYyt3NQqaLFiVsIZ4t0bm7
aH72yIEBCTNrdvvFpMYrK7Ony0blYpugmO2sLsBxEoB2lKWWnrTIekIQAViyFv9S
6CcwSi3oWgaHmP922IhTmmqChTa+IOCCDWT7cfTW8na1UWaAuWCPpxhhIlWYsecs
/lp7O/+EoNVCvuCpyBbNKxlDbjc3mGKCIoUrxXgdm/9RdyBFyKSG5yFSPBlORXL2
Qrg6w0r04rWWy2V93oBpDLjmGHuDrlKMirJfAQ0JK6OY4Z7KcPrz48BMz8gzYUOL
seppkTSIwvDRe3hxWYTR/wq2r2R111F1w13niB7xe/Y+EA+PfJH1QwYTMMCJxtgD
uPtrUNZTwWl9EC7bQSOP/pBkZfAvI14UBolTnFZ2Hg4GevibV2EfifK2KUxWIojp
bgrMTnrqX7kNCcmN03gPcO9OwVGrXiGUFitza0BBrfkg+Q5fVA3TZadC1O9QZSCa
wpa6XI+/MXD6PBg4/hLr5A==
`protect END_PROTECTED
