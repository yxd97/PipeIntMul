`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxQhsjGotHs0go804zE2qtWEA1Qp5q90vx9V7oEhIqzuqSNHgGP+da/Q1KP/d8RJ
/ji5GhkWG1HhDNwhmBNTBHoi3qNkVB/4QHcRV0CeKnTTxqr7EkZPXiCYezNIgV4M
Y4kCSMUAXhujwt8ObFSTGrHGwoMdI+usOVgto2QmXOImCLg8K9aHRvXSMNsiKRSf
wZQi19r48I6stD5m20ctIYgq2+86XoKPpm01Roe6ikfbRQFrfB45BYQ01PHNyiTR
jSCKdg4dm5Uj5o0CucNS+wAWl7PUYdWN9w5u+SeQz0cEJHefAej5t5ZZuBVXXvax
hsWRPdy+S5sAfBCDHT8rYUhfeF5wWlERSLHasAgn+jpHTjhzXfruNHbN0rODxLK7
8tKA2n6DGUM/DPaxfushH/YAKf9jQ+kekGKWK9MeBVxu65t4VrDHgePv7bzfrRu+
5BocqyGaUDccvBmq5b/VTAZMQOqhP5TivRKy8oBfGbrlXvspSim7IFSo2TjBs74z
ixJYZfRAYikUHxJCPZ7hm5Ft+F3AphwPEyD6mFL92BQ3Af7iwJuyS+6Lj0zatMxw
XIkRyZ8ptUt5QMjxxp7rt0gUSqPSs7GuDGrakUGoIMg=
`protect END_PROTECTED
