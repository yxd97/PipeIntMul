`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63aQtXZ8Mn9SHhvG9aK5zilHZW/BXhhlcHUdVJmV9nLLmtJqBJFJsI40LjIwN+kW
rKLmNHt/mYsLlklm2xEfCvaRU17n/Mu6oxXU82xXQ6lHInXlUL1Z0jXopiCwaLvz
CKGAYaqmdf1kYP+1GNflLNsVtkhHp6de+YKTLMMiGTWoXfdOzh0ftrRKO6qLEwhW
E/8GZu89SthLOn3clUcT3lWpQ4F5sPTqMkhfZb6BwNssP+93DGLBe11PXzei//iM
U1x5zhdkcbI58gqtm6rmNH/tNfsYlBfxNZ1tzhllULx9Ahnz0LE2sdFHRAx0BVqI
VHyxznmuQdeGBYsLjqiHMsJeRxsRZlOT4x9nTAgnLEdJVmehFEMCReNyJQHF0BFa
dmJPyQxqlQF1DtqR5GEGW/fZkByTOZU2OSifDcTNAH44I37ljY7l+JNGi+k/neX9
qaWUyjkoAkktG38Vt54djD5Q6W2ie9hRKLlZx8FyRFtZDIKxIZ0xO7mCzrYEzVUG
2dDKzK5h0xNZmsJ16Q+F8ZHqUPZ1DUdBQj22Q32v5h1bUZTBe4o1FUa5KQJAS28Z
YEXpI0Ied0w8Um4WLDHsKJ0fp2WpezuFe52K24mlomOark/VKv8woERwdN2J5+Gr
O1n5BtW8H1zbMOYE8v1TA4wNTtGhRNUoa7oWRveK6mdIbi/zwiA6uG42EBYtYjzq
MP8aoQ/lvcH0UHUD750FfUTNRpnycj86IOEMFBdZkd403g2IC7xzwi4uTPhSZLFc
i4krDzS6hB97LXiJKrEGF7Yfbq/tQ2Igq7b0UCSgJJODaLyJGnNwHnDJZhukSlIf
i0g0wOQ722r4WEKdU/oHWXHygfbU+CX9bSoPHpF0spGk4c4JcCM3jFkz8SurRM+c
eNfZvGyhVdHof8adWGVsy3fYs775FIjlwtynKcBq2uo1nmchXef2D+Mft0n3peX+
cDsfwiQxUUiFMP3M0/59uU53+r2/0xEl4kXHDLFIeMEmiA4BraHoHvDSNteNojYT
n8WWVKYT9v8CV+clhfyVEolNtCshsxiiNUz4mw+7E1u1K62HivwYydW+fKoZhxFn
R3/x40SGzMlgpzf0PSvftFO7BRw9I/f5QGNU2cC/MjFH9jMcFll8ymfpYsKkb95G
YG6GbFB79IVtQOiZXYrAkK9SFUaAm3rlkArRrDv/9vLe21QY5i627ForDzoNS2oz
wDrx636UmhYbXT2Fzws+tqeNg+pLBgnY7sxpjAUnbS5Pf9DpPF16P89SOo8SB2pc
hiIdEMMI2M5e+q4c1cw391c+C+f12V/xr2vPNvvXtfmLttcmL+Y9D3lswnYCF6eT
CEmAvcLyAAiEzLBLEoW73ohXbDr0EQux16/0fTZsqTr1zg7o4cWyLSi/IroZta+q
nKyPIO7sDFu1ayhgQV5AnJWGUoe8nzFDP+efg/Dr6kxbl5Z/MLuUZHvQl7Ke/fhe
yFvJ1E07UsRWH1Fd8hYBYti2JujgN9VSumwoXKuKTyP9Z4L+9DGD0x0t7uaX6B+h
rbHzLspTIIDUCj0YX8zHl+jAtmltMyTmsrD4CsEojb+2BKZpxH2d3k4hpVKbbJau
hDpZDi0gjRMcGd4vRJPKvxHl0NfCPVhQF2tO7nC9/qnKPWdaumTX28R+NbW1g46Q
LoEZJL8no8HLdnZ9JEmnK1oXJphKXh9WH77up65aLeYnDlB2PlXdFlf9rIfWAuoG
2TCb8DMYI2753z5It+dnJQ870Xl2Wtp929oxXudsB7OT2CVvyt4dElCEwxadLmsa
Y4BSwCSjHe/OpH7un2suNZrRwhseQviNgxAiJiHYRh30NdPjW/m6qVxaQdum5kx2
+NvJdcIY29aF3YGDmgqG+aavm8EUqYREBHE2A2XzLRb8NzaeDAqddtcq2XOFRmI+
g5fFmk7FL0dxp/9MZ/XKcNQOUY9R0wOhY9037gqRAH5nHKEkLWXTTg0lYzPB/AXN
`protect END_PROTECTED
