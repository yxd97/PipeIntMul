`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t05QuaLpqbVHwazHHANm78ZpVtdCPlpkLqk8FZEw6zLTps+HmSsfmDMFReowLjM0
fepDCM3gh1quVrUtxTt1D1+AwvcPZCZ4ZiE0w2J29+8FEdK8/D7Rc/RJayQtc84g
O3emPcqsCnIZmipT3AIGA/Af+3bYRb3MYWuJbezaoLIDOWh5dZ2OJhgN/R87W44Q
29y31O+orBujHQcas6Zn3/XQyxWxldDEYAH/c/vAN0dHcj/sENTp2S1L82CqeqWM
+dXxbnu+G6p8vgMSereXelUOulaCuNT9TJ79nj0jRQZfLo9T1Sd3Fqrh4zKpldIL
olFv3BRQjr+MDKL6dEihbpMVsnOofiyyyxXW5hF9xTdg3F89V+EU2Wbn5lNIr3VH
Gxupe9X4u5cs4Cnf2pJFJfgBkhItyUMP4ts1wIemNn3QLjL2jbkM+Xe+YkYAtd1Q
yfVBBiwpzbLmlTitzFQ/pu7jAY9dY0oISXQuypR5z4jB8CX0SRrOcQxIfmnpeCj3
9ZKp7QmrnqgEdFzMb9+yTw8rt/S+aqsfF4cYUmclEzI9d7BzttfpYTEzxsAwq9tf
d55iP7+7ieoAD8tP8KPO0+aBbf22KbGJ4rLb6823pURHlx9POI43IBzCERYNENgW
bACQU6l0FNmtgS2wOWdLdciTXJxLxiaD+OO2QyToab7nodM92qyLCTuHhxIjyZYJ
mnRwqyqt9DA2PoljDWkvcIjorHErtDgTpC7krwkB62j3rMCtGvzQ6q++UiJPF4zv
gXBlPYFc6HH1oFD3w1Tkkd7hC5p8V0oW5kLaqriek2H1mH/TZqlqTIdf+MimGHEF
fuLrCgJM5GuQ/VrPcCBmTUShoMVyGm/RTlLIWmwvV2ZvMOYVOGsCgXS1Q/qYbAA3
CDz5vbo26ngMp2/332FO19VKxPiilHz5rQ/2RuQgZya/1WbsHYexJFeAuJwbw6y2
NMP5h2luNWcDuTUtYy5QFA==
`protect END_PROTECTED
