`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tg2vNJ+0SpdAyvCx2Gn/ObLkcMFuk+m0dHObkfBxVpozfxt4QSrnAzvFN19rVYiX
wt5rq+ZdMrWN03OVst4SjXwGTO1fWzeciCHUsofcpFsXW2xgLQXHB+NYaTul953D
kvbMrTRjSUiYM4593YrHmA2Yc9J/FYsU1ERjI5q6r3UWiR0+SEh9eZ/hLXyJMMpc
mo2AbUWpqIoSUi3WQF0ZgCAQcMHdROO9RrbKTOY4HA+P631HfyUxtNGU6zHaFX5B
ZThPI10AduDQ0kC+7Ycyc/z2YxujKeu2o3gTDCUGCcZLdiMMIpiKnDp44f9/ezuE
b971mHEKGRhEmowbh3cA39TgnE85QeHjker3Yk6WvybRu3xcKg9HDxWIvKrUgmtX
`protect END_PROTECTED
