`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4d68L3tW9zLYUzt7Wxwc/prFMlrWQ2VyXot+rN4rXn2EJf4DCIdGEOhyE9E57+G1
x3HmJ2jjzOXTaZPpZ4YxCiwVMGxOOIjTDjugpBJISPn+MD5uMbCG8Lh4dgQpRj45
hyBRByPhsKQo76vC1gwKLYMzf4clVp+NgNrge4sgrPFHCjRJ5A4nTi/v96GRYAzj
rpVrKE6r/wPMTJbqJyRKm8MDXFH8U5eFonb4+6NyxzYWvDygkILoj6P06NpN80Xm
9cYqqX2WIB7La+JvZB2zOvR+VcFeQ0O+d2DKB/rLYee0sWveOtG7PPVXsCYtgb/f
jDY5lIRoY+C8D6ip/hC44i9of/fJlCTHF0+Zj00/J5tRVyp2WE4st+yPcpyQ8tfn
wPqszD+mC09l/1GwEUM80nsUY5to/rqVmh1G/JZDBvfs+xoRRUDG482OvgfXIXaJ
g4unssgZ/hsgHcjiEkxrLUH6lPs9asM4SpKZ1VLc0+4fM8bQR00Zvp5WwvyBnzrR
oFbWr1rY7LTyasGonYLMfgHYLUaHAQgM9aU0Uyg8aqJX8XDcMpzLtPqhNYRkn60f
vZWLiLjq7TXZ6lG9g3DzwB2dyXL67XW+qZDwiAGjThEZR33MSr5dNGo+4VoKu2qm
lzMWhmn5orY+cegh+iNnnoRNd5Ikx5KGE0HkZXHga+9XoXN50Fd7IfZKrZIzAGRy
Tt6mQAwMLfeA/iYnw+RwEB8J5nUtEEWNDwJ+prOYAZoG2xiN3u8bQE46LaSYmZKN
j2W8QqdA4dLEjvpYP3chpwQVjjfLques4gVavolsLpk=
`protect END_PROTECTED
