`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NFA/6isTa+HpmzWb3afFeqaXAoQHysq53wTc11gxUC7pxAY48jZc40fYcAgStZNN
6MjvveCD+rsLOmBgBjFpxbLOXBpCXhUo52iUmSj5bKjvnBsHznhb/k3fw3vgNg/S
4PYunqGu9ZkOfus8I0FigS2wGLaZC18U8xBBMFA4vZq33GeunxRrBxSY2Q1+Ekop
BI+nh7bigxjxqOKKew2mYDOgn6uwLug2bWGiC0Ip6WjvQe4i42XNbhXjkzLKmonr
a1jXpKTWL/6OBMJFsKG0mfD9/CDqW7TA+aL4SrbLmBBjAsBs/Vz/7W2+7cCtrV7O
0ny8WmkRpIoJSPqrfERjgCAsa+3E8FRxYbVVNpeHjlJy6V/4km0/O2Dbn4IlH5uT
BJUCx2KQIm8NE5AZWCXkLQcesw/VUiSZu4ASn0E3H38mMQBuBrd9khpbazl+wi4i
rB20WHAaBf1uqqgCILQ72MOH2dPdM9pEzkaDvivvjdcZN3Wraug5937vIKP7eoP2
hjdCjYg5G1OdLi+5yync1NZZgwY55U6VzaO/u2dlTP85+XVdhyQouP0PWr+icgXk
LO3EK//yeCapQAEts5mo4jNGsWs0E6Ew4kR/7WjgNGy1QQr1vAOE5xUUl1z0J+70
q4hNAOLq4SGY5rdyQ/vDotFoWbNe3oAwzayuImJVabZSF/7Fi+0YGp9zOTJ1W6yy
GUCEc4TEo1ZlIVIN4mfzo4DROrE7NpOoCVNDDg/nA5yVmei4xWAnEhVMxE8QWPGm
vQsjGWBET9cFm2ikriCz/HBOVSdgAVvSxd3iVR6XMMwJRx4gvoLjiX1toMYpghfI
MclqY/jLXkOzDNj4iEBYLJUdhU2AFHUj8Qa4X402LNrFoJNJc8y5xElbMPTiEq8T
n4LVDfXcZrES0ANkVQHudijENwyrz7qmQ0NcazrNvWD+43UYwNUyRTu4uVfuH1yG
LCKp+4rAR8+oscqPnkJXhaXHPD0l+pjHKeY1qiSDH5KDP5fJbCzCiMSOAz0yxwea
0k37OYi8aYtwJDruHoEnolHxqtTKBe9j232ASeHSFcQO87WH1eq03BpQelKwgdJg
JlHVf/Rw62OC3qn9D6sXqx34BE75lZ6s3RYyAKJwiiKsJCUCO27Jn1IZiNnvC7sL
jd6QJH5/OI4JF9ND1mjF5W4Y4nutqS3DQ5vh5tzwu9ASsRfxoDmSjlC6M+ToX7a4
8K98ue+tsKKEXspQo5z3Dt3b2/vG5RVX2mfIBX+jbC/hz2fE0gs9zY+KqT41HNgq
jobritBZTLQAxHf6/YhYsy9E8IBleCDVXZr5G6B4UNWj1zL0/ddxc8tPI3sHEUSm
xG7bavDAYvQHlXwO3GuURmXTbDohIysQxgrzI1wECTwVHGbpsLNN5guPkQ9/jT72
2/YLhPq7ttuG9/KVogsZYiKl1XCa3grbUaE3HSRDo74uVeypydMv3xySrN30CIMj
y28yFyjIvIgwiii8q3cPsw==
`protect END_PROTECTED
