`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1R0RMY2BO4oRM1LqozhGz6LhSZHsJ30vOmdhHXJaRreI2VcSxd53neqk95HntrJ
bJUcSwadZ/gaq3KHVNQ81Xh49PDhLxE07T2Stwor1qbAE27aJRSdRurYaz1Fmuu4
mSK505nGeFb/MPw2uiyJqzny98WD7uQrbrcMEjHechcsNBYpgUFexaNEfP23uczx
MyxWcAzI8kI85I/z4R2SifRcoJHfC0eQT93pjDTbUsm1EhRBGaPKjWkH6slxFGj2
C9KQRNoyQOQVSS+9CAO8J+fNpBK+JSNYeI2Crhn9TACbSsRfHqok+LqTJo3bJCZ5
Z8gHOlgnLc95bQMwhTmQ7hajr1WkKN7MsHAgq7PDhTGEIqhTd0jy2LM5EPsAMqZ0
siUmsuAdRsLHdJtlDMt+euWdlvE+rkS/MQm/zoPjjtFalj0AWniZ4mahPpbu28c/
YqjcEf+Vde1ht7cl/oE4hyuSYk7xFlnnFH+BKzqlydACxmd1WrNPfRgTaCZ/+tgt
ZxxhSUu3bpu1rRNNt07y120et/YQmLXlHlHchdioYLZZKfhIz8m+VNshUfEMPiSv
VemPLNySdwZ+qTW9gHNd99kFtX2eO06Ff41XcOeDAgheBOdfk32MUpbxRy0TYU56
Zu++uBhoqiRWfgEPV/xgPMQMHyIO5vEI2jpFsnMJ/5gTVDjkNMM2M27UzNsoVTDb
c23PqS04qpKJ5Zz/2WNyN7sLCVl/jQPAR3X3BH+gHNhLBo/NBatQzOOwWArNIsrE
rdn/2c3Ee/8XMJlqoaRHZTjl911CHHVKIpLrg7H9N4c=
`protect END_PROTECTED
