`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6hFuk/fYspHfuABEkECsIU7kGC6qFLmu3NvE84tRoqkhME2TcIx7e0MQ9rSEuX1k
viZfbad9zHdwIxjyozoqpS9S97Wis8sT2huDV9Is2Fe+pMI0vGbND42lGHALR6bU
4rPDJvmYDLbkhEXfaeTnvh6/iTO4+rc8Skyy1EvV/e1QBs8X7RWFABZMj/dCghh/
VP/Rymfr08+hvL0o532BrHIqGpv3rNz3NXe0pq7r5zti24DKA0buxoolrtFoE1uL
jq8hYJsQCiogsa/+hZluOyheEz205pe8TCcN7opfEDjnyZVEJeX4AJ5ukb4wlDO1
kH+/E6b1S3l0H4vXts9fhL4mgpLhyE2YK/RsW+wG1vPFHCGEqA/deJp6LxpZ1JAX
n1Bmb6MyzwK2NaKIz9qC6ihmSDt9vQKfALM+dtre70Q8frI9y6V2POo8nL/I9Cot
SZfkoBZ0iPK1x22zlyoFbMdW8yo8FQ3OB6qXVSGq9X8Co2HALvLyuBw1PuJbpEJE
XpoZlvG99SDtypfLGN0uJDdJ62MXcBOkqqKK1UkuQlmovzKuAXOowHGddRpw+LHN
e++o5lHTqaOOFUIQ80aTPokSfp4B6d+1MwKv/VZI/O22NnAUxn4sKHVBJrAhINY1
hUDVUQlxV//0uLoTL7ILdw==
`protect END_PROTECTED
