`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0GXaVYRUay/SORV2OtJvS1uMKB6UxiQE4FXyQFTB5IuIRJEsdA6HpRfnSz89i0VH
8aApAKmFdNyVdjbX4t2Vlls7QcaAdXCb+hy/Kt4/o+YsIquZ9wJiFBGtiKfuXBVE
hGDxEFZg+m4yfVA0W8MUBp11I3xVdHYTA3e5EO+1EThA1kmYu/7Zj52zKmDgQW13
DtcKqqGPpFT8697qeJnzj86QSbzg5L1T+NTBXDWKDODwJbAc9IMM43CsY8EnaIVy
BWfpiFOlJzxjb6PPXgbmPM0BsW6RMp18YiohDlXkTcSijHdckYwFAtfG8QnfTYp9
cs4SCTFpIgJBYfKLq4Z1EUyY9uMVfntI8fGd4ObmoQQ=
`protect END_PROTECTED
