`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iue6+7fBr/ez5/UGd/9B59H84bRDLFRAg5IHMkPaJBgbUq2PlvA5d9i5nc17xVMo
gAX/6LUdTxrIAuKXNDGgUmZMW7mdmXIkpj7eEb+vC4llxTiyNClY1ClgUyQf4wsh
rgKgjJkpAk1huWCd4ytXoz9y5lUypm1K3Eb5hdsCVbWukiRl6Udi/dPaZaz390UR
VIYsDP6mH+5Pfx/3vJEebNlz2E+n0N9hryO5H3C9B2a7YfMYxBnuj0e7IvHAPL2q
7ZCaayTl0rAvL3aVfNUDFsDXAVsM4m8UVVQcvQUix+jdnvxGw/OHb89zODZYBgkq
fIfbvAmoCBuqAqadS4weyfcRwC++nBReiFyNeiMvGdMFeloPZKUzIs0wOkUx1T3v
YRcBjpYp1+PPQNDhcwo9JJXoJ0+DfIoiy5j4VAfKzW8w5EYYVF7IBuLcTSMBa55X
TvMlfHUnVDpio4y8BW7IfdNiTabeV+9/I8XctnxDlU8eBnTkJdOvEFC2UMOLO7qz
pEXBjrHqnWd0VXiZT7IviZDF/VlS7auysMGGNRQxeFWDS9cq62uN8Q5j9QvblQD/
4bfOytohoxI3vVO0WkLCRT0ie00AIrYpvtj9CIouEFhqS3mMeQ0l7aXDJHcfI9Oi
1j0W/rqLCOMdxig6J5tRoYPJ4kiHP1ljZV7U/5iuEFZjIE9p0CGso235uhqx3VXc
01YahGfB7YXbpeGZEqV/F/naxS45+z+Zln4Sy3BQmauSq6KdQiE/1UGjwIq3oZiJ
SdZJvue4Zim2O2yob6SxyLb5TajNPPPzWX216T0ZQYbXkKo3LAK2K2Zton5HchtW
JhwJg1fe/QqAtdeF3p8bsHEUwd/k+Y9AzJKw/LSrL11vpDzKi+SgGeUc1JpmE1tP
1TiiJnh3tC5qt6y9P7fGEuBNy3duHoos27vcEN8EpC9+sQizz0DBVIvdOka/q6Is
Yv3rXbXewEnbn3fcoG8NA7TB1ntXEaSnz4hDPxlM3XvEwL2LJVA2Q1a5fQ0Y75RR
7ru38r4IjV6WeyM+C2+FHZDnB68WpeeP6EBEz4i204Km6jMGjvIeY4bRU6Pt9mBO
uwv8v2wTKtfx84W0YCzuHw0kFoxQe/RlbmHD+iBXYvgA0Tp4nfe3Y0dY81oEvj5v
nWZus77H7RzCVAiTrcf5Q0+pvZB4Z1rewns1b3bVbKihH7Uo0Rdhoax93fvQDagb
9Ym6zcfSH9zxFUJ0vlOEQg/gX80gT/AOsbG0F7PiHpbtYCVCjDiOFRSgZpGbEjv1
RkNY1L/h7RHtEAeyahJo6/qcAD8xBv4eVH9yIZGF9AgpsO4hVyCY6lwnq6u+F6lU
JgWjvErJBPg/HJ0XgzwIwsDJXp63YLh8LEpWX+wlcQ9yOVTh9HhL7NVDmYTf8Czz
8SmcKu7rLkuGtstnfnZ5Py9RLOiALLf+wrqH/DNKsWFaRBftqh/YbtaQb/y3LTKh
fl62KhtgngZBH8/vr7Z8a9GMp7bMEtuMcS8ZdyVi6+axFYN8O6hrXRTAwy58wfO+
LRFQZE7wStN+pXa/SIewgDaDphU51VGCADlrfkWlSsb/y9ZSSJw0o60EOT5ptbZ3
YlGdPWw359G0FGSv1Kfql9X5groWAx+w1+defN/XDGTE0HjxzEMCv9FBp8AvUWNm
QzNE230SaqgRmWBlElwGLphIM64QMrrxAKNW5ZZSyfXC4TdXKJYdPHRRpOQZwlKO
uMfEPHPAcChHzrJYkBdJnZXjIOQ1T75P5Nu0WZ7nFsA=
`protect END_PROTECTED
