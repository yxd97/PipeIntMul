`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O4sjNMQpp4y17+6rDzuyx+JRE/wOBhlDRmDl+c2OP6Bcf6yT0F9PbqvPSZnkOzK8
FDL+0g9YK6bdF2PD8TZdbOwq3aGfJgZgrUun6rZ8hfQi6vy/Ea8pPxXaBuxPeNPt
onIYyIqm4kkjv0WkrT184djWcL0NImT6l5yKzMdx43jv7BFYYy1v5gd7ldLS43EI
HrMOemk7/uYwYcmTogAXn8lUiLf1CFgW+LNsXH9/RoS/fmcBsfYhMnjsoQBy308f
pZ2ZseX9yaVrOrxjxQAXcCccuFZXQy5WvTRBghxpkqBJe1VfOMf1fyCgPrC5oYYB
nMT0UtTF2eU2Ea5nfIP0tuivL8e03H+rZSkM5njNF8GqPYz52NApxx75eC/IFMmw
rEDJtva6l/G1lMKBoAUOo3pTQ+WaEz8YlRAuRer5lAtBwnP8daCp2Bq4RBaeTtWg
gwX6fXC5kfEkcXDQI1S4afal5Cc/dvPUJ+Ru4UWet0AcPW+aX+7vLom2z7nDgb4y
4CSqHnf0KqPmFSLN51dHWRMy5QnezUBBXoY3Qrepw2tm9Nql6ZWBEkL7h9U9px1V
PRYCV8n5RHljdQJMNOP7GX9nAvutaU8C2NFvRI0Tmq7gSUfObHD0U48o4glfawvn
o19ooWSgnn5HWOpLslxSJFcl7boi8XzKGDZBTX3QfzzpSx1kH2T2zRV/Iw1Hvj3E
xEDRsYUZAAK+yjAAUKqGc0l3vB7F3kZ8i85mGkj+SIxOJ86uq1nPlPli7WIV+KKd
gu8fBVtA70A9X+etaoDzAA==
`protect END_PROTECTED
