`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lI5pXaFPYnqPN5gCNM3HUontssWsrfAbbK7ezF7eFbU+8NayJqBAl2vzK7/m3Erj
kDzelkDgylK2o96mLKuuB7XGycUCHMT9uu4mwl/se/8PHQiwQwStkEW7ZxAVEETv
+auNhMVrN9nKpogm+UxY9c31OYTHMDV1XQvZ4C5TDPbE0xUKT9IcQxGda0ddGku1
B4ak02KCvkVdaTomVAsNEUNbWPvsHULR0vmKikEduXEEev2Pp3wUcOibvOksJIO5
zqctUcaF9yjusI3CcpecojNHVPVsQq5O4D5JIc3tx+E=
`protect END_PROTECTED
