`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8dWPY8Siho9nixngjHXpFzKiBzbPQUhnlOB8/37enlOu4IvLqxMQJ/eoldsGopT
vMaNSo9L2zYlXIf9ehZTD1VRwA5f/u+VLx3NfCh58ppRWUXfhv+qLnhX7hT0vwKw
cICRPepgJb9Q0qiNvqw/znVbtei+UcWg7SK9V2Q/PxmjmDEx7b5uMAb7gcmrzVic
NGI3+hrTl+8qGh+jD+RYR0ZAzXD06T6pirW0W9d2ePN1FBfKn1lGkdjZ5TP6jSE6
xITGB07gPGhtrmDm0rqDyDRmhNBZfseUU8mSuhWnagGuEfZAQLwlvQ8Iqhjo3+3d
wBn4Bi8ZayAeSR5L9qM/kYgsHoCTgFDOuVLMvjg1BeXor900c7vf/BcO4e948HlX
OifH0xJ/+KkmYvwMKa4/6LHw9PGfmbXrzx7N5NuseDzR2EF9YVm4jy30ewKiQyVK
YW/nGnaEGRgnk/HD5b9GPz7dXEwNKUiPZfS/ScMmUXIXtVDVHrLzLeQVK6MvpcDM
/jumZwo/R2mgZ2JO/+MuLJXEde2Uqx27GefOPS27kzPsI7hl1GhMhooXq2Y6lfQS
dhhVBA3Bd/L/34/zcW6MkW0+J+NdPiqDV6BD7uKOULMCH2+vXdVj6qvi32GP0kE9
C/79Iohqfuyx1bBbPjQABsh2QcguxJGrxFwrT+Mg5SA7SXugE+N8CSkBBUT0wIWR
`protect END_PROTECTED
