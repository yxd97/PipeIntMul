`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9WB/4vm0d4keKQVnFpy/aTE+X+DTEAchT7MaNeu7edvWgZlsW15018Fs3S5VNPr
v/0sR66WoPdv2xOmqIAHNkIq+2IHuVIlmiDCFrGjOFnOAM/m6svgEMFqm7nkOVwE
/DSDX4IAtkfj8T6BxxBbccI+71V5r0aDdi91Gs/XerAoiJivueCWRUdLYVBbhODf
hP+bmCd5TQhQNu8GZmblyhxjxAT/i85Ju0Xyt4W6T+0i0RrLf99a29SKUkHPb8k1
vFFVgln7LZKX2S3jeVoDER5+H0usRt39cU3pLArL40YOYbYgSppuxCGRTRVmWOXf
6OuxB/ke7e4XoDBjkv1YguSE4U+gieLAxdl4Keu/TV5WNX5sRcG9f6oVDspwKxCY
JV4xmNjAKG0PUh5lFtxDnOMD8mFJIjy4SvGNirDcn2YjHRN1PI255vEr6O4EZfPG
`protect END_PROTECTED
