`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNevxJeSk49CuPl6dH2xRQ4V9fIUkcC2DqGh8Wj7Sg5hLWYd0pqr4Bc/Ufvt9sel
/UyWWenG+LEczlrRtAI9OE+ybf0Ihq6egpO+uGAsHz/2SZ8Ays8wgPXY8a9gYuEy
jClSoMji0OxpVS9pZJijbCUH3pk86DhaGLbDtaWiQ3VweZW+RqODAPYQiNmsVYTW
UMrSchH+iiwB7MjsKL2m3CYCBiIo4uZZyICdsa0fN8mZMh3X2dNTCO/WhOY1LKTA
D4AUcAK/ZiIXftaM1i2dxdjHvnqxrBBPpeSfUc+YvqE=
`protect END_PROTECTED
