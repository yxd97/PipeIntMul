`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TQkO2+lBsNSYUYbCthlgwMM/XAuU4xXWjB40a9K7ivntk1Gk1cPvzVMwfgUIX91N
aBVMPbMjnpJQ27IddY+p9Wo8SazsMjV6/7v3U9EsU+71QszjmuY+XXQ7qlKCsEHV
HQvXDnqQME8QKuTlgXBzzDZkWe04JJlwbq3OMEQfgMu/pS08Nr3PjAaackfscQ0m
MxqvqGcXtthshTyVsOWhX8DueHjPH4/cquyE1Xeyc602JMRNYTWDhaE04zirqvFH
E77llqZwNceYHbgw+pv2we2EO809OqmE1UaB8yI9NcUtLx87F23I7Hh4cPDQbtUH
I+ER8Tw8Vc8aOcH4nOdqoenig4Xwa3WXxvYutedrhexyzyRCj9bxfcwXfGCyCP9N
UWOex5uFB0zBSh61T84LOTDZJ5faH/MO6mbJjNjHmkAM7zKxCwmX5U6BNgYa+CcP
`protect END_PROTECTED
