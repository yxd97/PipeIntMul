`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEl5+zGONiaUcJmzxHV6s8ym73bRUMjkZhOQIBcDXGmkLW6pXm+HsP2xsCXaJLo+
grHSdntbVPAHDg0dlc0p7Iqppa9EsilkJGOra+UBxRLusCL42Phs/qqKmWK/zUnJ
8rqVEMeTzEyK8c1KBQ3NBldZjsdxmjOH8VMaZhd6lqGxJ3/ZicLvCn5YoTjQtYS8
XOTtO3BxmQL1lQhqAwVdCA2a5W62dKvPaTPMa1aWn59FqFoi3p1UC2UvzIJNnnG5
CBfWklqsdzrdrE6CKVt2BVahO+HdsgNIAPe3rvoQ2LxzQ3izmvKsAXiJrKPOuMgc
t5K1UKmMpnuP+XH8pkuGvQE12Fus4hG1oUF61nQIMctAYMFhgYmD1Wq7yUujba6Q
hC33Iyz3l+w/QtRhP5dAMA==
`protect END_PROTECTED
