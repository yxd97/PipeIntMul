`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iC1/BHOZzjQXng7mkJ3B7FeRGbFx8hZDP5RkszkLgqWcQ/5N0s1JatH6IitU7+xO
OgMvDGU6v95Cn/rkT6mY0lyoho17WmyT7hmfiplff11DUcqR9lqhQSo7KtSwVfkO
QwEDtkRiYkMMfMRSxfIeen8000aOm4ZTQ+yYeqBMj7WBm7ICKjaoudAKdrxZUjRt
lQXEDmBeqStbMDqN0qhLUjlzw80Rma1gDOhL++3oH1qu40UCPjQKlWh7SnIBoV/n
Ipci09//tkdJ+3T+NgHLoSviLSSIH7F9QJftHDf6fv0AzjOCojHlUkCxaUSqu9yV
zfsSj+bD7nLJkzvbH/og12xSXWG8lp4U4s5UpnM813tP5N2j0aE5SOsv65/kIV2D
YqivACjP57AN+hXqR2vL5zW9ijQVU3GFigxdtFsNRKgHl/RTtvL3qR3bKDrkQCLH
hzpAE8LOvg4kJ6GvT6SCyVqAvtJKOJ0xum69u8Rd8/YWVBC2iv2RiP97ib3fC58A
0mz75ZuWwRd2FOUt1TcU4QFHqFrDLxRziKGtoOjh5gtQWVkbVKUsJYkyldUNPBxs
`protect END_PROTECTED
