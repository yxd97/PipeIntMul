`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9w8hseViEo0ADheEXADe72p0CTzPwm5zaOxwtPd9NnNqxFEsz/O5PWo6qZaJLlqk
Vvt9jU7hY2mLHBfFdIioIGl89PIiv7ybdio8tjCm6iHZVZ6HAn82CThOGxvgUp2B
CRgFRarNLGRC4+EJXcYniwnDIyxiLHQVH1D6J2A3qx34TmxAi5Bb4yyL2WVZLrLq
ks+lpM43MX2MDcYFwoO+ZhRAmEX6PY3xlDWeD7PtxFgFELheC121gas3BeSWOam2
Bs3wCzn6FaFtfEqkQcUPua/XjV5sVyBVSODfnDZnHB/14MB47FaP5qxeyYJRHuk9
caNmDs4viywf75F+i6ObqEVVD73D+5gmhbENFluwXmrcWCKrBXpKOJDz/Aa8m6bd
JKlJNzkzo+qiMQghI1a7baF8WOXTvBdHsXaE6bMNtOmLfqIj6IN9DkE0mtKFRSsp
zxwO3CcE9OMJk0OJTlKtXBOFnipBqBjsWjZFSIG37Y0oIhByn+/TpxNmW2nzj8vk
VAsYke+Y/3dIJNV9TqD2Ed/6CkOmSQvzX0f2JaTwI4phgawrmMtRrthnYhISsueo
mRJ70ZvNKB5KMuFwlh5wjgLYRUgM4iABkuDlEnxCcpor0R/HxNyoeTk40OK0mKAX
OUdMlV8TPEbZswPaCCD6og==
`protect END_PROTECTED
