`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dIir5XRjlaqd3N4+7MnmpX6DQeEfIaeg8DpVKcSuGyfgbUDLbD/FAgm+yWdslV9z
Z2gg/vTUCpRNsrF0ygrCV3Q7prA5o7ydxEXJpSbbwDCPj3GeTN0EzsfEj7KrupUM
p3qShn3j4JPuF9VPUZjFiaGYUwv1mUzIPT5cbbeCaCFhrO956ddmKxcrf0Gyad7v
NUqUgjhen4C7B3YwSQ0sXWAPW0XRKzVxsj/PRSSh5Az2+IVhHPJuVmQIb6CzMHZN
1sF52foZ/GG5xiz/C3r8rFERmhvDVBXVeW4fBzExhfqvBIyLLZhn06dtagN4pYRv
a9ZGO/vCKLpjih80SKuTujwUjBadhxPKGF/aD8Gp8sHx9dH9WNuszgy5cd/cyS9R
v/0qemRHnLzOFduiwqYDwdL0l8JooHtjyE2Qq2JUIAhRTzDTwiLMJoMqle5uC+gj
h/FBK0rg0NDDn/re57oicm7T6uDeJ2cs4d7wdXEWxfE5PkUaKbqKSDj41CTZOhsI
cPk9BaHB0Jm/SmhiE8/coZ6l9zPxuWu/nQ3B+p50wAk=
`protect END_PROTECTED
