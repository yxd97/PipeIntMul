`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4l0d3mmVXZNeDOKEZvmY3DATxY8DlXx9qGYh3he4GIhrglXTpT/dUXtmMMpVrOxm
w+/FwM5Yn7YAoP3rfLtozGKE89eoN7YGK1FWtrT2ZhAElXO5vF13zXv8UlgSHIOL
CSmzCQ26Ojbiu3IkKnUfw+VbQzdgl9ZpQq0G0domWVU0nCkIoBHAf+bHFDirU8Nd
GEJm+fvHqQSIEVd8bbKsfz5J7uWTSzVprHMXdAEgMAV8lIdXgYrYas4i/fK/CS8t
jfGMOMP9POamkm6Blml1Np3Q/svg7jWFiyU2cWarswkD9r5MCA1IhwQrV+HV9VUD
7bD6aqLlnmS809TvMBcRvxIQaWLTzGhdft7wT2nykv8bigumH9uSMsfQFMhpPSAn
68TPVsC03rWUQeO7TliS5w1H1ZSMd6azcS7pZ1/JfGKxmLNAALNmtrrSqcERE/kz
mH7UOVKR2Bz/3F1WKDOiIYWRPEk+mO4fq9OL5jvPS9b+kcMu1dnc0tLsLrQygCzW
tTgbomn9khl3U0/NyiLA+6O9AzvYN/TlFc7Luc990Msjy3OaSDm4pCTvlVApwab6
baaYvyhKdCVHcHbDhQH41de2WuWrof9IpzX7KNiIQzVPVkGNQOwNnT5UTyIfTLzz
SZ+7jKDDu1ScskosAw4oYx0H5emfwf7H0cli5u860xGX6bwX+gi4bCA5AzQOuKmE
XFjCNS1XoA4HdfZoolq42bpeNTKa5r9fIMDkXxLhmXNwTYIyvxTce4kvFXZgIJl0
/Few/y/HfkRPyooiTkBG8QhSPN/hb45R7iSavzgTCK4JAIcOED8KVR6CodJkCZBI
b4vwsyk/yi1iGBKEGOXxFQuIX4QCbph4+Weq1fCJ3x2gnzoRCT814BnIf6WtpbIV
BuiHWu+segMUsClVYB4+5FTDB6fr+bSoFNfeHYTQcf+M2INCR493kPX5BswK0qK1
fwNsIiKjD0GBl9M5BdpbCC/5jW1sRoZcsOp63Q4uNvbh3w7MgwVWheM4nUGGUV+2
DrIlrwwqjDfEYBBhXLLKtvvCTVR9xQ7AyKnKV5n7/Rah0h1SpJKQMFx/UMvtgQJh
LgHGgCaj4HY84UfReuOCxtx5yBRH4iYB+wwdyMkoaIUoeamq3ySLw4i+V7qnKb80
AlcecgLrhoVbcyhatCC06PQA6x8yqEPiWupXPrVi+raKUBfFghYumapS8F8laNsY
3Gr02EaGTL7eTcYtTqAhlRvj7ysm+n5k2QTohPW5lsrFLgCrmzZ6oVWBOQNgxZKT
0/zsKTrh1Dz6kIN6FVeeqQmgDxDaRmxFCiuPGX7liRk5KH0fMUYfqDT43rvdHWxt
hTcA01Z5tYyVI3m/vP0vwoiAhgEyF3yJMFv5Dgm8J1ZudeGPm5Eb+n1pSrzgvbMq
g+T2TdBXiRrOh1mtWVwouzTrEmibBgOvVi6O63/ioVsz36iXIX9Y+09bgv6xipyn
k+SH21Q12uPoDlyYdef/F2EH5HNwGp1YV0aaDJucpNmwV9NLd2PLu+X/be7HpdOo
etYmZ2JXBvV0OMSXoGzWGXK5m7LoETI1ixwwwRhljLmjZQ2G6BQcGc60ZSOqfhDM
l3NtsosR5zsp/Tbm1pZDoAZVyP9Xh2kNXDhNPfL4vL8iN8f7qGPG7XG0sMqQzB6t
isuLZJjlbRgDh2Pd9aeij/tZoTuByaLvQEvks6l0gQWV+f10G7LIS9bqMsQJjKTV
YRGHI3sFbBUevc9QtYtbouj9iOBUjAdKbUdTTS5AErHTk538RTEkD3OuL2PswReK
UFMJl94w2vWjaD+wFBV/W+b62KSPH6S98HjovsOzIAAf6UBaAQxOGaTbiUt+sx6E
6vxfK78dkIziIxwQ80ng7Yk6osvR5aKu2Vn1LHLD6WSWKB0lqmw7Fj0A6/YW2YEp
7uWs8VEzPj8kwVDSZyvmZ9huFwLzvANtINqhptnxE8zS1ub+vWhoa4WopXWB+/bC
hqbJM/b6NOU2N3wNGawPgSPrnEgCxCxSv86E+4r/dP4mAMJxys3lWoWwN2OyhL49
fwgjDzON6oBcrO2DUyKQmRmeVHahSGX11Hom9dYZh9RU42mUlca8G0MB0s9u55uC
B9QIR2nDaPhMURSYw0iapLEVotvAPwYxWJbBugYpsymrzQ6H2bHLR3DpmmqiMkDF
lg6g7fRPpMD7urrRi5DGYVDnDAxI0xikAi79uc1naHxZqCv8nnKO8Y/PloMFfF4o
mKpYDExqf/8JHznZu1kN7O4OaBT1bYxgvrGmlhe6zHG6OqvAf1o4U3HP3fs6FxEq
EUbCxLHChJSvs1k0QZIvSk/qR76Nx7F1kMWVCNnvQ3ptRem46zEZUlXAtoEWOW4m
`protect END_PROTECTED
