`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybzFbY+eptIx4mPBfoyc2nX90r/W/lLMuLALWVaJ0mZE2K7ybE0TyeWAbaM41pnU
7Ni6t2bJx207/Z8ugGVMTK2KNEUMohWJWbj7Sg+zkucg4X9UkixGplqTr3lKvToS
gifoEeHGUlW8RVzIc9H0EUTdeUCGy8lwUQ14uGmlA1OMZieMuoqF+QwAQEPZR2lf
Br/oQSjSjh4Q9O8ktWKEWn0ddu9XtKsBdnnjRzRPhaS8D3NDx/pd5HMNUocB7APX
sWpZ5kGYVSYJxjhcf//ddTy/GntIMbunf/+RzKlDHf0Itu9nvNdFBTN3OwlWrCiF
0bg3BbM5d8bINbu+AGDAaw/31gK6Bz8ygqWYHT+DjGmset49Jsv3K2o74eURqmSI
Wi/0S5hXYTyUIXGNoEUDLA0AMmKV+j8wHZoGftp6emoRZIKRmJwY2RB36xfokVXB
RXx8Wqa8WWBWMD4VTnAj7/JTg1ODXAglc/gLrvkG65IEIeScOOy2rvrB1OuEsqlj
6UcZFXbB3MDp6pTwBPdUFbnOaDVIvXl7LNnI/oLu8JOLKpplPCb9nC3DO0pgIwHl
g25WV6FJZvDTQPr54Ml2NWHTxZ/a7xCS602bMrnkGj6It9cDFXmkdUW20k8ItV3W
7+G3nNR9O+k2ZXso0mRzdZpE0RyreFjCiQyCYkYPJ+rTtJUWpFD1ciFikmgqtQwB
qnTPdleCDHLLZRuJkf+63jOZIbiIArO2YKEOBkE4PzpRTajRRl6ATinLY/pCHbZ+
0L1IPhgd96lgAzj+/LoAFcV7+E2ZFLJzCYryPXoSgKJ+kSfGKAAjWhEoLqqBt6GF
aBIxseG/cZl7Sb7pkZyjwsOK0/XnAeNysAfN7JIFLchREO9PlCDCX3o9a6LANif6
mTEcD/Z+wfX8zU1VVXcxN07nFMJN3oH996SZefm/f5C3DEvqv6wWeUoFBm/HU/DD
RfjjgdBlEuPBr4bGTqrDk666JM64Czy0e2M+X3JeYBYq2/sT+dUnGRJgLR7CsJOM
0T5AiooMGpWYzIvOINDFhg6L+IWNNf6zDda4aJ6odH23w/XN7bVf++7qlMVttDUD
BUy9LrIpRt+kq4bW7/+wBkwLkm89iJCxOBjzDFHoLzdcXeeb3NczI5XgzSKzbNWJ
Ds3tybIKSTDcbXY6E1AhuWDDclIWZuM4hklWEs4kv+KRD3rr/EXYV9PTtww4mqqd
QUY+YzjVIuhdg2is22vnYkWfGm2+ozB9I7CuryaMrOHC7x++qgFNZK+DuXYwV6SR
7sL9QV9/WTLH56F0qXv2pSIYAjBHO3pOnemQLNMSwaOPit/8y2WWU68fcmGJTU46
iqoKXScQQTx/RgGVXf4b8z+LhMIoWEeks/RYBuLZ2BtY2b22qO/Ilec2FrUWSlev
Wjv/Tp9Ltar2gD1avFLJb3uO4aqxP4rcwGrCwfrpSrcSZlVnldjbsDSJzS5pMaPQ
okq9Km5fJah24d5k5SA6GpflyWYIm71zzlUaQ9tl0walJAkTI35WlsRZYlMVY9pu
1MBDqiWzPDeA0QK33X60fnIKERQy+23AxCFyZqcyhIsZZYkj5Yx5iGsMp+bpKJmB
m40otqyHmNxPiiaqwZWM91vqDe5DCBzCAYY8YEhIbZei8amaV6mI9yusbZOsCaLP
31fUEQ5Q4YbqBoQRc8bfDICgRAt7kaefFdp79eBqN8/RuHTh9MEmEsSa/A66mdaG
tQ5BDra7jmyJYXyDozOOM98qleXZx8PlFCJaammC5i9/yl7dSrG5U2WOABul3cu+
eE0gEXyYQRqakrIQqwKVOURdj+Wcmbfr7KXpTZPysh8ROUgvhJsed7lucT0m4lZW
kN71KWgQvMnvjZJWvd+nyrMo21MY09HLMdymU7yRTYOjGzZH6mhvLCSQJtkFE72R
3o1udJ82nfwwZ7EQj3e6EksbBwstAKpQVeS7An5P78ooE10lkubBgQnUzrsmjkMY
cAit9Me4KHq4UPEz9g2JYxbiGwu7bsttSU2MW0cG1rNhFQYZ5B/fDmCb1RzYIwy2
UAfWO0QZzbBrQREoPOG8RD2/MiOySHHsa59VkGJg2fnmnqqWkG8UbDppBcECiep5
+3GH1omsFTB9Z86DtSx986Ae0yNnXACCOCCIJX6YEhcur5wHSnKqPuaG/mu+aiw+
LDaPaNvSyzHWsHmlZjSJUM/RrgrzZ4W9tEgwkPuq1g5tLh8pvge/LteB9H0KRPC8
M0O22yc2XVOD4W5dSSNio3R+hDpiO6T3BpRklzabr17o2LOqrdsUwOkerMxQvww6
YgjmzMa9IAkPLrtz6tPMAGFL563rwY4ECel9Y5LzWQagRuSHLtATnC6ofZ8ggLVb
AH6JoGxAn1HITpsrjoR54PfOl6gLmzi2IJh9quXoFH+rtvvhXoct88CuUMo/B7Gp
oBx1HNthYCYoJxBuxecohGICi45otKV/UtoJH31WbPTlxGLfBO+Yi6w+L14kODUf
5FvDamima8eY4tXlwGkGvCOy4XVYP4xSmhP4emIGOdj3oasD7oYTkU0uwu7DKiCZ
HJwTfFjy3513BpUPqnOaw+jO5m/zps4OikuK2vvjgDguhDdShynOteRIp6ehDKlx
fuwhb0X4+JevTSXIxfhGB4eoL6fYGe9VR8Rdb92n4pn/LnzCDyuyfrNSZMbyxfwG
TM1ivESbEemSPQDRtLtKGGH0SxgiW3YIrC5rMYrs4skA9JEv+oAuXS57p0X+cCqe
v3taGesgS5IsZ01YghzR0iVyvB7pbPyrgU6X/2UOrTOOV75ZtH9dbkYlyQLi0fgE
EyJ6oLOoYUAj+bPDiCJqz9ThZ8E3Udh2twf7dUmPevyb7M6SuspUKo7GnsysJ5Sa
/xvkhOcc/6GUKBC1rzC/HtQXq+rv2lcNrS6+RlxdGkQbaHWCNU/h2ARsPaezaGgY
pNpQQYAmezyBxFhyh2sj3PSWGN4+3uQ3a1HtbTmauykY8YyfIgSXAPqaI8+NgVGy
0TBCHh3jUcDMGv6h8A4hOCuIM3C2fKvYD2rr+Q5t4y+DxIUYVBUzOEEAyH8UcPq7
I+CoJ8JqDKOgQMc9Z7Ybuw5POIM5ctIaGgVdKJnCmoxHo7wDqeTx9aCkAEh+scmH
pBuN2zpUb4mO5aBOvvB7YOc3l+7wp6cr96+foXo1t9c=
`protect END_PROTECTED
