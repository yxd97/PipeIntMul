`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v2iHu1djQj+YuF6fFobUvLWvcAHC4h9us+MmDF63qSEWmnoijjZoDxwwmcwbwErK
IrmSfLR6rPI/3TypRKBjlXOVp9YATFZEg79Zm7pJNbFjc9YwAt5BGHF3IgotV7K9
lT/kqbnMEH4Iu1rqkza+pG8p8/vc3bIZrXWNyMB63l8RP+zleL0VGujbWuOIcU/g
69AgEvr1BGiHh3ocWWmMr1ectjxr7MlZsK9JaaCFrC/I5G/7xD4yN5bbPXagnAve
VLNZ6UVtW/+Cozp0xajLhktNHlC+IA2Ur6Y2FY0ls5pwIkp1zDdhsUPxbEd4M8DQ
AsO3ArKT1sXl3dDTrfr9V4qdAmZ8eT/JWRhGAQdTJ5Dz9iNHNsquRChMOaXkLxzM
yQkP+Y9jneKttozMow4T7Io7QS7JUMbLT7ICwHTwuLuslpNeyv+KT677pV1w9fqc
UiER8iUFu7+CJpxzsYdLDKW+Y5u7bTbW/YMcdb69PqrSB+/GCccWfem2EApE+HIC
qXlX0pwmOOLGn+QXfpzuZZKyVFIFO5mFBfmyZJvwO4FuZD6eszdusvU0akWD9cjS
RL12tTPv/8N4RQIcXyBhH59WPv6/Sw3iJM7QCr42twinGVgNqTZ0ajICHddJOlN9
iN/9wli/nS31FC/78gH/Aqx4/1iGokkieyrrFY2AKN9IITnsUqfMM+CKRnVgha51
3iUxG3F+MpJBoClCwr3codxn2/7qQ440C42szcYnlJ1GuTcrEb0NjKtW3oMIDjE0
`protect END_PROTECTED
