`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTPaX/Kh/yWXDWOiZrrYzfCVvhCNIopAcRJczwKwZiibz5tkA/1Cke0g6nbacxIb
LvSgKVT+FFwRgYbXdwJpjNZOBSY7slqxxP2hsDz/h2kIpe+e+ZeNFUMAy2wMNQIP
fzIRlJ2pZJgreF/bFQoPB4G7ldDLHl4MDqoTWwcsVIB2AGqLokyokHj6jyqf0p8h
PmB/AHfaEyT+jKcbpvl0AH8RYQqVC4qarArWMJZIPTHJRPqQe//D1nxl0rif9cdU
W2rMTiFY0ihOUl/D2zX2SqowJVA/OK96VoxZO22/rzuUtyck5aY5wjsHCkuswC1w
haH9j1V9OT5SiDNn/K9CRaEQDS4YxJWXGN0Tp2YntDoZBW4HvYye+51lITYyid6Y
KdgfM/fzAfacmq8Gcf6zHPZsR6YN0eWAmsiyhITe5U6YAGDmk6ElPaOJXZX9t/yD
HJvEH5TZ7WqfbsiqW+nsgj8KEJNVFlR2X/LspKVm2GEBRnEGl1gILrGabwNOsvU8
dXBVFPskhid9Ktoqk0NJJNE0KCDhS0S8GFn5ITfBBUiL3TcXAvPlfhprzjf1b559
bOem/jXdNTkZGke/p/XKts6tj6AzAfcfXuHRCLsq3ORjbEDeWIaJC52RAsXnztbC
G7X6noHw2dJp/4Q7S86tNh/5ywrGnNmp8rtSae39jKw9Jq+xtZ9dS5a3lSkqzTR1
eyym8/JunYNFbO57Lm+DZNLJYlJqEgXoLCZ4mtIBoqG7u0MNU9EtlfGyyLoFPcvm
xbi0K2VYitBDXCsxTQnYUb3CPdIqOunbfL1ePJm8C9go0vJEn7r08fY5cAnr7ZOh
oB6pqln+2HGknraGdshPGnIDUd3WUrMOid5Ld9BsT4+w/iTKoJAZTtlTcDC7ficQ
boGRaSbP4kWyPHbygqo1GK4F4O5vBlfzojgFFxgBn13+pILwhb+M7Js/onLqkNQi
YF8irztZFMdNBkEobIOu9mWEgi0jdYnNiBqjKQO1mp7s5heyT28mNNV/HQVjN63G
khnhZ7tOWH0b17pB5GToplDfxjF7C8qwF7orafrxNxq0NOxylrp9Q/IvOQQihQ+3
kTryB58XR++nnizOmTui+9X7dErFy5Xw+r3XV4CYWB7KeanP/raH/N6VsSA9zMHT
r1wXj11OXQ9BV4mwtCVbZuUA/k0oOmV1uY6J0KcuLREsx2+0jPJg8CJH/gP70oxa
WkyzBPv+DFrE5pBjCx0f8jpqb+w37hbubC/tdLA5fU6mnPqcBl3NchBE5fhVsh27
KQ3Hug/81cJ9bPLDdFo/JHloyw/hcMrJrGz0ZR2RLDLDZ7jyHHYcON4FmGlawKW+
7XgxRchGeyG5DpCZpN0562QYL5m6+lPaSNsSTiCh4msrnxHpN+RqBBTpch+CsgFi
9+FIeFfJU2uq+UfCGOUG4WEF2iSaygXuGmpCg9gDgLrU65CfKsLuSAn84xfQQna8
90z0RcMlUpt1sAd6+63yuxd228B7MIb0U6hUxPZfA7+syY5rVn/PY56M6/5coRXc
8WOTpguaD5IZ/8vetDJkyLl//xH3WhDZBEeCNtOCUhf3+ZrUp4zP+NEMe77JMYMv
dqm7HaCqjwAX8bY8vgX/3owtlJ8OJXCNs4VsYWCsvHWkXSZaSke38cGNAIFhlLV1
0rWDG8fzY+m9YirHK8SmmXNh+7L0O284xk/9stH/d5UYz5sf7FAuQp3L/dH6QJdF
7hJbJCXsnmUENT4stRqAbA6gHwHP8Oxg2j6rhPsbfBmOq0Mmg7RmwcJHzhcXzU2n
KgdfBGCZNK2CenJAoBzQMqIy/B+pfgGVVYVhMJNfV8ba+OBRL/hv625DXl2osBBl
ts5wfIm9kqgAsdRxjthgIPDSIjXq/i4tGry9HBdgeHGWG7CuUoU3IXfY4ti4X9vu
hwISf6lAZ/PaOWycCG2k+2pL0ekGyVy643jl/TGzYsBlHVrKW97AtF3DAK4ddk/Q
hAVG1B4FG/fEJnsAbs71iHBLSL4CzvZfbvxME9c8YE8ptTMAMnslhV6uryEZy8Vg
XaCVzGtO+GTsNcYATIb+CUzAQXnwdm9MemL5cXF6BPTHcPdB8Y/IkRlL3KdXtCs3
Ay0EB+nREGkVe7beYhWGHA9fA6VRNfi3a0oX/1LWYU5QkcQoAouQE5ClmXRJkWR8
eRujz4FOHg99MJu/HKH/l8cGH5VKm+xhvHFA7xaGuvRyOOkYHjeH7MMchvma3u8u
uBQukSQlssMCQsTTL/aOrFkp/9gJRqR7ev9auUINUkAJVW9TTeAWEHboIZcIIN+v
x1KFrTDuPI+xmv7YohMKk7u+bHA84fL8s7tpXdvrY+D5kTHNLlqMwcr8POQOICW3
0T9PXU/wcRky7BGq1xEroVET3ol32dmyHAgl8WGg84SQcG57Wc3jzP6GvHMz08On
BWIZsHEeziSCOvKpBxqdtuoYL446F4KiXq4WHSFEGxgO4UvgXahEovAL4Fug0tC/
zLTSBvzW3ZV6W5aYqFnbhMh5TUqF8RKm4YLY/GhzSgECtpPTJjsAR/PqfKs3D5N5
WqlnpVf1HqWo3sOq1Qwo6xjcZFDAiSJc3yGWq3aio00RkpBG5obCrpgg8fnCLoLV
OQOTQCyMqe9qd8zCEm1FKwtJpaiW9znywC3b+7JCcwjIyfbEaGI8n7JXWTNTYwOn
mQq+09mckWvLu+nlOQF3XB92SMK6VMDODMTki6cRKH+EVIH53PX6cK8wrsSskP+/
bG63BTKu4K/zno6vCnXSFO4U80f1WvuD6T50rUtsMnJHmo5od1CqOQVpYrBrPQky
eWFUqsEOnkpCb5HDQc5UQQqpZjEebm4bu3t6dGU67J2dZ+QVQV+PxtBKusgAF4AF
+u4n9Z69N7inaGwtLXSdE5R7f2070vMfgjr9sMwwOpvMDVL1sRtHkn4yQ/yKL99u
tpcVDv2wTHZqFreEvk5NMKIQyzg7Qyk0/9yxEZ40lnvWH0Bf2lYr+Y4u3aTp1tc6
jTStakAF9ESmy2uIbpi8a6YbWdSzxgFKyaLruasEx69wlhXuuYXNhJrZokQUxYhh
0/rxiADEPWdbfUOjQ5Zbk6cBCvDxtzfTPLKd6CBxahMZ+tDKBIE3g4tsGJOlHfdH
vqzY65N67FqvP+TdVYqmYFh8IDVktShCE1bq2PWhW5rWs6x6ANnm++21lkcyMkKX
f6cLpyKlslZ8lEQZZXEKc8YSh9YntAexsSX+eajZt+3Im1caUSjyv4hxjI53FwXh
gOtvX0dReqLNSKoHOr/VM9tEk1YxZt9iBkNlgs5Tm5IQDollb21UtXiMZkeo0uYa
Go4QCTSxtrkLe20b5sGmBuxyqBLdA0+EyHE4teLeXvH0WQTBoZG1uLKRozgWZyxK
cz8H6rk4cWZLG7XezHxYDZWzL3n9pOhL4oby8jVXX45IMDa4a2QqvFBggUSjF9ki
riohMXUbBK1DDp47gNNk7Pq3TXLdYOT/fTgBcww4GS41Igdti7+IjybpLSdg8wn/
efCQy1Lg59psMaU97ibeSrhvAa8fjsx4NkJA2zFQ6WGjE3atAs06shSjEA+EEpSU
tZzz1I0qTluDx5TsiMcHM1PlbG7Tu7RKgHCSK8h6jc3ATOyyW+V5nthKHvy2dMhX
`protect END_PROTECTED
