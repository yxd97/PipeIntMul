`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gjqr9jCGheyK0sLPQttR7nFty17FZ/YF53vksRS/S4lB+S3fS2TWx/YJorROBur
V8O3ngLN2F68qr2RCHY2jzpLVM0YMONHGqx7kufrh4wjvnqXkbjdEtmFAgdl6kFJ
tmKckvIYIFpCvj3ARDbjhX3Kgzs6R5rBM6D1lm5qXUKRupnCYQxjV2fNjFu3sKU5
Cbro4ySok6KhO7sFIsAbHpTP2QmHdxpXCYIPbfpgXjBeuVgoPMkfUjDR52q+sB7d
wuSOUPM2ty86zN4SBmhD6iCw9fT+GpuQHaWAkHEOcCYgjL1nSdt3r4XZJ8nfv83R
w27djdmr/WgpIj49wptwQijOxIm4hhx2vO0QkpdTnpvM4eo8rg2LtNnpTHpSLOEm
`protect END_PROTECTED
