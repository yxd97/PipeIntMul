`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qmF8H7G8CYkrXOHyTzMHzcJZCG/8z5f56I0uOJFCfEzBuo/vzj/ZoiOSjga3wdG+
g9hLT0Km4MpoZJuh8b7l5SC9H1nwE9+7a5v2OTCxyNfenEliDoLP4qs2pPcbNkyD
wHiq0j8tNJXA6vNAQYeIzVebfl+pRJFC7CNNzStv590lfmbz8+waZxFvpWEjS2kV
uKmDlbnCV57k59SgqJ68QvhsvxJ8uiez3bJ6OuLCoLakXj99lmaiUhQ2wUdUAQe1
jw35GRsl5JognqXtLXVDhRIt01jzP691SvQWmfybGKXcKTPtpIH8ylerOrwWYlCE
CEW2FMBFJGhgp71GryROtN63aitxqDPw+zEl5xmVEjfkg4X4EzunpXyMgGo0Snzd
HxL5TVfcHmnKaClxgH+81SoD6vfuw5xwDHRFGKECjEvU+iii/Wd+VL+3N4e5q1aK
rTE2VLX5KfwSO79TVRdRqQ==
`protect END_PROTECTED
