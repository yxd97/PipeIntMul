`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YS4VBQluvxo5atVQh6mNUWE7jBXj80JefT2jxt8ak5mffLxGrY3I0L5Aw+FTgAZR
OAW04GOooozOdcvS82xsQzS5QljdJHsCWMAcHQ3FOdrT8D1Jpc56YUCLW0WjUEAc
CXqPb8HUK81RdoH84FrcSuSG45Kq+86lOfXIWmXHJisRd9zOe49Zjs19okywBwWZ
jNZAl8QY4AMH2xPXEP0V+MnE2lS6JkrE4YLNRRTRZVvP5bB+Vq45mmRf/qVZYhDe
IgqSR+Hi3eyIYT9uq5uaZyJkIfa3kMYOJyGJEmrQdWs2bzjdfZffl/zBRdEGq+jH
6K/UO5POhUUivUpgY1NVeh9EM1ZPF94pN0XlWHMatdoq3VCQUp6tIkqTK/yW2jBE
FowaRZi1wdh4uCBgBc456ejq0+doN8zuqm/BFQUC6J9WnZXRI9ybyiM12H8Qb/Ld
vUz8hl1VLj0PQIH9pqdIhzjw3neIHqt57rTGqJwnoyFLLamJI1coowumRYkPTyTM
YM+yQ28vj1Q5BSzMnAc3OUi7Ng193CoOc7/Yoej2ye3zXIoGhGBbDwT0/VLgYse/
DAJ57BTDX3p3DDbHnMxLRaQKu6/JFCbMnVHKrfqxIii+T8gHXHaW/fqyQUhjhTnq
w2FU7Vp1qM2104ATVSq81eQd+aHHxqUyCR185CMgB2FzsufNMrl/C6ZxxoguCbzb
LeaqD58Evy+NjlKIoxCTvdTlB+UenMRIucr4+gjSOzPFi/J+fWt/tWCiRMFpRF+a
wQ1syELLKUQTx3mZcKTMfolLbiEkPbguOOo85BVYv+KOfP48E5uZHjgfK5VxI1q2
yZns5ZCvMKpdhT50duMLN07NYJYhZlBjipe8O0t5KKPE7NdAjLeZCQFzCsYKAZ+O
gIhafH1/l6WCqGQq7NCDRNziAldjiht1FpgRLwsS3enfSa8ttZ+DLGDiLu/uv2BD
sI9AyKq5WUZ4G/wl0jUqOfM0mi7DJUb80XfRTVhzdBHh8ieQOX08JwbcGUU5iOB4
dlLloPn4ajCh4FcnAKIFbtImKtW32Hc8Zs962KDlIkxQaqh/K7Hl4hqL1+sqEVtg
R3twgukPzgxAe1HPmriQ9gtZ+ySkHW0VY+fL4bWVUT4so9ddFqs81ZA2YQ/VzSsM
ko0aBHA+lEew4NycR/KQZVJmV/WKuemuF9NX9gBe6oPVKaVANNAB9YXaw2UbOule
PXVpEjCZV4OyaUp/38/RDs6ND7U++r3DzDThyYTu589hrfdS3fgIQClqEIAlRlbc
E2QnTgTrEzE663sxxHgustYA9wJyfDFKoJz4ztU1QFoXcKg1HlLFxPzdI+U3vb4c
WzXf+nJms/IiPKajpZYRKnggeOPlzt+8pMG9w12RzBTpTdhioCuAItSHHwWUA95k
tcqiPmbfP8qGMP59UDwb3Q==
`protect END_PROTECTED
