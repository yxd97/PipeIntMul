`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u34RnjXBZVnGkRAREoVnGagERcwRNHlFjAewx193IOg0Dnx6byVgL+Ho0Z6Y2aEV
8o+wtdkZI60frmyxTuYWwCRXRwefEJ+SKPDObkVDz/uMomJrjWl9+DldIHTi8Z8o
dMT2yuOcUds9D/wFr1lC1KfMWP3dcqWGYOwcmY8TR0tf1SJcUJkmm/DyKde3ksBr
mA17/T5oTc0Yh/AoFurKEiipu7pnMY85ChGagUtmdgWQL6IQK7smzZCStnkZBTt/
xMu3LTntMrcHwQqPFtQGZh9jODhNaBdHbsqLqkbMz7cIbYuH6SWJ90VOpiKZFhfU
WAc7dOn6KkBPYnR1+LFeY/gHb7riL2MEQPGidGEUiNg6rqIj7vSnQmnVwVp4Z104
CeRJCeYbW1S3ICscLsRGdbUowdmweE50sZpQCV5x0OUBYpomT+h17nMy+dNRZ5GS
PGf6rLh1GxvfRW+ttWEWoZxnl0oMiN8KPhfKKqkRM/YUdtydKeXOEX/J/Ra2hd7G
Viqm7LvRzdGAuFht5RUZcbDKBU0CmHixTrxTDYvjqjOijuvJ5iCJ/beS+60m+Ass
3FYJxySQ5by7zyUCAaiHXogfhJc9VJOX0dkymMD9MYNDGbbihQbSvA70yRcqPzbx
nRl2+ktJoJSLKUZzSOjABuBVKTgjP2TvYD0e5CfkcnzzPZZuI0+CCE6DnEwo3RBU
p5kCdtHEn4LHOtjxc2RWw+FKln8ForWyNVo5aQUnSLDWLGNXuAk25nJDMp/8bSLX
H6K0IG6zt/bE82gcfOtl6gm4o1UU2aCzeCDOeNBQWgwzDiVGGyQGrESTQF2uwhLS
oz1sOctwSUUv8cFKY97Sap7XL/NHkSQsylmxuTb9QbPUds9+Cvo4vS+KHSzB9Pjh
Dm0dCe0mYYM8eOptELOJIhi5bAktJCGaKl7vkbedl/2cF6skeFaf1snXkDbr1wjN
`protect END_PROTECTED
