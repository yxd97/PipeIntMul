`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e5fr1XPnYk2leNvE2Irs1VTE5vklhzzrY5L+Z7gmQ6qiQ/l42uyKqHgS0J8yju0Q
7o/lzi15un0V11ceCSwMLMYYeTYt45UJWA/BPOfoxmQVDMX6bwZylExe5NgFnFLT
Q/IILvzinziyNpBIYb6lpPgKuWsDvRwv6brgBmD3R0IssBP9oEsk7Q5Mos0dFUsH
JZ1TGR/wU5tB6/wOmeGPVO7JXUDSuxF0LMOxT3V7WYcNH9j4lIMobaRoF+lt5asb
IA/XrPZo4P+HrhyO8zOeBffbukS5f7QHF0rEtcnTs8JPJWVs3UfaYH6msYOyaw07
N1ONOZgHHc/06QCw99UyuntO2Lwc/JAl1tLEP6bgcDI76lwLmRyckDVoCBTGE9xa
VGwbVzf9Kt4FhXSDeG7250j5vzEbE42hyF4vSsHed21loid4yDB6h1wQ/CpjK/3r
RmiJ1r9wsmnTwnufRwbYOSo8DdQ6dtan67Zksug641X26K8zq0wQjZcbEYXoj5WQ
aXb+n3cDLCiFJV4+d9K8N/Av7YlAPt18TwZJGGS/SrSkHOv5HgFQTxq9ndsRy/pQ
QyNsF+bkGmgaYAP2E9cARzgAoYcBG9cnPdJybf2PwgYJreJ1GuF7/vyRcaH5RObK
7wdR5aZCnx36nNIHX5Xrjs7QoCnesMY/Bvdc/xu87Q56XukCjJFfBCXjUZiuar7Q
UooGnUnqbAxKZ/E9xVn6BVBQdLmUIGe4PmBxruDCFftyonfe7/4JjavnMGLcpJcM
WV5h3a7oJWWsznja/YXqsUGPO/cVTQnwWLLsXgqlcG547SMufrLM6beRmS0TRgXg
cyHt+YCz1OzSkF+cXd2A3CtgK5sFaiX45Koylrj6J7+wYORIwr1URliq9O8iDk5J
n0nOuJCCaLOSX3ddr/54x6nGP6BnQkfPkvGG/TwWLUIwVhPGX9sYJb6QfZYeQkmu
DLjo6uWR9cmunv6GF+eruLtXrUSmhuhujE9a4X73hlG3DmaamST7B0omngiHu9LB
3EOglNSBQ10FVQmow5o4/0hcpRdx0HywF/SHggM3ssAr2slYpkH5UyLNbHPbDQam
ADFHQhhEhAm32n35eiex92aE/bm4pAHV7x3G3GCb1flxEyUP1YPJoYgDQkK37XmH
vcypPNWDCUW2NDDAWOF59w6jVNqcUSF6IGcxmOMIFxgAuz8qY4Fumvtqgg2Rj9Be
S370d6XKnALSRcL7Nk+PsgE1viTAAnp6HlrTdJwSmQ4Qz0+T6xqWwTPoT+BJMD2i
`protect END_PROTECTED
