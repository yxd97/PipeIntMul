`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t7l8xDMumYdd5NDt+QUA+PHLx7I2TN5B763KYNkpZDs8gPUmjB3JcglYDWmmZQ+Z
r0ek8Ipiyz075fyY29kXVD8TtI8/hB1ARXLtWW4RzlFyySFHlXVt+fSTTmrvgdeF
1wdp+vYWk5iHQruqUZRp+Vnm8Yafzm5yzziLPHbPMCzVCRlopf9Ds1ZLmSsbXGM/
icmTH3oRbAj2S0t1QiPkWfpv222iN6LKtuNxUQeiKGaDtq+Gc6uGIOH7jlj1Ktqw
7yZnx50fB+MfgWpJC0cMW1fgv7P1/FseYQqoGdx+G5MNKGnU+knFT7rKgqC7Yzf9
7GzsTCnHviyIkAXsRrkYCBC7zTuKiMQLye/KkZi++rnoSH9eIpxNE0b0RwLPN4HA
zvIT1fj2sI4gweLcBtfDShMY5eNpfvnHqlz3apkRPGfZtWW5F9/7ol3sykkjInHx
huZfIk1x85Tt9ykGO8u1Ka5dJFxAYIo2q2n5ZMm5XNTI2cQIz3UApes85x13OPLT
OX0JyB+ZXR3V6Adb5P9Q8bQTyu63yHnanZysRSZUyJ5q+yfjk53/LxSje+CNnB80
BaKbJ9BHszX+Z3CkUeLnVXi4U9ThBiAagkW9ehOXH1L9EEwSAL6hYVOv8/0rzo99
kGw29Lx9PQ04KageiOAkLFb9ZycvI9xrEda8r8isZyRuq2jqGAOLXtUegQAKemfR
lHiSv98viAniDtXE8eiRTqL/5R+ubJTK9KngOPhoUGfr4LN0bsd8fLlNvJhbaEnD
n2NJQVlwjntI9nthB8SfwMn/IjvhGHrWVuNfD5luOmEUEA9G1MfIzfQnD8dLGGpC
lEXlVQjvrV9AP5oMx/Eri2QtLPAu/3S6NPLSe+M+yJ2bgwG+Dd9zQfyTdxSF1Z9G
DVek58LvtGRaRshtw6+xZhy9P8RsgaIQF9BBXf0kIx8hMHvaJxZ2aO5uNr1uDa2M
39x3IJliOXAmDS6gnTGxOP63IRdyGAuHbfCIWpJsuxd61v/F90gfU7yfzHdHyAdt
/UWbnrchu4E1xfIZQWK7NQmKg0Qv8Zvs2YLF1gDNuY+/ZqlmE7vjOjizUWxQWQ1S
p6QV3I90skrpj60kIntrJUz28hWD4necok7cMfgHinsDrBfbk+6s+JMsxQaSUoa/
BTib52hSdx3oB+JgCAM9h4oJvcv6UFHy5o6C6rPBO74ZBwiSgIXhizmrEili0pwy
Pn/Nmr2D3T8LHZ018VmT6EnSN3hPeT/g0XszuDxGJAznNCVphU6M6h2e8V8sHUlJ
vwngRHDx155XCP+FK8YmWIgUs8rkMUSGEigSZ3vYBg1xLO4MLW1WiR+1N3/2Pg6H
fafruRA/miMQKni8zNywdCDJaWiAfBE7sjORvhnZQJaB9mAReP3poY34znp1jbT5
AiupNRKndAh/t8KhlQNwpytO4FVB3+C7oCmQUjL5WWiLF+0oRlR1lfSV/6gprw23
wOaZR8vlUqu+XOWmM1zCF9kev1eEkbZYHaDPe4D7UgYPDbNDidaIB2E6ZxA6P1V9
RVhmaqMAo2L1WMgsGFnJvt1kW5vnLGcgTGoWtlcJeZPAnlHkISCcxeUGlWZsAhzd
kjLqCc7d8Gd5hDAV2Cqg6206wv89uHH7GStIkam0j52n/mTXBT2+iUC2gO7TuRTC
CvE2n9WeHeYU9akeZapDEYRF6+l5LwLsQwF+QrVCGWgvcDdDZxw9bj2aBGEpVoUg
4GMw/NI5fhYbboPKDmzBqFjvPoFZZKyrLJzxO6lIrG2IVHRHuQ6yZniln3ppM63B
eTsNtMpRSgSB87B/giCN4QM/UdB7F01FAcDGuKjoo83v1Dz59e8wXOyty7kJYa05
ObCRreknoVDXB42HP3rkLaHjRmiJFZns6lW92k9qhzyk0iteHKTyGniGepnysWr7
XI3u/HHXZZKOsliIM7F4tTlJLaqL1Hv6IKwYMrhUd7rDVbKscjvroLFDegrFvhlk
B8rxC7yQ0AYlOrYef+pgW5+HfHHbkAEFp1HO0QRAqki1Cv34ZW2Kfls7CqZ5z/5y
Ecdu1INpw3ox+c+SmZ2lvDCkn0t67HeJZnUJ4pb+uyP98xI4iAgazD3xotoNscoK
jAWW/FGvT+ZRjh2wIMBD6YVr20O0qFOr+hkkQvzWqQfxdTPDtN6qoeimJ2XgLg7M
CykHXsBHB+KT44DZBdZxrhC380TNL0aFptzead+RbNP1Y2BqAxWVubHlEqFhBiJY
11qnkGIhvcV7mq2d9Hmv5beuINiCMUsHcIK+0q22T7YXBzpw68gcG6eJrz7YaD6J
de6or9pZNG/hwo8yK6TQsCj0hRellLkY/42Ynq1kwG41mdW92AwTotvJVl/e1Tgx
dStu69bi9+8MdpdGlIhjb8sUQVUwbQptr7YP6Sr3exisd9ADAOjxn9GiJLeprrB6
jMPk7ZkSwu1TB/CN3AuYHgR65G2mBdiYdJFd+Yi2z2dspJCHLxZ8ewcwxuKRbBCd
U492jKH3F0EmOzZOa0G7IHsryUMgr/u7poxf/Zg8xTNYtbJNM1EpGHKnSxxYgz+H
+KwMvpnuDXl91TrO0K73JT20qSNgkBDfJv+9EhuqboAVhERSbzNzNzlnAWLpnGBl
Sk8SPUR9v37Za+0zho7qp+P8czgr/UO/XmwKKXxzHnXxsHMgr7Dt39bOHSBScjm7
+qnKGaemZpVZHmlHBH2ncdWBDre0qMeJa+8V8vpIe3S9NoeVeM+F6E3dADC2PuGy
O7q5c/zIEs+cnI7+fu8KN6K6AZOHCjCnKFQiQ64SnGQnVgEeg9okkN1YdcXwK0J0
YyMEq/JE6T34UkJMQfleQU2hnUgdYArWu8JtvN4gPhu0bKCItXRa3D+YdCG3lc+f
1ylv6wB3DK6UWksMUJGpBUpnCm4Iz2YDjXBRkm7EtV2giuEno0h9/LVLI1gphZlT
8vXK2jyAJMDqfSivKt9voCU+PjIBrkBlJLpVqpWqBH4z3GPaGkCqw+74VrIxnhED
dgv0eKS8Df7Lc/goppktV/3zDHEvuDrckdQygP+Vm5lLLBGUj5QDszSmDFwsmK+o
9oGER6/i77CtVDsWRXfe7df2reN/CHzZ8f4yFtArN9WBgU05FxuQvfYwxtar5irY
WEUrDAEZgWbxut+4ecYN/6q8TVdBNUShIpuWejiYDRH6ubS94+4+3BHnwG6PKkKk
nknwwcysbpT2eDeSK5N6SIHdklEEh1Iv7akFHh3b2hIO/eUGsAo9jX6K3UKWrPyz
B9bEVcOTRGF4MZc7bxXSe+/aOyjtlW+8rqWTQDCJxlwY9iTQIH0cHADnDMMJlYfl
m7K8qrcXwwBLSiYQEp7bnEyGQiMirAyMl4ZFaRw3C1nzhUw1nLNV7nhtIqzLh4sQ
hMOz5jUr4zDcwQ4JvN360AD8ZB+90SxH3EGeT0vVBHudDobZUKl5LHxvQWtsLJ/D
zcTfleY4vy+eSSfVXP/6ExGFOoyVbvGQq/pqjYj07KijWl4FnA0WE4blwerj64wJ
C+5/BhqCYNg4TSi2D4GMxtM34gXkC4/rf/eMWQzDdyszweFELXZOId0Z48D6RMw+
kBAwcrkXSzBToHhibGBLQzdEKea57RhQ37o32LdBCKkKLYW1amXVu2D8hddrhrBw
Nu12F97m03aox7biF7qLZa6wilAATfFI9UBbO+eXgMWa1k9FLP9EFTuvIcvJzYXv
FPp9W2d0HmGSM1pCg7Bjeu2bkhZ0jKY/W4jcqc5LqMpoVZ04s1mFL8biOmUqNSn/
IF6+9XvoY24NAPvzILXOUf8BqWkCyLI77us3Y5rRVfg7DC0ZTD8uG5VNapI/ogEd
WugYqdL/SYDvc96oLYBpFY0yzPotIkPt6ENMWa+550Ft0Z69xNiuA5ucrTDbFTZ/
nAoRscohXGPvzAZfz1a0chpjPJu5vatMXP4lB0WMi2YyR1/8CDCg6e/bmC/Ri4Uv
JcPVKvqxRWfs2OPWWbdIfOdS0/QOmWeV9/vxNRE8EDYJQpeuf+0zheQ4n3jW9y5C
wBv6IHAlxxrIyZncbb24d/U/cWfSH995tr0eRUznijGLE9sd2WvQCfWM4aAAs3sn
1sXUthrRNuYI7MBuQt+bxabbR7P7FL0t38Kx7WQGT8JVHk+uh1Zh3MtJOSBxXyCG
PIHAGcnSGWeu9aYSliXtlqiU3XrfFmIgnKTiQf8FqdSQC+egzck3gwQckBEBtoI6
BCQajy+2m2qOq4ThhjBBDbtyf9Bt+ZTYtZBsVm4BYHAlVryrNqqhxxxY+wUyB69G
LPhWqGpC9We00AgWH1GvsUspJWOgAnd8Nti1v0pRC6/kAH42r5FKNNk421ApQd4d
SzXT9nnkNq3Fg5LeDCWaaD2JWus/mSiCHdPmrIPNIEH8TgrKicne/uXeIcAxd3jo
HpRsg1KNMqv76/DIUuE3KcgCfbu1primfSRUZUqRuBvZbcVg2y45oHyYQYUQO3Mw
goadpK/8pkrOZNe79ZuiR74myiSatPMdG9P79CBKtqaFhfRiwmKjOhxedn6xRgyD
GIkSTMf5/VTd+j/APj1AjfYrgh+q3yuW5zWihyDK7rAAW1PCZQlXHMT2GjVT9yu3
07UXj4ikfB1HP+OS93AwS5Ap7HYD5XlomLgY6zGeBv8GU2TxAh/XXeX+0Nxliopt
4BXWzRUbNav4Y/pOLEoVY5741VbJsYBer/KPNZ3oFaRGWofhmeK9wlK0GaPWsKhg
IysObZ3D/d711F3elyKFFhIGCPwsy9s/zB9zoPv8eJi5J3px2/mJ9fKA4sI51lC6
0LviG/PRJdBEzSqP8RI8pE9r7V6qFdz43E3vb0A3HoQcJZsvJZhaHvh3we39/6Aw
BKGVTMDbkHvxtxkBE9mdAYtC8dtG6lU/plr2k8ncE6jnAwk993Zc0gXqfn/oV0qj
LlhEHB7xE1O2iIjfd2jNCPRwiPOwfF1tlYDUpUXFI/zxx3X0FNb1sG3XB4EyVml8
ljpLvQBpR54f4XQfeNaErpXNTA5WQps4Oi+hOzcKwtUgyBe3FPSelwNjdUAbVzcY
qtE+QzGzryrQrLZgfCrYLCiHJZUhDupHkA65XYFU4bELl8E50vpV4CRGuXfXPm0r
hLMdeHLOmGaoww5i83hvLt62aFcJTUNo3fiie471xR2T8FSI2F1zAkbpvXQeV8FT
3+44zCLPPMlRfFplG0YUgsMFCYonPFvfWSbsxquHe3unc7LozE1chkjP09n/pk2a
coe4mZdrwMpXglSHcS7utLGvpiriWB3ydnMmP17N6Oz5RpGU8BQYXLe0DtMna179
ToC9tYbfn2zIXNieT7oSL80w/oGBYNMnNAM0UhzmftXPhBdVkUjxC31Z9L05pz3Q
e4exjSfN7Gfrgesh3oWZ0Q==
`protect END_PROTECTED
