`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YcXmETrUhHKCoGLC3TTMq+Hkl4uZvR7LckpspXJKw6cc+jBf9QCfzPT3Gly9V4zj
ZPIaGM9kiOREtwsaxudA9EDznAlYNtqqftw8Wgoo93HhsgCSgNvS+sn6NalIRzO3
hpDz2tWmH+6UKYGS5fIxIzwzfYf3iQR7sRaC4oTOF6GNeOatPcK0PBZd3tnTXIMd
u1XEr6C9eMwOk5FAs8M45v4L4mRH8hrcOAhEfyAHCSXS0/uCyDnZARSe23/qfC+q
j8vlOFKOCb8nMFFotWAzH61HSlpEvxmfdWLqHLeJLbOs6Eq1Mbw0R1S2AtnaumMK
58gPMGuQ+q3FZryYo2COdpZz1WJMZ0q9OjH5eImvbe7TbVMI21pMkOqLfNiIpfKu
3ENgXR4J7fvNVWPFiSazEdUdn4q0kgjmSbz2z2ePwzJSvvsHyJac2+SPHXScbsrY
M4LN9WHNPc4sNHwqp/0f0OgHOiMkM7C+jD7NaiVlaUU=
`protect END_PROTECTED
