`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BP17TdHCKfb9O4gwnbKZZ4s2+UgQq792LeoAJwUVCafeFHc9zhug8ws62ZCU1wLA
TJGzMGSiiFnFStabiEMn3igZz4kdFGzYZgT16YS6c8727nxOrvIjJd4lPaujc8H0
LUzw42RGdxm/cT3RwXXfRzBZ+Z+9nsmmSnEUKCCZYFq5Yf8kcy/JWme0tDKgFGCx
3Df1DMukZzbPTYG0M9Vwy+6/1OgNKEdLYxwcLTKcPQwSraa+uZ307DxjgoePvagb
NgqDi9UYu7UZC+3IuVqMIozeJE3cwiTtvg+aHmLvjxP1XAk3JXEkIkLaM/AsvZ+6
U8navN73DmQJVX0ciJ2J2R6yoxshHjo5Idtv9JsxtJ61yiq6CDoeo4qwkSX0BNtW
7h82TWiuA9q+wESLWMwJ+Tcci8gVfuLW2r55bqFxKFnH7AEWCibBph2ZIHs8O5Eq
qzE5RRuqWlUhwP7hPbSOHw05+9V7Srtbzp5Wkl+ENyfPc/u4vgEkketu2nNvIqIH
18uftEIKw1gCJC4ilkYAA+GhlFopoVXnkmbFPf6VZqWy/Qzar/dla+L4FMUpfDks
`protect END_PROTECTED
