`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jN2HGcM4vhFXCBB/AfN7OJXRw86SkFtvupg4pvmf9EvhVY1g8jNvnxDbsnoMtEb3
XPIlrKjzy4XSR4Qn0vMUeNEEBfjYuY/E3/2dTl3T5ObZ6k4YI159FCXHjplmcLc4
CqbfykBzW6S4K0gQjKmrLNewK0SzvK0jbrogMFEIjMW29RL8O1TD0ZHXtNo7AZ2d
qYnzaZ5HKZB+7X1LdTFyYTO68DYwaBzSoVvJ2+2W0zuQrGtLqfzL5Q2SOL6bo3Bd
3e/rtJIPKXB2CVY1BfveVOOWan/n4ts3puafse3/0Lsf07VeHw2Jnd1VmSATn2cR
vrxMIBwgMml83yhcS8Dj5HQq81id3h4aKFcKbOwLuS1gwJ626sl106UO4wTOeUWX
T3SX0sWzoHgar8naJ2cS2FNemjfWp2/bl7eRy/IQz8p+lZOhqtpKXFnBg0OStrnd
VmshpRHIdfUcGSk9VW5ZP3ahHVeqHthARy8tgkSpnJmuFHcErFcaxvMAGtaL8WR7
t1pgaW55iUV4e+pcMeAOTNa1psKQ29Q7ycDXSxiCsZkmjS4f0Lwk3HR1n8Qf+j4m
Blq6dLN6B4jIPOKOOBWE4JFjRNal2LDlTsFJfKHaSULsGwQYf/77d5RZppszv3kw
Uw0oBhgnKzNy+REJBFRs1oiDwfgiI34fu1RjTWQkTK3np9wSLQfz5Z27SH6mwinW
EA7PyXqhPcZYRBf7wbLG02cLEJAUZzgUb44udn2tz+lGnpxoWvSI5Utq3QdjMF81
pudVHvrJP6c4bAZr2tRYJsx/IDdhaVN+GNDwIX/42jdXXWeKZgRSJaDm1irWv0Lg
OIfJAfRgZYt5PUMCLvDubzFPGeAC/Uo5SAzjLZhPnY6Cqv2eO4Nz1bLVMEyJHl76
JTyFWm/vPWKm4/LSeU+uaNqlr7np0sFJolKP3Lr/QE9Q3oJ4Q4PXgjV+OQhF7Tv8
79OA1Xl2A6lZMN9Pzda/LxDIfsyRxkZ1z5EnCYmi9sn70RXfNPGDIc9C8upPKsRV
XGTaa1ouIAIhyA2NA09oQapIhl9ycNodzrTYrdZ7LbQnen3FCf233ACgL/tO8hU2
B9Osvq2u0zOx+ygSTPHADjgQEAAe3eGTPQ+d/X8CXOhIIW+pD00zhVDSOMcWxQ/7
Z+Lm1JLeLr5tyYlhVl46tSXUH39+6COoCn0zD86tMzMFDmsi+z1t1DEwiEVFGw7d
j0tzLgbxvOYsyCwjtOOFKB0YR2RNDTTg97e8dVqNxGDCWkMGbZi+XM3stpdEZG4A
Hp9Gq5UqzAa64zr+rUZFc1gCNePWmVMCbgUS7YcCpdj5sKAZsZBMjkSAS5zHKz1g
yYvnjkFqdMAzSogfCdwMY6lO0sACsUMN6Nw2Fa8otqhPIawvBVEhp6NUyWLNMi9T
Gm/5wibG2TQbewR98TTABToPG4rl/JJNWTTSkMWPGyxbL177E1j8WDl0jNCIYR4S
`protect END_PROTECTED
