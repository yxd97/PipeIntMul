`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zuPIuofsJfDoeQ/2OpunlqCeRw7CbCv+XlVZXDz7WmF5tJlqJkXOZx6b4edWnNfm
7OXJbRUeQk8uMJ35RGlR+uhiZGnA13B4gCiWCf8X4T2QqzhOlCfDmgwMhjW9qftA
ZpspD1ATzcqkhXDZVihGDeCIbwv7UsjH0zTnkDDuI2Y41DGjwTGPM3VxcbKsl5X0
HAJRlnFG13pXWDyNqYbkPmtmbUsG1oaPyCdAbwqBQeAJSIqV/fJ4JK+OoHWm2ghb
hN5D2DBDAxsbIhdHEfZzmA==
`protect END_PROTECTED
