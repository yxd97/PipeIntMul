`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gzpSCW1rYU8aiwjWI+Ra8CaQ+IEeirzwr/b96gZ//aE8x3pwtUgp5mQX6MAlbYl+
EOTac+6M9K+/kzav7d41LmuwLsl/Dl4mvK09vIb3vqXEcoELk5LtTOkhYyfnxxr0
4JUm6HCwdoQbrS/fdkSeFo05dCOB+UPK0icCxTNmNWtigDwlq1a3nG7Kkc9AX5gM
jEZdj5qV49BXyvbyza5l4wV1yEueDxHA7JxGjyQaiYlNE/rzCbg72TF5OEKyvGE1
o85JDy9L1M4VH9P5+F3/hNihBvk2+/xHYJ0qxD/QCjMMne/sidixtK6zSt9jLKxn
NDDDudhuyVPptaH1hUso3w==
`protect END_PROTECTED
