`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f1tTh/GtnTxJbJ3kW2o2omkTVwcQG3gpeF6hIVjre78wA3UHdug/bzC91fmQG9Qz
wpG8Ojy/7bvra8qWGU1HKDamqX6z8N6d7kIhE2ecW92Mcw0RzjL8VhrJ5tjEW5d9
Zf7hLX5qHJdXPJQlURR6T3eWsIy6jP6H/HfTnfolOoj5ozskO6YD08CxzS0S/0pG
G8QwDIQjgbT22OPEsR2qCNg1OBuBgcX721Vp9Lvt8UHOKvgM9Qz4wJ2q2JuEyVDY
JtI2dF4wi+03WeXkoCzML6jHK/Tes4gf6zWx6mhBjI0GcOFXUyshFXt+avYFl4Hu
xFm3kwKUZEERzL8hr5L1avcou6VD3ErZtElSgTRrimvi5idVm7SeFxC0KlSOcQtq
So9se0QYQ7ZxvbUFTMea/ejGBSy5BDdCu5i6T61+5wcQSm0PusK4LOYaJ9/E47O7
wUukgVt3hhIAyV5qc3peJxD5FzkoP/SGSKtZwGwhgu1b3e1iztNuy0O72rXcQvZv
9JmdgPGuzQvn60J3UdIgWvh5c3gmxuLs2MvXrHHyZsq6GJ8O+CO6j+PsJ5i5vUC+
GUKwlqi/gw87fsUK4YyW+ahm3kKZFXfKm33MXXi3IubAS9nriPNck+fVFXMWPupE
BKjJnMdVhHkg1m9npfSwP5OolE3sgJBYYnDckWDE7BCLHovfmpoLnv8mIGY1dnag
4iM18zb3/L6gMDIVdbovQbTNQwMjkZU8kddjUIN7+w6EiP1rdAV/VNUrUJJD8C3n
5xU/QKVtUuabHbvimlaDn3lpviE0TkXSXN3z5iy0UWKprhDy3w4qKwGod6mFVT4a
wXNODUsEYkwEOtWdp6QtoEcwrgZklZOsO+3+I2zJnGgtbOED43WIWMAwZTCbCcr7
cOgWv0A/JOZLqseQzQtH/LH2+0Nc3QZtVgUMr9yDwdJZEfDjCinr51s5pe+stSF8
Kq+QmB2t/k/2h+wjqH8M0aFGbK/cr30+j6yVKscYaDKPkYZ2j67w/De/Zt33NjPd
fc3jbBibrDnqj97yKq/zVNnthGtVK3YHrZOuL1giWZM=
`protect END_PROTECTED
