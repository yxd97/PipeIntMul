`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFpjSUXHdIQlcvQx1tuEVLtnbSlsWUttXI//YZG9ic0YmRIdWG5cERN0t0e1dwEf
qrvRSiMflC5ZxCBb4x/LF4Bz565idQWPH1natIirwweJeQKq3kR2IcUzBQXcFLfr
8XxXD8CBeRXmh8fdV6uCr3rH3K/TeQlnbgchnh+OnAq9E2NehtBK8lIjicMiwLxx
P+YNHNbGGsAGjtvwCr5/1By9ICa3A8Jr8qc02aaIaq+IsiFklAIQTQ5ccJr4IxKV
spaUn2TAemFm0s/32nLJwTOZWorSRuZ/AH4fyg/MYCarCesVV+bq2lUJZSklNjrp
apLyIMqQUhqnIvVsUpUkJMNCM2lNooORBqD6/46K4IUPdAiXlRqRryR2HQqjB5fJ
sIV+O++I3G4YvopsrLYvgZINKhN+FEzBSkcr2lyAOcc6wMwRi71rKBinbvamIoU4
`protect END_PROTECTED
