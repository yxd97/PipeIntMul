`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lFKG8VwuUW8Gw2q7iyx+1GD8Lrq2Jt7yRyIbN3TTgHal/4h1Ox4y0ncS7tyNkZsT
0BeUtliNTZJnpqnQzuge/9UGJrlRLD2joolgzv5nrVq/PwVMMtWUIIvm6ytRtYu/
F/CY5lihyd76dZXyS8GvFOJtd+Wywl/uOHuVrPP3ycwqrleX+rTWIb+wf0ObFLy/
xtuACPL1jkwSNPblumGGy+5/Mv99f1Je0YfoG5kBu79MnrHPuLKxYOC3uIUJ9SDt
Dq6BYb/TnRFi6rc2Kx2jwszlx+LB4W2k8v6BS5RnxbT4gyiR1a/f9xD02rEJtAEM
xtsBinxDOs6KcvnzuljwxjoHqXSuXRsCcTqLjPrQSjYJ89y+0jLtMJ5v0WM0jR91
Zj3oMNsEHZZ6doz2UlqZuHHM1r/trnfmlltQaqkn/lceK9gB0xEPusug6Ly/GFa3
XyoklHBm1aDUKDpDLdXpyuZHUgM9LqHhePtQ2l3TuwuuPKSJAD5Gyi87Bstr+00N
chqMSnAK8Q0z5jlvtyOeTxfRsa/SA0tQpGni6bVQ+C38IRJLuJ0xhtRyaeZcRXf/
xwoI5Ujg3761zimYY5M7WA==
`protect END_PROTECTED
