`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dj+W4jp16Hiq0yjmZD8vM1uTwAnXesk3ove5rORuzF7vtg8WPNB2/A0u4FTjf376
sMM/3pzxv77d+vfs2Z/Nz9X1W4qZo7YmaukO8SsnBigIX3RxmMWrilXlb/bctLir
W98Ea4Qo4FixZDLPC3LggHJjrvpOdTWs6M02z05lBEmY+L89H/sTfoT29/1QHS7+
HfR1yahewgBbGhnqQM5DjREPZCaZsUROLLYlyNOYD3Ur2Dg21VAMzA+x/jXAdAT+
ZAtLCQbluAFlmOaoHgOEcAy5x6+ze74cmv3kL8BgJee46U6PR0i1S7A3g1gwpVt5
IirWFAPtUxnbMB+Ok3dhmPWNcM/980EaLLwICGDcdeMBjEt27HnR3yn5lKlIB2yv
aF1GXFeQ2hBYJALWK66mHBF4IZGXMrvTug1bRihm4z9ZBRGrzpZ9+fWeym2gmxHs
pQSdxabfpVBmi7sRd2ipa1apwMoszMR5EnIgQE7bR4L7hIVpQk/iWhLH0twfM6KE
oXx5DNe2WSRjzfA/wutmdCwAqbw5O4KqPTQC3X1vHgPVby1kIZtsdPhlPfzjaL+8
0P37PgvgIO5wqep4w30YeINvKwu1+O7Fr/YZ4Vz5xgpZMLWrnxwkc4QYpwRHGqMF
UuJeyUGjEfKG0cVlMHAic2zRur6mSBLE/EZzrZ2jhzE6o34GSOrY6wz3Zq2jm27S
yGd3TzLo+vnDbwOURAeWglepO35K2FjfUJiXy/z5IuW/FwgoyVeyoFD7Bvz5HpjS
UyPK+yP7s/9sDr8YrJuCr/Ijvj32f5KhzpIpvBez8j7AJc8hIOPXoMKjccNsPaRM
xEMC5jwCN1pad9Iq25MUEqJHrLSAbrGe/os8AktLd5LVDYrFj3iCQl6RLcPkA09M
N0wRT9Q0QRHCL+kn/HGdG/p9shs35iFl29XATnNPg4Q2sXmWI6DmmeYJot9TRo9l
8AQWEq7DZ5/TXb4xAPMBTmvYS5NlXz7kPEECSNYzuoPxqgaVEHysl8UzeWq7oN8p
F0B9rq8vlF962ad75oG5jTYOfNLu0iCFl3F+buunuyrIjLw9fnWnDf5yqGzxoDaF
44Mgf2uA0mPpWdJcH/6jNkMW2tbYQxbjXpJjKkEO8tNgaBLYbPDkoEI5keL3CRo5
Ic9JR3Q/3wlEsQlgmR58HliNXd0YKLPVjSmqDOnAfQi74lTqsBFOHUdnpoPswOm7
ZM4dfQSqJ5+KISRvOZ0A8PsusKHqBvGDkFJ/Ai/vt8g2Tu9+5nuxDDHaSjGOJ0fV
L14iYRA0H/0IyKHi72I3iL6aopLN/W08y4AEHIDATFcIUfjccoEK/W6m0zVxxlcK
ip0rTT7LKm9sy21f8PjLGDFyHg5bPcSMpWeeAzvB4IGeaVKhAlhPCH593W1jot0+
prt65rqwHydSwPnFrJyfwLZ7JzQ0sLeLH3q9nlwPe1R2KrHPBQzk6otob4rVAiao
ar0fi4No0QhkzxLR95dK4DlYz+GoaTmWPbI8wq4H4K8y1Jd9cBGOLryTdv/y99gP
iTovk+ir2V+B83I6ETHs7dPqQ4uxWBb5tyPysM7botdrBDICBx771FtnaCVAnf95
gU0qHmjRGteinpp3DnUJtHxDfQJdwVbZeC1rOJi473WYcGPU69H/1pvmIGN70/TI
hZvF1pPkotzxVMD/Zk85EYLBGzHkYaR9S5BTeNPS8ZRoPjUIwJIEBQLV7BhxJE8C
kl0/ZpYJ6N0aSjmOjQSFGQIvtLFe4/2+gvUPLtgshQt+Fvig4Y8msQQfwwIyUO+P
Ul10ZuMy6de3TlQsaFgdJkLAkgifbD1XYbpBIvZXRkK7fOv9mR7ftUWmzYuAP5AP
DBxXA43WcX4tbsEQ2S5ymWTKamy93nzGH/tco7UjQLkQxYEYlBxpxZKWpZLxlCsX
iA7Cp35wPVbtjiDkUZvMiYS1GxAcBxps+JPM5UIGU75SDWSAF/72A6QGHsIsXkGY
VPviwjHEuFpBLwg0yQraXGd1KAnx0UjOwsCoxxqLFHNLwyT9j6cyCSgUO3sfcRV2
N0Ee5015Xvo8L6AMuQVhDK5OgiGGmoXC3FOJSNNZA9rVBsIu/7coDf3piWdUl9qt
roaQxfmkI6qwv3UwJBP9S/omD9s0iGW4JN7yHEUtY64tDvIB/0/nHJdO56FEBw1x
KCmp0uqIRfeBwhl1TJTMEmEu0JzI8tcxl9paXBemmoDlfp5rsMm7O3DjBxtyTqi/
QXzCz+bV5c+LAfUwONeXqcRLZ5bsp824aiWuPMXBOZKSyEEYEgIVhvYOxlLgJAWp
5D6y9H1Lz5W4aMA9NJywaNyazV4xMZCGE1SBEyHntcUxD5vKI9ORWigkpyDADLEl
FxcAFzDCCWjFwRWUffhJrVvXLiITinZap9AV+/FOxlXUTa09SQIwiTlyYfnF0Lf5
BD1jkFGHfBdI1DOZOptuutAs7I6IpLoRhwACdn0/now7wD/oLv5PBsxQ91RkOFNb
E2HoVwcnUlevO1lie+46t23Kdu7vM1eB4rAJncwrDccWgDzOou2ovbrCZLwg8kyJ
/NCpt94fg4ipXE53isUm1Sn8dnci64E/aOvxpS+Efz8cFFF2AcxWFzBhi4PfcmUH
s/sY9mwPMnJ7bPY69xjbLQ+J51Z6iU06k01mNDNNWIiPBi0rOn1zJ/Wd/f57H3dz
XozK2LnunwseVo+MkUjb/sQiSyrwZurNW5l+3mJVUUEczFk8Y437thRUoNsDuZCl
PjCynNf8Qu5ck8SFUTt67zc9xHFtmGEP4tcFfJ1BiBd7vC5YqaL1E+ZiiEKOtEiy
e6ogToFKuiuvP80U8wxd7uGdN7QMvx9jq6lsbZt5DPMFt7LBzZqUT4YjpNsDMFwp
LUs/GLNujLWXVW2y9TwL/wQ1693RDCC/QlCnBtgq7Z0iSpXe8Z+bH7rouxg/HjFU
qjLSxkphiJNxOItEGIzHbdO3kicZpeI2Xg/2BcsuKgan2POKYDBLazxnRtu7s3Rk
E1WGXXbsij+uvihpE5ruCqzA8wl45y2B0m+P/YMkrocEOKSq0yh7ocCUeLfY7ewK
n4DhdtQXtb6wpRXRjlpvzi3gnYwsGrhXTo29MZwPxzT26+jqPJKQQBUy6zL25sOm
JNShAa8WrEPCTsr45FMvJcifVlckkcxS4nUOXrTA6aLZjAyuA/U1NEbeU7MXeeEV
tfHlHhzUuerbDGb21G5TwYkWM1NzkIgh2xYM1l1I9DVs5mlGiRA5C+4yO6pdSbrG
0RL4I/1BLxnjUDAdVaZRUGIZfkLgKhpBg+bT+4EIMVp+SP/A49R+Hx5TFWBsZq4z
1sqmxAgBBLXlKXnQbIQabriUkv7SZ4Ju9pSw/Io+Z04VaHCBRL5DypeG9ks1TM0h
+7o/MPXPlpF3Vx/OGdZJDzoL7f6P9ZZzqI9llldZQ07CFBuJKW3hYYEbYVHVWOSW
VE5RtZh2eiq0chqWIapIsmTadGsGAH6hiEiRHgdk8TpYz/n+vwfZZfUc5SlC3Evj
Ac3qf6gXYFO6uhuJvILBgLXxVeH41zHPDpa/usXvhsAAJDokqpF0L8dPPYkyqpVF
h7XCgiRh7OcdY5FgkJiNX1JKBYG05pGEIQhu2ygTkquh0qAj3bdqyfg2LX0NJxiE
yvmhzlJN6AOooQjJ2/+pwX6ywRsa4GPoIIhWjle2JZHp3aLfmvdx/9fcjtquCsty
UIXffkq2HsDe8UI26X+xlP4ICqOK1CR4UIHtnEInFzD8RHOvdAyPj4nNE5KiX/Og
iFaU1xuV+bApoXi/Dvp0DQ==
`protect END_PROTECTED
