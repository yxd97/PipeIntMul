`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2UyyCE33lBHdaQ0PPayZAYYd2N0zmH3w12jrhM62inPCq0ciEwfbjyTsLnuNM7Jw
I28G4Yzh0wyN8PlGxcRWUhe0upGM/WOx1efq+Npx/eGrBMFFyBiaIUp413HEKwOq
9yAT6mIhqNR6vU9No4Ezyc4GNX5Fjs93aSrk9YedScYUyv7Og8PACzBFugTebmhl
ZjwSBgPgH0iFpPRhqyhB2CGZ6/t2f/ceKbQvrYtM0i2I5oQfdFwmSZUHiYmPDsYb
8Vwzn/+uJJoVowQWqtI6z7Pfzr1Q2FOXNktQtCjY62Z3fO1PtAOvFVf+zRr2mh+u
tfTAsp050gtJN4EBSGxnT2dVZASOY2yhxJRePArOwnXpkREQFy8mAiCAkyWITbNS
775IdlDedmngdaAwrEOYFOabgf9kbAtvvtToTIKPmcnxUCzHvSMSpJDXMUWRG8zP
lwuJF5RhaoxNFPVIexMXRQ+asma81QZw6O2pXkysxoj/Frqq32ooZpD7axH0p3Qo
OFX2moZZt3WtGnaP90o7TFH5nadK+ZBxIOTbQN8iokAeO0CzIWEnffTv47IeZ23h
VSL7zOu+nTkSH5OgTmN8UZkIZ+liCg04yfy3qanDkl+If3+VwvDqBf3qk7pTp4bK
zGMtTNiTQweaStNpYhlG+IzvXNfdGL9JHgiLxKyt8Fw0IcP6Zdz+kxi5gQafKopr
C+hDlcz2lL10X7jLAj5bgcfvHBpTTYIApnP4G1Ys3mHbGV/qU6AMfgKSbilidY3r
3bJsDfy0Rdil/vHcx59RQOlDQuSysQpIzuSqkhSNzdltlmaYqHEaGgsrhNcPdmEb
4jwR/fITXpPwlIMkPL50DsCcrkPkogphp9kagjU5oP3Y89xUvVsCQN6fa9fqM7Si
hXWQdX2EzPRZv5D3tZZ1jifwRaj+DskcAwtSIMm0RtkZH6xbk7DWxWn2/LwIiZAm
e8kNo7ZhVimVYl4FSScEKZVJL6FDpf601YF3AYVyopVL2PI30WHAUHbrSSxHcoKT
S/dKU9+VBGVq5GATOCci7vg580VJ32HaOGdXFwevMxc=
`protect END_PROTECTED
