`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G4USvHFBmHQMxcnUvJHMjoVvWHMULXOpW7zsFl9eWncSwJ0xStZVA4bL/d2mlMGb
kmxvRrqiyiEyDgfSwTf9NIGzx1Naz4D8iREEa5qXuGZoqmQ3s6flZtplI9CisaAc
UVVG0j1T6J5wWoJTmr0y4qqBVgYsPP6jKifqK3sMUMDnzxwaRb/SL+48gAqIeIar
48OW7kmnxZNE4F+4gSeKm3yWxCP4Kxd1fXB+0ebK+VwHR46HpwSP2vMTSB88ZkcA
5GawmcOSiihiXLE5DzFh9Uw9nKR4eOuwOAvlyYJ7pm4JotjuxnMhxoGIpCOmfsPc
cBNjOHCbda3naGVpD0x24RHIE48V9g4cijzxbt6/dRawsMHQvioa5fqQ1HPIOZv9
rPF9ciVQ3Oou7PmFju69MC2X+/26yfbTS1xD6NXbAOWCLYKrAis9Sxy5POCS7wlH
lskym0MtmwZr1mImpOhqibrKluKxwyke+k7RNeghJe9oG/Q6o4tKBDBK1F0aBShF
lRP/BtSSjPIXIjkwkA8v9li3PusqVCiz/7F33ZSd86LsIV2Dwbtl+Rz/Z9QyVF4p
W6freIgYVy2lXjLkUwFIJtLjz+dNYEKxuWgf5G4ixDZZ58h//uDmzPJijq4D6v2J
r54AJzLtiCjKwYUW3GysWA==
`protect END_PROTECTED
