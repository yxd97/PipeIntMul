`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fRgiWEdhiiObCuQhiq32LFXRY8AbUbfU9zu4HpNoey6gdLNQmdF2nnsreFX0XKMY
+dF3XBnAQxLT6ofNjyUVbW20oqti1B4tC4p7rnZFb/ijalD72oinCX+T1i+Z4VLB
2yahdOCgH/9l+f3wgdmK8JDqmayTBsRubhIsqykRE8k6s5oEqhVK7KMIH6wwkvOK
sZF/2dkq2Twq+oE7xOWStk0ruKJYgLLvIWUHjjwa+KLbnaN/lLmy7NkW97k0MrkO
rEWHyjsBJL81y0WcfX9cnQ==
`protect END_PROTECTED
