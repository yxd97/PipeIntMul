`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oqi4kPSHqFP6YNubHUpKwaRUCyUovS9oGitdbjnbHPUzc3dEHK6YzvgWoCNUBttT
GFti6aAyp1M/uuyXfvREV+st3LWEcEjaEYPRl5dmGM5cz9sSNBa4FcHijybt+xlr
dCE5OJIVlQDRO663dwOV2wq01aJ7L/3UE9K/QiVeDIq+C9bmjgCEzT0LMoQpjEfV
8ghkAxXt9Jq7hvVg4k3EdhtIDn2O149ib63Oj8fmSYJF2cXxGv6Cb5ZQPKsOr2de
iEwLTg8mVWZUFf5shEX7XVtdKyuhiLNfVzwAIGfr6Fes5QzKawIScm7269k5xySN
qPWwFNquYFBhXYwA3ohgcwcilSwUxyqNU0YPjMm7xziP44UXHRRqo4mxfGZSc7fw
9owKtAdSG+mFDtCdgWHPCdpcQS+8A5Reppa0JODo+mzNa3wEx305pW+IzT07MOvw
/t+nxapLCf51N/x7mIaUDDHxBhU3RsXSNdNk1gHtOjc=
`protect END_PROTECTED
