`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JZzbHHY3Z5Wk9QNHgT8QGAnxssVz2bJDJAhKonU/KxpPq8wWdNMZkCIvbhqXQDMQ
f0Qr/qA10h5q5WkKWieLX6rAlWh+Fj+OvbluRA9XaPHnBCgEWbQFF7i4mqcHT2Tr
BQ3jwhsJVojgRd5L6n4iidcGRwm4OmaWjD4y1Tqy9xAVnqGuPdHZqd2brcY5CA20
ztWl2B4VhQtZ0An59j3wVEKwi3gt27J8uF7icHhmBa41CFgjQdiuY4+cmVE3//7Q
e76hdG1WIQiJwZ9rAZno1c5HrMZLPXv+tgXRP3SfJqDzcKex3bgPmrCXKJiw4mn7
YMpdJuTsJErSaQu4V5li+tN6zItdEZNl6yO+jZTNI9C8gbFE1EaSU85e26KqNd3K
3EQOwhiG3Wlpxr4KK6tJDk17EaP65y4Tp2ojo+QkURdBIBNttcBQ0U8SsIbr5oxI
RkHRIKFKvCivabVRdEaOxAZrFtcMEvbFyaGIlKcB+ViQr7EwexosTXX9UWdzNqNH
ZOxArhlcjS/ZTVEGdyDk6K+Glslqq8MvSjwo44L2ptIN+JSTy3xiv7WUaSlsCba4
RmqagHnOCRMwSlfOHwzNTiBy5ZfnQtcBK7hoqJN+3UuE5Grr6SfuIBI6BaqUTGfS
qi+xgyquc21j2Bl+dBjejSi6YZDT40KHnDp8heFXj2usb8VhHrmtK7F96Xwwaqab
+EVwz64lX5r/6NbLVrUU2U9H2KFdcRWIqu7udirlIorVaMZkmcQD7MCpTzUleLEM
iPaszZea8/JL+lPujyPhvA==
`protect END_PROTECTED
