`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eq0YgVJARzhnxEteI0du1tOXGnrbqtw8ei4U29LK8My8ORQ6RGliE8Hy/YYMn+r/
DeoKTYt1/7DRuE5taL5r+c9sM53/rJnXQoL0bH+45nRpxRhNseWi37SVlxWedy4h
9NWGWBRCgfLFpNW+RMUOHaZjYu74/WONyr3dKmIjUM11SqXgdfJ5NujPST5ajYLw
SOjipw+ewxO+UK6rornY2tM4TkG+ZuBC3gJKGpI4DwwIICk1JG6aXlgvtliBxqog
33fiSDJWYsqmoVlN/acPb9sPe6tUiGgoXeY8b89mMKaYR3laIORNmjU9IcDv01HA
GY50A7lYYFJOs/LUlh60NlA5n3fWMAq4C+4Q27vMn6y50yfD9DjB8iAjg2ZO00gX
w2y7m+gVzgpdfXFBeNsEv2nfklsg9BQOSV52QGlRY5INy8hpt5htMmVbyMSTQmZ3
KUhOeiMUGeGA3ARh6HGs50eHwq0Zo6cmUD4+y0hnqdGPkkWr/TlnOXq0lH3ggYB9
kG/Kpd3U1RNIs5kx8ZtuBAgzCZjpZHnZRU3gV1HlIKQTwrgGduwqUb6j/UvGE0AH
FMw3YowGjlHZa56+oe5oG+nJJhvVyvOkUbb14XREEYW+WtOjPvg/pWZQqa501kni
GTyd/nGbSPBwTvD9NjfqTQvlbONOkAlOvihRBMN3lD0yTaRuBeNbjsOLkBrkt3cV
qaWS8jibVkoICeFb9WPjidBl1T915KNs1a0fZV0nI/81fMa8sNLnR8qQs0qOrxfq
hWX8YqK6jH8+7hR97v9zcCKGAOyM+81gJSuCuhG+tOwtV99PQ5Sy9w8FPS/92Z8k
b2smiODV6yLAzrpg+Tzl5AvL1jJj3Q/hVgLwgkqFKyx9TTOxVbhOMYudwnyU7lEu
qalsLp8ApkFmwWep+6x0wv3K6l9zhWqCFMFKwag7fcyUX4DKBjQPYqQTwaf9ThiT
KroA5iI+pu+jpN7yc9dYHlyi430lOpc/9cVr4p5IOhahmo5i778KfGxWDcN1EwSN
MDgOvBbezgBGHxTT9nLseByd1TBGDCRldsmzGZDaYl8f0N6AferWKuasJPNKVpBB
fveY+Hs9zjfkjsoqVprmkpZYquDDG1ZZNacxaS6ALVLrmajd5rxDjEQZRutZ9M/6
bd+IBSC3RhwoVa7wbyK/EySbNdmZU8+GFWzd1TKM+xEKzg2Qgv+gVIA+rasmZBhK
M7rL0sVN07FRK/fVc3OqGRe28PQr6DGp8MvfhzddMzMh8nqB1OuKZGhWK9CheNNT
vbT2KvbGNX5Jnxxk+eB46sEn1mz95a/ka98YA3ZoIQqIxsNfLUld+yTKmKK++kbo
3R+30VvjlLWcQ9LrJXhP4XwaZ3BG3T2z/iBZMK9kWHfmLbK02gPlZp9/WJsh38LK
wG9mypCf2vIstcJ+peu9RTaChAJNTVfXIdvgOsiZJPXjx+H706a46z1lmGmasYfH
NyKmEo61uak4TAQ2k08Hb743N9Q+8cCvW3lPwFq8XX2VkX5OPrezXV9kIlbeeUN1
ueJzHU8a6ALmRul1oI9F3lvjSX6lx3idgndiLDwB0Wvqi9YY8U5KnrbUDzWfpYRv
fwPGP4qHxkcZeALL+0YTKoJCqTrvJPlqbuSSNjHnve7+RW6CU7Q70wWexouzthiP
fFijmgDkLj1jsHn2Y23fut1Nrk9cyaAmSZvxCsikW0K6HZrNFCatYsJ1ss5APB15
5v6hUjcarqMb/hHQOcS23NKo9j2XFAr1z90rjAQnXDOgeCmqDMgC4NuuI3d+U6dv
Y/5IjT+K1b5V5/M2qSqIfLnxrQJO2nauW5eWtRY5xADXTD9XkUk8/BqdIKnI+KPj
Y5K3vVeTkzgylOC6ph9Pkbm7yq10Z/uf7A+pVvXRYwczW7iGCYJJ2q8pOlWEAhwi
zRYgrCbICuBMdxrsT8nysx2RlIctVlr/jqEzvBr2l0g0LH4fWv9nAmfcdUs+CyDW
IcvQdZkZAW9QaQL8+9uY0cC9KjKPjwwUq+NaBuJ9LqQjT+pBVO1I/O1Coa7qxwNf
oiECds81g4NfN6ZWc29p2d2hwvzY3BoR3HUE/It1w4AGeb0zAFJ8dgmR+Jdpl1sX
/nAxTkMlOp3piYE1z4ibS/qRI8sPcq8tm0wgzr+uFG5t789KCnFsfhS5jRK7paiA
R5WO83dUAohA2uRcZscHVDe+mftXUxOmYqcE9swHuAqvjVKX2aHFJzCQuu9/65bt
Vqwvn5r8h/SuHSVwQh6QbukM1Mk58W0mDULUNaQcf7IkfAvUv/MCoj9OKDMGepmL
R3LEUaa8oQUZwfDHzcdRWTAh1mIRtYmADUk8ENN33/9ep0othtQUyCpJek8NHIrC
UZM3ri/atmF+xRfpYutRNVrAQRfTpkMwD8fJETHBNefp5Lg60/LO8quGGDTTSgGz
k3R0+kn0d0zDC9w6eaik8S3hb057tOHNC2IWlOvdAPYsotW5DoD+eIfr1wedltiS
PHy0ac9nyyKsevsV3M3RPaUdgzyVrElUZNdmu7faZtwY7cYmvRu0jZBMadGf6ZrS
h32KzC/xMX+q1VGRZX+VrPxfnTPp0Wt36qTRt/YEo1IhgZaUVGg/njRY6xzkyib4
GzPvS0KQMFDUOVeprEKrNXRWRhILEVOmc8jrkS+fIxu2e2/Up0d5IbNSQpHB+YpM
8peOcPt32GM6nM5D7lgOoOXaQIa8zR+CuqItcFbNxcUhCWDEMGh3P3d12lFWHytz
WDJ6o8O1uwllxNuuBRny7lBVF5zQy9cTnsycoGa+dL4PRSwYRgs/dlu/sQ3emfM/
WDf6xCddY1EchnTwGVJ2YsjValHUjQoLebEDFQtjZLImQYgg6aJ/89/aCSKu6b5Y
DXfJrgAmI3IObgSvxJ3I+zKOCblYbgghjT1I1DHyk8yc+y3hR6eJvg2JwTvL3epF
1m8/nJOaGBS+CANUKEAa7O+q63dcHj56CgATRbv+gcXywl48AWoLwbZBGEeEhiXe
VIljmqfgV7xi8j/8zeEyMUMX1Kpk7OMoBQOfnoqZoG7gf34o4yI4On1s7YoUOfHN
yTInf9IpSgWq/+KIALvdpdd0iv/Vv4RVihbXAW1KMNDRR7i3oNBuZQpnCv9MGPaM
pl6Qhc0pzEzBkMk/BAvoZiE1uXFgrVyad0XXWbraSMgQrf4CRgOkbyUM99BWq8eP
+Onh6LhITSz0znaLvbiJLWha/nz+/d1RvtTDHxB8Hw4tbnvKEIcKdSM6hZcZrWA8
rudV/vFRQIqe0TCOnikoEX24FDKKfVrLilOpZxANPE8d0PL1xz7SnuUm4h1PDsFp
yraaaYR/sz2pZdrg8JYd5y4onYriHCXzSfgDgIlmYUHC8uTMlGhS/udblimvb7A5
j1pRXqhucHuIszedWK0oV5vV1qEBo7kH71gLhYTjoe6sxOmiGuY0n6DIRZX79LM6
aAWMm2+l+4N+4qeIkrXWxhX7rp/3QLfpFeXsyvhI3j4C/WKUY7iAcQMGfG0zCDKh
72dC07xZPcZ6x+QmUX6AinEHRkjEXeonuCuhHuAlJCaNZSzymCKAQp6A12xb4lvH
5ZPKpSfMIqRABEa29OY1E2/ktElMmCSvOv7e6IKaBVoGgAoYH6fLDpSTytNutarQ
QYfVlfujhXM47vCC6vwUt55l3PzCBRhfk6p4xS8drgmAiA+nyzv8UXcAvKDGaopU
C60cmFrf1QDPwDEWl90tCYY0EcU1iK599PX1ByHCoIIzzZ4GDanWpeSH/RAvsjQz
yK/eU9RHD3vpAjbyBrBauC0j6QaHA4J9tFF7e9wS6dKvhhNQLlB001s3y0hETvsA
zZDDSbBl5ZwL0VTROd0Es+JSb06CqINFfz8Vqi8vH3UxxxZCD2LoV5/HMpFvfesJ
v/Sps1GHdGJZ9zlpnj8YLhvMeM+9X0MPsGNEvVBLDNsQWE/NhGQcjKlrs/wD/GLb
a2edUSubEw90xo5fZ1iOKuHv43CUFQK0wZpBihOtao50kQPox/9G8Z6ZoparHJue
FZSFcbQiLjY6hwg6nLEnG94lz43aw1p8rJsSWKulXdw1eHBZZQLiRFTANd5MCF0Z
TN1ZZnX7sbY/1YNbdHPHWuiSZpasxmV3KUVeqLS5hO/LNYINZeSdCB2USCkkmz9X
0ksyINiPXUmVuOHepWoFJHiSuHdwdvHI6MFovKS/BbCRDt091FLZvShLou0BSoBV
Jl0JtzBtl3BnTiWFa13m5K1vBWJj7n7f9fZyBG5n1aidFnDHaEE91dDfpKLPGOMD
gJKUD9HznjNHzCyqpFKU0Mf5x1coeO1dglIfdsJT0iYK9ExI8+X4J7T3NICJlCwQ
fvV3eZgIzeEpqz1xsIAHd7z7KpPEdhjYND4KUK8QfGbIN9hOGahDkKSLmro55EXi
ITnrUDPFGJdr5Ive5A0BJlk4Dqz3iirAMTh1bfiEFJrGc3wCipRRMNm8R2UuNhrV
L1uGUOCeb8nAq7+8TYEB9BffjWFW2FhhYT2y1bL4k37rp0wn7nO+qZ0swrc0li0g
vBSgQso+zrq9OBAExeP5IwhVgeun/0Sm+pE9yekykW53vXYpeA6nWLrIghxXa36g
aawQ3hRzwv+a88rxRZJVShSXsqJZHei6NRTJDGkCR7sx/1w/g7fKy8Wse6HH17BI
lTt3alIMNS0eJO0jcqT/Q1BxanJdtgmg7yH0IcR2nfJNxG8qQs/zNP/5B19B5C7x
Moj0Kb5hq5/WQ8FEY0WBrvQ99n8j45PURt8SpRjpGTHO5u6hEPNZht+oGmdJo6kz
R47v4r4SDm6NfA7EpAHI2TQmYzS46uWzM0IyXxT0hVEw0lywDMqKgPdIwY1/k2Bp
L52KKcEEPIqUAsSsw42neQCToJWljw8ad/4FWp6dUYbLA+UtdpG5AkpiQ6dId+gL
B2zz7kooTsfz5shhtkq9L8enoL7aOhNcLe47lljEk2bCgmZ6KoEPEEnnYTfsv1Ys
Tc00kaQX36+FXSiTyA0H0Q4hGOFRkK32zYl/6e04GOtQsmh5NhtLlBdXqmUEEtlg
uTltppr8Obz08HPayxB/4Ef03VpFkwkYr1dH0pLsq3NnQvvlpmJNxxq7cOkHbYCs
C59V5waVuFqJwX0YjwMx9pmcU4zD6SzXqNr6YixxwoU4xHIJREAYrZu0PGpyX86V
hbnVT/2Ehn35Vi6f1T/huM/7pKHLZQC+2xF5UGNwacaHkcCzhmFuGCqtrmaurMZN
hRFe/JS+UqFTo9XO/3y/jooigdpgEIlHOSGWZVPsTiXVkk/f2tR4O2qFNLnoYWZ9
9bQGQRT06QZtXZi+xxDEstZjPWLHTEc8KG/BkaqV7ZZ0dZqWX/eOpifSMA0KJ/Yu
hXksgA6zk6NZrOA4dLJ/XYcqX5bpKfH4yJ5m8nqv/uCK17LzUmAFlen4Ld7pGDxa
4nwQMvfL2vPykIJkzIkQLb1DYnoieQjdIc/XHwPBERIrqXW1K1dIoPy3xRLYsn0R
RgVVpF2f9HXRmt86M87Qp0gnTbkgdaqR3BtirGYs/otWxjtmhC+oKKPYXPPMx9ts
ucTGEtPuFVR3Y3zSJcDjU4T+Ez07FmUfxVGo8vIqUyggNqmbTTRt5sPkkm0kbeh9
gj6cmluWaiMFGxHrAoqsTQbyvGQB7P2lseP7I5eKPqTGNXKknqwDfvTGioo1nsq4
+RO4mvcc8Hx5hPWiej/IDGRbXfrkGg4Zav2If1MfkXt7PWGXeIh0lJ2Kdj4I7qjr
UNopWIGBYc81Y38F0OKUUIcKxxhMaDc0b03oGxfdfTlNIqybq+phhy98KzpwQxr3
zn6HehwOTgedE+AxxjNuchMfYHfbWSewbBK0xTvv0x7cLr1Gnn9yRovM0hKdm1RE
2tekJF9VMVbkiAPO0DipX3YbdfWa8M//5da92yVcNay1F40ZnCikkOcG9Ho9GeUB
2VLm78oi4iQ54vUAqIMUmzCFM/yY35sLcQvM+S5hIFC3OFmw+WMsA+lm9SWqHsLh
KC7WRjPI4MdmGMr+T164EHvNYRmPcsih9Az6ycZsY0x1yxeQcUNcgT7m8VHwdYlo
NzdOinnElmBODPGfV5c+pQSIRucaHermdqdzxh+Wvk9x2/2c0y4dwQxPkpwcn1di
0lvvuKmm2KsvVKaO5b3CsEO+HHqtf26gMnzSyF5DFM6o/WCF9LR6L6gzyHD6bgy9
3bEefCV3sxKT69t+zRy3Sfn6LvVVsmbDbZOXkfXUneebyz1/pNNmbMX8rf+VuOtC
Iho6ie2TsxBH3W++UdR0Qtz3656GqGJxjnE6g9+c6XIFGzEcbbOEJwJdPugAV3vy
ga/YzSTS9zMHU4su5StxISyvKtuJP1KmXVGy2dQdWAAbaZavc1DMen6f0Vj7AL8U
x4NqOr5YdpVz7CQxHRwyhab0wmAYEkKOV9XS0YlChA0viwD0g2gxLc2EMu6cMok0
hlWEM7Fv6+4Ixk5zOCEtAMCrTONWkgztSL2LYoCkeJAwBaNHEiJjzRF/wSxoOpee
aoarDCpYYn1xQBYv6S56+ip+VRgZP+2JjvETi2Oor8gadARhl4iQYDB3Sj6QH8FI
Cn+W3xpzvCu9+TAbeodYADLbw1ME/EWXWd9ITGm2ZqgaoAmBir0dEZcHa6UPknNY
hrb18x2xzzb75gJntK34bmuJZ4cAYcD0vh4y7LgrksETLM0NdBf/XaOHvXgEpzao
o59niVYR/mMqdJvD8X2mhRMloNyTjoKeD2ZruY0Q57Tkde9jfV9wLB8dv8PYvLrA
hxDTUtzsV1oE7hhusHoDs5tQUkNPJ8HE16LgdeW+lZ+BONQMOIHhlkPrkZLzkAaC
aSjlPHfkZxpgkwlNb/u5MzpAuhoaBrA5XiJNSQqTo04O3nZw6n5msB7MJYG5lU3Z
Amb/1SM7oQIE5OHenznaow6TpCq1XSwI4IiFYxMNxPDbuMP8eb78/23zfcffb2qT
STn6UP6Hqj/F+Vp+Eq+OgXMw1Z/GnRvR+m5QKgZYm53vhS65vLAhVbwe5ftBNOv8
NUg6iDi2IxfCO7pqrFZ6bRvOL87TrI1ta0UmJsWnoTdjN5O6ZGcTtSNfsy3eaxWM
Etags6ZzKaPDr9Js1HLfYgCYYhBfkj51X08l8urS3hkIRkwBzjZTqKgjBXWFPJXv
6rlygrVfAOTa7Zh1vw6meZ21uWfdaVccWKOOdZZtpLvDBKPLl1LbGZ0I/UcxdUIk
1dWlCsHJENZ5zUPEsEG8I7xXETv6ksXn7QNGrpMdGy0610EeiV/mpBwYXXxUgIWO
Ib313k2Yr6q3nDe3i57KknoUIxI0wZWzyyYhr8sYqsjdZnhxfN9DcYDZz68Cn6Yx
Kh30ZT7Jg8MTu+AxqE9aYgkdXejNwyyBtNUqQOr0wA9KmVS5Cmnvi0Y68mSsHQR2
aSXaojNg9NvfENVkxy6CmHyp8opsatxSUDGFR1W7KJcNeqHSVbLUE+qbA/AgGFqn
lT/wc3haurwHeUCqKREXHkqhuV27MLfwrp7K06wMRiVQNhDZi02dsbX4zucK6UMf
AL0ZhNJQj3kUnwUFcJD6SET90As6gcG6uO/khsYy9OX7OxWwX/2SPV7ue5T4XUVM
0W1ifeA8yJKaRzR8tmJ5ouf6Ihg6+l+N4ectoxuF1EqrAP6hFlRH76URVTkMiINM
1KAhOKfhhG6eboNdqJrNaSZFb6F/kz59aPDNc0R+Gevw1UalVWpqbBOkHVc6rFJ2
l9dBxmw5yWfa6MUpJ9RsriqoY7FqeCDdYurkr0qDJufACl5j/uR8+PhEkjhYmxd4
t3DvCLlbZLLrEvV4EvMzaJ9VlE636VySV1XNLBDKKQFI5QEnLUjhj3XjmPpDuDKB
dTyjZQGbs2O7+57fUX8x/i3Kp9O2u4jhDvdIIHxMqGKj0iE7niYCDSvbgz99Rx1R
xZmCRZ1lQDMF9dG1VhpwugB/CNnfZ7wonFKL7H8M5OIcq9JZ1LuKZHDJnnHq/W1L
y0pFCnGHblteTq182ue+ra+zi/53YW4uurQ+em5Xmtyst/VJPRsuCvki9hH0D6Q/
PWHjOMVHPbHfXrF29n2kGhZyGQmaR8U5QD6YBQ0mwNufYbuzdMGEXlsOFFiZfFPe
lhbieMJxhGqLRyIGtdUJexV1+sOTqd1+01JOhHzvzXLV3OmMxTb5hr9dyLaR+yLB
CE0XXShFrUnvLNpq/8me5hcZ43Ug50A7YX9O3Ae0QgvK94k/Ae/JvaPzH4U95F0i
ZwjmRMPrfEVxfGBC2PdiyMQNqgeND8Z0uPa52xtL21U3sFUOp2WU81XumhND5O//
bH+dAUi3F+TvRlBfS0SukKxAlXlumf5wdM+1scsodeP01LIxPTmltmlLYK1NHyzp
mtHKb3VSlGfOHX7iajv/4j8AgzwkNSOe7YH0LOysuo8qRDdQ4T3SCP+r+KW1UO1L
x0h/8c+ULL5Xj5G6nAO4AFnkrQTCgnnHCCgjOMdXdmOq3GjmOSkmGfY2IX7vGpgx
EG90ywuZBAFDrcCOpLoalCs7IzxEv+L+yRZZ0nClZLBrZWqrpxdIt0H/UNwiefQX
tTV2io3sLFxdyIpJpb/hQcHUDX2oUz8Ah6fGCANhfVDYx0QtnC5QtYBkZFvQVfTU
iHXQbrjo5CE/Lw5tjuHOyP2qZqeA5HcOIL2EZts7KVc+SJZQoq2scQsinU6Wx3X1
j5fBs2dl3iluXmDtvaBAPMNyI3x6Vvovpe6MyB+3dfMG4UhfE+Mn4ZOXco30wjsQ
xnMilrcyV5igY8l4h6JUSgePmsniDctG9G2WixauKprYnxNJy3fRZZNLuLiehb+f
q1Z7PfqvolZOSyHGtApE3p21HUTBNNaCTMkisBz9U2D4btVQ8cG6GFZJcbQDyGPE
QY9qh6Xebe2JoPj2AHLR6DIgV58xbI/6O2utJCdfv81TVwzF35T+YTwLe7fUhSxU
lTu9VFx8/EAydTwu0C5bx5UVeZ8HR2CJWLjm+JUfm8yvfZWXQvi3eD0Fr4V6BM/L
BRTGUqmlccVfWopOBH67YDtb7mHG/P3RVW8qkzoL3ujeeWleZPVNCLWCYHBVJwDC
l/qCzp9lcv1rVytimcoRnzaQw4x67S9lGJyBGYF5kFd/Zxu6LXX3BjNroIhGzdl2
8evIZsJhYBhC0GCBObO7RKD4MikqsV2vS3TZ/lMEvWCC1FvrEv4MzNqLssjDmAVi
MJG5YYylSGKLEeLRnt+n+Dr5rSRJB+FfZJ9pyLqTj3kor8VV62C00bg6PHDBxUeS
Vk3dXIHljdtTsaUz6HmGDjO4ToDTYQ4Mz+1e88Znrk4KkyXZx5VbIUFdJ0QhQoOH
7EPTFxAZUBVQDvKRt5ssi5l2kSTGZIFB4SL+9PEkBq90sZchczzAhsg8jGNpV9ov
fSCJJznC1O8TycqEo3iUV2x1rsH4brKQSBTFtVI0uSVnb1pJra8fpl4cNUTG8mdm
kRicZSYS6N9QuUtG1KKaIE6pSBeXz3lW5z+8L89pRSADiT7/4IDhU0wXpyreG8xq
9eUDZCXBemNT+2zsovz/81VczLBBrJVLjLVbgcUlOF0WHiRjDrikTOXtccaRCFST
Ul80T5/Xc+CUEnSGzoHeh9GhPvU+etjBLCyMFUNl0vmlPeklSP5kzxUVB1JfA4if
KdliPYDmDUkNhN9mfwNMhMvnYskKy/4KenbZxzs/gLKjzx1C+12VsPDl8ol4QfL3
92dMObaY/vadwnh2A98R4x0kHNzElS2aENF29YwMY5n0ii/wAj91GSlvbgflXVGw
BGbsY7l/3AdIENERSxWpe2Qnc57wlnlFvAKnS2cQ7xwLICUAYA37MEHsKlfBGBRS
4gMwZ0xzvGVgsjrbyyFO8OAoIfI9JAz4wU2HGupgLa6P7p4ysnSbqTDZNDJPyWRB
bLo4s5txprTq7LVy3eXiReb2w19N+qhcYOi2aoKOYqxsRSS14wiul9lp5r0V+omm
3nYlByOmy1Wt5tjKQn0O5Q8kupiwi4JRK71x/qG1IEGZ8GOcYWQj55zBnx6D7n+T
YP6pr+VX2IrYbnU0wVsU2DMFYRsNiZvZ89Tfk26CWSm68m9YpV+0UYtSKTClVIhZ
yVN7OurHjBm3I9hLiL2Lq+IeA1tVPWctURr12/5/d+RJbOJv6aEnQMKKkT/xRoEp
segQZdENTSLeZoc2qxSWzjBb8ijH2JDRM6xCCsOLYKsVfnF/30Paej3iShDNtL6E
ydGYIUkAKOWREj5XpFtKwukSSPM31ofTNgq1O3OdUaylWzZM8gx8x9T1tK2cuUEA
GEaIQsBDZIS599O7U+74VwEDpWzmdNrGGhM3tV+yTJEGTsjdnATueQySehw6DCyD
FQNja4ZuyxJhdigcLDk4WMwpd0fbHoeUnxpaL4ISWagBgDJ3y2FXb5RlisAn1I3c
jqO8K292EYuqu1ZOf64O87IU3tbAfp7njskg2IJPHNaiGFShOmBs4+UDMcn0LuXq
/ctjnci/TuZlV3QzU7O7ik8tgcZYxvGZeVhottDj06Np+JZ9LAQUWXNuoGA0z1+j
9xKLKEXK/e15FwZrJhr23E/1d9xC8X8Hytp2LhQFrXiGWBUCAwhSqfaoVLousiL3
ZpisnXL7VzlQrQqz+y6mZVUOy8PVuc9RDW2WIRbkS/N3WzO1stfPJR/9TCSdeLYt
OorWhqSVZLz/VMQvcxdHKHE0a+YuAv6y7S092usRQqUOhAisFj0ZJz2Fl/munciy
yF+oFJTCkxz2m5MZQRjHUDHolWJDKsptL2Quw2NrP1v2z77Tv6kKOAZse/5tySBR
DMcJei2+gddqMBEgmj8oapTaGjVOH16wvknv7X4UFJDcWf+5OJJH/5of24u7C45C
7S1SL9yD5PC5Xg5dMhov8uFioPSW8SncsL21dMBgd3frAfA9zspaDt4cVVAGDk/j
HeOHBPAsKd/cTLjofNIrTaLbbZEUiC01BKHEOJU0I6H9HHkdniwf/WfaFL8daLiP
itL7CHIzvid8bS7Hicucaztn+czvdWlr8Ye0SjecMaN7jSHzoXHKeDJf2ZB9I35t
U6TWsMjykc2HzWFUcYf4pEHkoVDLbXMw3KUkaOPfsAzpGtZxenaY073QHlAakMmj
YubEBCrKvEmamjMhnODcyA4O9Phcdp0hPZVjl1ncdn9iKw/nvMcBptJ7xLs+PG/D
C0B/jRQOWzyWW9yfmYzPel+Iuuvl6PiPN6/zxcSdugftY9tWai2nChcrm7vkmWBk
I2kJpnbQGOOixEL5j3M5qrjdo7H9FiZOqE3HPHir9GQq71FRJdnbDiEW1ooRoOIi
tK2WUPuw3mMkS8JPhTnlMcyL08AsoxS2wXkxftHsB8FU1+cqeeSb+bniia1HX8uc
0xcqNC/+qQrZT+9oeSOfKdu+uGnnNumM2xR/fJqqBuidczud3xp7YyNa5UFjySoA
jrm3PSyKlzxC9T/4JNmmocVVW73RBGcRGi9tsNB+6AQ34EOjbCzZvLBhXhoED3dg
uNP/JopPOpct14gKD9OTxYgBwCkLgrxYh+HexhhrY+OTly/Xyt+COWn+fBSJlpqe
Vt1uhQQ2Lgv3+0LET/VvEL5SUQd44fM01FEpPoKUVrw5ufJncdrK/npuAb330j3K
TBqobpBKpiralxY2Xrl4as/D6uj+OuOgkQr4SysBwzLa0xGntWbTl/y8en9OsxR5
+VQl1V1qqK/in/A/nwTIqINU5m7B/9GTJ6FpCgLWwlrHMeNw3JBwop0m/g1fHi35
ceOpDQNB378AydtDaOwrgWZNcgSChFEHRq1JmM3xP4l841i+NC5CyeayDNFieT/y
atipa7T6dVpOrREVNK79d1T25R0rgJYvUvVkCbVREHUS3YaiVp+z+0dY0Kb1uLfp
1h8iMs8u1aLpiwMfxDiG5c9/BcvPd7hbcvGq9BxFpljVCmZsrhJ9DhYae+e8Oh1g
KdCyHne/73n8RRLF3EZMVlv7p9ZAgIW751BHch4CllpDLGoRK+oim3gEpWZOOcv+
7tL/yy5ZVOzaNpUK+Me9uz6Rmcl692//G67lOYxZzt5HQoPjjs2twwaQU8qk0sQX
ZgQZd5pZkjQYyy2fcJr3Y3Rfrl1h1cyYGCTHlgW4z7xJHQgYCaYyu7fpPzrLwxV5
3sOk1XrlVoS434Q+BQ4TarRtOb5afheI1vupffvQeeHV1IBG9kTWn+g+q87N+LaD
ccKADTXA15NPdG0x0pba0xr+uLF3wv3Z1ivc0IYVw7BNXPtgBfddQDs0nypq2QAi
IdCFZ8VIGkMyzAMvxJq/bVgJzRAYbJjR5ezCIc6+sHWmFQi79C++dYgs9KL7PeYK
/r0RzxCi77hVz9GdZc4nYCuQRbJGNJ1aB7vu4tvFqoCKrus+l25HGaCMoPLmgrBC
b8szyDo4YilfBknugStDXvEH7wYkZ8PWEJAEc3prV3T/MXV6Q6Y4s20UFEZ95MrI
dvD/I67pF4aDDCYUuXd0w92kZgz218Kbi1+YXQLpi1uvNHjTzHB0i4egmRzC4onN
IYtlosqUCQVke4gyoB6MKe5PHnAOM9rpJ3oQBRzs+hMOsrSjSf39tWrcHlR39DFL
KBnjMraQ7ntmiydbwwfY3kWl6tHLvyFX560KiQS3VJaX7fvQJf6hEh8dSCC63HUU
MLPykPnREIqGeHIc4oK5fa0dSP0dX5wHT+bLN5ShkPnmHrVoSyjUDKl40KZ9PD6o
KbS2AF6vbgMRNoGlImpO2VCPWZnuuaMkRgfyvuC6piFytbJ91p1Kw62z/sBU5QzQ
V3Lxm35A6SD8cuVjmEcOEwVLiWl5kFOaomGjDjAYWtFFP1Ujb8K95N4LxhPkvhQH
uWKGtQJHU7tthACJ19atyTh6w0PHC/9yWC/S8u/85vrBJMCVO881Cg1MK8IiGWYW
omgA2Wd5mZEVSXa8EDOKKfw74SqmHPQDG/14MaJOwSXznStyxgQ81Jj31UMj4jwr
SG+noxHO1RdbdgSJ7ZYrdTOKSL76M9mgocMc4FDfu+1jPnlqAXDMLaLyb3NEVgtQ
Oonkopi8OBYEH0Zd/jdaiiT4P13L4X/iiMygAB8ZUwb+zEp8LHwqLYgkb3nzix+f
wZyA7WY0cMJnZZeR7jv9UNNJ1ZWJGbUymQoowXZQV6gwF78lyReuzeDxzppdtq7c
Hu0X+mxoHr9rMJSjS9beQAtGCyqOee15UW6pTUqtZRZ8oggKvjycvxoUmrm+9ocG
QUj9iNy6txvi9wV9YCzaKm4nbqroPV6hMD6wySaFNR4xyeg2+WjxE0usHTxxqbQK
pWhW/6UyWL7WQG6xl1Y6bFVqYhxQAp6urunRY+eZR04mSxGUGw75v4xrCv1NwAB1
g/5hNthHb782OcCtWiUe5wa85eISmej03QFik99N3phaSDr3vYnaCSxKZ0P/HZ+L
6JEQTkeseTaFFxU2XbKZhTv4BW9/I9Hg/m8ycooZ/91GR3qv7Z3IUMXX3P72WAvE
0FsK/sjm/9oO0WIPb2S00g7HdW2PfL+a7SP7DK7SdqaC293ouNmHxpgU0HhM4Goy
gblU4dlLPMSEnrus2EleMkMDHzPsRF3eBACS9ZTrJuReXwJUmLT54T5a93JbJU4O
C2SQ23lwVX6MaUguei8/nTInpFxqN2WGnxWw6AKLi5NtsL4ik82bS5fGFp0RyGY4
f9J9qEViFnCVjPq1cJLvu4lWhpcmxwYDtL0XaeiXg0MOjI/Lib1xMS7oAv/VwSyr
ye4gXXZ/NF7hpsRwo5EojJgtOu7ymjUJezAdtT3d/TVIEMOfYZuh3NbVt9dmIerh
cN/tCqn0fDlC4Cl5tPrIgecJNxEK+KdrifR8BndXfgQcF5ZrzYiN/uc2Ap0+TFfJ
NmuE4rYUcHwxP4OJFJqgncNRboUHO01ya3ailQxZO2yKPLZEntAptJILizBNkV6d
Py8/Vkvqw5NNM6spSQRWA72FqjhyBm/sqYiTB9C4a2d9igeknqIpogUsNSCKItHr
TrTeNHjcI1DyswnOlsY9Na8KLNNR653416xW+S78Y3QqNsIxotkqRSlnhgYviWX/
+P7/tJIOP1EniTH0pfND/dvyHfPARp3m5rjXAZ0q/c2s5SeLS31YnbKTG5laZyTn
BNMrYX+I1h72SqEm7xUo2zCy/hO0o5eVuT6l4j86v+fo3GRb37Rwi89qji5CzGC2
g2z3B6VdkgT+Qh92yba6BUdUXE3a1NNADpLkl6R2G9mL1DBe1FGUk1/YyUSHrqyy
245iodfeGWXaYI1OQaPaX4jGZGNE/juOQsv+/ag52q4U5jNF+MpMi+LO/n25RQq/
95JebuomEyLWHu6Zitpk9qR1VcoZDxySpZtF9uEC9BG6BwMrtrNkG2J0XiCnmc8d
mgjTIQvReBYyBlVAEr8HOWNYPx1/Sj/8hv2qhANXgCAC9dLZWQem6uqgDNRYs6DX
taFKZt6dpxWnusMOxYCdqaOajOSMnfa5mqLK28JAAjMLP6grp4Fa9hGfngcSDUSJ
Y7QVFitOwXvaJAkqbOcspqosS477a/5+1JVJ6lDalNGET2pSAFv1KT5lE4Qi/Jgi
MGoDw08bPI4erB1HrIc8s/om6FIxd/XLBSCA487B1CwarZunRlsk3a5TI6UtBjG1
oStZSB+3sDpqwWbiuTJWjr7zkeEicl7FVGwbNJyheNWlP0XE68vAEnokqz9MRGXR
KjeF7nJmNuhoO+WeQ1xm1RaDBZGtcK5r9GnU9EJGEliS9yAJjRoDtclFRUcjFtUa
VT1/i0l36XYymOFCam8aeRa9eo/WFdeZjuCEQHOCVp4C7ZACg27lVDNu/PI4nt6X
+aRXHOGz6NKjqlcytsUCenzXPOyQqXAdhsOOgWuQwsg4Ce44/rF1uRGqciWJYVKD
KJeNy6bM6n/HY6I3gdOGOShBblokoKpX1IC6a8RWB7CzELyfzTz1sWLWgZT2zDQ8
412E1wK6+cabztRwnFAqsXZ8dngMvQpisVPzZh9FmHZ15CEbi5BvLLqRS7j0UETV
cxpuXmBit0xdsgHyjS6O/J0HDO3pV9draAUpftAk32KOyAjtRDfAkkgfQDgDQLDX
PvO0qwFTJIbghwgLZC5TuRBtizmJkTIhM1ffq6B5W+VBdnwllcjxHI2wyP1naAe2
FzbYqHutjlZ5+0n7LccjK5vB/75zJrrPf74tjNH7MGD9oJbxw0X/syA64UZ0cmzT
ZMRLxFaGzlV7ZRvnzYGBG5yeOUQlWTqKQpOO8XXx4i9Hi07z+PqJwEnCdQdPJB7w
u0Vd509vOA9tsKGJxhZld++LPPfmNQPFjWkioAxJUQzmVciyyiPdE8PpFI6y8QAa
PQ3z/ocxK1Ehx+ltbDqDa/lueNEt0myEc/TAsi2xqjhGtKJyGJ8z3bJSlF1wLYvG
grXE2sTvPm9M9gr5MK5MCZHkjHlqs3amMhu1lEKSp+sYcyGQ0f5GZVlvRG+81/zY
059vaprISBTouskFtrmTMnLhIpg0EOnRaBo8AFW2JPik98zT93ccI9uwjsWBOYHZ
pYhWhoTT4vEFMTqby68yTqazY9YBMRe68XyZas1GDhxXmW+NtMt9zk7nmjkeSJ6F
gtfUQq2td/ozClJ7Vv6a2clbeyr1OaGeIWC2ZJGNUfTJ5fveQEl0YdlugVhvwdSB
7DBUYrS3JmbZlYbVVCZAXEd1xmUo8xYlRaSXI6DYIqMR/1qjaWa3ItHbXP8y28aR
dnxPCDhhIacUqiwUko94xuvb9BXhULc2cHAJWg7y8Jm3SfjTDHSli5NwaFIZajj3
sGWBhjKNE+rHvTI4O3Au1uYodWG0/SN/3qOcqDk6Ukt+JepZDh26RiK4cFu/q47O
JvuvYi57P2o1RbpS6jyxUA==
`protect END_PROTECTED
