`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ql9nNWbG0ohVi/gniLaHNPF4db26Z/c2ip5pc9Jg1I/H3CeqtC2Q4ohqSLk2CYDN
qG/cNWH4gKzd1deUjvGDG713UbPgpOwy6eIj+XT6iNZoexvulkeQNkAVio855ES+
63BepF/VPCnsAyCpJ2of+Sm9y46OfgBYCYiP0C09/gQOlryQZUBd5AHgNv4AAUQe
xN93AxWMC7pZvR60JXeijHTKTIePt50M2Nuo8eDQbLYncxPo11eO7hsSAglH0wqX
uwwwmCneuo/i71RfeICRbNDR8GpBvW6iywbaXgiN2QKRX6Rl8e5bxWcaZeEFF+H5
UIhoPSZ0FIz3yBJpTZRYbTAAy3fbOd8m0lz2sLC7LtU3jQxZe8CmC7XdKDGCn6uH
0KkKLvxq/KGgfsLvJQa+kz7Lx4Ba9pYyh/8ll0I5zlWaJehcrp6bFxM8HjWjzZw0
cxzcQKzCgWgeG8dK2BxIbQRZNzhb6hOY2m2SmbyPXS/ut1K4zO1we4eKAeJrq1SN
EGWNwOPlfsQHEXm+R6DAw9woSGS3TN+9wEtzJPutj9tuMXaA0V8TmbZC9Lfo4xcE
b43KeTZhhPwLjOunVbJ/w5Mv4Uq9moxva6B0vza4SL+Q7rKT8jGqwyK4rGAB4TN+
d83si56BILbRgfpyUEEc48yjDbio3uOFKGCEryL65fGmjQwnME0Au1P9DtLJheXt
Hu+h2Re+bMeEgvHG1Zo5o3sb6ttnUdH65capLc3zrPBi5CUauPBeNzxx3GFg8PdF
4FSmSwVyrzdHop5lZ6iBP1Vhto3MrLP2TPfDnbAqzMmM7TMIZhtdoVvanL1c2lXi
IutGhJ9/+l7iK4FXWBPQLLi+NJ6NmveyFkGQGCTTTVQLpvnR72RQvM1hv3T3Ff4i
7jgycm375h6OlYOG0tZIPtXGF2wy9G8/tLbcE3Ga8W/gHEfhKORY5fMo8OQ0KMiR
FCtDOjPPUu3uTpIwtVWKqmnYeDcq2k2/fOwKwjlCSZ8hd6IGLgv6ge+7lAdcoLxI
3KhauF7xRHC/F8jV6mbe8/iJDPiXQcVy2ON0RT0azZ2YuONm6HJQQyW8N+wieeir
2JMY0PbIH+hurKcZ6uZ9Z9FT/+uCXZKQCi2Q62KaPMQ1zVBY7KpEnN7WXDo4Kt8M
3TyQfhKaRv/wB/ul4AUgsBxQ2ejvzBJjwrbxS9rzXr2/3WschNxOQzO9hhKZa9EV
f76n+UFi+3Ib4sj/SNFryzb0gOneIBJvdwD2dmBTAHN9KOX9Njs5IUC8D9cx0WfZ
X/RS8s+wAKZ7RtO+1on/O2dNbVB8Z8TL/8hV6P+pp3Me9qY8a989G9pioeLlgP7e
JRkzs6US8VpX5fX+AzAFCMCqqLx+SEXGOwNcjCz9oIOYJsywvrKH0LqLdEBDQxVY
hwpCNfGl2EIfJymAR8TjDG7RVG+isjqc9SEgwKs1vy2730OELW5gz/i5RgQQ1RUX
VyOaWE4+4MwQ71yOCt5yoaY3+SAMkD9s9VapDE7Q52DpqQowof4QhrldazcneJan
IG4BtR5qB7gamTcYC7SsGPXCszsVShisp/GUnvhA+jOcgy0UKuS0/xTmEGxNgm1u
dlv4gfnpnOj0p1i6Fxkbw0lecTphGeaZRuxhDX/Ezl3/TvZJ+aodJuH3lM7WDo5k
xnxhXOmFA+D4GhZ4s1pvWpzjAboa0yMCu52hmQVoDqJQJQ9TelmP6kvlkw99TBbl
aHXerLdjb9H5Jc1GfI5ebQzcmURd2iIeMX/Q7Xdea5HYsfulTD0yjIrdwzbi9/Jj
b2haz9YBpbspUq1XupMPAoBHn2QGGPGntrNHa7KwPE5okFG8F10Y57hgULG3N+Jf
bZpW2vMR6XkpyT7tWouFuQ==
`protect END_PROTECTED
