`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a67r8ItlcKn+ZMlptSBDOLe0zbqjxv88dZF4l4arqIiBVjVZBwiYchDJOpPeZDxW
mKqNEWhu9nagbsKvLsfi9Jabi3G70S3yQZtH5wzUmQh1AJC0nYPVvhz75guu4dp8
6auhPUh4Iw67mxeWlsieO9QC/EKgspwGqEwnuFx0zXE4z8vDhsQFAJy9Goj+2fz5
NE1nEEVMV8eus4nhhwUgXuo/f8TCHYBJjJl8yNGjwmz1XLIbYDABEv/r1qIzghol
ad+nXwSnsfM5XS22B+zbs6MXCn2jmW1kLorNctNnpglH3EXJ55y2ZgONJa5xxUAU
eScmH93Qn4jXrd7Aw521SQIBX9q3jvqHCh88/ARGcb6tkDpJus6qnwQoHZWwc03q
ACBcGfWe0oyotEb9+hAjqm4+7MXzYpFrUtzTIR0TRW2iVn02ukSsFDARozFFZCP6
Ka1umcoNDN4N3i7xWGijNQ==
`protect END_PROTECTED
