`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
le4dX2MH3x+inkvOvhbk6g4sZUf0PLaPfyFkXPTojhnYAxVcEMw5hqqvihJzukxP
ZhbFCvvh+Hh/2Vz7B+vlnDgpF3tUdYMzIlDRnyON/PfHVVecXBwciB81hDrqEwSv
/DqKQJKUS4jXEjmTf9/DLMb83SI8UmbI85edd4KUNgFfGpXxi6+E5wxRr1X2q8aR
nD/4TmeR2iBiQ+Zt9dZfl3bLnz45VCSmWnoj1TU/Z0FQm5D9J+7Yd3m0OVRFFE/V
UAo2Xh3GqsNjAfzXcXEihcU8FRomuPZ79SWhT3c+dGkT39vY13ew7GvbV5SyR38m
Uh4yOvx7xBTwBu/Nnh5hT61FCM9njnqZWSzLhI1JSqAwGMPNnP7EMQiBk0sRHlnf
B7rzxWlEpOSIIPTC26Z2nUZbDMAiaVvByfP1xXImXOPZFRywyTnvD3LPzk2XzER+
6xv5Z773MjM0+Ri+XPPzhdMcfSftNTOC90kbrrxlQjTzlgJLp6JE2Ag82KA9TJO3
cAq52vPJWISW+LTIUJYXdt6RetG9Hzw0zARg6s65FCZGaYrTOefhfGt0VPVqTt4s
f5fH0jrAdpMPqSKASZGk1jcHMCJ6HOXDW2hxYHrVG9ZL9r5pfdA7/t5PI2i4Y+Au
qYcnQd4HSNREPdICEEVAyFXfcRHFWLXpkWEm1wtBJO0meF3vdw3wFpK8izfTpOQw
d8fLMwaclnX54ao/xBfw8AphdFQt8JZTphoSMHnLzlz9UMu4RfkwB8JvKL0Zf2+D
ph6FGxcWrptPJd9FR4/BnvRNkh86kJjgaS5E4h1Ju4WuTq45XPwnJ7MlkQ3++Fuw
T7vRXWBVO17CaddCkvi88xQ+qfLhSlxhpgJJz/wYXOwHQ/F9JILh1vnb6chqJhIU
rXk3jFgQbijAVAKBIC9AXNM28DQfWVUqE/6IRhVcmtgk+BN+vopledbzZzHFLfzP
/sDdPLuVMnY34VX5LZVZC5dOdfq0wD80VKKiBJaOs35+JiBPFH2WghjCLomS8PKi
LB3ynSLhdOmaZa5FsX76H4EekCmwXivlrQWX1k2AuwWv6lI7cY6YWdHIljM//sDT
0LqiSPAi1ay+Xp5QoRY21L6r5F4aHKHelIAqU0hFBS9DKrH0idHpL73x0siNeZsh
D7Az164DAamNVm6ZErvMAKbYl+ZqK3VcZoEkeaS3BsIahpOMbQ3ndjp7r7uinVtA
aMc7nZOxzPPlbEl384IMjwBvGtXsVnFdlFCSqY3lAmYbFlg5N8Xol0Nkje/lJwnj
9VuU81gR19mDcaSyHJlrw8hqrnc5TJOILz3Y/jYh6CBMRoaXC2xDapHx1gIP/y9p
16qDf3WsDMCV37FqBhMWfBbLDTC0FbaL/Pm+Xa8Vd6ftIRAOdJCuW+wUPbZNAFOG
pEMUlOxAqHkNN87OWTXImdfg3/nwXdJ4tx9Va9B5adaSYkxrH4fvF5gomTXniXw5
LyogiAzeTzBJV63T6NIrmvY/mkZ13CCy3Sl04S26tBt2Mvteci1xGwTZAgTCVP/D
WFBnUKNMM0pWhFEQCCZ/FHZNhjvmKk8g/QCmyvUegYv2OdEqcBy2H9RxRI/pu+Tz
wrxYoLAXkoRKzfL8H/akGFF9GhtWRsEHNdXeBc5MWsH9TCL8We79dtWWpby49Rjw
Y7THwzDrNqOxSlqATg0KqSwBBkWuVgvml8PrkG+3GqW1ttNi4IphAACdFvDS9uPR
bchEo7OgPCoPt3f0wXET8JA5UziPrfJUG1WxnTjgXdzgtF6QaXFuJDyzWEfJzdeG
7yMxRpC0lCkevtfHT5Qu5j/vCIVRGde/o4K1rVyOUNhZwDk/uz7c0ebB0abjoLPM
k+7AwXtBfuLyNvQfcjXCtVjYMizW++UuYqLZjokb1Es3ttEhIAK6QCZrRH9cSlAx
kLQjRlIEIl/WyaJH3DoP7b726ZxrAa5gSuf1wgtHiGP6TGdZlV+surcyRFk8zrS/
mDiLuinYcsQkgijxy+51nRvCvZnzYGxI5sVyxklhODNrxXqAoCP0WoMl6AyxfMJu
0dxEpiqT/xIiRxHttkBnlN/8gu6P1Ei0xQZUM6a14QFlIxx0rHIxyfGQywGpOK80
6lDhLx2T4XOJlcK+c9VAhFihqlWsz4V/YxT3nUJg3vX5unau6swuYmQBwDHBFKzR
ChEQBpKR/bgOudeJk87K8hDstE57iFLmOQ0LjlEGp6IIuUO92Lvnx41N5/UYM8eq
vgiDitnmp+gkVds59PzweqHa6qRq2RCqoSWtg+IEN3ueSgFgBS6mUomAyNJ4xsls
cI63xZxipIgtjgrr/nfgohkC6/Q/n13hYfxV8Pw9iwGihPBkl2AFFcXxXp5xUwBu
npPZqA3xZLHhvYMSybOAS4qZIr+MWKyk5Lsm0YJB+v70SfkCiQ2mEpiq0bEZJG0H
FqNELCeC/L1YEgWSYNd+V88gwtytB2FWxYiT5omLPHTa6NCFh943smjMWrAOgH7q
JzTxIhecCEH1VqC05oM5guTXfk+dygd3i0sddqRJ+X7BbP2KcbjBoXKrWzAA7ocf
E+dD7klykLdRw/zxb1G2fvzG20cgId2faMp1VISieeRZo3cwsq5gR8DUlpjNkIrR
ggCFxu3y/O6BuzEGdRYjC557CmtZxLEFbj+Zz3+WGNSkyBJcQ1LUjsSIJ/FwC61O
h1WZ8QrlxjOQyRp488FQWB8YEa2+aBB+MyvfUEGav31xuigiffTVsFqClaTp8zxO
m2L855atOGJ5EObGHzFPhbZvAm5U337Kr35Nazr8f62t2ig+uBiGqLiYLIa0IgCf
CBqTT3LAUdJYX2qRIG8SrMJeGYcj7L8SXv3OJ3oOYLY65r8GS2ILSylcTyWM3fhl
ZdyRh5OoViFKNNcxyN1GRBgdMIMRzN6wOgoJ9B+95a5FUCNfvueM/4H5VT22MYI6
RX6w96vsVTb3/l5QMltNjH2Kpwlcb3xU9GwDasLwzhCnGtv9Qts3k/K3LdTIEtCJ
3tb9nind34LtM+kRwNKhxzfzcuUFyY5xHE3CsPRVdHbQv/XRItxwimFXZcTDu4cZ
CzwckGERPckL2Ayqg9IT5lqAr11M5L4ZGbHltvVyHW25D0DJVxOYfM0dTq/Vyz2O
FpoG18QXuCJxLrfhFmY+p2QFKVUak5DqxDfQvGShen78LN7FrT0K9cEGNwvOPKnx
vFWCE+nZboDdK0Zrp7Y/euDD1RUb3HEsPvYUg/FphCcFWhCd0RDLcAyG1dQXkBlv
68x1kqTjKX+MaOHR+0BsyCKFQmM+At9FsW2y1YmWFa/qdg0Cnng0jQ58raN/6pd/
0F+WO0tDVewgMSeNL+OUhR8DeZumeVTJOnnQ1sjTD5/RE5cWfWN5zqkxleJYiDR6
5uuhEIrOz8dR4IOhnwWVnxufYr8yEliZjq4aYYjZNN+tEe9jBUeynAL+aPtdgBiz
9rfFTJMCGWhZXkMspHtT9qlP9fHaouUsSOrEfO9DUrNrpiSFQTEHSycGuQ/LA8KJ
+SaWFeaJ4mO3boleX5mBxLRDm+YjkeglxqlETk+TBq2KKQntesIHh+KjjVEGiDQ4
VT8ubhsS6xQ6ASAU+YevGNokgbD6l7OUt6k2rQWWCkaskihXQpuPS8t45qndgOjn
yUQHJpTdt8pa5uiuroJEBmBFqwlAD3aP52NjRMDNCB6IYkT9x71AWpghiTweMThy
J4t4m0KDyahqnmDiRnHo9yKowAh6QlVT1U6AhhqChAXZ2eaZrKPJ+XOddECbrTqj
5/Fi6KHVV4VUMd1RPVuNLXNY61enbq9zbdL5d+Vtur+On+t9CU2V8FErEfSGUj04
IUH80ghjgct5z110szewop45wHRYgxdqWxE/kkVpw9VQdGebyc6lOVgOQTjjwvla
t9yI4XfuakeoeMs2yu/eJ3s7hDf5gFTscC/799+Af2zL716sBsmcWl/yEMSE/9/m
wVgXA6J01C51f/gfeVaa+2UqbZO2f02KvxBibJUeA/bdY4Fpzc83ImWSfCIVSneP
X5O9ngtSXOe77G7zPGcOFxH/fJrV0DaZniBk3x59BIW5I7pkwPHqEX3deG+nZYjC
PlRkA/zXhQs6wWfwcB4zrhOOYABMfdaSj7WADXSGKIC4kBu7j0uKnIXgR9PDUgqq
Fvpg5Vwkl/+PoEDeT+3KgvIXL3kwZC668P89s2OD53MUQ3f7SAEWGd8kt5vxQhza
Yqm7vD7eJorql4HySUqzDouvoiXPg+w1WtJA9vFOsN6Y320NaXJRMg8QLxfzZmVh
dMv7/yKJ3SRZqtZJI9ao7VkYoAe9HMwJ1xOM+fwFZ7FohEU44FRevYMU9JboFIUP
wR0wtFCjOrh3riF0/6dzNnqZVAGWiykR6sI7RNDO346y05WBwX2LWxRCyMTQWM7P
pRXM8Zih69TbS5YK5dXzEsDPHzugoUBAvgMG61gPY9DXJ0DdHUzpyoAyQOcO+xei
v+Jc1K+Sr5eTgxTv9EmyM16HEBSAqbWp3fwoWfVHjS7fFlrhyzHCBTG8bkpWbmky
vgeD/B8s3d7GYjdip9FC5eM5+SWixxRdlGg/TzBtvVa1p0NWPLsdcueTLBRIuhal
0GWa1hmulD9lnROQg5qqMxLyrK9Q4rObwUVhqGXqEso8e3aOj91hDVG5pfDNMUSk
/Z+xS1AAVNUK+KPY1JHMmdImNAQkwGS8Y5y9osWzW1g7OHtjb7xKGQPjHtNVik1X
277oYZGlY79JcklV2bHMuHoBhVeFYolmkNI5c+KGlDcid105HTrNn52NbSRtXRFp
osXmPQeR+MQJwU+c4PWvN980xVyAwFCb987TN+O6z+lHivdPKkqpCfgKsT+sHxxo
rNs57RNSqfpWNFvZ24K3eCBtDcLlSuTwdeADCi8zp1xiSYaRCPiCvw0YsdfrWR2j
DRqYMqEAK/Hl1GzQavIXavdWNxLsA5LM442WwdnoaTL9dQkbp7agIU2f9xPNQrde
qpelXEPc8GwnfOzC37NdTxS4r8wlwwyPBPH8dogRgKCIHjyd0TA/KPn4hIl4kyuc
jgVfLyL9U3HiJNYgqNEj7vKum0JGwMonED+drmWM5wuYAoXHbt5hCDGHn93TYB1N
PjyPa1jBc1FVW0ub+Dud3DiKEtRRGWrpWs8lq9JhR98tHX1dvdpgO1HtYR9OsJG+
sMnM1UFFlvFYFKaKQf7/CYA3mGhQXroQplYrfxPCTqJQjbxxgtvL0Ur5MC9qAkiS
QZSbZCl+nzi+3oN3gVbuRJ9dM1ngBTdwG2ZDwU+fGr41RqLCvgt5bWMmWm2bIm/0
dV7rsjstz7SQKPwqFKvX9xtgCmrkYpWmrdyeX6i+TdhFcgM3ZjX0l5GUbIU2+ngk
8r4SJIU2pdoxso1w2v/eict6qrlmWELD3f6Ts7gGd4uShfcA3BflV1cPuAcpR4CD
0IqHO0ysR73hH/pWZAsocISgqjUa53JaJlb4B7aNJCIkbYQJHzS0XHnb2D41VQ6b
FHNyXT2vOU127O9jnBWJbxAblr4oFtOcw7CJSNyRDhXKXttjaAAzASEnKNZAR86Y
LkU/UUdi44gWEWC8h0yNa2dHIlEy0EVLDqNbYJSPH8Mr4xUGiFUH4Ehv9mLOav2E
mmGL34ANpz/i+pS7Zp0GDpmfBC3lFeR3jTmSWJfib59V6a89l1gHFebm4e4tWJNI
udBLbbLZ8WCkDuEHj2veYWW/j3O7gN9QUwXye8QLeAE4Hc5uuMmWJCVOplDOjvBd
3XiZxnzuRn4lcJLaaEsxsYH/GVwqJiMPMRCGHLeORBcyFg0eMD6+jkXfCWRvZWex
wrjVd2TYHWrif1p+xzsozbocJbbGF15NpzkqVzxV+FCrty+AwkUPp/9jLeY8sHRZ
BV5q87zhDMQEEz/56gM0Kz0tKzGJWHbL90P70NEbCQnT+WAAbi73HLxdB3wdHLSZ
KDoiU5mOWLrrHlOVL7Itog/YKSF2uhTebqHHmYxw0ZlVE9rofxquw08ABVYNeOkJ
o5LtRy9GcD0UjiloA9DfIbAM6s+1h8QDKoN1MWYeQFGblfNtB8X29tA6YSrI/xfc
EqQg+AfaajdKbCGeKYcDeB9KYBE0QWKgLCZX39lQ3tkAJJg4hXLPYJ2YWdJyNn/H
w1l/yA2mp8XQyFo/L1VCwTs6/jNO5nGJT7Xpp7F566Gc2YHPRsvf1/YLLcv9jN6Q
vSRHhhx95/mwKsSSpZQ7UmsOryxRMUc3jNCOIE3S8rbzAzoGNPGwjMbeKy1qtobW
P49nqhpaNBkTj4HeThBm3aexmSs5jFfQiYPStu6brg+ZFwC4FUVml2caUpLZr1TC
FsG+NNiLioa9Y1KwD0fbW6k5J+AWp2Ar/bd2ifOwZqIgfTnnqwfU/m9VqrMAUk6p
wVWoHdY5sQicmkJifXtvILrVZw9pFRosKqybqBD4+0hswaUNpsFVYRnqXnqd1va4
rN+Ua0zoVoGvBqKo5LEREzOlAbxcBVmraCOsFQBqwDLHo2nIgS0cqt9EsTBmI4Q8
8jIwlOVqhFsCVKOPb9lNtGjT5VSNOf1oapLUU1NDm0zdDyg1LpZ4rFLWCXrALGTM
khhaItXn6sNaeEFgZlKCABblVCCcBMGOVFW9ZF0EEBtbUAMp1mERZgQ58BsVveT/
ykLzXuTUGx232ftF9RTHAU6qYHNw1IECe5CgBJ8Gvgv6mE9ufSgpIeHIDyp0x7pX
58qfOHRExq6jccgiyWhhODOkFIqBpXQFVsrUj9ZBauBR8w5+mM6FKpXMd9kWo5uG
zI6FYH5mCtOJIVlntvBC71QqOS09SaAAMf+9s9v0V3ulqSJCKF/HNKVcdks/1+lD
6h4jM3hWKaG0sv0JMLq9CojraYNuSlsrPRCgeCV6WjZk6T+jAmOwZw3ebdq4FLm1
Lqe8EIw+hJ7tBuNQdtLN4kvjxtDAUMwiaFSpPASQ0YMhdmRQ8F1TR2iPme1GSlGJ
ufxt+93e0conVR9Cz9VnoHRyOuZqZIBTaPHuMtxpRfjVsW4EaKMeqKmS6+3QwsRn
fJkKED7nhaW1xuBq+XvL8rH08HomWLQHq9iHQ8oYQ+DPfBsVRZtlVWuWPQ3vEbeu
HzzKBSGGFKBLilmY6pYuD3Ev5m9X3X5wtZTHmUaiOHIGARPN4wXScpYMIAH64aQY
BdWVD3q/NITbY+9EJJIwzvB9OvPGRCH9O36NP3+YfDJwxA9RMwpxZKEWKM5chEqI
O/y5yoFdHSj9/HlydryLWNbHSb65QhnpABZJXjq3tup5NPKcdIRaNaLtpwEti00k
s54f0S9oe23FYbw8Cuwx5qTJVRy5oD/q5oIu3xGwodAepktpyjFkYRQBilmtcgXG
TNGfcfDJlo0l/cRmBbr09krjO+fGKXlPcMn7E6pRWajDTFDBu3FnImKo4N9AIEzp
5Ib0MCv+qwzcEZRVXPrTOgK07tZBooUHJ2oYvWEEdt5KCmh2znsrejDebPQGaYdf
RWOwfmX1gh7y96fE6GmTv3RlYWAk3U4k/DNUfR4GdgFcEd5h7NMiMDKJs12YX+cB
dTK1krAaZj0g/EhOe7uAY9ujrP53NdBKfEmdZ1fsXipBabmsh7trGaFeP/odkIea
HmZLnH0FGASGvphBOAKyEk1dLGMR8Ujma8PvgRuX5mBiJwhwaQ0TBdpW8cjHCGPp
bkoZepcbna0ybdnbavECschs06hgaDm9iUZuih//+usdiWejyCOndIKW9bQx2CR8
E7YMK0k0ghbYqCIUj6Ud5B0siIsOjU0+Ou3ZLPomX7JMCeH1jU618C1GqPi3MAdp
i3FsLZVua6/V4sQfmheVxhr8SwoRpDOht9sXcFadoLhGcdgI+Z/oUjEApxl7bRaQ
cq2VQhLmxS1p7l7rStmp9rDdUKMhwtLHFTzUXBeqOXOKvKnIegxNR5NEvv4JlWIE
Kwzb7CNHvTpC6iayLjnUEIm79wzObR4PNFHnm1kywojQYHhhiBqJNEqy7Sx6g1ix
yzzvAgDIIUHqyBik1tHToddwXOzurBuFwWKLltMSchtFkphuIBSKkEUxxjVLB9HQ
TOR8qFnGmvqZRu5s6grgw5yjK6EhaqBTSErO9Gu1Y8akZFYvIS0U91SgA/rzQM8E
fjMQjAkdWgiq3YWYyKAXf1HmKNHA+KVl+bKeaR/RHyw0zJPEPYylracIvC5wzf0O
37mV/sVrTQ1QU2MGJ8c3uRVx124yXDQEQJq7Ucu66WBgpEceBn+LIMdy4JSIjhxo
zWhQpAVgAfo6DcjIKnLUEpW0IXLWqgJblHAUaBLBfMcQPpu8fKgaq66aTtNPME2D
2Y+lPuvyPAJDyg6QznPSaBhZEZXoauI5pGSmXWKuXS/UM0WkrSrO4MnIO/p5pocx
EYbMDKHnGQssTLC3VfnstFeqUTbtsMkXA9YMJgsDE0dM4lN6acDgqiAJe7/i7aJ1
tBUd87+LE4bG/sMXj1SABmFxBcuAslgTqsD281NhK3eUKuEIQvZIueJwHg8b3Zb9
tgyYwwj61ztrVIootzjTV9A21kMKhQ+2rQd0WTMDj7QbwSgAJ2h4OEAjOCh2f9sk
kTv06l9fT++XDDIKH99AcLbN/7/WGp0m+ANO7kQQjPIbzfh5AjMv6JL+1daSS6b5
gFnYETqOxVbAvtRR3kz/qAZZjDQU49kQWePOqg9ducHReDLoHYY1QplFe46mpgsV
TWPpn7CGuiXHn0lq+xe7Z8Xo2F+dMOQDHOK6xr+h174YLK18PI4qWKfZdnTpSrj4
GaJ6i7OiENWhajDuy6/w54ea2IyBGWIZlI0p9MjylxDpQ2sztOpf/FNRnhxIZUHW
kLqT6oqLfjnnorMIeKnq8FZYfAGZImhRZHrXyx0OIPmHiiAP04nZh+vD9fucBx5H
5Hgt6xk5rkU3QcSGxgS16r7TBJJv18JgsjMkMGstnUyVqPkOi/UNplkFTkH9ccaN
Kafz0tcu7yvF7IDL6kQU4UkE923QAaBbFAkK4zAFI8lU2fv3hgjbk1adWeyuoUh1
xMNGCl8nY9Yq2bfW+YftqxWsfVFClJ4PQYx4tMpCsoT5N8y/KI0qHXFuUlNNu33M
syiO+8MeZujAJLiigS+NeqSlm2jcn6upWSnuKE8tfvl8OBg45qY7bXZFxJbltQFP
JI+JQoHrG3tEV8rJQ8hs1BnAuzn9lUwDvckhtLtNkICIVAVP/jSk/ykEpOT9GkhY
hm/TzGRt9TXH9Kado+xJkcNj8/Q5QtdeOZNSk3emtVgFNrUfGvBYYPGyaj7JO6nQ
CJvKC8v4tN45YEYJFx/yEL9M+4RgCsyA2p39JpUHzMP0/dsRd+wFIXobdJt9EhfJ
iKW1OkxzpaT5hQ9ShBJjrd2KHxzsuFZL1aa55QPS5FucTpRZ3eHpsMQyPEwxbwUg
COhXuEPDv9T9SxE7uiF8MOsCJCkiX5+6v57wZ86dqAKe1OH6G1dIP6Z91VbEj5vh
MI96I2+Ytz/YuoCA68an5TlcPOMZUhpiOLNIu52+VhS2kdlt92W550zns2+JaTDV
azXYHVhebAvCsm3MR2VNmrsoEaaUp4IrTVWijf3eArT30LxHDo0lifZj/DLdOIMk
KMQXzIFTctBvhfCLkoFq3TehX8tLzK9Ny/qOLd89so+hKCX6dyVftusAWTPW/XDp
MrhFiskENxc/fF0Sj/tfLvW1KteZtzR67591fEpQ/XyvUc+Kd/F+kSQMpoZzgjLz
QXLmLgG/GWDCo9m4So6tIDvTkLFY72B79dz3I0kafJu1QR+v9UOP0JSHPXvCzq/b
S+q2ZrGicE7z0umfSYRzmVtRDBaxu8T1vOEf+SySdMT635IkHTE0wFB6kDs9NqXi
gvJGT0GwFUHG5MrR+SJ6FELRaIE9V24sh/fMlH9xHzO6/5QX0Vt1czKH8Wh0S40k
3Z+wdfX7HFaCgPuPjSr5lklYx94+J47fpsg6dTaiqU47r8XvcvP8o81kV9Zsfv17
HaS/loRAzc2nZCqHbzZtANm1rwP7hgk1zDCHCSccVNGe0eWtDqYF5A5e3/zcLbqn
wHMDAVl4Hhx0fPfFxIDPEFziPw28coiddULGuD0c8FTDxxDVN0OCwFCf8Zr8h3LZ
nv20w4VpEP/bCBzs9EWCWKB0CET39NScvNwkVaDnNI4ttHblCwpz6QApTR2N345N
gj3Ei2cDAuXXJYITMpjqt01I/GxnKcXwO+cn5kWGG0tGBUB3f+IxunLXwplTDsuV
0/ByQNaoJV1MCCN/WzfnEW8uxqBoChax95t9G+3XvASb/eRRx4Ytfip6+fDcO2tM
yhot8zu1Eu20ICLi5svYYQgskf0hLUdQx+R678WuIRz8xZGM1ySRnPH6YUeQLJNY
CpkIjNoJ1ln37GtTsWIijnYBA+SILN84StZZkvcEzMRyAIxWK3xBJIqZLXxcAUP6
T8Iwk8xJIcqXWzsd3v7k/oEl1ZGjJ2rPgvKUQEFZC5ixhO5UHAkBWYssu/mLSGm5
M4AQXCFVvVEBH5XpY5XXJR2BWVpzBgQM0UDIh7Oz1R6NhcjLLL4ejOkZersgtLGs
5VN1sJ1sgH2EG+yOGrB1V7mm7mcfkGPa/Z4z74DuZ1IxaxikTectX0P9/iPZxa1v
jdkYeIvWZ3MsCClI7EltRxTU9XAMILsVnpYi4ejP6at7lXnAmWy1JEBQqw2vZRZL
C/fZBFuNXiXfgXqeqD7Wu2VotGMWJGMruxerym7wWWg/QPcc2zOVdbmqG0a/xjlw
sI9meEfkTcu+8Iz8SrDYO3UGmimRZAmZNy9FLemPslwGfBpk9mWpYoIJn8zJqC3Z
Epo0jZavAifqgvKGcRosbPXxuhRgeo8YsAcFWd5s+d+Een2JT/tbr+yBvGtdF7k1
loyHHFWrVqiQn1OPuwA39ZcXQsmUYDUcrVIg7DlGQvCMlY4SUJvQ0hKPnweJxfjn
/pMczBh4yytv7v8gZmphwIcBhgFFWPjJQaOTHBEpG0n9pPVkpDZ1Afywk+Zm5hAd
0SQyv1WdcXgjjC2/Lw4IsP5I4umEugE2+qMCic9zLinrorshKawVWnXFSnk3cbeJ
3Ejpg9a6ejW4k5/ZeOeTxHgnEJdILu3DYYXX4h+OsoFzUkCUayrBRbieOGydw+gr
5VB24sbVJSVkHP+PNsy1z7Dc+igFRidhflzJ0iEgvM+8rKry+fiZUgtxAJCxA0dg
ujRU68Wq4IBwOfl1KaGiS6dr7zuDGPtgdwdBT/r5yhU6qDSh7Mdl36VblhGlk7vQ
QPXi4jVO7+Ni5m33l4nfQYJWxj/PNMxVYQRLbOJDZVmQZenvTluqryvHBD0xOS/q
ziwMlwE8+WbFFLOL4FB56MUelNUGZtRoJFDJfJzGttz5YmSb+oWyMZCzRVe53FPb
igzVM8nJ4QrDB6csVxQ2ADXFSOHlazjwltDQKLUP7opQn9Zbuxx5+kbXricGjK09
JTK/fRzUi2eGeZ2QtlIm1NG9EjE1TshfO5bIWCThJyAJzeV3rBwZoeS9EKZHETvW
hyZ8mKadgm4DzLJe51bTvDfu8k4rLDxplrHll4QvSpa5y7NtYVTnIhFt3HI+GbOV
arsSkoZnKwRypTK9X+5PqW9GH92zGwgF/4OSaJo2l1NrKWfaN0hbyYf7/3TTLPXY
xzYyrpSc/Y/TQrw6m2g9WcVKA8HI9QJYedgad3b9J0VDUISYoEBbZpxXR1rBG3DZ
bNR735kNXP0+UC6JgsCArmvTKbANBzpfUEyhUwj7ELfAyhL3668CE7zvQsVU9WqZ
QtUyOrB8klLgT6N6rgWfqoIIJa4DohYruEr7XfYYQ+ulPmrJN6VkuMBxQAC2Vm8q
IWwuaXokfY1mpx7UswzffsEPM8eG2v8VbYo1rAfm9eYObq0kmVkyysovRfXJp45s
d/RmlLGu285jIEeexlt09unt4ZoUx2QiGr+iaiccW7tWxHZhP9gZp4ZHcA6bwYkI
GLMEIIlDx523e5J+FiS2WNxQ9XbLHTPKzUQNXLWxEDAVNMmx/o0aadcJ5oexU5+S
i+3zI5Mw4Ap3OuR9DBk2AETmevYVf9b2hZa226CP4VHtNMxvOJ+eynku7vgkoCVP
S8h1pAVchBhyVTmzjg2kr4pkLwga5RRZ4jnsdF9EK2NiUddItmAwr37l+w0EOlfD
xp1wKoTkm3bFD7oRkUALpjSHpZLlcp4fOxqI6SEelInlueCy6ob3KZvihBr3zVM3
wAdff95mIGMuZVuMSbwlo97zdz+7fGwgXIJmJN3KK4U+Nt/3jZFXNSbBMyQL/aWl
uQYbHBTcfMJ9abDX2LgeJcp0wmM0lomC5/es22Ce7xETFg2OJpKQ+vU/M2KwbpKV
SGMxHPn/E0pkR+y/LoMKX9vaSbeM86H4YQxgcM8PXy9VlQ6w7i16wNu86D4MHHAj
IznLn0gVcS9wxN3wvik3wEhUq+7sNF1w7lvs7tr5uh4X07gre4Zs++K8i51QmCzU
FCZfDhqH2UWvu/yuHhT3WO/DE7nc4U8iYNKuJ/eejF3d6JhNTbqDDxZEjgO4yywS
KnTrJsMA5QVU9gizlqp9aoyfxL0ZRdtFPPakLM8N0x9wIReEZmOzJ7c3Jd3H8Ezf
1WoFGAG556gLYry49ASOHmeiPK8vjWmGxALf6SIBESFgoZ8MC+DfWOOnTASUh0Hm
hicpUDfKwo8W5s6RTMqxRCaioPl2koxkfTdoHSEqigabCiXEqRmT30lIneGBY7T5
3VtHUWSAACwmUZJSvLvC/a3tq8lJlMenh6onL2sSA7ybnlZS4S0g4BZhZzkuwQHL
4R7Otw9WbC/JVczJKMS66o8DI3hbm3XIowBUKV4Xg9of/xSSA7cOm9e5DxGexo6A
aVo1iZqt6unMJvnlgpVJrHAjL9POqZH93tes8AjqRolCL25thl4IB4tsQ6TAeXda
0Lsc8/FDRepVJJ0PoqaWTYgdp+9cB8jFU/7T9wESDkzvEGS/86afoOVPa/Be/iPX
pWVWhh5qHDYwEdbDWVk809ivHTvHV2HuHZo3TKASy/wPMdgoqMA+KM7lCp3JQEec
7ERoM5ou7rtbSIlYKXTnAiQCDgVGsyNuW4sYfj+1UYSnaF1/RBTtu8mTogPDi9QQ
v2KiujsPJb6UV/bqvhY4CIQ0ygobvbOsUijlSAE6E34ZSLHYxi4x8JMzZc/sFHF1
n04vaeehj7UY9jKEtOQVVqkifv7y8S0nd7dhsiBqh34M8XDCJ8HwCRzEnu1Ljfpg
NXh1znJhoo03pj2Svklmauq6cBQWr4LZeJfJoZMXP+uAQzBzMfRkoQaGOxPaRX89
rC8ZvGiRj0hCv1LlcVDMNUmW8Qws6OUXbjHYKzu4fU00sgDNlfAVp4kdqvkTg54d
44f1vfWflXE/BERdW/atCWa5Ma8xaCkeXOIAIlnUVqbEEli/oQgbUT8z1DR5uv8i
4DaShrPaTarg1Dyg1aycioFSDJCj4SwO3mB8TEEzUJefB2kLIzc1gKp7T3uVtLkD
Ut2/1vuur/lV9eL5J68Y9wm+ouIB0K7NuDmiXEyTUNvZAUTbY6SUAIGzX2PqOAMw
QSIw50OC8lqSCIzdSlGYsmsHkK+H11IGNgdoyhpoPbMEROzbqxeZRq56mnDZSRul
mUIwAfIBW0aPqbrMKoqO8KzsfjDgXBtxd7ysx91Ar2H4a8fvmbwtEYduGVUnaaw6
uXjVNpEUEPQFUsaiMUxBDu9l47zUii6lhpNSJVuiRORhLPw1sUrird105ldPm1GN
L9buwSWzN76C+PcMU9yGNmv2926d3hehZFySqGpxOyyt/rKm5PKs1vVNr/MfL3W6
nKfKP33WC4jA2q9+dvOPpBe3PCi6kLOm96t7yS7xk5Wdrj+t0At0HyhKsHWQuu77
5D+lVMHjSgaw1tYkX5CWGO3WLns5gvhOxlOzL+dm7xjpMJLKyz7gYrJ/EwOdghDB
VhSaCEpAZvtqiiPnuLJmWjjBNnuOjnxQSCmRMFQSC8gSbNDw+UnemF5J35zRozsr
aBAwIP8/dqJe4OkOGuN5mCMrTjyjN4xroociMg3NIhjeyATXovP3F7wb/lcGTvSp
od1h4TqC84f4RwCJzu8o/GY/wlf1eDl5lQuiON34k8/MGEmFrCuxkQbYBNpm/8Pl
oI5/mifpXrlNuibxwrxyV+YhPAhyrJ5jFSkETcU/ojBizQ1LKA8IY8CddjSVcDRE
zK/3aU1sqP6UJpHXrc68dMV+W+3sTo1nA61dE04Oa0IbWxa8wVJb9c3RaIfHyq/l
f3/UbN0msYdKOVix6cwjJSBno9dwfDiK1064JxQsYJE8pymTKJW8M4rB3JbIO33D
TrE8PIc360O6OYc6Ut65TuXyh2tCGg15qnzC/imT803CUVDPO86Rx9ob0ctH7sqj
MsbV69Po+wT6w/nfqUytA+B0h2TpzbxGO4rB3ZTO6iCBU6ZVEhBOQ49LBASXEmKe
dorBb9NMfvBKquBPu+SZ0aL6KbAH33t20c1GMYxiFO+d8h4iL6y5yWUGYnxYLbw0
Jk1p87Nh6uylt/DWWN6kPaddlPDVA0rjv4P6rQKzUbn6ncqfilKjelQWjBylqtwF
XmGtbgsEDP6V+kqdbNYKumGe+VxNlQvcjJFUu9H0OZAWEr1cMtbVNkM1MLZukSlu
hLMlubNsJJqGnfbdbHBHtJUAr7m3e8oeXtVTJORgP9RA3tWiY44WrU0J0oWE14zQ
T5IR09C2dOjwjfy2Klsjsc/yiYLBDLnTf+2zGX5hf+Jr3jbvFwhMcJjA8E5rfeo2
pLD2EYEobsgOEHgcyf9P3X+02wP8ox0W5gn6YFzLJcmeZ9cnsb265jZIzQrGh10r
wCJ1+zfpLum/yHsj/c5OWhb7oXyn5QOHFrPAejB4DsRHZpieZ+qLMI+f1oSgSMoQ
5H0FIqAzJkUqCNp/Ui6L4ft16U22DxAy11cm/TfxnYSGaKL4ycjtSzvatBj0Vv97
KEa3+5r1zYTYrggPz/Xp39HvR9T73r4P3ZzpZ58qyz2BUKFq+R8uQrGYHMiVeHQx
XmmX1m/HcOD3uSh0DtW+IcnWJ+JqOP5HiS0m1xJrrriIvNaqN7PJri/deF/F/yrU
qgeclZrep2xGOEt7w53jZd5EaA1dQEXyXloNChGn5Iv6okZX3hZmJ5suOqfFVlYr
169gkFHxUq2h9HRUEJm8k0ZfsE0c55vv2SyxmM+D39g+DJH9KJcXVn1QpAFoKx1H
0MaePU+MqZ5MDQuWxz9+1Ets0mZ3vxOT896fgtj7VEcT5YiGqslG6v4PD/jgAgpT
uXI1EIwdurvEvS4lyAOD48f57gxlLQQIrtzCKcI4/QV/9nS+F8dZKnlYYARhVz+E
qaWjp7ixUoGOGxx8Tt7nWzCfTnY/32VZ4sqN7qIcppzLNmImZttAIIkSaqO233en
mQ6FlMyXoiRyolNrjJKWFTHQYhe1VQszqJow8DB1bVVrdg83DaETUDcHRk7aT9n4
fYoeNfK5W2/HS6yhP1lDgK0al2MtxJoEFN6qmgY88B6pBe31x1gXXUstKuTydEdA
hFJoRhpABjP9NLs55OfOzlhcfo/B/z726x139GH5/isLT/dcdS0Y3PvyhdM/YQVr
C6xhAKXn4bbQciibb7baahnkVQwJjHpn70EI3gg432iOhOXcdsJLFTX0xZEwazBY
8y/KVpqvr35tW1I24WmCJxm9SzXsKTLJGNuFMT89+7CELKRyp873yuxP+ohGHlu0
XJea7USSLtS+BLuO4Pf+eil3Wx5kbwWS63R8qakcH4YkG8+q/N/uncbRKsR8oY4Z
/ldQSX4tLrpHzBnt0w6vikkH1fNx81zcErMkZ52cuaVmZFz+a+snAqvIctjwpjLH
ojPu6luv7Y74h2eM2mxH0sAQWeVoFPhRfzp5MEZZeazhsinvmqkATubLiTsCJgn8
Nz0G7l5vi33almFHlF5t1KOSB4AD5VD+m49UYRRm6m4PtzqEu2sTQjk2k3LyRgPs
EH0x8t+UrgXjeBG9V6WK26ZJxTv4iIppsug/oeEQOsG4Raz31OU4NnrCznQD+TUz
kHQP8cg5l2wOO5Xo+u4Pby+kG8oKi/APxCWnup86ZO5aJXhD/LQ1jHkOSq+0obWD
+8m+DXXh9erS7zM1nQ47kni7iQt4WErA5GlEBvnMmru/xTOVXOdtneWAmfIS8W/9
Aw0Ge6lji5xkBuCUeP8wZzBOClaYnXitKKkyhFcsYJDXR1uLgInNs1wufJ5SBmli
0vrncBT6SX/cNK6mxcEMS53zhJ492mnKpoJYAKYzUGTMZqm6qOtrGytU0/XxMJ4d
iamLQwFxRD93CTQtbVZXOUFu/pjGRiFso8PVOAbJp1zb50mSenUE8HlkGi/yOM2Z
cS4K3gUTp9RAgZ9MZ3Of+BhnPI7u0YMAt8+HWHrXdl5JGfwEllyx6TK9LlbV7gcf
tvyr0Ry0UTO+YRFjof8MvONqr8WTAi3pxMwcaxw78fOzWfJL22Pp4wOU/gv/paAA
5Aw6HviaY3xT5r4owwB0OefaWXmpQabp7IjL5l3iECWsSN5NUa+jbMHOzWS6jTAm
MR0PXXFyE2KfBoy9e9PPaFGNtlSRgqNP7214ZE69vfnt5oQUTtMywuhWxTIMK4tx
7dKhHHuBImYceSwcgNQdyvSCc7KxojbHljzenN4KoYYgcacWcWF+6Sp0yzuSL6AP
9F/n8ESPmb92DTWl8r4ReyNJS1VG93fEntKjuB7y+6oIZh8lBGh7tE1gELr87l5y
Wr2d8CKk63ZOJmjtp02PyQqTWcqaaQYmiPGBBEYMHmjNKLezy9ZxGVud0j8IqT7z
uXK9oQK95glQHEzfAu0jra/DDLZNY1SR9Umjj95W/Uf1cDOFNu9njcdwaypXOjE0
ZxrdfaO3uetrFpEhmr/TKeaNnLF+w+wt5BjHTNvRPfyncCxbH7B6A38xhAgIMuJj
zZFTtt9QoHQHFr/szKKj4MYCV/bVZUx2LAXTwZOHhtGDAJehYZNEqHKLuRIiybYQ
7sDEL2GfA25MqtrrupIo2L2YfgYHGgnWjaGTxVVeVMqkQbIhTxxxPmsEBA3mqttX
sW/dD3zZOd2LDTsgg9uko8Pb86EpGW9MIN6vw6or5BOZDhPsaYCCX7C/chX3JDdb
eK0Wveo5jHB22AM2HD/yD88j9KlvKw3TxvVTaDqOReQdVvnBXlFP1vaLgh0Toi8K
C9JhYn6RSZelQYtGOXTr4Ci+HhFY492xDGxLArP3t0i/5G7DJYlfjnelMmJaQKkW
M+ZaYXmn+RAxsIhg6h7GeOEAeyUWzyYgfwXu4ar4cs7N0OFiY5BfGhOf+cwJLtvG
aGPHwWcNtZX+Wyc7GNa29M65AMQ+04YVTC2rao9ZmPhIwTpg7Dwffjk5lU+JNn2e
ZfC1ylOhGlLupzXg3GQoYMPLIWMBJ+V5p/2kFtYMFMhHGyaEXUBDDdl4x4am6LEA
rx+kF+9GDmt59yf5Aj6p+sXeNzY2BHIjA6FnLNGWSg43xxyITqoxEgOuxphLvW4z
Sq6WFq/ZFdUeSH9sGwahuampakEzjYsZzwOjrzHlJqQP2wmQssJUru7N62HcW/M6
XYq+U2zyn/UcnZ9KaHhHzUr2mGKUP4TCyB4/5vM5piijP1uPK83FCuYeeWyUM9Cy
hlM4H/tjJIDvN/FrLLs6qAywtJ/pddf7Lx0tV3g7C65GZgezTr8TTbvQiLcbPR/o
b1/LsIeT3xqwpuzQSiMzqy2KiT1qlo9ArG+D8LnfNbGg5uGBekQ1OoBPhh6qYU1R
9/yqFPN5NEJx8hJkGrdrEY7+/wYAYiwDHAeZ1SxK1P2G2B99lf4timKefdBz6zoU
cZobBEiXv5o5iD3cgYSmVjmYC7f90/H1QrFYSMRnUGv/WlAFcoJBNXa1Ij9Uj+Hp
om83JvtfNNy05/u6l2uzvDV9w4sY1AOOSxLv6/3fnZtzylNzd35USEkIEdEAbBkH
Y1qnDzD6sllcMOzckbO2dLy9bn8pPlFYRutN6zgcLu+lG5aOylPtjZ4U13m4JF3X
P/c3Ntd4rhsWYVJ2VeBS5yGUQ/ddGg86n7aWaXQ/Ez3386bmss/5x0p5CG28GVjB
gXWkskuyzZWxF+m41eRlY3Yy4khGgPQ4l7ilVBpe3B/cd4IpzhspK/6y8xgdHJ6p
Dma86yXcNRUUYSxq3OrCBoGm0K8OGZFJKZGYVyB7xHuF0BRtEvQT49o+wLs3gK/1
/aogR4C2IPWC+XO/z1Z2SS4fQVsLai/OLu332L0bpeFyCTHUjMjxngefywiM7EKR
zlWbEFpRe0MA2wHbRwi0e3ZMEYY9LKeAS2kidwxNJrtsZ6TuZ7vm0+I5M2glDenI
AYSRa2inWOoL+wccfNe/dBckkTF0Wl/OPVjVrKhrd11Dti6VApzGDKgpUMSDiriv
WUqU8sXMLLw75dvv8gKK51eC1+HSrehqY2fWUV/QbWL/tH7Pive+4C/TtpDX/XH4
FG6OVEBGYaQ/XZeF8BMZD8iso3x6oTzOeZfrwngmn5q9VuQZ/JwxqeuoEbC39VCB
JzregN5JxX7/ABMPlx4IR4IryXrtIIOVixtK3rs0YuKdi8XUGuJe2Z3NTunqva/L
EsUTvjK7GcWtzw+9ywB7+R9KtuB5lN3GwcSVqt5h6MlAKvEkRQUHQ89r6XeW6JMw
STPBfCSkgiuvQVq9lNkprNL3EWGsR8MaORjSwR4Q3mbdf9OYRjRsKj4+pv6I0qZF
GPRqbbqNSFunJeNA6b5Nnei+8bW2zPFGwBLbar/CN5n5JJC9JzBv9OstQsoFLEtg
jIb/mKF7PTbmvtsfaGgJB6aXLwfH/U+8F1KtsuiXROSTw1dtv62GNVQNSpEE+1po
B+DWCp77yph2UnHice260k9/dAmm49rGAiI2jYWpWjSit/0JRpiby1lCPDO+GFrb
Dj3fpjsHpEttn1pdNn7rCUXy0UeaC3jHm8jrvaY9xUhsOQka8f3XFhUejJfp6bKY
t/MMrx7LGKMY5QIgY2KBi34XCgwS4vdVk0hbJmLJJPXCb79qhvbtW9b/RbB8ntp9
2y5ukcIKsS6IWEtKlq4Fe+bLlZ05D9qKcxAB9wdY3b2I2fk/pwX2s3IboIjDixBJ
APe87r2x292OQ/38wzWuR5d3x+p5CBARE9dvoUamHsUZIOsxPlHegLe34uQoEgOQ
Ooa95LAAtM2gOIJplx9gfJRG09hX0q4pwtgjCmSZIQ2JXyWJoMKjwhBRfO9QYCWF
+G0fQ1NmnIJDa1MIqI+8qaF1Ena6F6Qm/ji9dETlulr2005Zoz6JASFNSryR5ayr
ssa7Kr6op2MVKN2zkV7PM5ck0dK1nuDj0ZMkPSjDmG0feY+aWUYkMW44cvfjGsLm
Czm5VWgNQudzJhcg46id4DfbKeo+hNdibO/YOMoaFrsoKSytLE60XatFn/QAk4oz
rMc02JAslJouBBllw4RCeThtM5L+0nrdXVF8YOjyvVRSLPJKfzGvW5/A3S3FJe9s
MJ8TWZHgDa8hwps1C/FJ5s7t8048Re65xHFEng+gCXd86wBdSftOarA17uYsqx/g
gUrWWLbo4lQ3pBmWGCF+MqQTxA/YFiits/q6IdwiY0Cmpmt5V4pl/gnnUZWx0NuB
gFLzQ3usVNFH73r7pOnYYGQqWf4A44b5uZZndWgfWhHhNEqh87ZqzvjaRxWuyjHX
oEaKdaILYkAGKyTUBVSQQ36vIzQB8otHaA4L/XBNrjxCdWc0MWWVb4Szx9jI7nTG
mwYnRJIvJQgKtUDiNqyzvxxwn2HBEIQ4b5brMDywSrk9bZZU7qCINqkObCFx8AEc
P+gFtm6YmrJW6KCinxCYgD01YyJ+qcnA+7SQpf2x2k6RdK6zj9W2/YCpwD4wyHyp
Y6xh/UC4ZFGT6DEFulhN0Jt6/6QVk1XH/7+y4lyUAH146E2fYt32LMyAwYCWdzrY
UIUsLH0XMrBGr6CoYK3Z7ngeGDqrmTtqQP02X8zTQuzmu1mU//QV5iQrTzH9wi6U
D6itrgjez/EESe8vqbSEuJFlobx6N6owqbOh4mPcDlX4LSOFsBUpd4QvZO5nhdlS
KNMH+ttrG9Ewfs+KVGt8rO2tpYeMWvxQk0Qpy/9inekIjuG8CbFy/hoIEjGQB/zL
f9C0HF1cGJeWAHFsy0Rf+HzeOCSzlCCAcf7dxGPf6Baf8UKX4lkkOhy2Ojz3uBNo
nQW6kFRRX+OpgM99S7EehnD7GdmsNXfuNWliz0Q1llwewU6gw+NHlTgZL2V+uScq
+TfKXDXWwbgLrIUCfgu4atVJ2jQxovcliaUAYGC3Sc4b58qSVLOncwEZMgvqAyjP
UgRL1CoBrZuynFCNLj0GZg3WSZg1+c4F/L7GRIGIoCK3IU945GQK084u7nBIhYCD
qChnYSx0QzDXKSTksy9YQeI6d8AgqcExOgihnisTPXFGmroez6n+Ed0n1Go5Xcgo
BEqah4xeoNjhI4v90sl0STuSU3OHlipol2JzhV39VzxdaPeJ8Ls6YEBgrEmUMyqg
dNwHNPOb0QTwnxH1qLIABYDI2KPfgzR1bKpBrKH3TXiMEoAaStrQT86udTESP0U7
fi3+XF32jfRMv1+CIn6sTIZJkavfz0YKVMMpuHtppnU6gIProWtSJOl8GHbEYelb
m4IfbAXMBnf0oRDTXSoj9ibJGRHbYrdOgs8xeYvFjd7WcsSgmsbOgeM4gWm7e38R
WXKRQnhseJdKDVmTrWwgLdjJponw07kIMGaXXJerqsIRJ1xxRIFnH1laXgC0ao6b
5sFMcE06/I5GkA+B35hMLEGCwEgchtuLiYb/raLZ/hA9Ba3x5BzN4dOVrfpX4bj/
Mf8SJOAe+QDTJnPW/CqBrOPPnyqA4EwWxx4QaU/7xlEa8iYDqXOx278qemTT7Dt6
Duz+SCkdV1bECoynppQuIqlzgVSJeo9Wp9swItpP8TZBUuX94zxLL8pBKbxRZyrx
sD4kcrFOXHmYTSjj4rfx90lxAR4/VCQmFt8NWVfLpCpbUtyuWcMdZ0C509/EPSVH
QzTMMiYOiipmzA/07Aw9Z07Qi7SHqlqQnjPI/LZJ7XLZQrEyGwszVQH5f1KIhkI3
wfdMnVb2T3gbYcCOemUfD9at0JQR5zsas1+VYFVSnGiXfkZTbeu05H03o4OsysyX
reFIa+pASbyUl2zdubiBTmYi6N0jJTLBCV31Lgdkb7gj9gjqq4h9RdXfJ8PGiz3J
93nMgO4y3QJQe/WvERrI6Y1yZLRq6PxGJceSezfjT3m6yrDI+SQv1tbX2Ham3k6K
xrkI2zXZOlnfjQrKMj15ZGVj55BFFyuqvJoY2W1PGwiuqviz2w+Ld53wTzfM/8wG
FSVNTN1GkTxj6bA/V63Url7ks8OCiVh95Uz9jKuaed7M0blkIoIQ4ou8M+a2PJ5U
3JE3ppv0/DZ87tewaKiXTNPvznPy4t3MqZXSn51vc8ghmayVsuRGbI+C8EmWjWhS
u4Ldsid4yf8xQVlmh06Rso37U8KzQWBEXuG2YHD6G/OABbpaPGTkA3x/zQOZS9CX
MSyGh+emvMkATycqq7gD9rtJpsZOiOp3/CjdeBTmzUV0QGTZkCNSUJkk5YLWPziq
z7EuNzumAm8mUNv6xnT7/k7lATo0RZNJS8iqjZBXUxFFNbWVX1iXnGnL9jJkQnGa
h/LITbNvrmuu8CUkMDIxn7n3iBp9UAUzS4ZWS3AIp1zNgvI6lHwZECg6NJcrrh3/
lGjEUbmJ4MpqGMzcXMQu/N5mDZ3/kUyqXVb7CryZpcpJ8IzCOQNlVsU8igYykTNC
UlQ7ZJunZ6u4VVxTpKag96hdxWW7VMA2yaeoLMrggqt4EKWy207vkeU9j5J4yhqH
kR2B5wwox3vIJM6798sKvuhTB/9bDwNuDOILWpQa1bk/CUFWiXhEZ1xhXWMbF95A
JWI+RcC71WmjgSXVXX6/KHmUoQYjab56hJkRUYYBiv/yh8E+WkkYNkli1S+svnAB
EDqQggJkomPvdIWYvDjpjgOsm2mwIexCEIEIubMeWZUQB4GLRD2I+Ewy8kHIfOhl
QR1IOssRDYQuYHmGlBMsKSJhSD9mMJQFsc+DR2x92w2WMIkgOr6Hwyx7OwI3vrDC
BocKiHn+Ic4QQKlF4JVXxWC8ZPcS37vatSFplJWrNNb/100+iWYq9GiQH+396H/V
aw3pK8ro5dxLG2YWOMMXWZdSiaXrIqvsJNe3Gx75a7EFixJ5cpvNgHH3QneALJIO
VvAg4lcYM4reL++ZcPvteM4Ga+i0r/d102bf+DXm9YxUYoNK+jCdTfYzlsLhkPPF
IeZVs88sO/qi2sJ1I9Eufmuw7nAgyVA0ZXIdkjlYhg4Qspad1sv1sPZHJYMBc8Dv
/BVrecvApKMJDBoxxALMid2irO/etkINQTYUvtsm7MoS+MVd0Zo+e5FqgOHDAcN0
261O9KlJrv3p/INbFtvwFmYWKGpeSK8uNfPimKLRfZ6CXsdG0W8aM61OoaufRL3j
BYbkw0Qcm96HlB0UXXDe/5tXPsAVeSG0iLIwSUfsAG3qfGRCVcPpDl74FZ+cmcIC
RNRhuMPKnRQeksE2+gVOcxi2oj2Jhgiwt5AedI6lDVCKpqziGKDq1rKoaor48rDt
BPpUIGK6TIGx+uA3grq3Lkexv5RbpnJB5QjLqPKRYtKHthTk58Rvv0Enhcd9DPs2
UffQ/Q83m0Ak2ZuzRDx3yh4c8ALPiJ0H4BJMdOvz1QC3jxm3qOwDwPLbrKpB8XhI
UJOZiqE02qKN+aa4xNiZFO5oPyJRJZy4JiX1teH+7UPSdqIuh4yoHVlrEZ+Iu5P7
djI21lzmmz+rurGCuEa6oWzs7GNAfzqsfF0Xzngt1yRzozzFrmAtt2GdStvFVwZs
Yu0+R7pKsOGKhajxHs+WC7J2FL49MI6ftd5NOqk8rRw4iwFk8JahaC93OsZVbNbx
PH1H/fYyUbpnbTRe16R7wIX4hwDsaxjbFSPFnHZxQOT2kBLwCFURCeR6VImBVZqk
D9iIZhiyzs/tyv+5KgCVAu7WauMOCK85Ur8HV7mF/3MwHnp9DKzo+3qCklHyIhEU
QQF2heRPV+VUa9RYE16EyeyGYnXzrl0SdXERn4MMJJgnHrsKrh7xpyH2O3wZjPO7
d9wiDFud/vu6odcpSo/2n57WNnNXNEoixGDBldLSh5lBNttkxl0jN7GMcqekOLGh
Fv8UWoUcSfz4GVdzBOdjQMoQO0pDGg3TTBayO/EgAof6Kl8TqCFNmBt6jJVYSDcb
2uDDYnrLcBVkkf9uznW3/s3V4KjT45BfVeZ1kfkdkRN9PO0rJf0d7vr2t6yxG79W
WN+u2G+DB7AS72lR6W63pQkzTYsbD3sP/7PG2tKcKwYkTEH5T04+s++EKX3I7PP9
6NLoFR2G2DiKNehy5P0sIfIwIoxa5wlBi4xYpORDQ/uPUGsqKYWePH2IVL6cXb1B
n9w3mkkMET2mEXAX98c5uqRK/mbo4IaRSHEXnSy+XAoGbuFIGKcD5VRUsnlTKZRA
P9NeBmNVeqIb1cWo8oWrfnwJiiKFjeoPyivWwtYfIYJYqW2fRHRhtkf7jrd34zVA
erxt8s5W6Jnky1lU+u0wr3qa7tX18mH11qP7tXGcBV11Hm/MDtXFYKqgV6KUr8rA
5hO3kWpl53gKJwNKwVergE2aga3EYsONnAoziOtQMqd5gpjIig8L4qDIe2I4+oE8
Uk4ikvZ794pIr6mJfcUifz7c7tU9FT3ndgGUYlfdlj3qoX8rAlCjDXNvEeK2QAJT
QChISRVgx6b+Twl0MjZPabzhVlB8tfhHKryim3/u9Bqr0hpEbXGfhHKLxjGN0ufi
kTLgHJcc447OzgID5yWsfQxRXlkPKbi1+g4o0M+w9K9AFa4Wqicqc8EDQvyoo19j
QYiEMQ79b7cgs141ohFzXpdM/kerJ0xg7k47gZfI/b5Vl1hqokxdSG9nJ3M7Lf7e
9+S04pZQgH3RS2BqTiCfLL2oCPHAtMM/WoDV1Q5QQ6BZr5JPKNOSAQ1FdSKAsLjC
7m2Vyjxkq0uF7oNeuYlcgKjjCoxJ/O44iwMiYJARsCbwccJiTyuppzmVL9n0Xn+g
E4mXyEOBq4bMQaOqcTrW/d2viXNseRcjIFMt+BQrukW1+u//L/x9OStuVCPIt6hp
2W2jzt1a06Wsfo7tKzk16WhZqwFeyu4xO+IFYiA+PG/tJjGX23HVRt2qqHGH8cNJ
e7f3bV9JBU055P9ZWPMriyax0JV/1n2dKzcpFJAz00gHD6aRVVBGFXU9GLQ0arhT
NslK6Te9OeThkUHOUkUBkcJqdMr6IZMNWI+ToQNfzg/M9gIUmOnluROd+VifqLeL
kJxDo0Z+bKNbKRMdz+JWHFxZMTt8qFEipfIE0CkaMCMi1LfEFICyipK8EPB2dB1E
+/o9arWOKhFMiQ+dtKncrRj18QFTRkrqCv9irdgpeN/tn1AVQZS4Z11v4JbnTAWc
mbpyeMFWB2M/85hZ/NBodzdHAc1r2an9uOVpFib61XPKcYSCRyxaU0RuF+0cTq0x
nC6mfk8tXqadhamVD1BGYzSMnfeMDqgM4Dll2KEDOQL14Eq78QUvM/4l+AAlVAvz
/rddBIoOU4hCWdUhbEwgVlUVY9G+6STXi/4W2W6H0Z1FhCWaC4A54hUsNRvffY6S
wW4/8k3fSo0+oDlCN7IV9dE0UcUxZ/pqkBvb9dYq+jJx/eL1oQP2b5ZHRoyExytR
/tOLbbsd7QkMni5U0mFWUJV0eBM8yzsq5RpWhkmAx+Y8/Q0juSdV9Bq1YRaqz9Vx
3cfGUA9EJlTS32xas9Znlfhr4Z9WnncrqzDHrC3RiSNu3Q67H+KIYitxVaf35dJK
Sjh2cqMKyj0nEtSILD3H9xZh4SQasZHXpEGZrm6kuVAeVo7BsyHnfHHRNmL6nw1n
1tnWJegDmjjKzzruo6UIv4IAym3W1i0nGrSiGAkGgBvH+Oxg0bCXFSslky5k1TJX
8gldQm4Rt9zv1AxblenwlNv4BtJYpJ6q7VecUPYM6NusjblyiyyO1pDFAYH7Nv9h
xAUpEonb4H83POqh/2OK6KoV+ZGp08VKmaWTIdosg8nVyY8eYM5HtxVTup12LhiP
o+UthHhtJTQwODTHBDHxkS+YHwXmyctvE3pCDVW4fs9GP6t69kXmcrwK/FteTQjy
QxQ9UdvE7SFcHguSbYCjP/Ej6djjZfpFXFQdinicSzY3HSkV+o0b0o4di7D+NkZ/
Ke2lWge+guYHfHpwFxSdjBan+z1hUAPVtIs+NKeSb8434husXbYg311so4Wpuw+N
Ys+SvPeAv/304my3upab87ICNttX0JPxF5CXL3OK/SKcCyvJ/GCCy4nib+f2zKk6
ePkc4nAbbFjvFuqPxMCaQ5j1vKG4JnNbaBtstJjb8Nj7ERAb+t7We+OtkIzmgl+p
rS1kDisjnkKTqPrbjYnftIqOtn7UO5Me2mxQEbrXM93uRDrXb2CdJn6u5oiuyPcj
ibWVCQlAadOkX2VewtXvyj2dKZD0cqaT4HME38ZKBI5TB8ZWJwiIdtbgtKgaO3iS
mL2WOl6UGOjvdNmswE5ZHrSRUVcwTfC/YJYFFUd/S8rGig1zJORqW+XSv+T20Sxw
+FrL7cezk/1Khfa/l9HQIbI28MnTsOkyY8onwzBoU5WRlvl7Z0necTViayMOsV5o
v2zZLBGQnRkB2eEAO2jyOh8nUe5ldGinBt5PzxgOiqiYd3lxM0UC0JzMkpiU2rfJ
+JDidgtb07fE3bBC9cLou3CtTtYh3hif+Ei0LR2Z9NQ2LYhCFIYsoB8NPEL0NMK2
Uoio5TBAs4Aa9henQTrJgINTsMWm6yfywLcjotsXNReLryjdU08sJIlXzbx3Bn+B
gQuLNcQ8rkGVqoXHk0unW85jVhrQiqZ++DPLsT0jf/z2PP++hLWc2DgNZxgtW4e/
Z3u9STvNbnCkQhTsBEfw2tLoDEpWVTJ0iwSuHtZ9j8qo3AT4Qp/ebtb6Hu3PqTAq
sd5mahrnXqeNG+dcsz/ALdN3lEcs2a1coQ63q2NuF/7kDf3XhQY+n6UWOoyx3I4G
nLlcqEyROxFgKwifgiWoxtEpeP51L5D9HBD1Fim8k56rzf2yicZVEGkBeMcR9OA3
S0riHUWdGE0om/JixJOODFYsIJ96ZLOZO4hBXfAlS7jjmIUB3C3hkjyoFFQstSW7
07VEDauogxZppRFYdO8NDH49v4ilbY0fGhfzfRy7b2OT/YuMDp72VJVRRHSKg7Wz
2vChASWbj7FtHclo5efKujm5ody6biWN19EPWM2ELYyLxC6tvxOiHW8vUGjIfI+d
sS6KnYNA6rQDZzN+Vygiss/0d3LGsn5lQ7V0PYhMx7YqrUZnS5C2R0R3l0UqLQOz
ETGya7KoWXPR9ERWzkSSu5z2yFpXoJw9zMfRIH1JNey2hRV7Jp3C0BpWm2nQe2oW
+YBy9CYTVksxUQSezwHcquWm9H9oJ9dd90rZLK9kTRKM0CQCkyb27HQ4hqXV2+Kd
EdM1haDj1rrGQibSIVc4afn0N+o3BDpVW2wObwZrtP7V499BQSyRQPipNLpMrfOc
Tw859U6rZ1kBJ45fl7t4SR3IueUExCwjlFemdbZFl+9eyeeycimwiA47U3nYdmqd
gIxxwLEVOC3fOcolPIGHmdq6JAUnQIZ87lUeejHOiPRLuDyaAhsg1mFBaYXpWB4r
jDj3rUk9PXj9CiKShVxsyStvLCZQ5qYT12OPgSjSBzD2GOBFypmcgHQD+dv4+41j
D7cPx2VVld7h5SiGh+RGA0MZjkdX6IlhrpMAOpxx65VMaIr2zib3UDNXzdbfoEFF
SRg0rF3s+0qruyRr4BHLmtehs8hXJdRws+p4iNZgYHTWr+auINgG41GT/JFiLORi
BBVizmRiXvLLn1/UNmB5ReNBaHUpt07VchMRe+Qj92bn5n5q9xtuRh5inEKFBid5
fx/FJ916u6AaHdz5WNyXZJdXIizuADp/5cTl65j/08vPVUBoxXUjDYayBBOeW9Af
hE7BQr4to7qeP9OOiphqteIC+iemNtVIqPaPqPueaUqBt4Y5goxU0Gy/vvZ9OMr5
MLjtVfXDWIfZRu1Vj2mF6DbacFDqVs9HkgmI3+dEKlcylrHUEsxxXttSzvABUSAR
77ICLHdGUxwSYF4li27jUmuXLF4tjoeBbC4F+CC1A92ySD06sglyEObw9hgXmf82
Z3LpIv31gBUFrBTSY/jZzwjFFpNDV+MKrSAL1i8S8mnvRD3GZywCkNb5nZTgRqAI
D7aqggLJ5c8QpFNpCmhBuZILYsvK3+KXaNkPx96HXFV5CEL+1czxWglrFvljIitJ
V4ljzdfx39K7mX15NpZgaauSlkCUhkqPntaNAjHoVoxG0crnqaUEFWAY2z5B8t4T
2hXQor/afeKtFyDniSUh5SV881IvPqcjVP9KDD99oq7xxQyEpnaerAiYbG56AeTB
cgIYC462uzBdYIi8/lrd8b2FFqBUJbXydfb0jDS+axERZ1slyb6jtJcU8CM2pDvo
Ur79JQK/QVahxeDqPNEhwOVjKSCaSix7PI164ySe5ux/BadGM/9qzQn84c8Lt9Y+
BWtS5Xa3VbfkdLRP3pRH6Tb6/HfyG+BurPtZgbCF/dzg1B8rrozoDNNXdzHHHZnK
bNzkiY3WU5J/v16chhVd9EhHBP4mAjsFlYlHq/g5ycwdJj3TMW7bgW4ajKgPvMfI
fw+KcBKTJ+xNt1inNmmDwDiSTn8budZWKTzaD/jT19xHUABjfVsROTzAqsrz/yW6
060CZh3AxSM/do1IQ2s8mNsJXikNVow5CJk6eBbXGpf2wuyi0tzhG0c9T7ym+5xM
DboS3oFYR0nCqR8b4DVHX06KdFRLYBqXRdevbYh1hImWuFyXOhYB0jQV4BHkCs0r
aQ+BkrrLb/FFY8S/lWuRbKVfqXgFcwEQzrw1V3B39DfWO0Ortjx+QLxV7p8JGjZk
ovgmtFoqPADLB2HiS1/97vcnlQ/y+ohB5Fl5orTBgu8JuxF4GRPUIox5+1JLdt42
xBr1PvrYTKbPYyyWZGyKleL+IVoNFCi6nLMAXn8ruUNpYjVx/n9M8CLKZO35Y2PO
OK/9+X8HF5K/f7mK5HY3OU3X02GUKsJHF1EM5pPvIRhfl8F6ckUpnV52QU3C2CIZ
wZJdjSCiXkAQ7MwiXL4E2LUJu4qCaJc/gDlX//Lqqn6tuL8199xJQ7laH4t33FPO
raaHGNeH6TkHTDftFsjaaLh/NrHwPdXPXlcklacoqtx8t9fqOJ8N2lkP53rsOMJy
6kiypAdvmyk/qCpQTQQKxKWnsb1CW+AOPLh4V5JngG3EQagb4IgVybLTwcUtJVJc
XWkn/LRzI3rfyg2xR9RBhBK326w8JSOkc0OgY1QC31GDorEj3NZZi2/5wNRoZ723
J1+Wk/O5xro98oUiOLldcSg+pOFkLlxavBuKIFtUk5jK8dOSODVcpjXF4q6zuuaZ
RL3Xkmw88WeXsAcUnBS7CDBKV/IXxWfD5mWn1mkVDTS/M7LMDipK5PDc+AFHYghD
NHhr+SBUVDeaeIrghzH98dQWed80t3n0+WvKGL97+v8uml5Xapd7hvC/m47RZLW2
7HggQlSL1YrJFZaS6mvCzqcy/BBTtVgqfhX21UsRkm3QsgQv9jRJ8jz+nZSMhiM7
B5EFSaj2rEXOK493bUT+PZLVWkrN/cbmkAqGTM53HjSKKTAgPW3rbtOhlW4Of8Gz
Tr+pSYj6qDlK8rY6R187qcA9C2GBmj/1nipkzzYZ7x2s1xWniBBfXjrPdu8ikMGa
QbC12uscJmvu6mzZZ5lt5pol0fCFiYPkvWHCpvdv/k9K4XY1XPUfjLi1hNj985eP
REIqGus89xqpP/wxRrD7fu4/bZuaQUM5fm46IVXfkHHW9+x7EBY04P2E4XK56hzu
LpDTNbhBQ8Yvdq7GBO3peCvorRggInBfgS8Cb6eg5IDjyRwrGhA5Oazp43GDmHHI
EUHythKA6n7qf7B9B1cts+Kl8Qpphspu/QUwjttVNkMdUGMWBnZ7dIQAm2YbY2ir
DXs8TQ5gllmnMnQHREgszUWCd7+/RhWSw128ru+0bt5xfcjSvAPvAKX3kRH1ILMF
7EWzAwhKAmuxdJDmI/c7ggETOOzab93pH4RORYeLa/yg099Rv0ew0uQD+3XseuKM
qSdMHaKhE56jaukigcZqBhKOlWY31Wx+XANXP9v8U6xr5c6GCSyj1ZWTBd65I2/0
/BEn+uTAmfP8AavzaIznPO1LTtmeEJtsmbD3p/916bUGpSYrBxuWHFQwZ+3dbRX8
TDnOjyAkIW5DNCNagd8iilaBeH8PuGiOwDVPT85lTndnd3QVrD8cwxeLSwp1Y5pv
JMWFRyxP5wt9+5Jt3CeYlaEzGmR135n1niIkBDxOEJyIfcVW4fQyhsLADjwy16ph
WSgtUs8WamVxi/RYzX0MvZBCcmgnzYEXj/n8Q9PFBSq2FCFcUUL8END3t/59zcrY
lwUqrT833Ur/ZBaMWs717bKHhlzEGwbOTWpeAb11o65r69T2dGKwtLqWgzKrsUZw
tBxnz1bYP6XEO+wMoP0jdrPVV0SqgedK2d0CQYCWxVTtKaIhsVl7xIb6Y8rU4qP1
rZde+nYvjWp3h9Q83pQ8Vav9L7D0Kz9BLVb2ILht7LOWnX5Z6S0G5PwetUS8O5d9
3/f63YpGVnYe4Uhx2049eX7ui3crsP8di/a9v2acE6Iz0A7URbliTAY7SjpBlTyd
ZerR1VsCIA18sSmN5N3MIegqJZNECjmUorddT5kFWfocdzVEqaDEM7VdQXWNBQsV
KFnb5fCgRtCYRm+Av+jUWDfllA5aH3n8yQp6c/us1Ra3QeF4jYvuq88zz8niP+Me
ibmscqsDIRWvf2EIcci1VG4b2D540u0W1MhEfpTHCd9a4iCLTYXkNERjzcya0MFA
Z/BAxdtu1L3DexkpHQ2iAFvMEsBZMTLrZGKp4Jg/aIjY+uKaq3KJBbx9Kv8W4h9u
dPuu0/wSHEHI59CLMnTDeSFucP9CVtHDHOveVupgQaP+DhdodP2/QjNNf/Yl7Ick
/KYbz/XVVxVu4NTzLFVqSoa4KPfU96H4y9bXg3koFbqaEpqNoSHIyQoP7rJiYlrP
7zRzyQWgcFi9hXdYEoFlJhCidZAfU79wQbEdvxaGautaogxZ2tPTDzHCWsrSGlGr
f8t6LICI0NbQdq+mfXigvQ==
`protect END_PROTECTED
