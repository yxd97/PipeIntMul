`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2E055wegpjT9xyW0zdy3vKs6LF0g8Bh8jrEW0/x9Ke0V6dFhG8uH38s+hdWdCZg7
czK0pLv0nUgFBcvCGqJO08xc2L8gzDvWCS0kUeHTxD7sWXfBko5zH4ZPGXiBGe5A
7Fl4pofrYahtLcKx/ltqUBEd5vBD48xYzMWPtBE9/1K56vQIfpGL3qxalEk7j3+u
vYXv/itlcooj6mUjc9IX3dWhKza4VEB/tIlHd8eyK0wDjoew+Le1eJD4OEaDCQtm
oPSOp8NidbyeUR4xiNDu6d0VTbMxYwUQt8vcPMTNfICJurgxqQfHyE1SzVPb5c5N
mekg82Owx7w0ug1RjkbSZBWjcXJrK6rh/1T1YllXl+dPF9UaXM48KSVr9kICxU5r
IIc2EUdkQX3VEOaK3hc4qO7p8jRXv029y9WtIBH2/K2mz7t9b/HnCadqSnUlHcf/
gxnD03lzTdpWpvFZw1niDGdeisuEgCkOfAcLSWvBygaRW0XPjGRtVFwTZd7glNWm
wXe4350Qqs5xGwZHCiPZt6dR7OiczAzRupHnL/1hCX+Omm/3ORMvQgVSnFx6XLht
QbDqX4jNnMqPRIoEwy/yyu4OEIGHZ48lPIN5k6rB+ELtOd6xbLxQBRd1ujw/e+9t
1sby2W4cnnCpkdM3K3Wf6YAWes8IWb0zoenIdOJxKDf3Cak8Cix/CD4A97YaLep9
`protect END_PROTECTED
