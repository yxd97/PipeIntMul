`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AAPb3a9N62sVfZIF+oCbmjaUTstd5T5cUdedAX744PmL9ctwYZ1JL0MO53gVeXfc
H7heTQGVFIkaaC6Bf+xS7jkHC16Q2oWxSx91vO7LhLTp7yaKMvTYOpgFBUadOxjr
ZRgQtXz3e+pUqFXi7+TDqWOnxwCUwOZ90OZXVrVxrbpSptgIn2VTbRATzt1qlIup
uIru0oPd01wQ3RCEYX6i0bIRyQcItWzmkzn60vAnFjbIyrPDt3DJCtenLg9e0C81
lP44UY9AywLe4u0tbkU9Ew==
`protect END_PROTECTED
