`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DfcpImwvfPGrpF1uPg+f5w7A7IvmldWbJ84o13mlgd36FvPsKZ9r2thKJmBes9TP
KJlvgW/SMlKa5BRMbenGAf7a55syRtSJKhqzhlzpfQ7XMZgx/YfRSMXcjh3BbT2J
4SHw7m2oH+0wUUDaxWI9xp2+WbbPL+Eu4ZG7rHcdWxExXwfa15emHtBZKFFDXAsE
IAezeKisomF83sO0wIvqWxOpFa4ZnRhwb9kal2/QWsT6wOsn8K9Y7H4c98JvOChk
la0XMeA0V4xZ/UYnuy/LOgM8jN6RWo45EaVwpMPuiUHjNsOzJoEqUSBrFldDoW9V
q0XwGnkvHMOS+9K31Ecq1n5Tmu3OL2tJqGe+JMxttVSutTdaI0aSSusn/D3dj2WW
3/ip4AnpLNW59sEyfdvTIi9bt+80UxwwBkeMbycBEqZ/dtZJMY+ea4e68Wi3052W
t+4BRuwivByji3ilGgAda22WCWVp+5nPd76i84SIqso=
`protect END_PROTECTED
