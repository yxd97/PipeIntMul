`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ukwzfuWOfjHZ8GuuYUazoBcXwQF0NT5Kc8bMTUQWE+iIma8vG6d3suZ1VT6wS7/R
EdVS7kubTskt7Th48+RcpsfBTwcgpEnsB8wbGQM4i+t02+To3flFyqNDVjyTKkDE
tHkIIF9bI5Pez8Z6EqCciN+JRuZ54PWSH2EJCweT8AlVYtfuVw2svCeOxjwHf4Lc
8Q49emq1V06ema6jCBRe3rkgtVEuhQjC8WK06PDEnBfN9BAt0NojWGBtECF/x2hm
k5i1g3BYwtVcLSjLRypffOsjckHK4NQIMibesiNv6d53693dKVi/qNbILkyxOYKM
5jaHx6KnqxIMALQylfG6uh4mzqWBfBpwt0MVVUCKlMCUANC1jB6n/FUtK2XfvfsG
0z8J/Uv4/sh2n+JVuTtirhmSj9VHOJ77pLCEgGJj0UoA9pM3AOxXkcv4SBCjhWin
NulMz6afn2O0IO6Uogzo8L8mM4VR3dr4II8CtN54KJx/jC0splUTiGIidZV5+A4R
`protect END_PROTECTED
