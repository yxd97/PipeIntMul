`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
itXCK0fM3BwR/1B1IAemOmu+J+3E7jFNJNqx7nsvyB4RDdTVSCHZKeoYPGojNhht
WjD0+mPcqDnC89EoQ8v9vlkjGH7TnAhsd4rENMhUKIWpV087Ll7c3j4Z2PPEUq0P
q8hdNmop/X/YNmB9VHouHlRL5q0iTNIhFG9uE4KlTikok+Ymn5MiIANqh6o/Ir2Y
MLmsRC6RxJkJBH9jCwQ4K6SW2Vot9PkipmsKHUTDC36Vg/cDTsVWdKoX7t2kuvuC
NptVbvBI2qekd3qEU4T209KLo0Tg3EUKepXMsjPkcDBOmeX/njIY0QElilpthIL1
6Vm61oTj3mEovnAvM1wCCIa51k3NT4KScPUPryH1EQDa0o2xbDDL8a5E1JX6JbSb
tVmES+71k9duT5i4MkFZvtCRXu5xhYJx7zJRv9RkUG2gu++9G55WtTDrEdOh+wD9
12OQ7yIN+PgiBymL2mQUjcAW5mG2Ox4GEPVLQ20CEctXhUYls/sfNhk2Ge6mpQjJ
`protect END_PROTECTED
