`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vpydm6NQMh8axnXBgpTBUREqKr4w3nCbeChb63QXv0v4X7c7HeAA23fOqtOiHtIW
d8cNKA7po3KernesQOur6ini+1ozLLEm5j6Y6vN6nN6reaoYcZbwGY+fH9C4l3WK
+D4tdqiqBqCnaibO7T79xbsX5bPy+06KYNicLQs/HTd7XVWCKdh0P4LIecBjpV34
MkqGqiA/IijSI98lgPJr1klg6dqHQ5X2k9ejiGwxygBhpUQ0Zh//AhyZ/1BeXj6X
QNyJ9bGEmVJAaYqYCxf7gwgRhpdJ3QpmPgmyogLe3+NbHUBK7sYR7wCn9nrxJ2R+
99DZYDxUGYYqUaFI+VSGElsCnoeyNTdjovf47Rh0Q8TEdWBCY/pWSL2KzD8iOxLI
4n51lpcpDdePre0PPXqYQOGCZmwlNizyrxBID7J+8u/lX1yx15PE4D8NcGEhUcLy
keL3J/NBOsGPBObdS/BHzTZJd5GB0tqXC68V44ZsTknu71t09IV+r7dfzhh6LFTF
PLitUOrrYjdu2xoH0GhufqKf9w1BuuouDjR0cHHl2An2iDfntjUO3x1bPCPANsjY
kRWEB7xMnv5ehCvB1bD34AgtbElIqfsUnQppAmVLJxo3lD74/bW+Le/QrOkkb6vt
4vfzK40QMZJeyDUiwQGF9hho2c/yFx3lKsWK3FAASuMO0J0n8T3u4ksV6832RMXp
BziV8iX7NZi2r30PH50chiM+CvFCuOBW+/KHI2QAFJUzXTn7+Mbk1meABdu8GLOy
oxhQ81h+Ps+/DP7z4gAZCCuVEWZa5itpyafekO00K3idmMRww92MufbuifB/Gj8H
TQP6Khe8B6z17QIGaNOHKyIpU83GQIpbCaNlEBRW+MQFdkTGz2y7shw5HydV64+T
/6bKja4eLIu7DYKAPkd87WJ4xMOWSVo4g6IBtluRPet1Apsh7235bW+X4cQsBzd3
5/4116Z18m+AYDbDQPK2TxoGpD3IPCaCAEhLWprT72B1ngWtEUvJ9BGTIFg0+xXM
L49UQaddO9Cl5i+e2Cxafz3wqgVApF4GP74iQH6y3v95CcjTJiMuQ5+HzI764F5O
bvr4XQYa75YFnvbESWAA6PgARiqO43g6P9ViC59hHnNOdUzkjMdkds0ofnl9gUwn
gxCUAAPrqROrUzDLlILuCouRK691QxVSGeaZM/H9jbjHOY1FmU0JLYv3LB05sDTQ
YD2HT23EkiCAILND6IshqIZeFbaNvX1Fu7hFVwlnBkw=
`protect END_PROTECTED
