`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfDhy8kGkxmo7WUs5Ho1uP7sXxGECcbCAQ6ejlK7IKTRnW8Ayfu0PtoPu52U/cKn
BrqiKJT4taW0vK45boJsD+QYkprN4coKiu0UW+dUzAz0anKVTl7zP1HJKNGtXqRz
4cUF0eBKFAvefYOkDBwAlhBIcdhS9/KMrU4e7sNEUyKC9+TFqv+sr4jxOBt+LAGc
zTG8XsVAOGOUVBFdTq9wOUOqqd+b/+/VwQ38bF853gRugftxZN4p2NeMWRiz1Iu+
AnoOSSM23a8k10CJda3J1erlrUqQK7Wy6vPpIjnhprrCumE3jQULCGtpoMgdfSaO
GEzRBLpZvLN3bSeyaQ4JIUcKVxGZCXpkYvFRkoB2O9CKZAvhmP2LCcuYSFqkCjkZ
GS52SV1V/b5kY+yD3YfbGVE+OM4fhoiJgn4gQSVIJ8EIRDHrlfsf9BA5NAduz/ai
7ePa2ZvY15cmXxyhs7unfht6lvSmP/ibaJcBFfrtM0MUyfyv8diabkdD5FbpvhAb
k/UeXfbEesyLJ4xvd9m3MChKm6AaGTkB5izS0Aafix3OjgJwsq0S+N4VYNtixSnM
fljn694+62QYEtYhDpCW5YwZVY6jSONIXzgUNYJNa3YokDxySUmZSZAGLPMcPh2q
BrKSbTDzDOVfJ0c4cg4Tvg==
`protect END_PROTECTED
