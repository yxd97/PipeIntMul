`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+lz10k+EkSsNOkyRlZdhETsrsC96JJv4Md7ofYiGekA/uY+HI16w3yvlxOWceQB
Dj0ikhURuDKN/jIYcT9CL43XS8nYIOVhuVJqIEzCrKXQ+WV8aMOD5bkeERftHIL0
NZnQQBLfbdRO4/SmjIeRaEdsIiDVs/xQOq0QMJ94xbGFs7r48KoAfUVUNZwi60Hn
xR57hQnnY4mIpoQuFodn6Hi30XRmhcbFnDsLQWICvJ1jGFNB5E5mwayN0TUpBYSL
pS8Rg8x8U8vr907a8axQLCVG+orCch33+2vyGsAGASj/U2bQK1r8s4Q9TuBWlT0r
zC6F5lZT8Y4yUI5v/XBym1q1sF2MhlNNvzyOaI3HeoKxFguV4FcB39w68jv80Su9
UUmKMMOQSrN29ECiT1sglnKr5uCUhYyprV3N3S3OQOyQQGSEeyRnZARaonDje3Sj
w2KXBdNm2aSHtNeKqj6bKUW8D4rkiz32pZ0tyniknXRrsoTkDDcTgu+cU+QNF0df
T0oKFbUmBEwU86kNOA05wQDBjh5E7xU8XlBPxO0UJRzgEYlGgk6iz+rcJEdZKQHN
/iwzuwSUDY15ADDgtojV4L1v0spFJYtnI1/48hmjdutBEThrQbW0B8kgIKpLv69+
Quo2jjPxRzI4MXVzYZeUq+2zmNkLEIJVEh0+wv4C/p3DVwBaDFSJppk8f6usE0ZH
fwNUadeh2l9rY6/XBsYl20NHPrbKNTGqmDLAd1b5Lr9fTuhawUKp2FsppSeWjvdp
7ZEyGniFlANoiJwq6GSrTfoNJwM6c8DvPdJgnFcCxunFYOWpc4C0sPdEVQ6cLCBU
gbTCLKYmmn63xIRc6iKD71kQzV9/nZ26PApoDQKzajd2J15w904tY9voU/kkmRH/
euPT/WLi+Ja+Vou3S1xCqQ==
`protect END_PROTECTED
