`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GeLKaHVd8X6gZEP37DFpJ5RVnOKIC2ZbiYqzrEN8GFD3TxyaFclqRIjyIqxXn8OA
pXyl0lBPMI3+TBua0TTPkW6CIUmL9ReCG5r4ykBQrKPjK7E8fWym3sWNDwLiSC5O
foKclsude+LRwizHQliwh95ZHaY1Trs3pihBrbL3gS+vZ28sDEsI8i0fBwRm177R
9UiQ3mujk/RlMTirGkHN75nBq+O+IoF9Zb22VTqHZE9lTbK83+21NXHt05M4KyhK
oDEtIRwy8gEGzNQUJDMwMjOPk6eeHPdSxPWIYOUa5mng2pbAqB4ntP0UFxfmcbwQ
p6s/z0Qk4Gkeclzy+fk89W9y3j4sJFJSV4MJPxOI4qaJunNt0BIY7nReSltyozgF
ctOROvsNewcqI8IU3Od2GrmrsWWh27TFvNEaOPpuYxZPjEC3tLfItjyqCzdN4VxE
7bUSZcliFWb/rTyIaI1oCZcllvQBb4B8WQ8ukxuwiz95cmh9rpZz+hIUrhdEnqtg
`protect END_PROTECTED
