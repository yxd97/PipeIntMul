library verilog;
use verilog.vl_types.all;
entity OBUF_SSTL18_I_DCI is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end OBUF_SSTL18_I_DCI;
