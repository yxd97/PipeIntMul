`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yl4r/gUAbEzGeb5tFxkmkvGOB+JRq1mrS074XdCsS36gIcPpyN3w4FQDH7IEDMr
TFzVINtkRc6uPtMyDVeAfaFvSJDoAUnFF0Ojus57f2ycwKlaMdMtR7FR0VtvjWTx
WC9mZx/LlJqQawCMeNh35DOtrSO0Ozi7XE9nyUVO/GP1MhPCJCXlE1ytkfFMZDfe
0/QP5yxE36F/MFd6NPaSIDlTURYpWi1lglHLZqfEKNEr0+PZxBtHiijCKSc6D8wM
mlD9nLzzA7GROETrtam/TzlgsVreNQGo5K1NqzNPJEkdgOEEDY+Nl3it7YULL+kg
qRvYxhJUsi2/y260VgcboAVa0LlNbhadKzw/Jaf7TH1DGiJPleJj8r9A5xuQv7OU
69b3UJmYXKtVcjRjNgBcmA6ZaefHrT1FNuWD8iL+fVedautxsGQYfYsVhOG2yyyc
WJ20O9SEgxDPn4wu8XCp2FaIMxXKmdE29wO+XYDOYeVkE1uJ9LoSFoClmjzheCPM
XbT7Ccoe4Rc1yPyQJCGRO7je5Wjq45mqdMkeGxncdaZt/2Qh6FEU/zkuV49y2CIx
RUmZK62k5HexFV3E+xIyNHNqfR51z0S2wq1jaAVuKbnHZMmAVVbLNVqSAxaBgw+w
GhtxAf0HNw4SHk7yv0HIBdG//6O1QxI8d3wZrtr/UOvmJ3AA5vw8GkgzW6PIHSvF
lh0A7uZAjamFe1mbPT5FTA==
`protect END_PROTECTED
