`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3zS2lSmQsnt4ChElB7d0PdXiu1iA4jMD5R6IHIizyVcw2EZXqr8FFagGK08KC2P
NMsSPPoPAvd/Iq1MvyqGnf/QB2OwR/q1jbMu+tbtxfOKzGnYB/N8kM5fmVajpQNd
egPJeDrIrOLzwYjV0L1zL0tm5OdQddq3GMS4rYhRCEP+++RnLQtZYul7/L9DSFMn
xK0WqXau7Tlxv6Cw2WP5gTwPWhQtu9N3IRQQnTWcZpWUza+PIF3K9RTAZUrf1LH5
R3FR2/M2CDPko09V4eCo4Rh7K/PpewtdwocYflNdlkvUH0y2acW+MlMD9LMDuJqa
rJhv5diMSAG1iDyi/qvW80wpedEo0ndwMoisQbkcvFLol2ba3C/HB+HDCHG4wx++
trWEsErUuNty5pQx9Vth0dkNUSyN/ux25RY3dZLRYJR1Vu0uLQKuvP6xh0ILMnGK
844kHlxK4jaG04NQ6wAckUB7cGdEjTH+4C2snaLo2FfUN2dYlxxBdShMKgq+6OYW
ZqIReVeHjeB5Rgq/wBJJnRfwfNsuVqa2rsnLeMBp8QXXffgyKLdacqKQaVKBY9gh
AUckwrkEW9LVsK8BsteMDkW8VOlauvBw/dl9PGxiqwa2etxbsE6+IZBK+0M4cIOY
iyN6hWPnTqRpG69STruuqcnSXh7YdYnf+F1VMr9UMUrsMFqaxP+70mwBr8U6dz7H
MJnFluMkWdEFOVjeWtkzDUYzfrGrkknhH9spPX7AtxbK5Nox2OlRfZheYzZWZleh
1kBHEk4uYPhwblE2MWk0bG9iKaaD8M1Ple3NhoHEahdxfVv8kyAGiCaigK33R0vE
`protect END_PROTECTED
