`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1PsNnntUOcQ4IDrD8KDWU7aYFJzMMNgFE9Db7TTKRAOUbm4ZB22ktCUXLj+XdYr
8FRj3+8Bq0svZiAD+p55TmmH0VlQe6rY5iUDuMoBIweYuClwCpvxPsEwneaoAXyL
ZFXMPw6nlszTKXEv75HfZkLbi/uy6y1KVqL/5EtwIOVtQoHYxLKFDk+HS/ypXoPP
JARCPS3mT/XUnNXGN0uZUF3wLH4MwiDt3D04/FktX+8u0hIVvzJHPkEhyF7vbzl0
B5xTKzp3K2T1S+ZkwzZNgfq8ieGn+GU8krE60ekz2fAdogqvzBvTi9fCf1h2D9y/
qdnvLaQUt1TbM1u56wdSWwSV3MFu8xYpar5kncX++HdovhTVmabd8dw4Ay50jLd9
faOVqg3OwiYyr9CpbvkO9GSyahJJfwIR2+nxx6ffaNknaxwD8eGT2/Vgvynk1a4H
PazTJuWQuY2E0ORLlNq2I35sNJsWkX6KQiILWle8RAg=
`protect END_PROTECTED
