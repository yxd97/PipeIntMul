`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/wp1h8hJxOFZyq5pMQeMEifiNjVD6C7qqmQdJDCYEkuWaR0w4mCBE3jV+Y6zpPh
nxo8VYZ4vowFR9ToD8R5E3iXZIhwIjcxuWV7h82E6oR4r/20spXU+4UXKDapY8yd
MeMSZ3bUaeyzzyrA0Tl6vMK31zUFUAuDwu0RyFZHjqiHOMbUjNYOeVBWCBrR0IK7
3XUgbcletIfwoh/m1Un5WwkAUFXBM0+VgxihTQ2w4FrDdDQpASlF7pg4rxulN9np
Q1/AuO+Z9kBf8QkjdDrvZBD+snfUD7eg4ca8+YAn9tNtCa4/fYT9DEo+zIvuEmfn
FqTGF6NUGvRjNtp0Mc5C1w3A1C1vYODKuVry1mYROTupIXFNrcWyGRSGX8dIypYP
jUohZCwkO9OsRZ+881cTqOz8mu5o/9Vjjomv0+Y/zfw9BRaYNctM63C2rYFtY4Fh
e8HfuRWU/+Us/7HW3l6b6XetiNDZWHPaleanVtpznwrbOIeaaN9tuzwifO3MZZSl
9IgD1Ondit8SJDNeiu8lTq9xJD4I36jRVsUFge//SJWFMWZ1qQy5stotW8GO1/Li
QPTLN4q81Efet4S6MJSZOKvPQjH5/WKQrpdzZrWZ/I0DjtXIdYVfw9IQx4aP5tIV
mqf1vwfZl/dVb0GOw52zLNJzzIDAR4HtcMBizIPE4Y3SpzRjTHUflXA/jHBEl/Xx
XYEiIuWQCqTx/Aup0emANAINuqNQdHp9IdwU//HLv2Wp2YzKAvI4+HSoXVuImCgJ
/IXSES5A28DaU5eebtio3gOiiOHBVeFmzRy63TkN1KT0p2FHC8CP5AQmSXgSsFYO
3Vr9FnVCKxKPj6g/zpeYQLYrsGo0WI6vT7Rats4kaVa49bJbPqPwQ8AvP20rxfE6
7+RRQGJRiW4iItDXRZ978kmqcqEXgqjO/+YH1qetiQSg2Ha+mpZ7gvOuY7ZjpRXQ
Oxv0we1DuCiG0NZ00KNO3nZd6DnxW5hd9b4tXl6cEMTHsdLV0U5VAXRyKJUoPStN
xB03ikWZEvZiQBIY6hiE4RtVqVX3ugQhG5hMT46M2RsOx+RCFM0cmltISuIwzP3f
j8zEFaR5jkWYXHhLWKPGGywpwtQezdSfNmxt2pPx7DD6OguSHmWbJtt3W3WiQLQg
U15GSAIokyke5HNNpnlD13WRQIJpOuhRkPd2k+7zkkrx/2viSflMfdtdz7QcvWpX
lzdTFT5m25kkudVXcH5V00E6GwP9qW4C5LhbU4Q9b3SIlE3wnisEqE/Hop0i810o
rrSI+Mnl9fE56HyZpVNmLxA56Ftv0lW8ek5csxl8/jUSpvaWv9BtyxJEo2XKg8B3
gcrspRIpbymuYFhAEBf/T2LLi0EVjDN31az/YTrKzF9YweBu66ZXCSqeKyTw4jeI
EvQepTCrst/mlD9DqiAPkizUhkdPvkAu4X/a+aX4NJ+bo3mYw0jzMj4cq8yKoqTa
RWXZXcmuSLC5lWlHZgh8vqS9yA3RtEAHo+9IFu92P1Ds6A9hcbiH3FgLWEDAY4ge
aJMsI65T3R5rXCZXcKtXshxf9Ac4pumNJQ6pe6Kc0nvOls+YZP/aQUHbgxiKPl0T
kFMXAF7smGkp/38saiUVda7FdkpfDNtsJDLZn603ICaBcz9lxTRzyzzHNaxOpK/j
/Ivz0U4xTPWbxKRtIEFZde3JZ/P4wqZGBlz6/PXogJWqQLLp7xJ2mCHCefLwUfnw
VecOeR4t7783n+HsOh9TIziznLhrzrg/yz2NSGPD3MO3Ufsw17hq1VQObfPbpkWS
KV1C6G7Tb0Mb78DMbmPe/KXYBxwyorjGxeVu9pKYZlRZenxcsYlT4mdWE1QNQFSW
xNkLWAZSSQKJl74t8pl78rraZzEc/U7tFiOaQ3BT5v+gkCRoi1RH26YNbRAV1cTn
j06wmZI6lmgHVXObjJyY/DdSCvcXIbgbhj1P4g/t5D5VqZpZFBS3C28g76SFBqcf
gHwdkMUiYS50IKtasVFm4rBw3Mm6ydIHWsVaJ9mmIzCcT+ePJfVBiuJqDTqZa0Jx
kKfmyy7OrOXFxZ2YLpElL+ewlzUsSy5ksf/YOHDmyBMRekU2SDNjULrKsMQzsR2y
XDw+qKiHSE9v+VxMxStkiuCeXgbbc8gWSXyznE6Vom/1eeA/4MOB1IZvXrG2b0Rd
xnE3SfmvYkdP/IqTUmydDH2Q9iIH51lRKfel1RlHE0j916tRCQbKHTRieFBmEjXa
SyVaoPb1xSxaPWmW8E8h3CB236H09ic2CF7Py7JZTcg6is7zVdxwWYqL1NMyzN5q
rvT2//DP6Z8tn/yqyq4PUNfPmFhb1Eg3VjrOFmHJ6fL5rq7ZPzKWZ2Er32+zTHlm
MWVFOG4Hgy2bJWUHpAZVbcZPr1Wi2eyB1rAcAdCbbEWHpRvmaXt60X7l7BOi6w4E
cANZOEFpqYcMsXuUEUPmjGERvpAZMR/cUD/QuqMYkNhuxQn9yRDBRJC1BhhOzbUD
0orkTjGyyfpEFag0la3ng2IMpLReHeVvKHqRpIGFpVDT24x57ETOd+plnNLWQyBy
keZO1wEfKYJ04NFUx/KvJ3svyvSmYwXvgH5sNRrvVyZZKBZ4hvBC7+GDMEFXklp8
U3Guy9+VP/agHgd7wkJLK9NK1f1IXAjcQbKr8GSOOO7MiBKCjY1Sbr2b2rpGk0KG
/faEceYr01pHl50COnCccaJsCGpc6KbCMtCnKkUsh7V4XzcFwSBHydTS8wAkISER
rjzK0C+AKknDkcdyJPx+LxYfwG1hMmM7HesSrpHwk8mZdk8p6elOHd0UdGSl3uq8
Hvb04b2V4a0RQDBjkqNUmmdqzOUIOjFGCiB5vZzRIL4g10AMMuWEcd/UlPkUF9ET
mmS0FdmrUP+t/WMq/BVrp+hAUi9oklPgm3R8NHXcROkmx+R8bE3+cRoRDeR06nl6
1T2R8DZF0ewZuhFMPqTHI2YNcE3VCjhQ+VmiYoFF88hvgEZFYrvpE1yL3hyOp81H
D5/17tmB84ZyFN6SqmaPnNrrunm3tLaBtOCE3W57t1GDtkff4PVl4lw8Bo748ulZ
nMzJbvPipOjtoosh6qE5KBdXhhZ+jmM4ebUna0lj5pxpeNhx474O4xaMZj3psBWg
+W3E9Pe6r8+ot63GhK8af0fsbFZIzX/BUqfHxQ2V4xj0Qv9uVVA9ZojGHqloi0us
UPM8ZC300OHAKLcQrO0gMrK0TmjIxn/L1IoJmPDL/lcGRvPj5S9NBzXiGqj8AG1w
cq4s3L1HSmVKwLWxzOf8uzPYKKJBzc+1LaPdruA+EzUomLC/hlm8wiHEoBXlkAZ1
kLCCqgbvs8KStFC11ROXYIfGsZ2/uSWIiA5wTDkqwlStRqQEdIVQP25R0ndDD8yM
1+STxFis8+TZ+NUb2cox0LyYO7UPtHyn1xam6exyOcbIlf+dHa+vm49YjXADWjmX
ftrdovT3eGqyMKltImOBN7p4FbqrWna22P9zBFWxifAKt6m535CB0D/n2See1t67
+GfDM3DLQTWZ7geQtqL54Q5hcy+RGRmkDn+V71ipXcOwHpEeo1R44XbxXqgX0VN+
1O2jmzzhajD6MOS7Ts5d8X82ECFze53jCcr5ErX89dvdx/n7C5ANM2esymTXMk1K
7/JGTMPnKRKHhcCL2S1+m7BmwfBF5J7gpo9U+kbwfUo/qJ22TNafyO7C3CBE2Tqg
5JuRSn9aztWlCaI+22waGum/yFltQw8roCo1F8x7H92JT3AGII/EEz7ylWqR0DBy
IjThwdMPPa/1d9x8bZV47YJfLWS4q6L9ZtIo1pZrfwh+foU0erTyZZ7KeQB1JhkV
5Pk7IBL/H15Y89LvEcbEhlDDh97yecxSoYM7qeto4sRX0QlxV6dcKAYQ5w5MEAJP
63NuY6E7IcE2dtRIW9RkmjesZ63afwx4oSLdWyptU6duy5K5ERkmxJsSAJ2JizSh
crLzEVg4CJIr5hWvuaaGgbR8pO5rqSWwRPfN3gimSRtNJfU19iKAKlw/SEfP8rEf
ScxVqgJYPQvbH88U+TEZ9BGuKuhXxbirhaDxX/9iHg7/jZx3DQlPzNBFhipuRj1L
TAkLeNk4H8EzBD3q7sTUUPqZUokwMiESrGBWEdoEoP+XPy0Ss1QNuVw/Coklwji+
ba9NZoLnSfyTcwO60nZAGnrNyPn4U0mGTqrMGhIXwl75p9KEO1St0XiBPmI3Q7eq
e6pGsq9arLe4BThwEuTt+nR4MyTRUtw0XZqZG05gXpRqDkGIVMyIqz+xVniHrLb3
Yzku5MZYr3/DYvkf02WQhNXoy0ab6iD3WBR/C1+t9kshOLpSnTbkBz8hEDqbrFvW
NqyIImX/b5gjWKvZBpQTvSrxb5VWcLbmLN+8wRclCYu0yc75/h8x7EfqUXpHSlzB
Gku24J5uggUNyMlAiCCjxARoiU035PaL/S5zh//SgFFXc38SdT1AioEP3mQ6/9wM
8ovypoSCrQVoQkGLey2/jeTM2LNPX5nXQu5fq4AmK0VGgsz5Qk449as5TjoA83Wr
0D7kJ2NPm7nWSpVuU+8mX+gmjJ7HSs+jNpMY7qWZaeda8j9JeQ480vQ7nI2W/UGv
tbyYPvXu2XtrPU0NaDQ7jfs1W0jOFp5s4Qx1SQ4o4M0cggIValuvhestmO+OTMcE
fUCGsQ/GLy3HjJIVG9FBu2fOVGUlQek0P8R3vgltog8gwIxGzFb0D4O5Czf6p7Ir
TMBcao1O+azjhqtPCEWPTXDi5CohYO5SXRA5l7LSX6djiHxw+LPd9ySXl/Y+lZTF
cq2R3kcRdy16nUr8LgfVp86sMnhu6o1b8uLAQtfHACOakNnnInhxfOEui2qo2XD8
vpgzynr9yj/ijfZIKyM2X/BCfbbjgvoeQxvsSUPf8Gw3vnGgwEil4/VOrs9Hz6ip
H54XyTcAfZMCwIuxLUUWQ5sYBni+5vDnV/dZrdRe/0G7tboawPqM/v+h5oAnELLn
Bb5oBh68EEvLufCuxJGzx4CuKOnCIaofRFyMoAZWhaF9/07Zqx+2Bl++LSilrhME
bcDMO06HAQY4RT+wUkMXBNfif5hsKPXFBacumwjJNbLClA3cEYmJTvfvRFTjxeUM
GddMArOpjkhANw3WpniaJfvi5YgpOIr5cEFkltmvPYF9T0Z2/P8Ve830xA9lnnhd
c1t/aDgNfv1tQHUNzJl2Aa6hQbQsW4hyQptTmy0Ngy0X3h/ogkYP7WttYFkSKpS+
Y7Xt2GkUYdvnW4nWwC4AogHG9zFjomRTItVAp//eLcq4j79jl7c2109HgQZvy+M6
GTD/0tZMXTW8q4nr5Tok3CXNnfVuR+e2Xs/u3jbYF1Bg05nTcX5vnjQ3CXfMwfhv
uxio1gzCKPQAXieTGp6IQaNlI3Pf3XgWDAEyipMzrAW2SqV0bllCvmmg5s9xYhM1
t8cCFpGQw5BELs/ejSpES7im7sO3CzWoZkZngOb2A2O63pVDRLJzig5JNQsdmyP5
4t+SWdsmguozJ0KrE99ZWWlypbZGESXgJ2KVjDOXICGTruC8gJ8rp4Kqz7vbJMrX
ot+Mmrm0JmU7QC8b8t1KgKMWr21RJg2R/k8fW53A7BBshidqq7fusApjfAtZltWm
POjSWz3IFmA54U0pLM3+Y+5xGdPw+alfU+9THoeBTDkv+DaY14S/njn9DlPkn1g1
qmiahL8yMBs8Ke4O/kpVwj4fib3r24noJJdopXovGvQx2ZTO4Et/YUxdImdxhZ7n
9qsUB5oO/3E4+tqW9g7p9jEPpdHW5cn2W2xdsHCxT6nWIj+j/NoQ1FUOp4OusBsv
qaZixmbtdkc+GmOHnhtCVVUUSA4qVFbGQGx8Hw9R5IdRzVSYZ8G3gl4xObuRTOBC
FVO2P9pOyCFsmGjdMluDvGWo3/vOIDSonWFUk29KWgTnOmUZ2ivVtyXkXQtmHwGf
ruShLm5VvzVXkxcEDdMdNjhK6WhlTUM+3UjX28Fd3UBtuPNDXh4gTqRQDCLTXGsw
ojt6+2NKhcm1LlSa2UJS1npE7w/AZEY27VEKlWX0pSXCVteIjxCIE1SwULTm6L55
NpfELda3hMZ5XVeXlAxpMmurpObqytnSxVgDQGSgSvceGuDNSyWH/I2oAmYd2++n
FqIWjfL5tYTl7T1t4LVMgDA3x1rVaD/aRdIxBMjALRzAQny8qnU42v+UAgQ5x7OC
JUd+bUmntogrXvZjjTqeGsKlqIuFHoIZeBKamp2pyAj7PwG2w0mYn+f5hCvnuzd0
tYaZXGA5/EocmkbjxRGLIxl9D5Vt/uK18xcSPWYSImGMs94ro/zxvXd5f7E95w38
N275I57ikOJ0zJhqbs1hWdv7cNcYVFJIi41/tOAD0+zXOtG0CUrHXur3Pp8jTjVU
1VWQVlEOSy+fVf937W2+eVDzzJ50MM4SWK8neo03StSuYOjcD8NHDCP4QY+0LiUt
NVgkourwQxrMYIRL4jwdC87iQl+ID+gL6yOhThlwE6yIxgIDe25Vd/B8H0zHkdn0
2nS2TWFLTtjMguvKIfSUCGTgPKrlwTjtK7o3hcbPPG9HGuLBwwdm4Oe4zqL3yQWy
jlspfJWm1qIyKf/wKt8AGxYHOGPAohvxiu9FWQMZsAQJkAknqrgsbimIk4BWcixz
RZSIUeXnneZcRg8i57n5YjQGCG6P/TrOljzL/drW+3oBtJDtRKCmHTs8woZl2VlF
t/kZe7dS4n7jrFhFfGIYnt9qxTJjc1ukW5KkShJMw8IEcnA0c2fLkYONg67w9tfz
q/3DDu4X0BzCuMSTAN81QDv+eF+fYZmkCLI4ZnLB6Mil3cptLdHI+SY/A9CaOIIY
cBPlTCN0gxOvGXg9o9osz5ZPfCfM5NUxnyNa1klr1OnxmFg6BOlJWBFcEoQXMqiV
VAr1ToKVPe8kN6bf1DSH7Y0dhXyiL7H041KE0vguHPasoY3CvVvEhHL6cI1Xem7f
WFub36JsDCTBGpH4vcdVeQztwYHevM/Gw3PWNpvFLbm6sAjIeGypxIP6rY8rqsmW
52JsQ7rb2jpWY7vGGPCh1oza5eIcBQHjrfCT28GK02PEBp40v9dV4g/ouBuzMnjN
aYeSuQSj3fFd0aRzgQOSWAQOle3XVgLWaFpQwRLVKuZgD4gYTX1XmSLORjBbVJb3
vEQNOLZpM/gbcGcxKnPQ5BehaWNhXABGms8Q/CINLvv2o/AY682KkTT9cFnMzyNR
CvKeg26GRL3vLjnqxNk/fm3zxzG1oJNzTdQ79UVpKZeTzG26Bd5rpoczPmghWoXM
qoFCYPNviGXWyZeRuBbhFPtjXvIB20M8RMSAN09yQNEMT4zCb/PdSXne5ylYD8fM
g3I7jp/soASWHt+1n0UMiAMk4ja+ZpNf0TzOLJllC+y54XKlYq30Vq2Y2DW0kWhQ
13KgXI6w7oeK5ZaR5ZqUxRgAe7VxKdFhENahE/KSAQ4MvWADKua1AKhQZKtjdYsb
oo64tuJyQPGyCSqOgaCL+optArMvLeg0USWkdbKDdkAi1zoBWg5CxjJIXxiYPJsn
Q4zLm1roAGFUbtBliM2NbmEVVlFb3EPu8c1bXhRKwmaYzRtVpfWVP/l6IyOr40LZ
SWnHjYv9O0Vyhzw0XYeizALKa7LdRPo3R1Wwza8j2xP1faps68bTZSR6EKKAq7+N
u/uNCQuKj2gxqLSEJEbY4pxivrL5xDl7azSXXQtI5iHvVlCGgfOzMr4Y+MS0oPVF
1nr6/au3zNgAudVgqOV6hUJp9CeRA3uNnuhweSvNG30BrRssNYB6q3GYQc/651g7
TWGk8OfS/4851o+kxL1+SmxBIfWcVLodm4m2CnhsRVsuNS8AxeTdtHT7p8HsBXYh
Tme/YcyXNJf1GP2J9adjZXIg2DnjMSyeJxRmjvelFKiuUKnn9POvKET5vRMU0uJA
E/MlUbSF2aweq8Df+11pD3GMCzNTcg3nFeCZ4p2y7gvphLBucc3zLi5Q6dIxcldQ
wq2Zn/t7EFnFVKqW/sgNu7ppgiBFyJLx00HGKuAq1ArEt0ue073IPgM1ku8VTLQZ
IL9eoyp5V95lczN8jk+TsLS+EPSEG4yUH1QIG2rOGNWXSdTshjcUHkUXS8SvsLB/
InscRzPdCOWtflTu16mnbuJv8+f9w38qcvlEwRRMVXyWhcgL0dNGOTW82OsLtsDM
JMYYBAr3x53QSzseESugAJhDoaqO8WIx11kByPajGcwSVLZmAwgiznYgGQgo+hwS
+2L7W8Zh6uh1eLXmKg/UU6uNDr0wKm+ceKl6/sUEcke3daCF3iqBHgJYPDcc8VU1
vq5N8ZG2Smu7toPQoe32HZ8XA6/Ym59bU+gubAXZ6W501snsc5iNwpTFEwt2pJQV
63h6ZP36RGOwsNJVGf/Qf10POMsru48p1DmCZOi3+3wp1m5pquFRJ5kvGBLV570S
0I9azTOnceCk2WU/B/QDXndr19Rd77eQGicqa+1EbUXZchEqRq02mYCAJHfoa42M
abd0pqXEMDFVmv2xDG9OzVN4EJkqatofOBWNLGAW6QyBsERLVnHyRaN11QrMSgOj
LZz8uONX1XZaQsI2U9xJuURs32o4RTn19Jeo5fE+ON4LrLM+cKTye5jgj+RPb2U7
oD+XottIaXfpPNkqxdE0mXk1pI9AHBD30+FjJfHLB/g7NFDV3RsjeIzlFZT/Dndk
nkEDGxnJqu3r9TDSDcTob2Q1P9OLoqsclRiHY2z91iwSeqteHrx8ToSRB8rCVTCd
iJcM09/u9YqPR2Bj0AAGFBDv26N9G0hvTWI58GIo6Xkah68NIZaAfwxgNbgJS3dJ
fkMt8MVDiGwJtooRowLQJeD20BEycEry4BXoxcS/7yVe1VFkAiBfKLt/I/f87iSp
AUTGaRS30KL6V0IqoeHaCoTOQcWEkGdUS7cHYZMPgzf/o8i4yJwa4VMqz+RAZPlu
EF0uBAU57/BBUZWznGuhIWF1OQNkIbpR5+2yGHAslZK04tzPU4hTpRb4WFhTzqD3
QV7mOgxljyT2DUtTeNTsXAZ9GBU+QJO4fp4EPhgIT+INVwHSaFr0zLQ6WxT+jeHB
YyZLYSm7tZ0G6EPL52cdPWKcvQC1sdAM7u0DX2z9E/xBUxQmDWfnPe0bxHFgdww1
fuINC/SATMnPCRCWxVesvuoxbfN3fKIbxmgY8U9QJiqyuxFnjQefdD40ZiSfHRLA
6iDrzSUEqPy4AUlpwwkrI4vFiyP9GRhZuEUPdKzQqfeSrTUu9IYMpCqJH99bVLtc
CC6AYjluUJa74v+r0uIRySGct3k2Uk6zDk53641m8Lumy+Akqjyuq4g4VBcPNy50
n6eXZVWtioGalFLUW6j/DUkRGwip7NDnxVdgQsdM0QVrXj9UyPKfNo3bmvJiylE0
RlX5UaX0Q/au/sF3pIoVOc2k3rfZwZ23yQxEkMmtQBPUopRMxKV5vbuw7SLEnUYq
bofILeYzE6Vg5Exkq7rTJFGesVelH6C6eMtTt6F0SwKbxPQQpR18mxveM1/BrP4J
ClEryLuFjwKkcnZYrS6VjHNrjVCv8THDgBnH3MELMND4ni2KglzYZoNq+vNCXwrB
wnw10ejhawcPV1FBuQn/4/sMgVTPF9rWOIh93WNyFJUnx9/h0GH6m4u3jPlblaxw
a0p6gOIqFM1jUX/9QO1d5lDwaocrFVYVlVpccVw4U69DAVgLoRB/L9NiDixLayGV
sXcMo2y3YfDTRLqU/KhjVeu9h1+xQwweSQ9lzWpHg4bjJ5V1DshGI3EgwacF6qoj
b/bkDCyCZUS3hij4EOcKu6Heyds2Z8r3XCKMnNDtCHzYVfuw6yT7AFxCDFOpWIqk
7HBzFI93px2qyWTEUg8Q/fY0vIUsTi2fQHA3PosO08/D4vbOHtbgNp5kk53sQYLG
PCC2OFEM+et5oa24avCwu/AzTturyLr8K9oWGLj9M8xt2ewk00Ew83bITfSigzcm
K0mvuPOuhxjVAwCZUiOvv76E9GMr6JIzpdxg5dtgO3L1+euBxL+zjU5R2neDSGYu
mlrMZZH3ns0BmOSwOJ4cMtCR6B3d4+MhwrKUtv/qIjBd/sh7cI1ezoNk0m8y9VoS
3AoTnAuChFNhUhFUKa60MRnQLhcw/h+UJH//6R6Li/MIbnvU6dqXwcg0tEWM+beg
ulE99QfODWb2vbCYLG0Jwu6w12Nsap+65QAW/3v+28Tiwjw1pygKli62W1b23Aeu
TgcTh5N4hJh1GAIe2l90QR8ssdhLCrdDQUz9d5SnTd532c/aXl3YiO45yTwJeG6a
DP1sumNhd6EecVFhu7c+B70f2Wf1k6WyjvSzOuAtYKBj7MnYQYN/t5B8eeVxBW5M
fhMGawptRLSUXIsbxwEFVTOyRytacBfDGQ4oRrtAQktqYxxFR7aTzmgB8i3mphW+
aiZ2osFhRrAfufcnStgINdfbTii5tqQiJUIZwLtznF33Epu8FPo4V3WaaDgX/KVr
vEVNmQ42pSogMYvbsiHaPAHGkNAcJ159Hfs+Hq4AskfT4//vpjHIlFPlQPDHuYOY
tu8fhdi9UGQlH+QWD/aygwrY4s+EpneJY2Z/UrdwizdzwFtshdZlZLhYeOcoFg0t
0Lv3AOiOf2u4Q/DVBRMnVaMDhNZzg2wVBKE7Irdpyxhecpk5SrosiLqa+9kkG26d
wvdGdXBrSge45/Rk25v5jYd/xHPt/o24NMnsrlXxaZpCcuZGX3SggIHfzQQEB4hU
QJ5+WF8v3GJjlC6zRW5LlCpZhJuCnZankcspQNjPTG9pZutTsEb7/VgHw1oVeSUM
SFdv3bKLUI8PuJZ1QFQ9kHJ5z9T4PawVx0bQ/g6p4Kz3/jnvV1Q7ez1+zYb9sRGk
6F33v7ksbubGVBH/+f0Jnyp5mhzLLkr2t80io0HBOru5PrUXRndlNNc17cHaE6HI
LDbk9THUL1oycEAS2Qustxx69gcjvqm6TkvWYGs8oDPKyQdkULGiGzNWTNMCKTDM
M8R6RaG7NW21bUoa0aBbraNNQfYGp2ATK/AwBSA4j+dTSczY/2ytkUWbSDM3mCyw
Zz2MNsgEOmZ+WmKPfPmE5xhtxhhj/Z2xaybY9/kRxCeXdRwtQS4qBfaVhKnf0bnD
iMaZTkRxrbEpoS0DRI74F0S5mRhzFRKNdXeihGbIKROw6w2zMivXLrwWLJmEPqDm
or7cx6z5/WgiMPVQARhdIwAR1gEAzO+QozKPirTc7qzIYWSNtAFRNh2tWhLwtToe
LB+6/Z+BKiHsQuQf0MlJyvWqxsAlTmuVJQbNrfoeSZhlcZw1mVhGkB7fXUymUhhN
repTpB2frFVGMR0Qu2cFSyLBy0eHknAP2n56mUT0kmApxgizCoCDqefT7yWTt/wR
Jdaq7r9Zfr0E5FK9vgKdXiFGmTYqOAJ7DpyWPOVd9PpoJnW2+6qaoRvH5CMjCNBx
pXtaR+1fyRo+LRt3uqUSU5xNLvHFDYvHNql+jrS9cCcAoZ6rTJD9Esea8tv/vJmU
g85ca4WUr60BQ9YYMwOWew5rFNplryGISzIQA7wS1o0BLXtE+oJy0zFS6QNCHd+C
pOvp3VQEo84lEZkzjuI9rKZltEexHl0lwdt/V1oSCjEkogHSwLUWvTj7BxR0WEUC
KSSjo7+P++HTXfxs5sVhX1AuWQFb58H0h84wik2MlqlVQz7um8/7JGwIF6TshypW
Z15DlanEMgwQ7Ru9iMsie8yxgGC8Rn8R7Cq/WpiF5YvY3BvBZ+W3bpg3iweSgPrB
/Hh4/aXCBuIKeDhPCHgxATESWlJP6xqfd0Uj2sciXwB+aEGDxUU5VFOw0v/K4y5q
J/5TSabRkTFp7Q8N0fnpKJll7SPgqJkL37iLYY9VXS7iYmtdy+GOBJlI/wC0Gy9t
uzYXl2UyYizTWtX42cv6wrJ5nXbP5kh3kGN3LIjdnhnNk1utufBMWy5Rog+CeiR0
lNXSG4DadcA7wKvNLgwpg7lqa62vgZK6Udlf+3RDy5h4gqy55bupz62MV0pzLOb/
C9ckbEdzZtQY1B7oZSFrJ24TDv0NSlkH3gGxEy5BLogU2LJy1OdpIgMjNmntIyds
f5dbey6yQzdsfNfS2N4UNmWrDQ1No1FuL18U5aiQrgpkqrxyJS6fT4cQw6WsyOZv
38RnIryPP3DUytV5JgkI886mygfSdQDZOxgGZzIFwuZTFlun1ZgboZ+QoIO5pqPZ
Zr/tYvtwTigXoloz99YPvePtSsIE/LoohWVfr8WbNcrjy8WWUfvNLaiPOfrCio3U
N3XH29NqrlMhsqsWKPEZ7S4VeYv8gHA/g1kol2nnAkfUIuDKaaeD2rh/r2FO/IV7
ZjsGkffKzA01LMtZcmrboAB4eTxocJOgHzJo0zuxkAvIgwJ9665j2jVuD7xUMdNM
8hWzP4DVZMd01Iw1ELS94Mkask69LASvU2PeuOphwPeEkpT0w/l9Vbo7pjgxAZP1
gF79R766LDB6fFk/yRf+B5Br8JUcH9emmK10YnZgfS8JC8OpUzoOi4joeKz1BuH8
jnPRi1GbZDZt2ypLq7fomFGAPeJbPIhFpQVs+Y50LyOtHEJwPipqi8szV7CRk7N4
Cd00qewVOp35uYlYdGursFcamvq9UlYanutg/Bhttf4l6AerZEy1WE4GIlKCoM74
1UREEhlJQIjFb0rSJ+YEM3Syl+lM3ehtNkTn9I4EFVuZjW5/4azfWhUhSbEX+o8z
nFVk1gecmvv35US4UWQCN0nB0bdWwWxT8eOvQdruFfDdj7L3x6BeSNOy3Y091MaR
j7+TcGJYHT9kFIeNmmYDDYBIWmlGddBJ+dVogTZzgTAoMXCRucVcObbLO1nLMcbQ
lCPh5c23DnXhaH/BnSS0xEeTKoS+1I8Uw6imXHaRZLqGe0/Y/O2LUXMkx2rnWheL
ZvIZAOK4CnMsHfS0WttVlyQujniH/lDLp5PBMuTxxX8dZMy0C9h4r1VR82UAuNlr
13BXFdw4CKM6NH1RTAUSYgeoRsyQoIGUycl5kasEiq28fNSHDcKV/yacK0q4Drkq
+pf41ylbO9QvCbmE8prwnFwbyhP8Z0hVN27Fj8PrYJEUWiBTc+ozfsYE9+sBuIKv
ZcYOurYTT1wYqFzlSX5Gf687WLPhFVrtzhzzF7jlzcQixLOi5GHWW5ssKmU8CU4r
/YKfG1Th/yaodCNlioxR1TgrhDDdIM3VW9ieURDoTmS+Anw5FnbRk7bJMvINpeNI
kFTnVMSjJnQEHPR/2zG1rHQoQvGlRRRbFuz8Dan5w7HCNbs5CuiBj23QeXgwT961
ZZTuSIb4HsKdwaLg18zJUkY03isj3MW7t2bRJ81PQULIyi5ZwIoQ6wiDFbcti5a+
axp6M5gHFEaFI0tQSvCCyGd6mA1tfGiwbaKgky+8o1Lj/gx7KqiPq7QeT8ctFNJo
Q9HT+lqJjVHNHgj84M0KB0Cobbhsm84Z7cpz3i1h8DW4HXyZCSiuT2W1WRCabTtg
FSLPC681Vd9XHRCUr8KiHMOHg5WksN4Pzm9nbeqDRgwQ7pES+DhZi6vp/eHScU5J
m8oyIG4axr31NPWkckJQWG8eDLmfJYRSdv5ETFkq1fIVYsGgVBOhV/0MpXljRPHq
vSn3B/78nYiKIG4TIKzQWSKL4DPXPQ+qGiAxn2SXwKXuC/txLBigQmWhLqaEi0FT
JGAU1ljH0xVaGCC6MA9jJLuxZ0qj0T0R7OfWJoy6j0UvEDmk7TmQET70tOzGw1F3
7mlIqFL9ouKIbAp9SIeCBHZYkJHv/R5WatzEfXoVweErSxyT5A7719Hm0htazzWl
kDybuE8h5qDHNrKO7eAqdEgcpA1JhP5WKVNQf3piUo8l0pKJW26+lW2ivEwrhAQG
8Ceq7mU+++JzGJHMhNQ7du6wVkFOgJEgbNVfUGTHwAD3ezPqfypMUP5TCB0AdEy1
th2LxFvf9ANZWrPwx1HxbACvmY5x7nTIaWuXat0xnQTbXjlQhvjuhIa1dGoPHjgd
CDvtGRmzznR6oavXgpjysxmwsknDknaGyNriCo6itgExJOj+0b4BJKNzC0TwZ1o5
gc/vsQER9TxJkc74QDAGSLKX1q8/WpdZ6JlTLYcGdSwuck+Iu2yDTjbxUVI+uU8a
uyqmtfIu8kTTDq1EyIU7pkXX49Tkl6LpLF1oYJqCKO5GDmsOEebmkhlPGaX5SMI1
A3Umr7+jnxH5R3RqQ+qMe4udHuOFG78wht75gtADil2ZjVfkeADWb1JEeVpq7voa
mMM6K78EqvLkXe28sGNZY7Ji0HqMsO6Qh/R0RYK1ITeUsDOG9qfxa1dZbqVwkkPs
uPDnEAqiFN1Qc3NfKnYqER/+LuNbe0G0fMqiYtfJCo8cHOpjCDHG3whnm1DZT7ON
vEWAj9L81dC1J0quyaUcccS3TEGPn+rvrVjRfUgSI/c41gGtnnow8ybpYm81v5wE
YVvl4vm5o0Mw+7GQY5xSx35uptaZbpRc0M98wsSNZfmVn/S/dhInQErfj/Hhk+3N
GoG8T64dM2cqqJefIEALK0hd8WlvCzTG1ItwVeWoblQeM4jTuP0vQiq/YXqxbnTC
WlX9UnvCQAAP68YLwBifnMfgtAv91Ui5T3f60NbPy/FIgUrRX0YlCF9RMGhJl0vS
Chcy6hYenX4PxFy6STxIwO+qb8tdUFnuf9ImhlRUL9pYK7hfkfbU2YQT+wtDOfSh
ggT2nqZK+2wFR9Lwu+kP9SQl/qr16ST9RYAQ8gw+FgEVYVPpvNU83f8QLHT5BuKP
e6pc0HdK3I+3iyY/2Q6UF7KS2VyWWyXNgwptpzJP9HGx/E1SZTYFFvLJ4/ZnZSVd
FGEvNzsPM/vX9hXOSJKajGCcWbiumbBNO/G1ppcSpCSelwDmSpW+1ZvNu2KiWdwt
9Gr+NHUlsYX7w0XnnTBhvDixa4L8eaDi74NaLZfrYOTs4WYSuPVwImhyddnTbMtJ
F5kAesv36OsK3wTmSsINLWpY0H6B7zc2jb8D7qwXYipN2cJPZkQJJDbNEehxs+WG
pGzvSNNhALR1SbFByyEz2HFhATsI0T1k3zW8ZXq5mjGRWUoHIqPr2BcG6Q9HXMQ0
VhcEloINla/RETF1Xr2vWGYqKTed2gMcMlNjDdcqz6SVTiNZdo0EpHoZTWy4w1Co
We20+M4z7PsOg8triIKr1to5aJ52v7HSIFFmd0NEbmA+uHjleouXRXee3RjDnzZ5
n2jfhZLVyGPkV1somZwOXpDY8g0Zp2l0ZGmPA6s+Cv67caazgwXAkpMa6uenMS2N
kRScSHDlRudlKYY0f8tITH8Eln45yX4BOUUcOFAclJueYGYzYQLHwmq5+08d4Ara
ITR5uytanrHIIOAvMthR+wj6RFlmhD5DktQ866JhVIPbA4+1LiFVU5ntMO38GLd3
Ygsb5setOs5ykvAm9WckEMXLbClXfAA9LndLzpIFygP1Vu8CA44ip5Dd1JbzUxab
bVwSEpPHM3hSthQSH+xavyJQItZTv0oL34z/whJMXIyIoHvXI1UY80GE+Q9eayjJ
oFQ+E584jguDx049WlGpWB/wASi7KX0JHbvy1L6myK5fF3EWpfnQ5N0P9kFdV1y0
9fdmZG+oU2gulUBlghA4flCdv1UrY5qq8hwjaecBeRebxSGzxT8YX7UkMUX76PYB
tiCoPJ9Yp3oCu46UIYMc55K7a3Z7nTe1LemsC1+KxX4YSajU/Qt3ijzI0zYWnh71
1hWIDHYasvHhafeJ6+BvGiUadHiyFvy5b7cNNHHth2WhtLpUwea+KIfaxBW7xRlr
NXKhvEk7WjkSWV+YJfO2/o0dOGHqUbgAA+GpuqchhvG9gdxtgt6m/7mJK4BnYhk0
lS5H6oIUcojOEKW8v1f6okqgkrTkT0/MZuPMu738kiiQ8totalTtgOoMGVP4X8BY
YS4GW3onKinYhlJIgH+RyOXujqMXHGsGCIFA6U+7BmG/qCLrNipPLTv9Jqfrbgze
wFEylEC4F/5vmMoonjJVpPDECdPLxFh11AbcchrMe085glyyZAmzrXUY0sjc41sN
HIlqWKX5dNBMN2jySopdC4hlrffK8IRARDtio5uPY1LdF2ttZ/JUZjpCF24OleSc
yH3iR3ZxbI/zGXEZKxSU1NohbUFvYTqxmmtJaz0F1VPN/4WV5Oe5jARgTgZFjNeR
t6xp2Cg8cwggZxdKy/8nna3Lz9JTfI9wFUQyJkxuFichLkfjeKsdFoFRdVC9AZgn
zuq/sBIDNDrx6EphKoN+aTx7MskGVD8I1ITeVg0Y7fEub6gOAr5tBJrCNujkdWmr
ZXZcXzPuWphh5FrDlU69rEzZlEN2qtcqOl9ylHI3I9Rv206PZ/lolf2AQgbXFVx3
o8RqDTBXnKLwVEAsR8Enxt/lzgOxNSRrDjBNumzkJdCaAulzro2tKynpjqyneHaV
Fluw/ccToDa+lH5nbzI9KHXeG0t/2X0h5K1fNENiO0YrdfvxoejtJ86Z6pBVlw6W
ZnKblT+9D0ke15RHikOHht4oENkZBVQLbFXqbZVAGuXm6IJt2PvkshDd/jWCXe6N
RIkVeQ/KsdA9E9kc1vgMTXUwSJXLy+NDud+ryPa1sNsE/PwqFK89+GQZ8gzYzVZU
IHmv91bkO6Wt1oXrnQRHCzHkT5iFrnm4wq4Uu+WR3VWAwQf/gTEs6x259e5mk2w+
E6UiApccjuY31s5M+Dr7XpjGytgE0PNfgrfLntmLFZpscROi9hyPVfNFrcjjvOqm
6tuAzFrFv0CJjr+YEb+ryOxDZ8Z5+wlqjx2ajLT1guapPfQqRJwm+rPbU684OfLq
Ro7/5zxIoeqo/LSokt4TF+yB4THD78F/VVxy3XwKjkZq+MfE/9wTVcoRhbG/hnTL
4hpP09X1i1ofolBlcDpzsFER7Fs+4glIi4lwL2MZ959RAcMH5xyDf5JMEsZErBZf
Hcp3iXgNP+61D5VKa2fbHrzyiOenWN3hr/lYUwNmwjAlspyeIz0EVb+Jufjjvsn7
w5i26eX90JGzazi/HvEMyCfRYXoPGupi6qjwUEmY9zKAo/cFsQfVb9BlSH4PAiYZ
uVmI7j11dv0Q7Wu1LVt7sreUHWZX2NcIP2X6rBgIidsd6cc+ClZSj9H1Cag/QpbW
SmEdhKXryg/ruDsjkEZ41pXyk93tuBZawC7wQlbTpua71ibdmGQaSENqxS9Ci1E1
Qt3ygV7mMn7UaH9GJnIdJCTQxrJiojM1CEsW3s1TjpMu/FFzXQAVwjEL7X9yePGJ
b+7rEhiMKc6QRvmsmWiEcXMwB3Ynz7pkCHGj8XtAsuamkmfDn5lgBX5H2iogIr5c
pCkCAfpa29813IMJDz7tzLOBP167X+9gyWVoB/6jnv22yy5Nf4KkOEI0leSWamh4
r2ucnEoVNGRfqjIbssykO6nkddBa+/qKffEhmf/KNK+MSVzXKA9XAj2z+ffOZ0R/
feqzy4yOFsVNFuXIJPvIgt0jQQMbqg4w1NEbjybr0SQGAFoU0RveTdh3WJ1AfkZc
KkaTRfjmLu+ez1p5+HzqxX358azn37sWBD8zIGCs39+gsPX9p5tHczd9RvmFBsSD
m6IhBhViuXRn3SF7Md2afxe/WNNUf117vZfx9RCVUvChir1zrbpCmBCDrHD45eW7
zoRK/5cRdmhMdPGg1INVoTmwRXzfJAZpChNwHLen7WuXdNgkuwC3XsC+VXKsv1Jq
/cbVqwZjb/nvFOJP1Vo8jP8ejElzBuyhUbGsnUfPJFgeuxZZKewulslQ7SEF+uMc
x49+cAO//Sg1PMRhNM1wUgRmq+eOVFVlRKK/fM7t+xvuIwMa1Zas+v3/CdOeFbDg
UoEn59qfT0pqbkCzViwe25PZ03yWWPH66oLrMuzMWc2hP/5Z5/6OCWEYMpXg6n2f
EUedaheUlXSXNqlAR7jalYL1silQ5PudMGg6XFBKAyLAS62IzNsqEEw88zmmTSq2
QmswJYE07nFj7X7eL5XGwYkJj+k+uMix/hQelOLTHQ48uWwaGtk939cwu3mfeMwG
i0rAYsHXKyO2sRogUEVCObwN3F8VUn82a+2P+OpJxyk2wY0ZgtI53oQ0zN8md1RV
tBNvIy7qdHsjh2XnMiiRDacPOVAFKUhaHQW1rBRbpULm3J8FLdO17XRD8pbpNoVT
K4iMBGyhV1+kBi15OrAf3OQnbv9BDn3trWL8nS2a96G61QOc7HpNzD7ZpziiU0L7
Vh4q6+k88XQRvh9jXqWhjWVjwhs+LO6mhOOzDt5ilvJUORFiQv7uI8ONTOwyywr3
efJz+1mEBndpWCKP3WzyNXX9AHPO/ax4CK0xk8Bm4e0g8tADU1hlOjOOP8ys9KBx
fdU01icyy5THmP/RjRNT6cnr1K1gYmXRAZyzGb7/j5q7enTXIg8vBYcpMcL43oX2
WGt549owIUagiMI/LfAmd/p900SFdCwIkXPK2gAuIXRK21pl0L8RRacEFmRRS6zi
31sNWwJRIDrB/k+eDhPDl2XYutzFjczdYCjk/C2wsWbqKOw+z05J6O7Tp4IIFAnJ
h6O1Nxqnv7wdN/mHKKWUVGeZEn/v4x2JcIwB9KYhMTIHqG6axGaFZBcIbe+PyDyk
vpMQw4GsiHaBB4CGnMv+AIMAJD/9YIPq5DZAUbJzXzXeeJfCrk4RDV6OfmFwuH+L
lOmvKpVeLSCRCuvJbih3IOzKY4LYXjy64vZmkx/ZSSDzChStI0rp+u7Y2hi8oZI+
nbIB0YwcSDcLV+4IDw2s9DX6FFxKCZrlFKQi+DgrHLmWWH/mIsVt1LUsxMVsmuh7
FVWHRLqvCtryEV8BK9CMG6xCzPoouQdLwYlsJ4j2g4D2Xam3FN90cOd1kGRUejyu
k8BwCGts6saegciciDYqgHvI5JDzHstbfbfnYMADIg098tExD8Ea4cOAp3Kfu5tq
sINQCxYE7f9I7mb0GwXaVTRtwqzwrc2c+3xxAHVL66i35GfzdpIyUsVx5wj3FWPB
NRCcXUqIUA35wKZTvH3LTBq1z5WR/EVKDlZZVUWBzh7VDYtVdejgCycDjtLy8ISX
7x3NpgAimbiqddK8ZE2qVwOI3fIjFR1nLlmdW8dXiDhQc1UTDirliwJRxYn43B21
dUe5lm32j4309v+HdtLjayGql1L1y4Wv/LbEnILChXIWTZ3wBkT/g4/qnKusIamd
DOwfZyGyuwD7JcSBcDKpWguM+9fQGv2wau1cgx16FnPVwybv2Pq2DEfrXAM5kudC
eTzgREOXBLjfw51UGVz1/fHma3fKkM+Apd4KAOBQIwZA5WhFTzUsWozNSy7KyYHc
wGYag0PwNfcLKMQwIAyeFtqjhBbPKS7uk3j/Vc2fWPzb1C7t0t1LtLeYOGjTKONm
WUXW4ywomIfkl9lUqAwoV1iCmghC6AXoDVA9FBft/Kfl3+HqmkKINh3rfM81iBVr
WXy0swTxMg02A6UPASjp+iRAgkj8O5TMh/g+FyDnRD4jc19AJ0Wnoii9CO/syTU2
zA18AGNUTHVyFt65Ji10RzpZHHQ0fxxHjR5IuTdFAc35uTzoz9IE2NHX+OpjMk5y
tbfvQNbGJYozjfIu/5QGsWBYFlSUbxJ1IK8eOnnjP/K4vmdYpFSWkKNAVb26LLDy
hdIJhOJajGRH4xjOJisN+0f+M4R+18NsXW1sGe+lXikfDW7CWRfTvVfKVpHprkzJ
zdCe6x7RkhFdNcRK8ZTvyaTAJo1XEg9Jq4j9gx8233+NASP0jIsA8bgSvLIvzKOU
gPymtaPI8qH+YxHRzVr/V1P+ueFUcE2eIH8yXaPh7vvHAmpi4NGD8AYFIT+H0V9H
q1diOrwh9NkJ66UYiYn8cHusCBy7dhINGLjB+HLPEuA/cOTPRY+lQVxz9YckwJz+
mnpr+As0+9EfSaFmPoPNKjdfv6FTZVrwSmMDPVRo4aIKh5ime3V96zMZK0J3XIif
YCwK2BN5DP3MDh74yRh47MNa1naMKswigpkbclhudMZ7Ac6tABti5gag62Ir1S4Q
8Iqq8jylHzPbJK0P5fWHEGp3H/lnsCTr/fTSrvCGkolbHan/GWMYs8oAz2RIZh/W
VJIBHhB/beATmCBNY3SAlXOpMvDuKb3T5fMdviXX7JcIBnxzTdhmxX5+p+R+ljBa
UJzJvpL3Admflm4oIf+c5Y9o7V6FB96RYFV7NTRwNw4bWHzYBCM4pLh+tjZnpB2Z
PPPu9d6EdlgKU5tI2kjffVfz1T3oNDCVAxZRfT+VoQF878rhtzFSq0i3EZ3IPbTw
UkuNeWxR1qPWJLwkctEKnf2Ze5t+bNNq+RguT19W5KKoQUE1aexPgRyTLRctK5he
iZNQdKrQt4UzcfkHCBY5VF12Qp9ERmseqKl1qjchjeVri9Ocyr12dT8LqrpcVDyo
8UuRzQOK26rULRkl09OGsrAnvQvwVV/e5iFlHvJ4Y96mYgk+1tSUIGB6qRW+Bkny
58jHoWoxRp/2d9PIQO+NfjFFyMlv5QIEvWHjTKlSH9Pbb4sYkj0ammP/iBNfXNuU
ZKtU+80lT7lRKKcP0H6hNTKWWKfExdm4tMOd0QxDuIAwHT3c+NrkhEoV++C3TuMx
IxkE/+PeoKCFI0bbPdiCx8YgVrQ17yit/8Z7N2CS0BWCQpAUes7RKoEfV7XgQhCl
BMDZseXcBwPTma88n/TtBybJoLHuOBZRftgmYHuzKw3MA14uD88Hh6xIfaRgisDQ
km9VxEY/wJ/oVhIVXoxzqLGLUISQoEAfQoB4bZbZL3ylYgLJZOCECpi/F82VCdkm
66qCNEIkphlmZtHUKahH4/3XeEEZQCgEU11bdqMFL1Twpanwta4fflHiad2nn2MQ
OxOY04ynfhn0YHtmw6fqWMM2yb1yItNUvJxjI6NBCTV90Z5+GfnxD8B06aP1/Jmm
HfMQVEBGlbZI8RYcpUyWgVFM9ldXg+gJyanjLOlje8FhOXCqFoWImJqmrT8CYRIh
4yUmtTdd5RAN/Re1YWQe7KZnKsJWeXtVcvykIm8P7gc+BAxXu2kIB5MvYJjAxr5a
G5Ds2oM6b7Uxasq964XLMXJnc5WufV7tZITRr5WXqjjPXLoBcdJytUoAxY4mcHsK
Mk7voCkpbQdDD/wPvPlgYoLAfigLnI2HaAd2FcZXrqsc6EXPvoLDox/tYv2A6zX7
7ZaleP69uXcAt9BSXzeW5/TI8rJ7pMXndyJ8y6RpaZS7sn/QzPjMrCd5K7iXJ+xx
oYqAhZdImH/khH7pYt0kwrc0XKCMSKMDu+T79Sqai5h28YcQ1V4UYsIa3SfoCqR8
fO/sTyET23VVeeHKmEeVeAfl+625cEVovHzwQqvM3yOoWLEMicDyF9JvaYpAHaUY
0Kk+5CHpZCbP3BkO4jDwrRplWRrDQXMpPfstpxd6h+OSO2RA+ZiFU+Z+1FizRkXi
MUJF1DJUtfhw9mRkdcyBYJDAPjMndfNW8Fpy/sAy0+nJZOj4foLblWOnB8PrCv+q
ckCVqjOE/k0i1RXNQLotn4sLaq1j8uL19c+L8S6fyYL/8G3Jt/3vjZB3KIT3Dw3X
Gs7znSm3DfybsdKzB2ruAIBN49SHfPjUK+d9E2gfCD+RgpER74Ce46xk87Yf9/pE
AGqEpqGyCfZrYI0xEIjO9hkWtuCfBzq/VTypo/aKlaNvlfpjeORrtfQR4R3zJumR
KIbOfozd5o0S8bWoq9USgtVFMKlTD+W8Y1mEJke14y593aq/Ok3O0uv2L5nLRRyC
0YwZQxQ+X4qTzFmqr5oVwghuc9qXe902d04HV2BonruiaUjRTXEQqr+mOzQFg9Ht
Q3X8HMk5oSXpBJ1ddhibjw0mNQMtPAb2XznRVYvKp5UkfH72ULxzxxBvy+MMPOFx
XxY+EOw/CNViBoBeJNKANJrM/q/Cqcxr4eXtwKP6JmaAOvsTHMKZBnooMPAxW4pw
0c2X2xzZJuUmZMSlrG6wqXhV5sgjIpTNVNZJKWPFMbXAqW8Q2tILactApzDRjtXz
NqXB6WNOTdHZgda5tb9rzpothu7bhsAQBoUfyghVGzMfgrGIOBdscseC0N2/2Wrr
9xSvkQiZRcluVVfoDOYAczRXFNpPF68OoMx+NmPNg3XoXDKRr+hBoRA3hDwOea1I
7TJxWuyTFco77vmqCgpFkv873nwp/FdZ8ILNbDNFt5C4lK/7CksT2rqXnSkh6ton
L5ThY44mylCkv1D3PdOLvPQ8LF9skosL5V/A6CkJsmap++V5KNVgfya44wP8AAxr
K+yFQ6TgH2bFp0JGkUa/vXG9M7gXbLT6Hrm6W/eWHq8pTSqhNU7OJklNzWdpwJlU
GBDqTTDd1iSw6bBLzy12wO61sQHRU+xc+3JUyFVtlceDvcnOaY+7qjvxoiVOTnIO
SDWzOkDWkMvBt2r966NCJ52aCwlvCWi9JVtbZkd1MwL2hRPVg/0rmXEvOCBR6ui0
zCzt/YKyOrWGRIs8RRFJEJbGtwXTqCchV3vxsZy7yGE88xmZLSewYetmuILkGslK
ePkaKr084yKQUpuVd3926vsGbKrPupdS0WKGB219RsWx7lU3dBErYL/STFaqCWGT
WuE+vwBg8bCRXT3BmoUOM6VyVKQBn/QLqqIWtIT9JFLKHWSBJuP743jvblo8ZVLO
/hKVoYrI4hipLrDec1XeMGpUqOcXUMTP3Q/8LpWvDQbltTXGqbYCBzenW/FFY7Gx
5+1d4suwLVn1bedlBEA9VjYAiR1PgePnHAJYUlGY/o7zVs7dYgrHSAJ0/jcZQYIw
x2kVHFFyhPk7ykd6vRdVhfLbsWhTpjLwwk0Fc7GRvDIHSrmcS/eE+POwWe7XERBn
lK/OJSma244tFd2xxTt92s/z6upvDC07+DXhVOddpT3euMfOl8URTRVcusx4SSxL
gbPyZ/BEY7lW3jRK3AGZvakg8gGWD8OhEiAObSZnXEoNX6FrJsZF+mqpSlJeIHlj
04NhjFdGDbZv0fTfqqd9BTMQ1yJ9CX0sMb6P1XOZlupq4DQKyDFnCty75iKuBHuw
Vqp0flCEkaB23myPkwm9RdvQYeLP9XG+js9+u/cJP2ugZGLVcWC1y14UCSNja41z
HjASRoxa0S1mL9aKK9jXqMRPUINsDxzHPdcFoIWjizoOGOLh9qazuqE368fw2j7v
iqEc+6Afuhp/mr7MN7JkNn72p+MWqJZ3FYlkJAp6IGwkFyA9YMWS4My7JpW9eH3U
qTpatCPIIfA/BSAwI1O7skITijJoJoZznrxCDIUW6zH4VnTH9ZqZXLObHHvz4TOL
n0in0+jxIkBzoa2Zf79YneiDgDA0vhH21s3EwQyqQyOawwR8ydL5J1nOrtEotfwe
WNfxQivYvrGnIIh10IqIU/RPT0+pc7i9hiRr8TmXhHPz0diAwdZIuLEHq+78rvfb
P/BKCm5AJUwCdUDDVm4vHo5VJCrFuvPNKjlHi2Lij6eUrTPniysM1l9Krqcozwwr
WYut16V7xOO4WWFc8hGRuHGf/unbmJKze2cAOo/RO6CViIJ5+2fY8laMOuCifXQT
dX/g9O6rNd6RBs2bBpt/R/9MwU2xXyUL4GagV1Jum+J4LtCToHyu7byGD5XFhcIB
1A3TcaD5jpPBuRZz+OuupN6N3YiBUNadzyia31jWKyrT3MkJyQ+WGJScjI+gPz/z
nssVuB2pAGltCbhoCc4arLWoZUZTq5uMX6cZzTNojKgxSuoON7SkKIMLvF3h4KrJ
OjVUwIip77PZWtHV5kZ+JV+uRyAhZ03YS+t1xit4g7Ag0HIS3tLblbTv8wERllez
6O37fIIi4IdtnbTpM/lovaDV8OB6KIA/WJ5gkPT1nyxoShE3ZrvoAR3v1vIMMU7l
lqJvE5H0hiTaG7fwNzWyUhWFirWAjT74tfVYvxsoMvGSkLvfAUtHWYFIqssDLx4O
hY5elKZOxUj8zDAtr5Y9K/79E+wy+m5InxYKyrxDYFyVaP6VGE4at/sbrheFAFri
8y088z1zEqPkVGGzOcfKLia8nFkHnhZWZc2ZIWu15EYgKOlyxhfAUKRzP0UbmSqJ
LTuDp9mY8M6DDIHceUUeuU7xTy95dvXZhbP/qRVmfqADwEirTxIkZyY2xGHdot+U
jqIs2BuoaEcu2GDkMFVUnoWtkEYuCQgruLhW9On9uBVzhQIZp/yuXTzthi5OxF74
sI3nzbCeHMonoaKZLX/ORQRVQ2FpBPK6pZ/56Ax1vwm/Gk1Db7Aj0vf/UreBr6VS
/gdgZHkRXNPkT1j4woiMsk9SjhIxoiIeRML+n5a8NoT0JIFZpFKdCUm5Pk2Jpk3q
z7eFRkdW3L1L0TGc8vSK7+2v71T6Wd8sRcFUWGUJOyhWuHmlZNAUBG3+GcOojl65
f9HUGjdMUOJsGDz1Vtqf7/DpoJ9myNy0/42fDpiUkmrOjm24xnOHcSGiH9fCsX3R
KQwVhazdRfc16c+MOcfaZUnPcQFfsGd0FgGdOUwbjXZjv57nLc1wFhM19QaC8Ial
KMEt5a2ptnaG8OnlbqkMPlSqjiX009t4WJoufN0bCQVmFhSol+XFG9BY+5owE2+t
8hU7TEOc4/Zx0cNL0KbPSlA5EW+qiLVhuz+YS3cYg9SO+x9sgtch66OPev3J0fh8
KUx+9Z/gNYSWAPHFxWZ3XWhB/M4X9kN/oTIBIINJlJAIDm/BGJgS39Q6o5GZ4qtp
lOqGtmrVCO2znSa7OGlZFNF5NJ6caMS4KKrrWtn2wvQkIYSYEP19eCOjAYuihr3Q
lVtxEzUEwIbjzAYiwPEoxRVnix2xUGuVS+uj1NswFxqf+1vzKx24gW0hbOCvDRtS
A3tlkfP5jD6/+8jmVas3Wor8FYV0XBuqB5FUpRrWRp76waoKbht1/GsjcdLgtU+1
2wcavkVLl6AglCd0Fy6qHTbgES/nMMUQW+IkjVFIXS/3iSxQkH/lFivrDHc4cCWM
h5CbB+dLd07ifkZfek4FnzppMibMceUb860venPWLRcIB1sUSLzSlRUFAtnfd9C8
Iq5nNjlM6FUfORMPW1ufqaRLy9M1SfnXNsmtZCBAb1456uk5WNZVdDOFZJVn0fG+
9yTURP8OcLwpAD/EbdUBmg7KolMwm/McAy4WDpVRX+pJ3LoyNfXX9UbfJ0KjmdkK
LBejyl1gkhNQaqBnKTztDhGdUyj66b5xnT9z2GcrAfQkd6nOV2fw2A1xR4ffej0z
I+6npI0+7z72QIhFxCzUOEe8vLOWP5S6n4KvHVfibHPnOWicKZWcrtZto2gX4fGa
KBauPNziBScz9UXGhqWuV/zx8qxguL2TuBcmcdCdxX+FmhvrWG/h3sVJEoiM4HjY
6RF0xDlt8aWWReOY2zXzovjS/E2wtE/v4WxC8LBWe8ZgB+NAmN4ilbYCfE9pjnbx
OzPAougrJP+mo8170P5KTo9l0yNwDakRSJDWAEgOPkXFGwszdcQ4Ex29zzvE/0PV
x6JCMVsRpD6bGOeyLPdYnNjMciRv1VrrpQwQ62dLrOE0fw1rQCVP0/DWQvBig1ij
yWaHMRYXw+Fthrwt+ZGpOkv5rifDhxQwdM5QUhJ8jUDSPiaEUdOry/vXB5bAKZbV
Is1TrjTQ/60r8PMqlv29T3Rkao3npdH5PiwHMu4iqlGISWZ2/8eVQEBBmPv97+t7
yhiexmrMsRIvXahs0UKLMgcojqONGkZgktdv/wBLCbD84w+9q6QifQ2ml5DLcy6i
sHDuC1aCUqR2AJRy0mPCtVhOapue2z0UK2+KCbVFLUTpspC1w1H35uZcc+JxhcUV
jKp/SZ0buTmw4+48uwwd5aUxs1scpBMOp1KKD1Gfl6sZZ1RZ2LhkZ1ax6Ag9qC4w
wYt4e0NmupHw1aUjU8IMQqFLN9iLmebmtsyogmbC91P1KIccEqyTfgdX0piVAaaf
IDhZ6qLhAS5mjuHVizHZAAH66pJdFGQQHNpGApYkUTWwvtV0uBwWI9uBptHkn/L3
+lQ2/stwNN/OaKcwSNVOVBdqFItHU7RBehESVGGaVqXve+AwTe6dIGGPzpFR/HJw
RqQ1ZFXg/IPp/PhPR5LWjGlJFDp+83kHP/OgXnTDjj1EuumO85Zz6BgoDDTSOl4H
6be+VKn8ffAZW2S/tCqBY7pAg8BtqNtFJI9qm21G96VylsPsEJfTTYHYHjbjoXg0
tJNWnrF+qjMMwAc+kt/UuRw+H+R10yZAG6Ri6uKQSzIrtpYStER8cqKPCIfHoZKA
yUbDM05NMyw6WpsgMp55Y5HcCIAIfnProEoBSRhhJAol1fyzpNYtEiseREtYq8zP
WI9P279CK7D6vBer78oWGZr/BAaMRZhyEne3Uztrk7vT2ECZv277TsGgm6jetAGN
9+oLGxFD110fMb1BquX3+S1X2T3ZkRRDFsPRPPEqlZGmTyK4olIsEsRj1NxqDnXX
hjP3E7M+qzFa4BfvuhzoaTnjbF9hBACZArS9rlwoYrEmf1JVjt+dMViQX6Kfcxax
DhhcHpNXShk0Byn7VQKyitXvBjmM0VDBuJw4SOxrGgXyzqrPWmYmmqugbCH+/QyM
arU6ux73rBbp8hQiwt5YXRkRYTcYuuEnB4t+8K2QIuVMvZiDymofJdoEyD1U4TeH
mIG2mRpret8AYMvbSbApbV3Ii649VaaLcmL0au5hlyN/VABUpgcV/GB0gmIAfbHG
aB2aePIHBQuJRe72VWoky+yKGPBmCd/2yoWdzgLKKVNU7tP6XPs4O4SdR322WILY
IuXMZXARwbgqVc2kvy14oL65Ky+2CX3l7XXjse6Dg5FtCebtJa8cb+DPkFnxvu3b
+rSRxljbWBnSPWrAQgCorFF4XEHp8OuBtBq1/aWyHYeXW6Y9QVNjtuzxQTcc6Lep
6fTf/Npfps7m7L7zWetshrF5zFJpZ3t3TtwSkA+NOB/ydFk41DMzx6VDoMAnLdL2
J3CZOeeJWQJkC2Ks1sXTpn68G4jsfMCDAwggol9B4cpzFvT/ZP+bT8WI1Y98VeS3
gT7KjI4tt0YzmV5v7JOwohCjq4SELoMoJQ/sGLiKZ8rW+EoGe587h1Wyo/f0OJy9
Ec0q7OHO1I72193LY4XJCbqtGAbw6OWZXGAUerYk2UgsJeNCx/UGoc0DAzSFHjaC
x5qGMYnq2zg2m9hXXemnOuc6h4jZTNEkkFKGdHsQZvoF1+6+5DRjz9C3BrS8ACHT
WsGjFhKb/2RuCY5HWolvRLNXn/wRs8ZuzgSTNzEt6n+m+JIhGI4ckSr1OAYNawHR
xuw1Mw1tHx3XtEezM+Z2O7tIIhJPA1053xuA+H5du5CjEyrTI1RIoUGu7HGBBSVI
kbxh1S9oTPE9iti5i2ch60fyEHQVX9qGOBOmhIuPGT/AA3X7C/q9oEru62NAvU62
pqrrAzC7pwlHa24x0lxVyNV659+XmDjWr+ntNsr1roBW1iqOq+ONoMBIWwDF0Dow
cd0X+UDsCBVA7qaO7y1eDIm9fadq+WfgxoEXVI4ZNkDkmH9iab44p6dNQl32iKPv
G3Q8g9N+jNvfWaEaJRmZxqWVG9gDMc9tY5bNujYdJapvhaI/4dTOP1/MSJBTbx3Z
rjPs28w/YRpMHoE/4wQStGLNwwCXKUdmAzPuVm2Apyc5l0S0iLuSOAcsqTF+gBrf
3x3lKhLzVCAoSODZwdVNICI53i18imh7KBZZ9Xd3usXRcpPRQMVU4tF+R3EbQqcu
Sk8BuenkewyiLUVgDlzwJfTPxPePGfgP8vR2/aICAzaSehbHMZqXrAxzkL8VEkO5
pnmcsyHnxRDOp7WQHpLymmBC1WElV6LeHkfZvbIgeW+BmcrMP86OLx6S/Ch3qSnf
/73CdMzlQZK9HtT9uCMWEsnt3YHrYntpMS/IKL4JuadEVyJlTmxqgYpfOWks5JGW
jOwTVbRL0TkoLBXiSdWusFRrwaU03FwtmSF+HnyCkoMyOllIUNxXWBQfKQ57K3lC
OJM9lpGeGkwXItD/rkOEpPXSR1Pr6XlZtT4V0zMMLoK0e4/fLoeTk6z+7g8iQyRy
+bWyaCmafYR/IL9f8dCfICETIuaEZC/RI6JdZk3zavXqgXtbFuCdsRpc4rCPRSTC
kvli/Qdq5n2NmTGEay36hW/bdHRWMsFI3eLRYI0/ombIyh6DZKfjA+DV4OIcO0kO
bqHN0aBDx1h92BpFa7FmPPQ+nNvmaBKwgTGOKq8bVJ6hwmUfVaHPzd35haiCe5C5
N1TaSwInr9crcAgtqWCdiyklRpy8OtVES1wD5z4dDAgoy+Lp1gFN9UlCqHGmLHoO
JTFMk1pCEfa0splTSwgkuXfOjdDYFBSW+fNVdksnociiRnv06xdKMtx0MAyrAJR4
FiVcuSwKR5VJmQ2RyGDyB+Jb/D84ghW841a0HfQGSE6jql+BHMY7u60ann0RPMPI
1klhlyFUUBWFUJr7ajf5wFadvL9amhyaWDF+GWd/iC/P2c40JzdrPq9d3iqWJEYd
czF0JrNvgkHtjEf+TxGSMrV7/ly6OwpnWBHgj3/HE+OIHbbMk56OOpN7y2vixChe
BFPYh0PF2vunh6EpEAfx4Tzt6/4LOTDKg5lAtIhp25aF9ImH5LXAqhuEWenYjiUa
bG2y/qxuAJzdClI0tXGHckhfjlJdGyEJOq+hueeR+5nlXMBqB9nVd28thtpVRY3H
F+mYrGpezl/4Rf8p75mO8DqO1oPpTCWipTzpgay7GoWoMCe0QuwNciO7RL0yaZyk
aVM6TEOwZ7Sq6GjfO9+ox3myculTRgrLFKE3+ch7RF0SSwyXuS7Qboydi36W4HO+
klzWeiFLNQWuB0RC9o1eVUSVFFOYlFoufrC7tEd0uO0iHVknK0ytMCZmXrs3uJjm
3Wv9oEH6ewRR5uoKHhxKDzoTmbntzjHe4n2n9JIocRNKUW2sySfmbxTk+9wB5Otm
VYj44/D8vP+MqSDtFmbExI2olhk7+Y/GxW4FiAXchmqnzh9u9Xo1y5N7LGvKjtql
ohCOGMoYHt/DDIFx4Lub2PsCXJrXmyuGKNm5z+ORzuwliUpnpAzWh7qt0ggh0evS
Kth3SR0szzzuTFEibODgy34qf0NjA1Uaq5RWgzIEVptY3fHulHrCWqnxh4tmp+pH
h1eEhDNJjUpsh/lUfGourBZXC8rgNnfCXEyMgq/lEuvJTNASSwzEVUTq6gaJ8XxC
062jIIeBzRTfuyrd4m9z+/Unbpq4F0kD9LjKrh034fbNvCMGKDWX9BTJle6ZJgm3
dunobHIzFctIZ5U7GVhOyMYdDBqtk452j0aE+agE59MjAh1SvO1Mf9i4hEV32IRQ
mj66rAXgSO3MnH1b7+oSV8HuseblDLWn9Oye4AkfcBiLsKvsZYvwwF9kkiOwOzu6
AXoC31HatvM28CsVBRclQX4xZDFKkrkjU6H2WlG+XxK3YcJlAkVH1X9buancEwtF
GkfxgW7Huh3jSFQftXkfV8p4+kWC5UCLQqsG6JwyX3LXz9twqQEhFSl0/FxYDfyG
dlhrFL6Z9N4BrcJS9nK2i3pYYSbwNHOsCxAO1/gs/cEJFEKnmvCIKIxpNtaLIXiK
3AekGJ8Wk9CPjPcDUaY4Q1SiTlZadNW4LSsr92I5OhyLE/3eMxyVaoSij3GeSJTV
HGrygcnUpli+vbt1vt3XCGNthmd+p/UdXI/+C0XBAxqXCSDc/NQS60LAKrVDzXIK
SFFH9+OGkmDrDlaH/XrRVO7bx3pRz29hQqe0ZGXJeKUEq6utnHC6ll2iffDhvs7h
SdKjkxUSW/phu6LjAmLBe7ltgytx7JB48sJW9EBAgL6PRDWjoiRHV00ZeyQlcejx
p7RBHFlWRE+XSIpxByHGrzFyTzHt7ND/0WGLRS+a4GEP2ZAPMQvdHz/B/zVqQa4A
/SLTaJFQVEv3ScNY9QK344buUciIPYvlIMQi5zM1lv6r07vkiIrufOl7fNepWU4p
x+y+d65VKHXDcGlNob97QlKr4mLGU+ByMF9YsSWd30zxIXunybCCLaNqQCgWpATb
386JyybIkIjld+Hc4FkXOCawwvKqJXVNj9OuDkJhgLCQioM4Jyqw68g92lXvVUkO
+ynkSLYmlFSHGgK/Rjs5xXT+X68JHVUESbKz8YsrHtncKliCU1tjBIjIeqf2kPhi
G2E0xjxmKqnlkQx1RR0hxKYQECzAza5slOJQeGEW729SDbvK2LED/a1FsTmGj9Qx
bVjBTDd7fnsfvFgKtL9TYDMxEOvngZvBND3W4XkQroMWEkBNfiYjbo3umvriPGoe
NWoDL3cL3spshfsEXvd80sTbIWusqWuqmZGcB+2YdKptSLrjFjAwotjFSn2Z27C6
ppaq6sVuL3KgZPRr7s3/3w9qRrtMr4Eznlu43CXSA7ppQOJcJRNJ8LA60QuOD8L0
RncT+LwjUfxshpV2I6dV8daz66vB0PptsDQvajRMzcfwOnA4JWeD4nHXfdfV+BBz
AcAGiawaUTl9CX6iqTBwHZ6Wmxrgs1c5fPLhM7ngOGkpo0ua4oOmyIG3+K9AJhAQ
80cC2BSTRpowXpRSySBhnraSf8T1XJPU3PbTuBQs/Bo3ko+9jKSPAu/2HUHkNe/t
N1Bvpy19jvEI8EpZV0NLHOh3saN9leJIlfEb6iqKt+SkkQp3jwLvVUPGtNV8F6BR
piCtLIzD28Dhx6gL58Jw3ve0xXZFr31LuunMZFhZkowvnFYZMbGb78wPEZAlOLzq
EC6rx/FiQZzpsRVjqpy9X5IHD++gXuhwUKT6PEVibWsdQU42zrEA+2+Q/4018O5t
WlsNqUrKVjOFrkMdhwvXlFQI0phuTrAQG+nXtxY62l/gHLQC4fFUqXUOXJ3Dwvtq
OyVkG297uJiGnh2uMFXvJQCWZ8OsTO9bKuDVBiKrsNYvjK3RewaA7DS1DPi9ovc6
9D43qBCdFUl2DWN/lwUT9/9ZALxUsD2Q+Up1gOTJhDhQt7bs899YO3lNBg0RuxrH
DBIMq7Ss5zVdNud5jwLxDvQsGb9zJvbbvJQ6nUDqj2v02beukArKCztG3D5EgPLB
C2KIDfTNY6LRFNUMEXejjEH9dQ9fdp1aVzyayvPp0Pblta7qfobIGB/jiEOGY0b8
u7Ev1Q8+5vcS9UQQJ4M/xfHNyCRiZRVkrXWItonlVsYhO+7EtrOx2Q23BxIZ7yCm
k9XsugR+Ozb/onnBRGI270MTDGLbHma5eMl2cAFhfc7RbZEQ3UxYAk1IjzV+Vub+
rMzqcUqHREWcOHkiVcR5j2Y6ZS1he5V8Q7Ozc2mPNS0NbUN2V/1gpkc6ZxQyL70z
taSnF4+Y2mdIlJ0UF6v9KLOPVXTPF0b1K9l8ZH9rzuzZ+wNvO0aCE8g4UPgmoDKG
GMok0PWnF4XsOixeG+6uy0BvrJkuOQpmKefdM5bgXjOu1MRPgybTwlnQp2TfZCJL
5U5xJKasfS5doUyBVqqj0zYxAsw2MaOMJo+nU0dDi287+isoWutK4Je+yHfvR5Wr
aT1BwxZgiHJLWXbbkVrwHFiqxySiLD/15ROfKR59v5/HrVJBgy9/Lg8X5gaWtifb
OHzTPZDypkhYbmKg+sAka+wkmZrKc6cQdMCpi/iExx2FS6xQLvdSoTeGSdixxbFQ
0srgmYbJLHO0DI6eGJiJjidb3MZGQTB60H/gKgN8IGp37Vg+idHAaIjlUcDxKJrY
sUqUzbKLLC7g4y1s5VQ/oCsLlQle1YbXbF6fULRhNBHWSle0/SPBcMsx51E0P2I1
q0VN+tTiT4Nbx4PTUWhJ0XNa0QaUBGSAypTxCx6AOhqsnqlUj7w8cb7G2p65aAHN
ywp9ha2QRedWNpfDn8M0jPjSnknchLC9yshN/wC4QDgBsmv00TCI7Tw+9wVxhllA
hnAtTQ2fykLx7LvCsCchDIYPLqTbaGqIwcAGaECJ80Gf5JmXwXnYSriPTcnX9PZt
h/ksgwOEAQ1X8eklTtmvotYN4IJleTwai7KLHxg4kR6yYkw6e/cjYNdTuUdWoa/S
W93JYDpTm7NHIJiGJJPJtU/QGDabfNM1bmC0pg9CgS0LPoWa6zS7Fj4gT5dBdMb7
shnpuhuC6ZWQdBepHoJ/G3/7+m3RP54r7VwPSdPaQIIrH3AWX33s45YLd4CJsU7A
ks68yNdatHg+Lxz25nDD2puwHj7NXXgDoEL+R1LqHvfF1TaLohwbmdo0bENCFgV4
waZ7DSbmwKoYYKraYFhxj4Orax4owss0dMk0xIzDpsXZaxy1pc25FQ/dF6G+Wdkn
cDzdDAs3MlMmCg2Pl3fFEWQieIBQIzqC5OTHnJuBmKV5lANm11tNfHpsOaNoMztq
0kMVufwbdFZFFJx8HiPhLQ7Nw2sOV6ERYXg5kgJq9Z2KKjey32J2Tz6jvKqNfmTc
EC/64Lit0eIyyRI8acY4BTRNbUfEyKrCmofGwJsu99pkAh982Vw2wI4huyAVpW0a
0mTzMzJDq1e2lWcrtN/UT4bOcTw8tUlAQjUUtmUZ+tfF4J9mfKaEdgVoK85XLsC4
FnYyH4BPSjqSBun2RoZG/ElZmV9EBEWHP0jJDoVbBLe9VC4rIA60Z351F+DywZKq
IU0KqV2L0175gSW6kz3bKY542JbPGZCHc53gy31GeuEGxwqbPkfHP9K/9RMEAtr/
k+MgiLymuW4NmCfgyAb3au82TBc/KH1gIusoUAyjZJa60umLZH+lb7tzDHNMlJ3T
y4tSkSU6hujBthcyzn2OrYydsWhhaaurCkNmRZtVZNCOrkkxLYtDrq29ohCYV4hy
GAUKrG9LU5HZUgS/OjlV9fMpnjdOuB+Znv5KFaghQU+H2W0LpRRJLFyM0F3IydF2
KAahiqeVacs9casYBDZvv1BtZcAp7bh5ngYdjEwiTjifvjGsZZeQb/ABlyVyMtx2
aPonh7IAIyen2FDHM7uBwKkC/wzJyHSXHYlyuFQwomGiSzxLR5twq2k9G2XZ38lV
/mjG0iW66LXbMPOE0TXovWVLGm5Tnsbad4PliucpgIRcAKJOhO8O0ROfqPrpM2RX
EWvrzO/oViG+b/oZzBtQrhip25hZpYX0lTr17bBLUmtDdhFKLRgSpBPipubF5KOP
p2PHr447YJG/kcv7D2NNbSPgAd5iO3w/ViMYLJW7RJBG1MIyrdsGESpILnz5fT1T
59mgLMC+zw6Y1aNegXwPt7orzWhKf/pp7XzpqzyZSJebF09DuwYayB9CrCVqPzdI
oZQM0ufmIMZXD/lm7F4jQOcD9zAM6xBFVgAFrH5oBnYKjRI7YbyZym6QdTJfgSRV
YAQyoBDi6jmiX3I5jabSutSRf6H+0YF7Keom4Ia8Xy7fa1xNKlHTCdwWAU9aVhvc
kRZcNdQxkzxh6nz7z6Wc7CJ1vgs8DqJb+fQvh7niCRoNVCrMwX0zekHMRmEVPvvw
4XhLJAXT+kBXbG7jva0xxPEaU3nI9LDof3He7hChUFiIXgzVm8JNhf/4em+XQpN/
OhKam6rOjfauEMmuQrl+QJhqbCQ7V5uCnjY2jTluOaYUPlfssKjbdXoewBCRY0Ra
0QKI3qHA2hPZ0MxKfASOHWra/6KD2GE0P5OvQsMw9f/3KUTz6qEGy09bSqVyfadA
zL8olX5Tkr7GCaoj9GAWtTOyjc73yW4kyDjCjd4WT1L1yb5Q8/WhiHicNMokatJR
0DbxDQ7UnkFz9IPUY+30RSSr8XT35yZ/kC8OzOiz/h4pD3Eykv8YYe9fDXd3VJit
Ggwo3ZPGIqGGC67MuD0SlDW1gDA92MMZTFjivLHtYptkL2Vv3VM4KjNOxuJXBmEn
oZCkI+vmYUhDvQgZgVOOmvQEj0+U+jyJ4A1elNTU4ujJHd/JExL/wX8+tF+S4m3n
U6Z77qga4l4hQmEoHO7Dmc5JGeh1Zv+YsZZOPymzRrg9mvAUfOpXfHKSHUWdZ/4j
gPJlV53O2pvd7IdyX7dxe2DNiyuSbQiIf0h3zn+vo5n5o0jAzwGWb74gXHAlyHcg
mUcQCQhUmtjKu3qylMn4d9t4GIM6Mei9yIdcrYQs9lTKBGD5z+eHrO4Z9cL0sArC
uH/ePYdnVbDsMSwMtUkAjxtokVs0CHgHqPFI32JbtMzNcSRpT8XcA4glV1pjEVaU
Wpn7MrJyndAAHjtr3xve1206MfZc1ofj2aVCfYUDSvne/KxJdKlqktgfAOCLZAtV
TwETKvqDO8I3yW1jOQBv61ibe/NvIQ1NGrEKI+bmT2pDOcn52vuMX9Exh6BCjl5c
jKkJk9rK/SFNfyNIfELaOnkv542+p441iRDZeKvANDPVhnRWC+W+a/n52K/h0rNy
TEZvCopSDbSl7TQYiJB//xpgoBgsO/Xs5j9nW7ZUf+QyAHDxfrQBVWKMJY3JNXzl
BgES8Cld2N2HHUhy+rBN+qICdc09ZFrrXQbQDOMXYoIdRLm+/AR3GsU9HO58t0Rr
d/q9gVDbCecigjWm8+unoSJeRrwtc2o6TeyvhpXOkVNdcV8Y3qa80OZEMdS2QQ3H
QNzuE8ImVwepH0CuJx5PZXncCv4fhWsmbdWenYKAMMeCMzOhrpiVA8B/xFL7UjnG
2bLVktnUyRqYWKrE3/clYz1KbX6uecXDb3U/IPfWoj9YLZqwsj8IHX/lALO3iWLB
v/kxi8hlqhJq54DbOOOnr5i/3pHD9P9fmRihNth6CVfo/SioC7FCGqkmKubjmtq1
kO9zMXx3mZT45PZqSgSwppMH5RJyCtbDgOBtPG2vJzmidPdjPDsQH7ZflHlaFugO
tNNqyrrpcsfMD38z9myHK+yazGDDPSzjd+yrdJxgnEgDNy6DmtAg+Fh4lbhydIVk
PXewYy2BJYwJpd6Hu0rG2kS/hsr1YZRdu3ErUnue63Z3zYn4CLs2Cnh07C5j0d4r
s2Npwm+RLJym3fbz4P3D5BgfkoWq1TTR8qgvOZUkHZxY7DDnx6HkNHBW/vdgz3w/
dcQesLiNvatGN8sk9q8XlYcfzY2vqpK2fbozCbrIoUX6Y7Y1VlHqzHycrSetOF7M
v1cD468Hq1xwZhzOAZ9ymG992SMOtUGb2xM7qVJf6rG9L1xX6Uvp4eL95G6p1VBn
qbAa7BIvyPg2X5FgrirBJeJ2q7bhiwruN0gitBATYYqkWq3udCjlnZfnLqp9IAs3
5FDAq+0Gxkp+WKqrJvRJelIvMH3clIfKC32agRaEjk+NQ2e8Qca5fM9w+xUmBtst
wy7BVXN7k5APl9ICpGjYx8oilTFQEtfn00E1BMwtqRJZ1YpW7DLCZNy9m1629aLG
NmR0tmUF4DGwbrxKL+D1mwFd6PZU8VoBYGddZlL6Ni1PKK0ytUiXVLvXDL5dS17i
+aIBVChbPJgebrBm3uYMN7BTlcL/ktgEZbcftBFJmgkBzx7a4wyzRNndp8q39lF9
xc73nO2493jkjhpQe0LNjw5wba6S5ewc45QQVwVsqBHfQLGBfYnoB0Gka2g8YJKw
qvoq2m34qpyeZBXZIuxE8gGxRCTXoRJwrDSQOsGzdzez0rfBawRwJ9UTqclmf4Fi
yKQGpSzZxL9LiBd3Wdwz51Hkw8KZoj+jWtU/O+DCmDbgq79vcHSy8bj6oWnwRK0G
KNeNH1Hb8fuYI0g/V0pQ02jfmAviUhaifENcZ9moL4RR5bJvL7JDky6GM1EgBYEl
9907U4L3azK2j44L0nzPECoSUeKq//E489mhbjuTkKSidzeC74+t7P8wyUZJMb3L
bbNonQc01LBhfytEU6qbLQLdLWfGW/EQGSzuA0jfbnluIUsX/08HFK0g3wFhQH//
FL9fqXpwdjeE47YgXD31AX4Omq2BuIIXyQ/J3RO2ln1J/irNdENZj2HPD+kARnjA
svveBJ/3i61i8qKJ74YXviedn+tBtO+6IdguGnNZG/AtvzMLCZA9rk5MGdVs1TrR
GldvdpN+nd2sG+DUWAviUVkTcWLKqpPgLciktRV9KGxDdFfFZHmoULNJ3SqSQ4Ce
kQ+2kX56Dq6MVXi4ZTt/PgJjrJrbHK+huU619Pw7nNjJDSkGsAESkpLphA0WbnS1
EqDsLOFqRJb3bHUPiROxNiTbKngZq+Aln46ayU0o+OXOwJwNZigsL2QeNnHYXDYu
oXomM+DMc/J3HfS+kQohsybMRiI0pi9BDGg2ZbcVC6JoNTMffmmQ/k0upqhcS8jX
Z4Y9u4eYKu0FXdeOUAutUQvw90LQWzuD0EVCpCZBu7GGKb0MI3u0GBtV981zz/0v
MGNIRfA5KiiIyJvbLf/T5osEIDAgA3DLbe6I2Eq+ifjBh+gOxg+UQTfEhELjx+W6
L8lNI+IeoPbp+VMg1FxMDTl5lB/ILsxCH1bPCpuU6JRzPysU9/8NhDvue9xCyO5W
mdyoJfpQ+nsUeT/HP0LPDXU24h72M4+0y1XYlwBCkHcvsj+xm7uKv07c/14UbhCF
oHD/JTN+5MbSg0Z+L0VgrfgCqXzYJMNf/lLspSrnxb1gNFQtkARDsAweie9lkP7B
O4v5guwyeGkNIyqQez6TsWAard0ixSwDaRItWq/qM8rrxAeYvI/ktjkMrVjftc3G
Fwzqg3I0nfwrOBTLb6JdotVjQy9YJsot5eF5d+l0X2aku6cSJrCRIgqeQ7XLUQ9y
/UsM+ymqmXqN3DlYT5Z1vOyJI+7j2F/ckvQoEi7XypcCmF7IxDeBAV/hd0n9/iQA
ymueiQjVCxilwjlZcrC1X/YA0JEtBeLo5k8MvVlPY6mQiCST7Yj00BfS1e9TTIh+
mgp7N1joKhMR5Ud/rPCalw7njh7ghRl7Uzqp4/KacEEgvQuA/jxlYW9MdfZ0J4g5
R+npIzPBBhbanyZfKPtlZr1oyQxTpW7U+xSqh0cgRNbrKReuTiScHU+UiHJxVzXD
A8D7ClZEpkxPfpeD1Shaqjl0afN3bY6x0iSG+NWo/wci5Rb28ApuHM4x+qMR8/pT
h5w74v0W9yKi4fLSFBTrAlJqgFCNsJPlZOUTW1/qojBBiBwa0m/PvBh/7XFAJzTe
cYJJl0dDv54Q5rdJHvB28oDGSfsIRyD7LHFtLTRGILvyfYuptPZu7BqYKp7JJdI6
weRZaaEMIdOvH61fL2LWpIo8wcZEb/WqWMYeUyK7kl1arhORhKC6WqT79+vibyOt
chpaTW+OZBXP9Opxlgbs1G3dX1Wm5GeBdLQdFuzOGTWtwOy5q1Bp+oZLDrwyI+K+
u0f9GXEzDLAeVAsJp29GmV5XkCIEQSvvWDt+LGI7xWzJZk2++i+n14j6WrYj1Gto
85apWdjKPLjVknkYKj6AVYXfD8A2p+7Rljs1Ob3LqqUfe3Sv5/p+wuEo7NAmgXIF
XeVsIDejPwvVJqewzuAEKTOncMtPUrOHER8U2R+jXKf4IjGpLKFpcd7wN5XuUhGr
ie1nN7UOIzHTnpCXZByfRD7lFinm1D5BnlsxGtumB/NdGsYrsTwyjuVrrbWaQrIT
hKEHQ668C1t+GEym2y9q0IvZuOFvrKd/zWyju3XkKgCpwNc8S6tQWeXvD1ymdKsV
rxjuKc6CGHFkQh6vIarzWbSShoSNfON98z8WqEPBDtXZM25uxOXozKYNlj997Vjm
nQxhzG0dLPwezg41UnVLsWChkqkkFJh7NRz2fCi/l60Mrr47wpC9CGBgafwjbl5x
q2ZpX0MwdnzXL2NyLMb3oP4EuO83S/WorRVYzUwmuXr9p2rS2ZSu4YU0IRZBonDg
Um26oAkC0Q1JU6ncF9qEMAa9iHjRGpNkSyRSQnQQEJ2LUGH8zTXlHF+9fFuTcc/E
/2pMCUjuXIWGnP5ke4eb8SgMxLI9MQ0yMiJ07JKCv1Xo6fFGvWYzGdQRo7FZJPvs
Z12Zr/D7BnmS5yH1diGmf+5ZvpdDvZ6bmqt6yzn3ZrUCIzKoiPWfb2Gh1tRmOw7j
LWVHTZPexdEWcrN51uCIpMr4XIFTAZy382U9gbnDzLqmnzdyBqPJpbzXMhU0r4KS
UQTD1N1TBDEkQZqvLfPLLJBbUur9wWHqzxFdf/VTpDeiLqSg72VTMVPeKF2mCFEK
BCqhw0O63FKX2trTX2befxBMLypelcSDdcuOb+R1rjNYj2pB33ixrkosXDud4Vm0
IJOt4uOK9RQ+aD3tlmCXnsZbCmZWoKeUt2XZ1fEOaGYoazgcq5r7ufxfn13SEUKO
QG3UQtsWEQDXrhmEY12RxPkDJcUtk/A7XqQI5kZYL2sKhA+eLr8OC/GFfyioDuXB
3CImwqbGpfBS12UxAVqzl/x3yATxrFSOmijf+oidcSaGn8SriHr6aaMuEmXVqkEu
QhLcx1yR6AVNhfH1KBJvf8aJHCb9OOmNP8j/3+p/HjZYJe2fFHiKvW/qdpmDcInT
pj9Fy0ovaoQvtSwvR9bxUtJ/CgLKSAlACoAsWcA03Kzk0+JuGvVHBe9BcqM9mCpz
o2gkJJEU6nBqYFHYcTLRjx1DOfHx72pjTp2r/3XnlI3WUiApCL7ndQY1nLZ33J7U
rifSODmomY0bEyl+g17Zqeo1x6Ly8pObtcmlM8x7ZaUQct65X+qfFSn8Zh7FiUzr
HEQrfs1E7KCynqP5XxPcdE9DeGgYJCWzt9lu97I4OCZLPzlj4uV6TjaYxDC7Qhkj
iv+8acXl8vjnPa6PshDxn9HFrPOwro/Pt/bjZMnvZrG9h1bLs3E5Rz1ciR573/VT
Id6d2KQooJdpz0nSGy+X3nYYl4K9rsycYeMxqBBIja7RDLGMWxypIyXMeJ09//1c
j9jZCk3Q1uwCo4fsditXa8HwwW/sMDZUcGMQMOEJT3PV+edHhaKETYXjTCAkCXs3
iwEtxRpb9LgqgEEBVTbGJqRJFyUtsqYLvIOMueD5/kBZNzabcf+CeGH0MLAsPHE1
stxUkZV9U34VrKk5dFuhFRXccnaTlJtPT/xlmtj78iH505UkLJsuBuQ1b2gL5BuB
bYm9+WCrfA8g40QDt7P95Jh+B9sCWRj+wlruhou7DHRW+IfKQBn4G9F7S7ihxeU0
/wpEU+2fvOiJ0rxcSkN3t0+ztUEeee46oCU64C1VwoY6zln+VhZe1KCuiyGpMbfW
4m8Y6p1j4PZ+ex6DfRS54Y11uYiqMA9suKMYXgSOxMMq4T2b/wxX4uuasIaJZ80o
nKbppTBUWNYUVMY6H6JBn4TcGtub1WewRugWk1Z7nW/ILCAktOMcPieEfI0okoGA
MLkuHXO/DKJ7i3lt75HEU9MXYyedRDHwv+lSo/GJetJ7+fEaK11rV9gM7PzVMTD9
BaMkbWJRRa97NgOkY9CsxEVIQD7cQzD9SkBiTgZR6vr1IIZrNT10vr3CqcKKTyx6
yVTuYgJvloWwXekQh2pr+9bnbSvPDvf3SLfXafaOPfUakVDz/pJ1qPb+pOwsRbxp
jU5jS5i9FW4mFyH2Sr+O5LH3v6VJ8YMifPIIwtCH4Y+iUP72PhKO5A4ZvYh5ohDL
RdEcUS5gvOkoDau6oMaR44GUyv+ycRAckeN9nbJOubyHZUgT6Qo7IU0mA+WGDbT1
2s1phUtprNGhh2EGTQ+Ettr12meuBxxb8En/9Z1iAGj82ZF/VXSqTjeEa6l1D/Bi
ucuQ+KvNq6xc+yxGdExRnRL50rmXq5f1Qm6QFnIONRiRv18bzTqgFxm5XhPjFda4
AHTEgiTDs/+EQw2I3HzEo4i7KvIwHVmrUhkXx0J2wbWOBpf74Hl/CRvixTVSL2Rg
jBoNbLHH+HJ5/iLQhe/N85C2F143KZs9IddADyGb1SQmAK3aveFf3ozL4ahX4jSN
2UP81QklARHf58mcv/BWSmdcFd6x6TokiXw0d8CN7L0kmWaG4C18fvOoUofJjfXT
B5aUlBbfVvHb5/6bT9AJt9g+SB+d2s6ly8T8RStjPT56X/XI+zoDGuqumtVCr31k
zLaRPwHCeA2JqL6bwMUy/WAuGVcnKjp1kjX8bSCx9UNzuYfyj4xpLcECaccZb7m4
TuFyaX9yPIPvENrxT7/o2fzUYQBWYikahyzxZ3T9EgfDFCmZ5rojnc+0BfjITqoW
HDUHECVTX4hplZPdNcl0j25dcn6OmRKIkWePHsmRB9QXeNp0+v23ZOqYIvyfkhOR
j+B+Psw/W3MpTwc/+2d/vS8JfDwlshdO92z4gULDqYM60GjlUKd7tioCL5aSiO9C
exDY17So8oUPlwwbed/j5jSa5msTOGByWhXPPU1RvA+SwkTmcoloAzMdONt1WXok
IflbbH7AJIpTZClDsThMYhUIH/kwxRGyHFG1iaqIZ9PStUX/7OOTL67ml3S2JGSB
Ygsn+unqr0xi2HWhRJ/73XIs8QLKRXs4570pVcQrSkZ+XPlz6GQ8Ld7cQ8TKVS+w
1J/QwD0MPXX8SVGH5TdkAclcz1PvgQHsAAqByEhGytckh2Upw6gkaaEVGBc3krqo
GkdZDO5XhxQk7JUSJklfD9jvUR9kmpNcQqxMSqX0WyCQ1tNthyRvDfDyjHE6S0K1
Ub53FQYchxCjHlcFh+XG/ejGzkEF0wPOZyTEId0EB6LazqoGf2SpEVC7oReGpdqg
BayN1p0UmNxcmy2dFwZuSfnTEkc27QYJZGB9aSXVrYE8TEWa0W6wmrvd8GTnUeXD
5ETRMJjagz1hJDOkAzxHJDdBggT3/b03UsY2A1T4c2AGr1f8Ay46nyLgRBRRLt87
jNQOqqsBKKnYvquJ/hIzy1sVaRn2UiFK9RSjuagUQv+bf268WcsaaEZVR237GW28
Yi0PRH5pu4NUbxrFPODQMg0lATCkeeQUzuyoguniAxxRLHzLidvJLGPEL50Is6vT
+4bxJCLwQ3Pi955hJdazP6i0Ge8jpo+uw9vUity0/jOBC6KwWaL7xiG5aC8iUSWL
PwAGbKfjZeVt1zcQKnaUootElTbM3xu7nZGFRlR+fP9si1cZBz3DwnucDkwjYJWk
I+AcnkKLWiChLTdsiqCzwzCHxCoNCJWIXhjZTdAANJwkZR+ROLqSJ2RyQWeog9ei
4Igmc0gt43RNn3b0djGCd96woTpGTyGpDL2PqD/eAVzRDU9CCjojiFsJT07e3dtT
71elS884VfgWSJvQh2DkvpscivtriXuZavHx3Y2VKZNeH0pLCy75WJXHmPB9kkdt
tMC92oALvL+SfOlasNhSdADSG5r3xJQMD2v/F0Ig9iWmp0fzxIwnZV7y1QuSImWj
+vrg0P4fLV0YaDJxS3U3MLofZiBvLqk0IV7WuS3xudqtcmm8iSeEFIf0Qs6dOU6j
52tOQSbmoHr1VsH7x7He+HKdVVXUs1UnmDHuhLNUys1HIBUFhbBYmapHf6tvQwhz
+D6KjrbZ2N6jbJyLoGCNDtWJqWBguxBjKu5e8PHKXBVuJukfu8GIwxMeNKybCdRk
gV6WI8OtxgYt3tCYzf8kQ9dG3EHaFxc74WohmOE42MspjnRtU9URjmvCt6/8bcb9
iAzTrEqcc9Njy0Y/sgbCtlis/6t49e6b010g69+UNDqysddAL1zcliB6AG45TBPA
/ftqID9szIR7iNZTaoS+nPmb04UI+pxmNNMZC4+GhQiQ3EE4O/qI9p/noGadc0qL
8vUs0kTwo57MwbHM3A0T23LDXdsQJubFOjU+drxfCAo0gbOOcELDDR2fppSRffHf
M5z3pORekJ24KCDPtZnV5j6SDvefBLItSoMSLTuHGYPBU+vgjURR7fgct4oSqH1Y
EjDJARi3YmtJSm1ED6Ncz/iCQW+9p2uyCiIqV/azTXCtU3CC2rZE0QPWLKJhmwI8
ucYzQF6WuLSgDDgyIsHOW546uArZG64atu8Ms2RiG/bFutPPueLV0MoIwnb8H/lU
yEFZ3EoxqDs0A62ERGiD/b0woE4DW9JzyqRbyNayxrPyeMngQAGdR19MzUBcQ9gd
4IJqimWiPcsaYS6u+b/IJGkR0hO36UpgjdFVnXQtKG2H4ZB1oL7bDXn2l54sPgWI
QYE0/icXtFa6DOu/ZjX4rOHTAEtcZTmiDYKzStYhRfqFoa3Oc3SACkq2GMJu5s5Z
gWpdIILmJF/K1B+/yYKjYdwCX2WgPcz+Uvh1JhQmGKeD79mMGCLVqBf3k+JyyA8d
j+5+pCHZT08BuNp2NmFPvHi90UsEjDvWpqGTIyYEOOU32EAdeaamK0eowfuJzj4z
JE6nNNkw6liXHX4HnpXCi3dD/OVQaPxq8fKxfdFZA1CU41g25pyk3iKw8EBS6i6u
ZcRecmT1qq1qHNEV7y/X/EToNYKZFIkKm6pBwkUTwBOodQRQbn0E/6sZZ2NthaLQ
auuSlIZ2lUmtbGTHHK3f1nf3YMqljsbXeaRe5ZfW+GJVr0JE+te/DVdPF7Q4GTpV
U3gU6fS0RYw5tkGlF1ekHQAO9KtAAeMordfiN1Y5VigM4C8TnjjpRaeUKLM0px3I
w5Ie/70ViiXtUgpPqCrG7GybiOe5K22Sd2hFyJGdSCveck0gUWQbBw1jb6n9cFpH
BY9U1fS9Q3JYRQgBpgwTT7lRfY0Q9/PSvI8znZ5mJ25XIR9rJI80xkpja8nRPGRt
E+aJECxSXojW/JCuAT7llRH+3Zy5dBFaLYKvq5FQUCyuJ4Ce1qOzOR5Nw43ccJxU
cSMmK8HuXHg/DNc+6r11F+roDXvOUYCkf+VZO9U+brPp850kShKDnuApvqq6sXmr
q5bM442INgv08hFEwG1i6w87XXxf9LIBBCzrmqBMafx4YhP9qq1JzAFwV1WN+xdi
0zvkUKOKpxc6T+HcdzcrGIz3orVzB7pTG+lVaTEFSZdIqs3/sbdOtGZanqczODPW
+IcqNxT0xNj0iSYcTxoAqZHEiI+6nhMkH7ig+lyFcx489YqQN2cZPKCZ/4Groqab
CmblSonU7XOBSCWRvnDYy9S9775psScYZpxJ+kc4jXCM5JkYUhjtnKR6td/XLrg0
sBnoNj9SBGX6O6lfEYyvQzbH4PAlp/6IUoNjaARsY3Ev1Ps/lkeIFOTS6Dc5Tn3x
dS7yem2kpPLAFJVTNh5RCcqAABO67XnR5CuY4V3x1le3oyzTn5IK+oJ0JaD6qAT2
Sao7B+yV4bTkjpEy1uaiJLElrxajLHKhb9LEx9e5eyuNQEUSRl2OhZFc7aP1ezrg
l1o9EGctB69HpRbhWSpxE8CGUoc7+uCO5w9KqzgLUBB971seF8/xHBDtzlqXoIC9
YcUtFIYIG8S8+KcWWWPdBMXm7B7tZtgcXdVWYwPZZzGPslQvr/yVvaBXfAFTQlX+
w4cXNZ8QHdbWNheNo06kkBDwq3TELBD2mTC9p7CCv2Gcaq5B1vJyTChxkPjkb2gz
seeI5C32CEOMWQlvtw7rt5W6EK0YIjign9gz4nyRaszIBFQK8EX/V17eUFCtMkOO
2a7AmJbAQZhA2Tuy/bcDPNpZ22MQRdATaE1ahpJg+9T42UyvAlkhoyz4+xDwr9Uh
Ci0+5syvTlmkynZ3mR10v9IYDkDwdsS8AylLkRo049htDyTErao4BjBcIVbdsOSu
UjOgM/hhpQD8X1Mwlhp0X3PaB85pDZDHC+0i/Y2o7IZwpnMXrUnaWBdYLucj5U4B
0hPJmQS4vxbB5TAiIn6iTTcT+CBnUz1eTrgKKCAeHs4tlLaBFrFZTH/lP5ShSQtO
B6M8bYQFiPQGj8p3VXU3TRXJqIWnhJIciG62WLSR55ctmLjjHvGzS2NbeOdoojj7
xxraH6S4ciYHYJrq+vQJOXpYfqUMPUPltbz2bUldoirVnylckIQ9xqTe6lC0nHZG
idgHVlV6shqRGmVG2rh6fXdh/+yFUcXn1YFo9MAieBPoMvTxVFjJSLh98feK4FPA
poBmc9P2Rcyc9Vn9oMFM2vl5qUGIkni/uk3B+R2fBlDWBaYOvyKPhxhLE0M/OZq2
zMAb23OKwluncGxXegYUhn5Qj0A5HsCsY6WkwGv6+H1XPbIVO/eth+ne5lZt/EB1
TU/JZgReChPFaxZZglWMRjG/mybtEJHoOnFxS/f17FCd0HNRZ7ycVfZq8l35RrbJ
oekeCR+VVY/Rnf8Xb0jYc1cItejB7KxB/8t5DjYjWDr3ClfYATAnIK8vSxui6QYF
WfK29esZRCqxI26pDOAasvitI0kwmF1aY9F+C8a5+Bzy4p7axKz9B6DPhWrl+xI+
JKGZE97N5utaHQqi8CO9Rwb5BqQktN/PmIRLLShmrb3vsz7lKoHEpzUtfljM+6md
J8JPuvEGteHcfabIDJ1v3ehtqe72lmSNurslAS0s5StU0TNkLigMoNv1VMbR9TkB
g8/H+hGXPE7G4nEu8CPLhPyhqpwe+Imgbf3zoOtLnC8Wt2IL3HgGQ1cro3uaO6JY
TxJ6SuyNFrjpPZJOXixQn2zEV+jlYmvFdzbbgUC/v3Xr7JKnu1DvULuXgDrmGEye
Wcicsm7pv5bt1JU7E/Q9bAQP70UmTNiXY1QYALnfruAtXq5bI0SFh5wT/iGlM6Im
pMAzxw57jG+tdqdi1dWu+Wj6KVGpSxNGaKX07zWmsNyNK/TVNaTyeFWY0T86huV0
xFM6uO16+D5hGh12JmQBrUADcYJIKi7w/xFzYHuyRpR6ZVeF0To2iwu7izX+OKDc
cPlr3MFSO1UPfhViaMnZt6Ebs4Pd65L7TbwDINFT4xOvS/WVcpoX3OMYn9V6toKI
F9FTecLiynQ3Bv4yM2FSbDy6J5eERv+Dmj3Y8nusmmh0wZqMHK+0BZBcns9uReJv
8lgLTCV98w2zN1iWVVNwvaV5Hg0npccy5EAy735WV/yv6s+yoAHu0sRUD063xvSO
UOT8eI5JHw8UMzTM/CznRzS9C4R1Al5FK/qUXPePSdmYZLJ2zNcINeRzYsXvLa8e
Zo+qi0H8lRTHdmfkKwuacIzdN4KWckyFjLt3czsRd90v1IS0KYwFdKML4MkZWXzh
xMna8+1IQx562TTAVNwbLtw1fsYuIcG6ks7tzIoaX67CS+HNv4QmXqHLoeGUeNLt
To8lgrwgiDd3hiy6tDHezP8xgVTiXCC5PVDZ+kWAbjZ+UXd8BvCLyIYWRyU4eXSj
7VPRaQm80OGVkmIBAKYDa3jKbEC/x5O/8dXXIID3HnqqcGmDoSaTf/nBQAmviFUH
iwx+vmn73a9witGYZUtJ6AL0/O0YLqJvNAiSzC5JWONWhyH5sFpz5ph9dxshvYNg
76Gknm3RUnKqDTNHwIp2sb6EDcWZzQDVgF0feaqbpDa9QSXITu3Wh6ms1AtQoF9Z
Gg22AomFE8AmtXAf03L60MFFV28qUyYMxgxyVmBdECsM9kZi0NRA2kssulz+kA1L
VMIyLREN2EaPhL6vaN0xSaNq88HHaRUbnUCBOu8TlGXl59hQcbjl+1Uuq91WpUtM
RC7xygm+LwZ8HOK2c9hc5OsMyfa3N3bDH/Si5r0i9cMShXygDQEs3GcEYZFXKUND
xIDaPUbhN4hwYF00es0dL6zbh/ThrMPVKNPNoFkAPArMv59HWrJZrc7SqKJF/6O3
yP1W79DJDncBThhulvtB1ljq/p3ycyDdX0c1knPwna2Wklq8Na3gtAhUvp1vvUkn
+YavAX8myQdlBY272CUoSpicAOuOgr1SZZ2cSKmD0U51nWKwWrFtoZkjmz4GmcrS
jkO3R2jtEra1+8hCRii+lrs6nZftoofrQZJyV+6c+JYh8CaGJA4N83zPI7IgPK73
ztSPKzzhmfj5F5YdALYAaD3FSxYrfCFrrjY/8qqb9AAQm9nsoVoypmOdP5Ne79F3
Js/H9oh4gU+wdthDicFcXVAmlW5O94DjUQuN4/5i0D1s2vC6FLOYM2EfizwxFKsm
Gd+Mb9iPhuiAVIRjU/XVdjrdctUOQIExKu1NYnyoxLjItYldleBd85LUfcZ5sCMP
4QqhRkViX9qioa9FvPVSxO9KV/kVdCisJiC57yOH1fy65NaC5Mti/3Ey0Nu4BmQl
pWQWy91SXmeTHmJyBbi4x5sgDQoyeEODRUFIVUsOFpqX6MdXg9YRD6HNGRHhNtJH
Gaz7QHqA+wyQWEp8rIeeqZ+XUrdYVF8/fpKAhCYqxMlyrZczDaQvuu0pUYmggktw
HI++40nUXsFtI/dSkMiOwbyKozgyvTOUUKHoFMjB7ixGxugB2XnV937G6ppzLN/c
HJQLQXn6d619vFysjIQxxOhxCpvNI57OXv9Cxtm3QnPezhimzWmCK4LVhjmMgRSj
XsDhalr5sPeGOpLznnPgNIIpDLOKB9i5ZsmLYjVi1JhiEPXLRpltMCwddyngWD//
0EcMOG01aeH+K+HaKQBNqjr2WyxhwxLNIWQlPOGrCddrgdLlCUFn9nFVWhy68YN3
ppFLo9YPY+RFV5nz2E73EKiI/NL5UiUi95OOCP/ZQew12UlnmEAWkqLHgB8Tw6aE
Q39T4mebPMrHkugLgXPM04yN29hIntw79EW52kywLzrcXJSe1QIuXWcOWfffS3Du
0wtJoCph71F7UurV6GK3mRZZhbeMD0Bs5LN/6i20jnZWSsLQjBNoGmEqBoW+ht3V
jTNJ1ghPJAHDMq+kPgjQlmP8QJgp0bnOKteo22HCebjPPEAIKYq4an1PVZc8ZAMr
p6sc79SrHpVIrhYiBQah951OJ8lVXwlewUzvxvVmmOqROc//RlEMPzGjcHR7d+R/
q/SW4bdqyPoSnF2lFvRz834t+LzadCTN0Uo92At0YwiAJ3iRVyHphMFewcyBpfno
+iUltLbHjNIw4ONip23EIgoF++0p6cClyYpIRbfC1pcDgwdIFl+vYjtMHeuiw1R9
cU1N3EVtEr+LtHGsDy3pPIQclkj/OOIwjd33H5lugKk7X937U5m47sKH8ifo2b1v
tTXDuf88ly5Sc7uP3MXN5EyMQ+Rngg7b0nd8smhTS5Qbrkg+QoH21cXeCF7BWVX7
UN5nLClI1nGfwOwa7WxnlFAG9k+BSKOVFpSK1p+mY+J7O5FygIMjJbOpX2uYvW3s
Hbird6A7p7v8/p1nPYO2HFU8e22pjuVysbWUVuIszVZgmYTOTLvQOBMCsed2vpAB
xiKKt1cUzpmqvfCXzuAJZO5esBIOCivqUcyxAeCUub8vSm2QdbtceTSEW0L9TiC0
7Srh5sSn8D4WROvVGdHkFa+eRXBzvaCOEDm9PRT0j4aVWvP2AoHSYQ9DYGpZaf/7
Mq0m1sy2LwJZ8j5I5rMo8lSvTSrvC7/MM5AoXzv+socH6ZZ4e1l/f6AAtiZJWjjO
97CJCSJpyAvulo5Qd4QTGP4m97f7IDZ52uVG+QtgtoQZxSWbIZND/q0Ex4XhqaAs
pLqxAFYnRhfgoapIguqTBiWzCKv7yXvtYAif+oxSAggxRLsuYGrGE7aXG37GOEH1
rhvAE5pXVoJ2gKE4o7vKRbeNHqB4rbqiLIvaaq3F6wx88EJJIcBZQ+XbqGY/RIKx
MPPAlxIJozmvQBq5mSxCDOBzGW4DLJ6dOkNajilUq+qvZ4uXlClzEhs2AAD3Wus+
rmiWVVUz4/FqevU+GwpE0fSI1bUTcepv6vZr1oU9gFsOT9ypSMpCuGoVhpvL7Jpn
gYlmLKtrdBzmZD5MVcWHBkMOuMICkfpyp6zRIkuxYIwUmw9g6Tnm4i03xORIBV9R
IC0EeR+QSKhY8qDH58tbSQOXhuMGEvqWVl5/Vnv2f0utff6flhH3mqDHVX0TodQi
Iq3MOqL19rBLLp4A/BsIIfFY6jgEgJPYE0WRVsgObgZNdewqPqXE67TC2OAGFxhq
hhZAs74/c/Mhvfew+Kyvoxnn/DRpgX6x57PXhHsQKCcOkMLdRJ8X+x3e93Z2XA78
eO1XA4C49/VQSg4k4oJO7UC8bfDZi7ipncOKGZyq6t/1bgfJS61nY6H9u0x7DUXi
VKgRFZjrjfcD0xb0wH9XtDi+hP/xloiRZFaPW+zcedS3FQIfAuQcWigmeebZsOEB
YZnRfLnx3JMLfTORVvd+mWXLnlzTDU6hDKmkfuIG5eSmAqHXgSVUq/khr0s54oOf
Fs2ABM5Gnsj8DZLSw2JJgAJIS8PwT6jmDKrFVNSkS742wDaCzuXTvo2H/r9no53A
jQC77mySxmVbxHXnWQkIgjioQyyYbUxWgN7V8gZ/iOSL8zuDNMXiTERhOJKqQwf3
Q9TY43lJu+IsQ+95r1rrqdpQ9EpPgeXV1S9+AQsjL3ghgTcM3ECVpR2ylXYgtnTM
9fTz+NBeX+kNdbwaLkiXFxOXYgPJiMQhft3r8DJ9M7YIXh66jBZjXvRwIODNMUrt
NeZX4VjBM6pKKkgDJwjk4iNABt+kNK+L9W7kLKkQLWw9VkPet9Atxby80nD9+aLv
8wf/7DtNR8W6jnkgZXp++xgKMo1S1vy9rqZ11Sk/YTisenGFj41TF17lQGJrDntj
a4WYT8z6DlK6bxIK5m8wUK3oag51rmEUL5ne5vdOFcgDrCH2HFG7qmxkUdpw9wJt
rcujixyNwrpkR/69QjSA+nLrkvhiwCAN/tSYlRU0LG+s1jvVR3ZfntkhpPcUa+kp
vi2rWJ05TDC9RyrP9sfax8UlzdrecHQIGOy1xvEUEqxbRyt63kylhCtVbDB0nivd
hpgieA2dxlAJ6NpuxuLsudaF0VtPexflZRKfOvI5NefAJVRc9N4c1pchRBAN/14N
mAWZ6i5Y3LZxeEwTqYftdc5zfNoUWhlGUKEyvSqZZRF/hISXdnGN/4OTL0arfbww
o2u6tM4F9rNdEV7sNU1HNfIlsojmVo6fe/K46Fka7vSGDNRLV0SWkxsns1OOcG8t
Nix2do84W1Eni159VfOqq/WDLZ9bIYtUb9zVQ7TcHmOgMUQD+0lRcU3R19sHd0SH
jKdgypZgz08JN+QQLREiqdN0iEm7i4vHTXvxk6qdpEar7Y9f/Yh1czlKHL0n7BGQ
B27xVOMGdxvTFknA8zf3Aa09w7XuDHyMtOhC9Tcrk8N+rDajM7pYosw8s7iOfCJ4
i1ASCJmKzRIipVEgFlCnr4f8XR8HinACod8tb2y6Qj5z/a/o/nEr1fPf8+lajRHM
0CA06DwKJD6uSZj5Nqmx0OVrkUoza03iqG/kLRdTP5TzEImc1WNmsMRAsHXKrZsq
cpEgHf0YX455R2mwP5A4Q2Dd+A+xQXED+mBcON/cMRInzepGm9e55EBaz9xeTs5W
JFZQp0FEqm03kRHOoydtbVDftavjRlGHS572TpzNCpm1uZA3DmEr6NXlcEeTI8V6
lQQpNSY3kqvVMWzu3yI47EiGpc7PqQe+4RSVcujzNQCrOxauA3Br3JOGT3sPkIhb
HvhqhHB5rtKWc5u+4F1BwbrBi1AHIOWSCSZNFjkeNjQ8S41ClGtZ9WAXiFTYWLK6
71QA4N49fRkLb+EXVCfKjjMwbvk+HDlAYZD7DQlbuXJiBI8uhkdq2IIinfO8kpUW
9Kahpck+TSaEMJhlVYi/pSNybEIApsbypz8T1eidE4PzkwLpML43Et/Mw/PSXLmI
JC90jav0zIE0hVUOQuHOKA8D0KMhq1wYbOHT3Sx5ren2jW7GjJh4tzDMUlges2Tr
UAWhhdZ29mQWvN1p+cO8KKcCoYxwOEJ4DDUd1XGK+10LwCKnPjKbxO4f+msj6cjT
s0+UE457k7mQ+kloyRBJU9J7Lrrkgbj9jupu0ZZq0iCVDX9JoIRF985WzVApVwg6
MV3/92nRPcQut26/+sCsoIkZm0C+r8zANxluxw0aQ64vO6WW15tbgclPeh5nSB0b
T179Y9K2rYDQKk/wIjDkFi+ZF312MdFxdHPSyloKbKBLDxiZN8DFLGnM9WODbOLD
K5pfx/rUI27yuZag3gAmF1hzFuKfCHniABxwkFrWYcyTy7RZX+4XDZAWADLBgmrL
U0v5bgpWWmLLXDQMLO4JBaVX7MPllHMN6lsPCksz76OH1X2bQgTTmWL/HTr7HM2S
+19TWwHwNn+FZR1e9RLSLjYqz2CfshEtxFIGhObaCGZsFTb2weiINqjOxSEPLG1h
QS83M9Mj3Xm/qivI4HH1eGAcp7caLXoACXb7iksTj8Gy0cgELFYGYXwRe6UWplN1
R+sIP2Q6yrvAV0Qrr1FwXUbZHbIQUPvgMV9i3SIprPhtuZx9Wj/3O+BEtd8d5pCQ
IIVaMsEAo5nYozQwe/FDlxlOP/BUBrdlzjdtar4oob6sm0DVS1mXGEwrCD5EpUm/
bqlaTUPzkLaRgI6HRFet4L3/pBbo5vKiGA79/g/VJZ/su1iJqMZJ6pAU79ZS0mTd
rBRTV/vwTAaiYdk26MDyFFFXyfHoz640+rsGX34L+qbuk5KOkCaad8q4Mm8jwK1Q
HbCfGSHxa9HT68ZR/uWp4FW96Nn7Y1eM/SbeE+bGlK2IhwrJo9Gjye1XSTRfZZyX
nqIUtdxuEjQJbNr9viNeR6USvs/FQ3uuReaa0E0ECveMdgRS18Kbyx5CrUC7RMZU
5CItAOc5iCnK8or929H8AinpDX6/pADCKdc2rOldqC5ru/Szp5R/E0PU23HW9Q91
ed7SzWT1ccIGrvR+m0AV4c6rLKCjan3PoirFPOWr2/DIfXu0/6lfhLmfei5rHYZt
cNCs7rnOpN4XCa5H21P4Ko/iw1AecOsIguP3NF3d6JFfOLxB3BDnXwBP9QPDhky/
K3t6P94FYyzpShwDMEbMuUO29E5PtiQpjdH9MxG4F+iX+OAeMlbAcsL3MAtsKx4U
/kfDA3wcaIQcnn8UK+C8wsxqWFbIv5HhCaF1d04nJk0zJ4P/0AC7jGK4u3J7tVqy
t31fHN+02bRuE+rio+fgDrqa4/fmFaJpbaf0SwkitB4uLNTYbY9ws197ocDrGRYf
Zyn5RzppDir95T/fcqAQ+5sOVpxrnfNdozataxnct+TelcyckIo+PkDxpVdhnRrX
iVAWBtfvxCGrjy3RmF1O1LiSef6vBS6x+/cjIv9NEh9pMtqWmz6+XR2Zw5uPRvoE
Z2zJUwbw+AyCX1AwXg7UhB+u5ldlV5RFic1i96j9jRGPyO4byaLVriariz0QWMG/
xbbTbnj2H8VguQyoAorAFA5j9Zpw8YQaDbk9i7WRWQjgdouhK40A7aNkhR8l2zqT
xteK16iRcCSlNHW0OUZdX+rK9iW+nVbpkvFCDep7zPZRt7ZZoreVm6EcyHD/G10Z
Y+jmnemHML9Iw/biYOsHLczy1GHarRiVhFoEkC4ItizlZ8IKJxD0A0RY+YK7n6Ie
Jkkr2cAjBe2gTQ2AIOeYEdJFSY9pFV2oOQib3rF/LietSR47JRzIivJflLAlGNy9
ZU2K4GaLNY9y4niQz4DzZXUVByAV+DbKFfdwpU9ML5PKGJVht+0AN9EHvIfi9Cfb
NXfQIIkjejVCFrNC+PCrVCD9gr1StMAY/KXY0lONcQB4PwvIk68936rWuZ+fdAjA
62QEMXoITl8ZwJpepKVthrM+L+Vl1y4LGToACAqbQN6gxdCOkads3qr0G7jAVyy9
xiZbuXuYnlXo1sJFPyumRafwdNqbQqdQTO8v2j7zX8niuHrJkGNaotJgFgDJH5pk
t8LXSnoXihGLNUW74lJmTzsbS2JBMvH2C3t0D1qI4r64LwyxgQ9ShRxRbxo5vzGG
x4A3IUDjSLjVgp+a0/ClJLbmiOPDdwMJ/PudermcQZNFiLePXT9jK1i3CCzf/dBL
TkP99b7psp4CmKOeGz0fAiY496SsGHMyorm1tuKTYXhx1mR2Fwc1Ud13FF3vcrG3
BAA0vLJMaVWZRcvNunxC5XQIUdfShW43ZLUgLFkeIdzd3HpEVzo3JonQ3waNXoxm
mI0qFEZaYCHKyon1lY5fpy1IWoyRT+NtaDGD4CgFx4XY26HCQlQBbo1JYUEVC5ES
2GyicxWsCF/uvxV0P65ywmstFOhAmX9P0A0zZyRAiq4gsve6KXkRy685ctKFpPWz
5W8HbxcbobC+zZvxjf7NMGOajEuZcqkIUH8Bc0Mt7WYAxQWmk73RagetMg0g5J+W
zhyUOpabTKiKCxwnwt/5FUOHGNjxlis0UDwTksRYSJcJG4+23jj3NjgUkV5ctXXO
ZMz2WMT9iB2oDG0yQTMJzE/yWKGnmedDPBjID34Jwgg4CCkCCq4C9rCmBiW4Xw2h
VqkjYNBt/5L7KWzz5xOqL5w5qkdtbuse7JgtKTs08vSmiQ6DF8XTLkjA3xG4tqOP
AaD1o8C204ihV9GFPhxup5auJrJNV580ISOeQFjjB9JJWHW4lFFzYI8J+F7S5sfY
VXSgCukVFAxWxTJoEmbhOtUO473lnFIlVs4buC6uX8oUv/c8Iujo3kovyDf+9LGA
EgvnCqBBsUTIXs8AoiRsZJrBsc0CD1Ft1kNAZk8ly5zUlgRMYTQXq2xKarpevBc9
sBg1FcuUggD86C1Grrp9p29fov831dKHrLTOQabF30uyBfoh1l5LsNTR4Z3J6A5Z
V1ab3xskNKmIXk8VvbPGvUi1pFMmAONtRe2jdHW4lTA9P+C/APV+LCCRvoDcvJKj
eML7Q1bDMTP9d+deKuI4P8R4GpMJAouKkaPcmqfoUtfPdzmleHKgBwBKc7xUsLGp
67BFwLHzkz78gAD8JhBzrLxzaEIJXCX55+tGFfhNRZ1zwWTNy4ld8h5zVON4Dfa7
11zt6u1UH1pbh//KTsxtROnU0RKn/oN/JgMUuJd5VFpG8swf71RyMLbvY07DBugZ
Ehi0knq5rcf2kq0dNksP0FQ3I+GNdrnwfxZ+lwHKfQb324QRd+YsvZgE9v2LHRnk
ITy/XovC81JG6DtTfCKNcKeijgOz3rPEnWDNa2Dj6fcNe0lxHHOhg9hZtirdW9vE
KDBlbZuSQ4d8YpvK/bU+iE/iSJ0MXKhXqs0Fegj+6C7lyHup+WK/NztGT8vQyytm
XqgoUuptbVK2zlWH13Vj7frGSSbz/5NwoXEww968EKxE3SsuCyCNSIRJzf3leoDb
sfY7FHHYbApPTywIv0GNOuwZ5+8g/i3sagaYnu0yHiUcxG6UiRCaAM5HjYkpehgx
EjURRLrgzj5rLIxdiTpjijXtMYdgNEYGZfFV/fnUiAJ5oOyWZ88vkZhfiiELhbuM
aAuwTHNiXre7WP5gbXva3W0vDzn+aN7CRybb1q8DGOHzzOeWMXkMbpwaChRcnjbA
sagKyq17XvuBIPF7cIdXuJan6307j4rZbwEBln0xrEUD28s9/GAtSBjzYBYzf620
Bsl1UyTjWKDs48vHhQSm6rDG2ef8HXr2yytOghR0UaoJJDn0JpvbIgx4xnWMR++8
rP9sjlbMtpB5AeDyjnajl1klF8NMgF898BKeAM9UNnLyGZgAa1itOcFtfvzdwz7T
k72Mvst2wHSbNRgL2HXx/tKBZIF6hAXiwtC5qAau1xd9KT02KFgR42uqLSa7LY+4
sRJh18s3wpyY0GDlb0Suw0Z7bzkPdHwT/fG7no7hQG7ZYI+VKPJN8tqsceWrOyhI
8nATmHgJrlmWXD860bjGfAu2T78XOaf5RpTKfMZ9sSwPQr1RRBxvAM1RaboKFiWk
gRJsWkfTTLXdaJRXI2zwc65YeN47iWQAnd5wJMxHOz3DBjDvxGRmm1hJ7FaouWIe
+3L0cnuos334BCrr5mAH+Sj3xzS3553z7DqMHD1yz1ohHC08puMV2g38Bqjqueic
LjC39xgJpSlPWGvih/9V7JLE4F3goDAzqJRWMDGdhWlESqAgGqs0xUj/Qd6vweXa
TKDz5489lj17amMY/elNJDpcKs2WwsE/tCvqNOr927+Xk1KSf8Doi6THqdJakBoH
xzLfAgVAAJzwRgp+BcvE0CqgJfFfot6APKAF+ALAEgqzhE2ThYWDHUoSyelLU6tM
1RD7AnquB7julb7v/cHVApKZ2ab93y2M8XATe7XmiEB5C4PMQF7N+exuKlxbUPDF
8hnYM4xQKbFTuDk3YGnyXQEjzJun/m8BLqUzi43YCOy2bmEtXq+8wsMA9NoerQc8
TbdHkYYwG/1RSaIdpx+9u1BhdqpnSYI9Ba1uovY1U2eLHqYlIVVUHX7wNJojDtMr
rAVt2aO+3hg3ay3jWqpbRNGQJ5gg+7evP7WnrHacfC5v+Zmnl1/nxLNkxh+IYH0k
0fFJ1jjGdn7CWys3UCnim2e1oyRaNNznFC0BVf9+9DZI7HmdzuxR5HT82e4sYacc
AAnGJTiKEkULECxvHo/jQ2YYTBBtOYyA7AMM9AnqUbk4vhhOAOJ+CpPlg5LXf38B
a3nfpl5vUKSwlFZsrA+F4n09hyX1ItPxpt//1IXLzTxyo3LhOfgVRdmiTd7bwr8S
+cTeLZd0DFJFaImMjEI7tID7kf3W6aZoXUiWMhnhvnQnEO6Zy9ifU4asBTkeeNLn
bp7NbfM3/wJI2DnZeu70B7iKikLFFxzSeUxxTMQnpWP0zcjXutD5hcIoDpWNM2QM
lYE65T0KyOe6ue/Z7kWClBwVM7dVqaLa5KfGOU6d2OAfUN7K6y3UIDIbGZBiimop
dJOTZYwmXAWfp194njuan/pZyHLg+0oUci0ISHkw8NHUSC2ox6H0C1tVORErBkCQ
neBj7BkiXt4r22wnrLQB9cNU4GnIijm6Z+LyYAQZwNnX8+sPgHwiBSw0HkRydEjl
IKI+Hd3cNIMyey02UEqMg//1TAollo5UqkolWJ4+AWV3BcmEoFNgOMILaHg8r49U
B+1lloB1l9AFh3B7ycd6wlacN4tTnxVSqThZqaS7S1j1DdlU0Q8A4wt0RUswH6UQ
M1T1B431eIB60DEoQ8jmQKPyAGQO4/gQF7qhYEY3Of1/CPrxsaUAp7WBALIzOsLF
urpX5kS+vpaKg1IGIkZs4DPYMaUcJUfdlunGVs0ynZal5xWey1cZ5yZQClUy3j1r
ABspvVlOtKJyFQXaITvBGMzQ3zaEdsbr3F5/o9wWPmvw1RIF4vkPI52ZLq2UqNsj
hPIdqbLRHdaa2MIpz8d17Re1+p07DYYPZXQ+tGBkMy0OkbWwz5pAIYcyP+BKyPZ2
5BEEX62YS0nrTQE432BOi27vKA9sjIX2/cYhwC5o1vX1XrmvQ3vog1RHCq47p4Sx
RdgF5+myjIIKM2w+8pIfmw/u+wLHVSiNH41F7WlfAAvHxgC96mnJWvUDHmO1lCCJ
YM7IIyUEhgXoyFflZtAJihcQeMc7bxHOAemapgOv1DoZd3Kzdomx6Yggdh2Ki50A
eiqh3MJo2uFuQEShpx9jGht478mpcc6NiC9IqrRQ675p9Pj5iqbT9oTwplsIwulc
/YCfc0V/qrXk0E9CYYR98OVocnwt41IA507ony7BPZQwdwKFwx+7YzpIdrgl1v/s
y1FeDJy3tPQMZvB8F1PW+f1gWN87mb4HB9w9Pc3GHcoZ1ILAyI8Fs+eEeb/NiW7k
xw4fZFVlNpKtW82B+qsjPPN1xO+6eKYboh6GY9nooyeuj90kYcEyIstsrgjVY5Zu
i6iQhiDQ+vB7evz2jpymuhMTLUDy9kEoovP3kigpzvRub5rycNf+oFJFiqJkp7eV
6eNAWu4XDRxOvDvtFTQ1/On4bQVmqUP+AyZbQlLwSWk/3mG8eq0sEIBYzwXG88u7
pM8z6Ael1Bi4vjkHR11wyjepsryIgDwP170dYntDh/ErZVi9c+ax5KInBttvTW1U
pM5mrSuSmpUm9ARXCUtkfHv71al9Ht1oV0zETbkumzb3rqW2MeR6h9UJfaK2197/
QtxBbZqp+g3aIiMaQwm01c1UuaKQKEO4zTnaXba/D4dD755/Wl8hhua32Jh0DWQF
R4DZHkrgrj9/lMDeOsx5cc4XafSB2KcKAh5FjRuIVd7YSv+2jJPtinuCqXNCZwlE
XpkBjTr8jSJlJQzNc56Q14PJmkwQqQZvrzJlhOZASGOKtrjqT5578hXvosn9S/+Y
ySw0g5B5KUwBwS70kQfqXcFWw8w3wtlDEdlr+O37SPdjSWRKAku1WtGbhFICk7/F
oT+neNhVWzqlouZTb3jH+xyuFQKwOz061rH0vUC4d4f9BOlzx1JuVWDjxHRZS6vc
Gw8ZEP+35+DPuPOgEqQJCiDnLS2v5Ih4x9Vtltane9C8xH+yDqijMipqVFR0Iq9R
lyg7UDdm9Ej3F6qTVzRQeAhorAV20Pox7Rn2MZpKgLuBrkAWzWXWnzzjGlT61BbB
WuzqTixfMj61R6nhm9vAZyOXRYfOW8wuz3Cfb+Apf23AdojLpp/6oJmnwm3dHehc
OgeKLF6Pa+7D6V+ooSGUctPaS+gU1prQ2gLGoqG5OSMIWV1MCLjfqmI77qFoqnPy
RctXVZYhLxYtL034H0wjce1r5eR7zJ4MjgL/e1TMZBshd4KE6LPMJBEOtzlAz7n4
yNMDlAX2GT3piQzdkUKjfrYKE5j/Xe5ntXc/EloQC9zVPzR6kC1SC4hgkNj8gz6I
SyVQ3hUybllnZY974W2+cURt4fIt9Z3Nt4H81EEe9BWAXdjrUbhscaJt2mxWZ3pZ
4epuYKqrvAsVZANbKLEhIHPsybw0GxWiow9aYrCWTqkEPLPfYkiKEoqYiF86a4WA
IdIoxBKRGWGjm71G3inNGYJDQfhz+vo5Vfxp92qrUlSFHp8Idj5u4ZeMV4xut68B
s5VJsgou3+14Bf5cZekieFkeIHUGJYI3K3J3h0omgwq9i4qYYJ/yQ4uBr2PD++sf
/8L0uBMSR1GwmtKAYmCkstgCJY4VAyYclbJy62yDNz/RyAKlLBztf6CXNrxTpqIj
4/5Z5pS14fO8EsYKp32fSeefX+ZxhTmeHEpgpulRpebRcEKXl2NtEPgh1VO2L/ea
IyqnVGaZxK7Q2/CuMItcQLvJIwdqtf7aVesbYWqplwE18Ffj0RT+ddiVfCDC+Ju8
/K1/jt3JGjfzeHfLEilb3CQ6eLoiul+K6MAi3R5nsvyeitA8DPX2UOuTFtyrUo2q
93EICG6cAHIb+1y3yrpCaX96iVy/sstI/7pVYaSVhDZDUpmKxEw+MU+p+Pmv4ZtI
h+gj1QKtHIX6p/gF+4tPfgRYUsODRG+TtIETsDvKhY8x/VpJRsnpEwmjgKiskOTz
ShkI1N1KTRcm9U+/xdaE85flQ5Eo0UYFjnDQJT5sONQ59pAnPnyyY1hIuUXRGwPZ
9/1PRIkdadW6KyluhzTpDvj4hkfNEQrFPBhq2XhW5NiuSBytbSAX6PTME7tHyCB0
OjLrY0oQZOSVljyi07vyh+6xIlZInbVbN6/f3lCqImsEdK6cexWHj0xYbVlN3j8Q
IxoVyWm5kQ1RrgAjqo7y/XR1FobBo0V91aGuCiftrnkK248wVjK2Oc8tnPOB7gnd
o0O0GHgEPsGsD8rldMyykA+nADzs73MoSHyYMqH3tk2T4fDbs+umTBJo73fIy58M
OjpGd4ODLYrp/PKCuB2hItJ+eCwu04vrno1DVLSsqdxqQiALMFEplr/7C9TYTi4C
xrpKHZeoY0RhhZWtBje1OnQBxLqLxjP3Cl8d/JVVLuDIN2SQR9i07oe90nUr0W1L
QFHAnLbYrS/sy2MmzTKdIPklw2jbU/Nf/OuVg09WPe4ZtHMcohwwFHlWuM2oVfJ5
NqsBe97/z5nunuERza1TkYIb5bi+WawBgyRWKY//O7xSjtrHaZXENCuONMEiDT6i
z2ZJTpsrgTmehpDCUTmOLUd7CcnHatwhcP/AuuprQptJR63xMSWNFZ6STjy5d8S8
wCsCvqEr5eSOMXMxiuUMpbaaCYNn7BIHm1NQT+IapSkVBpPPWHspoIYNDxbS62D0
xH4KaCRCbks2y1HvTFlZ6xGdULmhnrLaNnbOdRtv1KRNNPYtEzqwNUUDlo2LZ4d7
JtwbGtfceb5WYvKI51azsyywt9IlB8OzFQBgWsVoA7ugv0OC931OB7GhwX+iXctQ
59q7WyiUBuGTSR/0fCa3Malq813IDwtmgBpp49zHkewvNYwPYQCeBn5+nIdSicpB
4U44YT1BqLTIshd6tozwc5S4xszBAQhzECzwHd6n5lrM8SRc9GzSAxR6nM1mNJGj
R5xxYV9p1fNCLhd+lUCBnSbv0YRfFGZKP+R1DtvKwRqimTjEmA3nIPrPsPkYL6QV
ieB21ERg7D6BDaSHAwQfrWxJXTzckVq+lakk+88hCq7treJajoWJpM2KvFeNIr2g
OsWrpLP2wxBz/AoX51qnhcTGKTssp7bhZ6JpqnMEld2zSRY5AWdvz9rpLVjn2GFt
hMmHOprRZnPhM/L8ZlxENrFsI046RQEZmA74zgZpoAv8uIii85AEsz4a5yBFcZhK
dZqOvTeTdAijgsQPXdm/hN7qlSg3nH145WgsM2pr6jZwV2+l1jG5/WcOPsA86XDI
QHaoSuEHKLwrm/T35hLnZ5AL8V4gRO3DsUpNBd34w6VDObe81DPehBXwnYL7kaDB
YNrM2qlvCdCGL1hmwas1ThDZUxdHhS5BbCV2UCWjLhgjRIKj9o5rQsy+e2LV79LF
UuUr9sGaTNydl8GQl7o1MBhLYh5zX5LhkYlMHqQELnZZ6VqG7j4kd1lTM7KNtr3Q
gIaeAa9dFb8A0k+qqnY2P+/9ky1t/+hA13mILIYosQuFmNdCHONi4fQNaLGR108O
nRTt172m5D/4Y8xZjXj8kQ0yTMHmXM516SkBbmXHj8taHm7S2rE+raDYzFS9phZ5
M/KQRR/4/6WmiNPCGVTDeaK+W8M0Cw73tUS3BfCrRNftQcRNM2twinOztk2QJcCA
dSj7TVlD8x/Tjt9BBr90gPAG34CQv608vJItRX1wG+oCnDzJXwxezr0I3TE2QySU
5IsGjnpPlU+j73xVMrzxINz+UX0oxIxI8f/9YeURMckFhmYIOui9QGIJo9ve+ciM
T+XpofzOiaolzUI8ij8ug5s7sHMI2gsa/I/IhAvRt6hz7yYECUnNxz8hTocOG4yl
jqCCHiEqNCNZCDV3b5b0Hskj+v9heg70TZtXZ8KCaYevjrKccNVJhYtvcIfZkm3s
1nKbgRPiTxULNpLd4YwDHmkL8GIWRIZTzBExHoQGl+fJM/PGCgkuOm1Dgl/PvgDt
AzYwM6d++TOWd77sEbIrJlv/rQgHrTz1dQtaoH1VAAkMHYMvkCBLqVy/KbJb2lS4
5b2gBk9oVvXKgKNey1PD6EN2I7AmhaVMgOoaigRdINxnflQQUarb8mppFWcGqJ8q
7LB07KT8etK9szaP9SkEahemgjVDDFrJ6X0h6Tpvcx1ImhCajasc0N9vyc1ZfK5g
y9WptFdsLyPsePrK+I5taii9NU7/NxvKsn/BBzv3gC/OdI0pjWTh0hzDbRDMJpiq
Lzop9YxqvV1m9mIpkHx6nHMxuM/QnPiPM7KFAD9yh/BKb0w3ib+6L03XbFtEOTgl
zwuFOTV3kFKmwJtb27WJ1ub5eNYkLgKUrTea8v0n8Hr2Jf2D3GnmlP4zF+KYv6u0
Xrtv3OF8z6/qa8OeQByNhcWJyAlKjWrme2+zaoGMAqLHcQaR1BHcxHUkfVXNqmy5
nRVsrLe+cUadr42BfPn01Uaa/Sqhn9vEhrbF5anCCT/oSjWnUclu7voxkThv70zy
vTncCmYOSlW4LoWFBYCgT+tYgxOYtBbvRdt8BpiitjcYIbE+XAj1nOyxxWkAnuC/
Ms9MmOg31Zd+jorf/EH8qAz6jrWotrAYXkZC9FM7dBfsGH9xBapHlj2OjCcuDgFu
2iATvTf+SUgSLkuMJQyuiqByc+OiKQ5Qc3xPzw2BvGB3q/OtpPcoTROp+FGMCaQi
1zLVJo4wy+ZF+WzhrSQQovzUnkjKK33odUFUJ+tbuHPRWN5KlRSO8l2C+x3vG+MG
+11aXztsbFslVYND7YvmstWoHoOcq9TMfU7QHxAomyJLMT2TVu3bmHQL5ThTtlxo
m0Uvs/W6pi67ZSYQcwcKAslMtvUV3PrV03kVECW4f5wpi2Vd1c1R3rIc7yyGkXo/
R31FyFdlafE7Ui/TmR6MGJSLdbGhsBQ+luhDyBjdlg4jLdCfmy3K7ma1NcM0OaOM
w0nzdPBWELqjixigpmDAMrQ3BlVWugkp84Z6T5n8/5h9sI0NeAV5I6N5meu65V1j
c1T3yl10juPEjvpe62MAD+39oeotQit1DpJROsfeekWVZQGnnZfmMECvt1Z5ypiy
rAlJJEkCrLmnC81QGtY1F8c1FMGkZ3n8rY8UIUlYgfppGMsme1OmrIcSkS0DA924
1tjjlOEG/k1Q088w/GI4c6vFgcbFjerPcqI5g4IOFWWVhpLXLcopu5LCIe2QFor+
1jSR5l12T5ZFEVQDTxhEuh9ct+1caz9+Ocq3Mk0xO3UzgMxxdcf+mGuGzAW6tz0B
z22PpM4gD+YhFtZyXelqCcG5NvU2JJ10syn3i2uljkjzfaEgt+7R1mFm7thMQclp
mJa7EqbLA4oK8ZQTNOhhigCyyevez71i6/Xkd9BcTuHLMQUAr4+mpRvkKqIlBVvB
21P+hcMO8sXijOL+8CeYpTR3IaYkcMUYlfLrCPcRcIaSW8XwTLIk/o3cA8vdpRm6
Px5UY9EO+b/e5z4uExoq1mO6ND/twY8uc6IUmdSmYxF0pq3NqAy0wwcKRAUVjW54
F266xkwUimW/0+CwID8LWzj3yeewMiUM7saNlmbRb/pxWMc5QoXYZrhLFmmeTTU8
8tQBjnlKZdmyonqcCBP2m8mtOdUFJpkCsJKS5KTa2QSlJ+Hx7dgzEQVsggeASGYD
HUiq1E61AXecI68/3fNGhwoWr+wLPq9P2dH9q7QZ9AoiRbcCJuz9aEhFom5SeQ55
FfzM+NHkGttCFjWqh9MIAPEUjYOHwo4uwyg8hB5ZthwnYXrxDjsft9tnLjtC45cA
gNnRx7EZN0M6lLTDEm6Oe7LyVD0wQ46R2BHZNEUEZ7Fr45G4UluhCaGyx1ixaS11
Flf1Oo3cftVRr3XzBYJZZdWh1duv78/iRJrNqbKRRAt89FjK7KYW4ZMoAL0F6qm4
1m8D/TRBygIfwVvhcyclAJIPHpjYW+lkJtrqs7rwLRad4Dm2tiqVpU6oHaEhHcKD
IONxKoCdlx/xrQCVqQ8LgnuGIUBueGsIC0lrxKSgwdwO3FHaADrJH0gPNMTp0WX3
RUkXVGNmnqGAHFFRVyCN3Sag4aR0Hebm2ksZOLM10+ucCaqxR8jmaaNY/Iqee5KM
O+yQ6L5V6mz5CMiFjs4brx/N65zltNIryDxh9GJSrOODe2HGU8rgzsqU7wKb5L2r
3jR7OIAFNUkl1VYI9n6orMWGoX1ODwAS2f5HmD+xTk8/YptvKnbR6TwyMgf+Zihx
sWnvGuxjmGUas4VSXbV5d2FjtmoFUCw9FWuxUKYTBtKThg2Ps2iHvBMYISsnm/2K
1CaZWsHJPDSW7WWQs4w8gkdj+gysJFzaFyZ5/xYXiZDBD2WAkVE/1cd4otwr60Ma
KR046StyUcIL4J8+cylq3R+QQcRIZggrFHkyl0iEpuAiOldKFHQi+r/AswbNff61
1KzWAKSofF5QZK2S39R/1Yyq2e61JM3uDvTlN3K1arpqi/r4cp2xtWvedgOC+E8k
nsO8ZrQV+zb/UAjCUSsKkKaqTAedNcwFROO6ZjY0TM5AjmtCxYpDBuxEajeElhfn
6hEXIaTen8V+Cen0XKz6LoSJJ24/6jvf2jH9yQAmSWi2jEoLvgLQf69i1vEcM2yo
Nran9lxwzl0e3kmoztCKoLAaFETBu2ZJhub+2MOg2+jb7L9uPBg9KSXWSBpwBUAh
OYbbNY+hJ1h4Rz2LZP9rKykP4tvNGABXtP2m8ruWYOc/qZqcfA/p/GhBF5RgLjo0
7PJKMLXbrMsMkAYKS1qjnu+VscOYlA1IZy1G5jAYWXFKlPnL5JeKn1UdjRePML+R
t2Ma1Z1grlaaTkvD0UmV3x7q/Fqp4q7vdZRo7zkxYcE+ecqcHdnOsO866fxTU4hL
kDl5uXQ68IfvZnZ7lY+o3vUg0kzvPg35AHrlSKtL2ORCe6FOzRwak9ByAtNQNQVz
LuQGyaRT8O+D1w5xtvUQAMohaviY19Gbusba3QdNS2I27PA+drPq0wU+m7OJeMQi
Lca6bdCJezMiDZvXbDSLFPdjWLNC01rnrZDcDQ+9LKk7/bX19Otx/DoIQbMcvoy4
3ZIPyVoWGicw/th7fjHNSpX1zY1zCWiCCUm6WFj0IS/KlR2IjSwa+9g2hu5IMEck
tIEQJqvYtHKyQNOzfCWRg/z7Dsuum6IMSQP9tlMQG65yTjTicCmGXfyPS9CpOK8p
+fBoow8ZGTGmq0OOw3aIcSjsCB+X1QxPPi/plwNAGU3nLCLbmvTG9VetuDkFv0VN
DSg+X5v6pt32a3kNeo55gRtOqPrkgYm3H7tn/qtcyCzDwq8aWBDsR9NmYRMxXpO+
DJjdPDofad86K59dIsLKuE77ThZRT6hzMw5yrl6iZtwx33uBOlyLnxokS4+SdBMz
LvuDpjN8b4UzP3Sn8P1BCLDwVrmasDHjOgpnrNtNFZWKKcQZK7Nib3o5VmWJYzGW
pLyLcbfxys38+MV/69ea6nbhVmPvpIWzD2fFY84qMYLZEK2o1dqlI1lkB2Xde/l3
koO0NSh/EZlCq6QXPsR1Nfw9JvOKr3pWTUSrdOtAUuUVrlsuk8nhznaS2QzDDCYY
MVN7km4pdlBLP1UiagSrkkcse4iN1lGZj69q5XwwmKSxpfaARJXcD43Tj57sPuqn
kJlKMQzeg87yQTYsf3rDXqJImKWT0OgMyqe3pxrDzQ1u+awFfmYv46Vd2zsX+i2l
5SHHKEzvIrX1as+J6XlV/vlwA+Z59/nTeWS6CWN1iKyN954GnGgIxuOmWzIehMvA
wDspNJeqJ/iNEpeAQSnrQQR92ZDmU9TQ7hCi9CIJEj4wX59CD5mLp0hgtvydMt7p
yhYvQh6yuqPFd5pUwZZ+SelOaQPgLbdPOeoMo445/Z81HA+cb8JCb3Br2RBws78a
SJCADVn7u9e5WljqQknZjC2a4uf/hVnkUXmsuMFAPXKU6x0PwotHnG1epJHBcguA
xF6xlNST1asXvHWSfAhMr2ubHbdA3EDsdq2WVsGURqJ7c0Kb4YKLvXXjVDuOGdrd
WmlEM92qSXsUDNEQxB37K2CdNns72VzAQQDKwnwmVPNkiqfNEEzchAmE98vyN9mL
48Q01uUA8RpoAjt8wNyFBfXDfETypxhmK0Pp2jasvYWxjXY6c4BgNZICaQrWPbCM
aqDOYubmM0OxuOmaP2YZMuqCyRZ3HL9d8RBQ7bH3MCbmnA4pvYE+KRMCP9Ag91DA
9BN77/kiOFZmSSvOJPSxSdQVffXsNIh4NlXED4M4iN7Nc9yb2bcceud5WvM//e/y
xGfaCg1Ueq/dfxLQq5QA2/ftm0N/GCja7RNj8QbzHJiRyH/4jib4JnwJJlBRwKkC
oV7MhRrwSNEqo5kkmpRHuYcVz5B+zYg5bkeDGOBTSfT2hIGeLSjGuYU8Ox3qE2QJ
wHHFbSz1bbel5+veoM7R9z9WZa+TljLcOZKGuqUdb0m4beUAXwou0OJCyvfzDE8Z
PIg9kMaRJn+S+y0h7ZTJ2/KnIZb+tRs8MXcD38XNkCPYnntzqJeXOLy8C1CHY1KZ
/Alk8mW+w4qJryR67bZxU07WHH7o55DqrzWmVpJLa/KL8T130HVMjBrwF1vXQE0e
frICk6CNJ/cz1tIfzasZFClGKyXa9FqhtZUUGlVlWggw1/x0T9KZhJIuyGVgySoD
Qyv9Q8/lK8z/KNCZUOtUwb0qlmDGy7S7+CaN0tdtLcmuCGhBv3eJQW9ZDdOXi0AW
M4CsNwEEhADtXNXZHjba1cSbfv/DqCMcpgufFhzr1q9pxI5jS/lSmtn5oGE8m/94
db+alaSS1N3Cb3eD26JIfbx+IDXLb/T+F1YnkWjTobJpyKoTqEMgIfgNXR3GqWi8
qe1ylJYPJ0Iit8HvMRbpEA9XAzbWgx1RINP/oe1Ktfdne7BDNBRI8i3uc0itxGjW
QGabBwk65vD27y59T+jzE/8uLSjbAFY8Vl+1Dg5eeBNmjPpGyBH4TwalAk5iXMDx
i4dRUbnXn7Wf1tn7gLFDiy879bBYbEfjAAVZwyH9PqNqMawKpQMdAx3xKYvoS1w9
irN4vlwPl+qAWySw1fHbEQlpqyxjKXgrHQooRvA8Bt0X+hnr1YviVHQvujWHy04w
Kswqsnnl+dmp504BKLJ/onB/XL96tAEgVFu0Koz2rdH7JWpF/gsbg6HgBYWTFcXa
uqZsjgXASFE6rInBBfEGC9MvDBOw3cRrHo34oH5fzrC2S1sZrVEUvaPnxkfjcNoa
0IvSCzYFapwG5lMMdG5omtKgnQ2s7Io7my8JUv+4/Crv8zESbYnENaEh48PIu4uN
KMi6uGvC34MvtMN/RbzJyNdIIvHsFeynTrprtVp02YZlG4yzxb0rjixJhqC+gFLf
CGCc/+t6RzuhcsTRwa8RhJJaS28NrnIKZ0dTlOn37PWHWRqnDqIeg9g+CYw0bjvT
ZTCYB2ptXWNh7oQywpnK1tDBtD829NVIbdZrV9t/cuR/xQ/Nu9Ld67+miI+Ioy6v
pAwTJSutjRkSMqzqXtf7rMDLj0MP+ecESqxjYzrgqIK/zX2wqfKBuI0jpzQT1b01
9PaNMOO03vKIuJn4+X9N1YNFuyGqt/kjmQHijcwBgGVvbQ3kmtDJ5HEiziYLl3wM
ctDlb/QdxgxbI5wtEJhb+Rga3rJCNVLavUHaWl5Vqu3vRvHNLZk9VjiMPVnRg/7z
WO6BcwGvM22eE49FfkPVVuBn+nDvks43W13GkrduI3dPZJzmghPkv+BYd0XEmU3h
+/yn7xCy4ffjqDbvNjWx+e9PIX2kvYC+xsu0cxvmuvRLhJn1zNNBaD7ZRE/PECZC
fXSbji6yqy7gbrCQaJoABI2yECd9fMvl/EmuZqI2oAjhd+Am+uCA9WksCUU1z4SB
C/VH9uLo/qVBcgpLeJmTjyfEmJa8EYnqXRYWBGmles2RlaArUbPsYi2JGv1NaJLl
2RGll+WpzYK/M0PgzlS8JodcpInEE5XGxB+i0tFhRDxdia/Rbo5g0/k1WIco0QJH
UylODrfF8cTHCUVn73VghcXeHa9/6F+upSeCWbvM6CulqQnn1LQBzzF0b9wXiDd1
kbFSJH8iSXG7HsKpGOEazzbNghJ2i4jDNoTsoJHHzvrFzbPDY2owFV4xbGccOSpG
yXzmUy1KBqpwnWDe58LgrncvSY6lXYEe1n75hleZS2oSB+gtmDbollYtXhdf2yLk
DgqBRlVZcEmgbu+02Tct2btuJEr2feSpd0lqlafPEIDyJxvGP3vGK8ESEmpQJOmB
lVOW3mITLmZyGaIbwv+FN+uwJgre9RiyaWYVh7LrzGO/MA2KIUM8xd9fd+El7QHt
XgSkzAwuQzYXBLIPZgVJJSiHQLNrpGWT9+Fn75A80giffgEvHlNaIQUxQvkYEy3O
ZAWzKZn1a+DbxO5RVWIZPLtxFMCIWvud542YjUgTUAr8QKphm/66AqrfRjtJo22J
xacaGkCIYxCNKYobQuZeF6cR67IuX2fjk8/wwTG3bP+R4AHEYnCdci/hgDj/82wP
buoCdM6N8sBn7LrvbNDCQn6/sYEkyAwIeUzhbUZEITzQ1+eBgcy83dOy3tXODZDy
Ar1v3yKpo5yFz4IL7cscwbSKL4Up4H/DwV2n9qk/cRVCDLgMkIxcRzkILj9ecgoy
y5SuSJkyfh9TwKquU95QjEACivFC98+XbdPuqZX2PVbcYIHXcyOsmFf9L504e2eV
iGM86A54JtVoj4jPchP5ls+W5nBQMHWFGzdXxMk83Dst/TvRQru7ksw3Cks4PVuw
1VupD0X26vjNjxI8UqAIsSxPKZk8XulSGPX6vFBDYzPXFMx/8hKwO+xV2LkOa4MI
SZDmb9AIhNebvixxuPo9uk3H74nl4mEUbXvimOYwW1pJ5dOwIdTyhEOKMxOqSP92
/iJjHkyxSzkvwWylQzOeyYgKFv7vhVePooANFQCTb0SngOXl6FLzmCmg2ZK5kqPa
erABD0IpdJZ+IRCfpYFpvgKdL6w4gpoa1OwFI0PGI1R9L/fS5O6v3LcvOvK1W0Zx
jAtmAMGNEN42ih4wUNfz/vZet124nqtmsdaZNq/M8xMbhcQanM7ognSbv1c3SKjl
bbbSfc33pCVK14uKsl1deu22aIu1aV9iGuB+sh7Xstit5OeyD5G9gFO7dRAR0lxP
RLecwq+PtQuifYm5CZuun+eNFJb/g2GToW/LeP/ilpAku9kLbhmbRgr9e0tYO/Wj
/QFKfe6TQv7hzwR2vT2YhM0c3+lPbv/oWIU2xDry9rTDcSr1h3txe+SGpFzYOtrE
b2l1uJa5cNe2HHezBi3GYwYgN+2jsk17zW3ukQN4isCG949+P/7eSiqkZcuWJWZH
1/aE7BT6WPl86kApxoZxTSJdjQ6upGbg7fFy0Fv7IMDyGhmO1g692vXheO/Qfv4C
OrKWGYuA3OBc5tEaef2F9EbEFbaY835qEr9kEoDeBruU1NI6ogWeqyHp0WWM6NdO
7kGpweInFCFYUSwsnuJIaJPKPIcAlW9VnUjS37HBM6d8xT0UcjZq3js2pGpTicpt
ePobatfzl+ChfAgplI9LElLAEsb/NuUuNIUUkX01IXaQLxpJhaTuVQDBbJ2ntvgL
ZtdllYwJ0aquUNfoScwCXtW3zNHMyiu9N51xEBSREErd8F5vaIiRprycmvMACfI2
QrFiUACfy0YRFett0hTv2uxZ5JbR4w56kfUipVbZwrGVz4oc1kbLBrQqeRlMrKLO
JXjnbEx/2nydKnQATnYdR/QBgrx7q8g7S3UH1vmzr+HXPUgjaybLXhfzCDAlVplH
JJ+mqXFBkCmGuFPQW3Nd94Jn/1T4OzlK18+Da72fCzfnIYSBPANfW49R8zROX/cW
LzobyI3nI+Nq9zlBBaJRJb0a4cZpIWZygU0ZQmnkesKdE0oO+vYwpDpxmMMfLwbL
RlUaycbT1eofM4po5x9kpRv1S04kZ+H/j3F1QW1Zl5wrz18i2Ncl6YT3uC2UV+iY
b9Scun458l6JS/78rxwnUE1GkHY+rGj6KwSCstZQmT6ofVdac4TugNQHUXiq0rAG
FEA+qU6wLf6FgP3p/4MHpfxIOjXp42nh7r/nz72gJyS7rbBaZQ6UUN8Sj32LKcMc
c9SXTeQcUH5t16jfLsBGm+anY8PlqfKCJ+mdE1J3CtGTPXPNxQVAC8xzMMz2AnUa
082DL7oyTMjWRAIrzHiPsMqMo+crISV+SlhCGB8IVVbS764lEP82ni6NG+sE35V9
CTCJ2KYK88EbqQfzkyvwR9fZkcQ+tkgEQ5yby66scSWC9Wwi9hIkfgmAunTweLiQ
CchhoIjhsA3zipaF+2VOqNX3Vmqz8HTEqt8WUyIS4I0Km4IBYaYoKOrOL4j4f7Of
xT78bihj40d2kXXduG/DngoQf5/Aia/+eQVxO4kHZLYbyzEpx5Zs9pOhvCuyxhj7
Oc3m2NoMO6nFJkR+rahYVtsWnIQxWpZqRJ3teM0IMlSC810ueuNZzmO9N+DzxFdL
rmFwn4/M3QjKzXNq5D7L/mvPKphV0z2uBnnk0bE4QrO8CdZbn74KGXCEdpZBFgCq
BVN/uL77wAn7OD1i/tykG11QFJZAXWZlc5gnKI93xZNlGlKCjNb6vVC+WK4Fgpj9
xi/+LSB3mMJ8IiFZo2fgbWmhSXKJYYT2bKY6oFeTVAPxE0zrHoyhTw/BV2k2mXSh
LbkO2teQiNIpkXK2Pk8ey53ygVut0XiplUSAUF3q53o+BcSfpcPtsKSolvDxvbsg
yG/qtMc9p8Kde9u0FmaYng8aRz/OboKJt1PY+7gC9Db/M1hrEMY97K+GLwX8c+3I
0gsE5vKlydd3qkf8BBxpIYEY607aWA0hW5q80itjc0L+MkRPkSS+v1t9H20IH+c8
Eiv4bcZtc2Tv54Wff/+yvvgVDy1uI1GdhPSf69iIxo/Oyt0q38Sfjcj19GKCFwsI
AHu0R0tCI8c8dse+yppmxrqcKZ0OprpeV0NpvblZpk+VqDnDIKzr/BM8GBH+u+MU
q8YVyhGe0VwQHQ9v3z06yWXQ82SDykl/GGSfFmianFqifQYEEGtRAibnQl9rAp6y
UAyE+30lbYEbVKny1DNrTB/5zcjO2YH5uPxVSCEgOIDosCYfrXZoC540HaTfubOq
0dHC42x7rW7N2/OzOXMQGRKevcS9ntaedyqrAVkYsyvCyXVYrL+wA1LBAhsN5V+V
YcQFrOsIna5SZTGnZu70DocULfgYG3TfQ46THt4nNFooqmoSf2pUZn+jUxx8f6I1
+dvvW9rOLUW97uwqLAhjhnj8rHWyfUPUBjO32ms016sXbBuqZavCpBF5iszYietv
HwZqlh+OdC5MzI7ialntFhrKYN65tf92bpKBAIruWi3Y1NbHEam/NIG2JBzJIx1q
XL+IHgTzQ82RnQ3kdOdyJIOC17AP7jvyAMtcbnx1/IpzBQvmJ4xPq3K6t1Lhp2eF
p3GGj2y/97V8X8lPVADg5UbUur5dsYGF/ZqsmUBILN2GwgC0VSLYjb4inHR4FbdO
fACkSg7A8v1WF6+UkiRWav3vU2+qM4KmTbwZwRAJglNxjQxNimx5YbGnPaAixQNQ
VjPP0whnvXNj3wXh7Tj1yzfOgg/xFDQYRMmO9MIvfEbGUPyimiDxpwx1N+Mcg4fO
kZG3s5Tl21YPhx61qpDSWv+5wHDzOB2Igq8DVGPeNcCmfQXaawBoZZY7LBCf5tJj
AGJpSthSqhdVMXnzySF0BxoLb7VWOaBQLoqqdiNP2TILmRKPM0eSmUDY5cXM7Kh3
RZROQDO3UjhrapghWzMAkyhD8qmaDdIEvvcD2MNvUzQ3YBLLNfl2eR3y7eswY1oz
iuX5dtyBkmjFfG4bok8EaBeKEjKbf2y1CIG/mkL7QP/o35MZwVq7r1RF87J+gntr
MVySAabsvpcEmVQW/fO97zfUfE3BtoFDlM0R2WPitFJXpyHkDWplnh4NxVlodIMS
EutHrp79TZmz2K5uW5NVWPSspNzdILd+X7a95CmY4KYNmIh6tK4dWDGTc2xB7dUV
FksbauSTqUoKS5jXRcwuyheyQ2DKg1KvIAe5x73QPQ9eUB+QAuuXHXxzIPyja9oq
J2H4dCigrGTrEFSb7wH4NOEQ1sCpdEcToX0sJ9DZkHMdTi5VP3uoxmuNf17WBcnl
N97Dpm0ZUV4lkIl3dSty6Dwlu83W/6AVkV8P2lUEIaZtx6ljbNbR7pMfnYYuBtb4
rxH/ZAblQoh0KfWVpcOlozdGz8q9mHwP6ZQ2FbOrLSppF5v9CjIo2eQtpcOq2Scl
uNczEqiq4ylwsxzMM107Yfzo6aQs4v/f/kRiN5Wuap+jBWDNwQlcwp9coa6inPGK
O0pYg2kjRHB2lc+cejYOaRhu3YlHcEV/ARVtF16Y/7XgtqvGBIPJB0gDiq0Wpnj6
4In5C/Nls2A6EXuOBg80Vp77lXGf4+yB6Q0aqCXsFx/mmas8VVeaIk5xS/aZfcrW
C25BOK4gkJi4K+g6Vb3eGXhq8orZaSac+GwWuLmB3yMCIRCwm7f9q7oiqUwLvw0w
cJLae6cHRHf1SPLGzPWcdC/FiZJfF+QD6mvHcBmbc/CH0Wjgelf3zteDqGjkaOyf
HZ9S45WIaV1UjhkcZKzpFpfPua586EN5fM5tKlD0NXnjb2xl74LuegcF/kcoGpQA
zwHO11IE+zg5gTtWgFaHUmwpyC2yRnAfxBy2kXFh/pVe5ugzdf1RITrRq7svefIN
teYFbg/TWd/1asLGNN+W7jHBKLOaXMPLJfg95nVtOMsBsrIOEEErG5PYqjN/Rj0J
IWsO3CDzdiMj3Dc8P/nT/VEDpExdALrRtiqmHUGWoJ+tyv0+vT1+xo8TimA/VtQb
g7Z8dr29u/7eFhFOCAB4BIONl64BmyfdrQEi6j0wC6hedgDk8pRyG5Hu5Oi/YoL9
yfwPKZ8tgx83oTkFS53sjh9tcCGkdljuJv8n/HIVHdLwaEmWEX7kJTe/3r3Opk29
4Qg8N/h30A1S++iL0oiBQuIK1B6Ml2pVCigPHhsrUpIj73H1prXs3oQGZgM5gUed
kqIC2HOVoSFYz9pkZpjLvR4lHLQDx8cpVa9vcOjF1GCF/2vApklH95BEwCf+zu8C
iO00FOtB3hEy9WZp0S5tHV5/8rAqxozY7tuxBdaXTDV9/WuYakwctM/9AyayS9u9
ubakJFw6HlDdZN0HoWMpZONiIBvDiTlr4qg2St6S6k0hX+NbVT2oBY7YHolw/gIQ
pg8MIb7Vqi5QpGg+XV5VDcjbFCHqM9MHPqeazx1T2hvRbI6QOuZ/Vl80xgsZJ2hx
Dl6xO5jocGUfsyiUfxg9nH6DXCmgZ/+1fdYC6Y7zE3xAkeWaBH+oddMSHER2MOG7
R/gZ9cGGeRoaKjMU8g0v2o6K978bzWpXdNXpVa7GfHv9/a7cfrM8XnP7Va+54NXs
ybyOv1ITg8qUP3Si5tDk5IQ26qqoHYxPR8mi/KfTUYcwLcD0wAEHr5x3OQHRCj9U
B3hR70befRTVk/DM7nulH5IbJabHC+GFGNFIFXv7H2GdHU3R5PykQDfXrzuHw8KG
+JYt+HH7Vmw0FWEwyDYNUMotIZgBshIV4CuXvfVOvhDswYy9L6Eui8BPLglHPduZ
tyFGSeygMZuJGEJ2kGY/EKk3f4ynIbZdTO4/Llm3HpkIzxLSQkNvJv8S4dkIXpKs
PN8PpaBKLhxaB2/Kafc+fhdIzsDab/cBGMFLOSI8Ej0xCzG+aGG/WtlSSrbDc1sQ
0nGeEKKXEEyWmK4NKrqN4+mVx3/fzga23af4ngwof986o16F/5jg3E1eCcMZ45th
8+TwbwFLMW+JwH+41fsDSeNdLKxg4ycgRKZnmPwQDL4SIl33VSo/4ydh2ZNVCJRe
5qLgZrGi9FMyg7U4peXal2/5ygDrgJc2/qQUxfU2a0dvl459gn02i0w2mTMMSt5E
pllHQsejwINDOi4XbMwCsmxIRD4lT5jsIVzLe/SU3Sm/xwqgifDQkq7h4AN/hTs5
2tAwkDXm3tv2cApBGuwhipkV0uXyIwXw1hns8VI2s+6gbo711ALrwcZlhmx0QJyZ
pw8WVsWphO69MZKd87Tjho0hd0oysNYfbXc3NRh+q2OnILhy/clOp6oQw3tI1C/t
WlH+7ei5o/Uz7TG8xEVqQIddEUw3Kq7nSpXvDrS5H3upsQ9gRcptGuTuWa3TtVxN
QwQ93M03/pJ8k+qjmGIO5Gl+vGPe9FFY1IYYnXGmeEb0FhJwVgfTaYjgIx8gPic0
3eeEj0sip3eGG0rN0XDhynUhD5W5G4aCxU4i6GhpC1yS10OiP9GDxfKmN57IIpO/
2BNj151s6M32TXi1JTP24LTci1bqLijjujl4oQdo3I5A95vEiEqtF6cjO1O847Tj
P7WeL2jgt5HK0ulZb/axbs2pLvbiBSFcfJRJNpCMMNKSVxLtWHdsMLwKB1C4Wai9
VCKHgBdumhQauAThQUd9lF9MpUMho9h6hIkG4Gayvy50Dx8TVepPx6lm8THo4QpJ
OQ4CncyzTCnLudjUNHjVKXPqzWhc9R/FAePVLZR7XbTTOHFNTo4RPJ87romfWKtl
OENc+G2IbTWo829hJ3PFbPdSYKtQY0QVTyHRgDcVZx+q5X1RAsp/NBlK2A64ZDzM
2bibYpoDupFzM6xQML0i3SmmM9evvghD170BEAeYoJuOy1gUuXIKebrt4ZYs90Jv
rQ4gHgrWq/oGUQg6oWhQkmr1KQRElxRgPovGwYiMISPy8+5LFwDoEnMJ9XQl5xg/
uZuY1de7dfdCtGT0lR0U1GUaVJm3mvXIO9Jby9N2zAziQVKb4iqo62GzFoqSbWsm
kUjOd4Ssl0/BAVzmfMX1BIs/91O6G9v6Kul1ZFfKWI+FJZ04uxjCTCIrfZH5iQgb
VzPNFYNNG/QgVmab5CFt9aSfxkNKuittCbCQdWhI1IBU2hlW6J8tE1gtzxIJFz9W
3UINRd+BwfisdZTqPMio7JXBFnxhbKE89+2HOs1VGkTiuM5PXXryKRazyE6lDmIU
nGPkyoLhs6e/n7rtXKJy5CoVIS2Os0wULtXa+jLbrC+zfbenPYWrwVbLcSmAAxmd
T6Sy2tmsp35Xf3CT7eGCq/S6CDetOId2hkTjHiJ+4rWxFVwDDL2KGlsGZ/Nkrwfy
1d0j21tQ+83X8J3zef0DNS0mvBAfWmmq9kfjXn36mmks0haeuHdlloXBkvCQ79n9
waH5xVBTJh/NTZka0jq4nQB5ljlVU/+/MEyusBjnES2MWtVrBiGe1vC+66Rq+j3/
SpkhIHrD6cGtKYA0HTUeanlBJ2nq7hLEJsdJmnjnFhTQ47aAWYx6B9Px/1x4sg8y
dBq09Gx1qkTtfBI4p9TeCqOKLMrlUJbD0s9fbKk/h85Wqw4lyNzvFxscYJzkufG7
SDrT60+pW7Wor9Zzak0DmHNfrHdvl/HRS+BNNKdsvwVw39ybt7OZIQbcIwoVOTh4
IhbJxImLo9h2dYkxgOpOETvm1NtwRCzJJoPHnR0kibIXpZwTQgmjPiFWHhkkIEjy
qk9qPtgUcKoHj4tkfmBoZVQtueFwPhIq00+TezTfjePtP4dpMfylndJjgs74LRRZ
cMKifEs1fMtIH+Sw52fsqmbb5VSvx7BqTECNU0fGoytLuAtI5/UbdwlWxeMYdQcO
pc0m2u68E1UCtLnPxpPd+n/fe7CojNCjoWiBS7nhssD+tGgVIbUT8Kzfc68sgQjq
LRDIJSk80st0DGcroY6N+76v1On5JfIbmlm/mT2nnYM/oVWh3VjH58LTA+5qGBWY
SKF4EYFWRGO7bm3HnJWe+haVHheLjRR632E7RuZazh5XrbbuWqQou4iJwDcI8ncY
OOFE4YF+nTUOHCOmQqVvI/u4oBQKb+A6Hjyq1v03IB/Q1bPTLb17OlGHEodtQsIa
neYVG3PqfMx7WTddScyacMCKE1dEplressicjifAScg6oh0nam01w1R2I2moiew5
Xp2lOq+eNFKf97BjctTfm6rCahn5tMHXIr9Ys+Ny22Tul6hiawz7hwzcs6Xt8Dox
sTfsgFgWnlMzpjkROsLeRJGbYrMBwlwxczGCTHJVqYJTEoYKIwAMYInLx8+8vbA2
S8y9MQ07k2Z/87AAICc+ijmmK41zKiDrFbW7Hghw4W21yDiKfKFWbLIqFpwbUGQo
ODUtAh/u4KlRR4mRHASn3YujNC6Hee+fV8bqShZHjViUOzqdlSuuL8DXAsmVUOjY
Q1r8T8gxJwZsS8nmN8Qv5YdNYDY678FsulLY58S/o1EXCJh7r0YzKGqCn1XafLo8
0SVaaMnIg7Lnu/Zc8NnkLMzWDzRZi/ptokExhFfgrh3OXrI0zuZODZ+65e1J8UsA
ApFHoVLMmQOc7/B1MXKnlsx51RsCujth7iWPUHd7qC1hi514RiLw7e0u/7nChStV
eNjtMKmRHLoO45EjQPUN6yUypCH4r1rGyo6OJQ3UdZnf/zr+4mwFOE/sPD9ewHhd
bs0IFtdaNcweEPkof9I/7TEBuPjWn40rVxm7Q56z1s+170h9PIv05+6o2HWRcxwT
uuezmR3yLMfMZiK8ghWWgwWnAhUIcv3RcTSOLCAyNLghtVGV+FjHZXDP3n61f3EB
6eui211h21bwlgCnLUXea9sbFlAFE17aJjDVS5ELZOqqHqI6dTWPlgRWQzFT+tRa
o/7XmjtxJ+w1UKg/CQcG2+aSnRhoD2sB7we+fSslEqngfrWP4HUTOwvD0aKenum+
2h+cDgAE+UOORUikgeZzFPXPXG3vdxm+yrDLHH4TDC3xlyt2bbpyNXZ3IqJ9gDKl
svEkOetcuxXINjhg2JQBx69fZ/m2gcCEYHGtv3oto/XOhIN9mPr2BufAx476xkQZ
d+aWu/CPZVpZB3YdsYdmQRDX0DWyWTuib8dcTjp/7W0DRzJezaowxSS3OqXXRJK2
hbYzp1ohVoqRJDWPnrxKUhbMitm1qntCaFp6KHWt+EC5S5Bl2dsc7Me4r8M7QpMq
DksPedjNi2sa0yJ2+SAPu7yn/hjYN1pju5yvN4iIgxDMNVTwOONMA/BQHig2Bt4t
rMut3t0lC76efNSyhotJlG1wwlMef1f5yKgeAMtmjDUBOaL7FY2dqI9Nfv1ywiV1
g8PWb+MAWfUg8EMBEBjOfvXTrK5F4lDXcm0k42EvwAA2ef+iFP+5U5hzdeFS6bd6
2+qqMq9qHUFJhjV3myKeZ3hYD+ma28M+0+crlaFABzIixZkGKn3h5VIwZHc8xbqR
bfZ3UiEcn5doEZ3vKaHrURFNnuf7xXY++QrYGPKBDb+OdU8Fjv4mXp5x+1VOZqql
kQjYb00IkYIEyl+8moO7GX75spFVLhk3MdI1M0GA0f8SBQG0/F8hIrjSRzynyDZu
Uw2BKzmEAczn43QEDKd+SN1wopn+uf5jyyNa9o1+ekkvEunLR+rjoBYZYmZdfn6P
spYgk9VFAVqtn4fy311/YlAXCnL8ksm1dgz8V+yNapAjzhzkNsVs5mOY6QE/RdiR
guSxG1//Zo0ODRi9k8blCbQg6KsB2FlERyvifeweAQxP5ecpfCRX7MRlsVXrI+Rw
uOfVszTTXcfkt6KQc4zN7EmTRrEmRVOEOweUsmUSg6d4ew9e6pXWKdScFHcuJgpC
jMYdCNqBuEqsv3V5beyeWCWpYKeU8bvufRxI8+XRe8FjpY/KtrPy9T95GA5bznf/
ZDBpPEzAE3ygy8P3HlxVsCZLnkBXQgfeYmaC9VKu/82H5aQzOjBwdz+n6xET+9xw
klB2Au6Ad883W9lL6TTZvvz5fuQ6LXmOPCuU/S5ZAwHB3afBthy1X8g+Ne0fe04b
Utor/AGrYeV1Cj8KAgco1C30hrEaQWuLMWmJmkx0ZOGAo3Bf71bB56AWZub75hDC
l5Md0ssLi/fw6OpcFqjPQPAuvx6HhaY6+LbRt2kgpenYy7A3d98nFXQGxH21Jl8m
GRkLXwe8SX1cWYNNn6rAdUdnCwlE+xJ4JVKnKuPs5aYvfYEz32KRC6WIOtkpNWzW
Bt+S0yWjPH5R0v5ZCcmoSP/MYG6UBvI4EBlUFsgueimx/GkALJWdUPynFIg4PxH6
aFIX3wfdRpcq1vUL6cjtnTuBUBb1YXyBYiMG/bt4vmx5+l8uM5ZsKSfUU8AlNLA/
4oe4RrNtHjTgpsgtMgE/6VdqIgvVDmWTotg90OevYRoTJ9npL4NrABtWVTKNCmpa
z5eTqZ3O/w6NQQq+tk5+zQnUW291dAUZz1xKdjzmD/zifV5MwzDzDCqLSROy4rrC
QKsWL5mX4DxsMeN5Fo22t8syuyd1bY12qwx/7RD7wZ7wl5Go9YyPbLE9bxUf8jUE
AajdCQ7RjULq5iIuutLfxoQpeH8U8qiBcQr4h9mCf3bfSix0cvzDYnyO09kG9jna
cPSijOEVkuQHTi35Ks9WplkV9y8JbWq8HjG6MP4FFk9hE0nFElOJhC/je7z+z4de
RNNWDAzk+ZKCU4NIzuLdIaKpyQ2+pFpE606+S5lHQvXuzkZJrGcx1WXhurLpnBFQ
grUAYLsRGfUCcsVyehONf+PSktqW1J5uknSJjQ9H34uDyh2s4Y26NSpPT5JDPBMk
pD1FcsqQqBOPK6pji2j9bAuaP+mCk4fV+75kILnFEWwUHHfUi5xNtaZ0nS7p05yC
juJImkDbBi4vYHlVN1vVvdiKvpfAdolHE5qUFXzY9NUX8QRFlAUXA/rsAiO8TRyU
u2O08yBDM5xl+CcSWw89EPHjI4GRdRBrj30wrya1DafhtlT1zB8IOaidR7Gs0O5M
MzdGMw6Rmm0xXmhdZTM8WdsCa1xcz9iadI7s99nwLrRLJletbAv6BgRVo9VJuSRq
jzVVub4D0cADpYTCeJ0GzviFaNxlnYmz45YOGLjGNHIh7geqzzhwCCeTZI7BJzQ8
MsimOxADNuTl+jRGFgzjZhk2PYeP4up4Z1cCiKWubTxm3HA8/l4t8VW4HNfC5GXg
uFu8AnsTg+QdqvRVTkXWWt+cu1JWVm7XtKhsTCjETz8yly7jqEz+Hgc4/eBaMbWD
2ICzkQpqys/uoz2/fWywSMO+2CTqcGnPLlzxBLU9PDZQYCUn8ORCOM4bZcZgBYF2
HVTARUHtXeBMetnSyWJjdrl6kaQ1j4DScvMyGSxZ6JE7/+LisWA9rhQGpz0gyDn3
uci+Vfd8wrf2jLVGQua72RZRd9yjbeM+mS2wCfK8/JTZ4vLZ2trXYDQN6Sc5Gr3p
UZ8uznpsBIoZ0eT7/lGaxiA6eiexbRW8nJ0e1ChNSV87h6Fiju46a2/uTTdnCYWf
1Assx95JXq9glGQViDEyv0vZ0AsF6gkUzuxVtEO5j1E7/e8uiCKdKv2QgKKIWNUq
KTJal6ZQl9X+lDSBFqNTsi5Rv6evobS2I9GtlS0uNHoy+qFVojL+um4EQX2NqAAL
eDmwiEdtwKxZTddFUEVv48GK6jtATnPIDMnS785SkAJ0qcJTBmXT2Q5Q6pE5qGZN
Jlfq5oTg+E5VMFrmxf1kGw9KhgPiWLn3RSaayO4NQ1BQnpBlaHSPTpLeRAerIQQ8
8DtQEc4FHHlx7K45iMzgHZiPLg9n+vU0s5uRQJt862y+nbxnWNDDvzpBzMDIZlpI
`protect END_PROTECTED
