`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/xPRmHOav+0DWlVtMgFYnkSXJkiGaJm7BQv2b96Ft24XwtjK8Vu2V6S7+K791Kay
aldUzgNHgEpM53rDMqpBQXyC5d9/WBFjAY6cDWLwLsaHTBegghr9s3f/jPdf/Hwn
wGyOp/cxlvgJJeUFff9SqQ2I9qSs5njAREZuL6Zp1px4/gu44ESRGTGcGZHvUTUm
ziYVy62D0jIORCCA7nUICEuTYSyQ2WTrnDmTfoWvZI6CdhwXw9vjc2zSvu4OAzfG
c3c0CRd3/OyDDF3PzRF4xepG+jHY2IakQdNhKLf/9sjAi3ElLWlNiQxEsFnQMOAL
snu9ykFqhRr05YEIhT2DNgDg6BUvBvv3opMp2i0ZrZKTOYSD3ZPRK70NVEK9GpW/
Ju/VGesnpNNNwHJyG38/cihtyqrh6tsNmsMCzaS4zugCT0QrtOgfQOPOD+3i5bX0
cwLd4UbvFtPUyeKHTlPCKSmExom2R4qCJ3SIdDrf7rckC5MLtuF2LglgbOCKx+s/
jetnE1BSHeMRkNDvaHioG0rDAPVIn2uRnWPlvEgJ6El9qbH5ekliiIWLKPm8tgal
4MB+IIW7d6sVQxuUJ/po8xMFp8FkQBJcUPDVTIRGcbLRWMjFIwCuFNMinauyg0mR
22x1fYdn32jTbqekyP8kI1dFrhBk3IeOZl9W7V9rjq1TrIpZ3Io27xSSazVsQ4wS
1og09Obis4LjDHBrAaMNhGVfwD/Pe0qwWDGhMmaQxV8QX9t9O5Egd5CqVIv/4egD
5ZoQ6NtdRApsQJ/oPEkx+AUenVK1C3UyHWyTmQjtKjOg0Dwvvx+WZ6FYfam/P+B5
`protect END_PROTECTED
