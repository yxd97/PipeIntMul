`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8T+BSw3vVi0wte3KaZUzggAr6LgXZqoWDSXCBri8Dl+DiC3VEowlx+5pcKGoYDLk
qbgyvoIPyeOvd1j/Sxh4ciuqcJJpZvbULrg2t9KtnpC90yNBWstYPlQ/BrycjWVP
qh5WdP3ig8ppmEsZdwjzPQG4pO5+ebcTAnn34QVecaav7+LJujI7tNqfWWmodLja
ChovtfwJv5B3qHe/jGTHggPBmWNQUBHa7qSnOXAtVqu1zbtSgxcinl9sSfRCs1Pg
TsAtz1HTxhQ5y9ddorW6b0uauqfGCbpM5ZZp730hQvsWcDy1r4XgukZY3zCps37z
eTNnRxM/3BjzGrtPq8Ib0M4Lh7xfgDFioLIDHlxuvvKNDpx6E4mHeUPdLoIx6w7O
RSgVx34e1n6bZj85GYoEcFPAtRABBiu4eTp7m+gZMrCFMUhKUZkiiioM/jB8JonQ
hE8ilR3/R+nnZja4GFk+Wcj9G2Cl52nK0/V560E/ac/hxx4x3zjpjd+n1XVYb/JR
`protect END_PROTECTED
