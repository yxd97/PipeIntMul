`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QmbnEnLiopowix39rN2E0aKrRzkgbOqYptAI7hEDyypH67syF1X9iLNFT+/zpgzH
2bWBPH/6zK54WOjEgl2Gc/6KvRqqA9CNt9gl8eEFoU+iO9NTq2zKT52Jsy5Zk5E1
U9AZRtFL0zbW01GIArMrlOL2dkU1NPPfCcEmt8g6LTiJ0F+9C62Q1CTFwSvYg9wz
OyL6kpNVqrH8l/99YlXDU6jAi+q756lZq9inPsq82kuuNQogVt5SbMNcG6+3nB9V
SK9KbepX2Rhg94jyj/tJFFrNR4cJqmXtdIPrajvl02xbBGWQG9KCHkbXLYIWIHTX
8I2RfNIWSYmakNYVYhRnEwsG+sGepHzrbAU2QzUD1InGdwBlKfrEh7kRVUBeZPIJ
JgfazKDMt/prmCH3vXXbzrOYmGGPiRT53BkkkX0CyymjeWXJslRJQtFBqlxDENJ/
XikA1/9x9a5aDzqieNDkCQrE4MsXySmSHkPjlhqhrDlYW9zKP+rUI194ZbILxcdA
+HK9F2gutxUukL++9fb24JOwYyw3Jq8GR26k/NM1vlY5P9n9TxCFVY2XrtkccM/k
C74Uzft2sOLaumL2RXycBg==
`protect END_PROTECTED
