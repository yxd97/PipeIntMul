`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XhJZVvWjbqoA8vNw61A+KE5OY4yGkGOwMIzeKZW/Zo5Y7OeJTVSv8fYzlv5nq/Ef
lMh1RlkBNlIjeOGBubX/3P8y/YNSMutNsqJ4ogXFEygEDjnfW358rIJab3G6Z/jh
pbEK8vtGXREjTfeV1+HKOPjdyne9kE1KmHwAadXHEdosqGhF2tm2SI19OYy6bR0l
GWLKFe/6XrkoPL8ZF5q7/paUTGtd82vqjyWSD6tRpi/LfnO2V5L0/CBxPw7v8bNj
`protect END_PROTECTED
