`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E0UWTkR8vkGoe/Sz/lBXwXXirGPb8X1s/l1DLMGk/jCb8kQgkizoNilvdAVTJVgj
O6PbpfkPRXldhvodwE4+xgTzh2gkLd1TFB5z7t7kA2YKxS/YBQQysO0Oc5FqWv8i
zDKaS3Q7M6HsIN+t8DZSU0b8Wxm38zU63P9UkusAuKCYUYGSKy3zuN3mrdT467jZ
hHlia4jSNMsicBkDoYpHW5TWanzivxKYNhbUCUrKLzfK7HEd7csy+cOALrNImAzJ
wdV1LFVNZS5ervVX7undM4b2g+m1mJ2NqDDS6hSr7s7zO69CZUzMg14XIvyMC3fd
`protect END_PROTECTED
