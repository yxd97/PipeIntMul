`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dlrInBbhNYwSI6NkylL9cS8SchTfkATlEtSA75WXBZl0YUm7Jwy6VovHZKCkbDSB
+LfCyIcAEkqUZ4txhCTnG482lgtFj9I2ESGsPuQm1LIpRaY/E38XUIBAW2rJ+g7S
KaoBmZgiCx6TVe2PwAgLhweFUCjtWKOVEOg17p+jvmjbh0F2ADimiNg+6sf3VO67
lnIdwb63o6juPCRN5Xu/4C5WPG3oHKko7uOEnK3bsxreuVH3obeAtkXJzeA7bYdF
ESbTCsmbcXmbab9a/Ko3Jro3YlY5ieMLMyXVfSCEzsC1pYrvz7su86zQGmPVR7hm
rxnhl83XIzmzQS73N93ejGZ1r7Xw8d3Cj7ZOO0WoMniDgeHcbyv9rnbntMhJOqo9
ortAPPTQFaXNG/Lp5guXrOtLLUe9HMfvh59/d4lfbasdPpePGN6Ua1I9dpIzGBnu
JYYezppF5fCj/4qeoGTivGBVtC5UzSaRJijUlnQRmV7MWntWMWWEu23lmxfocUfL
9d34lCyQNOpxIDF2y6nhrEj6Zd8sYS1xga0gfCyMx7MkalIHS8B0ccBSB5P+nvaM
ltlsR14LWNVoyypkSL8N4cddNqEPM7io7mNNOJuKBmVVBgQ6he8em+6EIKlGlAju
oYrcywZ6qg0CT9FsINStp4ih2+9g9vCDfc1zXDvfzwt4YAsfT0uJrxeRDXW6ws0B
Czw44BI8+xidFjvUUSyD7ooeln44jhNWs6ZNRNhOYXPwSuAaG8dqbPfSGoLU7lKf
Tb7L7e6RZ8nL6n3vsJ8JdE6CElfr9GHJICbC+4XPyNeUoYrQfqp2PjfO1rm/Flpa
ToGamwh2x1POlBRCAitVzIXoPZT0nFy+hC2b234Iw3tUQpHK/QCoSnJuSJqBfK+s
oGWEfV2kkT8gmKpcmziyBKUU5LY7IbqV5V2w1nQ7PLMtY/FRxo4nmV9QCjBA0CNa
TE4BUr+8inKYdA585j2ZYg46HlKMf9Rf3l1IrNWN5+Lahv+ZQyUd4ae17M+YfRLy
Qn2fJFpgUcmqY7W6Rr0y/WmHpQdgC+ENI51U5Bb5wcxmWX5p5tXZEkjbmKcSeJDk
UMOJ+u/BXyTD7b+ZcS2x2VNUh+b5z7djwlk623G7YY/TdUuwWmUDF7bvA/eYYhA2
d8QSExoVa7zFZkDjEbtlat01643pMrAQ+l9q5mPv9kwnabzVlfv8OzZUaiOMwglK
ydw0E66C6QggiPFHqdOnUAxScSYB8+kGb1xUWS3WCjksN6G1cX+4Cbitjnp999ol
7f7rFjfTHl45cFjeddruolq85RDQZW0QzzI6USVJroSfVDq20AbVfIrla+P/bmTY
yp3cPgz5KY31F/79fkOT/rzGe9S1WhZTDMLhHMtrkMCJyU7RvxD9Hj1DWaKm1pNh
834wGZkdvViXMjqjTws4i4gO5aIgL00n09XVBbgOCxsezh3r4ewR+kn4CByzkcBT
TOww+kciHU7919tngfXigb+vcEvydK1lO8ZPLZwGKNakZn19ZyPqcH3PTKwjd8Bm
dtHGQegCA3iJPAVLrvPBfKApz/MCp21EhjVUOdqEOtgrvzzJJb2VoCsaiW5s41RZ
SqoO0KdyALKOJshv1yzUwMxxIGD8W1M47qN1x6JNT/Z0ezroKGNZBPetghB2uWhy
85YtUA8MvdE7sQQdJhZqLhhRrvdnh8DNf8Sa2QqWYqWgqaVl9yxfz+yDlpUpCPFL
BY4WGyu25XpojGYgvziFGlzC4c32Ds0CHRO3G9yETkJV+xwQuaVMKHfKDsp2CykN
9hRKflyF0f8C1kfjUjKhWBaUdEeo1eCT3h7Q/oH0dl0QAdCsylt4HOoZa9SHQcAU
WoMCDm2Ud37+75aMrZiHdPh7Ak/M1ey6qPc3OrFrna4R8P7hSYQ5devWdqqvX+ZE
dZvwK5s3GJktSbOuVEwFWHg+MTnkw/Rb1etOty9+oRBwRtwMva3LoSHH0iiZ6K/W
s4j827bGQSFcTv3APV/T5ZmR9BjF0iLrhpP0QOqp2PX7QBeNSQf1MmXw04eflnDW
LW/iu5l4JjWhKYTljQ56P6j6RcxmKOHvCc93yJbH/hMbYImVYwbbwVtWBjH9Fvf/
ZQzvJ00kYQYp+0nSk9sGjrFIfYoFIBykBsP+uW3Emwh1ma+i5+wuALZuNQJ6hUCc
19nUFxryW61szTYRvQkcJC5hv2TFCVW6/Ca7SSwmkvE+rHlOv0RnNTKGPlUN2PaL
a3X2IgvwpgvYb4zuG1HOfyqFGSae3Sjm2NUkHOCaetVq37Jg4mi6AlXNIp/HkyW2
VuirECCa4lXbUgybWLMnL1Ntn492lQUtyRMeWBh+YlLj2ce+ZMizjXoXCmAZBVj7
JgtQMkk513ZzvvAd3ge/VFaJTIKdHqonwPdzcK1VOsogOfeC/6OeR//iEqxPotbp
+jFrcBW8DEWmHPZGiZWlhmKnX4zjEmGdAPEm8jO+gFykFAKPi7gcR6OiFol8H+zy
kQSvycLp23gRmh4j5gbje0TubZ2jRBrZSRdyAvum1oGTq3EROCR1Uv/SAunysxTk
0LzxYr3S8U7Q+l9/e6RIm8uAS11W4TCXoYcWukcuwUZQmmy2NxWOI22kKc9jTCva
LZ+XpKoS5jQBE57+4EqqvDi0J02D1Y7PM3KAI4WxxBUQ2FJcT2aC05dsj0m3Z9sO
+/YWxejh9fQ6W07LLBjRYeO+1pS5ebNLhbu6pV/l1fPpDswF4TqbbRx0OI/lXJE7
WvHWj5YALv7BMtIvXiHZDg8JWso/4gT4gYpkGbqY9gAGhA7b+z1juHYvBjVZfUWE
4pofm1qJhNY3vZRRXInu6uiD6yojHVLB7xA99WaKqbM8xE/uuIuq2IDHgL5Diawm
z+PdUO87WQwXbJsGagzqOVAnbZsJLPGCaZ1wYKZielctkcEOBgKWsNgpFKmDrc6T
7ZtyNGfl2HuUmiSALnfYTsrpfCJ9FDJuR1673/BzAuwehVQUipiiK6Skb7t8r7id
cYMWeGwRzNIsDH3AjtBqmxSdZvCWjHOHA0jalmgSzYQJSJ/admIgf7web7KHifkP
c8fkrvE04KpnObvQNKpmnMh1ogWIlqbWgJJm2IUppXaBsfKWuUBrpycF+LhRGYZR
Q8QQTfNpQkKwXDniwWNR0pmmZJPXX+c1Q7dup2hI0X86Cym65otimEM4N5MkmVWK
RUoDm6U6NhD3qhzAUuCQUtTbVw+vOTTDLlxaTwhJ60ul96rtJUhHoHmERJ8fyB7t
kxRs3LlYqxNgIlUDiTPu6I6pbHpfp9vLVvyQxTwgwZhU1ewzXQ7/0hxuavNH5h12
J3NtBWyEbV0S53hhXs+lKxyxdbOPPbRQjuBybcI5rmrAD5cHSbCNX4cMFcYyUueV
rHriaTp0VjQt9jrQu+wBpqwfWRO+obOsZA36e6kGAwZxS8WWu3RYLbJjvN59TiBU
MUQR/NZ+OqVL/Z6GcdqO9TEn5yQpHL/vICVM7uwaca430WrogT7HpgTyeVID6UrV
qi0eSHkTpB6Ank4jOST7RQ8AGziPj0DzNDgMIoCppfBk/8j1JM7fDrf0CAXnXDC1
DYAU9Bczb4LMvFM4BVlZCyoTYSZMJUyrxK304dzcSePaiKmw5IR/oWBKJV4wFQ2P
8ebbwyI7u0rytCrA0yT+U6+KDoj7EmO/wobY8fjhDvaDZle0xqP4UQmyPu8Qokju
TtnK4KI4GDACSjmeYD95GANJ/3whKCviOH7o6fHY9k9iKSYdR4K1j87F4YT4FlXD
zDOUI8WBiGqaAdNLSvemgGqaiTxsAViXqcx6HNxuWLRU6gZkdUX6ImGsOFf3JgD1
VaJ0k4F6Sq41e/WeoyAWA5GNWjK2ujDy1aCtgtpLd/IjwQq/PNcHRenP9uH0HCAH
wHRs4r/8JrI522skVaz1nQgkOdA/RBEh6qT0NwQmCcH+JfNqUfrSZWhuuVAAUJX4
s+CECoMN+FW+doJz0mpYfB1bCsCdr6MIVmVOh5NggVCl6CF8xihSF7/A0/hSLe0Z
sXtZ2/qxgoK8M53IT5thdqSLgmpaMXdseHVf4jfWFi3xntjdkHQS5uUqEFu0yIRO
Cjz/5sVWUlWcfBweofo+RiPv77SnWYCByGWirn1+HjgIQHps06mv6n/9qgkTitJa
i9CiFNK0nhzlZU5CQjJPpQ==
`protect END_PROTECTED
