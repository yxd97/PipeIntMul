`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JJ3lt9FuiiE8yoo9lEnYkbs9LIklItA0jOyBJSfS8bEb7VS3IDA8vVHUMg1fYZOR
1CU9MnOPSntFBIUZfZ3o87VTpuVnv2LzetToEZFSJeDnsHizE4WZOy8mVBbi6TJE
/5dSVNNH95Cl4agbtmmMFc752ciUTWEskXr8gDtV8lRYuStFpj/HEn0CdD6HiO0E
ogVTAn7nmVTQqj1JfuzZoNv9yYdVu3dYzrFIichgtC9roMxzek42s+DtPJmV+tc2
WDjzgqyEbkwM8laziHDbEJDjtzPC76sIO0sO08do9HSZt/WSy+Xro07k3qqFzedv
gzDb7cA1UZRbM3cViyIeJgLQayCMDHLnxB2UvV+VGaYksEJk6BzLZYWPWq7NKEcE
bCzCw0aFPTSYJaNMYSX0Q/2M6U71ldySU0mrIXCPB1v125+lyX2oz+f+GgvaYgHM
xtterONoEP81eZJWIDBQTD6htnHEF7UzYxOeAGmzSJCmXNEil6WqOHV4aB+NNKr4
olfmL0Px9shrdCTwvAo0Dk7Q8FKUih0jEdR2FJB8SnVTLzDByYHOg0fo0Bmd6Lue
GrH1vhFuRHNJXZTJKcrvYr0xBL/bQVtUlKKjIYOUFtbpEW/YSSXoyRZAXhcpvn58
Oxn/BIonETyj8MNKAJrYOxgfg6jAB/DEFyfkp+VwDng=
`protect END_PROTECTED
