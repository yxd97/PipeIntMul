`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8BdvAfUJ2IqQun76B5rDh36hdwiT6XB6JYxrT/JUqSaSRdVXEus7BcUL3auyDtUG
e/wH2iYR6dy9h9vW37p5DKQqb43+yTkmBUMhW9+bnhv9KqWHM6c6pud8nbQ5yJ6t
I2rS7cgUWee3azP43JyPcnvTjN6ZBWrwXN3GesqdCbIp2eAuhM5UHpDSYnkOiRAU
We22iojqTPtw6kRo9kjs5hRb5al3LNPbP2bMLlkZVQFxqtHI7/GRJlJm6cZCd4gM
Wnl65VLhsgaaiORAxISl/HtYpZYNDspF5yvN2IMr7x2PVpqn55aRAXP/zR7I1kTd
kSKzXJr+yYW9T1r3UzOjB/qH7iwg/LPRpRbdvuK57K0aNJ9JFP0OeH3TYAEobUZu
Da6gc3D6PxKbiFQyp8WESPQx22g+exg1mh22RSK32nh9Zj63P8HkKUpMm8LiJQIY
0qvMs1tOZE+DEDgRHLiTCB8L4YVhufnKruE85wrIK/7AjRTrQRfhL2fodeEBXvLr
66r9GFdXt9pQ6ITRdvMt7sOBJnFHrWnnhE7Ng6BS+00ihZ1lvVt9Fue1DhoLji4n
/IhE2/0RPzfg+2OwHtmIgu12YOf/Zf6Dlhw672SxUjPzYklLMVPOLexIqUZS8F0g
FyJJ37n6AcymHKLDu797vJKC/knn4Ap16iH2Dz7n+glSeMEgotWmiVoWqXvkkhhi
LNIiPTfzkwCMR1FrrSICxgc20Ip8IE9W7kxxRMbl6JdFpU2WQpFiOiPiU+OPObVh
A85j4AZPMr9pA5Mp5i6EXUQvBjxs+xztycwjxtKzb7AJcgxGDpyKElZu3Dbuhr73
yyJ+shPOnGKRIi6isPCg0EBErg14gnfV+S0EiEDWNevlmecHpvuGOwYutvAcCxwp
ZLHTSeEw9yn3k+mt8oL7SMguDD7a5tCnTvmzk2PQPKjhPLcJmWp29KK9OGzJ4Pga
WcWI2bf1RC6D4vWVz2VBybc0hZEBHDOTOTpn2Wvy526GayZo0P3zpbRXBY7LWDLt
PE784M0Qyf9tTSl0RjYe8eKL6rUmU3o0JP2r8S4ya2B7aDxdhSyjoVw32F9GMlAo
VkfGpGPcECGMD9uq6LMlOrV84ShcVNdRxgAOvsKLUQ8ljo82zMsm5fcc8csjtnRt
lz7MvmgUxNOYAu4HwAOTjnGfV0IVUY+bO9/6Wxa34ZmoSkPm15DdXM2yIl7Etb9t
v0Q8mqdwdIXtIueJ0eQk0cLfjuBGxYfZ8CowSZMuZhRQJOkggzZA3MBYbyVCUvFX
41yB7o8KBD6oodoBkl7XukDhZ1TrDBMZkFeY1UBLmflMLTR70dQe+qWVb2nrs/2Z
DEXxXIPODi+eGezHZYLqU9fZZimqiLKjHB+LQLeBTquLdBpeBdXuGkNgOs5rPdjf
FWHypvzvJ/0E4W2+xk0zMyUQDoO9/nreEqyznUvLWTgwUbFIF7WBHhgOg6wQhfMN
59h9u++nw0bv94AMi5HiDqbac10JX2IhMq49aojC3fZ1LnvoM2aSNNxXVmcN7ooC
fYaOCBCItJzzNpuf8PHvKMiS15bwEW/27+xf5e+FK6LTaLkK1+w+v/Mk1r1FDyi8
s4EtTHmWW48AdN4VXvFS//hUjY7BEtTzwHUprm9uUvqovZ8VPp8442c2xdEga3lf
hnOUHmdmFGQqhAEQHFDUGyik7uEa4imKtejPLLi9VjOjAU/4OFxLfuOPCjkk7++z
9U0hsNtfhWp/us2+VXmzT58OgaXGngP/uP9Mni09isb1nrIV0wprc6xIi7t7+jWT
e0uwOgiunEesGLAg45kQAwhFbq5U/Pf9iFVxRmiVF9HaCy/UsCotCtmvBvYUdHIW
jUjLHAWS3wKuBTT3TDwLGeBgduuh8ksNNIN/TV0aPJuIYCfEGtApM2xS57hu/zLZ
anP+T25zicHu3Tozut/vdhAMTmpfSN9X+4+a7Rkq1zNfGuagzZYIOei4RjhEpI9h
3wtsnpKnTObvcBwYyuokmvBaIToV/ryDBBw+RuPkhXy+FHGSQkF6o1+IKbORdVty
5FSfkicU+YfooUHgQJiHIRo2Vcw4HW4ccVb4HRFzgO26w8JQSUmqt1lLwAgORlDh
uNLnNfVxdRTYMXsfNg4NVhhHBkHnCp7fgpEZgz1hZ+j695xE9nFFegFRxUBgocBj
heqKMuf4zSxuiIYQsKq0oSoSO/vPOTi2qGFIinSH1sc9VoKwz2cuDCPaWShPDbMn
XI5xMiGXpFRAfdqOMA4LekeHZHIfsaLeZmitctjWynOlw51fQp8LHyVWm73VMsV8
lOI32AqadOsiha1wNZ9L1ol/NnyGCrUhcBGLC/vhKb1vFtSAPGFmxhkV0+Y58Ez0
xpue5lWAjdpeNZH8dvt/GlK6PPENAtZlBXQXkOdFITJe+PVYmsBFC2YpDia2rNaI
mqRrRiTD9SaIhHQaEMJVq6T94NKigt3D4Lmmf773XFlKrqVxeptUwd02sLNidndN
pO//yMxzvNH7Nrfa158EBChbZ/Ijdt5aKN79BVniBpv5MdmPeb6oksiUZY9a+/NO
yz86o2jL/iCMjNxP7K7hAwEnJWf8SZ5NXTzekkI3aMbckMbmCSuIGakr8vGtjTi0
HPtAsvXyoSczA/0xiF4vLxy5y0RRMREpPLxSwlg+isG5UC6uZBwRHNEclAfm26y9
zt/BQBeyqj9N/B/t2/7XWngQHqv7XLggkQpSO4bGPOOqDXSp7Ip1kJNcqOnu94jA
TICFZ4qUowp1KkMQIMU9ppnE7hc+Cgd1CCbd+5UXl10hoLTfuOvJDLbMfhf0Extj
CIYJYoGoikBIrzLc0I6wo8tZ4OGeoayAwFQ27u5//QjR1lPhDN4MqpWvKefxALLo
4rXrLtu5SFTtBSfDTVddN2opeucSU63vVZpUAITeQ/aK2GssqdD02xo3Ek5g5O9q
gHACReS49Wl/mOZMFneD068Yo3XhctXVdFAH11A7h9o3NMP1gL//Md8uW1oOT9kw
NwW9HUBpnrL/D39uMMqBZ4aNR3+USf8gE6RCsGnYglUZs42cS8qgsSi88OHC0077
/9qBsfaKxD8N4nqNxEMOmuAARgk9KWNRG5w/DmUo1b7abUPesS89xGRWWEPTTi80
eBz5ccsFdjUsEVJK5Ysh2E72quzvX6nU0FW3AfSSmivjlyBYO43kUconfNuRjEiF
kg0uvjFY57yvFGqtgjmpu3Ax+2D3iSs7tN3OmC5fdbpRQKrPQ1j8VZiwaU2Y8Q8v
mxOVKWeJ4+heMsvCWLc66ndBiJ0QaGYryt9RofoY/E975//2ybW1oeaQAVsUV0ga
`protect END_PROTECTED
