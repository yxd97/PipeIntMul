`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sVB8yWRoR0BZrdoMQhFN1uK4b1Yr2W+u2NbBB0CjDqYq3BR9JWF2gdleNvykcWDO
MPSLMgw2JOCQM+XWKgesYuvVfhuDypCOiSMlMJ8Gy8cxzLdkB0N9y616SprJNq/j
fwiI2TYOSXSEU/DXvq39Nwxigwv3zvrRdpqPhj+L1DQ1k32u+A6YkHACPr8oxTl4
mAuGmna1zWDEo/3IrJOxVWzq8RvvlRyyMFeCcMn4PR408iD0rN/kYFbRI3rd+2eY
QUG4WOVk9tZ5nuQRgP/kqow75KhaTYJP09q7WoMcSxU=
`protect END_PROTECTED
