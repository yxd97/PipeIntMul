`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ejHWZbKoZUVMtdNnQfTfg5BDF2W4Y8TCzj5gKfQBbdklHUz5r8jElHIK7fsLztlR
S6gEBofqNBXmmei9iy5OZSq8EldHgITmMKs142o7X0rxT2repC4HVb1OJ9lupsU8
+dzezZG4cL3O275TRO+R+iT78JD049aQ93uWby8KRS8kNNiW8Msvz8PkpBH98ViT
rxAbNA+xrJ/PzgiEFwCKB5oWNbsqo4CJiciKOpafVG8HOZhW3S0eqSsMh5gVkoJ2
05WxbZjyqT1lJsZQ0WWZ4kPEWVT6Q4r87CJDsHTNDLQpt5L3R9SWaMdOlr/P9Rjn
AGcMMsdrFs5m3wRLZprBxCW2IYA1O5GLALVm6i0YtMg0FnyVMn1FvlPApEGpFJE6
RKckX1/GuSTJmKlZqXLb4Zt+eFQv2Bxfw2MDIeiVa+xM3LWlsibQV6m87BQukC4O
`protect END_PROTECTED
