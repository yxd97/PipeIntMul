`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/6SgPnOBWYRMFLHygHT7oUHgCU9r/+TFsiwyI72huOKlTuzYq2R5JUwGzStwd/Y
TzAG3tZ1uEvkriz+RKGIAeDouF33KL//gWt21nQSTvCSRJkC1kYKoomcxNI93EaG
pkTzTOo0lyeEV1ZTLh8O9Ih6a6FOQ1ND3ngzicW6ZCjSgg0MRw+QruuImxtKPsHQ
YS9au/T76W4CuOSI5t0ntGpufvgIQkAoBI/QRvxTG8YaSRYSGPEEfhLPpqEHnWJJ
TiIuXH6GPJD2WIYpJ21HBaR5hxNi5kMygnswISZGHk3/NxEg4plhUZjASO2JGXGZ
Ra/cGywjfHnS+Zpzi6yoD03Y3XRbxawgwIdbUl1cWFBM47iBliaMmun4HV/PqKXp
lDCd4Vqjp7qO6RJZMeQ67HG7kFdradn1wYcdTOlBYlTrrlBCH/pMgqaMrXRUFf4q
ydKl3odtaS9zdLMsyPYcNiSK7GXi7KzgDpVieQXnk+m5umw0FGBkSt64Dq3ZpEzF
1qgOD9EHcFF/hXYZzhb2WS9K5qs1eMRZAeRezI1b+qfE2IfTM/dhh3xE0JN+O2yX
tpHbdGWKXX6pRdKyeQFydRNb68eCJyTNf6rmPvUSUahwf9okT/BfUdN5Yr6OJqnu
jUqoA3aoXWeXsdMRm65CYA==
`protect END_PROTECTED
