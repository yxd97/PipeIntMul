`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rE8LffU6M2qJ9EUr/K96IThkxcgVsrK6kEU91G+jLjpOLgRasZYzv0v+64lbbdx
KOefNMGH+F7SBGJrSAFewoP/T2HmY8R8WQo01SsvJel6XyBwOz6UDwT7QSSBIxJu
AVotyVBuGI/kbWyAVO2qQzZKrCpZavgKra/6Bp0bEn8uE4DtuwSbC5OhaptYExaa
hbOdbOPz4QOrrlXi/mmlyDOAW+3Zp7mgOUhQ0O8kTDTZ+1OOUF19sDrYmQF2IqgL
Wg4bjsvLGyoKxGbbSaLNwA==
`protect END_PROTECTED
