`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/e3EgDwYmRjiwMyctGFi5J1kcwXzXC17lcplFBt6R2M+xOeJ80BDGpg9GQCUre2
sS2UtPwFlgh0RI7TaWkh2IuIsSojE3C4sQkDBli7wX5G0o8i0A1V+ytXx/ilRTrf
KlETzEVUT+6+wpv6fUhU5M0FqAKftcdXR+W0AoC3AQVgqmM10FO1gxW+0vfcc6BQ
vmughjIZiAXCpJpxORS6USYTImFaU1g6eHsWumn5k4SzqDbQ2xtfxJUfWzXGZHr1
0GKbd2KvVlRDIUgEUSp6xKEiYPN2aRyjp/cErNYdEpWVN8pEySswv6vLJnggMv1V
LKs45xGgNmXOnCsyWSa8lmmvm9Vn0N2fTTwFzohmmzXQaWr9wTnRWDJTrWdoNBxV
agroxvhDB7JCgCJQyUWUsKOKiQpUF14xHJdQf/gojKc2cdz3i/uT4zCo1K7CS8Wv
Hk99yhZdakx02m0LzwMeKipiwq6lPJdRwLslfPmSv2oRImJIc8X1sVFf9BjmKXwD
2oqpeg0Wkpu0EQjyzkOawSvzPcsRdIUrAbjaIpRoky2DvMcDidM1T+ISbycJlJNW
VP71V8YV+TJbfEYqvOWhSlDOalEj/ehwYF11XYet+5MXmXDDbdga8e7ExLSGb+uO
YojUXbsfTN4p5B178dJGovON7wuLAHYJfKQRnzdVjpIDWBcb4SwIcAlifKpMJ/R7
7yqKJCnvlr09B/9vbYeyG73fv3Us399aL2rs8OwmCtU7VUHR0frKQsEyKkL6x58d
qeeJmwH+cjimzVHwEuHye41lRoGmiA3FTKpZchLY7gMZ6uFsX9Eog71GRjuPts/A
8QFaDAVX0sI6YOohAqhF9ya6G/v/CiMqOGDHatTBeyrhy8dB+gsUfbp+kAljRX+s
EcckjWbD4bZehgspBwB+Me0SumL760gbC2Tp+7oUteDVEo9L5FYIDS2Ck+Ua4dg/
`protect END_PROTECTED
