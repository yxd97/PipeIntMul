`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
otjWUBvmT5EYcNchatMy59mG3SwxtuBCTNiEFqdda95ssz/7c03IbVw1vLVkytTX
CON5nVtUllxgM/fzNA3DpGzoz9HVoTYrV0Tg6UJiyHNayHrJfBVPsTPENHYm5D3R
n9F6O+4fEhbDsKB03VN9bLqXLAHf484YvuN/mEbBPwgCYEti0Dcwf4CYiQXSOSyR
mQ76ovAEgkSgjTSPDWHkIPvBNN5dJKuKrVOXuXrhij+vCtvUCCs/m8Tf6wcX86V2
5iHDXDXVI5scPKY4Kar6VojKlVp0FN+gbHxEOkN4HJ0nPasbgQt3hQpAa/V4Wv9W
S9Rnf2OuLj5x3LWLhVzenDSPG+x/bhBaSTz39t9l7IAS79A6YfpFBgRPWD/LmJRG
K1icrQwTLLI+F5THjA4ut2GruYp0k8pSY7AWQn13aQ5Nj4wVmaU1KpJWqMPsg2xQ
jBxgS64TwtcRM9Ztq2Wapivp5sR2ssgP76amOPIIoCx8OoyZogGvCfBdrBah4FAH
tawZBudi6V9450kNh/eGw8qvmUJr4TvXFoPUOiJ+MwmCzHYR+uY0GXLv7bcqyqT4
39afOTuLOHJshCSHCZdbrbItRCl2yg7wNm4siUsOBKyA4823p77M3HDAWfJen811
ksktc/4G8OMeuwCOOWlbjfozonhYm1HLWcqZVnVtlj3J+9g6w0hO1Mo8gYT3YNF4
KXFNbcBJu0WOBZD31hU9QKQVnFBMk2Ih25ltCk46b4xfnyOjsY8Pa1Him3xCJNem
XrwH8VAHxYQ8NDPNYb89PcNm5pW776mK4s9FZFIoB/iLIjgrximuzk87kI3n6DiZ
n7GZNJP1MK+IAiNlbv3JW2/VdsSG1AfsfES4mdeLbvl5xWK/2st+Xyz4F4OgMruu
e9eHNvLhi6kTjZS9Pl97OBT18RKAuTd7z9UFCQvI/DWTfzwTWGrF+jh5MNULM8ah
TTF187tckBEp/Tb2wUXBOFMd6xwHszCYmkuthMlJBzMdVs0087ZzTa7RlnAg/6O2
uOXZvZw4RULZVqh9XfHbVoW9/UtIyKUlYyUUB8uXTG5dLwTXrM+xBX9eRavpFMk3
DzXbj3EDF2YEKnjo8at76IVBB/aryb5TWWSYRKx9dvlhRIvI5ZeWsfFEVAhsHAm1
T3yhTA9yf6toAJqroyDOeurfx8j0S9OH4z+vYfO3LO1NeDmh4ATDKzPZTHuP8MKR
lOAaAhDSoHzmDkbMjwRBrkAvJvmSvRiasqYksW+ipoLeIvPAQZA8YKo7mLVij2wn
2XitjmcDoBHz9ls6jyjBmla3EfRDhzQHdkBjeAJTw+EqHYjUu/UnlzVdt6xd/wC/
EyKsqQtjvnV13ysVpx2PntHFo3oOYavwzat3l/+CE4XfXBR7zvugERj59HYu86Hp
lvghvp+fjWVwGzIyEIxczSf6F7f/GrBkuSZZ9KGfY24J64ah/qmCJ6RdCC7QeY0u
e/LWsY2n/ZGwz7CssIKZT3prjt7RyJhWBeBDXSQzp4qaOJQOTehZwjDwUymCkbtS
+DNRurYFagiqBJ62F3SWzXGhUsJGlgHITK0KpaguHfnDLcz/Sc/NQPyDNIZ6RlOs
Yxq5rj+RhTtylzSOvaZoIaste5XoqqXaGQqmxaO7R2egcQv+7Ma6zsSgDhjci5d0
NB1Q1N/RhcTu4K9ePk8LZ5G4Vy/ji1nKnwQEVGM0Otx1HByDr/LhalgPJC9UGTMs
+7OUWntkCWP2eDlkI14o4l6pWzvDq19s4MMnOzxnNv5wSzUvjfpFp+qduEpGq5Mi
UWIm+XUhPQAeG/lG+hNkECJO3Vs4QzT+prFq0BX5PIoiCIFxHMSSQxa+xUS55/bo
CulaT/hu3RghGftQGMwRLcqZUq7C2j0LaLP/HmMGk6YFY3qBY+XWpsTJWziyms5Y
0uVpT/2reV+cDzw8dhpAtYehj8QhNuvdm9a1kiqM9J2hIzCjEIMA/tj4AP2WHrXk
/N2G05NkVTHwc5BleL0zSg2jucsQdeLxfK2U1tVFIsrWwhyWu+XqyZN3yXhckMTh
9WSr2VIQo8K8vu0TQ8EaNt1WKPWXZJyGWrjyEje+pWeSOzQaJnZDkHlhDF7smJ/W
DZA0XznJwe5DErNHoL2QbpFajqbrbZY37jzfLmrKIEYPb6mZ4yRu6tQ6mSZPk3Yd
9aZ3k5S1AzpMx0LvF3HA63tc2Bayw9z/sTaqSlyWjcGCpTeg0Ef/GQXhJioverJW
B4huEYw8l5BfPzXMUDQWysR2AxWwqFXQX4l/x95WUwFQrn6XYSOxmD35TWAgG1DQ
dmmA5G69cx48yUzj/9qSVfOOS9LOM4TE2btCRbL7uieRJkuXvkc+TFmZQKXStgkO
DW8XTGhR4kxQPhLsliTlD5RqPpNHDZEpVpf1RD52qLqbWGvV4Kj55fBKS01b2AW+
eSvQBQDNZCoKuITPgc8+EGYb8S09g/FwaJ50Ex08B5h2CHiMgIYRCpdg7cCqWbIs
QvzjJ/qAv18Z72yuiUMw8iuJYFfQclt0mcQU0loBLzAL+uoT0VrLcFsMuhV1q7ID
mTI0gM0OiQKJnvyfOm3w74Tm05GFfqqfHmBmf2k5fU+QNAs/aLQhlH6i2DPYaWfi
ETtr7yO8j/Dpr6grVBabrkket1aPOa5RCbNwzRe+m7AhjFodLETYODrSAJr2+cVL
kEuwB5SIZ3TKh5B9QbzEXLNty0zNQQntc9zBuUvntULgPcouCLzkLHfyQWQazlTp
JzPXXYhQ7lSRbxJkQeUX82BTp4DhP3LM201zIjNeCGZTtDP9A+2s47HaEK4Z/+rK
`protect END_PROTECTED
