`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/lmDLTASp/XP4u1Uf/aqNLPtm+ePwjIRFZ37vyiyT2aC5SW36f//XPHbxeGuilR/
Zn/7HMdnnUo/qsrDRRW0zAGj8LUHoy1k9vR9Y7QVPr0syVIYbfYOlCAqpAXbu3uv
U4KRyo1ZK91wvGrUc7rJ1bp8Jf0O6MnyGNh3aqX1dpwsA7PyOGboV5dYHexHqNy1
A++4gU43JeDAiocmqyJydFY5vXxUW9TLQwgtKboH9ceJ28i4NSwIK4mfrQcZNyLR
TIfa9DChHvmkPdM0E0DPkdnaa0xU9eVj4cBuq1xO3jW+hi5zl4ykjkD+VDC61Kx1
MZks5Kq24Fzj/NIC4R2wAcipz7AmLSJTarYoaa3Fi4kHiSxviDhxSsBHog1I8C3T
WnbryiJuHlc9AQC9Pi4g9mrlhniNgYAyaT0M1s7cZzDHh2SF4DnLpca4tDY/jue7
tlnF79TpaGuVPnAI/CbJHMFUbhEdRb3LvYciAsbQnyAeglByes2VzYmGPQHAJfOA
ddprJ8uqxbdxrrzNPb+Za94CixEKSd9QorIQaw2V/7TpcgQ1CuYvPBahyh4/nRZS
`protect END_PROTECTED
