`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XyAkJGORDPt9VyETYv6qek5YqrKfbbEY5TuqWGCLoqVamUoH5hjMuXUa85gcVpuQ
6MxCRsTfpdJ40HJaB/CYNIkKnCE2A5OKi9aJEcZEWX8Q3HcOR2fIHZK/pLoPz1wB
cz+7ECLLQBcsk5KwT+rfdX0llRK+mb3liTmfjvTtRAZ8n8QzWPXn1iTvZFu8aj9M
pP2PyOHC7cvLICwNGywuGx9R5RaYzPjO8bkOAnARahPUW8Yc9AkwvLAUfGSJiSYE
p/I4RLoQT700alSH2w1j6EReIF/ysF97Ql5QpTjWhUFUwqAN5UGDjPfeI0IQlQg1
X4g/jhU2g+pOhDo/mGV7LPbf+YkzUahecf5y4ryZiARjbWOR4YbgvTVAak7s2gIL
E1DYCXtCZoupsWWCywUCcAS+pipLs0FFZthiYhxzvA3BwWLzd+Sxgk1NjPMEdxOo
NbAKid77F+JRQL/1G5H1breHLkgiApceuTVZdXxWogYwDtVpEIJ5Fkr6Ul3PLkPE
KdOXfI3wKflGOkBct0/0cWlyAqLRoGnSxQU4t4MqFaVIeQy/U+47I+/xwdBZZXYw
JQk4o1ZHroULqpRhgUBpLdbmZzkBXr4KRysvZ3u4Y/o5M+VYOzdMj4UO4Jeegrnd
pNRqHI51kWqutBuSBUFh3A==
`protect END_PROTECTED
