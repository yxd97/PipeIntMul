`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzDWfl+TnEukhyR3Y4E1V+wBnymRSKHblLWzSo3Jp/l9wIrGFGQRQRFGgJAym0QX
YlEx1hGTUm1Pqo4yVZMhY5Kev/iF4pZgujmSRxrCL5z9Hw5wz3hpD532CNWMnUL2
9KREYPpF2mb8typakI2dlTLIqNBVaIN1VHqJSHf/XzgACNsginWZ5QV0OdyMI/mS
SEi8Mn0579O9xyUWhRpqmaPBjwkRq72x6dzxNBAXhHe57eMMfX181yeSUtWOFmWk
VulHwuf2puN9FC/VWSHKFjx+4+r/FaIBvdNqvRyGyUT8wDYTDyvnnQwniY8f13Jd
f6rRVVThZzSTAcvko2XsqqF6NtwGAjBz+Fz/cKQGFLW4O9LjiOtHmBy+k4RsEwD1
73BavTPbBZe2sMPAkptFF0NcjDECypXWHPvEuBRqOPvBVM3DfW2hFw9FE/NbwB63
lZJKKLV5GOmkAuYmhkzIPV9rUk2SoEg1Ru811QUzqjApH9oeDwFuZNUHFKDJA2hf
3V1hIilyDc23AJWKFBZPrNpd/z4R09ObPJ8p9uEccKBv2zFd6+nGdsjTaRwgtD3v
VQuakv0KmqFzPBxoVOtvSId6Q+1g6m1ZqCsZxQeSt0H5tYouJSz06pcSe6UD+CfA
Iz+Ibh8SxtYEWMDQxYbwb/9rN+lviqeCi5u2iGovw68r5ezoIJ4/uQiK1TyZIRyN
EhtulukrgOW93ul7p+kEPDPUUm+8zw8nOHIqFwXUKa5lmUU67KSttvndXOeeLnvF
OeAVzIQ+11jYGtQL20eP59KznAHjLn1FeqWpcvmXXCkNnqlcbblMbI6wumiNbGRu
lV217YZTVci51D7AXEDzKewo5v0BbtvsGDHfa14jlGqgebDe8Ta46+xe/AMx2Qtz
kRSQpoAxNX9/Cp0w/AoC8/X+XWGZW0oLFON6+ZNbdQW1oyL2Ur6nhdobQfg1EItS
8U5lhF51sSZuiB2jmc+4IncnGSRNMQvGBxrc2Ri3djYquJWanany/SHl1xhMFjal
+Qkzfl6wwYRlfBvrgZVrJBR6dGNuYSc4iGiRVw9xkqPDZ+aYW8+T7fpTJsEySm7f
/DeOBgPpt2srunRvr8HMLAgPkaqBHwAtTPL5Ppt77o/nqtWgrzUuXpXijOaXlO/9
EO5BGTjhy/Fyt0Jo5MGrkQF5zTuXE5JfPliBKzVvKIncds5b738f4uhAuu6J+0Ca
jATSq/zhX8JDfyVx3CHgGfDZYHnNzy5TOk8WpQUCuKe7Mj3Mmha7f6oxVew06b5P
Pim7m6ubmuBf9O+9pP7Fhdv4L3S1gZH2RE4myniTugzJw8jqNEi9eYu/kZ67PKy/
LZJB7k6+WWWIel3BWRW1RKk02gbL9pO0iyeuVsoFGuz4z/NqDE95/t3kwJBaps8e
7PqpponSC9MCy/fekiVk/iz1a2LtkpI+PV0DOdIk6ujpKkFayHiYiQkgDzdX5esa
bWNw+CCWR6RfExmfE1BIBj7n+GvIr0hVIS1Xw8ouzAw0XpfFnJANSU72tmYVPOG8
5uWgvAbT6fGbtChes4QcSajjvhJ8TkYVfUxIh4V8CWL9ENaMKKX9qJTbljDWRyeJ
4rM83vW23wD/7T8NWasrcoP/nktQ6gCUGeHGuPoNU9JHiRaA1X7mXk6Ve84XVtOy
mt/ccHhqZU3QPwlbV7h2zij1cVyCMb3f/G+tdnXb8p3C7gYO+RPeSq2kcvHGDNcq
82ru3pDEgEXLck0/JhITMDUnouS+Rc4fsZbGj9gOs+etgjFRroaoJAsYOT5TBhIz
`protect END_PROTECTED
