`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O/jSgYJsL/DOemBtAwd4EhThIDIETfaVC86bm6woGySYvybYeaqKL4Sa9CDki9Il
46WF7+SMA4aEncYI6z+LecA6DxMfd6U1e2N5aEA4WCtEKR6wUPkJ2jK/WsTxs/Qv
w3+q2nB/OXJzHt+xVlorwZtgRmYGng2NPRPAePcyLgzWVCZFRJ6BrEe1u6FI/CoX
1iep9ubHvn6mqKvopoP87y4zNVR0wTwZiRMcFVQiHtwNUKbyh1W551yX+BLuOusG
SVl8HIsKrAeNXf7oxbPqLEe/avZeq0nrwY2gxeqQq3U=
`protect END_PROTECTED
