`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gbrb8SCgvCJZ1zI0hQCoWqpUOv5UvxZ6eIWBN34tWA3IOwIQA6ZQFQI5sTOGxW1y
0/Szi+EYRE4IqMI7jnQFbZuI3YhAqncPBrIfOLyVe9MRN1ACw/+gkN6j3aiuNKUG
pam7YwL6+T0tI8oBZjjnUbctTh5tInbM3bQgIPxnzAaCuEd2svG8FoAepu2wxPea
eYg/zryeb+iAlXHwgTnI58sFu6s8IV8rOBxP2wZEBJLeoz/MUWGpwtKWuWjtK5GO
taz59HePJ0YITa3H88TEjFulA6A56HirrPkC2+BZocsKOWeeM4/Xjg88klfItPMh
W/zGgjsfJKs7TmFMORCfXwSPq2qNa2MWYeyOP4t5VmkATuh/jfGgLQxb86aeLbeq
WWGRLqtjNYk6MJtIda9da3XJPYUAF8E5Vq1m0eEeRhTm40b9llar4uMaxJejbUvU
PSYJE12UMStUladQIi73OC9A+PK2BXYZWIxp3QsTaRnQXC1rmfNqwhoj2dGVXykY
+B335NX88WJL7E1o+DqpitnZW+YE4Bw23OU9Aq/MN2MQ+aoci20K8A53cCVEI4i3
PGgsPqF/wBV5wjLKMsM0MxOTtjVIVqZucny6sfqoNihbyB3aMOEoJvtoavBUEXm8
/zTU5JKt5ZG2Vhmy0ynrY2oz5q7tztPrgsl94MuXTPRYtEWotuvbykVYuwOHWRlt
a36jmJW3/JW5DUgc2QsP+r6OqxQp3tEtTTP6VIdC/d4UiKc+IGXQiA07LjAJ2eb5
KoFrDMTkHG7MwscmYhyRoD+HW8eVYaZNTUCuIRUKgUQ+dvjCj0WdD+P0KLHUmJ+5
Sk/KNw/+4gTmPSUjByZQVIaA1U4yTQhUcMMnkpaC9Aq3GYSC8UHOvp9r7c7mc8tK
TJ4Am27M9H2HkSWqBRcPstGGQMHvW8Ing1EZGXXcyQ3grnJQtIm1/4lqJm98Z7TH
V/2GvaYPY92KSNeoghvTm1VyfyyTsFui4ibuOhvJX1y+vrH9LkET4b9+qIY3x+/l
cxwqwcopAWA6lDoHaXcu4MPwoNR8jXdj1vqrih6yd9Kt6fg/Yr3EXJ3KLcnhJoLa
HGJOw0B65FndW8mxLGeplHlbfhPtdE06lfdXoBh0jO//5N7s07RuhxotzfEnBtVg
0RbbkdXjnWcwnB0EqlO+morRiCDoGiSUAaNqD2wPgKXNausm407fCep3CV6o0HAe
MzzBLShRCc+QeuV/F/UPUcUnfEfqVlJys6ec07/4+u8RaUwQJcZKv/TBWMUVi8cN
tonS77oZT1TC9i/NY2CrMM7ggQyjq4dZGDIuvDTSCOggtTg24m+NpE9oAV2LY0Qp
lvA+FlaU51NuvnsdZGqVPNJPEFBmuC9J5fsISa+PIMxWfSROa9NRD0axIBbtybCg
2CjcL85ppkQ6qW6AAXXA9efD34T/pC8fdhpfX8XdIZKLU6Cv5pq27zkvfwcgncQh
e1tOulSj7Hm8zB3GfaeUUV5SjFlsY0LeF9nIhYULDfJecCTgghajdmRjS2RK5g0R
ku7yw3Ja1sgjHf6gCwiqbh95yGsJlsD+e+MYgoAfb4alSuB7nLj8cqQcuO4hSTk7
4DTcBJ2L04PAyAlr0lybWYnOcuTJeIqOpgjwU2yllOsC/t8kDvCQv46994TslO82
7pfutnySpP8IwdTiXGNh9L+AY7Ssy5yJ5UbKs/bUrd5Zm1Q0L7NEe/YmAJLkokQB
oRDU3tsH+5dK09ZzgVzxoumrugvTnYt5dLKwoE2F7WxX6e/QCyx1mSfW5R6QZ6pl
PR2siuePFlSPxQLGi8nqxQYOPfvIKihvOVuBdP6fX3EkYpejV07IEx17dnjsr7HS
/6X+wAMMG2hfG7m38F+0Mp/DKvU+/qzKZtGp3xDLvAFvp5C1u9vyrZ1KmlfwsHzR
Llcr43K7FESDeREExq/XzCI7s9swyHOLKhFXsyesXNZzDp3nJI5BJ6rYcsALqKjk
rVhCaFUtT2kSiBczTFJr5ckxJOpenfdgiFDD0AUo8tgsG6ra8r+i2gjv5nXLnqrm
mObl1d5YNAbpZOZ7xLRc92D5ePNJj31iQnL1Cn283qCx2YGsNWb/L3C7ptIQ7O9A
DUkL+m5I0Y6wmH595yXdwIh40lBXnPTHcFt22xJ3TUGW2wu1ThlOyYlFrozj6O9D
aPu4Jzcx25I0Yj/sTVZq3sY6EN8bMUyWAe+QdZ0mSnmDM5Ysx8/4garbV9HWM37X
vR+7LfmgmT/qlEXngbuT2o5PfOiOhWAAqBPKE+c9As31QkYXqjzNgIvmWXk6SaZr
KToJdJyHNyS3cnNiEyrtjfXH9qXY6PCNYnSalYVtpvMWDi30b1SWS4GCHn2JJNAu
SBbcifU60uhwPXuWJif4VhbCU29Srbqcys/k+ZFhQcqdZJImsKNHpV2Im/3MR+ii
gKMctwttzLLmywpf3Mte6uUWKUVEwIFo2bs4TIcZoJYwu8twxZS3sstfhTHsfn/d
0FRtpCEcMnkwCt/5izLj962w++lvOVEP5seVnIgWe3yKkBuc3Lhp8wk3K0gO9Yey
Xe1DrMXF83uZSO+51X52wQbdOmzZH+YT8JU6fgzUPTuAwae/jT5WK6CafesSLDIF
+x1jUmh+yycCRtdU5Ox219vVVf4zFst7yOwhsqimoYJcQbB4IIHhR8OM/F44J+JY
zrVmvPbxbSdpgO2TOpAbd3QND/Snjl3nbsoumCOkHET+RxXAq3qjVfg3/sKt/m3l
W9dF2ahbIb3wz9EjWgQD+XqpVNLsQ2IKcQQVF2wxtioU2fKy3juOHolMnXrL04Q0
/1qHpdMC0LLUmkcacJRrbG25Lxn6AGDzLrG1sV99E38Kq47exBW/0qA7ogzbZcim
hvoqUMrmEfhDLtPILRWBL288fWmgmcoNER9kLmM8v3dFfjx5K5UKf41PpiVsnfCi
R9R9eJsvs3VO8MYi6i6uX5/wc0OREpw7sRO1Q1CBjPQxV7kDD7yedR/CWGIWN5X9
oHj9bqIUW/hN3DREia5uXRgxfJzv38Qc2InFHOiXt5cZdFSOuHTRm4rCV3NpTb8W
PWbSjvVvQK6uk49QXknerFJiWpZlAOI1CYtS/W8EG0pvAvoBnevQhuBeozZO70TZ
2Zbs9eleVLW8TvuY4QzDoY6fD8Tv7zs4iTL9K1qsI9u346sq+jQt5BRdzcz9d/Hd
qWsWQjAgeeQUDu/DWJaY/ZJWQT69bqnJ+ncW+zTGbCv5D30+JEHOYUp0hdXuJw3l
8P4TJBtHTau2UZfzA1Cy83KJnp4o9zMrxe6F8Hx/fJagDL5M3KUXnNDrQjpJMpDa
pLZxtHyUaIIj09KPNiypzQjwAXZgPiZZivqH+FGYo+Kzp1qzNpVCdciKE0o0+hsV
gtJBBgkoFO+JiHqJM0Xgku1YgZk2+kZujPyyaruEn3DoX/06AZEe5u45kkDyb2RJ
X5lyf6l7JSMEmRpq0GcL97r/jM39d97relv4cvBwgXRl5QSpjtsE55JRKc4k706e
LzmGc/zi60tIVewy9a4DKQqj79XKrmZ76/8ZnQmMIykRAvc0tI3ApYpkqjbyT/w2
bFSj0K0xwwf2RyBw7A6ap3nTEZL+Kpmmc2yyxd9v5eRs0Gm8OQq/DmhWR/cQEFLp
TlK87HSCi6b6v2FCz+SBkaw2Isr9OkD36r8a5phO1WLN1MliD+ot8DxnGtmt8YqD
rrLfL7ZcTzIXPa42p4JZkXrhn23U7HSADXOFmPZrOgWV2/49m02afLLzWqaa2nnC
qmyWKE7KUh5p9PYY8DQjG8GNcY7Bu3eQn+9glSv76i7PouC3pbJf0qEwcX6UtiMQ
/TpV8eAacnMmxqAJvFV5V208EPEMMFxBm15irH0it3VZONDmrgglPZAy3fxpmbhD
ZnXD71HOGiuZHuou0cL0IZ5UQK/1JI84MSZGRGCij9cw9XG/EM2ABnOmBeOe8sua
uSWlZmOel7Hvh0kGHfIEm33wl5EMm62il+A3aMncdRfsLrfXaqnN096wFG3x4C5C
4jH4xrBw6luWKpMSy8FSeNDEWwHsboov1Ge8KT/LB1p6IQfz0uyYCq7SRsfnScZF
DixUPrLqxR5M6r0yDHwEdGoUk390f0ZLjsOfyW01VnzNCF8oWAnaOhBalN7/G1NX
RXjz+DcjqBXYJ2xyWpFmrrDzi5yRGc7NPsqnOqTq9J9ABbOdgDoUoqoUbMQG9zGj
RFv0Kqf25C8W7Yb9TIf+3bFV8fFct4WeWIgMXyEluimL0XGMzCUTxKiZta3sJB23
C/ikc7mc/Trbmk0JX788SNiMsHEfJnMTnMBodXmNLHM/sTXkfL41P39zPNp7bAHj
Y3stQRiYYm1z7HLBkhY5s9QfWgB/xlKFf7MPzk/wlimOXOA5hXPxQd5+t3UnTH4+
WJyTE/IGGB/KgTx+engbV3PW2gs44YCfl1WJv+Hk9jc51Ppq6nw5LXSr8gpRHR8U
nMa7ostch6wToxHj3sjQ9Gk22k9R+Zn6gBMuEk3xfsm4PBoobyOFWvwPu7m9IFqM
IrXdabPkFwPJxoxjINHg7A==
`protect END_PROTECTED
