`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
goFFsqjTtg3PYhqi8VeDhvEwOQpYG3AQM0GGW8bWiO0vuOJf1kYZnd/JdlprZK82
YxaJjc/HGcrQ4p5yDDy7wpkvXNjJgj28O7hZJui9LoJcxFO4ElTYAmYlFf4hw0gC
g65X2WbWdMTov+Nt5whD9ju9imbQJGOaSneUoBsiBRzU3rQQoraS3bamhzAChQGw
nnWA2+9QZQJjUmBg+gZkxeu0cb2vEql6m0MuZH/u3WbniwkOlb846OEN9k1WwX6k
1gB6+EAQYK45ohTAatIscZjX/D6mPMpIYu6aPBr7suPERFMQaA5j/ulniJ4M+o9y
e+CPLgu6aITUqdhwHt7hkYAcNLvLFXiDWUGQ2Dzt13oNoMxkcpZrcjwQd/JGCDHD
eaVfxtLNp8E/sqpPY4uwWLTZ4tei2w5LLthXmUXF7HuW02+/jeQhOlYjdIksRO5p
`protect END_PROTECTED
