`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCMRrwnAIOXEUZ/cW3MPkK2SStW3XI3JYqCdZRIwkNWpYc8Ggm8GbYCFY9Kd87/W
eVs1K2zXvTMbQ78MA+q6bJkeerbRf380Z2x8FbE7r5fThJhp7Ce3Cu/VuG+lrs5G
/dxEZLn9e2wE3MJT2wO8qvLQS7eVevP4KddmDbMSC4itXN0Xvs749DpnuLDG+lDC
znQPy65a0wZfJ7o9LovRaUzR1OFZIlPxsxO492SRNkozQEvED+AQQw+J7GgN/85+
ajaDlFFwSBuPsxK8/k8sRGDaGLgV+IrUZm0wyywlDAo=
`protect END_PROTECTED
