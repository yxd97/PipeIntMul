`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RwzxoBbj4wCJh9fx6w7cb2nrWEEz0pyK7Ux5GQGEUaJwvXh3rI0DcDNYMzw2jx9g
5LJ4+YViUr8G5V5ece8JHlECLFH+VRcTNNFoL+RgtKIxV0n2lsJlfSOy4jeuHJtG
WpBaEk8eIQR3NB/+1e+DRKqMd4+RRyY1uW9OdqHwSfBl95wHoVUsMhZRS9GzM2Cm
vViuG0mmDCFNkCMdBVSMeKDc1xUIQclQADlxY7UgP18zfE4Rd6AduyXFbu+pSYea
QeVeImqm9ZpIyBJP2FGrg9a/zCuVF8YcmuwqvJ8vT6I+H8nhnyULoZBAVEjWT3cZ
takA8ScuTBQYU64cj/WlGkz+/Kf93gVE8yQbUKJ1oJz2jC/V9x59I4z3rfFwEcLV
LtTROXi68RK5/pFZkDt9EqI9RMr3pzu3REHJuhXBnSkTdW8hn8VSvZJtPB4PN0iE
/XqTY6t4HjvVjPFNqXbveYP9xffpSSteoCFXloClUY9KUJ3QhalI5NzFYlIyZTLE
0r1Aup7vs6vV1vlXOPEAKeZCqpTn1VcOzZP8yDRF5iZNlFPJWcFnZm0V3uk/iaYA
aEwl2SfRmB6Mg06S/+gMx7N/s5cMigHRD4RAO0wTsp0ZqdMxl7gSVNYG4HI+/N7w
GzdXL2Gks3chkRoMQAzm6LAyJG6QefjbcyoA0f0aqDpdMneDt11y+YSCDxIBtF9r
pIm3DYHOqu+u2OnYGK0MiiugQj9oYFRttiOC6QBo5nsDIlkyDVhsvbh/luB5FJV+
tO5wVKEY9Q3aezgjWHaR2i8IaY81w8mIV1ARcCG/zHI=
`protect END_PROTECTED
