`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvvXpYMbgBKx6HxOEE4mIoIef5Tm6fPTNdhU1z3gMfq28kkd0/LLKNCjdUj1nxyD
LT+Pzsx1MpNFtyPNpObmXDDhxQ5Qrih5v9ZlGnwaUhjEog9wXuqRCtQjaft3E/oo
AcnRzFd29RYcBcyue4U3ZS6CIrS5phbT/xYFyQk7mrB+gbPxqOjwD4uFikMLlSp2
ZynkxdMGygGPLGsetWwCRwk5aNOAoWKuB+w1gpSN1KrZ0D1k723E67D2M5sCXm0b
u4WOwA3ScyiuIf3/DiUXl6cS3U5i+EN8JEmCO974TKYqPeTGBwnz1ku3Uv6+4KCl
I1I65DDeRIZOJf+cgoj9BbQ7Q+TteOX79vDnX6RTJdwZyqEERE2Gjv4aR+JBa2/3
/mFtOelJSZTiqn6l6L5HvofzDPjDItlylHCfTviACgYJxws0h0b6bUcz5nzd5PH/
VCyKx9dG5Yuu9noj2QBaMIs+7Csl9KbguNF13gx2SXPxyDBtxo5YWbKK8mDYK7+h
hO053wvKXentMz4+bNF06h8pGwLvGvwByq3xxPMMFCje/LxJDVksIbkdopJco9qI
T7eelkCx+c2JR+/zfr7yMrC0Ba40ii+KBD/FKjyy5rr1xoczw7FXEA1vhQuET6+f
QtZVEthW+ZLQVUgWWLkijg==
`protect END_PROTECTED
