`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4mzRfOqMPwMsM0hhroTjLKe9+P4rcAPXvAdjgqME5PL0Bmu0rhiTHN04KlTSu6Cx
9c1jyJFxwnH2Qrd+06HvN1D9KYWzaxhlrfhGom+4wRIRuo765bp9YLZyfkc57uKd
oF9BESq8T/WVQ0cTncvMLl7e4hjkcLIwskTl7XcXT24DPaz0v8/z1BCr4jVXTsee
b/pkaU/bXE0wkZBIqdHA25/TxEkCy+XN/qAZWYv2RtP+vq4HRZUnTpYeBSfXO8xy
0M1iCDrsoJz+0IVUVYqvxinvoBAqCZqR9uihrlGp98lCpF0fuk9Q4vJThhGupJBg
KXeLriqoWijZRtKCwYM3+UzKhUgeKkr7PeO9umDxjSHHGGgzm7lVWbGj4k06CU/Z
vzpOrXqwUhlXLv5wcu0yiDJYqTZ0NX29sQI4iTGAGnYxe82FHUs3ObJdiWuklSsu
DQjr/FNoM/ApbR0rZta1eFJIE80r2PLBHSLxA/+nBBcHp8fgJisNxr4HNzRq8ZWL
EFUrPuc44Z57q2766N6qOHocfPIqlgaym5MNP+vxg1irhlOCmKp1a8T/YWoB14f7
`protect END_PROTECTED
