`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jZzsOH0AmMXcyuCaWxr3aB9lWzRGKto2mWkZ9oWu43mwLmnKBRd2id4waJJMu9D
A/1XKWQkCNvgW5rN+1a0s8IJFjg+DOUWz75e2PnAr5J8h/9I6rzK0F7IDZ7UrP51
Tqn7CHuTnZjxYRbosBCtewL59lmyVrf+s+bm4/D/EDZQx/RFnOOP0ZUnglW7zKhb
u/+uMCNtiB0b7PJSV9czkN9Ep9azj26K2oZo+fm+Y5sxFT2IyWl7TiMorzjiJMJn
BoTBzgoOgTc7KOkqZHLVfLqaL+XlZQOJbz90DjbnJiRx7Nqt9GX8I7LuslSxLoUA
LARoCBYSIjZ9AqVYG9lcEvK9L05U3CTMo1iCyqveRhG8Bn+ez6rG1ObGc3xvb40Q
5I0Nlj5PYuFZvGsUqGYx1gLuW4MeVM4jYA+QIA+Kd48vXGbRnTBs6tiUe4lwsxID
cQzX/4cLQQoEDeCgv2HqmT54pGtAgXEOVXeDrLHTyMSwInFLlTLjjQn/JbzTU0pq
LqPnWRxnbN3pB7iZXMBZGmq4lst0XkLwDrpuKLKYONO8Evu0fomtI1V3SwIzWdsY
`protect END_PROTECTED
