`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4xeo0/a0Zt6dl6c2H2cABes0uQUJ8bizEfWTkDsePxfKDPkiQ69aEy1fx88AeIWp
axYO3CVKpMeDDr25469Ih2Snl6j4JFj1Ytf0zpPW9o5fzypE44/9X7U+6AnZ5ZRB
2qv1fv4XGHVBU8alu58qvQCyMiPDJTbXeBA7qdLXVTfS25jORjZYjOo1577ndKrJ
qpr+joFtrvyx6s38P54D4plT8ERhc2nO33vFSEY7kElF4bnS6e4LJ8RWvnoTGt5T
NZIqxAkoxAlG+qWik1YpqcsfpY4FxApzKFokeiy+mD6iFqQcTFFTqb9HGHsXAfvH
yL0Gpi0dxc9ZOY/YKJ03kHULIoOs3T4X6JKNlpciHyN1WOxv6pdEoaEmPu2aNXpK
7WJoOdycJMPyILRHcL1FfCnXr+OxIbdGFBewNZysdfCjRpex733NAt5ZX26l91um
ZuKnrwu6Ae6Qky0YIRfX5cA0ul7wLrB7XFm899htWb4Ze72Cn3/IMjXgIOZBAYrL
iOm0+FY1QuZtHfuL8VTcI3QW9KbMMEDRXljOMUGRVXHSu+CrYXqBwIys6GZRweDB
PFBNznIt81aTjvx8LRrl+ON1X9rMHCAY1hO9ixrhQhg5SjlTfws86cRzgYXPm+Qz
J4n8ro4eEJFjm6sbKgfounpHxfF2UVFNS+UjD7YAE5qKWq6xBseCWWgpwAhv9Rv6
RbkBB5kbJAXEZDlutyOi+oLQSvvIP5jE7kc7z2L1whlBEfb1tDrr2hcUI+G5HywB
bug185sqfeVI9ncN1nZghQ==
`protect END_PROTECTED
