`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1RmOyhYsYjRRtmBpxHQM7PL6Ex5hBZDt33R8P5ta1j5EasCKmf5azAuoNHS5SbY
0cM8/y3Tbv0NjzMZE79wS9xseY/xDv05UzWgbCFBGbza6oQykNoFDzicjU/Jbc7o
KbabTm81ZUmVAlk44gh84/clXdD6cUESHaNH5FOdWuhs4iCZRYZ+pJ9AFQMkVdkn
JWE202/79JcgiDg6mfphrYqZQpfxi1vGsVlRG5TiIohIBl9jYRin5tXtJ8ISkkU1
LJFiKGSgSsSDshvDJykwfdEq4cothl+Rg5qw76ail0bR8kL+eFWGxCScoelXL7Lr
g03e9Z4vZtY5yoNJSiWmjScixK9OgvwTTKZVz1qegLZpe+LO+sSFYtnmw2PTtwFS
03iyuWPtzCsMIW7oCUjSQ1IGCX6g7cxR/kbJhSNegjkdAjWIjf+1wdyJNohahg0K
g+BmUYLmurB2ckVQ5f531lgNKjyDXYUpv46SQWf1tpMCrHboHohyN1GxLerL9Km/
nUgvMF8baw5G4lBKZ2tvUKW8bksyJVqc+h6FxrmdE0yEgsXmdkc9lXaJ2fwI9aCE
MJlbzkb9YvdJaQO4/sMvtnNU2gDigMR5Ww7kyM86eVliMoAkuXvG9AgzqYk8KdPZ
j9C4jUohcU9D8yCHEyiMsMR7/Nt+P3RAyVHT588xSc3fGHZldr2OIwjXDdth6nys
svwDTQYo7alYhTNa1QB228XtILyLKYigV8OlrqXl7Ny039KflnzoxEEh4Bo8cTyw
rCPjMwE8mOallGIjYRuKCvFCo2ZjFvOL5MTeUxl9zoLftTI6N+JstwavLID8pXHz
GLjtsBYiD6S+pD5bwBz+/gbRM/NZRFpkOJe7rnQDixxdIUKffrYGxv4Kt3GFP3hG
qwtFBqmiAJkQ29KQtq3lrdxoC9/Xt6XgsDK4a9IaxR/hTHCz4TvvamCaX0swxsnx
QbPoXkhOpPdxA55Q2acD6xrlpmnH8gNmiaAOXCcyrVy3P4YfpeonyYseJ3fzwGfx
twKog+e21oH5+scg8hYwvq1tXmj2b4Fe81blO0NB4mT2OWP0BP8xyV02G6+c5DNr
RvXQNaw5W3q7gdWcCV/HxJ8T8QfhlqzW3n5m9vAVlBspUM45sOIXuixl/6/H4vSv
qw+OjKTBilQbuUyOf3FTc+AOAyM/J2B3Zhy8EKhWlGrGDckqQU238BiY38pQoYMG
Arn1sddCrhZ4o8rFhGvh2vYOBUgo43dAKvPYo9Gw2MNAfeAwzU2Os9R5jNn0hjH7
Hp8LiEozLZVQe/TwqDpMVF+CHdAnKrWLxLkga/ZXBKsbPz3Ur0srN7qQCbnGPHSr
SuIFrY4/YRaLEHPewtXMZ2Fj1fsrY76gh050TQfMYUWc3U8vQk5cf0xCaMIuQ95p
0A5MGS+vfMhGFULZJQPoEc5cFJ+5Nua2C8dT/3VCxQUkaL0q8Z1fj7kEiI0HXq82
jBQAWDsaNC3Afmk1sUZVNAUL9Ih9iKtgracK4cPLLEMpihCS8gW5xtZZWl6KKUJ/
JpiPN/7BFMKFXsKzmn61xfkJ3QEbGU2Wr2SQ6v+R3gfluLXb0gCT/12/RpI/XC2l
wTbFE/3v60SirE7jdIugxmw59PMnqR1TvKOxlOh9ukogYlpahUBFyAlrW09hR3+s
vcMz8fD/msrFTwf5Gk6RXByWuGC5r9SrWFXx1gnCgWll0EUq4vaVry9u7E0MOAU+
CJKz3mQhqIAQa0hUhtUFO2Xay0hkBDtaXIm5iwRu1kpRHczTXgHyp4PhFl6vyfB2
b/EN8W6KPlSZ8VHgdB1ZqIDVQlPrRf4jUGz84ke38WPB8aeAoAOOEP3EUAquPlgr
ZPbF7QUbaPUosZBwjzeqzOdGf/9kkWHxIusTt4J3gxUm85uAYke8eW/1GQKpEOdS
z6xm22Exycgf5qcd6wWBM5cbczX1mkz85yfQE2bwmFdgtG2TxMqAoOwr9WwDdQs8
csHS51OzcHTqpfGXrstHrlk9bELI+BnCOjNnkdgG8VBAzegcql21435Md/swGfUn
7Bf3jnRlal2KvFUuMv5JuVfOefW58nOH1hiKl3VJV9uYAnOjlVWzXNBULr6WiECk
4O4oM+ppR/BV86txuVlMcJh3icvd+2QYc5GoylJx3u2g2maJomJzKGcha/D1mIsx
BMv0vJaTuH9Ch4OXjYtnGZa1U8PZdMuvfFNt5ynCiNogA5SDIthfZL5w9D4dsFa7
Pu4EcXf+twwRRwUVO1h2MGN3jGyaYN1NtgECwTXKom5NZFQthDWRHk1X6vRndXbr
NdcvoVj8+icXKCcUnrtRZp/TwUBaGXQsAMA62dy6aIn25kwNfwnOA4Y0kLmLnXvX
v0RfQmhjdruevYgoE+uiAIq5ML4tv0ICpetA85rDiJe9PzvuMm0LPWoX18q9m0B2
s0+TMY0SW2CRRdWE3jq11SSldmGTKy3B8oo+i7yNWs1McjA0fiwqcwG57cPSe1KU
iI27yXozl84iukfIEp2LK0qW8F6zLD/xSlLKPcY32Wp2b+pc+2wvud45fFas1qjR
vfl03uI60tumxjQjUC/25MGbLgcHj7OIjWsqVTycFAuj+haDah1eiKwHN+np6szf
fC+r5dKfB575ewL3S/6HAStMn8fEL9F0IeG+nUht+xxyHfDTYn03XYhgtfmEPu27
bqrqqDgKhFKL/9pZMVyG6R5KBbX8FHxWR1kpB9r3YMHIeZ/Uh8RAn6IngeaooACq
p3pB3XlWHirK/rhBj1Hr/akBrnb4Tf+qKAdyf8EHQmTeRtFIVUOjArjvnP68pU3f
jvfAiAtBMwN4t5Hr9O8CsCCBbxCa1ZhYCertFtcQptBc4XansBlDJ6wBLQO2IuYJ
Yji/wlsU+ARHJ/E7r9YXuUzqMbTC/fZCkTvbWOJMxQOplPMFBzVT5A+BTYb1X9z6
f0IzC84DzF5cd0AQ1JBipx+kqBBsV69UkaOatrfMSpiC/QV4rZtD853hg7OLeCbW
R2KV3wdtfspTXgGN1zDbTm+YfKhtLuG1oXBCUwMZ/z6LxpCiRbEdNv/xn7sApHSP
Y056l9JEprVa5FSHgg+8S3lvm5gZsRGybFwA9Uavho9GnnULdTZjzHCdaS5ukDJ3
kw/r2cKjVy5ZnvzJO32h/3glTwrwQRW4ePiaXRJVXHiMZsAtAJ0ddcnafHPmcHML
9Oqx8sLwAWUOjpMKYvRYWw2N5EBEaqAkddO3BdUVO/1XX+yQZZ8LVnyKKnJJJIwx
YVNazhAeGk+W8zWIW/HF3nKMjZJjlagKr/oVNXS3TNO9UCAsFm3MeggKSuRL9D+K
vQz5v1esyjyAqP1nFHlvtebDGcUEzQE7tZro59IPjWRz4BAKpM9TmpLvh8XD9xaP
h9W5zYV09vsLDcSNxTp0WHlXqS2iUXIEqWcXnXsTEMjhlplnl+SSNlTvm0F+0kcF
ikCpFexbxX/JAEyoi6pHiJsEQ0F9izTbBMg0CA/w2N81/FQSBkXeY/3SDfObqbG/
wTskSZdrthCVA94ujhCZGLftLTzVhZSUi/SPwKer5aCDZLM6WREi733Uq+4ZHCK6
ar//HDU5Y1ndMrUSK6TP3XtoyslQwlU3MPc0fa0tQsMJQP6cnzVZrV0DduzjqZ6g
`protect END_PROTECTED
