`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kqjzewtqnEIi1/8i0o++3Aj2MVycqbYcmRtEhRo3oobk4bcLmq0+h9HsxxxOyPrM
KVUqbFvM5tCwwzjWyBT/B4YFBLKM9JCUceI6karsKBw4ZpJIMw4F/SbJHisiDsdl
XFnysj/D0x2XPl64z3P9thSQP/Tx15/3dfEYHV/KAQwuGoV0ro506ASCdzeDVCsh
lNhyrDFiQIf0qKSo3Jr98ZgGTi2awx8FNuPC5t1g3MPBLa3dWksBVyQPmQvUjcEP
9ABQvICu5uULOYjTwFvTN12ilp0cd1rPBqNsgO7pduwNgxAo7bTg3rCdxZy7DK/9
oxW2J4+rWzZr/he6r7qSMmmwMLXvx00L0XLk7RtjO0YyKQHrwmcofB0pKQknQ6Yl
oXiA642qbhNvBEUR67aARfh2ivrf4HOsZu7hy4n/EW7LpoI0W5qmhkJy1VG/C2eB
0oWnGVXQYw6xnTjzSeDovC9j8gMgSL13KIBr33vJ372Y/Ot99Sh31aRq2tuf8W3F
6N1Uk04Z02y6NZdvLYuDNW+fQKHxbfRTWhWz1DgpdY6cj8C+M3sWwh0G9gbhAs1l
1Qubt/Q3xMiILpvWl3+4mlQbh1HTyBOP12dRm8PUjOZyuaeyQ01S2vAKgu6+EsPo
OL8UJyjhI5V17iRKt0hrpDQx6aKukjpkXRVf+uXQIpIS/Bzys7UE4srjO9BancH7
M6daZIlQ3yHYhDo51lc1Cn1+Io4R6ISV0xcXh2zXYZ7jEozTdeEU028r15BQDR6O
YNWRzyzYKx3yetCl36ncGbFBeAs2+uTsI3tUD3MNunSrQeJAvGZ/KyDTxniHo9Vf
epBkNntqvI7zDRW3GXfErlGYOjzzwLKnYJIy7iGnnwUIb5R5sn7HpGwqdtuX21tp
FtHABT4RZRu6fjBaZYnVyfyut7uTYpEllrI6A1lbsvmj1tj8iZMyTJAfVhRPsxk4
vkKtbVN17PV4qEXmDpzgFK9oP7c8ekyvXJJ4wR7EzWeBI2AeaslnE3MQFPnuUPGo
9Ge1taqoBtvuooWrPJMXP6UUCNDdlHIjSOzTp4Tz92NZj04fzmNbX7fjw10TnwJo
ogMATpq2tTLGzVBRomfaho2UKeQGu/nXYcH0cdSBHme14OVh9s6FnkyO70B9RZSq
EBGgWiUSqGgdmc4WjJzCpgFAxZMMcpkL33m1H6dsmWvlzn6zU34mBspOALcUIRtL
/fW+P7V32fU6lGv+dp8JU2GR7FW34nHR/8fCN6E/e7ZEBeytCM7Sy2Vb+A3M4hX3
Ifw8LvBl+S0HXO9I+8JXViVao1g6aiAxfRqmYpFmLPR2GhTkB31RGbsm6dXHkAPu
VvKjYH6sod4re65oLQtPX8AIjaHBB+B3zbh8ljbzSpvNu2F0FHhvP8RrkhbPiC24
fsW15nnoHEB+7ENh++IXPtmjJF0B/EmM8TCLQdW7dY1zaWifPoFKhLViol2Xd1MD
OhNfb3OUQoDEkz3JVAsK3GbJlPlyDMsHDjnPyZ62Ndgs0AL5uNeAqqP0gghVsMBd
O51GTG+++9sW9m1hl6zd1DeZevdywjSeptjCKgqYMzDsJX7nV+s8vZ9daufXjKPf
Po+O3de0MAq5zI7fomy4TyFAnuuFLYVvssNAtmugXEzkJoBJLrA07uZWX9VssLOL
zpvVB28wuT5D6YekKIyBRP7obidpu/sEHk0dBp9wggSKl4GqY3p39fEDQj/PjtHo
pSU/EWL5c0XHsm9nuXyAOYAXqc2HONcpI/kSW75AB/xxuoMTkKPiILoRqrXgsy1f
JWcQSfktargMGIKnUIcxpi8k+T5BxUQCgigNzpFOrT1uq+cObpPrq6mMrkBkOFkz
arngp7xH9I22Weff2sn2zKcK6GYhd+HlrN0n9siYt1KbY4Brc/imWqltAio1FWZe
nmojTZVAG2G7Dk7eOZafFt3XPzMxzZvradiHa6hlK+zWRf4zWC9uDBMXENwW56QP
eTMj6JCJPwTPzy3XAIe8ndR7CM67km8v+sD7LKx3cms/o00qqwMaKCndOmRMOcOt
FcBBwcQ3diHflw86A0CAHjyHStmIFXcZVyTgOWWKF7PJTtC3wkljfysix911fKTR
HsDOz6C4l9w4WJHqGj4lf2WqzeX3GGUxYKrkN4/jau38D7Q8a58OQ+FoJKVqnPAr
eDrP8Ko17Pr8Dwko0JAvOH2l78c5TnKDRG3Xr8eBsi1LHNpwOHy5r6Ktb26d+JRE
QuLzLlBjEzXaJ7usqEWmh+QyAAo+U5gNs8pq6QY/zN+nj5At5gm/WGTUvq+sefM2
L7MHannppDueyXB/R7tHyKmuIARs8u107FvLNcc+f1g/wRf3rG8KkAVMC3RNMkzx
rg4MmCUrc5677wm26orY76bpNADGkQ1qq863qFE9+kwQ1NPrhVf3Vax8zQdJFusR
RtH37O/yIBCq1D++WFGGM/kPvHgVdY0UrtsJEOi9UPo4n9plQZWntHD2cJaRVvBg
OqyNuC11vuOMOQGgC3mgdBKuqmV32XpN8c3EMWKzgTLcw5eOObTgHD3UCSS2/PFJ
QQ7/n8diPQ1DeZC7UYM9uTehQ95M2Lw3GSUZc8YfJYwbL79zovZ8rkeJ6R3Oky0w
etzAm+BgYXsfmjtCySgtQIR3EIm3T6tdaQmI7o7xa5RHoF7H+xzp6WDDxYXwO863
UozMXFP1o8ExXqGYTWXpURLQqKUnlJjkfNVWykZBTUNkiuTT99Zrefn5zlmueijc
HJGci3Aj2IaZ1DuzUF328SrQFE1wPrgLAP1j8Q0vV05zN04HgHtnfFUD8C07UNN6
yiBvx6ek5mAiUBHYZ7H76aUCrydungM3/B39tU8mzzJc768ViLpjwWoBQd1LOWSb
WaUQKo3Xqcgb2DPXA+krrGnv0nxer9jLx2taz9g3371sL2vpZ64OsNydaPYJ8iA/
EtSYGURV+aYju2Op9rtXGX1N9yTgRIioMJord3X6NOg2uKRcZWAsGUfu4bZSg5tZ
s4Rx0UbN6qJOkE5H1jhLzjSrh7MVWzkswCMNdBkIGe3s54FhP9xx6sX9IzO84JdW
QgCvTlyuoqVNwL2QVmZv4ROtxfmBgkGl+UYssY8993W0pm9gJBJzk02Q9PWbGXvW
BV3Xfe94i/O8yP8vnQEdHRCU6rcjudDwmggBIslj7h7Kv0ohgEBtdG/kF3GL8hjb
qYuKQMiZOwmw/p6t/yWOJlSYwgHpG/n2U4l3kQhkD+0Dhq5cXAFyJ5NrzcVJZa2/
Tw4zHycKTlzFTFgKhS5uU7T5dG+a6dMPL2wf6tk3toECTS8Y5GeqBGntNsADakDe
euyrunTdtGtYuUyddJ9k4enAPOVBG4828IJrW7cgMXVTim9VW+R0wHpew5p6/89z
fzGXKQ1G60FCN/4NvQNs6YxU9wDgD/ILS4014yhQ7Hn5qKOxKwZ6wKrAEvpYBP1w
XqPcADL2yHsZjocVlTyAZOjuLG92esLASxoF8M9TsjIdvQiVBlpekC2s+K7kgb6V
2Qwl0TXxU7IyrbkTX3KP9pkhxOCB09zWX8iM7+AHib7z4m1Fjj89s0PellEt/jIH
aytIxz330dqNNiiQqL+HojozGg7PUnd1sCyTIaoammY7JhgNwdEP7cu1efXMLZZi
mcmoUMdMhoBHX4kd0nlllfEoFvk+/xuC019aIuFn5BpkvqhstCzyerW075+UhUS/
NUW95xQ7ppeyD3t6hIihAJxYS7eq4LO/C2LNv0c78KSoK0YDu2p9or8qnwaEZAJ1
1oiF86a8LvDGPYonA7hoO59oW/pnLusv4j1VAHAi9PAcUvwnJDNy9xWA6FcGQp/t
HdLCYQCGquixId6pUrqEAREjI9TQ+88ptMneO3B6Wik0syorhaYm48bKPFr1oaWp
xxic6b763FBVlFID4PXcoVJsCe2mf9KisEmKH4y5I5hUXREnJycasShbPXs+Av2Z
C6VwOC+EEKby19TcVmimosMBBR+ZAeSmfyvlORZcbQYIhcC6dVrZb0i0zsH27rNs
pPef66zK2f8PcE4L2KlUuI0GNcrR3zeOnP7E5a3AksAcqTKLqe7RuNafz3a6NNdS
I78kzcVhVdTfPDvxORUTpjsbudkvhhzukTZDQRQ4GK/AhN80LuIfhZzRWQi7IcN9
wwihHRZj/ipweUMBu9pDRjtakyw1lR2094xIeaBiTbsp4BXVs5C2hJaeEwPm3VA4
LKGw9lXyd5vvB+T368dbrof/ND0+Q5gxT9O9jOJotnQgSfJB6HLS7cYN1gFjJMbf
TeiIyAlv8MOZkXyPcqOCKs3jMoxOPgHpwkgwBApo+GvLDiVaTTM+WpNQq9iW0BIU
7YOt5gJpw8zQPBxwpB/JgLkx64Ef/0MBvnQ0snGtjRkJItgV9gFh1mKp17r8TCZ7
/Xll3G+6pAFKKeZXC4YXTadb0PHbzeuEwKvGJAqb37dRdNuVlMvMt4bROibAtIgN
H4fOA8PAF+HQoJdgMJsib8ivwWL2MU6JcYB/GS71OIjuu2pP1Q03+njJHzXiL2e8
z3UOkVdE6ySEKm3dSITum9yvIKe6l5kJQJh4k3DgOjx+IfvMbAoZ/Dd1tZQnpzwM
WybSORryjLsjv4qlWmsMkOuGuoR30nWxf3ER5iii/WhGw54grXo3Iygfs2cypBHm
btgxP8+wbdMtElb2y0pnJ5RA/G5MLrmxoAFN3MxfchlHsg2vuoB3gmfbmCIwuqxE
u2DJSFjvkX2zhelMAoFhCXMnhIXpGtnWhKwoJU5gt6yqHkccKdHnHT5mVzd3rIvG
CbDT7etXDPl9LTrsLs89+T3+WqY+x4SlrP2SGUC6/FCR/ZhU7ogZLafh0EoFGLHa
/X2HXWXT6FEdtuJX4TY6zMS+Vc9OXQqdJ2M+bzhCAEP87ckC53+nSs5xiKE6F/9i
tIcTUyAgOg9d4MmMSGdpKBRCqRUNKHMl5S2t9tMMTo1Ueh5yfmOmgkgCTSii8Nqw
pe6NkaxoU7WBIYpgdfluuoPHPy6XS3lUTC1gUk4jwrCTXdTDSetzJqdaRBe7IU4G
hXJ6W7ZIcIranS3ErMsLvWT132PrUg/aU9CcFdyuiMmh+PVaDalxk46iWG+HvpRD
9/A1O5fkslO67I5kXs0n19nOWsbth21bQoF6JmNH+w9w4b9MAjeL0DNBxKHPekw0
xFL9QNQ0hOLAqmvAUvvLojVZIqD1wQtG0s+G2Lh0XP+HOIVd175nkG+VEqfdEl5b
D5A5aFe83mYHgj+wBObDS24ROml/Gl4SL0RW9DNcDcXIkwc6IO//zZja9RyhAy1r
KdM2zlXIPT3W2BLI13pbx72S1/1V8sxqFBJhgOqKahLhzueFMitiqMeYRJnEiG9m
f30FL/a6nvMuoXGQX2axxKYPHEz/P3p2OhlzTTkrXPCHb05/swrFRWbVdkoHH5q8
Sejn7nKQiahBrX+Bgw9hgm1XkaQg2BK1mrGRpP4+LItCj/7GBI/6CCOSzHvnqJKQ
PC4rfXvyC9Yp0ewA8RCfLKAbq27D8MYnBzrxzSXUL2z9BVywVRKjFDOSJ9dgnaVb
R1bLYYuhIfYvCwnuIRQ//KI3DMGIjbSkyW+l3ggKj1iG5ahpb8/pYYjEgsjyuXfy
hChzRwAW07Tqg+JwktJoUIjumBTau2xVEamSs7DLlhtzfMoF5L85Y7HpdHZAXBMB
bvyU0XIouxV/61F3f/1TDDGhH/grifB9axeog+5ddifrZS1goeAAtOl6en/z25dJ
l3Obc5SK0FL8sYvjdWIrZoAA0GGigugw+ZQAnPJm2AybSJlajkoag1ZLmuA/Op66
yQakD0m+5i/6dt/SgEDpiuG05Dshn1c4PUuA9Qx4SP7YZVWtV5BIgXWrbAB+diy9
W+sK0/GR2d7+8Xwwt7esIr4bpIPFNVbGqhq7Ocsgqtz3y4C+sof+i+PtjlUbVfBB
isBuZXNHiqPI/tEAc3zpTz/2kikQMjl+ZSnBQUyoHQbjxi3epgmuRiwdiICC1K5E
0zL6WoUbcsbROLhvSgKJS7KoIxa4sYuM8EYLrUr0wzaOw+4b6S1bP4Q2cCLxE3X4
t0sKMrXw73NgyWDnUp4kmp0oZXuNCnpkeyz4aAz/59HsMqrKvoQN/z7Nzc/ItNvl
tYKlXj0tPAYYFS3LuT/eYDxXSeRWSwelU21O0hLBN/+BvPfEgy8hKwTExCMeOBFo
NuGC8Hndv3Q+L80sKqVdJuyVsP/gXH5/T30W8XR/D5ZCb+Jr8Akx342nqFXqfu9F
l826HOe66KZ8OgOngqA3fPXdN/AgLbpQmQlUMQvtJxw/bD8oa8ZcKL0UHV/mTR7v
OT78wYsg7W6SSksbX0OeyZZDStoIrNT+ozSXbVDjemZwPrn6a0EtYpw113y6UFLc
RLUGtPsbwZ9E+5Id/nB5JSz/fxrxoyARJYepoEz/Ujw/rLrpXFrJt7SQ1TwWdbJt
C1+n3iqvmMnupOh3czdGzZxgEEUmG4x4SBkLvv0YICvPbu2K6+MkZlASlbwFZfuS
QrBv6fJC8dqL9c3unI1rYCawaT+EGnqXWlaeYiO8/kIDVoKM8chFNiUar4mH2aip
yPxYJMxLnEHmCwKuhIPVRKOM5xCoIv+I6P/JRIORaoUtGj1E65DDGHowI9vw/Pue
vXII6f9BF1NPXtu3awIJ+AkzWXtwB5OTFtm21UbW7yGo5zyOtvuPEkIdfLiKAmoU
u1mXOuWMqT5yEHNNGYhC/c2Xdy5hyChQoV0EOAvxObf0yjPGLNu3u71mfxi+8phK
WmTeDuaWgAydWEORGEP+G+jyL8lu6aIcGKkRZGunWcHnJSN1QIU1L10sanDIjwW9
cWX94Fj/Gwf/THhID8OYC29d1qi7AwWo90m8mbeVLkut1c2lGAKAOeCEHe+zKE8v
ncL49qRsAz3z5slNzc02P7LbgGE/rfOfuggKR36W1g6mS4W5lhxdPRd3KId7U7LS
mKCDrzCy6BTEo8Mj6wNN52xrG54IaMAzAUx4x/Istk+6Dr9rjE9MVdEtGDRvX2Fw
OZMMz62G1kdQJEjo5h4YOw+D7MgOkhqEDe/JZexTIyFC9/urmDIfYMkzvIFEQ0U7
acEWE06K3VhMMnshDGHtrpPB+P6eXaM4CvUdsP/JTCv+O5i1002zCtvBNOphEW02
hiM/vT0U2m1lDHPuxA8u9qvxFBO43jsRFtwOvSI6jUdg4x/i6P5rWeNlqrMSh9zP
3i4UzNqZ+2T5gpRpy6uwC71qPOP0sWJEH58LILy/pXUiZLS2vtOJjYfmKQAFMCiF
kRgPdq4/gpUVqfc4G+L+WkIwmRQpulseBGsxYxLRHu1OWde9v/oqGrCXUsleqCN9
QgOdyOC7XsrzQpu6JQaF/v07KkW/kN17gTgqtMAKizKN2DH37Zr9BRKqGPl94/xm
2sJg2HOwGvNVMa/g3HpGLojoeBeYjsB1nBvulKqAeHzBzXyAoxU5ykcxMtjl6SWi
L4d4CUAYpqfEimCySTkoOHcwTF14VeKeFlTXn/ZhTjM7yMWbRmU8wL8NNe/BiuX7
WDA2g0qfHGqmpXyDy00qAAQnLygdTAav3fWvad5+oJ2/IcBNOUVviL0dvTTzLJ1I
5LVwuYXRALFVDW/bBTPbNhZnnf/wDQaXkeBclMGsv9jk2LQyMxKFvQaWZCirnu+3
7XfYjURUGT/z7azV/n/8EE/ZSPHe/hXeJtViy48ajasUjG0DUG6A8ZOmpXXdKZOM
YS1i9JGSPqd+yzfoKGvMyShiq6Q8cAluDBgyk9s2YfSM5wC/nwQph/NW00DWK7dk
GLD492I+fdbKrWX7z12hVWe4I08TCBxfbGER5+N1Dff4LZ8wGsRO/I9QOjH/C9Z+
lxmCqPpGvI3krHvQ4jbSLr9e5dKSMKYYScX3RyARZ1LDv7I9whbq8yrLYaZNchrJ
v3GZk2m4al4s0H2zvt4N3ocIzPAGjHp1Q8h9nB4x7HBXB/CX/brMzlOY4em3esSF
J13EkPb24jhZiaw+B1oUq8jnj7xwdY0aqjsIJje+042QOctgw5K7FtlEmf8S5IOt
0709ZsIb271HkdpuZwKkjKMNSUGGJ5prPgfdeIXira8nNlhKFWt4whwuGCitBmRl
xnu2r+f7+T5yoEcBuZ10TebEvrAJpHkiWlt7DN35Uvqf58/9OO5EcMATqB9fIVjH
cRC0T4uIVdI8R8qha+lGyuViUhaOfZSeDkFDVYGBmdPyQGBW9Y7aqyg73UFZZ8UG
0Rt5uFe1J6NMlX1o0HWl+BBlQfGcpEBStaHa1x340wEkSr/ul6J5dlObKemfGnH5
dLn23FIaR2LgrhWR7KP/Aix9vgohsleae14INuOX9O7Kc1CM35yVx4cdXVKEy7eK
H+M5sx8HKlrQCTd92+G34tqakd+IHjXB0YIYezLICt+D9ivYfpA7daCB9igWHomY
FOwgDvcFS51GBEQuKnHIIIaTUFJl/8Lfr6xYWPadUVlVKAT7NxV//tvkfTEMsbJ2
QSC/61nKIaBBTIH9upm/QEN3QQHWG/w36TeEpsVm5f0wtinNo0bRmYt0UfzPKSa3
GwGLzSfUndBpWuTdrDRO1ZImUdcGWNkPeKeHMRxw1T9G29CpvMqLmQvlPTHB2Azu
5wTXsDSE6+g86ayZqlzODPDPwTtz4z2w5SKAizTfbmz8pU1KnDn5GVWAZwdUkfXw
tcj+THqcc+GRq141LGrBExnRspYMKCNHcgBEh3vmKhK/yubHstR7YiQAxM37+Jqv
evIhkBo5itXiOZK8oyUUyrJJFV9LJDZjofYz7TqiA+t+xSAMguIQ2eJsZ0Lqr8qT
sGQl6ix0rKQtjcvcV56/ULGU9y+0QFwXOd4G1/iIxO0aJdHT2Z+HxQsR/Tb1AW7R
nu8ZyUp66DBhxJH2PVmomrFTR9bSeyrpjaEC4n0+DoOKnSDQf/w9WINQ9usubl8o
kBHYjfFunK5jX75wdMQgCXeM2ElqEaelqlADZfhLbc+YKAl1og8+nMHgGcjNgB0s
iZVXK0GM8owVJHX293ZUPbsL+jvMFz0XCprx6vHoM3nibQDzmPfz8cWTbqz5hG2a
b4E9mbB3suOrmTQeANTqEwY8pRJ8jJi5yDVibB6WSFGtEtc+H0yr7gS/Oywc4Emw
o7PjfotltdpAawEnyZH+kPc1iajHO+GbS4SHLVTDKR3UuZCaTbffCeGmzNDt3Tew
RF436XPiuvkQKw9HThdH9tdcs8fav2dvKNNVJqDeo8eWuPiwNk6H0ThOWOe20Rao
dMR1AZqps0TkWD/8K64jpAYCImCgw8+ViZIgLEfqHGzmo1tsc31ZyRtjkLSRIQAM
RFQpIsvOj7cJ6DxMkNOIQ5J3VHGOgdwjWTzKG06eg6I/H2tUpBA2uB+MmtkFP8rQ
07gcIvCk7e9ctfv5LM6c+GPZR6lPAHUc3ygt0MO1TbTSnBf5xxQ5iA57/HtSYz3T
ATNA3RnFLjCLh5eyIGherWOuE4s8N6RHCVZEZIUr6Ss2x7pdyT2rLvtPrpNWCsWZ
LrwNYKjJh8wLpo8tZ9aDeIwFz6E+rjmgMtDEVTtFhqwGcighD0S0GCmNlbl397cs
qhDglAzuajvF8/A4UrKuAbJd5Yc7xN/tHwxiOwL+nB4H2rUCAWgzPLTWLcKJzJLI
GVwX1HkAdLD6vnHnHysYH7W1QI2otmVYx9Z1CDwXOxEJsithoNTLL3ODXjMMtLzv
tfGy9RZeEpeMsryS4Ac8DzSWm4++YMofSp2eQMovloIq7DyWwmVK27VSU8p6r/8p
clnxcZ7kzLGrCLRpZwck/BGNDGOU03rcfdkQwubzfWprXTpxEXdQtZ6wQ837L5M5
08P6NMsW5d9whOYPktyMpgx1dp49FdpIyiJLoDwlrNTsYRICVY0JoqsQ0JiiWpce
yjN9WWA5E3zfbfJISwz+X0VaFSvq+i7UI6j7uVgw4FZmrO4BB2ODtKLD+2WIcvLF
eP93o/acuDAyDnRjDEmIfWhGy6biGwQfGyyPyyBqmbJGe6QS3FtNsZV86/ut7ONu
Z04dPjFdO09OQaB5+Of5DgRuHGPDgyZPNBDy5CQDIXm53cy0YEfVoU3cGsLdlZeo
S5H1Q4EE3yl9+CIvRWpnqV1QlnOHyiaQEyMZOlAZvsJir3CzXmHh/SCxowTbTYi/
tEjw3gEgNnnl79vt4w+GTY41w/VBUZkbGfnGbhXj2gLyAqg0pRckbU8B9N+s46c+
LIp+78uHqcphkeyRfIs+zFzBrCVOaXRmXfM2o2eCw67KDd6PJgD04FUzY1x8akLi
CPLXV7cwJxQ1v5oohWhm+A3eFkCWHrjuvd1Nnq+Hq+DZtBMAxJiW1A+FK/Y5KsV+
+kNwGblr51a0+Qjw4L9/iU/bRpKjrImT10lsIgBrHiJrYEl3QkqtUuXtfJuQtLsF
/Fcrv6MiPPcIAFavfgq+YdCdpjmWSH2Ot+OLaABBdZ4ddvxNvNJ/stE6sWcPQFaE
Bprkqf78upOgW7vCBfL+1dV/efexL230/rsLJvm+T+f3eKYbwrARj6ce7x7EVWRd
FRy4K/zwgvQ2unHo9ugVCvlcuXQ7PtgdIWJmYDdZ4gpi6Z17suhgnmb9uBwzufrA
mJAKWrkpj3dqq4FeuEQEMMfER8N9MbE7pdZeVpfkvQI+/W6WuXzYAfardqX5Dj47
qdxkRkygLe0iiQZSuabWxJnAMTPRSOq3Gs5JY7xMFRBfaNEWFT+sxEvaIa6Ej24J
9FksNoc9RMowuoH7A0gRxxpQO8qvn01wqGIHRV0QbJCpiU77jfY53ChG2QeUuDBc
uQ9IW+UyiteXEq2NCdauOvMDJr4SIKkCxuuoFNkZ1utCEC1qOldDK4E9end3HzV7
HTdXTXQMlwaGuVJF4pEkFyef4a23f/6HJ6YtIl0+ehCQeq3DWOwFGPPwd68UAKnn
KWDSA095F+1tnSZHnlGvJvXHKcXtNdmpUZsXGObV7RjxLxrlQIWAHXjfR4T5/L29
133F/Z8R8phnQ/RTltETgNqP/XCNvIV9nUslxmEuv2Nv7hVKX1KYRkJh1gpARGtl
qOqCOKoqPOwRIxirNIQJY9AN8BP9RMzhOjCYmJEj//36q1u8wwQrk3HwBBszSvDA
q0Vi8W5so8JJoICqvE15Kie47wAhwGrrq5gMwBjvWtUT/USP0oxkd1Vi91nSzWiD
F95QuoiXfd4kXKVcMnc26osloqeLSqGJbB5UZaxDPGRvhdrBrbDDASV3PcmC/Dtk
sbU1DtXNoKbHq8If+RaUKett0RvSMg2yxkenHu4dcHmWBlNH9paNDN7PrGpDGeFL
XbQI3bepte5EpFxyNVM9R3CYhYz3gw+OiDaALAsdF3keZTgwQgZE56QDPHiWhDkU
qKRHGqRgDRtHcG0xCmo3ELGGqajpM4AJFGHQ68hkaKsfxUjpouoZ9XOMnnsDn9tg
9fgIlMxmMJrPrGmzFfD09+ypo4xNb8KY8igkIgX/JON6UsCMV0/bGY4+ZrU1c4BI
4qUPRPqmKrh5st3ZILA80s7IXavuNxbyfRhqum/z08YrB7qtqzZy0dAXohAwZRrQ
OSFvfTedg3SsEjHXGTWjMnpyG1AyshExlwcrmkLt2bSz0ZxZy0zOhaKnmfwBQwOt
BMZUuYl/mQYtF3xOXXuGHCLT2/3bo3zBeC97/xT8CgXymb2WSfqoBzh8rGItpzcr
QmANXvWJigi7B8N12nYt5KMwJHnu76rc4Q3BdEwpvXG+5xV1uu9fr2MHg9pHWh9K
XPAe6dZ+h4jxw/R7llC1DOqXS7A75LHzKg2jsx38C6IfJzKpuktGyjDqEGFal/Tg
3zfOva2IWP6gDChXoXpNkHY7xc3BL3fp29DbUTkWm+QNgdu8CGaAnJHrDSnfQ5nq
UUhe2QYvel9BgX1P0uG7YN1ADcsR+UTyfJIJAw0+9Oy1rJdIqyL9lHNPQxq6IeE0
XzOsw63nXTwDcjZEJsKZNEX93DUGklDa9YCEEMgINRPGm+eLBrHILlrunTRIALOz
I0TQyuUK43lPqCh5gPIHmmzsrfEBbHnNPOqD7me7Cc2GQEPb/fzRGm1sEVL98Pp3
nmZrvF2Uhf55TSK8sjJvLAYezOkR6LOu4+PKVIUiDOtbKAMmnX1XE+k8JLWkuj/F
/ZwP63G9PeAtnIwJEddR6PkD9XI6nPwpdDdBu4g/+NR9LVwnWt7i/cGZlrjcUia6
3EYeLlZPx+yioalxTI4MmlSzguIsv2eRxsmk6HIGmxuHVPiXsHc0nrT+ss4lK+aF
uaxOdoPr9nLaIcc732WEOsgoW9PmXDNBkVmgk0/ciffFPTPtXR995a6P/pQGYXVK
PUYm/UzsX2koBEPG46H2HdqNBVu5Zxa2yqxO6H/ZBq6Z2kvaFxFU1J8FRuvWLq2W
K+4ewCc74AAa3YWbGp92ULX01J+9YtNBY27CY55LxmTvjVQ/WJOp+DYp9QEFbWOT
B3LT/M7YFCwpQL7o7Thkfx0TjIUqBexqkoJdv+mdoXd/ahw1keYJcNSfGp2kabtO
Kav2os71/6HxSKVnDzzCLFv5iWB6SNJJf3jxFGKR1W8rla8Fv44lSVtADWAKMA+t
167akuX4+ZfTlGyBPED01ns5GJFvs9p/0+09CNs3qLSTcuvfnWAyUNWzQrEJflvV
F8azEEcaAU3k2jAM3dvkGSLJrhqYnMyOzgpeXOzoCrFADfMZeTvmQd0pg3HIpTuZ
OpCzk878M8caCXRR8iiP39FdacviqEdMFgbX+mE6QeKgAyfsHq0QR7t3lu+T5jh0
GiMf86NY6anHIemP6LOl08Fyjzmjb4uH23BuWHnn68UjB74hNU7inHMliL2xy4lu
ra+NEjFs5KaaNQrukHCj8Z8gFN20eLweuBLN0iKW62mNhatywXJgttP3A8mtxMbt
Gz86TbT4ogiarUoyCPDI4XEhqhAeGxVrzGp0aAvQhml6OVD3YYWUA+xY0aRvg5Y/
DZ7quMUINUOFVe68j5ALmnCSshfiRdgJQ9RiRYADtju+bjuHKLtaz6nXTYyTlrGY
rZrVPI32EbVymBveAnhquo2ZfsAkGWOiBclLLKYPeMa/FtlRpKQr+Ml0MSKKLow4
LYaBJd8AM49Wi+hXpzt8ibPb77ehFHceMQNkeSHqTuKY4C+ENtrdUa79UQDtZDof
yshBCi/QAZIKBJxjQbxMzgr8wM2KeSRbPgJY3Y3IpQrM9i7sD7fHtL/ubsVFbaBv
0jgO3Em04k/pAbB+eogDHVjiEV32QKcEgcP/FbN5D7NW3ayQS3PEKNb0PQ2iSL4s
w6HxZY20BG2gffLLXYjlAs+1W3TYIgdOQc3+EmwG9mAFO3ROocitSWaDn4sepoXP
ER8Oww1ik0Ai30bsfg+FdYukr8Gy3nAIA4gJaOEvOKndsaoShBC4UBpTx8VvkXAO
k+Iw7Jn7lf05//7T8sat5BIrnRJGtRzofinkgtd5CZpfl7kKH4V4d7B1zULqmOkB
X7XcRGBSxt376PFVCLZqmzNrIJMvEY0Ow3yTat2gOuarZ/BErgPYALDg/bLZbIMM
4yUY2ytifA1eevq5NgRWpbwJNVs9BsJ3dsF7XrS4zUIvSEnMgXlSY2+wMFLNCHPS
DRqi6Z86K8I4qnDN4kUce0yIG8OAV1ukEJ/7Mr2Yog/km1c/mILfdflLyrLC9Mu5
B1MS5dJtVAXCDzxw1G/ClaiEdoGwdVvWen/0yjVdT7r2IdDMXSfuKB28Wi5tS+vM
CTzeeQHoH++wcF/PdNzrO4vVQez8yqmRt+piMVqCO41udZUBcuK0M9GBccysYiDZ
2mPAODPP3bodze+BV7iczVDZnQL4YqcNp2kLrS6NtwdnhmfJW1FDPdiFxE8vW2BB
c+gTZls5NySkSaN54R9MuxX09hW6sM3HPLZx3U+Jv9T40OTrspTziPdc2ds+qQNY
J+b5kCLyPNnmpgQfTUr0p3P2iyYb11nxjIaZ9H9qgnh72oN+JEm+T+xVrauuqLCk
C1/LdOomDOyfYlJ/ivOJRSJ/bvhH5yYjuSkjPQB0Y/2bnZS74HtNxUsw1LoAlPPf
4E0xUkfzKQvWvfPYsMCwIUlLTVfEDbPHakXLBp+DrrrxpFXgXhbOsJ6isOJVXNLT
2QOSxhvnl1MOZZbePfQSD3OsqHb3efwdijjwTQCqvhN66qL7uhHdS8Z1pZ0Ti+ZR
LHZBZRcGxvohDm4KADNazsLgfiszHAjWanpktyiavyTTzLgckZIAPCuXrhRBXOdY
rUkl/LtZGdYGYn9Dmzg9i9rZ62g7ddI7nr2iNC7D2Hi/6tpxgKUvebD/KMxtXqSl
n+8XedaIR0se529Vr063BCbnDEQ1ebkO0jVNv+2Ec3yU77RwllEl5yLEVpDgZs63
TP7DMg5kcxm5RppqiHu31jqLXV6Yg6JELnUP4Zb4s3tcid3mw+7Y4uUPen2CZIfB
5HUkcmZr6pZ0ONl7Q+7Ed6oKmXWZhStgDV9qbrmVuq9ZY84b/4VW7BugCiMyxn3k
SfzwQPE2r18XuKDImcUaDV7OCyaoz0OwcjPfztm6xAClBbAale0//ur6Tw3eoGuV
upmt1k67+BDTEUfNC9PFIUoFqk6eeOCppr8jTW/vmpWy9+iBJxaZGDpsjzOK1W+z
2BX1E6bv165bRzOoUamnBMpG4QCYlvBIP+I7Qo9krLWFaNvMVbm4gKNLHWYJ5ZfY
Ll/ABPw1qy1wOvGEuECVCz0bOH+JutrjD45+lAuYsRXng3nRLnOECPIzlqRe1gvS
1VbB9mk17xkH/bbqTMPYSqEojxxmsQZ0oDxFvrAgu5oNHW/Jmkoi763qSAOHDx85
t/NuFzGhEKffaXkVrOB0BwhjR9IVsaQ9tJp9k2EZcf8fLz6Awew4dsAxmbSaBPvF
YMyaMTMMNYpCV7h/tqQv5fOLYIdl6BsxJsma4jUJ1GV89Hj4zvs3QDDhPchb7UX9
on0MD12wdpXDuiTpo38KUJ+YCMKzGT5N8XFlOemGDtMfgLvp9FOgRuDSC13m4NLp
fLMqU0/NqpCswA3H5plTCgg9cgYRHoXjbNMXUY2dBVNzFZjlrQRFG+y++CHOGpHZ
lTTjTFdQnzRYmFh0MwPU8B47uX9Q1v2yfZ9wAmYAFor38VQ/thcxwjwq7kwPf1P3
UTIDz8azmTzxmU5OpvTZID8C6fGSO7ICcvsOjYZ/yWHzkuJQ9Z1sst4TqMEvhEU/
73ok0t56JGo/VnvlnpEyPw/JbmwZUVpf/G/vOqvUpAZ+vi+Ort6QeCN4z7KZUYYX
+BJRaBDyXOwmqxQEcQdkVBM6noxAdRmNuVaXxoeWXsAAHSHsazTwzGCaLuBzE8hg
xMe+XyMVVIGtS8TabZXbtxaS1fNnsG1Ch86r8Z3uueykWksaE1OSAUnwvswO4ihV
jiWvOuRe/YhtZLjaY3R7G+cmd7kSqLHWvvfZb/LmsxaxGv1z1X1hUfs6btbiAofc
nvnSIYrfs2hK8Ebsyd8zFj3N42t2yZqhK/cuntFqzwqSxUplIomjJh/5xmn2H3Dw
Zqc4KnOKzVmg7DTPCfMOQOU+u/oZ/MZsFOnoOdxrcfShq6I5eB2GCKr0k5ucoMCg
jBxL/eJPnQjH3CnP7emNcdg26+Ufw0kKt5N51DeV2u+gsPvyky93xJtlRsLb3eHS
xSzL00EJ4Wg+8owiTbKev2wLMv1iFs8JIT6/8qjS5qMAe8KzTI0sNLp1s7v25Zc8
F1UtpKwxEsA50tnQuykGlcmRiTiX2LpYOOyZPowVu58tuy5vi5BnpXFPbFBJDylc
7YYXSoh8bF8fkTvlxzVJPXnKHMyguDL2x/UyLNqLjgGmAuqxe6E73rDJbk08ugep
ReV07Y27EKr0W5HIEjRZqFscwYJ0YV2TNbn3s7uv7xM4g5scfLA26MOoKxlfiDDL
KxhoNB2TT5hVKGmZyEm/jOiRCtKMwNmwSOgarG+PdEZYIQCm3CD/eS8Xv5vgDyJe
0pjzLoAOtIoyDOQmakvYuob8JqHKb2Ptv0m8a7oF8t1M5EyfgVET5009OYvTFJoQ
8h8uq9nHKlxMXVH9pSPzukeDEfyxTbPzJyrnPbvc6ubqVsF+RarvTyGSmyMWdEOK
bHRdkQgo5GAIkGj0M0B5ZdFzuwD6niiL+1GtoGNcQ5+MFoKrIioU+g1hW9nyBnpj
WiidUfw7AiHM+qIV1n1E6R+vwbdAUkhQ4D6q2mT/zveCxa5WBRSt+5nitDwmTcVi
J+iPHUnJggny+POLKi4FSFWwxQ8/RFsh3Ps4HS6mKD5sV8ncgvXTfCirI1Po7UCU
CDi1tHwxL72ujaVeZ/dJaOKLZlD5DKbpo0N7nyEzcPADPEqvzA+d+Xv1cz7dhaLf
7wH3YNsUK3yNAkfbHHxO2RMSBPJ/04s5WHywNG9WvsIhqakMtK4SOhlwretlaRNB
QmliXlMVrUMv7PKw2qkRLNJD1R7uL5o3gkF+foHPkwwmFQ0tXCUGsbR15suVQFci
9upHj//Y95tXnSdVjL6WxtYdKqR3WKe2rxzlS7IF2xhd1XSkYkXkiRhK+NGBvULf
MK933RblkNtxNzeYPeI0KYsC4NyxvWjcnMjERYOqy5zvkwzyU0dA0i6XAUa8gfoc
SPcqcBSpV5+VSQixiuEx0eokhduanAH8pceaUAysQSsfplmU/dU2bxkZ12CFlFmn
3F7qGd09VsOjyGShlEhtinOBXnJVPkGOgd+jXMf8WrmOXw191JX4kc+EJKFmS0k9
veMGaxETisA7TDMYOFLj06lYodj31M7NxH9vo8YYdMBsLBXqYVc+JnTJzpAMC2u0
62cIiTdoQ03KdzsWIUocJuFSN3B5HShe67NG0v28vl0f7IFmZqcx0U5rbxEZQq/o
icEo7lDJDHIIKBXsAGuDoILDCO8snfYuju1/gbljlA81CXk7+0hV0dvyKZi6PK7L
tGceCXCek1ONOcqLJSg3ERSXvygXa+ymbJIEE1TYNa/qZGJvLBBN2JZKxxjUJXxl
8fMQZUEKPcrvoEAZqyP+iFSLvt2GAir3CNSMsV9BDLfFG2RtPa7f3AWfkwNBDIaG
3E6yW5zI8MbghGRinpvWfrXksUEZ0ny6a/iTauzed2mHK8o/a65wJf+yqsf2V4h0
ShIERhfzUv9a1KxJKSqd5fnCBt+6Kla3pKGEUuTHsaGHFIsKj3qQWS8a3O4EtC17
ThLCID38j+RJVbnz2IYQnC+6ySLuaAathhat6Fw9H0OOVNrSCH8W6yzdrzhzjpbF
DhbGRQ7ZpfvZ/ggNKQbLh9qPL0d8Hvg5ldHsbyyHH32tu1utrmBa0syaEJDx6mQE
0myZb21X0fnt3b29gjfjP4mo5J8MZLEZEsSPKPAhMutrpIRnpjPiD95ytAfkuBR8
/j5KOLjkzQqDmsakTtUcC9KZiMVpYbsV8xBDTmugdy5BDKnIt0spJpNZY6JH3I3Q
auJmGnAUebM8cGdZ5WtaD+QQ8aHDlA6nd+WkojJfd69+KMXFXpsvD5BY5/IDbpqR
MPonz3OM/yPPaPfq/gYoP1jFnQ7eQE9xfQmJmMgtLvBRoS37N7B8ICpOaROSOG4h
3uPBtbWhpTKEUf8GknShu0E568aeOjKWfNbo5tRu6YssUhWmmglDNp5jfDcBT0hh
FFLiQRbBaZheu58c8YKPyP5JGaHVFm2eBw0pSD0ySOOPs8tGvL2EboiVo9U8ELvN
ymvmp/ym4fGLAqDYUZFTqS+v3nBjO9mGtNuRibmZbJScYRHI603QE76cSrjgJCKM
M9vYNnzyzFwptRJYlIZcj1Hnh9Fbf3mVY+PkqufQ6GvI0ksQxC20r1Oyt9hxJpIG
GoM6EVwEFLZhk8BOsQIPfRVZotdbx2n7+cPBlUnM1zA2QiCOGCot5FW6MKvSLk4y
1wUaL2x01OAUbWfIKo9lMHAyThIZzaubwO5nJJCjcWvLvGJ2fqe6c4IiovSsa1Gs
2GhPotzImple/EF9f+GzfeZ8G+gr/zQ+b06YG+NtbWzBnWIVxZ8XzldwRo2xL4U1
juNieFvdd0lqApARKTDDwA8E+BYx+F7pUMUOwIEfbtZrs813xc6GceRKKJQL/Dm0
sGIXJPkzzJjLpkHr/61Q6Ik0dmHw/YXrdGj3uWz9hGPXgW8hWespbUswG2FhxB0B
3kH4FoMJ1wAyyghiAVWifqdQ/+XmiGJZzjVqVB0YXIIzlZQHIOIJbE4RKMXzFvH2
4NF+Z9hkWWZgntOli5+hh06wODaa8cjT39w5tnjTwBVYTM7f3IoTR+35cxRrvTZ7
kyANQtmOmiVr1ORP4JkIBpI7f/vCK+WZwWZQzKZbyd0c5lymZwzMGdSsQuru88iZ
n78MmCyZVXpoHOpuzf7B5l63sVBAQNA2+y69KYvf6qlqVmJEisKaLVbarfdVD1X5
CXuiCQE3lQ2cF/sGBf6yyE8qV72YmhJkHBNQT56f+oCD9Yzk5s/PKaAi2YvqVuxO
oPU+oM7KgQv88M4d+jZbDdoCA5NUSfITAlsxZZMFBGNxLyXRWayniuMTXAZI/5KB
yNmeJw/DxuR6WEVSNyJVRx0tCKxjuNA3Jm/+Ri2lwahOpqHNoKSYQbPrTUSgAYaJ
y0+LLCn634bSK7Y8CI/WsjdfyFxX746n2Q2iPQV5R536YDdJO/SlvxRJHY0+UY54
n1IeOPIRkxXPmsGF7MVrJkYlczMeydSczcnumLalvGcpcGG65KY56lzLuPi7V8Zj
H+okTDg7+UnCgaEV0JfIaGkm7ViTA2hZChfT4iTDllmvZ8xVwOaUitifxkr8TDSi
OcxKBsos9UHXiLRANSgoSsfU9+/o9xg+r+GSLItqNfu+W8z3t8qzP+l6vvkzJraU
E1C9WLC3cgJRTQKA6r3utjGGmQZtE/164p+VAlSFb6+w0xqXM1wyG32ArFnjDAL8
5putaSGHQy9/5vD5aCnLNSmjoTO+9nHz/XoIi6DWXY/XvOfU38eM4C+/rQU6VzL+
UQgVjX4fhlTlh0pkLxxcYKADXsZ2/0r4JLY26QK3DHanUMdIKak3bISj2XPmS6VM
AOsvPEZjWJ+vu/i5X91R0eRPytr/1pcZVe9Aa+7fFLxC8gm878TRcMnahQSkvKtF
pwa/In/MqcVGdwxeFbgATvC7msURn4vKqUaCClVGWOWYCBP3gIRgjRUfjLthwNex
71axPzyK2y569Gxuus7TKBNUhdy5jhpTUw+HOTid4MbnwPjlf2ZFba0IFu/ZpCMc
MSA12FHbhlNppg+YuCfjnnZQaT1qS5va79Jj9FK8xMv443jditeV+5K5zYTX5IYA
QCTMt4rdwo74ibIzUjQSrdanwBi1IAE7TZXdF8raLE9/KIt3YRqnloJFnAHIReGv
YYhv5BHRnTVi5MhvuwLzkEQVXzHaKlPRAmuPGRosFB+wmDry5ooCNMl5Atl9+2Ch
+A6FaGemwdPKea6lFsugPKHdeD6TJHHtHTs6LD1ftRB/2h/3nrTg3DSqqBDMYPfU
J0it533F5wdYId5wAYs5i4eZblmfYwohi7IhaPgz9x0Qt0F8Fk9fsHwFVIMw9oDG
xn6HlxU1J4VGBKeOmsq+/2SyjLJzpC9zbU5O+x/EbFNVuIGuTeUZmHxtOl3nOAZc
KsGi2QSUKSKPVTbvxkA7H0/9r1qy4O4C6GgVdZtdliRCvOx+YH9HDeTGTMGnjQZF
LrI8KYXgitc/o4Nk4SHRvUZB9878tkAQVs+StOZlT5OMMeC96OKVbg7L5OIiKLWA
8EEo1BNXvRr6bW2la+rwwSi2C175So4BKlSLg9D/oS5D9MUn7UcYs3g9Oiy3pGBp
qZrrmxkUS7fgltFjy+ttV3Gat4yqLDW4Z/REatmyC4BUzbYScmgnYqxc70ckT96l
1ovDBa+lkp4Dq+mM/nC2L5H8iwjJXy1Jyb1aO7bHLJRy2YJvYDs/hE/3NotUWu0n
zECWbmVwE37ltbWx0GqoPrtX+xwhoeVgsCYNFB/xZmR1pBXdS1HMRp6e/Tdr/fkC
6BivBpS6JLM/5xIlsALPaBb99qs1/dhIbqxSkLMR3R25GrKxDEhfZjJhtN8JxQms
olA9jWxPb97x9AwLkiapUUTDo7rj0hjOkMSewoA2WockmsiaSDeZrafWb4eU7YUR
eQreCdtcQHveGO7oD2Nd4XVZsrXNl4/YcO++F1QKfSbwvs7tVvvCpbF2Q9BTDHi5
/va5vJPGI653Xm23rmeKpr/MAo7U2fHbaWYSHmTR2kx1W9gICHiiit67GfP2UB08
HKbCDcfh5zTahKMt5DkIWutUlhSKDDOlH9hFqY+lqEaNFd15SUYAnLXxqtxFpuzH
wwInHk5EohjNpitclIRpeGK7UJubkDKTc2Em4f6RPF9Gg6oyrHEPjrj2MQITgEv3
ss0RjdQX+KwG6r/PdjM6H9he5v9WuVB4dpSKyZW1aPu5tCy/daJVbBkvpNVwRY8r
5AOp2z7AVxmW200YAtOnhUkBUqvo8xZ12vNG7sFGiaVHy/LVGOAPAHLnl+TF8PGR
85NQUjV7yXL5z8V2dNkEY7dDF5SOInCFI4kgm+rSnz7+yqGqfahD4wuGKKHgGYPC
luG3qqrIZxtaLmLH/jHyHuB9QDon+uX/r1zv20eea5ohKbjSTkvXZpdCmdVst4G4
kHFFI22ZAQAis3GrrpHxE3jJY5GXpw42pn0a2dcqYLXNMZ3NY61w54X2JeZh3OiW
jP8FV9PZobEJc2uh5i8vopcaCoBrmX0mtOyDa9jfPjznYeGHxYhUEwn7Dnktb1gM
cCM62ICHhNOugb73kQunRxikXm6GP4wb253+rr6QQ8CE+5a8eN1FYuBf+Mylg2hI
m5Ikoe32D5pcZnwbpG7/NzkV2ZxcOc8jFBRsTa/MMixcF4jKD5NTv6Vw8+mWijn7
sIceuLYE/yaUqTfOh4WhhCdyM7nNKQIudAW/ie0fe4k6KKzRn/yB/ljuFOj8OOYQ
BFLtnaPk9tckl1oEz+iEvDgDO1vInYcCXXIvsDujLUjgV91SGHcB+IZfUKZZMGpR
D5AQMRaz5Sd7vTR2w9XlHnjPgQuehsrFdXuBwTXj9E8Wa8RMiz0CbUCZY5uYfTFc
0gGjivr9e9HOy899oH8z1FfRgyqR8DYNp/lQ0feJHlnlqoztqOF5+ss9PHwog1nl
fU5nynKSTMbZfLNbbWrYXOE1uEWQweYChnILTFHhGlsyJ3X8SdoKwCFWdSGHW8g6
3tvSJdUr8L8gqCQ7PH6YnG/xe0qzdcz+y2I3jitErXe7zCCFrcGrq1AZii/LUQHm
qZkbCFmfswgT4ugHtAyFCXs206akmoUG+WBWCcI/dKvcDnCdilMhJ0yoHHVgoHBr
kfr5O4qSPjyJTNLVVrA18N/i2MkIb6B3zB8d4Mj3OesNMjn5S0KleEVFDnS9W+FU
XYjWyHHP1ES5Hhm6eLC1VdwDnnkyXfvxqboiPUiyHOlIMXhkMVoBCLnf49nB+tWP
twg1LRkFLkgptEALw8nEfTK7YzOtdEZf4VKAqxnEeKe2evwszqCF4chBOUOSIPKL
2rcfzFVuTaeyE52SzE1pFnJrSLxTpE+OSPzAIDmszEk9tCGnuMzF+l0K2sfWPegA
e6IT1hIWKvt25LZjldchbBhTKPTcCHJHZHX7Yii6dH7HwOPFaNM4/FCZ44gebCgV
SW6H+KMh3A4jzPHSctXsQhWzIEMEvI5tvBFwfjtoRD4wpjUzlY+9dC1tMoe2CSsO
JHlHXVDm4bcZ/KaxI4aryl9PKaaNbZKBrT9T6SKQXIB9LzJYZ+v3B6Fx9q+9V8HY
QBANXflGpZDHHJoySQ28yqGhXf0VSZ2ifeZiPfXy6ikFJA1jqbR2tNXNYzyo6/wg
rZ9RykAvqwo2X8m+2wVKAGvg25lVYlNFPwHSp4Mz4eY5kxTRmjyf490PRuiGE+g8
iQ51dk0p8R6RdiY7c5kpFE9g2X7XMzeFwZuqRx+if8DJr007QT1Jebr+nyUsLoHN
xhIzqRTdaaPPdXZ8Dmha8tsr8o/W4Z4SEAIe3jWS7kLg7OB24+YHfhPdvTC0lXIm
0rWPQKZhEoMbJ0sEj21NofNBktMx2rUtqTXE0eRquRfI7jGeLXvPlrfqyqoDssEp
peVGq7ixevXO9Ich7fyD57bOi78w6UGlBQ03MxhMRjv/eNuULeSuUqHo71zbFgh3
XMGtSOo6IaodV8IS9+LX7ETvuQmOqf0l57Uh1KUNjhoh85nDOu1dfS/R7pk3p1qD
LWjyfXgbzeJZKwBMQR9SeDh0lN/r3/ThwfW+xiDwZCpZqaDpJdaJ9/IXTzp68iqB
JowAKSE8kxPjbE8yfO9ttN5SITfwSGix0xNXfZOCi91WCZ78O4zMZvmCGI7FQdZb
7Ceq83Vjosf+rxOOBbztGu8j+UbboFvLQH0WjhjJKBkctH7t/Al0wXb6OHZ/D85Z
wNLNUsXYa+iIiuLdwxxqH3ZSfOQjoQLUiYwOcuRW8Am7fmR1r3TuATPcOPUox8dR
5y1+I2YIyIBvql1PmMZRbqzRtJliIf5cmBFngRyf0vQ0kEUWf0IvN7wXB5RCXUeT
SymSgRQ2Abw74QmwRzohr4V20xwAK6ww9whE0nuPbNBXFV1Gc8X0PshEfxgDmAjZ
dL3VH0Ur0iSJiaen0qgqJ4VU7xzksKz2KoxF3k/tMKNaH86ATnSet1EL0cK0Tk3t
4v7x9zQq54vnizFW7SwrAf25C3lvFTACEdPgjwAxRqx62z4yTSb/51DsMuw2cv7H
loDFRgc3oIMygMqJelPYDFuMvSnH0kQ+XIF/cN0ExlreP4nyjPD3mJTpDiYTcd6c
0Dqt1hVbOrZjQvpckUK2NmHeqJEuyI0r6SF3ezQo4f7Vp8MrH7dYkdbG8H0jisR5
xNEeIP18wG2cCvpEBGWte9GUWO2BZ9oUW4ISXfaQP1JyzMA4Ea1nUOmMUkGiutbu
NUHQsGXCYGf/OAlE/HaS/+wv/o7avt+SKsB4ZtC9DtXvNPlu8WfLHgZiGnurV+mT
Xh8LQ9s0bL9iH19we5mdd99w0fiXzEWmDN6vfsxQIVT4tBWbNhi3/eHm6Qk0tOsl
fCLm1jTLvlc4kI5zqsmDdXFlCeCuenMm1OzMVPw+ZqCqDdvr1e6uCiIUCupYzxfh
st+ubcVXkIeBSAa2o8DA7QqTsQCulNxWOy67sWjjb4jvpYJjJPN7qnltFlvaldfT
m0JeAlUn8k8I0z4Xrv+kpaFIzSO2S880/SZD24esge8A+uihVTca9RsS9o8w/J10
mKDs3i6VqGhKxo7p5G2Of37TBmvWX9uXD6QzaU7WqJZNqex7MrVnK4VesSg5oQzp
llEXkZgqsHD/49BI2MqQkdMymBjSGkZLSsqcJqqWzLpBJORp+VtMmEBUbIk0Dk0Q
N5WS46UpbobkPmlroTk81Bbc27f98zgQx70nAYEe5vrAPgIolS5XnuQgQ0zCq1pj
LkmUhaKtDz+i7R6FhOsSYBRucLbdXO7mRBYU2b1npaCutPyneAlX9bP7+fU2KfAd
qmSL1S/xYQnJR1CaKvVICFXeUmPIAfHCW1TqscxCM0KYKBA8dZRQdCT8mQInZ48/
CXiPFeMhmMy6wB1EawTVabkfKur/Ky+hvkUBfbr+JY6HpuqGNM4lu2DztV5ODujK
CAckkJeV1vujPBm2qxuHI64YUicjfT0k8YKWH1oIGMAjhBbyLZBSE7hUhIs7AHWq
bageuYmykIYGbas2BUPqeu/yBMx4hj3nh/1ldSKaddSqV1JJNWREmhO0inlQyWww
5rIQqzWF8gzis8ghlrU1xDmSTJ9g3aerBcatqWkwwfErZmZKr2C8TXixYVokxs/3
jY/ZWMvwVouzPCrkCs3ERKmz9plOYafc+yNfcyw+V2q+jhzdPamve0QCC004/pwJ
4hhfnsfTVVL+ayoBfDpVp3xPwd1QIfArJy06Frqz23+4wB0p5dpmMqHlS+T4Wv+7
E0mtQNFjcv2jS5LJyXt5XBhZPId2iapyIggIopEKSfpLwO/Z4ShBu75KJ/si9IIc
u3pCUcweiRdPKVdoCuI6mTAkJkWsTsH7Yl04XSUcDHZo7KBjgcz4N8HzxqJu9o0g
CEhB3J9ag3cqkaDb7soKg8X87qSsiq4gAptTZAJElzux8RmeHKRrEeuaibHo9Kn7
69ZcpnpSPyGXO6434nD6BQdZZaQSHdm73ZWBqFSne4duxHYWXtHZE5UbjxquA0mf
KmkIAQAg+V3/78E1zdlpPkiDAaanu3/tvtM3KPafD55lCCh5c6RNIHMiKp8X5SKO
SYakivwvKi/DVNeWCPpinUAs70bwf0WRL83YkWu0JSiSxeaGO9Tt6Bm0wisbVam4
mw9zRstpbdrSAnjV3XAbiKhywNOaflAWpLpnzgs2kmTdKbvLM9TnvP9X2W0v9NbB
2GowdxrASJXedC4y/VvQNCO5m3F8di+0iacBER2shlDUCHd1hVD2VuOPjHCuBeBE
C/nqHoU1y4IWikPT22+7ptPoLnBWJD3MTVdEkt1dXc04Jo/2jKFTVGDmgVWGFgA6
bC+bhWUqBiE+X09qMXytK561ws1USgrKC/LH/q8HN1oexVVwo0qYu3e4H1lpU3pz
v5fwFdKls0cS0/0xtL4ICCRsTN3mO7fF9RARxtHAeV4qQEAxk/zm4nSF6vAzgpXP
GWBK6MbINAxUVxNSeNLT5sWiZA/1tQK3Vc8SFPJ748CuCjUE2DyXlRVeidzGiB3B
06YWG9UveTMM8tIYdLr1B0Z1Z6Yx6tvhmLUacaImd+xQyoY7uPq3K2noxS3NhmyF
Yykp6sjcnj+xi/NflxOEd4bU61eWxcKRXtubaiP35Gbnapl1T+oCmjGlprmhFFeC
XGwshwW1TfaMrU07W0SWY+XBOO47BWcQVxIjm+OoUv36Q9/N3R5RhtAgLwovhrfR
FTogGGAjro8q2nF6AwBwMpW26nXJRx9YPk/8F91ZOKLJCS+HVoMQXUvbhZtwCoN7
GloTid08p8TdAuLgaIGbJRxjwEhe2akp87wXaKhoaxFrtFTSF2Q8RwoqTSGuyOhT
iTJ81K75iCUrLEMOJWU7ft05SpWm+bmWuOycyq5RVif1cYj1qaJAy8hiOE2usnvd
6CLQB0UL8lvd9g/CeLjZzRuRdsWZxCa+M1LTaf7Mni5Dc6j2ktVioyrm6zl71ryI
U27Otf7+oqT87sSDlhVVs9XI1TCccrs+n05MU5WpCva1Ii56N/7wX5T1RDhvMZkH
3WEThkSnxPQ/FoG3z1IHL4vhUL1OpQzXgoZz6BxCOpaZZkhvgM5jByeqPqRCCwgv
hvnJw4rMEtuXhKmQuBIfsr9LvpRSI9vlswDe26G5PcZgUy0Lk/uhtzvRnnHw5627
MoEiMKHF/6m91hbJ+sig3luZChV09VLCFGr6aAHb4zpjKSmlyI/Z48xKNGx5vu9y
as1G1OiTPzDJbozsuQf7iCvs1+dXyJs/3fF3FRjjHlcIXnqWowz8EwUOltqpv237
Pv29bIGb3i9OgYsLrld4UjBDXNEoo5AHUlHFx1Lip250gNJVXZ/aUdculsh4lCWZ
pTzwPXyOB+v7zsiksCgbAKDeuerR3BT6jyzjdUAZZVS9dA0r8L4+kYDcayP7IEW0
sFGXX/BY1d6xBT9d2tXHPWDsEsEBoRRgvcpdUgN5HCAuJxbWpC4ja0AgaNfWyZMx
ae8rxu+XvS36YolvJmbqNp+17QaKBpWF5kC5keWD89Oi9DxAgkzGyY+fmvkjN94D
LgbtHzzfKej+PbqQ+bDkaXvPQ1X+JRktUZwnF9iBde3z1VU1SQDo9CM3tq9GfqMe
LBMLFzwS05PqqGudEzlaSkFE8BzxyvQ6s2sk4E5gjNBRh9M1h2BQC2xcZ423oS8m
EdG5t+xjBk+D/YdoaHiuD6vCId7pAknKbwtsSgEqvJWYR7vtqNk1QH34YGoxBrj5
I5iob7zbh08zLVyNPhH7F28fVyK7dlFWS3eiBi6leQIy27u+0hGRdbuWLpAPGCQ3
OIlyK5ilHX60r6BVM0A2RpTzesjUVntfu6pDrOm+Irp+W332QExgzMCwSsuI4oZ4
4/04ZVdVQkaF93BUmRv0iPiLTfsXLYPcpx34ZCP5D4fskq780lCamjdlrBy7/RlO
P2/Yk8Curzj/s/NU7qAGazQ1gAo9ROfM352HBI282GDvPIbrt5NAqFSf+xIdNff1
mD8vTb/BPMu2OK0PvMsMfBWHeo7Bu7uY9xFhkzHCB7id3a8pXWHYmRiNMCM/BnsQ
p/NRtk9wCPicaRJgzmXsJEQc0LkTI7EoA+vrlQVwOiZWz13ONCzO1Gh1iKqeoBN/
626KtKQHPPimiJP72DnJZ8Gzn67hnWcOStlreaMlLpdUDlDu2IurZB8FrD4oT8Ah
f2j2E47Aqila3W5mtdTar4IAYIFOSN3wynwwg9fi528aFlQPkbHmJKbE6QjzTAgJ
ZXQxH8CvZ8+s1Q9MBgmYxZ8nfhnJMUGHwEqn7yalz9fX/zdjr1/OT0jg50/5YiZB
fzLD+EwKthcN0ofHNXrVhr1iuO5PtMknrxowMh7NHInRxvEw47PGsks7zk2bKiAq
yUPANlQ2V3V9n5U6lw++CZT0hsvr4tCjSmc7zNhpGaDkDvnbnezHTWqXccudLSQg
ZHjujDmNLnleMcqIUArBcII1gNCYxZuONCNKi6e35pDNm1O7wl0NXjfRoBPMXcQ3
snLHdw26NAjmntMmTIsiVUGR1t+m01qT916KbKInKERDyV1I0P6a25efytlM7s5t
sp5nS+d8lJ/Q4TaKE2Rt9P/q1WufJWcXz75x2lGRM+mBM10IeW6N5bQvzTfjr1aQ
4ySkVaEwj3/nYl5HUxl50PTnnf9QzNtZpCVbVwSFFMjkd2BXpCSixQsKkIW3xwI8
ZBrN+idjO/yFl6g2JcPurlGTBOgFsQ9BS09bvSlYpWDp48osJcXs7YUS9EvizAVt
rt/I3gKgstGIzdU4lIV/+++6mr9qU70iuFzwm1df21XLB1jMo2I5BMNLJclRwPMU
1qid7y9conWs4Pn+/KQ53dDqW5Ux0lvwXKNvtZFshjJQHSHYxhTzoVk5SI+8jysg
NhJ6LjAJq1G97teseyOnYawfP2+Y7/3TteJnKM+QZQKl7khJabcI0xhz2DOHa2wD
aCu9+kIwVJiCqmVgfY9cUcEQBBPiF9B3LfkbuIUJmaeO3LjpNUNWjwGoJ8kqx8rD
HByHBsI+t0LfwqQPoXcRaqjtf5S2jGDb20wtfRU/qVyepXHao617HmBtBW/z0NJC
c4iRKV+wrujV347QjxdxiJYNIAu/XuFHRRFg665sLA0Yc1asjiiry/nUczrL5Q3Y
Y5Nqs9gQEFx+jgM5gK7scY+mRHNfSSD29+rKT5wUptoeDJJTtQBlDemht9ClKzAo
Z+8bt0qaWZCi3Xvv0jKUMNY0h2OZPmhMYvnRR4AvOgR5z3gKOuS0KFti5aH2wQLb
KLXoFCJMM5gSvPtFtyqQ4dvsMkCYh43T02XN6FaKBVBKA/Pgeov+3dtxWGaJ2IKu
cJ1PP0KdIf+RS5yjjBp27+o6KDfQYsrOYePvpiGAMQ3/vC8N2kjnLV22v2Apmasn
KETz98o7zkJ+B8dgmnJWA0K4Db3W26BxYUNeBmRdrRG2CYeAaz1Z1P6HaGpm3xFh
fDwfa8KK/LqFVCHUu4yiyt6a066YUrxN7L5qQgskZtAP+CJHT4EKgdakVSzEd4g0
caO4VaApZ8c7YOvJKpV9xPOEQT8ep0Wdk/NS/s/KbXIr2fAL9jPiO1hn971RQRbX
PQSKlTNo4o83rY0bh4JhrpVRgml0FX4rAk9GR+hUGl4zf7bLx0GuazYvEWrQ0hi6
1lspPXT0O3g/p7Z/zhW8yIhrorICRI8BrsEFPrqn73p5on6KgF2XyH6T2e/W3fmu
kItRuMHGJO84Y+GOjI0ZiZsEXiXSdtbeksOMUpl6Nh50iggsighjrQEi8YlAcN4O
qp9Wzp8UhfswixrVCFXpd8dDFeqrGt1QjyDtrKe6Q8xqgXAaa35MjvRXnl8WdlMy
i+ePNS4WXeJrKoWuI8z4OnN5Krk4F0QbNkNEa5WcqSaBdLqZZmwwmmss9FSWDf0v
YqJi46tKH2hEOa6AYxI/Fw6QQDKLYxRYB0jX0/HKvJFJTktrkrcMJbsN7/z8TUN5
AxSPLdaf8J2Y17LRxcG0HaS4NpfOchGKsqQ1XgMthUyoKSV3/19YUAr/cM73Bd1c
SMVgsA5PhV549Ahb260c36YWMWMoj8CXJ58DR0I0isFUh3gSDiVBF9cL10jAKpYG
0iNIrKsVewaf23fTN2ML7DEzKya+Wzz/AiijAG/vbZGLygd1HkAgf6I40gHvIkHE
wKOlBtpbVybrjtE6F6d9//pCYgK4BB5iPrCPJjlLocKIQ65mk5FaSMTsqdouutp9
FiaQmJK/1XUDY/mxt3EU+IDRv2gBS2v8p3XkxgDpX4sWdQMK+ZErExXNuf9WVfZG
+Dgc2awQNAQ6Z+hAn9y4q3WWIO1KiaDHSFTdpIh0H6qLfgECUgSwRpCIL5SuLE7U
6tgei8bb09/Wqoehv1OzpA0qnHUt9qT4iEPDvGgFfgXbzzS/iQsmXx1L+e/ikz99
qDTgY7uj2wVJetXq5/h5yYElhb/KyDZq+hsc9ycnYbmMIBqf6yTo5daZbL6E/aDV
MicaDYAZ/PtiWxaba1csQW7Ezv+KL4K/4iRepzuLj6yAFbgatd3N7yJuC/0Si6AN
j6vWYk+K9GLOv1hF5TZQkwLfN8h4M6GPw+MCeTHWCiiAaJvCmstOnQKpcV9wQT+u
M41AKutP0a4IYdktC6xsmRWF7g5PCqdBpbngysm+iPdEdTTBIqj2jQvfZZjXWJvU
6+IzoHVlwHLN5Cjg/eSfEezUeXHAGcnQ+nWUMaHMpRvx6F/AL0EnBJoSYqiGZZBC
42NpeUf4rP3GY73NkNj+J1cesP6MNif5Bv84LCOgVzIDUMagPMZntYloubpIoGEY
p7KcP+201f0RLsokRVWGUDO21RdsykkHgvIckz3uUFo8Rvz7emHZl7q8WjF7ppgq
tRBYTO6fKoGXrZe/1HaA2fbA4GkO+8hfLvINh4YNWaOqDn53dDWSd6omI+xwASsl
FsxlEljs0Hq7RK0W4TaKIUXsH2B1lUQXrE4YYhNA+SvHE1lL3VEROGDLHNDCbKGX
VWkJE1tob7dCXseQbpc/lAMbVfzMZCnIyYghNsKxChf7gQGe5G2UpnkCCEClqbjf
Yq8yZA016aOj28sLIhgZSdUrG4lq2ZSboeRBqIRx6ZdsA1kKTXKuIHi/kweV5wbl
X6gVGa6rZye7cn9qW5zJ68WWs9Us91z+sl4MwK7p4PjY2uXaI24ufS+GTJPxciSg
g1MuDeP+nFjlvX23zVM5McEO/yFkQsMXd0OaIWY9h6P10ym1SUPRyZXmKA/bbgAw
Ik8B5d+lWNIplXvA7eY1LM3WbGCig97SC+KqDN9zOIZl6ijkSRH/kTNCV9YauhB9
jbJ31xPJICfl+hMDl3fv7mTe4/vhQwyt8GaeS4es7UTCSQQl/m3ELzMQl/QGX0fi
bgANMS5Ecg23gU23AZldPzgFeJkDRtvXbkzsB9Dj2XZQtqaHXuTvEJ4aylioeusr
5CHCB96e+QOv+ChsJ0t4phFDkkcfS1N2hvr9atiUmtFRNClR5spG0jcfw9wbLxzL
e39XcBpgjxpvgwEuVhNVEt/GQUoPwuD70umPrhr5St+mJcm0wro9cZajejnRwVW7
naOuoVo3BiRQnPfVnFgNQ2Y5qVfh2gM8RLJ8e4tTjxKO67XLF/URG2mDVnl1htJV
llziK5/nQTzrTjylY4z3XF4+PiWuOFlU7+Vu54fq22QaYpOSzaphzikCkZDrd9li
ZxYpo8faW5l0lDYj3pqFuMlT211hm80WZ8YH7yMhTW+Z0lTsBE0w1plreQo3e5Bi
Om8aM9GRfX6Cyq0ZCOIgangcgKVNqhpnYHfYiUz/Y8ZksvM+dUaPLH27QtcnuoZ3
MGtKvtuRTTFjLg30thbzC9S3IU3q5QENDvCzvtQGIy060tCfzAYgVXHZyDqh7jUH
g/GWJVxqmhTJahQfWHCJYcrYC4tZVkbSxFWZyq/6mcMKXvV+HwN06MsqVIi9U61A
e3Wn64B1vX/NGr9FIc01yVnO9XRHHO/WAfTFFLb8camdqFf7hOB669lrFgwwVb4B
7QdgpkKcTXXFTD0GGMFmzFyAWoyNvsRZxMpXlSjMET1jChoBpizkhd7Jw2R+aEL9
tT5rdqycJCVa6Ys1QmsIkIDID5ZT8plOmDoRqAT5nmY6O/nmbcEBP5I/ot+nlS/0
mPSW00If2Qis6Mbd5O4Y4tgYL0MmPWRm3GiHiPXT3fa1Pt5XCg/tmBPTAd09ZKK0
Hwvws1m4bcGjzgqlQvKzAUv3OdfjjcoBVQyO6HmdQAfKdrGDC5OZTmzjOMXEEr1d
6bUMBgbRUatUDYfh032iGIfbt8nEdGTw/0XF1XBEspaFiPSdGPe2+j/Ns7nH4iAd
RnVmqM9ODBnCK6MAV2JKxFfM7Y3DBsBPOMiSBEthZLc1n1OokGeBJzFTqw06ZCes
+XADEEY5eHiFFgNo/tFiwlYjVQDdb825Pf8/3Mt/l3cxHX6+7Bjl+6k9Tw9uUX3s
mGbs4u4RSIGC3KAhHu57Ew0AUQIraWJUM+oU2YEBPZQvSoxtk4R4Kx6czCBRt+cy
Tv0ISq/Q4N715aCKmwZc6yv7HJSK4qn8mRiwmDhjNkLeo8kr2aDeYrWQOiINWaK0
ds/xZHNQ3+9TP28Q8VQu0PEw3p5/MdjzaEa3jR+6us6QQdRiWFOyMKQwTJKjBszX
jspqgIpFNiB6Ra8w9kDQzag52j059doRQ0N7QRLGWHiQ2SZr/++dyVfuDNj+LYfN
WmS64mOwX71y4fNKW5UFFQ0Q5ji9/fLFGEopWs5k4PsLAdW+lsl0uwM0HpY8broo
8Jg35DggQn6I4zF3jWEVYcnz5U9NAYpBE8beb3WK+GjuScY+VyeniuCbwU/iFcrp
lcxUm946J93os8YqF9ZaRzbXT2RnxppH/YJSo2EXeRYoLybnLJ1AIuClr53+jfOj
rh6M3Yv9orXu1mFn5llE4f/mMlFNn6nh9M9cwX6yTXbnlSb7/wnD/OozEn+14YwH
tBwtMsVeWHy25ThuBFWkP1uM31b7SaLtg+cxpNAQ+enNu4bPqJWOQij+Oxyow3be
tbKp6Q/KM3QgPiKTESwWXnsu3GAGM03hBvnwDZrOh+y6jn/ihx7dfLyJjVtpYLCM
VsCQ5LV1BhVFZrQP63tUtmcvD7nsEBf7YCPAMgGSxEgJQCebebwA4H6oG2SCE1mj
hwlqPCov0CJcXYTlnOqfHpZuwMRjHBq31xT5MyDSPriPw60yrQ+7VLZc8dRDrr5C
WPz3/jQeiUvmxSv+/EZFYCoQ9opzuE2qYUr0js3wmpAFRReMUot4eG8xge1I5xip
Q4J9S4D7CuVminBVIvT7rYL5qxO1x5Cbp0di76TCoDoliOgeDJprOE8bmlCuLHaF
zzxSAnh46bnjMrPGzZyIQ7J8Cg1skWktD9wAQBmTEZifu2r1vzbSpCnwrI1O1qjr
+8JFk/cXbD1LfgoIBewqFRcFnlgBxtdcRv9Ym1yKJ9k0NAmmJW3SsYAIBWWAHbtB
d+19ykZtFjhy5XJA1IFiOOz0wjJU97gH93qJ6PmAH/isOb0XF1j+Db4WATVRZe7R
sMbdpdw1FZl+3QmrFK3oaPpDVMywLUHIt6LfUVGSBkK/x9HY5UUZNZ6QJUfueKxv
1H9BPubnocJ+l1CBGSbcco7lr6E7MmQuK0EatL9nKjBdbXJ/SZbXGke3g7T7tL2H
5XNns7qGeMmaaWlpxWJIuEXcYdGg713zyZC/TPfn2Y+pwyyWz+W+j6MIYp6VNJeR
2qngvGiImk+OPiVYPYigQamLU4GNvApTKoE784IGuMbaHRyzBxuOVIMIVq9/ZqOt
N7A6Jxc4JVlHyyDAfhE+iA7MPHqaU9Z4mzRbkV+8eNS0GGQ4BS1Co2ifUGKR/uXd
UahrFq/wtYp6g3SPyg2Fu5U/MyhFYEX2H5PQQX7NCCD1JDmSYT0SYOQJ8zUmxgBr
emJsQ7FVnw2Ui9aFUmpeumXRPNfYmPGu0ciSipPqA6DPSoUd3l/GSbO34/Y7sgwF
S1azL7/vS58loTh/IvZQP6H/SFTfIn9Q1sksKgS0GPGflQcVhXhudcjlSTc+1sP8
xDIpP/KeykSrCOToPVqSnZvcsng8UWWA7G3S02MaIq5IE2ej2xzejSaZ6sl5dTL1
wGSnpJgU2++Ko0/KWfVWXH8wel03nzhwjORmgasc8JhJVyiGAvhWEqMXlsMljsUm
X4rblMKmjqL7URs8ETo0r65u2tPQ7LPNVvwV7wg8DC+uUAYvuUK22fdUghYAUdEE
B5/bzcG89JLsCkGRy9zOkMs5NiRvoqloXO/gCLmprcG0wuLwyoH6eQ7JDqisnYWo
pOnE5SCOPCq9JWddCW8b6Pe7IQAfn2qTSdyKgDg1mCwYD6IJLJsDSkHZILzzrr1h
6He1fXyKAxkzO0B5Fl6dMKZA/nLmrS/MYCk/d4j4IP/+kr66mLb6FTbtG0fZpc0X
LlDh8YcqaTA7PqF3+pHyjV7yfToRvKIHOEV/8UGCDHriNLNQ+v1AZHKLSYb04HsO
UEYET2K0pcm8+0gMa37JtlOJXVpXpAFLV43FOdmlVbfFeZf+WgHbJh+rQ5ZExNWs
6rExGw5Ppu30IYo/No8opeey5ViwJ8tYj6Zp+512tTIfFLie2O2bztfquTAnyAgM
gx2kUod8c0MnWutYAXm9R3A+Q18fzkzWybQlkrPA/625RA+ILvrH56aZwQ+AVOGs
vsBaz95WTj61f7qyVmiHgDE+tphw/e8g8U+/uDoAZYalf1YkFUm7G2gGgkC/w46u
upU6LFdwtd796jly7HDlttmBW+t1g1E1Ab3AKjT0Onftsmkx87RUg68A9mAO7Gva
CwTBp7z+av6eUMuBMNv5jCnxgcDBPEFxrnQ9BRXDTlHYeJ+z9k2kFnuNR9VJbdRv
j8is/T4c4OGgDS++xS5ecCo8bixFbuzM+0433LJFsO+X6Q28dgYxwHInGH3gCF4d
E1wiDgRy3G067KFMRAX/jlBEKd/G/bIO/StnhDBJw6Dv3/MycO+cUN5xFe0ZD6o/
sJo+yv42z6Pq/kz/xFJOU1ugaaiChwH7OyZHPqcGyMRk7Hs/hoKn8O8OuN/xa72T
bTsk+lKLQnbUl2U4O7u2//36aPfzV7O5qyUbPziAqG1KLlYrrVxia1mXKUwS/RpJ
bCSalubwjcL0hDx018ZAz08dlQc2Yl4wI95Q9Fs3ZkkWSNGLyGHDkkc4ViKGeFhq
zhss/9n/cZxznSNg9XDq2cbmO7uNF0JNeW7totm79cDTov545DvJ6em1jdwEiltZ
kHLvoVs8nh0SRyXlP18q2kd5g3t8WQBGZMSARjwzNA3Xr5D8idaLC43j4GVb/KZD
uYPLOd4xmJUAK6sUOHxJn0yyabqJpsgsVg69z2d/uJSjeo90lBVdGPNeDPwsSpLh
hYl85oLfT/htoRjPVfM3+8VYt9Vs9Y1qBC1gfh6Jp1HI57g/ELChwTfLzb/kwIlS
XDRrzz7jkW7GX4H+1LtoovAHl0JeFahzhA8wZmDZreTzqB+e8DPHpvbslm7MjPj5
mvbqtGAKXqH7BBV47uVvYLLqoPrByXIb2poQbrF/97IBgDzAmKgAVFRvzYfmFNLz
J0gQDipsJOfpjObROp4AEcM21TU6KUS25OtbRHJqprm5Nebn0bS9PFbwSDnDHTdu
7ZFPDxaEhWbY6heZuo9fFn/DXIOXCUMugIGEk+pcAFwak0wMtMDEH9eYUhrrVfrY
8kZLxCZfH03MgtGnxFbildBf+SVcA/LnmMbIRX6oqhsegTWKAenaDipnyAJfHlCx
6PevmzVtj63w11HlyrNBBIz/HowziVTobBJQCkWjmyv+FNpFwmp+0bEfSPGJKZTk
+6s2KPfHpeTUd73P1/xNcyVTnVnTajpk1l+JRFpLTiECFZ9WRh6sqbjE9oKRC52g
Ip0lBRpFL81B1Sn4cQMAEGepNKitLbwAE5h5zgWBeeyevSn5DrLVOEmK1aEKE2Tr
3ULuC0euDgYtVJc4WDS7L8vJEigaC1FbPa1vLWgNCYny3q+tKI0eRt2DFWe0g60/
GLsqYKBIC8D1pItsYdcPpJocqGv+mwqVRI4R/ZM5MiAFU/ZzImmqfrLjBiCmCSPQ
irlNLCd2vB41a9yOeP09gtT7RQPSCqXgQowx2CvmcgiYsxtJkSfEp+3fG8QlN21/
TD4//9K8B7X0A0dB28x5QG9G635ko8mX4MurKiKNZLJtQKH2Sb1DgPsTDvZivBav
wrPJ+A5FrPeekMFOafzaxFYVii0bnby5XgQ/rX9hxvMv7AaoCj2aR+mxK018usjS
o9c8az3QPcMlZrP4vLxt4WSvk4GBM3O3785GIGgIZjw52Rha3YCMsv7XItGuJJ2h
YPwQH882cttxcdB0ZIYvOYJc8oVjIkORorP0Vw5dcAvzrv1SsUpaz+IMI99scdoJ
e5ajqKt2yKRVJ3Ywi+wNXz4qmzFHpeUB0P/6ZOEuO0Hpo4XcgqeK88s09LWVCfDq
F3qFeXAjuRGpjwsedSqq3hOMnXVXxBAWui8lz3XF0Cr6MeBOUkeYNioM5T50akf6
kTanxnHuA82KmxP9kLplK3p6RMBVGjQM2sM08wXBdiwpXKQ8j5JTP/oFWu3bI3Fj
F97mv9V7l5gSUKeObNAHrKYgfu5D9jVKg9i9OOSZb8htEr2YSQJHElfKgaJp+sQu
KgNdeDGmkvfSwqrKEdqEB/Hmn5aPO7IX+aO48H/xVp6+xEhrYjWW3Jo9zQVVyhqN
5szhyk+TqchF404xnh6JvWS7YsMD+oQ0VkyKX+o6j6P/zcd1G9zZ+uWyzOnacMUq
LDPZ6MqE70q1o6oZ4IAoYyQtIrVT5y9uY0+Xahb1jKMVNdPd3xmY7fh0yNNZ0pYA
4COpthw7gDqIkYVbK3nNpIjQlSru9WLG6t/mlyiJdjVZKLNcEbP5Ac5GLWNI9QC4
3Yi5uIoJbo9VQF3WMsC6k6SXFzTnY6SE7PD/vo11c+WXFEJhxJ4+qwVmblVDBFl0
wc71PfE7YI6YIV7qbAYvotUogYNijQ4vOhY3ey8383qB5OmagCucJB0wvuCq8OCg
lJujjjU6IN7f1Ho6m0C9a18r+q0SS13EzLuKivThGwFk9uBopFnRlMAImYnf4PWc
hv2k7WFDmfy7WNBpIe7seEpgjK0Hc7aL/iybttA2D05l740rhwgHN+JNPvQwXK+k
Rcpfw4mxQwN03mHZHury2Avdb/s81r2NJEz6am0xk8/ucOQQ71Iyi9IapwkPsErF
fALMmBNNj3xUl8My9rcSq8p6L6TbJ7iJp97QpThelr6g2y33kW4sIXDd7Wd7a+cX
NHYhQmV8HPF8TEEyuQDG3OkwLeW5dJwu1i1DjsMU2ChVcsalBiM5RQGFJYvK/f22
itbSV0ft1EtZwrXxusyEs2DG/wjmD/kuX8188cvAWKG7AbnkFBPTEuei+GlQP2IW
MEhsORt28jN4Gor9c7bmprT1dJTeYep6KlgW/DVv10/fNqnAMNz8EJ6dj4PD7lMQ
6Nh8AHmeHa5cEhqclHxzqtLaxrEet2eBMNUB6JLhId5xtgXV7CEBHWsiOckKstJh
uqA0By5NwtGRWbECUDcv8gXXFxLARcUKaWIaK2wv0t/fePoqacZeWqfwp4ZqoI6U
FgCgH3RdfFmhIhISeSueSKF3ups1DO6FQQO2Dpmdg2h8b91VIKJzOIDqfLHP7A57
KMRWUvHDVsY5ApQw8fbeuwVZecXjlT1e2NHlCCo+zEwraeyzjco6dI5N2GKudiVf
ythKzYuOP9jV1aeoWv4Xyr7pDUOVIGW+Pba5O8tDDlJYVR5H10dkm1zFuaHIw5ff
yGqdnDg1O+4cw2XtiG8b31s8evjzTR4mb5Gn3QIXl0GhWMKHQndzEdcN8iV8rO+Y
N/6e2+9WdnUB1+L4MV2TcKaUwEq81kcg3/GFGlT60FLkxeRG+rJjQhvpJbyAYEce
Ra5XYYcb5ivSw794TcqVl7SB+glIqk34PAaq4POar2icnm69+3NaM/bDEtqihBVS
RGWDnv3/NGo/L9XeOz4+LnlwAtp3pIkSl78jxkBAYsoZpzXsUpN1JFAkxoCSDS70
fhR/3IpoyJc6XBtE20S23nRKOBMORE93AfEkKKhlCgL5HzTPk45OqqVL01ePgkjQ
qDBnwQChlwU/8imXXY+tbiR79f0YRAs5+xc+GT6VxIsx8FcHhDacidlTpNKVVpot
IqfTcaWFVKtwSO4gKu/yO6y7mrkh4RkWJT0L8cJHFtXhwt/qt/VfDc4kWgUMJ9A6
yLh4bHgAF40w5oUNYnBVQNUr7RF+dE8CWy+d3qjwF56PP0CsoiUeLoyqW3ZdJa7C
HCk6QQmSgbnEnFKpjTMHGzS8/aVbPIRV2q6T8b8UCGD7+QQUnuApl2wQqwJJZyYH
seaHFMnB04nKOIDwfm8axuv9oBukKK/MZijUaAERY5Yfa79f91riC9vFSckjiVKT
5cIDRWmUYbANs3WRbKyvaGaEGrNt9JAM692DmzCUobtDlGXeNMB60yCVvO+a2MwR
LlSb1Th0fpDlfgLXZZrnybzoFA3apf1hWIlIIqXtN6tiUk4UcRivRzgh+9M//9DG
gBXyvwPsTASPMdd3q0mkIJPq4xD99g07UphR9PyONnuwgVeaADxL3tX2stZE/wv+
tgJPRP4nbjtElsRdByFLCePYZ2aFwpIweqHyC7qDx54NKJ3CAeUCceEbn9BvXAIr
7PQOR2NxZY+w/lIMhx57OQvNlgIotF6U6RJd68Punb01Dm9RKXZxZqmDJ4eO8m1h
EoH5uwLwpMDh/k5uxYhqXViqjYgzYsWBgWDNcW+ra0NM/0nHntTQxXR3vEztaaws
csEoZ1gUgMdytdhC3m0WtczSSMeWNH6ylqMSthlR6Yq75w+NQRvjgl6piUTNcGor
kDs3rEfObVSTRVtTk/bStzg/YVzxW7SnwzjmjZGRHO+wI/VG8enOICDSn+cq/8Ys
dzawDjgeWG1/6sjfyykJS211TjevjJtbK4TBfbItAbQ97QOHs85Q88jb8qgYXcVW
/jf/9oGAlyRFGI3mXxwvoxF0DiyjgxnBXgg6sZU5kj3UnTS5PnBCB84EKcOkaLmE
4NZI03GZarE+h7MFiUwE6hj8lfxwW/tJuo+/OHv+tAErU8kmuL5Ec4ZGU44Z9PBf
+IHMDG8BNsZTBdTVOZpLbhi5KdgHL5QlaojZ0nnDRj5cYN2WVLjmAzOG1Tx30qqa
eer+mCc3OH5FJ+B0gjDa0AMaVHGCV/C2KD7zys8UIdGMZWxQL0/ygkCJoqQnktvO
T/ebyR/i+yVduiYHuq7WldRRzplUMQhl6QvK/c2Umu0M/W9Y6fQAIdnFK/dFCxRo
93TZr36RfAJ3qFJJFX5pABYfOQaqM5YbqdATTsKRc+mGRMpbJ/fisQNGMW3pnN05
frSg1EDAPXutsWdE7kTSQ480LFRqYzeqPFUmyc7IXI22AAS/6v64yi68pnCEBJiU
mSr9sAswhZ4Rt4eSGF04HV5omgFj7GZqlmHaxIF8DznyXCOM2PtErnUJ/33P+AV9
GXCJ+DFhFbvnCL3rfkdymdwgu/8M+81pfOnucLz12D7qvVFFHFNsp6JQLIc4PTEL
ymrHOjZ3oDTHIIV7MOmG1Byr3BDqcPFKKN00jALjaU7OONYUyxJhXW/AQbvrkPgG
CQOR4bkS3c2ticsCiPBUDwF06duOy38bvu8JYO6XOYy/YWrBHghvPthR/JD99B6t
1uA6tdSpzyKCjrKuhp9Qkm8YCV/xmDsWXrRc1IKgYq9GgacDJ6Kvkmk0Hj2J19Y4
JkUnObb+5PfmARC9PUNEDrC8yntIxIR3Ul1ZzKZGzpsdGJj55Xltfl7L0Ande8rC
6EKe3XSB0PnA+ovHjmNu/c8zyBsmqVL9O7ZchZ6l2TQlG2e/QkqiF/WekGFZK5Nm
OfAqBSqK4INd+udtbKzMkkhoRwZaXTDRkZfapko2KoqKzUNN0TYzHyzxHQyPTeCT
PmRcUAngq5RXT89qGzeA9OFYEjFNLXsmekvNU8NcuSRB968U5QV4Z+cuhqk5xMNj
RcQWkIXtd7VF8Jk1yGvO3EqkgH0A84DDMlAnkWVbtLr8wXSQHGKdzFB993aCsB10
ElNH8k72MouAAsvPVHDQxAyKCa3DSIuvniMd+nMd5bbqWWT36Z3Yk8DbYDz0F4lL
ztJpm6YyLG4yjDqzLHkaOcBErUtdkTed6pdLfJF9L4jfSISqC79D9kWToVj//sul
3eM4VXZ594OXYRNEwibLt99uAlDA84p5X4N2VEPQvg945cQSk9ZmjOOBovb2xbej
m5TV36403opwH7688txIq8ygkI4vcfLQvp1YApgX0k/I/jzsQdBbICqTNvHEN5cB
cH0v/h1NMPyYMtzvfpG+uo2G2WnyIUgFtwih1uabjMfwR1rXkKqMsq+WzfUI66AN
Fw7hpY8jnDFe5YUzRqsF1hg83qo5UU0N79iCqS1sq4VR4IPRfssaMWyZarkmsIJs
OH259SjIz983xeIYaI5/lSXA/KfQv8vUC1N5+7quVUx9P3XFBfnfmwRDhFQwrtKR
FYJxlOSr83CeLdm7bZLENsxZLgeiPiisLXII9VZG2Kh6rOrnfzg2lTZKUZhkq8Dn
oj0uCDyzg1SK56ycHHYbcwLQxjjLXvZvvDTzraWAT7y7I9hMJX8caoLpPIAhsw1O
+mR9OiavGQM3bq4g/3EQbsl/+w4SbK7hx4xmKLtRz50yH42fJz9b9rC72h9n3JRh
SyQqFHHCHAyzr1gC3SEypEb3hyj6+q+HMRzj2iQw63pYCK4MGnTqIhiDV1vNqnaF
u2OGs2Ogzc/7dej/m1GRWrTnZgGrQcM5brerYmVVw5Jvsyohg1KrMQg3rJklZH0b
HNLKXNeFf7igIt5j8dJevmTXrPCKgpi987cVXwJQDFrVq178jXDXKTZFdaJ/AC1U
J7JD+0DCiK5BNn9RvTbcEDc3KwKi6E54BWDVpKpITaTmNCccmZadwl0lLFswXPoJ
saB/gy07PjHJ26RYegkbINadxbGlM2rltcA5qWNhNtvyu0Aray+xiwmFWSTxn8Xy
zT437sKaQTHswMpUC/64oZWoyEhHBcQtQaZjFtP4P5PtvlZzYIy19g6I2HPTmF03
CqL1RJj7Z31wpFqjQ6D9QvvmmkyefO3wd/42myU70/jQV/7lMCGabQuaC5su++yP
CEUW642m1R3j25VRTUZ5KL3+VOAnpjgw4O04qDgXC1o+kgQuQ3/Ts6Sj67eCpPW/
7r3oM2vdrju+IQRNI+wppCVmUnzpFB66FtTrDbxkleSysO+mRrjFv5vXLFG7rRQf
Q1594QzXTczCo7DoF03JElP/Utl+nrLCyJSktFpVuiZKOAzSuMDMRWwA+WFqoqWL
3L2LjU13iLdcQRx17ZoBhXSe2FWkeo+UCJiVX36SdC9RKc3AJfY272u+MF/fccLy
fkguhDmnBwtpATRQ9xK5/Ha4a0t33kuBBJrEFuYwIKDVHbYXUa14pToPP5duLv9k
YjoLc+Y7WpJLwt2G4tYtI5kYDSpQuHknuXvQIKEX/CXfmrWND/tHFbgIh7TfK7Sz
XeTQVTUVgeS77yxOTh10FXfCl81pG/Bqvczx1UWjfWCqKFPuOytxXq9hvnotCqgs
JbHg3z5awrQ8tpgU3y4vnZuu7G59uSHzFKldBH6UD59MmD0lSaAqU/n7LpkXaYcm
taTDAswCbscBqW3iAX6F+BpU5yaiVuB1OgPp2qWphmqzEqPyWRw7EzltYLZAjrSx
AkXm7Z8eBMGLtQuy2wOS/BIvv4PeJJAnq48s4e+swmEmueIz9enKA5Mg1ZaOmCuN
Nu6pvKjZEhsJn8fhf18MnNYKP3r2xgzDAVcp9UuoBPj5cFz/FUZPj2L2w0DU8751
dNTSSx1obPit34pZNBnTIWjEKZwUVeAuP6kMUtMGquK0NyCUsmp9BL0vQaQCois1
YQfI6cZs6NKEbW5fTB5ltvUNQYsbOeGBiBFaRntj3JiqJRx2wQEZIA54XsoeItb6
Sf/+uiHHjeYKKtvNm+vO7i4c6grEIk9APkcpOxvDJeU1IIjWQKNjCrV1LoRDRVIN
dkkKbNwc1hzrcqj+DT8RJAGjwg1JA4BFLN3+LmFZ96+V/2g5Rd8Jvh5Ora2bRX6T
sinJTiMr+ZYRTB3+bUyWgUEbTtIcQriyfK2GGCdwquoLm7xmrCKBAr0jVHsPB0An
+NC86Lq3CfLD0yGq8A+SfaghfISY4t9mrJ2vMjBn3tvfwUA3QyKSS+4tdH6jKz4B
ahwD/+mWWjk0MSCoAElZJjjJ9o/PnudCLBXQhS88t4MZuiaRYQxuHlEb6QDcDvEt
nXOqtYlouNGhd4Ur7M8zx6PUyN4tNivxqmpSWbP7f6E/jF84EWOpKhzcK1X+3rzw
mu0LEuhryFbT70dE/bxjog8ke96oyl6ovZKKcP6Nzz2YsIZzUuK31sv7AiRHdEnN
4FAotZY9QOVaNBOLjqMLGUZbWBrTCRDAxbKbsO/DkCAwymgQ9pm0VuOz43QVWP4S
D62v94pYovofZx4+JKDDMn9z8g7rgz7frzA3F8QbwCLpV6roQBAiSPa6f5pRo+TN
yyBDQbmUk+ECoRjYZiCOCyYyNpS2csUoyOTTVe/3EsBsu40ibCEXzreuDyitHyTP
vU4htbqGn/SYj2jIuTYMLQ8lZYIxKD0t4T2Mns4ivWiRUKBl+UyOHw9ZwlSt/Yhx
uMkYUz6IbWqQUqOjCQ3D1F/O/t3iWdiQp7O7Y6Vez+g5JNX2sVeqzWcBqN38bI5f
83hFBQL5nxIC1/VWTNWbAJ6kgzzJDPP6EljbAtPAleU7BjEM9kc1GAVutymqNUh1
zzMx5xaHV1RJyMO9+tJudpQO15Vmlk93ZtWLLi1aaVoS9wHkO3UU+/H9HjQxZNY3
sM6Wdw6gNaW7emOBre1Yv8CcCjezAzMRbKtybIiZ3NiWWNfTwsdPux60s1367m4n
GiSalp42NTJ3JIf8K5/HZ19KSDeeV//3MnLm6usftGrh4UpqedZeCvZhi2h3ERST
3KrlGXFwoBIRPCFX9PS5XFJmV8LaY+dTgA9DC7Udf7VUZSJdvXhj7oTy9LW3smbE
8COeyw8SDgdHX1EnLTEWWiVhPxejNCGVOWqziPU23WOgsCWO9GCrOvk3qb0BYj5s
SHeXOcwkTlWyjDU5lxItWeWyv7Qsa3cMQYNT0+SYI6HvCMBWqdlFEmHakGwIbRqt
T/vlFxibrpL1xUM6Plx4mvJa1h+JCe7a/ct55FkRBHhXjiBaFzFG3S86VTHp7ne0
7dREaT0aHUu5pu4U1c9KGCGXe5/rfaX+Us4i/mPAMU8Ba84sjgRiTCoFejoADa/8
pi7rGuXqaGAlz9ykpxUrsE2201EzDmrdZcTkNVYDXn7NXYdyRLmiMwjyOB6VJQWC
vC26JhAXuaZAVAUr2uH9sReGNeZh28n8m/6ZwqmRnRAJESnvij4FgkOBhAi6ufi5
sKVKpVCxY6QeSlk6IOLXb8aAHuMfkW+JqVkfZFr9TcH1mJYMrU5P9Dn6QjGndIWD
u957Y7fAPyjC7GQTj4IpJmqmDh4gFqfeAR93oeAIBBudTHq09Jh+qcRnT0iXfoHB
XXtbPTLGBOK8g+1UUV5OXppPYqQm5PONgl9NgrHE/AxOV2IydCPd2As3WCEx3mJZ
YiflCTrhbjEEwnZbLaVijdFTvrz907yYYYqs0R8po15iiGrERp85b107LUjjMa9E
VYPM8oUXpjfHMDkbP9GzNLSH2hxNXS6Jo4U8fNSfPyAS1C18iGc8z+q70MnoeDpO
riJD94HGphvjS/Rm2TZ5upSIO3xnAfwEtbxEodnZoTlr16PBVyCdc1cSOZxyotrG
nPYwhY8w8Ww1TLiyHwjvZ7UUdEsyKiufDuO0UCFzkD12CcfSoYqLLrugpA5pBN7N
nZ5k/WhPFv6fmt1t/Mq1xrrcqRyHCMUVIglbFbliWHtCviNf6zQf7jVmx/Df3ZhG
DrHqBq5IA2uaetMwxPYWm5irfrIiScif8FewYnxrzym3qI6koypGH0JQwW1cs760
ac0XOnS667qRmegtomGIAISVUI2Sjjm5pE28kqrhJPQak+2PwBwdbnH2rdIS2c2R
wVxVR/zUi1+RDb1nPjJRoADxaNTQGK1C8Zfm1CCrWaq4lESzTqCVz62gA90bfBo3
hMyARc/8ulit6gTTXPCD70jZ+CndqiPUELiiaF8+pS25iLpuSt7enPEPFIj8ODnm
qjBWwxWATWBYU36DKshdRkcsQbNPYvgiq9tAyDdFH2W5T7ejI3t+nc4av1qi3RE3
ih4p9toW3qidgO4st382V7I/ewpP5kxCVCdAi0KGoyjIeDVe5bq8h6gLHF7E9I2v
qjULRmOynRJETC59FOBwhrxccE7/LrBgh9xFxBt9RoJM2+BTMPWYGGxftK/5Ncst
CJlxSFOyrHMP825JbfSwKHYUmMOoMWZCQudEpJEUZZwib9C7QGZRG/YTdKdB5cTS
UQ6I3E/B+S8s4ZxYhaFuBIAdJ2E/0KYBHYkuyr2ex0LLT3Vm+yH85jmXu1xe1/zA
/hieGZmdKrmaeh7NNKgEuadhLKCy3/jtGQMdMKozW5fzqR7SjC4iNiXvUA0DMs+9
w0OML0mTVHu+flLN437z9SvLUFRCiDdjJSG3cnNOYU/yMX4MZX4Pef4zd8GTDvoi
48E0oTCWYIiq3SH//XJeO3tp08Oj6PpQLT2ghlRNjckWwsdYFMGtTGdtKu6V2nEp
isX6TTUgVRfh/eKpuku4NWxlltuTLODQNyh/weNhGEfE97dWqy+coIbDQcBrM3kD
9LXvIBhKK812jRnfjSWMZpX0/1+ASTwTO6hK3TUqHrpaX7NW8iQJn7LGIN2S9+0y
rKoMy9R7w6QS/fFRye3CAS/yq+YG7ajl3rYyQMHuGtkI8d9Grq7wVgg3YRThLSTk
f89wHmELXv6xXFiz/4oVkTeF/2iCDQ4BX0AK0l5c5BgaeFLzq/A1GyBcatgPgTZp
27rser5BuDGixf4N6kmkVYC5EHXFbB/Fr5ydIOo3+XqMgtCs+Y7ePQyig22W2C7H
ewI/7zE68k+GkHXxP2En8TdNgTYB/6eFJm0RLR1f6Po/b7UHcMKLUxSPG/rkPrmK
xovOEj5Wa3mWJQl5qidOvVkkOYOD8XEUrNLzVjdlvKhIKM+PmEPrR1Vwz6XIIfeX
PDGFlKeu5QVKS9pOzDJ8ON6vQSbxi/UZ4uQ1YDZiaRLiF44kKxvvsodFqNz0Jx8d
8duxExylyDSz/mEFjmMPxxp7ax0ertwqlZFPlVAxHteLVYh9SHv8Va/vWZmFquj8
QkZQKg1hNFSoJDT/yrAb/IDSP+3wbfJ9izug5iqcPC3ypnMgTk9XPc5FgNOjFjk1
1djlPGL7VsjJuTOjRpByTqvfP0N92u73ErutKnRdnlovwQOb1qrXMkICjX6fkvTq
yN+n5qKPv5HRchKpoTqmyit/deKDgSvb/6LNSCbnn2xOK1VUdU/n5cF8L+nfdxv4
9/+k6WpKmijfpUWtfoqt62YgaHMT9PIhK+TcCigMhOiwVE6Lri0tn0vdoDPMYSKY
iK39XbAcreTzLnzDXpBSKiFlQqmhfUJe9QRBrZdAD8dmsQTGMoZ4/QqoD1h4A6ph
e+I0u8ptZ9irg8MKbHybmc2Bro6w22bpIPmp7XGDFpvF9+Q2H3okBr2sbzc6Jxdv
eYbEOQYeVCwYu2baPQcYZ6jHbw/8JtQLJXjloUWjm+VLdY19w3UmnyOqgcEaF8sk
Ei45rNESVv/bfe96NkMNHcEhKwX6FjCA9X/ev7qGQVLEzG5vQqYOKGtm2TRs4bGN
O/qOc012qWa4+gsm51g2d/Pch2t8c/XzBeCB7rRh38uWn7AIBeHgW6CG5q8dYhgo
RxLyaUVrwgPGLLr5NeBbUpndwrdzW6Ii/rh+nWBhuVTYGu/0vVUzXpcjU+ibwDbz
5dmHPYTvovN+eWI0o0P2cGb7hj2NQhkKZkJshQR68uEje60iKD5DG38cB1JshHNh
WG/aCUO/N+BW0gyIV5lmsxvQfAKHllYNSsslmQm4xki6UBip0Q2Avz0ZQFMV8PhF
jrlP+Qh7bNwzyM8tAwKfUmPcTHde3kFagzs6KozTcnDD7mmajywIc0Hxs/27Iw6a
ccBt/Onv/LMosbQ1CV79tfZFmIp6digCFYgmgFrPexZZJxNUm1cDJCU1hMbFdm0v
6DTQr8ekmI9B6p7TLxUpVavgxn+ExcYtNzHcP6pkfJ0gCdXCBc7AiXuStOu4TiH9
KX7wJG9rNJRIWT2VWthz5/1l/JjKo/IWxNzENf/j3+fRMc5UwD7/SMQ/XGBOMkxt
qZ0jYdBX8OVlXrS+VK0onDzNtWd74haNdzHxZ2ZceKTdOfn89qWMPKyU8sURk9Um
MHdW7Pyh+sb2woP69GA3PIe9eiguQijwVCMctFwo71QER62tLj5cAz7sk0u8irqt
5yLrXHz8z8Eu5acPB9ziqBAejyLk8I6c3N3oOfGsugYOEaNi8JW3k3OalKgtzcWI
zLIlF/QMNi2lZsdWA+D/CA787gtjiGCp3n8/9M16XBIxPYiTPcsV3UjOxIwa6X4b
pZu2igV0ldtytGluj6yjsQWZhy/h0CEACK6yAZxkHBMtNnbivqCXh/ptbNFKtS8a
5/mTKzAx4iOkrsqt+KNzZnZEsytvrAr2AWDnyGIrNJLQKw+oP3jtGtzpwBHhHVHa
etgNSInMJfN1zparG6N4uKNAwQ2Of1cs6xkxzS+8NJMu1qYR3h12NundxNX2tv2O
D/4V7knS3G7MYF14gv4+ekQ49RK2271LIDCmhfN/nASwOvd3aKvqbgtEDcXU46dq
ro3IGVXh1B9B9fjFZDejdzrKm+lhvE6p2J8DeSv6r98nrQiZDWF+Jy27J5Z1HGbP
dvXgilbGg2YkWdExXVyHms3bJT5hPDeFz6hv4j8Y9Wsr8cdEhhbSx9Y68485ZvUu
tPNQ+G+JSXmjhYSaWrzEjjPJDOpBL5T3vh+W2BkQrNMTc5I8B0nTLNd4M//alcmA
yHYh4j0XdnDjRK8kYWuwn05UbKdU2mJl+bUzcR62lOnZNXGjtfLXVmDMtUAV2WEe
YmjuvBph1PZKUtLcqVDrIUtv9UKfwOGBfKzum0wCCdpzY1uzEr+IO7lnNAQRxSiB
zf+wStUyw4K+j5RvVAV9PMepK6a58JDs3QfVh7xb1NvF4wwH+2lAOZ0E9MBRKUxv
tJvP6tYJaxUnwQcb6PHRC2J0kCz/3gfFt7i0s36gOIhA5eui5svMzn/4o9hD7/+9
82K49n8nZDlsH4g0pJ9j1srH4c+Z4cvlxx3fF3tWwMiidyrC5zXWnKLhuUO6D9ur
oCe6FsrqHbDvmZy6NPxdgkl7gFD5NqsdsqPlb+igdX24zyhMv6a1h8AAz0V17Yl9
GRMq+j9/erYeX+zD0npjLJwAaTZvjrLhbOARssVSLO/LNuCRDLEhJwZ4FpLczLeS
mT5xBMryH2N08etGpKsCaptCTFwt4GYZ1qQ+5xKgVyvWJOuQuWns4XVVDrOWlDpY
K8D6/Vtzk3GuoxUpGXnOUb1K82GlgvQUPfXItPqPY25lERASi/9Bf0bQmyxIg0af
yOMxdE9oYPpKnIKXJSlNG5e0Hy6e91E93JV0az25odH5n/t4WyahdsSp7VDJtdOB
AEkJeJjyH0X57z2Gck+iB9RsSJXDOfwvmk+Cb3pjupXoeKsNi419fLtfzAM1C7k8
i7dRmoDTcXrV6diUCLsX8FvV7AbELUILx1liUnIZ30E5yJVcffNhi3y56r0XRZbO
c4wpnkFuLJBecngUfyDj/fcGwqWFjgeJawI7DsAxJgz7ZusNy04e22QvZfXqPh3e
6UCOH5i7ZJm6rsBvoWM4ez10Ia5Gy1T3app1L+V+Y7u9CnGpZv9D7pMPoT9GVZIs
zY2RDMFze0BCF1AA0oBbEtC/fXehbHgrd3rlBCHD3Ht9KdJZDJRnJWmRTPJncI2z
Y3QbcBek5BidFJvNgQpPldstdj7NMpfNFKQYi3Oel9JyTNFVVvzV2LtDs0uPyBjO
RoKb/IDUrRHXKcgIaRKLjqie8M1KKoteA2q5Tf77Ws4FX+HiFB5dyRf2L8eit13V
kvpL7/wO1Rzl0v8uEEjX1XgV0wI2bh1xps9AiiGL7bG+7q4PJpLK4dL37RlgNG6X
+GCMaVfNjsLTJbqp2TBG8Ascl0/vGlyHvj7Our7H0xW3H3edUw4+oRsczpbmEF4u
WpzwZ5D/0Gck2vYt3UpoRQSTzSn3EGNfWZPE0yGi+2oL8/mHJPjb5ggoWL7HS20G
dTSax30b7t9GLPaosfdKCaRoGT5Yz0CrFWy+5+hLC3GYU6vdp/LG/uaOOM3+LaSG
cT+HX201XDqcLWRLHQlD5rXHkwh2JEV8q8/xksvh4iYY/Qt0486hufMpCJHsRy2W
DlrRtHqx9k4piggMuFEP+usOFqKYwasxMJVP/H1fqipUIzDboFlqgTPXGk+wNPhd
oekEZ27E0kSTSu+ptAx/+HWF2+lbB5cX5V7ezJHKl+bJ6S7pm9Q+cxPnxOyoliq/
lxcoNthM/G2esmNdPovl4YJ3OZVgjjJlsclOzsXq2Fs+BCvahBFiQDDpnH1nMpT8
Zh44RPcYQ2m6dSo0VjIfpGoPIOxBnuH3DEx0IH5gSmV8fR27VlR/vULVQqaUTyiw
WMVNp3ACRdaGXQDZY+BYK26Qa9WukzInCaPae0l6LVtlvpzqFrFzP/yQ9zzXX4nl
7QLPKd7P5Js5bFG6LaNhx90gsNIRJ84/KS6rCZz++Sh0a53k2v5+CHVfPy194Dra
X2VNLNB+dqsPiBOfMfX5rHr+viD6xTZhUb49GdsbfXNig/jSzGZPEDkAhKkAKEEH
e4rHjLInvrKFyoYuWsVCTEuU/RH84e6oljtryPMxzC1XDBU11CSErej0cp7GfdW8
TCMPrXq7wWZoBxKJBMkh1WnD5SZnyT+bW+DeXHGSwgPgMamvdJtFbIeqRiJw9uEo
1ziiMd0IQ2Em5Cm2/vKy4Di8nCTFfGNOkAv6Mtdl30zEfysrsxCNxrshzboUaHSQ
n3vEVVum7dykhcDx1CXF2yzk53s5S4XRB0cTpmvSMZe/8c3fxGQbNhehoqC7kQMX
BifFGdRg0YixQ3zf/MjKzwZchO+/kai+9tsm75ZbdA295Wdqro2P+r8SHlcH4lka
ZQCrBJoh42wn6nZQA0OGZwo3CuFL6GCfGEWqI1+vE0dFd0zRWrariN4xCZ230DJs
s8lcDwKLIAyJKxRsxrd3mn+I6geU7zqjZagia8GOPdGaeoMiB3OEkHzAWdzEUl2C
2K1zUde6WHflc9/wmkgTRmC7yjueO62NTwxCEQuiJQKqfShhacePElnIV8qwrXC5
kLK4iftGA2bmFsNcU2xuwqUEW9HVMmdYeObIqg1e+6tFAo4AGJDiUayL1jUnPQQ5
CP4lE3qz04T6omZFH8t8VDLLqeAiudEfVaNxmHPBs2RYELesdwZsPXEOvRic9JmB
Yh6ONwjZljLLjHiVWALr7k6xFs+ZrUPxck9g6AvoGjkILgF3vEfEdtE1f6ZEQNWq
fyOS7xCOuW+C0Uyu8pK5stDA9gBYJwCcD1HUps56nqyU+QRYymxdQxVdUxx3bh8D
MP2c8zRxQBGmYFMksf7qBFygYnZmgFJ0jXicZSEl4qMqWDt5yBB5uyoL0mjL9nio
VyPZJDdYs9xyQmbQ7c/aaXIESDx2BVi2r9Ra8tgkiC6+phz3FiI/pSIKMueYWLvg
XFHT4MoIGnRR5euQ/A376P3m7toGermH4JZcV7aRJF5f94FOhGI6GaLZcIy7JpHc
soqXtj7oPfmzxNrEkxwTX2QINwoLhqr5P943X+Mbbnii6drqWf9pnm2iVq6XQkA7
nVqI5sqqch8bMew+wNIb57Z0mnedZYFASWKf8HnWUadA9QIk+dmp2HY0G3awGAbY
Q7nFjhFsXUucnp7VNYjDWNcvXIBtHK72pfq3RW3yWbjQJ3zHfZjAgLR+7fg9/Gv8
QMxLa2bQ6LorzIfU20QadI15ET2gT78QUcz91gDC3ZJZaPPM1dp8dX6FPDwJ7xM8
GZyqymoJdpMR7R4saU8grKYzQOQofWbECkJb7dn784GZN0B1NFWSVgA7oLLjMqDJ
8Yv+sDnffgFJvukx4hsoZr6RJInopqx2bJx9xhQsLTfCeh9F9V0eoXWUKLH62vbM
hfv74o22FK5Voy5tiGUCBUxQOkVMLOIpdYZCfPYuiq38Kvu8YbhiR54oE2mBB86v
+xjZfxV9lWTFta3YPhJQ+eEsb57QI7R/GYK2GyWHZshZREBt/smHGcMA6gjSubdT
t0bk/k6NlcBr6IN2e0OVrzUFBZgmZ08ZAlzsCi+wpjcVqzM8upQSfhaieHJZrTQY
Hv66Q/xB3rdSuY9dl3P9BkFML6Dcl/p2ZMInueKCAsngtYTmhFZUDTCsx3WTi+eL
VqUBqOiRU5P5O7BofhJzpD6OKF+Pekk10LEUHLLSUkLc+wTAKqVrWubNsSEPAluM
zy1pKkUVloGXJxn4nOuJNE7uv+PQeScVd5HW8PLt0QLZh75OCO2zdzCU1zTCKcAx
T5WO0kDvQvQS0dfpb/+j527CS5lgImLyHrGhBwBt8gP+HF3up8EjLnR5PQ2En3/q
BZjPsALq9aQXq2XNaDfsRVPoOuYez3DcvlF8im1cYs2MfbUi42mPjvioTsRws31w
a+CFSf38eO61e6AtdUlUjl7/MSpVZ3xFQC+i2pxJgzS7RQV/S+RMks1ONM9xdz+f
mV7Sds5cYLoxcZDXSE5Uvk6/7I8ONki648/Umv9ayjJl5GcXHR5aaBItRH4Fdsb+
FIDQkP7QNY09sRZUsvZR7cgZNwN4z9a7MAI50eCd/38ZhjIbKMmMyvtqXB9CMr7G
MmNvXJNYgJQ359MwaCkF95/cmMJ4hS29BOvN1hk5Wz03GBScPE0UWaITxzCS+LKl
ySOPJVimXpvdP7sGzuG98/oON02JlclTvHusyBgoaw1dFNCknvIUP7f2xEPZyxeg
VnEMJ2kOK6jbQnEXCRr3C0SIKuqqrH8zSJHGrz/j0zDI7Dr6S0iqJ/FbTWBIsBBk
KE8jGBy7ezFFLUSZQHcoZLQtQtyUCiy/sJbsQLK0GUqrMMbDp23TkKC+fgTtXkx2
91iztB3nsXuuq3M8v8cf9n7fxSKGGuSmQE14VhuEINIO7I5y1G378U0+12E+DKKx
4gQ8Gj3SHrlJJJo+AUaCwgL/R3Tdf2/fG+Jkucl/m38H3Kr8Ohjby6YQYosV5GIb
05Zh6oZZkIGVLz15yL0+hUD95xoUZXiD9joDrEKuW7vpFOj3+utzWMWvpnePsKMA
ESuSylrSCa+VX7Otmu+zre6dTTrSTw2U6pnK7Tg4aPlYy2OrRm2Sy6Ecz63LsRdj
xKzPKQUGbf2XXqEL1zvWFhHBxGpIbqjcsFa5o4rhop0WLdwJPbqqGkcL6e6LnIa9
7r/RXW3GAt4EOEMPabo7exzkTEyFHf6kjkARR6m+dovatGZ80gspwCP15w4zLWWt
u7ecDH58Ucb3+Bv4iEACZBBxUWSlOFdnp7q3OW17gPYfJ2VddRCuDRRq101TAPXK
hR238qF3sCSRELWLdCOIQltw+fTMPL8+BLVjh1oX3gz7E/J8eSMk+rYRMxAHR/Vk
hIG2IcLA3MMHS6k1eQ5aYg89Kgr+W36s0U1tC4NTFUsbZYFT/SFvezkfIYZ5xinH
IIGmrPqkJ/DE/MF6kO7DjunaMPy6od1dcMzN1cu9ceYCDQJ4l4b1lSj4J8jmGapF
0JbJ7zVIT9SqbTw1Hjy+P07ulhVYY7ou8MCtcQZ+hU2weDOcJA02QGBqpXxz0PqZ
JRgINp3Xjnq5BkthGYH66lGo21xOGwAc5zNWqkqktCt8fX78Jvp7GhPt7yfnSiCU
wo56W7aZm4DAb9X6dwxPuQDDuP03l2q1EFkTeTcVkR4+pGELvLtHMDb8NA12k04D
pINzUK+RcmHa1oHp7qCahMDFCXPiJQkbmc530tzEKspVdz9KqOyEQh6wMfZjNZTL
/FWY6a5J+v8zBIoNuU4sOB3APzNum7KBNt9qwklgg7dFtecV4pk7SVBXPFP3T25h
QqyaIELd/HjvCzWUnn+mEa2jCL2y146nX1R5nrOL6/oJ8jqllfAsEoLuCatI5Q4n
korNbCeesq7xa4lc/py6Pk/4BmxGQvlw5Og5OPMzCj33tLpX7/lukPj/XVXCJv6f
Ur+G54+R/25qYs2sJv+c4UYGrysecVvEqkql1rIYb1Pbue6J26DSD35tYx5qyyDJ
kXne7DrNXz2RU8DBaKKcRasabH049ap3TEaydj+PVTssSwf8fq92cAN1OQXmeabx
OHifC3SFtziKkigwdw8Cqxui6W8LO2JWOiwqO6YwS7Pbw23BhTu2GaOPENOrwedQ
QKASeQ07oRgV7K4mQ6AZUhRb8CTckIoRIGGtxNDUjmmXPulIPbj49nOAH+/+3Co9
GSPE5oaIHSeQAlQ2dcwcK73a1biyQ6UUGe2Sf0t1K2rVWhX2GDPOeHLXBrpRo36v
5rKMJaZlSaWn7q5V13D0tVe5IEFp5pP/XvDpIwP7W+npjH+dN51hLaQbH1V5EE0i
jMiB48zy/OExmy3dDFDU0D4NVm66EkFT8p00ikaCOtDUyyGNdULkrrfnMCG7nOzz
da4F29JLT1RjzIF8nwkxPccPnj90W022HVY3a2ZnPelqtjCCHjKiBiivm0mBySfo
mOrN6GLfHKKn++pift0YbkPviqclWTVZtEQ58Gd0EYf2nQyFneqHMPThXvKj8hgH
FtVbdqBTWBH96zKiwjBjtrtOZ6xODEZlUvLJEE1wXqauyGERFg8HBDewhQ9cnnx+
Hvjqt5rPuHjtarGF7Tu0wVdZ6q5vDIHJUdSGEaJkDAdshcbuZkBTQN4a97bFTT9M
KXHxqkKtawBv/TatPZZuFyhzE4RUrpvi/CA/X8LGDiXEx7CLKALJp6VWLWGN+NZN
oOnLngwOegny0oVE25UsH1JLTSFdgU6qKAZfyi/wwsxApEJDVvOBNyDY8HkuA0I2
3v90xjA93kQCqFpJWE8c1CNvLi4DPeqwgPefRvmdy3Mz5E2NJq5ZIj4yKFnHirvR
KPZKI9skama6FZcrVnhK1mEPQiX+TCacL+QNyvi6trbTNOBkpmzfkFhtTmZaM2n3
GE9KUGrXwoeAWrckzsB8hbaj793pxBTUD/FBnS8SBQmZ0SOqiFBaWlDaSXWoyQZh
S6VIqBF0qi+vM+GakQaOhKQ8qB2f2EYxCMvnISWmBWdBbR2AckwiAK0FZQGQ376W
y6hYVdj2b6klKE4/H8ASyh89EGbbxrrIMNZ1VN1lk7yeUglHR+yZcw9y2lU0WLq+
PjqmnMQV9VqI0QnGktLV0vStS3Q4j1ZwMTpvsVDUtMWmjoTxdO08FKiOYyeg/J/V
P6I0YeVat7WwPE42mAUTqcA1NaqImXKBJknw+ETkz6yHuPZFdivIzMRjIyFfeFfR
aXJH86bKWS1dRhhpqEVGOINQ+9isHyrJXuxDtQLWIrzuC/i5OcMA0ujLezX8mvkJ
3XKbxhpb3Pzt88as4oSB23WU5LadnhQxVLJYmZVAOOoWqgYD3e77ca24aAVzaj1y
FpfMzAI7zccb0qo2/hx6TN9QoMd24UL1NnF3wPDQUH9B8+fk4Q5xw2nod9FKPFB2
YO5cBxjjso//A1wYRM0PRkwe4IoybNHZgaqDURELI40=
`protect END_PROTECTED
