`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6XjT/IszlOOOBl8PzaCcZMCOTBZeiYKKImZDwLMxSkcqFItSPAD+LfB3zETcJMET
cXjtM1qUyksfTWfrXCK6LT6ZVbz5bKG8YtKwIjZ4cfZbAiUfuu9ioo8a0zgE7fOE
O+6K4PVVaFWs8YrnoLjE/NN3fwwM/b7ffJE1emLZnb0srIiVJ7tfws/TVWIdtkWk
XpK45MKD+tWyCgPXjhFl1NCQqkBrlKZafR/Dlur3XrXT+24hS/JXlDuS9Hp6QlOo
YKtZIplw+BWezO+pcE/NFnOmdbiaeFbccpiKrRCCn7hyf0JEzPELOxkitoo3LLEM
LQqTbZvnHUb0jcU/ipCr2O9YGjdGiBRwqUfzYOenxaQCIR09aPcmGDYeb+rS/CKL
C8t6CuQrpoWAqqAicWiiqexVPfMziT4RO7dr+YdwgAw=
`protect END_PROTECTED
