`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7I9f9CClXsFejU/LVInIuVyPISMFxFMvYOFimZ7pKl3adQ+edGKLhLxGH6N1NLsO
HtvU5CSU2iLUDbPSGQ+7pl3buz/q2W58qX+LKnn6TXbgGG0HqHdmuuO8KNJGD6+h
ONJ7vMSSnZ5SoH7jekb9wnR+GB3UQqiaohwCjasPTsqZQnpUA8XzZkQFlK8LDApz
QtmoODhBI5yKmG3zVHFcsQmNdKO75y+NkIM8S8qb9OwLarrcFiIMSNDYudSPjemP
vUrdrUPKOJC7z8FVWT8PQgCdjzdsDR6gmz/wXwcUEIp2z53XevSQlKuR87PqwyFx
SwxfL2Pbk6efIZE5rihdZvHjrM3DWiNSoWGDFAQV5v+TFZ+Aty7UyTdM6/04gtKU
NzRam/VSyoMgl3er0BYiFnMYEgBpcb/qVfoofi8Pa3HOhGJdJYdQmT268IJHdpSM
E6sgAeQRvdpCIo9a4hQsZkw5lBuAGhoKUieAIuINdvMgfyv6GMOfCaNjUvJs5SIP
fitu5yTfYjJ6YydJlg7AxX2twW5MhA3u2OlkZo5Y0i/TBgFEo1gyOM/FrNUT8hXn
pZZe8Piext0fkhtyPtsL2udQMLgKKKmR9Vf0BkISckviZ/7l5Z0qft2qnVIlFRab
I1NBILo9ap37vWsmtzCddY4P3LzSy1ch966JR8fs3AblBXcNvpaFovdwiQioHMiM
+IihWwSHVCWg8NEVq9We6jJ7y3GaSxeJD7Jns5LSL0Rxb87KL//c1hKRyZw4OCK2
F35oocwtzzDgZRkthLUdLa2oamH80KgtTDlDEKuMkf14IoDiPKOeN8z2B4z/foyd
NcGoLgGBYO9lBiRPaNF3Ye6/2WTaIvxcu93KzAIgKce+egjw/MhiT/bT2a1L0Eg4
DcX+/CbiLM0kJtKQe26Syf+PWDwBDZe196BV1nThr+mcNdoIY2/NHaWGZZ77o2qX
HBHJGx75fN5iHL2gKUB5Y1t1bIO+JivK1stQRM+fZB0O66sQzEQMw20nOsXjs11a
Y60V1TvU3mHIqVfypcyEAq2Ig/nvCGuz69NB12X258DcjibxGMmg5Zadv9At6nDi
IK1QVHN2nGeUE49pjQ0HpyN54HrY+iQnFWlwpYkCTuyhxl/ECADmXv6I0fiVKJ0m
pwULNUhkmOJusA6A/wWieLtidxUxf5PaxuZ43QlMvymolRKrVqVKzeomRjAxYviN
Amnc0QYlWYXalAXuMTqJSAdkXrMnBwYcjF2eJBDiqnXAR6l7w3ElxUzkk/sw1cJA
/mTo8xYXXyNUPXqNQecX92NzyiwBN6BhjYXO+Cqj2dITIpGyl52k4/p9Y6wMGStI
pCcewDheMAT/n5kjHT4ByrrkF/RvBSje+qKlmOPKDu2x5HRsCeNifv851hyOuRft
7S83g2NzZuH60QWZ7hEBh/lQ6MaZsQgEvFYkSF7ilpCvNcsGi75kJ3S3aBaevmzS
ReQU4sK6L2VHWdlfiVwf0PEhvN3+CuBLnGoeqxv+SV/zxykmh3LC5lHfeFGgsH3i
lEA1qeW0cNwrLQZdvmfxWLFeeK16FL2TmIuo/+bv3H3LX/3D1I6kgtIjjf7s8zTJ
l4zIQGVDftVfB0dd7FHJ6bfDUpBvvGJn1fFRK6wSWA9IoXZn3lCBlBa23InSaDtW
UcI67kvbz95eseTEGNIPzw==
`protect END_PROTECTED
