`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bSsodP+xACSM5arcyx0aZKKS+h0TzHnuONyGjrkRmZfJ93LFEpIz5B+HD3FmSgkJ
GjwI62tRHnHtbDx+umBzBA5XGTUtbMKD9UJcCKz16+i90zOv9F7yZBzPFCsSRLZY
pRbMO1RBu4EkVyeWXeJz5+AFqLYGONQFwCL9N0ydAi+apn2Q9eo/neV+wLzR1y3F
65bzPaP0p7AaYnEy2frxsjB/M9AR5Ed3fawIN+oMQywKJKhlTgMhSH+arhTLFSab
5Qbu5zw1Dbl+itnje20yTZCRU5AY1fZ4Ea0DI0zm1pTfrm8DjTUanvXcUbzvfPhD
EEc2khNX1aoBPuidkNeIrhKUIONkh2LfuOXIyoE6dE9fWoQ/nlJeQRLOx+cf7YVX
qKgpLilf7J1B1v6Hf688pbuoieZVn0dgEprEnKH25D74+OZkNzDTmsTnNf7sgHWE
5MnGNB3ibRLVpawTEQvVPBVZraavio90gelmsPfU+SUXqtGfRKd8p2PLZq82maqo
PgyiG6KxzlLRDDi7BgjlbmcJB8qR7rE9I+Zza4CdAxuOvaaCQ76jqisaeJ4Pdd60
FAec8wAj71Rgab+IdRTaMpsaDpvhmKQzK3YcWVLZ9VGaJr9cHCVDtGV7iS3fsFa7
oQAyAuKUqXxWO3sDOO9lDg==
`protect END_PROTECTED
