`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QDYg1XMVnWc8UDujiCDHnlSRgVtCL6y7iJwANLrS5CcYYAevgRqW7KX/GW0CDp2
8dEXjwDczIFGCM87Vmkk39Sn+u6SfZmn1lV+JaOYwqbU5JRex4bODZ3XsxLOilvH
4rD5mfhCU4uilU31NIwSwsQ7UDlz0UzFz5ZzaQl0RsUZyR9kHtcFUaHNF0X2Y6HO
T9KBH5EB1ilbKSSnHvxF3ao6hquzCffHO+Tc1FhJlx0yFBF8wTKF2vZYHf4bcjDG
RJrTQB2QT5f0W2553nuKjJrCL20ew9HQ+UrUxKt6cO9EECh3H3j8fhaHQDM9QY0I
z2TMSyddnWbX1XnVZSz5YzlWFg3zQg5VBp+YkwBUTVUyDodKbe8tiVO+/4g+mwFP
LGsvLQcSZ4NFWyGpkfc9/xFN7bTYR9x0H8tiD+3S+6cg0q8S9eQ/vYg1ytvIttkq
OmI19G0hVcZMEsVpFbW4r5TFOABi+jwVB2gVhd+Ew7bWh/FftGgAkc3/5ud16NAR
mCBesNpABftlr5xy/AcE9MKWQv5BonObxuWlA3NYaRF64t4ZVPslvsrTcjyOG+hn
0c5C/B3cJ5WIKhPKWpi6UjBvl9VTjPQsHe0xqB57UeqiMTz0yjA0tHf2gnKg1Do/
CjDgx0+BdmejUym+Z0HsltElIejJLvWQKPiGvw0M1y2TazkC75/f5Mq3UNk8eXAT
BU3q8uf30p6U237rVHAydwyN7Ij/YpF7zlKMQjWAAbE0NExZWKNbWaMSl3Y7SKfE
`protect END_PROTECTED
