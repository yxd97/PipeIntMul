`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nh99wCi9VPTbCfjmCemJkbgiyk9v0MPNUJjlkr49UbQa0z3fYh6D+23IL70lnGBL
BQaLxvvyTeyu87m1kzC0y0C88IprI27HHOat87mmP3gKOdy3WwtdBsaIqGHxBwHc
r/qC3UDISdPFFKld0krcEyFbhGbOtSzv+SCC24t0dP+0e4VtBRYCJNKqtUcDHogB
6EoZ6nTafXRfQbG5NHNV4ouwTWVxnjh6uXg4D6Js3KYIt2OC31S6tVQE0S4MsYfd
3HcB8IKYNeQnyrTPL1szrbPdSuf5glz9U5bRZcnXXaVoL4Ugd6TT9duL2VWKSIdN
UrnPduQvpQBdu1mpVzsg8Y6hwOs6UdCj5eQzqhrlCRaZfKaLE6GKSztz4i4Uzvim
uEbsSriZXQ1/YMrD7LDaog==
`protect END_PROTECTED
