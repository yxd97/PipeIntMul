`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rkIPUUsspJecri5IRCkx8nERWSoT4XKNm2bvkOcSVnQaMS/6BB99MaSL4Fvn6KLA
5HWQzctVj2/ioCYv+s10vvfZ4Ph7Tqx5nIb5dO+PFTqJiTDRmM+C+5OWCOR4z+/x
pJaxk3vORXtHlIDHQcfw1z17PtniBgY70tLcjrAiFpMNevmeM/Rry5yrEPUIN22T
88FJ5fbnjywCGY06gOEgBuUkVi/f0naadkp9K3x+4WJYnGGHAWmdwaH2DkvVF1iK
s50YEuAxkBM0yLqFDmv63wY68HLs7MorkX0+uolyPa2oQRG5TJCv4ICWf9SraUhA
QNd+XLS33xue92notN4AXZ36MWtwTWr+dyLEtHwTux9jPL0DQHzjRLZ6amiJb9kW
vfYjO8kHUXSY6VWvvvDT7ho+ket6VjWYkH29m7Mx9BL63emFty1vUm/D0t07xxJo
EM41G2qCAlhiU3cbRGjqMDgC8CicWCv6hUfVdt5KIs8D9ID1xm7hhdqS1iWLWMsS
PwNtQPFzuOgxVbhhw7/kW+N5/WohmYrVyLNakIL0ymSctd4tmgugQx+QZoLXGLAD
ga1kVvDUZKTieIAGWQwObNlKh/VQCCO+AZQNwQsKTb0Y4d3Jy1eX2HLttfkZXB2R
0UBBQxsTT7Q5Vz5R2NGYhnflQOUS98JcG/jkzGsLqN4=
`protect END_PROTECTED
