`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JCRd7ybvGtyxkVuYqzqND+ftaavKdsve4BOPWHqJzVrf0Rk8PQ/59loxg40Sbncc
Fn+Bsor292KGxOHPUsQr3nTSwbN6GDUOxuNAAvgaZqzJLlHoUtE+x1sJyYxabvwt
JRBDmMCWQGkODhB2RvwdRZjw8UrVzXRepdFDf8bpt6794mTmNN04mO6be0dbMf8x
txD/RCZVzDxQV29hvJWGZvKnu05skTzkVO4PKVZLs8yqRFA3jM72K684pu0IG6y7
FpleM4Qaol0ra8ZAvn6mewxtZvePNV33o46Ai8QZxXyG288rr5g2d6pMPha6Od0a
R8eD8Qrk+3uVsJjmNo3M0mgvw3K5N5xkLzGtxeMwO6nneI2tduYO2ZG8wVL6IFfI
wLCPqFHiHgFGVNXkx9lJ4sHN9wKl943OJMEIwyrlyov7X+/XsY4urskI/nG93nwL
9FwpXdq+WuTF3gYW+UB8D/CrlQv+rx2SeNhkAHEgT9297SR1spwYp9EPfBb+K99F
tJWxCTFwipV6dm63CZoQF8dwxuK724CYjbH+vAXweas3jMqWVua1LubYRxbolW03
aHCRLxYOu/+iT8GiHYZx18KO4SdWrb3BzAAqSOk+vUy7B1NQvW3WkwXbOA5rBMsf
lF0fWduyj48MfxwQEJKmVwMd3VX1PfGGWtMTLy+RFn7FLmH0T+fUCrx1njPGmL7J
NP8rPok6C7aARnqPbus5k+Y8fP6aT/+VUzTLXyiGxeMQNvqK/whkjGql323RUfip
JHWnTNbnDBe2M5EA5s3Loe3MNz/SOQ96oyb59l45ifxTnVOzy5N7c8SDDP85efbU
qemPgkWawrtuJ0YFuLbZEXREYTbfvCNHLHaaJGzr05Pey8TUWztUvOgiAP7nYpZU
eoFNvyBhE50qubH1nog/KWlU5XdnfCbr3om6k7SfY6XfPsy6E1mo++YeQtqq6lUD
wM3w9RY7jv2ygzgDtEZ9B69kWqKIPhO7fpawfWAhX4dgWtU0Lt0M1Mf3ArRFU798
yRwGWDRa5LGZwAa98skRBDE0pmuHEBLlGjMrn5DI44M6xRII7bMs3yLf1l+7bfCJ
90FkcBLGAgSysf+KAGowXp5SdhAjmoA/M9d7H+Cep//tg4wCpuKmyVekgOg30Yi0
GQDNo34lac4Yo6jjIdMtI4QUlIJsdm3OPbFeyyR1ga0TIFtuf9MQ/Rjb0RnwfwZK
NT/dR01Jbg2Uf29wV+wl/UvLrwzlyr3HBycj7WcB7FwamMPpwMLGXNDgwRa1pSqk
160mQlT5E6IPjPlQr7tpvjpglnI45K5uCvCPUp3jc8XMw57uce1vrjd3AvIuRM3F
pr9jpyis2FR9aYdYlKxCJX5YbR3fPU3AFqxMMvnMYzyzmUa5Vei1fsn8zter9jsa
Ku8qGizvijFLVtn9b5qMCfdsRtkxNp4QW23kjVHfTRNliK2+LkmsRGYdkH761sTE
bqX1ka1+xTY/3LUXd4jNU6WP2/jCHjsdMAK4InV2xP0RaPm1xuKmu7FaAVBr+iMH
2l1nArcBreINay8g4F3pd1124z+3Wr+1QkoFRmkEgNw=
`protect END_PROTECTED
