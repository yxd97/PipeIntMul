`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VM41jQEQCoIkJEliZ3tcssky2b9vvJAyVaEZePdWMxnR7Li3zvfpkP8RqA+EdOi2
PodjGtDGmfE64YzEMa8q46nBEi7ALz8F8i7Sp04iAP5+ymKjbGZnLDe5KdVlLP++
zztN5jK0hVDjW52fX2CrB+cHgVmS8q1GNZPKM1nnZoEibBId1IESgr7BvMPDJznG
UIhraCLNUsHxHHntQkh98d7sqxOHMNinrKrX6Mdhja5lB1elFNSgDCGNeDiS4z4Y
Y+sye2nm1AJuXzLrOKDWXfYWvte5Hpd2T/1n9DbL3PekQN4YB9KgRfB4atUFn6Ml
2Wa2y8RTzC0BVDeM+oDqfwMq4CvBSVmlOo7QZLBh+eIahHwvjIIy8/FaqnGQ5zT/
oog3k2Jh7fSQAYmbjqPHdng9fYBqZxwGD9MSM7blfb5MsWmgk6lBN5zu+HV3/1mf
F66iRrG6JaltH3EZwDVPu89TYsZLvYF9gXypaij7OiXugF09VD3Ek/TTWV/juywS
XUWUWa9XwSJwsGzdlFrfhHeYTHJHRB+5KjQ78En7wEE=
`protect END_PROTECTED
