`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kkTT7srIjMmQTewG1+BIw2YjLCDtksmZWl+n14a4EsTZbeaFfm00Ed3r9yHgFRx0
hTNVVEmP+KRC6P8LJVgSTOifIQuEdILp07Tm7SNIzwylXfAzSF8gRy/zu0z4xIRR
IgH+93JP5ZIMy/69o6HLfyOAyAjx5m7ioPtq6ruHpiSZM0YHNOyc4CYMDgQszMH8
7O8CUSAnFGMOIEEdev4BAjsgbEREQjqnpaXdykoL2e8rYuIoVva5jksStEw0Ganz
jnA2PBwtSzBsXAS/NDzddpXXy3tESFlwkA+d530exi48XIV93bPW2BYGqQI0RQAS
WnwX5J/P2fPSWjpXpsJzNUgqMxviKQHQZtTwvRWx6joHcYK6aNDgiolbuz7E4DOq
eKjxl5olzXkBUkGTNOSWBloKXcBDGT3owaicrLyCQ75rL0nKUSJSwGZnlE3QdImU
yOPgVn0jAobnw4zzHMFSSKgjy4OEIZE0yi8oPNDEeoIlv9hO9VqUf4XaHLdWbBwO
zpRfA8S7UtKud2I8yxx1spv5o/C7hLrTX/KuvZ8KfvrpmsjAJooUl9rmG8h0Hd4V
vG8faeRviUw9fvZiHBv3rWDlvCRmk+MOLMy0tiUJQtZgNIoI8malj9EcLDH8T/YQ
l2Hw4takDiyqkNVIZNvf/rIFIp8u9wFYWvUQQ+2vcYFVOnPuARAhbz831OercByT
2/qo3vH9waduBjN6r6p//AxNZjqk9VTZd+JNk3bHdp8x+nclzR3NnmwcpiosPLPP
CWWSA0uB6pq7Fhkwhz90YhiI7xRY83aVfLvC0IYGqASV6ymBUieKwbNPA++GYuqL
ACG8NsOMn93eG5KPwD7wwkS6DCcB8M0yINhHkyYYY/7ImGHWaBd5aJRE1mLoWxOg
D8q+PeLrx26VIZuFz82jumayDA+HtfMpRTF+9PpypkvzdaWaFyFEPuMjklvqAmPd
/iKytkGUkmG6aCQ0Dbe3+fOREVha/l4m3uPJXsQI+VhOcy+cH/blm8TEYK7mfR/P
11LrqjmDZuFzTAScGjB+B/OwKIR/1b6QEVBtbc3cablw1lniIbZ3fq+20NiluibH
rLk/yjggnPIVKOWjaxo8jP+mAwZ2NS4wbqGzM4ynADNodCpyjuE6RLAD5R7NnrSP
SiSn0mcHo1hziTO/g3nPXxK+c3IGO79PBIMCbrzuumVBHBnOO65jkGDX3VuHqtBv
mNNVfwGEQdz0TC5HN+CyO7+KXaHVx+/Grr6hqE6UcDImrla7hEPA8xUfiVb096w9
fheAMqDuXwDqHP9giHdmQLpH8dKyvHhTmUZvOKRD0B6rzKy47FbKbXz0ksjG9QhB
EmcO27uv65lTlYQsb1ytgOSDRMPQBUccnwsnpeSY00/NykI852HpvP9wzxjNXmDz
imSsjIasPXLJuOvts5wl3yFcGeKBaO1cue5Fan8Jv8Y19vN/HClUczv+uTuPs1vt
/MyIs+DsoSBqmwf8Z+fX1rnrkkjCXR4H8Xun4xCDkeO7nsdX38UIxrCssgtXpLGe
jmx/NJfMLMDxm2eknzfU4O+TG/QyomtCMZX3CBMf+sBk9SK30jDuBBOD33p57B3D
7DlyV8QPlWlx/skqzv5GraPTZGGbaRaBCgaNYVaUR4PC/ILdnVl98GFurJrwLVd5
QOKoh6nsKcaMM0DEy6sxj6oA08NlBEJR0a12VbTutN2PjKzm/8maAwrhMFI3MiC3
iaQtQzThS/5+3MQBp6NJVnLp/DxXaR6gQVLQbOubajo=
`protect END_PROTECTED
