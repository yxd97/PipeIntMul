`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m2Aq7lUnZFRPeb/VojtgpLJMjohrAoHafPRXSnQ0zp19LZBrhS6J7ugDD8w3aRqN
6fQRUmcALR9yxZKwTvECAd+7Qv2+yoInZ6yEQuNz7kuzVReMjOetaj3xAa0hp8H7
+MtkqjP3QXHAeUoe10+FkuQR36+kVQNlPh/akI2jhhBI5MzAUC9dvNF4ERWeGyss
21OKaVJTB0eDLv+GZHdTV+eLGvH10PcnJfzOLGbxK/FenaqmdtjGWB8Axvz8/mP5
17kXCKjwRRekCTEN7g6DJGB6T5ZALkF3YeZKpYb34ARt/ri8zIXgkM1a9cIi5jcH
SVFQsD1wcQC4kxI+XdHtMrp2uc3gMLC6a0MMPAcapop0JB/1CKi9SM2rgi8/d/gr
bI2p6naW4UZmEvftePjrC8EzDlbGgYwiIskW/W+DOuxoe0J6gozRQgnjIW5R/glc
5jothazOqutTGzXH/lxzBimKWizqsK5xev2r2ZZPJW4YUiG4RaoNeh/Ndt1dJd+x
mYBQxXC5x34MBTEqBlrb2kP+a6C2BAyL4B/oRD+7Vk5YFHT+dRzfQine3Bk4IUR2
bDx2SWq0V+eriaCoVvc2y1lPaGIO9lBvGuBGB9+TInSpzV7K0Wv72QPbHsQJ81X4
`protect END_PROTECTED
