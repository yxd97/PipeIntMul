`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qXOo86hd4cMeKyYreOPgDcCp40UIK+Uk8VpfsPym5DlKyL2faDz7psWfUAv3C3om
AOJjIxkvbQ1ids47WYZHUMaBwZAnX6ct7CaGNAWy/7A4188+B506QhY+TDGKum65
To8BldfXN3pOq5wNXLVEdCWdKZFluaO4WkXFCaVzBtwXKp16dRA1FqHVheJHDU3t
VA8Mj3m+cTMkA82WMybwsr9NqVtRYNc2FONyRoSGf6iHc1r+QDL511tjHQPQg8Vt
47AwVQN58ki/8hnCKKuKArJeWSFIPFMuuPton+oVdqmEs29yEGXOq3znD01+dHYv
bYF0F15DawTdPahDVL+h6WQQjKnTmJVVQIJrZxVKdo6IFhVVYnLjobOfkZXv6FWp
`protect END_PROTECTED
