`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w6B+PDT1N4Hr7OxwNyoP4R6xoVeCMJPC18vjlPZvdYYbrQppwTuH02+CyE0UziaF
3215VP4UrRoeCUmm7qevqqZG0ntirYg5k2X+TnFU2kPxUCpvdNAHrqnfp3Twz9dM
NSXYRMWPsARlUQQD1GUTEf/14VRrEFTVIRs9CpqImpEWdELw0lkNIjENrBPi4pZ4
l/ot7fKaVNvB/Ii/bc1F6z5SWbeNAj+PyAOFnqldQJiyRKM/W1DfKl/y+uJSz163
YST4eh689jUhEd9DJTCdEU8b1Sg9KurzQNUSefzL3skYCpGDS4UBqkCS5WE/7f1M
cs8ANWfZilQRWaGxNwedRA==
`protect END_PROTECTED
