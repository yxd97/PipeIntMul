`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
klvm6oBiEWCzynpE2KIf5nDcOCvPsVctZJYmRICCN6JdaZedQ+t0uepZqrxc8ZwQ
fm9Lt8gr5DQZl63Rs+pz+YkRJgqydw0MSS8L1jQPsKBBOS2G7/3r20mlIJhjD7ip
BEDJroTy+olgqy0N43YUSqWqyESRP5JnSu3eeVpqJL7IwbNhNfCaB5VnigHmjPar
P3oKcZRogaWGwyFxYDspoxI9OsVkn24/BTE2z89aY9N9Q8dcnwmZlQrna2mmbA2c
V7uogrp9lgjTAa+FpME1PmK4kU9o+Dkm6QWQqz5FTCOhZ2LGzYO/PHm8z/BQ1Fa8
ar8ELdtayVuvcl4xsVx/xflWljhQ2ir4wf261hHcbVj9+LlkVQP7tGxz4dw6j5SQ
le849z0Yamf63ENrQwXLd1dVF+5vwle013QGEmDEfGTTa7f9cmLQ9eu0MEWFjUjz
CQ6NvlILygpG5+i4Zk29VstAhjC/gylavN+6/wBjcG0yrz93goYpQ9TonIjE511y
xYUw+ab+UmU0GTAvlCETB9F2/J3+mh2meUbTzXNVP27Hr8FiB27YGmswFZ4emFvU
8sqb5WbVTbmh3gpatpKhC+aa0bEUwQzbn4vUt6zSpmgeAR3wQfjQB2Wg9bDfmrAS
kgxK5l7IfQGzWchSpMt4Cli2WNqZ4jBVv9Gb5pcLHhSfKdH7E4GCcBci04L/gDWU
zmFtnMWKivbBzc70HY7l9u2nQExrMhNXzGNUg4WHdjTTrVEtopQ0ISOI0xbZIW22
5xiQQtHnuBglf61O7wyX+9mYSfZgAup8sz5cI7eYvr5AvfsU9I7BEhuuCy++Cmg7
oZcoduqMFoyDfngWfQg290/FFNklp6CojbBQCnrRWMb4NL4W8JIUpELKXw2IyKA9
Lxnub9hTpDcMu4QYFhj/Fl7yMh0I7MGRL+AedfLRMSzTsicIDLMhHYj9vIFjMKK1
SdeeOc0/gMDrJt/mmwTx0Ayc0qNdAThpm+bSzfjHiZyyzl55QtSgBdwDIUsh1XSF
X1XOOENIZFlCbLpzsoqn7SohKl1Dkf1JMKEP/EtDB15RzUeKKZVy09fdvcB+MANy
H5Yc6xb1Rxxgj/WT08KwaNMiaayZVH9Cqo+CEeSlhsMuSnaRUbhZ9Otn/qod71W7
`protect END_PROTECTED
