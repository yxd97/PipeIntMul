`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RvIv7AS3B76BVxbIqkt8v5DpqKw2MUWLeLJa79RFWcqwxp9hCnHl/T9IX/c8ADJX
ktlnaXYLCi02Rnao1uhToCqAs7WPQfXIySW+5j2NrfVww8ItYJEjgEy+NNCA6Vbi
ouV5GoDFl01179HArzmyAvKp63fS1ituympSXwH2+Y/l7DoupQLsqIJkHuoAre0b
sAOyhiaNhAOI4GIvac4XVUKTDkfYm/OwczFRK6AprIl7jNCiImrpxtc0FOM7HFhS
+3fET93+KK55bvTJF7xvFS8SUH+fPSNADnrIoKTf4Nl8xgSgGGBsuCvfYX+dVSVC
s4xpzJqwF0ShPOjwn/KMSaWNjMVAoNQBDV9hqK/9Vxk=
`protect END_PROTECTED
