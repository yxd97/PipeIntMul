`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NCk+biyYBAKZHOntu+WGIX/3ycje5rKTK8ZG9FEhBqC9bp+Gv6oZ61LOlyWBUIX
IsOGK1MzbtmBdQG28iwYTVhNPmcY+fQeKPOksVJM66IVvbmKK9UEN7WbFgIF0G/r
yGUSffQDStAJ8sDVToNlGfJRfkJYLZ/3QoYkqPxe5UkxP4L4uFLGXV4wXdTXMXpa
nfsFBFZ3XmKQR8XaFYoA4oEd33WXpdpIIe+Vir5RD8xjSeuH1tVpgS1huC9unevv
xEA+ewqQ2YFPhh3RtRhikUk2ragNUiiYkl+p1api0JF5NXqbBpi4AYwzTDhqQvOD
Z5qwDOPaOR82fTkqtRX0RIA3BkFXB1R7//0BTUQZ7Qz4XqLVOVIdg/dWp/T915qY
uqkD7/lqsIere23V/L4F/H/SDyH8tw8LDUHTttGcHJNT51PqWcXnwdIXd3zqYdGO
qSrlvQd6Nsg0SL/FkV2PvR/J3osilQ647SFmIZ/FE1Odyczqg8SVHKpSdXvijCqP
F5MVEfhjSgSgTmG+0Wv2+/kdjk5ViGdzKQtJR+bOTby/zM4yTg4JDNFEUpJwW5w0
EX2+D235DtS4Fyq0AfJ90OyZ7keALYc+42ufQ0abzNmhpfIJNluFWdMmzq//Y9K9
t5I9uAdPt5AztLQjoDydPrI1c2GC0tI5tvbzCrnMYkjGX6fTVJWvqyX/o0cAgubF
9hK0LI3hsKID+kpibIiXn4MBMUepbDWaCovFRuZY4OevgA1WDCoFue4bAM0+ZMt6
E9zY2FvYNFNTWEi0jx9V3vRt3Y7NGOOiS0VeMkfGEBYhDIyRiaYjrxnWFmIldcfi
Sqwv2amHWVazOhEFYT/zon0eC1xjdD5daqipb6lgM/P5CQgOpJZhEaDSe55k7q+v
LNYFeu/U/bJjYkvPZl2j/P68+5HItPrq3W3q3ZzPAaFH9VDD4E6pN8qpboxAuuNS
7Rkg5It6KTtGDY91kj70DynJJMwIOpWFaWITADosuQ8wXBP5quTax6KI1paQpR2e
JN0gqtwDMhMujLX9zvogJ9N5DjBiCQ920pKfMrsS9vmoXksVk+RDFpQ9SwfWScIQ
9mMzVCHWfMeyl50BLiC+hkeL8G/cMSSDRM3NP3r3N3A=
`protect END_PROTECTED
