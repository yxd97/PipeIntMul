`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bpdd4CSjNu11OxbwDbxhBBTwdNkAIGVr8F+XU3WbX2vtWKiu0OTZdhjF+sX787pR
jKoB2+iMLuAzcs7ZFHYKyFRU0cnaIg89ehOsU0tPLS4gG35n+cRYzZKYm2u5Yv9K
+S7LMTL0IZ5tFP3Jfcwu6GZpXKwcsSwkboWOacrwTl+cBW6WBcF3XWO15XNG9S6j
feQOevybkGR9EXPQS3PrTt0mHVjr5qHV1KKOo6xNt7jMFxVKnA82t2GNq28B235F
o1hyBd5kt5j5ENoGBawGyAD6xSVYQ2JJ5rLjyYaO3/10FgrM9vmiGtJPrPsFtu2F
eFfCgZKnyOVke9hy/ntq7bTcjBd3DGyZFePNzXyiPTskmDK9rJl9glJfHZPfdCdv
cQGk/Cs+rmXsDM38VqBgsRdoeequ73WcZouhat9EakzXGAOM4MevbEZqt2R8XVdz
ET/+f8i1VjaGMaLswkXZH9nMbjtR7ddP4mRkXWcK2bpM1mHJbuhPUmgiCIF7lNpq
pdxZcSRUqZgDY+OvCzJ0YKEwSPDGUF6KJkHfjAXislsnNlPerq825HE+PElNJ8vQ
JKaJ3JoSpcTsk7dDVN0O/UsQ93pd0LjWMYyIXCw2RcwuWVmRf38OH2UX0cYOCkSO
8qEkfkTcsh9y+Ocif7NduPFawcRCMv0wrOoW8BEVqfez5sePTYRIam0vy88cQQLL
K5CpSuqLeFGV4+Ktm15ujlOJSnaVFbYDMDKSzj9cI4/FOqbxiwVOfxgNiJIX+D0h
rQQOUtxDBXN/jcGtAoweIcxDv+LtGRzDG8+i7s/TosHw0wY21045R8X9hG+wR0Kh
G7cLrOvF2vQ1IV7zsqLEIpx34KGJoI5wr20vvFNppiEcwR8bGHGTbCvd/Jk3nZtg
T7zjnsdJ9RGYdWnHy7IkyaLaNYhvl6TNcplrdnxJpKa4izp/ELixPWQIpAJK3ALp
tgTVbxb3XQ5L6aYZwlp+AJOX5MpWUusYxWdROVZobuFXdOUM/B/H7b6NQ9I/JplQ
`protect END_PROTECTED
