`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wU/RAVYrVxclgjtjDR7EFK2B4/v31W00WfcoogulTM5aqpEEQjJhy84mcxZwNX0E
/y0M3VmAPwgA1vrmI2lRgDvK/Gx70U9KhYRxpv5ftDK85W65Db7y3bCTpQxcR21l
Is+jEtq2ZJbyxc3L9jyVVqx/tN1PAoXf3oJy+LQdrHp2ItI1/QL6deR+bgHNL3ue
rAeYY8E9DQ1ij3599mWfL7XoOXN0MAUtAlQnk3zhq5A91swg+KWbW5TEcAtaZwYB
72k0g9Tbl/w4dXFfziBP3BfknQcKe4w/AH1adNW00OL4/WZP8QsvFpV1dh7qToUh
zC8CLO8z1u8nrz+0UR81vxuauYYZzzVfquUocrvm2baGgzubaH7JkQCFgAHNud+3
9BdyYee7UTJiZqP854AtGHdv7bGQWtN9U5FK8ND5vhwa2zr0QjOeTuCtEQ0UDOIT
75jV5A81tlDLe/rPWrOdnHcuge56Fn2JONZ9zB0Z8ffLLIAhQY1pjwCg+PK6u/fp
dfinN1JwfqG0tC+wi7PuDYtZSpFeTJW1D3+P/V717AuJeKaSbEKygi4Ul+8zF1KL
0LApCbwMEo9TdgEcciTQQpcYlx1wBgFQxHXEAAwiUuqYAl3BewMnp249lSaVunFO
m8eHTjcrSRhzzedsgjA3OI+zH16iA/BOvbvZJSZIn4gYb23NawVYxXItaouhw38x
wRFTDxDIamhMOi04/Ad+Nhunflk+Aov5KdQVjpTRhDSLLRQWOt60lKo0b31yWa7R
Ut7RW8rNYFlzomBvJFZVwiarp3F3eARr203V1+nXHMF5FFGBaLNrBJUiq0lRffYA
uko4Qd37sfctzK5mms4N65/mmJfrzcJzskIXc55OusOvjJmCS5t5eQVPj0xoqKes
8HFy2AwUAMMjMTXf+jBXg9s+VHdQ/YAudcfIrSPX6tdY9JQGwdPM+5y548W8YknQ
EXEntmRWT9QvK/AJEk0eLYagiSWGXBMVaU6IHgzciq9Z3f9NC5ywYtr9dEmhWpF+
pOc/qa0aJgUoVgtvYcBsdnybznWrNZulw2DFN3ZGnyCkV7KxRtYqkVT3eZH1F/HX
VgRpl6qyvuMBMf4JFVmoiM4UGboHY6HVlFefkxTZwgIbQh0kRtXOOJC1L81kMR5r
Tbmm66DXI3imYro8Es+nvfCfcQK51l+fC/TjOxaUTsRWdas70zH5yeeTHYEFH3IN
Htg1FhqrRrwoGznZTPEFcwkQGGsUnq3vgXFzAvLwcnmkoKBhmr3ztiJFRWvMO/Bh
8v6Wz1OH89f78JlGw0P3b0WkuQ5Jjmm8aJborPRg8LTfNr4rQVHiSb6lG5MAxL/j
1iTnWngysg0WDY1WO510NJPlWILXjYLz2ZauxwCAPzmFntWXZQ9XBmJnf+9mXbL/
+cu8Oubgz4dOd1J2xq+SoKZwMpcJxYX2CxND/b0jvOHam+HOCg3kkyYmBjksoK7c
1sb3XwVUrA8npkhrew+sZYYOT6Z8x0i57n+eApGR18KTjeDiYRLlj8TAVoUxc7Ro
`protect END_PROTECTED
