`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
glXey6BnTd0JVMWTRQGm6jPHq5MH/3JNGGXVnYFzukQJcPJ0d5UhRHWD/vz8do3/
ui5nEetXxPWUuut5bOn+Z7O7f4lEVK+4KF9ck8dKUcK0lyJAjzDmmbzCPxsskgGM
nqEsQCg+AJDI8uEjra5omMeuq6PZDuxq9FjN8E7JPUXna90ykFBgN4Y17uZYHimI
ZBnafPHMo4MOpwV0+2C8MN6Ed36jqKdIvO7XLbLg5T73oVSbZYp27HdouASGVKHY
yhRZh3nKeK/GiNZ1CEec1xCEX08nTnF0sRewwIHT6ZKMdumSm7ULKCKlneakC3+t
4pGjuEZijPRcEuU43MbujQ==
`protect END_PROTECTED
