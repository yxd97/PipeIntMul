`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nTEcAMssWjdEoXH3fE3mwxUT0RJcN/EmaT92VTaboNtAn8zo7zi6jfTjbbnvZ5Xa
b8ER5WgIDTX+Msxd3FvMom3wXi73VDxVWnHAOsSEK+ktdFYonNXyXJ5cqMf9d1fg
3BNRsZxw7Xth0YrENr61ufjUw3ZaqJtrZqQ9ptgq+Gv3stDgoSLLK+/V88XiUQuK
Gah3wkRvtOBgVFwGaQUSUbePz8oDDVys8hGdfkkKXITwRcHTeJjjwRHbd6rnv7VO
tTGuxp4TdM9M2X1GHTXKtkoDXuRt43JuPpSO/6/sUSLQ7TeHeL5+NkL7+xfoQb/c
eb6j146SMfqPjxU1/7FiENkCyuZSqPiXTAxMoqzrDXDKO3LoFhyuVJo4cwUaRXAu
K9l50k77TixCu8WNnGafVPY2Cn1/Z+vg5w6ClX1zLYZtLcMQG83jjMTxAZbTND9K
MuKd8J0T3+U6sc0zoUExFncqmHMeSCE5VCygvHx7sVEcgjGSeFRQHj4+BWEpT7gv
`protect END_PROTECTED
