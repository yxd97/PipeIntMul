`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6Q2TsXd6y8ZvdIz4GVEggxXW8fjiu8gpQwwzFJhq19i9BijKZi1BCK7VVxivxcg
6qiNXSzVfvRx62OAQcyLYZ2gjLlHmxlAHA4e+BJMP6goics2qXkT5GLEUI/KnNqv
9Y2BAbPT6xy9QoOR1vVr0aQGAbtwa1Y55ByrDVdeeV3NBux2/CNDx5IIv8onoTxM
SyxKsKSn2P6U9UoVrPif4s6b7YoLh1zXLkBf2D8ShlTAH4ES5JcHNIP6MhIIDCEK
sPoNtaW+aY+hTZGVkC/I2M/p0R6RCw66wDcm5W0Wq3c=
`protect END_PROTECTED
