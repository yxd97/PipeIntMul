`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cLqsfPNXlSel146WzR6ir7NzkJ9eswxK0S04cLVMTvTc31XCvt6YK2ST7LeQWMzt
PBeHal74tm3n2Kj6gNxPwoeIwob+eZgHi39ysUO2xU5QyruS+6pACqCCr+cxdn7n
CTkiI+eyZduyLyJvTfXSZ+wDeg5jBOenhrHuEh5hdQdbSzidjeicu8OZTYg3feq0
TAZLZn+GAOIZSljS1DK+vhetIoCCzI8c06ysXsEm3g87SKdBRGpYmZL9LxQHpnlL
YlsHidqMQzfP8EbEmZZu4A==
`protect END_PROTECTED
