`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evIWfN37lbfVao0teAfySrPIqOYGYv5Gg2sfc6RKSAMDcHXGSZNEIprLo/dZxRcg
r9W6JryZZIwq4P/SFBjw6RcnfEQzEd1jfS9tNvuFLsC/+UyvXCT6wZ1/2OKUi8y+
8yUGueycwg4tWLFGT82UOq8kQlNUfuLLE77EzMLI/oY/+zP8FpsESBzkU/of0UQJ
BfyJmg89VzKrywxFU52KB2We/kEBbR1lhsXA/UTWF8JiCYXJyNPn1GcTkFnR6XKW
G24nP97kkaF+xcnllHJZm7ZkoV2ZM/GIQ5sc2g3WSeWxmsi+kVBcT/5rtr1dmjWs
SJyD2Voj6Pgwq+L4tB3jAHGmBE6qu5XQDCME3ULu6BgvGX/STbHn717yBcrk3OAy
qTSrtUVlbV27zk0P7JzwAl9YsgM3RhN2LHyQgDhbnZWsowWmQEgJOFQvdjm8OqQL
kE5i6P1cvdlzjFNrQpmcmKm3gSG/JEX/aemt9+iLNnn5HYjTe80G6ZaMCPXgU+9B
g18mBxzFzzqNDN/a7W5NYw==
`protect END_PROTECTED
