`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlgvJFkUS0cFEWS7zSCcrzI8kJHLkMic8QWlv8SVplaQg+h2OBGywA+vHgnLKt05
JA1qCteNsbU2EiuXMc+QOuttxx9h2jzhnlJRBME2YoTSJPJECQugYZnuKJIPit3J
6qnOEHmTQ2KsGRcEL7AOJ/0zUoOHPNi0CbQW9spQIFaHmuIC4Nk9K0SMzV3tuUPn
S4gfIxC61o8KzQ8p5lbZMhNEPG+3nGTq7YpK1RBhKh3oS3fUwQRpmKFT1vZN40aE
elGuTWAkOdHqAJmmPR8dHOhQTUknnhJ//iYbPpOdjqFE5839OlGFnFC25Mu4X4z8
eeJqlFmIFIKCimq24SrSV2vMZoAQNIhb1k5LYH256PzM/WV3/Sog271vn+C5O/2v
GNvzu8H6PyXYJrZaUKOXI8A0a1r+8Bc8iC+fFGtLjmbQns8O+tA9orGctYyFEDq+
7WPJLE3Q1u5oVdNfvWazz7quMt5Sct5TKJ0frIEVv/nE2b2/hZcPWYlKOrRnd6RF
VIthp6HeQzemFzGIEGMuuBfBgJuq/B9jPUK+sfDOoboqOwfXjgsiCaRJHN4XJ2Jk
aVMnmax/WGZ5zpLyJidHAUsPB+0wl/utJ7R74uMuzBE=
`protect END_PROTECTED
