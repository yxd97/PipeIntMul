`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z8NE1tWA/xGbuFXZiaMmybbGDcCuy1shAHiYIkuKZTbDQFp9pgSohRClOGKZCcN/
zafQCtJ8F0kRNlolWvry7Mq4OF8PqmZkbJuxM/YJyvTVFKhtLmQcOPJHeNgUyXc6
V2CV7fU8GG4JVMuWOdK7vgY5n09I3IicYdctCqp2goJmicdT/vRHszTzsSwY1QrT
ky/TX3LSElKr1mzEoX31SlPRnSncGVCtlsqO7coJVu33CbSPfmG5RhUEnHMbuQAJ
7RKBwlnGI25d5zO3R/bLJcLYKkHOVWSXHSSTqq+Q/8sgHAiVOZ0+P4cpfzkBH0Na
8Mt2gcqtjvK4oNqo2LZZhMZl+6+FwAn5bug4w8VjfmaWUjI2dzqbIo/bpsksgXqz
4+w061aphHEet/VIbLyAPjAm+pYIT0/CgS0bmceeEx3jJBfCES2AgErTkZUGXaQN
JMOF8TniNxHOIm2/wirHKptUNKmwoUI9R/loWR1cZ2QatFcCv3pKduDdyd6dLB/Z
wnyjrmiDQgiAmR7PqIeRa9yV19Oy+FFutfkl9QadWWXuvDvtmuOK7qr4615kUdgm
njJ9aAh4tV9Dr2y6a2/HYwsPqMMCs+ZDtDnMhrYcYr3/dL05tlw5B0cIubcIkG1/
sTkGZERDrx4FJkkjxtTrFQe4L8IMiedrn5rPnL0Qlcn21V7N1s0wBkV8QCpN6haX
bnoz1D9Ob4dYOGB23krEx/avfS+ysnYPPqa5n39lWeRRID6QzRyA0wYjCS5YlOc9
bO4HyO3NRO0tdAPgbR8GBg==
`protect END_PROTECTED
