`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MNxM/v6VBoSw7vIDvyfcuu+mP8d9yD1RLlpXz2181FRwhc2VDQ/IlSnXnn+7kuxp
XAL5KHxRsLji3Fl6NyP/z/4bJJoWwSl+mh3oXfpMSrANmW3ubdbQ8fIcC27CIddI
B4/GhVnGVhJ47OZDKLLjEGhZWSP10CEC1QB1B1h2YOHONgM2ezPEUVEl7KSSQNUt
CTqjawhIMegpkVbvI2lkvoJj+9yMaU/0chQOXhv1gulihCwPc/UxDyA3KybnC9Gc
jrepUzQrubAYhTV3Ej98Zw3GbI03aZLdme6xLW1SthVZPNE3+Rh08mGgjrZg8uW9
wLMun3QEoDSB8BMkrgBQO2u6XUY0VYazG3L8Vn59UAHXs9WkN41+KfKkSXy8Hwen
gkyu3v05oSU2sT34UVkUS6c7e+g/pG3fMjs+PthuU/IfBG/R+jg8ciBdM4/FbVoG
ssWOvVS9ePFKAK/JjODMSBkd4c+n8Yuht+u7cRzBeATTdFB5yVdxKX7JdnlDpdKE
ooGhskmb/gd83k9Ip+1HcfklrL46+6AhFf5yVeE63mfxJkKY6RAFny0yPKe5T3op
YYBfm5rllfeC4LeGm6hvJAZvD0OENPwLfYPSa5egttOCg5B1Iv+TAJKlQdG8xx+2
AYkTclivv9HKog5CwKBTSgn+7R7qrFpppU+YFfNS91lK8gf/aCcYVsEYxpRLONqu
FzSvTHtpvWqPGzh1ZDZh2360a01iIdYU+Ph/Mxbf1xWw7FrcdJxKr60+ZxgZrcWq
tJSuQUE/EjLxczzg2nnNtg6XWnYDjTwep3ujFt1C49w7zgt7q2deItYofmBx26td
z9ZQ7KKOYc60VSXesqlEVeqLOehYmB7/i46FNNcQo2qyAJDX+VHd+zxoJ6Vck2jO
+I8VNh5y9A7AiVJSciMa0fV2znx18TRYsn6oIo1SXDApXYj1vx27KF5qvMutl1bd
+GxvVD1gkFpC5QYGhDX2og5QgB7BCNWzRLnhY/cj8n+Ol6JFRF+JV5WTaCfWEshI
P95JW7+ePJcBaQq5KXyUHSzXhcy+gGLXp4Q4JiQSeArVturY/OHYFiVvzpDDUUzl
otPY6JXLfoFwFR4QqbVoqKSMNMYqKNWw3UYwNw7zQNnbN7yGd2hmZxOh9nSlpXkl
oIOtCLYm3+V8UPaxArBFrMdfooywuZ2T2xeWCmqsE44ReLVv22v4AlbS11GoH+hj
3UpI1Z5xzDkYwRWbBlAZkJldTNbdhqTIhvnKB8+XoH7CxpLkd59RvTaLF6xuf02A
PyCGfkSDVhkBvFVmaSs5ltcHhsqGs1cI9CmlrK+2htQ3MH8i6VIF1u/IH8TLft6A
f1rcrkz2fIC1S0AA8LNGqun+0CCFaQihEnB0NHTxjY6yUUKQA+hCI8deUlypstfN
bC+dKYlLkvF+V9US6opbPayaEN6kzKTeawNlBJ0FaL4/0/avzzx1ijL4Yu3u+vvy
ysysGmwYxNsg+hhHWSYygT/hjvRUxrX/yDyf94oWuY7km54vasXT0tfMixy8L6lm
V/43Mm4Uve+HBTWmkEGN0Omaj1LOdfyk6m3CbAxUaT/5bxvNxwecngTQ0RxpdQ5S
nC8ggYTRcqH+4Y18c5NdMZFT9ilfIcWgg6i6hFflnymzPhewXOCBIjRIjwrf16AQ
jzznTRDuOrp2KrmXapsCKKbAbeNEHnId52uwS9ZlLzsTmVVE2wvZIzq/t073+QBx
rtKVllBqzCPPTDcEJACLV8ejwsPa81QIvuTqnYXG0nmNHS5IiZh88bHgKE+9HVSq
pxbF1NzAxs4RDpHK6fvKygltIhqOrKk/iRNPI/huMFbgSOf+PQhXVXkKZdAbmryy
IDJ18ySN3W+0fXgWn7nEizpQC8Oy59xjdN9nXh306Q9EZA3NOL5NtbBQQOd+6atl
DATxRsdFbBRpqqdkOQjr1FTzOwYr0vIIzJq4mJ9mi9q2glYSeJgC4C1a5B0xL0ns
NytwMProTJAnn/iQVjcK5CGqa/V+ESbsAq1TGgE0DxJV8PIus12lmCJ2qu/rS6gD
9ia1vVhjenOfXiNtHrgBla0atnRPjqp0E/FAe66T4p3ZWP5kS9LxgJSST6gekhAb
G3WE4CkttGG8ymvPdabECKhGaTHwYhW+j5IlcmcDlWP118oQKjIs2+1VZwYftPnn
6IY9MtDni/COlUmKPsPNPOoTZD/39bOv/V8sFnRgozuLtsBLeHG9ckup6Cm1PYlu
nPqc/+X6wg8GrI0BqQzpHulKlz8nnJY4iyq/bYyZO+pB65qRg7RyruxPWk4/WFbk
lff9POQcyAw2bPj29GRTFCJMk07XUdkJTQHYTqmNYGy+kf4oq31X0alntgmh+V4P
ZnVE/6ymrD6ivRn3LLOkOC3AEcSzQukUNbaui1sCJ8u1mDIjPdbVVNU6ajnbPXgm
LHjgRW0P07oQf0A7NuveJ4vY+mKQAazKbk7tr0wHhBPWwkOBI1dRzhhE9XIVgouA
GLEVdUYRJHpiDR30eRLtVtGpFPH2iiqzQMbS2kPwGUeIURpW3s20pwuXFldqsQQR
LQyjx5StjkWVIeZxSS6F+6BA6DfQIrrZJH+qUUJHxjnTQXJ3JByjLDTzdTMOqUPw
0+X3k2YLpCEl0KxVOsphW80+tBw3/yi94O2O7/NuscQFnRqlLcwWVbrLaIgtYWrs
R9eJGET2HczS6zKzYcyda83cyWSknTCNF+96lTC4QeC3mU80sanvyfKoP6Emnowe
4kUv2AC6hl1bNQFfejK+WNDDriDM2cvUIT7Hen0EyGpeb8TqQ7+wNXnQVRmZe4bB
aJGKymCimkpLls/sZr/1YUvS0S29FqDJVehuma/SgoQ=
`protect END_PROTECTED
