`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j/8bMTFe7hKh+cErtCAeHLyy9AWxkpILVUxA2Cjeqbzpmvi8cgPhPixlcUBf451o
qk1OaiEQAjmKtJtpkKLQl5d4hbi5HSn5hOjaslW0hpyG5w7cFe2Ek6XfS8Gf8hi9
3DM2cz/lhG4Adp1NOWYHzVOZKoqza9DGE9wUctDfbVk44LElgOUPwpcy0WX5Aszj
rn5kZevqW/+OYaQGY8CaA1Ssvyjh/SrjLQiKtpXF4dBSr7Zw2jPg4rzf11ZZAo3t
IY5p41TX7Vnc2erTSf0o+PrSFHWoUMKd9XD2MCFi4wLmILBZZrb0VW4ExNOk5wmV
jmOaRtUgdWUWzWBPKzIV2gUjbH/O2alAgmbhfVYS+AgMvNlWxTl22EK4/gJZP9bR
`protect END_PROTECTED
