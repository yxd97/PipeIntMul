`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DVJGO9WPcLNI4/tyX8wczXcWE0ofvOoonTbu3SMWOmaDtNIam10JFHvLQJvH0IK6
VICzhO8bgjDGWzmjiwoWcx5Y2Qk68yuMUd72fxHROTfIg4piBY14Qyy/MJYAdzFn
akcYx1Mw2A9Y/XUAVIRB+AgbMbWa6L6doNytPk4wmjU=
`protect END_PROTECTED
