`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZEmXP4CfxvPDLlPT3hdBod9GEhsVbgpzaOAm7Lus9y3wYSfPtv0joQK7o9ygPxS
mtsKSxb6BJDTGSVzMwDKCB+9phzAcuZ/9mDefgFy9U9aj0l5h2QZsrSmfdsLw2gV
MKVpSitPF3Yq5r88KI06AaBV8XhFWn2/2HCKoLGIWQt3UpU4AV83k6AVuWVzr7Xn
HGrh/KUtMcDYg89asuyFTALQPGUbcvdU/6ETXTPx75G5a3ZEveSB/qTgloMmzaM1
OcHS9OVrpwH2q9H9x4Yrz1q4jFSf5VIk2sx6vnSrz/dhV9Au0gs8x/0qTJ8oetij
oguEdQ3PKFUEe9bKc4EpbfTK6eXVc1XheOogVmVARqljn0QoUP3YDHnwMZ9IPpnR
M3BAWV8ffVArYP88E0HEE5nRyY+lPnjdtWNAAZZeFYoo72kvtpAH7IjXTodaml4e
sOZoAJWLK0dCmRjba36GcPwkiVdsXCkNHTTbFIq9aEOiQvmNnYRCU3cMtRHgmHuv
UXhWEcHGwwBd5hpUW7qDu4OUVSTvTDSg1itTSTMHA2jOv7LxmgtDmaZDEDffJycP
dpG5YI/tMvIL9/0uZVXc8Q==
`protect END_PROTECTED
