`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GaAoEUgk5UxEbF8DsIuV5+4hy0BJtzaqBcGfyZfVbkeqXrrB2OFnKc72eRQXQ5MP
+mof5PRMho60wkKjtPww99eUQhQbc+DNCBq9VxGl2TMRrdwy3I4Qh0p3PeJt9efv
cDvK1DN3N0ReWiXiRXdFqFtUtfWgOUy8OegeQeUcKossoOc4mueJk0lHkwKklJCS
+w8femAsMXYb81TqwJ8x8km7TJR8MIAzRnvWPATTuMg5u7rsl6Oxu6UmANWKmyEC
E5xlbMJv3RIUJgg0CsDqLZvCF66v566+IxIclRB8yuml8eATr5brjkVXi5ZfOa54
vFzar6ncQ3aku7bcp4H61cn1T1XtqY1iTmsc8UjmYmi+lkBaqEHj9mOt8pWuBgTH
/ANXdz/XV/tV15ioIc8uIG+VWCR9EBGDk1XDXvKdkOFSxf3FvmHklGeCL1ae4Emt
cGvHKYrBJ0y7pK/4rAnRFe09gFHVPGkJT8Ed9teul2o8oq1FMq2KS8hexZsgrnLL
BHrHE/dKbv2jDQ3HXYcJRY17toHtD8GvN4ny87iKpto6bUOc5kO0p8IiIR/tX2vm
WXYkxibNJQ/NcDpsPGGr43KIsIdfSyz5eOFHh9bFfV0PjRtN+KcCt8ZQmq+rQo3m
eMfLMHf/rqA2KQSfqySLzLU9Go8ADSnMbGIuZ5MGIrk/HGy7PunfK4f24cwG0JNg
jMcN8sJFMKBlVzazC90TOUgAFa9oGaHaINOR6dRO0rp0MyxVPtjgIfyHi0oaXLIr
C7COe0FtxIZ9KpexCOKlJwIlR4PXXSLKjPwbj2+7d9A=
`protect END_PROTECTED
