`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SbzupK27WghJPaYPyw1SFXuE5RW4D8Wf1rNKMSgcuY9TN9ZuuhHxxvonENRqmq9/
o3I40qH1YQW+fVKZrj2C/S84A+zEKLNUnk3EcGYVDRNF/1Xcc4flWEydc9fM7Se9
fA5OCI/PJQFMkx/oxikTsy8cq3mxtFrst/MpPCNa7hBk8kAv8WQ26MarBziO0coa
vMTGqlFK+rCHGS/Kky06IS044lH04nW8XjO5XFA3nM9qdQkEnNL+o3vhKsPuK56H
sri4Nl2a8vMThNAni4IG9N3y/lUZxIBUvRtK0znz4r/qaGKT6TxOnIhLOOpX+Rc8
kEgRMN//CCEESemNozkSIOrIMfNyxXsIeEeq261U6Fa7sppJS94f24VRN/qtwMGE
U+TfsB3b3ALPv1wuqxhzUuiDlOcrzRENFGIE6Vks1FAOG1+nTRjId1Sr06krVqH2
Fztjp8Q9tDesdOyAbFe6sgk3XY4zCVUppMapoOYNfmCaaZ0N4HFiYBd+OCzIQXBP
NXeeXjRZHMQBpwgaw5Caz5Rws7gF5V1xwZT1zJEMeqM8uz4t0vuIUrio62dIuS2R
KCC9O3lYokfIVsK4D9M23VbmW5ZTfW0vZJBAMRXsIwb01TFJ1JrnleLKqdj2g4+Y
sVR9VVoRggRAYgrmoiTgopwarFrudJyHmesj92EC+pXTvce0A7VfyjizK9ecugnj
8JjDV6IICfWtLILqOe4AUTP8seFD/b1pnRt5BluUJoaADDjKO77VnHsx/li4MAYi
/QuztUiVzigb3YC/uknpSJX631YILs2fTcJ5AEAtRj9J9F+4tUJH0NBADogRPaqA
FmPrfiKzFSRazOhc6+QSO8fAYYFFo03+l6GBUE+e0TZQj0CYYfPgcXRIZiVH+mIn
`protect END_PROTECTED
