`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/G+ToxBkhcE5yklstjJAHSYFRbAmYKfgW91wASZWhz58/LYr23L3tV6ESlZpukqG
rEMNgkX9zzF6G0PrAim1RiD9bRGALjgEi4SfmUVub8B8RZ92auA62YcU050MrEzX
3yW1jzuyspMQ99OVuVCRWr8L1YLX7eAODgBrA+RZPEuv1l8Kz2xE/99V2sl5daUM
AJMOAFX9Ivz02YD/78n+e+B5PFFHPKZw8WysA8R0Bc6GmOrm2i3zf1kn+kksoxok
4cM7GW62pQ5eqpeZcdARVn0Q6VPjaxFoFUQNFmIEABRTPmr4jXikJouUgSzF78Gt
uKLodVCuJJtO94JvYSV0m8BDpfhVCBPN8CpLhRE7iHJ7QbCnJXm5lWrryjtuw29Y
jFT3SuWgccFnjO0X3F+TWYLf2IHyK8PwUU+BNBcZVjo=
`protect END_PROTECTED
