`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kYa+UsGJ25ZrajeiCUmjzQcwyG+MctwPWPjlocGdiNUBbHTQ7QNeSJdKAlfw40Ux
z1KBMCDgKm1+tyO6v2AhM1FAnm6XHky2w2jXGCArqarJRHUvwk6WVhLNRyiMMl+W
9vR0byZvON+eiWyVXwgdN28L7XYfxsq8B3xIE+vd+m1rt6cXG/DD5nYMVWy9fqW8
PIquCl2VqnL3NZSYiQpF2CjmjTbhcRenVtyFY2LeKqWBli8fJTe/ZyBKstHB3M7f
3TT+Wpt5yJKKSE3I/7XOmSf4kbwBqRPIm8MQeouybbnp9Rip8w+XXtHqzAGzJum6
hcBOgqpRfhS7wUcbkpd2TOiRZlD16Ucy6CX02iBgLDNo3wZToPTkllNOri4xWNRO
48NHrb+cnHm8RSPlLXkR1yO5CybaJCTkDdRbHetQ7ZdGlUckzlXHFY4YA3lktdlP
CkW8aIX7oHdf9U1oX3vyQY59fX3JIVISk6DEE4sxuhm9AYiayKG1UeR2R87PK0QJ
`protect END_PROTECTED
