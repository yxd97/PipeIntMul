`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5VqYY1elzq/ZtYC20vO6wiFjBrviTvnALgxOjK5I/qXvhpeEv3VIJiptr18YUkWq
7oZ2+7Tjmku9GgnqW1C0D2975LKwriIj2gPKysr2rDGhxgOSVzTYQXU7RpfMDbkR
iRw/WHHpjSh0BP+gHjtk4nubJ7p8LoDfw8SbH44kzBhM4MHkA0LXhS7GYnbYcEYu
PZ3SvwWBnrMd29K3zvuLagYVdLNuw9OSNpZYrKRXQ3+4qgQrNsiK1Cd0sHBBEq0A
PfTzUKOa2ddZm+DIHR7VHYEpwwgEVW/HMdJ+LoFQ0o2Dku/8FXCWv7Vs3FJW9kjT
KPagX/WI5vQ44QQQkRF4sbAc709D1zuV2sWAGMnHs/998x8XuL6jf63pc26megPk
PQEeom77VPrAXmYVaRAYgLeeDLmuiDJubCzf5t6LXMhDmdSkK/XAIqdUOifzUJn1
99ekdpHjUz40Dme0YtNOJqhQpRNC4FLRTx/B4iPNwuravyRo5W6uNeidVqD5xq87
`protect END_PROTECTED
