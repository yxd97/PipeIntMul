`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yo31a8UaPazyB6JEfmyLGg+dWF0SnbviFXm65zYHeI5AgTHLSc1zXQJUGxhFIvCd
H5Y8+hKIcipnLAZ+mYGsOUzbfnBkJ/hS6A7o9cCI2l6rzl6Fah3FX9gTe8UGsVkj
d9hdxvafhp/Fn/Z+aPm/cYhkgSPS0fXFk/Y0AN6djSBYoxVxdungCVVR1sPmpPG9
cc/kZgELBFDXmXni5I8L2dILRqfFFzmFd671qv+8hods4wzzopkcfcEM22kAgYjd
O5pZPtlw+TZt5O/B2bzkdMhlhNHhDzZ9i8pCQTW/spVsIK3J4an5cZwTG0eRRiX6
lxPnHPBqRXhD/Z7HQCXqvv6CDGbdp29nchpGLjhvxpBeDEARdzICxqWVSibT1VKM
HZESWxglloplB1ZYJB0wDB8jUzovZ9E9nIdz1bEqTqzpV8Cyec0ZLW29SIRHOv06
TtGdaj1NXw807V9gTLMMu1BMC+b9UKi1ghbjKV0JYJWNC1xjzyNBC5htakKpY0jY
BywKG39zl82Ml8KB+0FLeFzXMS9mR1CDiq8Jp/+zVIoJ68CgokMNHSL/yUf07h7R
mjBq5P/jASwbiHbvwqzOXY9BJFAOFCwJwvmAJ061/2KrxFI+k/kh59RqgjlrryTb
NBotxtFwOVU9lDPdtUsnaAIMnJtelbf2gS7xIc2wxU3u9TvR16aBCzfe32b4SPcA
fwAQCpftvepZVfsFECJfLbjHwiTGJeZM4d6yPkJZSfmu5qRv4zNVdF2yIw+pPup5
yZuLQbEaeWRIGROP51kxdQ==
`protect END_PROTECTED
