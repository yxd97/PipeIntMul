`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tj/w4HUJHf91abbr0UW1sO4q9qR587ou0ujmpRQ2VynR5fghKMo1y3U5ahmZELsv
Rjxd6Cdu8IchnMFvMU3T0dpron+Oss9lAgLkY9RfzKEhN0eD5S+Advo4CyW4z5EF
8qvhuEFMJP9BuVGWmBsx/O9LicA8eVOqsu5knQCF1ePeBl2u22CZeWK7/fpE/BkF
Z1iHyhjQb1NR4Qu6S5+nXwHbz8IfLjwPQuDyzzuws8H6YBdq2Po2e8i7RcrAxuoW
stsN133/EXlhbqv9zjHAnANm6Lj+K3ArybVWffOp8awcPYE/NJKfbE1BsP1z6PKg
wahWaF5wdnhGFmu/0ToQ7i1i479QHmPbdVNAfMRbEvwB4LEpxbe3CYdhINln0Yzj
zvDsWevYMm3Lj8n+sn0MfA==
`protect END_PROTECTED
