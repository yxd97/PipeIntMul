`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bycucru9zzlSFxt+GzwhRfgHRJg2uy0238CshnzjdcG5a5rd2stOSTODObZoWyZ6
tIaYCpEgiMLnNhY+rwjYx3XJHQRshh6HGHB+/qibiUU9T49NwAk5oPP0pRT/l0Fp
CZIYWNLdGyESYYcQumWIzi1TqjqecD3jKwupNEsJ5O+DS3qUtteythCKx4KiFDfB
4/sBJQNvHuIiJvuTVmAYnHrg9Z7MMoFKNK3RwjDgNLwIQK0zYTdyG2XVSvZeY6vr
oVYekKYXFFkqWZrutbYns113dMTOsqrgNoTwmB6NgZlQ1dBxTrkxYkXUuZ9wkmfQ
Uu+k1z9SqgIxNchQ8oh7gced1UW86l2W1x2Rid17+W6dcyNvGphHhck+EpksrmC3
6+3O5K9x5KQgbHgL9FzE5YET5nJwyBRxmpvWCIT23n93VIdn5nXQQyGmgH8J7hbm
XlKL1yhWhlpns/2hm5wYBqy2EK1D+URj51kM/wTWRrwH0gauRziOiifamissV74a
`protect END_PROTECTED
