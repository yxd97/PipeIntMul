`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Gzx4izK/37U4vBwE5xtoIbL7Z6TNLUOMfZlCr93xq5tiqRM8OaKlGTDFuyQjbIN
voXEu0evw2zUTa7OS76RsrrtsZiD/9Kf9i+NKdsr9m+Eeot9vB2V9/ItL3WmWQ6K
iqDoy9azKA1J4bNLzZL2bZ+n3OvIkSbQpWn9hd5jHygjbKScagIgE96PbTqCE3t2
vDSmpqaNdOnIESp4ADPr+feJ3HF5Wt/n1IUo2dyNR3apD4jUAW6ZYDqqf5DFpTQD
hYyejrfAaLS0b4jNIQ7NVByA1dpXkAnrI/URxUmlEi1bnnHLTXC8KCt4FWQEbcLM
/KURJeWHqGrftpVBoo7rb4QEg0ShtSso9qrlfA8egEWTV3H6pQ6Ec4CeCkxMz3Li
tzAuiOWLZRXGZ92liXE8FbRc8Jm2F64aPYWA2kNP1ms=
`protect END_PROTECTED
