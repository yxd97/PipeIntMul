`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfWKn6uHt9R19ZPEGNn83g5Sb8KBDa+YGpSgCK0ZsG4NcO27AMCy/0HJ0TlrRRb5
Ye/JApDzi4UH2ADgP749vUtCOnWHfqSsdwArj2sPRbTocQEqPspjWr97cz5lqA0F
54WUm8YUeLIB6fXcZtlluqFkt2NICi54NXBAZEvBcBBGJaFGCl69iTlh8uAOQn5w
24OeVnv4iy03ys5yn1vqLBnwIVYR8Z+v73qY8D8m+Q7O0uCnqi06lEMKkazGeu6z
0Sj5PB+MS21rv9wORwgLIw32fa18ncVDMc/ZHntVIN9VuQOK+rr0caJ/wJtrz7JK
70BsxNDTlyekbwvZAnvyOfWeyxg5h5j6cowgfSrM2rZbf9Z1Qk/UNNLgfMcwFBid
4onDbwRlNRdIJFsXU9g7n5Ht37jYlztqTtiw+1komhVnugf+meWJTYQR9/+Zq9Ou
p8X8kcxj/RJ6fL7UDBXpBrhMk7XAVCUlaoAt36M7He7ZRTFAUA4r2HOlp7exM9ph
tv75KmrZGza8gkzEhYE9SoJI2VE8yyfc4fxWdQEXQos0ARSTOvE3u3JvqFZaIMWc
nnVcyTgQquE1KBedErjPxuYOJ8Gf+5i0T0opvsgq+bFnCkWJSykzLSSXTcNNSdgh
3rx/C6yo09gnJh7JzJJEzHPo4k1F1SaANpTYYqFdSLOzVdSs3mFZIrtT4NMkS44v
mofMuk6Qz8Ezy3sZ76X/qARurtZhuMSItmYda0Ihrd1qphJkmkeLgNqO1pDXl8Uv
zo9O/jFh2t52NTF0ctkHLqflNAIb06AhhFygOZBBrzNVWB7koqL/skCroUrpqdI1
DYZ5Tmj15vcEzusnjV4zSMZQW9Qjmp5SKZuEgku/1Y78tqHJNPOVOSlIzLVDGLeY
aZpTDSfE2AfToccg9akKnaw9r47p576KWQfdzleKhpOyCYKoRyv06b9I621owX3g
emAzkxAvJ83Vv+tKSuBWQw==
`protect END_PROTECTED
