`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OEWCqMlAYuMQxMi+/Q9qAlNF5qbmVvAYPvrbEKl8ya+cqvC8h1Taqx5YLqPviIRf
HnfVG+T1uDjiqkBDaiPcHmHlwmbz4RetnEiLbktF8/Zvpq4opptYf8g0YLczvwDZ
NJo/umqVA30QDTw/LM2yvyRtdxSkNprzvlLUaw2EpzmS/tSpU6AHS387aZa53Fv9
8aZOv19VZ667CIXor1YCIcXMlJ9q1+m5P9ffhHUjoED8AyMuBBmUi+88M6x4IZ7U
XwzlgPDNAX20GCNLCMG+N4GkpK6Z8lC6YGEPGwM66WFuSYHQ43gG+qN30jNW2G+/
cXc2wvTxBgtrXHJNJmJIvd+X4LmdN9fktjkGMIvRawFfYZKyl7fn3d0TRIWMQohW
yfFNOMjf0anuefg7dohP5IhwFY9hh7DjcxePW4IGajFonVoZIVEPNq4nVxhVIKPO
BKCN884zArdBYm5Rpj2eiEhqwXb8H4kU+gg21JXfcjdJwdr5L2mz3fURaSDULvQw
PRXOKTyBh+BILHztedXhSYHX7MFXUVMkrrGtzQVJyhgL42GsFVZ594jiMhDSFX8U
MqWil9ei0rch0oXhQDyoaE5FALrJFB4IxS1eo1/Ee72hD+Wbd9n1aA34TvRIMFNq
OFZcxzZiijzYYXKhxL3svbDUxiGjhbW7mi8RSuh81qvYoFHFqWvmoUDtJGhapADU
FyVoKWNYZocgPcC3q0Rk7F50+7we1yCwGh4S5UEcbltkABPbPJmb8FeGMyVNF3JS
5QlC1m/9IThojt/R/pldXvCcj69au0c/Bj3Cx2AzUr3TK7jgRbxqiHaM9qhYdr54
GwWOcMHunl4ThgIGzuEdniwMo7CKgQ9DKzhTS3F4MwMUQCQTnCjBDR3MjnxodAUg
5fdmnsZVcwMPe/ciSL0UR/Hdz321naohOqadOles+iuN+Y+vjQZiUxRFhpLZhvxz
1AITkJOCwrFhkJXpip3DDiRPOzm8kDF5fvEO7mP24JL6MgXsu/2YIg11EF4tHFNV
LksV+q/pD7oD82Mu/LQdLl77AQIIG+XiRjWsYytj24/nd3i14tsEyuR2AsZx93nN
XdiuhFNuS4X8TrQBBTCiti8EuvnP2lpz9Vc6jfJQ7s99wco0likMbQNwIslDKn+O
Nav69uQoLYw0hR5N+XGzR1JPfi8G8Eouxp5qjWDbIMfC2q2aJ1LOfeIc/dRMIn27
c8QLFhMULjq/MI43ez+lcfHZjCw0Oznb6S1bQK/rRJ2KGgBxv3f/dti1keXVK7XC
m16WfuBRdIOKfi86We+ruJBzHCI7wzfAAdhpx3j4HYlQYNHu6mUHC77Nv1QtiwH3
kJfS/t4dh6ekRUKL6eBC1O1DEgYVGg0CJYDOZuiokBfjOf0ElIAqS0j0V+XVV0bR
g+SfVgpdneoTL1UDVWSGT2trXcdYyyQnJTGK3mffmA2XcB6ShciNMQH7IF3r4a9R
aOXvfpJzihspmeX+QfFV0iEGLxTjoN5gdddqhWaCdRR81idUG/u1EvOx2BU6YL/3
yk9f9wouaUtQet3TiFF6/L63YavWYo+OJHgvmxwv9TnlfWt9kQmBw4wgS19jLJI1
iK9IIu7xOh77tiWztsbtZuOlGzuCr3Q0TSiBIh8k1P2ovIGGfENI+P/A5QicDLS0
wQKd+qeuuA4GJLhxAIqwfvtx60Y61wouUXWl38yfmurfh55S1yRALnPBoiRRogBg
c7HQkipkwh6x/UvBdgvyzTCEBS1/tr6umDEs3J/KN9Duy08F1uXUoPmIjn8f0UYd
+J72yrZ3s713JGp06Jdsqvsw+gwErOCsqU7A7rtERAK59BC1l0Nk2i/I/FEXhMTu
A6s3huXXuRB2z5MwBvY4u3XyC+I1z7Gvyabeb3ZVcauZ4OOq7nw4Rghq1AusEDg/
RW2/c5HbgQmnph/5QF0mdEo+b+MDP0FpX5gBhox860Zgaz66uZ2j5JBvKYQIpWwv
2AGZfHfxfaY23rKbMdoZioFj4Z26EGN4pkWhckSO1hXn7VHZheailtaXDuTi5ecr
L0lQshpYw1w8zxOJiYEs3L9E+0hW2uTK7KaLuqhLOnObqpVInIeTDoXrl+7F3mKo
gCrgB0cvggze85vC0viiFS6urWCM10dbsUnrMcGzK4s+bRjFwbQez8E0B6lrTCYd
xaBYpVtBiB7PROFN0BBUdY/pX9muAwyaH9TCINi7hnybDeBcYirNHXDl7cPLEghq
e4JrsxSUdmsMDoG2hWQ7BpsIlqu5vnbNdSiUkzrD7GQ=
`protect END_PROTECTED
