`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FveflXyV2faMvuxm4Mqedl8sCMY5pIdoJTam7hdmm2mhRJlBg43vRxd3X3JJIIdP
nGNNBj4YaxNUwYrTgp8+OCKiLDwOAkliLHUQEf9pJIkGm5nmEy3F7Pqxru97tIKx
EFMrZd9ZAeql2rRXz5FGk9BeASOZeS9Apo2mEO4hLgXGBd3I7xkDMOWhkVLI7ZNH
Td35O0RvmwPntH9epdo8H4GC4P8ccJ4BEj6J2Y6AA+gpcpgtYaf4GwzTc9BFvJOp
ITUqdU/E7L4bYQz1wUV/Jqq4qTbNYQMsFsaPjtgrtntlYO1RPIMJNOY4ZFj2Yv5y
dk2jgsRIPXohT+8HNYOLVbO/goWRVmQjdbPc6H78idXUpBh6y68AZ88kg35tV3L+
xrNHjO06kun9n2eQiBKYx5XceirLsolLT7iOlMWpOyjqTpDSBC/DCeSk5lHa7X7F
t0oTQF8Vc9VSliBXm8nhrqdQ7W6TexTmdEol56Q9JUT3VH8xA6LNjPbG5KCKUnWe
rKSDoxjgLyw8w/SZ0vgIQRj4ATYcmL/HACwLiCfddXUuEzlQXwKFw7ZjiyHCqQHc
adSbAunbKwYzI9c/sJ3BFP1gauuDK2RaZC8ey314xhV5a3kpYi5kq/qddUanK2Xj
BRGnGeYa5QSJOHIUbd1qwMmut11J3ERyX3Sn2hhTjPsZpV+Hi9C0T3SjiuYC9LEp
fQvNtTi3qCO0dik6IlhvZmqu93p8Etmxi5Ladp4QHQZjTxKDGwgyrYfH1krsqSye
eEAFqI5+gksVbyUHnx9x+q3L+rXdWVXSKzo+Svhcbag4zkrHF4Vy5aFKycp6zysi
`protect END_PROTECTED
