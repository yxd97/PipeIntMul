`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYzupu1aAYq3VouKf98XPgv28lAbHU44Ou4BLYFsEhvh7lZkk/1OTbA08ax0LGK0
1CsSKIbrlRBueXmI5E0VIuwW0b6ZTfjR5euD634Vz8cgfjownTESwRYWf56AG87x
4pP7pHRnfaONbNs3QeErEmDKPq9TjltVqo2wpZrPU+j9O5ixh3weVtQuMyDcHACg
ng0+8I7FrfWCzVozw5uUrTP4FjLD37keTM0rj0fmkrUmzWIc4TxTubEetDjTx6ZM
C/x0FUugHYQK/qNPy0f6aiHzha2y3SZmoEprAP2dvQPQqD98/faREzmIzec4+iCO
vxjZIN6ngPS2kjLuuUtD9A==
`protect END_PROTECTED
