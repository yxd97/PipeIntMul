`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VItZObbBvNcV2q4RLKtGG1HtphuVv65Hpvi+yYKPo3YJp1OkCDJL5FR6wxnYOzHa
icEOAmTB+B8xuxJsuC3CBX4vBs3+vCo1scARgMfPi1WrYy6jX3gqGI3lZinIRRyF
j8gTsZfGMT3/RxgL3t0twtnpLPh6ag5fkI5a4MY/6wiuZxP1o/6jBo8S8Ie9f8mj
DNzK8WM1whnI4cKK19lyDHUtr+YAs4fjgeZvBCOksZiTcZzTU8RucsWLbXFlCxc5
ClOJnshPpwFzCp0G9blMuB0NVMIue/VNxU4BicNitUdKeZ4Fdoi4o9RuvValf8aU
6+LeSzTjYkdYG1NZr0FoUIgwqRVzAac16u9Zerlx76ws8XfINZB+tqgn322Rs6FI
IM6nqxBE4Kc72ggM/3H5aaZ+2kL5Kz1WyQHIMg6poB/e+PZUpKuNZ1gNiXi8lhd6
D8I249AxNDnbH9knNqfLQUpecvFXQOJToOb1X6Xle5SwDYs+aLp9fk/lduGvmRBF
DDNZvKWYguFMsuvadagDZ7ttG6zRZ47a09991WG3XW5Q2M2sUwMjzpiPbCRr0hDL
i9cjH083tDGCQ9BbPI5EtUnYYpWILhbU1Y72Kh7Qv2qNt6aMDKxRorlGOI+/grXq
K73rmnBEolB6zcMuIR7M1G6e8Jr0sajTQ3nJGMMWuhm8N0c9rulBzt0NhiKAhbn4
Fn9vBdyiqADNMQNAhXkn9W4qvJ1wNHuKNQdrawfTePU3P9w2it/PwKG3zovfuv8v
ZitvYAnwmUL+7fHlx58Y5k5md3ubB75yyAT7Ao7jUWKZJpQhfdZr2nB2Bv+qN6Wi
XB88v38atdTmpNBDul4dhd2KV8vTdTGzMSyWDvyN9EwyyWb/n4bnAZUqBSwtH9fY
Owyp0bcxORAT3zFemWyI878J5axcBg0yvKNqxCR3DbjPgN/Gq1ZV96tzHo96HyEP
F/8QbWHVAwN9JkvG0NJWjpxxtzwiTAJyl773vI+d3Ec=
`protect END_PROTECTED
