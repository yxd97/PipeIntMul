`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dWXW1odxmfNhkoe+q45zrkuU30lpaeQcTiVR21UAmn36bUUduJ4h/xjsmecU/Tvl
Cwdk3Ab0mu9qd6P5FenQnsl9NZCtfxDWTXzjJqkTXXIC6+WzW6i3Atrfw2g0z8kW
pbThQW3xHExktjfaIEZZXPGQkUcVS5yXMUzNIcry5JG3CQl8tufNNgw8M+PO6x71
RdwvchX3bIv0jRKz2rrJKB7kcKjO4U+ysJg0Viotw0+/5ab6f1YebkC4qV5R3TQP
kP6iqt4P5v1Ew8pnIiMzyN3vyQAXLcueobxHSveHiR4v574MkXkh5i9N1OcVRenD
oE9+HM8MCFMACiRki54Gmw==
`protect END_PROTECTED
