`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qrwxdSvs1ZvqttvFEvpRIMccoyVy53dQtWisUo2kEIDStrqqowXm0JJbeWN/Jm2
GisobUMjBH+n2iGPmv06/rnutEsbVxGb51vEhuQzHMOFq3m5jvxNqITLIMBGcjuT
O97XbibSoFVO3rYQlvWiFsBDnJLVYXlXer0JnwsmMc4GIUTNMiT6iwjKOLiNCvFy
QAARWyUi4E4ZporD/A5EA9lU2N8Yu+a92wheUrpirmoUZ7FWp4J48k+j0YhYRe44
+WutKx5JXiOZkf03oPsq5eJwDkgiJh2aXwDroGbzJ/MoNC/ofrJYyXz91ZeVoKQF
khdHYXMofnnv8qYDmu5YRA0SQkbEjapDgFI4/XDWBihg6P+ZcNR4gXGVeIQ2J3wk
wxNWwMBhzAXE3rJYC5tutLPGVBB7h8a8uYIEmPgugriiuiVJkug+xWtcF3JpbWEw
etiXNhQLVmd98s8nhZRlC1aUESFXz3RFBw24CxWCPtMSiM+UKgBiDsDE/mbPzcDU
oWI8FdE2XwORej3qtHtBAwffkfjo/8NXePWBaRzqTuamBgNXBBkEdPfuNjlazqH8
nOMWtspYQXKec64rj3zMMqjSN8RspMo+vktmNB1OR+2F0so3iiHxSSCsYZ0reTmi
tlAr+YXjZ3DHAwe/kstJgSQ53X/h/C78FDprAfV/l3UJ9sHcJodZX2/W+X/u1NB+
G0oFRUYy4eg5VN+vbdnFqMvYQxichWkEQTo7mZilECWzTAZD6iENePCXZKtbFFqP
03PX9jdEU8pTjsqtUiNNAa7yK5BViCeWUyBnrm+tp/FY89ccPniLX4HhhNSfmJJM
YVeTlgzlMp/Cp/w5kddyww3Fsi5LTA2Q0SoIuvh0dvccmV1cZu6GzhzvgF65eDbq
PnrKBgdy56EepVPFZ6X75P+Z6WmzCmRWy9GggQHDoFMQo4n0q6gjei/sK/fVN/YF
CVe5hTBDLdaGk5QIDCuYTOliE4iTcDjYCDQlj5RF/zZoWqosXWjndSD0rupxKMd0
05DLwWMIQU3nm91ZWXgWQ58RAoLaK2IoluVKGqeoL3jA/Ks1ZUVbqHY68u8wi8YV
42cbxwqd+s+QlgcWopfEWuUQP587NhDyxdSrArY2VZ25knwysub4mMDYLm1AcrP3
aw5+TxnhD6H+/mvrJIyWee2OkueuIAzDFiIHjDBs6MI2frR7STTCRb7Gc2BjuOBh
JNkmzz7+HXk3T6JWG8UPExglX0oIKSrzOE/UQYfOZX2E7rKZs0NvicxpTV6ZS0Pt
kMLKENiaDIve+l3vt+IheYvvp4QqF6A5ExRTesXBUZsRt7c9qeiynkE0akKIUc1f
SqK0djHz9uE/hREkau0BAjzW/D4P7DY75sAxMxsoF4lsJyylSVt+cvYC7dsV1kxh
oQsnbTWALRyEDdTI8XjN+67CQde3HiqL+eNZS9vs4bKw7eETrKjGjbxwuciV21+2
6PdhM62FsPlKa/Hbo6rAnDL4b7/9wyhzw9JVLRDlTxeXbqI3tllXFGGhUqbxn2zm
CyLmueYJSq9B6K52xmloYua3C4NcDeZM2wDHPcFnVJp1LZwrBcNE7tz4DC2YeYPk
kh974HeNlrSJqOiMKoXfS6JCwYP36IXBtqwL/Aoef8IB444SFkCZWtlOIFdTRtwG
xOps8l31j9TE2WJqTdONsqfq6aSv7U4Gl9rykncBAFkLSqUfrhxXObpnKcG/h9vQ
NDD8TDKiNQyZrA8hALGFAZ+B++sXRTIsFemqXYDhcxBJGU+krX8K5FwneMM4BEp7
8Nm6KeCsvyhGeHY1+kU9OYRfpHMtZN8cmreFReOmQBf080nnpeENTR2utZjd15Mc
Xw9+TLchcWSmMqLBviio12jKIoi/zKyAVmVtuLavX8OOHk0cOdq2U84dKQzIYt5m
r6xv73plQe7Mmy00H/9LH9u0ojZ7AYeFtdJPG/k6qcC1iohDQQILcCUdMXsVkloi
2CO3eoLLRHX/LUn4n1Hcf7RPBRXvP7mj4fqMUNPmZpbhSQanFqOQcdhE4r/irhTF
Vs4TNGaahbeQ/3x+BS+Z7RGDj8lllhGyyGRlLYZBgIqC+VriIc2Ds7qskjd1RgfN
e1L2LhQAGYWenzJbxR1h77G/5orCDBFXzs3ROVOE0wwq6jpvFqBYzf5QWYop1pNi
yv3j/3dTbsAnxBj41S8nP/cpNeTVwelpPoqlmQoh+JeNIId5nhDKPcNMc31JS8bx
fpcxysQpI59wbQClPhA/CalVPKo8TabNW239xvONTqcu2ivckdZ0sapC+EehtRYm
Vetjf0U2tIrr9JguQ2co7G5KFp2Krkte2DShzfghxcQlFZh5P6RadWumtVoSTLYx
2N9KOXkf90NpL0p8D/XZ8113H/oy3q7F2KEhZRwC41OS7D8C0aOlmNACvvHz+UZO
jpN+wVRQ8KBfkjogEkunUxdNCLJ0Z+3Db6cmqPcMAzDb3uFdBEnOuKzsOA1JGpYJ
HIahXXxREB1+POUu+zCkP2WBGA7lzo6plXRavsT6LUrjpp4aI7RBfNK5HoQQiPwj
BkLEC6/K87l6rAk/+vjh+Xnr0e/zNoHZ3YVYMPsneMevacLgv2PAImQBOwxntk6z
WKEW4iZ2wdQNAzOVhI6OWzTJiPsMcTmH26Gep8M6Pk53i0mvvQ+bmAhWvaqiEHCN
r3y86mQY9zF5gOEEfhithbD4wULmMwYf1jFpWxxUKRJ4jSyBJDRBs0LXvpZ8KbJI
GYMKDlV2vzrCC8185UsRBQ==
`protect END_PROTECTED
