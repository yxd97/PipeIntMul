`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZAAEYcc6ZDB1ecRqKKqJCMI/5/y3WTlS80t9eGrrWCfYeHPqxMQeRk/9t/NTfg+
+OqoWTD9J0w72bKL7HW/A44wGbqzcDnU3jeNblQhAPDgt2K1RVN/Qa53a6hfqRn4
djBZPoe7s42DJEC6Dx+cGmmnPPi97MCx+nQQvugWxpq4RXmxE1TJyJt1p+4MUHGw
YUdW3Brf8YjvqrH6cwYIrhGYbJUr+37hQtnN9KwQXIfA7NPYUc9CTT65U7T2TFiF
Ibmm7d92NqAWiGLVpFylf4k6fJ2hBGwTCCNjMiH+J2w3IwwBmw0my/dWHQ7F0d24
cG+vHzd6L0kZVvxIXL1yvMDX/xWgyBo2PyMfXLkJI8aevtMl8c7s0LuexqgLWD7u
ayOt0MdInnQ/PHbo5uY/2jNSR7CK/cY5E5/7mIenkoKMSkZsW04hr7TEO6XRPTbj
`protect END_PROTECTED
