`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTVRy1Zrc1wEU8DO+tySehMfydaxur7UipNHa4ejjR+DSxxnv6xenP7Ygh/+CL3j
Unen0DbYpdF5vg1iTntHF0Byt61jmzKu7TtT4BpTeiHjEe5CzczPZbD+qlF2KofB
i1ouMQV1BeCBzYi5bSM5xXmgiJSLwdmpP3UsAiUOxJUWwRdIU0SYTcDPPWbzqwxM
H25lkl/RnqGQER8WXXYn8hAzAmImVc58uygDbkmiKW9R7MT4kPMkHa6RZUylo2lg
R4EpPpZRrsBM7ZgRlbYWyKIw2mAUGReFnFb8k4gokMM04Tlcbq0RAmridjG3vHlg
znVn6YMiJsQeF9N5BNHewepOdXXVR+VVq65aGvbXWSnLJaOdm1jqeDRQZAcC08yj
15tRydZ80gj5CJEiEk9b0i0jDVkiDlKDPPiil9cgPI+h8PK6cp99qzzqbDz0EjMQ
B3PERX8BjN25hsrnnK6tDMsAOOI51RAMtQq+3lJLb7lH2P23PI3ODWQ6ryxCp+Za
wM4PI226JCheLalOpFz4LCIjiLN2oGqCk8Q6JhjGN8aLgSTjXZ9JePY8ZI5yozIK
`protect END_PROTECTED
