`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVlU0Vsw3NlYPNfRF2/z5L1pEqWyF/T/sQNnCBqp8uZcYMGC89q4LUWOFR1uWboe
hpqdeFoMxe07d9wb6RjpM4GWNGvW6t4pU6VTl4E0A+uEXwjCSJ+SgAGQhn4bH9QC
rwrD6JqWcV6ymeQRZagH4PlE2KtgWPuvFG+Ijtnu7r5P6tmd9Sct5lJ1bfdv/gav
wX4ElmeJAVmsPSr5QzE6PmPqoaeNwt5UUoa+/UoeqHhi0GMfQkryqaaCtIP73Bu1
UMAvPjQD8vqmqyB93ymcc7upx6ZmCpYlClYtjUuibRifcGerLcp7uOyxpzE70/jF
xp8o24QYEfpl3F6EivPkRIlToy4dvQ1BN9FO+LuICzggfHPwOMMA/c+pRhdDyDSH
+3tIdK/AKQKhJxKQV0iklOGjOZ0+roZ6pJiEWEaXBdODaDJVEPzLWJcXmFTvGY95
`protect END_PROTECTED
