`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9i+AtT0Ivpaf1ojAVE6ED9Rb5naFiL0zs8LsR6JIIPxbs5thiaH5QpkaCXFD7YuA
4hlH6RAmdwhq9Al1RWUUGHgvn6gUc7kR8wwsyUvkI6O4za+02SMjWjn45EyuRXvj
PqgJ8Ju74phea1KaOxfieURbMv6Ug+NdmpqX/ba6Cz6MihBWJzGCK65Bx2+/xdXz
XQbbQcgHA8Fm7ShX3pjv2Sb5LOaT389uhOUEqbVflbVvXwFpv4YM5WoywQ65wCOM
uObVOXqJa705XzOUTHBt+shU2YTnpLNRun8nT72VQpjnXRSNYPwFHgpFUJhYXfhc
DyDCCsNxed7/a5qx03J9Bh38KrtrfHxBGE61W1jmGCoQEKREP5ik4XJF1S4b7VVt
x3Y+ZdVv6XZQxlX0JBoS9mgWFrU3MhFFKsx6SCiAX2Gfvs/BKfXApGHQ9eAb2L19
28APv6Xrn/IHUzO8ACLvE+pjX4DUa23pQxMBa7sOB2Lo9kO/pCK354Mv0GK4SpEe
zZFvKW/TtvZfSIXy7c1z6dHYMLucYCPjbAvcvtstwif/CuhL+6b/JEVgAib6Unkm
9TFm6OV/sZfZTRKf4Vdv8Sk9zxofUfqNz68DS6qIiVSYRyI+0g3a+sa3hws8QB3u
onDjd7BwWWJRYXV3w12mKkoXRrUIfHG2Zs2QEgdbiTpFoNVXWvwzOS1J6A7HCmNB
bK+qBVY5wu8tStbvu+vp5cQ1XSnm6tjctxomdLc4vsyQ0WUNPcoB3uMzf196yKWP
/cCHQKehBSjJjsZFUh0BA6mSevqz95cEVOUo0nDR3dfMxgymDOjd3rmnURMIUyiO
ZxaSHLnJJ9XcPQl+mMt3yQmNdttXg2accN4dGa32PrFGsmyOnTpZtnjt65k3F+yU
v4pxO5jeMWW7Wv4eVjjqDHi6F8bhuhxxaikRthfb7r+5kolpg04+IE/yqLSZQkNj
TCiEeOZuCb+rJf4lGUxrViAdA3apeuwA39O/S+msk+Dyv88JOlJzFe/cvWVjinGG
EIV3wqig4qri10mBHMvI15KAF8tWVfTOPUTr1jItLcT2B9QYpCmtJtfGmgVM9aLv
PYRi0WvzD4jQL1bcJIx9jom/Z7BlV7y+X2idHot9KUtd1t3kWx/c1VjDxbcHogGa
aQwnpqwH6KtJmTTRRw/jiN97u+/b7r+3yvui6OVrwzThlecZU9aUh53BqKxr6Pm+
R7tt7ho+VhkJyDjqADX3uVguwSAF8Eo4IvyYDaVcAMrnJ6mPUkhEba3JxuYP730g
7KuQ2qtG8pYNX2kmab7unnJrjF23BrvDsGQcCAuVy0z2BzNHYXoETkQ0jT9TGVkW
QpKzLPsqOtBMTweKI+SzXWA2bMzM1jlAnLnQD3nE2n4TvhOAhpMKoMdSbZkrK+y0
HgG6VrEEhyGgpYKtJvPLzHsZ0b6p04mQHUeFQf+47KuLEZkcoqFoH+UK7ozxeIhi
8DhwCtjgph8VQmWKeIekPk+716yRmoK6+mZAvjidxgkacw7YoMWqIO3pOmK5mZxu
Z9zxD6rTOo1UAhonpTDFnfOcdLFV+kFAkh24nhzjY9J+KC7b5mVUdQ28ibNu9KBV
UXMAJuBS9qpO4yAoxQuRwzK4KOGq7bNZF8lmDUBOqB8gMR+tryEEYgiv9A1ddBwy
IjPo8p1lNgHkJMGvfL4yKBW7kmHIO5VdqfV/UF4G91kzzkSvFnJkAE8BEYbtwEoD
SOCOOUK7+LUPA14vLUhvRobudUU8GU96UQ/TVLC+WdAPBXP+Shf59j2pyeLYZz5x
DjFuDgqbsAXKcJzcK+vXR+jBXrMj7Vyy+x2AdJ78RMI/kEyVOxSDHvHxnoBIOoX8
ihhnChvpdQ/L2Vz9R8t6zmY7tF7+fIfxjB9064cwvq5JnwNrViam3GtthONBsUJD
iTVj1KQ4F4HbvgR3wBdyeaP86UX+Gf2960W2x+nn61z8M/um3jbpwl6BJNUxAufk
TFvmXcxZo8hPT/DnE6dy6w16dDoiq7x1QP9k075tMLwbldfxrmFlUtcNBQsJoezj
HjOgoWDQZnMjajYXZAFBVnJaeXSMuiLbkq8graKnZb1k8ywbkU/Ur0cDh0KVCkB8
uZQM6s5/amsqbRfAYqmFL5q09NigKNnNi890eZkAOvt11We4aQ8FBG2PoWvTJtMu
bKIXJ1ZGP7TeCBuUWNFNyFTMW687PLvhf0ETFi/8KMIs+TDD6JIZ9hmPe9pTFLbm
Nc+pkbg708jxPSx0IG3E2fQ/77Ne6jjsDxXAFKIezKQaMmCCDPOAIMQvFep/761j
xn5GdkKlr9oN7t22Ny1eyX8IicPKefSw2fpzbqvYiUcBQkhkjSLcY7BORxq3Nukl
xXBgBKN+REvYNRndKOB/2kP4JPmHUYTOSNq6w/LewaNpdBlnroXQOuAkkjnuJ77h
XQhPpnP+FALohkgqjEZ0qwW2WQZ8Sq8Y4i+3tLM78TkN+fvkWAOlY8hXMV5KCCMt
haI2PZ0NKsDMjH5gisZ2cQCWAuKSrBfvAqm81zlOUo9CyYfG4jnD4GvcG9zM1BY6
nWIP5C0ZRUx3JPlduozoS+Ke3X8PneeUpGrwimHhOzEE0z4+qdVFwXB/edCQaML3
rmPwEn1sGBAmGncFLt2sY7cCk6o9FHylkwiAKULgznUQvmdD9k1GLrQoRd5xVR4J
QCjgxQezY6lY0B/BI8Aa1ubq4OeXAtfUikusRBUjSKrTXFBhAiN4WLGEpHvIv/qx
jxrDFHaI7JrWUYUBC5TBOLsZWdMRx2dSq6kKUXBemxGM+EhJk4REMdaIDrIwxtfu
0svxo4XtiLXog/8K+gqO7Eb2Ia1cTJUEhXHiaPwXjzKiTNjGOJViinpDm7Mntdjz
MSWM0Bj77leV1bv8Z1X4afo9rusywo6C7YO0HkM5S2lUDRSCgpz0vaYVP+of+ars
tqY7Z5cW1eytIbBbe1fRARuI7L/MHXNIMCHLcZYmBYyTsqP551njoFiY0K3s11QC
nQhOlOv5m33igm/4iydBJI1T+gfzv54YXXFGxxaOYg5b5md70Cdcn9NcQg5Vv5sI
Ylxlsa5PHWce+4xV7W/dUUoyGQ73u7hrqGIHRzGOR07XpmvxP2WZB0yhQXzlo1hk
Eo8ly/7AtX1M8QctSuKLIchFR25EScUUkPiS2Asmf7LIBVTyZQeWrzslecGvLVUR
U01A/OS8Fe/B0TsLTqlaaasKK19U+/tY8kEM8uIhQJ1v5Td/xEPL7Yw6yGhref79
oqieY/5NzklG1SjIAWpWGyBDXva87y6/A4fwd+YYbP2LTVTuzk9a8R34H+UDSvqf
w1QmEbwy3xqPyotVf0JseUra2Lbp8qr1Vybcy/0B0gh6bfVbluWuSHotfwe3MZ8J
J8MUiKEZOOCYkYTxT4iKXT2EuLPSKdZUSsB/o0cxuE2+Wh996qURBOLMiOFE2pyl
m+Egouq25zgOgkvqFUohZDjm3uzxURn08uE1SzX5AKkuQ6hS3WuHzexZu941NpV5
msETblgepATXkeZA8O9HoZOm9UaeoWqY6+h5oRXshuyYOJ+4o1IUbL8POPV8+5um
jraNkIgv7u0CeA5CDFH8e83qOsLKCdY7U5O+1TNOpTn16ab8wJ2oyEkdLuoGs0L4
1qNXaaeFE6BF0vTm3zx8GrKq6Ggkwfeg6ZtPHSHSJQS4XaW5pDAclKUs+RLxAN7M
E5FTXE1YY9GRHYMLW0byh6qwa0uQ7H1kvKYd8DNnkUkngDZMFzSntCNkAj5kOX7O
zszl8ksOnCfihEG6bUZrr5N3oD5z3g+ZRmn0iyKEZqfLjAU5xIsQYc6UKL/UNpwi
Uws/xIitqtG6fD/th2wNmDixkzjCa2jXKjO22DwZN1HmXCrXyJazvHXxOH0iQOaz
VGjIB9BvVciirCQAeqOR9pewqplUPgPPB/Gsvb/dAiMy6J9dR4NnbiQPwmgQPWcx
R5Ba5L/v6WPhPNVtKxmCbwLbiuZsKDme04V65j0JpxpGJabdFMt0+3h2reYopiVF
qV1IthlOY9joFD5YxIjYFV4ZGho7Y/SJlMXf/49EmwQY7xgo9NidwJcbDZL5JXnY
5uOARNQq8qsvsE+pD1kfsF89o35Agqd4Ylj8yjPJiM8L5341goBORtGISbg90t/p
8Mxs6JpVYCNoOT/teMbppkX2bL4LOCK6JYrW3uJiGqcXqlq0r5nEVskgGYD91HZg
QEwZFSu5N0HjKYpCKLu2bVB+QPw5gIOJ2pWqWkK+6C7rH+wnHtn0uNc2Mg2XLTbG
e8JRrp4rRKVYi70xduRQXnWoGsN4O9YkC9uvrSCGvo088zJ/Iyjy8nuYxHiQ0y9e
ZAgvQTpN1fdhC3D83pPvZfSvdIdJUy5MYGBs3QsIeuSgZj/t7SnvwRAJJLPk2e26
Pg0SBtPxg6sKA9W/jNl+A+RwCyU6ylkZUmg7te2kZKMRmk79ovGBIyIZ4y9SlmwA
nvYbhpOAMAT54qXQoYftu0+e9TJTjdnnyhOl0n2EYeU8STjUvakdjTCeOdHOq/qQ
/ilsSDBF+4QQdnEdSYxoredOO6pT/pUhtCimlWRj+1eAQJHkoFFmRAIJkXCsSS23
7yeS3+wA4TdLJrD6JcsmTyHRLmfUO1ZD3Ukc9rqya3Yri9RBOitS3nA4tgc7xlhR
h0c2xlmMC1dYUKHO9TBx7N7mR1zMmSg9HQrn9jdTBwOtfAJI5Senn1usXStYtAcT
zbPYUP1wr6W/Z9+Qjanv/bnJE6HVtRcnwQAtcfYwTkpUk0SDW/yC1qerBQ8yalhv
0HmNXh7a9EY5A0KJ4A1ZDVVbEKQh53Bku8qrCdU0MAWH0QeGO8Xu459SX68dD8Wx
BmzODL+E/HQJLoR3qEeQqIgYOA+OZFXn+y6YZedkhufbbnJSAK1GcG681E8APf0a
rqFkddUKYTJnkQ3JLNNcD8t6z7rYUCahX5eoRZgXms3EpKzuYobkA9BNQOF9ribl
C6rT0je1NJfaDPfidbl4H9Mc/UTXVQsYc8QuNTxdKqLBpbLlI6G8r+TCfpgGVLui
afiDc3A53ABadtT3S9CcxCzRAGM9BHuLFwkEGTJkfGSgCL4V0940tByBqTJr/WIk
9AXQ1P3wwxrrFlmz5JnkDRoTg6cZ9GNjHGj+nhFbGwdnKOnxEgDRVdPQpFoDK2gJ
frOfcHKbwWxIjF0CyoJBBvVBKrq0J5Sb0EF5c18nqz7X0dJyM0nMU1cmEcpiuZg5
S0+s9kV1CsgW4T/L7TDOoDq6zPeo12Oaf6B+5P7R/7D+3heh8nDL2TASiGL4FZAR
ztJ3CP+qDJbH3uHm3G5I6cXFc8Qz+3W2JwR/tI190+30t0lYu+gGL3dij3M7uUIC
v59KybM89wExUHZZ3o4V9VCpCTQoEupLP5ijR4NvYpiZaPG9NhpPthojXCDi+QwD
M7QQmOknM/R6na28YruCXevEVzOUTnskvmQk82id9SiF9zmw38BwlnbE1J2bugHq
OAwUph8W4cYpGwXaxkI+7p2Nu14EkJxCXEa8A2oesXf2Cz8zOsdX1lYr1y4cdwUq
Hj5rfHpV6JXT9iHvOna2D1h+nrOzFwN46HvS3GxaTM436T7G/s07eyS+b0uvogJj
ZNSuLFoQNoCLY1HbvtgLqdLNO4an+9H40WovxGjnE6OWShViZbTLMb0QQDGXBLx0
vDC4qJnBIVOiUIYkMDLJUQnZ0EIPwIWsUsYEp+PsgwLWInN0HSsJeSzfIBsqBGxu
FQ4KXUmLmljBIqVifDHeBoMl0XnRAafq0bIcMs8e/VrE1LGmcT/WtwCmw0mkKltF
IuwStKhmCiTpSOrLsQZ5zn/Y9dAwYBSn/I2dWwgb2ocTrS9p0lUFR9yAryoAfNPo
ra4y9jlFIBPAbt1hBzdykA4t/3MeMB28EujQKZFWuPji1CBmUh7nibn9s6ygh6O2
g3oFI+1IhBE9oG/M04XhXim+twDGl0Jt2zMNKDuwCeHaVPXGgGK5qon1NHI+h43i
OjFeqB+L9EC+ajVABBC3qtLdcmF4cx/bsgl/1/vx2Njy9ZgIT3dt7g5eT8+rRvXk
UrdYoSQXVUVkKsubeE/1F60B2kIb8Yh4ynIT+hZpDokGgqPCJrPlTX4KHBM5E85J
IBB1GH+UM01gF2YQBslkrVvQBPbzrom/wOD1UCs32+5ciiG8xT0X8BZeQRWSuF+z
zCxJ08G+Nat5vikAEFgtrvwS7SStGPlNOnvJW2U1EUBZOyKaL1tS8Arh7H+JgcS5
cCD8uAAch/N6eXByRVrmhgO8T/rWOuCxdatJBFrZuwg4VzD7rX5P9A6KlbyeoXOV
fng/XYhqN1EN0A3HayRJVraGdBznGG06Tix83bPXEXfsmerHlIe+nPprQbDGJwQ+
PNEZObCCaFAGdV39JSUEoyzyXC4uft3Lqikny5ReucxB2B07Dm/hfQ6ID+NZRyJG
GVIDWs9guhjNn+nqW4Gz5s3NgjYYP2jqjeagsoBo8ttNOpmexPIixNVrfK0Ut24C
VtGGM1wJeZv1jfbJ189JZGtUhkmWkBMx22RL+EYvw1jVTMBlqQZJzTVpjHcBJPtF
j42dfYsTpHfTbrtz5R91Pa62RgcA+5wYeB7qehWPdfir7hFOoCPdxcQD7bZrpY5i
SaxHO0kLRIBVq07Q9d1GsDJpLiopdy+y3hPXjAO8gvXbyE0RKrZl7TkPZ1m9/1F8
z3SeVIU3UNmO35U//c4NJdk3KmW0y6ru3sSOvy+6zIOLCSBoDqRhTr0XvrICWYVW
gG1fkrHD5HYhUiQsKnfdM1ERtZ7gRoHoPk3N02tbEv4AX2oFXuGxk7UcdSCQr13b
DO5jrLX4i+yKimtoJtEDXDjI7mLG4LIM2GP70pmpS0JoEIbfTkKFw4gnfyiSRVD7
US4OszrR8eFRSllbHCX0dyGf6bq+hcCVxg0Lk9gagDLnS9izAFoCIiOVFLsfErEP
iRFbpfYKv0YZZ164EBM+VlyvxHjpW3UeksMKJAY44uM10IjPyqhVLOqecnzBB9Wv
WuoXYGsORiPbyNE11dBFV2LoTXf8iqXxBQ+NMH0PJP3OE7X5O3ViYhRRCQ6y/oe8
nkh+aj3Lg0i5hf7HvAeybSL//36mBbzGzc0cLY7URAF3Yysf7JbZSxm7DxAOxxNQ
zfntfisvYNHA8qzdq5tn1TBb/VRHt48svnGYqlUQcBVz7WG1lLu8TS+83TcwMYbt
j9L3/ArC/5ptPyiOCissv39KMwk5E74oTgDytvvierDEajHi07riROj7vmEknXK9
z+FPnB+dO4nqVCz9z24h/dVOsYWxmfVe/uppmdAdQnVtKvO3sYJGipp/2TCanBAm
wirbG49sXS0yzx0C6Jf1mN87j3HjQdM7hq4W2HPVLW04fJI81umGVwNDqJbnk6ln
nphGDTxekr4eUS3G3WlxIG3EUw2t3Svr/n6VtQITwHuEhUVZY+DtZuWHSSOyFpzr
LpGYj8yARG03feVO8IrY4fB+oUD3rdDOGMXu9IZ7cl6t4wTH8Le09QzpWkTcRb5r
OlCyglOX2PkzwVlC9n3JKDO73Pc0BcmN3ZoIcn4q51AceLbNAkOKME8W+hRbMGT1
Sa18hMBEiX1q2/eO+S8zIWIZQVdVRa/Gly6jQCNDYjZ8zDfo6srCkCQt5Mrof159
TbCT+o009LxuBfAm/0rJDNwOaUlWGYarXKiGw6ACI9o/8Rd0ZoHnSUcobQnauB3o
JOjinF7gEkOh8NipmF4+z3JQdlblZyt1uC9l7rQ8VSIlmryeqC1f+1eRqafk2mGZ
yJ/7hZ3LWYuHrgcm9D6pmWjwCyeU39X78TC/ebwnd20NxEwpJNNR1UvU7jvleAXo
ZrU1xuhZT4C22w8xl1mPq7c/b6n5bDpGqB0pJ0txMaWLqB0sIP1yM97Ock/yx5lw
0rFW5jP125zkXArh254zH4ImzX/B1TPV01jFNsaqIY9G0584M0hX0mRDJCou0Fmj
jks9TFmcLF2F6C0lPyVPhDN+Pw3rjGzbYrD6LY6Ahnur3SjfGU7lYM4sjWofEekk
PnneslhmFeJ1Tl8wfc6PMSrS0A2ZipLAEVG3xNo0Id0zY1CIhXJKpIQxmYNAirL8
MlMUYyccQhX3agykNw7oEw/4GpCI9QEcA/LrZz/yUI6zHaNNFZhCAfNwYuwy4QYx
L4t/S/bu7gJzgQetMFbX+qp9uKiPboIf+wwQ8Pk8Ygep8ofy/MBLFs67nnvYctgr
E/DN5TLPn9WC6KSkBEZS0MStip+EJ92YwoVaG5wPWFSpeo6glD+5ImsHod4Y0GLr
83jArennVJB3KJdy/pFWh4IQGREP3qCmJsgFsdG2SInZnQxqKI9E5/uwZti+igtS
Lz0QLNCiex5XaQmHK2ZJOoQDw6Z8cbfQqQTc32Ee6jCEpft3kJQrT+Orbc6ZQP33
lbmYlc/AQXkFDLO/p7rg7t2BqhdD8eydmvm9I3/wT0dyYyx898+xvW+iv3y4u+gD
E+llZiT4pf9Up8dnfqerkB0GgfKoyoPUlFCZdjq7aJOtS9vO6D2EXNBylSpOIQhj
RDXuyzr1ZBjv98ZWI/IQTtNXYzGa54mHRLuGSMtK5IRWs/o4kLbyEWzuv1xJDSUT
rnh3hHCiGpnmmEhha3/GEknmSdJHN+OlcO3D92oVke/hQcoH1jDWlEsi/OInOwGr
trooeOcwBn+NR4YJ0lPb6rsl8x3D70GJItviS+pc2tEG0ig/SDl3/47R5zNblydM
kQnh/NZjXq/hiKlz7pnpBqSMcKOOLv3giAAMi9gFFNUBjIr0s1AvjehvKcnc1yuX
oRtZI1yyfMRg8nspeLtiv+TahiqNRTW+OX2ME+epB+3RmjB18tyzfOGp7+2FS521
oFijNDL3Ov1odoc8VO+6RYqd3nUkvytP4OMgyR4uHlfD5GezvCPi5d+1MpFjS1ri
rk2TTtJhjiOp12am80sdDcjez1HwVQC903DX88q9IhfbN6MMohawuM2W9UXzUFLC
pkjAamT5sTzGjCjFopu2s4i5gMrxqhVqyF2eq1D3NCnaX2NmrZy+dE0XR/41qMAc
u1TTDYxDsHLtxumWBEq1pBUqUKa1qjl53GBBrm5j3QcP8BAn9LrlZ15vNdUCAXUl
OfeAf0cEuY00UyT/MVB50+GsmoH3qTVdZC/I6qOhdg+jHujPbWNlstdJkxEbXqgn
xe3Apy0LSJT4fR/0yZdvois2RFFF5YazMmLvmaNJiEhaC7Hi5HxtBf+ggmsUU8PM
DCRyxF4al8BTMlhaajargSsJwZDk2VxOKZoNhgOeuIjqZZikhqz1VDt94XqCM5LB
KPzwMTHY8iK0+03dKyQzRhQHE9euI7hVZk3glVgOGxc/X3uNrVctwno/OhIr2tRQ
v/rmshmTccklUy0oyvCWwHL+1xnaPmwCp3kWPaQ82zHrLHgpkGnF0DE+mFoub+we
cLeaAEQ3Fh44duZ5maGUvVdigcTH4nTFnWAnpX96dNzqSqqCsD5oTsKUN5GlfFgZ
OATeQf0ETZciXIno+HHKZyXgdcgntCQ12UddP271U4EL3bzSrNKx9LVfTjwVYli7
N1WLkpTC/Uo2OqSoK4V40qh73yvmksxzQTW5VrcUvTJeQAdBs/wTvuEPhXNXD6cp
5I3GbE9p/pm0D6xckvsawAr6t/H9VzHebDbiebYjWBD/KyTphdnHw0IqA81jz0wE
W//CSZg0BMlA1Nbqr9y4gqu5Pe+ZrB1XIeGQ4m+8acBciCpawek8XP78GXBi9KOE
8vbeywy5xN79rOEVk61fg5NzZpEzeF2BDzbJf92E7RpJmaikyY8HKwTbNS8EoMgg
TEbsmTpQXViwxHLaGeAQb24i2+Sszqhth9a2tZQDsVJQsWl1YZtdeD7Qin7/aCg1
uBNsfLpioUc3IxeGCSpOOxYhn/zSa+jLeCg9ysidP2WUqvd2xkmZ3kT2os0KWttu
uVBTp29a01tyCkPdAPP+D3d+JaxC97myuGAeA7Y7jwrObfBihAzulHgWS/Cmo5Sq
0pmy6b3lkC93FQnEM3FLoWSPloYwfWjLSXgvWYd0Tba2+H32QUtyTUqE3NnzaWCU
dYNy4+5rnuuUd/D4UIn5l/5B0b1VygY7GjGV+CivxBzlNxeencpSWW00Dt1xD6Cv
TNLGxZ07m/JYHLVAyhhO3FB5h/KjwYdy5cLDM1LB67RjJfJZ6zmBhm5ga2gaYJPK
tdT6Fr9B0nirI+YN0EjxpX6J9eyVi2Kvzl2whp+B9H4xCGOOXI6EWuKWcqoLzvKR
kiwCG4V2xsH5ip00Rw9kIl6UjVwGZVMmBIJtSRS97JVT9y+6SODWYrlMsGBa14x1
kGY1Sygf0ZgMS3uFO277Uz6Uwwd8gdXmAGpiNoNBqG+xGGZ0ORKtukod17Zf9nwq
KTU9MrgBvFmrYKHELxXnkH5o4YyjjYZXKkUGHxMros3eJUc7R3IZFKXJAZsEVm2x
OtfsuXJnAF8sZa4Teg4Vi8MjhqgqA3KrVkavbBMyLhiGWtc7r2KvsTFAde990K2h
ioOx7Y8zCyvAz74ZSc/oVN8rTO6Gtpthnmjn2Hew3lCbYrvD/XEbRKI2celeNnze
kBGQudmJ/lfx6ACb87ZjuawEHGuOt0kJk45tkwnYuxphIYyprjLFD5rcLW2H69Q2
lm90FDE7moUx9UGWcEyIFTIyo27LRpJJNHdTapZP6/9b50LPLTMaXv/79ilrkGTU
PTiYTUAtAlJbWcUbRtP7sRAPhQDcQ1MFxBxanQhhnSMNnGEd/wU7FgKhvtMcUtX8
YwGgv+vi/j7bhub23BRWiQvndt/WGRhWXcDQNBKR/JtF1utcemOHsdeJOOS5FFHL
oQxrSppB1fMkAHh+Ymal8OETeYrRnS+yrFkKILwpyKd81flAJWOUMN3vDt98vVgE
gPO98cMCrmyAfvEJLX7UwYepowNKl94Up7GD0sltpNoEXtF59b/wqIr9pLXR7v/q
bbBPcZHtegv+9oSQkH/kLHUMaAFfWwIWJ89mnfA0jpGYRoCU+EZccavmuQrYi69h
qpz+r9ocgh9r00nS26rexUGmYrbLOwqTsUxIVbR/WVGYZ/YUMpl/rsnZscGGXrFc
fU0sKSCDfS+fEC8y5UZVroD2Q8NsEOo5BluAg+upMPy774T6CR5NZllg2Y6ivPq1
gh7Z3WQ9uvMur6bdwOySl11IPR0l3xMVzH/3RTsj4F8wCBTI+REEHXXad0fI5q7N
A3SVAmsO/LLDiuVSLtCWaB8TesP6rnypUcWExm94D4or3BnjpakBIHjGztz8xpuV
jEzEqXXeXtsXj/EJK2Q8PY9eHHeINm5ne3IOWTWMS50mOzmRtzirMY3qwUsvZ4qS
LA8vk4RngZiir2kvXKUoNavCXSe3lPpqW8WhVR7Nan712Brm9aEUyEBGjFmHH5mr
yFYnN4e/9REK3xjyd+PSXX1mFpnfZtVQv+IODXNJMHqfofeaXDX/4AmMZfeyRFdm
QplECqxyU4u1+YB11R7AFoggN4LI5us6KU/BPE8kn8cXS0aZZDBFT4emxRIfol4O
lCuTanRfJtV68BywMqh3CdQf7HtS9v15hasrihwRaZMWa//wKnXxqwMZWxuuBJY3
x14uTiBXz9PG9Qqwi/y1n5J33KxLcZCDt4WiSJ/TmAXIOzTF7IupLT9R6tl1R6Qm
E8UcWEXcTicZmWneil+xTqDkqFT5Y5H/l58smgc6rS6Iqeg06qGzsLd6JPdqOVo0
ZbcvtE+s90tYzAeDzcdfXZY2DS+py+eVZaAcrLNfSmbOQF/1bPRqBiO/MYFwHjNB
5q75wj7EiJGLNZfSVeO0fKZHc02Mh3LWDC1Gkiy3SIAvQWA0FC4kTml/k6UOaEMI
hDFE4dbvejebXet0CS6F09p3q6pRg9gbTr7ppMXonWZXHYdV1iVmrutq2Ip8vPkC
oCviLI8o7PAdpRHef+9E5GAQo47zpk8N8FZtsWmDjeWdB+H5s6Ba5lL1pt+RxtI6
SCINW9D/XLB+ar68Ark/oeIK2j2BAy6BdbBj/N/PLezfd4YsotYU05kMNot29taL
ryBcHlPMD9JLSIC2hkGMo7vnafKe8gvR+9qUM6tOzxOWlRQAFog7kVUGYpZHPl6d
5IYUfkjVYA1zba3lNz6F9jekggZfzMf94xLC/FugGLqUmUSXPXWy/8c+rHCMEOwC
q4ZTLR2N+nmcqnE/kxCXIm1pGW3+avSHZiifhJjbPCGQHCCFCEcDrr/fTc0GeUoO
Ffo/L7HIyK/0M3TGVbOGI4JwXwdHqBvL/he1hHcNk9VAtElNIz6WnGfxk8tiU/jx
QxlDfjQVPBDCPa7WX0Jfs9/WOpHmSFOfELc3zLEUDfQGxXjX+umC+x4hI8/tpmY6
9+LgH2fzjHJiejLJG/uNxAxR3zj8JtqeQrM1Xm0efmiKuf4urG3LKbNrJaGMgniH
2byktaAYmElcG01YviJfKpoTpJmYpLuvVHAfATM3zwAk9F7yi6d4SEEAZXJ1zKZg
lLo4VVwy7pXfegl8pZBCnifrTugM29fDJb90m8lI/4XMl8ezIi3LHbR0EyGMQafM
aWwnfeDgbd650X4Exqe1xsErDruXfdSQpdTVyZ+jfzXDKVCLzq2n7rF/YC5ZcehH
CTmf5QwTaevFgKN55mlwL1wtXB7nDpWS1ElPmjYTnwBW7m/vpcPpNFGJcWFSg5Mr
ZsADaocx/7Bsv0dFNXP3xdOA+GtQwGsnT+KN1QDOts4/2DgxhVMgYfySM6Dpu1n5
5ReAK4MxA4mRAYrGjqNNNOyRuIqXBA5y4ZUVYToJgEx+AbV162oRYpD/F8C60lcQ
W/lXnI+NEHHSUfJlz++lxPjFUptPVxLQKHKhEk2b7MsrDk7RSjcRwMShaKCFzMo6
FITmOrM2Zo9bn9i0rySQ1dHXugaGDzRT3nWENeUrPIvplH9wJTfRshYyzGiKSbKi
T/nZvnMLnNLo1HRrbL27vcvkNnqBkQjlmavS/ZS9+VNhw0J9BoPmxCK0bFFDXFYy
5o9s5IxS9WuLrdIWzgtcKOa3sDnS8IuaMW6+IqmsP/qMhzmpAtZiQxjnvD9EhyIX
JVcQaAKvvATeJubMNfoo6cKvaosSueZcQF6aJfqJvBqwdPq/6fU/0icVHFdvO3UZ
m26BGk/4mIPJO5UdlajB5BfEY0cp03jrlNXzO0g4EO5ftnJLS/lF4t7VtpJBjObR
DZq5afHocBt6iqoxV2dLCQPZiIEnwUZYjQjrgZHexcYXXS2QQVg+7OfPylQ40iEG
t8h7Wvz3sjbZxFaW/Y9zY+6Klr7m7jLz8pXYHcqVyyVfYmbrTfjqRV13Ldce1l+z
LmhlpEl5xrp8BCaDp7ToXRQCdhld+4zLA2dEXVXJypL884V6CdENjWSf9woJRLgr
genqZ5e6gaNSg3YFR5dRw5Noa8xCw9F6Gcp18DiQRQy8Odo4/0xM4v/d8dFZ5EGg
MLIXYhC2Znp1jAGqbnc9zL+XSt/zIlCsK++fdDTv8QFhWs/9ZtoY03ZLn7wXtCt3
EMLYFNka58c+M5j1gYNidsSHjg6gZ0lFYJPd1mOsUlVERvOCIqf56ej98obSgchO
H+cbjoOFs+Zg3rk7Rzbo1c9rVmK4Rwr+3SAkFMBdSPk3BpM7qFZg59Vhf0UpL8Zf
2Wo8eQnjknVltCQp6KIBw0Fyyb5n1mfqbJwbpCf93tlfDISApe1XXsE0nAYLvrhC
r1EaUbz1rEJzCt2EYHR8vgjkhoaCZe5YxzbWXu1CF1lQ0GouDa5oy09iCZuIjd+H
GOXGZTVZ688nm9WgMLhd493QA9FQdK2dqZknJrAUUO+SpWxspiQOjnePXnMtEgqT
UJ/kz8Gi7gVU/I9TbyMo32Mgyck9bZGHTPa4eCtrerXKIYiKuqU1eQcFb6TFvaNs
Fa2NLTxSOfvmRzMaBp12XfTApEtpOcTmT6DEeB3GytMryxDATv1nURWLMHqLjxPM
osNDgnhfKGHjuyJ/w1QjWsNr6bav67KGT20aKWPYzZhhdNabthOQXgoPnMkXiQTE
4Ps8GytSepF3oQj9N3vngVaJEPXXw4yumKt6KbgIQX6mR+MBogZcf3GijM1Y3gBB
u1ibObh8Q0NVxZOvahQ9G24SlNICVb/eYXHnDKctWOPJ9f/pYDucW3PsurnTdlHl
TiSq5q67Yb4MqYD0aYqugDrQ1NhSzzvosbh5wc55hrrZgPuNemxaif9cQw+tKm9h
o07MEKlwxzvW95OhLCyXvBkd9MaZLHGReffdJD8T7gWhpV4Aq9fZeVz04KIjLChJ
+MC4ArujYvQYm/xTxkgsCyGg1eR51i5cXsPuWqUtpl/8pEvsKobc7WeaG2clgtU4
gAT8pM1oAXI0Vy4cVwDBY1jagv7DEM+yXA5U/GEqZoBbf5Duc8bJZ7AEYwOAD+jS
gVlUkyy9kVmQ+ggCzB4+uw3eAQ7KkAMBCK0he+pNRy94NkKg8ONd3P5rsSBOe4Wa
hbj32g0xtlusAcy5tVv4HDQvrO2wumKFNLqmPP1McVbsbtHq7LyrMPK3wLKl4TS2
k4zmPj1lZjSK++cMlSrNb+rUF+IFwQSGfbMWpRBRZyGNFMk041172rdmd+2wPhOw
wn/dxZ8EySiVzMRWUFI89Yd4o73vIEp9mY/eAZF7xlDye0qTDoSG+aLTImrlVq4a
P8jtLaOBwZx3WsrojASy9VCBGd/VQ33+zNls4JJtOIeIUfhbjBrByjoeznEZJPkT
ydGgyB73Fk7kTMrY2FVGaPMjh6BNsM5DefnmdiDZJgCbxwZrGxNxhePpof0RsikL
8ZgfW5xSrrc5TDMIWADgDiFCLbz4uO+smoSOt8TThkgB814m6DYqQzmnbgzRx+VI
c5HwpKsrP6p6P4/dXFlN9020bWupNq8OBCU/rL+6ShAqYwJZ0w6xyhpa6qIug0bt
0JzXCgTj/cVKRL5x2RqTp7GPWSbLR+VOyMAUuc58XeMy/59OM577hFM6UumgDgOW
q/Zkg5EIe25G6qHBKau6DPlRU48UL5OyVvDub1DjqbR/bOjhvSQXRzU0gX3XJVmN
8nJ211Zz9N9LkyC07AM+3QehMwEVWihTC8+xHzZL4l/RfaEdQud6gAsxG46ZUKHd
u/4b0VqZJW++dD2pZ7F6wp88dDJI6GyL+BAnRwnh0vGwbsiSrErcDJPTH3t9XFQW
91friDe4KgRGNqyWkeDvc28BScGHRTsmcQSwnBgUNJCE4ysyEIWUst6TR62tj2xz
Tw39tR0XiCbOzcBAVuSe5iJifpALSoAjVR6jgUfzLnUT12WBhNe40hGKlpRSbiNH
d/pIn6i3PtoVlknN6XksPQt3XXahPL3TY4+sPHsH6VZdcyonKLBsxnTnxgJ4STVl
nSW58s8Sbv+QKNttAL2T198cqV2KUZhaJfLmNHwhhaHwYq1Nqsm9xLCdK3lPyT6K
on4oNJT7WJor0Gma0qayKPuy/YADvFCHCWU+WabBGA9bXwJuXpkPCM2sOyPD1FYD
skX7w/NBCHeWL9RFx/UPsVvPGk28OVWo0g4Xa3Do9kFWXtp7Z99PmNMeGthX10Ie
R6l7Kp0QeP/+nQmjOIopCJ1uufOCUdJQACWaj/t2xtbpgTgn5/tDT/uDEp2hwfaU
jgA/YtUvkwr4HCwUHNTkO7IhCTeedTq6dghRbpJ4R3UQkkDmYv3VjWbrfftcEyaf
woajiBgtCtNlYYqMW1okNGvhnkrDSrgFbsPHPK6CL2XGCObPhKcZqxrCRvvUJi3/
xFiLvDWINXTul4adWqmBYeT88jh03LpfINN9AFIpYVzjhcSuMP7JsQ9hTMsnOyst
2vkNRexuHyJ5uNh68tJ3rnPqMz+LpRLcuxcANXTXk6gdwd4Nx0mnP5skdHb9nR9k
tM4NzcL8bZZv+yewLoki2kI1/TDAfiJVnH6IT1FFBjA5LoxOvKE37o4ElL3igzVs
76wREeoH/YgAOPy6eN7aBEweU1u418cxa8nvsk4fIivjUtsVrhl/sILIQm0Pdhlr
0l2R7F6FuLL3hFrV5NtQTQfZa/Ke/YAEhlAojlFn5mOFsE+9vCJ5jJVGRehZrIfk
atNFJViGfjfrVZYiiADA7zCLii/9IddQ8ck964yZC+0EsEbQiqPiHbuJaISKfZrt
65m/Iav7IMIhEl8Y9MruV2MLzxmzNsqzNyqxJ7FS1TBsv7z6b4p3x8CU4I8b0XgY
e82saTRKfmXwEr0ogEGx/YuV7Sy/8dixGv53bUikhyLnfX7+uhtYZ+xW5BnFHoMM
F0S+q54aOENOrISYfGqDP95EdTMjfxqoW4uJRmXheaKWmVUB9oD8Y68APEWHUk6p
bhdxFP0L9DXeL1kuOmHiouA7bntESTWrzv+RvTsqeIMQi+yNA9EhCIoDtiFjSmM5
jjD6JqAW9O4JxozN+zbJDsDFS+RLj54qdXw/e0p1P59ApVKEXAEmhU/O3MIihl9U
6QsH/Sqzba88BxovTxLbRrv3KaMQWCXyolL55z/EYN+Rt27+4Ue6y8AwumS8PdlO
4Me3w4OhGmSbWzHoub3eSVn/d1VmfnNcffkXglftjouJSB0R1P3bpw9u7SB4UwR7
tNE3WQNdEfDZlCGQbmuTB5U4S+mNnu8wsVzK4JVGBz+pq1YcWW/ZzL9956yPT1gf
DEQ8Tqu4GmOASpsKiWCsIyu6TYOQfPuBr+7hM89rz8IKtH4ltFQSDxKuFCfr7GE/
TkAa7W3wW/zhcoPZdSHq25bZeSbLCw338W8xwVJ8x4gR3bDhEGoFkmwSs4ZS0LF/
xzRbqULSVTOrpftGryIBSVPtJEnj3MeBvLTqtCw162jhhbcWxs3dxpBwT3GWDG5Y
bee87JrRO8cV8g23rlXVvJY7fX/pTGoZPjVw/tGtlWVmw0qAKTLFH3DtfHQGkFCN
0H+rRoXr/2Ka9Ah7S3ST4+GWTniqcoALbj/A8HOwDHFbuQ5cRivlf2P5Gfa/8lCk
bfIMNlRLu8etIic6MxNJ1bU4VQNf6qkn+8YI6/6PJXcemYNh0uXBq2yWdzzDhuCF
KO3YQVzBfwiUOJEIbzvY+xUI/lN+gTW5yRglpMVcmLpGsAsKls5pmjhAP6rH1QS2
cJuYF09lzNHrv8E78+kzY330WzcRquTJqqhW3/OTi761N+PNIaxLiNAi9ok4DbdE
ZHduz/53E0GJn1ZQN7RT7hgn+JONycGyqr4KpmX5Xw11WMwWUAvQmAqRHiePbg5C
fqJV0zwLwhO/rJraJBtG77J9VTml4XmLiYPko5y4rFs4gT7+EBBckzTuHUYSF3zh
Mho8Vkv4OSrCvm6bksexCD4JwsWUBazkavl8gSk1xRcfCCMzuGVJaZItchHdB+s/
btV1kaDT3x8+JqYgzTy3dRC+DF2pm6XpSLPVMcxWhQQufrRPVMi/Wuduecx9nJdn
pOhzXou47UrCL5liwHMQq3Qw79nt1mDN82DYMkkB7WGTPUSiT0fSlPltzb7qLSdU
Awze4YPh8PM1wyqDy4miVn9FgAhszhEKwf5INuCkaqIFLMQuh0Cx9TZHPWEnemwl
HhpNuVpJtau5jpvUwxcJN34Vs2l2bpD1ROh/NgY7oX865tPDc1rNhGTIJj4MzMe+
hVN9iPRWVPKxIxzwpo9DaHf2tpZ9EepF5Bi3yyPxh16Bas5RGFZl8WGW9LRMVnwL
R8jvaOMeNWdFkSzjVuyoUBUQag40SxrRULHdpCEqCFjvBe4Q8/7KjLgpFegcNJrj
Ptwl/3xLvkffIMlZiXeJ2+WmROYhTYvcrdbqb6uBx3lbXbAhj0muqzEBJOMGhR0v
VezhLN/mbfb5B/rhyF/b0anhkAxH3YwStuJL63BVG0z15/WBugj5UBQt7d1m2ECK
z4xcMIByr+NMLRaZTuqtMnNMoHau+jid4EjAxkK9XZh8GtFlq5GbUerIQCi5BB7m
DQFvW9Pu+7IR0sHeZQkoAYMAcbhkcYCTMJimVdf+qFRDqZRf5sWIuHGB0HpfAIdA
fDZykkGUVwnlLYRypTsZUEzIDYZuEK4rB/s2cd2aEtKcR3U+NKBuZJBEVynIEDGR
6LUr7QlqhjAqrOeO2K0JN9yaq3jlJ9rOfCWGzSsRCqbIJZJRAS5Hxx2GFbfW+nOS
66Wo2dEqO6GxPIR0L9v+3xhBbr9PayS26sGjmvJJF+pI8vL/6nNQCXSWfoLb+i8/
FcLmHNiurQyFLYT0xr1MH/19QMK+E1w76YXfaWBhGnjqQxgLOaFWx63nIn+dqZTj
qWOWG54Ct2J94i4Ef7BCelU2hxfAxxGAFXVMwr8IotCch4wj+Q04pV7j79Vh+vxn
tqNAYDiFnOzF0MuRO7VNrX1cQc65SlnN/IEf+38gdscET3IiLb391PcfuoM32iKl
WrawfOAujtdpf7RB5IUtNmqArPRSEw2ETrT6WGf/MF8scqQxfs+55vhe/fnoGQP7
PIWGenjd/ywVHp2hIOZrQu91XLGVlfkrP4l35I44HFzJesfx45gFbFXyT8fzTWMp
v5Updi4pN7qSstMDh9fRMIaBXMIxnjKqoAyXyX+2NeHSktdL+24x9O2XBeTzswEw
EBWQ0n4OHQSObkZbkPvZTi0yYJue1FKhFkVD1B4lCzoZHYLUPoiIWNxz0rFmNzoF
JPscWdV8SfZfuJSWIZJlsQt5Oc8oVMVZ5KVTkWJsJeZYCxI+ksfqvCKXzWJPjc2m
dILAEHNAWF/dIp2ZnOughBB47MBQ8YZ7Q75mxCJUehKD8YgZTcuvgzqBdFp8R2J4
Iz702fBdJ71/1JJd9moBUkpShJQY7Fj0mKHYrBZpn66yuBOUw7FkUFVe6rIGhlzp
O4NB6MybYDH2yAlNLwMfwETRYORa8MnYlC5IKgXblmfviERrumNIVBq81trxfwJ+
GYr4ei+C9aVX2aNDOzcXMaP5je0husg3qWwyo6UdQi3fabr55JmtLYZ+vP6TA/EK
ojSKHvj9ggw6SrraLYOAIDSvuIWr/KrL9bGvg7xRBXql1lpE/gynabV4eUY22g5Q
Z0xO5fodbcoxC/8CTs4QrTo7dV/FvUM5MkhgmOkyO93mf6+sh8bg6pPqarEmdvjN
ZuauTKuToaUR2FsclZz+Dn8UW7xyDQeUAmpYTCnLRt0wtwKNyhgMTF85EchUgcoA
EBCA5OUCOVTRS9o4bCbEGjH8rWeQZzy3MbJSNs+dv0Ir7RZzhj0ZKR3yl52vkq4a
HKiEGN95EI+LZ6mV3M7i/bzrmhdWL+CkGA6HYOntwDzpq/FmPC4i/RNWHmcgOvVH
CD9rYSy1nl8xuWkFAG5VtJar19wxi/bJ/YwJ08UBJmh9knrQsO2mYV2U9vIrF6rE
QxoHThSB5z23bAyd97ztvIlZyqhgWCQhQVw4kJO2vDKW6xhz/yc8OKMPtmVIyDvm
pNob7yXnhVFYy3Uotjvsxr64W/vkoFcr3Aw9AnruhOSb2fhWv02YDq39t85Fe/CK
xOIKFLqd/FxOPBP4n6/kw+WwPYCDxXgQt9wFwV6bX6tFY+f/8Ji5K8A2z1PS9A6s
b8EWjncsoDSWdkOBXZr/ypUNAP9/2Vr6lQuIOJy+l4sJeqFEK/Ajb18GrkoeQAHw
6N7/bj8+3EmxwN23Qh+3vDImpTeISWg6ZUimA7jePD9cqlOMAZIBKut94e59BQNR
pSClFH+aC76StSBIEraeq0okmFe8FkuKbMo/y4tGCwDuy3V0C6pPxXryjGyy/3bJ
7/CVIgpTbCB/4tkm7xnTM9hu2m+5PYIzfMHKeG/kcakig/lob6LIiZKQHj1jGaBp
ztdZSYSaWdnR1ugytd/OLSpy4/dtJTZdk60NP2sCAt9iTTFnzOgBrLvJFYydVUFQ
LCV/qCG02TVXNownwxh6VrZjZX7iLuZQGLcW1uisi2Dg4EFLcXJ/1cQPIRTnPEdh
d8H/r1/TXr5dbup8Q9aLAFgvlgmc7eV2+eEU4/HWNAQPd7o4KglDeY6T/ulWhE9p
ePtRiZ26C3s41nTLgKLxaqCtltXl4TiEX0ViBpcgbLIGgIwUFAYXFitmQlljLMnV
tYsj72BeLOskD8YDrExAo+L1CyHWwdsx4nGc18S11t335v3TrDJh4UOMfGO/JIXa
BI99FaYEFgu/7ycAJ6PPXD2OOXFZdd4EbND6h2gqg290Uw25hYzgR92u2tuuVnxw
QoPnCGZsItNazfT5NxIotg+gF0Sv/0UXTM9yROviDIK7DSGYckEyIL7bW1WG/82l
TyYvLgWzNKz0aFkt1tF7OYNPQp6/Ba9ptgG31utD0j9dO5MLUwLIKL/5dcByRCcq
CiGspDPRDUt5vr55oqq+gRS/wU3XUDbiwgTq12MelWWfpmqwv9BzsDJcgyXipBTe
8jhZvcjzVbyD2nuJ4c1BRRkV8EUzfSTjql13hnvCYyIS7PfzhM/1VTiJYa8klp2l
PwB9WqN+6idE3mOJI9TRkl9I1XbEzd/dW0F+7ZUyFFqbIiliw1qfO8oLHD4rR5bs
+N5vvEF0OwOTOyukx7fHMG1EAaAQ35J1qgrcRTRArHm5UOlE0Zuc5ZSabJ05Le1h
VB8kvTbtfzFDGLdF4a3+LyegkeCByyui1idwiHVNV2eMipvidmJXZKWIWKAhFvIV
YbV8Jojz0/0ILOgEvpMla/QHEQWDohstd5m3ULdXoZQeou7RkFYXKL2bWnIRORhE
lUr36WiPJAsR5Hy2rAQv0ZsSPHXS3LTIJEOokoAh3cwMD2zMJ46B5QOTe0PN1Ki/
F+9z+2h+IceIudGqIU2FirXYqw/UVFbKp0bhq8vpRMqycf7YeLcgQTzXe9g/hW68
/GE8QdAJHgcac+p+zq+QpahjsRdzPtsR5mEGPFUlqVt2rDlait3NT61/ewoonps1
qHgTaZo/HFO297HXwdlurCzv1t7xQC0pZTDtyLV9apc5ack4C5yKCaMrr219MUS4
JkuNl79lafKiLm99bcKL6cxDpvrzAYuJmbJMPjUz6aLmg24+GVS9yez+YXuKBH6P
IJuayoqL3iBYhdTA0+NJaZzP+ItJC7oj3HNqs/5TtPgrpOjRapdlk/eLYLT2phmW
u3SXxX5hct1W4Qf+wkGnB4igpKRuVydE5Vlk4k1K42X8tZrei2Htyp65U0MtwPBz
RFO3g8v2o1ZlniS84GRE1y1F1dsjEDUbIJD9gwlVKx8acu9GsDVRZHgU9h3iRZ+S
1rNCsOUfnE6PCYYxvH6vIEq3Lm32jlFFMKL1JO00ACxwP+mtvRbFmMRSM82q86EK
X827i9PodCN32z7xhzH1TbmVjz+XCUBlz5BTtYikg6eajYy2CgXFcZyD61afxzWR
Zu5cLxzzEHoVy8d5N7/d2nn080lhAGgVG9WqQiCXLILP4dNCOg/iv6vKuNdaF6kg
2ojUL0tLN0Fcx9uMYSM/nT0V6Udsb40sMhzcnQx1+11x4Au4viya6Jv686cN5zPI
Ku69gwgQX2kt60W7uUwCymLvAQ2DvsPEA+UAVYLEcqoDFLWiZ3NWDYsND8jfNSfF
BC1tL3uIcoqcFpNaOXrJOBIPByT6EeKYnb4xvfZDDnFv60llpjt4L4MCqENU9jRQ
hw/EWtd5gBzTERAtfxyX3/yT+j46koiDvBHdVxOKqkID3zc+f5xsSUyQjQ/BSVU5
/vNtfy67uBjw9zi4+Fr3VXPfMPzSTLW4jm/c/KltQGIkTtiyHigtRQ1qnZwgV5JN
0qmMbt/MWpvcBxffdbjKzGMfpRHbkKFU4VD6vXu+vjY3bA6r603SmDlSQDRLFdbF
V0Yz8IteWzxWn/8/ns57Ww6lnwnnil459WTJ0TMUFgkLFzRJ3TsKoLi5xqvgfQHr
46nme8Mpa9FCoxBbE/znS92oLkFs08+66Pw4F/XRas+Mq4pDxAb1uDtmvY5QH1Kb
0RoYf5rfTsVbSlalqgO4xgWoAXzQz4/LvLTjzz3NJab37uGU9e/xUAMIaXRr1Rb5
z0zABe/BY6Pls387iN/gHZ50en3Ti/hXOM7iqXGPA4fEi1w+xeATkaJg3VQW+Kiy
PwBqv5v0fv45fofM0doHxHuEFpaMA9jOmtJfZrtMKKYu+805qfagSPOHyzfF193x
vX5DwLl9uLgFf+GOaIW7HYbjw9vnPs1lnvXg6jE1xR15XUlo2nX0tBnDZDIei0Gt
kKQRkF8JQGB/7CAiegdoMgqYl4rbytl+JitsFGZMUbWLZ8ftFS3x10Wgb3PBAU8T
jbn5Oz6mgq7kJWVQDITE4JuT2LQcI1Qtf2DGvxB6WWki7PXu98KjuN2EWMcXGb8l
0vw+kl5ib2z1HA7isA0W7Ct/H1Z2CSTYGhwDhR5WhtsMkaDq8uHsxHbvYrlU6mUh
UzA7DLMzMna0GSacLJOUQL3TAr5l86XVnf1Xi4QhM6avalFdPl4rRo50PCM4dRCE
E99vUxNmdIItPVhlWnevIyx5046fpeB3iOEcim2rBvWI26dL70GZahzVr/+KUCqX
z99f/zTkt1j0G+PqIBYJsArBC1huGrwhFchNro+l/wvildzofpeBS5up30QfHtEx
Uwl/KE9W9PzIaw/08DJHYHdUxZJjGNPPsGa9xCuQuaUzPGxl0dAHHp29vjsxihhy
waHNQT1FFibQWNNuTRu+gh9nws5ZqVXwS+aY0bWKueeEText+iPJbhQ6Vc327ITp
QT3CCdQc4U2dgrLyHDs3V5VhFbxRC+AoYc0sWGzU+ypERighqEPkV74sN9MX61L0
KzDfzT06uRk02JRxVxs8TUd/wmxHa4x3PWhww7zAJebbIR0efWse7Vh+ZKWyKbOO
rFlq86k16mBrmN8L2F5J4xI46QHo4Wy/Qw5bVbBK5DEGTrwEsw77ZbVWjsrE6JFT
wFJosYgpxHADcCOxp8h6gY6naPsagqrEoaYmW1ofkZaeZD6MzW2JXS7NVC2SnkU8
ByVrRZN8oiLYrt5XC4m5b8cD6XMCthuYFtnHzEbeBwj7bLRRwVmol96txJSBn6Ur
4eDLPjqWRYbS1SO8V6VAsVW2ibnMPP9u1dGIGRAh90iw4zMyCpNh8RXNNV2aMR9s
8jukGMwoTfjOiahBJ7SPjlorrY6F9gyqZwB4uBXzB+sSrrTrBJBRGLQh2DaOsqHj
2esELDDRMtpkH0xWjJ5V7fwDa7Ux8ZPkzJHUgBZPcUuycQjsUn90WbAoQ3d9+iD9
jBV9LnZYfJa3NrlKrAXlBCA2H8bwT6f7RjZrY1Kq+u8QEwrgXsptbQiFwQPBpOoT
I2sTzou/xK/DyEEwzubCt8nfBJQOpHkSjXizteij/McQAG8HkgltLUXo9LC6VWbC
GUsXqfyh8fxtBlIei7BGnAC57GvY5cnGR3BvbOawTX/tHuVwqcSw6x/0oA2e1gPq
r58Ekg/6aTeavGWuJAJSaYzdDVhk03VO2IpGmfFZRa5fylExM73Ctfj4HEC8DIN4
FyrMmX4p2J7yIxEahpinktswbBtak42skMmU/mqGAU8C08zMlXN9v8MCiNGrgMrG
JDlVL4L+sxNGi/ifxAT9XPvqHN73CjC3O3tEU+FRlabDtQ9MLsUJIWv6IbwtW18J
W+qpxWWLK7/QMNhcVCQpbkxKHfE1vHpNgUEe4UkgSkH4sYvEuAybtq48o0NO27uV
TsWZkY5KIttlBX8EIEgUTmT9/0GmaDui6puD/+cvCshQpOw+ZoblHYsJvlz6AMau
hlNqZYoPqCvWMwWnccTlndCJ7QCmKVCpqq3TSWDjjRvsLz3c/mFmgFQH46IIcN2S
QXYpuZLQO8M1EtPcdd9EMngclYjdDhc4REwN0MKSj4hYbUMvW0I7phmDGX25o4sX
0EPO16PRAxA2axAn2ou8c8nMBYzfTKJcJ5AKqFgdir4rMGnMsFBmbtZMZ12VG0C6
sOrMUMVaEnz7B+1GVDVF+GOpyUfqKKoQOhvbpHFJ76srwFVhXRY+8zb3dC/cwOvA
n8WtOS9CwQA3I2ZLQaWQqnOpyuBkDSeqD/4bzRxpiOCr8gCqqDsHmM28UOkVDK6z
+hYxIckaHvzUfZscokI9goX27SPLTf5VrLA9ph0xeBZP25lGx8mjWeHx+zsakzAN
TPUCH1hbZps+qqaWJ7yc9fbRqNs9QvL0dNffPFdE5v7mCko4ZfXn5+NPqGxorgOk
HJ2Z9jjKeJBsBxji818I+aTmkEeqnup1FCOd8OcQZZuCD2zZmcG1n1TLVHly0nUs
BWlznA8fy+k+gljS32KxF8GX4Nfeiw+PkhuQm4SfN5VE8A2mQhMJRLYeKGrV17Vt
sNgX56IcHNlGF1zidqYmfTvQM4qgSTqpPrA/Xd5s2pIfvhEg3guSoQCFT1qRqLcK
oB1LL+pSHxr5IGcOZiVqJpLNRs1bGu5xG30pxr+/oVn/cxGeS3eqFhvLhc2ycypn
lfhXxT9iIiY9X4ah5YIn2xnFy2TjNyheF1N8xDu1V/Nqej9t6bRmCGMhW1UE8rvn
zTCVHHovALCecJlUPKf3DxUeKks0j4ZBvkxlQdogmn4fk4PFKZ9xU+Zi+3iTptzS
pCvOujLa+X22sJrCMgK69ZTOO2wYT6Q92LKoL1sufG7GgzDvx9MXz2TOhMitUV4+
PT97DG+C8OaFLfCUtA0MzPNrU3yBhGqZz9KDWro6yUqXxIXtV5RAucM/rX0VeQhD
naNTIJa1V7dofr+RdsNm+XfUypDx1iRU+mg6s2uILYouml/lx+W7no9c1WTyTcJQ
+cGQmgNaD7pyEhqHZOvVWa/ItHQdaltlFbyVDNgWxHwkohWk+msF6myqyQMm8IWy
pBM/UuEwZBOvbPdGamWd4dCTQ3MsFhZ7pnTHDsjOAB7P8nSgJXnoSujUyBwvImg9
avgjGXXlyvs3lElne6lRM19QkrqBEZ9IVxfjOq5+bENWXIoHi2jh8Hn8LeTqqVrJ
ytIhiEpcMsnV3/3wekg5qZtajRo84r1IwpOia8BsLuELceAEh1uFMVPJqAtZ33CT
zOhfVX/wOsnWwRWEhRPMRv1FdS+gDhJaExO6a5Ede9QpEkPwW6/mDbWK0+1LTyU2
6l9NyvL8QpClprSvGEqWHGIolS2N0bINuJOdR+QQyqizWZO0VyDAt4YBvZpPFjAY
ld0tfJC48wbnQUfYkf47yQg5G2CY3SXr4khu2OrDzI7x4hvz/agKiBgvh31etMde
s/ZRH77HDGyAPrVI72SUe5o5QxXWryg85CVhmFas6gSoUShu9QoTelutnWBbJqMM
1h5hTgdp9UxdGPar/y9F5Wn5kwQlslEk5jYGiBEd4QdTpEDwF6FlSrRUGKTneNrL
KPaCYN5cmaVl8EY/KqxWODgQJ2oa0msYz6PU3SucIuBVJzJY6LtN7Ke179TGg5BA
JGVrVxNMA87quQQ3lZdsbNzlpAMLakCT66DsN7n8IxrajOepwW3JWaNONers9Qj8
dqBtsf3ND97sjS2QdGutMonKxYL5pQ2HgNsiofsRqNuUCe8pu0MkpCnWVJ84agAa
rLirFzK+72UAk2M2wUZKUTaDN/U2Ve4kgLSjGJTdJoyATy0CTYeVVitm7Y7xBzpX
F3iWCeuBcF8HBFiiPzShYll26oh8VPWwAha+HahCm8VNQ0hL13cZbQbq5cuWUN+d
7/g57wf3wFWY75sNGY2a96/XfhxTWtBYyPt/GJyL0piSC/QZpZenYEbNXnjCnDBo
VjzXHiMetTsFxw2k8af3DMsd/8/58RuyzpVQCIIPtSYy0Et0st8FKdmYIeKFd0G9
GUOZ5u8kVcfnmzgCOuOZqJTicj+E+W0jl2V7WLV7lAcIiMpL8mXVmMdnCMt4zqI+
131sQ4aUrYZfSg9tnumYHYAhNyCr1FwJmkpxGAn5Fwnm3rEFVtni0fOEy48A2IJk
vNFFL7/r+NHBzUY4kI6xmo1nFgwuqIxwSKq+exTq3xpuvzi2HeQrg/eh4bmwTPbf
fQw2oGsdGsXsYGb7il9d7ilwY9EyjGPLmX2+AnzEkI9nNzMOeJ1Eqm/FzoiRlMSU
3s9PJEqwAVq0K0v0WzOifIx6FuiaJE0XnbZFEdJpr6zSvu1HVoExMQr8zBd5+RYx
vlpyGlEgmF0IG+KiNVHSF2OHk1cuAFTLCxdRZdhH5uCUnIMD5Bfvzg7bk99tunjd
6YBy0p4+6tmmyLqzjk7Yz/MzaRzUa9ABoHGWXksKNwes6QP/hCOCebcBVLKrJw5j
BAdbyYbC/f0UbOJOOqQ4A58Msk8QaLJXZXfyQBFO12n1CL+jSO51BTc2nJ4Wizf3
x/CCRFNKL8uFhoh1qfxytvSYs7gHiGBqTUfDh7my6G26BttGscazjBuJAloX+1KT
Zaawy4kRbmrVoDzcE4G4oUwPaeRgM9TUmRqzGZL3uXH9KDCCsFJ5tul/hWaQKd2y
xFasd7e/a3/KnO9KVBthIk6kDWfePGfAo+Uprrq5XChEnNQoBbUrOC3CQv+awLqa
q994BJsHboXMOGh2QLlWSaW6Bu2UvF7DFhZSNHci0ScP8hS18hik6MlmmcP+O59z
98R583SKrifjYVfL8YnsLJEOrsyKYYh/jZNR54N0Yt0UyLFQ4hNPhzo38GUDvZ8e
o/znLRa9Hc1NcklrUsFh1Wf1XL0+8hoeQhVMC3UFVor0tRTjgtxqI8PxQE+89Xse
OSR82FV6AvPqeEw7FIf88o2+IpcsBd3PjuEAuO1J8rVlNF4PiZ4mxSdwsHaWgsST
svg9BHARZfuMowX77atuLrt2qw44gZ1X/dHoQbaME3weyT/3tnO2kzRYKwDTXLy6
1oEnDBHii4/PKmtYxBjFDCgHPC4cIhG4rzhunigFt4dJkkyld+HkcwHiPAlVZ1H6
A+dhXPdLKcKG7QP1R7q8iLnSsRBp0L3RjRxfAFuP9Lawm8znv/I2JpNCPBO7vAgJ
sQkNhLbazOaEfaCKy01UPhLl3QH+LX33Cc/A321nPdJyJ+EkTOjl498Su0uHlJXX
1d/72rIehad/sNFKvGGEqNp2PuVtR52sWxvV8B1yGAee9LjrldOIpRF4jfgLlRLy
2a4P1cy0ukNXQhY0av7YfEW2AZnxEiAmAa6PWq2MzE1X8C49WMpUkeQ5rpz+l5uY
O4Kg0P1ySNosrj938Yu/nkGzdumvlhoa9ZRRlxyB+svzLQgkph/fPYXDOXLykvnm
lzziAW509UfOLu1yEWVk/8aWETXdi3DDwqLUO5tu9mRAtFfRCWoFAhtZbz4q0GnU
004qq5X2+WHNyJXk5cnNHFn0PXqU5xkHFaSpLU4iK1CU1CU6dsubqrVou6ZWXmZC
O5SQFmBC2qcfPWFhxXsEYbHSGz+3XscfikIPb6H9dZSUFLu6dddoJwtlmCroYOGO
dnxTWCdxJ3oRe/oIFweFqW57d1KlLAQO451V+OxLfVRnBlGHhy3CutrPl7NLhD+J
fzvDybyuhfGQN0x6Rx/LkAZR7F514aGkv8GlIh7yoRig3gv/tGifxaZyYI76nKEp
BuCcqIrsuL4kr/a/GDuk+SK8C9aVhvKQMXkVIbKcstD4E1EuliNwZc2myLDNJ80H
8JmFTXgRqJYwQezc6K7fnBnU7xOlp0o9in7kjdrfiu6NG5qPhij/LCONvoZ16K1X
1zRw2KIYN7TAGy7dstQOSAdkhSpbxn38XIRstdlVTBrMaX0ZG7s6gAg43xjiR9WG
njy5uC52m7cF7dbZj7hNWWjcFjcU6+RVHqC828pr56m+KT7x0tLk7Jm4PvkfMLB5
wzwYF9sd+W3tEf2XGS/1VMaB2yZjuMnp8DU2KQKmT3bC5z8Wztarqr0drlzd2LvE
5AIiVVdsRYc3u3NBuPe0wEjh3NhtDuqr89FY02eX5czF9zmPepmbDpnU0BcDiCTm
lD7EjDwO9dIkpIZ91uODM2QHD5ImT8tCgIxLAmFzk5UrwbO0QbIUAKYTb+h6MIug
RRXg+Fviytkg8j6lyQ0YU3dHu+ijjQc+6mk2O22Mbbyu1/ZpcA4400U4umXH7ZZ6
4HCaqGb/4Yo3X0VwQqd5JELv/Uwztaaem9+Huic6hO4yn88vGIr6Y/JGwSbh2N4/
2g48UC9j3L1FUdmwpuKccGhp72q6K4cu7o117mi+SpXvasQ3cJBLky8KUK2jAyx+
WN7yfhaF4j1v7vyIsv7vutbRZEENVQhHgBtYNn2Cy5WoHjeOGca0VNkvN0zMTiMg
lrkwxWdhh0aXlOkIUHWZrmNEgCrwW8Ca1OiTlmRjUKJ9RUjshqJXu31aXwZ1956C
pJup6knFrKBFwFaUq116GaGjDHj1MksR9OqoYn5HAMlKPtdHjUj9ho/Qzx3owQ7h
H2j4QXxSRUR1o3j5m+wfHmE2ZYBzEq/7npjevBQkeVL4XPYBOewKliZnhFLAR6Jt
OiLUl0F6mWeCUYzfOhtbFMvZ8B5Z3u30ql0kq7JsTyBW4esB5pVEAIctQZiYSjyG
I+qxN7BBEskC8LyWQXjx5FdOnCs1afFIySvdo/5sZsb8J5vSBknU9LJMD0yqmL8P
cN3Okz9zb74FW5KbbahZ0oo7AJ6LEJUCA57LfwVZO6tBCzdI2pIMJRBYN/Vr5Hp8
owjsD0oHf9YUQeurOYZafekRC6NnDx5uR+02O7lFBxqh9YJrePL+9dGcnG0wDhT/
U8fM16/TT+BBVGqdGDzJArIykc9jXjCDOyykIs3gmBxOzREb/JjdrFkhrla/Y+jR
Q06Y9PqZQQdB9l3Aii+DA2t3yUVqKvsymVQPqeA+J8zFnt0vRGit2YzUPDypqJHy
sOAsFczQGzXL8Cr8gn/Vcv1lrtBtNq6pimy/szsyO44Qg0kHpnuTRkJ0A36hQAAD
aISq5g1dHDYYVsT2lEoCMvUG3hQRMGnJ+qGBCWiNux0FaN4j/W+hryloCCC+N55G
H9llfxX6CvfXFUW/e0f6IkJ1I9WoCjVBlB+VH3lx+MBcaJk0hr1zo44sJUHx/H6O
XC6gA1Wm7xpFXnON1AE/neqYkUHz0VQfANqyryJ6xaFc0i+SZJm/qLx7fHzHqpIs
aDTQmvGzk+TrkHyyetNHyzRTDhNX4hoZLNY4JyvpYYIJfy+71qhGuo0ftUfDhgaB
lGrUd1OXnLxzgVIlTu7u09ADLxDVGnicHz/hVwlkLz1/dd8eI9ifWGgpDuvMx1eZ
b+ETTtonuBblyyK7yRhlAqnjnzXZiIfJCzLLpT0lxT1zlsB+GgTduxwi35RLbUYK
QsDEPo3eYcnpQ5rPxwxlQuqD8lAh6XGxjVy1DqPxATLjTgf43cetslrhRE9dXaIp
Ci46YWr0EVpRDcVvOXa2AsG1GfeRiceZt/rS9kARgqOUaFY4y3DjrFpUBjDOzOtU
fnrHl/oF90VYOz/cNAi+o6AFumRPADdj1Mh9Aat7/l3VHODBGK78meKqq/TmuTUj
6jtZ30Mf86D/8dRBcpiAi1hsMT9biSb7r6f6JsiBAzRR2bNhTTTrUkG020DkccMu
YcZoPjJUCR/foR7zkiW+8LR4IqiR4h8+SR525AyEs2pUTwuClEl640DCdBN64GMQ
BQrllocV4X6RfGvGKWNJnIUTyPc28z81UG9wQ9bTBlLF6MWQh7JVrvnCk7ybLHNq
tVfA8k+AOEyKVdNufQmw4UuerugtEKh9cC9pjac57K7q5R60gHT+K2bVqzQOlaaB
0xCUcnVmDN8ifhtA3W2cMI7kUB0VJbaePOWYqrrLW5t+wUxlUcDANdMp/6NQky3l
WaqLsjZiLW4/8qC9hxpSr/zKXmx0QJS8CVCT39gMXSua+4XF7RZlGrEDdvZq10OG
40dX1zG9izezYQ9DbQkTsk0sRJJpJ2U3x9RAxNAYwF6bYrhnjeiGJ9TXHeyN/UeM
LU00BBULU3WQoJHGBY0fL1/x+ES2H9rPQcfYX+howFCDRhz1ERD01AAs7bZXoQHN
mXU8fa08aHKjlOI8rpcsF0VwY/OUM2hOQVNff0kh2Rvgn4QLFr7nfaEU65zzHMfJ
iWIKb5nNgwxGNruW/P80sV8v9SEnyFe84nHY5ESdtox9ElDum+Oygxj0OMz6rjqy
ZS7Kz3RoXsA83Ws3fXagKRZeg7ZiUl+k/Mr3D6ptXZfpW22tDN5aafVgQwtWCdo7
MPVvFlUFtMa5OVztT5qEBjrxH5uMiLbI+KDfdESLd64nZWn1iXiqnzStBWWRLLyo
JOMArH6ezx3VW6XQ10msa8C5TacFapvcPO0/xEdCuvqthPuwSV4TQ/IYkC32iXca
Nf6A0cB7uMbsCsf3wT5lhDf5PM9IKjjEE8F0xyAitcsSeWdvCTs+WQidrgGCIu8G
3fmyVtSweYzQ+OtO3vX7KBLl2KFydL9JVjgoMeLZpmlY1vpSOYBbKNoTyWw9ZnGw
mKr0wVOQ3iFAjVHfMwIJ9YkSZgzpkyQ6OcuOoBfoXk73hWPh9WWBNgMCeqqXXeU0
yDrEvaqx252kb1ZDR6Y4xTQcAWhPyCkjVPd/WumDrPfwr/UmUr9U93xMM122k9Ri
ebWaG2y+U0N1aUU90gCgzvV6HTZecJC9OdrlaCObSGaMAn+kagTtB0K+rGnQF1ai
apuekkd8GimZqYp7Buo29uCniq/rao5lXZmO3ANMwRXEeqd7oT0tsor9zpnD+Khb
xtVGuhwNMcjl5O/opKVovImH3tYm2b/k3CQn6Ji3gOeNj58E1lc1xm3N7sz7R3Gl
hYqjotbEmGdfY7JQ/bO7aS374UdRo4wdagMRymzKu30Ml9YTZGSTHm8LW8iM3jkd
nRRPK9ULYrqs9ePQwkazmSJpB0Zp15Zg8C6Wwfba1TC6wSTeWoEprHR72AUL01LN
OXNeOe63+xblKm7ONiUbxPDmDX42TSmNuoL/eN9OoJJ+mQMju0a2JXjhMdilFarg
FnJKnMpJGbcQs3x5CUSAvhFerx9nW+5BVZfyap/6rZCKPlPUiJsNxzlGWrfr8TZR
kVCFUGC1eEj6CoUt/RHw6V7fBgIlsZF3s1ie/R78Z6KE9lO8OuAKOaL2/3Fplu4r
9KVUk3Em1GT+t5X3NYsA6BS762NZABPnzr41vz894udHYclKTQ81wTDGBCCjFw6n
yPTYCSP0CR7uHQJAgsiWf8eyVISlsHSo9v7DszHlkUbCVT97Duv4gY/Tvbr88kai
bUSrfTi51QSYsS8GD3NARqrAHZgrnINx07N/JoSYu3U4IQxRvfsdbPaeMjGMnpvK
/f8o6co+FKQMAZYwlq1mwp7nHnDZGHX5s/KYc8yneQsprksOuhnBff4CmeECbfjo
agVcLfnW0Z/KkxKQ7ACVVRsHR4A+/2y0u1dSIkBGZdHnWmfx1n+DAbeJHjgWkw6Z
9sg5uzvNQlqbJhzlAb1+yAdNrLqmHrO/TSOeRtRDqropgL7Tq15vG6ibyyhZ0SA7
AsDS2J+D7gBVzMclyOuJa++Ndp53Jx+3DqmaLScnBsq40KsjqrHH1tsesdiw27NA
BBOOhMRyuRI5bgH7rXt3VjzH5JUyfQRoZ7OjBzs+1OdYCvSI68lPkRys0y4l7dpB
rkFCfd0KwMunYO50A9DBDY5deuVKWASHRUGr4mUBCdAYCjgxGBIgJF17AIs+3K9V
uzbH+C1e9GB9ZAbeUudzYXAjlz0Wye9xGupm+cxeSNe5wVwmIE1z2TbY9rqw0Dly
OAnDfszCyerXSTylQbPhk/1wa9PFq9TUpNwUVQZn/Mh2WNx2hzr8Hz5GdGjeXZhF
aJHaSem93WQ4fZA4qaTzqhtJ2mJva8x6RsOZRnIKCzJtgyNzemM6ksSdkaKAGlMO
xqfMbFr99098GOuDPvKSYdMQRPY/kNWveBIgapNPMCDkAL5Yjt5d9pBy7bHGIo3l
N/NQvNi34rgWiVX+O0J9F/oajTNDTp030pDvlYIvh44IjnEarBVRbmmfiGzAPBNK
j+BrDFRpaJ6VfHL9v3Z+LIff6nvysqzwtJ1IAS+jvGdtEgoGLBzYqBKlWaeg2U0k
ahxbGLFC1OJ73QAZ3vjVu9+YAK5E84i6Nw4VutkNaW+/hlerjdcwXUiLYO2NK6bF
bOmSyIRHVEQWpp4ipvhjNP1+jGHo51a8gdjvp/1jhtBpNIE5dBIQCSDwRMexFP59
MU1XUtgz/kFwAWR8nqPpFFbAqgjQGVs9fiAknyqNCAe/vBM/jeTl7WXREzXts7Re
mbI0VruW0B4tIK3VRUng+00oSixIMXzBTdF/MjME+MgOhl0JbWnMfBywWn2RaP2h
+wKDH7xfWJo0ZGWzOnZX/oC8H5unGJEFGkj44GDrcFIsGnTj/K2EgJvRMRSkfSOu
wUUVaTdOOet3bTeKYq4p2VjbnmcSEi5IdC8XcfO9dOhouHY2gYiBqWkH9u6dYwus
tbj/Ufudm/ZAh0JpjxVaPKNNvCDk7yAzDmj0R8o4Fx2j+gZJidT/6mCh01gMVxNm
6zTxQqKMU3IrnToVOZQmfjHT4bklsRaYaAQFWDZwT6bhIIx6y/JTg6MJBaW+TsSi
4GgsbUUuCOPBaVXD9GRtIQxoZato7e+o+qbKhgWwiTN8Ue4+KTV8bOEqxzudiZUE
f3pqEeKhH5clbGnfiMRastJwVuAKI+w6pGh52ranFxvqwzIOgwXHlleFbn//QBVf
SZrg0D4Cj9i/yCTxNGV8T+mHfrdpW4TlpbkSJKwIGOiSYrGyLeNhHKXp96oXo1ge
NHhBA6K6esU06U+7yHKQ3eGM0sJE1nri2ro4yu86yeBNLERp7aKW/e01c3040NX3
C+DflXAaaBfaouDUS4T1Y5UdGC7s8/YQlOIB9kPI3ETozgr+NF3KNo7wNO8DRT2m
RTFQJlQ8ntjBjCwjYH+3wA6W+OTkJPRSbM4z+EYPFJZQaDVsqSHMQ2h6JJ6opwhp
utsVYDTsxBsJLaFZrpMZZ75NzepJuxHQ6HWKb+lFjKfZ5VI0VZ8lujXnP9ww1DBJ
NQLhypIzOxOTAHHi9T2SoKABPr3QzLt77Kq2WwD0jwWiSgM/eWc9Ix9kX0HB4g35
gVeqkO3B0qh4cXXrjOTCXE6+W7l/s1l0rr+uwL+4ZcC34oPHWFMjLvFK85n0Yf8M
vlHxRZOQgLdEhFbaIeYC/jgVjyKo5GP7CGbBkRXcPv7lkj8HliV1VKKSZGfdyUNR
9SW5Zh33DXJ39yP9bp4oQGzvTelKPfOzP1t6Agx/apNoMIsOwFwpxdB/J6+jDrY3
6cDOU8/CxACWvHDQCq8bmAvWkdYD+Cb3BzuaFBUkdJ82fOL7/2MYWOv1yWG0K4KV
6qJQm9qWkGsPut+HymOvkTBvoyfzdXZjMItFa5mZJ9JiFAqfHLdTFNL7+62c8nAK
mWttyYZ+gnxduxsou2hzVQFnxIBDqcWRU6haTCbchkbRUQBY9v+ghg46fQ97gtfq
iEJGtv3ESVl2NTN7ituLOPdZBTxlIWK4YN9Odm3K5vP43Pc1ORuljcrntV4TDYU9
IReb59b1ec3fh9kshg9NkNcaTVRGZeYequMcJfQd+bea4Szk2gnb4zjM/aIumHFT
eoM6PPPyLMaz8bt3EO6vseE+DAgmLOseuhzcpqOuyuMi0Gy2r7YI5Le25APQPxtH
N/SfIBY7IB5rJJz79kuEa+rk3sgd5cI+nOvoEWEYlYddyUuouba2dy2N60j756Nf
YQWTiTyYecKz+2y5Y1rNGQaV7fdxBi/WQkElFmi8GNRWyNsF2azzNPlyYzOqv34H
LcBJNjTGZREry73I/nHcYX6Ivedr8TNDL7dXM1AFHrUtMF9aEoRkMgj2VZd7ui7m
f/ngkxNsr/hYMOex3mBF19iTF1dfRQ/zT6v54xM+o4JV855ObNx+ft4nHP9dZB/s
tRSSrQ/1xHlBoB3MIB83QnZv4be7EfmCbyTxdA12g4d6rd5v4CdQiczwGsn410ze
hakgD46Ctwf4JmlcogbqGqT/VAKIlI1UkXLjXgW4Xst6I3Axh1Pi6l/SPGrscoXy
AtwGd1t4F1lWYiRALmMC053JfQINcqJCOYt4VqFkvDgXmTDg2O/in/d4SYdwYKAw
aLWBoEFQ1gvkeICRHxLVV2MCRwWc8kf45Nz1deSoaPQBxf2gGPFUQmkBbU+V2ehP
/gS1tf1DThvIwqoBr9duTiNCPXZlZ2hbMhZAFZVP+oN4nHTYVgpBbkmB4sRMAxmP
NKMpgK5cUkDZATipJYYHDjQtIbHTyhcoigh4DK0pkneqYJCMdV1WNOgsC95Z2cel
F7W8s0P+e0HxfhIFigNL91zVnp9NtV+l0jXUGu2kuDbTvUGIy1jmXDwhwR7bIgmg
yvnpvny5fzPfA83E8nIGxyEc3UoBFcXedd0FAge1YWyFSfq+3A4FcRwpWYN0e6RW
Rk9ijt+DH9ly12fedQ3kYJAuqMCCU1rG280N0o+KmgFh+Qbx042PflfS4eRapW7B
q0VM/1hAYQWQkE4Gt2z8qaqHGSDrNFgiNEi0C1ahYglpk2n1rroONOv033fhU5w3
85Q7B5yWovd1jOfR8z1Tz0v6uMGSXUMa+QJnkwaOCEKGHeGSItSiljIjd2bxvhlY
/apLW5tK5d+V33B6LMUefSoQ99CkgNk1rk6PJ/LaB7Y+JQ9qdmSEqUb/QEUUiw73
5xUxWvFUm6rRFEaA+qfrXC40go9dLl7JvWKJWbCessXdG4oSCW70g/nZ4gtyLeAQ
nlm7fHTtdbAGESN/xk3mwiJNmAQ1yPQf4TC2zv0gUWliymM352n234UpmjMDd7Eh
MAdoucoJR6mxcr1MRyvzdDRPI0oURyH2Y35dr2KjjR8tkgNLcihsU8l+i/3ZjxBG
eGSj8J2cmPfX12guUBc7glJ3HH9YLkD8CUeQJ8OHnn5AmE6fDIvIcivLnF5WCdMq
yn5lN50kXWN0YDMNHk9TyHv5BdA/DIKRezzWVlwo5RP5/oWHTIsZsjrxG+Q8/r/N
bcQgmXUh/4Dp1QxgyKSzksAStxibwZ/DMfck2Yyd9X9tiVtomuE6/o0r7d0TT1bo
syAUg/vncEltUb571djJh2jIFsO1jAiikIPflNUpg9AAJkXxnEEr0U+1HJrdD1V1
tArqJ7CWVCLxKNfMD3vF8stIKco0L/X/HVU/TN7KcUG05+ZiFs6bF85651y+ukPf
5Hs/k16J1XGYFErviF3ID8OeN9zUzmzGtbOdVI4W56WzOsGmdQc6Z69lTHDgueaF
Y6dyRpGsL3ZTeHTZ08wDY0TABVULWgZaBMOlbvo0eaVOxkP4Y548JVmyvxsn7Xi6
nSWyi6zqzNtq73i1Ehv2hDF89nlfpPJOLIQ8noCQCVIC7GwjRURMK56yM+2UOJmM
0MRBu1mv1vofY8x7E3LvmWQTkWFQin/3MeWq0+8bab8qK7dVcpd4Gd3J5PbY6ynm
+fQK7TZ1MAeLtePDAezG0djTIPT/bwWk1QnRBw1vWk6vV1xx+ot3vWp6jUTLCBAE
oQAIaH3gQS3X/wLRWnyuiiaQNycS2EhZ7maAXYdw58FRvKRo7km+OliYLm00sIZs
aONiANndrwG61jNr+nf/CmRQj78OOHyXV38LFmDOGjhV+G1mcboFLqG8mApk1jXh
rYOL+ItK1dWn3XEuwRZnvZfEFDL3OnUQi0ikOQkeF8/+N5XEDn8p26WBDGWrFiwf
zDzzi+O1o025N6UP0ywyAhnxRt725mLjp28xXfpYhjFLA7s3/pAWFRNp55r7KBNA
cZf6jBSrCG7mbZoPHDHGYtd1HexVTY72RNg/GSQoUjK/l/6g3IzHVUun+QNaIp1f
l1QmDyHlkvih1hkvjBTs9Mioy05TqihhFxV49E/j/MhY42JbPXS9WFvplgjGQI8J
E2rmAXJNuGaq0FvRsG+mgg29LoCJEVeyYcIIj9a8UxZ/NToSR6EcpixkzTHCaFjL
AMQN4hdqsrVISGGxHshWytR4H2uQUo+BV9lLR7C0YtzAO7QGeZImMca5J11RVSwk
eAo61YbyNm2xZWovOz+GXfRCPr7Ay+jWHr5iny2TMzesaOXOawZnkXhVk8quIhso
E0XnIWhLalq8ZZmj+BKMBBgXPmKTsl3EUHOoXp/8IWwjgXb6TqCheYJ4atV2aLNS
rLbmtXwUeQAZ5no4UWvvABQMkjJpfEVPqzJ8njIQu1TWDg9gYeyMhmZKFrpd6B+j
xAUpgnGU8kldIdubOFBGQqJMY4Sqq02a97W9Q/sq7gUYwE3FB5+Ewhe2SORrc/1d
GS9jhThkLkZhL8Rw5bQ+8InHiAG3kdo9fSjQLzWHL1lr0ln51s8IntMSOclFhaQd
FSa/IhJ/7uIUTxKT0fxPYTYEyhHekyUbxeh0+hjgJZtChSgDzM5yCxTHxD2Er3lx
7qZp2rNHdlAknxn7b1vG/UdgH2N5Ha8qrUUvlmfAY6AwL88DzGXJuN2Kxfnof9D2
av1nCSorRxH3Q6RBBY16GS8EyIrS9rYhV88x/U8deZNwPyp4EQdEXrAmcwanKwC1
2ZEWLfq3n7mWPMFJUoWNZft4sIypYdbSRH9/gYrV/1DzlE0gAbpD+pFvh+UH/fW4
SZFHTUbAfotC3FNNXcQroCKP2fBzkM0LlFSbxnrjuC/70kNxKxOlqbs8TCyMcGyA
vLRnPSTb+tSbEJYl+0PjuA2bU+s8Jmc0wY1/9hkqno462p08QXKpvC2G82zbEBL4
8zzC2UgNOw10qSdbIhy5jMhq4vtShUo7NUOTerbeEV1bbBMKRQt2TMlCB4nbYglI
aJVWy1tD2YU/czaV4ArvAw3Omm3tVbE9I3dg2nAHzsByUteoVgQFax98675660Jz
MM0sFUbIJsywUxRhiHrQpNWZIL2o3PrEkS/Batl3qgayVnDg48dGI4UIrsRWU4IG
Kxfuwnc7xGEX6F1gho5+SvEh23sCctr7TSNbbB5gd3/ptTBk6wpzT0I+PgK9TjGv
OuDqMWXvZcFwDZKK8kqKc+z/PsgxsEuT+shwvxGqUuscIFylRQ9EO47pLq/QV+fC
Hb8tiNul5ZfmMPy4AA3rn9ame8Xfhnf0EtyQ3i2fjl1Fq7rehMTQDK3Gnlw8KO0y
XZfikOGWO4/RtfRabDp+HMzQ7y6kU9309GnLfj+CIh690itaXyJN1x91Sl2hcgAT
Q+UCGTlfB4pK7UAS3cY8YrLpGAac6uI9DP0PdIPQ4rmSrg3wyaqL0tzDIk5zlzNs
CnNSO8Ju/lH9R9qbx/mhKMhd5U80VYUQ3Vmvl6xU2yx0Ugk2sW4714hHRdxHvN8R
DCBO8Y0RC49HkXfEbzRjXkCf1fztw8uA19WS8dyxVH7Y7zQz8BCKDGGYmswJT0Oo
s6Aeux397JavlAfTym93TtJIp5omO3Vqsx6dtAJVLgNBaRKYhjXzBSO+4kG0izAC
uQ3H1iL74WU7ZCal+0R7xWWWQnRjy8VhDfrIHhVZdiI7rM6vQ9A2acTdlSOxIGRe
+rht1xhXLUwkgA/O+u2ZeU611Hti+oDWvXMJjMpbS9yCYPVofejJ0hPuqUj1Dh56
VR6Gi7Qk5ak0FpocujUT6jv/SImAHF1A6iC81xo56r9tjLy1MC7Ec8z0ABGdXZP6
LRfrdg8kutt0w15j3ImpgrEtHppPaXsUuvMALe05yXHaNeNqbmrGz0+RdQdghem0
fyDQsbx/LvLSr8oBqBZ+SNjEDWpRU9MYEaydK2bY8pFN4FETlIco+i5VtYlT3ZIl
fPko9sNNO7oSv9cnpDAsKuvfiKucCS+8erKCxJMeSX1T8yd4+Xddt/b0ENeq2868
JRyxxW6zQU1wtj/IxpKBxUgC8a4EZ09O91MqUcbsDiQ+SHDxUSgHoV1XDQsVr2g6
mIQ2h86bTZ40NRB7PMEOXHOrMqWFAfjODQUnpQDgYuInVEuCZ8Fb6QJuyyjjj9Fy
13KgDH/XEr9Xp4Wh1QZ/PwaV3e9a4l0Ii8RO7i+sgxHRRoVg1XraWXqh6VClYYam
mgjWg6uNQHG7OAZ4W2MhUImGbpHbuxjnXwBWTxaxLEhdVZjn1ZsHhASM3arNOPyg
waj6sPvUwvutvWblaF9ZBfTqcSviUPEpyKSQhxLYu6q7fr7GYfkiKrk+xAUdFmi2
nyAQxgdt07Nqi43w6aCwP63gH07IbyCE3junvlFTBYVNba9hAYMfPP7rcWn20uy/
H2NSEv2vIhcq0tesjx33lB1Q531P3xKgZSZLOWlhJQisdEhKo1UxN7fpr+JFKu7P
qCZmyG8Nj+fx/BTUuPwzVkJKK6KWvfA+ZQe7vfN4gP7wsaT3Ij0yA3tGJf80ivsu
PQ58JIwROrxwOMjW9QeQQxQ7a06nza03cUpfoe/i0PfWzixcFTtmwG7JaRXu8Wrm
lw57N68lJDLBsY5p9GiRLWJ8Z7NJf+MCxgGD+CHaadkVHnhJPx6ndtwVH2ut5ac/
fypqKmqEwY3mJLvjVq2qTc8l3fUbeDK6uX+X8kIKP1MqFHDmRP0b+SY90D+aTijG
acqrPBWi9U5DXXqKvXg3lPwovWQs4hHeiW5G9kthSHhmeUhZJGXz3033p1gaATnt
iM00xpE3v7/5BH5fz78xUgejZbJmaiAI8KELnN+s+2lh3FaSlPL6/v9jFoTv32Km
FTUw3b9PkzP/p1VgE/2cWzUhMRkj7996tLvXdW1e773XIejKfmiYjtD3bSKbgEM8
hI12UQH55ilsMAf5OtO3cL9VNx9hUeYVQ/6p1Qg5Yr0MM19phEn78SgRTyZgGmmI
3gbF8UN5k+mRaMzhStx/k3T9z3et/kO8DVceDlb7NdNOrOptopVCLLEaRPltad1w
55T6GPqQ2LNrqyGtvYSko8zmtzMXFR1/8q/bBTsfIMoH5zQN8i7mBN4VH3g8EXKw
0HBs5grLG9ZTXHDfPExyVQN9E6Uwu3iV0Qw3K6PS/xRwB8wOig+l390Ajlr1IEon
v3SZr61zLMQqtH6n0SsvI1KAGNosjU0Opxoi7OB6KmIj1V7AIRdpf81sdTudRM3U
+/N8Zz/hyBsF9+TKYqtHpHjO4W8kYB6M2BQBNB+uxAa+nUafp3kIP2TUaxm4XZPJ
MUldvFMs1HoaB2UhEONiH+pD1s9MdeIg+djmV/G9ZGJqIxBSq6NHCR/sdKPAIFfl
YlblpTZVFK0KZ0mCm/dPVHT+0V82ODPBclMSBvXTtgheZfXXfHnIitfEqYauUtP/
t/+2mxFBPC91tNaa4H2XhbPv/1sVIE+pZEquh1NknblVA4eK+2R+bWCZy3fTvPnN
YzQpQPn8f35T4wbvVWdWb/I3B6X6n/gOh82XwD53ZEX9XQGM0POWY52D+EK/oBsa
Fz66dX/JhKXnqJTw6djw2rvmn7c7K2Dqo9vDA79WhZiEtWZpWVSLi1kqYTv6WD4Z
PL7iG4PmqzOhMocUhcjQvdH+B99K8QsswE1N2ocYTmocQZqzOWiRnZ+t32Gn/R4P
DLlBHYqrZ3nWbseTwV/WOv+hy9haWg2ARG+G0Lq9GUDhHWUvKnrYlZJCetZnj4vg
bJF5JzHYWf4FhaUfXhw1rMINf8ySZjaFAc53fuODi1K/6jUBvVxnXTDbyiT8A0Xq
e9dOaN9+esJCtr+NB4CMfB8qhoBw/VYZjriydMXoB+lh6zNue5uy7JTcCsmNWoGE
0+p66ANXMyjHr8ol78UVaZXZvkOwhvGPzUW8YJh6UdLiulHboWHzIwaCVCVkZ3on
MhW6sicjKsuJCM7RvHOrVWQ+dQs4y6cd8Krydr188kEKC93onhX5cIR2n1yua/Oy
hi20OHe9DgoMM2YbR83inE/535Z2gKZb6x8wcl1EyIp9JdVisqAJ1HQVTcutuqr5
WX/EaituT2sGRG9CrJRim80bnrs7H3DbZYwVVXIxbvXBjSkZg67px3K6905YNFy6
oHw2o2amVZTpS2sQohcKv2DMBppx54jd9LzSKXnxMwpFpqBvuRmRHpR8FSNZa3ek
fon79pxPf9Uo5/5wduk+BD7ATzheRsprNFHz+yIzzuxi+rAiv3Z7KSWG9ZhfdxC3
TzqgC0kmpiQcpG1pEnbu+sYKs98dXIIPs5ylZBVJlgX2u2O/cB10q2/zOJLI+q60
9ctzWsNTM2o1rPmVcoSO+LPSwKe2DN3vwPS1b568pMsV8K4Hv2XWgOOWXNB/obCp
yawh7wRDQrNYXEoa6QE+4GQZNlWCcopTPUV27rGR1UKpKedTwtmk/wE/mrxT2Ubw
nGaSgCTMmMGIhqryDtfpYbcqR+kvGpsk/J+v9tBSigO+QuRF0oUYAQoP3ruOF+8B
mU6GB8RllxNgUbCN+6A3zwUJBjYUkMtiCbYg+AKyML5BBOJfZ8A3dOzOBfQ9s0Ur
36RvFAzyxdmr8fS5tm7sg/d8t4qOm/EAkY4rM88MRS5pm6jSy9Nybj8zBciShZqb
TSulSr+AzdZiWTwx3L2gcyHFSzGch3+pU33dWPd9QNWbWILpIonIG8/rbx1NQ7vN
aPGkA2gqEUioyCVCb0/mORt2E+nn2qV16/Qp0vc/i6iwtqo2wR7pkFjLkjjM12Pb
LfWd6wt0owWwZA4n2iBwV4bqfQ3E2x0I/uteXs3XasHW0+aCQU3ytUUp2YBtlCeY
tGlIeZ009okUAZQxeu56CR5weOB4Q1Fy7E3obZGYjpRMAGvCjgu3tEQIQyPJj2dO
uqr/4/gUlg/aDhWJUEZ+URomzkuS5aCw+tPs5de8gv/v9zjI6Wg4APJvc1ly6oHo
k4YsPIHl9fT9eLG+leLH7Za37JFx7cUydIxVWLT0LJskHu9phPnkrlp4bEXBTrpw
CjtvDzoKy4KkwaQnJzEfIqSKsiO3G+Kr48Bx4XPMTYx82hCC4bg/Ch3EUrP3ev/8
47yumLM3JPFMMm8JNPzEs6IQ/geTtyoc11gFc4g8taf4cgUvj7wWF+qTr680mDim
NekcYxGT9XymcKcYnBW6L4XzKXpaB3odw7417YHCcy/SCp0orJd11kPiPs04lwVd
vSSfWr9QbYenIkdSxh63zWDcp0Ez5OIwYr+Sa+IML97iW7DJvDYKcXqmI4ZpAC77
6sDqKGpqfHOic92A0PzZDlE8F+0zWS5ZkQI8JuJj3lhqgE3yefbY+2HB6AdDxQcg
1PgHf7dIDDuwhf6BgrQSJtZrxXgAbP62nOC7hEqZufBHdTNNR4I8O6sS9z5Jg+ni
zesXRCJ4X/ezpg4Ubkl0Zwqk22h5Y+K1l/v10bJbjPu0vBL3UHhOhflPbvZCQNYC
drvWpgVXG5ilvkCYKyUzRSR+nKCMlhSmD10Jq1fVw4UxMtJQ3qhxUyG+5qa6/CAC
F+2tisKqOfd1E+Z4siDfnEPFVKH4w52zYU3ftdcE4wggSxMn+uRpLy0+EFaAZS8X
FpgRl+MRC5xtu49boal3Zk8g7MOxCER/DCmwXXNShNBx/Y3fYkpv6yVgFbOdzeU7
2YXGQyM05lf5oknOFqIxqy5PT8Vp8O7Fk6qajfkEciFlE668aKEDl5YQhNahV00h
amlvl6DmuOdcutxmcU3KHy+IunXSs8smyWeACDjMqmYis2xEm81J26LoVZB2fgO+
r8IybGT3oH6iU//wVSM/pW9LppeUVKsggo78rrCxn0XuyJTkcUjhrGc/ype5/yqW
eKoxrmuNrIPB+4vlc0JNdXqoz+BQGpHX20/ku2ZtewEw5hx58UeomANfuUVChRU/
TZH2a5rRwYhC/gjirQiCeTUz4Hy9yMFyX2TIgbhEPUxE3uPraOg4pKDKEbDtfdl2
qf3MhOLDNWIJ+h4NIx41RWXB0d4qx7MNWOb7nr3usld02qhTz661vfSqQvHO/Gb2
6uQG4pPXBasr4Ejfrnpjv1FFSZY6VVn9nouT5+VLJvFV4/VnBDfWcQEEvV8zoFbR
iRoBpMD+o1SdPIPRA9oy45e96nofBVbnKJjtha4PdSZGaL6v/01UUh4QrG+TLQqu
Hiv0/q+yVrIb7Y/Orte+T4O6xjQ3oqGNevi0j1ioWc8BI6X6ww4EahK7lixdWWg7
yy0uCIHxW3i0kzK7arqjCGUz9Gd6ARSogEgiL72jPHqlpRD3iKBRZYgCnehxT0nj
np4FVjHRDRzMl6QE+nsnYngtHMRhwXrd+uPzuizGwZ8f3K1RjmLJFV7O+Z2YdNxw
IbvSkwEV/4ENEt9wxDc/tSdaHwV82wuPlatNqCiWo4vu55cVzFgdN3MdNHwtPMzn
KKbcmflD4u6rPxgkd641prf/H0S2nvI+X0sXkJ7POAUqosKzlZzgVqBQq8Op4V9z
Go/d+QxesUajtW12FuCnnEsEXWNYROBrwZshmeScnT6ZwoxnNxKsTcDLFzXjlIvk
6rcX7aalXHmfxTiT3XAU8KRbHTx/t5JhoA+fj9Kn4E62cvnwWKIGRcfgtWUkFPIt
GSTpQi5GlvqmxqC80VMA/uECwGKUAXpeiO/0HZF3bzg3pIL3MJVDuogyElfCJp6W
0DYRYbayeddBzhP6vSK/+bNtnL+HlA/D5KZGl5xT91i5wxK2vakh7iRD1BViyQWB
bw5jKB0nTa0v7gdAH0Tb/L6g3hB0psaurwMQF1yQ0K4YZVjAhMeaNv4Ezyq1Qd2x
L5aN0/Iyqk7JUvjDz7hkoHOVdyvciAx1IWn8J9N2RmNzMQK73+QdrveL8i4uT14O
afYdFNobbOyxoqy9JMK/8k+0RwiUJ27OT6ZLlgmjlLsy8LPf+EH6rHgI5LQ/t9CK
cD/FxN5rJGTRHSh8UPNg0ucQ1hX9MsoGfILQTAB1/MCR6jWpjx6y3dzepkdsSCtL
T7oTTX/aqYaAGmD5I4M7NTI0ztDXDjqDCgkmBbbbCwktyO3ZPEApc98SCEM7Zaah
YJOdjmmYPKnn9UB7Xh2RBlPNVOPEHFS7fb7D8d+WSbF8xX9Qs13Vcz2K59Vn8qDv
FH249FjdjvOViI6HCdJBnXc/UTrlLXsq9zKSgXBlBjpMbS+2NCLwSIbF7NiZuP3b
N4M6Vg/mbI9L0Hb5lCpTjEEZyNu+R9Gn0ykDi+Y72ThdIRsiCvsX5f7su+Jcavb4
Ja67isem341hZcO3iDuliyzfMvUp6hqMnfZw+dSG4BEjOSTrZxZDU980ImNmVLD4
w8ZnhYz26dOgbH+SQo6CCUQt6wavE7pEPLSZI0F2UyOZJJLgsAOjzdZ3oPXOavHh
28uCSN60PQ2lniWJ4FjTEoHRf9I3H4WGBK/LEi8GP106NHGAz7K0EvP8g+CyIThK
CXwJmUfZzHIuMagklkbl1Rdy/329x4t0wLK5tsJDS3Uc5L0AMWqOm7s5GxedGPdu
ruCOArQc7F8owjHikYlDfUNWw+9BF1qDBfwHWMlC2r1h7gwUBJ/kztLu0uEcmcxh
LTaxlsG7nJZ052aZ1ZQN2yqai3l01yJESIqK9Fjs2Jx+h9fC/Szat8Jhmr5vAG/6
aAm4pVrYVZRyqejavzAJPsnOxjQPt/RyGCoKXQX3+XgsuycXV2GDSld2dF0Vye0O
NfysBnSijLB90UHf7gGJt/8B0WvtjbPjNMsAf3ftnkU10RvOrZIjfNz3euZxmjmK
d8OO3PoyJNcapHXzRO1ktPRMFFBHY35qYr8mgJsaPBm7T5N/stMg1iglmHi3xdIH
auboIR1cjXqdN1LIlZM1O1K5Tu1vcHKQQ7RCAENiQ1SnmlTJPwtgXGWBtGPFmrD0
Xmyy0tRxts//tXGM3tmxQr1TNMuqeyIGbaMhb0/Jp14q5brXSfiyCzbXrYQWL4MN
tHwN0XxLepuu5uSMTcq80uH3u9PW/jIWIaIrlcTmsnb3/Z/PbIrYBGj6201GRiAS
P5B5lUbymSwL9rgFDAL0QLKUUSG+eukYO3R/cPJHzXR1HFX4hTWraxnKJS1+bypr
Lqg0f54thXMspEzEyYn8bVVBYPnLG5p8B7t/PNcbri5XiusjcYA2EslGXyxtlGrc
Fj8EIkI5204ZCNgS+Xo1oYC7/M7LIScu5GyZXe+IwXZxt70Y/4RHJUIW3CcAzg8a
JYOWP+zNxY7OjgdN09mM7KyKyKIdjxznAvEB5eAdr0uh57dtzfCbbGbYSo5Q5Qlu
mFcqEQU/TP/AOJga6USZfs9v+b+UADUEOcZSDnKldOwixdXCNrQB0RZiabL2mFfp
L3MYebgUlUDP4Bf77T73kI7zaSOyiBSTnTSt5deKTmV8Q40CU/VDCIUfgYbywWux
kKKYqw+bwKZ5fVAyAiV/djOPsLSUj+yYVSXBErwbtqf0OUyfrEdyxN+kPtnfrOIf
HtvPhA/PuvPCvfj5TkKvd1/dvfi2CK4wfrvEw327KdP0D0FPt/afwqw7IaFXfzCR
Y44Ib9T2/HFaWhrnu0oPzEy0dQC73he8fhNsRt47oYtiiI8jxymZuachXykZ7Y5W
ix8u6NJmyvKGlwXDVHVkDIfPi7Ol9GeKgdKyTqRdKkBUrSdFK72MPkmWjbFAV76Q
PO+2yWBkm/Bt+pRv3QLguEf3p5I9VtrUQOUmxZNUcFdkuzlU/zJ75+DA5UK5VKgd
pV/vKAejuT/VR6FM+hSX4sdC4IWDFUVeoa9XdCBSfDJ/5qHqVwBEXI6VthUulY/S
sEROUddkV5Y3+42m4f0wglj1jzfBgMfVLteMJb6YGwbBFf9icdYekKftFKGv+lYO
P3aPU+wmUOewTD5dusY6cO7+OV5Iss3t+MniWWikSFG3bPp2HLitKdmkFnUkWXJC
l0cXOutcLxRk8+mKiKvjFmt9yipmuDwMxXYdTpPIarPpoAmEgGEsYTBlQkPBAfqy
GYILBSFY9xMYs+sJxvPfOdSX78+U1O9Be7ZO8tsLqlvI8ck+BL242fElJUFKTO2K
pIdmZsQn73cwJLZwg7eC+jDvUoAv7gYB2QYkEyssfObQYXf9fl/qFW8z+dLTREDO
IcO3xyh5XQ2yhGKV3nQ1KtV3Ek6dZl9Ico4ZEshlvU6l3/89vgv1qCVL2WEm0D4P
poP4J/6hthxY9TMHAEpAdoTOUdEeJCFntiWxDeC5F82ZWcufr8ANlEli6iTd4gQK
dby4rOz6CnlInqSRiUEFTsrrkqkuEcrMmZh73TLVJ3oOV2zYclW2XsjpvsjOJWgX
mbn7hbKaEyslIqb1zWyQACDsvKuUWdaeoopTZRLWUsJwWxnVgn/vNZoxYlXAP2M3
y4EOtwIwG9eOVfPlTPGE/NvgUod922eakIgU63ZjOKLYa8z/NimwalcmEX85D4aO
ELXGitzjg3j4rt4J4E1wrBlMO/GXbu9wHfpTJLDYnPE2uhUZzTTh1YicDDis1HVt
QowAnFvUC+8syzOcc7GKweDMrejn4SuoqpMc4EPIfq5ADhnhQElsT+aMfyQpjz5O
YWNUy02eXh0ocSoW5MT2+OZk9gKvpGs7TRwfg65zmNcEiOIOZK9uR1CzAc7PBb1j
DPFvmnYnDKAIdfgNCO+RqRH2u1ATPOqGXtXOrmzLXSGn+Lfr8Ho4sqhIzM6ytBX7
Dj7bUXCB4UEUZIEcMQU6jyArFLMN3kpavTIRH/3sD6qYQ9MhlQQ1m/n6ZxoPfvCB
xpWlAbeke1ZMxu0qh2N+3oSkWlkqYet8M/TNrMMwWvUbHs2WEzq5kBpJ/iJFSYmV
0z7UOC8/nlGpNc9IcSGNxKij4MravZJs2QVLCAqfGU5OFe6voDwSyvb3WvqBZpNY
kl/q6tKNHyNf7tDPd+l5q0bRCIsRrEcFvcIDltXB9WI5/OlQLdsn57TUI+STEXke
kznXP/xd6M91LY6YDLANE0M+vUYGS0WdyZcp7+VJVO9oH94u4gyt8fo8sx7U0m4G
zqITG53Kx+hgf0kKycN0ZT9otytu7jPLMf5+X4gMLPxHuJnBRzpo4/I9s5Qp6QXU
83vMaxyT09FQ0OO1AUS2iheSmH+KNM/8a/u8I2gKE+1kYAh4i2Gm6KIXzQKKOfmv
w7CXo58hRpkj+wpByZFtDbuSuyrHJUmFKadPZz10Hi1sfsBt3T3VPKNNgdD2Knx8
iWHLbHEpeDko1K6nsXTLV0ADdyH8hA6lru6DjNz471mCouKvZXhOv6BOyp7YVwYb
N6fQXMM71+TLBXyC2KolcKig8+oc5+Q6l1VYHYHoAkFettknfe5K4FUtc/UKeY8k
y5D6/PeQPqrII4Tk5BbUQMA6yJVpMEdEUlTfcdSq3UQrY7i9Wi2vkh5a4WjhnS+l
n9DiZyKLhO+kx6OAa8YmSDhnrEwPE5fkabgVjopZfm7pzpJrJDw2BN8ssorlSyeJ
aBoVZ6tW3HNSx8gXSMW0Dm+itFkY5g7mLRCbdm/VFlGQWI7tMQbvac4JQN0NuyuC
OBg3N3twykq0sgG5eA0u3mrX6LqNSSUbOEhZu+NDxKc/SrUolczTB0Oao5K7+X2d
rBA8ojSK9snm9sUKnSwUHcO1NJCNFjQW+eIx5NuXOKEgbpl7o0G630VtfkzDT1RG
KZBmen1/4DiGrEJDu15EUZGihvd2GYNKk9YPruVHwio0C7GGTDKf8J9d+2F876l2
Ymtp8Earyhtmm9PaHE3Fxba5rXH2ZBTJrLiNdSG8bASE3ltaxF20wGTXloIcDkKl
/xSaFrbdJBvdXKMfFWSrJtY64eHdTkhKhAx8S4AEJAv1XmvbvGpdqgDgHBbfWwBn
ZmmeDJulGLEp0Va1naDdQzqCl95DmK3fcIVlU9xyqzY7jQMMOI+pxxTcCsurZZqt
EmVew7w8e4H8w0vhDpraxTlwngc/rZsh8b3WfwU7vNRe9Cdqo+dHr6YGTvkZbA9u
bLYLOJODgyeDT6l128Tcui0hlKqg7OOsnfwP+mxWb7+cdCNqS4AbtZQL15DP8Qfm
8v3VZt641/2to5++CHCk7eNM0mSp+HeM775w4iSU183PEVNmxBdl3pd/knyl0/TT
IcooN3IE3BX5r2ZObQBlwax8WwMy8kC4P0iUq+XRkKzFy04FfN3D+IlQsAfy5oRl
ADHGI+LHiNaHLzM7Tb5oIYJ/E7o3TVocqN9wqfV7iqX7IncJCSTjsom3B35u8zHl
+25m+rjboL+nIdyKqK0wV2T26ew/xi2F0vnTvS7Kf+t7A+Z/AZrq1d5ozg6jko5M
eeZgTBlb4S74CGMfnHIIxZb0S1bv7jyG4BN2upl/V1EuQZuzadWLJT+qSaxSz9XV
YH/YdS4SdHdJaCp4qsMAO47QkMCoCsq8p41cpa9oFwsKkOW35821bOSHtrjy4pdq
LyiilagMIoB12mAkKpl6UXR9IfcpKF3Q+HkYJrDCtnsr+oUQRTHAEx9Fz9Um6yEd
3S130eoRivXlUMKeq5+mtBAOOcsdtThUYGnmAG/1lsJxWJK0rEIdPvAdf3vx57fj
a6vx7tAik70gNtOTKNJZnGx32TDLPY+VIesaUkxu4UQ2FXpkvJ8YNyi+SoqWVYNk
JyuH8a88REKqtYhG5//rD/MabsF+tTjP7ICx9B1yU9k3vf4QjfK7AsRDxVXWMJoJ
/cOqNUCzc1ZsU7mGCFbm+059b5mhuH/duhIyWm5qz7HYu0mGl6AK/UISoqvIAJWU
V6Po/+3tRwv1Nx+o8TqgS1c8NzH0qkUMCkGRQmueTo9i9wRzCtVWajo/+ywU3b5F
5/QuJ5ndvIRZ7Lp1iqYgCl8U+bNXEuzXYbMMBJyhtTOs0AWC4MK5APmmXIdNkFGl
DyERVZJMduQBpbLAFZGWkQ+l1cTVyPJCU+te/HQgO/aoSnIuIvPQe6blayRRfCqI
39sR6KY3mxvlaCQpS+MChs9VwIS6hqgAVgi3VL+6M+VD6vIgdGJTouhtP5dYT61c
vJQsGQ1s1a+uRaDWwnpKAEpV7CtbmcDzouhnwy/W4j7TYMkwArWdygpGpgrcvI8O
30+ciKGE5oBhT10FGqs0Wj8LcmpgfKi9RMeQVcv/zfYpUxR2lbzyHs9ePnMjLxK/
f9zH2wce6wxGHgYuQ2ZBojQIuL3HyL1awAKkMLEGQBK0IM4ybXmbAAQkAHvQhazZ
4GHRgf8SfvOQDLX+LReU8NoCWZQrm4+6DBDJN7+ev6JYpy32ZOvR35HmgHsBM9YL
6cMYWLn8s1tGAxkf1SqY3hlBz4EWifCns4Zsh1ZVMTfMNmjS5D9qEmFKugtTMS7i
LmMWYviIWtAV1z1vd51DMZ6k19dDiAA/+z5d2lTGELyopOiVsZW8QBUFOS2O3QDO
qR8szJCsu9FAkVjcJU/HtfkRQ5a29D1G7y3ELCUofD8u21zKF2i7WuuWHM7PrDy7
S8TrZD2P01CDHC8BPqU25zZQkjhh0AKhfD61LppolvX3EH74PSCT7bUgZBa33YF5
lkGjQPkNUt8Gcgio/X91jNQHE2kHJHQoZWCLSzsCmXNQd4EfWF76VY051fS2Txcb
21YM+2ZhIHkGkvDhOmr47hW9l4RAx1tewXpaYarpOBl9hM9SLLR2JzKIRGS6vRKv
`protect END_PROTECTED
