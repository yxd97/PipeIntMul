`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FucnDekLin7K29C2kGfAlxi2EElp6Pi8y/deIlT7Hu73j60RlNvwBbSNXRs8J7kx
Q51pQd3DSPa+xMPWbZo1oybdE/26STEFoxVljdBTiA6DPluD7xSt04c7V51DEpAv
VQ+XhqkYr1A7JhE80wpoyJ1qpel0GRO9NOLgUOPRFNdAtBQuEjE+ctTAenjU7DWZ
cu8EZVCPp+3KRjZq7tyy8tLKdez4vXPZAXQP/Q2bgBc3pNKAzytl/FX7KJ8YsB77
VyiV8QPNYXXNKk9XHDqZQ3ePC+QDY8iUwM368qy4EPOyExzRNB37Xboe+IUACB5Z
lvHQVwT0OVdJUUSWbJravxsULNuH7lgXAEghssUmBcSU54x8srriZngWipZrNfsM
j1x5Ostyqcf9P6nGyKF8qrYcmgL0XX3dAn515MtKnHVW7/LLSJBqHQTtjrvtr/Le
gCtIJ4lfQLON/bhEtAsBhqBEznrhbikqPRLAkrhvnC8ERX1LVqh9K07qOdQRG0R3
1zuCH2wl4PqMc90gafSLTwAlBEpzNJ213esdoioW9ot7KiQpWi9lM1/4hWD97mSY
lnLbn8VoBzBjXhkcLJdf+rlhFj+q59XekqOA7my576k=
`protect END_PROTECTED
