`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mwc1nAkLXgtf4SaE99QZmxGew8e3xjTFXtUwABWSYqS+fL+8W5w/oa6KxEIff56w
QAABu65hwnEqpb1POcNh9hZZmvWgSGLb6pDSF8J42DJhNepdpGfczCXklw6SjRXc
rKXfVCDhah1vHuPq9GW/B3Rt6QVfx4rW6TL4woR4Su1gVF7v5D41ferfg1cy/sK+
ghPVE57JfiNmc2giXm0vohN0pOk/X+Sg35WIuELHi8ZtmErojhki542fkQgXEiG1
2eDyLvd3yGtpWWZAQewfieq7s4iHpQjBCh39Ri7KD5qOmP+n00cGfolDHAS1lJvO
K5kXy2p5mdxDrSQqFK1tBThtu+/VekKT51uGxgSRR+o77krCSyhpC6LucMroMEQ1
C5X5YbkouoPl6XVC/RIOmpcR/2Ht3Y8nhNW9ZgHwlUDivjuuS5xgi0jVIsEMSYqG
ZeS4mc/GaTNL2D8bJvhOHo237cSpspzlWO1yeSnr5Jk=
`protect END_PROTECTED
