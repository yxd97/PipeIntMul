`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Leub9SdgXh7G8WcjSDdOFfAvXBYAqFGomgUVSgzV53C0mDHC+plZxF9lycRPOgF
Lo89LB7V9bdEnx4iXwhiKlG6T2D98aOQf+EKiiYVA9UOgvJT/+LrmnxltG/yA0iJ
2kzSRuRle7VsA7wHa9tRWM+HaUON/rTON9Pqf24LaZVS5AawyNUH8iCA0cZwDSyX
HvFPGfOigOZxhrNDhQGHO09ZpG8T8Sujjvy5lt/ED1dnccRCbrf009ONx2aAiEO8
LOSh43rEkydo2PqJPYdQ87yMMrjJ5XnGkq/0P2rTYbK9AThJvb45fNZ+LInPOh5j
ija6Nfd2vmB2Iz0wnMFfv/CDoorhJnVjoZQwCgYFaTkoODf5l/FA6+vviys1xVuY
hQsTxyl3+OT9WJGx+4I6A762e9LHCa048fUwt1I3XP+UfYlqcmhTdwFiLc1d+Vvu
Njhwqz2Ws1uoJUGCqeFhIUq+CCP7YOqR/rRpZ+VtGWRuQkdAxTSutdDK6nM7HWCa
xMIb+ZNFhzgFwypbEjymC7Z36Y45NfmwfWqPaTxjki514Qcnj+LmniKNKY5QadZV
UmPa9NgS87Z/EJy/Cv/z/LeGwf/mjUBuoxSoL6pae+6i+VgzM1FnTJkNT7Awiu7V
uCsDkyWPPe+gYwGeuaIcZaKEvumo6KKIb7l5I/35qiY5DEK/G26+3wytiQp1lUKb
8UeHSdNkWATVqh/lu3jxfjr2BaybNVQSNHNB4wiHZ58ecTr/j2PzKv8vV9nKSrk1
Alb+Vf2k/qN7bESfFwbxxj7Hj/5aiPq5Lnt+jeTNzQHrdrV5BcyOgafrci2Z4RbD
9DlXzspRcBSbN08btRZBmePza5PyVJh6t3MghEygwzrpuFmO+KMsomShrls9Gkq5
xhjdr1CfdulvbIjn8CIQJnnp1BnzqlR+YjPdQHAjPvWCsequNJs8qQb66qyltu2N
OJz3JDnkGCW3WKweXJJdjgFnR2Vffd06YxZOTTaxGfJ19AzKbJmzYCeNm8N9xMDz
IibMKFajxeslYMg1XIbB2zWTQJrhtzAqSHBD5GjWXK5mRheHtzboN3vgeAX+lo9b
E0NgazEGUbGHNkVokuPTHwA7uTDNCHxfSj7J9kX6b5HasQT5qcnXKQZxEzx4rZxt
pd5JjS1yNS3fwGPDgRCl6SChh02fRSbmZzSPI4GlPx+F/ZCI0pIQPsblCUyjQKqw
tFS9hxGnvoN6x0Xl47wEf/idiQtQW/ZTsjEulnZfVDHWV/JG93XZdqcoa4TWR0sH
jONm26VuIlVG1yC0ZqXi7SIDZbQMSC4YIsixZIETX9jIQdxXvRREjbpzUfKg/m5F
XgyIrYSHKv+1XeulSK7yhK7qby8fTFKyhzobKE41ZMeH9lNFqsxEvl5ZDxsQCe7j
lnhRUTCJzKPKG9ADEcVZb14o8GeThdi/bUve/PTTTvcP7D5C30MGlKkwlQ6ehZYV
U2grC9YutVInmJzM0l28QpsdTVIJlxO0+dtoAtrFe1Fka8VeKP4r6MVJGJTmRiVw
E9AQkGbCy9IPGDbgwcwUBzKsyU1yCSad6yg7VbSmscZ54/MuPtjOP55bjo+03hMw
d1qohJQqSunI7DF+kR148qNZMy7+suJVnhAR/3QZKhuAtcsv+upH8usjgY1Q4iIF
dHBtnfZ3MHLjSo9Hm8nV/bsOzEGaMZx9mU6es9c3RADVXPkWA4IyzpFcR+vEMg+c
UfzSFP2hJ9Q5MLYzDgqBVmJD/6JZEdf0EDPGnn5Det1rLXpIdb74WUn8dEybxuYa
x+qbB36YPdMk7GZAJZG2C9azxH55nSBr6aS43Dp/HYvPTd8bGlfP2xyn9R9wnKkg
joOFQni0IWhAl/MbHY1Dwfd9YiEM2M3UE7kM5CEXqqM0HzteD7RzhS9XzIT94V3T
yPgRzfeF4Ptql81K5oddLZzL66JJOwisio0zHmL4Ozg1AjyEoWcJthuTkhNRPdwi
vr2/jGqPfhH9hgwQPjlQxmg56YRq0Wwnjyu2N14FDD00T5BFLtw1iZqI8pyocyr+
ZyY5kSTkpbsYskd5jUGP8pWCG+d59Y3kW3M2qZz4mekCLaARslf/mm3isFx8ZVqN
GPTlbuNWfYo15q39hMTSdl0xw2iJ1tHVR6QJOLtD/Uq2ErZU/UctcdYrfivFT7s+
hZyOBrBduSE8eBW3Y0D+tjMdze72F0ABOpcEKUxfC+JeQRT8WYkIkqlooL+gCU2m
T8qPWrvc5i1yPoB2m6ZHRKDRuLpkzcmYmNJUBwUuPlGiUreW36epFSRBGo7duwUv
EU/fXXVUqjbdixOpc/AzqOE1iK8MeQ3/VRlozxVUSEKvbFolESsckYIJmj5wrfIw
bPf31opO6VyNG2r+apgatANWJqN6fEtf16xErgNqD2LOsCYRTPuRn+xFN183BD2l
3cII07mxFMQ6eIkU67fw+EvwG87O/ou5Yw629VIcrZ7MxVP9m3Rtb3Aj4Ms1jai4
b17VN1TMVSoOGAD8x7l6xbG1B5a+c2hebU6EylMtTh4=
`protect END_PROTECTED
