`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dc1eW4nwtTySBmSPjiuZcLZ34fJUcwZ4pP/ZaizrxcCZWDp41v7mKoNEYMFlq/VU
uTI6NZeVp0cM7zAejoxpjejQGUSG0KHWJQZfKDvxJIgiqZK3h+73CRz/JERCENuW
qhNMYXW1hawLbEHfg2hEM1keAdNFy69NbApq4YDKUcdlNok7YD/UmoLnJglXtUC1
F1Oczivt+p0hZgv+8le4V7ew/1XuT9bkej5grjg7Irmbv10slnHm+sKr/TyUJLQ+
8oX+0vJnMRo/7gGVa4tEO8VmVod5ueJNShC2/1VBghA4aMrzNXP07H8N1eyCyUFl
6KjyYp5JrTRIJnvS7XprKQoDkEIG/leBlh4gaZQWJAWYF46oxnZbYjPZXTd7jya3
0C2JqgTu9DIPx+FiY9gzuOwLyV+VaNiPl/ZuqPhgp9pVyP/fPN0jy2ixku9mg3ic
gOYyWsy6CAOjrO9HBDCHFeIQXgdl5Pe4SF+S+EGRWhRJKwn37Tg/b16QrjcsjZBd
mYVT6GB+Y2JTvp0L4h5wj/VGlF7mwBVPtxONF816to/OpuFO7nKno6e+J9oZGqY0
qU4qgIY3HyD13HPf6Gd0t1z2p29kKYyOq44f6KFDfnGUmG2HoAfgAhItbRwWYNTv
ayiaq6rACJTLvQjBWHB0VQ==
`protect END_PROTECTED
