`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RFqVAZ0MnUiLDtX3Cq4RgN/CgCVLX3VZABgTxDWHHqRtdS4Ht4OCpGq4YHhLrh0
zaujqc9NUdj/IJW1tAiHfm4U2So8SGWptDnXKQhwmp+Alv4r1s9XVXfwdZ/UMNyI
t379KlS593IscimEfjsL0dwQ+eZTubfX6wsVdXOU9KMlBFumsXcLbVsIkdAwKowk
1vDAXU24+oxi5ztu2dRWIH6ldA6348TSi6Q4jKb8IFlStWmcCyb/qcmjeaTD8Rxr
JqfPLEiIriZm1tgt/zHM9kPL7+UXIVZYWFG74xG8whONr+m6Pw7BqT7gjDHnkdv/
hn8bZS9IvIhifnnaF0fTbg==
`protect END_PROTECTED
