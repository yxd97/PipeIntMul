`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOsxSgiZQXMfA4Vkj0Af1BppQINT9tRQ1Hxmh1/rwSP9QceNqWDovO4di0yJWTFj
YrAy9BGtnQ2725gJGbTVY9x2F9NED0eFRlXUtoUPUDt5Bhp99txks6ODy7vNSxcn
4Obr+e01Ys5agbPB0UNmXKPTItXAvaqhZkCdO9qFd93m5tr8nzxKZjJVDx84ZcP/
el+NrD+/yH+0xMjFLmCPliRqhVBfVb8u9olcY7K09a7Ed3H4tXD4bW363NXvS5W6
H3jnHwlblWha0fZofauXEzYyf84ciHIETet0oexwgOCLA+zxBc63afee+xf+/Dxu
j77jCxSvB58qk2vbXHg4/89dQyWsFuvfDMBObYBKe1dqp+DQsG08P4Y29fVdDmiC
yp1wn24tgGlOvuM7/zikDpkHI84XO3xocQZYeagyMpmKLg4KVCGn+EMlLwzvvg3W
CuYzrTVeKNqCHvfp9gwD4JddeZnx1xghZ6kAOMzhM98spIJDSq8bKBKh4/VFSLDw
`protect END_PROTECTED
