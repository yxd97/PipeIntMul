`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MLNegrsE8Gu/e69eFsbUuD+UpPYMW/1jg0mZeyNBwacBKdRPyrKt9e8GcYDDoX1n
C6oZeTxjaMe3hozWhM8Tl/bBPiCBC+deUV9NFJEWlTIUysHd7GULBLIiaYbLhPX/
rOQYkh/HWRfV4sDeIosN9mT5Xdq+A7Rru2H8iHtp0zsFBhkMbELbaF7icMvwm9bx
spQxAILXvzCOvrNJXoPVW6wKjPc/I7KnzztaKRZSVG9mAQ0hHwBro0dQvVjc9FQK
XHPAyjyts7PmotI2Loh2GqrvrDW60SyyoNQRDuTso37TasWchvdfl69C3/BTB6kK
PlCWhFALAl310+ihtWj0zYB0c/iPaAAOuhcKR0GMkOn3zMJ38OaPCWZ1jXDrMGxS
`protect END_PROTECTED
