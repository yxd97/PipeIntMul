`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U09gRzC5NTDPojo+GqRJ1yGDv4X+8f0N2vrnMd6XpWEsZ2aj5L4rPW0/tB1Eupit
HdCJgU8Vb20/gnmFwpQFTbqIixzhKFgpXfEa5pCr7KR7kiGIDc32fKpAW6RL6qS3
ojlvRC4r+6XTcmJBhgh0/cYQaxj7FkM+mapAX7mSVsDJ5FFutmf0eI+bYbW0RyX5
qeDPgAr4NMIUNMUhE+9DtvLT9M8LNCRp5RGhD20lBFF5xvIdIcM7MHExlq498VcG
2ucYqkzMyacvrB3I/4wtnBxPSJuVvQVGj1aQYk946wf+D4IPvMvwZ1bUDMWg10Wv
p383mjbmGPwAVhRb5rgisd2THQzjRdkw5so1pfK+7UJO0AAnTUxfQCqX6wo6IZi5
WyY6HW1FvM0P98eRAhkNqSAYNvYM/GjUeDXH5ob7BW0+Nxu9qDLA6+tVIan5iOP7
M2lOZfj+4i6SP3Yt5AmSWUNDzigv6EB1ScvSeyQ32JWxwaquNW7q466JLgR9yaTH
DkOOrQmNcnRjp2KuevfEyn7jYNikg8uuZeGhRhHPiG7/nL0A/3yN/bVNf+zwa2tX
vsiMzeSNlBvtvn1Phf98QRW9cDm/fVZTeTr8BllNJZbUZEgVANkgnOjWzCb7xZ4t
n5Ro/BfO8OO0xhK2P95c29GkqOp6fXzQOHGDBoLCaoNvqN2r4s3/g8V2Q2MWMN6G
4yTkDGWB5CH8a9oF+UqIMdXHuTYs6K2WyAhZPnNBbl+6/lbmY8UhpVjwIrt2Jeyy
BlVf98me0QX8JOkTcfxWY7IP+Ae3EU0KIbKWXmw3NO+fwceGClGO8cFmE7n54nZQ
N2gEj45LdGjQI2FzdkeEwqxK2SB6DgVA7H58kHk/0rbR6sSQWza12HO0wX2u2V/d
pbkMXYV0UaVstpVqPFZqsK7R4eDj6zO9LA1FACbzmClaCYPtsqvMRCSwW6eZHxBc
/mfSFp+dQwjL7KMsh+C/NSXDhecA1Ja7NVmiKbwkQ11Pg0RJ7Z+jdQMnp7uxqTqa
Y778h0MZEdj/5oXDy3CPcYLUdeF60+P/loUdXbKzcHQrdFphGQa2dcoXNXRuMhwN
BGfcQyre45xGdKrzyQHGHNmRWdRmfHxUML0Uhwykujma3cKCNgvz8srXkF2ONdE4
`protect END_PROTECTED
