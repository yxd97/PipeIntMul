`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uoa3pUP2H0w26+VicTdgWGkCKELPwwl5IvRDN0pFwhaOMF+RhL98XhxrpRV3tIL7
kKhj9xYwh6MrZX3fKh8XR8hDFeuEmxjShWyvtwvmBclWzUd+fEX7UIqyLcE4S21a
bU/YbczjAD4ieSYdsdI9cFOGqTMTLt9oz4dVvi5Oy6vHRCWZhouu2+9fqqaTCyGO
SDR8fSzru5jVEwRunwjTwruJTElr+Ur4SgBvRx+6PSM3WU5kEOMHOmFrQgODxQ7o
WluU1dDrDg/KPw8egI+5m2xpwYUUwOMtO/DOkILmfjs=
`protect END_PROTECTED
