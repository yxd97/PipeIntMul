`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VZxxu0SpBmshFNJDFB4b3Vq3SZfHUQLSrU0fmhb5BHYvLlnNGsLzQrNsQaPT1eQk
J5MW0J7XsoemELHOr/XYVh9arP0U87qs5ntI8k8xngAEDqATTPfDfnk7WauwWmCD
A6X0BPy4ShSK9q4fkyUQITBFe+EdlZhq1rpejqcVkvQnHkRKnwn6DJ1hEFVZYZJ+
eWvwJuxNxK9lj1kxZzHEuIbsnLBSoHYKSam5hp6796Ifzy+JTwL4C1x2RnmTvRxn
AO4C+kI/6LSY1r/ViRy1Axm3ZGOjqRWd9QMo8CWcrOpRvOBhi7TNu950n/ZDyiqa
3MzNINZ6GPgxaUec7muKdybLlzGnEkI8tMCHXzxbjbj/7dLY/1g11gxob04GWA06
3cv7Z98jlSXBdEIt1LbQ4syO/VAzLXriNYw8v48qXyhg9uAEljG1bX/twj3cqalV
LGrtkVuHv6Wk6jXvGA52aWCN1QK6Tb7Juowomp8aZcouK58j5vsBZrk6PRiO1KbE
`protect END_PROTECTED
