`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cB70/XpNeRZy7CvWs7A9jKgE9zoFJTB2Ej1rLOyfII9JM9n0edhpDY5WgsSGSmp8
+kLbqq7jQNvAJ4aCjf/n6VqXMKN3amXfRAV+yLaqhTjBdYJVyeGE60hFXNv1huJg
u4ywpNp/cMLLZt6qq2jSpyu3HLe+oB3G59lfrgHd4AbQLSjINeRW4vS6avTMuTgb
hxw0O3dTaFOUK+elCwFqgDgGBdB2357GIZA417HhWFvyQEQjORuuLrwoB0KLNXPt
vFPpBM2F6zyRbOFVnFM1UVEAm+OouigzQvyNMhjJ9+nXQGo8ZNSZj0PDGPmlS9pi
pXeUEid/caY0scB6R1BjxHrIpM3xbt3AFQ9ebfPmC9/sJCp61EKlZuDDgWz1nhuX
4Yrmjbd3MYTHM1gZs9AURucXHXwYepW2AVtyoSdPToD965aQ4AWoO/BSbtkwvhQ5
gxckVU3xejSwV4HBUMKfrCtJto8SZpAdW6cKIH+/fvzKRMMRgdLK/KnnGbwA8J4+
RqXIG+OCIDbTVzR5NiObZYz3cd31lp6ZDar6vFNUBQOtxHobXjgIO+FHvszfMns1
Qcs7PN3ZdiK/BNR0hfAVZRB38r+hpogOx+Km6L3f26rJhk/Ajy11goxftNHpSY7l
yuiXf7UFrv9X7Kzjb3FZJxW1Y6vyy0A9jLUsUc+CpYqcC6+GmezqZCQChru2OWDt
KftBjVWzSpEEUqrmwIi/RxYDXSPQ8jiv4qCCq9TlvM6bIrs1AgQokNqXkFT0PYCk
vdOHvgG4ANg/EhMmEnF35A==
`protect END_PROTECTED
