`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ExEVayQ6geWDz97x5Q+cxqOntU+k2ITGNJk/oRMkCw21yIOGgPU06AMf7z6+JO5S
62/6Ixrda4HVTIC9RSSUTnNWi5tcBqj3ENPFkvG76jgscOR7qIwsZcv4/sT+3VBK
KjjCSnsmsSKBXSBC6BIQAS0aZboRQTy5K45RdyZdgREizyqSTjCZBTeLltANQPrD
1GfKUfh7slB11SfYUnxfhM/RlhYjYnRQ9r6Wt1WsGr5kbJsrtDDR75PZFSdBjGbF
JT13A1gB6zbitxgnoLrhv52PXohVvx24YSLHvn30GfzzFVWBE4g6U2CnDVWKd8EX
2Soz5P0xUEvs+8hCTnv2OfVhUYEo32I7ljdILZyZy4j6oZLcROa+pYwZZV5dkYyx
E4nXdVYKZjGEekSpH5Cxrcts45EckpFdFFGkRDieHZCOtJCBe54QotUJA3Pj+Y3d
`protect END_PROTECTED
