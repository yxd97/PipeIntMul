`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
smi0QCKfPsMALTB7iysRdVWG2HGTgGLcUSS3JwcDVv/jgkjJageAXl1aWuGv4LtN
4ZvKlOQNpjW8N6LxdO20hTMMAvKLeHuzXScE5pUgZcDbcof1ekUmWK9u2Yl8ViGq
a2BDof84vCq+ArE7q3oeacIj5wF29Kd5SGIIfXhTflyR+YgrT5ArHx7Vq5hHgCpf
TTaNw36qCv/y5Ga4hw2/BnLncsz+AqwAka5hEi2fwHMl0h+eLD86bbOjP5Bw006X
qzK2v8dLkFq8ajA1Su7Rr6S2nLm3LKIdS6hq9ii6kP/i7lEEMPlQSD2i+CKicye2
iPxCOOfryf7hh9VuEv+/Oo7glGciThQXeMOpQ1m+M8lJI3K9RTJnDby41ew8wVM3
Z+IIpxoD4qLLeA5YkuUnRicOoX1moDS4mXUL40QF8Ik=
`protect END_PROTECTED
