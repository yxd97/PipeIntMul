`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/m1eJBOEGXJKYWdhBe6QLqYPAcUMAnaYNA2QQvu4GjQ5H/l+yoZCqpYA9E2IO3xo
07lxJd6Nc2xPqoew6TWsVxeZqkvXJdn3VMgQ6clOqbrF/nJKkFyoenus7+YhuLMO
hZ+zAWHkut4UAKxl06zpgKgAGi6jGVAm++T0P216sCgoontGKsZtg2GYnpc1bGMC
Dlq0bbz/qW3JVl8jM5n086SyUZe+aycOeqFBzN5eghk/2nqeAPr1/yOsCIRyOeXM
L5WC/2xTx6cekXghFgOeebFw3sYS7GY++kB+0GJaaG9jrzZWCK5hnEeNzjYCspLM
BX+g1+VS5DmOW/Qj8uK4mXaFTCtelkC/zdRpY1BhSN+GZybFhPP+0v63JPuIHCVm
l0UHEvfO17pZ9z3ELj9EWRWI79qkxq1xdwhlW8AEXm57xqPw/lBwcIod0hBk5A/T
ngBmPTh/NcfYuTd+lfe2mmNo6gUUh9ms4h/SaZN2B6dlsEYnRyaUUb19vni2tKF5
TZpREB6kU8dLKcU6Lc1bH7DPtm+exEjDCzZPvWzST5Gbxp8xHmYpZrW+fhOPQ3+8
VAjfUTEXK+ZXH/JqvzX+nQ==
`protect END_PROTECTED
