`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TCkXy7VLXPigrxWa0l+gx9E05/g1HMn9TE9flI1vEoqJM00st/YlDSs2lQRYJnOA
hpBNSVkHdgkTUuq3R5R8FZv7s/0UDb+94rCQ36U3lc4NJDcYklLJHwdm10xCuj7o
TsdwSmRW0+2MmrpBqU0XFyZkB5k8ulVAALuSpnUoE/TS0ZFprcXKxSVJC4bLty6s
UNam3mO9xlgbs3iEYu653SXKlFQko5io5PntLt+9bL1GmjgpOJUVHFx1D+u3GRSV
tS6YWPoZaQXzmiOwCJ0kQAItzF2c3pC+2fQeRM+LLUQSYj0q11UW4FvFcIInjtmQ
i7xyC+IP0zgNq7w+AV2H2qkPy5kdABECR2VmXYwi6K8mjX3osLt2qvPy+VapXu5Q
Jigp9l87HkBtDpfXhxuOE+NlAlJU6AK3yR1BxS3Jpx+3uNK5C0lskLbFYVv+wPsu
rHSWhuYQGDlowyKz8LPGWrDJE4TI68ZedaAqPwJzjX8=
`protect END_PROTECTED
