`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IzqtoMOnX4AAMHA5hoXKE/VWtfP6ZvtTAsdBBfVjOQlspigVzed0am/qV4rmc2M7
mT2pbjOhAUJVRTZ5O4F8fyzdDxy0HK6x9jVfDzV6lhEMspv21a5kCUtp8i2gxeA3
NPq0rZ+StNpvqIastGMF3JAjUD/ODKKxrlWtbypx6V4BNSo8oKeF/Ugr/xkMbGEH
8Oesk6hSgpNCtt1JO/L9ZtQJt9VyVDGTaBlYqDcRiw7iMXrH4Aqkn0r5kb0ktwo6
FxkVEQ+zUFfNHK1fJlMaJf9cJqne2X9f3nJ4wSX/DF7xkLMXACtwVAsIHEMYjbiR
M9/PQNzmUxclh/SROfLsUWF+V4BpjYAtW+J8raEmXlTVOx6BzmxHwMycTR+wVQlz
rVqTUSTa3HszSVAtWxwyxQ==
`protect END_PROTECTED
