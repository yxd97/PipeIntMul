`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFHaB/q45hHS1HbvH3nyMo7b6Y/SoxPIFdde3paJdANpgOrPMr8qMZDg6dBvLs8+
1xRdU6/YA11jPsU25B4U4slKpCzcEZvox4KiGrCVAcx1xktRIKhHBnvdqE9J54PC
+yLuVFkez2D/w5RP24P4AV+8P/2mqSF3uvYmJu90NNfF0fChOswxl2a21bJj0D4E
wvuhj4wrQ+a8nEihoN3pI8wPNrQStENnCabki5fO/1lw2Zo7NWn9jFUu3DwAmv8P
AJGtbY5JgRh3xdyvWEL2euvk7tX+QpyG1ISzkh4Qr/MDtRfhrXl2LzZr/2fBNJJ5
nYaDndl5cKv3PYMCumgyAkffU70TdaEN3p0B558bi67FaZyJe+lt4+ipSm5VfK8R
Klzk7K03OR0M/7ZoVo4tDHy+xl7WogHj4q8W928vb/Yn1KDUfk8gpjEujfANRSen
`protect END_PROTECTED
