`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nY704DWIWRvBswHoMFwUvInjkurwIiOq8Ths7XFBFY+TFflhYGSZ7SxwhE/RMEGg
s2ISqfiK39lQzlZrnIUDtlvltz8LlbH4O63M0w09WY2oQ4NirRfKHwTPNlJ7JMLf
rugF6NUJzzVZQwMHXOL9Kp+LW0K8F+4qjQfzf7mdNaWI7q7ooxw48dJ6C2mR/Xll
LbdaJ5pyUNTbcWySlt5LxJOKR6TeTev8ccr583DUjH66DXs/sCcFBETHHGMuAj3h
S90JQTZw2bbiH0RcwPbhC4dG2mTRFOIgy7REjZYUDxeTupl30MaCYcFo9BcBVaVG
ulX5axCKMP4w/0V3v4kUeJObqD1J1KPita4tNrjH0xsk04klsTb3mS5T8tjp6++w
pRLPbUl2MtTnu/wKd+ZLNuBOBM8GEqTWn62DG6SYPONAiY2wA7/0P69jaB5oxDWO
xcSVf2BFK3CaS9f1Ck8uPj2BxmDUZRtGO+yktNjlq3mlX/B66yeAffJQgHNqLLaQ
M+kGUhkZ58Wz/tNM/IOGNp3KuhBMSUJml1d8ZcekRGgC6CEC/JHSJmBqtxebAfmh
2xQHWGzn4oUdXBr7hb/XnDdB1nHt+FHY+GOg5TWc7b5Tx1qbyXm0grJnjtB2CiIs
+YeGhy2DiIEY83Fscebfe6PKLuBvQmBrnjvc5CfL39iQIjKwFjIONjy5ZcD+QW7c
t8jB55DbAQDMkNy96n3Wa32bEHQ2nhhnOoFOzFqJeQWvioid6sIGrwHtxcsptOfT
KTF7TLjY1nVg7nAWj0sxHLiECmzdHiLK41/Y+XriLNaIy3QqGL5eyK1qTZqTDPAf
nD3wffYOiBMR3OE9dyXWVfEdg2InW/t9xfUnEv9pfYXIjhVGh0f6lw4BzTfpItM5
ZkRsbyrrDhfMkpk++tXtKpmJnXDxzy2vWbSr4Dg1BwaB64pCNgW25l7XVoNh4QeQ
AN015MMZ2lXxnvDRlccE1w==
`protect END_PROTECTED
