`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7SaH71V8S80eO2JAQzEQbBZCVz9MgH7n1/nBNxsexJ6BGbX9V9tO33EakHe8tovW
UfrvT9qEcmfyq/oTaFeCMaCdbIatfLZaILmPS54qkBCofBj5KKM4Pc1x2g9jZLmi
qqrnERAkLpvY1XCxTKONXJQd2tyUfd1x29yO+pkU5DFSVlfg02fGK5bvdj8NwhAE
2pd9Dggn7pB0iN3fI5uAhEz+wMdzH9rdfw2PXqMU9E6l7WZsU2VBfpJWVLj8SeYw
+/mOxUkpTpPsSHQRo1NtrKKfsrCfkjWYzzP1LVqQjGsEsh4cU9TFXvoh+yaYpikg
XMg93sUCskNcimtQ6Std0/gQI1f4Ld0bh1CPILfFCVmBBPcFlvVtIWGnXCyDg3lF
f6goX9B494uqDuZSoklt0z+H12sTybBqYD9Ha02Zw0TvWtgpP5CVSdK5F6oBkiRT
OORypGW6veWWDcLScgyBBa2DXyADI7n5nztzW/q/cEI=
`protect END_PROTECTED
