`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zlGFTWbQKBEy2nHNX8kcwhGLPm1I8ZmI8p5cxRXZZi7DFSiGPXttV0rMxBuO1ouC
0sFdGX+N7gcQ80AxTuaeq16TcyfKPyraMEeJgmbKYH+1UYQUWVYNUhzFUpz44Dl9
JwEP9bjL72u65nk8NT2+AR1Nfom3zT0Tw4IT85cd4TwTjL+ik3WqH2BpQZP5QmaA
xhD1MDbNwOXs+Ig4+1uKlqzz3Xo2PJx5nESKfZwZv0JxP2AKqiqWPML81YIE1QJj
kHTFH+Ae3SnFaSI9U60EeMX7Wp8/wUxrUpIoXsBst4/r+cZSQKno2IFwisREnW+z
iM08Jv3OnK2Y5j6o27ag59FRb+Kg4NHpsZNfKG/u8Kh/1RXvCS6dYMVXGwj3zgzh
9ZSzAJmJRKNSch/u4WmRqKet1Nj0Yf/3sj1a0E1vla0aZ9hMaJj0Ju9grBmmmLwi
ucHL0Poav2LgTUWEDd3P6Nu0AnyZZFD/4P+SvC8OJRcnE6zDT/5ntuJRp9YooHaq
orjdKMeNl4CZYRZDdrTJLti/p6rsswI9DGFtz5W1eIx9fE6lawVh2DybmaFhD4S9
yMlvdlDG8HjXkchoeJhqDkcf4eWpYL4BX6kmxUR33L7jG5NZGD3lFrpk78Hm9cNM
xDJQjQHn6upGFFqyCX1L3K7bVHXG/EMFQYwV4WSke8AStJdeUlBWMnEQVFNo0Euw
PPblgIie+okT1qpISCgGtw==
`protect END_PROTECTED
