`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqepVruIXnqiXY51SEmNCm+q+ZKF59tZ0wr3LwlvNv/cxXtovseQ9Av3XHcNEIaj
0vjAWc16eMira9pz2l4aLM2N0t6RCxL8Ok9La/Vi3JvH25H+WpX3UhP03SRQuD8X
e7CzWCBnwbCklCVDj0/X2t11ZuqE356m7OY1jtmy66EUOqE+DvamV3YD5J2ESs/b
iubi8pcCpwyWqaJFVKa6HI+FxHDAYHM34cMxIqigM/XcDH70QejqchPwGOFBWzNz
wIlUBSbtFDvvRI0p+B8LkHb4NG9Q6sqJUQ7v8lrTres=
`protect END_PROTECTED
