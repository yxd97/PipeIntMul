`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jnt4V0V/4Ref0wPIxq3nP4hgQ2StKqGQJYD+BRfvPDeYkxa5viQ75i+kdby51YR/
RWIofYFMsHgPhlrYhTg2YhZXdD3JrK/MILdqVrjY/1MzQcy6Jjsry4+yZhcq4JHz
oQbXkXJYRsrqou3P+KePHKYswQ+FW8bclx0D5w9qq9qXGAEilpQF3Pz9hbR4zgXq
WQxNI4lTOnBysKnXGPYTKzXVf37u8Qr3+hVi1FKNHVzChwAzdQLCqYF/nXk64GN/
3/1gEp8OfM/I1lHoufxxxvAgowjODS9Uf94w3/2GPOd5ACLUhiuyCBl2LDoa9YQU
scJqBiNiZvoCSVkdMEvJ6RDb4a36C0g1uaE8XOuEh2836CKfhiHWxGuuTX1zvaf/
HvAuaVEl2A/WJyhf3zQzubGLeOnZGtg/lvQcxvwDEk3Snm4n5OJqKSzLkIRksbyX
xMap1crgv6jHyXcYMKf6FHAz/x7YEQIN9iSF5UFM5NC7EyKMj91wUVTvIyyc69dP
NedgSpdOoDyitjMyZFuXt5mJTkmYDhZlFcOv4jEiH+Zh3lP/h+dHSz27bALJ5m08
YAwvCn/nYfDp8SP/xauGHzumrjLB1gW/XHNGg8to7EhdZxqk44eECexAtUvrcJoq
Eo8X9c0FMmLJZcfkL3xUmb9B2/maanhCQs/pNgsKtjLCyw9q2DiqS98kAdlt9NMW
`protect END_PROTECTED
