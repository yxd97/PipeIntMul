`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r8UrEJ4TRa9PYVzxu3Q7Hu6d83TOXztnYVcwwl7ark4Dg41th/t8xXYmsFhGJ7kC
ZOe7Jlku/oTp+Iv+bk0ozCbSpGxaWH6GwNLXs35bBsrmPn24yOLVaT3sOxFPfPCD
p9yOU4oQ+aDbbtjy266T4sGGvBnKzdFg5geAYz7ekWJK3MxJ04/aBSfeWjLHKROw
MJH0xTKLQxlwc0FQ1ZJET8bTwBE5rjAOUB3LtXcasEObusltCUkAQCudx0oli0/v
tBvMAjcV7Va+FgrHkv0v9uaF/c5Hwa5cGMxnWPHMW7geecK9Yn3JMTDkEeNJlVtI
sLPmv/2CYe8U5jWdGgHL2bMCBafkZncVJXPEVq+3YJlmsEV+O/mW4SZQPS8+gRh3
UDbkdtUaXJfnssLiiz2PANdCY93fwoN1/RWh68fC0ti9yrhWbiPO5NKi5rhkpNdK
noNYow5QCxEaNnTztzrCo2khkwC58pCkwed3120KlnX6ihDjG/KvLYSdMZ1Zb+x0
joXaUAcynbdsNJEQN/EGSpa5oHs4i8L+hDEpFVVjt9QV7hVa7Ffiit1fVeRXUzxh
jwqxLrGhqS4uExCIsTEEsVQ6dt9USx2aEPogFeFiuUH86wxj927mtQ4rWiFto0bK
fs2mOnuWhmbtUhWR0Iki53egZgsQHY6R3HA+BhViQbLWgeM0hbIa9keTcSzfBH5t
kDbezCQWuHn2hSvMlzoS81kdUA1IlRttOl9B/ge78g9UN4POveRBZ0gEtZxnE9g/
dlG4IOXjqiF+BlEXXqIH6jcQktRQPr2o5O0CgQeTQt07oMRiR51sk/23cDF17vQX
n/L1NT8EQBPctq7SnjQYFwtcDzcPj3iO932TAPjmQzjeYwp+eIw+JvhG4d5JZWc3
PKMPE4BGyB46HSqWadErZBHOOYIK38KgL7qeHwKqOOrkgwNOV/982otnmrrcAp2c
8+S5vHclKMCASgOA/ZvtnDKBIrkkRUeDJRZZ7+kh8vGd9D9Kv3RLKTYcS6Ccp3MJ
UlNZ2VM3LP9a7Vboauuf8PloInUqG3C0oUv5F/7810iujD7ZrTdmdCXYMUC6MSS9
90Dmnn2t3QxHIfnqPuVKMIWJsDtKcNhujMOi1D7jiQc+XRanJU2LJsAhh88oJqvC
fjU6QxZhv4cKR/ZG8w+YflXX++5OXlFM8xl7QNz31R4+nAw/IWVjUV9URODRmXut
kDkv9KHityI+Ki7yUo3x5A==
`protect END_PROTECTED
