`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XIQ24ES6fMc39ijjnKoHMgKYlEhokIgMrQTMpslM0TuyUXiERZbIzje7ikdL157l
mHH/Do9oXgMSItJVR6rhgnVMoYd76ei1FM2ovTD7+0desEETEoQ3krgR3Q/MdCMA
MTK97gbX2h6GRr1BLUv1q6dSLMBGrvXRIkLuFlsa5OTu6sv661QSGNh9umWe+ihs
QP7oIRus2Wd7pYqVMJwX87Afe7NaJZu3AQbO5z2dAo+Mp4xUQkdh3TXCzvc/PjYr
t9IsyyhcX6GBXAtaDpI/4wbD8A6L0rmTJK/LXWoBEg2/OhqEnt1BpGCadRDIi6lI
XlVZ38v4dIbnlk7Vq2FFVDcJ4wJXxLG3zPw/7mc9aai4GIs/AV31Fktbn8rwjYAf
4QdxUplBzAu0OQCcu8k6B2G8mACKydRe26szYcjA462+R2pS6Zftonm3Ve46gr55
h7xFpOayIr7rCepanP+jKANmE/OB6F/PO9RJPUqUZWgXzZlUt/NM5vrPYna4kGQZ
`protect END_PROTECTED
