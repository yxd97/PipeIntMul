`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jhNbhEV5hnpufolTDoIzeWXksvsPg/gRTi0zfuZksof3gWkVvSXxhW1qHxagMl6b
9b3UTdBWogWOC6ipddSi0w3A68WFvSO6C4rjEmhuqTi81c3ucDFAVlWNhTmzqdPq
HAC+EblQmNrguIuiqnvEDj+qJYX6b0x4zLP1sgXUDmpT3Jv1wEFNmKp59EZ+z5Tj
ToH7qE5JMfuyfPE8eTh77HM6z+OAXc3WPDewknYWv1rvbN66jnIImo0m6a1IzNRT
QBhxnoQ54IWZGQd8UJhIIoPX0B6i+cxHvx6cjtqpRKmr+pl76kBUwbAUUpVAcx8x
js392iKOaHA16ECBu4aHQgAZPzgb13QL/TLzZ0Rs/uJcChGf8U16fkWhQznHdXIV
h5qw7+/NLNy78HjJ0Jgosg68l1Ie4RYD0FrW1iNVT0RlAzcFgND5qEItuqBVvzk+
vDoTpv6Xzn8pRZgmmG4DAptD09mjtNH7/NiCKeKgox91RY5pLlpnso/FyueZCGN0
JwGriL+VbOXkY1L5sJKerX1Sj4coPA0G6DyWJFbdyPaJFqDmKokbY/2p4cLwlPhj
d3QYry8Ofp4822WN1DNmg4OlUSZYkpLnQMJmKxGCnJY2Wo1Kub6dfrmZGuTn88iw
+RHKCqEa3eMbYQHa6UQIdmUpFNabmmJWH1MU4vMv1G1Q6M9PynLJxhoHhPkhup63
mlXbpohJbRe8J+Ga/93NbnsQHxW/+PpXbVMrPIdGKyo6lPjYJP1ZkM0OthVraHGY
YyohKfLXJThEcGgzg1MYAZY6pESJf0ujmWMmsbPT1cKWAt7Hn69+GLAJ1oR0b2cL
V3GzDlLJ8zWNNd+/EukuCA==
`protect END_PROTECTED
