`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EQh3xBCf/hSXdg3YqzTJWs7lhjc0gx5/Fv12ehlduocD9g79PHro2nXUDLr4ZOWX
Aekl3L8umGjjSfcpeEACGrs5Q7xwoq5ONrVtkWJEAPejHSWzfr8k+ql1Ckbzx7C9
5vdAymQtH9qqR2fb91TvHZdUb7k3olbS3MsqcKH6bbVsrl2+lsu+TcmqYnkvWacD
TX2LA6QeLAWLDdPqniRUKhnGKB0oY/vR70jes+QQPjHarL7mT/U7EgKUiZziM4cT
ZMrvpLLGKOp06X1D3D70ZL9oMB/7cCP4wc9546NT4bt8vLtRiAvfQTJvgF50Xe2K
p7ELfgEY7sYWyWOyJUmbsJnQ29+dsPKGfCZ4abQxHaZLbRIgZ268xspW7uwMFOpK
yr/ki47v5F1si5dCaJ27xZi73MBr7/uKFpYM7GmwGZS9SoinA3YxYuCkImSJBbT+
GlFMnu/sMR4JyFLLjR7dIvI2vYFMeVteLcEVO9GZbtpQq2dux6I0OL3eDZBoQHdY
a9OKkoE5U9BbZAvwppBef7fTz4gDrAVYf86kM8Pu9HjK3vp4Q4o94CbPs9XJVmCR
j7PVmv6SmleFMLvkwHLc2kAqLxNm2zeDvQBb18pCG1EQs0SepQJNlp0pfzWr9eQ1
U355RH+OjXKp+neYqXpwHfc+POZpBzPFqxvwJtDoJGO1btwQnvpqQcaj35qtyEbN
NoXIzAZqdBTHWh3PYSy2sOtgkXVTOjU9SgW14gTa2JY=
`protect END_PROTECTED
