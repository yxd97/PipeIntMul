`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ln+XLF7nZqyjS4lxHKiljvr5RklDSfBnJU/nyv9/jM+uel9Jo5+1kUfJKncwcsVW
EafxKnCdMSYNpRLFJbykRPMdixIRFtCEaZ/HgScIsJGc9q/bGZvB0tbHWbaSclWH
wGk0SMChYRx6vANPUS/n2mYcjgnpWDHirbbi3H28SDQqK9ECCbtU98a4FrroXuD1
9VuGgWwJTejyiuRyXXcyxIyVRiRNbMyQut8p7c2g3c3eArg+g8YpUETixzj+bExt
Xk2toEAMJbCjCKdH4n4LKfud8g39EVWjKFU+VQmLrtnGnZmEFaldfP1T4TUdUnXY
AdCy4Zvq2XitMKKm6Y0ZZid7BBoz53b6kxl1e6dH50A=
`protect END_PROTECTED
