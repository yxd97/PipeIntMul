`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQhlJZKzO56lPZYYBAgwrnADYKRdZwqcV5kQ3Ky7/DiOGyFg037qwJkacQxklEsk
2A+hz8jXDZEGCa5vygSayOAV70n7aPoJnYxo0kvxj3KdrT2fT3ycNVeHnBX9TYMB
BaaTMJZQaJA1fy1tS9sTaQKskCpH9084aJTLFuo41kCA7PuYvzQC5d3jOghY22/M
GmHi58bnKc3/fOmLd7rwOLfvDL6h9fmWRjLzOJ7xJsqWFL7X0YKD72+98sSFb1ZG
YP0z5D0DW6gWaObWa5ozXsS8ecRsE76bSCZFuuBDXgo=
`protect END_PROTECTED
