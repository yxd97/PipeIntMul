`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Wg0vAZd323k/1E/ZBrYrIqbNbKjGBKx+uzoOLfFcjVRKR2K0bU7pMWY6ztoRfxe
yQZo8bHH4qijFbDlYg5SumoEO8rKp6o0A8yBAykkBxseWn6BlT6lQOfeCzPOU3Ca
+9PMLdNkdw4yZJu6Lg6IAcBDeHp366sJwJcTDFjqWgFfxZi6QLqe/h46wRvFaZLX
0Oo+1q7M6/8078RzO64YU/a9sLKsR+zzGCKEOrIYkS6oFuLexvUXBbQlomCKsv+Y
rG4VD3p4XuXteNUQCAMw9+UqsUMvlaPC6pKQ8Yx4/Uz2Ev5fLt2NVrkvzc2TO/Uz
rDjgWwekJm9YXXo/baNOESEKLdSL80fjXY1+JJyHDRiS0RJBnI1FTEEnRoQz00R8
TkRZTu17dUhetQD4OSlvl6VtY9CADPDgOpZvt4nmvlwN0SYUWpNb9iyZE/xjCmzG
AdRmq2gjXfV1a5sdrXOK9WTTsH4Z6oo/Pd+nZ5Tn9IZq0VgiJJHEifc5EH6iuqUc
NoZqxh1pc5RT3j8lf32Z6Eghkw1nveaJfSePT8ZL7PUpUlOddL5qx/RMxGCKuSIG
90u7UZi4p8YLIsw0Yc8P2osWatBlKhtlmKWmAHi8Y2wzaY0XmQ0QUYbmaYWJ4Csm
KyP6XQ58rZjqWdgcCIF4QA==
`protect END_PROTECTED
