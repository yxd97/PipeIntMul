`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/E8JsFWtPNPCQombcvcJyjiBHpNz3O0ckVpRZ/ggN3SGvr8AIDsd0z1Ue3Md7E2/
urTZCm89BVB2KoARI+ki+LWwu37yaTW1grm/tPPp8AjzQIbt2qCBR6R4VfWqVwSJ
R/LXIVz4Zvgt845UrzCZ282cPCDViHnqixPtiqf8yqltLPc8/mo/eZQTo50DFkKP
vUgb0Owxmkdg5hbrbjj0zvq19wOVwXb3wBL+vNoIxZ3VDKSG8YQHRZxJghk1Yd2r
+5tkDuKKbn+mUqWUfLYgj8f/E4KoGOQikuJekac2Oh0m4KG4LLuScjbKoQC+BTDW
Jc/zXA28RvNxtlS7IfuIiX+N/OXkDfZNM3tIbXVFFWea1bQjlkp3e/RD1eWGTd6d
2n00sjWlg2TlsP0vJip0jQwGiKIgEj6ZTvGJN20kBB8GMYdep3E87jSCUonUrCBD
GoCY87C43pU/oTzSqdH5q35hLm8etYCEo/SoVulT2n8+nSq0ERJxTiImX4ATQy+Z
btfgDegLEA23WZ+pWgtqvCKnkxcFpeB848osaQg0qMTZlF7LoXB30TU89wUxYQd2
7j3QNy8S+vFR9I5YM9WJIw==
`protect END_PROTECTED
