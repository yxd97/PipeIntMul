`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pXBLbj684oKjlh7VJyHVqnJbYNTHE76vHXYGWlJkM0wOZ+q/UeaCsI5THkVwmUUf
+6j2u/FJdWCuZBeLET9A+Y9WhDHTtXNO8K3cCpOFcDB51DlTG4C4SHvLXxx0aQn/
VB+PvUMsMygAweIC8QpV4m0KkHpsmlQRYEuonP9A6mD/AlEzE1Cs45rT6SZbQjlc
wFyUzWS9nqtlwG5CQGPRWPyRXd03rgVX+AgVBHQZ8UP9aWDC5TSMqQjdOTqLrCwB
I6+qlx1gEeW+lrWVsjjtOY/gtN0uSMyLFdN/NNneUWmMEbaKLnujzqANp2MELTYG
XsLaCGQsG6eyuD+BX9bxYY1KL1H0VdJmZqmbNGqh3gWrYTbXQXFYProgdErAEBmC
1ZVm7xGIXJcqHs3i5pfc7DNd5971LefG++dHndMk7iFmNeOdv0Oa9OXpbWIJTOFy
s1KrxI/5zya8X5icFpE9WXaDkUu2GzZt/i91uWaHNx0CPCT5fHuXo9P4Nq2f3kPd
FnktGb4ab12KPOrhy+KjPLoEXT0Whc2Sj3QfFuf3TBMQkbS0RoOYBwxifJwgYg9q
bQqU/n+7EY9Zz/zZAZ/mI15gM8r3GxObLbW7uW3o+bvhWA6gv4EBRoN7XqQrM9jO
3BbLkM1tmeouepGcKyqI59MOJzsY4vjtjQex1gFPWcG4uiPzfWuolVqVJokhLHTk
/QW1wKA2l/o9zdC01UvpTxdMgZ2JnMCBEZBoE15mcCb133qiY4iP40d4OSAWHLzm
eqrQ4mqkuxgME31B7a81dZaiBUxzRy9QoTA9g5O8pwmNRT8e6NjAlPe4skCn8CEa
6UwOqNBcfvvpfsC2npeC7IrZeX2dlJZxakqdS9bX3ZWm3li1YnNLkQrLcXbqsLC0
ZOyzJp/sGfYyJf1ujxu9ficiVR5g3Mm7GBWbBLTe/YOvgxMr3vo83DO0SXaT+xJX
DSINEbtYhVcuuz+Z30D1aOpT28eYP+TMdsoeM7JzbX6ohUlHvXVa2L9b4yP2IVce
GOkP7U9nJ3MDgy19prdLIZzxDXIClWAoituCPGBj0RqhdhbrDyT0s/vGIIAaN25V
0oTXix/dKOnPtq/5vZgT1Ot1KIJrL3dIXViabn2ZN7fgN0oiaKWAXxl3+TR3XfH0
wDbrPXJeiJwFytqfxcv0vj4Dl9KiOuHxYvkAd83iUKunRfeh1QEkDXtnDm6D1WKm
jirzyEvXnQM3Ie3ox3U8xcFtuxQNiIYtZqvFRZwB7OFbU+/yCxIlxfufTAJT3is5
Wv5d8IHVSfn7t3BnGyhSBrk4LnTzFDfX8QJrwSkJFEgm/IfNEjN0rDclbOlTPSOS
acDj5bmgYm4de23o/hL5vS5abLNhKbvhNAQkba0UA2kPjBq9uNJgG3jSFfItutHP
W6SSS2KjBMlkvi6sVk8PvdXm33cSNR43rsxvV9sSEnHAb/WES4rSJ99F7aYCZAvE
S60NW735JQxBc0QQoqZ+vgffNAP+TyUCHtNeQr4YagHYEhtWssSsN7IBotW7EAwR
vxprApmb0siK4gFVL5FVV6n6Fanr90LecbTop5oiigOiMUqxEba3e09FURlsxjnH
Bj5HV4APH6Atw+t3mDWOm3bICnjGFAgeIF7bJRHKduMKF2JzeMiq4Q5sjXUzrzWK
przoq78X2q+ZosVrvP5JYGazaT7QYSeuaaHUNKoAvBOurN2VmGZdH67rTbbk9Jzw
Ei0SbgAv+9MZ+dVvocWrSAezD2jjQ1nYinPcVDqhjg/BfmmIWT+q+mz9VVDqiiVX
j673scC8fFO/iDHMkI9J/9z7KkeGuA0n4MjHQj3TT2ZxKFvRfekCsCWNahgEF7sL
MlsPSKRSjRNogy24a8D1S4RjBEUwNhEv05QwdXyGBTERL2oZVHJSupby/sABJVrt
72v4SbTAE8o77FVUAUFw3mtWhNdHkhjteAd5BX6+FhW/M4SEXDQ5/JTmchN6Od0P
vEMvFA92Ndjw5L2xAe1DeSIZBQ0/hc9Rmei6Crhw+PLhv/OfYAUpAa7VCg3P3Ez4
lf9Zy8H8mOmrh+0Ad8qC3AefG4oCEYlHb8O+qXgCtVDpTAF+k/oz2geanh5kq33F
b2taSX3mmjI1pO8ZBf5+D9yCc0vdQZXrCu7GzqooxXK7rTdw4FiqgNibmcAPaJVG
VZgpI20v4Gjia8JBInzU6ZsoLrdztJqiZ125gwtnqWp6GWeBRohHdlIf+Sjkpm5F
6HV72uzaxiChl2bX9NfHpvf2oIaLyVMA9tpdx7dEFhm+Q2o3Xbvl3lkWI4VaGLMZ
q10JN57LLb3gn+XIsCZZmXidQgHxAZ7rG0lNDu11kBbKqhDQ6pbctwOBAuHS+uRc
tr2vXNf8xupTcu5r4bBI15O3E07Ei+ogLaiauMfHf5rFaRXryVYsfiHseOzF/n9K
iZ7IIrIvad3LllfDQo7xGaufUdmbO/UOogFOleWfkfHwNXbSdjH7rDC3KmN0d/MY
a+GbeOygAFFsz+RoFEx3sOMZsYkRx8hefk7tZh2tErxd6WsVmrXnO6iXNIwqP3uG
Fep/mjjRBy7Gzj/bzfHw/Tp8ts+goS527yUrtotnmWVA5bZJk04ErMVTh6JTKO+l
fAfpgkseo2MhVvLGdeMqBxLpgJX7U2IBf4HR4zpufdIQsZJ5HrrR9E5DT/j81LI5
pqogr3wyAU0FiueL3fAROlXyMibyFxNImRWOOIUXQGXedQRyXA/tlSM49J7O/Z0+
b0n/tKmjANWiVqIF7pIY1vaaWGF0ukA3HiJwV3BnDtAj+rnepLE2nDAFJWsXhOKq
VrFdlaZ9u9SzBlyBOYVj4seWqVTgcIbkuMI84MOFjW8b7VEBjN0WoCsMhR5r48yS
MCDMZhzeWr9x2wOeRk5QjBQt/UokRjodWBM9UAEF+EyTlBaIPFHP9Y6EprksMOUn
LKy+eeZzxcTrtIXyTxCn5nYPAt/eKtmL5GAVsl91PPeBCJXGON04cNcstqbhp17g
HwL6WZi2dsVycaH4qkfcslOyZ3xOtonTQB+cmFwecQB84b1XgNQ0OkDNNfkO0Mfr
m/IJkKjVgyMD6n5JbtCS9/1Qml+1LiPCbEzfMAQYJQc=
`protect END_PROTECTED
