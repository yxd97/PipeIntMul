`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6M0YTIDKk8GwiHWK/IFMAoDn15omhR70Qs5owIJCB3h2+fRc6cN8TxsxtWWvXTGj
6bbWdu1msTfq1+m9PTudY89ZY+n4BVS0WqKw1BAxkfidpp/iK6vDpg5dgwhvZXCQ
5XC2ZF7lmVW0ZfLwZUYah2dRArPZ+aFq0ruKW1cYwLlQbo6PTwDztTH7s1gTovcu
iZtQAnYQ8SBMqtD6fujXT4AK/rhYmnRpVVbPfuUdasO5iq5wiwhRp30i+aWgmNa6
1Q3fWvQ/Y/gHgcXQcNmeZw==
`protect END_PROTECTED
