`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpbXeZURLQ7kS4ZKRGVpjZv/6UOc1MYQBijD0nr/5bLdt8pM/Ml5MKOWaC4CIdos
y/QpUB0nr47dBkvA5sd5sWEgbTshRf65qvrWDUkpyIs1FmrqMTYJ8EjIVOBigi2i
aCtTqCJ2n/xZx/Nyv7YuAwtpCCR4swDjS+oA6qBvNOHAKTbEaGfeQJqXG10j5WRY
Lh2q1EF8enPygDBmR+lzF98S70StZ7urbT8TCCJ+/EIdEtimct+fJG8E7O1c/Kr8
rYAiBsfEN77asE4ZJKWyZRjM4sTx/dVHJYAjw0kKnzqF7Ollmz8YXJFkR/8tBYmL
uz1j6G8OVtLPgN/kEZLGbvb/EMXwh81z4/CChoGJ3chTwCFTiDckgM/ZCuZ344bh
qG9jCzeXWQksJme9mCxtk6LwR9cBwfN4nS704FzHUXNirPsO+mgu55MdGCKElU+8
5e37PuAzjuvnJOth8+55724hq/C8orTDuJLgIdtBGWDFVaT0Hj2mfpXMz0MQocf3
FiPqo7u3sCVwB5O1ZU2thA==
`protect END_PROTECTED
