`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CKcAY9Kq8fd5pU0KygEbeLzUpiNguv4ggq5/6ScSGsA71LG4O5b/EidyyeK8qUT2
fw50B9nG6QpCwYGMHCwSH4yhIP0VziP/DQy5KH0PGQRBa38AQFjVncMX5nXsIwG/
JmxRW8hoSilrtc7GbT5NPb9S7PV3igxHY1sFbqYhvEyR37cyzb81VVllLBHKPn60
mVNAocOPyrIFIgxVjHd/gCjzYLG2LflA7XSfliqnuu5D7H/R2rYjv6OvZbXX+ibM
Ja259+jSdn36N3UofeljrFtuGwFI1XWWXpg+j+Bks/D0qI3IEm12XvAfMn1hAcXG
4UX0F10ukOrsx4MRNYqybWfamvbvyXNDukLqlBV00N+ePI6kIDzgbYbnyEmlifxe
INtUEf1Kk98NHbuG2Fst2GP+wIlmtKsRwTni/qp7TZeSfkpT4NJcENLiFl4AMh9m
YCY+e4+2yaYb2wQAJ4lnBPKzTvGdVWoi/MUarypglbF/fpz5ATVY36+mebIcVvgE
e9kx+J/MMqbARiOlXLTIFcJQ2chCc8FSGeSAfK3wTE+i26237ewr1y+gXiRB7fik
eWyaIq/hBvDV3A+SaibBv5RmmXR8p0lqthexrp3p/Y8JNi6h9p6PJhQZeuP2vkSZ
jMQKI9BYcx5zErJm2GkrPrl5Ni24hbP+Q3LbN7TF7Bn0T7FkazupV+LYSuJGFulN
hT+2Rl86QCel7YeA/3eVLsnhOtagsRdyePqszZQyxi9rywZkDf0HvCt965SM4J6X
1rYBkwkWhtQswu0iWsrL+kixdVFwgTzTCPaKtYrossoN1REBCS6xxly1TyrFXskN
E7UbpVs94pNrVY41yU//8EkQD2s+R0uqxklQsPVUVVSOn28ziMN+z1Cqzlqlr4tM
sb0gpjcVcI7OdP+56VVOVsA+ev+pbvnqktcolVnSKRe1AbXxqX8sEF8cTRs44J35
4DEidHHMNB3BaULKIn9hVuESxT5DfkJGuLh2WvzKjzbF8ZN5OX5jE1cLVxEhuXpy
ZhitCKJPWysHuygfZa7RvKpQD3Hxri+H4CK+JdhPrN6jRfBP01rAmImqR8SNn/Ts
9ky4YaB8fXkmq7cDnRjak71itW4X1vi32NrBdw3VwvBRSmq4nK+5XFHAPtcxco+a
70e1FTDsv5sHrxIxfsITau8zHMk/yD422PV/fcb7lAJqeaNlJuhjLfTaRWP250+m
7vQ3uV1sQQFFtLAb8OLCSQgfuTClvZbM5z5EvZ74uTZrMj5bBPDLEZ75i3wmpkmQ
m9JdgeBx1/0PZzNaagp4gxQycyQqCWrhBlmDyPWd+N8w3Hgb2YtDxuklAdIPHXtf
vB2hRQnAMTq5efeReJzNSTJq/fnjnyjXkJBmEM6lwmILxbJlybUfZmFtWuUOWJqj
KvY/afRv/pZCzYsXoaHHjoMxpdofL2Nx6jbPEfSV2qXMBfPV5152L4VdBED3Z8f1
bYubEFrvKSIYqlvqsRcleQPF/5v7SDJod7flFcKUafd657pw37nG90OygftIYj1K
CO0WJVCm08OFdxYqSY8oR//kARt9Cy4BoP4SUBHBAwM=
`protect END_PROTECTED
