`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50kVxr6L67bTH2pCLADQkve83hU7QejQ8F5nCaj63PePN2Q3uzpnbUgUYNMwRIGy
aEUzB3OSQxDC08+/EdkZ7ViFS5M+QNADuvn6L2IDObVlVfV/Cio9iRc+kmxIz5SI
lOKxmjLWXgSY/iOZaloCuXkiubH6DQ1IBcEygIFWjPM1zbOxoUNSZOd2QganVEF2
KibPUjM/2BwjMor0rEVyKvh/cP4u3HoE+Ox3ovlsXH3hxHy/t6vox1UcRJcKy7o1
tPkSf+hLyR8Art7FjRhz/SYqXpu7fBKpNKygVzatge/U1t/7OpA9RhYtrDjzAkrL
PuHQg5TqPHYDkfZ9wIFIJZx1O7EunmrptIcBuhd3XyLoeoqriP5EUmtVdyyE7vUN
FbwRbrj7QgJfm2VjTSB+MgqSDHQvXj3p7RC+hj6Ydsgs+L0I542ibg7si4FxEMxD
Wjcl8W+VWHisen5RDYL4nRwJHuefqR6zc+8n9XbzR4bC3caluH2OCBuG/eobY8bc
etZPsJyOplkbGWKI5YGka9RCDKyO8t5t1t+V2k7L+QmRnn0/5bmYPWEMsPhnTNn7
eOSOodUtzJRu+gzhzcX0zpdeOeV4CTOT5lhkmSaZHSp/9SDEIEhNmmXz1jYw9txL
Z8zsYTjt1XLc6NdvUIYlKndILA/KoxckEw/kHx7kEk/N8h+NiGvpZgy2sfRV9i7r
`protect END_PROTECTED
