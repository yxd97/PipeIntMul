`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/tDsshIK3NtRbk3AQKoytjtTwO9+NMHQ2w0w2nz+dRZ2bXlxY6RBJ0L3orahf1gF
6C43PVIs0Qm2J2XvIoBxjK4JuCoxOA4SL940raPRkf3WAsV1cy5A/YcRoX70HHs6
PtzTrxS6kR81oRfLPRXFIBubk5o8ZNapoQA8SW+6Nvqn8ryW0+ftMLAt1+vyInDR
HERAA1Lx7j0uaeOnNmBVq9kF6TBlWsYFSg16kO4AMRVZx1Mpl23KqPxxLOKQYDKQ
kS1znYqF8c3hnKZmaHoMSO6bcoWM7Q6zf9cgAa6u8YyJvAKAYn9NqOwx6djETZeP
oCEiz6hpaWzsGmY22Z4kmNIxoxyncMAZai/ITQr2u+aruhwfRLQYTLiGwAhH9dC7
h/MzrXj1VID1Hu/6+FHDYMdXDt8seNhuIibbrcn+8Sc=
`protect END_PROTECTED
