`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eR954ZpJliIbCryT7Sy/7hqkVLXQVYhcbznu0u3Fw0gnlcNjL8MbO2e/p3YA5unJ
1mAkz3uFKejT5xnc59ll+tWLOSyNaE0S2EP8ejF0fDNM/mnrxFpLmpK8D1L+xm5f
f0wwEPtu5iVvGc1wKl1JPDTZYc5F5IX9bSpRaQeK8w77tj/o8tsXcyXIERe67ORY
IvUqzzLvjYL9FqmHH5mFoWpIZZTxwh9IImQJw75UT04665UWOBWHhgxZkmtxt+9a
3TjE+VMQHNRg7UUQn4SvIO2SW41I/ohEQNk0sdhsH/kO+OjFbVJVynXZdGQ/HrEJ
+sBK+vv0Alpbg66oZGnK3le1iMo6yGrm8hGVCmZae3jxIP8OebbS7i0czqS+XA9b
ZL44kk20xJe2IEGZV44opg9Fu9kREZtaC66u9pPABSm047LLMw32mhSNyC4kMJYs
re9XvAJMi5+iFKmBpAg7ubKHnOh+SZ7SwGQ+8QXqwdaOpMhfWqRunKq8y4p0X7Vn
Xe6sLM6W6YvmkSPVr8C4cOuLFtKd2plU2blEApbJDI0S8It8LMVJX08LemT9Zq6f
93gPuo3QlgkTnX0e5G+3hU4Dr+uUfbYFyJ4v1USngaMUnqmB9SNsUJDdJTWAg5uP
8HPO0ZD6HFlVfgiXxTOZIQ2aNL5xygeR/Vv4L33sy9Y+nVbs+qh3E2Iuubc4H0h5
1x5wDmCO+yr431Xsq3emloswhy4Kr+/zDHNAtidK+YKzXApyaCIc7wyyCmraxFRk
`protect END_PROTECTED
