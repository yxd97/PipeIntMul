`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTKCLN/3btA1KGpXKKY6xM/9daCJEmBYClYgmfC/JB2Jal7yA7RKLRIpU0I+Baw2
PxrvpF0SKvs4oYBpBg0vNRe8yji1TiEGzSMbefDVu34cGtM8cpzIRzzjtD2q4fLy
IRfAdE5RN32vmqHHDgKbycn3KB0XaY/OFPjHMsjywtHR0g8WOwLUtocIoRbkohc5
eR4iD0p9Fo2BxfAysEw+GzqSRAP8dj1CqdADvwJnl0xWdAYNrYUSz40paVP8Nu6c
B/T456lsWevSzZJmbP9AUP6lePjuWQU2XkzH7QDV2d1AcPu2+bLQo/mgxD+qsu7F
XLRhEuxg81bcF1pWK0Wj9RlSS7QWZLR+S8l1wbHPRinsCszdkGqUbDrXRJozfVbi
kZNB1QwgDjT1XQbpHXaAgri0VqKebBmBvAYvubia87ogpjdu8xZTqpVxIPdXD5fr
iX9vccMhcbj9i27EG1sNo5geZdal6ejOVsjP72LG3NPVTb8QPxl1uUzHNd1bSSey
`protect END_PROTECTED
