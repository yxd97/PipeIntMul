`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1gcM7X3eYTbOa3I4jghrESU/hEbYYR19MlhmwlTRkdsHbQRIfRhyhzbU1iBG3lX6
vtm94l4P6ZwIIdycaneledjiBjmvEH+ZeUpOni9uFd9L7hnKVc+zLaUQ44cs6GYR
lzcJR9/7COZSN/exW1Xecux0tFaFXhs4VK1d02oz87NoWD3LRLq+YMnbY76fhgpQ
XhUn2Tv7+FwHDWJ1KqvNzha41S/vyU4Ed5+W5J8OMSsBJNNhdPPyLpSnc2sVSeD5
d73mimzPrKCG6MKDSYj5oFOMd4EO6JB9lPk5ZEw2JYzBWnB98Cv4yG1d/+APpgns
QzNZ6Fi8Xfo9ZtQiie2o19G74Q8Onj72+Ig1CIy33xQRSylZyeqOdvjkMKHD9mrO
nhh+bEZWyI1YYf9sZ3kl/qkCTrj1T29KfTB8WtB0eqDLUt+KvoXnhdNUMrnTkbFM
UI6FDzpqn7dRAG6imaDxfZH0Pf2sS7orBOFG2C0YjBZstAqqMG3Uyx626sA+Bqxg
5XtVyef4MrglxCufNHDyO6x3o+6+2qwShZRBr6fpG1VvkvwrzLiVj0odOvdCPEw/
C23xRkVpC/wEZ5fehGu88Q==
`protect END_PROTECTED
