`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RlCViPMycZ6gfbhfc2RnOmHRLmfvzZ6DBq9DTX3+jknvIVuoJtxZoT19oFwDRdqr
FU6X0aN96gkKJ1G2LAlVpH8044dofX9rA9mWXNEQJDtzli//nZVjz15dW93zL6PS
tLWNQoaAKdTD7UrfiFYi6bUCKDmKlpn+hE+oY2wQz0JYeHEofMTA92aq04/VzwVV
F1uIj3XJnYsXA/unIwy59+qaeyXale+qFxsiidD9tx5dGbnAAvToJNdYorcZpyJk
UVmVbj9VMLGTdLVzMI1j0TqfycnPPSwq82hIYc1e/OFpY4GUkLDFaGR6OnlN8L/f
YSEiiJd2M6Royp+gu49O8fDynzUNwH8qZWltSo49hkHCaON6mxSxpttN2mLkytx/
r5hsNpPzUbNZYYYSFMtw2Q==
`protect END_PROTECTED
