`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KEnW4lJRmXnVPsuDPEYRw7TRKWsOs+aZMJjPCwkK1lUjEr3uDlRSFFP9RrOMrZcv
Ed2QbeEMhkgaBOlr3bMpAblZeHeF5Fg2cSDU+JPsgwBfCFcokoew0zA5cgkJk51U
A6//ACGYtMANz5XPhQhVWt85PgCdo9dFs8PXmlfFCWOMGcqHCdKr/SLGBp91jwjV
mWSuooXCwJMzNIjh6Buaqf8L366wTf2nVSfMW2hkJSOVMjASdWcEf1Z2G0rQhn1C
JYpQFyc8pw32dzec2cXfpxbHKJT07zluQrrms1gOZQrRrQSlnGdDDJ8I+npRvBbD
Cg8kfrYZOOFTviea7QENs6Lh5/J0tQWC9oQsK99VKXXo2hjNLRIlBOtjeb0N/7ds
484CYTHqfJThiKPbQfvKrapX2kAiOLN65nP8mRPurFl+DVNzaStUrTXRxcbb+R4O
CmQtDWfYb/s1KFBOZS2yJhtU8oATBKi8wZnKEnFDMiuJX7lawkFx+26SD9Rbtu29
FaUjs2C/AWFO+UdXry2RTxkTFGpozcAqqtFTGq3CHdSXUGD2eXk62tEGtkQnZY72
i3po2Esih61KPUujiDrQETB4GebKYwp50JKrZbHPw/1QAs5wmKjwyNz2MXJzTjXo
XOjDccGFvO0hBh8Fz0EQ+h/VIz4C4mGRDdy64Mtmr7oIPj8Ag3Z5GKWfozIb7BGE
`protect END_PROTECTED
