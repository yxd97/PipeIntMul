`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wlb1FZRkTPhRC8RJc2glVHdmrEfN4WM+ZMOUgQgbO6fULG1SQUavjS4Jmi5cS9D5
huKUFCp8q3A3A0MhjfW6pPGTCC2kY6uWXWk9V5B/ue6XEF+YdvNSepJEybFPQOxW
oS0tYmApDfdnHkgZJ2r2uMjMNT8/WD9sxukl7jdBcA0q0wRSgmaGpVtO7SS8ovK0
tBVtIPG5WuSp9sm1HrlnsGNSIXSx0IUsmqOs9KA6qB8xEYhoIZ3Hr+FHReB1uiPv
gdSQ7JRSkT9mVun8FpgHtqJhphabyLiqjh8xx5f+lzpKH7qZBGehR39Rs48KHxs7
0PHWefoyjJZ26g0SQKv9iOx3sH5Txjl7mwVQgSEeFp5S/Mzdr8jRk8PPuCGykk8J
gSSagdprOam8Tln7tAUmdgF5+1Q3kggAWgjXLYfS9LzLFzSSisKqRJdFXO5xjVr0
RFCVI9wJUcDLs4WE7UaY6TfdIkK3AF10X5IOUlRtvYM=
`protect END_PROTECTED
