`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzJz8j9zcTzYQVOtbOGVtHOgY6w2giq7JOKeKoZPMy11n0gVUIDbJBm2tTpAC9yg
gCAUGDaEzLau0H38RbsubVGPDbBte9dgbW4U60Xn6tznFQ2isEJSSGVi6Bk0PXra
aU5BgWT3dJ60XzYwQ3oO5BCaE5R7SZJAmSkYIkVwepogMzJ19rFi/WYdlo13dC2E
6IH1Sko5k1BK0U+oBropVOUPlN3AKHghQrcLIvW/7lfHpvkkex3fDM8UtHY8pgPv
sDIHrqgGBpnFhIeHDmIFQeP/dt0g2fyufGd5es+OZPLVInm8MX/HSFeMyODOWUTg
GdbmR2Wp4PEy3br9WVKhcBWc3L9/hIK/Bj4DR//0aqhE2H7dTnvH9j/H/flQVGkl
k+NZqrtolIE3KWC3V257or8RlPbpOW8/7IW/zQ7gHnApmWAaxdLF32U/jHKM1hTB
OxeCT0daXbBxA07p2R/6bl711g3aErnLl6pTje+NL7aJO+BJRtpeXCLYqSlIZMkY
demxkf1naAto4q4uS2cWCR2AfAMPtIX0PyY3ojcO6eo=
`protect END_PROTECTED
