`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NwsOSGTX+c822HspFJMcfoNeS8OZKSXCWOTeEd9XWYpseTAsFOvOd3DzOZFBmNkM
OVENG4nwX2N6G9UVcEZbWCPWe2/2O+85J9GrWtXA3PZPUojxdQLI4I7DYC3Hul44
5CBguQ1cQulAQhSuGB8GhmPCTtgU3zJo8W7c7io25PHhuzPQI2Pn3Nw11HLd2Qkw
X4w+GG5umNfjI28exyKueMPG0DdYQHNcdvCJ9rgODwnUK0XoYUFHMF1GEDvlqGvj
QdakKsy1qgcwz3YzWC9PXKhhzWkUF4f+R7j6sy+OYwwVedtv8d3B1ObB5ZUBFv2J
0XzpVrTRtwDSDXPUroy9ZATeroRIsm1UXVEDbMdIdmKaGpy0wioEGFxDQeyHJMpy
T2V5sWujzndESA75AlT5QoHdLpz0AWII6Pl/Bxb0Z5cIIQyf6M67fTmKQ/wzu/ON
vh5mAkG4LcDvRsGuZsmd2KjB94zdJ70qgjZ4Z6HHky4t53D9CpM3z810gOudvFci
IKYyQ0j/tQWoUYzamIfk5BEuy2Qtmv4IlMdcCGkvpmvtOMxbO/GDHxrSn4rcSbuf
DqA/Tx1onBR2lnpmj7drXWLbdLH/4kiRcEEMSnzn5tM6BQdss23QYrQV3+Hla9xQ
rkA/qb2PHr1XT6cmGmPiisws9ZnPIMEgKV8Nwe+U81XbzlqXzCoHQDxOi4NCglXB
`protect END_PROTECTED
