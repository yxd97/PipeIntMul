`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h+GV9ThvwOWTXR1QGgZ6epIKSBWBZ9Ve/sc6Yels7kMLojy15WV+xnFYJJMWR//N
xMG+hJZax+nHY/aaxCfoj7ODCbEdVoRmHxJk9/cj70hCspF3V/tcAhSRt0oMUnOA
V7jB8cJcGiquCpb520VNcPkqEh0MLEe1pBwVpvqrW1AfxGtMGN3moYn6Ii1YEyF1
TzqQ/hjTC/VemlcUvYGTIDZQWAQEPAMNqAt0yQ7Ixl6OqdmY/pK8vx//jm4xTMtV
`protect END_PROTECTED
