`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xxUM7ueyvryuLEQ+eCbo4dYcellSanYl4WVPqc/MI2JUznJ3MkYVDPWsAp+tJ4BM
KUb952wZS2Ys0CwL/8+Uczn0Tv/lzLpwhSxE+gFai1IRqmOH58i7a39Miuq9KrGy
9rP1N6+Deato8UKbnwlLHWd/rUau3WE3RHYr4ZznoUIyoSVHDI08mM34A3Ur9UO/
Y7EhHSpbtqJ4awORGdlg9lGH22ggjOQxMnkMPn3hQ73AI8BMOIsnPghicztkge0i
4ml5cs3fO3MEX5ZWX4Gm7ZjaeLj9I8bp8d3Bhfau1u0mgI5fjDnOJcK45+9cV0Uw
+g8/ybjS8tlcL6AqpReT6izmMXv4RfPDdw8K6B4Wk2SUsKwJMkhH1bHnrUFqy1tx
nuS2DHRy2tGqG2IcCejIseXv8C92Bk+SN1a3jsC4UAS8k+94ossTZnKpplXL9SHq
nKtvZSmnvbWZWk6xa86v8HIgUkaWOrNv7+BGr2pbYodfDR6j//w1NxulKvpmVeY3
rJXQEebxLj73b89ujT9c0SKSaZtVWPStuZfdDwactKvL1ieRUYehKecq7wMA6Ccq
6p1FVU1h+PfeFMWfHzRmaegEBRucNOp7FQUh+342ltozkJ/cx+VHl+rmRyeUwj4C
Im37Ddhqxtr/U/S7/TyB61KzEP6nFZqNQo91Wp6Wt4jRIOKoofWBNiiP1st78Ctl
o2xfPGOJljJ0YqnUYNPICy2A91DvlhYLYRhYyibLdUVb6D9+sV32HDHTDi+qQEBP
r4aJj5SCJoiBhsFnTnUa5/NpbMs2PYneC3CXubEYkms/lU+/0gDVTLQ9UxjwYkoo
nCpb1/iUYtmfS0Q0bj0UK25gjZnKfVYUpA5cpvu63nykT/4/bNnTLXN8SOg1AOjY
WoVA0oCEcjLcwxLTP3G4tzIfAX91v2LMsGTI5SDML0jjVm6zO9+UMp9uG9k9t3tt
0qnAOhsY7cOypimIRWTWS/0cFL9hhmQ+GknbImanTvvCXbhkUFKvNPTYee8RXKtp
Ap0/CRcL3RLz52LolmlMPu3Unm8T6sFCqPe/QxsawzjoUjRNKmBMIMg2u+9nw0Vp
BtwEelVz7SKHYwJFZUqkGwYdpNhJbc2alAXcMHFMsHV8AkGQ8/1jTFWfSRHX6Uxj
r2khS+De3Xr9QZC4/rvvYEeBrnavzzCTmMxYb9wwug1GtE1W5tjQ9fSrGENlN2pa
+Cp9iN5OOX8gI4oq/TvUxVPB+ETMI72wX8mlWe8ExKqJrsL7vFfCLJZ6YgzVrrXg
aNTI7E2O79qfmg11pu/MZF1YdfADyrZn0CiDsv7isxWVQJJ+i2Fpdot+KgRHSSuk
qGCsFWHRjTCSMsAO2KeUOnOVT+v1yCjInutKbQxDkoNbwrZlribxLzy24SptmLil
K+s/nHCBOLRzPR+OM6khbX1xc3XatkbfWN3Ri6PkeQQevNl50LRqp8nZShhG4318
px3C7DXbt37VjMr8bKldP0JDLH3CeqzMWst2WSRu2wMD1ArTxLORFRiVl2TF7BAy
XVMwLOw8xtaXm/QF7sK2DkxhtGYRse4pgB96ypKWHT0L8+D2JQ1IJDReQcXZ2Cjx
Q51jkjc/5m/gazNuuLibPtQjWsFGd/yI2epV7sdFHGABHZATwVlgGqd2eAQz4WIC
0thzI+vmkiF2cLyQE0bOlJjOVtg6FiwDa8kRRRjRPjjxtQ9FGj7Oto3YebiEUjLQ
bGco54cFpRq9vExbnqCl5//HLRUZe/lRqpDxRaXuhuvt/+EEg9A4SxRcSMRosc3B
`protect END_PROTECTED
