`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P2AmNqrOatHBmfY7PtAMLbOzRuF84fpI5Sg4VcOf0OYUEA3tKqLd60HfyishglHn
FQTjaZajvpf9w1JAwvmybFtTjpKWcLK7UYw52hnOoEOswioWWh0nR/VE/FM0B0KU
D50kQu1inyuX7taRt7McizoHHif2cZ/U1ccrHcQ94fXxFZSSOZnzUn6FWdVo32JC
PVhIPIpM5sw/hlIIS340BiCDA+jAvIrnhrqijph7/L0D7qpG8x5QjYRkuIX/dLHD
q/d1wduuisryOZCmMJZxTDeZcRU9d2W3k+MZmqxffgoQ8sPZvCYv94HG8+ZATnrI
01tikzuUHEDB834Bq2vAvcoTeV+F78pquEn3whEfJH/IjZ/tJYqNzysw0UePqeg9
vKUufIt4kVF8F2nHlIJ8hdxub3rNX2ZjuyHL9Sizn0uLsbXSfI7Qt4pCbZLOaf4l
pIu4iFt0FNft40d6wXKPLDPlQmVQ4PNsvmzq+Kf3wYREqMtnZi6JEyH+y0VWVfeO
YnCYVaW6aI8HF1GJ60YyKQVgH491N93AL8qbBLckhz9BWvWl9Ql8PN35FasvvDaG
9I13UsVW4FNLbHp8WADS3A==
`protect END_PROTECTED
