`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
60te191/gAyIojO65PpEH16ZKd6vENYfIbASkPwJLGYXsSS5DzBLUpEYoo9NJBYn
SXZUsQM9SZjdOOF/IRUGnwMf6AhFRk3Mqh+6OyE0LhO55HZGBGhMV2UeGHZLukYv
501rVrGXRr3PdOHukyCRSHH0UpJ3eAB5OLUybblj9sQ9htboe/4zJ/uRfDIZ/Jv2
t+K33xJhZl6bSjIE88t1JZYrjayR9GcCu7dc/nbG2uaFg8lHBn/fbnNV6y1+Rccn
wGav9itJYEyWdz9yyw2VNNlvhir5XSiOhIF8bilzA9dpQMUQ0155eorDL/byCa2y
Gtq3xggqDM6fHdGUt5ZcUCtX6tg45CGRQvknFKlnyUY5K54akZ7NGDeJXGwCJ+Ub
vjiDfDoaiUw9ACWrg5v7tuBhcVuKw0bMMhHwaEyROlI=
`protect END_PROTECTED
