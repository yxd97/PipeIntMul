`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OdRKN74+Gz1QS7rQlbcbFT6P9dIlGAxcW80rzX+HxCg9oUgCPVVB0ETH3fTxId4a
9YpmReAYJipBSimbSIDsuxwdC6k0nYJ0luJCq5pUYOBzT393fY5qbAOgy8jYlf6M
fP99KrK6aLrX0j0NF4UB3RXqh3plPJinJZ7rCAlEW0/rIncB5a4PJxr0MWXUtovg
f4vg1+MABSbn0bz+LjQRnX+GWJXBF55M1+y6Kgk2yCg5Z6DqfJgevP5/aiQA7v6c
ljANTZMDi3Yw3ewiYeRYlg==
`protect END_PROTECTED
