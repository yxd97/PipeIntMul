`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgrVn3fPKtgQMVq2K5T7WhNhqqzahaqETg051Zmy2QB3QpBe5hWMALK9nU6Ho4iR
le0Eo4WxFoKKlNS5ArJdqXV7Dv8mJY7IHc4Ok43i7Rf3LdsYiXSBH2gnbNqvz4KB
BUCbKPGkajOa6p+xyiahYIiBVQaSx0Rl4BnhhTE2huDgAT4TmyYTPRTHF4xTF5uB
0ZfQNRjXn+uB6LQBf0eFI+nS8AMf8T0PBta6QijQuQXuHDlAX5FByx+QJlF0Hf3+
FWA7IMvSz+nloVkPVxd5uaPfUJKPiG3TITVOuS6Qk3Rbhjzl+bQ9TrpskvsPSzti
OsQludQ9O5zfOoebMG2N4L+pp+BcvVN1yckczEDaP1mYJ0Qx03oqJey4iv4wLWwo
4KvElBdfb6lEu/Q6QkarmaBF//9Ys2jC1SJ8S4PdbJeQcRYGqavMdZIQoB2q8r+v
9ks275fUT7vokGQtn9llTfU+KLcozEeG4rbcT92+JN2XO14YKSPqLyiBbZvQQx3Z
qF2Bbebjm2XD/X+cRILBQLxY+ohNcU9kfYAUtuLGQLlWH/Ts3cNn3Jj+cA/33ZSC
vOHs5pYaqKFfqJ0e8WCoqy65doRnW7ACyZeI+cRlomyI/HrcWBNLiGzPRhcUZ3UE
FUXb3QyAdT4Z99G1xl7t+qOLuH5IGZ9uAOmKKkaTPxEyBrOj/xQdgJNlM84o3j/I
JiGCqdRU9gDCuSRC389q2xxpuB3kkA0AKanOLMZ6FoTT0LaQdfG02XVxAz5IRCTq
ZqdKrglUUOidgspr+mYZ8a7E6pshBFdWyYtbs2wEmy2NNpCVtndVvV4gilya1mIl
Ujz4NjdI+2EQsYNlrsxQhWV7gG9RMgCCLmg5eS/fp/aVUKNMGGbWS9sphIyfOgr4
gIY9WUvXzsadefTetKayNPP0hjdVsTHdJ03v1Gyr9/gcdXHaT9oIVM3WN3VTOCKE
UlmH1jcRr7+Zvz03Fe+RS7xIhtDTRh2NHQd58/2b3aZ6dvMcmwFCsZVOzuT7XbF+
rUrMm5kdFGSr2iwGsRDWt9+Pk7Da7CFjdrOqfF6H1zR7vYPBBLULYIl7ub18oJqf
DdgKCNEsKvVebmljVUOI+qGZWeMT4WlIpM0cK8H0RX+Z5gCVs/QpM+S6ox9GwepT
NyCWONVczvmZuilQwpiGjtIiJPRmykpvs+opMZuc40jBuWIMow46+BFe6Cy7kw1x
Vs0svp6YEbShQ9YFHAn3E5ubr6qzeTLt4wyvVpEaf+JIOPLE+3xjGI1cZNX+xfxS
u/cIITqbLoL/jpzonEIfgHx/lQaIfsCCvLas0XrQqPvs8KGFr2jmLua2Hzl5UAmv
sXqmiDM5fKWhMUTmuTG3ApIxa8/h02RsF7A+aVDPMqg2xzPttJFjVBKUOuS0X9UP
WnOzDomWdxUSe/9E6+YzTP5jwHU37WUxgp/K/JUuA+mWytKDqBGdtACRSyZvOGsD
l5R8zpcA6VcaueNVL9sLhfX8zX7p9AaisJtoUQEvoXPJeodH51x9661/rpWKJMMR
DAM64lWghZfILNmRfjdpJNwSEWoy7a/p55vnik72oz1pmD6u3PfL0cbgyulVepPV
6NPbH6Utnqfi8Cpf24t3maSo4g03MfVOzVKPN2HxtX7mT0gLzVWc4UbqAD3hyi8d
gEctPdAYU68mqG9PTxIdAQMtD61TYpn4sks0uAzcH/x/2gIGd7Sm4tFju6sBK3Gd
tVw1usT8OjAoWwtOeu/D3noYkUZQjoYVXaoa7sxAcgV5830vBKZ7vcchkl8l5O29
QXkzVxykqO045L9omLNfTVIctjoX47w8t44aJnjlpbTEGNCx/s3eYZoquh76r5JA
azfYouFdvDNYef5bLosZBRMfCP/aYERA31RAYY7ad6jG8mv7vMPtsiq/26MR4JkC
k77iWr1tkauv37gWdrVYh3PiKCr0+HUfaflTKAX2dIOSodAz/G0IOHW96xXyMSLk
iaUM+4w5wAdQPhvJMI9zj4Pk2hD/qlnRNIjtJnHkfDV2PkMDinWAhuyDpOL/qstG
ytdG5VIyUFcp++NTiNSeR36NNmX5TnOW+GNcQm/TldZE+y5Q9UryKrMfoa1B+Tbi
Gmf/b+VaPrnNh9myn6cRfusRinUeIxxfIeQe60ZtOxsLgpndWFgiRmyCJhtaThp3
Jn2EMStKZHZcKbZFL3NuqsWebw1WYmk6QUVox03FxECoTNh0wHk9IGaLxhiF9Rk2
rQdbn4cvIzUo4pN02M00wfJxXttH1C3bubU7s+93cdfKYrOOrSB1SFx9yKN82/9s
UEqgDVxKFiPT+pyWmhbAvCwwhkTTu/P0WEQ8G+N6psgveUIdErkYCO83OWbc5/qa
HrroMgKs+2X3L/I6x/cNRlaVMwPMPEaOQPJ5m4s17bfibFXXPcbAfwC457lXeEkM
mObxyDxzgiKf1d5NkqTkK7YIu8kdglzVJo+Ynf6Pa8E8aQV/kLP0tJMqxttSeecx
R9biwpTXyXBjUuJyFs1buqyQTYR3QSMRCWrnSNSBdiNSJQfrOPdQhWZoHA/P5zUy
nBXNY5IIR8m7rrC7virtU/FT7SefkIIfnr+oN9TZfwl3lUioDLHG7K4adTRazQEC
p5s1FA32KQys+pKezIrgvkUf0NykZWJej6G59I8NiAm3m2FCyKkUdgy3tYTRX/mk
GSswK65W3obsnvk84xtmegVyVFANcdq07aRI5j9eQppkQjRP1FPZWpiwu4ruN0jQ
L1ax6spB8EMuZrYtoFGes/jm/XO7ZM1LoCgMAAsUM+mg5XygHYNvqJ3hBp7UBjYX
UOgHfuS7JeI/C8H6j+D1XeqqAoZOPFJqkc1BvHWS8g0WFCYV1ncYNy9XcHr/YS0M
8Hn5GgKYjmdyWX+NFg26rsgFUfFpF5txbfHyFpipLaI99CqkGA+q83m6+fkpP3i6
wR55VUFfO90Dl4NyXhTpW3J7uzRYtkb+wNeU365saHC/OAhXFf64HAK22ywtWEP9
BN2uuhX2Y6qMKERmSVr8iB6HYMyWLyHLZGMdDLCo7W+HY9nA/SXFDw5LqG5Z0vSM
2t3ujr5DD8C/QesiVnIAlgfd5LLLa8Sy+APP62bVfnIWmAf3fh8XM61LR47AMVXa
AlJAhvzLaoX6a0jrwoFwQIdqOxOsnRuI8j2SfcP384l/XT+3b8HfQZZ5BsRK2bA7
tpIycQvqrPrd9IYrKQ5g5psreNPJHufMuHxR56DTxVQLrBeSANid6idWERp2BtAD
`protect END_PROTECTED
