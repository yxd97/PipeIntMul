`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xTOKdgCsyhWPyT1K8iGlOqYtRxF4rbXy/CX1m2XedYyTPO4msQEV8iC2tKAQtAY1
xXK0423yizSlGghd6pMmxvnUL0CaE31r7ZtfjAb0HRO3SkpKE0zQwT9QAlf7TgIv
RfsiDsk8yeu38q8EWnLXNzuP+ZMauF8Jq6IDckEypnoM88yhqqLABZH0WuOEZM28
CwVB9wcbfxU5mZO3DjKCnDR7oSX0lUZKHojqTHqUa7vm9Zfy8Ss+AG/+zVLCPuL0
tNAABoqqLf8ez/4D5vsui+jmjumdkNDvWzDtsZ0xrjee5C0o9iW24oIGKo++9y6N
x0BGDjZpy9imB5UxEjeM0E8zBAHPnvKXb6zDwOI7532GuZW0bWSpPM3qmZyNSbt2
MvegyQBOq7ypFQU786eTUllTnueVfm0sJSd/3Nhc8XgxuZx+cm6xr7s2NGNxhTzl
1Lp4DpWTGM/XVRlSuQyxqgjp7KY4vWhX+cCIWpd2AmxFjyQJNnhVGB1gN/Ut2djh
GR8MGGrUb7QSH0m/LRW+Fs8pmINa6i+0HGuymbRmXbKSeqUaIyb4cCueANtPzBJx
VCtANsOSVggDCGqD8Tekn7GKeO8lVSWTOXsJw4s0HLAtbhDAnann7aPfuyah/W7a
TKkx0+w3BGboHnBec3axW1tN1NE4Z+Qsxjgu0JpruzKTsn27Mz4xB3WHLFxw8lO6
0JvQMOHnmxdZOStXtEYLj9EQCfIDog3xo8ITVaec6NRP7S2rCdfK35qEhNJd2rlz
XBOJjoenLxh1JGACEm2KwH37K16wCOIV337NN7/h/QsNXcUxiwAzik2GqwW9MNcR
jqYYOm/FHGr7gt2dJZCOn6e/ufeEQTvsMyymC0ipX4pbrhwSFk6jpyCPKWuCeSFz
S8liMyFuANUqM9flxoqlP/sJyCTHTGwWZ8iku1Cs0r7nlkc9KReGIR1WCn0Fv7on
VKQkwKYKWIrUn0+bayDxI+CCTOUjBaqi0XeBNPsM1iAv8Msg9oL7dfI+PDSc4QW4
O2tZ2OnBLx5bSewIbi4wkbMueauS8sjVZ525bLbt3jf7r9n3pJ3NZCU43ih2sYWB
fwNnIf7DIIK/GXodbFPVwUGbpLJp5v1zeCcYmk2Yb/0xhYN40weu1Ew1WQpM/QK6
Y2c9kWbSbiXs29vo2kaOGOWcPX4mj/Xvuu91L4NzVZ8w1WWcpFeXib51nDvbWfJi
WebzN7MgOpJBavX59AiO9TsX5g1DrSn5e43dHwF9rLqlWKUtXVzn3Fz2+rnd2xPR
6R6zmff8N0tpwSWs/fsBCfhoTp+vko2Q6VFrS3NNOpY2Brw5uTML233MjPyOMEGk
tn2RNJLSmZkm7tuSXGQ8dv++IMFq73LaTQ30Z2tDQKZ8sxMN/NISn8MYm3iaDAiy
mSFmlHzbLx3x/lJfKZ7FoorSah7GF55Lu7haSHv4ml02RDjGZiicJMbpxA6NgKnZ
vPgXhgzVSosAFXA2CDSYqUewgtSee8ZhA5mhOt9MNQd4cAVs2On6tE6J/AlqRy+F
gUuaPvTUgQ/TJSON9CXoTvlZ4hO7EJc6K849bWOfoLoBiaoIppYFJxoZO3JvHSrD
4QfHn2r7+UKm16wI1NQ2IIl+ckRoigYR8ZgVFGJ+v9qAPqBdHS63usKOH3QNkyJz
+nt78K3TI3v/oIsP/vL3SvZFMj6YUAXVg4owxlG6I+FpbBhWZsXxBAFQeFiTNyhx
XYNDsmg/K+R91Kv/AEKyBW+er2NqnCL9kOrkLU2B5tdspcH/oOhqP2gRBRX823s/
0/e6dU9I5FDnbJiK03wFWwUKOY1XsZUtRQB3pp25jBunm7UbLOFE3thAAN/HLOyX
YUAL9vTJUvPjFIIktpWNo48jHyp4OuqmCGMpIzf5CWRDOlVz3FErNqRxFKVjJWDO
dsWS0TirMQ0PkSIUWOyPk8nlefz48DGiVpqOvdS1O/gj0dA0ABN3fr5oG7OGrnpR
L8/5SDAjSCfo8biOgFSseXAYEOzDowkC48cB2Itd4r41n8qNmNF/CVumkHYEnZ2s
IHffTnqTtQOYfJ7OfpOEoWUpWbA0ZZhcRTI7gdphCSTGnTmIpam1WBsK/X16nG8n
cTKgvMpe3Lp0fn+QEL1XXAUu1gEhh2zEw8H2N91DQl5RVLH8yWpsKCZFWrRo+ECE
VxRfiuRuvGHIwBbgNNdPcD7i8UeBIGMY86eGJkODuYwtJdMdlFVV2oxBmt7ewSIK
X08lJhLcF0XfP9dM6rTDh5RYw8E74ttO8kzgm2wHG7JI+/RJDq/ATEr9yz/bK+0n
QEKl9D/BkuCRJ7ScNjz3mZYfiMVpIhzIaXX+wVIXuCkkMQXDUq8MrK1Q2GQwu0Lx
TfM85IXLKeEoSAjUq871NxdRyovP3kFYbmqQVe5GstgmqjeQnYaYyFCl4TW/0FdX
sCxJ0ZvoJ6TQmCTVI/oSs3NX+YzsMEh0QAtbHs8HbdDqBhD6S1c3X3zX69CT4j4L
Dpqc4MMksUEE9oBlVzumQ+pLaBjONJTCKcd+PNIfcAaLxXB+MbK/mibYNenwXMNO
azfQAtfaxXOMsO76DnIPxdpS6XoDFp8Laa4ybFCW94XDxsqUoLIGbsSCQ94noS97
aXRcSIAeVXfRcye6jVVCGQREgaauhK4rZ6Tj1CMsEWVyht+imqGxgJyfBwdNe4Y4
ZX4uem/ALHGs9Ft0G4Qx7P2ycYdrEIb0CeMRGDGxXZ2c2ZHNSIM2zZn9wZUfihaZ
BvHDYu02vc+a37BGAVOgwjt0k+U2y0ojV18ll5JAbG3Finx59DoqHhzwYmarNLKX
qMiwDRT51hFC1xtpjWdwwAB3VWgB3UWZJsXscup2qBjxf2AcUXQ5qOU2WtcHKtg+
xj+AS0DUxPFitj3UG2DwbXyXEyGuDDjyfGKp+NXBdcHqamcetG/WhmAtMGn9iUmy
bdG2lc/aAtNK4VkW3oaUBn4xVqxXR+cJyCBjpXEBbsdpC0SQ1lLNe5W4Ugxu9gjW
529KkTdbsMWL6DR5QmGd3OBzI3/SCRzLwsR5GXuGyYyqoWL7SBsryiOBv2bRuxFk
arkGfQN0AERy2Jpjl3krcM5b+b/vVnwzbvxZGYAspLSgb+QzsCw1LnANjkaR8ELb
mQCFB0PJXw22AzriALtyD7dLKAg07K7V9uQjO7YdMA7mARQqurEIlfW28/2h5il2
hdYBNknStH07Oz3H/mR+2xK9U2obtGoM2BqvRfP5vhTdtEuQimSxynQDbghN9tut
iYPH0vwWTwa8gSskUu+TpM0YcxRsSBQYGFyPVLPONyk5LgtinnrG7xeA4eW8swKA
6TFK1e61iIfJZS2nP+UoSozoflpCAZ3K2/v8rrviTdWKtj9jF/d2Zc1M1Cb7UFU1
QcbsA9Oz1u9/tY2YqcN7IMO7V6s94A7hZ5YDAIvKRE5b9r8Mcv7PIS38Y4m3b6pD
orm5zjUyUpC1GZ5DFJQvuJQgYCQ1TB+LoJkqBZ84RyLMdxVwBZPhR5B+jswsDhfY
9TY5g/ZfUikOg9a0Yti91DK0OKPRIW/yXh9YvcgYXFpYKSZP3RznILQsGpaPdj+A
hQdozwKkeoCIgnvxdOkkjftDlGG7CePeIwAHTEkVzHlNlBOT7fSyKxa8XCp6c8dd
B0DHqhcTGMXpnJpfqt7qIpc4VVkm1j/IPY/p9UnZh4aX8jbx5wnlvZyfEHAF3t/u
dNMDheAttOxDTK6JCtcNCNEpSckovYXUL/0pzXsE69/uXIN4dVh2CGFwEr0DMdCK
9XO7hT+cyoPF0bcaO/KwVl7k1Z+2mdpzr84/bsd4vWQPYK6XS6AlZ8X3CB5a06Rg
TiH5jt8YlmIVFejC7wlXN1K2iLphPpCMQDYDVUhkRBUFhpsA9bjltRiX2UgB71YB
Hs60W0jH0TT5fjo9pGk00MUU6RgFzTIWItZZF3g6VrwLF/CbfHR2r12S/ZJBHAg1
+Z/vfcXi1YFjpE/zZcXkwNlLJpTeNQmP+1PExi/RHMcmyhTmOnFbkVPADqpe5BuD
OrqtlDflkCpQsEkrQ8cRaL3CF2Rc8eX9fSbJFut+VuE1VNOPfKIroJTqVdVE+imX
9PjXvUkTGfe/7ViE4tEuqt9PDeXtfYvi4o0P7SiJXbDKXJMe4o0KtnmCHAAVxprM
bK42NLs3j2sodscVOgFLvdsbNmFzkseRnEJdzF7T0DdV6eQ5HzH2a5mdo6Xo65Sl
tmQVjs32tOcKNH0OsvqwayTE1TJImHx/weIdAy/m8OlWPh2zjbWJMFesBV31Bp2m
pTesrKnzsuQ+fTbQrhsQqDxnTOdce6fvj0iiPknyxBOAutfyLzPEORaIiKuMC/KK
VS/DIcvw6I6NBXaeMP62laLhHroi3+b4C7iaY8iwzeuajokNvXd0poj5wKGHrh5d
3gua4rRSlcHvtSZGFBuEXP33PJCqWAPOMJDRoW+Q1G0C9wxQGz4XhuP4Vv7GQNxS
5yoXM5N/RDTIm2/jWBb/pVXD9Ew78U+CK2oMWTzvqTkqdf9AlsWh7HWdvOQtxcJi
HL/Tu89IwfzjAy9SHEdKwLvkf5cb7+p5FVTRIAWcvvC3k9GrPDbFXkh0P/GyPy9V
04tYp3vOJsq2lGoEMt6sjHbF9sTOHLPO36mrK+6UTWxn0/YyC9OSZ1HAq/rLuNXG
qCY9hbZloxakVHTRB7qwGLksMAf0heCYpn2vO9b6XkzvWWJCkQrejTVVT/esqvF7
2M21sJdtws9zTDwfkdWYI6Iz6Kfw0w3mQ6sPmcfpOxRkVQkFmkT9InMJb//NuwAo
0hH5QwZUiJ3+7OEHr4O62ki0CCKq/RwaKyt3+xha5vSN9IeRzSvs4cKDJDnQ1J0R
EzW40683jG3errw4YAEJhMLR/X0kb/HZpOdfsKnlgsuQtC1l9z72VCyJuxde9os0
vpnANKwXmt9x0lbMy3gh1nC4/HzAIeIKxwU+QUI67SGurKw6cejdWOiOq8gLNVZk
VBghpB3VssAaKsqGh5UGVGFOtsYoedUMbAf2OfNsi5cSbmiu2F1AERUHxkpe3sbc
m4+BJkw7k9HfuJXuZ+kg+I2nc+Lw0CGVOZZm9mduRiWvwZoBfkuw52jhLcCvsRYH
/K71ohgMaPPMHpwN2HNwDBeVpFBiLbU02sDS5E9DzUxCz0M6jkTkEJ0hXcZQHP3b
fiN9EJwG6iZypezNdyZItJcvLEhd1DM5vTQtm4A+SM4sL5qFbt2qcYFAqZNr3h/C
AisbkKC0a+9Og9n0a+oKGoOaChbJ8YySl5JqeWvQL0/paDemacXbhRe2JhaJz/o2
l2725JxoBTNz0CL0PkZos8O1Gpbc1kwlD+6/uwU1m0QgvBA+ngMfi4ExbNyxZu0u
ckVbAbK9+IUVmKd3avM08cXbOWIDGQhaWF4hJ1xTosXtzViqXcL8dx+3LtPQGfcq
S9rcorJ6b4XfEfwaQPaAgLj8WWxGG2Awb7tTpmJItsNRVooWxMD2TwWChZhqleH2
ReA3W9v8EQGxDkExIRF1izq5umcLIRhMxejQCXoAoKX3P80EIJNh8UwiphQZEPTp
hg9jlGjsL91jErneC+uPM1I3OVBGafp2sPk2S0rJl9gsehZ25YLm74RUIOdgH28l
CX2Z4w7oEqZSM3lmnhvaBz7j5WGkY9y4GXag4FMj7PXsUZJ/YOK+xV3zu50YZX+Z
`protect END_PROTECTED
