`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QtlOTAI169swoYyVOlx/mMKtYDRLA0ybqsIqG0dseetQxExaVyOhY49ZE7HmAglQ
gqvsjFmB8zGVj4jCJGjsxQYVKmpR8/y/EYTnxklw/bUEr8Kfb3liNZ+40gyyeQP4
N+3aUE8XEqQdaOZsjhEyS/3PXki/7JLUAXWDB0tVa41zKLSUfeQoSofml25PhCnj
ykzZrzv+3xfB4idKxB6RaikGNvqIAzmXS60Os+QZybHCSrhwUR4SvU2G3KgjGoGa
afWrgyZigatN5bwXIx7roA==
`protect END_PROTECTED
