`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IijwHao1bbq8VGOww6Clepx9LhcxtD/0ntnYgZ5oUc+/bDmjiXPyyW/GClXCGlpf
q8qFrVUedkTBsr9CNxkHVZ0Y0uta4bt2Kg8+H8d84n8MsF/a480MdFGL3naIxhaC
GNXZeeEmtoQka26NH0MME4Yj0P9Zqaj9oJBZnEvU2xBXwLDNOr5062ItO+j5V6ab
DxzqJOon8AKMJ3rMOzDl5JGhTLSUjbhaMraMMyoFLMBY1zX5phRT7/I416fJ7s4/
t9Ev7mCqePx4IH6fe+5/YVA9iQ17dgBHBLDFhOY0hFWbuqqF19k2y6IwHWUQVX5A
`protect END_PROTECTED
