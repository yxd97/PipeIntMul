`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V/W1NrGfzjWL1LfwG4a5O+B2+sKqImBfRcMvEI0H0uZ0YKSj9QbsY0L8qjQ8XffP
TJl6f+VtGNQHv6aeEUBsTPFZ5Qu9NCjv9Zh5CSj10YUp+K48AfYPCbe4k+k3JmCp
bjAIzZ0Uvz2gWKb0d/iN3rHHnWmklxSUWqGbqN5QooRa9gJitcylmF8aHz3GM4J0
9BEUOsi2s1+U1og36A7Pfpy6zje1JCBDe1Rbz4NRWVYWZEMZL1RLJwkhtlav3EX4
APj2kh2lrDLiRvNq0okAYTp91YiVOjOTOKKEV0NskSPFI56Fxhxsh2L5vN0a3b8z
RvDqHwqxtxT3e8u5H5wMERT6HYacrpl4398CQMMluAk=
`protect END_PROTECTED
