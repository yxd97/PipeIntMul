`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6kPkdmWGbp2OsQXQ1aodbOIoNAh1Eg9eVUC8W7oX+XOdkwe65iwvifRCyHYzC3A+
haq3Rn0JQ7HYv15uP48EsHo9UtVoD7vFfmC0nvujS9070KKLH5QqGKBLkd7aYPGX
ASWE1v8wxi4dJLgY7ro3eP1aqV0jO1BQDug0YgHqUTqx/kQET1mjurGnyO1GAhCF
NbqC9GT3U6lDpP3PUiJP8n7fyC/L5ktSbs4gCKDLDxLEfBHs3gfhAzYhYUQe2SOT
fx9ko8RT6S6a1f8VWrxqaLPZrsln+/Pw6+3utzYOXs4zBQHM2v6gyDVUn3cpkhNU
`protect END_PROTECTED
