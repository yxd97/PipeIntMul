`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oOrLizGGQlt4/a2OQIK1HJLB0vcI7SkUnOtCBhmwtURGXeGzr+7Q/xpHribr+eJs
fdVYyOoGa9y0Xt4uUMP/CO2u6SUaarkwyJe7xXUo2n2NDPQZEhXuBCFgIN7ZnzxO
hUoLFmWQtxfz4CdxFtArclKu47IpG4PrmfQRuuwmbF3L8ThcbQPGtR2s3KILty77
urSzgjb482MtHn+ZCuBeIZA+CW0NziB4jg1WUA02Gh2Zn8tRumXUsHAexXmwwCN0
2Wli3HacIlcHv7YNYb9OdkFw/Q9rMWerUaCyC4TC63QWK109RZTV/re/x+yMc+ll
5QL8XC1d+XJZQFAlrMl7J/0H+bOdx8obkDjjAwdeTkQ/ObwRyLUNY/eeloG5msSX
avYOC+Y6Z1zuyokp7P+EJE+Dum56y6E8iSlCUsQp8GOY123BENaJ7yfR+/02lwpa
kqpcbx724Shv4f7N2UU9ZNXtmBG4+FevK33Kb9v84X1TJ7h3LNh2E1CWYvGm1oM0
mCAa5EZqeIgl1Fz/XJNjMVJmTWAOurHEIP0hvOCPR7eKZMw6TuCqsuApZ657Sv0C
qradWln6p2iz3c+gPQFK6Lg3M/UmWeuRxfscFM55zUgyZerj/2j67njtzl+mae9a
O5of2PIyt/+27tk6y3qKFQ==
`protect END_PROTECTED
