library verilog;
use verilog.vl_types.all;
entity TIMEGRP is
end TIMEGRP;
