`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p1obqVTSuSXQLK9ixZjAJUa/BAohmnziYlEWBKnUn/VDHkUkNiGthqKuw3oxuNff
BGZsjOBHXuLCzGrYN6yRpc7GwSri0p3hhkA3v/AZnR0Tk7RqaeSxQERsgeUOkTbO
cIalKTRuJ6rmPLWejCaH8Y/FTMVsHs3+px9QQckVWoZUOoLdUnqYGjm60NbjkhZX
dTk2HyfJ/gAuJkKLjj6bObmLqzUMq0nwg3H1u6tnhGa+3DOosmasJiD6kZw+OzSI
ZAIesyB6wdk9NJQcVYeV/hvcIynxUj/c+YJmxo2HfbY=
`protect END_PROTECTED
