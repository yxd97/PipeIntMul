`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dqg4JBPgcSchvHOjUffMMkfidRWcpIFOCwTqlPP4Pkx2tsMHa6haDZCdbZM3GzCf
ws5wWEHD4zb/OAEEXfTygkwMQkTkItdjYA1FEpi1mEtLzkuzTCdnGd3ijfz7sOu4
HNexKtwiLEJaVnHdCqKNssNmNPu2c86owgAoty/0BQmU6abpU2bmiQ7E5jBrRXqX
ULKBUGx3Ljuj9u/KhASLbIY9Y733CDloxzhgOfuhDUfUW5c0hOW/n2Wrk5QuELsV
KLJIZFz0s7MOq1gXArxTKFQnOxwN7jW7hUNTsPTeZ9KHTPj7oMEtom42okKqzhw0
ny+dm6aPkjvsjQEU+/BFn0Xn/ykoVHWcga6/9zoJyJM/FLm2pgEQDxfH04KFc3y/
y5o7UvEHOrN3C6y3Dws0Fi1zvPrEBt3WNuneb5bRhgtkeSTEW/YSJSgI9qW2JrbG
tPvRuQEnIZuREC2s/1ogzMY9ImijlI2LftPsy+ArPfjGxEU83zLHEootj23L7Mf6
rZ8PXTZER/7sVEZSvHemykxk0DgZwMtNAmDc/bL33G90XqWLjR6vMhNX+6l10bdd
2wHYWW/v+gs1TL8DQXwgME8GUDargo4WASWCUDsiH33OS/xeOLRO5w2jhxpAJ1FZ
chmvDjEkjFiHFSFUEkggl2RmnJblGPmHLDWu4L6sXXLh7mjGT3hWfakEURFtGhwa
w/1lvlWq0Y5WDCqBWM3vmj3t2ijqsVV4f8czYvdnCwPPyRDibMji1oqFU3J9KXWo
+3vCX1y2tE0nWG4w0Wcbl6JLb/5CDPEkPkqeEQJl4Tj2WV4pf0UcL9pyrfN3D+2k
ZkcTzuPzLtwR66QyNbqK5k250hxGC0/TvXUqwTA8WAx5r6mZZCMWkcXDy3oRar9b
NjBlap3uPBF4OSDwj845Ke3aVv5x8xQ2fJEUQNjVLqlpm4XmjH4PIkbw6COpEnv+
gVkPHXQ966ygoVBwYwwBOOTPw4aLXtlHDoIecjB908h8iqROqYYtKHjCKVqAIvcT
KxMFcXyoaxUMycHmk9b4mYg5Ww7W8rjoK5MV/ca3KRopNc+CPVYyje7g/HqOtNsK
IL/G6ZqeIyurtw89I1y0dVTfdSbBHMgkQDuPVcWS5xtwacupXe38ji5defjnbCPg
wZIMuGFiOo9Y2LqNDGND3sMUfn2HRvoPqBYdSoE36SWffFFtMmokvQMk0+ZOy6S4
1Eb+0TLYclRoX/kIfaJUXPtjWtHLhmV1asuibeJy2F2OuwRF/g6MDteIuUHMrAaY
uFW/u2Rwg1K6frfH3LfJbdOvTZTkL88yOKHUBuvAWJPRo3EAE+IXDY+fHOa83Ab8
Xj/MN+eGaqQ2ygG/hNDeGF/ZWY1pLQUoQN+as2M7ok1Y+friTrtl1LDwj2AU7fLS
XHQx3Sv/GTNrp8SFOt5MWPNRvVp3wK70L/9v06Q5hAJDIjpnxDNcWjdNwmvxaNiX
y/FMsTHzh13q24ilK3vqZ5XuKpkl7GUltgxszguXrJV+UE1CiVG8//zjGcmX5und
l9r0l6uxcEfnrWSjduJDZ5txemRaj3KdcGCmkAVZcpFZPHq3DllmzBn5vjiolYsr
qCV9mEvLzXLu3oE4DcMZfBr/7PCSI1Q3flIyDnuoLDToHhmSTatwHnrGPZqFavFr
4o7OnWz5B9x0ZkFT4V4XydtZFsJzgKgF0uX1e6SDZ3FXifwNVLl/UmGmgAthmD6x
imIXShpjAexDrhnirGJmuNyISNRX2TXs4t8iY/BeM/ARStQS6MS8plgeG3GfMHN+
NWL2GpoxKxBG/G8QPCKvw1sJCPwzdwn0XPLUS27OgA0na/+1i0zlnS35aX1ehlCS
xrN9IeAJVAsV5If28Kl0VfwuwWhrj8xCy24NsVnXf6IAP/SvhL0TpCPmQpOfxhbi
Oz8Swvh9sWql8ImPzgBlYSPMMvLVYl5fvzn53LKDGbqAtSk+gN5wtl5sT12MsIyN
VbERGsg0+zyIRiTNmy9NzUStRAY06WU1Gh8EBladl5+ndKudjqDLIQgkvGTHaVOk
nyEd3T/AvuvWhYqzjzNqXi9acSARmxzio+cnZb/EyvS17q3COY6R8oguvHAoEY1P
gIMs1zWllfkMk5vVJ/gt2GxpzcwBAKsCWHLtOM4BmEBQ+UG3V3CYbr+rcgNjzcqi
ARC1lt6Ar0h3cYK6JdZ1zB5hUlz7E71jQxAa1cEFK+dFo+mWF0XI01pVPDLJYnS2
EoC4Ha5AnHvbkRkyjJbS2uoXk1q+3p0+iq8Ip8bHI5TZvpK8eAsGMm4E+dxmeyw+
uXLykFK5xfbONC2fQ4yTxANmxnk/2ncku/44Zhjch3Hn09ZeNGL+nrF2Sa6Qs9vD
egNKBaQ/SVhHVzELi2oFJGbjzn2j8hZWe4nckiKjBj+0aLVuXT7UtWvV/HOUXkky
5O65PP7wlfZiO0DYzNu7WwiLMgHAfye6+XysyENEGMe/obZ9xlmgogJWOeaOAlJG
ldOFOc3VoZ12rpHqzkRxc2fZVvOb9JUlRhAGujGr75+usoASwTr66CvSbj5gKTRz
88c14IpFPbVdjxyq7CvTSxYu2yS6ewFFx67TcxxkyfFExYoH6jS+Kr1Al5pERZ7Y
9RCwZVuEynUah455yOrpApm0HGKH6g17QdDjY6JmQwYkn1EsNTDQbFFY0IwddCt6
lDUydstTFiFkYLFMQU3fd5ydVEoy/NgiNHBdNt6KZg7dK/huf8tLwQPcMBTZ67/g
PA3ewwGQ6uDGkV3NMY6n3C4bKG4VcFqmRfbAL3p5BlWRYwAqCvbqxx3ie06kb5py
wnexOuaWx8JSkHf8MEGFEm363vqMh8RWncx87Lz4c6JFQTcHs09GIZhFXg7CoNVd
1L49pQNiTlq6RI1kDN0n+x/Tzp8ikmXSVJXk08yOTvpnKkpxszhrtPPi9ANLXOXV
/zRzK6kfYdNyjt1chLSuOp+3cNRlkiC0F6C5BhZwoXxKSgC/SCscVeHlZAlP40WC
HbLa+u2qE0n924ezpWDMknEk4/LUCB/f3p+ysF3Fpp8YEjVN9Y5knVxPVFGFdSHD
W+VbN9hwh3qLIaQJqMdpxAgGMB2cwCpBC4TxdzkDYMHRhQfwCPOcNnPspxMVmSmt
Sb0Xw23oozxZlTuQSjoBHHv4dPNNsAbw2qJB7AGVVTkPtNCQy8val8Dk49K7rEPc
lFNrgMi8uVWNM7dE441ujDVEuovzW3ie6flg9vwGu6Ha/Kqr0GIFdjwmtVDeAAm2
brIFj3/gVpbjm1nipAfULGg5sn6T5U6+i22xXPCWrLeFwO1lmmSGH4BfLBzXJZu+
EpY96Do1+QxzGeRgkgYm3EdByOeQJ+QgJ/syNAW/5VjeRoujRK8Q5leGXME0a/hY
sYXx6/GLj27umuD0WJUhoml+fWRnnGpKIenYgfQC43o+ZlkRwIgW0xAw2Y+BjOJy
1m1ZmkScH5/Qc5GE4iEfq1mRCkz2UaAW/Qktffswh92TbTZKZ+rlyJhy3PqZe+eo
hNYh2IZtOrjGjU9hH6ONTGmhJbakLdR/kpBqgoeA8PsnnB0FD/8amWa1oGWi5gbS
Rmk6hY8Sjl/oPq4dIo7v9qhDsZWSPjcbFUO1QJKHsnKxvCdqab77VeuvkKb2kpXU
4NClf0bIASPa24jEYwFYow==
`protect END_PROTECTED
