`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a4WDbP7JgWgEK28l7FxeCMmcgf7BaP37g5rh97QZITgSAztAMjFji0UHw0UZIZFr
6Ckb6TLEiOWroEjfsOTCjGwVF6dcmzwfzMf7FpEeFSF8M3wruj15arsD+LpJnx6f
3UW5Khrcb5sSBj0qWBFs8TEGYSwZUouRHpBGHTDWY17D4cuKbqRJ3My7n5Quq1/Q
kkBg4/26G0pzaN5i3vqI2e68r1rYk/G61QvwQDSmz6hn/sC/8bP8NOrXhCwkAJ0v
OVjqLnXzLnATruYpO7nc+m44XPURnfX7HHfXst/PBuvgvMnBe96snlpFbEIz7xrb
sOZxpBNo8z5mYD1RM9Hz6jef9Cr7d+UIyv6S+otMLJVKDCQhn5t7Q67ifiTybGqT
p1D02fkq+iGy7J4lOu2RiJCCQEPm94k0hEQT+cb20bYLmSfNj+JnsPDSe0fyjni4
`protect END_PROTECTED
