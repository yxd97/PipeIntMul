`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1JRMa+MeyFMnhQSeKR5N5E5Vnb73Cx6THBTJ01PuKhmRJCVfnLJapHSgPLwTDAH+
cuyyhEnfoQsHaclviW3JWYHQMjehZQC8oQ28vj6AaioAxi/FD+TiBu3ibBtCwO2v
4qiTE53RiUGsYcMhlVodOxOATXm5oX7xnoojZyoP5vfwiDtzj1KP+P8/z3gzxTYG
DF75GICqEWjpWdEBSVFYq33C+efa00bfguTa56efTikMulN3Uw9FCtzdoos8E6OS
DK1fiN6Ii/KlgJjgY/SZFvxBt923SS6HSe3z6s8iwvBnglMcdCQM8/D8j0LVrATH
BRiEBm3Zh1Xtr0r3TPn/6USPeirQhHtj+DMsiU3XHfIXSvty/VuZMD2JGTqGNbzH
MrA5FV3gmMTvJn1m3OEqfQ==
`protect END_PROTECTED
