`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1aChXq+4cvispjV03zHBo0gOl2B0/mpaiO51v87h+Pl3+i87+El2NPDYR4E5ldCr
AUwmAczi+LR8B4G74YlH5ukns+oc1I0gKWDUQ5PtHA9hgcOipSxRvrl8huxOW6rA
LdEHhyMUetYr+sEFo3/y6PIJ4DvK+6jorVYui9evutEn1bMyY27x9Ysa2Y8SF1S6
fGi5wXHHmltPY0AKE7L15UfeeTnyV01MtzSk3VBqe5h/wm/+LYRdBIAIye1AhQuQ
qZ2rlN3obYfFNF5GYRiJ1a+On0NdsIBhGx7ajnlF5yIQorPnNaV8XN7+p9tcNpe8
ko/jdZX14ygMfDeVNEdDMIK/I0fz0gUhd4tNZ3yqAFl0doKI6JkLqAlvBaKFNbj0
3ffC6pJBznN6ptcEA4F2EChvIDjg1tAnbUg5H7h5uFUXNU1LvfXfnUTCGu4NJaLl
qSChBbIa1DVHjhed8kZiZA/Tbxctn/55duJm8k/ncJ9SVyf8uPtRBP4TiP7PN4Jk
gqdsTuhih0ZDchXan3fRved9LSSwWaBz80lua7NeNZ74nph12Ko6Jgr7iIA44AGg
20kD9Rm0NM+C7G5H/pReIG/bkZJVRojdBf/dTZsZzWRY5iW4bW8EKMIs+r+H0IG5
moxqSI1/OaCE+7V8p8gfMgiFHM7TD2ApyUhgZSsaal+a2IwRjQSd6LqOjwf3FX2t
gBc/M08pTMpJOlQfDjWNCFVQlLKrcoArwXjtfH9VYU4kDOZeWLvPA+7PPOj4sYmU
oXIAIYnkKpXlM9AM/RBNKynEhUCnf4VWY6khg9la+hbDKSVw/1noXlp3drx6OUN0
M0BRgGK2RdSI/LFZ57spUyjKzXeUwV/cVxHk6znqDWvezZ5C4qDD+MgL0H479Lmv
3s6Xy78ptTWwD9/7IM1hiJDkvwBxMttJ8cN+AJ7xINAo5calakNqbyyn+beFFv4q
gOKv/mMLtMMPnH9eGaEpVh2TzmVhWL0+h7fkxPwcVIa+l2x7HbwkcZk/b52YRDV9
0YJpZMLs3TB6qJp7T3p5X/W62NMZzUzi8iYe/u8D8H3yNvCOEugcvINt/rC6iYl8
l2+vEkqFZkQW6n3zpSTjzYcJIANGeHWAzfaZ3nA94HKizK789P9uNAezyBQf1QHC
NtokUUbq1QTwnGMdpc8S1j9Ybh5hUeD3sLcetirJW4FDAQeByZ3RS5Dw/1xy5ClX
`protect END_PROTECTED
