`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uUnT0+J3VNm742xEUCXR2Ib5MRJK2oTSWof5O3qQcW65KLikcb8UIXwKO6aoqpYo
yvVdl9j6o5rUp5B963LxFSyviSI17VP3atl7ALFThDE89az2zWVHxmiM1J1/6mzH
bXwYYcG00Kp1WBkBuakyyUM7V67z8wcGrygsjhrn5how8RNrxqx8+fvUAzcBcjbu
1QhhZqLtRkOs4zWgVDvv5SIj1KvzixPJO9z3XIuThDqA3VK7C7Sv1ABK+Riejjr6
Y8YfVVb+aEvCJAJM1fUQp/UoOjY2X9CkLEHsYSrjwisZb+OcbP6ha2fGaUZW7HUc
jHf22AvlrLe33KoLNqkyjlUCJT1cwk4YhThmyW0KmwDpLuugmdUQINVQGp61Xc91
iHgA8fAVXdQnzdcgx/NA6Y97Sp/eoEgOPidwV0nnNqJ3vTR2UuMWPLSUS27/JNMg
CFeprYiz1HXLT0B0td/2Psqp6NcAr6+YBbY09YNJO04afGJBE6iXmMpcS1ie/YHh
wp3OIfMGF8UTR8vCS0wGWxJJpZWt8UfvYYoGRbooAL1jq1532RBCelvLPIKx01Rx
`protect END_PROTECTED
