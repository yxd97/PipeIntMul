`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YmTVyUC5YG9EH1wJFedO+cgmpaRaulUCr4wRHh18LpKnFyZaQ5dHV2l3FM20Bh4M
fi0eOlHgd7gwtfRt6RTDF5I7qWdud00xMJ85sjiKHN8vKrYtDz68yRg3Ge4ROjcJ
pWGodXSyqTCkiabIgJZcdGKQvnjJRHPThtwe0J1fJPGexorVxWv+Vd/yjNIN443N
WJp7M8Ygx1ekDxPs1GkfpRjGVrBIDSEqYmFqPsCUvrP0dTWBJMe6hjCcymHlSZmd
n+ODbn1iyoBXqiSPUHV9rXvjUlWONB1SK8ywgsCJKY3AROz+abmlnIiEsiXQ0MLY
RW2i7wVPHfIAKMlr7yswaw+BicsZInnuLj/u/mz9KzE=
`protect END_PROTECTED
