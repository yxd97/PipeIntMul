`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aXyJ5y8b/MxGYro4cHAh0uS7wPQ0Nlizlu2Qi9kowG0sjCRJzMpUgMUey9cocUU5
nB7mNgWM0OHeQMfBt8PCrUZv+CUmWDK8PbGfJ8dl/oQQxT4bEv/jX1jfqisKcjdV
28JsyOX0uoFXLFxawe+59nGV0bp0LNRlFmhj1Dy/Pt+SVoelToq+O8FC+zkZk1fe
jR2FB3cTD9+QEh3KhCZ1V9BvKo9WNtd74igWcd8f/270jvKytTF9/4Y+BGJdjs/w
1eX+ODE6+l6FHWNR03O+Rdmo76TKXLxxh7unZq5ubBwJJIIG6ssSQgJRGYVgRKqV
B3YEkqXeMbyzYwt3JyqkDP2v9IqQ3DC6sOzv8zfIbpx9Wxa/DINGjZsdokEVKLsw
uu7KmWyfWIrYBwnp7lFCF6H7O29amtG1BwBCEiq0IJ7sRVohyERSlTwPinVmM6zP
9XxPSi4MRLpVlve0I95fMgDy2v/nK79LyUOdb7HGZtsLcHjfzpGvVgkuBzgNxCVA
kXU56XiyqLQRTwtP0EjedoU+9W7e4SlQm7+uh5uWdwbHPDdx3PfIlTNP7iiZSiLE
9EzbSbzEEe1Kqycg3UYlL9sAfb8WJxeh8xdZhXmZjf52zthq2EMJjml9sU1Zll3Y
wAh8EpMhwfyDOv7pORK1WVlgBT5A2K5d7LiQWA9UE3gYdv9V9Y9494oj/GhSV+K8
denCP7S2kcBTBSON78IUt0I/Y/WUnufoV6ew7GQqeKtIIXlxZxyf3/PdurlvqNMV
+iqxYyfB3FbJohoS1VLeeVN1zgS+Ax5wDe/DDjut0xQfhhdyCkVZSopQxqz5AR2z
pXxgD8ilU2bS5nS5HmNW+7zqmDE4oma8HSI8scsm0JtIG5bBUMj22JD6ct+NJOnL
WChYkAJSCe3Iu/qqrdpHQgLIpTOev41Yuq7oh0i+C/HVRU36dK7lA05G73x16Vbz
`protect END_PROTECTED
