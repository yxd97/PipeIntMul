`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OWvvgRvjajUpWbvFFknZVe1MOW2EzM3/udD4Mhiuy/aFRxef0MayEaFleZoV+V98
ZVQcVljLtxXmsX3gw1AzbobrpLLffAM/+5Fn/cCw5mrZ8T8xc71KTiVVloPWi53n
AOPl+mUAC0pU+v9YHQ79cxHyvczBmJdvc8eT6m2cYDPcGxIgDGyUPi607mQCSB6E
HBYuZHzj6WE6w+OR1uFILMwzPmB4cjwU7e1wI+WQoJM94h4CW318upq41ckB7J3d
ti8RqA9DYoKlFnff4LXQTRHXF/jhgBV4bJeNaUjwdt840OLs5gI3Y9lmJ0vCLUT6
hXWPovxAs7G/Bdt9qETb6A3n8CGGKnHzp1zjLy+s2MoXJg1NIlB/Ohaz8sl6FSPX
4YCT1lMNZn4wsvDfThieynvCEPc+6Po3YPNgeYVXoUalXJuiH3YuHwqBo7NRunkX
3UtrJ0MVgubF+zvmEB5PC0HkIBB1kT/apHU4NiKWP7c=
`protect END_PROTECTED
