`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MnOoORuR09I4a/+l5D5B6GQlKW1/AN9nN2t8Lq3VPhpK7uDea9BS9Ql+lG9Z7zAh
QgK0fSzy9zLOBAOsaVYN3BOFxRfvvZlsa3vNwuOWVKkai4Ai1V+hkcyUO10h/xKH
H6Ggn7sONt742N8I45e/WJBIGVJRc/uJzN0mBJFdCDmpGyaUbncNzNdi9p7hnrjZ
h/XWMmTcL9tNAtPJzFZU62kQuYDqmRq0MrzHoirQ5P7nSQFUbkstqL68xrFxnvHk
KPfQvKFZ5BGmmMgTkp+ab17M1opLr2G4BkkkHCLY+vDIXkyTWdEvx0QQ+E+QKvz2
n2Tom6wCiU1NCNNxX91Obw==
`protect END_PROTECTED
