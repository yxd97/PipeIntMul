`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LZARICpj2vvZcbG3AlIat2C54oGI77nIC3yIb1bFXI+q9ehvprzgU73PHF1qHNGO
8DFaEN83MYDd8TV4He7/Rdb3okN29QwaGGI2DqDPuJjp7vb505faVZWWfaRPTbkA
TIYXklqLA1otDINoCQtSFnemVlGYNlWbGsd8CUwbDpGqIGlhRgGtdW700laLQaYt
5TRElIJG53AlX+c6telpZKPCTi+Z/QYRO9T0KRwMMvPrqYuyp2kGdhZ29g6lL2ap
FvcxS+li/3TOD/M59/fUt/6+4JwNJqAWeW8nXJZv7poufAR5LOfHERrPMt+B35Bc
UYKGkYeZzE/WBLtnIAT3NFEhk+tWuuBymPKNXM4HBUvlsFjf3BkwZrjfC+KkkWII
JZ14oU7n9WsU04Kf6bskfcdsCUe0OYYTzADptsH738lAguHZOcJXD/ePb21dtBcB
Qnxq13qNtNROEYpXbY/ZgMEtDhb3VbsAW7lphI6vPfXcOFY7gWFrO38FGVHiTvse
zmRUBfCp21WdZh/LDdG5zBpr5nmKQ9ivhZcH5eRK9dENQqVUp83K94B4ceq4AxE5
TVK6zemj3qE0lisxwRw+pi5B/wSekjicsK+KfXZ7qv+NzOvzuRx4+x7j+pM09vy/
YewIjHpF01T8J24FA+rpSlDnibARMaIfiq6Q3OxLzPNZ82a4JUO3fluQnagfXnpA
mOwrk1D5K023hcoZzTZTgQUrhUplg9eqH84S8DJED+zMokZEorQXRUwkk/+RwYfP
5fVpO+9gsvzsaiUBalzuKWI0h3yx13nzUOLaidjgX+lANgLDLbQJWJMRgedeg3tH
WqUbGLJuqtDoT/bUmFaUCNQ3GRPVEQfI08+CIcoW4J7qSD8TZMC8YSKqsze4SvEg
O7nPvlsJNJDXYZNsPr308pzL7bJmKMbz+ZP74rrY1m043R1Teewy9Jf+BtQkAjaL
6gTOt2Bd/ohvffJtc+B1R/FVJ8sOInNFaMeetvUGOoqFpE8k5RadxTpxN8uZgC3B
`protect END_PROTECTED
