`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qiaiWP5RIB36Obcz4vU8GJWqwWYJLSMjfPu8+hkSfGLqBhh1dJavvcwN3eeO9MK
Ou2/T/nJQ9a2PaaDgAUIdhkEPlhI32m/5jaw4TS6Ss7uL8LPl6t1QPIEJJ6vkppr
g32xEVwTlPCfYxptYhffXwuuRGrelsEa8Cd2exKRN6LWh1CP6hff1tOIcarGPyc/
cHPotYRsKFZvMx+gQOm9+rJoPvUpKrMV0vvosxD0YmoOQgoJ2Py/iD7LU6qT2aiX
gmFEKOq4qLyG0RXQW6VNhlhfowZYUoRgLGOKw8eS1Kkqgzb6bTJOEolXuE2J0okW
0/+qv6r57JQiIsTcKtVB/SL7XiHqIlkM/Sf4os8O7U6HpquPFFPUFfqY1n0ZS4gW
EbRvPmvaNqGSB/i0+PmQJL5HmeqgOwE2+/lQjA6SDbikEn1CC0/K9p32wiY5J6la
`protect END_PROTECTED
