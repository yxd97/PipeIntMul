`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rifXm2yjUKf50wGvF67bks+70upf4QY1D5DX7S/L8UM8iSEBo5QwVWc4x/KXwgdZ
QAv7PVfE6yUWTv96hXBLToLqRRt2lWsNw95+2fvt9KqkfzcRK3EDdmPjZtznDoNa
3Gpl+1lwE0TydM08FCWzkJqQxPMeeaGzADN16w1MJYuatd7MebdD0SbgjHfZnmEH
PQW4dsVTO0YjfHRck03Gqx2mNtQ94rP30tlGV9qHVAo0iLIfpkpUn+rqPeE7rmUI
1b+PwojJifG77YEPUwKxHNFfj1FzyuFgJ4RGdghaFF3CCFIbcU/ErrdnUbqIQnLI
QTacn1y8j6spP2fRtKLN3qntiCMX+9mrVRyzlHVbetorzzuRlZvN7z6d3Nl9tggn
IKYV9HRcpNmvJfV7phtbxY3tdsoth2H+158YEtad1elJ6m8b2fdEOhDuaZLQDwlX
IC44ck7IipsecI1bFuXH8wCWgwdTS2u33fOo4RV8i8/rbDzDwYoLGZOV2p1Mvv6f
s8We+hJZ32A7VSC2uil+Y1q5n0WUl12gLrAsvy1dakUJWbxABC5OgPF9GixP86+5
v1pw6cajAW/K0cQ/WrHpLLXXcRaq8O8zylBkCPQTnwExbhtj2yoo6SljLXtaFE0T
RvpBLrq41m6g9GxWCV1OkhqHlZt3iShgd628VSlmAclv1pJTQ3lCvVdjs2UM1x9s
37cxTzF3ApXOl7toS2b8YwjW5P+Azqecga4JOwanfG2PNxmWMbtXliOHvPV29NQR
mvaIZlGbtdFDsgachuhXaLLEVFakZw0pLZmsmnN20AlTHRV1iKGf55atUQrGgsRb
CKSXJW5O9EeW4N/ATml+7BnL+/en9Ovc48ztZvhXX4SCjlVgKLAiXWD5qy839k1+
3b/O4nsJIVmIKJR3MGDbCxkHEoFTXq+bhfg3osAVYoOHLYzU8Bn2ojWER3PcNMs/
CrHC3qNdv9AlGVPQ5h/Iak3qND4Fs6Xj3RJmTWUnWtK1bizl9xfeOSQB41p/Ge2t
qHUQ7qo37OUdndO9iZbW+dG4NiutnPeii+28xcSZyyiF9kwsdPBancCrkLMc91SG
yo2V8AOZFtrZ5aclL02Ou/Zjcic4HUYJGs8W09ogVlSph4U+pcD0ihzj2AJimDfL
RE1Qgpoe7qik/lgEhj98U50Q8+iQUT4mz2WiZFakwPxDTpFCR9LhQk/HuGmnegBg
b1bdOawKnCvTZ1R6KUvmT9rH044thUQjH4wgwkiKtBJbEhDVN2Z4q7kN4XprrxkF
jHrEn2uAwXt9+HjZWnh9xu+iHuISsH+GxnM4MiIwpiIBl4qHO9J1Ylyl0qgDQPLL
Uxg4FkHUzschXklqhvErj/leW06uUaXsYgPL7k/9uzql15FWcJXMNMfHW+mtPmnY
2xj4vD+ZdYLTRBZPTw710xZzkocirOnRzCulpt4j6KQeQ3CSjlJA5ELbWeZPzqiR
PpJ2fYeiJcWlT1B72XCEs1VIb67T16GIrGRJ4xJLgYZQVWjRib8tHP+zD1G9yR1Z
gEEjz+Go6BDrmF6hbSEvuUv8htLfg+jHW/rN4/ieOhWvOB+fLxatS1FC24wIzUY3
kRpTSa8Zizg3bMfYYXBny1VmhqSyzC/bSJIcPQQ56GXgCE2luBozVLsE1ZIMuATZ
IA4ZzvqPFrTKZNSWBv3EihVAthuPmlintjEyvnbgzay5oGAN+JdpFlTA8lTq1R5f
kFRR2gqYg/vszvuTSFdTVkYHMSzICx6mbViCLPZ/osO3cckU6Wg44/bOMdSZgALv
47Y0ilirTGVNKxaO6L9fWRbML7CauGbrcRtGgH6HcnGSGVlbxZcYVivLuU6FgNAM
MGDd5RiSPfuNrOkE+RZc+VELiitDmihV+troiz4bfDpWuzGUDGklayQSi4zIMeqS
6h+22KsJThg4iycyhex9yWSDQZczPP6vr5qw4lb/2UPIw3jhvJxbBRzgfDiGxuFl
1FJByUm7BpZsCQ9ppqPlxvzsFTvXccxN2eHTezNLYFYgW5U+rAwwLAQU5gMTrrxc
s3zTyomtg2OY84UZjWKIPD1SiQyqcFK3foDWF0o1Dd1QFsGDevynZnm3L+fQVxA7
8+XM+XkkzJLcrNqixvd8aGkGlp52GAb3aEpd8/hywf1xebV++mWhE/vI9pIpgQTi
CpVB82lAcetXvaERZLWOCbgTvoGPgLHKLE7QCa3HPgDKQHnADtsaPhVBDC8MbDIj
Xn345IHG4VLFVzhQBuNGW98Z+FGTZSaSFGykX+VNzSYVRF2yeiRkbpcoVL/8XgeX
Oedod2mrlohhNANhc4T+ynpLKbcxfATfPiJQJ/HlIz38X5JNN9V4YTG8VN3ZpHZz
VR8X2vzqT6VxNuJc8pqufEm4zh+FK5uxguPFliCY3XzL3zLWwdRtUQyQHM7tm61y
hr682w062+qDdX3dOmASiDZomTWl9ttf1MY5/kYs7tIovtexzfp/TX45cEHdOtOU
W2+Qi6N4yLvMLq35EVw3pUa85mXkC6Hh9uaG+7RAQpnkNvDmGvGvHHPwwfZj2NIp
K3OFhHQ0bA25aFHVaCtgPZC53DuzscMe4oIbZ7GdY4U2b065tujRevUGmg06n157
uNIiA7lwhqRot8OiJDy6CoEdcw/qLKtHHg22ieGdZpKW0hcKJ1/ufJE0181dqiqv
q00sT3NZ2mHG4cmOLbmmqV2oLn0lmqLIu7Hi+WMqqZuEHWtpmf/pSP3wRkeWf5VH
0lxMsKfu7+a8+fVXE1ecta/siiQZK1RPiTasYMylSThxSPMs2sXoHHkdJNjNPZGU
jkK70bm7xU1BL+dXTZpqnVFxs0g5GQ2fRzW5zhbG+pKS43eGgpddCdAtJibf93Dl
RYh5NgodZQufSJ8h2Rons2HnZnIPvXOOo+TZOBSgbVbLAytTmTaD8m/UvFjNNRU2
K8QOkb1sbGsTVSEV9B4Cujfn4IEunRJje0J1iQKzBaNxP9arS9LihOwShG9Cps6D
yxsPpZwqM7SL2MOU91FQQlfbiSZjnC+Ct1i0DfC3vSWlVtQsA3x8nplxH2KCFbVI
C9g+IpwF5zKrYxTtSr66c81grJ1jW15b4oOeGObpF7C1FpIU1dPttpk839rWxU0k
z4xDTzdsHsQsx/pwKv1RFIS30djWUANJAKvvM8TstHF4nlKoXjb2NSqBGkoioC8+
6Ic6X+BdaOojITshpPmUz0wcIUjdkh6P+X1RqB1IEjoucEHnivhBRyPgiGvOYC/D
AZLBaryBKN1FKA0MfalORkTEITCjT4nSBSsDBcQyZ4FDX8SENLrNxvXWUKHDOn/G
jVst4r8SwpP37tNQs5F+GJkMfqe32tVfzl/XuPx3Gncvkbi8nOv0FTsoln2bhWhi
CzzgE6DVm/muqQouCbKR0MRlJXMLhzWVd/EtzY1V/zTe1mW0n64HKOltY+JoSlCb
BhCxk79gKRwhRiIsT232Eesx3b4ZbGMfsHby7LTSCqnBKI64ZBsyKOMnMSpJPKtV
wBcrlpBWeQE074rWOPTroIg+nN1j9OVlyipuPUmJ83sZinqAbDOQfDwpwrOFB1rR
3I6+koUM0N9zLu2YizkdP1ZWnnnVwPAm3xIzN6FATa1oig2AE0bLCTlCks+nUCKY
1QeJT16M2QSwg4my4UdpMUjjJpVD7mzcJf5lBQRos3eubVzutxdE6wFwFlyBTFa8
f0LhIK78HgSqbTNVJtfxXE828X1nwCCaxl9mb2HNXVx8ltqrr8Yv5BQ4GjaiKrUA
Pe1NEQ7WV04YET5NbhKGI4xr7K6K+XkJdRBcfLhTj2iAA9tMfpXIVX4xO2VAr5J1
pkaY1LpKQEM7cZFwenr9PyACz0sRpEa72BmpQYPhS35cAJzal6FttancgVWGftwm
yQ3Ew1+pLU7HOCt7UJJpQTTdPt86zn6R1tlwOo+FR8GLBkppNXAv0ZQ6e6cuS1r3
nNkR//jifDvMlT8SVOOSBTeBJyf2D6S7UO8EjNMhD+detlMfndtV5YqxoQMsUZQ2
NlVBlStXe6iJp4+08DG2+sdgO/kFlvGHN/iBGdBnPU3RnyrJrzXwVb3go5mpasWH
Oms7QnoaFA/231s0qdi0f7NnaGCMgIWHEdRE/XLdH1t0i3MMcfuxkIxy9pi6JMyc
FCLOIplw1MDJkc9zFIuwPH67pIp7c+MIaCFy8vhXyhX/wDFmES9lSip7oOck0YGH
veokE4Mkxqg1CcdueUie6W1T7vHnQTTg+2n9RPgqrGn2Gqy0FTqTYVDpJl35wkUo
CbP/tgZQmFHJdTYab+1NxE6wgMoHwVDFhwXjmeTB86Jqi9Tao/6ZgIVPTsa2x4wD
2cdBwCSWus/y1YkVQDElLRzzpJpj9zzmRoNqT11z6t33cK98iOV3aYvkCLimNj0H
g5m2X84eGJJ1YMWlrykdxIeyAS2D2ON1Q1MN1Er5XsOPWRB3fFdfYK3j3kJkqHPq
KlFZ6wZBUsjXjq1kV1xsVuOLjAPrd+rp3oCGuA2TF2dDjrTO7fmDPzn/fLIzyToF
KtMx4wCsA9KJ4ZpL+ByViZ3FWRjrcHZUlTEFHGx+20qrR/egfkD0PXkCaPWEPjVy
0jsSwd9oipFxVx86V50E0fdOnjVZH/R7hirTmljhirqBBh4quWVkO6QXx2ZKb5bQ
+jejZfm0SLmmcd0D9fB9BlTvSWP1VDuVjnHfiE8Q6tAw/e4qSVI/KH8jmX33hsQb
uXCfpd54mnhocwJIgiaBLu9gHIFm+ZNuDmkYsgqc7VdRZcNtGI7zfc9BjzmzIBfr
wns0BveRXJdgayqeEeAPeSuzjaUV+Lg1Kx9ODzmBkmAWHIhagCKG4m0m5/lf9zOg
Y4eeeY/Grdf0JrGEjcuvZVRPz3JgtCCqLWKi4IP86YLeFiQZKHUxRNpHOChMHkHK
Y26s/YoKdbtBU/58aPBuh7gQYzzQurw15DlMVYQQD7aSM1U1wR8I30Zmaneq7gny
F++HrjTT8M7A89OFO6N+D8a1eclYRpw/HL1FNnH2Z5nXyamBvx/REDCCwgoFCAOx
4kTw+mweL4vPe7VVSqG94kBNIPCdmSxvMgExuu11thSI6u6WrDjy2GbVMNd3ZpZG
TJ7Ef/ytU8qtkcyASVd32MFkcSjKc4hryFNFzah20Yv3OMG3yT0xIaE9gnWTprwE
7IlNdyHjRXBnyeIMG9phBKTqbojNhJZpaDrasfTLwaZSIcxFgwe64ypfEBIiV2qu
lAB1hq85kahm+Gb5EQ+V/v+EaHmJcYgXZLaKXr0qSe9Lbd4szeu8IQv/c2rtI0CU
gERkXky6MMYBKtqIlgUprFZY89C0Bvsj5rvhy4fcf5aPajlRy+1yHiYKtA4xfzXi
lp8Ny62g6lH0lilkJeVxFSi5JSHRYMHU27Cm4y4aqPuvzUhByAOW1zw7NRMHXfI6
K2nev1l4aeQdydp4uNe9E3gc4GkZR/QKCdglK0dqW1l6vaMYnf9JAxOdI32l+ccj
lU7ubpmOu8tq/Lx/5tZ8LU3bJqTWkSMfzzm2Si7lkEo=
`protect END_PROTECTED
