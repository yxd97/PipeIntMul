`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UELUwAfi1MhfiHieOV1OktKawIWBaPsByoJwF0kIdXe5h0dJ7FShwO58JapQVvb0
Ng9fDGo4BRCrQCKJ2fXmAcVZHCeOz2iW4CY/X983dnUJBLSBtCAxYp+NxgfB3kfZ
EaAIJptiz1mNwkqjJmNIbm2xboHM9869aCBoEB+GJsFAJiNQi3GnsHAlW1/qN3G8
1yq82UAsqpCcUsuG3yiWnW1T9sIocfB6Mym+K61elpBU44Z61BBeTed2icPZau+r
a6Moxtui2vOGzY6j1CfHNRthksjQnSxaXwjQ4X/vp4FYwQc+8Egb7RJ3V9lMyxMy
oxwc+3D0rfzYJAh+KDBjFDHpWLOJM4V119f3WObOTX5nXYDp71zSgq9ucWLqn+fI
RQ874b7QMNIG5hbn5H9oieaO2jq/9RlUHli/Sy90RHU=
`protect END_PROTECTED
