`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XVzj1ErnlllT2PNRm1jPfoVm8rc7nR7V4lOzppn9NVnY426FjIVX1DLL/nfScpNY
XAsP873dMC5qCcfy3B1BqTSgW7hFq5CCkzRfgHTCWyCX/PBg2Zi2wjjpmTe0eEnN
SqHTzziS6Fthrxgxxo3zcF2ynWBZM2l/DuLdjE2X7QBI+gIKJ1joOtYCH5bkl04z
5lHZJbR7plkqHMwUz4Wmqp4IOyaTdRIImqO85HULRhUOLtVaNCZNGJDPSeRLrgRU
K30Kz+qcnODEFKuCnsrPeiKBMLUpFGnMaOaxE4S/Yq2qTkX1KLJvu0u/OyZ/kU0x
sWt+4jo10mrSZsZ75zdwP5OkTXKUgdQA1KALeiixaT4ozCYQFskvSv59v7UyMsZU
jKyjrqbbNPJwSGRt0Dbanc3z6Qjrfxdj8/vA1UyrI6AVsjeT0nCAS45mAGTQKK31
E0oMafV4u83n/ohp+/Pu9Q5KO4xshLo+VlcB29qgbLVZzR+uYgNeh7xT6wpaTzg5
b+rxZ4gZ2mfOQ4ZfWvs7PxadMVGt1jEbTY5a/O9K2WVNslB8s7/ILSLQ7daBDJS7
NMV0FK4sRSoyIA99xaTRUbKpHihEPRjgSm6LRpERD3s=
`protect END_PROTECTED
