`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3vQjVTY0AFUR71BqLMOvDX9KzW92nERpyetm6hEZIgOh4KgKgq6tY14q8B3u1x4a
hzZSZe8md2DkkpvZw4Tf5T6P+AdgvjWuvuf5YkbImeCpJPmS5s+md8iJePh7OGgg
uLZZysjjPvO4I/glpdg6OsJWVa58VJNJPGEqrdu5it6TrlPNkeZJuSvmVj/WXMzr
xVQBuHZejaw1iHIQMew41yv1ChvFwBeWxlWqgRpuKmIe6lnfV2djq0rckIQH3SER
fvui+XJuRtBA1baQCfUxwUFc96pqRAxF75aJa8uSjsJy/Hm0IgbSxTA1kfBwzZso
`protect END_PROTECTED
