`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CeJnoHAwbR5JNplyOLA9W0ZfQ/WJmZC7P8Pw321glmT9aRnYH1ZTiMC75fXwi9y6
+SwsS6ENj2pMMe5RC1BiUrfD2rLck4RXqANwDnW4w8vkXOjbndF17siyEEikfS/g
ONQQfnCrbMgEb5HE6ho7rLV0ZbuKu1WdE6yyRvmdoGJQwVvoDyw9WmxwBeVdkJLv
ouNJ0i5pd2PdR3FL9hT5SPjfUDp7Yf74QGIpyoCiGiDOXfZ8lXarrchSrUJrvcrk
MuRqfdcC/f2Z2ajqAg4Ug572HxL+r/+iyFYO8HDWmpLSommglzHEX0k3aao+WlkF
xQeSDtHhWkSSMUiPJ1DbTgwSCmZwzVMSERzo+V9shXCKpOc2ODXHWefMrNIL2ZJH
MA6EP4DJt08FCYpl3hRwhTzYLDuDDi6Sm1Dr+hZi3K8pvZscoRiQ5o3Y4+9IytB4
ZmrJUtGFXqgwpK1TEI44EhyGfpDF2R27M0qc/6aUNcPXJZLv+AREYWIhM6EnI+Pw
uyhj1J8yekvI5NBHCzaCmzsvo2+kP9USv/OaPkr8zwYzDwK0wFta338m76fJpepH
i6Ham9vUQB5BQpoxZOfHOtCpMvktIdNV47Z0rxk3IVjPofRrKrSXzgj1FoU4ZTEs
NetDkTlrZoiVxCEh2xum2UAKkLJLmtpjo9EF/oBwzCADvv6Z+K0zm/qVjCI1gg/w
kJ9f1/CF61lASXw+napTLBCP21M9U40TerFlqG8nYc6rwuk25Akjshy1ZOfwLkV4
JibaXdNC8gat5vd928bO/A3ZMUo4tiqta7f5gpQjDrfIkPUCOO6wMRCqQ9j2+J+a
/QYg6XwXEFYqGTXSPyqy3rhwcGobKz+pErEypG72T9ICnwtzf4zhMUFnUb0vv5qw
KhQ/CCNXgvbCd6xEtkTm+CfNIs/0BvhwWWMBBpSY/V8p9unMgal1qZ6bMmUeImuV
rQSZGPbU3zl0uWwN4nyHzFpR8Vwt/TgtyzoEsImdvh/h2sg9IbRegkJfh0gGM4DY
TwOSqF24/NskLMrRhnmjstPTOOw8TQlGh1AQS8KrozBEvdvdE+ydnYTfATwIxCPj
gfvcse3AVaHxuqRvt2E3y4DNMTUV34z4KvgggZlhyAvGMqK/7visa9pamb2xMwIq
vHV5BNH9L5MmTNeNI5PPWS7jGx7lIJxvH0mjK764eyxP/1Suqrr3I4/QKa/7dIVm
jE955bf4po9qnBuZb5dddl4OMvZFXxLEHZXMWIXipkWSxpY217XljtbUnWdMjpkK
o6l8hes33HPpfRUZ4+nSyRPwGuCesJihEF+pGqykNgDJPx7uriTNj1aaEjp4x+Jy
/WnZJiu8WWHMnhzyK+6mJm/fDscVDY4qqIjI9lxZVqGzjCJX4fjZgfUj5lSTEXM1
wcX+kHt2Cip56DoPVAi9kd+rFIVe+OavKzyHuDaMjAaL/X4/r7Fql1E+WvdY+9fI
1J7u1aPiNeU3QuQZ8afZQdj2LvPSC2rIaSqTgy8ZE1v9pAZx+o/0mtpzjLfYs/r9
hEzqPrRANoPySOXl3yyDJg48y9UcgDJnCmkKSjK6H5UpQjY/r/46iZlETvudNe4V
`protect END_PROTECTED
