`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Uac8s6p5yOVJysFJfmg87ii07m7mfeaIuSjj+OKEuZjcydtsO/7WO5byC8k0WjT
LD3TqQhdUKYZDlQCUP2U3VC8EcfsTE7wK9k015hfnla1tomNAvQkvwz6JyywhXS3
cApFdUSmu7lZ4iSzUJV4dC/jXRFbpjKpPLjzzT77DftyiFp+qbw0J1aCz6gOiLsa
U3lajw1JWkLTWxM74xpThQwu/jEP4OfMGTFOoVyScWjJ3fXuJvqb9XMG2MNFmAn1
hRC4xkho+Eta+N+Nnin/qhzY+GaJy2Nt/r2cpPJ4nri/dAMdZ5GpOoJoMhhb+VPA
NjlYy9BeTNLacZ27i9o2l2NGwxopT0KJgWDIJqSOz+7DxVrQB5b6WjTAsKsn1K6G
9R9Iwycp3g5DidnDgzBRR6esFy9ugHAHhGhgXfVpIYvk8U/S3vkw6X5TIkKydhU8
+4MqCSXezmqBzlI9AD+fM4+ZC4kWawoU47mY92cOqv2nxqYW5M5g0mwc9YYftgyA
uVwyjCv7TpEh6CZyYw3jm8ESAUwDBxp8N1TTI9XtPLEaE5QDvBdw+lceHDZYMqGw
2/zyfCads7Oz+rK73cJtjP+fwiMqJ+FEmRdyc3k2IoL7Ya6YQBSy02/OD78YgcYE
N3zyRQpwl4jJ98QEr069LEecVbEYCPzCEaJ8vHYn8sUhedW4jp0sbUAxkn+PtIV4
FkcnECt16e3cTq4Z8SxST6IKLR+1Mj3MnrEnZ3bL5MZtIFaelxjxBBICEt9Q6yHr
caBnvSuqkacy7n5YMwJK8+rq5V022/Btfs7wKRfbKIqX8cfXKWI1pDjQruGrhI8S
Ygphm4oh5wJgiA7+stLK3J1nu2Vu0E9IzBB6a8KldglBuG4ylN64Ivx2mxYdfbKi
tO9//dXiWi7+th/TYk27x0c8j/caBMpurhgDfOic1NoCdszwUlVvpoORcXpD+WqZ
e85Bi/4RaCkrn+KAfJhHzIENWIRLpYVFpIOELZBqoZ9qpaGIiCxfBE29BKaY9wyG
lr3/FMIL9PQr1H1WRJ9IV1y/HEg4b0LgHHbxe073CZiOZ3o4zKJuC6nzcLb5NTUj
GFom4tMOFyHK30ht2GLx/tc6XXWynXmyFaxOjNz2Z6T5h4ycHvRt4vPW5rWjAJcH
xgH/JIAIEqseN3izmZQwAmRS1Gm2G/vR74wuAEa3lITawdFpmL0IhzSrxfkgi6N5
zCJg/GoZIuM6inCbURj1zY9EPqw39NBjQ1HXEow3XJbpLSNmS2zjReVAV2umxR13
gKxsyBquIAjgXEwIxB6ynwbstqVftrZ2WnnhK5pi33AOeH2n936Mfi6Gwb9sK4En
ISPwFL+MfR49nrofE3xigilBN7lTTqp0tH+/qBr0q3f51ITTBVXx65Orzha2LIKi
AyON0qZLovGKXWXKY/h5dfFkP9an2rqMGZZVrhH3BLjgkxfT/r0xpiGTXvBygrpY
gKCoBzgNWtM0X4hpHJwDX0wNBTbFVmxOse/IlbuCCsakuqet4Bzt3uDgfvhO07XO
HtwCtAIixL9+xNZDXrJOC9uxgVztZfIuNRapNRilG3D+oFPE8931rrz7YN3wIJKs
S41NRI4x0MhNKQGBcnSarqqeM3E5fJ1Cx9gSxN1zB2zi2RRCrDxCbKyk/TFkfVhB
YfsAa7+4wgfxd82nVNCJ2fyMPyKgMFLfnLFZcg8bvZg7GtpKb9b8yKYHQ9+XpCHo
3rrTigYk9jnCEfnVLiGex+S572fhKVjDpr6JPj3fGbq0APoJlF/yyIy7ZUAJvNh8
RcsnoP+8wYbLKA+FKkmeNdfqAPBlxAVoIwQgdVbpID2mdC/H4t7qmlkpvsS5VHrB
bsOcEhwXcAI5TDvMjVh3MfVaLwffUCd/ynlC7ROkgrgOg2VtTyJqc2GLVoOhia7K
rvWjI5x6/kPv8Tb2MoxFxqVxaFiB2R0Pv4JFF5WXxG9l6bQRhhYkmuumjT6OE4Ln
S+542pW/gQDzwd0y5r1kIAKru45XnHjlGBaqCUuid28T8QbU+Qho5P12qnpVoDQZ
ltGOubVBs6RggbBNMYLXn1Ex/m8+F9QS9K8yKjs846YVHEk0oa3SQjFpABGqfkNE
z8JMeI80IPLfHZ49mT+Inhq/fOvLdvfoL/1IuKtEwcYnZC7AfAXhJCKwhSYAR4AI
Yo3nK3OsDS9sZDznF+Xsq2Ye5A7n67MrVKzz7vORI2ri2BlteKNdHufZM9+RSgXW
uhoHf/QdKU384+FwoeXPkwbDcOrBUq0qZ/+L5taXtxp8/ipWJJdvzoJMQXTtKAki
QgqFLYUomWWNC94jMF4OX11vrGXn9XfP2/P5gzO+4oic+rXy2JBZlqE//spgcM4A
nRP1Bsu45xgOgnejBNJma+6gF1jq3y+lvCfnENFnNtV8l9ksXrdEAqiAt2iOHcs+
zcHczAVYs9unYDYUEPUWIfDpnNO4HbLIZGxIj+HZbcIRbHVUCuyw8OVXT7FoOAHS
sj73PJ7YJIApDgXzGH4SEjgqx6ulqNmaJF6QPmKdNLu+S6LhMjQmDrkeTD91f+KC
J2Ol3JPcwQXmUxLA5q6y5aN9yTqcNR7spCtc4FdsMiJCUn1TlLcFltr3j+GkvzKo
B54+SDvIFvmBTxAfq1igedcYxSzOU2IYX1MkjrjXMFpr9T5AK/fSJfGQfFIXxIJf
hHhS0rBgiAuBzDigfQ329eKki6V6SwpucUI9CRwzMO0wndj5WPA6EVAyRufuisGN
9AFwLvBEolyNqR7VPsZT75SDjj2GliMME4oLKt7R98SZTeu32fUTidID0gw5qYJ2
dqBmBCkDL9ztqeg8gH7ma8GiUlqsMmc+n/yermBbjC7kkzYUY5ykfalVFtYcbtUt
HHlrZ5dEn2iUDRq7zMQ/sHSlsHXEDxWg3yWKKpR2K/yqlRS4KfgN+Lxu4e+sd/Yv
TdtC8KdzP6lZytb5GhhPnxj4uEgrJBobWi/1OwCl6fzR92KvHY6dYs91HgVzaJOO
E7MBJ9qtYSeDTIz7EPpUud+oPXbcntVpYJ/Z0L2Md2AE+N0lU/5EwJqZ7nPYohqo
eKpphSKNaYILb9WgBePp3gxMeJuR8W8nxHl2+cLBdblRVCNS8iEZzVJwNDjJ/jEn
KCztSBNJNz2vg354NzP7NDulpUtQfkPy0v8B4CVLi+O4waaHlRXsOl4hSGhE8/z/
d2WWVvJ+pqehtPNe0+emfj0zGVZyoboCOjGygX17bG6dDFU1e9xBXlIAjxkxtVen
jE95jtvYIBSvONLKEt6y7PonIKd/8A7VBfUT4SvXrsO8AP95vVhgYCnab01Iwsr3
QCL8rl79YmkZkPs0Z0t0G1XsK++nODHY5vFmSEGyvPCbFeFMJsTFKXLle7QNUB1L
AE330f1x8Y5MQYz33XcCymWXRVF3pN/faWAR+YALbawnXtwJFWHMOcbPjyU8LRJx
Ux1CWP1wJthU78I0TNZJ4ih8NZfKsCkYnkugOOe6hL8PSLDylvJaCkIjmIWcgTmo
YTFrQ96k+Gd3iTfuBoitfNszknK0Kc6xqSEWMK076fPEBKUDFZmlKCaesvievt1l
xeF+JEwGTGyIjx3r9zSkMfqVCqz6mdbzuPiuBrQB3ebYwv+3RFOXCl4vz/+Wjp+Y
LYsGHbBhbaSMoeyUZVLuyb0ZCOyyypYYoUs4EdiopoRmZitSV217o/O5isvWD3un
81VNFOcZXM5p7rjX1RYHqa7tX5XLm1J+B3wPwhd8x9x1n6WVQU9rdb4JmmNAcC7D
rMySCASZkcBT7ahAVad1TkxREYsx70dwB59GnPctXa4NAqA2GBBkhdZF8Ea1x7/t
liQCaYhl+c8qC/wMEioldiri0JRuCjqjcuhfAFku1hlc8phewrTy4S62oSL97m9L
bWx+UpRBKmskc8aTdYmf6LlroUhSoSy+2gP8cMrlTReCF7rm30yDM5EL/Q9uEe7j
FystsKibPcdS7x12ZIRIB6vB8P+ulY+0+wwZpp2/weLdf5DbHWT5RGgG/2ncyMNl
gE0NcbzaSCGmdnyHD3CI8Z6u69zTHo2ShEiNiCxOOa+1ZPDqEMWCp2ov39PC7afG
vtfvwgaYs71nYW1VxHDPLmEnjI9VL0VeGVnGYN/QHEmGtJxMIeRbqcXusJ/9MkIs
gOBEKlMV+vhZc1T8ZDaho8Y5iwyzcI+BNLW2jFiUOkIymIta70W0jqWlBI+ZCvxT
PulLaa57uzMpczRiwMkWUErRTu49Jf0oHwsy4h9qZH1lcPQvvOVisoJ7WzZk8OMZ
Uu712+ZTUSaphNJtdB26qMxDc9uNmh3edf67FFFgd+0/2LvmQy1ufExniRX3DP4N
4K9cmBOknZx6V6fPe8eJw9yCgXj5XvybO8nMxVLKwz6SrGvS3ZXvH9f8nXAHFit9
UTGMIPAmhPnpvGCk43J67ANXmLef7EmR6fq4Mzkiycr3n8bhBYQJZFiheD65EdnW
Y+mma9wV9LY8WEZqpZCy3dHcRU+eDql0sismo1wSpw4XKkiemjkV8imeHCXzbLx3
Zo6jeR9tXhj4z1MEDcrr1sAMu8hbET1M8P9cZV+T2LumD7Rxi12woaY4htm4nZVM
lwVRIGHTtrdg6TnfrQQgVK/Zc/P9N9ELhRnYFprAmRoxNhgPPwlmkE2h/lMOwcn+
L1w64KbXr+6SijRo9DoktW7wqAixEq6NHpShmflSAwToQruhLFD8tSQc4lBntuYy
+2a7o45FvvJq3Kq4mwi7q2fY9AolP5a1uiw0VxBJhi1R1cgd4noDGpnY3GFAkmvF
USi0sYrtzupKlwH6ipcW2W1LWUPsfp7JLyeBtdjWLYehzRjfgDTErXPwr/+9w9sG
yl0eCajCqZ8MtErPVP4lyR/xCV17KsLXaS+7OYWGwBYOGpViL2gbaRp3ozy89C4Y
qahdxJrTBDGT5OWMFMaWSYB2bEqKdBdbczPVe9x1LbD1hisd7n5cCfiXCbA1d9Bj
sztBcsv/k7g67IGBcXjCMsLfD2ImxuIQcpFb1kzC1ct2YxocfJ0oikzIxZXqxpH+
LVThiq7HdLcOazUYEs83TvQlTgUX1GN3zZSLZudoQeJ3wGO/xhN618C2jTJJXMEY
RFAJ2GmqV8NteGXjlz3MWyVRNy4oxBMJzs8ABoNJMj5q4ntxrKh2aGlpnpVB+e3U
ld6xCZzK4pxfR8rrjkDOKY1GsLGbSagPmv1ofWY26w2dBL4UwTBMgVIRU1TecrFl
/kvFlGfHuH1QTT9bDf6fcLyLWsaF+XuDzuEHPJZvHW1FGDdU4L3pz3ypga7Rs2xl
0zpYq7s3+0cNcN0yqUWdw1ymHnIe+LNf6SHr+yGp0ROcmfV5Oh2DOum/vNQ0IXHH
zs9rzRgmZPhGJZ+7UKuSw7EZw4EPgc+RZ67iylnDtDbZq6PfJU2fvmjokCwFbj2H
LlMB9+mDYrphivxYVivKqONxFKQTQSf8SXZ9uPpp2Evf2fWkrRPnACHrgbKjAJBr
LbK9kZA70WR8VlSd66dCttaQHnSlgKDlotjFJjHWjIRS+Ms3ZdEanQXdNf5CS3X6
I3RGrvoK27MvD780w94hmJHnEn/NISi7tj/zzmuQssDJesQ748gadOfgzYZ3u4EY
8JzuF9sg6IR+KxUjlXx5qH6kmMvvMdVpjQf1eQQsFtkWKoFZqWbKWSuXvejvhhGE
LpbqlbGUC4A+2nK9k615F/9p7nTJpA4qJH6HGDJMNDT1soauiagz74tG5GLiiKnC
g2t7op9xM4vL3IFFrWxmK5Zi1y7rO2OZQtjm8Pz3e3ZrmrR5WfNUnu2yhinqr/tY
aAyN8PJHTiDbz2yZTp9KeUWLXAF9Qz9Ld5voy4+wWcqX/FigukwpPbj41/yzlksO
q7OLB7SER+Oc3mz0NfkR37/CyHkj1DpCtJi/sXFkzDGmsJydnBF7mVR5AKzXpDDy
CNGI6RAswwenLV+TOERomoS+Ezvz7DegRvf1IqtgQB5LzdmzD8nsfun6gDzyyeF2
KEeABSveDO04a89CEMzs6p8gKiaHOrb4Dh+/7AAG7N9mZB+0/Sl/O7jIJJU6Wu0d
lKG0/2iha7VRINDArF9GHtYEti7M8xLsLWbUK5vh78ojBQdXbbofDvuMb1wbxnQp
YMe16dqsEhyQGwc7+O+PVq6Ict3qXLIkhQu67hE/cxm1QP2WaHMKDnU+gTIeuRkH
YINH+Fu0Inqw8A8lz76ZIafpGiKhDAB1UEYqWw7f3DiETYDupUMSWSmfx3i2Vw8V
bnPLKShFeZpPdhyAoqyaQgtR4ri7j7o5oXw0AHw6yLs+6Sk/q3/kL8Ucbzl1uVfc
Uke4CxIGHxSuCt/cLxSWxsZBc7erVVgmgKKQc3xYKWh1NmLSLG1L9jP2vCEUJFEw
OjJ74fvFi599x1sU4ilkJEkpnTshF9op5WoZYE6laV1fkEBckpGUfaYmnWabuLWo
dIakWWEGimlikpWPhi0106JyKo47abCRs7hflRKOZI7PnGou7VifkVaJMW1rtgeQ
LFqVZsf+GDBDOuZZI13nH4EgJeeHE0M3odO50nTQwUdJVbhjmSAASECrTm/SUfoh
ehcmhKp4hKf1n8p46ckZAawjLfGgO0R9cG1qgFo+CXCfwADipIyqmld0otp3qsBP
70TfoFYQ7YL/by+TKqpq6BMf7mbNk72AiMdD+wGLDncO/MS6i+0Rurq4HbjPpdwx
pcPRFKUERqcZ4iSwCVNvPnfhe0ZoJHl6JVfDm7TUjcEv8Q8BfsKGZJVaexhjsMly
XfhaPfBKW2w/Whj2Zu1QcYD1RxtzvesxfSfNwLSeDXdUKJF3DLd9oZoU0OQAqVZA
rbUFmgZ4nqCijxldT9a/FYv5tH8NY3Oc1QJcHbT+dd55SJnkDeTMDyZhM/W9IzSW
NMX51J0y19iAHhVNtZl3GWXOL5yCfPwIIV9IIn37RbEIjjJj2rlTdd4R7ktpgflH
gDTj9BKGQ2UsJ1tiNUKhbkNIJITjxf9bN3HLs7UuBH6hRhJdeUneHBP7xlh5zzfY
yT1cXiJ/96DnFyya0vu8VJ6sxBdzaU80X58QQtKbCkKFlYILKeVymNjqxygBVEkE
myCYyi4Oke8nOnY/og7rtdAAUrhuUR6m7RkFJYjzETJxYzfcqtIQELCvzKrgRw6l
UwfRz0pFvGTZRxsKqp/tw6Sxyvrzb5Uc7SW/wDbUGY2VXc0KcN02Mg50NL0GXlSN
nlvMbNicCtxsU7AjL++Mvosf+hEbeSMWGqOE563WKtfwkO+Nti+Qi0saIlhZxY6P
COjWsOkhqI57dg9RF3H8OPHnhz/oATlzQMmOCZRsX24opvYNfspK+1sCikOb5znJ
0VRoks11bp6ASgPZTuetzNoOFNy22l31oI5xTtTJsS0R3UtZUPPPcpMOTKFX6wB6
qETquqeKzDlP6lSzFZTsMrdv845EX3v0n68Sf42hNjJKpIrW6OAR05Dz1FpZUp3F
xww30r1P2oI1uKTnkzxMDJELxze2BUaqRHN3vIgKRaGBZ9HL0ZDL6RItXrgcmo5I
p/wWzmM2ErUsNKBEST2Q4dG8BPZhNaiO66X/kdEoIBOW+e7xUavY6rAShEbPzAQy
A5X1CeTSGkwVaaLQTPt4fu3Ob1b5jLLI9yS25f+ibvTd21zdKLHZG5FoMvxesY2O
xrgOqi0ij/g39yS2sikun2M9tEQTf/k2cXDtRZuBXo2XS6FMMbwIg0P3z3ae8rxV
fKnv7ljvkUewYcr2lMLoW2jQxn6VXN4pvyrAPNc/eEDqSYnyxMvAwHb4bQ2pcRWn
eZkNNMetwES+SNaEfsx+1hMDKXXb0/AP7V44zqDKZe2GYNfnvPhnU9A0eLVarv0n
Q3pUDv6WhMyIsnfzV8Atxb1X1Z/fIeLPDnd5hdBm3s87upMLyUUmHXyrc6n0Kw6h
VTWdiDH2L13IQm/w6DtgXcmd0q2exwHUy0qfSmnTTvSi7wbmHYlbAn7MYRYz5JCB
/JL8hids2FL5Fdf/XUWfvjrcLKRocNLroxOfeI9b6iMNjE0pGVXctDF1HwIogtpN
vX30zwoGNtJkCcVC7K37NOhjJrAvhOlRlEIIkhW25fCFGyOUUeXJd/u4TZF1zL9f
At0+Tt2/ZquswQhvaucBDEWCeVs2JqMlD74Ba5b1R5QHAcAOsXr7PHi91iBUkn0F
qhDuiE/eeJ6/j2h3ILAS9tzPDgJBLXy8YuUYkhG3/9uQ0/g+rDrznWP7wAd5mRNZ
tmonPxkb5OeOcj+7hbCwc+tX1y+4fEIAdfyEAGTF1WqycmIyXSI5RuotOHKIW0Xb
gUKqYmm1/f52wBmIDnVtVrFWz2P86idGJg25lE6th3dhu6DkgJV4HWCp6lPVt6Gb
U3KqTHYezXauA62cXPjc1r8ay3v2hb2LnOZs1/w7GszOap1cQ5CRsRlxog1s9vWK
ZVMqC+KfmfyOBw0GtKQ+DCTlC4O9N/6ZVArjO6zwRN3fJ3FHk+0ZaSsufygRS33p
vNyN8EJD2JRI65BwJTJlz6Lxs5jTPRJXX57QCXHMgKWOHBYS3eI3CoEkKMsmOuO8
NxwU8VJ0B6NkhaHsmBYbPigP8dAotlA5tQ+Pj1pE8z98C42WEFdEJNEvq2OJ+sfk
Ug3MBEyzEeaLMa3DgcdSuugCyOBCTqu4vxaXAy7GJv6OfBZXdWwXmtAHixXjj7QD
XS1OfSx+dRXGZmiY3it1YGrJ0IytH7CxPFJ8uggdWwfcLrJEs+EJhJzdRUSe5zff
AsfEqD9kN34TbN792aCsp43NNHRJMtB89+HV7vsZ4raFLNfdtRfPluTWR3EIW1KW
DXuWzQ/Xi7UPa4yhWTMeEjzY78sjQ2dKHu6n5c48gcBJC8NS5WxvdU53BP583KTi
Q56SqYenjZRCtNLQwMF5r7OZ9Y6QDrxIXqQdz0sSiOJo8RHPqP0OZiGRRhz3xcGG
Px3OalI2wLEpu/+MHvwk9STEfj1C14vebpxR0PhKJ+hv48sUDIKGNzo6YI3rP/OQ
Y747o4vscJIklAk27zaFozKET3UckEE6tVG4cKLznZMpre3Gy6VhD+sx0X3kLS0e
SOz9gtUME0OQNtAqoKvoCDsGSIBDfxQPoFWsfvx0wyCng1GWB64ysyZegyfFrzvs
TbPduFNURQWYRcJy+/2DU5+FPuveshfMMZan1Kbsv760OiOZhj28BhUzviG2xXMI
yQl7jkpsgINYVCkYdtk+oyd5nj8TRU0erhvQAvkk6PWaAc9fXdfUKcth1aY26h8q
eAhH2W0hrLj8h9rkM53Avlx+VcHgvnbmHYdWQ4DTD39QHjOO1bgw9LoKxw6nAO0a
S63jhYeQPgm4zF19Oh28ZjeoYf67Ss34S1T72So9yvrUChPY9/1DkvUzqgMiuvXe
C/wHzKnjAqUtKhnITkz5yyjkK/RMz6if0zbW6GmcrpPrd1mt8zpuBeseJTfO7x7Y
Vh8+6pl0JuttHPBBFs/gDaX4IaR80w7parTHkskrRF1kkhOJfqAkiDFwfQMBHcTp
/Yg05Fmh8zF9MH5j+HnSRbBQjvMJyKij02iJE2w11IHIJr8N/NmkL6wtXoFZ7IWp
u482MR9yJXVBPitKJPZcpS7ocjt+HcMOCQv8F3AUXX9TGqS9IRdvcOKr02NXHr/3
zS75WU5frLXE6mAxDNelnwXty7iShKMA6z8dXfQs8b34k0SNR/7ziSieGyEQk3Hn
WDv/rHwUsunRg2afKgdn4zXsTDIK8jkLJDTs5dmPfHCkyYx5xECtL61JIJurX1rZ
AtkLOaq+L8BXnud5smxm4Q==
`protect END_PROTECTED
