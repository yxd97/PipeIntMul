`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K+qHylc6Fv/09XkIiI5JFFPcPjMQPH33laAWgUeHJJam3aADYQyAHsi+xp/K7bPg
M6yHaFoD8mP3KGFVBM2vvOeQ6QhBNdTIOFJGaH7cZIj/ZVHpxNObF6tY4LZKW8no
6hVuen3koP2xLUwkfmHbRCbatmQVnEqvU2JJJPsAIn9tju6I1XmtvldRxbxNz7jv
7pEU0E40KZrz8L4yTfMvNmCAlsS6ANVbSdsCFeQsaR23F0RHxVZkb3m+LH070ltl
YDCR3qQt5t4IGqitQsjwjEsfKDdktTqJcsPk7caZfG519/q9+q/S8vw21K/y2bgi
044J95HGNNirbEnlQNd6RJHKZ4bAi2xYiL4PVvJyuGqQtbOJct5RMAOGo+DYb0j6
dQrHQgoCDJI4AY546PQIUKIDLGjIp5fMfZBn2JB09Aol78temkAZ+b6GQyAhfyys
s8XoWIPVhI3kZx6nRV5MczYbiK2dz8zA4/TV1Y2RDrg=
`protect END_PROTECTED
