`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7D8w1MDgd6qWVL6lA7D5WnGJ64VAAaPUqWw7TeH/WMluR22aNKK9qUm7LDusEjNO
gXE8KbGhxTS+nj892y14oKTCGf4/DPMlyDdqgEVz/RbN8RroXRsF4hU2GMFWkMob
bQfQrgmPi0j5AUfxGfEdGvUX7KcfvICXxZUQw23VkV1+WySRjHEsd+sWSfI5MPjD
CdMwzO14tJ/ZkYIyimCfwhC6YbIVCE7mUE6igNvZeMgBywjh5ESHDg6sQ/GusvzU
OoH83opM/10kQzRKo8xcdVQpbAINeioSLeOXApagQoQO1FjTc1WvZwFAlIjKxYPQ
4NZ8VY1Di5ACvbMfjz/lTQjLWabDqEefSa7wkyoQlJpWbLnPF4UKrLpmbDOzER4m
Nghd9dYJKKSQOmW9EY9AqayTBmc3n2D81JoBH8f9x0R8LYoBrYVddM9+yn/WjMHl
r4Pn6P9kkvWAZ8Yd9XLpm/d5mNmHM+RKl4NluBLQIRyzooTigoEjR6WpfLzzcp/8
`protect END_PROTECTED
