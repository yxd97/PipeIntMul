`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DMyQnBpq9O7B3U9P4WN9yUizTvOeWGCP39Q0+5Kp6DVWyPmqoddUKLusNx+DA3yw
ug93rIqLb1LvNwm/z17uJaeYg1xGKbyAqxKeJrd2LOpTq4H99KHV5lRQ+UeNl9WI
X5BKev/c2ATDXIg0VuWPVWI13RyvG3cPlwumPQBZ8SDelbOo5E7IL7XFuBzaRuiZ
5pySKQqbOqkwE82kEIhIgUuXlLTfSnArJTcC2D/gJjPBW0J/Ke1XGsx1fdoAg9jB
71Yy06NaMMTZ+ffzt2IcDHEjYUZv8cCo64RRBWWSgUmM/X0e4DHngQHdlFOvd0dt
pL7UYAvc8kttcxTcueWw/g==
`protect END_PROTECTED
