`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MeAtW2xlmNbfKQKfq7CfMAGZrzpovW+wL0i5IUD1D81nRlVj0TK6iQw7vyqzc4cs
m95iCUw4wO6aI3csVM1c4QQ36rxAC3+n1GfZZY9Wcui62KisSl1QB+UG5Jc2o+nR
QI0iZ69po06IUSjxdFZwhis/FGglnT1AiibW97+Rfz2RRmQPBdcxCOkXlLi9DAQy
d06iAKRkhg0aDPGMM6RF3LyqiSoBYDgem8+omudj/ryple2JA07FhjJVshfrf360
JX8BPiE0j8OfTMHi8MGwnsfT3+YXjLeBXVTp+nmtSa+jYfTJQE5jiKV392TUWhRN
ol1OaLWkArcijNlherswwi07phqnTxlD/B0x1ErJl1Zmwl9ZA0XcPCMc8L49dden
kGgAj6p0fEUsFf5bYYqD2Q==
`protect END_PROTECTED
