`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EcSSgEOBYPzLzSx8T6K/+IXstN9CcegHv2TNB8pb0tYBH56SRuAvsJvt8UExAMsi
RFiTZqqQ8WT5/bW1GFFGOH2kWTGAcrAX1T0tJ6ID9NK9cquzyb10cg9D5WklQRqH
bNepzMtzSGfIWocFZzAYYvlCoEyvGXM2E3/dEOpSf8TtUHm3SKAI4C1YNe6RC3Yg
GND1P9zKE7o6cJ4Gnymv3SFqWRMhLMIGCJqjSO+N6MPk9WpzVAU9T3dmNODc6vMz
/FEpng7mdVDgN2PKi9uafrm2H0+6/oHAKJYtzTSekCxGWAD3sVFkjrSBebfjboV6
2zfDdKvr9goIv0sPFDhExP2H7kcUIrigqrVhw0PhGOTiyE23eXoEiYbDp5x1yXoM
LeoJFG9WaqwVkRthNnUrbUIOx6eON14jxuZ6KY3LwIO19kpbYS39g0Tugu9yu0LZ
ZIe1QsenVgmC8Avp++0BzZF54CWkfqPOv8EvsTsHqe4Hmycw8u0FOX1w0wwM2Uwb
mdqaNtKQ3mfTQiXndljDg7h+CufboY6T6Tmy4BF7jLRTm004PPAVIXHQaZzYHkt/
eufCbRypo43ur9OGCkLBp+ZsvoPYWAdWvCZWtvEhXAy9VGd1IpyU6hYF2W+WZQfK
DM00xanOo4tUQYS93CJRatAooIYq+ZHtrAnxdR18K1Xin5QI9Mr3d+NjDnj98nZv
83Pc3tAg4nKVOKpJmcOp+kzwzYlsYJ0V8iQfVLVyOSiZCvujd4DwxpHVk4C1i5zq
Ytzk5Wu59OkkrpMSFJYliSccpJuMpkI4N5F/aagE8dZtTRs6SIVi6Cb8dClPwtxK
IbpMZVAcddNjRxH4aGYp1ZypWVKpYDfKpEC99HwOgqQH6lwh4ex6aNX3zdsOea+W
9siVCt5pKqXlNWrSDMWnwg==
`protect END_PROTECTED
