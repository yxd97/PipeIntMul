`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IG6WpItDyPoEGyBKAlPOZ4aFTBTUMQgCUZrQWIlwz4CWeMoC5k7okIl2mlWERi2K
m0eX4FJ5V1vKoYt0QF3u3bGshhzC1/AwEcsRXbjF5T8b/pXIaz/bvX/gB6eSO0YQ
Y6IWFPg9avQwRkwjnoIf+cb03HsAw5PPtNWveFlC5BwSHq25GxNG+YKBBAuTz1UT
kIljhUryY+mW4XPY+OzowezuXD4T+dnzq3aJMYg2VwgZQVYuHGFMbOK9JXGDdQA1
BBylHXxfa047dPa7k9z/D02vQ2JpLKog6mtOkwHBkdzCR/y1Oq73GdJUR4rfnVPR
RNVg5BaKdOrDqzFJDerWnasZzY0t8x4eAwt2eg0ZJPNA+1Gnr4i3E3SAXBtrlNGn
qTg9YAVLgFbvClXlacxqzDIGkGPY94M/87M0YE3scndFTwB5l4qoLCl8MdRPI3QC
A+KqHOx6pzhrA3IzTiWBPJljZMpbvGqX2YkMsj5e2dLrtO4Iayy7Ld6aA6CYcstx
j5iIMhyHK5qfiZyKAnYVYRmcZZFyzIiDTEwKHt/IwPRKTZadE+eJwGJIHkqE3kC4
JyrhDl+/JyQG0qw39M6QEnP1d+DLkD8/ZRiELs+aM4fEsyDYwzjOoPHtRGIsQy++
T5TEWv6eoKY1lY0kjeB4z3tcdZ+4tQ+kC4Cw3plHz4UpB/Pr2caykDgMgdIJ0BXt
NjWsluL03Lqxb0hckLJ3+AH8J7GBb/S8PDDyT2qz3rjK5VsvGQOBi1SzBnP+aizZ
Ihbui/krnPB936mbfdE+M7KEAeThf++1a54tsaKhMp0a84GcxpoleNdbh47MLed4
SnLkxNYj6QZBWQWwfjsOOAtwzWZeFWTUTuyUyOpf0pZa/JjVgIpngb4kJjJeKPJR
l6wIGhkJjxj1NTlmxiyx6WtwW6wek0oRiuJQTD963vVVf79+BUrMpA7zDE1BgCgA
1zx0E+gwzOhKOxwlVpQJ83KWmlmZK9Xs7QVHY4EzsUtpB6EGkwLo1+Q47J+GVQUY
HFYCTKFIiwJo2jJ0fmhwqfERhc8Xbrx/lf+w9QSLqUdZE4tKWsaW0XMw9Y3vKHrI
ZLai8EWwFj4en4/qDQoEGdjy4xvh7mm9B+PQdWx1iKKQOFdNArlruTnIZxZR6BU0
zCXLoqCwZHWKxorccCd3eYjZk7zhDrbv+Zrgzbmnih9Fcnj3eM374lAAiXhLg2TN
ekF5zzFMQ9xuU9YIIpbleKe3yNJ6kKWoD3ipUwkKRpSHPuC2CN7AOtO0Wnu37Zdd
pJewO+1rXeWXj/FC44rcUcQaxNjfsp+nCevAQhrzeYdO5FNLkl1iGJh8MZ74YBln
tOg4eHViMsnEMBGw3aT6I8mJA3bYT9ZZkv9xIRmdJJaZiiMfjmWad3BlcYPN4sTL
mmh4yabRGwubXbYfGll/9HVyloqPxjoVClp/8YtRxN7T5gJHm6reseR1oGN9U+jQ
iFIwFWWxUONqgL6T0+C/yKFxydp0lhlwodEaXwqA0WXTbcKfOxguNbocwJn864S5
OT0CKI/gbJF7x8aAuyRVe4WZerYagJtI5VVBDqXb4kfAEYtCU2mLrbEzDvI5SbNr
nY6zIhF/WKptD/pwjgmn6kp7cYakCRpws94GYCcmVpU85itVjloSOlzR7XmYQ8PY
kLcnCcuiWK+a1WKzlZ5eoc8ASJvAzfhnSYtXMFcxRe37xGWzfip9KGoqYqI8T3l+
fDnrrQrSlVkfzETKLwUJEHjJ19ukd3aUXl7RdMgQORcI3HthxMRXaOKRvWZHnNx2
w08Bt+k1tHH73Ma5DF6qtTZ59XNLXazE8BCMhZ2fl+6BlDVw6Z6MPTRauMdhe2gy
uwYKu10+/Fm8IppkKevV4oB2sKNqZHDm8aYTHbDfkkI=
`protect END_PROTECTED
