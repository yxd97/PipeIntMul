`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQkHyIgr2poFgZYNlISihCmUbFqo4e7k2PBraBcWVVlIAIYuTeGn6vIdPSUA6SSP
HeBQmi0bLRorAlkst2D0C0GS/vGJWfEVU2zp67LFbpbY/TymB2ASsb22KQ2gYOl5
/R4MvsVKPlwAsPeoN7QxcaJt++nkb5Bq5GAEcahvcg7hyLzvgceg21/G4Y8bWIem
3sEHFyxdVBQSA7TUc3/bi9/8tRrnVqa7SamHmE+iAZc+oKkyLnzfutenvgSFwWzb
On8mmBjew/B9V8QCZia5DUfSPNAGbtSKdiz6kNfTbED5NthxiJYiFjmC6bf+QcJZ
ULZ9WJ0lXZ2kyVot44lAnZtK1MrbsOtqOWBXgCjNTcfrOkWXYPOR3DkxRVFnePru
ZrxAcKPiLmuclXtj0z2ZZRTpLUlHzEPsWGYnQcWdb6YHOYtahbLXaZxlUzpdkTHr
`protect END_PROTECTED
