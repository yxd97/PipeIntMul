`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
70O+m+F0yg1v30EyYHEAAtoi3zufM0xDPIggQ5BzkH9TF4Gm8wYHxEIaRdlcDu2O
E5tWUCZMdPG6p451J2wOBEdpMnMxC+XJS+N/8SpIdjCNDHg1FyZKuAMi7MELN9Et
GcfGoRPd/uh9FdULFCArpYZu7IbF8J1UAuklhpJckmgiE3offeIRNbnE1YpS/Da+
Y7sRBe/mxh3GzBBFj2MnXEUTQ7iOLH11w52awLDHE9eDJ9qnjZVp0mF87+aRsks/
8hTknOUV4C9q15BRgOXpFXLtxiBbHwkquZI9AM6Nb0LY2zH7eNqlkAtFOuSYezS9
DjSQupbk0ZPdnQb7e/xhyFX2Q8/LB47XRoO+O118MpzbmQ5HrdksDRoNl5iNMdKZ
JugSQ3Jrqw/706mpSbpLhWmSW3K7dCITV8tr9LFkTDsW1AyW1PBObBICBsA1I1ft
CufgyJcTFBTeUkiwNCQ37UY58sdiLaEM19YhL3y/TQ7DgR4WsJX4BVHe2EA/KKvu
YkkenUx6HPbQueooem7j3xrVa8U2/QGJXLHCt17RsrvMJGk6Vc9wknICs0bvvRpR
H78Oj/PuAQvtfTos7LQSG295Z+vmG47L0i5x7Lk38D63vKnvwMTCbQGy15eH0dNC
cQE+v1GkaMa1JcQwH2afdSPIYn89BISln9A/9QaE0DPmnSAesG98aVB2s7haIbtN
g8n5MFWKDyPLv6C3Y+1NiMWFdEkT35Iqfarnba41sfGrkV6kIYrP6rAPeecOSTO6
WRvPGb4wL88d+P7KI3mYBz2ikqZuUBUKODKCL2CldTmgHUVXbD1L2UvirbJ8aUeI
Q/NFDTaau8ncPFVSmY19GVt5Wg4BOQsuqKB3TcoLHIR78fRoMwtoUd+FBI/w5Kyb
qLk0J1Xdrwx/GSyIk1ZoI4kHOFY1+L+EBvec5lwAIg8ypc1NKbev7hHiVEqbdPoj
4TFat6HxnpM2egP+LK4zNQFMlQMARSD1t4qiq/WYp5BpENVSD4GLG7Gs5VsTM43T
Eae8zQGCPBw/wUM3zSBlwfqFzn0HQmlPIuHvsv0tdA2Syqf116uljwoI97V+KL0i
CIFKTriGsVW1OF7iteFRQbAkUu0RkaLHs/Z57aDLQKA8bLdAh3VvTKW0I6Hh1AzF
BCeCeNwZD0Ei4+G2uuodLP1iGf8BCyjeonmjcWq0V7V0UaNvAlpbWMAAS+1sUzcK
`protect END_PROTECTED
