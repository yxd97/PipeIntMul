`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9s75ndeMZCOTulNCGhsZ3Hc9o7gpsPQXubNluG5HlLIui5fpYlEacYM+1SoHkHY
IVQfGIusV24YKcWcj4vZ7Sh+nsIDULF2bnONgQS7zQZMU6s3k1QKnVHPl7F0U5+F
lFi63JJhhEPOcB5dpZiD6V1DTF2E7lqqFtc4VvLtNgXjtJC9S+7EzuQbu0rau1tb
+dlxNMn8cCvjbgtInTViK8KmHWEQpIgauE0RDx0P0EbmJ3/KRM0V8vW/S2sXt/IX
PYT53RjeubtsVQcuOMkYIxlGo3zvjy+pfl4KDBzgCA7Ta8iRigcx7y38kM9iydM9
lQRVoYKB7Y4bJHZD+wdfqDUxS+8X28rFkPYr4lp9Qv7m3AgF3UahDXPv6HBm0Wb9
IHqa2kfid2A4c6f/zKG3encjwslnp/kprwPr04bq/KVvv2AeOvuU8TV+SSzvAWzy
rlD+KJ3txJI+t3ANNQhJHvJmR+btOTZ30/OPVpqO8Vk=
`protect END_PROTECTED
