`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d3clkY/Svcp7t5ID7ete62yFfmZeraw/lh7Euim59r5HM16ru+vvLbY8HSj0PQxu
5XbKZy600UAY3lje81mk6NYLcX9yxu//1mR31cIGMVWpw64CTXLghzqDv3ONHLk9
ekHBTmim0t4a9pmIiGmIUgi47ynrv7benoZ5GFAfFzI+oIhy79+w6bN6P9orUEap
9cXN/JDKuIqNwkI9pU6tUi5ElUxo/QnwcVjGNRdrZyAbiBSbgh0QMOHSbGmBIVQ1
y2zYf14HgO9lflaHHuy2dhDxKaP/N6cANlW9ARaSigejlHTs7M8fnWfie/iN+VQY
`protect END_PROTECTED
