`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hlb3qrN7CoC9VjeZDuBL0Xf2R+wzyKWkuwLOtEpfNhx6AAw2fow74lKDfOI8Zq4S
2TmK0cmpkZPnyhIQ51FGFre+90bI6sPECPWb1wYpRbZphg6Nq9W99+X4gRZT5Jcm
acbpCW2jqnpa+Om7mXqXcVyhEekfn/wjRTykJVNDILawDiWNYouZxwKilajKlm6A
Bx3eNZQCnZ3GTkB2sfiwM+j2e/QrXqaxu54LyMdp+fFZtEZKBRxrd9Pa2mDTm2NI
etjB00bZM1xnC+logfOwigjMk2MNYBi98jcn3TaiR/o13rIOScsjMv3P+uHRhHKl
sqLlOTgaVcHbou3UQmXEYMuyl90Hh63PEAjlip5M+68Dmjy9nJeiofe6xOjq6BOK
1BuM8a80rghb68DhEL0aLM3p0B+CuhH9O2Hc9v2Lb3Y=
`protect END_PROTECTED
