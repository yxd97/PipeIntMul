`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5Cka0b/IYS6yPZ2uHdjHMoHasr36BVlTkuvveNSGPNLCBVQAH676mFZtwMEGOMp
7NNLRtZKh57tjbAmLGvBg1qGcgYawQc+IlMfQYMsweRLhZeFGXtArzmKh3bAf5xQ
y3KYS1POpDtvNmMZ5i+wXVP0/jbyAZlZmYn3wJYwoByEIkO5KndlVCYwMXQ332Tw
nUsBAYr+kEnuuL3XtR6Idf2uv4ydfmO83R9nrfzHfr/AMOpSjGis0Pm+Tie3VxSv
y5o7/DHhNIXaQpZj9PocOv3m9WQaXJbwzB160wumCzCDbWybFelJYw7qerU/xR6R
bvfeG8yRzGT8UfC0ZE7GhoHR/l0nCtOuEyFr+D1tBGxCvFpwx4oTashBFXX6IA/a
KKi2yjCbfH4sENwctWwYVTOWkMQW6gAZHHpgiQq/RY7Jlz4JC8/fG+XQqXs/iEgJ
hYiQYqZtTCMHr/Dw36TQ5A7NLSzW9m+oyCjzDk6TKxbPu1H2aAgfVVugRr+qgaIV
aF2jaIbY/ftzKLd2+I0xFcHt1/YFIfqOWfHihkdVovYVewMLELi6rXup2ycTus0a
ghkmQoMrfu12eaq4Ks4DoQH4l9EkbrFlAr9zxTYfDd6y6XHzZoyHsME9J3B2ekxf
FedSp1OawrVAcwwrZNjQ6Kbkm4PWsuL/BQniJDsPAwGKGp1dft3UrUO9ziPkV2Kv
JeDWNPPYzVzkEZR95871ovSiCOeifrRdV4Xzfi0+LSPstKDU7ZsTAfWALoFFeOc2
RG8Yrecr1uUTrPudiROZABTho2yrH2E2U4mJ9xY2R04ilSTdqn3V/NyqzXd9mJJW
W6tKHY/1X5Qk3jggL13TQyp2DS0o3eIKxUWIRabgoyDIfAIxQyvNosSVp+CCt7vS
8O7Xoy2SvkgRzT1q6/nTmMxt0QZB+Q9HUaddEg26e8yD+p129Ke48snGNbiwjxrr
ztOx8LEfmme5dqfF9YMNdaFyzyH6rmxZYh8e4Ps/uPNW65iVIGic4wF/BuC+9ykE
v5zYY+PUOY5irZiq1/ePacwWfI/FhR2xZsfefC4swLuU1uvgiGGpiV0Ih0TpPrBO
R9IbPqlKjjIolkZ06EuqyeQXGuuGEfjEmVxSUGKGrkKmsL6P+c8DaoCRJ2Gc4Y2s
JD4aFssRDLaNDYwHzql4GqcTIVJXLdUX1IKwpGyDMa9xh19AbR5/3k4v/a6p1Wcb
sCCump6W+EZbjFoTeh2kNEuMedBj/HP+a/opgPSfrHXZzqn5ODA7ymyUBAawaUCk
M3IEUIOdzKIauXk9/kmFYAqVKFPEarJYZ6d8JFCd+TGPKF4jtaLCOv5BftE2C2lZ
nqsAX5WgA9UtMO9QbaU7nmZwMazw+8y82AwCAip25gJ1bbQZNEnfMkV2BCaSuBTV
GRN4QeyP/CdykW3/A21eVyghSa7COCf8PzpJLbTEltFt9GQPYVJAa7+vhmFs7bZD
1KnP0Sec05+CaWRkB27xs4StPe5mPsg0hzWERC+WVRyOvii5m6NTvrHh6O0/gebE
CAqLpheLvwh67iU5Hxj0lmA8F4Ml7FwR55d+PCYwPBWjmL3sBcOSprnBCk4BArhS
VuJQwZHQDSHK5PkM8FTX4Cu1UvhVTAoqd8oaaol8Hlzu4Boj8GIH2vHXAaOIfiTX
MFaVXgDLH/Ig1P0gxnxsebZPJ8q5OFsEL21QNirngXcQoPa7Covbb4COmjI8+wr+
QyDnmaKdkb/xEm50DTtt9O2BXTlBadbW4ldbGaQ2G5ZN8R+06YEICrHoZDeqpbG7
yWMafDVzKXFQH9OQ5LO6egiIcNrrCO19p75ObU/gtKMpx/Dn4OZIeId8pu/LquVG
`protect END_PROTECTED
