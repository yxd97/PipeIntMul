`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OykZtnJDTYxm4UnnQplFguPrKYZ9a8AgNLx0Zpl8sBSBvahhfUYNd287QJ22pmva
441zt+yG9o7CvwC6Hu8u0k1/4k5uRDS1h1hX+ZVyoQvjprTh/aeAQoPw4VNgYoau
+iz98gk/hTOBYiD/Hzgni/PnAppWWjZ2/vgbZm3j3dqjhfMtH+ozUzVYD5mqHQ8K
HyId3jIzLEmNH+qlRu2kjIXrNTTHCEs8xuPSqZXiGq1i1tWbimfDVMzR60FZwFcQ
iaaimz5dBVx4gDA4FTPfY/EMuhpTGrivJbdaK9XuKL4rdWFCyoT5gxXrxvr4cK+O
Iqxm5XGVbehBXI1MJXMAXScZGHv08D73u8g1nih5W9cDgKd2fa5o8bN7oywngxNk
`protect END_PROTECTED
