`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGBACHE6qHiNT9NOQ2BhpA8SH7JaXau41rncIrVjFNLMV6p2W/pZ1jx61dZ9rKVw
jx61PzMfauL9WZyhKznO5yKc2Di8///oRv8c02Th+EGU2hg0YpKHvaW6FPYoRQrx
nU90zKp+GAIXTK03F/os1fT45YvFCiA+aWQPUXcayqe5oU2GPfDTl1kh/tFYu2jM
J5vgiNNSd7rS9f6fL9bFJP71OiS+aGsarjxAydWXEibK5Gem7VtTbq95KaaAQ7Am
7rQozt7kqbZ0iUVFnh1WW1NI5xEYuM1K5LXkhwFJBJLuI8eOlqOyrK8ZPl8S2YaK
0eqR1Bk29n3fgpQk6qtpzv+v/glgpkG8icd62cWhyDTvVeX+ErLEhqo1f71bkwsS
/3IeCyhL25r4gYKmzdTpbIKhct9Qht7zCT2/I01X+fBpnDopYU+Ap1BUYLQuEFST
qjh+GbUdqkJmV/jXejdvvhIaqml58MBSiKVkMqATy7pGhKKf4hCD18Do8jndAD5j
3INuNKvLimE9+piR62KdAGUoVxfXHAKBi6N28hmP5jI5gH+S6jZTxetVpCdcvffB
ggbRMTMPXgQUggYR4E0KVOgLXAT0pVKlisSHZjNfq8eOuWsyL590OAvIH7Lv9Ti+
TZj5eETIzs23Z04dW21CFmQv5FsRmTAI1EgiKAa96mmKwVZvZSLwE18a6l9VANP5
fj01HrUXNYlla89BR5hWa2Y6FDTdtOqFyvP3RVtpCEooV10xJ/hzfltg5AqCxnoG
Q20C6o1q37BI9KRsY7+9DiW4rz+rRlfFbwn0H8Qt/o1QYn9ixLLD36B3xw7eXYx1
U/4dY4+MyvqIk1xbeB5BKQ408Fgg5fFpudHZG0MwiCu7LglD7yjjZ6yEcPrcxyQs
3ncgk9IwnQybNVUXzvnkb5E4lAEzUFvyG6skxfjPzEXe2g7H4jIVmSFclvNUzM0f
w6ZfkJzJ2rwRKavPa2X6aMRg6uUr92AaJwM4nx63hP37VvC8b5bM6awiKNZfz0j4
wTzBxcStTlL+kxKF4bSanXUTaMI1K82FBH4f5B69fGDIKBQCokF6hzLgVIAfNuo5
0sJ+kduiaz5tSo7w76ec2/jO4Pr3RZaV+/Z4Pdhhu5BKqe8HUEKietmfYz0sSY5j
A5cTUpMiOYMMMJRuY1+vTEvhufSY+EjuOiVB8IUGE1GX+1UQN4pv7urUfZiqqePv
v1fJqfADqlRW4RIivksfDtfxWT1MRdAWg1JTSxL666d6J8L14OeYIoOCMVA8xwUd
lCvPYNBXz7OII5CldHImATyMhzNSaisQoMpBd/azycv4ykoq7cDGiu2LK9xNbSnY
ERKdWLubuKTcFxqSmJ2TCDIJfM0SnaSVFvFtvu8lx7bW+X5IsIl45DJWFCE+JJaO
Bf631F+J/ewKYqZ01dABywH+qS/Ugup5N0b8q7NRgT8ahQPObaPLUOTxRKqH3lgk
8BghDnFvTY+Er1hOM0VvgL3p8CvJRawgTkoqnS2cHqIBQXeUMISRjdrXvzpUNxUL
MBf5WJ3I2ZuQxRho+G8wlybzaIJYIcgRNml6JTDP5gYk+8RXrH2O6WgyqOAHrB8Z
14nIKFr8HXxqIiVEheXYc6JGL0MfpeGQSAmrAPdGkGl05Mq1NdrNdlMqq5R+Klvn
Z2flIC4p1mBUHb1WwFqBbYwx9sXL4d5QaIbngp2Ou5tqM+OaIVQFfoE3NmYsKNBI
oUdDlAa4DJxpGODJtOcBxip9RH3eJ70pTwuIK7o/UPIpNsImSmKd656WgV9OnmwT
+2P9PFpcsXoQU0mO+jyRM+1Kt0n4dNFpygyuCxDXBpl2Q9sLftqY6Gm3/8byTtoE
2iuLnbXnKLICT4I8a94IaA8gmMiOdoL5K9DkEV1n2GwlIBtEfEqVB2EbyRdUBnaC
KECVeztcZvbeGqLKXZ9hg5rU3tNp6tpZq0cpMl2TK2xFMplVRmxZnb5M7F5TE/9U
puFAjVqKO0uRRRLpC2KVu90kdn+4XkoccYg/Rm6YOx2IRklxp54ShYjTqkl4gBL9
/28oq8QEELZOy6i+VU/jz/R2HCG6E9hL92ZNhMvmWQqtfoNHdAsqOnL+4LvEQES3
AnF5ky+4LR3kbdUb6itwPlEuMl+y152XYKhgWFZsguzqZY4pGgfb05GVX0k4JBbW
U8NllWte8zmuSpHdALI82LTQ2pB24rWVN/C1KzpFRCTK6LLpyYdZkd1qAJaIxSjB
Fe/gGPGNZe0vdhMf58BTpOQEBFxHVwXN0dQPZmAKup7nTM6eaH0/Uw9C03umJnnN
NWwErpKbO2Bai8wCyhygpTgdjj3If/yo90JcWqpW90eel1OshYIBYJl3bgN3/ycc
zfImMSfl5/kGfJlUI4FGQ0m8KiU3wdK2xYPd8Lk5Jg+ywrm4Nh2Lw6g88VRN6HCc
soCwk0ZHTr+Lz14SaT42VPe14/fPB0JdxWAuuoBt0W3ttJ/mDRMAwdfTpMoh57iO
sD8nV0Sd4jwmFsU3Soaydxo1q8gXHA6HHQq4Py1R/Jsv9A48CTA6RXRnB49XFIDK
ix1NTm94Qk7+AWadYiCIVx91PJqmdto93VDmcsc01ECx1cNny/zEX34hU28nivrg
Oi3xN6Qlq84z6IROQu/lRg==
`protect END_PROTECTED
