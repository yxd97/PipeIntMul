`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qTyOyI2iOLqKYoBRm9hv5p9eW2DjUu8cvB1VGthDF+F4LjtxGno9xan6al7Mqkyr
KxVpFoOM6J1avDSk2UkjtlbdzZNJ3+QpyXdM4rrHXJVBqJIYff3/FM3F42LgCQFh
NAIdSdMKkJKTX8F0L2qPaIZveELXXTkmm14Dd8h6S6Y//mm2TDHdPdWY3oXGRk4f
1jpVHIwzcwbmLP8cgVvss+IBINZsF+IJA/KIYUKQHkUZ+iE9sj2e6gJBrG3xMVq8
RzKoj/NfNbZuMA1hrjEvHUbxzZxFdd4pktzwnC532Jx/T+B7oUHPvmAeQZ3rsTrS
pD/X6c0YRjDs0INv8F0Em4uI66FrrJ7Ep2KOsP6EF4euHCUDk7BFJbT4yRUX1qjl
OBpnCSefFviQsX8Qhu0yVKfYk0PvpA6gaTNxwlVo9iJKSqw+upOyojdFgRkQm7/n
3uxDAY3xcewCGBDgwPLYXNZ6O8WOi1m2ee+OFdtsXSu34l8SLlHChUUALe7elxKw
sCFyiDh2MIZsy9z9Moj2NutuypD8gA3Aip40HMbf1DcOr2CgJqF/avyo3wABiI68
IYl12adfcOOTmjXrME7PWQ==
`protect END_PROTECTED
