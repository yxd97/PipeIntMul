`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+l2MNGOc9oipynEbTvr0E8ZV+lZOcBOHhHwGs7Mltp9fjUB8ULTyQL++kvVXy3l
9H9BlLKAlRNSXIWxCOJC1Y9dRaVX9TRtu3OZZITP0BYfJh1URGn3mRwjXs7qWZP/
Vpl0rg0Fmqfy3isUqRv+Zu26znqYwFTuzv+Zgkh8Etx2WOxN64lnsTYBvkBP+MjM
KM1sgvb/ZEG+h4CKXDpXWaUSSTYf8W8RRq650IfhjVvkeVPoCt0MQcewFypGJge7
gGco2QJjXIjP3MBLREYfQiibEE+/tRXn+Ythho8zvqcYaGwEs7vLeSBn5pXrqNcB
Q1xIr7XkH1KREBXI2AszruNcDBP2GuxsXCXMO4YM0EEP/lpNNrr6/iQXwpvPJJgm
nUUPva1xxY1hAY5MuqRiGg7ptakO6TQfZAu4V2M1JmryOVQfQMgkI5L4nXlH+gYk
ZMcaRFAW3Rpg77wv/mH2SbCLclIgjhHwD6HJqdQWGVUxPv/qL4xsjoJWMzfQ97xy
`protect END_PROTECTED
