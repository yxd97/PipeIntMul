`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AkFO9D/5zxcibSxrugD8XpmRkm8XOzMaIIxGqTrh+T/iNGjulVYvMkoCRbuaaLuJ
FUxoJhRpQaFWa8WN3ZmIyAVg81kD8Rquh4aPSO0g0as017Eq+nKL7QhIVdRQjQcj
9gfilY5u7SAyjYiR9mYAh05rhH4DZlp+8VZyXhlNU7Nd8taSClHc82GzPc+0z8/b
E2BaDTnNyQVj4wdO22gnNMYKO+XSJUBgyJxY09TSGap/CAGNM3BwpPOMIBtUJ51n
Fkg14iv6u5ZrW5TQU1mF9wWOhZyn++YR/yPGahYtbxS7S11/QgqOLN7B0eLq61lC
A/jcl36x+Gd9Q3ptb82LLNvZc9bl+THEJXPAyBJg7vVyQ8JwlmDBMF80h52k9NN4
QRod4E+3t1Xjdd0shFeFd3fPY/MqZhq7fvHzYJdeook=
`protect END_PROTECTED
