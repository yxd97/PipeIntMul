`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N+77Zlb7PnpWPa+LwWBvsscAd6zaeH9+zjJCLQwo1fXxdDNrcz27a/NET4YB7POd
GzjgjJkv3m+ym36BF1ziRQwwVSZJFT7b95QeXIelsczGRFcHg6mkUN7xBAlj1TNY
z6SJhBJ/htZCYcCGlykenBWaKY0nbw6DWdOggCJZIUXq8mv/SlMhzHhA06zV6XXv
boc1NsRPB+NGSzdQbbrrcJz5PVzwSJYLFbqNdwDOYNCbA+WzYDjmE0bncyjaHpzD
VRL9w7CQWF+0EPQC10mo/xt5Z0AF69IJEiQKRS6Vu/FjJEFrubWejz4DiqWw8zk+
ug/L9zP71ZwIA8382muXNzaxEU/zdWCcimHsd5/uKHeSCpH88qdFH2rncW9foVjO
8bNKl85JAOO1VVBLZsFcavqOmSuPKIcBy7qybJlBx9/HG2dAvoH2jOrEMPw39vZq
w144tkzvYVHrFiznyF8hCwyx0aKy5mw9theZFeoRaPw=
`protect END_PROTECTED
