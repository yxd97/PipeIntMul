`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r7XF2Re+ryB9WxmK889GuuR3gVH6w19vlZ0OM78E63N83Kdz0XYPASwzJ1PxxYSb
6fDJudxph4qv45TxtCsk0lnJZjJb76pBJ7anDdfz7eJxC7mKQjYLButn/81Uo4tV
NR0YqXl2x09AzQ0eW8OlY+Wx5fCUxRmYuJybPLj0mfYPchMKG8pD/KXiCy3VGku0
yBvYHXKoOAv2Mp/qaFV+HphU1px1uVCDoc4oXmN77qxbPp9j6MYRzIl2C3OHycGQ
f9C67g4HyACkbGWgn3lRdOiN8Psf/UbxNcMjJY1jXvbwEEf/Ft4DOCchuLYCuEEi
Hm5v75Sf3nxEqfsl41oZ26Torl3vU9lw8UCnx5xpb09vIeAUM02fTRQijZhBs/Qt
+rz9TO/ZEabMdJsy17eIOWpOz/rSdXQTZ1kAHEdmrUU4eJfdBAifuUc/+vMQYQLJ
lUuEqU9Tj6so3nl0f+Bh8RffNCRb5K18n2vkNX8sDB6OOnPs1zFhye0rS51WzzEf
faUtJ6Vu0Us5hkg+nGNn87d3X83imjYiPR5qViakRa0cCv6SqI/FNFw0qqeFAnE1
+yA1RhYRhq+MSl+0ZHzY2z6gcEYNM7XyPZPAmL/96uso722e6dshG1WDq028iEX1
LkRCYDH31cetTQsdXRCqF823hocMnbOC65AhjBE2+Vt5MWS5oUkEnh0/rYXICqcx
vAxeXXptF++A/IxO4UL0amacQmQUXWTwyDn/Ylz6bqjQqn9u/zVaqOztnT5mF0hX
jj7+KRrt5e6wb+SksWdUQnaHr730BMrPP6o9vfZuh1QX6XVcbd0BaFKI/+Uw4+LI
XbohRtNGsUzW50JZox7bZLyo1drEd7LN81RnkBIXsTr9lJ/hIvVaGcehXzd4MJdC
Lrvu5pBZMa0ZkqnJ0OCaiMIE/CeFuKzgEbPuzskh/F1YuWtZ6Ek65iybKi1RxHoU
khJRBYx7IaIa8N6uvhUqrpYIWLwjNEP/Dr5sAlYm6QVkelMW1N6wPEEo5hFi+y2M
UkXTWatUlTAeHNyX5F0bQuP7RaG2FVJYU9P+qsxdMWA6jtGNfdoVxJ0UECuvUXmn
I+QXB+G9HaFBoj1kDl7fT43bGHbGaJa4RjfKEpxpuIjWOsbRxn0NZgCCjGF6eqAV
IoghmzZ5RRmgYMJPHmjHGGxrve4VmGHI8huLWz5GYlriNOoqkLUK19KcIAtruM90
htbWntN44RxCop3KExMO+R04xR/gP4406sG5VZOXLkwr6IDEhiD3Rx2PNrXXzdvz
cjVYKfmmyrk7Y6RHnldnBZoJsaMXuoXcKtlT4l3qc/jc7WbI27LUcHvewc1t2yQA
RM1CYlcptATUzdkDwIZN8u41nHnvZ8azmiFDWogIYDZHmQUtGVnJdL7pNd1T4O/z
IS4i3evLH1h66QWlYBiSinFTdIru41BxcP2uFRW+iQNJkNO0sz90WQ+RYnV7YUJ7
O0/numNg0dRaFHJyKDBmzuOwd/R2f4+817krBDeztpqhMcN6qW0a6ii2vFWRFOJO
VFucJYHoFs5fm35J3H0DeeMxw57M18N4Vdke2deAGHoj8wE0EIiaIZPcI02+kCGm
gIAkRBWfmb8NbFkOdR0ZIJX0hgMWEk7n1d6g3w/XMwxvocRpxY0KITbW+vj9xzr2
7Kyv283tMQ3ZRvm8KLyg2VkM172comevB5zpH8/Inybb7W5LhgYgRSqG7PgHkrp/
YublQy4GC2RFAKs0jsODwFzHJmFQcbLg5nlTaoePUEY=
`protect END_PROTECTED
