`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7JQVV3WrEtvWjP90iBTZ+prCYq2VY0fwC8hsk18MF6b6BMB9hPJsMerQNVQmy2cC
TaJrsnU64bRrkWaJYsDnyY2VDyQRSrjoTRe7WIAG7B4mMAnaPzTWyc8DSng4T5bz
777+sUyN2hJYo9FEexleEF4AslijxxLtSzt4a2U8nyNytkCW2w1mu/efYLBRVUdJ
KpbeTzQGKHx+tHRz8dOM3/7U4W3f+CWh32sCbb16aIIaaBtxdnCpU5QIEoFb0yUb
MmUHyjEnwpERPoKZzDn6xQ==
`protect END_PROTECTED
