`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z94GQZfnJrc6t1wOT7Uh5XNYxMo3qXPwbjKR/spq6IOcHP5yWPVhjypC6h8fTbF3
TNi8JIRcU+UUMtHYlRV3a50ZXjJJTEApMS9yle/gsVo3d4+d9oRFjMZaoGjlJ3AX
+HPB6W1/2IGa5DEryjKZaMoLLAhu5JQvdSYmEHgTT0OUR7PvVjb27C/OaMkIq0jo
upQA4rhvgQRjB/rMjujBnnTYSWjvU4AG2iDBzrvxnig62uvCsOywEWJwG13o+2QD
wCuzpC1EZq4i/5zqwIIJcAT8FTh75RdJJn9GZKkEWBwZZ6NFcbVR9iWTOc41li2X
JddhE1opVEVqTZ+kEWFpSDkZe/VfeL676EYJo2TP1Fvd+P+8Y0TG6RdPJKsxP/qX
ITzHW/XTpYXkIrMrhuRMSBJqezsFffCe+dVOYi/k1ENSX3VfWlBTDdbmY/6lRI9G
ATo6sn6D6+kan3oFDQfnP7OeGEH4idh2dzNTypT5gUemwH7cgVhNGaJZ74YjR+GR
qDNPAUGV+OVE05gFK0K09AlDz4FHL6Xcso99m6VUMoAWnnwmxfk52CZSSysFLd8P
e8PD0asmCBLK1vr3DSUzFJKgU8H6Xsh/YUD1pFpqwBI=
`protect END_PROTECTED
