`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DkWi+mHwKlzP2HrVJUM0CGx0A7LbXGNMcx+nBfTowIzwC0pQBBHFWMh/FTci7OCW
dAV62Xm7j7uSuUipdENJIyKktGOBXToKhVl73qGAIlmlOwirwQcgjzwujpwaK+0f
FChdCyaUkUXJE/jsQ/v/rP79de/OUE0KMWwDTSxs5XSNtM67EeK4X8wKci1La5/s
hbjy3Jp+htTErBS9ZJty2rF3Cdd8CiuRLo1yU+rlfWSDggugIiR+VKLRxdpOW7So
mpkPqTCTlbXmnfUA0bJXqygIxYSWiDvFTCgLFaWMyMGRkccHXemp292Fkbke07TO
Fb89lveecR39ixO9vG9mJBJ2q6fujxYy5aTVfackgQh3pINpNyTZ9sJXp71YAVSp
VZpM17dawpC2GHmdR4WoxrDa8Mjjy6fyZBUd3Naxeg7Nf3YUkw4atMZriIbzUd7j
xo0O4nS3j3zkZYcp0GIQQcxygGIJD1oUTwkroXscUyUDfhfVAHYAFl/pgnI3a+7B
EVl3gA8WQZoU5ZWk8I5Ya6YCBFWKG4nUr8NTMciaPSwbL/2EV4cv0/1e4ZMpDxYp
Hq7iaxa8xGgazUAsV/PBjPnOl87ubddRLQzBc8HmjMtrdEAXjpXe8ggq2W9Iyo2H
/TcIuupgPlrZTeCtoMf8nCkwlW+tMEECo6m0i/wsE5wLL7cB+oUXw3cSuSQecpAQ
3VbfcVyLdZPmV9kjA8ai9j3loUPKm3o5fisLN92yKNrPUy+UQ3kWtJ4jV+4EkxOH
3zsOexP1nVAt+rdmMJEnXJojdrcslSwNynSMvV7ONG3a2R5YPt/BFKNT7Fq/gpkq
e1SdS1MmK8yudctC12rRn3w9YW/6qdXgZstjK+jYBbdcRHzoqlXh+ViJySaSGcPz
euZU6sxfR8DazppFWfZtN8LK2caDSlIWJDKP2b4S7k/nhg/S31JhZ+EWAvPVrv9Y
g/k4/+rwVbHtq+3YyxngFm/i9tNlAf2tixjgWvDXMdg=
`protect END_PROTECTED
