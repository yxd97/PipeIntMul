`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMO3lvAq7HHwbc12dLhidjj7mj4sPR5pWmrOqoP2ex1l+6eTo4oKu2774WdSXry2
60pDvmwf72aA0yJDtrnRy/Y+Fj/2nsSlw/PJqD6c0nKYF2BYZ8pOWKYmOQi6RmOG
m5PfLTyu75716+Ux6asms1RntnKvYTvp98Ai1jUsZ1wJTdxhmsnNEmwvSTimUMg/
TDDq1+JdeYjifDXRjJhs2xFesH21j0oJM+h5i86z09p9MIyN3zm1SqnfCDGItUh1
L7gjz4nYvDY+s6yfU6NOscS68DQznSWDQ/Y0c5GAD4LO/22rGyEHGjto7peXDdm3
LSITX8Uswcy2lSC+G4dswXwJcsRNVT1stJg2Bbso5tuq8Kxe2hEAk2Nkm9jBjzgE
UQruWX4F29V+Qk9Cy3U7xaCH0fhUajyPZptnVQTYtxmWU2RIVw3pNA1GMR4lDvjv
ZcQYpGqA22DKY6cXrd4l6w==
`protect END_PROTECTED
