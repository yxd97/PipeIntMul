`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0s2HPCl5vXMIHI8gVkWfDhwCJ39f9uIvfS6Us8f9B1SZIAka3jmY4dSnuY2GiQ3f
y0hIdQWYe5ifZQumAryj2hm3pQ9RkHN4pGtVogfVOLGiizPsvu1ImpiJyVtYh3lG
mQrF+q5gLTtwMuOa/fViGSOYTZutETHw7RuJxMzgZCDbRNHrOleoUObzHQJaTN7R
PPzFSo9koaUPvhi+5U9/M41G3XiFpBjEJZ1uBgdXEVQ/gB72QiU85CKTsWqb/alF
EOYueAUMZOkIJlvzDLEwUIqjsfaVGolfZsz9xS25NR0g4tJc38k0D9vtUlmuCPyk
m0/ao/Nguxvdaz9fNQz32RBzU4ANjVoxJPoxgIXEDk/wGij7pJiUAYdimJzLMsyo
BviXy5js1HccUcjAjn7XbjjJ9MR9wYdsrofcH/cfMJaGjzg3Z1Djje8dOplEYKlE
b3l5N+ZaqixaIir+CpsE4RT4LVJ6hvIHCsLxNwdbVRMZFAAEeJI6WXQuCIzzKgTF
Q01jQlU/X4BiEqdafWSujIp56MTTE5S+zYpnKUB8bA/q49ckshW6zR7FfG/9CjV7
XjuWGWnK+2Anx7qJ/rAcf38e1u/+LnO83GqAD6jloGrqLbTVWdb+Sf4FbuUGz1Yb
svtuKLVPCDQR0WsQZ0XMuQ2a2A5YWRjIaghJlsLDEAqea/zzN6VU8cPjHbLYdiDW
IQVrh2XlHb2W1q4AvtCbgIsbL+S8YOh6MQsX2p36BbmoCi/ySGVgIaPSdQuZ7ZX0
Ugd3paU9d2+PaXFHR2VdYaC0ULuao/q/OrQ7pSWBboXhrfjp75EfVdfoUID3b6ok
GEXKZesCMgDRPwPnDjfG00qSmWfGwUNqxYp3o65keDNqEhrSCVMK2Sa9daCJYuYQ
cEkzXghizulG3Og4Zai0v0DVgDvjuLRyJPxQPgxwUIiWtXdAtMf0wBhGW9gwA2wj
1yzbWcRWKNlZRACOCrfQr4N/QIIDPbYuw7phjYFiq6Cmmu6E1VtYOdjAXZWHjANW
3Ri2P0ruI5zD14SXz+zn4nQ45dT+P5pc2T69hKKXqQSR7xg/2Yh5gdvw5eNyquGZ
7eAayTYh2M2puDCP4ObxO87Bfh4B3ldAIGMPxkxNc7k=
`protect END_PROTECTED
