`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NADZ4cRvlDhFT6jHrOZ5GGEgR8T6v2FCD3NX6KUlYcw5MiDnE3bFfpxtBdcA295b
Wl/dIV5cmqApG9uaPR+rOceDB671rQn8iYcGFNArrZDSWJd/NVGfu6cAbGt8JGbU
uvoyoWEdHRXEco5UYrUQhQkPH+gjIwOEPLveWqFhbjYEz3T8jAt+f4y9t8YdfnvQ
AYvh5196Xb/WtPRPnF2wzlWG9rynQL/80thYV7LMOS6QD1a8ZQYkb7gvMIsJAbNb
tzcCsXHD/y3MMGrtd82qbw==
`protect END_PROTECTED
