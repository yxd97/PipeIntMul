`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b6VqFuuB16g9E4NT9TEFeptL8CuP2Vmh1WT5ANLZr0X655lVPl7WpYe9Z2IWMo17
8YrAV0Q1+tDE6AMh1hZ4wfoIVyikbxt/R/GgL1Hzw4+Zgi46oqXNuUgrO+xcIH3q
3+RWRxkhzmlIuh6TBC+2YQDKsBuPFyQTEcpz9dkZCcXZB0mrlF8KSk/l90qf6KvR
VAgSQJIJ4rcdUu8VMRH4/8cdA9cSKB8BMmdUBxozPEyWVm6Yhi8mxB7KBoGOmJi0
1SrqSzbpJMxSh0cS1RziJHp+7d2GPp7ESNkyjvk1pdmPoEqVpg28+tbHzNzl8/8+
jwuJRUbHtWfiet3MLYYngRn9JsofZ1KxksmAEENxXouEUSHM0vNcnYP+vo5i0n7z
VfV1Vp0QIvORDtwBdRtyhcUroOzwbndGNSX2HYAK8cLefPl6LOJSHKkvRLG9EzDA
aSis2WU9pNOpLnwqY7HJLrzsJEcnwKxZw14vMDAuY95b/v9t152UHjgnGvNlfpjq
/5AUnEvpLUVjeGn0KO2pWIUu6I/8RqPLQduG7q1DZWuGs+g2xZ3oLKrlbIwCLwsc
oU5QBSaT5EOxM3XnIa850FqoHrSbjmzYY++xKFve9FWXVLV2YObtfEzvJTchp5Zf
SW/aiLnKHQ1mRwxEz1jA8k5VmorfAPpUC0H2AcCfF3TKxXtyJZgEH94e3nI1FStG
cOigrQeBMtxGKAdXVM0ykHUZdICM21+8IUclfrRE4PITgAtJBQLWK1oLSHGeh/hs
RozKSoJNc5RsyRq/JH6fqIc+fHpoF3lsOOQgmq2BQFvXwp16lPqdv7FRjUu9Mirg
hTY4ERlpPJkLkgAxH1D2HI3slBtZmg4OuI5LUtTt17RMPZZl5+KYnbjqnN+XSkto
ZAI6oqlCJAbsvs8EwMUlZ6I/+MmrEfCGIiYfXTmKAmYoduaTSDJJbFUVQd2cezLd
AUAdbaG7po9v9uBb6rbJ//o5V1fvRtBnoOlnHGX1Yh2L/VAkTpfiIc46RjJYC0VJ
JzTJd2jQ9YJaJfc34b5gUj/25yAj9kGNxHm9w/WzId+WifrvW4acRMgg4loUthNa
UHapPGfT8Tj0AI7joXB4GL/3MCWYt8tlDPuItVJQCK3+H5MtIFHDXiXWQGqVhSVI
bH4igCMIXGoPyN2ap5gEYpI0Vlpeb8NdMjK9Y08iQqxqhYQknHsXvuzLqn9qTXTn
yIdFNcrtDyJVmWtv2dO1NRFNPcbA6e3GmSM+tX1YIXex9bUmY9ekwPPE/gOpr2nk
BGD7cc1T7lsV/X5u9c7aOgN0H8jCpxFf3ABpNKH4ez289oUs1jkI1V2WwgUYdVVE
mEzkrVBflPLh67LUuoyZX7ijJXKedmxVvSqaBzSfIljmQit12MJEbU+eqfEgNXe2
XBNNCr7uqchbtXNPlmYHe4/vdnu9ynzYPTT3c3u0rpIkJvZSUKwQ3FVbq3tN2xv+
uAkAUfS4fYSpH+axZ2hQX4lLSPxrrxbj5MhbshbfVyaaCC0hEf7Ob7OxlGbrf7WH
xE4N7H9yGOAogFvQPgiVueg6zIw8F9hg6v+wWJmK73zrIqeJQAMQPl8xT1+rvxB4
EYOPcT69oNWOqxLcA92PgfTvE5CIO+K4KZd/BlQM5XyeVZQ6EbmtN0xcdszHfWZX
8Gt3IUUe+EIsctQhPdUstVDg6x4QgfPlWwjQEajJBumX/QEXQq4L+dHO4uaAx0po
6IN0UYRZ0JYv/XND3oi6D3TZEEgrzyQVuWVY/VFGEjA=
`protect END_PROTECTED
