`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x18zY1tS6REvzNYqz+LCIqQcnXfgSD/xhdu+efjj/1zsWMJ2Hw2Dmi2XsOYzHUN3
otS9gtwVqHKqsXsJL7VHUbVwj9ktfq2FLC5TBZIMFotmCJXxRcOwJDOLPZM8q5NI
dg+uksbhgBhAQtDXHggMLnCpcwlCBtFhNyaiGlykCT4oolYQ8ciYg4bkn2CL0GDB
zwPgk11csaPPbGAi5sWbDnPIQ9ML7Hv2oLEnpYsNOUrIC43/4mjYJoJ7FgfefZJM
9sfb9MnmUBZaZeoNU/ulwAFCIVbZqZcZdGza36GMIFF4Ud1klH12LnLqdP9sWbsA
AL+jgwBZVMlsQwk/RTlWQsc010x/BJ7NIlyI0FbVoqxa8dgkLM61f34q3lzV+n5V
5HdGFVNij1OB3raHDZjc+Edc1LQTwxL0KjcbKJucC+V6JDAFDZnG3byGPUQjipSH
l0fz7VvAa0JAcCUWFExttZve0WHNaorX/WgaV1I8xMQGSg5+PLxrVxpVHumQdoAc
`protect END_PROTECTED
