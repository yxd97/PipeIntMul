`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BzIclT3RmuaZPBZskz7TF6ZK9VMZTgBGbBmtb5mgiX2hpC6IrBOmcfPXKlSrHJsc
zUXjqU+WQ9Grrl+gMJlOD2MjK/In4yEO+VgV+s4828y5hLTWpeRTraOprv4+7j5B
7BOT0C4gvbITTF3yOxmqrJUYEfHFUcCamevjJJ3Kaw8bR8kM/FyhTrZfGTHmvbPa
JfCl1Caa3Fapi4qBmYmkz1efULUjY4h8EOj+65+c+0N2UWBnN5+5kfC45gws5Nuw
7VI9OZpvLoXqPuTbI2qjyaKihqr4GxLusMir3BQ8cN8tV/uCnihe33DLWYZEFDq+
u9lfpBgMkuY8TQk9bPq+2+ebkr6Bb/d8FyKGQ+7z/4V2g5MK/tenxzRzDfIG5ET0
nmUY9Pktvm3LptuuokWWj6TTzM/E70UZAm3cxjGNSe35fosWUCtPdaUZZSxsBi94
`protect END_PROTECTED
