`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RNc/b1CA9gmciPQleFzqH8BceHgKOyCTD188Rt1wNeK1HocGqCzFk8qGIqt+e6z7
PqccKZ26LeI0EWRS85/KnaYjOqroiEztRIrM820HgS75t1nZQzpJwa7JkW7QMtAb
3nf4Almg88nvw1wrHxvJyy3InZlMX3JFAtHrOxCpJUmQmhGQqIr7mdIW7k5b/PMr
Z1BlE+Y8F1jdmWxJ8AlCUv2J0JaZhAqaCX3T/LFLt2FDnBuOTJw7dNLeUCyOJ6+s
yVeiiqoHpsC9fNSir7brtp5vifPWijP7GhS7m+bCyl7sRbcU8hVddSUDTufKenQC
gPwfouTeVk5zY0hJ/FFtNbAbrssgoZnjB+wlC3FB1W2f1qP+GmFJF91PJ259Z/N5
7q97zSE99zF4MTgCnJaTWSBa6sjLWhnEDHlCqEP3hCRiqjYfaqUc/XeO7KZ10BdK
Q0H3qPW6xqDGzpvbLvi9CcUtkweT2pzlYnTud2U1ed+vYcuckRTL7J2YC7wJwKkp
wEMKuZtEi747lK70MCaSRn0pkazJoHTgIaiwM/eGvV8b4gtv/RBF9XKYKPHMh0YE
XdWVxPm+4ZVnHESqVDRZH0cfuFghFPeuzSpFaUAmvYFulnenQYsNJHljw8YUYdIb
7QC+9U7O0xrd4QJw1PUbWE7gmYoB96FzOuVTf0lffqpbuvoPq90/S/k8uRc83/2J
zS2Q3k1SYRLNhHaziVm2hw==
`protect END_PROTECTED
