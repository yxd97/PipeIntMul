`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
paLf4QO9+u8aYeY/h4i2hyLsu59IWXeRiwJpxiZGor1QzQ5aj3ieeGAgFJxPoNBL
h1d/ycbU1bsG2bz3PjHOyMSQatDjfY8SsPyfENe7A2Xdp8c35kKF1P1/e7Pslijc
1/kbfreTIqvpTY/sxfEACY/qoB7nKc5WGUDhJiXcIE977LFARrRmTdtfQrAMBcoM
4J2NOais3oFC4tXjRt+xlRJ6x4q+4x8Veensi2qh5yo72hpk7H2h7BT3FAFpSriM
tL0buymIkH+9PdT7ZmT6HqXXf7n/TBeNDFg9LpsIJ2hKc2fMtN3WjpXzZNauXijS
uL8P0XRQjaxHQmOv61jMWEz3CQyAMZg40YaGQZYnADldzEMp6vPUzYkrQYmoPZWd
ZPHzxRT06VkOkP/EvCEoc6RwtVWM9kADexZMZx3vfdq/Za0kWS7LcPlgmREQxZIe
0pwWJ0nvB1ZAeUzrPDj6LaM8h4AYk9bZsdNg2uI3jFk=
`protect END_PROTECTED
