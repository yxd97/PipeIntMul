`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gkSen+UprJpgXl+wa5gps8pPuaHnYbmVcgZsns7ZxH8NWsSnJf822+aa45ppQX8u
KtPIFKSS7WwMv5eG7h7cx3jatOmpDkqqQUCZ1V/sHThnAkVpVtU7Dk8e1IVaaGMV
Ppl0jBc6w1lSPMvV5pwKB20Ly0NGfgpMvPtieGLiwtsCeCYr2Km8cJbFYtwhv36T
VnkgJ1FPpgmb5AgINR2cZz0xjfEcdEQnoORjq4EudwIHvU3V5teeF305SWgfuAx7
691+b2Grp09q2ME1ArdDWnJT5Bo/TDFlgYAIeGD1j+Dga6QqvpT2gKhuhN+fBU9D
MymWHO++mVvv+/goWnwY1j8CKV7Lehf95Ukxt5fpfEENNt7t+xGXAa0/5jYc0hsV
fu4GEYe6Mt/dSGCp31FEVZdCJkoEPxR98VEZNosMIYOOjzSjHfs0+9Jtj/DI5B3W
e0sf9bP6u2sUJRQnWDph0A7YiW1eGJr5ExgjJPpsrDIvaMRvMdamfOebnrKvvRLc
x27sYqEEoEgrcsC9LjR7Qyt8U/cINK0XrdFZGEwwcp9TG0yNocZS6QaeT2Y24/br
B/A6BrLhBo2Gdj+QF/VG28qNK4Le9k9ywH2CkD7ggOmz4Yiki6Cbhq4yjkcWYUGv
ww9dzXAKIejCwYeUyTZwvlwES79vJEX2e8lpgq1NCNpJrToERJw325aIAVlPAzD+
2M2Yb5VHUFj5S3S9keuMJMHR5MjIJ+jLtYHn0F2lWBnEF+u2PHKxTczuZmHeoiVa
BCUfLZY84Qx89TVK/gtdC6QliwN8lGFKQebwbei1bZbxLrrvPdBKfl0rcD5M1fEG
Sx8UwlB3JXmPFjqrTM43LecQN0HYW7SmRbzP8SY249c=
`protect END_PROTECTED
