`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+c/lF52w9/4+DIu7ApYOsaVPTG+wiJiAvlYebcBno3OgWDq7LMMVYGnpFCAOPkqx
RrWxhD+fdL5j/E/3blQGA0hDTaciCAiQs6A6UXzVg6gmhikSiwycW7/hDMqaOSfb
z/RlpeTM6ek6A5HxtCD4icqhNsz37o5eBKD/E/gP5d0xChGigZQWPPidXDjC5DlD
6boGCraqcXISzmIKZYMNkWCL2D5NEdxSJHRPj+vEuG0SY6oxUsJ8RbHHfFZKAAwZ
hmBETeY7qGPP21sgZeADoj+zuARDpa5wdf7BWxoiFKBtMGwsBgazMzn3mm0rQSD2
4y4KNIZeQKteo5RygzfGIKlEjURlEhNasD98tv87rcKuXHxTkJT2OC6zjvxBld2Q
220PSksrOj+XCDdZyy70vg==
`protect END_PROTECTED
