`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3GaVCpcqfqdxGsWSR7YO7U3g+8pb/2HlovN10AwMSVa98cfJgGeioafMJw1Dxi7H
ZLioFR7DhivIZD1DieJWGt5p7PTLqpBiytZoDyjMLMvDcYDqCALAilJL1vNreKmd
+tjDeFxb7zG/mi6Jjng03goOhwsR0xyGRfRfYj8d8vjMDSxC6M8uYynAGS68riEg
mLXiQCnSC7H5EKpXL/2at8EDk/Fy91BpErnMCLtHZoCz+gmOeR/mSRQDvq0aaQlR
H3DQ4/SyJ12FrSapxBD/p5qd1SNfjXglVv6QQOjNf72OZwhkyjjN/YNge/Vo5sEX
G1Cvy6r3TvlhvVFhTikwsQ==
`protect END_PROTECTED
