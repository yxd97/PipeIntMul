`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XUHHA2R+vHA75ZQTIHw6N24y2sD+0iJxsEtITXmxv/eURvnQqD0EjHPTK1yZXZy6
IbyBwJ+UmyHDaM3Ffk+XGMvKYiNYFU6/i9DIovaruKAuc3znHh7DFEj3HfRWdxM2
hmSc/so9MK94jldzqX4KspeR0a6YFgEN0qcu2uQQijqBn6S1HTpuX0N6e7p1Ma5W
8rEpZufcCZ31Ll7VSgcxLyq8SbxQi7FS1j4NX0EVHUeQg8pTt7EWzZxToRGM7aMF
zAUUmSwmSeC7oiHIRavdZEbelJWLMRaNJTin+Z6aEciww3qJN0z3mAFsp4ZDHKEl
/R/LoKW0TcnvxVH657wP8P25S2g1qX7asnJb2RW2ev6dsnRPeg6Yia0206mcJ6LY
`protect END_PROTECTED
