`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DKqWRCOrL4gKp0xX/OnTU/83lCjlNoF2YDnYwI1lPNh1J6tOUlq7nIEb/rGERXQI
oDC6v/z/MZcqaryIHj24G0v03WFN1W0etCYf4vtHlWyjDosRrLbbFvfhEf0OQxC9
09ajxik3Veq7EAhhjw/kW6dP5MeML6C/3PEqYZVxIVZoLFXkoI+Fm29TJWbfaiMV
O/FPxr1Ew9yuYZNjYe5H42ix2Jl625O+e66gsKUh/oHE38fSfBD3DmMlRKeMBnXw
/Ztdy6I1YkSm2xvMP328kgmrP0abdvH7y+DWRKABu0B8naznXfjYHSIQLVR34POd
ul0c8ZuKT4K8/pEfGJOZcjRelnag3+qXRHBs5YyXptdjOreYYhbwLNVvG/NL583A
V8PBKF2hFzml5dlTa2Lv3vPheeTX+DB6Ssd6+/FE5ZN+vwaYH2yBC7g7dX3sOMJ+
QpQ3UBiDYbWvUF5f6JYXCT8xY5KxfDgreUWi6UceAdo+72rmLU/PV6+NRalND8++
QBmud9Ao+oziB/lL66EbiZufa7c+MROAW9I3VIwmiYc=
`protect END_PROTECTED
