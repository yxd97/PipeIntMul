`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
270wtujlSTuOUz3XxSKiQWv4A4qGSQ+Lj3TfZiI+pujwTbL3vM31NnAwzpELQiyB
U+ebHT2rAepvIt7b22d7DiHIvhSMRfP8QTQ5PT/3PLRzzm7xBn35UGeSg+BaGXdT
Fid4I4CZzYOSmMQxZIwZqI4e1VdVOyrX3tBx3ctiH+Go9Ed8cRKj6fvoaWOgyNMI
dwUmjfSY5P7DtvV7HHrO0IC+Dy+nkfkuM3JJXbF1MnC+nWCo/USc1zmZ6nKeA1HO
b8CbRyjog4GeiyopjnOf+N4lfeYvuRL49ZM+25GBZ/jVcI8CUU4AevpQEVGy+sim
`protect END_PROTECTED
