`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
foLTas3mMc+rtQ3CsMz387yXqFN/njox1ObnnIjyCs55x4JqstqiS5gPZ8gw5i2t
dngJms/NBueUsyZoAQ3cb8wFwjqzgidrAZUa/vlUEeGNFVXPj35+A0qrCa+W8hQZ
pVk1jBMlFwHOcB8mrOIlDhoCOPLXoGjXkQkV7i+AF9XKGdyfkcKoREiWXOlK3Bpl
w20Zm+/H0hTxOJR/b9QROmYW2imODyGFhDIETGyD9TG1CFjKsxtb6KvHVVl9dMdC
BxXH3cxDmk7nstCZoVSizZOwtr6fpVbjfZSu+bowRbY14DTtvFZ4vTqC2mk8tDq1
lmZslT+QWQvBpqlbUOnEuQUOmHefjziW6eIhF+KrBjne8y18xEhIYOM7Y3EPFzkI
+BXiOwwx/cXxezHXstC1VbIecEpCdiN7sFgI/C3Nc7QvrGNuPtZwcc7CGWiz7cnG
51rw7u7K6zbu8HcQB01n2LgucAGbOb7gvu/mLH29bBuG1l21o/VJHjUOvV+h/vhG
D1o3zPS/gKr2jqSs/nWmiaq76IV3X8bln8I/K6qCBJKh5QOPOm8K7RF9jzhSmAIu
Z+IYt8XCeNK2K/BTR/LqpZmfuE+ezv3hcDHEgODqRHRjmK9bM0ZZvwVTGxs8zciY
K/AbWBFghnVAleYLSn+lwA==
`protect END_PROTECTED
