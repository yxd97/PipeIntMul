`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b7minp4lYD8BeZxzhN1g5FuUoe+vt5OQ4qoZ8lszJDVWH3prcmNIt/UGsJEnol8r
BxFCUHvsJedkw43AWJw4fVNQckaOgah7MxeJWEWtOcxiA/JsBO+rJQRQ6XUEZc5z
NrMn2gmhJpCuiZkkKQ+/o0x6+PwSTvINVhyTV1xCtCY+2MoslI817PgF+uwwO3QN
JQmeeP9X/59kOHYgfh4jetAWuGSABgYCfuu2zoWOXF4sWqlOn0RBxge7ocu2uvWn
+iUDbddkm3jSya4RUG9bQA==
`protect END_PROTECTED
