`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7PEgy5FR4VDxpnrkIy2plDSRAKSF8sEYNWpHXZQz1beS0HzZQBCk9H0NmOkphcRn
bUpVXncLnEgaN75NCZzz2p0PZSZfNfAsgxPbMaCe/KSw3MUIi7pS1U9E3C+n7ueK
GnPEQ08WLzyLc6Hex51FtPF8yZlOfZPdh1gBLhPyiKXh/zTGq43ktc0NzzO8FzJH
KAQclS/NIqumns0Uu2TayQBCP3TLmA/fTq83Bzw5acWLYcnrqNpXaUV54qRfBh++
rDVrIOcjqGdUzWMJr4sNh68+Pg2Ce8XezSm3IKQS8d7C5ecqNQMvF1C+r7JogCjr
/Pj/UKV+CWQtwWiAHugAQHeeEHC4dgK7ROUYmn7Q3+1qAAJPpZgYT0oUY1FretQ6
sM0ZkAsJ/li6jMKwg1m+GVSVzvyF4IGph64wFy1b57K1Hsvx5ZizpYtpif5NpbSY
X5TL/9urFdaq6DVJoma1v/rjeJJEps12wm3JRPR76YcrpavhkSD07iYUX5btNKzN
kK4RMuf+eew7uZD1enVIO+6qtUtbfLXBDYtxQABI+4+nT37F6qDGSkksoSn41o4T
Sv2OVueLlQsBMbvJR20GfbFL/QI/X24z6iVq0E+igiiRCjibeeNFSdeNKhtjuMKa
ke7h66uTtJJnNVyhqGbPGV2LoF1AnWTfUZgUUnS5d5KxBSepyVS57r5dVhia9Bma
oW5H+zR2RqFneLfh6KWvG6qmuY3dwY5eCCLEv3lFq0/n/G15794k8Im5Q8cPWLXe
`protect END_PROTECTED
