`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EJZhoG/NQTBPX7dn0idPczTvk20+nxrgX48UXfVxHPuPFHJ1qU3Fee2Ls96WC4jg
N9HSJyNEozV6O0g12bGHevn1sgvrjtIMQp4MXdkzdOU5WKyRQPy7U7rOChF5Wtrg
O/m1F/VajjzwZMljCiaG24ySjzbq1XsMDIUjeqj0u6fa63xi7vfkkmRQ2o/51k1h
bmYsojre14PIUazd1UKDjIwxv11gqWhLHlS0E2F0SQ40qtjz2Cr1L/V5I2PvkORb
4FVt++DJY6B+lSvyXvP2njEKV5RSa41Mf0S5p/0Mw346/hXdkbq8KEGEEbfK/94c
nT0vqkjRcVh3bza8eXnlwmT2VNheIn1ykmk0cP1xALjgMAEFJyL0VbVSGi6wEQPO
Pd/3fNG1IHvsCr6yiCZtnuDtHOzhFAPNnNajwyG9834=
`protect END_PROTECTED
