`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7DOtEBJ+0kJwTJCpAq5bCbYLIyIC9qf0lT7aMyUn9xRfZDiqFg5+1aJqTrQPHtUz
0LkDOPXmdnM29yxADAOlu/i/qt5+L23q0XIjGo8weXNHr1IIZAudeIRTEX+y/gF+
GXjMcVL+MI1kv9Zdq05fJSrtLwtji+G1oWS/AnQcijG8kX/yzgBSQSPuqQ9sNjhd
HaEooBmcHO/8QVErMqrvXeN7z/n1aGCJF8/2RmogaIANdrQuuso2YMsyPHvyTysh
Q1WhtBN9B1SmvbkFe30ZeLBrpzQQ93Hx3i0QAEaVDI+cZg9pXFfnXtQOquJvczDI
bmUjxD7nQKwhGsNPeHEJdvBXe67QfC1yor3MGvF6AYfMN4H3Wjj6NnPf4Ph691v2
f8/1pIIdr5vChnA4wOnVBw==
`protect END_PROTECTED
