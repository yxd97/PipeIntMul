`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3XQBQKhc0+UfxO9tuA5iRMg8cs2/TgJRMUqo68t66avtNuI2JeaXSicUaaIMjyY
ZltanhVyA7xDonK9tlYGkmGk69k4ftX474pqmX4fXdlhx7s84OWdndOTveCBtxLt
A3lZoeirubwK0dLH4woGJHoO1ybXd2ah9q1uUqdO+EV8e2cvlX9dR7WLuH2OBem8
ODh7Yvk5fcVXvHi0/2JEM6Jy+nhsy5HhUNn5sABv+2O4z8Hk5tUQ5NiUM6UGU7de
4GpFlIOPYK8I2aphTbGcMUhGUFSRKBbi0sJakTwV0uNHydbJ4D9CJVnQqFqzR3GL
OUQ9I5wT5pPTIQuOIJ7/InaoFsHEFeXO5DCXPIyO6/JEJNTOdqK3Osa4RlymDR5c
8YIZB9SDGDCPQTnVkZzQk7ozQx+5nyYf/rbmIuzR7qjQirXY3ZDBTEWPSY5sDmWk
LTsRF1wDlJD/X3Cuh19o89PXU5JeZPmOofp7hZtBGqc=
`protect END_PROTECTED
