`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7WRBeJikdl9HX3OUG0D8WMeeOrfioqddbFeKA3cv1YaJbWJsY1twfn7qD4cAQdoO
qVPFI/YcQm5jZBZR3Sd4d4L+IUqr+HE2iksvC9XhFUhT6IZjiARqpAATySAIB1vN
gQStLsuoLTPQIO5l2lTrG/e+U8lP6tR+hXv0ZCCfwJC5QO0xsPfnjy53XnFukpbn
hX8GItTQI4jotaZ6ZqnkCxMPhIZKe0ojlSXMxhZnL6BAhF2SEYy+ypLaMbr/3UPP
ViJ+MivFxeYAU1Ap52OFcA5z7RKdbaMDoXAKKuMFyWPbREp4Ib6LYbEYvoxyR7mi
30vRhm8NqjZhoGBHorkKBDW3+aFH2hmIeIDO0U1dPHaoCeQKUFbNQdRezSxPCcwb
uFePxyCNg94HYy4Z/OvH2yN7T3ILxvr7NkIbr46NZPNWDeOZ/IhuMaUVWtCnDHF/
S1wWTQ9qUQN6gdm8OH7qmX8JiyhMefYaxwd5YutGEjqb5djQI4Nte8zQFHZQfF6i
e7kQlT7FRuMbihy06JMSMlEMXOYECw9/8zh+Fk4f7tDlM6daOoloUTOyC+s5fNNm
6wDFa8D0QZm/8aRwVagAMpF2I4mEGsGVh4VFtKce5PzI5El+gx1D7g6aRvqD4Di1
vUjDlRT99rqzrHvYojRrCsy4X2Lsdm+YwaOLCGl3J0AriUYEBqBrHfoDQEdrk/hJ
YvVjHA1J2ka9zBQ+mwb5v+DpKGeG7GdKFm1uuiEYoYFlKETnbwKinPgiQmV2EOY3
pCDD0vKv4uAQJQTLDhIzSg==
`protect END_PROTECTED
