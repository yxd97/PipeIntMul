`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tj+rF5KR5nGEYUk4N+yW/QM8ihjl4Zx17Gle1hxFSn8Rykm6PGLJrSUkr8Cqy725
JTsHkLOlvXPOEeOCUv1CeUbyemu4J4M0uvrE9WXEm/Li7pn4itQktC7eeuy9TdnJ
z4v9/QNSxNAvQxD0lF6VVIbvjiHCK0t0PKPh8Uq6AbwDBcj1ocezPvhVYCRxd7Dp
QWDmHnXm6wz6fw39TMXDDD1jDoSWhj9XeoC+hatsDR1FFRXiSeSbGyJM9bSirVxt
welP1KpAh+fjh4RM+GZfBhNl12YYuh/H1wuvbIYYG0NkFG6ZdkXtWnudjVHYj4+M
a4TsSYYVULyaVav66hT4f+bAlmHhG/BO6dE0MeMJI9u2ihNYFPYht5H4RVoXW2+V
hxT0FQYvz4ert3/TnzHbIhrEgXwWP2pxyyEhaiXjH+JNRiwGOAH+tL64jRpLgNXp
P+nQg0d/goplSfENr5QZtz+dqWgOsUgdXQRr5kl/Ix8VdMg36/dkCZZKcsTIHz6J
dgthhLxDgnTYZgKHV4iOv5knpjyiqKt8+pRbKRPLjSk6bZIqXIm02LbKLIcTHa70
w03P7OYeACdSl3LAwTP5WV4LQ4bRLJE7PafE0IDjKQOELdPQv2fTOAyaEp4SF4Yt
i39j15/IxXkeUMBfNagLWnB9aYDvxKCFpz3nARSFPQSbsbEW931LEKj03aNJk1xN
FjrsvCIPiqVauBPPrE+U/lz438OG9LSXpe9B6kPuZP4OKiI1pB5Pd3mZ8muspy0f
uaBxTncMq62OMJJunCHNYyAAWV0HKvwqyEl6kapOCcrkbQaYDkISnNTFL5jh159X
5XkpcoJrTpv8vGzLfhqrrE1E41MgSGFyPmTEDODXryHWncyT5ed/SabWTtukprGf
n4yza0tTSFYt5sOktQHGfm8ThKblwF2eHd6d2SQrVsWlDW7WEgRqpn1vZqGrYrIE
ft0DuJFBpB6SVWE7kOq/8Zh+zMDxV7yc7F/4Ha3/WiHoFhdNkucxDJWWgL36eq1s
4AMTIFWefXOb/pRvkkD+Pu9HGwKNoOPHILMytUo45ike7Aq9ucdv7QMSXtaPTPmY
IsXV3YQsFr+Mk1eXpSVX5A==
`protect END_PROTECTED
