`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KgB7DINkYvrj1x/tmS2uKo6MM1+C1tDIVTNRmi/9oU1WEbYAFWSRm0mmT2WVLOtT
KTvpW8DIbODsZVa/weyCw+aaQY45RKExUB125UgR0rxezyiWb4pS04H8aJr4/VDz
KvJaKXdt+KTcrJmqP0TyNiQNyR1leMBcRbIQlHT1NrZuXmqN/+L9x27fjvCXOkHs
DXtIJLD9nESnHWyB8AXgTMwi/ja6uzlqRhp2AxcVfDOui777J9+bQrVLmn7SwU0f
EdXMOwmbvTC034wn6hYl9k+m1a6yHjn8KbqaOsLsnjE4M5hXMB74FfpuSmg80ePc
pP9NCbNbGZcbOmTkyI4QK8AnAVYHitS7FT/v89aYOrvVOMT2ylPWFrPsbEeHYX/Y
ebgU0jOyJ8ZZTG80pUqZysIdW47VN9QvXw/2RPIAxt0GvQXHLxblmviFoREBeOCx
EEsL6eMYTLvsrEGZv3OxXtWRo4xRpenjbOq1yC8bO1RZvzIB2dbOwoeq/NSKGRjd
UpzntKn+s+yNhlBzA1n7ldMFmbA0msb7sO/1h8fSwzTQrMLzVesp+j2dkdhx8Kq1
b7+llGGSiwa++o4p4b0dwtvUZjJdTYdrKql8kwQz3GKg+h4cd7eozBX37RmjI+88
54DiaR5yCMpF1bSAR2rRHsT3b51i0FFvWfypTx0qDSdwebV6Z1enGVkUfazBINg4
4e+8mjtzi1cqpfQnOsdbt78LEIY2v23j71EW4JsxXiaGdeK471pWpKxVHHBFiukR
xvrZurWb2utmSEWITVOhwnP8nyptRgY3AlowWVblT2IZZzYtM6/Sr8NKSgZVib/t
muxBZTBrNIGWMGJOSIAXA+/DE24eatERCARm5gpI6JPTv1z1zYCi3lrVLgXFpM4D
9Xe54fzBhLePkk61Qt1Om0VQpu8vqa6ZgS/gEVn1CZYqagVNaHhdALe8nKrMEgG6
TSSlbs9AeuwOlOrp6CR0A/WxRJBM5KJdC07B3U8AZLWbCCipyi91mqmFnSx61Vrc
Sr7YdCGqS5pkyZPV/xW5VNhDpAf9Qi6GwmXRsRr74nIa/pA7auNVNXFm/uG4UMqp
3t7e7+bPJwE62tqmQhKiJjZUlgW9FFXgP1brD6tdzgH1tmBMJ6l8zqm9EXPjhaFN
FMHGRzqVZdLkTVTOBGnvp/K3RbTg6U2hOSertqflonnSLE+VyDnZE6VqsPZsikyp
YVrl5I5wP3A2CgMIoj94BXSm+AzZExtXpk0q7A9qMJLKCDodMUmcmXms9PqeQlcy
FB3KfwA/jAMJl4CLw6Lw4ST6ww9i7UksTZwz3WDvK6L81wd10U8OdLz/GaSNh7pL
1pPvt782BXa3u/IVaCtJPV7RZ3DgMQFIsLK6LyW718/Q3wipPG/FD6PFrEs/NJty
Hfj2dzVMSivxLQNWHmKBcAu1Lao/gZ66stm5GOsZjbf7m37Injb48e6FKDXX5gGm
ylDKqaAEnMPMyagfj/qJILCqaEQUPrvbOem0WYIwgqkSFdOzC4RoYfEbVQz90WfY
FiHtuq40482RmR7NAUB+AsLZXy88W0ZY8HUQ99kqBtHZ3gdC5MTNgqDwWzuSnDpP
3iySa6Q6WDmb/dZZ8U2Q6NBLajJZCvXLGNb4dI6cwmp1d7mTsY2tIRc6z7dDRkoM
KyynMLT/zJ3Tnl03Kmj6JgYVs27KZAA5zCGVMTgHUbgqVVODiUa6wdsReEDK/uoq
98tZBpiLyRa8eRjtnr5t59o+Hifp5s4RpcUR9yS54IWAox3jkr+LYXhSze4Dq9AM
Ea4Hua1G2W2+bWKs8sAbtSznOoGIz7JcIzBhfP7l5jW9It990DHw0AmyykKkluKP
OXPljZsdFesetrz3nGH/L2hvywE4DuzzrFBhBM75o1Pf12MQLc0e6IFscM2TGnGM
LjLpDwDdgtZ4tTGmEyeCO05OcqAHb7UYqRg6OQH2P5LOWp7XqUlq7DZOZfEG1zdQ
dE2yghScnSZMsjZCQJIZefNKjfOyMV/7vphiXtHz3u4mZpxg6ovDq26WdMdkNP8K
+PPiwvsaDltanm30HKRrtYqQamh1ttSD1w9EwDJhJvDzsv9hLemvxopzpTOxtNwJ
xcv/QY9KuArn4UihDvA1L8/TO58tw0iYnzqrMEDC+rSvxPQreXSL7Re0r0qsjitD
SP79/ZfrnU01Hcy/1JIl+sL/tyng3c3JpI4/i9Bmil76IxA+uFpTP0KiIkjDhc2M
SdyQpD9rjF6oNjuFRPZC/7mPftP2wTxjBCMPlL3dz9QNi7rYpKllNExZNirkZKUf
GX8lg3pnixsmE3m7NsOEzEqmoPrS6JFHrHq6h+iTNsWxqu44BSKHiHCrvpRWLHGC
i3SOMnv7prNiVzSp7NWPXRCImW3EycRbbqs2QGGVdsioNSlxHq/zArpjEv/MFIVb
c7wu3AS13F0Y22Ggd+Q181y9HdNlQw00rrUJoZNaIvSbiN7eEvGNk1/Qqlus/Ym4
Zoqw39qgQXRiWBalzSqq3cFVnPM6o5uwBGfvxWuiXsxHAJK8nS7Y/7qQ9GVW0RyK
AbcmZTz3GrtqbMOORsWaBc5W0co3ftiqx1cFzaTPm4cnzFFqyN1sOcHFHRuY/g99
vu5Y9YGukFtJmUhGcQTlDuhfW9qI/QL+eY7kAOxCvF32o3JDmjL27KkDYsqS4qBu
HUvJCCSyfqK3WwAjbyeSNzZboipXUme7voeoU9JZ11NIIlq6qHnkz+Z65b0n0S8W
0EoxiK9ImbLVDCCedn18LODj0sqyUxttePB0nVbfHNeOM+1/Flrh6r/TDErDe4EL
`protect END_PROTECTED
