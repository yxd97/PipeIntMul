`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWTZZ9W0yGgJqBuQx0gxO2YdT2wxed52ItOOKuwLcvY+4LGNowrY0yfpF4JPDjem
eBUuKHz9d0oQylKBcO5UxXCTaNfE5Bwry9XeKLU4CizSVw0hQ9/A4pxTBm2oo/Jz
7kj+QlHrme3yJMH0izHJePXuloxnRAgNJtE0UdocP77GFYcxnfBwgF2FEy5NFK1G
ENVUU9J3bBsurJq/Q4QNETosbBQ74QibfjMsf9hlLFmiwopkk1k/ieKGfROE7SY2
3s7YqTGqQQLOoxIR12FzxJIpBMzZrMIKlFvy5vbHoayxI4UtrMVLbwtTPQ+Qhr8X
orYuqcOqDR6mLimpB273rV+B8LQD0IHy36BCmWv8NzjRiXNEIamW3AEvR3U/Ccef
`protect END_PROTECTED
