`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/qGYvA5h6snMQhw4tA6xCsBJpuxr6K/eq5t+iS00KbwEhHLNe0OgY9e4mXhv86wE
Tu02mSrZMoTDc5EcBkvtUA5qOYKoUapAbihx4Lj7lVVOEwlE3bjcQmXGpdIDEVL6
ZTYG9orV80LeQFbQ6JBqjFNEWnIJLUBJmJDzs5LkAUCtwRbYrRHHEilzBEQJc+BF
plKCgnGw7ac4nAPB573OPVuyXSVGhhaGkR1+LMlWRL56v0Vhs+GDhcCRbgzAzThz
CZTbIqEGDNuj/JKc0H0Lrfp9wQBTu6DsB+93pCChTKQJV/TPW19dan6uYlrOEexh
L4vk0lHNjrZKTQJRRMJ+QEmoFgT4Sk4hDpqkzUB0vUe+EVmQcc110gC0+6f1/u38
pFZMx67wWgILS18vyLEvP4qEoPQu+P31ZKj6T6g/uhXy8Ei6PQeeBSVUCSKN1iuy
XBJ9kopcgUsftTgc5j2MOLbhX+ormL1D8umtyGKPxmxehcyIM0uidTDjgQYGBJUl
7wjpDRlH64D65Q8su8ZqFrshhziitThmeOtrHP2QB9/U66A/Fp7qaNLjjl390kHK
dP0aASZ7aaV1DTTRwHiOcqpNLKcljiGqdlV+DVluUfB5+HveDXejwNZ85IIleHa/
3dJ5W7Ed4gS+f6GLSB2QCA==
`protect END_PROTECTED
