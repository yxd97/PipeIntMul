`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OCqGmaOfZbuQoSH3mPwTy2Yp7Wt9O/gFQ0sf1pKOjl5a5Xzu4sRHheK++GoZDrWF
mzIQj5IcNf0dNBFnXfQ52PCxf+Eb+Re/0ZPhlRKPOMxbp3cCn9YYc6gTLENhDpVl
odAi4m4YT0t0aRuNYXlkpnLf69U8MU4ZrMVyfn9mOuQh/+JH+h3A1/TgMFRM3ME2
eoJK+TuZQaz1yEXvjYRdrnCUhicd5buFbltaf3XaY0NZMxCFNxf8C9RKm+dM1eUR
PodxCkyrZDEE5S2HjA2Zx/B0RKvbT3M3sQSWP9hcnkt6ea5TBD/8a9N0IaL90Pvv
hBzeaTmAvCrSCFltmYInT/tWfFBp4OhPV0HLCKYf/L8IkChFObUUZaw8hVChHjcs
3EmCxMNgH54iz+ZqFPZAodtWwSiLurdVdNCf2z4EgG5iN9CBug2wS2J82DbDBjdA
vxIsTE0oDo4jLMfxz9aNTKNuBwOODl3T5nidaOZBwUaD+ouvXYEYoib6xEheTQlt
/Das3kQcLIPQbjRet4grBPtZB9zdErFcU+s77dVYyQmOhOUeUmzQNanPRAzKb0wI
1sph1QnegUGBh5o8vMoeAGSg7DrboD9Mk3iviSby1rAKbzaHUNQcycZjjkkNCXmF
Pm6CC6kaaX7oXYSEXFb28ySLycu22GieHLuVA/SYi5M=
`protect END_PROTECTED
