`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k345tIg2tStX6ZpyiynrrkEAy50QF7F92huLTGlcy2q6ALclgOjh8mLVoi2iYR0F
hkcKYD0Zng94qkILG1IAoygqi27xYketoy8f0hD2hwFt/8sDln+TfLTM8iJFpwB4
dnQoNoLi1Cn59O1M3RnAWHqP2i1moZ1U31AN9YMYhOC7uSqTiO6G4dtOD5Uh+3fC
Bw6kRvL82wc4uJpAhwLultTfX8/RAyvNc6pOrc+lW/NDBnuQnlHk0+eaqrTgDg00
mj4zJpPfWicrre/BoHO3zW0/2G+zpLKJzvIjfajXW45iPEmuUnT1OMlK/PmRlkrV
`protect END_PROTECTED
