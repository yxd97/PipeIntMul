`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Ziji8BubY5gCzktipVjiskpegm7Q3sotwrMhX/TsHQNvobiRLMY0PO6VOYjLiN7
8JK8V4D/Si69Ga11LYoBQnnFFbGTRpjS55hwDAfg7ZE7baLazctDU3jmBC5BbOhg
2iwfw15PVzBP3c0AskGOyga/0Ua8iQfjaIBDPmuer6GvPwdWDp1+k0sUMfRYEx20
LE4uCqtCDw0BYSPaZaLWFE0eW0M3D0mcP2eMSmnx84wf54xstvYZ2+YmDJfBqMf4
8W2faSV6u2ucoKh2RTmVAZUe/JSnhtDTYts6BO4uAwwusobaJpda+Va0BNAcgIo4
BmviL5ahF0oDlIrAzSdd00uGEaAIN619xpvMSk1rctNA+h0FIPtraK1F0XM3XDOm
utQyEuj5XopYgY2Nx1D55VNjUaVpoE2D0Ic3prEZHJ/RXoG5leQ/cbxAlVt1t7BA
NRtSOkUgjYVE5u7yyADEOGnn43w73wHXicNeCz/zoCnCneYywhEngyGYxVdmt2/u
9CYPyM+mAQokMaxoVW3wecgIFTbVhK6xKN0PLrtgXJfzCjbb9JUWZ/nvZNXgLg1A
+rzflOg1sH7QT9pGvEZ1XJPK869HPPtWVfiql7PzxOztNbKX0pmKNL0ZzsVHi9ip
H/slg3VZ+PVMcY7Ost57a4bzuIg9RNrHGMPcKsd04Xo=
`protect END_PROTECTED
