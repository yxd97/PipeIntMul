`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VKodBY/fyo8kvb0Ox+NwGwSBoCZH5UZpe1M5gCkBqM+UQQ5o6gRtPSANTdE1ULa0
fi9JbYsnWnYa+T3nAm1+bAr7wNqZV9Yhu8ekLCVNWxMtBHRBghM9/wWHIN78wt4a
rVFg3cNdfKUM1MJzUjR/bTwiOMsTjQumJszuUbALGBWoeONs90Cfm7boAYHbyc0J
7LWtQlkVi/7O9KzrEWdxNhNNwxkFjU6LPWtyaHFHqa7NWv+A0mhobTjoHU1NSZKF
BxyWAS/nFjWwnsBP2PeD2gLQIsXeIFLpE5OvIZCs1N4RPzj9v9fZf/O9oksd9vb6
+QqcEMV4Yae9Rr9IyscnwshrXjAsiMBrerILV/dm0DLLctdEpKonZ1zPW3mD6+an
kf78HDE789dwS5ADFgJ3oz/BU+yP6MtVq4roK9IF2uSu/dO0ZSzCV5uqaAJePilQ
nkDB3firy+8q9G8alpbvcjmC+YJCdqoAAZnUCqI01ArJSuWxw5bAH4zV+OXtFh3N
ZqtLIX6n3y4jG6R5D1wNvCt8XJwGm/nC4piIeRAvW9NaKz+DYSgaNw1vfYvOQxWz
LdecpBVU9EFPoQWMaCvQsfujAw+ydDJhxQui9o1askEHDldIJMLPpaNP+6+pBo0Y
`protect END_PROTECTED
