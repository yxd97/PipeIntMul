`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7tTCHvTpNr8/Pol0zLSMclV2J3BltWYswA51k1D0j3QZY5HHddvqcCuqGSyK2iW0
49jU+Wss/WASW/aH7bgTDMynz2gGUfqGybdVPDC+1niVrFxtd5GcprF32Ia65NtK
d+kR9cfxB+kCSrb9piQrmL3iO2zzcOMAhnSky3SU00G0xi/bER0hvvHrRguSl/uY
RzaK6eDfvAozlv3zCkCuY4fQMicReYgpbzUAVy8XkWJ+u3+2ATCBat/UHrVZ1qD0
CCGLZOvpom07U0X8BMESqJQc4plrXcBS2Zl1FHW8Or4fgvfxY0gIIv5xpi4CLwFA
LtjEVzfJlMi7psP2+DjMZFUAhuB98A7rLJ2LfeK3xzxSjIF7fiRfxTaZNqcZKAYb
0PqaCd7txci9YUgECqEcQ4P35XjWrzqX3aH21HjsmHh6v4Y4cXn941xUi7uhQfUR
TvdV4OIfwnK+vqavhBPB9X3ihHztKhz+jvGICxZA4ZXDREj9ZiNjc4hUvQ4aHCDv
+2UD1wvv6/JS/sXwXLI4fb0P7nVB6kM8j5vadyxPJkvDnO3yRsWq7lt4d+KdZn2V
ta5X0QJaulWg6FHdQiFCfkf0XduOKrjUF3N4bqXD42WAhdLY8shOvMQFQC82XRVQ
9Me4ZxuJknBMJ0VM2boCSqv2hZTONmIxwGxe75PqfyNKKnB15naHt29QGVaccRBo
BgpnQ2ep7kczSYsom/JCqCgNmLSO78wzHwbjvGlddmo=
`protect END_PROTECTED
