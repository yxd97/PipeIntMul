`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CH445slU3DOYmKhWrPBmN187/OuQ7f4JiGRf6Vd1kjmeYvAxAb7m/SdPW2guk/l9
sIqNw+wQL9UCsIg/KGeAF/miq5Slc8nXH3u/Pd8EnQHC+clcXEXDiB5in0gY35AU
ijugifmRxzuuC8sQ4mjk0Y5blaXcRpJl0U/eO8k40K0EqY9bIdDsXGpSiarspACI
vZ3yFhuG9Nh0E1sgTMJYOlW07NGQowyp9cUUhmAGPfGg1TOGiGTU1HzvE3iMgtH5
4Gk9LLYAv3fz0YQOOZxTqFbzS8pQ+v1cKKEEwQjmj5WIa7mk6bSaM5Vb81wGeFe/
8UXA/VY7oMwFFNPcQEe5Nb/M5ZOZma6GBcBvSADYJ65Yffs2ymhwDLyL8IQAZcAU
Jo/LJrw/gwHbZgT+/auStZoD0Km3do1kUydSSONYsFjr0gVCHZ5GY3+C1+XUCOVh
EQDTBXAorf6+V+5RN8p3J4HMHmFN/wcxXVI2HExKmHqv4eJrP7nc3WX/z3SWjqLF
jx9x5YxpZyWNEJ6bmbuRJXZtk+KJRU1vJXem503YTgme8HucoIAKrYkuMtuEtwNl
Lb2E5uiS5jcHJsj7BGXJYkzUGgf7qKY16fQIP+0nUP29+5ufVsztravyu2k3HG3/
alIKl/wzPbCjfmjaSkoJi+ySavWc6sCFgjcEln6FfjFtUxkyLLqx0MML5IZruiWr
p7xmuKIs9wr5ZNUsGL/zdYUurU2j15hVWkcrM8e7Uj9XvijL0i0aZF7QvLbx+D24
sNLQK+R6MWRkCA1J2bwMpAvhEzvZlI1btr+rPmTXbdKJ0TX7/2su8/DF3Sdxlv2s
0Gdy2gSCiX5abecXgwKpH9+OZq8ngIOWNazJJuf4am/PJ+SrlUlppakVu/wGDyV6
dKHVeA07/pS4GW/1TSX5TFbjTT452g8VIkZwcU+9mrilgM7qsFxFJnS8yPIbZGxy
pb0Ktc+K4VP/oQALMiA6iqUZ3BFjFA+g3/lzSUUFF59+6naeUtCwXS86EMiaewtQ
XgIOh/OuKam02/aj3OaI69NeQs2qKfQVjX5oQ407Ey4wlU/ukv0et031RzgKQbSU
AfQv4BgY3Vh3X52CmYzPUQTVcZp+aNSGMoX2pg4qdTLYAJRU6RVr8puIHNk8N3ei
UBjbzBabPICiYeIZwQ6i7EoeeFrMeACjfnO49vWWAqew1KIckYrOw9/8+aKs9DxW
X7i/AeNrjseoL/4obYDf7pblzYKRwqt3pSH8Oc12blh6XdnmtsCuvoVnUK2G83WT
3S6ipczNSnn0zxwRkK4p8hXBoejwIpoRhbzPAjl8yOQiRJ3CiIQ5mbSEcnUREkoT
knjNrspzxs86hWDhHxHdwQMXVnvi9qErvu/mvYSyYeFIz/bKn3UrXBmu62AQhOHS
mtSHVHNHxZTa+Oa/lsPJeTWygaLoKp+1A6dbPG24A+AX/+YNEmsU+tvDNn5bqpLb
C0XSDxG6BjdEzFMqagr5CZGBz/QzapdbYK2WNV1Q/hbRKluV/rjC5Eq7hwnpXr3a
+n6F8VtLtSGmv5Do0HvrrOEYYjim/JgETPTtpntZvu7sWLVDoYCKSN/XfqWXfovh
lJj6A1be26eKBM/wGIBGSQ/YRP2HtXeJ2npfvMR1+Gxb2OmK49P5toF230s4TLcC
zUf2cnI1aMFta3gwNY6NNrvHf6P7DE8FABWNYMQmElmT2wm3EXt2dtrXigtLQIhG
0igtrVO+RVyHPLsMBYecdl0P+lxsKF7l4eq/QlpG0sxXdK5nvOgW1hepL7EiXEwU
lVkDvoeSWwt7mZoeJkMI/VtOesW07BSIOObwvq+PkS51KyhunLlsjDUXzSKqWzPw
88fu5XxJJFKNZWrXuRPLe4IPIWBSFZhuIej/n5ycBe+wZ4nwRH/QaLIxbqSq8WwH
BHeYB3mI7Xk3cJP1gnva7wBCK2o71yISSbHaH7J938UPYE4KZ8h/87APGtbsaUt2
AcZ6F3Rdg2zZ/qKYscE4uNLeXGl7XIMhqYbznNU4oJ/pySIYMei8bzHBZJSEwVh4
8mscOFkJSd47ZAgGF9WpUrm1UzTKAzLQp6rBDivfpiHpYvaxLpTz7+bC+x+4mTi1
kWNnqGmtWFdTXfkNAzlnRiOrNyy+czmMOMo0c91pPeowLPjSaBEpQqN2Jrm6+TUD
H1IqC5oo8AuUXP60kJuD12fTC+oGbVCedrKanZ7oSplkptU9FVB5svn6eQzH6tBu
QWJAyc/x+MCAiWGM9mKv8v6hKq5l0N6p5Cv+TrEz+OW0NBN5J5xzp3PygsrKB842
YvdCFskxmRlcARi66MZVIsVyIo4h8P+9LeTQM07Un7o=
`protect END_PROTECTED
