`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
98pckE5cpLPY107un9Iy+hCJ0clOqb1xna33R0NZdiqQBHtJEHw8iMvBrEeaNvqs
mlTbCyajDeqyOzh15ptWUBX30885+FTg2DSp/o1wMnavpfRUatD66RIMiDR/bQq2
SgZPvmwWF7Xk3ePEVqWknD5vLP9LVlbx7L1MKjf9hD2cCTnNuagDCChYy6edf/mm
CDj4bP8BtnS/5Scbm9k27E9RX4B7E7OaEZ37CYapmeWHdoYGtZkHgkM/dK2IzUVF
ZXt6XmcqPreW0UMEjVCLpPJxi02cqSr4vs99su3gZnZ9kNene3vEvCj79ByifbgO
sLcHnkOnHinRYP0zOgmIm6OG1K7a/pm+Sjtwdm4knFKYQZ9vVQhzGBtF4Td9QGWb
84T+C0bKRQBPp/EqDI2AyTcdyq+YxAr7Wo0QGyhuKeun2+QXNjnohI1DMeRplESP
ttrxfEIbWM8GsBLwII0J/ySpRzNWZDFWkzBMrCoEqGKtnC8WtAduABlnxMhJkIu6
`protect END_PROTECTED
