`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Z5i+/EHiJwUG6zLT9IKtZ24kBbOrujIYiQ9wEnWXhIUKE3CXuEsEGhfkyDYuGpd
d/IhwVwHqdkwSKfW7jocpEL+iGMrWIyGt6IDTTcT5jDfXdzugPqaG+3NNFUuzOcP
eMNSQImGff+igvRUanrXY0E/gpBrQU0ibA2azhgCKPwPg1iYUMPYIWbDLsy+1049
o4s+KAY/mu83DWmTQCA+2EjOH1MH0HZ0dutfUeLT8V/cPGbUQQfI13VLmPUPIlPH
/4JiU77pv7163/A5721zblZu2mmrej16tXyrZiVK1kM=
`protect END_PROTECTED
