`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/cKaz4ESYY8dn9zcvP92Lq/UJ7NEwRGhYeuXMZ+5zmnNEle66sTdtj0a4Myd3Hq
vF1uuEEMnXIi1NnBxG85VDZI9mlBZUrx9WUkdxuYSLRxGa0js/IkR16/DdYTxXFy
P4bfYuB7C1xa7iRKjceXE998A8VGXRBC2VRy6YiGFfvegNt8L84tI6govx5aLA4P
8tFildalFXGtTrR9HbJw4nWC2pti+wHl2VYakILUyRyNAiJbXKa3ucf+4cS+cQ/h
g8X3SROirHRAw6EMkkkJ0mofpfgM6psRHBxRrWLs6ON3DIKFH2ieNwDAIRB62Ho3
0IaSJ2k2UhqUjQChnSQKf6aVxrtoXK9gLMX2QbEqjX7DpyOruz43wLV09RD0N74U
VMT8v5f9t19f9HFS9w6m61ZsYApG2yGQRIVcOtb9HWi591zxLoH2gElHB6MNWS1q
QFlRFTnlE6FfGDuUBwrLEETnVFYFRGxJj4cVvDc/qZQxjz3xvcGvdcVI1pHsIKZw
3WmQNyG6W2McSvHTYHod0Hb+zGxEMU6ca51ySwqI3HfOOC/u0EQ6rm20Cs4W+5xt
`protect END_PROTECTED
