`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NIE6fTvxsYQnjd9TV99TFH84cfH84MOxRFUyoAVufTLwXiKJJlM6sGLYqQlkbH/v
GW0bCGNf0ZrxDTLthozA0GK69kDSsJPpcr6WMJNEA+CqdherRq/S3LLoKSkEm2oX
U8iNm8wgD5WhbV046x1AduqkW6J202RBlxd5R5+JGhpb9IIQWtNPN37hZCfXE/em
PCqy+3tYrF/rPlG5aPyvII++Ykqhon8TyV5I4GoiVLKMFI1iaZQJUSGfszxY/LHP
mX4Lzhi8qCWi/jnzpqd0BshqE6XlNhGeEQIiQYYUbjSI1o/HlVRgsChflWafSZ3z
xgFgqlkgmF9f8wOpkH7v8I1m5w38mG+xVsgjInwvC88YjYmKy425TiUf421vN59/
8Nllqb9zzgj/H7mkd0O9tk8vac/auDQQJ/h7E3CnMPqMbrDQlEyqXxwZYka3fZad
7COvXdtno+xugkrnRx7DVu2g0+oga6xDz9DdX8+wcox0uXX2rEPo/oQtUjjLwxJ/
DVkUFzP7OLmk5074128++w/+11d7SKJ+eOpJXeOs9RV0B7ogFWzXuTLLfW8UXdxk
18ZmxhuFS7Qc22NaUekPNVgZKcSovd0CrIrxbmDnJyfPY/kfOOO0earYzgiPG7Wq
JTcPjR8iCZWQ3FCHuOYKqUiOU4XOU8zs1dEXL3OnCYDiLp3DBtOAY5PZDWvUReO1
YnL6Gz3q6v1CUi25ppmIzFeZfqcDHsEeH+3RSFTHj4usIlg1TDYV/uN/dkeMBtWi
Kp0/uJJNk8v8iMgWDtK49evC6OkPnij8iTwT4mzvA/gqYFiVIPUpLDG7d+UNrxC4
BFEeAUcMrPcV0Cpzj9J0kQ==
`protect END_PROTECTED
