`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEPWAzJ9QId2ipCLkAXQT1vbh/nJ4BXKFNcEKWORD4Gr6l7elnymhy95MGNPrn5D
3o4yulcIbsSDMVY9KQj6wQh8ef4z4UlxRcXIEyWn2rkwhvPUNwynrHmA44FAr7ve
QQMzIZprygZic3U/78pzkYuCMUcZIA5WrFM51avKod5Rh1m5B3nzQ5XGO3TT/KvG
uBrzPH5e+4o3VvCw0sv+91z/jl5tfvUceIOJiPRCYvxKAa32iznm6IYKiiUsrqL5
vAhn90FblamCDPMgn5TD8ncOYE4eAFHtEhEQoV9/Bnfm27jx4LxP4/pDxFjpNgo8
VRvXf4wwLZ/nUe//VzAQ5bYvk2/xsSKr/1PhQGkYYg7nOYKbN9wD1kKXbWDS+g5r
LNJPLQDnzLVrex4TnYps+ROP4Bqs3QrUSkqE9WgGETk7IZDuQZm/db7QwIhnB+fe
rfk/eBqmPUAI6NlNcNGv6vbccddmREnPcj3c2smghy9RIuEohwcoKYH+Ff7j6DcG
l++vuKe8VAcLG3UvnrNlXKwIH1WqHP9HIKwgbhNx0Y14YjCZcl9VbJSzsQ7PEmqw
QQVd8bAeW0RG7bd49VvowT6M3YhoHrnE6ZMVOv5buXklVKv+zq2Ipdfoj7EpYnvu
iBtURpuH/dbAj6Po21aGAkIhzblmfF2jGKqfTuFMo9jP6/MEZw0P6ZWVJvvFe5QK
z79Ls361pnn7YK2pjs3RqexmmUdcXP9zOSNNGakWbS+Z+jzEPoxF8z7uFkVdj5Ex
VTMe6Xkm4tdtfUAyppYpMw==
`protect END_PROTECTED
