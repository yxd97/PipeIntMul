`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wCHV7cgxZwyzykCXZiezgf7703Rgs1+w4ltsEKsmeAYaE9WFRGs3347OORAsNLFS
VgR1fhOan7InRqCsVgbdnWPrj6UNJp44X42ZStjPJgzIDy1FlpNetoHXN3dztn4/
2q4Usi3+rMbyq4io5CboZyot2BUPB2K+zJFuI5svp1XLtzP9v8QaQvwnx3pPO6dK
OSA2Zu5qNo4vAyAmyPjH2qq+2WqDUNnJFQPDQFcuUYHK4aApVKn9pGIlOZuwGFTm
HwxViYz49ubfcwSWG9gvmN8nwViVunHI02eTd2eBQABSjNTJb9XbQCbid7PPtE7m
VRa5NSCibR/FShZNgL6cWg5+VjpQsDT/T6SWDIxv8TxapD5PgyFZTnICeOP2+vhK
fOH3wUbQ9u/80HDWlYDV+9SnGZlEBqeTTW4EqHLWfqUArgbaixurDYDNMopf2E/7
`protect END_PROTECTED
