`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xv2aw65NSX+pe8xC17oMWm1t8TIwJuWKU7thrKS5wTIBOW03uPehcMnOwworVMx0
qji5xg7FJ8OYOQUo5Yhc5cy4Ec7WQPhXPl++jZS17WXpH9N7xy274b/0U9JSKIca
UNohG48vWqI+niUQ5WfhM6eDErEIZzpaF+bZwaz5Jw4/LV8NF0uuEuuuRghC+QdT
LA42JzYaoDnQ/hfzeeNPYhSxbLxWixzauOEOnKA/Aedezy87s8TElvifWF6ve05Z
UmprDLlFGVsNSn+QYkAlB24BvqMRvvLndozHDrtDmeBklegTZLhEU4KhIRX68OdM
wT5HALjAAUwuP1+o++eE6j61+YdtjIVGyXLEOu+sq9CiOK/K2p8QPkhikrtGMKmS
FTmSYzRgpF4JAGbHznmhjCFqOGG/nhYxJ8gkVc0EnapJ0b5AgjvzGimbf7OCN4KO
n1AgEKIyYYYqKLoNwgtMMJdHhEpVksCOLbjb/MsVWSvDEbyCkgZQnGZlFbtfiV0i
JnoHabRZIiJxUpcXm2Xa2aF9Q8NP9IYrsReWHzAFuUPicqTy3QTH9Of0U+/ynK+t
PhVM8szitHJ2FbflKJn6p/An0t2r0eE9KUrj77iLV9uyOyjSt0N+aheTzXQHk48V
PMsxw9nJCtfBMwJHrOmMzv4koImAIdDHgE7koo4IVERnCsfm3FAKNMZeP6/nLSHH
pCjTYRkcbU1v0+YnO85jNP8s+k0U+OBmqy6X1biyxJ5j9pKjMBxAPZ7MecFFMc7t
FE34I6idZA4HEEnAPfNUD0T29XXMXXAqaSxtVXZodIY6J6kUOLhrax68E234xjCK
p1PiTKB1TbXA5v7WTO71BXuYIBwYVE3xUHeKgdCVEG839igtKN9Cm2KUYCZZI4kV
gIjsD9k2GvqtAeWqN2zTPMyc0Wp3hs0smBci0fLSIc5WJVZeDQT856uGzPBkKUet
nmZz4EcXZC0Y0SlV+l4k6Om/WKk1qzUFs/LniOUwGTPU2wVClQuTTffXOh9/99Br
vL6yv8f0Nt2Xcs5QJRjo7ofXLqlEeHpJv8dh43Ve88nJcYWRTWfd219qabnR0SNI
7DA0H4whRQCbMpm9/lwSQ2bsqgYwr3Ewogii3lPORIiON6TWjdIK8RNns33aArzm
eOkj8cxSrjNKuZf0X1wC0LzL+7lgHPxoepavkbUE4jlLryeIbCc8lYtR3Al2H5iK
DZj1FpsuLOiyW6dsXvaEBboWikpnX1EAmqMA7UR0ZliJqH7fni6AFrPuXegaVxFV
7dmOh8/CUN8WWDrP8NT/3W1mVOEE/AEuxFNM5jEWaitgZ/C1cUyJ2FxEPcLl53tM
mAmyXX4LcR7T5FJRchMfmr/ovfuJOurvzEBpLLAH1UZyJPuC4q3fxHquIZMIgE4R
YJ8bBOQ7uE2h3FsmWkk+2r2+RKgKXvMKtirp8owkBk2/DQoJdZ0vxNQkPm68bQJD
cMjb4WZKux7SyEng7HyPvOjj3p1wGLE/vv5ghItp9yAy1GyJTfvVfST8miagNRfU
n1zM1EAJYXJujxskCIWwuYe8LTAcoixobuaNH+TApiNDeVaQxdMpiM+8GA/tAF7p
Pzt8BRYD+3Gcx+x2RbF3R80Y3IpIw5m4ZzjnWd3E1lt+4pkuG8v3pxMx4gjgT21l
RoBFfRAM9nR6n0QnUZPjkzkGxs21yPuvRWCvAIxYuVgwhJvD8+4qOYuYsIFGpI3U
3a74+1VSca8NV4m/UoAO851ybrg/nd/ibB1ZHvM0qDX+y1FyRMqiI4TUgbxmB1uL
Y7gJ1UR8pq9f7D6RN5ILro+A0yZQN8GD3OGkbkUcjroH95Du0yHOxABkzDHIgllP
d3ce3N+/7f2olRj/VbU+esLEjAwOLTWaRs2N9UN5rqZu7rIs8GS2p6gb4DfQ6Ok5
Oh0qpjn6yrzE2BDWLlmDYcIggBkAeeFpkw7me4OrBeegQS5dziX0DpukiAs0/XNj
5hIHd7XN7vn+bW4swRImoneCrvyND5ie/H3RXtyNBSu55+hFuaa0fw0WX1RUFKW8
RA8ptg+eiYFLGTcPrNdjxGsPblKmYTj4Al1vlA20V7ZKw/mPy1einEFJpHkSaZj2
9qnWw9aWJhnbkUWsm7uFrgzaWIZ7V8ZvG9T9Tlq2BcxqIaQsyY1tKOUm94xCy8vf
NFfnKWEy4ssT4Jp8NDutZ0FkZ04qVo6OKkCqCI3jCxPq3Lp14hB4D+dzCLgBvpsH
erQS4AnvbX6KcG0D67lhkG1ZtREmafiSji8EQqwapXV5UKmfxld9n2fmMIcEk46N
/9lcyJ+Bv1bkA8VN2SR9ifdq5PXZs+IpAUUGOe8CUX7QRp87RvpB5NTibH+oP3Yd
eI2fPIvHXk+LDckITWMRM1yif4z2dMdRJ/3yTQfWt4K/q8hbDoc3h1CQ2+K1W0FU
DavRUDrSmEsj9myjDqy+F9py0/nwmqIKakNzy0xrIvXQ9rfcVsTBS/OIT87t2STX
vM3Ad1fLuO96ZCTIG3HH/1qWB8cTpjai55AIyTkppBHnBfHDCkA1bPW6/JU4oTuD
qHquJcZqk5xSKj4oub39+02lcTKy4vTzfiG1CCR0dcX0XW9Eo+EyADBC8Ag8npOK
P73yJ6suf8QUtIPd5OYIeFHpzwEqO8nOG2Eu4be0Pa0Nr/GpPwulWSVwKCFLX2U7
9uNm8hexVCa8qEm5FzHUQlillCAuh4duN/IPnNBJOyBxpc/qtjbD7U+c0QAITVvt
kp/JOlRB0nfjV0PA7tD07c+CSKl/feN0wL5P4R0hUnLYagPy2tZdyIkyjwns8Bad
EPZ09v+ul0n/VlyuMASVBxLJBzoE9Br7KgnJSerGA4baGB2wuLFlWuZglapS48PS
N/WVed9J0I9EQ1lltSsBvC4QgdNOyNtwAwGj1qesNnXuE/OsudbuA2VUDcRSyOW9
ueGODD2AFwBZguCCNI2MzHckFVSeh+DBqI8of18xD49NOtGKjsDuhr3pUgFawOlb
ohfF5vW65yrgEjjv7mhbyF1vEa0tsnJowSIjqn++c3yUcCsILrn4UxJlT123cRAA
U6jqQR3DXrcB5FFV6XEbdinIcM4knfc7YLiVzXHNw2LG0q+wNl1uBbFIW7xtuZHg
RJXChszqpwvPyGsXVpnNBF86/eWgSEs/BRsxYZ/49N83hIRM/J88CY/t9/ZOPjKi
X6RoHC0MbByAZOytq5IYHoRZ4pUjMuiZpHTLPo0EqCUL/09Z6n4RSZa7HyxHh+Da
x9B9Wtgt7YMutL8klW9EjuDIL9OJycZa9w7iSNI7xJq/nDUirOII5wXSqw34jybG
xu/rot1g0iRHNv9FPS+qTjjkjpinaIg73TXRqquJtnUHMCnC07wEc8RcoUdv6SiY
ajJuTU3P86b+RyVpyavueWYiELTTlZiBu5Mg87SHw6uq0Ory3BthPbZuvEZTCkAm
CNqcwQbQt3o0T2ITCRTbkkggi0D1FUOW2+cfFdpaDD9LsZTZx3NHIFbVNbqRQx5n
RCGZmVWGXC+zNQmq9eEhS1KS8Em1BjuSYbGdyUDoFJbPbfD2G6iJageBfeq2wne5
scfnXftQtu1KeVkX8vysBsKowEtaL1vhpzz58dAnQIM4RrBTBXgtwpeZKHJ8wcL3
BiCBlNOjpH9RrZn5WBhLX7iO3wy4qHxA1Ddn92+DFWEZ2AaVBiSiWhYWDT2oe62S
iYgG17G33vbRSH4+LOTYoxlf8JeZL7/D4nM5pdepr02xcC5uTwHH+qhzphXPDK+C
qUQc+hQviPatAviX0R5ZdPLz3Psv4mtHTVUlHN9mTDfFqoJ+0rsG+YeVO0Li6Cwy
s9uIJACif43igo4VcrgY6YpH/j3BLUJHuaCHwEX5vYFEByyw1ok7j37fvY2Y5vaC
vtS8rhp1vQ4/YAgocrfk+yYwvormtDo3rNJ9QXC7BDQba9fQysi9ZPx4C0XFqag6
S5GRdcOjwXgB3ecGx8BlIHL0TiqbZH8TFgM5Yub2txQX653BWFPWn1NAgAHur3YP
yrzNM5gd6DGLIAdI+7Tp4E5yGg/aGa81LYJYVx7ekjVgA6wg0Hua8qvxiPyV+Qdq
neWcGvuUnBOn6Z+JMtwZf6LrrV6U96PmZYP15Qy4/96ui5PWLNTHHBzITJru5MOu
a3r8IJScNN8soEKr8FbwJbqMtUGV9JIbz23DaXepd+X3lZFqYqL3XpCjsjKp+AUV
ilSRpV8SoDdlECplMP7JCee/AvZ8S1Xo8lgYrtw136o0mqZHquvNMYYAafY8MTgI
fnif2rmyRWxymrC0bPZdMahNdk3nd6cs8mOCJ5v0HyO7BTTmu4qk1VfuWwwzNFu/
YpyAKO9NtEpO8Gdk4K+u13IJyZLpI3iJtzbZWFoHoAXQlfBn2BobWCCgPxw1cQlk
RMAb/NkPufBl5f08GcBbyHVTDR9g9mfv7vE9P1O3e07nx1z2/cN0xAEnlbVrADYN
G0Gex64ZDyxeH4JqQyUeFGKfEyufpxOHEcqOBYh5qXQ1bBN76Tx+S4OGuX1w28yH
CMyJ/sqwL3bgDsDxWrOXWYcQoGIWOUoS3cXVDstqQN8gUU8ktPaz46g1HPFAX2kc
8VY7Z8IJ1KocvwIxaiZsCn48DxS5C+cPvGoeU5fW2Fg8r3XCXTSWKsOttCY7XwL7
YZB/fQh4+CEBjg222C6WK7BfnRR55P1Wb0G9PiXba/RL5aLvPtHoOjqXTtf807Nx
5mwncP88uMrKU8YjZmdHxCu3vPNOwm6DeRIJpyvInhR/n9gnus+cE+1Hsxt9ofT/
xirA+mLZlWXCaYr3PVVsLOVcyrSkjY2wwgfZ3cIF0vVrPHVlnzSAxYoKxkN6CfFc
CV6b+oCh6KGLm4wECCIvyFjGbWBZsfe+8C9RrmbIQslZe0H9WqkKpEC7jW/RFua6
i8jJEf1I+LjKNzV5cuZPYlbnF+bmpBfsWOaecb3634ueAAaMr/uDuVaJ9qsK+Kdc
GQIK+CrlK3K08sYRZrHY7rlLd2wRCxUFO0coDurdP5dF2EAIKgEnZLI9OU/98Emj
n9rTaJUSxlcsEMnSCz44NWW/aiTtdDHndPrdcGjWfs55pGEEUmu8BObEM1o7EpcJ
JvDIHbdraeH0itxzwhFpnHd3t4/F5TOLKUrOD/+hD5R3Dq4Hi5Hpi2fBF05Q5m45
WWISIb/7tDjJFmcHXutLTQW9JOlXqVtbtCMkGnkRcE1CJZd0EGMBxIEtsa7Ay+B7
2jKYTilmR46B0FIKpElNaDY4Cp+ytnhI/V+6cg7ep1RpvjuLPZlZ+u6SCUEILQHo
PRNyZLEiYgInyQvzqnYvaIzJP3KBfkc5n/z1oDT3vWl8FEKy0Dz5SgZwWOoVKJ5q
S86FqvVG1whHWJfegMZIzANJPba9BaUxzieaIHEo/ak5bxuzTQcf5y7o/QXiLTw+
57WC4Rt7JbxjrYca4eOy25R5TR0v3TtwPWpXLt27lE0j2uUpfays/K2ORo2kctov
Y8nuIbd4M2ET73gIceqOaqFb10Ey4S3HgsBHGMNNMupnrbAr4mEGMWROfQ5RIvwW
njwloD/U4XncMYnNchKk/hMIeWbPAhQhJaAcLG4sBnohl9aeDRDvp038THfKfwrt
Akw7HkJ6wWNKz8ueGiXzNHo1mcYP2aN41TwC5qRD0LFJRT9G1iR5EiwJLRfwqVEt
cVCY7DJUh4jk/m0Phywzj8LtQ4N7MFaAMaH28z3pqVBw4gEX/di63hlHDUPfyZSl
N49ibDVuO8LIW7YsXMDxI9u4BEoDr8dBSEkfNG4AUS3BLrLBUfuNFwUUGzRW9KDv
TmseBf6P5WVW3IeaezsbcBkXbVQ0GqXaR4UapMAMV3uDWku2TukbVq9ZL8OS+Ig/
RUqy8BnF798axdtIuKwkodc7X0mP7vpA6WQXF5TJfK87Cl6l8K4+Egtp6SKmRQJv
COAvjqMYpeaAlgDtqkJ36yKVw+dRJmEQlWQ6tE6GWsp5wZ3Z2Gm5IhM/VKTujHqi
1YA73r9RxYibSSl5VMCMBQ==
`protect END_PROTECTED
