`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHcB8SVxKMwUAeBveSThuT7CNloqzrvYwE7qnpmekfj12FNiCAS2l2UuEURtMf7q
EWS7E+ZSlgI9mpS95TcmeVEsF/1/WsFHJt9Hg7hJLEXAQ19ljeoQEzE24sw90pUR
jzxGJSII+k2+U/G0j65l31E4eia1gUD4zce8ztzPEgJ1PE3wN4CXhw6QCWhOk1Gj
dGnkdnZ4o7X0wVl0Kam4vppn2dMjT8eVpfckw1AGeubc8l1ENrkGAspgVnb5MSlm
MY9yjc5uAE5EoVNk/b4xBLMq6Zt5wRoQk66ZAUPABFdS3eB00gExEy6zHQgma2ES
dzgq/ytGopyM6ER/51teHu7UvQqm14ufGLX4T4mLonNCRS3Ndvaau/KT5OnEkID1
iZVBkXdMbYD8cDlya3/uko1ZxSvOQKcSy5FJsOw4WpExsVEK6UMaQ2JZmOr8f5mf
`protect END_PROTECTED
