`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cozbR74xLOkTiS0CcL3qfPMs86tV4Q/INkP+UMY6tVydq+cm2GEeX+DC1Jouawdj
voEqQ/oHi4VThBBKZ9QX4T2TGEpN8P5k/J0r/wL5cTXkWs27taSquOgkKT8MN9s+
sIUbsAG7ieshmtKRMs5D79/VyQR/trQhFqy16rH9t+E/CmfafOpEHjB1hu+wGNzq
OxsW0+9BlQ6PsWuW/mW2Kjav1RPOPxS+iyLIF9Vmy1CqrBJc9uE2+VL1ilYfHGRi
DT+BFAEZrPN4D4sm/oebFTW6p+c/VuXxznZvZqv3p75JvvoaL5C201QEx2YoX11l
LI/9LAgq7fvXoe5DNLoxNziP8M7U59LVZ8g/8wm8emRvzEBmg39VKnWNqrkM2ncp
OtAzo2Q5BhZCcp1HsHvuNAp0sv+Lee9k8zlvYCZ3hIAp3ciIFf9j9SxCSwLtDyuY
g2FddmGIasnhb4OUMYoH4f58yJej71EXgORPjt4yTZBeKMLZLH/WMs5q3l0mleGN
ea7d/+nmpSDE5EyveTcfzEIzP+1niPofAEupDkx1E8pMlZ2iBWbdqZBKmfYBL5Ic
weyRtUCyeujK+xfECfedBDk1xp7fcG9TyRC4JlOwm1vFxbxwtgifg70+uh+/U5of
v+0PSu61Wv7l/W7gfxdqw5QUPTQgud0n+JYeMHBs0kMEOaSO7P2mLDsuq5R7Q2GU
lM0uY6LaYXKdkUhdkbUiU5XvvPnezX2bwASpTDQ5S0I=
`protect END_PROTECTED
