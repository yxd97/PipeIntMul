`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzX1NoTmyNc1/CjKa6f08YBxGzR8CZnplwXBcU6igHT/P5COUj2iTabq9PIC+dUc
en9KZ2fmvFL1X3vzR7v4/pqLEB0nUxUPsqbWXWThVylfwXfdw5PP7dY4JpqnESiv
7EfeuqdV/j8V1AgLwi29CJcqUuV0JZP6SmCGKuDTqCqdH7Q9K5wJnPKywFK90PpR
U60i00WXr3aj/I20+VcPNqliRyw03tyPF+l2xWTZtJwQ0IXFHbk7qQUOFutIx2MJ
GoTGV6seK5ky1eaJlZVUotUgb9QJwie3Jkp0PayJTudHC/z2EkAw45dhI31TW8rO
5uFMJlzQzSIFz6w7YZtltkJ5zMrK+n1Sz1d5zzO//bEmLshllCjb+Za2+3cPzjyq
95uvFbobMU0oHnz9frrl9Hi7x4I+RLhBXnBj67+tIsyXnxuy0T/Z94R2z4hwgIE/
ahsECklcjlA03py4GbBT8HP3LSe40MJeG+vcoUR/fycE7I6/rqwfaN4CE7PCzLkl
B7KWrlPJZLRqQs0a5SRPXruMh+FpYsYOVjRNz9ONatwCw1NPdi4S1/y7MBA9JwlL
YUg6wSidipg0VMXjeD0FxwyFY0fF4Z2u23Cn9p2tmJyaGmaR4EtlJ7DofaU14nFc
9bl6zMyWPQ4fqVgPG548SCJeZ6/mM7lVLc8G4i3Au22BNgsSO5PeBT3JAblbjtSc
0Nl258/Ke1lYLECpuPdunlOY+kPmughU6mirB5rOQX0AyeXVofox3Qo9VFj+RptA
wBj+vEBAU/5o7DGHPTXAFXyb36Hz5J7CYVWIDEccRDqY38C/oeI7YhsHg+KbuSK3
0PTh+OuNa5ocjZIN1dKHkVP16kW16CW5ANUyURhjdGMQ3RjdUp9TaQy6Zq2R2s+t
vTwck7zZbLWy5MSBI4GtdNHNblax9CABLRTVTXZVLBvfrd7Hj1MqF/E+enXw3VjZ
ZhSeod4IxVKVSqN0FTmfqUtOfvmjX+mxS+pz4RgZY7lKA8mvd2kyaFF/r+49czHg
mpJZT5c5VKIaXXCcIvmgIYrwLZVScKXJruE0izuAhnSan6/qJh92ugkkUHi+L8w0
c2ILlJSUI+s25MojydFGJLtETyUDP41cdaKf1mCYwf0OflxogKaW+xqfEgmrxLMW
yoiy8cAVzhmlX/Qhu+y/2yt0UZ3KubZqQhyRBeJZl8QfhxBwLlBjE+rp5YZGsIHb
capf/ux47AToaB2V5l3DjhPcr3ft2d1RdaR+G6oTkFnKetO0zcUSwX/E7cxVhJ+o
r0i7VvLI+zz2EtMzpSSpqR0oJp3WaRl82Mts5ncuKIHjtl+HXOpbl9PnfSP5vfIm
CsjYfznxZcxNXfG2+Bxm4iTfwTnJ1nloRAywe9Q2M9P/6/Oj+CrJjqQfUhqs2fRI
IN8BGuLZD3kCZ2IxRQ8YiqqE/HaDqXywUo/ASBJVRqbEqX/W0O7iPTxBuEvTBAtu
GxiUDC40M5rj/DknPtL9lvnHvyjICJStsMcdIcJO2pRn//fIO8PICKtr3Y7243RJ
V9g6Q4lReS//q8tD+lXGn4pEb9psdE5+UCCTJvADHX0Fc+n/qzpiZkKv5xho+/gp
8z0PuHkuhp5dthi/3a/wdnMyKrySuwRF10KhnH+k5kHC/EtOOiaWkTMOd4J8FFdV
DnnGZiPRgQHthcIY3B7LpKe++0KnE69rqFH2jXWHjNw=
`protect END_PROTECTED
