`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lUC4ZthyGQeQoS6nwg1KwBDckubgFgGYNOwQd7rFwZMnttT9JhVUmxH86WxPNPjr
k8LAReAcTufFZWc73yT+yqWS4OpGts04oKgyJpp4fMi2NNJQ+cquAxSa4NlILBqM
9r6Pf6HjEPP1GZBiCMup8nrlRvXfS4U4r+Zc4NWJswnaxyTqOvX5jqX9/arDMuWI
MsVgMhXqp+VrnLlqfpjFKSEybJiqxzl2dDkc9B3hCTY+RQ91fgXzulMkga/YQJfL
YMshnLum1xVyJVuN8w0mrHZTICK+5K+nFoJEN1WLS43C3J6mJKbvIZhVs30jfPoe
`protect END_PROTECTED
