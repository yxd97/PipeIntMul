`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9DOws48J4eadbrO7Avhh9UwOBcZ/SA+LzM7642nw88QbBtS8tUJok6Q6L7CReFv
3qd1Z5Lv9s3yIXli2Z+W3AxTeQLmpSePdKklE5IcNQbT/p9pX6zYm2sK45Vdvz9h
MDFsLW+xcxZV4m8/Tv7X2ZVTEEwKJ4uCtxua2tMWkqFjKuAUkLgBlJhpOffIJFAI
6GAPvlgvagGyryh2ZMBcEsY9M0fm4+DYPmRbxI0DmzSbNj8cyB88dlLZe1u61Q1l
M3xvUB01tPOVDET+j55wt7iUk3i9R6YeT5BI81EntsccwO3VV93pfPArHbP7e3c1
XriSezoA23RqDpKvG4e9SFHCT72qzG53u+WFfGlHhhWZj8a4qdt+kRe1zLQEq975
srXOBFbLWnqiyzjv7xMMlUU/+RQXYho79+0vmU0QGc/56+E8S34YIgORkOeXr281
6JLAc2uKbd52A2YruPT1KfIKU01NAJG0yMTa0JmhFKof/mdBr1Fzt77F23wi2khY
gcIKs41YoLApY+W/+ayvH1VYKZZEl1dGioCvByWvOdFOhjxTccXNY5c90GwvEMUN
Fpns9+HqfbOtETduwQYXeCb9fPCtopsFIxOUb4E07Z0z6sj/AzoUfCRfifeXIlC0
WvT5FysLaPT9vdFS0uzRFQ==
`protect END_PROTECTED
