`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDt4FPrAk+wvNBvYzKVp36QL25K+I0i2bfHQ/Q0zPlY9+MvFS5cExwmteNa8y120
OIDWxAKS2fw0gb5KQym3RLqjVeg48mZ0yu0ayeadQVmKac5A372QdWp0H9JDfGiC
WfsB5CR/BTEG4nZ+n9EbhvhGozK0wUFYwNATEgXlzNQU1iWbhByVxSxXtgGQ60RI
iq/kgpg6lYZH1IiOwaIEAa2Z3U+RPHwTVbRYpWs3PtXSOwPxspMScwxYISOgMKFH
MRepTzNeT27n5kJNvkBYB0hreDjy0iTudeGuJ+m7lSQ3I+urJZNFPlD7Vci8BAhG
vYe13RU3qMUwf+DSdd+6HEVOAIlM0/63fShdiAKtGhnOKhMZEx36SNqPnEAl0k7H
hDMKSJbcyYwUaMDzruswZNykxX3ft9QVJKmlHIpGxF958Z8coFTXbP+JJ4aH8QIq
mIJ6jDy28uroqtbnHE5wfR3ftHeQw02EG9rWz3YgV3+Dt+KjqCasd8MybJilvO/L
WKIoOELl3P264DjYapdVY5C7Rmgut9yw//LmoE106D4PzkKZtD7rhBCmEQM7iQWp
s2lxO/DkGXDVzYCWwC0ce9rafI1AqIPNZPOol0HIbwP0OnTke+aE3dcvsrPcpboo
wp7YWWxcqQJjsalif0k6s4906lpJzYtU3Q0nx7kuFcq9H6SGUFTGDZKQjvMQQ7Ti
`protect END_PROTECTED
