`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0zI6Y4gX3wYxolpor6g0QkjlMiA++AEeTvu/+e7zx0LvBMPiDpJqA/V+/si99DTA
Wbz8fywUMKe9/So3CNZ4lpS9aap34meTQ60f8bIDz7XCk6dlMaKPfZxUGNhGieK/
QcbgOBgMNXPZmyWkx7lzPstQ6trdOGlOsxmcoYFg6OK95rYKkkPXeuIQSm7WmnSU
X+96CUp6qq1mDFKbpZyqZFv+wn6aNBXKhMNz3Y0ofomZhobb9sZkZ3SzaCEbiZRY
zu0RMbiC1/xC+k9sscduvxq68nPs1zsuhSHZZ5ljmAmBnddU8VhjLErTcujGCu/k
+kfO9BlgxXSsrH0kgkBU2F59Cl+H06m+mdnzWbDcp5oNzJO9w5D57Rd960MzAC5/
Gg0STqqjifGOUj+aRs2gVxf/DSKPIKbz4KrLJFjBToVEloKeCO9MXdHbMB+Bxvxu
5LhsVhQAoSHk4E5D5P4+CTmPVS5AjDS7oUmfz0FxvEdP/xLZTY2OSGU8C2Je4ypT
fioKvGuyzrTSsXZx2SSCn7DBnSUu/3UYsYY/090c8cH1oQ0BdZ3opq5mx7yjUiIq
tdMo5QRbdFaV6mwQUBHYH4B/ycbf8FsUS1/A7y5j15ctDYv+M89qEmD7cnlPR1vd
+iN29lZh7YupPN0Gs7rvsecacGh55aT2QibiqytcjeBzbj5/PR19ICt2dciRoIil
LLOONYdRFavDNgQ81zhti1GDVzEtWYu4vUa0YR09DBef1dsRkwwkIkXolaMCUGkE
FE3Jyv+Hf3OzAC+Ok0KQ2A==
`protect END_PROTECTED
