`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f6za0IHmh0ErsXpGkJy8fUQUz8m5bPgLJEKY2Izibcm++3gs9poF3WpfVyKbgQjI
Pkx3WkpfI15sgu4gA875IMJzOMbcOFeiT94ScqWBalH+H2eWelTT5CvgmoZ4A3CV
R5VBi4MJvMRwFNPh9L/1T9ybjgfWK2qSJh0UcDZimbGCHcLPIhCBIe2FlJyAljmA
vaZ6+LSTnUVUG83LRkxvGxatSRbUszzQm/WjI3cKG6+l6ovfJHI6C5tWd4JhMibP
GN3xRaC+GtuI25VcF8wXtHarL/KeQ2vz+Ez3idcgdPYHjGdFM/wwETTlsefa40lA
qh4UiHccH2Bq/PnXeLyKppTlm68KTw1nECIW8jt4/v3H7znBt40QjVLdVLud5O1w
`protect END_PROTECTED
