`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dh7jMJ3nxkVIdGJ/pp7bZZskvKKsCc8EIKZRbJ0SS4j3TNqhDh4q9Vsu1+3mQDCq
mE+hoaLjGxN1OxxLFoKGgGgz3h+8PEJu6KEeombSSFqaCuOpa+q7VLOrttg1cVtf
88jGG/M5wrPf9b/WN54VfYFpPkUBwKzRj6jkj/0/DasVSoK0ciwKxlq+pSD1fAdk
x9y68DcYaIs3j3scbBzqeSzEuy7UpHcdg3OiYRtH4oRM06k82IhnXzhtCxqkXX4C
gO8jA58mDZHx5rmROQOnPPP0bZBT5we81Mhd7S4b2Tq7D5bIrG5RPIwywxA3VrDH
wT55FreIXGw7dH8/LopggO1mMHTzz3ild2VaXVrmojpQjUd06H9BGKKlL2TdKN/1
x/Dk7vklLg9CZkU5Lfk8AlSH46zgxVlpH5jZsXa01Wj9hjOSiKPfGfqRlQPnbJll
oSEa7JnqEgyTArJM1AvxOV5B6FLcsHqsEB4wgDS13oPbpMrIJoROwTNhhCUFnvFk
Q3AU/5jmaw3r7mlAGXcSg5wLl8KE3ZHXTF3tcQmRGnr0VmkJf/UoUJ8y0GtegKw3
R6/AIZiXtr2kmzKJZWqG+rZuZcoh/v8niWyP+bz2/1Z7fNI4IOO3nS1B74VHoIKO
TQj5MOOYbyt/4d/dJ2NFTg==
`protect END_PROTECTED
