`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/nUkAiB3QKBLOVf2MPvX3/yxKM8TEBRsOWVsg5WaubLqzuPm7cWlD2GobM5YApf0
2PPRd5M0aqM8oGTeHv0d1ocUI5vAR49eN2R3TtQiuUxw1AhPijAEVkDMAE62TWUU
3w2Re8CGC1au+10Nl/rXEJqSvm6gjo5Aw7IPaJQrmC8+PboQ1emXWD8/GvEPimov
d7JWb9eYwBLh/PDc0ntq0wmn9Td+afnAdaHx2xBqMGXngwwV5y3bI5sQkunP6ruo
3vv48gTx8BvVCsj7NMEZikWvOk8g3lvM/nfHtX8U2+zfLCxZN/JPcMEUQPzC6pY8
9Anel8Hj0Jig5bzw9rDzqUh1yYRasyuVnAK7OZlglUS5mqVixAdZ3Xhpt40PhLm1
/7YTRbM3cDOuRGjuZCI62DHLbsKnKgHfCaeqy2dxAk085km/IPND+yTf+/+86+rh
`protect END_PROTECTED
