`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5AJG1Tg51dShSOb0C/FDjSfe1Pq70/HTxx8ED/ZPa+SQ/Z/aGbR4uSB4v3FLzux
LAqCRzcQatGmw6wjW/fsPatw6W3bN/ZadEZHdjmher9y5rzoasY7E8PCzFQfMQWi
ALObDrzkJ4n/LGThgZq9ro2F5Bp0ZtAAGERD51beDbx4YqzXlUOa5yjRvXDnhmHo
djZKuxFIRGI3wkJcUBfNqql0Agthl8VZRa/izlHmE51/2SLJ4ryh1UOeMKnFrpje
kIJHA4fKa3RkfUvErTZAr8LVxkORVXvHIgoV1uQe3w8o38sI7iET0pNF85OTSUUn
mzj8aUvwqkmDuqqMIpJAOy4dFGjxNm++g3+UAtwZ/0enWcULlEh747Bm6RwW8eDa
Qv0P/oZm8un1wfdJ7ZTJ6Cw/+YgPKFRdWrmS6cTZxCAoL+RLy6Nx/qNtQaLvATuP
JJmaqBysJcZTbmF5mU2Hp7OqGBnweBM7Y3PH01ijZEK8BYyoqw58T+Y/OyXhEkyK
ZRtsJ8FfyJM1zlNFFBmL7dAnbBl7AUP7xS458//4Qm+eieEzsTTAM9pcxkxix9w4
ShclwjfduywsQBbLALJmCEJhcw9d275wQhwtAwkqo7N2DlrejEsA3YZCEQ5cOhoV
157+2JrgzWqu5SwKMsv7hNHTaUKmhdgCpCsHmPx334GLZL9aP9JybSCaE8CDYsge
GpJX7fiDWeBarlpwsztTsGqyLjMo4Vad/dsu3vYglMMSUMt99fa5ND/3zhPujuo+
5BG2mIz8TOLxNIXlwK2tGXmLoj5I9dSxSZjJyZEzDExcbUhdhCCXcuxK7E+OQRm4
hJEmwcw+1SyTVLtZhoNyIzEabWvXK5+I9r/y0UbFvuEaFUT2hKxZZsjroRvKuHCX
YBOQEufV7lixtMjUg9gBTV+Rkq4pmqvqrbN8iouBGPB/uCs0qVhhg8p25w54pfl3
yX7D8RP7ib1Z8+TE5+EoQFpgwizzc0e3zJuLfJ8pDzDXhjY7k0NfNomcvc0UnHFl
pZxIrm8NHziL2ZHHK7fQ1pTfriS9AmCDwbgEdX0Y6vF0R6MQTeytCrBiJ3vQmjfy
h+jhZ2P2tTCZwbH8Rhe1XmqQf/1q+idQi6mYisMAauVT3yse0pwz9Qgd1TCun6Bn
wlJEucuhliW9bqOeVdHlf4YpndYz8whAeakfrXnvY9pdLOWWYk9fzWf1f8QnBXqE
m+awYndyI4sY8jFwlj2FniWIzOp86AUuaQiCsk8uFQ5rdC/lna4wcFdXT/nLpDWK
K+yy0Z4EDUGZYnzbVVcxyLDv8egy3YpMC6bD+ypRmE0TbMJ7HZAbhb+AwVh3ipr1
e0dRIDNE/3WdHNxTtgxvZucTisXU8nHVSu2swU417UU=
`protect END_PROTECTED
