`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RlyF+Zbo5Be+qRIiNBFYqyvd9iYn7MtHvt3COKakZe4GeNX5t194rQAHHcgEWrco
yYr/Xw8XcHrr8CXxwW6u0yFKH8HD/KI/Z6TlFGkrfK9pOHwzIIKNFEWfqPqJ1muy
tYh6bzSqJhYA1peYHzN3KyWxDghmCvvXa44+C68O96RxHEbvBo5NvgY63eQYnMcC
x+Ylr2PQMDyBsjj1+wHTgQWm6ZJd2bwNUmPf3xqzu5OHRluhnx4pjrpjZ/VAXUQq
L9txGgivnQM5CplAMUAdoYIMGqdbZHIcriERHnS/f8FpgSAyB3ni+fY28w53beb3
jBxbwnkCqNiMA7yN0rkW06evyAIxeWa/iuPhz9tGHK9R4o1n564xemyFdk/7H2wH
/aKYDuz4yFmmIA3g1ikTnhninaBWujfEV32HRO0Zo7QTr55hg9xu6ECR9bnlF7Mu
ojZPs6al7fEzyCEZb4F1qppLnjWFn086iBXPjrKUgDiggoxlRhd+JmFLjM2j/17K
PNX1y9tB/grbm9TG2cpX0012jui40MAACfSCbi1jY8ZRAUhL6xUZIAf1QF1LupBx
Tv+oYx8/WSouLrX85gYtFyVJOM2sjiB9WNdvycqSRF6k9v7f+NXHiw1LUC61Crbl
y3hUipCzRP2H2CACPV6A4IOw5raWEmugEc638qYwl+nhVsT072JFox8oNvlftXTy
21nQ1UaG7ISCFnkEY+GP6xiyGNjMkuLUA0+wikmYzGh0JWec/BmTib6uF0sK2v5e
SHLf1mV98aTP26D8vdxaT/wcuxJROsDlL+JeUrnYfuYB6bPLT//yfYL8PgMzLevw
Nzij/PTtRKyJhfsWMDsfVGxS4gnDvBB9y9JoZW7Eg/Tn49t17AM6xItHtWY2OLyO
8yUsf+ZJd74I04SfJHgjoMk/2udwyLlwiFrXHhBNjIJEE2akbSQEUWqG1JCl0Lf0
WnTHWArklPzgfDR+UlnFNoa8gbQRW50lOmAX+/urlX4eds+yHRpFNX6YJpfLs8tu
vRPJTLAySbC7bUz3agq/kUyDEV5hpmss4mhLQsWWrEa2a5qvtNHJoMYRhZkRNJ3M
QfSPJ7RNX6pMCpNzBdToGEuQFNYAY5TPIto2KeSzWwMhWob5/tHklRpnNxwj35lP
R7fNtOHZ7WlRHfVKhlUnm+vHB9LKbc3J9fk7WPP4k3ai8RBDJAaDV1cfhTWjr6k5
iZrgjmRsspsML1CV3RcO2lMoIG/YDxF5kQRr1eAJNCnXAhKaMQ3ir720LpFWg1q9
8iEZSJrjaN94HdY27vtTi+ajZoW56wA1rVLlQa3TQcAXW53HIsZJBnOGcmzvbOni
1Vj6u25Hd2lCWK31ZYrzrtNlAEcTf1y47L1tQTxhH3S3eCrWsE7FiRzevraZT4Rc
WfRpl78+K/dwLJs87kXZdrPKblI6eh5LCzDRBHYZm+sOz8w+p6TUKZbffLle/7CF
ERmJO25CY2hGLuEYLO1YG2PzBX2q97Vz6LiPjHgSBESh3Jdpi02Gc9xfOz+bDeWq
3zYzYtlirK8BAu1kKDYmW8IEBFz0TExAANnGLNvcNJBcMkifPLTi8Q+9ST0+hg2r
mSXt9Xf0sXrULYhmHVaK5otNWNqFjokcVhOEn22YwJt+UNuqKNyeDSnbmpsdj3cb
Y9hZ3jhTGYFocXkuOiriCaI8jGxrd9IwQvYxoCkJks/gxE7UeyUCN6AOtxQuWfof
ZVwa0+U9urLWVylVx6cI+HoL5MyA68eJmqAsOMphWJMFo5oD+L2unZKvU94scF56
9TCpnr7YALEfdk2IMgSrBhS0veuDWUJcY0YGes7nKXt+RhHAWvXd08VPb0DNoWkh
1RV5Zyy4hqisWI3XukffeQUfF4DLZtwo3AgKR18VhKA+bX9BwyA+ciVRQwVOJasc
aTjH3IwA/cmoms5ymjMh+KndaSd6v+L7NiGr/3v1Iw+5PHQ8KslfJiWjmxfQtJmQ
b/V6chud7YbAvsbQriZRu9ckJjIKnERe037WpFKLnOGj8gKlVDbR7zNuCSuoChCG
Qk6e08LQTSZ6lTm78IWXwUV1K9H8kWME4dDsRWwwngEk6OGVFyd7ucEQaV35sjo4
DEKt8GTcIq5JOV7jCU2NBCmu9HA6jIeqngiI2d/p0AHU9bWxzhmbJjRxaQdLto+b
ZPUCylEzLK0zaGy2Xha7WY+H8S7s834uhqpiYO84Zm/yguM1b+x/FNq/pXfEZb6y
/sFJNie7hMPwF7Lz/UcRtZXd21/k5HYB4J4TzpzNt3LWiyvHTFk/h2PvTvg90iCu
iFyLcNB+m8deLXPaTTAJ0BRBN+kxJuk4cYbg63TlGW4xUObwdW/Syej1Pc0g19gM
7qfUONSGUy+LVwYvtqUrO0fku26eV+Y+/eiiQzicmVjOelkRMflNGmgMWNgezeRs
PKFHHah8pqymntpDxexB9RtE2FvrnvyKhFNYqC+m8w6gsAgpJAPDBheDQ60ta6tP
oGRmMcQPoF0WhFuOHOzYL8wNFdv/bM9kKCe/oCdTv0mRblbvMqhyTs1OBy6J1RDE
f9jfdxnN1holoTAY2spzIdo2f3inLt1D4axuLdaQrJgPdQf9qsMSlNtM0YG99xoS
ERj0QqHYh7jZKcHJbKf4fjsnwxXH++wpUq9y6u75glRFpjTlKPMgphfPlWTLudCo
wUc7+W9s+LawKm+BQBGr0ZlaANzV+sP8zhHKdgV58IyTsmjNYqp/WUDXnq/UPO58
IeI//04PviPlrESQ8aQAFAcPkV6Bwn8utjuQHkXTDnWmvjRLLudNT6KTTQOymQVl
lsjIZb+FKbY5G7up+/asNpD7rHyVst/ccq2HmJiAmuHaK7+PBSqbKwDnICKo/ycL
Pgp6Hh+skwUNzIGDIqF7FKaJmE9AHbZjQkLFT7DbNp/6tHTYGu1wPWQH9Wp/b+u6
Ikktw4Q03QaVl+ulvGjHetS9Ze37IS1aR1OqSQNCI9PgeMHpecdtG+AtjLlitBcV
wEhIWt4C4i8hKyJPnwVh6cxlvWgpdp3sEMkXflBk7IMB0RrGsKDvXLGNRTMsCYzj
Uy5igKkriIe2P5cC86cWWspp/i9mp5T+usefajTJLzVVWAe6SfF+ahTfEdeTgqFd
luPVgxlL3qmyI8YBBoq+Cpc/rcqEU2mT626rPZLBhp6XS+LwCeoQnOiLBvU5sT6v
agszovrNCrvBgrvOiMBoiiCheLEAO6a9iKhgmDXYGA+aNZHZe9TkHGQc8dPhocbQ
bRlBhS44k7gjmWfDK6PoO1z7j6mpC7ohoPcGkta5yw5nXOTzNBJ7VI94osjIk/O9
vINmJf4Nl7CIDoK4ETPg+rLJYzB5R08MoR8ElYWsnTtU/eLrjbegyJmTMMrYG/Gf
1pmrIKbcfEeR6tMSpeiZ74lkm7t7Tlvq/mkiHENjaBkxtD6mxVmWArcWYiU6adqr
tFjd7wyvzyF1Z/SEz2avsndb8pfJlLEEZsIS2WAfluJ9laW/PZnXVL+ET3K75GCW
GzDRAXlIo3Wd0u7/K35VUTXVrRIS2yf7EkK1++bI33zW9pHbs/8pJtjxk/vPmpam
YW/0bpc+fvqNxcvrizRJ/rRrNT75ZFJoUBKaSSmhZL8vhoJVgEJ+wAGV0gpHpAgT
Jf2pzIOkbdUAmUeyeCRUEzhmlPz7AsjR8pVw93GFyxEvi92gA0V6WeByVlIvUlq/
qC8BeYGySSEv8ccHrSyt7z0MzKa/hHSTlwlkJ9u+OAwVOmy0ZL5WSvP0cvpST+0o
clOGvuAUM0tBkQ3nA0iZiN7hlPVbc3p1rbBoSLW9nwSRMuWTIvqo2OtBjiffwJR0
a/ciYKyB/5bQ7vIXl1hYNp7L0MS+kkuKm/z3jmAoR2EIDO+aNGzmYBeJTjZeKC0H
+/1W7LJbIJQHikBUShEJSJ3QTQpLAH1f/6PxZaeMO4IoIu5/SpzhAJw9WuA9pzHS
1EUnvcxwYHAuDGQDtWTdty3L1Qm6NS1f1qQPhMGcn/JxBW/3yslZcjx7PCifg+qr
Vuv/ncx2xkkMbD9l8jwldenBDkT823bV6sD8PrmHY3/F4WgxFl5ZZ2lfiQxkgHNP
n0rIMru07Dw9Gr82xQdpn5O26ZI0XXLX/tbzxgmvT6I0op+4Zsd8Prd3Z+nd/7Mm
wMM5qCW/gwVYr4crjb89k+7hs75vujdoZ/up4g0KgEiji1HuSlU8sVtqte4PgeQo
1fMaNbm6hzasM33vlfnvHAMl/TzifcY16QLPRyWTCQrHim93auT7kAdESj+DaSZv
zHfrAjphzs2iw19H9UVZfDzN/bZ+kdr2tIwkugwgtlPl+uH/pcG3UJIkqn2VDgBo
ARZ6NJtIcrJ2ABDCN4TGLVjc4d0b2o9/cZQ6uKsqL0J8xIBmQFZjodXag7blxyZB
`protect END_PROTECTED
