`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jEIcSaH84nqyCiiiDo/KtrE+ozaGJgUXL9Or9HupQzuKPhSj44h/Kgtb8MYcHXJu
O3VEMyMBLhgVuKSK4VUAE2d+q0GqN/HPhoAbqpxBsmRaFQWDenDY/m2Dtyx67vGD
WvzD6ikYivTtXiL0BRw1AkprtHrQEcU6P6FtG/udu5BjMyZZnRMBNMqTtPgkJ1bj
78x/frZS6HdRUju8r23CMmaKkxHCB6li6BdJiEm1RtDTp0BPqRhz1X0qh6/s4JWL
o6pXkjNbcE75/5Ij48+ULRTafGAwXnmDuU9RkEIxIuWpfvzVRWn76xuGp1Z8fqul
IS2bF3yIKSVD8uIu5pVoUQkRBkKvqISDIzWDn7wsMqNogcr7gG/jtiNlfrjc4Pvk
Nx1K45EXyYtEoZqca+xmysfrzDnmZOI/U0yc0wbVQkpu0mZNthDmVNx/jMI58fwk
bB8BNcaAUVHmRrH8vZ1vMevNIre/0isZOE5Kh8Y3lbMPD2IuCGqTtzYJp1BjAmn1
sC0KApRi6Hc04dnaUUmGk68o/NRbmcmV4C9yk/dgyUYfsoB1p63kozJgSpANO097
Oy+JVfd1OCBb+ogNNsdM3RVFpNNqZTQuGXP3k8rHk5UvOUsl0qm40j2XHVmE3GZn
zvS/fPxFondoJdKUobaI/ylgHmDH3O6mPu5ZZRQyGfq4hJxhqOBGTRpkhYQJlvJk
7AXJHXQNF6pU7LbSrKDAJWpkdqVyR61fqFd/3MAf/AYoM5FOPhg0O4MPcsf01Un1
1SyBAvS/z3WDiJQyOjBaM8WG6B0PWNJy08Be/WgBZwlArWRxPgyiLUhz/KiHS4pu
zuHXgAhZNRs+OySg0WPEQpfFq3/NEMwAZdOpEoMmPBBRVDLFGNnnYEH7T2khN09a
poIlLU7f5q79LcNNOIXjjuIKRnXnHUJAskCIvJSq4bq3W8X+3hWIsTCvA5gQp8r9
RknXNDupkSJshruVTlL7pZzCffUJnmC8/5v2L0KSHJGKh3GmETZi2luaPnPh8Qvb
wNcIm//IcNxjjsLln3e37c0ZWJZjxs8mDoM3U5UXK1myBaRKQ9MQdSvoA1osKD/R
QWPxVcGmGDrNY7H2HuaUTWPubTuHKJh4jteWoMQiKSAg6pvgWGa4cbJZoEdGQ42x
rXVL0b5LW6b7meP1GGKB608QzkCqOJJUc2yxkihKdFN3YQqD4PPg7Qw7JxdlyzYy
MdHLRLB90bg9mQNkTi6cUsWR4fbGhlNAJKKXAjQW+1OVJkE57rNFTEqUl+/D5mlE
rTtxYtafDon7weuSSgOoBKIi2vQxbbRent2nJNGe8gkOPJJUxrhjxdgjcU1BMQPP
iE2+SuLzRY6NDFyM4xYVBu8TzZ/JmnzSQGeGPyuc+1tOItJhWC8XxdIeRjs+9kGw
+wOGBaqzdtd5Sm1F5nsiElvDMr/EEBSAlulTfMohSqvfMlVLfWEXn6j0EP8Rm3Gx
LF1oynCFdyM0qoznpD/BwgElIybRXXWnRPdM2/wlUupG2286+Rj0NS3s6sUXoPyI
EStYzn7hFuWs3iTGctzwpiA8aY3EHjRp5xpn9MuqFIcL27MQO1MAw5cA7ghkRyOV
M3f3VAsSDgPvE4grcg+LuJbrkAAVJOhHJzf74DsKyGdr8tD0odg8toc4EO4x7cla
IUnysumH4mnO1za39wUBpu6C/1ogIzAgVjrP2xc4BcOxNKImZ9GrohBCwOTXzWqJ
I531mrO+gQinz1/l+IJiIktqPiqbRTV7C1kZsCrugJP0LC7bEUh2x7amZsM7xhua
wJGcKEz6niRZ+ro9N+BzCPcJHg6ZdqWdUC4CC/7hE7D+5MLBJYuvaVRakGu1JN29
htcNSjmx6zP93uBbxUaQ8YSXV4L7cOXCsTBWAG19O4ZjAW97BLjit663PB9Fqz2M
y6C/dQkIqh4MflqhwxcgAASUMn4DXrjze8HVXX50V4yeKL1ZeizQn+8Xh7CzPdjN
pUU824hLIo+Ji98IT2kg5woE8ygAVs6U4P5Mif9HxnPSX1r1QFm3AlAG0rfCNwsU
ZuVBgwXkxB/vQGMZ/7U92RE8HDqTDCrNt1836qSWy1gbdg72I04ckFHLQDlsJL6K
DayGEAHJPi4ErOy0pPT/ligK26E0oyvff9qIYZYnCbnSXgD5dxUzh4S8NedjtFy2
Z4rvtFsEOhpf3ZT8Ej8zFkblUX7OR+x+JwO+VrJBwgXUljDFgtxenWcg/CgXPUtz
yya7Wr4NuTqgdMJTypvVd+a2oijbQIT6p6cwHLEZk4zH5eSOirRQMqOAJdgjK6o2
U7jqjhggKsSykJlMBeRueHtwbnZMt9W9F6lc2tkptBHu/RmLhUqeizGEZTs47swK
0J66oNu3NKfx5XgAHiiuwHQVT3DZ51F4RoveVRF03ildEBFpES/OA/HpENgL60CB
1GcdRqq1EG8TWJ68/OvrhCYI2tRIG4iwF5huI9YhRM9hV6Vd0b+FTxi2Nen4cr0K
jOVGmHEXYKL+dT7Ndf8PvGoul9bWsr1CMsEem4PLuy3X/wijAajyliY1BNerOh2R
Ktwmu5VybIDkFfxPRyAjZXS7T6P4lklO6TXycFRv5bnI8uFTUhue2hglMKlTnv4c
a6dkHDJ2xNGHsVAw2ic0LnEjNxiQnWR3caE34BgE0c7at6SOU/etYd/VuCjPcHyO
wAqeg5Nv/efmX7bVN+ohMPLnj4MCkNIa+YoJqDcqPDVMmiEBKh7C8fc63ZnGIwjT
qNgNmKG0rhpDAyXTJToTotS77m2M/0/D7JA9CwiknsZ94AOOo+AB9BrH8T6k6Gor
kyL/C9h2f9A4XwNQ8mkTRmaKbLw0tGecm1tJ0ljwLhJKGNrhb9ZoUGV0bi0N2XBz
z9OMzxMnaH0TavOqbrf3pafXq//iyOHH3eUUiTGjzCmDQZgxvq+I1qC6MzTGWlUf
PTELjBIU6iKSPb03r2J7AcWZ7GOepfwT1oAwvFbG2ebRL6jbFRxJ0RYDrh5doLqT
3tA/19cncbMCvFBiTG+soxHD02xnTdZYj583ZwJRTHSGQVCtwb49Dpmq4wfpMKM/
qG9XGUrqppT6tmJrasYFnowPhWFgWhNBy1OQgNe7YksaLNbb6u6bdpO5tiRSUn4j
SvibrT/qMJej3N9DY+kvkh8lXfom6wmCNIWC8O4hqQnWJG40aImfqS8CMcCW07c0
IQTqfQUOeayHY/B14IePUf6r0I+fUwhSFBu46blQJV2lK/idM3KuHufM2VlaihTS
J+A8r7XIcEhfcCjpGugqyhY1+ZM0HDHPJyxZCaqLnHrSHjmYA/lPgiCwaUmASoVE
KIWJ2E3AlOEqjEcOeUe9ej+gsekfXNDwi5yEKICv5YYllYIjTR99aW6OS73mr5UK
HfxFZ1c6BdG5Wj+9pEsdLhBTUsfR89Ncv7CAx4uaWhjae989eoX68OPggetz5tp2
dURP2yL27FSfmB76BayyaEuEk4iMnzgQB17CwpxKEb41P9/lsaKsA+8Up/AwAS/3
AF3PuqqNA0dk3gy1vi8UWAe++NXM6mXWbatrXGiMTdGINx8YP2BSu1umw5CZcgWy
`protect END_PROTECTED
