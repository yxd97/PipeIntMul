`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H8awoQYTcjyyVINrd0+rTsPEkubyKY75bjKME7F46UMbOB7iXV/mWLgF30E6xvlb
akWRkPwhsXe0hRDKKzYslNGHG28qHNg5i0YO3Uh9xMC2gEvi0bh9zQXJwWem55Ue
togaqEmlECyH1Qr0ZGKdp/E7eR3hJK9zZY4XK3YtHhEqyYYCme9Oi8CUP6tgivAQ
SfE1ACcy3bgwFgpkG85r63wydAoj35Ta7F1VAR9v92UydtsBLR04XmpWnJ538yaJ
L1obxAikXDLswYIFCR1R4Sf5tiTW1ByDL7bOlPbhMnNCNTw2RMrcGmcuBmbzvu8r
HWe9UBXRc45C+WihpKS2vqS1iETqyumBXM2YzqVN+7PQDAzgSOkvHAxdjw/azhAy
fD7fVm3iHvTKHgkEcNEb1hZH8hZ5wVn54Xt7IpEy1KEWvuTPE+ldGAIhsT9iIxNc
mfT3c4qhxifHTeeoJblz73/G30m4E0NdjNFBdNFBQKxOYOqN1bZHwyJKF+2l4UpJ
n9VuCD6HTmydh7BPbzm5rG94J7H7XtW7bQ97JHJU389Paw7+hJRuNPYHiddAxXLS
cEEKK536IrGxswS3po+lgyMTVcqiT3db6UN5HGZ+h4yog5OqUghqzK9+dTyoZwaF
WjUG993VXZqukOFKDWnbO6Er5pN+oYIzkTJXj2KjvUg=
`protect END_PROTECTED
