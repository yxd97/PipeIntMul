`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vsq3M2yBw6XRppBKDhfv5MFDG7sgNPZ4sisw93xjGTRX7PA3mP5o+t11cCqwurm9
vgYv/tlUpp12Ab5qmMaiUuvl/qthL4Pgj2VwEBI72LVRydLL/gVjmsiiMBCC7ni6
9S83+kS4asCB1nStbx+26IfxK8W7bMQid9aEl/RlDfAwL8kTjQv3XISOzORVajHq
HNrhKIKkCLqhUDmcfAC0C0erPg9PcOMmyIYbsmtLQ3uvlv4cMYuU5O9sN3jfzxES
JGauQ8HWeItFvbJZKMNnULUbuDOtdFfP7yMaKtLHuBmEJzHj1wwoaEaXx5vw4PVo
FJWiG3yWFLC7iOs9PI90N79Hb6qV1sX9+3Y92n885mSowx5hEGI0vmQKsbZ7ppum
9lA76w9UjifYpo7v5eqJ7i1vRL/FmK7nQ8WJym9NhQ31aJlQikm+8gKrN4XWtfA7
TWn6aajQ4x78KHwYRagnLFafQUGQeqfmv1xgDctjM2ygGD8xWRLC75mVKL3xNNGT
pgB1ies/QBOCeaEfDmTuCaZRX6fYAwHZNkaULfzShJkniJwHi0y4GlyjujhX0qbK
`protect END_PROTECTED
