`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9O9qv4kge2598C+8noCsUPqch8A1GNaHIlQbQU5uk85FvGkPejImjMpAatRvr8IH
MqEFAcSwP5nv1aPQeFWWrAmm0cBqoFmaMRhbzNWLBgPHCtSd78npMtMXVAX0VwVt
O+foc/TI+3tKUdg72mp6NmGmFd56414VOBKnbXUgg7pYuIFp1Qu6w31AZAhlNowh
NSUXSTwDAGoUMaP7HBUB4kUFTZcWF+Ds2YR6AiVO0z+Xz5PDvTLNfM5fmYlHo4VP
vRDM2abHdmH46iu+HCW1VQ4mrbWmgh8YSo63bL0d5YFM3kNkCe6GhfxSQpbfgH3X
R8Z3efnxkbvi2/3IAuP4BH7DlBcavB9f4Yu7RE5Rovetj4+BpcWdVZoVmuDGCtsJ
+/pAV70Im0bgn3r2Kl7GSvi3aNqVrX4WUuAYeTKH4+V4Xw9UL3fzJKHwZ+0CLhC0
r+4a/ozP6Gym2bWLLLTy5q4Xyis9z7iF/B6MgoaenCbAWWmiCwiiAnRknfLpP/X+
ChFIb1YJxGdu3g9f0s5LPF86CTWeDZCaFInrZyl8iJK8xAaOxvWIe+GBMvPlJwz6
3hUBbtc1u0GmwLJCXlmb3gHSHabUBeZFeSeVXx8+5jBi9MIOLbDMLTHLc3RO9/mv
0EGBMI+w9uBWsabbqd8gAg==
`protect END_PROTECTED
