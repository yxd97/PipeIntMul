`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7R8wa68atc4t5JWjCIyWMmQZ4a2TWucW/1OCduAdt0PNJANUXS2Gh6wRwxVWbCMJ
OaRaJ4fKXa2cwO5hUr7hatzHmFOwQk0ASKfzM1+whUw5H7bgR/3Ro37QlDvENy6/
v7R70BP+kqiozISQtfRrQAy38bRmtM3vk7B0g7OqHluHdnHdHLi6q/82BDTb1gMH
sG15SoQKaonNPuLynFY21J9uNR6DufeA47X4AKJCaqPO9VaTUO3mObSDjS5Z3Rcf
wph/WA8G/h/IW1kg5h/rDRtvBfL2WOqPJ7e11Qi3E3Z718JAaP+/6nAiDU8gY5zZ
hFPD+4BaQt4K/fwf7AjY40tMMbwb3IViHeqn/HviwwefDng2Uy+TAKUJW2WGQ6Yw
Nzs5PWu9GCFRRcetaOH6Om18+CkE2CSpUy0Udjr6SsiHwf6Q9cJqYd8xWDjn1WUP
shRzWZOxrq8wHKvhPmLRuh9bpP6Lh6K4cxmKsKzNSWolKiJ5l2ZLejOkxTQUMjj8
ppZurftBo15Y4rnh8IkhJ6b+/2a+eT8BDd2yWxEMNvXwQB/00+d769MLs2pIJMaI
MiVyiDHQ3DDkZRUu9/Nwm84V5L/z8sS6bRY/mIh4IaIYk6W/eKigwaNvvjFlJ1J5
lQ/fti68S8hXhY9kWalzXYYGQEciK130GiPZMy0ew1Ah5ciTiN6Sy78Ky0bF/SOo
V6grJmeVwI25xjAkNR9ueJXZk8N0WwENknI1PZNEIB3dNGUYax2EtYXHo7ammh2H
jBgOovFUttVFxb0fxWr2QxQkkVaKy27TV8Wxu5N7G7AmwqV8ySeX5TaOp38GcJ6q
6jvaGbd+odeR/9sFTQphrjEFkVupUZaLIyMEGU1SHfgPw9H8FtVS5wRlk/9V+q7j
BvIXx6/UcXaIm+g9vuuAHz55vsADxBwdOfwCqdiE9Oz7KY019tPEUMT4770yTqKk
HicSbYiQhQo/AxWmrfL4ZYtvGjRcz1cu1mnccIDduQaXnLN0vNdDXvDc0Cp2usST
h6YCwbUkLipberschCE/qL1AwtyRsC1CUlrl1HJ1JXZyvcCzopBI4aK6p82nrkco
xoGHzrvSOZ+iv7NpqCk5/1bqADEPgAXC1lw2BJzxPOXKbjDetcp5p8k8DOWWBUwl
RLxEi/4+WfE7R0l74DR3w1fY59ozvpLJSq/q8XKje2d36SVb0m8SzS0/VGq6KwCY
5AKGvXUhbX1+NyJTq/Jp8ILqcMGjZ57fxn1AL9u1tSezfmNzVFlRu811N17eljty
QZBlOajJ+oKwH1mdhzo6twyvosdsy7f77xDzzOLj854BnPPUYlSYC5oQ7egyso7s
Y3ISxjiDBzwjlDIwj0lWHnmJ/Zbu8rHbW8eoRNgFm+M0DGmEawEPF6qMgJ750zQl
jOdKqxFeE1aptAL25yV/mfh6BpFvYwRP7KkrE4czcvpCG0EfsiqNSnldpaghKWJB
LrSSasRkbWzj3TVL61mbWogU7qtg3g9RMhbkI9dln785W56lQC13AGANzOraK+DJ
3+K9D0dsnLmW6KN5cgss9hRmWz8CPxhiatmbO0CxsfaYBazW5nVduf6IKv9oV7ln
OG7e7O+m+0osoQzLXRxkceAA+GEd8+U/MXQAqGwOFg+K8VvRZZXhh6M4slIuT/b9
zKCFs3NkVe6xQdP6Yibfj8Sp2OsWwQknjCM2xfiUj/MhvFBlox2C1dAr66f8KBn6
nU5MQzUVAEedPUc1PpoxBSlw/F9EraICUx5GuURgSbn4V6qgHIRuwnFzz4gWeXvh
eKeQ2IKeLI7UGTtac25NgHUuzDquSkRFoGE2tBAv98waBx9ODJ0G9QA8OrHZBw8f
5mZiV6WMDRdkD9O3G7RBKMgbH2n562Q1OsnnIzF1D1A/N5PbR3bNxQT5jvORHLad
DmjlmtV+b7Gjeg/1gtwzehgd5GDP5AGX8A7VHEE93sFD4VyyQKKGkCYEOhTB8HSJ
Npx49rCMyb+PvHrH4339SOszbhYg+sovIE+sXOuqRdcQaBEedM8yey6bmZ6Odqg2
IxebuKybL9TVwwQfRQ0DbUki/v/fbNVQ6+LgXoQ8Kx2E7lhpzwOiJRZrYb3XWgzb
qHigeJQVPkZdtOTXnApmTEUjyAaTXS6nH2NhT01uLLPW/whFG71HhmD2hA+qMXVE
cPptP+vNmQDrYqu3npYmc5K5PDpDHT/ZWYj4Wr0wcOd5kBjkOENPeE484hsNw4ug
uhlp/8HF51j0Vr7qicefY84gaZnKxewfLC2oieZlBgbSdyxgxrMJ1kXolXA4bN0/
9sRG5ANMwheR4j9iDWPGndepADefVkev+SdQbxSS2BtaFugaf6bm1SJ/aGqmLhaQ
/oJQMEnrkhhDcVI/VT0Y2ASSR6Aj88ZBWndwzTTjdMUvMPzLaO7hIhwNvF2fcS3/
CW1WiiYk2iQKA1hstdsGyVVSePQm7/PVOeKtKV5ERFqtrypZdys8mZ5QFRO5orZ4
I9l+GqEXW+xnh6WlOoS78yyfPw1t3XMwz8rboV0BdvrwYkCt2iqnS3ZYEDtv6ZW2
CCePQsGD32GoYnMK5tMM5WWI/FSHqmyOhQcb1tGSxBcrPT5tTAqfxoNF6NtOTMQm
Txv3G+FteaT1vEqBZHX83NviI1T70k5yJ++cgK31H+TvNC0QwEA3iJ8Pxok4R4aE
u9dC/C6NP1IFE2I5eaBcC0P4W+3gD0E1a2RK2ZGCShenxrQd3TeBDaxkA1z5j2bC
bqNFdw/IM72aLLe3dYfNyJLtjfRbkkxTOfeA53nfmuerJRG7uI7dN6tqU6S7hy5w
BCeotXuR8vcvUQHoE6Tyv/+ZmSflQ9uu99XnrpN1K/y6sX8rxE4zIsnTZUrly5LQ
TYBmPBWfD7wSqhBeEj7Tampj8RREwQhe3sBx6QLBjgvvmi+s2uV6oJKZQhM/xZjk
LOYxoi3fA3cbAbwsHLOaNqValSr4N7jcUsPinSiUxwpxzwpR6nQK+gPR1hu5TTWF
YVW6ySobH+Dq0SCAN96ADPuz0o8+X8+AtR2TJPmrSizfYAEiv+HflamG8AZ9bAd4
1aDLcji5uQd4Jvt3imU2HSTwrX4mpsSsuq1CVz5zDbZV4yFUnZ7HeaZ0Prby9q6S
+q2hWfuEg6FKZ4CgIfFfUzO5c/3qDIVxjteikXC2ibHH88sjuLxA6/sURlKdRloz
uZ78RSAGdCg/NIrVDs7xtAo4Sw4YY1lcq1sheDgigzW1f69hcm2IP/T/XV7ssD9e
0rCS6MSSOrOtRxq3AiOQ5u2+uxCQqK9NnzVSTP9d/YFCwRJJXOD6z13phUuyBMrg
EXKfYbHpOWzpqcx4pREQeGRohkQpbzr4jPK0O1ADVWdJmjHECAxGv8gZYzJQ+WV9
MgTTaEIkbI6ykhzPik7bzCLsZxmG+4wHSQAdgi3n/71lZMAiRBFN1IOXKtltW9XT
X09u2i+PISSZA8yzTobjx3JYsNSEf1CKiZOfMVJpVSjRNHF9EyWsyKcEO90KBS5v
DvokjQWNOOkWWSn/cMYJdSZa8Ka3vOlIUWCIW5pfZeBVA2jb6Op9V8Ls2bWJ16eq
djL0Er3IC7FbPkMv+/pbiruTAgs9eFTmJSn0dMiiJY+1La1OXMYDX9pIOH5zMkZS
/SpShRGi+U/UnczexQEyl+R8Q0SUUKZXCmf7JJu/DOyE/rwh+PbcZivOwG8mdcKh
cmsa620lGaiA24hvsvf+dd7kA/7IKKYfkaCmc4fidbfATztk+BX9vVxl89DlmAJp
X/PTi5NXpFbDsWpNzQ3hOwqMg2Vuv8s7ZRXutbC9eYOnXnW/IGg2kZm0QUlpdkqi
JlnVXczJTolCE9iaHJML+p8YWDKl+qVIU9+K8+JVBa1ZNRW9L4UzNI1H15ZFppJE
LuxWTpLErSL0sZcfl5WIVrN/FEbO8WWDtTUBgNftSXMBc3XaztabSVW/egOKbXDC
Pxt8MQWJgx++dY36EGF3VU5ElKT1wDlfu94CsLEBCfb3oVX6+M9OsOiy0Yn4iup9
gHFdgozzLni/76uxIz6JBQBJkTGDaYXhVSMctl8FUWJr6wFdv34DEDK5hlwPnLSW
3HY4xdSGVTEM1ONc56iZGA6mLHqNDiZp977tjTnDhyEazMuOEE7AOQT33+jLMG8c
h8r1L1U4mYkGYX52Y0Xpi6XHi1Z60GZAmdDd66e8Isye52S/k5tuY0SoTNi5v9HR
k9AuhxZdpjGkrHiDhSm0bK0ttkxAb6wxI3gJjRZTBCWGX+mlhZdr8j3z7DMeLjnO
YuhbiI5HsiiIOeCIOMoO0ZeXPNqCmMfTH+OCO3w+eVgohl4bHOMu5J6nkNBdkPV/
QDub25fFIeWJ2wdUoREsGPtC5N/cPnHJ2ZK2mxcAFZFlVYz4UnDT6+St0Zq8nV96
yWSHGQFlQNDbOy16FS+91Ub0mmOPo2XrDVpPcPMP6EM=
`protect END_PROTECTED
