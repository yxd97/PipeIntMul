`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i98OWiI84G1GR7jyeW05wYldlXhwiOsiWIZ4qJ9XxXy7qamrgzdTujkABWq9wSwA
e4XqDtm2qcESfjAV0dQL88iGI4VFkswK7iyMP9rIh1YT550neTAl2oolulNBlL7c
xG12Y60IaHpd/r8sUWK15I351+BG3VJOEbfos42ZqRV1VL/vsjQ2y/Y1AtxvGKL7
u1tVJ5CdYPbGA7n74lE+zKwWs/e6IMs667hqPywmT3JtKRsO5MVl66LaBYCX/IBM
NFnknvb4gPHF2j7e07hyN5jar+DNuo93HiEyMHuUayecYGD2jKZpqsYmmUDvNwBd
K8o7YaeVDHUuKeWVCwMplVsra5Kufw7ZyAMp3FL6WACAO+NpvnG0EwDbCJT3AhWV
2OKpDNzXayzGr2lNm9rID32ZQ8/jbOjUxaP6apFNGES2/4GYoY+ANXsFsffSEoYt
YoCFGQHywdn3eL2i66FSu42SxBwTvkYZZTuCFJ0iHiSRNonhy/d6Gg0gTFcMXsLW
9a28vt9amrPe4Kg9yfEpblGDBuBs5lESztjAtSCIlxAEidJv+g/5RUEMJryV53vR
Toq6lqkmwBgyvUPxhFfGitOCjvQqaxfXP/KANFHwvvcVp6Flaa0D0dZO/G8hkkzG
ZEpETGbuoQxn6oDnUD+mNjxGKbGyrfxdmHwZIlurPYFscNsvVtZ21Fnsc/yXw2EP
/ZKcGhavjoZ4R0K/zqkjAarJ4ogoLiRQP7r/9grCVLbNyMdGffreeadpXZ04hAH9
USJwWbcgFO08imD048efaqvZE/gKXeUk8702jZLARRlvBnzvPn+IMnEWWxA4r6aN
JFvHjPEONTNPYg117qQhlcd8KkguK/v3X+sRNcqvyvdCiS3Te8XvyiCel/KO/jkX
mVWdibguXsJbRYwMMpGBJcg+FX77xzOc96Wn1eXkYO+wR+ZM6uAx7570+Vw8t4vL
t7bRv/RuhTW7ZJ0D4TJrwtLtcq7W3KXeyQYecDAJwhMcNoJb0wSlAx6i+ZTSzxPc
Q1IdXSDa65OJIyEu/1KVL8zwq+kevwLbPYH3oBElPMoyxSQTb2GmHwSmajjcSGWw
+mYx87VqCq5OWQ40sK3Zy7bBPi1h5wa77/PdBSjSl1yug8RFXOtsEiLc7xESrMdu
RIA1tRWoma5h9nTfVtDek/gElKZ5iwUnu/JF2mYsmt4pN9gjgpu6dFMLmdEvjRXx
9uJT5YSajwjPy+gZguWzMUZI7U7lmJ1fY0A6tgwW5/FALO4ou1YmSi7AWQZJ77JY
1xCDYjoQlRPnTjtRETwlxSumWxFDIgylX1rwlx5mp2rvY2k62QXYlbawsM2vuZH9
pE9HvbwTE4IwOcCDVNUqvSYievLLeWiswGhoPZzb70WdS6WJa/yvqDveOxTV5VRi
P927vPAdTngyQF5AtnuK82etAvn3+LHCChsIXUj1egw4RCs6BpM3og8T4p+VxujG
KJZPDIBY1jSw/K0/9P6LALf8Bl9p+3D09C15Ny+7edKqwKYQcS3+l2VsQoEuvw4Z
tZ574oxPkibnXVh6F9aaPobdGN2VRSLiUE9NcCSpnx/A/RsLRnjEgKed9StR6V/m
IP2D2YZ7FLULNvE62QYW/4Z7jAWuPQoIJiU5zMRqSuP5398rCCdffv2OeOWbmX0O
NEaGCxQyKs/V51Nn7wNJQurFw+rCX/iFYGtZ1fGAsXP87GOzA+mXV7bmEBlQy7ys
WZY8w0sMzWkfqQqQzlUMO6J+h7SprB1k6wKrpJFY8kdWjVQgD5uuTk5/1Eusiykq
4nvkfBn9J7erQ01k5b0jePV76Wb5dPCyktfm3wZLAqf2+zxcOpyg8AdytDdUC3JB
j93ZhUGHQ3s12LkOWVxTS+hkVS9JWtNUAsNPtR01dsXvQ/UZn7fopzpOwvX6Fr5y
EA3QqMVEqvKMd8YLLYzQsI+wlg/C0/VY1v10fHfsgUPO6/+811kFHvQFjUR3GP0N
Qq5Oltwe5qYa74Z9OHDFITa4yLRBQpFU+lM5pXXTbcKQGF0Q6ULUL+GAFI+QV27P
tm/EjxosUNTKRAfrGOtA2fNnXfeZC9jivML6PvD7NfbOz7VI0xjYqYn7wmedbs3r
2WXv5/f95GCADm2BXZ3XOPcqyKSpJhaYfgfRs1h1Z8bk+Nqq4U4/6vhSEfxmdtxA
rnc8m1JrGYZixuUBcoz3HE5/tkRVE2vtM6pidVExCkKYBkQ1Cq88Jea8v3evVlu1
3KxrJh+l9LYCQfLyu7Uka8mENrA8F/P4w5No+LKL3lxKLjDOiwGkMQS4pK+DvZ3L
D/51OQ7Q22VFqwHn4gxTUAAuj6TMOUTQsB4OLyHCjj0NOciATcZOjRz30cKMkZl9
2Qoyzn2m7bLhPIwlb5Q7cmconfkovpMkPdkDGjOelkjn66gdqBfce6w98dwE9+Er
a1IkhmXJFTU9jH2BolVIBEBe2FVKfFI9EOu00EKyxl8aMmiNaqD9IaSc0zuP/rTs
lCQDLbBMhFohKDnzyvHgSQ==
`protect END_PROTECTED
