`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0sH8Hwkimkj5VS1blQhGZYn3KnQsPuoAKnIC4XjxOJNSwHaX8lUcJNOF3yDaX4ns
n5CiMMTNySKqqhLxwEBl+WK1YcNR0mo4WdOQfCu1josafcKu/NArxTkxwPqmlW7O
gbWGRAPbJMjJLS22lLlevDAx/n0BBj6ts2X1t+6HErVSDaz1uischUf/TbjBZczt
awJR1xvtWpitD0nyJgJ9WLYP4Zz4CIB3c9K4mRdRXGgdhnxYVp6ScSKtT4YC7MY9
iyixxZ7NcbzBRhlq2PtpvcbK0BhhD17gxEDqpYMAT1Ux5zBNRPyGca2KDY4KrD8L
jzW2c2TofKVEBNK6GxUyuB+vDG8yX4xU9PGAUtLfO0KhIS54O+z5siGD3vSsD5ZR
I86KeuNQEy6ncWUrDmozbzDIa+Z/10yGRgE0MZYGL6qrhOXlBrsL+tZENbj7CbAX
fRBzqc9kOR/xqoIbnCofW6ph/llxbFGqJgNoeE8P9YziBkPthmaIl83ctKWhRQrv
IMcVsu6fzSwxM/3ph79u+eF9JYxkWhldHEmdyDYFjYJJgzTiuz8xjYCeK7JSQ/FS
4Ob6HMqdy9qWIgBe7r5n1dyiw/2+3tRNI/JNqU/Q/xignsMo73CSGIgseqO4V36j
9OiCMGRKNgRGO8VZC7E6pMQFRQhWXgj8xjMGTHb5X1071Q6lvhKmcZwYLGPvzcTE
VioUensvb94OEDLtoQE6H/qudBTEohAqYRssEmSx1C3AoulA1k04XzW/gO54p+a/
a/smZWMmxvRxeBfUsY1AKTxWVEGX4IIP7MD0YtUB7f03iOh/QYj/hYaTqJYQUdbG
x6LmY37qqtdgXMXdnKaYsnvMaP1sV6l0gkHlbTtb/8Km+h9zGFiS6DNGEWAR3NOr
R3Xq4w9STRLT/PkD6stb3MefCcix5WpE8NnIa8tfVtN8lqsItTKOQj2CYfB7Uvzt
vgzjf2wICX4gdBEYb4IWRb7WaVVbaX4SM4UtYu1+0XlJ4KObGYFw4jd0hJZ5T3nK
1aVM7TZzR5UD6SZTUBzGTbs4lUNFkThVgKDMhpy2EUYG12pt87DsdBuyasFV8cou
gr4J/LDlVwK99bBpzQ+0Ik70MGfkpZhg3kOlyXj+BIpNKYc7kTUbHlEuWiVdgIT1
E1MhoISCO1DPoKefi7R16wMmtv1rWGrPJfxxopL4v/C4uBK6Ee98R4pMX+XAGJf1
nBI3DClITGX9A41CdOj08FVo3y8JH5GhbDfGNAaRPhWMaJ2VCmhE9BgPNamCetvr
`protect END_PROTECTED
