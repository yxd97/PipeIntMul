`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fh16oGbmbCJi+IQdX7ZdaI1OouydG4Xv+UCl9bLfrz8/EZyTvRscHmKAjZ2tK9Xi
Z3H/b4Ag6GUoKUhKBUqUdYTwy1582QkJtO9kj9tdU760Otmh5zu2HNqcwSIKXVUR
6Sd7NUqbW71bqw4d2bH/bU3/vLOWP74qaxgecTaQxpqNbriNmgD4RLMxnqiKe4zD
6eJYErr0yZ2sQnjVkS0DDQDT9NU8LPkPLXqcgY+ea2gJK1Cx2OovpA0+3ALlAmh+
uf4CodSjZOFiagiNTVydLUst9X+88X6ui++ZtAgG23cjyn9T2jq0919xJnCZmEyD
BirA8T4W8gkFYUSmvABYq/QoQETS++WiILpM1WitooES3nvilvH9VCILMZp1b22+
xTSFz+YxOOp8gOFDJI2NOg==
`protect END_PROTECTED
