`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lACb1ghP0xal4wRvxng2UsV8rzIEm/aSxQg7AEApWp9GvDZQKUcNdTaKlRVz6Yyo
p2oVivK+eVWzDDV950uu/pd2XDfHX8LiWhvq/jAuonlhdHlBZA7LrzgPEQChQ6jB
agGnvnPawGz6PvSqBx+vZzfIrJEid7kyPQfn41UiJq3JcVT9t0V+1Ijui4HA/lJe
Q/nQWwu/V+2uQHPW5tcsNiGfIKRo1fGX5pyhtgght0kyT4RiuWEAGsgKAvUHdGxP
lCV9iYRZ3gHof3i9jMXo01+zyTkfLhzKLH1/SsZAfubzoM4gUi2xIOz/CSCWPomk
MsxYdi8MWk519XmULqYNacOvkv3BBqjfZYgrIeNc8qHkIFMyqpPA2EjT8UrdJMHX
9Gz+acZ4gsYxBm/i3MiteW3lfEZKwg26vxVJRm4PiiT8Wy49e9scKhfQMVzCQpGB
6n+vhoVh5joGZA9UlANVFr2zl2N82kuM+VJertU5NAlMCWEUcrK8YPHTz4XbthYJ
`protect END_PROTECTED
