`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
baGySzkzVVqpXarNnamFNv2uy4RHIxs24AFGaWx+xCgLdW6NraIZIdZKOZeBUwng
Vjoekal6rmM/wCMTIydDkesyL/fgggu3hgnCJXDmwq++2f0g9vAXdC2/cOQetUM7
+JAeQx453HzI6YEGVLDudVdN77PMlWk9OPD9VIHoEL0Ta9vPaz2KVz1TxXqbfAG/
kvb6O1OjhldFsbLGepko0F5kKvV7/7StyBOe4VatQx6WROphbrvNYHdmnwO4POB1
0yJP8bAFVwkWr5p/7MnhoSc/yiYYA4FH63HTQ1BOap9WOeHesofX6QekW336BZx2
VaU03Jk4q5Bkhh77adqnUlqJ5FSdK4Z7u1sv1+pQM+jz6mpjMCGErgrSYNWJqYBu
0gbD1RoV2wj/o5fapQYhw6wYr8Vebcz3/IQGlGokMmpGxMWIUCr+iwppHJ68GEgB
0C6yg1Jf+mbayqO5RfO3uw==
`protect END_PROTECTED
