`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tZORL9AGIj0FtnwJYXODjEnxZUqG3gbQPKiBS0bggbMVNArNEVhDTOVwYDGRF+px
PFykF6/oACBTNaxPVs0qUqY3kEP5zp100RontKTYmaZd5L9pJkyKmWROKI3qD6tH
b1gE345bLDgMbC1bdtkK4AWUj8UrJdIaNVbqby9cOEEychySrLawf07ViqfGUKHW
uizUJK5/mEHx/Pmwd5CqvOdV7QIhZs13r7qe/h6xfGPgDk8HOs2jOdfNyeQcWMia
AtRp1M7VVdSs+0JQsL7XjyKwgOHv0LEHRIJid8qtvLumk6fyCPExZQeSfm2JOT7B
nLZoYqwZ9PuF55CtEPI+6LZnsAXpJOfuux6yO1t6zq82i0LDyL5OXXg1VbjrQl73
Y8tmes8B+SDklwnSVNP24utS27xfGWvD8UpIzhxBuTcJaDc9B8IwDTMfoO/nKA9n
py0jS/O07BXtNM3CO7f0dFc4lsA+Pn0IXHRhaq/1bjS5w1jOZ0ADjOLLac00x2ry
zTPyGe0jSHUHvnQpXGtOFuBeCSVoFEerb1JznNoj/IYbqOwrHf29DEMsLxNhHzfj
7hx93Ro7s+M246lQQ8jQRQoEoZKlJSyQvFtvIqbX3SgoLyChbe2sKKP4PRpAD620
Kt6tuI3k4PLV+xkzOWNqdA==
`protect END_PROTECTED
