`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWVJbsYF8yDff7VuScn7I3xfBYDeKZT6NmmtwPCk2cJuCqXpBH5VJKz1EGOFLEva
UvjUoMkPXxpDG10g2SSgiF9JBYcUhiMnQ/TOCdIIikbLmk6XMUAFNzgPUl9sxXDL
ZuKh8CCPwXbEshIyrTVF7FPNKz4CqLF440+MARjkJoTRnQZqjvSnWmUKGw6c8Pay
w+2nY1nCeKNFtQKsi0UarafkSC/igwTWrqi1WAYLSapfqbM4CVvoKZUKfoPn/FVU
9YPsqB+ZHW3W+BI8t0x8c6vki4sK5NDVOc59XnT7q2K0bAlUaksGNzGYu/htjRpP
jmmfPixju2qMMolC6bR0whNKROArBQxG83X9hufEDkUErHTP/9CGdigOxPNfybJb
`protect END_PROTECTED
