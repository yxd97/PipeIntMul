`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lWC2nQoHVbcvENM+9loG6fBMHF1n0NM+NePIc0TQ8HFegqlC1L3tjDgfMn287Jhs
IlT3EMB149Nzcjb9vqasd0PRFJmFh6IjCxtUZIYeXRAo9XmAWbbtBGQ033ma7u9z
LzhsLiYRazP6CdHbU6JDPt35xcPUWKtrnPef8TBz/lWDavQ+Ltx/cWReCrdgJvP/
EpZf+7ApC+ePy1GqgEIfBMxPsGWDwMj5neazmWwayDtgUwQppBcySjXDNMPLeJ9a
ZXRSRI3daimFiJHQXc8dKxDE2GWMlfAltPgRTpGBpaV+XgpxkMjxK9RfXYcKrWg0
DvM5VCbiU2MR6rsbT1ftkxZkDJK4wJIyyy9HenjW5mHruL6BfvYejiPMYpO9RWN1
+KNebk4iENt7ENKvSzjVjcRUfHUWifVXB6iSxW1/vuBQUw3Hj+OZ0wPHyWsOOeRX
N8g+iJdKdsVVPJth8qrkjTfBKw4pUbTrNSz/eT2h7jTUPh9A8WaAz9zVl7GNK1R0
QsnfDQ950Qelct+3tnP6g8tSged6q9hlmxVRNiR9Y5n8uiM5DU/Lg67ckIYCqgt2
`protect END_PROTECTED
