`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kX9Nqe2EPREarIhAv9Km63+3KiekgNzOW3d+nAZLuVtR/8zXHyMLWUivjvLJJ0r+
MmBO2wuVNOZznTkMM6F+Mg6BCkeZnyoovAGWIh4LnCCBBVWKJ7WefGxUWvOlj2aI
y0HsZbnU28hZVNJCnj76spYPXACtIyO5DibSAwrLdg9ajAXCrk6t+6fqOvRmnTLr
5eAlmCXGyQ60F1/iOjChfTJvcsejF9+iqOB4+RYkG0gCYl3QsZoPQqtn7W5NYQ1l
ehHJOYkFQu2nPUEm1gasLctjUmWd0BB4TTBrrAVXfTy6Sn3ZBXvzMSIEM9n0wZ7l
Tr+uiFenGYsVwtAS+met5GRtKYW8mxvMIIQZcJ8jFSCv6Cg/y3MLHZnnFJAzBYqr
ShBm6ZmBJmqQoSV2RRlebPCPFi76sLpwHLVUyZboq3dP4XfCUdDRxDPta8VJq8e9
syEh4DUWTIT0LMuo2faSxtHtD+boWCJ+tgNpY2izIBDDnrc/EcfyPXvYt8iSplGG
`protect END_PROTECTED
