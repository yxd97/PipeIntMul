`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+Mg1rNO43fFYH5D6Wxjusz84jgNP/o8jvCzLDIKg5qd4XJjrPXzQvLmZl86ZVpL+
qYdHdg7yuxkosbhhs3oALBu40vzo0woeYxQikf8gN+xsgUv6Mn9joqA3Tgu/l6iS
JMAt6Clw+FGRFuLMNUvdoeRggJq0+EDxqoIreYTw5M5WI2IhcxPpFRe+ecms2vsV
PmNGcYueg9KJMWQp47VY0nZNdhd8lttbbrzi7/+unzz3fW1g8qcV0HLf+Ag6ccHu
zybe96W+QLu/GOCVZREJjD7zhSdylLEds3qpvvuvZ/TggOjC31dytj2pbSOJTSPB
SzctjaKbKJoX18KfCeteoCfmCpNuNW8nSitjvrz1M0OiChVeVt1WNGeiGTJG01yq
XKulNJybGecGE/LZEVrgmQSYiezqfa8/vKIxsXxrFFdVK9Wdun1SBNj03PgCXyP+
Hdeq7rBiafMSIVNMIkHBNgRKtFcldYxmydzmg6YL8gW8huMSlBKYCod48DnjfXJU
Wy/0EAzKWjqiUyOYGQCcnqG7Ima8ARK2cwyZwByrS2eRe+Y/yJEyFnyQ8Xg8o4Px
g6FoFzYc4iYOA5HrYK/hxvSJHEClMqs4E85JMovAu3LiwJtnBYc9xTji/b403K2p
ptgIiAI6t2FUZ03pwHZetjDlpYsyoSXu0z98YJVaETA31kWxpr9+GX1UeSRWwo52
pmcA4gOKLaJVOuzVI6jdxebqIaEb6ALjRYWvUZ+yB1gtul2F3fYV5sKnb7+SdEos
Tj18CRdX68Mx/6FAhwYDn8mXe6W/zXHtV4mRculK3LKq/wwCbTPBp0kmcGkNRHtq
Mime7mNr8OE0WsuhT3qG96kWys8cD2MqeA1ak2KFm+E=
`protect END_PROTECTED
