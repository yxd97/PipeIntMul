`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bXCVr75okwGoDfxGTYhFtq0q8sXtB1hPMmhblaVKeH3Ml33Uuw9a0OyRipvjU+RJ
UsOt0n4eR5+Glz2KXSfJj7Td5THxg0LMbbzeKj2QKSRvr9FhGZ6WYRzyeoauq1lp
7OlHsf++rXkL7GdzTdzrXv7kZimrL5WMx2faKwM1wx77GbrqIJXflfglqVqHC72l
wrCmIqRGBBYyZ7wVGVjGOqdprZouLLCjHHCg9ZYdGVYgLSLF9P3ucRxvYRmc0ZMT
KTq8i8+Z09rZyhg2Z7AQ58uxZYUIitCeYN4n4cFo1Oq52U4Vz48M4dlzYmlp99lm
g1Q6wScVPWq5XjZ6EmyBjypMAgeVLDmmzBAEkU0o3ToM2XLhRCoAe5AaMTE3NgrU
qvFgyLSPrnGh/L/ui6DAof+otAf/72RoTbRv4yFFdrBw5czrkfdx6KGFzdRH18EK
GqwF+T3RhLCdLyazt4KuXa/l/cvWYXl9i0AKC0zmvaNAvrgc4PzpRflUHUKYCcgI
6w9tUUkktSo0nDHIBTvoFkJnZIyvjx1jnaUjXowbY44=
`protect END_PROTECTED
