`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
045+95moyW5nAH/vuCw84M1hkhw4GcwjcPO+/gRv7Vf2oxHlgSIlaby+Z9cR9exx
kVz8nkg4YI4mxeL89aeLKLemRiyq7UNY5GoncavmdmpUMLRMt55Dr++6ypmBVto0
1/Cd5t6Zspjzgi+f6gIZQjK0tPUJnJG/2yg2Mfl+yDGTn0/oLKUIDu54SXJ7NBRX
0i9C8DIWrPkrCCfVG5EyOoNPYV3xp8yuuSQLXAyVjSZjm43OJnTPSq5tyjTTb8fU
84wnlGnzxzJFUGOSDg44qnYZhk0FGMbFGdf2Ekgo/PHKZz9+ZSv9gb5Qi6jHosda
FJstGlfl17q1FM5WceTpKBbjNWJc3rE2emoihg/++W9RJcSt7O0nhOIjKGQg7jq8
MXiSPCK7VqiVIFyr1HDdRnUWKC/URWmFT/GantdrH2G9FT5WFBzsTulXL5UR5YVe
+3m4WxlTGp5OOTrgE9RLgBllOFfz8LLox2SBGycJiNOUtSIpVn63tPPNwTNHt5nI
wiHaTXmSl9ze61wANqRy9xS7WOmnhbLpayU2G8nIMcmFhFBWb/cR0oigjDhyGlgx
XZfuQeKwbmAd2IWAwvy3QC73y0z5hmqqn+FOCyHHJZc4APvHwoe9yH5evyIuCZ1G
`protect END_PROTECTED
