`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Lp2goZfTO1PJ8kN+XeRagtH+H4+70+fXn68fuqsAqDI83qUjJswxqa0Vi7yxspI
9mdLI5kDNDrAFpBrI18sAS/TyPrVhpr+loJlkXF+Q4Kvxyp8KEKwfcSf6//nwN0w
p+pbDxuvwWFC9lQ3a7X+jN0YY36SINZ3XJFPefmVL4Lus6QxdDp2yjMUP6GIoueY
gKaJ3/kP9bbRj4LB6UbF4g+8niXu8hSuuLt3UAqE0P9gYTRjax7QNkW4g9cWWd4O
NoSvYXmyk2XvAz5UuVm8GjgtCM47XtZwG39OLDNinkUdB7197fDHKwHtjwmNtKE7
4mXgPj/jyYWAHHhCzmS+xBuW9fG0BUvHEOxEYc+T0iyaS8e8jRvipJgN+ChZsXT5
ZkLS5ESmhLWMmJZGVZ6NCx6Wd24jNgyTZmisUC9ibbZsW74i2xSBuijkcxfQV82d
BQwNKZKAidWt/gU8b4fOZWRSzvTE3lXkGNl7RAuVojewS+vMMtVSjlg4w8n86/mB
QXU9tw4guh1FgRZupJ+U7SFbWkWoNj+aap/GNgYyDkVhJsgvmR8lOMn5ss1CCFSf
sv22osyKxOzl2d3n4uK9d3is29igHycm+wNzXVx4vzM=
`protect END_PROTECTED
