`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2ZjXQoHvpgaO0k8nMsT89W8wgUc4/50HXOI8OTIo4DaH25e1tTAJh4+1EMOM9+d
/sTUp93jCn4IPSyOogEnFZErWN72ETgMQ7pGqRPpmyYyKyym07AsNwIkec2dbz+i
mbeGWT4t4CX/ip8LTmLmegRTO0W+1TUN97hEKrAtnLdnlqlouoTkXokmBqnfKkH+
Jl2Zt8V02XalaYdZlyJdg+1oQfad09SlttICj7rCOGlFcRdHuoAX0rGne9LUFAfW
j+E3y+5knXbFo42OL9eI+f0IFy2uvb2mpCwOw7Sr2UU=
`protect END_PROTECTED
