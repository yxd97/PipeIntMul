`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UThAP9CcCYV8sD5ocOtWv4P9ZyXo4xiLEzzpzCRe9/36ihLGoSb0R9UlnhAhjWv+
WcP6pd+FI7iDfY9Gg0zyVy3XdEPhSq4Q6WQ/s6q3o0+Wh1oy+gfPyKUC15ZZUmxC
gqT/1sUIfoG/p4xVQl1VOKNtV0/9pcpgUNdo1BnLsuHuOONLf5x3W53q2oiZhH/k
Gawo7jA79bMyFZn+sTIHcbptXYWiSm+rOwlZ/fnBc1GA5VFPMAZMHheG5BUj5mQx
LCSsNzh+xc6Ya6DodkiKaCpiTSMtqoV5XFCUeQTmz29IHt2JpqXH3oiWI6lOWu3U
j/AgKGDVrEjRHi7H1P3ApYocdJ0PJpEY8ZfnCldPg9PnSCfdePYTNdIQ73UUuE2i
kzTn2Vyc8xbHPEwJ6Gu+e8gP1FtjiirCpyGaXncBZ0lZj24KObt7zjatp5VvmLds
3rAF3SAAR8laINEMeYhJ0ly9aJRQidGJzch5a6Az5g7yM/MvLMknf0dBX1wzWA9e
goiPrru2jsQ87yvffUrY+BNykq5S3mwwnqgUdClDvw5kgqzMK4Elum2m9+pZWAj7
dCY2+k8VZPV7Ue1X85/yV2tsQ+v1M8LLi9xfOzoakVOTEZKSZ1xHKtB2jhm5B4Fh
EKO1oWHwN05z3j4QkCpa9AMytXw/+Hec5C+8vcnMd+4pVwgFMPT2nMpe8V+Ytf7H
JwZmnDM4RaBgljeZAo/kYLU9tKOEQcs7/LUAMpXiL5NRjdP74QxSZrrqNVFSftXI
6bLAwQSYEsiSRHX5QnZGdhfHyRPn4VpLmnrBV+3LzK6bnvOehiuhcXBzPpld1w2S
7KgduDSAxMMdCw7Fb6GxzhctO4LFPOtZt2v3Dy6lVcVxKqdRkUPYUhGQ66So37jX
1fH05QavbLlVwivjqSZIi5rSGk53cGHY3EAGg23d1hD00ZmIovpBo9o5raPdYkth
+5K8Nb5YlxfMT98A2oCi2wR3dZzufESxsAZacSjuDeuQ2kHOBSKyH6cnFN98cM9H
my0RqRrOLqXHnOGlFl4OCkkXKKPimSdkPS0qtuVsdG2Y9dXXrORPmE0S97BSWZRa
IaJweEqxx+BLUs+uDzb4ngPtfa2gFTd6+NSIgOqBqMKKre9XISp+QrXmGwja/VV+
k8ECFSWIvxGVxTwsz3iKnxIwujf16SgCgEUHJuyd8ojVOHlq1NMAX0i/UfYLFk22
qjjwUKDV6DFYlDf0RI3hddX2blS0mSs31S3+KvSoBJpQHCBGot/eQCD8mGcSnXEF
Zzw0IwbGz71WWmr5PEv7DF3VRDMUb183N9ZxxfftojHpRrk6pp7tTGt3lgxL5kaH
zbQl8X6gbu1sbG7sJN854AlZEwCfyZdI8ZLVGDFzTrLP49xtxgKM8Uq/kn44NM0B
8K1V5EQgEaPxl2JwzFTdkTCXl+60nX3LmtYtgCfKNW+HhU1y1JHYylRkaFP1lxrh
n+gdO6znS9HR+S5r5nk3y/21I89kpLxs2NedsqZiJWYnticfpVManLRVMMCpB2W6
djWki/zohIk+7LY7Xt0/gmlQVwTENdkzDCJk23QlCaAETiu0+j1o77jowsWavR/J
1t3vBY7+lNOUw1N13ZpArVblKGQKKwpg7YxkuoZUid+vcD/h3MuE6m5FLyjrqlao
OzzYnpKPvWQmsIGuiQuxS8qHDrA228+9DLEpAgqnNccIqTNo2RfJyP6mYxPHHMaP
uX0xlE79tvUkRsA/TtCqffmNcxEJXDkDSUvWPXKtjLSQMYbL0wozupoZDkbB0aY8
Cjy1wj9vyjPWIHqbOFUThN3Rk5fW50spzQBsEfODHL5+mgQ1gVQ5VvR1p5wGuENx
+lx+5rdljy2eTZOYu/RKKLSiZ/KzmNW3ZQyVZ2AzzfsljSK7gDiISlvq3RGcna4b
qUBsmm8J/FYdunCeDAX7yuz3SovY3qupQAqRs1Jxp2flOizo4niHFQqvf9R+Take
Yw1hIpr+9zAlD64s89qu7DenVVmd1yzyCYCs5iK7U+Eq9A0HzyJuk+3/lCtrvMCT
Os0u2N1UR9nYXS5WkuT8UDLEDq6yDoCv78h8YfYYCjVUNGLXgblUKygtm3ZSLPV/
Woc6256bPyG+jCEz5Fh+DC8qkpVF5Ne1+9OFeymGPJikGv/LIljcbo+RT9SDlTpS
bnx8Cyhtn2NuW0ynHgl+QYSNhk/cNqCQQfGfj9mxw1WrqUmggj4Sc4mZ9MLOtNWh
3W9gFNlx4N4UhQoJFFfs92KwpSjE/FIj621t1iiBaPzbY+sldPycBk869o4qJvvq
RYpziWeZm1rw3Afvy1p4vnuc4h/2rG9kR/fZot9GfsEkamiKJdXWCi5JY9803+6H
wagU7PoOPiYQ63CKjCcM49pnLx/QEJOCOtjKeMtRkXPWeePKz+ZHLV3c/la7Vq3n
Mun0p/DflpD7+df+0Rw17v6rwz9BhzrXGxm9X4PdW55N/g/LPnMM0f/1DTV+4lrx
iYCtnkbwMF1znkbCBtb+0yPS0xTlsu120chcnj2aBGCPllc1QSWkYRw+8CUxuCJ6
cN0wlLSqHUowVcBCgX2kj3PEhm/r2AUTHE/jLGgnA9KGhJAla9wEqVlrSznW9MaM
Ta8LhR0k6ljlxztq8oqHiVVGWxScP9UqWX/wX8PehbN4krdt0E7anqXArReuFG6Y
Wee+ydzq9e22rjV3OfuKEusRr0zXQCnhajJ4TOaNU79Ql5m87ve2C6lsJi0sZdX8
QFiOyvRgrkXF6J06TVLPRRgLm8P7UipnmhDblEe7NM1tkDVs2BLRcJ4v0YgPtxiD
zDA4z7askXM7RtN6zJSM/+ktpAFzp4s4000eJVU25BpLX/M/c/jQgJkGks3FNxSW
YvG3X5ESIlClvJj+rEqMHy/ThEWWeJRSPNYJX2wCL81pQ/vB6CRVdLWcwC6r1HL4
nmh5QLO82Gnf65v9fICcJ6Lu+kmtLihIA1y2ex0J9qLRac4rRVAUxfn6ETtMn+4B
/07RES/mQpvhS1h/z+mwgecew1wUrq2yGlnmC5WDyLSSJF2htnAfZUpXo6sW1h+r
iY4Oe7WJsc/+SyoNCa8NFEzYKgNgGftD2pVvGYkv5ng1zfdMcZptbOg8I3Vxt4YX
VIDpoh5KJcX3HKeiS5efCuqlUWqZrRDxJp/hzG9vU08Zfyj5SoJk7m61oczvye6x
QyxZJSF9dghgF7olryjC2K+7RKkOolobvZBVsFw6wEJ+kHDZ4CEaQXBmDn/aFxPT
xHfmDfjTDscWBx4B87hgQSOCAgh86Q6ODZx7SXkHM8whMWitCDzksQcjDMTP/OgN
0/JP9FAd2nqR8EKxfWU1JsoKkAvk5FFevaW0o1IfGy6kjecqXt2CgYPVUhBjvkOR
iRQaceWhZfTAM8o+mb6Wwio6zRHK66q9Perkn5d2y7s9zAVvYLO441uE23IPB6e6
/7npdD1Nfsku9AT/xYUwVHhq3eUZx4VwGh7TSCBzg2zmDpsqeGDnSH2GQTOa94K2
uR1ywhexkgHEVcSIOBkNPHf4N01pNgyKZmi2pKeSXKf+Q1Hio0W6Et4Je4eEfxOP
6jvVnSXNIrekwjJg8P9UHet3PcxBS5HpPy3m6WvMMwaT2r/hNqtAKEt3i5vwAZEz
cNyEk9FWdIiYX6A77l6u6HbxAGfmFgXM3KbaoXPw/GQJ5jhnECdxzRNSyol+WWcG
bPjsu6zhu8fNQkTAp6ftCMyFC5f18zWNXD5yXdnxUmQZ57qHlyCY297bnyhPt2Td
ut/3fFvHsA5ZueqPcnzIUUsnFsKcLelJScc+8ZgsnI3Tt9ck+1Ql9duI6+9fBi8e
JHYzk+mtmrOm+2J4/RCL/cjdO7WxaKOefDp7VjU27td5aCRBv53idFeAfvzXITbK
82PPvnjObhPtYcQcH2ZTQXQAojTg+Y+kX6DKpFtZ3xlW2EAanoIuAccuZ3nd0nfK
FUAxgmyEtXfXR/IJ4rACFn5/RFjx8hmyw709XNseONaYuFcSVtl8o4H6wwB88uts
zdBNL47WBfH2muAludtSjN1vJGnESUDV9ZCMHNsST1sgS/g+KWk7VnBGnF2J1P0R
+i7ppjo6GdK0VjrUOGLsP0i8BZwOxF6Oi+z7dnlvcuphK1nG7YFBsCdTI+ROokvI
x0/MKHcmcWOYs/0KZT4bMh630Xzc4Esmx0obuWvP6T+p+YBb8uQbRP25Vgv7MjeR
/I9KfTBZHoyBch6/Q6GipZSWwsM5L+SNxWvvcXEZ2/vuqlMVIgH8+0wdi5phBq0h
rC29QXJ/V6JGHANvMFEEySmJZxt550MRQ/PuXVylR9YXcEbUt4NeGl0K05vKHdNO
ciAyriyECI3CZ26BlESsxGe/xoB4/qgtcaF0oPhtIEt4prlQv1OsJzfg010+dSGp
oyfWv0ZS/esk9gkuY1006qvfEnJsmCWVH+egE0O9MOqThQzHnNECumqGnzGmRDwm
TiOVmfXDdJdrz4LQRMLnHFwOsiHtSwZ56bk1tP1BgKcjoYROSGjNrMt4yKIM44lU
xobi54qOyhDIy0cejOPWRgAZabkX07eYFyJdZvW/nYaOO+3QWCfnUo3UX6V0JLF+
F2MfvnjD2dfpdsrk9UdXNkc2kn055Kg7CmClpnuIPvaKHJzGtPvHl4QkWhj29Oc3
WIYgyHYRA9w+cUmwDMcnGQ==
`protect END_PROTECTED
