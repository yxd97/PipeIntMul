`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3B9LdFdzkArPjb6TDq8ZHF00AlbSH7YCJcWBmnD+JW7Efert8/cGrqNY8DNoYtsP
O9y8RG91+F9zxypfQRNONAYstfwrSfYSLpWZ+OFcg1VWxtdzS8pZYiFn8QdJK9/L
t7whouc/54TTlaudDQSOU+nz+wlmNKmdSaA3BInTtFpWiPlRMT9g5yZcpqHNMcfd
G13dZv79TZW4rp4rLzITdNMqHFDJ1cRrIiFguVyuYCK05YauK6QrEDwZXeZuf7yj
Nq/SJMdLiqxb/Dgtz4OSkJX9U3Hwm16tt6jrELlgpD1ODkkm5/FhrzTYkBePhdpL
qCtlbIM4qjZRpwPtVqAWGOc7Ufp6ls5qDkuhAAlhohmPjbVF9gFg0KX5JqUdmvnO
mRzTHRFStIBAu1p7887SOQ==
`protect END_PROTECTED
