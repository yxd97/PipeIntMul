`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
By+PH7R0gb+YGUiWKx1H/CPQZWg3KgKUmft4eSANDPEkl+2kgpGsPCueEEo0AiD7
xb4n8F8eOWrwAPxG4hi17cwBX1x+vQLYBQIXN8ZC1USko9D7F/+aUQDHGdPihvOP
W1k8xbvurJ4fZOd46uqPJ0QlDDs8FIAo2rfJB2onVyiKlMos5bS1PVmya5aRDYgK
BNfw/EJAV/JOFLtFndsVUENxZrK3oTcvCmuTxmfmPhk0KTIY/zNinJcjfX/xnbgy
XFSqFXoUIqbmKo8lH6iKDKAzUiDj9tIp0CVg0xe/vXOJ8mS9JXsgF97GAnbD3JHo
X05cfiUMSWje2dkK/zVCbUugZqARohFcFT0z8bvEYoq/yxXv0acjbNw7+cC96JGG
q6xQ8/9JOb3VDAYQXb0nXv3+jgj/PMdzP6/3T76umAFAAR/IFtfcJQUfgPvQoE6t
2mq9b6m+0qeheHtcr/s7QVx3pzdSThBReotvahifRPOFzbnMBio61KHlUSZoYvk1
UL5/gx0o+o4XDbCGjKFpsKjBUOzXCPN4qTYMrqN8xFe21se7lD3kysZqrzUb8baa
53p5EQNHbOi2RMQo7bZtdkCEqQNpYdXefwvu1K2gc7nJHWRPBXNRxHqztgcqlImD
PqCbb1j9YNOLRhueWqaUiHfiuT1bdLLXTacftnNmJX9P04uCGn3gtVsesTxMR+4n
IHscneA778Mly9AGy3/mFet0JAJmtzWVLFbDf11A+/MVdnWJ5nT3uTUHZICI2rcX
GMLzAdTc8YAKZXbHGdavx5+YUAXj5LYx5Ky954RnlhNuPB6ChY0YxS1SPwzxrZj7
esLubpWt1MjXaR+invrjZh/oD33DWMko+WqGZEk/o25HAYVVMTfAMPcWCmqcf38R
dwDBf0/uGthb0AQpa9KVTM6g7vYxUOI6JvX8IEYD3qwyNyRbHbvIoP1riiMHyMWL
j4V/WS+/HzVpj5WcUqJ1tCUZFvBmkpFtMa9ZbiZo3s1YJ5r1iPHJ0ZmPJZyYTgGf
`protect END_PROTECTED
