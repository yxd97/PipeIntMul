`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VqphBTykI0vddtAGd6RpBjf6C00aweuucc1Gju1hqFf6OZtCgfoaP2ZPG0WAlG5b
UIgWm2LRttIdm2ct7APzQbc575tU3Tks0s9xLJeSrlOfxBx13P6KyQjM7Sby4FSy
eH0YflvGBgr8uw7m4Sy9ggc1T6aCtmAgwqqM3Cq8LV4UdmmOlOfdGARPSjozPXh0
YmwcYSxM/rdfiaZqWx1OWXf2hYxscLAnyea0cqg9m+eS4lMF3P9dx001qZz2SIlD
/Gmn3h5qq/reN7ZfOECWzCOP/e2E9Nefs2H9HcvSgXLQhN33Gep5LwS9DcwHdueh
ebXb0Ih0DOpD5YfuJinrYNgfn/l6nPhn1ESnRx/tWhi/iMOGxpR3PAfYF8JOzbla
WLribctVaYXivIk6nMJlp3M0nuOQ0f6ptTi7o6ND/UEMaqCqyF44s78hJZNqPw4A
WM89MNzdCBwY749Qt4PKnclMBvJNHwzEMf2k23YYYX2h74TswuJQvFhQBsSjL6UJ
vgpl/jRAe3mDlzu+uhAPlY19eXBkjym+UcmbCsJO7dTXzAIGv2ZCZRSFFKgrULKf
c1GeCFhl6dl/AwtKuVemp/evoR4pzwMxjNGrjcdCe83dqe00Y4ln6pVBeGHDmc2W
u/sgPnEHmDZx4+wYg63oXemods929uhy4lS0eNpWfwfwf/YvENDGy0ZzW3u9bfNR
piHzW06ubiuTsqCXWNzwCs9bH4SNLkvW5aUTa1hFJlc8FUPDlfZ2Rpd6hVLYdJ6m
i1kXwRXRUQxsaPzTGnAR0GxFEcQoRoidJOCD05tLql7rh3a48ncBEJyiRpfmHQKT
M0gNZY86qtXgLpIsFP7msjtcUPajDrVQv3iDAUkSAEx1vbsos1XensQY1a9T7UKa
FiwmySKjH3UuaviuT9OeliaVS/hqXvO8efRPxw7GYhios5ZwUjFvRO0LtcJEfOol
ci/oZHKf6eQCtuiOhobmN54M1EYo0zmG0g3J5e6H4xOuyMy6pzBPHwKwaYrK4VQR
ViYYt5QJjj3v5eqFpatZaUGxuOl9vnZGHTz4Xy3zQK9g0z6vPu9cRp/cIvYoOQBb
yNrQ7d//PiITQVnzdbF071XPV03hgK4v8j3mrrnH4NsML8pTm52H9Pzw8/m508Ai
rGEkKhjy3O4q//l46atOx6DJnR1T+9vjPk5r0Gr1RJ6RiQasC/p4onVo4MIks4PS
ESn0vzXTgoP72ZD/21VZ5knpFBAI/+wWpuUZitI3WPqbEe1k+zq1yRpjAuV9f5B4
VdaO1h69p8rp6kapUje1rF7XUlM6pYcAiBw6LiVnaH3Ztc/Pz1RU5f4dwYle33kQ
ialxGGQTZfzRLGpZ0e8i0s07ReCPadAd9ZprP9+60+Y5Hli/6gML8l3TU1klW6a4
stxWVpt72NJP/Dkxt/c1MdSxXr1olKZ//0cNq56SCeWrNOl8/kDwUYGmKGCSCJif
jvUAQ90dEqtao1+yS0jxmXG6Cq3qYWndxCVJS+meiCl8w9gzhB8qeUqUIsjUuOM7
YL8pvCIqsJR+/azaHIccDsdmSuaPnpHz1E3s+aqP5a90xzJ7z1Ciw6hJH6HJeauF
dtv4q07YPtdytLTih6fFbtI3KSXc2YmYIs2JAxAq4RqvCa0zq0LQO2qil5ax6UQF
8mYlz3iB52RaueV2Oyb/PqzUzfHg1uDpHpcWJuzhXCKf0n+PkwvtVGRCKHtjqfwh
ezEYB67ORF7lqx3OvKI5cJOJO66fDauS4+sca8HcZnh3rx5Vh2te7SS2R6c+8q+h
HktJvJWoXYskr1nv6AeBUQHrKmBlMDgMlXG50u1Tf39+DqC3IZBK7vFY6ztZVLmY
R3ZUGLXEEtm4velXljH4UIR6/H7HyC/8NTdeFKcHNmZpCHOMwnpTbWqnQ5Pb9pr4
b8j/TMeyosMQW4ZTtRuepCSngoC4sx+rWgL4j2rRU6fTIMrOg8X4Qwn5ZdhXbE8w
rWmkt3/Fq3ndC41WLFSCznUYcpLYw8mukZ0DwSeyR5zdaDqPnD06cZvEUViUd4Qy
OkC/uUBcCLa7ENT4+foNnh5DuY/GrB7A0dH1sU/MG8lyy5e+HdIqepCxQRGU9wUe
Ks4TjEzCQEiESd/ijxyW4qcoK+LntvOT32ldlMGH9BAmIkFVGgsGI575jietdh8x
vsigfN8zPev5JDci4F6jcAfIkrtkXeDaBMXc5uwbpqALKAfZGnZPiWxwEbNWnzfw
oTeFd/1BL4xd7awy5mGnh8SbCNHyjAkByJjkvyvMkf9H/CeY+TIp4jM0DQN+YJ1g
sEHV1lmAfM709lo++DRSf5CpHXg0lZyiAvslBaoh+wHyK1aNLxSBvlT1wM/vdZrY
bcBnqpLhvIjz6d2L0Cn+0ZjRtJrCvXmSDtET1x1t2eK8OG7hJKMArP5zYpFzWk7I
X7czS/Ne8NyHVPjX/+yn0xbO6blmfTuPKulixgXqHEI5FSil9VBmju5+N65W0WbO
v7kLtox35PaWvgJuncGTqyLXo6aR+sipSL+Hob349JJfFP06dikqTcDNR9mpDsHQ
KphuMKGwMa1inX6Kyu+s2rR8buujID8SJXt1/n5KvEZBXg55mCMfYndf4RyPY6yD
pN2eHoE1qd8HTvYDBjHaPid8+sThpBPaXJtWz3tM+8m2qMa2V57mZuu9enk97cFH
K8IjrZSaKZa3Ar/2CIJpbLXxlEUsnakJky4gRUrZ4RYPjYlqXymRLI5E2VzLbSlS
y+LUpoY22msaPioeO+X7YsTh0CA87zP8SVFLRvzKPj6xJRbwwTq0NGjYvpnwuM3X
UfgmhnQeNjxXJcxcYcoWcglCcJqWOETT9LFfXvwjui93f+z8OjfTkRdlKlxWEjbb
0swiq990Ik9hxHF9/Vikte2hD/rphlcrrNCdlnMc4k4LNa/1xn6hWwDO7Rnpe2Ae
GBAhkqXl2964yR6g9OJjOyHwJOKRuG7EOqHlYzVjcHi3qW+DDlCth/HLn/CIKKH+
pcdpFcbo+TS1MiJHAzfoCfWaLKsVp7AFaC1b+JjuqR1uBhxxD700EgpzVfFCoPxo
XvmrLfPAV/ZSCnYDixTeWr/S6UQrIyyKdi295uQY0uAVUF4i71q5Ct/SEwXw6S6J
PTSSE6MdwpWe4g+9eMUyqfV/atRmKCb+GVICsOaFnzDVvlxPX05EdqF1Mp77w9lO
YUe3KlMJLILjrGPvFYZvXqsx/nknJRAR5PskE7GRvkLdm3PmDDBeOuPWgPQqJkKv
UdAjJrFOlsTRal3WJkky2yphV4MMn8ZVil/vhFGcGmovMGXzysNoqVklxakewMvH
R3HaoaFMhoZMoVLM/Et1hQo4ff+3edz7NzGw1I8qIP50YtaapYozWGIwAJ5SB9lx
X9VCcX0wBdaZoLf7fhuJSkLkch6kx8+4BMiUax+foTOtR/kJnFygWa3sQrBOUvjm
zrvHoWo/ssbaB4f+4M1o5EIFHyugRIeaqbJ69cAN1CDjAgkC8hkl5WsCdBKv1i5U
lbgYcg+FIMKs12AL16H6SBegacBjW5tPcc1Zbt6YToczRHF+fpmxXQs23Zjmu1Hq
RZu6y/Xv5LtCj7tgCc8Nc0MiUHcyM0Ksc5v1i5+sCY0CR8JF+34Rwh758V6p2Ris
1zSJc6YbR28BoqSnj175Rhu7DiIwdjmKhLePORYLnD0aekB5kjKt0tTAM84FQW/C
vdjX4cJJWFdAXD/ZT84qAnRWbZ+LoTHn6DvntNIocPUt4WjAnmj3M8XEaqxXbKMd
HNq2RpNKowO9nWPt72WYXl90AanyICibYBZBEuo7h5JnuGxzsafxweuudLV4NAHO
sZzGFNFizr2008gV2zeoB2aDAl7KyzNF8fJf/WQFpoeraW6DX10D5ziHB85ozaqV
JLrdAKflLFqMdy8yee0K7lGB36S6uwnJP6NL7RM8LcjQn476QMS8ubfMlYPWIMwA
eQ/9vxXCJ6AJl0+EBMLROce7gWlcI6Wi1aPV0ck6JpAz9mD74i5Gasa7/U96r3TL
HvDjafPtl3020mvWig7kX2kxbSByUvN4gbIWIxXDfFqyDpneiGsluzUccG82GrKJ
tDByoNpYzI6GlTYLNcanKL69L9LogYvCkQL9tQ/MZoD4JOKL5AETWhKTvB8M4rF+
fDUBosZaH7B/b3MHtECWHdIciOl7ql1Gtt0a1bsqjDq4/lXscdqDLbq7wBZhodXJ
OebITaWP+zV3pnL7z64xqpSct4xYFJiwzY1OHX2GKiwQ8ILS7o2KN6R67qG96/lT
Ar6/i76YBhblIesIothLTzx6AlbtL4dgv9Ol2rtHkF8Lef+XYQanBlQAvmBaeGkh
Hq0Vqf3UE/1HsLeI7DmugIuYe8pB/duynF0RMW6MID05WTEwWPeoFUOiokWafh0P
mrAxRwhpFznZjoJTYL7yiQglSMfPHk8uCwXvfqeKHVwE1sFstQ8VbxLwTxKPmcne
jbR7ClBqBgBsBvpO5TQA3olqHmWZUSzkwhVJcxgd+LjhEOGtGnD7UnSpU2IofRyO
6x8XE/BfQkcXxdOSNre5SMrIDdxyjsHZKBUeAgPOZ9XIkh6fQtqUmG3nBZwKmrY1
peiv/2brqLNBHAegtncG9eMbN51q/rR4v3o/KFNJWIrszdly4V0dnT1xO67SzgQR
8WUfKmIni021KM939tgdzmBqJklLMW7DCCwRggMjNx2FNJRBkOwa9k8Frepf1dM5
iHLXemT2ebrlQX/CZQdmWV9E80tLcc6ABnP6rXYLRhLBIkHdYQXDHp87mW5FyUE/
nZjgju8NssJ5YBt30MD592oa4Cav5sUveCRhq/n1fYmGaMzS5dhBVRsC+98sClXb
XIff3vUtLV1MWKLk27EACz3t175tITKnftf2GGuXsHhMDtiTHZZilD/UmN8hc87o
uQ+z2j6quRBkC+/gKhJXBWFOTmEtSV/nt3wqu7C3ceLly8MCH0oDamhzd5W98kGf
l5TgZIGP4bFquYAKGe6QWLTThSJsILc7f+yvtJlHi0mZ4a/aBBxdE9PNOMUrLaJz
Wbv9/w/qRSX1wtO/vrZ97GjjFfNXym5iXzl2iitBZJWbxtPiyDi/R7rV7baxiFaL
SWrCeGISrq3aa2wCAovnU9mqeiZLtOrSH/SCJos+g0xFsRXx7HcsxgJl5nXOn80F
DnA2fevF6b16s65Na8ljGGm5diEZALgxh6dewfdBxoZycmag4IZDoKigB9Y2Aqlf
9gJ+HZvndNC4h6XpHXqOi2VsCeCs/FrXvmA7Dr9XTo+vCvptJog4Yb7M8niDT1Eq
GBXn2j/fIfSywrGOweZpey1spiMtHlumrJyrwsuEHyoDCDS/sAIMwMgttAviYm4M
FcQuWN6SZv1sB7gFputAqok1KBKw2xGrEc4EFT23PsjunUvcrearL1fnr6jB5AcV
8MQyNo1ZscAalOXH082WRvlItrWCInpjtvngwjWxlVTg6NCa7pwAXCcvqjUDk2uW
+lA2WkjhO98Qst0MiMmdbomvvTiFH1PO69WkAzlQHHEi5tflWWDl83ZDUoQddRgf
wAw1CQnQTiby6S2Xd6adYQTSpi9CccDchsafxxVNMKDlc2mWXgiJ2GhxLLaMnUPu
2zNMDVpYvpFeLcdhhUPTX/HjqIFcgj9lDc6eEAIAiclUilifbVlqiJHsRaszWwi1
LR/UC+v0v0CtwW9TMAPO0gpQB4JA9n79HTMB6H5Zh1R4QA2jcstt64IVirCC/Ywq
xaqOGJLrGV5vr3LNraZaa4JD5KOOSCHSRUVV6AdQRoMMs6FvEPcvsPOB7F9txTb0
mKBrMv3SbxVL0lHW6UzPzdq0sr03Nm+TWVuK6oYdDZcYnQ8ZEgCtBC1nazLon6uW
QWHU+qxCpJws+zu4VumP9FFhfyBNAFqIXtYHHFl3o/sUNkR6eocux/t1OqF0suRP
PdD/WEOltqravzTZo1rOSMVGiLgQIbfXQen+7X0fdMJibrDpmrn20/lGfLYwjvho
+6mfyfcvRO6932qfKRYbjtAHnHogGZDO+OhV7EnuIyxbR9xqaXOVSZZSRuqr/bFO
kqvggtsNp3B86DBMKyH0ivtFx8n9gT5Ci/1Bk7i7Xq/Q/ub1rwE/15PAGVuSbw1C
UCaOoCn86EnmF06dkU63RHioAkdAPme6R09XLAYTizYSqdhDMXLO3Dtx8MNlarMS
EibHnB1EWI/SGtjcidZDwqpGiJLdJ2DN8GeJBfdv0aUo5c4BkXXIeTS8sFxoUPbL
ly0JoYwNcGNJuJNuB/gyqzxTWRP619LXWoRfeL76jzSUQv3gDHfNxvV7+AaceOaR
uyKnadBfCoJSOEoHRoTr0ugpiVij93IOu0JZvwbk3MfnRfY3mvRGtt+nBkkM38Lj
OGjIE8JxuNvRTHYBxcLHGJPWgp+ysoXAsm1AcoKLjy3o5XrmOtT4N4nE8/5GdFfh
AsSN3hL8DZ9cvjuzNJJrWtYMHXGFJ4/i3JRIwrVI+94V+QX0Eyt3/ewz44rEsW4d
HSU0E7QX6np9+qWJ7MN62MDo2vJLZsKcHU12EsMtRtXlG1uB/u/VftmnCw3JHl5g
77awCNNx5I9wrvwY+lk0XAqLTAZCXP9R8D2Q+HE6Fz/EDb4wsJGsLEgoZwEjbudi
UMrYH7G+g0Jxuv5DDri3wvplkQGbir3AYIlW+qRcIaWQYhh7Kju6TuZ1Svy0le3k
aW0Bu2aioQvOOlaFLVMwhDHBvrXhdTLQwNB15d+Y0S9Fue9m4SP2SStv1yJPwyD6
nvQ16VlBRMRqH8C6F/S9OzDrct931xkIva+h35YMj+x7x2mhKpRKWiW5TsAL3YrX
EpZTgsxO4+YClrRnvQn+zg2C9hTf1JhVv1ImfZZXkBCENm2gN+9krWv8FOiV5Y6e
tO0RWHWCZQjlp84640c6dFKOWf/hZPyIQnWkEkKNtZAmlsTvwRwkDDKtNgOu7dle
PusVMfdNaYm9jobpukDG+UA2Iqu0r9t8kVLn0xXJiIS38fTcuMDF9RAJyb1++dza
E7CKtS/qsrIYQ3oohAk6jSj36sRV1G2eZ5DGOKWigKCgKanYwwySY5wCiRAM6LR5
wJzBIDVGXWfBnBZHlrLq3d6L2oW4ELcop6Um2S/yf+XwxmhbctQl/7K3VUmjlZFd
uInuCqiFskJlBInsYVFLNifaRQ76LDV8SVcM1CmNGnqwF8FeI6377j3T7B2l4Bcc
wMEAvIHEz+1b9NkXuj2pQmk4rnt4eTXY0C0+g3FxFG7CakkaCVM3g+uORc/ftdI6
OuAU6hk2SwIvEzDs4x35UvBtz24GW+VT18imP2Gy9TRY+KMZY6A+RDGxW3r4k5XV
R7cm00/HIfuO1B3mTyl8n3qOtT0WvPFT0OCMyZNY3pXS/ckforAPJIBClqBSF+vG
E+sBuUhYUPjY1U2UjmyQ2qLV6sull70fDbWr0yrfWizpDQv1w0vkrjBa+cyXQp/W
1ULn3NOLh33yuecTJlHjBiRr/+6p5Zlxb1xkzzF+6onxyLsQ1UYFUUd9tMjR8NPy
D1CxEmwd6GFnohxXun1Dvov32DvO/KqCTCezQDnsxyIlFHSZJcHCqCb3O0R9AkmI
EYV4srfN2hJCxelHuf8CLu+1vl9XixY/AD7HSDDUr3FIKjyLw0wFIRLuXTha/Hiw
zvXpsX6UDx7K+Is0VivDUibi8C9O5CZMTpeZGJ1BupxJNuwpr4yMhZ8i3tqT3b2e
DCL3Ub6UG3neCch35nqSNlVR6vYia+jKzVUeVx7kaxW+8nkmyX8u6NSNhvcdWvbU
Z6whVJD8gQwK6yvqqkM/XvjYf5A6X1XpDBuJO+eEXHTFqK/KVD6z6fNNLxg42yDG
w+Ham8UXLcDwpgr4Yucgtukg65YyyoiZLi5r/3aaYl6DiGoPptTFKSHfDKWz1pcZ
Ng37wE+nK4e/8v5olsco9ySyypxXWUxfWw7yaJvIlsbX4MIZrqqn4OeJ5f5hxa/b
lC8SkXIPcyizEyefgnbozXZII45qrSkMRHXsLRj5ZDxvvh09U74SSxwzXDqFsmgx
qcFHtSs5vJIkqz51qxE93PMck5qMcG9G7j6X5FbyYpIPGn7BVBMBEaoQqWAmcnBZ
hlHi6PFE2n9uB4snEVTvlptZLu4DNhgVjTxoKM6yo5+g470PDzEW1oVO5Z5oohaT
L8vI7nqAI6LUI8JHUmc0pOpu5qJ5k+8hRsLYSK4tFAL6LUR9dJi7a4lGickXduXB
D4uWNvuZ1EgZ94sgFYhRYS/Q/RW+LFa4JGcXMT03Tp+BdZKeFMEkhUdnhllie7Eh
FiEv9Ew9SQ83AlDxyQ174NlmdYZrvH06ISpzQv7AxHq2Wt/Z7gcU8uwv+Iju0tU+
FSrdlvIpjc5Uym7WK4Xi6hnH6RxzVy/zO/cfwJYB6ktnEp6j1dpm8UwvvF/7Ryqo
Ygo+xEHKFAAteD1pSm2xdwHD6tB1Nx2hFa4VgpYCbtFYNFLpYp+Ysr2L8vnbYUG7
/tlkL4+7+EDg0rT0IY7KeqQmCqXGnrtOT3ezaTvklKvd9mDGfNL8RR/aWAXbcOGw
KrFtP+Lt9kgxlT0ZaN+O2ioyHdlTvkiNo5fQBHaZeHjAWC7p1YtPdHsYfDiD3zAM
qVWP7fbI4A7Wjp0h31Zi6mJBsg/TT9QISf8/gOH9CaOFqmOcI0zmmDd8cw73qx+Z
1yly5xGkvu/CwtWqoWWYNWbF7DRf4n0EELmyPixe8gilJfwu4OMnGkrRYrClY1W4
VwHITXhpEOo0N19QvqjnnKOtK+z3CguH1LGNR7fGMRa/xGb7OL+7ZjUEbQ8xpVON
s9qcIykK4yTQw62I4HlKJU91GhJjup1yaSGaEKHwU6UghC1oWRFum5M3AlGb9ssW
+k+B7sDZLdea9Eh+6JWcno4uJrERvZisDHGwyCQ0MT1QKiOHFugVIjowN+BB0Ori
dT9233ypXQdosoc94kmKLGL3k59UXfxBndtDxRN8oHRUVdGNjgUFITghAz7CSlxz
izHKnoG1i+XLC9jsO/WJGfpa6tpEhi9lHDw1JaD5zpbYpObinekmB/i7TVSKKrKs
Da5Fzx0eMDGfZe7die5efvLkYZKiqaKYYTaU9QLGjWyh+2jbrDY05gFsdbMZxLLo
v2QrYhPQO64E6MI2otOvfzCkexstQAenE+drxYrV8Qf6YinhgxGmTAZm9UEyCUrp
lCmrvizwkwlk490qHDG1uzlCxUINN2DPTH0dN/dvfR/qYQujiV5bW8auyQpHwtW7
fyKqBifN2dKJivItuXHV9rQ/qhze81azUPFSv/eEw/sbJtFYuqxCstMsjyJ7c9vb
OO/0tj3Yz7zK2MPgjENzB0fL38MQqz64kpYxqXs6HRKOPVQ8UnIRLxcz90/bYknZ
0gtRN7V436tpFX91CwdtcdiEU24dFunoKgalRoevXgw2acAZlZNUlUHQ9cTWBI9i
g62HXwGQgzovRyy6gckEvmDiWcpeGwb6zYhLerPbpL5g3pt8KZF39z3T5xUDGKEd
F1UACjxeOPgSnPewAY9AvjsGuIawO7PEUaEYa3mM2E/fyoiM3uH4WdQvM6+QrqFn
PKubs2VyTTdIK3sP1ur695CfQ6dGSOtDc1go9LywTNJbuWD7pwA950942rSS56xt
0T24nFXfDeAdjvVmIDSxEnFSOV/1/NjMo6VRlvUxDlJtasRr9mL8xkMz9wTqWvd4
cgyxGVPJoHAcoU1YXSszrSd6o7HOYYUg7ZhdFOTSZfQkmTMy57RFv1P3LENAjSdj
Ut/2JVHM29P2HIo4XnBXSsbWCpIpYmqa9UxmL6yUr+k7JCEtIwxpbMnmVjYPqKZD
NU5KQasq3pqg8j3oC/+EQ1FCWZ0gSEftY/3J5jb853CZYoE/D1T8RlAZN3xOECyS
tQXMqvQC7c2eL7EGNvzfEhm89Vcn4wxQdgX5jyzxYxxln7efQ+EoJweTnlrBLAuJ
DDHw/7AI6YXPZUI3BrgTAo1/y2HJaEg1ioi8kjZM8hw8nRQWUnRaTU42WZ/4C7nL
CJOvgJZ5wAoYW8U+WgeLeKrru018dMQ6aEn8RGuBGfdt130dAbBZv7qUoTbDaZXa
xvOUS00Yo/pLaFNOxzHVa8CnqWr+5erTeW2JjR9KTKRCnb/iZkpRm+D2QNWYhfb4
olFWTl8lVtfGvtK0Z7ywphim6hy9A+7laztVJy6tNyGPQ7KZE2qMNPnzpQQjaBND
pRr9rRZIy37KvgZua8fEuBlTvndR+nmPmIr7KRCY906C+5nIkMjf//WsdUxmPqie
wNDsRVivbhfspOriLQEpeb6JEXZ4G0Ybb9jhHsZGC4rA05R2m2mwQaQHQZ4E4Nnv
TDtXMZfTUNrVw5jcm1G/XHBSJhQSDirpXf02fIiRUO/9IITs2DsPYaPKlI0ekIsj
VA3uqE12U8bxDpxgrj81rnxy1DtT6jtMIowISRHtEWqjNrUnqR5pkzfo9BJZKXyn
CrvmMqkqaSrQjLdvHnzJXyhgGQtvAksA07zLQbOfJbD2MuTZPSYJZwSzSrdigKvd
M3uNpMc9vZTbCwr7Shnc1gGmfw5DnJ0nnh3HvHn6x2YNRIBrywR/BHpU3CBwGZXw
x0WmD9kgq7Xw4l7083SS3KAgTX+93iZ9AZ4NxOFbBS4f/IWlQTMrCIywiEZgWsqJ
1hLdS4VXqmfDVHjSXIW5UhsIFa1ZnRCd6+uwQSiul93aKJDnHoq9Hc7JVRt7X1Ii
nkLxfCI1AdH0suxzapmnkEEWw5Q0e1ySsQn+YgPxZVB46+vfRdCayf6hIJueP74E
JhmvIljGNR+8Dq5U8shr54zF9npEuuHlmz1bA++o6vqzsETaGNru0X57RnALVrQD
GUDaI/S6h+vFd3ENP9gkQo/gNR6JlcAYcfcSukzfSk8Kl6J1wigpDkjVmih02FLa
flpJzjw+9P9HlzHvtCyY4gaNk/XZBExLflMLIinUcTQNsMHgxRxhdkJjVXiL40KX
kwpXNFzQSh54/vqBFT8vW0RAZUYH+c810vsMd1Wrl55kkUv6E7hoHiFqt5wAHXrK
gAnVhZtQObm+jGEA3ZTcrFCrz/4RppCjmKvWaAVNd/HEigz3B1NWf/suiF5SrnG/
0XCsQznPpGydL8gApoKJmtmcqHbamptoFM0vQZ7kY51OPa0Q5QCJdx0Q6lPbKl2R
TvPCVdUkrj3PKx6IcsVDhO2pOrHPZyKkZPALb2eqiPM7239xBY7qh5YVrNNPPohC
+vI5lpYMwncjpAJdJGzV3PXWiRVTL1+/oIKwvRaT7NAyD+xoaz1nlxNSl6UdOxLG
ZkoW6FNUUEX6eu75IKdX3z4B7WXOXjFpsCAvAfFVrue3ujPqm8MQmJskIKbCX3dr
AhBq5usAyu+SAKT9O/z4zVQWRwcB6GfaDiIkl8Q7HNAGuW+oNL+tJhp6WIm7bGph
mbG+xwnoiNV0j4De9UEODWnAezU3OvDp9Otzdfzgve5sCzJbHOr8y0CPajlJh+vG
DKkSjn+A+vOtQKeKlJtUYYkmzorTa7X9H9mVr6k3tUAmBMLMdt4e8eTmo+bmZa3n
7lUVEGoeCrcef2wnZygeJgWWI3MJm9UtgZDMl3C+YMT7eMjCzmItjPbQfmBCwN9r
4llQGzRLFi/Scun291nIyKdepIPDu8LCKjp/aMsYBtzjf+pfRPerDrhr71VoAQHi
boGwjtFl4CYAVsEOv8T1tl0bUINHloCkN48TIEcdqvipOcfdkapAg7qnOgEufHAp
B9hCE2LaGQ7bvGz3pDp1+Z6qZp7pN89Ijm51ZVUN1ziD+M/0Se49NuQ9qYPewHnK
6IN/Ja40xTr5Xa8Q59nRy8HNMWzlkYbIZhU4YbP/jUl/48m8Wd6U/zlPJKTPmg6H
6I2orCiafrwkeCXQFtKAdjGvjL7JTixQN9li3jBw+RwlCIE6YvuU5UJumSmOlT1z
OXPEDy9z3a4DxLvUsNypEn6616SH/m2EXXKEweKNqTLm0Lg6AWkMigeNCocYBp73
voLBxSX9pQaM/AFN8EGeAWRSwtzI5Dbc36rd8uAUibncKbe/nQoe8bbg7/EJ9pTA
FNOKEOK2WDlMJxu2DeHlwIHXEJOAA0LkUnQt6KcmHQr34U4a69JVXXUhARSEn0EQ
NiVPzRwp1K4uFW1edZ1PY2+O5zNSzq5nIQZUkHxG1DrwXnH9gc+XLe9ilFnKRrhI
ElNpkmQCHzaRUH/auZYnchN4tcfYG6Y7sRMRemfXwxsxiAsL0ALf/j3UbGr6mE8O
zXg24z7WNVHw5D3SKdVtDAsfyLd0Pf11UP+h+dK/xfU5pQ9J/V59KyyOTzEmBbzs
BGAZsMTnYxLs4fUWDjOroWZYwpRQh6mAs6R5vqU8aPfpNmemCvCLsr5HVFDr1K5y
5e5rNPNmRvgSyf/PHNhhLUjGnR0g7HZMseLjr8ft3b3u46f4VhZTOnrY1layhWUQ
TECoJLTRjfJE3Sbi/ODjqcb/JLqvEc9LUYszaLc46fInlReA1veOkvLJ2nr6lJ/K
7d9RfeMbeclyc2qSsUVqTUfbusYzBB64wbbABZhT9WiBz6rDyiVCZSL0VFl/iGOO
E4linqqh35VuWVaRxp2kok/be6HMxLAnnVLeBLfsL5kMUcq3/PN/OhlD4riRtwcB
8HfYDi00YUwWeO6+FxoQk1HQ9UzkVycke3YtK2tth6DvAtnRtp9Gx+QvUX8ZMzAC
jgX1p61EkpGDK9zfzcyQQQfNDhEkkDlMoHA1HzhTEsaEr3nNitM26gvL+OhhF+qP
EADO98dxWGyvTuG7JjevWtYErOL4Y9dg1Z+ZAEEKF67FCyl9eF5WbVJyeDtKqjH1
XoDdz8dUAhdZ7xBt1E2SvZxiGuTcJIrnyJPUeoammivI3slH6VpPmCmerEfd5Pp4
u8GDeEZvbd6J0fYGHbkNMY1X/Zds1xharS4JazYiu5r/lvjI7R7lV/2j5sc4UrIW
rEr0FIKLyX9n4mCeq2zblXmLZ9PXp+mq4Sr+Ou+jXj5zwgUU+2uAzDs/UvVFoomR
ovkRfGO8TCNMS6Ck1QSUB7TAaa/7xacvLfPnIbfcrdgSWzlGOJrXFDuNfLP2/WDD
Bp9tdFX0JTsTP0ykW91escwl+b0bAhnxTO5oZzeW+PPaD1i046e7bT4cwIh5Rf5+
L/h6RzXFPXJZchmcbLc5zsl/e6VuzfuLZkPcDM1FOzrjlz14FggPTfdrxodxezeV
1cGsUIC0Z8vTASmDwCEnOC9FewiwSJToosi5n4Hr7TGuxmUGGbKh507ArHqHfo+r
lPVpQ61KG295meldoFEPnL5pdz3t0GBUl25OzYH4tBM=
`protect END_PROTECTED
