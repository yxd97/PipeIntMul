`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pdfLBZJuSqmRQIyJaD2F55PDsfABl2iLYdzSFeZI9SluQfraTL97deDhqDRLdxiB
TO2pR5YRIGXFGlSRj7kcrgnJKFydRGcJ8tiTpe8IE8Szq3zTICFQ899lwVue/QxH
y5Qf981Zc+RBFN9ttMVWZ2NhgMMBvn8KAS/CDeXZI8LqiHo1GwyJlpbadZzLDpQ/
eu04a+pA0/mid5f3rrrhpJ0Qjk+z/Xkfo0NqVlO7jSFr90vtb8L57opcNIzhWVvG
Mb7S8zoW1khYWOccvv9MDPmnPmlbimDke3616Kdyt9kB+PdzkuMciE6mSxG3nUNU
uiOmPN/eEkMMN6UuAhgc8vuTlBTjurciQDMZkJ0ElM3TqvyRNox7d2ORWHmXdVbK
MLtyirkBEOFJSSzQIvnLUNgtiJsThj1FMSo+aflEqHkjj7xk3TLO9eyU8TGK6tyk
YRHhLic3JMSmPchcQVeoQMjmjpPOf/yBvDg+kQt+NrH8FcvAsd/JllPv7j+9Hic2
5736F/hTzhAtj75hWqLn4RjAw/RQDwb5f2lCcU9MNDHmqeeVOAx243xTQuCFE8mT
qQBIBX73dmwdO4WTrOqW0CjuJ0aeGlTDRq0pjuwlfOC6XF9yjajq5gIcDqSd9ScE
XjZ8Hst57PglNXdrKkR41UBKr6WolnUZf3xqkfXcfGI=
`protect END_PROTECTED
