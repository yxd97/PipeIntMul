`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NDvyI3/y5HxAKANYkUgmmag53gJkw4i8X4OYeEj+0GCZezKtfTa+0B1JAJ0ZHRJN
SFD0syJixK+ErmP0py18uSAarPcPDvfxJo5t7MBoxb8bMxVYYLiOLghXLvGI465p
cyDx4C9hiWX5YmQDnM/tS29qlBa7qxtdqM2D2QSR10pdaGdMbodbZ25NU5Cu0JUB
bz4N0OF7LkX3bIsKXveLckREZXDe4M1BO2i2p343tzKU8ThUNd+vKlPl9bctnEsD
WOgObP11KGSCYgcbW/fsDaZF8ZDM+p/ggJaOHmOF+/xo9XhT+wuTiUoQgX3VwT8D
KibsUxNyWE4TAi3gOHAEOiLGUVUxgto0ZBUhIxZlfJ/7vJXa2FVcJ1M7sqvjvvq9
Vyd1uuWlte31i0qZ80UrVmH9G/x5sBR2slvMcNzS8ULIScif4NXxvbTjTY7KAoJL
6sL3eJLGvJWIxysvyYBzgH6zH3rhdvaoqzjfuEXYU4nD+syUTR/qwcNgyhx/kaAB
9LI5GoWzohW8G8zrHXSRzmzPuJC5Al0m8xJOyofBTTWC0YjS0sdviXNyOZ/TAEdK
A6YYtI8AX3iUq0r5GdaH9SVDwyTAzkuIDHZMBwv1NguvCrtqJo5PvXz6AlbF9jL5
cnRae5XHdsqKe+TU66sdZf9C2JMsa33ylHtCALSqq1Hdjms+mm7n/DicmPF/PJoZ
M7P1xJMTF0XzTXdQ/O5YOG+kI1A2wqgvV81JjmU9m9jKFnh7kixxkdk2Qs4CTog/
G0ZobFyTPEaYwHm4vYVGnk+DkWhGwUwkwpM1XtPMyIoV3iU/Tiv5CP9vRYt/jfat
eoMvjG17/ZzUHlyJKRlttBKgoSJ4R/xJKD7mEI5UzGhicBw/o2l+dPqSf2GXItUY
agxokL/1WADa+BIBdcmfTd9GTsTs/zbYlXq9/aMfHyByUlg0QxGpngkkFA1RhDk5
jvOYVP9hdHYJZ9vgMk89/CfnbweyJpO5/9XEySuE1hM=
`protect END_PROTECTED
