`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qITAE8cFF7bCybkDRR3wkmtPMABVBhxT7xleVqoUVD0sxB41hIZXEdiuvxkkNoWa
OSkROspDSF4fTtLAn/+Q2HmX6eHwyNeeu23MmDl5DFqPSD9Kp9bmVU6/hiKTcGsp
HHPBqJ8yz4A1n40LFLamZyX9WFaGAa8QGRx4XHevhIEbnehj+1mdVgGIIe2v8V2N
43ITU+e8M722kjLIywIIi7FECxFiWCQ14ZorwnRVwnK6oyQJOIqm2EmES0LPrma9
oQ7ovJcR16mvg9iOLlEucTXvKV8nM4aj3i9ILtgsfrz8xSBfsJQBOv1AWiAJSoq7
chIv6EVpm06cqIJiop5uX9+UGeiSfMkvlux7XitRcLbVY+mQXsVbD7eD56DuXAmL
CGVocf5hDQRRiuwjA141XN+AWj2Ra0g/8eVn8p/e/9wy2gjXhEVF93fwv3kg8A6/
vGTiAVdgPMYOg+UC4t8Uiz/FCuNYmJzfO3Wx0MJxU5tLYvJmwB8O9gwq6FLInS56
PADLKpXbPwepogsks8H2BYw85G90RQIvdX6E5HOCoe+RnOGrsFnpXGqwi7o92hFj
3XuUv/BO9HvyGjCXNU63BBYMt8Jw57sh3V1AVB/vhOORSPlGgyZtkAWBK9iG5eoN
E9SqjsTG4W/vAmqRundNOEyuXVrwutcCnS60mFIz37t8MfXCRczwBQReUzG2nE6M
QA6kJaC1XWU93Gxc1cMGBaK69BXtZgXSEnmkBpEejXKmE1d3zk2PrJpjADgKDf4N
vWb3sXDCoVxZN8dpek83Gf2m3ly7BgBNRjmvrTwemFc9eXXf9qiWKAxlaEhlGgs5
k8g3c1DYCMhR6AjJqi36exlJZfCsu6Bu3Htdbvolv2N7AiTttMmBgB96MCujaLcu
Wgsgl5EgkrJhMwjnSsRb/VZEjp+CLvHI+HRjCyEu49sLR0KZfZhXTnjA0xrSurCA
nbUEQ1yEz4VOmFHKiBIBHNDUFBnQGGYU7yqXeJ9MwuV9alzU4k8eSbmW9s+Yfo9m
T0muQFF4t/6yTL+2OZmE56eB70srsothBeLTFFQbW0gYv/nxxpN4k3+lQyDmE+Up
Z3YFdVeTT/sDeei6v6/5XYEkIlOGAYZ1zxqvBmsNPOwc6vjNH/4OZbTR1ud38G9A
kqN4baPCpmfpQz/nCRjfb0IGLl+VDRhlwwy2zdO+XnDKgjMQ5pzdtbaCheY7RzSz
Qh4wkhBncOhy55olMpTZxLsDyOLJ7wWDTb4dD88oGJCF6FH7t0X7KiUm78MC6dEd
VjlboXJuWjVNrBhIYJIX8SQWNoRA1z0d+5fTuvp2ACb8bj3LwsnwfD8P/72g4Oaq
TljT4COjS8qVTYBm35mgOVGDKg3tSN3fDkyaHkzQl5FKCxlwAXk1iIwkGGEiaYWX
kA57UIQvd3ISAAj5TItJi+oLp/e9TqiuZk8tTj+1YbWh9fE44gTp0hnOelujxFxg
pcGR7GF9gyaBN1O0b7jNcp6tf4VA5nNXByCGFFplU0fwRLc9673K1HTEpy2AF4AT
G1bOtPhzrNxb6HYFS/s9gl8jORL3HmPg0xiwU8oyhqlhrG4GrtgMvg/S8Im7siis
8p5bVd6w+cW9HAWv+I92sKcS2UKC0Tx+Rzp0kPWLdG7vGWTf2zNymJ//h4b5ZuLs
PEbFJstC9hmSY/VIAGCCGeAv1OwG4nkishJlN0BzStt81oMyzsGFSIx8ArQpzgsW
tfgnzL1qhqqYAXwyMTjpuTZaNpbO8vwACGguK57byhP50H92ypXD1PpdfaKbPYD7
1a5+4AdAk+0T9f7uMDiNe+spwk02g1HVGJNNZ4eVY9SUk+vfK7Zi9/Tz/bSwMBDY
B5JiFGQ3CD7zSq9KPxhQ3pOsR0kxwdZQzG03fJ6RN4x8c2Z/STqHobb5erdwCwKX
1qfKkT1PG2gpVDuq6zFbDddg+RToWvvsC6Ttjm+JA+i56zEBH8s08dIdKxxUdjpt
fqb5PDuFhEY7e4YZS0DisubaN9GHjiNb883mOW8jDkFCjR2Gxyzrd3+847v9Au1S
8X0tf69eZbigYY0eXnSrgA81nEREc5p1Un8UgFMziRp17ZfRDk9MVhL3jlg+MWLs
1Mp8AyH392ulP+Df0izY2KJwzHt6WrmTc8C/ifWuPOq/uZkIueDBxhoEQ/BaQnO6
J+2zH6Vi3HifXya6qxbpWBCqab1I6b/QQI3OOMRActBLNX7S5BBDtnZS9LYULAjK
kDsR588YFCaZ/EyquD5oaIKpO1IODUWIYiSpobkTinelHdUYYNw7JNGRQlUDHUE4
OmtzdgPLuK9khO9XJxCKGvpipqgaHTydCRKZwKNMJ5NbRncacomwnMEZeADXmbq5
bOc5gPdgf/+G7iQkKc0tlKQHq8N52TQQLI97RbcysOwCiQmY2ttu4Hlch4IFMQAU
Qroa0MMJaN68rjqNxAMYsf6uJPbegBOo8lsgTWJAeVF5JgUqcEOZ1rKwgIxu6sTV
y+fvgcERRSjiLy104N6/euXxeu8jkcbKPDHZKheG15OItNd8nhB8TmpFFh8DMuyA
GmDznAWpBy7c0GNLoNIv7G0YD2Ck7DarFkz5K0JGCxfXGHBLFk5pAFrHOhdTUT06
Wa0r4L3d1NCBgFdtxqKcNb4Tr1elw1KbbaKzi2/8nOsAv1+AhUdgjVo2Crm1qE4P
JxQwxYW2OFsftmvBsZWCSiXl149AvTDMEZh3hIaPYFoc1s7ySidcEHTgPlacP7XP
6ladZpYtAz0JqBOm1O4n7SD1a5vWQ7spkL4aJs0j+0X1MlPVnG+o380kL0vyHnor
nM+vqfcIsC6w2IJi9ahlJjVRMEwUpzVbRWCbj3/JQvgcncl60mhnRVD0c/7SfRvQ
D+UX/g7p2STgN8C9BuJ9uov8ZI6KkwUsd42Uesdiv0Fo9g7MRuhoEhKRxOZQCC2H
Vb+k/q8FTKlkVlbv04Yhv0MSQWQy1+2cB6w13KWleqXDn5SacvOIR7zvFG9F+V4m
mt9KbuvUcaQnzjIBvGe3Rp5LAU3A51awr04tai6wsPYT6i1C3y6xQ21pZqQyNxkt
iGoHZXtCxXYWUUM1WrYHsB4PQ5oSGELesLfP+rU+CMrr7OVJI0nXWhGXwchGLDv7
3J9JRCEXd0S59Oy1sOOWs6lCKDngIg/9Hb35zMA3c2aeBNCF3G8zYM3BabA/2ivb
V9mtE9MtuKRcHWmhPqaYSCh9XvfzzZ1Y/58YAIYGlM/4OifcY7XCJk0N7ptWPiEI
qC5Aipr4sxidyhCmCjn3/uXmY+t/XcTUpgP4/xvFOdjNNlYRqgCbZf+146PpuMoE
ESU8Ju8C5YqCmGe0+hOeaahRDbiiognGKLi4Ov8AUmJmKiL0eFBRjq0l6sDXN89N
+k9P2lNY+E6UTWxB48yxpaFm4Z2R687yGBofs6m/TF3AhAFyMY/nsWf+bb6ZlpbZ
QbZzTUHjy2JE0thajcnnpIXtt/T52F/NA/YCVOtobv7HP69R/qNI5q+QLenZ0xfY
ReiILR0yz3On4HurxiNtMsFKDnLHUdYDV6jUKVbvMxT3qTb2aGnrT221UvzqxKdw
i0PDJv75g5Xqu7oef/8J3+EWW3P685fFJno2HNqY8iwjI263oRujLd4id3sNRJn9
f7uWLO61rtYsNWyYGTHJMnA/gY8Aj2I78J6xmkZ3ArEEvIYqKZaQflQT0nU489KP
xlxiD7BJJK1dHFGePVHVPKlcjmyLIGOc9IXt1vJVx6Fcl9687iR8SxBMOeC9w3TI
yN3YuYMk6QBcX1NebFxGxCGPkPgYzg2OfqoJjSL9EqIAS1kAB5tc0vGXwb4pvpLz
dbA/nNVng927vCWCY9vfVFjKqappvh+6IAIiOkMv4mHrAmLBBt4ZfKh5C0WxQgq3
nxuFyyXdCVt22P69aVKxpj1is5+Vdx0MmzxYASWSNz13sqS/UkZYmS2uhpUwLVbQ
/KlTaQZUwMOc3rndWa4ZFa8X8wHJuoFIW1B594SMldklIPdv/9nIcNYv1KbY5S2h
EJHQ6Ar+pSmEBjXP+JjqEEX6p+g/SxJLrdgCbBWDfpxM7KQpBZEpPmQMfsQU4n8b
+lz/cWQRN54tO6SdxTOnqnaNCeLnefgAiZyYgk/MCb0/HL9vO3SnRYSUXejWWXzU
vZKojRS3n5VKkcBn4PKSnAkNPUl8YpH0VcZangerb3z6qwtFBmLqflSWnIfRY6Nc
MOpQQPkIE+Vkl/7ig+5alD3ImFLf62/4kYWNhhQkSXVZ2obn5wGnzdtu7j7lPoqa
nQ4yhUFntgtaBa2WemPV9ftBsMUCENjY0wmL4LFhjxO+uuD4YhD8F9RPW9fk1vuH
B4uBALHc/xtY38GhqdE5ePZl0uYG/lvELJ6JRe62ncu9di/9qNWk5CLwhUDwOi0n
88oe2/IswDR2IZkRR2aXbiFatcZRtin7xlTnZ47gAwWwIHd86/sAYY7Ld+5HZwZg
7fPJUdX5z908zgQ7sXt5jcH17G5BS6bZtjA1GnjiDnUWWX88ipiroRW3HiS0h30U
Q1MoIZEgz+9PTwyK1jJSJohDG6fWLaO0+znXFM7CNiSmRJC2Pz3kcMceft1aLRBV
kPDkJ1VOWU73p80PavjG2hmsqZ2jAQ2ni/fbRGBRrbafbtEUZ7TsxVe2VUHnPzmV
+vvdh6MPkj9C3VtkwizcOcaiCqp1ZX1Ta0LE66DGHMjdgjVH58oS9TH0LGHZZGGA
j7pNXJKFeTz6fAvjY38HWuqsrcaAILG/zfBIYON/Lwf/51OBNFADRiwRcMOFMW59
ZnZWpGjCuKz+NmTqYfTgoVY1T0YzilNp94dcz+l5yzG2r2hk5wRzv0uAyFi6PCOP
haY6TeOHZ5YMFWr4eoqOQwDuXv3TTOAA9fvx7qKbvyVhJVJFLt0iqRjYeAbg7qj2
x4BJDGxCiCFPQDDbgrxuJqdEKFsia5A1y8GW2VdcIZaDJRDG83Uo993yrmcff8ac
1GrWPS2y5VW9z7umTu4P1fTbDjNwvRyQ/OeBryIbUeyX1OiNSjOrJMSRzMztT7Ec
ymNqncUs4UQUBV5o26pqtijNkHAU6F4CqQcuwjYS/3iB5DYME2fPXokihHrR/Xuc
w7M2Dj7F0lxwip6VYY1T7xIU6ICiGxlrtCgVLVUNuX6FBPafgNltTPac0gwu1I45
LYQZDwkSYTMG+TTbFSHrHKXJjo3+THuur+xVsgrJfdkkJrwXzGi0FxMlCjUugXMy
8stodJC3umqzxOZq54j7kP+hbabwKWNUuk/VATI6o5O7ZW2v9GFaAFKnEaqmGAAJ
8esSH/vVndja757iAO3El19tAPylinj0jh9nhOUFwjeWDIrCpnKpcBUNpscvOY34
e18Z5t43KNX9nEYpY7NkUO2B6qxIW9T+8rBJ5QW8y1W+3KanWaFCLanGsRb/K6n2
izQ37e/DONVGx65uZbQNHi2W30Lb1DbariOc62ODczo0sNHK1oly6yz++uH+3QyE
CnbrQjb70LkUwXbHcRKeX2OoyF++JPqn5oWZbJ5KwZysZ3H9ekyHCYh3SEkAz+1Y
EATC/JgxftvUbMcEtO6K7dS1vZzgE4XC8OCi8dO0VJn2WxxjjF6o+AlF73ytHEsI
QVxyanREnAotwsr3YKANI+2l93T5zViXuLRixEHc5YBBXP90zClYi6nheLeWQhCl
kZW0qTXqNwfaHNJF3UlIwZn47e/W+r3PcTV49BnSAQs+QJ+DMXs2R34zPw2iBYv4
JjpyKOhWOO9sNDLHayg8HI2ez7A2r10PqOavvRX4PToMum5DNgEZg5VdY1REMn3L
hEVF9KOpL/8rGwil30L389vSJOYM/qktdCOHMzbO5zHHil9u5f5YdY7l4LFVkMn8
fOyUEsKpLMxDHk+EeeRmXrzaGCpSHB17dtZfW3mJRhTfEgEEv3Hbo1+pWFZ1F0Bc
X8bUsv4DzemlkQ60dOoAGiMVhaOJyneovGskBlzCqEPoenOqFlmTvx19UIE8tjMV
pjtXEXDRP9OpFa0HjE+63dQN+zRoY8JgfsDrM5OMBik7/nOYPqK44jGOewLQ19Rp
zjatD33jU2JjB5sdP2FWppWrtEGsHIN8qaAX/EfuyJ7iuf7Cf1XM22GTP0DbsW2p
vrR8is3WCSW6m6ZkKr9tS3MaQ7cmCc6qpKyhJhBPNIg9b8MtroVowbhRBlH3nhnR
TiKpMEB5heJWLQC4xUYiLm75fX5FNJPyaOYZpro2D2URmhGwM68pzLM2xJ8yO54y
CUM8R9m+OdYpeo0Tew3U+a9YRYMj7ElV/t+3QRZhRMwLL+oDfKoomU2FSFwVRwWj
5V6MXwT6Zq2tuXmZ+EqHkSW/bjBYupEADG2FZdQ0PQmOWDHgDEPJu3gcGHawJ+Ys
RQjfmz7Xsd6NooVdj57t9XNWJ0o+1hmje3jGSxuQii1E8Whew8njGb3BCegRq097
T/eOyy3emdYiR7netMLr2PzbSd8Efh68aqV8fIdtF/G3Y8jNdGKSFEqoi6yyZ/vX
gNwxlW4pX7zaNtgp7aFySL8fJ7PP9FulJRVlOG95bD66FbHPtgXpQHgwAv5OCwh6
OQA6a1vjfzW2xEL1AVGLf1qTg/dnyh6jJ8XLPykzP/iilJHkA8zDDhLhBVc4udQo
CElAEMQjyM3MsHikv+YhlN0OPj2gnoC7stiMQwHjkHnmM8aBGAuBSZfOqfQd5X83
wfbgIYzhW/630R4aTKLCrXMsbB6Fmh3DlPuYDyOJxvLUVmfJ5VRKapt8L9e1iufK
zjqnnoN5e01uF42GP8Wx7737jjQB865JJ0RrO0xtz8GSJFiYoWQgu1XQlfSamgBZ
amirCwydCQgc42sBA8deaEBpaLIX8qGY72slWp+nRlsjfrsB20YrQCsnMyrQKrs5
o0j967eyIVIKuyuKQnfLtg97OpJ4npaYJBpU3S3WkRHexdQ4Cv0h2B2LHAJ+fHIR
pOMeLlH8juFqpZSutoA6XLRZpFVzmmVnGlo9akYiaBhBbQwIulmiZEhrGiP9qDgL
QaziW3vw67TIOiinllC69cq2PBqVZuwePucgjdHhMhUS3WcHd7BNMUWjy05hGOcj
RRRMEPNAkmX8FS7yLg7kq6bKxLL9Lv1vo+54yCj/hZOkv+x/rSOi75Hf5VlExY7A
KR0rCPmnqcmctNgAG0s+GntZNTbOlxtq7TgqQybNu54jQ+7MdsxfRhBjL6l9QpY+
dyF4V/V7CbMGwn9WBqhX5ems+mdaEuStwJgzradBFFQhvr3+38gqlEHv/IyrIfDg
sI8Ws79OW0EWbtkCmJptIYBPj9TIc33zbtkBZzRZ7TbWYrj+26F/xrWO9Ra62xF+
0153fpjVvNcxYqMsoSGTm354RSf+6V9K0QTitwJt+O6jrxATy/JTx+GysW2yQETR
cR7Yq2e+a66m1PjW3pgt0qBZATZ7x//Wz1BU0TCeDnRZD3pBazE+kcRPZOG83ZDa
D2IpzrPFE8P6+T46GdaDkmYQwlcbTiG1nzcCLgy+OvtGiaMSKxEWSNdywI5npcXO
rsmY/vcQOioZVfsMpvhoNw2ejgIfOoDlcYrfVhWOAL+2jdhM1FkGNkPIRhV0xYme
ig/5Jwd2gj/nkD07Ra8XP/4+aAqv490kl/cAoqnyR9Xq9i5J6HlHoqktqLIgB5N4
r3SKuNWBUz6PJyIbVaEOORBCRyuPG9XCcZQgomFCWQFO0HJ7d+MXh/Pa9X3ZeUJV
+H8exL0D4Ff23gh5Wjj9RfZeaHkBjEHfhSuqpiBv9xjMG1aHDbHCJ+o5qIUDmBn2
CE+AJedes+wYAb0XZJZ0wM8Jk6CACfg0M48vf2Jfr58VWWeBz/AR5xwcVebmgRu6
JQnT5KoePDFPEgb+PIEX9KbV0QiKzOdIiPa4nd6ziiNcKoAO8eA/vuz89C0wve6d
5lEDI7dZjX2XhvjlUXnBqoz5/1TjyhPipSBTKnIkcSMfK01e+x8datjkTiDj62v+
ewCGij2DotuzUl5bxyKydbQ0DD7mT9eeYX+r3mbUW9vsrNhmbXzxkv3qIbGDepTZ
yyG0SXmXpIhhCl1AjJAXeO9dDQOPcGHG8ifrM3Llsg7V7FieWIwoIW0nyDTO4ssm
e3MCgAUsPE/6et1nDYvHymHWbH4oDr/ofdNtFvo66Xb99uN7PFWdD7+ACihFesNs
XYhcPIV8v27WkIHwrSIArkFnKIk25UH1TFsgsfH/K1IHbhGM6qU1Zh55uXj2NBEr
tGw76wUZYrQ40q42HXLPzGdRnjg5hE613tf5D68xq/JQwA7ROtWa1lWplW9eus2E
cGWKhF1sRADYsRnSdjmpRpbl6p0fFtFVJjzlXvuOg+IsdI1XkzQp7m3JMKpGOhRj
bat5pVATWEpSnZVR+EeaokeSaOSJy/42QhAD3TBFQw2OREOFkzjz0gXdcXcdaMwJ
wJxwt77vyw9x8z3HattqeI8aChMHDaGIZ0+FQZwCY/uPv3mw0olWz7ida1y6z8Uk
7nKZI58EhZboU4Hf4iUV7dkalB/xqZbc+zI4b1pCRYD66Rgdg9w8Rq++44w7edKU
fnRYJg08OgUp9YM3HADaKG0gSs+IJbKTHzOkXLAh6b6JI1UcyVoBbQIwbbsXCUYS
CCPH9tVt+YTCQ3EAH9brItSQdgf2avIYdLjgmbXxsUChQrAqqEJ2OvD+nikYltJl
u0Pf80zlSkN3N0kes6uzATdGw++lb5q67u0z7N1Vg/Q34cvfj7eogzRiRXk8NGlN
2vFtHeKrfE/JXh5peikic/XM3yIYk9/iH5rXi4+3K4bNVyc9HCYNugJv48vts2Uq
/HiwnwUEFli7jsons0po1+6ym8QaJQIlhoSvLsjc/u8C3GyKisUond8EkL3o9E9B
G/WwiPMoq++GJ890pQBihIxea/wf+crqWZFtK4k4VjSrhgZVjJPhtGgV3EtWqDRc
qcy7DpYlPFNhHyefB/ZCKOUnroBsJ/hY1cfcHY9Jbl0fkpfIaxZYF4/2SXWLQYK5
AiX8e0UT7N2WkmDtXeQd1KltvQVrwarsjGpKSTfNbr6P9AAVj2KZzibWlQKXknWx
zb2LfEjlscPTRG897b+LK5ra5s4j1M2rw4F20kQ/BNGEphhowb0iosYoIe4hzRLh
OGD/Dkcbb+YUs8Oj8/9xE8YXHdgQIuLaHC9gznv9/tdM85eAsz8h67j5blD/6a4R
Gl6t5q0fFWPOyFE0X+q1est1/Qr6RDvN3qBCgepYrg2NCIL7zb7DmH8XvNM1Y4Cj
/D3vRSS8eZWW0jfLLkD7P+5/XSLSKCPfky56YDSWetbPiVFL5dBFb3GeGSRX+2A1
NBr9TD8gkyfDkitIOQ++Mrt7POU5HaA9XNrSBkUvWBxthavKg0pc7W7SDtmXE9Kk
jtHBvJBjEGwcszIaXB1dCbIeINK9xmfNJ9z26A518TZD6f7sUrJ983lLUBv3OXXG
B3LxKiMYhMdwjw088w35jrtRkkGnRuswGF2VXQop+Y/pCKUNJ/nisoRuQkIol2CN
5g/zyWBxt0OM64PO+x3pv2yrA1FPBuMJ0nGxoNZdtZs5MEKh1Tl3Nv5h6EA22wC9
Sn9PnWqo1BbxNx7wmtNcDzK33VWyfrNcFzv9j/FZzr5gQwqH2XK/aItyZfCJkd8g
NbMeI7kfUVuzI61LKr3nzguS6CXSj8O0xj6qPxNoZc5DvHCXpSLqz/2DN47pUcRp
yMZqELYNOrv8KULnGlVZpBnpPSBhvK8CMIKklQZi3LObpWhWIH30TDanIP2T6AAS
SD6XbMDNK2rCcB1JzMw73FWbF5BSmw1P4jiYkUHtJLXVuQ77/IjErq4fFk40aRdV
0l5uZzvvUTfWj9RlrH5944LBI7PMwL5DFWXp9nzz6pl14qGt5InWoVfB+lzhZe6Q
FSg3ulqKuNYFChD0yKlDsg55HLG/ooVaP8yMc7G5+0OSDXQ4J4phyXmJtR2VuwAL
jkcHy8UPwkkGyfnHzJjIFuKxMzU+xKKfrkMOHpv9Vi8viLWyjLLLaWuoP4VyVchg
6mabL1Gu67P7Sl3DdInyOxZmxmyCdCrkTEiR8rcEmbnGrnmzETNQadvYe2s34Msm
gvfxIRaj4QbH/GAaOTSCDAknI0tCuhr2opVRr/d0+0ZhcXPc6FdEWHQgvhvDDxBH
oY4HutCuNaTkd0GsG5jQbMlrzrab+bFISgRWnahS6Ejy+xXwIGVHYBWYvnGgH+I8
JkyWei2uqZmtJK1DNmDJz5wiaq/AoKu2UOTUYzroAM+1C8RnEV9kc+fPM+hKrirB
0gHa0fUGyIjRwQTCKVGQWqUjfjeElu6/0yocjo8P+78vHWb9UdXPzBvwvnzP4hPk
oIEotybL/qNtATi0QtIXmeud62mtpYSe/UNKUq2wZTPZ4sHk2j0NC6M3Rx7M3/hk
LMdZGGe0t/fWI9jeqSxNSLS83zVlDk24FUMjW8+LNr/ePiVnz7YjzDjp5TTm7lvy
XoNLTpqgxs/zArxZeq25pT5geXfxgiXuVqUgjZpcTPw+nWyr7CNxg298XN7J7uON
Kx9SwoM6rzn7hoSd0H1wD3St6z2lccJEQB5Jo/GcC0PgGgc7Fz90n1FmSbN9xK6y
smJAko1DHVmZSytOmmjTx1V8GQPCllw+r8uuKHGc1JbSHfK/hqcgyikwAy+M6xNT
zzHrJly9LOq2slEAZmxdLdj/omUV7X9emFiD+Z8c3nhiQr8joQGMmiqtWGUW0GrJ
DhBv3gb0OewNJdDIUknNN8+yLZVW58+iOJrcoBSXKmDrUsdf4wckV3rkAw7qtxQM
Mn/Znj4+B8j6WzaFsccSrQ8xHxMF8/PR5tl3X/xPKs1oPzKeM2Kkz6pG53GYV/Cr
FrFsPqfFm2HNE4ql5lkfClzF1bLKSkZl6reDd/idfJDuFMEPMMSeS5QTk6qFTl+c
uIIRBRJ1n1q71s9Lbzh1bLaZ/oJhhDMQlB7JM+hXo9Q4l2j/ynoqWWhJ6cgLirQg
Fiq3Z9sh0jvVEyK4aIWA09QjrZ3IfskF7T/mDFUJ5IjqkZXubYk0Vo7PIw0APrHn
1gSfWdILsFGuCWj3Twu9bQUyvz3hCasC5wEGga4SVuXKQ4QkH23X0FbbEA6nhGp5
B2DpLH52L4LGkt+J8OAewydrhywB7mnJlBT7LPjaZtw254UBe2eZ/szNt+01wDyh
ogoJ/Lu4b/DmW27bKxNiMnoJL0jVC4849RmUsQDB0UTbm/YX5sfGcymwLtGF45DA
wKUIkQWUZWwhXBP/01yUhMynYeS3H8fiMu3itPL7Qm+5jHfvV0IUlxTS4a4H/neF
Hc5EBHw2j/KvvCelAifm/t3A5zh3+gMquNtomEiwdqrorCvioQykZIYDYWL3GxLb
hv1RH2J4hFEidm6+DMQs2E5SFv/6hCnAXRMOlkYSQb081mItoOsWzen9ih9BIhSX
oZeeg5DVFFKAWJ1SitBGtb+qK/PEE/x9cBMQxF5082S/8mc/eOdbkfwf7B4X9Vgn
td71Dzi4JDx0Mm9VEjujTlI6c4PjMO7cE8prknmCZNYCxTlCc/YTsr0PL9OMFMSu
BMfZL4je+cNf5Ab8kzzBkse2Ed7q6gFvDkObDECE098=
`protect END_PROTECTED
