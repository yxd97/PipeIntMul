`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDlhhPdJf0g4h0qXgtpDqLHng0cyJE5V6Si4KAiNhf9r3TQ432YamSLc+5P8UBo5
hRn0porHwaBjGiKjZeNbflWh0KAnJoWx3dYnAm5LFlkOtatTsv0PQhFn3/bHaWCc
lkJ7xo0uuLcNIqwTxx4bnIxHVdt9x6BiDGX0TBzPDdK8/x1dTzIEDmFohxYkSF5S
LI8D+qt9qjZlu+ZZ2onHOlSseT3zUpHNZ2F64Co9Hef9FrOFkCx9fBjJ2+BsRGMb
14N9dTMsm/0xnZ/nZhuPJiXOiQJffXY6y3gGqoxK41xDYnKaTFCp2imbz0NhLD9/
fsWMfTkWsQfmnniW7OauExLoHS+7ZVzG5KRvOgGt/O7o5tS90Ynu3XXtfJOoFhnu
0idPe5cYRHd9NI0dhv50esLCI/HHz4z1TdPhG5LUAKlvaIHdLM1kOH+YL+6ylUDc
owkl6yrHz+vMb1dUDo0aj7Dn6s5JRy6W2UquEUjHA8lD5mbiWHC/joNOhPl7iSjS
aef+HIDg4IM8Afhptr0DVIHpFHATDXq6fSPVEKw8IuksrEkfc+KtPpKZqpB9CnUe
ZaQqXjJEEO+Ta4Us8WY6LKjp1CMVf1R9zJDlpb/XV3gibMpgJzX73SerGB4DK4FX
H0YJJdBQoEww7NaCtSyPTN9Q7iVgK7AFoaMQjwsK2ojaXCMh6QPsIOKsFfQHAagn
PCETqLZsBuDQfalaXiuzqqXiBI0aeJVZRu43GB+jRGKHWgXPeMgnzEkAt9JVSBLJ
WModOQ5NcAbtwSIkxsPWWQ==
`protect END_PROTECTED
