`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AC/vgZhXnNPoaL5OeHKyfSNe3sODpFvQthYkcbqh4ro1SXockn4SeRFbEz8tI9JN
r9m6CjQpmMoKYISeAb4PVX4Szj6q3V6NG22pLZLcrNGBYIRzw/nlRB9AIu7xTTCx
dzXY8GcQKbR8kmhvhw+zQqMDi96rViU4CWFBX3a1l0e6cw8P7uro5gJQeoNMAvj7
xBM1AHvNw3y0M5907N3yVxXzQFnO0SatxFdPu4ga/TrhVruykExJms67FhO9lHMD
Yqh/vi2S9Ti3sXn/J7xxig==
`protect END_PROTECTED
