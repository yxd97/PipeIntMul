`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qfCRetN3eXDNgmyk+XefbufpG+xqCOBlyFjOWSllSg9sSVjEuBDDxug2uAOolByk
LtUq7PAC6ddnw/dv4TIiP5VV4zrRINLpUz+SI3/WMHb9kPmSDJyV6ALmRYjC4I1X
mGjQWNvxw1emdU5kFfkqxZu/k4NGLUrhh0E/rkOriAqDRFglyIMJJrqcXlnLOclU
2Wcf9PKi2ai2uTrwdwcIdBqffb/neStI8jyUtTF/Ideiyu/kRX3aeFRJbVCTyAwa
SLpPSRoZSMQCOsC2prfuwaTSg3DIA+0v+EXZ4gF3YjzMH19ntqZdXcHya2UN1J6F
wuW9aj25VbWyJ2PybrieGaKUgDfUpzw8rdv9b96ytXzRDK2GKcn3zflKV0H8mdUu
aG0Z1fsTqPAjtgSxExMjyr2v1QFEiUmGCMs8jIRBDz79KMJxlYjx04tTy0Ei3WVd
tinNctb9fwqZR+eVU0q36CGb+ggdbYMZ6Rt4uzxeE2yIQ1qvSxxb4ysBBLOHuX7j
83J3uVufi08R6u/lqwLThpTVOrCz4/NOM14Doyw4LiOnNLs9U00hPkmMIUrBI/KX
RqlyG65WUW3PHDolvS5fTqJgX50/zzZ8Y/4m79bcaUX0pWRWVufbnUUPa7Yb2Yfh
4zpUvHDQzc+CSFVANc2ZVIzgVja765aTx0Mu89y/gQ4evzdcR8SxXSzhu4c6P4nn
Zoq1rqBmojr86omzmrfIhhm4wzqY9gvY4ro6/XFDAy8h23xR4VNUXhlvZsBnUAfT
2HfP2kWJFHb2wVirfPWUi302Kr6E2XXVBwSv5NUKf+gPftF21OSA6rUcXy3kZIpg
r0dgV9edcbX6atRm51rH4lW3AG/Za3utxzM1GPwah/7TF6wTm8JR7S4aY/t4IJGC
VlqinMHx/HaVNxqzE9D0r3Lc+3BeBZSaJg9r+yI770QUTz9XJESUGzxAWPAL1Gp8
WTj4bievzM58IZhZjsWd6ivAw23acvp+JbDU59WsR3Fox3k7Yq66q9xUh/AZu0B+
JhDMO7cIV47L0AhdfgSR4OQCRj51pwSdrgq2e5viZSRhM3q4F2ymedlVeYPdVBIz
1yhvJRQiJiir0wXrhjMabLgygiLk6d4Iee0oRb2wNok0CHvCN8NJPsoZIZ/grSgc
gOt2+ISqQ60+Yp01+UU/6FKze2X0NVqPRlN4jUN0EjNg50IAQvyEdHhcE11xhsXA
Jn8mOSgJEU8KBqtFJXYvs76F/FHtyYjjuivdvSdFJDGhWGxg5cWgaN9AvRiRdd5a
HHHFuGwBG9dwktkRwIh2U148MkZUe73a66LpbNsqyT9fjKK8JtUth7e7EI4yDPaP
5s777VRQRYxnxxLKv4enVri5eBC8eOeTJXgcq9Kf5eI4OAKeAQamdmeyEM4q1hpa
2sHfZ5PAASshjetjRiy+2vWNGfPtTHQ+Br8aIKmDgiaewjPsfTrCPa8lMHF63gxj
wiT+qicgMVfHfL7RLq8MxNGmOoMb12y6yPZoH6GH0QAd4/jPwvXjjffbzx1YAi2e
Oi0spQ1pWix0uG1I9V52eVylUoGVrHYNeFa+PXyx7HfnaeQm7uAfTwf1uVFb+H1A
ZUveFRIJtXm3fZtEVpK8VZ7d+7IyTsGoguXuSO/pJFYRO9Jo4/BSnNUhWzRZNI0T
1YcgZjUgx4HePeAzXYHayR6YAp7PKR1qigzDEtp0QKLVPPBjxxZ2fCv7kP2ucoC1
xTkVe+p+MWOfTcvLpqjqHd18RSBrjKq1FgHzP0pYZM0lGC+vvuA5RRQSM+UITrre
5C+uPBSZRGNEeH5oQ7bo+fAj8XxpdbhchfVovUxqANALuZJY98yTwYm7FFJy93FN
Ydv4KLbs4GYWjFvsS/HdmnWAKJqsKLqX8rzqDw0SAlEOHULAh1z9p7FHrqmyy0T4
B9QPT5Yy9WGzflKkjDTFuytUMwtFEhrLRvUBlyq2x4CjJ0fY7guOfsSvUhPSWznv
/FWclsqnb/sEy84IeB3+KfFitifRRF/YW80h8nb4Ry+c1r/BH1cTfiTzm/406TBU
USZHKL1z+pzjucpRDvCCggx/inyGMql7Fp8TNsveM9mPspvhNR1ApH09V0ZZEdO7
fRkpEcyRxVesaPS1kpHZa5NRx6Tbgyw4CFsmaVOzhCuaOqq48PuYARh575bxzlJ7
VdnOENr41ArnJIMDuhWcw2ddztRouz8pNyLE2q5nu4I98iw39E6TYAry/Mrm+aWB
xAln9rMt/LfvThG1RJbb2Q4NKxOoBUJpFkkpH0kFci9NwNOmUQ/SSEJE82KcIDLR
NtkAQ7hk2HIh+C4HkokRUIqF82zHmB5oGWlD8QLQKbIWaZinT/vaVfrzAg8wysf7
dimiM4TA3L4+hKW3ULv7rLhfZRfndG4c0LcNdozGC4GI9WijVhKJxTEe8mgmpL7f
x+FW0Fwk70ApPimaX09+yx1b/uoybwk8LwIlH7N5kwi4CwI5EWQpL0Bhdu9ga6qL
+zJgX9aXX4m1qaryXlQVImV1iFCeHAtKOS9cyChi+T5YKWvsPX8Dxp0fNat+EpoJ
OEMx9G8I+Ha+6Ct8uJhJhBgO1WJ2bZzZhovkg7PM9hMngzYdDEjKbm3YIe5TKg9O
pEGuhYIGiH2FBI4oQS6WQS0cLGY1JYlN8B3T3CByCRIBZ92+Ky9TDFHj/36OC2Aw
xfeRZFT/Y9jnFhvN+G0sOGyad5Lpy4bRoOa7hps3Ltwo6fkcuHxurTco6H3qucpG
OiA7gbai4e/G2UGXSicnA6v5LJxFVoFe34ot3vYVAOgDXbLj5Eobp5CD7wXpz5qX
+VdsijSHCWKQwalQ9PbURFbuAAP4sxi9x02WubiigbMkJXjNdfOBZe1oUreO3IoL
qbCAD/kX1wOc+8tWxL66Kw+AkW9XW05mQZMGcyK2YK1+XjbhCjDMOww6VHJI+8UO
c63zHnGfpHT4a7lOc8vaCW5xspSjXeKW9nLS1+PTXX7zlcUYpwjiyS+E4pV3ytlU
h5Pn4qGYyObe+Wp0hb3QUJvHkWCAFJtumzW+Snqh6oWEVfleRQiVAIeEw2vZ5yHU
65SDjZKe8wPm5svj+t512w9o0NyiK+9hOocGY82ITOxjRwRFI1QkFFLSlrIhuZid
fD4noSAn+tSqC9NagQw3A2ercWgWd0+ium0Z3ubfZX7zOXGzpQ4HqESE5hqd95Jl
kWA4LvU5Uy+FBr9I4oGfG4F+r/eYKS2g9G4OG5Sh+p9pcH/4XHNim7Ff0oZAOO8c
drbwCfn7OqLYckDRA2Ux3Q==
`protect END_PROTECTED
