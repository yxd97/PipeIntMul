`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
at1CHigh9kqQkgv6Lw5g8Ho3IBgOj2gENML/VlRcsbpX41fyBzbOk2HEb/SI/nVb
j3LgOjh17YdONZP2cM2e4e9VxAp9dIGl2TP5YkF8jw1in7ixKjEEIGBXbrWSt5Ul
0sBdOOz/7Od99pl3dPyScuaxxvAEdvk16BrEtsUHrQrC/kBtGPQhM7gHR1HPeKGw
fXhTRvTevt6PBjSabsU36Z+1KzSR/XJTnI2/F9kjUQyRC+vmrSOHgJ3nF4S+RrO4
f9w6lkIjMRITCsNWNDLMqDvEsH21MsEogMINISLdUtsWqBaXgwG80IP1ZXKLyKl5
YABUq9ATSP5BQGC28VQsTADX87CWCht9Ini+J0fqZ+9nE8bDSu2YfSmCWy4dAabG
Sq0EaQmj2/NXbueNtrfgmgJxWghe6x3oirh/GqFaNBtA8k198WlMmrXwnDPE1Ptt
e5MxH+5rRbFkSRV9l8xxejICuaHCw0VkF3YDDUDNym5XkKtTJfgKHlyUYUFcLYjy
gzuo3Qitm/qWEgn6jGfSl7QWkcIxzHDrVwXb1v6DfJrhLsEqcEo7dAU8LhUXPyhu
q+4JgzdgDP01d+wHvrBXARTzPdtpmXD503jImWEqONB5FluODvu4f+bn2QEV9sPf
uVWTgI3K+LAPRj03uViPpTP5dx64JOU4XmpM5QSLs8stHDx08PpcBmqHhJ/SBmCG
omG+OoAduXcxdrYs5VObK1N0mR0GIz0JnM/9lfMwoUloRc/w3JJDYyMLryhrH/g0
EachUjWUzJvCj2bmYA3dx/6lUfWNBkm2svDyfPs1s6LL4OqiwocgGou+Qw6GcsEb
jlIVQGjX4WMEKT4IGJgVW4wWAosdtjQJN9AmmZnGNHOFbFKD99W1OJFn22IMoTCt
vD9JtfQ8ZdjN1W0X+DSRtz2GJZW/nfRKOxonHdrEjyqD495plPFqg8tjl3N8he0/
ZDnQ6dJ/mtaNKC/imf7FeQ6EwBQiR/vkxndYbgexFUTQY2ykhOF+gph5bG9wrbL0
dpRJhkm2pCbMsI0a3ILc/+quNK73Bh7Avv+Pz9FK4eHCuxDVyqdSdw1Ykb8BUZq5
sEEA0mia9wLR1HsqhdwZq4Qj+Lk3yQqX7Rbq7yrPi4U846fOkvU3uDqx7CHkWT/E
jnbmY1ORf/PUf87ik02PKGNYyYAXaFAgdVs47f14uhbgQZlUalvhuTqJkM2QZN+N
TLCYXmF1wsP3Y9LDEBI3SDh1dwjoYUAaDyZ/Gi0tTrZ0QqDfbcQzbfhjsi/gdwcb
aKUo0QYpTxG+UBjZCT5qcKxqfZ4t1eC0NWS0yTxEnmg=
`protect END_PROTECTED
