`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzxIZxk9KYvXDlKugDVLRx25m3p/5vs2Katd8VtNGTbsw388/JLyd5vtt6ecLet0
N0ceUy9oxJ5eQShYYJJjqUn4m2Pp90ncWbTe7XuekZE6RFdpJ2omusWv/tM5gcSX
o8la97iosoDpOE0DBIr8hBfqkZL+nxKMNt3jPrg/+T7YcBuztCguPcjvtQ+DpveO
2wtWXzA5TYzihwO0dW47PR9ATL4od+nnWKwtZDBa+vpXmc3ZkND09ZluCrXOpjr2
TJ4is891qXjvqpeNS3de8f/T/wg9v7XxxO8t3oTSqtHZ4uG1KCe6w7fvLLUNFLbl
V8IIbDiVo4YkiBgFgsWlN2wwhnfC/E6G9dJNptukGtwHYsbyP5hAVFEBz86AUBss
530yW9AXe3aSI5sCEJrnjUB+XxzRfQ/sbzfI3r9dDznC43EbiuT+htxNYCZ+n/vf
0Cq9Q+NrvwF9xt0sBHoeUGCZrxCKSdh84wz9Qe+Kofw=
`protect END_PROTECTED
