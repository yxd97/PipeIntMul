`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xQogRA/g2eeUivtha27K33IAzCGOSTPQPG2we9OrGQdbwl66l69Lu8PKlCCb2e9R
jZe4TYfbOiNEPEgA0KPPy8hcviVDNi9Yx52sM3xXzNl0PiQqQm+qI/+BNeMRNt9g
XulylFd9k+0PUSODpkKHdBdLTLqKdt/Dt/1EUkdLN3V9k7aYQ8JtmzSGwrS+dASP
lNYBoyiA0V18TygIqn4NlfNYmg3wxRImt2FC6Lu79o96btrx+D3kDUZHcZmMuf96
3ndZ0js++h8AAlhnyl6r5xhnazilN298xz8jr/vPp7Sd4iTaWWOGGEXP5VgD6Yp2
02wKhqOWi59p7aeeKUN/h1vHLVwdMg0i71whWVxnj9ZHhYhwPlwv5G/2m1vmbzGF
CT9Xou4UqYoH7MJqJ8ZTBJiEY8BwD+/rKsgDVJ8OqG8t1Vg8VUlqQi3jIWoKyz3P
0Nvc6f95mLWSi0x/rbArNEyHLGvbNYSHPZ2h3ZcrzygZSXRjuoM8bCvJAEPoOiSi
xUDL/Q+RaUy+wATIVtXkLpM14t4J/HKxIkjupFmv4Q2qYLdU57J+YLJC1QYTiR+m
QIboAwIJpjErm5yuj+xnbgJh/nLgAb9echzAWZfkskrioeHhIKDuDA1SPYFqRNV0
qS2qSwM2TKum3ABLtd3ubg==
`protect END_PROTECTED
