`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zdd2Gp1Xyuh0pTRDyJfwrFKaEJ21qVz6atRl0A5KPIWu00w7z/ovmAYVdJCb+QW
GHUgqeF83+Dhk628uONBc9wJSkDHp1fr438Pj2DR5Tr43DI+1VrTwyZ3edZbHVCp
lRwrdOl0/tm8cfwU8rdaXffPB4QXqu7u0OHFEq/DA4LkdeTKSb+uQHM4oVEW8Rs6
qNQXzCsPko2B34tbP2F6lnBfuvQN83TmZZ51cPJDWeL3mNWa4KNGyb+/SVU7FLMf
p6mVjodNEYg/FVDYEMHwAi5EXVWRm7F2xMkgQw4DINsjdU6d3tyEDATO/jOftw1g
XXqjPNUg8F/+xmt2h/ttSw==
`protect END_PROTECTED
