`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qOv7Gu5sJtgj6if1BkkFSMgQWzeB/1CH2t3AFJwbyrH2WcU9MKQQhs9LTuTOSc5M
+gYWWnKj++dEMZ3Vu7NIvXKIfW+VXT43cLmxOGkjkfC2Ywz1X9oLyNkD9mfFLeIq
Rwr85B05wOa0RIEfgHvHMqgzQkzMrmLGGKeIY5atmGSkGR6vkrdL80XwddZY+P6R
NdyAlc+kf+FkhORF8UfHzYwPbeUSuDETUUDZ9wxJpt7J6kJMGo94HmRR9pSf2Az0
QwkMtrzTrUJll5vxWBkrRQ==
`protect END_PROTECTED
