`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TjrUldySeedusogNVFGbw50Jlt/PcU1Nd/+4RrWNp8Jm6NzB0c/PspogiMMY+1ii
ty1yvsQsX2Z5OBp6UNFwaEeB1zilM/JmJHs2cLmf+XOJsNnM5r9WCLkUe5202l9A
IETtooO92ABe7IeSMRVstiE/G8uJ5HWCN8FZzfbF0nKuoabshC/yA1gfaWH2jU1h
XCKrTCl2NpStorwIus/XBNfr+cbJAdbLhDON3kRLQx5RQH1GRsZWK/F04QJ7WCT+
H9JlrnmOxQr8X66nn1Qd97SPfKDG7pYHi2jOG9QSV4nQQhl06gDdwmvGMFCYJ+ym
D14PI9ZbUW5cScTN8elK/yGCoHsUpouDJjzBSP7IzTyVtrpifui2qEmh4HpqyFwf
QLe8YcaD9oWZfACJzwv0KRFZtWIHsZt6IKhl8+1T9L8=
`protect END_PROTECTED
