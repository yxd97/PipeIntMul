`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TeetN15r7Qh7y4QSIAf74VGJRKyHgGe0mn2dQJ6CLCeqdqrwmRexDFYWdws8SiA7
eEr03FNyYuUF50TOhVcujvmHfGWniEzTr6Ryk0nXNU+pwUCFc4yoSzPheb7B4Yqu
mlAT0xZmJA7hBmWnU/+c9L3MMcfV6m15HBcliibpcU5rZKw+iHxXMJaVbpe1UVLs
Iat5WmINEJYJm/RR9t9Ivc+GiQxF6RFIUUCiCwYFpqmDjfFqmRN7v6P6GLcL5F74
z632VBOppj55wMPFqZ5DoRAEJJJ81t8rBQJ7XoIjosAEdCX0QgBs+F3dy/qrWKao
Gm1jivRxSvjcA46JAZzUEqnwcIknZXc+dm7LNMh+HB38GKv1oWUe6RV0/8Q8SrXc
yxN6TyBezMgFQCGowGA5F5qMMVQnvjdz/R+HJJaHUzxFupQAZWLuQA0G2buppJ2g
GyXPe7RoKSiG8827Wd3NOxw1vItBJGk3Z/A52utAdY+UnXXBCcedtSycDtnWThlJ
2vLMBaUujfo7XlvwE1CPxSgnjidKzndldi975XGEm9bK5JCGSIZzamQlJr9VAAik
THYJfa/cjWR0IyTVyl2bkwWlbTdKWUjPvY3s/90IPrJpancTeyNB2AH/UD8qXKdb
2SMKc+wQaZmZuZoUzudfuHmNGKHlg1VEceuMqeirmHM4bK8mSBVuMUp76TYhZK1V
cdN48/Wk2PenLe323bSE9yEe2fgUzxt6PyIGGQyGptugQwpAb2lPDxl2yfhukE1r
iSkVvzSwCuJBBirT9yQq7/dCpxhEL8IsoXFay4tog2+0F/AEt5gDthbwe7zCHS5g
U4gUTQiUvHp8i+QSCGqtPj2ZRk0YljpgDXy3bsnCjJTkMfUFKqJFlNFX2yPRpeUh
1lLmYbLPPK4WY8KBcMhOKnHp/k0ZbPfJDDmXMf6Xn3ad/MnxDLN189AlDQnDpZ9+
QiSwLJZjULFiJ6Xv3x/xIj6mlk1B9TURjcIKATjmYe/SJl9JJNYgGaYC5/u8aFJg
RCXYnkR7L9iQPiOhpfUsgiftApsy3gFdDh40T7vrldA/LAnAf6dtpNZPwrVAGcDH
ElWdNmGG1+6aKgQJaH2TYXIGdWHulk+2Bl3oBDn9h2rWdX/g7+k8G+f1t+lifiFz
u+mTxdW/CqHYg4vxINANeR2jpPl5YWXvkYppJj67lbsv+V7kvIsWS0o07bgLO+Bn
LwCHN0WNUayOLE3TtNzTHnXu4cTTVFnFv8QJxq0Xqi/GNoyUv5eeu4SuXuBimowg
8aK+laTnKZ1V+17qtuaadL0rSqvmkOSDJs5thRbqaXH0h5fhXJnbM5/k0waLgbk5
LAiJG46QmJSvDc2buvdF3iqnlc0C7UHoFvTt7FWG15e2lfHqDilf47jHXDxL911E
aqDU5arNT1xFRfnm0kY5PivyjV0modlWYyS5d3stDZJiHTW+q42uyqTEmSMmcc+R
`protect END_PROTECTED
