`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JxuUUbuf1Joral9t8u42JL1TA3EFaUkn3qJdVabudRIAv8z/Xt/pxXOsmij68uLM
BXVvWioQmx9olNkbiHjZASxilqrzRr0M5MRV2f8acyFLmv8HMEPX+BZImSNl6/sK
bkDAQp08GxZiV6cjKibHFbPWjcAFKJygEvILjh8Fqd9jC9VTiWNl27XJZQuidGZl
qaWtun85XKQ46IqArgUk5rNkUoKhnclTxDpwVKVTCcoH3bErMayqSBBxRDWp/Gyg
jg44yXm6OaU8Gwd4kZh5tI7sOD5bdWEbtfj6KYe20QgWNAMfuR7Pgx7qwIT+PUol
5BFefZ0bAOcz3sm8OXPMdjXRExipYCZh+kszWJSTIyrcHQEQOfiIfqWZlh5JSNwR
zzyYayS1XrmNJO514Zuqv006ERETDDzRB9+bAeplEyk=
`protect END_PROTECTED
