`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/yUn8Zsh+imJejS4S6nBGK5jkiCiuoSfATzt/Zm7VhGQyMALfJ76TtquEdr6r0T5
CaQtf+8ggjNlLVoTMt1UT7yIII/XCsZw5grlErw6SsqN2nbKsyE41F6MbBqEF8rZ
cRBeB06kJORrduQfgXZco01r90+GpOBsoemGxWnkqULo4avSutR3dnXzKcJDbZJX
v9dclGFsZ9YnAHF0nI6WWY1HCD+qh7YIpcirsiyK56Q6yFM1PNZzvUhBgOKD6LWz
+uOjk2nwUicJXPba40DSG+dhtbnU7zursxUeAE3tnT9wL7pXH7848ewY+msMdF0x
sRdE2H7sseqtFBQsX7a2tk0iihPu7n7S9x6Mwq17Z8mjNxcHzZ3MKM5v46JfzMm2
K0AeN6XkU0qbXHOzhsHPps6k/kxwznnhoEgQibsDOIRyUrXQT0Ab8ek2GpJp75P6
xH/rykl4E3655XhY/2MRRkqpxwtQMkeCk2zK/2hbW7Xqm5pmE4duK2UlBZPi+b3x
PgCygGeIrDvmufz5uJg1zqzoz8dx0sdvcKJt+78Zbq7iMPv1wwf3uNHaFLDrSLQs
Z61x4kKXaa4osreKVYZ7wdNopLD+LiKuZ8llEuO1AurE53QKLfyVc8TUnaaEMu70
xoAcqbQPrDCxG3VoGqPipMmTU9U6kfGDvHB6SDeibmE=
`protect END_PROTECTED
