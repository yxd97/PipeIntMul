`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jSpKf+fnJo32oG6Zxz9asLmUSxc4DC484b1sx1y40cGSF/D9tRJLyAVWlGh9xxC4
VVnXjtDxDPSEtOM4Os7YdoXvaBCBCq2sjCeIiBes1T8vT8IE7FWhpFjEzZCkqKJ4
6KZ19gfWSxXjt+nCnS6o80jriEyTQq6vRRlv+fWTp7BPF+U1XRP2nU/m9yRU22XX
7RjClLaexkjqm0EcaqanYntPmar+MvCXLXB3Ho7fjcdQxeckM32KWnufy2gx+IFr
Qh1QYDHG4NIZbbN34C9qc1DtMT3qMAz2xBG4/jktwNQSj8zZVb4mFsHsy5zcEwZc
Tq3As6RaZo5zndjhgQ3DCHI9hy2zMfERqVdi5K5cTSP1814WiW2xzaUBxa1S9BHh
Hr2UVMlgFeQkb3PMiJn5umTXMtO53Mflh1VVlWchBYK+zMh2V9fioTYaCI4O10dy
JXhR0NWcCmS8uxnueHZWi2wZbbACaIT8V/FxGa4cYoDUY5ZdW30l7dliMy/mNq8s
Ek2KcvdPrDTPQ8Y+/0R+KIBO+7VvHoJxrPpS97VO7bT52xEiVZDB6eHnQQr6rXVR
fEvmhi2WCIsYjQXASriWzx3j363HWrRa6qD1ToIBlPxegI1hpmBCJ/+/J5eqKoeq
yjT54JxXm9W5/pMiJdKbO+qFK/xN4VrSg1uAZ63Zr2+6sl+y+soegFgBgO5tsMHf
j3TBM+7ucOq9u2HucSgFOApYKigw9MC0a+OKGetHa1qpIkICXm3e85NTeKHIDpML
FH20C1qMCf31KZRvfUJxXA9oGJhB4cKtXsX/At73taD/ahW13BOs9Up4z5Eb7jT4
E37cGWAit8lFc7nVbtjsXmUoxThhFd1Zh+B47NgZP2ydp1fIjIdUmljNr1s5CxOU
n9f0Bo2E4sguz6/O4qt2k9QmXw7k0BCRsu+N1jglRUvrLVIpgARFKzAePFjLYJoV
4LbZ+p1P/IvdiAMS3Dn6zH2lkS1HMjAcZJRWRwMI919HYnwCHnWMi+X3UH5RZXUN
QBTW3R2LlJ9zPXHZURcJzQpF+Vn9w2KRqt+DbCZD+gysU5XpJAOeLTnhhRXRZbUC
a4Je0GMYhLSYGTJdDTy0P5MWcDEctQqjfC5QaIoxFsnaWhLT7G3Sb+HoZ6HFdATZ
M8qfD0VPNDr7+Aj3MBuoQkRvtRINeA/ka7tfgWnC8ddJbdkEwqvpQZNwEdtTmrhu
dEnLPkFANf+HK+dWiQWt+2WTUqx/R7MKYKnvt6oihKw8p6lGh7O+noFb++I3UeFa
OQZkbICIJwq/O9Q7QQgr7aUQFwnuLPJDZ5o+ekcOphhWwg237jwdSI9SQcOXtRMG
S+6BgV5/O3g1pvcJIOJXCuX+7VKfb+N5aBcmQLWMzplLFVJ2e3Ef8nKEKzYoSJmD
RWruDdh4LgCs4dT8T/9LvcgkKW30DltCRKtXRmihXK/s+z+oj8aTw7Pev4v2slCR
Kd4w0F/L9zcXe/yvy6jBwQ8VmzfIXVFE2kOsS3VkMSoHgSMzwoCWNfnrjuBcGmol
jnwnZW/Yzl5x/cOOF/BzpZpnRehTs3kR3BKNM53O47Y0sZwf9RN8AW7ZkQeCt26V
+KX/oyGwr5oZ24NUiaCz7uCVGaDmvq91KVdRZkc9FfwxUMNAzM9g+a8U/TOjmVbW
aiQYod6OoYPKjp8J8kdopqc5EBxKMN4ILu4jnqFLrlMFDgj321rmV9rYy/5khUKM
XTGPfwt6MDy9YQBdL0JEuHUfFyE6uPk4CWGvhkzRiIMZNxQSLf0BuIKouEfpdedP
0CrOdrinDvDAmMUr0mFEqbzV/C3h760v2kCCp1rQZCNngqC7F7Qp+towWiSJ9zyQ
64T1p5RNBkDyk12f/61K1wxTlsgunyFgl4AG8vVmqtQ05GWw4wY953yfnubHJIaP
Q9KJPSOvQvZeUmwVNN5Xb94xF4CRAjGlQbFa3t/cofsmAsI2tR0xj445U9GgdGm5
R1QHIeTr+THYdqHoTTChb/Z+oj1wKQSbow2CzWPeBPkgm29dd3T3wm4Fu0k7LE/K
wm2B1crQ2OZKqJ1j9115GbnkCaX6ymAkIZeoFhKLAPIQVyGnNVkIcg+GnCMApJxw
Vfvzlb5iLkTi2ypawtix5JoHZO9DkLpHe7GjX47S0tAgE+3PH/z1hy9hAOVjOCe6
Up/sE3oIu2SrpuPGM7qXalaeSp4OfPIBBTKZQ3c0EwN91TLsYT1FNmh/T+AzY0og
+vTsTi1SPlHcjQn/nznWN8yYCI7yRAFET3VEmgeGzAwxmr0y3fc9Jf7lJ42grQa6
1g7tmUlFaEDIZIK64bHe0m6hzPppXaCYDYqwABHLmjc=
`protect END_PROTECTED
