`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YcKJSJWyYVm3wvl0FO7DDxTTnhfQWy6WFuT6cQ5tjBeGMgojP7g7LplmOShbZQbh
BmZNCTEtAzH+mK+YfyOOC9LGf0TRNsZXDQXM4bwnRAtzPWOsDS4Dv3kWFXGR8H3q
YpSPYMSmsPeR5S0Uru21JyLGkjUYRZ3cHbnDZXyKTpzd4AEMrY7z9Tc5zBeeEdGH
id+K9BYyuLATP4CXbxFvaMgb22R1izG0ZFLT+3fQ7Jo9vbgHRlD/pRGjxZ5PfNiE
92Q/uF2+OSfAiVxb0CC+lg==
`protect END_PROTECTED
