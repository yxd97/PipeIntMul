`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdfIRT68vXwUaAoKE57AKiCkVNu0GXZeg0s0Rl9QvM1b5CdVzP9HeIz50X9rHDRj
w6SgFJQQxZgago15wCBFPivdkye4hdZUDjU7LSziXXkujKZr19wBz1HfYY1jIWRb
EmJE8Ueas/iEz68PGvDULoww6lqBoxz4l8yNFFn5g9fIwHJi0DbM9Jkas9RIZld0
0rHvcFFBvkM68qAjU4EzQdNXzm5PGEPwlgmtKqhE/hqrfddCPF3OEhlulPq+t1fv
SpjzJMh6Z8YIFNy28qH3GTEXGTVXweaMzMmuTNTmD37xPrIF+D4CH7zr5bb1aBeB
6lHIwIoq0IyO+EFEZbBBZcAFf0/vimMzGRMbiQbv93JrLs7IxPga2mQCPeVKqMku
c4HV5eWs6xbiNgRAxq9AK36nyY4U9woXpwW+RJ+kGqE=
`protect END_PROTECTED
