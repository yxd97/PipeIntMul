`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uH2ZyxElT9TPkAHOtH7Vkr/At/aZyfckw6OohbLzKEEdiLwAJCtqk7oVXKZcymAv
bIAHf7cAE1lEzKgnJdLgGIA7AnjXuLp+/A+rHmXknCqE+ga8tTDqIihXhJS8UN5G
kJOK4eabuqLTSFn5k6VyZLWb4qtCNlH/cCzDHFzHkRCnLk+m9lfrgg4pH95XadNu
nPifpYHe0/YyC4kKjkRxSRH38ZKSjBbaKv0Mb9hOBhskoGdBdqWKAVNa08xM14V/
uOKWF2nVjzyYDKsSHH/x8XRwbYY0ol1rIq5oD3E4jIUp1L+1CH2DCdSA4C68xsyB
2NpJg8b5oSPBMQUWWRK6+CTUBpkJ138b2LJAM+h1fZJOtlqB7BktE4OH1BRdqBbi
nnGfSd2S5cveyfTSbAkJlw==
`protect END_PROTECTED
