`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n66xdZuD99HcbX5oNm/HYFvU2Qfcwwb3VoyE/jB4a28uJBAhCz1OSQxVAOgWJlyR
wJXQ0+MhGbQZqT1seJOSml9sTZkznbDhcQgejZCat9i2wMu58mWIS17OhJMrDnXE
rxj+cqtqpq7cfvm3AE7uqyzWC3U24rJ/CI9Im+oys7XyBhS25tO7r1p2nMY1PUUo
zcAGTaNFLjQUNuErd8iD2nc81L8/C7rOOlKEe17dmvZ8X4CnxIUZ3ONsY428AzpQ
2U6ld0doevSDrZ9cUjFGeoUdd0alPCZ8QIF9ZOK2QA4hQmR4H5yygyG5pwuHPcVB
Rt+f/q/M+SQVdFk6+4Hp9feLmM7Cu8L4isDdraPjLPEEskCaqqUFHmdB2ZJt7ieC
DyMxzKpwNjwXQPA++fFCVJsq/rAdKE4p5X5EIQloXTxtCTSluSuVL0hLBEztZR13
RSrvw7mac3nxvLYsK7HYLk6zzxjlSftCK4Y+x5MS8/yAQTruE/lyB67ebpABoEpp
xEuaj7rqdq93Siq8m5+zQz5gtK7lNmBKno5WuTrSuVw6zJBftlyo/RLp/roY6+df
tljBto3aWsp9FlK08cM4ncZLVsyo1OKu/gYdRBOt51R7kcoiaXo+0oZQU/+Z5Id/
NEZDukArFUAa0PkuxMdDwDUFnI1kM9HQDmSPHnYD3JM+aG9tkP3+2WDAT4NhRDWn
nFb8m3SdySyAO7RCH9+BPz8yepNzQ6acGVtEa+6Mr38optqlFbNukI1Sm/Zj5Abd
31rDoD65jFBNlWRRc2qNc3ht0N8M5xsOr0BI0jRvbz3zb5Y7X3P5DVCFw/it6BP5
UNgjQzbkPoC2OkBMZ3MUEpQE0rAR5W9CUvqYdpTBnfOCBxq4yhCZwjUTwj5QKbSN
pHbgdSywSYLhuJiwIgM9oP/yZVWvUTGKyfgpqgfXzOzUv2+FB51IG0kkK5NGKUsS
gd5TRjJROxcdO3vG93te70w8jio30ei6VUOgspasonpDTxr9xC6V9ERUdK3U8Etv
+S3b1KmbuW61/sMoNW4AtTSdNNjZqO9vXIGl2b8/jf13vGccVQeW8yxmwAuwadxM
dhwGxAD3jBBgI4qOkh9fgyBtr//uzLb67yJLFgMJP9XHmN8g4olrFm/SfFy3mnSY
a5j2Ui8b2NpaZQT46DyJaxBf/XSrVFF5pU1WVVYVZUhHzgCrae0VkLhmX8aFOcdL
4DPdiLvuCQvL3nnj3DhpLpT70OLd7rUbcC4ct3QpkwE7H+oBL/tKD7ZCs5wDCnst
p6oUvfFvYqvuYsCXLrsPOgAU0kiqrs4tVpundbaKbeO8CvWF/Ygb2e9tObMwoAAF
MK2YJYSyTU6S780V/10avUB6v8bVUXQ42ducVKlwCLQA/+RiZPG4QfKuBoHEzSC0
GWZxdVv6qOHlzC5hOoXostkhqbnVYPv5hOTHWLCqZIrEtf2657RrFEP10h6f+nmc
d6zeItwmAM1sZMIJxZpZsegurCPBFX6A48BnruCmV1iGEhYH3tk38Jf0G011mIpZ
ol/8iW0oCmIIYhP73Xc+ByhPZ70NOFqL/9KtVGlbv/Pvu7eNCDsvxm1NTkHiZTfx
254+D0Y8DT5WZuyK/J5U2WCVf0CUCXvVFYILGycJc4K4xPBTc6kjSQvBww0fyfDh
7f4wgngzpftkxim6nBc0FEqLz3tD2GNyGhpliMH0xz0Co7u21w0HHtLGS6UeCUQ5
TBRIYeSQ+HMn1f85CcuLD0ZgfZmrgtBQw+1XId2pRfQv+6pG+dSKrAFOEE7W3NxC
S0FlIeOlQvKPrItKRsc1xEma1zaLBiLRrKG729G0ZwPcwUYRzJOqG39nHKN8iKIC
IyNv+wwji+ezTd2ur9seP8oa6Kv3hyh7tuLjEZbA/ucJYlRT9T2oEbH9VAlJULdt
H5fApw0neihU24pIAWJUmc7w+caVZ4jC5o7jULb/9tdCVY7W3C756jVMAfgqJC7e
CVQ2YLegYXBI12WLKzH+6FqU+cHHWiIslRkvZ1CtmeQT250jvskAtvQFtNE3H69n
0bo1wFmsxjk5aHKqC0MrNDLtlDhj6j+ZA31LPyhA0S55kvtAbhrrFFXCPAGWWvt6
jM2P7q9g51HqjWbu0F+Yuyaxj1OJE+KQFC9wc4xpHfAxzX+WoRdCIFX8i12Nordy
7sCKnRFoZLOTZgh6sfbBjM6SVcHzrnDokidSIICCyEWiwf6/+0fbZztIbcCIF+7T
kKPax6NhzXlY9k9NRwhk3CewVQXPHz84X3fd8IBWnr9C0yKCQIDQS8e5KVYtpMc4
UPVChXfz5UwpAPraGVDeGStploxrKxdgdFJWAHAJLK1YebnDq7M03hkA1H9lOtF9
3G0A+B+KeoJ6u5qmyks7QIWu2xuwWaDAg6fa5ySuG2ARKq0k6nzfej3Crok0bbw+
tSZWCInmygWbVW9Wr80Qt9a+A+CvCkWEiGgfjG1l4ZGhAokIEkmDGGPeiFuJ36Zu
LKnWGyK9tQ3qCVFnm4nK95ZNxIphlzZHATXq9j3VR8IBXfdrRcWFor6GP3pZq4YW
xzH15EuqVFAIhgtbAy6esWb08MtbLS6S4Jgrt6pARxfZ6qD9xyvX574TAhDoPqvo
FAjmwyz4+KA7a5boDmeXuO2Kh0m+ZWg5qY3v7TPOrOHegawA7ABOA3s4q0QgTtbF
wB/CIAkIWiGFO9vg8oXqiirQg/+rA4OQ+4t1osxsvaT5vG6bvvAXy6gxYsXR9zUP
BAan6L7E23Mft5hlHvFOP83ggQYvoBokO4J9V/9FFH4w4POCdKQ6PeAy8+bXdcQk
KYFs9XYVDak2du6BVTe9QRDBSqZ1qgCnfZ09OnhbtqX0NHe/9dM59SEuVJb+kWhn
V2D2qwEhRiot912nOjaswtJF8hTRTuYz3cy4hokY3DRiCKtgNRMJtnjLbLlutHk+
3e0Hbm1Dva9DbVKkl/GiCoMjIQ3nL2CSJaG1F0M6PLd7a1vu/8xuEjft9xDBejS5
sXGPRiCKREJZfIwkpGR77jPRwpqN0CnA/sxZDt2Qyjj8uDU1tRmTUDRJMlLnAkpg
E+1fj3Hr9ASnOtySrSRXRG9XpM6d5EWv6SbvgFrn23JWSgHKDdPUYaKLSIA5AgzK
qsgw79Z0GJnp5k9FAL75cH2H7FreQWCnseYZ3RL6KNgkXhpOxZiPtGAnplhSrVlZ
dtTc/lAj29tMrg8NOc1pL0LUByhQ+yxa6MJAUj65aTW6twomTz+6eIqgoRawo6kf
oXjy0LGb2SSE40aVU3Apb+bb+yoma9a5b9J4ASpTii2SN9/swWFfyn0sCeVP150W
AOsUeU8rojXBV8jw1ef2Gi+5F1r+0Jt62e4ofMoId4EZTXveK53UWh+3cvr6dIGU
FCiqTnRNBIAV8AIx/N5zFUiUGY53sLtM//1x8zWraF6KfgghWZZ2Mo9bS1XkaKTI
MHe+yXC1oZMbSeuP0ljocWGzvpMr5g/LRGUTJ8REdYjg+SR1HMo/jaaZQ4PBh7n4
7bWVEwHvGnRAq17S+hbdJSrvZOd99MC6nTp5oOrmbJ3yvGsvtfN4Ia9/UofKyd0Y
RihcKryUsPaChpqwNuJK9gAwArPOOXMqa6pcsn9vnVsOYaBT7gdM733kea+ZbY75
Az7Cc9+9GDLT+FmM5GMXCjnQd/Ue9mZoUWnRvTeP8RkoYHc57FTq5a5am1pEFqh2
OOsB6ox1z1VCjfyJSZxKZyRrcOJ7iNminpE6Or8G1+Oc6Td2VH1U8DsYxVObvbvW
STmb41Si6YaIdNqkIEIQDncRhgCRsXdEHjensZ+tkVZiHA8al47ZZqRv8DFtU4Bp
NgJ7AX6uHzYxyD2pCWqSP/B0InFjpsnHa2oAqHNnpuz52rfB1VTU9mShmifIozUU
2IQNhupDTN1c2mmMnCvRzWxGW2RJzUdM48BWaqfBGnO3zFeDJ42B/Wdopr9UdRW+
tRAoBZ3QCYYIpyvIQgxHjF2VchESQlAMY2uG+Xab59eretumJUNwx7QIGP8slCR+
JcZdabv6Umf/9ZVzXLU4gp58XqIYGP+y7aq/ywNhxESTsxTb79lUZZXHotyUOebi
tCWgMYfUhL1VbGDjwjfFLiGfmP7EQzDm/ptaUNiBhZOGdbwq9SOOXRqtF/7DC+/n
rwSWYM8acZpZPMgRwdNn5KY4f+O/De1d/CN3SqHOu1zwrR+N+CeszhEw1yRNjsXc
9KKGB3GiawvmRgkoImMpE4dKbCjkUgCQJGT7i54sf/H+BuCY8ZcuIl6YwU0Ux56X
bYAvI1wUrmIdo+/TKEVn7JfqdhjhUL7idxYhXZ5oRgZzbo1brxFcO1qWNA8/wKJE
NrcyDw8KktvSjwxqLrEx+4KCsNStbNKCUAtXR1ZPs3IYyVoMi4+Fr56OW/0gOBVP
ckqH846XWGJeNFqe9gVDMhEkN8BXJYr6AGZdTnH46vSQ2SAvfeVkTaT5qignT8tl
5Qj6NHdfl+0ab0lq7pOKui4rBF4QgDpWErL8bTD4FrnmOnRNK5F24c/bceT/uxyD
N5aj9y5MtlKq/vKd9q59/qWW2le0B7ZnNsuV9bb0drvwCEjQU6bgDKl+u6gb9TsL
G+u4q4ZJzhmQVlug9ZsMd6mM5Td1N68DnxlyDOScqkXVHwgo/UozWhJdiEbo/zDu
XKulFaA9DSUuSRLEc0iUOvkjGUFEzIma7FHcf8Zf5TFaQTbuwkbnuq3fcti25SNN
i7Eke0/w8ngeKJVlq/CCY8YyyIsqguNkNJK3rLuzVANIlhNgpfd5UCNcUhsIRh6L
Bi/ABO7PGn9IgJd6ukDxjAX/HyIFRu5y4hy2NUT0iDqXXv11mkJVI8czTIQIEZwH
3hSluFYUbNv/21Wb39JVbu1M7MApYQ2H4B1EO3ZZSKVj5AtLAUPHEsk7e10bJpT/
UNAx6VLa16+9X4ty3Z27Nt/+BVJ/TCRvhEFp1Wv0GWv80RAt3312Ey+HcHbPtIi2
iXp6b8VhLTs7lIEZMolDKLvH3CBuOSEigNOcxYuoWaFTWrRgXnu2m8WVBi7tVYta
wspL2Qchq1J4U6KZQNOE+WjKCuv6W/wpgVKdnBt78jdD8EP8km2DMWEjun/dqVEF
8qWCT04w0gFUQNxCvpIIMtgf4YRMbid4tuZZThjpv6U+Ca6ryF4D9+GB9gi86xHz
1QkE/SbUDzU7cfqByo6Nm20IoJDEwM9hIpJT5hmzOUQ9OrHJuAjAdWMayX9Wo+vW
64bGgLXFPqmndiaw3JEJb4SOQmaJcc9CNY0vg/Jbp6gjE6HOYkN9JDg0CJTNQg/V
UH1+PXhAtRqep4Khx5Ukv0LbjhCBvGQXHFk8qEMVhJykIIrYgVL2yjGl/L+AOTan
lV9ymPTP05HkfiQtSU5BT9x0aW0IRceGr55bV0CpHmwrk/j1Q7XpLCC/CyHY/FUy
OoJbfvX+IdrajQoMOXKzJTXByg6O0q2G8FIgC3ZLNAtZWqny2gbansbk0pb21pqx
fXT0gkUrFa7mxYi9ASkEdFbbozfXlYu8p4nFeFo/X1IKfr0Py22Wkjnbs72DmV0y
kJAFkjd3nCuyq3xol06vzcOMh3WTbbdUx3ubiCq7RLEObTj3EoNfhH4nUZb/4YHp
dDhxsXyeue+wkFbH0vsInk10XiKaiui9QuDxnIrzDfUCIGAAKsoPmxYtrGgmjPtz
nVbdxvNDcyKi+I99Rb8dtHA7yYQ/+Cmw8CiEWDlOkiKvdY0cKJfP5mTAMuUaEoRV
8zqmzKVs2gt8C2LmN0BCQu77L7wNjiQPQAGihblWma4VxJbDWL/BRKxqZe0RW2qD
yyNYGyDUh1sq8bwKL3+2ze55zdgpMqvAITd+CIMmJ6NCCnM9SAgDPmJQL825QvGk
AAe0S5YSo1NM2S+piSpPvg3Hxp+LD/uOBvERVzTlgkzElNP+1n8AU6d+ANuYHHhL
+KvUPyfya05rufDfL8koep7cBV9VqkLjEx8hXIRtLLczSV1HQqbkOWUYX31rh5go
7AA0ujI/xYsvum5NBuW6lkrHaXmFndFhE38MVdUnKtH7WvUF4iztTuNCyUTUOVDF
B937yHdN3grhWsL3ZbdHR+WDqns1FniT8lgIBjpEDGStAo4YiRu8esbeEyl1yM10
HzB04Pqv+krUSluioYqnghd903Fe7zAbEWOhYWti7nDrb5b91wb1KyJX3GbhOl+o
Rkhaj17llLjNXw24/iBHdV72N+l5Y/hH8XajF1ub4jAXWn1ogzzuJeoW8vebXzRI
nGYeM+Sipic89HOMVHBhUkB9km4wL+GsAg9UgYkfC6qtwRJuUqHTwFd1Vdu9UOI1
dx7bGCiJ65hXAxi/5lCEm8lPGBcuhhzrVQujj5LNQhpp92V/4h5vU0X3UOltgtki
ybEAmcmjAw2AlTvwjPfL7UMd6PmTL7I4e7ALYEnAWN0dawPhlK5xlBBTp+evfTAg
0IGxKJmaXIAF+bj42+2J5+FJY1KUOBy3ue0AA336gKjRFZ3croaFkYonwULt2FRS
r/zB87YF3Ix9doaU2ASUa4PJZ2BFy4RcXrQCPTbyEPc4CZQhnFYyy0I+R/3+D8Nh
GojdJzoUyG9OXqavNZnXovFBsZTWpThEZPMVKdo/b7isEe386x48pGkFD1MlWII/
Ze6hrpbTCyx07mbLCpFJkikG3bFU1MVHNlUVheJ8p6mYOloQQmbs6naL8slR1JEn
CDcx6olzRp4dZNNJFTjCfyuIR5WYhCXAb9AeVh0Lvw5+myNFWGQlahMPdiqDDr6U
T2xU1ArEjLs57v1QSjyOKpx0Sracm1MWNrm1S5fK1DyP2sCc4gWKhmAenz8OSqNR
ZfvZOUn43eUCc3INpwvXkioUTBZve1bMg7T3g52UxZ2vfD75B69MPwBI7fr6xHkD
YN0MjT65txETNv74Pv9BLKukk9q6APJCeP3rxGbl4YxR5RAZqmMzT6Ah4d7mwymA
OCMfqQy3M3ulTwcrJjAaackFdmHxxfnxgNMSlXU89su0sU/Rk9MnYk0vf4cDVQwN
VcRWnZ1JpRum0rXjMEwq7VP/ILUPuy8R/eDLTOE4DEzwr19rFPvvqhi4XCHARbOq
bqPbj/SyVtTaqmEeQbxaIHkVlRZmlt6gVFUlChTdFz0lM47OwSZW7m2RLxOdjPpY
2GMv3mqv2EWbKHIWNG/nWnZl070RSwjf+wSJcuj9TVwj0b+ohpovnDFfRh3oETpo
Sv9aJGrtuvWgtTEdByb3ISvz1+A0c2FFd3kY1lRHDHwK9EmB/3xRPBomyfiFMF2N
pgsDKTnfEyCgDx7AqK+qKmPaZiR8nCR8V69QhshX8IQB+NAk8umvzMBMHCG/sV7C
D4nyPGF6cL6/Fn5K9zSEkShFUNhWKEx0N8M/nI71+BKCpxqJ9o4sifhEGJvDvQmP
KsbBBBe9vrvk8vZy8Lc8nH3CWOrE9WTag+5Tz3es//RMTwzFGFTF5EDh159zx3l5
Di9kN6OdhX1Tgu3H8bHwITuDpRLmiWu0EkFsCrFvFJc2FyqX5WcbMG9l2kSjeS2K
fBeLKUfkkUKOi3R87bDOa778P15e7UACMZfj8BaxWaqC4Jp3eN7Lw+2EH+H+l4ea
LHUhzDRxelIoMtY4ipWZa6MsI1d50CD+QsBe3ZKoU7MhvKfZueAVYllqkx8kww6V
u00ieSqVD0hAgeDwHCOQjl9AUGDn17lnC+PBNIlBH/SF4ILgx80CIPDoyyA+fwat
A/iq710Ob130/Dp3UnKiGHS5yMrdtOCx4FuwkZOhBxD8W+5H334Fo/Dv+W7bY2lk
jb4dxLG4X7o6CVF0XMz0rKfQBvv8b9iHM2lseBs3TWLQ5VtU57+OobVljkLeOmkb
fZ+S9++ehqscl96OnOr8Lr8Mgnoh45N9irUTA0n1ceOwffV1eNdcARch8ymxpejL
y6rYZs3HiHS0GzTRq6yGLtVo5qO8bPFkYawShWvdvlRzA8XPay3i9Qp5pWjyXIsR
753II7iQe+tuFVdbTb385XnDxTx0yQXtkga7l01sXkAkXqdAvE9R+XqJYhkwfOe4
tsoUFABShbqrz5Na54ssmGncoiat1cDvglP1xL/X3jpnWTW0J3ijC8+dh2+FhmsE
dfd+hpk/knlHzJl8GD0cz4F1TcsYBTPqpAeWGG6fqVgXINr+8p1dHOrezwy19Pto
8LpqicVVYjg7uGkk2FEEb9IeuQ0dPWNJwzaRYX+ZogpBBGE+UG079pVJW3kanT91
RWQj2p80zf8YHvZi7+xqrAUenMj1tG6bwD6lggBk+Lw3FoA+jBTQhoaFLcvdUOPN
TVx4wELyr7WlEIT5pw5y9wVXxmIECbwbelOcV5QKGA6nFqroP1N/iACYqXV+Hj8i
hzCBh9mqPzo86HDSlEFtrtFq942HiqNwHaqd0xK+f3/p0f30+YYVVlhFbxcNGLtZ
27n3/x62EvCjpZyXNTadgcTDoneLMyz252UqtzMeyQOCtOqH4qI6RzqWsGfywBi4
tZGlB99G0PWxRg0L9XRd8TZ2NimMc0dDjKmzO81p85CveikTsSLlnBEsLdvI0a7j
+XcgHUAqlJ26LYZUJqlDQ7hAVC6AJTyaGh4dAh4ptO5NslRi7631s5cst/9UgLJG
4ZzmTa8N0xM6BikAt6LhFCAP++oxZVuznxGBQiOsdljfHZdB9eZmHxttXxirjdo1
/Qdpqkws7GHjVdwkh7mIgDLs4tVLf8XW7ql89mxS9vX2FnZ7e6XHSz1VLyb6G1Qx
Mm+B2heyDuMNYO1135X9iA7gTbDNEeLjphaz10qAsXtd3X9dGRv5lBjM09ZazRzJ
eAdtt5QCYVc7vfSdWvWzxyiZLO4n4L74ZCICtUE3flW+5Viejvvw1feaYiOshtzW
Lm/OCoQGFEJFLNvi3Tp46iYkW5Zu+NDg6YIM4q+mLXY8z2cjioJS2dHNNF0ZzKZ7
Ij/TNu7hqmRn2ChFYPDyTErrFLYIRSI9aFZefW+BF+Su2QlW0nACba8ZeGGm4MA1
+00mQCnBdStxxPL/kXUd5ZJVwiGkKLh0CZg3JolZPgXinMupsAE8CvPmIvf0BGGS
IRzsbSxG3EaOqsT34JD2amMpryVaxEGlaGg1e0WeFr0F6xLSQ53qmjerNfqWzbeJ
IXVn/y3+UBA9xV0TrlALxq9Pf3+FimnbtX0e28NyMAq0Ve3RTFyWIccOWk+fnliu
uUJRUSqIMqGZpFRw/f9iFDHTc+flqHF4OrAN6GG3K+QBvgfsMF1KzgGxcgGiTXab
cVfiBsdGAkmxGrzhAjaQ1HYyqL9Dh7LM0XxDWgHNvzFAHc8yXuSsFwGLeax/G7y5
/NXMj5iedLZlPLgGvGoq0oJJfAPvCeiEEyW4LBJ2GKuweHIneb0f7q69ExIJGagN
oRUJ8GQTzPYh2T35Vubkn/2mCvoiy7i3Tvkycc9eTPZf3MXZzIM3XQO1qz8IO4E3
HadRW9rCbNw/COYTA/dYg7ZyeCdw9izbUDxAix+Iz+2j/C+phx6xY9C7vH8N+6ek
rJCeiBysKtQUDy9YRqcCyoLLf04ErYtoLKCxYx6W6wa9DaNGWRvCDZ5vbgI/ADWo
Fb8Dt0T2YlRXIEi/KpaX6HnKUjze37ftd/X2j6xYQW5vWfQeudr5h3/OYxhMJ5sk
oggIsm14JLJvFjKacwO2WhAIzYJqOr34OcpxAPDT08FPjX5ujYEx/RCdL9xzfGpx
Awwr702z9NGVofUK0oioL7TL2S9kFwnRlg81Oqe8+/6+ahx5iQ+7rBXSeLVfl6Pj
4VGPcUdRXCS81XL+IGF3wlveSGl542A0EE9EGCgTh9hOJokYuFfS4fd2T9kLoUVe
UyvlZ797tp+QwfCTZtj8P7lKd2yvwf7VVF54moGG5fHYobG/r8dczoFP9izztZFV
CzaX6rOtbqTcgaZBBfDF9XnHxrSuxkz0/yjUzO0o4sLH5C+YgXurYbIZFj3qi1f+
Ort5FiNMHFRv97JeLGeczF6WGRwUcQmxeW5os02PXeOqddsXUc/5QtRHLwK4vR8G
zX4xnBXe818Di5D4rRUYRQdPEj8Vy/ASL7iU1DcvZSWc+hEyJ30SfQMqwGXjY95j
i5bHCm7tULxXJyOrniKAu8AWfP1Olh4WLyexIOIf0qk8DZs/XMwRsueC9JTdSP3e
c9iC3ciIL0tIbsQBcMfccGhGrazdTo8lFRfrtrV4lGvSJRrjWOGE1i8DV6l+8IFJ
q9x6X+d4mAQKTlYasMmxxLC1CwFgTZ+ZayXlTMMmcZ7Ckj3yTqeABax0REtSl9Cr
OH5mKhFDbYQr8tYEOkJ1eTjw0z4noIj+mQggmtoZ1UkShE/bgIE4cnntqn3DIu1f
Nx5KUbOoVzOCHwtEobJZd3iQdtKPMS4D3PKbkM6hMSlq1hW8ZlYqXDby7fRfFcx6
PJXeQOWQju/rX0WLcICV4WTlGVWenzs8hSDalWHs/HZihI7jGsqk0MjHgT8rnXyi
Xg2Qz5zL16rGFzW+Dy4+dOsoOucaw98CXT/sgx6UXI7daWcwR0lsHzXTFehbpz8G
Dh+0ISWE8+3/YaqOI/Ny+5XorKPSx0AXdp06BPJMGm+hW8T/Wqu2Mn25ajd9u4qZ
9WxGHxeSpwo3HPl2tyyggcOuByuYCE+uohKpIjybIwWZcge6JZMCuN7ZXRrXLn34
mJcg71FuJuMVZq2mkV8wgidkE2SB/CULvJj8XY59GHmNcOZ6DvsWj1KaKg9OoKYJ
x5eisRKb9rxGPOHylObyPCswgdPM/jO/NGPcAJYZq/5FgH0CwWcLRmRQA4i+WPxw
b0vPnGe5+ecNGrf+zOb/SS36GzDCogPJnbQ3Hq09Q9AWlBP5ITfti+/w4BcTbi9w
lNQg1v8nY5XtLlfGexm7YhnA/P1s+gg4Z4UsblSNQIhtiz6QrpamL/UhD0BrLt2r
wkHudWsMsO5vDOzuXqD+82gDL8CsEUIrzIdcshu2PYtMVe5fYwLiiD8kiat2rnnZ
9WEnrCkkdqWMURlhT/EcxeBsp7VQQeCnap/XgXkNvkDl7/m4eIXMMJhcN7xcrEqS
saFfQjD7ARyP6SqfKq6+D4H84dWpfHP4mDP9D5T10WwGZ2ugNiTawJqn3UWpCum9
C1RsWgCqVQfeVFZc0+seOq2hsCVjQOcd9t2b1kOJvsDkn7+tG8bWo6HPtQY734tL
YBBJrjUViYOJXCHCXf6FTUIAsJJ8mKdSzwiPC55AVJoZQ6JXaPAzMFTLYgnHQ01I
Devq16IIK39Tadh7We+CFtLfnHyd+uJpJOez7ftaQOY=
`protect END_PROTECTED
