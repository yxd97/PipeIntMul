`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVyasrYpvY+mzzATYORUCbtYT5Iac4tq5FDOJ2B6SJXx/iXfqYw/O2RC/8Jcs0wy
5pVjFVehSxcKaH4ZHSbxwjGXFitaL5KPofuXWpXOtrVwj6XAIK1ALgG3z7UwsDtP
fouJFA5pvBMRuNk2JkiE13tqvbrggOiRcqyevDmhNgDM/VckIxFZqPaE0ftnqN2s
e9gPYsGavhjBlgACHJFuRllG1dtnvrSR3fkgPHfyXlgh6Yjz+kuldLmxuFV0KoBm
wXer45kwYMlYcnKPe4ELAL5q2LIuAEn6KZ7O+/UdJzQh2r0hrmBXDbvXe4/+MX/J
p1ITXusTMXu3O85ybpRO3VB9RPy06Qzlsw801ZWADyfpo9AiTXcUpBrO1wPOIS3X
KS176qh/HZADLGLrgBepT/Rh3ck9muvYggD0j0xhp/TGrF/CzDg/lxlUMY0L1MVc
aZRXAe0jGNAhxC7dCZLrkWVBUrqg1OmzeHO2PWGiOwgcAMYJePnKrjW7+VFNKt7g
gNxSJPJ9QQTv62n0pgi4KE/vBNazUi5ddf3g6zT4ev4m7Up+pjmG+Cv4pTI2QXOi
dW+4Jm/GNRpnPBv0rj8btNtWIKoFIeCXWxx/2lnOqn7glNcWT5Hs2Jr+J94JYvyz
SbbqP06rheZgeW1kVyJVikikhUL9fhgVYgdrPZZIPW23C8OHXV7PFa2hi3pqa7wO
9q6N/ADe/M/UnWxr+tyHJM/h60wgH9IU7hNUUNIS4xEs5ckd2xrE2QsLo8ib4OET
lKVFpAuc+Wg7vmGRzzmIXJvgDopvg0iN/2TQHbydgoRBxNNUK3IbvQSOFpcGeLQv
7gu5muHjwlDhTNOnlazlS7r3AS75g6enVbzObCDPn0KpqaAa8JOprHTKZB9FNN85
OnAGVv8sxltTSNgs4PBqjmGnEs8zks+flvxjEI7z29Uo7iaMzSlz1OSeTS/kQiq/
`protect END_PROTECTED
