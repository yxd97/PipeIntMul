`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
965Ihu5RdZblC6TnZxeewHHtxtpIbXJHif23ptBJGQi/g4VHZWG1SDOu+LquNQs8
pho/eaiZ4WDO9YRS8h0Es0l6Bkr4uiUbDEjOMX/BZq5ygfiMb+OYaX2iNzQBnZuh
loN5D0ObkAvAb5y4A+AVIKAHWn2YpTFubXzKXadAOTy1sYMmdCWq5xqyBLy/WKxN
V7E7VC/MSKKPrCvZSkki1GcAQJLCeL8DsTkOjpG206Wlxcqjh/r/Q1g4HwWhSpur
YjaxuBLmOYbYSFIebGdwmcq9o9W+oOEqJpwcibKYfIJeosiC1bhzw/jSy4kPt5PT
Bg18Xz+R7bKg9mrdf8VznYc4hxN0/zduMJ5+BKEiutoteuDb8MkaA91FJTaf/3mA
F/DzkAZpV0nVKt6T7E2loLk89gP2z6W4Wfcw5Vcq8Qn83umLUYbkijJ14UJCSRyO
`protect END_PROTECTED
