`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w3lx7eMHWXTKpCWTzVC9+j9tHN5MIXwTPOGuMPjVz7+LXckn9leX/Lv3HPtbNVEe
tb96TLkI4FZTexFyd1lVZ7WBYkfZAx6G3ObdPj+LGG77gWs1muAyfxlXSWDuq1Mm
GZEINrYhDwQ6xjL3Hi8pJ0orNUcNsyJ+lHVcNhrloG++nykhayZQ+R6OAktdwUhv
7cN3pe70uJ4vbk5axF9VFbvjQWZCToEUd5+RvqeNJ96FMhRD+MES8Boono9y+WWs
RVfvtMKwiu+mOOhY5NmC+b43eIXR217EHqdPUptsaGzTFbbnAFmLrU7cB45DMrTJ
tZKf/3WvH3sIxDXFOXT64f/sz5qAHOmAD9lHgkw03wOqOaQzDVH6BRKP10HuLQ50
1xZmn4mHTJVd+7upj2rwX3maGisNfZIyU/OrlcbbQX0vr0XzV42eWahhUHrYwkM2
`protect END_PROTECTED
