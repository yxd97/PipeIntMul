`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MSft6e1MmGrzFgcDc+xxoIiEZOPcgkMH5F1zRkpVwuuTNw9fAiD1Mb1/l2ag3e7q
MDjaVNp5I7Zzqi84RSlCqcVPnEm+hx2E4pHGQoZFl6iXKtsfZYSQPk+yKMuEqP1D
hPOoG0Ndi3RT1bCpGtMyKKJhGAkVcAkeRM13PixhwDmuHPlLChhSYPQePPoxNxi3
7xmBhFe+d81IEVsa52Ug8H0ZL3BMCbGTe+Zt4dRS+c7AnmYdCCyfMdwQipUKfsNQ
tjX1KcllYedAianlWTLuh93OPLl6ePY31dAJMygYk1N+rkqNONYnHnZF27ZxPZfr
wdleNC+q1JHe/pId3Wv82SfDf1AkWSFCgRht1T7JpfJgB/JVugv2/Mn09FO2P6Wo
cwV+2hl8NhFOpC+evKPUtuT+gLxOcUqTkt34BCvIbcEm9NrqMHUhO7FNJqrCdebV
`protect END_PROTECTED
