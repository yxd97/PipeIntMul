`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DXd1VoYJlL8rJizTUvVHP6ko2LCh5RFw9WHwre6np3cNsAThuzX6NHr8QKD97Gg1
g9seG7YltmVG38Wp7Zemdfq/fvNFPUDLl4fKSaKONfRHV4iCQlwA40qdCtFuMIki
76rvhV3hh77Ke8u2kjMJIw9HNxYCItUMYgarM2sKRMUJl5vkqKogYSl3ka7PF28C
SKSDMXJ2xYKDCeExlV/0mBH4PxDesuV9JHgu5uytwV5RQzyfzrko9bt59gORPw8t
S5CekRJt4PNalwprKuzT/VZdy7usE8YHbZZmUs5QOB8=
`protect END_PROTECTED
