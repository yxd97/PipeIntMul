`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fSWAVD+ukiBOVM9hvM2zkfuUYDuIvmEsxQ/8HwmQ49zO8D4wi1pJuf6V2VKmG8Es
iq2nQnMRE4pYOWBCCN4BcqgyEAtF1rZsR3lvWI5oZ/dAEVE/STraQrZF9IocW5qS
4+bojZTk0pcYUFkU4uRGdM5I4EhzinyRDMhYqZQCG8lhVdUhjCA4rnBFnmGI0yOJ
k79WiyEgADinXrLBhtREAs0wb9iECrrVAaulH1b83yo3KTOwaw7g8MBwcccXSptc
7iWZuLuQ37zQ1ptTHn/r+f+TBtYqyuNSTAL59ElQt1I91QzTscrXuVIhevezHeXd
28pwwA/yqLbDCjXBm97YF9uvbY+KDmrkVN9/2GotdUrnatpwM2evjCRXGbYlM9Oq
s1IGo3WsA8QcP+Yy+D21zw5W5fQsHpmfu99cTqgDPBEZqBxdLiJ5jB43JsyJfseU
NMPZhy+2q34tpTdBkzPO2AvtO2YwocnFVYbLoV5A+0smvglWtkR005OhuTrQyMKt
N+Y7fRHMZ60BFROjw3l/4xIkWRovdv1g8RO6qfaXDjMkEKdJSBWJpajBXOYWQHgc
jdEmaYFC1zx3JqZtFw6YNhJW7iuY7pRbfLuI6OXQ98eTrdgwganr+ocDZRfllZls
seRBBmf+pPlNpE7lUqOzNXezMN/B9BUYcnDbHOtUOUm5psfONG7kJrbkYsPDgy57
VhbRoQTV3WKfwZij5Ue06+VX7UAKuuYc0XYhQOv57vUcPpIlD0c8uKL6uqNhadwl
nh34hAfkMaYXu9lXBHDT3EG1Ti2sgUz11OzprMngFl9XxvRcjRxOcrgy5d9dgMMz
71Gqs0hWx7f24zF8aDEt7ndzcM5hc3BNQ5tN31NPzvDmUb5e8RsCdEooQJqDYdCH
SrHuymANI33y1pEacDmsq1W/0bUAiAIbFgeRAN6Vh+bLjCUsBVYjPJ+PiiEdi8pK
1wPW4Xk0enFHRueu/Rx5X/kQz11dsWWwm7NMMiSAeP2bDv4b/Qiz2Jbbj6OImCrk
vdLfzU4gPRB0BMSvK+ICPDnp+z+DtZtXgqpNqrAurrpZTafAm+KDeqgmyJAoHJqq
XaDf5ErpF10EvLirKd6xHF6IzaL0SyTDrtuUXAN5TI2FmB0546qgzRX7X4IUCsT4
TUCthIoq/YdqdtpiOgRJozJq39wZkrqoO2UPEX2vt4xltD7UyT6yqf1VOu6dEPUN
Ud7Dbrjc1mQ6p9WPfM0KuI7KxuupRM5gfNA1NHfUCgH24MT3tQ3STk7vqy/DlQCU
`protect END_PROTECTED
