`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SU6Y6AJT0Z7NloZBgwpOvzBM5Zrd+IBFL3PdBaa9i4iT3hBIPK3PxBaM/01D0z17
j3yX0rYxB9GrN/2kmZvO8kL6Ut2zGYgzeUhc9GyncckUZRXWNXT5oZYv/UPZo3r5
mLLCiQHhBdNKSS6kDJdVlsZhvUmd6KVL0o5BJB7d1DHp8LNsOC2DYZeLs1CjkL0H
89hz78dhVkuXebTWX9IJPxOH8fXWGaYjmdQOqIvJ+Verc08LUdFOo+GbPgSdsxeh
6bMDUZg5EpDmr1Hf05ts3/oHiJUMyGrwrfJSYfL7fkQDsOfKNubfyS9BYDsj3hb6
XbyGxSbGn00L2hqe0TLX4p8xIDeV7NfuGfKGrK6TNDMcgWX7izG6xFOqHWKRTom3
3IhpcVI/FLIRNxd/cCm31q6ntowa976CF4a3MDrwUXbbPPtz8UZZbI/AonQ1TZV1
M3e6PrDmzPXss2mXhVEHvfVZcylCuQrGfyf+j6dNgp6xzb7jIx5GElwcdD1qg/Gy
iazTLqpGefuVRJHEr935zW0E+YgNpHnNv3oiyQqrn3Sh+q0/I72/g9KSF8yAH3En
XBJ2893g23jKX1QYM2bmpshWR4VhE2QFJffGxBVedBFXKaCp2ioI8Lbp76Y8siLc
`protect END_PROTECTED
