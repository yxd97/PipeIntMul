`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B+vFYFLaxp29i0dArPun0UJZVpnEsAuicHXWXa48CdsZEO4kmNVF+hFWZQeXVOqY
IHSJIie39Nc3UchvddritjVfKZoSXaovoq+eHFVxkNbw2hwUWFYLnx5NP1xkoRbf
RqUok3ZMbaqd1GHyHZWarJMh6BkrMVZ3zfOq495dnAbr49AHgt2KGiCgsex/PFYI
muY23h+p/G93boNBbNM7Trw0yRpLVZgzPIsY4j250Ut5HsHS7TKVisV3/ftqXheF
ktCAdSQBjDRWkqEXZMrwfxvGsRjtlCOlr8bkwENmefz/IwBp9K1mOLX04FxubDqH
akUazue0RF21XyyWyEq7SAWXYd/fhXsp7wfIRidnrUMUZ9nmkTDTtP813TP+d919
ZWPxDYZf841wham55J0hYGKcPEhZLkFpPiXICF7SZBtdtJRSilnuGH6Rj435WnHq
zf/fC3YYDQCgccu8eqDAXkoiXpt4W8ANX7GzhXjb++197lafBVc2THOgaHy4nmjp
9LfK+x1qwcT2hIv9iqfKjCeDyiUuKEv6GfPfgQuzRSeF8AUZ/+8Ks3jfR5BtezZi
qfRqTilrCcv30vdRHEn5BQ==
`protect END_PROTECTED
