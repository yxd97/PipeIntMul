`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZhgkRNYkOnbboIAvAKBZ+GByf2rOtbpl/rAtmiMDK/I7qAcAFt8aArc3JqAjInnm
jceaFo1BaINFVTxsh+AkRFxXRDwnr2jtvalqBk+rZBG8VnuC4tGWgOOwt/FZiI5R
uSlCsX6Lkf6p3EDZpN/Lz4zVPJaPFkTAFf9fRHeRH6UXlH+XP8YL+Q41b5xn7uLm
OaAZoFSNwfFSFfx1hPuKO5ORVjUwyE+9Jlowj/I7etk4/IpUhDS6V59wsTliUjIv
dx/McxSQugDGRp1uJkwIww==
`protect END_PROTECTED
