`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tm+orQQF39FS68w2QcdNAOixQ1elzoGJGBCry1O6q7IS8hOG4XQMOxBHZ6H9Hjul
viKEduydsWv2sDaeAhjWYA5h/YmZlKtQic4Q4VpfoDFQaOhnfKmFfNLxx/I+RgLA
zmcEXoFTy8pcbDEpVX4oYYLpPiAatu5U9KXSWcixfA3Aa3QnaDcIbUhbBzPkUmRE
8HjF7Svn0ICL7i0K/gdhADegAvhq6Xs2vNBFYkdeHWN4Z7dRmZSK8+beyY1zhBUY
WHaqA6Ncy8fUkusqMNRLUEDFUmPCQ0tCdmQRQCMhpI3kMQHPY2C3b8Ww1YQXFD96
kDN0bzR44AaOD7O8h+oLNg==
`protect END_PROTECTED
