`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v1DmmtgkH1gD0arAEVkSPKnK00CxqS0lhPEftV/xmlQwFd4sWY8Vu5MA6s6eip8+
lHMgUE6/4gZRIr7CH+9LhO437IZXPhRsVVbGyoHKwetvRr8ZmMvoRGtN7vOcvcqM
dI/iVhhX3kKzY1wDoS6RXR3eScETIht9QiqW/o4mkqIi0Y0aBmhr1qmtLmmZa3x5
CUBUeiWlk0R+8DkUZ24/HbhgJaP6iuxxxtqxxMDdUV/ItOXGw5N6wr/bGl016P/W
Y5XmbUNBvY4RwYVFH3MysTsgeZuFSVMWMehj6rYQo4q4PHIDfrDTDAHaKt+ofkFq
XM4qdzyUmM1YfHzkyzSH4cNmgHul4//V7DPoFGOUUTEF/OkUVhWbtQWT0YMFCaM0
O7h5qrD2VdX934802e7L/INuK2Qm0kLhbmRLXEP6+tAStS7EB8U7EueEhElAd74E
oY7MBZHvYS0gCNygHZv3BXuOJqLopEM04tpc07mh1WYjKAqzvlvfNUgCBuarAAe/
VumObBSaChZVE9FQFJfpA/D3TKHJCZ1KGHmG3dxbdKg598LTGLbeThqvG2vNtRvl
DNTgdq0x31QT/oVZ9yKdKkQre4b43qJ35G040I67Vh1098MRbVspPPTsTAnndNzI
rM19m+4h710GpPONBU+Fc5DE0l+1JejdWkbAM65TdboG/5KXK93Sel3iKv9ZD9pU
/YiA/xspx1L+4HlMKrbB1Y/1SpikVzu6+x+5mrzlzqJ/+tZkpFTpBSPn1RFCq/vJ
rctTA2rp6rv10D2/wxL1uIegLXu5VZopLyJolEYOwZO796Tu4XcaZhr32YfXqxB5
V4BFabig6PxF5BV4zWiHHJEZvGJx9WAMjG38RKwt6V6/CDId/GhABxaWrENKvGz6
jLV+8ddP1bkfd/mBkAWlwyB8SCavOJih1qbA8LmD9t3GTOot5qCDR2w4s8iT0GB9
qCpcmkxGlONT4LYtVbKAUohp52ox60wq5A0HKIyv0FMlhnLRmhQsK98JKhANsV3/
H4xztsrOBcQHLgR7y0rpDHoq8rUqt5hc6R6bFsN98cCyuFGZi469GkjjN5pL2v3B
VnbTE9+toQRnVtkqEKLXCnGOdkYqAAnoBEiwJtvOchy6YXNO4XlA1i23Df5p4CQJ
6PrCT+bz61pH1wue0YLF4bbPrppJ8+ipLzOaMCVcjitDgbsqPNuhmXeHciUZGuh/
bPiyAZdWfR3/4o9sPnTneOjpF071xYBhZVfX48sBqpUoCh1ZkouAycXIuMriXZhm
J0q2xO2RZlzdlWaZjvWwyTNNOB3MPu8vAzApl1/kUMUFGW3pafO2+Qt85B7QMrAg
XCmTVfU1ALgT2vN8MQJ/dXRNRYa+Q6WCl9WxB2wqXXH96b1yEtTgRtkxJJtUm7gI
SlKSqIKza57uXTTvPJw1TPcJ0vx3Y0VMSFD8PpLPiBFSgkcEPL69ITNq74hf6KqU
vFAnQRMc2TS0Pbw+92i6LSO3cCMeX0yNdq9gkeshvqRdzT12db0siCwslfw/basa
Vr+zxafRLDTRZqWUUNcmIEWyFm33p0li4Bff+vOkSiMDwTWGgHZkV84VnbVer2/Z
XKfiIJO0Jx7XFvLAa0kUwdACuKO22T8lc63yRV1byZZhyefLh5WpN7+D3f5Htxf9
1130j44GWuAWSjxoyIZS7G8U738ZNfkiHU29pdxZteZxTSZGsAdR/QKLYu4SFeMC
3Z5py1YW2LRQ4Gn2HReZErZAND3T5+4M0vPnSoUra1FYuRf1ztub2kaUfuNAP7u/
CzpW5rdHJPzhQPT0lyp+z9eEhgl3646rLAPZ3pFVDb0lKkTHS1/5R5nhgippaMS2
ILYodlmY73GlGB0olbhDQgPevgHLg3YOkv0UvFhT2ZgigebEsrRqwPWpfB1scHA4
fuwRQMxGkwTwZzvDFMzsK7DONp46hFYQ9GZbgTnekZDJZmBCfTbhxGrrlZJ3T/rF
/UdhgNlSKVNBh+DtvOilhkU950f0ljhVMpMsBD1MkB10BCQKbSF3Wp5scoSYFcbR
s8wz6NXXJMjO7bX3216Js7bOd3BwNEUlgPbZ2wqncXVFtdXAC8I9z8vzX/k/eOqT
1mYfdhi8UYrIiM9/fXwqBY1NfzYHGo4s3zCJGXTnz/SgB55NrZFNvf3B2wZzjhSi
vzR0AZSmUdMkF58rFTw5htrbY8XTXMY4G2r+lyVlBvZrcHv6Uqne6K2jkS5cEocQ
fLpJ5ffaIYO+poQESU4G9GSD8Z1O80naQGFxhWz5nTqSQOxf70t/hsTks1hSj8of
IgL6E8xWtk2F7FiCrIiMFcQHwe4xvtLc2y5+fh9QQeVXS8NPnQAKUVPV9ro0k9tB
efOShNNaWh71dU9WMLBrFgKTe9DumxAWjZzPdGrSb9HebsxsU1LEbrf9OMHs/d7M
gCgQyiNkMnz/yis/Fkl1a5t6+bytLHE4swQWt3/Tvk4/iHysp6zQaoQoSMp2f40p
wS/MdkAstlfgenHdyCiSwgz+WR7FLIi5Nxh46mOnAew7FadJGYe5WyHMSd3Yojox
aCw1aid7Zrm0yi06gu0O4Jnp55BQGn+SOM+f1k1QZ2yDg6Tmf9UdIDXymlI9y0yq
3oAsKsIf206sMWrUg1Gkzmc/UIsB3YST8molYG/g2tI/bz88EfYwFEERCeuAxjMO
YNRSupLtjKC6Ck25NDv5DjfA9JnmmvU6hHp7PUDkEOluPV2JSlOQAau+HUJ1eHBh
o7kFgc0M5kdtoI/kbUsyfcU8yrpD8KdvpkLAmZjTD0Rlznrng3EBhDzOaXO7Omas
VzKTsAMLVwo8XI4Q3PYHQRS3X+myXe+nJ0wsd0Kpw3Xon7Q+rT5MqgRi+1L1jNVf
Tr0//8pglJjE+jKyQS3GTUXIkGnOzBp/zY22nZZ2iTGQbJKPZ4ZiUdofBoimk3MA
y51XuiZQBa5gBqcpb4kOOUcLCS7gq6lwjkMup7xJYT1VBqwYbU8vmzlNGik6Cbr+
C+BuIdBQ4HFHIo9ZQKqudIAxxsBfY1Sybq2vmK8MAI0MWhiwHzZcpSIiCosCozqI
nIopBwDfabec4OutqWrSc1ZH7linSsaIZzkEVNyU/0izHwQeKgTuhNzxD+ZacCqQ
AyXokeFmOkm23ryciKhbBL431hsZrDJzlvR+BYXWJ97VgwCSEaq03jhkbb7yInbp
pv6W8h8hR2vNdC0aplI5MkmlKhL0ELteNa8YfgAbSG+0nIVDfyT+4acHBKbk0mjF
aAHTGS6vPp4Vux7u340XwQv3LX0rb7uv4EzWgBE4DhE56alUSvThNU0ef3VK6nSL
yWsihYVrnLVJKfBPcQgFSfrppPWXQTACyPHyHVWuEqs8PylI7Cy1IOdZNtqbxjRZ
cVHbP1uv9gl2GNuiyero4rLL0JStRn1a16YZ02W8nnHW/ajvKQt2Ay3mbUIGiMcq
ZnZUollnv4pl1vZHabpRkvd+y0G7l0Ks0LYtWFtbqBhkMJKbukeseNis56UadD77
EK0X7QF/dZxUTfqPRLvXhZOOxIz6IP8y60V3X9vlk80RcKPnEZdTYC1gQCIKHmkZ
Z7mlcZqQQIGXl5FjPwtpRglHmRmCxsIZXXae5zsp2+Xr3riUyoqNSXR+rDIBDyuz
/OVO+OEc+DaXNIivpbcUnq9kvab+6+TvIvv4KbKJGVdL3CDb07v7LUNSZpLeAFj0
7raiJmgDNwFvRonCwEwRDj4zhcgj6PC9qB7q6fAPr80VVcxCW6TmAwBPk6t2Q20B
Ly8bnD/LbPXOz5LRja5dz1R+b47lKdhp/ZM4COTA2UGjotA1SksI/B5O72HG3lZJ
VKQ+KXk354y6s3HF2Khi+h0xWVShvr8KD28n7cMAQF3g5mLSQXOPwc5k1C0+7vkz
hi+dxzRV40u+bAya8KoBhZdHuGuNO1gDapS5Q2sBtcJtGPIwf43ITiVkq8qSgfXY
94x52uusHSkPhB8cloZs7f5Igvv3eKXxxrukDKdJ7934mXq3FcwCx7Xm9o1yK1Sd
gr2hmcxNCGtV+IHLqvkohcp2rpGhubYoqCQCoZUubBe7+spoH/JZCoYHUmMrORI/
v7jFgb1ldoVZF4hBiktNoOPzKOjBQEBTt+4F5mb5x/EPMrecLhp0gDU/dBUmFBld
Uh0POWhf/gTqFDIy3I3C5AIUjJEI1qQlCOq84kk2YKN/b/h3VjidVghvMeNgEvpM
0zkFI82Qyd8Ik6YRfHfA4ffQfyZwIyCrYs7TkI7JrUsJqIoZow0GshzZqaxWFX8U
G28d2QTKXAR8sKV1b6y4PkV5QtB7/bwyHiBP90EavXBiyRiUPSr3bd++WoSMCHCU
/zS8paRa92B5ZuD32SAks+EvPzSTOTKt+1eb6FQo76tGnUmuTugkRtjn14ssK94S
qEnkehcXZh0mH26I0QRaFO+1uyIDF9Ea+JGptSMH7Ol/dduFfRH8t9BWe7P0AXUO
Bxw+HK4T2rEUMQul17y9ZxO2xzGdvIxgBIj81yvD5RCWYSMyiZwGh0W5VFTbcK9s
Jm1KK1g0Xab9ql/osIVKhiw5a2jVHZkMSNwg/4Uzlp9zalXij6hfCIOhCH5Xd7KL
2jKzTxoLLTBCLyANahsH32zKl1rBxJ7nxNKofL4eUAul6LAYP8TCF6W87/G57l3c
M4VxYAuLSnlh4EVVvtvyqX5YBLxqGr/JJLYMjlFHCZ15em9aBUl4cn96JC81rfDu
KnjoI4Lrme4f89N/tEzV2zbyHewXHSlfRsQgF/ZaEQ0am9NIgh0Kmr7d9tSHoR9V
t6uEWFHZfRWXx7nyTIX1391L6DFTmdGDd5D3X3kTSVGkiTwP1p8WvAVxMV++uDx+
ZQtwEfY/j3JTbd7eGs5AAfuK8DXrp2EMZg7dED9yicWHaqIEicEAtcmJbR7KvpfD
ngxfjaqth7zuROllXXV8fn8w6DIwYo7QSOFJYENx0rzfeB8BGmC+Rw47ZILAlZrB
04ujxGJms6yqWIrNUk0nyhtO86A7ItgQFfoU1icCA7+WhdZXrrVuLX5rBCYdbcU+
MrdB0DxlMpHPQtBd6+Re/+Qh4JynZ9Kxr65CM480qCWM4TvKfqKOKoI1z6I1Staq
LWfdZj9ESbnSbXRD/8JBNwf/FSN5J7+XZguJEII6sBjHbW3KTt80ggipZjE28z86
qT9iguSut402/dtW4YjMQvf1RMQiyts5ZIkuTFq4T+l1ilBOf7dkPEf1MTWPMKyY
xokLgC0V5T/T0OJHMc5WZ8YrVrMyaZWG3Nbxgj8la1EQJOgBTqW7R2YYuhsV/XmI
ohvbMjK33bhm9meEF6b5T/zi+/OFdGaz6t88YQTgX4mvxGwIVkcX2Vagc58MfcI+
fEZLfUSKtFl+X9bhNRawYvG7OnOdkmiXdbQn4Aw89w8VCeKYCaX5wVjJUdZAS5i2
/j39b1guCtyn+9YY3aP9qDKmddscu4GCuDtJTVnZMbCR1WeIt5uqzwrS/exDSax0
8jV4U6ncWkL+LxvP1mFmCvOAMEeUqu7OPzI+TVgihilXSta22O9tQlEJGhlj+I8i
q+CvI/3ZCbn92xAweyiTRPuFV0XdYeFtWBZ2XGt94DGDj7MLHsWukP93GYijVwPM
pFqSGpHCOnHXOpEWNH3PPpVcfCd0nWlBb5xbqsshgQlnLqj47D6kNLxRJ2hg7ZPA
cYm3K9dD4ItixjIQz7H6+dKUqrVejFXzavtXf6F+eWcj5qZLKGbCGa+kCKgkndrk
xK7h4pye2ePhyyonYZq7bECMoGb9IlqtpwQBUzixiN7L4o4K5kkLGL4LvupDv8gA
7G1ISPx0sqPGaJGnidydVAQAKnuqnNohVzbqheTVqc/vv7LqkIMpVdQQ0fyTrEDf
W1LMoTiUmbdb61pnmIxJQMEeizjXh7WzFSjuCbSwMoVkQrvTzW4F0e8cYWtdcfAY
hWv0ccmlHRAhqF4XENHkj1WMGIavSNRBykoenLjoKsjdtrfl7YMuGJFYjkIUx5ot
1OL0up2ja9OrfGIhbKCFStrg+BYbkyn9gCQPIrl5OPyL1vyyYNqR2Wkeoxh9D+gX
meqV5GsuZTK2ommLMH54h5KAOb9CWf4bTB9/hbF/wcL0FyQ3dGjvt5+uxEiV1edk
/1qPAgI1E6OXNIGHh0VLP/HPlv94XbuhEg6zKEoY5J8L59K1oA1vYJI0I+Gzwhlr
k30RrMiEHpQYzgzzlK3sZpda9S4o5wBuspTuXQ4UMA7UqMmpfv9AvkgXfwRQfKLK
LK99CTCwatqHaPHQ52vJddiUMMCMUVZCoR3+bace1hfmsFUH7By2Jy7hcIJ7PssT
MtnYYCByvzX4lxPbizOJNoZ2VmlrWO/5EUFfrIvCnMb3/aaiTcSciMQq4N6m8kw4
kI1OuisgD5rEi6eX0Ky14O4xtay1r4d0UOruKOa1kiXTY1q9xiBksGycuHUBjNjM
Iv8SaPKGFJU0jW4s37Yj0J9UuCMDiH7ZYbP5ze5K7NaoD4mflvAaBE0V3eY2iXDB
2zU3LVqzk4c3Lr+pPR0iqrbvwRXRnb98DmBXL6GmNulUWIdKfSna4qA283A43CHR
JaK2ovD3mYIr8wFJ6C3tZnJc2u5Kj33l3qbwXfpSRxQuwTFTItytbtDZ/7W5PL5D
iiRhaPUt16+Syx7xrWGQHrE3cFWtTPPaBNjunnnltkjnvvyu8Tg5VHSksLv577r+
dA+gFLdPAkWKnCpr+mYrfFNJxPPdph8w3mIX0dZpVs49kKhizfFbZl+SHCbZWZle
uthIFuqY7pr3yuF3sLzI2+WU8Eobar80Zcy3vcsh92xcY/4e7VXOwT+8iShoPA0c
W/bbz4uHeUs72t2gtT64MUdhpE0c3z24Jsb9Nrt780a3TEgfdX3EuLTfms49xzkA
xBim/9c0fPDjuD7EkApnVy0f6F94CppnKOfQ9WGELJ6dtH4WkvP0/Ww6d4AlPgMr
n2Zgybc2CoJFs7WIPyZvw6d6J5fC/PeKBxMb89hqrTGJbqhQcd4RRbhEtQ6lQwKu
FAHuDAsrzQzbzVCjvSQIuHnxX/Sr8rf3Cip5ILo7ZueEuPlvRJuyXpUbDlzB6ePe
zNrX21X5N5GIyudbDhAWxEiFQJp34VWM9o8Q9DfLlb7Uis/OOX32BgPDdyURKbCr
HHyMzJKlYv1f1LrKPppUOCk2LFmBMUEMWym3g2HM+nQWsJbxzFn1T35Gx7WlfzKl
5IyLwGroZpTSrM3w0OxCYT8ZdM7frazGTWJJ7soJSRuqOfW/zOAtJN3yVmPLD5Gi
zy2XvPGDjjhRFSbnP/OE+Q/cSftwcVfUMLOa9zY8yZYuAu7X9gcNd8pie96IpClA
SIZ8fUArOC6KdO8cJ9C0z8hjcBVKhO7yPO4AxSBy0mpUQM8u8CbKrqxb8dCMkLBO
SL1zOsewU4+1FKd5bPkXRT6BBEkpVkRWffe9oDp7nbVAKVcIZqA6Keg6Oh49QCrs
Ly9CXCSFvwqOhDs2lZrBbkkmGmtfgVdXsGYM9q5am5naghWcjoGS6E1UQhXNLEck
erGMy8IfAS0+XL6Yw9bF4ZBuZvDeR3InnUPBM35j/ycI8jTIqmozHhs3Tn+DtkGq
4McNgnFRPvhvlKpNtM5QYryB8uBAwSPJ9rBQ0Go/6yT+GTHcT1r+XTvODnMNilgF
Z1gg2k5GOuNWniLBzezmKIbPpzEib/JSzlizUVFv4lj21Vo3EdAXdo3aFztHobbC
TD7zOSi4qYtq+EswHjiV4KJkCd2sTxXV5Q0JiL4rWZeAHjqHMTUSoeVTbqMD2dvq
kFXv99b67j2ICJQ2MF+YBo68Oq3+vUDrJpigDEp9KVFrt1QKAWAXglxCFuM6TCfj
JN2YTj1pg0KYsMspCdUgDVhtc1U7ORwDOXtTZSYdrIC9MT0HSpagxZs9/x3Bn8T3
FW+8hK0KeimacFa5cbcGd/hOofDszriIrVsn6RAlmH7Ur5RM08dIa6oQcRUKmkYV
bFoSYttm2QO5rOfXLMofD1xgPrgw2DONIJdV9e5NSgma+QlfrTCp96ozDg8bm3F3
LHhrG4wBAgDu5dYumEs9SjsOG37Zuwza4n43t4fnYzrBfY+1r2F56NPgUb5BTNut
fzYE9gOMNqYJ2l9ZKFyAALwvUNzXzjCmAMig27cSzUSZbYe1yq2R1RsI53ZqzSNX
jMImyh962wbcFArIoNZogfOGWtIuuiC4yVL+AuenJO0NPMnZXf4za3+PHxfooR4U
snIPas9Bk/EgYDVCYHs8bGPtJz1O54tahgAqcFxqsOOxiSQr38eQLsFc/HWcTiv2
XXv2Plb93SPd+PJ8jWOj5aTcTjQAKr/qKGdBrm0iAE5ji0M6N6rYs4LkGB3ZMpoy
JYkBZmpVJLNiIyAoBdM7T8ABW+YF2YnmvOxFPz5Oke1qRbGAO0DK8Zcd5OwdrBt7
DHYS/T0IW2wSmG479DjF/FOW29xSlen5rn+YVBTeGXGuxWJ1PbwJDfzqQiwjp0yi
SXNXAWqRWADAayC1OLrWlAYCAHIyPrHQznR0PJtSltal9BcmoiabJAVojM5BruEc
v04GLu2sFv6Tjk1vzPa7Ny1zP2+jHl+Hhbm/UUlwWBkftsJZzRZdp2XQhMbyP0/n
MXQjD/2T+m/F7MlHK1/PXwcCnm/Tx+a+TfT30QrPo0d6/aOafjj9oR0Fgq6pzhhi
CEbN63E/yM4sILRtmttRyon4nCNKAYBrBB1FaKDKkRE7xxmQyyegcaOoS/DtVAwS
zaQRGYoqcEEAfCfKsClwp7SGsDXtQyKcOCgvA/GUK0OPELXwjKravP2zG/IecJi/
1hYm1ZM8oz8qCaWUKh5wxGk7NUjRtJMIqtPa2BvDLG5eRsLQJI1Z2lkT4gihoXfP
O7LzJuIFj+i+1S0Sf/oLIG1loLTCoG4XcjcMORmXvs2YFoNw92mQCDzGey9Zrck+
VMw8H3woCYGKuX/lbXHSEssnWdYEM7erdyqKLLjlNeSdDPVLUg1IW0nYInBixvPw
/nJTuqLRKXF6++GKsWR8xLVtx8xdPEiWyQvV9tCysA/1sxF2pQjX40qN9GGU13ou
MR7noYLzA4uWhSXZYQTdv8aWtjImIcB1vRIefMEF/npKGHwHwFjUR95vZrEasFZJ
GAuS17Xpm8Qzcj4kZ1LCNzv/p9qDwDVYjZh2ePXVTQoTrMmLW1jyykUtzSRNCF77
HsqKFkAkC+jAqINWH4XD4auuH9o2+O7bQ5bXs0VZvV6IEjkZwpsVqehX+YpLx8iv
XhxKIJcmUUveky4kQ5pEPEXGVIj2J3ctkqABKlOBzhZ0CSwSkhxDtFjnfVq+IPc4
b3rBEhdvdnvLF53THZW9hGRAFLiAJ08D9DUioi+Ehij0i+bPmHxpC8EJV/c5VXt0
QQWvgiDs5o9Yv3U+D0FgackPtLuiyg+aiwjCi+ZIFIuuvj23PgWEdqz8PdiU4UbH
0kO8cm8vueL6rKQMZYR3xZeNvEvuuSJdMjxAkMMZ6ug9gxVCEvRqslDu+zEwCjw4
lYyfRnyWfprvmBpdMLsBodpGAdss4vmoLPUqTPeE9sdfyEMxjVRumCWyStA4sk2O
ZAGjha4AVgH9OxyWkDG3vOqDa5I90TCa1mR4vc4Tv610l5nxyjO1ppD5sTkTeVlR
gY9AstKn4hKFMLqaEaB7MTqsQux7br91wGu94QhxIQqOnkwoO1ds58QeLO+XuESv
lPTcQIDnNwNyHdrIQUcXnzdfFWIEi9TiFndlMB4Woub28jFJp+i+jB2A00JZp3V9
GpWYVVeH3itmEvicnNKfhKopCjE55T1WPJ6fF7V9hvUaqTI0z5M2vJ8V1n8aqlqZ
c7sEuvy8eJJG+aZmAjz40dp9EbShdh4fTpM89OmwqErn75ZIaWUloezzlu2WoVVa
O7VmxFRf86PYPwiQOaTHk62mwl0oiBZ5ZDqhcZqpHJU9M6jJEPpVNKaw7PnEm2rU
kR2hDibiAsxQfu35sXVvENtTfw0YUGeIxotpL4JA6844rjitcbHsT9m68C0ZrHgA
/PNxBL6cAe1xM4lQy9HNfzCHLZCJz7AEf8XYO23exxdp6JMm/XM1EFeReSoWW870
pIXJoy+EIqbTWCDJ7mtpzJXBJRrgFxJ+sIoW7J4UB5to7Ph9Gz1qj1vBbTjoWXFb
JpK2B0BN+7AxDMd1njBfCm3YhY9G6AZNpeSm+Ftorn4/2WciNS8aVmLAF2vd+CZp
PREH3sb10M1iUxjhSU/lyJrrby2cVDDjsyXpLTmnF21NzNZmtI+M3YWLUgWIlaM+
oEyXSusB0NqOoOJHObetjbOAUjctmZHHdlJEjrjYy1GIvLkSvrbREgD5F8O3Kj6M
XaK9ze7Pd0btEA30/OpJcqYTEZXBO6POTlXpdktWc3lHY/7rY5nJuBMtBbSeItXd
gzkrqYRFvFSWgB/flJOi+fgkzsHq+UEetHej8fxGolOAS1t02br/qk5KTBv2paq1
5iGMjjxvQEb+6kR3hWrccplJNUKePaBdol8QNKNhJlNaLTXNoLeVf0U1mAObyqzX
1GvAcHdh8Rr2Zvv9NRiTM+/Lzc2dqyO01iWm92C6efqGQk3zbyPdKGMznxd3VvkS
eMfpQJ7NTmnWDHV2LYQE2wTZsoms+wbARuRCbySeFRnCUUncBf0U5P0YDifFtS3a
kWS/0DMOJh3MXoo6wHYQQxuH0jqAYTmaxuk/078HQdgNPFoFSA2hIAKgs7rZ5of6
cXMTetN0btuJ7juimjr4h6XwsElHRoxIrjSvSwKCW7G+MZP7vTPjBGXgn9Jv19W6
COGjjNtP8fZbcLtrm33C2cWWiCoofo8+PVhn4sw6WFJluKIdUZalJErbTkBI0goG
xSggAGnXy3Y2DNsWJayLrvImSI2m3c1MfGE3+7xRLkoy3N4y+K6n8HX7bj7hV5oj
uRuCuDpG5DizwfZsOZ5kcg9PhdrYO4WFN/IVDVE5x358ud2j5pl9HEFTtsg9L/vz
pJCMeB06gk4p4RMakLU8IaIh4GdQUfWQxT2s/0ER9vVAi/kR0chBBh6z0LJatmqg
OjMc3tarkfE2ONrJumWcAkjpBxyw6wKPTAqj7Hzd190awopl4CQPlh3a+F9cj0/C
iWr9yCV8I38kstnLuLr/lSjpT0ltdtZ8WHVprGcaEvhXNWzX5gPYSgoI3EfZ+N1B
ZW9GYe3AdO0F1lkfLYZNWxjTKmAU0G8FBvVT8Ml49q0juRvCjCQFFEDvlSJ++dB/
p+tnYHCe8dHhBrHB0cRFsH5nvs5+b53mEETA1cJdHnEl3tYEoxVGJMMJtrokjVEF
0hP3alN0cCyouJQu7+Rb88/F3kz5P4auSquc8YXQhtReaGMP/Py9SpDEN4qyR6yd
3PHYNx74JsmmM+poczr0p70p0DjwoY4GV4A9ie1ErlgxnTqok6MjIiB4X2eEMnPk
YFJkt8Rksqq+0bRYepScDEzI2tEbkQ+qH9hisw2L0836rHfRbQSa3/ALw65M5vq4
88P7f646PM8ZgCk/duHePEEyH3kanC4EOTn8rypFfZjatONHi3cyXgV9n9KpPoK4
E/bNMNECjtyTakjqzByDXyVfUvjsvc7fX77xoZ8huNwa2h0ZpSzN2yjxeQRwjM4Z
yFa49oRsh6FRmLmy6BHojfYiFQrtCDNxU7ylAhQK7SO4tAQo/DwSv3ymwXDFPw5D
TUvpoll57MpoJW+WpVEHZ5VyLoVTn/b2zLlm6HgMTL5h0l3yfBfj1EwrIasmdlFL
Mg5PaO9UuvRxKQSkc7mRuGPxrORr3tRa7e0BE6/9e7knIAWpFOVolJc9UsQJNe4s
l4iEnwz+oHpem/AJz4ZjgAwT6l3lSs8DCQLcumHTqWEhgHf7VouwMsylmwH8Kjtw
9aJsreJ7jnlD0q8cWQH0lQAD4yIqKXI12YAyhxKzivQL3PcCVAJw6RCJ4uNOjZOc
HlKLIxXg4mzelIzkWe7/zYG/mC6OR0ZqqHNpViaP+NRXH4JbL7YQ1ICrPWNx2zn9
Rxxm3stzXPW7JPWjUG7qKlgnQpL/9Hz/mruv/sXttNZTlDd7wtfoWSfIHF/kNlXK
yetmjW/Zh9F/3wixkEuWCAEt/KSk79OagvLjLLVPa5pgiKq+lCxJeqlU09p5CndT
CR0tJE/OpUdcxB7yiUV4z6gegsHjD0M/hTKj9OAWWsg+JNVOsbGcyOX5xjsFSmOn
cMnKcHb4oP4Yx7EkOwIaY9dRp0apeaMDNNrtfQmZvjV3GxYyRzbN27GsmhDs4h41
h47PW8f2LQW/WMwPSYHB+1ZMQZROYOtYijwQWSfi1WDfuWZwnXLh84zq8OqXg58S
/e4BGgi/2fTF/RHbPY8yQvq1hTscv0vRuj31HIu1HgMS9jR/jkyY5QNNShZm7mdE
0djyTWbcI4gxhEUkSdlp2OOIzGks6ytAsICw+HZ+eaChIyjCxS3eXA0wMwFPb/8q
QhP7F15fPyV3i5N6XXL/E+mI5bgtSp3qO9lw7hNNoG4hlImrFCVusbOcgB2R8Dex
mXmTRYhnk8DE1O5+Ru6R8lmAZ9f1rvmx90Ijz00FqyiLnhGvbwjWDzKEb1JmSQ0h
HmOfgfAqww4aNC5qfoKsAh0GFC5nS9wk6peu+Mv678irxLgr0oABzkVSrv7rp7nh
TdB8iOX1A7tFBEp38BiJJ2L6Pa0Tmkjph7yOET1gg6aP8gB+Kd0QvGIG18unebph
ml9UdHYd+ltJH8f4x7OzdmZQDcIpnZMBAlTMRLsPpa6Hu4RSICxZovnRZr3b/T9i
lZPGDB0uEbMmgIlJw516p3ceyf2ouor9P6VuGhv0bqJvq3i617fCltaE6vnNOc61
KIezYuwVvTrH1w4MoYFVhN2Hq83a6GGQL3pewsOe6eiQ9kkwyFQs4dGtRR5KFWKm
m9yKpDEyqN43gsetEq4l6sM4hDf0AvAQyQpQNAOHqcyO4ZfXj+GZdDCN2dtaa+57
COPjTKeQNhyJtiq0bDM1+sQtpO3VVGbsQ2d8I62VYtUn7Jj2Y+v+xajkYB19n5KZ
pm3oSGO0w1HC5Ne6qKBdLgUa8VS/1dUTJR+Nm7zm6pnv2odgwzSDIzsqHnPj0zFK
Qd6G/HdAAyYP21Dj6qyCEVikwtluWE9eSVw/CIv0VcsdPkasi8w8mMlWjv97Yqd6
UtskXFeSzT2ymVGiQYck+l7+7HZbJ7M69kc4er6Ar/vboH/cPWRALfzHVQPwlFtP
TtXhp2Mb2Ab8H8JvQXqmkwE9HXnigtLxGVfMj6HrBghxt4HuTCGpOEbIteVgPu2u
Eq33OQhOy6cw3xafpfykbOtzzjUAuR90fMnpAVPWRXTSuc413G0/kam9rUw5Lz/W
lZ1uv/oWegkHvGFmv0yjpg/4HWvjJrJhoazj+Q2UmmGiCcgcSE64tuHdhoPyie8X
Bl7yW4B8jBRUuJ40rvk0hnT1vv5COQhLyvR0rutcE8rwa9HIzwXR3Frp9tcIRID5
mvvHyJF5glfrCtYv+FBlG+1KUP+zlx5K91uGrTbr2iDV/cettRAXnSdu4UXkMMol
90VCm22PkQH998fQAhCHYQ6gjA2LNWq3QO5CMNJk+IWJdNYG9nwfKYP4RfpxpBeN
u9Pc7NxJZ2feXEK00fQYrohQyHozm+iTZBRD7wHlcRoMsLigXI39dqzAmrPJczQ/
5zLc25uXQ0dS5+UcrMeNZ9aZWN75ae0aVFUr/gSSWdcPqyNR2sUyYFqg+UoK5Evz
Iy8xvv/lDdJ247eGWr31n/MGOkU/scAv4jYpYHOCUPIUofX1M634chZpL8dPbCgv
qxrIQQj7RkIwX0SE68gqAW+LXndbFsyBbyStBvJ7pr0YM9yPHOL/3yCB4YatIBvb
Ve+I9n+OuZqAOzwR2w1bs11ywi+QksVWzds/3r9g85yDuV01UiLDgQf1C9eRtcZn
P1oFml3xJ8182/T2BcpkqVur+Bae83sEuhhUjfRseoS+6cpAEHqt0HDdTSs/vJF2
gKrKvFBULSuFujR1fZDjBiNotH5VDM5InwnuROEFapkqs8EofRUKai9M5YFJkbh+
8ToRZQTucJb/PbOEmU4QB7VqMIUHUot5h9b/JsSzFXfus2yTtoG+6Dx2MQXb19Fy
BUzq7kEXaHvVyBhNZMeO17EQBLAXX9hLqt5yVvz+s7hq2c6KUoW/cCZSqs5jMhHD
qwokwiINzrjqqH6qNVT2FzyE/wh+uojvk3oNn7Yn0DMg1LusPZVJKq8EoRvFRtSX
n/oQ5NDC4TRnYVahn0+ZtA7k+NuUJ6v0PRJeWu84U7kOs3LncYQwxnrToWMYQtdW
3rg6jt1kvGOs8+DPRtpkHDNoZd5hdQKzLWdyCKrx6UTmXuEoYBs5FAiSvSf0PTQf
MU/6nsydF6Gq9aixmIWPLYs0dQ0QJm75aGRd4UkkjW4RyD6EUdsVn7tIRD9fMxYV
d68lt0CbWO3mgw5bpsZha78oWSSBDbzc4DPZxJXKylrGZvsThR5uX6AqgQ6jhIkH
s08+Jn4e8LWKx1+sZRhNJzyWFOvACZt2Qrbx6/fDpWHgaHePO1QstYONfeWhYShv
Ovh5zms5GMgtHC/o9C0ZEqu5+MWKAtlJF9VicWRnE+S6eDIjfG7KqXzGNWXdaWhW
tUCRxM/MOTV20+DRkDI+rGU3FEMRN42gq94isBKy9qkQT7q3BK5m30kk7tGACTEk
6nJ4+oUhp7P0sDAhwkZ8uqBYX8bftQE8TT3aBQf+6DCvcWzfrm1AsNjZwwlv+9SI
sktxa44qMzHaTrDEKKUTTtg7uqYA9aoSCzVOfvX8r7+NYuEmz7XscwqqBQC5UPFT
aRnKzysIFkLB6yIIYTNPyuJjgPA2YbjqH2PeYRNU1y1z3FzRLVPy5lU5WFicF6m5
Tm7gMUwKvtMy55bo63JNr2orRRYWaOjXSd/LiYqCLIQThbGVCCRsOWDrutPt2k+v
ig57D3YkDdpBD/noSNfndO/bNmfT0cIikR4EvfJvyU6hpc98VIjidPrzezS2dlI3
8/ph9vl2m91yFkxVHW79C1A5dbxUjtZSUlpQ52H/xogQ/WOci46QvvUGGRKPmYWX
E4fXOC/EYWxoiugRb0M97dUVupElazr8nTyAbWHtzacfeJFxD55i1QfKNkQ1XFEo
3uEEI0pgaQSGufzEhfjjg87K7gJoD93qH6v0urfo3k++d9TVtyoDkjoqtVxZQgeY
4GWmcdGa55usdFJd4Djoop/5V8bUHFdkFncmm+TfFA11RzyHt11vXlR7xiptLLwe
q230qz2lXkSc0cBdbcRjkUnjR+UWkTcsSEvv8rG+dO/8H4vyWSuOQoldleOCLmZ4
br3LmwxUurP+31fI1urEyl0faGYjn2OHZGlojH9ADfmVq5bpw/9oOj/lqnVqcqGO
+JtzFj/Odt5/iRdsdVl8M9ULQP1GgIQ2AIo5KzeTHgB04pMuFEZj14m8ZAr9ab6+
3zzbl5Qva0DuAIsSVy1p6VuHvwcDmdrlgkVP2ci+2tRg4VW1VWZ65Xx8kyrTN3kX
Ha15T+5+SDPGtvAfAWBKnjGasIRU9po7DxIWuS/nDZvgw+tw43DaEjmkzEPXY093
oGAFY6Bse3Fj/V97r2PhKeqDTXfmtBrnPjyWauyYbTqj9budUgt9xr/1bNpd8kC5
8btofdx8kaTeB3EhZIFvOoXM4XoamuMKYOMKhIkzJFA0SYG//OZ0AwU4yIkUw4RP
fXBqBGIfXFezQXyq+IKeRbHSZ08YP9nVIFleEKsQ86LDR9uOdL1GXpQZGHKY6vE+
afYc/TDlCtP1CbFz+OR9P7i+bI5DyGt6YqooOQhUg/VFrXJP0k1UyQozLWg8TMHI
mTnIs+f//d2hnfh4L/7ST9TpHLGbVl/zvP5LSOTVWVN3DHLJCPkeuqpU24yJjo/3
APmGP8uQltE/ziZnXwOamiPDG8A7PLAWZWZ9nSwVkUk7tjn6f5gr/OasTeD8qTce
0xdgoDBplxllWS3bcRjm3+rL78nQZioq30VduEe+WS9wv1/xElM9M9gBenU32csX
w+xRZM/xVmri3mmLXOqIoKA1Lmw2MX8fnnwAXmpDC91RyoaioPj/XwF6dCZPDj8x
1B3fgx8HuqotwJVgVwQIepHcuBGZOWBbJLwG8qDWhamd9YGx7FLb7IcAXot5Jqtt
8Acnu0H9tPzoo3of740VT8/g7j/cgVZ1EIVTYfdtlQSFdQJS6E7aRAGmmJ363oJR
70kh/1jvgNecH88oDUeFQfHmZT4HldmpnRHEM3wrJITMIc7C1EGyWzpO/0qMAI2h
ifBthqvqoJ+MPmQ4NjnbSAYgWg0EocX3RKJ2Tu6m4fBA+2eJH+8MXVRYHMkPVpoa
M3RLOCqQIBOycr0FTzwRD0F+HPLEaJIh0vVST+CGSJrTEA/Sk4rezzvyoz+RPYX6
ixxZ46X0PIGYqsXfF/bCK9Ikh7kW1e7dcxk+3nsSKgXiOmmtTNDbltaD5FrKdQPL
OmYCI6n9Wlvb9Wrsy0Y32QZn1CU5ZrcYWksSCE70vLD9wSt6FhY+a8wTpmevJXAQ
tGC4zu6MbknPaCqMfmySUfsJNBASm1I6j+P0fClKMfXd5BJ6oJi7ZKHAWA3/5wJU
EN8MR2HSMX/pSBap6KCw6+U5np9tZkUgeMltP8KVrv76DY5ylS4m43eX3qyN6G++
BRgHVGYDE2YYGdboTIRan3q/4sZLzLH2pUAIgyfEmtd580s3SbRkzZx2FarDyR3a
ziANqiXULBV9lKLrdtWq4MRUoYSzoKWZQXxxMlbpis2o6VkRmQX8ZAU8dRdqk1o4
i65+5CXf5ACtaj09VTk66ee4xgUribfl8C0fiI6lGgoHooXobQW41pUW9Gn09nKj
ecOhukrSqUiOrYxJ6vuLr+ZPUK41DFRSTRYJnMDPf9g3YmLrDsOnk3oz8QMSWp4O
RRIBG7m0HflGQFkzxilAN56w3W7wYCY1XplgBt1tHodERGH+wkGAonUnC3MA4Lh2
NdvnEmRX3ouInha79CZ294K1BtmCsG1a/Uq7+gDELfXdRulSnU68ZD2Rd7dbOeZe
UQ2bL+9xLX7YLQXZ+ar2GgBsJjBEEMnFlqaoVOy8oMAmg7Y8SpbUlqSwrdFOkIn4
6vDHsYB2i41nOzkvHPPlYd+op8osR/blN2Py84EQRhFaDphEaYjNIGwQuadsKjYe
r/Mc3hfv/6G5r0bGJ+Na44azNSEjVOprtTbH6ZabIg4/9h3GF8OAt2yyfnqwhMbE
N1hNqEwIYMoXiSiCIJcxfCOrutxvfiM8hikrHmfRbPj+eD6kW8Cl2TmMcA0TiZXE
PFmeG1HAWMdQ6uOay12d09it02/jSGbkyn98F6wsrJF6MpwBjCnPNx0SktUiYop3
/AHW0RLgUrW4qAXx/pD1ji5ZrGChSbYhC18SmidZUpcwB4l9OOI/ailnD5/CW24+
F8iOUV+ki7gHQLm/aLe7TVtz60I8xVyTfcplj0FRgPHLAVgMsoSweufBmT+gSDup
2yg8zPYzZZHKqk4peVqUT2VX5kXJNHrskhnyoHkpc79cR7uSsec/DxYDkIFWqTJa
LaIl1OQ0m62p8eOIlOqsvRWL1VGazdZ7F5Q5o9/1Stcu3ngiydYdCj3xR7UUbjYe
CJdjHDx81c5VMGVXIIIZYsXEgpx9DbatghBGrOVf91WXf+fB9pDpcmmnDsCT2KDy
bIPfN9yqjIyYoCYcNCmNf/R1zQhLKrKlffE7YetKN7c6cY7v2MSb+wVz68Br+9bB
BBZiVs+fAKeRbo5zvQlZGwVvymDUAr119qfodbYPuBHyS9RxZfhyCyxMHmvMS92l
yER2V9Oywa+WZ+QVpYrgwEfGGtnmEE7LF89x9BZmzVg4zF8m0gx97iN2RC9K/Z4M
aq4L5rOpsmDeu5YP/vElJqIS20o5ibf8/dxIl8nakEfBabRhvBKb+xXSuVZgfvU8
+0kE8+WouWJvnXdKaPm8UqJ66ZoI/JbBcbpJFufpxMl6NJhWYBgonbxm7kUegDYH
sLWlaCGQiXgurHhRMETxEeNQJVK5BYKj/5qHV9UApS1Xfy2QNCwMwz9RtUNgWaB0
JwJXFaVOnB95l0wMWysdTtWX0PvOosB9uRu7a76bPa/oirzKce9LAVVa1/bd8fwI
LOJJ1l6n9DXKXs42KH274+BC4nz7m4OKHc4aBCBmv2Ada1Vl0MPbnGLH3c/jtcXx
GUUfWy5n7XOIJGa9K4f3sFMPIqaKQnmogi3iOm0eZBDVgcj+mFE0kUM6wRN554lg
y2OKiNtWfZL7J9I5h86Dh/zjENOGt4goI6BH4TccSlbSjgU3i0rO/6n8lrivd2Sd
/438BJWbZJR2ArSfiDRin9356BLjwaaik9vWX6RFzAaUHeRaezh+buMN/i4DRsbm
sCa1ejchODndYriT7opp46weGHyrI+6C7NbBB/81g74AjpbZ0L0AMkcv9gNXaz0D
DEWdE+rMiviHiD6nCDtFvgcFal2tWhdBUsHCG8eif76BEr+Z4Z5Fn/QAC9wmi+s7
kwZX67piLt54Lyoxnrg18s2YKUKSNi4+qvcWxZ9eFNN4SMYGdWVEU1CZgImNG9yt
hGhoG9QSZL4jxHp7HvR0pxFeNqnh6ZQRK2bVzpiqlo12TGydg3aFOs+7zuqVpbER
KgfBr/HhiEqeO9NTmhixpg8EiQtaMmmP+YKot0pLIf4NlE0QnM/kUiIBF6VHMGXo
WOdokh2KcpMrXrUm85KFjqYA8HmDFTg5+a4AqM8l9Ey8/+lE9rDiC61GoY8sY7xh
QGzRCBM+zbr9iIxI9lZHP7WdDBaWf+XNkI797lNg6QL+qq+cnYPrKOhReuo+VOfA
dNLnCB6Vk5CTjvELYNfFbjzOnQquPRqa7+lnMENsJNSpC3tny8B1SCD7QkLQpbQP
cN9pnst+LOFWjWLTm05b0Ah05XuXMEIF1j5MBXqVkYxpjb7BUJf2fNWwkWqWUvgr
usykyKE9zPMQSjy6VAf7HamvS6+BxQmUHuSZOo7kv514AKRdaVNk9QC34pyVaKNg
OhcE5xKRW7k21hjMaCxZhZoMzK3W3vupVe+iVUQ06Lqg63bEzaaCxrt1kDMbPTcX
TqPw4LCthhgcwQZXe4NTcoILxq/b/xZWcnWayTX9Uzvwmm7dP/OpvszzocfMQd8E
sRIFWbpKD8uR51YUnR3qOIV+YFntp6WYuCoSXmFQVxsDGpf5q4fKVaUBRUZucOdB
JZT0gk357ST547gp7yqeb2LsS74K18+75DvEtsqYnsl2REMfsA5JievD1IoekSaP
ieXmHzbEohKh/3AQSGBtyk2RVgxqAJWziHz74OlTw/lN4/h1z1ddFd94q7n5BVc8
l6FonZelqaB7gvzvezsBDcC2gSrkDJu2jwqkaqjzYUp4kwn/uXVZpeFbTXen7jx5
xT5OHkmcZdyM+p8vIVbTczfFacCFoeLBCtzUpIyVnpIPu9q3o0adLFN1WNiVMpix
Fnv10gXV1jLqlt3gJkUoyMioaUdJjFbMUzPMtFExFvAecm4qfQ9DZM8D5xbBrBFP
rmrPwZqCQzpKUxHQqhpXSl3QLIk2BtVqQQaGHhj3yZw3f8tRHu44XerZ/31/T8Rc
Kd70e0ocVWF3nkCHybarLz6Vpdjvs2Vy11nVastqmV847Ybw/wcykrWP+nc8tzsW
qotyauCa/oG5pC+SJGurbfcNBBQUACGj/Y7jX2kzBCk5OKzA1LFvAjEHdIz7eXiW
DA6mrpFhgNTl6W2edbjb7xDd2GK3fvQPyh9dRTjJ4zLxz7/fuVLvWzcmiJhnMTxB
f1vIwB5kyAW7PoXuJT6+I8LyJo8+57XIwp7iolNYU8TN11UC0zPu1E9Mf9b9ZJ9n
bfuLJp9d5kHbMFK9KIzUoPW14qWvW5YvB7vuvyh68snoaMW/Quj4UK9MIrva1bQ6
HcnmgafmbCIISJaKR7GHpsLgkEBWG0eCYaLDKH81LWSaQKO5Si0fC4SbbkOdttJw
rP8UfGwv/CXVwIjL3kOgRN53vaUpdlkNs3Bhf62fAiBC6k4JJ7UWEXENs0x2tYzA
vwEhcZK2PB4RAQgEaC2OQLPs38VBouxGpTUBhWznQESy9I0FBNKTv8lUiO7ulMFg
zOXf5tbLnXtmTJYUobsrd1929/4zanY+n1oBPNwZiuScThvxt9Xhc4usGda7Z8Cm
JeYS+J1O4tS3iYlgMPF4jwzs5LRtn8+NEMMSIqk8RoNpU1oMXkM2IxgSuJFn8FYv
lVaGyKuSZPFjzzce06nWzK6BdafcUE9D91CQT9mTTr83+iCzFmBmprJHK4TwO1DH
EbYjahejMBJ4bLgxTgCeMQLG6eeXqvXZLBCCJRvMIzFSb5Vvlou97U7KvPG01ijw
iJHhzFrZrHfhdnPjvwX/eX4JjuUHxurV53FLEmnuZbUFYpXL/HQSD0lJqVJA9NIy
98lfu2FIgECaRwjKThK+bPoTPw1j7z8Ixn72wFOfROKIplPEpP7hU84TKcoyO3FG
pDYZzf5/H9axHOiNtm07ybgpBzcnWU/UCGacB0ufLiE8tpokuprro/2f/uC3g28+
XtE6wqw7qvnxp4JA/Wl5kyZMBoWXcVgptxBvlsA8J1gpjMO4OgxXZhf5sOKnM+JZ
m9JWrjrZ3DGDWq3HdDvao5EV0fAdh8Q69fAeJqOUBV0dLoZAFLuOXXbfAIlgqQlz
HcgeJ9NUJ0aNoyNtDgf7kVWzkVZl28d9q2I8XadsuydicZ3Ez/EkGTZSF2BJtAzQ
yv3daNIUVnhumGILPy7bYEVYJogT4X9lnpP67VjEeR4usdhvQHFqbKg40oOTuCGL
QXJWqL1EPdUcK9ObN5fgpOhwajRdo2aMqatbvpQvHLJ1bL/UOnH0Gls9Sooygm34
UtQAX//ZdlcW8mfkgNxlXbAGtkomeZpIiWJiyzJo9hCmZvisd4fV8MUFw7XsaFKI
YMr4IFVyQSnwIMrVdir92Pj9+m3vJKyNfKerTheh9W4pUr2RbfRmO58tvRUmCF39
reI0J9D5sAxsw7A5CKpmYdoWDc8d9ZClHuNdBU0q7PmywawxYwUtRHgITHtMtvUS
qJMTFNL3lcIuRMTVGuaxPoUJHwwJDR+fz/VZFjhMA1WoTuiSXg/4jEhcr7DHymHS
QnvpLlw/35P0v0dyOgaSzOEF8VKFGBt+oWquq4A7Wx0aUiz7/5KtGq5TXe+Yvz8j
Fz/19yu1koqhdc1acX76qM2piXLz0ME13sMwfbyWdkTRSgSFe7DIqoZ9uIfMhJYb
GTzrjEgFrgpvbtnAkha7z3e08NXl+OG3HAn9jqiacwPfCiXmmfat4eTUr9yDzDYx
ZEJigk4lK5qZhcsUS8jP3VEbWKI+Pw1/DpzqOBddlN6DI+71n0kblrIeFr+2sJba
v8H2n5Fn8VAiIRwMmwKUCKw0I2XwkGmtBojtnwFSSm8D6UHc2jGXhhCYIdrTRGLC
GyPh6nv6/CwaX+8IwgNDUmGTLNW6eoufoVYr31kt/SjumC/nvEf1K4mKdhYUoXEK
ANSdM3cb+kY9ddF/PItOKghbO6+67elwhGShDPDsACGlMDrS3c6rAnimAu37IjRw
URyXWTD7Rn7+4Biqp/tPr0mqGmjFQJnPbBAvMXJflZT4Oc+F7wshmsUR09Rbt92b
ZIYISxvJidtkxG72tnXf81oayHs79XdFqgF52qpK4MVLhQRPypmiex952rMHEY9j
obYoK1Yu9O6ejJFcAr6RFzGfYxqpKG/kKd0HbPnjInnSqqYgLg2sXgkg7/EukKSb
z54rdaa4hwSUyo/zup4nVkvdw9HgjzkGAcOgSvRU5VvvasY7DnCGFzRdPsvdARQB
BkUzfAzbLeZO3ihsLUSGgvK+LLVMIL8E3QG6iAyTXl/Y9TQoFeYdJxPGg61i5eBd
C14Le6yiuqhdMCTFBvaiPMfbIFyWkIcm/sBTofIDlT7jFPfQjbpq+5Z5dAfq8fgs
L5q5SwppCqTuDRyDtj/K8u1rdpcmjadc3bNt7DzpYSEWeAJxJ4uTg2ECWD9FMWKM
cAGfU1BHL6mRfNb15eyUp7FJU4s8FlrIFIPN1ckCb5Ehcm8i7A/nL89+PKWsY3QN
l46808yw7Sjs1U2r802S0806QcfspG0/PVTWZPWwbGSfnUPZ+RoyBbD/jSu2dXAJ
0lUhRXFEcF5rJJnLtc+0B4a9UlfUaxfbF8aIC1FASY8fGDJ+OpT8jx0lihNW9jny
gG9UlzQwanx4vPQWZyXv8OGe+9Q8zP2+5xsEtSkD4GdgQzTsUUuOkjEjB4OjsXLv
0LXihO1RczOBaNSjbDIHfekDS9e8ZoeLLd5Y0HuNDpjvRjcyTkcAKnWiDC+U7xBm
LoEl7pFMwD3Hw9C2WWdsetAmAj0WaOeiDOavJrd4OzUI8QFjSahQHXUR50pvQZiO
TNYFSe4YJRuHJ9eeppmWhkx86HkqUWwmh9C3J5FHYLOrdEXS4eK0xFTd9SFLPdy/
ZOhsekyIVEd87PIFkijc6E52+G+rQiwxzxsSmPXWQqxHOgXBxLCanj1ACYBKQrqx
HJedQ/EPyaOYv4j89WgxilzjDaPltNz3OS/LklbOIbD31Uuc5wmPz0VQHJHwFQKc
JuZYr6ISyAVJg8IKmeMh8wAVn5U5jfyZHjTtWGHgOHpUEURlzDKbWjewpai8x7Ly
EN9uGfX4NVJJ59WRPayguv3Cdcxv/W8L0X/diegN1hMsg26So5kb5n7iCrYvLpQp
gkk+H77y+Wd8SC1UfpFa1pb7sVVoFEb1nYiGXyCCoXPyHFt9YsjlVJGrS44wtvi3
v1pKm222lxjV5n5l8gCWvQFkY+mueWY0TBsDTcyjWhEYEUe4/3RSPiQEAEN4RhFM
/rP/kdz0o1Utnp9Sij90HBiHIVBm3Qi0edxai6vEUlIC25UzfbBdU8bbEKlV6hy1
ejaeBsFRwX5pOrs2Lz3+MD66yr58xZrBbA6pSGwvJccVh94cGFyL8f3tDDNbkeZn
kH9OYrx5P9VgXT7uG+WXQeX3xD50AJTaQPrTE2gYi3B3KNUfk2A7W6xN2BJzolQa
JAI4liaW9bQai/KKcwDF8/xH/3RY00frnh0CzlY68hEiV0KrhaifOtE7qgLCFvku
SPTnxWFhZmIFoVQd02njX8FdQsIOZ3S0ohIo0msGgJWm5iCOMJlf4MpjQFJVut3b
0MxoM0flFy2ff3Ir4gtQ8w2z4CwTG/Q4tKuMpBHcOkWPu0JF9j3MOXbrqpeAp/5y
3+0kvz0CKcg7usZAnE3Y3REThgbeqxIIDDxqn62zhy/FWj2yDTlxQfivBtQEHGVS
Q5jjNYTHGSymdax1syS49j6aEO1DiDVMyGD9NG9xKZetWb9BGp8b7BsdJz1f35uL
quUHOIIUBy+E1/G0YqlbJh4hnWLu+TXZkvQgcZtZFqadLV2JZW3QQWyHVoIm9Vu/
9cM+SSVgNEKD6iewB6y9MF1EmWPDQp5xDBj8K7K32idTUMxkRMrPI3e8EVPTRi6e
oziE6SpRlwp99oStgCQzzbmKgeaUwFFCMapdy9Va9UAGC5sv1iXB1UxiHJxNgm1V
96XwO7sbV3eZt8W0yYoG+esmP9NSEcUrgjo9vl3yoL6LcaoA6SUL+h59N4GwnLLL
+A9Wd69QCvp1DI+UdeFH4fOEIYt40pFuulFpTZTBFG4yeRWIFrx425mIooaZCQM/
QypvdiLJu3y3HkBY8GAW42HdOk5hx9+g8MewKwPbSo5/ZYPfaitXt2WL0JQ54Ty8
/mrK9S9Jt5ULThCWjKC1DuB4zgD5wio8yZDU4lJIn2yLv2uCBEjoQ/NZHj7VMox3
zjGebyuVOmz+AwwnDLR7cAIXaB6KahJkJ/b7PH303AsVCPbRiiVZAF/bk9IKbt50
9wLsGQbAJHEQMAhrh5QOM47ZkaaBQ17wocEwRXR8jxaGv1fyaqK90hvHZn6ScUDJ
iId8nBHajd5/j8hgd1qiLQ+38ZX9oM7CJiXQliRnatW2AhX8va5HzJmaSmNgA55q
3xCQi4UuTPtNgdKnnHKqtoDYT/SNSK5ARKM5ywsEfgOdZK8mmXiNt2isLix61Pie
t4rV+lD1SikVxUtd0nThRG62gk73g9XgrptYZsHRwZYhoEdbB2xF7mTxOiHBJ0oZ
My07ypM7505f093bVR143JCicxh5Tx4TFHkIsP1tBVqtq14dDmdfwTQET1bNy1P6
Ccyo55NSUQ+mVeOzvKkWzj9tXaMU3ebtvOn2wFMBaru9YYdBASCZNOOu4uCNbWty
SJwNzijDHQbemTq2HkhnrD7NGYVRRZRbOW46eZpUJUvS3u96iyAfztoNcmgaHpsi
AZt/bAvEviAt/eBvaP0PGJXvG4yo7Scrku9Yy13h9bk4AqGRlnPt90Hwi3O84udi
wS0EDNS0Mjmko73tLC+R9NDHFZ5f24YetmhQXD4XDnh48uKjPiTGM7wLl1i2dikY
TadzY3ol2HdHQh9gsiDnBqo66vnH8I6JkT8nmepSXGtcbtrITNt2nKI6vkH5hoyf
zdbwM+Qml3aWbz/MUWVuD5ztmdxts6kiasCQY6urBC58huPUzZswT2ElfxqByuBb
oaEhnEsSsw7D84/pZdsdrh9JP0JyNjLCo+TPGQoOdHikUx1ZmP5yT2jqpuqeGHRm
tH/AEWXt1g7l3G150cERSJW0GvzxvRGCom7/5KCVLydiCh2uuJ46QVnfsk5VES9f
4L3GZT73epSUSE3knFCFdJ/rkZw7QUUSvIQf2o1ioZWM48jj8ZxZyYK5bh8J1QB5
wkHkTtt4cqqkY4ZrUsuTcg9IfaLvHlc2CPx+ZNyW+zoTD4UzOnl4BKC85iYNn6WN
t6seRrKO0nOspI1cxFkeMhZFo2ZdNA/plT9Rg/UCjlp40U/sGibN50boxehGj8/z
bWKhkPCiXk3F7R7ciim3ORR22UarWHFLMHR29BfQKC6jDhdUby5npAJacL9moq4p
RHFJoPv9L7GPbjz3YqqsE0bM2g0GxlV7Zg4vRFwIz+c1ou/kmAQ6Ai8LabDsoAHa
Y9JWFCspEOTGTwNfLAg0l0VG/Fm/4lh8a3pnRmSAwATeIxn+DRFw7dk+/tUPdPgK
AodRRlRaVK7Nai2c8jgjsr+eysCc94VAIayAb9ZPnnA3rM7t+mx/LYPAH44TFZiK
9AYYyKWiZhFBYJ8SrFqL35K2BmRSsHtROGFZOa4No7Tlq3RAm76N5EKvfJLz3XSM
BYf0ujhUlC9jgiBJk8YJME0QFAgvBpmrtnrQ7NXuF6OBV9Y5w8Tafe+K1/Abe2db
MgibQDyd3SFg6WPzAVZ4e8HZC7yMecHzGjc46gcSPs7DUZjDSQLCeqlA2iUPGLo+
4izqNPnqf4E7fz56K+9PicPC+38uAOJ1lhX9ibDncKZE/sFvCFJYJQGCJohNL8hC
B81/obTH9y4FHGIp4joABCcF7emZPdgfEUDy24NhZ5PT6AOnm5dmK8+Bob8wJdoq
NFD5M8Wti9O8jDlJJre9ZCz+6zb4EOj43z+Dhk/dlW7qqPVQMl1el8B5eNmkhoRe
7Qha9K2M7s5XYiCOj0+DfrF/QSCwfjLfKBB/KpbwuMyHpbwV2k1QDSXUsVZiSW2r
JcqiIoFxMqHvNbL0SlcZiiOWm/m9aGA3JVOOchajIxET6MP2jGoIyeJhUopV5DBY
4GhhiTB96e2W8fpw9/fuFksyyBCzXu1FHAO6A8PTPNxzl4Toy03M2Gx9m2EEm6ni
dEQev0sx25oLmyNewkx4DQ5MLJD9LAEK9YR3J+sEowc5o+pU+Ey/GFVoDGT8H0Yj
W1MBsajlSvLyEc9lIDzJdQJ3U64Ye63eXMaPMWcm5XOSZgt5AK5DM9JU6RWDx4pe
clWs9SRuEWyUznI8mmscSihI+jSuWthTuv7It3fnaUufoE7je/0Ev64YTDQK3Y7o
SVzMqR3EoPFTbYOtNftN8KQoa+ml4DZLJLEDEsxfzKMtb2uGugPDw+AR1BKRhABk
1LVeVAQxSmAAdJCYEKuVgAFrZT8cRisNKOPyVEAhWbNwTpQYxCswejXypPcGpjg5
dRWRicdn/Nz3yPvOqWL5ZW6epXp5NcniSMwvUONDVUc4ZRFDjAnIyKDvkLpakk3X
tHT/fWoBryo4CDHx143lUCRFiLhhh5p7huVm176XlBa+fPca5CIGRqIJhQhK+SxU
oqfhwSp0EwWoup0JczDQOyf7hiVllwq4nTBw9NIn67gNUMcRXf6OLwoJ534t0LAL
e6GObS830XprO3h8+A6hiQocl4eBcoOMXf+ei3rz2XCeHlBGKGJ791Dq1CXWnDC9
ghegFJyG2WzhKhSPAbRjfBAeN7U8tuVFN/tEGmCG/X1KCBNkHJExNUS9tSjo2C5d
pN4W7zaJA5+5S77KQ3wrCyQIJssujtZ9iTDq//NfP5sn8J+6o3rdFxeebM1YCWtn
Bik+sJ8+rTQTTfeq82RukOa8tN0TfsrT4Lv9lQ3/wK3U0nGJeGY6VokzgN6cGxiZ
pIlwolyq+RQ9chT/WiII/tESmxtW70IvjAcTGRftmtgBE/upraMp/ONVgP3YGet3
B6Xy0u8FVTYlAeQmug3zFH6CWOsXJoSRWXcBdNAFKJtpS67VjeMwZU2i3307LHQG
B1iBgrAQSqEuLV1zes+Ezf0Pbe3bXBNGMsoB3HdsgqSz9o8cDHePGFugcPoop2sl
zRkxF4umr568E8W2cYwlQPSHfUbSXuIpNDla6iz7ElUkLbjg/qn37T99/45JeffC
Wz8oAZdrkX8KvStMamL2aL080YaGv4mPcTcI78eAjxB9eoGAp//ezWns5AYmgadK
rBEMhxQTZ3iG2NJIldBD5iPOdWinEy750GwQDJ4ixWO+glk2uNeZXodv5ag6DMYu
0uK4RcwZougV14BVPU6LJIaqOEcFtYmMk9pXrAcAzaunawd4co+F3fhxgLtH/Kn3
iHKBBR3oMn8QZv3Z0OojQ7tNgYoM3+L9GWw0ZfEVMe39GBCZvEHKcRURwMPTESk3
PZQ2IDTj86QfQai20R3x4ZN84cy2qIrQg6sAq1VeHRvDey/hgxbotMieOLWS68qH
WXW18TIQ97Uhx8RXFTu5AEBCiX9zdAruAyr57umATeARE6wy8LbIW8v+3LnezxaS
bCQ/KXnyhUT9SE+2nftjDezfnfNN8W+xr9Or6hALoF/69VHpUCv+C2x06l1Xin4e
Q8qT7I5oH203vYVsABv3jm/I0pIzEk4QrKtp6B/itz018ZOysCM/lN70DDZsmGaR
baSNv6ZSTP+ZDZHmPmsEa9Hocg7SxDqduq/9gED8EXQaj1vv6m03zNbuaSN96M9P
ha5eeDfkim66tcOT+CfpljFesidw3h1hmItRmGLOdQbM3dKlXEgJsrv3OujrueqW
0+biQjWaMM7VXC709FEPFnIaENQzTXynFQdTS5rDxZKp6lWAZrDVjhjmkVSN/lJT
tax3vSQm9xr2sW7S5P7V5Ue6falEAFPYzmw95p+P52ePkQxKTQu3pL2b4qFpCtko
ubcjdh8jYLN5ogY7PzVC/Zx46aHixssRKEC05JaETbRH1+imTyKwprlSnZM6e7Gc
UYaUftH45nuwG+mTODxCDKmBXgDoilTUiDJDaKoWpZCczXlaF9yoHZWY0Zv8S8wG
X50U5rq4uo+T4/elJ7dg58qyOk49LS/OGvCpEqlLMHtuN2RrePyCsRxpXxaQbEcT
4g1UZIjor1BFCJJqKbBTJPg30Ju2IMUdz6W+jXSv6jYzPMdrCW436ONrP4tlekfl
ln2VLtu+PHQqpKABKZ6XDapnglDORK8KVkWOMJDtorr/jZFJTSIIvULus17622iU
p/6v0ENjkRZckwVPzlYGD/KOv6+2dxnVHPHYT7zq8dQhO5YYJQJOegWf6qPNAnpk
HY8MsCHjtAg4wBovsx87V1w0pzUITJiI/B9G5Lm9JqTqfBmulMBc8OQ7Mqxko/a2
ETLUO/r+NWwMoO1NQnvGi16R11wMvITZARbea7e44XM0lhRQEou4u2LicyjBCMyB
hx1yYK8qrOL/Us1D9saVhpiQTl5MuMv4c88b9k9O6axx1KMiQeijv4CDyMhqtEtn
KM8GORn0G0x7CfDPW8043ksGXkQz6Kh3MAsStTQ4f2Ce0hQuj48ygQa5Ng2RwTmI
dhW1nQDuaqeaz9BWcb78ooZDuByjh+gCpGvQr+WKjpqy05CbERQpcq3Nw3pXUmrY
JaVQ54mII0Q91pWGpAmJeTZA2FE9S6CDef1PKPdbjs5gKB3YS9Inix4Z8zdxw5ax
dWWSdS/UvwBaXy1iADnFjNzo6aYodrVSSymCJArdGTKnJI4Q9Xsx2uDivE34GOBC
my/ig0h4zd88VfSN6KtQu1rbLB/gTp8pP7HRysaBh3fyafZgq50OckG6SXJiVSXK
ocj8ciVf4C5vCGnna5+nePAmSQk+70n40QumOwVWdWV5w57XkD875UYiSKZ+rkMV
Th3s6AKB/yLsafwFT9Ql3bWPhruv1CLtIrfCkDMpzbFpIhd2naFZ6yZU+e4BGCaG
HdbiPTmDtb1o9xKEs2xiUE4UhczHEUimIhSB8BX199p8W0yQ1OTz2nJCnyIf9DYX
310LZ24LjBZOLtGn93UuMwx916/DhOjYcOPILni7APG4DXN0L32OQenqBwnhXgqS
LJh2DYbKo9sbIRLsczme4DX512UANfe3+FegCC6iBTyRKN5XJ0vBJxa/7yNCs6D8
fqCkcso5WHcb131W87uc4wTXr2wadmUPk+nnUT6L7fv+iMlrAkZFp2iPKkEgNjFw
m5b6FJ2uznOqGEkRtaJ8NL/IUkUb555dV+4+h1Xn/Vlkp9GrBjzMRfvwbDmqOhki
DY/0llXlndLs5faJ9v80Uxa+j7j/8yIzv1K/kECCLtyt68Mo1jB78lC5hzZ7qpxu
/+WRjzkls38P6roYiqLhPrwiYhHIpWxkyoakaUSAwsF00kkv6BxM8/17eAqjF58g
XWOfq59245tWZXdojhZRvpZgp/lNxRT6xRsROjuQE1YSzXmBB2rC90sYSFXJ/47T
9PjlZkUo2LL32oCgdc6wTuhY1DdnvIdv6UxKw+808YmO9iZMJqZ3caJI9KxfM6nA
1ZfCDNKkpJYqbfwVWuBplKaYL1nV+WcX1+q/Uo9wCHx76BF5O5owtiNu3camO7Zp
SUD7RwFu1CsGrmA7YU8DSpDUSliyKb9YyjgJvZF7tecqBKU+lfyAPWSlMud+dtvu
j/2UktgY04wfJBsBTdGsUIslptXbyCVYBYTZiXLI3XET9cj6MO/6GknZq2uFjzFb
sj7k6ej8nyEf2r6bsOkCmCtMvLWB9X6CkXumrVkfjyzc3WY01sYIhPGz5RR9qZR7
rUIXmNQIGHjK98HmUUtMp7z5E+fUHOE+8nvAYaxf1OrlZJvUgSODB5xjehILodig
XTa30iNp58BzEfRHunv3kKR0+4pdiZH4zT/ATNRtGkLUu6uVfsyGew00sGo8WM5M
CKXhLYIdpLduEfy18tPXBhGYUkEB7FrYUIAz88nhATRYTqG9q+b9QJFxJMTa6aWo
qh00+nnVKbwQ8j79XMkNVifsgs22J91qsQR/ayRhZmMvkHuXQ1YjIYUR8efmQ4Jj
CAP1+R+ZWhfAP7mQkd9hS2H9S1wXlTknE+JSvbrbiBjr/yjc+NQsPN26Ralh2HiP
eVsavScKTjF76FyDjjZXjUsODi8zaBe4zO/Ztn6lf7YQz/g0Y7VIUoVXnAjNBtOi
AeU1BvCtCgdoAIUnuoCrorTSKqQ8yxbutUx3xGvpmjHY0oX787QnI9G67gsIxVYI
k1SVCxyPaOfdtnL6v6B3OwDDpxuJfkcgLjHHaZEA1FOjw+RpDk6JNNXKiGoFjf4F
e15LczB+eeZKN9ee9S3m/fuCbscRlSrJm8Z/fPekSHLMrKCJcvRTL1x9e4mM5D57
PAOKKLoEw9JgJRqGbMwHKRGlbgLeolubwRZiBlp6tPmU4hgvHURldFhSuFRLHxQO
tW2Tmd29mMLct5a3tO2UxdwnSJiwzPRTamKW/eaUmIsmOdt5V8U3ZqZJ/21y1jjY
l1sukqUPU3rHZLRT12pmi3+mXbooUaBDCe60+9p+U6GlMXcTpCniMhSmzx4swkRT
88DF5+OSZniyKy214fHY7TqAIPKK64rqQtfeqRPDaOwnSO2h+MdNtS2RxmPxxehU
DBKoHWSVO6/pQZUWBuQPuAzIgf1XRvgJ0E0WLP9kyYxQ9UexDbRmRvXbLQacvfS4
7z9nB+nsxeE21uGFQNdRQHReeVlo5mfSNGcbUmIRApc6G8wXpxTDnAc0gHe9zbPx
Yf2qjm5Tq8A9NWRGqXGrmwfm7L4nz2f5gX+qO8xQtBRkva+EWCQ3ZCjb4UblHCoh
ZmxQcZ0r5qpislBqv/Bn4tajAVqpGkFIE70X1ETSElDIMgFh4/MsQTig7cXMomki
tfUlGfgs81yRrP3OCiYs4O3z2jPWpNEViTJPYMELbnFSKZdBlbqvUnO/Qx4S6NiT
/TiGEw6GbbMzyH7948oYhfiav7/CErvs8xt3MYaDfWUZJB0gP+YBIYIO3pUthASd
O1J12RAFrriWcjPI8+7R6Gv063P4MvrZIMCgkupY0pAEPByIxcSUKbJ6toRzDOcb
/N35afbneiBc+RrpWciFXqLi8OKRrKemFQ00H7wW/ULswyPHbvZd/mjGavYPKPh6
XRtDYPWHpnXaGTUK78I0NhpUYU6zJvRrKeL61t5/1A+Z31okl5nMlSz3HThTw4Wo
IoARtprbl5xnyI9/+Yps+ofQRea7VoaDYWTvA/NROjOpINR4gQD6KuAks4mXdXbQ
7gy0W8M75TXSWZXLhG7pvohSHPYrulkxMgahccgTgk0AWp8CsrZ4AMH7RFaVKgmU
VENv2amWRi9igtaF0ZdffrWPlVzLZlfR5J4FBrksLSOYa2twaSqOi53VYQYWerDS
WaAM8hBYTPgWKQxnrUgX/mvZZ0g5PHMUCV1hdFT9rHQBRmLkAR82vfvh9iJNIJO7
tiRGkEKQEqY844SVc/uhNNBfLndALueQkXpDj7QEyFv0b1AtrSyV3yvAMiXDPHKn
Y+02WOnv+ZNkWG6Dtw7VIfEFSqI3dWUylytZWv5awTAWWvt+qywyVMgTPl6jfW1H
FM7a1cxzvffFnZs05c/ayw+I2rAC6+FLAVqFULnb63M1ICHIvHxEPoMbOt8+SVdb
kv90JIroJMlhf1DNDXhm5J/H64pUjLIM6+kQ3Z7wJZKYwRZ43Chtg7fDM2cBkhyU
jjA+hlgPhsER+oYjrKgambOFqgVKvkIeVgBhlPb05ei4z6viHnKL/bN2lZ7ISfv5
YD7mTd55Y9OsFIWT21OXzC92J3HJx+PS8Q1WILQsgsopcqqS0p+hpgoalXfpcGlt
Of9NKCFbV95FgSN/OwDX+WvOXTXJMYV+n9vqiyEvrbtlyqXsk2oT/6TrRVj6sWIc
tFySag6+6QT1kbH1IsXtaBgYV9K8eeB76WhuNLkjRPwYpMiWpDBVXwOcuFx4yPeR
t3V/Hckh5LYmEIvuGX1yG3SkJQ6JWRk0OxrCguuZdDpy2f3fxtw9Xy4RmPT6vAMw
Pk6exg/iDZWPXx09Kj5OEqIdWzfcv5Fnq8l4lWsRao7mB3vmrvju6kQxK4vwA4R4
Equbs+Qw+tn2BN1D6ttaEl7hCOqv7Ft1yfwimuXzSXbjCr5R2CbAQlKsimfd8Ul5
j6wmFOlV+ZUPTNOdibb5L0xqWvemwYkGJP/2486Ll7df15bJw35i3MKPKnxuXCkc
5RjdoUy7NY4I3ngGqdE0KG6RvdOtDBGUN+7jxC+7Guz6ySdz4GYaaJ9pU76eF/AS
0znG8d/WSLfNyuE7qN9ihSLj5hWIBfptA8s/tUB00ert+JWcjNVBddFCqtRjoYNA
auKUvfe5O0yRFIhBKmxkKr6rr7YjR9FXSvM+2LB/KfYzaI4Q9iUDuU+6TQvmxvVN
hOwJ/pBcqAvuoS2i+NVLibcTMv/4EqlM5upDZdm0N2sSDYfqHxMQNdPa86sV0bm2
Lrp5lVf2ix2/Ule0rFsDpoPJ+zdAvreW3o3lo/Asu8mwzoj8fYm1mRf1qSGRlKbH
Jz7Mse61b1YXwLC3UwWDEn4j2y8cALRUf34i9UpN5xL5siiYJHtFXaK1KlQolWEL
N54Iw+15EmEMcD04S9cvgwDCewuLkWHwzE1kns8Lqb2edipPBWm5krxE4KkS8kqD
C6ZNSyT84eLCRkJPoxuiOXN6TTXt2pF5hADMTgCQ8R68ZsNmp7O16f7ERbI0v9Lr
5+LdhNRSebIm5ZQZw9Bh3eWuOJSyzTVRL8qE0baQM2V/x+TgXaRNJkpnHmVKtnKy
E9oODZ1hQmZ7YOG0OV0kTAPWzr+Zn3Ib/GQC5+iBRqKjR7XV8sn32pQesZhgYnzt
z2LQNvb3gKqUZnp92dPrgmxL0cByNd3xXkvvFOyXEp5IisTNDi07nEHrdsm3Ze8Q
mOZ2Kgk0oUwySclQVK0S1DPRjOKYb6YM+0qDzkn+ZuUEFAvv+1K6crTf5ziDV9yv
cTVNy+3f+E2LuQJaJDXhWD4MxmQxpUGvkqzKAGyTl7T6JRuVvtgcwUmPA/3O1SKY
UH02KIQygxej3CYGb8KL9cdomovc2Lpy2HOiY0+rwKCy25TVusN9+mi7xKEaQxsk
XQvBCcD17t9QmCh70UmBGM2bN8dqb/yvevJBHdz4CyL3ZIFcZzyI1hE/Bl5PTBDf
azdJBEIap91wEunZih1enZZn9bQ5DjuJtcO+buZANJvPegQMKuFwxFEFoHzHw+hz
mN/0cCDE+lGS9P+G5ALFxikHSWlpZcaCyRqrSdaH9mJGfUD4xfcjqbIHKoLKpbDD
M/OZ2jEbFAhc1NMU34OZUN5lTz+qpE7FFZxqnpGCWpPriOL1n7DV0ad8RFyWWUa7
vfX2+URUAfkAov+AczggqHCfMKsQ4LDgILI5S8zaagZeuj3Ov9aYcwwuigxjXV8X
+E4jZklyWParRlLmlsKM453jnm1ykpSTkxezzis66oreaz9mZeBrdzq1Sl7ePGPm
wNkTFLIe/MEZsQf8kdIGmgGub/dOhjkFw5fI7l51yKVOP5sGOcT2ZQT9bbUQR0o0
HrvvgmWSTTGKx8nodUqxH98kasAGliw8VdASDehh3C9lu1CEfBKi1b4h94g2OU3B
Y+t87lXQtuqooZm2NPyfOhsx/EKrZyLxpYE7+T+bSWLb1HcNvcjdxKK0ZTViOPbM
b27dR+hQNlg45LPok8V598AqrsIH1ZACm2N+FLBSOhMZKfQEH6LB+fCPKpHurvzD
frOh+NuITOW/nK7RxSRMgWcMGpwPdYnUFb91hVxZ+5tsDnw4U4OGBpE4Jmo6WNrH
q0RmrMHV+sLAkuJEE6T0q2t/kDCUQdq/EKBLXXYhAaFo1dqjdrh7oH6y8bmXykt6
0cIxH15ZUPivZkhKzYJJuah/AriE+lC63FA5oCPETTeXYbznXKPbrlS/shnjanOL
6sDZC8Pw4zHaTCKvcR4vp9x2o/HyJZzYihSsBOz2pCsdijCkY8/3+QUzfXKeeVFW
xIbEemOlsrNq/nKOzCHl4AjaiLHE1JU/Lq9Y4z9HlHuOYrol8Or9u1G0SLeN5RyW
7A7WA3Lal07+HCAp3x9TGxiabN3rWHA/zsnMqFNFfe4/suIavuKVKklp41vji6wV
hHXmhKpkIg1R/AywdPuhfuVlpEkjFPoia0K1RGhtLT8=
`protect END_PROTECTED
