`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
USxFeqBqNNSLYfO3ZPAHpkKrRVfq/8htOraimfmYyPmS3N3I8vHYLlh1h1X/P/wr
xz0VdqgcCWeBz548XbL5M6d6Qerepk1QfKuWRHrCACqoKKm8Q4v9GxbZKYcXjgXt
tstZQtNf4vSTA8bfdwJ93ZRgg2AU9BEIpVtBwEnqKFYatr52BwalXrqOdYazWV6z
tsp9nD+b1KeR+QL2zRe5OnvbKe5sBOPsMv1d4d4aJxyAMJHXPXG+cBG4d9xJU1TM
MGgR1+jG99dT0TU6FmvcZxHqhM+Z/ecsg+yxw8eJw3erl1NSZvjzPWtW6QkkMQfu
cSkjPj4MRgUUIC2hTehmyYkNh/2cN7UsAZ9RlxbRPl2q7zu2ic3wHnZ03de5Jh11
iJfZucnMvqe7HimqBEC9Dw==
`protect END_PROTECTED
