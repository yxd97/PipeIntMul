`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCFKdbq8Ys5CYijiIoI3HxheJ81m/Jxc+hWEYrNhvudcGQXqblG2A8H/rcSlVIym
IDs2yogQg260FGpaGjEuiYWki4RtXaYlYwvESfupalzugTWwxunyDI4nITLUOGJw
YwHnyUi0AtUtOOKTTdVQ9X/6uZF1Pv43fstDNJVsD8FxVqxLb2btUxJkotUiz9zd
XjDE2ekxwB39CNgFEl6nKaZPrNSSNN/Sm6ilbxB7+3e95OODTHWk8ivJYrLBOYtu
volWL9Wp+oS+8NxcsJDFqT4C6uJQIt9OsxNcEmy//QsyW2fNWj+TN82fa6Awy51Z
tNHbgeHufPrOTPC7gayk/70MlndciUPWV7cqQd10M1EnELe9+GT4IWouUo1+ndia
9FmxQ7sd1CNPXdf2ySeWcBJECq6NdLoNECmvHX5DxycYCwNEGcAKuXMMWBkA8H9O
8kr/XWbn4Wkb9jfXcwTjEVp+1zbjvRykMWpIHxv923k=
`protect END_PROTECTED
