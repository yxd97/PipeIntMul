`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eR8vWpXSylzzNROe2wHoQ5Ty8w/HFaP8cDAqEJCgR6Wz63UV1Vq9QIv/dPTIJUdX
bzTtyVsWb8dQ1J0JoTd1DVqJKcy/s1cI0pIN0U62DZsOG7i4FdFUQO4/MP0IwLDa
0kDSOszLSMNv48wZ4FMJlhpZg5GCEvoIq22FM68ClVj0x5q8WuJRjif6QtXo3xxC
eXbfOQxLGVa5APiS5P0yX2g7I1jVlNp6VzvWm0lQJ0DdmmkFJRbe8b/mowIlxMmh
6psRSs/XEFwyCJaa8ZoIhGPFxpPs5wftCVMRQzoOEYSaEghJO0cpAC7+3hyhmmq/
RnBLP7kv6++4/mCK8WYn3GU7wwhF4Y9jBpVnKUmAxxlra+2Vd/muWly8lxmGkwov
oLKHx1SKIeE9XhXcNc+m1tkQGBi7IfP3ORqIcO2KtS4y7G+I8iES+s50WVOviPgx
zIJhYOoxe7f01JvaFpR9UuJUQgp65Wv/rTYRUE2oF3yg0du5jclOI32wXxYMA3SV
D73M0ZDXSySuE+jkdJZIm86TgYPq52el7DN0iY3vApdv0Fkos54E2WnvPHLJRfD1
SE3GPdyMKOfHr+nBdxHTl0Ziozp99zDwlyhi9ggIwJGhijKGVjljcQI1Cu63xuty
noanrBQTLDX47t3EaVX9+itIWQw2AIck32KflKXrVJvTlcU5xt0UfnF9U/KY20I0
UGJroKMicXizybKocUJ9rw==
`protect END_PROTECTED
