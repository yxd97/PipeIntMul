`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GfFDaxJbyoBQHx2niWEbx9GM7EXUYVLEgZtbQjIVTZ1cLS6Ek0NOCr/UAPQJ8sqP
xrClteyGPmGxY/KaxgtD3uFcJx04+P5duhwGWoiZCMdquG3jipSn4CYy7Vs4ApAo
tX6r4J3QBVAv7mdW9YC21ffhq83dkIRhJ6x+spkM76H/M24VgcFsZA7/YfSQ+VGJ
3dub+TRKUap1QOOFD3URwtoRh9juiYNsD46Bzk1shaghIIunxndaZRi6Z71MKVtP
0Dnfe2keY3ZKj5OMWe22dx8QuazwcCmGgg7HZtuOelW9caM+UtBFF4YbJf2XXBjm
0XyNR22auqaqNoEyzH1Ry082t7HUTx52bUwjBmLez8AVQA0gVQFmrMCf3NeZZWov
Hu3uHyZVIty7a/q4RE3ouuZTaBDGficcSEE68XmsXLc=
`protect END_PROTECTED
