`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NU4OhmtruvIcO3sWUrfWey1+OyeoMKhciyhbpcjpA2WqR2QGntxjHZMoZzSCCCrG
lwvOsQ+mrtZ8u2cIG1pOHXD6KBYL824fZmf9abqb1RvCy0Q3T9tVKiBFyKjVAWOD
eK9NkntNXff7iP34sNMt0kULVTbLZseWfMGTDQXHXM9+dfFg9FE+KZD69bpGc5xg
CkoiO+i15Sjta2i3fsCJRLHZHWmSbIgZjIttRxHuTkjUM3uRvjUMwGSvLJyXXCr9
m3cGmbEXn82hltCkxQVBtFalHYD81GHKmYbuyYHFgWF4LJ5qcmU+EUMfxd8GveS6
ymIv7hAadl3sAj5c9IvOhISzIHYtAeQiN/2qh2hlScxCBJPIgL3w70FYytVlX5VW
9J5SKVx8N3N44enu4YE5KDjUaihaGj46n+1DGM9/2HVNiQDJZwSMwXPjXfXAvCWN
Gdlo3Az3V4g1And6UT9TDJiYuMpqZiysZ1Tx7jwameSSq2I2ZfwtmnaJV48ma9GO
vVKxugfKaiMdmKhs5DRlCYin3MqXAtp0jiA3Rlh6ckYQl1ucgi034l+b5we5cK0T
9h6o/hNISncLRQ2oj51Y+txd95ePnl4GzpFoEhVdCc4=
`protect END_PROTECTED
