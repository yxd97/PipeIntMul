`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NLE5CDscvCQ5dojlIA16ri5BoInZMzt7SUgz+s8lL7ALc6MlwXnuKqFWzq5cUX3D
U2H17uHJFVKVckvVdLhGsAyZbDNENOylY8jJfcEwR2Qr304IPi1OJdhHxcEFrrMV
lkXMidxHTpdW1u3sd2Ws5oeVUQ8MOptxL0Fbmg5U5cov+AMygE/kMJDDpgmsX9RV
nmqVkIyDwzi3DVyd0pOFJCaGhOIkElPFchs7xjVXvg1NBb69UW0mgusIyp1dGy2f
NNeb5C570lM0pUttmYilkqNhDlaCw4y81jX/C+IEJW68bKsOe6pOFe1z5crN8lK9
r6IrU7+c7lbUW8un9yW0C4nqM8JO0dniL0BGs/N35wqSunIC2wmMqlGAuMnWkoiT
isPQA145lYeFIclhuTDdjH47K0VAOuFSJOGUwZXv7P04MyGwL3XXfkKs2wpIb6ma
pIkCHeiPD01+/BnnYmfwTl1hxNfFF2+GsguHrku94EuXQNOsgS/TZTbvOWdnf9Q5
v2ljv52NHqm8z+jRZI4aoJkCVR4g0Wf9HEij5EZnvIZDTkM3F7zjjNvt0DbxYURF
kxLY6kNbOeDFw5KfiMAP8upAtNS5AZ3MymBlQD0NCZZ8e/L8jqM/LDW89W+PMf+O
Ihco8sYE6wp20X6RzPs7k7dZECIOw8LO+b+bkb8GZ8/ySDPEMBbSrHyVFJGRlPgv
Q7mxeLbBl4x+gJDKO+Tvih0zSulQPZeEvvUmsCdEo37ZczYxXPh9PT4K80XAgNtQ
hh/hM4M80rNndZTIbgQ0WPf+aLAO0ydHTCl1M1IGb6Nr5Yld68a1WdrFyvRElIRS
2EDPEnRLZWmX1fMPl35efg+DGAIjGV6MqYWLcxqlvIuTdvRHRPfm2G7SfxHq4cfr
ryZJ+jcMIy8UZ8isvv8967KAOonizwpE7eXQDYlap/64/Kc9ivb607J5NXOP24xt
Kq2pboxuFhPPeOFL66VFAaVkGZK0WhyE5/Aw4nb3dXjNBA7UgaWyH2feQyIE6UZJ
`protect END_PROTECTED
