`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jYCUvDAJB/pVOTPXQYY2VAgefoPR+iCxjMBpIpD9yhz1knmrEE3AmapjpX04vD5T
cXSFYVMsgk2SXH2qD9dYRdBd3T54GxhMWvqsnddxrS+TmuQFdTKA6YjOUXDYZ9b2
ouQPeI8258/dMrOBNRVqdkC5CtdLYJ1nDU9kgEUU/ZFK/XRpS4aRVdN2zVovgndi
mIHfEdFpZmr5c88Jy1edUKM02XSx9vULFRkH+TqVF3r8yC6MhGhIKd7Jps+2TKIF
sgYGyWvMYKmIbicEsSSymBhwj0PCEAaaHEu3k4pmraA=
`protect END_PROTECTED
