`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pAOzz/ClQ/j0Axrr4pW8+yYJcr3auNiBwnTg+ISu9SZqkFUwIEVfnIITeAsAiiz7
NvdApBNXUXVST7qqxuYeHFJHrLyMUF8/Il70VMIK4TKS0aMW6LfN+bD1rkBDSWci
QBtN1AN7K+tBcjvDNtsPBXYwKytp8pzoFh3/w6ZnmrPpB63clEDUyWx7dDYQLzCp
KFHLWtt1GI6OLQi3K356sVSmX5XWKtyKjJX88P1Gzc6JdWkudjokry473FmzsWye
IQsOEbiVyh29fvXQlFF2wimhYSwx/CEPqE/EVpna/JXITRx4bDdc3vAQUeEmh9jt
RyW5Wogtf/hv0mxYDGHOEbvLsjnl8O+nnYzzpXZ0lX6A+nfvJPAfXAZJr1gGg6iq
4hqXO/+0zxhSx/bjBqu4XYvyGljYBjr2mqmuxbD3BZLUBwbCYbest/3KStbTT+rf
bfstJ2lS9dM5Xu8FkKHG9KARhoDZ+1X3Bcm3W3T2MjBD9t7mN8Bajjkhnc3S2GOS
fsvzT7fMWJ5JQdIDD3SY5exDwwEmYKHeKMedEYQjngKYpSkkFdeUS8xHJg3PRTIZ
inhno8wvRqhws3S3R7QHljeV7fRbY0WZSaMB+bFCBysek2QZE8Wxs1U0KGcbLUHN
oA/1aqkqlvMZ9r/mdul2WJG9YBWtsmdn9smc92n0UDbsrTKGNXcBusios5avIQOV
VnwknDtC7CPvNFhulSuc0XJMlyI7lUkfhYXuJLorycmoHy+vxRGI7rTvCg6lwg5V
AFuISDzjTPGyoW139LO6yZ1teUFlZjA9AGOzoiI6tlzfmSsVAkdnwzwDlw3aW4fQ
w3goCgm1c20qFxtZ2xUNuDwwb+vI9cF6FNwIRSOSAOl1jnkylRIUqVkCL0OoGuG4
npRX83bq2wODU9B/aETMPF3CXyp+FCQig1Zzurw2RR3jF0BxZxM33XE5OZF8BdBK
OarMAQJExIOK0oMQuYUk6+Zz1ryA5lzzfXtY2MNraMwBtMmL7MGkyANSstTKoNcr
b6VCGLaWGtCSmhIOnh31lyxwyHU9WqJLmnoarvMTLyidDYvB9I5buaK7w0w7oeTZ
Uzti2b7vKAvhEqLm0HS8gfY8U/W7wA7yxmptBN7TeJsceV8o7V6YGHv/SVJUEEzd
1yNdR7ibgMMEswNi99tYDQJsyWo/1GDP0StABNyafJYU1IW2Hic1Pm4nlZKInAaN
SzI54aS3jrtmqHp4VEaHZGmVtiRwBmMwleZlMNbs4bBCHB2sCl1xmKfrlvpEeBiX
1Wk4iT/xUkRjXmBnaOyXGIAhKh8CvgzfLhkWCKJryXCjjCob3tDgZU3syvHFiH/h
C4FgYEJX3WW7oe2s4agBcL6Cuu1H59ab4tZsGkDYfRKHEUIUFPy4bwMkTB710fEA
odzr7A9zuNebIDXxEceSiHMIzqopHBA0PcpUeRncVgNpP2gg/svV9s9jiL8BIk6b
No2Ql7bKlsnzxYTUjxeQgXtS17IR+dGA+CBLLgqQCRd4LYf2dkaS1vkBXtjOTYzV
PYRbNaar/6USmJR42Y0Y6mONpLUdRkcchRxwBPFJ4VI9ZVHuVMyraitH0e/nJf3R
dPo3YHNbVxKBgH/QULSxeQ1kzO/HqUte95nD/SAF2SHL243k8dcN6Q7DlBjqR3B6
ZA+qTj7bLiMqNgkoW0WYj2Jiy2X+16xmvMTMaUWo/KyUIvHT+f944CaGsKRyWVl3
N/vzU6MQpRiVO60tcqiKvVWrn72mdYBTOQu8UyBWLw65AWTBaMQceQ+BxnBzsjV8
ZM19J62rUTCbGBHkJy00uU4BH+YAie/on/6BruwodHWHFzlxwz4od/V1H2sbGchV
t6jrM24bYAoqCz0ALjAwhqnsJLro9cO4tebrZLvnnlbfg2nwSBjlWQwb2kOkITrR
p3pIWYQ4pAGYgq9/AoT5RiWyEiG2BeBKfhWZYHcIzdAIDL31AfEFBSiDv8JfAHWM
Ix6rkev8m+M6NuAUsZwcRtww2EzaqLOzEnR7zf5RhT64tdH3hX23WAM61H7xd2Kn
bC/63lCLTBPf5jB5Fq39U/91kDupbVBavEA008Cy9+F5/bG7Nr/0MoEFAu94OK2K
vJKlsbB+TQwNBSaT/ErIGJNOhbb7gQ2dnAL0BcX/vO59fVehkhW5TZxQJ9u8cMrD
rID0JJewuKKg9VqNEMwm41lgsZvOy5MIf12ZHC7rHkmqnSF3HcOPf5imndMI81MX
NLsTReUEP4vPtC8jsImt4X5jw6KzvRjxmrszw2rMkzysxID427T7fJqWPCi1smuc
9+kGBhN5++bDCEfTFqw0Wb+H0qmO+pIEek0iYubnSjzAGVjsQgjAgveA0HlQuC5L
qeVbfV8MbP/lqsEwkhcAOT9Sdhk6c8PTU4fMfMJV3ulPT2sz1vjuRvEGOYZM5oCL
P0vyBWwa7iBCkX3Vf5cJZy1Q/KDn1ye3JrLmM+rB40EaGjXtNuLajiIpxXhvhWqt
S0RdgtORJElo7bhVrFHAYAx+24LA/nt6juMd1KZL67B7ZkklRWd4RsJ00+i8m+y+
OsggBDRo67zvMGO+qHic3VT3jdm1UynsZMOsejYvkVRhWIInfJbb+lcD8Pp9Uus3
O8p1WjT874LsuXE3wah53rfTSAv2Ck841CvYz9+AsXvlYVzt2PETMYJDr26s5Rag
6u8Jh2QwpNkWTzzy2XMSw8LNoFrN90pnR8/wTX7fHgaRkZa/N8YAojZNqn9SAEZv
QBrX7j4wCyWtaYPNE0QCAW9E18hANP8zZ0+s7EkmFNz7ltD8607GELN1AUokzY6J
N6RucDAAVcC7pqihsGodYtJP9SR8SCG6LWn2jnQebk4CV9zEYziFOvgd3mm52kDK
oFTG6t/kj7zxhXc30InLQszC2+BBSpilj93OBhtTV4WPBXkT7OmBZWGihkU/LbOM
xWJlEbHlNBTXUhYn2f3owGKqshEVsSzEzmn9mhK0YLjEVdHjTCq92XcmbXCWhkMk
TeSxcBhd/V4YvMJFLPBcdg7cxuwBhXp7V8P+Qbm8SeYrRzChqxOaGRL+G2ZzAZUk
fb1NkWciNMpKrWpk1oHBLx9ARFT10L9ysOkWIJtiUrG87vMasQzMo4G9iRd5L1QF
RTUXuihfhj8bJ/1/BChnKf1YpR1BUfquLZ1p8haRfCHTTkBLBIkxB1RMLnvhsBJz
N9QfcxV3IMTXX77k9/Sn3JjG4r0TDjkLuLOkZA1cAl59gA43yY794HRwIUhd1I+o
ROFnm9G7nPcJcfOrcXUnaQ54G4Qh7vo6d27dW1YMSUIFD14lDay0Z/FxDUBQx2uU
I60Wbet6cQjd3OoOHg2cJxzaMuN9S9IKqtN3c8HXWHw5GopzyVTnau0JMGxtY2ag
GQxeTWvklbmcPi8uct7RPPXdyLGP0w79pqyrTNSkSTribiHXbnHN30WRtad6Yov6
S0f+ayEnm95fUcE/qFL0fjJ/Ol9kepjDx66BtqUIF/qXPdgVxRgXoQtUFwfSHHtn
orJNsBNMEX9t3sjpSMNE40bTERcL9KQ0bdhZ2irdtbEIRWMfRmsEO6X8c0o8z7X1
WML6Dlxck8dINOifl1Kd2OEJhMkqiN+zzyT8BAzWC1ZJ2IlJnzT69Gn8c5yXCLFR
mWGVXWb4jCVhpm09XaqWJEzknLxCr9XpqkQSV/1tR8sxM0Wjld+k3Bb8RWpYrAZs
zEhrNjdi5sZmGG5J1VP+TIgfjsdRM355mgNZreWxo9B7nrVsEIN/RDESGh8J8Y1X
UDbe6eGxxIPCEpoBEZjS7YkWBnV0EbC3aD4a4htL1e8Uz5B2hOg0lBJkAXFN2jkp
dg2hpD1+ets/RCja8do0Qd0hp3/FubpPnujVMG/nfJcSKnj1CmAB+HxZ+NrKM1kU
rsV472tu1EH/9w8AKSDPnL2B3KVwsuskfKjWSiGFQL4W6tkHww14OGmCUnNID6h2
YM+9KhFn+VfhL8cGZPU+YrXmBe0KeF5f8J7+BE8Mq+7/Dt/RG/wEvjqDt2AiV1gD
JpBNGZg7l7f04w0DrZBIkUvjQ9MTDTtIVVDUtOIBlXgiwF3HqgOX77tA3ivzprK4
zpc3otQITyv8UPzM9mtNkgtYuvlGopEYXVrb3S8c9H81hMRducTLS/sFCtM8f2lo
1MmncGC9wQ9K8SzvwlQDI15IVz54udmAk5zqYpR7aPLAm1pCeVci6j66H264pd56
2QwMWJOnHQUAcOF9bq9TQpR7QQJeewm+RNxNGwx8HyC3TW97qPq5FbFUxLZkoHUs
GwINeAPhKsD7baw3YVi01BZ/3QAWJKZM4I4YdheAMauKi1/AjtIO9PvpWPxYQkTo
HBwDlPlm2YPCa47tUwGnrELBO2hYZQCt1WdOwrYIJ8/CLPayWZq+N+WR8uDR8emD
UyoXkgpfby+KdBzID3LoIMFU0Z/GPKaJLo95/VuwiD250m7YMxYgKuCyCs4jXZnP
KFsCX8xXNX+k+jXGTxIGv3QVWuDI6O5xxyqyM7VnX6mXDuO2v8oPxPSm0KHO5EHm
dOFD5Gl3zO/0T65cF39ruDIVSm5OTP4hNi3JX57ViisQ3x+XPClLAqWuM8mhWPJn
ILmQkR96Zaj+f7y4xuB2xJAMbZgI/NJfru69+9xt01JG5yQV+aOfKnqJX3uPPAFw
txF9GQjCykBv3fb0cM9JQfk/DTzzB9GR7qAI+/BLXzm+9J2gaUsAJHU/9aVJ/LfB
x+fMaz2D7VOCwEP9li5W0sX03JSl+5IVqJQ6OisFQM6Xt+vU6JpoXR4PYoWgTADX
RDZr+bCPM7Argi3gWcv1ELglFTZZJvEess7iFgsURYI02RHaBwltZmqwhnRQPIqm
vWjwYPvGlECNyPA7wiRKHDUkfYqS2XqZPYEBJGqp3z37dHxT+3dskIfG9dPfkVVX
V/NKRVb9RAyjTvVveafynLt4LVshGi5AokMXubrOGE1Xf4zdn7d7oeSRMG2SZlJS
Onnb731oD/PY3Z4w+ESQba+RZJtteg8TEzLFBq59eRyDd3gjZTxcWup1JR4vN4JD
cGNReO7lDeY3tkYu1Mx93mg9JNN/ffs+PpnFM81iVyIcHZq17QrAwfcYAbbkPWl8
lALFaONfEDhdB9IM6UpE+Y1CfNiZskIf5Ls3wCtqFu1LaOZmTvg5knazb1gkgfz9
XH6o0Xdt/nerdX4KEJQkQ3Itw7mXFzeCtwRX7lUJkOGfnQ8GHA6Sp9IKptZyStha
HkadwLbXaSPkq/Dxnnz04zZd1veCTr8CqpkTYeJDFTN0LGRuWiuxOdl1n6imrNU/
j/rBG69VN1eXvdTOdjaJj8q0It3ZwnfPEdnrpYv8D03apzVNgsOGQB62hzwV4iFX
O0kHTVywtMXIhFZ9f4fWIgX48QBJ14FpjMpZJj8tfsP069oK8ZbXJgBYqOGYiVQ3
uMEHV2RRMYBQWQUasePLhE7h33NG4b8AvJATCg4nWCj6ozMh1Bzbk9Ow6uJbROLT
LvM27AmYk+fKv417mhe+TMltO+NKbEJf0rkPMyOAl84R3dYV9UGsnFv9gYb7acEe
Sfp3DHh8TK0Ti0z+MJtxZDAhh72W9MJCH+hz8Kc1qIawSvob1CyMbi78gi+ndGAY
3Nu+pPMRQ64qDfvy5kVLRc92HS1sLcu7kuXmh5gMC59oTL+LuSXk0xogycjfo/e7
+r6uegSE/+VyHLvGX53WhQV214aRT77bY9aDbBx82Z678ov24dDXSXrCRrn6qcDW
T2zsf0FXoCjAMKaCXLrJDckOPgcoZy2Lx/NfW5ohMAhpYSlYRAK1LvKxWy5zWWL6
rEGYyhZgTSso9HX2q8m59obF2fRctPEBrsjh1B1MwiNoGJFW/iYoK+y61QUmYseF
pLYbz9UubfYPKNjggFy+sCLG4y21ZZJm5e42nWvLncukMLuaIrz887PgX7W73zEM
iB+b2buOCdNDeIjfMybPc0Y/kFjNvEnq+jQ5C83hjtKHgU1ccj61hStH5WQUvZuE
TASJ29Bl6hjBezB9W5F4/T3JF2GfQzscftJfcQaY5H2to/egRWR/L2rnYitlR+JN
OsigcdfC8s8jSv7Aete0K6jWcLD3EsTlxjXcqeCBIiW4rrwCeuaaLPIa1q4roHp/
6u4gzFibkz8IyqON9c5mWdfg8DxAwd9Ytk1+gznJtwZrgASki40wITv81MZ8f3mx
tanl4tGNtxGmLD/llXE3aiGG2Ts7LbBzMdmXrOH7H6IKIf5B/KW3/JLeLQt54BTq
z970ohvTJ3Zml3Yp45cJJ5h7obeAFq7jYuvjcMsH22OWX4cpidDfJ0/kuIA+mYoT
AxnrXhVJp2qK69EBveerEH6vcSow4OD2jCMUK+PL8tw/4hDEka9Y1kozbEv7l5Bq
yCFHYisgO4TQKTis7da519doZNorEodIXpyEpksxT0nnzkz4URhQE4oWZMXsSOry
xemDa7lTLxcQAvxXgOCgJXb2K5f8z3GujQfH3HG6fGyLlb2r6M3XhQxvbINFBaKc
pNGNE1/3j9L5kNMcFj0PdclnYvOng+0mpM7gfg3wW7UBBPzBp0iP7GgVLosvJBpW
ZDV5fbz210JXDwhjBAe8UxA7k8XM8Lp1tMfHFb+lIkAzvJ3qwWimV6jUvRE8tRfD
H4ygS6Eddq7gYSTNA6j7lt4hlS9hYugLWNUQJYJs/i6zSDEK+a/h1A0JhXxl4Kjy
3dJ0cx4DlB5YgejlrgDXma4JqlzyspwMFkioUWGDOl4M2WRKa0u0LxMzgMCYkszR
7HANvCpcIk4BLTNK3lIfMcKy607LFdiUt2qx4viMTs5smOYJZFMf6JzI5m23EObT
geU1p/YYR6qlDDGHPk/McyTFzzlFaOTIfe8Wn6jmrWJPQXvQx0kJs1sQ9UpJxuGm
mHdOqH94e+3+LNjoAqkYRd8HrE3ondsgTDur88c/XyxCAx2A3RplZgddLwIAa3cy
gZgF0/KckQs4R1qOnyR0PmBdEw1L+gFER2hJIrxJV+i1yDl12MXvgqQSL/GxqeHM
R62RfuLzbjfZ7RVaCi0QCJaVeUsNilcMkTlP1nS+KazRZZUZbugPCcAluF7zIsJr
wdOGv4GjZg2jfO1x5K/d+Cd5OVY7wyKouRmUVFgxQnZjHVYf6+Q9DjuOpStiZ7q/
HBu/yo4FPvADaiswBX/ggefBAnyy4gcCTxR5aQRGrGVRP55wmnJNraO7b5zsp595
m+gSfqeabDvRm1xa3I6Wkgx4ZLLZftQt1VOfAyOYpa8r6j7gUPoG9Kyt6AQx2yKB
Bcv/61rGS5r0o8L93T8o7txH6V6ZTn3ABqeAcqyB7N2K/YzAyxBr8UimKVvd4A2O
w/0YFxorEgv431oVJZnPGz6tr5fpjqj7OD2h007amH+Jc+E+Vq6KjyneIsfDsHqn
wEAM6GFFU2Qf7KLwlVrs7ALHGQ0EZFwrDr9U8EjRR66KHD5LO+D5l22Fr4zIb1xT
LxoZffmGRyOOaBC5GJi33aSTYDjQ1yfn5wV2KNinpOF+3iD7UyoQbik1XkT7zvgo
D4q2URcULyHI5sgFvqxrh9oaExayN3LZI7/fG46WW+OhTtLEGCte4mwxf7nIvkMF
u7VB+/pJri80QHF3w8exFF+ZoxRvSJv+AIViDiRq7d0MvMGzRAMoxeb45Du2221h
Z7P80wqigZDtnqUGxc1YzHBgwB+OlXZcpbd5TIg3/4XTPZAXfcUMBxClwZ0uwdvF
YdwIqigBVjOPfUMyEPvj7Y3siYWC3uvxS7dquPd/zDXeetq6YoCNh8WMYSz1COj/
1tLrsaiJg6wtsQLMVpN2BdGmL6Nkn31vV19UIPya8vOzwHYssFloeZjgIl/YJSdY
Rmd9uVbXyRGe+FlB5MbTnSV8o0PQ3RyfU3noqcQbTlouVB+qa6cLam9NI7oL+X3f
kMWyDuzPEvYR+vMewVNjIaw4Ltu1jlJGymLD8mH229cCoJin3wcRqIuS+L1gy1RM
9dYh5tnVYMXmPmuY8oXU7NTrLE/Ve/itqpC9BCtZS7YJtEqWwWjrVjJIV0miuQWM
Uj1FM+CvixwYRBnvX8cLXQK/bk2or05Vsq4JvbwfhSk7zaM/XEe0IOEPg8PqUJUf
Mj8kI9CDaqtoBIMLN7VuyJ0lI6cSguFkkrEOn/MCbiGIOnJB441uI/H1WyELYexJ
4QJyhP4OxjQGc1E1PoT1K0f6hbfOCHu1yk60k/iqlBIodNdydidfTlYs5jwmf8YO
73WgheH9e4sDTekvmWvc/Wda+UnRCoixrCpGjVooKv4eNdWwHqDBKPtos9rn2oTg
1bUuLSnNjgqZ/4X3Kv2dh97BPCqhrCkb+X6UF3rErwVJYRjVaWogEPUgZGhXaJF3
0XWayJI2YrQLp3nut6UyhcfkW1y/CTcagWblDabPu3Vc+7yyyR68FXoVNMpvsABe
766MGOoWBePNEmrJlxBWJjfB3Y16P2KxefBInj0I1IPivOZCEKZyN7pt5WA6q2tp
Wyq8/k79yqvB0DkMb58a2VI499xTzpyvdW5euCvXQ/rlAW2hWWn21WGWoaBvBI/s
ZYSkmRr/y5EMkSPjzENUDPPfUxqkmwFwQHtAMxdhQJcs9IIQJaolQAcKhcGvU6AE
4w4V4KOg7DUQakEIm71MlmF7NEwHAnuwLkN8luetJY5nqHANPqLs1T9Uko3ynlXR
ST1d1Z8tLusRvuKaHP/Ms3reH5Vfk049YZFxFbnG8oJHmj5Z2eVvKKE+1WWR70U+
bwHXwc/HbEhsjg9xCCMdTsDMLx192h3rMoMiUM/RX0kRz+xXD8JpQiybWnxIspdE
wQfyPkvGHI37cr0O28sZj4e0lebJ4rK+5bZDg2gXTPwnCkwi1BB2zuqoZ5p/cx05
rOkxI4A6wDxZ6KArxkvQvUdiOdy5qoSSg187SVyEUy/O3njX0ZTrbw9D4ItXvHLK
QfTQu4A/4ejyPG1+OP2cVMd9KkmQgW6DYKnnInWWidBxr0sWictvJpFpeQEBPgHw
VOk2yDdX+ivPPpR6WWNZN8Vw6e9V4b+CHaJj+wTfPehMCrM7Y8BxRmeS6MUB7SQi
BYOliz+avgBVcaf7PtWN2V5l2/EF0ccBoD9WiMHM1STpuTdz3Al5nm2BqNNtsDoB
0g3kAgP/XeLudjSv1aRK9zvLQ18SI/iH75ul4Td1WIdIwDWWY0DRLmjbkikTlr7a
pJmZRVxG+ANcKdv+zgcvPnmgIwM7N9uM06rhHiiaQyyETiLVW8uCyQRNk661hcXL
oO7dvN7Ov/1Tl4/53Kya6Q==
`protect END_PROTECTED
