`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoQTPVaiodxLx+xZEbe4sTEGHTAM+eGCv+vZNdRdtYDa5Dw2JsGSe8ljUpywDaAx
kITgSg8PGjox0eslEXTwxcTniGdNse3ii8RQS/lj03038iHhPOjX1CoS3u5O9fTu
eCivGdSztSV4zDDKRmm0ZYDGwUAXBnt8uMrPrfc+Ic9jRWEEdazSOZV5VzxrBvNK
ZO7PpdL/Sctegqgor9LgUqs7Y8zRniP7iFS3MBv3WIHGcoABDJA3o324z42QTvV8
jT999k4+0M2cL4oZern5UWOWquxsw8CbPUQ2IFiZ8QuU+1kPW3wBJo3zbA54cdW1
LXjuH6ItUzebtYsIGBf8Fdby33AIuAETZ34iYmBJ0t1nk9bXz4iaxypKJL3hVXXw
dLw7a4tn5kwhlU+1uEsEyANhWmVDcIfrPnD/bGj40l23JUHWlPl4Oef430KRJSLF
t6d8FaYGFOj44QfFS35Ufr4iF5m/iZEQAhkDpwt4njo=
`protect END_PROTECTED
