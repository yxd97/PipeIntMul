`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYFmeNfE+/+7hkFqBm9YTlkExB0JbOmKjtTx4kxhZ6HV5LdN449WsXbQYOVoorwN
UcH9evDHGhBfj0VmEN1lniAkNvaxoRDql2e/JrNyTsEZ3wtegGsxbQ+cVk1hav3Y
c50+NwrzbaHDuR8SiUlaqLyo1+FaHqFS34eTcaGlr2zgOPda4bJ0XMajXLJbeR2x
gRxO2TnL4AFdeAyU90S+KP/Wc/GiLL+6vABIjWX82V4GDrsOCE9ivZK+orFKOUEY
3HUCVPFzHuvXB0GWM7Rkx7h6CodmLLFw/8s3lYK2K++BcUr1JDisFXgeknvGIMRZ
b1YidifllsNGOLm7zQcsb5hzQszYfNBMr76dmVXDc3yNg2Nj/2pE4NaUssk3+gxk
C35A6xsRUyJ/tkx7qmx/wfXAPeuMGB2uKI9EfqLLRAgjQQO+TE5IZtgw5GURDGAf
SWa3E+DERGi/aOKG1kbjXWdNxxanRXu8TnwHGAJUJHJvASex1U3GQ0pGkJgPs6ic
EySljFmFWCknWX9gGPJnqR22PN1KAsY3Prlmsu1hyRb/cJDfRO7C1oDIks/C+sjw
hZClO7xftSj215Xjx45Q5uy+Bfz8cUsRNQmGxTU5g0Au4IuBJrj7IZzH4DAf+2xQ
W8vJkQxWsqhj+S43A8hYofhijmmXVE5ABoOJhkqeEzJFssSeWMDSqxSUBvk3BLvH
oe6aeVMlXDFqEnboQ53adIVDB6JTl9eBJd5iB2+w1oo=
`protect END_PROTECTED
