`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7zaa2yj7IDsIIXjlS0ZW1tuuJiVU5IbXHP92/mmcJ5SwPDUHqa+BEIhi6210ItYZ
osVxUNb2+WUk9wA/+zXVpM1zF/LfVP6UBPKDcID0sZSPLvVJJDgdoI/iUCXplE2Z
dz5SlJGDW1OevofVDjgdzKs4jugeyfStG+YbsmfjVl1LfiQZbfv2+0hMO3NzznNS
JHBAASWIjL4GESyNKgaWGIy6/qEERx0VfwDMoQr5z4fKKNVZFklZa7SVDs/OIVi7
QPASOhBOAZFSL6xTNZ3If+Ez6YccE1RjXbddJh7VDPOG0NEg889hLsIZNMIzGWr8
FqKHmEx7NlJzVyJuTUys2HG4NBd/x4HJKtNXc0CHmbl6t3cVW4d4+aucxcWaDOWQ
sWvUyJ0QqFPxZ+rvwrCU8NV5kDKNZeZXh84xcgjVus7x8qn19X8ai/+orjxKudOs
lmtlMxEX9i0A7m8jJshR+cwiP3kdrjtMa2JY2GX2Ur1K+E+eBkaHAIGiOyt4lVpk
Wg6yr9fMzGFDYYlf44ib33JiNs+tcpLEYOM/A1snR33zu4d2vVDpO6nbBkwdXAQg
XP7QpD/qvJ+rvODJYnQl30pxdmzKwLoUd4cMqV3BC412yjX3coL9FmgSqFP5wCt3
i4o5UY2GbtrBSjd9uqMAVpsBOVuNSCF4e7/emQ5NJaIHZHiCijhuhX79BERD7kv7
4f8c5UtmVdfOF6zxSzNy4tTET5Y9ldFn2IgU+BO3b4+01ay+FXnpwUuBiKspkv2V
bIQb3c37MqRk93wiHe3R34w7ThYOwUvvTorJ6x1quEdKvucwl+bcBlqdZf2f7H3r
4ixChC9z5qplokPN+JKpJE73qCOzZCUzCac4b8WGmxEZMx5txCP2zGTvlcA/+F0O
rS7VJU3z/KFB2+NCucKj0EvJ8fhwB9gUEY0OnsqsTXqHzyxTHmF4LABLcurDekDS
pk2RTyOED4EmxUhDQNTDmG3B00UWuDXd3ac7PWwcw8EwHYE7sZEZOqiUJVKUjQbJ
`protect END_PROTECTED
