`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L5ZGKiDbpeQ9Oz6StceTgddI7lYywuErjfAg5ZbUpjHgbv13WZ5JPEPv+1brlr1X
NxYg9dk7tJgFxgE7aJXLNSjeJMLKPDTeWzQFysCgK7SiAcM369Lr2ysRG0jBkF9n
39d6HVnsWPkJ6hdGozMR14ze7CA1YnJdFe3eTjyFwNr1bQkswJHF8EdP5n0F9tLa
nqqmstKRVUZCQ9tmmVvGIfRZYeuZD93AaSeEfnv0cPdm78P5WeWAF0mH9Ms8BmlU
25CQUub0HxcXDLGBGjPrxeoogW3Qa1X4XvNpx52pbtOKKzKe43g5WrOLf2mRLUb8
j3n2djsqcNYC8Hoh01/ABtatrUB9cDJjd7nRjtfG1NRC90hJMWaY2ibn6n9/i5kB
5gQXw/olUt5GteBLl0tWY9YMPP34kQWso5mUrTyhCyHxYvO6wfMpQtICdfzE3QUT
DR1CIpr3/X8XfWkEOzkNSobddcI2mIMe3sqLXC1ZwTqitBqOWufiL175+Dk4IIAH
RRj7jUF+73ebjyHvcvmkxV0bexdI+eNGkleuq/RDmLENGh6uw2DfM7L780Gr1w0o
`protect END_PROTECTED
