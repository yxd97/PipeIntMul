`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jk2NNp9vxEOr+vvFwMtHV5zsEfNSemQ0nMtAuHiMXwRBUu7DZffxh2ujodPKDg99
N95NJecxywkHS2i/s/fj5lYbZfWrdq1dzEpEpYSggZHOjNyEs+R8eh7zHzY90+2t
7E7GHVSQaybDwJ3kbcsi/Yh6Iv93Zl8P5tige4XAFtYYAoiJ3tF9V6wiL8swaoPQ
+F6lrtWpt4uMS8xeTjOJ546FE7ygFVyrLs8BIYFaV4zchKUOHCJlQ8lFfBCRAkeS
mqYd0WGQCc3Sixrgrt/4Po8asumNr4hYs8bBs6FmglcI8jykpR+wnfEtM1j0M1jr
J3bsND5F5PXt5sCLO4k/x0/adVrWJ1+di0UR2RbhKDcAOhU6YBG4kcC54HsIJ6Kz
UVgQN4QF3EgZObYWrEZNjtB2j5pQXqNN8AyNnhFMKLCsz+FpTmZk7uv+nU/xI0HD
hdfkH6q0E8mkH1miWZgR1LH3YYfxGR7FDxuT1iRJ/MWjPLqd5jCHHI4+0BYuJhAp
dVobO8uMuKfS3xWWDYMHeNa/coXDiJrCSvH8JyLro+RbQ3oJGOovY2NXSYV63EB0
eXPt4umf0VKFTKJxpY4vj2GczA/Re7gdGWy7VJDIRpvGyG1jy3m+EFCgRk0dQ3SM
RlT9jPK9HVBZ9cnDZTweBcT7vmAKg/idWNQRf8m0+JXTRk8/3Dx9pR+AF30JYuiK
S2pF/XRud56qRwsUMrrvhSMhEdeeB+I+E+lyhAfrxgHRo9d/btxrpo98bYsvjMhf
h2iORQAPLn78BUw2pavP6nhS5yQxK/hevzgF6mXUuJaL9EfGRfYmNLpd5vo9lbwx
kU7VPMetU/n6OH/jrYreilXPXIL4z+QHQEEwiQ3w1FM3now2hXjw8tkEgfC0bDAE
chEnQKodCv8CaN8tUKJiPHnls/LxHVcGbKgPhr+sSXFNiTa6rhwEB26h1slDgsyB
I57vrKn9uchhSHg6P1ScY9N/4Iueha8WVdU4qjow3FYZAuJIwr38mp87d5aFeHgx
QG/UCY4pMNrP0GHpsn6pp/k9/3QHl08IpwoCMW9fyDVRZFd2XsPev1RZl7cbKz0e
tFegksQZnHuXlqNyzubNoNcnKdc7hD5J6TMOcenoWZOKCr01YrCLkDYIIpkerDdW
KBp1iNFa7JNeGgTsTj8s9NRlK+xwHT1G/RzuO1UxP6vTc8B4rjeBsXHCiQcuzQwB
GaFtX1yILTYRKj72PrKgdXdJ6oK2BGxs7qtL/PlRO1MvdRVSIpxQK1w32/RToGZY
uUd6QGd7OuE0J2ErYmtZAty2yS35F0qgWkhmjhlpwkENFn8z6UPWFopxMz3E73DE
zsUtor7PxeAUA/fG1fRAhHHaH7SWDFAN9HnI86XPZW+P/BnqzUUzHm7NanzfQjpu
n4OLwrgEx3OY2f9s5wXD8AxGMsmFZtNpNOKxmqHPbwa53Lv+jZHkfp3+Hl/6PkUN
SFR9QG7/p4RW0G7p4MaL0ZRbTMmttbtvQ8DVG7KJqWc+ttEddS0g0sod9FJ97zDB
CEHk+P1MgNR2JAIn0x5TKMGEI7Boez1pr0CijqI7l1TK0WyXS6S3S6ZgO2oB+H6z
Hzl2ULPYEbwyGTCCYDqPqEa758Wdx6ON83nhmGgOkrT4D5pz34DSN09ZAXKTp1ST
PyCZLMPB/Q6K2n8pzb4Ca+AhWmSvLUgDXFA0QzqlvOx0HAHXd9+q4eU1X8Yl1czj
JS6e5KFd2OQ7LKI5zwqS+rF5+/1I+t8Pep3anYfzupCD9+Oh3ITyz80MQZ8r/AtB
b6cbIzUQM9RLRhwLlXjktzgG5MwUC/cFepFCZkb37W1hkI0Ui2ul8qN7AD1dvEqB
ucyJRenskkSS/xtX2MEkm4xOgmsOEMpg4UkD6Si2WZHJ7z3/Sy6xfpJolFqzb7sV
o5exiIpVam88yow32xFhS1A2PRpYpzv6ZIEJ0A/k3uRq74eCRTf2DcxJidXnUcvK
w+17XJALOQQ5dv/127SiLM3JpAL0d1LrU/tNTXuAA5HucBZcBXeXgVDpiH1oWkIH
+BhUeGkI/qbAv3k8HI0V2WhXPCMCiLGY45Shw0WUyAPOiHPbceY2zdZQwMNqPoaC
9G0FBfQzJO+PpE8aDZeGWF811gobBM8MlxU/t1bz/b0=
`protect END_PROTECTED
