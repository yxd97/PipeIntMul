`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pd238gvXaI8OplBDETrN1Qlxmb8BibabWeseyBkKzBBjYIwgmcnALRbXrUIgCGX0
1hwEmEFO6e18YCEBwwgRD1Ona+scbJZWmmJiaohB4nC3A7vd5z2U4cL1fy/nZTqn
RUkJ+GiROCcF7wlkmotEmxDpEThVLRbdT4BgiZzbt0JhaCr2Km7jf6dQrXOrpaRc
XFs6uE5CJfqWPRPrqB/lKs+7/T/xw/fWKlEyZan4gspDjRNaz3sB/h8p18oArtwT
trYvdw/elz/fIlXNoTcXEaYP/5jl9boEHepvXwRCuLIB/7/rBYyaiiVJwX3neMtu
HfDp6MxzB2Vuo3z7iMcdJMv2O0HUnqvnoVU08v0+GxX/HiA1ql61xUkzgbDFnpz1
5Ot0gYhxZY+hH4eH4J5qPCXI4qtY9N+9yShcqedpBLMYCwiteMLT2pvnM74jaXIq
6UM9ulIccdJaqOWkPUXBJowfbh+PoZ+1xWMYn+EeJ8e+flLEiHC+AEAWMj4nTxLK
`protect END_PROTECTED
