`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
agGXkMiHzYD5z/0+YZ+4ijBAs8uZ6yZuYWa/CclSIy8bcYYcNOB5OhsQXc9q2TtG
4fLNbM2d+mTLTLFKo967nYvARda92E7R11VABYuU7BSHVQOZS2O0qbrEAKMJOv33
poY+mNkN9bLAHSYO8Z02QM04bUS7I4LByj/XPdWFZ3tjpI5ZifXN9Kq/CTJvukrp
l52lgupBmSoExPpz1UGLVs3ziasmiSbOcDMWw8g1GZrmLrEgPCTxp2uGGYS760Mk
KnVQX8D7BmJmqxXYoVRPyo6taLgkJcScmL5cX0crgBAmYDs/imfz/nYhic7wXBhc
VjB12sDQJRfLXAJK2BcBXnxhwK9cPS2LhGHMDnL5p2055GaDFcTmXRdtlVDWZtVm
qNsjjlkBJ79emhMwlCt5gwIcxt5wtqjiBj8GGM2KupWazY/BFqIAFd9QQpXnsiFo
FjRWSvCd+PUpunbcvlq3k24j9yR5NwekJg3uvsJldw9urNMOS90OjsO1wJrb7O1i
w0q11MX9Y7R5zTnyfpmWYy53NXMztcAyUNjmKJl/87+hTLeumr4UxDKi6C8za4CB
dU3ZzEDFDrwQPtpfN44R2Pc6J3ILmrNGC6znL2ajyGiMZ4Ky61Jjwo+Wm36XZGy+
2wAhzW7kW92d6pYqjq3J3jT/+GBCJIGF6JXnUvOvszg=
`protect END_PROTECTED
