`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3ikPHj9QzFUhwCbw7pAiexUVvy+2jQs79phaQap/dFPpk8r0YODRtH4vQHfAb2p
kwwvbjWKmKjqgNfmDz1OPjaIXfOQqVPLgDvzlj3hgZZLMS24KKD1xTivXOmuuZJW
ndxMVohzDyA0G54EU/z3iU+scyxgkUum9rB/W+yt6tFK6Ko4aveDK5qTgMZ41SSU
ZPtjQK5IqghkrpbGQMeR8p6kCN+MCaeoBvmNoly02oPs7tF24o0PCY8AFeDo/n+V
A6Els3uNCqH12ytVuJ2lUyHSi6GsxWEcDM+Ujq94ciRc7WCnrk6uEqTA5zMP81Dq
DGOnLTNW6r2VWmmGYiXaNyRT/seapJ2b8gMEXuNH1I3Q0fywdRjFnhp53t+RZ1SL
`protect END_PROTECTED
