`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JpsHZx9foOzerwW4PcW/Ut4RRD6lb230Xmt7Z8+ZqVA8FNI1CpxOweYO2pKxwxig
gYgpLxfoeGoM1dMu7rnNlGoQa2m7I2Si3V1HyvFCuWrJb3m7RIn6iCovqCbslPv3
0QkX91kXj1CLaaie50apCpzP5HCkOD5NvgKfxskQHM6+G1JGBlp6AgV4kId9D7/A
rqxCbLGzSPlXa3hCBFWCPxweOB4de1bmrFBpZoFEtm+t8C7ooUAyiwq7N7ECNOmM
7/es0hP9DrJNfoFyssAeD1bw2x/yhhEcKpVbtOTw/Lj7ea7WDAjQpdBzOvl6kYCb
wmOsnTssrVu7XvhNgOFhzmuIUa4pk6tUCLpn8E6HDajA0WQqFt/c0Inh5SkHJotV
G8O9+3bmbozFk7ftfH3SKTQ1moUzEzKjPzTF+vYJpYM1MxpGaw4lmBr4cJDRo09O
FXGFMyiMmg23miAnaqovfZU8gHMq9ImfDVfEwkA7pSU6uEbmv5IvS28nTbHghsyo
lWvqwZMicyk0uzEe2EO3I1CTvKc9i+nG8yCPziQUIW5E6rVGtjsljoiHzNJgnzVC
/5Jrbm3N6fN5llnKFnOs933khcS9a5FjqJGAs+dW+ZlUdT41irjw6X5QztrbYR91
/CRHsV2OIOieO/wcBpF53QeZIbDEXKzr8nmNwVkyg3IuM2mm6/LfqBZJ2SnJSeVP
7vYn74GaRtPGPNDBlTni0FvSxrb7pl28LTO/KoFeCHT7lOXHjQ2bamFe7rAfRSV+
/1mekymYUky9aP4J2f9cL9zC3s7eEjGKPPR7ruoa5nyg1bMTjP9eUR1U8/iH2mQ4
cyDamwZd+gxlGkYJROenqPydKykfVxlronkq2uBB23GeGCHH2W1r/JjRLWslh6TW
nk+xqWuFN3QhowsLEgDo/XEsruxEen3qXMmpoiWCyxzNQldEJr+Vr08h7Nar1WaF
uQ4BCl0k8lvKWljF6v7nvCdqZG5V1YDtvgG2BY+HFFntOKG/akBullux9bmSlzGK
Cqt9X/L2sBqrnnMajairXjrBbKF6MtXohUbNkJZHiwPCYDaqi+owPO/bQkMvNr/r
+zI6PHHZvFmsRrR9B7Bwp+m0ohsmXJv+xYYwrtmNpw1pyNDb3aPkGzgL7v7A8nrS
SuXmpTiiWl1xImHvaptAOoLifCKTDxnnZroUBqsKaTeRY+tkrUOFI0ujRnrciywh
aVQK+N8vBsrJ/I7Nci91iMimo72DOaR4vV/BTsQwGt2ABmqPBBc0M6y5G6Jn4GD9
kcO77Pi8zc0ewLCkdsFsPfMQjfvCwAcpwu1TPppgF1jz/7ua6P/4INuyLtwR1zc7
51AIUM4Qt+RHjtLTMVjdilGI6jZkc9rTsHTTiVp0dA4tpxjRMhumbbrJWV46pl/Q
7kAZsAlBWZWGPeMsNQAquaHR08qcOt4SDFfLLjhpsIudelywgQ5Uojzx6oLZcy+G
t2ICHbmcIsmzeXi8gaxYtjc7Yb9zl6Oz7MUqQPVLXs4qIlFIgi3/JoVOZeHqf8mL
JgL2ffw4j73jjhiJ16ZLxHSIKKmAZOtuH2nQir0/QxC9rh76J+SAUyqnYifw6oV4
9MAS5ojRGRH+zIMksa9CBvl55BLfKVa/aACdug7S9i+sqOxSQ+EQsR+gC+Kz7qAL
7KkgzmJexj+ygK/EQjrLNErISb9q06EoMWWaljCQ6LTtTe/Ies8fIiWxECEO36J7
YjrhTyjC8WkdFsdmXCWSPGaYcEA+8C0xq1jCV5/JLNF7rI9nCdKxPdp7anSQVKtn
6MZQsZQ8yxPXM7zptJbhQ+oA7TfcOMlhZzBNW42qeguFrzHy1KBnoLhakFig/n6d
TIaYg/fkas/Ub8N80/OAYJvHN0wX3RArou3FoF4VKoc9E4Zf/ynGrVLAxgOoY+0h
rDfpGetp/Szui7n7eebw566GmBdWq1REykd9spGXEAeqM26DIk/WHrc+7BZrvqp8
NnDCNQvvXicUVC+X1zqkDIvvpDyBZwYUjvzvPRSHLQSxtMJcIxCzhzA59Ij0Lh8x
meto9v5O6Cp1h+zZU4BCzkztmXh3Ym56JBkkJ/LLQ4Pa34v/ftCDSAMIO7sMtVF/
8roUMFhRvl+DBgNX/m3cUZZ1t66z+1ISF9GRNEw15ARlMralm3a24D3ooTstyeIy
`protect END_PROTECTED
