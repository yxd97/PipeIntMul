`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e+6+vW01lEI3wkg3h2zxVcnSoHs3wiPNxTVZw6EsDyGG5ClrCKqGvK5z1gO+7Er1
EuFQHlv5VLQlUduNtDAItyrO0kjIyebVB6GLafKLwmw/qz7V+i8rTIxB63k4MFIz
j5SDflaq8/KEQVawGV6hja7MKWHAc8iDNL0zP4ZRoh+W8nNwykeSqbpkFc7xTG/8
Am2x1pMHNQj2PwE7k0HcSsON3ZtMGBhIto0CLC3Px2VO78AEGHat/f9Af4QSl1dY
ZkEumr4gKK4cLPPPg9zVa2QJdLWZ6rtYUN9wbDjURuX2WiIqlAR7sMp3H6lZDEaP
GOWdXyK8tpSL1ek5LPdUzPo0BWjEuNUMblTEKQzS43ibvIAOCGxjTDYoUKhN1O1n
NA9w8WoEIXMsv47MYWbnLg==
`protect END_PROTECTED
