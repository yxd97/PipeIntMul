`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pUfSutof/nrjyV+/s416XjiP2oBbRkFvZVtgORjfKB1C6x54Xkt1BGkWu4u/4W/m
4G57SroVyuatSvgRH6ZwHLRLkDhYyhTrKEl0eBtgbHI2rw41qos82l4+YHfrBRSN
TxxouUMdagh6Fz5/y9urt92w6Qr8kS52kmSlkA3r14RCzfBhKQv2GPrid+7eWLIf
uziYKnMb23jA/LKPCKimGQAlnX1evmQfkhXbqRv47+hUc95K2UIWuK2Nw2SOVXdC
OJQq+DN8IWUQFchl5SFsyp6L+g+dQoqqWmGt+LOInmW7MJRXY4GmwKGMfY/8esN2
DkP9I2oCBtUC7GE6AzyIB5viXatXRrAzLHYpw7DhL/DVIN/dptZVXMFq0r5bxtDd
AIXDM6SIjW2y40ai0CVI7UqcXTGS8Euqx52hDXxZYyuqXlybHYP6Vscf8kfP23RI
RRbizJCFVfyEBQxto4j7iUR2G7kRhWNH7bHoix/+lfTtVFTY5X2XZc4otLz78kT5
`protect END_PROTECTED
