`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rBfy6B1OWZPcMwDk8+9mwg5+gYPa3xv3Jzp4O+u8E6B2jARMetVezmFKecoUwaTx
STzTOt5TBD6fu16o8RwANIdHI4cQEjuh1DCUQinaJUho9MhOsHJBl91qA+OMB2oO
pBraH9SJhNiTJ9LMRrChTXoG4+5DUr/Qdka3LMBK5PAss0xPEzLTuQ169L7fCfdF
YC4Uv3NmHhmrNnW5SE0qBkTubx6AWKpsQOduWsFdOAkSFtBe+5O8S4iZmxxuEDlK
I+wSdmcgl6kn/DqOPcWdIw3xA/0MaIXef0QX0sr0f0eyARXUm2Ek6Z0sgquwdrWE
L31aYBnzpyYjdokxv5D9Hh021Xsk4gAuAv4oUXh74GBR05A79w0HIDNV8iLvJ+HI
cIRXwYQoBrl62LNAUVwj1AKadz3Wf2h7dHCC3jZ+5MkuvMyeja0elgDWj3B7/RE/
dUGIXvav5tz1PthjqK9n9hjc1s6ynHW/O7h9QKfxpyhNVzQDHLZ3fW+1niggxvex
lr4A2BpeznD+bDUx6pBhl8I/iIF8Ug7uqpX9aBo37waqemYLBJ4QsViCwOm7TooL
kt6Ja1CBR89wMEChNXZskT6nh/NzYsuahwyfZvH/jWCl05Az0mRd8xjOuiuSbpoY
owFDnQtF5bMVolcQDFrmO+Pql8PjDkMVhSxVuxYXWBPa7PiTHlwL+qPIg2tLV/WE
xJA9CRevrGSlwaTjUXAYarSnFWYk2yvDadTbDNcl12VBjyVqpxkQIa4KnKvtOsdU
+0fo0zTm6SdYWFRUXUQlX3bygXmgdQOGXGxD2lVkI7YCU6zTGntHrxuNC3yy2UGK
QR7FbzEtBMrTNosK1c+xUM4RYOoV5Euls+JtQJs6RpkqGwejZ/xZ3aWsRTIsOHgW
XWdFjVx0al5XwCAWmHH8RvkIavLBK8Wuf3+msBw3TnJpoUJ4tufFkSGx84zfV6yZ
eHeZpedI/x/pzia0pS4Ai2kxeA291ERNWXGfy+q7kBH0Miuswnxmzkv2wYxUiBDg
YKdQsDa1rAyTkM8QXxQkNOW04Sa59wz0G//+iwZTZHo1DUCD+YFhS29YZAcBohhB
IRTG4pZaD5Gi7FwHSwLpvM4u1TS/Qe8xDsEH3SxRqLYFka72iPHi7fLG9wkO+lxU
Matru6uj2J9zyu049nSOH1KNPi/CjvtDdCXK/4+di1dtJVyAUZmvZWOe8FWmM45q
bLlstvzo+YLal2VOy9BeWXA4kKCXAHOUN5A1jojf0/cqlBE1eC3PMNbMTBnPWPLo
U1zh29Gjo3bzD2QVgmbKb6ZlhKpEUgS/XOEoOcieB41ShjbVFH4a0Kwl+M8rDVTm
gQRru9dKTg3fxRcrey0yA05j7ty+H6C09NtFet8QogmWovdA1pKJnRAyvX1GhC98
tP7Th64GWX2WDVaHMDxXZU6YaRZ388xyuwX6oKxpdwo61KPzkzT6o1I2Tp2hmDAk
BnR5ZrZ6RhA86Jbzow12bK89be0ItiNLrafmlSFgFX6zA9taH3c8GMlgAqAUIe5g
O3zAOCaqQmOTiO0gyR2h3aMIF+M2mxKwKVfRuBzA7sPxeOf9YbTWZAT0HdoOMeKr
kQ3Cqvr2UQ8U6z2ASRUrlx3E0sjyKFfwpr5Ha/s4wM2YeLGvgtoTcKl4Z7m6tB0k
4+OP4lmWVUUQlfDyl0PBs1oNESkt5MdLDhCTB0ihot2mD08DzMMVJd6PTtqsdqVp
wr+KcEmRBfp2Qw5O6ezi81tj02yyOEi3oWP/dElqdqUBfmhnXi9mKF69Mrw8Z/CT
nQxTmHwwZwOJF/mBzKBfo9HJEXQQTmMFgfsWx3RzO1MNe3qus6EMrfWuZmneGtJA
PKD16sVkmKzJJiVUefCbE8A6KN66WqfOlhu9BipraiCaESN3YQfB2+YHqOS7T5Ed
JpS7C1Ovu+Z0iN+tNyM2aqdyRZxiR9a5dK6hJs6QMUdvQshbbyc7UkJ0/j7MqVuE
5OmWchUADEMxKi5x/gE0Kv56sd1f6tYQTHpJUvy2pkVx7Efs7y+KZ5+vwU0+1FP4
9R4BFvCQUrU5UEYwyklKaN1b4l9/n44UZ6F04g2o15x1VPe158XeC8t375i10D52
HbF+mlKnZYt5gO3KdNfptvt1GXuaaYEn1QFkK1M988Fqwhk8XxNOGflScCnXV60B
WjRQP8jtvgVuJobw15tc4bEP6IY3eEWLw8j4986v37VsbKn5z+j0XYBkFahWdoQ3
2O+KLT/Jx6r1khE30CZAfy6JGHnf+dg4OH4iY1OvjNESFCgPKj5R0obwAba1wqyH
+fOSuaEJvHPmYDxIgU6foKaNpyoElpWkrx31QoYVV7cCP93dlz9J2JADTxRNKaFP
cJlh+PNVSnAusK1u+UInfYMobWZDgT2Dsm5B0UiSTz381Su05t7EGbU3fo7V+/gl
zobUtfKB5AgwbZbpA5RLbIr9vgphiawzjHpDyDrnLOr+2STIPpKZWw4Sd+F/zQBi
tz6XBpE0bqriOqb2Qg+7DDOlnSC0zrSXiMa9Xt2A5RMAHpTb+jSwgymjTy3dRy1E
+P/VhYKPnUwEYwqCw/eMlgxN+10XjoRu7CUSsDWZpxdX4haXrdyBdmS9YG16HLwW
1SMDLygw6COsbXgS1yJiEPrjfgfR2Uu2KndVAb7PF+9BDKv5vdpeYrHR30W3nz2w
AxFIV9xAuCNBFmAkw1uC34pgkFSE90xLS0UndGxRnQiotMXcW99V/mZGlETnJep2
Isl0v8R4hve10jo8M+mr2ByK0smAK+bjKS+vEGrSVcjhKO6YUAMOdMmjTbrWXxub
16bE9eY98QXEtQXOJfiwptftMJKfqc3+EBvQtmRdx3u9KVYcxdJy7rGBCnNY0/wu
aHMDvjddguyAXYoh9pVPamDhNuYplLLmmwVWar9biMU7UWKhsuWmqsJ+lwu37BDV
bCbuqt2Ko5fy4OPufr400L8fhG3mxr9avryJJNwkemscQzzxLBHu3SS53CbcUHk6
WrPXX4/Q5oSWE33HvC3B6bDZY+p5kjJijjoJ0TZ3zG6MzW0To7qI8sdw+SMGGy/x
dNstB75aMFcsPxJc+wZn2tb1sUwKK206USUsths+3QcNIIwXPNc72/s/0u78qcxJ
vhMetvDuM/plp5N8rl/ONGaseD6sMsNNlmtpMIvihUCkmyN5P/DvjHh9WKOSkJah
iqi1Cslesu+zSeQoDSRpxBNkb872PYYmRDk+17ofUDS7KchwC7dM1iPhWlDZOE5T
PZJc6/2lQiny9s+SZK6IiiHKkyF9DxqDMyBMKceCnasf3cniArhwFFwiT0vcBCAr
oVr+InZOkA/YNmrA59Fddhdzl50wtC5l9YTl4BF/NZEceaflnQ1HCHBD0L+0BoL9
3vYHBuHAW4Q8ne4Qu64Cv6q3MHhED7qWnFPLcC4bmuZYiOK9YKyhwe1XUXqndX25
2ZCkwPPqtHkyoXlV1V3Mi7nxWiDdTxanHXZzvNFCqaT1fhEo9vXwJyCeftOg0GXj
dZbJAh3Cc7mTfVsx4jdhMII62DMzvEkBD4iYoou7mdOmDNm90j4FcmZS9gTUnJls
NV5ewfLMiGJn8dbuKONhvH6NT0cz8U4dU4+QptGoFFgZa8ynk8G1Xbv842oiEKAJ
mEVFBAQv0cVBOSGOZdUg+DT/PG87HRLwn271q87mJEptVW6HP6q5Fc8NBxUOYL3Q
dqPB8ORt72m/DV8rjfYuPD+REPhdi3b9k6FivAilUJmw8fryfevkVc7BiMBimmLF
IzlSiFRw0Lb0bHRGJTp4VsAru9Ty9aXZBaYaTY+DThgGUzNuzcmTT4zrh3+EZ+HP
cF2HXpY7R2cHs9QdZ9xqUcDlpK7LGnINOij36TNybhD3YGX3DBxmDiDI428L0gQM
SNYhlRr5sxg0aia0NUYKzYRszazajdrMvgFbUvnCEExQCDbBNhmWy9eUxCHX7RGj
PUZ2d4JrwmXr993CV2bPUKGZ2j0+408wvZG3Pe8ZkcJGHZYSZywwGZ043a3Ib53G
ZUqywUirIU4xAqCWx7d048JM7cfinQA8kbIubAWZhLUcp4JJtuzY955dQTtySwXo
PN3/3eAhBkQXbA+aYzyV8KCiMt6HoirdrRwEuKSbhHlaVpMrV0xc3yKU8LtTy9wY
UK+kqY4RY3Vk0zPpmkWs/jg/ISxxz1wMLkWi19Tq65D4uUUrmjc37JOlMe/2VmAv
NX8tL5uBr6qdywDZu2jK0hjYgFjt0l1mkDhnqJv4dR0qxCloIlYbb1Y/xoKfkToD
0l8+hsnjhO4UR86u00F9oWAgDBsFVOllyuRHHXQzbkcVMacknZe6mIjMocYoqRbd
eSU4HeZDu5l7nxQ0vCNtCGY5iPNnxf1G3oAg67Z9lFOcgsii0RgJMPZmCod4nJJm
qkiGsMgShzylY2u395brfEwtYE2o8p+oiLj3BXOPjjvppwch2dAYg/6PBlSkhWeJ
WUysAietZ9OU9pf91VHUdt5RBVAqs/PERlwJPpl1EtxhCMXOP3WlR1EgKMrIwRcq
ib15ILOJArxKGDCRdxrJMbshf0gN6uvBdhcpzC2t6/XauK5dsPX3658zyHcw4Cfv
SZpUUFIeatkDbpifeV8lm4lFlXb9k5T5BhvnT/QTRWilj1ZoxOlQ7bKoCl23GbeK
bjfgTXVAulxVFDvPFm0ASOApjOGOrFjemugYluZGDpP0I7SzlzZRNczPV7eke93Q
O7C6mA23674YAzIBxa3yWVhiwU3698JRGzOJJu24lEXIWJIBLU5PkrIkhZ8DY5WC
hcb0c6ELHcNyx9eSwYA0lpSCVBaXceOdlCe/yBGXFkb1djqPAbYGR7O9lUEKIGRY
bmcTlKFRAh4v5GyGNZEM7FsZwTEawg91ucyWqEKDqO9lEm20UUDol9tGXFLlcFCC
8du47MtygCRXPxwyMBp5qglGUX8KB46eu678FyiVuFpfeThX1wvMu0s8tlxAjm0/
Q2FenwbMUR1wMj7vWlMzcJ6C4zVT6Yk5Br4xKTumVGX2UVfgiFh0xYfy0HlqXu/J
fpWPiRM+7qy96IvnAqlYr9Hhe/L1N2NnEzuixg7XoBgowkcw1xbt6xGvZ2mEazM1
54+vUIoqo8nOvXMwVjlY8cL4RvkdLncBL69kyMggHh9LPT8n9UrJaT9flX7V9Q4d
p66fF0R/3IKOGxhf1y8QC7ulpXPKL+meEOQvYFGqtcFPhH4Mf7/Opx4JaxESuBY3
WQMHJ/iOu89ZQ3VxPEUKeCCehcLlDI/GSFMVeYbKH8rcNPv6H8uIMAA14hJQGupz
xcebX2u+gznCyUnSJ8bdXBLh3YJBjnTWL3zDEkhn2a64nZ82LvUwApL796IPwxyI
javaqvFhfAQ0CrcHSb3tWARnj90yHWOlwIqoCKCxj7o3/3GlkPuNDl4gK363853t
lP3DY9O98CR+HqZ9dz5h0g6Sj/OPmSRGzAOLUCA0RZVnkmC2q4SkWlVWtYw5wUBg
j3nue/MNd4Z1iC7A9dho09wRx2E0qHGoTMBXon6kosru0oDJ2n63uATdd8UF6kbX
lfrTplSldo8o25182qLpZrDLqrYxvL/FS3xCND3uhT+HVM8YKTfTdmh9dMeUnYeN
lmT1nv8UrHShzBbfXiGfU2T3W8aOS3yYMXkxAYfiAIG0YPSAZnW3x2uDfCLymB/l
js56IKLuMkOw9W1pImAtIltogzzzRQisrCFX0SOivSrOxmrQZmZOgfVFxYvlZuo8
LxDD1vViflfMQeuAeBy67U4m6NQHs+bWv5iuv9qBj9OpNxBFqq+aGC0rbPSey9jy
z7lLbGzhYi/YeIrYTn/Wtd2IC4K3L4Fk4a88A8AIH+8Z/gaaiaqsGscX72KngLYG
ffe0QvskrXL/gG9azdEilNckjNh2G/8tkFtcN+dV6KU/IDq5kVa39/UPpwNnXo7v
mvF64Fe5UwHdu5L9zrQ/deroKzSjY9W+77eC+qXUBxoe6LIvWyguKdMH5+nxCF8k
lUDrKcfpJHxMJK5t8FRT6E+zUS/q0z5/uE2l2L/mBn+TnAmXvI1t96oypwa5pnBL
zEn+EPzs3IaAhaz4/34wu50A7j7LfzT0usyMJM5H8ECLefBMoyXeRr6KjetdL2Zl
ExEm8PVqcrhTw1TN6j5ylN7DT9hRyaEh2YlpRyZwzgFH2RYlaRH8xcT7Nrcw0sue
pqn7zeAs/4g05rAG/rAmuhwtkRTdB9Sq3nDtNdQ5IG1bJ+0jpev2YKHh6Vci4Y02
1nhyfRmq0Siggw4+BbJb0MH+hno/4IiVgxvjFZG7f5W474DYidEYvB/fm8zFhz89
3YweBgoXgvqBRtlevR23TTEWlwfDovtD8KQjSxq94s5EOzdaGwfBhOtLVCGaXOD7
iTNcIWsAaaMTcOTsyEJEHehFp23J43IrTovXYIrC+y7BmBwIY6KE5970gbVp+oCe
48hgRf+VVv6xaZCc3/2fZM4bn7sB0DOZXkFf8cu7iXgLnMVf7FbOehnf1dMcHScH
ggmnOd6FQmT51n0XPAMtLvmI9zSaPSEanUpFKRrxLlMBO61qZhF0V8zoauie5Isj
yUuPFbNpX/xtoFVCVbg++iUs9MJrlNKtLI8/GgFdkm9TBUGRz0Fh7lAHgb7LN/8w
vF919sqIJbdp/Ff2pCp2dYPChu/ZxJrxAGy3qOx2rXOQeOXlDuM8nrQ5vO8zdn2l
eiu8iTtj7aDouiAVPgIkA+pokh6KWdMmf4Ey+g7BzQ3yVyH2AQ+XkKem7FFHeze4
TGWJWoNBF+1m8eXef2v/hVXQulg+hEe6fh/ZJ+0e63HurMtMXB5iWxUPf7Nr9e9W
3HLsO1QHCBtfDmlrJdytwA1hxLywmy3nYeU9ndhZUQa/vcUxm2CqgIORr51tCKGJ
C5kVaA/evXA8BdL5Bl/0rnLEle6zBKeqycu0c0fN6pqOpSvA64X9rWFefsUqBWcB
79phhBXfGRm+7WXZeCjx++MVgIfkCKUzL0TAfy4hrP2Td5oxc5PxtKNccoNrjd2F
xFyOVQrGBaVQW87JfYqDsuUbHQrXn/TqFx/HeDDV91MQPCLF+p3ruX7Cl4h6M3Gj
7QjT6gQBVhmuCI78+kNUZhPwtG7iJZV3pYLg0XQNBniYXgHj4gXZUoZ84/wx0/7h
uiu/YBYb/E6jd3SaVlXUPAp+r8yn+peDoxNieytBl3BDPpf+EsSjM7Ykm8fW7ogu
AiIkZSWq6V4jWcA1DMzC17eRUnDb4gJRW40ZctgJyGNLkFOgPUKVYhdhmgbYUgWQ
hpew/FmmZY8u12sYb5Yxvp4FPoqrGV8iMuNMeX70Lb28RUcWGIwWzDlQaA6T7GA+
Ky100HgtKC6NZqaAmiKoCi3wogmjBZTsg6QhhKluCgJReGHrvw0UTSMPBaQIEH76
/mXYYReEyF5aslJ9bhym5UlY+qozzGhrCy9rWitH2BHl7dPmt79qY1JTnqySv146
Odi24ceUfW880W9YRdV3r6Vpxk4uZLYaV90xHDVp0qM2JT/KNlCq262bBdOaerk4
fc4dWDRtCAmdvSwHqYB1LNkIs5ZomjFHImtNTvAkJ8jPI6/CidlKBg1kLXTXtEMw
ZH8N8uRXGH0Tdo+ETO94SAPY5sUb0emunoIma29CPkfheKkg+7a5yXliiwYWccj3
AQywgbE9G4ZsCwAVCHZACm0AivI+sq1Mllo9AS2PH5c9EgHKWxyVQEfhzOqxC+Aq
wT9fNgY7PXMkjlAUI9tx1IhjcKc0X23FVxzuRhdeAOcR/Ij3GWAsFAz2+Qb/XqvS
FzXnKX2OL4d0lsnLkwzb//Pnj0JkMw/C927ikRGS1sKoTCdr9EWtpiiEF9Rlt+kp
ueB3kIxUVSx799hxfderWF47cfsfdzmAEx/pl5Z1XQn68c2B7CmTiqqZDbXli+w0
fR2D0qHEnbauAHNNMLb6gU/N9xAf+INi89ixYFuacY3PftsqDuo1fWEc/PjfmdsH
S1mhPSTLfHi909ASQaR1M1YbLV+sYVvG3ocRNwUtnKIqE94KP3vUap5s1QyzKNur
bpQf4UuYCMnb0qvbL0ZK2JlpVgAYuy8cdZdmH8fJE0CKcbl1xCa7RzwoQtMAM8lg
+z9+YH8gCIw92TlwZgmgqUc81JYimuQ7EoVC00gh7PCE6fpAuzPEwpywwgHlLbYh
SLva6RpFMVAqddQDLrW1Y3m6SXkiU+8HMj6JCTQ3PsozjOMqoVwTwpVu7jwypXe7
KJBY483DeoSer8pGSuhDBA8OGKOCsKK/SL6nYqh6jY7j4gSQUWwI+9EoszFr77th
31pgniR4Ad5d2XhOeinULSx26CgO5daYmrK5zusmM8RL/hF0zZ+AB2/3DmXTTjp5
r5Tmxh+r6TZmEZx86ZhbQjzbAvPx/GWD0ebctYCDVKu0NJGkplexFxBjuCB/usIu
jgIcwdGYu6b/OkUTsISZC6EhhF2AJIkmWycp8lg0HO7tzTDOo8vL5GAosvnB9cJO
Ief2kJwDlKzWCHCpFIgY4kXoNwe0d6ef5T3oZokYBPm0UJbvx77s9cVpyQsvj218
r4/yw99/8zjd6HcC1tfUuL5Z3hSiy/Es4W+PKXZGB5aZcnDrD0XF1drFi+9TGlwz
eeVr+xg16DRiO/kFgaqXvAS9MAY0RVh1d/KS5NnrR7gDqb2STD6qu/za58iw2y0a
VAWZAkRvdz65p9N7v3Bb3BN32BVUISSrmxq5/ugmd5QJc7rk3/P/I1MQfSTzFZpp
rFx3W+fLdyVhtELfyTKCCTfLBhZB81GIminw1mQ0uiRLJHedwL5upFsabYWvX4Yx
DSMO3pAj04q138Ho00zf2VlB8Bd+VdDzseb/6OfcjZ6rk2v0DSBsNrJmvzzNVpk7
PF2s5UtUR7FAnk8tB9o55PFQr7FCPGcOJUDEgK0uFHW09fQuPj7rsOKZaHDGqzVX
o6ZJJR6QvI8YUHLQ7m0YOPClLPqEvMXwKmgCJhE8Rnz+6yB6k47+hM6liMzPbEc3
WiaCuY2tLiT0dgD3iqHBAzhtvxFfOvd/ju35VMYLkAlmFsObWmwyamfVJQ+P6oiU
UsKNRbyq+9m/hLmAd6ChELTUHz2aNrTQkNhBQURdga7QqJSn0crxiYVuF0r48BNC
D3zZ8ZRHLzqIdJkCk7xT9HGFe+zmUSZ5L/tnM7cQAKuLk/oNkkiCobfnWE9Zgnxe
tR6buCN+4vzPUaKsZmkWBORL5QEgZXza5b5sB8THjW5v8GV5y+aWbz8WKk0OR0xa
l0qNVak7waM5lPbhVVFcl/1muCtS9OGMd8KWn7d+c+UdIJbXGzyOZzHK80DhB5Ma
E1rOegBbb3uKVClp9vbeCxGhwg53qPLhB05ehqQq8NobUfC/FCXpxnvdgb5FiURp
GNAxTpKDKQun5Q7Ou7zFSi3r/ty6VCbXQoSgGqOOTw+ptcOklRqgIX31PbVP7vYl
lRIYaksoRG55hSrjDUQY6TEHnst9DmxoZ1hh05G4/OVzd7bc9VaSZOJkdNEoQwO9
qoS/zTjlP2DupSp/OWlpv2K0nx1ldj2yArW4d2Kb/gDbeFuXqtYY307KomK7zCWO
djLx0K0/42PQ0VY0KIRA7ytz325I5qmwJDzKBBr+OnaWIPJiH37JLADANAMr8mT3
DcrahOnyXLHjWMpT/lvRyJyg7LxdWBeHncANY3SvTX/fxNbtS2ZsHOrAbbfMyH+M
KYATEwSc1tFlCb7IOfNj1g48FhdaajtoHhMlkhcAmgn7hGSj+UCSzP608BiM6unn
AF3SmcuFJxQlQ7iS7H55Xdx0xpWrsf/3vb0THJK4tMzlVgtUQgKnTuPrBaD2Y2vg
pLrqEsq5Sy0RZhMNI3eFvIb0WO94uHjrdzhS3eQEzzsnYMGIZgLx97JJUrE3uxFZ
tkUcwlQCTdlxvIrKsdwDml6R6ou0XzvNUVS8gxXMkgQnDAxcC4ejEjU15v8cBWRa
xqX2ImjaD+T2WVBYNYiaSheAW/KCgU4irvqzSPAyAv2z7L/Tl1a53vffwbYftIiv
07H7LpJaZEzquRGffiK4SOwwYno/UAPRuC+SCLeLHTs5283P7lUYiQp9ZVpT8lil
r6Bznj5H4dQ7+8gsOnEGB8nmTw9GxCmRM7hWOodWJyvOWAS3GthXLeqApjtbVtNX
yI3jbVGQJQxFy/rdiyOxgdpuj0lvshzxb5Ui4kcouWdwZI5uLzwT7PmComLsRZOe
yW/bjMmoFU6H0b5dVD190zc8v0HEtwtUisY7M+u7ZgYunbKrHwVERrwyvY67DvCq
QwymUfVq9xFC943nLjCsOuHLOpVNIRm8RyyS1v1VJGi/EaN5h3gzVaP3dtdwroUm
pjquPAY3AVr1uXsvwhilNHJY9fEdYBkcZFARKdNzJOlJFvl/osVesgeLZwTDtpal
WDEYtnjyogGpu/BOCOSMNj7AjuQsO4xmGd+w4mgExZPa+3irriEfI+xavY1elvSK
wGvwYbcHhhCI0NruKE03xQneunwTsnZdH+kp/w2XWahHYzANA1kBdTzifmS3DjyH
QsBDNM5pdg7W76Xxemcd8RsM3lkw0Tl1CiI7cIE4DmkhkjUd/neeGCHBbhNR9OPM
TDGVGBwQE2MANQSAXeyNCQafMVSSiDhukGRzOZU8DZ1r3xBE8M+820GGvLK/R+a/
aNSJlF9ug2Vrta32F7VlVgwXEpPeimFFYUM6aYgTeLL/scPuuDfCqX3sFY4HwNJg
4QDI7fBJJP2tc7+ZdSjyCp7WY4L4goUoLDqXjkTZ5Nb7L3jFKoEBvZSVk4jMaZDq
VuqBtiPy7u00rKR0nyFIpzFUiRzsRbakMahB5m3LQX10ZLE3ayI9OwlQyTpHljP2
ve2jvLRFi+wpP3DNdfank6t7EwXSFihQaIFksiKXmt/+9BPBvd3GIP1vtwrsdh+k
`protect END_PROTECTED
