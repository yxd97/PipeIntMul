`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58fCse5E33DK7uPZBUbllmRUceHwp98RoCHHxEUWjHu8YTKsb/iLoKppfz4xM+OI
WVypHs/oR4+qTLtNYqhBdRFEgFv7xs6bQ9XUrXUGFKPGvE98WsghhYzQC2a3DddO
GM8Al09gdbWhnahrAzWy3fVydcfkgsobYgRc7bdCE0vysBJ2rCl6pq+U5c4v/CWF
KAJxztDmlrWTIZovM7cuwAu8DmDv1Sbu+R+rLlGHvD1ojqOJihVfrNiab4Sv8wKb
xfxLZ7rzPlHCYsoDdWbPAXUt695jbRC79VsdxQFuxaVKAoOKHWYAeNppDyrJQO/F
cntD8xOUqwejUd4iQSmfrvbw1D7H1jJyd2rmJIRpUaQ4NgIFiMJHwPYAKNrfaLkG
ZffTn6ghTSYC6g7ecB84GADg2J6pxlVuqsMH/sIF22YPXxfYYs3M7w5rheJXPu6K
z3mJIz60c/PKqk/LAyhH1XWVFHplDxAvwJkyY0C1kwOHr1I8qNIEP2rWaawlc9//
xyHMDkSXotIUChaWVCrR0RUDWGCxI0syXQ2LpPpLrQcLVwrSTdykOGhOwgo5N5Ts
Og4CB4gua+er28S1mnfRD44hHDlHAf1KY0YC96CGQKpQ5le3mipjMo7M2NHyxREA
s9GEvx6C2k4mahYOYgocoybBhJx5jVVpaaURogg/4zNp/BtIIMHFD+q8YZ18zMCR
lS8P7zA3hNwlw7qAB22bkvho65kx2+kkVSxjZvAxkQJU0xq4GyVi2o7CbZx9IGTf
`protect END_PROTECTED
