`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dwdcdQPIf9g5oG7BRHTABxxer6mmdhZ7nk3we/iikk282RIsfkWss+4DMK0j4cwT
4wWIFS8r2TICGM4o4nJAHKQp0/9IkuVCFQjRZHybAsD0XbT4jSyySaTPnqs2SfCR
jboskDKga3PqHmvHslsh6PxKIuEdMdAI+A94pjitz09PZhANu7wnhc2amS3APjhY
ie1CVqEdLYju5o1TjZO37OgHJTynUoNyHYVAsJs/UI/pZXn8OPfhqrGLLLPEuEEt
zZhwVSleOv2UgZ5wDMduJ/vTA079Cs5ekaA+7LNXkBVTYtU9R6zk1moCdd8T9Bw/
pYplkZ9QyAg02sDSR4CcY0fu8p+DQTL9X2ciAcde0iETzJRYbPkrHe+wBkW2yyqu
oH4OJEWO4QZ6yRxb3CWS4VIFUPj89jMotRuCdmYvwwlA00I8um0tixg8gTJBdkKs
bE9KdM8NjFitJQRRY7EFazvZzR/9KoqQphTaLtdo3uRwdOktkKx+QjGwIbZzztsQ
6SYpgDPrQrCwVlJXLFjV/A==
`protect END_PROTECTED
