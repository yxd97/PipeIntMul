`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6XBppaifcikJT8M8+NtozBpMFz2swVFkHJn2xyvUyIgIgu4BIQg+p1JP610o/nt8
ZIsqrjJcPZxL2G0e43eimrHbWrDBu3w8mlUEOohSqHr/SU0Z6PSvefEpSz8MCtmk
KJtakhGHNdr07AKJKkvZMe+9TuzMvlHxD8ah+26gjuOwWF+uhhYDT0rOlFzOcNtG
hqsbeixMCYbhw+sA8S3+lccpC3oEDR2nN+wDfhGIf8Uxsf+YuTXobWIUK9KSsfOM
Yy43a6LlwW/10kUqJj31b83hwm5uT8ZhjOpds12qXvsFqAuCZcAQ3XZ5xWFkKJQe
6ACxn0uZzy7MiTMiF+YaWOlPNkMm3LKDtGmPvY4uML7Mwz9qmluIl/YQ1vJ2VEdQ
WJBpT/rkbkH0zUowqCRk20AxPJQf2q7gItel60WXUe0=
`protect END_PROTECTED
