`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYN88DkRe3YobsaDLh/5Wa8nHpsTuzB+B1LxFzYHfCGbbCre42cDxPkMKJvOIOHd
cGRhZKYEXoH50av+GQ01fjjd0T6Wz63ZI+mDc4Mp9M9t0Xb6vCJfWokyauZFIgQz
OvtPxBlR7hryXDffef+aTjlIkRIwOofBDZMC9W+zAbDMEdsbqmnLLEszE0hFbpeS
29S96hjSVhVO1NdUeHH8vKQ07NEC+l4DjBuSU1TOVnzp8/LbX+dO+cso85zOHL9i
OJiGGbv4PDQe8zAO+OF7010OqxeO77R+UhIhN5vti+tbFtrPgoXB1S8gC7ICCq1/
TVSwHyY5c4F76WQGxZZ+sFb4RmWxKJqVAqVW7wRysCJVOs6uLs9HYcH/vtl8I5QV
rO4XR3taVZfZUf0G7q5R69Xo9zUOEMGG5T4SCrjOMfIpfahvSitrIy7q1hkDgIND
eUXt1iTqyv/1+0zvIeA8dTKDjWLczjaRgLNU42vP7mQcRduBjYJBgUE0K/bALpZm
GHxZoLM2MBVgetHmTtiSCXYDFKLkovrSTbWJ0+q3WAWc8tF15E53th682lwN3kfd
CHtVVGQfe7TRV4klDDs1cYzKzWQQPwnNUpXuEnfD16GeoOl/j4YR8ggJj5D9Eoj9
FRwQ13XHN5tzEO1UviyVZZKUvCyhUDwJg3xez09uTy4F3sdU9nGKwtkFFlMkkJt/
9yzblnWFZ1yXIkHl/KaKbc32v6hcpD2daGtW36wBtVOEYwUT7uwMsuFk1LNTzIf7
Ki8v3wbg8JXoBKFUQtIGHEjxhqAjvx3A9f6PqJPZCRX050tw6wJp+66O1TPfmHe5
6tZkpqf0Q2ezWs4Noeg7HGWxVgSSi/a9vxHOJwCNOG3gScIbu402PIdgOF1k+BxU
PbnT8+NLd3xZ5U61X7edSdzHU+a2OVknP9jXyNtmBT1berFGtBZ+XgzkJMqP5+bA
w2AVySJF4nyjvnvRLGr2kZbT7+iQm6zc9e9b7q+gwUqNdC4KQ5YsWvRUe42xHoKx
5vX7CfPjtLmovTC61W5YkzonwBw3ch/Qyz5IDZmfZcNFO1GhS2acMUiw4D70N5jX
h/UpXpZKHRsro2cl7zmBxf2PSxEsOfWqPEwas2ruVtRsxDq/WLNXWGyeKYvJD40l
x07Wwmkjx4N4pMPoPjJenTIA5MGnB3TbUMdpSAgPo9UIxGQhzgnOeijMiM2J8g8L
pV0ZHZHjsUi/rnb607QpsNRUPARqG0X1qfgJ+PMKaUYfqZvXXSA2RIWuGft3aTwH
LD3RekRDZwNcNtpu8hcEuo5+onGz8DkifR2nzySgb4bx2E6zoNhwgqQOjJIZJcTl
zuW92ffDhTU4oY0mxfdw3+TXMFO2ygvSvUplaCf6PKIgYARMKNt/8i2+I+EYwR0u
2Vn9o5axqQiY5Bi1SvqXUh/PM7sp9ZRBiRJX75ETt9U7pykEKF4/ChnkPLDn5vhA
/rVepgpJ102ZXkMpbnUEe5Gq8x/5byGF2/uVpErwNnj21Z8xq9pVipQnG2L0bBu7
61Wbvr0T1nVY8STvZvsWCHXyCQYbxKgpTW49/7xDS4I+2anoSYdtlywrjSVoSduP
J/CFxFj4V3BaPmeuPN3HaxXu045zM2PtCFMIgTVgVTI2ikWlQSs0M9zOOLQr5RGT
HiylTSC/KXmZ7n6KujyOcNZR83eBTggLACdyzvj/K/0hnX1bEpAreUZ7Z/Hly/RQ
qO6g0z/wL969qIzPxrtoDl4q8pUecifkMDF7JIVd2giKIDJbvq9iaGEE36acJRt5
JP84js6id8mdXfDbG1uChA8+aX6dVXM70vfmWNYDFPYVagXHSoiVXNBNcvX7Bxj2
rJUBlyQ29kkh3S9Q69Lr+ifM17cBdnq3gXHCTiTLVKnLoRcfO2Bra2F+3kyE9eWF
`protect END_PROTECTED
