`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7/8rCbRpWREIKsBrrqQcJEUo9uavpwxbzKk6dm/vCc1Y6OOXaoHQaoxFWUYwKiE1
tI59BHpHZePAm/JO9UjJ/PHngbfS67PcEi89k8Q/9I9Kw8rDrWm63HZU1e+DzoWw
wFLUFHnsSEg+wvGGRVsTH9ijacK+UsbjWDEoUO/owuDOMR5aRths2OIbIhKFq6Lt
+i7O/cc2zL2eE8dYXYoy7jnnfy+wm1P27S+2kf9HuSqicNek+rBjn1Erxc+kq8Dx
fKYfvwOhpL9TiRNVppYEph3kcknGASVyH2AK3HW2iIOujcGyXafQNcS9m9YsOWaE
t849hisba70G0F5eT9Pm+vrUL8kLTWVLUHKlV5fQlOAccrO0CyzcdUvv0tQ+43Hz
/EQjc1OKYpEsx2WFnSO1ZmUKo8PxWKRIoKW9arsz+om1GNCTi+CplsMHT6AuDYNN
P/sS8UwzGRmDNh6aprhOw4pPJtg/pHoazzEXSAhSZeGpvhk03XJFg+233wW3YLml
T9V6DHNCh2D2uud4kDOq5H5FVEqyVTxlurPOhBrO0hB7QOabZGkd2z+FEC3Y5AAc
lsgxbq5ER7KIil3kbzNb73BZvuQwMY75H6PoVVJ7Z+foeMh2WUnKA5xin9bDy3l6
XtUsk33kBoP5LvsrrnSK2A==
`protect END_PROTECTED
