`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sR4xLMt1kUpF2YIxT5OIj90VrM/3kV2ErF53Kuh7fI6AplET3Nib0uJBuaHAupTr
hD8cB3pATR3aNXtcImfVUGlfcHyirx2//0SXd2kTv0nv47xlMz7w3ibYJxqBTTU0
jBRybZt6eByzVNJq/2DkexN3/wkDW5LDO57FtjTSB5N3VKgDgQeP/0Ue79dcI1NF
bboFcDS2eRURVYoR0/4f5nm2/+FauL7RkZftau3BVlFKJDg3p0EyAuHl7NuGvZJi
zyYx58xYfQCT3ICvFH9t52hlcgIAW+EULWejlOuckUhHA/BAR7Ir3QvuecX5xRwc
/4Z8Vimej6cnwscqpLHbclj1BVJZS8ltNCZrYaKBDNO78Oo4mU1YE8HGqYTg+jve
7ngOocREG+BfnZBHQKyQ8Q1nbZEGGQ/OhSiwRdzFjkJF41Yi1J29dpLyGUAfdKVe
DfVw8+xQozZHtPwLkny5oHz2ACqNe5qLyNV0ywNT9Cdt+FN8kcXTuBcXOcPnd9xa
Ug6bCwTA4Y1Kc7JdNzGpfMSIs7KfPtvGTYZBncKJvOH74NNbRMJKEaBYtWYohXNs
Fm3pYJS7Bf4C70iCcaXO3z8FxzEf8uBn/evnyLyksBRA+jodGRmi0Nq5UbfGAEP9
xzvzIyjva+dHUlR4mjiBdkrJmZSrNOGWO10Vg5ENNUL+1LKJUBiteBkai4buF93a
ngn5J5Iv6kdHRBUwKJ8ORQ==
`protect END_PROTECTED
