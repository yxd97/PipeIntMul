`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EMKno283tCibEOp4tcKFO9vNpOSb8ag14zl+Avyhds5aep0xlLjNwPY6QpvagOm
f7WSy1plxUxhjtZgIWqHxXQzcTIX9Lz3IXz0bdX6rLqHfiyJeEeXVqIM1bdFrr8O
RLkfkxU9kD2CVBv9BVvtNNf3gd9Kgu2/FoEHm+chhPNPPcbg++j4aDx4bXoU4zel
Ko+AJkyTTz9Pnc3tbgOtq08TZ3OOXpiR/4MiQIYLSoeNexrcGxti9Urh86hvDHt4
JZNOzqA4jZ47CMX8cd0zR902Iw0r/e67rUvhklM54jtqO8Hn+ZzqDPZCiEh4aUu/
J1eKn+9Zdl8S/8Ezh+2sIQGFhZI397YKD0oGutBZx1Y=
`protect END_PROTECTED
