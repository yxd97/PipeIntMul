`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8M5Qo0XySWPymTb6gUpZg3jEyA/TiZpO9WDb/sy+x/++mt2Ms0cYcHgCdbVYoWw
ukkT4h7f9UFoSHsRciiHVRzO3Hl+RtoZX+MPXwQpcaIjV3Wz2A1d1NdPI0hVrhEj
mB7NnfbvPkRQR/X91JPsyG9Oc+8CswgQCrYg1lnSb2nCMjRWHCBXrLFbIEntneOV
dHdi1dF2u63xURJNVtPjXdCfetfE9ExvwoTUWxk4G/CCkYUM1mi6oqS+5PHNgT1t
tQp2/zN0jtySSYUA7H8echnkDKKTjNRapZHuKM37DbGF+qr5p+OuEnazJCI5aOtN
8Jsov8FRoGoEbr1eLOeXNfQW1uU2tT58+JtbDhVU7dXYw8+8KH565/m7aMyYXlle
cjIZXrVC5j7A2rTUdNrcjK50fcGQXLfLmcbJL58y1Lgj+DrYSAQ/OlprV9wsHYnp
rshPC5NPnQoz/f8FsGd1GpRYULeGozo8ZZDKD48lq9tOPJG0BA6FzcGPVOKsPdh/
owEQiRnq5Vk6pD22Xol/zOmhicu/Eg7EXE/UARkIc71vt4z/CBI7mkiNnVGsD4tx
f4Pr3qE2krZP/YFF8Z/VxSL2/7v7oF8qs6oiD2AfuRE=
`protect END_PROTECTED
