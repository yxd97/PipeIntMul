`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5nwSHe68O7WhcpmzY9lrmPgFt/Hj/H207YRPJ5gQUyA8ijtUgW14HLObj2gITEiu
L/pkXfqHMRwrpA+8rzokKieZCQk7x0jdraxaOSA269EbERzcUDkqMUJrSHbtKdPk
5+Kv+nzRi/iAyr8UP2sGom75+mUxu1D+UzyWN5zOyX3jWbyydENfIDTR1HJ45LDT
rtwE42o75DtiOlcK39qzhqKPQ75iKolVinlAK5uHP4npQkvcv4rU0d5/zOVOw7+F
B68JCN8XHw8J8MEHKhCqCNkTfh9mwixC8lL4JvyKsbfKimQOA6Xd5Kkh1QfMp7cc
IwQPxMzEXPb1kDtftaCzRkG1fCLDatolcmJ2Q9osw2WifT5UHDH6K84KszDBsjrV
2uAhBofcGLqR58Ts/YIHyujhzrkjTBbYfz4QsbPzvNs=
`protect END_PROTECTED
