`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LWStTJ9y1O/aAQ8NbpLmXVNre6NcBrczvOUyHMx7EMzbmSyYgA1DsNUossbB0rX5
yjetjGMEXJTOZDWQ4g3j1yC3ZrUxiLjvzpdfOKGsQo2J2ZskMTEw3pz2wrG+YqtN
V6hLDC9nYtD9uxWY+kVpsLQojd09GMe3R2wkear8sENRcL9/XWAdNDsJl/ZmPWcv
Fgx5ZAeESKXmnfkgW/QhT32ZLZBRoH7kfPMfK+1fjClqIiLJxRcEHJHxdtSqhJTm
AGCCp+fe7WkA4K8NdVADjQO+KVS+aP+XORdmGxWfgUU=
`protect END_PROTECTED
