`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xXMnbY0eyrINaXVd2r89PvGmzFI8arPIfkHnFTr2c0wU/fowfacAAZBKWFFnsasU
vI6R4C8ay4n2HfFyYjZ0D8QVl63VAvJ8n+qKZp+rpf8cRracZ8zHUOiTFV8vLVAH
hFXbeKf3Ge67GzbRKVpZ8ZnqgRT6Gqi0TlOF3/5f1k4hkfQHriOcgDG97rtTSm7t
4MBHEK1VWU903VEbXZM1jqNnihfNQlAjMRVHA9aXgGHMdbDinF9wvN6hPmH7NvmX
lVo5GYyjR+dv359kwyawQUJVhd4/RfTNCG1M60z9TSTZPLn6OjDW+Ap3yO6wTcnG
RCemBm3Y14qBjqrCe13VsQEIVl1J555WlIn9XJRdjbXRfuKKeOZLGfOARMx7AzTp
fQ+aAbfwDjuFI3pUbegeQ3LbFu782o/iKvi7ydrlCFSncAZV6pE8y0WqekrjaJN2
xOiGfvE2jrJJ5G+bHwJaKRuVumivI8MICAV2RzgWJPXZiQPUKCSceupC0+hIqOpE
scTIeb+76whXEJiAhoxuLLOEvXomQLwuXLY7K/zBdlH4PmRqiAvPjuZq1eRpTJad
kH2ASu7PW5ySqUtkUaq+z8TzlVcbX0lXQsWhoYD25R7P2LhcJ/8O4TQv4SYzT3aL
Qv4pG+KWNe+IMfSDli7ExMYnt9x3yZksOZZ+5th6fG/e1QDka6JdXm+G5oh8RuZO
/rYYWo/WK5nD1xB/pXSJPqJ1epajsM86ql93hMqbBSYeNCJvwbVW5OKzhbdqC4J9
3Qtwi4dkZ/Kil07VOSPtCJFcdAXeh5hRr7w0aH6RaVmpKtAQuV1tYrXDdQFNbh34
6uBjO/Ss1nI47rbmsJDWv3BNI2mldfqBdtATHr+uzztIuAFIWKUo9olODX4MXjEk
dMlj4XJm5a9W0gFy7SBprHmvgN1q9oFrqNNBT2R1G1kVoAFu/qFu9neBBdrDBGkZ
4EieBcHGW6OF01yrGaAyFlo1VVP2UqfPqN8ZlM6pVZEg3UYPIrAQzYuZpjoGmlrW
9HNIZH50kFAXcGzOvkSSeQB3tCMGsbnlLzmVp98gYbM=
`protect END_PROTECTED
