`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/4IDSOTCsX9H3c+Uvmc/r17BdBVah9yD7JIgkIcvGCYxhnCMjPjqYrkDz9hVkOkt
0utkQmNXju47rzVlvhGJGZ73o2aw/5+mGsxsgBB0PiuiXHFkpwogiDlfmUSHlRp2
PYmrYC4FUmOL3Gv/6JtuqtwMNsUvzqBO5AJ1o+/xvR1dZErmck6eHoQiOjn4aSY0
15RqvzQT7BwWYX51WaUYfzrXT0Jq9MObJP+mMCg5wq0HJlY/djJBW7yvDqSc+HOL
oAsjFUQiuiqRHVqqYtP2Aj+CHQeSGtEEEC2GmhL5bMTvh8t81iLTQDTxKlIJvxlT
fgv3zYVpU/J+jWRZv19YZ6ArGe/i1jYq80aCHxLgwnT8rjhBJSGKPltcRUjYSLbw
BYsGNY7+r3YxEOnTVIg9A6zxwMvkTDMIgtuubSzbfpIXvOHwESl39BUVK+otUjQR
iVmS3mxbP0Fo8FJYrX2i1bIhQlf0X/K4XOKIpbrPwb7G/mXcCQ+wgj2xw5Emh6YL
0OmYgfPOSkr5fAD2l/lECQPGkM/U9UdJrHB+TuDh6ZEeDn8eSLYLBGQVpUJLcBws
d3m9bLIzqrvUoJTlUjJQhWLxwOhtlrERm54cKZSSdvzgnXG2MFn0y9H06vieUine
l9yGMpWu4t+FDv/SAI1xQ4jPmS4qhyJFezWXOTdxeVx/jJuPRH99QuHCDkWmLwfi
9o8qK4Y/h7yGAvxkVmswFS23YnyzkKmXbuseyPcWF5X3PRNQJQb/dQULP3bBdZrU
auozO90Dv1VC2G2wgu+vpD9f+S/BE5EoPCugwvGstup1sB5wVbIKwjqnTuvptRFM
MQgCuhlxasBdFxcr3N1AWd9tpF8K+yeUA36M9E/J9hU=
`protect END_PROTECTED
