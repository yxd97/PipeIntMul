`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOxW7QBfdmQC1hdzKVMV1ozedvJZinEEKDTobfB68bskuclXvi4tPcSWo/5/jLM6
EkVD6xoafNbi6nXpTSowCBu9gyXRKYdZf51ko4Gxy7H0pKP7dAyihoCetdvXSr2X
LiQpm8/KPk0Cap1SltMc0zIvJae+Qf0dyEQimpRDlgeMJUo4yyuN0OkqFEU0xzT+
bmAWK9n9o3a73v1+zwpyElPPl5QWVdmIDtxO5weLza7IrjoYM2gPaHLukF//bGx3
5kI8Qq6LuSdofPMox7JC+Zqso5n7/yPDwiVJIw93fn+Ah0b4rEjTY7gNz8nRxqQY
sxxGUjS07T0h/86CEU1lGHycMycvUQiFJcQT52/pYCPEebevigkJlGN+2a0183lp
IjOLldMGP1b/Q0jX8e3KtvJkH3BKAUUsZ9NM2Gn0Hw9dZ+RhwzkZKrmJQeFqZ7Y6
Me8eirjlxNmnChZ2yDkP97/TaHyJxlT15otnBajnlJV+EoyHUujw5Fu5XVIUB5+Y
tRyoZUglzeu7eSRo6OX50kkUqi4weOJmx+mheaN0smw=
`protect END_PROTECTED
