`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MBjkMSq2EqYPwbGbmSUvjgN5jMNjHu4PKrLHKbQMPUlHqpmoCCdnRQ0Kif9tL2oh
HKQ8aOSQ9pMam6xYVax3zVOjP2MSHndaRLdGnEems/cnMXZDGVHleZ/YwQG/SU9s
gkKGiPB/8OykBARw+6o+2SImzYXZKFg6s/DnCqwTdZ7FqKnUiLUHvhUjIv0hz6HZ
49oopeLLQd10w2iLMoZ+GgAWSq2/aL7oFIVsN4bRJA/gHF83nJWBsq87pd4+f2Sw
WK3NmWDd+Vbxg9SQ3+TibY5lhTLLlviqaqNC7dunT47KHJHiXZhv5zZQzaucZLBV
Paczcm3+SY0x6dS1tfAh6UDh5IghFx2WOTwVPfLpYTC8P7IcMS9BlFjvv4SMFbx0
d0QqHsb2n5aShLXfgk70ZHt82flcyBHBhFXf5+bueXs=
`protect END_PROTECTED
