`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EScVdio1eiaKRrxOKOQXhMGCp+w6TBAELmH7lfCY+gF2uD857BookTy3cxeRPyeQ
oMPjpxSxFs5DX8IMukkCC7tJ7ddec8R/zzTQ5AcDz47+0mszNqiP8Vt2FDROoeMa
eHISfz0By0ydk7EnjAZVYikXNdmir/ulUQUGlvP7Uwm36SRo1TgZom18/il9Vm8h
OtwYRYAw9K3koX5klgjMxmooP79dWohGECld4YdH725st5RwUjekDM/BoC0egbxW
k4XMh9tjjGY3GtCJj1FAZYY8lkKiKsyrbCP7tQuAgC6awUn/J82LbVpozcysWNWD
KT5vdYHw11qKtGZTZ0nsfds9iNpVAFkyfAAJ4uzNOWOK9LeS3t4Ai9xE6ZKKYckY
MYeI18E1P3x5i/y6e8prVXIfdGwU91D5hE6iPuTnGpaa3TYRnfaq6DomojOKoO/g
BFFWgy8oVXFb5yvCYyArh4UT/w2RgVd8Unu3CdY1GPS8+uuarwdyIAQmnh+HMubY
hZ6vPgqBRlpQkT1Vx76T0b/TmWC0MkvyGMSETLUG2wO/Q6TZ2Gdw3BI41lmbD2JR
8jASBtB1mZHsFmAka8T3WETOxDBU/rGJPRsMGm/TWR4=
`protect END_PROTECTED
