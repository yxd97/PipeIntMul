`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WYISU6gC/VJmXxFY6B+JeYlD+6o6oLBuednCgQ5ahRFaUpiWRC0xvqxDqHiSsons
fHX27U50S5J7sZUWKN5w4F96VV7ykZOdmGQ//XhyEunfDGX0z2YdMyQuCzvcqg1t
PW/pHFVtOuNZQk1cmhV1QK4iKyN2RPfD/S7z7jwYsoxq+xnmBcM0mmexiSaoUuck
y1Xdu5Vh+cZPknNQyZ6GBAXCxE0PtW+3KpOW0+E1XNE0Za8nNuTs4FEEi9b3FJAu
EQZiGoSF/Sop8fzGzx0j0plw/+rgsqtHT9plgzQy0JU=
`protect END_PROTECTED
