`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0v29T1jQNUwsE8GOth+iDa2M7J5zBusXr+nuFlre9Fmzit4OONX3P+BmnTzvPQUp
DoNlWZ7PT1eQIJIOqpEcDFstGG81kKN/uD/L8Y56JM3weGfbin66HOmno83srHlO
d78DSfzWx17tTEp0tNPfpKSuj4FRNmqwr2KCM0JwIHY+YndDqnXOK5kPn+W2RRzg
ePNPhJELdkOctGjZ49ZrRspVqiJz9V8+rC6B6xUTQhfXxLHW07AdfZ6dvmsZRYVQ
DG1uPyKYbAjw/mEgo6hCWYgNPpORLeCWrSyjjXWBLFESY4OqA3EVoVB838v1bsjs
V9bpqZQIi9+iaodA6OzcQtxgnNZsK/BmGgpFHOWctCrkULQw3lVKaaLm2WWFUpwc
PIngYjKNGNP/d7+LN3Uo7oCR/TJnaWMJeW1uKkUOh46I6mzZIITnq8Y82C/nyaa2
/vneWbjr+7Wk7FYGY7gUnu/eIvLI3qBc/IwG/Fyon0Y5skCddbAfAKHup9psrveX
veHgHeBJlEQVS7M3e/xKnbLtxjf9sOkky6Z/k2uryKs7bmX4iPTiwSnQjbKNfnWn
CndDxKXI5AjDXhHitlRHqM46vIPXKDxMz+3yKd15yfNjLkWw6m8pQH2KFyTsAh5F
L/83qG534nhmOVbiA8QZkAUe6frEycPFp88TnYozgrlMw7pVggUSotaDzG6l1YJD
hETTTo9qVu6wVF4PmIIPea1kWWPSahw6KYKQ4YBmDO7bLg1EKw308LA/nwVwY0pk
/dyTygP5+wwRmh2lzTerF/kpLpp7LKYmMgQgVCp/9bYU0LW/Bx2r9Ojkjq19M4/O
6jEuWNqeJJi/mWOYLPFewA4x1JXH5cXv/aPbyCCxcBPo3wS2jVeL++HqWqHTlikA
8B5rGSFNKMXXpc1mvBZj525eaqWMKqJ8N8GwEbMQcp7p+7q0U2am0ENTgEwgcKfP
QKXHaU40m1S9nRJArCvJeNj1oDqFUzJpIGYZB+BmKkEnYk8dJsJYUyD3FpQa3K9I
UZs+mgTkPDmvIwigVgV2c/J37KA8cTgog4YVy8Ry7uMa2upN9Vt963peukLCnQur
WJ7/pM32u6DmqfbRN9t1YzQJ9rKw64vvmeYwdwBg3FM9uts6xkjXMqMdUpKPBdSs
4L3nKmiNxYG3Z2VGN50gueUBp0n/QHv2ZqbHZaC4JH1cC/idoLaElFb0gV6k8iBs
BOpg12L3bSrKdefXoR+niilVl+0NTxYr7VsICnrRpvJXCDX0gcml9PpjJJVXW07y
O7IRaWsgBYiBpPQGVnudmJ3kAeHviwmx6JQT1EFuiEDZguGn5IIbd3aSWnFNvdqo
pNqTmeya1ypgTr3K/ns2MfPqAW8AyyWrdJAIYIikuKZiZStR6Dgh6uuLoSa04dNm
z8Ja8Q9098aYL/9iW2+xdJnfqwRqoNNnOhC9SkBzCz7zBzNaWgF3wKtDdAeviKo0
x86dExys8JUSurC9q2jJOrc+x+G8XeeJE4wvhdrNj9bMZSg4OTqe6J7uQO/Qts5q
mqvdj2RVnsl6MCMwaGKJfb/nq0P4nW8oBMVI3tPpCC50ePhowv/TAa+S/dYmh9A5
SJogYzyCE4IwmjzxgWTaCBxS924GmGYZyoJBL9mCTcH5MCXGX3D3NHUfzlnvXXYz
yy1O3pH7OBgrZ4BodAUelW4pKYdwGlvhqsm6Uc3IZNtGxpEoo0MQdNuapNlZj3ZM
iApxMU28sGwRBttBF73zwiS5oJkk7NUM0cbgoB3+gRUxY4XqjISeDplvkDmwG7YR
kJuqo6l0T2NOmCcsgnhbhrrAHHTzNioEcI3/UNlP2HLQSJ8ElG41X5ErpXr3MXZZ
2bliFeAQ+NNbUzE1d+6CaCOvSMib9fyykgByUulSjf+tTI3KGlykXCDCz5d3tIhc
TFxSL/ZSBm5Pl5wIKPXbr93SyPoUkUzDmfayXIW0G24Q4gfqiJp8ilN9CKmoi6bv
6fuEgBF10cg4vbusY0ypNKwSfgDgDXJMI1zg8R/KLKhUVRQXGPsxq/C9LPO5S+H9
Bh/UbSXIrskIQO6Bco/PPVJEeylniIO2rAObSYjRzh0N58LVaxxhr+kvKlz9g1YI
ClKRbOmrfaS6XcZ/0TR2cVHeR9fWL81TJhNUiT6tZdyEK+aJSpD++CnmUhL3zqV0
9YpjBWzy0roBo7DunCAEJfyFSlxdhqLRyEMaw6JOpNLpBYyO7erzZjh3MRb8gtab
XR0vnY3YYwevCR7KU+PTSWVONvEse6L4Ip0u7XW8sSZWYItBpWy+ebOPXrsvPBxM
jUmYLbAJZA4ZD+V4TIuPZHBjy6M+ZxkKcR69nomcRk3Rsa0biCICMQGaDg70uj+s
Y/+u4saYMiXAg1QmoCpQkFsKPLUFlD7NbDNrgSfSM4OWWSFLaquXI/Sap+b0wtne
AvbfH5+LXZzC/CQ7f1Bs7z85JaBizQE96xTwJI4fUGJGIXqwmqiEXaeDwTiFwoOC
gRcN800ZXzZMdxM5gNyfJTcrWo37qEfvzJlGjU7FgY0fMU3q8CLBmVrQX0OKjnRw
mOzzvo/N0wvNLPXk8JOr3urw8I/PIesqdrZtqlvwg71ebA2H+wxCiP1d20+1J8Fq
qfsOQtFej/qddn3T2nKiOVM0SHIJAgEZnzdh3RC3uPLzRW/t2wLQ9+pDm5h008i/
tFKiEUcdXUf17PG2nbgWQMbvmP5KU7KHYH4ytiv/6ljo1mY2p3MS1Wwkw/9sxvqT
KmNOyBS4n9kDintD59aP3TTrXQdTIe9nSd4gcgszuM07OCen9Heg/AVznqYauvRb
ORrnIBob8AeLiLB4TKdGYnl5Q8PnuaLi05UW9MOPeXZfHHz3Swdb9rHmMn9pLclx
0XMA+vch+2pDvufJf0AvUYqWsWo6KXysge/xNuA16CJdAYc7dBRdbgGPWzeK9px6
r5+whvPEcnKqVTvls5NWR4gSMxf6mAswj2ubTO6ELS5iOuJmCk7dCBpyBYU8o0+m
W6iISu2VpABIS5vDyGIUc2O9notF2YFEWRXlXWNP5TpSiADGE5myndeN8XNYvZFu
EjF12jh5aAdMQg8pFBQDkd7fJBQZmzGRG0LTLB0l/4b9nA5LjBc8z9qs3Iphkme2
6dnqZLKei5JW/OhuEzpwdg2ZBw+nU5NnDjXzHdKn23qS5o3wXFD6O8a9la1YlWJ/
f29AAQlNycS3nX85D3clme3ajEBtc5cE3bzwjyLumnIQ44W1M8EVZatOoE1h8/UZ
HnNdHaBE+4pbOrbX8d/6er3cx4ZzXhn0pI9c6W/Fbif4S65gJjQUSSate1TpCt9X
06hrJh5sg20Q1jxZwuLczU1qC34OzoWvgQDycwTcd1oTg4qLED5TueRxCArDvbBX
zAfLY64Ae+4UOvugwWgD6lzy1DNgWgwGYg4wYR12u3DDbPSg7HOZiUmcR1WEy5/8
v3W70oIIb4iZ29nxWUo1D6022HPxJVhHiOmoQtOddRyD/J+3w/EPq8mGFHf3GaYc
6EyYWePtMuDr4JxIR9QMp5e6aOJ6BkSmeb2Il54zfy48Z28dZoEqicjLC1k1E9tT
4QX6H2fXvZdTMv42z8wfVKsM8gzbGe5Tir7fDcVu2hNQoUyZrUvcpjfGsiYymNtd
jIMLSLTT5insGHjnz1bHfWM6qwotFPkwGegFTo+Cf3s/0B9Gz4Q7nZNQczTP8okH
G21AIW3kYr00ab0nDbrLyNhYkvlFSdRyXxKo5QqseJJ2txOpS4n7X+rnRHrmvV0S
zae2G5GMadE4NKT35rJ7LE5LUbN5j62UG0WFa96/gFpRnBUayq5OnxIIYhB+QkhC
RRz3QtID9Nb/nQ47i33jdSKtlNWb4iRBE6dNE6XGmfl1go+G0dT0vE9Ue9N1m3az
wh23SjSIPjhnTvhS7qEDygzg14vwGzXe5bp/E3nTd+KSIZ7Cp1hoXzA8C0USoAGO
Qb4CFpJMLm3ZkDFS18VvH7WS2cZ5/2MbMY5jZ9fD/G+InjDQxjFsZwaBqjN8C8Z9
AWam3w8SYGHLFQ0N84r2emVNT9L9DRRGv31YptrJKSTcciW0jSplj1VIepGWVbKZ
tVkd/a2DYNbu7g2E+MYOxXx7PI5EfY9kM1aveIgfN1zepbEAnrIzrDcoF3SUFTqL
TVN1BvUxZf5F7B5tlc4PrcSw5vEoDbqiGenRj9PKHTpu8zoeHB0Ozr0kr6EsCg9i
tpFIvmgq43eMM2iCRLgx5jpiNLsYevaoyRUQpPT6LNzUcoBtbNmYL/Lf+A/M0q83
60uMt9RdverLCruw5fJ0/sZxubPiyfpcnILy8LL1O6lbaULEdd3CXxj5DTeA2nko
cJID2s3cM4+TqxuTp6/LEwzOh+wcykW+y4jQ+BZuP3ycuYVzNC9nG+rt//lzcRfj
2Et7qU4R4GmhQabKCvwE2WJ0r/Tf/1dBLwyoNF8X++HMQM8GkZ7uZA4yM4+5iFgX
8EnFQWihj6YEIAKPdBsYZr2MaHvyd/np/E+Gk8iY+ztHVZTgHQW1SgDRkGQlUOEI
VFE/ywpMUHABk445l/3mWnb4C+dEMbOyEmyOzskx0HgtcehgmK32QugEiwMUhXV0
jNUuoCOiVY+R38lmQwZcQ1ywi0omBGhzV8JEtI6jSB77lHBx3CEoyq7yhURM8xjE
VBJLKYBPEGtdEZAZ7Lm5vwGPBF3Jlycdn4ly8H/tjE6DYo5M8oC3ps6bczQagOl8
pPyINrEQl25gMQ8QxoSLYyqYpqgZMhZufB+pUfWEgMTYCFDkyoGQ2GOtLcD/vqlq
uKOCjO/uUdlxwiWGawUTiVYn5jIuUP4+lOHpA1Qtz2ay3mgKinI2PdUVn8qrRE1v
YDVyVNiIl6g+sQpyPtq5WweW3gfA+uMC3EwDbxDG0t1LfjNNvafe4tZNFpphjTDX
tGe9cXYULI/YTyhnJwDkHAV9qnTgGiWSaVBGlBTm8A0k2HXm/J1U+Afol9JP4sWT
AUM5h6zXrXMBWOBFkDhNa/70AD1kU7EImgFJ0+Qcq+zZQ0umc5Q2FzgWXVEaGUNC
ur5p87/vJYwD7PQi++Jk9WKlpcy/bErKPgHHB2fgReNGnTBDOdcWVvSsLmUIfKBL
nMkzljk/ENvQRxQMBuKIA9WRZVZN3aqCvYOeRSKjxL8V/YF8l3XDsUOYNhNzHOp7
fq57y+T8ulyeWeO2yLGasWxXlFX+eubaBCnaSHUE0fTLLQps2Vo6tt9oc+orj0I5
zPXO62MuDs+XM3RDxJ7BmSyqYgsvGtMVJ8SUFjGtWYTvTQSV44wtUf/Spvrh+nCV
h3wi/yPbT3nLd27360Dq7B2JHSikeHqUhyc+WnNo6hlu26LhGpayKZNNNzI+u1SD
eB8Bhq+0EkVc7sZoqYPpms9qcHNyQDDNgFrvAy651bD4pBS06zTvg0SPv++B4WLe
bfnkJORCCDw8cfUJr/8u1a0RaeFW2gb9A17dsOvYxjpqualpnNjjFxbcTNxeAjy+
2CaKCuLPiPGKd4Mi/HzcRqMEhYhJZX5lBv9z3iWgf9Z51MSS8FOkar3iXY+EJhlu
6CyMqR5rT2iLE+2MywM0IMpWMHDSQLAU5r1k8ZXQyn3LlPU0P7G448/Uwzsh6Egl
Jit8DPWhEcScKEIXMRbq7b1nqcCGbMyHeoFdUTlvBe7vIXfEP5eDb6bgUq6ZY1Tj
4caTfQu/bPthP1Ymb9FtVa7/cMsJC+eBAHKQUIa2IekJmogNdaJKR85ISqYUh+eX
P0SK8PMJlNOy6c4gN6+Q+mwQVw7e1mJf1eTyqEgDshLGgOZi2XJZ3VT+kap4Bz+i
s2m8sMI2dLdVMiQJzKgS5qfQgfCd+vTfgY1ZnxpGRGGKR/gmCUEp3UCtX2ypc0Vn
I1riF520EvWs389rFrIQ6w1GxbXXV7cFRGbiiwR7HrHDqOxYsd0eVizzzDL7d0ce
f89IXCc1iEsaJR56Ser0CmryRiH9VzIo40RjrnFDA8pss9u0+DNtWpVitOGrp9vO
5ZjVWElNIxvV6AMUtP/sLk44N9MeMvbvhJzFrpZykOIX9QWGQ+tK92jKpgoeGaxe
YwbUXHvA6Z6rgVhowIiGy5t236Y214KICTmSFyGdIxOG1DbJAdqxa0FRpLmBWp0/
haXX9MqkEN0laGyLUMKSeWKEyXdKOJ+RS8W8sncwAmKp2uwtEoHJfTzjTKc/Ugh/
TTcVHsZdqssHusUICtsphtU6Q3qMU38zeTqTae9MJxEFr4l5W4pfBw368oNzPHFP
/ZcLQ2OCoJzSU0DP8zM7rxS6ERcf2m7SHBj/VQhtxfv0rRsbJXv5IMtzeq1izjxX
fmAJGhd6dPKGhlHRHhCAwqfL03cXv7iFTeWubI6hYwULqXta839vZSyzlhcb4Dch
ZBoaGWRYkbmknTqAoLY4uqnI5N+evE/aHkMnrjh4csPm6cy9rRhgoEcMYQWN6934
qUDsny6F8mzOyYpvjKLyNIepFq+939hmkQwQjwkjgRRhpv8YIQHV1UFi5t9du1Jh
8xLZcY/HoTTN+1rEZpY3X+iViSOUSIRfX5TzXhBhDgz+7k+hShu76y0gFYJggCVE
xtYEBk2g+8Cgdt4kyokJ2ApaepW7FCbhYhFFUhC4ICK/OMCSoJfDcJpqGriEkp2p
TJjaGaYJBevbuzK4UjiimB/m7wRvvhCFafloslO2xFH5x6mLZmNyviSrG4vZpf87
snHJaH8yLPkQEACf6FbejwZIW9l8ANjyHZmB7LhUBBaZ66xvf001RHxmLIfXN9og
NJ7+CwHyHMdRivDL39Uj4A3H2Hpfb8vQq5pYJbEJFkmxk23qPt834TGfutrZuodZ
kObkfwOiIzy3em8r1M1muBzUlkv5Gp7rkB4fqIOxybxPM5Y6bK8gv/YjqWhvYECl
I1HZfqyXmltUo3oe/NkPdPkSctd0jJguBj+xfHNb3NYshRfTtzAVNvrsUjeoBK3S
BwKv6+HnDo27l4pHAQzYhD3X5Xrk5PRgbO+7hhmCgC3QDQPqUp036lVFBauzpPC0
1FTkeWfxW3yJlsu0RVToubeOL6UFbGXpcWAwT0xjjEhkiZbXcrIsYt0agr3C/O4t
SHsXn4MqxKWxU2U17hjTTFVAj6KURzpaK2zibApJwMIwX37KtKevUA6qcIj90Y0m
hC9/rd0jj6tdRGz0Oe6n3qsec84fwObiLkKBXjs4LE5csway8Mn3OvWohPkf8E6F
aAi9e1whRJpdSRY5K5K4Wy8hJrtjZVmzl2YVbq+YoIWOLoueUf2swT5Noge16fcM
ic80860oLUUqfoC7mXPCnHiN5dqt88IqT+RWVsk7GzLRmvpNZsCrslZwso84lduK
63lvxV/rH7bV0EpLMCUXQhGq9nBN0u7/Ue2P9b3ohIflnKX1eTtpS1IZerPuuNBH
FyYZTOIlg12Ox4Op7srf8ECyvGeS0+3Dfd5C6pfYjRibuE+w+gVn0G+tWyXfTCPP
iuwgQw1/P0eM2HfMaLwN6G2fgRvfLZgGhmlvXwZtzrKx8uFr4C4atzqYqn2/RxVa
FkUo8S2eXZvWr/R8oYTS4ls49yCmAxnI7KfMsLz5um3tDsFsS7ICAI/3fJ43yP8z
HB2KScKZTfieHhpw5b7JWQbcQycNm6rOWlE7eME+XjGCSPJ60y5J1a0EyteI4jMS
Zw6dCNuyCONEqBWcqzPCUwZDnMBe9/AaNC37dTX1rkxsJbuqMBBfRN9qWWDQzjW5
mAOZLBH39sqonlJTK1s2nLCTwhzIpxs6sCXM+orp+o7HOp2I26gaZt5fHwWvWFf6
HaQYf2izeo+T7dwb4k5VXgimBGIvOi1FZC4egFzwTropGEsoOGIozO8jx/JXx0e9
YqOOiOlqAX2Ejp+UPKgdEIXgZEd7AuE5mTbNFZTctVH/ibaFHQfiPpWZZ1rOhF/N
+2GXG6HKL9WY0kEKj619YrHmNYD26b2coqPm734jily5U4+ugYesANvm5KqlepUr
1m/RLUoDWbOfjjDf2+caJVCSHWvqDBLkL1bURYZOjarZsM2eaXPkFciHf7ZJlrXB
OawxV9m4gJu+omDe+n3DLWDFtmwJq9SgvmMAczXHeRRH2CUbnr0hh2pGlb/693Xg
B4i7DeVd2eUP6AU+zUrXLj0HVN6tXc0QUFivoMfdmpcyMEPD8B9wbITZf+31GxQf
YJxMFrJvgyEk+f386DGKZVXEetEvjbjByqhPAfBsjOZtFx0Eo/nOpMDJ5rJBwUSA
nwEnGTId5C0c6hY60KPA1K8bKCn+AX4ekaOqS4sorfRq21oVqdCXO5lEHXRoiEr1
fnEmTVbhYllAQOw18xIioQhWuTxNE23tJH1bfi2xlbPhditBjj/YwSi0mJBQ1jgo
XanjJCl2L4bv7MzpUu/d41i/UKfq6UGDSxqkTiBHa/nYx6wNoNf731AkfHgMLdoO
6UTqN75Nkqjl4uzn4CyID0dWfc6fmJW/4wRP6DPigRjW5mnO2TYEvLh64Ck7E/q4
rZuDUMabPKi9QOOqIYpGHAqmdY3djTjLiNW1Niw2wfwBnUWqOAH2cBzaJVOCNuT9
x6JwN/Abtymb0eqO99OtUUaOLAph4sZGSQ3GqlBJO5xkM3GpN5QhIBAuQ1anxH4m
IDwQbcuG4lp02KabhFmldFAxudN3wa4UCIQJYQBs3mOhCXHFLQn0vfklSR/ufA8n
Gc7Sdd0fJPGxPccyLksD42UWWPWrgguwwNBHD0wptq26KVXggmT7bqehdHLAEeXJ
qKwzrIi1oz0MWNBOk3KE8sJqNPBF5uRm1x8c9Tgp31zGXvAHZdg6y1wgUl3rB74T
8Pu6V0Z22/a1A18PyViSQnrVqJSCrO40pE6m2ImsLQDF8snOw1ODosNuF8K0cc5k
pSJhwTAPOYvR3NgS5O9/wR0O0Bz7uVc2tIZ4tZBpkxQFWeypI6JwoW8avXZytVfO
4ZShOF+9qn5Qra81NY7CKusgHXjGjllcdO0ysXti1D12pCMR6Ijb3MhtvdcKvVWY
zK5ZM4NovrIdhmCv9HXx9Cx7Da9XQGb08+yaV9SrapRbZLGzuAz1YPOV7LBtzgzk
l2Pb+i8sSCIQXuLDsfgjV3uInLGBmcnfobG4lst2s1kYQrGipY5Ipam9vERTmjmb
hulcsMKsztHp6xyNGROvSuJFr+2UX1yDZOFNrxyJFJrDOX7zI3ROwsjRlSMLj/3s
tDThzbP/9S/siIWeMR1A9hX6BFEf16po0R5aMNKzm9Q7R31S8c+qz5aiveiy+e2K
I2vOBKafqq+DsOFjWJ3r7NmRnabeK1Y1/6rfJsv1Wx2OL66EBkb85zOzLbQAO7s0
I155DmCtV+PjQma+KdAPcLiRUd/iyrRhg2LXtF7wh7Q2k1cbltSxxfvPOd0x5/EG
+w3gbFjuyNr/+T3+sG3yrmSe1GgVagqR4qnBD5xHOsGewj09wrGu/kAW34yCn0lH
p4qycM+fEyB9frN8lCFKxo5mvapLF9tfLvAhQQOV734bg85dfW92i8XUJDavDPWo
yxuy1Vx/BMq8aJ4NxqaU3DTDDx48e2DI0513Mr49ELSMtHEzAlSOWXVpqciUHlft
bl1+E55zfXHukq//2LS0T+EhxGyJP5sg2MR16rtnhKdy0SL1E0n6saBB1mK0xDa4
mHWyCx+P5d8Kt9IZjGV1PH3upY/Cm6Q/tSTF+rsRqXjJzhtBHA7+X6RtyCJHgse9
BT81LjooT5A0gV6r9I5nV11Y3lfpvx6+vhOwGosg++T4dGmN5XYSC0MTN9VNuULG
nVdQsDCxtp0qacELFcv8k8PvLd2HZOf1EomHQZZh0eGemOEFydYGLLbuVDgx5U6g
JrSUsA7FUr7aD22qSAB8wPiLpKRGLroYR71yW+zPj+eYj1WDFryfyGZOji4CqSa5
UrmQzzE5pNGnZQAmdJq/ew==
`protect END_PROTECTED
