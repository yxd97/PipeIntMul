`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7hkN81VV49MahSBdUyz799ZZdMxcAkrdccVxmOqgVz+euPVIXotIwPMAI8F2aYFm
lA7a+K05XJCgMZREiCAeN5RahnmfwW2/FRmP/0S6MzvatBfb6A8MHB3qD5gBI/gx
EJK9rNy6LXdjogwpfR9JFYO9AB49EZatEWaGZ0xbZ165oMsHpS9Qin8zWZUJ83m5
zMQW7IOHgWOf4Y4jozwSCd1VhwsRyJ9YYxled4wu0bijAoaDWwKoyB2D/Z1aVXu7
QiGmwzlanqXrmAj3nZceCjgltJxlmebWZQWLFleU61ztmRWAxzJDrlJLx8emm7CK
rbpRCwv98sWeNyLHOW74M/JmVEG9sTrK4CjQhNLTiY3bk4OuKsgkRDG8BfNo5rrU
6xlie5cJO7AyBOwJwoyE9EPU8DPFYdQ00Dg3jyDDkOO/8ZAGy7ERPV4+TzMOPRXG
jfTSxaQYTpDyGYWgIFRMqTIGSve2QWGX+7EtL1sWw5xDCjiP+gBdIGI18AdKCcLt
qMP5RtS6+VyLYhE2QD0aMwfvPuAQzURdgjP5qZwqa+w9geDKEA/z81J7octCsJJm
RfSlYjSMWq+XjMVze92+HNEStUa2dryPcDCnZnLMALcKijjArleK/sN2o6N+PBHV
kEE99nH56L0RcasPntIaH9uS+/BdepVISG1yyZwQPZRt5prHAo1kL2SOvXhWi8ZF
N3C9Bfuf6R3uFhxhcGaoC7UmCF7tWgtGuyfkIXrNGB38ervtKIppzGum/XFZ1r/R
2FE3Qekgth3vNKzAoarYDg==
`protect END_PROTECTED
