`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qnovXA31AtFmwaCrOC8s0YHDw31aUbUTkcYbSML5fgizXg9uI3BwWf3RN/EmkCdv
UBAs8t4fhA3Q3idrN2Q3bTC6w99XoJEziHEhgRXbyXGMqIUZuJky8UnGcLw/7Ut9
IkEfCMUrvUGclB/vBCDqpI/nrp4bxgxChuEv+fxcFJ/RwZkOhsRT9tJQjvsFLXqa
FKcr+LWMjtWIGqPv/MjI6sZ0ukn3tq0kp6nP29hWVhij5YnjGNnSShW3mJwaydEr
UJ0HC/Lo/9SL4LntmuX2UBcjxowwTo6XK4Q936dW4AftU8fJCHbGU52/f1oEKMZt
YrBDZ/SMKJUS6qduzasnQQ==
`protect END_PROTECTED
