`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+AOFf3h7ndaYKWS0H7ytpDserPv/QOF70bidwi6OBmVoQDlIUI7i3vJ4pIIhAOa
a2/w5Qae8MvnQp3l30r8cp5zot0sZvv5PvJ04rTUyJs9RE6qOWewCBZDa8GpOZcp
iV9dn/kABVKfSgBKCuibPFcgCNGH5wCbEt53NiM6jwMyVDNNVj+9q/qHQSv+L73l
Ukr6sBWFuRiQIpPs4X9VAvdqmgUK3JEB2KeJJytBJco=
`protect END_PROTECTED
