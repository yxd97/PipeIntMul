`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
449oidHXy8os7v+pIqGDvyVHuSx4U+/JIg4zIrif5kE8WlQDbMsmhLLiJIaIBC7B
Gvi8WuajC+0WRr2acKgSRY5tTFqB8eu2/5v868y6sL9eVnFgJ/s9jqnkNdXFww1E
ztkFklwI17JPS9EKPvqju3cOljmG718fAsrk7N9onGS5SxaKj9sLlmupoulRXz6+
A6rzXkFSz5Izi1qQDfv015ZHQoTGvv2e7SCBrEX+r8wlFnNjo7dU7E9w96JPEB/J
T4hC397Cm9LAbH0t32Oqos9AjBfEK1xXcpyP+hYVzlogMlPZ7vTf0Pz+xs9tw8/B
sFW42Tmfr+/VYUFzz4izXB3CHBP98t61GWa5APaRMIiTBqwnfoLg9UZYmoKv4GRs
KWwAhaQ63VSAOEj4IlD2dr2CQyuKMXVUdualnUo7tYbIh6YYsxO1qU+sNu8Qz5Ij
uXClhlkE+X7txflBPTtrYSzwLwSKJySTbLaQKMHfSzpsONMvkEwT1gSzX17KBbMl
+OQd1FxEL/zm2Q3nmDBIcQ==
`protect END_PROTECTED
