`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFppMoSts7+EeKhnIQxwHzG85puq8890PtIg7EA7hZEy3ddhadOoR+TLxFHXqBjJ
3pk94YKAeEiImDb9xCoAC4y6dXxVgbGYaGm/mAUS022YMUZmT+a05FJsVWE4VJQp
nDDsO2sB9rXVT8g7rOI3WLhVzTpoig4YGgWJqwKS8+zJUtLW1GAFpM6+d8B0SoBT
MYJ6d3EY4hN7JKlyPkbAnURknymWDFowpP7nntqkleELXnruWZMbYMb2O61XWhR4
awgf7FxDD92bzMvhydZkC/y6qxhp1iVyaiSRJ/XNhAo33S9gEUoiFNeFwp9ItzcT
F/bp70cyaHmyW4tZA1mChvpZGH146s+td7Cc5YwJaNHjxSMVX/agyONudC5oR+DV
myBEjlA6lF2cgnKZVfOofJC6GpdN5KCEQCBwth85KUk=
`protect END_PROTECTED
