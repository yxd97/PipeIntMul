`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sDSuMMsLlscbpV1CFcl3AhNPgQzxa6ilzJi7wKtiptxp5bbeTVaL27fGhZMe3SL9
mhIHXw86hQ3rRUFD7QvMfZrb90hJPQUWg/F/J0NKOrDpRGwt9cC1ytzc30YBrkWO
A5rl9NWTZuzRrCaLK6XGP+NF4ahpYY5R79h/B04y3EXAF/obNYbMYqCe6ZONmIv9
GDfoXP10zHVI9uoqqXM5gB5IdsUmtpnxlqEG5o3YvSxGa2e3JEkY/bUZj8aw09S9
p+F5fyp85dbgajg86HB4waTXSQF2WyArM1rigG2TWKQvQfQp09f1mREos5pEa7Bb
GOnFw4O8TjWxCaPrzrQLQwnH6KkIuL+EFSLsDxey0naPu09KkyrldhzMh3kP0G8J
omwEqJp6G3ujefIKgTPvrid2jvR+bw4G5aUQgYADui5LB41eC6KR8dUSpmviZlte
8CndErXhZ9kgSot5YSrMq5KSrmZwq0dtXk6/S5cUWzqaCHaRohRzwUJcU8a8bhZM
NPpiTRnMzZKmylI7EEDsJaumN+65V+FmAaLRVe2qiW/Uy/kQBDOAPq4Qq8C9BIEV
PY+q3ICxy2EkrkN1QKOMWDsbyht1CH8mMhJphe7b//prWVbUIic90oqENaFTkCii
O7id0NhzLtNP1Wfkqn2qiw==
`protect END_PROTECTED
