`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CCa84dlBtzhikEZGwuYMI6wv5drBKF2CK+Q0qZtSg4qWinUXDqwpZm9WLpggySL7
YxKz2+z1/s0zeohvESB/6lY+D6oIcaQDbm4/DEJUIv721J0NHd0J+JB2Ed91oiot
hxYUg0W5ljTemFsSx6+vEYP15I0o+RFrcW4uZ++YZKQywHjxtfWIHKd0erHYkJOy
WxCT19SamYqYMLyD3D5kJAb/2HjdHL3blZ4i1TZ5gV5unS4rm2hfJq134DdyWp92
07IvFeqEiEP86qqZLpiT7qtjqdCOPii+2cVFaLssZdwHGLu2H1SYzFySv4D30h5N
tc7AM8uSbYXpcwv+xLOjEAmrZNwFT68SHCp/Z23+Gkzp+EoXu8TKj0hzH7VFUQIH
j+PZaPxI34Pn7LU82545mk5ZfI/QnDRPbMNhiOYBcy3bBoSy2cUNosstmLVJ5TDf
bdQVn5M6dDRnL6h4yWLqWcZPl+Xz7oa73+Pqr/bZKzxjW+EQfGcRbc11NgHl+IXS
ZJlCmPcHoZ8qG4rVu4eBzbfbCianexD1jL10koHNDgvLbKFlEELr8qPRNAz1lUE8
RqNOAP5mBbwO0GL/1IojTcSw4BhSXe7Ru5iqbczzCAYZ3YI6WXfabFwqFLHDELPr
5nc4ZPIxbhwNKHN3AMqaQQ==
`protect END_PROTECTED
