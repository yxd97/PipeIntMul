`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGucyGhduwWnl+EIi1ZwwBogitV7gK8IpglqLjM+0syafenzwlvQekYIgo8aEM2V
k47nbkfkIBGhURd785FkItaxnJ7nHNK5P4KrLuoZE1VbnNIwfYy3fRODyxmxX+rh
VriiAg7wy7LS9ee86tPYqGbU6JcvsYQSQgc77gX9mvyUAIt7akoiYpn78+2DhRag
jmr+b+AxbF2EYrI62HWB6xKyMzpQ8I9CO/aybE7Um7wO+CXjO7LGWUdkvuO5g0JL
4BvocUtdlb1NwxCi2CRQJryrKcPceBegJMM2z9xoJxGL/Dbk8t/vDAbJKAy0dH69
aRCo8RZn+9boY1KXbUcXwaXl6zy1EZz0CDollJQxPnNxH0SrfcctOpIwHRspwwcX
9b5UtpmMTMQ1x/U7/E7ipqlFwPKiIeETOdv7wigEOY/geVlF2KSlCS4HQDGVcqLp
`protect END_PROTECTED
