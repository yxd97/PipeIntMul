`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P36fTKSnhB5crjPeqVczZd+mGtgK9EFOhFJ6O0/hAdCcbUTXokBUKWlvRfjWS3bt
x1lu9qqCFncjS1h/JqH4esWvlVLdIh9tDn4C8kHHUt29VyqidtY7Ou2twm29ReLI
ZEw72QCZYgesyRtvf8ZO3iHK65BeNORXsiTcv6mUDvb6/4NS1chlEtmftOT8Pvv2
FESRpMncx4MKWegIzVDjgV5FaN0X1cWrjEFlK+H6fA/8KdpnoPiF4rHLp4zjKkGG
Iu6ZIyYiR9OQJfG+vS6x417Lde0yodb+vM6BAUmJ0Nx5nMOgGzY3O2yIOyVK+qXC
DhnDm+oyIrbl5zCjAEj44P3RsOvDBiky4NuQBWXRMZBKaa8t3sNcdKrrxhVPR8vG
sMQkbh0QohNdBn3taIrqobkwfkT2wD9iffQpItSW9zb77JY6zD1h2ujPix5Jr39z
1B44MMTDwHfmGcX8j0QKzlPaTF+iaUfgx2R/ibnp6SWHrUu0Lt8LL09yKNEOUaQ6
4c0Y46cyG+Mx4KVHqi2x7G50Rd+jbVBPlXZeCFkFzkAIF1usOt/W0IHdLXII3YMK
FE3iUUy4y2XmVr+/bYDOHm+3+YE5CDcsovnq62CREOTD+LM1bRRGh/0wiU+dJfGp
IEBKOxfA6q7vLWxivP9ehP3DRQu7w9+YnRp+ChPgAiA=
`protect END_PROTECTED
