`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4L6wADkfcF+sID+3cfZi9CnCGI83HoYLEhKqfcMhiBshDBkvXaKkN5NkH28fDpIC
zG4dbnqVRZmuGygTkOW1xvDQW+PQpvDPOPUduEGPcf+k58jum2TkBeepMsOBWG2F
VU5o0LFRCBR6HvrTso9P1sOMYGQXO2ULYUGJuoXsLvXUwwGzgZNVkpBbSIv7Hd/W
YQMaoGGpok0mTT0+7cZDcQF65N2ymBLZsn3ADg1LNqjJAiqJJPb7YThDJDZGRjsT
1LyYBiQ9G+Iy5/grI/S3uQ==
`protect END_PROTECTED
