`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJV1LpdutXi0Wyx3lHQ7dDTrdMrYFelX/dTPH9yGgomUyP45xCtJ1q7FMTErz59n
7XFePYJp3aYZfUtPcV7NDXaZu6ZI456F3V++NojvPtqRFEjTaJTkuI/da2nqYmnl
8uFtTYz+Bzd9ijqtd/uevRiM+b1+Gptj9j+Ob5J4uPsxkvl1hDSjrYfucTGwnTab
E9qA1QmtJFows3hH3i5kZGSuicALkbUta/TNb5m8KzlridOihJaO+j4n0Iusx3Un
cL5y7p15KGPK5Iew2NZ5xIwIZC6W4U+g8Fbn5RcZqfvHGVQJ/U8tsgjjPgOZ7tjU
tBd7WszuFeqTpyfl9SF5qPBA/WTs8fZsqti47Xo+I6IjXl0aPWiWHoOelVNFrZLy
fn3EgTcTY1YIyEgrFIEoKPlLPEIXNBktWBx2sfShZkwWkOpk74ZKlmN7A5mKt6oM
jBtxvIn9coZm0ODyNfxDu7vdliHtW9oihm4+PULCLXdnTvgiavfy/Ndst1D/Vu+1
9VomgcclTZB34JQnpI4bO8gsicwYqgawz5KjD/ljtZewSYcMWVCnGgig12Gomb5r
55WrO4ln1CPEhfvaF31/bpgR+CmaRcLuRXDcmCk+YzkANunokAMOxQCkQRIk0zeq
+oyaY5WGIigLo3Fo6hmJwlzx7IlSjgnOM7GEAeOoQ5Clz4N1p1gXQguq87yKaEje
VTRCadb5PYgAh49ae7hvNhC6FHBgOTUPaB2wxI64vU25HxAF+X9aZygBfaFXHs+J
wwsIhFYc+rGJlL6HNzaADSU9/F4GdEJc4VrCrnKb4GMKN+KZKJmn+eEoMPQeZMaV
arZFStdq9UJ71ILi/1I4CB4ip+09IDM17C/WtsQUPjQaMF2tUx8c/Nf4M1VnJlZG
3jy9ptiR0NiYPHhCtHcOYjYEZ42bEe8U3F5MwcWomeSbRP41Kv+KNBCexa9e6lSc
ONk+tutoPLZkejbJRlMmVavq3glFz0jW5VrxVGoHEaOzW3IppeVwQOaDq6uak+6I
M1b7m21wx/LPZVQbAujFFihcMfpNNY6OHMgs2lsr2ao=
`protect END_PROTECTED
