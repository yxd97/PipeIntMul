`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vwry4W2lGDfPILgm9jTwfbxE9KH1L85KF6Y1fhJ8wM4IWEVvIEOIWhfvU0PH/xSX
fsElvvSOyfwsA2XmuXRU7SWIUJNAoeGsQYYN+TFIp4hdC8RJLYSMm438hVTNYzfG
QW/VCXx9yN1mXLu6goeUAJgT6o7ecieuRi7Xo6eAj/CJ42PERMNyiNpBSnU5RiuE
YcvHTYpxn02qnFdATvMksJ97jGTK3HDc4t6Z0P+TVjWtm6MFcmzYfgAmQjBR09ON
KbiGT5SHU9KineHRrDs5KaDFlrMzMvyGXi99kAMiPQOPopuPDvaWflPv7sVJI9K8
QTThdR85+vVu3mryN+2CIduq58MVGxgLcwI0bE6VpRWByGpYZ0vPwfMAS4fApkEt
S9yzeTANS0vrmQxN3W4Py8wdNnNiqlDUjXztN0MKz4g=
`protect END_PROTECTED
