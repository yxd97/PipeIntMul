`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s33yYZALylY7Gnj9ZXNFKVBUkxTUjxlAGyx//PyAikl9rTPrGGHRoS08x2xfdGZ2
8lid6LMiCP3rNh3dekxzUkTBP5oVuUACACrCJE+iHsmg+fB6ZSFtkqqlMl2UTgmI
0flSFMGoWYpQyxzFtjUbvohU7uBVYfXDgYW5cEnQ5BZj57nVKjm4k8T6AGN3jUuA
7/76rDTX5Ew0GuBFyWPDsKVTuqcZxZ5TsRkD0puquR9o97TrFGzi1an91V2CXmtH
jHf6xtA/Qpz01kkvDoJ6RtCobY9bRrYfnow8uKbu6WniIqprmEit3FTJ6noXR0J4
ciYW8wbeBFGzmuceGnPUBpqftaFzpm1MNBS5cMBz6/ll6z2rQftSWG+rIAaRCK9H
K9Ps5oYcUrmvzsS1r3ykPHYkAp4vLOxAF1gjqxBaCwxAnpypz9ayu0bHsTmxWaTm
8fdFHAYcH4olN2zIXl4zs9zCsSfO/XDCnKsay5eSWqO4BVi336ougChB+pycGd4l
xSeuLqx2AF2cUoprqjXl5J0rFFJoJ+H42D8NrlaDch3MYW0E0NDGAtQppATCecKA
uU7TTc5lmVoGo+vGdzKvdiGaLR3HMK7cAHSIOkipxyvB7VBUIC7uFfVumDRIgM31
0r355ic8kDipmvJvpGC5Un67HAeGY+MKdHa4RUm3Fh6D7WjLemiWzXW3YhR3eZc0
B/RrK3GBsKEFSVYUFyQSUU0TSXNiZNHvc6/sNMt81Q4OIxWRTQQsv2h4WGXLCYTS
t0H9rttYO6rao++Jhq36Iz3uSyf5XFVLJEnOSPtD5sNjMFQCRplAf1MreFV3x9jB
VfgYVIc65aHYPCQbYUr1thjqqwz3QSkJ8LPK6I+bcyNCeYWI5J8o7EJbJp1N76M+
W5ZDQxeiVqIpXwZ1KTw8GWaLAxez1RNqqg0v8diZLUmo28Ecanq4Zp91OMM7pPXE
Chfrlr/n8ZItrqVWU7XOEa8M0mg6fmH35ESK4lVfYJD8r7w1+GPRW9MGDz1qTVr0
AaR+Rf+oaAD2y8ZH6UfIQcFQD7E98dGBhGoaMX6/Mufx9sroO4KxBGs62zOmSyNB
zE2jXKsXvHLE5nSaHIWfdWXjUqoC4Wp5IU7jp39MaVdXSqBT3shc5dHzU9hEmhPo
p/eRiwUYiNwTVBdyprJLEIOtlMzSiIssbVzIe4lv5+lXFC0Jg1wEWLLqO0v1adEb
iI7nYXalF7K+LN0ork0cT5PTaJtT9QG2FQ5HYd1JmZnPcujTch+yIqoJSwDB9JUN
Me3nqEgtHFrHvUWh0j7OIAAB4jHw2mYGCs89u7p4I08yA1Ld5G48PyGEWFhHx04t
bU4UDqLzJhaARPUZVvJ2rnH4bgwzBsGEJ8AX481ZQ/B+ecYowR8WDaXrj6z5InhM
8AHogC08vEAurQ+k6kuGfSnWVzxmoCtU9VWEliurdAoPN7zkmNGcSx95hl159Ru4
wpJSKfEQ520BXb0tqmdtsfuYDvJtr2kV2dBdD5mKhbur0JbpOflqz7Um2c+EVDHa
DAw85vTcwUelafAzUdasxCnJ2smfj6irjbjgjfcudbuW/u4o4S9ZTT+zFIR+nAbT
2sWleKAR2usLUFsIvb1FILYc1zhIrhuB/OEM+SdyclkEG+ThrgvcsjyZXjfXBuxt
aGNY5NFB3SqaRtt57DK/hryspe0Iyt4T8PqTgAjlOm20sfrKtruZFa+Qk2JihXmh
1RQCDe5cw+PEKbA5/SQ5lR4qdFMi93LI7k8PXskU3JzSizhNsRtM4yzU9EFhdQlV
vUhxnCNtQtJvJ4lwTaLzvO/kH6OmksZR7STiVnngdxo/zBiFmCWQTT5iX3OpDHYc
MyYdzEGvXqu9KgfvSDLJv5I8Fe/bjEMlFwsFWbdaDxu0aNqCJTa/C/4Psran5fUZ
HoAn9VqwM7F9VeJaxSxdfBRObeo00sYdWZTYLkyKHD0pXKxCzfYyuvqqraTlXZuK
Ctr+CtzvucmWCfbat9O0NwXo8pDraDGkg8u+AZ83XvcDfJ7NRHsvdvrVx4eRx120
O2m3VHzDsn2fmAl2SvIIAjIDZ6Iot3FPwb4G2tmjbp7iuGk3NKHxB/ZYC6l8KIJG
Oj6233GXfxriJr8wgXHOYPLRklmyD8DvzfFpmrnpi4GXaDVqq2fHJyu/0+c9NbEr
HTCArVHzX+Easr0GiXGgQK8rF4oh+i1SZN4mKJOn/Odb8syV9Jxy2aE9lqnEbPb7
t+0Gp8mAOgJZuKI8DCZr+mYxsep+CEmjA4R3S02o3sXxKwIMBv2ZKlvXZwjjIyo2
ylHHssDdwStKCT+1hJRKbelZV7DcbQLq/J+tJlDMYxrdiTLnh6E2NSM/zXqqo/fx
sPsYl9WMgoRu3rSu9IBfzbkowyHHIMKWJPdi835PggmNRplhPwG+WOdwtY/iiOA3
ESOPc1ELhzHQfGYcCuPCDhbNgyGE8JFoeMJnIvGmaVTWQ+1l3a+fFTM8Ueu7sgUM
tOfKv5egdQ334Vu1zOHbnFSwWZ1b68TDlVDEZdatq1zonvZZJoNaCZZ0IyEKeH10
lhQsiO/P2RYCzkHyAfAVhddGCUHgzLAAAUebZ1MeJuLuaEHHTTsQRQv6nkvyf4wm
IyIpCBtRZB79ZqrzYLqRArusSj5Z33hcUEKpu7G5l/6DaHJOKwyJltSAPoSVS6B5
7fy1nYuA/KcTirfbNTLl+9W1rc2HNboW7n03hmdCOG2f7YJufT+mTXVg+R+LAxmA
SpZnuRIy4JY7V0ZO7/cGf1y7Tt6aeAElAWuo+O0B4mbBsjpjlHkMRZFdIAGkzWIQ
LyIg1LhixN87tL/yHyu4aEFffDSDacg+D8WbejmaUdTiSM0u+j6+FG2cc1dEEspX
HNvSk/H0qkFEajdoghXmpFubMzkZZmf/Am7DaAk+QULP6Vn49zyI7KD1iWvrJvVV
U2NxXzOMVw8Rql6VJbJAHVdd+cv8u03HhzRTBE4CjwJJXMLAriHQ5XXDnvCGLY/R
WDq3+VUdaUiWX+cG63EAM8oMOoXZncbz6jR3JfIYC/ItdvvW7cjxeWgkVfh6h2Os
V8mWFRMgZdlS1s5nyktjaCZpea37nRw4VjbIE9xggQUmiwYoGE3EtvN3mkA9AUON
piaZxM6NeGSS+5rrnki4O6tQBcIGzx/y+HIggg8d0Thb53L3e2EqcTl02kH6FdHI
wqoWols6lHHpc7lpJ4kmokiVnY4535XXZpSRxoox+4hOp+kP2wTwP41Wgy/S8iEF
zRYzeyq4iYpOM2vHEdrnKlSxoCLpERQ1I1xQg+ELXyH1knEv2qZgFtDGwfvoXP5V
j0939Ub+67vAw3aHn8JLfpoKLH63hsapeOw42GXlCGyJ8sGav70ieGrmeRGs5OoP
uTzfLSGG+KP7bRKT6BGfS20s3fEGuiERvti/5QTMVOlge7jzHV52kGXe6VSZh5bk
r3n1O9UIK3nbvmFCUOYxvL/PRKuiXH0GJwAEKpt9TKyb1H14vX2Up7DojE6DU/A3
wyvpe7g95FpW0DVQKpIUB2t2FOQd5gu88pDHvuBmkOdnOFZZNXUxqVgCV/BBZfDl
od1uztpq/617p5yfonb5XgcsYrsuWHK+mtZPsTZp/4/My52z0hubuyBdL/KijvBw
1vOrl8p82zKCMgPNgWJURRjgGbe8QEYopYcUil/6Glr83u2uTPOUFVGzJ52c9kai
/TQPoPp88CkK6n/o+yxyoH1w8cfx1WZhbN9A73HwLXCY+XG2/Z/vUdbKyllR9/Dy
dH3R+JTq2ISGGvv/tBnwPGj8dplHRsfCLQSYvayaMkAUfVWjbpYwAyucjH0WVGnr
mr4E4JWeMaPCa0w/pVvqciJJJJEvGbY9UMVqxKFaFBb3OjYZqFKMVCqvBPyRqBPZ
iC613KwIe2BupVSHU1VIj+2kTHIej//9nAg7rLUDiereBf3k59MBgh0SHxkwPMB2
jgU07fn/QxO6P1eqxk9hoCw88/4MZUSsfi+uHmsCK6SldH2qoOeK2S3OhouwZPPX
Nm9nWPq37BL5u0CoWkRrrxSrAoR12aAZpXYB7031MefDaefI+a3TFtKIkfqyhJPV
DR/FI8SiFUVOAhRfib/vTMAc+JR8er9oZEA2D4M7AtFmQFwQLmoKLiec2BpW2FEn
Y9rossERlQeG+wyno7m+nmMn6UjzPCw5VIOUKOSfPcz4NKovNXbMnPuyvvciN/Wn
g9jPnzeQfSA5mbAC2/HQyR8Y9R1sQx0Q3hkTp0KTXP3K1Q9Sg6u+t5vX0unaBpxr
jLRZHtU3pzmw63jONb7C+ry/ihZC3FJ2wCRVNgNAyIc8xFHBQmO3uYY0VUyDct8d
jgFsCfi85R0gxKaTV04/F2Zs/cf2EoNT1P1nKe2g/nJKZFC5lJX4E9o33PZMb/pP
7Z9osVuxQyjXg5GKxIkMIVYOW835KhnopTurnwYNLx+LWaLNJnoNhJDRdGeEbp/z
EISonrrpmNMQmHxNTKFxn8PTiuFI2pD7XxbkWX1FTkZTIUmIJ4BUW99DnmPbz8uk
cxoEK8UVmT+DGYQtgk6huTkloufzMFjMHebaXQ6QzgzkFvRSdZgbSr9qqJY+Tsts
i9yGBtn+9gFOfuLwKDLZKB/ZcHh+MAvYUmNEh/tFMTv8OKjtpheLqZmrk9RByX+r
YkhySJSJl0ykLA8sX7CvuKE9EFfeHod+WvLDGq5NjggiFTxT45kGhs5mgx18/qLo
tWyPpcE4sl5o4ADbWkskDN9cGibdg/XvEU2bCdLwUwQSgSEunaJPBaLb1UbzcfBe
rowJum/gdmhW6qimKxmJWJqNZN4L3FLNptW6ZXdHGt5CrFLr0T7UWSrf2PdWg51z
jxJxXNIL5CxH+bGW3obg2i1jI8mGM/s0KhG3ZHhU0OHNOBnAu6PPCpmWXRN0gfvs
w9Ed+ihv9Jjqo/IM04zS0ztxN9fyVuQU1pKXw23/6HEnZqDtFNaQNvzIq/p7Tsqv
XPWGyIYqWHn6aNl8nprjVqlarzgT2ybzYUTrv4cpu0WF2WWRkbSscYNyYUgm9wUQ
Mxxl4vydgf9p9wMesquM4wdTPFEljChZltPVMDhzdG2oxmYv8t5dSo43soYweW/w
urptyWwDt0xYQJ4blvFsr5Qoe9w3oAtkIC+JucekTqsGfP/hwjW4KMoQRhmywpXQ
fVOZON7C8vM4SaUffmUoSpscrHuMxS4f0rrqc89R8d5FnbdVl2HRWbT59x0IUuEH
8+7LBkAuXLhUBytV3BHDdM/dH0iJPNPyFnRz/dv0fjqMUfaFORtx7I3L+nYGy2fB
7HNcIGvl5K2Puh57fygDT2xgY2QFKWl4UNYmxh1qHkXIpcUM6CGVXSKW19pQR9NP
3egXO4o3E4s0tGrKMuEy1riTFtiherDIXq0RaunCb+hu88SxWYeKUwMKZPzPPQ8e
n5yH1Y84kkW9k21gQFZNKrHyd8/Cy1ul/9saCUlIr+F58A7Fy7aQTY0YKsdIcMeN
IcN2c/mN8lqMr2sPebWPYmludqsC+MB1wYZzACuQYRSaJlgx3phC3mM0C4/y2j0z
BK9Pw+59RzWnwkIwlrM6ELuo4MW+L4eZMUU/06SbDUTDS05OhMcxIBHSVUmHXNO2
IvsvVt5bj5a2bYOBCxiDtbpVjhvQNcwhojfqzdvpwi7vJ3qXop0RxA5Wzop2LeHG
SwIhwsiwJhO12he4hJQtezmq0WKAlNpqIq2yTPlxDtSaj+HtkcDBQ2D42e71Ktsk
zt2zSDpoiJj4XiD2U1Ii51j11aMntaQgGADeSYPdT0HB9re/rr4Ydjri9sprQTCm
Y4V6dBdbvWhxN0LX66AnnqSI1THkXJ/iPAL5htDIxxySfPvFmcCyQLkNBG12cOTj
l8Xj/Vomp/igMVedW8LzZex8J9ummcxTzTdcntVUGTcjnE/LlmhE5KDnzwECHsmF
e//GwIQ+0VLkPIjPN3wPPNqo/meyKEjTVuIFd+QPi79ZOp8awvwT7hk3vxre54zh
7OUQbCVOiJCp9SbBZoa+gq3ByWeJYA1MprQ5S95U+6TxQE17O55OvYjhFDww/3T2
02NCBRKZbzPPh8u/Cb0t5cJykB30AU5RHa6TmM9GEMmvP9YvNaq9xztqadZz3Zz6
NKRwRSFAEkEsT4fZ0orYDc0r/KPCM5sJWltyLBsn/x6Jfh60Rhm3HoA2MRYnYP+z
jLSC9KeUu9jndzwMfcMYNYIUFfTHRGn+0jWbF77ttevK6kqLwgott6qlmyuTgrh9
4OON8QGIuduKc8fagCWN6b+59o8QMBbpTkIhQaXrfNy6VGyvtcT92QiMa99CJTpG
kkooT6HcmBL3jqdaXthCPCDjZ8T8n7lEmG7T6jzLTHfGgqynXwWt0UWsWV/PL5X2
DUTWMNj35oqwIrDAV92CXQFNbmg0gnKwT/JfPpJQ2ZjODuNDydWDsyAf5akrgPDt
vp1HCyh/5HFyW3Y2P5VUhtPOmjTzfBh3HgTQOFLUYlY4l1ME+zcsGhoViYK0OUou
xd1geOGMjjMMONGf7KFdJNizTBcKPPmHG2/nb2Tvw2jqREA/7g5CehUD44v+59mv
M3G0CYiG7/7edotq+jVNzN6jAZFxywwpu9LJxuEcCwkA1tw6IzK9uyAvqAAgSP1W
PaCSr3NjXKtZt0Uh0yRqvX3gCer7tEh+DCzj7Hkyo/tnHoUk2RuNDrCiPCqwW9LA
9UE6+0Lc7IoP7r9ZMEvuggYnZhBTJbmPBuBQ161QRzKGqWqcbL2IMaZSuWLOBPz1
BbFxm4ea8eyTHzupVec1ci/IzYRmx8Qy8qfWAkQBVHivG1pyYUVeHnjUW/KKkCZb
g0qp5Anq/LDSBiIC1fwlM0aNqd8mrvPy85xAeE3hZEpU8kZkEwMb8HLzVIuzHYYU
Jq/it/wWzOP84AGwqEphyZzjgTctSzX2yRYouXn3AjowdZgflCJ6duqTM5AYoFUL
2Pb8oD3eRO7QVRqxdcc1UN15Q72Gg1DTMJ8NddsNT2/fWRAKk472OVU5nwU/Ea6l
9RAwd2OjRDkg1e6vNSoEeBgYE73r/9VsYJx0cUr/l1oPXxiP4N4NUHDDqOMlKqG7
gGn8USG+SXhPp3iKxgpd2TYZQJPo6XeRKtoqsUnf08Il898eB+om5PxWMgDFl2oc
r7KE4XlSXvuws4vfYqOOt4Z4djXEBbSbf5UDcpsLVTA8N5LbvxRVbZWp5jwhUm1K
vj5sOVqyUyvhnd06Wl95f8Wf5TC7TcJM3svMRhPk7FL10tGeSbv3tqd1t3M3nw+A
86CcQvoHwp8C3zTO49HthmyAJLGW6OB9PeyKZF33HCDHR6YWb0g/qOOCPc63X2p5
Uu+KM7ZoZl4iWnpwcmY9MyFtaP6OBDKw+0ikU873Ko3EJ2hwSSdWpbBMuEx3/0iX
6tG9c7/NWCABoXnMMJzvpwkXxOmMl+b+gCysrBB5XoFo8dyRQA7w74Xhtyqf58OX
qYz42lwUthMxbDCNOWLK/2OEYfBlNhWHRbiVuq1H1cDR45GuHpPFmkavk2H0Us0/
gBEyWKvDvJl/9gk3wOXjF5lOAU6QmuXlCz35myM7FtHkAvRaIuJTQSCB2vFgML32
d8GsxHkv/xLARVnJk1z4gRQp0iWPxTifPdfMjSdMPthxunCxzew0hTNP4OiUzvgZ
alQV9+j9Se019zucxJFeFGZCtlgCisrBP+Dpi0A/z/YLBMsEJ64K5XXIL14J7wyd
czkeVMPjpECmEl6pxki5czaKmnJgwCUaNaXorfdwor+9ZOy34Ni8588f5Z4O9dI0
2DHBSCT272XA63CzTjUF+M/agRri1dvpqfVMKvydIf6Zn9pfH3hPUWkEhHNkGvZf
Rp3arWS+Z78ryZ41ysJEzAOvG050lcl1sgKizlOzBGNv09dT0qKGidyPZ7FVgSTT
bac4E3wEEcip3+gte6hnTH8SY9kSHZZvQz6xMxLk9CCBfw6uZL8MnJ0t25F3nFLy
/eRhSa+pCU0AwoH+Sg8U/IiuRh+xePF0pMC+BIpFRE9UIxHUuR3XiEBiGvvGC6ZM
1hmdQof0oFyJhK8+bEE/A8x0m4DGlzFEnqCdQp5M0g63rw/L64hoLEWN+LhDgNXn
Djd68TR175sk3j0DddXVmZG4Ln3zqsfZ3FrUoEpgbAOz7f13v2e027gzdH1u9jrE
GipZIi4r8RyZvaQ4RozMD6L5fy0MIl6/HF0SsM6NdYYJUb3hB01h/aNZDwoSAdYc
CpP/rKvYwtgXa6ubC3CxtMhuZ2PiPZkP+avWhtMXJQm2R1OHFvuCq5dmYwYi71id
XkC8iplTHIW6EU5CtM8ix8czK/cLd36lPH8RFffZll9l3xz84w1J7ll7qLT9vftn
xdEqPYwUdNuxyxkq9IctZvgThC3fIXd0ieOMen3OgF0TnjOtsFtfnGi/Cpzurt1d
xTu1NO9kAncJuoFer5YKX0Ola/VcYvDQ8LMaCyymVZNWlN5t3SxSLIhoVN8gUk/p
18ijZuhxoo0ad35OHFjzfJnIVnihNWni4cwITJg3fg2s1Va+WbPrK37sdvIbqyR3
RI6KcEFKee0kd+4FwJwBWq3jRqIhS/sNep58nWxoX6aoib9H6ZOybps7/YxsMawu
u6Ubz3t9vmOmeiGjMWDaIY8svmRX7+7ZOccbZn2MI4XksBA0M1wcgd+LxYRE9wXn
RQolup3kHr2Jiul445u3/U5hLQEstf8ZxzeOXPDbIbRuCPOblj9mDNGyuhFxo5DG
K0KgoZWybWHnjp61GDS2qHFq71dWe2DW+lgCStrHXc4ZkriT5/3YefFgLZoqfa55
UrlLnYCYwqgKZAsjp6bP3Z+q5kb7VXgBxjc2dumD0Atfg9bqlm5Wsl2jf3C8qYBg
fSaoInEDZEwbcIALIqbyvRapFOYvWoM4bPCwqWXotMaUgFKJI3UZsiRfE5pdDCwn
UNzybpedMb4SLZbeuy/WTmZ6Rx0Rrr0kNFA0lhm8H/3ASTM9U43w8mhNuNSIgxqo
/D99b2wx8cz3cqZWHMk1VXIjns5ti0fg8wzsJmkl3EOkZSovarplB4mt04+YPz3o
yzkcniA6gC8EwmDx3iORoSHh7ODwr8wbPG8PQGh0ZuSEMOrMnsPcCCm6hauJMIJx
UZDCgjPJv+yByd87u+FyYJfJeaM7rLF0eo0Wts+x+EybeaVEDodMRBlgSfo4Rayo
0sIeEKEUu6DudguWyDwEMmnTtzj4Gg9J6yqI5Pjdy6aXyZNcb8svhRx+GreG+oTR
j08KQREOsFJ5psCGdQz2iI9AMSeqi0uYPlcx+40sDaYWAIJBQ4pcoEnuNENUWMtZ
ehGQ2cbOWA52Zg9iJtkMy3VoqZcjpwFiynJg+L+TsQYS5scSDOpzsnXZloz4v78V
SRF+5lsK+kJJotCO+On5gnxxxgeq5Wqx20LDQi83nMwko4w1Wpc7JEVAmJK+S+gQ
t7RdkU0HJgG013yK4T9HPiwObZxUgUDYEKNkN6qoVyaKHgUntXBStRHCxuAcshDB
nfT855rBrLq19AdSWnX8XmrP5wBt/0FQqSx4qFJ7imqHdYkj81+WVHsxOpTKTKb2
SDTQ+a0bJdkZW+j8Y61RYS2UiJMl8zL1Kfrs61lpxGvaquBuGecHoNz8WzqPJ4hV
HyrpCmlu/ylwvr4QbdNcEnm4U8x4awdFuiXc6IDdKbWDVeUTYQGTO3oP7vuJKWXu
xPBsAE246JcxQqmfOE1CpRlAal6L29/c9YKQei6JeSHxTfHYv3OvxNZKOVe8s+Ly
pNJanrTl1EUzjNjXvmdDRM4be1QPKU/madlLEb+rxSdXzdBxhD2eXQlIXMBE5Cw+
NqtnZ1AlRGN5kA6YDNsuPJEWgpA2CuABeFrHHcsDZPRWCQiHlzv3dBNn4ECdPU0E
ibwvhRBp27oQlM3LXy1d3Q2myQhdr0dlxyYbmVfOj1i/5bxQZKuJ13MHSd3KzEH/
e0qy2Cmok35iwAwLmG2x9ZIRE/HDFBnBYctsejISpVJeQ86orDjd8YBP7eSD8SaX
/2pog0vwbUI0LNTYOMkpx6vL0wh/uEVI0AG+7G9/uPR9qfjSs2LntSYn6oPACni0
NSV8aUX+Yp9MFUgy52E24UqqYdkFGFg0MXI28oEFE/exrrfYPXikqy8o0vS8p3cm
Zz3Rjc+9i9w9rcV2WWNms9zp0j3z5xYdD/Nq7MNDU5HxC9o+qCQ/lVMYxq0bS+9Q
PHqog+o5Fibtc507qIsEiesWer39dx223JzCvZnkddUZ7QoLYpby0R/nzIxbkI3M
QnpV0LO2IKGI1oEaJNT4WkyN75BvSRsI6q4s+Z0EW/RivLEwTZHHCpk7YxE8rn2R
`protect END_PROTECTED
