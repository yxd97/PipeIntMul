`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qMBSomShpFj77R9EuGadJbDL+r7DnCQBcoY9tVEKGtNlhl3mkFpaZFr/tDicEKey
GMOJjbYa5o0CWPktpveR2wpJfvG/Efs/NJjxWJRyRFoqnOj6P5olll3O6xCiflbC
MQSkFu2w5TpdzIFWMloZiGqbOSHZ1WF0r5vNPwc/42l5j6ahHpMMS6s4CAwZt/o8
7eNllhxJmJrYrfT9UGuqcBa7wHZF7tOnBCQmQ6Z+03OPZZ4J2VWf0yQyGC/DSBNs
Qn76kvCZ8l6bp7R4dM/01ocVjL1ICco4dcik3CBfO/L7YAlnuRDr2VHHBwwvcmvI
jfZRw/QfFydsvk+hCZi9rgpctUxn/WpeOoXVVUMc2/0Mbr8MKZdZ5vglkfStEoZ9
`protect END_PROTECTED
