`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5o8h+P8okjH+RxzytX+wYnjGpFe2xnWMfAbq5bKMuBS/0AiK6gB/mENFpDGvpxrJ
6CUd7TVqlZfi+UNQZFcDuC/nAlC3BOlx+QCdMSKqxLFJqc5XRHDl6Dl3d3t3xAEl
IDgkO/JDz35y2ZpzMDm/J/Y/JhoaO4Ihv7ZYXBaRgjrFwoZDP1/5phv4z6ehChZQ
rR7JHZd6G1qMNXMXFAUraeQ4OkddoINU31c4WD9s69cHa9NTPSfMbSmVgHYM8lX0
4PppcYeoC3elOCFfT8tk/YT81lbGjLyNQWGCmaj8wQLaN7oUpZdCZAvkh4UhwksZ
E6nsqHs2ZZfKTV3hCkllI6vwjYhbtzTzlkdxHBUxY9S3a1se/a2fqfiXeo7XF4qL
1T24ExvgdCGvmbqQQPlQYCNUXGMIq9TxvgYux5TG1GR7PO+nzA2SD9+l5U7PnZaK
JPn1eYVD32uU9MoTmMkWha9YWqBkmLI4XEzeuk4HcpCwEkyHbxqAP5Bt++76VaH8
YLoDIxzUmTwt13l4yTsYLW8SjZ1IUCFmGchngU9BioH6RpHQOCxRR+oKj8reps0k
twsZlP+DNClC7CzFVx2xtpF8GEyhSvTNeq6auGEQZaM=
`protect END_PROTECTED
