`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgUeMK/xnoVmc3yAyKbg3oGUInGVOSndYcnJYSSxaeL1KHxeClXI2fOiHMvXyNMg
f8oTpijzcjT4bcUaO4LK1xa2XCWry8lJOV9fe3+Xd9F8KfKfY/ilKKy6nOsFagEU
BRp1GuV70rO/yuTQ86cxENLnzNdddrhhYoi8w/+eNf7D2ru0wyvlN2ox+i7DATjt
1vNaLMm9jDXHh5IGis69B33Tgwzvv84TWvdbM55AOEQDydnSW+aQzjKbHzm0JA3w
JokzivNZPR1xfCySG1TIYg0o+TpgnweePYP54m+E2HgilVGjlvinuX7t71XPhTjX
avLqusBUTXeoRJtEDkSlxDv2ZSDikJYErBEPfDme+BmrnppUKoEq84KLL2U+RDlv
dWBynKtAi/j9X5PUbQKLbR5al0dKl8L4WXuYWfVSh7IeCrdWeFJmOwsGBy6O5mg9
esApRpKY+wc4kc4a+KLYx8ROGt3mdCZ9a3XWiCfIvsiFXsGRRj/edyFyYlOKsXpW
MzLWw1xTnGXNqpoD1XTBuyr5JRrjWWwtiWUqmEFNbJKdwFQYy6BemmntCmoQr0Ic
++9gKY7GpH5uSXbUaim40s6nx+QQ87RUrF6e7lEIR2Ad1+IgtcYSzH5a6ysMtAPp
u8YcnFA1m6ghqdQ22wkxe0v6J7NJbqEHg4W7untujA/GinPobjHYCb384ygnS5Ju
o7/juN8HAIsbrmRSF6LwmIXWTQ2AOkO2kSZXj696vRdBuzVZnhV/hAGTJwoc6TDw
eLGjUmttJEDY3SDW7jAe+v5pxr1Al4cBfmN+thytQyX16hPddqCdLjjM12bWNRFJ
`protect END_PROTECTED
