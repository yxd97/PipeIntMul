`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0gPMJC7HPBvhnhbSwknXik+JWhO8btQGLsng+2lOqPt7MaXDoDkieU9oJmSLPLol
3VR+0YmVZvVKvYbvP56P93sRpzcplVup9OuP2CJS+GfKahc/GLp9XPfB/tiHYBBE
IlyzpCNL3CJD6zoYfsAx/BMI1w4Y1YP69vlgRz3cJC0wdjdgf8Olg2VxznAK+ZZY
svJIxHywYBDPoBh+wn4TmuHBKtJ7awzInumHZu/EuADnvkkRUbzt8t5k/DVUhqch
4bJipTEn/4JaCy6MLFl9uHamVU9V2RGRoyYktewq1MzBIRUHQDtlFPc6GYXROSMr
e5XyuXq1tDOyy57vYrWk2lKPHwDb6bwU1gZ4gxBhJnSnoqNADjTg2+aR/BmwjRUF
6Aok67EjhpvgT074MiasgU2PuH8dKJM9lomaruTdLPDbuqrAGUbDbRxM3A9VWGSE
LUSlPH9iTESjkpCgAdcxHneDHRMuo9W3KTc/4NUDLDcQ4RU+5D4OGpvf3eKvZjg0
H3qckIrWvmLY2ZGIj2QP5rccXRqOAxZkjTNGankjMjKrJTvSuQwTC7aPIHuuBUsz
Wlbh1knUTctXa+OCIW3GNga0yhhtnRGLeZqHKLGYTCdDCiWN7npDO/61TCLOWUMd
AvoxgfLTxI34O/Lvp/wWFOCg3zHwjJk94i2xqm3+Bua4T2TR6v3j7iWQJH8n1Lti
Q2ZwJwiz2N5M75i8A90yYKPHXtRToicCskPQXh0HbQp+tNRyyPx2HqZul7+UdRz4
U7/zNwOMGbo8rWF3XosPEhw9FcnXDH3HAISwbzgsJ3ll12WFs6qiS9dXBL1/Z2nE
7g1cFo6kH4v8WL37hSr9/G8FFixoh1B9JuxN/BIhyFugKob8LxC1oBLkscmTm+0k
GlzxNP/0ptDmIkw+gRHZGDO9K/F/f8jSewfl+TxJ8vX++lTLthroXO9N+ZHqrzxo
qhU6DcKmpWKFaK8vBvJTibb+sp9CScJj/GtVanP8wJhr3rvlhWUTjN7nnh907gGC
7YqsTMAnQw5Wwjgv7XD+eN0k9xx/cWGRSy0AKsJLGYyyxhnFd495Pf2lFXE4YjWA
99LFMe9cfX3w/ZWe3W+Y74xbNdLdIKfKVJRUe7eqmsbfiU3Qv86ON7TBop9qEysE
zw+fP4cz1bDqHv1bJKH+NltfLFExQMEnMCgTRBJjG0gm0huw1cXP1+qZKXj3hbAj
a/VyZc3ITfF2S2LhcVE3UE/GvImcCnQf5iY+33nlhfQ=
`protect END_PROTECTED
