`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3KuhnSIbd6Wej+RCJoCoievsjVoPJ+BpB/mwbxUdIRoUZ3QZO4Y1E6X83ZBxn1OC
ydiciHwaeFi7HoiaHNi5hvJlDJGOTv15CXP3EQ31Dt0sFhE6oeYQCkgX2UCtJlnn
zELmsCU7rkvYsPM55Y+thjr9W0jtmRTe+MhxJwxLJGyGDhz82iDwOfoEJAnpC+St
ae58gxdh/PbFJZFOZ9S7BEH2NEuX1lsHmU2zobQ1kpF7NMrc9phzQVm2yD4cbSy7
V8t9nauwHxSFkSXGe4WSFiJmgxxhc5VdYgkUfxVBED1EJE7ZTpc6TsbQS7UcN8Nu
VaE2hyeITGuyeXbh6YhoX++m4xn6fztM6zbKnwrydpxpO5Di/bTbHtoyXJPiuRKN
NdIaugNjaHipOgEleZBQyiXwAULJ3+tVx0ts1c5TU14=
`protect END_PROTECTED
