`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I9Q4LpTiEmd69/KCLAEnZ3E0pFojfS9jqzmxm4alniTCQ66GViJGQKYieCu6Ge9d
J07cCgSu+D0eDp14lDg+aX00iYkpMPrB6ZmquNTTNlwdAkJdbNGkJydgMAcpimEi
ZAYRtTmcLacDrDkcCg5UYCGKfBR9AHGHjwFUa6V7Ob6N61UIlGLLp0vcf9FAVnYm
GmgsVSmPqVzEVHQ1JxX/AVvqHAe8OGbgHc8aWZN0VD9dP5U66htrxIKDDGl1Je5S
g6HLIgjYREmOtKtriDS88pzCavRygcSTUvLi3kxdJnBgBz9AiTKs2mcFDRorX22Q
zIfpRuh6YiUhH2yvofh8b7jIHDyUBgYURUb4vHS/pnzffmFodAiuxbNc4Q0sYJvH
rfhY0ZJySc78jd3jzIcs3N3f3C0gBv6HUFJ36QIq6Hkyavfx5+IswyGP3c3+Zjoy
hhI8NjZoHX6M1XuIjjjyE5Yldc88lp8u0D3JE39bM+LUQWOhhi50JBYbe5hyOt5a
RmowLmzHOmqfBoFm6xJHfn1cIKPpXOvCssJr5izF1syz/KgcmvV/C+ZdoHdttKWM
bxa858fdbkIMPVEQt5HZ2U9FVjUEwaJn+IjPTV8dguF9AYMUBia/LoVhqJ00DAWB
3CuKwwL2c3/4chRZgFzZWjUBS4IyUbDSCjjIGS9NP4yi6NqgCSGonWPqqI63O/AW
ds757ioJDuQCqS5FEF7VKcqKML1zl9FRNqxtwCcAkvwEqbnEfPLJGs+1FC5MHBeY
4I3IHcE2UKN5Lkdc7a6g5X1kzc0EqhY4INhU5CjPbrtOMvge869gwz/mIaj4UGf0
P417Xiz/yWpxozAdlhv6Le1uWed5lqg6TNifBixQMF+ggNpjOHAgz5NzP7DOb87s
aebJlmjRUKmrFzidpTzNYE9fsl8UROOYUhY48FnYRBGxhdeo5mdRkJLaxwHoALwc
BRa3QxXr+b4JNkz3a7EUO4N5r7dc26QjTEY29MwNpehs6QiMJDOoofqZZkFlqemC
tVXmJJhJ9OswkjL9fGL61pnxONfovShpqxjchATqMoqGNBPTNTDnpjc0UCM3bIcv
XtDDA1kW27aBvQLjMKzZTVMEjPk0vc/pI0HGIWa7kQZgReHA7iwXImFA2tha1+1e
RHfc1cA3pUjXfncIndgs09QNAarZigMcafQ0Oi6P4hOeoH9IMHc+8DrXu0oT2u8k
4wpV8C06p5t6V6EF/qLUHtpyFhTXPZGmXzNQ8ByKl/0cIBTjk58QmiLkkq5D71NP
tV0w9v9yfHrJY0qNI940qbChc7bgurJTho4kDoOfr+1HOWlM7zjhibsS59vkygwC
mytgxC3yx7FS9rrHDWbWComHE3BVpBY1hn1kNVrtj4wUaD3lJ/UgdV9S/g41XCKQ
DqjoimZmN1zvPqAv0DisGYuJ/SPdMqWngcsnwOyd84kE3bwBdb7TtA1wVknY3Bzz
jGlrBPWmTyNAxAuI3boIX7mCLUm6DISoOLQjeaOB+mqkiql37lVmb4bMmmzKKJS6
gsJgmPcwQ6cFvYe/uVfgK2UdxppecWhSlWxc0yysxNpkucEeutjhJ/LCrlUaswUC
oOICC4El9G357E0ONyFrDnxIkBPmRUpPktq7g7WaELXBnDBSSnw4EMXagyn6m5R2
LH+7LofxHGkUI450wGU/pfAca+3Y/b1oWM2EHNaZ+8mxVAakRakmv+Qcac8KDK95
K5uVE199GcybpyAzhcw3IWLsNwLhs9CaU2Mww1ZDsTGvZ5itiibAr+/mzcLfEzsV
OgZNK7LI6Az9Jx+tKIh6Vl7z/0T5qk+nszHlaSer95xmZI0bL84ENF6pYuZNdtxj
TLeI/ZKgX6XOnEyyINKNkh0A3T1hZaTSL7Ud1gaqtyiVvI4b271JIV8JGD1asvj0
h5NIGsHDfVACyAaiPsrTILIrWz8TDk1v1hrmqzXZMkdg8rC0qaq3ubxzWUojDity
U9bDpK1z8U3LqsaYnqXahg==
`protect END_PROTECTED
