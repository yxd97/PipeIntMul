`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yzFIVteGQhJPGhhqJxNzt3WQna93Ck5GtCQaViA9te/18RqSuZHTAm+xLtBEcO9f
3kEIkv43O0Cu0AuC4v0Ku0BUlqSnY1376gbOyGcefOPoXbE/fZRIsOqT+2ziiwKi
4eVdCrMuJiBHDtZ8v8eGihQh8XKscH4eA7HveMxk2zH5lYYPFsd/1MJw/ZGcWPfO
ryaLBt7R7X4ByiiSEUJNVbHh+rpxZ3L1MerzKSxC5qGXS3f/EyO3i6JVYJ7xGOe5
92dJhOyXSq6sp1c6gY+3tPr6r4f5uA4QkYUGz/qYBbMFg+rP23v/kVoNkdNmsi4A
4D1m9+KMZuIA+SgE8tBUd1Ob87jIl0QtUjqJnJhfTa8jWX6/jTkrl4mOgMjlBEYJ
UaTsVdp4R45M4r2RQHxe42TxUnR7/KoTbNTYQo8FJRI=
`protect END_PROTECTED
