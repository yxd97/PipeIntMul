`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/osxNuz21XMuYar6Ss3JcsX+J9NZ7RXhON40ovomRvmYM5uMJBCUvFFat3FMGBqL
q712gGeFI2XjvFBcmGD0084+/3NXqcmeufDhYfSE5eJFotddB5e2O5zVjOMOCEWf
OuhByvmnvzjI4kGYbQazf4b7Elkx0feuzO78dhLjNIfbaUvotaoj61rElBs3hpRv
v1cprBwMkGrE64cz7H0F8Y1t3j9RmlgyZ1gP83rG8754m+lDYq8ZrzW9RST0G/ib
1nIlHwrIvy0q1J/UlYZ9wlYQbha7Jwyb18FLoW1Pf0L3SOJbZ2ye37/00Phdmfu7
mT9/zqus7NxJCVh6HiattWbixy8xWmfwF8PmLWsIcn6wM0j7M7Rnw6sgUVxAla6a
MUKFmcEPuvbDClW8LYf5oB79/tFIJGEL56iFvzz2azXT6/8bOGmY+nHuVrVnNsjc
jZrste1RPuvcj1ldpk6mrM4kocwS/IjsOa18anC4Aevkj3IscWxivZei00Yul5QK
85HEYZsmSECinp6T8uwRuqEVoR7GqIV+yibmQHzWpwlXNZ+4Tc/mU1vZ/r4Egx8d
r945IC1AXs3yxiMmvZlnd4BXEvNLdkQLf0e9cNxkMew=
`protect END_PROTECTED
