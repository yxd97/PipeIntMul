`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MlwHUPWwjgBCFKrsGuWcjND1iG56NcCVotPe0GjRNlM0Yxsg39ZLNpI8nJK+Va6m
dFUzejM2TTzpdCFc853XtMnRhU7tRWagwrZYz2aaHueFAywsrq2m7xa9LWrr9CgI
5/gbjJKE4L5P8pJZ/XiCLm6TWwqUZyRg+j81qF3pTD9SkVxCrQ2bOd7mfLQRetLr
Vq73bREU6/Adj7Mkj4mpgiXth1CaginPHoT0b4BnPz+QRFvYzXdgXYzrC+z6UaU3
Nn5eBN3lyB3j3+rCI3VTN+u4j73IPoq9BrSn/21VTvWWRx0eW+SlQ5W5TOVDOROd
F9qXF/Equ02hMPgc2/mwY3MYCp1FAR6stA2vFXyZgLQCaVYIAaYW7hxNucjCcS5o
aEl119VJUf9pre7aEcMV6mxAuqACjcIW1ajYiOXXuR4G57KPcZRzWNAofOqst+vl
WMF1Sp3GDWkdLaBLH8NoBjoINXl8PAp2MOPuoBOTRqNRs53Y2kVLkxss1ZQYnB92
GoHHdcAHmiD6vl3WhF2QILj27HMlVsAGi6JpTU7EauWl97XrYIFc3g5Rkpkop+de
9Q7Toe8+9NCktR2X4A7+UhPwfMyaho//Xovx2k/c3Kdwj06iToDcF/q1jI68qIQB
`protect END_PROTECTED
