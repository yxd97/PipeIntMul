`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uAzbDIMPfRr6DJ5cI3LNHFc1gtb57IUb6BQyenavErEK9S2GuUugsYeFuIK0awcN
ctleKL5CtgGsJG8eEJL/Rb3OqSvSdrkA5iwFdBjIMZjuAlSTBeK5clM9TtNPaoHg
Xl6gTkGto401wPFhwE/o6KtEZPXVh4whDbrGWM29BC0cUJGKgEdMk8e/0NIIOT7U
tH89UDGkhQFoiWp9rSkrXVno1UtM+TnWZ6dEZrdTtOVAcC8i66xBneQPh/zebU2M
sjxuVS2qMgsUAkvB1s7b/NPJJK5wje2b1K+/sRZeKM8TCHfC+cJisRrF69HTKuR2
r7gNwCBxO21eqjvPrj6xY2QckiEfoTEIvmmydb67HU/pzuPnVeFe3y4r48WTd3rS
ixFO41BX93yQvxhbGgGujoqHROHU6YGt5vGqycxw8Kvtix9FYiv1ZWrofYYZH5dJ
uE7x0/H0jfwqRMnizpt+gHePZK/3raF9JKvvudAtpwK0JmI6wVyPZR0CHfs9x1Gt
MtZlodziwDc1vznXI86ia9ryxLub/3Io1p2O/ODUQAZR/oz/gLwEOYzdJ1/7TJ5V
NKeny0lhzF/+kGyfKZ6goqXnSZcPi7z0H4mvxi4lOnkgkv4G3WTC+OT5uVh34qbl
IXhwWUIR1qWbVlqDIjkPavBP70ISznnmOaGJ66OATMC25F3KSmSZvEYZDKn/O1uw
R+jzu/0+4Zmd31buBOSZbkUz3la7PJmLC3aBNDJFv/8=
`protect END_PROTECTED
