`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5LDmSqQgYM38W1nk1EW6OwTgHpZElW/ArFLcZVOZHt6foGE8vVp2O6WJ7/z+o8Hf
6F7w448vpkHtL1aTsM3zLh8QGwvlRjbNEBzImW3rBFq0Ra8Ifl+RoVxNIMWtZr8C
nn3T7iWefXVkN4x4KiIAipK216mIt/pcZCDqxyoDw3o0sl+cPcT+QquCQ6sL0Reu
LzvVSKLBlKBScmLCLFFclYauf3QvhIKKa4YnEq0PE/4vsEECLst+pHuPoi6Hf3XZ
B/1uS/ZGpQx70vFYPRIbT80QVuL4Yg2JG/6W9FLnQK1bxuc3czkYRpUFI1XiDAtb
xxOJwYSDQFyHvzL63UovOBd74oxvu958UQB+yP1ZuvhZm6gsnCMK6nwkwx96uoD7
hEgR64eNbAWhWDffkmRXWmqVT1a7cWWdtaOd2ScvkJvaMGh0DHkub1MW7NiBuAe5
`protect END_PROTECTED
