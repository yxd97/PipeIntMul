`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+qFMnyNS7sdOMqQchJe0amGSe01kLXgGTAlvyLZ+k/cF/OFNacWDf+mjVzlqY1dS
M0jKQQ4x5WTb+jGen2XAfR9wudLWCpOn2y6dD/8bmvLQ/iL8wVvqwu7kCeNvLKsz
Iw2sZI1vgVWV6Gw/TrtXsK8aLOb2WHyOg5r6vY8I3QfSy2he1k8ceqFquqtke7c1
NOXj3k7zBjevK82dKcihaLQ23PP7I/RVu8VKWC/jpKOCFtvI7AMY7jg6X01A5aH6
SdQaiRI7wq1/mVUkKY6shnbTuSCGpO2lX5Nqjg1O6w+ceZ1hSOAyLKexon1iEsLj
MKwJ6VVzIVDKqq0zhG161Z/U0GEkPqDWPJ52109AyDh9iDF3Vx18bA841CdC29bc
4q/khKCRAzWwpAUV1sIUgA==
`protect END_PROTECTED
