`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+jBXzQ6lNAsp6ddRIFR1v19lkYVKcrZ+ItY6bc8c1tc07nYab5CWtbnWOMRPw6HO
PJczMKkap8a94lYmqPJCBvBJKdP2YgYsCqFIdSpEzSx66SgLObs0OLKWeK8YjOS1
HybCyrHJyLGO030IRbsj5NBjiAeg66FjSDiZUHHktAoY/DcpGoN8oqOw3cibe6ov
sPb7NDms/Kfidirhr2u9WHoHQSrwHE0xDETJhIXgA6Xeg0ernFSCza0X1G1Msel8
TDmvweH9ABkSG+e/25lDjqdC0mEEeZx5LvegoQMvCUOIdTlCB3ZUa7IJUtKvC4Sx
olZ9Yohxpcgwfo7OvwJAKoVDKz26e0KzCjs3K64ClW4NISkArIPd1yTTTny8oBPn
Oqbk2eGA/tujWRG2vBI5gkeziCMA2t2cVgjJv0YyR8Cjj2G6HAvxv72r/dHfhkwh
y5tAWNiGcwrTgGFVfSA8dYlbW8pWjEQi8vikXnS5nmziX2uOMe7BLzSueVeArz6N
`protect END_PROTECTED
