`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VK2A5ptxlNPB9exmaY96JHBGjseTYCoNLi/H78MnC/1/2aCPcPhgafNE3rLsaW4F
DZlk/lal9Df4ibT56Ugnl/QP3ttvn9QP1jp7tANX/cZxw0wstn/TISvyjuxOb8HL
2UQwIF/XVrdtOwxuXRP3pZpW5aKzO7PXeFuVWupOqV55T51ZmVFfHiA8dTXuW0fA
7x4eU6Va7N6Q7SFbPIDpR40zHDBC6u44xEeh7w1F3K3GW32uEVLxQSLkGeSBZoOw
E+e98WEjT166RLArJleKzu0YIyni5368i5Xkc7J7qFCKq6oWp3zOkcbDgPqK6Gp7
2LkIb9Iy8segetjQkMYwS/3lSXKSJhD6XqMSlALlHZgrBJ9/z+b7qoxvE8TqUama
30n/93jxOtZPBxphegsazTRMO/CWbiB7FFJwgB3mb9fHcq55My3ZmU4xx3sJjK6B
z3KDNjGw61wEwUzR8v3TIpa9vle2YOUnIU9CjSRNpQ5vHnNyuJCMHgTggAnMuPUw
p9F8gTi9Sk7+6rGmkCHstso6q4lIxuim5Z77slqyhKZfnt9lDhXWrGsmQE/QM1BV
Ob7quUkA92nMwIcjtbyC7ITNTyOAMGtcjGQZEzg5MXDOPTuJs6yWSbO8Xm/xy+yD
Y3FdN5Tqw7Ocp3eKzD+oudG+bKCXnCFn6dS4K8PzPoKXJpwQu7JBNdDXSzRBWLA+
HlSpKXFgb/V+eAayTxBIE5y7xroUfIJ7lX2s37DRWEaxbgowY4A0TIJ4+9yzH7eD
O/awE1OsQsxjfUsjxkKF3sx3onklnmhIRw7UA3gMIFmkntmz6j0ax02WGBd5hzBS
7tQPxEYP2ZPuujZXHbndNw==
`protect END_PROTECTED
