`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkIgCfCBHA6yWF19hJdcVvWCEdMT6YEXBo90sB5WCEBmFFs/WUDFQ1V5DCIrVGEB
fhK6H8mj0bzl0Ssp+Es+BjlClkmzfcetim0aS6whLrPEy7M4mTqmIbR4YGc05KGz
L7SoPrYYxDuXH/gMnRHBXZq1XNQLEfOUkdN7S6ZTAjFWNPPxiyvWtE3pnqh2Oq34
aSSnvNwfWB6ozXWpuiF5VnDZhz6p/KmE9wHaTCblAby77jtwntO9tJuTltPcZ8CA
G/mVnVZP4b/4p+A/91/oYa+wjuCkefUWg4KhW2uU1orIvBdJdskQ7XJO0LJo71SD
pagDUkrz8MVt0CVHWQfr/OnWM++fZ3aoeXj7VdQJblEpWg4e8/mgeTGYZqmTw7Qg
`protect END_PROTECTED
