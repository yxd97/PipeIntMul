`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74Qr9yEV/rzjP7lX6r6d3fIfrP6mLH8QGFoaXgsfBdq4lxkduvKV00lKqoUSQGMY
ufPIEPUFdjIjGpsTUGr5QNrdOsZaycCpC+o5/psp3kzeicD4S4Dbk32ApWOLMkYv
m9ltRQSufh3d8Z0rWQZqPjKuKgvETQ7CLiNmQTT37xLhZfholxivhElM4UyDhQKp
G5qio/TswWPal7pt14tt6X/FuQzs9zQxYiy4wx6GLDq0Q5DE9CB/hXFJuAiXPXcb
MlFlV1E8yowX0TYM6ub9VOIAKS6jCsCmpsV81JmOh9XUayBerTCe/uIiq+PDVhkJ
PQ53JiJhImKatnQqRLCChy4ou2tDmV2LNDemwjN7m7JNS4WGKMOKBBpOb27IU0Ux
fGDIEznpBRaL/CiPKl7iMWpIHK8rdKsA+GWzumDFkGNSZVSlx368Kz8XGHBf+2wn
xyMWPa2Cel6vS1YrqTavUsSDohF7NDDY9jAHqYd2P6K16HRvtULnWGndEOL6E8zf
61zyno7ZJa6kmCdyQ/Zqjw==
`protect END_PROTECTED
