`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2MpNv7+bWZaVLSwsT62+APzrA2lts1NzGXpp8V1Ih5nHxDWolh2rP1YQZtsYx40d
ZUq+57gPpexRIUFh8StiwP+0v+emGRaNnkG0JbivKrJpk3HnF+uHhR8okThkfwR7
evv0MTDfxBLdfvrBJ9qP65Pn0Yi08/es8MzpB2WOTPYAUn3cCC+gcGZDQAur+D4q
cWQG/UmlKn/F2ThrLSXK/tWCXlu5BM3+Tj49esafK+/JtvhPHWcB2ET5lB5XXOkH
dkNDVj4jeJrFjdCzIGO9HsGRlfrFbdn46i9ZT5QTM26hcsDp3jvt7Ad2poGWRNpp
OvLcbhuLIReWh9W9xZVEsQXTCeuGWDv2o5cBMm9+8RXPcMtwkbdI6kFYQcYn2/Da
GAIc9SrYpXPgd6u9fIW2CIppLN4wTL/j+Ys7LFGY/s2aP5BOmRAxvN9IeRcXOuOh
6RonJ+GvQSdY5gQwqQVKr0uwHZ0/yWA/wQJ8/zKqgQPHWW0XHPxcPgET/7qtZQb9
`protect END_PROTECTED
