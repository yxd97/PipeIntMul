`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rjUc7cYloB4qg6W2N60cclwmGYJYhYHMgX0mp0RHCnUU0uhOWmXK53F94XPQ253
uyE7h7RWZJ14rqoYc2NZiM7xhQhkFAHLnt/NKKs//hJWZ6Z7nxVJ9DnqO7Bvgje4
szFfssAYdo47y2viVWHoVJerkrQU/g1uInwEPc/EmzRDQNhoUFP7bQJQvn3BBfnZ
87wNudI0Fn08yrl5458lQpOmNweVmp5TB8fT3tlu6f4uCanYQmszaG7R7lSCq3QN
zfrQKHsPeYAeL/nJDvi50SZZGmsuij9yIYyXBrzfZVaHQiQeQWOUUWtf5BT3SZL0
7ygsY32od08ENUCxEQFgZD+aLA1LmixhGD3ctyYGyGP9IdNTPC6zUvP4sXksk1S0
dFoha6R7n42sVKVALLoQeUa87zjBbitYhscOoI5g4v2nWOIT1wneXO2GEjp4hTd2
ZO9ddiKEIZQux1KMPdtvpoQO08654uRYwDto1M6kyaIwyBBPo+UDFbXRZDt8z6Lj
eJYCt8e6Ia4C7R+Vk/C6lNzcSltUYMZtlwdoSHXV0fdU2FwBm0sbLqDHoxMD/xb8
+MM1NHVHhiGwCMF8GWJ/I5pizdZpM2zX6HbHpWaFeVAKHFPpzk9dEt+0VDHLbeXK
Ui4y19uLjv88OTYQQQGD5w==
`protect END_PROTECTED
