`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDchCg4O6arVBhZK04EBDzizXr08fkTcZpgrV/80qw1RqIKiYJCn26Yq9S9UDBrY
jg+lSs1vKnjzWPRrWIPTlNsrZbXG/jTNrClcaCJRwIHw66Gmd2zTjqtjwapf1FWB
CeHggeqOfkEWwt3gFbz7JxrRb8pbdi27nuR/tgolKuDYu4eSvqc9fjVpGHlauUNr
dG5sfdbbegk0h4r4fs/jUPuxa8+56ByyZF35MSgbpfn+vctACIhlOBGIROzlytfA
CZYrXHmz53uQFpR9l2+QDrYg64QcGJacYn+3T7JBpjVq/MAWZzCJXJWIb6MhzGJP
4t2+qZZHJg4fyCvWGTYM3qLRfAG7b9/avVu+OB9OkASQ0mhfznoMj5ly8q4iK8XG
zh7t/Pnosj12RTs7xVgxNFY9yPrsSKNmutwdv7LLwtjg6NW2L99t83DNgQnnXnHQ
MzvSkpeYFETdCJJRSbTMXcLvboxGHCJGAEYyZ/TVFGd4hFnuen/O5q3gsO0e/meC
MrOnwmz/ZgY8KTNc01Bg5zom0KtxOOiHXACYgGkrLrljY78RmenwEmrqV29BhMqS
LDYDzQaq9H0PWbFPPXR3M8fWU0bQirg8Cfdlm2vrQpO3Ef17lr8wtVnZ9PWfQPOH
bHO0LE3gUpXM2itQLd26EPtQ4kbOYhC+QYwgi7Dht+vv+Ey+OJ5vTW8IlqAm1MWN
3ANmrU4PtPvHRT5+ooPkG33n8taVMqfuivtTqgETtohHM9X7alb0RsJj5JrVcRNJ
zo0H6y/0Fskola/mq98qMXxhaM2zp/gWAsK486D4udpjD+/+SJSQMyixBM0xQwXO
zR5/HBgDAN04/kV88jfqRyjTzO/wYJgI2FPJTHu15yZlIIAfkKstJbZUceo9J7So
+zDaPRo64WbYZBPOOWu13BlxHt+ty87+Lxw8sP+8bzWpkQh3uhSsSxGxdiKyMuE7
G4Tv3pfitqoBKVZP1FKIrBTudCbKKNyQlBG2XWM6HYzfNpiQL3T0SacwXM4axZAm
YsjQdcSBNl/40Pb9PQJi0PpB8xsD1mZxaEBGCqxZgpkor/Ra/55YHXOgt13yBvCg
uEvm9CUHIdn3sSSO0XmRBFfG/kvE0amzfYaT3KdadT01zohQPkPWkgpYJAYTrvvp
BNSlz4H0NYUGn420IT0yWooen6x/v+pALPIF5X0Llujlw7QDCNlciI1iKYkrM++h
Ij7VNPDa3bDgdCduDb2AKCFPtfTPIY7fwH991sOIQ/xriK3uoRG/aGS8kQXPEv1T
Cr2YIyN6JixYQG71zjcpkpkrfWo6AXqk5Whp71NwK7RknSeJa2F+MBPrc7b026d4
cK59tzq5s7k3U3xllvCdxRi72sFFgiuFQC4UOY91J08aeZvx3PGs3ZIYihJBgZ6n
YyH6FjFmbgwiNLzF3edAdPl7EeVlkZBC9KbhFdmth+nNSKqi0f74BBUuFjTh6cbj
3SZrJygNA22660JzY6v6QOaXV2piBQWS7XKD+fkm+wHTp/9OJwfzOQ55S2+Z8S8F
jwVTwotBRGdwStE26F1oBSYoYI9KkB6iaNsqg1LT/6S33LfiRVobUgdGgod9Ot72
`protect END_PROTECTED
