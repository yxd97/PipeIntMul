`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wJ/zm0XQkfZimPNxCUEG8OzRBvjEfLiNR5SCVd9XtD3V4yKJ4sTvfGo9xw7yLwwh
xFal8iei9JbSON7HfXEfODcXSYskpNG6lFJ1bX7HKEMQ505mb4JwKi71tIug3XYL
Q6LIkzLE5CJyGHruGIfzbsVx0RCZ0oB78j8QFU30gPGRNpOcR92fO5NGUKPGWsih
kEqDm+XMaMAuiTgSETN84X3MGo6iMmjwBe7ZL8F5fU6jo6MPOgYFS4ZEvQOg4/9N
7AK2E24ud7V9LxRZM7IpLKi5smhIHbd3hTWRV4ib7CFbSXeCHJrwjIC+UBp+uCR9
H5f/MJQBfPqUQsgins647Bhj2HBkeh6LyHcr96a9D9Lk6cpmU2h3qV2MPBT/BEKC
15DYRKYTIJCAtMwKhgMuGWiVEFSwjrC/SwhSKkVQR26VKGhdURzEYkXIuSv0c2H0
UuH70h8ecoc0o9z/P57d+qMQ8hIHHkUEywBnm9ciJO786x3m1WHf44BzOXXq6Qwy
Aj6hYHrSDswN9EWUNdVJtcLk8tpitjCQmx/Ltx6dXWpURrehL6Is3KPVqZ6zX49t
tgSRGVPcKqKW0CV4rj4e9mFc4UPY91C4hzQIh5Auom6/Vdfzb/vbeemS6GFxzW4b
6MGUY/VuGA1x4Dd8AL3VjALddCB0cNImNt1HqSywQbcLJQFpKpxd1LVecaKqRqAQ
6kPviaGRSQQ9wxtv1iGRZjF2H4K/2yrEHTqstzye6TCpkwXvFGmHWwZ0Wv+1Mp8m
DYnVrOp3yvwdAp/PAaM94DyjF3MCyBF8YcujQ0HUMC59zfARGvFizxEmls6+H7kG
dhWlNk6nlWrn9x/IOm9ruQ==
`protect END_PROTECTED
