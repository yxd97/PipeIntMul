`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d//wo7sn/uJ60D9MM397Ysx8h20roPX5nIuNcKh52gTmAVb29O7Kx3Fwesa1x6Tu
5hq2tizX4c+hHeLtMKMcJ6iUtXHrPV3ElCkYGL7zEV/PvrbOKpF6vmqaJRJwLtVU
sCbj5E+n3B8m4Q0SZz7cJlndnICDOv69mC+k7XLsuXTmCgGjwwAG/roZwtOryGUe
N2LyZCpnDwoadSUJklTLgjRrXqfIqxsihIogqrTkGOz3ghJ79xy3m4gzC/FH7AVE
8TuNRfDh0eZojE5sAn5tj7+TR3uhjj7uvZMVSESi8bil20j+oTwbM4PnF0tpQmCt
xH51ifqhid1JSORlbzRaFRFRxLon4bicusqD038+dSPrOIHgMYs2yAU+KNE5kaSY
bq9ixE1JliUUax4OyqgNba2gvsiuzreFLLQg2+fRnoCv9Hq3iUvSRtceUV+rVT5d
gccZiAsiRoLTFhGSYWpJUPgcbG4UJyG1EgmG403H7VFtxbI8zv2RnbwLyjo1KbQ6
DWWP74HU7x1GD8xIk6hfjUMUOFnNyQ0Zi3U3CZPFbkmP5Qtp1kAhohkCbe3Q6l5v
lm8oBnLbnTNyOdx3T6Pr3+WKze1eZAUDJocwgDSRAbPJcQO+leh3JQhNGtVuKvgS
UgDWgoxiVKCtdSAzMkTz9Hf7BYhurm1H0Xaxala8Hgpht34Xh1ixYIx93PzUMAgO
fQvTFaCnONvtDd24plAnvTIeJJwQg1Z14wn6+IecJtoIANxnYE7eKbImt1X1h1Lz
wwDgGcM1yYAR+k0REpz7/A==
`protect END_PROTECTED
