`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GYuzGOVBjQyvWbogJX3U48nghJeyrXSq3yhcXao2BXOmvn4U7QhrGPDPIiiJ4xQq
9gU1wL7/pSnLKBHBDMHvMhv8mH+d11K5nszdS3pAQZvPbl+kK/dGKQzCAILKAqqX
osaGCP7a0xt/5Y7gOBOkl7ExzfWIA6jV3tG+FIhjJ9c3gTWYLkradjOo4BhwVuQx
BoZY6Ciqcz3OrK1L1Jz8kqvOwlN3+bCCmdh5q1Bro+kDYsMYGhRCzN1x0hnIUsNa
9sogOGFAc0wESBnWkxM4HTGYsLi3UewK1hikeJcwW8e3WctPNEq+qWYT/zrCpz/e
W7HOdceTCiLA0x9E+BZ1HPXCuHdcLRCTYtQ5S7j6zGst2boYtd6KfIBPbpsHbot3
4X1F9Ra2m56o/mC4X1nOjwfgl2jNgecLeY5d37xki9EMMBxtKU2i2FSw+OeJmnzh
LI70hwSgopPgxZS5fq8DMdTauxslQZu+1o5UZgH38qLb/XpxMLHmp/eY9CF5nkXr
TdMtO2zu588jgVdP3LMm9ybrfgdUxQPV5Yct+MsprxP/hpnSbjdqjueF0z4IMdur
sQxMkuLzXJFl5904rpACf8m6zRmfX8EggdiJAJGeXnrE8KoaqtF27NsMsvDg+mo6
/Lz7nXhW6SZt5l3qBd9iHw==
`protect END_PROTECTED
