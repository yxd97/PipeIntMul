`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UIpE/nYiUt6YDCY0D5gEc8y9UFXmL/6ryrnKk9TaDNDhNizsII8UpJM1M62fij4v
/mVcOnAr+h5Q98I+15XU0LiJnLGeFq/cdOqvo30/Ki2iZ6TlW3yQ7339vaIlyVah
CNu2UIXXUrNJ8KGqD7SDq795/X2YYCl1p94f2zgq0d43SLSg35sGhxiEarwuKHpD
Jv8b17SM+XKN9r0TrJ/9tLw7InzqR7oHvCVkE7IcDHQFDYJ6a947cjHwzMR9utX/
O+i/CRtANa/W9MrYQx5km76VV3f6jP9MQHSFl9cb5j4g7y/lJiqdmLyHFoEZ+AF9
b6diHcN6g3ql1+YJH7nDLEjTy4LNYEdjyqPC/7hDRLq5AcXbe3PTCKT0XeykRZMJ
3knnshx6gjkhKTHctCh7CbyWv4/wjcuLPbGLXioluGa48v0m2VaUVucIY73XeSY+
s3U+NPSWckkrCpSLmKgv/qFhSJBLFEM3OXRfTz26xlhfJj4m33OlLE9l/mMu7p6j
P3jpJmG/Cq5ruufy3q18I0JE9AuzFHthkBiEF+jUi7nz3lZFd6E7inxyTH7jWCaO
K1qPsMi5D6XHuEaYUcp7TFHNY0yoXmpEfVKiaB1y0lwrOORGNASPrrAhRvNxgJOX
56heOknazlAKk4y7QKzqPBNSc6ufS/zc3Kn7yl1NRhuyBCvdSDE8/JJK2aIUF4NS
rmYbgXK66ckp/MzQ9DW7il/hTEGOHFwbO3/tHu9W1J+Ey4HengT4B2QuhnabywZb
RBPU7l1WFk/SLb+jdiokSPjuxznBelnqeQi9/H0QqFZM3fZwJRCfgf7cLKHndTBc
r2ToZ/wfMK3YsphbIhYa+KUJU5foWj34kg3uiykWu39HEAFa14IkvJhnO+B5Nxt6
zOilRS98XU1uTklf53XUZy0PasFKOMCcXFFNbC4Ks24wQD0f6DiH0+FYvgxmB1ZN
ZmMQSYLSwQDwz5LZcmbe6djUvH423dvIOImUZgSlrVpUleTZT0vOpR6H33f3k1mK
lA622ELrqk14SgJdX+QAaRa5FZwiyv1ov1OniBfW8T8a0IXbV4uyh8NIc/AN76K9
gfJVFSBhh8FPwGC42Xx+n2ycMTIBTgr1L3NV+2/TbH7iD4TGvE3mk6lT3z3TePFb
caDOW0YzZrEiN2Ghqm51O++erEV6YzUxAk98/1GgUJzmhq5+rzd6sIyeECsLW8kB
koAykK96Nvzr9qRJmMHm8mFavBaHH79JRAH3dRaG/N4F7OT1bZzu6WAWE6miOg44
KdVIcLYAIdb9jZmPP7TsO8lNePQBh3rrO7CFo9/ec2HExJ861vruDE7FqZNu7KAm
tXkLG1eayysn+mCtOz3AdWDemmXR0fwV4dey+FpTfL2wmFHnMiALIfIzoLhNZABL
q104FQgEzzCKp72ohJrWI8Y8brXUV4pGkiUQA/mwhOavcoaudRaQgmxaoDedRmck
run7Ecfx0KLisIVk/2gWdTNSCJOuZHUSmvdS7/ACKw4oLKoaSNwaeu9XW3MJuI0/
Iyk7pBY0ZilWpRsFE6wOtDZNJFgfm267NyyZNeoRc4ZDV5xqwS/+0y6TJ5Yaf4WV
znAzHOe21Am1P+lsyGZcMgh6KrBDWb5jeiw4aeWsP/ghm+kZ4NRiNxT6wk3gGa3P
Qr3FGKwTJEUVBMUl8P9A6dG62byExNdH8pO8h59KlU+5LCPKXkPnE7vHK3OnRtb7
bYB7peJoxrTLjrEOuR4vsM31woB3XtBPOf2WgQO54o9FQNIsBt8hGxAVZjIrMepP
ojwU12wzUCBzHHF8iXHhKrxrf2EZhGCrYmGrmareTgz6VBRs7MjDgDz6tERYD7++
7hgGVLnXbBEv34PBaM3sVuDm3MkYO7ZIaGOGqVo7RFrONAIXfs8785O3giwa1rGk
mV0LnNE3vIKUUcBzpSK+f0waNW//kJSnrgiMxfgDvcfQqXCTusq43l4f6V4WMwTh
395nZ2TiXJKnU6GUNcsS7sEMiDSN198aZHwW+r4ZZmX4IX803DSRO09cyl1PFLqo
erGGRPyomSHKeG1qdsxWmNGZlJ/c/zvo9kk78pvI6yOlqAlQvNB5hwp8G12HxliV
4tLdeQfTpc60FZSUS6B4Q6u4OavWFEdc6MEb7bsuQgrhQbbyH86lp0I88j4bmEm1
KkA11pukRIFEKdhSAiAYo9vclGyqOGgTXk2+0qbxtTOSI0NCKHGDzxXRwphtIz8L
NzqQfh/YK9tSr3jlBNSbhWZ8bkyzBrL057seT7jgSmxnmL3JGsoldISP528HwVaU
kXZtGL0GSQsZWtD5PGdY3H7csf0jFoWHFtJp3lERz0BUmPgYFAgOBbFbfNRaxs2e
rPGbNkKY0q81Ss4Am6OkTS/5Fj1Hz0AV676f789aAJjcBkVHt0pmcJiRRqedR9ar
OzHMd76tBSdeDStC/pYCmUmg7l/HzOz3WEnbd68OTz9V2PTnU20tFLQvcj5e8QPj
iZeW+abc9FI/JiUV7jAKkkCTRX1nc/0B4+wtqWO9IlpHWw842kzChBSCLc0t5mL4
geqJyAiT8VgRkdnznSY08EkbOSwgQBxeiNEFwGpa1jLsxYKBl3O+SiuE9ui686NN
buJkULwpReXHgLsKSbOPmpaAEz4bP5rujRdPWPURMLyZ2hW4pMcqmPS3V6Xcf1QY
0VJKDUJYtMoAoi3oIsCsYgiJHcxx3TrUMZirU2NbLmbKtIdcd8PaMxKLaQ+uO0KE
ebqk6KitTKT0TqsmfIKJdcZoUlHmjN1peRb+5IP1NdWYpbyf0ZRkbWzZTl+OsAqf
H3oRknhzY88u9ZEQ0aUkkfODmOdXFnZ3RmAGd0cKwNviXLhPXymC7AzawQCwfVAW
y7F5Rwu7gzLL1Dviob5f7vhMmSLIJHC2KMuwrARDmERHG0n1Nt0Vr+NPLFdXJubZ
fKsaSmoTjrEGshP+yW/iiV9ewbemx5c2RnRKoK8jJtUsCA+HxBSDdDFMHd1zxiLy
UuNJn8ydgy9jFLRWvtYki3Fh3h0ivcXnpgZZMO+T6Lg1MaJ8ua36wlvlPLl1gnD2
7Igx9sXLMZIMqSpIpBszRPIob88gps8MM8VEi2UkwCXzHKJdVcxX8kLYp7AwlvGV
9Harl1QMQHDmB+0KexZFHvHH8nglGedLOk6UOnZW6fvEoI+pvJQduKPnd1+sezZC
aeR4f7DIKCmnh9OPjEgP4IWjbU+WUu83cI1GCxgnim4crSdh848hYBDi37DuS9fw
NDNp5PvjlBIp84/HHldc5luDgysJxfa1YYDAiafLbVU9oRkhCxa7x4jlm90mOnu0
8tTT9u7KKXU49SvspLEjOfmuqdmszVfYsugIue4b0PR2SlfcrVts0aknNMsFyCgh
EMz4/uWcUeD48Zuu2csJpGgL+yY+woLT63KXCcczE11MQ0WCyBjQvN7Dc8oc89Sn
qSAAiU1SUFE6egh2pNPaC38OLHbE3ZX91cTGkkIhF+mSQMHIbyZUtDfLKrTxbqqj
55wx2dBx3vlhZ8eYN263OoizTvxp5tHI1dVHGkqr9/Saxt4Vm6fW5b0KDIn4O8Ej
SlIRlew2pKYqtWfDF5k/iwhSu5GkhJrse9YE7psi/qSuKg9bRYwnN6oGUFx8B/QY
nSmURf5SzXdlQDCjCexSZWShmxqzHNC/LiuQf6lRccar+XoOB0WgjOY2GoqZol7g
GU12eUO2JURZIKEefrx9FgtJcH3BTBN0HzreVCUZT/b2Z+joUqZ5mc9+sC6802c8
HTBJg2n8tMbYHNOTw4kz6cZ4L8T/XGQgeX9naxeYHVd7zGUnUPAgI8ysTiTetVEP
mUo5nnpZ9L/N44SBQ3gUDaJmQ0V5JA0NSkms7H5TqRHamPL88I+irJsZohDcghcZ
vcx+W0/ZaWEvn2hk88wA3IofIahaOSucvqH22Pv6O21t4nwpwXRksUrfhKVpoggJ
9BOEIDcsD4BgNWtbni/QxXVt5/Q3MI6kRZ5nAfarzxKrMAamv9KdPcMyB2QlZLHw
WnLil6YDzbmYzGp5N9Wem7AJqZAS/yq9GNNKjEbp13ObocTWS3QnCao61b1xlVm7
pmt/7esrdnar0yW3np6pLN3bjajNomp7KooNtGK4RU4r5rv5eGOGXM45XDfSn7lB
D7sLQYMHRgJjYq3Th5SxB+sxsDVWKBeIkkkiN5tbOr3sCGxBQevooTzk4bayirjW
VUF61IDioMxNzjH00SJA/lvEge+qCi1r1neTPRqsOGNkDouok8j7rdlaSrAR3fzh
I1tR5qPYGF/otHFkzz/gLK5ACzbtkukwEab8yozWeerBpkN3/Wv/BySU7CNNuiwB
Xnejs21t3SIfPkuQosMF3uXJ9XWoQLD/NugKoqHlk0IuC92KRxEGI0zJvBGrfWTX
c4Vil/DLI51KlTFxzvYNx2lE6qS8oLZq2p8rRkyEQjE6tDozD90PyFEYx7AZaX3L
PiIjL6TnjTMloaVxSwfqekUqF0aaTFYozgstzLOJQ4EKy17ZW6WcZf20EEtim2jb
+0qghtcuws4y19oJFgAbM+WmST0Bpd/ZXdyvct0LET535AW8usdDlHQBaaEq9UQH
FDpGEDthX304hjRgXytd26SDmfj/PNg1nxbO9PbS1Sjdh82L1OfUcYNBknc25Xke
u5uNbdfDkwvHmHOZltG9Api5M6ujQ1DNP8PELw8j2LNrfNHOoPjiGknt7y0Na8CV
1Q9z3v6ia+n6D0Uyyossf66ts75VMwhnNqQZ/KXWItrd5R81W81gudDCdbAFmR+K
BxlevsZli2NcW1I+/KpQY+OLl9VjnONbyW+/OC8vVoky9R54E5SFuLTsKJN9iIUu
UVnZhBIGHs0qelJ85FOQx9Jkf0tVwONgnpfMxiL6AyP0wUAPiMTDjud/x+eVqs+C
aBIiXXgWLm6Jvkb+Hj0VoUAZGpeFImIqtqnmPHY4t0NLcEElyyxArvalHZY8oo5z
lABTPup4NbHeDL65AF1BeQ0V5ajjeGtOh67fjDUrpsxlwB1GFP2VNC3ZmKkU6QYY
w+qDQ1h2x3uz9g+9y23dVjv2o6Up2tsadCMwcIqGct+DUXuHxGlwWL/GlgA+K4MV
Jy9AE9FvGYLg2RP7qrJZzci3lduytInfat+OVk+qRYdbLsNWFLYHUQVTBK4HP0dj
bvw85ASLeIAzQKHO24y0V9c1auI8f5m38KtT5ZX7EnwjgCScrzqFgewDWBoo7Aha
DUgFcezC2wZB4EzKbqhOd7YKCdJhR8qK9xog9oPHIdpRAk6ZlPrCqCQHSky+1Y4V
qTzxRVWAI9zbKupfB0Ly3DkQcpJjv/jtmAvd30MV5kDVswVZquFTsefKSiI/rpsY
ePbTU1eakVx+j4R+Xn/wHXmmHzCedUI0jJwaGHFhmIA9j1QCdZg9n6/1tK6wR3oK
y7JCMBWFlGXuV8YGrz3nAX3HyTXZYlvRGpLIMWcGwSVK5gSYdthaYR4tgDCVCvEu
YWQTLOC37Zv3KtrHrm5/YYGQFQdpZXAz5pqicxbssnSjBy6UY5okueZS+otq7QAE
ZgzCfjocM4RepSsaYwcaQQVTxv7lrT++E7xY8PeClaXIhxkG2PgoH0IXaSquBtiK
n3ZyKEVaxxRp9lh3ROGnIvLSC0f9MNdi5vYVnMEoYA5uLyDtbGnIvUVmX3Y4epWD
aSsUhOvQ2JLdNdQWa4n9QeDNYfakRRCG0m4+4m8kzx4PsKHl1ytAvzUyzDIsGCgp
c6cReZNLyWxXdFDS9Aze8JLYNqMsNlMYs4nFg5Xz/NEZAgn6mbZ1P7u80xNV7bDE
M2cyzm6bQlezF5H4S8DeemYCh7F6uoZ1bRR/3aaBZ+K705wk/BPYiaK/gBma4B8U
ptXunrlwgTKmY428Eco1nGfn5WIbCGX7t4twKepZrbn3CDqFKAaic8w8TUkTgVLj
hO2a2N6Mm9mwZbOZD7YB0uNyWkU/sFPD47wPeDdwji1Zv9jNOzHPsGNBaTe/7pwy
lbRFBnwzUpczzR/2/8MSxYgKdjL6oXP/p2YtqAEtwfLkEoK8dugEG6j9nIwU2xk8
aeRF6Hk/OUSr6I145JLAKXckBo9+T+KqDrfLhBLf67tasjksO5HKTf561m4Eqpk+
SYIRPaMb7wxjsk8NU5SauMNEteEWT97sS7qNl/IuadIRJ7gwmaEzL3LJIoXtscRP
mWQ6c2du1IzR+wEbK8kOEUh3vSBPA9VQUw6Ddjk2zcHjwKbj7JDXzSoOL37p+K+F
J3iKzpg2+j7nXGayxUvla4YYjf0rI9UoFLhDPdvO9+2AVrrxAzrEaB+7HME12rzT
3JW2VMt/nrxtRBYhsZnijzf6hb9nJrzcR1fgxEuTvMZgHTT4whBwk+Ka8f9n+oOh
gBGMvM9UQHnQLdlzmWgIreon1n3czKxG9jUaW/ZRRtpArvd/0HYGLf7alkqm3/Sn
sbZO0KzTXOudmipZQEujVdJ2iolK8QTc58hFowab8lsPEk47Kqnn7mKPFOc/6STd
mE17SBUzXrPfmyDo35J3fyglSE4zOZ3jw6k61zZokEgGyls+1yq2aCMZl810HyBC
5ZRnQ7kVq2b/xJl7i59SkaKYGWDrWq3YvkGvrgqH7J3OqkD+9Vr4RhU+BZ6102FI
6NHIhQPG++lck2KtFJRTAG7D/C8yyUWtEYD2/jo4G7SkCY9CUztojdRk4fiL+ZPC
gwK5TS7d/eZzS5bChtwPsMbCjniDs2lX8u7+Z4N/wZK+x2ojCdqVV6o2a34NDLL0
8GHuZ+D19qkpkyQvUnbOO8mv2ylh7/FFZStI18YB13S68q0K7sUtDBYgXXODdeyh
mIBQAWK9W5OopyXahdQk85wDBhHSNTZfk4yYkZoy8znwrav612HWTioebZUw+HQB
+ut859n7jEhH8tWNcGhuO5g+ontCPz02b9dxTpwgXRwsS+PLoq414WKNVf1xXO5p
r+PgR2QQZUmuBShvmNHLSKenxiQL3RK3moHoNcKbqyPVAVuvJk0gZlR23tI/KlbM
qxvjknK7qAG8HGP5FvLtj1+jCYsYzZjLnEXsSb5Izjzx1F/2l6KaUBlaDtmKOfLc
mhzeU+B5moa+3B7T0VK6oHRze1xWgLWyjUEBvpBGAn3tj4bKIVvDRzZovGYbbJXc
vFy+MUxcswer/CUzCpgjxJWsAZ/nO85xzZ9FPU8ptgr33Vm48rMWYzlHytnJItqq
QaLbvoY8rN8/nKVH8VtndFqZcqYw+1W4HlJkcHIHFtPxlSoMlAlwFX4yX0uGI2D/
vghbuRsEhlEayZtlkiPiHfmmEKixp59sDkT5FNpLjVQR3imGUE4/c2DVGzjoYuZI
xJRPg2Y+YQJkiyXER+wcNE1f3vbDzaFR2iHuWXR2lAyhQ8qiask7oWiIqjgc4L0Z
7yrhGiEt6drSbtL0IRv2xe425aX9Dq3O3NlrUzl2gCILYplxtdZs5syF6nEN7vUE
aW3Ca1+3/NucRi9gpbNeCV5pNpo4QFAv5p5xKd27JeaGo3rx3DWFwvjlMl7e03IV
bVH7WQUZlfcVW21ew6kkxtcjUT2IZBM7HbOOWVSqvxUTMFxYwwW6YURwt04J50X+
om4eCTjMu4pojopsfUxa9lRkrou6qclLvVV+bqZX4oI9NZY75iImw9wr+cRaaMTH
+9F5ampK7bSEjiSbl/Ckj7Er3FqoIJj9NE8WLB43SzcJu/c1snIGYsrFf2vhN3Nq
tJgsB9y5niBkQl/ih/9RgYlK7Ng9ABq2/4spZYVAa+t56UL3O4qKQzpS6V+9vrSL
l4AbtYFlHl3TpsfccvFl0JFK5fffgHAMQnDaU9Ej/eU3jZyQiWm/tWTmk4TIOvFT
nIPE3PZWY+1cpUTGZ1lI81Yf5PfRnCFR9/ZBdxUZn/UVzb21uiZ7SiH9ZzBbUK/t
WcHIvWY7bhvtJGJVHBXysNxCKx0Tt+hfG2a6st+60lLsSWMj72YU6j4+ag7YvUfh
Shnqeg1ZYQgLxfe3Cuy47gjh77fn2ZJTufKMZ4vnTmUCYhzhJrCKvEgce0K7ktO3
MBQLk9hAzO7msMJ8KEdjAzvU4qYUw8ROwGbROwc9eSo=
`protect END_PROTECTED
