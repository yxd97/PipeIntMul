`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59Uq0wMnHaGvlex+DuHQhfxv+H14cV6ZKUjjiWpOY7rc7jP2sUYAxuhQqO0GwvG+
gJUiAF8h66mmj6KxzjDiZk+8qHAuwFl+ngIbd3KWr+5/CCeHzhdrDzagReO0Jmcy
xvXRuzR/c04XYZTHh0wOSDWD3Y+xzXA6JaI3SIzgvTncl8ZuCROnohcGri/RqyG6
M5RbS9CofurCKgCC0vGfB6RdDW6w4P9ridZkiW1z2oVZ0WGgixROLYR9Q/JlY2Zb
xh+Co3d4aQ0VTMSp4oGwbNKKfujfQpm/Tvg4aZZdIHA=
`protect END_PROTECTED
