`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+aCvljyp0DsNIB3EBoHII59/Lqdt+RiAN6iUKiuaOGPVAyEjg1Ii2ERzYKCmc2W
GP++GBioQh8Z4jxYSNM5wVVRQ87YXCNxtAunDCG9pMjH7Dsh155fRdecvvkwRQuG
Kc96IVoLIgQ9bMYHPjzgTk8z44u6jXQF91Ke+8DVmfmr4GRaNKU0Tg33mQsRcdq+
IOpLRPy9CL6IOhDvSlLOXHQXWvKhoxurKzihXgxR2ENt2xlLsiLsL9pBLYatz2RU
RH+AFdA/rXi25b+Ci2JSg/hC3F1YttrQ1e8q/zCaLTaXK76oOXMf5HrqUczujZN0
daSm6V7QTso2iRFpzqMen/YxlpamQC0l8wcLWAFZdXdJ+MtRxNzC6SBk6R9gdez2
O/n3KpHgaKPEPjTwPskFpc0wa1M55lRHehOMhqUmtHS2I+Tu2QK7pRlSNb7C/raQ
UQ+l8O9fQN3gBlm8djEaPrwYlPeuye+kxgkJ2LLopBe65Dd1q2mW5+zo9bIIfFch
uulb9cyQtF1T22qFtU/rMB3EizhsYccHG4go2p2Of+vSaM/ajIKmS6jwbAYhlKwS
Kx3U/VFEkjqP0XC1gM+OTaj2gFa/uj/W4ucAVluiMrVWJBtlPfTPF2WaUXj/6t+h
d3kE73BauGo4xAf8500Q0adGt8HNE3PChBZVCNv0FEdWIjC1rDV94SpNNP+iFTdh
MZK1qm9Da9BLGQn5dzl1c1+NfY8WUSfUKXaynjqYVx7fEBVNers+nHB4AAGU20IB
m64krsGDmjhpkyKhFe4f7KBNaMGzp1JRPsgabut8j86bwOslMYNY8cBTOoWMU/Si
GWYTSWV8Gki5/sdHkjJGxPmuq1PapsEdlsu+VTQkICVJAiZ9Hhd65QkiK8B77ETs
EhvLXtqBQIKqWdxKQC9NaVMAOX4LEKp9M7kpa5qlVvuWNTTeUYRxmyiI6ysS0+QO
1zgZjG8zhspcM5N9K+xeV3d/1PZw731yUEA58W6PgD8CkzI0fWQJ793TyUuVuUKd
RloMXqzrqrVnEQMOUd33Kvb1+R/swLXr58qo82q48zG3jRwo2BKmaVeXWjVdA+Gj
eyOWOOl3dA55JwtjUAMAgZeO+tWFWcaQ2q46diUE4sjI74k9EkZ70VyllG7fsR2j
HPOZ+BOeI4ktwpeytRRUdvEXoYQxd/aI3wMH5blNr6+zjkYxJsEK398ikzqWQRD7
y48CUKAjXd7kCK2cRNnMCwHb/HMgqrvdO8dgyy5VgC9Pju0YUzPWj5QR+CCv+PTp
Vn418qJaGXN2TyhSTZu/fte1e+NcJkBRmLp3Tv/gqvx9FVB//bW5pDESCD+RE0AI
Qygli5sy8suJLSwVldgGIUP+FY0eqCRVKYjMUHlr82dZTpQJ2uC/3lHrTNA3YpXw
sMDJP/yvJLXFZQduUTSJ3hXw9RZ8PRr/9dRQODs4/pWXLfuVgYqDhvAx4YKP5zJ/
NcShz/ZUJ65SUL1PsrVhnWsMSp7Z4hhs0fBHiK1wY+2zPN0aT5n2dNk0bQIjBIXO
1dJQ9eO0Tp4mQUfVLCjps5KZ/lUOBJwHNUOJt1ezeedN4deFFUTaYzWvprE2I9du
mqd19j2UEw2IRM0XvuVmRDWgN7zkeh0MbgroB4ff0eyt5lwQBxH8dfG85A9a+r1j
/T+zKJ8wTrftOcln6URuJnDAwyPZhbj2/N8ARa0ZRTGWdktWN4NH53Zh26AuWIR8
W7D/1Vuo5aGGJeGIpMYlgZfWWyBCHbVUtiJOgv6cEX3VZXcxrWDugAlWyuFCViE5
uUgkuE2twMH5UnSEM9dbETlZACmOqU/ca+30L8R5KCTb6cfgjgdbWqIwdPaDYEaP
n9cIbmDTLWQUGfwvsvtX2/mBH8TEBJ34UaHU3UHEmqwGJ9eR6Fr+pB7qWc9QtpSA
X3ZFWcKZJ19lNxFhZwIA+qPDOxZMQaIEx2wcSnvcM7q6VHS4cV6Bk+KhnLo0sn8T
9JK2mOHevIdoSteIEy1kdOJPBbREKFlWEp/NpRnn4vL0b3EsgF6pCVsWiEy3acgE
qO7XMS4Tth+9CuqK3dbMh8r7CP5xAIvwyQkXZ3kC69u45L8DACNLD6S08vjuOMq1
6g1oWLk8Vd/Q4qssr+DjiAwI/sxOrbPML4RWk5f1NFpWdF4crdWaX0pj2/1HGb/N
GRNzl94ygZfstVjpvxskqnEsoGRL0uKNqiPkeyVv2acUvhVfO9ffOUkQPR/JBlX7
4l/8ayH1kUfEdumNAz/sNv3wV0pYSgWzbpKmvEjoV90=
`protect END_PROTECTED
