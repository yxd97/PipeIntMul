`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nyWnJJDQrEVczIqZrjSX5DZOjS7mq4mY+YHJV6foIOowl4z5+7bcmgUXglF4Kmb1
MBWrzwbCmInn3lNXip+LIifS+6yQYZ01QZyKmEMzzJM5J7KaPhsrVTxS0DtZcVNz
5QwBzlZ55q4xFfEBsUhyyYa7CTFyNZxSJWJbSUR8MKUhMth2TGu2oelJiVjmTi4w
5DNMnzGCKFzieVAZ7vfJQ4y77Ec1fVUI7PNALI8AX3sJNsfqWGntgOCngAWyMgMK
I/zZGWmez3TiREe2PYZQNlFC8DZW5i/FFsXGCqrS7QFY0WD3SVLrfNKeE1+XEClD
xxeb8+al8h3uJ/AxnCiY8sSUuI5MkGuv4S05L5THj5e6BYE5QI4Z56HPQY5L/249
yC0cfCCdXQRWlTu1QFuJ0r63z94t2bfEe/HOQuj+y0vahuIjteWZ10LMHcKLOp83
YsD/Kb7DVKFv4HGIdzox8tSnt9msk9BsWRPPlogL756HEAWznwpyZJdJ8n7kogqv
LhsPsrRl+jKy/iasOISfUw==
`protect END_PROTECTED
