`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ow6vPQSfU3UG+AwDDppHu12B3M5u/dBDp+i7oXIMhKXAemGvhaK7mwKSm9ClHXJA
LFP4kmR6Eg8nOuZyrwAv3dt4CHCEs/ZMa+/a/OEEUDL4OAQOJg5PHSPnstaFIHu4
6JXEe/A3CqW7P+r1zhqtwYRbjtyN1LYsowl9KQGYEP2LFsJsKG9TWjMvOfVyA8Ri
OsbRpJ7aluooJyRKUtYeMYy/l5We0wDqX4NTp8+IrLAffJp459GmWcrnB2BgfqCk
`protect END_PROTECTED
