`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URlQUDBW3hFi/0y0RkxjhKmGCx9RHDnE2b/dL1FSFCCbIZaFPp3TTjzp+0FDVyIk
t0/IIWIK0TWgp8f4Jd/oc2G6SfqmOFouDHLO3Zpg2/jj5Te6BBINWXD4nwyxb2+A
O/Pf9zsniphNdx9qyR+eZ0iNMII34RVIPfwuIOJ/jJwvdqt+yAckYKg0DkL895tL
FUUfDW/Svp7HihY40TDNz8rWbgS/IxkIYrJJ+L168QQD3DwP9IOs2tSRolCyJl9h
Dm7+2xRKy3MD/bunDMa9s6wJB2OCRRvJrluBU61TJml4Zq3Ot+ctoeSQ1Pc65mfG
N5ZOqkWEOeV59Cp22n1seoneL9VP4iqNoN8Qyxt5ScPQrp/sGz6wACC0oAsrnpan
4mjE9a6C6jX+aR0x4X/2xKQhx6CdrxANWQby9lHVWIFWovx/cjJWPdlIgK2k1hPX
tMn0eHUTOULSgaCggEcmm+GP+5qOS1HpvlzTWTus1dVMCZzv3Zya5gd0U6+1x6IV
VCX7tVMs0LcpMEbF8TRuqKnRgxTdX93js3aVPSAm8/wrGtU7gBACVHGjDMvnUug4
GEyEL1kD9I8zAeaeHo4RkYlr2E/nzcSd99DBHgay1h6awXemZn8y1hgu8wGQI/OK
YJMR55Py0QLtWX0Ddu+NoG6FGVb6tvEuQBymJ8yVedSHmAAwKJATE/QPJqZ4TCLo
z3PAeDvQpOZVddFnHIV3dC1jVrcPWr2HftR+JJkeZJlqssVonMcA7VL7rhwmZYFU
2Tpu2MukzSx+OmZWZ+xUs4uxl8MbEWIgdS3tDk5T0HLPffzxROYrLBvimltyASRs
e8IZ/KaW82hdwYsOEdmnkyn2nW7nx6dF0X2YQ+horqH3Xk9MVMhX+xgnbo42yeC8
iJZSuAI83qwit21tLFdh10EP5KrGEC6hndXYK8tUgT39NgKYCsNWqO5IlaFNASXR
CaCUYakJFaEHQ8YKVGna7G2OVQofoiCIjGo9b/YZcGRiE3rDB4ohlI1bwvsL8k6Z
9sAq+MBbkVYjEyshofxRs0pd2pvwUReDM1tYx2wwRQ3b9k8fgiBMnvC6uNg1MRsm
aZWAVogTgwI2tkpKQbsMINuy7D42zX9NgY0GHzSfPjc6gQdPFqwY8XO2fMh9m3hS
KCSZpOdk3Af7uupSnoeLWhnEum9v0bbOarTvmKVF94cZnDFEBAkkTeK8RkNGBPw2
k1Kmr7hnSSWjtzdA0RS0nE38L1A4XO/sfCyJv5Ah3q3ArbYK1T+F6flBTPNFfMPv
od6YCPVDHCHr4VoKLAvJe89ZbOH7bzuWAmNnsXVskLpVjotEpUhdBv+W4OWit08y
+Hpp3EEUrjowRJ6knpQ1RS24zFTIsujUJWq2F7xrcVu/OOfBziGeX3VhuqpMMJPb
pusb/M9TSOLUvg2945vZ01m9uxlp9BfL+Wo2gxRFFk5NsJxUzx9hHThhl6Twrtnd
UTWzv/dgNGksYXXzYAb5IlJPozczEHrLPM3SoRyv/AA8bZ/YJXL5v2Swjf9Ood9R
Bx3iOyh7rb4ISyhzuB0R5o53h82vU6Vdt89+dtUGlo3L/Y/46N3eKLjFxqZKXfSr
L2ouGTBRADbwuY692UN3R6ejjg4jgEa5zbztSP8/R3OiLvUuYZ1DBfArtxPkPaZx
8A4VfahHWIwxXfp2/QUnz9u3ry1w2Yba6vYolm/QCn2d1PsaRyIRCcPhoay1ZH3+
2sgvirEnnZ3KdHd9ppLpxGYNbnf7Px0CTx6yyR6Vv4TFBblhFoMJSG0svybim1XK
MI9nQ8oZhZQVVMibYU/toOd6ZAri42HQ0Tk3j7obiztkYgdmNcjtp5+IXLQ/D3sD
j3T11cFlJ0gDR1lY2djwLSsw62w5s7G9PkTsSlTKNxt5Rmz4dGbE6W/1J5st9tmk
iR0trZrtrshJygXncndRNkDB0X4HfSWIvUFpScEgXj2AtvA8SFtidpv9ddwAsOph
0HIQe6j2mPUTbNwA/CnJuvCcOQ2U22ELxQc2F5p1ZgA+t7JmaH88ADQM/ntJou46
Nw2vYy69kczJyfUqIWjPrhFK/cnT9GU1GOh84JPnwPtY1o0+D7hyi9DWjVu0oM8L
X3LDZpOF2hDWtSzEWCWmYbHutMokNtXjbjQCGGIlAJ8ZBcneP/1xG4Vkj0AO9rSK
gMoF3ZxhBN67S176zqyDFbEjSYUMcsiCIQYlaDMravSQ8+1muv7Fg3ZtUXqEtNSn
ZVAlHTzSW/ABa4RiQLT9Zw4WwV2H0Tb7l1ew1u23ZXN0Rw6eywgj833Fo1Rc1ZSw
/yEL0zyVnUMU3pdHnaFdtziJtlyS623IoOYN1tKmKvaDn8R78rm6P0OG3aOAtgJO
SK9a4ENZJRm/DzTpqP1CEnqneD8+yKhr5qKAHHg0JggA8ptGNzWyqKM09cq+dIHQ
EZWegh/w4Q8Rpuiq0Cvwat9LI0d0wM5my3NyA5R4r5ABnVddwvnyNsvjkjvI2JZ+
U+MdFDANAKVUwQjdT3HYNgzOzXR/SXC8tdWeWcraAl9giRMC8aq75/UQxYmBOTFt
BXkEP0QkIqTsBUu2asIQqppFh5ukvmtmmwK4vkollOLQpsmAHVskiop9FNXfdiIS
vFTbfF9x9ud0xdBnZbOrI7AFG6StRvwSbOyGr4c4sa7InEufqvgrG9g0SApYVv3K
rgsIEt4LjAAW0FOh0CzR3DaL7aYNiA4wJC2drV0cpNo2XTobpaALF0gRHLuRSTR+
J0t3BIEUvuC0/skG4iavDOZfoHayU+RflmqHUaTqptcoA3trGdnLux2KX6XoKtED
ySdGFOqRT4CydVUmy8HbRMudgiQ+YRJ5tJJZSfP8gOysEfKQ0uA5k9IPiJQehcfe
K46ll+7F55ZOBFyxQHhQOqYpL1c2adtdREuAOXMLXhqWIORxUcnFoYxYXKJh9au6
Y7ei6+aoT4pxyW6ZFjUuqGH1HBCMadD5ekW9BRAiof0=
`protect END_PROTECTED
