`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92UtHjgHszW+RCJM+HSNjqazOXBc8rnBFmdgRC6VSmrGhbYyhYcfnPzBoZthU8Gc
N7YaTCQN5ayDsM2U3Tl5vGSeroJZHABX9ahrYmmHDkSeNLaY+L1c0Be3CALRqqOW
X903iR/QpJNUo0yen64hSxwRLQ2mE0VsdiBnZ6zWpq03aqNQy3+A1oTdOWPwlYXQ
ly/HRet3AjUCMlgS3PjiFXXQasUfamRsED0SNLE/osrfap+knT8f+UifzzRGdxDa
i59Oqks4L83CGqcuJC7LRNcN0K/NdFU1ctg0zc38LLfOxx7gVBmdBJBHUAEXAlUm
FmACg1AV9f5ry7zN/BaxKe4wouELwVjMV9D+8IgcLzN6Mw+zw85AT8MU5Ru3/M0J
hKm+gXJ3q0KWVsZlof/VEST182Yx5ylFLahRss6iKJa/jbckXAuvsvDW9aCjuph4
/9haikVcWo3U/vLtNmSi/JaM2koyvZFVnYMAeRZBah58NiPP+2pOr/gKbRZf6adz
uL+HJUbLbbKnakv6r8c4Vrqhk6LQPYxNEuREVLkBmNEoNEkiBN/7uY1Z6PZw9l8a
QC+G1DIS8P3FGl3N4ccXq3WWqDJgZaZ7y4+nHYUr/T1sU2PkHSI4U+7fHg9cCsU+
7tFCt/3mhsLQiAi6QQc2MxqkFJ6J6OFApPAJluODM5iu4bPYeJJm4AP8uvlV1RNj
NFP3SbFLounh/RTkF56nrAe8yHG9zSrkTIpfApfpmbO+jTV0iR29oZSCE5HElspr
AfbsOViyzAls86Eato7dHcsp7E7uW48cfCYMy/9Alkg3U+5KaHCUAlQNpj8e5JBR
dMblP7lZgMrXuD3DBX2CjhYJX3VCz84t0Kgwnzjvo3rlHN8O7AzT+rQzPYJhbMKA
q36LBHv8j73oWOp5mhvw7uCwmdUZjsJELtPZjFITsLj9fi/wCd2NY6Bcyc8zofWk
2aSgZvVBbtWG6v/tbi5K13HIpq0W9fXEOJEfNzKlQeWQl9ScfTgkMlf3WvQP+1Rx
188zWkFFvS6bLf/WJhg7+On4x+xF+PP1KIkswBZSSVL8Axs+QbNxQhfg+/s9gY+O
y83Yu+geFriirKDW0wLyQvMAMVqRyX7OLpe6gFa850GBQIyrKI2UhTRSKcgWDGa+
38b8WvFGcm/FOx7a+RdHULqCdFEMjaxl3jYoS0bc8A+eAOVJdQqXUX5p5aN9u1JD
24xGjZoNImIkv7JMzeMfEVb3PJj7BHJvhlKtr4oNxP2MJWk/D7Ti66rhtK0L8gXa
W1e9fm94ssCxXw2168IsJSch1lBuV+PNkri8+F9y64Zk9ZRVpHCXlZrxD4HlSntz
Qhi/1etH0NGQ7Yct1o6mB2YIUz9u3X4iZkP4FwEZQVM3EdmyRSeA93D6avVfkwNI
sEJa/VjZdMYaN7GwA5ixr4RF+XuyqtE5wkI3fAQSmpgpAq95nuDyu3/ltgOZcaf6
JmuTssO2zSLBbpy0FFQrPJi3Hfp5T7HbL8EBBlD9dvkuzrdHghIUMsLpmUgXa2FI
QV3RMPsSBusbyWCpDff0Dad7N/xr4Uii+g/TnyVxAo15x+FsqIJSJFcpqoc3r6iS
JukCP5UgNfDMj52+ZcoGPRUZLr0qXePm3IT9ixDGA7BTPHNyXYtcVrcsHQrHI9rs
AB9FGuXWsLQbzrpD2v/XvJU35z8yTZ1lvCsI4LClTWNDqbNpovQnRXaHuqv3vE6n
Y77otK/IOUrKxuJ/vjewDt71ajav7M+31q8ykvlSvckP65g4hXnD3qm9FW01y3So
eCKnNVct/j0cXU7IkihT9z2TRBoAl462e8sWLnHLRkWBENJ5wRMzVuA7zD3aFWWE
nnG6zXcS5jCrnHIVvgNXzqX/BLp9+ZmblLwMEnS3J+uByjTpSJ4YevPMDIjlxS9l
JxEXxKOX/KSOLuYaY7h5I+hF8OVp+JivANOiRcm0HKOoM39XOchCiEAAtKPA3Jw2
fAnLvlRR1kZMVYshX9pY25jCzJ7JzK19e2xjXUR4KEHTMfRPieplO+HLTgHxVvSF
5k/6cRdbjlWDRdxaLemZ4BKP8axNQ1NUhaPhGhplX6lbseNnqX9Wq7ZelmzAUo9S
hy1UIyT6J5BmLkBqf/PtlGmug783RiZI70OkfMQpTngVDL9A92wti64+4KgTlaI0
ivAph/lnHnkkjr63vA2bUPVSqZZ23H8L2hmb70/i6z4Ow3Ju3FLlx/EAYR8acEB0
6Bf48enPAX3xZV28En4J6LVHSiwMekinrcimEQxzFvBTUwmZq6iEj9nlwG9cZMHC
R1UM80GlpVRQiFsmzEEwr0o3va21ZHWS4HDbQIEYWZf/ZmJLZB92223QllUpFbtL
I/lxooCufj66604CSdRsDC22QG4TmSw3ScsxAK+jaq+I9YQgiwY313VFIG7qBBf0
RQ8QqcVa6IQnZH/AH2VHsGJ+pLw0xNDFFzzUI+nNta1+UrWn2G4UQhrD6PvydpVC
jpMhALK2wfUprHSF688/XrT32xanLynn2GvpjoCIKWqB/GRlxsCETxYhoqBWftGT
sx2P0b6GyePTf85muyjUcJ6G2IiqMaeMxbnqcsPcosGLKoJ3lhyAkATXPvQMAOqX
Sl2VRLbMKbLn041TDw+F6+RB2Ye76mLdxMb3j4OzNfSZ/qXu8OT+v5ItCuFqLRyp
6M/DhmHFrOiRMd3gwU8IfeQRbAeC0C6a9vjNqQno1tzSbw10mOfmuBZGQvv76pU3
CenoR4NE8ZhoVnZnyVRIHnVYUcjSDdBuXRMjRtiKP9hdrKM+Ml2cxe7VVudNmkWb
HlDsbrY6R+EwQjPY6IjT0QP8palRS9iniIH/ulrBZutig4Ro2+4OP3MrRmZmFp1A
eGv98tckleAew1uvxGDnsRJ2aiwIQ/IuaXYk6t2m0KboqFXKQboDos0tFZMSH/mJ
rJ+kSJDbYt1de3gV18DGxyFzAD88mSmTe6GUF5/EYiHuka+Z2+Wu9JXdilYRsLAD
fj8ftwvyqkXU1LctkSwyhNfbHT1Alz2hSSJruVborgMEVy6Oox/8Ll89OUXXuPRy
joDg/1Ao2vMSJQ7E8+0cz+FUXQYjRAVAZ5/5F8oBUnLl+2aBUVS85OmUWxYEXB3o
0mBPHrHBjejL5iT9FKOO/7yZmT9jXWShF3DvUy+iSLnNrUeCQ6ps/j/Tq29oGqJa
qanFzKs7LuiV2fbwDzAeJDkGttViYP94rbA1BwM1FpMQXFaOqGNSX7r1fP84qSFl
g1QKifTbd0JSu+y1vUK6T+03Ab6jJneCOTY4iHXyNJaPpBk6I2mFPfFvg8FkLjM8
d77L81WkvUzjcIDhnEV55PRTZ+YLA/FlOnt1Kl7ZzZiepLQ+l2m2WNxcl3syk3My
ApXsdKm9NG/w2tl3FWu+mdymjSgvWXIp5CMZVBxdm68+CrFhlIxhSJOcGaU5fKvC
nLCjewYpQe09Ars78lBltDRksXJlAIELpxQoh421Px4ykCvI2pfq+1ZFD8RJMjYH
/3iiFq3aYRpvKBIj3ABLkyBUwUjrYiIMzV46C/cdgFGjrD2/pIa1Q3jWEcIDtrKL
PmDh7e/br7hLsT4UdQJLteh2nW8SpRbhG2qdUhi0xW8h8za02ajYtXiTrwZf5Jo2
s2Z4QF2Iy9O2P68psuc3d8HDn89S82KOSNA9Odc+EITZmzigmySY28DByCkEmCa4
G8pmm6a9RlleFDXR5WgfOihCjcxnNPat46Ns72lyO63e3BAw4pbT9Ck00VA176HS
XMLTdQocWnwY1tlBbCUlwISptxrTOXGDWjJotY2JAC4MPXGjkaHCJGvXdyUTCpy5
nSkrdNRXxGFUebgLZ3eg3FoUvwYPabvExWw6FmtRYhXS1AOH/Nv84o+bj1bValGI
hEMeQhsttpeW5SUldOUxv+EIuWnfnpEsC18r3mdWwmOvCFUs8cf0d9Yk1F13/d/A
d+/qmllses5BHNa0gDxdq+He5jBP/DTI5MGPCu5G+62Y2gDzW/VBl1qP6dpkhkoN
nc2l3Vh6FnG7QfOhYwNAEeUyojj2kAqRDEYIMtNyGUKTaeHEu/hGHG4Tnz1NA9ha
yRRNLtRKMevC+beOE7WnZA7GtL84lS82h9Svl9LTPyWA4mf8vw4W/DI/LEUXK0B/
KiIktq9A8RyAlW/MVp8vPbCe6eEf78HC2TyHSt7qA+3KcF8HCA2xrsLC4i8c/Opn
dyLOnJDhR7L/OsEtwWFHIQc9ss4lJV8SwMDB2jifoX6U3dw5YEViQMtLLGHUeK8S
VRDHOWtRx9AdOmB3qWS7hzayUaikStZ2wAKqwa1lm0LmCD22wHJbvNubJTLOlNRa
YK9uzVBdHZfhKd6lLy7Hhlaw32/setPnJkY+VNHdTq1PmB1YRUNtJEVFNU6ZGd7e
OAu/39E4ptLs3TILTEBkHrdudvjVkaHwa1wqi7rwyLIhsBkKZP4xloiCTMmQ0p56
kfKPuT7flNIxm7BEVID+BIn4vzExOwIA+aLlk2lHjDMyf17MSxCa4HZ958tTcdW8
PGFI45uvfMBMIVlshqsUvjWHmyg0JgHoUbNf234nFDEU+N5/qWDICW82LCrsUuVD
shwGyX4dwK1D6sLNAWudKwVlWBt7WfCgEvDpVOpY0Oi/+UkWSmxn2msdzJV6rcF+
Wh5VL7XvboVyFVEh0mItKZP0qpOgotMs9OSV1ufLXu1yFIkJu4zfl02aC4WiWFpS
G7pDn/iNHrPA7p7NT7m4YI3amzFI6LroAIJBjEJcfrLa759ZGAiPXCiKYyVJo6pB
+ZtGi4mQYFYz0SJllrxd6YAnUS2YX7ViwVdXSs7+mOTzIkNV5INKpdYvNYzB0xec
zi5JhyYSLBPr7hIud4gMsleNnTbTHo2udrxPtdnu6+XjZVjFUozH0tk2hrOUIiy1
KLmtAi1OE/pOuqNoWPWYzLRKbzieZKz2+MoTu/Y+N21qLNUWFd5pdr9hjc1mt1lA
Why9ZYd9CFtzXgUrJluAlfECCBZxk8QFnhmh+TDYp317lniqLjVkJaYera+gTDxS
+twSUDXHbu79clFkDyaMmMVKuhqOWFq7Skn7sPYXc5/JDVQ5KQEBN4DjMONDGvuP
89Is31+eLcUo9o2voCz9SfvRknAmc+I8R3tFnHq9NGDxd/A4InEurPqQRCc86vc2
YTTQ7VrcTkKxrEZoWAkXN4ozeNOL2uiSa2yj96/nWU36KZi2bqgIOydHTB64Jbvy
wUGjI98y7injpX0thJwikAUbd3UGSwU2XU6Sdv1wGzyKgJf0XwGxK41MJSHWumRB
1rbEY39ezZqWmUTjJvjKjsYp7fUbRh1MLJkWLcwEfflEnJPg5tPG/a9Q7hQXw30w
OeYg5CEywH6L/JrKp4qURzjCf2yWuJR5xK7FBSZGgejVkA1D6E2jBNG/w9jZpgm2
q8YKAWIQNt2a1xNXReF0+/boKu5vehJFUiDadlkewfR4DE+gWjOaeGJOVK6pP+/l
YPchcKAp7Ka0Gp6K9hfEmLAR4Gh9tfTxHYTOIAsh0kJru1Ab/6X4C/qNhHmM2iDr
k3aPlLzNyGWPwg17hrDnz7dYMNZTAEZzXjzkWeKxvBdirnfvSegD/dY7kgMOWh/n
nUFvc4RJuY0qsdNlQb9BMJlcIpcjoBbXQ7QoUHZzSAhh4iUbU4NMGKy+/+c5M7Nj
3hpxiyHEh+ZBRvtlhSrCmhcaHWEEK7pcTfj5FnyUcgZlrMq2uFCqbfuj0+6VEZMa
cvqALgBNWVbuOXlP0Kjl104yMIjnOBOObdkUB0j+qa0TiCWsiXcUnHfNFu8mXUYM
UfGUCx7HuiRWiVjsWu1mJH6oEf/tfRSLDnv5Ug8qpcM6XGXmzC2AHoFVA8xzZo2p
E07r96p0eTWI7NSohNOJ/OsDtEHibguofLKe2+QFo/TnkiPgPT4rronatrfkMk+h
DuAOeUjez7fJUn9P8sbWd/NU1Tsntat2a04sQwtahWucf8lc6Jw2KIjhwIt2jdF1
HL/TS2kPI78Iuqsh/kWZWDKAYZX0NLhP+MYpfsEWMWvRUWRPlVBhUln9CUQynTZI
Afv+iz/RZkA4s0nPwRCD7EhT4hP5gAPstocwk9YCu+/Qr3h38kbKa+49Xco1t1Xe
x5Ska9lOpNwN0LrU7RBD40YRXz9tIxZuCT7MTIBXUHeODARADhaYJO1B+On8IOi7
dfCMI6/f5TiQD5V5UxHrDA0PrKsJi5wylRmSKV4Z/LF3MVy2pSNB9VVFC28esOmK
sb7ptYmPA2efcNIj5XmqXk5GDBMzppWq38+QO00ffzPUVVqRHK1V3dl38yxer3n/
JA34g+4j+eKnH9TZLBYiZ8xGvuMd5daaUSCIgqrxAV3Vi6vdt7iRX9ku9dfy7QyI
B+dsUM7MVempR2NJw4WAVPnb7kKqfWQjXkix2qGGUK4XglI2LdQiyEQ5Gp86mxMz
NleDMdsscPdZzgWvLIdEELH5DfLfsI2cTaZadJeZ8Od+TAqcWFC9te/LJ8XpjVZc
yrp61GPWi7YVEKP1GMTHu/lKWoGBgyApQw0WyV+01yGR6pwQHT0hjDL5rkPf4Vct
kNjqIuyD5q34vAvL9U1mXT+5pYzhIcYrmIMOTD6U6neZw1KuHKcguOnOjcRg3QUp
4/ZpCOWQycDSIBJ6t4e1EnpG+eLaV/tlFU9PBiag7DiZDPDWJxmV1Ccq3WsXoo+s
a3qkgRtRnK2z04qloCz0v/LmB+craOMipwdWddqTEHoN2uf3UwdMcRKktDjiNxVi
pdRb3iZjGFKHdjsCYDuxXv/JQ0kwG8Aq9KeiRzcWERn1fc6tf7jUAeRJ5cgajme1
0oX8A1oIFWWmdpAo000kG3sRQnXWeehKZlGZ6hKHkEbAq+zZs4DKt9zFqYwEgJLz
00u4xPmUT8Bb3LHT2+hM3UsT8Uyqw3hEbgvR21bCpZqezwVrZTivM9E+sNtg3XFU
aeKdEfltqANhSHtb8ZUWgs/YAvL7ezvh88bkw5uAAnzxTGiwR70qQvJ/8BXhBxao
JZ7o5FQybsBFTQkAiL22MRivaKibXpxH2MzwfbsnFkJ11CJrRX4dyRbbODYEph3w
zoeE8wpbpRzYDntRFg+U2NDkPKpXeExhEWSN1MSh7KRfP3efzC20ial925d3OL8s
tj38HRROdwkWoHKF4yR702UMHh93gZviucBMYis2JjMoBRyq4hYjJpG1GBEi/Bz+
q4QDSVntUbNYoEutkqVrBFGD17pquU6z6MNiwtHF0fY0QWga0aI+E+4Fs98nmEbg
o6hz8VqL5JQIVSET9WukB6cV+1NPWb55d0AYEyKRG21vpQ9mifoftfV7nALH6VG3
flOqxLH2PA8M1RF85apBRwEp9dID8Yjn/LI2KWPCa4sL7vY0G/2JEs+S7btMKuw9
rrA2mdcaTwdc96qVayMKGsdImYqO6Z62CH0/1LStXr7kiNWUgKu5VCTy78g7X/NN
WVWogpCH9P1ykTW7cIc2czlb3Ngg2vRRh99vH6GDe2MJnyB/J+MUMLJSdWREZZMR
2mcL5mA4QPGRIxPIyFquwvc/pdHjLB50p2+XA4xobuUiFFhZwWjYYLzdwcgjsAOU
57YG/abBEP+oBEu49fuLBx2RxR3ijMckjND4dXd1/QJ3axsnvxJcghLlHyQtozZp
fWflj5luRsoQB0WY5cTBgvioUKgtd57zye8wkdrIT94QwBy/eJRcSO+qhlnPmxQa
OxytI8+kEO3vXruXdQcIhFk7Saj7vMP23OU+yucRFGp94u/xEXEPTyh8oBJNybun
GwNBpHkgXGTmPEPmSt97fnCuZygv+7aI9dp4GjFOyGGd9spdFBdjEeDQDAvypiXN
pQDSoEuBCiqedVIf27ks8FB2xLZoBBieQunPSJmDr97JnG2/wuHBFEANbQOxLpyD
xxNU151/jHEpyb6TrQMxgocD6aj3O+3v8nj537dJDQIMaKT5x8VRL1UCLHxFLjK/
ugYtyO+54dBq0fkszVDANTVCSvsa4ndDFAGRr4eCZapvGWFZzXpzZd+K4ddUPhye
EPTZGAkezINp6/PeUR1s7jDp1A29PaBBSoODK9dY0xelaeWhDXPqFCSGMqA8qJCE
5iN+OEjCz4yhbzL2RgMJ9TNKezvsinmq4FwL3WJE1YvwyMxOsy+GtpgwkktLDdHP
FumUkEqglorSKSXWUEhYo6BWC+W12HQma7rsEOPkticDVkzeZu5L7kKq0arXtnE4
x0DESrufm54qcr4FcoUm58XmjgEH1JoNHOuG+ZO+0R5upyMFghanIzw96U86s6hV
jCpHvJ2Jr7dFWUpwyNRz751bj8lGXBrpjnVXBPrFI5oSAYVoPzmCEkZ+iMGtobnC
92LyW9b/hdnXHadZbDyw4ZXZVYpkgfPOfqEUVPSC3qF+Kj7hkbTXFDBzY5SjNMjl
GiE+J1wDyuWiqdmFl1I249ATCdX4SfYyh7eh+jGzw7vWhEh1gbUkpyw/TUagGL0s
X7pcUWrq03rbLL9xowOb26AsNff8RPE9C9xsKjP2pQyXpAizTb2xgAYRAd4kXb/k
loK8+SNfaVFRYrOb6sGyYtI5CLXg9zhQYInhvwy2wEjB9AY2aKB8p2VMUZFev7mA
6Er03avjx0VfSDkJpo2ZzkfKzY59nvGp+WTH5N5cQ49xEo3HaLmbSNsmcUzkcEUW
RvmbtxF5tRJnHetfKvcNoJ5+SFfG4VJ2SNGmCoKAw+vZsjNonNmoGyEJnaICjkz5
Hwfs8rW1ZWt1hZd98Nkl6aGpIQMGfU/cjaJUOVeww9WlofiaZvXxIofLvCUnh9j5
szn/3CWDrJ4QpwvaE6u+Pe3KsdlSTmOioE6t78U2/u3BCSOeTiF3/J5QKKdLoWXh
kbdf0iX6xamRDHPN5rjj8Vr42BDRD7rIYSZuUcie9g9CkI+Z22J65T5xJ+qf7XBa
RltetInfE3prnCA84j6EuRrOxKXxD7hN+FlJaitCroEhO+Z2pCsgU56gdqtpLbI+
N7FybN3btfsJBGs95OYtupcs+m7SumO9Ioz/8aKu+tHDfuxhAVZPkwJfDflbpmaN
qgOr5Y0xOQCAAIQYfDf560jpF180JggLD/ifShehDIxcc5ptXKqL5mwgvagOiV7e
6baqdVm4i4+X9Uim9Dxwxb++UAhusgLQHtTDbnpvu4/emaBjCxntLzurPPGa+Pa/
lpi34j4kTCbvugZe2fFyveneP8xHEOi+dXUWmGvz+RB8hik3+f5iYkZzrLXLfpaX
M40jovCaNu1s/pplKaVFAJrV5YJ/hQyXiT+Z4dc5PM0vAzmxAkJcTN7tPfTsZtuF
ddxjA3ffT2STHTaWdYycaYb1QfCn66YGiIMiJOGoW8MzyVp7tbMOlwycnuhUyfZz
zNSv2sz1vbNg1h5BdIO+V/MDSc56f45fi3gTnq6tCLBurlUTAJd6ZGQtO1l13Qf2
FI2145Lleu3DpBSFxI/0vmoqix6BWTJ8yUSGBKhlRfLskX0cyWy4oxHHiXm8nO0V
bRvJIHNSzm/VcNo/N7QT1/Dp+jCf4TIz6pBEBru5WyzOCeA3BTsJ25eG0pJ4arTm
zhWMNI0GuckD1Q/tn50/g/myR+tsoSpKb5ktXg2bbPaT2ZSNPIRy01Fs5xWfVi2U
4xGceOQCfr57kdZrjChJIEYI8Xot5z6Sku0i6yhi+HBQJ3uW4gSrfVV0ECHYI3wi
VSJrtLHsOczqClNgp5+AZZyBJIP2nziF9f3JzxazT+X4luU28zO0U+XI8fwu3RJD
5SipGN8xgVePZ7LP0tsBR5xS3bPM43Hnu16/8z2FdSDWEnhRgYY6CRfY3FI7IAaT
jCaEW8h0+12K2IWoWBx0nC1+JZLzE9IVyCsypzt6iTbKP4w4RhTFpjDz0R6Jh2bH
bvUqBRFP7+MIL3CPqOTqGsUbuP802/MosNYv4s2/bMoj8kWlzs+m7jt4Pt37uc9y
1MHMMaaqIcDEIutI3Hy3QIRadMjwDeGj1lKCQWAWBQE4Q3NoBUjkIcLpgj3aNJwo
Z3g3LRbuuks5x+JhrujNxud4DNVHx3wTzr+sdDnY30fnKDwUxuWGnOAoKe9m9F5I
GnlMItIM1CIB2ZFsP98zqPGwUPPxk1hsMZ3cP1+m6oCiHob75mCGc+gXN+hrKyI8
oy5dRigxKVkgQ6n+8LdyM/tirGepwgIIbe6O7QIuLssmSKx/R862G/sWke1/t5XE
vt52Fu90ahmqTIYAsdcd7ZZaIcYbXvf48QynYG3Mghw1iVLIiWlIE1hjuFbDMjv8
u5RHkUSoLKgBar1TXrGhJw90J4vzpZU9lunggTlcXCa5F4tefz/KX47jUB6J2p7E
Kg22voNp/rl+P7KDo8xWq3PvFGriKWQsKDi4TQy5FMwAln8fB3eCOxPFlrbqFvJL
EhEgae8+CimQLTyXsFCq5677THgCwgTH9OKX49CmPegGui4eZkAncnW5CFzr0jcI
SEILxpyui7sLEA0h2s7MnlzV6678t8OcAKznrzkTrC5wcxUbJc6e3J8flPg1cDr/
LxL6SHoBjm+hfxNhhEXnGOKwm2plybM35L2JT9Rq8j5nH3uT51LRwxS8XXpLmFIr
LR1ZqHkNfcFIxXiSeQ3VxFQCxXLHcdh4GZNwiBkf3Ct/rireuckh25zen762drw8
ZD1rSfjgFPhKpriggnFJYtdV/VV6HpTP9w3hmdyy3sg94/qczPMldK+RS9KZS3kb
rHbxNDCd4W5lHlHyaeFxKDgGfix/AnP9twbB4cgkB+cKuxfKgqVdr+wJpUgH1cm1
zHlY+fhyQdfCg9De+4STjg++7wTGz+TBAKlvfzGbchDTbRA8XDuH8LWAqcJxkShi
R/2eDfYCZ503vHlzjDv8n2/tx+ltu9u9JliLVr+qSvwTRdN2O1RC+FIjMpqJjEpk
U5qnLlCLJzXVDzigw+1WVeDb15fa9t/BNBcXhyGZYyo/xexBqbQO/eqKYniNI8r6
8+gCiWQPgIM79RSozrZWIdGfMyTGjq9dO5W0ZO/vXM/FpkvFRSRtjhtZ5/TTlPKt
puWNb+Mt8XRrxlVmcNEq/1D9Yn+dBdltnkcNbhGhsgL6ZNXdNzVGfg1Gvygzcod4
Hp1Miy7JNGirW6O+fXPjojQ4vo6RK4IqNMvf4iYN5H0Ch86o7+VsO1jRe+J+ymCA
vttTdrRv9hXNkZcaTK7UoM1UzhPt+2W4lWPIU5WzXRRFA6/4LTPg9ndnRBDOLvpK
R8wBnbVbfLqSuXpmZn29CZzfstqFCr/Kp1uOeiV3jchCXRbHT9qSWzTkJioDKX+S
O5fVK4MwnetPrbwCTDvla6vWslZEgOradNLwxtZyKU/aXQnmppCehuqwwcvgxPDY
8C3IiaY5FVTJPAJQkjNPQyz3+IBQWH8Va1zeEhLt3qSkjMyUiXoRpaVwerRdNc+/
XsB4dPwU1nN1Iotal1StuwRlCalbvpVYxkLRYhFS9nqT583nM+5ZFo0EjONBmJZf
ds5gy8DQ9EPpG1hj4QeR1c642bAlxo3ARUlRg2cjee7NJbJriH8+h3buoESHlEfU
9vHuSzuJTel6v/fmpObV4xiYR2W7SOTdebSjbu8BHoubzjP9JcH9MTg35qy6FLuj
igaPcx48I9iTkFyGFNKqk24eBjTIkQXdBKD86HAF2WeUDMLk9S96i8O3O8J4on3q
Ay5ATdB3MKLEHW3mBAurbirOmo2+rGJaHl4DVWZE5wi7xAu7eH1vNi3PsNlUMz16
uLirLUgeV3UZQGQMpntGofr8uqZlkcBF/sCaLmsdiHJko2hmBhfFny5KWAY/vhGF
30tcVbvx6ksLP1mxAQ8n9JMcpM6saoI8pvdXL4as+jdU1qSb8n4P6O45Uc+Rayjm
teeUl7EzYg4RZBccaS3yE8saBmUGEBfInCFnkmLZgXIBjMtaZBrEyuVBBI4v+llb
mw0Ze8Qwt7JcEdkZNl2zUMqWCHBN9rdD6fwtyIGSDPegZxCvEXK7zg2tnpik4J9G
GQn32S4llQ9UgST1SMu375/lsXAwHusYSKobej4vcACFKoA17pMqDEVpoZTUayrT
lQf1ZRMdQwC3FPegk4o+BtLVupKySVT/o5tSpLPV+8G3wNypiBedJshHSXUsaNDM
wJR/2b/xjn5WZ/YG5lacwylcz/B//p3FZFnAeFTzngmGtq/b/z6vtKjRb2CxHjfT
Vhy1dzkMWcEzQM/yh6N/i5ug0aS/93DDQeFmlA5tRJi4IEu/TdUyQGzpjbxa7ImJ
/4bzwxeu4QMv3nadD5TGYMpNsbKwxVxq3yRlGh6F3w8DMD7PCTCi0ecmBQE3jNOK
MhFcVfQVcvK6HhuqdwdKI1ggAM5WjHpEiPIbAinmbwFueDAowPPrbWPfIrQhUbQp
rLKcZ3Yesnzm3yVzrwbAXoEqFCFrpp4RtoaxwcT2wWU4/mYMM5H6Sfc6lpNpkfQl
gALmHhu4KRAzz6U3tz5Jlm9dDYg/iXGpn/UeZ4N7WXJ/O9tF/CyHOwFswCNd2xZb
4QuvbgH9IYGShemASUfU4UhT5Ui98dL8saWKImGwr9jbIFE2RAIwxOr8yfDqEDDz
FOGuZqkNG81cIb6BoUT9RnpbDeBqIgCvBq5fNpLiWQf1iwLZdZmuwjVQ+c+cTo4+
i36DLC7r76LWa27nYqiY45+kbDubDDbsXcgR0O+PaIXOn9BR1W74WSXgKqp3wXcL
FAHKH7pkUH0YfYDJsaPzlHJAqP0v53dLXP6cjn6WfG8spKxmm/r0NMhMWD6bH0g8
ORAOs2uWkRUtnxStgJBve0IQ5ABX6lfL2u7L0VaT6+MUTP8cskCbdQaH9yqsh6E0
utYe15KL77DYdNDz4M/nkdyG1+9MwI/z1RC5miKkDN/uCX/UWfDq5VNhVKZsVdX2
JwhOtiYapVyNsTnmt6HyDd4/O0ZSokEOIytiKswZY0CyXOa0pd4gU6YEQeVa25LT
E+L6arOYKku4Ir4hcDBfQy0BpjVx/gL3vUNnY7BNfZM+BeFUGwPlfybsKxswNcQX
WDbiaJD6gtk+ULnTqkBubU8U+j/gdnsZ/OSKNTfrTYle7qArTE4H05ptGOX2u0ab
nqhMbFHSsSVdJh/NfrTgW/ridRmq1LmUhqKLjMxR/w+gfIBou2/WhEp/QflNzYJR
4NZdn2Vj1ohBo6nHGPG34mHd7oxpjsAOZzfjH3St3/X7hyhHBxwgBAZkH+5LpjI4
Lt0lAQsOVEJyOnCZ/ZQuX1ryKSLfIdDSZId1QBapDy3felJb9HK7KfaC+ezVJqMs
ss11/tL2ton5IcHHVJmrbzjncL1mYur0WCJPmAz/VnUiasdjh4ZLOTtfRglwCfnB
sWDVSiTjer3k8CVgKHbTf26hgTJxN0G53FQUnb8cVF1Vwb+TLJMCKMbk3LE+jDch
1TuA0b915Hw6K3C3fx5VpOY5RJUmmuklnhHSkcplEsuHTUzbcnoch/LzAoguFbZt
HEDAf1KAXmezv7UkXNQy12uiA79QwHvbjMbuSwoeQlRIGWZSZf8rqUiM4dj5gNpS
1t11ZENCPo6NJQ23s0bQIcfJuHIJsGHWYz8wQaOs4puZD+J50/f3uGmyV8EvGxAy
/oVlBrZXreVMXCPu+qj71L6KsfQnOAqWFvFZHHl0ImAvnvyiQdUsxlZ1ss2L78az
IyJesIM9x7oNrI7HVbqtFBseyE67amVf/xUH6Y/0WMH0PUfPk+uAfBYgWfIvye9i
rJtus9MzpJGyfgXgoO2nYMZTnl154/KszO7AC7kVxkWT7vex/BAQLH8OT9Xk/SUj
Pvh+kwl980Hv27bbwmXWOxMxA8bOLn4A216MCmOAePLdhlpt6KphdNmskr7l2nbr
L/CeAlxhRmm4R+f9/XmIzs9ihqWQgzTX0h+XvFreS6+HnGmR1EoVNsF/E3cKJ+Me
jQyynIdXWmtZql8tnLhdSIAa9c6rdkMUTdXazJvS2lnopsD2kGzz9rJnySzorIHh
Lwco9LNdg0XZSR3z+HI+Jp9lICCxLM2OP7OeV7qTly5IF2Y7UmMTqVIWsEQTtnA1
pikaheJNGZbpZHwAfvwLZSvxpa2A1kho/Ncc/tJHZlUPpUUhNRM9HrR0ETHo/rGi
oiTGtE2VLwnzSRmTQlu7jH9ZN/bY/bP7FaTbflFwZlmrsiiUxgMu8+UOLOLGcasJ
M8r1qtm8cxk19IHpYZQ6vZIwJq/Yp7vft20F6+DG24zpU5YCqnAWq/zx0O242kI0
RONVZQHardyTZBpj8UjHx/O51O46wEB9qD4vebEp9hDxUj1aP+8Pf2isq8mArwB2
4GhZrXCDecg5Z207uuj7JPnxjJKjK0ariihpAjeekSuv6orkcl3E3f7rHV0+olMQ
V5/dtlHXEqyCcYKd3kyx+yblzHj8A6ZK8MahA8XbxP1OY4955kPTXJySKHULOPfK
EJIqCGFApt3d50JmtZMfT+gXi/bh9dtUYBDsASlbllYWIHJOBc+qvTegZXwCthPb
i3PeM846mjXDLzmLu9Ng9jOHSJii7V8CjFGgzF6gcuOdQkf4+HZaF/SelCCWWZyP
V4VsZIXn2j52RIwUt49ihkPGaZ2WUzxq4K0cis4MWlKTKPEcjTmTQ00ReILJKTTl
MAPizQce6u02eAcbhVdomMbknfjaSY6RuRltvDkW/uAjgZhlwqZ1mlBFG1Z0leQF
3altMxN8ZXQAMJosZ4cyhiWZ8QDOGcPDlqEWH/eHUlX7dUDA54aPxSi5+CxWnOeA
NSD2nLQq/nqH//ndR9ov5i+amzOah8eeBlvL5R5kBKRiExvTMM/aN3nwYz8KxO14
LOQZqivlHXL3FdO5Tgi66MUBce5PlAmV0nIC17IiYOKlrh6L42MtHyBnE+jwnDyy
C2Mn3o7Dn4lilHvmXY/UqYnQ8frIa2dWfnROmGy6V04eOEc6daNSo0a7EEnxsh84
+UIadYI79S+0MeinAa6dV26ez+EpfGGUdCG23mzj/lOFUhMwwl0e4AtlCSIVp2UN
iDc7C/uUU6sU0Np24A4yNxmrEcsu4HelDJJihoD4ZBau9Mw/7XA9skvp72oG5p+a
KSMwkc1c+p0JY92MIeqowrzL85C1sth0zEFVPnNxsIBTXOKEtcR44aqhSG2SYEyB
cC53JhNCMhySZ4rs/OCheK+qndttKrkf5+ajVJ7/ZlPLtdkSkziFtAaG1zUUG+Ne
7suJjZSfKwEHdvUJ6vyzft0jwEs2gd6fYW2TudUncq0YVQfZwu4b+SfnUlKqPVd5
/JY2MdpKgWqiSVpSlbDb4hWEptLkMjip1SH24kTLF1JOsSZtIocvTGRLmby7dQud
ufb+EFiF2B3/vF5T1o4NaMKNwaDgp4/nG7tVSgquqOdLj2LukjCBdbfGSxhNGabF
BI7x2i7FrOMQIbzVZDZd4MxKytar33HCj9qxW+jLvHAlMcCFHM3hVtsR09ffHT2T
owJLrgorDGKmqCDXe0vpocz5BGqz7UkUdrahL7z2omj4j5jTm9sPCbT26IgukiKP
iD6Haxhkm65Z09fQocREmQVPKSQTa7Ac+pUoF8QaLvXk/m6Ayoc8tC+m1g8uOfCc
TQtqY1JOPxM5LQmZu8U21AZOvBqSxYxtmUL3xn3WPtW++P0llXzd+l5tdGqtK+SR
IGPzJR1aUK2r6W4yrdsSkXg6tIX3yGBZDd72t/a+1bgjcVJKOvViHfp1qtZG75x0
+Eh352RLm3gfZnYbjGw/tq3QTWCkL/FV4yDrQrlWx8st1ZTMrmug16OUAndnMarO
ctlzx2rIQrF3ZhSxd5/LFdgjyK/GEsPWs9VhxvKS9r06rEdDu2lTzNEuIjO2sNnW
JvDuy/HZ0sbXc2KjFi2kpiYwEzzkRmVzozEXlez+EK+TJlUHDR6z/LJHtSZvJIkU
HC6/9wDtNPMlyW/Xf0jTKXN2ZaOKnCBpx+SGmXbW02Jled1xiI0i+DRLh4QPZGmN
crS0KYpm0MBT41xwy3YFuTRRfqRcyG8Dp1/nUFOG5RgGTPSKaeZAz0p8TUtL6tYv
OTVRfqiOdKmEO+FXJWfxsEtlBxDwSVO8GcKTGr9UMpVAKsjyygCHvj2tx5YNse4w
Pnj51z1J+Y5JwlAASUHgEkD4ck3RHvrFTRRmJnDK+5iMQVqTGT8Q1FFQtwhmM5Bf
ZRG+k2rcJiDeDrx1DFMdKwspNYwFAoqYa+tm/0tF49GYTqxsw3AOIj9t9chKHtoQ
Qx+vHWktqzd94YrH8MgQdFIY0Eyy+b2LEfkiFB8ZGvzbyCsRYPg50IC9WuBP/H6J
zBzZ4y6g/YPnsl8A17aFvoWLdvDGtWti0OIgz7+1aRQ6rqNAOqazcKGg/gk53Ou+
siWubp2QYPgdCzqSBDDO4Jlwd34Uy8VVgHpxlwGcZg+a5ywtztftkv1USc6xutsh
DXszSgBo7jhkSS0RHqnwnsJl7WTotE4A8wvqDDUksRVRGADkdAnHwS2V896HcDju
OVfiS9gYSdvr3DlxcmTyO8bbd8rMjPIcGZB+TA62tLlDuMlyM9lEycevv+zEXO14
5PaB0bFufaAXSiNPesG830aX6O5oPbrdOFmijQnTpUazKdtc/Eg7OXT8eeKoqgN6
LOT01E53i/ybiAxACz63dbBfKWAhh1zFYl40X5xTSJqTYSpy8HSBl9PsXOa3hrp/
J8IShj+D5stFqs276BmfS5nytOaInQKc4jU/lEOevfS4JntNNT7qfH2Aw8Bo9JPp
9/d36WMlX3bgachNcVlFLIpsqfaJo+MGNCvfVTkcqoS9ikZGA6iToRbaOeBt1TKG
47oWv1IZRCvL9LH5aIIW/Ew/61cETbPyKPpZraUp1E+hTPQLb/GdCWL6r+E9p+WX
3EBqwdbYIuNZTf/THlY15n6tTUwhEsiDSFHpnaJ+k49qvokzh3Ek67hw9ggcwKaw
ONanOIYz4Hoxz4mmKQZ68tFgubAvPrEPeKuPfJ11VfxJTI1eXtAbX+wc5x80JI72
0hA8lZKJIKS9Un6CEGkzwbXEdi4D/gVNzqhvgZK48nXVn2uNAp7FyN9XqgFa//gc
ZZzjDAlOAhousPUHiL+jyyYu+jNBbxOFzboNEK+z/TZDhLAExt2uvPfPOZ5n4caD
+m0Z2M5xSFgOa2A9Hxdh0uiwRRW9JJVDTAUALB3e+B9vV6Npj7jU7R+mSBcsVpQa
RC6OGyKt6aYBhxNt+ojPnB+9TIvLpCnjFcQZSROwiYQ2mbQbaVgzP/G+I22Y50T1
VftSEs5+DHBUYVpaay+Pk0AKNq9ExYNfa582CDLD904yBPd3Bmn9cpsbzYxePQgF
5IX4OqFjmqU7TOKDCYdDDsqDb7q6NC7FVDw9znL1plbcVfSDAuQGVokpb1EbmVcL
/5jfzG3QZd6kBmBc5aR4+Vp1GDIcs9e3u+sZC5cBsoQ8kARyYs9YMfgAgwphgnWT
jGfFpyFXr2vJkaZVEIWX9YO9TlVMTRctF+EeoRPcEo6mPwxCoPsr3iNkQhwqsV2V
22CJcxaoj5lxK6SVujqSy1I1SG/E7mGpQBy4+h1uFNENiQgAKbd8mAOaSB8Y6EcP
rZUbguVONGgVjzUAvuR/QEK9xQ879QukPU919YF8KyH7eAH/1YV53TUzDnzeRa+K
1MpumN+8ecND1z2kWmJZrmLVd1cCN5FzJnHDwnL0hDgTnN8cw6WtyiHRUKUGuKPW
SFqm5cKgAzs5EQJUdwPHcL+W/6RVLloUzIrSUKb/h5ULshyzJOGaDeTWfCpu6YfE
/HmjaCox6JoXMjKNsWJQVl4zefj3+uwKa2CndLi2GA1IJE4jzV/ME1jr4dl8wp4F
GtG5nhClMexaxNIGgG55zBU/PSwS/OU9fzAOtE2sZfGBMT/p4n5fyQ32A/SGTdK8
VgpOiAov/AWFmd8WS/205QxWHwxep0vAY4qdQugbQYICko2H4IefY9I9HbjGSkIw
2AgKsYiXIXBEaVWCTtAxNhssksV7c+QuOHCE1cfLNWgy+4RAWnPSbXEw0xYjwsbj
tYiWwfbeW29eu/Dh0zLg38TJNTw3UFrnr+aEqD2rrNaaGm/+OM/Z8Q52rkdtvdut
zn8m2CuV34m/dOVGZhiyoeHuy+edlX9iiXzApqejSpZ9PphmthtUDyr8gNYGGb96
5uloA0xPigiPYuw52e1Iu4v+296ENnZelOrYYbIgj1k7QzwzdSckIovWOrm/Mgfz
jU6uIC0WAoowxxT2zxrLsEgJsbEikcH5rr1PRoeWIA6JMjs8aaZ6y4R9YgFRGhVH
m4HjIrA1I5iXYpKKMxWctOa/0G7Y2CnHXebBljccgjfDMrrMBBwbz6wK2PYiasWY
5PyYd5wBI0T3qDyGwbHoI/QQYRo3u3/dPY7JOl9nmT24b3JfyRmgBPv8/+w2Qi7C
3eoNhXbha58s8Ok/58+sPCeh1AFcs5miZ7juLCrmIn7bMGFcr669xTnmGFhEoJAk
uf5p2IFltKyKWZNTMMh6y9b0sWR6i7EYJHKfwtrfNsHZPrz/F8fnmP7z1vhkLv1f
Cnr4i2M8mMmnHDCla+3pino4KOvNT8oEDgeXBD/g3sZNeKrMQi3HHVwnCDoE3NHP
yJI6njOCbMlz03C92xF/THhxoKN/np6jky+lr2MQiadAlTMVeijCIqsh0LpBGf2O
EAbPxZw/DM71UCu8UCeZk+FGzuRr8/kmoESrFic+WLOpNOl07QKEAJMrq3okYPQA
FmWHAKKdvGFJ/wQP6vVJxrBQ4lSG1rR6aCLQu08FK9kSXhk+/HLVlvbzQPn/98TU
F07zlG6XbYTGdJJgrIFNKNs9tAEPX8qlBqDpuMovJRzDc/ZrwY0HB29piZ7NMX5u
yKQvhc+/a+n5g48xIiXAylmCQpU9yaGUzoYrAe2hRVfY4zS97PQn2z+l770hdPai
cdKLHK0s5UDBxzxenS1KUXCI8Wg3+7CBFF4Zts+bPmlTgZ5R9KpJu7CudBPmlCdf
zTdQpUKBBj8Vim2nqDSM9ERtypWhFAwv3MVeCwwUl3NYPOJf/TmXFYSK651R66lB
kPASJwx2dHc5ZZ1n4J7VkXQxa8kOwh26bU7PFvxzZV0tKJOd1+KaSkYaa85om1dT
vhnrIISBTCl3+kas8rh2LDvU0Sggt/+hlXXCvzaWrqCf8zHZFwYDD7vzbIyBBeJ8
EbhmjNKDleMXDl72IPS8nsL/GPc1dVw3wA2ifD+55yeg/5ozfF56+1yepHI64qj5
3DrHeIWhSGPUrNva083cwuz9vmU0v9IEAZ85wHMfKrgD3uDQelUnJE7JS6CAiWYl
DBsiSxo0PQ0E3fSCy8+MvEIzzZJy+R+8jNfsghKi57hf6T9rJSGjw8fbPSLj/NPx
rzPVd08FXYvss1CD2mWIs366OoS2z0oiG0g9Y8wSgOzwlo6azL2YL2qP0X5rLPND
95KeIuz3jS2dICY9iwuZEJLDeyT/dLh1DCb2JuIhrZBLTwCSXbQco8NJNTVh+mDx
Fc6fwlYcF1jhhi+NQs18rHV9lxdKkFEuU2E1f282yhBkP3MhiW2J39Bo7jK9w4uE
BYqjUhlVEt+0MLvoFt7aehSGJEYkUTLnS9+aHtm8BbKC9crIpJauP+DHWBZybZCH
A9Wy/XPzEr6Nvox06psIm9N0zJFOiEBxxeorK1T44oGlhI+SWYP2Bx2hEtbsbbxm
/f0uR8yG25zgKv6j3puXqEByycRM8/Aa/Z9YD5FwcIbHK8PKTmWNL+D3YESC5d76
qz1E0f+KNvcingKhbAAHvllhBGGUMYg66dCLllOyc1aCzVYAgxnS2Y4v4XRDiXSM
C0QAj47YnHZXTRKn4gkvzf2BijFxEKj/nlBEMMl5K9P73xNeJtE9kLm01HWM8qbn
VmL1qjTJ+aIW0Op/n+q0GGAl8r/ZXiuTxk5XvDXYbtaTgFk6thCqJFqf7AkWk6vY
eQWX47fBJe3/1UxGi8qKrLNfGuon/icRv5+fSjzId3bap9F4r9gLMtvOG//YVeFr
57dShsvIfjpnNQzvYLKkL1Io1y7wEy1csaHbTI42LrK1tVEtywQP6kLsZ5o2d5ly
hbZx/wocFqJWh+wB9JsVK/m/tAWszN1K/y8eh63PY12+LYDzlGNrFxA4MpLuuLsR
GyD/GD4L1ii1OKBug54Kd5Dp+umWSYSF1Qlk6TaM+hCLbpJWBNHx12ze5a8SrPs1
FdXXZVBUvh5yzwntJHuPt0MvQ6FpLl979R1VM9Jot6y4jOpy7Jq7BuDaQGh+YYYs
8upKrClSVbKKKGpkDTduk4ViSelxTnbSmgshMbz8slOPugeTjj9YAAzTZpz+30Yw
3xXUax19FlkRkFfd1sl78l6o79D3iaON+9bIOqU+whAbaIf4SH5MIQxH7XvqykeG
jy14IUERgsDSd+dzua2P3vhjeD09fv8ybcT9LjS0Xyz18e9k5lQVfD7pJ/9yxFaD
RzwIu4Q8Gdjr3FTuosdIdEJ/cRhsOeih1tBUvs8FfhNlAHLM+XtjNniG/Bj2Clv1
XhAyC4IKQZeEZtjh2cIQXPWFJdptdj7fUWjj/Amu6RAHag6MRKmgA/KLqlvFEXcg
xuHqN8zYbyd8KULfgrJwe21FQz4p32Kf+q0Bp25yVJqYqh8C/fRVyO8eLMKxinEN
egt199431i8xTGsyo8nb8d2u0azqNopCam+5joXDCyW/mJPgFaOMl3x8/718P2sg
YprPr5UuqbfpXqb5+YezEXPR90kDdl4/ZVLHCTZKiK2fsIb8oTjBS61vXwnQCalz
beaXa+USKSnLfvmNNclLR1XQQ5dVumUWOD3fo3VBUdXUXRf22bTE2io12rYmtqH5
5AV9e+xxF/L0wLm7TnhDxSzMznGhamQAJev+FKZuzsSPjoc8KbaiGmA6yp7hU7Qu
xwnVyON70nf9B9gDraxFl1xq51LpAiYtSZdHWlOieKzmHdrDc0kUqzatzNbwSmKh
OfIT9jw42V8CzdOygm51YJBP/2ScvNQqfrMOSKuCnC36vMo23PEVPnmb0hU/cF47
1UIpX8vdmdxxq9zc/0QS35OvJ3F1yNPR4H7FJPl4E208B10XLUV9fA9PwNqkeFSb
nBfI5JEkVRyAwc6ryolB5NMk+jeXl9zdbm6bIjkDloOFpqQtHqJVSc+XpEri4w8b
NDzBCPCi9xvTqP1fB2milTOKQB3JdWVS7T18jHT0MW32GdkHwzW0QHmJGr9LLBpL
haqm4JlAd7WP1/GUx22mYaFh7+89LBK0AFZOS3kY+k/SjyqUYRv+kqekD4pRenOl
tM9cJdA5DnU9OYuiBYUQum42xtFAslYCb6s1zD0CvNMcZtZl+Ly9OhunljE7OzmK
KnOOMjMzMQRpWoFuK6kf6U2Ib8DTKoKeIqsb6r8ps9UqsPIvHmsMXbrzH3VHfaam
nqJ2BM1PL+tKTfqXYWc3eRtaoS45MmPR+FoQSvEBVXJgcGEKwf8rD5H7Otfcf/np
7i5gL3yJCzkORUmIOVo4vZ4sPJC4LcgJDSGP69KpvLw14VPb3dTWZONfqO/5Qwbf
6tlr7aASb6fLDIwvICOrR71v/KJM/+OHd3xDkvADVpYDlee1cpkBsTfxBCV2yj7P
cwaytJxWUvrx24tpctAvc7sQm9r2AkznpU6Sg3cfeYNrZFfIzozkn9lfrqsC5GHj
8ak1EdD/lK86MhSzG2TaBi4bZ9yVS+KTmgwjNYdWa6RN0c+EpX+E0JBnDhN2OfVV
KSZrLL8qIIoksN9Cz+/eDyrd2jhxLIWcJumM25/1t5b/7dXV8MhqGV8HNT4Oq8HX
zmKK/J1eFp3TkgBx7Gs0l3tEDXkaH41hy/xkzoss2Tcbi/KIoW0TLPsK23LMQ4YA
7eMgcBiR9V2vTMaFgO+UzpW6f2f4duht4GVosJ+SM+luVkCyyECUY6vlRbayvWQ2
UA7Ei5Jy10oa62JisTGNOLtDwbFSR2XlS+vcBlpBa+5Ij/Pn24ZqXDy83rH72xy0
TowGhIStngPKiORKsJyoOip0OAooOBlhjffd28Ts7ku1Q4BeUm7gQ8He8YwcKdWt
vqsC3crGDdWBf6ufaDFby6icbnO4U8qgSencwx2nM1Ict+CICFTSr5yYmdEmTmz8
eoSdV0+YFWqa1GqqmREa5tdoxgjDQKpOU6qzvCbBChUgltr1fL7Dz7o8GNqpfsBU
9kVA5YLdViFXyJwFsn7A1jLzkNFWifvLnLUx/2nTPBQeJ5kC7VoM6dsVRqEcxcup
GvDXkLMAx0BfAAASOFWxv6bKU2RIv9KNEyndc4963JskAEdse+8I88SgodXh/TtM
EAEkCP3fN5qcZE0Vx2FgNqWW9+JzOfHmldH0dbJPyTMw2JJXPFkv5CPU97ZogZNq
Jzh3+kgj27Um9Ma7tVd/ajV0qwDuRIEbRM37uavXA3XMWVh75BAUxW5QTakU2ycq
iUHhQitYXatLJxAN2qjrdG0Mu/X5ks/2KTSbGRiild67mnRSyFdjczUtromvkZA2
UWZw4hbqgFmlpe6vA6fg1rlFRfyDWwLMWvDVNrb2/AgeThlvrLxnll5JpYVGkMof
CmRX1JmQZGHxdEmQVvmSayqhsIXhufSQPStB6dlTQKJ0p1eRYP9PDv9xPrxVIHSb
TCaeXmpkHHR8aeF9kTuPyww2e+RyM/n0rdYl06Cijtvkx/nsW3NCU0uQ+eBiRYxL
l0qM5Vl78aB6H6b6TBP3LchojPOgT2jWtPRArn/aAfBRU6cozFZH8rtCpo+6XFBo
j+K6II9TevJu92A6+nWV+a/3QmQaVqZnByfHWOunTERGMFFSSfFDMZIlehfCJJkE
KM/IA0npLSVuHRYjOsQz+Q4kU0Z0FUoYjcC5zarG9dkZ0jMZBjfrwN9iN/O46SV6
JK1JOs88DvhzCLRYQR3HOeO35syFIkk/aIv8waVYSFO5aix1LipXfE44yyJzQLo9
M1MIETSlaUG7qaDl+SKOn55MeVJuw0qhh87/xAYTgvT6spSwIkbWpp9QvZ0vQxOn
xGDmhmuoDZfVfxEV6IoQKP6syo51Z8FLsbnSL3HnS5b5ttloRijZRa1jG2uHAJSw
Adm0D5kGtibAOA0BaZ04L1hFszGVL7XDypSWCn3T9l3aOceZYlZwx9iQPzPXGfy/
dRNC53R1h6q9C+YGvfWRVFgn5Fs3SUD88dzOuctHbzN1u9w8WIWmBXJcUG/7fQdz
Xy2WSNnGOouhxByFxk/1svGtK+FkLYHbdNVqapJvNb3q9KlN0tgjmD2sVWqGXCmy
hCehtlXTxmgSG+hLaaLVvERujxqxpy7sgAF4ClYrlbOT/WvbXXbEqE9GRczIOdYM
t8pukoG8+XiPdyIW95etMO1+ZsaN/GKGHo+td0psF+CWcIUMYB7V5jOnfVsgzgpr
+Yk+/JMN1zJU9SQ5xp+NL+N+rz9loG+oVgafcWyw3Ms9jKSFW5U8adwJUxOlIh3n
GiAzKde74XJQuCn1FLvoRdllXAPqR1ObIK9ZTvM2oia4aVCwIEO12cpr3Jt63Ed3
0aMPlfsNBn42ArHN1Oa1xfR87uCUeYqrFn3ra7UWexTjSrPzsx/ibziYyuLtkREz
6bOs0Z5PAPtuwQVHaJUu2pt0DQ7TPpyAsyeH9F4qZ8O+P9FdeDfuZJhKusxDMaVc
r2poPHnm+jbx8uugi734z8cbaQgoiFHem5+R40UV+gARSq3AugYSkPQTXGYxw1M2
8zgQ8OZiYH/jMOtfa60BK5LUi/XGcaH+1Kh4nfWAjZMgO87tjsIQZHn8mi//AX8B
CDN3fJE6/Yi+iorlWkQuU3ApOwWrcqf30U8WTRju6Mn4HY/95uYthirymMRwBs8r
CaCHf1QS9cFtFroqqP/N7XgCjrbTQDWQ3HQC3yoiek3utY7CWJJVdv09G7jGO4jl
4YC26JvZWxFxOfyt+G7MV8TPmSwltEWrtGeC0SGhRsEI+DkUSXzr689WB7KTxE3/
8CBIIUmQl0ObjHphcdfugHtqWve/J7NVsyd7JtUd25QP7SGJzyYqGpZhoHUs+oVa
8s3dntfIe1dS6NjexOsUqGe5wlgxbLZazGaaH3nXmv1Wif6ID2GkkRIWHLCJSXOo
B4kV1X7oea90dCyPeuKyXTLIRRCGRbAC/7WJhKk+9PKc4+s7PXAvfXfgGjbpV3kM
LcUAaIEVBZSyJaGeq7daaSPX82e8vsMLuwqCn2x4t6iY6ap7OD5rstz/HRCCSqfJ
IPxE2TlEMDksM/p7+NmadEjRCrP7psvDQQjuhyeCaam9BdtBE7vYAOuBSDamSzj4
Z55AIyYDH7t1wlehXDq6ZUv2CPxZYy4nBUyO9qZZdYLs2VyaIqlcQ3xbYnhNOH+f
Vv+mXJThhNzCwVHTsao0ZIYqPEhEhgiLSjE7tsVh0Ze91UvNGS9Lz6U+DtS3qwlH
DA+NulgmZz89YSC1ybRKBUlvH++o+LOMZCqjna7M4ZzwNaHfEGwDvwJWZSd592FC
UicRG7r8D1mwuHWHkKuzD472vuKikkEn04NRUHin7LCnpEnwokqh2DFCN/yjwO4w
/PfY+ppbuGycFvHUWpVZJd6XqxsFwQ9XpFEeJjcth3PY/z5jiAU8ZedS9urv6tIe
DMYdjmt3RTWsQacVghwkDSrGvo0WjjsvX1hDnmPHTIGRl7qGwL4OFDtVzfHl0yxS
qywI8TygKABRAetue6qL+aF2cvNIelkbOINttnP6ZTO3TckNVXy3H/cQGARNlSg0
FF6mP1BgpLPgb738shxjtNDfXWyRn2P8fGBvhXl61fdo/wdtxfa14VwttkfuJ/cG
xpkFdPoMZEWQ7TzNCh2qeZ+RnK5NGCak7uG/dfmokKhmPGERFLfJlrbUSm3Isp9C
Wsc4+4tGUkmNzJ0+N/0Qa3ZAaaK9uM1mFGBh9g/UDjPj4B8GmaduPAah37T0VFdI
t5F0F21r2wC/Ua19647eCQEbc/yKoVagjpjQcOo22R8E5sfLryBgoEdCaDwZPy0A
UMt0Mm9yRzeHHhbfzquoKKlyk1sEC+cKMxDE7khq3c4Q0nYbkBwl3zguhcGUImhL
54aNX9ur6/cWh+Ykbepwh59oCxwWBgbC9qnpSY9J+R8ePiaIj00l3h4P8hYY6Nr9
4wf6pqeKYAS2Z48pLDtrCR6o1Xv/aPIEPUpYSwDKN15912x+V4A7bAmFoB0e/0hh
zVo+Cd43XuZlNXO6K+ChobTKjVsmM+Pg+yG663T2ASQjThz5Abeknb4jqcd7okTb
3c9L6jeWr1If9J5jOhzvIguZyfN9lgQQsDQLm2T/KzXHQJLc8EYEUDb5np74XovY
trMs6reZ5WSnyYDtFOEcfoV0TbE6k0hEgscf9breuWwCyVFVpIl+zqmRkLP70CAr
qtNrILozPl0TLXFq4RqzS7izysfPJIOdroaN0xsgfM/zYB8rvDOys1z6M0G1m3Sk
6TUguL/ZSMwhjFlIpfyAYsyePivUfMu4SWTw0WpbB/N1knUi/yj0oRa6LEbx6Jnm
wn4fdSBNW7UIWgjpeluWIr4Hoemwx3OVtPNU0Y+QRMCv7sHkU5Aq3OnA9M/jBW56
EPsMwsnK3aevVVRFQs4H0GAFY9UEEnfzMjYwVc/WceuVH6Clne3RZfOUSskF63QN
HeJ/s0hZxqx6gINzigv2xBXN8IjNxvOLcZ5ldmP0Hm5WXgg63K1fAZi7JFRCUVpI
oitKwCYlq4OX2V6RVzGhn+xUBeI+Wf/b3fazb8az8FyIdLG1ezozVAiqpkSeHkFi
gL6/5/dxmsT82UYfcTJ8hFWcagMq6H+uLElBZFi7jC3V5L5LNf9dszLl69Vji7yG
FEZEro+P5VE9NnjQdBFh1gC60FU0e/4XFg0t9bg2+ycNdYwEQJhZ70k7cuoB5Tmf
iCJxtgZXMI3oyerqphyXs3VgMc513WqQr9IDAQw7llePxnEyum0YnnFQJPzRJc6/
QnEQ5cysggPSxWPorZtDr6sKj9GXk2MfJro4Iw4I4JdZNHB9nQjYky6C8d/80HtK
Jzzr8uIyhPWNV+5H0yAa+n7wEbCq0R3It1WCaUTuaX0VFNU3KuK+a52CYSWfC05e
WcmzdJJZaFfW3yW8XQX8Qyc0CEdZdrpFtN8PqhKSMN6Do0U62kEnJdaKOqtxdGXf
nFzloSJC343ea9/+rpEnZdKjKzhNaVzUJ6+iZwO4B3pu3ULJ2IL+MA4egJxMV8Eo
wArOi+M4mxaL/SIgRbiKngZxMVAikpwRvBxzK9fATgDTatKjb13mq/BjjqTRIcB+
e2lMRoeflOqZbiwJsVXC0e1GfPAW2/8KVR4lTIhTUbb0BTAlPrZ1o31SdNYvkPtx
jln8hbRRkqD5OPep0RllCGCY+eU/5zQcV7lIvYLstEFzM1VHgmeyon0NC5T6kw5h
dUF1AXWW0l/D1zrsUGzQr51qm6VA3FgsoLZPfXBF8HbR7LtURj9ql5I2q4u8goBG
I0N2qC4QrY41VNgdHvIjprrYFcfF4PwHUKh8zWQDHqT7dWHfcdOfOVeaXtvWnqmQ
mIsF5IvrYARr/sXmbezjX9fMWXP5DSa/l21cP7MwbAxmS/ng3MQkmhBTH/g2+XSX
XD9ajp6mR1+K/xXkZ2pmpSXxzfOiN5xT4QcoLrYiPBnd9P8Ky9bpsxFiuwrbntLh
sOPGm06UoRi2ge/bR9QaD/He95AQVp3n6AkGlmmR4A2hF0sM2R6ZCeasToGxcjBo
bqjJBi8XmnVylyNlgRs/Q0A0pDVrSp2K2fyALTsVv6uDIZ/jTFSsO2Mpx0OBcarE
9wquwziaZUT3isp7vzNXjRr3A0RlL9i4scAne863gtvkKxS2a7csPdkIZddyb8dw
71GkUNa4MkqSrsmkx80EXtzxRpRcnqSN19g0IICGzZMHsEYA8gL+WoO4PQ6QrCyT
JnV7MoOpvvflTQq9Edlw8HdDohRtoiYajUXYaW7oD+hZx7UZgVe3r2Zd2bHZWrbS
OsXJBZUFJ+uR9S60MmL6M5qR7opbGysE9GqWbYncNlHMmlu6PrvpI9fogJj3Prmk
NhJOSY9Ma6480J3BTdiulN6O+gqAN2gPePhssXNzF3BR7LTtNVoIQith+DD+mdVX
wlJFXuJo5ARFCnqqkQn6bnxYQvqbR0iFf8VH5dRpGmKRw6MKlt5Z7TGkVRQaSq6c
4oWkyQjbjVZt5QEvKJTE4JsGrLTysMNHFOBrVreJLS8XLXabuP8k5k074FZXGaM3
4Nd+iKdMc/cXKANcD33lNEqWzt0yRNC4QMhuWuJs6M4jnKejoTmM4qVY89qj5tdl
8FD7iNcYKMFNzlmVcpp1Dcvf/LPhuKYfFUh31dd+CbC3k3o0qoRiD173g9k2T0FT
yc/pu/YMdzokFBiRy+OBv/aOamUuaTex+4BAsLOwxXUTn9CUwhDymvXvG50N0uQu
aEWuwni2ZhG1aUl5758MVUktDz99uZBgMVHs6x8o3cqp4Cob8HN0uzaoQDemyrB9
IjEG6atwLq07norto2UupG1Z5D5oMj7wcMvtAm0rqum7xdwBe6cTnmEC99fY3gVy
66it6IkbrGBAFbQ+NIubXnFXxu5Ia1sTMOuLqdHii3wkQaV2vx8myQ2JG75zUsCK
XYkuVV+YldjOBtxPg90Mp4Tr0OQzRBYj+VxvRQKEyR91M58DM5OMHzo5UaBOWEp2
POXvHbIPiFwapn8xfqF/fA+b7tkN1aMJbz0TFpTAnr41Xe07+bUsWWS+Xct4vYLN
dB/aPO6WTHbKzuAK2NuaozGrhcgfAc5td9uzjoeFG4LbZBQUNzhZD9KMOZ8gZRsG
lq72PvLRwoqn8X7PsgsS6xyyDvSEhgFBxT44Q6Czr+wppaByvZRGT+3bN/3SaPwX
LkblMqiKDyRP+rMoHIAPifL6Ao8KRld1ByIHfvvn6q1xS4JHUC5vNA4+ouQ60F9z
mdM9iazZrBVWH1v1yL2Pcrzh3rDcqCBYxMGc88pCOCDlIDHr6SOWFF8q/4YbWPTB
lpRcAvtTVp2x8NDf0OfImqUM+icajHDlroZBPRBEBxzCFe7scEdRyLJFGJ1Ao0Mt
dVazNUWGVErbc/spSrQn/7XOXwWP6gK/r7ADKb2GxEVlsSpbhdX77A+HWUZ9XfUi
OjlcoBNanF0ZS65N3RhglS4OcoO89hBE1CnHzK9rocl6uCV59qXdvMww4VHfbxMw
pCNlCqAoV7Ha6fAsPIlJfcSVqI5H1+d5sqyY5m5KUtpiWj+9Wfr39JeInGGMsF30
0JvBlyfhe1wo0Nxq7XAn8l47B1pohwWAaUoWDt4B2vRC0gr6uS4WmG8ZdxtWk9i8
+tuBMa0gqoIDcTZfgpyZapNRhsyRrIJ77qv+89obvrhI/DgjsuhPYQ+gdP+Ed/0a
Ya9JypC58znXaw5L0vuwvZ6IhdfCWddNRaPp+UGeUxgaMScLNeIdg6lgevYnwOmd
cTsee4BeMfrZun2gmOf7V9cev8o0nZNjL4bQJg5iO3epZe5if55LFznVHS1DDIdE
l3Gg5kZs7TatLYU6+hP1ovWEZXQIN41jfGVy82BC7/lQ+uxYKwHsW5+pDVU4Aefg
MNnl4y0EBeurLqTkNhzQq+QmpkMR0e1SzQpp6TJ62PiaRASbL9b0MpvVN1i+Z2Ib
IGp2k26lh+A2bl1Xt5GG4Tsq8i3A0ZBxAjXN653wq9iVvphgYiKAMKaUfvs21/iu
GLeDbheYre07OtNFp/G/lzWBnZ3/q6UoCdOgw4i8we6R7TGOnAkteyAn0oxSCOx5
spArkxwP9xRanfQalkIMIwqlceZNSzE54JBUgX8vkJAkADYKBNUhoybs4NURs4dC
n2MCO3ippKACS2yIxZJzPEKEpvGG5B21H7Zxqg7ZDVXDI+tx0NVptmjZyqctsSoj
vsP/KxL7aA7QMkYCkSxPprLsjX8aIW7qy3H2vCrRibVBUamVCX2dDcyPhOvJnZl3
a357FhzgpGH2UDKIPg+Q68X/QoxI++MaIzgX7Bg73UskfR2wZJ6xkQYBD7x834DR
aThgYz6SP15X5wQ7psLjX8oQBgPHmXt5nBwXq+gf2wCC3DctKW2Fv436FxszxBjs
txDH/18aClwrsISNoIHfuq1WNwS4wbPt8bQIYrAvjNghnLM4a9ZPBrmujZkBLKMJ
CEMZkB40BKSfvVu8tJyFUGICwqInLhHm8NanRgQ2kni4/UF88x/JKZfGeE1fOKJX
2P6tOZFj6Hz6eVP8VxMPQ+T0dRrBcZkxrSyxu3XBTyMdrkGgWqDpj2oQ1aOxtvX4
k2JKqPGGDfy5OSTy5sMx7z5k78mzTr5kMQRYNmxhYRqnacaPmp0gjgLqb3GmzSDf
/LW5Hgh+tWB0Cr32kCETIVYq/VE6Y+cMwDpt+keHl5ErN9a/VRCbqbjQnAGzkQrX
AIJp6+qWpy17ZGktc2kZfo+eIv8hcxCparK3Y4KjwDIUob4hom7fHXgGNA2/2GW2
svLIVsYHlcG1Wq3EJr1O3Q==
`protect END_PROTECTED
