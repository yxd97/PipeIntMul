`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xhHcGWha2FyC4KF36+TixuL0cfe8KEW2vjb4HCnJ36SEo0ppNPhhycNp+iJ9+9I7
y8CTxyBlAwsYspTkxYbfz7RfnrCsQOgdJx1h47zypBx6TzefNHPcD5ytoLzMMhCt
lk1XSFyFlNuiLkI56CkBU8OzVV3mnaJXDDSigos1iTNhFjupSAxGMt8TLPUhWyHu
zvz+iacVsRijOfQopVhbOrtTbpkyruM49UDKX/7D1ky2t+bVJhVX8qdppbOSJSR7
Lj5/mml9Zrs03nIQ/U+9tFIuhwsw10R33+1jf2+bFqhalAcNbayyQmX/SOXRLWFC
lR5eWdihLkn2NZKWYfFv/Q/U5wW7XzLDdQOK0iuXUrj9v1kclCH7/tERGF9jXYPv
zs8BrTJ7RNxJu9sl3GqUdS9CIe4TnkvmwjFjF6QAOLcnGkOiTAceRiVGDg+qfY7u
YKh7p/uUbE/B/FTRc7c8heDHKvw9alm5QmWyNakcXjmRjIGNlqGqXupD/PTHc6qk
`protect END_PROTECTED
