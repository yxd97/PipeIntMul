`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZnNFB8KSqWO5EP5zdjhkNnWuUp5LYP4tY+SxpcmplCAgOymZV1nnfmFEKFOaaGc
00N+Ix6a67G1h/ot21kjyChZoFPa7y6vbjpS6Sq0ktkhAv/F/SM6mFe/cY3ljvyW
FP1axIg5rVK/7MGhvShj6Q2qDINDsFX94VsGDp5hNkEfRH8Yw25urOy9vvRZCypQ
13YsMeajV+xSb5m4f8fGV13uAHQnbynBAfCDBBpl+TTyPjHgBhHN8mW9xOEcMQ/d
fEb9tBIzP6wLbtoC8MH9H/BWf6iaDbLXgHBBX4pPsDfzObSD5oljXgELzs22vN8C
/hl+kfHJEb5dzgPcOfH+4T4818Z7RBX1Wy7Sr/g7LW1HHCe+coxuH66Z2hEXj4xa
oB5AmRclPMJIOubIKQNFie56ehWNtFaU42gYaG/cuNBnfKwez/RnADWcL1eZSA7R
R0D2eeDsbHX6b4rampdPCjGXy468zJkdkU+Qbd4EIC4GbJAPQf8dOb2GpnJgzcgn
ULb0f58/xDJbMjogM0m0VpBvNY40CrI1EQ31OcWA79VyVVDOvVCzaJqNQU7dxWv7
TYe3TMuo6xCOJyJY/xMwQ8ZturXlb8FTamHptgq7TvM/LFLg6L+qSaXkliEcyH2Q
odwUdKKUetG12Zp556vrr9vPp5ikmnFuENTTwD3w6bFTiBwFWa3n9d3hNVlO89o6
DfzD8M3T64SszrHqy+hh8M64XtymuOPwKep63MCEikuLUCSoBu9CTuI9yePUPoLG
V7f5HBtpXx6vG9X02I6Xm4mhLxH1hIcGW/JavO1s5b8Ot0uRHP/asIB8bd1wjwez
sRetOpRLC/k7YKFBkMAtzPGef4pAv9voce1tptXQZ7lmimmKkx8CSCulorNrkoVW
3fJ5+gzBeD8Yrfbst0z7lOzwpy1iikQvggyKK+1V41kjf7XtQwcVGWitar4eP4zf
mvWr4J8BHxpgV9HdqywK9eJmEpemAJIyIVHAEF2PJa/NZrBKqvg49n5xLy4s6qhR
Yi4VF5eHWt/dIPAZ5bGDpkvILwPxc3uQwBMrZX4Wvidpt+dlVyUrO7IVNFM8UN8S
+oy3dgwMsAri0po77zZvboZv9Mnna62YPQsN5iml/oC39hQMrY7XFsbyJPa925Tz
2tQ8TCinRlvuaO4OM9LL/GBJDQjrfaB26cEX2KA+xvUtfinYweREwSHr2FJTgWRd
`protect END_PROTECTED
