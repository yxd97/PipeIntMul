`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bt2qTIdJRVUV++zp76p7BILbjxN9EdpFoAsDI8r+QqS7ApoUYMhBV+Ob3Kk/NLY/
I+xeheOKnMhVlc6962KZMjWqoMHgyVqic4KR9vpGH55VCtFHgoNpcqN3VDjiVBKZ
0he46EkpT96qxEJUWQpl/wy7/upifv5vJGIsa8JWRc8e66/sjyE0IS7c7n5H891a
/T7nrrz38LlzQdRdA5MMI8GEBG98X8YxsMgiVNbUcHIJCuQM0YECgY9KRUqQNC6O
6/coG0KlzuSM0OIQlag8cH4I/6c8xmCEpn7xelgNkaM4JCxQ7ptnEN7/vlAqpcvR
kv+xP+BtAiUZ9/pQjJb1mH51O0UpT7nXDadi2laoVPd/GQdWw6ysfkEeq7QBX5N1
MS5YvPMSTKoLl7v5Y8fGws0ozvW+VWIYrSZ3xMl0SwA=
`protect END_PROTECTED
