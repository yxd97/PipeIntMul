`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/1FuO+FuUk0S9R7h5GDhOd7cgw+nIfDDVGDM4JJgY00hlHUZme3RnwtkN/sSVEiU
tGB7akDVfWAWkPegpZ6wMlp1Ygs7bwOvDgZs5qO2/ZUVJkijugCsOj/LjZ40Oxhi
zdrDG83fTxIKVEzTLa1jvKCUKq2yRqbIB9KzlntDmtlZIK6eAodby0wsitvrH/jo
LQBGFybSH84blj6AJnMu0WG39lHzQXzIcT47+ww6f2I7VuowGsZ7VHaOWrNMYydg
KryJhgh4pPcnYqMqvUgBHxQkvy0l9WnxLXpYBBY21KlieoGFMV9b8AOI+VVEepRN
6U6M5O/DBdWWLxEqa/NXmnhCyrEwKoZiTVtOR4Z7cmCdLdqiL0pCr0W2NE9KmSda
Loa0+/jW/NTGo72B61lJu5oD1h5jo1Jr8dOW6dMxnfpnFVdUfG11gSs5+g00AApo
uRIucyotXxfxaNHzmzIcUjeIJWKFFpEz1siIjdk9L4WpoLFiSsjsjvKg9BzwNx4v
vqY2nNh/uOUfJtau8RvpuSO3c3jacSCQhCMN6gU23D1NhWh3TwiqTVjcUSsFar+j
ySMMdP7CQ/sAj5mmGvaEi2tFA7k/DB/IoJxtsbi7aPo0tughUuSTdItWv6T1hBiP
TlePnz7PoUFaFJmkc7mmxHjMAcbVtXue5XPj58vRckQO5fN4El4y1XOjchtWk3zA
XcELqiesCooPXTmAzFsJ9ggSe78cx4TK/q7sthFFOgcjcdWEaH4iWpDi0TRCMJwX
1UwXj57r4sMECFh48S+Cgw==
`protect END_PROTECTED
