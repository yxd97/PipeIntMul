`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMW83wSQjFAwbmNZAkctm5lQZAl0xs19IEE+n/aHFe8YBxcoNVZ1BuDUyuQvThS8
mgQUGr+LmpfltFKGRj2P+gCfgoUX254r0FX45JeEtMYrmZl83TdvEi5YFdnpAm5K
edW5mkyG4BGFNdDY+GLpi6DgyJlmpkpsxwOfFGhXpk6adbRq1DDPtZ7WxizHmO3d
satyg52gb2/zhhOH3TaM5BcFwytHviE3rcEoJF0bQQNi245nPbeFs1lNmzIzWIL5
9xNNhb3l5z/d+gNHYSobS0C11BM4BSNrU+sBxi+0aoW3qzXaoAalkVXsd+TPSuIi
Uy6t5JTkxxRgxIJmx1QAo9VVHd3bvdMxfdUayOfCZZIu+keIqRaR5A39qb9IyCta
1aVI8A/cTzwjLeGfNkHeviCw9t5ru+66+vDUfGnBvQeT3i+PV8KA0VM0kNoGOvDH
UtwVsZ8Ldhg9Ec1sjxH5pzn9yXeT+pCjlMxQ61pI37qK3QD4HMQvya2jQ3BfxxTC
rRID70g7AriHZ7Ub6sSq0MaKO0fJLPr2ZpvJoFopNGJDMbWiUtfDCpDy30KjDosB
knPW/piIdOsnHeQlpmfxe1DzN4ErDr9lMbxxJV5bJW278oQH2lY793ZjwZGbxGlS
E9VOmQSuLSVK77SUxnS9yRlvKkTUJDgqA3yRpSsF9G8yxyct6aeT1GQPL/gv/pwV
OGJ8ccrM0Pgij45bSmgqpg==
`protect END_PROTECTED
