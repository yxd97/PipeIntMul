`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BAHLywyoArdKzIgsqjCyjfZKWaqFzxNKyvOQL3dobKl30j3p22yW7zxyhOp6NApd
DTUxXxcD2pHQ40B3U8hVzje5NVlAeABpmcGUFtEWs+2/K4OCVCdWlQEJnRYdfV8I
keolW6Eqy4HL8PfTjj2xMFcm7Y5z/InMgbSInO+hZdzUrzI0nXfAI8MbBUdzNtvw
5IE7QF4Gu5Jb4+V9mlPMcB9ODUfnZ1803GFE3GZoNJOfGbl+apf8TVUunCK7dS37
RQlCagFF/1YITrkYeLV/8+DjxicqeSnjmU6pPp5xI0wR+1PZzN+aQEQoa2l+0UIV
7Ejxvuxl+KrkPzxINRJkWigx9Ih/Ap7HS5gfMRkQCuTzn7ngQmG9zAVscuSAHEfy
ql2TuO7bOo08NsRdH4RwhDl3bAVg+nyVb2ZLofxPHSM=
`protect END_PROTECTED
