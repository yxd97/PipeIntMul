`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YGuHWuNjv3vr1t3ORZ+oRTFWOXxdXUdFxvSfXxNhtA8zIudt8N0t7qCgDNwGZewJ
44SkJ0YLQEAnk8o9mTW9SW6AOE32EiILorVCrg4fA/ZaAKPWJP3EDtKCDJ6T5Ppf
9AplwU9DVoZltls1k6S4C1qFlTfPU8p+mcW+ayqPRg0vgl/f7rGRZi4YSPyDs/41
nKnDHSFij/OHRbOk5rw8YBqKOKh28v/5n3ph63X7sKa04Qt7JVjg5GlAj691ATSc
MB0qFWFDvuORclKDj6Z+ugnvJoZLD9OUrgJf0LS0+XLI4/jJ7NQy/y8m5Qsggegl
sAJ9T18NERQGOxsA+SqM2HXvAC4HUqk9D2OfAVMZAqM9h2qFOslop0fFSqrQgZR8
w1051pDYeo/MQDFl9Alu6Q==
`protect END_PROTECTED
