`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOTm60zfy6iWaY1Ww3unppKhnQ+r6YfhnXN5bUXYeDsOeQ05nfIbOLWvjd8IGk42
WBwcjVLCIt7KZb6dpdJvD7Ihm1sPqsjoVOwPVarpUPZ+9eEQdBBduvhPy1Sg1+f8
GSc5U8pE8gjw3pAlNRjQB9Hcix2ZxH4k5W5qzw+SnmOj2RKJBkYu73SPrpX0115/
1d+SA/IxKUP8E3cL1na8ZrA3xmwvAVS+1+0XaujrnjYnX2x+Hcmn6uJ7KN5/0HrC
Z2iWRAbWMXgoT7FCYiC5/v77EilLuaP2XTvrGpP4Yt5PBVVT6wCaAcA/AK7oCX26
135Zd+WwGyQ/RCYFZ73V1H4PHMXXMWVD74M+gzqz1jHiUm3rn3pvfFfHY2VtQGgC
juQBkA0AltU3C6FKY22hSjRx3qYlwL6QhTkzTaLyPi10FRdftW/C2lDw3WgJA5G8
u6V2z6OcnPbGlANE/gzP25SECfiodohJfNMzAiiQ/60LZwQNMs3jIe+TRnrlVfVM
SL2XMs/Hmf6nUzOFjF99+FgRqTCR5nOA0KWv9L+NR08Y/dQqTX2t9y0I21Rtoigv
iOorvWI5MmoJYzjhzM4HHfbStwVpY7WKD+SDOMCTsXp9Gla7yE+bOzCh9Xyp+GiD
78rFBDwOK/utW5+0kucIlrzAxtMKq52M7gJlGDnHmeztfuUp1eL0dEAS8X8nlaKp
8UxjJ6CoDLzgKErvGeWNRteG8D/Lnv3le4frFXAwQM5XoLKa2lvnrB5U0VpqgZA2
kFfjRoAdzHmUUw960YGcjWLzwMi2eavBsCNXPpfJYyMSL0HzY3biS6C2uwupxtOT
u+MJAOzHPerCARnl0AYmAVvOTNmyJ29Ka3eOx4/fkkc3Vh/gN7ZnkeAThsV4Fk8Q
BpeRrpyJFPsus3Xznbj2LfrOQM5Ydd6S0W3OqB4/j79v/B2rUnnnhFq62LGTS/Lp
yYXcETFtBoJzFypPyFSxQizoWlSaLeIL4AIV/J0Rv0CgoIbs0UkfIUuRWFf20LMC
`protect END_PROTECTED
