`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1tvdQGZ9+qn6ZdNK+2aucX7j7byKwOuW4EN0DRRoPThwquYfzIHc25rNz9TLq/SP
ZgppPyO3/0r1EFy04iW2BoW0STJPDn59OkrDeqgqkyrncN5zv9WzggV4dq5JS9nS
VeCaKKWLLGpR6HoBctIIT/B45laEcRLqApEOmUnTXolTImepDIZ8Q8ZYeqOMVoRg
uqC4CV1PLvOH+ynCkJjBFbqadIc6EiB2F9W3YRJw+tfMORDxh+6VXuj/sXAgzTzp
1Rnfw/IjCGHApnibesW6TQ==
`protect END_PROTECTED
