`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SmG+eJsfWQNx/lUfRbJQ+Qv3vOVtT26kwR6HX3UoV3Hh3jO5mUhBM209Sk2mZdj5
ml/MyVxIlpR5LqWSzgOkSgs7/K+RyLrE0oR6B2G0UvBplAwFn1G+nuOJLgG+gd5y
8MsZpbmCWS3sJwchfF13AbuTyzvmOnbVzr0RDRRRjCPl1rCBFx98I69l+AtDFx98
jxYdvesW2kTD8XEAXMQ+EyF2vmrB8dpBa6nBybwIafOAbkAfbV4q71DJuVe7KjY6
+xJlFGDL9JPi1JA8iVeGnqFh+9D0qnpCdDEdTF0STHSgTqZ5N82s2zK8okSw/quY
8qC8FMWuMBfIqdVVKxYYEeoL5DpoeW12NpSXAgKXQsUb7uf2oRNnBakjd30y/h15
KavV0AzyOvarC+lFmIo5Y6eM6DsPnsCe3pvWEEjgP1N3rVgQH365H0rODIaXmfe5
UDgwyEpeS8mO5mnDmf5I4WkAKbMrXePmkQkHGFKVFmxwm6wTCRUsO8nl1w2Okp3N
gFqg6atay1E/wS9hyd4O6MaVSVV/QSjTmbAY5qVg4BCj3mwaHHWNlR56myUABSpr
E78pRu4CyraLfuoG5+WrXRgnM7N80dep8TlA6/N9u7ynympO5umdu0B60uoBCc7q
2PvVD41QH7ig8x6Q/vjwFArbH5GgfFgbMpOGCSjjycaqD8+SkXu4Y9HZlMf4TACM
vlN/+11xNTDPpEJVkWx72w==
`protect END_PROTECTED
