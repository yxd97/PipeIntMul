`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5tB95mfXtxjBU4g8LtwYxVaTrsqBHeKm9y6Xo6kOc/AdTyT2DbltIzpsijj7tlAc
S2+8YUoz6kJiBZN9N786Yc4bRa8TIsdE6pSfvWKX0kBNsoSB4pQplzg+Agpj9qkF
ldThC3TT+Mr4nuzty6G57qJexGARaMDfeL0h2UIqeVRyyvamrm/NkTah5A0n0JJl
jsCE7t+VBptvr24BrtJ/fHiyzP3vJysU9RY/g763tLrK7lvDfghiLgnLRjpk9kUM
70AZgECAzfUgvGj+r8wwKXGVuHuIfb+gRZ8u1Lgn9o5irgS0dR4QfVLeAE8z2Adg
8Tm4SGrzj8UKLSpdNbPW4M/JcDFbr1Y1X7f9BbsFo10fG0qECLbF4n4bdwtU/fQm
LzXF7V6KkBGSnLbSBEuoREBDWjYToW8uUHDW+Rozj5bCXIELo+TbABNemlL2miOr
hBi3oDD97vZ3lhuCjhfoNl4hcxunHx5E8lmlxnpgDpUEjIuXfbkOfThxIaumcw6I
I1uYOVE+QR4Zi+le/oUF/7YXVmeGkvHKNu6JEw7fiFiyCHSjh9SOTTEFcXyLSBle
cIgHHmzjnIjDWpc4jfvM4fp2LaHJAhkv30E1RR0Oo58lVpxQ1VcTNcK+jjUUmS7A
em/7EEsshqy8/JMNqnqqYXdKqTNZbGKEPsfUw+8s60urUQ4x+OoWmvQCDoh9aiB1
icZxu8e9fgXAfP4flStT0lUq3TWG1olRYtCmrdduijv2vv7XQc3YqzVAPtNz3phk
9kT15s3aHdRuSqXwaIVvO30PfvzF1J7nLuZ1ltDheiZMhyYHJz3Ko9c7nG3o1iAC
3LF6Q0Iou+HlkkP0pex3UR2XO5jocmrVLLuKMdr3qF84Zk6zLsNcfGtnywDpSYNa
RuIaZGttzXny9tE01sVoW4SMFIxc2a3fQdXHCuz191vSIjlNbo4gxqVnThyUByPo
NpvDgglx/CP+1UUTb8zHWUUU2RnO7lbzCIj9ev0UqCddmcL+dvmGr1k2s33bvPMe
3phs0NWUXcIQjalCy6GNag==
`protect END_PROTECTED
