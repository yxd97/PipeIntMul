`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7Y5PzvcPZ0A/gPHDSLiZeoBpzdCLUchPuDvOMXcasA88mO3qkebXByNcg7UmgO0
8yCtY/IRyKGr6b/PfuhhLEnSEV1gj3MZPwwBQ8s8jHRvaOsUFkp3Zl4Cnq92lBpT
n8ZuMXB+j1xA2Q2AhuqbGvuX6eSBZmHo8rncHw1ladlO1WqUL9YMxpWjPiT0E815
zWJMDn6M4+TPKQOt3FAztLnjY7p6O9jDCn9NJP09jsxofHvDDkva5boeD5jfOmuO
zkV/zHQxqvHr2KMCi9r/sPEmfFph6+oIj5/CIySdUYvNtfjqQW1CzMoXVH6iilkA
//xpYlPKApzCOm7d8TZp/2QR+wUVG3kpqqxOYo4kQIv/oc0fu9SIzze5IypbGCkk
qrCT5+DC1N+52Skw+vypBkQKLz+iUKsaA0vDqfPnW9uG8wEGu6eEPMUP6NMFFSTh
A4/L1usEVXAgSktqbEojToskZ8CBx9LFFjP78tvC043BAacoNmtoHHR60IEnzU8b
mSgC1qXNGIiLLTunHoZQ84zLc1w4zBr0VBwYKdE3aOcMWbOlae2MqL76REU/Z9Mv
w6a2uBXQpq4BmpibVmx3fjacKIb+kCeS3dZnwQDgMHVPR/qQSGt9x5IZOXx6OjVC
nNlsGv95YUxIBFGcCOreJ0gjv/x6jdOJNa/KAjBlH3axJ5EfnpNS6sbB6icopujH
OJOMPMLSVFnSvfOOTFmpECWllnGfhXQyjOWoBewXt05zn8ocpVHVG10RaJdTyocb
2fJuU8uZyNhKMBNggdbS5akV2iUGjEWSzmuvMIGy4e2HfZ+O96OTTn8TzYd3lZ3I
eTCnYB/WRDvAITtbhQxOE8ChjcKaD1kIp9QldhfEk5PfdcX/VU2lhBIJunIWtO4I
TaqzVXC+XIuVfUFmpthZDQG1A9gY/OzmU1Hqp/lI2n8G1KWhNPAX9ZqSZvluo4KR
lCe7UhfyVAFrfuRTUYp6maTXoCfts3TUov0mmwnmJGFanSet+oSf7oFdAun+EhG3
okenss27sfqByGFJTReUXRicxPZSDL5RrXRIHsdTznp6B9jfz+Mpq6BRPZaqGa4s
Re4bGHF9LfAPra1w9f7Ul3/kibwb6kisluImYbUo7/rfmUh/DWG/zOZs0dB3slu4
P8P5XG7Ctjg+VdcKVx09nguQpIgSjwySIoseyLhRcRodCkQSpxMrbmE+7Nthpxr/
mAG5UKs5+npkkuFEchzPiEQ+vEfRYoOtm9KuP498iMVGoNIDuj6cGaiwoSXd3O8j
dqFaNFX75sugq5Qm5zyAo884k1mBub8IN/o0NwpykziaAdioh7CLNd7YAKNQPC6G
voNDNZ+hksv7cRZfJ6ujjwsoMQPkkx1hGbwPgMXliQZTV6Q+e2oDFHlhw69p5FmJ
`protect END_PROTECTED
