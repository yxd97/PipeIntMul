`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VzQcX0PnMPKn8f5KF+viipxdk8n4fi679kuq3Ey88psdG0Xj2h/4lgc8rnpvB6sf
3TrGDNxlUMWeoP8T1nZrN42HsG86Dqwb2aW/o9UJTcwZQroSYGwGlhyRYxQogt0H
pBBNru9lOXv2l7y/ptjYWEkrt7pwivJQIcHBkpH9No7+s+kc62RjjJbbdjvIHbdz
HnIw/hiRmAHNRwhAQYx0vSaP1AB9RFade7VkwhJZUoA5l6hb97Az5iWcyrZS3Yjj
SlSP7KOh8cAKmcfvfeH+9RkjgvwrBjIa+KWPpb1oxrKafby/yEFdksq1LXJC9Hph
6u2T6upfi50AXkKmtt5Yde6hfukNiCPcz6WD1Cc7UGCSSicvEzhoCMrC2+75JC3r
BAdFR/utQz7Lk+WbAwzGDG2EBwSmnPx0T4gT9vJKJxpxINOzdxe1rA7fEZUPSE0e
`protect END_PROTECTED
