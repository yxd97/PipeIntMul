`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VvVw/2/5MjWeKds0GY4s0Soa3C3X5r+S1V9v2w1qIEqm0EAxoXXhcy/CgOoq9dAD
OJkGCm2AY5n01gj04IGfEpO2o1htxswyoWYIdBYAGbaw0vkiZOwnvjHQM8Cj8pl0
rIGaKmpwt9zYkyYUd0T+fYX4WzivzhubOljdIKCu3U/nqRJeEV1PaClBVBMNb0Mt
Njs+Q8/oHo/UqmkyJxcWgAtTKjez7obZC1I4gO1vjRvmv0ymBIwqQeHDRvRHTl0J
ZxKuDwqvrrf+7rn4KVQqYeksucDjmdkACV+dnZneO5mT/kw5Efasyj2JI0FD2fnL
R2qFUuYeN8veRBJ5xnfF6BCVFWQPSAHhedtl5C7xm5j5vQWLBQOdpdle+Y28ad0G
dQtddAPTqondcyipfYiXwbk1yYmzoXDXL1dt9h86Q+21ovk9dF7YjOgNhjFmY+dr
Z/P6hcJFx2nJE91WooiOjBQfUPk2zzv+IzgbZ0q2Osw=
`protect END_PROTECTED
