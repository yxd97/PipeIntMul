`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lH5IAotVB6Jl+BCoy4SgZBOGAq+AOrNpob3x+zTFfNE67EJGhqaICHjWTHuzZTy
XrMWBGFMOyIexQsOSdJJprdWs2pHtmNgS9WcB5CmKtQ96dP28GuE0o/+T5HdJHlf
NQf+VeFPemKt8i7ySA1NmXZ1buBkFIVDRnxAAO9sAXaXmlG5WuIkV9BaLQWmPKOp
OvaZjPOih+f2RQoNDm38xtWKmZXsZb1bxcNb/P6jzEivuZcXfsCqAzwo5llAkbDh
nelSs7SNSXyk8cyqkKJLfKmR+bAB4uD6pIQBLZE5S580EIiQPAhstWC1XU9Sw1ew
KAp/ILlNAQeYeI0vTSt5IfnLFSticWbHjcaahxRaDdXvKHgzqWchml454yVgRn0Z
CBWiCSfnHDyOp2vE8ChLwocFZmGx4qf3rigl3Owc7rJ/41GlG1VmhLvTbFxg9LQo
tSAbL1Uukr7WFuoeNrxBSrcCGinXjC4Ub0GlK3vSAL6ZMwY0bOC4EVJavpcxOMi6
8RiA6hHHQorOLsgg0DLTGvQeegEhewD/2eF3tZnByfW2C5XB+ZOVsQbrzxVUbTov
xrAetjC2Wi+mhnagpucZkw==
`protect END_PROTECTED
