`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VFptxEznX+tiyLX/52Tvo/yrAqzqQmQcfp6MqhjmPfK37UiFQshUGQ8iAS3TwaUS
ZkLeLirpxVym/WOgrO/+koF1q+tBPhSirok4DDKB8/hPuVyggZqRPZwnVnYEoCZn
4rhkSEFdio9PbWgH4BKec9ozD2vBqtGat3zQuFrj6wyGTZUTi02SH1TcnrL5FDw5
DvhqdaAVaza332SCUgdxxuIXONuyg8P8I1kNQMhu5Dor+ukA+uHDrpaUu2fCe09X
7Ev5+aqr1shU49v5qvpvb4v5KI9mDKTHzYqpJLN+w4aBxy05JPH53ub1bLMVW42P
rLrzcVw/a0fRw15CvWaLEGhf3fL7sI0AxlmO1pvEOwfkPA7JL/wMc7Cyp+n8j0Da
kwf+u6Jvk/I2Drgsde74ZIBgSYE9y1h0YiTlnbbM2XqNHbTD2rnEKbHqEnIIVyS3
JCYbs5USlAL/LXR1dY24jn6G4SBCjXPKinQ2bg4gea2Q+ymPqJBK2rT+0/ZomIZD
WvfSlJqMcMC0KnYZvPki1xoC+td2wpA2ig6MJM1mJ3ng8/Zmyc0/2DsJKvghHAsX
Fn9hH+If8Lx6PbhY72cIDdpg/vv0mSk8MpGrGyiBX3AWvnKNI+aJLF1lffC6cd95
uZv68YEfUw+eswhTc5DlyWt6UAH26KV48DHYavnXdGjmTraqtBGrujNCORJXVEwT
GOC3f8bAu+B5ormEuB25mGBspA0W7MEnDCptKIdkMzY574zLDbSddY+TZtKPdHHA
to+R1vamABLX36py8Iw+l+9wkvzGeeAL1m2QzdHMw9oQ8WaF3F3xqoWBmx4sP8HC
pGsnukoK0TrfUlHklmfOdbG/Yurm5yzHWeW6L/a3Xd+yXW3++CjRvnMOKfmQ2/OS
7XYviyq+kkV96oYkFoNWxNdgGUzEcL2zdpvGOYq/hBt0y3Rm5QShC8c5rheZ7DhW
ucFxSOmME73RkFwK/zFrAKAkYlqwXE7CQaObG+maKwrZ/53xK+iAsh8R+v6tTgsk
iCnwNwSBNaF26mQsOqitixSqgRsxCgcn7BZa4ipWTMC3qGrUl7eYRRoBfObOsqm/
RMNGeJXpzoMmW1JmZc4lmihoe5gUfYuKMTAdRwZavuvMWa44XG4OjCamY9fUQBN5
+CJQRnOyB0XahxgQ1WsJagGOkksLsnKMoXC3leUS0PTtQgxWZdZQ3Qe7/jNk8v3W
vJVjjxvnSUoKGRfVG2hpT1wAbBLEpH95K/IL/mWYQa1LiWYaS0P5iR405GIFEpMQ
t5O6YXzzacNInFn3N3/4ZNBaRJ9SFxGlhJAqVI9kqqD1rc96AwON3yP9/dw4k3lB
oZdeDogS2mOTaGpRidIAtkyU48s5pfceKASWbezsRxR1Mw8ZDecVvhfiXLAIaPRK
XC6mbccTEi0lPk2+QVzAFzP8pfz2zeMFAZf378zPCzWdzKMA3RqD57WmkZ8C+JIp
Rj6qACF0j/LZZTwMsAfYpnxniLMYi34pxeuzVu4mIVPbIgouBE7L3eE7faCgElS4
NdQRRFEoWyo9H88ZyoosWrL6YByxHRHwnkTM3DD+7QIz+fv0y5mmql9LKoJnZpK7
qdbaqH72KonYNrD1nHpddp7YedRlC+HPWuG8hRpuSiQV6tsaY6ErXkkLRA5ikMBf
waKOVA3sAHMqgm3aXkJPjhVorIPfjEDcw2jx4vQezqplG2l6CrRs5j3i6LVMjOGQ
5M6oukHzM6ItcdKUTMLqucFcwsoIdi/2UyNEq+f6T4iBkxRnl797LjAwxodaOn2a
wbJgmhXMbN0qeYdwr9yR7vuQZ0/l1kh2pOvWk5DxhXAbOmVG9tUwocL8PMrIxmJT
Y2/T4dFBzaXQ/GorqEgaHhCDhzjJeJUqhvtERZfiBZjSAKHKKNl4+DcToQy++Cvi
lzFvB3aRuKDQOfYAtJDZHg==
`protect END_PROTECTED
