`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PzUUmHOYNLZsjNsZSDgfTyrw+qsAZyTsHvYovv0BR2ReVWSm1bJaiYAHPXu3msPy
0gEThTs/cM7NJq1Jcf8J1nu2nDFhjzLOpdGbZsmHZfLE7NiBrcqIfMYVWtQCzMlu
2kEl0JKaoMcFGbsq/JVAWNBbOw8n1HQA7654aQs0x+doz/qgqlPSzgOj5QdyS/bq
PV2n1fnifymPhEWsu+sEu6OnzT8q7FhEJkLt15g7h18YTNTYhOl8O7791B0Pdyqi
OhBAU20LcAh8EK4WHvDln/BoI/QK0g5tsSy3/lHv2DE7frcXW9esaNM8eDOwZ3Gl
hvJzCU6kHCh/WhQrpmZxsngGa6XC8Bnnb+A78ApgaEKR/vP4ELN1kurbp/wycezq
i+GrwPu1/tfmSg4hrgGwKg==
`protect END_PROTECTED
