`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KJRcUL4V08h1DRohUU3F0KnZVMEE5oPDi6VVb2P/bNId1tkYh56WPijgmxK3eZ8
VJ9hRNUoHVyLZ7Neyx9Om+qA6EhGtJoMWhhMuxy6bpc/yPu6+w2x5yNhjiPdR4Mo
S/rl6RYtj090I2iJzHlq+ptKftlWHj6i8VnLvNmXVGQOH9VRpZ4/1NeDlnSsQsiN
/c4DFwzOv99Qx4+a6DMdF1AyhsREJdWNrZt7snFlAlPV37Emam8rbP0gmyNAUJi8
uoVmqZuEBiLcm0VADxSfWKEbtqpZbLusBOxXCqFDUZijUwo9EZ93/5Hsq/EyHyLw
lg0d5elmtmoTcV4OoHw9SxrgmALxOcvSB1JkmJByac7UVeWUictGfUaANP02d5Yz
q6wh82macS2fWcETNNH3F74Bo5/m7qYddnvnAcFAR5fQhiHwWMbge3sTxpp9OvOn
n+iZLAoqBL5aFcBCBNgc+TKJEWj/OqzU3HG5N2vdeqtSJ0VoNLq++Viv6lZT6C1o
cAo272bMeWHNXSoYJMD/QTbtDiMB+m6B4UVuuwyeOcuVxaPI9xQEWA0lvcfB63My
6tNGqMqFy79Kg+KpelGbF81UzLJgWPH6Z3H1MvOA42QB6eyWWwtZYls+dgJ7WKiL
NzWh2vvnap8amhR41v95n4OHxpB8+dANsakErieh2kCD/X/3AZf/qYhWx6G1tXNE
UrmdtOpinW3BDoqXa9heTV6rUnERlYrkjaVOWP9ACKczuwSE5pBHbBTWbq9jzhOM
sVTCq7exdokwvz5slnG9eYx3uYZd0CRsXLfwu75rPA+6grz7tpw7Slu4DUImQvrq
tO8oZ+jFegIywuTLKapUYA3/bVSdDXohCXHSoCFOwK9/1VKP6D4MQJ81fw9fjWWT
kTP4ScuL7gtDOs662EritkGb5fXusKr15l/FCcCXoJ/6bzci5Dw+9WLoo3y4nP0y
Ij6RA55i56gUZYGhlGKlF12ysPBOcjVyRDVGzCcztjMtf8s2UW72NRh4fbJoIjQO
bMb62qUs2Z7xAdDXzkGpYuxGQI3bwKiaG1r5EPODrwc=
`protect END_PROTECTED
