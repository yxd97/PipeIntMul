`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xChzTn+sBmie5W/PJnxAUdWueXRvkS9WpwOqjlU1l+jOhS6Z2zUI6DF2ciecT2pf
dVQZLaDzfGxKFWHJ/WOsVF0x7VEBwR56KkcnkakemCixkz502vzyquObCEEYsC7Z
nTDMV2kgNJvmIne5wqurc3b3tQ1k4BM1y5GibyFV1S7KMKAeVs8rfR2QMVsGsL9O
Feo2P00s7rSo3NX3imhQVDinsLEIclv4jBHt9ujF8ble+cYxuXZOa0Bv0+OCfQXw
SdVj6zE717I7Pgqa+ijQ/AgG+cn3/kZR+7el1R5QlYoNDhNr8K3W5anLDOwgVfa7
XkVQ7m8PWYtzTQKy24ZUneXIbhHNKQThWMwf+IqRfu/adXqb89Ye2iqM1zrG0p6n
rEA4A/pjPf76EiVyQzif+BThlN9WG0K9jtwKOAucpvm+ALnJNRzI/JUHBvOaswNO
`protect END_PROTECTED
