`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2/Uo45O6JFHJEIhddSaiiMVU5mhP3BZJLnQH/mTSlgbzkU7ycqvCKrrQp31gxMY
VnW1V/bx18r4rPMhQ0nNSNonO9ZY9jlCzaIGPT+LZabEmCipl1dJ69xKDq485EkM
Yhi1YvGIA1MgTAeRoeBZXPhhMv9HUnhAcQ3cR4c48KoDfI0jqyL6UIcrex40lRng
X3O8jZ50d8aj5qN0th2/qxMlnTXCOj7hHrOQE3KLq8RGairo8TH+nbwg3T5piP9P
ZIh1NsbAjmyyU4BeUfYiiAUFaWwXkf0D8ZZfXmhZq6BiZG6VLKQdQXjRVu9s4rqe
uMPkntcqvwxrhjwCbnZ7icG5IZTUZqmUtiOmNRyrIHJ0g6gJ8GnkiEH8YIWhdF3R
dRnKjgjziOIvaUKwHtvoIEGSCKLmkKWLAPcPsJckLYVkw/91xhJf4Bp/3w/x/I2z
o6NdwGm1oYi6gcHWQWhz9pvW+QrXfyNIWdGfjwYlT4g=
`protect END_PROTECTED
