`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjBupirHiyCRLvsbo+cgMEgpzBhIhndgftrdbPRClCZmUSeAY3iOqMAvXM0ft3UB
cLHuOoF+bGSfVS7y5UBI3s+GWX28c2es0sKj+Ut0wfx9fiHBlzQgDWWGnniFoCCJ
Q7UNxGSrgwpzirnx88j2lHSFdVtJmlewPqdEWG/cqcqg9dAxFhicR5LKsdVEUUOV
Hv+hwgn/8GlpVHxB5P2JF4LgiXjfPtJ+Hhs8M5pKKao1ojg1IkTRWbG+Z4QbV4Fo
oP6nYOSn+gaAZOoTWyjXYebwdvW3ntYH4Sxf8s1JFLBHZ4H6ObCuARxjil4CCvR8
6UNjB2WOoy+SZDnfvA5I/Qv6VUNfPU1/G6aP6/lMfP5ueYTkU0F35aS+gwlJvIqv
EqNMpXNV872qj0Ap1bkSQMD0cE1XjZyj73wulRogIt9K2GZHH3e28i6JI+DlZvVP
`protect END_PROTECTED
