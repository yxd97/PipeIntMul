`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L1q2CEgTNNN6cFlSQWeIBotrWroIVqKQRgcyIJPohLMYOBQkETFdQZ2Uzn3Zsx05
loBa7PyfYS5FaOdzKZQe3zotP5OWz4Uo+2JBgTV0zczUyOfHFSQZAaRo0/zHfO00
MWbVp3erF0uAC7AvDYbbU+dcrMPZi/IaFJIDoCqEv+OH93TkgN285E8Sm5Lx6Gt5
AB/2G3zF+btzdZHkMMR0K9oV5DyfAMK1eib/Zjm75NDmlMeBXNe99cbEy62iXSa3
eusDjil9cBsP7cG3MSN+qzpPqSZtZ9rbrHRD0V+wn1iqnUbIwmf9ZvYzqMheb81U
nsD9Y15IF2F09LZY+A0+d2aMUv2J+VQuqREM7t5gaix20n+k3PNHRH2csT7N5nrm
iYJPkXMeG43khBI/N/FzoCfIZB7HvOiZ2WhZogT5kBgTihVoN3b9N+t468th1rET
2rXdSai858DqzI6YvkhgUeursfQ+BvSsLHgabhry1nkqAaqwIr7Ex2BqOffp6n4n
F1Us+efYXf+avbQVZFczdha/knEWKR567xetn4cB7SoGqi4efNjJfJApcrIRIg24
x7PmGqOXpJcqo+wXHXaLvucIdeOl5pcD8DCUo0VJww0GEc5pqMkyPM0kVP+7ZqUm
trnUMxVmoXEZAKzAkxLvpysTdaLQbN00hQCnfr3pfou6arODpZ7w5TIbTxdKSZSg
TucMN2bn9SPTVZF+mEX+h8u8MF4e8iJu87WBzVwN4e+ic2fOlke9RYilLubw9zQh
v3qvhX+tHqKfHHDWbhkXuM6+9jyXJsTzLDospvDma/HrSeAh3VfXDTpw3+x7iDFJ
ifHKkLPLaS63evrprn8hbdeqRE1M1BPDtA4GDUZ58VoPp6ikcwpZFgCSLKW6RJi8
aZ0WzKFiwiVAkbyh0rQkqNhMp680KTGuQrFZhOP4+t1lywl+WlJD2bgW5S8HXzA+
MibstHIQoK4S4B4Ziq5auhfRm1HFuUkQtSy7eEq6VieoXp+f+3BYSU0S9A0OgDmC
cOICuYRU1xHNLkLKfhr8GsVEpZKndsSKSkMZOyXa9ro1z2ddcJrJjupFnUTxURco
zC0ORRj+10S+3sHFAfODQ382c84nVupILXGIh2Ed/IOejiu1zhRH/woZpDv29net
ruyTYheJvTn2CMGPNH3v4G5bm+Fs/k7W0BoKV/EAekfKQ0knObwwQ4RJNExNwE3Y
gdlP5eKEmaiyFG0yxMe5IPNwqTHjGk5YT6EWMi32GDZRRxyrum09KQqcx60Irhrh
P2BUt52VlviWRW1/OzPZBQMZ1KR2a37lzQ9BFZ77eRZl5qFRWqWy9QppkFAyj8Tg
ohoX6CC5YnztoZiV+nUAjXtMPbFqbuFpShoket1SjrRgwHch82x6FsFqpN3XnrtW
aY8qL5J4EyOxAd0KfoPfyDDzo65UQ3pdjm+QUbQ6m5R6cTPtoCPkqkIKZ0UD3fAo
rY70L1QTbC3NSTjOsxqv6X+urEhetfJquImzTrrDT5ZKPvMJIcVJ54HrwS7Qbf9q
I2N7K/eAjqUuOXhprOfOXFWO/65JiYd8UfTXP8HKOV2bJPxq241/Y+qAqSUOo4jP
0xGBVqLNvFHRnRH7aXbCmS4/OQaxUYXGRgsLLmPccPtq0HuU004zwALh6J/aNBr2
CL4j7ECuDfODlKU5JvZ446dPom0IOGzjAKrUGWqyj8wtmFGFgwWh/FlNqFbPzmX5
VMWVUAbJFqe6AGQsci6m50DNqNFW9eSS4DKQ09ieRBdCR2IuVWqSijMXTIdbTAVi
Bof7rHStSM6Duvx4i4ZcjVkKdQZNIy3YfjNtGiUZMiN+u6iuEwFYk14vxVOqtUqO
FzIIbv0ag2+ScbQi2Pew2pkdf68k1FFQofY/gDhp0wSbDg1bsw+oms5MTzYI7tx2
PQtgy9P30hzUdoEHQ/l5b3/oiRZpPFffYrksSGgfDa5xKcvT1qyc20tHT47xhdt1
YBsmLLch7PkUz1Kx/ap7VOb18jboXW4zMtCHsylshif97wicFfRB+XiBqFUeTHsX
jJdkMZsmIInL291lyTLPZfBJm/75uHtDrbw0XD2NtPpUgMfZJoCO89VPXeALeHbZ
W0qOnsGrLBsU11K+NmlAhI3DJ8Mz6W0ShC8ek/LwhLe92YaMCXreofRCxcgUtzKh
FNevFDKxR6HiIM8o2OSWtrfclNxCvRcws3RTdFo8a3DZ7/X3+5agiA053iWAaeKV
bCtj9/1yXY6ijgGeZwZJCQTKwLTjD/i/cXjCggbuAS2djFBFNm1ApQDOGie/dTox
f5tdOlX5KysJKs5FgXJe613XhaXnY9oUU1wTUtIBF/Qnq0jMQ7yeThhL3kX4s/NR
ResJQYBVqufNtsXao1fmkMfr3aaE/AfqNSts3b4LIXkE3cTcSajsQ/QHcSLwMtTD
1iATQhPUcPWKkIxg3Go7wN6Vdqklj5M+5n26E3BBBmp1r7m2mlyWm4H2oGr+39mZ
LyKvz9+bUifL3kglYX5pMOuB9VgEGdYvB3G6XVaFTbpZZoNaxSqFQ1FZ8iTafDAZ
jbDwI1FaqpOj8/GwkGjASFpL46KRK2Y7L9sip4wdqQBUvzUrh5xuiFGsdndzZk1O
faQmPlqp7Vrq5NY5kK2F68CiNg/pwBwpKPkSR03gvUGzP5yarbOu1MQrKRBbSYSG
EwXLyNhqtEf4bPDM52d686fBZaB2M9dTO77PXrQmYrBG82PH2zU4wQ5xu5+BeYZN
TItVGgUFDgEKzrfQTFwjQ3kFr09KItWyFEfNDmbvfegDD+zN9JjQAXS5JuGexpjZ
BCkxjCm7pa4dy4YHdbP4AYnXXHXiDdD3bOGeT1yOCHttLknR0GRcB51sAaBfXBVF
FEEvJB4J6CzlpWtnmLidWJHNhxQbXCjYRDfirxJu6en54pqQvxQLbM+hx5UgiepG
o/FoBphyIHlE2rJuzxrGpQChnlSBGVvDcJ+yoZbrHCALzvgswlt+Ffiyydnh2jL9
WYpPgxdsw7q7aNrhoyTOE8QLXhbGWIoKRLdnbORyLydVEyRJRTKs1akH3FrxP3h7
mNzBNSyFxtqxzftGBwTjqcdX+gY19kSWx1WrR0xORda8pFDgtIbH51KhlUwe6nqX
S9QXMvAtKgh2wkmJ/ZdU9LgbzxhyV5jKEnMTu9sOiy+wPVKA0LW4Q+hnAJHbY1y9
1ijE6KejO1gEDh0aOxqG/0qTZ4J1E1NT4fBA2bT9I+lh/DJV+x3ju7G1wXqnyhDq
qYbQxQ2wW4vZGGq9JIbOU2z2HiHARmsj1GAwojoyqwHawsZYxwG0GoK2HIJlwko1
pdTRRRQ1v3cS+LVJFaYuFt6f2140KnGUkSQVQeBQNZE59Zj8arQIarlNk0J71CIM
E6ARd9vdc8gk60gf5ymZbxjYjlwnpc2reQN4KhGeC93ClNc+8BnFPtBWTejweTvD
sEGjKRplPTbZPj347vXM3twlpcoBFn2GeS7S0k9WNW+QXhzoFfecRVwbbnfLMS3R
8Z0GdbuF2rmM1RySQri3YTyxWHjMLIPaoSenJvcOR6rZzW3f+9XYU4Bu89w4v4f5
TBzX7A9MALooCmdR3187sUdISXbz+8NWW4PYmmrtbSnALsGgksuBABf1Qv3+SkFn
WZ/iv3A4Fz+t6/iG2NUo5OEnM1qiG7EoeM1bnnaZ5YfyX3l0X6iPa5M3+ckrcF3f
zCy5JWZR7aoTR2UxC6c4YoxcXjN2qtQhZOpho7rqmuIYGHkzARm3ujl9IuGT+Qsk
IflyVst4rrvMe4u2o0PCNch2BZcRP503wvm05p6Zr9x2FJ8YglZk3lfVm5tHMrmj
BV2vTBWKDLvg2Cwn5XxR6j3FhX9ltKdS6YZ4CWJ/Y7qszL8SyrygxiiG/nNHT6Hf
8oIWcT1279vPquo7qCNK//91d1YKYeg/Fzr2sCMgjFxj/dM8JpR48zDhVrC+5ZOy
xGfH6MqbOQSmDbQH3HkJrSxbTimRqCj+TT+yc4nCqslRUpB4xedn0r2q7xerCzXq
4gioQc9FYJQRyykDrI+YTQEhenF5QtTBBR8G5X1Q2y6RBwbO4ycl+1d9RWcLsH2I
0APSWXcez2yCiqpO4DtrRe/j/jSSQtxSg7Rbpw3+/jy8gfFVvsZ8E9r3azscd1P7
4vpssjIcouZ8GPuH7tW7u6kRXsL62EXfG6MXQUK86D8fnpzJNTDG/UdCG55ItWBu
tu14Y4d/Hg4b2dyCKPG3G+Jm4uGPOiBK70dQF1ds4wGUWJZpjcmtSD4xNUHDs5gj
0dsWF9tlnM8PVW0dIxPD5cCDXMfdno61eAKLIKtnYMv0bNskMLQl14PQtpaM14P3
6t4dWhmeNWQAsU5QLNw0VUG7iAc+D7F64hBOHBpGwGBopkbrbjzcWW2OOlP2bfPv
O8nZ7Bd6d+onaDy8j0cGjEp8qVfulDz6gfyien/0YHYqlZzRDVKjM9G8qMEy887g
TFiPzIOsK+//ZrCdR8zT5lJzn5PGzy/JIBeGyW1a4YRshMHtX/jIlyLzk3YfXPdY
nilWcJJF0bN45ViVQP3ZqHQpp4pjphimRDVj+Cq8DdC3N92E/tbpaY+fwBp/olOE
y1i3hesOu+i+EhhE81eb6wQyKc8aWDtsMu2S8q66W2hSzuv+B76d670GNbEnKN2f
dMziGCjwBabV0uUiSl0qZU1hl0dYo5D+ZDcSv0pk5Vpd6V4eJJOHsrQlu1Xw55OU
SCgg1RJrdXklLVppGTl1xvGVOP3V52Ph849wo6awI9LGA9zpGrRwFRLNzqpkllm8
NJ/dP1FUof8XH7J0gWPSeSfiZJoA/KuyRLfet7J8boNzEnRuon0Pgw2DhBPyn+iO
ByAYbmoc/0+4nezcN29+AoMKLy3sGGUaxNTHhC3UpH4=
`protect END_PROTECTED
