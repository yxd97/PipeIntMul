`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83Ua/tdkgFMd8/kKqWxcgRZ5Pcy7LFPROq7aSo5eBzwIi8zpV3VlqADibE1N3Uo5
F5fw6ovF1jaDHFFR+p5TwnyPzWsXOsa8FMJL7zGdFPgsoTBVh787TsYIcXm1PjvE
hyDOKGqa5kURu9GuiM8xtnmzEXG8gUJouY1irHviSPBaEbQ8Oaats1p8DDJQBkx4
DDzpGzT6kDqJgo/J1787wWpsBxwSAfLyxrEgs6E2Qe9KuC/RY9SOSlj8fOkX5xQe
adeUXwiv1wUZJ32D+9m5z546UPz7NJTLETyNXwevEDLPp4bpXsww8jYWPMejBWPv
+GY2y4kjmnFgUqYd2AhsUSxbgHSYJrDTMxedCEUn5Q0UiT2ebKwvwxkYhd4DTVa2
8gW9oJcePMNJP+nWKfbbMA==
`protect END_PROTECTED
