`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0KIIzfiPhKrWeeaiGffenAsRMxecZM3xVauEooQKkR7W6ANSfC6v9suyu6nUu1Ld
SAJAa9VhpladPyyw8t+pCvecZj+9sS0mzDYmnDSePrZceoMjcqnuJn3mCIXb+d0k
sW1GP/9O8WbFBBWki2F8rbtzQyY9olaZK9ngbKI9GWS0fnzEJ02DcSBjI60X6QMb
RN1OZvo6OqpGlaODB+TXH7jBZVbJZ4F4+9vbPDrbn+mJwM0KpWhR9d/RUW4yNEYB
/POQREQyrUdubxKR7iKfwS68uDfKXpkqz5PgXoD5DxPfMTpeWuKPGXb87rfmecdi
72nTP/xhSnbzMHpQQBHhBI95cyD59n+2h4AlGlzDbm22RNNvztSyJ/kZ+QP7JnXp
SZt+zyno7gQeRRVt+/SPqQzoT6Qy+HRli6fahb/bxaMR9a7CGCk7UVAGo/ABmX1U
`protect END_PROTECTED
