`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a+hpQlJ1LYt+Km3DP5ZTx+mkFog+SRdOkZaCCIqNqksoRnCjRGn4tHb9OFhnXVLi
wEv2txs+veU0M6Q+kmAJ/Ue7X1FDMHTpcxI46Yij5MsAQ/ajnIgd6AQPD/H5STDQ
Pp6pOgiwRRD7ZFTAAXrQ2YuQxfl3paNyTNqcsWEyBxbYMno796KJkzEsW2tAo6PF
mGjehYD4nQdNK8L6EdQB/zzXEgEPFK0r8KCDoT6To0RnwyG9PkxMAOiq8Nb62yf2
U1NaqZQu0UWwAfnyLZgXO1/UUjzmmxcCJFSJspyntqa4eJVmFZutURsgZ5d7at2n
tDvRbAbaIygH37sT2hBDsUmhA+8fiiouQQ6P3DP6EiW6HmSk+M3AL5yBsl5LKFVg
cl6SeaCj4KJ6k3vcZ9Fuw4DXERtzN7J0sL6cTPuKhEvQvga6wuoaK4ENvjZFsb5+
pmVnt13Vsnpun6U9cmGlJ68z14LkH+xlsx8idhNo8GFq0kJEcS7jN2JtHDCRY21+
aOuj/OmbH41Ilapg3AInUAW5DqNmDSqrQO4jrAgJxiDurYmlLX/FKlvJVgh4aZKj
Z0OxQJF3Gf734pjzMngeEy35CmYCuscm3+78uz8nLSU5Ryq/Jiw1A7pQfu8Vl06G
yvelgMkmGBF3mZH6FW0xQW4DbFWbmJFro4F8rXWi8VhubC52USMXB1meZn/ifIzA
cyuA8avSA4instm8XK/LknKiQrbUOgk3OvFz+v44H6UwvMz+VOM6HNkDF+K8vGqW
R43MDyAeFiXL9y9b6lrlAGAeCQEJbi5DnkERhL46aXgXmxrQTgEKI44fpB5yodPG
J0hft7fUWkz3YwxI1Ed2VHkXZwn4FBc5ONAqb3XljPu+W2r2izGtV4/DxF0nke18
Fb6UlZ5io/vDEc/cLsfM7mRBHFeEyeaq4OZLILN+cEhhFW3g4KpPXYaCJzrorcTS
/WTbYNBLNhn/JnY+bzNGYPe9BAw8t3zDUoFVDbQimLQk2j/wdngowFh2oItarxo3
y/cF63OogfKrI5pLd9uKdRb6yuOYrcAb8hlI2FOLpICCzB/J4nhJlY7GF9mhqv0c
fbDtltE0ptVN8Pc3kgRZjPmLbd2ZDT3SDr953beoM0GaN3B8YY1hAR5l28zc++FV
sD0Rp+T3gOBVKeXKIZjMD9mmiE/eSl5jffT3DsIV/uNlk0Gmh+M3QSmd/9HhBmQ6
tZ1LR8UKJSjHKAODm0h+vA2G76ZiEmPYOYtu6LS39vZoa/JJoqa/YPGZs37o4Uri
cXsKSOa6gCj3Icj4ERDacC6MLMymFZ2xA4R9cAWo881TqnpBrrL3ONBObwgq4E5h
Kn73cZojEZILwz99xWQT1SqHib3w/SusDCz0MiaoNZq7H5DSUZDwl0v+5Qg/mxpa
S1Ykl5wFQV6X2Zc4vXrL8vn7i+9UuYEN1hshd5BdqAnHQ5XadfxADX2jT7SwtELZ
i1tJCIJ+ke4EB8N1/G15l51qA/jiyCOgaJIaP1nRpQSniIUBsZhnqSLYdwTlVBBz
XXznw4bgr7blQdMbavODcoKtzDqI97B5+M0lfPy0rPVEUhTMJnXuqfvRZ06VP6FX
PLfqlhHxRYCjMEW7z7oLbA+PYMj0jNOj+QtVwm307mkMFG6MJ828DMb9ZriZpnGl
Em6QeEIX6UjPU0f7LdbEOx5lXyz+mSUn26l/iAL/U5AA7r0Jcl58PYTSXFPZQ8lt
xK317KT4joEgpIXPGZdaNhlh3ukYDsPlkfHkmqQblM8OdgJikclaiu80p/qLOi4l
3bZQUEmeYVV4EJsgI/OsueLHNseMW+rBmatfFaMMVH5eVOa1FJjP7pUNiUHpQgVA
OcIicAA8GLDzt0FjK59yU0k2Tf8yTKJI3Kml9dK/hME=
`protect END_PROTECTED
