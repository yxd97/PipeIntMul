`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IQyaCjx049f0MZ7BRmlGYq7pvlVkG6VesxmCSSFVv7fPiVZAsH+d8Pdt28qBUij9
3zCWpCPqaAvftCTJuZQ7uAlXp+Z7BRIxXaYwha/Wdav7LjNPHPnaAkhCVvhzPHh9
IxQb+CGHtkDSTo3jQBJA03pakDF29rxKqp2qBPvZ/URDBc8O1WRK9bj+fSZm/Z0c
VT8LUW0avRAqEXMZ7tmcgcTuCxrf02h0moiLp6fISp2U5BWolczBw+WdrrgJ8/Kk
Yx1+gFHY3QG+4b0Pl/k8syw9eS4mrh78mJEY8k5fbKUDgaFY/a/KozxX/BV5suFs
nxh8T0ueMKN+By2Mc42BH/JuYSCuWucc9gdtBbz8ucye4rJ/+zottZar1OUy4r7/
aqcQ71BVKKkXtkdN91meieSmsq/bazGJ9y+AnQPvbyUNtATExdwsGy+2Jxae4tmf
jkYuOGyjEl4F+PfaZtwTSh8RaKI/C8Gy1gHkoZNXZAtxqD8wTtFveqI9Job+/PGJ
irft4coI5QvXBIRuhHEpfUOrmT7FNL84JaWQa3OAmM6d0vehFUskcZ2R6h/Ojevy
amp/9N4+k5VZ84sRkiT7o3NGNwUSCUR/yM1SOeuFznlzSraXJphqZ8AL+NQ+nBZf
v845AbH7fBA8K4xSStfY4x3di4ZgHPrnkOLZ16caUEUgyNnt3o3F5tnmO+0ntiTu
TVNKEOAPqJ6rw1fmeWkbWLv0Vrukt3VQxiUnSx2eKKMYStRGPjD+DBYhEW7ioCRv
xBG8mT8KdU0GCj44HitOFmfSgjB8WUgzOeid1MNbuBXBZa9SaoI150j4EgyTvy7a
1cWrpAMD5TY7bLtutXssLizREhcewXygZBJqo8GKQQqhx63qWMWV806Tj8bCtGP/
X7TdnG3xs9gQYfZ5g9hOTVahbAVdePWWV65h+M+tUrYHIw2pmjsgVNtcgGJNGKqg
5IH/wdq9dyoZg/mOFEiQMjqC0J+SyQj+ZHBs67stuysA5AQjckoVEKr8bbYHz1X4
WJnIWKcpZnX4dP1Kuwt7GMJDW/NvnLQ0njFv6wKR5IGSA8xtfB7OuAvGi6pM7/do
`protect END_PROTECTED
