`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SN+y8O1W+C9j8cZ1zVPkFn20kkgirwtp7Xg57AIl3ri8MmH5W/LVHwMwRvddl7m4
/ZFHn9HJXJt1qV75v533jLe769gnJgCeSwdeFqSo7AQMrF7zPmlM/R9fDoBUkTS0
v9377Ffq1CsH+xLkyDViyLADz8955BB1rAEbKNJKGGzVNYtU6IG0u9rHPWDGngHr
zkaWzXTVxWx4sBhs2HiZSUQKsvzlQta0URitHr234zo2NQBBLUUb1mNJupVcK4iy
HwTVHEY8mZuMa1QeTKBl2ngGNJQf3CgR1VJ4VOn81L9AhKkVG9HyInyBIl/T1iPX
IpLm3500mNkphkD1leB4MkPd6bdM5r8N8LFIqzVNuEX+/7RAapNYuh4RlNOdP20+
7qiViPC4PxhlySZKvDVA/oSbhnvkGxDCR6A6XeN7TTOh+SKwqgivuhow2Tn0S0W4
X+jmzR5/hve6g2PzD4yn8EvaYp1og+8UaqEufyPkOSjFpOisNPs5M3oU0V4Ct8D2
GlhzPlbs9KwSlXHtEO7ybohUQ++SAV140QkGF4YtENxdQRU4vjag8WewVbzDobV/
kKmgK5u2jokILCB9hEKl06bB5gdXCyZdMgRRUWKXp7RQZnjAdtU4K+6KH6CwNBXc
8c4DnsliOf7PWn12hPDMG62U+uJqFNdJ5yXoWwgl0/BVgIE/sECb8sp4wjPUQtgm
ih/bL6WB9168Up94deP9WFPr02hNeeBOa3UjByy4Flkq9lRmtlvzr+DDQIgPj/Jc
54ZeEnum/MwjcWFA4JRY1X5PktuGcmIIQwF/WzVAv0YgvqIyhXSOF5HP3OrTYvks
XhVuP/FI4VBO1aQuCDGO8EIj/2J2xwX8c5e7Tu17v/YkSczEKArpmUUlI/cK20Do
MJyiUc0MrGZzqh2ZewFyr/0bUwSPpKFkJs7tiZ28o1Vh9ZdJhTgfHHDqGSIOOdzP
`protect END_PROTECTED
