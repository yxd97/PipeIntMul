`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
flMoqLkn6RZMrHt27midZKj1iz34+HGgOIUC/ED5Rgz+WEz+vY8Y4lGNwTRg/SWG
7qPe4kKL5aAT3qwV7vIM9nfCRfZkzIzHaG+8EuKQh587X5fWUawrdGVjb4AvCgmB
yy1jWOpyL/K2zgS2aAMoxeAWxbwtuplEcZ/UhE7IzbIkYIiXsZ9w80ggdd37C26O
vEkXBIDxXln+7c346GkRGovWdggs2A2MdUfqWekEAn2pOwS1pUFngDBffVvJFkGq
FdRz/a1lQGKh9K0J+hu05ufZrFsOSkmbS6HkF7ReVORmZfWI1z48noJ+M3UncI9c
BW+TDcL7wvTvcvS0a3145WlIFImgSRzjMMQ5nbNyPHqnJ0T6FpIUZS4fxk63mPvK
MOqfTPGPoQcBK3PNx+XulNfbN0FL85DHzpp4d8G2Y52cNpDY/ZHLgLHTNy9GMoTU
`protect END_PROTECTED
