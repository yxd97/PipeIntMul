`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7UjZ6gGc3G+J7rDiXfht6D8rmaFyN7Z9uRjLTRsqqMXAlf8mhDeQipWXwGo5jbiu
q2vzkM8GTyYyyjMlncYQ3ty4hBUEXn53o+VoWR8SYh4FZ8viIbYZ6XQ0x2THAwgg
vMZW/BsX7+qNi1I9dFnCFji4YqglPZgp+OBWQfAvHWFZOnsaQQb5wgvv+SgcZgHO
dzJPx2lmU9bruceDTcekz6XNib9VC7d8jxQHG9lTWOxEROEthtJdgUl7WxAXrTYd
f1UolHEjbWrtIcPIZuYvTem2wH9/BnLa/iyoTu6y9CVjDGxj9O69pdasCOL1pn3S
/c+zNeH/CohUdZTDNAtJKEmowg8ZvX14oEWUUX1GglFVUkqdlH76/Z/ITsIpn5WL
YMI7V9SaRAo01cuY1CxkOoJkcdoE20fymdwbDRlEgxx53Xn5VePKeG7bsKv8fxj3
UaKF4nfbSVlI9EBIhIUHipE5awdBtkJTccwBdRiY+BceQ75QiGahQ+zhlGf0Lmmx
iCf6nuHH0RWLwEbsJVloSh+yVYgQhspTvPkBTiTjKgGA8bTIZT5axpJipE7P+M3E
Ty/uv+vzNV9TopQj08T4psB/3zbdug1lxYAAATfIWWKEm+XY2IVAqJ2ky04fRYoW
OsnVct9EOdG8XOzIfuMap2yG8totnEaM08of/QLmMcgdNwd7oDdDn1JOuOdtRBse
FoH9jHga2cjKrl/fMPfVIcHamgMXDAhqPbCnjiq5vnPc0ywEKJ/npb2gwHyCc+A2
KPzvWkLtcz4IfFRvk+b6TOzoVOTQL7Z5Uu10VE7QOJyhDHlCghB0yNJZG589PJAZ
zFxHhH8j+ve7PqLB+GHBNjje9nTG1HxnqLGxl+fRLxuUXbvdcS2WLSdHlU8SBXf0
vwUxQijC1lT/K+67vmtlLxliSlROwPKbaj1TI44SbmMyzCkzZNEElwNc6T3nels/
YamIjBQrBwmaxlR08jVvj2XxwZNYDLtk3pr/KhZiDxE=
`protect END_PROTECTED
