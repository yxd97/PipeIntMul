`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQ+9N91Cp6ujrwC1dLjm2WiGPzDvw5X7nEDPXa2oFd0Gfzm6A3Y+y90q0c28XSPz
YGotoigBUjkAtCWnyG1Wwryb6UvN7p/+EJZ/cKleBspfv5Mwbit7k5nM2/pspxPF
8oNkDirbZcklwqZwiE151D/tWzydtfEvFYzKdDYC5QVaH4rNbCthbgZV6KfwKv+Y
X+z5I5ypt+x76tbPm0OIt8QIGVTuGZkLN3WI7lJvkWkNvXihOmd383ynxqd2Xoq9
YWbDDlY3XKQTNrMBTD1HN4t0RMmCW0jB7nRJNdob43PjK8DmYPEq6xy/tjFvcrrm
Vu+aR8sQLEqhAbZ/HuZh+BBke3DrNDxzn39+363PwBZdB0pLQXM3qkVpWSGUHDut
amHJKpO5mAKIDGSQfdxlvj/2BEsqLeCEhtRlw/pto+AWrSqBODA56B2fhvRXCZ6W
6EeSV0qpzMPtQElwogxNUQEaHPD1Hn+lRGfdBaQLN1MOX1mwxPERQcvB64tgO77a
`protect END_PROTECTED
