`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Sv21HSB85KnVkpjNn9TkSBYQdUlQWRtiqp79dy9R0r0o4WIVoxhOg/zegMDqANM
ySndkTuBo7yZrsdotVhWcAbyAvA37sSrYIYokSKLGK6+VM8eYwY4T/SJpB/1gvz+
W3leweZ1xA1Qd/E3wfrFwqV9VWpcIW2Tmy3HiD+3CxkEAeSDmrCydz0yru3fxLkb
7doshyeBIxQWhb+ffA4PpxYNHVVeZPsP4vA5MXarjns3LqtQIIWmAbAnIIVL5Ub3
t2TXNmycW8U0ZRMe2RrND9FzIO1p0DH4SFQ3ZRAWNP+FzZuDGVh4tnOr0T+ZBxQt
wAE1udLByUH6K4xDCULeF+XNTXGLTuF+iLiLovg8J9oyl5Cjn4aqGLFgpnC1eRmy
0LNHP73lnUqlIp/W4kzwo92Xl3dgcMZdhsOgpmcIKy24wBXjlMh18zdnmuZY3GGf
AAgAbAQg5tLZZ9GxacYRua8LWgG+1+ASjrMoJdxUGVa7PtKno5fjFilGXUC0dpt/
`protect END_PROTECTED
