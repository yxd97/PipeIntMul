`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ks1Mvdo5/D3T2P11mJcqlE2zV550s3uIqWQc7llf1tXI9PaqSnOhZl3X+HX11/w/
rzpFXBNkG00AD9//qK+9drMKBqGhz8VihHZBx/44BlkiLSrfcxe0JYPWJsARm/9w
tsslhlkFJez4Uu6E1Dkta2UWfRRzDA2EFu+ZOCSlWUCtbeCMxu1anIOd//xYc3L8
Hxp2Jc8cT60BIRWRFxga61SDOjYl4CjLYKFkAitRikPiESe3Ilfjwf5hxNW3lgv3
pEzS4T6HDX/91YKe15gjxYUNj6AqAh1+CbEFV3mHUX5olqx3i2PM7MXGq4YhrtLQ
EF6mY+iXfF+yOMi5KcZ0Xn0JZD+Yh1kZQ+0sX2UvMZwv9pqkGW9+q4kQqifM4CHm
1pi907XVrhrpcNKy0qX/4rAOt+4fIJqKKNdQJDWEaDwRrTBO4KS9hzK1pI/egOG5
Vo2onXwYk3U7TAhdSGF8HsCoBagtFrpn0VGBGZY1wTpLGvIgX/q6txvQoD2leBig
Wzjcp7dUH6DNWVJ75DoTyUOtJVdc6XHHlivl65epggIiDXcUfy/p9Qa6zaT0kZvw
GnjU7+vw+AgvsuUXg9o1OmGNwRgRgbDP6i6MphLN51mboyN1/SHuOkeRBKS8Fm1n
TV7gcrfOLHvWeSzR28ySNA8IVa+3FLOMjngHjtX6OMYIoixl04/MBojvZpsZYmKA
5Qrp/fOzB1FUAIHw+OE60Szpg207tcXo01IexuZB9AaO7eKh33CbyGx8GrA7USeW
HQ35o6gN204uvwZUbvP2PEbC9pAwGcWi9TGBWSTVo8jLfotRDjagycbBYBuNK6ZB
5xsOxB+p9f9yKTr/rGI3ISh+qMR3PTkYIRQwE8NeH6X38rPAfGNSuNWWAPUu03zF
lvm0psOSdHrj/+aSkwHrifDZ+eMcNNeHfaTZ87Zd+H+har8jNKuxVfusnJ+IBoB+
b6jk1L1KYr+cMDftpcrURiZDlp3PNJwNqtCTf9rgmyxS+LEcOqRmT80tuD8ILE2f
SgZ3pkrfx0Zoe8hdFNOtrOjIyH+46tYAMW6QwLB+ezU4qReHy3nHpTmSL4Fn6ccb
`protect END_PROTECTED
