`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
88TU/Vj3ZGvlxisEeuwkeumoXKq14s2hLjX7ffS3xQSAKGLy4l4wbohEK3pSNHYB
lUpafUwMZutA9E4eIdODf/qHQ2OfL+eXKVzYfOidm02ttqox6nnvvnfLToaTj2uv
WcjJ0cPzt/i3dBdekxYjl4sLGxCPgqzC48g4JWUddgoQ711rDY7nFss/lBBF+G7W
nerT3N7CvHREtBwxDx4XW03U3vwAQRDwPe63c4sY8NX2u1SWKH+zM6V1P11glRaG
ZiZN+U1faKKSwSo8uC1WtaqjrNmolDvNj9nerKnksItnZ6vVCACEjXWkydnmXIVJ
/hc+J6m4xT88U4htCoF/8WEvp9RSGG+xnIFl4Tu94FleERpKthn+mqxV2bn5yXG/
+HnYndXwh8QchjjwUw27VfIs5+86DO3q3ZEIRHgczD0pE8fnfO7mtg6382/Z4dqF
WL5otpJG/tm8CoPioIgAW8SywQxAgM9lhBu9eenvYouGl4CXDIf93so9rNygtw7W
h5fwtM28rFjq1sFYi3ig73vDHNZPzsyxTlbpLYYt3ZpIWAw+/VkNVmwW/A1Dft/w
atX1H6l27fYpCWzFjKeSFLgzo1ZlZpIPlm3Mm/NfOC6S6gYaoIQRyOAW2cYiEGUs
9rmEUPdP660WSvUNxw8dI2oT1AKzeqM+RqBy1EVUN2zkO6o8GRNULubxaFC9+Zie
TykgbtoxxiwAUzyy/kG3h9H2wZcFisONlxlI6oW+NHxFAIpPAcjTSm5zU1PNFmws
C2ebhbhc+fuyM35tbzbUW4kP8q0eriYrRgqVkJ0KQ9hkTBcEiEHwEPh0a8Jm0nm1
08koOoikGs+1G4aPLqahFIdotnCEjijoyxqkABiRrjIZN3DdiAiI4/3IsjuW9LdH
sIe7bn6I4EGLVxLdskFdGvl6S4IVV6jU5/DF7TBnoCHGqbrRGiN5tQ8KaWDwSxHb
+yZYJx9M4MjKVv02dytfp7nbG8iAm3aR6NdcuAxDIbpA7f0r7Bs7g+WjLFgVnEjr
v4Fs3TnEO+v2zq/SxoqMz8CuSXkpFvv15AeGFya2Kc1Ip8GahAVjhUzm0fOjNuMl
Hxto4fJYXy3xOeCRMSo5n1/HAMH+ACr0yKSn2IvFyZa64iNpeiKIRwlKsAmKk1I/
WG7X/mG2CWXXW+oz3dlEKFtMNPLh+gzD4GVxm35qf0Nc/9IhPy7XXmMDfviPfomN
jRk9g8J0wHuXGrGzjvMleIH8lHNvpt7FluYzCjKkubnK9E0NZCBE7cpM+fgsR932
hrMBebqxcsB5zF+taTA4ovlXaba+uDRQXpYE5RLwyTxZxCLXE+rhIUpz2tLXTM+k
i8z/7SbjXgs+NzPzLBOjkyb/Jw6SS1pCY1+t02qQnibuMsZLNbODBV0Lic4gs8bs
KyBrGnbB9Tcd2X3qPdDE/nY6O6lBtLMkCeP07jQ9aPClw43uu/1EYAsh9Bevl2ha
2/XyOr7R/wpg9mt8kGScWGxloXKENZDgV/Xi5GumhruFKIbDh23MXV4PxWkn8FPT
MnH/dg+jDigL4kJ98VoDBOEWUgr7qHn6EA35KxpDcH0GRygGFTFGN3RjXhbjlMSy
Un84Ilvgy1aGG31DzPuSCJXWj5cRJsrMEoL7FWIqKdQxImyXc6CE8jMWFIjmHPw6
ir4MzS+BU8ETtTiyEB8wXVi7Z4nBKcIjl6P6ija/0VXK4HZd6yN3xi0Lird2XB4D
GpKRZDcvmCsW6ad/k0+HT68prHJhVJTxAveVH0bDWwHpd2RQzH8xXZ80pEBUDYqd
eCJStUAHTW5+vJw+QOibA/QlcUd/xY+9P5p//8GplSbG5H1uXvHOhIJBlHS/fjZ0
tPUUTtrfn1q9o/kAJ7t2S/O9S9zfxDlWwRYafvHEbuNj1DK+yNiAmMZxGaVPQHw+
iMKhhwDfJpwVcm+Fz51G92OZxoLLKGUN89xRmctfLHQNqVtabMnKt2mGFX9PrvzH
5rsRDgOVpwK/xUHMvWU9WW8prK8ag3a9Ug3xBv04d4itsyHJTBbv+C5Iq/OrYbgb
PRWX3X5pxV8UpnvI63U4hTKNJibUClGpxdQyHWDr0YFfDPzjvYZ3fZffj99yRaxb
4yyh1nZ9ygCB4BeR+/iWz+CBqp6IGiIVfbP6ghmcvTWIMcZtfUA7IrwLi4KTeQ8o
Ncbbn5ZudAd1/izcCFG0vAGJSJ8CgD1wPPM+n0rG5tLqUW5WiDm4owdrBMYWc343
mmdl1VdNKf/nK1/27h7m+7uws3kwD55fAEdA+9VSvwWvqQVjN74D4WqkjKwt3tNS
2xNAwpLELH7ER8Q8sKWP+iZLMGPGFLdRK/YGanbC9jytaAnzIVcmpUpzf1BGRUWZ
B6e6rJKBWpfiBwEeickiYV4uuCxCvUl7E8Z0alZeIDC/7oyeLdC2BgNUIzYhA4fJ
jZPIGM2nDUj+siW/Rd1UJrU8UFrCUtDep095bMlwa1gabo0Fc8/FybxgrVJ1PUz5
2nOIovfcB7lpWUAraViy+JG7YS/vw8t0VrK4GG2WcjehJKV9Ewspi/TQ59v+7WjF
DQCYkwANcqqQs/q0m2hjZVgJKJmeOiMzwC5DaNUFkBGrG8vXF0Wy6tdEKwmeaeAR
nSufaq+QR6Dg5HrUAl//npKGM1JA1U6EKRyB+AHrCJN4lzoXcVUjTNUlLXSwmO2Z
RwvQDsAZnR5AKhx0CipoGv6oku1eVJOnynOSi41xQdOIEkwjNDJP/1TP6DsB8zo1
9CH+VB4uvk5e7Vdn8BLYHe7KXllgYACJV/nq+2yFyULlrY0dN5oQm5iRM0MFnlMJ
r4LGnV1yMf5rRJj53of7HRmPsk3cWWoqDoh49x6SR5arMgoWMwdVIAwExomgdOyS
EsNrsTQ45h0DaqzgJMYR09xG68ys8eAeLVf/MpcSUvaZGdKaVBDOiRsJYhD+JlhB
J8VFOwoQD+E456cJj4mJB0fGha1RFEFdkDHEXZnMC7gq5hPKU2MWJ/aFoeZGp4N5
66VCgSlLAaedLEsLZfxuOq91HnQ/L1gNbs+rV6VHtC/PjjjkGHYNBbWdXYz8VRIX
6cCTgp8qc5rfawtwFWXcdvVC79WOTgCYzZDiPoVarDxY9L9/9JCCof7bdyVx8Gqz
HncVa42GghEm9/XUy8pulRudllSWu/xYAhrJZhmy261g5OwKC4+vp42zy+Ppw10L
IzJFi6WzF0S7LIEVTOrZJy/X4F7zdS+ZcDdyzpLh3NuwsGhbtfQnzrEC0HWFOJ8F
cLKUQI0tBmN81b31RM3cWfHT5LtM/z9tK0Pa/PQFuJUtYUheoukV4RV+F4DEqOao
4pdAuRyp7qaeMmoWjzGWeKft9yh/gXKkeu9ktNAikgRqzHMyLQWACxfwHT6oknmH
Pdekrjzyq6QvaojDu2krm//FasE+SylRWCV4wpClU4AW7zJLrcM+xFIKvjz8Ml26
5v/nsoESoGdBAyZRcMJonmR0/VNf0aUUTvJz23HC2+bwFxmieJma87Xi2brfVeiC
rZlo8NIAUE4ERbE/SfvgH+qJDowSe44hatUpYuNpebxa+DPUfBCKg/uh3THG13gd
FksfvlXkN5FaZxHae+qcUPFfYn5KCqs0S6aoRAD1Mo+J7juUr+Tfj5snZ94EalTb
vL8Eh/epwzdF0FLSFnYuELIP6mPfz7S27NWTo2yivDRrj3J9ha7MjNe0vSibLcaa
3OWARXUd4nTo8O34UO9eURYM0H6GnB1R3npc5EfwsvQT993cvyH4oYn4YFkIA4eo
xIRvjY6FK+pWvsqoGFLfOjbt5mt45v7QY7vBAAwQU8gFWd1JD6FTx+h6W2E78lyb
KzZtC9ycZS3xx46Ke8X1N9rZCTBM7Gp27Sd+mqK9Q0vL2XZmiwNZ1bc4e6gggolL
liNkSV96Pa91VIp1IOGKO8wbsCSwZYaCwPp/qAOrAkhxgqNA0giKt+qQ9z2S4E7s
PSFHvGHUuzcDOSNg50M265OHA0ZE7AAXQf+FysOP/MhvuOw1HUUA7mQWjLrPcdct
v5tf4bRYfzS2n/Gy/LZs5He7uDEqcj1FeRPL3aXe2wBdtD8AuiBx1FOFxcqYpePo
Ibpi8CI9TfloK511VCvldKTBpPVcOtLmvF7spSxWYbvD2EmRTxsMqsPuppcOAWpa
r8RiiPSoJftWi79D+jiH8QxO3zHnlL5IOn9LkLAEGuPoiX4KXT1qvXN0s6rG69F+
jKRCSVmK+3bpGkxKJVoECAbygWJ3oWcKdUvd/pMxR7XNCHgjV35JwO2zIz31Nr7T
LW8UXzO1vF56DoYVAX970FgqTbT1rGXx8cw0V7IHVgjfWo29V3y+wpHWA6zaihIr
uBJyGR+jnZDFCbNLgv0wiaVlkuIcuQVrINf2NyW7PdgW1V1tAs6X/H7uxok8xG5M
pOLw7MbVJxNSyEJgRAnPAqM3e3mc5wA6wTXzFBIbyAZeYg446QcaM/H8n1fgXsba
r+5mJKeuPy8eggw87nFG+vzVN9nBag6AYD5kN66tjpN0DyeKNjaU922xxUMGOpRq
0ZCt3KwFR5FRPRtZojwoVllcOqX7h2aph84/nW7qdU94SX8/YbJ/uQxqmtFagPdT
6y/wRsSTfxKYIyKqC57M+tRe8czEbBG+Rc+wP1gtk78PpvfFNlgBHPIMO7PxiG3C
/ZQ67fopjV7Lx0zyTS7nXcmOjsd2j7VqDNCtYPMNF+BM0LA5amiElUoiuLfhIXxl
h5XTgHh6f4lylwGNqyKO0vTZK7ozfM3xgSo0m/DkOOZYQN4zLW62SS/xcn2sC+jc
TUuXL7balxIAkhNQ5sscJCiNX5kFeEB2Zp6+DlWfmyNVe1QdIJB5fV0eEWjoCCsF
LbuBN1Sn8zwsC+O5GtybO5lynjKU50sYqRG3+8BAH7hEkFE31xAI8RHYNDn0Ygt+
9B4MSMUdemY/QbYcXsV6pxmK6nj5XxlNqK/9pXVvBHNvdPBGMK0XyW487hC5EvWQ
BJRKvJzJI63EIOLLirLPENsgV1vqtTRVUv9ESD1IAFSkinI1PtnPfYOIdVXPpKvl
QL/0dcDiJmod1R8cZoXJl5WwTJu/Bu/3iV5pCQGQNaTo5iiRTrtiOKQ3k1igYwBA
/TIX+YH1Xs55hkxfqjUOhRbBJ5wczqEpVnehSXVS4Szq8u7s7xlZMwXLbk5tLNZ5
SWoyKdzE/WD3emdC/c1SJ+nQ0VpK679o+hL/r5ssRxWZwHSKfe0rkoooTnw/VW29
EYsPYfSJYUDzKsnpCVZXkYTzlcoXlxRbUy0YDmI8caJxWpegQqa3lBmbdgwh3YDe
9nG3WTzaBjRztu6DmUehEZck6ckOTmOL2Wsl9le5xn2PSJHMXKDqq5jcfC0dSPiF
eXQOX0rDZChBh+jz7iE1zTEiDxmyeVqgrBz/m06u/FQqijbr82MPKpFkjeIclXBR
Qi2Z1AdvzD5Gp688dS8wUbLlSCRsD7wpViwX4KywWaf/pHHXpsjh68DEo/vl0UpY
ZsaruNnEzfOCI2xMGK83x0ocaK6AJtfU0/sm+X9N8xc4dPDSvsRMuhFHAzkPdtL3
y9QuY0j68OZnmcwEJVO8zpvj+aG2BBUHTMvVpyYL5+uRyPd63GPFuTH6ldtJzXvY
509mNxX/DU74pwgKjIBeyrdvlUYiEE3Wun2yWiPTd+BzgBktZ+5sR+X3BB93r1ZD
5mSgrCMRK4HlHEajIdXJ7a0D9ZQ/alismp5A/yWLqXF5+LAsT4cEdcbIzSN+c0N+
wDXrfcQ4itw+eYYLM1gBgd6AMq9pvKUbgXx5ljHu3zVvg3FOsBxJ+Inq6Yyvl75L
sX6Aez6hz22NEAfLL+rzDZta/zghYmSdHmjd1TdRii56F4CbrRqmU74U5w727CQ+
JB17LuJCdnVc3DUJ5bjPnEoJwZqyrGorDIPtyCaiSxdwKfXSKpyBv6ivJcfY9Us+
yAFF6NIe2oDB4H4S8SA2taiZ1JOWDzrKfvNnEdbC+ppZeSQjlere8iuU43hVb07Y
ziOnyFUJyHg9wWVNJN9brPmF50/W7m0HHcc1qqIBMJ7UPX5BgvGBhRbu/oe1cZHd
`protect END_PROTECTED
