`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2btqHLAVDzPm8c/dnzXAmJchPIdD82Y6SBCwPm9UMMmC+O9swnDjYe5Jv7M1dO8j
ooj7aM9pbBsh0p5GG1HH5WlDW4HKmoJnMdQsGEqCR7FV7IAftoxdccMlyJnIttlm
Y+cI/QRLjzrcirQgAWwLPpvxetygWgUnVPHe6mn8vJzof/I+6j9u3ZA7OE1LF/Fe
5K3aYF4m+pLj5hFpBakCbr6m0GrpUBfv9B+X2d6FxANT61+gqfvJ0VRcvQtEsjvH
78E+fGu/rnpx3G7KL11LKb8LfB88OpyLB4Ayi/6QR9Shag26dgOok0nF9hKHs8ZG
/shg1DKa0Bie+XMSz4QRxaAgCvncnfcrIoORHROtvP5DL8rwXdvPWH/yOioJwZJH
JlIll9SK3KX2FUyEaJz23ndbONpfxGTzWuoSr1IzNQEn/aM4GD0O8NC3dEcnLVVo
bdHMU5OC3S3p2GghU7JGxLglUzlZQuRTF1MdebN1wG2QOl46aM8db6KngANpSGc4
k4DmIShsgK2ZuoCKj8YW1f5P+vS7vvXLCFfiPBRzHyVfyzMtyHadccffKYAlJ8HE
E5V/VMdqqLuAoBmIaqmAUqVXvjnY5nJydXw3L2LfI2d3HmMaVuqxbq06cHO00Msc
udBp9/adxAlkK0G0HXY18e1gRS3+tGHD6VZi4cAIJlnJyW+rKeho9PNJAb55R0Ur
5YbepWdJY0FqlFgg/QNazrw2E6nYEStRtH65iN84PZ4FrXHoIJpmo9hq/2+d2/NJ
M9LPHex6YsXmZFp8fIiDLaozbxHEjKrYcVxiaYXt11Msz/icFONlrRIcgOWFm0Rm
EuDxKuzsYm8PTQ8knINtHXUhP9WaQg3IJNw9LJKN1SnIsmA1vQbq5TDwXb66l7a0
zLABzlkW/jK9kWevoEe7uwda7gCvTA1nQe1kY5cI/lHMsUwm3VHdFxskYl3Z8XVY
5lIa4aQ3tsEF52Q7LDdiwp9AaIfOm3a/PzZ9364kA0ee+b2pzWXvgcKJ5WlLSTw0
1pwfckvIZ8mz7PNa66HbkYl+FFEEIju4v9FJJCQCtbc7/Ays6aO8NWW/KMITj/Fv
aJc8Ol65glTwwtyQrAIaTiFUlgzEmLoREd97g85RXboFmRnnyGg5KuoMNpS8ndq7
HplO0RaRY4P0LTVqjJdqWeVfZa7LAVKtm2sqWmBmbecwvsZAYY7dQNSYkY7l4TjF
`protect END_PROTECTED
