`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5F8Xcl30dvme0q8kFIDsAjBx1UVHtXcn823zXz75eHJ2ul9pZwRu1boDm59Z7rDG
owhp3CIuV57uGsBU5V1biSQAC7vlP27X2TmrUBDYbM49mfnxfEkp7rvQOYmITI6G
yoQLLbcvxXbcOXaNBsZUIlVKbPDNbjgz1ibbRBFwzMSENvJTf/OX+laKynqLldTF
M/lTB/IfJy2JPs+xk8VZSm6/tJ4EFkRVobzg9UYvJImi4Bxb/PWYxZ1kK8idbGQu
zmW0SmDv6G+oVa/tIBNs75XqzcBdIaD/88HjL9+8ioX3ysv+kInb+nG8i9gMTHw2
SEJqL84f3qfM2gz7rGq8+B9Rz2sVu5BiA5OeUregbSJmmpCigXM+YM7fFJawjT3J
+Kvh2Udj+KwMqNM5DDVOC8nSbmndpJDb84BpwBdLW/Oy35nu1KKklXqpRoCdTHwb
bBcnaUewTWImoYONW/7DNmepQzjBjNOmTNAoTCbZGVnuUc3fBr4tSlZFj5Rhe2y+
gGD1pmzW5RbjjBBLptX91wLzKh/YcE8BKRQMj+u/zX9k5XSdqOLJA22CwLoaLhL7
UbktHaIHEu+ST7KxoEkf5vV8VN0A42Mfhq/jMMtjZBagW2UwL6ORPOprxUJPMYgp
OgR+lqnZDLqLb4kXFp2ym1H38I9gQnqBReu8ySh3Tk/OdiTu6yOHTtDqEz+XyeUJ
g8UY7Nhtq8CP/PlDNQpIFzipIb8+3tPipwB5+SZWFOzxwqLJKt0Snf2MHH4ftVyO
2cSAL0rGNoEa3a7BL7yrgA==
`protect END_PROTECTED
