`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UApfuSsdYNIYsAdxA55bfj6h9ux1GD6WsII+s5GWAphm1t5EL2eH8kJgTH9XNV6A
Q1LhGV69ZMN7LGf6t7B8xX2ozE5jVsCE5wUiFNytwRj2ovCZnbv+AiETrjFxh2wg
S3frKjagZ+NgRUB5o+DTNMeuokaHLehjXN/yuu20hKmPoAVmN59JDP3E7bSmwvkf
5ti9AyeHqIi3nViWW0rzg2812VAlYL663Lfc/3XjRICYF8LU/JnUJNsjO8tW0sd+
hJZqQ8YQ44ap/++DScbSAGWJu/Wq+Tw9V74ELYXyGNAx/Oc1odTKtSz56QX5ou3Q
zfIYyMC5m6Yh3eaS7wDdJvsX1lh8/IaW7VDQj2A9giY/HybW20L5gPwkTiFtPbZe
tzkiIlPp9s25KMw5DEKR2d/K3wJvO+xIS21Bfa5jXmZKf19muUmEYtZHA3B+6AvA
lTJnat0m2JzMfH8AiJcZPpL7RwSloexhoI+7EtkC3AO9ZDKMWdy4GeJikEKof6Sr
s2zT2y4jqX1Mm9R6JhkobpSXBid7UxNTUMs8e7brgMSowWdvY2uzFDlqsaJsAtCd
`protect END_PROTECTED
