`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qO+FIOyAP71Fk8AsudVUq5Y5u0RWdr+xWbXXsUs8ninHi+IvO1YrbRmHnBWRCMtL
TlNBOT+RWLI1+885oZ3GtokPNxJTz89SpU06QEkHorwVOwhT24MVC2xZc+Qi+dku
YWWa5G+WlwD2X2ib19kEF0xY2S5ud2YOvqae2wrSxvw5OJXCbLpg3X8lOOmpKg0J
/3BTJv++6yjHqtDXXqGJHaIZxWPQVvelgJl3onnSAcdAtNop5xMhM6PRZC4aq4ZP
8h0zadiXLG3MHspdrPhJcZVrP5lJgtffuB4/zInywqCVtbZ7ssVver4cdX70DI/S
TJ58mGI8dyIF+Gt3BhTq7dBMrTlSXBevhoZbx/qB3oGBy8KLNIZLQ2YjtL5/O2Fr
++xezzJOdAZqpnhClxfNFR1q1lbAiqc7DaLJQzZg9MZ3saCvR9m8CysG8D/3Xe5k
RtpvPul2l0xrW8YdRTRIPpgOZauFBTH1ms1ww2S8IoH4VSI3AGpGBQXb5DJg94Uf
2UVq5XPZSTqoTbH0f9gJgL6oWVXqDVzjvHn7gE5+u6Xxh6VKYjdxgKZCh4HiC5nU
AnrheKAnuPYkfI9RSgbHMvpZnfQZ9HSG9DI98QN4nnija3h4lmwGNuXHNsIVFJHa
jbAtn9uBV7q8ZiHMPnI9jg==
`protect END_PROTECTED
