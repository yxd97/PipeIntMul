`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LAh3x65fuordxO6df+/WK+JFLvtoMa46gfYwghpIfon8fODZlVwrffTi1dRxQBxa
HYmOgY+9XaVpWpel4KWjb/ta/LYKHZe/ZAwCbdi0narbJ5KWcqVYaVB107vaGX0J
mzI6pUJ6iU+9DkrEOdRI+4i6IQwv97GtR3oS75U3K30nCOPxED7LtheeFL1OGnYz
ixc41ID4mHjUcYSM7wCdGZWsDhC+H/jUZUm7GYfyqeZIecKvjM1+jmpjtFdarn7f
j9Uv6DlQjuQJI+YChe6sGCFI30QunJVHQZru6fs5YEDKw6H456hNQCYYGWejY3z3
CYFgJ8gqqHekQnM/xjjqblO4T0RBhuBPeMrB/oDb0pH5iH59NlAtuDyaTA9bMoMK
g4GxdlWolSeOsIkSxW9oflKccP0cQyaFFjUAeQvZhiKh/x8RUKSulx38x8kJBnei
jhyK/W/RHts7VHQa1XAZu9kkjH8RLKg9eg6r2AiVgVcr6jilhDjab852qMxPVk1/
GOEK+lY/6ByMDWxC78MiyuZqZKx6o+B/mFtNy/dafcKbtbr5I6Bvwl775sNiupms
QsNLbqr/sWmdE2LCGsg5r0uWqsr9H32Hp9JT9iOJS1sMKoOMlAjQ2ArewmNbtQWd
D9h8Jmn95uJj+Tm36KuGCQ==
`protect END_PROTECTED
