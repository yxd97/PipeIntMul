`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GylkD8WIgF7Gas671SI3syE1m0mj04KagY7aea818zruiqZouonbukVkOWrNbo1p
q72mtvFvDMr0tA9a2kzhkUEv/0EsSB1LsEiDCOxSgT1ESz2gGiUpY125Fy45IjX/
sUiU3yfb6IQ90u6h9EfebT2APsxfjnz0Fw9VafHcSfgYsUX7VJHLI0JacWc4Ui3p
7OJ1xjr8fh1U5yiNABc9itSdN76COCvi58EC6TP4BIyhs8PUud2xztJ7xUun7AXi
UxpOvvgJPKY3vy9BPP5cmcOB0/BAqm7nQ4ERDy6CowfXjzr5THB0pBZxjQD4T0IB
tdrb2luqiDYERhaqRWC8nNtLjIFkwNMFzWo73fz+ZbU+nYFw2/aoYQlnevd7LosQ
kNFfVLAirzl72cLsfhCF3JZXC16jh3EIhgusr77NXLgqNrtK+idHUHTuXj8mE2pp
cvTEFmrWV/cDhW1x8m5jD7NlP1EQr9wfL3rV2O1nPTh3FfkbG9b6DHDAezBfNaO1
VDN8RoFmWa6IV6UCo8Enad6Fl1artGUslSYySDxfwZjrp4kOY/GOFnXHeJ2F0cIV
kZorudQpr+18OuBLFcC3sCWiSaIvWWSA0Sx/0sYkK35DoqPpf28AgmD71HtTrVHr
GskvzfzIird3lOMgjcqfFfz9WYjoOwkRYVIomys+6arII6KHRr69Og0k5a9Fawpg
b8AKXkXddIeK7odybKvdY3yjVjenMuwowMlsCmOGxNGWpeCT7GniMrkeRnIU5eJu
bjFEmB5AfjAlsIHQYAL2j7BLy1YSD8mb947tWcdhRy/1sO0uEKqZMGwSD2G5PuQs
wvduHUibP4z339+AtgUlehcl38DOVW1Eg7mFaHuwIyS2L1XLyHnTFUmrC3++h0Xh
`protect END_PROTECTED
