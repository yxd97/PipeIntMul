`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8LF3LsblUHL4+hFuYNpKIqq9QLEBPbEVVYN1a1WYyZrhCoWNwkqXtMS+tnS5VfYz
dgOA5m0Fa8Y4O9NxCLvCCnp9r05CxmJECkqnlOWr8WzbHz0003JO0LW2uJV3ZDrP
ml8HDtKk7kJLrnR5dl2wSprijwf2boCoF6wC6dn1T36/1LMGkq+8iSjhKLcwdCu+
XW2erJ1ZFC/ZHU1EBIzSDmmhicFJZrxNsshbIB0MWM7vED9Htk7EDqJuHhLg+QVn
5gzmc0sqt/m3+rsMfEUIOw==
`protect END_PROTECTED
