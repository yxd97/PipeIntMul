`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LwhwLAn6YFG/tHWu6isC2JQDcP0QOEfiFO+mqAv98gF0Ppo9H7Ag8St1/MIKU7ze
g5Tu9HAGADKRe6Z/MzIzx1l7Z7R/8V1doXmxR33VR/E43LzX7RX0DcHYINz04zoF
lqn2J/ejUUdRtLTj4c0d2Z0hdJ1hM+GXp15GKmtZEZerTt7rR0Eat2UkIRHE27oe
orfkebH8LGbv34oMpm4NmEsH3+5cSBcdygBrNz17FCViwX/CBC8sOaiecWEF6Ztc
HcEOGDCJjaoLvBLgHQKJPjhj/aUHkgAFcM/Ydik1B3/XcYSB1YfIxKu6wdmLT8D1
YDhEtb3FSQkesnNYTBPNolDED/dsFAwcVQvNyBHTr68VRC82hfhb6uCORrxJSe85
1u1RKkyB6HPMtgRK3DI6hNDXjHviv6ynC5ouXRn4gZ9kmmBZxXqctAmF1FqdkLOA
`protect END_PROTECTED
