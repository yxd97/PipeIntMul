`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8JQLyE5yQR1vP3tu+4B2ma4WUSKRg/efvrnaQfkqs4GMBNFKbw5XXvg5ZusyTYoK
3i/0UIqJR7IS5cy6zQK/iMN694nsX4PlUAseK1OVEJrIDBgmnF8scb8LR4YRt/6h
bm5VK0pZ5zHSsx7DKyEphzajf6pVlw7h2DYsw1P6U7cG3PvrXwsj8Mm84unQQEu5
o9VdQe8wxhvIbU7bAmkDeMolWCfb5/b5bwjxRKciK3zrZg4LMuaMOfGjvcAJ+Wu0
DUCLg7fTX41uNxCaNy05KzqcoD145qwl854R4ViL4k1L91IuWyeMce4mDObBNMiV
9ssSiOPWHjLqRxI6uXLglGHyqPaoGQcL0CFXXjAIlZZKMdP/QOytKdFipauGsDb9
7CFCz/pRMyp/R1KsdhAp8i6EJZUoauiZG6CE6vO5oTNDNd1fA+DnXNRa+8OFWOU3
`protect END_PROTECTED
