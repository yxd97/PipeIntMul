`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7gWJo5f3s32QTGAudAWF/+BMk5IDTdi4A+XAtkeA0xHmgOV53kFSrGLjKRoYJ8HH
vpGqjT2oT2JO4N/Kg0ReDYSTjOMyTcs8afOR3c2EYndttBkoadvKiTSRI2ocSJoX
Qzqg3kyN7bSR2OFqF/f8afBlg1AtEgm/31gGw5CgIE4m2iAbpzmagP/raWCG/B7E
o8hkHiHKKXQXcLxUop2nPw5AHu6D5kilDdvAgOSY6DUnN6zds/znOBa2Cn7mew7k
9ukykYzQbQgbFjIAzVZ5qNYYNPrUZLbB5nuKXFitygyOoAlHP0dhLGXqGIiKVzoK
pIUQN750YzLuc4cx8aZXBPtMjYciXhkaRGTJ8o1Sgps8hoBl+yRlzfxSzgKXE0G6
cjhsh4XFZzPDBCoJG2KrCnkJZGSOcPQoWVlot7VVXdX/xgMGpKUHbGR86fMmnNGs
hWZK3Wc35bD9U1tiPFTbrDh6YL6D4aTyCK1oAcM9xTlEUt3bV/ObX5tRa9lSmZoS
ho08whHv0z2phIzjl9abixIxUbMdD3GAQkY02RMOQuRTuVHthz60j5eQK+tSywPf
HQDLrwdypl9GsX7Iq7SkLzyzM9iDCXAbUIA/bGt7cvn8nl0AlKejN7ErV8VnZ5QY
`protect END_PROTECTED
