`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m1+Psz7c4eZHwlZu1DzPSQ30MuU6KAYi2w+XQqNwz3SLkaPrvl3gt1EVZqbyCtPz
3dkgPVuEsO8+2oaCq0SmNoDQl9bs0Z225/IMNh8kSirFKg0bc55POcKFR1vQihS+
SmiB+26K0nf2TB42NqN+W7IsoEDrKIclLqA0F6MZ9ZsAg1UDhA3eB/pdxEAjBR5B
fBjkUkPeNnkc8+02SUA5kC+PKBR2ji4m8x4IG5iYxdsWrViIYprML7Pphlp5rBfF
/WMEA+zl2amoXMBHoV7mdLhZ3Yk8sFO/geLvAEIQvKSlStrUGxAwNOm+4+vcpHQx
gFXvhZ/xKFkBDMhe02y3sJrSgQ/Z0I/Fg+rYqvRKKsROlqpeOaGY2EY/KhVtZzTE
5Qp7V6GRf5VDKIWGpaIBh5gRuMzrk0sMFs/82fY5Ge7m0ArhugMgDFyP//XUCBh2
0Kfo/Uzye5xWW20DBYJX4Vz/u31azEXVylTeV8/14tk=
`protect END_PROTECTED
