`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TOcgC49JowAfjCwjGraCjmZSEI5RGwL7TCDPBy3DqFssNllI1YJUCgzny5NM1ZlI
oFZ91sxFQPVpw75E4MY1pJ+6LJCOlTIysXdgey+yZOooztceeQa8CvAwN70Wu0K3
DKpONMEAf88LbiM1MMbQY30E6TdEF58JzqIJq4vAGTu7pb/x3jeyTO/RxsfDK93f
sj1Zg/SqFcoRvCcW/YSiswCf3L7NcaNNXtlLL7qaPOVf6I743n1nT/yzvEtpSk29
zKu8nA24TXoJTnHDFK+HD+bafU/CTF4GxtyGZOYzQETWO8NGvQsPdrBe5ywK1Jv7
u/GCiY4x4JzAp0gHbLgF3Yy9Am3W50Bt463BHuLyK7w52t+wNozatK5+7bw9yCKR
CPGkYnA+hW4eYJLY9cyyss9A2aNoIxiRbwauTuVuMGOZK7HWJ8FKPgwBMhqGoFGG
7/GzhJAswnOrnZZ8BwWuWROLZQfsHabFr1x5PIGMM9n1VJSBIlnPeGIoCX7lBOfV
2CCNzKNSYt9Rqv7kNmNAtyy0Zt/V1NK98AhLaTAvfK6yKo29ZZu825m1aJnK/xux
wEaRE6aZyPCRr6vwWGmrKlLyCS6w2x8vd3ejFaTutXGUbk13EMgKX7JP1jJ94ULQ
NIYAbTu4M0b613WU+bc2cVzHeQxyiCLL0j1xqFV/Ltg=
`protect END_PROTECTED
