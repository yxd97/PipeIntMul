`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XD/96Q5nXgq/h0vc+kNEdPgD5ehMpWdPvcvPjPZwSXN2XomQHeT0YSg3d0cksfvp
b8qcvMmeXe0p/zMaNnuMh+PF2s7RBMOJ+vIaF84wsj5nEAUvCG1YC2PBFwdtLkH0
gJgqT7FTwhEkWEyez2cNUU0rg/Pythl79+GyiWg1Sy0pZQguGaeKW3ujQdr6lc7g
LZoZ5Vt7YKzFt+THU/WSSnZ1ozcTdvFrft5EoUSywl1KkwwYJI/SJO14WdrHRKkp
EaKGfV/8scqZMbwY3H+XoLQugALdfXWpbSOryWhYx2x2naUNPScjH3q4+J/erlYh
8hVfLGmCHuvtuYzm5eWYJKkzgRSSYGMipbxVB3YNLCRucsFHaYeFPKgiTtqnwKd+
3YGdy5MYBaDdp8UqxN6/nEEog9d03DdNAo8hLJGFgmBSz81MT/Ts4rcSxICDhBue
qYrO1VmAv3O/9TTeeYsvDcYpqXbnWLnB1+QXPSBiciCi3CWuGM5YE0l0S5E8DaFO
pASNsBJLqg0sLjbYt4Pzx1MNKu0keeTVvZY6e52vBG+Iy53gMmPYzCDgbDQBuv4T
CKXdT6pFJOOcqDgo6fBhQSnemeB5MwfNv626JrvLg9fb9vXfe4piGvNaMfganQY7
vhzU4r4Sp7hRkI1pjd1VdlIQ3N7XT2/hafmFvSp4qrr372BBonE/4TxZ89g+cd58
r8hhOHCV1LyDugcQyx4m/FSRmGqnjyOVzYk/c1raSNvmECOGMge0crTTkICfVP3B
ZhyA6Jzm5zdDS6jTC76/4tp337SToi7FN1aSt1Jv5tulNGCxUZLhPOtbtdoPPqra
Bz+LCkp/EfaOrDsnLI5tLN9mDpmU9z9elLuyc8rnDrP+F2g/0sPaAHzCUfYaINru
BX6EtPandDGlWx2rVNnja6gWOSPkRGekbXNKZzm1R0HdDaTb+O2EMNo0zaPOjwIG
OJAHXfYP4ANmSr52p1VmohgECBY5wr3QCIzFJ6LieDei79/jPx2EvpIVFuI/P+qr
LkSBYNEQRawmQsneF1mk08znZaBbi4kp/YC4M4RmC3WcGIfZ94xTNn2k9Rdem1p1
wsigYKDohbVmo5Zwyo9/H0gHmo/eOKYZ/rUNV/wHoXdxmpQ7RA5NFfwTrDCJ9bnL
N0uTOQt+n7zdn1eZeiG46F2VeQXIY2F8l/0+k0hfUsCsKY48SOT1ibUaLJjfYB/8
OcUrTAgIMO5h5qtLIMoksDDnGPbrILHUp6VrlAZSw7h/9giF6XCJIZCgoq+SRKSu
sxivXniVeHzblk9QZH/NTMbnv/tt1TTPso15FT7jB/xXaBneidOYFDbH9sdbErRe
TdzGk8c7o6ev+MwqC2NNDG6iwsuKAMT/Nv99p0VkZIvX7d6XWf3cssHe1M3cZW50
8U107v7AfWwpdZIYoZ9qaUidyiFvYb7apc6soqf+xhnDm4H2DquSGsux6fNMhGOT
/axiFhiI5M1JTtmFhSJ1FkapfSYwoRzrWo+9rol41dE4cnENIU+TJEvYmluSAKPl
nCn4hVpQ7MbMwRRDggDbmgwEb8n47bOzh2q00vFIax6vVLWf+HtYbNBsh1NYSSeA
UsSZ9tp0gRd1Lvf6MiQFPTVGOWXVfsAnsNRxj1/MWbjmN8NI6Fd4aM+OLwJisqsS
oJDU44go6SSgxn8r4QOrbD3OPVMTDRBeUvxl+DyddhD9UZ80zwLWLnLNZo8bDZgB
mDA1pWpjAmXEAUpGA7MolzLW7+8n8hr5XspT+i3iXMxNOL82ys40GCOM+fgH5UYw
iLXTsesbETp5Gmyh/kwBArYiF0NxGMJaJzaWdIglndAhqRBKjeJX+t9dxbuQ4FF6
RVHh2p+zhP6keO+6OkPatpeKRn/hkpXPgaPLGn22POdqatnDnwq9oV1as/pX0skg
s9VrjHweXFibFeSPB/MlRGKqs7FKqNRW1cPP61Fgm9A0B/Ef7MqI2HxIa+9eVCKJ
UFs713B/gstdinTLX41AZ8VJaGkI2pElTvM5eOrwKDwwIfyuCcCAv6/jkk+DhUca
5ReT067FF7KtbkXBY0MO4q+t3pXXGqGBVM5DFO0S/5vxZkzzfY3Ok2GmUHvl9ISp
KRp5BYnYl2ALgw+6mpnH3SRdRVNgtdT10IhJQsI6ZVaiOiqagLzHesTzUF79fAde
WOy/N6MXgyUzEjxC7oR5ymnJE6YE0vcq9ovDU7oLUyAOBWUo5IHziyBNhvr1CIpc
YQITJ6EzaZTKtIVAgBZngFmXewyff84Xryd6U3+VLEZ6jP1IDPKNwJX7/fS2QNCi
e7PN2rw57JXZvsyqimMsIRMd3xF1L50zgclTxUuEs0Wu7ORBiI1qPMzfxlof9GL1
wjtOWkR/4Z+JqosX/ElGP1j1pqYiUxNT90t6cMQM+oRDYcaSJiRzDHj18DO6+AAI
ih9+K8s9uXmjLsInL1nBLkLEzKl00G6lKbvzBCZUfVRMpL9fT61w8NuSV3dQIqYb
uJcfr1kdpnVcqskcDYHniVAjPw89upIz7oxyID/iHsyG2HSCPYecIVRKiUAchhXC
ulqVCfHxiFobvgSb1T6pvWepLdzbBGbHWzEWT7lOrZ90klZkFxfNolXx/GFmmyJK
XX8p4wq/JVbYJEBbs/e+f2xnm/KNThZA2Tk9zo42jE6dYoXK2NPG7LJc3TfbI3is
ZfPe2BpPeWqaW9V/PFeDWZ5uijTKIuHn/jZzu2tn0RrZLVUxRfl5aYv+I2ZB/G7p
dgEvUzMljVH5bdmOQKGUzvPMYcNxEDLDFGTpmGHu/OpSDIb8eo5yiPpyeCvccpso
sN+NJLTx0Rk6RQ5DDGJ/YTAUzj1qyrbvM+dpoUci6or+OvA+DNzp3C6RaVmkfN6h
e172UJga7Ms9YCVuQI5ZQRO2NkzyRJ4dxyp8uTnGexLlq/ANV4FS+XIL6VzizbjE
lS5Aes+K6r9L67tJvBPcm2t6mlOis7RjhhzHaI2hX8ha9ONrLC17nJWRfMuuj47F
1QcZeHARgLXHWFBWnKxmlKIZ5j/lWTPmVXkRVOYRgmQuSpevuYSm2vQppKnKdlJw
5KeikL55AFmzLuTtVj6EeZQk5LeR3j31GeIm/pB27N+yEawFVltOMnjlB6FuAFsj
tmqLPu3s0QY1gufuRe8duFkz+AbowYa3E8enFSB27/2qlBANfHO3NwkYHKwjmYRN
BDVcEvPE47tkbVSqWYY/ueGX+Z4tDN+lxoHBDSAT1rV38WHCmf0NBTivhtZtdUC4
gnoLetwTsfVR9u7BLfTdegV4b6Asto3jwuJV3mgAxurMIgp1VI1mmkOpP0YTE/BN
ldYyvNNI+DofSp1ltGlW38uKENuqqG63zFjvoqRk3BCBq+QsDZd0Ii+xEwH3JFs2
0HNOgIADyIX57YajLRvGoqrXnlrPD8vWJ/cvr25rAa2684e3HpqlYZmk50yKrv9w
rgZTh7nyMY2rZAwfPsL82wZpwXM3B+RO9z7Z/Czf8ivJqDhqk327FkJd4HjkrH7q
i4eLRORHv5tNZ8ZZqjCnsk+vofNEwVn3OAXtglx8CGSgHD4KF0ljjmEYiC4qlzSa
FF9mmlxaA+eOAyRW7EsZc6A4qZHXNFJXLn1XjaGCVpFxslpI5f1xaEmIwF1caejH
BtxfOl0rlM/JGSleRE6RrNRsza8gTrhfBGfmdGvgrpgdeFusn1sZINOCgFiPGlTk
c6qCEdCO389DXc8yxn4SEwZmaId6EAYZrtmXeUrzzzzcsIwmiTIFaW+wql3DS6Ur
LDPJPlbiT45X5MMvANS0nGCwDEXOfXRr3dYclvWSNVnrz0eN4okkpnzT8venmJ8q
UAuvJmWeokq0JcQ9nESujaIner22sHXzDbCcg6D44j0GUuIleUXtMdFqneDzjG5P
XqksipsWPBLhH/WY/wjZH33TuBlhYRWZ58sprCDhLxUjzlSi59snTajtpCTC1WzV
jaQO8PlPH0WLxzEyPwFMHgo3Hzyqs+/RCJ/ToSTg77S9s7rvKObEbESQ7eL9z2Tl
Jm3cPMIafTnVUAtNgKZHoQm4RiNedKrKL0OVUCb4PdbYgevHSttRWAgcXEwdUols
jT2ld6o27ma820zggCU0vboCHYrH4Rj14yBne237mlVaQi6IKqAPn+PhzqZXe59g
DgQP923P2Z/LNAGqlw1dX4WGNXq27iaOcqb+VNOo94tO5pF+hFMSuWJr0P92QsY2
B54kQZbFHS16oB502f2YiSRw0zLP8vnvgf4FKPFvL1Cy1w0qdnhehDVds6d0RohP
e7hArPBfmElDCeBC9rJsVMC9u8oFJJdbGbrXkG/qmBWVO20lAdkK2uKzdpVKk4Nx
UritxzubHc2wtVv0LDt+aQKREol0R+7ux8cZGU4v+pvYKlJNYikt5/BfWP/sJIkz
NU56AwlAx1dSSkGTZy3yb8lkBEbYRcyizWXnjnusKr9L6QaSwnSZrQiVzKFUxN3m
xmESaC8Ut4u7nFaZK/BUU5MYSscPXvTnAnJw7xBKNewYVn7EQGkTC9uieuw1uo91
ZgdyIEYKTqzsMeUyadgx8khxdPU494yuDpRbk79js4Xf48zkMYHVIP66G1brQkFy
9sJNDF0KBHPq2SOQpyoZBJVPaWSVMQ4moSW3LGMFkG0WlHUa4DneE/QtuhnVeV1x
qfHrJg3GlmLhwWXcHVfq/w==
`protect END_PROTECTED
