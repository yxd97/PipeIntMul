`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qc7M/rOtJoMbocoTwsQeUK7fYBiIa2XGISlPvFngWAeD6GsCgstk+dtMkz2RM++1
8bHvAc2norEtwSxFFOvCR/FpqW/04fOo9Jad9VAeslrJQQQ7H3m8TZG2ICAj/Ylw
Z+9hFYlfcbAcM7EtdsRX+do5l7YOrrd4bXngb1Gd6vkZdJQ9cCMugvtEF+TgtIlu
qR7hY/Coi+A84OlwzrDPlYNHucFR+oe4WorOfZxb58vHBeR14E3+aYYccjXeglwR
Ft/fGZZo1nO/Y//Go6bpXAqadWgdJOJB0BtRjiqSfpItZDgIeYTTGljaPXljcGFp
WpcscvvOI23tB8oNTMtEQc5rBSPCAjgeeG2By4waPgpQo1beFaZQ80hlL5cgev3T
kSNplvsPy9P0sw3j/IaOPLlVjRwCbgS5iXbXXkITeYEhlU2CQdMBLCatJ8SSTTBJ
0zakVmvBnzoIyPb7CYxjCMmV78gEShMxq0iF9ojmVlAXXPGRTY/7T1qBfAaBtkvP
eQXDLhBP+MZDm/s9u00FknTrVLnO8OUi2r0ROcu9Q7pjyMa7JdU4oq7YNcL5/zT/
XvxkdtDcBs9z/96NEg6dcHI47KZF1TMHm0Dq1vZ/KGoMIuxFpnkH8Oqw9fD6XsDy
hfRgGiohxYZO6ZkfL0HhH9KHMjIJWj5WBv+X+0H/s+M/kcYEzQdIXo125fa9kGX5
xQc5RSXGY9dS/rc6snRIXGLkkFlfw6+7fq0mafGYtX8MO0CfV4Dhe3Xa1ZUbplqa
OzQ3nySGd7AO0yTp6iLS7/9cvkQAN+VOsDE3zWLwCzI2kekVT+A0w+i5Y7yaG9zV
dDyA3XoIZRMIG/dmpR9ZLg==
`protect END_PROTECTED
