`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ICECwkFmm1Q6PQVszXxZsA/p2i6TcpUhY7bxz5yad/h7yD4e1FIVjNmxC0MetUp6
jeecTelf0L72fBUaDsPTdZLQCm0XyOye6JUvGg421Ivket/XJoAfJulxvULoBfCo
HRIC31ooZ8MYty+FWqINYQ3naru8i4zhOthsWCCZ+trr+rByQXS8K7E2LMQuSfxj
z7cUtnvkE01OcAOUNu9kV6u6R7oj36hyOjTT7cJPH5onWXPtqrfVBIVfnNUj7yeW
v5oNFen65Cnv9M0bVXbi/iErf48oJ+kL9wQIThHfGEJ/LeYfVc0cjNfzgEt1kTcL
UEtg5xeDj/OxlZgd9Dp9psZhlPJUqbmC8HJgTtX4Z2Kr29bRAxOMPFBOHbqIz6QN
tiQTlNBqkuagm7mJeiiFuGr9dR64oPuD1b/i37KwzP9Bk7yOfc78C1i6RDzGGqvX
bgFCLm6t7NAEb1qNnf66VAdH+MzJD+/d+MEt1Fl/gDE=
`protect END_PROTECTED
