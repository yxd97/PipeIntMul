`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
42nNJt9bV8hB35q2tzFMm3ayx+yyCgwlMUpeW3J2PR0iiVdPVxIJedFw4WifI81x
avM96teHRcFwi89YoKBfhuHmGRraLbd3Z5twaLA/8qX8T2JKiZuU6H39WpLYyTO1
Vn+GvGTX5UI5CFZeUgjmpz+x29c2Ioak8/Df1J0btTLs3btBCiO5g0OIT2p0QE4l
5xRlTHEkYv2StHmzZIpvPZDnBef1I1zZq7feQTwhMq7/R+AQ81ARy0FbZxFqu8vc
pvsTXye7xMlGGG/jqx8Qid4ufHGmgS7n/LwiRp53wSmg/msE/EAnriPJfhXVAtiH
WCnVq+5mTQuAkBnEC2cpll3hxfp9U0dsTYrXvhZ4E4PJRQZ8s41+8FIzBal7MWmM
dmJ1aFhXC2LhYlpmkx4HfYW2gOGvudVo/K0PWtSsNslPU6f0GhWiXZUnAsLV+imn
gJdEVqhDeGHfrcwuS+gp+2R1ebhUv73NPFf/yJMBf3lfLKEu4X7RNeOkfdxDyDX/
nszAgo44Ld3tmTqkFdi+cYYRLMVZ6MJIWe+eGT7EFwS9mJtHJ1FMQmDv+oULoA3B
5jDPRWPXEyIS/vWAjWfpc5J3D0h+SwtMeFTnzyWFl15CODnTT+SjQ8tiDvJjTgtc
bL1Q7DJrBiyuwKeSi4nk4MwSdpcuan1RN3hvpDz4EtDV4BPD6rO+7lR7wSyTvl68
aC8MD2WOJqOHLw7R25Jg/UGG25YV+0NNs9KsSU1vrQtsdZipaJsG9CiH5SFV+Wdl
FitKLZ/jITiNZjdb1yHVDDKVWb3qIVsq9mPMxiC+8+FNLHkUoULfCafLY26ncfr2
CUuRIXhNxwKBzgOaBS3gek58jjRQ3DHCCO/gVpVqy9xLpDWTZr/J3stljHzCFDUB
aBN1o7pIgYLFD48cKJ6gHTZYKznthLMt0AYrYVl7J3qtOo8T+25rKQWFYseI32e+
bAuAx22lO9yhKsVTi5uCNrEAJ9+AUd0QBgymexHtZWeObjqE0AMSLkNqr1BAwjCF
uannuSpXQT6BrfAlp5NKNa9q4Hjuqw3qi05U0S7KFNPFRklABpMXvpERUwvjgOcl
T9Dm03hKwOXRGJ8ThL8UHciod6LVKBBzKafkb3XAZ/4YCtOo289hwoXNz9KQZhR5
h+KS7jF6dNQWYMhvtCO8l9VtRdGc7ZLatqRVfRTUp2i83QdnoUreI7uMso8+HU/A
/R+yfWoHApP3jTYEfrYMMve8fKcXUco2TTd81Pdz14TuufRYZ1MlexTHkxeTWM47
mExcRgKnqOEGaYCLmD3ZAzq/FTKoCcfaW6bqi1xcO9z+9N4JEJDHHnFeW2JVNaQs
/6vPtZeZmD3iRvDcUITXrO7HCzoIDnnZAckkcHA3i1ot9Bxg2HJV4ON8XgPPweiQ
hx9IDHjXfB7o9GBrdA4/VWjbHd2Yi3NNSStaQz+06QdHZ3WotvQ0xU1TmBjuS1BF
DvAwe0OaPtVwBShW9kV8lVtrxbUADYWSj70TLm3NxoNddqaPaU2TftR+nFv3QHbR
FtxSxPt0xT2WfbqW4YRQIYYSVFp4N83XHNgjgdeLNoJUu/MldykHZbJ1BsnK0Nfj
k7zeLUfNJAX7xW7RsLZt86AVZNvB9PAH47nEfwyMMchY8sj0Q28IMuuwLO8d/rjt
`protect END_PROTECTED
