`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2+nuo7ZFWYFfwdoPhUpd0eYipjcdfTJevl3gjTazpbEUCXyZq2BtuwdZNXKuv+mZ
OaSDXZqNCJ6Cz1QFTnbLH6mKP9pnK86pxYGEZ4ZlcbXdvFQ5HDlMC07cKtS9xgSj
cw1DpHGCHR5LoNIAzzvx8BBjQpmpiXypPXONbkJW2ZRKwEgnub16qCw9yNK8q51W
6lygXBYeQhfwXXzAHw1P7MQQViQeCvYDDlZZcGkyXq40nF1ThYUDN3KjfRbvzcvQ
qWnd3X2rrhnvwt1iBkoqMA==
`protect END_PROTECTED
