`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bWJHeAnvK4n6eL3vOlkjmY0B4JytL5CAoKzf+V8eeollFnp7Dp8uXKHFqV6zmcnx
+jErJHX0wrUTxBt25tokgXcGMXdYfuGJbaUl/+vKZUV/Uw8std7B6mHDGgz+Lx13
UaK8Jh4eSJY/6iXQuQcIAkvDhZQnrJTmlKScu/2eEIHXX2eKqpkqjpE9JV4r4pjr
CygpWAlCrFlUWRDu176tGyl+XFywGp3+ldHmtADzv0LiThonEp0Gw+sBIcc3xMnS
vTExq3c/AxAR15myI2mSXGfiES34DKLxqDWySh4PkPUaYXL9BAWmW0BKBa81Q2hY
NpivyxXx/NjPqhCwr8fWCiapA3TxT+ZwiPvdhW1MkXQ2TSns0Cy1ae343sA2tlJ0
2ew2D7IKQtmzkpswJeOU9SxaZmBwEY/ZNV25zb/9ABd3OBOiCHE3bwu56i4xGcBb
uY3SjdKZAytB2ln4jkwrnjv4u+DD0QtFPedVtAWbphIsBBiHH17/M8XCfpEpTnob
3O18iMNmWUdgD8NF8j6gPPSzo0mibwVeAup7AYY01RW8+M7VwCQG4lHI93MNMxJl
V0UTWMv035x1Zhl/CVb6zQYhPuZh6ReHJu+BIso48Of0mVQV8FUX4SxLcHWru4Zl
n9WfU/XdrKi1BZ2e0rL1apfAGkItRVFwbYrsl7Qz3VY6P91djsRX56j/YwKUM0YK
y98maelHCcxI5ok7iH+tKbnyr7a/otZjn8CS69aobAn2Uzr0TnXfLhhUlk9XMqEc
`protect END_PROTECTED
