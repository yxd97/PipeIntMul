`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fKRCMBZfHG7+vsX/XmzhzBTcK9+3SI9day4JbWJp65pmgq8oZTlzYNXSNOrXVVzD
IL7vhTGB/nEtymUJ/vWRcAg/tvoza7weKQfJB7uLoZvOW4SiSEqPyuBVvIv80myb
WpUCudh3j2/sLoTSJROYJibnoxxFw8YlOnKLO0vXd73O2ZezOzec7HzVFfvlGp/E
s941a3A7AmChUt0JB69XdjjOseaKhjYjOQjvbUtXTAoE/BSZy53illMJ4M4WclV0
VfUQfMK3G4843W4ONcYArU/Mccdvtpxq6M5aEx5CoKhY5bGiaD7m9E8rbKAS18WT
8rQHi4LgdVulJ6OhlniNgeSGUi0bapTrCY+0apQze91PMEPeap+mxqlOsXLMz2WN
yJPFw+h2JSWvSDTOLPyrHKt02FnoOYam/YWc+gARk/QzBxC1RP/vCZHU1ZqEI21j
GqGnWZ6NNdMQQ4WFst5ROC0+BiCEE4ghS3D2qfAfW+o6GnuHaJwveyOvOTRYh3CN
+/mBQScrNRO2SLEa3EoMLbakxoqz0rr+v7FnbAXUzLU/hO+vYl4YTpaBQIQJmKN/
lcF89fPavsiBX0Ld3+f9cAZndNUoP/9/73IUCw2pFSFzA1fzAhyH3Hec7rSe2cJ2
0cz7kDQq+6HCz44yXkQqX4vB5gr8mzdxuG/E30pXjwTJsbIIb9pqPW3LDYvnMpDz
O4IIHR69sJUu9vtTZN4mCHqnYLX6GLagJ3AjvnW9Mk8PSd338YadBEUwphPcq/W0
MDD6VQvys67H6yXJFzVVm8xjeLT5TdvdiI1m2mTdqCo=
`protect END_PROTECTED
