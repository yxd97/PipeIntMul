`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gxx2Ua69XoK5DWN+zDtbL/28lQStxyp2lV6TNZ6MjLltiYXM21pF61B9awR576xR
GPg0LevD2TcPfulQEewwOs3Rg3zq7zJDHOvtrwYLCT/DsGqt7uzqUDTBDTbBwLWn
vu+g9Ozn7b1lk3J3ew9A7DR/mOX8t1VXglb9y0T9DxnXY6VAQk4jLjwhbwxyRVEc
Sb7T/nzUWWUxA+cKFcY+xyRJIQu2/U3lRDN12xz2nH7+LK50fsqJzBhb/1c/T5+X
149tIgH/QlKgFsZoPOiTRpwbROZgYFEYhPxLrSoudzhJTCSLDtorYgFSYBpF60KY
TTpMW9MzDNZUIQ/8HtGzXZbUPCc3S1EQRPLtQW4SuDS6OImNAzPlhtjcLQC7roSP
mHIlG6ZnqsJjk0lPPtyGczKA4GqTBpApN5+1qq1lYVUHx0Q31UTVC59PcpO+Dr7O
pbzOUHUMMVNo6++vpOB5dtxl3taWTfe1rbWEz6svtXB9SbJ932W8X1u/EtFgA0lL
o3FLWpf8WcYeVWCk2SypXMveY1XgGPraI1O7c/ZukaDT8S1NdzNDOSLTaorOfQwd
EQLNpBwVsxannExAutUTiqkwXXZgaTAsNs+Ery/1TkUQATuQYGuz9tJzdN4whi/L
3aLdP3Jr8ZHuHmRmWi0TyIIRUtz8mUlRqYqQo19BvfWTUVK2dT0i057r+yt1djyn
ktVlJbqjOeqOIyqLYOeXH6zSc2SKkIV6uTQX+2CFOQELbNiJANCgnvpkfu7XfgY8
7R03ryDd4tRTPjZfIS00rA==
`protect END_PROTECTED
