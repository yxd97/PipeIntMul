`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPbe2wuSN29LUUud66xeG8HAQujVpr+dejlmktpXhLvFSRUv8DqsHX7klIlP6X9P
yYHRd4gkZnC2OC6Iqauc4wuxZ7eI8Q7yZ3kBr6xQvlScIZub6jJ4ztPFaoRfxk1z
Dl7qwwXe2UjbMHoi2bwvAsIu+CJhbcORVEY0keXmANTUQwkv2h43B+vnYWltWo62
yG2XYE+lcnVaEQ/oCEvOLAliHa8jmexKvSFMG9OnPmXocEr6LQLPsLbOFH+SSgse
Z65a63rml54JhTs5UZ/daIOO47wKUL58sz//7/x28lwgCwF1YnOcF6pD03n8mqgu
VZkIDcCQcYA0gw0EwnHeteffVIP+6gUsrxhVoOXMxFwVnS9boVksXXs36PqCfaU8
/yxxA2wOVeJ8Ii72pWDwzs8ZJR4yoE97yDqxRxoNsgKxUtOUdKVU1cNccrUn7eTD
6bcWeslPoRjoXXptJ10E0DqQNPWxK0mV1nTiJDz0FJVZiepMQGsMs+859msFJ8iC
Z6EzxeHWhkLRziTS1W0upqKFjcV2MECzFumTLGDuY16XQ0VwCqso7RTM19egOIPj
uDs+JSg0/obLQqSG/eugLtxD0cwLbQzAzBlt4dUE99rjkf07l4rfoaUMQn6vSqsI
8yUipVT9JE38QczlO2hyH7JY8ApnjIdMAZfJvwYXh7Nu4CzEOWqtq9VAgGdueKhV
U1kW4frQ5RA1J0WEncv5gA==
`protect END_PROTECTED
