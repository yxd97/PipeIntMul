`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAPyNZhge/dakXurnZ1DdeEqrSESWEpWDJLHhyauXPATcg/7pMiLZtEWIyp8ZSQm
AXXdhsOubxQ3usOSRwy5Aez9yIf1M6tbWpOHBPLQdegG/yRZ3YvmnByAPBX2anvG
J8sVWKmkdfvA6oNiKPyFQC/TYsujR8p6rbz+r0M54sQncA2mMPr2c1IIFZ8ODoJI
JQTLZvkMDHuxL6qStLn2VenEeZmo6xi6WtZbmimlMWYBATFvk/xXyoiHcqGkbc4u
l6oSAFV9PYA1C0i/hTgRGwdaVz0YUrVC1o6PKRjZ9Dp2cV7766o9ue5qoPr1i1gb
3RtK/Wl4bAKbyQpLlxcKOx9fPv02xcMYDPl6MZ+UbpP66k+6me/K821g3wm2B111
KOrG02v6m/OKiypIJ4wFurC62OVRbX86/dCElne5z+riQ4WUsmlRZLesCEYglhEu
QNOctrOhmfOwN4njN+cFx9xvmt+GoJOdHleZeRhD1rpnKqKsyCCmXKVKUUM8jK2V
B5PLG+l4xnNaL4tWrBLXFh/QZMSojCmSsJvW0jOdq5YtkEhPY1TpvZW4jkLpc/e7
p7YTsj+WnpRN9g1NG7qaVCP3HZG/pCYcZ/4ObS0pkf6miQwIOfA23Oc8jlO2NQqQ
xOgMqx/DTaM7tlXG9ymQLsAwKEqqhyj0+t6E6L105FOW0pfHdtoGhr0mJKXlpPfl
p1Mr/+AKbZdQSYvMZW2HwKPR9Z8jpIP0Xw+zVcm5sCzaWv2YkI1xqNc7HXugmbdC
9UJJDB3FACllVIQwe2Ao7+Y8sk4C4MaYMxRFFgsuUQUDkV+4tHQKnRgs3xdtH3vw
mMWcM9ZvoN0+Sg7TxymzKANGVS5jhR4To4XYckvhJIA3AF2L9aW10I2LAE1b8QUZ
PMnekIyT/Snb9YTkG/F1ZXkg/TCzJnWc0UwCWx5ry6+wwX0k+4oBNWDBaqe63Zbr
pT2/Cj8leXlKCm98+ajwGcKTqJvDlTGMV8DKco4P+zzXSC8Q1RuNHQeZRL4mg07S
SkkDiUSPM3u0QH8GojGF70AZhOm1BkwwH265EECY6K007St3OdmGIDdcAXiKMk4Z
DUidCPNaC6yvUGMQwHOi3NGCGSODMpDlOPFpnWsiQEamTlv486PLsMQ8+Hy3a4iI
ecMKVV9xRLzCgaFVCCJxgZlH66JJyAc4xjlmoys0cD1ulF1SG7LtECqYmLSxXqHF
Ri/D5w3Sv/1V3J1EVanD7j98+pq1o3/46HrA87cUlSDYJ19J4gCuQBEFqMYZ50bC
p5gDh0A0EAfwCQ+Te12+VkTjmxwSFRHd1O5b3EvGMznh3vv5pCI05WhBEm3sMllS
/MJmvf7WzYSUdTOwjQMMlhFp2Fp7CR9tWCRsTk/U4jgyIl0oX/8lgjCxmw1Ha35L
yDQh3S7+uWIdvIuIIUPFOcoQdQyW0Ep1TWItetbUvI9h0yABB6SKmAwjo3KeUL2B
Atsehpajs9mGjKm0ANn6p4Rj6DWriThhe1m9wKKKg8lb13LLYD+fVJBGzF+6NfC5
YYRYtEyyKcN+kXBJwnnl8FFbfkC/A1BqjORGwvZY3IFzB6T1uU1nL5Swkkw/H/XJ
DIPJlrluF6DTXy5v/WfKTfMGLIg+E89JdAY7HEiHR0n/5C3mA6fTj+rGujhEnsAo
ZV1Hvr34sx/j9fkwagJubf3dmlejNBzVdsVsOIDiG3KY9DWCaQ5bYjldi8oWNlHo
otX9Bm3MbcwivCLESD+Js3HENgLjMY/4KfiXoxIosAzAzsTaDZFbpcQlCloABw70
a+YLwKe8wrwBCVkuQlDIMea9ZOBiK4e1iozzFDIYXYCZodFh9JbMRoPMBZEqqm2G
JBjuc2Ayh1hLzV4+bQi1xGxrd1ZXWYfsGbFEz8wkZPItCZg3O1AAnsAs/mEA5RQI
9xk6jkldHmfTyR1INx6EIIFUSr/sklRIKkr8s5aGCKsTZhs02PXqBD5c/xSoX9HJ
J2RlRT15kiRgsTEanJ6DCKBsNNVgQOhIpQte4wZ+tZMx5wVmyOOStHgxjhzHGbRf
oFrfFqMq6czsWNT/NIzzd8FpHg/VsCyBHu5UlqSQsiePlkrZ8Uzonusl27eNmQhf
fSALosc1P2ZLIbRArrrKWk+Thgrn/Wt50QaaRCCoGX/1CLktzGASfUnAgrqi85oH
DEnnhga/VBO3W3kdVQD1c9dQ6WCc6om3n0lHXm0ST6kvrkfRstg7aOH6wKc4EiuH
jjHh5WJA/DZWk0lyW6uTEmbGI93OWD3IdAQGym9+/NIimtnXxbVUvFBwzTBNY3Y0
DjCzp3wBL4iFwPhCv9dDPU8QB3tG28+qcNA7ZiWW8Asr9oY1Qj08zyYF2a0pDQhf
`protect END_PROTECTED
