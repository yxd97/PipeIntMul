`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N9PvM2naTHCEiZ+qTshB6tc0HpZJ0anxcUQ48dCMXU0JD48z7NCPiC4OcLC6eEyX
zqngKDSgoxF+Qm5PV7pxGkOT0kkMefNawp6TkEeMPJRo1wB0hIchV7VeFk2f4X93
AkWJk4r8fUMmzOaYrsv7ycb0owYwshz/G67OISMNvlnIc78w0Ayp7nJB3bgsmds+
rtp7rsFAx9ZasPq7GGRk30TnqHucnztyJ7odijIC/aUY0v96STEhfbMnD1n+yRcZ
We0gJexsirg8OXi/B0XTvP29S+/y6mpK7XvutXr/GN5LybYGklMin77Zmjis8WtX
Zfzt4tPNJByHvmK4/tAZ/OG6RmWsb/dcJ+IRH198ql9ycZAWBdA3q9gBPDsCf6QF
tgbJxSCRUC0z0HuJ8Q8sZ2PvyIw6CWXP1iTExKu2RGqIHQC0K9lssmDvoUBrNmGd
S+IRLZ30It0j+pU/onx6HghTD01wnH8JxsO3uflg852I5IF85hR0Gh8fmYY2xSm0
KOlYjhOprXvaM6sq//kEfB7S50HeR18vlyNTV1eaT8xMRo2bot0hUz9pTgAO3NeA
+oN6W8ywlXWpMV2VhsMuUwQ3SsQFL5irMad3+5dLrDWbOtLVrGPanTJTXuNZs4Fy
Q2vTxhzW7fQFkn4RrsQAes/aDu8H86BHrIHZKo1uKcQzA6OjSRJjEsTPqTb0W2tZ
YU7+XPrrno9l8aydlzf0GAtgdBS5ZnPqMvzhfal20UP1UqOqBKkvLfgIYkd3qIgj
77X8L5MLwc3301VVSutYKSWvuxc8S/qIICm3Tr8rJoYW2pPZZ8Yj7G4mzxVwAVJI
5klR1izzLP0fLTWY934LNqrS8MuPnEIOQZ/ZONCtUZhAhrQprrrm9Z17Ealqbsi6
IiEy2ljo7yBbKvrIFbZRyJYrBNGT8/wyYQGwJS0eam0=
`protect END_PROTECTED
