`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ILf9llDMndmoQNN2e3ibRyOchXIxOKXcGBcoAWQ35bKuCuz8y6a+QvpYuWq3Bv/j
tUisJoW8IbZeZiCEP8QYg8yIGRoxSec8azoK9/RYpXtoQEEVPYFuRvuhIXL7vO8T
F0SSyZZWKm6YbIMVvZmYBkp+yqJP06yB3aKtZOgg0njWPwB1Smys3vuF2PaUOZeQ
S5HySLvtzy/5nFn2SDWNRpKJnEUbfPemofugD3qB3TaCyrJQa1AYZwuvjrVRMCCO
V1EHia5sDHXzOzgQXfsM3gcVLXJpcb4ke2t0itCeyZocv3fOvfhwzLy2kTWoAO3F
nQHd2MUlLK3RDgLrfWexUhn6j7Tm9GUqJznUClIcNHeld3UpVyxsCR9HuZ2eXxJV
L0/ruvyA0oQpX4/ppWDqJqxcH5POoYZTJa8DGrFOAvc=
`protect END_PROTECTED
