`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+QYdoYT2tlc4CVeoyVZpHQnJDRK/1gtW0Z/S3Ueu6HI2Iy90ZVKtBcez1r1r+kT6
ZfY/U/GsXiiSJaxehdnzxzwcCGJc0ne2r4M4E9VpLx5QvPxT/L7otqDcACVQhlIS
O0vb6N8ZCP/vv3ew8WhCwGFgJRp8mGkXhu6mBzIXfMcQQ5SQ2EkVMEZww+UHqWa5
WHTyAn6CsXywBG1UITa+sA1XAlApc4u6puYzUPFSJpvpLOas5ZHyhHaOY3fNkkgM
g1hHZDI23zQBW0i2G5cCMd5sGXm0eyTCSoR2B/oHBVo3xw0/SATxrFZXe2/eb+0t
yLOGdvlZOEy3IPxImnSZaj4/xU8E51s9SlkQN4diP8segysfRmY5k8Iw+ZVPBjP1
L/PqMKlFTdsxMKseBwaoUhTKyUDKTsQzMMz3I2Gr5HjfZkD+oX6z2+EucdTC1jkV
XtB0iD5lFHwxVbCAM9ms6WxKoWsd5IxagxvzioxgoNRnV0MSUZdraRqUtstpc5eG
xCmyWewAA6yPuBSnYoYBcKZ6TW+rQeAyFPYoB3azyrFCp5PcM4LS9GMZdrnAVmoy
lmSiGTryzLXn2RoEHvy9LPL3beVc0ikKuvpwKF2oA52FOsld6iSa3nVeQxA6VcTh
MTGBltKoK+cdC4Zw+rzyOM7ZqprQRyBmRS4lvs+ceQFUkoYliOd5myVSCkKo+PVE
OBkExe/h/UAzcogsoTQWjqAQksWHEt/9LLIWjz4oqbRUiSQ+1xmkccvcciVWVEAs
1CJB/PXCy8UFZgGyVlZgzo/Y6HZGI1zpDgeiFaYUqaOjhvxLHJy7bUMMLVaMyiyW
5jivF2r8AsCpAtx0BotOetQIgMoFMyDWGvbH5FyyEjM6UjrH3hMYPAePuJOyqJAw
yAMs1t9B92V/RI1CV+DXJG50P1x9N7r8W65p1A+093Vcukai/Lb354IumcsjQaBu
U3trLthKJCJg7n/aC7sQNI+O9AgJtBKnBHxuys2H9GiJs+xRan3HJXEZqtjf+luP
8X6Sb0bydxFfJVroQrz49jA+812BL7Jqh2vZ+E80Wx4J1IqNjH3kZY+byFwZUkFW
IVbgzjEX4czJPAkpfY3aOiCODqRBrESTW6bIYq0ScXE43/gPFPb+OOJoKF2q31s9
R7cVsvf4owxcB4LUtGkNqvzLCPebMdzKCqqE2enNRoHZhZzumMMeS3L7EWxL09rn
ktdUDhfbh6666lIUJFOoxPxQ/1gWnhuEM7UsSIpHsbSx1fA1cx8wRDMqsnaQIdJ1
l+s2fw3exoGyhTJUdobaDfiJMMu88pO1+rKc4jDseHew4LDCKoc8E4DLQl/iZ2fs
WfjOR45gKQP1qEGMWlLolhYYUpMrBVTnFHvcFp4stonzWbHBo3VDNywzfOMdGrdj
b+qGvjkZ/h4cFUyJQ7NIj59jw5bUbBc5E0MsOmGHOf17WV6xuySxUZ32spBmhgE3
BV7dhwZS1dv8FenoN2/CjRLAVwFsMoUFzlzm8nUDm9xiHCXpjEswjt0b+SukMDuV
guyCVgFrlUeW0KlqCDs/O5z3ttWfVfodBwyMqlBcUg4oKktmScNR6NUQm/+fGGM6
Hd1KxENfE/DYoMkjdlZYpGPlQC5bghdwglbNH8UBtdvOQrmB+aACLKH1KeVD98X1
Wm0AxNXWe4U8kgBnFXgNXhDlRf1IAQPVYUPU8gQqVZR5jEv/ZjU9I5tcBdC6p9gp
RUAf3Xw8EpQl+Cbp60/RVf7i8b/kAIsS20tmX93D3dS0/RRUIbFuINxn5zhYdgHI
dU1nRWGPvhcwy7ZMO+LTEpY6W8sNxte7gQM9C9Xh4Vr+oPm5n5hN0nZ2dsobJ+6r
VIs3S+CewuxAttNM+bGIVQIB+04ma9/DIyXg+yH+cxdV8fDqsYRCYexna6N6PME7
Boo4zhFIDL6O4lKep1LZ78oecKmpiemgcEwhToMCof6s8pvAtjsF/sbX/KyrZlCT
U0wKhkcowQzcCQgLx05/aFqPzUTkCtbi16kFH9q+QcdEdrg5fR8ULkFHLmhjZyhA
ptReLTfnVb+jKOlQScw1y805JIdlCZxZjZbF91XdtdGlvYuwSta8mWfPLxO3pPoA
aoT3EP7mttQ+H/0RJnVATnakE6D4Yww7SJs/jtpooAOfk94hzxVLertXVXLex68m
H+v4TYohjlX+HicecRwvdYW5tchLHBT3egayFjarZ39PpDdXqKpBE9sOr0/fzAZ4
mutR34rw1TJTUMDHRUn2CyHeGq6Gilut7ayrbe3VJUwfrggsM/nWrm9tHdfi5KZy
jV4icnZSCyGehrnIiQrmubph3NGM3er1gg0E5CO2Cny7824wCH0lKRdHRcH7TjUf
PAjrXOu1SHIkJkI3WRtBESxeLU6Nc4ocZylv+KBzxJjc+fq972IxuW6leR9DzhyL
OoTjGm1n1Cmu3kQ5jLfZ7eUnKTpIYW8j9h9o9zEAO96kKrJaVD2IurteEpszrPBn
CSVsx/VNWUJWJvcocDEQHxn5sQHBJc6NGmyCL+5erVFOUaKtUCXPzz+0H/aWyAC/
HZx+PgZrzvKgILgdJvNML7uMik/mOBCBcNI29ulEp0APJUzb7dk7YBANzyh0M8ai
jxmDD44kiKvaeNQhYRGdf9MpGH4ibxrIb98wECk8yRLF9LPAsXT+vKjbmI2FlqDY
TyYglbyYAzzf4q80XL0fxG/u+xEQLIehnrXYAVARQBwzNshc7qIzQM5OaS6Bh6n6
02fMtSG9/wINN0GVQsSA9EZwgWsYUsrOGleznLsPBr5jd6NFZpbwfAzj3V7z/J1x
HtiGolpjJXFa3Eeqn/qwPYl3m6FJfyo3SSOq9+T17E6i1mFLjgL/Rqjg98Q/pave
RX2miPmR2EjKIAyuQuetidRWbNKv6go+IrWdbG+upmshwv0UWOuqzBvPTqo0NMws
UqpWmbsixz/uiNCUiSDU4jP6cJpjN9JOagNzoGaXhjFwnGsfKaeShd0x2Y81EhJL
NFFlvIAikgA/GPLmslQPmzyEhvl36bPKHDbK8UMF2D0BcVEG/8BSwGYsBDa6PcHf
c1sjiQEnlfSPFLIpXMUiMCCokkg3nC5ZMzoVMrMtBq4LGE5WFTsNCe660DR0FGsT
EyAA33ow5pCzVGcLYO1Z4WmtvqXRjV5ObaGv5oT1lAlwKdV3RNjD1Hg2ucEOjTSy
tCqArp2rAKm73Mw193JG+PTkq9TR4dFa7fEnVczHtsH0AgKYPMpQsspPWJYwsOee
kX119HTXszB0xg/8fR2cJrd5ZCPLlB5J8otwlxf6dUmIJRa3HTKtHbRT7IOYPrNw
NkJk9qjkJbwof+1j88/I1DC/o2/YwGLw17BYPie/SPVwLq1zKmVnrwn+JDy0G3gT
ZHUiT+CQr8RxPELZpCjKkatjHCwcSPZ8iooEd9TOLDP+uPTR1pg9r/lOmD2M/1gE
wDAH582+GH0pvaP4qfPw3A1kYG0bEN1/zWsCLN0momZVUVzy/AG9nACRgar5hhV/
UHYfvwGzbA46GZN5d/2pGZVJOgbw4ppsdKYnJXT1JV+aGVLK1Cb60vdItDkvsi2h
78eAG6kroq8/bOED9UfErwE+GNUvBKlWE1dSFi6WphCaWOnNlNbf9mlkwzJhe7Yq
JFJKCr8cFjGO/OM84xnBy51F8K3VcdjY50Uf3U8Ok3+sPEY29LKDvZ07ijAPtafX
HeAv14wLBBMsK2FZ/kDXum/Oo0Y9bEUlLx41kw6BwHanaAenfpNVGlQC8HU1hpSj
gYN7dw2hFw4/2dAl9U9QrvEkFxkvyAHR4iCodTMMMMcZuzT+A7q+n0S+TnpbvXcG
wQzxdIAbMNVWbhhV8y4AYPOub/ZWOQuiln7iXiV1G//eQkH783RQGzc+J/J83ZaY
28XInGqIooyidFA35INQ5RD9RpEVAPrsqCwI9jv3mjJ7r0qKMGdytNR0V1mSqt9U
p1jMJ0uhqxTZxoVEO89KllQOTDiEZHVqsxoSk8u1FmH0/Pv8XuOEOKx6zlaURecp
li7rPsENNO5b5d1amS498luk0nZ+dp4nwecpC9/oKlyt2Z7zHMJfcUiYWcJ+tm1X
6iHvvaa+ZLBQloqEKtWax65LKI7A/cRnuwXEi1ZShz3cYG5xPWrvntLrErl+CJ9H
b0GCsU7o1RIOTXbGp28aeSfJ5M5NffNYxmvBNS9hAuZTygy1LpRbtzcmR24bf9A/
W3WOYZPfSLiFGqtqTrS06FbpI36UNtR4BjSf9FtE4QGWwSZ7rXo7hFsZRzbWxe/v
n4ppc7fLsKXC/1Z4DoZB0MWCZhiOeExHgrg1LSfSFUE9DLiVPEZ9mnPu+w7teG2X
h1gGEnOyzofQWQ3BtUvxvYQbjzoFTlH1jXf97T+DM2R1AAIbK4kCJcx246WJtwVV
uYcKyxrg1TLqsz4NKvGgwFbtAxru9Jt/Kt3iEsjE2rdH3mSRVhGZeQFIIVOOI+2/
HmF6fWkTpTcilpw0K7jBlEkvzGasJMgWdbGKnhcrFJtPFmLiNKD6UEQwKo3q694C
RNRnBOLIQP060BrObC00/o/3GuyhrzWJezJtIcYw6uvJfL47S3Xn8IqmvwCdgzPQ
Vyu8MgX3CWLOcNEA3PQ448+0X4u8BCCoM3+iENkT9QmYjGiHel2l0tN9HNT840jx
OAM3ttLhvtNabDvCnQcbdtTSwKXrWtFV2Jz9heQ+gXWhiF9YUAWzcRZnJmmUnYfs
WJP/tIyogBNQ5ov4/zoHsjCv00Bi6OAypqB5krMPWqWb19LFIY8EuKQZFjaVTfQ1
HuCpn8zIK35/irrxpE+EAptxC2Xv7WBQmDw4M7iuRR6Z/odznF4kKCgfPN+Ngt+W
467w/drIEyNBU/EPWd2xy9QYypxb7ZNS74L+d1CWopENd2EhuvAZGfJsE2fc8W7O
757tgPl968ancbQxMMlVhhYfI4Nfm7XsPWeXOiaeB9EfD5lnEcPD4gXqmb1Ghap+
Ha24HKktQ/kEWx7qc9RsDt2h3Gw9Swd00aY2RbIA3bJWDPvz9GFu/5WtIV70s88E
FHOoVc+HbVKXiz+XXOCDfPY8FJMb+YDVmPlxDZl+9QucZtPy9wlnhSX5jUfdsNJw
8gpBoOgs56DPkdDs2m19ZRW1pwgtu8T71/NFigL7F5zcA7KKBfiZdqIdyGzzhJAa
zYK1credqPY+FlpCSz1bBqSbAjsk02wSHEC9N7CW18ubvFmoTzk6jIiwBPrOGIca
x5hR0wS2DtjyLd8jUQHrKejjboaP3DmxbQnR7YORDcmrUFgNh7fQfeWWKXYyREUp
xjsVVjTpyHH6C68TH3dofLiPi3SnVFktgjbZhSH06ORtkh4gPlbDtAr0Wlw57Vth
GE4SUV7xWs7HIf26H+2emeCPljgUdlFcZmMlgD7BICV/5HOQS9LN51X/84qmyN9U
2TbWZJaY1y5fNdFXDJYxv0r70pFppxS7EmMW2wDX+ROl5q5v9lbzkCZYXGvy3r62
My3UyRKDIS3re+4IqYsB4SmM55oJruma/ER86PQLsF4+ILsq/cuziJ02CZzIgbLU
suJZPiM0KApbzil8YJ9SnpXhvxMzYfpL3w/R/hRIdh5/qt8HoSSuIQl3112Mowpk
zlemqertewqOBITIKPKPqRzJXRcD1nQLfeuJ302pLN0FVBNOQV1DxeVKruoO1FQa
rePETF+2XW5xublvh7wnL2GOBhpCCxTZl7tUIxhDVjw03bNm0ZFvo7SPMeAm29IF
XtEP31gT8VcVW6pPxqGd1ZYp3o4YyHROKulkbZfd4eBo0AXcSMF4CVS4aDOjzt6K
V0IZ9UGehQ36iGjXlSydQvagkf4Hv901a5ynVZmI6v76LKSb+pHqv4p3a/wbGbg+
uUZga7t/tEOEg9pTEmk0NWXfKVCIrvFD48DvL3WsIMubBKH6dGMj01ZRwpmzadFj
yRrGV332Fk2H1OZhLrKEPL/pyWFkanjq4msljXnDZvpGyQDDCvQnsnD21aoOSnL3
tq4qownVqRLPUI2nBMK/oA4Cg2tx4PpFYSEDZZAvsX9/Bf9JMS5smdTCvcLwM8pU
8Vl2snFtGJYpQAmKXanOL+PWsYm3lzdPrQk31bXVQntXtW7g5lBLriVF+7JvP+jw
Wd0cf1gi1LPV6WzsokUiO53Fceh0cK43hWJXHXkNAa8pd49SXGeXcd25Miusiv7t
AfFtUdwSFQ2Gw2PD4cFUJh1b6Sfuswrqsc4FM7SaFRFHYqt0iEFZi+IkK1S+dqu+
KTbHw9y/Wb6JIvMCZUeRcbU65Q2FzF4XQH4cTGDjkFo=
`protect END_PROTECTED
