`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mevLSJQD8W5orQiD9FRg5mbBZeuJhjrF+99a0j/VBA5nkO7U6LTBS5guEtHIrTIb
O/3ICTyitODYqimIvapANLgeez/upTRTEepI7EZbWCOcPQkLrvuyehc/fZMGOCy1
X2fX8uc/1rVPKUyMVm+23e/Nrrsz34zxmhj8Fn/PflD4MGSPwyd6wE6in1uYC2S9
UA9Zr80yeJu+REKxjV9q2649/DrUg7FxjgpAu1Z1EmmW32LQTouE3+PHa/P1YF1f
N6TPZ0qyBjBOPa4P5vIws6mbzE4YMzIhHD4OLZ2lre9f28iIJN9HzlKIB++XScZa
zB4k/jOvuAuRBiPLwUlMLJY5wIkmABFr61KUMpJhd1h0adJvMfGC8WGOYJFG1AAX
HvGlsZbNH4SC1FIZASgIJlxgom8DvqWNx7b+K+CwacdEoMea2/1mp1wtPFPfn1nm
`protect END_PROTECTED
