`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tg0xkX3kyRAWzirROMDYzwjMZ6P3rSEIlSSMLzfwS1bV0j8nJ4iSVpP9rDI5xaKh
D0uveyCh0t6afT5kjkOVp6eCGomDVoS5HFqTR56WpBxQavxGBvqQM8ytYh6Y5wly
scRHMotlqUO6ywrVZgKC/fZHQ0RY+GctFF0AwpBIe3UFCBNskTQwjYcFe7AaLdm/
JQr1d1IaD8WW1K1W/xcz1Job5Q9MvtBz6+n6JCBsSP8irDhib+gJbQyfuZ+Eh/ZH
JjOxDT1ySPTyjAisVG4/HjSHkT51erGMr6aC49q8Y90ry1YgdbVCmtFhRruYuZbH
QcoiSkvBsyRLx8o3z/BEqnHwijwg2RypBgh1B/i0gEnI6MRz+ohl83RfLeG0Z9dw
OvApmGQUBMgWub6thaPXahlBnzHfq0G7YDrYWp3XiAW8XZtMoxuFyOd2YDSjTUHo
E7ib/5FV9x4b7IqQyG3rkyVoiDiwyQICK0PnrHsZ+1wG3fQGj7q8QG3mzCxEEsuo
somqOElxKlCR/0PNUb1V/DqSeyP3yOp9A1mUvBO/jnyMjM9hE/Lnembpgrgk/9N3
O+hrlppZVkMSIm77kRL+5mOdLalVz1x0A6IWold8EV1NSGFFdkMajuqljE+Ng9DS
uQHuGbunGk6dZf78bL+hfFnvZqQvWucRxyr3iW0Py4wEc/K/Ah/GUVCkcj6VNgEI
1gbwUm3CZ0RIHCtiZcHCk0bjptn60QaGpz7E+Nnb7pnE0K2uGZfXP/WUEThtVqTt
k+xD2Usq8W8HvZv4KyFOykoD2tsBahxGKr8aiiIdx81VyKXgb3/DQxkn6DyebhDr
XwSX++cw4wGtjlDima3+fc/952y+obJiq/LI2ME+JB7DEP3GVK1u2GWDFWnFUUr0
IXN9h6gKwC49RkBPMmrOGie2L7HiEcECf/ck+8kFdRvKesg5W0IpxJIesDIYs9mi
b2Wc/IG4kykgUzQuhqjodZcg8pcc74irU7mvbisyQyShoxumuuegTpjwkS2fWMae
mq0ek44Vci4kBf4c57yHbHnpw/POfO/6PkC4M0oVy7oWbFcPyXQvtT319+pyZeBU
9Dj6AbC3yAh+SovV4rx3y3/8N8xw8Pxe+LZ+pUfMQ1YQ+DpmM6kQz6OrAwqIl+dC
AIujlv5zGjz7MSooAVHbOgB5RTGGy51S3L0Sf9xB13BgbFlViTS2BsZG5qL5vn4T
JxOVdZ1l5oP2yJkBTSuQ7SGCX8LOost8FcFdfLXmTZtSBUc4p/cqO7pfZeNosR5Z
nDo7b2DZt9m4F6cJSLGtPABxPkg4oMdh6NzEPW/VMpAOZJ9U9ZYmVJRVAVHpx52+
sQmYh1DMexMTyWmJDeujwcFVD9YWLvZMc672xNGGLeHTWPUyG3w+7zgQTwMmKQIe
g6ufl+cU91JTTRATDVVl/Pnl9cLp9aXorP8BYeeBOVYuLhfujUxTaIVW0K0Pnun+
MWtU0RHj57zQSckdTTvE+EkRFswrnrHNwSmws8QYHR9D04F91KTCdiw/P4pBlYMh
QvgBjOXYtvGneLbiB8cjyBU9g3nkdW4bvat+dmAY4Tuc5TocG81JsP9zGO3FMiB2
9oKpQwTxfV3gZE7puU8rQCnGiId2/0VSK38KvB/RBYWw/X4NlOktPNNCNLt79+kP
lQwzD23/1JIrrh+DwLYKSzKP+HnjJuOUIE/nXavHx918IcmEZbGEGY7vHJpinnJY
r2nGPEv1UBm4FPFwz6UYYpGMrZq6N3NqFRqn0YMU5/5Aoj97Cix30llHym07+uP4
0p8RVrbkXxjtoFszKfojCAxB5PRwi+fBEVnFoSwvIL97SbEl92cqT8elT1IO4YlC
lq5L/Sz5LWEPBiTmNxoLjbLpgJ7p53iXfxSNi4HkbtC0g27O73gw71N1KDQD7rVe
B0mMXcosrvmil9baWm6U8CKO/RgxgJ65hYgUOJzHKiZgSYlrxXQDse5ztaPYEfcb
e3hpJOIfbxzV9P4N+QYcgQGsbucvPKMLi7rqKKzdUxv9shCKhQW76mKRkkcWQzJO
c8N6erU9oYtOeY1FOomVbKCO+eLYfe/t2KMTMR4Q7YnWD5iwhybCa4RyzpAEieQP
G9gdU8mr15X1u1SiSBplr42csFx6xM+UUKoDWyeDvb9OJDa8UG4zKCTsLISxywyK
JaitZazUHJ/tA70vCs6Kn38xcCs0xZDymFHoebceg+wVKWzoSntkY2pvwKTbGb4A
+Xra8alXVIbUbaUbRI2vJU6YTAiOnRjzLEweFyDj/OmAPca3EhDkX9991Q5mgpBB
ly2okj3k+JS5MHdrofSnrSxnYczDPsSz7RzOpyQysizwTZpkuxqvbiTsUkZPIEF2
KGCxQgJxFrMJsf8taJF/KcOfjXFBDPKQkPuwBCLSlodkahTRzNy6dTzJy6F3gkah
7xmJl5xczqxG4orrU7dzgBfPutQueaCwOsdN3bRaPn6B93LekwGh64x7FADU1k4n
jMGbLKIO2DzLQnRhdtHWeIlCD7taq+dbP2o1DcgGK06UYhgemWhj5tXOjv+c0lkR
AbqC0WwLVqXtNGkeazWsXvlW8QvPa5hXK5YrFU96fjiOnVzOM+UFjrc2YfzPs/N0
Y5Tiz+c2IINcjo6WBbgez5EchZqM1ZOrkeVR7x2ofnwBUmYE4r6PyyOX3nRRZoLN
UpBlv2hbu+/fjK6sKmdrlzoGqX8hbamLo2utjWKRdEQwUq7tvZ4/clXK+3t8OZYl
ctO6oExRgG6bbyNywZwyK+1glHP35ZXGnwc0tIZT4EH5drih2ew+5riM1tnn9BZb
kdqSo1CmBL8s6W32om7+ibFyv2lRCl1NU3lg1K4EfT6FjCOgXVdbbQhsT2rkSqjR
KHTXAyrctxMUkSafHfbEEHBsUAe4vwWy8d58umDIh1f0oR4MRS1YziK6s6AJQ23j
yOFrhqAg91kqYhBjruL8wzlkD+cCvWkCRHiFYCzxS1+1d9lK6xDCTpjZQ5bzp38h
31Ppc+qcrnaQX1tmwGNNsIoIDZ/c0HfB7wU+kyVnQTd/752yVVmmlI0AiWj35PoT
ng65SRnPRrXUhxtjJ2G4szfdtsil4FFlnAENpOBlghQV0t9YQb8VsAgC1BIeTYJT
Y47PgJmdzh2RZhHQWKBb7B+yL33J79jjdbq525vBsQDqMMeOe8mvh/bgccAvWpug
u/XsWFqJtI0K0jDq8xT21xYEAT6HSTylmJ8NC0L8L8RGIkFQQwskEJSR9PNdEFjS
`protect END_PROTECTED
