`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XjzK0rIY2pyE1ggb3wXUCXVzn+U1PQFY+oDZjprEXpOEWbg4YKFOgMZo+WTt/MLn
cCCKEkMm/SOcF6Ii1ObULYDvvnjOutBnZ8AelvJvo+nqeOBe5vTsKtW8tvRAzXHu
BiF0YJ2bABNxZaf9DMaRdmATcbPedeoARj9AcDNSKMdKtv852Rf6+v+8YSZow79X
A5yYIHUh9Wv/3ugUPparPopse0XYO8zVUvfn3Wy4QLfm49QrsLUKVXTggDkzkZZC
m9+JF+3JQNHFxmjweDLBZ8Jz0OT1NwFXOkRPYeFL1hu0GRyIZ5QcKJpmGN9jPyRZ
jycNwXuYILTJpQz/IWAg1FhkGsbHytJ349vgDfim8Rl+WZh2hBnElKevKT7cUpOi
6EZHF2kiT0taau1Tp2IfEzDcyE8d29jESu0N7oddDVYidc2A6RLhedTn20tS5Woh
wOYM2B9mS2lRx26RpyXOQnVMlRVg3h4gOowjUCF7ktSZS2YxcZKMCOyc30Xi+afb
Ipc2VJMiZm3wB/MfiE+JY+CeHgZsY9DyifdkzpmHSOlnD3QPM/sql32Ej6c5umFG
ZmXeU1cuJhP6mEkXOcBeB7sL5KLT5P0mKDOSXBs4DaG9TE6ydzdMO3biTy1LMzrZ
yJfRYJQk6dGM1D3h26RIfFih7bhhOalZ6WcZhxSxKCrVtvyNAn22PgsiLkbY06os
jO5FwfvR9CDnTnAD6V9g2kHtid0dZQpd3kCXywrPc15rdzGQX8/tpJ0KtqDBHU73
eLFNtKbifxIZxGqW3K7haQISXOe4830875701VGhKY0+66VyJjoqKnNWpZbWi0Ok
TfmkUKOYRGyjWQe8K8b5vk6eKIrR7oFJm5RpIwyA1Nrz9o7I9zQvNkIzALehrd8D
Sj+A5xb7IdVKzZOZVy5yPNm2bUK33SnB7I83Tv04+VOoVbOOqQjrHf8rKGlLncTS
WdzpPE9jXvJKyyH2ST3giCEhdtoYJZyEkBBgdWtC4jBkA8yvIJO1YJDPuOfHBVO7
551Wq2ArQLRWzT60cMOe6eVH/l2Ynuo2QommsFNXbz0xQs6W3gMvBgTNrm9huUqL
E/HhPMX4y4vn4FRWMwzFiB5z2fwS5UBDpS7GurUUj68h3Vvut+Fno/GxNeAy7MCf
hp8PYaULiQTWJYDnbtU2/b7EyIMfKQkUO3qGrGVi/G2at02PSKCZvXAKtw6CxTe4
eKhczoExoz6bx18pT9hACu0l3PpMw3OSIevn+Vv3Ejc6khYOK6J3OKydLZ5tYIuo
EVU8v7ML9wS4cGDsXrILQ5ykxojDk98KLGR+UeshJdN/nzKXCcLw1/eSxg9NihP1
SdbaS0hA+GeSWR2s9+kzt2uou8vBJHcLQTiI213T7A617PKxbZT0QIEfbZdVS0t3
MZL1m9vsEAUo1J2xEWZ0ftUt2UlbptSTGpXesMn8ZU78eGrFetuK4z2rmD9dlmGA
/XmKi6HkmLiC/gp+u59aGWAnzB/v65aqWz71c11+SCvlHOrFXgGlB9xCmImU0x+u
ERptf1Tlby2UP6rQmW8cw94QSZNlLR1IiirPqxI1p4U3ez2FDzt7Yxwv2Q+GKH7I
s15rG7la2qbnKSsf9e4exIJj2zM5cKnQpP7HQxxDDrlfZs699yL6aRcRKvjgyidi
JztrGjlqguIrEP6k/iEdFf+2CstwS1/RXZxK3fITzRH3NMFPeOCoiIV6HMmXhYbw
tzspMGWUj6uS9w+BlPAGY8Hrb+zaLcibhrQkzkzChjV7q8w20ZeTV8Y56yttc64i
KiObDF7N7S/c6ZZxorsape+NNMS04fZeJiumNZfLFQzeaC7BU/OwFQDegGWWB7X8
K1wTBlQAZtwkPySYFLXUOejK0iDAu5Qifwaab4oCRFnEZd+Ya1YdCvZ95r8cXXZK
3BWxeGuLQcOSNAF5aagPou9nwCWKA8pCvjHcQmfG98wU6Wa8XK7ZWwBYq9UHVnXI
gnn7QIz8F9LWgWIpa+LaiF/3QcKZm9NFIqQossmRAAxHKyEYEUObRYTESQC55USP
MggcRBZusRY6DxGDV73xYEIhN7nd5tB30GC96xTr6NAb5iI4x909TE8IjIzpcEbw
mhVfLtZqW7S2sjnMVCH2O2+u3QURNNdvMGT3f5iCv3dla3wfvXD+yOObjXVvjjCN
S1hD6VffkvdPTNxk4OooBI5mlVn5hmBxloRwrO8PO+2kGL5psW2BiAZhsND1D2pm
Sknvfs5De9d+2D3XYXwj2F3Y351ij+wegMPvdBaPPBNgs0st+xvqmYcEE+sj9KR7
lJ+otSvOpFat/NVAVrgLVDCOOVXPJTkxY3IoZ9PyhYH+JlxSKoGJ6DUgFEd1da/e
mlKIScWSQPB6TikmyG/32yxVA1RvT7ayIYKSdUXn159KiZtYAp1HXBKlFfn3s/rG
+nnrlsRdF9qyHKb6hkubRNpwFUZ00gkA+t2OM8JX+KlBjpo4wA8gadGcjzoDOLo2
usiAbix47d9lvwTlyZe5WS/mE7q0DXH7aIY02fQRH9FhL+d6ZeAqnMT5nJ+hCfdU
gHSO6A8dk9p7WkWAfhYIHEueGfsn2Xd2PY9wU4yANYtsH7MrtFXkAurK1aaJF93U
EZoH9CkckZSwn5UMzhk3mNELDCFFRaXmc/oSM57kfoIYvLzpw+nkQZm4sOE/YLQg
rmEkJn+y4QBf1Y+dRTtmq97nzwfRMCzV5pEMGL8cJizPznh/rcKGWC0/fJCUEoIh
/sfW9zANftnOvuXrjxJQTfMRVhHW305c5pY6OcGBpyjX4yyecqhA7nU9/qx8uUFq
lfxISE5cpLwGpvkOZ/jWtkvEiG+Ppop7oa1247W6FxA=
`protect END_PROTECTED
