`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
esLtX+BC0x90aC9WfTTbzJGzmtrhX9w6zUfsfumRXLCfNcWlwlBPdc2MVA2yPqn1
gAcRqn6OziMExHmWHDISC2xZwRx66kWxJ2yIH0YKsWIrSuG7CzYWynpLjiPSCjoi
dhicklj8qSRz+XhyEEZlCARhGPSUEoA88GUNQMbYHZZypn1Mk9qeimFbUwQjN4Rj
XiA4mJOtKPKUk9AgmUJN38O8FQgLd0Wcyn6ZwIgaNMP05/HnNeZyQ4tcb2XAjCWq
w/wjJT/d0IvT2eV6S3JB+v4oLE0Q2qOBgv65Aa43/eaQ5QmHLt1hK0pYLRsWj41e
gLoeks6EsAAMdvwsNmoDyiKIvPqM0ca9dW/3keEyM1cZPm60GKK5KdDfyapgg+ru
sXdLU9ekcWBxzB+8B/q8ngQ2O3flPiCdBOqr28Wwyanm9Qxj60yE3Ak6WcRwNIi4
LqBmhVRnKil5I3+wjVpbc2wJS25XwzfHJ6nOgWef+wZtySVmRCa71mTsVxLXVcjz
`protect END_PROTECTED
