`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dBrNzzUCJKKL4sXeHsvtfve9/W+d9e/4bqJNNSz609KZ4AEHl7WVjwQcfqbHzRwS
B67DrYWbML349eg/2aSdbOwQva92x4cCh+scdUlXCpnIrptP0dy+addIf+ppRnJZ
SxYGHEJOFpgc7cld0QAovo/25qh6MV5Nwt2lNyK5NtIweOvo8siv3F4ZJMkb0l/q
RpCaF4SgXT8BVeIqri58TUuvfTMZ/sUJLf8/+qBA7gNG5EerwdUgkP3kCKcoKM9U
1BSIek8Xo0HHEAnJBUk+D66cxLli9SYOjR3jSbzwUP0H7PVoF5HW5p7IJqXrOlgv
DicjkQLFA3jQrSX58MxTxgxI1SHGMBjlEcf9nIC0TkhrHmGKmGqGPLQIrIiVTij5
tOrVJw1V9aR3+D0Hp+1pXg==
`protect END_PROTECTED
