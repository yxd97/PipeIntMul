`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GDYVEy+Fvdc+wmVrQsqH1BsPqZBR5bIKWDXVal2A1rLMzPT9CT2DoNXobjy7udb
8j89TGrp1+dkoiMLQqrKVOxcDuKdkr/hUvPVWKTzfiIy3SMY3bhgTqD7AjtMdBAI
/oQZrftxBn/DMWDaJkNSSvH9+6nn/h76iQ6d+QnQkoOlRBeoZNpFFO6CqDA5pQAb
8y9BRCFpYxFJVZ/xCLwjOrElQKHdZlRuGU+RHYg4SETf57ABu25hiyjN/OTGqWBE
KBV/T5du9CHkdul969pmbXllmTUc9jYKaNQsO6NdiODFdSUJNFftZtFuXvf9QkOt
2B9bupDtoTZ7MLOFHPdLhwi1M3LVpar8Ng/w+CKiW/p2NSifXNMaV7I4FAdhndi6
XYzciLkrwNQgkmYqISrGY846xm/3d6aJKI/n561DH6yYzVM3PxVfnI/Bq/GhxfTA
fPQvjo/So3Oucy6n1bdVvRXA6DdxWCGX7PVjm6MiM1bNNXNWa1q6wSBECH6QvKkj
5NUe52IRU7vT/ndFXWmR4Tssp9pGXambZo9YIeLj+5VUqe8ynpdHh1z+mzirnMmV
V+MuvawVTL1B00l5rnGeO1Pt4XorwHIje8C1qDtdKr4TV314MKORF+CLw90umTE3
j0Xgjp88Jwq/a0AgzS+bn4tsE5MH89VWIPbdtshApdpYqiuVhhlOcMCwWdwoI0sf
aki1YGmKhQZTgupgfcbFMy3xjHWOi5GbtfGySh6i/zF5bn6xJuDR1Rx42WFupvsJ
SxkuxRVGFYMczlsBNV4shejMydXMe4Hm7OcQHSGNCb0LCO7Y+mElvNGwAqVZkvaf
YDfRhtvgYizYYTjHhHDJvdTPkrlKEgszq8odInT8paR+OmN02FVO5BUJriULw4RH
RfQm6vfGx/iBfc2xWqctfJkBrAc6y6y1iig5oCoTIs6CGovyGf7qvjmKalg6Zy1d
hiM/9XvyrWK4rmMu5sho1lzRTBmUvz+yNlG9eNU2/Utl2WJLeGarz3nwqyJY9Ldm
irG1+m+B6RkGf7fXYkF/cXNz01YLK4RhSjuaudKJoNA=
`protect END_PROTECTED
