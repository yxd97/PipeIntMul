`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
daGJpXbJweAJG5wW2MeVnxXFRuPMYxdIUMkNC0pssRCM6/F45f4hAKKkz6+RMajW
P9pLE3eHqHDjigSDoYJCx+Q9k1172L+rtnGK/8T3gqrF03Iru9y5mnf4JdQN10yq
Gr1r3ne5r9V75Uaq9HZxX50fJWletAH5AsciCvFU4y+wpJm+VX5knQWPICZBOz//
iYai1DCVqB5BQwbU+jWHrW7q7oLV/eGSUYcRBzmpyLqhjOQ6hhyFmM6Lb+cHaudf
W5G8USu8G4vukhe7kvfCTZHOs9EfPsY/UXou1EXLhhYSem2I74NdPy2CWWAUgjt1
ksK8S9E7aOMQwyOfo300bcOwKKD7wxf8cmUSAHOao6lt24Yp3gYuatVTXiiwTqPr
PIWMzl4C7gbMygzTCEVeF6uIRNdTvh2Gbkwid6QJ+jjbOfTTmjmKMcGgvI5C+JZX
+AsmYlXkgxt8gYvlglYc/k7kqKYVHPSElf0yZRmQE0YqtNmPriJM+2HQ8xo5Gq6x
oZsq9Ajy6/3r7jhVEs5msBsLGizH/utDaGDWRqaCCyH/jLe7gDqPeFVr7TrStDYS
xe9Y2WlvthAmRupw4tC+7R/TijzRpavkebBahAIpRgkH6fZ/O2SPQghdhakdm6Fu
pKxHBC/OUVWqyb4EAZLV0Us/CIv8GYy9GCa/7+7cO+sUdIKO6BNlPN3xJkmBcRyy
lk6gp9ajr8juPKwE+dLUoBpq4UbFeEyNBOoE2i1W2i6T8Uk+sF0Z7hnoLxIrRzHR
niShh4kk4qGULncqB+X4hBWGNKWT2iHur6qfdVq+Si7hSgnpxsjtP+/RmuK7DNJ1
zU0vlVoNYThpuhv7mXdPsK43+0jrCPD60dTZgzbr2hxYlgoqzhrrawKpgnJ07H5A
RvYjh7CYTEjYB+sHDJyBv7+w7znPIs83zjQ42JKq4/6KdkgCHi9IxeGZPlggYjBP
+EKVha9qpmN2eOexejTQIMYomEY4Uc/HqjYgtMPUZ0p0cHLmH+YJuUQlpFWXPE5G
Ur52M8g+88VB2MKeeDDBhvmhka17pVA0TvW/x9aNQI1uXEXYZuQGeYRJSKhbbbVb
DjaUw8WkNNrikOAjXg2AWOvFQHuvzCG9fUPOveftK3l4NzAeJxtJIIxbLxWR/pTH
/Ciau3lCBtcjS2Yuua40psSp+ZTRQPYn0dCwZ72Yf0gz26IE5HL7tChS7r57ukrU
9rUpSSc+ULioKgKHvmTtOybYrf9QEhyMGHKQSMv2cloJmIwKIKR+k/E4N82jScyu
KVoI2DxzKkiC0otpd14yutgwMZ6m3T9X8BweLFg4o8GXPBit4h4ZGjkXFwTl/8hV
PmUw/VTWwJqyl6i2uWL9CnLDGxM2xfX/NksPFSf4mCE=
`protect END_PROTECTED
