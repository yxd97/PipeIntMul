`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8O/lt9wpmi4GFn4oi3AaRvtdQHazwP1VAu6fU23y+LWQWTsnZcBSzgLVSkzcDEuB
CpCAiGO7oq/GIL59kzj6mHqR5SjoJ5yipRbKdMoLT030E2jwzIOcvXfPeyIQws7Y
CFBOYwPrMmotNRwUoPcg9hMXGCD5jAtgZWWOcVS+tB/wcTOgeGRzrUrW8NaXojec
MVdjShOazWLtkfnYcrONniSyEGha1KC5Jcv9ni87uYQU/f0Px0269GZb4XRWBfSR
wHArZPqU8CDdbSQO2zYmSoUsO1rtnEWNGUCnNYP5wmQyaqx9LA4P5/FCWcdlPR+R
R9vkO5TIjBlSYRfNO+QczzVoXPTrzRzqUM+OdGgQ9mj2wt8/Lnv/c1e2QRYE2MDG
DD88Cd/Ft7ohVahk7ao58YqhiiF4H2dJj54seejtCkQxBr0AyCkDE1U+kedIlMU6
D+38MMsIHdFN0ZFaFlE4/l7ZH02StCiO84SlahKKGiT6j6iH9GM4WUllhz5BY3Fx
lrZeZmqEhhAWsAU5Fqg44nUzgiV/AKfRIfoBeAH+Qwnm0fLxd77SD9r5ZTNYvI37
UspC0Rh4XHhWeGkKunOFDrUQB6LF0fxfHftJuIJay7AVPcMEOLA12eQmEXPjGpgn
iaMKYJPpizlKZ/rb/itPEf1c7MMKu9LRdiOSEMWYD6HFwuG3VUNOVzztuv3XOr30
oOiUk4IueBoeJ7vgrVICxA4AxnUpiaTlI/EhPZbeoy1KnZ6iggfWG5KftDBGtiAc
x1FYGn+ZPFD5Li9DdDgojukocfV7N857L5JMdSvj4vblN/pMd29jSjfOVdqIdz1u
cC674Hb5Vmri8gxPiLaPJyPZ2q+JmxKtkoKFl0OaWE+a6tc/dpVlOh7ZNHNaF97R
rBaR4wGhnYJSnXWzG6mHZXGyAXmd65ZB5oPIOvlLp50DWo2xZN4nGinLs/h8eBsd
WvFMIm1VUAscaChW9Olxrv4ZcYX04u6YH5R3aaPQ2sdAPNOn15zeBBpdWHDKCAd8
fKiB5qwmblJRr3RZYTydx0CRO+JTkcCaWfEcti0u23tzh7pwgBKCrNmZ993fcuZS
7mahbrtO10AbdZnrVXESyxLMomJsRFCYxaSbVnD69Y7tN/OWcYCbfOHvcZeUrrsD
wko3219xobjj4mPK4bEX/Q041XqM53mqPLXolWQBIfVH3lWM66B67NO2XUNdLA5g
fg6S/UOM0sztOPfn71rO6nw0TOT5+piSJca4dFLzFZgsiwfW0LSvhWLeEYEey2go
UkW6/MEvQYgjxvFt90colJs3xhNKvuCjl7zJFpYG6SPWXS1o50aMWat7iw3U+yiX
WDeq06RayVYHEjFCCaXtcM/tpR2wWKjOaw0P5JO66Typ+ak+/srGNUUDsOmUC5JE
DSQY+oM+tGI82EbeHl44jMDA8to+R+O3abuHbyxrfyEvdFZ8VwebUDrx/alOGVjS
6tGcA1HCGhHUS+8kUhnoAgN8VUsHbZ4RVuRCNVy7l9IgudqDvd1U8TFguCN42+LW
a9cX3HDG1kN2I3D5VEfCANJz9sIuWOqEM/CICy3DCx1duPBJuvr5IK4ni8mjj1KZ
dabcS+e6cB78Ew82XTmrPLFU40PvagLQVbnA1rOlh2GFMx+/9XjKCnBG4B5Bc3hv
GKUYqBkIoeLq32chLqaCuHVRjvVSSNoUVnCn0bZaASDqLYtTBzR5q4tT61AKmNm4
MBbHteb4cwviPEf6t8lTNtdBpzpuocMMPVteGArTq9/mw0OCVbab6HbNbOEoN+O/
LhVpkN8KqSZ8LbHNwWXSGIe0bmv4RKEq4x0OqO3PnI0zTFRbfjxbLlNyBfSd/Gjg
6C9G6SmOEOhaDL1q9rvgGhwx87vmqt4FfWeMHAVHsWWj18hQMNfQdhG27vVpe3+i
F1SQu343EkFX4Jo+38s2fimePW5OveCuN/u4oRu+xmPZkVviz6ihePsKFWiaNEVF
VHFdZNQ3Q38MZ79U917XqJB6rJoKP0/IdIvnPwcvUyZpcdLDDA8iAZA1Q0pWUqa0
66dbKoIlbVxS1VIgm8C0lvqNRMVeBaJIW9QX4N0EDRypAln7Qhh9GYRWUnb7IgEo
1UN3MlDXJ/PWtHupvN0jUHcyMoigNITLmLGoysWx9vz+OT1AOwDRO1iMFViKRmXk
U94OwaoGuDP+JOeR8NrWhDKMNXlXOlM6y2ql8CLz8crzY/dgfd1CR21Qp4nFD1Gq
F39VfZJ0RxDXfLZtAke1kKItMSC+7buQUOvCns5aaUQ2OV9QUAgMEksY1NZ61gSQ
+BP3Rcu+PvTF5s8oh9Mtl7ZEsgAFKs8BEV9bUZuKLqqecVmIZN8aVFf5tBcO+WVy
8DImQEMa+FkZYD+vY4j4Zy0YAytia0Bp2WXlEAwMlsF3cA37ZpNaZxXDGARdx8nA
TPYdqraq/S+Ui+K3ox5oM/XX+GHNMyxSKGx4zlFwzd+5aoF5i4ghlv+6yI4Lpksb
Gtt/HlBKDwzkondBzc0L4PnrsjJ7j9ZlIuXs3ob1FUh+0iuHsoRfLJvVbKfV8Qj6
e3KQXxRowyZtiafcjyMdQAoThPL1/7AFV5U5UKSJ7X7c9NH4ZytLSilR2wgyVRko
sXW83pd7/pGG7gV8b/xge8VjTJ4igmv5Vwq12AQNV3H+ZI2z2cpDEL6mdeoYuRLw
iHccBTKQe9VwRnOK0rQdXDOgjy0GYQEwoB9xoPgbaDciFsxNDDDbaUSeWFTLrGdW
PgEGbMY8rqeF5oEKv3Wef1v7OOQ638DnUdJjkRWKf74qyMs84g9AueV0s1NWYkzC
h9msRh9IohlhN5KQ7nH68MRUcW7yalUQBG861WTC0SVJHiGkg8JUStJ741fKbYw8
/0JEX9jC1mYqVcwdEAOxwMC1Dx2h+sSdGa6O0FwVjljYzXTYjR0PwFcHi2LxCdhn
Y6Tfe7ovoyZVpCP6dAC2jDzQ2gNNFd+2hJwVE3XNgVkvghMANAEMXn+vOjoGQyNn
JIaUgCaYs86Wr6eRTbKtqLNlW8x1KoFWUnw/QAhYHf7kshKBXiEwGEv7kbr3jork
25zHOSJob2KTqLIDnUYUxfXekbIwkhnopJorAgF62MnfbKiZcl5FZX5JAEhH868R
nf0b+DWsXViWERWRvudgJz4bA6H9V26DxkRUWLrmcIHwr3awyai7gyk+h2zNqAfC
gKa0J8mjkniCwFszsn+cW1okf0QwyBm0uGlkIZ+JlcJ+Ro1m+c7xBfjMF6rb2mDa
JImUZijyNUvUEx9AmoJvxFR+qg5fIuzz/WAORCU0lDR327yhKgk+mo5yIaNLrD7j
dZG94Oc1DvoASfDBURcwAAGOcOpAtubKhCT8g1+pu8JjVdSSHnqObJ0uz7lXtvVa
J71hXkSzranEIAvpQaz5yo1UFKQTEZrjGZOwj65giLXhiHzpvWkJZ/8ccClRKmHp
m0E+zhbn6TytoNWRmHg6DCQ6RQ8vpjheGQzUjPvmAP32g2TsZRo4YKx2EjvmPe9d
eQh4RdwUTsp3PWHczY4dHDLjb1Hy252CrxY4a6DWCquzJSiTyc6jxKYWv5FIoPzU
vNAadrleN4NP1wv/JoAucsHL2+8wW4qs9nMG0UrVkasntsY6UbEOHmolCzkRoEYc
`protect END_PROTECTED
