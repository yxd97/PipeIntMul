`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aj+cH4NIW0MnNOIRw5qatuyhFZnrt+43iefsMsReeeyRGR/MUCfyzhXnVxBNcoTJ
p89YVeYzDe7JTJeKMF6T6ReiHFWNjXtShxaW8LfBv0xt7SIliTRs1eikDcU7jRpb
LKJAAx0Zi7r0FZF9OD5aimMxBNFfCaktuhm01UtYmZrdMHhH1+zvHXJbXTYChPO+
cp91MJYysTcJFidU6ebuxLCqV/vAaKsNQ67mptI4Qnf/zulN7a94DyGqQAgwAKQq
RKIkXymA4fQjljNz9C9pX6ZZ6jWcPyYwomHPTo3Edsi+tdeqit3Y/5Xr8P3kNf6c
QGNByAWWGoUjzX3k2PXdcvbmdWIYIbXcyzvmLcStmvc38hi8vZDTdxSoHPwQGgE6
ITjXUM9ILj23Y/1k7tESmN7vIXaqPE5Fv4F5B6dVmyZcF/4uSEGPWoeA3d9fBXjf
lBaRSrb1lHyq3XGpnJy1KECxdrpKcGT+tzoi8Mk5tLO86zHI2BzzjjvktV0fSHZd
xyDKrApVOJ+3HIAkPdDOpMhSStMSwPmmGQXn/7pqGdakHddCVEmsw6qi0gHtLOE2
`protect END_PROTECTED
