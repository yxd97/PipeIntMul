`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D7TBg+6X1BVhhmjZDBVEbR2vjc9zcCws4nxIwAB3LbEMJmR/81pHlWuzclysDfKw
tynjy5CvfRvSjaO+y65Cx5IsQaPKhM6mcsYhkx/3Ck4hsAxdbkTt7w0EC+80RQ9u
GG+c/mVTnxHbO31q1VgQbFHGT9nXU7Pzhl58rOukhQCqO+6CLiNGPty9mjg1yMdJ
y9JWSm0pIXIbHS1stavoOciq4Pg+xPa2ab/Da6u/P5Z9B7aIyj9ZE//+AOudFCoZ
G9r1JWSb0smoD2SQIMlYW6ebOkasyhkeRt5Hu23Klp8T8nx/ybOQI55sgBBQfy+A
+QlICLi6r17+NJO1OwbnJLLjqBitxHnSlB972/WEjN75Pyb9y/Lugnzt+2ErYcgz
/vjPm1Ii++hC6GcJB5aCoQeq81wRUqMUveJfmQTlm2VNkwH4O0zP9rS9mEpw+daI
`protect END_PROTECTED
