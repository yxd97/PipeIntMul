`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XrjxsIOesQkB48/mM3oXU3fsAfmaYAGXSaZ2B8PkFNO9F8vItb5+QGrecFkfEhgO
BWrsV0Ws5z0u4wP69b7Az7+n+QJdO0dVqE2fkbNbj82y/YqvKQWsCMBsy4fa47iP
dKKgzY04cIAinlHI3Apnet8W0zX1Hn8l08rSrwhpUc7p7VPa1+8UFFxbkyIVr7nD
mNKr10zgPFigUzsdRiXvpxxCHhdXZnz/qEbYsce0isaMoh2lD4e9VCOuUJRbtPcV
6krZfCADy1hmMnKdW9EfaYWv2xVdGtMbGid9sjy7Zkg=
`protect END_PROTECTED
