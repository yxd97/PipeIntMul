`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/5NzOJwFOn319id99q3+4CZzdZnYgAwAo52YdF8yKp70/LX+/AGEh9qGgDB3BHqM
MvfLRZ395dBJ19gj6+3w7/NCyBQKHQVSLsBeSkRzvRjZc4rL0+6R9NJ5xLorQV0o
KsOq9bgK8RTRCRfx1q5TuY5njXWQcee7s/ILfvKpdPhaeFkdSJ87YAlHxGOAbTpW
ujagkjO7d5tB9nquAHrV0yO6ABp4gOGwdI+jqjoiBA3wgKGu5oUigFn9pHB3rCoW
MZY6/p5CCjzw5XCJJfzyA+64ti0cG8yQD8qpDZVUltSW28DCf7a/QGr8e/PuSyfC
nQ1PP3pnJh8IlwzmmpnsbATGaYjdJ1SseQoXOkueYOSAH/PrMa5qjN+q/zVXJwPJ
mhzyJRmI7myLBKilY7/zHh58tRZEfANOfYqqLs7Vlr+qg5nFbqe2dZ6usfjTDv+t
nCG5llrPvoa63uEYBwPsxaT+V7AJSW/UwcIvWdZBp6DPVuAqIY79N9lVFuHEwx/L
vlZBRbDUJdbbCBcCDdcgE20/9hKcus/+g8LttsefxWtWrqV2zqEazNrln5I8mzcw
aqzEesWhpakCAV8zPT5ViL6GfVQMuMjUFuB8pAkfoDeQ2rYtyyG5DQOxZnrFSP7h
a+klgvHv9Bzno2JX4gR/nJDSmEwri+4rWOQDWYZjG+Pj181i7kB77QIZZhmZC3kU
oJQ86/MbMByfnM8qda1Kce7vhbT/ld6CaUAfMl9M3SLWv56hxwuPRfSM537pjfcq
VpFPFvs/D52fYTPM7mm2LxtRi8tApvyOA3nLKaDFXQ6jqD1uiFGZIyalgKDWKJW7
TZ4UD6drz9mTqM7CRz0O6AyZl/aFz5gmLNDarzbaC7oPKEJDObuiE7Y2gtUst+TT
G/4ARqeYPLXL+RajFR+IbTDjgt2JQYQnFbSMq2Y12B7rpAFZ1n5BmrhtvZRrG+bR
cqzsBsZuoozWC/CkgA1xMqroLf0QfPxlJH1UbsBOboSWUrcx1buGns9HgX1Ec8JM
BqwMGWpk/EZQNztbQWPbJfL2dEVFLKbZhoKaXL3d+LWdMD8AcEPhoVHDykRkVxKK
SaC7FUwz/AtdW87s3aAxbnL0yQnzZwklOvR4QBT2zauPb8srxgl+pHaZhznconL0
UYBoIUzD3hE+RlEEgrv/QuO3CL6hSi8kNDtlxUY1H15hNr6TpG6C8O3c6kTkBmoB
+KirJGJK32KKfqwubyLVqfCxEFwlnHGruO0z/bU2j2tXz1ea+fbptk/fit7eXGY9
e+jUoIouwFPAG9m2eVThvT3o9b0QDbIho6NgKphX510tIira9kPyWFC8BXil1rUe
`protect END_PROTECTED
