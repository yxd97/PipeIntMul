`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
92VbD5XQnzaftoaZdHJLNUPTmFjKdnHKQOGZbTszRyy2/YS5CbRtxse0M8ajwQuj
AioAVQTLpJWUjBciv+l6V2hF7MtaG6RjcEBwqnaUrRJ0V8ui3V5S2KH8hYyzqWM0
HgYTZrmBzTeTr0OaaJy/GSuy3c1g0tkiCjzi6O0/sUiLI8n8/BS/VyK48wTtGeWI
HQcL22Hz5rQlGrmBuJmR+2mTVZr29SXGhr3KrNsG5lM9UU5MIQWJ7aL5ijf0LROv
Mb+tmpsLM58hiElN8rRgYzUWhbqxAdmHzMg7iTrItYw9F+kJekml8VWCSdH623+m
/4aQLHGOg0HI9MT2rJTLDFSWq6kmycLEO6EscBBJAaJwtrvbDPZz+CixNrX6MVJ9
AJtFuI+yatL/rnoTkJazOA==
`protect END_PROTECTED
