`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P3+TS0ZamvrsYE9fM5Fm/oBuD5QLbpI57P+5PwXcJAg5K+wic3ZlCgvfiMgx7B8l
bVH7Yqr9SLXfWrQ4VXpE+qtNd5waVK/+8a0k09xjFYRYC/MMlJOr9c44B3Zq8F70
BKPY2MHYY3Sd7ZzVS5WFjIoCpA5yyKNxuiQA0vLN1QVZB/lhIQ3YXj2N220zRvPU
uc5d3lcbgRwgJSI5iMhXNPHQi8T3BLWZL0pl+sFW3vExxAW7Yw9G98ijM/KnGE/j
uLtH5IdNadpjm+FUvBDlFRlil2NLAbz7ehn4R7tvJvoS8+auURZe73UcOieZT75H
T6JaY/Tggj7YbgPvoRdtBw==
`protect END_PROTECTED
