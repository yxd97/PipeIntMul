`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POz4mf1mDOdP58rga/aC0xC/SVNcl+anQKlx/zipcJ1uVN5ljrGIyWg7sFf4LUJo
evdI3Ake8BG8JRUWZg3BVMnjVeyMMPIXEHWyGO7tUDM7FcgiFxu62CJJgH8MQ2hf
YZSbgI70fRodmugqB4J50eVIkaPFpdrzP5UwXVlnKDseVv0YjsZA4s12LTXtPjJn
LXARnX5TOg2GL0MokjwJ51jg74IBNysfJxWhI3yasOHzx5ZsbMADDaN4ELdzVQ37
/Cp3sdmIu/b9xaPG/a2k8AWn6t2FV7Xaj9VMTGNWZIuw0XnregucYIyF0fbbYmVL
sUmkPK2Z6POIxW8oMjX39FZxD0r2z1doPEA1VmsPulmX9vHbg9S6HEa0eWRvfnwx
FikQAMrjbu2F8mIb1QGHPw==
`protect END_PROTECTED
