`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cayrbpC5/WNbU2EXO5/H2oGslV9fErbaBrCMNWY3Vg0B1GrjZeHYlOZJPrkKjCgk
97CbVUlrSs5GHma0O3Rsu2e10Uz3KOGePw56AJwSfNR4oKsmZRSfCzXKP58gh7wi
9Ikuh2e4y+Y7H8G5pQjet2eHzJObilJqj85QEcmhlVn9x/En4iN9PsUoe7+GuJWK
jZIArjuq1NPv9etQb2OsxpqlcgvTBS2RhZdSIa6nAHYnjrEnSSryL5Q+9OhuVpWg
gTlzinDTFEWtzi7LF/d934XNv5ZqBUT4roFTuFMF+CzDoXzmSyUzmkYFLTWAwZUN
Gp8dREsBPNgOpYLJ5P489qQfSHqqBw4Tn7CxIc67JmUa3by0WyOap/mGGxP2mwZd
An+mvwJLPjwkW+jGpJw8NIiNCOZtMYdBa+5vnOxQ1O+79xdk7QxpA47+PuTwuZRz
LdFf7swwDqU1GTgICU7Mhzs/Pf9tXH2zQ8ppk2nwbs8=
`protect END_PROTECTED
