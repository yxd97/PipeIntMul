`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RZgzXlDJffJQFgvK+6C9yXnFiCrjbmry6ANRtnmzOHNxJuyVFXZ+I7WslJWX5lp9
pS7dfRIdnnkNQgq+YUq3gYLyBueDylCqoKi8dC20EK5O34jp+BL40BNNSRA81svt
C0AUTS3XjdBnz3uf0TW5eKthx3DEA0l/CMbsI+X/1z3i9TWMrWN2qYGkErsnFa1y
YaRQ2Pl7pxuUNWCIUWqKqVnl0U28P9odeKMyLSnpc5BDyjg3Y0iu32LN9tqG58o7
n4fs5nCgKd3nUN2u/YepLRdmr5KLVz6aTUOL0WRiUkKA4wWzDvvRghEbzizTDmez
yGH/MSPJmDQmBSoQUH5dWOu5ufTp8TCcYSK1KQuwdSlqtoDTOYZdenY/iSuUtBJ1
i7EaxjCNpZsmIuR+yMC5Uz0cRzsAs33n5R+NNWkAMek=
`protect END_PROTECTED
