`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RY4fBjViyVdXeo1eHZXhJrvFYEJNdGx5HZDTWZ9dGkffXKYe9AOouacmO2+1gAt4
u9n1vG9VKdrK+68XaNKNbr4Tk7NV7yyScBMZardmb7IClyQVNl6eq28XApv4Xkc9
cwCbnqgcIdB2TMCqLfhcKEZwm2P0uHYhTYrigN7+uboT8kKmNxLFiZqT7X2lFGOj
PmpUxxd+9Czm9XxglWNCIlwLnFMocgazkYt1Te3mF8DAOG0yMIqxZnqzEMzPXoDk
PureHjMztm4CAyu7zf3tW3gYn5yUFIHPHLY2+IwaNU9bKaAAHBJD2MSntkC8YCWU
0x59nrSHoAImqmOcDsdDxLdzbfP6vlsdX7Nrf2r64X+1SrctAs6HnI9ouIvjxT2J
RPnFi3EEP7ioph1jxR9Jbeb+HQ3N44IkA/lU3AOYq1ZW3bIGikE6+Qryl0f1/aUg
zDSHXWz5CYOL8Kb2KUsJwkt8dRff1Y5QwiDg/XNLysTHw5w8chznzhYpyCiEnN+T
3gPISfCSoR7dg35dCLA+OINZeKOyFnFfdd7aZd86gPCWVAtEVxyNvv2nUkAfdT6j
`protect END_PROTECTED
