`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IaIrBtYzFS1MMvi4dSkDhdGUkrHXGkpJCfMrb75G77whljjiyHKvSun8ifUUkM/B
fSz8ljgcaANRm5W5MAdSy/KGvAiYiVEqBk/KiSkoBuZ9enkR9+RtOqx3nKHqp7dC
vvDarSMhCzvGjOYmjoKl+SqiU4SAp0Drykdml8l4S5rLnaPtH5dvp6M01sQRDB9I
1Gp8qpc8wD+/I9KlphCy+FbVF4cEjQXq6yk7l4lGmeLDeVasPOOZaz5DNGhRhsIN
0XL51Ot3woHXoElLRePNqOs8z7V36V0jo1YVkna+FRj65HcoNJsqpPo328mQ19+b
yKMT+dhuLqck2fEYNg42yw==
`protect END_PROTECTED
