`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UYgqT6LT3mLej6NIUrxfW7hAqyypC2AzW9mbu3jO7cVvDu4oTCWZpphbluMy4h5/
gnW7c1FSaBpZUt2N6bQ4u2g6dis3RoJrU01/ZoQjLhYD5wSmd2Dz2j/uIKo5NT3i
0xckrrcpHdBvEk8lNy6ndiH8vjiq3YRQJdQVP2G62rc3cUEh6a1zsuoMD9OzlZo6
VwdHANnilpcx/ZtZlJxndw==
`protect END_PROTECTED
