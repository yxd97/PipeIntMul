`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A8XYkMVxEGGGHpn94tppkJU6Q2+FJNdKMcGY929uLW7PaJDXIeEH32f80QmuUNPk
FNcIhciUB1IoYbF960YAgH4OTwg2zV+ZRh233wZkspqvQ9ZFpxXTGJxoC8f9LYXz
wdK5dNmoPH7fMn1+WXr+fJT6rkwsmzWw4EF4RXKVYymNmBMf61wf50DTSPmnGtoS
9wzbXaW/gebuMyZVC66cVbH1kkCwP4rVd2YGxsbLkkPe6NHwHuaTWHDoWtuZOp12
Ft7r7j5ZR3fFQa5WokAm1L1E3EQ4IGwb93WLy+uS7E5gVjdGNKS9kM1G9VSEnv0H
/70+yWrgyyqKLrmJwddGLsBQsBQaHE3J9JVtiTe+SMGpsIBJAH2bajV2N34xxcob
UOS7o2ZCGL/4d72ooWvCxcXpgff4fbYsp6J748L0PZVGf4ojyfzKv5LyhwlmQTcW
8e1+VndaHNsJxeltIoyJTdwmkW57ua50a2Ee/ZmQ1+9SS6UGK1SJTS+ISNaqWe5J
NEg7M6ayr1KFIc4LJNUcqg==
`protect END_PROTECTED
