`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kqt6LSjAH9E6Ne+Osb3ibmyH2IayJZWCTbIP0sWLiOi3kpWzGJD8p3WNS1JEBUXI
zrvYpvObsdHQqAWRHt8GLGThrG6AN+2bOKg4UgsMwK820kxCeIPHdfbGGx2m1Sfz
c0BnK7E5MQ8kBkDWu4uIi7lF+rP9ac+tG4zeT6idPmSBicoDWb2cQsIeSwpS/Qny
OUsOXI5VjPbDguWRMZA7J7OT2gGfCoPWhP3uidSLkQJ+1gWo0qgQdtYBikM9H9fm
RBHlPB3MB+0PNtuVLEZBQ72wulJDDpq5G3uZEjCFZxg=
`protect END_PROTECTED
