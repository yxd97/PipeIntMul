`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jxm7ka2z+HRYm7ox8S0n9roGBrVpgrLs3+eFYYsyJhxbWiW7rjuEhOVxpNXTaNm0
vcWT3+HM9YypYuhiJhB1mLYDkwbJrSRrKB55SJ7KkBhpuIM0aP3fLFcxSURNfmp5
qkE+dF1z/emjQG3rG4zhR5VPiBYine1izuy3kzUJ+ANkerMMG0hVKlMr1WgPpjWA
m5nlIVA1eRxuWfm/U/MaoJ1ZpOhJS9iYGhVXt9rRL/t2wSqBaJ7rjog12XhURcXH
075xNuI4ymrtv+i01CVWbqUteETBLE1CJLa0JkRMK4H8MSibdwi884PtARYfcPIb
mCyyYUeEe9Fw7BvSlpp+EXtS5DYc9ChDzUUOEDUqQ95NSOX6T6ywitU7xBVCWjbL
OZcaycPzehFP9TpjkPyYLAKDnRn7XRUBwVHOmU76HQAaziFsuyZmnGqLSTDVrNvz
H4oRSDQLiobdHYGH5Q0QD9Rn4y57tNU1E/MU9ZqJUyESCbwgNWqF73sUOYnb60vt
RicLrScXzqs5MTSjPOIqRRdAMyUH5COL3FZjln5czgP/YYo3vvFOVvSahSjFZWGo
0F49hP4nrK3YNd8M05kIyi6/O1z4NjY5mX9NFl61F5UztQMCOHCbITgI5qa49nq8
R8sq9IXBye97yev1oA/ObXtRA78NMaDDsVqtW2R1CvBj5LIMXSCxa6yvAIvLvv4Y
SDNLubgkA4d6mVkmB85hMGbQQPa+j8ady+SjrXQdVUtK2pyPL4RiHXMIwWwMT2LW
NhkRX7yqmEtDooQiqlHKvOqzqisaj6K4mGC+1pP7CsQI8RKlCJ5cEf4w3V4Hx/fX
NNUdbhknhQO+x0WTl4elZ7O57L3gR7SMLoG/DQIUKwQ=
`protect END_PROTECTED
