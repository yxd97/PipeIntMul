`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ciZHPgEzoPkR3kZcNOdH/pzSaywHYPFdXOOGS813AHSzQtyQ+P7XoIPRCp8LDX3L
w2boMTDT2VFEDquEx4tN8Vddo/8QVfqcrnCJdScKoqnXQ/OKmh+OgNQHpKTq/2yc
NYOZPWrXg3XDrnBomeiQAiO5tv64p1KZ0VKGp8oeUWLdSqS7eUExARFytjHSM5wa
kpqvjc8Cu2OVJUUpgI397B4samQQvLeplu0rNfB/+Ru72ZdUdJjnfwqqggf4Fr6c
Wm0oWIsOY0WINCM96qaBTZG1Km8w3HJc+JfcuFk/6q3UyxGOiOemim9XkhdMPU5y
M52fjoNdtafhaY92WnqYj6R0iV+Et590H03btIVf7uY2BNZE4BHzjU+Lo/niTjyQ
SWK8MC7YWOPbmYv7IZliz2HGYWgaIVjkmDBQt3sNC4VG9zB/vGn96RRqJd/33fjV
50YmQjeQ9BdXzBeGrx985AFjVC2rYwbPeQVEali0P1he4J1Y0BwjV9xcF8lrR0uy
7GK4R79RiZ1HAyouJKPj4f4NyB/SiqGQi0cBw0OFME/j1Vcer7nu8nxSoWSi+NSR
5v1pieqJ5i/fKExpbuXwBXLt53aQceUCGBMe3H76JLzzeUASXe2oJ7EcfiE0bfLo
sItgwmr52h5h064WYPA+GvDChtnuMjT24c1uk7iXoB0SASYpFH88tIDTV7uNbgdD
G4zOCN9ls1597IniwV1O4DaqiqUrKsqsjUdjU5AJDGQ=
`protect END_PROTECTED
