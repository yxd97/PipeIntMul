`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPznRNQyltG5F+XmZlePNlmoe+U7NyMlkf5TgeaMcPaaQwTmV6HirFouMu52PwvC
8L664e1Rpy6wC3rv0qh8LE/MAbLC5onZQcnKlFKA5xUb1q7gXSKQ0q6FkxEeMFh5
QlRA6bWwjWL+dvs3fQaQvPz28NuMnq52ifjAe18SiqBpISCOPgrUPSV6gwbZMDpj
0pdQfff5patHiaokMLEkGdfMz1+UIyN/uYy02KPCnQyOsB5JoH+bbLumqx2MkLhE
nRqjNwoYGYStS5li+/8LJ1Flu3tMwVPqx1CLFA6V0xfaeV+wtZbr4JFaKbVq3kj2
b8oN9ns+6iy/yaEMgHyZSZNPOsL6hK9ShPHibFj2BM5k+B6Upzh0f/olSDx22eRm
9oVhxj7+hRDKDf2THVs0w26t90z3Lp4FjKXmA3vGlGwh866UmYZ6SxXYK6TVfuxQ
6hrvOHEOUwSwNVyCdkwiPj32hiLcew4LnJSeNb06iaLK7xZ1Tu4Nmn4/1LyfU8GO
c3ZtL53ZouUrPkjjCqTM/umQb2NHzGNA9QB+pcdS7FSU2JwjT6H74XziLEeiqqSx
4dd0GF3l7wcsVBm58lWqW4mV2o65mFAiTqoTE0v4I2b+kx0yDo16O0nzt4ZN2ax+
5nn2hh4gpsVjf/PmLMFfEJqJJNBvVwd8T0QiLYUt95jroYlPLHfPLKzuWw+LGRMQ
i77MwcJf/xKJqr7bDX9H7/oVp1BIQVGiSTU7hJaoojaUXG1f87BchsTpalweGj+6
qL3lAjHO2po917ComWl0GItQgz9N/3fgaHcJtEcsWGWCxiWRhluWWOOPh7OPjGHe
VcUHMH2IjN5XS8cVbOeimI3BG344hFMK7IGFt1kZI0ZXLitFCawzv6Lj0MU+TrVJ
MXahBmCVU+iUs+5ZHALyODY4ViZk7F12huGyVtnbVgE1+OQN1Jkaxhp85hQzqd3p
KXK2KQNcLaNu+dxxBQTdjOEBquGus+VAhQyTmRsFlSxj2/sgb/Bq3g+a8PcGZo9Y
a8YFoTWJyDyt11Cjcb+CuePDvTHUPa+x59eUxZrKNwZ6NAZnKF5ECgoccQ+YU4G6
wLiu3h9RbaVsyGi32BACVRPZAYpx8NoSNtsYJXs44e8bIrVmH1TuAUOPnetUbS0N
+JXVish3/1f6/+hBYEnMrPKyfBlOPSlTl1bXFsqTXmcO+OjoCw1MCY/RZk4H7m0o
JZJ8rwKSOhS4uRgON/KKvSe12A6u9bLxKpilgSKdZa8z0rt2vbtYwQBkqmiJMQob
xfb1YWNkWKBz/qFHZidLxlDMGA/waSB04ppR8sA6QQx8m2EF4P06fEPqxuPSs4x8
skqDCjHtsMwzIQILawqoiot66vLp9lZyMm159ze3/A9fwD+SI+/WxpFx/69B/+wl
h0ysolbgVi5hGnJkl6n9Uj4bm5hXka5gLWYEhN41IeXOHxZGYo/DSRiOFK+lTNCu
`protect END_PROTECTED
