`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vFafNdHZLF4t+OCFm02q+H0cjvT3thXdpWiTIGI7etVjxzFEBvgNkB5dfdy38F4D
bLkkD6mp/3Ql4GSinx6wBovXnMnEdNGui5VJyQJrYU7jqxOgL49qq+OyihqisXR/
s/dztnw3NcixrdXQXP8CPEhLs0MpFLFr/dOBYqIrvUlQJwEl0lPSk6Xfcd0MgmvX
jOPRKauISk3OBD+0c9N52yP26UNZCQUBdjlqwLHdryfDmXlRMPxF8UDJ2VvlRdae
WhvKwWqFE8Nsu0VufJOSEkm5+jBj56yh9b7bf+J+7UcmFj+6vHNqzbafPGMwmRAK
l1OXSCYfEty2Zwb6nkvEi4W666vQPKscNRlj7fyJyqzMBMYkQMduteS54RkRH0Yf
b8I4o6VkQTP6oJ/DYz2wXfZQb0l1CNno5ZKAZAiklJkZsydi+fKts1s0PhsXHVEJ
j2fnC5hpUtPVbnVnngm4MYMsfOUuqP7k9gK/iYBY2VG8wb5Dee/Qiv5RSfPTj6kL
CbJdtLnzoYOLHRCeUKcuHo1AV5gl/XnZXtQcyVUuqBtI8P/0V8z903SINkUAxumz
GeCYRUJ5Yq7JTXAAorO6QVkrT8S9cVb0V4NpIubp7ZALzK0Bpgqpu+EKtVNlbQm4
b5/bhpyQ5TimVSqLQD0SkA==
`protect END_PROTECTED
