`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sPkFKHlGg7DRBC94XzkcBnmpvnI3QUjDMKtbH22JeojJRit+wuYH+zIAUqS4kLpq
Qp1RQLOMdioEHGWC8ZCa95PcOt7g/duggki97aCLNwbncG4gAPAaxRJ68oEHIX+S
midGupi13I0dteePvi5WJJXzTfidQBnP4zKyETNobehKhrL6m2F3J3sssqtrfYSr
p454qcHqPe3WJ/fvgo7+y82dMaWGHmyEU330gj6OTZLP5bj0BCeCK+wZXMKLR67k
Rxkuow+deOSKxtph67NbIX4q0NC5lLNVIH9DJlC9FM3wj+yIzQ2uI2yEqIxIB+ZX
SBE9c3cj0Hhav/EgpoapK8D4ypBozl8hNLkE9h3wg338hZ/Z1NXn81bhiHV1htBj
tPbxt+bSt6qJy1Qlb59oN5PYmxqLhb1l074W8t+Jg4B33lTWd0uZFBtvSkNpLtMK
blQxXBLD8QAzEQCnvv9dQLrNWvziP0RQgynR+x75Ws88/NNKR8IRelybtCgYNHmi
2MJCkWCTI7IsKqwkkMb/Cm0XlHc1SCTHaB6MmRJznLRyd0VA0svXwFArx4eShoPo
FdzZMMObp1D4h2s36FK8Y6tTsBJamKtUn7Xt8W5uauM=
`protect END_PROTECTED
