`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7yi0sTE1ylTVYfl8d/e1pGYePZfjs6Z59rlCwTd32Z4pcw+EG74Td5q9lJEvGj5P
q9fpY9wREy/W6kNIcmSslmy49uqliiG3JXxBK32y3uIG4sKrxKLzwRVhdYvmfJax
FQkCM/hQLJUdZ9/02YOEdF5JZHGaUtlALPjULASyIafy1iIyHlRslHiFsdd7nuad
HV11jBsjeRvK1tk9mQgn/yPID81nQkZNL5CRYZ2AvRMRbtZO+Kup3oJZj+I/Ehf/
AGKiO2yALO57psuRtqUo9jVpOhSORk8JPlooEv1sgjQ=
`protect END_PROTECTED
