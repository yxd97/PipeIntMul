`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvIAl/sVkxbn5qjsK8FG7ZLYm0nH60ULCMICN9dSFjqrbx+zlVd3i+muSJpC9I61
tCICyn2i+I2QvqLmaoKh1E1DJEEoE58dzY7WKnkmObqxF2VyvRZbbao9cA+9cXIC
ut6oU8OybzfeFzl6kkEEOQjCN9hGlql+l7Bi3FwgyMRCfQGixTsBmUgEZOYMsCej
SpWsbPYbhR3Vl2PGbvKWPL+ZLtx3X7QsIPjGxImL91DBC6UU0tSMoIKzsfI4AdkX
Lhx+kDmXvc8n1NlS9CnaKLyoex6+MnWuJD2e0AhlJC/Boq4lB/5+7RACzFi6Yo7i
GtLjcTB0HtHjM7txd9PzftqYSNhmq06B0cK01hickxdk3TMt/SweRwBIVz8v/+g2
H/nLktYuidnUastNJ6dZ1XqUI5HMc0mvdjZWah/8XiWS4Q1cqP0UwekZNXk1zHH2
x0ekYgd+oIKhtWtejxtVHYOz+WKBoWa6GhKZepSw9QQo4u/0UwThBCTkasi3Ha3S
SEq7KcV6DbEBg9qlDeZNp9B/FBNcyywaXNdstOxYsIEraQQY/P5pt7D+VOFpF5Zh
sF3gKTz6LtUkV3o/+MqqzKx8X3S+nXpUv3PMpOhI7Lns/6n1j67VRE4YBHKd8SiV
umbzpLDqipO824zjTuQWU4DVZl7ORumYh49IJf8NohAON7PxxTu9Mcyj/b0AMkF1
kwc8QKmAz5bszpohkBRKdrKFHUb2PKOE8QMbPqIka/pstwmMlcwJ5WOdyC7UjsVZ
VIipwxRdRYIvKjnf4LVERFU29RIXRYwuyCN+4Hg7/O2pkks01ZFqVjEOdYkdwF4S
WDVL1W5fVmAdV4YfmJUilQXl4Q/wz/JfV5sPKQB8SevyO4SbymACjris3yHSLGcH
`protect END_PROTECTED
