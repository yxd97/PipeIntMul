`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
43w5owRvEs8wdCYqu/yy284J4n6vDqHtXNgrcXJMP/ZdpQ8wH5lLKR15QRxFH4nK
Jp3Thg4rElH4+C5tOjfhanoVSb5e9Bp40E3E4uWka8gGB6ekBVAdV+dFFvxysbFT
+aZvGZ+8zm7hWxHOnQkYiXuhv0A2W1qZs1SoYF9EUy8CSgXA3dnC9rKlefpx2vC1
z0jVKvFKklsgxUKJpKC623GMBZUPRxYUQ56hLTj8fvCavjD/CJQoqj4K0r/8TBBx
gAmQdR0oBOBzGkztkqt6UMj3cFrdgUZWb190qKCDokUnA+IBN0ySzmHmlVGOkJ3k
`protect END_PROTECTED
