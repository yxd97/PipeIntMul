`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0Xk+Uq4UtPOyV2k6wjQV1UhF56m+560iprF6NPts4lH7aGZs+/omalqGTbBG/xak
jmYVpYTgC3BjIRWRWvBN623DV8+ywcCzlkMtoT9HnQo90B/lj/W+NxneBqlgQU62
KKsAAa3H0/+ZpByFLwRU46k4GawmMbCuFEFZSJdetWTUL1NU7iadtEBz0ggVHdK+
QJq6Awsn4ctCLfLMKrEwdxM8TusmEgZxZpIbUpNs9kD50nG5W2Z2nIGiNxUOy56z
mfIi90soCTKykOmFWuEdU12KQokc/BZhHTy3J9snEzzhP+bEHB5O/m14MmZgOgjm
8gpdZv4qp+0uBG1ZIS9HnUfpEueJhxW5CQByultzpxXQbdi/Ada30U8lxjUD/W76
Btq09HZxCmzKZ4RWrhPb8Rhmb/Sbxtf3bhYLNeoiE5Dvxtkmv95UMRZIRURSN5v8
/n9G78S0kWmiMuEP56ROmFxn1wjiPVpXZa5r0r6MSZ4miyrfiDh46Xl3qQyDfa8j
eOB+h1s2bM0DXZ+62b7dg4sTTQQDkuI7hH79Fgdv40Wjs1wsh5fn4mCeZ/yaDqWA
uCokLal89uLQfDLYkrX3+GexRri5azpZzscLWB9+j8IzOhwqASfQbXtHOu843j98
HiuxlBrJq34oXB9rIR/YyE8ZQKy7dT8zqT3x6tGgc4nVcWYz4B5fc+kv/ISf1974
50ZKrR3xL/RX2cUmWn2/Qn28nHHA+HbqiFf79rT2Sxl1dC1BIfQiti11wQ70c71a
ymYVLQuKpeHxv7MdPO3mwngQPwmUuvK4Ibr7NKALi3va/Q2ljwa0M1XvkzxFGnCW
PWKT/Y9m6P5YSgXJs2sQv4UHxAo+x4FgKhoJqc47pcdkGfzPlM03qRVHe504fFcM
JbG5Z/bVYJwQ35kbd1L+eqT3Hbj15nAcvmsCa4jdD2rZB7EIXwH/Z2xl6U4xOB28
FMPzgJby2rcwXAuys1aLxutAnqQEfSUVknwtUIUVuRwH6QEGAykm8r6wzKmkzvcY
2aAanEXanz4cME/ZmmhgQHXer8VYNAUqXFoLO5cxqdl9QlatoeGrus9HrsV7YBS9
rwwif9t8o9AjBBV5Kvkhu+pv9zgozu6fdfQjQD8qdxN6g7WXtqc9FHf43/YOK5bt
3FiJV0wy9So8FElXfJdGZfIm7E9HGixb5smSObkF+SoEt6X+LU+oWPm76UHOJ7vS
PpwBKkwwfcKVFX9zD/2KLcdCryXDJscW4L7EVhCnNkiHErXhbOCoNgz6PAjidmn5
4qIUNwMxX7F5wDpgPyXjCYpeWdjxFULrQd36681teoS5O8xcKxKCLglSo2Pkv72d
UHzwaKzDwCyTj2LgLl0/HPVye5auI95vTeuZeRLT/dlMHH+h0Lfa/0cD2LdNnkIj
Mi36x0upQDwMzKwX/TW0b+1MhqXbnBfYrDT2sAuXurTroa1vSyeSOy2Wo2AoRrCc
ZWPsysWIATzicA0GCMBsCxggFhcr3aEhJY9iQctfelxK9tY4mG4f7htni0GosyLn
JY/U29HBN946UN030w+H/2MGACz/QDVaRQEnF3XKYki3dlnEkWEwPhEJUnZUDdtU
VVK3RoNv5t3kSjf233S7ugO1d1yMlXV42oIqbGUvT4+MsWKZOb4OMqh5uQTJB5mf
vpvbf4gvbrllGVDrkSwUv93YX4V8t4OuuJGUy2FxJZkK6YlMGElpIFEm8AkwMZWS
84f8W+heW6vwvD3eCOkVvoocgFv7mA3U7I5cs+k/11aP7nfS2nnekx9uYh7qPbb3
MDFA0kTofAOaC6WS7TNh6RKXOYtDoyO8Ds5evF7zEDPCpaMXMxdjJWKTn7py7N8c
5Vw3t6uTs2wW+FEny4oz7vemdZD2wI88Fwnx6hvgXPdJqC6T8xXQLPmYyjzQOIlu
6J5MMCsEP3S7To0fWM/LzdWXxCNA5glNHoUUptsnGuuiVUb+87Itds+9rbdNd1HA
lnDYLzcX/mSDR3SlEDF262q3SdnkRfABpgO5ODThLLX0SMgD7QayLySVBh0dkkiE
WVki2aNvqKiCwV2A+FkOQQ==
`protect END_PROTECTED
