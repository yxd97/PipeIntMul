`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OsMhrL1iyH6+iTwVocp2TXFDxO+QcP5FGDaIbBEk0nEDycoCCoKWIKUjQjZGZyAJ
ZBK6xvvL7k/HuQLbvxfir4wSE657RhdqKQcmE3B0NXjgy09NE2RNeSv/3tqcS2jQ
QwcgGzWjbqOvC1/xU0xCEiuBbF7gNskoGaDb9thIeisaBIOdSWM+45jhFBY5vrIr
u0TS99qhZ25j9woBoSVyQOVJxsS+VlmdphNN8kebY1Muii1kJl0LSrKlr0bMxgK7
vNtnW2OrGYaxMC9cozjs0HSAp4s3Lw+Sth1y0lax351mElacEYZm6BcWxBWfC/Dz
eAa6er0G50x5HjvCW5hf31i2wQmDu+/jQYwho4jQCB0qQIOm0LzvNmm45bJxDKIL
`protect END_PROTECTED
