`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kZLorAZshfpuvkHCAP5qp/jCf+XSq9WeOGRZLPLriRLYePos6hkXWVQ3gaWfyLRW
xvNwcvqqE/fXce3IwX/lWuxJ3txkj7kHdtEJcll2nKtECKC8mjwjLwm4y2RUCdtG
hxO+HupngBDMOnan8yuclTvFkcagKFTaN7GJJmA8FdijKsip+AOrCwobaOKkrH5L
Qj265eD+VqrWid3e6oRCJOG4k9s+mocjzemS9g2syq+IPjC71MT6k9stte1SGIrG
i4l2HMqqPPJg6XFuV9HOtg==
`protect END_PROTECTED
