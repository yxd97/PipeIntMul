`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7lqOd7gOGIG1wMIrYXTj0BLVxMvg1W5frrmb+U/nBM1qegEgPwm0M8Y7+KTwooDi
e8bnA5NSpx4fuzHiVbor49qQdso1dGBzbPr7MibwWZOTixgc7r7KuxR2Lj/W4GXP
lHlbGFTXuv7QuneXh+AD5z3cvQzLIWSgkSBsgn5SewIwTPWmE2JmhyITTLBuPQwL
0RSH1EHUbjdtG3qVFHfU+0szNKEEehYJWjjsfr2J+sE04c/leXkoYSnSQwF8NHMQ
U88hUU5LRBZY7HRiLSKSC/QcdQ+5N73YWPiEDHon/MntfwBk4pF5XcfXhA0o4xbs
kImk1QeIOZPbpmyRWxggUOlJqBxM9bWoQo1O9pqCOq8f8hkaBTtagxgnRrI4KHR2
wTexXCn75K7HoYBDAb4hf31f6gf5buDnsSwePkAPtbef5vm/FyN69Kbg3Cgt87tr
B+tExqOYuo9DnqjD7leUGmRpsB3jQLuTCHu+JEPL0Waxw0n9nHLTePjrh6QP6OB5
Wd0WagJ0Ce0Zqgd2F9+oR1xiMW9Ud3o1po0H1rksjW+79VAhpDkbA/bq7Q/QxnEo
033jN6Jh5RjKUbhMJ3XoB3xr1z/hsoVOYx5IiKkAi79VIoM3sVMA32t8xopsNmfk
D+NlfUUcE3HfhxUff9Lk1Q==
`protect END_PROTECTED
