`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCqtPoJcxFraOBKrdaPrk5Af4nL4QoAwTBLXMcOYhfrhOJLrrBUbGaiYQhxdp1uo
74ER3j0gUC/LUfao3qYFdkBapxo4zcliZy8dDh4Og45Ko6iyLds0XNCuYgS9pJez
P8l9ggUNVOKR7S0lJvR15TVwUlPO4oX4yjkxcDJvLC9zxaWWyeLypMjssZej/zWu
WH66DkCIbL7pvN+bCckTzaZbzhvniO/NB8O5IDisVI32kvOQXJjc2dPPtO8Dd+/D
4Ry1vKdxIEVjaYlNWVCMdVPhzOej8v5aK7xx+sDicEePfe/Hn0+rndsiJP8DWi/V
9HADot2yMDN3kjI/rfybNRM1SjSY8RBAWk3vSJaeI2DtKocQB0cnXvI11exaHDXA
`protect END_PROTECTED
