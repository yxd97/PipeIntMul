`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JvGWz2u074NsXGy0jED+qRgKpRk5UNO1CZVGMJNYUsYZ8KBp6TVRo4WRy9Jvc5Zv
OHBpMHciX9jAsluMQ77OdLhbLklSB+FSMUNtldk6RwHLy5rlRqbw51HuuHJuno7l
yvswNglBzhvcDkotwoQxFlw331dYG3fECo4Lh1L4F30ktm00E7HiHN/R/Cx6uJbN
bfaQ1897fwMS2g2NgXrU1/CEQNHu+sPWsE69Pl0x8arak9jY8V9kw7v9izLbK3N7
BbbVNkqAOHamnH7ILaIDKg==
`protect END_PROTECTED
