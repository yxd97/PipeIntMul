`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BbmH/nnhHWffbdjoxUFsC88Pezb14n/b5eNhwBN3NRPoY/ksEVgO2h5Nm5GOnv7F
cRZa4FldHR1KGUXvI80d2TCFujvcHPfKUiw2FsCsURMRS4kiiNNmMXIQvByoGMxk
7SUwUPp6bKRosTNpFQLjniHAm013veO5bx3BcvzL/KpIohotQCZG+ClZvkG1WJ+3
CS5hsLSC4NxTUpBpFknVEcxAe5avLfAGMEWlaVxp2/sFWDtZYxUQa6EopfFtwNHp
kBEYW3biQXGZ4yKr9OBX1g==
`protect END_PROTECTED
