`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8SX8dFte+rWF/xEIfdOZeo11SDjFSOdsqsUyzQbHcn3bS1YQvfB/8u0hR5VgP0MF
3unKlcFQ325lZClddigTkVX7x9d82av3JXt83HQFcvQE32vsQ2OfxjeuCMR4EQb4
ogEKILqu4feXPno8wi21c8a7n4F9z5Ul89D61yZOLOAQNuSwgMJig/fuLzOes1u7
Mb/3C4z8xHLPTxpCbe+/afBH31isTnqZrLUzSRqi9mpx92vhyDpTVJwBOUb/CM1J
UukSLY8wKJuDZ43NvGng21RR28JHnk4AeVLAkJVjju8JyIPxBN3BkQwJNZVw7W8h
1+etfQpXAZEcveQpad95H6oGR3WvEfbUV7MykNO2RJ9qjzIqBDNnIQD9WAIIxTky
HcP65Z0TnsCIl33pRPzoaQ==
`protect END_PROTECTED
