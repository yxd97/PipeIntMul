`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
280P5Fghf8OQ6/dMYlMsyfuZdOMZqklpcSpoA/W3OrTMo0iaiXlIf93P+Xv3Jaaa
FGDxj3njj+0f0Ba5ggiEeo8HkYcoRLsklhDz16LM94KzpgTA+8kZaTA311H/FebP
GBwUTcRP77hrAtfEtWwEkoD7mx1LYSfGTajdkFJdzZgESnZwcubwWDz2dc63UhH1
YmeiWgS2aH79G6hacBxJmWjG+iOzlyWvUWaaLEdacva3PYw4xPyiqMZHg5eGZBVS
+cCZeUSNQuKibyxWZyv1P9r75uil0ewjl2EPmtY2+q8=
`protect END_PROTECTED
