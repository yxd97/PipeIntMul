`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YiaS3IE7uAYdVbOU6HYLAxKD/7m3ZLW3xYKpkoLhHqXnz/FwCO69x8pDj9F0lUxz
h1V4AXZqZF36J0gGqbXkaVFAdivktSyTF78ThQ8V7mqS3N6Lt49QGFsQJeqzifiI
rxnI90Iotc978ZAnYQFxYGgukL0vINKlSK6ziAu1E+chXrj5m5k9gZnH45CRvZ7h
uu6g1UzUJ9MDrKtuBUaMdyekuJubvUuU8a7gzGp+mYGJsFJGl9AB88Urc1EEIWix
kyxINZjd5KE/KGDXRaBwjsg+J9FvDAVGdDosSklF8CyzIJu9KI+OquA/xD613wGf
cmMEZ6K6EYmneUnxbVCCp6726EcHxZ+u7WZ4kqHTAxsNF/recb5Vl2J115LXRnfg
q5tDGtUf/Uw8CYp2fvUFop3R8/fQMi2C93ZtE4XnCLTg4WiO8KTsxanSSA3ogg3D
BH8oP2dM7egzeHk8O53Duohhh9Uv/OKmrrO+NfrmuR9kzWwHwuRRsaKumUa9fJ59
ToFrjXqSbRW4ew+D1WEpiDMduUffokMA0bLKl5QP/Aib1ttqyv2MMPrySD+I8eLc
O0ZOtbDmQwqkLDsriOL2vOQAgmge7BxOOri88L/MqmlkWxwT3JPZ0dGL33gt/ik0
pquRmERUlZqlQQ5jlp/jR/A8rrYBOHd5vuwM7LcK1W6J4Y0YGvaXUR+Y+utyeNkj
qMM/ygZCAsTWdhYPWzJPtsE9FLwAvQTe+OPIUYfPAlEFTmJO2RGknvomd7BZtEjh
HlF3x8/EyfqAp9bltqE06dVo/zi1oIDPboVovEYa3x3y0BOuI66uY2N3qttJP7P1
wtnaGwiJHJt119obe5lYHO/mvfLOo2NA2jwgNhxtBDolrZOGHZsVLe70ZitFgwd0
2qn6mqytPl0qDWfakkwWlQ==
`protect END_PROTECTED
