`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1NWG0yn+VvCjIPjui6vZsRDlYpsBVcFQtW4sDTNq3EbDtF3RtOSwmvyDU/EfuO3H
DgzewJgvZmgwIXTJ7dax2Tb81hIM/QuYBDiaiNrl5h6WEQttRThS7/IauIKQgRVN
Rdy9vkfXGux2xtA6lND0+MzreloMil5Y/F5wpjZ2ovnuaaX5IEQ2s+p/i34Yx6PC
wciItR0shAk0492ALosx03p3iITGhwPqsxVeMubbutw3t1d5PtrOPtR5ylxj4PII
6279LDO89lfrDewmzNs57a3r3xS7+AG2kOh/PW9pApFf4OE4pIHNe/E7uqWGLBSd
dprqXD4tdlpftBbYtNVBkIgiOzTsrRSEMdY5jvKwg90JI1drjJr/hDYC1N7qib16
eKys2modSv4GmKg3F1rThpA9XpjCq6tGM3jpcTxMLWavaS/4okKBPEjHUodg6X/o
lES8oYkbwYXKN+ueMfFWFaDNLdGxdDc7RUMV51+tM7qE2Gho4X/Dx+aQzPRP1+IK
8NwTEtpnzWAQ75f3lH0fOMethCAef6SmpXPzdj7RP8ruFggT1pDC4h/3idKpUxMJ
ngWRtpaPfQC86TZFjRtHwBvcLbEFBlpTs56qhRstP21qFA6Cl2DxiENWER+A9rrr
1W4MhJzVaUkomq/Fu5rbc0kvlJEZBuO3Zb1Lq/sTXe7Ci0FX1eU3kS869+C2dF+p
`protect END_PROTECTED
