`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iDDCev7APizJ/Y++a8PIpG+dYZT3riM6ssN9GPYTWxAEcNbjFawUmuc19XjTJCzU
vXzu38l6TD1kTxKa8ruLV2BCXiiYdx/2XFuHBhHxybFlg3fxUX/bCqzNKtqUPnCo
xhpEOkeTvzX4o/P5/GoIeqZplhw5vusxDadY4nLPIWh2yt3RSm127Q1rp6ux+oHy
wsBYZtCqhXsH+PbOEcX9YOJI+Bxfay4+0sZfbTui06nzVpJWb453ghHHwtZYu+5+
thqEQsXy1ir1wRmcnP0Aa23Kt7wHHTAtciFV6GmQpfYEA7A+sJCofbV1eqf8uO4A
O4wpvnyq/5QVHSuuWUuqWubwhO5w7Es3obtA+/LSb56OP2QFTt5e8LoTxGtgjKeW
QpeI8VK+yYpt6tT7n3QkeNNKsjDmPPmXm49UKL6UMRaSiJdVccO1r/NvMXmmvZke
QSu9OGtfL/Z3UJEY07WfzWKq7Y5/EeXjC+YMRE3ABPg=
`protect END_PROTECTED
