`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L5mSyuh691PMuVcwULpSTqidzP1XNlmQg9FsWO548CUBmeppBcf8PC7ZOCX1HGbU
UOWKS3mYVYIwKoD5f0OsWZl/NRyAc6omhHrCiHASxiYZSLyH4uOO0nVIdNsDOD/m
pDazfflUx1eivWrM9zqPwIJ1PXkEAtfUbtm/lom4QE2iGXcyP7fgEafj+05eN21k
AWfwr7O8UN/CXDMh6TRMods6LUvdlCqVkuIEBCTRpwXs0dceMS5buaKRIuGP34+v
zY27mN/2jFnqA04R6vKw01akjXBlhQwDIaeF2LlThSgY0IjoPQKXVfUv5jqU4Gyx
9TkrwnMIgIfj8WqrkkIuCczz3kl/nuEvFdYoCsiZ5MxWDS4P0rG6chK9RRjfkfph
r6GXqbERGEHhNkn+vGeLSiItLHZdZfpND03Roco9cXQla+bI+FA80GCVFoGWPQ5V
AovymfzJj3VYBvkX1zM9hLUxouGWtRJOYTuY8gaQPF2/3PeFTaCzHhbHB8Jp0193
FLq/pU659pG2tVEJUbAet8TJRtyt2ElzlBI9qLI//X4iY2K1qqVvGUr5nVejHz/O
RRIHm72cJo0v/sXu3puij89nQkajrsKGla9F/Iw/skL2LmD4YLNqd9OtVTK5AFyN
JH/6OzoI1wyNOubR2cwEAo/e0cz/N/5kCw/ZhaJWmsMtQb1u/afOFBhFZ/tA42LQ
kb0xi9PKR1v82gStcY711OfZTyWe3wyZejzhVNQZFZTWB4+OKPvpGe0maomOz3Fy
v6RQTL3MXpFzlkVU1AuDd/UIPGmPEDu/hlGeYnRtQqxFQXYZsdwKYaKzH3uCs5Mw
qlD7BWSOPIioWEKtdeDHY0hNNJYyGqPW7wsq5V+1mCh5xQP4jHDE26xcaxeeO6+Q
a7UlqF0v/wsUXDgDiMfYnJ0PdcccGVHICsIK9FEdVbrpwg0wNOv/S6rcqblD3byS
7Gsa5TgDohIx9RoGl/roseY7Y+QUDkYgbazmIi3EBoNIaMVkOYNw6e8ggUjb9+hi
5F92lf2VBrViX7jgVySGvFpnTSGCF8tiAmyTWYFqINyFQBzD4WYf+ARhvx5BRt3B
JBPhcocMEcSY33KA15sVA28VOY//+wLECTcoaYNWyE301lcfa6L7YiY2ntQjkDgf
`protect END_PROTECTED
