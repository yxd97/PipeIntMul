`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4y2axvtDjzGS1PDEq2raQmbnEZRYZezN1Bx7PvOa/y2S9/jsL41uYMhId8UGMCG
AHA7d6f28l0RH0c5CqZAXQ6ONNcWdyiMxpA4sQk/uBOIoh4OHmwaw3aMSh/vHkwb
WwHPh2kAAV3rsfvxOws6YMVZiH93pGXQVLA8QCB1ZKnc1D4lGaEakuDe6mLLvy8J
GdDEfw68Ma6c+NMyf/qapfxZcAAXQ1SKC6A+qxmialpCDa9RwM+PYdfbbdAsRd0K
j1ftMW/ntR7nWoybMZnkrO+t+44QoBh54Jf6jiH9Rv/zQm0Q1yZEFnVFAsTW3x5b
odUTMAJs9uulZjqCjYfpDe4AbXUkYu5MmukWOCUYfMy13MKgS0KnDVhpxA4n8Y61
Bv+U1fIHgCyKzgDZBMHg2tZ4q3tEmX+5ciV97VNbxqKst7NrQSVaBFqpSpmUV60s
bPOYAfv6TZJmOPRj2ma+Sd61cLwFWbTISCXUNtOO0LP3Em7nWlUFRX0y4ROB5Xn+
DWsNFo7gJvR6BTdRN2ITb+PlbPdxeitrcQ/qWh34YbuikPjCFwcJLh5/XHY/q+/G
pky8rJ2gzcjEUAs90kZ6zbGCgyaMgRvR+62oOC6qE7WVfblWawuvzR9AA8WrB4N6
JnEfB+EFYX7Yvui4FfRZuNbQ7ZdZYRZPTjj+jznah/vd0hf2lkoyzvdxchXCS1vA
`protect END_PROTECTED
