`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4BauWG3Q16WeSxViMkKAhaTDdXojyUtkzmO49Cs89J8eD8pGjavBolHZyWc2s18D
aZWeOrMc+2UqHs2KQDJk1gV3/qrzYfDHELAQQVmJrFv7lUxa1dCwaJoVH8R5opDx
vLIzeEXDc3Y4d7azrAZprEaMYpueYgiDd7M0GuENQUGAEZ9+SODtX+aoqhQ+x84S
siQfAFlf267nArsjSiF/r3FFC4jSqq6ey9n6N0ysuzevtXX2QP9U0W3bUd3BYd0b
BDJ78JGcCwS4ikRj7z2Z3dLyRtGhFCzve+v4hxrWfI2RFH6J+k1ZQ80Bh1/6PUiM
LjtgD3XK1nPQxTO1/2KcoRtbKuF6ti8EYCNtRvBt0yCjzaaoQzTRPKeeNW0chCl9
9n+F0UgGpiugTlnORqZiK6G1UQWlLD0GLUmOVMbNhig1cM1kiTkf9XVgjtX/rzdg
M2Jfe5fx+3JSsQwzykAB6IC9Ke+FCg15hwyuq3gUGYY=
`protect END_PROTECTED
