`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+e2E12wLTY42cNRt2egf0+wPaSIt12HOd5+fO4VuE1ZNYkOg244IWdH2RiUYrmQz
qClT75N0jnLcXb+di1oPZN38YsnAW62+lITahQbpChqZnJmHgpBjpcDTmOGmHfYW
sIn2fHuGl+0E4+MS2pLdDhn2WBjSGvPzcQHov0qIHkz8vAdFLi9DGZYyHKZXjC3O
FCFvt/Q9U53MMYgyG2N4Qp4c4uFU6hbx4ZfgNfifwAmEHsPE+2q2DJcLLYvh9nvg
dvMjtQ2EF+dP3YFnhoiBuT220Ldl5BlrswIkRI4ZVDk7Noee4oyCR3lCgYLoz64s
On8NS/RYzCQNy5fzuRyVEg==
`protect END_PROTECTED
