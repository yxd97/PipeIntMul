`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SiVkV3pVLWCbOwwcZiXDTfL+LsuN3lc/ViV0VRJNr3OeKeo1GK5K1TxSr1oomU3x
UGcABfIbkoyJHZXcjrpN1+yCz4iOr5X3h01uHPl4Vo350wxGcOUmX7w9lokfARVC
Z2nJy++sBToc44ZtOw74QtbgWmR5kFLJkW5ieDHO+WfWKu95YbyjhFU6gOluCD+c
zlt83O4NrXE0AdyM8hFgacJpl3sO51+wp6eHss1FJmpv9YSjILKVLKi2Qy3JOB/k
lWjHTjZuqRQ4Y1/qBxPCQtFZ/bNS5Xf5q4pTlIyMlOpMbVusQhHBeWDk88wwmFUl
LTSuv0327y8lGDn+Kovco+2pdVHI6n2H04/9MPVse8Ur7PtiaNpAHZUGdDjmxGGu
9THMK1GnRedYy7VlZf0Zl6FuWwm4aOErCfAhR7bew3eQqT+sAM1C5GxqAmwNCsWP
oM0EXrGkGjSO/Vl+e3ZmcjErL4UObUEkuzFY9lW0Rdv0GQp9MPGp0aRy5Ge2Ex1n
LKHw2GIS1PljGK10LMe+TnBRKggAbbf2EZJTq4WnAvK7JnjMlalaWGe23ips5Laj
KzmzlymwqrJyTMTzAAcH3Y0exZr3d44bCmAlMkmaGSH+LTC9aQQQYkYuNbBFLsLL
Hzl3yrBgu+HpWWPkLjlKQbNaqcxcC3W65sbuw9o1AkalVgET2wp0LH/TB7eey3Sq
5UyFcKDgYOw13CjUflMUwZ3tSXCIXE5QboaCw8ePHAzydaP+hj667IQS492f4Asl
+j9otCAHweBcR1BqKax8NHQS3kcx6P/Jqig/CxJgZJKZiFx7PK+bsiGwIxI2XRd9
vLjNhUpV6KEaV1Swtwisvp1I4j6texhNMnKRIPMij+tozAUUTzWw5+4GGGV2x0w8
XbzuHcCW3a+VpZUZAW6nMH06FUVJzMzpBh1J5y9409qjSIj5LbY95YeQn9spGqj7
w8PQwtth4/PVPjuk4V43cqzi89LRkI9NlTCKmY8TLWy8g5ZMn5/f97ZfHREIVjAr
Iwl3rz1ah1CtnVMWo78/uTq9EhHz1yx7zwwXCKkO9BlfWMWee3PP1hwzqzaOVFyy
lPwBiJ0j4+aNtuVqYb/+oI4BQfL73/vnW5Vbf6m8I/RtRsv0G6w2e49UzyKiXv+H
yC7S+4uoPmrGFRYvF202YWtUDL4Ic3/os+AegC86wbeZNGrMryaHviiMXnuXFuHu
dhR6t64Gy6WzpMaRypvuOFLQ0WqdApJf8fA1BBzXtaeslAGZx4T4czNpw2vWinuO
kme316Pf/8OSidPv6mx4XhFlRJNN291Zv4ofl+nggHJ+oMzOJGJQN09KGQrPSI95
+jaD+BtDLb6tasmfame6QIjEdkf6vcW0gxcY+t1QgCh2vx4I60AOHOJVl3GDx9Ax
k2QhgYkFDuztXujDlVq23grRg4vusneALLcIP57/oLzTsbHY3uE9PecBOkoWivXI
SGIXBFTERVwHVt8oPB6DYiAxgGu4BtPQN619UH/xwe2EFq4uRmJxqOlZ0fOe/+pl
OGTWkfqb4nYsIJZjQ90QkBwUx2sc7OOd1eAsC3jGpGyRD/ppkLLN07b2+Tn2Oak6
IjkxM4Fqrns9/zJyz0Pb0dp2tcUY6Oo9Dhx3NPhvRIGikcTl6MVwmMn1fTAFpZG/
g11irFTRvD9c8PclY/v0tzCMteI3UK/yEUtEbfrbZsU8B5v0gNLMEY697bL01Hej
vkZDrlP8EDJ/kBoaB7dp/lows2B0c9YxyhgxDH8M9yPb2SFYsozKucwm5WWmr8Bv
lX/kYGzZQwTpZOg51i/k8LypA7Y26qYRyYtqgjy/OH7yOP909Q4Y1m342B4HMsrJ
3n/TNhhNiPFzdmb29dtGVYfJoLn7NGBPV/uXNg0u6mgzytVkyd8otKbA8c/hklhr
x22SOD78luFEjF9S6YjRQbWsFgulziZKNNuXJ6tmxTXxXsl/IBXR57ZWnfN0HSs8
pqGAEhYnDZaEBX8+ya5WB9dMuygCwWeFGiIXjKup0+J/0YGlnCjWhLqBZjdV1Q05
TH85pC4TzKBZrjoVWR8p5hk04FrIzbgKHaunonCWffkg8UVhemNtRQh/FsAIx31Z
W/PE7bzF4ZtrlEtkRa1Y55X8Rdb8NM7YJ8MAXAZ4ZYSCBhsOfJgNLJToGpAKDNDj
Ge9XOSxYc7U395XJ6N1LFdrMEjiijIyhgB4Ao0hvxNwCTOvATDDWTWCD78g8YxUk
bZRQmHy98bQpU3ZCQRG37G2AEV/E3UvsIREpdYqpCamNmyc0W+c9oM/HbrQBCUqc
GRpR38DVF7MPqvD0pEa34FNOzY2er3ksZeip0t5/MvRZHGNZcefWuR0x4m7yiL7O
AinqeRBg7/vNdZPfaXMygNOjTCzyu1vsq37FCKWo9PhY+4fdtToq8aRfChCNurJj
XL72KFuDq82BrbXykD5CvXfTbpJKsvuiupyNGrRVUlM5gvaTgpGAQHq9+k5WnOGb
xnRjDpBPmhQxhhIhJSJyBk0LyHA9YR2HsE4bjiwjc5ZR8CZ5ME1bIk3Se83bChyc
UyLdPaT5wk7dwo6Lopk1Uleo4m222ZlUHYuDHozA99+BKhS5muu3RouIIv9GBTYh
CUK0L+Fn7NPrP/ISwDab91QpI3UVHi2pBeKN59+XoZpIRjkGjVOu9XATdwqO1S98
fGBo2rrDANUT9WGqhyx/FfIKzyM6PZ+QYPz28EtJ4upOhOaTniOdVO48vVRU3aw6
Ql2eyYXt//95Pdua9QQZ29w9kI21yHF5OuulGAx0Ji5RiMYf57dUyp/hf4FYWeQs
bL88KwXp8xCnyfJ26n/FRErLxCrAhUehB8QoEr/z4kxGb9jeDZlO8LONEXy3l+Au
t+2s64G2gOrotvtrBm6CwPfbEimXqynU1i9tMzdEBGA/RlfXq8/DPH9vRsmbK/6l
7zKwmubHFFzSPCtsXhwmXzl6sjju+Z0uOkdSd8hJ4yOTzml38WYEUloZdvAt3YrX
AMka3lVwgmIboKCVELwPzv1SX177Ks/rXNjguKvVka1Gsb9xZc6q4siMvdXigNr3
zdBCJmFgY772tZJ2MmtEZDl7VKn85VQgq2noXTn1IfX0xDWLlyNcXNBffYw6D/Jp
g+tGOOcO7EdiOcWUJj2e2I7vbrDBdgv74d4Bzp5zPSZJPOp5U4yNgdNumOCbn50q
CS709qBpM1ljVJThsVOP09bNUGrpItIGL60+NsXQFKBQfQsw+yL6d08MZ0G2otTw
5fID62ScZdjw1C0FLtfw1GzR66yi2vs5mh+G/GBWNHQr9bLObyG9NQbhbkRpAKSt
c2FL7e6wYwkA8XfoL9dUjazcbGQ96+46HVZOmADfnyKknLN/p2EvP5GoxoRxebWm
XerQDe1SD9xDroTHmaEmMhaMI9BS+VZzxE5Hpys7mruwl9JbKTdC42/++ZYksa1+
9TAUOrCfC6FDM7WhTkRQelNOewbYEzWQY7gx4NkZR1VdI1TVKcOC2Xe0hHOcyxA+
zB5j2BsvsU6tyHHf/WiZ78ypwwwt73ZFLZeCjYYTPUfnpcWSb4NL7UAgUb9xpwkT
+OvydlsF/k9/tWRUiegG1ak58qvaREnG4ycIk/Hw3+QsOkCx8x7moencEKSCue5Q
7BCaT4RnVgvS7oEA18pQsAndylkShe3on9NVuW52aML2UwvIxGLg9hF4OHgiVScK
/9kX40JS3FymYKdkHuLvgxuNxxvMDxjnvUGoixmofLwNepz0BSaHZ9GgKsGjXIzt
DkD8sWUm+9qrDEaRekEaH0/Y3MMDdhl6Q3yCIIcjjI/SAQpZNYoZ7/vpgmTW0JSD
kZ7JrdICRxGAQO1jyRSVcqfSI2xNLTfecQnMTm4lmYpSU8ki8v9Y94g8WHIlmGey
p4b2zvw5+5VzIMGkd5wSnE03qZx78ZJGexedEg4skUx6bZDvPDTQr/z0bEZn4nT6
C7q1acZyPOAfBtoLr2sy+bA2XLm9fO5cZK2tiW3/AE/eGtYH/6LeZ6qYNH0bbudn
NFBkssCZmUvnx2+/SqRElsez7foGkID509xZGYRpA5pdIAUBOdJhcHANUlmzLZ91
JhkP3hqRjNCJmwVitlpOubrhs5IeCdD54Z/cbp5sLtbrDHczw+9XcW955JEgXdwO
F9SgzgWY1uCRzYS4qltqVHeubgcfGxL6GflLfkd3aRKx9u+bOzgUwLtwaPyYTKco
3pu22lwyG5WkkYe+cCn0gF44K4xCvudnYrFzktjQvmT9rRZ8CSwErkZTD9FvzUpk
MziV2o76q0qJaqKw0CZDSTXyIK+U9c50lu771Tzkld+aQcXIBV2/z/P73XZpy4iL
6KtivvD6szEXUX3vmEhBAMI3/hw7iSasc45ls9FjWe3dvtrY7nEYQZegkfpCc/8e
Z8HM9MjpGWcgpHKYAfzXTQKhHWzM2+tJe7fC2PN97InzuCIg8tVCNW7MaBH1WVuu
ulsS35WT9QArs/zh/LTfmPbCrzNf7J5u1GDEP+yeprT67bJRkexg9XA/g9X+xl7O
D5BKy79sT2NX8f8h5sWRzUjH+HJ13G2Oce/A4qgfNU8=
`protect END_PROTECTED
