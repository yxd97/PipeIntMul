`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u9n+2jt1Bec39PxP2RmetJSazOoE2z+GGp1MCk7VgK0X7Vt+BiVV6v3S16kGzpM1
lJpZ6Fz+IAJPe/smEdJRWpmoEsvEqZJa7xY1MIwAT9DT0GOOB2ll6/CtS5r8+/du
T0eMbwiEyT6FivUy5MCxmyD3qaelRGoQxkcWvyUSv2UL/Q+tydyAdPAHffg/sLiE
0tu2UvC5YSP79Vn53gOkh9S5vTyRGGXTfBqZVMeuoa/MW2rOGBCf1T62xFc/4TBo
cP+PLRKO7Eg5I1k2DDW+bA63t+v2Dke6Hh9f1C4VyOfBPXwafYIW6hIY+4WQ/gYV
WSdEHMQlbohAMUsUP0Wz4EGl4uXs9nT9Wr0HzLwJaxSgUMCN3hL0mBT94CKX/q5s
IVd/hHA9HImtDrdAuw0HMthBFBfJKSSF9pPTod4TLROofPkTPhsJ3r98nkrhDRUo
33xoIGCNvRuRqU+c2cgnA+ZFOhwXAF85+zL+Fwo2LUeayB0QWbUylhokpxlY8dXg
cKboqggHSG0xpY5Ogjay+dkzQhUK+wXmJYjExFqvdRZtEbbR+a3VdHDmJBL0Qvwr
EnTM1Y0xU5TtPihWr4c3j4EFc0H2q+0Ix2RWYHAxGV9TC0ggLsrwphQX0FSH3u3w
Nb2SzSLoaHOlM5k4mCQWLLl2axMKi7bYODODe6X70ykXBX6JhKvAyLUI9OoKeXxb
kHvefozThjEPQdIn/joDYU7LsvXeAop9UjnO31yv0kgeQDXlkQVAGYAGQXvc7iHC
Rd+/rFPyZs4x/VEcjg7U8gJLNRdpwXPYfRwwx5zP6vPoY7G0BvzFAuB2Mu0MJ7Z/
`protect END_PROTECTED
