`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NWuPI7PhB1gaOZzf08A502OSLGeAxeAhRP2GdSF1PcIxFeCm5hxE5ocBeDA7Y60l
VOoONgHaMG78yQgNWjzMTFSIKk18ipyUbsHFTtI5RZz6eItkfwJlnY2Dx+zqNrZp
GwDiNBlyOjJPolIhSYYLtetErXczcBI5e977EPw3IKDsTJjKchGK9/0KP+hOoxDT
7J22Jrxd55QCeUdfzeuAkV8aEO2UhAswRoLUcqo60HDfMUhf3Ofrd2oopgscgJKy
7LOjcENtrEOq2Mx5ihLYLC29OGAnVkrnT/oLPePquzqUaWvxqwVfTHP9iA0qQKUG
SyobK6RbtgL1aZqc9eM9ZEG12QvTGnkL6GlFAbl2TGWHf6Ks7+YaRKKEfacC+bwh
iHKxXPE0RH7OT/2bwf2TLg==
`protect END_PROTECTED
