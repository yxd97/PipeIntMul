`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hbTH9W74jpA3uOqiwvHLmcOwesenWKMnNTAdCd4Z5qcUnwl6SNhSga8xsCPS1sOr
TfPeJq96/5ytpiXjpeNywvnr0e8V1Gs9av3x91570Yw1hVv3aOZnyeryQXbEu+Nz
EA1yGR4XqHTwJ5UI292H3dyQTjgyCy0m1GXvLyHhBNI21R+7mp1ZnhnZghYZuDp4
E3kvHw7atZ2hlq4Jq3aic28Nf8qY4sWP2VNhTivnFNufi63xl7ffWLDHLg94Psov
lT58hQmDhRbjeT+6rkgItTqmRkRyeAjhOeE2RchBX+dU/Ya1LljdPZ3STLDX3R8a
L5S3LOcmgwpOayfhyt8jf/jEE0/wSc40Fxq1EmywoYqHzyfBKTKmwyt0JxB5cuwL
TsBLFr9o/H9NdAU7c8gNzODviefFf8NB/qbaTcdbSXdCIBrvYoQjnm4najgRjlnQ
Hhi2GppE43QMLLslHoe88hNRnfjQVFlQOqeMrBCt4ooJ2/3UnqUW0G/yqeqSxpSh
dLNmLcuX+TVZY7o7SaSG8XW/ajzWciFG4sWS/XhH+oJRS8G3GxWNr+a8raAjqej2
cC4XMOKj5hkbdpNB1P1A/GfjwuN5B/5cNBeOeniXiESX+//akefr/PFF1eSn9OSS
bB5kieEPSSdY4dO3MqcbZBHrrsYPGyD6/aZKdtzp0/Zl1PKIafxaukJhhMWP6KUE
OVxhxCY6lFB5ssgviANEJyidwsZAdcRhPlgItNtA5Jb6pt/MlqwTzjIfM7oEUOJ+
7qJL5DMdEinZpMqLoNESPOsBMgCO4XleVuyytp+Tq+iUvlqViSscgJhVkuM+bsfj
XcnjSGGoksxHnY1WW8wh7Ei3JYDe0+ndSkq7ZixeDdnD4lYh6FUmzDLhLTP/IGXl
LeZXDEUe9DZueQRlPsGjTNSlx1RP/GVr9nQaedSeA8TBwbibe8w2pbjrJioo9chu
`protect END_PROTECTED
