`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RL32y9GYMLKsB0nt8z/GP50qzgt87CEyGgZvxRA8BPyqhb2NfwzTh7v3SLEtEBxx
4qm4wlm18Toy7UHpVl78rkJptn/a+c2rFSPhnYlgjqkmcjg83Le7npx5aT4nwi+I
bW6tES7xkYBGGsxAFQIuNjJCRIWre9npUd9LYvTHrfRwQnemQ9QgUIosRvTbqB+S
FKFMC62VYlwyqxYaUrSw/u8yYv6jTORwxovmX6kQbu6OgpF4FaPKyZ3zjoHpqpGp
CI2Njr68tvs7uPJW9rPq6A==
`protect END_PROTECTED
