`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fapGEvngroF4Zni7INkn3Y53tkCKRW8uLu39QPWa2H4FdUPAGfkcVcACxSrD5Lf
mF0PixTKtr50zD0sPAnl9Xlf+W5lMk/BdvXe2UmpGvR6RZOhWgLzCRbvzlqJq0hH
G73Gc5k6Z8k2IBca2U+9IDXZfcnucQSkGZeS8FXE6JDekC+zGW1yJC4mPgkhuXuo
7mYuoZX8/tfTlOqKBYZXnwkTwRAXBI+mjXOZtxyQ/909ItOL5kHFKI0qR50fKgT+
wX2fbZE2jHGOub8bDr/V6w==
`protect END_PROTECTED
