`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d9ldEF27QJfvcy3gAYIP2OA4Grkk9qI43hAXIM6LBPYSc3evLQyA0m5YqJy4ls2g
NoXsLmPCFiqUAGdiw3VmeIowWVYnYkR973c+H/li7XLuEi/CVJ/IvSth38GGdiPH
VuBDesAlPks4oqNCuz/mmTw5eK4imLjATKymLC3B0q5wHaA4QKBaz5FuxisOQdUM
siKqkZjOMI98pB8zfBsCAUVI96T5fSLDtrlYf4ZV6lw5YK3y2ZEXW70zI3kIk7Mw
PCqWzKkJPHn7/Z7O5ZT/aw==
`protect END_PROTECTED
