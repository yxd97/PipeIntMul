`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XNbWU8p0Oj+d1KKxOq2ezv9mD0uFfOxjr4SgkLyR2fsaSDxTwsT+xwj6m5MpLwVP
5PwSFa9tJIi4/YnP5iEAQDqZ8zgeoIBtZ1JQfxBUs5w2FJB0mz035x2IzAVZyCNh
9uB5En10IhOqjfWnrDm72qKABXOIci1egyExi0SIumE2hs7EfHcYvgKGq7Ajv2Gd
DCfnFDKRc9XXNxfkqxYr4rZHjDDZgIoZ2mQo4ACkl98iii6lQNZClpoBPNFBXD84
GKFuiOGsnQ9hY++p8cno8+iHOTmNfNtE4JsqS8RVqcUCdhI3URURknvgOJZMzym0
YFCXQ3yWKCfysEAbPH2qzCc0v/I7K6pKib8Zn4eSfTdX2Njo+Xml0OWXswZclL/e
`protect END_PROTECTED
