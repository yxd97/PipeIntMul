`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r4d+qsPDOx0uqan0n0YJlJM3D3LBTvzzxHYjc7kOmhLRbxbqRhnrWBdSTSJDoAdl
zDNMBdi76PmE+nxX66jtx5O04RV1Z9gb8BhLaHrq/c1WoWp/hmYPptPs1yjROvQ5
uI8QRh4p4S4jeQyPiCywrgi2dPG55F7u38iUSAuCQTw9Lxo5EwiumwQrFnu6N4eb
JtRr5NU4VCgQuhdjEixbWgeWd0FqhaaLSMcyyUS6kHv3NWOFovSUn+eSOJ7SwFvN
GNWnV8VVVwl4waFHO/qArWAec5//dN8vcDu93F9U5+hGQHyeH+MWHyPh9r4MBPX+
ZFyGCe5fjhPcj52vpf2G+2PxBoPUfJeUK/4Zq4ep69IT+WttNraZyWRqA6rqgKLP
xf4IqD+LLSGisHg1Khse2uy7eUF3N8Ir0XOjZ3e1zeARfUg8wtyFPCXGjB2UN7ll
icmMsmgv0ZE37IOh67FZWcRLzbncj/rPR71xfu6swB/p1kH9skFQfKYur+PA/l5H
S3FYZ02h5Kzq7O0mu+T32djtNnEGU9OKMEV0lqCUaIQsYXe0XzHEcuIPadKj40qn
aVSR8VUw7XuinmPqf3JHP8Vnqr4TYh5VI1k/9Hn4ew7YhOpXtzAYa5iNKEcrcsyl
8aWWgWtJyiF4vpSntm4Rt51s8rmMqT1Nw6lKT6Lehs0mY+NJr81s66abh7ueVQNI
68tcsx3LLeJznFwLr9kuYNn/Mn3NIhK/WolfV19oy5e/LZsaCq8V1dv8K4RtyHn6
z4hq9Ml/VflTAvoXz52R/A==
`protect END_PROTECTED
