`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DffSmdNQFeV3fIe32m0CwvC68wCNGKhE+ErC+zIR/aasR76pqGlcQHNh2Evb3Hr2
wEikl5M7OuTT5qIGv6Y79rJu8x57bJcj3wzruKahWk4zISjKSQmM2wEEpX9x3b0o
WXvoVhtozUjhQY9Y15ULxRllmYDbcxQD133XAr7anEAdCcNaMaHEkDHHcGDf9swZ
AtOl4fIeQf0q2pGZAEELa67yo0sUVS/i5GayUjSty2bnRZtLi+clwciGYV24lpPy
kAlvIZksWedWosTNUL8gpdUEY6Lnh9aREKKlMgHUT90EfoPzFnUmHPFOktCuih/F
HVeYz1Xv/zJIOIMiLP22gPElqkx6D1gYiK7rN+0kKJ2rWJOBUQTVEf0mL/qmuGxi
Vu2YTtSA0aKKYZsRNwpzevSuNsmfh+33ToRCIog2b1zrDbtvFqC1YbiMP1ckvxcJ
zqjOS/mlV/cVaLvVtkqN1bUKrPxlq9vi4W0cEJqM31Na4JQ81qrr24kkaQgLHSjz
CY7zIWP1Ix6Org8+eNbHpgwMj4qkiP+yKR/YBlJgb6awnueMIfm1gVqNcMuBASGP
wl3hrO3zIKoNe52Sn5I5l+CQ8TJy9ZL35h01IHTSexnyWWrnJDZ/7oWByNegR9/D
GaOMVxcFTULNlXBXMMOg6egnDCP8P71Rgi+X84nks9O/2I7X+cgcayswyPSvtEsO
aGgEI7TLHJe5aUZiWAECd7c150D9B74KDfRM9BIEIYXydf3rD0LW71xXJWWznQ7A
m1q95rCS5OlbeYo0TCIeWiy5wwWY5bldoExqrXy421xY6TNyMXov6DYxb/qXZcBD
O8ZadW5TDVBjG0WJrxx5taiL9xBmGRBAgjWwU9D9wYkJL8mIHBdmxlnslokp33PW
oT/mBB/OhiIy7otG8IXNS+uwa5/Fqaz2bEmAvfU3ZNE=
`protect END_PROTECTED
