`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nk1DAKFfnGKd8LxbgOr42ZGvnlghg+zSBRl21yWLQdj6Zd9btFAH//kgYvb9zlck
FcUurM45dRLWG6eAPni/n/8IyK06EoH3wBGRQ3R/gdiBHxnybUWHToa7TxGV+GCy
DejNW3aFLZhbB6vRiG6wHEchT42Hj+GuEbnVtiZ2zY7y04t388WYldBlJB1fl7PV
7zjAVvMjAg4lX+hfxaIba1QSaIWfguGO9M5p5Mi+eJ65W4gFu0nOgJJod3pFIp3K
dIEzoVAYO1vFXru1RyxQPA==
`protect END_PROTECTED
