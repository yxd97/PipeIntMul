`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lCj/BuH9myw78TqA/AZvkHcZ8t0SlavWkGQrgOWJmNQeOI5Jji/xqssoq0BuZWWB
IYqI/7wCATRhj63/xkhDUm+yaEk/+03HpQRYvl0AAT7tiROLpAlmnBc6Y1UNI01X
j6j7b5RpFJvHOqVbed4okNggpWX9kZ5m/PMZARd+d7tDQfW53aVoLSTtTGGeXC27
zXGG0wtuWD0ElomVpeh8ej5x5NcWouImJIUsre4fuWRJ4dcn4ibWPnvaZvWpkeRE
NYAoQ3A9wT1AUsoBbdcwMg2T1i139UMLiFdcbLDfQNTfqs1B1V79lwtO7Z4URn6e
s6DpeuniGo1KJ5azGII0qQcNgzB9vPVGHCxxlfUsjXKaFd83ypVbfLt5AerxThpl
pEM+6+wt8eQSOxDAXW5ddDsfv+YxKPQ7ciLkyYph2plg85oLWZh358ZCUx1pbjGG
pikf5+i45NO6898Lc4U8iuw7kwe1UhZpzMzoE0VF+hFtXL3hNfeoqInY6hDVxdMv
rzglW9SY87qz6Ds8qRmXeYkKaSlQbrHqFYgYJ/A18rMmbVvBnksr/YAZls0v2Hcq
HnBJ63T5gnHrXJ3aVa5mYXqg2rC3jIhU0NdCSH7ePwIEVj+IWwm8yFDnP8THbpw2
M3my/TVQSviKK0LCC1jAbUiDlMA7hNpBlp/RR+8hE8mbH7EmiELXYoaDlObe+RgR
qryyBVw1TVf7yF1Z4uZBaiCROa9gnzMOkRCSN67rRF0grOLQDsQhInpXbcEJIYBV
cA1ZE2s/LujS6j5VVQpQBBzLWmypl9B7t1IxK9UlG2NCF9VREoSv0fyBuA3eKegT
gwCmJkxDwOI6VKEQGYoPdg==
`protect END_PROTECTED
