`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eUYelCL/s+AQIMrrRXAobiT1oFQrA/GoXtCeSDuFa/EUT759O5QCqC3bDnlgKO+Y
B80dLam2MOu16Uca92dcyNo64CPqrlSEm9Ktus4wZ4U6CCXaqfIcUzrvbbXU5WjT
XaAp4pPqiOOaRfFRqKEU5ZzqkQxLiKOwQi4rYeAqFKBMNp5QSM28nZmWOxB+d/UA
NtdHPE1AEKoZPpncfB/t+3pf3XFr6tgvpcBv2bt6vJx6Yg4JA2xG/VyZjJ1xn9CW
sYvT6cpgB1LfcOvd0Vp9u+ksXDZA18soXswnFhDVkddT8rZHOzlE+D2qYEZJ8ljq
uya8Ttp1VDN6VWr7p/DTTAYyyyUGTejPjYgMPEkymmxHhhQW727E7EDx7rzJasNx
PYTMSzdT7PgEfRYHx0bMyh8V0hdvEMOaspkyFcJTF9N5q9CN0oZZx+dewixPyHks
uSqDX0FZqU6aWE6UKml/Z+w2mq/DEf+g8s9nUz0qrQxlRYtwPWlrSzTtiKeQj5hX
oLTQXZG7XxWreJgAf1p3NkgC0C2JbgHEQA3kIo4IJZLDN97pAOzMRyy7KHeFThh5
MiAhbs34FwXIC5h6VZv5QZuj+cPp9ToO4/TXxgYe/zzKXIYdetDZVX7LKadH9Zkn
gOChbi44ff9AHdn+Llt1Zjy3i/h2uy/j7MgFG90EgylGlNO7dy9oVY+OjbJHd3f7
0T8ruhne3eJcdDHgRkES1vzHNMPNlWc+RQv97m6eeuQfu4sxuQhaZGlGDrjCJSTt
j/hb04YuyBeaEamI22VOYEBtQ1anddWwWFqk+i/sQF7LqqBL5F3T41emx0gUiKHj
9yAj+2qpPEuYpyXBJryT80GlE5VwW3bflsvoL/NMBi0eUZ1r8hi6JIDFW/JWyxOz
/PiH+uplvw2+oqtju7lzpZAw0DsqJWZje0k3IQT48I2JNlaP3LkpbDaxHPs8YEfK
2p35ddSo0BQDed9LcuW2bXiAVyJOKURCy44iNn4oaZmNRkzFf8wXo5VIpDyr7E4g
Ig6MgK42OrRKXOMKgUd+IOAwai+zyNEhULuyD0DyS3c+mxge7BwXRWIe3Qp09HUb
n5yizmTrMeY70u+iqNmFyL+fHbgIQ7NUkECliwo43M4dH8dCikYwdUXvDfSR55SJ
fNJq6JsvRLz2dbQsLDcjIk8Fd7tjmOCn13jZfJpyyAXC9h+TGG2IRTv3dr69m+AK
Z0nUvb8YL9ADwtY6QDYM3CBxKe9B7dYHf3kXekUHc3tLgSjUVxAB0N23JwbtTMj1
Y92pKysrKmIRd3nk0AwPO3IEZXbo6YbAK6mbWb+SWHfx7+E1MSvtTbrMYZHOY3p9
+SqNsit2Ps4jOjj8yIX8KBG/ioR7+XOwMC+ElhCfgH3g3xmP4M6OdDATjEXEwNnu
pFzRvl0/PK+4o7JCAvP7cSC9qQP2rDcZhLtUOptRk0SLeaZPgHb4dK/4tFh2yE5p
uurL/10vHz0/Jm6oQS/kHTPnj/9PG7DPzTZpaeltUjGj2IMVRcjra3K40lvMngXh
CoLDfG2nDTVcb2FzgUKjLk+uvQxVhocMjY2fBsQL3I/mrXQt7pR5lwZBD689ETVj
ekvlBhIENmiU4YbzqEeJnTi8VoPE0vB7ebkdxQl/eQDPfd3eP2DGDpaK4KBOnAxi
xOCuUzD8Wb+ew8eppGJjyPx0IydOZUz5AbN4cy3hcVAn2OFV691iSl9qV34JTMUP
sd6Xp4nqPIv09hx5Te55BLMZB3L7CZydMMJUaR+m+6d8V1gVe/22Ee/CV3B5S0Tv
fs9q1H/4ICPmg5lLTv5DdXJklZarqTLOs4O7Nio303zXnvUxKT1uZX62wL2isDhI
TqEeQA7WnRHJ+4gXswtZxM9AYdqXg7SZvDK8NIVqJPZkbaT6/Haemq+8agOjlRng
hGASrvlIHkkPmJz+wJ6lSin9/X48y/LJ0UZLeSSXkZ3zffcgxrOkY5DZAQMYdtIl
Gc5ON7mDoBkaLLmWnfOuqIPLaeL4oDbikM6oE5/9s361CksOCYdvxJ9zSqfmVlwN
dRjCYEVhfYjJN+32daNLwFTcVKK/+xtYCmxqWIzeMzIivV8YVv2D9VOq8Vgsp22b
XKW9bcK8evV6kHUA/dVXqh4s8F0paFUvlFASWQdbx+LREoctJOaNjmvYwugxsgHa
rwXmCU0AxyPEtaW8M2gcY6i4AGajnQymXRp9Wa5WPeimKv7XhGycHf1g9MGVOPee
ugiqnj/lCMkIMeS78VOgvTiag+jMowVx3yAz0QVtHpY=
`protect END_PROTECTED
