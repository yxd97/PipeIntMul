`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0boKK8FuK8WMtNXIjVnp5pQ/XSp1IK2z/fBc8l/IOQvsuAAKeBcQ6aUIfSela/hb
o9euD4d+e69ze885ZkwDvjMIXsGee/9vKFFw56LwUNEv+sBSJdjZ5CvRlDSWPOQt
YOefn+zUuwswMJI9zpFt6qjrnpBYCVMtIcxisxnWOazAkt+nxUfDnfG66SOMw8yQ
Ams/pAmg36cdPjD3l3MYVsGSaXq2qmIhsMCNJyDwDKETBRl7IuAv+lhPedlcwjZq
DilInK6Av9CNpwCJjzxh1mwHsm1GIQEQi97eSo00XZHT8PteKoCvNMkxWVvGeX/U
zjxX5HpU+2CoAeY/ZOtE5ZNhxkJpaDLes8TxQbLjxeE5p5NVKTH5gJWTrnIhrRqD
Klx7uWY6worJI+NnwE3Aek8nF8ssoMoTLlz7idC8vzKZcukzRmJLRDfHvh0pvNm7
ADFofc8KQozawr8/ZNT9B+QvJAKANrCnc7beaitx7PqNX25SBA5rg917Ff/BeLkF
ymRPrwJLR+3d06HXHQxMkN7B48D1hGjl+RSwCkz717IeUoNsits8CtJgjYXQFBH7
lb4xw+dE0Q2uxafjtJ8qz3RfwhhlUNUgsJ0FX6yhAEudBJOk849SWds9nrKGi0eQ
WbH4Z8gVdS30XUgNX/g3udvY4K2/x/d4NMdWqLfG39hD8ufODXiHo+TIZxwNWkog
w/7S6F9LWLgw/uOwtcS68R6hZKAbgQe2oqpEPce4dRR8rBk5UBG0VVmS21ylxmp7
Uo1igA9RcooMQUTe6IG7jA==
`protect END_PROTECTED
