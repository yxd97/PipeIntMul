`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6BXy4q38XXP9FU0TA0uyZawzs/8jClYvm9is48LeOc2PVfHm2EOm7HQX2qWZlYnD
ezXcWwFSpCKiebAFT1xmqCI5K+0Fho30XFd4lNzKNxOdak2RZKChg8Xv4rB7Qumt
9lZ999Gm9YsSU0wwC/Nbbx9jwspjLAmY6Z7sfH1VQLb447Ne0Curu/piDPoIaghF
t0rayIV84XvAVDsQa4yXwhRd/PESvBZDaqwhfvbZAuDlcknjJ94Nw3lVQeVH1uDA
uuD/GqDWorSNoEbV2pyRlmN2vTq6sboHFuy27QMqPIl/o9klpu1OxVv0zTv2eVaj
FHOssli3DKPsJjGPYaEOCQTfXlTU9dtr+jGMAIPf6YR4pKHW1uGUG6atc4BIW4im
ZKPIzg8r76j+3SoT5CiHyNZ1PIbLknXfvseZjrAJpNXAVAtTEMIjU/Axpd7wA5Aq
1nAGBkLu85HpHAhozepb9zy1ZxzI3NLzmsEJ8bhpG2+D+9kUoY0gPe+9SWASOfMf
AGh8nInVlQSfdvOsJ8sAPLOS1aBt7FLjTFHzhSUkHyCYAlRvIUd+oTDP3XCTDwBs
J2i3qnNMSvUcmVdXw4pv4/gGkMUiOGgsddYpxIstQMDoLHfQZlpmRwP+U2+tWqfg
CbuWRMQGPg5c7GPRWVQNudsmecoXdoGFwO0uwCQpc4QEdcKq7J5BbVLsUrewfVqx
9YjIm5/K8RQeGcaWYjDmUSg3SIGgn5TbFLxGnMiIxtgRmN/poZZwmLNmfBiVn03V
ToeHZJYQgWaqHPxG16jKclvd0qePX9/GL30RpKsTLkRpbawaywdQ8RaMz0+tN1eK
uSeflct17rh2UA3A2p6LXR4aqP4CUSuguEpr/mkT6Z4=
`protect END_PROTECTED
