`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aU0EgLGghGQgqF9KnnqdVdn7RV1+soGW0umJZTMmS96FTOo1hRBipCfahe1T6fNX
AuVRaFpL0A6GPv6TEZmA9vSeJjPQiSasa2oXdm8RJfc3xg/wh97kdUmSSFy7kBgA
OEvhjWZeIlNk7byWffOWViOAxocC0K1rA+rtHgaqj0ez6Vr/FE00V1tlZ36JChvr
LyJ54cWChzTqYJ5znGdHz1nrB7E65EdCXhRzW7r6lcmDdPqRkswwKQgRXz8yWssx
kPCi0IwDHDy2hsrPQWWAH6xb4UW++xOyFlb1vx1FCZsjoqYL8YM5U2OK33bHMoyK
8KiB6i17Qq8UHUVVDoT9XBqKRTUqbq9wmmRNZO1klTZhh7vO5aW7VBZakodbWf5s
`protect END_PROTECTED
