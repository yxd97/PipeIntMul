`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w2uw7SDF/X5QSUmz6zWkw+yWTqoCGjXgPZ4Jfa8wl59UxUKN6b8fr+Tcs3HziDsg
1YQenbROgZaQqLcJ+JhFJtkFntxskDt6VP5/MIcxdW7yzpjPc9ZgZnWmCqk1kK6Z
N7l2y8jcSAknf5B5heLM3VUgTn/9ht34qTcymV9aTyCPKXOnz/6A73i1srKXXSEG
U6rH4fCAqzSe9UK12lJlu+yH312b7mv8pRnGZljMrnm4U59kVLl2hDt91u/VQB+/
TNKYmSPyErh7fDJDcDID5NWwtDXqR0b/Aly3ivrW9BE=
`protect END_PROTECTED
