`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AHodL+tV0+rAPAHoanyXQb3vOw1BHYshgOcoV7UIl9YTGs+kx8oNP1IS5xIf3aFe
THObTbNe2RzrX4//hjCrwE3Mbd+gzq9aJjcmWhsYs6h+EQJ/UxvSSt/cEj8YAAML
YfbjE9aMJwKUKHvD9NzdwQ4G6xfeMlCM5hx/WvL9o7xthDked3NHM51yAV0OMV79
5aDHOYmw3vRi2VwWqpj1bg2hxAwpYMG+aM+plgqkt9JrYr6CngHY4ukgv7uCxWeK
5BCO7EtR82b6ZaNmguuK7oLuP82EmvG9mo5a03xyHeH0y6NP1Uriu2MqiAjr+iIT
kXq9mMYy9LsgdFlHNEO2zVKOvme84JO5FiH+8NKndrn54wMtKPv1EMk89DViOCIJ
kkUieUKLbDBtL8fiMWDp78sD8TveVUf4CWOZwA+wHe2ehabt31dPuBpG4UkO+RLZ
c4Ar/3VSyHHLHOav7BQUEVn2tWM2VxiHHYOjaWJFwDpo1XLmbSEpUgxmR7vdsxRz
KgW28/oYpwN62AqXZP5KHmyUlYSpra/IWjmPuQRt1LgCjYhvLRroB/h5plwULDby
ezIU9btSuIxmN+mQztJFtmlajue97r9NzHMJdnIOwWuLjlBk02ErLxgnCCbhYfI6
RUx0K8ERtocERqH3C5z6n/dQ378IMnWlsNbihk9MeBJrtJiZjXaBA/KCcFFUBVYy
p6H+KLTANI/zjTlagZHfDSbWRx2HaYAIzg5amgBsZtvkHkUTC91xQwD/7StAjM2V
k4GHP+0/8rJg3pAUvsC4cBWPfJFoCbejB4O11ywk1p6XVJniktqRF0bFq5Tia0do
hqQV3f2CtPlXNCe8R8f396W7+Ef9v/DrmMdOnphwkx4=
`protect END_PROTECTED
