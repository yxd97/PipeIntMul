`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n181G7czd8hSmw2mdt++hsUDGsKukMp8s1pevq1HRCiDq6+Fk2Tv+Z1OtytGYvaQ
/6E+5H9rKwbW3LsWQghZRrYsB00nxXz3SvXPl9ppBWvUumTEt8ugeVi6v7C0kjSZ
ERbIJtIPTf799EK0Qgp60F0p+lP0TJ8pXcSrJYJOQ8PHCLiMqAr9SyIdAgYmttBv
lGJV9dIEyC0lY20dFKU/7aAHU3Kdu+o5MRSc9RJgLtu2OQIF23VQiWF+o13zYXeL
bMW4lBfigz7piN9hssnnmTybWfco0cpwlhX7Oc4Vzy/SXkoOa9Fbp+zHcrJ8Tozf
10L4oXnUEcgG35cHwhHsv2xV1VF0gfWOfMPfW1aCCAAm7i92JThLg3GtuGD0uDV6
HSl0bxvY9Qp1RtEIAYmTVfQ1SHdP5EsmTbmkysH23I3gcFStNyDp8A6s724xX3xK
cwIeSkFQnkE2x5+F1T60jUcoItVx0MUu8ct3U8oj96twpeunQabeFQsk818A/nEl
4qSsSn3eYBgTOFy3LNkDANYjErjTifX6Iws4HdK4ixj3yt5LxhlazdoFxwyYKLIS
LXLO5AyW5VTj8WnkFnseLCzd9m8mB04gVZDukffCFxZnhuu/pzBgO50V+NdokmPM
NzSx8glHIk5etX5Hqb8kulkU6sTexioTd1CtYWYvdo+5ZVCGVeBoYHzrEiH0CdkM
I+2cbqhu6x2cMaCTk9dIewQgTg0gC3E4ds5B+lHTf1NERXyMBtkMPNruWggXDC9h
P1ewaE3Iym1ytoJCDjB4FBcwgwd2pjWzt41KWz9YV/3rb2MJpxnwqnTDYX5QsHdq
KdS9n8j7ZQ4u13Q7wqMtKGbMGgs0UZneTfxob4CuPs02jIkKsRXEqTp7juIive1Y
zFDfTC6sbXkBbJpbu5xOrRO6u93YsPYtQgiTIlJoGGFu5qd4dtIkVair1LWrcYia
GFxQIPxcoSPOprNsD8jrpj94RZnC2ZGA2V6y305ZbZiu/Ql1Pq0brvbfiubWr6q1
EMTaMpjxI9e0/ySwaCbGQSKWj8kSfw140pEmY/OUtUx86pH1FOhWSbo4FWB49Enj
jlBMwmRKzO48Gu5NyAcY5IEJ/W2iRnoD/IdTyQf+TzxXLs8D9JvknueaAxnay/rH
DbSbeX1e0g2UbU0bBpNY4BChLKeuKlf7I++VUK4Ak2pPuFAVksBQkE/wQWEs472J
59Xnsco9T5KyIH1y8i3BF7P+LxXhZVh4+p3ttUjJJoVcnhLX1382NkjR+M/CAhwY
pwfTTbUiFc2+E+UTPtTlCTYkAgxL2wU5NMyTYf6jR6Ts1AM2dkbYfKKNCiNKjndh
WeSVgKmzGG741rr4Wv4LkaLY30EgXFwE7KGZCQ84B64iz7n+5fJ8yMIOjWquABp9
luJY3jqnr2Bo+Lvx6wNTfZ6rEcqTEHcckkX0op2wuNQberiyCI64+in81oh7ZqlE
7QAfpl5lL+XHd7FyciCT8n9sDW9i8yOJKw1FU2l+85fAKzTRNn/n+TQeoHkdIz3E
76VBtOL8OXSwzqW+dYBU6tPZ8cBBM6w5wt4M3/lkjyEjEC8YRQtYUppxAXJSPxkV
6R4p0lXOwvT7rc61ZZ1VHdD95a27m/sfWjPiJDFEj7RK3n3tXvV8oa0ltZAOFgdH
IYvYTRRxZpL4Q9NCuFtFR/T1TdeDD/viTY9nCRuHOg8eNGN3Lv4OzNIKzHi/78sb
BdMIJD2fBi9nK1ERbwnOEfO6CbzsLFOangsXdu3luHKhmf+K1x/vSfk69wqYuhcL
+lnKCZTuflDoi4Fp6AH//fcX468rYztKV2COkmJAKfK/wy2WIykpMQIXcBbXoD+/
VpBNJdRwkAHOuyjNaJvATjUiFm1qajwyw1Bm3vNzLR5tYo4PqgMr5pl4CvvuqqU2
vCfD2xmpM7biHx/Gvo4oKSVa2rMvp6nQxmzv+Kt06AyR129aUwHrpWbmDalnuXLO
Myf49Z4TJvkEg90K0INA7RQYua8BCDMYonVbcP1AOM7V+TXroee8OUUOZkDtwUhY
JH3hViYsCkt5Qa8XLy8FOw==
`protect END_PROTECTED
