`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOu5JxpONyJusyMQq3a2EbzS8gDgE77Rqkx0NGb3k/o1IgOzxgkhGTGUzZ0n/y6f
EPI1yvIFj5jHbM78fA49fo04V+8ky3l0hKxAqtno+t8X/745q2kjwoX1dewHNkWT
n594OWSQZWslhqiqMtnmDAtBzyT1Jl1cfZRIJbL1fAq6b4qXtI43W44Bu08wdUNq
NRqAXYBte4u01uWk2G4DBeP5p1ywdl0YsvC5LAkJ/lAbPIHwTZXX40av+R5IpFTe
pJcFv+rIp9t36QiizhsOoOTgwsVKXzp8uRttI0iu7OOls0z6LvqSitjOPM0pwH36
vlw3BhTo3As09crHk7ldnz185kWxKZ88ZcDej2zGjUT2E9KNK6gZWYcHctod5G/d
GU7qNIPIQO47gSjBB28H0kZIIgFPQVLR6m65fUFM7z8=
`protect END_PROTECTED
