`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U/Vbc3bb4Pi2FqsNUxvIq+N4w/A05Jwes97PBefaPE7cBSRth+MDEZhxJ+9bz7WT
lbFRDqN7egHjAcG90ZTpvsZz2JQ8EedgU6+NlVihcikc4JcekZMJp2W6YVseHE6S
okkB3t8ZvSG7A7WM65PkVuM0haprWstMcNgY7XYFPcdq8zJ9VItsa0xng4d2Px0M
y4fdF/+yakYiYPt9c9ty5F8p0+8yVcGwjArBVJX0qnbFpmw1zF/onMSoAGLk/raB
yIDt0kqGW+0VYF+9w0Z3h7VEAnnW4PhKGm9DNnyGVAl69BwqaljJrY6e6UdRrpnR
h5ehtNVL86Sepsb97dNLSRj07nxo3u60dLBylEjQ87tuZb0O4G/fxCWIcfZ++xMe
6JZYwbsgNWA1JQ04v7fDCVpgW2HwKgV0u7GYkY+XrLviRKFCLwGWO4pe2C0rHdU5
vVcFOiAEE+A39z/pVb+TQUjrTkK/O77HIgu6OIhqpkj7OpL4F7PqCDd2tIqIzflK
hSmw6PDvgF6qX8QGkFah3i8FEYlGxqj8mt3K+zv8FIGRO4Ip0KLlmb/jl0IDLENb
2XZt/q4/258ibCfBmHTzTFhv/dVJRfqUuX/9Xe3AvxeoKbB2Y3Se0oucSswTKiS+
JX+ZNrTBTw0iC0CR7iCuXUE0r9BE4EWkw/WaguRU27WCsyKl/881S6BP9PoZzXSp
4pErDILKUL4inOSjeRAqlxQ/h8szYLsVMxds0fJrvECILjxJealsnbdgJvhB0ppc
OSMDl7GXuhaN6/9sZ1Z6pWgqTw0E7u+7pMj3oXAR+vmrgt9/UmDUGI06CyxM4t5D
8plye0uXqOa3nxWpMzNdhCwjNHCeDV9Ki4HQMZQQnzjcfiGqIPhVWsTh/8G68M03
BUT5E3jUqhFhebkV7DnJZQuS6AZlKeDo73SyIES0rSYgNOq5EhBnMAjZ06uU6h92
SG4RDqSzymRjG3X2aHJt9iNWeaaL8vV37Qin++djqF4gQuQxvsbXYf/JKC6sglPC
Eb2/FDASUONED1DE62Vz4wAQUHVX22S70Rf4OUy02zaNVNZ2THN998wiOniu/m90
9YSWAPeGFyj8gIUgi129Js6dmV/lWTsgdR1Gl17gLCgWoezCINh+iUBP6yb4sMiz
`protect END_PROTECTED
