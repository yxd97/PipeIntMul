`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dFhg6QuRwZ9shVFc+nZ+WUon1prQXyVjuz2bPwnS5SKW1+PWwOCoXmqhW4EHHVBK
kwyxLV2/aNYmtd9sxf9Pwg7GmYZXCkqnY9gYrFocItUfvrzklkDfHFawCZbvyuav
x63ZfWI9wPc0UhXr/zM1E3sk2nj70sWt5MpBJ/wMEk9GgadWgzATBUaGInSdrp1x
dI9ApkxstK9/IJX+oljvKPvhbHVTf1IaZBsMZUEwOcgJMqzFg2N5ReiTX+bWjr+5
JtvTVhghP1o3Kvib7QudMyGDiusE1kJ0WFi5UdG1cYdlaHYGRyCVIjilFOo2yWj0
epczFzUa+yRhbD1c/cGZtWle1S/iIeIZybBQY7eyRUsYgBWCHevUWjF3ZqeY+qaQ
CherTOSaXPHmrhvs9dl8ncVe6aZviDoq2WtBwgrT2Kkhpigb0Mtk+pTzArBM1jFk
QUQwQ+Z0kCZ4NBYkeXbAFuhLvVGm7BLBbDyzqotvNuoECnKawdwVsS4YEjS67TYR
2fihTRp1zMop4bPEOYLCOOOF/crWEy+XUCG+84gozO8NgPb7a2s/F7TYIVXdl9Oi
C02TwZhdzSHC3mJKMXn5MWRIE7gF3keEGP4adHUfGCd3iXUDeoiEd65q8f47Ise/
3aQFTn+fTlKbZNm6RtW0u1SDyQN322mjJSC47KQKmlTohw42ePi5Fly4W5eTjthE
UN2vrhYLydWKkWbPWeTAlA69mJuRsGM/4I0qMy3VvHrA7150juL5VxYaSFohoy5+
SOXF1jMRBy4bGedaXfLNzyKCUjK5QndjiMYs2FJbaBbd09/hMKrldI2JgmjyzaAR
wlgfIooVIRDCDAf3P/SR96YQ2TQ803sSJmqhvOLrKOB3HXRuSSyy6QSZdzmkI+UD
v9FHBUHc2f9lpBsZ1lECsaV8M3KT8sR7Zv5gpg6omeIcb/9HTTnr5s1uM/ahVOR3
lyWUVL8khYFNsjao2vBMS0dgMU33+NFlHYazwr2yGd1tEiDQP56JNeg5KB2Iw9SC
oaxx+9Hb1CsZdq59LAO7fVwTaCKYPxQadeMPG4XPmtdumNBNf8f0Dyya/FCq+wDq
sbKnDmJU0zSchYp62yz3vhUR7VUCU1YjgHB24yRCP+AVfwp4Xn79oxxMyiEIlLRf
wKqmllwMKVIECWbOmA5LAn51TLiBjCNT998DuhHyybHyASkbdNU9XXjqyKmC3YWD
dCaGyCg56nUloD9oKycFKHV/7M/rhuuKxQcHzoCUimK0iuyeR2CpAnR8nZZM2/Mb
+z/qvh/vXkw+WsWQ/BblR1raEwDqvBc69lLkEaX8YP+3BQCym01Fhmm+QrmMfNr1
Cg98WND1iTdA8tKUiQIlBluVN3qqxS1HkfGg26qEG7SjIFTkbxSV4CDE5271PdMb
47t5cHzWvvcolJ/EJqND+M0oUaQ4a2kxV0NFguGXBsxUeBRArWdJKIVh2wPSMoSv
prEs0qIzB6Qj2gRiKxLqq8tFO/D2RK71LPmefXmoiilbS0u2v98LREH9Zmo0j64P
QWRwhfEyypFlM6INv+x//G9rAAz27NeEPkcS9N5XbwjtMfjFiM4W0CRrwafzffQj
bGfEONZzNKNdyiBH4O11PQQI1FSiOu0rdSjB7OP4WYliDdfEY/sAEZTEQxRzPR6l
u82fXREDujGBttwaSTPjds++Tt3tCycNqJJIyGTxmO9j0/AXguEUqANQqCVlFUif
a0XF6Yo24KPWzYHvyG67tAxbCuMPiV8p0NOz3AqIdf2s1I0rYmLLFYBGay1rDWBV
BmUv/wLJDbZFRpfjRTbqzugouZbju4+HoHzSYd6aWAqFgxe+7UlnNYgL5/w/bLqX
fb9AtwfA1b3R/E4eYdTse8DliPKYciLM8Sd8cD2M130g9cjVPM8UCCWdxxencWxH
RnIyJkE26u5xZ6hCnQF/rSjfj7LX0v7wL3AT8ienZmoPueJodL3/HNzem3Z0lTx5
iaxQblRWJ5I76hlB/d1XMQ==
`protect END_PROTECTED
