`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPDCeVC5AV+bBjXy1PrH2Mr3gxDJiBRT+k+ypEFJ1FzIexBrScbfH11Ac248p2+G
QIwIg7sD2/NGvvjWtg+z8nvX0sTyPxIita3Rq+1lsza5iRNb5MEcmC0vGAivOnfk
eHCdKpASCHD4O7HB8n9TnYqSQI7kWbUnoLg0elbXoADGZCG4/hQdlJiPLF1F5uqz
pWB9QvNBdZLVVwFv3s+dJGHRxn8XDwDmx4PZtUk1j+ZSE1sFZ+dvndX4DxnAwhDJ
Y2/B+ozt6nsgvIF3650AG2ft9at72y43ZnxUSJ5SnBLV6PfJ0qzJOA4ztCwDzeK9
8gg/+PTK5423Sma+tH7hBZ3h1tm+okQCAcjImR34STKx/uwL2Bjtjc9zd2GgaUiv
OpXP5Ta2xgnE3p5WD/HO1hhn6Z2ZwT9FGs3Ofo5xkmSbhmNeXekQmAKoaotHFm+L
Qpc2ALxPZjc0EAaFZT2W2SHl2ZctZVFrjI8tgBT9/354NRnPQHrrK0rFlBeDHAAz
+OI1VOhAhp+mVN6n4vKLtG9Lcybo6demYHSCOEBS6DrvvdsKH4ddLe1np6wKoVYR
8gnhw50FDPP6SqAD/D28uQ==
`protect END_PROTECTED
