`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zX1cYGZfL3QrM25OYBqg2kIXmArktcD4cvIQWT56m0DHzDK63pmqCQrRDrmaSx1U
fIihAzWZPsCil48cN+TwYr0wfVZ19SOV47wFyK39Ctxiy7TgXM7rL7A+p1xeArVB
vHveVOlbx0mr7p1gp/l9lDNrH8m+6VVQm6W74eZ93BnY4SoR2Xwlp3l2yO64BVTW
eZUqhbkL1RueCMw/82deFSpBirkg6vA5lf7BsRcxDH6LOOtSDiehGoZTCfd8bjap
ooI/F6ptEgyAliVOMBpRZBikB4rUdyF1fTLemE1ubnJAtHWcQoZB/pA6pbRbXtr+
Z5BMYPTCMXiAPXfkpdX0MQ==
`protect END_PROTECTED
