`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVdtP/pIQHVA7lhV8V1U2hQliJYcNAnvaA3gveP6r21D9NnuVYh1vFHZIxjN6T2E
Q7jQiZcjnSAWgEULXKO6oKn3E07xYCLqm/VptxnB19SZlG2lacjsGDckFhxDey6B
/3gpiTk1TJskq5kD0gniYRCC6WlAyz52L+X6UNbjHSTqFNuo8F6X6TFe/WYcIm2x
3dKN5CBSvD5EvjXwE1/vfRzAdKWKe4Qz99rKzmUa88mI92CIawlMLv7wCfXBcFM+
Cy0RXHhWFF/4irfrOHmTi7KJ03CKMc6a30y5ZtxyPveM2LYWMmhatIebX2tUpPjR
X47N8dlsZBJldOKZHw/Y1fhFAoSxcQiMsRuas2fn6na8xskOJFVGx+GNsJoOwueW
d7BMAPd188hhI8VZWYmJP+zbmhIhiZEtalBtPea7p0L7jXl9zCV6Al6kXfmBAMYu
Ph24CrZaaA14dsDaQ36zoYBaurIFrF71/mbauI8g5kiDbIDOuR0iOjInZhlc0PaI
jXUkwhHQ7383PYiETTgeRXab8j2x4ntcg4KlFFOQ+8g=
`protect END_PROTECTED
