`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5KJd3qdXhKoSPRPqGyeSv6XYwoTn3hSfCD+SIM3/2XPemKB+KxQM5w5f6Ho/UMiA
/dlYoDq/anLyahzy1Id3fUeVyc9dFCKDHuu0ZNEAXCXCjvYXD55OTZafuKybLFSE
D2c4cvXt1Wi6sGngKeX9TKbtsnZh/+grwHXgnbKvdRf2aXVluOCFtBq5Th0y+PEJ
aLOVxx6Ja6QBidjGNK68cmb80RLfld2vz2Cj1uipooqmPaU4rLslXxu+LwKQoD2R
i5gDpGBWSg4fU7itZhMA4DsxFBsxpVrdx3zDqvu29Yuxmdyew/h31V9g2Cf3t/CQ
NjFaep16y8jFQ2s4XICO0l6Jd014kzcOYdoeWketfZrHBvMRRBu3Va74zfFkB5PK
hgdrfMLs6cpyzDPqejgc3G6nBnKWw3T5R4WWhM5VZwW+AT1hWEGVJqAkt490BK6C
OkmFVC8o0P64eUbfOUZvYXG69n43mjgNoVUAbZOwvfYqVrWm+0Bx0aFYOkya7DTW
MaZJbgmF/T4qj72MRmt7/+k1bRdRL76q796FmEoWJUh0EqJFRZ2p8bxXhcPT8rt3
Jd0I8zj2faDaJUhL+YkW7LFZXmrqr0m5jdmSwgulsMA+39Q0TdeTtMvtHhgL3nBG
6Vq1HUx+i0qW2+BYgt2EYNeg/BAXGYgnjJLZX5xP2a4=
`protect END_PROTECTED
