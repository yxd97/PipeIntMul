`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YZs1qPnxxKxQ4l1vremStRqQ40+Yd5rG2iKtb9Vocw3ENDFPFIdf3EiZTPHAb1cj
Teub5jpLoAZziX0DOwNtjxb1Vs1OYqL7J9b0Q4rZnhpVl35WUarcZfJWmARUcKRn
WLkqEVLJkVUq0iXg1SyjPDJW94pljytsiTPxO004Jrt9IYIir+h3XLU6oZS6hGvm
pDEU7EoDmcjmd+7ylB5muyiZ3Ce5VmlMbToRZw1X2gop6zmRHKjhHL0HAu33VZc5
q8WblOhEnoBXSqWR79SSQgygMPTEUPK9iEz+evyqMixDgtWISEdAopZ+y2FqckMi
IwZJQwAajtD8mwPdJYidKs9cGdcZGQqAIsUhw9sswpg/9yJ4/33Y6V+P1R8y8Pp4
gVELN3mKqUi1o3o/TE76+mOE2V9p7gqg0S4FQkNK1BAUxgL1u2TOwqblf+52CsmM
AdwiJzNCq09OrozqwpBOu17Fd1iKoup5qfjkeDURrZA3F9cxgUv2tX/C6faufTgL
`protect END_PROTECTED
