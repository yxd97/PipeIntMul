`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9V2V+/WO2QHHQiiZG6ijgH2beaS077uMnX5j68ylZ0fbD2p9npK9LOYei2fDIpYu
KBcqw+owC8zY4qUz8fdmfDhgoxonx7QDExzC/Le25R+2q/24QZhsLLXxBfw7XENN
Ny0UxmfoHBnU7PApioB2efZL9/0STaa7olCR+ftqOT7Q4z2k5ZqyJX+8WkaIoeEe
boUzIlN+ITzmgVzEnkpBoSFdYviC6/bbYB/yFiXaXu8VdulMTDA9pNEpTbRuyVPm
ZqUTHkAgVDwegDyeVuTaUHIcgJs4i5EpCfNmuUmZOSNjVhr19Y+lYdGwDev0v0XB
29S5HiCbOjVOtElSY1b0Em4x5VCy+IwUhzUu7vL/Puzo+P+bc62SRF1Oz0zgn7H3
LgYjRzaSwVH6ETZ0g2qZ6BaXoNEd+POf1l6ynDOypzinx4ff0INRE7n7kQKHpPzZ
9UcQGdEEMVdNJy169L/p0BniEbRPgP2olQkXcFaoLXnk3HAf9/WE2HE4rXQVarMV
qZX+bQ3j0S63/qfTQoIxeQDvvgd87QJacx7GULNP1B2GQahYMSQvG5GbwPb+eKXI
Erm2KomWY4NUMsFsrgamPj3xD3AL813xeQbnW/NoCALZGh/8U9lfO+8EKVfm69+a
E+Y6CQrXnf0M/sbcQZS3Y1PeoTLKxd/w4OEPS1uGqkxanUaiDJ2hXf6LVd5UKwmt
uE1a9Sd8IWikMaLiYCGJsUoCL8AH5gCuVW0GfGsY74U=
`protect END_PROTECTED
