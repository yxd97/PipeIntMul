`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVEdPQzulluO0rp7/zAeudkWrsNvlRFgKGDv59FWtdSV772nplqN9Tfz4wYGFccB
qCZ9oUwOPHk5vdF810uXEoprSslOLzoBxgEzNr4eBGpo6hzh3J4zAEyKpKbxVg+8
CvD2q6ziQb/DUx9O6bQdArd66Gy+Iuo9a/OWxLvm2v/JGj6/zFPj0uhBMt3yUJ7u
2dg59Pornivf/n3PxbOCItiJELtKNUFyCAUepm/rKczEkKwIw3zdhtIDbewZ3eSN
g2Z2H3Dfoz1+cLft9L/tqNXJVj47YcCEMdYpVNFTeyy9NTGjEs2gDuBtnL0B3lol
SE9AdT0k9i8Q7pzf4hymQZC3cHK6Qb63M6fpDHS267q8S6EUUnuG4/MNWEOFvg+m
IZwnxUfKqoEmL8+0Uz/fXHFln6C5K/K0+K2xivFu32X5QDj77MtC23kxYBOehNfc
GZrVuoTCHl7Id9RlvSgGolFHy/B/yWqaklMFWXnJQqY=
`protect END_PROTECTED
