`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o15NASUrCEXpXrMLEuyfMSZqLH2HvCqOWi82Klw/0kzIqYTyWtdSa/xiFRptDBKX
hzk80XIGJYo3VSzoNghk/2tLxm63gJTIu8ykbqx68qehcLcw+OMumcz3N2B7e6r9
yrUex2Wuelvf1DtyKZZ+Yd+JORFWNzKfm/36YpnHyW9tFyTGMZ2VYDryu4ky8C7X
LYdfdaw++1pI7Bnz8SW0euDCr2ObJhoC9O1xMY8NQ1wwKTOzy5Mi6Vsh0Pf6Mesy
TR0KuOs/MqdqfEsuYAJ5KbFMyLLwEsdFdiQEtTdfOEh7DQoZPHm6PDCKDLZITeTU
cPR2BGYcZTQ/2JJeC2lH4RZeabnKrBGCkCicMDc3R/4ZEP+sls5qYGy9dMvpjkZ0
ncu/L5yX6g+w+fsU2xep5ynKkRhB8KkrAGJ6QYL2J0dnMCE4vCle17Wsj7ZSjLRs
f77jsSO/XqCohiHCKN+Qk7CU0SmEVBwkwNDCLZZ8mlPl8cvFpmoSeMPa33vnGtG8
IkA6C1bd29arXunHACExKFQb/2mrPW6pJ3tj9XOHVdkI/T00SOQ0L2+gKhLz6YJn
NdtDrnZcgDn3D6T1J3lxGP6BXOH79Glu60AClZDG3ltiuZ1egvRdgnWo2hXYT8dn
djPYGZ5rA3hTEBYF33k0xCPRBNnOjtt+PPlm8F75dBtRhMvllLeJx+lmt+K3Dy6q
db3lNqoKgNfOXGQwRHB7v0qnudzOI2Ors3KvV2tUu+Q+57mumGozPYpe9ZBdr/bF
7JQZQgXBDP6vxVdKoyylpuEtHg2bgb7z1pK0omViQNz5tphsBOWBfrJfJ+IYms0i
ipcFcuIx1NtqkIe0BqVid0KF1epAntw5Iqb3IFJyzwzEJVBJ/7yJ8ij+s70dP+Eo
JO1Gd1e7oNWcg9Yz5BTRyK4+i8XL66sBQCA6h9tRETWWOujjx1O55LjEXMYymZqp
uAHFaxHucYNd3raeiaqQSBY5QbTrI1odbzRj+k204oM2XxeGq3Zn+qoe9/8vSumR
`protect END_PROTECTED
