`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SEQU4CrCbrs9BrHKNKrD+TByzfEEa/sNqmxXNO4/fVrVRYI/WEIdgZ9lc0F6TJAb
XJwG7WL1Skths//LULfGHxtw91tsLZiruqph5ZlzNIj3OhBa8Cx1ItOSGjPPp/Dl
ccGcCz+eKp006wQrZI9y6L1EhnirJGMZ9DWmsVbcjcxHLTTsOkDvq3PGr3NyzBEu
VOI+A9m1l4B3vCv0G0GLCGlCWJv6lUbkDca4szvmJ8GbPXF7L1vXBB2BX1g/3aKz
3ZBuRA9NZvpBUVDidijr825EwJ2uF4lyVNN5/lkprzy15AAQXn44TJ63RCHK+QkI
KXozww0ke3lpmgv4McPlDGaa/w3O3mpQCwvN+ptFU0t1+F7CnxPamRv404A2aWih
DSDP30nsGVPcSjd12uF4yr9i6zyjYlIyeFGBhOqbj9t9ArOAy5wdM1O/NkDsXIJ1
63O8OhuY/ZNq1kMIt4k9aOgko2PZp5NK8XLEjiIqT8y7rloi+zjNdu1tzaYqVSyl
oc5+sAhk0c98Ns9sU+HYH8Kt666snaByGKXLn9FV3uVwdXiM4quhhODVmHdRa0Oj
5tedp+P/z0vZnHP39ZDSgZDu06XdlcXVGi+I/3j1nMTZspARYK4UNRGiHqWjFY/6
YEJEZRmMQkQ8OxJyGC6R2EeBS94+e3QgkGjUE8UpvUDS9ZfEtNkrhjkiZpZVVOzO
FRCq4FOBCf9UNl3tdLnzW2aA7diLtJcoh/WxdyTWZHDgdOwPQMzNKv5zrgJkst1b
M97vM//zE0SifXpqgTgiCTGp1dqa/yqbmX5BK72WvFZbeKsEXp3ntrJ+V5dsjDSX
LilpEgKeeRi7S48/4tZB2g==
`protect END_PROTECTED
