`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgP+NB/e6V935dHh0n/oeXbbMRtMVt/t04Tz5M6O10g4qjLpTyoIm2UkG6J1YDEq
YiedW85pE61rvP46DTxfo4YhP+zOiSK8XauIGBUY5cn3RCQBsyDgPx+6Fyq7b94M
Tv6jqBSTpR8kcBUMCFP5dqDmu3qJL+NVn702nMnqUEGrgrkExBerE3d7ZJDVHhgv
Yyp1ejfSO7gr5WQRsn4JupsRNI/3rPMyqvzV6Abkd6BfhD4cfb+MHHEigOKb7Tu3
CqlnRYiCHzeJRaun4qPHEsVlUJIpsvkF2VBFu7PmKBAlPOien5aY+okb58BzCX/I
RBlrR9Z9GOIVIr8HHXKRAIn+i0a5JBJYxCnhqV8NW3U+dlcylXLYuB3PKramYjNF
vx0MPBJrEb1upgthYkbUFfBRcCXrIWSrhYd2UtTkEyO02hu97eUrqzSJZUl2LVpc
p/O4R/an2gFFf/YG4E0nLvo58h0hxmZ38u9QlxzCMIwc8oprelbRsvYrARiFJniA
dJgFE3409yMqMHA988BUwmZtxZY50JhjteJWvP0Y4AEguHPFdinfMJmWZyXv56In
c33YUsJWUV4sztCy4mYjZp2gBrE63s3GB3fGDPiBaOCehWmZKpQQBrC8MC3JXPZ+
L3LExXDupbIWZ60ggVhhPH/cIqON0OuH6L8v5Y0sBvnLJJF2C+zw1Ph9zaAXjNKc
/5cI6ej3yEDJeIgXyDU9/g7FGwFwro2Md9RBgd+4WtCqCwrkwMNDCZntTSXOFtfJ
`protect END_PROTECTED
