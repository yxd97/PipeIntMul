`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVzbvuf/t9ffK0riNGf9G70dWEvoQDRwpD60ocrhZZ3De5obte/AOvxwTzjRWjsr
ptu9tSILPF8WJPMbq08mmH2TeuJ2qVwF+bmaEVFM9ddnEQnuKD+FM1w+MLBcoeHK
EF5hdbzTbXc+V1ZhgLi4aN/peZqq8/dQipdO5P3HJwgBrIrCs+jazNdwVcEkG40v
7S9Kee64JL3iknp92f/LlwIvY+AjL67GmBBPbY25txO226NkPVFUHt7k0BqxpzZ2
F+uA5Zioxl2pNxSf11K4tVX+Tsiw6GYozrSXoKXThyqFpyJoAPMRF7Oda88mj2YG
iZknbkUaSMoJQHHoHkmi208JIzaSt0V521njF9rZHA2wqyKNwT1voXH3gnXOoL46
y3ibtECiIwGXjRvEEi4yv6IDaWJClflX+OSWcfSC3iRPLecVEIHR2XPEIjHSg7Ch
g7vSY0Zxf6TReLMT+a/RTefvqWI7sUkJhCGHdSFY0iBvIEmWxx6yNeC96aJr8Wwc
X+qa2Hffm4muzNuPl9sqixmlUcbyUhx1NiU9pFqMg8IgC4P1gnekPCmG40gNefva
KbvxwXwOfBFejt9krc9+K15Jz0SE9ksEmCOAkJniybT0ie/eDk1KvRMDuFAgXbXo
7wjcjmirxf7K+htmIubkcjeXgECFJK76supjGeBSkThZrlnykNlyZkAY9tZ2qzs6
Bzx2OFLUPs3WeUDL5oJ4ZHT1j+jbd0e9ITh6zx6N0VYvNFfreU9a65hGCiHFrE5D
g5dFWxZg5hMLLwF8h46a887He53TyWwKtZFZYKJzTNuhQSxWz6Xvy+DXdEA3cmbo
tbJvKhv+raSpYmGk3SuvQZ7OvSnFdyQqqhvKCB67mOe/8k8yf6hzC7yoTTweg5Ag
i1n6xyZXSxixe0bdh+vaM9jWzMOZ10WJsCERfYu8xDomXpFxO+ofst3E8YKIifHS
gwl6nQO60m5koo5A2AP2XZt8ROxp7cOBOj3pHsrXRZ+a15K6YwoLRpHFWSkuRZXC
0Cq43OkmrW09NQtC+hhQfUDA0dNtRBhXvmjRvcquMx6HBE4Tq86UQu4ZZxVjvhdJ
YTmLV93kgWzPPSWUr1gljl5LV1r4mnEfMhqoOX33Xj2+AUrFSgSsENkyOldvvKSi
pzSBBfnt9WWOh/18Bs3o4eqTLUr9Q8Lbo4WEJ/IDDBz6GkHrSB3TJiRDMh3pCWai
EfqG485zY9cPEXOTBoXpkkRD04brCiZAWMS3/5qW9CGs/0+uNWtIIxyU4o6wWGCd
xkB/mbitShfL7evehIS0yA4h5gnaUm88w3otAUkxszDW392KvtpAvqn30S2JYwHU
Ytd7NFCC5O+/NwejXpQgGnbc4KToD6LwT4ywcWPRfM0e4fPUavuRLiavtbcmOczv
HDjoVOvh9nza4G0XZHqlOLdEwduGB5sZKyker1aNtQZC9TNrZnl+PawUWBYBnXn9
x9hRVuCSRYFe53Tv4x8yvxCZl7WdtiT8WPYckUoCGt6jiLEkiUzifNWuUbV+QrkI
706u9HSS+DVyCb4e7U96I9AReCG19adXHABRlLj0loGNg4eXcfU5zuq3xj+pdfCW
Obb5MLrau+5dXT9hfDERc9F4cLFoXVIrfa2RTDkl2MA7kGlhvoc/o291AUcH4NPK
Cw8WQcnZHN+AWs79x1Xx6EuuQRyVNPXbV55UAE9poFDBKFNNspzstE3gNvB7QhOf
uoX5uFxAloXWJRG7cRlI2qwK2ryNu2vyMKBF71BYaTN4rLUNqEiFMdvu97DPgXga
diqNkwaWiSgD+P7tr1dj6kb9n3vidCs8seMzQm/iatLa2jRWYvo9obLIwaVyBIl2
WNr8yywlRQi86lIykldUef9ZsrogB4cW1kkfKAaRgdnULlsbTF2kzWNr+ESfSd8j
WMkzTdz8ZkcI+Lre1cZO60EZ3Ti/vqId42yqzc5xwGqoFns9kuHI3V4rOXRBdZiC
LQ8KdBYroHiBRaDUChHt5DxZITT992yR/O2tUOHRgLSp1+3MuPVrqXObbBiR7Pyw
5Yr7OXDe6yhOS7ARiqrAZRYZ9vBLdp2ApZQlbRyMsF5wTWyAbI0nDWioTl4Yrd31
7PKMg3K6ImkxMtyBC2LHOV+Lcd4OWr6VjrSYj8Eelx2s1Mq8KJJbsQ/lImDSlvBt
u22HrovbDkWdLuOg/u5vgro7TmpkBDCgB7+vyVmSemJFcL2BaDejE29wYS1G6D6C
MmMAOJJ0UGbZ7C9m45y3ko+WbpxDgkf86itNz6WSQ0nMqGaFkIOS2fN6aq4AfFBF
txreskdqOaKD7I5EnF38rirCJA5A6YhjCoKt2D8XOmnc7yRPttpE+303RzxP9pkE
yw2+wumuQZNDYlKZ5Gm/FB0989xV7ABBHs+C5qAxryhLNQY/X66rF4zALBXmkln/
f/VEnloD93MFgp2NQG6/OnUPVd7A+kLD1ozkmg7wTlLA0Jt8CpR8J9s7PJFQH1Na
777QCNaV4iEyft5RGFMBCNpPIHOe26WfBkz90GtnWXdQ/VNcRHYc8kHgIVKYV9vo
jsI6pnMmWs0S7K1j0hp0c/RY/oamkXKr2hGwkB/CMKuNbDp+znYVdtcS4IenEeG9
xZeRapPjnfh1zaXz21m3qPP1A5q1cEDm8wY5K8H3QqmnPTdZ5pWzkmX/U7fIHxY/
oojD/C+gnJ4NhM4XpS4PPlZ6Nt6W3pNWdTYB88EOfrxtf5j/ug2z1TI01zNHyohq
qt5HUlXwsxhouV0T7vK2jLUTcJ513keMXpWs6irG+U2OnmNI+i1U87PYGN8kA8mX
14A9sacYIRwknxEsG2R9qnZe1C4eUGgN6OdFCDfMvQ/36DqVeDK5s3/RCZJmP79E
McsMwG1kyiai17Nnd+RQDBiBkL48Lg9+k1ZEsc7C7Sbl7kDtNnqrOnK7o1H7JSHu
Y+FFHwQ5F7G0PcyqK1Xmf5SuqdgRIXHQZ0pPr083yShRlyj8OnY9uKdgvg1zZsaN
0sCKkiOQbsnLKlvQCHHWP92NnJ2XsAi2LFPSpnVlEJCppOQ9+exw6gzTOUrNIZkJ
rzeCrhQnK03IZdEd47LJdk2145jXQT3n5OBcOYlVArCimrm/n5KZ8tG1QczxG9Db
HavvEzoVTzIKnBFPGtE+heYa1Y118Q38J+1HQx5Q2h7P2NP7JgDXTmSgWcXSbEMl
ECDN1GAwcYZ9s/Wd2xds10+mKaRAvQzxyWpwkdoy1a3xpiE/28BuvC3g+OaqlCm8
eH7wUge+fYEDZTgeeT2JvwFNDbIgxpRJEB7ryJrwnwtzsplD8jHVhjz2irgaHlWO
ZwpDqcpldE43R8O3LRv0E+ojyQFCKs2+CxEsrDG1MM0xD2kelZyHtRIB85RjKdAH
cejqe+OfkUjWivwcBMmIo5s+RLHgyQYu4RmbygGayAzO1Pfj8fobP2oxSwIeu2uB
FdLDIm3wabAVrWPjzb0Ni1HCaL/Ua5+y/8Hk07JarbVqBt1OkovsXmbYF29qgFQ/
2PFEUFZJ8FCh2BdY1Y/4vjDYv14vCE86F1NE2XJOLAuqlf62mntLH9QRSsjPQZTX
qdEn0NotCq5nGOaItbyy/nBw7nvyu6JLTEnU7N9P3RtucvsPmSeGKY/BDoot8UK6
huue8BqNOUP1Sii3JOLj6bRieHH8HQWwyUe/arnQ+t9ACgUQV7dtCScEOALIOn0x
+K56Au9iv3oa8KNV11prnx3HebI8TL+B0uEgOJB1I8QKMVWIHP8dRKvkPMrPUCOJ
ona57KHg1OCtOFlZX5gj8SN8zjizlAuJwtr/vGrR1rQXBr9NIzsiOH2gYiv0OsKX
2xPTfYFTr3yJt9bu21KdbO/FgXIvQhSwUVgc53z3a2i5OLKxzt1rAYvF3+XCiQl2
3g+Y0/4eNQUWBDDuXO9yFUnUFDpsUDOdp5+nRQR0OrfS1+l7m9P0vPlH0QQx3m2O
68W5rkLyq38m18TpQ1SZ0irXAZAmSfVSY0pYLIezEyKq0TdV0oisGnvdc8V1KTHn
LU5qDqZKh8Wa5ZjSd0+YO6xuneny1fPL9S5As5+8RY/Po4GULxIs02/vZxI1VhRp
jyoVQeRHtk/VmzGpBkO4tKsQlpj2LsA2ozrufrhLMKpJXmDsZxQDzRJkUKMwQf5o
rz3x86P/T6AvO+h0WBf89nHLnNKJDLQmTJFRODhTMVWAO3uxkddts9PISJY9mZo1
cR+HR2rRA/Pxv3zlTz6L1Jtc3lTrbnnGFuBojj52YXnlZOvNCs6e2tkJUiHwPZkl
S6Q/H7GXFeKkH9I8Dfzxg/9csSh/fecqXQGWUzMe6kUoY8H7czlYPZ6A62WIfd5B
3cERiViTCXjCXafbM/PjMGkOgw3e3R76lBBWw0Yd3lxc3JF/sVz/xUq1hz3aPKPN
akJT0E3QqA7/134oLIYdqhnF6tS7NAnzh0rAqQ/pbD/oK7z5C5dapkEmyy0XqsWq
IDWm7Vw8Lt44Y85OboHqLmGZVBL77HJb2/ejuEKW0H+jCzM1NgGC8YLhrBJdS39n
YKF8bEeSe0rBxr48ea4T/1pJFOkCTFc2s9ia/sK7DU4Dupgt4yjTITwPpz0zLZQc
8mvbGdnU9OSG1ebiDqo3tcb1CSsXHrC9r0Wmvt9jQdSQX+X8fHdhsqprGWcyHBk1
FnJO/GiGrlRGMNOQ6YvK6v07mMBCVE/r9t77gdNTaornyaJxEr7Pe2RSzwxe7O8D
LEXTtlebEMZ7u7K3XYluJytcUogpibgREZWHKfp8L1EXBEwC9GGE2u4fwp2lJUzc
yusjubTkqbeA3oxPUQeYHavpTNPZRlQc9n9iETrKyak=
`protect END_PROTECTED
