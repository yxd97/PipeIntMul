`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YprmanqxnDN+KEZ8HqQpoYrZ9P7LJ1vh6bgamPJje4C8g/BCur5eJWcXjorcH3yB
6PgsA1CjpL4hTUlSSUCuP5y7lMSKy0iREznio0w/rfgoT0jU3XfIykT2eX2d3Uhp
FoXGUGd40odAWdvUT6rLJrXcDCviaPG4eOJA+CPyXxXZNd2+TNH3HiCKHAbpMprL
/MoPgCZka3tOL4rDqv5/EdV88T24W8p+BU1Ddb8r/Bmnz83oE+E+o6zDyaN1pos5
q6SVBPpVI6/kNMtszwOfBIpq81lvyb24Ic5i1RUj0JbmrPDrbT36Mdqf02d5YZGu
vDZb+aToo4peRG20hUaDgWxRFyuhzjglvqAPVQ/ifavqIXrSPgPy99i1steJ1/ry
HI5uaN0cDEzNXfyknnRYFUlF3d312bV5SVxkR+JzCqpbzoP55ZRhRTv3woVgSxwM
MMdGX48QGAyyaRQXHsngwDDsYaCXxJYI0EaGcclCUdqFIrTQvI8JbTpEvpjdovEO
FWOycJNZBD8HTfkrGApcB9NBT+tFEzYCyq6lvyOfJdkrveg9s/Y2LUje3Kl1uHFj
b+50JBCu0XAtqGixSL4WRc6dX0AkQQoJO4Ilnh4ditq8PxMcF5uhQAN5Yzn4cvvK
T3wS8nkbsou3gnSbBQ5vUnlfpg+XPvwEFTdZoI9oSEKfYXy32D6KewJ47S4OfDoW
YiMBNCceYK3bFGtQbsM8khct+z7gfMUIlGD/VseotjT5hy7j88El4THARhnEF6Wn
dZX//1MmnbvM4g86YV4hzkyuxKhCKj7FUXVPgu8SJnzDiMpqCmDA0Yk9rGmieALY
KCpwgXDpCYhTlJ2yjW0irsC5OD+jQIjQpN8FexBbSPIfT2t9f8FKHSRYZhiv8ll0
qAw1qfdHd6GONNWQsh4yZOZaYAlBpN2cVJjQaBU5z6RfnWzYHm9J6yEouR6HshX4
p5HJeXZgunK2BcGz7JMQHroQc8IPdPQeB9ywl/VcaShbxkyb5AtVZnAB+ppFJ6kW
44AoC8piI4a6LfFOaoNGYjsK2A9TSTrtg5R+zMse7mBv/Kf09FlzQd90DA8e9THy
p8VcFkoLKCOOeZGEwLfvfOYzGAx0R6QhnhLVK+aSMIffaE/z8qP7v9JPYEKH1nsr
Luw1NlXH45lAJM4z8FqTNRvNRl/eA2hUGwAJvZIggxW/RGBrmiwE2hbkkQKNeRB3
ZVVTe5i/O6Rx9k36GagsfV9xLKJT8D2NCra9jTaGkwEs2/KrVM7qooaGYzOfftL4
9DW6pnyxkH8sLZ+PLlyVJVxvc8adET+qPzax1MNpGG0Ihi4S0JKX2Hvz48LfH3he
OCwKPDZZwDd4R/TBNOPaVOQJwBZlo2/KJuz+44JJ67xCWc2hhRDTNvPxN+GcmMpt
RfR83y6aykRZFKaMeYgeLCMwvx62Cx5Edl16s3MmgG6UUkTSmN2bTjzetxMThmK5
5W+5pDVTs2UFguznazTtnKf5mH7JN2OLByiW8x2MEeCUEzSF+5gxLKv4x1wtkFej
JsokzfeKh6nNTXU1CCla0+yYsN+M2F8PZcMKx8Vx4zl+aRqNlLxLpyRMdFbyjps2
kw1DT5KXc4DSU1ybEkKBbwX90+02AxMEJwZca/cThZpyojGMCxavOhlZZ8Ej55tW
7FhLRw54FASKGW10l+sO3md0QE5QhdXQO+HSDGFY7jSvC2Uc7WEDhFl8jiyMtSEr
1U4Kgcu1s1G6b2fMm35hAIgJlrP/95oLAdeL6mggvRVnqWh7QMzcEzblT3Te5QAL
Xmd/gzck9BnKGfU+BNgua9g0uawnc2NxBN7w2MDwdhbSz2N6kkvvL7QQP74KRbf8
pkdu+x7NusxwxcxGIhW3bEmbVLggvCQJFoOKRBvwliW+aPFcO9c42EGkPGZP+02N
dfebIDxgqLn23CT6mW6XLcsIuQQOmuV1ugw0IwPvjs8pf8jL93k+G+LnFKWNnFMU
VmD4uFb+I/DYKLryJjFxj26YhWLtPEFPFNoawCQmFu/+BQrqOWr+Am2rV3eXSTVy
NHXfaN41DlcGQewMTq1Wz9cM3D6bE4Krvdyl4CJ3/A4M5dJClCPgMFEAeZI02gKE
xsI0N5JdHkXebSsFl/LnDlm6atwIMnfd4mxPrV56f66NDxBs7BTHVEPp5VT+QTdr
pqR1LtM0ff+0VMFf21w4ksj9kZkuCJkRig/yUmVT/Agb+Zz0uQHEIHgWap6m7B+f
tW1cJZJTFMdZHFb+T/V4L2t6qkkiYxW/8TfiNgfoPz4KJQvhH0yKyFSqI+qiI0xs
4RGl2QVus3rZgPWC+N9sA8u8LJrN+OatT1PAuCyq1Hoxir5Qfv1W+1K0VMIOTXiZ
RMnrYJPx9B+h34e8mNHcdNEyV4ZY0spEigiwitJuOE0eQxN/B3VRQkM3XO1tax/I
AJmN5ZZxm5R22wqnQ4DJxtTbamwFrAtwbXTtIxb9t5pUB9/br5dZuSr/NDkyiqsJ
RWQT7MkfoMnFrqsz7zaveFZXjD51ipxwVxDL5WqwwK72p5b/FgoUHT8RnMCEQDq9
4C90Wl9ju06ITl3JkHB6tWLYJuD9OcqDS+/1UBSy7aePfq87bSNYn7DKt72wBZnU
SzJEBAT7nqh/MPpOOozL9+hbKCn5fDgEivL9IPeBH24wL4lXCG7REFBQGBCtaIjg
6LwKPf7GKU2TNsY6EPRlhpDAd7tMvsqPU5PMbw7hsKae4V2eOBeBLb4e6wdfSa1R
GOihS0hhDMP+gXd267DyBMOdi58IgsiAms+fS02M4mu/U/lONTX7OcLmiIQRfa0d
pQEghlXrQIk9WSAo+Uh05XBGKM/70/ThuddCRX/2YPpnxcuNcGtX8X+8Fz7Y4Ja2
hNFJwrlUzxTzx01FMRi4AePQRrntNyZdR7h8Bp1yIYRItNhacZ/Kud6KVuQkfOw9
vgpow2CuAvoOQUqOBMaUo9ZKM4wAlTqIXKdqm/7Anye0kfLsXqtxIhE1tNxWxWDx
Io5TbU9Ul1XxY5P8VcS+nd8ryIR1uWWskH++/OwP5iVVFFMZ37k651oI37k6CtzA
jtuBgx+B4y5o/7if5tvn/eBds6lwI8ckgTm3dXBfblwXuEiEVMNNRZIPfCdcV2o8
ghyI/lwyavUQSM3Vxmw3iS+UzFTdACYDwPrhLnkKMEP0ht4wcTDb23KyVru4WuGS
QDnfBRvJFCgVKTjAjUV7vqxdMXb8LsWKCZvOm7rGABv7AtRp8os4Y8tUcgHGrB+r
0F9zcTjgpi7itstGn1SL95Ah9GGMxJfEaAOo15Y5biJ4neHEuUudTxnKT4N87zax
sO+1G9hxmxVdgwjllspMJDzjZAvSieBEnnlGSj8OPJKM2pz2As6ryY1P1o6BEgUy
kjeoMjZC9/IJimEZz8vdJLbLYoMzUo8h2k4zE3WfpD+7VLNlE+aTiwYb9hk6qLvP
+AjV/RzCssQbeDR4kOZqRlmDj1dbdv692VAgOO29QR+P41WjHE1jOG7W+Ea3ZcN2
WYXFa2j1fsX2thBd6Pf92Yo6nlGHI8JEHAKwMAOfH9kOHNxVqfK61/cJfaBQ37vX
r2NzgOVpHRi9U/xzPt/TLdI1mbTwzqFe4QiXu+Jjc//8N1VGtgPMxwLlHd4WZNJt
hP+bEB4TWrqxdYz7H8N9rCL2JO8IsOGK7p3iDbLbyYx5/bq3Sqs7UQWiA6+viz/q
gzA0+PztVlb6CorUV1URd6ef54l0Rtd2oqFSZqXasNBexsJBnrbWq76rensr5WDm
LtMhvAqjRMWxwE5PIneZxR1yt2bfDNxPOi0fBgezutarg9Atgr3TA7NtTcoqiHBk
3jfE78iwn3lz4ZdABRwTOWLtuA+NAvJv+oW2FWbnijkHClg0v+tijgtokHAcPYdr
oaUFETDPZ17xpbX6zYVFtpVHj7fFALuwR2k2FnjVKCK3G0rwbMWQyfwRXU8vyYAr
0J6Z6PF74JPF/HpzP8Cnxo8U5p1bm3yythNLQhrmu8x210wcTNuWrYI/xgaq7YYP
VLRxc2hcobKByEkjKoqqTDlpg1f936pdLv7WCPzq1NnMu5ZA+r9/zAigbS52rZ3N
N2QuhHWK/fFNlWc6ekJ121VMh6KiT/niss9gnRQKKxIpmKQU38KguJZtmVnAd52b
9rweVUnpfaXoxlYfiAAX/jwmQm2gTatRXV8MPShonzepinikyHaVNBZMbGrixzOm
Nukaw5AsX8x9kUdp9oILM4nKyL+N/25FZxgA8ut59magOyAkERmjyu8ePlBtDwlg
bNwwmBX+mpv3+XbsKSGNoWk77Zn97zXj/pYokrmbFBQJnQNQJ5vQ8i+UBg3Z+iZU
s97J6uOqlyJ/76JL1+dfRnTG4u168Fszwb/8ldpwhIZt45iW/vOm9IeMCr8s2+bF
CeA+xj/Fzjzq7i/1E+XsudOSz5MGcUshgH/fi6Y93LoYPDBfGm4+XVNAiioosEwQ
6pdZwDZLKVEm+fOm/bcV4dcyU2iBoZ92JiiuUy+uMg0Ny76dBiQWrvIRl1SIpHQb
2qD7/1/JhQ0MkZVQrlcLfKY0vxrEej35gnSVrx1cRWsPEyvur48G25PdMJvio+sh
rsKmypQPNZCz8qd3jsF37uMwBbnugeFm82OocIrWxpAxSq5ZUH2zVMztd6HKBX06
F1A7elKDQbOD0iRvkE4UBKiB2h1j+XylJSMi+MC8qN3Fy3eDOQ46kjZSdIQSyxh1
tDZWGWX+T3EKFkERP0DYCKIeNOtdpaSCiaUDmDUpszSUy9qvwTMYYLc8uiedp/wQ
8faCAHDR2rMFPsdujgdPL/zZXzChDIU3E2uJ+X+rNU1DaI4Jd3QcHNk/IRA3Lmd/
o/QAONU8ouMZODYtGZWElYK+e7+F/myKIYycSyCxSwOJukjWJJxPJ565TcAtTnUo
apIziIiQFogJePUEI4ESdXcP/Shi02L2IfgeI8E222ee+NT5ToWVd7cDz18mSjin
IB3z1hiP31JkXra0qk5W+KR3hx8wY+kA2VehMP3xKtCW+zapbQQSnifjWL3lPjy+
lFXz9xium9GfOopO9MPj9bS/hoH7m6qhZzvtWzy9APjTbRLbTr3l2t+dXHyF+Lxs
aj2SknP4UUhSjUFg5NWon28stAeHoU+OZfxZNGtikEy521KNOkB0tQqfKYj97w0N
veywXCk0C5LaBzqX88b7Ae3aXuOvcOHHdpx/HfavnOM1Qsm3cUeFSP8piHYNxUcs
k5AGzQ9fcUXieyQZQYGdqx5CSnQ7GcGKTRL3o88mQkHuRiM18sWgugFth5bVflNw
/qJ4q1J2pHwNDfGCEXurR4rU9YRWcGGg1wJn50gdzDs2uLsW6rVP/9hm8vcouJIz
zg68coYrQ3h7cEuBNVLqF9osXnNfGvaXUJh9x2h75Qn4asVduNpgl62iS6AWYl8V
lvyRpIfG2PkDIiX5eUiITwtqE6njVRXLtqX6HhdTjURw4sqGZkvHh4YNAPPVQOQK
1ReRT+vmERqUQRbpXFEp7J4HfBxJjsD7rRhFLlWJ6wt0r5NkTbbHSof6D7UV58et
3Yrldpf0KdA9rlt7AhHOvKHURtBHDbcoK1TfTHp/UzIWrBKIkFY5vB1quTlKS4gO
5wSVHXlwrIylGudjruWwE9FJzCgOJf6PHCSP+9SeFItsm2FxrNqRFkKg2U1pCeSk
MamrMcaryazHhvLenfodmYvcF1XHfld43nFHYM2bi3f+fwnEggqqOAMKgyooRjDM
uzE7z8vDTDitl6nLRO6gSpGE+hC2F5p4j5uh5FvW+xqVcwfmcsLSI06ocAgnQ1OU
vg7Lt/rp2dIPKApa/4bghh8GDCWujo3jPWOaxeORc14HDCdiLWxidqU2IMBL7jqN
qb9GQVlW68z/w/t3f0bcPQDaMPoEdCm9CbcDbtvYnDmAuAP4ErSDJ8nw+Sfiat9w
AkT66+GyFLEJMx+D3EVKSoBVEJME1rU1N25dpqVhQ5VTeuQ+lLqWabl8M75fdw5V
352AkpdiKiJcCBo+gdV55Wigf0V8UMsPe31vyyyYzRcGiCc98+A0JrkeIAOZ7Hpq
jX540b3FhP5W9sQ5SpbSxPBLU5TydeEXwZtSByf2uJtLMY8Rfkxa7+b9Xyo9A855
8XPOrFE5sBGeoBFU3DaWKdhJbeQi1WsCUrmeByR4rq383YXdKwlPsOr8tCjd6lq8
O7mR/VcXMTxyQ6uau5Z69mqyWzekp367/52kB7lTzyvDiWutqEVcfAaQd8n8k+A5
/DrP39Qgo8WaJdKdjg3blefKA8FYG4Eo7Epnt6wBy8OUJviZ3WsZKQI5UAosG1Tz
P5U9yJtxeTan7rA7iaWhskrtjbf9Q1MoG7/JKlwo3nxvxaKfjx6+j6LAh4lbtt23
/4d6rtt7LpQj3CUWMgVY2x2qN+DSs/Hebd5hAwJ7NfCcE1J16ZBIK2dN6/7bvibc
buE6sHBc6Tuk3ej/WDaRNfgb+xN3DoVNDtBu5s9r6C+6Dz9FMhCyO8+WW7o9eGjv
p3Q/0b/oMaKwmeKTBpuiIXBdI7pHkZOsgKch94zsKJT8sCqKyG/Iu8kGk+rmSTlp
9wigBSSYNDENXcD35l/XI+6KPDRC8FUte2JDEkn8oeaHRNOuhhxS7VER7z3pe83B
AMiKMW6aN+6S17J03CEcZfetsISI8XWw8Oh7q/0bzyPhmlC7s/Wo0LwkK9GGfRc1
3gYK+ZU4xq7zS6gYQDE+ZKhHL8YC1UhxQCXLuV2/nJ3HTb+s/jW32w4Kxrhdcqnk
Ri6FSdJ8xg+W8BuJxHSgsMiuf4IoqlMRQvXVn2WKnI6ITKn9RSVwD9DXXjDYPv2Z
3b6XaF1DG/oB5gsUqEy15t4uabJeU5onxh0XbDy+6fxHLbImwkE6DyWiAqa/e7vd
2BwIYvnHtDS2l5RVo6JipHjCXxJ0rblc9eTE/d4vaJ0pj35oZtdO7EZxt5YIR6we
REKDYDh/9T7SgfMTKRjikgFv4AYG6t5ZxQIpWaQvMSqI4+Q2c+wewHO4RBsnMWa1
ujSb7flBu5rVFyDHib6tkhYbmV7l5OUG4z24Aoj9EZrQVjXZHiZSUVe/u5n6EV+X
E9A5rOrhpdO0aih3No13Ar+dALHFdUjccbc1FOvsVGU9tiUToAoJ4bePwfr4v0wA
5HP8SFXOXxL0x3fbN2a6HTp5sPVA5qerXaqXjugWCG8FKgYjCKQs5FvvZam3jRNo
AQwi53W025xq//EzD+nnEPTfIqVi+SDEEPNvT8kc9GYt86FrQSKbqLDXDG5DeN1m
5CWCK8TxTWW6kRWqOVnKmkUIECoJth3YwHXrQy9+mI0MfTFSdT/LYLanjwwQ0uv2
4wR3o4YfbRoRhLLGk3BcfN69QN9kze7lK0xGfCoeZhvQdnjMvGLuYEgYFurfNR4R
s91IQcDoc2a2ACaSjS+tchNLpW02uTrK9BpM5wVYYOZ68wWEKRDTW8cxr79xDe/9
pdaQ/ooQ5kpBYp5Ml3h0mZpWnPN2bpLNfsxbuBFTM26v/ipO6U1D65QlYlJKK6ma
CosyUswJEVBFRdWKVhM4OczynP/sbF1dkDF/nCrRYEcSBSUJjHN5VjzWmrFt0Rkw
jnzG9G0Atr2xx+oTXSyKDYhCXUuoG8U8fOuHFEf8z3gOjCq+1wMd7M+O6CNXGwDA
TOqNq/BYXpqXSqXeyOU1I2pubnVz4lvJ3OJn+5W1o0RVVemoTWyYd2A+s903zyxU
YszQsuVfu0Tg2neK8KIhC6/Wqpv58c0fv9NTkxI73bd/WQdnb9PTTVUuMolQE20q
WszHnTllbfBnjUaYlGR8oLo5H9awp90TImKhIFEAOsmHW+JABCsHV1jRSYGfXQ3s
4s+Ac5JaM178fZxa73CMVkABOHF83A4yvRBmp2s/yv3iPbMvF3M2utAhT3N6QJHh
fMYZG2k3j3OZP5NoTfq3in2NnI/csSI5NX3I/ndhimz0yo72IIzG66U/QMe4LM4b
jD/NNoJJtgweeHDBqPPHDcxbACmN96LhdP7b/I/n6TLHAQE/Ywjbx2QLJzVemucv
Z4bNsBjFAevlQMQs1ZEOWcV9dQbOCdXdDGyFM9fFs3lqTQguomTo1LvaMHqRSVXv
vFviCOeEZXNcD6wEIC9LuVHtm7bZDlA7TM0i2TOr9LSI6zXYive7/q9xixJpYlj/
gKdZwTIdZfqBUGHyrvBUXFUHqf7q1tq2skt8xK3+6jrgGW21P28ynOskgZH1srFw
UbnYu//HWNMRBKgq0SHm3D8/n87EzVDf+UjdIiiha1WtPZfkTXK0uuql5+d8ylSM
+4nrZty16e/95uMMOi6zyniUcrHjygHFBh95VPqFEDraQC2CQiz+rLVgf0ZEXGR9
rFbc/bBr9jw0OnfPaHOjt4S2q2wd358a9IiN/NwR/PsYjjNfduCv6y6eButGXvXW
/hxikDusZj1agzTR5CT/ce+cIm3PVCegFBeOjOl6J1A+CUlM2PxrV1qWkvoU9Asp
g3vlyTjxAEYT43e/FHXUkHt9WbQteX/JHB24z2nK3Hqp6mjerDCnfxw+cYsvczHU
16MLZJW09A844dIfH9KXMrbYQ/TwyOdyEeAnB4bJ6KM2OFd+axWS5tNxRSAKb6J8
GqymbonCuBLaSqIkVHyqLLyCulKibi2Ekz5AG5h9p9ErUkcuqHQgJBpjYSMuYsPF
niyu5Son1fAMPpv1vxd+VVP5hM0ZrNP4YPHAg/jsN5g0SycKw5lT9A5sheCP7bWd
40kKfSorpFxtuN1JufPiXLi2ezURT4IPLJd1ofb2vDwf5ows2DoXwR4u4GSlOD/T
95mnbD/jYOAFLWVplz9GkgNN6M10SPgV9F+JXF04X2WIXn3TedFeqQf8UHwdFgtY
wrRaJQL0cd6LUoc8bTw7AvgD+MDM6tq5IojzRo5p7zSWLLElYThH5O2KiS4Mi0NA
FlCIloyUFx33g/2Oj5iqJ59Vdaz19NfQJn3f3Ufsr84qUX1Le21piN7tT4ZOFSfh
/Q6HXuZV+rUP6P/NdB0ui7nLLel0OfPbkZopOEJWbxiuVB3WiMIp03WsxQQSpBmj
L4Z276w+2LG1esxgLoeWbL1cW859PrC/koH/9uyWg/BpEIKwnQcEdg6rA3YjSnG2
6nfX00I80oyTs3mZDAby/e6NNiiAnFLV6dWcViAbT1v0208YvnmHevs7S7VP+ELE
QTXiEzvxjMd2F7iMJzvtMs5UbS+VTCXreqRnYSAL/eNEaAeXvkqtmNaonA3BWYsf
6vT6aKrSNqruPIibFO3m/s4FwCfP8goQ9bRXec0FV76rGcxtm4NH285dmmWKzbn2
CJ0+pVmR1fUbPVwtHsM1hRU20x3q8vxh8X86Y1wpNb4rKZkA4YYlOgsUno6LFU1Q
pDg3FytbecPOtu6wGj2FkACddyncr5pkpgQu7KIvpliuDsVDKVw3im5LhPJWfpT7
848vx68QIiBVC+1MbjHUzWU84s+vs5eAdr0dtNQHMirjcVBrZc0V3COKRBVJcxPP
Ig+6p2VJ2h8qdkxj84+Dq8xPGJsShdYZX011PUa8u19ZVvyg7NaNIKLjdg8VeeI7
h6CYfdeVK5Op8KGP02xy0swK7EysoTjW6d4UP4F43thnbv50nKhJWSTofpKx3ACa
RTLlXr4Nht/m0srUSwF85K0NC/jlUuxkiwNl6aApNe09jxJwvWOxGjwjY6mycmQJ
dxWXcP1bN8BD+Cj8aaupmzTq8MO2G1Mf+DTMC/FjfRG+pTlg0E9zjyD6yvhnx1Hn
QfEEJiGMqZ7U9zSXW8eJ/6uii6Kp8JGMMRaKjXaZUTaRMf1wJdSFgzaD1XVfJ8A/
S9furcKluedx919na5Kx6PHBe8/XocNIVoqm8cWU4GVQN4Qek3NAXDSjR0WwSTah
47/VUP1UJSQSlY8J2fmdG20wW69CUODxDzUXDCQYO31AFn7z91QyUEX+zaJr4eqG
yrrsNz/l8wFWdCv06TZz8kmipL1eXJopdKL9L54P8NnE0tWQhJEimKvubxCxaZaf
4y3JPLpjeaRzOfW4N3hbOMP07hbH4+3SDj+3tLVnn1zkQWev+aYRdgK7GW7uMBk5
Qrhc8Fs0n9sxsmv0EQDIjPblt4Y7nPYEMbiJeyF9Ps/ARwco3NPuHzQs9RFVeDOy
FIxi0davpAw675Rqkq4/Nhaq1v0S4tBNhmTbRhGq/PJW3hUxWej66ARTdj4a+ahM
bz4r9bPDSVJGf2Dw70QlyegLBqHjPUfQ/rxaZNUetVnuIpiMI0f3wWgTvocm7ZqV
iqHzX6Va1yLzGhEVdU3RXSFvt0qrjVHr4mOX3uMsJYNdSmXzoGrc2t16rQ5Pw+3U
v6M3b885H761rfp3Q2azVxZtLHRhrmk7KKIpfifwJaQnzgs3G5WJ6t76RyHkSs6H
+aSS3XFR67B3GVsrKCuTxlvG8YYRPq3rRrYQCuHquXsPmukDi2WQSYHyXZZ0P+YQ
Wk+YjslxsuWhTt24BnTvRFhP56PKzb0r6kFFpqTzy50Wn89ma0njRDPD7pgzlxqx
m6uBRgV6xM+ILf+7EzI4S1YWeIiAPGAdSNm6EWnAeRzGEo6doHW2n+vXYNUva2vo
30rk9+ujxq/B9JVzIekkmCqrC2mfyU/jnac5XcnVejXD/9RY4wF6f0Y8TudNdl6k
hJs2E/9QNaKi+4x83+oPeHIeSoFRTxVWPYmx5GMeAogP1Racc13ZO9qYWNWqFnFH
oKqy0iUFpBwa5m+dz5rPg9FHkqQBX0na+jdzLUVW0p+9AGAzNWM69FC/Ho3Kfics
38nT1tPSiWveOsVdqkNTl7TyhMDnE4RyVk28+maXNWa5RqgqmXxXeWmm8Wya97Vs
LJlX/kcwmV+TmjxkPacipqeQq83svnVe+3ypD4WcP6qRre80Vvl4dRlX9ylPkm8a
hW2Oo9CyKsTKMOoOhL6CSjbOOVT0nE5lMsWac09UkTd+vErxBvTs5c4iUnHx4aPq
PhJK4x+xP2WSHCZ+v28wRaaUFP65XhqmMpH3Z7pmf5M29Y4c93BGK7b5+1ktDhnS
FhHdIkm2cDXzyHhFDajr1lE/u3XyLtk9likyDNrmUekDktHRV2eyEIQbXxntUGr2
bbzw2m20MmQQ/PxjSg3gqlZC5WaqzwU7jb25Gzzu1eiB5DH+bjQ/tTL/u99kwL+q
Z4dO6aBQ0BCnkxoeQ/i5W87BEFAM3Q1aDb1W7C07uosx5tLrTLvYO3iyv2rnpLNF
U17GZo7y398hKlt/kpE6DC0AeAQtEjNrgZ8Mb4yARkqzkOsCfqC9rW/5XpoOFQ0E
X2vWu2a+yH3o+XGTqc/xAvxvI5qIjKtMJsQHOdDaYte6805NYHcaEQWtVWKm/EK5
gGRH+l5xrELcAI9eg0FJgN+QF28C8x/vujw+YXtzCAMAqSDrfEVhgKndIfnoh6y+
1oorECyc5nywuC8LBTMM19/4waQTKqDiL85oVB2OgmHlnPULbhYTKSJi0IPJQ8xE
+tYLiORtRtfph1bV15j2BcT+0BH78jnRPF1sY8nEQ2Wx2YtFTifEb+H3rnSpusVp
vYSjnWj39W2H9zZcWRRabmAVEggUEpQhfXksFci7E+IusNW4UocfJcYvCsB5XHi2
2WILa3UhUPD68VmWTPxcNcBZXHTJyRDIGfpAWdhheDekyFpY812wQOgwwyiYs+md
XI8REkZBxaIJA17mI1P3bAmZf1TOX2PyokmkNf+2x/AoP78OrQ/j6WCS66mrYJRo
r5IXEUTyuuKz1/jMBPa/DEOv/vMs9XkAqkEitn93kh3DYqKOIR2koMpdoOGELEIr
968ZRk27UjZaf0lh+Ps0eY2n9olqrwXdqyxAgp51P2/nia6/CFLoTTcDQce/Td0d
D38DqV+3+2AdzudpGRg7HuttVEh3G7E9E6O8d8XpftmltrLFX7EaLldXrDMeKfXi
wZSVeOmM0gDT4nkqENQdOoV41pSxHD/a/MkYTNSANskyeG2PnjdS19e5C9m0NpNj
U+nROp7UNaHHQZve0cmHjIyp1Xv4IbZ3bYrKMcRlCE5o3Vjd0er76pl92h5TIVQy
rUDsehsUumoro2iUTdLBL8ht8fYRIwmNaxBvH1jlLM1woMUXE14pTrpbT3ZiqsB4
E+02ngLRdxMFqc3YY+tVA7RtoLCTJ+1u3+Bua6mODPDi+rCJzXajZv1oiXwH1Xuy
70Zny7H8FPgpTgsY2Mr0Csq5MPd3KkzKYh3hqaMwYTRy5naKv8n3VbbG4mw5rKYO
xrrvVC4eajy7tdvBDH1w/OdOx3L2yONIos+5Amke75SHZkML4gBEXWXIFZlGnCLl
8tQCLch8CwneD8zM00jlahO3yf25TH68wmsVM6l6r+OIGc1oHs64RaH+B1gc7xO2
+y6HCkP7X6ZBTayVUtgaFcaLqVyoXgn7BWSWXQKJ9f0Khnc+1f+whB8FY7KFoHln
gJaMB4UrHBXXJbNjiFQNv41W6hmNxBMBPYnKlq+61yr4UyFec6zi9QX97tY+1kGm
f/NhbdZ9gAE/cWMrzIJJ4jEF0MY/nQoYZQfH+V/ZUNkscYBj5Imis4SGPwP+jeFx
hcyWNW6YdCRd9eEVnkuK81YO13RJanCvbvNoB6wPtx+K3OajlhVSu9gQsmoMUuBm
CV4zvjNfoqh/2vKwAjzgXn6O9eBOiyHRJNdQuLhbL0jpbYINNvsudWZT+fZr/EcI
ZoFjXJPNUU7mMMn7TuO1vRAssxZ/cW1EHS80rRcQEaOuoKWNInwqKUjUaLMUbvIG
oEhr3UaWb73R/MmMEQHAJNtzOw6fv6Hir0X/5rt2j8CS0Sv7i/crxZo+bfVDTWzz
H9Psh6tWYwZjkkId4TRk4+xxTEVZIhy7o3ZcRdPnDi82WiniCCVeyak5YeH153O2
gfRCH0/k2UPdcJiM0VQHKNcMw0njMr+gfUwl7TIoemcWU1p48tVgLgZVzzFvnFmF
rc55m8WSzJYlId0kPH+uNRAW4LHhg4gxOZMx+mYSmChBieyfmETeyuL17JiupaTs
HRcCpe4Zq08yPuev9CBLda20iA4nj77dPSvkp3Fyst+U+/x5wPOsK5VxpIFc/l7/
l5YSP6mQ07nuepYB4RwUotaafAzvCoYrSMJBHPNqdPhXTVjzXMM3q3zESg1se/0P
LDrc7srEuMluU9ecbMjo/O6t7yJ091HXABpMYMU9c4Tl2STiCfm5t7AgSCq9R7i+
e/QWzeBthHLcyG5MHnOJDI34ajrz2s4RadI2tDUlQt0Teb+fd0dT3YZWAgk/B5oe
qBV+ZWi8wxlFzBYxjWWqSMV5IwXnPC9oEYFiH9OaxGT2cuo6bMn51Th0P+/KyPci
StTtEH15s/33FlAep+/lwRCAgBmlUJAzzU7usoYn8DxGyRenTcpIPzVgsQU5ByAm
IkqVZh5vx9/gzmTlC3SWQdKePvMVKxXFyPVxUKO7jQ5V7ZHrfGP5UyGZ7NYa/HDD
z32Y81kPzqDSJbsnDZZCvnLq4LbhiIVeXE79vrbuHGXsfGGNB+jh1IAsDzLhiYyS
B7oeTkhmqp7oXAVGfm2tbmhDOk3nxQanOTJehajXw5OunDf9c4YC79UDQG/B4xT3
RY/JytgGYF+6g1TkO5hjziFcZP9H13ZH9hu1BQ3+BjEHlg8/p45bIk3KQkS2PLku
9vFMxCg6SAKgWNOQnxR92YJRQhyHxIIfk/HF1zQ6Orfjo8QyVcVtEuMyPWnJpqn8
dwkitGy6WSCYvYIs+xvepdbEr+3Fd/hwHwlwL+BK+b6PKKZVTpZu6JuUZK+6khQw
jg72t524O3eqYVJRgcbZafEo57MM5c4rke8QSLiG2piOeTANfiKxUKHn+PdKckOy
QUtOM6aaWoLwE0xHNo9QSMtQ6VEQVJ2d3R9BvVvBuzG+g6/RqNjofKJTdjV7KilB
JqdOSxZNRjjoRYtQAZEzvYtQXynkkBkEyr/hnipHA/7UNneEvsfGDtTeIFy9mo7h
pGTxaUsYUl2bNYgyuF49yPHZEPcWsEUxiW9yTKHR1Huz06nBcKYLHNU/c+FCuZmx
0DCusFrQZ4I2DP4l3qIai2ocTPtTiy9IxLVpjgqRjU/fVGszjG9t+fMD+mmbbA0A
Xw9u88PM1ILd5gStbuW9oHO1CBIGzTemnUzD6XQkEZdgZpjpONQ2KtE8IDjwYHN3
fyPmOrifzWt8qZCmekNT2gXjikuerMTTf+6PB2YxSGRowu78Y2tJb9LWmF7IyjOR
wyPqoy/opuTV8lJwHjnzgpQJsoGwocGRQGXneuBIG1gcZxZ/zMCb6KCm2yjAdNLH
uZ1hsvEMMsbSK0ZVX3UTjbs/d8qzZ3mQDAc4Ci04hvj32qS/3FPSONIxk4Ychdjo
mzdlQ8uQ9y4KRyCa12spZoSUIluhLwRnBLLEPgVgely8Khjw57S61WwTIghdh3tf
kocMijyAZd4SrgflPVUwukG900BJAXdQFGKhQluCPtEnelaHhxF8cYzgHD+Eit/u
1TIeGN1i1tDvu40h3LRsSLRV68dhyIrRArkvW854iZKe6NLHToNjDBjzP+6nCZ97
XES/d2El9tDa9Vn8rgV4L77YpurnsPJ7q+bdOF5e8phTwK0CML3k9IQRHoPpzAOZ
Tj9SP5lGkNwDlZTYUpa1UC0zuiQhXvTVTUCZJgdyxTu/oQZhIZ6m7H7bqlt4UlME
BFs1vAEvQkjl/YJ0DL5nLXySRY23VHm1FCYJPt0757HTtBtlCON0H8Vix9J+vkVO
1A/9Vx/Z45xOULEK/F4Bue3pB2kIwTly9gKKPpoNqf0QzJxSJkoGx/DQN4vma/kP
OXAn14gNbb/2+MdzmOI3+jvL8y11r6IWvbXOPaBem8GR4MPY+RYmwb46zIHAHcHQ
9S8Jynk/mH4GjZLabIgK+KhlzZVxhNLJzOO2wHmBMba7lKxKZabfLuKu4Uc2uHcU
yRUdI6oCu8hSycaitxsvIzv60prd/LU+9bu8Zn4ZfupJ/7yXZ88Jf3BAH1xW5cgW
0nhXFv+MAd6I3jEqtp4hXspa0wPNn4k+/UGmp8MBA8dTGrbJRMstH1v5owydTioC
9vj8550W++FDtYxoa74OaVD423xXv8in9RZ2ctPsWDR07lj3408K6rmGpO5CWZ2x
02zAd+5qUWCyXbf8zUdHzGM80GDHkvh1gKa9ZD9/styckGd+WcVISRhPaDhC3VI2
inC0OSTJatIYEgTadxjIYLOLuX8RsvAK4ApzVZLgY33BssWLOl44iHdCXih476X9
kuUjRNe9cCPjZmS3BTBJJCn0eLBi/ynoNcIrRCNSGDK1dnpXlTmDRxmyY75tCaPW
OCjPX+tyfenQo8fsKvntCmcW1hRbx0y9YxepD74G+uFbCfBtfzaO5oS5ey1nXOeS
rKkKQkd5ZCk66d56bEtXAvp8fgDf6FPaanOHwubnKvx3bodGsCcodPKJ8zwc2wHm
VNxuJRzjxiaxeID1eab7x5gNwdvG/p4DNb5d0lTMkRcg02qmIf7o6x+nRdFvLG2u
Ac0IS+f5h1aQOXXwUw00yDDYTJzIZEVZUKAuFz4CQmvPEccWBJkFfYp2ShcYIlXj
1YQ79eL+4zAD4kM4k4Ux/hlvldUn+S3dg81WsRzNOtR75RuoE978UJSQGjVC7N5P
K0JQovcAvumDaMbYXscvE0jE5Pus105KwsVKJRLDW4WC0Lssr+qpnciBfEC2TW6Q
X9AScMrGvyM/c47fAUhwAe/czSiiEErTK8EO+hXKRi7egMixzYW/+Bnfh6QSgGQ7
xhGClJsTzHZQOrhnnQQFvKHosDs6xQkxlyOdtYH2V7qTLMH3qk2GsCz4BkcNRFwf
iuLctBvVqmvwt6txLnT/wn6ycg/m8TYjmFiHhrrYXfyEGNoai8AZArAAU0M0fOOM
fxQcJ+pQfaJ2INLlhB0Tz/SuYjde9zPISEhFyDv9K5v696rADtmhysYsL6hOQaHp
gkQShADcxgAxMNPkVtU0aR8TirP4tw9oL+PnPhr6fdrk7xzqypW1DH5pESpPnEMg
Ozc4bSazh3wtcqJif/aRro9myth29ZC9hktsYeEgOaqe5rTlz+CI7ApAwwWNQxjw
33SBAFN4hr88cINCOxnsh5h2x5r4WKfKBM5HWqsR0n+S0gIOl4067Z9yRKGWIYT+
U5MYtdxmmywPxJryLOe4YTnUjX4c0+XOs7dZv5QYwb0RVz5I0HgAWuFIddsOPyf6
E1wRv26VHUsSgxJIZuu5p1umKaKwHUfPzVVUZjdOPHYEAYM89gI0ReWO7jdx0T9j
s2CtleiWtVAWcnJBxj9RSbANnvOIy6Tu5LNmhlei+A6PVGVRjoLDofQnQ/tgEZnt
xjkLAipBfliTlaCXi2m8ev/XIogE869cpt7FEsH5+FREie/HHGVUvTFsxAHiwRza
njaP5rfGPLc/naHAQfbg4nIyOQ3w23XESlGXkecghNqaJf6SZCUhUDOlNnRSfYTg
nuOIm1J9CnM0oDaZ5TAZTyvFKoZnw82CmElivvxw4Tdd77HpJzOAUp+zsbeIXJbm
Z5YZJTcLngKM4ZCbtvvrudqXKh7wvfCXntdduQuf9X6HU9sJu8q84cCBJN8mNGAH
gwW1jkQW8vTiIljDiHEjXYumZ1aEm17erULqVEgYqfrhUdlPW/l2WFYRXepsuUdy
B0l6/CuwIeGPI3VNQryylndMvZwcJ5ybKU0Ge0pFn1smNlqEFFDYc5VOnXyRevhS
f6WdaYdUFfKiwHeI4ijiveQ30Ewdbwt7PN+MT8/xmhkudGYHXzw7e9eXF+PJzR8Y
bz6aR26gEmTD8TzV7mGKW1Ln/JLcocdoSjPa70wjGycRcNwsyHIzLKYEbgFdz6zC
54lf1oAAKxf76IRdR8h/TyzcBLXgwNU4oHZKAswGlodW7xOwnuiCvLgr0yHlKR5C
8BunkqmOhQDt/f2U+7lmcjRMQu4nlunYCmLhRGoxrYz9hZun+rNRA6k+O932yI3Z
tWOAcpx26PtpfH2/CAEiDua7G2Buw5rVwfd276po2Rgj6elJP3USV1grFtCrrN04
C++HmsdyZny/ukYBl1dYrOtj0mFfjwnUr2t1JbHbpTQG/t+F9mwp+VTovx24o6Hi
da/RkHTQmjkpZ5fhZTBchWXRtSaC0BOI+eFeDSrv0orXy7kT1eAF7LB552R4XiFB
31fgM9R4chmk1dGt9p3UyjvxbDIgMU7U7HDM/h+hGdlDaBzWYAjQqPOeL5RDeOmW
RWKLWdXBJO/xCWEM2PITAPosfefAWqKwE0s7TQv94t17tcyPfqY2VjvS/bwQSLm2
97l5Q/CIOnLYNNe88hAoq6BXWS8uTGnaP3EN7V9eVQwbiFwFruYTJWtDk9bhNlAm
uPeP6F5bve4chDFaZ2EU+Fy++zufMEXBKYt3bSJ/YOL1b5RUW0F8ATnNYveJOPS+
N05q0k1O6otKET3BC3RaXca/Xhx08jnYTeglbKiVztOl/oxti0mYB9SryCV5skqc
iRWodqkRdYwB/HU61gfhoXucvm+viHmYS2thRnAZrhkZyxFKOxOIkJqZdfwTw6ft
/uSdUBbjAICZpMZ5/OD5cckRuA3oeS+5e+DYvBUhu3cHUCx1LhCIIlJbiwTjZqKn
uTA9alR5z1ydLlLr+T+BlZJ+4aPkKXyBIjIfpx7QRmeKd+9M/iOMy9CvVydG0EaF
gkulVWwNc4n9rSkgpPv7WMls2UL9k5o1EuktXyPsQVHLOagcw+SVTlhuhxcXAve/
KEr2WwVu6ejK0sH1JGsFldpHV2Dk1tig9WpkTgikw4/EiXD1TofS58EBE275iDnh
ZBiYH1xPjnLO6qLIleQv/CckT2q9QbhS9tNsfyass2ZhlNQEKZyA4YdZN5wCwZgX
MGvWujWVHYfW/awF+g0JOL2Tk8R1vlAjSZs0D3j/kSNwOYsA4G4YW9OCGB2oV0cp
Kuc2plzzr7ELr1czwSQd2txTZV/MNZv24CG2hMzz4DCY1CeTRURQQkA6R1Fy7MwX
Q/Aedqgu/MqDt8kwOXnTwSS9cHGMCaah86Z+gvX/+OPbMAF92aTgUSytmRtW6Hji
/fcxHhO6FL427pxW1DqYdy//WKNgiC4ixIiYZO0UEBXjggiXG4l+yIOGp0Su7TsO
bzrrZl4yTNqLSCPvHpn7CpZZhNG1NzR5d39oO9E1GQeip2ui9+FbBKyi0ZBrczi5
OQpFkaB4vm0SzUjjRgtHo4eIlIu6C6U7d7yU4VMe0ZcQ4jMDnMy+371Q1VOM6x1M
Fen+XZ1uYvGIUuC+V2HYh64417gcDhW3kPa1HF4RJgTjLToKn8CAZZiZTG1NMdlb
EFbO5pF314rW6eliGUKySBUXGsesAWgpy0zNtWFxVHNTAdv5iVZPs/OHIAG9rFU2
7+zcozek1cSF5RpqYYsXoSTIQjUI7ioEDNVAPPIbhpfi+f3jXaOBgEfgW3xvqeIT
4HK8ry9WT16t4I+Fz04UcHw5U29Z47UFp2CxW0sD4V/NEMVVxz5NIm8s8HQnWvWS
GkBpq8aSXgeNtZim0uX08iD/QDKsduqTGu8dfxyP7aN5Iso2mFqO2/z9QO+6XDzV
tiuwyiwpCSRR811cGi7+EeJg1B/Y+D6PDSlLg1m6cOzt+NgqkszsBMI9jo4gEKgV
OPnHH0qtZMOfCZF71ksiaOEqVWJYFH91BqabvN6R7TH67RteIcEazeOjxYOEyUlq
VOUZSFHC4dUaPdsE+36dzDzPJWkE/vtLKm7D6wXrn3l95LfRDbKfetxUvd7EnnSo
3Fe2uCqt9qoYZ6ABY6AL3D77MKmqGe91AWNRSiYo29UH4I5WMVx8aHqyHM9G3CY4
qY0dpIQePZqZUoqGgq/vDFjxeUvpc+Tf+VxZATDDnPKuOwCByNy70AUdOWM47FAo
i3nur4FXBozFXIc/5aNk66Pdbsm6vK7Hu0F1k/b24xvLpIEHF8wwLoKwUHdJtnJu
PZmQlS146Kzyw2B3FLKFt4Xx5BEPkCR+X36jQajPdN3Gtw5WfeGD3DwZhwZfRRjR
PdyM/QeO4xjOySZL8kmwsqNiOjGKssYnLSSTjmG2sxXlk2dtQ7qhfR93tO76C+4S
YE/2wwq1291yax3nAElpRu+gcOTojarutlUyTdx7JlNjYgR/AML4BgI3hdqo+JNS
MH9NYZVfvVAi2y1U6xvOO0EOEz0S5Cfy6Y35IMaeYPhMO/WC7pRr5m6Dj30A1Z7K
+QWHgKY5034OY6n6jwg0qMQEQx8q6WC0y87z0QE+2uffKW9la2dJEQ7Lr5xPZYRr
1Eye9NvGMRK1kw4FuENJxK08+vKtc8vtVfGW2ZVLqhb/nD/Z3QkquM03R4XoDq1i
/0hentdOW7Mz9l/ah9BvpGW/zFQLVjeYal4yAqBZd4Q/WGgtjQlAOH3zsayc9g8B
6++Pd6rgkjQw1j1KA40riD9zCm80rysMwYn1C4QhaJJWe94sWcNubCrjFTTX/ZTK
rA1kn1OykeX/+g7SGhtd71n7w5iMtMC9Fp76pYPir/PqQhcJZKesqGSts6XCLhVp
65xvUs6K21cPe7RroIzMP0f0xomkWrwG3qeFCtLudMFJcWYcNwMSlaAd9XcT/D0V
Pd/6gJF3lH8sCQa94FO07hZhKAg2JRNpUGB/x1yo3rXtucu/SNJbQm5wGbPORKfD
NFm0dWw36Ya/JyLcqqs5bjy9RzJjpuAyN54vwvo3NRhWHHfJp0JSbvSKow3ay4dY
j+ud7qftkGqZMRshtMEgi8vu7Qi4oVMmMOuaR3Ne//V3uaa+Tmczxo36P8jo3foE
O8/1T56sDN9XkHudv2vMkBESQXTxIHR2N18jOV+NATQrfedt5GrBGhJmdW/1NvlH
AY4UiJEJpYdjf+5kxi5NznmaxJDTfiaiwQHsdjWhdxZAECh8FU7ls3VCd0cdvshs
WK0sgMGcyxGBXwyS/G0uChld5cbJAPGaNfjG/Zqrp3kiMZqSnqDzhrva9Ho51+YH
+Z/yAtl/80a4ilhjxk+mh5uIbflehExyRHIUBzUalvGdHmT3B1NVTzlYc2KjCzKB
q5lJLfz6TDT00Wflmq3OOKaJ7y+8vVFUF+UF4GkfUOTE2aDdG9nc1b8oBmPlkEfD
UODyPRgyz4q5x/txTxn7oCXZIQUUnFnfonIxClzHRB5U5B3Fs1hdBN+fKik2YDV0
qw+bFMpTu0s2XDOG2YvZm2jBjkxddODSq4AflvkKCxpnRoGY729uk+n3+0zEKAqc
l0SPzW6amZsOEfkef5xWFSUtOW3s8AB2kLDYpZH46Se9kR4Yleze7Q4lB78cNfX8
nYPeCKFbI7tvHUz0wSg1L3IH6JpkInP45poxtMgX9aWKZwogQ+oXzKYUTgQPbitg
4fAprbWDBcCz30YO8Ie9R3bNOeyVQ1H03bUyWUMh1x7bFu2PSNxB9lC8zbTGIvHL
LSyNL8Tsp52mJL7dDc3sQwvnI8+zbkjqe5K+nLTAZY+G3RgEA3jwzHFi8ZzNq7rk
dSrktIwcrxMct6ybmgWujw0xqIh00Kr7cWoIAcPdhdw1DNJw1yXe1WSdA09YkJ3C
Q84QANA/7iVz13AnlzAKMo61UardRL6ojfij43yZEjqG8qp6P8DpM0L2U2WEeWlu
GAtULQvnNF2t8IA+GFHnJY6DB7arTscLXnCoup1r9Ii7GnJNsq8dn65MDRxvc2kl
Wmgqms/dWWxBZk+KT0G055RHgfG6DGEtXaComAPfqU1vWlr952rzwZ8pcSfpMW12
ZeGCtuZXmZ0Amnta5Aaf8r+coiYSvUIcVNCo5HeRcwwV2T/kMobI3e71m2ibCKnj
SnpP3eBU84Ej6RUopZohEgRrY5xWQAN1D5sqjX+7GqPtEcvQgocOfhU9B6urganW
gpRNHipvNtFIk9YK0LIS7Ls+33LAIAnW6J3mAdZFrvRL/eorvjpi/olBl7Mb52Rc
0EJXcnrzBjEhY+oX8ruIv2mVEqvIx34+QrByIXqt6KgS/uvh0XOby42GX9K6mt9R
E0b8S88O1hNqP1PzoCtYk0ZHuYpwOwdd7Ulp1wgDS9Tn6ZKzTDe17mnPn3QEcPcF
LRGCi1R8CnJwdEDbc3jeHFYAtGFw6gbJcxtlIoUIJeWGuefnMwbFv0ff6/4PyPh/
AmqB7dONpnjcQN8DNfLUh9kvRciB4daUXjmKLw6ebz3+5GN+8NIWgQ9kav42tqBg
jioP+YzUuqT7B9bQg/FgYldHb7pwG+2ItucWxeVNLGS24vVE2R35kRjcaDiqzia6
WHRRCbb6QUTKyEDBnLjH3/euZuJ6jsCKN4nA8HgzO1VL4mAtuXjUzdcsr1/5pBIi
C2VMYJc2h2ONm5Pl+976tnK14w0BI6FZAyxDxHLK2yGwoM2vffKdplC69QaTVfO1
tlAG/WiTWiPSHkEtDMhprOBVNDKFRdTl7mqKgqHa+z1V/Y+VkSCeN8OhVxsYJz+M
cdiCVcgQYeMkWAjE0gtgMYtE9HqYbvGiL+ijG6vZg2itEBMDxubwIt0FowvH47mC
ELa3p1nFFNXZyrmLt2D+D9DqdvgK0ODmd9bR6BEYplMeAq1Cir/EPM+BRxOKZbEn
anvOqx1Qwj5M1MA388k+McemMjr+xjO33XagDlvSTMIYcP2BVvCCgGJ7gG71Bt5j
W41Z3Bw8TLe0aPNcu9fkEEZxRl1r+SAyXXUEWexQW1fTP+Kp0khRN4yVztMKY7vB
01quQ/vt9ZoDiOltrDO6ILlJ3PYdnm5LWaQtNb6xVghRpveEGxVCeRkPWjCDDmj0
q8uaXyeK4Pa760m5TtX25dMjT61EXxYs4BKRT9wp7qkbQVGmhUA6atk+rvPN75b+
ueizx4v/HffTmVS/781CNYjE1d3BZC2rblyhSQxD4KVUHYx+p36h10/KIrNn+5eO
sU+YDCUS55PflB9AcvcWir1zsZ0L6qYfCgtE2xOjoaOp8hsXxuBYMDYgHCMYpPww
UXL6f6fYRrbz/xdlOowu/CSN5kpov8BUvAsItNUMZd/HznxkPhul4NOqkT3C5zSs
oKIxXi+CKMORBLOBWP5cuUUndOECrEKbDFfg9RhzZv+9ipgwSNKs0Lue3wfstaO/
aqBoKcL/hxXSD65uQsvEY/sz9QxfIwUOUfX/jgFb6Lx4mMy/O+GVawfpdHkFfOT7
H4d/VMy5O705uCRADRczbNqnPWIyCGuy0c28qJR9Wv7jkx+wsoTl7VmlziUHJTzt
tciPO3/x8Shh7QacnguHaw/Pw+IutFTCyB3qvnYfWJ+mNBBhuigeyXZom6pdwb77
wTDeS7CCqrAQKiDBdw3z4gYTr1rmmvAuIWgeuT9yTDaLLRPfbgsaqZPMNSN3ysQ8
A8v9rYLyDY8xqEcRGOrAibyzA7WN1hvZ6T/nb1KyJNi3r3rB3T8fEEV5MIslLrBO
+S9Lpd3URT0otfbWoeB+E3/YMNsClhTkUC2P4hLUWeKAuv+Mgf2F+1bCjN9GxEhh
A0RaKbHlrPRDdIvO4DBlHJZNZDploi3k08yLYgZQPhmt7leElcU4vvT73BKgl1Z8
Fi9NfuO/yQGnNNxOk1inA/1EAXsFrtdYWv25GBojxiTgEs5CI//41n1BEHPF6HNG
6yojXXXfhr0bVQ3PPFzrxtVO4sb8AViDh0RypBnqqWAy4HAwv4aIqdnyu0Am8Csd
LmN2gsVhZJzVyJWZVT/BaZBvvW+ODOhmElTbnbndcMsjpkAd249UxQdZYZ2PLBI0
GgDuFm2Ok9tCmT6Rp1hQzdKnbQLtlmGliDpU6U90iHBZLUhLOtS2+xpb3l8XfXUG
da0ilz4fwedFLhk8J7lJS+TrpqJdsum4yk6mBt9f/j9bzyqSTU3WNpMI9nfC8a2r
n+CNapF0h22tl0o301FkCiTzFtkSLLMrI6EVkgSiI6kjFHRkWtCHskDkctUqe90Q
Yd4LmaeAHqvO6cnSkoMXDRk4fxuPYQzMx+tDZaEC2QmSd0ryD5gyavwPV1kB6Wpy
0YfiEeQT89AGpb3YQ9VqfTW+ze3jQ8uLe3gQcVOwq98DAb9CORHL72QFjKxCOOUD
/qfzSkyCboR0ecTRdJi1ikawbSyYMzn8aT1hzzc4n5J6MSY1FyCVduJCJXIQLTbm
PiyReXPd3GsXQUQKvM+CvRrTwYj1WU+6yzig6zyFS1R1nmA2teh96iDhKJfepklT
1wIUEDdyQD3u0gVtqNNu70d7ykOfGZYW3SiECAW7k+hw5k8JJm8YLmVOGUR/Tcd3
72NPDiTE1PvOQIAj50nvssED8jIEMAO/Pp6t4FcG9uqayh/eikYeB3V6Z2vdbon4
Rm0Q96Dyj1nk+AoRFVr+oYR9xs3+G56SFfwcS/OMQeiQr45INYTtJ38xeDKA7GhY
t1kANwDp2bLSY2gWuStinFGqurgQ9WjohTfyzNh830Z2hZRqqR9HG6huZA2C4VHh
dci35bbHsBi1+r/8zQ9SxmpU4QSB7V6jfpsRpCEJitvsO/ZfaAg7sRdBlaB7bhx9
/DLpooVVvVLw5NoBZOSS8tOsGLUBzoJDuF9eXG9xfzX2N5UBe//WdBd3u+6I5bMW
lIOcQW91Hm+A1uzYQzx+V2vEpK7K4T0U1ypVK7hgcADD264Xdl/1jxsPXbBG3Z7d
PJlVcGoWW3Ug6rydJikjCR1G2ptQJcBb9UOu1tdVolNyMMLWiDFfTKFrLtE2vhBn
Jsh2qSuPvOQAn86l6dKIyjDHbHoMSqr4HlROf+2UQJY8Ujs+gwktE9a1aeKqNLdR
qy/G71rwdSO+BNOwr1XXladpFTSiuUPED/0Jj/JqckOJcBF3ip4TMSshSkXbSSeZ
AF5p0BEiBVoajGiOIn+9ZhBcZhq1vubOfIDIMlWqzerIMhPS6jZyolleSad5HGE5
cIbPwEZm/dv3FGFYnNTvmVhVlL0XwC1msz3EQcoTDWWqkeH1758/MhJX7ffnjU1D
G9O5+hAd9IaRv3fusAeoRLEoaf5OmyOJBz0RvIWxtL1JYptvNzmvi18fVg4oDDIP
cBxDscZ4fvB7KtQDRC1hEfv+iMHGwi1fVL0lOaBsrn5nZwVG7r4shiUuaBci5XjW
r6TqXcv4NwNka/+k/0afIlnVju55+fkcQa4P8SlI49rDE1NW2dZ1l8DPpkGWbB1L
hze0gSHAYmRQ9ocqk4I3+g1A0R2QAIhS0BZww2X+eZq7fcx0Rq8Er/F1GG/twCiD
JhElDDOo7Lep9Ig+aAtRyMaSJa71IUAznt+GNNPc6gYjIkajVXDu16f6a9nN1IUT
pf1+UIArJEGURsl6rPXEkuEha+5fNV8sXsj5Ja0qVKySDYYyar4b6BKeKaiuUfvw
0Io5JY8MAIWMSch/HjszwabRp0Ks+tTDTdplzea1elkVvfQwMTbNoH+05eOCK/J8
S7ALBBv/LFJbCw/cHMNCuW4irMUpCGOlnHKPEemLnQW+cTfktoFm0TJtOfJdbiyf
9VVwJUgtkRJIwOuwsF3GHcpdCTGnfkSHH1m5FxtDEWN5Zs9n7Tlbammex4GDvZxu
S+5XK58UsQxWjjJtwwHFhK9mHGfpiLM0DbnWw3RSwJjW3CtKB2oF+CSq28iEkDPL
4ItgW/K+ZYr1Li5i+zYY0KCwmZXzfCSGj3D5NonyiBZ9fcZr9Jdts/jzurT4HZba
N9hpokzYhbszbTp8xlPP8ao9+VjJeit+qpSHB2vfSVWmDtmn4InLRLuwOjePtBw8
/I7Brcb2WzfBz3ExcSYyZARIdk+GQhofctoE3d8NCkbdKm3j1pLwshBW2Y0XNXoW
mCMscbCIMIGpb3kLnEKFrxyBvasdZWjNWDImYBgm4VVBd4AyVpw9xD5SxLpFO1ka
c+FoK9F7n6OLFhrvQAvvkMuWCGlUmf1tr1Xgh6LMx24GFQvUaFxG0xpKbryd4oXS
0UHcVD8bXmg+zaV/oHK3CH+FmK//06PYJ71KTWyzz/NgXLDCLj2MnuaBv0HHv4Oh
lG049xOPVsxnoP5xMBIBXkYLw4/+AzChYnDU1Fk/5CsIf+5SelRQektq2Ifs6Sxv
TkvYhsudGMq72W3wz5bEfNM70U2Wwi8jHWEdU4oNRI4HnX5XkiRPcW0am1awC1ng
wDv0VgUuimM27M655rtjHiiXiAUNgJWVDGLZ3rKVWNz7NBXlLvgoSxe8eyuklML/
/1XhVHekAcg1IiI10Pu95MhSF5zSCCUWX2qVqv/zYhP8qubs+Zjj+KcxS6l508Su
7t7BROQarbu2+yOrg/yg68d3omfpn4iGFG7zo9OhU7aAViQGP96kQYrXUmQ9k0wX
kv3maniI5lNsbWwbFLl1y3JM5+ZCxFBt7jrmK2e09eOLZytfFlvt/6Zpu5xdw6sM
eAqFOCIlXfD7PUwt6O/L+vlKtwrpwq+mSeEtl9/D5SJwbEKVMDogdxxvlX/R9iEX
6S34ACPA6n+p3bG7BM2xmJkRrnjzori2XemDTUjP4RKsA8huqvYDwfwGhuA0/1dq
EkkpffIjtaKjhdTWcOjqo0/dadUOs+8etilw0/ANaJYYY0GqyB3k8z8Jlr1ymLCD
Qhbb2wzqshxriwIKDNPOXSrOyq9kY821248tQ2rbUmsZp31oqNmxFMFcKU/9zV6H
5BuFoJWXipseh6Y52iLBl+caHTEKugcUjSIUMN7TNC+TIfG+MyxPyihdSZD6NI2o
ADgfnNKDoOiCqfiG/RAbL2PYCD99JwaVK/Bp8GWW07VpILTMNbMuc98rulJSrQRQ
KOur0Ox7IPhH7TxpO1Vi7u9E1K7D2HK6Eo7JWIFG9Dlabwe9o238B9hmQn0wBUgb
VYuDryvHsFPVAS/IVqEpWY4uwKjMpBSw6D25qYFkZrf8bupL92AdJh7CIdO5pGVh
j/VfYP6ob4oaMVmIpJnKeCUYLs07MtMDuiDtrNQDdTtwnHKQjWMkMKXjJiXOmrBn
WQXilBZFwucjh6cHq8aJjPTD3IjsB1q49AFXfLv/PXVOaT4y+UtK0Mg2vyv66Vxb
bTtWgqe1YdOmh7ipnm8HOLDvh+EiHISnj+ItmdFsij6dMBsHWh7J2uwAtgsDxygR
Iqh/dWs976ayUWjFOhR5qKZ2NDXZytG3K6UWh7RRB6Rq1O8xrwgLYef3bflngryG
9ddm5R4720W1HAHKX6mwhqCzJGw685cAoseILxyc3XH9I9Q1di+oic4IWFNBXOR4
ipAqjnLiY2lr7O9LVSuYBgMEVMdWOND3aNWxgpKhegJPp/STsUGnPmX9PMhRGoiE
tHeaRXB9lIDzoaVpiR2FtsK381j6sT9W/bsgF8yBAivDj1UL3shqBcy6t3bI5+n6
3QUMj1ME/3vciW+htIDs84z85gFfcUn0jA1N0FK25akxGUhkLA0fEW5d0FkYZy7w
I0Ek3tUyiZauHcW7AB0S422CHQzb795m94GwRwjFOxEkshGxIdh0KzItG0VXphWN
Y6K+BUu24WgAtpx8JIYiE/AZcSv1yFL/wDp8a3O0nOFXsD93gQNh07Rwh/YcFJVN
SaLT2D21g306RgW7VKv9sxN+R0ZETh1jPYu3d8GUUY9Gl1vp2RQeKi+xwMMl6WaA
45KGZ75R/rsL/cUXPg79hrc9lHGcmRFj9bLwJwp/K2oIqf0uYWN24jNYaqWi3rvk
jpaqIA4386M1IcWqoByKO0/wHaqwuDBiJc1J/1NR4KJZHdH0mjXhrnlRnpk/JUoK
79jBWjTXP+a0TazqDV7U4gXAYv2f0dL1Ho1Zco4t4KUOx4U9Di/+9v5RgUwh1kRd
Bhuk5jHs2QUW87TMJrTG9AjlLUFd+kGsm6cFJqjZe4Fl4nrXCdZaT6cRk6w1MNff
Wr8csfOWM9gYnhxp7m0PZ6UWxNGrH5fT4MbPmILgZKAg7rNaK7Ny/WcYss4Q4P9S
s+Mspn5lrkWgstJ27XjyX0vVrWogDNNU2Rt+67U6zUjGTKuZBwoqfvw2VmA37Qaf
MAVdWzES7dWP+BilWzj+DqVVSrERFlNHzvr9DqY5QGAxLZkQJYNILl9qmTs5pxto
cJtc3QM+M2Wx7PPTCybFVc1DW8gctgWqlUljdEZkhB3CaokPGsKT816b2GIsimkA
EYG+Xkcn3Nx9mUYzExC8C2auyUA4YvPT7GvtGhAlv1ubx5LmUyAV5peHEUa0GQAU
CvhA9nvuTuAftAm66+RbiGU0ou4CY9wVkzTDR/UZPka9iJRXtOyWgIHbDZwTbs6O
AaCl2A79LVO+ZSI9I7c8XT3rvKAmNy/y1VzQhrM4BOaF/tPqh8dJplLlkqu+dDVj
lWRFmTSSxmogykSzzK19M5nGtrocupia3qjwTlqouIcLSZwdWEUGow/Tak6AAruL
qppVOhosSwvWFym7EViqcHH9yDoiXpXc8hJXBGPCX0pJcgmXb+xItRkb38qfgECs
5UphlLe2h1Wg2raEhp1DC6a3wBSoRQtJo+z0CXjFRpjL7+t7xuKkXEcCt97VNEP/
OyhYaK4zhu99Iq3xg9RNZ2HXEXgIowXT12fiL7MQjDZdAH9QDLkrnwV6Qm30IHWe
1nlVkhuPWMltiJ7hdykxsX6W0aPuqrfohZMLX6c3/zBDzgGJq8TB0IpmSNR5cZMe
5kTBMN1YNxOGbs1wY+Io0F4ju4m1/nE6u0Flvo+fvYU8WouLmq4dBXj24YQnumZv
cx2eHmAkpAm1GuZV7oibxwha4XOG7tRJWOPvjMkDjjtItuG7c7yJVc5VWo9Xe6OM
SCXnoy5dV++0H1ayytQZ9mt6MjhnAms5pqX/jn/oKWCQfVBlRDeYfJJXdFonjx56
0psyna2ls2EiDcIloRMRmO1Q2iXOCpvjhNEZdwE5Uu/ZZPol/M3/ugfCvP8K+onV
JR+2gIQ7waHq2XMgziWuxxH+e6zDS/u6ryQFBz/FJbI4Yxv1p1de3kUHz+x97Ci7
1PFF3RYxop8D5xE1ZxjQUBSWCUr8xy8gwXYyvI+QaEKwaHCR7H34BwoeM2TQUiK3
8xqaijbsimfPBGhM0J7hrT9vGd4HpRXXNFeclzUtwnvtvPyjTkcUA9lZKauTrddI
Lp78NN2LdAnpbQTET7ViM6nyIsGKfSDjqy8yfeH69oE500xI0m2G/BgU5wpsY8t6
balQ265pdsslG4roRzbIdSlBjGTE9fPTp8HDm5FuvJTCUIU7wPPkGdnUIRFVFMYo
3MX2u2X52GLiM4W/0N1rHxpokj2rsVOxLk0QI1G6kL0ctsjDgIRyvbRN1wiDjGGU
E7pM7TWZn0qzpg/JbR9BSbJCIcMBxM214P43zh0TMQIfKnITmDCLbOnfiHTdoKhm
4FZaQTIxFPUGg5Mlv0heCnq4dTt4wovfxKOrkZTza8+6E3/uSUkGhG7YQ8uiWQtc
qmfsiQJ4TfZF+O3n2KCdMYjECSsHtbAdoyArtbO8XCaOik91UfycFIuhDFZ/vYkV
91KOrMC3oDv1KNgK9vkmbrBlMvmS9emuZcLJakSCihudnwOvQiC3UYtWJcOv/xov
p+WFd7AOzNs8zL24epgbH0HV8jCr/s5BOdFnSJQjqcqMb7tH4bgiZHx7ttOC7ovv
vV2hjQoxKCVWIceQ7jB/mJkgR+/Zyyrm1XEyCL9XNEvxWGnIwBDq3aMba+9zg6/2
kqwm4xAkgAf3poQqJn9D51UTtGvUy7poBPUmAfUyVuX13Zu7KNSxDO6DNOgQ7Vp+
mtiHtwINSXGG91b9dsA+zQiUYShjuMwmK7jy6HL5sZ7WK92Sue2UtlRzec50IAP4
jAR9SRT7FGy68XTVct580J8gOPaDhRIwexs1Da7tMQHPsdxpzS63CJiuFf3STeKT
lTN+DuokuQ9FtAE6NKOQAT+8i+OclVY0hsJrN5/9NyYzNmGeY9DyNqW6JgLwtPb3
1y+A3PT/QwGvW8k8Mi8qk8AJoyTybMdVWQpoonsTqUcLUlNmUqxJHeZQHkAjxzT1
UofLtAP9HOE9Xau0jGh0TLODbu2detBX2Ie6aL9v+VMiLjtwtf0I2lnzdVdQruOz
r5ahlWizjIPm0ucL6jiuKeMh30h6IxDA5ujjB94RmVuq/J6DaowCxktO4YvCfiea
M6hxZo5iBP79qY2QAfE1aG/TV55uTYJzj6vUZlvFwby13e7Nty0jFTpgmsBbkPP3
RhrVjnG2tdo8WkeF4LoVp+zR7gp3Jm9bgDNLdzxmTYMAeDODnjUIcK08i+aHuPq0
55EhlLxrRze+r+m5NIzns1dpSnAfs3qGnMKk0qJqUdvJDWQmNE06h3t5DJqP+nVL
mZKaB0ejQGOwQXcOvboeesYL/7Y8BPoLRKJDc3f7NgvPEJZLkCIcem9uwqqhf8it
8ehBXaemhH1maGKsbSMZUiR4rPfGKY4pRtaYEZf5KHNtm6u3QSsTWn0wHxs04ZaS
sK8arOQ4x4CnDbYPJ0vOouPvRqF4CwsmirmpWUtZmvSGBxBjyr1/qsQmKbmi56jm
FtisDMKMQQ7uKZh6GSQwBgn/PCMs0FsgzCeU6o587iBaqHO+Qcez3uK/wX0bLGdi
bGGsAMkAYA1hribzPn0C1CjvhTpmtXtaOwyIkbKisuLXDgnkuTmy9fVy79WMHLzl
Bfv4rwQIiAi3WuDqcb6AN2kv3de41eUpHUMd6EgSRtGOOcdeaYTiiOic9BHgoYqm
6fPfwwYageqlr5FvybTnorrkqixJ0yE+6zIN/CMgMhLKBnMHHHI/REhaZGmhl5UH
+3ypx+mtaqg6P6Qea/3khFS1P+AsLS360c9yQWTpeoucReAPN1cvxMJcXO+MTsxN
Bzl24N0SxQeeSidUbvWsoI2bmoEQYlFS93R45gcQI+jJWAPQ9h7VvGtjWRi8WHeD
0bVV3luzDQRbRQ8HL1Xy9yF254PYgvXzf7lrcMqtFn2jjwag4CKfKR9Cjv9G7R1u
9L4Qb8Zxr5NSvoaaw/Tm2Vh1D39qBRm2JkxetSP1K7XTsbukmm4H+9086jPH6zVk
m6Sn97MwU3hC8b9H8hJKxUfyGboIGj5BBo1OTEf8wYZNkLx/H0GbBk3NYxpsP++j
jJ9O61cjShVIU7FWcQFyrUVqv74oycTr5jLOn8YiOVrJSbxHYynnbXd5UoQifcQb
na1p9gVKJZB/9wyGqqdQj/SzvbzyPID6z457Pm0D6QOiZqK0CAFVtBWZeQfXiV3M
EF+DyQuyPLAZr7AF08gXNusW75NnJ1NtiG62UERewisBRRZqu1/i8MEJIXU7LE7S
B8rtv3Bh6dvHfzFHQS7ekeiVjLTtLY7eUOiGY9YfTRA6YPaJwRa5qO+STu5DMbQK
Xi61ONEPM5qBwpTG6UfFBohfQ6OCjDsUTpjaTMt1MCB4zURkHkoquylyFcaUdhFD
k6yDskWiMWLtxDKwtzshJUsU8+h4s+Q1Rw23mi9SpIhH5aJYmDDRll+6mb0d3gJA
LJvPf7axLLRk1fsDJM4pbMdZBvvWigxQK338vQuE3qxMYYbMcHRJsX64+1VGmY+c
4aU4fA7wxdpwNf9H3b4yGFcHeJ5w2wyunVWO7QLI6kr/WlaiXYwuDTXpQy7YbLTK
3W08mCGiIV76sCa18Uk3pcrcmVioOk8GlrfM9sdk/AVXUssfgeqGQAgnBTE1nL2x
Yf2gCf6hXEGh4tK67Dd7w//Kx9a9WR9e9eCdyZm6wYQH6jXlalaycGdjXYk1U39c
ekpyMGaNBALvRCM3540OApqtEq7iKXxRU52nGhKBIphpRFXWtud4M0PUQlbLd0yZ
8aP48/zK9WKBM+pocvfsViI6by+Dx1KBlHTz8v1mdbezZnHMyv+MkcDtf4Qb4P/c
NyjbAkiMpheiA/myt8JQtFZWM7Mh3lz+5sxXPg3ZJF/tQUz9FGUwmo5gljGiiP1I
cujVDrDwJQ/dP8MkYAkW0b48rCOHEa5/AufbKJZCjf1OwWW15g8D3Mbu1K7G9YEp
QgxV5Ln2oH7ugtA/IeNqW3Mqz5k28dSYDGkuB3uUi55T3bAulpdEHsAxFTPaIbg+
k8vY1pOFLpgwqVgc3TDU22jp/dH57mnVA/FpIVdiw4LvzNqs2DZXOzO0xvVoYfZi
4iJr2V6gYw4LCXyWfOdO83QMMmNjawmXqYAfTgAYgHdHncgVENIER3Y0zZNjVFKv
xrqXBkT3Cqqzr0HlRke6CTNAyU3tRA/q8uegIORIzKuprPRr7nvYyWbLKL7wsV+k
Hi/9yPu9JweTz2eqRp5F552OkeG97YOEj3pPjfSLj2W9x6ngIJzOHJgNX+Y7HLo+
C0PI0iqAMXMbuGzZeBmgpYAdbQEbMp1VwZFgNOVD6qNofpvUUdjGAF8+4QSXW+HH
CC/dyjnJOBoQzWcV8ZsWRBsnG0vItDc8BbmB5lCqFhRZOC/LOMLU+Xr4zL0RVvIi
X5XvRgzCRGGil7qwzeb53+VS3hKG97udBvrLWA5ssH69J93UYj2lrQIp1H0MjAMv
+O8N4SiyN9FkZqhKAx4WI81ToE9QYJgM1LnLT4IMxfsSoHx6te2KQzAgYMMidPsq
hKmObbll3b7r3k82u3JONNMv8SZOrM1pb0VzA5fqYWiovBA5RK6NIZ1c5EGAnPTD
J4lOlIuDZs8F5jaa5yPiOcaoLdygqJG5wcmhKpIjV4JRXG8DGFggxmW7OKe/qg0O
mD/mmzCDU5tXygIKSLt8YpzGNlTQ917vug2Zn1jBJ4ae92Cmhbk2IdjWZzc98ZHC
rQa/yC7bOnnlClYJtSaCfMzsPIsL2hhTnNiVL/7QyP5f7NqXhFy800xu2+s96Izi
i7lhljlkEfDHJqCCkjagMxWXc+5r+KuixxeY1mLatCxWaDQCmhwK/laROlDhbi18
S1OT7Tl+Ez5nyMCigTzG030T56s1kzsl6hu5dY4VKAbkYX4LeINMNKEyYDPu0WKJ
NOPnctoKjVEIRaoJiLr1kjC/0oOVllPeE5pZ7yM+41RTDOwLOdXDWFscMJWKovyQ
fCKYCSu0VmN3/Cr1DyR3q9FQBjbzd2VsXMaHLi1VostVVmJwOQopqsKgRHmaBLKU
7dFd41Ur6CR2RAnTnlZY2uftIc9Qja63GtTF0OJsHiTDJRmzsugQnO0WeWhi4CxD
soL0bkoBZYIyFcWVbu6nU+JkUgrkqmFzrOJcARPycWe76vrEiyPWL8SgyY3Kfu9M
YY6wTDLf1ANCDPubmcnjOXVXhOfiCzjJsWDL/Lxb4cqaEwIpxSpdipRP8Bn7IvRP
ju9hZXTvduBqp9KaS6jyjvWsuZ4gJkVXwoYAjd2d/PBdvh7fUka28gfKyMDyqKvP
EdsaeuO5qTey+zPIW5UOcWtJYYu4fqQaxHu8UM+VN4/IMEVb/FER1ZanDoXqR3H3
OLBI2HDtpcDiKnE8X8zx2LD67C7uO2NMqwNdGR6V2c5RCaG7RbcjqYRU3KlhdeAS
jmYJFC81P6iy4322zarKAE2iuljzZM+D1DaSed9EqROWQ7e3uDFPQ4YpmEafz+w6
MVgpTKaQy4xsrg8wCzGS3eaZdH5iQkuxuO/toS4ZoLgJzCWagkDil+XdNWenT72I
Hm4UCZpA9jAclx0szBFnDahBCv5bauOMQPPVaxzTGbAqfzppwWv2WN1hmRzE/IKN
QIEWNsfGUDDDtSsErb0R9t5VTi26MFNw2q8V98/Wg78NQE66UkFqBR48dECkskYy
PrejyWEdzg+wc6MTp85KX8Znn11j1UpPMdPRytxdMxp402syBXMr9t2odiL6lnPk
JaiL3E42P37rIXa31qw22K+NC0qSLF67kDTEHKqJuei4pFVtTDtpRVWxI+xfDpPq
Uvbe95fPx24uk3wC4s+X3mvO2CHKT3cfUL8Rqx4ErASJMdwhJHre6YDeXUk0d4nT
aw/44EolBUCgPO/5zVwiH+cocWzOx9C3a1fygh0x7s4Y72eFHUbshdp+UELAarOm
mrY8jcS61AXP62KWCEMFIIg9nLZyAal9Zf0D7I4H/Eac6nQMP9U7pMxMXs/AhmN3
sXCmXh9yPVfgyRRB7Xrs19RjBmW6m3T/XsnAsdinJi/e4xdL0rotjxA9eMihKPnu
Jbzf5BXWleqhVW3t8SXzlLwL/jJgchrP7fNIYOvrgIpmx6VQW6DFjuDNdMPcS+vA
V6byP1z9m839rsvFHmMiOzRj9el07J3cIgt39J06fzpDJqFAxGx5WgdLphMDA4qw
J69XDgdePn60v6xVFW1kjuS99olhYXmFEVoxq/Nw521NEdDLN/C79OJozCNZjVV8
yhCiD6qrh7sBhfI3e0WxfrobLEXqiddC3cuRa0Bv4BWc0uyfwnvLBIJLAQa3jDPU
QWH+Sq/svEFg6ZfbfmszR+nP3OcTn0i8tlH+50zNG1wNJTfRgQx1L/yPLwiKxy41
OIPUTwzgZsVkuShlgT+j6MRqyFBTUjgYFDKEAw//Z+IM6rp56D9wMBW4SAYpDBkS
a5xSNdh3ysmNNS6/QWayQ3Z8PurWagLpAgYfeLHu5QxxILHbPfs9hlvJ3DRjhfrS
42nEnItjfrWHzphLg50mpsNbqZn1IM+PUG015jCGxZtdGwYhX/iZ+IemZHoYdHAq
/PNYinAUuHg1gz286DCccm28WUoaH9KeF5hb8ELRAmwevPPRN8TabX3FFgWEA0ZS
faIPvK4xY9hqIzmrbdFlIVe9dbCFQeD3e87/gE8mdnun7U3p+ew4hEDM76wpNWAp
mDJxhpuMYh4A0UJCd287IV89J5/FSO1eAXGa4Sr+M8BQjacYX0uMm2SxKDHERpGX
1+Jh0qnCSL8pRCY++DL7nzbIBoAXT0z0WsGONP4ImE9M8x+BLo9q+q9D9SjstLnA
f1Z353LjofRJE7BIqBGKktyxYGQl7PBp140o0SoHywe5axbIuPYc4igZZtiJRvc7
FQ2xDqrcazErtFeSYsn/dbsss69cn0U8Rn+ezVhMdiJa0lakdPE1b1FTY3ciAVmK
Wifc72gXttupfBnFnIzdCDAgQiWq+XAUT/CvllMLl8djSUr6wBKPUyqOMstYCZst
pbqAxN+iJaJE2paXGSWMHKoz+ykgFns0BQMEgIcdchRM5in8xd72kQlNSHMgff9k
7QzCbiJKFZKB+fLtMv2XkM2/E9TNh5LSEFb5wzJSm1kTIY51JYBBt2WpLzmWq9TK
Erj3h56kcWQJl2OGj/HM9tYLO8V4c2v7/xn5cmzJKz+WpPDDKXNu8tWyU3XS9m04
AWnpJg2jE4h5c7LfAAqNbGkz1edRWA84uTJIE1uVH3dYf3ok1QrPhHT0AzhGgOBb
y0dgmhTApLdvke7SIGTmPfQWgaTNyJnrhFOVtGoiLc5NTM11Y6KkaCqGgAMmsgog
s6jJBti2QCiywW2ngCVYFt1RhtfrrZSYbykrrlnMFBvKO413A4o3Bt0UrKin3CqZ
zZJCArkxr8cl7dC6HTjRKlxO28/CmDf30+eNRkTIwza+uSvooGamphRvPtqjA5HM
LIEiwjkaEtDe1URvausKNqWauHWKSi3TUNqguvLn5N5vWaz2WWx95k0kxZUongDU
0ofUivedL4Z4ARJ1gbR81tuYOKKhAMmBaqoZmBO5hbTuR/5Y3KhfcQE4PXOet6DQ
igNk9RWgHJVq/9B4ZLPAIrwVNU1INK+cz2R3NiBFwoXfKYDokKad2FLDcKk+LWWw
fm9J8+sc8Z+fHkrtPwRDbBLe7R8Knmnq2asFN1AqnY5ALpKT0ct2mRNU2uJdkEzs
uL552VaYR8hwSANYEfh0ijqYQ24JS9tF9cF/s11418VthgEwdeWJt/HK/63991Lp
7z2Ua8EMgy154KHCcnwloWYRHOVsR46FEkeq3kR7j4QsnNHKgkyP/UfEl0mVCRmX
Vu3twO2kb6BCI6r+qu1iniq9wSkPa4i9belQyMxyNCrHIC+xkaG1UWAYHEyvvQrh
ChhcEqPZC9lQwcjI4ih2QuUOKjRpf/lauubyz8KqVEHJZN8d0nktUb7becp2ovln
ix2YLxw+hT86w0oOO1hWuXdgrck+hDMH9NpA7KsY+gPSmQTOr3r1qhia9xOgZKzl
QWp8urJNgz8MA3Sci5M5ZY9IN//va1o0k9LzD3Ryml662nqUu/VaLqn4tcDEgLyk
7s/nhnXRd8Lm0aClUplrwBzgTu3qM3xOWoEMyNlrxlyZU0+OxEr7pF/6ar3ab4lr
iSlsdkTzNUfgJbv8wiwF6OAUE9SGf0U8F6gc0xlcXJ6EnF/7weCIkMguCpCNKQR5
uNsI8C5PqbfWeCySzifsDVTwQ+0YuSWu4GFlxRZURaRRuYwdq7f0+KJmODwgahcc
Lva5hgVOMpe7Fay96Mdqwy95migzJF5+QhXRj/2dS0TLiLetrcMPm2d8TwOgunrl
j4WJlltOi5EJJH6RjJ7E41LPEWJL4WebzPOuqLcr3qw0/Hmafo+fGR9hmk2CMMGb
bDgdag4j419HiruGq8/0a31z1g/mky79HcNBlYeye5aGKCmKpR60aLaF/2zPAd8U
pybt35CWviUuiPg9cejx9iV6SSLltz4GSWixyJoG/NV2B5sMeb57BivLkkF+L2b+
SnD0OQu3W8G21+gPufrGOg63fmQzWHVbiot5yA3PYkzd26YPOidIwdlGiVRYwIQI
3KfHUQ2CdLJzHb+0B9cDBNkwdRRDVnBMU+5O3Al97S36nlmM5jSis4FTeexGdM4C
M3STOCjWC3mdCUFOI4nZrdc9dOb+Zx8FTtSSPJTZ04QNOAAlFVZq2BbLvYFEL0rg
RjiqTTWWcsLjBBbV70fuoDo6s1SFZeYTGUc7vq21tyenNZj7T/8Rh8XQ90LMTliB
lfAIr2VaohQ9UOm2btfXOYGHSKMp/QulbxoPj/24EDHppl6+f30asLXEZmE4BF7k
3+Bz83ELrloD16raGBx/eDeW3B2bfr0CQhrVFJrmDisIfUXoDZG/Qu9AMUi0LI8v
ABzmXZtWq/XAXgZHgMmWl/1aUiuJSbEhHj27HRPn0y5X5zY7i2N4Qc2EYWM6RswX
A2TMHPvO6XxtPM1vZSsMvtoe5U8NgdN2THJG4aQR5Rn8N+z+NcA5ThD9pHZTvDgX
3BcODB1hhIvjkSahuRdCYUABKhROKs5iemI/pBfzgAgALmAHTUUDYXfGE5zHSHCI
pUwU8hiO1OD1ETWIoUXC8KBIgb+6Bwtw14w0dgC3BRywy68XWq07rkGxVnBchAwC
riIBegbuY0ANeerfp02jY/nUlrPRdOnwGVrXfjH8HUGXJ0BNRn79CM5OmVq1aJd6
byOfCsy6KwqOOGVuHZZ2fNUAPWMuIUZDnDHVKcBOAthxhGSmPbqlBU552cE/KLG4
/Dz9AP4Q5GCMtv1i+WYulVw29pWaE9kjBgBmkuKfRLjVsS+IZoE91GZKoGBYUqob
tbowYiIAmrITuZpkAEv2M7EhlibB+UP6iqlZFpg+0+g82QwUIeVCnjs7Y1hTicnG
TLjxC1aazxEdNJBJWxMfABSSKqHW2903RBNXFBjQpDjJJ1yyx5TQBywYaE0r5TWY
2a9qa04SAiADM7GImt8qudyr778ko7K3+v4WCBXVvyx5FZAzB5D6RfC6iVIxGJuT
GV4k7FZBnVZwtC+0ewvBj87xmqPrFe+QPOvFqBjv+hdAsqp4qu3/yaLozlDGafjJ
FXlPnN6m2Pme1zN01QMyLQ5WxAIbFiBQXOAiVnSrpGsC89+b8hJXgsdMRBESqoeB
lXiLu2NMdzlywzAHy85doBkWnTuxZ7U1tEbuFE9Ka3AswPa1egX1cXKmQN9g+zTf
htHxYhZbwf2EH1S25mSEdgri1Cz81StfHgh0vICwA3z4r0qv/g/m3aByxDXG9KmN
r6daDp3uk9BVVfAfxZX9AK+jz/NR+CFOC5PyWL5W7QS7SHl3Ks4boOB0r3rgiD2W
4owqQN9vCc17Zg4Hw81MhjxoaXvDQFMYKiNCgbuvJA8jKt2Z7eqLvOhoBJmYjUeH
NU5UWYIfwEUHkL7BvyAzsETZamZUCdwG8AfWt6CWB+U0nHJA97RJWcM+pkqV3z5Q
VQS3ldqpDlKroTe1iCBrbLf7bSygFMSRLqGWwVfl9G0Q8DkEKyn5cfGFnsd9BXgZ
oE5SCxNcjUfoq1zSfv52VeTSYQGS/395Ps16Pqds4bs0gaw68er0iJnjRP4S2Lna
WKn6JZvsvBuTeORaQYPE4j1Y5c4eZaSrzstB55qYIs/0/3Y3DBvC7EhH0UjoSd5X
FqdAAFh3d/RM2aSliIKa9dkztbtahIsFN/75AcNSeb7MSWfmODh2CHpKOWHrh2pN
sg9PsVdVR0pj3PMA+jlwjOmGB1IC2hdEeRoS80sY66LNYN/6dy5epQSTMH8gIb6H
btokcFVMcVJEXrSYN/uoACIiyF39/kWruIDESWWdBeBo9YxOHR1LjOQSmhk2TzEx
RmJqOxiivAfl+TdA2CbOhlG3Xjr3DALwmFaQFimBQVP1E6VOyKZPjWbRRdg8kObO
dBybeSbzkhE+h3mhgcp1rGQxAD+T2tlumTvEyomYnKOWoBJVvntWwRGkPa9pPTIO
0KCww8xyOtmrBrJRej+gkxZ8HqtvLx+jiDRMBgL029NgkY8himqf0YiikJ0F58R2
Mqv05nMmagsBc2X8eHy9eg7KHLEVvh1XRGiwo8mlgKH9a60z9EL1Q6WLMmwkGmfW
bxgc2K1/MpKqhdN2F3kyamDYvcC+DtOlK9g4w8hnZSort+v4fA63ioXTqbreir4A
VNwxnyCaVYueN4lds7/V7nU7WM0Yi1dM2Iq1I6hTQlIVitEvnNy2UfNbncAz6/bL
NjiVtdXMf1qsmpEquClWKIBjfsKvwc6KK/ZKCwTh0fBv/RajsTORgfRQBSDSdyda
OCk7Nj2m6nCjYQIUwUEYiqN3GdcwuWsURN0My98VeEwMwkH/QFb1McqDnWATuMv3
0AFRp6U1C7WqCIMXnr+jG4k471nzBTbi5wkn0i12RTFkTU1OpXkRd5cdg9NWDNc8
1xQ9ojxxZQbsLjE2Y2d09OshLKa8Ug7aJSxuhD4jMMgfg0erPgrK5i9CyryntFK5
NdBheEwi16LRlhsajz3uQGfoLnjEwDozc/EVKuKaon6/2yIbxzrwL+CzvMF1+uET
BSNY01Olizdwf1NAbDqPhvvhfL5v4++224XO+KiBmMW6y178R8IdWkisLnZpj8CH
FCup8ZrKAvAe1r07OiQQ22eDzxqlWhOLv2WHDWIOwVYdW5zH5nleTv9Wak45RZdh
K9Ko/P4qk+xKShEJEFel2HyzqferoKrcvMneppr3hAvrRJpgGSoItsY1BQW7XAM6
Q0qtYzWxE6v/uBNlS7UeuUV3gUxcedtyanT4xTpS1kx/0vs9nNpfH8fLnYMFfZee
3WTlArtWjVR3hctwX/P+wMmwBOi+3Pm5CeaR8fKIdPb3qg4p83wgscxnAyg1+opG
7Z4WfsBmTPDPc9AqmahUIFHqEApk3R0gjCUTQlCKcQ+pXarPQLwA5dlejbkRoVTJ
TVLfE7yDrvk+mPLnMJylt9Yb1fLSgxuu9X0de+4CUJ1NchshXwk7jEQ+HJhK3II4
vMGxcfEcl3Azi8pf/l0cBZe5iynshlU9gSX/hG0Q7QYYIOwS8nWkFh/PjnzGAcy6
My754yuy8+5brMsap5/dByIE/SGvD3IjcoVZnRRjtnSwR/iwzeODYfN89pq73nXJ
TtLPL6uPn6YIIqHwoPYXOOAdKaPawaL+yoMeKoIcIx/GloztcQu2iqdykERiDh7N
UX4h3iI65Gyo+kL/74nx0ymLirkS71QVKTFWDpbJVvaRuobq3KD/QtCluhcpQQfA
kfWy+a+a5pE5d4KAWGViA6HR9DIk+6aIfH9Xp7K3KS5mAOu8zdtG2pIdaHNl8Lf9
bgh79nwAqyyztyiuuhWKIW2Nh6HCpWtlS9ofbBWZHqNJAROM/fzitd4SLyTml0nf
wDuCaMxV3+d8PRL+Zyk3l3l2LaHwLGv8BiC4fKmTZHI/p2DIoU/yfuIAz914Eafm
yfle/lkJyhdyHcyotXpVJP9K1OIMDvgEWwsl+fO4VrF7672hj7nVTpdOXQvFi0xZ
PJo460BfYCrBuXxon77F/mAnLwQuRHEAS+pXjD9oK59+7yx+QBPWPPsX9vaaSlOP
d+NmwplIHm4FdWW4KwloeOzU+gV1OfzdC8s7gghNWPTnO+04jr6a2nnYjb/PxPT4
pZ/yMeUFJH4Wv7Ne7w42LhWScTJPc1HCi+pkpe3+oB8itQID6bzYpKEBjzNL9OPB
rfmk9EYgKDYyoAumjyyyuoAc9RM5eyYqsyn7LiHaB4Kuo6E2iAka4l2m2iJIsmL0
AIicVuEVAHBSvpQtMvHlPW01vVyREYugudV+tWb71jzk4Si/Znd0W90b8U7/FY/X
EQQBrXoipjOXJOxR2LychVA5IxHgVyMROC8Vq1bvlqtuxJVEwk0Zmxm7YD0ta0LQ
g/JbZVvtLAaLV7IArvXq0YpwHPbn0L9az3D6gZLKgB6qZ9HcJMLvTFZKljIG0/5j
5DjrJrM35EheEafgVEfd1WmU22OIhkavNVJ/kjFHwJzHVQcvkrw3knGtfmEbfXvi
87XOvb7GRehDUxsGtQFHBRerHyzG8nBQN1wo4wp1qaQYncffWibgeyJhpVicSKOC
vNyTbWqQ/xz5YNJs3F8dipxCHJzqQIPlShP5zK9OiyKrqAmwEhdEHxVwYCUGSGPN
UAkiKVTm4LLkMiH3cCUFB9D6FQYRas0sWxAGxYWM9g3y78f23Nm8X4Zw1f0S4w8R
DfgPNPi7EoC2ykwSXeVh5oEcxXNUxwWkan6U+ZTMduxVBXlV25dWAtGSPHwbfXf2
njVsY/jIpdn+BGS9IcHX4sn9w4T8gBwQwp9DZ0hVRHNx+ZtExIT+bHgTYLURL620
v1Wn+0uv+e8Dnm+I35cdLhKrhjT4Z2e9gzm+hFZ9cDowwuhQkDqQ/mYUWdZuVRiu
3IF19cbYP75uKp7q/OfRotoWbw8yKf3+ZnGacFf4w8YrYHEQbEWzAlFAvCQu3v4r
u2JRy7y+EbLxbGtfIsfqgm5HVEZSckWR4ktY93s5l+00ibzIL4lNCUomjFiu8bI3
qn4fiN4UIQd6To9/pPUHMV1p2p9Ow54GifGP33LmwgRl0CmvUXBILFLi8PpVFhnf
u7cg/V/yA72ptlrx/8abaRoeY3sM3MQ3Svy7nN0BE/h+eECKMEqpcHIxL4dCDZpp
EBoveIjdwkbz61noJpkQvLoLaBNh0zgtQg0mw8RTuHQj0hqfRVwgOxauhHOaKg4K
voZ3yD9RPZSDFuy3SFdM63Af1CzOwPO+tZ7oLIfmTx5XFE+oykJVoBLmzqS8Y6SA
knemXL+Rp7dnJFAB/6TVL3XB78Rr7fjt0gMDdhxDjsFSSPpCeyljYsq4auio4NM6
xDtMV2/eWTGGQ2qEiozfkr1KEeFBF/iXvCrdzqN3M58b1HOe2wfgr9Q2cn/4Qvn7
VKF3psqBs6D+nSeWFUviqjB9gA8Fmm5fcDQk7Hdh9WnQCwhsSIdqSWTJQhsawRZE
aheWs8IKDcaC0TeZTXlYNm+FkRZrNfL03SAx5/nyyH1BNUY5L048YsR5J1RC2ZfZ
O6qWbISPTX75HI72/kPa65wZi16AT3J8eNjTCSAI94OdnXRyJANZ4DmzYAMuEeHm
3LXL1R8zQOHd8g8UeVNFl3wK5Eo0b6qGiRLPAKES/SqYZ5B68BxrQUbCTZOLbh3s
zsHi3nfo4tQapvn5/FDblqcVMDA7I5WP9rM6obe2cJJcrgvO/9KkUdKh5jwPCGLF
9WVbu9q6JuMVYAKumDcfhGxLJPd7IW9WwYKucZgtHiaYw4Pk+sguBso80KJwLRSG
xFf/LNIoFQp9dMbDCVTli+5+AD62WhVxPmyE3xlfrgl1FWyED6i+WfesGRHIiiI0
of2J8YuHqS5yYrwXdldiG9ezCJsLj4XEDkK2GWkVgkug54HbVK54IGJ/ygycyDl3
0k3FXO1//ZoDE0DmmFACL6MLTuJxnVLG3A6It15C6AhukvLZiNxjH5adpzj0yW7o
3dSsRuZ9CvW+CcqZP8137nFDlmUPvUBNAimhI+J/nUCdpO1wDw9RnWWhlUYM3SO4
co2Kzu0ZQdbIq7gn8YrQGOlruP0p2l18L97R6c6QurfzjPAIGIqESSaBxNdgnXt0
m/F3lCCcr46biPZxqC5OtvwcJEBDIPxyoOgTSgAXi/p40CGVgPVBgsnW6SVTSxO6
0wPdnYW75nMvBy1sn4ZCQY4BaiZJ1UaVPxGNai0h2F3Pum32AtLggas9fb1OC9UT
1AIw4erTKJ5KzE8yyzlV+d3/Sn3rNu781tMlmj9Mw/RbEtcycWAluB6rKq1J3X+G
s+kuB6Lyo5y/iA1zsVPmPOifcYlyJERmd5MeKMnA+uiGLv2ZiESTfyFDp1Jd0Hkw
n3mLH/XLg65biImG3KrV2QPvsE3W0+jN3PLSmaNn6aOvbS+0/P4iuGggmnh+YXZ0
WIbcKzTUo73G9/WFG0aOYAFcCcHODUg1oTLd6vHYJDvW4vZncv68EybpSdcqinTE
V92OT/6HLKnqSq3esnWCuZp25XK9VuV0kriF2H1VlAGyQo54LGISD0Te+tePveKu
Vrtfeo0eivvdFcATNZJLb18wdbXoiEFm3sJhmjNaqQGAHUHvcr+W3mcxCTPe/NbD
QfSd1N6uV1AeXrCT5QPYMgSUAIIOnhZVgRv5oDF3iqcxLv8UIM77fvEDJflytqnM
40IEd+ZL96a0v3GzKDt3zATB5ApGkTw2+LrsfOLL+8wSh4MrZrGy6FzguJmV/ZPz
9OT46ff6uuIkqfgjUjPP8iKjTaVkp4BP41tWSP8JqPlpUEZvr8WnbUkSdPbAMIhE
qe6+BKceZysj7IXzVFWRpONypv6Q0ivRasmFgRTcbl4frMMy0hMNrE3MhOGjjCf+
6bM96Yet1zKlJwSKQAtP+G7pzUq1tqm3a+CeN/C5wTF2RLI+Cc7cT5DmrXjp1FAL
buaCz6c18R3Mi8U8DA3h+VhuQVHV+qEHBDd8bIDZDdBhVuMuwnqOdyZyR8suALiT
iseDX26FXBRNCZK25ItJPnhZVb0C5udv2mTXr3qSxiOowDEGqnApboyDkQsPlcJ0
BSWKRkXOizEA84/yWfAzIM4wRvCJEiPrKKJm5VJ/AFzHf/eRRMD2E52SUXRvveJu
qujkSvc4ae8X/UKIIyxmNRcNom7A+rcKh5fgtDaCC+51I84KwtdTKonld2OXZ5Ep
cOjERduTo7N7QKa7Jj7hXVisDet//GFw3ayf0s3Fv/pri/y+aXEcObdPLBgFpt+H
u1+w2ecN6gSH0ES4SELXru0Do4iXSYw7Az2LY/DkIA2q8BJ57tbUmkpYKZIWxPRv
m6bl4MV+eJrrl6l/Kduksy/pN+Nbwplzy23Qs+fz8nVhtDSM3kr886j19VMYUpNd
Qisc3zQlmupDATuucH8JosQR/vGijrHn6e2gW2VRCsMAhq8KSBLfroReBHWx6MIp
ZXxjQcCkbhXKwArzTINyH3ofphuu0llHEb+HxFMsoeOVoSH7QCcCxsVKBZpOtd7/
ZoQ4FSH6c7BX88v6CfKP3zDDapHDg75nSXrV8bPqb7RJLa93YyeNEogyMwBr6JmJ
CHWL8O4BscKWzktk33kPzFxN+jpYnqSlWlp4grJ08yTUd4309krap3cammhBZA8P
RZd196q+j+QPuwAQlX5xC/6HQRFYNWIzqT7wEg+cTbefK4oBaeosGJnxjckMjEEd
lw7lck9rfA5vi3obt7mb7A+P7ZtnzuUgn9hG8JHaTAY2mnm6cdqCplYY0LGQ4ZOF
vH2+wBPQ5jtr5mOavzZoUaSCtTpgq6jw1NvGECS+ZZpV1DUO2xAwBvQNj1zCmTI8
0tLfRaInWkfDGlGHplzq9AfDmtlZogoM0+Z6TA+Qav+ke7V7Ql42/5Nhc/uNKePK
F0rpIomqausT6ZtZJbbvMQul2rie31E8N5K6PkI5xbdcjx8F3TZ3FChBVA5a0gAn
Gamdd4qtbfhTHhrv375qRN8/4PRKkQ7Wnc9c8PaL07g2bQ3mxC31ZKtCF/OTGN1M
twO+14K+DcEQblO4SpFxUPsPwgRpAGLUwi3EL88xO8FDJdrBgu4Stp1gsP7C9DFS
CK2oApcktfSkHNmFoMAbfCZLeFsAwNbR/b/jopF0vjlwFxr0PMEtXWExtKLlv/RQ
brswNe1/AtqJzSvNqdjjGYhvyFICLQnTz2ttjbv4jXo2bj5faGaf600MMv+CsVvT
fNXdo3TgEVD2y1A57/Y3af3Tcyo9ZpI8y1u+b4Ai80oB+Tq0U2oORCQFz/+NNPmq
yjWXjZ+0tEcRacDgsR7XwlmoltUHK5caAKKqAHYq/JYsj6SpZeMSVY1Ro0OMKVe8
ucH7HjHc96WPoUMs3vcw/xzgChCoebYF3d2QXVUTOpU61AFGD1HWtLGhjH6osIxr
7As42RNCr1ZiMnTVIlg1+1Ve0/KeulJmi6gnVekmBBrhwWPXRPVGdnGQ+qD124ob
EreP4Vr6oTTkkiSu3NnpouhYv/LxBN6NJRd6JLznb7eHWigFQ6R2uNSaSEoWJKXC
vtbr3E7RzPUTzyDLmZp/F15HrCtgeF0sU/dGIfsUIaWzLn8y3ON5c4oEzpSJFeLy
wf1ygVRFkgCMp0tfbuiTF51zxzFxjb4MXkkHtltbBAI8UWISRV2qnKSiIV9SyAke
/mO9DjMTrequDGPlUevSk/MqkMmHg2SR+P65ga/p7u/UmVzvJ9alU6k1LtgKfWuz
zDt6ImaGUDIttXjHh4/5fH4Qs7RxzEkkehtKwKZiQorD53QQr5tu4UazI7YdpszF
BcCW/EnD2T0ftEr3PYlUYJuFCzVN2EWaQLH3EApaGDrgeES6/tieGHrH9QzOZigp
y7LVAobNAoJpZ7NRKIDNUPAfCr9dEc+h6/Zi330nVKyblGVWd1esTghwa3wI8TUg
Fd2hIaEwaqX9dKWjJ0STzxnziBr/5u+/ZU/kjDFzkwMfE/qXPFnTNVO7t2xADOLh
AMiLWlYebSEYCmNA/bvNqm4LOuMsk0N3w7HGZM4t4rfUKslObYGMIhHLJnm0J15K
dOgCpbGIisGtkCyvBCSt/j02oCtndvzeGV6ZNPve88sIqib7nCZ8pqkRMo9jnkfV
OzRj+Xxwi/6rsQZgS2xKMxXmsq+peKztVrS+RukjO0iRnt9sZvpgfbETbKVSvb/t
+RSVjyN7z6OGV2p0yUHkr1MItsuZ7aWkGO06YcY0IMIfMM9zzWfy+9ZdQ8p2x23d
qAa9iUkZ2qLe87mowUId+QmSbdZfALPNH0bs2CjoB9kYG8qs3/0eLTrageiHBy2m
L5EqQ0JQZCXsLZSyTgwPYASHyLyt05Xrq2960W7ftezG76pRsY1DgiKxZBBRgDdC
cJoCsW+LDi0+cxMIWOjbwaKU9rm7+n+imc+qfn0i3J9n6J6RLQS65HmpuB2SKEXV
EYCsapb/SZfGBd9wxvFp0AnWx/SfFV7C4qX9P+1JX8HsiFsWTZnDwSA2OXNRhIKT
nX9/PLeWi4EeajJ2brtL8i6JALBeXTVQk/F6IzYqwE6Nbez/Fg8ITJbQMmQNvOxF
bm4ce9hSViWO+0mixuKorzQHKVNC7vgwlvxh4uSFCURnQNsi8PLjX1c+xHsEl+Vm
YFwbC6VrBrFKdJqSjkJsNAkOEAxPM5cQjlZH3izAB8VqiLpP9qAEno5zus/3Whko
lYTJIelStGLmhJHs3Z0rau08Lk4ZQOw9fiM5m0SoRaGehsBBVOKHeeXku7LJbtWO
bKEaUTXw5c5gs4HRN4tOm/1bDHpmT0N7blxJW23IWKAIyMhzDPLB93uMlCHLxHx+
FxT8sm1xgx+oPU6u6k7GjbdRJt+dNl/rlt/sEnpA4woOoSYc9x2e1lV5TwHG+FJq
4q70cgNZvPhaOc32BZzEVimJNnhBubrk8fwhmSxt7n8LqqkqfMgs00ZVJblpCJqG
u9WPxQYySeK3wM50IQCv6JEelSinaGw4hca+NJ1/12D76RDYsV/idDXbw0yWL/G9
3XBmBVm2VPcjtEtkr6wxAkz2hqEKLMq4YkrMqSDKlDMpDiMocbjcmIFK5ZAc775/
Qjx4LB1jYKcHlXVFUNayTI3wGPHwnnrjieJJQpG+rg8mVNK4qvLGKJvZyaskInx7
5LVw1g29HmJIzD9UkNqpHWF9peF/tJ6Cw+86dXR88jRtgfwxgspdeuKh7oqEOJLV
yBOnwrn+gqnZbgDUrKXPvwTuvEKcweCIFPorUxwWaldRCE8Xd9U5qIdwTllp05WM
34vq2wV1Dk/BXMRS/DChIkKx0tyNcqCpwPSU/cqRdQ9KByzYMz1HGAXdxCl5UMcp
ey7dJRpPTdcYOi8TI84TmnV13dVcn6AKoE2N9ZMk0Idk9tPKKh5Wn0nQYsU/yimB
r9N+5gMECHrhPUQA16j1+oTjFe3Fsmt5yqvlVFtGgnvMasTWaxrX1f7idcBQnTtl
ccfJq8EnzfkwYZgTi5XnQQd8BXJyTPjNvP/lYw+F1p9zMJz23oVDxCIXIJ8wz1aT
OXExfoFx7anfysmVJ84HD1YU8uRBrLJbwGYkVU8ASPyWZFlpsYAutwBS9IThPCy5
8UzGkstgrVr/hQ2MHKxYLlCtoPPj1bjoKrxYV5wfbNxpxze5Z10sQP9WzmejwSiB
Fx4MtwC4bCrR9pJgAtWfztakZeSXYohKbJmFwyLbQgvZBOzFVN28MYZA4y5IAkG+
XVfGl0IJczx8gZ1+9FZ4XzmhczUXmMWqOUaIMKDYobRSKy9YAPPvIdVeXkt2TS4x
L4kjx3Cyo7Rp4G1+bl0AFWVhkkRnOAAt+myWFRhxi82q/54In+F1jxIn+Cn9UCXD
vgkO7QdkTO9YyejN6NhWMe9wPnBDIP+OXHBg5dF9OXK7yJkPkUUWEBrAGJgMNRaO
KEXieFS9b5vHR1aglJusyECTmFLy0J9bEmNb4PcKzWPgLukej7lWnOvhkOObuZfp
B9dcQzr7Mmic8fkyFlVWRm9Q/N5ufGECErXta24pUwFRwt2GVen9Yzj1BBtOmNzT
qhRAYNC/zMw+zEeJDCE92dtFo3l0b8o+ih22dSAxdhXMSfDkoGOmkKZq5vTSvbAn
kPrLOVf4D10Hjuv7iDgxFGBnuA3rPCP1BlM+XfynPadyldwA7+3k39JnXmuit1zO
Bq7iGVc01bzUF81c7GOfZp9EBBhbjMgcUbuui4dA7UvcjIUJ0/ZpUstBCa8SSyxj
+qsGQtZjI/70eYAy5s6wFLN4+feW8y1E9rqrQHgciB4SxZYL1verpNJ4DYQPWNgg
bI4kQaEJ7iijfp/kXxYijEr8L1ZR292o6JLolLv0ZKm0P27imamwiqOF3w1dCgeB
HVjHWloVZkJztUt+J9TL1XgrEt3RYKlHDLzeWXFP7cpmyJYwTe0lyVDsMPTjXt+l
obivndmGuI1KOpe0HhdMtD+5SQCmFz79TLNwnTlttLR2Eo5HDuz3YT1YVX4O9fpJ
txSZY1AkuFbtPKFhEBrQWIXd3KHzog6RjDaA6ovo/hB4c6ud3XzlHPoI9OnYNU/S
ZY9c3KsZaoGETWcmels5kFbkmUUBuqjA2edb3w7RnODlst3/GijuHHJsBA6hVTje
f5e1DojY9iBGiH7JijMOL/SliOAghHl6CWZ9fBXtdL9nMmISaFji81rna7LRfeQx
BOluu2U5M0Jr4+qhoxFnt0ufWdQcgllvcnHX66Ywds/GjutmFqtym5U90eVui9G6
1tv6jpj7GEh7Li4Scg0mj5yuhaZ4yZQ/6+I6v4mFZhMbgEy2MJMzKHdLA7ykb7qd
M/4BwEPRx70fnyppgLdAmGReiT0mD1Gz4VCur+MtqeS61KQ8I/WXGokaYBxm+h6y
qo/zCAissgHXDJX+sbsAjXHFzA7VdJr0ie/BUsnb7xaXX1AP6R/ML9/Zb3xkS/hQ
OBMXlJLeUDfVuJRMbQwmu38KpMuotIWRe+jL1mzqryjmObLCb73BfocqMH/SUgQU
jRwepMLX+WgOSG+D/HwK164oxnC4Z+ZN68qAoQfSJS296bnRKHLPV1gN+XcRgJlG
Axn8NCTJ41RNrRutuo3yguT1KKhF/sQuYIs0MzbsqEsq26clAnrjoq6xKQXbJTwx
ZS9X3iEDa0PWZlP0GnjWJHQLn0jedymTQKZUZXIO0V8qeNRaa4ubao1dNU0U++8X
+gE4Pr+cDGLLbJY/DDGREQWSUSU2DScILgNsi5AWvGw7tJXjmUnuAGqm4eTE1xCi
ZilPn6dr5P2DETe56Gf+4Hj4DfLSswz0nvLEAVsWwBBgOaGC4PGmny6SN6r8HHJ4
vqNsoFhFdvlGVQOiUjafVYSgcXw1zjef7ubxg1eRs50ZkoRSMwMVpBOss06D24x6
RwnSNLgrqxjfOAYzesgFSJ7NZZHGZSvR06hnKrnSV1OS4IMvKW1ZDnmTnloL1TrS
dP0pKrbYx1l6gI3SuZpLMaXx71Egg/BzvV5fIobL6YC5rbsl0OyxxCMlxgAvrgh5
Vw4MmyUx5ywApyhbkPc/PFuRPhS563+R1XDFOjUdbpMwmd7udtEq2/D7280BuLJi
uHxLKVtFDwGAsjUyjjvfvqA+jCvBXMMAY2S0oAhDX/EOH1PggqkAkPI3GcUGLZOT
ZptS4E7g30SmFpP3kHOoWs8HTSRJDwTRn2ya1lXR0dliEzq0L0veA12PWIV2wync
S4TSt9o6vlo8HskbB+EmZNqLw2Ofd0j0z42h3Wt1M+rtHOxOctKPnS8pMxoQhIt3
dW3H89L6R1schAcekGfiOQhf53M7enteOjWoTjfgyvPWXnxGjfYGNpRhVkZDDHUK
Z3Jv3l7ex7TxnD1GT7HyrHBpKCZ7gSSkxFrlxwNt5IuxHshmo+HLf+IoglnbpZLx
2tsbWq8Fw15WbJtE1CHuUDQGClLNJmk3ZJSRephSEcwPywxY1C22nZR19haM7yj1
BQ3UXA2vdGN4sOs/s8SxrG1nk53WjRkJb1f8WbFFMFIdKYXzChkROMHVkxYtQ1bg
0x1Q1+auILMZkIKURDo2HMvzAwDktjF+z+I/CRP9epZGN2lgipPXaX6TnCY8zF1L
MRe6yraXsvz4bvJxCA94mgviI/Lz9cwOFZy6eJymah3LuW8jHtCgxP3HA6wYvuNM
9JjTyzvATQJuFvCFwmRTibzikfD4QV/WA7lerFE2nkWJgQ0Hg6Ffk6i6Hh5LmUwB
DJUuDhpgGzaqDztlFgxSToIU98HyLmBBDo1Z7Y/YFoGojlSZBs0FhI4XfOpgA/23
D7y+hFj5BIGXjYiHJwrMnTmRwXbaIhc6VeAL6c4T/x2Om72EudIMwWvtKQhfa+HA
phej4jt1o5a/zq2K0mU4eUXLsIK0CnwUkYax4RKDiwnnJTiTrOdS2DgcRZLfcZfG
mD7xu9iWcAJsogJZg1X1olmKiV+Q0EfYA9ce/jpfrngvf+DrHQIU+CskV7uuWdiL
Ak0ny0LCWclnPmJTYUavwmkdP2HhsVqROMYQ9JhHx0mQylSuJfcdAwFLoAOIFfW8
VLkl3N/RyGkRbXe9QkbEsOETR5XsTBKUaYQ+ZS0Vicp91VtbQpIPSCSSff5UEEBI
m5pQTe3M7T+lVznaEtMIzLQBiMurgFegtehL/zr6zVtnliWBMfmNv8Y7ncgg/OHA
Bl2oaSQGDilJR7p6/tFGug79iUoJqkcKPP7mMKGjohlFMjIHaGit+GYdef9sy1iG
PCIIlBYOggdNoqvw/C8ZSphDHCuNUURiyLjuU6OOaz8i+isEFGzCUtBFIfxVwijt
vDBUTO1ye2u7D7+qEeliFAk+/KDLQvAwcbmdEJPzzP+fa0XR+pCnnt5Hge6NiUIP
Fi0d/2Q+eEPTcz0Zg3FrcPAzYSf8zypvDBFVgd/baRQx34pj3sczVSWz2zssaCzK
Tv2O04JC5wGOxNbtYPBwBrH2AqzWkTfphiegzaI3BkZuNpIibXpH6V86eXmp3lBp
XviLiJS8VhGmcGVuI6PDEQQZTTasF8pU15MDIxyk0cnT/NQSSOT3BF0F6eGas2wQ
Dq/W+smMAzt0lvSr6vVBa5DFovNhS3/0MLyQkRqT3lhzD16AmOvdj1Dit0w9gaP2
1jXg8E09z3P9qumCGgf8QfTVaDD9WbD+ezaFodzeQ+gp/VKnc0t7UqgVR3kNzTFA
YlYK+1TqezjeV+qwyY5GdoZsAicbLeZ7x5FfQeA96wsEw3BGs8Iok/1e7Piyx0b+
vmIpcvqIG6WHlqmEerGMRJlCxTl3CQfg0QHwYNCLeCzIioEC1UHc1X468klIHgpx
7kOIMkfoPNdJKqgxi1qtO/rIv0nVq5h7sVtrvpPlR0BScrusBatyaxktjk8JSgv2
Gv1q/95QOV4wKpb2J5OSkI1UEErV7r0pXtY5Pd4+YuGtSOsF5imR828Tqs7+s4Sh
7v0Wg00LvXa03jR2SMNjolQID47k8oVZas523Bv9SMHiL5cEvVT75zBlR0h8m53/
cRkMJSTJrC9+Lq7tkzGyDwEq1tz2UXlBK0sjZSnl4ki6y5xMgx5C6BV1pRr/75sP
osGtytDjIhi5uVNw5DN2iAa/c4FljDdVGrDJEKLmqhk9y74MtMia/t6eNfKncIyk
sF9d5zuQwbvFRCMgy8z9LPXk52eqti15+8RZETyzvxXqOL74FYkRBgxILFykvNWT
YUQGizq6YfD12EL/tYJdNN0szA+S0v57ixrAdQeMYKih1hu9B4kFrQ3kPtZYWOyl
aFoYtxzXJcbxeWHTeiGLaL1bMIxzAPjmUjBaQOV/Kd0aiVpZb4yA7BjvZm3nfk41
WZ1dcfHiV3PnwZGIPeyUXFgPkgeJVffUo2igQxgPiavfMGRSZWBVtoPrARRCCoTx
DkTqyAGi5UB5izTuNCBP6FdOHiwoDtA9UC8XF2NHk4TQEZezvFhtgrGd+eBlA1H9
huo+MJbHQ6mr3a6a/HuHfOnbIOTbrfKY3OM2JuB72RiGDbeXRr3ygv2W/vykxoNZ
1E1tOElzcA3lY7zS2lJI901yn+Z3K4y4SkqtD5hFs4DRfIL7Ezimuun4h1KqnYXj
0a/DnaM/KtWZK/USTIyZ03KUihQ148TPbMC7zs0L/wz8wZY0BgGkHfAFwWn2cung
Qb+PBgyrEt3wlCWECh8uNPGkQw2leMHMkqegXvRjfJvyBNw2Y+xORTIQ+sydu5z8
wEi7o4voZhwlrzOBigUIxFjMOVwkNtD/Uh/ohg07Qqsn8+YtSo3bxkkITBmOX22s
SOKbTb8lyc/d10NmcDsuynfj/20vDNqXsxKFPTmynF3rg8F+X+nBpCr4gKCQeI8B
iyXYhP0sishWLDIHgiPc52P3TWjdGsvwbBtMDsimIYEi1/VOcqIKr95QxBqg4Ltg
c5qyuj38MziXwrOUUJUIWaC5ZmIGiLDAQmGpHkmxHUHrN0aM5+R8lMXK+e3FklnA
XJZnLGEcxiC6FKvQ+2MZl8kBH3brOTF52TO0LX+k3g9c6stFBN+FC6Q41uJknw0G
mLMomVsJ2xIktWSq9Hqp8w2ys18wepgf3PUun0hPde+vkMeA90GAWci5GuU0D/So
youMUE+p6uDt2R12QvgTSmBqlH58MVp+Sgxzl3QI0+S0l3Pr8cErCIK1ldze9mMX
fDkmtZxkR3GfpUhex5Ovo6G/6dZbxvELHhTu59Ot+HSRUNhULibQWQuTcwr/nZhN
YuFan+S3UIoxvD5i+rY4e+cKCn6+ihcOeSmiFkpxb3A42/dUWoll6qjw0Vwt5IZc
Jbx7Rp4qPxfqv0vzr/30BEkQAWf1OKaMaHr29DQjocBIpV8A4nSUvUQR+XtEQB8U
fPEtjg3uKIGMyazWcekghTIuSr/4qdM10USJEaaC0rRo9kMP8pJfDBaZS/cRjKAq
oyR3dtrH7f90RMmnDnZMeGHa8arcKvwaqGGePrVmJWVgxTNnF0U0NwZswpM8OW5c
gduyTehzQ5ThirHHalUwYJTPuDdTvFh2sk21yGmUopsZO4JJOqjMzIXNT4SkdGd3
K5RYG/uuzNjcoARMSEqvkDNGQfPUbEq1XZ9r8PHVq0arR16BYTnJ9P7L9PSJByMa
pgorJPXAUo3mEl2baO9LS2gWtVoXlMlJmjDYkSkNPMDxel2FVbnYqBBsCeSuBEh0
gMobAtgh1VDcInLlE5dfXz84Lfyhi5umKkIZwHtxXdLulMfNpurtp9l6yBxfe1bl
nfAFpQeWQs+QMj5Ge4gGXdzgZ8PWwOHReTRj5h5swwtfQBywNVeY20e4K0rzCQDj
hnNfpugFDFS2es+NpPptGsimKzmbizNJN91MSyRrCLPStLkRJyYCV9c3dmZgOXC2
6f7tecFVPloRK5qXezKTUsqwFmnZ5o3BgjVfRSqVPh9P+Ejd8wArWH+8k0nNwe82
8Yqt4K29NqDDHyy0m+tws2Xa+oVZI2IhzU7gNhJb+ez8Sa5M8HZrrXUTrLa7cNnn
dkijmhohyaNhGm1Ir2uopmG7jgKBxoTwe61/2Xc64wvgnis9kaAdn4c1H2OpuASa
tiuFTQlaLG+myE+wy8iN34GNbmUr/wk1AN0z6E319O5QeoxR2Fsla/KXU7BzAYKs
02N1s8JV5DUMSY1GFvMrm89dMov7sptE+qBG/koj23LqJ6ry1JpjfbNGAv/aEEVy
Q3npDJ4zbbbI15rPtSqJADWcTnZOewU7OD/z+hN0ba8XNVskTgZPba3tpa1zFeft
k8qiB+9NkYV1qGxiUf1Kws/HLEkHx31CVg7AmRVwMHX/mGcxcoHObZ246N3B2gP1
2nysuQJfG0PkOjGd0d+CpFofLTjUUzvCBZm6JQ31Tg/RSq5hIiT/901f+kf0pOzc
pkOCT9MbB3rZaO4EJ+RIeNQVZIl04pKaTIbowh92xH4tbkGscLGuy+o5YlaumkFB
EJZ0OqWZh9Qqj6q1xkzJgtvI3f4EWZZZ8kZsQaBrUAmUwrXp3a5vFMbTtRZUYJS5
3Lrt/dnPvw18Kes/9va5y78K+yFAkWwgOHvGgGewf4jEwnend44wILdaDFDOUpe2
knfKJbaAm+vqdMOVXFM3dVDUCXSqHlafkA1F3+BAmTljTOhsdDun0+0u7XviO2ft
7qsEbdGQiN5qbh588L5eSg6dtwvcLZ/3jNoz9AA+mlTf7yZakI4kbFmXYgaJ7XAt
ZkKRGpMkjYLp4Vz3Nd65EKYt/RDXFVbw9l8hc1CDh8mOe6JFrybDT7eMmF9M3TGo
Z7Sd/fxQH4JNF4MhrhkLyCNNsHIIWHvCcN5XpAFOH+tLfsqdlQmPSHH7jnnc6f74
Y16tMF+D458Vw/7wjIucALv30aKntPvTwWWjMDmI1Kn8LIXqba8XE5QIbLXHhirC
aXpDymcWBvZK3dPMDH8D3rKEnvRWr91CvqEMGAcmWdRtshQ0owoxS6uZkqrMjfHD
7bMPJ/dICAuHfJmBnKNomjjcbEpA9ULLHAm7Op2ZkOxMMjhf4+wxm2aPjcap/3QV
kBQ42AST4+NLNsdmaQQNZttQn3Xt5zZalrb9eAu/zh0asbSbsTgd92mzA8OsDz/v
XEZWASWneW4+1ztHWIPDtW76xS/5KBsiAzViSY/09T5sWQ1nWJscyvjgCNa5Meh/
zQ+7wnl6cBwvFSkPebbaXyXgj85Ny4bAl9tRJsc31o4uHvTfPp55cQhQlyhDiHsB
FrURL5PJcNacnWSbWB0oIKy/EufkfH/rdtVl+1Cg/cs6Zefz9g2XFv5fVB4LXly1
r4O9QbDOYpzWZj2IzHRh2NHqlGMuabCT7Oca4IEWM8Mvsvm2vhQC4AdZvzHa90Om
udA2/cO7V9Zez/SkRQYNtsNzcYd7BDVC324oLdOvdNoLoUTg28PEKDRNAqniqyHb
+VSMdBt0/RW72SlE4SxlZsZr40DIjivdjsyXirEkmOqsDxP3x1jh/bpVPGzgguz+
+/pBY07+nG5JVSkXYyfw+VC4N83cakj3Ai7NoWbgfSlFlfqUZx0UMJMQRxE/ZAmk
QDySXCoyL6DEattrXq1x8ixyd1f0Lv9RYKa74sm/XWI8BcuxbqWlk1J4SKLyaUDZ
HckiAvUOKIEbYdA78/2wOcAR9XvhRaU1lyADKkoOKec+y0mFDuZDidgddhFRRXPT
tfnbarbisbhiyhjIo1dFuXKhvwyb127Cj841Duu179jVpjn8fOMbOvSgD4YhuG2E
e7xAfq7RRXFncuD6QB+k6pYfskMrtupAQ/i4Nd0fBQRIleYFrKZp75C9jpVTMMNd
bDcOOa/rH5g0x/DJggVbJN7m72mam1ooZn5Bu39x2Lpbo84lh3O6y056S9V10qQs
QiWUX1ZR8fO6O0T/kxErA5UX9YS1OrGUKsCpONhbbDFKxR04rTrBRWRy6mf/d38/
TZII7mjQfIjs9tRqwpd/Jpn8ZKGkTc47fFlRj73ntd1y0EVKT1gHmGiz5N3eQ6M4
BnVcLvnzKNEfB4S5StRtB0Prk4lBnikSeBzy2UfC6XK7oCbGXH49LVARVP1v8QPr
4O3B7lvzaZ0uFKHYl/GzM3p+W8GqpT05gtFTh4sxIbPQ2kTvRtbotf/+5B5ELYNC
fDgYr5AfEBacUp2ad/hu+dgJlZOlsuP8tpEbIi630uAOR1CtXfq03qbfby/yOApc
XvMIHITT6Kxm+Ed5w4uA47o4ioIRvu9WEltRuOGSvrrvPEJkBg5CA+FEdMdDLk/y
VULTdxBzLfbWNWhIAljbnjS/C1xtepTUgoBt+r98HlSf2q9DtuZaBnUSyao+Q+IP
eAOvx86LOv0ogeeO0x2SKi8kZPaF7M5Jesu91braPsrd3PMp2BmftY6hCzAMG2l1
K0Ep0CKCsQrKDUKBUdzjGfolQw24eP8VIzynxJrgpw9hfXSK/xE1GRlzvIto8Pb7
gHxbls/NBirEfmK1PSmqs13k18dD3L7Flbwv1tcC93KLJTpE8SS9/ZgAPlmZoUud
gJjDKK9+2fEjM2POXjFuExxdQxWIxn1lFMGaIynyIvaPT7Gx63/AFMGozV1Vcshb
0vKOxZXsO2NBeQLykUthEi3fheNRBitsg6HODz0PEU3p+tv0KYWVgibi8sa9fZ3k
UzY6TLEB3+44l9uggaNnRIuhucZ2QvmbJ1J9YTOGB1Ve5RZePWvYVY11pCCYp4zO
dZKemA0m05k7hdmSvDljFa7htXKdHqd6ZbfpPBRJ+jO+SUpWSCInNqmm2/q/ECYY
KjwcOkViy8rh1ApcAoPzYbYM29sfwgCvanbB+e5LjZXxd47GjXI2Kv7l2Pv5n3xi
EsVFJNysqvF+LStbwRsaDVf2G3nc9NYCBIqJxOe9B6ih3ads1Ns3nFeR8EdIsuOP
0wQfq+dNBe9jHZKXfvPiWefJVS0nuSwiNBvU0SLQx4IHZkYak6Avwm4VVMgNd9v0
ZtQ0Q/RrCTmVM0Ro7ctb/nxyA5pCsNc8Avo5njE/Oh3uV5KaCWI+XlHYdDxbvUQs
Dqv/y4KWu0sx3Bxl5L7G/fKAmHg+S86j8Xu8wz03JOE0gmrSjdomR8KcnqIM3ykr
OOUI0Y78IkS070alMEPZkVxLWF6ByZm/1ZOlcj+uVB8mjBZyn7e7fHqXl2Pr8S40
t2HY8khIEriEM4FteeulRMi5K1u/4Uo8fWpuA1uYv5g7W1KAmd+wGNmsytmkhlaU
aj9Pc312WgraLQv/I1ojJX/0WtREKbFgVE9+hdcLI0Y3GaxQqJtOzpeWIc9VGXU9
JAGEUg9VKluLthxg47q1inDltpPbyTVRnNyyqPquArMWcVj5gzwC8T1yb99lunyI
NWaP/czfKIrpmz12rSrVwh32C6ua2CeUM+315WdJaH+pk/j+akyGyv7AFYQLPoMM
5wnFOPIJmbTHqwyuOmEkL3dZxPX9Qemt+qUekoTq2w7vU1NNcYk+x3UU1mmP53/6
WEPQ+L60LypihAHjEyqERZPaEkVUKtQeXDADbLV23n9sH0FCUp/beN1RWkkI9iiY
+g2bqXzvDn2VEahq/3HvwTYPhGuSYBx7O+0RcKWmIMGRsxqGe0eg68ICIA5ywc5L
wdnuP1ZCdXkcfaq60sqKMrC03VnqQNivYol4V/2USkeu4sSUzJyIQnmrc/tErShU
QT6vzYgUK9eH7qMTOw+OX5TNs3xX3nBy7+jcsIMJ9W0hZ8++AhxMVulT9hDz1nfm
rzpRo3Sj/WZ3OgH3FSvVEEBFKzaCE9w/2RsCtqrJCkdVecA0Sg+gufocllHL/T2L
dtHSw12EwEVABFwHxTqy2OaHaTI9tv0DrT+mhQdWaiECa/iSfTIs5kSkb3TWYao/
VVkRXnEjE0lZB5OKbXPEMcQaE72lN9kQbSRbZoQ14rHOt+UiQmhLVQT9O6SYT8Y8
jqf+zCXaLCzOThfLwbkQj2ZCT3RBIzda6xlZeLAMrIhP5TgJwUCeVUzv/q1aSKVq
McUgFkpBhqEONThZphDAZaYEnjkOYdNwvyzViWyYQ9gsNTurbr3YKjk9qdR3N/kY
7YVEqap+vLMBYGszdWl6cQ/NB/HJsf5xDTXr4sIeLsjeukPBSlrfWkgSXB+yUSKk
N6gxiVI/XEUAs5HIqk/SPUwKNKW2/YTs+Cv5+k4792bwcDnjIkEn7Pv67n/DooPG
urAb6dFrx/gmSIBaD7wLVCl9yNeLbqnfy5lzjn2YMavWgHcuT0JPLspIsr4sQFn0
maZ3mOwbtrKKQpb/d4yjLXWYqz6oQ1SyO8kwou9XNTxZgY2/Lo6cywfi/MDFqu7g
eDMb7g2F06mw3oxJBx80LdCFMeqHDXIzlZA6KqGEhdOftIohWlu68n2WkGGMJ4Yz
29KHteKNAi73YrK+w4exHOlq/U5s+xKLVg/3k8QFKdVovfxbV9FhgcN6AQjvYUQt
ckV/LzqHAj5c1AoShZDBg3fzKsfjRrlYqDQI87HryJwQQSdgaF11fU92G2ys14rA
15H09tch7Ox81nKs6BPnTRMVvDlFMNM8BtnDKtlrUVGwPDHF0oQOCPqASKSD4dHQ
8+w3fvhwpToVcRLttg+eVY0r9zPtUgOd54EZ+DQ7jrP3T4XnPalOZMjvOgmIiwO0
wJIHAv7V9/wlky55BALHIiGNhFIRYqZF8mWnM/ELsJjlq9yG1j1n+smMTTEx+Wbv
+dciXVbyARoMgg3cfzD4OIFm9/smU1qWyJ9mUzF3nBz8acub8tc7aFQBGpF35g/a
kj2942WqNogTi4lQXlO2drqPWglxRgfskun2ht2h8kwiv7k0GFNxcqRMoIuqMA4o
XShlyOffdQ5I6zs1hCuLVbSf56ilBWzS5QfBFORsJ5jLkibY2t0BLRDQPotQ7a4c
C+WQl4iOzkGiFa8rskez8gVCAB6pY4gApL6t/bX+HNQD2xZAwvcZ+ouBnjtozunR
9Lkg+Xilwwb0qPRJe3csmKorKsR9RTCTaNzYvEPyw0QV40J8wGOI0mdPsn6jvSl3
i4qCUifQ2jlffT2ENE4ENQ6BRle1tbiwplUHy+ruwwTTiunee9dObrgnMpHmH4r5
8OrGQ1vH41sbu1AetN2XAdg/nZSV9ycsp0UpEY0oGVetg+6xsCWZpOjMq+wawtb+
IxRVaOGz92Gwt/xVioG1OIKtfpjyGNXYEXLiqD/wfgDTWVi37WptApPHa17nJluv
+3IJzXyGW74z4lhiRkrILIbAFHZHpiNfhymDC4AzlI9zfKRpemjoJdigp3mjaON3
gEHFnD+PfYGrvYLppTcFrT25K7LoDZz2UDyse71V9MUIZrjyBj39cob7OKrygSCp
K+c9fDj03HDry/fLZrzOXqmNfOweS+REH8ijq3Cl708o2yZGqP48howF9JmMYUyD
TJUm5YmknJk0GvYToNrwvqnhvi11PS+EuAlHVG9IsTykYPEMLuYrP2x6qemsNCDG
v24Isz8c2OOBh7yNVjT6mAz2KL2WjIqePt9800zuqaTOvpLxGoFWR4JFeMfqEJ3V
g+dw1Iyr7ygn6sqej9xeQ0CrDRkwLqOkBmUXd2oZBDFZS6/IvpqyhrT3Qg52Qzsc
viT133LSlB0PM31ZY6oXOV+Uaprfb+sFws9cJoZ7XEu0bijAEbN8sKOPAkSHpUOt
Y8jCXcDZdDgGhjHBm1c8buDL+XiDAbjJbyCU4qLHuFAMTM2CbtXe3SITaZTYqn8A
59Xdp4wI7+uc9XAIsWNqEgIhOno1XERLS7HnHKauYsul9uio/eGwHOTOwl3/Ptey
P5ZcG6C3rzns+CGjZR4gF3uy4bfq45xWbbh8dDO1XQfbHjMqq380Gi6bz57pSIj0
HhmFF+RylQnm0G/O/lCU+1lzKLiXr7TjviQN6yZxqMP/6RtnrjfRKYFEW1RRBXFW
VAJ4Hl+oCcrpG2hQA7o2DOmhQUlUDMNwPFqp/6RFT/bLm77rX1oqRPYtheMjA0/j
POThTzXejLOfhMdHwuvSiLaAVUEQgqV/B7bOaNnBf2AUeZLCD/ALN3n2u98pivyw
nD7cgakolqRkMVGBgSSDtx/H9Umas8oJdJyuP/HjmSBsjKEFg2lj1A7IF/KZlwwp
W0ll1iccxVW5Bc0S51gNUDPQ1PY/OAphgGJeeXSRTq0/aIvYbd8JtQKCjAhXSW4B
bhsLzsFLfqtF+kYSY4T9dJRfUpCFQfNY4Jix8Xtw06oXOpGexoHG2tUliHDtOTEm
XVw6IPbVreHA33gghMTiSRXaapaDXf5iFBwiPjV67iwNRnA627zTDptgYGkl5ubH
SjBFlrnMignaq2Kz1bq6FzaOtQ7gJg7QKmJDXDYkG3CHOuITyDgWvfYY4TgY159U
b0w1w+mD0Wbe1AKPkODIxJPGwQbenRzjMKjoG1TxevvqjaeILnf9EMhBY/jyfiI+
ezHlirfGcWrNEswBvmGJckufegtWGJF0rJ08t2Qa1XnAl2B5EBCrP/PYkBORU7nb
ulmaurjX45Z7SvmQbeOzIcCIhi3GijxcJ6oCTnp6P4pRr69J2oDP2oA1AGrL7G94
oXw6uclvTicE75CxO/rjQRJFwOAtXlAFbIi1NYtefpeCGZ0QvoV1HMVL75IyyvCM
DBwG/POyAAu8BbtolySWIxJABgzGyenDKFQPd51q/+FYicbjcW7kcOy2a/b0N9M/
rQcQqiMK1wkjF+nuLcsZL1XVIL6A6ut3xUa1j5hvIYLf79d20vNAZcyXMlEMnKhk
+0C/8liXHZwFfBR9owOXED86YXxZrdUBk+pqNYOfX0VVg0Qf9LQGVzOdwMtVFiZy
k/Xsl27rLz/4zfQK1oXK0zGeS1y/eFGrBSmxPA7In6AWefWgXprd9aag4tRQxeL/
sotfDT4BDubXkAdlB4NyFj5sJQGYkL325+KNxNASSYnV9FEBxKxuHvnY58UWmP9j
vATHMfRAscDmDXQBJaR7Tx8/QCp4MNvtfvv85XR2XlZ+nFh3kEYhwWb93NlgCLuP
+jTGJa3EpaMKjNDQIoPMJ/U+nWLcYPoe+RBevsUuEo4KZaZZ22L83S0cNREydEHD
3dc0NE+gyosZn06uTsl88xIFzQ4C+R/QAOHqH3eNRMnOix2pfDGtph61CDmUiMMv
PJ+KIY+KDzXXse2q6t6bfcmeX4ZgaK/44Jc40COkVR/NeKqmIah4IrC8DobQhjnl
e49wZUsrs6r6frZI0KEpRQp2G1mOphEi3NskzFcG2p2ftjDbQqgzNsT6vm6fF+ZY
tTzAvfWs/qkKLvPO0w/3b/FCkaQrP1cxWLOY0Idu2T3yQXFm3kYrkaTc5ch2JhPW
HKSG+zWHmxuzT4r+6x6qqelJgZ+z8bJSAPp3g4y9/mCIzsmfeBXqkzjSDHXux8AT
w/lUNZRgiiFHdVRDJ2GdXdj9b475FJ9o3a+M40exE6YtRzi2ZIZbdT9QMyMaa2uV
3SISA0vYb+mbM5Xnns8tPjRTyTcZLI6/uC9W9uTzuDAVhfnPZVQlevpWmgzE7689
nUzE251BzVKhJamtKjtUS9b1t2yPm5y4S1auJK/vnoxwndQSettxrcKC9F3GB7z8
15xJg5pbxMHslbIbclSpIwjVEsM8wOoi8XFQ3ykV3pg+Q6iAodGBSZeMCdGxRXkR
dbnKmuirZOEOL/v9p1fcTiojl6LzrWIZ6ZxEMviRkVSeafVERdY2jNCEgBz9Q57u
Q2JLTelTr4EzC+aRwPf0YHv32sikJcn//zEhjtY7nT+p6MI4XrJyiWSFYDKOlh0E
LksvsPmBxyd7kyAnvYxsZ6YGVvl/xhuHKfshnGmIr44Vy21x6slFUwIJ49a3vsMq
8ktzUsux4ARfn9OGzpleA/ENBWuNX49/Egxf1b1RylnYNQ9iH+g4vFMwhENeNl2Q
LdEc1Pdin9nfnJDvjAmUtuZnBE0Uq/a5p0qf2w+oEg44jy0OUWCnEpqfeWFgCzSp
IObWV3Z35NeX2aZqMPu3wWQP1T8ekJtGfivIvcJg+tCy1Sx2yX//O+ex69NAHgch
gZD80v2tizkZQhrnpH9RSeRGJ+pk2YnOBrc6dvKLepPiyT4o36p33LicMC3WxkOy
5zkp08oGBcKg2lJlEu+yGSdtPDS+qMsd+9mw1BPHXSL5PYCSpJEuAh2ETotPYrRU
bgQrVmLK7GJlFSUalklbrBFfXicp21ohHzI+oDmNHgDRYJvi4Uqp/26uNrZ9xMqC
tTL6fa+P4PMXBbYz0xxXPBStQAfa89/aKdbK+JhvUUUs355LqNUD+/bb8DimT9Do
B8GmRjdZSdaMKHkpjoDOF0irsSfq6tJ2lek8tBek1gMZDJG4xtCyAkdm2VHSQnrY
9F84X8riDv0lIAHlGDxdCFcJlKarkk9kunrYOZv9VOqokAOHrZt/nF3Xy2Lz3LeP
Xx4fPkV3mtDaHssC19WzFsau3VfY6dRTLBDZ5/VGIbcxhBe5RLZAXQ1ZkfSgqN9S
U5D32xoIyaXH+1MpR/2Lliv5d4qLHNDzZuDvNxRXjzfAc4xf7ixxpz5Mb01Lg49l
HNVMilkwICEymNeDMq+vugxzYOEs9gbs+veUQjMO0P0tY3QBOkW9jUCGvf/w6EkC
/ieu8PHEPSvIEX4XRGDXsRqEMTSIKcL9Fr3rFScNuoslFIS9rHYUBvgIg5aqRVq0
AoPXYUdpxIWQsnL6JGzVzxtw1cIvASRt5CUWDTQhX+7AX1UGMs6+R8y/T7JjVy6g
aqAVPzQCKDhdqhHiD/sl/UVfaKF6HAtDj0tVvr8+I0ICO4DJYSgB7xJLfVDZo13s
8j1t8XsnPT/Ap/Shpd9iB5rombpfA2ViGO4EKWh/dIrIbsZU+pRnnyBctcTnAYlh
V5TUyNrvuvND1G6Ug9FPVIw9wufpUXFqDI4daLx+vUOE+BcilOx73jmxKqhJH3aj
eZW6OB7MgwkJUFgmr9zw31w6hIugP6+bWO3MlitrPzPVm/NHePZPp6g34n1LOE5v
JCSh3YXXlYPZPdJ4VQFMBRhmE2bTFE8kOSj0mt16byw5oHXiVHNACQlxpjOH9Sa2
Va3t11D+ziFsohPXkLJBURyADW3mwIEYYH6hOuy6sndKlyZvIOUbLUc9s6r8swyq
GFuoKtLVw2+GZSyb/RG3n5MaRghGJRnLttRb4Vd4+m/4TQIHAWxr3PPd3vitovH+
18U7xnEZLDrhbgABjIJIMOqcEwE/5orABRvyL8n8/KDXCTCe1/gFuyBdIMoEEQ8L
PSttIQJELCsi7wZxgLM/R+pNR953fC3yuD0pvVu7DXK/gkeayRq28gxCrrzdNAh3
yAi7M480liAJfX8RBWrVc46ewrXHrYIELtfnhoC/tMjzLcjwZliiTAcBFzg2IKPV
u8QX32u9oeFdBTIHI081Uxpd2b0f1C/DtX6dWG01a8PbMtt8+P/BLbUkSxL6+5C5
w4gMmXOQbLYY3n7ZpmlsLlRvvZP1slhOvPZxpnl8qfBD5kT6sZBjpM08NxG/sJKo
aWZe3woV1g3/O0ra4aTlVPMzZYyuaRUMrM7dAivhcubZjVL5ytm6+xdSROJFn7XF
BhnWfXY8hht/Je+In7mSmptH+y4KfHa9jMoPLhcv/L0kUQRPCgchoIXp+YaRpGSn
EXvfrixhK9Dw3ciklC9Xiuf8/2VWihFvw/2C8pja7jfptwxRX4iZewjHpIWRLPNu
44ACkwGsdhLdtamoZhBtu5H7JsL5Ra4Ci5HIDcuqJafDiImJlWoZxm3Esn3E9rNu
k5n8h4+PDyviGFyHkrGx/p9ihvAnEwDmPDHem3V1y+nYD8fsMGvILqxrS1V4O6zk
HkcKH99NwfsyHhPQcC6ErzKZ2oVVKI63vOS0FidSZhpptiAa0dyj+HL1hBBJsV0Z
Qw1y0wRCW7HRdf4DAgs5xVxXFXmTSdZWA4Z4oyuCv2lFCE4BEXkW/94r+4G2NhqQ
JJxHEE1BgGl4WeOSqZHiGNrR5+weu7KUb4v+nvYE0lsZb/IbFJCbH5gPYZ0IG9tg
0gS1AOrDLjvIRDbKRs+mu3kZNII+JEf6eVPjRMl5X5RmIR2avKKjX5hMvxG/TmG0
cmtoIv7k6woFmwotbpXhUBGVYrcgwjgqo9lgJafe+qQB8Y3z2hI8hPDJ2HJ3RrHo
IdpbSZpjx9ZnmxECuT/vXtc0xQrWnuRdkNquxFoFkpZtLqjXyLJepYg3kbR8Bxhs
gYJb181Du5xQrp6HsydE0+mfzCGnVaIHuWppdDwECobFfI5gXzzofAM4iHCWYU/x
vfT0fh5YAAOjY6DWTzRQSBuV+rQQy/BdVwFhJlMUSxwkauUiQhHSdnFjTa51qa8P
sTKJsI6iWlBkeoruThH5ErwDXcYTzX8J2x5TYi9p/0Zs+v1dKG2RurnnsOHJZKbx
8aLLM50Vdj5AXqWWOjfLAYkOTpGiLpTSeQKZwcDo6z6qPZ0NVsesQjF3sOStq0i5
AYrm4RIz6Iph6d4sCw3exuHSP0YS/bc2p9MyD751+dNjHOBrB17zj6aipT2s2a5Q
YnfUq/2T/P+vn1AS+2jS6o1DHD+9K0yMD0YEE+jkvnMz1i03tIMVNVnkyut2C5CL
0AziQ7bjnRerPlNylBsLv5flrYlaTzoJ+vR2zMswMv0YKnIJ8aMxECyMUZoPBRPP
qSXz/W5kjKmbm+0grHjv/MAhIlJyn39e+nzyaPgWfAxoXOWwOCCewsEWqo4NlAIb
rwixZoyIcbE5zz9qT12DncvTqZzNda2ZI+KhKJb/G2aya6QXZjMc3xZoLNDFEL1I
L6854JYDU2vyYo1ysTahlRhErFdbmU6e4Ez0iZbxEac789BDXX/Xn0/VOnxbrsBX
YVyjR8fG8hW95yLgOIpe0z9bK1pfriz6AUUyU47UIR8v/RNQTzPuayJdfQGen9Jt
rnwL1x2x8amU95nJnYsmUA1f+gAjFGp2jXmvLKH4Oety6X8n8IKXNLgI039Fblec
L6elA9Ew3Pl2didbG/n3rt+ybGKBf8q7GMpkf1gcENptHAP7P/DqJzJtnjIzeFdi
jW+xo37oKlTOCSmYhhoqXhFjwNITBaW7xxI95QotWk8RZdxkCE0oJvmD4QLq4LgK
Xm1tkNDqK8OBTjfWrx/ZZHrrr9K5z+u+5duF6KdHWVfRd22v9uf2vSlsIUD05S6B
MqK/2Bq44X+UP/kMD1584B8AyWUmGmTsfLMdBR5KG7SJVdLa9SuUkgJJJdo2I9H4
GSweW2WzpfAlCZw6oct6CwYRCAVY5+W35EI0vAoxWBAqgK/lSu8WztrgiPbjA7DS
Das4OU7tz+zXRKsXEesCwLhU0fIR8slbz/frkxBdM9+oskQiul1VV2TCTtqPlpYZ
cM2Rk9J01ZqMYeqe3nYWvIqtb8kYwAXJ8kVWhHLK0xQVqh5IdvaVpTaPzDcxkg+v
uoQU08YuljZ29BDvvlW9xswPaScxwQKJzN/Rr8uuXa+ZcImSqV1/gGn1x4n+1jrr
jir3SfPCSW1Mf7L3O3kQrIBLUxZ/w+UyXwSSJSOjD2HhYhcDf+GuF9HXbP1EMGL5
K+uxAEoJaJSFp+inWSqA3qw/vGG6g5DGZOqdfR+cLWf0IXMDpkEGkfGaYXnCCNKV
RCCrI9XF0PXu1dqrbV9GoGuPSiaa+UqpAFRNXtOq6YCUMTd5CCI04++ygA6tx0Bq
IBq1rig3TbQTbsR6Z9xKh734uj99IpS3xdrsdffGFLa+98AIY5rleDWFJFhIhZKZ
I2VHJlzKzQ0Zj4LDLDW5bPjIwv6LZC7iQptDJfUIYB6Sim8YxUbMR1vlAH3dVddK
X0MnpsVOoHnpgzkuhwInZAkIlbnIvnPCTOJaXmsOQZIuoIo4NwK39NXXSyEddTMe
h6+WSkFz9ihWXHQeVTBF8W6cpB/aFTtCp/Li6o97A7pJMjoCAw5K0QHsWWSRUVTu
A7ofuI1/VgetyKO6FSw3CY0Qzbs679MQYQ08KlOlX27i8F+0VdWg+UqmsSVIpxwN
ra/0QD2Fgy3QutGEk0bo43KR2BgeRRS+nPZnPeNdlogqT9gXh4v/zOEWFWtlS3A+
W4GztEytruluFXDeCNI4mifTwvzYFWqgKDs9wwDE9zueaqCiP/JLBWyDSyXve42Y
eLuWkUF7sHkBudpdMWe28T1nYZ71rXWoSipPf+khwDqsII0418ibCC89fAQVAxXx
aqiBns2JALN+x0u0VFllCSLq6/o4XLyb8wh6Cre5Ui4iFFGiSdbD1SXLJmYXcU5P
NJIOgD/gbHE5AI3NrVquWpzwH4H0FCq3RNW6Emx99MCDo5O5YoBTRxPyuRGXj6/V
SppBfBf9NZ2+PvN3XjJHPtief9Z9d57dv/IwBlOx+3sBt6LNX/93VnSotMxRuO3d
KRNWvWZU7RUPrOFJZu0vwTK42mRwePbTMyfpj7pnuU18kdO5Z2VCb5l5jSdc6KvF
vJcwiu1mql8Nhi1HhgJoTdvyuftETk/L/2vS8CrYZkGIcA7nnsQ40LLfaikFe4YE
h61w2cux6OwKKdVQkiQw2zh2JlGWJDii3bIJgPWKhf3D4SRRh0++tNExL7GvkElC
ek8KKzx1HduwbNKXPpxGB09ZuMQoiFYENPKb3qE0c5a2/ou/5Sz42fWKmNGu78Nc
WHdn9Fo/6O3n8BeCVHaQ5KDYY8LwLuay45Z6kLzFaxJK7aBS2VqK6kuxUUb4lwfi
6PVVgyHRXDP6zpSIIB2YhCDLwRZHaGqyBOx464bQmczufY8EGrcGcxNjkX1FJQ02
IF12JpNzCkpXuk2qDZ+cKlhXyWGYOwzHS4DIWItXEDC2HMmY+ZAIHXUItNs6SA0m
1UD0fSVtUo06HGxtmtls69NcZY3HERu/E8fZnBOiit6+zW2oewFYFEPIsJgCoVqY
Frp2gGCoBr0fh8dAgQUmS23fZ92xrfRgI+udHz6uouBmbg0yp9ZfC0VF/VNnFxBp
OT6gY/VbWmCheYp3ko8XEDk5cdpTmjUiBJ4IW1iKceHkkyrDuMBV+DCZTx3cOufv
vw6LpoL0tc5/mvAU618tWpiP4PUTBxnZoHThXjy/d4/sIUK4pchrOOdQl1GBxJ7W
cgz7KJYZXyLajBeR1RdIbg4JGSUoUBvaXPh0SxN67NGydMIRQyavyhGo8y9iI84M
lnJwKp8LEKUyp5omyuSX1ia85SZ8jiIF+vot8DFykM8WB9KzMu+wjM50lVEsmAov
kR7uGUGqlpQVGQyqhz/RZy4PK0AVyqoXtkr1HcVHHXFmMkRzsPKK8MetAq5b8RW+
cpP8H1uCZNLv5kkc5LJNS967jmOLULqrJaECxTz7967U6CpY+sy2siOtFgKPLS+B
qG812GU5XakpnD0kcoJ3E2ihHN6jfjsZEncQpPpmajEpsCjO5QlcM2B3HLXFCWbm
6xQgTAxWSpGVttXAXmWw5dUPCMQsYHgnJd4HtJfTuMWsSWCQFiPjZdnCZuBkb9hW
waeDqVrmjBRM+83Nw2Iupg7RKXPcpe8OMMTCqvOvTqymDhHoMBOVfquRWsofkU1k
97HjAU97ZpTLeiCgQSuCNQyofRGJGKK4xut2MBlV3SCIG7ZjZRc3O6HmusyLzqW0
gfUXran1L+semjB3Cra2Gl8uszPzQ/MkiN2eR8mluLbBzoudJ8OBxUK6Bo3oJI7W
1E51M2gDVB2WQ1QMnDuRZzFvZV93K0FXTLjikKr3PtNpk7fBzvZk/EevZ6cD5h3G
Nvk91WP+5IStgQy4laAlXvqcPVHUGVU6OmNmPb8FuULXvbyzmFu08I3vAkmxVLCx
our9tzzCnReiE8dBJfQGHuLjIO/SM8unISGHekMA8V0XB9Fptb2OA0Nh5iuUKInL
DfEQ1h88cX9eQxpfO0D+/4kkvCCcOlViwTutAEhWG+xKAQI7z38HzIsoHnBtE/RA
NPVCquGSzcZVSd3XayBNuimNvSm5WXzjkaNVMnRDrxQF0CnihF67bqM/5+drs0gS
VmIaXR7OVTIo7sQZKIUJuCCjuwMr6FDeVEOz3ktTrZUy012qA5jwVyH8uMH9FPyq
PJj83Jwrr2cxfJNlf/Fm1mkB7dMTlrNgDR4zTu6jSFMPFB2IoFN2UteyLJsRNmLP
l+wVu5dduVqt1/f95bMRRNyoK56NyGO+dVwH5CrAEc10edbeX7KJxqQ5hODt3ROD
yMb2NKnEIsNhH9S49Qcs0A4ylLRdx4Ho1feaOJpC28HWmDnJ4jLfKsFX/aUaS5ST
CcEXvxArTiF5EX27HxL/rdLgGCviGu1uh50gUNDCUmOyGuYuOYeMHfTIC2Sjyr1n
H1oezhqrZnClZvOTqyfZn+8aIDPlSHNVabwcuxRUXjwztxW0QeCK7girAHI3x9zt
7NxdpkpNDLMKh7TgeHc6mNOrcskWlu+IqDgjbEhiUhA9+UiWDO3ZjIfYMLYXSOFI
7KRtOHu/f14FKlGEsVaVbKBFpoKWSQXSoPpavdPCBA7yFhfiqFNOImfTbN6zXpui
GsMbWx76t4XdBCyXCOaSFo8sRSgCdqAq/3rxU6Lf/FCZFVPzjUq9Odado/qBwNfd
FYloxz4jlwjKKmvHXinK3Ah+qgCEcnXbF4SRt0kzP2E9MKUU5nuWwRefgjqM0Rpj
f1Br8ab5Ee6DvqHYrKtEFQ907EB+GEV+cO6uMBymWU3uWxc9O+5Ppc2pUAz0FMG9
4WHhs/+yihYw6dpyXZwT/wSP8JcKZpazGZwXXc9d4uUXr3H4+H10qTIxRx7nNH7P
a5XtA6ExIYWLGx8c1HhPEFp+C5n+I+bBFlWkVgRBISK5TdLY5fw+mmt8CdyQOif0
HFpYPSq/DEZfherp3g4TMZ2IPtd5zbtLQ+TuoXdKD9Z6/gemK++nD1W2nqOlKSqt
vsbUJPpFRCvhnIJTjSMKv+TWtGTxKMU4HowVOHkHsSvNCdX60REYdfEHDNtC0cdy
FrSA/i9xD5DndSm8AUsHZNbwyRL1zdkH3f653tI8ouJuL4sPGazcVQ1AtRVJEpLx
DWJn1lZnTfPFG8/7f+tSTY0A+vh8g5m764JNHH3I5GHlmoqcKBJSRqorSdybJyaG
Kz7WgubT3Zj2JOARHaqCqv2H/nXki8EeRpViG6D9NCxqlDHlMeXHaKRqA82LwCfg
eiX9pBbifeXoSlk2GEFBIKY2krnZyY3pDSjbVbpWEPSnkNYiKEAxNor1U7vR3ACO
fVNmYHqOtP/iYJ50Rss0nWcAK+M5BcneGc07mNjOC/sApAyDkQszmmuYmRODDnfv
WOKgdfpBUvy09deHAYnMaopUDhIET5WmSqaDZQRAKh4WjE3VMG3f/ZUEKuH6q6Or
V22CHfhkhbkNu9IJcT+vY6LvjR3bGvMfSS5RgZjXPQhBPR3d4F1ORn9wgoOI8+/b
zjsQeT0pwNBxRkIDCwwz7Vr5AWhPV7pnQWLHAogFNPOkTfxDX6bsiIXIbreJoupO
9TxnB45eTb0dSEnLPhJGrL44pNIxuC8tzKgypeSr2eSpkJHNUAiETfunHPb3AOaW
+X2egvLA27G5XdAT8gy+4YxLQz0TWmWPUAPhaSDHHOUjUa6EpODZQ+TAxLyWIGfS
Uz8nGj5KhptawKsb4Ose0RAOjUP4es46Mp8KCR7xni3CSGSufDeridX2k9bpCsiB
0aLkFf6pkmJ7ez0FNID3oaTl/hQnBmRy5QRz+nBam4JFL8ZHWPuKbVGwX3QkXkZZ
c3BKNdKqy9KnoQyIvYmHUQvorNnCj0a84nn7ZzRcFNQwIf3oCRBGeEJocmJnNgJQ
8REFH5XIVRvKSC37BQ/Vu2qwKeufuZhBBjnH2I7uCYwNW840Rxpzu7QC2EvGoDTJ
ZZe/rKpecIVHTZupqHaDayw1tmvl0sclJKf9j4pKJNoagfCR3580YPpKQjTlS43f
wRl0sSse8/4xTQ++eSz/IbsJqxUoRazh4rr8aHn23AjlaW5gAFRisQiFs0ZKCYQR
mXaQr5GIXv21lkquixhiyesYWA5UGb2PIGsTZCDl4YILqXTMhzdc/xZZT2V1HyUB
NrV0CpnUCjkBwgyjMkvHzHx+TThoeFGwaCNzUJnQbZB8gb9nYBiZGs/nqBihmxVi
YRmnQDY5LBEXlQJyTF57fFilzVcRsDRsE96vsK7vQT5v+T0RrxktRH0fGzefk/WK
U6h2TaLGIXLSg5RdnEYlXOolSzA7eDxYcf3ZSj0Wr7O0A1uTyvHgDDPWdMVHpDBm
YapNie3eHoq2zD9AQuU36qDmoa+uCe25R6JiCt43iN6cO9LdcWb5XS2T6hcym701
2CXxPaNvAJLGQ7Awx0OWsNQptLiiioucZiBZmodeQcWhJVgweJfm1b3qFK8mYxwz
vszz0iMFoEVD9JyAXk8I7KK3hP+lao16pXJey5xevsiNOumCmU+Pz3NtuaMHqQvU
TwlLJIosK3mNXYw5EaP/PGUDmcWT4OFDpSSG7aq4rB1nn7cw6JR88Dy3lk8niVwp
gJk2SlLYE5tJDaIRt9MVquni20+6wcNa48T4ONWibqgP3bP/kU9C34sxmQs9Wv5q
CFRnKK50yhGF4JQoQgdI3gVenGdefPRqclXY76cm8XVSj09QzWp8P1pgxAsjViNQ
//6dkaXfcGjZYtX+PEanWmbx9n9k6nWRBUg45m1VuOUfprvSssbZgY6Rb9fkNOuM
zIVdeKiM6HRX5lqQ5rBMsl0PIDgAy0HlLVhI5xYtx2fvOByW1nu0gbf0xMy67Fv/
AQiLzRYkdolxZpfqBD7SKhy9lIn33QYL4qtZfNIKmvRdi0lIEsFzidytoNEJJVU7
7Y6akzKChLBhCX6BIUPu37lcOeB4Enm8CaCxp0ns955EuzUjdH8D0diLRKaeM2fF
VDr7QdhDBKuu2sZBR6irM6Vd68yQP0Pm2SCnkSbmfwAnmnbf9vEKQFuxgGHti8nK
REaX7IQR7cnDHUeilbK7KHo7PelXnuMZH/RkLS13AfSwSh6sOEbLSFs13MLKrQQ9
Z59t01oZ8uP4tLytmFNiMek+qGkXd1c2OZWA1D0jhphqRZMbUlUOgPvQ5v8TP4nD
EqzQt1fdMLbc772XxAC/kOTqt30Ndz8Rh7ZgS2FgePJ0kQu1UxWqybQ27b65Ca30
ChR0Qz3+XijLwMtyZNcrlwjw944icKqIXladLopVSwuIRWamRW7vq5aeFmOyMgUJ
u1hhUvIoWoJ0vvcY8j31spfC9f9QrGX7wH90uDq6HtAhE9viQJ/pJCJgQYv2tK6y
woP2LiEud3vw+JgMfKJ5h2KAv/sYH4ycENfgbpJtjdUCHi18z0w0BfzKtBb3DWyu
n6V0IAWxg1vYdh1EtR73ib39ovoT0EnZf46Mqx4IuI8anfHpvPLQh6KGt1ckvB6w
JlTNB9pFqrQh5JcNipmf9sAnO5HvE40Oze23oFJRpgnQyZG+2mB86is7GEghFWsc
mXNSf6KAmpALs8gFUfjwSSIp2g04a8wXTCl6J4QZzgx4Cg38GtHSa+oSBE3r8DZg
Vq14A23l8k38Acx19APIC3hQCX5NBqS+a34L+a5pUpNbMXU2oWaKk/4V9ese0NiJ
Rv5NNtE1gd6GiraVLFeGyk82kbzdudyTDlQB3G7mrbGrYMH0jx3//FN9ZkVnSHFz
WBf+yBqzbJONhfY3v8XvIs9wCRoG5NkOX5/2Pk7cuD7Bg/KMjfrwDVL4u8VcX/UA
1F+vh5M5j1o8EouvUKQKEEsGMuc1wFOOHg8vXpw8Rms6pHBbJkLNFA8dd2B+MEh7
2YRqY+S7E0yTVwBCJJiV3JEI9RtDzp5a4fKD/EZKU1n6798SAvINh1qKZJKezUGz
7Zwc8WaoOgxd6aT/qzUMdBrMse9GoRq4y2ji+NWbkdlPUI0Jw66+/+Bx2W/6NtJd
A3eLoqdXKEXKErAoiixKH0T6tgpRxhL9Nu+h3Yq9rnb3CNY4H9wusZ4TFoAAhLxW
6wU83Dd4mZA+rR/x9QyouujxkIEs4LydYmLtfCXbMxuB6LER6Awl3T7/ppUwlZLS
AgH+St/t3GrtaNei2/IoKnSOYqVaaXQxxAQBTOVctImyMVDzh6WU+sUnZiwgaoHG
VUCd5RxPsJ+cCxOp9qTDElVQKLSNOj7z+EHXF9swMC2Vv2l1Wd767rPnXhDnlzvW
qWb8nizjSsz6yXHoPKU+OILHkAFecAcatvv3a4zA9JKqJNRUKwCl5nUNg2OEzusR
YHes6SNvbVs78IZ903mwOZrXGFMo4RwTjph3cLyMGq2dC1IRhzfH0d6BIsZnTMu3
bzLZ2Spi2phFlIyhGz2TssTuqt6OAnRleZNAlCzzHI3HDbIfe6G21c3aAJ6v260k
Fb7I7j9aHfSiG74vfjvi8Px2PgzkHGMBa0sNl0RXtiOxR4O1z/z8km53CmdeMQ8U
eQNWdLZtx062UpS1eWbXuuSy6DKhpF8fFg4uvMemZsAPg3RCBGQHBUJp2L1sJSva
gu1/NtNWuHwkk0uVkvod3mC9dBwFzktXKEHGZN5ySNJTlYZDM4aQkyv7cGOyC0IO
7eyUx2bs9ICUvnbMyyMnHfjyEk/HOruYW3LVDJgXfHswuHnRBQilIr3fcU9jO8ld
dHeewM0CR6lhca/AD0hCcG1L446XQIH9uQMdfHMfrDEb9kavclkVH7IHwA2AGovv
uPMVErRxkS2SOuSxZKlalvG94Gy/zMv7c1Waj5eMH/okOGOTV+LHd1uboZQGXEDd
9UZlY+WpedGCAqm/fe8x4aMP21ohYgOWZNDmh8TXlddlHQgvcWuIrEaIZaCDWZOr
6/Knt+HbmKz299gLAuBiboupxH0vTZoU4Q8jO68UXvKTclROpWack4bt1WnFmymP
jtgVhaVyOlPcb7QTU9+ax4giZiNu7To6CDIQmzsfh0ULSi+u44atxqkOyX1l86sj
Hazz2RKY7uyKxzDjBb3uvrVeLWhYuCjHZF6JBWV6hExnqaoh8Fm3hzYoibdhZj3J
aCkdDhahitngC1Y9olASuVIytwmatRM4x0x+fpCMD8v3jg2JSkjXEwRYf4u7AdB9
oJ58sNcT2kDzZSVQcQC0R3o+6L1a9U+oG3OH4bwOEndRTH4HyicAMdVlO1nfvkyX
hNf4p/+GlrIWp7+QsvXZIVylVrmCOlG1XEbP8WoPA6fzgo7NSySQyijd5FQ5UrUk
ut83GbEG2pv9E2P+Rw6L8N2tiBBNPaXM9B6rMWOLeRRkalK07zRh5Ren3mJVHLHY
ndBo2Y0pX3a0Sqab+2ag6WrpKspJvNduqQCUql2IVO6W3dDAOiCkzsFphSnjwIU4
Y/8wTG0j5PM+ntjpZRkntp2ETnywrrkg/KP7cxnIinUULko/BQwAiSqHv1LNGPNk
qLBBkBCNqUfktKPHHUQ7pcnjy1SoK5xAOGNkwOk/2TyE3IoCeJqML3n8D055WSSi
zB1puLyMEG1VcekPfzklTqSgYM2X+MRO0UBt8+/SPAQtxIFXNJaFp9F+awsr/8P1
Lq+xDfrAhucQ5AuWxPmj9ZLlaAXyRYx0w4kqetAF2rW2eAZmsidCy61N2TSvuMXH
u96sRzgkCHaDYAREY4c+uF/fOBsaVG4kDRTKoTmOA8Hvb4z8asYiJaMLh5X/d9VP
IObeI6zHLYtePLSDCwuH5Rkuu0F1AZcBwRADCu9KG1T4O/VIH+ZuCidUM/tOn4Sy
bh9ReVCiGsQt4a9WtPqInC3/MlXcgbrZ+mW4GjbhZWWzS3QmyxL2LRyT4c8GQfU4
A5iO/8FpvEABAb/FpwhYlEw3+0ftTpiUPzfqGTLuNbye6Z+XUIFelq7RY5ZpQryS
g81f4zsSIk4oJO1szOZWlIHx/0HtaSkcCwEFlhv0CM1G/PQLTvSZv1NnGPg/69oS
ZJRinJ2ligZLRelxezgTVqkgzdvTtQThXowZNmjs0noSQzHptZNwWQU3IxGXd5Ji
8vh5r/elol8YAwnZOpCjzVWF2XOjh1EUXHCy00B7LW5MyhBnRJoHmaYZ1Lbqi4oi
mkdGvTLS4I0XcJzU5WY1OzLll6+iMn+y4sBcJzvKb2urHzIfrFeksUjU1q1VDavU
CcYH44tkGOjL091YbZLPFjekXU3a0dD0aw/Zt7Tv9VMzlg5T9HPa7/12y26fL0cE
IEeTEpmB8zd3HDklpX8nOHWY2v5d8CFpqx0QEFeC3EqowOd96wCjsrXGfR5lux+B
FDLfQdH93hkpGmYxVAOVuwFXrmwnuBFvfyeOLrvvof8eLl0uShQqnPj9uPXUbVNw
WKpfi+zTRspCAQqiyJzZeedOLGwBof1VXtNTHKJexV9K8O9tsTFfvSwCKxzUHCJ0
5Y6XHu0yM4NrfEDYG8t6nnzLkMA5lkNnCoeOKfyFVPFfrAwc2E6+MSn1r5+fmXPL
83YR6QmYck3+sVHHPl29eCVz9nEj93dnIQ+MjVmnnkziCtkk8uizyZMsrICXk/fH
eNqnUWla8KUqL+cYBVzGJkCLowJm60D8mKlzIrbtZ+/1PtET47hsBLArgfXYwYSH
7edIy+puxFRvxLvfBPxRUdkpbLvQE02D6kH9rIRClHd6Xxb65NHMux0Lx0ZYxzCk
jJLr/0uHyOpWFTah5lNgJQXgIPr9Jm5GZIWWHlG5idPA3nYRZdgA6sj6XoJkhDip
SyAO9l8peJ9i65Kd/RW9KhNZfhiMh88NAVr3RJINc0Q5GgdlhI8NOZJyKlGoQp54
kWcIlycXMQ3odbyU2NwQVC9N0jrqCei8fiAkmaxZUEh2SluUYfCDXvrsl6Gb9uW7
9OiUhZtpGhRc4AafN2VH0usRsDO2kCI/rqtHf95syXejC/mfRxAqx7tTgSKfSUNV
2JBM/U4bV4yvvM2GlozDfRgfP8uaZfZVpcDvXch/tvHW6UtltJSX9ojTj9T/Wj3b
tOPLxnGfmt3ljED8dUpVMBcmc3iwnPsrV+GJ4aNP1R1VzLyJyh0QXcdgQ/cD32qb
rN1OwRKMneCY2gADTMj04zkuMpdTQYlKvEkaBlG5OaMssUCD+7EmeL0s3KOoHop/
v/2XgpLi40H3j/1Pq8wx7Qu6MGGHX006hvvpSYV/v2MfIC2oathtzqvNnE2NCHPn
Y50g/PbB5fCol+wdcKulPHRB8fhdthYaigdVQZBEDLP2ABOUF2OYfnssKip91r/i
x0Wue3/MGMQh6GmKSwbWjO+KhtrtmIVk9yi7vjOaGFMwN1kQTDOkg8Lugp5Uzz+A
5RoLt2W9xQ0gs0bDbgR4o72qPDtQ698iGti/5BXBhkUfXKO2s3x00a0jJIzsk7jF
d3DpJIbAqe7qJyHI65RzuDI2HoqK05TQRVfqpmUZdNjye17d9mFYxy4idmTMUi++
xH3sNYL1tfndQGIfuGGtqumOmLYjszqdqLRA002OkFFYgrROTambWuI50U0jS+tU
uub+2LhGKz9054Gy5bradwvRCW76INN9u24LIA3HtOAyICweq8I/AOZlkUxIZzxf
ktUzyu3qabkrODFQC1xx+a1FzaD+NHjoTMuFIf1rcYJg3bmjyY+13LBBS2Nk0LQP
uU/sGkLlN2WcDkVDf8IsgXz9ZHYFrrATOz6eaZCBQXHTdVzW5vU1enVCoPzSZGkZ
I8dcn1ZOVTXH0ufy7wMzwZ2yXePfdHvs2DexgjMV3WqKKueoY3jA98rfg8df227r
cs5Wn1pOGK1XVz2AvPNptmyDFL4FBP5Xrr1Hk9XEtEgnsqtUEhypO0I+/0wu+G9y
9g2cMbh3TseMTakH3JWYVfc6lbks21VKIS3XnU2KxKARjBEbyiiRHJXu8v/fTaks
5XBNyYOhOS+YQXuU0ekxotGJaYkH7As11UJzgTbM5EgtktOYjybXuxZb3DPRl5j1
mTYbqM5GFmQjnak3lEiWgHe8pxLrGrE2nAB25FgSI/JHjm8vhD74wk3EWI9xEFmz
TptbEqCjCMcfU9ojLh0wn5mF8wEpF4Ac4VFEFOL5waJ6WSmOyUfrmo7Pmg4AscK+
Bf5Jcl3VfmDhoDUd8VlTj7Kte3G3Gv7JRZKgFtIKzJMhF460IVvOVHkCS0o83Wed
jrieRi0eROw69h93pLFzs1SBhdHU8HvCjfznHmL2TNkhkvNSV2flq0eZllu8gYiX
mXGpCCok+7eRmG4IWCYM+il8fPNHYzl4fPSr9oRBc2PE0/ejG9LR8sMK33XD7Fcu
8xZQJOK8g3mqV7ojhfP+BMuq7kIxle3/G+YC//CtUEMqtaNuQOCkaR+tn5aNy8Ll
c+2mnQtG5ifrqvfhJ7RjGzszOCInogcA2bzSG3Ur9t2d5cUKfNvL63N3+7qTr1PI
XRHXeXs6ZKOPWqZozhxqLQUjvADabWaKzCNB5MdqbvFOk8m+TE2RwtzANnymFV0M
EED9N+ymwvS7mX2JeD1Vlxnz7iGoW+MeaU1BTcT9UmYqeigZGH1Kym3pQ4q6Oeys
qs9coE+jXAWBFSMoKPdd7Le7JnwFHyx5dPssNhbbxNSoCXcpLE1EzMHYyytHdvSs
m6lnVST9aY9px6KAjg9U8u6kpttXB/opTNHmqJd5uG6gAwCzySj6KatyKYB42Qsl
LCt0R5NOKbuz4onUZzDSPlI0l+Cw83cOyaDt3i8Ee7OyeMTLWRGdvH33uNCo2eCb
YWoCP8T2qY41dVxEXMlAA8B7Bvm1y2pCwp8MbXxpRJz+xOO+jGr6LqD5oq8RnYvq
X9ysjG8yyx3Il9eBjyNYA+Ej7wLJTaANAyx1zhMGzXdzxOgvHcw/x/lzR6crOeTZ
rejmCNFSQdk2VU5vRp9GvX0VD4IuFkEPucFig+wrBnSxOl0jVaCgTuI4sSOMq7QL
8ofoP7wIOhYFlBH64O9InWBFnNeXtvOEVma6E7XcO5QEIa/V+Cj8l6fJWmYfsRsu
Sngndo+xeqbwJwNtI+UtLkezgUJuHrQC0znnicgZGtQ4xBPpo4iFc+a3/z/cf9IV
3mrYCapkWKOPYPZQTrNkiyhbSTcJMYkKyIZybEED1A0NkEVXHAZq7Rp84SfNdcUL
+hE3/iM5Vej3ZO8zisKBRvPkFBwsQzHULzVCPLOeQNjscZGhTt4Ic5ThUfyAr7wC
SrwoZby6hhMc0MAwLjyVN0eICo0j568ONvJUniFtSnC/2AckOTOEu8wx3cwtFtjI
OWOmK4SIngvTR9Xf/lNrEgZV6ovnqIYN4lk2PtYwVDVTVeHxMHdI+km40Iczwjgl
Qe3GSGjkhdEnyMUY21NgqCi5ylLMWlbxARXKSWNsPMnw1Uz4rt5oVS2/DJOr/9KS
qMuUWzFG74opZ02tAdsrhs1LujUYojXbAj4WpDsO7UOpd4OkD/fHhNHrFM51Ekc4
rzCUHTUbKH9lD9F992xaykBaqdG2w/Fx6CMZyBLnLLiQcu2KzuRkR7fO6AZO54Yj
wIfA7Imcrxcsc7NRe1ZYqgbOpP+8+OwDN5bddWYTRywTucHD/wl/7ApMnMzbL06l
c4M4suxhzGumowFy3HV4lvy9aZBWIe0p5K5RIpMYDdeT9Pc2cfxD5F+dh+cFQrvO
AOzBWay0chaS9vIqiMPta4yadsmpuUVGNlqQZU+5qbxjNZv77MqyJZ9PL/7o/NH3
H5ltWA3qY1s031WpoWhNlVAbXQTlOIWmmG7XgtGoojBPqlsA4wie+7ga+t1KsfVT
QvM3nvKbwG5VWkAKa2kkG+/cOKKZadwfb6haErbAxpI6xQ6UKMvSyLc2/YXh1RFx
0Ftt7cJ+1dIEzBGcPsIAOYEU6RhamuoyoePz9AJA3gyf0UHSqxGjsdw3kUIq5oKE
T+DaVfjmm+eHUMfM+/FIiMPE3CisEi3DPxMWcRC88OMIY4PKjNHo7IZt9dGSPGOC
qsoIsdtSiRgLwmi2OEOVasycLOCNu6XHtUToOntwGEAzGEazEkILkWtdZIl2XgI6
BGeDaQ+zpbc1edbpjXVviPAYUJFsW0difTP51/jYWWj5xMv7rboJFp5kUCq9aRTx
HaCFx8hpHB77xjxZxSkJCYdH+TLrYM2KSopU5Vc27t/Az5JjnBPGjIBnoVV4ku8P
+AWqv8Gvqs5tvViY0DiVIx7djx7dS/osgg/rdkUtdxqKznP53dnmMNZGqF+wz+30
M0nBigI2CIeJ9RLv1SGWYAZxWhBzkT2rDx2FHuOofJDXhuiVfpn0smf6cda4pphe
Z4if1lbzrcFpLZkvMKJ0V38p1zCfbXbT66jSJGMvYKwMcf0mssRhuFy2tqN5eF7I
TfCg2KTTcW4ZykWJcasTSF2AvUKB8coVMDrops8LPLVoUjphajzBgB2UQs7bEhEf
5uSZSOnJ0BbmN0Oh2bW5iTMak+Hc5bFKT30i6mFP/5PBM6F2UK6NaefI5tbUvUUm
V2zK3PVNHmt/d0GbFCD5ep21+OGCDBqJQFQbAAdfrMHKQ62TiUCy5u3KexUA+aHF
kNAxn3+4EREn0l3crnRkbagJJ3bH0niNeEhv176GVOWqHVDYsDPov70hByr4HLZG
GTtWrbB8x7KcuKBBPtNMGgnk9BQD2Rdv+YY5JQ/mxc2EPRXG5aQYqE0pBEbnpEfG
1ltGcE6WD5fzawTRTp1HoAIs7xW8BbuSJWjiyCTa5k+BMuAyfDbzfNiREbiNgPAj
4wW1P8YxY2JhsPhDvSD0I0Ykh0KEgaqsQIxIkyTTZrPLbp9OAEeA5mc5ia5imCHA
f/5keGZT7OSxfeTgnETfbOhL7WSZpERG+OIY7SOiFUiRGWIJTQ24nDhQhVWCukOg
2zmatI1TQUMCgYObwJag1dxr6+yK7heoi+JtkLItVn1YSf/uLMkSqe+qLX4dVDHz
5aFSDryx+T+hKPGLxidxyQcVn+IAoy+K+QgrX8u9SJKAGN6B6g3UTcQo9A/dDYQ2
F9Ar8sERly9z0Qqzfu4uC6XFAPhRQePKc+So/OFTBYWS8nHq0OGL7jqJvn209Mip
in0u7SANzD+507qx0c6dp5Alv/RWxeJ70kHuhEPaxzl5XcH5Rx0IzGoW4L0u9JSC
gFruaR1JtrUclPFZibULSOQY0DlvaJ0RuO/0QLiBeTwy/dUjpak9zIL1F2GXCUgl
s1h5E6MZNItBP1kmFuYOxoVQ8c8YZUxF3vC9PeIJZM8qxupSq8YXjGS3/M8fekpY
FTXQnvbvnr0+OTdyK1yckvUTKCcJePWRlxiDrh/mp2vPi6uTe7RYKBcFGrWM+Jev
rOznxh7NTAzw+Ai4adEqOz7Cy4BtpOOYZhrjS045ETmZ6r0Z2jekb5nuMGbA7s2j
XiH+ksuEpPWD8gHlmeMS0mvY1QAT9SrIppwv4zJwf/LJoijuba527zKYiD5ww55R
ia6YeTCDX/4o4MeRuqOXKwD5RwC0dZ+ePZtCcMD9U07wM4hxgSkRWnYjsU/ES3wZ
qTgo1XAkPpe2THNBY/p/41Mw/pH+AssmyEgnVzXfP5KXQdSDXqp8kqmkP4HkjgEC
HRxYQxvSHY+zGUr2INGpLz49+kHLWvAes7Q1jbrcipwOKHfnfsgnfuLV9rcprHMi
VJ8AQ+AkNDHFnigWk6wbqID7Yr0o2LDP1oq04Tf32eY4oEY6qpbC9kNmoA+SiK8G
g3OKzMdHpYut+RGhsL+ia81OqBGHyMpcm0i/rgTd3dwER8smfr0hfOUL/qWW4phI
o3LHPtjduNsAFwtDq+pPzSkkKItNqMQwAkokWxagjjnLccl+Ptpt7p8WMTyPSKkZ
/hatPPYXobi74Uidfv1k5WzmvXLeiDQrJR4RI8m77v7hwT8iMImWuvbGrQo4vhD2
r3m17M3/z+DVRxF8/08WgngnAG38TXw5gDV2wA43ewAn2+wMLW79msKAIlYeMe4w
wsj0Mz3rk2qKItUN+zrxmmQOx1eKPHR6W2ZmhM4VlFcukuRi61IzzTIiRfYZF0Nu
qvNMGFsb6tksHH1XTP2etcicUt4VA3s8LX8TYtmDj8YMvJzsH/kVc6QWngLCgKYJ
X2eYlit8UHVmMVTNzLt7R2wqDDw5pNatU4nwv8Nf+FudvCcvUkls+UIYs1CLBGfu
zF+yjr5rRQGzbt3m77Ro/TkPLQLjpib0b6fQGa2uLB63RnzOaaC55wKQRq4HpT1r
9Yiy0+gtYrKCq8ICSYfhg/gaf5onj8HeBHcDdeAC6jG+7UYxxUDEuAvm1vaRIsbk
r6RTe7iqqBxWv/HOllCdD9yRD7kKsbsRey17hlnB56dK8zXx9BrphEKELfQV70ZJ
f2f6+HrKEVMjIYtU4UKrhgEHxcihey9WvP0C4MNss9e9rWEZqjfR5IMXQ8s5r4eN
hdKXNRXZf8kakaPDYv1m0E0t6Ft2m6kJLxx/CgYTl7lGXDAW/JETHkVkdp16EaB/
F5T39acaHDXRmySKWJ9XkBXH/reLT0GAsJpgGY3UHMdE6RuEpNAJTBQkrKz4IPak
1ksdpCufQe8Oi/8K/cmbdEbgb9et8wHejan3nAn2N+CaR61CX6luCo+8P/ZFO54I
3eoDDPUZQcjI9YsZ+Y2ioekGA4v0HKozSuZ4RB6yUvrIfB0Wn6rc05S59W7HNUjO
GhNyp+DckCaiwFc0padP9TVKZT6/45Ib9HKcvGdIAuHWCz8PJ27BylVGR39CLHaW
eP8F/Q9RxOWNEAh76c9zrEaosV8DZvn+7FYGuZiSQzuHWcCiKDE9JvS6j9P2HUzL
F/6JDczmXuMiWbhgTPZhZXGfGkiHVwNRJXjDAzZZImwZOjwSvpR2UZpJ7KpIJFfP
guflhaBYPoPoLrOdZYzyKQWWjx+PTMQpfXIgrYduy/QNCJ3xlk1YxMgv0lp+tYQx
Px64hJCPTk/HRK3oILjhB2wxzltOcqfMEm+jCJO6rQ+2WsIJSQUTLN7RZUmM54nA
MPWVd7mh2KbZ1AlQqxn5TNtptw4wqh+Kt4xTaHGp5IbcjXusdVdYRPl/jvReVwqZ
XggSvIL8O6FK13eykT5l8Sv1/lIdgRhF5UnPTYYa0aIIGn9AXb5wMPRHojxvIVNS
CfjnPccEpZsF40Cy2duIMQIKuXxEJNNRB75tuXKfCFsWgD5kM0acx4L3xNHMCcqp
CVguPqz0V5eP+VbM85QaPZUNE9Jo90ythaZI4V1cesELtMO38v4+kDI/Pnjzicbc
PEKn3MPCMrT4tiNNQw2TmY0TBbdaWh6LwRbkpApALvAScmAWX+IADE0xFbBSLMkV
bY3X94xs4jLxRLfiF4Mn+qDTqR90kG404ylW9GjV4VTUA6ZWk3kdoRCdQPFwdkMc
mw7zO9/Z9JgQ37voD0umCXErLU91lq9eoggKqX9nUIFsO668l1CpsN/39qZR6Lnk
pAssdo8eGStlfqpLQvu8IuVaag+qV9TTz4ok1C34Zm50480GKQ1Y2sxT4aXdRbFz
KPQwK26Fa2/HyHJeGPi17amzt+cpt8/lJCjM+qnNH2OAMl5PgI0nnRFoBMy/dd4y
qso66kB30JXDye6p3Hhw6NWJRnwkaevZXo54c+ereoel1V3YQyIaD1kjzhY6yDDq
7eisYWIXu6/mrpSqVnG9QiMuWzdAUYjTiBtHreDQthSTQGPPz/biWBrLsViQjboh
G72iuq4LAI6WJQUl5iaWnmZSh1BJ9BT3bQXVOKhZlxwlIdLpgYzIBwTnVgHdczs/
mntTPoCeIPE//CA6UYyr/eoJJILXkKNUP99qUHXLLS0kHKgDiLGsZwXbd7EuAHtX
4cda/EbrtK0n6r11Tje5OL6EMsOYk0y98Q3Zbsq4YnEabPL+InBnfraJ0jgsj+Zp
uJoeORedxjH5l7ZAlvDa+gSvln4xlhcQS/AULgEPIhDvEJJDmo+7ds3aXFphc69U
GS1xHIAGLhLdN58U5Zsu5S0Y0PyOaaqFXTRF0YBfC/puOtcpimRkHnZvgn7T8Eyy
RqgUiS0Lf77YhY18jiLV5iT/WsNf9WMk3F1GNvTkUOti1rJLcYDxn210LAfM0UXo
CjJiZj/ioh/cV4LMOYV/KMFMjvUeLJpcsyLS04EbqyUa/2KeBAWih92CzFIAiisd
NdK8RzTWUl0DjSeLcRcKfJCcrzt5U3CJaaXJRwFsOv2/RVTuokAcXoseQjmB6LaR
5701zucQKDyBG2ROFYRwp5GLBFmqV3DQdGROz0hxYp4Hrx5oEFODBIdMxd3qJIy/
PKN6qnQsG3xs8zCN5YUwuV85vZVmn+LE+aSgZW5rb88UVBEucVq0bDyzBnb8H2C7
aR4h/hMds3Aa6GMe/Oav82UJx2NrpRqMS2tShed0j4EiyeFFjd2mFnEDbi4e+MZ4
IopM/tA2oFEOA3FwEFFPGzAWdb3M5tzJwrUhRu7iHeCjPCeIgC1gDMt5UL1D1Bj3
PCUhsgNF9BhB5jbiCJ7YxbiiKiBCv2ULDLwcclYOSe/Y7uvE7u9jX5ZaFxf+fz+1
OjMdqr/J+eMvJhaMdUsnhj32QtSjhxhUxcFkKvCLD6Xt+mwGCH7UnMGqDAFx1yIz
3J3HiVZu3OSJ7gXOSOxAYiJKDoJA3hrHhl1jzsifNd1z5yKKtH/CIwrBLDAHBfqe
Ve2T/QC17IPuF35J7M4s1zA/Mc6PmkDgqmWbzOJQB4JF126QLeZdycZShBZm24PW
dQpUkUZHh053jET0+uVKhkIyMd7BLGfnOrGRT8rCqC0GZwnM8xFohgU+ndx70Jhr
/L8tn8VehttT3tj/tTt5AbWSf13SPUFMbBNDjnL7IAksFhqBkW4NlZGlJdgr/dy/
L5aIfGTaRS4iRdaa1H6ke/GYe+JL+EWd5Ws2ofnOLMBcUhRQweQxDjm5vHqX5M4R
56m9GICkc4ewaVXPnk5OUY7gaGtFZJLByedWFvCMI9SHALoJ3r1jV9hiSrmQObt8
+dkD6EgTbpnZP96e/BY7W9DSG33PRwUKatVjlA5b8Sejn8IA/4KjxDShYeQRoB8N
djLt6+nAffWltmRRdY6b+n0B6HcjojX3qmx35WlmAPWEBsh/U3b1n/OPhd05aDrF
rGWwgBS0DwUE/U9XQ7Kl6yskw2dK54bpnT5GbnBmYFkXal3lulLJyUo3w9aPqxdj
fRjX6SmEr4W8LcNnceThwPUxN4p4YAr1JJgY3C+KM4nsG9ZE+HCp8OfXZSwjo+qh
/jh8tBKPVETLkMe47fLhWt5BnjGu/72t0BHYnuP6Hb3CPMN9AcTBhiEGMgSRdded
tEjwF2W88b0Xhq0JF/SlFjp3zqTAdg5T9FZ+dmfBwlz8WP4GyWuW+OV7X9zEssyQ
FZ3LOPK6y3OAx2fuGt2tBDsE+miRYHVxvKTwMiyDqgsrp3yu8zkxbb5d2dwh7+4L
SoL+Ejtgloy+CDN5Hdw/Zjx5aHbt7XG9sTWQEMEvNJw0nd3Y3VzDlzZQSCXK7TTF
K5INqThVThh1dNWxMsvwxH8GA0CDvtLpje6TIKwc7/vFhw+5MJ6e8qJV5JrEQ+Af
MUtzX78Yyza9yy2yJsTJZpztn0HNco6ntcHRbKggldFRACSb0sNZo0OsF0OXSaTs
8rBZuM2jkfX4WcqmY9GdUqkVbMh3v924KiaXzxLJ3SfOwYPItBDnDHTC3XDA0rKe
B8yB6m2sx5KPjCgyBIk2AE9yiEQKZmTvYQdGw303fVGmUX4ySpKPDyNuGFg1a0Y8
R7VKpWo8mR3khjVLpw134F0Y6hvdpAFcSaTst2x4ORcSyjtQbXm5kebKFOG47Er+
1CRJsBlkCfLLiPg7RQv5k9mkkHS7F9KruqwNrj0ZSo5/U27g5XLGRor2bOABuo/W
iyxHtBZb0zk5z0FlB33EfGaJIxT2U0AFXYI7fwly/UIF2lU8QLFV9Q5vdo9N4JRL
2ZzaNVgAazlH8Bseh/6ZV4FTNG7DagN4YqaJoIpoLok63iLzgfGGMZJUqNfP4/2J
NYwbxdyh4FERT2ZUKBTR08Jn9HZN7eHVVwyQN0heFFqjGQdNgZmA4irx0uXfgo1w
jEhegCzeNGxbqjEADFhlnT3s3JK214DCoP9HB3aRLjCp6XH1qUvE8X2bsS6y17QM
FIWPxvp+Bl/hW5vYTZO+6AXKhuWrySe+qZGoTavR2Io2xA/lcb4QtiscEIUQfFq6
oVM1f8hgDNpSaKqp+oeXGZdf+kBAO8sLjOCfUDClvS2ehq+iVh+VEQbnjetdmIpM
9sDS0a9wL0I7ZEz49WT2jk5o9CwOe55f8ILj4GyonWqzQH1+p/9/uGp8CF1ytFL6
cnMNjmfp79NtDJaVJk7h1GaY9/RjOLFbuhO7JLiLrmRK/fWM42xLkcKpA3/sSDlz
Z1YyoLIp4le0hsuOgitTbcF/6Qog77EDUKXnm5Aj5Nvnjwp66aXaw7YNqaagISor
SYlRztMSmt7PwKkp3uTHKjk6yQF99I036t0cSDqSVucRyf1cDOAcPbQKkyXl88kj
uq7jh22FfkEYRQUvGBtDOvJyIo7sFLksg/zHmM6G0qHTxA5Wm49uHgt3pINLjGZ4
G2VkPVdfH2omndU6+IRagXjylHv3ybk4FSQxbu9DGsr4rKvhAq4nW5cc5vTuRvLl
GcMynqmGUqs17cuck4eUIfUowI2Evq0ik3ur0H6fsvKZCpHTK8jzRGsXAVESTymN
k4Hj9V0N5wOoVJj0hlIEgm82KRFYQMHBizL5CMv//gmEiEFcAteyIDAumObmOdtT
Ga9P33Au7u2EOmNuLTJwlb5SFZaOIUkMaLShNBLkiCfBZIlqPIQRvuy/5Sia1EHC
k+zlbGT3lAqh6lfBc9xOdcttZvBldVSibpkM5mmlz5mx3z0gJo6z/iBBqlvOYbIn
3UM9o58hmcQx6qgwZFh4X4DkjWa26cakv3ybL52t0puZKr3rcN5G2BZULiCQnv9/
LlpfI2NTPWivVVrzzfCRR0DglsieSeNv0WEvKw3syHhxn53/rpgDqaeyEMZ7WtwU
tEZVJzkjkeAu55zoC+OPTvnzIRn12VVHfRCyMBmIOh/0xZ3FezA5vL515mRWYx/z
ttoYYdPE5kvVd9ePfsdXSwG9oY+dU9DYEtxV74dqi00Kwly/ywg6cdxrawbqxCsB
YXAJ12WJlX0VYCq7ACVhZLmDChgW2K9sKIBlMjMo1FDHsixJx8CGtHA2605Z7fBP
yDeXF0kdHNiO2RaLZ0KEC8+7isqLsOQ+xTd1z6RFNyTxRfCr4mfiniBxSPGQgOcQ
x47ULgeJ7MbFTwO47JJIGMQYZM99ftW35ahK69ONlDq0NREvMGflyolMlGKadsrF
R4uCWBjqBeOLF3BqyZpocHu++KEChslvrD4d53SXYrOGyJpeKArxQ6KJ/H1+1yQK
us7zBTLdERxL5/qQNqqEjRp+OVTupsUzw9M/B6p4Nm14RmEON4A98/1XrAaFc0Lb
hrGsdmpXpLxUpGp+zSMMI6fWZVE+pIS2CWxiCz2WFw0nmwPOwXUweuvpi9uiUIlp
xmQc2+l5LJb/MQuMsi88YSQlb+iYZM1Aul/ZVBIGy/KnjOmS4mBQcs9saQpPiz1X
/GTMPdhI9VDRWMMZ/KhCBF/W4IeeicDeCwwmjWojnk93Ojh+luy+JF4qvKx5/Vlp
PS8WkAgOV1JP2kyGDoW9meaQIx987LPZB0njn8bVOgO3mUFN3brSzPcUxrNjiV5U
kPt0P2++HJRMC8qfVDMOQ4DRSscxzDmtQ9in2HWUu6C41CIc/90d+gRfXB8+yTyq
NRaAZmdoOCcUb9BUYWhgZGzLTsqQuVWL03mANBkGlgeuZYA5GPkAf+rtA1i+nlSQ
2CKPMvtZGr8Pc5mHbGCoilW58NNnIYU6u7tv/rmo3XiQHf2cm0hF+cJGmgtAjpkm
9zxWmZw17GXQM1LGQrYXQJed8uFkZpliyHdmvq6mL17i3cbeHHfFm8s+SfkTTOfa
bVMSeL2xtgJTQ6McEUz5d/xGC0QAmmtVQZUFcIKcYGbd7QZzlwm+F6uQ6jeJRhme
xwmKcmpSWVdTkOYg42ww6lDVGE5Q/OyxIExm95IBWHbRUMK7fmgXM1lXwTima4jk
XWr4G4AzqNuReK/ffJLp8RqmUbmltsGm27CO09bv1OBdnmCd+T6zb1cvfr73kgvU
Du96cJWfozBXvG6mJzais2YZ0jueth7Lrz/dZoZdsYv0BO8Z4mJt/pS78WEE6rwF
NWNh8MyPsyIyTUSgaV+gTe4yo4FBoJzkCJ6AWPODCeZAmgZZOZenh6vM0fdNhn+D
r+tHDPDPoezjOsWKCNGa1jHGaMPd+1xKvUaE1jqd+fldKy2IyBYTi2qUZ7X32cf9
WZ2vONrmj+hjPzn9GEIFYgdfXi1yQ4rf5Wizk0K8BMTCPKI/dEXL3j+YMHN8m7aD
jufZ35SE0V/LSybUpSL9NpzOym+T32U93bPk/TzlNLnNLsI66GpYIiD2uR+dHia8
xsZoFmvg79NfHHhH8PaMwPEsjxxwVlsHg0vHGNMFfGlVxM53wTvhZcHr/oEbEGaj
7jAIAGUmxNHdAuK+cwAnW/Ap7YxIRwRgiqvEAJlCEILPz2301drIgiwCNYLwqMTv
74RAqfW+G3r6SDMBQ6LgAkyC1kuHTwU8RDRNepdxxE7K4RnG1+cldVVCYjE/mJ+g
zcyXw70M5hs7/wAZi5G7gs4w3YSkSVQL3+Ptx7Y62ptjOx0/36GhxDBYLqqlUM8/
kHqVS+bk2qFqZBOg8LRA0RlRLkeXJgV+JgIVPvtcmL7TI5ob05Z4zoNf+YTpEYXP
oClm3BQXPyATV1lp+QtFTV+e9kwTOgT6SZrcIZc3LtgdyUFhHHzSNfaiPY+FBXhi
L++Ca2ncIbQxKz6zEL9VYpTkTBo8ys6kMkQLxzWh1dznmXivkGxJX3pueIpwIjYY
XWm7knOl9mGjB8ObFu9Av7mUTUCF8B9Gf+udsZF7mSQC6MdjxveIlY5gxfVj3wFF
Hw3FbDVY6X8Pb326ZvCfLC9GEc1SSWJm+7e3/T84payX6baNIgk287fp4HyWEiuo
aQvgYkVAfN93taVDfh0OXziGge42vpqT1SuFwaI+6VONbhiYYZh+Hc0GpolDdZnI
idNRXT+uEFIj5eZ4gJCisbxMaGEibxattTXoYuuw9xf0lfR5e16OW1OwBjrodCWi
gtFDTWFylwGCcJVi7zx3R3ISCychg7iwLSrY9oM/T2uANpw5JyUCRIYNMz+w3Gc2
udof5WexvUs2ZIKb7hUpu34ur1YO/lqRG4tq+kOsfM9yyk7nSAn5jsEZuFHHIFkw
P5KryBEG55tr/M6zzm/IzjOyC9rjZ8Y2HwCNTxmYlPlDt20+TcYZStrDy4aMB0zb
mSYYeqnWc79tcfJYij8sXzsxUIlgAnIJXvXQYXwfIR5Wua2itwQqUyi+nYZDWvQV
ICuAdg5eJELKzkC6AcfHyfhd5rGt6yG3u84JTdjIhHQLWK9AH7aPn4bouHaaIzMD
PDeVjL5Ev7E8yfJ9LpczLNmIeikh7qugTX0KboZzBQ34Jgx27CdSa90hfL6Mah7L
pKxIm7OjyZ6u6wpJO20AMFKOY+g5r4e0RwGrj4jowREuraqBeiSjzBFpuz6qsMqG
crZL5Ib+ppvsjJd/e8T2j5KxP+5+H5QSVHPYQ9+PHjC0+ousV9wLI01AxREX2weT
ug8jcjqz4hUbSWF+TsetRNnmmr04xaE+UCr2bawvCmpuaTw2sFji218scgwdKH2T
k205NuE1wxiSKtkYkozu5R1iekwdrnhz1f1iSvgMm/MnSi6/A99SP0i1oKv39sil
TLB/qK+0pgjfm+ijCacirfGj6TFNuJb/U1CW4Jbyh1+t8Un9PzL+YkLucYSXGzKx
qF9eOREI2Duyhhe30RbVkELN7YMiH7RrLzmWwwjSMqTKurK2i3GKyghjZ92olQFw
UcQyT+sGU1dNPFJdQDqZsb6EuhmEpm56paSSbJHxM4kaCcnMBKGwymHIHki6Bsig
il7VvWUjdKJbr7dU4VkpPJLJmIHkIEUpFt13Fss4epQJw2quhPo1+976n4VkMp2f
YGe/T5Qe4rEbRQS8sClNMYG/nH2jyglZOT6mt+P9fnB55oarsF4ZtplDmJe/MaF2
7/G5N8GMNwJrKAvs1CS7V4iSIk1jqY3WPTIamtiz8aEtFrflnOyaI/Y09v4MX8wf
LsENqSnW5hAzPxS+VjQqis30sEaCcW28ZiOtvXazMHfKDxwcJ6Ugd34EZJETB7Rt
ce10aZO3dKQxtXscBxB07NHnjZjG00x50hYWn8K9U/8hu7ETrnowFW3nK7kP6oK1
K3lFpIz+L/svmuZSKHe1TSK+qXwLm/K0kIBOTUJOSuCbodJzbf0VkRLJkYOfol6i
SgjWN6BTDQezBDOe6i22vU6ZF1l9dnQCcInY9WMF0TkAaHAh1WNAW2JZKhVVauaF
uqGNexYELGJ4yrSHvFxz3ErYbFwt5SUb72Enb0Fx9q/GPlDnJCm8ZpIbvpJ32Loi
QtEVP+HaxcSZWVWrTsnY0expbEkqMw5T/rcp2VuAF8axHGgEeCqD23fpM/N2xzhc
MEhJx+fxgFqXVmSWPY8tRxY+OhZeZkJoGYJbbdHQRWK4FjdqCyJvX2kGnotlNE1l
mqI47cYLuRtZqc60GAzR9HtE2dqxNPqKD8XBZ9LMqUiR9W2TpK8tjAkzv1+bDVJa
qa0p29C9feorHsXESnB2xamK4WpKhBEixHCQhpVIC3BYXC6zKFw1TX8sokYUOERf
i7+X+eavF0W04YoG8xw/AFDOfOsvBNWJuUxoNfy5H6P28o0RdJs6HKSLLfCdnLby
HH/3NKCOANDmBB8G23TX5n961hAtUruRPtBiNGjgwpk9nGdfEfdQ6W6ofqlp4GM8
i+atrQUiD7PrVOMY2AFXB22aJnEzQHA1WhSaMgTDRWWHRathFsBx+OkKhA0uwXut
J+tfggW/1fxh2CSC54SbgLLKMYlyNFf7FUS+tbg0T+Jz9qctpAShqDMnWW1QXkXC
RNQyK47kQmG2kw5PonAqT4Nod1h9EqPxH2SrQDRqJAzELxzk99/m9BHDnHBFUfb0
K4yOdn3JrWbys6mJ36TunzXsciZb7PlZsfWS2L9bpfUVnp7XIZ9vqoaU2uCP63gU
8H9Qp+0RJiKRgZqGfnydVVplNyDS4HiA7jOidPrC/UD5/xU4qELv5MhGiomvXXH1
TVuERgtQeiNhTe1mUW83/6bI4oM5z5v59QIIGI8seiGv4oR6vjmHdBkHoabHIHQW
wASzt/VED9usR23JjuZqPYT8wPjFKxIvvlWzy20kJqUVsKcuCay+hyvzsAMvG3AX
THInzktw8N1vvdFUlIZAbfIwYYyvXjvrxt9pb0gMrL63OKuVSxBaDaf7E8v/sFTn
9qVoW1zNwP1HDYnyjZSOwgCHJbgiM2DWA3jETpqqmwtGnFgCzWKvu3zpgJzQJvew
dgxY21QODhAexz54FIj4nP6DvmtnpoIIAvBTv1IcQE4QmCkPkNz/1KodXtFhFj1O
1su5F4a220/O+TZO8C1uNVf2RjV1VI0MshEZLj9ZMd1EAHcdz/c/pgtSQLa21BK2
Fll0JZ0TXu40GZYYxgO4qCniYvDXiDTpsOJLiGID4miJ0gv7FCBb25vThfGFMulL
UjYx98WwO+AJzZqKO2KBGFHXDlSpkVa81MPEaYOpdLDVgiDxLh5/4UwvQPpyyziN
BDmbFl9sWto7zG06mS01gPyLe5kpeMJ62p4ZFhyPYLUdMC9hMEHJWMv7235n3Agw
4a+1kiDtM3h7UkDGWjkYiBsAr/A9NqOG5iVFbIGjC29EsPglsqzOXvQexj4p6xru
qYooonoEsX4dKCaJk98YUjMbsKnFiNRkpPu/LSxDGqnQaQUO0+raiOoWkzsx1vHS
zjNLIX/yxh0aZ4PPg/xCRxaqV2rdeJ4ky2WaUDwkmKRSFnz/yoQ0KAS+CcFqCOdR
bi+/gDACdIOffYS8wjSDnJ1sr++i9h2BJMYelHzMCu0e26gY0ifbWulsbLXybLVo
rRN8oB0VXw71PklU79JHW1vZ0UH9jdydapfSNQztsp5GlD+hJVulMY+wBFt4fuuZ
75O/gJUJWZHpDeh5SfEwTVMnwQA4mHuUZBgWGJKvfpptskApxqex1fXDehKwS/UE
RjSvDJNWdDf6k5H+S5teO2DdDOrGAJIVzgNsnMWmAnyCEN3n4Fy5T99r3T4SJrQv
YbSJpo/N8gREJk5sbeaOFpMIaSl5z7SywbyZSX3xAdXDWpJZKYEUkq9ujjSW3I8H
t76qnoEhM6FBO8+1S6gh/t4zCuHR9Schp6eFryawte4wfvoj6+bcXhn1ybbcILhF
pqmK5g6XiNEm3RbtxMHPIsfUQ7pvRR9FBtO/48vvfIPhddZpAavD4Spm2nMhjPKO
pBAdvGGnMWQCFdASiMZxwOQ+a5rzgORP2KjbW6dFTNbhHCPKMijxw0JFUSx0hoKX
GZY1gf4TdBcf29Y5K4+5pZ1JLQ68U6LwD52EhBnuimPzmup4GJAbexpOoaKV21Cx
38OCabbXY/EoR/IrdBl/5SQQkbtRyGxrJIRc7AKOZ4VM4c5t/Zi7zchEXw5q892q
45B/lHp9opd7VQZO8kWdX7Z8JzJSWvL+Hiivor2+AuVR+DRrzbirSTTArZoDHr+j
0RVF7AWMre4DSjr+/ypxPdwcqxJDp9389RXyEoGmbySo9UfuUVr7IVgCstd2820t
BP17wKLWlwZGhVM0gDu60qxTAERgeYWtoYKA+m6PDHuabc42ZJKBv4xnOPJiamck
I+6sv6Ja7AIFdNYt6KTVptXWufNxsxNhiaYFl86p/Q3mKdB0n4xVQCNMxk1N9qCe
2cakHim7obfZGox8thwgQQbhROatyFhv9KSHmV5XyG9+08CJwHphhNzwBLfxD/7Y
xaJekv09E9G6dQP8d31x4yJnhLNVfl6DTJw04rMGCTar+1/Uop/dbqxtXdr7UYBB
hOoh3btP5bryoLu+AzH9hwMUWARIDawbjOFEojhcXo4UGKz9OhUjyGI+w83mcuwM
wt3krdfdcS3xu0nGZ7YM0/44PPO7XiwOgVW4CFzCBw3XxkSB5RAuKHPOc8TUrHSG
bUAGF+sqwUbBKcfn6YeSMPvI2BG83hisG+qZ80ECztsXkCUUfX5bYsY0Xpa1sJ48
kfsuvEiEHbbyERV4tBkm3xbSRBDDEWVk4Wj8UwHMLEss7G1xkpu/WlusdTD/xNVN
IEXGZDjhA0mCLfKtBw9ZU23fg+RwIkGOAzDgKDMX/kuIKw5OshGqPYpW4GrQRDSz
pNM+ZMZnFyD8DVaitfBFENqukHsVdBLBguFchmQSlnYRXY4+JaALzar+lemK9W4Z
o+ZyUuc/p4HIThE1/vfhHg3UzGk1c0KPLJO6khaIiWXp3SgADmMNvtSaXGvxWDGH
fK1SpQUnPXD8NE5ZPDsHoWPLXBaRMmx4iQfawqRasrH0dy6U/aiJO+1sZCdqLqFz
hiZLX0SfzFV44F91XG8u8Dl7YcRSODNBhy4K+8YqXlNZkfc+a+5j+RCzQf79sM3K
R/d6zW5HunoMDhAMxb5TI45WuRXZUQ9f3jbojm0ZneSs9CIw39tTg/rPmIA33SjX
pSNRUAiX43wSe8atx2lL8stsFWZe+c0QOEpIQpqPoV0eqin5Sx9XWKAfFTYhvBEz
VnZRpmuH0f/R+2995WpaNlHEnipIBr+7aUHJKUZvIaccEuNhjH3uWCXj124O3kX/
2CX68omChWOK+Nn4yuidKcNnqouUQkn/caL75sVD0UODq6V+Bq9K23myggl3mcgg
x3BXbHIygIly1+16bs41F+Ik0EAJTeoE0rloEe5Rc1+KS7BuRCHtjactRbRU5usU
aYYePoApP3XdG/TCOQwTG0VrtGzIDKtBlCRjAhen8mak3uUrNrVrdkoS1zn68x50
7nNnzEwsXmOxjwga1u0drJQqvSdDuya3H4PwHe6s+PsqRGZuUTUgyZLIcCisq+1O
QN9q5Huh/wbk5fi77gF2CD0dgn/6VGMXXcT6cfFtyY7zTplTLbHKtiq28EXekik2
kOoC3wGAzQ3E/zQnf4IiO3ur4XjF3u0hJJNcBwEmEFpTHKDHSTiAWGfcbGBGfQnK
xFqr0GV9yMKO7bTbnV3tvJ03B3DErL2vf1MmpL83PyT9q18lCWv9II/yH1GK6TP/
lmopIVRy6GLvpe/KmnCCtKfCWF5QkwZS+0w517iEY0HmMCgVoX9pR7PVPEXZfO9P
l03yhy10GSmIvBJevjSojDPrrdus7fJVv7qMDKfypis8/W172cGOMgiiff029zyE
EXB/z6KK+RTVnvUskWv9seSoVotJh0HFHp+nsjR3qWZlMPapb4aeClAHW8oranQI
KSuj+r6QWspvW8pj9Y++w+mwEnoHujWyOxPk/8Ry+Xia6tBiXikf2g98JBqR5aht
wL3LpFWfxHILGYzrCW55OuidRluvklAlZnTahVthwPHnYnP0OQN+Mfns6rJ5fctO
NPnge3Uch5uI5C5tAREWp98wIGPZrBka7+f2sjt39JLcUcgdgliOCqeQFLoM7YUv
iTrKYCmciYCuvGNq+cBPoGmMuctPVndrhxDYE/jZ68+xOQGdk0po1r6f3LnxxuHS
Qo989wkK7y3nYym0ncPfjxeOVlxrX/2VPIMau7qavCg4+kusHauysvA1ZmHDCGzQ
sn+KQ6J1+YQGQP8MLGsIc2yYTsmmibh5SEenCINKn/5qDuv7bY/XOk3xg/6XqFpY
VRgyNPGQ+PCzpqxMb61yZgkjxZHTfZfH4wWO2SZo2pfoNAy/PinhlJy3i55wsMqq
AqyZGpdNrRrixfLdzvyWz2jYWwLr+slyCzb0iKKbrlRk7kFkJALse9GqrnfbhjTb
Dvt8i8vFz2FJQyO4xNKf26SHBcqXOv3jeXnM0ILF7K+g3Z28l8RHnrjBQVeEOo6N
4/pLa9DPciryaT3wDioQA+h4zuo1Ly7XgbEiJiWMRxDyR6hFLetkK7iAl107u1bG
kLXymbiG/KkJaAlNDZ9/8AC5TUlBx6eXpRx6G8Mxmd8QAbPRiBPJlPU42NFPKsJ3
hf9XUXgxwTEZcqw9axLxKM0mayngbCKtjKkqPVSvHLQ454ss0TbUckl9LOfW49nG
JTGAZgU53cqBw3ayUWWTSaoCPe6s2q+9iLnkfzra9MhB+rLVOhq5u7S/UoRr2I9t
bKMmpchu0Wla9U4ThRsRoHlNEWyJoQ85pufCXWuR94p3cqGgNSP61twAXn7boT5r
slBVx7a8sQVq/exeWY9ibBy5g+LxdKc2HRFvawV9ZDBxLBwyCxPAi+cq4wJcG7Oc
adewuji2suNmv0QZjSiOxgwmi4Z6cUcOukiA0Bv+XnraggzBnVyjPsYSb0uGOTzM
UXERiHjM4XHxssHHW2YgwB3y15YpMPiLyZAPZbkAyE0NMGRWxZEY6XW0LmiRpdXV
7MfHxSK0xAj5SwqDeWkEa+twDuxtozmqWmQsIdYjztmqsXgIgcq4L71x7mJT5MHp
8vz3QEICQTwTNoidANmZ2kgH5DkcJ7PirC1pyjEidLjDYKTpeDi8VIC82GPYJEmA
6SFA6xQg+rcRnWAIubcHdIc1+a4l9iFgkiYOLhz0EH8w9gMisQsRr1u/Gt5SR9zl
nPtPXzFsyxGD2Xsk9S9k6/ZJJVwLvXAjTScTyoBCRB/5EmHlF471Cvdx8yTI78tX
Q03YWQbRs2NobzUl0Bn7/kNnqOrQge5se+TkrPNqF2L7uQbajAOPhr+GlyIgUTcd
Oj57cmcWIbYWM70JaFsblI2pdulQFHU/QnqP3c8RCD2DBInQ0mjp0ipp+ISQAVo3
/cAJnjOWUJw/IwZ6fc2d3CfoRsrgBznqq57Dy+c0kbdLpcbnD4yp4HSYhWr0g14m
CEFiCWUlkALdeByJgKBBrZRMC7NETFa67daV7tKxkVjLE7N9l4lXbksvt9u5Pry8
ffbG/GQn6DCvMl7pFkbg2LCCIQgLmwI/t4qUgxfpirwaPpgpc2TKgQsdbJwaM1aP
3Yo6f5maTLBK7JpdQiXxRWQiT3ksXPlRcFRZp9QfGdebKsmJPCvECiVDXuPrq8kt
Vz8xfi19x2+Wq66a3nrp4bVPWMYihlEn2Sg0sf1L4MI0nF2gn9+eWc+w0Dl1dhwJ
2GDMbQtz1GrTdAQvEo3aJ15Ucc7ogu+q4HV6OvT1Os+meA5Uz+AefSx6fx8eDQnK
4FZunPtHgy54Y8jis5dVFMbcA5SQX+8BaahUZxkl1wmHXjHgAcIAOoxmRm73kgTz
VrOWDShxNqQBn6NT5+oR63JVnUA9BKAulyBoxFe6VbiN55Jadopb+El72lHG16hu
79so37r6USYiJU5PoczwTEZmu05QUA5JmCtlehtJYdPjijwyl02wZEkMDXhaKsQ0
u5JawH/T5KRTVkz1zZMGdToJji134c0APKBYucMCXXQyn6B/8WtidT25QY7VbV1e
CL46/hEm1RvDRjuKAyTsBF1cMt+Ib9KrNEc/8w39jdjOXcPHjfplrwc8wgSJv3Cz
msaW6PBmoVferDJVxNKAJh7fHRi85DoE6K96GnhPcBkQvxvFnBznAxHYZWmzACD4
ebyUBGnn+2gJMgMly8EFgjSwlKi+5iMXvYRKRs7MOT/2Pyo5lW1qCf7rmIcBZ6eR
FPRGj5GNBZEe/VG42MDkl6j1peznBoWGRZ1d3uLdEtaqCtm3yI/FAyaK7FVZifk1
h+oKwmzTgfPoT+aTssbZUeFbINxJGAeTEG6yhw0N/bBVfCfPelGkjZUukz0K6SQG
5BiiT2snGiMTj+Uvubnoa5eIe9zUDpvXDiswyhGnE9wQlo8ha0hKgMzqenw2Rad4
IbnwUGM106Vsv59KdXi1p8DKRkpMxuJ/Vg79CED1t5MlUt3RgNsKSLmU0tXtkJCQ
4mlutRGltAt6/sRNslMNlj1+3Ar+PYv0i+L1kVfvck7nw+PCMG/KvF5MGFyfnDt3
h6eQCSLTrntfSzfge+dRhOXslvVw/46xAMGOfF2m+VL7cnsQ1m599ejIrP3kNwEC
7kOtnJVlsI8b9Vi25ke/GU50odvk2jhCrvwvfRyA46m82OfTtYUQ4gZp6p56sSYE
ZxXmfPj3BRgSCgnBWhFIvP3GVnDEfuR2/wtACqDVz9CmG1XmFkZoBRgfijquV2rE
Q8tcdPb8O0pkGqOM46ZBm4P9iO2EfoVVVNjjtcz7uk/grgERCQPY96hmvu2Dt/zJ
kX/cMyS/E+5H7LtJPBVfcdTJw3U/Y1gI5SLjNOt2frggCeZcs4vWRElQTz8guV56
mY3WF0vzP3+f89wSo/mqTz/fRl92hfSFHmMcQ8R4aB+WETrxELIVPqjQbQr2vzOh
dMcpi61iF6GAHDw9aSaeqwUrtG1F89wzS9q8ywQHSWJywBXd5Nvl/uMMA8XCQoBw
TRUyLQV4FxX2I3vVmtGEhD0tkS8jrEhknKTKU2gGDmiGUoRFZ8Asp4Ve/1XFXV4g
QucEarqsFcl+sA/2Tv706WnfaJQSniMsil5qyRyIdFuOO1p+9GcYWL0TvKx/nrlY
YAx6SiLnewNJ1iQo4fOA1uL6MCmuayh2d1iYMIEkwALvTV6htB6pWJ/KgZJjBxoW
d/G3hilUA0hkwAgnJYRdz0LurJPlMxyyvjrEpNpUnyU8qhmRIPsET+tYj9ktEsBe
hrzLHjOJwToKO9R+HBhtetl4ICY0e0Ax3PvIRjSlVu8qD36hX1Qc6JqFhpT7mIpE
6hFcZmHoezePIhlMmbldJS2U9cJ+KazPpx12ejpVnUs/Hd06nvEd9vti8kPHlH9w
DO99SPvG/TyuJXKK8rl0+eu1/hYuaf88K5jJxEGpgBMlFg+f6jlwK2fB+oQ7K7vw
SeqOlohyCBjYWq/Jk02ysJvhDTAZHtip+zQ/fBueK5vCm+cPCa7qdLSlcWzibUUv
Dft4n2cZnh8gVYsFu41vWp0hOAXUKM1/rEvck0f00QZz0tjovObnV1DaVY0XK3KA
5F0LdAvHmeL1FAn1kPzWXsp8tsyxWGICZF6vQc/X1z49N2pseLHmgE+20yiyuJVA
FoN+pVNvLHZ8PVM4tAhpWsPNq7Wry1SUsr5FbTSQsmlOpNYNB6eh8ofQOAkoa6or
1JtcMsGija2zp+nU9lpt1YAQY2AbIctH5MfHlSAfouOreKERETrhVSFBm/d0QSp+
dgtSBDV2UnZwMlnMroSHAtleeaA6lr6Pz5m+jD7p1s6eb3r8GfQxma7+hoyvi+3/
3QdEa1wIiJb6M67I4+g1OlcW53NvqgBhrWSIg8RWl1tFB/ofh2EZbrgmXTDwJO0Z
UfeZvLFwBCgK9zJadBHQ/fBVUJubZanXYyctjMi6/3qxlMqSs++NJiu8YACMj9PS
Ccd39x/K1XqGoUhDzCqgvGdre+3zGk8qJb0b0pOfjAD4gYaHmGRAlF1RN3Q0zDJ7
JDVNPvd/IWCCH3el2gjDwpBtKjGy8RzEGxcxid5D65uUieW9TQ8OGSPn9xQntJBW
QtdQgs4X4R4ACTYwBjsz5LP37I40jWzm8GdDRjqSWATmNXFl78c7Of1ERY49CxFL
hTkGHY7Mcq8pEZt+02oB4N5iwd9hqInY2yiGUd4D1FKNuCqT89kKFJFU+Deev7nF
JJTrJ4C/W6KmfV6LBmJw57QHKN+tg7997FMTKUurpdjJ6Ch63aoyZkMXumDDSrB6
OEKiUKMnT6rlf96bI0g0ibzpXlp1ia2S5/A1TIBKh8uC38qLWwK1uS15+Joh3FNm
u8PrZ7bBrQFrGCkCm7H2ZdA1++YIjEjcV7u5HYRuwNnpyQI/oFaS5KP3jz1Uz9rs
OIIQhe99dQdWWPvSRu7JX7lcKvYjvHIh9roAyv4NQv7+Sxz8UQ7WLzyQPyDWBiWz
r+tZVKw8OdEj7mbjmJswpRX3258GSAjeJt0uhPoqLr6iU7bcqwKB7DAAoQs6hkwZ
KgXobkn1+fJw3v9RSqsfaH3TGRIZvr3Z/GLw6gYhWzaar7oimkZwTQiHq1ZmOAtn
VgxRCxz94BuAmAPrYgmRL2V9vQ9I0oAaMlovqr/ONy83rXrI7ZrzKclbgKiLYoFS
k29XqXL33yLcDySRw66T30SxS4WGQ2ClCqyhDWvGLx51BTyILa0gzNZLHv9I02kM
VD2gU+q4ljF5Hcvo+uRc0mQJQbESz33r1kpgU1JBl497I5BY2OPmRmuzps1SJ1XW
aZXO5zj7/V7uYzOWfqjCOGoQ1oHRD55GunjcDa9jBF5bSnDktRmSYmnp3b4n3N6x
dgBCzN8hIqkYzul3mDsJNZIYX9P2FLatedJ4bN9hB0bpvh/sCtWUumtNDKZXUODP
0krG3Aw5IuKfByOw3o5lMunjDRVpC0pMkW85tUmI102E6Wkq9reQOp1HpepN+lEn
5wYR9rrNkuOBW/j9uK733XgtZlKIxIfbd+12FWBHDy6DPaJyB9azDXscBCfy9cBo
ef7CHqHKFP4DEml2t6P3yf20si/sUtMFuhFr6Kfa2yhQQQQ+DZWptfudq4Nk2aGK
us00DeONPmQOxMvJYZWG9PCI+cWCES3aOj4Clr7J+v/qLqUKDJHX9PGqguKSYm6N
WgoneaFKqfgEaDUDD+3km9yzq3HWJDkAQ4afYCJ8D0j49rNuxqNkCH45p+5fZUI+
ZLFBcFGkIOkqWDNFp2NSAy+/6V7WKtHuiyTSLDrRuBdHIQLUsuxhdo5MoIf2PHFb
XBHsax3DRX4IRUCvlfIWPxRN9/v63Og/yFBgNoVVTE4gsO94rTuI3xal5Jdtj+8P
f2ZaH5SN5NmzB4NYrK8NHX1T07pVj2tUSFeAhs/x6L7LfYZ2npxljDIVL7qwhfhr
LJL8Mm7DZncmMNXXd4NRLjfy/TWmSutAOT02qwSDTfiiVI949j8a5pnQE1OttCpi
eErhuijofGlhEWjOH2ITNO298/PhXH76VK7fGeQFPV/ZZai0uCDEelrK4ZyymPbw
FfaufWnjbGmdb27Jito46lUCLtIOR032A9HvrRTwtlnieRnZR8Wv8HlQZcLdtf4E
xkgXd8EisH9db66O9S4qRW5dhI+kjkbb3MlVY3b8zAMzxAOImKMsxkUqHmy3uBIY
wjYEkFVbrYty2Ii2wxaxsOzqCyIEcBJb4rXBJQLfbU0eAVbG66Yq82rn+mzUDCom
83E0trujI1imhex/fmoyiIEscA2oAKFO3uhtxK3ZJ4yEwXpUc2lNcr8XJK3Sk4s0
fRYEltOIpLEYNw/zXk1MVeicjuW81y2hgTC1ixvQ1QYMjyLIgPh85yfLDrp6CbRg
7VsA12cDFW1GQbc50sjBL955GpUoXNiHsGC/2dJXTJA5loeFIf6ppvXapACkVDmb
zfRaPBSlBiTYhZ/4IJ9no8RChw3r6piUDMUo56MbPAm5p2TWozTrlTpVIj2twPf8
K8IiGsYw0kMNFnAXSehdnbEOx0NgTQoQdUu1GciMkB0EcgjelyXRFAZVEtLPdIBD
LnnMJ8Puz4XWgWH5wCo/DFwYUGWHvLT4SJ4kSSculs/9ed2gpe/Oi+7iuBpV4OUj
qoaMvtjeK6fz1TCJnFYo2U5mFzBg/VHW71GtWQ3zS2kVaLT2VfsD9+qHsMhe2BDb
PoAyvfHMHWFkEz77pLgVODbJXl/abrf/SW77blLbkmlDSE0rEmaqY9MiZLyt+Jzz
dVem0h2ROf7sF4XyEzYJe9FypIeF0NIqY6764iMb2gVoVbxDuwOfoOsPvgm3y9yp
QDRH7ziknkXr6qKjVMJWNXY4TkTItJxi5TRRkwIGTNezcgO8b+PWlOyVZjsWqFf6
zQKoEah2NOcT+/8lBnoDbPZI2T2YZNqlR2txc//8OVSz6X8oOKOaNXQJmWrjPi37
IbvMDzkdyGL7Pht9pTjeFARNAxB4dbIZVzz6gIv5Bz6rrLvrrbgbnvgsuS9j2eBU
w+FaG4wzyxoSD8Gfu0fhmgt1/xDuqHwCrK89qhVkiQnCXhbZ0TP+UoTMYSkUHljs
sP1XmNSMJEGOceS8JmHnKzZLeZtCNfR/WifUii5gyccD+UVHydAGzeg7GZurQ3+D
a992tKMwgp11rVSH4L1cr4r6xGJ7ktwVaek0lk2oVwnNOcjKScoXCSz7QW3HxNUJ
d26z7ta4cZ+Y6aUOYXaMla5UJtMuYg9J+7xhe6j444duI0su5Ei54Jc2JOXbh+AP
LsLuEavffGT5/OZH7DpzhZmRuhdugO11Iyqg4Iu1sy5ZJymgaxguYRvxg+GGBuE7
kgnbwZLkuYLKUn3qiJgaT3EA/Zhcin91BpaNak5eGmy++VMa712c6F1InAZWKyrR
7HkZsZ9rObv1H75fLycCB7uzeteaWTYomhC+2egVdNWH241FC871YQJ99rfWflgW
AO4LouaPpTzRt0JTaJ6yjpX1NArqwchVoAQXu10TshHiNywQXk/E18jTufpki5eN
5NM2A21RiIJiqOaGjW+Y42OZbvVWaP/yptNWHlkWIwgrRx2jSn5a7M9VZ689tEEp
csHcAZXmd/IramFqTGv4kc5NPAwBkSAm66VPzDJKF/nGnpXLQizR4qx2J26ieHPf
BlD/l0J+q9Gv+r+d57BTaoqGPMbyl79jSQB2+Eykoa+WRSRT3+bvd3zGupfxGcIs
USaJX2f+A1Ylmnw9A763j5B5wW9i7BmY6o+OgvqltwoEvm4PrXWPBZqcBH1vU24w
10u55e/FFnO/sUMsZ3j82GUdGO7In6NFeRXU5ZEEr+a3i1oy6rQcGWKUCC0LvqE6
GjA+Fb49JrJOYZ7RVYOhmyc3jPAKwRh6dj4lNnumK8QwVqrOc7CiuVgTwdT83Mir
WcCaVhM8lquRWzKSNUc6XMhDWTrIQGwm8qHAqEFBd/D5vNxVsFNw5zv0Mzq/Mj14
rz4aIGM0HoU7M/K590A5AVuRUWl1PngdaDzHBIHa3g6clygyzinyxLxSe0WiZsYE
bf+UwRLdH4VMMfHK57f5XIoQksVVobvCg9KBYx2tf2cb8adRCxKNhiXA+bZpsoyy
dQ58hP7YsyKWndi4OZGzUs8Gnzq47rzf7BYxfea+2/6/48rAvihxp0sMXZvrP+5a
DVFvN+Y6f0515z4pZKxTHoWP93TQ31c+CqjST2w2B0ODyWY0lADrkT0xoMMk46rJ
t5TNPvT2HnWRvGicKym+SuEf6UGvvJzCKMj0tXnn3NvmR6NUzhT1ldHeH24gFV6Y
nTLoAeLKxxc0zXqJ/GDn6vajhH+kR6Ae15lOfSLVOUEFNnGkmQMhb1MvdSNdKZeo
dhyGkkSTOT1JBDWvPJXPLNlRvZLgiguo9xDGN585jAKywiWz/TOBDi4BZ21xfPGX
k7Nm2ajz1D+htGgChkJea8SWVJzrKib9BY/ucc2/cfm5SQhzB5RlC72zmmpAwzlF
Dhxv1cgwknZ5bek1+JZP3d42Bf1HTm9Hn1xa6y5WXwrxGV/fA7GSrRQkxyhKFkmL
DqEAD7IK4zqOKQ2GT4IWHD4pA4iZ3BEV/KOvKTtRl1ay/29fIsCo4dD+LrMh+Bor
1B2dMz0ESHcXaPM6rERM11v2VxIAts1P/eW2tKtPosW//4UzNr4T28E1it7pjMw0
kAFaCBWszytnv98jkZTTT50K/dhs/RwD64oO4iaBSeOy1Y6eBM4tNKClv++/W9lF
NfYjxIBgJxC18eQPGlzoZ53HuKlf+wMZbNCZvbHAI1sIcNJrt2HzN9qchzT7d/dK
+qZi2JNjVUlZErNp4OJfX//5e61rpkAWVy+f/cg7G8NgcSFtC9DdToPtGY0khtKt
mXcZ9BaYcxrzHRYa7etbkabEUo7wbKefvby1S/edTGQc5R0qa8Pz5aWvHy54o4JX
3tSPrlkaUJopOpFTC2FsVhG/NKiFsq95Kqsdj4VrRjXHm85bN5kgNDTyNf7eytgL
NTJ9kQApfVa6IAJloag433HwHwHUXrUDD4h0q6pkzpgiJcLwBhDGDPVsOK7T7rsf
z7m1qZHpyIT7nWmknWlsHtMUsCwpH+FZwwQ16L/7zoLNtCVzpjCgEtaNcMOuCit2
DsRYkF2aYkO4Dk5ACDshqY1Tvn5qBwcdKDrxB3xftBCZ/jYtc5cR7uMFTw69/QUz
5208Q1bDiLD6IpEFq+JhkV8I9d9fUMae7l1pd6clAagjFrw8Qd3wHthWOPs2adVr
OYGP9XFERo0qXa4GhkHU/L5C6BLPiBt8jaykGcWgL8FIY4REjglXUph14UqpTcO5
yV3t4k32dZj/lKZ/9ZGFPrK5BZSJPJU6BjZGl1xZEAaF5WUiOU5HD98mD+vDEA5/
fTJ1mrsPgmHI7dhZelqRtZIanwkPCrgFHhuDZIp1T1Mzc+RBd25IEvhogggzRKfQ
Me9F3sgMFL5VoS3jpPqvKhSnHY4v6KvaW4o4Gh5RxpcgJ4g0yBAkdG8umeeha2ek
b63e+QVxJErFdCwZiOm0YwWnBwTZ77zWNp9abiU4wXOCPGjMGm8cEMugeNqvVfRa
7g5OEvrH0ezPhXbPOPI0MmucH9LrvDsM8ncS7K5omj9yP/or3roeiGqOH+UIImX1
oLFBYOQnGZgZXH76WmmzUQk3JbVPG6fjk/6PD0fcb/LqJ6jw+muFa6vk/sFMeMqm
CbV2UF6H1aJRDQgoeJ5aeV4bqdEkgSRPaj9iux0fSevcKr4s9WYQ4sJRm3Be4S9N
2SHO7ulmPiNPjaque0ecE0dJO4UMA1pJy31yz7vEtpejXwAc2vI+biICh06sw8VY
YEM3Kww/zIn2H4QPfz4EgGBZlIz6ZH4kxnHBj6Nz+KXgNx+GVrX726nUOIVE5h0V
sVIPzJQjYoKLN/tLCl4iB09/Iyae2TwkbB8hoJRs1N2mFJchlaAG4TaAa4C/IVA7
v8VmpO7xwpnmbqxOU4mMYUU7lBEI8oahIS2OXCpKMvFpMp02VuOYYZ7GXG0TsXmY
BDiQBJVJkcR9eDzEMxljl/jyVqhl+6mUYkyV6kJz1vtClnsfcJiScp3mSTLQdENa
SnP4zFHo8UubSycgXqbNntG23txqEz0FubT66Vgz5sH+cd9lf+uOzPLLGybZOgjm
F7ASmWWGJfI415X3IZ44Gzl95ivk7XpMwKjuy++mIWKjSP/X4PNJU63UkuoTxOb1
6gmE6E0CKb2Sdj5Rw6DqKrRZJG8SRX1GelM2Gk32nTZkmBJlaHx2OcLvvPyDt3xb
f7eHKHe0X/2BIbWskwt5sLUi+WJNxFL7cKGbaBUTR3xCQtBsJa8rXfYiH/VP5rCR
amSAYWrsJ/s72sS4slKyNTsfX4fjrTDOx+hfaJjEKsz4HyCvzd+mWCT2BWW20Y5Z
Jegb2wqVyHWzhm5NIxEwzkyCuoHuUgbRrYoY+FSfrPyqjnpYOE7rZ8c71eW6rLUN
ksZsPRGj1gxkiii6M7fSVdNsXcYWNxITBs4bx+jkkMnQg0/upGebzzRxHVArn051
xzEhuWFpNAKXrURnXWQUKC8v/IDPPHtrV4H3mgBX6dsyZPQ0PWjS9uRWgJOLjdaf
JCG1upDordQZGQaPo84FVBABCmWpmJw1xb0u4uoLbK5ay65/FnoM1ygJnHo3acwp
gHQ1/35PPMnpFQ5swP5rP02HO1B5U72gZUelkjxHEG7Y89qh6EVfZxTo40lrmDuv
28f18kj7l06bFuwCB3wUGZ2r9p1dshDFPO9dk5ensDUnIjTK/mSNcrjj8wL+2nEe
zjL0zJV5lT+fxVu5A1YuORnll4th0EKZbbvoEQ9eQyLmy1KVDNKxo4G3S4YeqpOf
aisNoRit7PYqScIMtQoRMd071Wg8XDDpNPYljapLYX4WaQZPfa1bNV9mcuyStiUM
8S9BAGo8P02yK1YJY+dNDZ8qW63sYuh+Ci+BQFCE079FVPONFZotxo5BOfrRzes6
EHNkKAyJh9alWMC0gPxh7YdKG4Bsm4Soj6Pq/yKhVeCaWbQzodyIzx9s7Z2EJxM/
DL2wAaeHQ7K2KloOE7IqnzyOTCiuUIUxVHCnUv4ykhlisjE2Dzuqk5R+5nzFrv0O
PNUliVLkxmI2b0v/SD0+l38Q2ag8hcAq/lct9PWOvHwSM73pd7VcM8wlo4oxqmcw
+fnzFrApF9vdzNkPBIFBDfONkl0mB3k+2ZDG38q957XdCJ4ndzHH1z0riiaDEyFV
zGh1QxWnzJy4lTdLaTP/hqOWj7Gw9cAyrZEhtl0CREw5+QuWx1rqf9x2GqR5Ft2j
elEPyQ53yLdScAZvjWeKdw==
`protect END_PROTECTED
