`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CymU2rBDWV4AGIatFEQ7pTVi+Q4yuAJ7tv+tUVA1TSGOFoQVu5v2PxcE5fZ+L7Vx
y5fgfVCIpsvnfOsG5ri0ETKrmdf+ElhiacHcDMQCL9zrbtdrabWr0JIoqN0rtK8t
6IfXumGVu9i58HnDgkRALm0oEqY2Gd7voOK4Mf446g5cElS6JoRl98qSq0RzNHfj
VEtE7ihooxGV8rP5HFQUAKGextR+pfRsmjhoaNIxj+W7q3E0hOWWe0ZTssODrMCf
V4mUcwoiRFcFPQezP6CLt/I+l5bB2vtph+qdwfiJDQOcrxJzy4PlA0kFjHMfXNHc
dskdx//RbuUIvCV3+3sW37BBAMhUeUmXwTODelrt+mDVlJUnziSLnOMfZWhTQ/Jd
w+14QH0UVuB0Gc3vKV2Qx64t6zlEJibc0bjH4//ABrnBabEV4tu+Z/y8c676G33H
NhX+4h+s/8EI6JH1wMt+7517IOQRlGibYgzXhwUtM0BA/KBos94mBQkWmzNoSRzR
132R+384pqXNqHBfCA97Kyqh+qxoxa/I+R7MTz30jbF4H/tTn3MtlCHnYR0kVf9t
eBfjXW61tQlUSxoYLQHL4hMvtFe3SuXnFmTHDu8cAwPt4hfmOlYmX6oPCQ+G9LFS
jetUE+VyEFFsdXYOwLC7sDW70uQ0zHK+qCFLGjIjExm7LJMiqUOMpNE87b4UQLUS
HJ4o6Mb+BHpEXFFVzMvtrSQFlhBbwaTsElJwUzXfz6SQ2CIpteYr3CWuGa/QjPfF
k3f5Ds698h4eTRhjxOIO0bE1YosTio47yvxfbXOeQ390LUDqSEbNFSpqn6ot7oqv
o7FwMd1oy3f3abiiL9gQSSEYO/yYyQbNRNlsQYCpnxy/9wR4hi5+xgsjMF7u3HOn
eBKNv9r/eyAEEmtogtOPmIJ5suBYdBYat3ucJ7aBnBjicNYysF+nvZzWlb5xDr9o
`protect END_PROTECTED
