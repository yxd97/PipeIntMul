`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QjwdKzFUAUldgcjd16Ah6wp5XcbPJt9jGaswsG7cwyBu6XCo2Z3UWvfy8z05M6Bw
FOsZHmPYQ5H4oIvcPWVsOGHc2YnjIsaugKI4on4vh8B6p/S8vnvmSPdXbdNE2IGJ
HtaVheW4kwm0cd1qRC5J2bqz4s2ONyLgAONEymvyVb6r/dbQsk9LGqEkbAoBPYiE
Q1Lp/v0nv8V2WMBc3YC65CUVUvAd9yxpedvFqOhn9aaQfs8y+VptSHsW6BqBJVOX
ehAUf5ZfI2sHxObKpYcqDhu6cxsgvG2NRqSrrTfCxEdJXdi5QDzbNFneHv8Jg+BB
H01tvbWyFE8eFLey7QQKV7bTsIuaMWZKEDSavn0eRlitdsqWL1OW6LCc8Ja8j/Gk
DmZLbfcYLB0U+ELTiArjKQmJ8GG7JZCSQPj+8wcZ58A=
`protect END_PROTECTED
