`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
om7IQ08bIMXRzkM/xpc5M1OaiuyoiYIrHB6IrD6iEpVNl73qhs0PpDpSm6CwG4wz
6NyY07S0PyKvWbOnCTMslH7MHbTmsoZ6WOfmSarXUmQVzVnjwXaZ5Fiu1+Ssj5M1
rmx8ldXl8hCVRNjzBv6bSc1rGncj7FrFUjsB/NWfjqjk5PQdQYpJDAep/SB1pLwI
TJZmy6GD39IwtCKWy1u+C4L3rgWAOrZzlgnQQedZ4PjgAvQIODNpjbi+9C2WWGGm
rH51yOBIObw94URI23Qxb52WdefWERTn8iDQAroAQZ23IqCqEoIpaMTH8QcGPEZh
6MN26EQbjFGIvCB4QCyG7I4T/uEIonCyoKhZe3ol4WJUrbCOoE2ZzuM2Ku6MQWaD
u/t+gsw2bHNYoFYpMijb5dh0JJCAmoxn0MJn+gBJM5d/fc/et3LV4MJN6GbHU8DX
`protect END_PROTECTED
