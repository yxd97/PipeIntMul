`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S01ydFVBVx8ZzwhsY8XG83ug3zKDqBlBVZnA2wd2/++B0S0J5GMvXLQMwuXTrXGc
0YiGa4iXzipRVub0KDgcIOpryAUSK3qc8hW9ft5tExcP1K51pbqbjJ8VGg2Rv1bN
cgdIZr9be4rOCdcrWOixINvGgNq/Ro+qFgAVarM+mPLMuf5M2mmbYxoGzdC3d+4M
6k1X7waMxNlilBjmw8VfDSBmL1m7nn7z5tBx/Bh0Ef6GpyQRZojjoHdxOFohzDg+
CndMhUQMB9pu+prLppDARHiCnqAhl1JYd3Tfkyhhucgz6Xgs5Wrp4+ZE2/9gJcuX
1o1Vy4Ulmd24+dqdqxKOYGZxnsI/Ejq3OSjTJts9Qdixm+xuq51MUWdVmRstGUT1
plIIhsv7FkxKraOwh55qxNEX1aLxtpU5uh9SpzNowLtQBrn+cnauE6E5HzB0pTTT
4NqWwMHq4bUG3dvsmBtgKimuJAwIgAvZaqYNjMYFJNhB6uEtk58Tazp9ir44K6vJ
crUTzJiEFqCJG3y339aaY18NlNrxHbweQH4Hp38teRe/pCJubUDUaidczVVda2YA
66HStrjJEKd5njyrNGHuS0tPK1KL8HjfLt1G1FgyuHnpKbg0sZEJ9xlVWJ3VZfyW
cs8hi0g0+eVoI4WAUqZLI79IEFYSEDzIgGznBB4yQ8gIbdTutG6m/a/aBs9npH6K
cbAusLe+cHENHmLM1O/otgtJkbtfRUtqEq7bEtKX6K1hJUQaponJCsPOykkOzGxP
Q/D1JKB/OnKgHM2mHgXrcgCGCSZP96Gc/bk5ZUPW/Nu8kvfk1EByXop2PN24TQ+a
7ikmnq+gtQU4eYbHowEMkIkBu6yeGedfjvIOGKM0STIjpK/kpBtBEaKY8Hwd0mUy
TbgeRCLZJ8pY3DPZ0My2lifdTH17rxF4enNgQvKj4sO/xJF9DWwebVmQLUx5OtdO
fztBEjZ3zVZwuJmlLDTDEEY1qN7xv7j8baEGigdXoWxHOzO6qRffd07WXwdNSMCo
qdr7TP7HpYZEC9FxyiRPBnQRqrMAu6w4H8IaHwsV5Og7AtasMHAniqvbRjnj9iyC
xA8pGcs4za4mPprXBtHU0srIBQ2un3aUEzsxuU0ut7+zp2vdkT5Zcl5iGPf40gGM
zjYjEqBaDDuhu6r+D7vB4f6bZjBJwKZQt6aQXA4n/C2lSDT+UbX6q7Y+EtbJR9lK
YuEfxh3u/GZzsQp4FbmZuOKa4TjUueaUd7xyul0ykin2710aN9u4jMZZSY36ns1E
aBgHkTBKJwOOr6QtwNrGpPdWTpaaFp8/MOv/8A68gGKI5IIwUgrAcnUAMAN7Cm2v
gIgEDnYiXS7O4EQ12d7esgxdhYx6nb7wlwAtH9onoqFiU7ruYgc6DZlTxQs7qija
tZ1Cp1omtHQh6BmoE6s/2RBvQxk3+zU6Ho4LB8Qf2V2rGFD8Yjqt++CI+m++bBbm
S3mlheUWJwl/7sRw5NFwIAvYk6yBdFBb68LMiHTsRwNxPfbav4QzXZA6SJkBCyep
ZokA8YCFFL7hjISG5Pe70fFIHSORIupP73YOyi4s6y0VKMwdPljnXmZd/w6AuU8b
6iQPB2CZINVZM7a/EZpYQX6E2vU0PSCH7WF9ZhIanMEvvfSTWxb+sMGwQOD5Qolr
9wvLi2sN2aWRa7O1Nv8OKA==
`protect END_PROTECTED
