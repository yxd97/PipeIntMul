`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qs3lbUt598OV2dZBjo7IGuXlzLcqN7Orrb/UYjbb94Fpg8uLiF2SAlpTP/UPHUxi
yWk4mCz7JG4KoUTleeme2ze8Cs+YZh9oMq9HDqD3tRT3yYWVKf71SWMJhzGIUYxr
JywOHpcRGIuCwrt63ShTu/9ex62GxmPz85qmBVByeQ0O0PzBcya6mwiJ279foAhy
fH+2hCxKKt64x2LHhkUwkZAuEWZitL0Ruzi6uSs6cKXdtSYaXKXfnZFqUiqIyKNw
tJo9oiRP0XMQ4QvBToTFPw==
`protect END_PROTECTED
