`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YYWnvljF6akU+BFdhco9U68tPFZ+DBf6Ib3Y/T2SemTxYV150RYfChM672SRrTtd
CUZnncge/Y3AgLBBZvbD0/rQS2sKYHhwghNcSoM5yU7MHmiAAO6rZ8D/AZ9zdCOi
9SKW6/NYqtcMqKcVu5MkejwAA1OEveZsagjVkL1o84/gGxcrsvUmK7RLKjRKL2He
MzLUlG++ZYTHAcr/6E+g5rE6fOn3Fl4lvrCk4UTZoxjRfWXuaEH3SJmsjmW9jG+z
VyFztBFwsVVnrEQCoL9mTaGy1UbkWrrkPqzDcjkBDAIpS8U7RfklliuV7i/17Qwu
QYC6I7CwqvdAN+bH4D77I1pMUPeHncwVtLEW//uhMX0mh5YyBth7QfgKk8eqqAdN
l9oAxjHaMIN/Nd/d4Tk5qdx47WF7v13hZf7TIhALeGsoOky8ccS+K4F8Cj5bqkWJ
0qOCiVHZT0SG6kxYfs4NHo28D797jVg+ksFPb35huX1qMNlT6ey8VzPOHtVIcCy8
3gSNz0meskayd9C/PGTgLBYgH5m+vSirS2cTG2go58NTuyy5w3tZbbwb6bQRGhvW
6v/Wryzprf/VAkJjNji0Bw==
`protect END_PROTECTED
