`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fa9jR8OvGS3m+qqqWwbqsIfJboJMXasJ81rb8pymF8idXCM5+jA0EaBXkVoFQ/A8
mrBSSPstJkmWxOzyG28/ebEMOV5Ob/QduaVitDhvatsfz7sMG/52hTM5DrlFgfH6
SU3zHJMB3X8gMuBE17aZE5+TKVZlub6IGu9YwAJromiVWgB/4xhHreyX9t0uniy8
PKdctyXXyhwhCz9ZYDUFXWfMWROWsGsR9+uif/LW44ESXedzq645AUx2IuEu5OdK
9O9W/mVFtggrkSY5gAwGYfmrwS/K7CS6m0jxcXg632scc/LsQf1Ikki5oPBopbex
Lw5lMOVYCfNVVRzJ3iMAFYIInS4+LVDZMUF2m50qyLvSw95IkpNDGtlz6Hm92n0g
dGlzaNitNrl3yOwNZWdfywTtTjYh+473Rh2bptWHoFPVqYFZ5SdxgKZgcqXz8IqO
xz5lrLP0rqFevXmfK5Ckb7KSugXGO7Ad3J/ctTEglqYKX55i6MrQStfsHDmJfiTo
WB2gYz3ogfFkptIjgBxx9b2Z8eMD3F/mFk17rY29buDnyy+L60nBTCq7InkSKyTa
xj2t2Iyc0tNxQPJqxN7C4jbIlsOu7rT6boPDRGAxg0QWLsgvpYS6rV408/SlhUvh
T5+Sx15PowYyu/F1Otr/OVRI3XFnXd6ZvSz8gCTVVwQ=
`protect END_PROTECTED
