`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qT8zrSa4ufXtCLuS5PRSepy1Nxw5f7ibBBhZq8Pie7RRbyfLK+IujyyfMcWCJjEZ
HmxPb4wZTXfWnLG8nY48lvsXTKUZy2kR7oZqjhICvNkj/6MfXGfWP+QckG3A8KRo
Pg3I3CgVjkbjmh61D39yO7/Budy+fn/vcqQMaLnxJWt2aMy2VWGPIZt5IBnH7GFw
usvaArE59P+po6vbQu/5erXvL4Y8PhGSQJUN5tChXfSnqPKZT84XMdkFvZqdjhHi
vbfrt5jj5RRtyAZoaJn6W/WBMwvQfvcduyWAp7Ns0gGHKOI2DWrqY6xW56UCgcIi
fXRzkhA1sBX0vpXMxXnWhpFniZfj7d7wo8bIZTnxbWWW9o62USU3xvXBzno9Ou9P
MfXP3TzavuTT09YmgQiuUg==
`protect END_PROTECTED
