`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/9A4D2+od0zmhG+DOQ8GtHYT2DudJ36vRwSuP0Jgu1OEC/enbbq/Xvx+Ao7DlNy
lxhI4Al+MROZN7eaHC1PC2xpyA/vNl4dC4fZT4yCYYQznv1OUYC9Y1efrOdkQxB+
J0WomryoWl12J2Mo8NKdVOccoLMrKtaScA/2LYAixG+NSvJG2ZezNsmhl1Jd7Gv2
s1DhjdHu5lU1vKlFdpTza9EgoDDiKuowiEwNCmrL8lCFAgrY1bnwix3Y3fQrsdam
lBmqFbPVTCC3bMy2wdGZanLb1xH4VNxydxdLqhvfoioSm5XujfdTa6ZI1W9kEFTp
rAQzG0xp3sa0odT1S0NRrZc144QO+7sDpoSu8t7D+Sx09MEhKnv84yyIye351tQr
jKGxShwMZybm+12iBTp057zCeqcrCe5T0vuygmTu1yflMQ1bkdaHqAFPfJxs9Z6D
VG9Yr2p3sI4yn4wn6ML+GbnKZ3rxH2EkvXLqo3mzWC/Jt7NP0Y7HO+sYKlgRiCZv
`protect END_PROTECTED
