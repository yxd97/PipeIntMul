`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EL2T8p30lQekIZWDIncBZi+h9zgXrEshLhI/TkqK/hSF3xaBIaRQOSj3eW750YCe
ePPwU6FjjLZ0MHbSWP3ewWYrTsfQ7ML+CjFfac39m7KF/WygiNmc0GN0SL5kF2KC
VMbCZknr9TTE0ylGQRfNcqLl65zwJkufPlIjIPL5EU93QFTt9yBmSzFvYgpgcLZN
eugot1ntE2Q9lzH3utX7BV6iYxINGvOpoh/HhFGto5NDbGHIpPi7W6dN1hpws52K
3VjMLBX+g4o2AQHTSBhgtFAmHvABbbg+5uGN/dl95Lb1nGR3Qh955I5h07dAfs+G
2eERbFXC9a/z2WZdYnEQ8CrqB+LuGcO0zHYKQ15IOoDRnzBE4bfjNYpzwgx/C+9w
I2MoEQRfMtkfhY2g7GpU+dCk312ybs3Y+CDp+mDK4YoPm9qJ9q/wFx3S/NAwkzDE
H+T8a6JHdAyk2Ti0K/7uujDHl8wCjQItfIsbr70wRBY=
`protect END_PROTECTED
