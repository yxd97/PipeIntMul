`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P9DVFUiqJmnH8phpyS0O1Bc8pg1jX8Go6HS8XbgXISuE5/1/LUT7mrnfpCq42SW8
OhzE1lwfQwPsqChcpt/HEBwAay503aj0vM4CqWNuw88NZPPTLnc+LOiDL4kUQHSb
A8yE3Z9mY666HyL6WOqnS1cwGct1MjhUnXgmvYy5N7PScuJ+I5vfcHznB2vb899D
pfwremoaARlZETv7WNEUpgHOr5+n3NvI34sWAk6gwPaAHke5E3zLkumEfo0Nv5P+
KFTaLZ4eLU6+zLo/DNV4F0Sr1prCwokGHAiNSazv6D3Zmz+IfD1B9Xx6tOPiyd3u
lUbdB6Rsnh3ryAduL5cvnyxEXfjeey/BQ49mixfL2Ab8aVdKsRxHVqIXQDaeOp44
sLGcrYrjPUgxDG6NpVJIhemRihw6S5XEHGBOnKPfnKPN4pZKRuibSz3sAABpRiBX
qX8BNFaIhRp74LodqDTJrYxlnb5zkWRCzutrKrkoqQOB6/nClcVPXS4Mbzo0GFVt
SVsbX5xKrc8tCsNRHm4JgXvbsoyAiSxy+fiqUG/mb8VAzLMQ27OJfR8hay4msLOp
KBnT/uuibqu4MSwcisqOJcuGjwD03SSTwl6qc9JPQpV1/bSTzoBznIWmDCNWj+A1
LfrXFDGCVWxgB7Ij9yXjjM/4LK8AcKdpfDHBq6eflFjN0oNbmOT6nFw8IR7neydm
EQLasfiZ/6UwQrttXdg/Immqm9A4WGUebywgxQdWgzEuUxgf75IL1F/abPBJh3Km
qsOd0pyPU/G6YofCWSIMbn570/i+2m1gwMKJRdL7rFZfL/gaaOAI+1TEhSzQ+sJJ
cfVmHAM6ReNfNvTzxuPG2TVvEmZveVZ2WJ3s4eHKiNk/kGUueC95b03+udPd0zYh
uvQQayTQzUIZbtViCOTY0BEJcieqc79TLkmLLfozc2sd/MsSQKK3XC+4ReaiWDgL
zOUU9Q/woAXz7swIWW2Pt+rPogcIeGgEKdggAr9H0HOckfTDeNIZBBuWmEkARu56
RzMt7sFN+MyF1Ag2LfUn2+MKI1prs6RPjRy37RMpndcABX55rVuwUzJpp2NaSafc
B7wf4oCweE02r7x9OqwQeNzDspG/1ejbZxbnJ3pqkoXPOQlVuCnqhWwiVkvyaIvn
O4P7yTg07hee/87Uaz0izFaCBLrLgL3uC8xtlWIv9f8MIrEPIO1jhp+wKcIdXEVl
WBXqhYkl0yUUl6dyUdV41RmRNZCrx0hFiIhFa2gKF0cj3eCFogg203N+sLK9ZZ/S
0msm9/7WIWDlGc1zr5TnveE147BoHeRTaeqOgJJzr4mePr0Gd+YmTNVu8GUX1yHM
QSJPw/ennGpuqT06t8dhsfSzK8EAo2IafrKt2zmnTAlOtxEUfa0qzYFiTlx/FEkR
FNfLalh46ybfFe6OKIX+/ao3HgCCpPpZ3/rZ5Jt1x+Gxi7/wafD0havHaZp87Ll7
vL70C9u2ws5Gt/y12bMWE1RUk9It+WcDUbK+5DqU7LsrlVzGFF4GAk1bwxPLTIFI
y5CCGoZ3dClGEWRZuKloZbjFmlT9uBAH1GOUXtwrwaKjR3clklavfmyGAOpcewtX
4ZY7BcEt1/UTgVTxe+U0QtAP1KwGex+4MoBMrlR8b8mRPZg43c4zRp6p5c+H/6wB
uh7jRFqmQFHL6DEihcLgkuViPRfUwcR9Nr9k4LLliFXK5uiA58xbnte7J3ZARJEA
Y4Q/w75PR9oBAIA3ClMqg5swFfed1h9tOfupfwE3rhvFRIZu2+H3YPBgmCzA9mGa
5WMYKc2N+oLbkJ7micV6n0DGGXf9ZoU5Edd0Q7Ble8IpYXRXm9pOuk0/C18fjTPR
Wh38bojvPT34aG8cdUwFma1qXAMhKL47ddO62aoz2Gt2Y1KCC6MGn7b2LxeyX+Tk
BkSIgKd2NErSqo0zap/bnZa+3TZ2NOUmRnaBsEJn3DmNM9kHI6lQ5r4iSJgAG0bv
7/L/CHBvEwPOHlBUyWhuHjkpPJuwhnvQx13m3JLSKH5jmZVkgzCkwOWfR1RgmOgm
cXmCsKdtSji2Ndb981hFHPRR2ugNrVD/pTpruza1dxbIAeewvgUIRLZ+RIOaS6zZ
L2aT448u47bsAoFcKfrH9rDDgX5/gc9TFIKdNSujNyUt7j/uVvn13zviv2SI1ANI
pxBtOPV0QFElJaISkoaatb66KxxxKzBS4M4p4Lb7WUZ0OMzzgLnvQ+jdjOqtZgAY
CPVs7tJ2Rt8hVt+mSOW7CCWu04wq/tiuRcHXGxdLcH5y4ubJB3hocW3uWbIzjSBT
70PVMxYPoCOLaLJLesDzvpH5ZwMyONBaR6giKC/Bqb8e1JvSpS8oXg8FbrgBFpVA
Q+LE96s5PrFWAA+HqoiG8ORo9s9/W/4FXAQsu6Ahny8HKRVjBQjRrHnWcLPyljwa
73PK96jF199BnIBhEXX7C47g2rg1Nu78B0ZX6L6+F7y09bpL+mx94aLi6mIynMuV
vhy/2mUorpwQYYqJnD2FcxLGQbj17KYl9wYcfsS4hliRmI8dKL//OvDzjicu4Sow
XiUpfac6K+Pq5Q77GPrO0dTMIbm9/kclJCAb606RniugRIL3plZURv0XXy+AcmKV
wUjrLUaG9RlHJpJPsI2Ht+zgfOadapfaQHWQ0tHqAyWNqOHnC/vkr1hiEujqCHup
eVIvlR7dIf4e5TTXhA0BTw284BlmBtuHyymRrsjn0qXcjvWzHs2ZXCll3lqaZzKY
I4i6BKCBWT97zIvb4u6scV4qWG8Rp0GihUq7SD321DVU1e8FWKj+sbhn7OtEEzeC
WDQJmAEiW7eAwmxCnRxLHquNAxRkcMmugRcOlnkHEEVXpt/3kwwk8mvnxOS51OwQ
ByhqrWvmVXbjvtIX7zde4wgYnMO2JjJlb/nn2oX21kAk+C3qRQLD2IvfH+CpE8IR
9TN//oq5sPwONkvrk+NBPq+udag70nWTo1JNjarew8G/VsKQ+yOPkNE/In2YB3jQ
ugHr32ytrw7LjUmw4s90mchD7Aq9/xpLseoEBLvaeByKaEYieEjqMQFOSTfkoPVR
aaDo5kKA59vfXLdebCIO05AaYglaWkvbcr1m0B9bjjxQSbQ9VbfJx6p4w+laAcn2
sbGEIBI5bfyw1C6OsVDTdxv71CYkFJESpizJJWd3j5L26Ksho8P9lOTx/q1y18jQ
YFyxtUaY6CoXPgXjh+HsTESj/e+EhNrrhDqEAP5weSdaen/zUTzu6DAKNykBoNhz
WrpDSqxQpiAyx1nEyfT66YZ+rcB8MyxZ5h4YBWSyB1h6To+6AIuRR7VEqT8kVa8K
1W5gyr79vFh19aOjtZ3plR+ZcACZnhjtZLUTTKduzkAWfmzhzXwKqOboACxJo5WX
f93F5shmpLfTyj+srBNuQGPrU4MAtoeP8W6dBZ/lDdigkczo1XwuiZ9YG01v6MsU
UE4tXzGqQpeOSQdTWrWFVBKbYMQPhVfkYN2qQyg6dqkSNLGWgrVYVbUnSXNfWTeE
GTQXescQlIru0dJduWGIkARB+6TqSCJMXaYR3TdrFKZLWKf8Wti26uYS3pHuylyU
81bk0h2jhuSwzMPkPgy2X1cUgm8fnD6e0uHUCACW7nsVMFfH9KzY3hohaCcO9frN
9oP1sXz5PnPn0VD9ZtRUeubdUG4tDB6gp6ntlljyZ9xYDs4BjtfKbt+w6Cu02GdF
3QfHW2cyGxvxQuzT+0J5IClqpnPp4CvreoMeeVYWH7/2nUYErFkKK0Og87malywz
F40uktP23lkYFAEapP9LP4m7vMioSipqwnxFD6SWMsW6bNRR62J9/392qLh4rf7S
Q94qFUCmY/9XuHrO7HgxHQPzJSk3+qczjrOzh6fRNuawlH15Tahttu4LHrMb9o1g
W8cV7ihz5TOOgSfROnbpkuDvUXsgwqJKJ1eunsTzjDEjbjsF88NywBPLUJ3EcgDx
0lHq4NiOl+R1fGnfPAxB+3aXhRJUI7ooj8ifDsXfbM1oHOWhnCYBhs3aqRehaXSw
55MN2Fv0posVzsYYqpAk3iLaN/p+fca0YH7mFZ8iHWwLP6YxF8vICHwy63R2BEG9
2YzbVrdimq2CZfrXzoK3KjtLC2mvR3BmohNd4av88GFMlDkqCWoDNfU7w06olUNY
n0MbfW+Ba4r1bUCqiycvgzeUceZq7LoyO78dn/XJbZh3eHxAG3I11H4GJpFjRbkW
7Xe/va66l4Kv8HYMQi5ylDoigjZTblbxU4IzOAmxl/bXrRuvV3Te31nT6WE/QVdl
N3ld9kXFQU/K3Hh3iqKMlif48DeMeLnXiWbQYLWvYt5qgS1wj/+V86OAldE0t6av
B9UaPHHCxUJQ1xdHW8YLUsEU0kzFCBOJrxyeTJLWhUv41PRtdGelx+8q9DWd6JSr
fUgziyzEkKTT0sNFKQKKDgggQoPFBzD6zXo56HEpQI2tsiXB7kNhfWl+Rf4PWcz6
+zoJrEB0uW+eo9EW3WzZDyGl5vlZ9bcQTbRjLcYXyQ6y1onPzcGENRe8emIY03he
5QEGC3jyKG/8VZ36ayFeu+v55Xt0SZC3eW2ASU096gmopgsoo9YFNEOeXBaxIwsQ
kTxpDPyegwzjXl0HwmwMoJ6ZKTH6SrfmxqoJdIliDcKLZYVfuHxH5eY6vQExX1PY
aa0dotE01Xl0Pf/DN9dPFFG4J0HrXKAtSVWewijhvlwIquczqy+F60SuftjbZBsv
VudKrAcp3xFOgSo6UF0+1Ggl4kWK2/z6S4xGu8tWlrq4DcOtw7GyyqfkJyy6BxIO
x1wQZlKDERbj30PVKUu1J1Pw/IWrdSUVcnJjO27aQIDLhXfccL9zFuwZ/h1YMLRm
R0OzlxzpCefybArE6b+1dTy9Yrvfjptmma6Fu9DLzRiaHn0OHcY61qnva8diOSRH
SNdyyQp3C/fXuPATOBBZEAQAXATcu/63+mssXkZhXfVGXNm5Dm9RXkVX6kQVp5xc
rwLG7Gs0eVqqilv2Vmo2UUYv+uPxW8VJXeiqRoDTov45nU7yZ5idMqV0Gf2ODFTn
pS3+DyzrSlRLgmTWGo/Unyh9E43TThgYblIqmQ8FKrIcG5LSEHlUyIYt3z2h4war
ThXntfvZXug/zaP8vDsVdK8WyPp45mMFYDCoiFYYLk9EuKUrPcmOVUdqiU3+eSo6
csdn0DqTRMNTtTalMImrYWNKmxlAWFRiC1QUoPOSTK86ckix52s93Vpovk3udaG9
SIWwQH4kcpG8cr2rNAQhRDlYJeSWQdXFMLgAyw78qflBe0nlSyJM/zez+2mwW6vB
h1rVMLGYte1PEdvjsADXCvXyJNqnFPuKa2QVPlcBAFbIU6yXGddtV86fxzfeJhBf
MoVoj2HXMVILqbsv6pp5Rpahhr4c+UfotZofjFlA34eEn8P93XzAConBx+OLUZNv
H959/PsnO4uyf2QiG0R7NgDKVni87DvnGVwe7FgXFMR/E9f3XdLfctS1+Zt5olDB
0tXbLcEXBY/jhZGaV5ivD90MPwEp+W/xCUoJxMlo5EM9TVxlIkOt6pGX7a8oW5fA
9ZFkw8MY/gakNgieaBoKa3M6AUMzHtz5sy5xv/4XRRuoi7AzU05dndBNOLNoJAYG
AMBWrOcfZByo7p7oFzvJV3Kqwh1gD0xlu/uihktGDgaCr8VwqiG6BJJj1DPHMF8u
KhD+AfnkJETkDcrZCmEKlCV8W/lM1UEiYfcoEDu8eL9YAqMUAbJltnN+jE0tvB48
uIGgdi8Cf8nG93OrwazSbwuSB/tJMcfY4yhtk29zGQGtVESgSrR6UHVXICRxt8o1
vYTvAgjot04aM/4po6uA0j+iqHb8vdk0AISrL5TselXMhcME4TGA9SFG3fXkEcm6
8wDWqSYW96BvSKbUZW3egnDcjpWqIqCvsRq0sC/Qg+VkJdqS2s1GXteHsvqili2A
yORUETfH4LUPuykfZQz/BdcjbWe+iH+8auBLqvDUh5yeRQYgdl/SDQpsga8j3wo4
LYKqRWlGde64D8CQqBIVLiHQznuiRFrSrYJ+zmJm9scEPtc3lQQsQf38npj09q5K
EioRf62MEfxh7/KD/Vjpc7e1zHlIykizASWGY/6H7Ollvue3xfg/iXecL7jspUqg
NQAuNtF9HiFEBb4vkWGwKL1nrTJyu8C/Pe9aDr0RS/Y927OOsVj3rzj50/LtkOpa
4zyiuJcxh/mkcf+lDVdyfYndMi2R24F3A780e9kSeumA5aHPYE/zKZ1qwyaNMVXX
7ESMLmaw7OOjooYDKbQIhxmKk+mUKkgu4Uh4DrZuv8U9izoVGmcuBQcSuo7iXMkh
e1kHG1DQ/3dM8+oyHu0Kw7kyqz5tdfSN9xV1Bi685wg+/WXAss+fY2ecraB8K/mh
t8YmizYmWGrgUTI0P2KBhkISnlT0Ozp0H6Kaq0pYbEXBOzPsX/S+XnZlXc1eKE9a
IVrjePy5tCFm4Ak66uL9DGjwcerSXH+J2OMOneKZKM1IPA9hhBwSQMtHAbp5p2pN
A5cRlXBAlQA5K/uL3o80XaVyfyTiljtmNrt3fC8jH4bJQFn9K8gmbgKrihLTmOWN
qwDr1fVoFwl7hg/VEdHV3qNwEEKT/5aSJmE6WQHVphjvqx5WAdQtP1sR76Ndcf3W
Rh+2JGfg5EHvrq6o8t+A/W/4m62Aa9KMe0YPeLa2ZBEVvTJC+AyRbf1Ob0ch8bxf
FM3qjtrB3HpCtRHiICdRgNEeHbn/LpEcwe0r9VDo+MCxaDSBAkngxvN/pv+NGUhf
r2xKnyAy1QiMvBvtN6tofcqe1+4WMnxoxJ1aRYFd9DKFpUKpPmS+ayJSsx8ToQHp
Wc55VGNqUtKFi2E0ORBa4VziSOkecL+ec8nlL1UlYVdqiLCU2jBqGcc6QsmZbz8c
k88gh7ACWvuDp9qRcQtNCs3DYgxMLVhCGjqdJfXN/nBqAPpVlsMToOTwz91z0poO
6UbPHGK63SI7v5rhdEgdsMQ5tOF61PcsaziVpa7G1gTZUD8nWbGDmYFuppluwZ4P
dRFT7/J/0D36fUGORAJQnicX/dlilSASK1t5hdzL5e4A38o2D5b6wdStCcDLBiKK
f5cAOTEXXNiqlBqPU+8yRireM63VlQVR2/7skJ3WNfu7vkq971/HV1usp4mqAqDS
nX3kmk2q5TuA8fD1s7kxcHFqry6uAfxgvLHo6GA7eY9twZ43AAMzhkfLaDfr/0/F
G0Ye5htJITUjn6oAF66iP4MKzGv5i9Ag+tjwURR5xd0i57HqYPIPGHaNjlsX/xgx
y3ORiQLGKTsTjQt8Sp6INk34g370fR1AA8XEGiVoaf1cXEK7QFyIwGo0l6dzpJQL
RvtRau8jetgMl2uc+SLbDEZLIR4CfwXvPxEXqILGYozg5qk/uDT4RNYh+2kOmVze
Gl/Zmi7EqnU8tYme5wlJEm0OSDtqkS26J5+IEpJFp2xprSpwvI7Rwo94kYybDUyI
uaQRB8Pk0BHPTC0CnYKCOMQZnwsWdaTOz0DY0FsoAFAxNQgAeCR/GPUO8jotDhqP
lmt8t01prEJJ1It8QYNyQS37xHBBFoO1rNd+OWYVx7zsBt/PBkjClOTW4sPYu77k
/QE/dXjRPd09jlQI3GfeYtLzUUaPqsl35dqHzTzfalFNGjsOaxhWCZNq3zvF88ht
U1GSKFQMBINhF2PIZQ7MvPypTtgWjw7ioGKEq6YqdI3lke91RnrZBFrxi0KwBaLn
RFPNG8+je81qQpRQMBvY7KB3ZYkHoyFPtSIIGMN9qUHfxBd5V0pIugbIUa0lMxOR
zITLkXGr6Il0n8h0kwf6aNx0KEMBCZSjtbmvut8k13/iUwVbAuL3x6JWGO4vxu6g
cG4OImiPMMwlePk3/pp7W28isv7ccAXl0FewhZs0Fnst21GkXAMquGLOGCNw+I/E
sRBh3UF7nKGsl6IL0farNT6uRwFI0tH3f2EuiWvBUHBuQ2Vos7tppaLKGtS+wh/o
n4sJrFthBXeqUx7WhQqJWliZsiNWrisPb2iiWXNidt0jeVjiraPh9SD+/b0zRc/H
z5z/75Jp8sNN43dqDbN8zPWnE5RU7iB4osAikWGrNUBuNUZJX+0OYcGnEdYBVsoi
TqgD+Ri/WbSA+dZ1QkvDMsA8s91YbiCTeRD5Hlev8QTK5fEid4wrN4/wDu8A2z09
NT2eTdb8TREElcLcWPC7mZuH+YuX789uesEeaYBWpuGcRk+GnWtM1jvHGbAvphXq
Ls9x6YN0QX79dQSu/1+lNHtTyvcyZyqqF3kowFmsFLVEBK7cHKSu9EGN5QmaxmOT
hgaiXEvCCzXJJyMHQYFwihXjHHJMP1tvvgkc+R/coN5BYcPEeLVC47aIwf6j4QYN
ctWemcv08fNMUupzMOmLULYtW0nsg6tdmYpApUfu5RJtBn4nbbNi45jqZ2IgtIYM
PLs62mPd5qd27uvLruW9rR6I+6ifPjkOillraKEkAb+2r1ONB/5lV5I4mNusJG5t
2IENwi1iCLoLgsVcJIxOWjBtAniCs7HK8hrcNl+C//XQ8kIl91LQPAatLpI0QYQI
Dh4RnKArv5IWOB30/43BqcFp7siOBI27qkGNQV9RWO/TLd0odL6tQmfyUcqaFId7
ik+5i1c2XZxt4LKUmi/Cj11H/XVkrY22m1CgIQnfkf0UzbtqtbZmKvMTApJ39MZA
A3KuinqAIgX2R7QfArv3BojuHgvpJyWYkpnjOk9qaoPafsUMWhMJfOium41ktOpd
TzCCJ+ZiqjVNYxBPSWoT3EA4MnbCuSmoAwHwwEzV4wHgOBmTW3dtObwolg2qjSBk
h0dLjn6HTVAgccmCq+QNWcl3TQ5oiShlVcp8uj0+HmTBIcReJEPbhlHNRy25aTG6
cAY6LAN4gQm5yx63jJ4vlGaJxYeVR3k7sMVVeETCqLPc9j2VWCjGMddHOVOaVr4m
XN637iBFVZRRUj1h460LGCq5Wjj3P87eDhyi742sJpVFiJpqxeHiUTV//SvxlSjI
zO2paqpzHd0EOuDnr2OpflnBIVFLkXOO7YYbkN4KxLS+n3wYCEdobqdR+Aeu1z1H
WM+iDOEWWvQRywNFXRGvthgDrC+4dQ3H5m11IYl5H6/rWqrYMOVmqw9wrLsHxlJI
x/PWmOxH/Ba9jLZkCbqUlElpAKboZfORriL8ECDmrOTWTX+HW9gxSQixwgbCsgCM
6Po8/BOToM3W4okdz38Dp7NhEXjN11ArWw73Ego1mcceSzsnU8FUCMEkHTYXnURk
ixS5EvaCx+jaPIobCTzYlqlsCkfgJ8DBxgch3e4IDssR8N42iLzYzjNKurhuD++J
kObUmHYGmtV2NZNAT8UQ81pd290267PwSZJjGL7RRYQK7ssj8ibOU9mSA16IK8sN
o1a7g269vk8aN4FGbsXrXZzO6DwzGEz+KwWlQiSWA/YGmyHn0BSIOneK8paNM200
YJjGG88juz9YjyECkjOVyY5onH+8tGxev/WyFElohhJedWqedPKdnglEXmauyoUv
S8SPPWi9b7IL45t8u1QVFXK3Zn3YPADNswTJwuBDMzHwsC3RwE7ZaokBVQ/U1dhf
YGUIa93JOpQgN7vhGbLB5W45i307U6XfXLRQ1g4sMlxaErVSpcwp/GMVdn4nfz5a
RlCoca5b6Hn5o/K82mt4LYyDRN71wYzr6QoCnxnVJIFrfpHMTOYIc7D0GfQri1Kx
nklTJ7VfYE9KDExDJNoP1Ps7rdyxa6khgrZgpPfSzbXkY7DrdfvGcy0v2PxDDoOn
wKhSTF3LuUMJDoai7AueuUlSDWLyyC7b89Dcpu2b0/4UKLXDvXGRZyDtl9WrzI35
J82rCfmw/ugSsIyIbtr4s2fFiapPOyGQVx0iss+UjsGlbgBKuMWuxcnrE47ra9qp
v2Vr3o/5xvpyVNXohmcj3OvJZRxhkhuz2hN3nZIeaw0nj2WziABM4nTYmKbBIRi5
CcCXGKco1QXET1Q9Unh+I8A2T0MAVW26Gbu2jTKuCA2XvGIvBfH9YdSwdtlEIQWl
0mAE3bF0VezKXDgXFGpLjcBcg2wAoLvfjSrNlDrfai2vOnSDu1ItTDJrzmTvSbc3
CnNMZhPmN0wN+XJ4LcWRskywN9h4Z3RaOnl7HOQsMeNhuZu7WQeXAgLc67S9eInw
tqAJ2xVx/IayyP16L7DF+OI9Lfz3Jb0ZySNtyjR1a0u73Yqtz2IJ1m54deh54uR6
kIjXVAtjppWqiHhyFGsFNdoZU1GFk3+1bWOnyE2S3riIKjobTRPr/HtNMN6C0G0l
nqrhxyo3qFsnIY7/u6mi5d4HgVx+2KXKQUxRmVW09CfVA9ZVmtAsOpdWrL2l5Pd0
H/n+OkHbirbRjjmkad7UwlSnNRYZlf3BYCEhKRSKymmcPxJjitvW+344QQ0QAqgO
agKzc/WkhSvD1ej7mkK9VYZMTXH5qxFZJVoN74NgsKsO225uKT7KTMr1S2nSNz4E
kX+BzrZNUIKQfsHkDc08mWHiKa/cOI6zie11lFQ86vvVa/Ok3K1AUEk1d7R6NGEP
zS3bavpkk3+6bKNgfnBpGVwM0Dxo9tnrUYbXrDSuPm9qDeNfKEWF2PWAmiH3cSqw
Dpv7/ofzOKyeFDKVeYlUhmrdaMGSYrZwbI/YMqdFzlYgrwd/wkxOQBVFEqINSs5r
eddTszHOf01LaTWsPozxmdeycz0Ziu1ELtZzdOR2bTxIEoGk0H1XCxOoykiOIx6y
6N3237Y5jAjRaTWXOtd2fczl5ifRHwbfW1KpFmpLs6MwkOjhe1rBm2EBh9YPoj4R
q0lm4IUxWW8MxyRfKas+F58IEYDTgsL4+ftDG9zeCkTWzqgPEmt2ux4r3rJ3FrI/
0VMDxuCymwnQmOVbh5b3nijxqaM6zj25uLYQKI3I894ad80qk34fdf7YK/2LmHKD
1J9MOEChRHJWblMLtcSa1rFe7no5GMeXlnkPdL78CYQCcPB/gR2uBIXHhP9s8CSY
qXTFbpInScmQF9M2k1/mOxNOqX5v3mTReQOxawfuUr8pUqgbj6Wj01RHsQ4rvtj+
G1JthlbrRupwmAvPmpqtE97Spd6H5JZfPXHLYNH+u/Ym45GQxB1OVQ3bi6DtPBVN
8RTnFPL/hPeFvN3mON4BUEM1aCuimzpd6bO8LePk48mb/rMOdAUaEtB6H8Cu1Qc4
KRhpA1qjiDKZ4rnXz5uZGxYyx5DPipbw2XKEP2fwjbcPGAFKJRDTe7wi55K9p4VE
dCuR4SJ+RhGukYLP4lY56M3/rLEsxTwrEximjkXlU5LSQb1OU7d4jDPw7XkSFlGB
Bgepj3rIEqcjXlyz561lDiHHjQ+MZdgVK9HxHWbTgKDNXzjgtV9MCFBD6sIqqa+X
dTWBvSoOEV3e9OUJZt7JyQYEQkxUzrS+EdmLH7tE3ciOlrDDc5F/EapcDIWv/Rvt
TEj6dZbT/u/gj/Ejgnzze5EnFTLNjqIIAPZGmod/Z+z4TqnH3y9e04hyl1GkfMlH
ymUTzai4aQhs+e0nSwSU/gZIBza3ih3UqGjfvWQNhXPHItgLhqghdah0JPzr74I7
pyUhil7w/wO3Dgd2Qfsc8u5incUMae/ydAEHK/nNE+VNgjCAGj6nWA/Ko8jPKNrG
4U5ElAfQpFJ76sg8Io6DQt6WFb9sbV9GKfokL9bA6Xm1+VxbYxSbw8wSgG3lvvSA
OMCnpscSeujjYYTFENVQ0+mlVWG47E+dMU5GeMANJrxPR3GEo9DFp768Z8+x+fPy
zmycT0IA9Y85GIaBotlrOegC5lK3opJriUDTPgL6zIBdcniKFJATaUVq3P/aCXfy
n4UQWtjo5uo4BG/16iPTQTESLnDUWuMoB3OcTBU5EhLhSa4jxeJVWBPB/PoEJJpb
tZZu88FnbTV1Gapwd4yLazBISGTQRcU+Uy97OPk05act4mG2QCniYZgWReWFQSHv
k67QMXp93kiaFNau1Fzw62A9zj52DbWl6zGjC21wKF5YIlx3JxitQov3UDVYQsIq
iBAv2eLcOJtMVRkCII8ucnlcvN3qC2dMoS5ijgh+fIWWfHyMM8OMAnv/kM0+7Iaf
RKdFQeba9CZnA+Cd8dKgx0e48GCwo7jFNAQc9NWPpjzSmjiMtd03nBZVdnEuJyXS
L8S3aT6mwWQWiuCtJJrmxaoRDyQABpTcQ1UL91+6zFMJmbwUjCtV95CwWSdyrrrc
NnLnjoRCxRMayVjCMT48Hs34WBawxDGsMg/VGKQ00ArG4C27JritDewOm/kDixV9
1ugKQm2zM3g75ijhu0dAc41zLc6ipiuk6Q6r1RZXY8DdJLEZJyEyY51Phc0eVhnU
LxWSLfgCbfXMym/Ek4pUn6g41xzheM9deT+JYagMcFLe7wCUA6DaaHcYSIZejiEL
EwSX2teka2H2lNQXTIRD36cMjRDiPl7XIhLu2wNJfUZwUNCHUTaEaEz8JXoUlJ6o
nchijN///ByLO/zo/QTBG8GecfxTaoiPJnD61iATnGXpFuINrxTwwqagxC1dQr8k
9b4GbsrJSnfalrxocbEV5MjceUioBYSV+PG0GqrRvY9LKvrxmgNWn1uhPZo8K1w8
NB8dJYUTiUB16DNfbtKpwlYRPPMLC+F+xeEFGH+v1c1r++GWqT7skKAheZyCg5Sh
vrlPWCubDn/kJGQ25S2FsTL0MRSHY/LUUsLUYN8MOpvAvPXhsFBGQpv0i4TZ/RR3
ZSg8ZDtly9qaA3Bew4S6a0tUk9b6Knmyqu4uatbEZ91skqCbBsiPMMwhATPA8PjU
7+7XTso9lTxv0+7BaWx7GkrvNG0qGzBFcEVJ204B+4yp498fkKH2C0izerhxVnK+
+t6RPzdEz2wkfig2qNdnimFaChLB2W+4+0j5ytifx67cMybJ+EKk4HjA42cFxMmg
qmY8QMKmQhEAyZW7U8SWNrKkup4dgJonLFRhM+DQdHJekd7pt9kScOZx3gCQblWB
tQ5ozJILkYXl9hnWmil8iPMtkJjjWK2173mFnw6KJ9kkZLXYqk3DMv6nuWnOueqV
iDFWDe/ELn/waZR31C6xPOjqiXo8LUUWXLB70YTOxHA+6k/wBXuAFOGVhdWPrQG7
GWImLhdrqAQVGyFEN1nXeA1tTk6KFEBGx2S3iQ4s4RxVX0WmkdEvlVWymP3c7wEl
P33HiMLtaF1jSuGPBtkLCkFQmyhI+wWFJUDk3GAzJlA7bFqDOprtMK2VVqtIONX5
Ma6tb1cqSyFYAXpG6+c3atIV633gjgyRU0Kvs1xhbOTBlHZzSeqFqQkLlRdKKQXG
M+Bipu3BbFbsxyqD/vAPEJdP+8BvL/OGkp5fcoyZcCX9IoWLpUjWa0JjeCtQTBvf
qxbk8NFyO0Oh+H2j8jUSJ4DhtdrW/XhLhHUy0uQ7e8af2m8fuxOyyD3tAiS319dQ
pHw8Xyq0zSkUu3dsOJDq2GlW/9IIiquCtjez5xvcXut2z8TEvN9AONhhG8UW5pZ9
U2dct6ykOhqss78ScDGVTuz5vIA+Q79b+oGgVYTPljb9jm8H9IOIF6IAjj3T6nGz
gDHuBpwJ4AM+35j8hoakyPluXpBTv+ccB2wFnYmyk4ghskgFN63lyGst3ld3w3OV
B9vtnewOrkn4F626/HBed8UO4cHD37VozccWlqD5DrrUmbgLoFwzTbOqwQT1SPal
/M5k1oP/IqUMHGo6ARFAsT/LWy6pAnvmTkbnrk5pkVhlVUlKA/Og0WSDFx96F2uz
0Ni19UOMJ9heZhbqQlfbmwoWuFxV1mh/unI9SYDsDlplKEwjzwOmwYfW4GxbsztB
Qr42doRWZPhc33bepslgTAsKl9PXumCKfTfRiyGxpR9R7AhV/EgZ47n7k7Y7zp1j
f+AfTw+vRl1FbalEBJTRiP8oaFGI61FNTKPCUO5GmManhOsRLrUkNBVwN8do8F9r
feIEoGZ0HF/GxwEubgOt+0riJDv216r6K1TD8qkggqHubQwMCkNI3V1AfT0RTlLJ
9GgAi83nUk8jgcOzLZTXcBUIwjTR5EZuKEdzC3fKyjmGlFdw6qrwrjMI6oyK/yyE
6mKJUL6N47yQRVwfccauUX4OKH/T0vBWtVgwpaF2a/9rUcYk/7gRjSxhCdQ7/5kS
MqsiQnn0/h0vya23C46NYkHSypfoINCfXod8eywnT7W5ji0MC9yifoeRb5BWycGB
mIbS0bQ9L9QgY4o3NoS4ct/rXQpOdmSUDATZKU9IKpAUZjdm7Fw/pZ+bCV19Bw/O
eLkfIvEu2H0tczn31Bih9dmg+cq1pXx1PiaxTXamGbKhBR5+e5v4alXbZpavon55
qOgzyxkZJ1hHglryWFiIk9ZY3TRZfavdhCAz45vh7f3ZQ99tPZeP6s28rmUOIuqp
+8cW3e1PjUgbWt1XJoLk/1Rhnp/+w/11tQC7586HJbu1d8ZSNFAsTyFscya1n0Jx
YN12/8xtnEXJ5aRZZwysoRvr7rIMOC3bPavNiosEWo6QePslOwb68XmFi4Vje5Jk
vhi6HcZdSkiVxmwjFv96VjvgIzkvizTm0MuQlooZrO58hDBPnLz1IS/5t9KumFXp
RxRHGm52bMTItdmx2ydWz5AykjVEZMV40rWvtKdWR96GEMFMJbr9xzDN+I0gBB/E
aGQBiquRFbvGZOaNkYiHCdXzLbGMsbv9+WmrLhS5p/AYRKS/jJ3oE6Cw9Jos0ER1
WMVf/njC5qGHTnisexLKXSX1QjlRA1gE0ujopriFbx+t0cBSGGz2GxmS3eioqDOY
C0KlfxGecBwYdMSzBZh8p/fXg+AU16N8p5Ku4PAv0+IHNSZo9ZaEF7Hz1lk8OlSr
SOrNARobcjP01ac0WAtYc5tktCAXnLvy3lFAVw3dflkLXxlAwjcg5AnNHb+qjjIX
KJqDdoOM9xZoVuf8mxqKRUSxnKbpfRX9sFysXkdV5cjVYSuZN3T5q/VmDsLa/Obe
MBQV7ng+Zg+ju+iF8ur6FN9Nh2bP58WNjZqu0Tijs86nFF6T+Na+FpJzpfX6aUrJ
5OSyXxri8yVY4Cq/hBD3koAHUg2hmAroFQZVe3SGE8HZC1347A2Ao2VFvw4dD9kd
rn2LNjA9FdL3KFd9hP+AMEjW1KAjr2yC4NWpR2KI0qKpmvqZtu96NM+r7tJN/y5V
TgOx2lSmGmwgU8gL/XEktzfU1Qsydzcsdp56ZmrnNnKA31JaSJvCEZk3iE7bIc9F
rD0aAuOqRLpmcQTHckDGLDXG2uWCdzHNIbkC2wAfOSzys2ukNyTFNaT9JPqfVI/R
iseT9jUyN8V+nXIcF42UjyCCde67jEpVn1qsGHCyxK3r7OXxouK8bV1MvZQHetgc
vWSoGc/lzVT1N1ogkzdfX0qj7M5aefg+WInvuCEP0agBxjrD3hC5hrgMd5H49vb3
zwwPgVInSRKmX7fPJ1oKnxjKMHdSdSz03swfNP3C1lEpgHC7nFHxzyL+ZIYT7Fhc
w5Nln8/gNwrrzr9rEwm3REq/1PJojQuVpfzt1xzeytJOVlMCEUOJgNS3/leILpjD
pfdWFyF1HXhL5z8gvOmLnTdHgUWaTU8qgLVTcVuSJ0t2g9LYIHiYPA3UFJK6wRw6
tD6BoQVEhjcYLVSWv4XLJrRruakP9CdvoujJwUL2LLDF1suTfSEITaK7UkdI19Zd
DBOGt6tbGocV0HbXC2/dDJ6ldTHxdXgtF+B92KATgP1EOe61oUoKkvr9GTT//MH/
5uBIVAH04zB59HNtTC5iFMmPofJujZcMmqplj8al0f3vQNNvXPZFs4a6arI3aPG6
dQR4urxLLf4dSHZ2aYgkjSsOR1ftC5+rUQ/viCRlHzxxSvGF/gaGWxhhyaPaISK3
AKby6UCriHFJkSOIw43ZtM5XlEJzD3s0y3YLbJZByvyDifw6mUY7rfep9MbWSLPa
T4K0iDKNKeKFuJyOdYODxah4aOwGteuYTcN7z4PgTL8hHrvkTAv9ZF7UcItK0xKF
YShSHbgQUtf8VKcUA1BEdGvLcndoMCsqB5x7hcpoSi4pBZ8a+2AvWfE+4eG+UIaA
8ZRo1g1RwY37u+zqOUETBPdL0dDVMzo3ufqNck1GRTg4vsglovavwacZuEc8Pqcu
lWYBTweuXq2/n0oD+f9H8xekizKD91ZrXGZkMwhUmEwatCtN0n5rJ8q+8U3L1erE
Qn1a4UxBJ0kOZUNTd5PGxCd+LiTuc3U6sDSIdczlo/0HDyuWZTh1LL6ckLth80pe
zKuuZ2RB8aXZGa/aQrNDsyOb6boJkeRttgzJgwyUff4gWkr0I2EyR6QwBqA3mrIE
R1ScGzjtp8HvJ3LW965DnkgwLt5lVrmwwa9lD0F/PyGualDlUI5Y4whX0Q7ilIa/
YXNmCzUylr2g3354KFM7Txj3xhsN3rUrgteq9ygcQHBpVSEZGGr9QMrbeXbO+9Ao
Yq8pDqOmP4rap9WHuyPORUTh+TSfOG4EuwNBk4vH1ZXmI3Qd/5/9pFhCYJYiA/81
L3hklOozQKoO7jXxhGN/MVdKudf1judDbGtfrvGFyFEA8pvraKpp0QuCfiqwP2G8
/EjwtxI0IdQRsX0L4NEhl0BSZ6j7ANv2BaXbOjUibyClpJRj0/Y2AAbDOwzm4/Ie
HzI/QBxeP0B1P+q71qsAVqv9k8WuhurM+7i+V6AgGokLi3r87PBC9zOKoDkPsF8E
SFv0y4us/6hrHSUfRENQrB4jyo82H3HNwl0TqN+4utm7Gx78qhbchGldziJuvQx7
E1HLV40PuAGTBiwWl7Qo09n9ieXqmy6kVX63q2c1i5KPQjlD0c/hPzipXcGZIRc3
INb7gnp4IpVFT1Qq2IC09XFuldNcU+3c0898rFydk/XLVX4v2W382PW2tj5quE9o
d3Jull0bYqqCgNg5dxvvc3wyQhjDJqliALORk99pcG9zDv5ajlTdqewcELav91pY
ZoJhZySsIg2C/PlcJQxhwKPUDKRpf0Ruuc1014HWexDBS5rPhHnoqnQ4Aw6ImPMS
AHPmsM5OdxarFcqY3NrIZMo8xe2syUYbBNksDiW/zsF1ylPWW1aNAXzv/APtlKCd
OWCD90alvj8Pmj58YobRIMwluwtFvm+9pj/BftIGcVukmmH+eTl6Z3No/dVsjiA3
leGx2iVTfV9/unV3+cqn09OMwKALODZTJNdhppi+1Kyqmn0/lfveGu6H90eIKXYe
bvndMXIUjempQDmFEJxIwNMJHgZDRJalSs+TbCuls1pK4pI75CPPwnty581ZGM5E
sCD1dleMuKNFMS1RGhUhqZqnv1VrG+r8C/PyjYbzc2YzrWNg4MBvvHO+iYmjjmqJ
HKvfrpYT+sW4oXKyh27wD+Z2YWsOYcjBPKnS3u30nPIS4MpsvPhmbDlNND+QhgAH
rsZ4b0P6YE8vkam0sFRz4SRVCfG7gXT2o6QlcAxgQboSdDSLGrK4NytvuRcGlXVk
jhip5TxbQs+Q5PnIuC5Vc7OvCsjBnfTVmwE+JkECa6mAiv3soJ3uLxkYPOEAo0mY
jNiKLNAj4T45J5ZX0R7gcvTIzIA63hcRAclz+H/C1JHVwEckchXC+nzClP3xhb54
HGpItdHnLHrTszOiu8dVoMidrOZV5Mr2mgfN612S1fn5gymbsfLox4EUODFPw6eI
781Uah47xdCknKq2H+GBBQ0Cd9kUDRYubbXbT0X75AFaAxfnd+uY9tbyUgQF3UNa
Bijgq6vmPy0lPX1jl+yvrr9DUQkur8SpGEdIo/YQZG2k5hie5dpGxau/Fwkt+qvq
6kk8/H/pPHfcxigsCgxWX2mndQcaWUomzAWi9hCYrmSyXDtBl1A8qkuybuDYbf0n
dNwED2C/TNUDWykbh92xs6DHJHcbrc8fT/pQxjkv8tB+Pwl4nL4v+62wmas9vFF/
2PjH4cgas1nt88bRxR/V0KzKF59ZpLTrtMcnjsyopDJNCcZ0LY9S+lxm4LC7ZRyi
1BkCTYqZPNqQphKhZl3Ql40HvSByXi7XZLT9bWfBjqn8lyzV2zeegf3iHsjJA1C1
o8l3/fOc13BALl6ILYHgeQ==
`protect END_PROTECTED
