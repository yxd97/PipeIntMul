`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4OD91Gb04w/5/hQR0HUarZFcy/wYElxU3flb6c9qXj4t0tcYFYCq7VaXj3KKWJp2
Ic4DBtGzBUsSiePHqgjU4lRr3IPDYtlRfBCuIoFedWYTVUNuhdRdCSoY3wIRG6Ry
KYyAXtHyz7ucrlDg7V89m1k4JfXe+qtzuNnc6LTDxtbAx3nB8h+pZstfu06vBmOn
2IFwTHqAZS5g1AUlcf+RyZiqhkNz/9u3Gg4/uiW2CCR3Kmjzx9pImUoxhGhdoEsY
LKaoyR4o10+OJoyMJryYoNXeNnXuaxvbAnYj82WrIYABbkEXcleJmzfJNlC762wC
Xv514OavnKSqkMwEd7csXdTJqmUt5QNCv4o/Z+CYUFHLW9ewuwzzLrazRPi9F3b5
fBWBqxvV8yFj3Z0WZoc1qQ==
`protect END_PROTECTED
