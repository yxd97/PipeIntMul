`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WG5f/4u8BR4Q1DjSKtDxkJUkxPQQ6CxShSvNyneQOwbRFuz7OwhFUdmYZaAegLS
3DIWyoHSEIjiRMRb83nY7P7L/FDgUjFkiZXdhvWVSMEpAyyvzlXCZ5/9ud8dZJoE
/Dj6r5Mq2PZbfXehx4YU3VIIL1Pk1Kh1Ww9EYI3paAYQZdQzX5BXLPMC/39VRADv
/3SjPFkR5BFkUqVrAxcQFJn9+zf1gpQ7B4CERzaBZ/3CL9H0JoSlzBVBeMWRdDAi
agDX7I7EHoSfFa+ME9n+qFaPsCeRHAGrJMqVlYegcVCHEHYH1r0bOve4ux+LSztr
Nn/owcI7eI8nDbYVBRm8ZvcbAMZKy9PzNt0zKHByQqi0QvS9iE5aECYJUHyn6I6L
iQoNdzltrQXWwYgKBiPFM9NbCYoB7H2Qd5DMLmK7t+4BMpzRdm/XPgb8NzUdoddq
QRW7bor4SiAn547gN/EQu9OhHvERxWHtG1790+V+T5U2Vz7Yq4JJICnLjYnKnCp9
itl+LRSRE4K1NNPCbUfdRpNer7RhZJgUU250jkQbPLwwn/lmXCyX9QDuF/OZYGF0
/9+14D84QJN4mTdqB7zY+8VVgsuxSF7nCc7UZKg3RUh0cMXXzaAO0xqPUZPCSOxs
KL4iZNnFjuLPgPJGVhUGDw==
`protect END_PROTECTED
