`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQUiM43iY+aNTiP8AC6hFoj85MDd30jT1N3WXW0SB9BFzwfCJ+QZmk0txceZTsAs
5HmgsEOI91e4v1l/Ar65EU3CFzjpy6aqGgqoVBBG0OsnC+CBhEeWOx55kcXSk8W8
yMprt1c9l3DVy4Hdp2Ozfq+B77M+hRgVzbJEZLjT/cJqIGdrcNh26S1KLlXh1eGM
9yXbhd48iOaDugQCduL6opCZCzhXSu2V9lXAG359cnJrchXn4hs/JsOJWU5DrDDF
T8TIPowvD6WUjcelL6d0UFV5K4oBUzlUA/JG5egQCIKxFi8Bd6ThbRmWlaGOfIST
MuKQz17lnVbjOQFp7e0xjiUHy3e0dMJIY58wNeSjC6VkoyxOtt0zNAr/WwYtL5+o
`protect END_PROTECTED
