`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zs9oDrOJsog79piqKFzHXbU2DY0SPcPlAeB60Dznx0IR3uMXTBqZFVarzLeTo9pX
pj8mBfI4rIl337eT61eL8ZFYiK4ihzaZog8KFHXAJjbSSLUVZp5X/+JlymIuut5V
HriAUZ54I1Gaz8NjzuFpxbhSUOr+dZYuSJ/npGwsAPn3TvHrMqE9+3mQZeDOsyO5
A/E+BO1ssXDnPWIrdeThoOfLbKADoK0mV7QpwUUfk1o1xqgcDpWyG9IO7X+khLs0
CcCjP77hkHMDo67B9X5SsJebUiCKlA8ZyYIgkw5lg0RDIMXRMtMQlWlg1lqscxPm
wMM71bTF6yrqd8jlSHhlUA==
`protect END_PROTECTED
