`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uDsy/ZGi0LM7ycHeuYSoM6sDfcWHnLlSWfcdF2M34CjOgqIi6JPeqzKAWMG2RZBE
bZFMsJhnpBcuLhFXqv7LRveqj3JEoJMfpdJal5DUc4ZwWxYMwyCPDtKTt8ODooFy
aiYVKm3FyhUqFLTHi7GE514CaAxKtnjQgM2je3ZNcTy0ta5VVp6GZZ+TrRFuYja8
22LRjVOBEUASc3AXM0Wzl8X1AeIo5j2g9Od1Ts3D1bHsfAIWAGvOCeIBB7P4Xk9r
wnxTKXp5RxzFiUYvJ7NzX5GotpGB0LnTxnufclQiTmhzsZaYBFseRzLbRXL8841n
zN4r0z0R/iZNAfi4SFXFwSOZbBI7+C8WEBPxAfECihU/uIvP3RA+Uv4VwV/xilD3
RebKyjAk+PqkV/BAlBQfKR15z7Z2RBW2cZni8IT+3hOZE4TU6ocrjsWCmtslK/QK
LgAIm0AzVLOLZ0daspnEhQTmdxJo0pi1TiRLaSZtUfw=
`protect END_PROTECTED
