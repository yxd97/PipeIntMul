`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vrjb6sAGBNyJsZqqL1XpHBjaF7WL/QuAPXQ2iwksp86QdwYTmLz8flFmn+09CPEq
cyMFUaopA3x/WDyk1myVGvBEubdPuWdl6Zw0fq7/Y0kUGG+DRzmL6Pq23hd98taI
KlPSTPjfyYziMN1rZt1PGFQf/QKkwhJ9dWTnjqQju+GZRygJPTunTtSpf08lolTS
knye1T8VuoeJZem0pSrrOMHve478bKNymBR+zx236UJ3fyBbZ8QTsoTNoaJ7P2ON
5TaQBQjcStS1WQ3BDINjRLNyxY2tcQznmR62XutjWwOXcCnw1Inplxj/+5Tg8HIJ
OQnjNJLa5ba12t6aEfF4lRP9VDk0sBxv8LdrLQe8PXE3z62ZrVXbUSyu3f5V6KsD
dDaD+JNwORmHsq4d6Iz8NfdO5IypqY3a1dpV8RB8z+VA872GiqcmIS+sBgiHVsrq
mllrIssUAaD8S9WDnhd83MjxO0tMHGbY03nXRbrQMDbzPNWjFHdk15oO6cxrz+4t
eTsVe0gjqRQYRsl+6VzKPdX1hBvM9Xcu/p9MlgPWOUs7JKvSW6KroOC+gUaTjdW6
ySaP2pXPdUCt3WI/43TqLLfuKOnEi1fC488S++YxYVmsD6K8WW3GA9o1psFVfdWf
YmRQZSRn/k0usDNBgaDj2aXfHavkAvsJbMGM/QlQUny0YiYuSc6kEeVFQXr9HFHB
rR/X4hOCpr+b70Jx3TqzP4JxL/cDgk2eNOv9M8yNnZGAipmkmP0RK0jFfgZBRrG3
DJ/EoYljkkSsSWSNqX4t2Vjtbme1Pf2oAsdSBH1/wJ3GR1F0q3IbC8nDegMhlSzb
MOe3hgLoI+fmNTQ5sb8wFaYTDldAjU+JhkAZu5520PHO2oIrtRzRwZAiL/8CZHGg
qiiA1ayi29yAPuNcy2vW+A==
`protect END_PROTECTED
