`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pGA6IYqrRKFT6123YxVzMilahr+EjQwjHeGPu0a/EO1VTgmVU3FLGvTQvt2ziV9N
sqlxCxiRJLXK2H+XNyMFp5KS4Zq+PUMWWBw1zWCqerUFNvx1Ovhlr/OhUlD5CELt
z9lw6RkfwG8PjjBcZpU31Gw0a3k1jxTjRsQznFcXlfn9Juur2IZidMk8kSjrjzNf
jhRTOVjskDBPsPUeu1r8Ox1g15XfKzEmVe9XusfjfrqWBIZ67V4pOf89D+RqgBhJ
gUBVPX32/EDtTXqHzdnzwfhQfM3vMOUWT+pmWfmPgFcLhY2isrPB63uJra8+TJhe
rGNRQf5PJWVZCWhlk8p2fohyitTTgO15PgdjGwHboCBvTo7hzkLD9I6+rX5SUfaT
4rdQ70wO1lv+IR+WVe5JWEtg/n0rRdrmQakODQpfFs0=
`protect END_PROTECTED
