`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5afo0PorXZP0YQk7/KPzrsighHclewwd60xyU2ciq/O1/mWTCQRz1aLlk6mSd0fg
LrS6ZnX3pN54cSyNdspFPfItBIrb86aBJ2o0pkc61T4sD2Uxa+YIl/0ySXSJcuAg
kfNEoXnz1qWLShUG07vnjN/z98RsKKGMtIynEq2YiWS9oXzrZXL6yZzHYcaj0m4r
KmHXhI1GzLiV2oMo3bF2HMgQupU7i+/I1O9vq3pOwQ4buy/Q2hUcAJgbLDHku8vE
wSCyJl8HPEbiOqRwGts7xZMMvbr6XRZMVEFq7ycQBJ+n7xEA7Nd4S9KAHYoeYQ4d
cRiIvAserZUwkWsNmT3eXnkqWYnxKla6lmdAg4Bezsl+nmLHfbERBG97MsVIfdNk
Rx7Hlo4lWaCJiqNfwBeDy1d7yIedhgAMF2DGKKmdQzrT0+bqi4z/u6QugBn3uSYr
PtYSAZiFVTKYtiQlgqfEcmMRW3s4ONpzhLOl5WvJD8TlgiB5J3nLVo0uhtF53Rvj
gR/g2iAp9uNDD7LtBwIGps3wCwZ4MIxC13GW5khgStI8e+HdJdFXFxFDNBcSXuj2
`protect END_PROTECTED
