`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GZCH/Af7M7nGHwkHEJhDPUJl4LZogy599FFmHSdRxrN0OpesjMm1S4rHA5D/ofjT
sTPS5c0Q0OwXQ3S3sjioqKS4X2eXN2e6nbxd/OBPhbaXmzwSD+Bo8ouKNLCn6H6n
QiTF4zQMoKGT/uw+hmOknv817FOMRW30rW2qzbGM8ccAdoOInl8VyfgarKKKLACJ
Oa3eE7n8S7ljwuwKRG8Igo/0sykVhtvwWDlx/0qGrPLUgYZxcb9xZv/MG69QG+Ij
Gff1LZMKPXd+C+Bsrm6hrldgrAznBoHoGo3n4+wejkOvPQd7/0l1RmfuT1ToSEfj
OEIrM0vLgzArV3BXhFU2AmgX3X5CDOPLcJdiuUw/Cy62jpxzKsnY9N1kRJUjTAAw
WmU9Lz7/+gxugDxSrYvGSNpyM0S7/qT3edJKDM5DnxoA1FdB2iYdorY9U7N9uYA9
4P6W8MWsadNkxlUEYa0lo4NFOJdk4TtohCQ3sUK13WY=
`protect END_PROTECTED
