`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wFxYswnr5U3RDunw2v2uvuSuh0A7EX+mzdM6k53m+JPj8AVFMnTThzXwMIVRD9Wk
QMIsLYUeeV2R4XxUPF1qryMavawbj8DJAEN3AEq3aUPR07WSU8NdO6ngUPQU4Z3C
oCzpJWYfasDaL+ivffRnbXJf7cbg2LlznKDioHTjxqOrBK82zsRCR/tWOaxap5bp
3KNOheg8z+BifRj4HQ6oZeWgnXCC0NYBBN75WhL/eln6Xm3qpsuQ6q9zvS8OIS7F
Kl9nlNaWbiAMDyqxq2e0YHKg31e7Z8xAyjCPg3n3XZebERJt7HxBGtEjRevVfsEC
U7KJqX7IJDheCwA1ujN5etBzI38bBf4e/gi1L56SAjpz5h6Q6/GeNzugeu97M+F8
1N6NGPbGg6bPUUkLbZPEB6gv0fPx7cs62LPkSO3uCc6SXq4iOsGY2DaBxnuObvfx
UYYY1anX5jvR/yfVy4fVYLU/adm32BC6G37HwTBx7gYZcFRqZDm6IaWyFdyQBTsM
/oyY86bAVLC9qgJmb7CFlgGnicCpXw/nzQHlPF54RijykXgRYYfmkTwIH09gIYpn
N0g6grXEkFsRKvszK9c+ntQYPPRzamqlmgffNxzMSE4KzOELxsSGehnbbIjBNPWi
ABTtXJWMyMnWOm06n4mnFyC0X3YsA7G4y3mIuBC/w0cnpwslKokr+RZXIqSFE6pl
PD2+kw9vvJXHr47lXxYcFvGgkUtKggSMLh6u+i+RpFq5a/yi5if3zqg1qPWhOdGF
UzvCCKNhG30aY0IEJb3VA41kVDxxPc2J95ILEzLQIDmbdwqEM/bcIQp0aVu7Xdjy
syutKSz38AxlquwcUn3ajrlU4KItV3U2SYkXMX98g8LPHRfSG3R2otq4+Ad2iF4G
mjgzqc4l69t4kEOBVL/W8lgdc5kKeYN3v6cxFdPXJr8kMtoYqNTWWKwBmmV4fYES
8rOQ6Muao9jzQn0+F5GQDBJzn5WzlsVNRbaJdpjQ46sD6074X5Ri9tXClfWeH0QR
YjzREHZeJEBVh6qQEh5DTHzsk9zVqi6/KYXTPlXEYSNZs7CxjGcUJ7pGmh7XqLjR
ZkzpSQUV0VB/QDUB7B56pmUyImJgcP488ElwOf7pDZnHlmnd15T8SNDS5fiXgdnP
x+EO/0utvaKq5nyEOsXwKzbAn/TD8n+ljF/okaSmeSY0+EknXRGaf+Tm0dJQTrO4
JXuP8PGsF3MinQ/YjMxqCmdJEwU5mYCdCTxMOz8adpGvZP4q7K4/zWwqhYAyH/ZV
S10WsWm0O0603i82KV0kd8TEgpHw5jSAnPzjfgI9s7l0Xp/iu0o3s9kMPL4dFWv5
N8tnhGt3vySUtdkO5pBKL2ccEnCOql1aY5ixKbveqnOhJLPnn+gYv7faRP/llgVR
ze+IrtowksVq18pyWn1xg+jWfZN8yCWgGm+kJe00bGFlT8rfigbd2aFDsaHwuh5P
/IFAeNPfIezzEZWrRkItWUmz0TlGfbJqoMCmmwG1r6TGU2B7BbuYHV8OkvuN7Fb0
JBN38zvKI0hSPftK3Lo5HM4YPwcE5kcqWgMsKcMQc7k=
`protect END_PROTECTED
