`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pULPmTJSkBGDgX3t9MXihytc/McX+6ch1CkTpFij1YMwjqZ67Y7of0WQTHtI2XB8
lriwFT894J7M7qDH2+E2QMPREo72YAx86uxOZNno402NfE/fkCng9pldlvOqbCk8
ONcZBqmcLxaOtTCkEa1B28ubTE7ezBnZ/czyZxkT4TNgoJ9ylAe4jdDh03mPyJD/
MfWwp/khEBIcF4vtr7u45IyeGgKWbW1h0qhy2qfxl6jzVxLMASxXcMkbLZWsZQfs
8zb73SSPEaUs8syIAfIlJLjA4Kp7MLgV+aF4WloaG/kedWJxk6ekUS+DbGoNLE66
ZxLNzqWT66OW3CUgacXDAP38F+elzDvPdFBe3uWx+Ag7+QIssXYf84u3LP2PCr5B
XfUoLQbB4E3VQq7z4dOjEqMGKzNaOvwxA6K0KP5KGyKIHpSqD17YxpT74owaCX7P
K1Pu7ERPI8jY6rm4bSfPVx48RxV29RzGACH1qg/2HxWpZdFj3iJReLejQ8EmePSi
2uFPL6s+0U/y8p6xOYGUZQPdNjPk+UovnUWiRzu+zHvEG4sxnE042DAESwQ3wMXT
KASHUCtdze7mSs+x7SzlRz65RUTHVnKFf9auGJJf7/q6cgoJFE7ftxXKJ/osMPqj
QTY7C6Zv9o9Dv6jaiCYa/ehyMyB4lcVLjoUhlZgaJZjEVDvErCA9RxlDGIW35asC
fpoGmEXdb5WK9JitGjBCqPciJqqbqVaZKgHn4YGThVWCPjBFa9/MXvnwGHYi4kVX
bMAottwVwdaJuItZiuqPJeLHfGDdybHU82RY5Pw3tLPhZtND8HN+wZlIE2lniyum
lHkgcbOoEXw4EWj57DVM6HYpUUmrhKqGFtZqa+BrMxB23gMJmeG0Ppvjuj/welOm
A/kywVB9LzqMJ5PtVGN8jXUzENjebzaKnkjXTpw4ytA8uWxjobP4xzUCuPviCO23
0IIrEaIw6N6CfVMSgGsxASiEN1DbRjv8OZ5XDHRVdUc=
`protect END_PROTECTED
