`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ul7J8XXNrIvkJ9JbRKnmnTP6eYoeOqX5TkXK0j1DSquTjLQu+6sSLTb6Vh8hqOHj
tFf86aZkR5Wd7FjiR+ZPap6NkIJxq99Z3u+7yOMZJSXSMu64c3odUy3342emYJMq
CmvAr4A37uoyQV3jg1dI7CHynzVxId/TP2Rz9WwVOgE1gHkEsju+tkC3HoQ0Tr/9
Ncs3HkwsH8ZFQ6c/Ki5LHRC26z6f+6OltFDYcIh4TC0ffaS60/sZir53nuOtvt3V
TGF5LDlmpdk1+I/nA0FiimxM7OAkFwW6mcZUUXgv91eg4IEb7vlfRQg8bNGSL2B5
/vWFJl3otkQ1yR4Br3+KpTzU7PZtvPbZswxLZHT65XLSHOzkGVPWUdfGoI7W1MSw
JD8wCWnzidk0TAbG5HFU//5qvbE5GMU5ocehfEVk7kK5x3BB3QttIB8+c6NDxXul
`protect END_PROTECTED
