`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yT2xjaVI7beHquJPUPlOx1PqEfXLP/mT/T5ovRIeatqBXksQWkLdod4RDOxxAgi7
HlIm2OBm+qCpjbQ+IlZTPvMREFU7E+sP+/sLNDxR/q2RkraZCAPB7Wrx3QwIXT0P
pqWTrRTrzHugyPlC2ZPlITUnpZMKI0tljRNsoOSNuuEOv44ywX3xB3aOHO4H/9SO
W4rm0sL3QvEgyaIhNY72KgnaJv4JeNFSCOfqpR9S2VZmNQn8yYMu470kX4deXuP9
eS0BfY7XEoL7aMNIXxOA5vFl4MvMqtv9q34zn7CG8bnH6pTUAqj6BaJe1DeC8X6L
JRgODa2bMpTEJCm5MW87TlG6A/6JTvmGeyofpaQFw+vFL/K6vOzXUK4P4au/OPTQ
14rz9xNmeLSblj4hjQPyfAVwVsMoPu/MBN4p815/cY3jMhAcEU0Dx/y526SlMnot
y88szU0dVHEDwPyL+Gkv3oTUmNqwXK2LDU8fpoWjIOsZhL3Jw84cseBeLNOsAddf
h1LYUB5c1cUzfAGFPuoefUgWPdB++a5gzhwAd5QZaGR47po7ptODKEuq3D9iYEKR
LSNa4PWioJLE67yFwbvvgCi+5R1eHT8ITkzu2VZ9xY7PXYzPZfFXZBt1VOq0L7UX
TimLgrPPjt6bIUtul0tkjrrLc/7fXqhyyVY09SRer09gFs6cmnwNwn2MtseC5zwM
Xx//+/GXhhj15yfViWINTf6JS944CCiJS70tBmrZ6zBsp6CJUE3/n8GKDKXZJt0j
1m0XBKjgMTh6dcnFQVCJQjhW4zzeQrG0qSnnTVsMIcCyqjyRHvpdg90nxNT+06BM
+3DFNANvmdfQvlbvTVc2gf04AqHpBrGgcftCLYaS3X5fha7u/FHUQWmfXoVn1MUz
+7IlwWGkjCflvwb3qtbCsXxlDqHTefisodZE10lyXzKT3DirdXw9E4O6y9/oJjfQ
ASwlU5+0LRrZioPC/Uawwxkfu+d4bri0E6T75d5R/YjdyKwwgZTbaFgBzaYTulUj
jNHOeUMDJf/8AHJYtdBS1cUR3SDCFoY5GgcWXbRP2OjZG19Vq5qKDWQO//zim1Cr
5xDHqdLWK+JQNUpTAXrWLDExDKhIcQVrU5jtBmBKMBdygyjoUEsBg3yaleLXtL2I
CfZnfMBK/+LSWRP0abNi439lHCFOjZYWx60wYTMeIjlwAOXYRbG/lICHHP9gCb2q
L4hRRwHcehJKlX4OzIBQDppo4rS0+sEr9qGuOxgtXGdMelLusX8P+13QBMuu0tt+
FAVEBUs4aF/5SfcKMBtIXTUn3voVGjfTrRTJkVFE+RrFCBQ0R9oSvCSILMePvfdv
78isT5Ubt6CLTh89p4VdGznVqg+rYxUILy8eCc0bc2VcKcucBzOwNdC5hPlRcRUe
5xqfa7fq40W/RtJbZ5Xeo2/qVacJNTaJxpKICd/36KIEIx4mnDepOAlDL+GfyIQe
TK1yvRB19uZ6o7wpe0Xm8l8mnJjxCiTZUsJS6URWBaGu9jKzyPk1R6fvhyVDbKqJ
WyHM5Ayf/ymLrKui5g0s1mLvnno2wKWt3nXFQRQAduT9Sv8v3aFmzQYjQYQwBpNX
35SSOPiLw66w2ubWuY+KDaggPcHUlJOcI+VsbYHPMNq62Zf1xuQ/UgbS8DejJY8f
i9aXpo4SmUQaH20VnU53/qgmsZsWlv9mzgGx/lgp7GRj3ldZ+S6D1h9efHFGDe47
r9n9t5St79LLdcJEkgkScZoxxfHz9lceDqjHu1YqlcFhHMlhfKGOTh5fDVZuNX5R
1A6P8rt6+F4BHcY3BqQvEIsl+CiDEw53D6cEmEgSggw6gR7HgL8dwmyznVBFPTY4
5UfYs6bvr7hUbSmXsa6DjlO2wW+LuB8ZGucjKRdNMsNApRe22xt9gOZq1TKe7hgM
FxneVAed7ZxRZFCcqrV/fE4F/BXQ+P69QpfI6e64bDMJgWpz5+G+bD6kizAs5xDc
DnNAQWml7biy9wu4c0RMqu9SMx7JLDMtGmxhJgQfE+x0+KdZacQHxaVC9Jtpc3gE
d58UAwMaS98fagPMitEJb5M3+4Z9afzUzRocWp8ool/rvLpR9Tdfjve3GNC2FMFF
XLqUsyxr/XaqoWpx1x385efxjQ9NjkXhF3gTeyuE/GNvNcvwki+4ppEiKWrdSofP
D6D/NjWxocXsM9MgGNRvJ7T1UPyN6D7tEBqE3HuSsxUxTL38QiktZyqZCCRZ4pkk
x7099x6e9I/fdAABhdqgRoePxqwjUhNXpHeX4qXuprVTt8hzHva0T1FW43xQ2gGo
j8Z0XVPFm1tbfPbtbLfU6LsM2iYwk46tQdFYjw35SU7nTar7vmtYbBhMbw2zX/K8
GnJa7YRknGZEQIxmzLGsDWasz+ui4/4Q25XfARDKGEqXfEsf71thswARWhGpfech
fuMuCbJ/nPzseVXx61Fh2MQ2l950VoPL0Kgw/Ub+d83leVkRWmQnpHzO4WDgMuoB
FMnYNL/8p76ATizAR0dow6obRwo3zhnrgfzciBRbjQ90DJQmFuV8IgxUXSFBRLkP
CgEZ9y7sqClnALN8/RGfJNQvfsfVdUu41O5O+nk+jpri4tjvDARJYQU//4uH9/lv
m1+1TnmMM+NQQqv0kwmkSjXV+KjFs6OvQwJSvtJ+KjtBYhV6jjTo1MMpIs2dJSdg
DnDS21hiN3gzrUTSsPt6MU/gw1Q2kRj6bJX21qGdUn+ojudbIAhPIWJZ1g1fNNn8
bqhJ31TTMbiuIQ6FSTYAGMRs1GVZzTTIoVgDeDJTjjNA5be/fsJdhMlxF0Zyp1gX
oRUdamheNg4r8mDXNM8VuVNlwvsB12+NioLBpzauiWUAhXNK72LhmiYToVOpKWBG
XZypv0G3VXzj7yd4XUZAoP6FZYnON2BBq4v3B0B8P2odJAqaqQgIr7V2AY1M/84u
2rYoSe5z92sNoSQj3Y23t0w7BP7F7P4d7kfClRsvuUJ/LOSg34twK2ydpmKEEviB
zYAl//TZUF+c3XKC/fH36VG4q88f/UAgF+ZjgMFCGNeVoaGVi4TnN48OXePNGjtA
ZxN9S6a07SBRaD29W0MiKsoabFwUHvSA5MRZtS5tf7tGBuRZ9hwTjAX4G9UxU1WR
SMhhJu+34yiMnYLBJQYdtT8m/yj7wTMV5EJkTEu76OoHNdG0V/ivd35r2XjRDJvm
38RFlLh+SYBqPDHn6qnhCqLUWDKJOyuryneByKBGmqvYCeyzzARuFBODlViIOG8M
/vr7WMBHqVqFB9TMxAAVih3RO2vVgQ5oCfvUjYMghEkowycFcLmX5vUbGwox3pio
7YBtcB6eoyPElxOvWI/ioJ/rMD8aNGTjkT2cn5bh17sb0fvrk2BtF8Dy/L7hRV00
PHmutady3mV0cAgl2nKYPHbpePiyuMxq/6itI8O7DvWpsDtyqb4DIqy7fJq8zTDM
2OKsmhBoEyFHQjLOZVXQO8whluGrFtYVdlXzISIoxwcFbLopvmwEprM1ZvF/F5cL
Kf1SujUEcdfvBFJQxTlrNlW/8D+7BYduRL6ytTouOs2yZVriQ2HcabsWpAVwANrC
RfIQRkXgbFhVt9ctzLT2L+Zh2h3ZyREQYMC/1OQVVEswZXqkcM14TZ1gRdt/ZtEA
/cD1vcOzY+JPwdkP3gxDcGPl5Wv5QNhWOvadg2gP8jTuKlh0VjzsrZlTChqLvt9K
mFO177ibpuxVxO7qYeyWog6uvLmiS9Xjn1HAk3eBmBQHBNvtlUOMdRsVl0f7MeXu
spGnLwbWQWqHwQeoQ1gI+jhGxrl+Goxhl9blrvqQoN1DahlOn0QaJQzYCM3DLaw6
4znpWVLdSwMbnAWMch7Vu7uA67am98b+NlvivbRGaQuDr2ns4YcDcaSbmutyZ6mX
KIjyBcxRdRDIZOt6GjhnSkD6fGVH5iAbPvbnyQ7yeGNhjVwEImasX4b4GIrGe7qG
ptgf+029EjcXRWrgDTasdig0DsZDINnZvBCARdBUGm/TEKht0ajYPsxNfbHRrbcE
XO8el92OoEje/3XLhIM2e9yk3L6/GV/OwmS+z7wLFgycEl9KwHQU3/5oozr8nCX1
4P0dqc4787PGd9R22kelZa/OzWM/Mti0LCh42a+uG5Xr6QVGw/k98YaZWYx6bDiK
DNH7bJl5DBnsM4od1UjLbakQm1IkPWnaMZ0jBZR6gzu4j9mdEzdoZAPQKhloxb5x
LroB810YwoqIQ8inusYjiNCskg+7upBQ/btYLA2SBVb9LNGZsFSOq/nzaa1TTDzG
3mIYKpBVX3LpY+dPelJNpkkLj5QowHr28suohwI++wumQgqfhrOqHk88HtjQpT/t
U66NQNZkoN0F1USuPJI0AvygStDwPOLAwnOiOYKjw7JyTI5n5BNxtUEOB6S7VhoM
GYY/YdbEIMYL4xwUve4s2doIU6/yDSneRpKqtA21ND3lNDsZF24np1Of+vCm1Zc/
1cKS9VU8lXCRbwfc8q5HNtq7DW7mZbkUakreyHJn1MFXwN11y3v0FnSQtwBme5c+
72XltcPCPGSv13h/JF/FsaGYh6NY1HQGEqNOwzTnbVHV4CjnBN2sGrSDbVS3PS/F
LgmXDBO6MB2+E3P4BzKUrEIauBpcjsdYTvDsQfUfiUR88MogUG50IZovQpPUdcg4
LK2sRt3rzcfBUCT4gMaHy+or+vrO1olGFIPzxK/N6PKuV3K6Nzycnn7LFeCsqHzD
35JL0lEhI+ftaOnNmXUNtF1mgs9y8mYFQgTXowDPcFwkrgV6Q4V+INKLN+OdMtQv
gYeFXCis0t43lrJWiEs1CZVtSyiwWUNIz+Ol+QX9k1QuUdAfVv2jtBFyxu8dAcsN
09kAIGgtKs0gWoJAh46ioH/tDX54dRM+PYX8QrVDNXqnPn87ZeqvBpF6/EDLT1CM
zK+SLviN+BduM/i166FqvBoetOM8N/7zM/gTtT/1Ze/d67QYJ+pcJvafLl1nlaCa
2ikmsY4hRJ8MWF3TtGdXjHedhlUzn6wnYo+UtSGVq3aKnWjzJiqSmiiJN7/DNk60
ZrnqRxennqwkXeObGyphMqUhaQyyhLhYc60BuX7QqUp7Z+CLIbLrnE/l5yl+r48A
6fhfniMRbg/7OVWfdlrTtOEwIRqkChW9vnmFF/JxDXSWEqFlP0u4DgpJDEVv+MQv
QdZsw8D9PUK+3KFL/eakaAhPmcSEceTtAfWskMTKhbUZScnH9p7yGU+FAuPWNSRz
sKkZSY8unlvBcYz521WX59l18AknxT4sCS2qd7QrRoPPKiBIy+WMpjNzr12tpAt8
Of6Pxyd+F/unRmF7P3u7EN41Aiizyvxq8aIQmPaagqs+VJzM/afkKSFCd6fwBoA4
B8d2SIIFHzViGEgHfsTpEbGIgIa6IBqDQfx39m7Ygq4xAA50Hr+OQcOBeqLkdkL0
JADUWvM34tA3jQZpM6RHtUoOzmLw2FjvhPYHj+ogOpt74Pmj0DfSDYF1DsqPngK2
wSHVj8oX843aYbqrVfRYT9KDKy2ngflNdTudjjMEVxenDPhdEoZH5eEPcs+0yRLx
8XGzXb711Wkos2ZBtStsymYw4ufdqYTBDyUdNOj+mnppIvrr6pS7OEwGJ6e2o4BU
qX4I2Ms3als9/e4pYiYHLptkRn/NXnB1ixh+Wl50/V+2H72yCn+o2lgIoUrZYXj1
tamRpyHayzjvnKGaad1nBIs5BxVF47cBuw1XhMiIfqBUWtdbk2o0GIwYKKmSwVgq
iOu7i9B70iEU40p5hNexApObnxS9jqB0se57D809EMvvua1e5sWQdpm48IeRAxb6
2RUlY1vbsqzCIAme54Cwi2IZZocJxlpaigSu9hK8osKJ5nreLK6v/FXr+Qu9E5l1
982J/DkEeXOHpEM0CoBu/H5r6MwS8XM+XLzXNu3R4L/m4Jc36WgdJrLFlO1Exk01
+XH+iUqrkF/S1xd2HppRiWCCJ0oxu//3Zaj4WH9YPLZe0dshgeK6tomM1AvKDzMl
GSdk2JoZCL22yrSZfkjnQWsEVUDwl6Tk0WcDIrwO65WB88VFsEJtcmgccPOj6hFu
4DXzF6cCPf1WqNAXNi3TBTnEpfVbms/K7g0VOq1Vsk8mLpHn+FJza8wCIr2nsAAv
nciJc1kM5g8cZNTIZNE9FrKYEJJe5k+xhia0v97JS94xHWHrVRZlEkWRxdVApM60
9DNYG0VGwqVM83dptPXiKrv98piaZTByHZ16VOlAC0hflzX+0joMCunDTD3NA8VP
P2fR8CNRkBuScgTyueJCcebCvqCjRzwqqLh05SDjmVI0+Zlw7fUA0UbL8S/smz++
nyos5vEwdhnTPc/OV6I8q5ooJHOhQgkzI2wvFBPB+l8OLNmgCKhkPn1VcA2Oss5f
tz1piLpqexfMwCEesjjaFrg3uMK7/AL8D5kyPuY+jb1ZFPC+HefE5OAPKh6vpwKP
KM8jBEQiRcHFSBA4aqQ1rleo+oQo/WPH0IwS1IFOaoAqz/D3WdArZYq/mxTNTBn6
oQZnDzKR9dyuzv+2LfMerWyUrYGgIXrgv6OdgnC9fvGnz7E+x65P7451HaB+Ecju
mTVdrFh8CcIzyOauUoD2JUfqv6M6t6/JJnhezdMZNo0h/TCqjena+Q/chD7IP91Q
ScNv/KlRGFcImiKdMo3e2LigruAsVbW+eYpd8sImXnPODBGQ43h3TolRlpFQMITI
/yw4AokzkOirMF4vUjOHq1G9neSjYEuvW5q2rdci/xij0Qu8nyX485yNqXCQg4ym
VdX2+BhSMolQeQUyZuXIUzAAj3Gk5mNHDILSuXA8VqJD37Knn9Jf5QZmYUSRjDvh
HEQ076ixJ47G4Ecm1OyGXcQBtdZz31crxvttisy5tJ9dyw3xvw6bzAPg3zozmUy8
/uybuVmq5e6n5omRh+cKO1sGFzQH697wnmmwhlgWSd7Z95dDaNlhzKuzk+c9c8wd
LyOmu91FrGXF637saeFoIGkV+et8ZUxuvVGYnteWjwoqXli8SFexdVw8yxcowkRh
XkSl4h05fNbB4KL/Dd6cSF/E/98nIaMCMBzgMTklep26XnxC2jj8f2s6rZsSxOG8
OA9TMzN5q0o7IL06z0h8u0Mv9KIYo/yLUy9GrwgK7NqBcgY9n4O/0iw2A2YuCt84
uGeqtVSmuFcHcawXFjcfwagPzZSzhZ3UdTAXWEPA0rZ1n3hBspeKLfLks9m8HLRV
zPU8SXjnoTQjm4qHASFYMVXPBSfwpI2Pjp2jB4wAe6hQE2pA8PhEbEjA4GiCUt+R
9Bg1+mjYrZrNhSccP3bl2cDCHmtkzXbgK8+SnjZXvQaderFHgw+DJygnS0Weo6x6
kZ80z30GS+vFcknOTNBN8EPpjEEAW9p83Tl6d1hYDVX9tPMv8eXVctPqs97SMsKh
cun+qQqKExq/BJwqysY0h40sQOAxWPBqLG5U1Jqu55OrCQvJd/5aUtgM7E8e4Iv8
dpjeyPO+Z7gDFmnTsUCV+dXpWdMwIJYYVeByy1Jb6oWyoFY/+tMYWuRkhCB1PhL/
ODp1RnTikJFIugLeBNxU+WZ6XxBJt6KAKTqO7X+uRNVZLQKUtlPu6Tqg00ge6I+K
KiwA4gdYryD//y1aAjKElENjpoL5lQ3j3eglSBCjiFDH1uxX5+/5aHtvny/8dLZs
znpNTzZg7ENkujlrA/PdTZF4b5QfRiC39TDpZcpQAEQR5v/HphUPs+gLtiHOkH/l
wLyzDvQEQhdYNm7Ti2rVFP7C8cjftNA4Ks8S4A67KW7Ea2b9qCXPY/2K/41NLZre
3MwbnTJR58+AZpwLoUWoF4bEDhVEwZ468UlrmNpAmHWM0BJjOfZcyD40RtF6t9gR
HGHu/56zeqgpgoxE8b1AAvpRaGALMgcfNvg7qwKHLBygKWyHIVOjePOqNgJQlkZt
NAJ4JvbRBqYjLUlB2Ccvl6lap51y4ZnZOZz/JyyVymu05pvtH2fxBTlUDN4xHaxf
IgJ3LNTH+K+LYw3Y3xTYGvQl7tNkCbNLG7DkMqOmBvqIz3VrOafIiD7kifd72tAf
SmGPSVGo/Hv8402qLUy18W010+cvpLPFCspfvMP1SXyJecCzoPtBhIM4JYiQcWIS
SkEM2ZKvXl0SR8QmPfUqW1FFQTQgrFXW+L01GiMTRRhd3GvpW9hiRIbBMjPymp3r
DSMvZmgcYDnds4cbWDonY22vJwL//Un7RwOLBT3myfk9qg5iFKlQd+tFir4Ls3/7
FjMTi4VzLQMNbdJn4NVQ4Dd/DlLsDWApnbbxWDPc+fQTPLpPLGM8AjBMAXbkzvAb
HEsFe4b8w5gs+Qzf4OVBpIx9XImdRZmRPbHozIVKffvv4vZR0HUnUtVaRolXc5Lf
xtopo11I3LRH/+X9m3C9lxZ4kamuqQCqBDJbI+6lz+UB7iJcTVcc83ccmG+xv+vG
W9IroNCGnswcwz+ueaYjRPFf7feUzo8Oe+0jAbw6W0018NTRcjPgTEjpF+drHO5m
jf3+QLrPE/iwUKM58PopdU+URcACKO+KWA9DcK9U9CvYOtc96/yYBIh4N/qexNeQ
Mqc2jvfi8p9v30ojmObPPHPa7kKCPt3src/wzwDVusqNG9QRT8cQBuJ1gn3p9+oR
XUlXPQpIybuJxiZ+qdbbM1lcSJejiD5kWJRKI899q9+p8V+DSuQO8Sv7PwvtjFBT
kjYAeQNTO8mgThGUkPCapicZHfkr8fyd75PZ1Y/VhXFBd5rxJyjcrNgl6Z/vow2Q
IZN05qrdrg4GlazKHajJBnAmKWdYeTgJ24icPPASorDlJIjN6+7OO6ZDCR/dTZ0y
bpVP/M2gKr3pLEV9woH/wI3+l8KV1dLiJJrPDENpTCNWt8golL4D9JEMafHmGLwO
Nh8HHQ1EJdOBRtUab/xKYYy5SFIiEvllRE+jvlTrtkgNdTouJvV9+Dt+OK+SwBqF
3voJKiEmz17qsBWhh0REOD4AFgB7OPRvgR18yGdc3YnPSFTVnsNELznz6Xhg8rw6
Am4Bt55aIvW2f81wWPOxxR8DoiVAvKaaKfGDDxxXwZGzrSElkMZoEc2RI5dLuCIh
xyJBghfDInrZQKVrWa1QSQyetnZCFamp1Mvll79Xk5OppDJ5E8qkovK6B2b2o9+M
cdhpc47RnovxedY5243u77ABQzOa6Id5DLA6cLxclceQKUY72koZW1ErG1w8gzNN
b0H5T4nnmSAp8zcnfxwv6ZOJjC5ZOdZPAGwkxwt/sP80VU8EWGhBeHVxdn7DMWCs
jpkXiMqyc8QR4xnZGHQkOeYwv8QTLhaLyjx8jkTqlKdm6Rp320u4QgEzJh5qMBJx
YlAgMZ0ueOHP0N6AhJQHxnqK9XumaPH7cJpwRUsMMIQJGmNHL3SvzB9CYNgG31wt
TZXPu+5Uby4BoVjogDaEckEoiiCnCaT5J/FWnMv7egoKkTlz1hP68vVMa34wZ3tM
MI0KlAm1oaAar+uRW12LNxryuv9lnJuwPs/mQm6y+J6w/tLvd0AYymaiQQZKeLLg
7bLi4Y5j1lKKFXWEHnTYt434niLv81L6GIVHuZ9h/BSf6MFfkEnC6orhK5FVroHa
GAoESkQ79BLmJatG99SczfoL3NI4uAuS++UjNL87q6HTsRILRRxPkjWBq/tYTG6i
0bdeOFrjbrH6gI/1nhZazO92+vNdzP6OomJOK51Nwsd9u8IihM3mI2TT9VYZgUZt
IQ7tg4SNV4nu6ri4p10/3dld+M1NmlbTUU2j4e5Ag5GMDjmNGFYvAPNBVxpexw4O
XIOwpg4BCsVwt9B6zmZY2BT66jqTdGWDU0H3zVxpJdGgUzes6Y0PYlJ70MnTkOyx
xa3KXr2u+bfSz73fIN0odxEpABYFnFmIl/2d7TL7vGH8qE0hjJjkJ+bWK68voxDC
LSeT/1Tw6u7RSBf/T5+kZOXc1jzCx+3BdCfKxm4pXMboIw2vqREoKEMVsp8sOZMY
TJjFr3iOGz/dHvJEhG+D1YmWPX/ZZLaoxhCU5j9zpNB8HBX7fezMRqm49zEM3Ay4
Lslow+2Bg0keaOcgAwGN+XJ3955JTJUliEoqqiFQNly5iVfHV9G7mJwqKYew+hKS
RWO8WaCWVNm4orl9QiDqcJhVta2aok/Lswb54oAs502GBhMkwW6iKKDqmQ9s/+nt
xQjixdIHcvPOn9ycEMyD0t02q1/unyhpNzBsDo8XrnhIQRlBh5GddmNiLu+IGRbN
mAxm9G4XlAirXC76yxjiSAt8XRrG7G0SvFe9LgyWsSPw6BP/sBUjynD2nbvHzo2y
6OSPWT7o+ofD1c9Hh2b9oiEeRVmDoSQVUzxwPwlcXrNcsGJn2u6j8d/QiZguvPKZ
PiN9b81v8lAkUHh4l7uiK3T+LMJdxpOy6XsW7YoG19zDQM4Htb+Eq8w06+R5EwEx
rMHyQrOfvE3w2SqPNHHoKYL5s0U8cRjZBxPgIDk9i8ymNZ4Ao5XOk2ixhtUP8NNf
6r8Nu1oqO2DBeXymZIp/Cvlb4bKGdX4rWgU3sYFCu0S8pNiKH6+VOBRuB3Oy3Nt0
rPg32j4vjAeYJJ6VlqF8esQFFuvtqmETXzeYiYEYAwBDjwx3QqXagLfTlMVszQp+
d6fwuRx3sHiHa5zOG+1Ge8xBRAgOZlEMcyMldL05ILBJLLQBCb0DcoaCLhcd9tkK
sxRgXs4gJjY3gFd9sRjtigFxZy6Wpy3g4bXnafuaoCo1aAEXmH5WlGpWFRyFLCcu
34+YzMzxZWtApCMzWa/Xxm9xIxkvGFKo5h2ct4wiQ+2j/NCNtayKCqji2WgqynYr
ftXaB3NBpkC6lqqYXA4ZWocUbW7qPkoPwOfFrR0f8C3Vxmi/J+KdW+r5EA01dzA0
WJwvpfdpjxn0sSTulF4AY/07z1soeGjSQ9IdYeIJPu2rB4jIcp7UBKOM+4rISeBf
tKMOGtEnUaqn1y55EaZAVHuvXsjBDD+fHltUQy4Utxq9f7dI5f+2xFHcXL7nVJBq
mWR91ipGm3CUW1iLtfff45sqp8ZK5+qHXQaCJ4M/hi2W/GZYqgQCp2+om2ApciIj
rIP/GkgoBEXZfRhTRfDYKPy+HrYmf6OTulnF0+0HvToWdJhbKib2/n0M/47qprm9
7eKF3UF3mXAPLWrjcdIpN3ImcvpvwPn4JDO9PEr4WWlEgVK5yG0vvEjztijCCKIP
sqO+R2s14nrev01EbGqjmC0rf3V7kAP9jgc6dKYAB28My4aHG9FdHCTNCITHv/Ce
yJwEnGwPvicZAffG4YzLuYfhXTpukvD9aRJk81u3bHlgRITcSS4VspdVSqQpZf0x
N8BszFJGtO3cd51LodcQ9C+sa8hXGbEHLzx18zDX7qvlzzz+G0CaaoiKpePFg69H
jKuikKV07b9WxdkcdLhevP56OizSWh7CmZFyiYKFXpkf4WbAFcopJHEwSs5vn30Z
Lya1v3N3Ygfbm9ac7fkdjPccnDqVUsEzI7cgKfFS9adaWvexaOiIskV1brmHtZOx
ZzNX4QyGUTkAzS+AaDwIfQB7V1oDsqiPeUExJSHUofVIslwf+u7MD43rkK73CM2Q
gghvR148uL5ThrmW+0vTPq06lKRGC8zzLgVmHwHnhhWZRlAk+U1vNCOSJu7mzbz7
ZWlzigA6BAyRoPIVmLIz65eWZyLKKc8Vm07TL5D9IsBVrVEkq2f0A3psfqElUiPA
yXq0GPxPowoKxEYOYzsVl5qO5+iGDGpf8ng/mf/2/SW/EizzIDQEoibbW7VGYxas
4id/QESvf8kcgcpmsz3rdY6Vs6/OMrGj8JcPWfEemVhgLp3V/MWwLYTOUXWRrlYg
MV+oZXmgVbkUfzJvnIqPwAiHNN+s3ocWqfytgcXmk0ruzY6wjE0mV1HLmj3iImxI
be7aMhFBUgP5bPPejNul3U5Erbd/GBzkUzrk3lZmrma8NtdhBOpnr2Jw7VM/Y/IB
wCbF/rBvnrTlIhYcWwYhVYL2uvxPb6SX2MWJ4ESN2ovAKlNEjw6WPDOP6YO77fWc
kEDB31qUyeZMLC4w8sur9KLtsgnWUawXSIx1Vaw4Pgw2Q41AnUPUOGZJCC0etEGK
Rag1NO2h+nzDMPgGqnQsE2CbYw+4JYv64bOfQg73K0KYh5Ii1ZzwCmzSqBnbYDgG
wTspQQ0UvsWBawzcud+V7Y4GkmueO384cW+X68BN8wKoglfvVAdgBY1wj8PIPvmb
0GptVwfhqdg+3XHkeiaQAccCOLfhVkhoMPWysywmS6ty5h0HUuClM4aI4urwtG6A
yL4CCM9lEUfbe1htPE4H1gi6IPqtiJ7Vc3+5SZPS4nmpNwvB6f7cJc3RNCVpylfY
kYMf0dDiAtBI1YqOjV2m4RzHXzLeg4n14vfNjbG4N5yuwt3LZQgGBwliG8WDOoMT
74RKkbK5GP0ZBShxxDJAsPnxy7Lbe9HXk/OnJUVEloH2vBumXNH1sqYUYbzr81JI
nNQpdgsuKwl7nGw9GpcVcK6JLP0tsH+QkkD2Ci0KOCaq08qsX6Gvnk5NQVu8rCzH
gZmf8QGxpMlL4HXRe1F518XiGv0INe5LlHGSAlVGztBlYAhsxA8j+fsUqjMyOrFy
bRDNgn7ZvfnBuJlgtL4spvK/ETESqrvHric+C9B0MRFJbtCb5MkxXX2HaDGrHEoO
6aNGYeDMeEDwIsQHa1zpfw++EZue8I+gM4MiaEpR4e29+2Kz8c6fSOOJNYYNVZBo
hyQJlpfH65k4gIDcfVW3iCi2CNS6pajccYXWo6/iFOqfFobjDMoimtHme0sphbQQ
mtbuGY3S5MI9i4zsnUxA4BPeVnOFgpwx7IueYZYcT4CYIYMKuXZgQu8+und5cnhj
H0DZ9gyMbOZ8aO8tPjNraVAVRSSL28a2cQbfdYp/eWrk0qGEhKwrqphEDwYVl6uS
XW0EIsaVylpu5kg1lyf/Gjg+mE1JHxy77vqRlyDvGY8=
`protect END_PROTECTED
