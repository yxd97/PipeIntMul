`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GqzYlTFx5MHliPrURv6ADJ2hFBRQRpdvYHbsOejHhxfBwWIiCy3isLE2anrthNHT
qy2wPEgDMq4Yau/H+JlynrV7oPxt+0/sJbauiBgZ24bNOyd6OxEOxQskvVXIORaM
vIsOFO8GkibJAfHV4PC1BAGdhXXK+KNowEbZ5uhQsJKF7B2wxt9XxmcyVPhYyUg6
U6X3fw0r/Ts7QDP26xToNp6Q+wAgDErcTdg2qOaRPafFGb0dRGIuGKwl+hSr6nBQ
w0nic/i/h+cBIbCk0iGtsgL04AR/Adv9lz2JjO/HZKKCiGrZYbuRM7YgQBCDz1dR
xK9nBxSjyTXGk+gtSDMeMxnNqBFv0PP8JyuJtCTH1dVvhgCNv53Itvm8so10BXOR
goz9JKxl8yduTFNp8vzAE7YJuae1YwzHd2li883YBhT2/SGt+0U9FVDghJxGc+OV
qxepdBo6NhitgLjG3n8OQZVsHwHCPR5FK87sGzRIspbNAPz5sK6nqWkVwkU0Gqqx
`protect END_PROTECTED
