`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UQEXc7z3ESUPTk3HaT8/VTNyGwunD3X1Of4/6fa1r/xjivB2BxSii9dTxf07naEE
R4caVXwrVuZA3zQOVmRqaiQckZdPMPX30n7glrQogkPb9/0XNUp7gH6yqqcs+YVk
zr5bu6ie6q9yrx/KSpPM7OOoPxiv4zQpm6K0AzihT98O6O4FvcZIqnS6jc3KguXd
LDzXAeyansbQ+PS6yo3Zxq52NWLzczGaMf9F5lKbM5Yvr09KQ5tH+ZIWxNkFigbq
`protect END_PROTECTED
