`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M7YISwPZ7OKCZtfZ8xpD5mTnk1XzcNUNAl5iPTvM1MR18p3sf/JsuJ9lUrkrqNTM
wEUToIlbqIQrt2oXHdYlDAn0ARumLh+TjnfLgLkFcC3MuAhge7bXL5YTH5m/Bca2
OGCmC7x1jnhEZuVNuqFUF298lC5bqNef0kcA51ANdFpCiO0SPhxyNrvT51WD3EhE
PVxw+wJ1o19EKnQ9p1mNd6/tKMZlBUlM7sJn0O6cUDbAqtVNyYgE4geLJ7lWjtmu
SWyuajTS2ZtD40rx1JXor3q7bbO13NHBakkyZW67MEqe43VJ0HZaCKxhZflG/vka
69fNdJBJ0VPwziAB/v2q+bDa6BPnfaOcI+KfOfFp0l9DPjNhNCYuhk2om2jrdPbg
OheUorX4tVnjgs9/OsF9MDsvg6ogkQrihooGaYq6UL5UGL7V41hCAyWpg1uzdp4t
+vrGRF3fIiS8KI5oPxqlJUjcFG3PEX+N6YlnZy0ltqNu00BD7GHizm/HF6BPJqUB
AoaXZTE199PYF1PMn27k/EjCrAMn+y9MxGcgE/RhWHchWkmB2xfTkqq0+zW0OGBl
7SL8afs4VoIWjLl6vUyCpv21pZ4MH9ATxtkeJgsSfraBCoOl8ISYOg6ySL5TGVCq
obkrctUpbPAD1aqUzMve8yc2Vau6SclKkLxKZSOORjFLxoJdhy22PfzOWFfdf1ru
axetb9O2gUKswJfXLlQzZXYrjkIxosXr/IcJaXiNe9qa/TSVRpP+SEsw+i0FpS5x
MYKKa0MgiEDQgQ0IT0XDcEqpBoejle/D1tTUh1Lkmhmahmfv8TovCh/YugobkB5H
T4OsGBGC8IiVz3aFJNrEiYtAAe9aqh+IQspA2HDfyRTTdIs0eNm/+BbPWywszFcF
bOQUeJcQDAiec4qbCz1sWdZcpPCsPppj4kkx1+3nIiVAQHYDc7djYtJ3taysaEA2
1/adKvDXaGj/uqn46ePdzczN5+OIPp8ndQpuWRbN8sE9iQD6mRJJ0OENGOOzzU15
eEtsNpmaA84dvBkdBmcvMaNIQZaW0GWNjTmSxmNFW1g=
`protect END_PROTECTED
