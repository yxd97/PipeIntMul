`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6RK6Qcz3pdU9XejX3NE1H4aFL7g51lnZ1mU/TWoTfyMrSQ1gvZtIEato4UPKX1W
jD1eenQo62YtWiMKV8yNu0Ds+H1dL8AyubxBl3nN6poACNCmfTQmLLpVhQ5n5X/W
ZqUWT/S0yewyN5OB481W9855rYmALo702fGNDZbFgVKWilI3VMyFexgi03VYeHkZ
TllCeSGFHxD3BOcVSIEWM5AkQADxCyPZfqL7Ik7zT+TdjpUncXw1VRsfaMSnobzP
LbibIocLg/eWCVjGASCrO9db9Z+CsybyfGKlg6sF1TuWLztN+t2zCxPL0+BdMmDP
`protect END_PROTECTED
