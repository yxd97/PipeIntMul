`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nZKHE1JNXqpcjsqauGXLxty6P9AQtye0ABMzwa4iOKYFxJGtK9nOMLpXk/1kF0Dq
oOSV5Sc6mPnpsLA60jejabcdR6zoXBV1sw7ssMgRdO5sbqy6CatWmGBT8DS8Gj36
Os+XnIByNTpnxbOBpZsquYEXXhxlb0eoJehuq74jcQVh9pgEugwscC8ohhljG912
4PRkz5RKLLpL3IYQkY7RvvyJGP/SzOEbdt3HXgVWTtHMo4m5E3tHpe74oYOP9XpH
UlOzmHEUdVBIHUF76BWwqRASxWDtJFpmFofsaBSx42krEJE2Cf4trMYYD/NRzRSC
Y71RG8HRJzF+HLAZlMDwte5HsMIhXWM7QNp4bR/65e9xtMA2k6Xk2yh9AS4smyUi
`protect END_PROTECTED
