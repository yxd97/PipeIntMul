`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQpJgpf4dlMuM43Z0hfO/FnMubeZMsI5o0XcXlvR8Nh/OPbsJGfzL0JPrGBTlxYu
nY1DnraD57ggBcHK4DE2oQ/q1CtzPNa7PqKSQ99dV4QDa34ls2rHAuM6C2A1x4XR
ccgMFES8ny7VUb9VvBomhzVBwhdgf/8NbT9v23oSm547jkMQ1ybZJtFQhEBDMGcl
KI9X/MQq2TvtbAxWcwgX5VPaxYkPwVrV9N04lto5/H4iQHVFtGooNBPOapsBzfeg
c3JPrJbgs/AfEPSR/Uik9A6iuDgBcDh8PpvOA98/j3P3pw6Bbo7Nadj6n0CVa0eO
aU04P+0v/bsCbJWbC3tx/LVP17r1lENwbwX3E1Uv5kfAyrWXjnIbLUB7lgvHp8I7
+H/FdJSV+ygWrn2KLt3nR8K9388+Gic0e2DB0d86UN9oS/j1iuQ7nNpNkEa5dPq8
`protect END_PROTECTED
