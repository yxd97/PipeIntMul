`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u0kqig3qpsp5MywoQ3NNBwC/kXgykFEF5+mvb6oHpTlSMSwGIaHVn7MnSvIDurI2
VuCkSXXycbLk7fuA+UBXwWbQ4xcFz18llhj9bJF3A1JhLV7AN/kKRXZclIyNkPrg
979ej9tMxVsLBklLIlZxSHNyZgmZ0K7LRhXeXLlJV+OIAGzYggK9P1lAR+BqGDY+
mVTEtpd2IXKmujEkB86kE2p9fSAUBqg8FYkzFoCr8sw9m3fCIPXW9H7aaoDFNmYF
ro3+PXUghD7W1qKpntYd16KxwQPFjRDgO64QLUdzyeovQfPJpJw2B0+XrwZN4BmY
UaKrzGfh/+GFt5IwjBT9r7kUOsV9uCsQMFandr0gXX5oR2l9gXuqDShuKLXvsg9x
828g/KrSva8USVxHuq++jfVmD09P5Jvx77CLw8M2AMG0JYB6hOYkSTwRdyk4yP1I
ENq8cyMDmCEirNCqYsGoYaOtNOEd1V6+y0CaGYlGodRB0iGZpj3Dlj+w/bnSJkce
R+Scqq2BWK6jJcvMekVDOOVRPUtQ/BCVIXSEM6+5olcxlK4FtTsP3HgtmKnM1OTV
`protect END_PROTECTED
