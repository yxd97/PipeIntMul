`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mUzN2lhZXl1kQFudADBpjLQpahmIXZNzKXOLxMyCzRD1wHHhX+DJ05xYZGXHQgOn
dWJrOXXBvW8qnfUPcUutnMhRhtY2/1odNZjqNL+W+1vK61pkpjUk+dV1C0Opfe1P
roWqYg5heRDE8JKZqW7hoXkFb9uW1RcuocUmP2zF25/TtBYwRpLsGwfKIirSHQss
dogPwDDKlVldgTBOOhZbc86McvhfOTdx4jpCmd5bF/NmDFPis0PoibZaMmxpArYW
cm1SxG/zYLHDRqgzcNQgTy/qZeP+oGUU3P2gtrsDyjUeqw4Xj6H5NVE07k7vzK3k
mScZeowJc8vVJ7Q56v2SEf3Tai7sqZJS3HX+F33jjN280ER9dOQd+4PylaIpTZ2V
dNYKwphdFDB8mkEJcOQCyM09HJzrBdMgr3xyFhdb5Ho=
`protect END_PROTECTED
