`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1Ws0+sL5NEgmxSBsSnKtfh6Kw7NqoO41vhGGoIITm0Mza0I6/0zq0KXZl5tI29p
B8RJ8+sseVhcrOh0zaL6VaVwUWUABafC/0JUuYAUYSuNwd6Te5l5XSLdGZFMAoeC
fyXeaOEwN/iFdQZUCAIXupl0mth/tyxtmqhiMEMp31Dyi9bAY7K3ffAHRzvcSJBr
U6G+mpnreMlYOZN/keIxr8145MqA+XRtZ7AurEV6F+b9PWmeibOef75gLebObLMA
IX48xYGhCPo7r8KsQBROXF3kXnUmalsvAx3dhTmjArx5D0CN4fP7lN//7LLnyb63
CszYDgScD9bKJMMpe33G/afhqMfdVrNe1IqSMmJV0xqYvmnqGsat5eGxELvNhNJU
1b4c0Mj6oLjHOVSkb795oV4gpRv8hOOtUp5stksyaSsmDp9JqycsgK4iyUZnXffc
VgyN5BgzfM04mv0mKfDOCiMMweeoEbEXUZywBrBLhXjUFYNNBeVbLEF6IaqTyLZZ
EzcZbQxXl2RVdECn6weU4jnqcBQjwfq/CnwiZezyAT3sfEYGGYZUy968GSMDJjTH
hw0NFATkh+IVBbrZdK2RidLkQEQycdtldlCLo1U5xvRmkl4HK/N7hVadvjrOukM8
7np+0f70AZeBkGoivCDVTx2dg7xxSJoYBj0dw1j1ecc=
`protect END_PROTECTED
