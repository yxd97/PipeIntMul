`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3ObPKrbcI23+Du+htmCmggXYgkYewcPXPo+6o5MLWwPNgaqXrWQwmNNfJjysvzVK
WxW1U7YRG4JyeROIXRGDXYxFh6hWVutZ+WbKE4CsDbSfhLI1AZFhLXpnii2Xp156
mXzLSqakF+ivhVxotiIx22dbGlmX4R4iUBdrkD5dErurlTYx5+tHLChkWfezdi8i
EC3Eq0zqXaMzsqXyUL3gGDHmvOOQLfOa/AkI/JHxiBJfYVLW4XhcS6Fqxav0tZiS
pLaacfb4/mBrediE8UPOUzd/AkP3amChAlXUgYP1wl7mmI/Zp947FyL5bVorXcLz
qBWatHPSuLNg7jqRAHQmA81DalTxiOZx57Dv2/C3WigUJpwcQpjDAR0NruL00p9l
DqBzVNhurEeSrfA5tSfDqdA1cFGDXSpdBUxtmUxL6EOXro8sUTTNd5+apm9d9rxp
qB97xonZD0OCxP/sucEuMblRVD4rUw7vBK6KTQ0iar8N/XoVnAXr8GCSUgokGTkg
HdIYa8qbLMarq31Usgwt9JHHQCTuapuguXBQvw6Nrc/T5LUS/sulv8yUWeVr+VkV
efkIrXHjMxkJEFMN5uFz27peV46SNzqCdL+S/Auj1cr6DBOf4IrswFRh9Px5tMNz
`protect END_PROTECTED
