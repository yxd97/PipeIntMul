`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DlqM4kXGypEqqZ8+Ir3JBoFv2rSFy8WZSmcpfL3Yz2ugtHO+fxkEngLXl6Yl1PEa
/ETQzQg72mxtNYiZpe4YwFxlqzobsUKxV8WvMj8ZGx2gi7K5wPLMSkJ/4BU2nvix
d0PDUTCxlTPn6BNXyFOsh/QCzRB534sHi1O6fkIk8NSyziXgsWvCAymtEyTlGp4q
9LDRn/V5j9y1KFOm2zS8EGLko6RTD44w9h6+Vt++IdgB/z+5LOQ7GkXcGiz0nW5U
W45iqkbpkoWzuygSRk7BN05nzDCeyx123MHjUJv68UkZbgkZTE929j05NvRRsNb4
J7yYuswoAaj00PvcunVrmmhlA3Ryw6B1pnmZu/0WscDYoXLLaFmcMBgJcw1CN1gQ
x0Pi5eDjMXljiBRLOlJKUTgLxdAZ2K3Y0B6IMH8js9ppAlbDNaWbtAbD8rcINRNA
FkdUXnt+/0jmBu5ZJn0/9T9vnFrDd2vuVeSKhJ2yReKKTcjdfPWFl09xZm6etTnd
M6s2nMqYiKbfRHn0YCByKJTLN8U7pCIaIPU4SkAkyPck8RsfE07+rbEGzZsDXv2R
oRmKN6IMNeIovpyrI8Tq0nrznH9mHuZWYFWRVtXEETw7+TzesFvfm1Ev+TxHiebw
ddxVDY/Kfpi2jUuVa0xbuE1d6/StmhZmixtUWnYXK1Y=
`protect END_PROTECTED
