`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lUIuO6Vyb8wu6FeuNRQx/1maaGCjCjuTmxcRfz8mlTiE/45VO20McgkgmO5NglWn
qGWKOt1fApHIM1Xbt8ksaZaTO7qeE/JrUaZXE/d9T86x6fSm9EK8Gpvbftl0EPd2
i/V1Bs0YVGlfj4F4xsghTZ8x17L5orQgcuKtS4uFXKuHKdVqtyY3XepsLv5Mwykk
3xr1NtVZxl9Wy0JrobcIDWNgxwT6VpndlITXO2opSmJY78f7O61gHBhslpwGYc/T
bpUSCD0CAWH6a7give2aluuxLYTXKaGuAn9knE0wfEKkdo94YrsBz0CGOt8SY1wn
R4jDWxg7yCPpIkke2OVyUG8XMlBHjEfiA0iwbUvKtLtuVN/WY5yeytEjn5Z3yCCE
HRteT38TUep7xn20kgSjccpESAmKUL6QuU1+aI6RNhkPU0GBQNZGrNHzrBCvvTB1
aBPHgOHMi1uDQxNrFm0ZC0ALyFFlOIQimQAyfhyq4WmefE7b29eCQurlfCF+2gto
ZEeDi9B7SRiQt10KqeNuYUI5oMxDf20G+ARXOaQ/yeYmmLcMUKzuWoUKrsH1h6My
N5NpqpHCSNhVMiCPEfP12OvhIOkpuZ8bnGYNIvGV82jHtw6yPVjdoUfaFfohni0C
srepZe0kXMfO9BObFf+ucs8Skn5O8hdt8OVZvBEr/Y0ducYPjXZ4kP3JJpjjaJEe
GM7WG9woALEAne5SoUHqxC2nWiDVTZbiX/xtG6kdlQismDswbAOxYSOxRua0hE7Q
4WgBauaQpi3Q4hyQ8rEESVNfYuTuNFJmYw4n0OvAOJ82k80c3sttKlrnYy9djxVR
ohmMn/6BI635jCsRHSgOzbZPPkUcCjiSJQqiHYqTTOVbchcafrQMUrJnOwEpjfKS
NHd80bCaNnO0BhTWy2wOcBJ72n+kIbehjEYQl6Th12dBSkhqAA0NTMH+dThZhC1d
CEqk4wOcgVVHUeU0uu9bnouhwaoOK3ZrC65IJgZA8BBdt5Mhmz6D1x2FcMmf26bE
4iQZRbU5IcBBdFfd/MNxNZBwUtL2qmCM7LrxDkj0VR3ppum783cu+Af/H8Y4QuEI
FSHwKqplcXMMIXaIduTP1de+1yPFQ0wyPhyKCw2v/Gl+oe+dnjBaPS4et1P3xd+0
RXEVYYB4Dqt7eV+QVk7ULeXyMilI+6kNM40p/l8DbItUAl2P506mbKL9RIyzGHxj
QGH2p0/IGF84JoemrW5CCg==
`protect END_PROTECTED
