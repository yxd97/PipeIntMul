`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bxXY9TSL4AkP/75WmdyWRsm3TxDzSWrTAnwWYZy/2LLevFJ2wNSn+G6BjrVJ6oHg
4auTfMFLICGgj3P8FKz+eLndMdcQhqVN5HdFGdkVZIHwojnPFpjlUXTs/5y+uOmF
Ixeh+Afo1OuZ+ODxpOnzIp7PHry+A0finrzEhPn/JIuchquAStuBsgBhhW6uEWqo
7k26d9Drph4oTPtCr9WOyQaLlj8j8Az4T80wVE7xDzMMGJRkwgKBer+Zso4K11bm
5AUujfAAIeiwqFatath+NUMf8dzZmC3fk8wzDUF19JjvKfo65sRsK0GWNSL+aYAG
VE64fpa6PRkaN7hlakW+EDKbM0AqMLfgNbcxz0A0yhf7DMJIj5c0gWS0IVsVDkxC
0C3daR+ymgTf0k1L/h0BMhomjLn87lCHUVvWOsWhocxDRorpy6YkPSMq0AsKvblI
utrTGL8QVjmdE3JLOf7Gig==
`protect END_PROTECTED
