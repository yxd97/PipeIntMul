`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mPOqjgL0Bj250mZhffjAnmTWYBKV0KVqjSSNPVluspeaXhWQM6grVCFIWjfxe9ZN
GjTzmnHBEn4UoyqE8ofctVTHo9aN+0v1nlAmwl+CGDVoIVwTvHWifAx6+Ak11bQG
hkzYtz2zfM4AIIr/bDUuxkagqZEAVCIUtLa0OHwoS90uZ9I2tjpA9zlhnEhvSmGM
LwqEGPUMMGrds6MgZubufjq3T3DDv9iRDbslO1klJhF5tTvYebtZvUo5nfLA4GuY
Tvk//kGPNacMjriIBLntshTWwPqn8dEEiv01dF7hMyNVCSLiC6aI7mRW8pQSU3FG
MLg7IROLIcnd33X75nNGzw==
`protect END_PROTECTED
