`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdXd6dC7GWJJ/rtyazswPFtwNBFu/UB4dzdU2RFksDDnCrwi9hB4G57yAWq7naDL
MReoU+hg+/7/9ZF8/0V4ZtTumUW4Cq4xD8DiIPKbmYowbe85Kf3d+fEW56n1xKLS
pw7muM5vLPxFQ0vpR4bItcua2LevczG3tL4DNVmpHh5YMbjPJcTzqIlNr1h+Ja8b
rmOUYaNe9at/LW1gfEmqrdEMkRl1H89ashmAbvVgV3uVBsXw5iA84gzaL65QEG4i
CYQMuS2OutxECOaX+bvn5IRpsqnZzcNKht+ZLvki3SvFkwTgSA7CoIdn1t37OI3s
QsxbVHxG8TC0/y8Duo9T9FnwUeKjHHgBFf0eR0Qu7PhqpRii7S7nB6UMjcG/YwtB
F0qnHTBCmWrNFopq0e3Gs4d39Pc/adXCXlrUzo1Vg/DMWK6pKjXtr7JQPn4NXlYF
JaVPSPN4jVfw4yREEWEF2Q==
`protect END_PROTECTED
