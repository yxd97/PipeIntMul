`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7HjtCBWljYRKsx9wxt5w2AkOd9yyvDvqpr5tF7lgA48oJf1McQHMXX2NnayAoJvy
TaCl13oQNKkOt3BcfLtdFyRJhy8GfmWkpjBFKVVpnbBBwZ3LyOr1ItuFDdTjtr+B
Of6yxKgupNksTzVmc53y3SBo814Ibsd3rh7NbNB1Y4gawy0wdK/qiN7cNbQJDGDm
+sXCJHyUyXOWUgAZ/lStLRvC+zpIXmDhGQSItF2DS7R0tnXJZ1yF+RMlFaouaT5L
z/VgBFblTPRRwY1JGNAnmrtUvwI/hUj6UjkXf4dPzdhRpmyNPJqGJqtx2qJXEED+
5VyBW3AsLMsO0LJ1PGPK5VEXn9feAVUVs8iuslqaRV6cFLSXUqYe56ZBIqY4qEDD
GNAdUCi8PXtzPHK2bVBWE324zD6Cz6VBFbjpmQ5b+PdPPszIKYdmrT5B/dbgz05W
EyanXJF5ZxPFknh2UJhK5o8LRt84C+IcnH3jS7I7LKCu/9A2V3R3Tl5FuD2ghgDA
ncfyU+4Jey7YQyOX0uXUSG1jpG+BbIlDtvlZLFc+F9MojsD6rEPTHk0vb7o2rnWt
pedKrq+kUoL3wCKvDhKC1P6E/02/V0Ikmwu0kqrDIEFUX1uzs8AfXhEBwi3jhq52
v7UKCIaNqnOwCCSXUmKTdc0le5+pqKWnRXnuyGMgMMPNI0wtSuJ7WkcnuW1Z+faw
UCCOzKAYHKR0RaYJKiTVjoh09AlACxTKAoQiPAaJ/YgdOstUN+AG5tGZ8IY/w2Hb
klDp1NZ0dOaMjfzrabkw4xAVZpdqY/FFl+ySHdStVo2V0bytdSuijSGILlWsQALs
q6v4k6RpTbQjGmrxZYN7893Hoyffx1i9lNzbeD1vGkf0aKmSIwux2W51Fiz4bh1/
xIoYA3nKm/tShkrf41UpgcjYHECnHZ4D5qmhw/uJEP6TvIpLxjBXGhAedR25qhs2
NqedHcZEdMCIoFXKaIZ3gx6t+T0+wOWySbhVuNmYHNWjKXw8miesQokY6qt6F/uG
xdZvC+vOisw3kROM5rP4nNJco7h817QvalwIyXe/lBtsnu3GzVB8culV9n4QI+UK
eQgDj43MgVJMW6e9vUUVdbXktNilN3verkukIuq7moq2ndxe2wsV8+kfmRxi47qi
NmhOzFvCXPgfe961p9GXl/m/CsBXCWx3a1UUu+I56PNtr82E5SbR4QBM8oMZrHIC
yjeCSdipMQOaF4JmmBcJ5IJfW5fo5efDE2pV87nqKpEVaX2QYDNA2XPCwBXJgLf+
uwq2fgIgFzb9qNRj11AxoKmQZh995vCewiyAtoD7azRsBAi87VUnOirz0LHcrvyY
XRsi9t0jiSLUdnHjgvPm4JY5jjWczUgBiqCStMJmAUdH3nC2LaT0klyb/BeuHHUG
EX5kqjfqILHLbi87MClFr4TvrRLpjqhIFRy5EGA5OIKFcailpykUmOfSU8Fg4lUp
Q3UsRsNLwB/lcEkhihUVzE9BOCbpvz5vd2G+vGgUZwQEOdEgKo1w0q8VnvK78Suw
eYXQFZgELBLA14U0n5MA3swMFYOgtP/zeNhrvrm40SOpvBWBYuiKIoXS9bQZLlK+
AE1r0/MJUczHrYxNkEX5vgfygf40ifAqZMew3Dvzc2Mu0jk0bso9Qpm3hxlbjCqp
yNXiY5jXlyVI3JBW/0XU9gixRLmKyLYhJd76wTUCYCLDE4lBXpUnQCN/sFhL2zIQ
S9Fnur7A7gMI+TrPjKKWeF0dKDXRsHITjzjO+q/utf5BhGYaohZO1ROCgQfvh2q3
22v9qylqp0Oko2LeN/Etm8OSRL11BvvDgJOZvi1EByhtrgery03JRnzKWR2fA+Az
Hk3Gms5gUeNe2Z+XNTbXTVVTfFgHV3gJLbxJZbuAEKPn2wbyY3YIZfvTZuTOl809
FWVtUhCvVyRpHy+oR6FvYPXrRkS/dc+9F9pEDQ1/60o6y55OtuLK9BBBzApsZNBC
AyzT6aJyTD+BuVSqyuJn2bkUJfPDURWehW9S3XlUiRLTpKux3FLsoa8wTsEK3B6w
JYlYtd+eC8wsa0DdR+h73wRDsJo+0Tn/IxIkLmaCUZk9XFPUnwQBAxPAJC1b07nE
glqjLixPVha9fZOGfK/628e4xkFyaVeDvYy8o6ncTrznuP2LZP+S23nVa264PG5Q
UZ79UMTKc+y/ggF+ACXF+O9oGPy5JDNbKw6nUkeJgRwS4wVYQLvj3nIp6KxHG78t
5e7Z/trKKcEydlCaib1sKOBjSK0gsQcB9kP0l12Qy6j4YVyRBK3zdHPTb2pEDKXR
0iAChVkTqAsTxGpWTubp9HJkUJC5apUUTLv+/MCZNVC/TUFKPd5/Y6Xn9UmkljYw
aIIvmtk600gAx3INuCzCGTJPgi6An6zH+FB657sW1fE6LTRilIspnm73ppqXS4qK
8KFtlRfk3+DpTt3vMUWGTHsB4RoR+G9femtckpnThOj9+o5sEylYlxfhN4fuxRb9
3L4qN1aBoW3M2+gTRS5S1LB1IjkAI/hm2Q2wp1xG+JxrQSiNfnwGZwFO9YJZOtRu
w/fHKr4NNS8r/yh9UO4ZVCtDxVUkxLK5Qnuk4VAJD1SMjiPoZSKTTWfAyot5FW5w
NCVRxuuJR4mc4ikS0KLoGr/tFPhQDDIgfoNVkmEY1XE1UrlM3f1CRZMvQEZPBjYp
aI6VLIp45aWCYfIYitxA4r7+Qkot2xsMqfE4kaA3Yvzj5jx6Zt9V/9y8I7dBnKA1
BwCPcXOGb/6Pit1DUMunbt61KfNjClPNsnheifhcdGj22ILCi5EuI31rqpk1WrlQ
CCpnNihHEr+a2TGcKUl/OXf/n9I3wrMzIZOv37oDo2ufpfHXxfu26++6CWK6Nt5K
Oc5IuJHLXg3DOfLyGDW2at3Z0GYT8Pt127+V/SqJO7/oFV3ZhoZlAwb1DhB/GxuF
Fy5TGcqJiHOCV9oI9L+EreExKlgouYktjmcxl7CGjyz/3amhTkGahpvDJSQy9CnT
QZCbVTf8ipVonWKz+g6+pAj7TxF4i4++K1YHw7BLXuwizlWxtNI4EPPZGLrItViQ
49KLFff2mATGMbFk7ebyZpmag3QuBdpgML58lC2NPmM8tVFDMkDMNF1Jst1K9ieZ
vawGbJk+b2eheXWQdLfHhmWoHd8CfPno0ABRV6S3dwyw4FC+TPHMsRLiteYy4OBi
4f3Oq9eWORSXehZl5jpfq9abX2JMwwzkUOwpxwz+QKbJ0f1xjQn0wiV6YlDGPsn4
bEZhvoW3ZGMTwuqJeBpaWFKS6R5U3kId9KNfoq/l6XXXjseJzNGY1hoYFkYoJo6p
szlqNBVdKkx30Fnr+ZGPti80AEebwmm8KuUQY0J1LUN+tYIflPaxuEulo8tqpdaH
BNOWy63TnExKSuiIvGcgSR/9Id502mzijXlPo2/MdZih0GU4erM58fExmPf4GnIz
M1GVjpbaQRd4oP0zVQW+Qa6gSYXI8TSUsbQLfPzevj/V0Gy96KeByQxhhev9TT3f
P09IYgdm8IzRAJYH3sImbc3pa+tjRj8w7hMk9MkV1BpBF8oshAxP6bpNTXaJtaQ4
/2kqueHPF4UjUBGWti7DPtaTGn+YTW6jKilymaJqx5xBlVA71MDu7d/NhPrcQ/a8
VCE1XJM2UqaKrXSTJvIAv0A7I5y3N1V/KTT6td+OT83nkdNeaWv/+tDz4GGK5tfX
okDCfByCesJFjn6p1OKYefhjU4y4u2GM8TjgfDDZ5PUwKtjvoWlqA43ZqYGmpZYR
XRP9gg/ZzG2vL1wDgpA+PtIluGMW9mXqh3eCDEoTpdDjEYE5Ti1VaKik2czDUcgt
rBQxQEibASiFUxwvrWohroj1yrdJFu13302PT+0+ep/9z3CsOjXdoPM6ZsQGpBDA
Ej1OtY/ZiCsML0zkPHQTSJgZiNrT3k8v8XUUutOtnOf1Nra/0ZpsYX6/wEZiPR4M
U056gH71A8OZA8Sga333fIKs6+/afwyyf5irkzLL2pdxxdj9f8J8Y1pWmoy3tmq+
YP+CarsSCZRqN/T2jIt2rtRmJC0/oGk6Z6+cJ1cMZoZIFy9JPqFWvsBDRm2Bvvhw
+bueQZPx+K7ulAwIbSDBXy8xGsCI3iLpGSyskLClr1B5Q5O+ikMXcn0Vv1nCJBLB
L+pjvX+9+d9ZF/36Ekx+ZoQe9bb1t7jMtE4AcJv3npCVTZG/ymeIligDtEN38hYu
vYIvL8UpyEbxZ0U5lXDkAuRpEtRIWTwPRI0sFLVGn0wjfYlxP/zB2NRL3xlwxkSG
z9up7LoB1g4n/GPLYF7qyq0u7ACBo+tictJwHXGo/pMfpxIeGQlYHL533mYvx2Vp
4l4N8xSY9n5jpT9yCM0ds2PE+Y1K1U7W7TvDc2i4ts6BpusTQb1pa6/SEQHgR11g
vv2r0uDR0eTTm+yCQy1YOGWjybN4RIdtKe7eVQ2w2kukdi1LePwxW2mHcbTiBQQe
uxHHyhYJd+yCPXUD7DFv9Y2xIq4L4oUOcZUi98sKp0HOTKGNQXrqmWTzxfTNMeW8
zIxlZK7HPYcdwPe8oJ56ul9O9PufsLsCk33sw/BnfYvOkCqv4EZi9F0/Y3TW4ara
5JIwmYnHaQBa1gcvTRFXXH731CnaxWqzq7Tmzar78s+dmsY6CVBVpS3nYoIErgJm
8cPFhf5aD2wlxcT9zz9YJq2LDnk/iT0BV/v4B4C7uBAJ+1oyAojwoELthw4esDPC
FjhL6tj3yYlVfrD1nckzRPul653cSdZF9S4WAN6T1sR2DIgoLKsD6UnmIYJi9RNQ
/D9ggFKU4gIwORq3TJU4reouhH+iAb2dr+WsNN5QzQqiT6PRJGbV//Axmv3Hz0SH
FdRSvgqhluI1juhABOT7EBkLE/xJ0JduDFZ2NF8RkKp1uuV7C3+cmaJP0X/ADNOf
uoH4TpWeY5GAC1jiVe0mcIMve38guCiWfbHQFX6QsST+fr75uhYm9OIa5/hleQbI
JTrlzkCHak6J7yL4v4190olMb12QX2wp49KnrpSOUt+nGdxmsDs24t8cZnEtFc1o
TqMi97+HsOAYygNLBD3i+iWWAHfYSpstnD5NFYMLjGREe8QBNxE0dB/77vN7L/0Y
GOmO6zHqtbYDOxjsKJRkCarX43HkdVo3UFtoLGcrRTBvbhpzay9jijf2AEHGqowB
NDywDUYgHpS92Org+d7RQ++B/4/64Pekw+BxsKo/bl5PHJXNw8io8CTmCG4YqTqH
sa8EiF6cjZZq5eOGz+vRyRvDMZKXyOyf1ufn7Hhuw+EIXOtoh/Hp4HT6loPgwgll
GyQOr2aEjovSsC9P1xamsANoSe/SvAjvenbb1VrcFV9xhuXuPvY7MbnCVZyOGZOY
hD1aSRkUp29UYmFYXeouWcofniTklSAuv5zLBlRWFIzda59yzv0BN3zMgsBBux/M
mDYLRWjXlNKyfESfQIvAZ45t7ljyp6F5uXPEcSgHbKxzjLeTmJcOka6Gm83sD+wh
9LHiOMSAjQrzJEZhSXiFkFVR7NJDHOH0oMxn0lPw0Av3l8CgjiV46+U+57Td9DG4
2wH5prgIj55luHVKysBg44/HpVejAflsl3ALtGHC8cfAIevjZSR2jV9fzq2+6+Sy
QdNgcI7fkAPDbPUudEoEd+q7xOwdJczirwA4n4K+BLDCbCCJomzCY5iWzRcHGkJ8
gSLKD60iE1Prr6bMvSPjciGvy/MIwCb09QZk2vSJm7nRlm4dIE67DH4uVIHAygCs
2nejzTHxuIEBVI+PgAdx/j+o3WTq7bGlP5vFsPFYu339bZzRYdEo+lsg8I8cAq/9
YMLverb31ggjFVE5dEXarEAxMTwRvDVUX1OA24xaNolFI/w8pCl4qsyt9LetWl9J
5H8ZhBlopEvid+GdCIev+QqA7voK0Cu4zDWrqQvqYIuQknSC9kbSOeXS52uykXHz
hCjVfbD6LXuglge3TVqttahbe7kTir2gfebeH5aCSr/hk+nG/RHdd0Mkg9EsnRi1
ZGfXOaQ7kn/Osa9iHOjQ1YM6Bcm9LP7WNM0NTODQC4yBqtYSOsK+U6vzq1wVE19Q
GeLYRP70ZWKBmOY0YeOx7sM3HJMkZpISlQ374geUx6exAAqKBV8Pw41ol+lWCp8Y
f2lD0lUPTVGQ27r30ZsUfDLER0t7EIyCWeML1v2BwLF21Mo1NudiDjedDJkE+3/K
Bm/3RpaidrQ2oGshvhHSjQBFY6sEZ4rfqepi6bPXxkCe26ckueRvngcjFFe79eK+
LLStKkK/XAWselXwjwpQYHShvRPw7BS33Of5pC5MTSPc+SAp1po1X97f7HC7Gh0+
dqwogMnSVFcB6FWWuN56Ohk6Nc/8IE3klNViWA2rczTpfCMq2PyEt6IGS5yYondk
TvQc5Sy4vg86mbSiZXk8rUk+nBJ6xL8qb8SaYBBgrLr2a8vEcOJ0HQ1ceD/dP04U
2blPvnOxC+BcxfAJ+yS8EPm9/GjQS/iXy9yI5h/CyRknkF4mkt/IKNMgQcAlBYfb
ZpDUTYSfZ0pM7Om2elqOZo8bqrV8ntGL+YMLD1YNJflPKJn5CncYwYPLeRk682Z9
yop+n7RyrYYJuNRvGwhcUEJbDay7E7nbAQyMvPiHDE9n+rEvl1AqU1E/Bt/Dt9wO
jq8wsVU7ItpyH2Pu+YoXWkG91ZsZjxJ6vZNvnoxm0Q/G7iFzejkEC0fyLwAyHak0
1ACm61fbq4b1rIHCdOMdPmzOo4amYeV54GeshmUZgtg+zG74TSSoilr3gR27tg/p
Wbpsqv0MrYm+9HHzwbVt9PwQxjoipOVRx9mG2HiwYhx2s9YfeDqTV/bhGd1wA9vN
1WsmrIs91Bm2lAewdYRH9G3zoK5Zul0o53K2FKR2kZHdyYUOZCBO3ZOWhst2pT2d
+eEaT5APlJFCxkxKnohHSuVMUyA1pMBZMWxb9gyLkmn2WIepEXyIdLhdDrlzIkbE
+2qahFri9wFQ3lUKfIgW4gEqbSW+Vfw62sWug7sehUEJVUfLu1c9UlwWlBewVO7u
UHSuPVHAJlB/0gT+SmyB3hQGqrcfUygCjCrUSvgkHONKV6QjTmxRBX1rjY/aZDQz
0InE6KbbsG60dsMlSKxNvhsfwskQZnXJf+RK/LdiLopdY44IG3IICEtDv3uGkqBx
e547HNjdRD0N9mQzbXLRIQKyAqICUYm+hgXAPA6KxQ4sRY4oWGxhxzj7wi85OqkO
k47bRDDqb4WjbB+FTrM1roh8esHt2Z/5IudnWF778U5WHuulabiTe6GiEOQJbpjQ
m/p2VQAGT5W/2loecw7UjwQ7i7eJtZwyJgAYAQcr/fxhKMQeEWKLTsa4HMVtc3Ab
3yQt1/bNOM7QE3/wJkZ2cq1YHbp5LUHcQv0/D+Xzy0yVNcF9KJiTplvGX8y1c8p8
BI4lOl+Ms7FTYASi5Gyzv3xF1NW1m9tSZaCU0mpXL1De4U5jUOXuAbVE0pfk9Haq
zkdvCALoLZ6SLXcRJKLvg9+ViG/3gCCSRKxbcdvaLkezCamIFqSEDe47sfWF2wbd
VI2KhUdLmhpvezoKL2i9hQfjLVBkJNK2FydgpdsnHxF8xPSDlIoX/xTiS1voY/Ax
viE1FbOE67RnxnKPplUID9ndPH58W6/9ftEpa9bihMVF24Pttbb3AxBumy6PTRiG
QJpjTqBrijOoQMh26foeo7ooFiWUe7tE2bf27N4beE/3JLOZKPOzAF9/DnwTRfEc
vYBG2pSGJKulRlPKcs8haSiqtHf+bkh42eJL1ne7n9/MXsoos+OxUpRvUYRlV0Mw
/mbtcI8+3tvWprHdAf6CzT8UYmKdQ0s9vnqud7Cz28tiOR5as5SbosnU0urduq7D
bKRyx+IYJSvU5nw5r+58jPsqt1VKi0dpXpg2+3/hb1bP7Dgko5vqTMXzIEGAmb68
jICrYhGNMFS4PZvGumbi9G9A6Y57Avqu3YPFhvTuBDTRn9Bdx3EiEdYL6dKchdJO
j83mPCqm8qBnFZ0irY++nnx+ohEbZV6qi1hve2ymhBXNddki9HXnzCVlvAibmg5G
OOcRJmZDnJXhYMXHKXb9+VFVvWtkoPDJD9jnXE0neZcO1mDpSh7BoV+mCCIs33OJ
w5ZdRzj9x94ZGnzAdIzCXPxC/EnfObrBAXk3C3/C4ymoYXFjhDvYE3Y0HaeHE7mz
h6l+Y3S4b+jeAdtPLtVRlHBbhkd7qQM4ce0dwAPk4Awnv5sMTXAVr6rt0dIO4anH
qgguRHykUcj7oW7JdAKPwvxuLqqkb/nkp72QfU9rDhlqopHZUgJisLwTq2TMBBHi
JbpX8c6y0IeRCzEFMTUbPM266BVd1KmTkA20vuQxhu1fHWajh6GwrZCJOo0eNJ3J
F8GdirSKGDaZdyH33/0mOyr8K4faiET6Ku3LZxnljbAzOqKU1BCMMPkQmahESSdP
dH52zFOjXrxhZZg6m0o2A7SDrF3X3m8GwgNOYB6tB2N2YrYNz7bU9Y00ctSBclAj
2oY2+ZZc5X9wjOkyxIICjtjVo/A9XUqFooxWFuX0zbd+LRz20MNc3X4EJzyFhALT
ubuUES9d1sPzUUlfxUYWNQD3Q4tEhiHP860qsPKw0fTuIj2xb2xAK6JgyFSc8uie
S0j6JrGx4Iwq33WyIBFEfKBSnxSxrJh3v7TAHJvRcoj8r/adyVdWSVHZuhoM2j2p
zzz4D+YDvzZb1AfO1a5Ajg+Z7YDecgEqTqjAVgY54/CUhldUz5g71yp1mrvZMpNP
Zak7+1VVNyjkdL7xjqKEfVK07e5OhZMyDLsdAEAX91YHjNNJqclycXnoMoHVXtjn
t9U0fTtrbFgpEJg6RPDjF2dFV8gDwccq4/Q8Gc7akC8PxTUvguW0Y20YeFtCDWY2
`protect END_PROTECTED
