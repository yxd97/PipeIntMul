`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gRABI2hD+tKYBs4L5X74miL7DwY+9jLMHS6mLbK3k8f4wiPBIel1rBaV1x+nKetK
rmmUwiIGZLsLegmSkdgEr5TyZPPf/DdDLo2qqegazEpcpHwQx/Gko1gs4E2QZBlJ
Jf/THDBiHpHvCb0XX/VK2uuqlFN9fUuwVBrfe08djbMMiZTL4znvJ2MI5a00XZR5
GLXITuXlERfmG701wCgchzBICaikuLxFOgc9EjSSSo9bQx0VL3U3mM6MOm6kv9bR
9euSMevsMu7d37x490/CCGtNOXIehPCNq2YUYgt4qt3J5DBbubdl3//dhic1lOvw
SvUMyRGvLCtyT9jy5snTc6RLFF22gPf6ITQ5IrIb7JjRTVDCJkwWUK6pOJIwMQnl
U8qvJE5VdZY4QwfzLHowygSZWP4b90aFCaOph2UxmXwLfArQB+uDUkZQCMvIs228
3Sjbd7FUikPmvtxNAA/H+Lu4tXmxipQGJzzIBHQCYyKCl8AHVZ5sXCW4KDwZGMFw
qdX86ETBpjeV5WdhwqQDv3gL8X2LTjMG6kj8giqjJBIPdRbG5gm+lz+2i2Nlxqx1
UVzZa2dWPwE5G2UzxWuiJWyHpZe/QjDdwFAJKcqgBcFxeu0nr130oeP4B6+zegfH
RO+c+pKKEhIJ1dUDPTgy7MkMs2h//JDkDhZUeiXDzPINFq8lF8DqCT/+Bo93zMgE
8C1b2FNtqsilwXhNVVcfeP9ewRDdhusbDVJnS19oiexo8YnKg/fUJHNQ7FwQa0KB
yEDWE2hbMfwBvaw0nGMuguTCpjOxMd5E3LdbJvF9IBx0NmxylsPLsJEEZ7O4OQrq
s+/iURODauUomB3yI0nPEOetH2z+AHkxtPO2AcC2ovCRjFPeqJYr3w1jooJhFT20
1ijKEzV66arU5BUZB1COtz/rOQBqkhX+2oI1g8a3LzNKwGv2TAaNmze/P4JxotlN
hWEjcngNt0SB+PCcGKGzb+cA7PAfnz70150zj7VU+84Pxpk0JlZFFPMN7pa2qP9+
`protect END_PROTECTED
