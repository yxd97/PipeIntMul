`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MAFMjkmV+g6oaqJl1hYSI7BbQ9kQ7FdpMyu4KuRe/up4Kv0RJN7HAvWQKjEGHZOf
YToM4wURffrlDZVQALpu+RSK+81vXLsujkQoap6vq9ccP6YK45J8pnm6+ILtxWGR
3v5j+7csZLB0+/wXF59WFRaXsxVTmAtoBHYGCp9/t4nazOfDbyhdu/mVDzu0Vqhp
msY/KilJAOHQcx/DmTcLRHioqTYJizOJa0xTD9Xr0hcmjS0QatMt3yaydh0k5qKG
0ujwA/ODcm2d7wEzpLYVpGv01QUvQ2Zq9EILanL2TpOQfIumXHjyNE413iAuhjh3
IOgvNLYv0u5D2Ryp5pj/2xWc9l4SD/I7t8N/061vD/gWi2Mnd585h3G9Wk/mj5cF
0qxliSXAG0OlCt1NXpWUfYiiFaIeQlaZYAqk3KH4+Hk=
`protect END_PROTECTED
