`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FYReD7imS9LlPjb4dyfBzqqiQBgq9+dxgYKSLY8M5wk/fwq/1cznefOHM0TDTCS+
C+ArV90OKIG0l3vosEf3ubYhHgNJWcHTNvR1Y7QOWBS+AEld0qjmRd/naq7Axpw8
ybbpJ8tQC+AnkuVxREhtCNqKFGmA66GJFUYyFhMOpfMdJdGF8SeXEI97libSf+NQ
obeMUpcuH7/hDXlheyAjKAF6Mjvo06qOMNcZAp8C27umd41Xv7dilMjf4z0Kcrsd
Asra75Mez+X3ueI7zyk2zouwINokrBARRN1JCcjIkH256SSKJtEm2Gi0PYazL+/j
3NcZBZWolljzhbSripzv2kTucujbEh4H2NMf6FZnDYivn5Kb9yRiNZKyLTV/gPcT
IE9rjYPzi2Ke2d/HvMEwijvwZEMawgZlgDx5K2hfFzrZbT1snjY59qjoIi/A3JMT
O09gOX/yt+WhcQKcoX7c6DVKaRTneJiryerc0DoCdIUQJDxo3Zy+JLtjXpVCTtYW
`protect END_PROTECTED
