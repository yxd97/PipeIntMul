`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TmBxh6qu0OR2pW9pE/Mu4P71udo55ImUPejhQmSk/e1elQEgN/wJDxnuGYEy77A9
LXVnYgHuprk0qyhz4ul3VYdG+EQy9rBCSF8uRcJe+fLi8z4sUk24CcRjkS9JUvO9
9yvJO42Z9TXV7aXtxLRRLKvXS3YChW71L9BgyjtGfw5YLvaZQQuNKx4QkbTis1WY
oaJkNnyYnIEN0AS85SzlieVax9zxegJXF47e4H3HevnV2lCaIrCSTbrL8wP0aSYG
i5Z0bfMvvhfekNEJ/wSDrCL9/3wrf86pWf20FPU2xtLF/1rm1eyG1L5jE01vqzSM
AthEIyUMKtKd3FQIpJKv9ggoqY8a8MrtuHBQ39+KsGPKGRCyAgts0WspLbeVN1pw
ZHP9l3apiBdzkueEjKmpLjgzk9LrVVITiYTyyCIDN+xF5hZE6Ssl8rr0zVmrCAgG
QKBweHwr3EOPZALN7f4GMPOpysENZzEzwrJ0bqQ47QdDftcb9lqj3U2TsAHT0uXo
d+fci2YFG3iqyUUn3IpjMAEaokf6MOUkrjeGCWWxff/rezagjY8PMC/H7yhdbG40
a/oBR30jA5vMrYpjsBp/4X3V1LxovaHf9wXR9PnN9V1UsXt34MgqSB8s4blrOX84
GFw8Jrlc7W4BsuAhpsVUMSA46ECb92g0AWMZ9jwiS2Slc0Q2Fus4bzpZspvunnrx
uxomrjt9KH49/+5I9+nP2fSq7+wS7hAPBQG2hoTAMzJ4SshrfaB0+AOhrfAw4PJh
hZjbGO5HIgeMxiQ1xtNTTFvV0D6llV/vP+kCGy57srTPjI/j42Teb4CvhehxBDyD
bxuf9NcZVTWjBa/J7s/LNAqvFr4Ff7pnppkfoDOHWa+FGLJ9gmP7in2oNmUOQZ5N
lK+OCYdXXd70YUJZbn04ax7j3bFRLR1cJpzIS3IBvp593cFI+ARaFV22f28/3/dq
2NNjFl7Zf6S8TNNq/ll5m1AZWol4AgFRp2eELre5VXwxJSNAR+nOxLxAaYXGZnPC
cdS6g3FzWPRcpj4LjAuIOZpotkakwVKVTKWCp/Ujv7xxu1YGfDdWdXcwAx1PyzTW
vdO+n1WUIEwST2qD3EOYES/+Lscw/UiotheJEitfBGEdHxSWqIU+ZgXeHmv9dk5a
zTxMIaBFPNOeJPlxY74cFlSygBSr08gugbxh/3XJ9poKgrglWoSoKONrLfMrP5sJ
cQUsNM1NSxalQjNUdQFDb5i3098dMQ5MIK6KSRRUJN29/iPw+vzuvYh8IO0fdEhW
PbTiaWq9oE0uxC6dN4+F/Ehh5feKdwU0bSvW3beuCTcUkdXzrpTvOlGPhWOLfWrk
xva+XNZ8ZNmZfzMBUAHlPX1aVD5O6oWerTIH5YsU6BkybAN8plCabd17WzUMNQs0
VurE0pHOgRAtKics0DNWWoUj/BIedXqVc0cS5O3anvpyrpIlr/nS3u8HZxvxdJ1t
ZiGDxE9bVXugx3VQoTYQ4hpo4ioVaSLavVZr2d/p5/SrbD/nRL/mb58pxwMYbAH6
JKwN4yWhCKSMssKe3tjeZZWzOl93LSNIz6jtWK6hqZlVxyFxRfgwPL7uqN1Oom8U
V5kh1aXmeOKi7d+LyfpAWOS2UiN3udjfh8NLv01jobz4WdQN+rkz0FIZyg/YrgzT
Fk1Sb7h6OMppH23E3UTb3qpUE9b6t+x1A/774hn0WqOWs5owHuy/p7tpeX0k+9Ea
VwrAgnYtwVGl1j7wZ0lxPBnkREKjI9K1wvl3MTOfVeWgMtr3nGrp7Qr0biHw6Gxt
hXPwvkPurgjlT/CspSiz2CA9BnRxOgEVHExcYKd/tP3zAW6WMEOGPz1wHUzzXyuS
CpHBhPogQT+8J0Wj3RuLJTtT21xyJVHHEOcCvKZF2OEXul2aH7qo7BcA+sqex8BX
/76IGMb1xpYYNqoNPfH/01YaBA+A+EOHH0jMzszQevHSccHwbAwt8cmVM3iHZSmW
shbbSDTP3P1yx/o42V7pgpdhFvuc1jYJLqMiubkvy9FD7DrpYQikijXhsGS8zlRr
/7GQccAvDtln3rvLjvV2bvReuNC/2GNsijA/XbLWQqbCOX9PJRMKa7FUxKpyTCNi
7GpKiOhfCzVy1q1dis2qrCAuHn2aIsBDwVVL4tPimwVwizvVjMX7sC5IJxxhiCvJ
H/1j2IHYfmX9zbuJ5dwz28ay1ZVDia9bZFDS72Ql77/5soUTupdrmkjInAg54v43
akqOsFeptaediH/EsO+jGoyfKE2GrTdapeK9EjTbdMMkCqeKFMb6WBSxqPAsR/C9
5X9lDVjQngWgp2I+7gOw8uK2BG+a6rFORav8RwEa55Q1b6huZGBTLj1V3ibdnYVG
um09DBsN0PsXtZtvQZ+h5IJw+bJ2/D2G0rBQrClNgJy/7TvWXxeYA/reWMW2wcyX
gAID3DnuqXRNSLf0yafd7m++wc5EZkDuDm/utjST8n/0MjFuFFntE2KLzJX+cVvS
H+A7QGZ3MGbs4M0WrYWWYkBf0Lg1/mNitYaVGMeIm4GV4Ek9OdIrlR5LSctlPjAw
WQ47CsxpI18ZNzzn+ffBlP3xvj76ZWnQxNBpzcGsi+1nCe415Ne4K1AmuhbqmK4Q
cXy9zWoGI7whO711SF0phc8ky8WcteogySR7lsQKAolHso0Nq/Jy1D4JQTbfp1fM
EoQlsjKL0O9K5/l45pU0+wZorU33pBWnk+wgV/t3H3ZB0sRKtpD9FRcNutJwUs/d
BVwA3Bzs2tfnzOFcIua3MAHedLwoCpNikPxznL3kH5+Dzz5RY0R0mDl5uumVKOSc
TwgdibUePd/Ci5l/Tp7DQwrp5DlK3uHDW4QxlfXEWCtB2S023wvYrgjG6Jipibgp
XhB8jYyWcf2RMvzU0oTSrfxaZIE8jcnvJuSxZa5ENYw1Pg4g5ROtfZ/71Mwed/m5
FGZq//Hn/XQGvytxP8uIoKKOQ6ifr/c0Z/9DdAtLMVZ92USZE4zix+IFmFamcGBE
97D32LUNDSDi0LySitFXsK8JvOQYfCrCAxJAiFJ3xOdfCTH+tJBrIwkAb0tG1Fbr
L+MmTT9vtLapx5aRAtE7vp2m6E3/lZUJA8MWKZT2l8jA9jt3osveqDjAD/C9Yl02
prTcBNXVYLbWgxSKwno4MOwvx9yNJjTtlkM6lqtOjZgEGkMEIUoRrwJe44nbPSaj
B42s77TbDbDkf4B/mbf5sTDcIZb0b+BWk1DiNrMCpoh4VJQ/6axuqKff8jj/kfAj
9KeUNkQh4CA1FqFUO6aYQ7mgzmhCqalY2YLgCu2iX1wBzWOwwE8dkOJdwyp0Ielk
+qotdLk/n98uP12whbetNwox1P/BiMnRM8DcsQKFu+xGSKOxVKhr6RMCmsYQlHWt
jOHxROixaDD6qI/pZ7OJRt5ZZxlbodoMo64EOVlInIdZutv6EwJ2GjPdkGEg58Gj
vleaRHJLNbReKEP+ToLyCboSPBq18c3rzAuKu4vXNzNXyDMKpth5uxuanO87bqft
uzi+KXdQT/sdoQRCVdbQLwPglqihwLfhgDe1F2Ft6/xhXKHye42wFUI/Ti1iYjPh
Nky4L5cuu+wpf6a5+XPlDAGU1WTtR7QJr/PWg8iSaJ5EtovqZVJBOesW7q1yZCIu
URTdEhSUSCk2rRFtIZkux443+ZzFTrl9gRZiI/uvTLTR3ntfuA5Cq/GIYqG0F/Fk
ZdYHhIWG7iEyDTDFV3I8v/V7+gxlXoCEv37o4bbdM7NCG7nYeLRb3eD39z4TRP75
CF2r6pEZwfqKzzgW1XW5ivr8l8fEnEXpsgArRwMzotLTe0lYHI0bZ1KPpId+ReEB
+L4q6Jtb/VMjJ1flnSxoMKTfrEaIGynbAesj6PRO9ArA0QcC09k/aibrfkFaZI9p
UM4FEF0kn1HtEFjobTPIrcmOQwHc42ejs62z/uKA623wh2W53hpG9Yz064jZqdGS
lQkXE2zYj/3Q0B1jscWiL2dScWP3fmzhLZBj6RIhKp7A171NOr55Z5UeSkgXl+t9
3wc1jzNPb01hSVpilJ7g0LqSS/llYY+nYxarJIq7n3snzUT5jamnobVgcc8uo0Kf
iJoygJFXp+oqhG91rbVo4rMZdY/wPFsWDWAkyx5OZV2wF4VrT13IuiG81v52AM66
Iqzh8JDF/andbVY2RX9ccxUM+7ElFjV0yhcrvwUQ1iY90J/jQIKSJKGubaRPJnct
0k7R3VOaaQqxzJOTJPEJUWO40306YBbDJ2FPUhHuWP+frWno/nC0Qm1Tptinqhiz
`protect END_PROTECTED
