`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C387en8S3UCCDLNFyMh8d6SCcGipjCj9ML7Lu/Er6of2i6Q6nFOrmy1weyUyU0kM
7qbkLj/SMJftni9SVL4dHx24aQkaDedydBy5Pgqqlcx65Veu2Nwber0I+xkqlqGp
b5s6smENLPY0XOlqMZo7eCMmXHbWrR7zBSdMnaML69ah8UrSymbduJIcXmspvCCG
iEgRYhTpofL4gbuzcd7zYqFhR6ywoWRGq/pHwlIj3MUd9s0D1uvzClXctDxy1j8V
kiC6d/Z9o10Vn1gzEECdmfUD9OTm2pNaheW8Z0dEuhARCgyhtJqVkoa7AyAEexFZ
QCQwSxeUZO18czxFqwIhZ9CTW4wRK39HhYucV6709bohQcZc7sRi/leA4+bH7EJv
fDQFfTrSSVEhZx70ROSKBWjibZI82DkcXVXolWSs6GSPx9dQ0Kg4RPPXhd8wYjrc
hv4trklzDdaU6MKH9oYJpQ2Y+GMmhLhd1zjBuAUmEeUjdgipWbDNH1/Rcfxg5yk8
y6W6OiZTSvXzIsZIy1y++QYnwqIHNgKl3zG2Mn+5/fWJQOxWbFKNvNYLzVSQTLM/
/Y4pV+zfxr+u6xVKOvokgg==
`protect END_PROTECTED
