`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u4lvrszd4ItPLMCqCWpJ5hKG+rdZcyuEqHlWORpZ2Yjb/pA+aILOQllJNmfvLLmy
OzoMc2tC4wYlcRc77yORCj0clXqulTUuvMvejyHwURCl138ZegabxMkdcoiIN5Qr
LXRp/tVvMsWKTTJwz9qcyxp+jbAiEbtyB/j7UsM9RtrX7WctnjqIH7mrybxq04x2
EP/CW9/MnK7H+xO/unResTPmJ7i4Kkz+gd5QCmgJi4eZ/rUdwunEC2h8gbvfYPIN
8iWIaSF5yxPKe8yM5uUfNPeA8yp55Ej5bFU+bmqgLdIVQZV5B47S+U095d4hq5Iu
8vLPFISXYJt77VMDA3iCDDk8E7RVQK4VKIlb3JsOFocU7vZIDD2z8tDfVAc4zGQg
O00Nc0Iew0O2PwSAP3jSt26xdDZYn5i7MDeoOgHJIcHQBYpAWmKv8VqMs5tOCMt2
KGqOHAxrJNYX3qMX7NkGNaetzIzeZwvdejMTcR0If6fbEF+3J9goV08z+C57hj7N
hotHF9TWSbYT3laLOSdff7itRjujfeY3IIMqFgLyLRUcYbutWWjGvkdPFTrRfqby
Ud/fbvO8W1JvFuS94j7TqoNbign/Kowlo7h0fMTFhU8Uw12HGR75H5vyhiPRuVWk
PFRE/TjJt9mbDn+gSUgHx2RCVLQBWWtQHFi+5ci4sA9w98JisIUIme7ZUHQbyG6X
P8yr/RU5apHrSVlxInFhnQ==
`protect END_PROTECTED
