`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SOieOEuAJGi4ZXO/BktrP8hDwJH/mbagUAVwfYdGBK9MTo4GWCVEO6JaAl3PXItT
D2Td7Y0s/8p/KxvtVb8rL944MYkz8OZ+BX9yt0+bjNfNWoc1wBWFqCblizSu8Yfd
3SS5TZmNy+uyuLqVCFKbJPPt0RwGOsOJ+kDsa/RADB98VnNtkNi1+sl6yRb1b8M/
KAXw/Toc75A+8jH3pWO3Ki+H6G4ZfHKsm+PBOnrIEHrVid9y9njBg7dAlQ99mRjc
PB3Gv5vLqyjhAPVNhiS49BJDxmAIudSDxFuxfhzZxzbLoizAu23mCFgbLVg7o0Ax
IrXHChIXezlfc1rr6qaV9n/vZS2zVYqIIrKqcZlnW0Mg2paOGiRpZBv/dTyG+Xmi
Df8OCQ/t/0SsewJ87OJ+uGRd4mTNuc9kYFrTz6UxN6YcxXi4D+5bEzB3B+zrik8M
2C6IHX03t6oFirvPagqTFTB+MaTopE9hy0D/heniegJc8YmIlaKSP1KnR2HTPSwq
WJKPt3iVzKXcvBkUJoYWog0b5Da6q8OuO1xQHhH1xRrPQa45vx/r+s14cxOHWZpT
WkSfFz8Cys28HicdZ9bb3SU0xGuMlvUqIbLh8yg/I2BZeneS/zdDdDnW4jVLwTtG
K9AJryRDJX2Rx0j8sHJPu/Ul85g+Pa72bl4/uV3MDonM9HNT2BkdUopwv3iKNx01
/U0cBuoRHqmYLQIuZQ7FL2wxHldICu4UfUD2LzEg/FOB7SSvkB0e6zuZyCmw2etQ
uvs4UqN/qNrjniHQqMHa2w==
`protect END_PROTECTED
