`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NK+23Hy60zj0TsDQUWLN1Z2bbuhZt+soZb3mj8Oxu9lOYpGQ7AB9OQedtOOwfWaH
S15X+8n1dk0T5BBF1pQS/7EiOoizXh6viYPH/95Tb9OvEzgA3EQdq9i0Zorz2IiC
7iFc7OsEVox/0HbYW6CaLF0sSojx+qTZ+cVRFP0aHJZuK6OKjdsgnnKA2Sy1zliP
fQAMkokXoqzrmM4oThh0htD4Js24CVvs2O9sh0ePNK8BYWeU+YTM33BTM1UiSjZ2
iVbwdl4A15l+/ECJS/9D0yyKw6icWt5kUAkLBHSKqfFMB4Zm7nkvxlhuADZGq8Um
sjmhl/QHrm+m/gWvWcy+LFZN6r6vTv8SKihoaKm31InJiMUiKcISwiC9dlxFtPpZ
v7siz6geuVN9qxBKkmidAhDfPIqDLxRh//ndsCGk9HW4prCXUW8kvszj9d5+uqxK
s9mVi0y2i759aytZ2y4R7mUbNeHcvBoIBWvuOJ1dgm3wNGQdHJB/e7GqEbJA9dkf
LoPbHw2VBL+FW7FhLXvO2f2Nzs3ghCli+pCELoI8+Uvlb4ZSBWv0EAjRqEtRuZxP
SIdMYV/brxenNiMb8ILiFr8R1jWuzLBm1pUU+zq+zSI=
`protect END_PROTECTED
