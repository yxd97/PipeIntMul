`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HV5GFOdcQ5BTnuq182HoLFRRY4PXebG8FlwKuwkZ6aRQrw8fOShXXlsWXlQFZGSg
YVH20MDgcG0XHc3rVXHRKODALt1jkWWHRs8Dg1hgKhY6arJzDGkpWDNaLyovehgQ
RsyLxE4TIcgqCMg5o1HX1GF52LcWF5G0W4m+oVitqzE8yxq2pUisGlnz8cgZjVIu
ZU4l2dsw2pAAQmbVlkeawDzejbTAPEzGqhdJTGMl6juQMtUmCjvlt6fJShWmjhDa
Dp+lK3IMy9caUAU7xCznnAvWgOIqSE+I+uJeeQ3Dl1BUAFwLi1bIoHAnVmtPqWhW
VuWjpoUEDiLR0+DlagZSAN6WkHxF1197wW1pwkWgIYCFJG4S+e6G5a5LYRYiiHE/
VBiJAZrSJ/taGIynPWQTuTibaBGYYAyVKRoyEGx0r5pBmFfarVm63nsCMU7o1nWt
`protect END_PROTECTED
