`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3TLcXushjrhg2mF/pCwvw3rsxn/oag0UN0RFZ6qSn/kb0iobrZKe9KL+63RZGnz
wHMEn2XOIeH4meQmR9TwNvpm7pHv38dr/qLYHJfd8JmoCbXrUUfBbY6PYuUoemWl
5tePAAF2AWIChPFOQdS7ZK/q2u0QRc/ZHQsqG73ah0yuFp1ppakblDPImc8oJFyt
brJlo2fwhZFU61rVkuzHQ3Fi5ez6m3Y3niqK2EtRrU/O1kWr1NoScODKP90B1/2O
ijgF5SjIy9lrj9n796KlXSam/hvBpLUfGxA4ZAGDo/qZcYB6MZXXEPbIx+AxI4/8
AlL3Q+eQgax+iiUsxUGZAf46f0+q6KbC5Q+cDS2547F1CyhiHR3DKeOciKaebmDi
PV2o76wM36vrWmoPfbsZk+saoqzLWPGdBbgFOrBWl0C3wCJYXbWwlo8fVlqjb52K
DuIQd9X6FKJXJ93q68aPhdBcPuTUGxj8AhmlczCdXl8BQMuKo8MNdzPzC0g/GIaj
7CVjcLDvvMT3NWISAB2msvQYnyLYR7/W/j0VhVGg1VU7X09+/468XAGTveYR57Rv
m9JU/O6jgcQQ5MEeuGM5mjZMhMSyfgmAXarOnCG99uqctdP4/ZFQEgO1TviDsni/
EL95WPzPBIvjpf3xRuqa/Znq6YeZcl9whw4ectxY60fnpNn5+yAPGjXuKvRuNwgs
d7GTD053EWA4zKlw/z6b3cv6o0udQSoKTMbKftGtqs8/If13tC169gcrdQwuSf4U
zKGxuUKMAw7mwQK86EPTJPEPqARjG7ShCAL15zW/c7vQSIpzIe7RD5LknMvGEzmA
JgGoAjQKWYN55d5e+TL0oj62Si9h80o0tmzaE+U+YngLq5upABlu5kZwyPRLo7d6
5SR0s15f2fk2nGZsjG9DedHn+DBm/5f9c+zT9TA4lUWqXkOAlmdz4u1BXQZIHN0y
hm5LRGDFJNcanu1pFoKhUNU4vOhI92YhaQiR1SiraAhMet9DVKa166XEdlkoEGWF
V/PbxCjAD5LVEcCit6xaq/jfh/1hWmxAfT1nE11sMOAyfRWPpVNJo83IFt6gERJU
6k+voL5oXkWK7LlVEoWOvVAsUujH8tgW1DBP88cm2mNmMtl/CamAPRrcb5eefZw1
87x87D0Q+V1T5mKtr+DW/+lWRK9f8Ju18lwnDK0gw5ibp28uI9VwJBwLvATalrZM
lMhyDOylUs5/BA8Wn3Apysh5FsvSehxPDDv1RdiAC4F0K41iG/eMBHQaBeh5W2yN
NkYtHlkjtOMUjhXfUIT0JHGrd/NfDGCGQtjeeLrcrBkTZagTxDdR3VkWsf+++QU0
RaRwtNgMAMvhRswlcRaTnBPTwclasfRbS2/0iv9YuFRP12EpyzSo9hQr+gsaQrW3
Ne9EJnrh5VXXvxqbpoMiGZVnbp4NgnIzpIgnj9jGJqVcQP9il6tdhW4KR90peMOg
ycuNJ3AziCKjHHSXKIASeegBu14S0P37fnwbgvYPCmhzU8IXdFisbhx1D/Ftotzb
k/hY9FSR9+a1ZyBPfHsm2lzxhehu/72P1aEltcWqDRx7Bxu5+JXuPi2u8xI+ZsU9
c5ZTFYDCagSJ/wVW/Cm5vA9RQVWVUuVzyld/m68oBoQpON0dH+lF3rqxl9By3ZFV
514/3gxy/gc7lwkdp8bG95s60ZbPIY83VIk6zjb98pFRXz/aEySZT3n9FDHOHtTz
Fl/HG+AP2UR5XfpB2C24DHcieOVoiUuqUiUTcj5XEQXPHcuHCclaH3BeyHkd3jXV
KSjRY63sNRt19PEzTm1UVz5g5jewXR+FcfQAg4L9w8c+aR/i67Qm6rvCcbqaNQnS
YuuYmFNTnBAtLIT4GOQBZZEYdjais+Tl/oF/W2qvou/tLEf4qQgUg3k4gOPEHLkT
ZIg4uT547F7YmmofWbbOg8J0OfmR3ahuvo+mHo7GnaWncSRzUYoTvumRo42u5r1v
41oORXbVTtx+yNPA/jQeM9M/TA56rP4I7eS3uC/tiGCHrd35R5RlSxTXY4fxklxD
cniV0LBj1zRhCetJKV4My5JE1XygYQVOnN3XUFoxWZkMBIRAieopcf3utiu+d0iO
vkzavK396rsjPT1NJAkuCiL8wxGaRWHwfCOIqDt7SfGyQ6V1+E1blrtyRzRt2bUu
8YMHONG/VzOmzhTDf8V7TubUycyCSKjbA9/Qcw7yPVFB10fGd4Frg/0FywuG3ZyL
hS+MiK2SKkAzyLsSwfhuh4dHw5bBkNPxqXN5tQpjCmP04ZjWhBk0CXkES9vqcARj
dJ1UTNRuDJluAYAGXEc1BvSIi3Rf391nbg8x+aRuqYqHHazoWYop8ocnUOlbmd3M
G5R35HkyQTSQnoQXgwDAD+icpmsSF/WssyLdLX3hQNMPrjasnyaBhQP+LHrJ4TeY
udA7y+RDgsxYfzMnpxxa1CrSjr6ywRaZ/BguCZPVinP+arWmOIEb8lebpvEkEnpu
7z6Ku6VYCes9TmkOzdK8K0H4F9rYVojmFVv1SuIyWAW1PkajRoC1bcbc3LL5wxiZ
YSW80J0vHJpYMOARxIpkY7cpWu4VqPRCmBXpE0GdWPNnkTH9vCGHJ0NgTI5pIFyD
tdftiBaQjhD1mmJejxPYuwHixPzAjTTwUJZDqAHyNngHrcS/sM3gQGQEffp6woF6
CyD22ygk08FlaNBv6Hlj4/pFaarwSL+vQyMyrZqguemip0pswZaxpIuy3xWo8p+H
lBNy9n09AB+MTSLan8BvHnQ5r9cwd5Lcf9Mww0Xp4DzaZGDiaGbFssqiAAYDRpbD
oG8AR1/uxhnhXgAqKjU0J4FDaLL2k/behAfux1qB+XsPvwQf8+2nDQvMC6iQmgK4
yjHIdWGH9O//DoCFYdndiL9aX/CDMxWQtJyR8sSvYL8CTGO9E3Kfw3FZmxGBAh5v
zLMRnkqvzy22RvHNEszXtWzfgP0ikk3kmISNarkWqugGo6JNs4DYFRR0KwBcLA+p
ENiWn2pM1rzGscfx7r3W0j+C0AhBVhlTPp3fv4Btu+tileje5isiiiWXl1EEr4bs
wWoODLE8ZLKoeq5Rr1YZeTIs0FjglwXGeBiz/B3r4BwK9fxhVF8kuRcWYjyaEcBn
aq9rDimm8Rmo6O4PYvjB2O40JHleyC4hqRacBMmtDr0g1fly7pP1lvUSt6TL7vPJ
mkBimY++KnzvDoB5Rxm+RLPzO5qMTLycv6M3Eztpva9gHGZz4okBrTo3VoQtIwv8
a2ZDgCEx5eWKhVw8LvE6fHQJF3/QnvRvjCg5rJ5XYfwmkw9Y0U0R0cEUumGOdOi9
AmgMMrwmX7JRKYigIKV+3q0NZ86oSB/D/Ys2+Vyo17hV/52MbbuBSDjZo1s4L5LU
wyCQ8FKd2VsDpT0dCbjSjabLHqF++I8NpWtnFNXQhkVPSMggAb2Zaa4rx8oA9eDe
vPJusgp0HXTueKBmvHBfte9JjK2aajd+i/vT87j35ncZz6NQ2gq+tstsgyJpySoO
ofNfz4rp0/sAI5YsPykD9ggtQAp0/tbdks7btmx/UP+1kL4H+Yk0QIi4DkchhFtW
RXwS0r6IuUJ5yZ2opzNuq9QlJpXyZRKMNavlpK4pnh+f9mXpC97mcxbAuBvJ/hRW
RANkFGucO/Ss1SciG9Fcb3i78z5WRobx/c63giLFP57v7LI5Kgz1RAt/X1wmAHpD
v1b1a6bGS3+SbWKRxQK7k2eOV7Jd2ggzYNThGTc/dwIIDY2TeRR7x1/g8P3Ro8PC
GsruHIJ/uMLUmMT4/Xr0Vqhun4RxqhriWc6LeJXWJAS+aVMLqaaSzjVdJCp4Bu/e
lRBDeyJRwEqumWnIuX8WnBmMcq9bOFu4GAmtxNOKpgI0t3dVjVxjakcIwwgOCs9u
7oxixxAAEQ+uB+7zCCwfrLQUl9j7vcsj+/4od+LXsVVjs+lEG54zN1gdW26GNR3y
F/7PjW/wzg9SaLeTMlOuzwnzsBm6D772Vc8K6+2M4ZIk8a2lenTw0yRfbPzp9PJl
kWsr1gUnnHG5fMI3jrC2OMq7DnsYj+jZuejst1mnUSDSsYkHFQ1v7+u2Wsi+blWf
L3l57jtnKkzRmcXGWkB0X69KOOzVnkFcKHwRYuvxl4YVKmh9qUvAnFjn88p6YXOm
QRtYC8FGN3z78uC9oO/S9wxO1JITVb7YIYj9l7f9v7QX2jpZx0xpEAhoQWdP6QE9
MfBcTsOW6RIxBqlH8WZAv+yjpOTfh9YIv6E8qjA+FzfPyjaptxrav5kwehsjyuaW
Jll03uSDU93SoXwd4tnxXRWFAdcca2ws/GK8DKgshYxwnPxlfTg7U9OSSkXkj2VO
UlSw9wzxtVrgPx9YyXAC733gyFTrrUXLLef0RcIJCBAyBGpwXBg4h9mXShz4g/q3
YD6bZehRDBqfLklwgowUP2Bwek9kuw7XhhEhyAsDWI+uttfcBrZmHMN9uAjDKnea
xLHDBjELa1FhMR5vAfX4YlCeNWEk7bS4JE9S3SMs7zKsNcfJ/pH5Cqh4whyxifZg
OCtehAricW1IHzDHvaPoIrJb7bodV+uu6RphTfmaadmUwflD/FbgwqV34WnsHNXw
o/5UqidDN9QDngUlcLrbyEapBbewm0wfjSx6uUyYwsf+1Up6LrHlF6hNMuzux4nR
pisAZt3p4Kt6rQadlWw1YxpaQR0ayUCA1aO0hpA9Oey4uk0G3mJFmgs+4RJd9p6X
Qpyvie33z2HTWcLZkAv5XMCxh2Sw5iD/76ma2QiPuv7IkeisEtlEZkG+hZnV/dgH
9SPtrnJOCq8PelJ7VkJAcoK2JUGkXJbekKw+Phfc8ahBUo0FHUf8U0VPkxGT06im
btMbkWdhg041N9WbA1V4TBzyBt7hGX+C9/fjLEG6IhEbHWlLODwhtDjgKHXep4WY
iGAjgCDUWqI9nHvB32iouVV011gSYpRXN0Uh2e9UeiJi04iy0RladwJTxuAAAhEk
BO9JxzVMILU9ZYh4bIHPDyUq/KHvlCZSQjHVpxDydaOvokILojj39ZAWxQjrOaD5
03NyKajZ2GvdaX0bmdIJVrAW2apAILgiMVJ9y/twshrVlhUgogLcJWecnMtMprSv
d64eW1lhvwD5AQavsMRIGQ7atxeozLjRGPp8NK0dJ2YyGQ5BxxZNcj+7pP94BCAI
uCcWy7vflOtlc4oJPfpkX+iIkow5vwSaCfBgoJCb65wJARRvvpWkQAW+LcHY2VuP
BQK1lLecS0cfGTFhl3oP2/17PfWPHxWoQTchCi2nMn0Fk+qTJ1mo915LEjRYEFoD
GgBAjRanWCMvzlycSC9u3fkQ6IbNZebLHTWxhAi5VePNsJ2UG9p8tue7RQBE5sl/
FvmiUpLwqlPfs2n1j5hzd0DMyz/Hmd/cKUA0ACwR9eI7wV5J2eNb+f01Z5KHAWMd
HaULFAXadjydXZh8rRyBL3BQiupMQC9ZeeMr2tL1zkHbXRLsBfIM2TtP94BJJHii
9c6gu/g1exWQZXVHCM3a/qG/WK3LYeVdBauWIh0GqIoGCA00ltNEUyOdLnZ0+V7r
nTxvIoGaLhvVLmlk7XAxbrGHdx0XohJWpGh0t3KyRfpFO+bQC/iZGiFF0xu493Iu
2pC7HS7TfUfFV95pTMmWIfisSge0U+vjop8fTnund4f5uKaRa+1kU3HEPRp0J2Mo
MM1hRAzTVVjSWVFXFUbpdUURWydwxX5Eucsi4nAXOaN3t6a4Ec1lnOT9FO/ElitZ
K1+0tjoHdok6ctrgRYaSZl6hi0AGHn3LAeUEg+sb/FhoGGxKgjSOVZTs7IR7vyVt
DGEUpvMFYyeFJUuk3HvdxdmzoSdE2+50QPLPqFVljjZDAD79QNoDkNW7N/4vXL6n
0/CII4aFgyCIbLq6qTTn+zjgT4fzdSRcX0dXi1XsP6AgcNZ7zpj1wAnQJfISY1ei
1WFR17dZL29aHmxnnoayzNd2PBxQ3WbWMIp9zv1qLELrazju2YUGskanfuzS22sw
S4LKCsClMNKsdcWe+blWlry00OS3dbbETAumHaJ9dZXAaZXwxNTx9FgPzKmgbkAT
TZlddUbPKtgY4TUXRkaACfzgiQxsCOM3v4hlpUekwcJ+F9hBXT1tI/Ye8PP6ML4t
ubRb5qOhnJDySoqEg4yf9hud2Px6oVvJ/JnMIdJba8U1JU/IKLK2qmPViI0LhMcY
CE0X73RXzgF/h6Jt+h9lhpdl//jEOAiTFl1VQMH+gEbmtkO8AmWNBPhyGYDRDTk/
pKsbLT7qJeU8Dn3hGTIvWrEkXdCFiNsWVVCirDMquKFMkgMTsC+jIKFTeWucvzw1
MI2Qzw4j3EovHc5dWMPRqVhvvgEGvEP5Sg9jdTnemVzHWsEjMqu+7JvqmC1YXdot
bCWQTwnZk1/pcrlRGCOIPPXbU+GLZf8WtALXKMpiCT4mbdG6PsxBjzNDU/6VDzt4
B5XQwqCk+7cKD5Nl69LRkQHfGd7Xk9dN86zFzqmj+hf39iMs5SzoSunrbf+obU6J
VIQNKKamqpZdmgaIVx/HAb73LTlmanWa/fFKnqaPuUxlBf78iJCbGeN6lkufdyXU
RPjrrCvQnVBKjINHptvR+3wwm/PoW1Mr9AbTjbnn9jlvG4Z+UDPZKcjQ48fwsctf
3heXovOpC7xWbl+J+bEUP9afwuZjXg/pt539OJ2/6CNPW/spSVLyd8yZg/JoRAaa
WG9VEAdLmNJHrQKc6wvtYR7kKPevd3K9bVGrwpZxp/Sp2MjslXo/ukd5fFrH2fjp
ytXG5D6V9NeapsUYwZSHV9v9xCr9+xGKoe/IBWVICYX93rOWsz926nDCq+38S2Zy
kRc/19QV+8DkxZ3w/tsXCuLXrVu/6kctUXH511WVfHbdyzB9wmii1ZQA9y9sZ2ut
/nUk7lmS6G1v4Xvsz/6dMh8mysGAz/uzKGbhMhtTL8y7SC6K1A6RFXvbrFvU/BaU
jgd9kHONNGbwyrFYoap6v5zUt26YhQbV5fYO/gLXbfBQ2KS8DYg/ziJ6K5z9u2eO
JO92hNtSqhC/tliZZxnewqsVs3FghvZYLFZm/NfMe+JIOM9eO3x8HLQOabYfHTIf
uVwrV8vXYcoNCj8+HXraYIDRNQ5E46ecB2xwB3sLXwzmB1PIlx6yYIDVeZbFO1AW
1PWx4jG0jHVGM+1hguOAHIM/745iuRzu8VoTxeo/ECqyIwlJp1FeVWX1HRuyEIC6
LVLZwe8G4XW6j3YqSXcLPFUPTvP/KLJ2RudaBxZdzE0C01ybqtEbDbpdTAJK3HhY
qcwvZapaXUTvg9xZgKbY5L2PDIrPT7XPOyA6FVAf8xs9EI5NcNoHPVbVN5cg23Po
JGuD6+Q0D9NgTSbo41/6LwGvURe0jMD/O6Me3mWpYgjybrysS6lYB6wdwd7E6kbk
Qya8f6VzPh8fR0pdLAYJv/l3egvP821xNPc49lQchib7KjDxs1HreULmn/7zJajp
nrxVDrW741bXmM0Y1XyNP4dHXvBhyXc4Crv02jOl+wuspA5gl+LxwmH4yltRT0tm
uZSa3t20i6VkURjat1Bx65L7j9h+qh2sBmGZBiQ4GchcskM9m231lc7Txofb6RJx
X0kSMeMIbN2sASO4a63tDpwBOsGu+Q7GSskbqGkdW/q+c6KvMlaAu75FwTquie5t
pAtUV9ORZROqLAxyiYcmRycdnZZoNMuAaC85jInZAjElTU1RUIdsr/pcZLoJDTdm
o8nyn06grHj95HzKrK8zstLTJlqmeduMrlpjAl+q2Kybx+4K4xl8UgDLoo50Ub3b
jp4gZfNDILivJN3lHRov3+rrhksojs5qi/Jk2vat3wKUAwkNTC+x6zr1tlDEdtQp
kZU450R0NBsgvV1Oa6a+jJy4vQL+FLUUbOe6y9U//+XwrcL+ltYMYvyUrcF9afRG
GCno4/ixW0bkRqH8bGbXC3CT5n60vePCOxvkYd0SjPyHmXL3mbKdxxNBJS3l96P6
ZEKdkwXclt9ZZ7LUwkBp92n/xiBVMWLOz3VzVmrUoOHhCFqYgFbIU46Mm2mgQKyE
5o5YHl3wVnsQEYvA61gxgKtnaIAGOaa37ZDoR7P4TuQ3sML78l0fQ8nCbKDjj67s
QOpLYst4aAM4PsRNtlOo2+MHaxvB3WzaCOE9HE5JJT4PBe1Jl+6cZSw68WM67yad
PQKth4eX7WJaZ8NBd0l6vImaCzgo+wMrynzI25VlpGbAzTqxzzY9LGs6bym/yeRa
S/+DryCSmqm/MkcfIOtTso5L5gdR/u3h7gH7ALeODYDdFxu6VJIygKUKOTpNH55T
lJkdUlKvBYh0kukUY8DNw8wonnqH2hT/6ing8GwAbbxCqc/6tT8Y/ysptvlETmIb
JlvMkWAEXn4jjWogENE4ONuwLzMuZC+TpexkdHfmmlYBaSvzoJQ9wNxC+esHB3Ru
5d7rQ6ED83AIKUyELQX+7RWC7Kus3tq5FJT23wOI22wvR4eDN5O9zTIkPllHBe4d
I2AOPpUO/+YJbhN8Ud+0NoQ3ZK0kcqa1SjzGi9MfIA1sc0Yakzn/QMiNEWVM7d4q
mcyFw3F3USHn85KCBF0LXT0+J3djg5coWjJEQlrGYsGD0gMF/XDVzMHY+QHl0Z30
iWSjGbMuE1stLH19oO5Ovq/w3ovs/qiX81SrmmTBMNFvWfB5ASyJ8FHsTGIpV00c
JnEKko21HyNFb7eb7w5auxmE2slt2A1BzYiplK/KjiC1M3+qBA6miMd22hRrdEaA
O8l9zadHmkRywSS5HBfSYhPeTXuTcccaHAZKeebIxVPEGo6WSkuSbZ/4NW4sWbhm
ctcA7jy9KeeNOd0nTMDb1XlShd0pW1ajhz8RnwiNt/FSfJkDpMbOwO+vZwayBu6v
RuyJ4MSZnyBYBR5T+1lYuKqGNpG1Zpv+Qp2PKRIXD19m5fqpkc9fyYxH0be5YvmV
u+4kvN00BGiCEqBozyccIFHIM05yA8h3lBJG9XSfscmL7/god2u0Mu2Zox3PFk66
hm7l47hM6lSyQW6QLo7AJYF8gLX75OPV9mI+P5YQl+iShRgAcwv0YxOBbIvve/BO
Ah2wrenZTe6saVrNSTqwdt8LTxvvf+IB2Wdi6iQ5GX+pg+IPBJVsINutNy6rJJkv
TBKRllMlWLDSfBxjLqJXzg==
`protect END_PROTECTED
