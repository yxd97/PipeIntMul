`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZQoTFubhLn6KqVhtL/3YwH64Lh1VeOiOfdoH2Rc4kUiNP3PftfR/ww4eNwpDLLwR
SdNWvKkzM7/knJvdesaSsx903EMdJ2sJreeLgfooCTRQ8g7ocDskG5tW9Qc/Bupn
3J+wbaLnjPsdJDZpGi3vygoG9zgcvtOrl7SR+i/1l2BQOxIIKTcr5xwxgRpSsqX3
q5ei9wSXpZNLSexwBYG0kC8jBpK80bgHJtJsX1A7UxuWOz+HDS5om9QqEbFvKYqZ
idOIcfER+dw/qQuHoeae0mhMS/GvfsknPg7TDyZiTfBOK6+FmGDU+OBIQibprneG
ML1kkcBqFmai3Q1h+7LYUCj+uKN5VS24TLuFCfNCz5QQe3Oll9w6RfDM6YbjFUk1
fst5/WDNnFFsLWXQK78/mpswx0Q4vjyjKNVEBF/ElhDQcb5HZkFPCQXrlJnc65/p
DXvPzWHMBdgPG60f8UzCMArhepwHBjwKNIR2r9jXtR9zOuPdOqjLwAPjnDvyY7o7
svXXPWMT0cIp/tnmVROTdgwqvTDTXDKqJmJ8kvvDRMX7LED9QoyBzuE4QKvYdMr9
h9Yg7VPovQDLGm/395gpP3WSZ/tnsyf6UzrRHdfOwS+0nJqLQDSuPfx8yp0ejXa+
o6jz0QuXDtDik2qhNnnZolNccMfKtnTLntK3ZvX6Xy276YBfmP0lRneSHMshFHpE
EM2pJU1CGnF89vVsvRuQZ7zLFo111EogGa16QeslWsTKj43DPaIoyM+rKLHT5Ucw
a+bxSiKUPXjdfAuSXoxblXwIkufpAkI03V99jhd1R3ozwMIO8Or9uAa+R7QemfBu
5tVsWTojZ80AzLumFQNSeSpM0MhSFfMqq8glyA4rlzlfdsg6VeDFkt09QHXXn5c8
FRH3eo49096h9b3og4BRug8iXTdQOUuDEvZgJ/JcLfx16RSdKeF3Yz//ao27tViw
8XsY140i3nc6tEzAwh19RJn1fRB+0YtEKiJs7Q//zlbzOo3XkaUL1QO1CcOW+2C0
1+rfUR0yRvuYUl5/Uu3Q7YjhccFSxcFJvtrrtfFz1hWXVAhlf6P+CfacdtwR4F1z
9egA3VP1MilAvZvQiqGbzP3ZwuDs5yBVdvOnQCLms7mTnQStiWlcQbmIgHIsVhyt
XM111K7TxUIGGVPkBFxqt7JvppB6N0R4BZuR661WH2qjQdRn6g0U9DgIZWGwL6K5
isLCFAdRkjK+LBQFZvB3KBTTUpKNqzSWsNyHEY+MOmOSg+vUVo5+fC0GTs7RwT1Y
m+6TIFHX0THKqozygAUwVovuITPouaJVAYEMQ8rxtFYErKxJP3EKJP1BMWuIFpwn
DBBrc00GLezAgvSIvuwjH7b+dRd7KZlSmpXz2O6VWhaLXf6ejsaEBFYzyhJZZoX/
orga/yxg2l1P0AbdhBFEKhgA0QDPsMH8LITJHUWLXOhFSJGnZ6yeqWf5y1XkvLzG
u34n4+f2aktbSU6QGcl75UGtu0WMYp8XRgz1iN2CqZ3utvWbo5+8X+fYvBNHesLv
bR+zYG3kxrpUHsDXf+yeWd5mVJXiNs+aEdXJE4AAXoeSpU68UOfQ892nC67RfES3
IH1MTSQ7FoEStDWGXL7zql3WL+e6oioZjH0oaEdVM9AOPkwfdvxcK7hsnI4yAwQf
DjQIsWVYCONLlc1x9ELIShxjZ5blDEuuKHWN9ONoU5RpKGOgMKYCIRVgQHAho2aO
e2WvJ+ZXqxKnUnEbA8qm/whoH1ztPUjkEkxS0suJrxLBpqMVkYoafDlFvfoTfoz+
1S6M0NrZNsV4n5qO6gvKx08uL8a3tGHNdakFIHMZcfZIKspzc6gCLW3gSo97Fsvo
oNrw9aSP+xLuESoQjJawbrsz+yY+l3zzP+eAbgMvbn5KAjG7nBCN6BokQx+qoJQs
`protect END_PROTECTED
