`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7YPVaSRTOhDHv1f61x5rUAV0LyMGBOs+5FjH45GQkXqXwoCumHGXzY8O4ofbe4An
uDipKD20k3eg4Lj8QraOr470C52cJNgAOGQ+4oM8CPKrVU8guzECxbgErD+Le3bQ
RnZkpI8RfupZh5zwCk8IR7lIq299lnd3VIiSOF9skyw839XYKZCZp3BwjJQUqTMZ
SvPpoYcQmCck65twrhme6Q1k1YHan2chQg0a+taABVPcHl/zMVqQAS1FcKbwlWnk
1iOKleqCLMGUBiWqoPm/pcEbGMXfRSfy0+ZrLovH/zA=
`protect END_PROTECTED
