`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oaDXaX00/MZd/XGdZqjD1ZMdJivWbzw8+ghpiMH0Zm9ZzGBfuBw2/urlvTgQf8rh
W/9Z57GIDu9nC/P1o72YqIT2IaudYt0otf0ySoP6VWkeBNzQ/L7hl9qkDP7cgm7d
VgyXS7UMBoQ1wyZ1v9reGNJXHMUpYJ8aLqxa67jgBst9cjO+q0Tp3l1bd8r2NDxV
YSmVfm47dBsqCZj77yl892KiNAnap8ux7xGbXu3OnCIFPqgndPCOGXRoPgcKIho/
39AP7o3f/FunyreVO4WpHh0lH5LOMYQZFXi7tYl8aSIl6yfgqPHw1+fB8I1TFaIm
B2LMnOrG7o+VtEAsma84hPgJk3Fo4s8mhkKW8nihgeEb8dhNbW2zEIBtGqHOocon
Zphgwak73wsMGrIhIqmbgQ==
`protect END_PROTECTED
