`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LlKHBGe1g8/DhghRdUev/OjgVY/+LHbMfS0j/2vcugVM2P2rSVSacvRtBKI4FPgk
ucvtmGdY57txuINhB7inmxDF5RpcaY20bV/IIar3M3yY5SK9wccRrNg38eNuJ3fC
/ovyuNx7iA0EtY75OL1/O+NuteilwTy/s7nRfQ5zffIrmtgegyhONZQfcJFG/uWn
E0d7EAMuNJ58MqVyR/6fJxkmp71IpgOahemtRPCRl+CI/pSQv6hnUTGWXGDo03Hi
rnGuOr0lo60kfKaGpaSVT1Hzpw+fmTadl/n2vvtv528qn9rX2QwnIn6AqZk10Tfo
0JmMcutNBIjfoVyU1+Cp4/xikIp3QyDBpacBzxNEa6u5D9XNnrVz/qvNBDufK/mj
utPjXbAXblX2mZbPmDR0uvoZVXwXXAZaZQmpOBCgNDj/yoLiU4L1UbstZ0sB4mkv
WflPfkkrrU+qlNfxeMfFLCBIq731lzN9DqFr97b9LSABKkRqPDexSgiQTKYEajGV
4fZbf4SJ1DtlqhG7BmAMdmg2T3sok7F20xZAoJurWOkyO52gyDJXXfJw5r+3Rd93
9nLzgKw28AJS2rDzMVsJeOxCDeRrQPQhn3jkSGiBUyBeVENvlRMpzhRU+RJ9ICZP
Fi4Udy7EKsz/keSj5uIi+ZH7TzNT+ampn8eby+Q+5QnKGEkGoCUwzZgcT7Fo2my8
5Y7Do1tf0X1xW6NYv/MNpNraXfkRGEKYTx72qhrTPaWCn8U8cHonT56PV8k+Rhyq
Mv5pSSzLrBqhbhgdyRxgvPK4QF1eK6ifC17//vvab4yjagbCs85rsfruba6K8sWI
URfjqWAwhi81BZJXE4E/ncAgXCRwIUPDpoCxCa56+cVfqK3U1TJ8Dz0dnKXwL0O9
1VZRRyALpEw4dTeHPXMeXBc6lrBt1Fw+ou7cSNBVlXoy2uRr62inRlAEdb7oxIW1
uGrD4k8lnAFJIjn16q4W9e6p63HjivNcraUgYiCpceAIvC3pqgoHGm7aeWmPYbjF
tc5pAt9Z4k6WeivZho8t6M6+A6Nu+UPOb9h7pWpKvh394eK8A/2nqUpOhS7hKAWY
5kAetdF3TgrcWnUyV7ulm/Et3ubCHNQRqcViUqgaK/pqXSHvlYlg/UTSo6DRzLMb
lbj7lVJa8ljrJ+MYi8DfiF7wC8GYm2QeRzPr5GyEsQWXfmYuLs8i/xtuIHY3xKrx
TKxbWKSvWs8ZHb5eAZM5sWihx2yWXhtwIm9Kq/MEBKVX99itfVLX45v0vt453aWE
E7RswDaCJGs/kYpQoL7Zu5yzDGLVOt9x0xUjDCq4fpbL3YX58bswKuMBpO7yFciM
u7ByEmXX9doJi3mc3rRca0BqYGqxF9HtTxtqSREdlRrkyNgVSriZsk56VKmwGOyM
lb8wmv8KVMB1/m2pRG1M4i7hXAlmvEhADXdsg8ukhKMI0H8CZ3h6cDvkpmvxqJHR
YVvDZHstbkxLKzGlJ5TJl9UTpNHMjX8/L+LOUFvWLX2eVIunxGH7I+agfpMJBG3a
svsf70gn8WNZzbX0E7SQO1HHdpPFha59gakMQ1fmD6FkhaWmsGRCV9Xg5aECUvLv
Q6aW1aEXIKzV/rKbqZkiEcnjyhGDHDo4LB3uapm7wCEdCsU3vwU2ybaLkgIEFs85
cB9plW4huo1MKiugGDQWhLGyTN4uaaMBkxD8Ch2Ms25oOPw2aXM82qxvScEACeWv
UgWHsl1f0QW6d9YoSx5B722mK54nh3qTTCH5QQYGbZ5S++vzZhYrsCemPG2u2Qgm
f7y1E10SMBOFvWeGQwHNgXIdwVLjDLvlT72MzYwq1/9fV3Fg5G3+UU8dHqwhAXBI
LPD2AgBXLa7vSiDIjUrpxq6u14ujx9o5dHjPnPcS1dupkNT0Cs9Kg6VOJXogKbGd
V0eyc6r12Nm11yr2uAdi+yQYBXFHYElzpJmHAfWtRsTHwYYI6x5aFmw4raK64JP8
xW1FMyE89Fe1WNw8vJJz6pNWncE928tQ8iGqSjrbJF/XehNX7OgKwV94i4NibYSZ
moqYtn0Tlmu5Yh/CNMdxSH2a/Iibf4olA7ow7PmN+7OwOr0oZPV45kwE/K3tgx3D
imz742qlukBkAcLxCPK2MjkIiWCrrfuYGcjiUxx6U1+7FpdwlklnXavPN4fcYoY3
vqNzhL4kbA4uPUjsMj3vBxahNFXzDnC2dAyoVK0KeBnw6i0+TNooesSwwYsxLlkT
yV6D1cT5BbbmRmEK8ASBv/X6r4GN8D8j00gpPtHrj0lzeWmpWAOpPWwcicTgNS/m
5HoNEPDQ3T34u7ODwx/B2i1RP5BGdwjB11orilNuRsU20WkmioSQ4o7Z8hrCQh4N
9L/24MZyyB6jzf7BJARXb3EXb27Qth5UKtjrEQSGC0IWezonC/crpLyuIAhWjUa/
wUGSspTu+B6Dt2R6YnJJEze0zXP77LEMZal8zFtS29+8he320E1aRn6aIOl0ylEZ
kvBOhaplSRNbiZaaSkGIi7SYRD2Oj8IfuqI9PfZMCDnV2oqTYxoFT3Mh2Jq3PZIg
FddJ33DWIcm589fUqeDTUn1T3RlOXMbZioWXgaUtr6RpOJQWQ3rEglYNiHSV58W0
tf8RlnIdb1pFu8MSU77njLIErtq981qzX2xbF7+IhfYB9jrys1W58OZ6I4vZwIBI
a4TcGPkt4HI6hXzfxlhgfr43F20GGetd9wafCsD2GPpzTZUPcGJgaOWXDWLLV2ub
C/7aLg07sJhkKpcuV8ETWtP/PyU+9/4jrEeVT4lQFY2Oo1PrNSJdlzZjOX73AC1A
Ebxwr2em1y3dC01xkkKfjewUt7xA/ztjVw/pg1fePYOwe0K18Cf40GDOBc3xWh4/
GtmriU/VvJXck5/VLEzgb96NfdBo5LlIhIlFM4zTg/8xIpmP5+1FId0p4F8dTcgz
2ytXOKjtIeSBCvDgFITjbwG/+jw+uMQk4Z6Bv3dM1QY85Waq8DsL1/1Es8PC4nBy
T02cIuV4LHZivmh9LIu2mwk3nfE0MaLusvsadbWSSXu2ofdaIQG+d7o0i51RsH9m
LdMdf+Nhq1Ua55MW0ONXUQqFOuHOnZwWNRwEGufbVJ3jobBphzNl9fD8VpaGxS6n
6H50bwTCFCFqZHuQqWENko2G5kIs735W1Y88wlTOJrM9PcBp1Fd5BdSf+5BmY8/y
vX+C/5a9rF3CI65Z6FT/5Inie/blR7wwcVvX0H8ILaedBzOW7GEjpvrOo4tl+ALW
ewsGxp8Y1/KaH91WY7K6U8BYbqJvYnR2/u3OJsGRHKo018gDpK3eUxfTIamVkB/A
lUuNy0NYRGCIUstOHTnuMA==
`protect END_PROTECTED
