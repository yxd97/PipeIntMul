`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xAg46DZTTCaD51B9lj2WlAWJmvUYam7vMFpHQ/ID2U2bEFg6MzsqqvH+oH/JmCAK
JpBX5qgI6paGlgaZv/evmwfaFSJ6+mswi+/dU/MMLUoCuHzAXHaOBWXUx8HB1xMm
Ad0LxgU6UPraHKSz/kMkBQkPH+kxKRg7ni+fDJe1+gAW2FoROZYKecNLIBTVgwib
5EkmMzIe0ms/JXp53StLtqKpSSXbYO9IG8UX/paGgCcsbOeNIkjJ+g+rm36bM5Ev
YOnNx7hH3VObxWSFyeV2LuKBozLnnlWpgVj9UJhKRQKnOV5qbPlrk3t5oX8wMZ8j
KotUJNMTEuzcT3JKcli/t14uxbGQirhjor3bvE9bC65jjlWxs3EK0fQwwAyYY2hu
dJ3Nm6n6B4deg6ZplDV1G2rHyfuJkZjSKAqiG9XKFK0qE9x3Nv8/HVfmWd+MRU/H
IPHrKigPm9PUi36f6sDzSxWrLNfH9RdXysW9yYDoCPpGwDFP7q7VTtfedOWRb5ct
e2Ytd14kVGMcYdPlwW73JS7xXxa8l5wBr1w6+wWQdivsCJZh6L4pvmC5WfirOdg9
nV8r2U4Q/pQFZfxHka+RSO5oYYAB0FUzQHD7jfGBTddwkQa7OHKGICOeX+8jdQpH
SNL9bLvB2tTxSwqApipe55nDV89eUOYqWDyVZYcLHtkwSZqrN8Lgfc46/nkW96KZ
RYV1fT9FGEvGCfihI2niy/VK5g5c7mdQ5zXuyCDSQ4wwon6i2yEu5Z1Sz/VlF9Ai
0T2tcu9GMAercNIaEc6Z6oLngGuLOZaTY1Chx9BU3SODVF5a38LMaZOoDJL9xRW7
1dVzfADI2lUTmb6HCqsmszEZaP3yQHclbBQfj0hnryeyHxQW5+DUtSm0lo0VeKv6
Izsnf/7ZiBYZUuYOKa1b0gBlL4YIjmn5k7OeW4NUayZ7BYpfEAbhlSBZgP2B5t0K
1xa576M1Phw26J+fgjYepmSCqIonby9V0agDPfwi9C+lKqPWH0CimwzoatDzxD7R
1mBARej7wANq0d4iQpDR7DgeFfJcTdA6G9SXYkqOPYOM73IXS6pcjpKomyVAkIQF
A6P3gQ2Ve/lORszVUVsgOanxJ7YRX85PlPfQ05oohCL1dxy90oKzacoYusZirt2l
Mz2dm8szArI7ftyx05Sog8xULS9knorPh3EwjwFCWdaMU8+Td8v/PQWhfAeJA342
BgkKYpGmTSkRgUEnvdmVHXKS6/2V46yuKJoIn6xMQ5iH1sbJT8+mBlp83lEeF+Oe
xDOPK6Bh2ym/Cp4ITdrkvaOZGsRUkUNm+GK80zbemr7+b9XWH9uBy+1vWw6/kpDv
2uiveubEVeNtjM0puLbiL18oWhTAgwv9Vz1rM2KNEiacr/HJu1TDrd4lCormdLzP
ZSowYGJSzC+oKq2WNjhWEcOEeqNnXHXQ3JmLh+IynDuOaEPanrzHzYGC2Qh8HlfD
KdjLZ14Y2WmrSNbd4dKkLysLtcNxENo2xOYmxIUF44s=
`protect END_PROTECTED
