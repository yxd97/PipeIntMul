`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0Jp2P5Ffjef5rS8YXIi91wXCzzha8ZVFh/N3B4dUr2i8C2KCUU9fvRQwxkJh6pJ
CK762d9azks9DoPy74SfgGg65U62t6Lj0XDLiGF4tzJXcLag8/ylX12dS1Kzofrr
yLlxatk0VGEDY5+sNEkM4/KUx35yEjOM9qYANxjOXv2fRW9gV5Kxhpj1s4wNE+4Z
4/B22moFuA2ir4rxJIwGdkGWqTG1AelTB9hnMPjq9qqntjN9Zd9tUwp6yrK7KmXB
HPF68PYnUR0QZnjLMMNuZRb1nUUwZwcB4MX/eWysncEJ7za7KKkdVn6i0czIajRP
euTIemprqMnEsl4n5mRIKQ==
`protect END_PROTECTED
