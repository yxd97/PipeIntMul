`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zS6IIZQRLQkQSUzUVJTIf7D46FlAO7SALcM7QFKt8oZqlJUN4sZ0lO59eLgLyZBT
cik76meYMdQVlg0KOOwyhzpIYzKwFcklVnS0IrSGDRM9qmHZV0OWZv5nGQj+53c+
stIags2FCxKzuRRUot/9POff4EqKFxOpnJ572HxuzNtBLJCk8Msq0EG74In8GM74
85KXD+lXLTLk/OCAb3ElqnUTc1Z+awk1V8J4oTwShkCQbKsepo6L4Wsd4izrQtoC
2CSptUX86jlrJy+OMhmx+HRq/nJzFNGVD1J+a1EDjA7ZjzrnvFa7JS5Ns/zgMAsJ
PxRNNvnJf1zcdsEQ50ib5WPQOtXKillXaWt/D+S7faNveTMeYwdTcXWfISWP1Hz4
haVzuZyYXlwLvcY+CM1m1Rof4V6i+RyYNI87ufg6xDU6/pU5aOcp6rRLy26DPN9z
V9f49xHiJyW/iALsbSBu1deoe1jjWaVbowhGDGC7QTEju41rBGCjSgdZFu5pTCuB
PQVu7J+CVzEhoHJAJ4hnoPCN87bYYSh5czukLnuHUEDKw2u2MfSTySMyTZojje6C
CCXJKhiABFd00xMk3qNkO3YX+M/J20BqHfZtcCvrVmmDx34eem280eIpyq14QOFP
MgYgA3cPv54Gbm0FJni2jw==
`protect END_PROTECTED
