`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VxGDWMM7FMh6oqAo4zdxLR4F0IIS8YD+79l0Ewbp7A47T3kUExOQ4Ygbn+KCW8bb
WzxknyLI7T7l1clTbH0RZK8bLkU44mNOWLutAtnae0dcIzZjEfoKvEaj/UmETr5c
oQJD0pUEe+w1BOj6dRjU3/ZefFWFXzUIMhbTW2jKI3tfXGlFvSLXYcKxiwj6a/he
J2fch8rHIK9IgjE3XQTLfVYKfUWoz5gz+Wz52j0sProY9OXP/1i5zuBRDF7Al/ou
DSzbwnLvIGSLhbCMu5KfBB7uLiZgjyOVE1iyTw+5a10=
`protect END_PROTECTED
