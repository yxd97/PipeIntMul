`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hps6W68iWYW39i1GdHClhEGvQVgLsWAv+6sLc+WQLvd2pdrsQ4lT8PZw7cIpI6sE
zEmJCIPMczkqPZztftZXSpKoJ3SjwF7IdzNMVRlxhxv6SEwDMv1R2VQBupnHKi80
OlrpzR006qnbn5Y8Beb6+ANgOq020vD8PiLQs4mIE9baofPHL8Xg56erv4xlOiD5
3vQzTKcGrtzK+9mmsNfscBrb9esd2k1ePOiIiZknirH/q/+Yi6u3i7luXMenfTig
e/YkNdSVDZF8E5Ke7w34FfK2EkfPWCW9tixm182YvxTz7D5lHcZ5dOm4hqm2aI9Z
6+1w8gHFI/7vOyjtWAlgyqttzna/9be8MEpa9GEFisFexEJlLBkf6StjVIsKKty5
5ryvN98ET2BcaxziH86yrb0Un3++sB22YbnufARMvG1pzPZaN18+HY5BHL0FpVlC
mbVXed5dY7sq2oH2U0JIl+bPA2vDEPJWjrO/Y+ITaphUIdGW8DRxPyubZ2YcNkVn
`protect END_PROTECTED
