`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
91Bj8DujiY0UdgGJTmMK5PUJk6pqdHeItdcrCR3bzCD2wYkQptjholavTj22qxOy
Uy5LunStWPcMEauXbYrQoP2s8jlyiRiBZVdLRT8vrSaHAV23EF+kyg4BGO0A8cK8
JRd/OGmmk0He1vcfozR3gXfeqM4BDUZwtsjtiiaIRR3X2jEXhrNuHn1z6b4xydry
9NnPPBvCJOhwbswWK+wIPE+15I3qRSN6edDY+MOEhaka0R/boRV3neQQgyUWHDKH
CDYmMdbVFKqLzk0V28yIXM9y/bn4gmFY9BfttKNAqwXAb/yEc5NPf8taG2plSq+y
+xe9gECh1ydFyy3vqzM6LBeRLC+ynKLVqWSWAkMmQCIJGle9XPpK8ioDUJOESn7e
OQ9UfRWf5XT7hWM5NbBYLrN9VX2WORGOnPMe7wpT5WxVVTk35gZWt+qhx+/Cmi0l
H4rZ49nzUwr7idj5SLbXZRiayffWHISMoFrPuOcrfAnebFAKpMonEXOwU21BFjBA
uHTMaYDt1EEIsN6s4DWDk8FGN2+ud6+THDDBE3zqGGfJR94YwZ961FELngXzu9+M
Kn2tK+YBaPwdh+INSUD+K9khBzK+xmDUaIQ1k+aUOJE=
`protect END_PROTECTED
