`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RFucSNmTABEebpUjiLYa8lQx0O3Ekvnl5TFvzRWCNXI/8YyTlypuorQwGtfxN00O
VYCn7lrSJIHmaM0U8RE2Oa+VFJapBBbgE8uPJE968zW6O17+0TT8E1/WfzpENSEM
Sy8gg0hmASSQK5V3xdJFDvRE3hHI+w3NcuPGymP+/AaP7DJkvH4nBE9JUw0hjsvk
pNQK77fvCymaKZXewW+TS54lJ/eoAM5ej1EJvYEMMPjVTX58bUkm7+9hM9B5jgsg
TiLHSMTYOAk9k6IUDbHE17KT7wwa+n2eu0I313m53oSbLOdgWxTD0l/vzTXlOn03
DpxLCqyVlZ6pbF7wydK+wMN8/Qxfa68dO4iepcjt1kNXhf9t6u5OS9EivhWyzAYY
S/RzGzbLQJccFW/aJGmCKnnVJsgg7pfdpIe9PL69Lg05cLlh2Bsg9CyNZ/oj6FsI
r/2+vPlpvMNMIivcLwa1MoP03K4mZI1765l4e3EuwylkWYvwbWfKZAyPBzIAo94/
0A6vIf1wi1Ks4NHJiO/GUjF0YejSsWosPrJsgCKre52lqq+64O9QfxYk9x7e07Zl
8PwQWQV7qcd3DnLqBkHdjvmDq197dZx9uDi/bRwOzxAcqD3ADACYTCBrTe43mX41
dy4ZA0MzZ51vTKVDLTkhQywe7wox3/hTVC0eC9djILXy+PnWT2mSFUNVmXQ5FKCW
Tt/IvYzGxn0CIHWAvRwzUghWJeEJuT+AxOEEpVycAR6WVkrAGzisyHx2ZE2qqA3Q
DNH2TOWjTv4C6TkVIySK3hAgtzFK42x4poed1167P/g9S78V224JfkHX/659xVNA
7jXbETiZKHPpTlDHTCXA+XbP4p3G/bmSTh4KUrfE2VIH7fLKd7FO6Hg5pkva020m
3OsimVtL8NMOax+aNwpH9wgqbLNwN+jT821uId9uWLQ=
`protect END_PROTECTED
