`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lu6NGmepbdS3BhZa3RTrd2sG/03Vm07HO1YvBnbiJwukK2m1Mb+vjQxKxU1amNpq
9zbLDVziDRnKiltmtLs1hpUCrzYEpRmrqwj2wNerYlVlLyuYu8+czj68OL3tkyIn
lv4Nprkz9WZSDmWl1ENOAaKjhmC4xEbU4LDm+49C40dH4jaaaqmti0EugP5V8n0B
/nEufLmUtBOMK2rz3qVT3laG8hGeSDqehAdV8HbnGLIH+8R940nX79d77HvYbceR
1lF/abqE5Mkc8ZBVKB0kqhPzKDCBoRevOY9kpj1mhN5GJNHH53j4grMGdIisIcqC
NJzfiaqC3Ai2IRlfh2t3iGnyynlSIPqiZOLCa2Yr7taZjowSFwlZDXqyZwe9UlQr
UfKHch6+86lu9GTjd1OsHZ/KgwgKCzj0eEFl83MpK/WEsJNLHRZP4MFUjWbmNVUJ
UwqGZc8niYSnAuJGFPPZ8nQqAw09/NmNdwYfRRFu7UI=
`protect END_PROTECTED
