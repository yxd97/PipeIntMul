`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jWNOntGHb7JVmB9ntFav8mMJRY7yoH0pbABS7DQ7BomKzeDiDTkYV9MXrH6jGVEW
kmDgNTOCvQHGPz+QEQGjof3J90Ney7CTIIG5uEgKpD+3O25JjRmT8rmIUB8AP5UG
H7WxcmjZTwBKLlCZZEvI81iGwopo7NHIRLAIiyLNBE373bRok5zs2Qz5CrfdY5iS
Bcj9gaC0BJCYhqm15cHFv10uqU+pTo5Cd4BR8+t/w+H9+zEui0Sadw7fILTGjNAW
TnDA1mIARH851LGIzASXHNlXhn3CviEjOVaOuMyAfx02Y08IwBpa7K5UyHMcGwud
M0tqCmjk81GhRWwUPmVo29Pevb9d7eqfZNv23e8VteRoDmLxFc5Ro43dqJRv7AnI
5k28ra6UUWsYDUdnFU0sZg==
`protect END_PROTECTED
