`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x+9Kj6yezRJz69MUSOQeLL2d7FIejbilWTZpovq1Qyt4FTn7GLWnRlrk3O4ShipZ
kbV3I1pZbr6l1ukvETL2/v1DGmLO2gH+VaUpitDtKalk3bIatlkLjAorTFaHTqGb
PX12781DhWf6ZW/BCl4g0Um8CyoS4Um61wj8WQRTFTOCFppMmTB/xQvYcZNpX3x9
cYJ6NkN1Cft4+pfarvqqn4e0w5YoBfQsLEjM3mBOmW9lznEq+jjHqgijGHEKoxbE
VYeQ2vobn5cxs+NBVxKmhc6EhroFcpCXcamP7YQR6bqrMETutxKdnpUGXGfMkY6L
/fbolUDOsSdVpw/1xpC8w53DOPlS4jdWuoJBB+a+QaJNgPMOvYJbP2u9CcLOq/Du
BycRGg39z3SFeM2TrxeSyCjdbrJjKbetXPE4qWESupe3Dn47XGvX9UXBeOXpgtXs
HI+vjfQ1CcTMWgvqKaTdbHVb8Gk3BpflDtmVM2mnLF/4xOXV8PXJjgmMcBXmmMLX
a1prb5lkggOpTPJ5M/a3x85XR6H+knDg1zWy/k/JG1c0Yv11sv0eKxTYi4vohYhr
bSYGWZX8xf6mlJOAiZ4vb8jhVkrkZY/f7uAuMhTDyo8=
`protect END_PROTECTED
