`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5mHm9i0wYzbbJluW8MKY2gFpW2v7x+gRNnnRS0DYyIj1LVs8984Ia8L3AYtSb6NC
+XNRnu9YTuPHivHCpyXJJePGVqMKNarlkAcQ9IS7SWoPlDH4kNhqf+Iuara5tHrG
+0wRY3Ff/Nr8K0jhg6vC3Isrdxr9zDnUamV4hc+mv3r1uG2uaGXsQF/TU1Jnqnrg
lyQ6w6CY5vBPKRpY+FpuHzIf28azSYCBsuF5ThSb4up61xTGaGXglCzXyS0qeBAC
XRvyikz4yJ59TPdxPQdkUV1YFxemBkwrHwfTm+DzIgRneMablWEfbXlU50aJJT+j
DOEEgDRTNgLB40dX5aynis3AkqWj9Tcqqg5dwgq2jaQG/x0CpZf/7/33UrSWNjCq
kKcajyOlOs2QTUprqZVLiIZn7iurxAzCwy9Zq1YcdzUoWVDjgDppZRUCR4LiT3KC
maMIpRfJKNYb74ZAC4wSY9vN5Hg2kDDGVs2hVRHsZo2AeiHxWhNdZ3vnutAbkY4k
w99kENiq77HdKIivkWnrT0Q/RBbgXUKN5U3vNCpDCnn+i//P+ij0HRUAwjir2Gq9
pi+O/VpG2HqsifoANUWTIOtC/0qqBLPXprv1sv2ZYJ8CtTrR3//yrbJZqKcUb6Au
vXkSi/rU7vqif4K+L1gHqaAfFc52pS3VrvZ2iPgG68fCqgjM1+3PcNJTKzfwq14d
sDMrGvWaiq95kaAZMqbHW2aIkIoBP/XjVqdcFLyLtbNgC2FjQ7OCmY3DFWviJfek
MW5rCmYHJaXoE34CGfKMSSnE6UCHNqX+UJUJRBL6VIP18B82UwL7lUEpcaN4+Dg2
rg58XGTCUJprHqs+cNKMQlIZtZrwZ5mQ3xwHCw9rk/yhlssX8x6ocLvsHR3MS99o
kaePmfNR7ghpBs17ud3YqxFs8P0kPKAqAaiyq7VYK+8zvJHnywk8vIave52KY7Zp
+k9tdTV7ypxlYnW+vDWILOkCSdgpubflfaN0uVrs9q0=
`protect END_PROTECTED
