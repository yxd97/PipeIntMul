`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zbyVe67YcrJHcXBTwRhkR9BtWNJIXak6KO0MEQkSYN2Vjs+LpowPqEuCzV/QXLy0
0rdfMkeso8Pp3wSVZ9w6KUpnMLV/aBROGWtcf+EFVwXHhy3QFxNvQiEui78MihEJ
UT2iS+PcCAgOq/QsP1fr93U1aI56coBiX08D+aKWOFcEosKkFjfjjdiJFqgGnmZp
HWA/OiqlINsskR477oG7VX9a90ZvcwGhIDL97fONqFXNnk/on2GQya38v+SaY19/
+DD+J+jCSYzuxcJ0apnx2P6d2hC1U8S40yzAd325m5FZNbt5UXCSVP6HyPKSarDp
4RfjTPeJzmgbnzOsTCOX0B9Zai4RPL6xMMecibI4pc/tj3PI/vp6IvM5vhhWIVnz
TRn/Tbtl1BgWAL0KQ3Su9mpSwcv2WYuJDzSV8jxHesU=
`protect END_PROTECTED
