`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
il3uPV60puLnVDyD3tWT9TNWf/HUuJCGD3iTnNawOS69eJx5YC8RYwX0GfXM+HOf
exce8a+96t2AXi1PmDdmzkLOV5K5AkXsbpbf1Jnbcd+s5GDWADhoSzROXA5dUj32
oqqm6M98yqJ4EUuspAUpjVZfv62GUEkOcDObo5ZZN7Bs2KWGfB27meULFRtPSRDv
uqgUCTM1sUW/01ZKSoWxnQS4BO98sNGksGNdtOZwdIbDHUl3KSPLeFgTcfuYk6OE
uaKLqJayiQRl7aoWZ5cR6BJCw7NtwP5Ki+vTo/5qz2yrJoRxXr38r2cBbiKkL8dE
DfJvJcYOb7GesBMqIJDn9fvnZbao2XfsfdRy9UsoS6mO53S+YHM5EKinEckXMob/
KSUsRDUo6flI5W0Fp7eATsRJrSGazr8mi/YxsrXjfNizrtQ8TxIJiEcStEHhbPu/
nHglPC1C5eBVfPiAY3WklA==
`protect END_PROTECTED
