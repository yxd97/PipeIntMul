`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hox97N54bOmgpt6W3hl2lG0tnchQhYaLtDf5nubxpvjaLF4lOyFzocgB1NSCQEAo
LvSRE8+rmeiiwR80Cng7L992avuYwkuUTtAOTj+11wE1xLfgzLmytGkFvTMXxv5i
ps5AYh/SGdi2HRB1zmWcFkl7c7xxhIMSHcsrZ/ZnceonFSXTBEV/AZ6FZauq2hTX
mYbygq3xuwNocIfpjTQJM8HjC1aVHhhuKw9HRNazFfzRu3P1BBI5UA5mLUDAw9MF
8U1JE2LpqbvAnXZrKjrcVeGYqUc8qNm1f131m0KXNeMM3hcCLiLreiiQH5ax0ffW
CJ5etNFloc6h56j+cypjoOHfR1vhpsH+3vh11J4UBF4J/0cBc1VHp5HXbEtoMnWt
ckq1//WsmIHYGBHDRde6Bjz51UyiJz87SXdWuEUFl5AnS6pFjyK5r3L2ps3Rr6Cy
Q5hrBnA2Nj6/oV1cmXvcSr5QAoS0Mtj/8qeZpn6UcUvYraJr7U6gcFqa546j3RG3
03jxKZDWCVlIr0NKTd8atcSsiEBbUiytup93ujb/Ps0+kuPyDT/SFPPasAZotLFv
AVxi2+Gu4GXV68XZBrrhhNx4qgRqn1z4/JlEVp0SFF+WJZwpqYE7jz9vIl6gd79D
9Kl3tMu8segvF176wzejKiYc5/AUcaiMdaO3o78Fj4yuXa1/OAhhCN/P4oKMS6QX
c8cAq3EVb7Q8PH8JInx7ufMnpOdLFF7QDvq6w07fdadQKBxrPME3SYybj6H13D+d
lR/empO5aOR35lj6I6Hbx5lJy1xPn59/Fd1cIJhwd1cYeciEsy5JgZy3QRtjI/Xr
RxJlLKi6n0aEUFFLZ4cJa+qI2s248eAzx2U5CeGBll7zEPHIbVlWdK/z6syC3AbF
2V8gHXF3tNTE7xfFfI5awbqH7IUsDf1qu9DtoGgNMYZqj7JDQhoq1qH4XqkXGf4B
5/OE4RgYuFK6W29rcDeMvL8rKVxI8lkhEX76VE0uYHDxG++aa10dFCT2DEuIpq/H
AiGs/kAgrzNbQfwkixnHtFDrSjmFLI06auddLpeWaJHQwFZCQOUyndzjjVbdvK3l
RkcCkDtpORtUg263fk9CUljYCsngRs1erFagkB4YWoX07yEWb5U3/Kog6QLHK/72
M2RVYoZbuG7lpxkY3RibYI5kVjrwXsaOZxo1EExgy77Lcsl/5w4A4BUgGQ/nm9lh
R3yTru7uG52eeK+hUWf3jdExHbxU5ZSE24XDAiMM0MmYLJlyPlwXxDhcv6tI7nZm
ln6SN7zWD8UEzrzvJLFtKQ==
`protect END_PROTECTED
