`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pztuqL1AcDW7VqeuMg7vPc0hSUUbIcSU9+Kz0ivY5fOX+o0Gep25Buh/ybgY93S2
c/GaQPtKYHi8O7vamXXI66OgZ+fp5mHWbyJOsFHuE0ME/jAHSfFjD7FjABp/4Bft
iReUXXSUFJ2S6tiPMmsgpv2YsqdyNKt7kLFdrT9p3BeJhB69RcBU0t3WmV1yISCT
WRBkIMhKt07wKWglJXn1AAeFe20L/SvEVBILcG+U2K/fbwccXvXz/4dyZXmilM8q
YYkhej3QLk+DaciCUQKGCJNHU2/ea6UrqqIFXvw/QW/mBmE788HbLUOT1sD45st7
VyzsiC7KzvpZ829dXAAyoV4/bwK6iywhb03Ed+KD31eIg6ks/z52AWYgCL81cm1h
XrsaCKOOJBswBlM9qTBgelOjJPe7BW3jEDWJgrW2x+6fvAOXRaUvtb24PoWYDRYp
0FKXhuG0M2N9pDNaYCepbh5EC1IGie1jfpLO4RqOHSnMCNcwWVaCQ1xBsxgmYji+
Ona3Hqy90D9oidx7QiPtJzq+Dxv+MZaly1HCYpjxyJsuVOqdgv9Go7rsvJ4Yn5KC
t1MJklq1gUPp3C39wd2lOmhs8baZwVk0twBq8Trt6QYVYU9sQ+WDBiIXkCHFYGsK
ZgIrbtGOATkPtYgBRXmQVmC3ZhH5zg5zRLyPs/kek6smYKTp0yjwfjnCGKSLou2q
`protect END_PROTECTED
