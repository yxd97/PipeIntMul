`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Lmmf8frTch0DwW9sLwmCdQHub6hKVDmNUw1eKk0sCnjHek+TxWRmqsY9QFkqPwFM
F4j/0WKj0xY0rmayQmcjTx1xP8jUKsH/Mg98yiBjjVZzpd6PYSxiuhKUV0bsyIvU
i4kx0nG+I0O8KrBxBp4xpBh2GqPFDF7DNzAGmJ9xMGoRbBztzZSxu4VoWeLjB3yW
d1ZUf2rygnTnSmLHTntV5v8ADsIEoXCvdEHBjtPTpnoRS5/sFDSUQIxcP4+5xQGp
`protect END_PROTECTED
