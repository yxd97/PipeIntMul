`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HHBzeyeFizn3Qw9a7b2M36ngaTUbjhNUoxDdfkWjuqr7TCrxmgZ1T1HnLTPF6CZd
bqiYmZROCYqzVsZ28X05Y5U0z1d+Uz7Mzj8wDrvCduVFXRi6XWgzlTWjpvF8WyWx
SJFTSu7ofQTJkTGCitWuK4o+O969JgEPuYs5iBsDruWoKj2oYDRoeamfQvIIyTdA
X/dnQNvcZLEMaw7YSgzbluUBiTu2WD1thApjQ02w0QVSbywSVOcxTJFEdm6MkQ3j
yehk0H0r2L5hUXBpsUIj1KsphDqNYqhBcls4llXC3RP8EjFg9sIcRmz2LoM50ELL
eL/jO1y9MOpIWlhJ9UElEZRKylujdA9A49D6BUZh0tnBb6ZMzw/QmSOFILl7R5Yn
BtSKmvToOpSTPomH1HUJfAMg8hqf1RhzVtiWtASRTpIvApbU9sIal36qit0ARAED
GfcrTUQi8u0ohIdGwZLKwQekqpcQX9qkobhVYkAol0IRy56YY8GpjrIc1XAEgkEB
WZTPMMw4Lx9NmCqwac4OFYsMHXPI4Nz5RwIUh+s77OjBnRGy4O1RN5zhQSjhOZwS
77XMeGxXtu0B7TQCHBksEip/bMe2hzBVU0OqxGnnIvL10o/ayoG68vfCeGfaqaXm
btRO3SyR/mUhJPQo2e2Ch0xKfqj6szRPYqLw91rKaHwQaaCWLVJlgGdVqYYs0Vx9
n7qtR22ZAXA6M4fsqrm2CVV09cV5JrYOjmd5JM+OnPR2docV7YCydd9SrOMljHCE
F9dZ5BQpuwjCHhbYlBrZskS54t+v7u6n9ODClZZyqYiPzgkiAcusty8tOo4mMHYd
qL6FjTaDeDfCq4GA6TRdl6UkyuYrX/kAe4Qwtrlmv0K7qebGLxeCNUYREDx3wgZ6
J+cpfePOeupSqDhliqYVlK4wZU9feEeJEMke/MTEqXq7QvmrlMUOErXD6p/6zNNV
DL2PFN5yuMxc7kOpn9RHC5/tQYmaF2SiC+hfieuVLoj5PXn3hHyR/ddEdn04CBRu
SsIbElC56t8AIXmSnZobWkQXoh5NoacJx9igem++uging5kzfDJNRQlJ43raBE8j
Q+g/U4wgya9dYVKMALrVW4EUSbgUqteRL4eQnLTY5j4+p51efcFvdNrfTlW4tHlH
24I4UuFnFq/YbGRgV5nyc1lC7yzdVcgJLWmyuF6/2A865S+NdvmrWa7ClPo+oISQ
U80yBNxS+7UJUUf8ZJatXtGQo7VMoWePrA0MC23sl0mah1VdP56RVq3G6KgRmIEF
/+T19irVb8mgovJZFNfXDzJJ17fqZoTQl7ww/BPAHznEexrxri+f1m1SVB9baOkE
UMWG1ifw8rybVtD17n3unqIpgJR8X5eEA/jz0QfwsQjt5Liiu9mnThP77egOD42Z
JCDIEqGYb1jmiKZHaastylvbtjX5eSWi2LOLs1nF+XM0ua1nroV53dEESgjvZYJ1
wnACMMVqV3miaGV3ocgl+VEXsHUdB0slieXSAV/2y4IcOYPkwvLS9wSBXBUvhTeT
`protect END_PROTECTED
