`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UrVmWCZdnNs96ZSJpK4xqPa9ThHxtFbTBFPCA5zM9n/mWb6eEhhPl/9k+EKkZ/dV
X5R3cc7nDtnb/CHI/ASdo3UErzRulJyEMChEwt1lpwtFIYsg7UqZBm+OyhPbrfE4
MTSDeX/PqFCsPnLSWycdO2TQ1vDPuckfcqhuhOYazZjTy2nQ3OJhGU8vOywfM5lM
bq1VCyKi1znzhQy7EdgRewlIa+sGL+iT770w0GSD2gA9VZ0hoE3Yj32it8t8Ih2F
uxOldzuksCI2DdMnCvSNq0BGLYc2hrDLfWce2Umqb8q/0UWWrrRYdcRSBclwqcZB
vjJT1lF/paaFFsTlfkP9jClJLQOg8dHmZ7qMOKnKXEqFTapZ44/kMvf/Dhn1bGK5
9FGsTytB8tf3nvRz2VRaHafmt1KCBkELStwePWxq3qioW7PcM6+ow/h+ssdu1nZM
9b9uC0mRaIH52D7zLBfsu29ifE8KmPq5bxLwqELe+F4=
`protect END_PROTECTED
