`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sak62Tc4bFJFvR3sfbMo/rkNoD8CYP6O5xUoxGLI85FYVvrYMsohOuMwiSIo+as+
YHNEMqsDCsgGT9DfdNLb2KuySbxaYgDFu6VoWdLa6h80dD1SCPkeQdRxxaQSLaaU
is0cCaQ+juoloMN1+W8BWGJtDGXvlifDYY2SGlKSZfe6pBellMmvTnIdK3rZOEu4
Akn/qvEAgDzKJ2AUrB0xkEYkKVvp1vT8kldz0Ysz5Kipl/Mis8fLsRhHYum5J8I4
LDYSO0sQIAyYDuQprC57u7kqqtt4nc5UXXzowtEupBHq4mv7SW2NqidJSn7aRnAq
g+2niXX6PbES3y9VJEYDJbO+EY15vJpD6VMNuUEYxfHBWYeKKWu6RdN9SCxm6dqN
LCyW6v3sDxrtRoQTNcHqSPte22e7KNNpY9Zg15soHiMrpoFgbUstccRFhhLfMN16
EiSTHZUUQXRlEfimS9ldKXr40jO1SG1xlwYDm8fhfwih7iDYabPgv9DsfC6t2fJg
f+Rble5I4pcoYNWFjVi6q6fxhbElb/shllPneRwkio5dcu72Vo9iEi6kMyMD535K
lv7/39OeylybZCljnWaRcjN7srzoJ+sIhiHKl8aC5iE=
`protect END_PROTECTED
