`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfkKlE+1UJb8sxYQRE8cfSZAyaLYHIKzcUr2bQXJpW5uPUJLhTjwOTsSJgNIalmI
KW/8h6W/KR5LManV3yccWi4qvdS9AOJEKR0y6JDyCAEc8Hwrv5H7F1idIYN0P3t2
K5n4qzbjI9F+RZLtXSRef+o2BDHQTw8flR0D+v8IIagXq3EzPpHUhy1HQs4evySu
9luIgfUR+5u1O+Z4rTTPFpUnKycj51Uv49Ipone9ay5iLOE/fPf+oojke/lMjoK9
qWnuMAfrguuV8hvo/2mjBCHYXqgxD+AZJ9FKSUf1K8r11MYPpLu3KivljBAtsUI+
6Kd87p4ouR0l786rsaiSSEaH//5DC0IxBgGR1xHzCa6ZdjdHX9lo09S5rRBEgtv6
xF88IAM/8/5BOkK3/fkto+YsLx9vDKmXOMyPTkCBuZre9F+5HypoHOzEIehplOWM
vzGpDXj9+K3k6ILXjFjlcoFw+zT/6B0xTUGqKaW/iNEosBJQjU067lQ/P0S+g5qv
7GX44pc/XUMVhLnfbCwLvuVi4cBeJhA7z5CHSSPLh2d0ijj1p8hbp5P2JCpjpN2y
4UgSN/2RbsHieke5oYkulVJ700Tmfm/ZOrtLwFCqKDu6A5QW3aPtZCaRW3a8H3BA
ZwJOIOf+WEze/uA7oT9Zjc6CWK8c2tx9GYtPOvEUl+znOA+vf9v6o3Oj5CnyM+JD
DmKs56oncUWFhob2AqtD1D6tFrdqqmYHuQA/JFSKtP6liVjLTfPnpWYZEIa8DAeg
w0Sko6K16Shk2j00Hel4ww==
`protect END_PROTECTED
