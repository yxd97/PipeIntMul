`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W1gwOogm/U+fiVpeFYxnQgMkwvomjhscK6ZfAZpbs9qCsM9FPAz4X/QneVwJpgqX
KoxqvPhmObiIsvezvUYEBZxbF2mnUsL/0h14MjXPioNrwuDITMY1AMwOQ79iEXdj
efYUIbFpqrUcF0pievZNd6Q6/3wdP/HnaypoKQUfdpxGqAReNcCQwq/a5xzY1yzJ
3GsVNWs0a/OFvy/VdZoZCRbRtOPDD3oBRnlnEn534mjP3RaCUhV6zUjRHyXvsZYp
WY185w6D2y/tfKXFPOyDxmdNhWHLtWvPt/sHgYUNBVEeCYwbzQ6oLOENvYWwwXb8
zqsMeQ4SvBj1aeiPydKkxoWD+jmVoOlsyz62y1jSn0UlQezIOalPmrdKOGtrIyxh
n6poKMn4ZbeZdPyuWTJpqA==
`protect END_PROTECTED
