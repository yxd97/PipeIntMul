`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T0Iyiy3+sn2nJQmTLgxs3AxZVnpFyTaqDracaBLadY+KGUd6CYywjMypOxbBeOeM
M74MlwgypkwJtE86Jl2nAGaUGIgLKINY+DHdfDE4PuHtKTs4nk8O7MMU/dJ2tPyq
+B5/DbqIhnQz4Ck+wl9AyGDzaydyCAgp2kZFcaqrCwt6q87neKqZjUb3D+cZQp2s
r4L7uCOH4qTgmEgUKQj5fH2i3JD6qXwsqD/UcyqDnG5kRKAbIHwVmiQ+8Qi/ye+n
enjn2XvtxenpAUulvLTwfq4ybEE81IvpUa6CL4WaexthJi5u/TD71DhdeXJ61yP3
2vYI/6Y7uUk1FTRaGoOLZyfqeUrEPc3xpgxOv4MH26i6OFDTV5o/fAFiSZI58lCw
hPH0ZR6hNu60IT5u3j74zN46PlFZVYROfssxehG0XlxneaBV9iyUACZRjT3Nm4z0
hXJ0bnYfuEuxzyLXKWhGXlZDBCawgBXS7MuUIJlzK0CgeGPgcVfOYajX/ftD7R1S
LDmJkBBEwYLTq/OpbED5qlG67IsZI8OTnn5KUJQCYXSoobHeNKGKqMPV9YI04nWq
DkRxaCdPCgZJbzLqWvPWGh2iChQcVOOBlqxUmZvSJs5ZvzE3wc/FKSSYqlWbW09D
gc4celhd+sKLEMtLw8+aOpE4jHu6FBhpkHCsKio5tNTKsGTMnH4CTo8cUFOQ+Hnw
vEDPtlvR7mndzGUxNmayHSEeWju9FvSvgVnIw5qzsm9RfXXzvGQnVphLdcntItfp
rW/u/NFSFjqSYFW2vWEiaQ==
`protect END_PROTECTED
