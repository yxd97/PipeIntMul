`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nMNWyVmKYz2epCxv2FECDmSd7bnzP6SmzJkt3ZeItCkv+4Flq3a+HMguIWGLTmEM
SnY9hpti9/gV6oPtOuKS/82UOgE7lhSBSknHzh9v2/byaZVt5o0dwx1e1rnbs5uX
MFq7uql5GLB/qBu8jFLeNf5IubsAfmIHHbBz0V07UOCUA6wf7pncXPbE92eU8WF4
78l/mZnXwNvK1tUKW5ZNxRtPuLYr0Wn9PGFxmH4TF7bMhG0441Cqri/hmPms5P9h
NbDsMBwzXFM/WRvdZ8yB2rEHZQGogYbkW1HjiREPaG+rZ78t4fA+2w5TBRuEuJ4K
Ku+Vpaqd9cF9In8B35UgbTS+TuIzTMrVdkhT2GhBZBa1u9fxTuaqlTZk8NRcKl9E
eQ6tSOs3fA2VSUyvn3UBPg==
`protect END_PROTECTED
