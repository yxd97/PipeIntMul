`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+1go/h9ypCFrI9vrpurYY0gxKHxISmpc8AApQdKARHzQPbuyy0LwOMV/aPO6ltm
g3h9U2z7cuvbpiYFHKwt6NUyEL9Dw2/h3OttqjsCp4bNHiSutZ1oM3oXtRBeep6m
MoO6bMnaJa2wjrB8efjUdliKBOy/jbf+05c0doBkooNLAsn/uZA4W+0AQABpPI/Y
3rzBkgysQ2a/hda6esacLzwH4uXloAFSfWUVKarOysoLZeqc5Zv9fHz9t/kl/WnX
78T7z8EuQHrCG4RKdWnLz9MTZ5gsVmOVkI3Zu7DQxwImVrV6zrYIKsx+Bl1+dqOg
c1qM3OEWVnscsm6o0W7iVKeWnYvWob1ljaIUy6x7Fh0Fr/j8nt9bQ15N5mlSaC2f
t/lBUQ8YH+qHDlzxBrfQrfh6a+tbyxGibR0CB5+3ZwCNn+9j4ZQqOis1jy3E4gxq
70DxpQs/1ptj3lNlW1bXUlzvERrYKYwkNJh+x3a+3og3SyRU7vO/CYMMbASC3XJK
2qBoyTbH0UyucPNqMl2W5e6blg7WJcG1qNAvtk86Kec1a05cFTpG2M4ml8Ucf6z3
eI+34YuQM/3GwsDnGav11SIkylxYRl0fdXDLQScVVo2Vy3ISe5kNm13Dhn89oyDe
xZlZXbmyHtkpRzvocNXcKb6Hd/UqX7M5tFyZBwxu8zYVkGPsgouba9RCAI2Noz/T
Q3BUI3B/HriXXTcu84qXYgGIBLrjw3aqeSYMkOrajTMpWluTi2TQtlK4nhz2aT0v
AFICmsMbVNgY9BNf7M7sy2JCes2P+DPorEowt2AdVh3pmlFlvuiE942fowhDLaFM
pXMUS0dLIS2lIZfM4tyyrMRWcQr1p9PMYkOivrkkJVV0JYRp8E0VvE1utxWQShW+
1BGQCvlWjIQHdhNOaI0WF9M6qOia3obmuoDalDZi8nG8l4t6+BF6uNU/s9EaVPQU
3Ina8KA7E4GnHEGJC6NrBBSpzvZwrDE9UYi9TmPb9YkwPPo4nzORAxc78aQf2VPR
W4AEziEORCF8dXxD4XXZ8a42ZCtgohECzB27HgTHd2Ufi6+Rwa5vE+yfFr23y7KQ
amzp8kT4GiH9d04fQzIAbwLg1pdGZewSNJca/M3JJH36rIFcPwFiNr3lgYIl88m7
dpt9yDZAkktXHtRSOP48V3F27p1NUzdu4HbSk8Deih2Ia6y8sfJMwjYZNZ4YzHsF
l1KyXdvnMvYQLf98ldTBQDI8OxxhOMCMFU1DhigKqy5F5kF3r7BlMEz5bvlOQmGk
hroYZvI9QbuIXpbE2xnBfKm/Vv+PYlCaY3WDFrGd3EhW6Fb1/yui11E+wcgzyICr
oepRvK0pBYHYn0JFDtLYnJy/DTRmSLFNIVgMAPKzMPsQz9mm0/TtP4nQ0glSsL1q
PFvz4pd5X/nN8rtVL1UGECjW7nsZ6+ybDQGKK3xOtBacsn0GXldDdgiUFD5XmvD1
R3d4YMmj6BBNsXEvcN/5P3Z7kiO9jyK4TNRtAAz+rl6eNl8QWP3E7NDbO6qZlgZA
IZYBV/6ysrfx3w1LFGWajPZS2LzYS6XtMS1kBFaqRGPj1EeHW3bdIbSw+/YzuQO1
YU92DfJID0WSRKbKdhKPTBCFkX1zQuW7BuF3Sh6FJ5AWjAXxrGfS1GqwEMRkcHsN
TtT/bUlJXj09yA1wW8MSsOZJ5aA6IOpcUdIQMnbOY7xxx8OdHT0fGSfvS4VFBoC3
iGigdUBV830on7R6GGp9lb8jeJUHVXknxJfbyUMeXYyBE8uYV91YqC0uUdR6TshB
cfAHGMCqGxnyGhadXgyokWVL5O3UJEqc2KfkFs8KZJjhhK+l039/uf6Q4Np1rNkq
/XkpdZhf4UT9NoJ0hElAsdq5e+fzSIbO4Wfkq7U/5B8PSmxV6xU6VmFTenCwlTaf
dMkJEQRs9+EKTp9nORPnpZdw3d1czxayZbVglH9plgmDrAalAI8hGRzm2/1Vvd2P
EIoITWlkW48GmV/wiuebmcajOR9Ww05NpVUZMdh/Dh3bs8zYDQOhL279VOx34ceY
g0s3RNgz4FuXIEaiVPgZgGTMXf30sJ1WKlBxKTjHRvL5z2J2n74CCptohmkwYcTm
Vll9xEF+ekEt/aWcQcbHIb9ISa4PmlRIo8s6ikxaxJrXQa5pMnaVA1yNKYXYFmPR
DCh/cCa2kMSGBN0hAEgWBjUExd+8aMRrcNVWcYjsotAfGH2FRWP6jF51KTJgRZT+
k9cSBl0IPrwIpFx75yYinD4Niv1wrZDtneXmyDoqJOxq7NxDvfxjDUJSv4WX90xW
eHOegl9ZujF0/P751Qvj4aSbutGHCumQEaVPIUBUA+plsvrtvaTqizb5t1Bfddgw
mgl4U6VgHplGmtFmV95RgWdh10NBn1HjUPLMv+ZmBWAhy4YeYa/xKFpz5o13/P7Q
zFoHC43amOUUf+w2qanBuCPJyC+/75rGkGMwUynExxkYEITHzC31R4FcNQ6XbVpt
+WivFaSD0KVeuVGK7cMlKsSwnOc4VXWkitwz+lk4PQrp8xty2JGEHVN7IFFj1JOk
Nlw/MtVWQPhdCJoL2x5GG1ELBapWAN0IvS7d09ZGHwTGOimmqPhyF3SRhqpSxv5C
WHhi4QhMsskowxyQ91jI6OwmG9OCM4Er4iVPzAJ31YEVk5hogANSyUaE1gZo5WA9
1B7jmPqD+TWUEJH8+7WcGh6cRqb+jEuukU7T1NVGfKYDQWedhXwKstdYZCzD57/v
n2z5DKrEgTghHGzEz8yOtEo2iUjEPjjpYfosWZGUfQ0Ktw5UrBrHi2Yp/Jp+9QOh
AzBGB4nfRnveJGQRrQ8YS9c936WBfPaaY4heXZp1d69XTj6EVqTMI86VwLqWeMQg
tIiQnZgcnpRno7QJM8vYFtuBbOkSmdhKG5XPXbkXpDQFtgSy8t172/qNv0bF++Yr
cMCQCQbuVBdKBvXm7BPCfkOmTmoBifsrOY+Z+0GcvgbOjIX8x/pVBAtB2KjkCUAb
VCZzD1Be6FapGVkSLTBIdNu874oU/u4Tr217YkBpAUxdxO4rUzQ6IMRbfnJMeLGQ
owi8lo6QzMZ4bp+B6RqSQZ1IXV1GKaG3DVJ5DBwmBzjjPpYZMw+qoBz7/RvCAPCi
vPkZnfx8o5hx7OsjLOfRjdv5wTPh+W4CjDgHuL/r7YhBDR0sAILY137psJHQ41dK
NvprvmlhD0L7ndWgao43SNEIVt5gjt3VbU1WZdKSOKYIt3SDJ5SkvOfmvT9fjYf1
hXUWOYjuClcETJgMr45pieISyZVeOpd4O8c8Ef44MqIMCnjYU9tMMtE7IcVNTCCv
uTS+7o4ZJeTPszCsUq9TF9tw8vS0MGYJ55HWTF1oHyctkThUIxpphCLfUpyYrFqB
D3td6cGoXTOoKdaKj3TASSOCYW+n3FZrD9dEvQiMIqcTBOPk54m64fjcnOg38AnP
F94OlynArusIJboewmB7dDoLClDr+adP/bMgFfL1wI3uSnOAJMRooBdoOpigJ2yo
8Uo5St/l4zvaWpLzuPK8jNtEEKihgSxcDdswICvne8q/rh+COCrHD4KdiQO8rAxh
mKowhWU/i+XlTDZJs4OqNcaZqlXQ7A1T/o5IRnh0zSwm86KsgY6ApYFIDppdHkee
T3q4dwxl2pGnDNtPQHjBO1410g9cBxVStAhjpgaZHF1Sy/D8K0N5x89Jpjf50d+C
YobNTelNd5Dt7VoVFTr3S2JLp0Pr63UfihI0koI4IIt05UTFYepz39s08d2muad9
dznIo89cNJNkv8iOu3YFVatpjbsdMo052+46bZuJp6Cscym/xDAlWFg2X7G3h+F8
MY9CkbKOaPrG7t4+2qt+Cln3WJbfN6/eQ3r/MxN7N35oeBnzMThU+GtuF0Cm9/TT
xq8vXwKdyK6Qp6bHMKs0ZQE4G7n9l3QyXXqPR2IWHRA/Z98kIjQjSEPt49JzdJiQ
Qi0njJ5iaB44iqI7nuMFNHTRUbB8p3kFH2B+vXoonVfuhZ+/r2S/G+UNkAlePjs4
/19mr1LaINtQJkDHeePyEFP7pTA6TrGWXKt/Ehy6dM88SWrG5KNg5YCZWAcO2Yuh
ytXa24XvuUprhIRsOh3avcIE72YYldDJpvXmtWi7AHaa60/j74N2A8VUCIH3x+QY
v5ZPhBOKbVOm9HKLUCTtSO57j6HcVYA+FJL4sbwao1+Nu593g8Kx7QaS3+gvpvuN
yyZVQiu6fKgCJ4EypUG55YJt1MRIlJsd9Qh1YJb7jQU44K4NnxDFT8prwEfyrZJx
Em31SiRMhNu0dy2U7Lntl+DzixrcNspIFXzRZ867OVr7b/JdwPZZxHBuOzROus2V
BZELA4k+nRyUi8fZE7FQrK1VhoRjXn6oYqaZna8keoU=
`protect END_PROTECTED
