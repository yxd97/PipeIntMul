`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pmZu2vH8bYMfpE4/H+D4FztyCtPxPYcwpgpG61r7oytCmvfEm3e8vEZOzySFY/3x
y9q23gcMXNVy803zoHzwXDGyHOl3ragPJ75NA4hE40Mts2PdlsGs+YG6qi3cTWjP
6KMIbPnYW0DjJA4oBdwBZ9q+3LCzRMbVOIiKFqcFHT3nmuT6fMN4KI5XmaYP3OCA
jSU9bYTH39zj3zx+ipB8R4ABYY58wXtatzLurL6PeLo6WEgiNxffQq9i8QWJGGlp
3rgLfHmZWpNuZaJ9AyNzpQNdQcE5CB7Jd3pK3fM3AAm/htfWVSlszO30oOU7yILu
oVNF43w7foM9276KLbmdKdHvsl5YFPNkQwinfExcgTlOdDQ6ztyZDd0+abguK+9s
wh9tvRZIldItJy4TXyvSOa5WpQaruB4DbEwyASQ6KFhFcQMOzwuc3cOOK9f27Whn
iKY2WfFPcrW7n0FpG7wcbKZbdniprFRKzo7Ifv9WTV0=
`protect END_PROTECTED
