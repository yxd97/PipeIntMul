`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F4+CRNvr4aFthRViV95pm9vjHy63bc+vrAljzkuvq4ZUEU3Cs5ap/nHb6N2p/UGN
COzsG43RYaSiQU54H3VOZ3I9OuBnLRfujYaz1nNT5LEq1Co1qm4wST8WRp+TTBtq
V31gv27vw9tPSAeFnC+EGqTaNNcgPz+DPeMRB9ApjvknKqUeI2JHYiTCvZpDFLX4
Ylo/4l66godaYiLq+yDNdTxdhxt88foQQRkC+BtueuxqRyUpPUvWvoByPcmCW1xV
zJywlhddk5B47E+we0AbNJy6FlDOSuk+DNEZZ4zvMnbwVP56dIeXdgQ5nJmOI9RI
y2bOvuZ2uAzjK6IbKlM3iRuuC+ZAwSsrkDR+HiHQQtdTxy5ZPX2JdrhJTdJ9wOL2
fJJcw8Y6hZWLYDobmtHUcBfRVAV4j+UVm3ocvZnwfczV9kW1njvc65b5VACd8aw+
fA26KCf7jDVhvLKngRIliuXI93fF2hQXv1VgDnkn+cfhLVvBboeadRm4Ux/J0cAy
Kx/M3/Lkp/mc+BfK6XFR+XtiSjzkab/Z8t0L2V+hoIte32n8GRh1kYgHwMw3VFEA
bzoQv7u8qUgweB4sdztgE5Vom2Zvg8ld2iyPOviaiZhLn2BUHDxXoE3sPPvPbo35
X+4tCEQgBQ433agLRWtM32/KA2arONBPdSZ/9pMFZCVdsfQ3GddGz/ImM7gbBKN5
mdmRQ4Jh4pd5RQtbW9Q6hZtca2QQ3m5GIh0ns3msuBCrDqf28N4vPGf3IXrTg6WE
M7SM1dq/DMPlPsZdRe4q/u0K0O/wl8jKuRaoyHkBbB9si1AXifjMBS5IOJ4VAzge
`protect END_PROTECTED
