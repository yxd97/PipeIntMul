`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2b6CvGkXF9onMM3g34fS+KwPEHiIHQfYTGq+l06mOXG0V4TasZH/CXp4npDANZ1t
/L1rw+HWCKaIggly2aiCEb81tp4nc40cSyDMkBT6ukSqLqj9jxd1Eg/IdrbBoIPz
Te0PaR3XRky9JWUIPMXh62QiKakisV90cnGdzwwoky0yOpX9ooOsoHbm3j092YC8
V+0oDCwCVAk0i1FtVM8oLycQJ624y36xpPjxxEPFlyjbzgProdx3OuCBDM6pJhR4
n6T3xqE2/ekYV2yRVXFmwmoqgCnxtbM3AZnoKmBUuAtuq/UbxStqZEBYL1TUePL2
Ce33EBElJ6SHmYp/jZMFH9Za3KppPfGXCD1kEZ8xZ/9djoKfPadMmdDUPmezDeLU
Jfqt1K5PdaGl9mgEfhi4CNjkTDVTg6u52QouPByU3XUfSdzyYxgfG2cQRf8WllDV
ZYPi07QT8YJDn3B7fXG0v8tJhS0/33U9eFh4bA2PGLg6eYWp1g55HAm5DUSgTt9J
oJPnToF8KAxJQvtR2zeE0HD0QsZzni1DKyAXBg4zBu0jROr2k7vbNfUTtb0A1SPi
FJyH+qVsjS12ybckssIH+KgJnqSGFmOC9luGY+fi794Y04sWXo9cIlBpkI1GNbG6
`protect END_PROTECTED
