`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
piZF6rwkrR5M0wmWZczRLnMGGEwfxNDlw0GbA5P/vCxI+ZfAwjC7trv5t/mDjrYs
aMLUtpD7zqyK7VACO3WEVrYMu8Ere6FFHpkQPsBgvIf1OXNiyKU6mtm9PBitbCqM
sih++D0bWXYo/+wwkA4/JkEVCryPUFDeu9tkUBN9Xqy/LYy3rwLzQXXuogoVlFca
nSknndiGBKvqpMvaG4VA5ARbdguNzYzqkVRz0g29enzHp1nW4TbHcCthoR0BExJW
rD4/TmJopvgnNF8ZWzLrRjPulqKzIumrg/7yO2eIl9SatgJoWNAEuenB0rb2sRwU
YB+ftdlS2w+zlEhjClkJDCyMQfPDOItWSD2CqGAW7sAy0GNRSgFi1PzkhhrkqymG
CiOSor51TQcbDgrTnVeR0r2exuHAuePzAPiW+UhugmnkSQkt00b7NKMEO9kMYVfF
YE9lLKY4pNBYLDi8m59WjZEPKnvLgMBMPh+bipzZaJ6HWvenSvJY055L9Gp8EScF
sREUfs2S2ktGt/36OOQts9mWb8nlrooaDil/LKPHUOI=
`protect END_PROTECTED
