`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BoO/4EfH0WL0BAO8avK60J/9SAcTUxafu2m/5Qq6cDlzt6jYVGHkKEjQE1x5JA7B
22ep9ivsfIx5pEHlzpYVtMMIO96TfNYYGPZJezSmKgqgieqh1OaZrp1WzvulE1Az
S1YcFC7QfioWZVM1UoNZUe0yfiBtYdlS3/FR0lSh5JsxOmG25B3z3Dl9PUYtP4Cw
KYkZ/ShoPntMW0sVwPveytel7oSjVEio6ZZpRr4Bad/V+B/qLM7fB2x0Y7YXZWih
fmJz2oh4eCwdUr1PDPfyT4Ljwlhu+aFUfsq8E4fSh1fb98kg28NjxIMF61OZBIE7
foMsakmMJx/1INXVKXyUBrkBVRTAJ6fJB1kS3rQjEbVxhCwN8PnrjwrucQdhGOWT
kw9N0K4ZWwH7+GVwqcDCP6E2LO5yLW+QZfME0X+6Jujr479ImBxmRXeGIoJK3SzZ
wXIPesVM+SH3mEOYU0Yz5GJ25Tu3kLu3eRAP1aPJb2+o4cqhdOuWWH1JMA4IUTW/
+c9MXeXEfjG5WcQCxHVnCXXaqKNcVTavhR5tMMXktTxwBS+XtGC7OJOsTnPhrjFf
nDvB7im16R2juWKKUOUzmXLx45viQDfARQBcYViqB50w9Uq5cwPietvyVq9CGFEK
U/8SO6eD88a/lXk2kThd9qXwH7ua9xf5l9QYpumdwiKWUOQgm599wxCux9DKZeV+
bUHcJP42e9vFRjPQS6tuvbuqN4p4kwSuWTZOFQx9kcNst6DQcImBs9GhBUoFm7kJ
4tA/aaefb4wbwkejxbkFdQ==
`protect END_PROTECTED
