`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fWTJqwAdbTvh7FuqIqjdJw0PVcdJQh66p1uenqVgNh5Gil01cWFVsDF/aVYhYr/T
ZXL4UKekO8TEqw0Z7XJVGj+87V9xPbbupSr2JqLUvzUAQ070ffs94sMSpjPUD8E2
2BaAn1Oa9gwm0STXcmldbGZ+YExo8LBH00F9Jhjx+jBBLzVDPewyf5YL2u1e63nZ
hUvy6jTHuAHm5bFASu2nNHeW6UI4CFO+BWEfcxMZu3M21tyyJQzLUGBP7H7fb8Og
eqEB4/hU/+hBwEGleFgqNbDSn0YnHecXVZqiRV31ATKnaXHXr0ZZ01bFRI1Djh6i
U9MKFba7fEfyDB7pA6sOa8ZZq2kLLJhHq5uZFYzSIt4FZfSFPFn0vorJtLQjF0Qc
KgdzZAp1/+3t2Po79MHgK86Rp4sDYUvMOtD3azJM6mKmrPLQdRMJif7r6VRUwzl8
YumhHfu8EUjp/jDYIPcYDSEt2saWQiw3RsOgjhI2qgBKuVhGeLDjeV5PD4X40zfD
7HCp5C80IdyWcBCuqGXwjGBHOkSC9ZD1ihabIV7INQMuCP9QlZ5aZA1xS6UuT7Ls
4UB2HUcd3fGiY9P8aLkK063sVKgUu/IyCvs8g19swGlN53Et2X4a2MmqWAQXbe5q
D4ZFElaBZr/d671cn9CNsnkTtZhVjV/Be+7gdz8i8Pco/3MKbH6iDPYIxs8lJ1PO
VXjbh2GIU/ZjpEwqjXH6PJYX0nvIVJ1M2sQYI7HlOW8K01Xn0LFpK2Emvnk95taj
O3G2R9/i0tx1BGZBpFD+nklAWyfrqtft7u+toIJ+MZhX4yE9xzpe8C0AH1K1A5g8
Jiv5rrVPVdI0Nx6LuESJMMOMlUAm+rbh5UVWbYPyEuCgSYRE4fO4TLyvQEeQEKrq
LX+95sKsM4qJTNOW6tFKz00ofEPcH828hHynkBDDrnHlq+9O0GcCNTeM0oIj7LRC
2mmjE7l6Vg6evEM4rFnHiQysgQDSfJi33J9xUZ1xSJiCQir0AHj7jQUVk1JVXbEo
+2nMgLtO8i+yZ2yCkaHrARjGTxj/zI9SknI3gRyik+il7tKtFyrFvqmJNKzgRV3W
HyoU5klx5N0pER/wBEPjOr3S8vkd+/SFFacyMPWE27k9LSa0FPfbmtORI95RZvOi
YlaW6d7Xa3g61B/6XubYglahUfax+YHsQ8vpQ/5saZ+uYt/ELk2fwshv4z+SoEYr
wnTFqywEcyyqn/07yD/0sUNdLkQIkbPhRoN4/N4VAt+f2OBM9QmBglkgeHPLfIjB
Q9uN79eIq1jFdFV7Uz7JvziS9ue36hXzedAoTtJ9817BrCyHpNFzZ8AqKblk+KAQ
AoOvo5h0k06hm/ZVL7msvpKGIuNTGUU2EdAKmK/xTyvGKUt1ACY2Q5dnWjkEW7FS
o/vVhQH9GNmTDPfXqKtGb/BDwG9UzwL3XurtvLgSFJeBIxxyG9xRFLUkmC2SbXqC
S8orvDEohiRl/Xd0a8pfsXiLHfZ9GyFnKRs9IFH+XA7SEQcaPcN7Unoko3LDLib0
HGq5avGdRWHCtnOxIC8Ach33muNsosqmn7BY6S+BC6UDMb+srR3TmGGcNgo44pVM
pqHbie5x9ZgbofSfyOjJ1cbj3930grb5FuAndsIbUYvxQ8+wonFu5x3Bc7hlixv0
BsToxFhBz2MPuzc6B7ttAOMXuIU+bplN2Ugn35L0Kk5z5dTEDW7Rb9WkYr5F7qbv
ckgdhtGP4fnprFUbX/ajnRpTByXwQ0Q2BkOTiT8wAohRMfpzGP3/mHquJ4j80KnI
BUE8/tVMasF+Hdrb840Y/Zf9lT/rvLap9GuF6H/++l9EIuEcpFOBDLXDyf1w4xp3
f5NSMTrb2zZTfmYaqBlb1iryXyHdzaMduzP1ZWObvoFd2tRi7Z4T049PCS/wueeI
HQ3gzhtGVfhMkKRQqEgn9ZDsx0x8ULYM4f95ZaxosfnjD+wEUZb3ZlEVn9MSo4WI
gKVMi6bUnxrQC/kbJE8pcrpKCwgMpMFE7wQqb1b+0EnAnIweAevBuVHBd/2a5Wev
fQDeNY9xwrVkzTPEv6Qjeii9/JRXWynJ1z3Ht7TGtPFHy/HjxH/Lc/Lu6qH8vFcN
jgM52zhGyJZgpam25EYmMrYXXXZcajQTC9g3shdGH6O9VVXmRuNr5I5WY2/e76E8
KCVYOA9TbfHeX3hgOzrmZr6w/SEKXn6+mKAZhGyjHsIyKng1VyXsZut3Le0p2Pur
ai/pFw/RqLsVq5ZDZglaCWzK81vtCY6UJL3z9EqbNF9XvkWWcPxDszcjb//vastx
p6V8MqeSOe9ZMNUfc4HAKzSqnm8RNocTDLfXLkFBND70MqlkKyWDbvZdMnLL55RQ
SBFWSgwSUqH5787DVNBoVdbuHpG2Cds9QsvVnuDe/0gEP0oY/c+DYHY9MCCdB1q6
KUnSTuSyz1krTT6JpgJt/GhRM3iErQQG64bvsUJUvE/spy50ihYHOWaPA2VMlYFa
aRxN5PxqUzeLUVVOuinxC7Jk/Kf1tPkwrbCRiaaOylP3eqIhWFDzuFCzEhbocSs2
1y9zQq8r/nizIiCCIZNCfuETYUi82gfDgDBvDdzMXYBcDKmfQgbZpopRjHSDNbdB
m2z6kyvIgZf5x/Vc7Nv3xIFYJUuclPB+wGISVxnU9wiX94Z85p88HiXeC8R3HAp+
vHfDOthTtfg5O9zWksJgX2sCsPlsG4MjgIcaeVV3dNgLrjZ57cR1epaGQHGuw9nx
jQzhE9NpBpiu61zvgHTJuer6UtHEpezTFIqXmLVXsBextpT2x43PVvEU+ydEdYwa
ORVbE256Ph17yh50hKtMz5YPYjE/fngf5mTzC0lDtbZxgIYd7U2GtetrgsGue5nV
ftLwb16TKr6up7lYfxkZDuyfJ8zBfrj4E5Th7XxxFLLwH29a6N409E4Bj3vvL2wW
WyVLKornhp5U/E9oPgWcLer7tqsregFxm9r5aYERyjMTefbizF/U0ka2S/XzUJBr
mOCTc7CC9CW4tdsWfZIf5Z60FrcjSZDiIYa0U6z7A5FDzP5viSsIF4wjoLhV2guI
untmvGUacr795KcjYun4pBL6zmpxCLIjIlx9xVJH3qA7nUDzcU0q4tZLvW4s64B0
8k3zjhcDaGHP8/F99kHIJR9+Tbjid7m6kZWSn6/hW0XfYTMgBijSdUIYM0rJ9dvK
jWvve9YQXvSw5m2s57e676E71bgkmwhTT/YqCFHPB9Xbr3RmTfYuVtcCx09qBCKg
etVrQTZxeUVkphtl+IvDGfvrtAAJ/8K+KY6h/pLuxLC23+KhOEI3dSZdLwxyPIqY
pCGLUJWGcY+GI1QxMBFsM+Xt5rgsXoCHDWqfWUx5gROe6yMGtKyhvSpK6xP1mFHX
zxJVtAAp/ezkykevMVRfs+gocdUbaMnI1ekykfAkjuU/Mj7zdzeVPWqQgsrsGxjD
kBKcladfGFFy/rRK7c7VZ5knLHTAkL9rro6cx67XhqGYxqXmfiK0zuQPEhc3JQHp
Uv7S/mjjERryDRGsx7py1RKlHWgG00HRM/jAGgBTTXl+QSnOsQmSf36lRV15GbSD
gjG9Q+UIcNydQ4ooJ57uaZL6/PUJZMAD0hpp0S8AKEfCP6xiPSPPhX1YD0wo5RFi
a0DWP5/qtl4KI/d7ULc7wniAI6s3XC7xWkcdJ2DjvrUA+4Rvf3qIzVvO6/zio/Rb
LCiLlAJjrDovmLS+SIfAoGKhJQXSgEYvdOEs3EAi6Lqp8M4rXLLXBg3ITiDmxv0Q
HYidEKLRUmzTScuiNLbGvodma3CPJtpsou9qUbrNMrKfjzen6MW3qx1w8wQNvXRx
VbGFcvPGayytydDoAwtQQxlVuQop0SBKsvHjifw5KdbNMrAUJwjPhTAAecE95+cd
98CDB+EUOywvfDF+k4A52N6fLqeMB5pwU3OywHz6+/PoW+beHzzV5IxL5EJqLp8X
EEiPRN/GiRrjaM+TNF52oAM/8XcB+oiJhRk0WErv/NorKwTH5t9pjqQOdWcNZj4K
WJPgwuhsV4vXdt0ZJLGnFECjNOPUEOHGsTDLQ46OsC190ndfycQYTRC2QaseXoRU
v2bQYCc3V03EopvKP3k3wSsOYwzy5+4Xpv6XCEzJBwWZ8WvC9ecMY472JfQSgrtR
xxVv7CabJSwnwbnr1P2W/TnZ8RWdUI+8pG4/dD+pyvGwEzFIN0CP/viBSFqLuN8f
z9A6GiUH8kKDU8btD+Fnjmsy3pWf7nNRdd7GDg4J0zCY9Ac1+7TrKJVZv7SIOjZs
jsHmDnl9yE1x8Nd3bCERAI4EGe0wvTACwGcc5hgEDujNuvCD9tZAvu6ELOAPrF04
okpyEzgXmDlBeXxRx4sehrIN4vizvkBP9qTL9nm7oUQACVktgOgjyHIJC9T5yn6v
Uc5YBHxhR4BNp2rIAyySVGmo8/KUNNJGVOqU9cd/cRSi5szYRZaeNTMRIPjqcneo
f1tmJqhBOvdlEXwfKjc64PRSSpKbnfyADi7Mt5UcOrgBgCWwSndvnMpzswOJ+1/i
KiF0Y3dVW6Zrem6l+Hor1NGnsb2YpEek2J12Nrkhw23tpeZOXBU+rSKAZoe8Jb+/
c4aXNv9ttHJhwUtLTDjm7rTfUVtRb8J24jiJ1ojDK/rvz+bazp/FgbdjTanUIhLE
4lsmtSzdGuZl0eFxm0VciyslTH0AnIxefG4tL+CpwYu8as06bdxJA91xi8RfWJzv
Rp26m8t9eVrXyGZkvJMNffAN0yaevCy3x/gTQ3I60RmFYSO0CUOP1u1YAIp0kWNf
deFs2gkkPgCQn9uBvcKLRRbfbsAeNvEyeBfWVkqt6y4bvyP+G1moxZIZr6hOe/13
CcMcCp5jXkBXajLoAxXNNKLb24GVxdCSmpxPCxhTPlbkhWm9VnH19CZQm2Cy9dFk
ZvqBPFECWTO62Zq8cp1zYK0do4EVX8Jqg6GNQ4WKbVZN+RpGgGu7oyyah578Fu/W
HZ0Iu+p2hfJCx9ZqDYJu0a8UYTJ5tntVdoob8JS/hPtDdPdmqHFjoA0txsGkHzHU
j9cmZPEkG4f2Ds52uw3sQ5XII5hoSJQfXpef36mXP5yEJMN5o5uNKeY4gwO7w0G4
VZuOlmjf4yse4mpFFbPHHVly4BEZ9EsiZ2GAzX3tOEJMBMKM6G4aX7omQ2hVxROH
VtKNNTuoxm+5h7ZCTY9spz6LZsisTkGYizGs2Mr1IE3q5psMzc1yaPf6cIZirIUI
OQbmsH5Ta4w43g+eU974htJsGeRJ6GC60pdbw31zZ288NEcVdZLMNqWihv6/KQ4I
eanT1QhRbMWtAbDSQc8WAdIfysjL/2m0HUm+LD/UojHpZWnDU3CHrsbOwzgTLg3Z
aFhFiGx+v1dROH29phu+y/NKQ6ypbaQZEDWkWpBKdXOeboizJDGOgLHAek3c+rEC
16d1WM8sKXYM3GsjeqAmS9R/fNp5vx0wh/REzAfCLfB7C7JBT41qXShpE4j42kk/
Irpgvt2c9eYcfOLD7T/2dlprGTt/cYNDrAD1GpIHyY7otO9QdOWJb7GxGo+fADTA
PA/wdfuoARAX+vVbljibXBMfLJ9IFGKpEZifRfDMAwJwG1RTdLntR/xH31EzlH7/
dB0wmFv9uyLLek/o8nNSlW+KPPnTrKsFF2h0FJqiYTdqxl/AQlSFtRWbIcPRYueE
BMmyd8xJoADZgu5OJsQjT90KTWY9EZwS/DnH/nwTFddlePd/o8pCqbwVEmFVGFm9
B6wS7aZyTRAcKjNu7HA9EHRHmNEPVhDfrjFp8mzCbns5d54gWf2TDtnbSf89WxzY
sZCzgXYIguqfqJXInSLij4qOMv30vTkHU5lmKivBNb9enLl1cj8pDNSoGDiuszlw
NTf56deFtt4ORyIQ4H36NXUafdDj7sTlcFfmZYYGCLDjnzS491XQqJel+jwH4vcX
TgL11pVgK2wtG9DNnHQSRNNYGEBtWclg2PosmZ64ewP3KvwOZeKX9TIyag3iFcjL
+3OjyHJ1jZN0UuUum887NNiHhXxy2brBhsK2BiFwsFIekpnkilNUNdQPeTycbwIM
eiYOS/Q+OCnHsIw4YGr5Yr0hUYVQSatBkUneH+2GKNKzduy6QkpN5yqG+VjGq++E
Y/DMCeyjvlCiyT+GYjCJZyy9BNVRjT4U5x2VQtXpny9lLV/+C6cmZ3QX0zoePT1o
WZ1s7l3zpjEkj57XnNLw04RgV9Vt0P75td5K1WqMEKkhsBV3W7qHC5voduuGOXrX
Z4QKj+i6gPrj+czuYXo6UiJGmBob3r2Ph/SHdeb2LBVnL3Kfoc9/IKyJrxTNeSSg
Mkuuvq7DoZl3JbnBYh6G23C9ya7XXHgsjtWAp7xudWRT7XVui9gHBtNxBdXvtM+0
Y64u6ww5WUCT4bIJcxULHD1AXfEODYVyGhivSAekEA5TWUOwLAsExKS6jj3QcYBD
9YbgJbbvy4fMYvvmL0t8AKND57Ri7W5gmgBe+4x1Tlh9uFhRlCSj/HWhiCkL7PuA
W1uVwuQURT2TKAECLffkGUO5WSVPIn9m+He9H/RN0RgbOKRKnz4HxwycmZZCBb5z
YSYFXcXVS3D6V+PU0cupQtIIb7y2uQ4+vaQP18vjyRq7a4zN4KQ5Ti9eBnICtvrH
6vy1wPevhHWmBfUad5BStoAPrMivPvjDjALUCa5xJHUWQt6s1LiLg3rqkWeg1z77
hb7G9tMOCOnyhUvCND13h6fRXYmqLfURddGanYZkN/S8foG/6AyjzQTiH7mAgsUr
aogwcrWj13mifcs1ZwzDJiVCcHhiNacSwgFNDfWocMA52EoKu2t4Ee8EABG2muPa
OO/tobTgzn2rSvGl/BW2e1l4FfRZYUEDrzVAcbX/AWnvPTNRVU78yS9PJLXGvYQn
YETgmt2xS3pjEU5ewQA1+djiVwovHjPTQOtZsv6S8r82bhr9oemHvSHqIIQL0qrR
6CdoncEi3saUGIhp4L/rmLzmF4GqmTdvQl7FTluV1nntU1qm7+tvVGoQWfJ4mRgU
24wbuEs3EyWc1GXZ9bdVy3MKu+JL8fO+Z7zGx4d7xIFf0wNYlkwbwjRZteur7nrq
to5uv7ivx/a0sabJuccnJh0L+h3LPLld5FrDlyhToX11GF3SufHV9yDbFfVM05gp
WNG5qXahCcTzodmDf8zsb/WhsmgAETdfQf0zS/7Z0615dVY/imq1yGFaZlgriVD0
JjfchWTDpf9YY0aIa2oSTXxtztDP8uO4apOTSLyH67WkWykfcdJ228jf0+p1h/0s
vKdSWAcovNGeEtB83m/v6pZuHl34zs6ip1aNI2RmvT7H51wz5F8XTeDIG32bjy9i
yCS5MJItVy1i5YPV7k8cu96bzx10fkXaDBgSCRnsvGDvmJOxaSAQaSh0mMkk7Krm
7vYjBCKgiBtLQ6uHMntZ6UXRQIlHHD/bIVc3me2VLvLqEebYL2+Qjkr0uE8lKPji
bI69pASGJ5mGIhtgv7b3F6/XNjB4jvVuA90c0iBjCPBhYc7Kd8gPlrrwxOQnsAcu
PgKuUpfxVvbnJ7Igfw3v59nYwqflN4hIulmXiqs//kltT7RHlcp3Y1bQVgGZK64I
/vi6bC48wR+GB/Pyxu3UkJWCfLO5/HC942H1oTBrjDvKn18lnMtRe7ubB9aAJm4x
P1A6sU7CMiQD+03byLPyPP57dsTWPBCelplFQ6acIes7DwNXwGlUctS1wg9h3UZb
bIb/GrIj+T3EQo9nygKRcE5kzJ18xMm06BHF+kpFU9Y7BlIx6DuibGco7gZvGRKM
vbaN/oS8b9EDZxa5TflsJRqirQqC7i/RQUejnMfwPK+5g7wyfgpkGqjRvJNWbCz+
2ZwLkzU9ueQgBoHoBoehLsFxuA5lg8aVfmAiO8l0sfGiHuFYm9OM7xNGRDAK2lro
GXVzbpZazsk23Yhjk7K8PhGnmSp8x3biCtomJEUt80Dpg1k8zUrQGOuEBQcnJBGn
Gki1+suM+RTDzYb6awUUllE7qgJWCCUp/4go4qc6HqoYndm7cPsDzy3m6D8Liz1v
wqEfd/n4lfF+o1FlNhY51J9+FX4nCQGauZQZg3DQ3k8VAzG+n6vwwMy+hfoEWL+N
BWzrj75oxmkBds92BOs0WZgbXUSjDvjKvQ4En5vqhSrlfpeBUwUDkAzvtY/pqUbN
B9g/bQKko6aRDb0fhFQMidV63K953cvDEFWaxBTHyb4ljEXG5uwtW0mqDtzmVYP1
gBNYH0fglC7VNs5K6juH35KTdTjwNaIheSlbGal7k3jJRXiq5nC07H7SRxuox1+x
iTbcw3BA6yfRV2ffkiaZW6JEp2oYjKrMCO6D3F8eJPCqZyXIS7QoD7pHo+wvgTCN
HXhlAWolm3E/EBj8qca17+PUJVPxXYZ/Hh9ObwaRrnY+P/AYt1fUAOr/3z/wXk1V
/smiVdo0Zt1e0G2lbtRJ2e1UBdc/WwB/kxNq8aDnGJL1Nb6Fn6F6Y7GHF5w/hMLG
QPCrxwHap9RHcHm6eZZXC7JbiFokbWrA//1KXX8a5KcT121ALExRbFgUvqf3OSYv
b84a0oUl4TZvyXxYN9jHickYHUfp1HYHaohLDMjLMPkuG1PTgktG6TUJ4p+rVm2o
3E8pQW+oadPpBIHkSzL4IKB+XWkPUgvfovar0M5v+/FtCOs9RWxNeRspPiVedgbo
ifTxGUO7KBlYLfEcux20fNG+3OvM9NkL4bIFJAi81xAalXZy0i0Ipv2q73H1CpUg
hWECkXKCxteGjJdsAHSYuuBeIoDB5LdzgHRcA70+A2tmI3aOPb/ozxZFlEVNLkKB
D1CeGwa66C1wQQkQbBNct7bALgeJewFRt7VVsNDVgWQ7FOoe4308xsDrwwDoHVwO
zZU0E/14ZeVIMGIpDcqRzosxmS3skxNCIgVuD+DGHW2WE3NVawnu6naF/F3VM7qT
9edKv09FzfFhSf7Y9kdyORBJV/O7eJM/hTpzefJGtS0WwhZbwUBQ7lI4R/Pr0byp
bwdDXNzcDjysQyxtp8ihbCh3BUyqfIRFI3KBUpQB4c7jgesRX+Kit/WYAPKuf6LT
t9/UahuEsugmx8HG5TlRLQHnxGQegNbj5kNYAGav6SRhfM5lzdvLwD3r7x2seqU5
pwwsT0X1HjdyvNsti2eaIQbOThM55KyMtoCS3VhZAQJYrB0ct5e5jTw9QnZEcQ72
9Z+kRKprks4riNJTO5rXmirXOjgeaPvMCpT1tsM4UON0I8J7IbocQgqHdZDvrJj3
z1mnj6bXmHcacLa2rxARE8JfpIVrylaeCM01D2O6fNlK7ef2k5KT1V2qkWJXwKr2
9i87ciRKssj/8TKO6ZSoNTdbKrMpXb75L/nCRph05f5BkiKmpnOVsXPvdWqq5Hc3
Jom03UrBcQ9BWhID8D0j8n+yRHXHsqXj7qvHsgkSeCgsGP41Z+kUc3lJOy8B63H+
mmgiIRbHtjE4YSzqZErWPKr/keJfLtbwVH3+KoJXI47UBvyyOUj6k2amMtSgzWKg
UKw+un7iFPjXZfsWrRdeXBAMm5LBhqOSsnucbrnjMhpGAQryP5ZR+0Vg/RlP9+Xn
yNboGr8T8Mtn6Im4KaFBbFzIItP5rNKAQF/D7mRouoL42UVWqOhAHaGHL5Rqp5/G
+kIuR7RBsw9XOuOWOQuVOwEVJB8CeuicovBWO5y/VLM7Kfg5rgMJ6dsxzCSR00F+
f4rDwQ7pWeTymtV1Xh10o1tmoRRKme/jP0qvjfeTeOBHbYLQX/Mylj/M60yhu0xQ
ubUoDI8x/lyW2oOlqWBD2cN5MjWSYE4wU1yIdamb0GCteoEkr+/4SnhrkwEfiOcf
I4fVIcl/4IfmUk03sB5C1E0jgEumu3Z7lJJwIJkfY/rWsfkK1W9iGm5a82A2iED+
tISy6alO2oJhylzGRKuRdzm+fDFjhWtEuY5i6DatCxuYfjnmvvw6ldAqOC8nK6YW
Znst3pbsEfCf+AUe0BG3BnrcNuO2WnoZBlUJgTTOEc1CY7Awn9NDx+1zuvdE1SmZ
R30KkibOf+2wGmukxLlFdR8PtMUMwAtXJkllCFtEVLaPDCj53M/QyQFYq/M4xaMO
YjsMm8ICIQHpSikcXM2UKcrTb8GDgLB5FTydvdRkraZXcCtaDfY7JTHrYonnBHLy
AJA6B3MNWVIWn8siROeGv5S2wkuLfronyOQzux7pMO5kYLn2rhxsF1BbtP+EEkSx
+WoknXO/Z26m3HEhlIAxlbFx95flUiSY6CQp5yziAncEK2RQ+0RG64JmCf570SEi
0ZM0ISaqHGvJJ8xphFrxEG2Yn7t2R66bxq5r7ZLF+h8J7o+z/gzDKpqOe/fP+O4c
qYjfECpAKRWuXCEHLGX3WP1ScUhSl3L3sw1fUXG4qGElATU0c77l4BtVwip68NJx
e0e/BhibjeIykzbRGScIO2AVCLoUpaXioFc/KqLrW4PrkUcuHPYTaA40xS+vtfuN
1agjI3pb972N67IWKu5fco6bkZQMT15FPn99qBpy7kgPKxFqBl+0pLCYqSPcv1GV
G+2OEF1LXijtKSvjLyJABI0gByH/1TI01yySh7PngDVl1dLFRjMoV4Zt0aN/JcJv
NztOMZWYpODiIJDzhxdrkBhz9wI6ayQgNu+IfljtdktTVsUZJIlO/1trV1+OWEn7
lwQmR9RKl2zDXV25ZQmPlijnzza5xpyJEVM1BWkQ8Zxtb0KBGBW6EUHuR+rnSQlL
GtUGeyoQeOdFY7riqbHWZFtUV0l3ljk2fXNbMOU+zt3+wmWlUnHuqNbbISIQ75OO
OvpF5zrlasemN/pEkSY525yGsXPvoYVFUolzUkNHj1h66b/cBEHIPZvXqnB+qbkc
aAJYyfYYKQqcf/ioHvN4lL9uBoz+A9q+WLxwtE+oZQlBiA9cJB+lQPidrrcQxpVo
qYxt2J5wb/5VdbEk8KRVfZEzyYkJt31pYyaPfbRmk3z98R5HddvrzLTSvfolQYcf
lmzmxHJ4ZC4k9kfxsHLZuYz+etbT0/P855xlR7SPRAYtnOKQMELylpcWY2SzSHgG
8xvycNwBr159ElibgA4FZrHoMigOiStk0ctwmt6yYBRPJuMKxD6Fcd46BSsZBaNp
f5yJo2OGaRAD23daEcPnpeFq6+s6AY7qHD7v5nx58vE=
`protect END_PROTECTED
