`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qPNLHUVKBn/OHgn4A5K6i+46jgYklnRGmxE5phnGBMpUL82pFV6+tg+3x4ZPThk6
7fIrRC2pRLN9G+p4iyfN36M+35YrXILRajbp2goaal6QqlF2LjM+R2SxCR0ZRTuS
4dFMhMWdi1rGCHnfrTBnw8KGfmHMy4kEcxRu7rP5Sg/nMssSNYjdr0mrSzkSxM/L
f5U9SzEbnSkFYgOZPcrChWgFCSYq6e3/NtEFqCgUBE9UIiSdKLfcV+6ugi59ZmxO
bnwRnNDz1WJiuuNNrladgTrgnL6s3C7ayV2dw4c+VI2ae+FA+Jr4+SEe8qNrrvuk
6FyAiDPFi4OaPjgaN2jXNl1uAc2YfkP8gTFTVrhGOfZJRmQGd67PHYwcAE9uWuG+
HFounZLOLz2aXkLPN8PT1kajl8kQtxzntLQTz2G4bwZRBqFtAIuXj1b06iOakl9I
OHuW0jcwgyn45/NvLuPHGpTTbwuH3BzRaqtrDi3PFQ25pY1cL4047Jq5MnomHXdd
DVwuzl2mxYveR7mEiY3n2YDP/1T5aSH43oq8WVOj8RhJMQodtxSdTdn5fpdhO5sN
gWqMgGWvjA/TipNhqrcDTWa+CD9N5SOJiHiXr4srbwrcu+LK/xytDAcxIX9yl9OZ
gbw0EhFqDZBtGVWhxEKxey7Ml6sm2hDrteTe28YRjgWX6ONhNBxGqDr96C+Wv2Ct
HYWVXhtOC23Y7yHgq0HBNae95JtUK2jh3+B2C9hC+XOEonsv7h5ACltj5e9EETB9
kbGNawXpmcK0rHYuoUV0DAz8gvzuCwTJdGCb9UFJxcFV3bHjLpGO9hJdTUl1vkMk
MDLPJQTXJGLkiVWaKDgHTGhzoq+uBXJ5mYpvXfHcGpi965RnuIbCXxTmsyMJtCMB
4V0e+NsH7ITJjmEo/0hTXX29jxHE9yskbDOT8/wMPYubSE7SywJsruIIjgKMGwlv
IMJ2jRT6dlzGwwmGbZJTlOvHspx1/v3LJzLcFdrPiUCbMCXY+FTlUs45yBvjsjRX
cBiCiwdqvRQNne0mA8bKOI43Ii8btqdb+QOCkWeiMpMBAhtKszSzBbzQcWwgvZaQ
U6iJYq51W7l7b2cSkbS3iJqFO+faOnfcDo2cbF+9FE/+1we2hCbWjw+iA27M+tKr
S1HjwwMmiDgtfNra4zaPysfPZ1oap+ojziqlIh6JLO2Fn1E88IjGxe+fKUD0PXpS
vZR6g3vQimQ4+hcYApBq3cdU8ldqP3aHtn0XklyHrRb41xIoNnCX+MS4o7v/0e40
9aKnHGa5XqMLPxBUnGLunUSG5YDYLyOhBAu8LbFCwa85J/EQwvwDgfpG+fkoW9Fu
e87dvIsgUsF9WlW5ylapGENY3jKd/q4D03JKBHqu9u6uGxJgkjQa5ajpxvB7KEof
LC+f1TGmXogZ/fGMXF5GcZ8s9g3i39uHZNjH6mTkaZ5pZU+x0m7RN/OrTXJ7su92
YAsVgf+DkvbES5CfxQlszgN8HYanRh8JFUxAPNazHFKsiVSJkmhdPgmJX38cEd9m
b3V1G0Chr1rM4Uj5WGn1Vg9R1wKTdej1/YfJHmiKKfH5JRyglmYLfktpGE4EHUOv
zcT09gvd5rNZUdwpXEzuDOEKii9FbKFCSMuTuJ5OufupnXQs4z+9umu25OeWeSYp
ftxY/UnOctFa5y4x+UocQW5TQy5mOgOE7X9bpaPPBs/pCR34y2HldpUNX+RwPZs+
WppCwFnP8E2mPhgbW+Fljp0b6D8/ZgAabe75Orh0HNiV/lZDaoBXBZA4AnTNKuAm
PcntMaYaErM23SqV6M+xxD7/fDRqcWdxTY9ihzeT9hpfFeRTNDrZRHoxXwcEUiUN
a/TzVUPpAA9reprU79Dqwc2gEP2iv4JbJ97FT8GSNhJVjsQv7k+z/m33ktIScuoD
N9nXW5sIGRxnHpKX7MnJ8h8sGn8DvouPHI674VeTvQlGLgof45QM/58x7U5cyrnJ
jMOVBts5nnKuwdPJbsjIOZAJ1dAiBhUZvMz5g6NNe1g1Eqo0otK+/WhCo4Xoibgc
3+zpN9VvoAQZF6jxDKL7SVjqniO1b/uUOK5E9wHptwiJ5BOxrcbe5Byu2vexb66X
0oRl8IdiZ55vc9k/lB6Lno/671nyWNYQI6j11mMifTXAFe39QS22qcadj7MXr4vp
2mNvxc0kS70UvMbCzZonwRU9swlH+0z3J3d2ykFOk5RZHACjTUq/7TaLhaoiv5rA
79RmfOgSLWSA5K/aTdpPpwEKv7JrfhNGnA0tzfLjxK/SEtYz2GJ10eyy7qUFDB17
NiArWEYiw/huvsPttV5TwZtTPBsmgzOzmH8v0DpYp2MsJk/lr2ddqJTsbryVF/Oi
WS1Du3X8B71BchW8EvFwpChUkSqHy/QUTZB1Po/Z/7obVyalV0o7DYJ+ZwRWzr1b
7gZbWx687I5strplSN+OPQoRJNc/ncuiCTePqNc9IK6GsYc24tXKSJY6ah0Z97QH
tQMPu32TDeF+oXFZ/f4NxhmF9p8NyxhY4EJKFWJz1EyoGNydlMV4+yxM0oUWb1Pv
Andqa70B8sXv3E/XJxOGOx4dZn497qkaVXqiJzD8lDJQX8QpvFdC+LZ+71MIP4+l
vm3rPeYhphTFr5iOR9M3CeZgWzf7sWA5Ub3DfF3oNKJk8tMSZlAuHpGrypBLitCe
1pij9IVkZNWJXgCQJWTi+U0bboRduzw4l4fggOgI8patTB65I8mftz0bugNWpf5L
ZXr6jilzzfn/WikOJUK/+ijnEgHqPUrATj/MB3SeNxbS/V0LU/HdxnOzWMOX0jYH
+PC8pxuCaL/Lvd/j9hGCrNywaTKl++4fnTG4cvuUZWjpOJtO3oFGlkIQz30Pcamn
FZI8dvrewX2lcBdP3vWLT/LnQCEwpuzK8h6Xp6FzY5iw4cwC3glXFdP42eIDW4H/
vSajhrzxCU4aELy7wCm8k5ro87EVz3am/nBA852u6xKjdRzD1zOKPvV55fMk1kQ/
Cv7f1pWODb8ngcmy60ggAjd/wLxwfwV2eGD54H3eI4Wozuu+FK4wSLFOiG3SOVfU
RCGm/Hkh7WiSQMDFMeMozqPCMpkwDV/pVr5qlbs9xn60qMeYXDT57fyYDtTS8Ybl
tbAx0BtPkxcdqJtkvfonftSz8POCFI1zrV1cWuc01+3anp27+uQKwTx4cJViPKD9
jQNzczvkDbdFwHl/h4iCcJ+eanL62RPyqhI7kd/tyWVMSy80wvuvZRUGg6MlEDqg
gBT6Ao/LJbZKSLXyv00W7EyC84daywCDlkCQF0Xye472oDaEl2HZolLcAPXhBF3H
3IoFPafbQMw14lofGU9WrHs5xLgdGg8RrNkfjrKgF8MFL8iZctwSFVeMoKjnSyT1
sKq7AiPdkWqd+/HQxQEPFRwT/sA4d60WyMG69gFJlK9wqs37a6I4yos/S0ua18S4
H7bHSI0EaUw4LHdGlyz2ImVQGqCaGimheORD7qmPIklmguXLUhKfDUdaNSY+wDLP
iYFM1tajJ3U0NpI8u/0EqOE0VyiNx3hNfYV2LtbeNbOqYI5PkX8cvW82bcfgVrUG
xSWvd+0o+WVBoebca1fIIQ==
`protect END_PROTECTED
