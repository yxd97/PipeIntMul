`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETpMHm2MpHHka7zmQdX4z+awWaK7TN3cIfzT/5DAR1NRnAXW83qaSBltuRSJlVAi
mfwCcUs2XolTG8dqKXBxz6XCYdG4dtc05L5k3tcVjmmIZM3RgJbLqLqP46nW/3A6
zvn54k6bb7V/PKKGVp094OluNjcyBcv5g7Nk9wvEtGKquPukkq8Y302Uw5Ccz9nV
RpDETmHYmXuKQmCq0z8C0V1UqvcvML5iMJu7LKkOENqRr8L51h0XbhNbAeYIa6i9
gaFyqqGR2gOkTiMlripThFZiZLTxBv0Mws/emxUhAki/foTTy6S9EkallgHSn8bh
`protect END_PROTECTED
