`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B13bOavmDlzGok+3t5NxYGUKZDKWiXcPg2gFARy++3qSY0AmJGAjudQIxR6In2vF
pBd2rK9nF5DHFtMwISygqpH0W9K43I1WltTyT/Ij2bdGXHEKJ1iVj1o9Gsed/EZ7
M/3JKIU1B4ZaxK2xmyU6eEauZT/Rkk0nLEDauYERP3yJV+5g8SFnyVIVl4MgJ+27
0aFB96kEH+0Vtiqd+O3lC/8hAtwZtuUuRSFRNbxfgq+JxnjzdG0xumxAN9omF/Op
GlPtvOakZ9n5boPI/XJ7gIFYzhN/LYG03E0aAzY/j4zBpKdmGMLeasVRcFIimFvR
QHwmfpVJtO2h2/k3oZh/i6exWIa1nsfCUKZkG9/EMsbtqFjV4EL1BBylWeea/F0I
IJJdfi0AVve62cLye92k+fAlxxVHKQTZuk6xPm/LvBjGx/Y4MNMMcwJRFsF3Ds9+
7bekVzbCBFtKdqvNOuVPCx3mKrEzFTk79321VeEzTJZbHpftHJkVWVysSimhrwKM
LUuZQkT5vXwdMBuCutqI1ECayBsgn5+uWtp18PIsMWl06W8DUg/r9S3An3TwRcQZ
2Y+yc3gk5f67rvXH1xTMoYsCXnNrh22N8fGcZPjN150DpC6TUhdSNnyl1mwMX5rk
1BuiIVRdWcHjBBHnduvhlnisnhfGA9OdBYsTv96L3eaCRLF31ewSSXnis60uflMJ
GhmUwUrPhy+/vxVbgZHj2WSmG93hSwZPcbhnB2IGKpuFZ9wITqwtgMpVKyI8yqrN
UjTLOIndgHYY7jFBS1xZQmFB+uNLG/F3yQpqoaGMJMucF/4pxEily9USPwV5vMf8
qmEGfBp7BF0DhiM7gW5VR8v55AoRb9pb3sh4OYa0sZg0bS9JoWaRpS7BAKbS3eQr
CuPetYdMTXh4H2XZgkUmrtePTQoCiTWpBYgQUmeFqMcZkvDNQgKYsLHkV40mmp8S
ZeUCHiBFKth+SpwK733M06J9NayztBsyPIGab7BqKC8Z0DzaS9qxEnzfsKmcgtkd
+yIAemvaANhaGwq1/8n4yxJMZWO/7S2+mx11Q+bYah/M70QokNwFAmuODGcJas5M
XnTtaMaUcGQ94dwkQoqfqib1slIH7Q14jNi0lc7820cmfHm1MDmw8tdPqpwA2qWs
d6JuT0xOyX7IHF4eItw/5jH/hzO/XYtVBFPk2dyNl5E3+Vsa7iK0a5z15PYGWdyE
jArpHyp9LHJDP4RFz3whYltm181Ie+UmdiU/XqhaYyKfcNX+leRVkdPZnSNe7Kww
mviNJtJqCTJilA8hpOT+J+XcSziAr4weSmodVxQdGYhFr9IM2ZoX1++Pkm0QdIah
ct+DKqE2NLC2v9E/cKGd8e+pP/a3dKn9H06C4OtsX6c7l0TDgPH41uCKc9+Fmwxu
AklCps3VqrrC9tUvS8AT0QRLxkgWOBIxcqkUxBk3uosCQfijVondUR0+8rM2TPvq
hjy0ZW6cbSrfgVKtTZYrGcwI6MVA0ZqY3RSfdCiqkC5rVnhNbrrqBkusSfzFPNCp
s4jZ99rlvUpaDldPqE5O6VrFTcSt7vWVFlLolwFwyWhnOcErUyYuIQWGIJm4ThJ2
RPvrYgp19JKuKw774f/ApjqwNvp+OtJoLf+07swpQK+J8E4uMd/GYt7l2GeJqDzr
sAFBlelHNqn/UL2bcd0nnQt5lJgaYjDIzbXAbTNvTKgg7ycXf1vxtxbHaaYEQBji
IHUhaMPYM983RmjedEviFEGjos4d1fh/zVhgoc30pIlyV9+DJm9aQ51bUUN6nJ1y
FdTdaYrW+w1YxunMmF/6ACGT4bJe9mrm7WOqSrZ8cTy6XsXP2haUUi6J51gj1XaG
ut2yRHfX4DPbxEwzlp9g04ZhsY096hoKJb7cFpjssjZOIFJ2uQ7T5A3mABAr/+hI
ld26sDjpFW/ip/FKXgIi1FQ/K2Kc2KMy5j1Riq2LAYz/MI6Ee9zeEYZNukK4wABw
fwEKjnGpdf/M8jRozugjuMx5l7y4CGwlJB1trRWpSExu/2fZCgtuhfP7Q9KF0u1B
JIkTl8IupWflPUHu8saXHWnelajyhNOKsoRousdmnJON1q+mqCC7LjGtbP0gJw+R
O5fyUdrAQ5QMX6iFy8KZpy7mXr8ZRS0FJyPZex8FQLTHF0pMRReSEEUc+Np3FQEP
`protect END_PROTECTED
