`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UFk43bgf49NvXmmZlniarsB2vo4w/HlxNlI3SecQh0DouCLN8+ZnZyr6IiogD84o
rPsPLYuLixXRQyxDeh948ZPKEHXcb3/BA7o2B9S+Lx3C4+3hYC+BTQGa0VXp72GF
yfBgSPVZdiiowC2QdhEg5/gL02oBuTy1+FtFIO8ezqNHGb1ENGHZp8BuF0bjj7IR
oKHt3jXb1C4NjLhIxcSABwPCmRvKIu1qlMP6y0TSMouNfONCN/qlSH9LubMlqYzA
E1tRQtb7Rcf/ON/si3DAJTctVtXYbWuvthGin75pAUaUFMGvz2utqJnV9QSnAwmU
w7QoP854N8NBANQb3z6bMKtz0vnAELyt73eJpC5XTCyfIhribhWdVfLS0Bb4oEqF
QU0J8M1h6W3J5I6b+CavWFEB3pSSedlpy7hoPz+Ley8=
`protect END_PROTECTED
