`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
25Ti39FmqH2s3AglOnKE8Ozp4fXbh0fnt46J1cb/KYJmEDav9zByJOIBCFjBNsIN
ASPRc0mnqvliOgGwMUWgt+M+7gRRUuMCrkAZSn+f39QdX6WRl/yG+HeandhT21GR
oPD2nKvxXe8smaEG0OmhbhHKygXPZRw+vBCjVlBkY6Pnk87wtU9S7vs7EtOEcTca
cBOZCHcm6rQ0Seh8s5Foev+ym/9h9KjqyCQ1pvcdDqpuw2N/begUHOYUU0OlG+rG
OIKeaNHfJn0rERUl1LDrVKeaqxCUS+/ynuu5k/Tqi8w=
`protect END_PROTECTED
