`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85zkVw9QEJkTHVvJfXxByXUMjzhE58Etui45b9sVy3OpQ87ae7zsGaTq4bDE6z9+
EgobX2c46ImilL/YSJHxI3/oFCHERdGTGzP4h8bpntjbaLhf2FJX5MEcn+RRB170
la736Ps6nf9jfjMnKAj0er2GE4wjFFXYTBF/tBEjdnWI7+mozADYHE8xSw5spA5q
k7gJ7+j2E/zKngMz50s+rQOLbW13qQEmlRvbKPzoJwyySqb1fGsmUUiKsvc5xs2y
rVTEmEIQrMCEW0x+Uh410e/Wub8a39qRaLZL8V7H2OlcRYu4IbalOMpnyAxxBXoV
Zba4QFdzg3nsi1LZycfRTmONYMQQkBh2xVokcDTqrN+E53R2iUfMnqpzGi6cupyj
q4cRO/x0GygPHuM3zrWqno7tsUTrM5sYFUrg4jXfwbw=
`protect END_PROTECTED
