`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sO/EbWKB/9tFg2a4p8WAW8GO8sPUm0TDP4S6Qs9nIn6hh5FhztjiatM6lymaBivP
HVUDvXLjxhU/eRWZhTSuXzZHuIHb05KI72zO0kjk6Wr3cxehK/54CKsd/Lg5c2cX
2VIcgPUERdEeDEgCxhJvN0Ly7idsJQomOMwZ8ptt0GEM/hn3c4yqxHKmE6km/C47
toK5M01JDeLA5jqCxPVlp4ZqeQWHy9Ce003f6X2Sib8CsrLoqnJt/Ycf9K5UP3VU
X2HEKKgfj8sN2KWbjpX5SKUPH7UHt0yCxEkxM9jgQylDf9vcIMhyWWrpSzBbA0ej
3dTxFX9SWFlLGbmZ0yvUHj555AzJAwhF5CGVRAtx0Pp2Zze8Sn/6UuwRlpvwN945
/Zjh50hUMflzUkyDEexP1EBPHzI64AK6fhVHW0mA0p2acVpPZbKT5jpHI2l6hAgG
6XT8D28IUMLeSYkG9CQDtEQkoXSp9Zhk7zBB9eSJL61TeQd6XTL9SLwu/36xzAJs
IqhEGeFbenwUlNS8Z+dbVBd1NLzlkJy2A2hMPoV0tS7reHCuAiMocgbqpQBD9Jgr
YPRnBVkNYrKMrjKYMplvNPCY/E9+qPCZaw5fJoRMx8YGhnkALMVHc/Q1LRpCWSE1
QZjBYhZJkXBn67aqe5k4L4PhidyX7J3S2TXWj/rqs5TX7g5X2MUYXzZoq9tratuP
vxKkf06IK6VXUr49dkYylyAS9mgZY+06S+hGUuv2kPWDlqOuC9NpFabgs7iG4q5d
aoAtfVRP8Dfp5f/9ng7edcyadIBNdTDkcvdC5gG6ABxj/EKOPAqn/k37r1n8aOHi
yqoj9EKP7emRyWiPJvdcIym9L2AxBqT8P21TLpYRZOjtswEcZbFjSNpBcNbHDPwW
ZVliyJptpEWztl3VJkDIE2XNIu876FjYZNek01FocMdNJPWlR5/H82Xx7ZaqWpSX
oTKYB4ylf0W2DYwHWzHcsSgFcZdQVEudA2CboBB7cks4/KnohgFiLhf4pjl08ohB
85W2FBECUhzT9RSC7g04fFnO89j6t6HJJzuSHsjlWPt8LzW2lNRVSbdL6VfwWB0H
TTN7Uu4GumxT3TFRjROwLfUlfps9Azi4Ud+87VwcNP6sYSpbl/HUEC36TCgMUXa+
GH5N/DItpLPftAsYZHyJAoo9ai7xKfCp0hseMXEKnjZUVqiw29aaONwmudPiCAUm
quOtnZv8/SNRvg4NCH4ZxWSr2RQtRMwmpWZIwS0E2cp7jjjdHmNAf5XYg9Zw9rMF
RCocHT98aJSfGAtRT5FMH6UXTu7whua2MAx9En7psBfvxkJF2TQnII8EExvuhIMK
UPhHu6Dfsb+YDUoty+VuMA1IGrIzYltn4S3iYKtthxWyqNLkItC2j7SG80BGZzGa
xGFoRe6s+m9dYcmHkL2l2WWetDFTlnzjD01MRI9obixzi9FngqoRu7f+sPq/85rq
CvOBp2lpXpydtjuz5aSbKkhht6im0bmTsaWba3+30WE+UtgHTAazJXj3YFbk+6xk
JPh/VfoYebvTJdCXjjEdItkFhl1zAoBdsArXUxG+S/UwmsE4wPMI7nF7ExTjURLY
l8xQNt+t8oB1IKX9HrOvZgSv9uRyAnO08vRGpj7GEKhdpzkQEqo+flW84PSTmRRk
4HqCHa13yuaFikJXfkVaDIpuOWT6S4472f7sZ0Sb4jv8lpFnsM2bCMYWpY+j/QHu
gdY44kRZOzFtrZHs+nrI14tVbbs+K6iWSSgbE+RKzLQrpJfaCahy6LMegu2l3YqG
pDarItKdS6z11i4sHcloek8uMQCzFdaZtlLDslskC5IyevbXwNhYjZb7Zaf9tAwE
6l/YaWPaFtliqunBCEKobtpBUxHzJDpUaQa1wJngkc/XMjnmDlSSDm36t+AQS8Gx
yltepDwPIs0TyUOb9CLVkSG5T/v9wa9B3SZSqiQDjDQ/OZOj3zwHIcnip9gk6KWK
6VbkH+nzebB5rcvSTd9QKes06hXyk/iTZTeloT6LQO57Jpl55+Ut44KowvmENemJ
uQ9j9YJqQZsLRhvFTQyE87G57F5yVFbQeanm0emtiKGmXwvJ11PHubnUj8Femtkr
`protect END_PROTECTED
