`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gEnQDdctDujW/NjxfwJqHOlHGdr7ckJGYEQSnrGBY8u7nUurVobmD8e6kKUxA3xN
t/ZAXK0qMvBfKB297dE+GhwTSiTQ9i30aUtFbuWusIHfplcRwW9fYyQ59gXvDc+S
cjCKfFOA8noVql8focjDIJh9gVO5KK7YZcVDSwAyko8Hu9KivMynLT3PF4AcAbBC
ULZO8qXjwW4VXSxdytYHgUEhHm/Ilo83dn26pHy5MDtdFMs0TklY2uDPj4bAXpBx
wMtBEOV8cg715Zx7yuE1xI+zI0eyEu1jhLvEnv756UtoSKpTUqdsz4AtqreFejMX
J3i9Kv3aKoYPpz2ZilOHTYiENKDtaU9+rwkslxGeQrCOT300QgrtPMaJH5YPAdd9
CL3ew80mFFn4Mu14360chhdJx2+T3/TNvWaBLozLsATVyQGg44UEdMVY93du3YZh
nJvpfsicX13kVsMJIKksnt4JdDyrKIEz+A/hp5ngqQasZWHQ5lSfNF0/QGHMB5b1
6+BJXPyVNxWO+yXw7fUlT5HIWD5k/3qynKWnrceX9V1ybbnWB9E3XOS2qehYn2C0
/8Mo5o9rZL3ApM9Rx6ujOqobFcgIc6JwOhK0zOHBdEUyMGLBVm/0TfmqCacE2stI
jbvxaBkM8gsfy3Li/JTDMzt7CAkGSJI86OpbGy8aWIVk8L1aa/zXay47AmTicM2a
LKklAPIkGY4XugNegs5g7AdMir6uLzW4IVCuMrCMyzZHjz5WNfP6GpbRA7K3n9Ho
VRn0P709r+L4EHCLtJNiNQP7NpEmbUxrgIFRAnuDK1sGh9xg3YzsplWQqIiqYADk
YnXH0X9slujxDiW6rARj3ZMK3UHfAAx8TZ1FHKSgYw4WiVQVycm+HARi1HWEVuYx
GylS/hicSNZmSUggjy2fBIFlDdswc+DIgPuNytwsFrYIZQG805HURLhd9QqdAuVo
7u94qnKFEyAkbe027QBCJ3t+0q3QygRBSWd2ZpYjcC1L0a7VGQbzJdJgjaKwTOMX
pWVOpjtF2oTRmKuuHHiQVMbrqPw5QvP1bObelPE40fPMNTGp6fsfxZIFDFWICA9t
Wm8m7U0BSG4ZrBoNMRDcTvHDXjyPGb2OlIttsGlypNY266MNPuE4JkGle5XuU9aH
512bSsa/8j4lbeWx6YishtiEgACkYvFuP4vZo0wU6QdCNkQBr91w1cpp5KSSbP7G
6VIx5RtPV9I+XhoHPliccYcRovJFcB18WBi20kaNnR98E00QVsmbBAPSXq0TCEn5
6mp08sBLQStdYXEMvr559yWN6Iri1TwDocQGFQM3mkGYucrcBs04tAcl3eBXiAN7
7nQrSc/1J3/T/kA0D/oARNsIYXcaSkRKVf7c88TgJ7T+9WjGaQpfwjeDtH7MSAYr
tQHCaQYw/Md+JJatrKflLhcp9mj1dUWDVtGay1zQRoPo1264UpS4Kw4gLAs9tWE4
Hcd0Fzw79Q5LKF/BWB/FmqN/l0B5Qj7hXwNrKxv55ws3CRY2MipySvxmSaNvZbTp
PiF9Op79oXFV7wqizQAbGcjEqjgFZWOV/QDjombLS70ttyyczLgoFY91x3RLOtLQ
+xy3oo23jRM+dbm3XAamF2At7D7G+VRKUS5vCFH40IwhKpPSOIsdmeYMguBbFt/d
pmRpkzI6JFFYTxFMoc5GQm7E+U+sNjJy+DBlCPUlySI6Chxh+w7cU00YDn61GNCr
Pzt9fqzDvx/7skQsbtaIhUDl2cYTHimtovHv29Pl8secmfCaMneXZo39oo8H9kTn
7t8q0C3XKka7t4RkfD8Cw81PMBbiOdCqCn/86lJs2QKqlP9Nwp+dtsavoapCBr/u
2sOw4LFrQkMFY+cCjrEVqqzgLJwFgH6OfS0ltx7Gw89Tl9yTB4d34eJOjwV0PUk9
JFzAqpt3gYun7Wp+5ZKFDKl7KAsbwGPvq1wQ/Z2yfwHPwE4HfaozTgYTO/FLgQ81
AMU/mZPZQdyFVPe7I0wQtw==
`protect END_PROTECTED
