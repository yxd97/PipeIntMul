`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IujC+qZYGaTcFsiPR8nVClcYBeTZozg9w4K1AJ3QWFYmBdFTlM1pVpztbCtEmml3
DAWNOXKQ2k32E52EorT9LWnLg+RTvUCWUiK/UiMOh7T9R3mLafLat0zARMdPukk5
HAA/KA8Err1r/2N1M0VmsehwkN2e2V7quz/7LDudVyQ9yYJwD7ReEwpQEiThK6Zd
/aKk5H71NNTj+QdDSgPuy+useC6tMaCbpe579G/22eMG8F4IwHSMpDe9HvEs/fbk
DTQlNJDxZOEGnyQLXKr3lQQCQWyB4hUdA364F4Nl6/M977+CWzLaDgZdzKXWYNRK
ikw9UK6eqa0WhyXR357CH4Vhr1+IO4641i7uhol2zj9q4ESHghg9tVBse9r2Ec6b
0uKgB8LQzkb8C0JQAvBInjbD6xhkub1oHd/61fIQqUBUCvlxeOlU1MoEAT2muUI+
UTxAabg0jtAv1yxnyBnv91xHpwo6z5KfTj3R+qyA565FpVKWamij9vH/Fl+G20gw
GORKN5gmRUm3y0lx5sUxgH68BAUejBHzyTPZ9A/VzfUZF8YSw69s3Q0pcpawaUge
2vJBobmH60Ckr0VSoNDdjzGvFsubjzf6E+ZLfh136zHB51z0/ZBqQ9pJFgbwhOvC
6HEt+gOOzlpGHra6QFpy/pjfg2vzXOKDaeJlryQ7qNSU0iwEsf7zSoraR6+K/BlS
f8qHFA2Mb+VeWoA3cnBF9Ak4OOrijPxGdOnJnHT1UCYkKSwUZCaZ3crZPRhxtvRU
2LtBcQBXUSyhH+S9Mdou1/gN9+8mLnaazbhVCtbbun1OpWU67veIm0ZK13XwG0S8
3mY9ZOXerA3yofvnqVU6+4dwjpt+MMVmDglpBKHR9nakuE3w38Wb2uLOyL14Yzdg
dqTpHo64+PqzMiA5+cZuL8wyc9YpE4J4AGGpF+NV7j5CU008zboEQ/+18LA0Y06R
/ID/zcOvIMnHU5czx7q2QL1uJvfXwHgcgfL7UT0rJPxKkE3C2j/DAAAW0eHVqTCS
wkwmVnmchKgz37f1fAVPwlqQ3y1QwXw/3jYq9CwXrhWNxh0933deMR4MCnkNXlDo
RiF9orpm9YuJq1tShVfP0iCkm+kFIrfqFev2jqD+QVF6AbfUgReVD1lz8hwouHum
BUu9HD4JppKesmS5126gYNTNT3DqTr21iKEC1Eb6FmFhe71BC1xpiRpOqCxJcqcV
C8HM3Swhof/GR0onskYuOaVkNeBepeGEP+r4bzPRCqLmMf9oMz88gWJBgOJOeNyf
xckl96wqdZS5QDV1NPQYGK3TEpGSXo6pD4o0Xf21d/BGjWKFQP9SHEgOjo2N2j8V
aePHScK2+F9CFx7dIMIfoV3FNP5DNWLMZmJcf2GEP2yp5I7SkMZi2ql8Aat7N5df
/WdF8ghZv4C41i6ZrcfX2XCMk2Vm9ia6Wt2cfRCfML2ppqC0HN8+bQknBmUofFf7
fcHEHISAPWYRfwZLvY4ELEY1kTCOB3X0lEdhaBO2kMEHdafYX14wCgxcDVbFHgCm
6GfZv12wHTiq7SYHLdxM3+yUvbeDsH7mcTI2S/hqIn6bJita1ef3VXs9ObgFYDKq
Boq3vw4PS2q5/9lVXIKhzX83ycZSzwXy9So/Ft4XWlm8nKFywLSXA2ZaBS/b7PON
U1un105NDYYeHwAJQJdN+GXDMXJVcY5dss8f+XgrcBPrVd1R+MM7J1Icw1SPk+uk
6Llwf32S3Dzqq9QON1gxHXmQNCBkg4xLdIK/iYwGe/+5pxvB9gO+xY/a30wzeM9K
22h50bgdRcjJCUpbc8E4Lln1OoRSl6Isu/01FG0OZOEpA560RwyCSTrmrku7pElI
9jLTiHC8jihZcQ0ygIuG0HyNPMtcBqnG/HQh1/Ndrj38+WcnTMtfVOGeWyk+atG+
4gHyrAa9JC92gFqn14kYwjyNoFHNitPvdU02x8l/vBbcBG0mq0Q5/AVF4qO3NbMo
2P+pHomNFOfcXwZD68HrnmjVvTtFPRzEkYk6cToF6XZoxCS0aqy9dLc07ikuuRJd
6eRn5UQNPT7Vr9JVNytA/CucFFu2KAyWlaAiQP+NjDPFiWt53JEBNQpvRP9POdEB
eo6xXJY5+c2PuSjCwTYU+RIaGvlFSemu49ax9B8BOWeI5/CjPgAOBaXg/Tji0Yob
GQHp9j9EVNvFkhc9acArhy/yqoN0goToSVUZCDAHyDOHdIsX9eA21NPrz/Ok0qYR
Ad2pTIR0w0Mk10ItsiBPHwrzld7exBMyZyGYCPWGGakbpd/EyzZj2A7xw8gvT3x+
Ke2dv3ALUaEPsfJtieeXX5MxGv9O/6zmv8KnXnn/ivkD85F7zF5OmmdZYK//Fymk
jcwJwxNW5QYalkV390l4y5du2T7sxl/01TIPl5P6Cuk4NtOXiF6u7Jm4RD8ehZn2
GpBkBHW7SMEZIYf5iHlfhP5MTz3HWRsCQr0yn7LXeegvwft7bAmRWCVdJJ3CJ9YS
kAOEz+EQMuK1GPymO4ovFiS/7Gmno609V+xQIZIORp0+tDk0HFcMObXUtqBa7Oxn
Jg23sU2hNtqCl0IjVkHy1Jds0we/aEg/HUGSdTaY0AYcHfSMn1i4NcpzS05A0cja
5QRdHXLkDXFCwq958OGb/9XAxWx/phtkQoGhuN+zDx7+pCV5Y8aM1BHHDTNCza76
a4b8nggEG3v+3+purVg8msWzBtslJgP7r8SR4g/DIMIZIuz1eNJ30ueQHQcpT5xe
dl1LlO4JFFebpjuqJd10AU9BJjk3q+dVnVoHSvQ8sfWU5+A73WgeO9N7PrZ7/sdW
2krK/RXzbAN3fUDh5CWLOsxeLiNhuvkC14v/LOQ2z/Geb+XGxruhRidDUM+FT1qB
mfgdUzCOx5SqxnK4GMEk0ly7mohdCuEbIXPj1jQqNU3NxT0YeEJeAy4dGqshEj4Q
Tkw1Ee0nTYb6YvOlY0HHjOmEJgyj2nk1cwXMyfkIi01jHtZk9MYRKr4nTwJA6R2N
iA5ebqS3yXHDOhtdhDCEIsg6ez8+4+QqJ2c1OoIskTLkQyIbJogOSOr7ChYRBBAw
s2YgKLZO4ygbAvQ8exGNcH7gmqJ4rdvlDwD4qkNsG+5NmHfqy1qqo2yVcRXnGV65
kS+I79Uu1AaeOFO1fXPLU23NTqA+qaxjMh1PiytDONMo4opQQL1n7eDN1zI0AvfA
lKkTKBr3n15Nzxrobq62vDjNy5QNRNZco99JV5LwTOEis0nE1Zt8vi+zE3LcZ0A1
hqghk7f/xWhmPvRbw3wvM1Sl7aWWh4SGQtauAwP67VcGELmf23vaHytlTd5cI8/i
ybort14ux96JGc6lGu9vEVdj9KG+A0q9kR+BviQ26IUapFNC1VDWrB26v3br1vFJ
UmgMgFnw5kWUzcodf3DwgmmSCwvdh7iwXoSTaDfA2PLcj03BbMfHrebwsRI5Lk4x
Os3bQ8MR0/CJkrQlzPjZnpxbXD0sbfavkajXszff01Va0Zi2AVKNq9MF50BHiK8+
wfakjvucBfDXaW6uVKbZSOzZiYiCyGAZMLHQHafQWhGLSVGTgwEPxKRNE2Jqc8q0
4Apa8uif2mA6iSIBTChpOs6gZYSf2DfTCXdeoXuzsJg=
`protect END_PROTECTED
