`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C6o5iivbnYRhzJBgQdUe7/bpVIcsPo8sH1hJ0A2z+EJPxGPEEkQUYnwov1MUIppN
my3JMHjCMeIRjFc0H/MVen1hG78oLuzSu98MQ4mooqEvWXld9wbOfycWA5eBHG+f
soZW6zC1lvlx9TM4H0BwILEeo9oe5UnlrCkbea0DqLKsKoETV4DU/St8bkHYabG8
K3q2d49a9n9vFyGk/gwRdTjQElFsqehy13yEkQ+XX0wifkG64EpB+Qvgtiil+Crc
7pYTUM03ErHUEOtfsgjWUYyWCfRpxRMDUxltkncOlyN1Ias76TWQyjL2iRBS1qiP
wpO4rKG8eZJ+GUWzBxfK9SQAkX+tGvescfV5Rac1UPhGdxeyAPNryWA5PTFQwOL5
bWY0xBbhyThifaGL5RgIPUcC4SzJxvPYyn1uiYBANPCzJjOFuhQmzsZy+O9IuL7H
HFWkN5B8DVLNPHw1A8lN9MiDojczhY6LEwyb8sx4p6EJ0FvRqQyiLiaPExBkWjop
iBSrBOlAUgIe4O4jT6w4M+5p5WaT7SNDP0AoyFamHiYYuOUBcviaECqt/+ggOA6H
QUBElslDGTnxNxeI2uNeAWDUWvYR18vQOKKGm26e/2AjlQOwyG0ZK4IwBTRYPRPs
wPC09Fd/ts1okFjNTIdny3EebYRFS8dXVY3annj/QOgRWRGzGU64qC/shNFGERVr
W2wHdGM25pXYXU0cSYbkTRzAFR46MEyp1mVuSmen0+ArKMGcv83cT9ht3yONqk/D
WI7BIBh+nKiGZPuSA2/8DZ/QKyEc5ympcGF6eHHUGu6H1GMHDDStNkN2JwsqTcDm
ZfEpZ/i+ocE7CYjX9QZQ4qfIR6RDA+zzmkrwMKmG2MA4glsOIK44ibeutyekG2k+
FkbwHV78pSaybYMQGP/HyMF0Sc20fe1T9wXjuZ+qIFlr9CcUtVMy2sJXb3HfS5nz
76yRWm0mwTabgcs3eJEZzDyF7qJ9IyDybHrOHThX1/0nsiNGkxkVOPfQ/m6XNtJ5
DtjFzN+jhImctGRM6pTYfl95lJBwPewsVO5a0FAZrCRlYypElylcQeQI+r3YqZIJ
S1zYtjG4KHTxkTl5wI2yFlqXm3CpwVVWZ3oa2TVsZrA/6plZre8SyoZyHSk2GtV6
C7bIMsbCXwmpQzRGGGRixeV70avBQg1FlOE1IPEJbYlJwN1U8auvuw3L+usrH014
KKXXk4LqSoyztnUUTyXtW65bypELQEjsgVjU9El50vC+A8Ha4DvAFS/+eXVg4U8F
ixy/zgzY+Fs+Zt3GZJZeOdm7Dqwyw59tXgKt0wBIdo5GMhAWs6sp7JZrh5O8SksO
L5DGs1fZ8PRAqsfh69MoeU6gflO9CBPPiDqoBrl0PIelTm0rMsmk5pCLU8/G9Kox
XgGkrMVX5UwanvA0DRSmqNEcLKA1pLAskZV1jbwttZq/15/P1xMdEnUFDZme8hB+
k+Rscl+kIUzif3qkeEagaYXtPURE1NzEEALVcHjtmw3CnaLZMT27m74STAzjoHzE
IlE2yQ25pTy5oks/Ir/4Fjqh/ghd+GTmwjaZQwO9FnkLa21y7hjHR7W1r3CI6myt
0KPTfRYLNXBoIqKw26NTA1ksbhrNcDb/qgbT3VuiUVrP2rIOQBHX3FJMAFe7ofTp
P0ky7WTE1Q53J8cCmRBLCFOs2D8jET9lR1Nl/gMWCPJdBYzRaq3kvj4yR5MhFL/k
MEStPSZGmVr0fKySn0xiRulG8oSjTYkJDmirCtmnQkg/mbmZnx6uf10hfPvDWCq0
3tr6vHakDMynbH3diWWl/ddzxUDypil63HcCBEbcOzZ9ygwdrCqLzfkhxqUW0s7m
Hsxb3JrdofrWzFxB+gYMeo4lDbU+7b21Ig+gTvUodbRV/Bh+wDKRcf33VFOpwCM3
2hjwbuuclTV5+xk/OMOh2Hfy4FV/JH/FLvFoiYwXss3qNEcpA8M7I8whi3X5CvhC
LpF4AuAa0EWa5xiXHEXacad9K0dcihi/qtPiQByiGCmwxAqhFDhrOlUziByA2fap
`protect END_PROTECTED
