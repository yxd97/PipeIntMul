`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OO0LuqJLsDFakcKuOIE2LSMegGElOZGo9grguE1MPAdZkq9jSgdpkgiVtRS6lW+I
FI3RKeO9WEdOiibsSKfSruDgqhe2b2drubugQyfLxyocyvKRcTXwan2u63u1scJT
uM+Ets5/LtFcWMFpZ+bZ/b3rXcUJIfbb6CiX+hRHc8WPajjx57lA/fQFZBodGzCq
P7jSpyMJOFc0AOKkQiR6Q2UNhDT4Inrb1HpSK6vuS54ZIyg0g/q6Zii5Au5EUx1/
o/itrTGjKCXSFAjCMNuxJobzP5To4OwBa0cAEIW+lSyX7s62ibHgHnR6W9v0i0DG
hQtdEBFMTKisy1NjnNh/wh+dtAOMX4oQVeAbFeW5rfzqaotxhVwp9ueABwduYdcp
ZSPrBPKyhP68lAZY2feLHR+3lJyPIPAxRmQPzMVqNt5vUIWGVhkygzsAlihfWa5A
v52FPGHFv/3cqdVqKyWzG1hpwIEhRLTqKR4rNx8F0+0yzczivjHQ99IraIImm+zl
`protect END_PROTECTED
