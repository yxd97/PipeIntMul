`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YxA7f8QlqvY6NjF0sC7btNa7YQrviSt11Gpz/VJ7m6cXIfm1j7zpfQEue2zu+sPz
f4fgHxbjLCVLrpIxo3bBZpiaSA06dShPMHbJ+FcXniuxD3mH93ZJE6ntrAF7a3OL
hJ9qOvNxHOeYCKsVs1JhJsjUIOh2a/LCMUs/hMx0/JVf3d6n3DQDvo8aBTKToNtI
fzQFvSH+vw879ZJQLKqMXjxlXUZhofNc8AWPKk4G1YSNn6GPMbbjC6WRDBPIqPnE
ZmdrBRx97zHetupJw7PkDg==
`protect END_PROTECTED
