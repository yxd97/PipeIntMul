`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/rLIt2TsffCJWZKUAuB/sD7+BhX2cAs6Y53pvHM4Uv0kFcYl2p1+XCfRUCy/9D2I
OD/pXpAeCtQ5oX0PNCzQK396Vasmwb0xBV103r2b6XV680Hfc2yu8jZ8u0xauSw3
WeSpZlRdqCBWCmTz7255Qyvn8DcoLbo7dyYW02NHz8PaGbotrbsUzfOd8fS2A0nO
IHv3hoCjIT3pyAEPFAEDN7FESw6XzOP76X0iGL9tw0G75ya2t3qD/tW7MNLxD+4Z
q/GRl8gh0nfZumkuPJN6+Gm81oAxTmGyGa/K+ZBAMAuvANxRmoGu2FCGseHb9dgR
ohXv7GUUr8qcPCatgaSNNg==
`protect END_PROTECTED
