`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MeDZfhhKL+PsySg0slR3gL1YXkCIR1mntnT7pCssvpZ0nGGjZebg5HtN2F3vTG0U
MIRTrVy2GdJDK7s6+PoGYkNQHB/eLwfGmfJpRrc1umyiDjcceD2Un08Zn1FFH1Md
leWd83qcjooq7Q/zdGew3A5IMIFy6QYOV9aHh4JRASiJuv1KdRFZAtDbrGtzxFpa
dYQfceOmZ2Nxxu68ivvixK2q/dpI6W5eHfouMGVOrEQJy4IFGFvM7T2GV5l2S5j5
SzMW675IMedEiKzKfryPUo3xioWGKl6E1Z8USr4gw8p/osStceqAt8zQ+N3zMFr5
zUfX/t/3ixIbgqcXwlluzg==
`protect END_PROTECTED
