`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
axFaI/XP1re5x7OYI1QS58lpZZGTg/utm/17mrltIXa17u6aE1MIDJPxjEVNi3TO
uYioqmy7PD+MlCHlDLTlxCLUbICsf8itcKq9uWzlQ4Xhui5QoetToDx1uqAIemMo
tbYoPwctXMOc0DpdoIJqWpz2B1yzsPdolZ8hGrZg3ibvUKmDjC8WdOU90q6dt28N
oigoCo1xBnt4W3rkZCmTmTppqunpgBRpskFWuX8rTaKHQO4sRiju8QmkqlrQBMYB
NYJXegeN1wHus8zx3OxK9RGEMEwJ3OqMKWwqrEBvShgeAUMJtjfc5N67ttsHWDJr
et/2UW2CorOfMFgxGWPOw2Sk6nmAwZzyVs33zm0U0VLVYNGLpz7RBly/3HYkOp+w
7G3kAMmxZeo6p852uD952aMn1vBQYS0u8G2ZF2rOjprIPArUbo3p+Zad+/B0Y+Mk
fBZVVANfwGHEOuAUvP1ku2ZgzBf6dnK3Dcytn6NjXqaEdyUTKbZ52rWa3/S/LscQ
7Dgk+vgMI+UIxx3csEwbrBkvoCGBnktaGULDzyfKbXeOPEDQR02ub6WndWWmZWjI
0dt3BoTww4gbDspTLl/FQRGfP3I2q7DtC8kxjNB3rXZOuIR3YEyRup4gYy0wNBhB
N1UkfadOtdE6VQzJ+xld98/T1BcIL7eAtEJp2O9mBv9+0XycYb+8jPz7GZZbKIU3
DXwDd+FL8LaGW/t7Ub5O0ddKQtU3Y6A6XgicejEyWQB0jwxHP0riYBoYT7JL3VPT
UzZNezZVfy/5bJTMSxpmYcHNyxrj9F5maTTbcL8B0Xnw6mA/ZV4rV7aT5UBTAswV
vEM/Hd+OUGPZJq+pp3OFmgJzEubDLxue3aAPtivasWFMCjXh93uBeyKG8kWCfY19
6G5wG+XAFYUar0jpGkBMtr7ebgbT7p7lvFRWmFlKGnDtf2P9MngGgFS409EKd92y
`protect END_PROTECTED
