`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NM3A5NDqef3bMBsOU0oMqzKXxP86AaHqo+3vtn+F9AHI40hbBNj1snRE00s0Ybnh
nR3qI60w4Q/IeXbh27G1ZzFciE6sQdXHqd08Ts9AMh/fZV7D8wgSKF1fAg4UxqNK
XWYr/OVeUmItfVMaUrXxZUPzIVPV4gN8b0CHDyLRjaWrOVobbcK0Z1FuCycRftT1
NKCuyPeH/rby05seCD6w6Wt0ic4R7K7j5EWsU+/0RJXjNMfLhInaWPvRJDi0irKd
Qb7Y5bljRx186T7Qs0eElSU8zxaw+SKaGoFG7ZEUPFRbWsHXNkpUMpDOwcgiUfHp
o0fjLndNF/mFLEL7ppVD0KB1ckK0SyDkQpMjds0agmnvKnGVqOFJF8ScKZpq0XDK
RxxzTvAO0GT2dkqkskLkkvd2rwF9WvzBF687D7GhyWdNTsz2Zc/jIkAXlSqMUfnE
7VarZYZ4kq+NTpwIjnVnf25TPZ9j9vGto+Dp/Aw0czKnp+NaqRu2gz3TITkMltA+
K7v/P0B1Fsyijru6RpeiDJE2in4i27fKbHb74MnhGOF9lQSLpGWj8mTxJGB4hhXY
q8fZyPb6zNg7HMmFjt41yfD5hBBHujy1PWzkAI6YHrLOF85TonbZvu7Nj7rIUPHZ
evUYP63GmkubWh11/5iUdPUxb1ZpkntRDRH5sBm0cGymDQkpa9/qYax3Q1mF/7+X
VsJSxPRPnV8DywYDdgx8aw==
`protect END_PROTECTED
