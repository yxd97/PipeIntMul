`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WH+3M//Wcwmrr1buM8X873ZQET2CYrTs81T1AHxTk40ThlO0m4/l7/E80a8aau9X
7u58zt+H0DyqOfO2VFSXksgQpzYHHxssduDMM2wD0tsde1KujJ2rSSCkwac+KUC3
UY4Vvq/1zgc4ZxW77OU8HiA7au3SEnGyb2rGH7j+JV/Xs/3SMIESfi7rmBHjXzAF
DHA3pzh2QAYm7O9HOX+hl5eiULv76jWgc/83BzRocTSkNlItnkdN6ITyEER3MmgP
CYzsK3b6ldgIzZEC7C1UIPqzbV39l/ncUyPxjgjJGVO4J72IJvZTzLJqdw4R09qq
qK98rfTo0VIaa+rwoAXt8bP0/ULMns2NQJ0G/GXTWqitnncVHkN3Yomybgnr7yhZ
FlUv489yVOzPtd5u/7XdBK9WwFVPhdiqFDkn23y+xJbPYmx9nJSy9Ke4eWhn4r5z
32aXCNrieh6OrINQDCWVlGN53PIu8+CZRjOmNpd9uCs9v22JYMt4JWDXDHwCrhOT
EwslM335PqKAdcgUUfMz5lymftY8qVWB90+ASrvwhw98hsC/eVnUPkYdCWFP3s3O
grsNo05WeifNmXwLayCekJDFqseJ09qiCxUwLA9UhJChAh3+Bgvy13Eec76VDyyL
exxD+BHL0xReGf7tpRpaUL+lUxkhemVcokbi/2JCWrkF/y14KWekHEHHqKQnht0C
Bdop6sHXT7ssOq9scW7HhRFI5Hdpq8LoSK/7htWAcU0=
`protect END_PROTECTED
