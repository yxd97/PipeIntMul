`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
++BWE6yfLxrd/q9MIkJtSDGR1zHfNghc4VkzcXHC9Bfj6UcVXrKvqtqwaVf2S1xx
UTvZYbL6MmC7HRnkQAjasJJpk+OY1UK0R5vYe5OtoUD6Sc+hZhpuvbl2zxN6BsaP
aEs9gzo9XOVYCQde1DWNtI/WLvAbN2VJQs0PT6FHgP8Te11YDyQXcM+NiDR9jEaB
NtFken2PTX2kjB3wkAncW18iLu6GoI51dr/E8bZM4kR3OW32SyjdRaCqV9xs6gk6
cGkYIdWhgIHv5f9Xwgz92OVpXt53DqHerOAmHzzycjiRukLPnI3ZdTzARTTFn+WL
ah6R1WhRYkn2/daXuUdT1A==
`protect END_PROTECTED
