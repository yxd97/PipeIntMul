`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Qu0nqeoAAW4F7go8JAaMtNTB6dF2kxrhnzrgs70Twg2fKBsZhHydSO4lobBmG5f
ka2hpmL+gDRFWAm5t0FKYND2uGQOxFk6sxsuNWrrOXGPFPKVud0ic1Md/C0kEmeD
RlKRZ94bdnG5jUekwdw6qz/JMk8HUcVlgq/+E93Sa4ZkxV3562XDYy3HpQPHu+bq
wcutae1/PQRcBTkFTkJW4ENy1i3IhC3vl2MFRvwPbJMg2KnqudoxXZGgaNB2M7sV
GFBaxulAhiOn/h84BQH6Qi+HlIdHlFXeDmFI27P5y++aRLLPboIBt58jRBCms+DG
YkL9h0UnbhJSu+YhFj+S+rBSHWFxAafgXg4wEUznZfMFcXEUyB2PROcFYUaLVfd1
gGEI2Icxa3lS1/+xqy02ZDspFuVcv+Gs3ksh7FDFu/9CAhKoThOn1KBS91NoGRgV
H1rlqhbvaVtrRw4NJCQI7Ubvem6FpFzxHiO5y9TlWxWTrd0mKv9HLqpTcHicpBPP
COs33EM4zh+DAP7xbifrGgPQm1WPi58M9/qX7prAPeQkGC8aGS4gCHn7A3cMwTiz
2UYVApjodEQfYWLKrCHPHhJxQe6o77vYjk5v+TyRxr5UGIbu3cERjBSspmdFzVi/
4vbbvQllXIhryDLnV8ZOQIpD0gqh6Xxev3MeN4R5sYooDLXaEFkHw0JfpBPvSutL
p/g5pFI1RvIjbO6Q5MXNvmW0OnJjBCh1l1t5pQS/6BrxWnix3NpTLcTRPtBSC+Xk
M+BCEe8xyVayJtVLbyNSL3lxGFhDUhXV5/SXVrcA729DebFnn6EmrPUd0KoNCe5/
1ZuWD5cVThTwDyRJ/G9WZDwbmz2+0N5ZHcqvnkoQPcPWyacUoy2EmVfDMpK9qqiC
rwJ7VjVXFD5PbVkPb3IUzJiLRqyCOTTmQ2PLIizZqLVk0lfLm9GJABGjXtPSujv/
ck8Q8ZrmnGKjWFNCnYf6E374AnvIlVUHQQzjlFQgcLhMCCRG16sL5ysGCJXSgDOu
M3XcooSe2qxm76DS6m93Dr3iIssP6kD8vIWtKyE6LE1lLusD3CYz83eFMWeXZFBf
pnkE6vAPtQf14dPSRB+oNwbxkr3T1WlE7OHRBiSPZ902DIfqvBYDw4KZRjuy4Lkt
Nt+qcgvPJK4beCgBcI1c/J7EdfFobe6vVY3DtIO999EOco89JaA+efJVqzGqPfX/
wIbkTVQMaMcVcU1B0QDoKiVQG1xPjCHld0PyNAX07TBsOWX8RnGsvSLQzoCSYFD8
4oBgRh6JfAiKByNyjjBzk702F7q+LLqj1OjBDoXJfVF0Msp4xR+XkIq+30oHWgxE
ppLesGhzxGPpTkwO75eZWvNpMeeMKP+cAXM3cRj/wr3w+FRGr1CJ/kDV261ihdXW
rJB1H8yiMm3tzH5Du0ugXiJMshILRiFdjnmi3K9KYG9U8R619/nwWkttEtBEzWVs
/qkv2XAd7zyh0X/eSvtOiK/tOYQuW+AFBtMsNFXOHF1ysnT1BcPE7WaEGZMQnNrG
HPWQxoSlqlLLdo9+2FKYy3D5d6KiObMcAH0iwTQHU+HRj8FuYpMg9xw9B5sQbrvf
`protect END_PROTECTED
