`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1x8a3f+FdLKpzWjhJ8himv6ymdFpOE9T3ijiPBm3NIRO2jN2nukqJzR/7px1NvO8
eE4ocOYNqn60xjGAVEcoBmwhV09clHr5+S/JDz1PXePPtvQ65PSMSTl+AVm/tWyD
1F++LZLdSsHTcQaT7XgTpHCZyMpUeZ4CONkaw1AenKWmt1bNAgL9HJkgtA3DqhL6
4kufvwIeTuDXyHLCt7eo2LgEKUzF1yWusOghJpURS4fiUvsZ0qVlu5589sKFg1JF
skjUTtgWsViDSGET0d58DDUcC2QqCoYVl8Q/fvqoAvdhngp9uAqm93d4wm6o2ypW
vDFOZhBoYVIGzZ/qodbO+g==
`protect END_PROTECTED
