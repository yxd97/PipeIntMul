`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rXepmJ0CmNlDJD8PCyTkTwgyAsU/5wQM0n61TmsQh03Fr7lzJOPm+3FjfS3I2CnI
lHeIShbsSzPr0ttzatzWaAQwf1dJE/W+3z06+NvRUZ7wMv7FGtjhi+1pENJ1qof/
ZIztiWPNM8FzSUYCyzukurFujY0cZ24fF9Hq+lLYwDOhi+Ul2tNC9jWkeoaksZZb
DJGi8rzfyax14lLLyYvpvLA02nDPbY4nWqNtEYeII8jDADVJR1BnG4SaidyIeFGf
D0a0aHbrmXAlr0v/UIQf57MAh8XgQpkMEcvKQwWi8477ejt12NxjAsm65bJF+nKZ
z/saHkBoJH1Y+s+NPnKOUtlbI9kiBWLyQM5S43mu22eMAn1V4uYDzisvHVhend2U
p/EeAgCuV7FOPVJ6BI5d9BhKWhdVUX+yI7NIY6rQov1PM62WAQezUjj+0ncKykpn
SduucBGPtn/JpYCn1x3FTI5VcAGJbEgxJ7fkxlxGOccKYrXam46b0YZZFzjSBZJX
5U6OTgvjmmIJmUCQrkbPzpKaFkJsQui5y/T5bl+IYFiLGWI0/y6+z6SWU8hZDT6e
bJ2vPdCyoZ8pbwOD8irdLdbSwjAzMCNIJAkBJxelu1V6jLNSJnkcddR9le6jimCu
2P6aD2COQeF1oTtFtZSoS94qHAytAwJx+mgoTJsBWLltHcN5p4RFoHjDu6nhIRRV
yAeBhEcM52s8suaUq/zER2y/03ndpQKOt7FYb2lzO9QL2dZz2a3/km40ZHqR3Rz/
t0+pnGCFau1pNxhE6fOkCYBIZSMycU0uNayybU0axMSei5WUs0d4okc5BMgEGspQ
`protect END_PROTECTED
