`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RDqPEvnTqn+jW/Nek/kHmmkv8mc01xV19uM05owpMo9UaCO13+Jy98hCAOs5yQJX
Pp3NUQ4KL1NtkuIfuJxbT229PuBfZvEnmtSeJ7UFfHn53ReOKq+reHqomN/ILvCR
twQtZEdyPgEMZ58vj6gf0LG3ShvTPEtxzHHklwR/vUqZ7EIQ9DESieudKs3klF6V
4xAn07v2FIN/7P14ihBa6tZOhzSIp5nQfNh1bpd/FwEILkvOMaxfOkf/fsr1wAv2
aQIZSm9DT989VUEhM6FgCG2thS9OLlq3lO3Jox1MTFofVGUt2q+skl9KHgK6ZLIH
eSbKQiL2w0rKQBWuQfTHi4lULCFxSEiwftp6ppvJuWhFlwwvIJADQwEhiJaVZyKP
`protect END_PROTECTED
