`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3zR7knIIXrMASZDH1sW2V8OJZbxPnNP2HKanps1pTn517IFMBElF570zDO5+1tpu
5hkn+VW+YKHWyocmelM3Le9mAZ4GKItIPzDvOaS6lgwgOlFU1fkstQ58YuFXQjYR
lWwccVGh2HdTNIXK5z5X+VGr6hCSRIYFtHN5T9AwRi1Z1kxEwMMoZSs9/YYZhPV3
5RAgdthN3Jd/2VBjv10+0wNTNKS5Pu7p8AFv8qI2SwhPb/Q8jmclIuxPiy1hLdXG
Q76xHVE3QCEfFj8o21PqopG/O2RkG3Pz+D1zqg+4g0c8qkovLwJ9AP0q+ZBiQnAG
1JK1x2CY9jquCeelVpOWLKApwWS9rKHspsVg00vZThmx+2XJtgEzsc3u9s1fdkix
YdWSzgtZD+PoK+zWivXjoPGAPbFLMZpwI+TlsqdG2oshElrS+3dJdZ61FxtK3yWD
otZOxZuEaXA90TRk/VBl/9kPDuU4OPkCVHAq/xjub4sucmeQ06laGWpfOeGL88ma
QJxtm6mek+IJygdHqHRhGZYuQBMi3GolC5p9Yj5PJfJUJaUcFRCFm7I1IVB9bcrc
cbs/cXCFuAJjhkgjx3nRCaeRkl/fbZSpTcqOyyMfCyyXGuJJW6jacpeghZrG6rAw
x+O22xAE/vnCJJ9JpIoBerNl5lz864TLcMJ5kk20OpjLxUQ6FJgVBIfkB3wSH2Hb
iZYh9wgX1mdC4yJpP6SeiLg1T0v+wPrECPYKkCbuo8nL64EHz561FEau8NdvtiPh
lLtga0PtUN+TKE3WxvSk79B446YA8z+knBSHq0ovR6dLBCWVA5wJ+1KuFFFPoUCI
fewM3jaDLoVseHY8t088l1A1xldKsouLa6CkTRErX5+jyD1l4PIsHzgcmy2UD9BA
nXaFpii0Xp+lIuHDLzKK/+ALSaP2hqtLqYo+vHP1vMAmmVRo/3dUf6289qNE+CbL
iQ86d4gMgGlCrXTj31590eneJ8lK7dduey8mBwnTyKg7H1fWidDUKDGH/VWFm1JK
jAQ2IVH13C7csz5F6BqJpd+WIrWY14KXQyk7dlrosVo+src/wJkRVKWUehCMaQUq
CmocSxaMKJIq1DVn8W9mymjQs1KWHDyKX3J2tgIE5F/FH1xt6MAGxGkx715+Sgkr
i6niGBojMMMf+KNcZ8VwBn8+9yUs1M5xpBcCUBkzhKz4CfsdBrLTQB1TXOQKCm+e
huFqqgQvu/NhkCP82m1elpZISJWlh/ZNN6IbZ4Mi8lLijACrNOVfgL+4WFZCnyMh
d2VsmiGy2TGGpeX6GXfUyKzQQa0uj1Yx3egBZRWoameArdb7xUCkzCyk/LLiE4O/
VB168uVwCXJrWS93s3Ojd72sWzBGvWteW10fdoaeZaEnTMwEUuXDF/Yj/OHBHULP
rJNnJEqrqc50ATu/t7wC8+mr+UGlpHuhOAbq/0/VG/tfjER0jqTFHOPnd6dvTiln
TgDTiJiu7og9XYcDoksGoDC0JMFqA7zEi4KCJmOYZZNsOIlStOLL2zjWMjGzrYSo
cucLG58z2O2KaVV11tQjxSsDwxmdE58ALV/cmkMXpZWmcXYrm+FcsNgC9s/ip9Yy
VLKoJ4zsHj0hJxqWCvcRmKqabzRWHOW+BlTj6HUJvkv4OHpL5tAdp7iD0WuNE7lA
32iL4dTbVDFVwLkFCQ9vInVooxKHuIoJt4yzMstzmaFT0PVkx21aAt73Cj4+9Tut
no9GlnNWAx8DOExkup+tAU3Db/UP+cZWQzzEoZGlWRjyLJSePzOc5AKKjuKFiUYz
MqHghVFkLbTGrgoj7N4aJmE4zvuQdzqDMs7j8eYqmfWRhN58GVYql28FElVho6gL
`protect END_PROTECTED
