`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5n0TFgEF7E2VcAOzr/GDglZBM7fhsD2QXeNK1qMWWMmIJlG/4sClbj0I9YUpLzz7
QEPGibc4Yx8EEC1wY0KNg44Z21fLB7E/zSgGKNyEl9mU8bM1ekasJ5dEEzMg1znO
UjY3XG5NuJfwsHG8lNBE2hvRt+vBVceiPojMLcAlQgITR4zve4YUDbu6e/mmEk8R
LxEio6IXenPeLj4ngXSPTryTp66bmiEAAyrZ7QDOm8wHspL6h31ZKLOLyvdAVTgr
EWKpWNUOJLn7FoxRYk7G6DWD1QognEZ9Px1R6EZxZCVhwDPfKGg3YMd0cizNNz6j
IasnQCYKIukpFl2DdaQ0J4kQOgtW2Fm3DBSLNtPox4s8owQ6+7UJupdNsxegcvpu
d/1GkTiix5vZ6fhmcDCOAoe885rC1L372DPdTk5FtghOWFJ0ds5JjtXN3xcTkTGE
9d2EhR0MWVWeRs+w3H8HxFNODq4yDkT+6l38KvTTJttK/vsG9l0pIVr+lx2+ruNm
wTHYbiMNqHM11ASepE3SCAnnaiQQdpVIsbmXCrzFu8jJ66KgJ7te1DWjlL87r/Y4
Zmn/bLZwUv6KgWX/oL3PUwsX2s4/MJdldT5VXufFnXY=
`protect END_PROTECTED
