`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wU80yk++Pm3kqQYpFJSir/Mpg+Ph5+r6VbiMkzinzqZMsYy3S8J49EP8cSzFwiB
+4Caj6ft+5q/jUhqoAJlbn/Siemt4hjD08VVrTn4OcApLhuGrh+Zr5OQ6Q2n+QjJ
lHGk8Hyn4nvSnB3auXaDFf1b+fJmZ1aPXpIELic95TztQHJaV79/n4PWcoqT6Hen
doFL0kIubtC2UM8nlow5cylp63ni7tul+WIknfifG7HE/JQbmIxkLwi1OXHmllsb
cjSndA1Vwo54hkMQ/UAX3yiqnJBcYiZJ5biQtk6axC6hRIqA8yOKGg1NtAqk6UQ+
gJOQyxVWCuWem7LK/+c+m0GeSg4HcKnUYTzJ6OFDdzM9nDbJjKn0q2ZrBff/yAzW
u3a0pnKrJC6YYso/SWxX4NVLtlX1pRw7eoncguSBGYa/C3HziQW+mTG+rrv6MUvB
b7W6YyMTMYqiBdKeR1cf7aZ0z6zvVqAIcWNV2sakFM3jTZA+i4N45FYmaeuNPpMb
hc7FpGzojwPIpyk+Gd8y5HOH/JBw1USdf3OBHp/rIXguZYmEYb8j5tPDsbt4G8+z
sHITrKFf+aWu2cMClHM2nmSWiC7Oy/J+z+7oLWKYvBHzP56a8UCqDkPhy2+gKSah
i2Hm5FZDZV7kWYlZXu/hPkIV0mS1VMXjoeFopPuRD2tNb2/WVGQTKsQeDtXyVQ4O
lYvS5oWDO+qh2pRCMTbKVrAXp7ZajWfig9dJcJm4zZZ3s7x+kuVg3H0//3XfxvHm
rGjEO2B3gnXgRs/7npsdPG6PrjJ4XgOleuNFRqOmgO+UMqTZbD/2PTBCYFy7NARm
Be1YX3qBE32xnS7LTDsrDqrRAAj/9TbDzWglvYp5j1omU0admlVX6eBAUv6Pcy/0
pKq71WcmLSeQ6odF1SzP2oa2Zhovu4Eee94dmEYSJ7Q6MOIjBYRIRs6RJYCYDSo6
amYfAMWo81JxMlZLJJk/2V5JpNFkuPHOWGtywIJ31RBdUNYwupIfOd76sDTRTYEC
r2TCVz3drAu+OdrDZhcY6mDsLoQP+5SjcbTOFsjGA2/2k0n8Yt6uPjB2950L+Ugj
7siEDI9p+tsLbFDHFUBZ2MsVgtIkZD4SQ6C2sjWoDIGhVi46qv3KjPElm9bkfI33
bsW6PlCvodgCJS/6Btl0zCI8Gq17Qd0BGb+6jAd3FqhZWBQURf5EWNlF8EIjCcck
1aH2xCFwrx6H3mDmJxJX8LlwjQ5Xkn9HTBkGq4BxsOymP4T1b/VbSAID9FLK8Ao9
qICo0LeFnHJSCRaCOnxArQ==
`protect END_PROTECTED
