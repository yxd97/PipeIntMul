`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u4JRltIpW8sLe5LKz93fcmocrVib8Kfv02PDHt8hGDwcvE7Q47RNtdOeeBOjj0Zn
/jEyOw7sTd4vDh/6rp0zjgkxl+AtsMfqAHM+SA4pjIVWy55sMhfL0WafVTyXP+UX
kmkGQQMcgSHSH8v7bQytLd07s7aae7sOmabL5lbJVT7p2n5H+jew/+N2R8naf2ey
5e1Qmeld0Urk0pqV6zmqIlGUZPAV6YTc6jPDjaxAVRChbYl7rgshd2a6fo4PTPff
ajx/feBjPLeLMTc5DyHEG5UZ+q4bVPSXTDWVUIFGo5mKEsOtBhNv3Ac4tTajFDx1
YrSNJx3v7GjcLnNEBsW0sGjlRc8twqYevAtfMqDMkc0ykZvVgfIiQsKN3TxtFSs1
+kXnj1tuxNlRCDqKC3JlICggVAawYziAjfssGeAf2SuLr3pdDLVT6pO2q7EdPtpD
JzQ4Ri/2kJ7gi9Ng02rLZK4m7zWRI8ZkKzyWOQO+oRBm25htwp0XOjuDvmmMPlMi
L8qFxZpL+zz4pxSNKBYN6Z2u9iT+F0wedp4F+MN932tTsZx/CU65R3UUjdNAPffo
GfR1L4wsoULnQqT1O7hwcMLbbXe4LWNy5k9tda7YlweWF/BBivQPELqst8O7p4fH
IuMlqIDwjTJO4EY5azAiVcFyaTrBsp6o1gRqJEt4oWB1grpCejjo5aqL2ZsFQ7BV
MV+sIzRojQ405uv0lezmFsylRIf5ewWTF9TicTqiGUkjG+aZkZ4o6cG3K5MeqW0M
iymvCJP5fjHyjUm+hJPNIEW4iCXQlfKX0Yai4Yr/4Ymhq15Q5jE/hfkjN78bMqcZ
LT2sNhBDPbJjuxnrQ4quKRuZM1dm6h3AGQyizu5bp6fhsuiq9mVN5tgmBZj4Z9Z4
IsoWwAxDlAFD7sMGZVPgASHxdto9RxjjCrSuLdpXNnsJRk69n4ka5iaW+xp+LXz8
yo5TokBvUYTwsv00FbxhlOYaLlWgWUSKnJArKvGuvIAkElcz+YafKXn79Luw0EGv
/J2Qb6mv3dinQ1wtlPagaG+KPcxLKVvQfMO59m40F/yPctm6Z97cIG8Eum7uG4HY
j0u111QHnawQbDFsEmN7+KMi5dmbHtf3U2HFt1ijkYlfhyakRlAnfVdLi/88vrkw
TN9bXtVd4RnHQd7GX5X4Xa3R+ASwDYS56UwGl79Kp2GUKaGlR9yPwT+vRIktdXHs
W7vMu2PvjM5Lt8P4x/OI52axLk51NSFRexDmyt+LhcIkMBXzVtIe5GxnS2iRFRzQ
2e4M83ugP8RLQhf6EVfxHNuzfmPll8tbmvFRON6pptO3Vutb5dx6kIN7kVlYu0A/
mO76jHAenMBXYAw6GGOLa6RHa9wlMnJYNuZXAxgLxLqsQNtvTc1ChlEvKxuP+DLs
HPPIsH2yj/QPcACNf9tn+O6+raMSNTSkvd3sSYZN4tr8N8OBVmrFZbnpvuu/1XyM
ejHmnv75PFOUXjimu9bseoppYkeFvHjrwx2uXDSbNW/XdU6k2oF6rOvb28n7j1lS
y2ATbsLJY4rgxoZVOkoQe11rUIj7z9dRxcpsHjJ4usIYUA0yZkQh7swupYvcp+p7
asHpaHIAEynmgzbrtwaMc1dNh82XuUwBk1f+Qed+hM5YSzqZ+Lq/s1t67UpX6x61
0bMplPD9C57ZLCE/7GzZMg/Z9ikXPBkmMdJppXrCeQetf1T22cZnl47VhkJnkUcD
HcyTIceRV4+tQCFjXvkmDr+WxWEhoJ/Vbflt2M+KpsRhTSEpEhjtNMVHmWNESiQc
CPvNAetyif38hr8mOAT1kQXV1RP3UB2v5ZA0ui+zvmtttnbtOFGKcBnpwbbk/j9Z
dIyKil6Kvm0/GTZYXj4qJEUhJWLVH0KrgYx/XAzVdNLL1bC63XlmuWFPtbr98d8j
OJ6mpytcj1/txokeRb+W+mJ785bJ3oGhV9pXUZrIti/pW94IlcVwi5//ecVA44ro
Zh1dz+6/G7GP7zzVlxaccSzGd5oNyXbL4iiLNgeBAmcTPfQTjeCb7QjT7HuOxnEi
p56/0wCkCyCJPgdBRGsF2O57sL0Fa8G6no1tWCwMbgdXow2j0Rg5erQYPithaJqs
AB5tCp0KhkXiV4YJcPS0bVZSfq9HFLsaakCFb8+UQ8ukaeSABELFl8J6+kUO6M6m
Xk/Xx3cphDo5O3OzQLtu/kIAlWliXGAt75NqfYWg3fpJzUNtrgKVojBBACuAREp8
w+qCrVtMnHALBvhc18p6sRjnQFyASNvwS9owSb/BPXhYMOR57ndOvah24VdhDujd
Mj07gep3HuLlYKn2NdJCXY5RPT0w0f/LnVcaOUTHx3KnOXlq4OyH5yAWFonQGrUN
BWNC7yTVs3yWqQqCm6JfPP4CpwtbOrYwwN2g2pr82YB8HQObt6XEG/nbJSAHmE/M
AZDKTMKh5DAR8wNlrf9NxOksajz635G4P96nc/nCrOV22amTIwQCO668XQ2gd/XM
gfVYLhhiaj7iqW4X3NGefAIJP/07n5on+Ocw09rUUtQ18oFFNhnXtUqtMU8NmExR
U3QUVxB43Ts/PR/CLNR3cqqT5WMI7KQvcGBrdV2PigFRdaJALhbq7/hseIx7lxiC
3RQoxQjQ99J7F6uFuabcQA4HaRYO4xJnst/t9bFZa3AOO8RUw18IUCDVu1IXh3wL
YMk30iPS4paLQAD2Aq2P+W1gSV37rPZCoVs5NiJamNr8TxrOBBppVrRHqANX+hDg
OuSmjxTg2aJzso3yMo0kFiSQ4OUnBdYVPv2eXll7ff5EbdL9eIya2sk5bIbLYTMf
WTsBTX002F/A6iCYZgq7dQ/oHqKwQZ6vX8MuJn+T8/7J+lQiY62CiedwhH2I77L7
vOP1s0kukJCdlCTJFnpHfC3ZnE3oF6J4XScQLLL3c3+EYz6AhCgbJm7YFFAcq0Ji
Hlg96La8BicYy+U9Nl9ijyyly+VS5ru58JiVY0RCU5nIkoMELu/YxULkcOh7I+5G
9GM391Voyz2TKq7UANE/UT0OumoB1xL3EZqWikbkM+vtZqpZ6R1OaIzf7+SSRvmV
plrLYjvXrMUy1u2Pe9GZI4StpwZOK28v/01LnZZHVIiNPLQduyRpz2M4+paFi7MO
b73Wrb1kL0mgzv74HdG73C0FWoxGY2YmjD1wIG9pB+m8cOGVBHorG18O7/3BddR1
XY8WoJgSkHekm8leSV+8G4O5PCA3bdjXFDkYgaD5AxUhd5ifveeM3zbTx8uhy7Np
72e+pvGJpeF2jFafKvC+C9esMQUCiVWo4ZOdj/GM3zWQ9nKvUm9Y+mZqUOQhGaT7
0h6fxslcbAZZV716Jytb5dqT47gGMoMw2ysANtaU6bqsRQ7Q2lv5UIBMDbXb7MGa
lIkc62nrZxksJPCeViT1s1CNuahV0OH16hA5l/zrMs0eqDmoiM9TxVzLqR0NleFE
e7QVvQcynPhIvKX+4SqzWeVKBOvWst97iVgW4l3BjmPxoA7z3LZk0g4zof79L9gT
tWI49DUioJOdCbcDkKjQ/XtBxLghAxQ6mTR4VoeCKC3kNPZgWk/JlZnZdJf7CzS9
uYR39f+2IJZaKIBBO6kF4SMIiTjCqjsLqm7o3RJ64MM/v06tNtMxzc8lp6FqCwsM
cgO/sZcTuXyZpJtMJ4tMHvPVRlZKXtcQ8VyKW+xFNgmrwetOEVDt1uQ9p6T/NiLJ
0xd15vTaMdDRxsHRqR1Pg49ogpNAkcGOodzyYjUEOHiMr9ijUPnPilJC6Hu8hTck
g5jZPu1jBgzDfbZKGB7dMtt8PJVzEsFZwiaZ6B7IQGS1AtWzhn31p3gUI8IP0Hbu
vrJ5IFGmH7ZVD9tCG0WqlW9KXkB6PGkuvlyKzUMiSVYJQEIJORbDHOQTBDrOscNd
+Eb1YiJ7Ge3xd/lvHeVP64w6SnJul7RIa3cXVwPL+zuNjqCBfrWSmtuU1EUGDu/W
aoZ89t7wfs2LMLZVbtwYdO9bQVGv/ktKxsv7FKrSXJEaNYZX5EjE8BpNrC7lc3Q+
Vut8LQ/UihjrV517ovpIuwb3FnSCOD8SpSntUDilbm4kdR9rRiN0vfml9f2aDh1W
yiuUe5n3RRDwbpVsJfnqToMBSP5KmBk5nF69ZKJiisaqpORvgRMIL+G6ZvwUrqqu
tsOk6O400aloCXEEmz8ZKvTpBC4uX9KdqnnYZBUn7V+3zbq+dZL2P48yEGAvKLkP
96QIgiHVwamvaq37ospDOML9vzFRwujtiy0Ps+o+7sWAJp8Mh+RZlMrJ9+iFl3gd
4/VYpqh/Dmuqc2S0PpSMYQqX9UFvoXK2Q4iuMIEPKsMTyFvJOjvyGedbdKgCJfae
ll4Wt3XvglgHJQSwtn8FjfLt2P7mzVJECSd3fGSpCXYDiDuC8E4rgvA9IRNHIykC
i05OSu9UPf/RGsH1BkpiP754dmiO4e9YaOW/WSlR/RWqs5jM9VmgstmOv3PeGqrV
whakbQqyf9pekoc5EQtyRSULw48BRfysdHWDQ96mj5DRH1LT9u6ug5rjTwrh4aF7
QmsFdzUO2mqU4CJp1O1CVi8id1R/Jde5k7bL1d9MYzjsuncOSw32spM9mu5cNqR6
WgHboBfhfPkTl3g+b02gqoTeGP8WtWK2+bSX+B8Uiu692LMV3YD9hgRtyo7hJscC
qye/D7SbtG1T5hLNJlrevw==
`protect END_PROTECTED
