`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ryi7twKtm5u9BsyQWALRjwSK/RTHaNG/Drmq7/62zrCPSf3q8ybnnQR9sriNa3S0
jaFMctbR4EbnS/5nbrDm0LK1G1eefxGT5CfjzfmHDrBgCPdpvq1gZeHg45NDXR9C
mQbYyrYlf1QsA7qu0pMbXFMUpc1GS09q3kXqaaXOK/obB0G9npSsn/caBtvWDR0t
L7YN81LR3GYaWK3WqjfVFchmz+kUEBp6pjpIvNse7DjkPjN0HGUxw38T/VS8PHHR
3TSrfBaxcwYMP8AIQ3mMb3fMVsShd/VE1C0qV8gCojpwr7/NBxMI5JrRyC5wAS0o
k9fhVoCAv9akabSY/sVO3h+gjrg2RbUjGSQVaYtSAeIy9p1pghnZePBhW1ZKr7BP
wHg8UgZaGt8it49JaNq6LOGGACvXjTRJ+pdRXSDLvQpZz1844TiswqULKt7tk5cf
G/f94tQDb0T4Fag44gA6Aho+GaqM6V6SI/V18Vf5tZA=
`protect END_PROTECTED
