`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gv40kCsqTfsar6T7JurbX6U0HVPsomXf0ut7iNDCoqHtQjl6FnsWPO1Y2GHRQ8/Q
ctJ4jKR7j6lKpC7bKU6kmKOeTyrKHUgcSYNJ6i05qX23bmBfXM9rpeT/Ol/Cq2BG
0JRxTIexRSCejY5kYQKdreCfaEYb5kRq3Cj8QHgVbBvT0Cnt51mokZBQsAK+doM8
Az2DJrqBUrincV9TnNVmoStuv+r8e+9JbNMOY/WFkem012z2w38tYoAkdTlh5p81
I3Nnwf1vlDopiDzKPvxAzXnWh9fc1m8N4FdIW3xVxQOBfzOqonmn7lzosK4g6Q86
scN72ZXUOpIZlEDX2UVBEG6Lydmk6aoqGALBrJNzKqVNutuem0Piak0LZHnsfNIc
4VGisae6z0ytJqMqnryATknn+R+pkRnKwDpQgRhFgAt1wkY8YjA4jhv0MSERfZ+Y
2RZCkXR3RztHFKTgouH731W9oM9Wp1covJxlzc4iCIE=
`protect END_PROTECTED
