`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FfxOne7ENUWcvHtMM6ucXHfNrBA+VPzMHBB5I1kAHbWbJruEaXmq56bwuhaO8eI0
v7XfNRH+enavExharCvdY0hth5jk9d8OHMALlKQ65vyLyyDZcvWmXZvprHIjP87e
dX7Xc0rn0CvrpAhVVE83l2In/cMSv6tQGyONR//4p1EcswPlcIbt5EE/XHQ3+owq
+UCpwTWyl4epoDAMiYD5dttPmJVOuXegv5R0a9DWoEkSk/lqYxczy7ezgtrIl01C
MUZGkguGbWDRUs+ZLivjFR5eWpRJFfuZgGaW1h7Bm7BEonX2MksqMfK8C7urvo93
qZqB/2tP0KSa4lHuyJc2aD62FKP0HX9vP8+IFnnUYdxGn+dxYEhOr0/Zt1djjkxL
pzJfe8hrMRmO9i/pTfairQLOqGZ6xtShhz/eDzAr6kg9idMH8bFE1GMLZB2L8cMA
7APLflppG9aNMVSWwoBxCCKqjkcymfg+sNFsCbVD8oPs982OBNZhV7g5cj39VqO6
TLe+MC7ldshWtGiAB/I53SW1o9UYTn143xVWS292uHe19YzAWOINa4LLOPr288WL
WLNKDhrZ6+yCha8h0Mf8UgDQW+4X2UoipZzWb8u3HPzL9aZ9xWcrpDWIvaH/y51f
EnzvARX+xCY8mT9N/vFx+dwV0Mp9znmw+B8qEFt8Dt+UHnUW9LRSnlKKpDIKnhoc
y+/QZyinaQtJXUY2LirVTowXqaNMRvGQR7wEkJ7/d0wc9C02BfhRUqnBfdkfXiiO
ZAZCerO+tFqzWcfscVwIWmMxEPiL3mM1sNc9crXlyEXxaDW0PgJEDuRX7cd7gput
ZY+U9Xw8V2yXr3ea6lXSB0mOSiuG/WwMlwippZjtQw/AbEy4L1upZxkg5m4QNdYD
YwklPcZvy8ntE+b0Y5j0dsNQhtRpRaQ9EOs8yOItMcM=
`protect END_PROTECTED
