`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7K3hD+3jWy+x1D5O+8kJdBZnJ+OCIBjursdK3Mnhvpfz4JZ4OLZMfl5JUb/OCrUy
eYEjQFolpplUwjbRnLpZsYHqaRZ84DWuMcf9hYYpOgPH1TG+Qb/PyCmMCgWprgTo
XUnErhqnOLZrvYrb3xzlFx2QLwJm3lmgtFj36BhDMiDMXy5aMbtGvZohTeDOm3Sp
N5iul5gWHHh7u4X0ZD5qEXkZ3PEzsf60F+UGGcdpUIfBfaHGOZbstbL1ozbL6V0i
G/kpNXmqbSeAUrXPVUPUdgQkoyRS4vQWX44xb3Kh11qfOI+LkKYEHAJ2nsd30Ajr
neiyX3z26wzn6w4Z2R3r83urIY/SwNA3K5oLl4PwwgPYxB3xNjQk1WmI7eHVEjPc
NCQC0rD5Nmwru7Q4vJsFhYE6LhN1C75jB5sfoGLi2/wgnwHcMDuy2d/AI5vgbTRf
hCkqTYvAMqQ87qWZVc5JJ0CPFI7S0+7TBXMbY5+FrkU09T4xbHral6s3tKeSidcE
gW3AiZYdcOR7ZShUt1t+wAh/VYXll6ce0vmPR3W6NtO3lGFzR5hseQCQHBGl1P6u
BXSQ3t6ybNSESqIO7Y57vgB6PQJLzREjvQhgiGjw9hDlNnsZB7vwdJ7izfQvRU+m
hlqOQECZxmX06DJJ9JtnikOGayEBGFBcBb8Z30e954gwXH0EGuQsJO0D5nSffIb1
`protect END_PROTECTED
