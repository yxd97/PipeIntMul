`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/g8NQ1t62x0MLmm8sBfxZmqqvFJbrK2KUp7KhG1WjfDui4c5FKEpHElK6B2hUTnT
J1NJNsD13lI1kOGuIEaHiW+zA/YRIXaBJF7jdg90+GcKPs/do9gCyQ0k4VPPc5Sr
eMN/zKdNwx92U1ygukyR0UD62niCpieP+5NkW/RFXEvfGoNTy3rjZAW9btqsZ0xa
pPc+Zy/U1W9xQkypHZGIt0tqDYpij39xROqCFjYK4mypbQj6BOqFCQ/jB8GFNFC5
MDwzBlmnl/RuSHAGoUAxvigq6RRMckaWb/I2x6h231xxB0w1UzwC4P5jz/pl53FT
WFnPqP3inmp+MKWpRfIJ3bcneIjba+BA4QDjTWLPgESTzgpO0+Jci2gBiqZSXrNe
dUr4JhrTesjilhGD+Tkkc0SonVlYye/bckG1SX2yz8LWXkqDLTEyCojY5UZSaAsw
s5FadtmJEmJ139kJO9WJDisfR0gdU7etGJ5coaxu9pMWvh1PysrOufqkh2/JeIs9
8EIWvi1imY0hIWFhBH8c61wOtUurIekA4Dxmknk/jyDO5zFJxTYSBWXLviso9LYN
EjXPzf4p04Pl+YPa5N8NAKDgNk5U6xyjScJVbMKplGaPbzW9Ckp7kj/NTi4VBTaH
vxOnRvABuOPFeP4I13zRXoBKIGRS4FLMcoCdw955laDNTEXMtKrmbLRo+e/DbJ/2
kuwr3x5s2RPuSD3bY7+D9eo+Qa0xyiNINcASDMlYHQ6rsLBk/AQx5h5Hv4Dn0Ww0
`protect END_PROTECTED
