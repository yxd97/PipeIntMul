`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ij7+xKCtus8W+MvZbK42T4rNL0Fc58vTv5UJ3vEzdQ05TEmqyiiK7Px1mt0Osc5c
N8lST83SNzPA4mHfH/FioAc4DOlCHEp/omC2dVzZlOueQMyxoa852iL8Dqgsa+OL
keEOLq12xcQVHzlDe5V/ELxFd/v7AHD7wGFqgj0GDP8VQsaikOIHFs+6PMxOhcsz
ZqVtT2kZNxAKwdqWEbleadQV7VDKBOS9xrNt+6WVvygLrzpl9fyxukBrGh7+tVEb
kkBAFapSfRublwE5MrfTlIzws8+tSc+NFaYm9u2wt+ZPXLmecqZflRc5NS0QEcae
GG9SHb1rXCOcfoUsJoMuJJIeHGidxTxyQFS5V9iZn0JBPVXhOb93YOccG0Jwm0+r
G5X4f392WintXs5WgY63+vZpNPbvCEqA46F8+9T47CUZk/IeD32EdfqUVfi5GilM
wmTL+qV5IpQUdXECrJgJQA==
`protect END_PROTECTED
