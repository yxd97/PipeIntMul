`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrxdvcCrV1dwW70eqmxmGNRrSShyZ0oql5K+vK6WRzOd/0PNMpG2xRWlUOegaFuv
y7VYxOxqA8zxW5Zw5n9XR4riAANsrJOQ/tcxEeIRyrWlQloNDCgDGYzEpYtxrBze
l1pLPrmqV3R+4fPX0qOE4gbfI60EeAAtlYzzp9SrK+xlkpXQsP6Y0JMiGAH/yiAr
X7OO0xxVrOxKmbWnb79CK2PWXTgJXLH5WDx7l2cpMWV5pFX6dtQ6978+VHRb/MVy
YTcV3q5WwaDNM4s8KPtwI1j/FS7cFZPV6T2YGAZIagCS0N3eZRSQTzi30q3zWxW2
vMAuodvBfeXtHdpQMSx29BSyp2ye96finpQmQguAIRWhAt4XxemPTrbf6fCcG2au
/D3JExD2/8jIorovyCrkF3T6YwHooxQUo1X27Bfx25N6m/kB/LRI2oRttBOVMh0D
JWBO8bjVYuYeryySR4/0jjdG3/rbozE5792ZhLlX3msHRBieIQMyLAN+6k39QxYC
euDz0S38I3vdVRlVQCGdp+/kbRj4CBEbGZ4MGAeM8wxU+fK5F5znSw23so4Hlnh8
BhMYqM1ePQqWbNtMoyxCNq+v/aIDLlqHfp8oVjRr5/rVUSajyp+t6r4io0ibkrzW
r4x74P4HmuV/WNAULrvLCYyCzOsJY8q8rjYUUijfPfO8ecc0hbGpsXzTAvqCzOht
TfurL1URX4pae+o+7hbmE4KjkGgiONWZrwSNpESp+ezEhLfLKukyvjEUQDDHUVIT
W1j6Q0zbTq9x8rVU7fXTRrizGgT9KeW7FgtCLBlyoKhPVQxyyMO1qYOJqNy7kpqt
wsmxwF05kQm+xKJLAhgqhM7MkcfywlYbBwEi/n9XTJA=
`protect END_PROTECTED
