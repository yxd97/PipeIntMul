`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Twi6klkoGOL64Apr8tWYLXHEVOkL34IrjydgNenTy7LIxzJ4lgc4+ZhXoqDC/7r5
l1fqaXPclW/eXxc0vfxlPoBDNsQTxyIUEVE5SymAO9cf+gJv0KD23HTVKUmRuV3j
bVGaJ9FvC/Nxfo9v3Z3WazpWrelS0CPTD6OmN6mr5G0LS8EzJ33MwfSqSZ8WQVYA
qjpcl0QFU6MRntRDfhVnfmVa0ngnQ3IDgPsEr++Sc3nTr3nCA7KsGQ7kH6sJzVMR
5FC2OE1Cg/jLnkOYtgfTb68oIdI/vwrI3SLtiwm3tfXKwe3Rz2Eseb2OmhiUqLTN
CGuTWeFSD7MfUgiF88J9oHCGqDNcSqG4ijlNtv8NbmjQkmbzgLtHglaRlzjBI47q
Sp1k4GsebeBPpulREnGViCYINNPRH5oiOLtUEMn26fA=
`protect END_PROTECTED
