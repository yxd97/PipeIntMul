`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eORM4PXhVpplMJET9EEQ3lSkRae6xHl7hxOzpUgXldmVJoqiPOdnucSA+EcSuKzJ
rnB8KIbE4a1NzIoe4po1uwu/4zx22ronB5mnte4w9Ub1NYPRK/oQZkY5XQqTz0Tq
bsTKExMAjM8wideNjwmqnFbzVOeOXm9UGJ+05oSAEaiORRnRw1FdipSWsYC91QeW
fuvXpSBOYb3LAuVx+mnkie/1ro2WFPBqCNTdWRpH42YkSUu/kHfzah8JHMH1NGRJ
+MZsLXQ3WsDLmbjG4cYVf2x8V7ewzcRB0wyZoxQJQl5EF5d4NWL8fSWtcVen7SWy
nvqB4J3HngRNjbZeFrr+KXNyN+ZlxQFFDT+iH7GmkJt03a4aMzYSRj7Q5tNy3KA/
7kL8UxnUC6ca339O+bzVuJbcxwFtSt4wm84FnCQXPBPfKimDOlRdqCQGZ7+89idk
QWs8KWFQ8SL6OKHU6PUYYTFhTU5KJqYv4rStvun/mCswVK0vyBNufpbZCdAnj3hS
x20qmC+wTr4PRBm20FUzub+Yv9Twu+FNUnPwNs1p0V1QghLRcQPSbZMY4FG2L0f+
IjbQvzby40lGm/8TbIn37Q6i6StGqdT/socC+H5MsXDaLsZZFFjHTa2lVua5pYlB
cadZuEEKAk/psOdfFOtiuvBP2u6WiIqT6ru6UwvJgHPYZ8x4B/2ANQxGwqu1dI9T
YManMWXkRSuGUm2/fi0ODbw8zMrOLHY2OghGgo9IqRfhRN51NkOxwoYEaB5c1Kan
kaBM6OepwxG7AWosohcJFUJYBZWf7tn5K7yxCgPpSpmnGibJgZco2Xey0PRkImWf
v6YKy8s6ZjOEiYN51WT94K6RE6JAc5N2aeYDgvwEscotMkeacBJMYnUzp8Nj8kWW
PS4Saoaw4ToKUdR6nkMRtTh3GOTaxS/APUbidtJowRaYHeldrwHiOH5U8beHf3Jj
hfG+JyxiLtzkqqVPwiW9a8fNqPGwLGrE5QQg5sb/VQJsauyDAlVPdyJJdXQEfutS
hBUTiuHzPwZKOupZbXOUsL7FzqUqf7C469PRk1PtYomkiXnjAyigF2b4Jp82fTKg
ttdNJk+l8QRth/xAw50PIlm/BPOTAg3MlQPbqcrSXrreO6JJBICdSDQukYI8AXBM
gM4Sqc78P2ZHreVlGjhfiTFiar0QXPF/Jc6STAJoecg71VWo35zS/LknTkVSFBIg
/7RQjprDPvCmHF6q9SVZmSoAtnND4hwKE7jeB5SSCk3YrU9P5E3UzAmNZsPyWKvj
iSY+r/j4QSp007Is+kdLGjP9Z2pCk2I6S85dHSoZX4wKSGzq4YBGw7wA42qblXKW
zHNWZOcxikzg8TmRrROkmz1VomvWidlmGrjLgoK1jsbhK1AF65hF1ENbnffflNGb
dCEoHVeMgkuXJTnxyV/qh/oh+zvgBP4j8X+NW2EDK0Nez4S+f5tK/s+AqVeOCRo7
gkxXZ1FRlp9FxzGqSZ4nY8Or5aEv3uCHJ8C/8jlAMRPwCC0ChnRGY9RfR/4W6swu
o7wqs0nnFQWKNTxnmUjrnnB7eNasVtJoBNSDBPkJKia9GPgA8YqFWmECY8Wi8bv+
5pA6aoa3o5rEtCxTdIob8M1X4yFwci3XZl13BNe2GREFsX1TE61yGdh+ZUzDTOqr
NbXsKYvBQIKK/BK/zeKF9het2v7+sB0zIehuDKTRPylt0XjKMtskJJL/zPMfrDjh
oHunGT4a1Tf+HdaA9RoyRmDkURCRJuKybyCH2hqUukcsvta5DUdb/5dpCaeSDvgQ
6rS/yM7t50tGoftjzZQBtqusI9tyZ0DE3XZxebQoNrHLgC9ne5oy0UAMlD9aVhHx
uuomoXjA1Bu7MMNYxZq98WVTC+5MzVy9jpZo7arx5qyB1BpJZAYU+gh4L1SXaBNG
w31ugjda54f623rjbqyaXzIuQ3jjJek7LAlItWTuypA6EWMifcTAo3dSCe2FRX5R
EK+jBnduM7pyMHaQEOsBT273CLFWal09pp6olo4TIlG4nSHqxtxcNwHcRwmfwUQS
Abd2V+XndlWWqECtWahdRkHl9Oy+sXIchpun1j8Pnhiwa1WSnPtLHnnnolsY/v6i
KvhsTVSOOK8Ctvwg02tmAHxaDshRm7oQ6+T0zLlD9u+Tm93LJwgPLp/GfeJ5wUxq
eNEnDA2ONwicQT6kQSCiAuR270dNCyTotyUxoz2Hlo5L34SZG16mEGd4Xf6N+Rv1
JxGedGCCW3BJAeNpWXOU0dnR9vJIuIQmkwElm5UExpWaLJme3BnJiYaHRPuHlKFZ
Q96yKf4OpFuRPmfP2HpNaGc0dDP/cbZJwt1mpm3s12wFbJ1v/DyfbpVGmwWOOyi4
H8luX8LT3E1aC0qVlAMb60dOufo7FIwAb9+zDhgpyBX6odJxx7DR9r938uDUBUyZ
mrxXq1XXMFnlt/9Rt401lmnoHIfPqMiE5xNB2/LN6yI8tOxzuBP86Wv9ExGAymiZ
Gflsjmbu0jm+g99ioOa2CCWpJiygdROkixYi20GeEK8K2dOjFa9UsaVBWaJwQMeW
1YFAN2bUroMOJ9bgYXLKcYDMIxxn1zMhqcu6QGsxe80PH86wTNigvQWe9ivaTIVD
QQsyRpgL4EikX4z0a66CRUVzSG0aUbpJUlIBY2DsWEBDUf9jDv5Ls4HNANizvtSG
7bEfcqhtShXtqRj2tHD7nfHG+qLQQM018OR569jRuQQYuOlGmFxHjcH0YjsLV/y9
64X1o7rb3jVR1hUdBR8AzXHVaK4hXF4wq4ZX4uMmop6WAddNNY28n7lNWltP3Zqw
arqUtHGyaATUGDEkV+AafHIh/424d/GsAH8tj1oS90DzbgFCkW/Eb56tA2MfcmOZ
4Pxd9wWUplm+EyeuiUyiXSbSx3OKem5cJq4xwGkqD5SxdadxYcPSpdaBXnFE5zli
5sDn57mbbtkP1Ksbs1XcVVR60wuuXS0w3nqiqfgXlDUfSJgArmFISv8+2SKxRS5z
IQhAO4imTmzMd3oA+KjNz9xL/AndJXUt66zb6hp3m3wE52dQsmsMLVwKfE/tDNHH
8zzCK/N7ZnhlntoMJFHRpIY5rxwGNQesMNNIBPDoQYrNAfUokL0Rs9lpXnMjrk69
cVALs3cqOatXQfHLCaUWbOhn0JkHFjSNts9AUCxcrXefJZJFeN0fX9wj4LCYdIZz
lW4LzHLvhl5V8vNJZfbEr9AlW13AITDmJB4c2cg17YVRwHASMeysrE2k9MwX2NpF
AMq28aL5+a1icnmqJX8mj8jxncVOkkxOHYYpAzdrD9pY/d5ojsn5CYSSp9HxH/su
5Ey4IqKcyFfDU0cJip9zs3SH7593FTrAqBF/cxJ8OMENu/aZTCjQ9mcmJWmPuurK
lzwbUokFBKNdorpePfnldoYn6IGYHZCnPp7v+guQKbvH+HCOFjXQAw17GTxceXpB
Efp5wsfzu2D8J29TqE4AKoqcSSHhqh1sKZjXSOPnxLaTWIND2n91cSI4Gd2JrBiX
sdc/UzyFLPcq247eDMmp5dPmoX75S5ZPWzS5iRHppSGtzUWsV4KbRNrBlTQmsDkv
wGWcrVFLjNNlCVr/xh/WasG4ltw0CSjTPsG1rXDmd47DGtGWX09eoCckhoA/OYzZ
cvvvLo4QJvAkq6Zfpkm1kuRm6n2mEeh3zMPU7uZtdeeqy8VvDJGV2ie5ciBUIWxl
cfywJmtIJH/mi1WUpbmPUJqxxp/bJuNNe5VrDEwMP7mlANvB/dXlttzaQ9YlbKoh
BCIy/VYdNDpocNxwBFY+jGZzzwaqekoWPmvo2eid7uu0pdZQmKO4jAoG0puiHpYa
Ejlg9WfSYeRSEgzIaZaJgoFL77Sbx9cg8iB1oaPbJ8ilZQA12m/WLYre/uz2DmjN
3ylwFF7QWYbpQjWGCKcPnfpzSIIEUsbAR+P2TubV7LsUCNNQNLnk6hY1SUubgjc/
U+4LvF+POmxXQLpQu0YROGeX/nNP63Hven1BCb/Bnv/dTIe20+simwhiTRbgjUiQ
GO5hAlipkjdppOkgvCuJwb0lusmyi5OYLSbz9yOT4Fq5/0fubNmCcD9YB4rA9K1X
kic1nrHQ6fpLWLGhuSwmkh7kICLCJ1LdvsZtWrPpMNTWAEV+3coVO7wzEMQpnfAS
tRWu89PtyOZNnccUvCuR7++3S8me+EeJgPKSC6gYj94UcGZlzFv/3oDmnpUz9yK7
ndXCdNGxM5Jd1I2ac6aAe8yL/DBdZ7hDp7HB4QdTHlexwQXEkiSkz66CDGMpCSJt
ziq8l09p7DtlrpLNBNFLLX8KFOSd23ax5sUnZnkPyEqk0bsxA/YBVJBsT5YETwks
5GtaERI/Yw5hO8Ucy+0TedyRmV6Ur3Kfx02qFdsz0344L6k1MgIlzhaauu3Dw+dB
1WibgsJLTVSTIpr0ioFESxhZhnFVsc54SbYmyazYt5zwbZeyQc50UaOW/mxmUTTj
0bJadQUPkQnd6DxVo3sWVK0c5W2b/FZzW/NHHp9eAFmEwuJYSBhORZjMcCtBCif5
ctXWULJsIP4kk1+UeWZ1HlxYoPy2IbNPx+a42FUQh8txXWV8mIuWBQiOelvLv2C6
3toY497dO5iQ3gdnnXiTSNMsHzzkpfPjdBb/OTaeXYKA/y685rSLxUAttnkD0m//
5GGFliP9QeaDWVRi55pfEy4fhkCqHZUNGfEUctB3698hvf97mvPrwTf3uBwwO3P7
yowu2UJHFFaDAF/8Or6HtKn8wiwWL8lxvyoMvFfFgNbyh5D1Jmsl+7EK/B71KJSx
PfqMWetHqZKddhxjTSrBtXnsdfVyMeCjAUKqt+zz4Yp9LvyvGgu87N6Lr8lczNOd
d79H6fYQtM4AJlqMCHUXiPAHza8Z/655obE2/7hLtPce5+9ouk0dW9rs3n7CgNRR
zZYWIDfv1EqLd+3Gb9rQ+XZkT1EVTPWrIanG85gfFqMrf/wYmBFIxH5r9l7lQSWi
ZxU5dwlSWrbDEql5X8t5a2B6wjGe9sik5sY5Sjzxn0jKxc5uuxTuSHDmOU0ejJ7s
Ku8xbdJzRy5yTMSrpo94iQrtBQRyATuj2GadkBF8W+flERiMArP+SAlAnFyPVbJx
RC6C6GMRuiPnLlX/WiFFuN/MOIlxOAdvzPBfhhVFcKHUstYStOYkntqKj4d2brma
3eSXqWXo3cus5HJ3rkevNUAAb/Dr8CCkNp4e3lHD6TDO4sV8hvfqGaz0m5QO9OiM
uPHuWQ+F6Q35eqOL23fCm5xH++zrlhYNTQpb46yrgUv9Eq+uWLvEKXcdTkKcprNJ
vP0xQi2EI6W9+AMfaaec+XPdZczwdl50b8/+ug8CeyM0Cj8vGaaohZyIul7BaSSJ
GijxBH+VAgSsd+dFrLX2JFAI8mfmChRtNRjLDTV/ORQgJorxsSD4TB0IK/Ut7Bq9
R4UllhU+c/erOHwBlyrkpn85wRcYWmwnjywOc41B5w6/fKGbBNyl9werdrOP2Vmq
KQcHQEtzYChfc0rW+e2Efyv6/hd2oNIyPI2IMMu+uQmzkZZpQnt5TF18hB24kSpK
VetjbSGyCkcBZ8FwfbqpeB6btsPSZ3YWiTAHUSCFsio4V2uor38VzM3eIQLUoqIS
LrFcDDvBwSttyEOo2gspATMbuufzcFEDszj2nljdk5yzv+OakAEfzn7YEfnDhAcu
Vz+NKzwOeT8NM1OT16R89atm/8B8YHhMEbAFZAdSTa8IxuCIN4p6o0nIvee1btFQ
S/HC7Xls3jPmH4hTWnMYdfzu/7vEKd7SBxQqKe3N13AvCBlrUiIYa2scJDCufY14
3drK/Vckn9gi/QU5WdqY3gmp4aWM1SBygfX4X0iLp0hxhobpm4MbfxNWtPVEISau
WWnbTobA+69CO2N2B/+cNJofYmudNH1ruFky6hdNhxi3WvAs2C2DKvTyAzN9jqY5
f/fpN9clfrkOoymI57zr5oVQzqVBRu1I68kO0gK7hDikoV2cBUillWqzuEGkoh7d
kYeCvoDyKufFCrYMBF1QR9lR112OIlJugd1dL9zGJyHoI3lhhRDso5JsE7wj2+9n
tLJIihT3CZHU54/6EFzvh/eMR/jVVTie05kV3500Hrea6/bepncnR6tbtGMIRPTm
MIiF6g2Mw07nubtGoJSjgoudpisv0mEbjbSrCZRMKkpXhdfBSScmpSJkkJMKzWkk
/Ft4MbTzCh20xzFZmSZa00o7dBJulxQEadDp3jkJ9cV0M6GA+gqtxEgkcnl0g3Es
P0fimkybBJFCD77xbeLIFlDi6FpbNFhcxtd6XEZa0O+IHoRlvNBQwDReAARh3tzO
azkv4TDYxrjRVgIl3hpneIM72719APy7UNcqp5lhZBC3fUcQ1Xn5XWcKLsA0VUmR
xFocP8stVOFiU9xekNKhU9/z5OPhkL30m0ckRswrjQIrUtAHeqqZ5G1lJ6w2jgvN
nImYx5hxTRJIrMKQFwQe2R6fPp05cZ5eG1tx6vkwoxDMYXXNljquw2zXjtOiJbzu
gCABJqlSI2HxJtBK+HPY6H8UrpeSYMBAcct1xIFk6nrXZ37SRDrUMcbedAa/DmmH
73PiGYlhcWbJwkudzqBY0SoKgqtyJ5BC4OdoxZ/9zehorf9WISyw04Hnr5VvEtdP
PDoOtHyn+a6hOckSjdUTbECGg+1jrcNRLEtSmvU0kzEUtCztQxummpSLJqnJrkOw
fwqG1vwFMtZrrWz3+YZs8qao6RagcDaI0kq/k+9dMuEQgJFLSUt4yCpcanQ86DF6
hbp7l89kRyfohXMGuBB+DLB2gOOaJiIyZU6T9ne41+wCzZKDsNyLIGo4yfW92ovM
F5984xHks8uojL22edrly3UoNDcQ/5n1No4h/pjx5PqZORyj1NP7R/w2s7szUUg4
3BjfeRfkH91JgeURoGMnNaJ0zXnTyfbyjtmiYwxB2SpH3q1VoSQPiVZOS7h3k8vi
Des3mnlnSOCA7fV/n8uKWdHPNjz6RSE5Q/iOD+HW+OR9NH0Wgy4oWHG2/H1NZJ3W
DsapbESupwEbe/TfKo0W6whbfoVV4Jk71YM8pAzn6wboupzLhSvIg6euLLQRPI9s
fdA5AT/11iKbM1VbAFwc1rINOljt25hNa+wzJufTUGNMX8bx+5B3tH6Svd+GMIBz
ezYum2NAQBiG44Q4JIbFxJhav8dtLrVPv5rqFYW1+TALA3KirwRHFR4aVy8bVmLw
P/v3O6FU7HsrtTxSFjzS/0uOEFeQt+IpTl/tdYpyC4R3AgH5iuc4vtndRT5xWx5g
5y2o5uMFuIcYEcDTlwcTNTUV3VLhVFZynHf4Nrt9sTeEzrA/59tkUE59u8uVneeU
d6Q1UEcowuUOg7LLkO3HnKqdsDSbqC1WX9eE8GEhm5PgFORzReXS7pwi0ewKpxVe
XGwgSSu5nmk9BiUz84qKgxjYaUjq+oQNQiu4Pk3B+y6FpBvHpO387kdSH62dXVFy
GcYt16CePFP2paaFu6LKK+bUgxxWpzBZxrW1ICzypC5XtcYzVzwGenjS/wbLnmkx
t3/8bPlW1TS9K5qT1TeQ0sQd5rBjDw7YAj6FrBvGRNpX2A3fiyhh4rxLBC0hUMfy
qrNUnw1/bwDc5u7G8mtWKK0mF9SfW94X+ZYFGA6ovZxs40WuimAaIjwKW/cLuNKa
qH0QNrnfURf/lMJ0CJdYrvGDniMv25yxG2DwgDOroy+RNmkRqe0rRGvD+q8BJFb7
dcxUrSuzdcDSF6oidYlNGHhWJMYSJkyww3rXIiy+s6eCo32oKe9DuekD8xTafZwL
Tv/8Xy1xIBpNicHRN/ySkakgUH/Dp4URzAQ3UTtUSDNcLckCVG/8JhdWj8pJE0cl
4c4F08vqNseYtL39nu5Llz28lAqnWdgRKb8Zm1VUAcDtq7b1JUoza7wU4wNL0agH
ki4yw8NItBWp6LRwdiV5C49CKGgbIlIsTQ2O9vx76DmTgOcVudQaV5Nl2wrFB5NB
4owEPA8jpYG2PUTfz6f291mXPgIg2LfSVMNtI5o3XW73xahIwOM6rf//mEtU3nsi
s2hT+OUyZX9YLhUtLabn2+2LhH7gHOmVcJB9Z0wcKFjovYVcFlBwmIg2mwzjBVEh
ywzEEJthSqal6wTBdX5dUjXH88rLfOfueEXDtQ0ZjMgVcMw/qFyOat/CXhKrQ/L1
1cly/SyGguFPP1Tt9AcmW9Cs+wWGCSrJFeGYqdQJgUfZ0PMQzT8b+H4j8IH0HdTk
VtpJKLwCfzdD4W6uhiljY+NPLxYopmSYuvx+z9D9cBMmvWtujXvBWqsKNhv/3LgU
Oj66nzoz60OrhoXbPpl0A5GfYxh9z/4F59bqsTpvd1x1S5f8b43l80igUbXZkMeN
lf5JKZRYFcSnkxmaIj2xjPYJEwcdpAZhi+HBXHLMsASFRGZccMs4noHDRIZWIl72
0dY/mi7Ram+6DMKTucimciENxkbo/JfTX8FGI8Epse7Jm5OqDMlVB7tgLeeoJbbn
JICehSto7fOHIJNJ023slLUJyAFmD903AMHakExEj8mBG47DMrRSdToxzbYdIIf8
X4nCu5WPJLElg+V9elPWKTUbwWY/Ysfx44h37b3EL/M6fyw1ENCcwgZun/lJalGo
Ts1c9g13bnAzvLMSuc6uduNIqAxIueO9MVJmrwN1SrdRdo+omVxAah1SZ25Wv8kL
uYRYg6hO4ZZ/6lTFa1HIjebQb9hpb9Q/NayJc4oOSyGAsWnK5bX7sYPRfb8XmDoW
VlRmD4viMXh9rIeP8um4CrLgh1cv0t8LkY5qkuAhZpyKTESACbizXhRWWDaaaL6G
aiWzthyrAGkYTFejLW9huJgxeb0pAW/v87l+sW0p6hcaHZCPHJ9Kqggrczk147ih
5HVkmLBRBVzZMoT4mz9AQ+6BmTOv53VB8ygty+a09ORbCHY3sogCd5ll/M4esE8/
z99ap4HoOfPnorJzRegmiNVAwaerjv3DxAIS+6ESib50l00rk5sWRbXjrNTvfKyR
uZfY9icMe1/UnORz4DCccV3GAw6M5yPXa0B8i81EY15VM9a12W6Cn5kfexXF+VLF
AR/Uk4j9usPPk4wzAh1qQVQ6jWNy9xEIunRPi7JJ5yUZYqK6zdt82CRe9ib75knV
Yd25pyCUQjna1f2LgLxZgyvXsyraPYAk51lJzRqIS71dX4WAUPSNy4gf6EMB39Dc
UokxglgxVCv7JKdapWrw2s58xlk0kxu/S5DC/pWWqeO0PIoIf742AwvJxUgfYo/O
P7X9CIzmji4SvFr9w26OTyWn3O4zfdPy/qwSuirZuQDEoz7/qvZFojAKq7qvV7gt
US6BkGz6ddZZ1ne4YquZawfGY4dIBnOYFwAKeG9VQDmkueM9/eMOW42iX8Gs3XwL
U0+rEMScCXVOBvk+QjJh36RvtP8z+OXBIEUOgo/Eb0wR/XrJ472dvONJPCIN6C8x
e8s1XsNhttqwq8uLeZkxB2ivRdrqWh0OE/L13zCMhsncR7UhqlqLHfKX7mo6V6Mg
+7QcFRqsuTSsWy039iO1SdIlcLVpIcA+EP+r6i/lAQGuUESsrkqkRxfaL3xnfFs/
XJt9nc4L3th350zbPDBV7QkVwlBAAa/GE6Yvm9PjXqP/6OiyrY2nG2p03qGI3n1y
DVMST9VO6pVw/7sjPqLzLy6T5GLMzGxFIDNXTZ7HvN6GwhGkC9+XY55BPpqBsqpI
tsaK1xwFIR+ITvgmrOvBqBJghzGGCL62csIi4aCaK4SlFBzmLuO8YpAy3pYKW95C
FfvF67MX4x6Xfndme3XMcrPtnatbHoWnNUol5CZfu6zpsvhvoi5TLo0JsnwSptyn
4OUuThvh8GU5cZ6ESql45FbbWsb6MYGaVu/EmE8NXDzB6ClTJYDy7J3dPoEWm7yv
6Nv5sVL3osN5bGQSgrhoPIJVsNiZwuA9CMBar801phEt/KT6VWVJZyvGa5icsT+2
Ous/spH5PsNASH5R6qTihmJLpAmxjgNDCpLDYaS9paE3IGAVfLj/IzOR1HqeNU+l
/8amADgWVYf+0BvlPscThpufwfGUWt/hRka6TlkYoV4XoAXILIdJxdz3OToetlGQ
0u7f9ExsLIT8JMjzCFlMEar0CKfadYoLW3fENkR8yKVxZD8IYVLNEVF+A7RYblUr
0WKOmwSsqYftFHbsfxD0hOfWIjoh8NfzKUlXkQ5BQkkW0XrgyfsAVcCzJH/Nvm41
uTJ+aXgvBsdpZn/SzQpQTuCM1nHury/w+pV91pJubyV64qP0gH9vQbyhILpLO4Af
iu8QMtkLDavBvkMjAu2NlckTbv/h16Ce02xrOZJsDeSkc6N8r616Q/diGveSCkf9
faqrAWBP97WpB92D2hdkjiNuOplR+iryh7WN4hn4FB5zCRDKdlAF+IcPDec7q64R
xJwKrzQrSAJbnFzPNqidKr/Ua4yjUAfPG3+25ieEQ2HU6r0sl/WBiipkmhjJ2qM4
T4lOTG8Lh/k8jDWVJfj1o0tMPYDc9iOWM11aAFwg/MGQ88XC39CYVW474y6rOYnt
tz84rtFg9qrHnnvZ3MtQERJj16XL0PVm9LgP92LigMyB88PRKWE21uqZhNP7mnfW
ItWSX5IvviSREKu4uNdsQBqMgDtiFjDcgvAcqJ0mTolkTgdwIvcGhG5R16SJgtEK
QzSH8mSCZevcWFcp5itjdM4QZpKUicpPO/sBcFlOUhuSrjnk2CrjLlnnl8h10Mmm
PVM3GgrNWCAAHyC6hv2qVhm5rkVyi9mnqzJs0xwiY13KNdRkyEon453GwXuJUd72
NAAJJNHNYDX9Bjd98lLtKsgji0Gx6DtUdbGCLVj7yuRP0QZSRrJyHZnb8Jv5c2uF
vRtvdi1t/T28A/5JOG0xfgvYUlCnM29cgk477R0EpGr4DrSxvsvVaaiuyWxJMrIo
1J9fVJt4Er56h44isk0NTuyoRGDRrEmnoVex8m9Sbu/+qmshcADUQR6NXijnOUgz
95XkOzLmMn/jfwI5zyuht4zb9iWtIV2Uf74o4LZArYaPIxkWPq3hl5/S4SGaeK/b
rzetcNbQtNfR6A7Sl24pMmbLbK81689gy1GJa4G8bDxPhsfJpRLU1j67ateIXvm8
M2nj7FV/YOu2DE4qn2ccff71FAzS9arzZuxwcgn+ih2MFsCJ4iugUhnRiGZ1dcex
XigB3KX05LE1n6tmv3hlS0fWgmQa01nXOJrKrB8l7B797oIQJvAh2VuXmagcj+Jh
3kCJdsIsL1NZBfCX3LuKsTe+8PNtLRRe7c8NX5lvQqsLLGDVHDaKijC99GuP9wTi
wumeTZIGJtzzzrMRcwphct3Z/i9gH7jvYgi5t0peoj/Qu2BzksBObih0XqxlMn13
GK1teTU/jH+B0aRQj6yVFYbY135OHRbfwN5z6WwUoYdrZWwUfNwYrWZkkWEawBo9
qZOKMxeT+TdGxraJGcMaiPPm7HurhnpSgL/XabEbodNupHYGmP5p6TqlmLHKxeQM
l6i4gaLzV/Ho770DKd1grDJkfVSVQBoBMWMhr2+MPQ8VhYjO+jBry3ZkR/eG7BMF
OPuJh3diIRiycg9BuHHHvNnWSqDJGolx4SL/B1qOw2kq8WcPHFevbv8dI181dAjg
DnVVgAucv1jnD0IWrYflr01faytzZBQlopURNOwuMNZy1T+EMqIUyd1jgF78mqRr
JHqP8IURxASrXKKqq0XM4qH2X//YGZqGV/IYgnU3mn/O3W/dEs2DSRFl/4iyYfJy
a3dbGNIJuLi31JDZwT7N2Xz98RnP5SNIN/L6jqTx8+pzDX8Q/mHD4wu2ooKPbrue
D0FxxesaRfb+rtjWms4i5CUEl1zz2Nl2ThAHokI34mqFoTwx7Sr4yFORlm7s1GBx
N8PF4D4S+xcx0RviuRnxVOZY6Aewou8t+QRl45EJTOo0pbDnrJmeLknNdgciBsD5
PRHeRbKUIQAUkWXIf+3rR9g9HhlEZssSMi5E0uitWSwB1WsvRPEhtr+GCoIB8P76
FLwtfjKqA7IfriDdHKwgndwPilys+t1IpNivTRsyzrJrCsyf09r/P6T2OmEy0fkj
v8UCN7+Eiq4lKaPGAOlFJ3TFRQXJTQqyS6k02JcNQDKkzlR5wkrRVDgryg1GAqpH
nlz37XE/pjcw7HZ8gc+a3U0lyvg7HDk2sVZr8cIVL06QZ+Oz/Y4FZ3O64AowMr+7
flY6Rm0zpd1touj10iy5nkNT3lSlAWFvU63t+/GW0Sn9qaOs87XoU8lFvqergJmb
Lzckq2+k9l7eYsrAW5UgJynsGmNLoLlb9ABgwbceQGYbJecH7MN703DGnkUVengp
R1F6vQNYCSv2kuiCgnC1kogNHurPD3mL2/fbfb8Nr0FLq3Ga3wpw9aWZFP69vFbV
tJiLlOLQ/9ZueA1S/WEIKrKv/QePTFiQUI0npwAa+7OawAjeH5fmXI0m0l/EA24I
IlQXBhbS51yoz4BZjqohoVBGbS9zvP84QCQ8nMv7jR0EQKb7jMU43RiLuaf0jr8X
1jjhQOPXyCyvqIh3dOengIBCML2i/YD4bPk3pCT8Wn/AlhuxG6fdoEA9sV95Ei8n
cVL2iqikFOR4ux09xuIOn5ml3Y+s7rGXIyG/dC+AYyGdyy52bbV+vwRrCiVoHFe1
jxAY/jAvFY24wx5GvnIHwgrGB/vPcAPgQbFhFYCKb06feOihDUWj74XAtnubmBDd
IzsY0aALeCqqfNBvFRTR3JulLQ4moypr/F3yrxvX5RfBUA7AKslI3WQX3knzQo0L
wP4R16XoNrrUWSltjESmpSrRMNPcVy7jNJas8utcjVuhNEVLor/ORqT4JyT8CltU
rpwzZnqsrxOMAPF+6LzAV89Zy2DBjk7hg5wBUMbePU+/4nKTMqj7aeQQtiSrQ6ye
N5rfd0nkyQHV9AgzjW6LSTdT9hf7F8WyHm+lwP2EaArkKCZuVcyXyb1+hHrylWG3
CbeVHIVFCeDNnbFMmIaKEXuwra5aSdFKcNXlUGaCkYY58rITwYwX8QGVuaiuAe8F
VvATuIR5HZ14x2BwVoHS0QbrAm9Y2cIyQKkdccTdYnt66LZkfTEym9i3WvF3KqHf
LfpvQVXhQTM2dndISpwcOl7vBvtWhE2896VrMGzmzxooO5QKSZgrkWuLsAbyozmH
HwtllNUBAlD8EKQJJinNur5Db5tHa/uBT8n2jmaZrWEHOwWGKnJMg3R4H6XvXrj7
pejvJuBPDEMVac+BElXM/ZefWMOR7RyzZn/7NZmP9Ok+lj7dYKlL6dH5d4Eowrf4
/HVYwa5lAtMsDBoI3wLVmHoFV6NUeUBUyVkzx4iusiYnu4TVdk7dpBX+oudzE/bf
CYFUK42yKeR5esi5w+Te0sd3zkoBM+FBzWntWtCp4nsDOxOuR/c8EqwPWNfJgDI5
qE9DTlNf+EmyjmbflBg7wDuvROu4GdgTFjW7y2Hr3bMb/Lp4U9Q17uXeMcTL1WCh
GfxhTMD37MI1Nek6ezfRlHmVA6YiZ/dITr/DEaOIKkWnA0P5T7MjBjs66v3pXYls
IATX9Ngibf1Nvq0kKhA4usU8mc5qrRJUkDx0LJbv7g/wEfdtOcIeCspGLakY7+rY
Lbms/3gr7TpPEhb/5T9DwjwcGJ0C3UXXGQnWOlkX46NtcADLYRhN7YWCoIFhmMG9
X/TfvlmTgs+hIE6ooW+nI2QNb2kxcKe3weYKzpIyNJF+HNRSZ6C9eA3wrZHRtYXu
txwZEnvs0UyZNU1zDK0Jzekz2zfct5Rv/If513rtK19Ou0BbZHKLnB6kW9eFGdaP
3RqoQr97YEb7Gpkl2NGIGqWMcI/rNsujfowjcYhKtJ0AJGcXN9lfA8gD8Zf1xOTg
x1V9ifj3SAYGUhYRFjNbuCfLkLt/9eSy1+m7uZTTu0aH7qbwRCAE1yGxeG1F6Ge5
B469l09M+MjIBCH9dpn6AcoGWuzNpj7AFug42gME8GlaYf8BdimqBwbYY1bDcwUi
LGNW98X+PYa+mnyTGMyCjcuYLZWtl4zoZWjYDaHxmeM3xH65Q8KBbAZCh/LaNak4
2yxP3iqdO4HCQmxR0UxPEwri76DiYQ9Wddhgdf+l3fXWJLy+AYFfgQ9U9w3BjPJ9
ZMAFyBZnpuEfhQg8sw2wZw/lJu/SVyh8AMLlmMbXvOwszi7x/DSNf2jRBWo2gAzh
PBOMBMYlOWD3hp5r6coAQoST/Z8T7hhozSjfjMUjnzz7aRt4W1PTW07ZNKixsTmh
NdibCYGm/J/x4kREZZD6myBO21/2vCO8aRpFE2RHynrBYCWzxLkrlJCNiRnMuRLh
ib35t3nDJWlYSkJFNyn86Ew0tVj3+U6K9+EfHgFWbWknT/sxi7FYryNS+Cj3BO0f
Nm9kKXzJckfGFLjJtlRiB7h9Y45XXkVFysBZ+fGpjKaOgc9B+GWUW1MU60YivN5B
YxazfujqwuZLrwpIk26W99EhcIdVB3COE2mvAHYpcZlsOF8CoZyyLlJGJHceexyW
pKC09gTEwfjAl9YVpeyF4T0UvFpfY4lJS4VNn4pzksat+5+2FvPhZzusYBYlbzeY
iu3R5dqYch6PAi4zKMSk/VsnEfH9l1aewDJuHhrczSzeWzf8mfDegdWB4F/foGL0
4U9sv7wjlPMn7d/TvGQPRYelGmWDPYJ/QoSt5h3OBDlIIl+cxB0IlACadDYbHNoh
O6dact52iHfLDoT6oe6W8tFXGjiV+0svVnTYJ3Fg8BkNlS4GpX0i+pzvrS8AhtRr
wfHHjHvooGOE55AKOraMhF7Vkjr/rFRZ3muJxEFPnHXN6w7pw9/bkldhq4jtg8UM
R121Sqm2JFnpY3mrdQ2Obb9dyVZxVLvS4eOQzfeoZy6XjeYo163yJPg+HTIqQMiv
zGGpXMrtaTzkNodtUZjK51bSCf6bJ7gAqnIqzpyPTlHQCCC6W9/k4yWxKWLO906C
39ncsYDTboaiACyo5Vi2fLUKiGbeNbujxv0sBvmNo8DocddMU9wHFcgJ9wtdBvIW
4aukg/sWPQ/WQA2S+imJ5IyZPyDYDU20fTgMPzdr7HHQ9lhPPebyMwgM3Is5/Z6I
CJ/S8t4z4g5D8kfzvAwity3cNYvUYrUeXwAbC7emGZBNOAL9LYVsQyINlMPinaWk
i0FfFybhjG05aT9BUeruAWtl46ZaKqhhmKRW9KC5qtNbwlxUDGkC+EzTKuzxh+CM
+ge9eQZFISpdqF36E94T1Jdz4IBYsJmeTk+F2X/RfsbB4+NkQD94ss0m+Fh5Luu+
wljIegcClTXw4ICkMhcnvAKH7r5pVOKAlkHklEBrsNIxQn6gNFQfqKui2arbaVt9
k+WpB1LNPIaK2lMTFur5siybcQhnjcgVWlt5EN/ZFolSPQmyKyIQIQUiUGCxhfUm
3fs3neRMhvADut3pAGx6Q4xszgQI7A4trBMSI4u4A8p7kf40UXaEgoZftJZqYn6F
ujrV2YdpAWtsPhHlGHdE26PrRHTH3BoVjDv1xQyPDTq9/72DSZ6Ec3PHEBhdci4n
VqJy9IALJoP41ZSlnWdFZ6laXgeO+y/uHwKTxnwWpEXEBEU3bKabQKR4cVJsZgYc
Epaz5M7OXugBVGYIj2NwPxc004NQtxsc1QHiw9kgfcgw6l+LMYmlHoG6ZoDzoM/F
FOJ5CK93TyASlU7MFPshRhz7xErIYOYXIQxINAcuDSALa2fSUYwJoH3ZHMz5KGf0
PrpcnK8S8hCdbhQO24GzNCxRSp1iYHF2JGYflRo/Fn/5L1P0zUQfkBZJlez0e0Of
En4LAwrzHzjIFt/JmoR2P/cfT+EVWlnpzs0WvPPlq8zu7IXAxSoQ8gU7R7nMtWSt
x/GjMonMY7dovnad+rZRZv0fpjGVRkf5I3/DmLtfr7wbU83y1cgGDi0qDPmo+aQe
pNFXhYwEe8Jc78T9L0lnawbrKs8i9p0b2mbLyLKX3dUcZ8MH9v7/pKf5f5u7BKOt
Go3hLMfM8PRjSUAnTdeI+85TK37jGJAuAaMaE/D1nz5UD4LkLpWPLAPB07Ir5tFJ
ibNqmJAbVNmVZkuhlZz/bfshMdIc985onEwc2e5v+Szri3zl2D1L3VOpu645N06o
wwN0ORcprUsrq635C/IKCqogHvrlJowerbQE1qzTW/5zIYb7JzzpuvbgmVd8NQWM
LmbfmkprP3zX/Cddvt8T9jece7RcAtoClOJDngwLbcAbGXNLnRqBBj3cJNKHbvoZ
G5uNH/IXTAS9mOhPpxOpaWSkbuZhF7/mK2/sU7HYze64kHPkk/1tqM+2i0yuCcQG
XYjTAv0rwSphSHhoSQcxAYHWYCGYh4yVl6ONgufZsMhIJ9Ksp9WM9gUS7Oabmzng
gXPJgc9fs5AsRM33oySZLSEe04w0OXHP+LVLhwbkgJipJxGJy0cZBTwiDtdr3WiJ
fhRJ2KBbEXm4raowV5JWza+aluQtPhDsN1yiCc09LxJqb1OOTp7fO9arYqxF8awf
GNuGQ62qvE+tJ/CTYAYAPDj1PeLITx209/pV0p+c4RuyT/qpjHDKBc/FS0wXo1k9
DAHNJYoaK7rjVT+GKj6sY5WibvF9bCqlEVK0ZezHR/eyl/VxYxxsfCupQP6FK8KW
dDuKGcDKCGbDsMVUV/4GE+l6LXqxzyKNUIb1G9IxJMTDoOPQ0EC5S9epx8oPk7Ox
aF6Olkq+RTeDXLS46uFohWTILg0WpmdwGMhPAq8r+6h4g8sRdcgBdzOBIG6E5ajZ
zJOpnCK+BBHU2VELvjfPyWxMJ3aamLlj3Vldpi8/cfTzTrBjsT5jWur+19OMgg2r
YkgPLyFbcnO4xsCnQYXm40vmrDLqGMvAr2JJ2TN74GYeDP8qtGtPpmcXBisgdndd
lVI1/PiqYw0V69YkAglDZP5/Vnnw1hbaX+CFfMYzNrom+L+HdeobSmgMwG97QhXi
G6qC8Q9F9WGBCrAfXoSON/7vOgUHk9AFIxhKtcIM/jARTltk0cimT9TGEVJSn5ki
3yH1ggZAdkvEPeyoOijo3b+nQMxbsxpOQecmxlMxFYMFC00/jySLhjezXBJ0XU/n
eKeQOs13kROciTfuSCCRK3Wzre4n54l7lhMNseBoJCCtISI0bDEbfHapXwZixgkS
BQ2ROVF1X2WP7xDEDDtiT/05pCbrzQVrnUDJsN3dHJLJC1LQZEJwDnddCBhtwyZi
`protect END_PROTECTED
