`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HI0rhrEnjmi6YT2Sh/S50I9vLJ/q1ZPLrRsvGIajNBaHCkA16C3OK7IZDRDIWa22
MMV6F9VZ3P0kbUXx4J4NyMP+P302oFbNV9lBf1NHVbQIYOYQ4PPM41x2mAKhxg49
jEEHN70yWU6PivPFcXMTY7+LhRF+KmUlcBITKVgXqlemcXIyU+oHklvy2QXfYjqz
5tbI0guKhaZKrr+nbB6yGVqMmEh+asUYLMaS5F+TaOZJ9LS086sHZ60O3ySaDNR9
wyLhBzD2NONytCEo3OYgZolJc7Q7PJBuXklSvSpZriHj9pM4Ca/2+Q0FMRxh5W7v
S9RGwHPxMGUb2Dccj0GzYoynALTCOY8/+sBfVt6LLRIwub/S/abWsJ3uWp2GqcN1
HTCBQEz26DO+P99WPmi388em8ids2y7p7IDeOIqQdzQ2ikU3G4Hljud1fx6ybquR
+OHlJbqAPThIB6WhDT1/mUBIZ40n1H1m+ZZSK/1adURYDRSvZColK4hxFulwkBfQ
7jtf4pHFbL+AEb9W53+Z2bRcuYjF7LG0ZIeBACU933TsZ3IJfuuqZ88uJ+tZ01A1
MG+sfCwFl/228yx3NwVHqM1+4wJcCroB9n1X7RclVz4DM3bWbKDDC3ZhgsL7wf/8
jyA9XsqUL7Zp5pp8yje84Q==
`protect END_PROTECTED
