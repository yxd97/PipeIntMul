`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5vts8fkHDf7uUliVB+b/6AACjxfv/vNJQXCU656vlHaTq8a+Gq5uD+cTtbZ+1OW6
GdLsCGVMx6Rd/7d/lFL9baqt0duk2271Ond7uGizjt9M/2TdGoFqL5rI1f8R+xBh
8r7iCiezb5EeDVxdKSxwVo8y7OtCxdQVUfneN41Jp/OzBKClbHdoO8pVMHlq9DHb
SPU+xuybot/VOAByL23pTxeDE705UORHYM0V3cZ/k9M6HNtxA5h1mOz7LRmijJ9Y
ewv4HECe/x/YrG8Pkb4fUw==
`protect END_PROTECTED
