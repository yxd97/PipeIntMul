`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73a4vxqI7J/J8rCM6aFnbC2TEoltfVze42q8t7ER6yDuPpiM0sVRkYgkxqs146uT
4mht51x/VnS69mRyXlP9AcSmbbbE3aWAmXTCIcrDzrFLbeC/JUzdf+8/LY3Ma5Q6
QcBzdOI8Co0gaArzu6JHyM+yEZq6Tmg3SYZTMwmPrW5mjzc+No3iJlXIVnl4hCZe
lQKpV+EOK0o+3uE0qODR7ZEA1HWhBDBZX0pCpIw9VVzb7Ti1yBJZCr0JuOYWckwd
0Boa3QC7WecvAyw8zYA57q1cjzwammXR15r0ljkHoEN+6vTfKSVO6rLvzVtjrkUO
MTMqa6aPJs5kfwdDqSL9pKCc63h1EwwdeU0t6P3iDvqjSrSTtoS03/QvLT6ULiLD
rKSdK9aXS0yLbwzeq3nY/BrQWKk/tRobWOU06VnbzjmtUuYhTEUrq3Ix+kMeN5GM
TJoWqfrSwC5i5VDR1eUZXmhyqiXTzi7+ZGPutGRG/wVis0qqxe3nK/uXb6Tgz6pr
+a4weDf8fbCWdAzaPDtpxD3fX8GWeG4ZhQHnW9zbCNID0QZBXLMopJ6EZ7Qhf+WZ
m8qhR1DlRh1JYpLmT9SWag==
`protect END_PROTECTED
