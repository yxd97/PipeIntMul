`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6LNRzNnze0UEbUmN9zbX+DvZSZkmiDz0p+fZWQHcgvKhNGXIqmhnpUQtgMYQNeMb
MeMHg3ZDhyENwCp6GUek9TRIG8+TI43PUOqRYI7FWy+loLcirJ1vafDWO9NjwRdT
o8wdtEDQbfK3l1dazhz3MiOVA9TcOBYJX3htrqnu/M2YTmtFvwhO/nKvZTFartND
zKgrG9H8/ev6WJAPrjV796dwSEi3vKx6CXLjSxruF8/YJiQQq2W2WO2/LX8ioz/H
DG1FwkDpI+5u+Zqm4hK8iKHLGQujnOJlwWgNsiV4/mKSTiNBKsRYHhBflVjHjUuU
EES0vmXxiZkEPpvgbmyy7U6WI/uqm5e3hTmnVBnNN1ObVVQgUDedJCfGU/HIx6Ni
lT9Dkc5J9gFPD1zrBtaPqPeTW48dLwNduZo4cpjocfBqIzvbyrmhNiClXJGUwxgd
724Z48oxkGirldrWFk9iPadab56NWwV2KUbPTXU4xtk=
`protect END_PROTECTED
