`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/2P/r2DVWq7c/Vls2x5jprzPwU+uzId+mjQpUW+7AsgHgiq722HNmcIvqK/fRE7v
aScd2O8xt2Am8baQ7xYuSf0amNR5tLUGyyV1KYxBtsNFuZC8LW/JooIp7h65lPKd
8SbHp6YK2q2sp3pt7j9HfeMGotj3YUXkoyfrEqFJOxFeeqZGojXsw0JcAqMuvAke
nYAQ86PyGbC1gdx+b/pmfuCepoo513BblddsrrqNGsuo+8nmwL/64RNGLXIA9Dso
j0lpBgFDsfTGLj9WGKB55PD1NxlX068IMuAsOfqCCctmcgIuQY2XPNoQs2cUUgAv
`protect END_PROTECTED
