`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPIFiofnZ2E+T3nCU8LyyXujdjrTCIL5wEaE+CGkdc+0qkQCcFcFdqoZJqvFrfbw
JafCq+Ypbk+HNg+neQ2TCVqx8c7LyrLqB1j3r5zilLIiSVyIkJanSvPP3lPJbYgh
DQBSnyccxbvXnz6Lxl8LS3Nnaf7EuFV6XC2WRdhBJXyh+J1SJXM+IWcCd3Bb17SL
lCFAu2bCn3WjV/kBd14FT31JPIx0REVPPhITpqApU8q2HxMERpdV2eooMq+TdTfU
ahAhCtBmGYQzuyM3Jl1CgR+/BIQKL4IkTztT5fZJ+grye9B4nEREcCDAtmhKzxDo
+xvmwv2b2MHK85auCP/zeV5hHksSvBG8TfGTg8pRMCE5cdiB8bGF03v26aPZvjmR
11Ua+okrc6LOHv9tzW5EjBoI97UdRgwgQLC0E9QkMgxsO92MuT31/86Fs4iYd/FC
XFf12biy/3NSZo7cO+zyuOSM8Wuc+uWRZ5dkq1Z+TH4xI+7o0KpKgdTixKFfYlfC
L1NGhWNxr17YyRTRB2rtHRkZ9AC5zC4gqBeaXUyZf2paNfB44KxB01oUrOAF7Ocz
qv17wTgYjj+eImDPwyGZm687cpgPv3zVntwcAuis9B6PEeXiTp+dNUFSqtWFRHe2
Qg3UQAD+d4lK5YEs/z6k99fNDwHh5mw1atum/hC7ArlZgB/oLeuhLVn0oTdfShuI
tEMwYeYoiHwPVK81JZN+oHdiyY4oWqXXZ0EYnPjmDisfupbi0ZH13XKlUWVR5yrk
gac4a3EZq/S4T6NmC4TmLw==
`protect END_PROTECTED
