`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yljlia8w2eNJ3XZlTy+D0ItrPx0JDiucNkPv/6DUBe59yvUjqAtlI70VCkQWRtTi
5xYGy9QBttETf8Hqenc8RvWwG/bdhvgnDsWtBQGCthDA/HgC01XmUw5Xyfzl09/s
0vUPkcJ96kGZDdMtSeYOFhgmpwxFDLG+9f1StDoEq4afSBXevb+EwUqTjOUku2x6
qr0GvlWy40O+OMCHpt35/hdVKQXZr061m946oSdvkenym7Tr7fLB2eljRPsYLvk/
cOgWaElFocPGFRUi+rEi9iW0mcgWHbRa7hKZ61RDoSd1HhAHYLa0xmOp/wQzLJPF
HAIQRbxV62v58owTRAvKzdWPCLX/n7R9WRijAlOsibnJ7Q5aWdDXVC1BsGEUEBeP
4zFrxU9KXIpC9/17MppjrexnhvwwzbGc6pqSbuAOdE/A656HxdgNGC1JxkX27G9O
70kXWVNBB+2NZtm2N1AleBdzlT+bg/po/xEhPEgGeyJS4aMHwz0/zXiXXt8/m3cO
SNBJ6uFHDOMWVBDLPmc35Q==
`protect END_PROTECTED
