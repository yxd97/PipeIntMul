`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nfwhq2wZox5+gyVbnoHLZ1zn3qa9jEixV07MJEdVO/7Zq2/bJBWkItHk9Uj8hsvp
Sx8PsEwdNN7FlJ8J/91l8WNrkyq5lsU93G3VDCOcqyfDm5OZhbQNwFHAF0Wdt9hP
mkfJpQ8GwayUA9bBpSsbyb5Wchf+dkwbOgVqJn2v+GMygc+2l16HGFcRAX8MBvKu
df1x1Vpjwi6OWooUAK0jLx1HOiSrEg9zFbCMM6vnLhAIYQNXBeZ+5xA/1UEoaH5s
uvs/CMA6d4hkINn4xmPy9v9Crv5lI0EwLQIM+Ch096sRC/B5BvjOaT8o5W/KYQWJ
WxSN4UzB7DUMPeYTgo92em7Vaae42AlYvFeOrp677SsgHasazSdiVhP6oIHGdb7z
/3g8+6XAT4lCcSrsrFla37Fn45u4WxQ6aUcvhv76aVmdLRn3L/HdGrF6BG/wdBWH
5IcWkjgVvrg24Q1hXg60oRhaa5ckMJR8pcSGnYpahPPcGbW8maCXVnvFyguQTPJv
U0nxKObnykP2HJpC3UdNZX8t1Q4uO2413Tf5C9aOZo/CrPR3RQ23hzAx6s2fO+kw
+SF+WpnCxb1ymQ7DIbuCFIlwVwYu8dIbnEGwrYdl2l5Iz0aHOf8fO+0souecFlQc
slw1icukqzAZpE/O/miyJQ==
`protect END_PROTECTED
