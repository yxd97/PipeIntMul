`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1SjGkiFrMFASEkvQtmr5VPvjpcSqS7io+3bAigaypodfNOrjF7DhQSqRo/QaxA7S
Xo0qEvXQUypveKkBo5JaTICsNw5PrwneqWRZzpseB/8+PVS5mmA2Ph1ux7PxG0CP
utTJV2nnnLTWIt+sUOiHTfs86l4bqLLLeGoZuw5nNWQibowFHEAroO8ubskJvfek
ojNX0OHAMHZdjl+oPkveP9CcKYpcN4dYozxsPSl5JZvbfsrQU9UnTgYss96jaEa3
sAYt7CtdZjEUbOIQ9+KsxLmtKhNtdmLIlbMCkXYVirksA7MY9RCgkMP/jWa33PiS
QaNjrTJxVTrN57k8c1gPXNHjLNs5NawFKm+TiWNgmJXpRp6A2bll7+mN4o4cmM2Q
`protect END_PROTECTED
