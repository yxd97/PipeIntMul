`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/1YvZyCmzYTKjdUpKiLjwheRDG2/S0FywSApGXDXk11zsHzlArwZT3ZUYEp8Zb4F
hDF4nL1x1qHQEImlEQ9xlzKbzqeLuonnqTN+eyKLT7PKbi9UzHB6GYdbF5cvyyCD
LsL3N7bhXlF13G7/CdmFXg2rQPWfibsQR2Jru55MJ8pF5rYcjeJjVWXxK+jS5C4M
nvCHKVZM0Ish5Ci2MLPhYc7P41SwxOaLlTp/oaR8U2qZwveZ1/tks0r/aF4oTZld
o0DhI1Q6WjejMFsFU4sXJiF5bKsL/4PVXyFqDJoe3A4uII7idIKsTKE3GW313Zfr
3kYttOUApKUm558xJE3tDYztKhD+nvUroZTcaD9rAieu/TK5/urnsS6wJvZpGphD
ZavNWkXS3dSdVapcbvmyDUJs19N+t05MVkRsU4gGyetPZQ7wn7/lRWTTFEdVcpqZ
gZwpsIBZpKqIsoYF5ceCQX0+YDmjf4304a5492TD2ur6OiipzigKgH4mqp4HdmKm
OMQv0Ew8xDV3hzqctZ05GjE4hoHt5BceNUCjQp/qUN12maDpl80lXknzTRBx2jLp
1EgIzpHuAL3+8lMxM0lS94gm/vZZFRas0WP4qAjx/YQTD8dGYxL602RTpGv1Snx9
JxQYXtVIQHir/BjKUuuFOSm6pbGRmGpqmM7ZvbBfdsmHKG50Sm4WzEeuLivnzSHQ
R0hiO5ORPKSxd9oMnAfzcsckiJnUGLxZGGxd5jbTg5Vyff0jGf+gVzMLQ3nACbqE
easaGntPghynvsrWqp0jjdobhDXOvrx4iibOBEUdDIDr5UC/AKeoUprRYgI2bK6Q
wOCJZSp+fZCkJ6vYFy2cR4ezJayHtIh5Xgknj/90DB1G2I5CW11/OlLOPu0qsTIi
gdIvtZEtHqSXXWWOW+MvdsObFpHMTr+PoGOL65b5rzZWxDNWGBpS8J0CwH2VVenD
OUyaWtwJ7QQ5xbk+T5USxrVqNwh11VC7WN3zxjkQRGdEyr34ZsPFNDi6XoB/Sttp
glqCMWexk/aL/nvfXXji/KRO9vnNLkvYleNxy+M1jqwVXuWq3rXedwbNDgwf1miV
GpTaescUgG307p4ZtmuDz908Mp3cYb6+2Sa+sRWUyKP+H7/Ct0Sc34GYPzpbbrJ9
`protect END_PROTECTED
