`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2cUfCmLhXs2GnTUzKGf9l45ZF9i5MWdx0ShF7zNFx/5gGCsUV6BVZfAH8E5H7M0
DMFCWaav9RnIkfXHIQ7cbCepV49tmZ0sSULPyM2muHCoeQRqSKn+AMMMml7KmYqU
Jbk4d5kLWHD8JB8w9/zjLO5HXB8mJDiQwWaraqFnf8HGXMYSeNtcuwiwrqfJGGmq
cVBzPUUjFkeiEzK9B26z/XuQfYul3JF479LwYldoPJlNOawYbhqJa2zr+F+WLOhz
7RP5n7/jnntu12r5NX/3MOx53guFWMJRh+XVWoa/tVgyT5inPrhF0MHCHfuZBa0w
VotiMa7aRsErcFT8diq/V/4FJmwwa58ZMN5XoHX2ARDrKUo4e3Q1x8W5H5VLdxmi
/2nUat0KdH+wuCPdTgGsEV5/TYxr+pQFZHPIoHpWQG4O9s1LKvVRrvv9aFmuLGmY
`protect END_PROTECTED
