`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
23PjqMDsT2G/Qp8KA4xJcVUUnTDDUaShgEOggiLz7F3FjZsmyvkLMqel3wDXBr40
dsoYg76VXKQP3PcVj+QWBIa3lSQmTCsN5R5Owqc3D7snjpOunWBIbnM8C/vyMylL
1+V9tK8wAa0I0Fw6rSGoXL0Ngivzqb9I/TV4PcRNDA113nigWPhZyBNlq1stIULz
ZydmOYX0e+8MtGYgWdjsUkgIJApcBJ5X+lzbTOqZwjieuXafB4oyATDBVhI1L1gQ
GGLzxScOX6YaMa0oRfK7c3jxNEyfaoYsLI4AqjSB/rjODJFrVNuXrPAQPmxB7MA/
WD7XKvOMvYjj3lDpahcc9yxY+R/n2hcQOql8FUxbMACkV7TdYeb0REAhpR8w7M8W
w1rM049VD+JqmzJwe3PXt4bRzIMhQ03XkLcozqzL/NcowHtL0vkjNaBtdfyox1k2
SMcfwieDzyndTn900vL/gmrjTF6WQ0VVfJgaWhVTZ6aakfTtFRQBxVkAneMk3q6i
6dniTIMghsOx3wtzmP6YpXk+lXA1Sk2W4VeVbYK9fQZY/ObEU7aq5t+q8qhQsHGc
WhZ6eZbd3X72qjWeTdFAe2+g9fHI0HkrJ6/AqXW3eONKGVBq6DVScgu+yk3X93wM
p4uhV1lr580lgjnhluyBOekeg9dZRURs6oDjAyzRiWt4SznEPG8G2/j83vWMZSdC
V2UwHUH9sMO/dJRUxITpXM0GVpOH3Wcamn4+fsQVKDIP5hhCC8sxz5PlK6yDc7u0
w6Av7FUfCMPm9ybQf268jza38SHUD8A90gOjJibnAHaqiZbESgWcv7dIDBAUJu8L
cKgJVuWG7S1nEMRX633FjfZ0UlzeBPyMR38WVDlGvVfhylWOw+fWTO2fwX+TZ6QM
HzMPW2nktm1lQpGnVErOyz/jOPJE4cpQ0udxnGZk33CEYRtLSg9qCCJwRUjOPmAv
ILneeF17PgIo8Lgj7PQSzIcZANDqWQhFuYQiVWaE+XTx/rbnvPcv7FEt9hq8xbDp
AchYQxydrcVG8yIZrmn+G+k8IkGcbV+niSd0Vlouj2JdHf1B1kJFJhS/B7okegjb
dVydzf4vd1yGSlmttFy80t1+8vAKQqB6jXTGxciGTCTFZiOyE2r0QSCztr3xlw7e
srzAhEk+wEZkCr3G6taG5ULsM1Nx/TvKEaOOEWDQJsD/y0aBFZqbTX1NHv1UUBEz
4ExOjbYu8RMVV1eI3qj2MUJyw+Tfbr7A4XVEWH8gfqplRLho2mdat1P+ll6brm9n
f1Bi2a8S0HsEHy2joipPzCtxxQJ7nnbBa3gA38jIhb0ioGn1jjGB+84PiaFd05HH
Yp2QrtUlwQSL/k3a4xfuTZ8XjwXbrYz7uzherQMUqX/uZ8Z4rm4K3esBI1/O1lhr
CD23IxglgeuIsabV87cAVYWAkknaUKABu/wp19fPVSGfSC18HtLMYY8PcLcuE4Wd
/9SFPri/yf2X6JhpmI1/KszDusr+W7wa9pgYys0dRO2xyvPfhoy/BWfajtjnSs2o
TuZbJH4cPJR2+7xQC3/yTfyNLFePEnNS02l4fry/Y0pNQc88wdRAqSfVIMMP+J8c
G12e2sP0D600tDJ7rl7Vpn2EKkoTMQ+cqv+9Jauhz55gCF3xbL1lfKacuih0+/+H
QuwkB4WbyumrVhhFsUblxw==
`protect END_PROTECTED
