`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wgwk40h9+IZN5X2GILbc2Fjjaa86C8E08vSsplQUs+r0hM+KTzPaWPai12LrYNj/
mhS9v8VeBxLT5F+bWtSUEbOZRpAKEt+LUmvisoUT8ZrJgCSmjdhhl6nbvtal65hv
k1DINiEs4WJ1pPPI32zNjuCKoFW0LN9jCVqwXZ5+9AfxwgtHgt9ZQASu33nSXKMS
hhAuyIpV6ZKHsoUlDxQrOUtVReWGz9yPalgq71xaQ4LHHUpf90Gidn9SSckpLN4V
raYvoNFM0PSK+F0gv53OirPDv8U1jIc6XFdAHmnlVvpeINGeRH5lHbDwsFFXvEiv
Fxpc9pUF6kNHDfR+PfXexg==
`protect END_PROTECTED
