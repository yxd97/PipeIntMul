`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uYNf663DeVU3cwaqQd+TDwwuKtdm/mjMEXQRB+dwTvtGNqdU2VYscK47bJ0M5K9f
W7ujLmsEXPOpqoJ5ilQEX3fk7uXszjn3VNDtAfuJYQb0rgEafuLpsHdpoMhCqjOq
dIHY+IfMwscO22RSbQlWyOtC/Zttoo3spFd4APYROF9KBtOW9vlLTrQphkNpiE6Y
daQ9/Kl1m7V3FEbcL0pXg/Kn97d/7gHNXQlm3I1Oo9YVXBrm3gDv5lFwtAOsqwBX
b26p3G+Nc4z9McY05B1omDN5H8BeaQwBbberSzWDqu8=
`protect END_PROTECTED
