`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiKZnRZtzUFgq4k7EnoeN51XNlaWLANPJ8XJoY3Sa5Lhz/ziXB7t/peVgWlTHcdn
ouG56gBJOpGmcaGDqrYabGWOT0lLIo3bwTPKhuG8ybSDKGZbiWTLArCV/OgJszZP
ETecbHl0rdQEfg8V6ScQzMRpuFHbstvAhfSzf6Wn6AMiSoKZpAJsPDG9GBSeJ+Vm
VdNFSM2UWaQXRkohaVE90x2Ken0kSdLdcbCwTiYWEy7P4xG6DwrrwryeigBjRR72
/Tec/o+kBhCxen6k/91pN3m7L+cPjFecV2iw5j62/4RtXrJzEuxvJm+W0jYH4aEE
9Pg7hr4MEzdMwpvWGHXeJS80Q8wuTtBWBYkFzvW5CrG4ln3xYmhbozYdSLgbSu0S
Mbh1BWFY/2OIHG1w0ADK6qcmbnwJe/N7DdhABSNhm+m8G8W+4B7YdOf5MVVZAJRM
KlFhWsrzFWx034TNpm79CIsUDmE3tVx+/YsulLaCFyHTgUnOhlcoxvbg4GYF3uzg
416pl2jAVR2i9xb7vIR4ll2WKLyfJ4tyKRdP47LwjQ2gCgIcL5SOgYZXPxzdNVW/
i/4d5qEj4TIqs1LUFHs+9c3SW6EwpPp7Q8JfKokHNk/5MZRsj8zyFKbsX2qDlRJ5
e55K2u+/uJCf/ZMmUzorkgWc+93MFct1SHPsAXkhglZ915o4jyGgQOPX2T3eKmJW
+S78vMdPuCedcVfrMm1OHLS9MOE6tzSsbLV5imY2sQSeXHSlKmppZU2+IczauqE4
gN6i1ThRWGX3eYlTPc4oS+ntCqCbVA374pZCzut2hpHxfENlnzfje7GJaTyKQqTo
6/kgEMJoDzGI5vorcU5WieRY1epfZvgH6XMcWkCra8xOtP4Qoj5n8q9Kq21dvmdp
isiWr57o++rfkP8rVbtWz80akwiLbk7VVpguA20EArxXVEkDpufmQzHq66vmWJR4
uQM0aM89nmw+uUBOZIJSdLR3/vdkBV2Nl/bZlDRdLkBt/clnqBab3RfmUlQY7+DW
RnSOrdyHfJSmG09uKZumuR8TH9S7l1wJuEutRIPckaX3ZfXa5M2TP4suRTFNENWd
YXw62jGICbTLGATONlV2gMC4RR+sFRdg+Ei6r9MyAlk=
`protect END_PROTECTED
