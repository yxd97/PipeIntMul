`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oXlFSQuQC4lALBuyWRcJX5KDg8GZsPz16Qiwe4S3hLi29cSLDj0WkTjfZJLr1JTS
jCe1GYgphlKake6LGrDfJyuA4vce54MhRkYkAejKXujCNj+wV9K1nina7O6csjIj
sYH6ifbV4+wRGNVwjDhBpGhyl+WLf63e9Paa4v1olt/kWg9WWHCttTg4YPQq7Brs
SzUODP+S+Qhh9VDU/wfi/oD1c9P5fB11KriFgnVovSzImgdEpTzbvWqXbIfFTcvK
yUGxYHFn/N/M4Vh+uLUT+NW8tIlAo4CLijSU7PXe084a/bXrKnbe725OUUWy1zEA
IXAjpTX9QPoOjPYKIYfYcXKXlenEg+icgPSFoQE0y3CnEGjr0oJhtVNzlA+Qyern
p2K+6vvWJAhRlyPpj+ifsqCl6WoQ1Zf0MIZBm6eR5akwP4+NK78cfuPfx6AKubu8
96jHSpKa7w3UZgoWZRLTukDos2R967cTYwzYTBIVTFPVkoG/w7KOWvyALaD4Adyx
mlB+g52skwS1Jp2MpolCtCDqjU3ZrOxh72kWCmHdqx1RlsRMbLuOakgYObcnffai
Mnyv0ZvSLNC1eeh6gwLGiFY/lw0LyEeYNMp5mesw8PtpZOvNjwYAazME3h1ln3Y2
lkKVa1YLMa8TCRUM11+casr6upXA3bfsGprK3A22H2A=
`protect END_PROTECTED
