`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p01A5m0RESHR1pZDjv7YvofiIYCC4EpXGu7XmoyYM4QtOC7EDIqUBhH6fX1miVzI
mqZSvquAK1y4zm1mfMpJAUNqSlIWmR5bMbKItcosFfKyk1Sf3mb8d2JN6Hd0B2l+
k3QIwRok5vzIaEtTTgRzVGd3SIVI3K4i+/z0DZRb/tQiD8CL4vr/N67MU0MbZRNx
umSp5VDI2I2wCxEm5wclX+QheFdfBEAonmuYxvjSRjPHbjsFuD1/k3MwHYZI3k1e
GJU0vWs3U9OEBj49UFZlYIthj/fDme9g2IAEiAU4UvqJIqwzG5uapoPvLkgQjCzr
vWDMK+9wNX1234GSiDK1cjlExSFx+e/JGvzar75Vz+hg9p4QxtjdmToh9tYk9w95
7He8vZ0bLvgDRhXV3o10Sejx9E8RvAhxNmnkQeflMEWm4rAlylbr28DkBSGx+K/x
sBhP0PjRKfy10kxEApWuaeUjpCNSXvZ3PSSXYhQL/QyJS+pZzvdZc354u/F3QEO3
UzlQTRMpbALf8oKjOcX9N14dP6W+4qKHSMF1YIEebE4qqT5kpdL5TwEZulKBjOiI
+RVpcFbd+JRAK0UdqOJ8Yc3eGwRa0inKiyh2jJ86r+CYYZtkR7Tu27AkWyeV6k0F
X9FLabKMyMyh3GOH7/N2mA==
`protect END_PROTECTED
