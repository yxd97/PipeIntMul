`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tW9dD3kTJ/2P14NdashBZ4FCC2unhd0GKs8R7WW8OXEfUAehkPNfJHLRyXvv0O5Y
eHTCt2qz0+nnMDOibMD9lYMlN0aU/G+E5whE8XF8XgCQH874GhzfJ5bYf/RO48fy
EiustMtz9MlYqJe473qfSDH5dWq02RdcitifH0oo3LgNwkUnEZshGnVU5lt0Vx6B
eI6ok+r1mN4wFAZ6dQNMybMoABIoueGuuzT5CyEuhyi7N/0pRWfamFt1vAuQvo6a
M4F4oYS03qRfipQPE0MVMCyYKPbuxJF9OYn/oiG24IP1giQbeNByBzRp5mrBHa2+
GTJrOcCOMo5XBqd0m2UCzQ5WuJOXMeKxtucBluFx6S13uH0d46qaBgJHLoQ1p7Co
DpJ4LNDtuVE1EK8PilcM0h8JLwde7YMS52W+6ZCzIA3g8z9kqrcgS5cMtg+g27cg
`protect END_PROTECTED
