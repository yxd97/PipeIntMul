`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uZG1eWzcZAL3MK7wZ+Ky4iIQMWYrSENJmn+elcXQlU5A/+xrMgz7mRQ6+yxu7iq4
RCBAJCPie6egNH71lCSz7l6LFBNg6XuegDSF3PZ5qJ1Hfjpw3SenilNikRcIvHaW
VjMSkeeUW2Uv+8S7FhXTGeLJNK7HoEzA/SGBVPzny/9vt7Vhvi2zCJfQ3vw7S2kE
PpJTojJfGtkF0ihY6OX12NGBPmAFXTLYcHwhLsOq34y6zSRmQ8v+YEFb0H1iBS74
JBqwTyHJTJvcrFc8tS75vejabpyJdd8z3g9eYMCjni45vJ+FK77uIbSJW/UAywUg
TBRI9NIshrHNFB7yyGQmtfwpS5Uu5C+bqH5tOVZDi+yaDLWfkWsqPchpL4BvSFk3
DjqS6r3mpNrQhGW9hzUomDxz+n+oM4X5ntmy1IDfyDWUo1YBFWWLfEWGDptmJpib
hocYe0ASIzNLHmmG4Mo4gqWSmzkhdS4bGgPeq0c2xjhxRlbaIMV00EkDIo2VbaeH
Cls0cL/yYQKQ55tbLhmjpXkwnFinRi8NkgDPuEW1gWEOkxJN7jPTlxHg0im9vmhl
L/YIlJrWGGeTs+xOuJWr1AgNisRIlyYBTo3pgxdDuR5iW6TdZwT44kKoGgVqz3P9
dbZ31+6MSSrCla3PsvzcxdNHW+hsJmtoqYr3NJPtp5EV2Ycc5EzRGu1y8DGJVrRW
CJGYZg/3hXLkC2gwokKLCoR/GGpfgpb1Mo2hy3+OWGS7MffykcXtMaradWAMHAA1
YN3ixTQR3wMAZxKEdcB2D4xQ4Nl8R+6UU56BIhYIiUfDCdRa/6wCxgwnM7zFi89v
eBg9zNoaPieEIFihZXNOFzJYw6RSAdsOQlHqgPP47orBifwRbwAaURLfuedrZ15l
Obl+HQIkC946n0fZeTYn5Hda33pEZX80B0Eiqa4JV665UVI3BcDd0S/x0jZagPaK
4aKjPoG4DVPNiDX+o5l0rwfB2HKcG83Nfm7gQsATV6o=
`protect END_PROTECTED
