`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
szxjqq669w9DMgwSYVysqxqJZ8GmJM6vtCjcfPKOcm5XIbmFXlGqlg3RxTDSznNd
/B0XqQ4bxQspnr7sw9byCTynLOj6HsZ+DuTNlMm8lQuAp8Y4TNrRVsV83cG8mYTt
3KCHoMqVASBM/gitPg5cOwAyirsSi8ys3Q33Yfwss6ZgbfC79OY2LAFQ3GF29O0+
pKNlSakhPdbDX2oYwgFXiQqU7lhBcIsJug+rKANvCavElQaYgAvqJl2DgloZaLhN
NmpJvJsUV36N15Nqqwm36jEtFpf1VZZQoLMedegKvPZ2mFMud57YCPrUk3Y92V6o
18rZe7qiZwxnHi3uvexHnye3Rxv7oGcCPE5bNtQqmghojJpMfvJ58pTgoATjaMav
NsLJMihcAbBvvmjUBg6S3uJiN3iJyzKiTQMmy/BwJ5RJgAnu7c4rEsIsoGTKWHol
LreHTVPc+PrRA8T10s0L9M6U30HB80QOK6dVxJbYCgOTONnHxn7svks9wG9Du8SP
J9V+L/XFBZuzZEfEq7cUmR6cGh6Yv++eW54n8/V2YZesVI2jLlIeOaMEd/L42Sml
5Zs2Sth8NGsTnxX6aMFFVa6kULfoboBD//uGfsUae1nM1XXRixAKpw4FosTMmdV1
wNXOW8wMie0nbaquZe2xAIwSHztNrBZh9v4cCPZqeY8V2jARpl3gzPEgZ2K/yLOh
ycaRCss7iWPXn1gcdq1ObkJzlHT8jXgGxU+pD1xKlejpOw5qXIfPrP9bj0I4eTyy
02kTGERqCzufCePOtuMYXw==
`protect END_PROTECTED
