`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6PkopCX7z+ioTuTX9DMlp9D2KcBG43kq6NWH/MQRRX2lnRm3rZsPm/sKJPIgaNUD
cWvh/aofFrAtbceAO6Lf0Mwm+GQyTox+Ut5w1CzTOTICrFitX5bW90es2Mu2zrpw
mEugjDZ1McD514HtbYNfBVYdnUZw/JGEmDIYI7Bic7uOUmUyzAo6OI8NRcVa+XZR
sHai9vqEgubhH7f55Ry5fICUik7IZXK9GTJ53K8Yv1dN7CuyA7M/boQtc1NXnLds
TtGuNPBF/HGT6tFfCnz/y1ujS5AD2VHjSkgDvORzRus5p4YFx1kN0gFEIINOh0oY
E5GWvAme3A7XBVSq0yeVLXoqDnN7WsbZe+opL7nAJ62IWb1agrwsi11k9zoXv9HA
9vRahIFSwq3PR1b91P4zXoMtTrJEUlEkPF1cF8P3XY9EUEMpijkZUdNg9QrNCLUE
0v7YdLvRpEjD+Lee2AdjWkKIk6yh8mpaJeUit5+5Js6XgjRb5zyPpL8Jl5AiOQ1h
ZPr8YL1YcQvjRXS02uFE/U/Q2mizKhKCteLz8sR7GWJ3RHOLK976YZr2Ps+1G0N/
hUCpo4xUzbKwZwcI/SNJ9Iy9tG8E431VvAbg9wHbQeJE5pnRpNN2KSeUX2tJAiw6
wdm3MqsauXnkfqW62iFjVzCz0er7Y+gHwvTgB+Lj/nUz69IfcpNbpRhOl/JVotzb
U+aiffXW4FcrZfRavxJoO3MJSwoko1J4CSTO4k+QMFiDx8EN4BMNjlFsh+vaCipH
h5P85FnQtgjUTiC9bHmFC718KHt8xFuB+OWi/8tOuApzmoCZf3Hx0E5xBiBCGtkH
v+0E9izPCwlruLyFXhyqXJiPEIn7ImFWayzkCgMwhrEa/0JaXUsh+gPzDSUFexvA
+DiA7iwqPLFotytwn8K5/xMyGmWGLxcwMPGCz+yT8PHJudczqRHb2uP0Dqocm6Af
l4c1gCLcwIdBr9nQp/+h4nVbKy2LUGfppjJXYihc6q+FY35hRaGAb5rPo1+UmTnL
msIe9Jv82mOAHsV9cc83Qn+m5WWzx11lSLtjquSX5VFarqXTzY2xaUFTm8tGrKLM
Lrhi4FOOIllKGTWptAvPFPAsYn9R5cQX0VV/kcar2opYQSMGixyaeLoHm3tuH9Yl
lLpjGKojTpiABigR+K2Ucuv0k824p8hd17VJn4gi9fcX/11UFzPcB5TH1uYmlfAV
TXzRVIFNVdyhsGskyemOveyrocaPiWlOi2lZ4f4vY8SNPDFXlxTpX/f6Bks5ox45
NxWReQTQe9SgoI9cf/PUPK6cKL8ie6GwwIggAa9Ny/G/JrSiuclG4nJrtiOPajfd
jr9JQC8Kkratx5xP56VOu7WE1iJe1P0fKgFA2hjomACVKTs27jSYaOyb38Du0Y0G
YdU9LcayVVKnl8V47Hw71YEk8LFTHiLnIhf/DBuh0jIvqOTAtjqG12CM+kTJj1d+
INripy0KMfPdyLzr6QWWKMsHzuxfWBn1Za4Kn1O5dbKdsGrC/4/r04NyA4ZOvtHE
t+U6vlODVLDSd3br3pl0TXu8+IAc1yt3+fZc9dDnn++teWGHwGWUVLw3d919oODG
qR9nRDatyD1G0xnSpMbWtZ30MoU6xWLT0hrGn9HmK0tOzG6RvJ+4S73179410Jeo
F1dmvvo/2mkOvSM6PlS6s3LkVGzp95/rPd1PPfkziWy4L1tsuQAwmQ/7Qqw3UjRd
VOMuXb5MACluAB1umM2R6WWz6WYK+N9djXq4RietPrTa6P/9Et+4aYAqNtbm4q0Z
vS07b67TUpbtRqpythxb1BuC02Dxvq2yWH+Ci+WwRQwlG+W5U6WuiDzzchncDPnk
Q7Q2URaMD81N/TaDwFE+94g+a79ISe8aDt2nuOucYqGsNBlLOsWU/yByHxF/ZMWk
Th0Cuv/LMBkUD9vYxH9Qri6wqNFv1xDBDqfPHacBzOtiVzDX7Ls9aJkI4bYCpWBG
oJqnKhDQ2TOEAE/7FIkryUcyp1GlJljjO/XvHPdJJaWtm+3waHXYDxXYXBV/IyGE
rk2rH9AMtxGrd5Ev0LMfsj3ncDplsHHsoWSMor4jV9PQOttvCawNQEHHA9vmAuU5
a1eRvguaE0F6OEgvl+QguEI4j64SmeAcqLWuWG0zl4ylnB/2Amm5mhySDisorH52
Wb2Miwm9GFzyQJ3MDuyOD/ZQVVE4d0GTbXjixpU2oCh/jFuU8sieofomKZtasrod
0IM/IEzKH/BVgrn+RYD1YtZJDoJc5OQrKX3ID4bSJ5R/VXMXXbk7Jr/KqP/YafXd
P2MJ5YX6q3kYj9kLRivojOi8Y0y062sRdp4DSDNUdBqAWuh/Ira6vZx58XNKaAqa
GAKCTOA25eFqxRtFBB8XSGICqDNrd04ETNs1Gwdyyu2+yS5X581f8lI/ieyMA9w0
Icjnh/XliXhlhmVyXEet8zYRQVcJRdoPhy1/YaVgc4+P7JX89+qD2GTwAhmiyL3Q
yViEEm20Je3b0glkT/2la+1EtXgKZl2IQ7RSY2fUwyWAc013YOViO7jyMQuYUxXb
gXPc8IJ6PENLr89XKbjmHInx+Ds85Cbbw25yFu3ZtCtMb679+Z2PFRiMGs8yynRt
+a4RSbPFFYVZANfrGfkMEm9zS8/W5YqG3uzQdfm9FXCAdLYjwdPg29J+J/RIL5ud
EBBo/BQwvfofJfNa46Fn16TLqzVVsxhcAXmn1deFl3em0++JtQfiLq6sw+p/ln3S
bAGm2VDvaoipu7GZOMoLLZFsgd66rKgqsOUub38egOnUl3moOFtTVmNXe7f+bI/T
ZIZC5crQsqz6zjAHjjez5zFxtTnifFx/KWj+SbUUQwW1Kex+pnndk2Z8LhlYt+zB
bV/H7Ko9h763xnIOB2QhBqxtb2Ihzvf8B97GcieeEBpVOeb5NLRCX0vPUE/YqMlU
TWmKsZj0z8LsT2uB+ox250wyQrymLnjEc1KS9XGEO1n/92iTjy4xoeG3MFBZKPYb
DZXRplni5qMwFSaV5Z34FhecaFBNGP2tm1XkUAmMK09+BC4t4F6YICYsgEOIVQmE
aEWqkaFcVIC6+VVkGH/g5Azb4hnA8PKt3fvytFut++ruWaDHUBPdnI4g1UhqBqIg
7K5yEqm915vlk+ocQzEB3HuQvPQTyiN937LfjM9eLG/om+gxGKDPXzD/mMVCVfrK
VmOIOeVlOvbmn+/eQ+eMVKv3Q5s3eubxuwKC3hdDtFYc9QwJjcKGA2LJThI04Vy7
2Pi9+/Ut29ET9ZWLAJ50ZRLg7ryJ0FUWxjVnN5gvnjC3ivwUFnEfhgzO8hh48ODA
bcRNfn4cPTE2iJsUGQx+MQaAGLExKViBBdzwqIDZ45XDXm4JBY8YA5tF9lOY5lt0
emhc98Lb5Q/ZBL27NZmNzt8smpyUNIcpq2XHmljTNNg6pbBNmpDgftuMBODhGD/n
XkacpU4QAY90OJm1g0j0lL34Mzyal89Yj80YqgdJUkoBdKsG4Ed0KdnmcWpCNgrX
rd1lya5qY1pJVceRpdDk71opgNyVPOh1xHCywkrrvp4r/cY6LVtW9wRa2sll6TAd
5rOMrnEx0K2SathbraVIDgymINEhluZwKOh6JmKw7vWe89EmoGu7/6jZViuD/AtV
IaxMih0KC8TDY5bs4ZuExwMS5OAc7fIt7zfKIwH0iF1yqC9/F1WniB8xpg80y4bZ
RRI8Y9OdVbvOAW7ECL4wEDmeBbVghIyPVrV79gR/ICDozhoYE4z3CcxwrDFvIROJ
8jJUnzyUYyaN1pmnAGe6iA==
`protect END_PROTECTED
