`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIHLkJlj04PWCIzFkd7qPN2f4nZMLOeQGlXLVy+PiS0dx8Plm+/r7IgkpkPCqTSX
cK5w33lAuVJjWAe0aWoIL6HQyYPhHg9yyUihmIbtDpEj1bPd0mmAzIWX+CGvOq0E
cAzfJgP0QsEFIut3deW7pcox7fe0vHHpc4SGOuflDA4RpHratA7ov0axaqaLACmw
LIufcZMn1NOhknioEAIoou0q+jXx5/JxjYXAklMwQmRBvTdfsbs9wDwga1KCJybn
I7KE2FCFfau0+6RhllcRC/YEVfS0x5yX9wXyFIBqSfeIpjOyb7yCKxdhPy4WEvHd
sVjMRm/x5y+pnTO6cV5KqFJQvRSgK0gL0mGdf6wuCrKGHcc8ryVc0QVbuVDD1NBO
`protect END_PROTECTED
