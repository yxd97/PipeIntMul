`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o8SflDqT2Ng3mYDGqMZBO5sQiHkIBLcPDDSp703SYrvTJuKQOG1p6AISSuY94f8n
UuUoWvqCuzQYYAvtL5z77mLbYvOdHgp1u27wE9YEJomrYuIfv5PnGqSrDFSBzmWM
gxXzk9WFANNdtk9LXzk0Rs6xIhjNxmGTNoO6lp2K5Q/9lMA2+6qVqiXohHAWfSxB
sNrjE1CbDNaq46pmhVCN9oiJ2JBQuF2Fl9yyoA5aTo5NgeQHFYdQL8S0F+bahpSw
GtlxoqkkwPYcTRHQ3GkQA1iqgS5VIKhGPKS1/OA+gM3Ze8iva83G6uJJ3Awi3zpE
zUT4N29rNWtp8uW1XJ3vLEhYPyZGxNSO6jEDSy02oqVHFtcmjJRgDl00Gg33juYm
Cy3Pc6qW2Wu9TUMFb3Bxq58P0IMZj/IY3wx94fNGylziRtCmEHw5Am87lau4HaV4
BQvUHJwzXtQP3pgAj/6MeS23yueR/viAa02VvFcgyCIRdGIxi2Z4WdzSI5to9CLT
vkGYb5MAe9a/42zb464b+2vhVQke43mUlXH2Gaftbp5dhgqjfN8gKLHN2IeXKpRZ
9002ffaa/CL523ZOrBtptolbhaEk44GMB37GVNmVZ9k=
`protect END_PROTECTED
