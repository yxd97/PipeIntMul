`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W3j7Gfu3ED97BCpwGBovrHk3Ri4T1R1onHDB4E6os+PTG+bX7sv36r3IVonzj5g8
p0IsBaRD83RDK7HREUSRuG+/+fy/EVbEBdrLhwBhAIUuJI9L4ilsfH9Yr2RNYgzq
BpQ1uJIEsrChqVhK3p0oc8LlufvW/f0UN6RbgBvjIst5znoX+tBADLkEA9uBnAbk
RXxg26ouqB6PzZQdBS2xxBkD5C211e/lW6wfH6Xj3FY+r8DTf2q/vieLyIg/DEhT
hCyFKVKwaYpPD1FVNEF8AFU4lmTXIB9ppgt4I4HWaCbzfPIDJh5Moyva7DWdLlff
gaWRKN/mnh/SC4i+7ZAVJT50KFw3g9g3uR1jvPOIrC3dwVgZcaSPMmVih/KGjaSX
V2d18cb23h93KnP/6DT1tvxD7MxbnrkFsloqlMxJONpBHMx2fcys6nTYrcUnZaVI
XQHARkH74ilyvGBYVEF9v5eOs+PvfdTgTi9ngARjavULIIl6ghd3aVZZHXzSGYtw
8605rXn2Q1EBWcq8Rb9oxI1pDpLRB3pOS+3fn2uL7DJRBCoblFpDJiXAeabEc8Pj
hL1LhH7x/38S09MADfivcpMekQAtFr2lJaJ+X2QEwNhWc7i+0HBc9tnQbPBWyYtz
UEgamQpQP9Ibm+dggcrAXiZV4j28FNG2jMwkB0D+1B+qd1oARRKjzky8IW0Ca8ws
gFQ922N9uDn3f7wpZcEwhvsX5l3/a4DtdzUAAzPzwvdqe7TsAETRi3oYyiNx6sbr
hxFf3dYFbrUWD8kQvEM8SgAGDlYV2aOAo/MsjbMqYWVDh7LCYoZvtdgvEJ8lTET0
Cr+AWMVmybqHT+AEXKpKINRJBul1SeHwsfLHKuFcXixI8UG3m+YCT+iqBZFyzSqG
zwjP6Dc9hJyOjjf/PbSRr0aNbn57AkAcjVtbqnN+/0ERpTzqk3TeyBjAzVJJqr4W
GtonRSOE8BQ6YNfqdqJ4J2+EwjeSBY2wn/MvW8gXkUghutvEpFM4prphcfJhJqvK
NiyggPtsuEfzuaDdRiAQ6fcXlGFBbzTaBr0/R36vKxzMeL/ENo6wKSVwjl5ysKdA
`protect END_PROTECTED
