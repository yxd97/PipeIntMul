`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
umUlEi4erIWD0CW+rIDtVwkyzkHIpe9DBYoegrojFY3W9KROWfSWJaq2sFN/Rb4U
CMc3S6GqsxQDiKWtTB33+XmBWdK1tLf2NcfTvOxmSYTPW2XsX2AONy/EXm1lHYfP
4FX77fEcTpJrWJ5fwsAW4LkIRwpuGqX2i7QkZTG7PjGNENTeH44YPJkimVgjHhns
agWLZvS0Wl2hTHCVjxn1uBS0wMg2/d8Zy6y21djtkkz67ty9QXytd1r7ABKb+7ek
9gjHrvpueRmHqLz0PBa7gFOdOQHgynM22z1UJx/PjoM5Y5D9xDQ/vaTVxjl/PRFQ
HWMbizi6P51WMHkp7nq8e6WxQhf6y729OS1LVrX+NSY1yvPk/VlkE5YBe0O4rmK7
4B0+qAyDPEPFqO+/2jp1ac2ZN3f2mWAzEmIBLPYrn9HuU5vjs95g/3/JyiIbK9wK
41G8TmSfaMAMr2W5Ia99gRTmVhsaBQm6XbAu5sA/sl7wSJy9SqeDPo7BnFy6yK60
xB9zjDMgjcrjYjzTj19ttzBi4Gy11K74YSgyOGw9yjPdyuv8ETnRTsNqlPmGQtXB
iAIf+4KbUs92gt4id/n1DvlwRB9eYWWjeNrUcV9ZjVw8UIquP709mu1CqU5zAMHg
GveNNZB6eznrWCTZlCumB2iGDR682RoEV1QKICNyBgZPPqUlRBGYw8vZbIp+92RQ
`protect END_PROTECTED
