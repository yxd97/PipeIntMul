`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BSdCrU1VXmBVUH8ZjMQopj7VOPpWeIjcejf6lA5QoKt2XtCr6GPtlh/cNYSnVn8E
X8+ybxmUhFHO5XobL6qM8LXe4mDdAJp6VBLMqrJikHjLy3mgMZEl+ljoVNW+6ecE
cS5Nzh57MFB3CPVF8Bw/TvpZ4vnqjKg9oJcsr7czMdVNTgh3v7NysAKFnkAslwUY
/j/x4gmdAq2UyCX1Ux9MuijKtl1kV0UPBjHV/4UufynN7MaBrSpyQJyOzgYj938j
5xc44dVwl/cSsvoJ/YEpi1WzI60kzpFYTip9ycbZMzUNXqw+rNAIsO6yzzzg27wM
pte8rQQ/lxiOhRnKyXKZfIYTZQe/4LPHdGDcToabGOI1Um79NQKrMOSLVaaFxzmR
XYc4ONABqW1giEw6oBPtbqrM2WVDrP5A/9oUWES/3El8RrBW3Ocvf5dT8BVF2X/I
YspqD61GsMhBf2CnUTe//BqR3uStPwWQrTWa0s6Dlj9FnTdk8nSjq1+O9VycHs98
2pnTZif09wgNU8J50l+X02efd3tjpj17D5wVBLTbljkXnuKYDTpnbnwawGeTvIce
oJePI+KwsJe31NzLwCsCqqxthQahT/wFzOJOb6TyZknWHeye/Z/4p4B7QmIkQEaI
5qw683+EqSGXblKVIVhD7953HppYn/8KOm23A4ItU1g+17QOXITyEl8x1gKlsQNA
Ob1nlIYyklyuF1+k1sPYf5ZwpukxRHbWZRhiRSoA9+9h0ysqt98o7D2Wa6MpHTP8
leS+x2/qQ/wAmaZ/Z1ucSjW0/q5vgQ3crcStAA1U1Qn4df6Ze1gaXh6bEi2w6PHn
uqwF/0Id7gqjalZA0GbUftlxhGmcnKeEpqJl76xULeueHsE0aQFBjsDlEGOASALm
DPSAElX7/d1g6Pxo8w56SWG8tMkghDvGyJkKzappM7puXxSvd5+HbXOlFvoNL03L
34iHsT0whE1EPpMoyfQRGw==
`protect END_PROTECTED
