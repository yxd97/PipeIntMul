`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PCvalrt86bJguaVXlo6Gq0QdzwZqXFHTfufMfFhgNd9dur081/wxu6cPBLq8FX67
ivqTpTcZLFgvj0duezqSusq6XmJDfIdKL6qpoWoz1LVus6VCcFygWOB5wStUdpFA
yHYlenMC6kg8+sKH2OWsCDApjFsogTfRdQ5aeAirGlQQLIMBnOBwscuMMPjvP5Ue
m95h0fssQDYJNC4diOTGu7hghffBLCCMU9MNOwF8TMczyo57nnokV25vJw3HDXU5
nmvORMML5IpN8R1Oj7edEPeZUnaYR1U+UCNi87J+n/1EYL1TBdW6Oksf1CxZ0LuI
CCw0E8hv5Oobheg+9IPWGkG3fvDNuXsGT45lGLDgstdd4PCmlzZr+t1AbVyH805Z
8gmBxSt7av0gNRg2nHRqN4pCz1Nt8BxWbUaUgrdXG+3T3fp6Ru/xzHy8/mXZcCah
aZYKfb+4vZiMPOuNhJk+5b/Ntytc02rB6yGL+ecPIz/xm9Fl1kCTuxgbCcMOW2cp
xWhaksTjoiMraLBzzcIZ5+NTI9YwKHFiU27e5ekCFWp8xi7LWrzNGUtgN9wcEcRT
vc1x/OPeMblHSlHLdEpBO6iuweIpV0Q/d8jiAPuj5X8G1IVfjU0F6JhOI40bw4hB
ZnEsdvMgFaIeBHk9V+aoFLpR4QPvxvTev/ynHy5U3MnjaUP++PHCKKIjvQJstMEk
E2VuFDzwRgCZcU8wyDAodTSobGyfsDYO6P/4xt7sdVLhgNgNOHM5fNQQzoArCBdH
uw6MdJbXtI+7wrXx5vFBeQPUsrjcqS26mqxdG4s1RQJzjeegLmm1NujPYGeguT75
tObPrwXuZ7hah0GAVwBoQ9A5AAEfklDPSokpBufbWQezj6jUxFTgK5UC6UQ5+JqC
06dIxH1QYB+5x466OeQGuQ==
`protect END_PROTECTED
