`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1bNFQ30EUt5FEYnsUfBsir13UH4MAiZROElm1pXX6X6QydrQScm5uawiTdaDmv9y
wmRB00+c2eIuMW+DSwqESj/VzyIRKq8+c1GZIM5/aSyRslljltt2XnY+sP0vG0hQ
zHZNcGODs4BGfxfIddQE3lHtUnWKfovhNQqXfAJdXfHa6GIveNiNfE8GyB7E9e44
zlxBQYRp8cvV54uNSts7rkOmlGxT7Yo3gY8+oVYuTf7AwGW7g7EYj1j6n1fWhczo
dmUBG8Ji1FW0TLgH+2JU1ePM85m9KRSIhojZUrdagKVtS+BUKw6Nl8gs2Z+1Iylf
nSXTKU8DkJeVdHb1LX6p2Q==
`protect END_PROTECTED
