`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOFeQVDlBKtfYlpotZRYZcTLtVn0jys/9a9A63HqfKVjbtfN2+jfn5R031thKvAD
mEz0GK3Izd2RuI97lniKUGnNNezSwYbkE2cGrUUmsVQ5hYodXWmwCZzBBNMzWXMt
1RdsQJla3dsSq9rONgWHGZceBvPnK5z6HQIFpsPlU/uBpftvCfJ+OnbPFPH+M0qE
3M3vfrHfNj1LPJmj6PaTuLvRKH/ENCa3qWdov1xlGzRCbJ03Aq7VWRGTq4DU4UXl
IG+0aCaAatdk0J9VyVef8Hu/SI5q0jNtdOKvb4/k7gF4AZ27uAZVk7egM21Pyt0I
F80xofNrN1SpxTzVk3oJBbPbJQ/9+Ht05IHgKOeYk7mQ0U9lscdafeRgLCsofm2/
wqV8INNawxRl9vJhJDHTW4k+A1N0xaQk6FUX/veo0OcNqJmZxXvBCyZUCb/oK0v1
6H3DbL3E7tVnjvYl0W2LbLB9e/CEs1f9Z1/gKz2Iw8Y=
`protect END_PROTECTED
