`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FWzGzTle+i4xTVD82M8FDNkkye4V7ei/S/ZOmi21/Y5BQjWq9SmIQ8xPX8nSoW+x
j9uyqAKqV6X3mMuQWLcRyfC2t+ZAS6QDVoIBkSDgUmYqyZivA/C6Tq61eOjfsN5A
8kLZmHhyQz61j6d1Pnc/hbFTSYVWlrz679irb/QFZGUwCUeB2KQQ88skRtuaVNb6
mEfcW+6VzcQmoDWM93JjEMICJzIw8Ucife5yHErB5jdXjoqmLzhowEPwnXouiFWh
uGnrZnUN52F51p/pLodqNQ==
`protect END_PROTECTED
