`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FTwp5okM5FcBmA/BXHMk0luNt9G+CR4vX4sU0BYD/XIRa3sryCxNgI4COAf7OIz4
E+6194Cv3/XrlcZ0Ef2RYZeV5WNFbKJSLUNzWtSDQK8lZue2rFFYzSOqUcvlplfE
lJMqILUxXW5hU3T8eyVJm152xWoFJaMbkgBxEdFy4hvNx9/L4Hk73MZFQBgUxVwF
Vr6WDHAtM7s3hWRgMP/30CNlJtnwvjYlYlBVKdLNC5My9vCL1qYZYU1ikjYo6817
qRbpoX6MfqWCTwFWpDTI2t/AuYMB4ffczac61pGaVyoSN218J4dZ1T+fYRPjG+65
0BKaS1LE7dV84vuMSXvlXmiJ0KHrQn6nUfP9GujYOGArjJxGEREhKXoqKPn30wA+
Be2D8Yy1cHEwxzhYM08Zz+ISLOY1+QuvUU6gvHdKfBBjLT+IYTdvVlQwWoBsXgzu
`protect END_PROTECTED
