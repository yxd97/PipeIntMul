`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JkB2UgnCMGKgJQymenIAE8VEnU6sGkaydFYPeIwtAWEWRZp5oxOOSdq4jvfDKF/p
sgoAm1/yg9nhO96kJHTqVgKzUR9bhfQG0Wary1Uk5PFQyOe1S/elxegX6nvO1WVH
zOf6kK0BQDFA8wciGWi6eSrNuhokpJo9o0RpBg5/bNSJ9zgrYxmdNQ3wuDTt77+D
ZNSmFPAbPRLEJAh0Cu8Im5V9Xzb+yKvV8uFVO+qjXBzckdcSmM0p5OwC6KCYxOwt
+yMjmh0GYMZn6ptxN0829h/RPHRHikWazEUVwbR6kiBaEGkvZeQD1qXiQgFlcwBw
GDugJql8gRMibOjYY/tlCLl+zkOyOJH7LHBuTSMVgY5UOMV9sDMdpF6cwJaGt0WS
deYvJcApCeRBMO3ZCfPbcPuptCCjk15J2gr4eEXYaWI4AgzfngsXooDkkmSPgFv7
Rz8Mls7gkLJxAPpqOvAZruHB2GykayxMdPLjWhx8LYJnJRGXz2IC2V94oWBGQcer
gKdYeiMSR19rfjVp7jCyHB4Btq096QW2wrTdhGQgZrzcp3hzVf2dh91Ct3+gJgUe
blqzPEzAI6AK3/SpEmBxxCjuziPr17OrEa2Abb4OBELf5BLRu65sgJIIJw1f9c7e
46RryPhwTcUD1JC4YFY1j2hV9kbKFuHkR1jAixUd49OVcIpvPmiOlMatKYErWFEe
xJ3lJD8cSG08RgTId36d5xqgIO9AwWL837dxAgmx/COln5W5NPMjm/n7sErHJdtU
2SyR7czXiu9UGTU3DHOKTD9WbGLHKuL46OlRCig3/mQ=
`protect END_PROTECTED
