`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
udwjNJaFwYUkPOnDNJEuz5NtektlubmjJv9CCsYWqoISK20bDMa1tIPqGmyloBqr
3MrDUL0H8M39Tw1GgECVrqR1wSpaqcW4WHjWrCcUrHJnEurxUwkdKIDhskFjatOa
CnI/ltzOxYjMEsaEGtdipuCNMLk9v0n5tiYeUD4jWE6kbKLZE3D9NYSwceTOKsUd
BObcKhgHB7W+kpZWClZehFqdTgc/xGX0R6GGjmWTiRhOW/mtG6/JXdQg6raklOUA
EOHTOGv3vD7kAVmeugR2B38YuzIWzDhltFqWcClGPzoeQ5aGaZwp4+SdOwsVhRhW
aPWPJbMmuuwfXceUa/shNrV6PrQUUGZ7Qq/8FACJPawDwAX2onpSkg8HpSt/w+hc
zATY6AAIoiEJ/nRY7hoyeQyX4hs6ySZRBpiTLFKu1r/N8cC6i9zac7zlonyVFPem
hEWDFUkHydYYw8uBCYNzoF/iSDQqScFL78jI4aNU//ZebcVmdGknH/V5TJHcD2Au
625D6WvhstHC4+XOAYg5R2bAvQNEfkZ9OdbdIF4hWAnyq0HgDLdHofr2YEYtpqw+
/u5a9WsdV7CJdBMhCWoDOEEqjvOObRCmlq+7B60DJ7O1+fYUzgPnIJwkujwl8gVo
c3qW9TeR28RYgIQDxyTNZ6yKlCJ6i1OOfJ/i8cEOf4Fxf46bdVNIp/cbUe+pfSd2
uenk1Q3GbwCsvs5AC/9wWYeocyzbYtYHRsUJlyHLU0GuEIgFnaTWtW+8jaiVGSLE
`protect END_PROTECTED
