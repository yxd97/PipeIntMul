`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VY/D5latupoDR223Sp6lIR/t+zQKM7NutytBEifbq6LqrfiH8vkn6bLPdjnW+GDG
3JCOmycfyHqXm+bc8w/5nA5bxaK1oSzREf1D1ry5P7tJNNDTUQ2ghuJ4m2qvU1cD
IdywZxNDoBAAFpqaNr4PQ9xCtampXmSjjM0o/izOY4zj7aGoDO6RDq6NSUwzp3mK
0JZZhTGglksPGvecFhjwkmkgTAmvi/6rbF5CjZwLTntwKXSia3NH9OUygqhrr+Ta
lSRZFFjEo312DklWOSDC3LkLnuzm3XHZKmKNpN+gjZjIHgX98Piyinbf0S1/Wc7l
GcYXz4iT/VVmkeRJS2m6jGIr/MhNsE5nsFM9VLSQ7OX1L+i1EdUO2ugE6QknObSU
IMu7wW1heRUVEXpgEcZYs7B/N2zEAwzVS/D0OOytanS2hJXKyS4aQwSgiNpx2L9Y
u2LRdNR4mhKDZM4ySMnTYkwHD29skpYzFLScgV/lBH0neFWoxcfl7tKzZ9Po0xqX
Gw5iEpgGNkzc+8+BViHDzfzY+/wL0CQq3i66zq30s6wVCca6I8TniGQMqPv779cf
JkBIfoadkR1GRyzCID7bNO400yZ2xu5Q3zY57vK698QU4pSyq5FeI8a/fXgynCX7
0gLX5bA1mkYPa4rgHb+fFAqY7BX8JA9Rjz7mHarLL3c+DOTdDW/loggPtPEs6qYK
ZRhgAnKG4vk7sO2nLwqrRo4APbW04+EGymc4z/QXwipbz9hpRplFYjNICGp1uqz1
a5bBVM2wxNENa3qaM/GZUNiMAKIUy06cZP94XoB2AsZMG7BioPcVPW2CSREU+x6O
hsURIrTaujyrVcqqp3Lg+z/bR8b6YuPwFhEl+PL9xAoythI0ulo22+rL0xvtNcfx
ivYEMIkNbnOOznyP0+6XWd/DC3PP89IBxCmYFuHx8XjquCayKympSi9KUFVEQVmS
eYufjz9MZ+QNszv4EPtRyMLuVIBl51pewOm+XHROzECRUQN5toJKMLn70Rl3SfGW
ulXJKyg3soE403dPjgfLfrd/vkDSqjqu3aw/zOHT46Yd+ngA6bBIOKMUK+eDxqQc
LPJzYIUoZeQBw8qKq0EKOGdV/EXoadwVJyg5cCqnl/ETV2IuXIK2sySClKf5sJpX
pKcFzCWznz95Foonpn+pu0iaXfY0mqMbc8e2N6+fVdzhALHtrQ9xvdXe0eGpYaRi
gd/qTdrgbV7f+c+7DjoxSSU3bN200csiyCGkiOT5YER0habVszTqgq7c4wxzuzwX
`protect END_PROTECTED
