`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fApeKCZ2lMsJ6YvpS6Zd7bW4e+jrX4v1n6hag91C1rkwYA7c137GWMrnxcfWf1yW
its51d6YFM+q9KEdGpbO1DXQdSwFJIMSa48v0Fte3lprKOJyIxV6eNCWX+AKC0Ka
JmgNR/8pdtcvcA/9lSQt6ecPcaes0AO8HDlVwGF6uL1KmSrj1myAd83vakv3h/4u
Kbpn3g63AAnUU1xe4/hdO1h0GG/67WrOC9GKq6V/wJFxF0jqL8cz0GLAOjtsC1Qh
RyUT9PmZsgnHcy7Yudrk4KSApqwYpklnwx5TJmi0hQrloCh+wHu826O6qP/HFmLb
izSJUE87gKMRJ2m/1RYHpKai4Y+EY9R1H+SZ1NoQv9cd1itQUScESi0c12LHNLvz
cqYzk2126z0w3vCgcti5FGoXEODidUWjDGdbkI89FB5gDqXNXuRlD+yTUlgh/laV
LO69o12p1GOH8y/cFhKfCsDBtqlzWJSqGHPxkVf5058=
`protect END_PROTECTED
