`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VU8kI3+qTTJndtzzf9YnblvHhcJiQ827nSv1d+9+e44sBkKucR+GgGI1Ni23hwSJ
wXEIVp2KQ9gSD1NOST398tvc/j/t5c33DiaZYZkEQLCyRM9uXubFNx0lG0hFhtmn
kNkgOey+P/fdcZkp5jJWg5WVGNxk9zu8QlS84UYzkybFMOvUq83Y74YnDujESqLm
424WOis9VMcbg3JjjoSTUhOCXf2eRKN5lB1KYvuyRzwcSRd8MIkhl0EkokMi6mY2
L9Zpw/u66o+6ridZYrcVphYJcExcxHe/WcmRjRbOifBwkgtf4e/Eua0qm3N0nZO/
yIydpgilwOur5r6VU8af4V6E/8b9ORogaPeiy/yOrkyRJis1LPRbt1yHmMHn3liz
RyVSvxe3kPO+nfixYOf1l78zSHblVyQ2WxZuLyb2BFYCs4o+Xb3UBISxTtcb7d+S
nJmL5FKQGxYZjgf8HC5p3tERMu9FVA+IBIWMLZ7pQBKtvBEqfkrEUKmIIzLMg2Ix
lxi/W07sbs1An0Yn7RkAmMGYyqALkPsafY+qy7uABbl1OgKZyIsKNDkiw9tbafLT
0Qfaw4dxaFNY3/OhfCG1rBzo5/ru/w0u0KgLQbQGkEL7XnonDcD45I6bCGBQQnD0
oiMj8MplEtjX++ZqMFVXfKXtK8iNwpSf33VypN3oYhIOj4FDPap22+nyflG7IxOI
Wtm7twN02ImGMGn/uKSF/ZpqXniw1A2O8QzRG1ZTwYiI1rR4U2L42yXdJThKaD6G
ItS5h0Udntaj44l+kP7JJA==
`protect END_PROTECTED
