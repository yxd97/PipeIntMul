`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unrEMvCwtCUF3tcHrgBLDssQeyg9a8ZW7W25HspQxwzmE6yP7eDUJ91LZPf4pB4/
GATFIMaI8wxsEfuj2kxI8mM4N9bSDtXRD/DHe/pfoDPRIuMH40WiR9zQs0KzRIQ3
ajVtkWpp+5x04EsdJCZrf4iRpooUctfIG2KmjLbbSQPfO+1/guwYPGYKzePSaEhK
vP/4kmYnollbYpQ98TQeNUWp47glFqfXYNS7+OzzDNYvcKhF6JspAP3+FcjLlNf9
F/LftcMUH75w96JpQsjdqnxqxhTJgHKDudxyh8WK5OaDgjPsBK+yLFnOwJBDtvuu
fQaRY9zjOI+cQKpsEISAQC6MZ6kQvtAk3DSqnIW8/56NbfkcDTV1wvZ/WXv+senF
2GJjgSWvZpWPHmjehb7s3R/4aAi62JeFd7NaYtMS9y3QJaaum9HHR753l3K3xzpL
cAoLhoIHbogG8yWq4cqwENcDAVIA4thLL74F4a1cEkEwQA0HO+qv6w5rzfkv7ZMK
43SlIKosbGGFikXpm+5VeQ96ZQ8BAcBask1iOQxTXTa2hZan1llJqWshKWu0lolF
50HeuXUCGn/R0dQFlYV5TA==
`protect END_PROTECTED
