`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QCdIuJs2i366+Fob8hpou2rzagr2vtgo3nSR6eyYbQVMfJfix3y+77KxzsaDN4CK
KCytKjE/Tnw+xY03wL2HForwDT6t1aM1xuDCc/QcRL9yDwEiiW1JeZOdZw+DLgb4
2oMLc5ubmqRty9YjxEPc9R9hKJCvBeXxNzYPXEu6WZB+0gAfhdBT3rpplVr3h5HN
cClwUa3NjU9V5pASNAaGez11tOKXV6XwQcjFiDuVTFMY6ycrHRgcBFpPzhCBgBLQ
yNAZgmndevkMWLsHGm3EUGK5Rs5ZdpkNl6QTSpDmjBLu1+3Eub7Ox0rfFInqjXO4
gxrXiQdcp1mf2gx8weUU0jaRH42lo8PgE5V4LuPYccU9ntoTB9c1mlTy9OWM5NF3
1sxEB5I+mk3NapaXpCGJbfUX+rFRvjuBjwoH+DX1djZkYzbT8NYBjqfu1wkfpzCR
1o5afINLJq7cETf7kUn1KmKoQie/s+0bu9XR2JDr8pvy4ZbOFdpEm9jjadJHpevI
UYdeQHDj86qmgvYedddakS9+DmsR5u/5bNnOl6ljz4j687/GgBcIb3vp++GKo7/q
jBNpGJppAPdtjnEWcCIDUSX+DFr9yswimn83B0xyj2utKHrWkJQ7r5k+pxMgoNIf
D3xmb/BN8WbnQHNacjwVBxkxhxQnu5JOlK0uXLIjpXn0i6JTFg6GU0GK1U+aRlbs
gDLdFPKOJkiC76GLT9mUYtex8OAkL2CisRxUfq1siAAYwLRLsWBJYcfsDd4VfaAq
+CIB82G1Kr8E2P5hk9fCdhWsuV9cxDNA5khckKBYYIXyc2UXnKzxwIbdX1lAritF
BivF1djllk0KnG054SwCphU19eKoDOeDUl7XyPaf1WN/bJoz60Tub+Wbroin2P+k
HbqjelZrSFdYKv7LDIFlIe65XwKbb8u1q6FM0X0eTbtKtbrcgpi8PY7PQ0/iumS9
lgwcmXVr3L/xB4QxR9X9/Q==
`protect END_PROTECTED
