`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oFIAdTaaPcUzD4VyvDSbECEydTaJ8ovlxPWMA3HfOgSKhwGFivW9KdhiacL2Tx/m
uQ9gST7HW9Gd3cw7QdU4QUmi0qa8y8cRrHxraSU/KsPb2rZs9EvhY0KqNEX5dDDA
ODHK80SjBU2Og4y1t4Q2YdSEZZQ6o2OD2CSACZPQOfCCLjBJ8qpi+h/tcNwUew8L
9jLuoFslpTm4rTn15tERYVvLNhYRQnKBtJWymtqN+dfDJYeh7MfdnykUnC+t5gdh
eZDCZ2Dde88sNM7J1sjcdYL6HYGlCSmdzRfcNbyEdO0hzimM9CvTWgQWHxp8zaax
I7S8/AytuBMO7NC8MkJhESKnKHnrGO7QvhZvmRkY4qQN1Mm9BniscnJdjGsGLySL
C3nRvEaEDt9NtlCMi0Fu1XA9zXbhhC3qRB5UJ9zlEnn8eCY5HSHtcAnC8FMtWqa/
1tc9UVtnpio/16Np7Gh/0KiLYtSTsFQbGqCjfGcBsUOGD+62oxSFEBbFuZLgUat2
j6hVjTNq07dyd7eM+9I8UkTEiDxBODoegOsxy+LdxtAr9uhELH5BuceuyMShCpiE
`protect END_PROTECTED
