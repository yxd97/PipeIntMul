`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6g874GKPvmgncr5ZlZ8bfiXEpVzBAc2LAgehvWsZon7A1cfZf42taFeIxT6MfLn0
n+cYgkrrDGDcV3QrQmy3vzE7u9BbeLy5F0AKyD4zV1NEbOKXxZuqkpDVUwLVIaIv
oVnJJ9MLqRlVs+9OoRcZC6FA8jh6KbgDWeD+Z3SF9MbWMrnHt8aU0MUps7FW5xFV
DLiRhIJhCUAs2y8s3lkvV03OFGjKml7wU6BHpu80qd9Ux92bxVfssoFJVqj7osd5
1HAcEn8jMJaLRMzqpXdATuNHikQLLAbwYW6RneAhSYXLmU7dt/Bhhp/vyAcH18oo
`protect END_PROTECTED
