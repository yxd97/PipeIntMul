`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4GWrHvI8dkWgk7la2CRHHKchXauIsqvHk3ihHYpWiu/qO7XBcnQcHySeg9olZVoD
QSEJFf9LsSXAAKGHKFQwCbN08up1HTHNsOt6HssUySTeshAFa/JMQp1HvQF/6dXR
8SmoQIh6id+flNZn5IURU2tXLnAsrSWPhFJnN4cD28vT+ST0ZVTaXXSw8QZqe4zX
LC7mT6lV/PUbf+wA2F5mH53zFClkixSkh9bfsWW2zTO96aDFA/gKstRzCptyF3bV
Cc2DLRdN1HAiSeAAuGvYH+xglMmMFKY7JEEWyq5KjCX5bb/TCpfZeVFUKbtLPEDK
rHpTgLiwmKnpQjlVqvDqaY7PY9xsec8/xswUmDZVJ5O2jX6Z/TlVF2A36nNz/XRc
ax0SHedHHYgnrSO1678pEkX85GbEftM82ar/wsFXdBsB7MpN6fSsavWl2vEqJr48
jBHNaHcd0aDJGzd7SH0D2PagDzCqll1QHwhg9eOnrUQbFjVxalOQKCa2w9NCVd18
`protect END_PROTECTED
