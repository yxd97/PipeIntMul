`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EvTEauve16ydfxIedAy/k/6EUMMlecnp4mzpWFxbnPmgSddoPMEEMi0c0PlINzXV
z+m2I5eTNXwBTDU8sip0yreftKNctPufK9Jigco0F9IvnPf/LSGMtU17lQFGcbM3
ZSa5D2txuLOdQnjm2P9PUmtE23bnQBMlD2od8Nr+M/zC6GO5ITceNTTYFVoCc93t
gZWaCAixy2KpuNr099DS7TD8anQ7hIgQyaEa+p4javJY7o27lRBUFny0PPvpi4pO
jzr3jxfXI+bBmYjmrrg6Cik4OW+IzIVgMXF0AlGsG4MPpWp/15fBWklytJuMoFtK
/D060NhI5YkfQ8jYswpYoTW+CGwXtqQziplymRYzBRpC4egc+r/JGjD/wsOi8liA
2fR++5BEKTnoEJRQFHNjnW1LetTGqLfLeuqp6lNbQIAZewuyOVy6l7I9K8ARaP3k
mAnML+V3zruqzglq7t2+oyTZ3vGS9PWTg308GEqTO2h7pl25u++vNj2uLHDiRwy8
Z4pPLPEUToEyt+nIL2mBCt0LCZKxuGdT1oZTCkUGL3LYh2njvBYRjEKkFadbK+kG
jogFtKMiwyMSVeWIBAPF70bWKKTdZTehlRCb0hgIibqIfxcWhvC+ynQYRvxN0bu9
CIk0Xk3dPSPU+voDUw/aF4Fd6uFQPQtAM191bruXLU6pPbv/Wqdd/uUFBd8QRw+K
PD3giXHEKUcNX3x61c9De42UBPISEMtEXh7IexG4HyjD5vToacEj+nZi/MQlqesc
FoIPK0pBFfRnBnfLhJoaB2rlVnV7q4jDFyLYAWI7lRekP/5FXynUbsNjWKaExw+T
XFsIcdVhNFedp/H8aTDeUEh+qBVHX+d/KlrQ7nox1JlHCghROQ3czTcxnFqvERIb
EE+VnuSRkiNnpDJ+nEOY2f/ajFGPsVB2dpPfDMfrcK9YVKJSuW6XCHeE/cJjVGGw
SyKMbqMDTsCPiP64of3bMsoA3bMJVlTqgyAztoOj6Zz4ua4N/WnctdasKw5uxOat
lG1djEuZT9OihDjqSj4+D5y77odnKnlxWfcD0XQWCmpLWaWIA2yDzSYU/jYLLIAT
kESuS2mf6G8U9oaVvDmYZaeczOWbhOTqapgh8/4E1ekSLIArz5kgscvS8SUqZa0c
mAeqhkxv/+4hQLN8HHhOHXXRPvMlvyYz988KPLe0Gv4DTY/L3jZcC78w/DyYeztC
1jTN6GCLGBAYT2Sjqg8STmHN7X6ldNhQfPoTGmrl7VvN4tsuaahwGbvA/1Vi/6K7
Gjo0aFaR3sQeisjmbTK2e2ctJjpqj4D5qptpGARRy5VLlv8Fz8rI7Qs+wT3ouZ0X
KiFqpx6R3ckP0axcWNW3JoQuuhC/G9sVPvtN+/GHUT+2oKnI50YCRlc3VhshHfoZ
PzGby9xZF51wBT+e2r3ThGDoIDQ1H85Q0ZGsHAAhVKJmZIxVTxg3T/Nfom3r5cpi
rx3ZM05XKz3w9KBP15hgXGiRJRnkTPMe8rYICOsJBA2oNtfNjoVvwJutPpE54jfF
UL1G14lZw5oLQVEIMyQyX97DGjiqr7IyRszdbOkQeqX8Bw39tBXB4LbCe4eyMjmN
RVDeF0WYA+vWaF7v+F5x/RoNpWrUkpD3Ujmer/Jsuv899FaIZzwkMS1zNPQ2IT/q
oyqJIi1b23/CARa/L27FOO9rpp+wruzF88z7u2tDBWOMINt40fh912YxmjNLSee2
LDMQ0QrTgQhgq2QL/whJwNGStSDJw4ZOhmJyhTew/BmKr/VyFJi48LLM3yhSk8zj
8YacHGJovpAA2dwrdw+yolTllcwp8QpkunBZjZktvcffeQCQ5BLkEAt3c7D8lQof
/fO94gShIkzP84hqDJWTpONcOg50wBxdKudqLNBnfGrTkCSFzmMZa11XjmBYKdSF
pO4wiI5E1mnADIwainRIpq947TVTVX1y6UvbylZKt3Jjo8s6Ib/wVFjLMREPmnrx
YiWgGcstnx7wzh7Uq9GWnp7ZWvszCc2ZbWr1g15k5Mst9lUioXxzlX9WjYamQHfd
HGlLGwD+aiRwSyv1/Om64O19l3blPBUTnP2IbIRxCw8=
`protect END_PROTECTED
