`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZvXj6oROnIwhoHjNKnrmy3crHAyEgOK5ZHmFA5kXDZWGOInV61icHfi1zSIfj+2Y
AIJBAvfAGthnMcO2kwPNf5mDuzUw5yCwnvoeqRyuJHytm2wzGxmrQKfZS9LP8RMm
WYC/0YHT+muPVx6WWbCk49EyhLR0eBOAR3Czs+q/zdancfiBh34R9rjdptmOfV0C
yhkhUgoHJiFjwONfhy/Shlb/c/y6nVLfLYNx8QMgBXJkzjhHePIGCWEGSxuz/JEN
EeFtcikDzZmvzo+MAAHm8ss5QCOKQIE70PJMTUPznPVNh0SMvmG3QpGjH5WZhZVw
+QiEBiFpq7w6imjIPPnovFc8AOHbN+NDI75lMSGpZK1+Zv4IU1gtTBGym86S0pCR
JD53pqnbrQZexkvtQTzpoUE9dJVWpK49MAOFJEBedIFZsZh87gCsK6Qs4RzNAN/f
42xU3jaIsZoin6L9fs5AeY9Vn0INLxu76Ig3bQTgK6Zo5n/rdiF6Bxi4SMupTKC3
NgK3a3MJgT4XkNovVo69ScMGgykcfPOFZM+V83AksIcvmVp8PY+ci/A8LI+m2+Rl
s6N622Qzrs9pVxj/vjg7uDuAX8WPdL4rKch216SU+p4=
`protect END_PROTECTED
