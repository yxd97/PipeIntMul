`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p98TiLE0M2RPvehSJjLFztxATmFD7scj2REtOSJoFiAfqjyxn4FFy9OJ/wzqUJSY
PEvLNMayPoCZtx3V4FUuDBXrnEI5mo6GFTeFh0iwIsrcWIIsaZTfN3E3vZ/el+iw
+94d21mFEw+56Wb2AW7v1NplGIcDmKJOGvpZ9P6FxasAa1FX4zd9KQ//piRWo2o3
ncX5vQN7Matm53uShcm0gdCDnqDsyw80XRgJdLZYYAxcUOiaIcmHTVY4G3Z6D0ap
CnoVn/f0PjOc94cixZFxjO0M4EkY4aXK7CSAWVLNiJ554FVjDRB/J5xENl+gn/ZH
XpfO8DO0vpGlZrkOSXfSTS2XXRBIjGKVGcP5M5Tfn6pJ2+sHJhSVquOcADgMlANJ
wHUtYXC6W4LikTktbnUx3R4+UjZPClBt1erv8MRX2Ob34TSh46Ej+7AARS9eCW8D
krFn/YB/gEtQLzQIcVqSUz8XaQzRgaM8k9EZTHAwdS9LdX2GvidEmtiY2djpKDZ3
v2C86jcQjyblRc818CRWf47dFomozwUqZHvyeZTR+YKBum2HfycmLCw3ttlhiGaD
/5X/reRY59d03QyGzFejhgsEXGHH/sX64BieuqvMnpdGo3rKjLVFqEq5UkEXfyrt
LPzDb7632/agvxs+2XU2KrQ9UuM4jSgC7Az57ICkic+VyC/RwGEVALX1GJjdh1oN
5eQq2EC7Qg0qtBiWLCzVelDYeHz+hka1RG8zlrWpqLOJ/ij9iQW563GlMi92Eq3A
4LwqHWW8gx9SRn8ljiXLK6VpDNVMpH8LAe28Pp9cjalzRpl/+5tskFGscZnYrnVS
B3+MZBCee4pp9WuNcj2Yjoq2SoEpViSsYcMyqrxoqJv7zIj2z3jdH+eyhTfTzx8D
Wv01rQzoNbEQayWVfON81tZ0JZ0WsZzmegBA68ocxFYVIe23o0+XKFbMyaNShvqt
YD/+34JBHGgRfDxfjjnbRQNmVLf0z1dy45mXQsu9Y6mccZlmd4c5j9EElxTYKT0o
JmCCZjcoIWZ0v3I7bGKpKyyWLOP8LgNjRDLtj5uH7LF5W8oc6Ys9dFQKAJNE6i1W
rEkdLFMTsrQMBhSmB7sqwKgF0srG1K04nfbd76UzLECTED9P2hsbm0zda5hbVpCX
xLFT0GXMuMYyE5/Ovyt4xfJrGWyf64i9L7kZ32ms4eP5De9r2ppt84wR7bCj2SMi
Su8uTKAKD3tYa5xgVlcXMkXkblr1VMkVfqHLlV4I4ozmdiwJY+YOrq9P3mxUQ/iQ
KgSQkuarrRzonZSOSRpO9CUrrj6oW6FMrT1jD5MlQKEUw3MwNxjBuQ+1Dr69Md8L
hTVaYagZKPC1ozyk3p6pjuJtVwwgTB+MGu94yIPaPBgXPl8OZF8qpLV3b+8qWIKD
B1cgoNC2t7+gOu0nhWropY9XHG7Sv6hltzr5HhCzqSCN8jj4iaL8QOtcblFiRerz
BROTTeg5aDasE9q+YpADZTCdhZnpcXkD+yNfcwZ/T7ZyFcJdv0GgzaMrLqgRWFjc
E2MaUfcgWHc0qJjyBRnaXHslwvRLOfXz4yqNAmUCw1iAbGvkNZ5SuvGKnQy0phla
5b718hTBR3efliifCmtzCT2zuwnlly/tZyBDijYbXVKCpKhq0w8OkEieb9AmONOS
x34l5Z2rcXJhI4+sg1Z1xafKfHRWq8ftlvcdMM2VPPzX916yEVwF/PF64fUuS1Ao
`protect END_PROTECTED
