`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yEiTFYF9xjh76zP6U0fjW7bqlOiev3lXDZ/eZy5ErsFVhn7O51J5t7qYF/CltHSd
EQbDRpH8G43YPhzsnt+RF6uEbfNKcIbDnH37gwnT9viWj+A2iyv6GEcukCBSo2HL
84IGsBPKxhk3OUnbO10kfXrsEPZZ1evj23mm1fDcqZTzEPMXETs5TXCuDvtZhG22
z6eRbXD5R2wXrFfhpo5L6X0agvOvQaBU4YmSa6/GB5VcU32W6by1X1EYeYuGwKBB
U/AnI9U9RG1WxTSN8KjV751JPP6tYp0MCIv8MYr7TKdbAFldndwc3kRcUPFtZsTr
wtBmtjSxlME1ixR1I2Uu2JtTcxjoLKEoWVXFNYZkdYhgBPhgfvUNC26J4P2uBr6m
Ap9NunuAj5jHHsRLPu/8EZWRDnGjBJoxzzyGp1MncMw0d1n0vqGMrIWjeEt0OCp9
zQM6EeIpDpccSw0T4owMH3jYHH9GEYLDZzOkF8FqPsceOfb+vjO9V8hP/b0nG5M0
JCroabOYXhONhTkibf8NfeRYdJa0nVn29LkB7GEsYlzFMOTuSAibASEL+HtcEG5y
TevbVOV3bw1qJcX6jcAwHVULjCme3p3xkIOz6mSuZ+od/xI5mpOjBE1c0SAVjJ7t
K7Cq9ipcddEOh2pJTOBVTAI3ZnBXvrFF0NQS1WAOvCl5oUeCCzX8VPbMRbWpeUOb
PWBpeRPHDhIidWSVPtBREqyslWA7TQJSwYbgymv6i5BU1ZRVc7rOKsqE5fT/+JNz
`protect END_PROTECTED
