`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fI4u18HlTggyu3NhCMsdqUDO6CGyZmzXRkXXUVvLSjfh7P4HfH++96sjWKnAkDmA
FTVW4YHIa4Ixu5W3oH9ehOt/uqAefsCxnfgi3or6U0jRvz3Vo4xN3IcI5WF4GhVZ
JMT7l9w88NHxQCrbUdpt8251ZsZvVpQBW4ljpyMLUaEIyJut/71ckpJoOXAFDjNL
Nj2fkYK9USAVzoD2kDU0PoAa38zmqChRDu6iL+gXm3PXEzJX/6JT8rqx4r/ObFoM
eM2i2MDWXn0svGpk4gJacrfYTygmjuoJpMmT5giZ6Sv2VvTJd79XmJo25XNNmb5H
HkKpKA1Miyp96/Xw4/KS1K3x6ZKNRMwdy+i5LeYauEYJ8MR7/tVWEslcJeHW67OK
sOtak2ZV4tM18UhuEMlEnnAwxT2Q8l9rcp2AFNSUx9cFAmTINoTZUeTmvCQbJSbH
rtL10LjzEVU0e2c8sfr76KO/sv4PbTZZ2RN/omEKDaV2MYB0N7RC8/bJFO8R0u5V
Sxv2CrXm8r2VSGF4E0vBpng7DEfOUyBa1ckq2qVrtYPPpfvKMFfMAwzCaqlc4D45
qPVwxCnWHk3LG5ZcptGlFDVIPRlCNqJz1UjzpkK7v59fdczx4Rq+q1jAhR0WIU7y
oEBOpCzsYHm5t30FxtFD3dXjYL1zyAtUchvY9fnezbPBhnRP9fmDSCWnzxHCwShX
FwPVzsFN/kp1/Yo5Wj7sLn7ikuKmpXho4+OBk0pJPiDNc5za6Y2eXlQq86fhALh2
2LTkTNuvznz3mAw9zIIoKIH39FbobTVfTsg/j2r9g6k/0PR9h0llkPsBE01gN2PW
9cg/oWlDJvu1h8K1pTKEij3pd4o2rYNzOS7YAvA3z4lgiiIMCzQU0u6xvRVTeIrn
0QuKB1E+sFepN+NZlkMOIXZscDa4W7fIsayioiITBg8Rb+2EeomrwiYLAHWnkEdK
RCGwacu5qsvhl2T7SszugQ==
`protect END_PROTECTED
