`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nfucz2vCzCJtYGbDoczzcgYIPp+uWGzqvWFeqjlMYhITQGdJEBwR5KNFCxfffuCn
ClR2P9wEGQNxzqyBKdYOawgA+kGqJoGQD2nXYxP6K9BPPOjFCmQol9WnNky+WIxw
nHf8V9JHimZjBWHwy1MpCOh4vAdoWQJ1T4LhGOI7i+C8TD4vgdmsd2HCOk5UgZuE
mIRKYwgj/69TYqpNJ8tqUQygFjI0t1C2Y5+weuxTLVEk4sGCF5q34+GsYU55oMUv
F3zg9JXF6IsmQRrzcKqaRc9paUqCm1mtRsaK31f6JytMe486X+bzPBU1GCFDVus0
rBOp0i6TTy6MNYookN80XM1q7mSFLjx07T6jwsJRnD4nocQTcJewZv2F/IQQdekx
+qrvqOV7dyWMqJWWDKFIc6AYV++RcX/a8lNh59QR57UVobBDhrsiitj96cwKvsmJ
8k9ELcGLznHdSUIdYMLVSIRuQpOrNL3MbVeBh2DMYMF+Pbcb+CLo0pR9GyWWEVif
7zque3z4A0uM6HtswWwWy72K+2GaS0bSbeQb3WvPS6GEGIq2kZ9C84KQ5BUiBrr1
8jKMtcrd7lNp8At1P+DbYUVDHHeoxcOAFFd/yjZ9nnrpwahXMMP6kfcdQy4Z4oPL
XJyDxvbqVFtKc6sQ9ye8mqWxutkT4UiHbDDRq6QCvKjZp16Qk2HTEEMGVYjFi0R9
+fY7d7yA4XxQHv5WPXnwozB89vOhpZNCgyCET1uS0cct3DFMo4BuZ520ooyhJLTw
NKerS+AcJfk894tXQMG65Q==
`protect END_PROTECTED
