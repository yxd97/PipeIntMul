`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PTTZNbWj8gBCPNAooH6NN4S5n0Sd5Vrq7PJeZQns7/4I167jIvXVUCZwzsH7szBZ
tU+MXfdd7yA73rBNg/oiOFthyTXWG0Y4Vb8RciIiEl1PkX9D7xzBXTojloZJDZzZ
IreoaL4g7+CViUNKfsp0laBizvyUgIYQqOq6HJ8KXzAzcH8gWyii0jBVF1oGqCMa
l/+i5IBOuLqhpOsiulacfSC5a9OvAScnIn8EFJcSetOHj23bfk2EUmk5V9PjLK2D
zgvb86i+dHzprUDGjaZEwjsTAIbH8YHer4CCff6ntB01QCNno+3xXtXBU/+Ra3UB
PX9Bi/iR6/k7yYHn8QE+lgj7PX1yyy7Hb5VXE8vusuPY6Z2u+f2/e2P2flwDFExO
kB2cXjGKJcXTgFdCkojXQO4/D/4tVzYyopYdTglFKbOSZ03A/LCTqteAXYQ0VSlp
2vR/2bQUb9JaYcxgm/Ryv4/EEPP4Wav+9vWjexhgijA2+U7FyDoTRkKVWZ2ga1y2
Zo1Yd25O4yqsVASyyQL0Ll18KBClt/5yTRWATaTsmiYHJYF/zdgST64DAYNpZwla
Ri7kAbXqfZmq5KDODtPqdrOZbwj09MxAT+GOOcs6makzk8HyRhu/5umbSPE6AAmW
x+Yyqy0LXMMd8UiIMdt5iw==
`protect END_PROTECTED
