`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L59Mx3ie6TyENOzm/QBqeXfNkMVu0ff2RDTdZot1lZJ0s088qu5hXEGzk8UIEB7I
f9gY3PzoicyoiCg649ImaD1L0r37Q+NZPHlx6iq3flK7z0u1xdu9xYUI23GYApr6
pnVb55Dycd0QUMLqVHnWFjfBHVRztJzTp1V8fXtgCQPykQVe5o07jrZvKwa2Dbk4
kwnkp1QxB6wszT18XkUbU7r3tr/3BFyYU9hxdWgpew3fUPy2oLXHKjIYDUZaYUVp
8Enm19SVb94akhaEr6d+B4ghyGhHnZQv9VmY6Hz/ZtUiR5FRWLgkTgtpTrVRdrLh
XL1ZSJro52D8qu9zwbjwtA==
`protect END_PROTECTED
