`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5j6AWQGASKipum4tlMK1UsYtouaSCsdssiIadgpkv6tCfC1I8d2/p0EuwW8/rHbj
mhpo6VFRUvIVoek7md6pLkQ/GuWo0Q6cbKdJ9lx373lBHeXeG+zqborXijxWGvWm
5aJGJbbO0H+LgVOgnvJDXXVJ8WNBhMbtNqud0WgRpSDS/lt2siWzKu2YKUsDnr2j
8Ko53VM0mNxuO4Ie9dpzNxWTmp6sSWX4JgXLUmo+iKOZ3dQUdlMMLkxhVVSAqgCJ
Ir22kzSPkGeSyioSWlcB4jJdiow9DbrlfYVYGy6q1DktlpP77aCViT0azGEtgd9P
1WC1nRe3wF2Fhfwt2REe3lMW2BEWWVsz0XFxiV704ZmFu9sIkSTYrQ3lG8uWXkA0
CbmMz/lefZwGpmy2Zk0oAKDz2A3Jha9Ns6GjfvWq7hU8WCCYtW2evU95yElclyvi
VjR7aqYbkfSjwX8OfYuSy8J7cRmTSUchNSDngE7+A9WobHgMQclk293crXi2im+o
FTDL9iKct1mfVyt0ALyv0qIu8M9q+GqwXWc4rNv3KceqWFaoR+MpLBzU8nVtR7RS
jOTYdF3Rjcq8RIAJ8oPo2hSaZGAq+hBNvyzpzF8bK+zQ9SvQkLYGuxDlFyds+jkQ
5nIqobMTd84jv/xUtUqrrw==
`protect END_PROTECTED
