`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OOfOMFgisv9ijZhz8QdYq1lbI9+INvdfVc76esibpy5EYFXnw3TqkmejSlWlNe0c
YdR9U8Hc8t8plSWrrIHAHHFA6milKEWdlBacq1qFeApj7bfWnRDUuL0ovzxupfgz
+11Jg7jtn1AEu1w/87EmYUlpYZ7ifZJwQb07bCVv+cDCDN7dtaiLcBjCxIMiEcvG
CLqwLpqiYSF3AvhvxRqDIJaBWJWkNgKc7z9KOiNv4jY92sWu3ooqqYxtPgOesmr0
Y1fwAPpXwzEJYgvORHT7F7TNjQ/S/Pf25oEF9ICTDutnlposwLaQ0CCM6J2VTjXE
2h8lKWC+YpJFR5g8JXDSSj3RGvs13vlMPljdM7A95JuH1EuUk5C9HXePLHYwX2gD
imjAm1tmHgYbXoud697wpk2lEXwnih88u9LTnn8uaR2pZa246pttXYWq/0b23Dhu
MNuc1E3M0UK+BOipP9CmBlvvTN+GgFI7tlrAYhZnLhUo2gz9KQaKTiT6sMVZ0l10
nEshvKmJoNKUAx2DFwW5QMNEPzwcJVechcFA18EFW8Y3sL9DuQZwIf+bHiWf4EWz
lZhcr8hR3Njgc7SYLoK38bxGLHKHZoaYKQBdtIqM6a4URoGb3MfYhEmpJDTMoHQh
WDoFMradsUXpCtjyHYoMxun1dRvUPupddxu8EzMSeRy6yyjIJOLuJUhXWa+SBb7E
LOU4vUQsXwgLhSYMEIH7Gw1k30mnrSPLqSyJafdLXHg1ueq2DOuPBbZUGcbL99UR
ZkItNIWD1vPvkl7mE2N3LUQUeWzqYmzrsW16zMM6h6k=
`protect END_PROTECTED
