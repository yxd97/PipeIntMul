`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EAVOngz2ZX4ESr5Sqyli0qbHx6IfbMrgks7eYuU67Q9od/Y0/EnGMH7oYJGDjcSK
YtrBrn77Jdwg3R1DRVLat1ViuegsLPCqAe/6YyKQFGbAaSdQtjxzOSL2lp2DGyOe
x8Jk67K1TVqgzNWOQnOMLmWgoQZ8Wtfy+4a3pq31m18p4rJwsYcS18lBvydzr/1e
vPpFP6zbFoBcUJnaEQzbIK2Dsp1HM8vFB0wfh0kPvv51+Jf7sbrw9PzLonmTFOVH
m4bM6pLS13A9YMc20Hsh6LKjZ43NDD/Nsu3v83fAC1lStx8mb7W7LuO/Wl4fF1xW
NqJQbzUbuN52sgaC5y90IIqBYa6Fohf4fwcOxn447PcdNnsDv5RMDnkOGUvhtucx
NOnoYH1myG+MPKCIo2E58cfQmesjRs0QP6LBN+aaMJe3O2RD6+tZWw2gVj5AIzpD
LL71NLgE0aG5LhBqZh0EkOoFFiC/FgJZadduWFpFCoAghBGHf/SkivRsmyzYlv7U
Ymd63oxkD2uuMijFx/MBl7b4UhI5LqF0WGVVtnIlld3LTIp7YwHy1fiVFWCFD1hI
7Rp4dlC7UIvHHuZiPbqckbBXdrT0OMLru+1HDU3TodUfvgamfGgpSKCO0aCDtBBw
2SjZ8UXmAgIeUEygjly/HcT/WnG5GdOz+wjZroc7OzSgqlP34jPsyGaUh4D3WDR2
jELaXQhkwp+6VuFokJ8KSmCI7iFld06yxPWln4u9pi1zIDofkLVAEOn+wUS3GZRS
AZwuPn9pFyaGz8On6OQtvzQBghKqVbpYnGsa+KWLWL9+vEhsgVseT+X5ddWOTeOy
owxOuMYBVMplULJO3cWHGdVyZ0Cj9LIdwISEjHQDuxiySNzShQN/m+ls1UOorCqL
JVDoTxF+4Bj2WRItAfFWJ+RTw+oaCDl1DIzhrIOzCpfAEz8gZdqIgzfPM+weq21Z
CE+LZEq1gEvAS8nm7JstV/wMO9QKr9GY/kE/oaPstIGs+bbIj4tJN1DGn/auGWcZ
X7QeehIyqcbWCUksc13Dt/pBFx0BE58ejuLNn+NRAXtWDUZGrkwq0znMCvnVmKM9
4Q8LY890K/htBL1BvZ7BLMzeAKrK9A/Mmm4f6OAmynP8NOMUwZb7VmmNGH7cai1M
2aBac/VgHdJjUjxPf/FOYTV3OyVfnJNqkR6xRPZGGioeY4Nx6CyuzZDsk5XDnpQv
rkchLHvCrZ7qPdCrS1NXQ5pkrTVcB7BAPwzJQKy88pni4htew0gq36dpR359uNrt
zMOhR+/epWFWc+tyJdWUmWTZVCR8aG0GGbxdv/GC/e4CzugCCUd/Dk3wnBk9Okay
/IAgenlIArK9cYgWSMLPwEh6cjDxVbOOPwSqzXNIIl8+PoayZEkqptnKf1t6lPTL
KAyQ8k46jTi/bP/EGqUAvUs1FSvbsBEnZxM8y47dBC/YkmsFPlolZDvDBmcYeIr6
bCFIR0vfgGyS/SNR9mvUggkoHx6lSoDn+oXCkogP/ATA64Ghv4+pfRSyGrFE9Top
JTt95G3YyLYwH393qkwtjPFUS8erZNJk7s9dgaxB/bQbjTYU72xU/1Inp3mLxwom
OwMMZb/PAJ/FNdfz/pRPPn5eh4o2Kiv6S8r0UeqKVYqH+1ZmlEfh2zYDLZWFDqly
pNUXTogqSRXiniHN6zIS9ULD9MVOs6Q9QbNayvXSwChhRhiKXv2muu0V5LcDi7CJ
xQWzo++rkc8c3k7O1dIGjvvNPn2ObMB4Bjo0pe9ACAt/5cMQVKC/UfyXV1aRm7H+
MX+gcDwGeL5tC+IXTvw2REVbnLR8UwdzQdOTr7sFNBjS8690Gup2HtPzClz8Y+k8
sIHKAxJjQJAy9zbRdsnX6q0shIJFCXzotpyOoRHUlAQ4WvdjoRAoRG4r5TGxnP19
0JcydqNLHLjkI3qIH2KCzVQc88KZEWrloisjpTKSHrd5hvYFv63F5O7urqeLb6XU
1jEf0EI/Uixi2zo9zchK2W5wXIxJBWsgAI/LDsfWL/YDk/FWyz8K42LzqK6UrP8O
OchTSMO72g9rrWfgVTU8ZhKYuOAwWt+gPMjJX3+sAuTmqkfT1uFnBaTl2NzLFEdZ
Baq8EiDPScaWIJefImrHexsLvrhbgvx5KDCX0a1bhCH93K2F8CKm2VKyJTJZymdz
ClTb8KED5tTSoGaO6NRBjOTvuxjkqX1FUIfaxb66zr6oKbKqv8O+boZBBXDLbklq
T55KMqdGPU84pNY78lv0Px+lnk9in1DcJDS6O2HQnmQUI7VFFYnmStWOzyez22H8
vXW5qf8Qbl62OSc4gXnr3AthJlKIZZCvbMD9wbv8GvUoVDifPQbz9TIyMypP7Glo
HNIme3ErAX5T+gk13pI3WRPLgz1fUBQmKYGHy9hyTObjFGXOgA6sEqSGz/rs1V8Z
xGf7FckjA/QtebwKhB9MUskdy/ACyYV2CEAlZ3/Lpwgm17n+RUENOys30lXA3v9g
MWDCwCVi1CNIhlkQoHcPCL4rXtfmz59JnciIoHmp8DMyOrHjB4OwAQGR8JFzfmeC
fCsMVVvbFpqkDX36Uewdr4koVkxm8ZzhmFMffF04RNDQ6V4qpxUJK+FHkE7TdMaY
gBDq6lwsLbPpMPXIC+9Nzksw2aefsCIF4UwGnjtFt05PQVoR7KCmma5YE2mUzVew
jltlLuBKAxEgW75Td/iz/ydU8XFyviP3HKBtbAIT5VhJXgWdVRwEZpjOfV7Ljpze
bgCLUrhgHn4XRu/V+ccEwqNf3PBqoKKa/0UbGO703NDMuTpObxJI2wPRLxuZU3QW
erRtCtaNvf0+3IZ+lA0SeV0TzokFxlF3JSgazHN50Lk+It7KzxmsBAB7gztH33IL
xMHudD9iubZNlSLwMhgGPirSRgrFIEsnLCBTwt946RmDB2z9KE/7I+Uu+P0CiSoJ
iTk6ZQgYtbz4GFlECKG1pKV2x49jvK/y/wg5QQM601jfQEHePr0Z49KY8YwVze9i
XVzoNLmVlSbBixi43upvvE6pgJGDLgtl/crr+3XhIr/7pBLsrZ8R50t33RIB22l9
tDbJTQPM8s2ql8IrJ2gdURW9aE348I08dCwkGO0xMK9MbfPqo+LWonb4+v1O5Hgd
tO4EfyIZRLtgIzZgEOe2xxy8IJnC/ogtePflKaUURSzjsfNu3ySNdWCp2Al5oY4d
MWM5QjMtXItk0oad2lr79tfD0bmiOwMceG3B2l0rEJaYUTPnrZmTAt9oxc9Ozmxm
`protect END_PROTECTED
