`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/bhMFOtdv3e8Y+f474drGXbdJr4dc1vgPpy7ibNAocv4HpIcuPa/Gd2OzyjK9sQS
bgOIm0lUDO4QsJWHFcbB/cPXXttmQkCReiWIACASUeswU9EGGPhn47LG8uPnst+T
eCFxJfeJLb5xmoRKq3jLiygM8xgGmLdlKMvzu/A7Fcx58JxUvuoHeC3ulkSOed/X
lyodEVlKY/yqosW99b+HtxJDGSYix+Xmzt2Mn5NnhJpF+MECrGVyBIuJ06AVcRrk
pqWCV9Hz5RjBVGrau2951QDAF35ngHcMB+IJ43RR8dI9ZbxGeqeOLDF59xX+6d+q
bIm9ydLkSooIpStCG9O4bt+n0MTgNhNT0fCJQOKiItoU6VQ0owNMloGsu357KJyH
hWmHUYY8sBWdTiOCFUswT7Cf0m/GTUrXccazQSw60rw=
`protect END_PROTECTED
