`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
224PAfyjrovvRKHZERFD0A/mtxbZC38D1HL9aqpE3WnWQgwJcp1c1jD5QIg+wp0N
TVwh8uML9HmwIMFhbvswtZys+7kh3PwZIvPv9o6sLYXaXQ+AgaTKiL5mbqub/Q9A
97AcERNNilKNVtxNSh8mH8kU4DDkhHaCj4kLBhARLgKufFhDo+QSB9UOiZF0KrGi
BRb0xaJF8SlJrp8Oloy+KJUwkaihlKmKSR/GFsygmHrwDPtG2Sor7/Zg1g6Pk6me
eDIDOSNjXLs4dn2GbQupxz5p6/tG/vJH7BkUXeFke8zT8K40nfGuwAkNxnYbINeD
yVBAeaGVdAGUDU4aWbJPg61UVhasUgu8Tjn5bzWHBiOSZ2z0isR0UKZZajICiBuG
TtTmACC+UMDD1lS2hs5hWySwNv1g9OYRXfbtEXXShkcXD8wI1KTqjaEnUzEWNpEm
M1nu9V5yW6zPquKR+JsJ3w==
`protect END_PROTECTED
