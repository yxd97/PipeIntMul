`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VVfpI4/+No/f4lfVCudqkorMw7hqKojCTVqWF51tOshoNjOh3A/kHjQ/o6CFkEp4
v95ULcuf/LzoNgDL/1EL8YHnfDvl8amv5lePp6hOKamCslcHqOb8/CsEEaOG4dYS
IE5RzI/VsYLSCoXn2RWzX5WUCwZnqtaYNp+JZ7SjhXr5ShdLj79HCjzhmuHzFTDS
4lnCIRZ/ZJPaIjjimj9MhXYrzy87pJSwRdxQVg+LqAm1bxAL2C07+CgLsDpBO+pQ
4eJGR4QHnh4J4HkKywghI5DvWhmeOVqjJgynS/P47RvkMHR5a7KIlsPMSfgfgyKT
q8iYXxINgEBsHcSEL3QB1Ymqsdh6unPdi1EIFrD3x/lrwk3wKoJVfA6KXOIzGvko
xjFoEpnzP+OzWHHzcqTRRV2gLmes8Px4h1I7a3lSSz2sjer8Qr5UJC9dG60s9yLs
Rl4LAaep6My3iS7CAlA33rMK/8XsTgkV6tsYZgbYa48=
`protect END_PROTECTED
