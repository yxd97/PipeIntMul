`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ujc6OIR6SkUGL1dqb7Gp3OAPyHGXID99IxMBl+J7vKlYe3AsgirLfh2+9bI5fA2Z
O2aNezdVeyx+JapIOjkx6g2YYgFJrdFAl2VKqQLiC/VLOK9f0c8ViADf49rgE+qq
+0fGXSzpgCeBwT7z98Sl2B+a2SKq7w+7qwDL61J64rBhztjigRwvrdG+whXvpCjw
obM6LMOfLrj6B1o+/Y66r/B+l5re9r6lAnlEJAFc0sBJYbJlaXMRPFviLNGxWjFh
mFprMeSB1lILquUT4tDp5fvcAPTk+I31SrbxHbd0Puq7mNjo4iCMcjZGDClDw72Z
Z75+dRxnOooRb0F50ft6Zy7KQaAWDUnLRLFZ0A1Pvjx06CKAh5TdJEWptvm2j38h
ffVDMCOHedsmiqTZxjXQ6OuP6W5uo8qfTDTPbOQPT1qgtJS7xEom0MGaPlEYo7hd
bnyj3VMMQdoRJSLcLN1bBxnQBvDodhOLUEtZmJkb6k3CGxWddGT0E4xTA4uSxMyr
qfw3OOxFz70Uoidq+omMy3BgjwEzH+STHunVAFjFvn3QFzJXsb9PWWMgXzCZTLd8
uLJD8bULGh6yRv8SiUDGxb4UvU+NW+AMUnVj0lxbk2kodB5w5SF8YQUQEudrO1J7
501ikIsutVPxqNVsjWsh2vsPjdfapM8UapvhZp/ZOJlRzuwVLlpU641lXU33UK6Y
I1j0bW51QfKEf//SMG77zvlKQ9us1mdDJlwsJD19T8Y+1B2NsPLa7P9KSfU3Kz+Z
gG/yd4ZZWeP2VU4XGKivcAH89rhAmb6yvaIQbzt1n29EYaBrN3SIqOOCvKUHncDi
EM+/xJNCzw9kEXuYSdaoe942I8Aavfvxb6nga868ZgHTGM1w8CY+mWUpo2NZZxyV
Jhr39TPLw+0aXLRWcx9EdxlE4tWjHv5KbeE17+JFW71sMyihwDoHDBljhlingatx
PsLe2TdPJEnmSSM4OagRjA==
`protect END_PROTECTED
