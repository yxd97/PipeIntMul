`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hd9W3Cd44Sngq3nhTGssms/5X9629WPuSmr0d54SmjHHNYg/CALF+wN7cVf/oERM
Bv5YaO4Foo7iRUYuWerKQhsUYRv5MZmqH4LVBngsDsMrkVU991nnRBlxNDx4ESST
Yp9YB4TTzanFOV3cEBhM+aelc/QHw3hJEQElTcGPMH0p+U7XiGHBoukJ7BwBs3yK
DA77Hh/HlfxbEF1iD0Oox99+4O+vHuexOwrOcWtwMPB5H6EPO0yw03IqijTTPDwS
FRA4YabcObFsCswATdCHa4BIoiVemDPw/f+sPOWfAdcC1eNz0Vw2Rq6U7CAiuv0L
HWA9Sx5pmlC676kdrnLDug==
`protect END_PROTECTED
