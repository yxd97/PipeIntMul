`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ynka4WFWMEhYnB7HJR5qHD7Xl5iTiuBNSA5b0mMDLkm1iUcm1gJK3Rv+Gta93zDh
layv0TytEHCUJ+fn0ju3ThvfTbkWdkNU2ofKymQKdX2cB24qjAHC+fapVGI6/iVU
dP+/uFcNBLNQJsx9GVx3rpyVUPuw+SfFNn/BNLU+GKVzOJVLlla7/tSAK8bPKLra
w/xJlP9mZwVgapGwbrELOGM1wiuH8Y1g4e2sOB69kqnsWEV1jNy7guA+VXlF67Ik
EpyrYqYpzK6Yq3xLPRayrX1oylaXQD+Sb0u2Y5IKInnzD2eEkHiAkmhib8Gxo4jP
TxMgKgK9eS03xs/F3na6/f1Aj0B5XtCYvnLXcaSxe8WW/P55Miz4+L4n9f37DmZ8
fFo8MP51VlTMeT0Gp8B8PA==
`protect END_PROTECTED
