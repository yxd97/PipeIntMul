`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WSz5cAoKqVClghllJM3r37iQC9N1KPhgUMrisSA/er/hbsUxwNAVhHd0Moatf914
EPvh8+lnK54iTAZhln0hfJK8sK9/xhRukYoRMifDLLop1cqGJcQWbpy1iFKVrHLW
JDdaPRjQjm3UOi+08u34q9wN/QMFF4hfksCUtUykNoc8pmIpDeCfp9onxIXHqMia
2K0gqhErj7Sn/rdwxgYGk0WdBFsXzjdeBUTyYdhph4Nje2dMb7Y32vWO2BU1Z35z
gY3SINaTyNbRyUnWpi+CE1AT2tWNtKD1B3gqAA2n0+azulL1SqWMAJV4i3H9JAYB
e71RDJePPRldjwqdh5NtrFdbQgwc4o+NA5a+CwEi4Ne1OoPrMstO+y+dzGaucvEX
wRZaBmA6Mre2eKX2YzHejdAS1Ay+vK8QZUr5p+F/ZzJPbs0curPJNEFi7YtNFZb5
`protect END_PROTECTED
