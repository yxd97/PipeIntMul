`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vLPjHXgSoqVLVXcONdMUZZv6FMxc2UxHoXeCpySKPi1UvbALloJdb5DUZMvdLKHE
9uMWxeizZ6lCXm8AypQZ3u3sO0NzKdulgpvT9eIPtGxsjPctP1YWzXDgiFcftgzE
iekYsA2t0HQZnXC3E6rRGOMugeKHl997H7DdBosLQP55LdPndn/1uAx72JkDwm9G
n1MoqJ5IWrVit5Tb01Cw2TapGnEcynqSSjPERjZ8r+eCj1lL1j6AXX9axFsclg4a
xiw7/XfoqvlG6V8HdW2SmUfX0vSR9zzZMfhaEsjRDEvw/Y0JJqG8/4eLPSZk/utC
Ndeb8DaaswBV2Gb9TXpiTcyTMpCZPbM6PJv5lYpxRQ/8jGnzo59JCXcP0xHPJ401
7k9mtdD9tGEhetIJGjw0rYIWxmkV+wJ3OZVXblyP44Q9NXWq9ITxs1ixkKKf5Az7
SrOByMSnN2vJD7Vit7jUtFDQ62i2c3ZQwUVgnk2y5hk=
`protect END_PROTECTED
