`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiyYymAjD777xN1B0OnLbGSqzaus5RqWWCETLaBPxndLLs7BIMlhz0TRXDHT/msc
/q3zH0z/OKjsCnwOVpjxmgtnxFc1stxt1Tp7L1h1bwWVj8IhnMIisQ+HlfXEUVrn
vug5uw33QSV49CzFPj/z5yBXH765akjov0v7cyQpa7fe/WbgSB5zF1GCBbliGCnm
dNq7CI7Ehr55oqAnJPxzQ1WOIzIUycjh/0FKge2oqUlB7DhZKooKnYuV7r0Q85v6
lI32R2pGUHlYsFjHx1Zu4IVy02kMCxA/7imF6/njVgSYHwAvGC5uw1b+6lbfLk+b
/X2G+5V0wvI00WJliECukai3eJlWjqpEm72U6nYnglNEdlat/gckVpo4Jc5VI/E+
7wJWTV1Vn4uTJcNecU27EmAGvnx/gKRC9gTyKcWFUfu+/NuVBqA2zC7aEZEi/Joq
AxbJM//LCbJ5wcCXvNZF2G/juX4ffKA2kYrAjgUuz/tDZJ3+BGTVqEgksn/wlVQW
1MpgQlUf0nSTYt0CzHbL4RWFVp6Ogjwl5sorZTCMrd7sfe9QHSrVqBsUITHNy7VA
fKRk82i+Mm8w2TboXG6ayfWvlRp44Ssa7mVPLPy0MXKJ2x7igRnD2yu7DQ5sjY2J
RRYTAgjEmsbUmQRH9YqRLHQsCy1dY2VWpiTjy6ieDi1Iiw525/De+0Sx72fDHcH2
uymLsImXEZrA6Qm6vP7hKxxwgburxaqh7GQ94pDmcmi3irSu5Os/rNncyEVXpuWT
RrAm3GhidIRRt1lDq/QcCgA8GwrXy2SmUg0t8ATeJOr0uMoDGoZ6v1tW9bxzXZIa
xH1NatxonB4FIxwV/bCL1MGEwviP6+hcJ/mqN+7QQH2xE1RIkBDDD0pxB+TdvAle
8DHL9h+KXEA1APkxTxeaTjLBWZ/33hlGKKjN/H/gTWmb6qBsLJnhQoX23XloAUT+
804UO9MXjroYrh3Dzewl9nSr8vsrvgqJo9F5L9KpW+sOjVE4KgdiVTyZW/Re5nJA
2ah1vcy34Qx5qAiuUJBPWSWAOw7IN4A+qSvd6Kyz9vf6cBekOmzNI+w61o2aDiqo
AeD87q+OXjwu6YVewmLf7zIo1siuCZ2l6UJRS1lArXmK0NaNqfqwNwGTDqDI0f3F
hPJtmQDoq4ni0d6FkLURWzRrkW7IHOLE+SCYcNtluZ40deEUvTAm+Mkp1a1cx2N2
Z+xtymyaGhDFSv9VwAvmHpAJJ5cJIlJhrZdF3Z4y/907oX8Wv20t0IS3UZhIXw09
rz8P3G0pmmlmtTiVRnyQHyDlJ7OK7akdDiLnfeEggSSrXxr829H1Hq9bvZ7lePjV
1kTHEmydQYWjRK5Y7lyWpZxsyMuC4sQ2FvSu+CG1eU14sZ/LUMP2e/3l1eDbHwBR
N9XZwwTNlxU6glY4ULCT0WXI4k1xWbOiFD3eOI8nV6ts984lrEz0tzqL2DQx39wS
xad4vckklb0J3bpLnWZfcm92fKXy4zvq0qGpZFxmd/7uHY/c0BjllKv2QzHms0P3
RgF/B21prDXDqoV16EMxybzFADdejA6pBHg5Y6uMFok7xEXYVhdl5s2a1kxvMMT5
KGTjQKyclv6pMEDzqnGrthXcdh95r/GinQ8rvXOvEY5R6ZI7TaDZ5mKMqlcUOGXB
NIu4k1QBvgiB+glAe8BVyTKWEt9NeddH+Np8O5aoqgQzNwoEyL2us/jWX32xSBCY
rYOfEogT1ccOTnmMmcQKf4t2ItmVIqNJXpwDQWID1H6Qk5cl5PyBj2tLNtlD7qeX
Mk8IjqmPlCCQ7MDrWiVT4bq4kzh1nDbckSY/7IujuIOsziweEf0921UzuFHRnyNe
+ZJdBbHMYpFWz5DdUnbxhvfUGKEZTebBQTwa95j0OEGIl9h1S7/sIjfzk/c5ZsVU
4cgJOWHBIkIeJnkwZLcvzbN1ZJeosYi2BwkiKbGXlWyrcDE6Z+aBztAcTtLumXfN
rJ9W6aq1QUOLIUlgMXTLGSQlI65uoRlTmE3VCtFHFQLEsA9DwNct/ha+I6lfYUYm
iAC3wQuvfzikHnGMT+xtwcrGFI87Wa08HKO0GjqnCAYpfieB8CkjZkxSjmIZ9xQz
LtAnbJmTt5pn6rQFMwqoK4FJ2cunjXk4S0bxQAmLhwd+jHBgCRke+g6deLF2wxIM
VsJvHPbwEw5nFjO1z5RtJYt+ZrqGAfuIb7FCKfnvTKPm6zlgVNAwDtpK+c4Tuqlb
qDG+T8JZqCCaL8l+mlw7OZkEdaxqz66kLbiK4KOTdlUILInBrUUH0R/nkZOAYEpN
/0fGWvfCPF4uDK9g9Xcwskns1q4Qh34P0mI0SYxmfqbf7+/hXQk+ESTTfMKd4IEc
/C4uo2MR7VAcGZsirvZxkwYJ4nFSLVLES3F+5ZFMcZdNasL3ghoBuSwpt2/A8u67
VapROVpOdI+54aSLMtVbdNMGI+kK4o8QnmsoensHL+Oe8M05delfUg+zMNt9gEfc
aK8SPZt+PLdrcW8YkEuipYffmLWjwfxLmEVc3axyZXGDGe72JDiiUdfN3v4SgX71
/UIULe5yINEhpWZLLbSqYuPeN0UjihptvXChswqqEjKKh64+23JzTY+gW5ilgVcu
NxN9TXq6WI73G3F0+r3ParJD6+SSPHfoy0eCAXLME4+yP3kQXwj5L9B6Gnqyt8TG
y2HmqWBPAsEfvn2dSXaqXHTcwyFN880CMIXiRlxhhYkCJ1voSqaKflSbkezjYH/M
Joo8e7zb781FK80C72jUpzdtztj7nW5ASMgiogIRyz2nHtS+aR0mRlUZcbl2bI/w
XxO8I09iAbfjp9SiJXdVohBd2VFKufzunqwS6Sakik0dxnR8zJor87Zy9mA5LzxC
BYjGGRDQcPHYQUtQQ7378WD+bjkniqWGHL6rlXx4/DufAkgfwQJdNBlm3LCFoiYH
/rk7Zyay/FKM/eE90+9y9DDu2sllPxKCMWeXtcTtGvA7NHYn+QOeRvenbBrYVHcE
GZ95VwXC7roG6xkrfp4tzJr8+25UcnJqO7Xg5cmnMD8pLkZxPPDKoYO6X+g2MJqa
FHjY5q6VMsxkHPkAUCBDp16wau3nUX/eoIDTB6oX16P3avH64JtuKwU+ygI+hU+7
su2WffqWig48jq4Dm0aaMe+sNsYkMB8DnN3vNo8vAIQfDRTB9Nw65+/GU0gk0qKr
lXJdaNAK2LVKF0cbv/jXD0eGvOTYWhAO5pcR16VTFFEPUUi5NWA59ubpaRc2QmAN
esmlK9aq1IjamevPXQgkmmxpXDnVDxoEHm+obMbGKoJ+wgjuhfOWr23y8wPoHs2e
zGnoFtRCD9yFX+qb+EqmRf/tNH/hXIcUajivaDKdr+Jn1zAKe2J+uVS7FvydOVXy
VIU7TD8hJx6Tl8YalIZe8LwssxGDeayhcZhZgJ8ZoMu9Igz/h/w7t+odvai+TQUE
t3xpMbtar3qJ9JU7JXA0PT2Je7nH6No0OTYoxftvuS/UGlXLIH1g7JBiGC0iTrYi
SBPG75MM8NNNiDrOiCxT2/ddthWJHI81VsOUZwtMJWEk5hywKfVAn4iD9wL3Kjrj
cifW7ZQ3ebzoEKjRuX5XZ7X/d6/JP2P1eLPPCudVHweWEl9Qld1LEU9X0yrnYJUP
ygpGF8rB0RlFbZcwUYW6tre4tYUUEL60HMPB6BQxUbKWdeD9EoCJWrmwgoXKBxRC
vZEAQnTSec0ppioSiJq+1sW5rE69pHhP5FAXZwYAlq6MWOUdZG8sTfdzEpENB2wc
D0nvscoP4d4U/SPtNnCq1Xb+s+br14WjcGRX5om7E9pPaS6j/NXG0SiLJxKhJ+PR
hQL68ZheotxySzaJx4PIUpzYEX750ug6PmkPlgwqy+rkr5EIdrTgVtaDNKgWe89R
e19L3kYsv1cfUzJ6xpiN9cb5waDNngD68ntk4wSm5XjH7lHp+HLIa6h/erdoVgtE
bWiUVw58Q4h0Xt+blLroQ9Hk4CVaSpjxHUytqAwxVSKpQ/ZOMrFwQ2LkjbxVkGGD
ykuo+k3tubX6LfC9xmHPG4IO7/YI5ADZWx1Bfndm5Cwf2DhIAx/f+boB0YNb6SaR
TuLdfUuvZlqMElS0Wr0AMNWO/dzp1V/GLRen8hEKChEN1XhEOsK1hdWg9G0rVcrI
QtpZJea6D4eofwQVmRnuBRW1mH+Zotb2PUfS15yTxU8RldgwAhjpAY17rGdV6hlH
fn/xVg99TdYlNaoreMQT749JcWvOmlcg7kYqasOVf3dSv6h2zPDH6DJbLmm/xSlP
G8YMt2T+/MvlgBxzsz8UEJi8mnKPJAvaEbODNYTURu0dSeRvWLHSMvVbslhhQVEE
cLcrcahYFcTIJaZFuILGCCk6TD7MimwhzTb8bhPLJ+gHJmFicbvqzmHJDliQ/aaJ
DYgx1BdTYl3+DY2WEI5ErQaOdq0cNMXUZMFrwF1nqBnBhXcpI52gpNbX9ORl7yid
FmgE8hP4+/pptQDHYqzmDFW0ir/CPdx/MAweWQRixPI8MMSOK6JTTqEW/QUGEeKo
0brCJl0t+3NsrCMtSwY0qLxfds0AB8cpH+zgHHJ5FWFsi1OOP7ukXCt1Af/lsG/y
q1A+KTd9Hcsj7aS5cKqXLNHbKU/tZTeRvT6fUhccxZtnezTn9HZEQdY6afGfXyPU
3gyTOL/4FiJF0kpwmAtl9/w9sFu+4O1gwRAERqMmr0l1wrICBVWZHVAZDwu3isFz
Z2cP6dOlFvy0Hi8FIQOxW2/ztNZ8fVME+jO2oKYk6Q1WuCgoBC2qu4t6Dcmpi15z
inJE1OgwAV0jPyCu4FzPorfelUy73s9icFy649rr4rUyr8wh9FLgRS1nADiLKJ3e
f/9jWNmd5NpmL73MUoxvYFD81qSKoOLRBkDy0whnzPORfJXLXmHE01/FETP/YyqZ
YGJkFOKfLRxL3ZRJ/46EIpZgG3qoBWCXMZeXk+4ukDJ5FObuCVlG8eDsa6drPbER
6he1cA0GMPA3LP+UbuARRSIFD6Bi2/qm66NFOTrpzx04x9U7dIIrXxKZrdCD3LIK
vmIuj32pqiGjatW+1nLWXFeLSHrvWGjb9MFxZGTWTSfVm56AV43Z0+lC5avQEE1a
VAu8ao5/22cAPXlb3RB2WjJrEqowgdhIiW/oHPg+XEGCjjHnAUPJSMUj/27BBf1c
sSTVcEyf7piB2qGYKrYHh4YhIgLEwNGM0Q7zPPJMIBhZAAiid0pR9CTh7RCqWjAH
SDucLeH3wTTlTHrd0QO1VbrtmTjLWEyHkiSDYxQQGVU=
`protect END_PROTECTED
