`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FkxI3zqV5cJ8DPaYospraWfp/ynyIF3Q6EujvOsHeY4VTieL+1bvUfdYo3FgLneh
PR1OzOsitQ/J2eyx7a91QVpogRAI1e6qPgL9hWgi1g+X0TFyvvGsNJbF9SEtkeDS
0w1lyhMI9DjQr7mNU9SI3ltAP98HGT4z/wuLwNy2fSeABJQwgBjUib+97XZxFcmy
qIbkPkH99CUGsYZW6ULEhs4zA2qtWpHsjt81qPlI4SNgwZz09BN78UMN6IeuaWSo
ByTy/vZuo5BcD85vAJ7hEk+WovkOI9kvi9sdO6eWHYrxdvu1NRGbITcJwHHNBchR
bW/Up6vpo9qYdIz/pusvs4iyq8Nlm4px5GxftjQMMRM3PxzJJhf1DraEs6Pk/HXa
PPEksS9XL7L097PGkXN9OvZYonqYfX92S2uJCq1qEbKluxvdelrMVjxIhvoWTseO
OEJZqXu5i1dbdiuqSW+ONvsGJ9f3sBAqW3K50yKutGhiszMZHz6bMbiNla2/h5Wt
ZWzhwOQdXmDjSh9R2bIZtfCeEM5AwtJvSP6nhOjuHEY=
`protect END_PROTECTED
