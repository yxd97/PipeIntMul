`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MQRGDYGLp+hDDNHdMiUVK6mq/vL6iHuajIsAy1QM9uGGY/4JwmTm5jhTCzELVkcF
DmAIPfFk7h2lgcWV8bmgxEKLDFey3chiT/gaCZXmofy39pUfgjLA72QRrbdbPpjq
LmV6in3ZzulgUM14asSfdC9Mr7l5ftbn8E8KK96qFw6wALmE6Q7Hj1Isps1Ov2+R
WVWU7a3dIihAfCzo6CNP/Z8ZvVRAX3CGno8dkHUbmtJ51pwSI9D/0qUWPY3RfEtD
p+oZXq0sDqAxfqKdtUfIl0Sqr7cKw3uLtulWwCUKRrrqNkBK/J6x7QUTaccZjXLe
O+8X7j+E7SQgPPckqQOAHNUiJIdxhwV2Nqry3OeFMlTfn1iaVgQIpg2dtU+i+m/x
ChQqxnM2xLhtctnI3h+y/OzTj9vPp0Xr9A8Z86oUrRDDlLUwLORgHLbEey+8MNmu
XUS+EQLeBvW3ZNrwJlwHvnD7kYUi9Td6zgWxnM07VLRgE4IykpUqpa6sMLWhv5ve
HcqY4N2ZCc8tzcUWM/ZymTXh8GxGXOZmV/JKupqkwM2dTvCBvsvqCKkinEnefN9d
1zW2/K7Ucwtb2BxBfzRe4Vj/3Bnbj2G1by1BdYTXbx7z2MvRg5i1FkxJTxdFe/mE
aOuYwHwgLwt99FWHV8nz0i3LoNGUZF3WDNmE7oS03R6Wn/IxLZaqtW8yGPIEqpCA
eqNn9iOs8kq2RPByoUTgaMWcq/7hlB0rbo8hJm48eIo1g1dlpFPUyLdtSbfwa5At
aeo5HINV+9R2RfqHmAUb7YoMNaLLQ23saDTJqL6MYeZc5/uuZl3JQDkGvnNnozEx
fbEsh0CPsh8Xzhc036BcLkTx1lkA6BtsESMq5TSsay85xy5K+D+4BdErfJhbtXKU
1eybJPeQRt20POScF4eH4GFsFj3IsMfYneod2yURVEKwQZ6VFUwgN3lY5Xk/vdyX
qaphzZJS4PYu4ROzKMG+ukKsCFrKUVxxzUHLrx2dveAeNKRubFAs3e+bYViMll2r
jNX/mjygCyeDRd9/O3VXlsGsWQ3GT7JapqeKmnIAT3D8P3xxL+fStFs1jHAsHo0M
n+VURccJg6MVLm3SWu7lYrfhAfkgiKsmN1D/JcjUxPCgw1x9ig1DJdNBQUoiy7qN
kguOQzM/aIJVhmJCoLjJB3BsmmQJE8FrSOwjYYSAU9sUGRBrKfPFqA4iAVo7QEbi
b0KisqswvBy+slIqMzWVvuq9PkmmqY6CTl378/op1iaIrAQlm3iNLlA4q0GvBIQH
gAl5fU73etzLa8DaOM61YCcQmFMMSAoBHXlSyFwipVhFtkVIyjSvTccc+t86RO64
nXko71Q+M0RxuMGNdSkQVeN3EBizMKvXWHhYpFdoEvihq7D4FdOUguEyRc5WITF0
HCvwiACNVI0JKJWupmx0CdHYf6NKFYHpXyi6jIErWB0D/3hAC2VqVMZTw0WF4Bdo
yhTQzM8RKKQNDhBXqSKhIjQwryevAl/a6TGBqxmsNn85u1YLQ8y+86TTgqPjS9IK
aGARPry+Q/9+NRAeEW4ofRhGFAzyuqteaVaWKmgKcvF+cj0T775MejzsoeX8wnns
j+1Wuq8lO38ftu/0YM2YxZ0KSsJ7Wn2sCJliKdsLj2GyC+PyMDO/4+FY8p2e2fed
WpWcS6AURIufObEtdK5sP922zwIh2M4xyLEKkiyuPErX2lz6W3BeuTvohCxHhMoh
8qLEsKICn2cwGTQnk6T+q/PegNS2ZbG1r5Y4SDqdTP5cIUlQmeTAOVQLMqySSYaj
KkJC2z38e+DdYI6KW+haxhXR9HaC6UrSApxgOQM3KKtyjL5vZ70J9uNfY4Psw/q2
1fxJBCacthSmqr6ZUAcXv1UzjT0A7FahZN+v2dsFHB8RATXcwOYeSqoDDYuzOpr3
GZVKxi1yFE3Gx/UPUxq2qLgiR20qN3KGlqZkXDTABvvXoZ46rBadgH+XLeQnXJGR
eqfwESE4AjagYdsF8I0DuKXKtPUvXDrtxGuGpXtO9rzy0gu1Cbf5fYVuHWoAH9tv
N0TD5hP+QyfQS+XJqbnCdHPP80IMM9q7nEvFmYcOJbSuoYJtQO641E3NkRhymb/N
++Y2CpgLsgWLIDNYEfOqkBlC560djIjg550mW41SwaLKTw2fohnqK0qvA+/tareP
ZfKbMjxqwu4a9atIeFpApA6fVLLeETHvYsgDr4YE199STaVYsu5Rbtd2hTzxawNX
DBuq9tbqkYl9gU08hgtfUUzqL1lq/HR4/79dkTe5XMf/EMtldeZMcO2gakH0CZX2
UiB/7+wkEXm22Qs6lMUycNdxzIYtvTEaUcfOO3UMhAZEMuhYzGL2lBDs/Ch3T06J
+W/bUWGmMtKll2GdKQKz92TiAgLtXzPnFaJjIb6ar/dgKZjeVFYZqRs26g+tBUYy
8GcsSKH1j97mAiP7w2zth6Jk3dNka2dWgmkvynyQDQMKCZDkkfS2WkC5vZVhkFxC
Iq6dyOxsdFGrxb1gWwBdEy7cQNqG+8yTUjhsVm5Q0sDr68RxNzd1vTeABuakK+zz
KxahuceZ3V6rZKJ/pi2alKxq89S6psYQsZIpsDJnZxeG3c4ED8SPM1mfhYvSdvaG
6Z5/Jixg8AG9RbVAn5LBlrlipaTvOKW+dcaGhGqPYAfoY8GU/FHNlUWAiavHTtMW
YJM5sH36KZkKZ2jaFoDl/owZudosNT2veSi1zjmoCOye8r7DvxxqRLW5VLzIwRJV
cyZYiw5DydMm0k0gFv0v5NiNKh4KrjYKt9MckdZKFIRL7iURX6qVfiID0tc1LhDC
I4R3tm/HjnJkiOsd56x78dF5OJH05pJXjUWWBP5OkJKHuH/ZANq9vIOiDBc+JNNq
+N6UQh0vD2YHmo2dQVX2Vf9H0tJVJTTppL+cPbU0n5tNOOoplcN4dbt2N91YpXqB
YSmvN3K6FpjQJomhHJ+imEivQtd9UXsBF5DOPqQPUozJSlFekUoBXf3FSDa+ZcIH
ZsAE9aPahchyWXansjbWnFjTPNWxOcrK+VhcN5VZVRWbghqJ523hu5SWA5mnq3IT
M10XSTKUF51fHHic7p4JdFeq0Rayd4ldp+HrRQdsPGmEz6/6kbI4sX6MnDkVhXmw
FnKC6XAG0ne4Zn3wrjrTi1yesHGVi40X4AXjIxoTdBkkhpg87sSbUllZLNbjSjXE
jAX42RpNj99ChDviwU4P/8WA7oTY7del1d/7QNl1HyBiEGFEb4EFDCnvNCALi90o
IJnX6YVs8odmaa5AZXIiColbslJMVD93kxw8P/Ys5pjlZwYJPTvyghOtmEN6gA4L
/COwx9V3otT1POm5V07pmJovzOf6T6ilAsXVP8l/NdWpG8SmS1+qsX6F47Q+zt79
pKTGoiZDsCd388y9uZX94rTmNwJfBlizP2NIcmDhss7I6QIIpt3CE9Ys5WQ2UVTf
xypGnSizDXez7aPznlwe5U5dy1vhyNZCQ0OFzSvHumQJKuwQkF0FNUOJZRtiorir
5Lf2MB6KuA2/Rkqnbj6yTIWsmcect5SMMuWhlRIHyfTbmE7OEBNV0opvYQHHy15g
1fm2AAayvTO5avqCL+11PhpHXgoxx1b+lJfwjcHFeTHxdey+gWw9tr6hNQG9O/9T
JqsFSVMG804quNvDXeWEd8jzLxm8ve4wchbrRMF0klrICXOLTIafzEuPmQ2LHjmI
codX2kdLf01pEk8lJfHqcjaB6ZiylsA1bUMqDIb8oCJHUVk0H11J5dsUIJunJP4V
UfT3P2iYw81oc1omIfH1/pXI4/ymzEVCprfWYBD0S3+Y3h3XpUpf7nDRVpc9fXzM
D5Oq8nY3nyjbg4+ettSHvIs6wMV/8rvd6Tx1eQnIk3baIWuujZGjSaBc6Cz01e1x
CvcaByvUiAnc2w6GkbVJ7u2QCgFsy+zyFtfzGM1rJAntAtnqH6QME8A48q7qRHAU
96SC9qzW9QOXjYo3F1ie/hckpdW5aLIqhjShgViZUmEmj5EVbrUoDTt896d0guEn
l35Ev38h6ChoT7+tf3a80scowsod7JqFBrnxiZta/WSXti8C+/TYLQS6eoJ/JCTp
xO/RHmVC5Bw1ElocEepcvoR5wSMhom+LuHxUZaaRhRcnF2aPuC+YyES1GuwaCeNO
vZBbFRnFP0tPN7p6obBvRmr7OGbud5xsq3+1F9KgUVaWTL30KjAnwzCXUtKgKUcz
PAkH8KFwJxfPQJ4rLrPXRNEtraIW6M0Q1q7zNEgYfieIpXYWWFwEEb5vxUWGs7S5
XqF1QZyJCnVkAHwuYi4n5GgZD/RaWVzm2bZlxo8QhrK35kQ8OTa32MxWppMaRBJH
zQyGe/dMUzoMwa2RZIvKylp/ZDXx8P4cSxfkdWTsd02zCsaK1yUysQ/6EkjCZJ2k
Yawt+sL/bwpHezhoFGmbHZ+sGxHIIhne0xRhd3QnVXVeiZMXUf0dTa4jLPVjpn0A
MpgdrBcYnJEA93pYuMJEst+nGj9rua29p2w25dG/z0qbIKEMknyK7qB/+KqS6uRm
N5lUOYRbgoLj5g9SaK32DJ+qJey8+Xw+xrS8MJ8VjIKicsojivEsPgyzIPJVdfJM
v6GAuu5tfHcb5Xahz8TjK1KvX9nmkYVLO58RtVKxzDUQO/MKszQyZEN1x8J6Zb+x
/pPVr4865+xHAgos9m7bYA0N1zGyKiizy17bxnWoTeVAPWo2zFBKkeiO56H+upfO
mBCfZNrajqsQkRorEbdLTB0BQPwCCVOW8jgutp30qtiaEWQXId+LrcejRFBYZYBi
ddhnOsa6uhBkRyjnjAA7HtZLWVHSgpyqlZbruDOp4r21ODiSGJezLMxzpvXqgI+t
tgWMy6zd8+ZYYJWcAv+DNOU1qXqvDvXxbdnsLZFjAzwSeJoXLOENtJqRTOPLFLDQ
V47ENGAtYwuScZruaFE3foUUGzmldLNtqzEGvqDEg7/t3kyOcUusT+gPNFVkk0CQ
onoNZ9kEOmoesumWGikSrWdfDaiXlGVXNO6O4RP3IuM3+jd9F73Rffa70PFmmq4i
9F/HJTePyeIn9BbyT/fuodHs6kNco6YeXMUFgz/KkdGL6+6wgfsepcS778wefWyf
znRFQk4hZGA7qaEQmYOse0d9Pe9e98qgq8WyuyaADMAIqO4BzSiLXHajvoUg2SIJ
L1MPQr1ZxVKnAwGCMZjDU/jzrL33dPq+JM1zg8uxjtzcFj25/WSRVRr2c+M88qzJ
50854lLiCRl5IcT/3gHI04IkzfoPoaluDBOjC/YouVm9Bmy5dO4N40SDHKDsWNET
RhRwhIZmiwG6maSMbqGvRE26IpTmR6fBjSZbMj/Qdv5anTpGZGzyDa4g+gGoFhT4
dTbkAM+MpAnY/Nw9g/UVW1vYCwRgcRUYK2MIcI1Niut2QrAQZ37S54CRHGTx3OC6
ymeOHO2RQYFx6v5FiGysLTkjvd0cqTC7AD3DxqdGM4QYDskQZIKtcTVvHDPkwUJQ
z7lDnE4lRwSMLXsBeHoqzvq1mxAYDiz6LaaoQSyoi4BVMrw423W9NY9rOwjdgL6Y
2hSYFrF97vvxBdCxA5pHKlgjqfHmeX+9ZoZWtUirKvsidFQchrL7Hsrh9SjZbz3k
X6soRzvxcuBBz1apkEYocNy9pQHZNa9AIqsFU/JfMKfhffOX1L46Yqr6V8dHbN7W
PJvO3r5gHrKm/pvKFb9GAmNfup3TCT8tVbWrE852kaUyksNnubIr7V3S5djT+OJS
7tlswDb2km6zaSsa1jQvIN1xY6s0iN8qP8iv6JBFF9C1T1hCT6scvgTGA0hFLSTX
/VQ/gfZhE7j4Jlpi6SLvAn4fZ4AqDdqKwMuDv3T29A0uIAWSGKIToVm+RMbiLxMr
rS8hwxp9DGNgMbQptGapHoG3uHS2eWOrerPZU8TLrt7FSw1AFpnIt9l1xK3iNNe4
5dI2C+G5c1rJGZUrFRXBYHnzJXaLmUVDTXXH0hjnH2uTZxR5wqJH1ffoDbvvqa/5
1oTHtGHx0urJqz549ObIGtSjBn52HYrhJleSdyhTFwAo39PZYzT4VFGamFTyT9qp
ar/lUsoKahjLEWMEhLZYqN0NMRR35AGXjyue31TVB+cqlHHKVTIScA1FaJ/QP0xd
lSqT7jZgEyQ50665KJbdPKZkhb3tVaGVZyOh/TuRanPXMwkDAeeLLAaE4qH++/2Q
GyjMn3LyLGnp7SNDn4THI2wNqVIMMFN/4ksgEnnyElrLPMLgx0ChpswZ2p900Ae4
BtFUYNBs8pG2tU2oxYdFXVPocJMPleWs12eOiw+FciMcU/J7W/XIvtmrRWLJiBzc
l8kOJO/6ZwfURYtZbEOqi46Uc6nHDQoxcikYC6kEZDgCPm+Cn3A07XgIGu/E+9sY
vWoWQyHFgd+7tftcb2yCuX4yXUWm5MKaet1zM1LTSe8ZWxlcQW4GpLCKLlodf+pL
SdCBQ1BSSCZKS89k4AIExDKm/iyJC4NW1HQsV65jmCwvStLKjY7UOLIcjZ6ennHT
mg72eSt3l2Q1COq1DBEdgQOCBwSj+insXjDpSppk41Nh8ylgfh0F2KMfLu2M7xpv
9MQ9KBYGLDQ8pywyTycjw7swGGzAVGAoNQEswfakGt8WFe73SkpGN+hVZgbkCJYI
3lg/4Qr9YC0FqX6c/H0FDl/xx8R7MvMxX4CtnrhzLe+xVAHjUZD5Nhd7E8leThrg
YnZ5YsAVDEE/mDZcu3o7a6zcBBghis+NKOzLCQeJXSA+Q2a6mS/IxP/WPHAH8e2C
Q0tHVuqr3BmRQxpF8xyS3aBXL3opvDo//FMt3OZnSQhQ78u5WsGL79wcbQhaKaTP
2JxBVUbtuMUD/OOdWLbNfNCIi/YcMq+TtNISbU0m91SM3YEAo4ylrjfJvjTsWW1N
EOB5VaCtA612gJMXelahP8Ok+jhZF71IAarHh4wJ5bGK+iuYZNXMQuxmPQy/PfP/
MeJ1d+Woue4IoLf3N2G4ogSADW/rxAesQI6Gj/jdQeOytfhJU7SMkujrE/egpokf
h/zuDantyfoGYIONqCtIdufWFmy9kuV7e+XCdPC1BD5Y/h20Z/5sDJuWRFNLyeYC
A9QLGpobC1BMgm/OsSUbFoIWCSatmPyGK5YPWePDk72o1jDyp0xL8gm3VgAI/0xw
a1GXmqHC9fcpstXatnpQEZ2gbh3C/Q/eXw8EdZfNgtz2VCVN444EAu5GMGqqqTyN
/NZvCeh+hUxzhlcgV4eZ+BIBfJS/D87CR1qJIdgTEwnhtkx0FknzpFIc+eMqQ7ez
MWgeagRL5pODotwItKk24DfxHAacB0a3PkBaAzPQtgZ/xqavXN8ppY17b5xOQrH9
FLczvF2b88o5fdHyoStl38h5vHURCzWV7tB8ghSobmmfXIJr0I5cYl4cO3vuNFPn
31j9pqhWA0Px/Xd/aCUDJovV7Qnnx7eHlzKJF1DnHJDSXs8UmDvDduejEaTWUOWt
MaSQ8EbF7KiYZI7azRxGKnlyBFtr7RhxUG/97oCVTf5Uyf+q1obmQDa4W2T7FX+r
bPbkd0DHtV1Lj+Js+k7aB55PFNz4FMCjqGzlE6Nwp84IW+GKeynHuKYrneH+z8KG
LC44Vb8aDe4pQFpRxc+Oi6My60ZO/wSOntHA8QxgrqRQIF5wQmpklU3z6VwwZzrQ
qLpjFhnyCA/VfB0ksVaWGQq/Ee+euJguCFi+OMo7tfjOAmPrOHvZurtw1/9pdlLC
thMuilhTKcYZuVkUc7sk44DONpd+oX2fDq52ZoNuOwYzexEnz4zLkTU1jk9oU7zW
16KXxcvV1y9sX1UJYZec+1c/NxJIf+PrcVdw0BTLwE0ezY0GjaABcronhd5ovvT5
ePdiu82qRT8A8u9ig/tbtOtLGkG3BRveKo9NsT9iUtbkLf5G+TURa4yZXXrf02Co
oB/oQ6S3XmTEOG9tbUwt/XW5bBBcDEkKYzp5NBQFopPccxaWHrvt21kPTmgv5WH9
paWeQCUHHogG9RkKSkoZVz4LWn0m92i1+vaQcZyB643vwDFrTRaRAdeQTPjhzmPe
4H9YbcUw5Odkfc1jwylkbC7+wC7gBqsIm+Dcifb21uP5OSxJGBgzN7Vlq1/vxsU7
SmxV4DLpPDZqJaFecEvfBd6+yLgATonM7zbFiGLVDrwGqmYK2w3XEJxZ/sWtioKB
pFJT2a8pA1R33iJpEA7U51dNcoV2QN1ONmh0b5HOtYtprwUtaNijWy+zwPLLqzfY
OkOTqLCI3Gp1pvJ/z4JvLrMOU/GuBIaIa3TVfGucyIv7oMmhVgFppUe5/7epFB4+
S7pqWBQCksfcitRiLq2HH3xtKzD1vp2gBzm8sRAoiX9tWzwRjvKqYyZ3BjwDOc3B
uieU8ay7IXHMyjPK6v76KYxzjnuFUEH9BNAU8qPdg6ruvYX5oMO3uQaiqvbpKtHn
Ln6QD9jygtqspw5FNA6ay431JrQfr4qvHMV9hhs3R9vc+9H01M4fEyC46sHq8nsl
ValzOakC3wJ4iriMffQvI68Ssfph9XW26lbmwG1l6YbHS8KEqa9+EnhpoTwGOjlX
b1Jca5x4t6EUI3iYBUvFP66O3MCXpbt9PgwjEPqUkXKV5bz6Y+MHW8PVc2nddVUe
M/Mbwk4GwzRbpmMlSHdavwgoh8loWpLO8CPEJ1CKKRMYRVrBwRzrHZ/SF34CNRy0
UDmG46L9URHFqwEML2gsibNusPDTbBiGyf2UvmdzW/N06kRpiuVpwS/KDUOpThq9
NBjjtPtvkB3xTzwsvpcdxIs7eu9bGcdzIU3nrIGhPJ0f28YNoMdgdhaXS42knLb1
dCjqQTLVslvzO46DBEV9GOKKHxUa4tM27RuUFLgSHJmVLhP9cx45rPjbjs7lFqhg
p3/ABNzc5xbmbKuw7PLMVXW51DjVVspdh0KAtSyTvEnX4Bl0DI8HC1nDEo2ufxp+
M+TAnyhneYGsBaB2v1M2zQto8WiTEMx8uQpO70ATwP8ISdqsZdkqirbfccdRRch0
v/RqS1QdbAKUtYIph3SlAGygaSvXJlv0jXCaWCieIczxUx2Bx8d/ALMCFkWqMzo9
RHQ2fPeZwxEekSlEcGJoYsttricZJnLHmTdtYV6faE4gxfnjYRhhP5TL9KKRHV+i
uxCLpKpPOOmkjMIMMKSwmravOzNetgtHSr45jHeyfL3W0l1J2JMGoonBCTygoAPp
Jirza6RG6eLh8ZTtx0ZePJDEQw/RktVFWk0NtycxzSNfYtCmIvgPII2SjlpxS/Bq
MyqGHSOUC0e3Nu3OtyfIrx9xQSAaGkkBnO8o+ipiHxW+LdvWwJJBO8irkU7ka1ux
7SPzn8ZmT2iLsCZWHgJ+jkE89PJGZjUiQApYnILEqj/t3ZLbp208XKS0Qr9eng/R
9srbCw/ZL2+1RzFyCljWrSCGJOQ/n+ivp79SUvsNJFC0HzogYoiJlAh3D5V8JzLB
I1ouP786I3z9BfhiWF69htHM3Gbo8GsVnt499eXqySb0IeB6Dg/6KWmKgQnQnIK8
QF4fXnb4yXk2hp54abb164NFSQYa/DBbYVF2y3pypzO5qpBwI9s7mjAFw23qIFx2
+D4WyvB3QYDSVm3/dcVpTOAe18q57Gpzoj8O/ivfbRIWkp2vFvWc4/MkntcbAL/D
M8/6yea4yP+XEFs8NIh1yOGdBnBjHXKpbPu14kcmg3AZTt3MlWxmorhb2qOozel7
jdKPIUlT71AQygvrGyUdGRsz9SXIFrbKzrKeyZfBdSY3Tx5r/fLvgkzzhlzx6nmt
TwD9slGJztJwDn3/N4i69PC11RAAd3DlfHtsOe+ZVUP+A7Q3d2flWT6LSkbtuJ0j
OFl5QmNIQLj/1hGCP0OH3KZ4Z+kPgI2lpUjXFtHmTPkenYQY7j2GPC6DSjk6gMFz
ssshqoNbiBF8VEzG9CfpD47IeqHwKxuXn+O6NvkYa9qvtk5oD6ce6w0Xm2GzJkSH
ztE0nhG8nKbdOE+9Z49srSiwuMDECZNxDiXSTbxGYQRGvP5Yb7krK3djcBTtyiWx
n/iRAdzwBEPnEqKjHlK6fwD1uXCj1igFqno/cxJoxlpiByrO32qeQ/smtpYSkrVL
Ex5uyp/KqHLzajEasoMBzwfaYAyEWwiz+Wb++fH35rq3spFI8bg80G80V4wNmu/Z
+/38eKUM7qBfjkMNmph1BhUUhNU3JbnN/QJqsrNSVtSN3exVO0gijcsy+Fie8CPc
JgLwVwLb+pd5+lNw+T3/KCINWNFmTSljjbwrA86EgVRdmbkcxqj8jlIjZbpppMum
VSb5ms7QlMkdxTdi/l6/7Mpl1AckUvMzN1HTAxTjlPaZd1nPCKnAWMq0S69iPuLd
W0pXNx75xzIEVox46cd0oCzIEuKdDHCfPwI0kjjymOitWpPIdVFmXGJokyH5ZtNP
ibDAQioo4VmqlSlO/5bFRy8/bgJvyMz8gqjlbQNFrpJ+dQVvJQbnft4+gzqYIbni
uTJYdDaO9mmI/Uweh5bg53NsC2TvNgcvuCF+vCauHoW31V45cPjTkxBuFiq3f75I
M+jV4aP5hw1r5Jpcw9pyMjnh9lnIlqMxseCNg3jrFYqZFbhusLBv72Rchrkcp0VN
jVhZiMqv85ZxtxMXErAHNR8DPcGAWLHb03LqH6a00trTM6Lch0iDxge+l9FQw04C
7Rmi7bXV0RPloMC9c8ChSFvBIu8nz98qqqLhVJdSQorUP5sfrQkDHy6Bffexgez8
+oAIX8LYRM1LHa6hY689uQgrPjn/6ntXu53zbR9jWfh4DA9/wMhYFcQswCkDz+it
ngNsrxDpJXH78+p2UNMGkbL0jVLt2Sz2gXKeGPy0A3/3lj3/rfPHcIQRMsjldUG0
uSC+U1IAWhDF7oNynHWOE2DqDi1aRhAsguN/vSM0gc+oPNDfQ9IQOJ6QrHNJ0167
81vewgEbA28jB5PJf6h3BJ5eJKqY6zSUBVeKiSUQ6WuuPyi9jAawoH7TPTj0Vvi4
cKF+yw6sZ/bM+ZWeWyjVJ+mt/Bz4LyNwHCrxLqcSWmb2UKeRED7vpwiMFdECLPvb
IbSf0aGRFkswIsVgM0Jij64cJhDiPx4q0vwGcOZVUkOAL1nRRHmlX4T7RpJ0FbQ6
RhfQ6jZw8+M0MzuV0UEAoRKVqGkxvDMo4T+hnaFu35Y6HsnCTsfMHzomAjIoGjIC
kQtbL+IARUw7lDHH5XgY4sFUf667hYmz9soNueVnnlrkouZ7GGmafcm1KRmjrY30
X4DKh2mLlGRhBNkcnslNyc6N6eX8le6qieQn4F7Ko4ajVj61a7MKpFnimWHYSOzb
2JeNaxd5LTKaM7GiC32evc4lQUyZpdH5f5Cf6deN8vGEmYnyzEWVnq8lh7hohJge
Lvb128cyDzvOALahxhAhV9LaRrXQbRuc7iPa+7SrfD+PgaFAudJXlyc+o/aDcsOl
j+0pozYRwPEK90AJUAEDNBJb4XGApKmWsXNTkfHwwYlrYQ2J8XBKDysxjl5MD/s2
bnvuVQ/1NaOL5EeS04Be5jCZKXall+yFG6df26oNaXmXKXIrZVJROqDV7MbXCD5P
fq6iG0A7yfSM1jspEwyEL6Gk/r2dFDU3Nbhapayt2Y78woABmTfnJSf642hkP4ml
rlKmb/aLEUFpEQ3/S4dhZ9W8m2KB/AROd2GZZtil4mdUBUsIGyE2+vwHvetZSPg6
9gpKKw4FdGtQUoO5OF82uEXIE1dJ+90oajui0s/H+/eBnc+xZqSnlm2mwTRmUp5f
dRwy+6xzBCMY4dtx2aT24YwNET7nLbtZx3PH5eeclXxbY/02gTYDBXyS4lFgdP6x
dKmx+EtA+c5+9yR9ryprB8mL92X10v8y2jsKiutGwNAk3bjXB6r68gvAE1gEYVzM
vutuHp5H0Wi7QuB5BZSWkqgaDOpILnSyY4gSWpU2m8MCRCj7do66zqhPEwUY2L4K
N3IrXeTGFm+YU9ydMB0q/LjQEW+BC+2NZd5TExqQ561M/sJeWIU4/sUNKnY0nUQq
86D81Ggh/m+ViddUVb5RcOSMBwWO8wVP149GMC3iVidzwLuozXP8Y6yVPjisawwj
3AFun3N4Ep5JGGN1zsvRqFza8JJpcydyLeRVSk5I64FDuzY8/YNxpbY5p9cC3xXq
SRTeDZA+ZHeL8O0fAWs9LCV0KPsW/wDhWCNV2mHEHosmOdCJT3aQ9ng7GiOizM4T
yij8H/lEcwpTKpmR/BK9gc1bOsXdV+YVnja+rwjLJISTyMgn5nylq6RgSce7Hu6b
ee9qM9a8fPj0jZtlZAh3FLRt5613yPB9+u2AskpBrQZb+YlAKn7mtBMwqNuijmjc
/tlen+RjFUP2l9gezQq0uCJrjE7P142GMiiLSfJInBlBcxxt5FpuiKCcLPPWjwPl
9o18D3eqgsDoXtoKzUuNg1sa9QmOnOHttGw2Ml/wERPOduZeGiZkrwN0xnUh8Gxd
Bxv+Vw0wON65uDuBI27bjs6e8DnCQSYCYakeQHeWZlfiVnSc8wPDFKwtFwjqWJy6
yOOVQv7iGrA+YWeVH6+7eDGxEAwkhF/mbZ3Po+TM9ib5x2EaPn+TIOOXy1I1JTnP
MX90eZ4XmSnq26CNbxgcvlxgHejsOYsCkzDXRE91Vq2cL5hRvZ74dAd1uW4ymgmA
IQvoL/j+EBwKEv1SIajfA6r9+Arx2ug0OIlavuiHZ+XzGRAUyfIPvFiD/umt/Xx5
vd8pCqmQl43DS0JBvWYW7cdcPWzBCaE5Bozz9GHmah1LD4RtefA8BwpMUJI1Gv9+
Myv1aOy84/i7ltATohFXzy4AtdeBVyyKhqaNinodRJUWeJ36Uiggo9G2k7MG4a/A
0WQRGtP4dBJ0M1heiZwUxCCobL33Hw79B1TX5EpkJkJLnQYzYwrLvKYexOOYfENN
5EH86P85MunFh1sSXiDBNIbOoqAyc7d+Jb8co5CAO/ltj1pTdF3IAmlJkBsvsOg5
1savbx8bSTvJthN5sZmQjkS1KYNDu+W9m0ypkHFjGA4+Wl8Fn0HgSoHhpjGmEXYF
+uT2V2Hi9YLVFjNLPvniAeQLTgPLeMPRgZ3zyoS2nQu4eTbSln+6Y3kRCg65kEHz
2fECsFwUu+4IztyRHIEtOEferS+lK1W++c7Xu5ykGgBzjSY5O2tcpwbkiN0U8dZs
nlyzRF8SuhmYf9Hqj28s0u9n8eyCGg49r7GUNe+m+KGlGUWzC1TMybqkLtOaib7E
nPxhTIjHCNvQla4z6TzrT547r1iEYhV8Pzy47Wc6MTL/WnuPq/Z6HxL5XOeI2CtX
/CvHng/QW/XepGwsYGaYQeDy7ryE3YuHl1Qr8mKlf7Soz+JW4R/0EvIfNJxqybB1
lGrtH653DpZ7Ls+09irLMUYrr+TXB2CNC+wvGDsvxPeX/ffjB9FRABBXMuc4On4P
2Iaie8537NoMnKMcDxpQpmaVinvUUFhphmaCoJxuLBMkS4uxx2VG76t72467dMOL
oU5Rd+4QWCxU1RMxYcBcXlUTSS2EO/eCbEJ85hiuB/mF+qq2G6YNVYFW7ymwa+rq
RGWGIeSU7epwOH1oA39zyUp/jiF89Lv5XoxjAsjXJ8DdFCDYhmnfBCG3k5qLIMWX
RcW+IlJqhpuKiK4zYZiboOZN3n+SHOURBEX9sNKuACZ+d0Wwvk9V6WGeVmURKHVg
0gwZzAvMx7bmCDRp2+rAx6l/TnjS4XWwlMcvOfPkXaGXgpD9lIOolHqCieELsgnH
EquZ6DJrrKLfxBExAw/kne4e1zuQfMs3mOaCVfz2svpTU1Mx6+NpHzYlWolcEPKt
ePABb3Bc2gGm8hJHhAWT55Lb6z6BCVZRJ0w/K1RJSzvpBgD/taB48BggXA0QTmK/
+mJ2vRJpTYQl273kLp5KK5F9vCANMRWUcxf3Lnh/XmJYv88vlLsNUbatca2YqdEx
+g84Rd0iqKWaCW2roCwtThiSEOI+YMuI3scRbWZonkx/LDoUpDrIvD5sKFXCdHNK
LDqI7L3hjXF66lXVEjLRJOGaCVZD1u4qA1NqYgv+ZFxQgyDvZbi3xnAh8T+EVpx4
wxFeSzuz2VMAm9awGsfaoYwT8Fi1RtM9OhHFkfuswsKBY2Q4cjU2dQeCuZIS9zpL
4+1FT9ISf8TRfCDalkKTKdv0lhL76YeSyngXSkMASfxa0DRpy7VNF+K37PrC6lN+
d8VFTktIwaFoVnHZ+JC7IMcsCHaHO06vf0rqnEdjAbfOAIldd+LGt868nsiWQP0r
q9SMwyKJ5rQIvd2O620C+SMqik9xW6vpkfWMd4HAcQzhGFlbijHI4rdPcWqT48x0
znBuecCwX90ql5Q9XrOrSBqr6jQXOvnJDgEm7F7IE2Y9PXKTR27gxSionlTAyJd1
L1uxDk835QMzEqxv6d3iEX6VejDpTZfAUc+SKVjArt5Qaw3xUht30fjfd5+RIs8v
gHppMd9LGrttLKDKf2fS2T3q4H0uP8GQEfEylbkJUiXASv/EfyF8x6gnleEBwBFX
7jJw6sdn10JlTIhZY68TRsjpncVlxvOUwsaDdiPLftKN7V/CxypjZOEAWUWXMoUc
3Yj1mhjuttAl+0S3XyAUR/P2XH2x8uZG9WO07H2gL9RH23FqDB03/9euyzC9gk/S
2iNrpbnSGto8VTFPX+jTt4auT1VluKTY1KsWQYvgMEKT9SmqaeN2xvZrtavGqVd9
Bd4Je9OZNPey6Jho8XTbfMYqRGTqUxUvaKtIfrpuSBl+5pg+VR/HwOl8qHiTcI9o
wRLb2OAJhRtErAlaqFwUzXL+mgLE+LqndVPupeVRiiq+EG1gfFmdM5ceut0xIiUi
Oa/IWqFJHQhSEMFLKbTxjdy56N7vU8U0tveOd7bNIkpmOMR7F7JLwBVGj05KMER/
STo4km5/sTiq8aLoWAPkrPzmHkrU5QUn7AFIomYHkh+UanpwSh3Q13kFbLi6AHaR
m9MEaCrGcKa2XxkeoxvCCLQfNBZ1Zcpfr+jCY/zbaNIB1gBAZxW3Kdg9pnoy+B3P
2UfTAXUH6HhcItilcukBAOczHjdZf2ue/Cuck+FqSDgL9OvO/zKeoeTjyvvK0Mgw
Uu2aSBdY/mG3SQNYhwOBhaTSqLiGF6NYw0mDPojLPh4kYzMsnzMVHkk9WqVjkINA
GIzh2xmC0xek/CBOEFuBj84r08ox8VMZIGG0PglZSWpQJlq8Oa8ZM0QST/ZGrbJQ
UE5nlIBmo4NVLOhV3fQU7XRCKW1a3jIqwpeIt4VYCFuM1A7Efu4qLGYQARkrAvZn
ZPKbgNkGkmrvlyIPtJ7U3cPVVbDSGZrUiL8BnxKcz6QcCyNa12HuFlTvh216kWuj
IIi4i3hp99KxofgQ4cyMiVHp9erjVUAhwyXDI5sMXI1oh8LWrW7AJYmVVtrgWU2f
aJlYyfAZ464kCYolDL+Kx1vPNKi9MdmtOrpC7D7hctsPiZ2yp2EyL500gvT9Azc5
iVF9U9WrRVcMInhnr8OgXgq+mrw1Kljn6JcjuNCZ/fNqD87dTLimmJZQjXi/8+oj
CMZfKP9KIRdpIclY3LIfZ7RzcCZ1ZRbDChJNXTkrSXg2lMexrTrllOLULgAafqum
SGCsEip4iMMYgfMwxZkbxH6Nd+EsOKYiAimKMw5R1nbWvI0/KKyhOLFNsvBO3JRG
tOki5ZnVIB0Vhge0Sr5swZX9W1ykVn7Z4BiiawvAkB9C2BlUJQZ2C+DkfZFvJSDS
bzM31gTKgEV68v9mMBzbu0InIG3PB/4ndfK0gtvFyMOamCes4JBHJF2P0Hw5CcS9
ebj85gVFC/eZ9Dw24PkOBeRDAr77DTNflzdDp0spdhL+BziKEcuVngY2qGp9G3H8
X/gCsaOjzlJSB9oirBqlarcHTxUd6dcDXje5b1uGLtID3/K50KaW6x+9hppUsK1Y
Q9DYV1JE3ZjvS/zEt6lXmejuNm5uG7Xul4w3ioPpZQKW7xgPA2SIFyjCX0gDG8ia
0SZvarQMZ1OdKHVLq4e58eizVs5HS/DAnMRdyfYK8AMgMBmPNrBw8Ic0BlW6opjW
pIPRFTAHnlmvxUhWgXO0g4PD2s+I7hdJh+k/a2mxMKQCAWKR3+3ExYIuJSSOIrmk
uwJjzqYX10SZbSh8v5XJUM5OAtA9Zw6NzLpAAynmRSAY6+JC/IYrJVi4xCxT5BuV
T2kGlE9wYywAGpzWyAjHmPJHvgIGwIBYRA65vvDeraDUPNKpHScVHojfpvafhNfk
3T7cWVlO8WyiwMAcPE9oYVEQFDAMSD3VUEA7rvlCcox8bIioaDsAiNVnCp6xmbLT
rcHqmAWDjwIzSzj3AScXumeFGrdyi+QpWxjAasLkbwWjk5P420XFfdk1OE/kFvBZ
F8qVvcaC4nZTBE5dg/d3AWkXdBEiI0zIOPKvqt+A4n1d8N/rMCoskfH4aybGprrk
xJ7CtfbJrnZJlhuo7YsuZWjYpiNR718PmUhNy2VrxWkC0zfo4qs6zAL4PFFXGc5P
Hys3NzPuJFTIMCAjelK+SwJp3RAetqTAApHe8WHChQUnMGQfpAafrbnTdU3FTaPW
ylYloJ+bKrk5sRxT5dPAXK0Ccg/NzLjG6p1qFnhmNWiRRRAGOqP/ubIUCQ/HU1tT
ka2JHXKUyikb3X+ffUjWt8XYwjdRmMqxP4+K01wv15CU1sKz8YpY7tldi+TJc8kG
wxQMkTs2r1uZ41oVhQ7/64KrRtbDwuQtBsFXeWM9/npkrZX9AaShLtdErB28hg/q
S3vLlJNO/Q82MKORZOWBhxnTR83qPAFJm4KGG4P9nQlnIlfSO4mRiVWGY190CeX2
qiiU38HkODHKB0lc30u9oTiRaOve/FK2NNy1Lu5PRAGfZb4jJr695d5Qe+FUZy6h
NfnkKX5A4oeBL0PHaMbr5BTwc+3xPEUqFVdujf3OlCI0jHqtmGzNv287Cp8eT1sU
gwhvxuwDRifoKPs+mc+suyp+9xBeAVQzWxuOd0OFHjrJ0quriN19cUo76S0PezRw
rcqTiSzrvnZdjljRbCRbcjPpBEoRKC3Z3XIn4D3bCk1bFpn/u+IYK7RNRJOawRWJ
01lCK2w1cV730iRmgILidje9/yi266KmZOjzJEfJhiBygZ/PwTTC95saZmB8Xo+0
U6RcybGayFtNzZRSdF9dFVZBcd5lqAQM468v1nSMKooBAs+OtWjypxQS1S395hKY
Q8OoU/tn3+JA2tiDAzrc16C1y2Xp3S2Y1K6IKOdG281fuxG2vZuj3dPlB+30OaZl
MhKkQ0i8UukKs/k1486ff09WVIae6eC+jFRLcgJDNdRuaW4elIbftGxJD53/NyyS
JV2A9Y1/dl1eP6TN7VVIUYF4bRZLS69ettTjRbOH4jI=
`protect END_PROTECTED
