`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xt02p1hsttHEAwY3YhbFVe0i5pGCaXrsi5SGLnvOh2rVjTYfp9DYQdAUA1Vn4GZ/
VRP3B+yiB6MifEKLMZ466HyjagvRd/UucCNEue2tqrW+F8LkgbxvtULS6QQfkUUz
7GJlnysyQiCVvJ6r72qbVlMS2VV54iTsXUnzPYrUvms8wm/sv0j/xweVWqiLDK0N
MRF1N377M+v6KpJKYJ3YTCP/6F2ggjY79hERgkQk+qncDI4K6FI2FBo4+YB5rZhm
4yJi2YvYVP1GHCGxH2Heq86OCzLmTRl04auLSaWTQouQDYS34T58INOEz+N+crBc
UiGOdfKu0zVgcqp0RqBIQlscoB/Hz/Eywwo+6+5KgXM0ihfsuPEHNHvuWf5ZabjO
y4RGWDZCT8KY8iDA+vdmpQ==
`protect END_PROTECTED
