`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LH8z2IUPIHSzE3vSKVDNWcRxbPerapj+5wd7/BJK/tEXMpCCTLWSTqY/X6l88add
kTq+CJ2cgK5ahmStM9XCxDA8W7b3sEJ+Q/DobjRJ7G3llIaWdCxBCRu1QMMGja9m
9yxc9mQb4H7bHpFhfAL+czbgtpk/ItNau7iJXPZhNHZLly3bijMe7xuqJDAFBMxL
pc1k/PuoH35mMM0IPWwM+NK3u1cbplF4zgvGvyaYof6pDVaA3ZXDuVVHJcKzX5pt
gpjt/DBmbyk1sj9Te1HnQwLPZCo/O9XrJcC3xhEHfC0XNQXNTBTA240T6M/Xf6Pa
G/5sMQtqlaQC/HHsS0Z1o2rfpDqsEvKuYjV/5skjF5NwJzFgVY5tAb3Owi9sMjvV
fppm8XIXekpZGqxJbcbTnchWkjrdnnPPfe6pXgtwMZnNFxvz0BIsfA1y0IUfVd5w
hg0RJ+sgZfQk6UxMckCdS26JumqRw2Pcc8mskrcH1brWYoDXUkDQ7qoy3SUXhtb0
4p5AfM6aE818tWI2w5o9sEzIMSc3ejTJClXl8ROr/2Iw0pqJIpca7E39dIikynts
pStPaVLj800gHzr4SjkugjN0yNLYl0qWsUp5ZGGeCmfo4kqFKQkyYaFobWPdL/lZ
eldqHxzE2caFL4IVNWSdKlA1lbZWS5OcPUYX50DKnjuWqlFpsC9GBl86lnCu4IMl
uG8Xgcg0RQCDHBhRuPmD/qftfBY0hcz/4ecEQHPtlP+ihRYXGamwgtTQr10bZccZ
sAyHJU7bwhbHo1glGvOvEDQqG+Vf6t5pXvygP/yDE2gKDvfE02pk/XoII0OL/cxk
EByzRPH1+hUknkcqU3UefFWSCvixR3TjdrcjIzJpYwHKoqHIOxRoUC0uEwPUjgYH
T0wS+83MJ06DfYOWyLtZGvvj9O89km+5E2tdZbAlSerz0gOSEfYa2YuAT8/OwGdU
6T1rC6FYxnWsoVvzudsMhp2Vhg362NiL3YOEEETw9hDbTMKjp3MsL23LY5dSHwm3
K8W8aH0sTH/rSCYGr3uqS7CJUKQjra/0flb6sEaJRKFaWqnd+DIHyvk/wxCmZiYc
0bOTWBm/RjJpG4UHvkoyq+y72JXD0pQit5WLEWnKqqptu9dAlnHUrKj0VheoAXXD
mGDENdPkj73He+1jN4mbA+XChdFOIKjuiYdXI5ObGDcqNfPCbXfWA0gufgb7lQQ/
CQVp9qGD3hVorE2FCM8ontsOpSrsPS/uIbzsZZz4XUGa+ePCmTOtyEvwUMgsCM6C
JniAZZN6MsktmL3CqdvYuA==
`protect END_PROTECTED
