`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmk0hXF5grae2uOqmCFSbTHIZqUlaFR5i87X1MQ4+2TJcs423SYRPGc3zfQBGT8L
mEucMBZRwmYbmqP2rV6ASe0/VnKWPp/r0/7s3EvfHLRXWHd7sZjmlt29zh65tvLW
m9PLzyXdgrIbCjSxd1E+Fjc4bFNrAEA8YEn8OS754INZArAQctMdqr0sNWoWN+a2
f1yUo7W/jGOMUetgW93567miHzPihoJweYHsjzWD2Dy+TqtbUjzPAx7hwV9g/v9h
bJ82t9obpKT63R4lEE3TPp4ZWDfUgf40ps7ybjoibKLMft941i1HXoXZTP8/6chV
EwQyUblYo5y49u14zUgJA2E8SK204bC8OAE6g8Az4UYgfdvxnNZGPVexuRvK68LY
ZUOVdYXyzsExnZu4QZY8VQk2ApWiJODaHL92IMsJkwaEGejL0HZpfumzDsRImxfV
PD1LKhmQZ+P5JCL9Prv+3eJpfvGOOHErRAeNCLJYcb6kkKCdrXv2JrVQD6f3U4TO
EZDvcePDpSR/MUYBLJGfdOn+dSEzuQ0i5t9QclNuJ938o8608XuelOCpXMrgjKiT
3UabAxv3szfH7Tvwe0GM8Cq2d0xmSs/UlvK0WYXycnEwaeEd2H6DByMhY2ODcn/6
KaDIlgmHno+qc7YzRLW3ug==
`protect END_PROTECTED
