`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RMSTipmX3+gJfn0pAbcNfR8ikCnpJMyFB6hEbB+vUOoJRoOUFN6CgEIOZDEom4f5
NOhVo1gnchVM8f2g8GfxgBKtg3C7wIzHmlxmwWTZ1lCe904kQsT3DWhEZaLqfnvf
0RVqgTBmbdelqRpbm7hKLRdUVTIXtxLzBwN5AemGglHnEHvdJZPnqkY75raUpQyh
46aK68jNo9QPZqjgcJN2BucTuGYNJg0u/DmqUxYFkMOLByXYOjYuUJG7u83TJf9e
SfKfI1IP0A4hrs5hm6kQ0cWemWPfcdysvHNGud/yUfUnpIsH7dpLbjkaWv5LoXaV
DX7F+AgU5l/Cp5OgwlsUQCXHz+rQLJzHgd8MqjueOb9n9ydPZLcI1PqDxR595Qh8
+DcBhoFjlescM2ZKCrHRdOLFMOMY2lTujs6Cexa7wWiGtxisCQT5HMFGgAxdnUS7
B7YDCWibTYCT2w5yoau1WfQIQcm42E9vewtT5lkJsOj5KM6rTPvlumLWvfx4txdJ
9OU0w75mSXkTENgdNBGf6HItFRuLirR5oi4HpRJNiuMoiuiXe4KXh/vDFUBZZimg
oSXb1522IsMnWsxezRADTSfbE2QHv9K06kehwiNqlLUxGkATioAQdS56VvlKW2ak
5VkTC0+0bJRKvPCfHcct9thvX7PK+IqWWPqnqqGlTgs6c2L9puxRs4t+CfSxvM9w
I0qF7Zu/bpdn7hH6o4CrdtLm/YAKHH5V6AB/msdjEkg0/If11UClLUQCfrHT4UfU
W2R7NC+BsVqcoIoAihxf+qDoLR78mFMOwVrOXDtdViojqZQFmVxwRTzr6ZuKbp9j
pj7Bd/SNfgSJuBa7byzUHyiYCNqqpyz861guYjWTC7XDVSLOt3CfmmPORWiThHe2
OTnaDZcd8LmPz5eeF9q1MU/gEYsEwljXFYa1+pGBjmKAAcHZy3hvX5t17B8reZwz
ckJoOj/f4AAkH0nkS3Zk6iU/sCPll3liANaVWPSpZNrtVjDW2MmpVbYJUazv9YJT
W5bAer+fMkUJeAE89aIhvBsujjRm8B6D8QCY9HuPe4cnyGoDySFHO2OZp3TKdD7m
QgMwfXMY78ceR95OuKkR+BI6JKmRY8tRONbfE0VWGTDR3rPxr+kfAN4LLobXoJrh
2rsCZvqSm5SBl6pXeI4P1leaNUGAaHUKR24wkX+4bSGMWCU9H/yhAduMEcxKWaOr
a06DYrF9b/D3UPCsI5u0zdwltUKx8Kc2MQWalZkei+waCDojrnERyNleRb4Fc2jQ
7PIbzdsHPuhvtZQWpL1iUFbQrPlFooDrzzWk6oGYrsV6J73ja/vARD78sXCnjfjb
cM1VxAa0xBpc5C3OBKB70vtRZnZxNG8xcurrvPHZDEvd49kzVAP3jonWl6qICfC+
zfZ/EQ1MpStuCcs7kb/Fh/pYTKI9ejkxkgCNx8dD0mtFn0OzEM7kaOEP/XTE4nJk
BHxS61zNVpihSUs43ZWcSA+/R1191dY+I+BxQsszf6Arv5KaKobQTVpGnDEX5cLh
o1oxYVLG36SPPYJMo8t3vkkP1u/yr2uUD/zjXZOSFFARoqHfp+ucvL5F1xOofPiR
`protect END_PROTECTED
