`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DR7rM+FOP3JRO5DCAhxrq6mGqI+sY9czuPsfW6dUkP4xAHmwiDNw01tHno0rvyA9
Xskqitx8OxutEw75PmwS01vSKGYHnvy2Z8BcRQ+HLdO72cJtrxqUz26KOgBDkRRy
D7UZM/UH+vN29wu+EvTNctS21AGUNl/QHibTjdULzWlNIac1k8u48hA0Xz7W48bx
ypUA/W04V8Gl5x/dvBXdsTXEuk7V69PHBgsHIr0hpeLkrklDSOM8nFmUFZMVSMog
SgpdkU60FEk0l9y5PxVag3ryb9iDokUOEpkdifGoUq1RHELPkfiguf+p4GUBNgE7
jT6QQmzWZQz6N7R2e8yS5AWnVygbQVUUI7ZNmUNL+7avb5GklpM+nba26pKzi1Wa
MJWDBnWWO+jDCvxXDcZNao5YsB0V4ZEoJuneztwaBU5EPB68zkLDgYm3BdbIDE/q
9VaRU8ZkNWGOr2j4ftoN2LV5kZt49fztoFNW7HqNBPLlAb5nd2X4bPFMzDNiy7ms
4/4UX0y87FUYfOJjBGze9oq/R5m4hvk7vUdEoz/Ty3XOwDXx5LLOuBlgN5jDTmUl
XGVOUeDHgz/CoaYmG8rAP2oPv4kANniOulWnBT5dPM3DGXkM41Da3IO0d3wXkvu2
`protect END_PROTECTED
