`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
m49FiwfV/etSTBWuKqFnpMyIdtc2wUiwTeOoOTAy9uchcZk+5K/+3t+k3VSkv1/M
9snae68ctyT29Onlz2G++GsSmei0o2aGN6nYyOqoDJ1+1NFkAXouxCFbJSCcIa40
B7INki9dG2QlvyZZIXO55KcfUvHFW+pszdFQbELoMJzuN5OcVtlGbMkKDwA68x8v
RXvi0A1GiGuo6WoTS4nc3nWXBSUTLNKTwgWEVSDtghBw230mzU7CknV/Qe+Kuv1e
9Wmv2GqucfoXWz+gjQmbdrEIEfJQPxTc15tbGlVz9YY5EwJ+ZEmj1xuxP72aq/tD
piE0oKBuqrDSIehJxa4u0dE9SLjgMJEZUDFV3vG990q8X+6So+6Z7o5kuu8whAen
oyB6Wc30GhaCJ1LFTLj3oCYetzxP0EObKu4Zjaf4lJ2Yn38RUsYoMioOQNH1gr59
NiKpXfVVGO2t920VRRWkm3gv99/4U+obiG/QRhnMe5Y=
`protect END_PROTECTED
