`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
emy9jbVc+YXe1MqjDN7D6LGH2i97ghPP6KMKkkedMwMjW6H0rlAFC3IwhXHgW2KC
VSTxefZ99kZXTDoyWpqnWSYxObLZfCxZssgEFfDJex0NgxJL60KfIg9BdpYXGpjt
xz+ud0Yi7ZT+u2e5vCv+YgNab9xQeDlldu6YjwHUXwE7y+MRijHi19Mf8Pnf/XwG
syv3Fagb/8mAs2SNvsP7H0HCdd6SlnLgJlJU/4NVni1rCCf3GLB0QYXSPMLAIQ8c
GglliAZ1j6qY11U6LnW5gl/A1lA1CJnmHqW/ZOrvsZ/hbBDFiyO+P2o82fTiXTSu
gtHHa5HuFqkywM8yo/yTB9lYhPSjix1d+FwEjs9wsZqgRwn2BRlfbsQyjhe2PjFv
YV3ChkUpVIEpWZYCyRo9It+hxyGnZwoz9rRq4mI3jc2bHlxM5V7ZLbzsrFch2G7a
swvzB75x0NNKWGvERG60gvANV5zlOXCIWVuY9XaSc/i6RdAvPwDXgbTuQF2skADN
rbLmdkdWvQUO/w4pcddVI1yoGS8Kwf4jMdhU5t/amb4WHVVXlqISVze4agUsL6Jm
tEp7h6DXgobRuGiKjlzFe12w23baVHhU8gNlbH86VsCTpfr8B6coeye64DXg4nDu
OipjiWKgw+Jg5MDeNLXUzA==
`protect END_PROTECTED
