`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FwefupVlDuCw9nKmcgwBW/VsrZzdT1V/6TcP/AysGca3E1J8544vnm2lPYKeBsgc
mrdhYf7Ri0HV5/o0Yb5yKuadzOWh3xSz+SGJltZNbsEkT+1UcUuzOcWb3DpvEue0
E6LCGQMnZrPc5Db7vvqoHfxbyBQLdBnlVBvLZE1LLiNA+NtDGkPf9Oczg8OsyFo1
5gPKKUmKoRwlSxbCXrMDy5FIUA08outCfi67aCuJg+X6a96GitQFINYGuXrdQ59c
6ljUjCyvvmScYaA4+HR6w0KHcTyyd/yUuQM2+K5PmT5C0srsJ65Nz/dU7nR8zYYi
NcNdVcNaareKDn3BSLlA1oB0iCfZ0R07DJvcLw7TxnwjE7szhdsUlEQKxYoJrtuO
CDz3LSOVduxC8OawHAuGea1nQ/MNApuu3fQV6Fg+7k/o4VZd3RystXgy8Opcq6bh
8M9z7c0uAZT50D+AMg8Iih6Paj8/2lRD9sRYxcEXXylmcStCqbQdlbWlSDzWB9AY
O73qCSV3zYHygcQoeV6VTcGRKVxv9QHvAdyt2onYuZqiOuaH6MaaWrF6pgpzGjXz
gen97n9KxVmfGbOGenfWAZDRWyK+fSCEj794MQ6QRq0IwYu+b/bCoMvpg+VVQ1OT
mu4YWe95SmXX1xW6CA7Cng==
`protect END_PROTECTED
