`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tn4ALdz8kEQrabQZG4OLfrOFbtJmTnj+YBkNKggVs1jChW3hxagk41/A03LqBv1/
c5J24vJmfBMn14fbcJooHGVRTtr+VqSIv4vZ1pUge0fCua714VdfPWCQsKjJxRL1
fJOUsfEuR3TGMM4uJKEfugeps36nUbL4oqZZptBBEds8M5zfozKx3a9zRMPTZLed
Re22v+gD1U1VxMjGXY+SdsghQouRFZ+3QqbpD2rTrVX3aMXRyIx0HO7t0ypI/K/W
LasJTuWQLR6JqB5eZdcSRBeFAt+z6Dc3M4Scuvc7HgRu/d1YoN0ktks4Godg46hs
Xwik/S5NYFrB7u5I+cNQkVhH6jNR+SQ7nF6VRi+fOOzquWdMfFbtf6cE9JLKz7vp
hUdI4RhQ/3T9KCi05kUuYK8aWTrpU55Cy6dDOC45KsNCKI+P5ppEnUeDaXgGzmOT
9rz5a0+n5fE2fo8XW2ba/VSbRDCO97KNE6C0Y5JRgEA=
`protect END_PROTECTED
