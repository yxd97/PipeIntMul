`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vHXVGa64xGA5OH6vwftmay5yw3lbqvP8yxPn+2CveomDbQBsJ++fFf24q5NJCy6P
Pe+AiewW1UWbWgXCN1QUriSyFjYPSUEMWPk5u74jcb1xEPsqRXqfl9TzvpOVMACd
o1dxVklOUyo3Q5VX/C9o8HiM2o8fPEjqFarmEz1ALY0HnbPz+/99SozEQEjFHGKf
zE+gJb/2nbKwGVL4Z8qNZMSsOp0ZDOR3N7n/Q7+nqkEc0ElwiI0GE9ZoCXQIVaBo
jNoD2YRog+dZbx/Yo0i+hFhBlMQ6tgsgDHduFnbcjVLRUt8w0cMqeqQgDh+G3bUY
OdBPm2dBoIHTo+mlPDLvRcACnfesh5I2+lTSD8DNzJooEuFGQhXKZYsEiTyVzqpY
NtQG7q7Qm0Ha0wKu3Em9JMYOMhCWacf00BGQqHSglGT82vkqkJzQGZA2melNQZ+y
A68dS7pCF2C7N1cBtj3VSWl3hjwfWLFUda4sMjD+mB2DTlgEUDiPPKr3kFZuUOUU
ZF3CtSrU6PeyxTa6+iVKyQ==
`protect END_PROTECTED
