`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+GGsvzQ5ZF3/7K0+fp4w51kFdwAaFx3N9Hx44Tx87kr+Y29seCIdYYB/WE90Aq8
4yRlusAnvBj7mLJr9NZnAvzSW9sI2isGmWSwFqWOgy2k4bZtMgrkt26UP1N1MhyL
zTUeBLhyo3DpeKJflISh8zRUN/Ow40z891iqTSJf26OBQ/ssJreIomwusVLBGHAC
Z3nqRY73q3jGvF0LWc5gjzrc7uYRriuWsR+qXRtcvWV5fLIF2WoViJQadX9AJ3Hk
05Zk8KNWBCBrFwEzNs/bvqqHfqUr4C2ApJQ3tyTjfsz6G8RmJlHjQtgBBxsXBTG3
rgB2V6paZq0dWC6+1wrqh4CvH161GjPPKbmUeJh9zt5+1Tp9WBokAybSiIvHOxbd
fJ9hQRJmd+yZxVtsgjZLuA==
`protect END_PROTECTED
