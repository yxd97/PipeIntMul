`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KiFLK1P9pJeUtIzmj1SUnCKqyosRGhzMSVJYTB5LpwcXzNDLPtAboPqxGlMzi56Y
6PumV/+pm3B2Bxvsk/QO7UvViYhW9oyjG3X01C+O6dWIJmYZKu16b9WZR+AYQyIf
ycvendImE6raVGMxZJDcMQR4rt1Npa8n2X8hzgH23+DlkSOQIZyWocb2wfiHtmrZ
PJxsANf/DTpUPIIs9OtwemK4jPRxier4H6vM+7R3gLU55fMhgCZ16Yua+beze8Cs
VVYigBGr6nuYlvh5Q8Vj6jSTbnG0eogmO7KxfyZ4JXLcJziOzuhboIlTwBZ0wWi3
29CBfpR6AtpvrW6dGG6QU8681TnrXXeOiQI3cWjisr24baNsX3S5joWz+zL0Ws1l
2/Bs1k+gGOXgka/olbX+pdZw9y4cmuqfMJRkbA7jz1A=
`protect END_PROTECTED
