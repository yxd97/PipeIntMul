`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ED/3G84aG4gKyjJ/uwAJwqZ+FVPxRxz0E6ybqoHtAzguYBhGVgMS4xIszD59MIWP
o5g9vRGC24TponkfKZte8WuHYawflXhgJPpfoacnR8PQaWv5OxrgoXc0rZKK3D0S
/lpTXOjtuDxCphINQQmTl+GHOen6b7E676AO8sn8JfwNOtk9gn06tqM5mM15S36i
wGZyh7E6IJ+r54JtV3sTx52lqvFUq1V8T8gF9+YGEDlVowa7cIav29RWmgPtosoV
FAojMLPaL+MCrm5PpGGryA==
`protect END_PROTECTED
