`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HDaeF4oUFii1A637hh2Wgq6J1g8ZXd6WyBmTsuL6j1l8/j1jR004SzPYcJ003Rcf
/I2tdIJRVhfV64PQ9xWvI9i/zdJQSCJCYQjHxTjmiM751H/ZFvYC5sllkZOxy4f1
pX60H2jjHgle0zSNlht6QqPrhEnIVw/7Jms9Mk9slF8QSJswypXl4umQHeppBUfR
1Snq71i4Z8NPPo/5vQgquR7JCM+fcgjBLaqi7SAisDEMBh1MkQZF9ZqJck3/vqbm
iCF/vQ82YAls9qhJLpj0Wiz3l7RZRfx9ovBt2SvuJ8Fb6OLJHE/pj/j5jpcg/JxI
9aEG0C4Dw77BiWnnBDEm2WHXa+mNgSvZE9PSPB3hmKywUDcKmfjpjtPBpb9qkW54
FtQRYEoJ6TE7h+hSacRR2wvwBb3jcDZcgQfDbHpLC5esPdqEAoHmXtZ6QmESXhp9
Su0JHdBDTBf/4h5vadJGtA==
`protect END_PROTECTED
