`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JHkDFMeJt0cqrxmkmAMBUuQCt+Uuuq1AP+9u6PtDjdaM6JhO9HkZqE8fmTtuj7dX
GI5UJnUBdZPRIGch6N4DciHEWW/7AjGZFUe9Hyl/4uFq3BK1FkYv8swX0PS8xXuz
a8ku7Uma8t4q4/rlWEOR+q4UvHgfn7H8F/EWKINlcOwdT7iW8vouwt4a6r63mp+S
nKBVGHY/AU8VJE4ZJUTjabV7awmZS9tuc5sy0l9cg7TkYZvvuUgq/DXLtK7SCYuU
YhnlnSkNyteM9csCAcvq0dedGz9Fmpa4n1YIQU2VHdpWsjEljsJxvLv8T5y2FBGM
EwcpmtBPWveIVRlwR6Q9YdLgqzRIGWsX93zmPiOPBjgzFveJc9ZAO10XOVS9NVx3
86biZyfQdVSqEgEDL6SJHQQ24OOfcK9aWieNALsVvE6nGL4w/sfMBP58uwIS4/v0
FXPOsaa62N0g58CTy5SwahvxZO1wEUQ+hlzjtamJ+P/sOt7okGYFQtQx/7rUj9SS
Ik0kopdt7YCRPbpHMLK8Rim8uL0wVicNBgyN9sWh+CqOUdfzEoHdUvCcNVO6/+dE
TU1ZImvdvaEHtqpzR8oKz9ad9pZr9ilvvBJr7cp3aH8ETM8bd3Jzo0iF+PJ+eOTa
TqM2xFJZcaqJ5UHGBFln8Jh47Ym40vMBumNNxk8hdFCisFTAmuFO1/UCIdUe42Xp
HL9BzhnJGl8mZc/dqZISWY+W2PxJkP+kjJGdhnj/6XE5kj+ahzV7CSX1KYhdyFWb
thH4XmklSss40H7BPavhhTcErsHTakWRMcbnFmQuDZIg0X+5Zyxzt/c9ycMazU6e
i4xG/LurGwzu7YxtSjEnaemAExN6DmSyR7QjW77l/whjtQB3WxKyagqR2ytw4Nt6
1uMlMVjqhLWaUvT2Wnaw+6sIyg02IqTueqWZqxMytE2T7wB1PXsxxKGLCFQKPyD9
+KfsJWUPn9JnNay9pm5hPcdSvDQtq9lEMDMk/DAjwL2NXcJGJHCMVT3OB0Lrze3y
xNMCCbamS1sZa8Tznsk/ejRbECq/Jjpk9AhZHu6fIGujVnMhuqkeTHiKbBU/wl5f
7SEInLsKuui//VfAMrp5uHRn9WlkjVMR6b0VLIjA9jAK1oeSHj5pGbO/UyhMJY1k
9k0y1D7YLRL9wTiFRA51OEt+IUlZXCDJZc2SYRQ/P1W3FRP2AZYOJ7uIja4llFCs
sQi/00G+OY1xCRUCpbTDa1dqqxv/lF4JkaWHtIv5oLidU2zsIukw86pICyJkLRVu
Yd4VAgkur+2YW1FeB+hP9OCAP6dUjZK3GqFd4Gm1kwxvxVXaWUaqbNRo/Yd7fiZT
+If3/biSac1hPiTg7Y7O2+xsVdPabCC+QBnMht54JDuFJkOd9WVrJnRNwKQB9LIt
FNmycfDo7VxK/blfWhVjyADUjUQ70Ek2jYEIuts4BANDjI0OAyCWKEnDZ+wwdN5g
9LbGgbYSY9OQ9cOUveQZBoHPkXIs6PzbRcgjGl5W9y0bZs7nx25J6BVaz5uar48U
XhG50MoMvcW/zL5waVQ8uEGIhOKhF7I6kC8Wel1IhVFmZw1Nq9vA1kv5QB2j0WXo
8yJQAOnwOHNFGfL/YlPefgozC/kmhhYS7M0QrO5hf/EYD2dA77OTC4BOzLio/Y3C
1JBXKx9lVWu8jVqwxU0OCTDKrMu393lIxWwogbRXE24KZ2Jv9VWnHi6Hp5FVeyBN
wzMZcJF6yxF1dTR9+ohR78/ooTTLsZx81I3d/Dgpxffq/3HWEIJwk9rkxOfEWKud
j4V8lz8fe7xzl4jOqfSR+P2UaZa4DUOv3HID+stJ2X1nZB5dThP3I2gwR7eBEVOH
OKYg7Qn12vYa+/x4eiXOqqhJ9ElRsUDEUzr67lXKvV+y+/eXrZTXWVgr0A/e6wu7
JHRspK1qGJQUw42QYSwNPYtJiSI8eqAIohKkVQbnEaLwgd8NzsvAXhI6pB2On8je
c0Z65Yx3WwBQ0U1OqmEJLaT4/Udf5J/bgf8SjlDTavm97CuDFnsM0dNVLh35F0FQ
9i46IeUhk+rLH8Wt4cfdrT+C0KTJeljF+X7jefJup3oEFrIk3QWqMac0to2troUU
HOCjoHQ0jiAcHoVfHDJqujm7rlMCQq5ySqVra4tsL85IlBFKAW0JPmd0uLWimjzf
joVWRgtXtbP2o5mGNmLSBDZ6pZ0DU7SM4Lpxx7+ZtHU2Mjrcjr/W1urkw22B3/5i
ygrBjUWSGJ0riEOKjIxeYbsvxRXqYwUXid3OFBCvDPx7mLuNdPFxdhXBngH3gUtb
2GQHg9VF9tkOj2Nl+qXkM7xPJa1H6KEJMOHcaajzNvqqR1yosRINtMbVRf4Aw/nw
GUs8qginz6l6UjTY6nguTIFzoPdSmF537KBb9Pe34A23GO3RCGBi8p3OufZ3D3ML
6P1dotpX4gwXh0mjZrLMR/NERoCK+KBO6v5efSa8oSQo58xVxT+aBQyJwUrwWiIa
x7Bl1/H+DDMBtS/jR/3KJWHC3LQp6clBDwYDUvTjZ4/L4TwIki/peJZUF7Pvzx/E
XqHVwTD39qMxFr+1Ho0xT2PcGz6ZKu/9ZAi5DxyC1ujfIRP1N+wQfFBFDSITRkqk
9QRWVtbBM7etcwkkr/v1E6co5wUoGmNBiRlkQv+u39KhXJ21Sq6kcJDLrEI5kCtJ
wz7LyyoUWB8Brf0WPDi9OAkT1QC2vRN8Q0900195YH50ZAvbOX4/XmRZrJ16Ji8r
NN0Jr3cjkIX5SWKxL35I5QT75r0UUNy0NU49MKi1RjyfqFNMUjpa5Xq0vCYeVkHc
uowoK9vMdZRSUoA0JaAMzYFqvgBOZDqtrxOvF3MfwiwPB6g6s1/xLq2X0DUMUthV
Pj9Rlk7wtNBqiCjZDZMBPWlWaVvV/X1Kmiw7TJUg5Rz0uyUFksqrXAlKP+DDGh5L
88uzw5/omyRgMqqvJGCPMzDa7y63hGBpK/pvD5vCIvp83Z3zEX+ZwouUWiM4ooRc
+lp81tVcth+cxM9WOVbf/2pxqTtSXtCy6CNUSZruWI6BJ4y370bXeCcBAuTVtYpm
Z9GMovSP01sMGWhy9LTEgxt17rCptgq/EYIabbPPUOklpywPcx31wZBNvX6p70E5
pHlbC9Vm+0mXpRXJmlWY95eZA59HlDetn3ezHr2b+tuDkJJIbX3UlC0aZVvajOQB
HhfETQuQbjYnXjngowUD5lM5gwDW4+qw02OCWvdwtOpoNzdrB7iFoN9CNt78CHHa
ZV80L553MCiIOOo3ShhefKayxtIN9xpYITU6FdyrWuRaBBH5psuF2NplimKm0oE/
wCD3jyWth1uSjjGmHcHmfAjgwSpC69OXSsdmKventQ9CJv7cUT6d2x9CB51wbPR5
sOoIcQ/ULQchoNDFi1rRdyg/OzpW2jr4vwIMq4NdtWy9DmCGQCPD9s/eQiGW6gJg
ih0mfUPbk0ve/VRLuAB48XyMzuh/+Amc9msLqHE2YctgBSrFhJ77GNaM3kDco+/l
yneoY3dGuJwFkpWwwnu3Ah8zEnHwr/3YXWBxmfHFw6rL+O6eIDJJ2PcL/FtOnXq6
EQ7d94Wy0xm/sANcMB/gQoyyudnRLMeMVGlY4AWOMURRT88iaYR5oSw0yByx44FZ
CFY1Gi1WtNsCutn25SKpVEXDbS1Q3TByv8VAiYVdCWbLPcgn2KT6h/Z90JIpIAqt
GZU8Zzcgax70pY0EayBOXl8l9BNw3ahHi3q8n0nMwhxPOp91Uv2M7gVHCCdy7bKQ
AmRpqHrBTdH+BYsxZnvSkSp+HnvNwFLQrdTExkSQ/d3Gh6n7+g2u3qavQZVRHkir
J5IVWaHG0gGBof4mgg1Wf9ilsTF6X71NHxja1LR2uDdTfcPnJq1hidSQqftawS44
2II3JyM1XoEseX0Enu47hQ==
`protect END_PROTECTED
