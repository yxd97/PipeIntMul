`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eJVhZWVPWlcwzQgeErj7vO8ZKvo3DVZX0mWFpwr6e8Sc3N2eNkTPkU0XnoJcx+8n
KViB5lmotL+eyZcXGG/VDWAHdq68QRlKRGGFUCx8Da7HzOe6I2QOZHSKxc1lFyga
QEJ67vvs+iWLxJRHTLHlC0xnjQr7Cg42xD5c+FyMQ1mD/WOlFYeSelP95b/zNmuE
y8DcgVrHEkaOcnvrDeEfXr9eg+T6eMyK6j7//MDbC952SbxA2sdWEqkZWEAvExtd
2Q8iwqjtzWaWhdNUgyayhGhblE6lznRCfVGA+c+hyz5ZGcLka5bcRmUzzMpYJ6nt
1N2jKnS54O5cFL5lfxFqEi7DJGSEKEzANDFrN/q0xNLCJgvYCJL/7dk4/LsfVWgw
Ek9qmYVQzRNH77ML9qjJP7TT93tSkht7jgwiiZMcWuScedqGV5lq1l7yg9EXlUSR
zti4y0FM/ZNiObegp3zkMbKWPy7UEBv9LW+ualB/FcmxEnyalUXu0yn2Qn2ed5s1
ox0FqkNtMz27MAEgzeQAJpRDiJj5XxIz4ovZ1MhS/8WXRv9RZyBwb4hRywHZrMqe
VOPl4oGL6cVJp8wWkeBERL6B8svDWDlvcTQfkNhX/z3wJKgCoBhew58R+euMyzgK
dtt8mgHcM0jxuaZg0l9IepirKkLk0Rnr6mbGzPdbSas=
`protect END_PROTECTED
