`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HhuKPabokVGilhmoqH7x5ABIAb/ZAGCo6wJNv6OQZ30WX8vzSKNRaq4yNpE2iW9n
V1qM67PiU5K7FrqPueDCQvtq0arITbfpJkRrLAJrqlGqoCgvpBG//cYYfvCvxcn/
GarPdpW7Xh4XTQjEFU2hAed9nwOqaCMEVp1S2OJQ4DoGdV+ifFF5OpevyN12/WbM
u85vcadaD22PMBuiWIWSECsMvDTkU8VYdZ8qTCFW3SV5XBCLOqBQXXY6ZjrvHr0T
lGGzkHVHwUcwUWvq/8qYY0tem7+BRtYaZ50EehZDirHXXkefh/hnH9iWYtnQLULG
AbvMXQhvotIpOMyZadw0oURz6j1TBvvZ5K1KSeOQXOMtwwWFpC8uQ7Pbdu78uAkU
LXd1e86HeAvZ+sEZCiaqDoI+zcO8HbOzwY2/nITHDc0=
`protect END_PROTECTED
