`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d7UJOGeNH7kpBMB2v/9j07Jy5HuwLKe2EKFQcvtv9ZbxGvXQGoxU71cXUSKbvKZC
3A4szJfbqA42qX4hLbQ7JKYtvgkeRX0Q22ZdFDpslBir2u9OJ0rzyv+lhjuiW180
wIg3QcATK5EqOMZWoAnX5DJQ18J6o9DOgvhllUKLALejQlXytg46I8U66kHN+ADX
yjPcvf1RPlkQroAmhAIYCUXLNX6rAOhzSl+o0tEuMelxpk00mGvn8Pv5B8kuqXkT
DgtfcVEG26n/ncF3iQSzva1r9sZJ95nqRZPAW5M3BPxtG47jlJRtYKnJSCJzMO8z
8wVsUmP3TjoqWlyS5LQE1flvuCkgD9Z7OWPVVPFFaLntidFoxGfxx8j2R1FMpVdI
1RVcwv1BbI9rhN+SyZXW7oILy6pchR+vbuJZDg2hpc2RNwZ/vsi57+6O9PX75lJF
1BW7b3AsIxAKerruMTkMMkwKR/BFjNZfGITEIDMHHpqbAmH4rwPoN2xKW/tmxPeg
is3dASb3I+pTvyDV89pyfFPkHeL5oa9hDnUw5MFQOMaPH2MgWDnk7GD2MUFaOsKw
4KK9W9dr8795MY/JtCjImmRgSw2iUeC7rznPB409+gY1TRN6E3co0UZugYXBlPaL
Qqc/pNx18L1whEm6KycfFVAuFshwdCxHEwmFjEYAqUUP7wcQBCbUie5NmtJhxrCH
pd2gvGN6mG55oMmz9g39ZsrARNT9P5CW0FAuKFudo/9c73fz63bJwA08019fwj6V
QHvjJnNhCho33uh3HAuiy+ic2HrLDpVa/xrz8mefvaAk8IfXFd651i6xMJmQJHFD
NbfBZF02un7vFShMq7eXFqP+1uQnyP1kW8UeZiA6Cy9d48tVt07GmEEG4z2ZQHmT
JknUfEXpSkF+hZgLg6KV2gv1tOOdFHTT6RSV81bJmNV8vNIJPlgvH1LC/4gfukY9
2F/zxeVwJGDEWMRhaTL34cMGByy9ok/QCkMxqLbQxyLSWAVOEW7AVZEz48c8Ac4o
fS6NvtT023nfJeLV6BH7HbgM30hjjIYLo0qjw777OlCX3I3lNuxCPOMRDdbJVLED
LvRjTf+F7GCNe8BGAJITc7WxHfUJjQXAsX0DK0EEGFPoMkf6yNESzeZ+QeHv7BbV
YnjvExQ/UsWO6kqaLr0T42PT0sKsFcjEgeihvBdVcNzozcIW/rwMLCPDyd5zJp1V
jiok1Xw5otOBk3Q/7o23MEnuzSd7hG06b+JhJBWeWnmRDJb/4PpKr9aodtd9QDXK
`protect END_PROTECTED
