`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B4oMVb2KHuC4KzDcyELHicNTt8OUW7+bjsuAz5QRZxMh9lMuQh8mtAJIOPGGiKzu
NtGyj/ImQ/WuHQ8ev4amhclWzVkY7YMZvW/mNjG3E4Y/G04/tTAuRauqGCFBf0Wh
YzDfL/mGgqX9jotOiy1wjBu7UxGqXQyPdWCxYBwq6wmhBmLJaeISAOYcbmsbS25K
wnaFJ8Fi5pB7/VpAor50KwbqQ5948pkC0C5517qEkLKMwgguDMsxic3tcB1KzzLC
Tyt8Sj7YlzCeKHMRxohR3Ii/WrRWtBbuSY76Wy521hg492fWryshZUxXmskqaQIY
soYj5NCXHV9oPRbvURH1LouijeItoD2MQrIFyCXadFspX+SLMMdCR92Md4c/EnZD
aLWPpa6qxOHV/KY4ynusIi5hixBHMQML/imIookMh28ECkaJkzyBHTC4jQB16aVa
ayTbzF4LYxR9Y4avjj9sGuw8/ljy2y2MdVyqWwFjWCBoEgYYZiUUNFC0UsiL7EM6
Sx/fp+FbI1cjj+99QHbbx+Amq3vjemM5xblbdFy+Py275HPUnBBEVy2MHesZWHvQ
vP6jC0SAgLe6CvLpHCay0Q==
`protect END_PROTECTED
