`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DoHW/zj0PgEs1US52Z3udf2w2ZyfoBh2/kwQYSNGumkKk2AwoF2RLfGFPR8oNWQs
JcjIgLPtHQzDIbsVzygEAhUuA2Puj3au4gu9s/Xu49PRnXIGmleZjnqr0GxLypbF
dLoeT3xHpPou7dAnIAIEwwX7jYbKTJ5dGDawiWKLTEhuiFZ9I7BpVToysXzFDzob
zYuIhaeFJyqQ6cGm2hDdsd9HW5mR0YQG10S+sBYwGdkFydQDqw85YvRUKRqGk338
rmVCUNPLYVVVzb6vcYyCb+vIh0ZgyAEbn5IMvRXWUyBtuuc8Q+N6ex33JEnV9anQ
jQSqc8wmNr/TEVzZGYH7XRZZjzhYs/92J9l5Q4risdlc3MJIWo92DlpHx2C9zLXC
D3EZB0lU8zFbRmpQ8eAfNAFQ5wdvpf9d5TYDNDf9xy6eiFMGh7xDwSket8wFpniN
+KbklADPr34DUGky/BDE8aclYz3dCW1uItKZDrm+bae2VT7B/JhBKkqN48WGgdUo
2mm9ZX+WD9BxMluDpDZzhg1xfQsvRY8GMqf0OzYZoRg6cny0rK//PAWcLdriFnrK
98jM9FI56KxMN1GKaUvZKdhR9Gs4gTFOuofaoszLeXFWao5kVVboiBF4qsoQRnHR
bpajGcGB72KPVzryporwZupQAS7moNvzLkqkFra0J5vFsS+eE72SscUPDHfu6LH8
WtECdLTXJIYFN8chjD6GUC1xis+NJKsNttzSj8i59lBYexz7uy8U1GRKRCVyQZ40
IM9kzroWfP/PRVwcDufKhacgWkRx8a7kBYYf4AaXn6lOJvqV0zTdXYK/lZQAC///
n8Imez5Qw+ZMnj4soXKAbFkzxStkH6m12ixEBABSG3TcAbGT7alO/NuK1zz2TQaR
aiAeXOforod6phJ2otQsiT9u/ZU7KxU5Al5rKOr/4r9n2Fo9wfCKihBbU1v7d/6Y
`protect END_PROTECTED
