`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqtJvl22WjVkl1oe9CHF18EB7c+RtPkHljhYiHUQvXUkbx3oZxrGTYX2T7gq79vp
okc23CnJLovhz7hXVGXmh0KCfcnVWWUu+GGeZQwtaNIh25eqgbU8dKYltiO/5a2u
/FSraWnCACD3FdzTnmDiEhCPtrQ6L5tmICIPCIARq960TW/oEHrV7lzNmkrGMyem
I3Ee8R48E4VlY8R74lN7yXh4QjdXPFw8mZU6J6kr7Q6fIrZ5zNrGlF2NHn/5G7dV
0NAe5lMh/b00VMvmCA4euDqTnPmDyaNTI0u4oJp2ovIp3K1lEtRbke2t0ooop/Lz
/X4TvTBCcGx1Y0Z5tUdmSShGJDckbBZOBbwq2J/IHYI=
`protect END_PROTECTED
