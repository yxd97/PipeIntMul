`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yGhM52yLChTnJZjhtbQlZbVWa5AsqdGmDZfP9CPsKDlomF9BdzYDbl7HDO2NjJY/
rwSHHfprlTAE2zhSKKLyTEulrNdo9otZQTTbh3pC1YrNWMKODr/lyL1TgK+sVnID
f/TlGVRdBU/C+1irbFp0xFkWFsyJuRBjIsq6OivX6tZTcvw9BGjN0ToH68NmyLOr
3lrZHEGvL4X8HmJeZs3wOnBxyrpfoS4lrYggfhjVJ43klocAB39cR4L18NoCP3wf
cKIn26hYwz/694WVDmP7yr345h5poYQoI378wqUHcGbPs/3jNTPVhl8hQsjgncUT
SulV++QcxwpS946B4Cpa58DPmeRHCZT2IJ1G0JUPqDbDd1wUd9XRfKxGGvhQ88zc
8bgUry0WG+UKDTWNYEn95j6FwR0HJFoJ7x+eGDfPmvU5N5aJh868EK4henPDtBct
c5ww9pP3CraN6cqkfoQILlyT1UHmJ2140REDU1gx2epq96Nwlx8ytCyI24b2R12h
SQ1JBA8fn4jPdHszgH0fuWQ4EXJnkANA1GNrJp5971X96Vn30x5Y65YZScp7a1M1
O9ZVfDb93HFbm/fE5XacKooRjBc4S7RZH27ugNj9WB1bgRilqh482DBZwH5o7Wo5
ESKyeBbQ+Q2bf+NcynSq0WNq7STfaaA2H94LOoszpPI=
`protect END_PROTECTED
