`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fo+HMlWBX9Jm2s3oOwU04kch0+g6ZHmQTkp29/8KWtSy0WSx5y+UoGvmjTpPl5Q7
faCcqvGsl5cNIsFwpzIz1yhEE8Mb3B3r4EgkCeeSTX7r8L5fRIpV9rsN6L+s1nO0
0CWOtdYdklRZ3HYCRX36IXeawmOpwXqParVBKnb9kZJeX66IhO/b/uAO7C5M7eHf
8bKcjPgrtlEqTb1uYDaWJlq2Bw9O1VU3YPvPwFE/T//GQq4XBoQxzRjerEMZaW4y
9ZIQcflgnkbVzBwW1jlkO4f01PTIJIht4EG/QfOf1lY=
`protect END_PROTECTED
