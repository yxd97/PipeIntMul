`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+xq29M+caxY9yWCx7HJsVGsXf3jouiHEekQP9zPlwYcWWfOYsSZwYc0vKNi0jSd
meX9MrV9FJMHnig3oi+UDCO3t/g4IOF+bKfa2WSG3mEcEUdYHkKLGAXpeRquyfxA
8tUnQ/TeX/4ydEf3F27doBtqegXaJguVfKbi+EkvDUDBSxkI1LJ1uaxR3fpU4s5R
inT62tREMNiXm+5VA/mBA2Ym9fyybfCJ0HfFVNZAOcOA1JpY9BUTK1Y2g1U+jLgQ
B+XSlUbjHbNDycvXf+uNGH7SIU0MoHHRuHiKFHTOVidbEXX++8jq3Cg4KJSQFA/J
MDc02Tzxz+YPdaDpCexEkt63c0YBFRQJE7iuCQpWK5ZPSEWxDq9Xo5fmV7w2QA2s
1xARJ0V6DFhDIUZ8f+YTPIRiHFoFbQHp5drcHkYir/zcnFLO4kJNzBtkiFMuySx0
y6uOHgl2iMwy6OmJIxZGjQ==
`protect END_PROTECTED
