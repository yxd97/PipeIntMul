`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jzj3+SDGSJMqOR4iaSUVBuqnNiDzx696NrrwRr/KmmdgalUsM+nKnVJgTYVNcTiN
ViCRVKEz81A3sH6MhAWRVybnttBPDNGUckibNNO+3ID2hB/ObETFuQlIAtPa27Yu
ggpW4RCkmgMqWnBRdIgbhRFLD9BzTfU44p7nEpTW0FriBxbX1JjfjCyivKaeDVjC
STlhT+OivIoCInnyLixzAAQK8Ckam0/PJDbLU28lH/PFrQt/o9I3ii8EksWDXt6U
trjznYKgpf5b2v5U9DwKsgi2vxSA6MUf6IWRR7y4qLryuJjihgE3x44m5uEJJa0x
Df5sgntkNx8NKG3pJEaiRIfmFyQvfjDLcYXMmqnZThaR1jzZJ9qR764Ds5XuEp3z
MLgIgfzei2bZ2DlVOfn7a/OET6AkdgxZB6c1DkPG73n1yaDYpicWUp4Xne4QHzbE
DjTqLI0KEbqFI8S+TlS38Rij7nEk+626Q9l/kztCncy7AyhjZ37sap6X9F3uJlqL
FILey22rIpgViKpXOKKPAvNxc2yLV4HvHaGrxc54LEj3lwC9ZoM/mPGYgqmHNZxE
xwZ0DrLsYybHc2/FcS9jPvvncTwZwbfQLESwXq6ZRVUE1+VBQIQCvPmpDrbMLwTO
qTpkcWlXTCq4ewz+xDHYTszE0JL7MXfCOjPm4sxNfLTZrubErCUzV+9S8MUOXD8U
UwWPeFP0R46hUzEFGDopnGuxoKb6Pjy0tDwdfyImIGIRdEpvj7ub9/94jv2vKJhM
Qu9WbpnF7f8hiq5btFzI0a79qxUTjnbpWHqdfeX2XTKUKASHme9RJeaCMqqrjRSJ
8I32OjtIkeb4Ur6MSsnZLAliBEvmDiT0a+sgEgIM91HpSIh5g/lrujLWmrT4mr2p
clvFDbcWh5cYx55pNlNJJC+uWLA5cbLAA3/MuiwOiXJZtLFlGsJQGCieAuMGi9o6
qDs/XwGw+KbbwA09fEa/6UXUA9wO/G8OdLWuMCaUb1QT4Rdjwiy716vE4U4nILiD
7Wv3fh8nYzZ/EzZvJwHEC1lR3/waAohM20sbdlKUtDQfaTKbCsHTAQZWYsWbh8zh
ROs2hJlK0oDFIARaPLqOlnSeGDP2UtFWwrObZIMBqqJ4jMaOWfWt6KjcuLMkPOmC
1p5Mk9PaDZ/bZGKMp9dt77D5ynLVW16xWAB+dylolCoz3+p499etk71kwKeul/AN
YMoY4hwQgjMMFlF2OE2o83WbJonm4FwRpnckIlmXCivarZWjQQCBmKaXiN1WWEMh
7ErLprpt9Bt8hWuYDsXlpgWvLSqrLWQZYs40CNY+VH3kWU1JrwRnuN3KRL6ztZ7B
WaYyAajqPFDCtpga9rgh0hRi30FCECoJdUpslI3DAimjJHYvbir+X25/sTx+5eXc
+D7KtylfDJqdf5IGyDc7/sKuFc9R5NcnLKAEKLRXGcQCrc4HkQarkrNxp0L6bvV+
DoLPGsR79p/IDo1Ox9hBzg7bkN2qXrirlyhIMvWSPGwunPwaVEOaALDJxdJ7+MPj
eDtxoJuxVJR0h0pYdV2IVeCrdsvOVcrcK/6kLNQLXOOHiqQVB0hibKXlE79aO8LM
2d2P4Rh12lSTKZ0Vd9ECfOq8QvzDs/9wmka0Z1FyI4y0aQTBK40rDukuJfGIkzzg
hrG+bF02N6pvBMi6iqLNBZZ//Egr8YblwNfX+gJvydME3p0ahYotOoaOT3WRfjhd
t98B/A/BnJux/7NiLyQmEfaYq3Ldq8PxlDfdkS+hIdt1lJuHZYGjJ34BHEX6Ms3/
mZTrIPvymGuMHKkxk9h42aMLLkfDBu/aVuM/Re1BktFAnlas3H0RozeQ/WaGS0pl
IUdYm+XSkN7jGqjTVc2+GnPtiIqZD5cp+mzgpPB1/2rn0RLpFNkXyxiRzu34v2kC
KTrEtU99UbTTa0u5a6/1O6C0zJQh5ZwNTxXaSnHDx1MZuObTbKARmbTrRnjPuPwA
h5KhwnBb245sN8aY6Sgwx5P3Diya8mh5Uc3sW2kuug9647P2TbcXXPYv8MQs1c+1
UwwDpFbJ8Bc7bf1z/8Lx8PrqZEJ1TvXdTKVy+ZNb/ZnB1ugLd4FVuviAW5h3Nckz
SJuv/CplkO5M9CNXQdvNpn7x8gyfRc823h4nzmCa03/rmbFMt+mIZcArQUiKTomS
ikjuA5UDGiGCK1GCQWrhSPZiXRmc88Fn9E3hUhMJkERV87B67AziW2fL6d6DrtzN
aW2U3a5ApRqv2a764mmrKduYim9GTpWz61P1zYnNPqCYDSflNAZsiJZZy6/nnhc7
kKx2lOYPFbP/KMkr6kFcTwXXdWgyB/m9t7OKKfahO2yDQUN4bUUKQlx/pfR1VUeu
LmFimZAo3kCuK97AtCWtt6++tLrZup25V6YmnsKajhBu6LA1Hfi3TgvovO43GzQd
8djNiHpS/f30Af/HeK7KnlDeSf2EMDSqajuI0zsXKXcflgq+LJkxYbi8wcrRKbuH
QYK926y+guyCC0NRLhuhFuybaE6dA7TPwwlFHW3GcbsCAQRKi92Qpl8TE+vMOTxE
toKiHSp7uXnxiX+5/ej43pAnm3ANL6LVm6eewkTLgJE2fVg1qmStMHRALrQv/y/C
WhueP4tdami/vZfgZN1FjuppL6b+/2hpURbvA4b6Dv6RFenV8szUWSVC8HOYg+py
C583xPmJRqIY2OA0IvBd96PO6ZyhF+nWnbfrqIZS+G5thst/G5KG7wyHK8kUQzc/
cAocaHQdQgP5cY3wKjfzNEGjDrNfSegl6AbOz/XH09HcxzlZ84OIpnzFQP4+32yy
7ZcqmbUAJZf2o/8FR7tpx9YnrjxJYpZJ4GbfpnXwHmx1M22B8W0TWJpaowyg6cKS
WE/qSjheCWrxIYpwPmvK+nJ7MXoNd4EMsmU/5lnMiWL0FQD9LVJJMOYsdwjggejJ
sQHXasiKVW3phAYw6VmIB807QlvIvl8rN/F+XHI8E7NiTK+25zN95pDHYRM5YOZX
e63/49nZBupGzWu2PJ/ui7P+uKxSExTxdn6bKbZ/G84Ajd9NNQHdeY3Whe3ei+KM
`protect END_PROTECTED
