`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3X/qq2D8ShH25NbK5lhulZ8dxg6htCmdHzCPxvAshuJdHK//pGEBgFFCuWbwY9GM
pAk9zPMXqs4p/KTDKPbjeEBy8dxcLAqvOTb1G3Oj7pjUsAU10wFDB0lliGepsvbp
n2mzWlR77ykrHl4sbH4vAtxmeE4NLGtvsR72v0k4Tsw+MCI6zVvdsHMKwkcSHJSH
aANG5ppqBp54fOYni/TQaqdFUHp5RfvS74FHA7psyoeE2v8ZzuC3pqITAjdDziAK
0UgDkYCEtDG25N+i1L/4BIPWFZqxLpejNGb1BNDNkfDKvgvuMoYfJp4P4Ncw2tWZ
ZRnDAJvfgi6Gl2QNCPlk5KSmSsNxPrefhzKULu3YYz7U4VWZT0umMbaeLbr6Ih8O
7rHHvBFNOxruTkG8vzhAr6TgjBIUn2C9q5Xt9eCG25GDHL5suP/1WZ8hJ8XUlG3S
K1zRCpfaD4reVY3xJVyvHfR8BsAUri7eTfktTvyJxbi7TeKlD5Z+Jqe2kH3zW9rd
dKMQA5GBvinZclXkG4IWI1xQ04ejyVjFQcrB+Yk85TU=
`protect END_PROTECTED
