`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bD2Knj0f3tdzYVEPu5i1BTrcIkE/xUsWQ4XUKoa18brXv6uT0Wkh6DgaTVQxgLPS
Ghpfre11aPNaxY1URQmcvgdPjLPd7j5DHPmL+fKha9IEOrAAs3YDE+OI3iIuojNA
pUTlX6wtffbiXNUfLmHxqFgYAK/HypPAYD3NUrl93F52rUf6S5lvUsAmqjqMpLxd
Ohkm/zxt4FhaaAay7b8MbKHJIebH3OkUjmoxyxNTihDeKCIPfOPXD8v1QHwscwu/
0O/1ya+eySnjtx07s3cZjSmIehYb5eQRhkleV62PirUI7Qe8AbgYdNKy75K9FQc6
FMBkOQKAIxpFeM6v+o+EEXpOJea6mLw9mVq/ZNxo3f5D4vh+KPJl4AnpIVoY5cvC
QmRDsDvBjeiyG1dE0z9vINxQevpRxxcDJchR+jjk/Eok4muV4HJ0x/N+YiJ2oIku
7GQZKvNOlok8FrHJsxuO/3mXd8VFhgOtQR1Mar+7RP2V7Klk4uXF9mDGbqvZOgRA
KvQ7VfgTv/mxIklmD1kHseMOZOO6lImVSJ65IAD3ynec9i0ZwC7sRN1c+9LrR0Gn
qReiDDNifW0n905+DfGTe/5CgXAR1Ye5HudcpND2Rwn+hPHtqqYThBp+g3ZisgTK
uIVmiCtimyPGoKQ7g93yVB9vPTFRjJDaifT+HL9e4BSUW8WL9ofc5pD6kI3BCIpN
TUw+/mJTvaUosF9RYBVBiLFa3E3oL8hFo2Q/1ZHs2yr42xzVNiHemD5gpgBYncrI
eCLtP9RZZEPcKZsf/yGLlaNJSz4ZfzzZU+14fqwJbVYvicSS/IAX4DuVzJWT+Bdp
ZtkLHZYSKG0wi9ovU+qeEDnPnfJUoVwc4Wo4QsPMwyJyC37lWkua7s5naFT9dVlg
gpZeNpBY3lOCXbCC1upsxX/k/3C62FEYsbjj1iLqSKb7JGvGOy586Qig1VXx+2b8
QME7z+De1auhIfYKdgElkaFyhIJz7oyvNEAVFztoOELcLAn5eflsGlXeKQ+xs2ih
oCJHtwE5q1CgqvwP7ukWf4nsZf2fI1FUKnKrTiSaLm3cLTLGxdfPxomikN0DAdmt
2Wy11YoWgQS6Bj61pJRHEGqX9jfUeD4lYiBqyXAfiRBWLKZnaO2SEVSdLqQVOryd
ipn4dA21qr9HBvsb66AbZ33sCjdTyNd0Sq9R5pKoXEUp4xIoaNPXCNSD0cFH/IiL
PK4NSRNwTEcge4gWg6F5oGpsmaYOrYFTSq4pMI7080kLIkn5QOTU/C6/Aoe8wu47
F9I6EpLAdnDvglHIujeFnypSlsYUGmY4FplDPuDMRGqKc09JQuHTvIZbAvktulT9
tOpe9f+As/Zo6fYA6KUk+ir045+MzMT4rfsNcBmTRR7ArRiVLdQpowy8gLI+FVZF
d+iqYleBJgQEhdP9DgYSUBiscpmjC1UYXmsAgqRpjKpa6ieObdS6FoUcHcYjkenA
hCDpc6rrhyxLjnFFLzBNl1PTEiRRSLvvslZVLklfRbOW8+yT6xl+GuMc+ZxJo2gQ
waCkinTq0L48rx2Hz8RdX+TlkrnCk+aOADO6TNWy+3YSrAfvY02Jvy4I08Rwjhix
GQB4GE3yDnsIeImVBGpB1KWfzB/Fc4Wk4/CP6S3FQhNlOAYqhYC068YMhM4h/4+v
A5IM/srcwDoiafS8MLOhrkHmE5MdQ7N37M2SsMBeUX1GF3rlXmVVAsZ6/iNUHMRq
bTIy8/cO91IOh/6kuS552ImwjgO7QjaWMWKZaM5AAgvGs1088j1kjMWWFrK749Qs
2mpP/hoohRkScJRi4sVlImS5txW21+d5Z4lWCJCwbc6eq9kpcjXZcSBG+HN50ark
2HAXvMqoTVtwfcwjhlY/iX9THkII1vRi37HkgeMc2BPRuf9Qzfneyefrqu5QH7Iz
raoABSgCHDIB9BQa+N7k4wIek2VYu5z/TiPrcopvNnfjb+a/nhUuXvhPWehmP8Nu
3sSeXmEt9pfWg/tzv9xNiGILJnjgtQMhuVLZ1VhSoNIWr1bYHleHolSgbrpHNJV4
Nb3IgjnrEGyi0vr25M4EDl1y0qgzX+axJ0ptgRpnGK0rcZ2wI8UBe6YekcQHKbiY
GQt97H/LVb1ia7g5xXDMy+q+oH6MNO/XG9L75GBuGfP8SohKmmQbHAIWnT4V+00M
Trqv63H3+hBI9gGlkN+sWVhEGY2S/jbE8CSwssmuCXYKGfUpQvaphs6FjPD1NhCe
eh+UaiQEdWomrvzf/5NkDgYWzD3+H8iWwUU7czxIsucwOJjIrmVVKaPjetvjnCR/
ko62WZSQxwF0UBEQTXY54fS2axo9H1VzJYdCZcyc6/k5tYAx0byh+xewtNFbAnKz
7nf1pkLCE9Cr8NNUL/tPqXzZ3blTUwR6AZu2RhbEQvHB2pOwwnDGvazxDXBlpNGP
/7PVu7BUtqorAoNdu8gUyV4Hm7ERw4icVquTSlDnR8F944LQfTT4aopJPi8KKWvy
Prw2mbq+gW9mEcS0WAxvlYp3WbVztJ12ccD7J3a9WlRpDhnnp7lKn4IeAJHtuI4O
ISyyGy5b8lRM9uOnC/phq8Ek3GPBa004FJcvCRkS04vKkN6MP+hOd9pOb7Pwqn9v
SNoHT1CBjjJ3piMZVK5yvBZ58kpk3yq9qhntB2TplBsS8GCsj3XOUmPz4Wdjata2
UjYvStNtNdIzZvqQtbKq6IZP6wo/xwH+4cXhj4zErlU8Mo0wba8rGu5eB9FUJseD
4MlpYv0YH3dH1oiQ5+UB3GvyNpDJAev7ysPW5PsLaHoqIiVhhq01nXEXu7akuFBV
qz1xBWthzfovqjCFJPjmKpfuTQ57Gua1rVyYnCwOSfbfOzBFoYIx/fog0OkvFKNM
TBg+GoNjoikzbplngH2kYGsptxsFMv1HVQUVCJb7zvGdXYTGWXXluAIFV5I2QyQN
kPJv4ia8qpyTuvJFtuh+A+h9q7siNikUM0TSY1w0K3iYoYyYE4cSXAD+7lmiabNW
5fWi/Ez+NaqM6J19z3H9RPHBYWE4TSXF5vokjGyn39/Tt4QKzIMnuu+inj4htRGC
Hz/BKYpeBAMBQ8aRvePnsgpUkZeypXBYVsvhFPTnwdOCNP5A+4+jfYlzpjLZnfEY
5q5oKs/LI677lX2IxhagwM6InYnT31zJEFptHqzgG7HZxIM9pst5Hvc1OAerGvvl
mbB2nCJGWqyO3qAX+G+vfBkEQSjPFBtVtFzF/nPuQB+k2zHFjiydr8nOa1Id9bH5
VYf/mu7dzlryOzjONFHG3Ime2Fgu4q+M9MJNtb91YX9exsJ4NFLNORsGRfjIluF2
rEWBiHSePO+XKwEAhhCPIxxJgbxgnEXtwO0G9crHNzq3+RWqq0lV1h+3w4eSJVKi
RwXE2qzobcZLh2Zw6KI9XqWaRHJWAyTcHkM/CTBD/edtYTya9wm9NWPa3AgtTsZu
jEhHcnD58t9Mj5C3Ccj1cG20KgeZxD3+QM1jO8J1047O4SWM0HrWTfjOSx9YMCYT
WRtb3qX4QQQm2WiOajJDn1N94aSKeGVC6uPfTfVCRdoh/LJI5G5+xhAn2Y3sWFwn
XBHBqv0rtpGzm1/2rhSq8215FtqnALFfxQ3Bw2+SUc5TxFZtn0sCi/1GIUiYdnps
qLp6aeM5K+d/K+WFbldNO+tq6lYTezo46j8bNhGqPI7xWTBsPWbbW73iBsCQ8Jco
jcOynkYYDVolBNz1Zv2/CYQb1tTlrqLwI2s6GQLkN7KsBEabAfbJLuHKy3YzBQfo
UVkHd2tB3btroD6ojF5UREA3SQawzQdiVdlMRwaUDymnzycLWjR2DokKKk31rUAt
ukWnCQhMTbIGFhxa3ERTHhOj1mN4W2y1KF+6SLlM7iOafstmt7Amn/LixxQ8uMfo
gU7bMAxTQajO0PB6ExJUBADxVeza45JFg/PO+wnTPqugtaLZ+P4ycbHWvcHX4A4n
bcsLvBTmcPAUQBl1CZRVqDHVjmKdmyox7RDnIbOD/yIOozmfbUSCCYczzM3Kdl/L
Up1DU1Zxrm4sHjUbcQ4oPXNc3D3mRY84GKs4nHwgVDGOEAteurqSNnSkpwzHXvTh
XzDnFEpCu5TiLeSMFuQF6PLjcufo78ghwiBt+arICYOAwatATzpIBAuFJqWEP2gz
y4dFcg0jBpCLSVbRqH83IaPMF1xFSAD2RO21gK/FK7PKkMzBm0DaAVOTErUP8lYA
JdaCkO5yCCzAzucV4BkwvDPobMlCcAaEGsPuxjGuvrscJQiJxDtuJhDP5qtxccoX
fLnO/8dc15XkR1EYXAv9KQKuGfiYCThya+iW0nZG2kHqQs914HHCgTDKGmBp5uJn
bhqEdvHdU/NS1i02NRlKeinJwEQaiOv6uQlCJsXaYeM+vf7JhBnJdFqAHBxNzdM5
rnZaZU+KStTzHJw4MpbWOSCNh+Wkvoa2jdjkGoJaRRO2A6eE4c/NJP26OKArZMdr
M6U6BKsblGyBl/WUjKlgr/8nmUKNmY/MCaOBxtUigCZjEzVMxuyKrQz8ypo9sI38
qbaCQu/QgF6pacUdKc3oPEREY66aTPZHm4MFOQlc4wxKBEJ5+I4Zks9vqnVf6fuY
zM/bfRrEFgZ6pFqX9kx5gsW65gL5tjYJpxZGJJK+3a85PGpyl5eSSW3iirEwgbAe
bSmNQbhP9OL9Y/rm+o79Gg19kSiwBVWh50a4aQfD1DsJgG1KMBO7yi3WuT7YoD0A
V13/Wo2vRGZTnhDByq+4F9dKq/CO0odhoPmWkA02It+c36h7dzg7CM504riFvD1P
qSOvKz4FN1uzPF10vkwuVDHLTyovoWBmtKZ8M7zjmjk1TdhsZPfLx15+n+C0JCC2
jDaF1Hs2GmI9/rX/1seug3uWlMfQ0CzLx36CtY6N40iIEGeIqm0VuWVRRCm5EMjG
ILqAD+TmjXsXR9FTA+P+GisqRMnKczT/lw0wBDb1w0K4gCtR/ZTGHl5pGj8jtlpK
itfsENp8HVHXjg9WnhxoxqBH+VGz9rf0SK1xeSOXwn1TRroHcCMbPLWeqBn72HVy
YIccvYkRvQVgR/oKAuZR4qElu2Qr3BFdv4DL1JuwsgGbfTuD1ZiU1PRxZfcFReUg
HzBg0kcaN8FK0gKmY5LSPsEbh5P+KEZVsRKbPiR3EVt2FqjerT3BKGds5LUgjmfQ
RvDOt1/k4PnWW78NeKwMP4LyLb7tMx2YVbDDt3EhugLjjUR667+M52xJP8tndyQQ
zwSf+YKc52NpK8AAYjokELwie/4cd3XJcePmbmsD5AIithQiYEKg2WvOlTUZLouv
aRvXGL/11qWwdTZCVhC7xnOsUWPsGzNmtCeKaefuiI4NBWGfXqZr9U6GEKkk21uR
CwCJnYFfCDDdTX0kUHjvuB9dOFIrlYlZRhgazwfEF0WuJuXlv5Hv/GPUEmF6/Fnp
j+574fc8UgGG88nqfp35k5aPiEHgi6Gwb+nGAvNwdGNljY18IRbDESzG21TmkZOk
spKQbq8B0VgjGQADJo9omO2zeoZbg9vZU71GJh8pbDzAft6BH4+hF1M8Te36lAQt
4Q1G4ar6kbilHK9UK++rV31lGei4HrKzKyIfjMg27nhkNa+nNTfPmp+H+ehLut8h
2KKf2nOahEdQug+hli/FPpBRinZhYnmVXOctDuo1eZ9PYOEZ6fjDyK7USLhVZbM+
YmwZDTPZ+DFpZ8Np5mmz+GwhbuxUWCf86kilypkxsSQJLtPpX/YS97xbyLK8V2aS
8SMs1ofYyeBQNuURHonm6wp5CJsR+3fl7mxHnyf16/6weQJnaoFHh6GK3u0rsJJZ
sNfyAsPqAAZ8ukTqrGpQOp1zC/x/JR9fBihAYazgoRWrJsJ8ImkS7CUfovKkmHSJ
p6GqFB+0d3VM9NdNy3nb9DA2ZPWWFsl69XOisX2fZ330EfJms2c+p1TBBCFIeGsp
ajqrsrIysegX9gFcaZdMo6rRuIa57uYA8ieIYLE8BWxLzznfDfGxYly4MD/dbH6l
EPKZ1r+PTjaQFlVNR99NJUUqTPvNUsMoRUaaewq8WqgefzV4zERFgimv7esLkSB5
thdy1w9oZag/1AS5Q/k4vkU3tAzTKighP7xPzM3xUNQaFAUUDqkwaP0mMQvE7BrX
G8vU3VqjyXmSYKQYhbr4Avtp/d630aCJUa/O92saDM6Dcc38JWnR7nD4J6o/SW5K
7D0G3Tzim7lpMEqSAOucltV/BIsTqnEmkz7jRZXDK3fmCu3l0EXjGM+YjWcTOC2D
9+ORzerhEelK9qfaCJ4SIY/X5f7A9ANsM/3/mMOepFt13UMCLS1Ur8uli8lD4ewJ
t172vIgIcVBMIU/tnROnhI9RX7zwxwBJjnopyOTMah9kksR8AgJF52dW6QSH6BCN
bUx/8UGmkF31clyX+IYBWLi85W+Quy2JngcaW5+JfmiVCSZUU6p8nwRzNoGBT4aw
jjqKLaJ+VZSkyo7vmIQtqWEtm1XKngS9jMQnRXB6womqHNTmaxB8AGorS/Eonwpy
iyQYtiQZ+84vez2rxCAOwMrFnajgJQ9onGBd45WSU/WbG5bSslLP+k/rGE5ShXDR
E4taRi9qCcGTcwhN85VUqXYVAds8eZPa9hIbVJ2FCp3rsgq8zDoMQklgB4yHCOVy
MxxwnXoLiXIqsSyVC258WB3EcezW2U8xAs/9iovD/KU3X5iNzh5PG2R575VXPRr8
VKorbxHPpaEzn2xNCZnk1BIiwYcLnkN2RfwyqA1t3vZ2tMRJ8deq8AnzP7k2XZ0u
tG8p0KOluTIHieXnrmKOSB9zw6bECdw5q0ILRD3kJl0tpkWWE09ZyA3LThzoF/f5
teyNB/qIIpraFH3kyJJFKUO42cqk7AJT6R5/AAvd/Jrh1cTJCr/+NhAq1BG2dbUC
8f1UYH/B7LBFYakVLV/j8T4ZhdBRJXWD3jwumROFlAMmae28mQPOwJGN6Ml0D6RY
YZGpDiYr3DBg5ecGzrzeGAYMuorNxapCu6PFoTFHI4HwKGfiAGSaX1l5FTy4ONjb
eMwK7u+9QQ97+aZgRY4Wsn/IoqIMSh5XChCEfmila04wYRFnffO5ybjgDm8SLkY3
r66yMH3weiGaFpKYruJYuOQIS204mWsRnjXCu4SK0dQH+3BcXdgPMi2sybMNkODw
opFl90D9ZqiB6UB/ROVEATxqKMEqesRv9HBjwlkPfQSJjXcprFO6XxjvtAKwlw+W
xpwdMtswxxNswrBpHNQoNYvZySkzYdhr4u+vDoZ5qKPHRUihstrOBnXR4ZPiazd7
jfUFQvj2OK78ngV6xol2pnf76TCMCd8QarEXQtjFk4X+NIzkQxmkHSCyfATqkIxu
uhnLlm23sbcc29OkbCaeZKOR846qbkRdRyYbNnRebrszJ6O+37TCY879AKj+/vD5
K8i/PDc6OB9bG+yZUV3tRUAH4dapOEjobImQV00/5ET6j2vnQ7zwnFGnf/NI/yky
NaC05qxU/pNSuD5SxNMJURQd8Na0bIDCAN56ZNazdZwzUI2ieC6C54y+W3lEsb9f
gPlOsnQue11p5UEd8iUsMtZiIIWOtjQoM9bavt7/FDuF2KThE52Cs/17Xa5ep5ya
Cl3D778h/yEJ93gmNazWmmxPytZOcDOjEYojDWgNRH1BRbkv35mYMrkJUczih7Wn
MjI6Fu1cV2RLPsvLhiZjl4+fNfAgtvvWRYyDx85Vd02AefvvPCDgzcJhDq/Ki8UY
XdoWNfsECsTbE9+ALszNhB9/gpt8zf+VcntXtMFvlUgKFRCoglqS6dqhAZAO3qh5
vvAchDchGh+DIrJ+6mrtX0DEAn20JfM7IArdp69umKAFda9CWdkgGl/2jAd/SjVw
Cha8hRJ0iuRovHPHwrXQowQg4BzQgqFY3dQxft6BxyiwJsmDGYJRP3YCP88QZamp
JZ6SL3shZ0EDQ4a2UWoXXHsflJApNeFzInBOfJMq3aqhCIvPTddwcPB5gJ6P0CSr
hIrA2k/lTbJJIMF8V60zttW/i7El/tQujh7R3V9reKMzrFx66Q03fhau98pxnB/o
MTlcuZn2l5iQDNh3wgbf4JkgwroNKzA0PFB8qFy0M4ASPnkRH0ymMQfO54vPG7Wz
JUNM55ze0ncBO+CHLLH/VYQZPsWO9Hyc4O0A+ps+Hm6E0bmC43cav9yR03Rv23u4
B1PF6Dhu9CaN6J+65NCLG9Uic2Rz8pbjKxJCkKkziCI3/mnzLsR9esyW04sQyVCX
ZvLky5jRyyWgHkOG6SGoqos6wXBiCFnuWGyaRxUZJeMyVXCZJ+Uifj2LQ1KEWuCi
t/IpxhKxH+z+/6b35hsOLScEAd95furnismVbtdd/jMdwgYrrPKcQByQzUsPCbUE
E0KFizeNHjjbky7kijciiXkR1bkiPyl4mv1bxdCFUbHM2z1xiU2dwssXAdofPGhH
y6r8nk6I5nYPU994+q+yxubZwuxjNobHA/cMqCeWmi1dCl4UYxxXgX3xnE3gMDxa
NbWUrta2hfw1o/lcfCT2kpbg0Vs4Ml6rrU3ZHleaom82PfvyYcYRF850xrir/k0m
XUXnBB572ZNDcUmiVGdJA6nx2XfQunpAMWh11AA3R43s0ZwwZLouinvBVKREbjnv
DlQbi6wIYfWeHshB5PkxBtTZOnQ3OOr4LShakuSZqRxeOyPg6UtBmELu1ccmpAOF
QIowBBknEfe1SXk4JHjDCbtnLja/0KEfrRV/CxSL81g66AhorOaTxnK95rkIRmkB
cDvUCeFjJS8nKSSfG+dcmUg22KgL+z/GQDiNUHZ+6vrrA5qqUxisVU1YEGUtsrn1
3TTSK9pUGjOG1V8sQGQI4BHV+levBvGLv/ZQ8fJacqCZSQrkoj4WX/wqXFPB+jcQ
LqovNqUdMGwDy2D8y2ryIewyG2uifHbRtpmSEeAo4FjsFAyZJsloKm4kMNvupPzT
chg9R6/RfIfba2YNpiuPO3Rpw7BcX+mznmU5pA0IW0wZDlJ3NnHbQzH2lax+r8Am
8IhzYBjiFgDQyld3fUpAW/A4AU+oKPRbVzU891R4B+9UjSC5fFpg+CeGhRe+1XT0
5eGdNsGKfS/KzqDVk+zfKwOpTkQ/fhvFmG3fILanUrvvoLhk9x0OweEch+uV/Oo8
hqr8uTIrazblzRiS7f8TZvetvAekj7/R6iLfVYOkIA0URzD7YmFNes5lPlxOnoT5
fRFKQF1ICcACDsSFZi4UmHgPLVM75awDOulEk+8JJvDQGm+ipI/rrmkGJvYToq02
IM6bY6r/rJ8SFqkFkrkW1lixKtS/fnBwW4y57oeQs5bDlNi2Dodrgf0iHeoV9+Of
+s56Y2epiDhvSDTLgAss5Dmh2Yc8gaJUqrTIJFmy5NxwSaGC8n+49/2FPewaJmkL
ZQ6McIoqcpRePwG4SlyQlx7vd7le38JoUq4Cpd7YoIoRFj33hJKHY7SwmpXaC6hD
lZJ6b4aD577Ufn9aUtsueBOTP3R7aG/uBxyEDmN9Wq3CAWkW8ZbPUm4wvlmIZOop
Oo9syymQx9aONRPIIqX6vQtuySqL/TCmYY2622mkNcS9MDU/UBgthTOjKSp3tzbS
1xBXT9mQKVsxD5KzhXrODEKcaPI8/lxdMuG1HPB7OjuWNDCnAawdj6f3oFxSAQhY
2wwxV0K0xDu8f4ikOD2ZE+7nmUKWbZbDxFNs3gzwo8ID45bleXe7rkMkBp6Pk5bQ
xeqVCMRyseJdOh/8qgbzYrlpx9KIlS0QdmNhaJJs2k599POd0qV4nL1uwkG4nfoO
17BWYYEzA6YqEbi3YSkDjUvdaP6mga/y/Yuw68cir/WwescukouzBCXroMSk9XgC
s6n3oJXEDMatPZyH+Xjx50H+lA++C7zQ9+jGICyQeJ3KIninRedpl9EoqlF4/4Jk
4Lejy9YKmx/313WtVkczOxV7aaWUFZRF2ZoVR3PnxWTntamDuuhQJiEPaACrj2vF
oACBSGkjCvCBgNWV8rm+Cd684ye+Dymklll1rpNvteFXN1mO/FWfsgwsdHURgSZ2
OhN4knVguOEC74BXvr6VSot6xMxfZDNvpeQaRdiwLLojOjJIucdS7tmZ4inBut4W
Q6XasqPJtrSNEAJpA5YGCSY9/yvNuzDhM6Aq83Z+kTlwuEuhqK5CsBjCVX9W9yQh
Td+iAooz2fTc8FphO2ca7QoZ+6iX+5pdiTX3DPCaH8G/Io+3OoXS/tIQ9ut7zdSL
vtKZbwsqzMUgnS9O7HugzCUEEK3oZ3/GGM2E+X8fgBwuvb/n32IrRCQ/VoZc7qD4
of9deU3wuwr1YdmzyBthiom7YGo1dADVxayCiCgInAty6phKiR6bKOy/YJ8MbMm5
ziydklSL2YB7wChBBJQ/AcYl33oRx5Nel80yCFMXwjKt4Pn6K2AQKL5wlzDBzRhr
adZ6rOmZavMPNeBrEW2LJcD5t5Ck6ldND6z6maMNCesWhs/9gkwnnwtx4PJZHf2J
Q1OuatFjea9yTe9JIOE9wUm4CUkgHTmsA1j+Wlm6K4x3FkMYPDuYKVUuPzCgkid0
K6kz9AwH5Z0HDPWbY3bi5ZPfE9DcpDnwCY/Wj6pFuhTcs/jX4Va1rdIuc96zmEUd
ZzCCy7Q1Q51aBeJftcwDXmk33o6Sc9ijbPTomEVYmfoJUrt97s0Ot7IMHdT2/ZVY
09Ak88BINdGJpVCL3lH1GL7ppetpNNj2/2CF6QLM9Rueo9o5imaINa5tL2mGMxX6
fuULGFl6HcBcEiYaVRXpM++Z81tNEv+HnmojFv2ehd+jdCsZzh68j3owkRhqViwP
IPGYJOGAeCcGkGXeyKSwXLn31gXfsb30wIQLHFPYzkGEchWID/K/VJbQF9mjx35J
xJJI9qXd9j1NsKrLnKJdvT/5qavPOZbijkb7OUFKcgNDHa+NIOgN8+o04tRMiZMJ
7HzfDnVoa/hDpBAZJy7J2F9ftAnaE/mukDeQvcVoTDwjhKUcEDGZFOm26FMtMQNA
0+q4IB2LsoIazhvgB9in3koL7iNx2L/p6gD3Q5EA3ZU8Vy+KrEl0Nk9Xl4HhP5TC
dbnjQPVsq5VRfsaxqxhb07lPt/ZhJETrJ+8MfDQfpqQBhX8XJrzpWxc2eg4BbzMI
IRUPNlCrJyT5lJ4BpTCwJPJGp5Yqj4cYNdshf/8ck2c+I5U7xmRqkIQ8VSUXm9Oc
kOAGyoxJeAn3jDRK13iclB+8Fyr0XEs+lI4MmoZFtEH8HGFaevJkWy1pJmKB1Gmz
11uJdUwZUn07L3ixEGYEodAbkCdqIibPc/ptLlxImdWNZmcZGAMq4/qMAVHtqbjH
Pg2IbK9gBT6XLhx7WhlNE+dHtBf9E2ySnVZ08+iI/vI84iRoDaixMqvYqvDuakIm
fAf3twa7OSNXwwEhrDHxxMkMb1HKEFvZh2jtWdhVNCAbW7GgSWLROXRxBH5g3Ywp
YLjo0HGogACjchBGyuPP+UW6kHL13QePSrRGtB8wyZ2Bd1l2nOxXPxY/djMpmKHA
c3Nfs8QGy5JbH4fBx61bEt97b4HqWZE1B0mFVnFO6Kuu/BWERdyYaJ2PThk2GQej
/WlACeJmBdxh7ggXeGBvo6UrtSsuaHsiBv/GlHSl8ZgaNXmcJVcCGPLiAFlFgx2h
2suwxu+23z1zTvllW2tihuWaCTc4MYHuBDAmbH27MIb4FAIyKuSchskQBsKv/Oi+
lWyBCNm+Jfp+PLAqmEakYybmpW2LP2zTugwKTHnOfXBp1QXI8vBp7tXBXIEP+x7k
3wuwELqTM5yxApvNUbZ1O5XLvLeYk7UsIpRWN9k8rgyUA6XuVrkCXoYW0nSH6NVm
cd4nSF6FSL5QDAnxuabSMjJbcYd0btDCjWr391Ub18T/LBikWnq830UyIk0x0y55
k1SzFxIW6TNfkgzioaB8jXYSwz/LykjE9pLTSXLNLDgC5GI+rWVHQWHQT8SRb0gc
0cC+cdCb4z4orTTqSdKX1s8HahZjRjJeamLdTCkTUVpVl8RUxMYww7aok77uQhfv
fo5/CviYMWlKrMV64A4QVsmmbj2Oe7p9ZKWk7qNDtiTgcmvraMTpapF2fExpUa2E
jwhoR3ou2S6M1gvWPvrFDVh+onSSRqf51ogSApV5F3q5km5Bb7/mjhk71yrYrl9L
PKk89+SZ21zKblzWwXsX1RZvrBwrP2tY4vc6PtOgd1PtTJDiANDNitzFX45GOr3/
pKUMk9+gAFkEp+csf/cnQfKFiGIEbdKiuKAWVB5Nd10x0CVQMLUstjhi8r5A5ofN
wt9OyWbn2GbvejilDtvxbW6h1+zjj5FHk3RKnm0Sz2B7Dr6CQ7uz5UvafuZwZmON
jbLZPKDI9MUzWcTL3IVb6c2YY80dFKyy7tKMWpqkN6/ygbo1W8IwBclZWrCQG+lm
BchgQZl7lcuc0236u4hhavQCNnLgp7OxzA4lpweiIWWukN/jzToCTmrLQv5B4eMg
gjFsaog0zl8GUJO+cSGDmhwu+8QksyywxnBw8qHVnVS6lkycrJEtPeAkYYeXJU3z
ZUwY9EuD585pC/ajCNkC1cKfJzMcanHfHuRzy5dCK0H6PsYuVo24x+q4Z9KYPLsd
s83HJTMyzFmk8K0ctzE975rQKP2z8eMtbqTeqjz69ZpMnBLL9R+NtobEOzr1p9q+
poHr0JdicUjFYaDxkn5cQscN46Kr//7GxDtpZ22p1A3nnsc8feJWOhInZkUR/L9k
PF4/HPzzCfOCVQ5pgbTkWx2ZR3QBGj6w+640t4wo8QbRoBY2VXfRgSdxJyOothKk
BQEPaUeEyHZx/GxWxVq8bMpmz+48/0fDRgeuqU64DT++iea9TZIQcFbgHRbVNc0V
XSaA5VJ8SfaooRSTIwhtfQVzosFP2cpPmTK0+aL6MybmdzlfkYB/Kp2lbwE7CRNf
6geI6YReBCEYq0xLlyhrNzHIePrattZG4wFjWGokzsfgMcXSQjsR4HTLawdlHzGa
SwsvCV/cN2UDZLZURB5Nv1ME4yyMuVVOyf6DWBf314z3AWXKK8dXW/1hEHoa2u7k
t7K/QAkDDD23E58kw9FkskniSSEWZJqnlXl5YGg2i6IGJhd4DMyhC81MCIEAvG+O
YeHK6Vpv3n044+ugfgfXztzqnCtAmgOa7sTRFhjlQ18C9TJFay5Htv2Tm9oS4ulZ
ZXInbqMHxb6ZojL9qc2YEAgMPTVjxqBVP1vcDB/Gt5ZicJ3j4sas/xbk9BwntQpK
FIxmSgmUsEx1YSohqqaO73RU/03Edei0ZQ7zC2jRZqxeGy19Wfw2np8Dc+2C+j8f
1VNGvhgO3DkDMx1zVipTKDIKXrKKcAOjNtKDYxg2H8U9ECAeb5VBMKVpeUHsp1Jt
4ymrXc9jp2HVujYZFMbSJ2wMtqN21txrOXL0IO9weM3Am9fwCo6QoW2BuRX84QO+
KbIm0hcoHxJCh0snhX/EbQxh3ovB7veyX7YxxjIwzMaRRW4QzqUP9fsshhjT7fz+
CdX8Kbo1/5hncm1VpBixviX9erL3jXiPa3Tb2SbmCbvQsk3zWIVPcS9RTsSwPj5u
pMY5mlmCK3sXl7EdbQcHDUiM7hgH4KSpZ7ijKRpYN+ag8mFu86bHFuLf6diyvQGQ
HwjUhwbP2ygIlyJ08DFr/O34XnZdmb5hKyQ4emdMX4u+Kgz3Rs1w4Ijmwz3pRniv
0LC6inBs+wzcoBfkV1jWyzUdsnPJyWV8c/GLFCPGAJk9o0lyMp5msw7PX1dTl0uV
joZ7YDt3RtBqnW73obVPMXj2Sr7th386kCsenn2+/0846amauTg3Ju2Qhdz6Nws6
b9vbaz8o2aVLx9i1HAMd7TGKjA19k73174+AsEYTypZRzEpyZVQC0TA9mclmEpJC
AKix0/zsu3I3MUvlzjRndv9OkXT3m7AsS8Gec5scACLIVNrRKI1uR/oH90bjfaNo
FJpqekJc2bzDroqcwT5c13NH8YdZSByf9WQOJN+WFLDYB6lX5VawEdXuFpg06n0g
XWk2Oy84EMt9jDuSbtfT3twaoXDqBF8jlhZH1WLuZ1wk65uAjepc3LfitT/3PyWu
DKJ21GHotQMXnaNIzVfGjRW1ET6yFIfEFzdrx69KpaHPUUICF4/Q58qQCjRJbYOf
lem6kQ3fz3H6CAn2+MJFzwZvdBayaxl3PfV2AMyCGpqiTxG4olLODBo/ksAsBq7t
VfUvHX5xn5+HONALXUQctbN3zsd18S0KSV1BiuIyWbHawL/eViXnA1GZZylaKlr5
/brm4hzFXg2pSzXWL5LNVV1UHlcwrU1FxRDajGh8ZXWogx5vAmkO+vqhYQBKGdVG
E9cxgQPG9DfNP4Ta9cwv02lMth5NgNs9QIjqxJdYropelSSLRupZVRT406Obq+rl
dB5jpDhK0i2w9+tmwRXDgEocC9dZGnRovMgQTsEMLXqWlotIb8atK8dGG6dzioYV
dWmataCYG9zlT6T3pfMj136TBI12LecHdpcwRZtV10IfFZcxagv2uDBFykeigXsG
BYR3L9arP8REVmeWrOfsnfJieWa1oN3EV8reldS3hjCf2RmvaLKdO6grlG9OAw6Q
i1nI4o/zHFaS8+DQLH/tR8hpKCmBPb2iGUSOzi3lOtzaLAZt1Wa8X+Rnc0041Lyi
t0G3Td/MQmpmzafigewcTKGUb5PmabB5b8pIE8aQaU8HnaCoogJd/CGHKQUy8xOK
9m1TzikafuogtmnnZgafwmzwtsw+mmj7ZCu7N/lGpJ5Qd73cIdYOEMztdeJcxbIC
f4hq+NECIy/hj4Mbzs1TxAdgyxFya3kiF71OjDZY07RiuTmoc+xy7BtRnMl8Bth2
nGRpdriJyaBug2nAr62H4b+JQyDyLg6EpXqSPqygKPfvbnckSc0M4pAUuVlHlGgS
H5ZNqw6+qSbD3+NXDW3RHfTFK/wE+5JSuw/on6iNmS3FZ/73fraKXq6gebzyMR/4
d++H21IlKu8dev5ZhMdDvYdl6VtfjU39apjfkWOBVgHbFzBsBUQ4yJybwMSTnfkA
UXUO2YUP58sKJWWJ2EqlhjzneYARmxsJdGFqxWfwi/3BU+0HwD0NpoyjZPfJ0xWm
g5hWSzecJvxoc+gmabC+omS8PjlNdyrMp8VeHx8QLVbn5SUypFDV3EQcB9urq/D0
bDXIJIVFn1tnTfH2tYR9MoEJp2JBWrEGNZeWMf669unASPNbOF2ZijhBvnRAnozS
tHNzH0NjUHsg38qE6qzb7LUW+4x+y5BfiPAqwpT6zh9poqvtlk+6svse4dH6GIuo
RS7hzuTnzpKzVzgPeiO0iPkn9A0C6VNlynu5liu6+0PjVtciDw4m6WVJVxsYd2nQ
9PhB926xMFhedF0fpFyuTo+yWrLyt7GcpIn2AHAXvd++pd+TM61NG94jw4rE5iYv
2tMMwyVhacaUhFxQs2M5Uas4XZF2MmxVyyaVn3bSIPAliS1Zwhlo0xKb0n/eqrVI
aqtfWULEGwNGtxpXAv+OIp+1oXO9gSZQDRyEAM37hocrTKEWaxbQl/EShUfab1FS
PQpT8+WuqUg5b6YdACKT9hbrzgrs+yF6PiSTWTQv5kBlAMnv7DOofj13QPaOHBoY
Dq6IzlFon+8lOUzNlR4Elfcs3wjiP4QzRb3505PADMIJx+QVXXcj/JPhKvmzin4D
lQqRv9BqAFSJa5dNSkLwp/QSn5kHeJi84YPQonN9y7So/hro+q2Wf08+swzdHEGo
qZp5n5zdpQml0m+s1mfi3mHS3cpFhvi123vQ0xSfTbvqF5xjW0YHIXN8wFEBZSCa
JF2dIqhvHsoxlBKaMwTYi7ICVXF19sl0EajPXEXfEuUd1WcZtPKDxQxwjT7y3GCP
FQe7WID57SRonlba++2TMoAfghnfrMsh4bWlNJzad2eNyHpqP6iFrRGYPMYGNLdf
a0Z/BW48FSW6CoIPpZ2jG4JO7aXR1l0xVrSrXzX8DEWbSiw5FcAFoJ8uZtRZP+WX
nVcNFkXMCq3/sIkryhNMJMkSkOEW5tlstWjo2TCwyqQOL18JYf78houEml+u9Mhj
fp5npMci8cY09n151+r/0iZ99/oEZ2KNDddGZNcq/0whnTQno284s4PryEDN6pJL
4L7Qz3PCD4oCkV6DHtSmH3oH5LDweZ2UwJlpWsfG4kgP3orl+nECXXfJwyqO3IIK
1OzBscLubZndBwlSJEbVXdOgGcyhfSp50NYSQ6/O8D3RgBDoCla3TB9l9vQncmqj
sF5uaKljnrMJBpr/wqLYq9uPMgOEDDdoVNcZcpfzJCwO2fDTA8uSALOMcyaduNSg
GgT1kEWbZDXWzRdNlickCjiu1AKwAeG5C7Kg5unODD5X8IMWXMMpCdp9ou8zxq4h
BIOevO7ATR/NxosBxPXDsR83WdugSo2H8EbD685o3eq64mOx7gK3Vv1uBAZMfwPL
8U/MdRee3UYv0JJeku7jpCD8NStzzFgKljXtr0Y5T0i+2BQwrEehkkVoFSLSenHV
nTfHg71CDGztj6Ufjgv3UT+VUMYgoLPmzGQT2W6xSAgNq58z11fSBHBffc5FjW/W
ytOOa8CMkdZMPt29TU3otfSKhcd5Z3jJcwl0+pddEhMflLPBAugrAkKzbqFOJHm4
iigWEeQqYd2mEpnS+fLvTal90AdOJG75EReBJC1m0jIGu0j0ke0j4hV5DbRyVH4k
n0qShRqIhvJHjQ5as6kO6FUSMWx2qtXsL9+FSaIkMmwqdui2lk4Q1VP+KyNvJrbw
OwQYhQexFbQPUW1Byc5q3LFs+l/AIcNUViAcuE0lj/77j/YeP8oTn3wcapUNODav
A2qEc+zCUEHM+WagUHOLlxKq1VtSzz57tDx4PJue5WnMPDLPME7PVR+nyubqGtX6
iEcKsTAKQj3oSZtg5FUZBxNKaFfeOm7UhGNlHQ9PfBpElIxxpXiMzbLocCoHcom7
YYBq6VAm9mUJwO1QE62HDLJUPBP42SnE7hp18Um/6MpzxRvbMYmlOderBlBkN4vK
NyT5LKfJWNAW0ImTYNeM6eW1uIjxk28TjEqbcLeem4Xje8KBIVOhLFKF9XvTQ8Vg
taYwnWjSMp4t9XHMiQZ2Xy4Ez4f3esC0pl42j1wjV/rz6z36qrOvQ3hVVqyWvbhi
ygTi3vP7sBVgLtl7M6eRpz1mKBSt3eNywxWT6Hu2PPUoze0FhXonlMxc6n5EKr06
nndvCqBUecAiV/dAAU0mfRcGuEr76+VWK4tmItaGCiuGNdmnbQiBgTHzGKvWYb8Z
VhLQSYRRGg4FruWOVC2kepTOP6Z9ZN3BX0mzbI/hoZPxv6UgaHyvfxSSMxEMvIzS
aZQNBmV0HvsPNhGbB1QV1R24s/5AtKngY8RS2+HSoTbMDigatRL7nNUmWCP4Rid/
jm6GSkLC/oXPU/QfefIH5n73VEsAxn/YiLsCgAqYfQVhGlwm9be4+kxUS2JyqOrc
ZdOb9AS1UQX/9G3n9eRniZPtVrf1WCd0WOKoUCQZtZPL/BJs/Zun1HKoI87naRkP
QByrF4scASTNN71yvVP2931cCKx8OKCRuom0aALMUlFXR+QqQ73/0tSEOB5s3jJm
3G9rxNhIDzH4gomaPHNYrK1HphEjMoOe20k42YdjhbGUOMPHat91wy5SP2SXdJbX
HUgNqIkeo7VcbYnW0eubynYLei1ADYTTlnFvMbO5a300ittYXSKfER7GtlV+OesT
K+Yn9KBJeTm68ZRc70Pf3wVXYhEyv87EMHT5pEK0hc72stJF9bxkFP2/fq7TCDBc
kqmByYi0oyuw0J3cgGlZVSHeDfPoA8COUqF5XcEwldHt8Y62Y7YO+w251ZAubvHA
DVBzHyurSwiiQQng9PVigM0WP2cZRSCLyNEyEV244wRRfnWOpS0J4WePNrMPiQCS
G9t1mn1e7alPAH1HWN3mmJP4/fG+raiTMUhF7lIfP4SmNKz3WzXPlaec90y662Ul
QBFHYhUFAan0ClK6hMKe+2oi9L/ffju3qke947AKuQqWm8zqn3fxeYBkEAuLQUT0
igTL0Wpxavl4bu3Vh66K6NqIxkTUlcFkfyzsbEVAMz/tSi42qKsSFzBcvSK/EcmL
++AZbS5pmFpXYrapyeMBn/12dJjsoGYn6h/rkga1RMhSszz+Eg0ZSW+Vq4U6LHxY
IwHDxJ4oR2L7g3DGBjrbMtulCgSO2WE9HrqOrUK6v/kYRCef7Emc0xTLKeita4rR
bFEF1KyflTLT16F8Zw8LZqF7MwwgOGip+zCZIQatRjkXRU6JkQtftQRr9dpg0xdf
2KkCDcBlEJKmzqFmRdYySUMd5TqJSVNF+Y3Hznm86JVr+sLeh99+YUltMVw+1HMn
kbn5HnXxUhdXLDpjhXYDEanMo38SnEHe8SgI5w+QC4knB5Mc5H6gPvCIZrj+f8qT
ymX3TVY2fqeiTaVi7PlMmjXoP07+thqg2T1HWTExqnT+6GveDod2+TQi/kM+l4mV
+7/mEmreDfz+SvCs9FUVwrILPcC812yVNRTz6MVerUWidNTqVxpStDpB0pOYqx6N
a+bN2UmEuZ0+QkETtgZmAi29eIvbJhNc4oa9EeTKq3ytzaUVq4QFZ2crk7PyxJzj
Mc/IgT0Kopugk8dPRflZfrZg+fJfNkV60YaFenHFu2em2CDlUhk3fQVE1whQMZQk
LYL6YdHlvljYz4GpxpnVp1HUycgokh/qUARlOEDlvLKDY6qLuYXW4FXt/rxEJz7r
A8rYYfedUkGWC3NPnaSQ3wnaRMIOrElEzKudHOVHxotxNKRbFbUMwBQAhwJlokJE
4Gt1HJeoGqyLc2uuYJEaPUW49iymHBG5s/xxq48OXvOFBAYWklq8y3h79IQQ3PKo
yh0zXy1FEjunHFbfIJDkGPehGyO+OSQ9LDIWxHyYuSctMEnANEFpGXTEydp5Vlyy
QwLTq5njbhUIQKowM1FHHoil3MFp43LUX2g+1OULZbY/bbfVZDU3vCiXSzF22bZX
kSKg9DiZOFG5WFBiT3x48vbKElgnYMWjlTjtRxBQoCqj9Nd1nq0xi9ztt4PYn8mz
ryo3ctyw7908he0ahg1GcpJ6ds4as67o9KC5L/ECY6Nr/iLhS7DEmPeplXVANF5q
Dk+bB10HvlbcWk9c/OSIRO3GvHMiTbzEnHRdKGAydJOZDWYo9paXZ2NViw/uBj9f
BI6B7IDenXUb37Jp24eTdgc4NHs0gjqoMm/2cixUcDE6NFBEHd8LahwFPNX379He
3KgLRHLVY9FlirZQkO9XMaAJtgkBqUTeAkWdkF5iMByXs/TdJVgGIvnF857UG+r2
TYccNNyhA/IcKnHl0KovgFKsMIt1b/sr99mi+71O243KewJBpvxD45mmSpsAjoTB
mNbDMS4EFq0C61Lq5Ju7hPjp5VZ23txfnpU3dybCRxb3daz6k8lonWTyZJcPmkeI
Ckh/xzv+nLx6cmqYzMVAqEzgniYU8CynfkAAGic2i7k/SggQnKHhgj4sDsKRSlCh
sVuYgJY5UAxAoVL47Ev7qyN36WZ4WX/GWBPy+rn/UQSGJR0eQfLexMU9OH23I6v/
0ACp9PntesNaUxqjOauMExoDac1n5UlTUBtZ+Tfk3vG9b1qPE84BwG55IuE/IOrT
esYwsrpnDSgUGbeqmm6xk0B9OJxP+dFMNRluYXhftwu++0C0nwkxQPYSznMvaFtf
WghGrObzN8c9zB7GPkrkHrubA+hhV0+ruA2dVkAoT3rcgrMT9HSM7YtVo16T6FUW
osAY/ges+Q810eiGn9bj0LjLfs0k5SMnjzC+GEl2rXVGcr1zSj+gfzziMX5/hSWh
o00QRvcT+ifGCFcKmBsxVbI5oQfiLPpxrlWXbZYck8RSc5rAy8ONRaFl8xtjaZyL
IcBjb9gkk/C8DDOmMuxljo9XgqPYQmIYVNN0uFxYDvDangEoIZxnLgS7QMnxdXmc
eYFT406ibEDZ3oaXP1lh7rXEPte9VL/AtPXu+8RxoqsYlAiC1uC2foc+cidrT0VJ
/499WU3dabGWbEt0dPseSyqXa+hiohpOZPFd6Vrrwhl/YKwR76SylEWPXQJdcUsk
d4lG2mB1Eo7mxEhyiYHI9BOmAnz3yTmJ/MDy1yCIxH7Wqy+Z/tDxuWZ5g0bftbTX
PhRlvw0saqSJb5BlUWR1MVA/4tQmlpkQcuf6jKCGiT4rvXojqjbF3sx5SfPpJ1Ax
uy7qCe7+ZYVvvz5H+YY1Qj/irSeTcwB+CQjDosvD53ldXGSYczvDTlJCPVKhcySy
1CU7CEXO/5dOG3fGesypmYnpSFffM5/cO50MoBrHUbNbsYAVgzqpokoQPhhYLzxa
wnwZWNxBwCNAa2BVfFOrWKxGpBUv7/Mc+Dan4apA+v+BOb1Bl6Dc53K6vFJM73YV
0nEFJzE5g9Xr15F1ELOFiqY1Ncstj8QDpbJRYeNVY1/bs9uyXMvEwuNj9UGpsNE0
r+vEg+LHe8vXD7HiWbESQRwDsV+4uUr7DlBQ6baZ932rvsa3f8SHbkiehtCm2djM
mxmObkEH9IvfV56+DI17eDwDGwz662S9+43UvB4MyrJn+28knCK8goVnH1T/buIs
ujy3YE5DzZ2004/kB3qnqo9NzzjeKhxnkvS3XvsjjH9JBUANtuz3enqCO4t5kuAn
lNtucbgTadf/fz6VvX29rXOYi4HSiQAhV8dKHWX8cJNd58MLrT4SRyrS8MgV/imn
k3EHNHqC2U9SBbVXCga3+b0kSqQPjnrVmCmrTJ/Q2K7RFbecVcId0mOFBOyuRcUg
v7HtHesLVyEHkefqjmiMjCk+hDpJgnUWlnNf+RJQucy/ywfjHMhVtukQerqW9csN
ttDpv7VKbOTQoXUQg1ayhhI30yJcf6kF0U6mkwZGipE6hZCrfDTODis5irZ8nygJ
dBadkQT1e3No/urI/pdRrKYUQcjoIdBabclkJY/M7xPh7Hz7B8W5obyZB9M0LBw4
vhr0zu7AFXviKmtWmkR5Jr+dc1xF4wR1Ag6Cs5kRUi3M/Lh/lym9jqd8tiu9Zy/K
Cxvevpz68ia5fXl9E1KzM3mTGD5rrGEQcnxnb0M1TFSgGQwNtQRtZLPqqQBBqgrp
zw8Gs2DDhkOylfEh3qv/psWkwoJLY0voagfRa9NdQ41Vz9o3MUBIcbMdfCt4xn76
4xZOwdNHbGvIJhq0BHvd8sPl/I8eMauGpuvw3axEgy+FJgWnuAuGw7gwlJQJLIRh
+6Hbh7zI2lfMks+572rJ0dvUJGOpX80DJH4hpbwq7cwgB+4BhfBSR9j1Chi9aaWP
n31wJNS5NGL7SIpj5ZEFPHG2uXolpPsGbjwLFN9fwA3a9Ksc5XOQDLnQ+24RURCr
s8m6Xvsj0Ema4Oi21w0oo2HMuPEim1Bn8nejhh3w5+FPx74YL4pHQzXxBcePS/Ld
ouIN1PP5u8XAR86DvYY3ryNY6b/p28ylMirTUT3aVuO9vDrpXfHZxQG5cDU4ZUc/
O3j+5GbBGqjYt5QHtKcLQsNs0W4raCQxOjboOScpZIaEArEyzMkS95ostTLp75BY
cfAKRA0IrBOnkNT1BYBm0J18I1fxAk3xkrjT1ryGcqNwJTUNUeMH/5pUOSV8itFf
DinB8blwKKzkaAMM7tKg511VV8OQpGcHPPXwxZzVtxJrwCtrGsMINHbHcoyhD6BM
BqqvIwWNsKpwSVkEIwp1m/RE2g8xIz0bfPVrk2lx7WkrrBZrnU7SrvKxkiuO6QEg
8SXAic1OByB/B4KtT/0pNMUzNyZliP5KM62gAQcbnmH87cnhIv+C8MOZuK/BEm1g
gYGzdUPvQ9iBEf2gbiKkE60GDiTed4W+q4nwFd6S7KZXBY5lwLtpg1eedBsqbzSv
D3uq3ov75f09FquNpK314eMyeGWDG9vzXwSZ8yqW0sOtCxDAuQ2cosqGcrNBHR8i
5icRwb+EkbJW3WgnBEiyD89VTtQb7sOTg/P81FmjMXVQISRdOqvGrybnpX//3IKL
lndZX54HG0b5rTPOfg0o+EeEvVvIzHlEHT9PoGn3G8julYZqi3OMMI0n1/p7nniD
IuLRJZsxuBhgf/4WshjkAUa4tHTUHIY96gH0xpeZV08X0Qim+C6SVO3F/WmSKpll
M6WuJ4uVZ1lwiNUqy2A0LNpLuQYOTyXKsVJ1DTIfUTicaV1oEqjjoFDDegeQ/IFd
CewALcHe74xNynZ4Ut9BUtxb2THdYrfwP8y615q4S2MCVw9LhWijoz4fmimsmXXN
Umc41IkOyQ8FmOoErbxsQJX6pcwgVFzUec0ZYgF44MWtYwTxzQBzWO2I6+b8FEHW
zdAb1k/S5Mwx1YC1FLhFY/5TAYgn8nZiu9b/1rjoYXh6Vhrl7v66NcqM4Pl6PUg8
fnEnYRXpLA3RfVOuDKFKa/UIoa2JckUMeLufwfQmPh6n8Rp94Xn3KXJ5hkEOWyCf
/Efv8+vScf1KDk8nbaBI7SApv4JUwV7IatdzMmIi/CbcR2p5ZDwJDNEapPoaq7TV
cXyPCbrXUce61cVrO5oQtpbb+EozmCqwEMcgGjQx6R1rLhET8UBpBQa4/W9mFRzl
AI9beNkmsKebXDqCsi8iKzkZoyuFNfkaXq/k1eNr9r9N8ink2Axvjl5xQLgjNd7m
Tbi76IUe3k9OUfw0TVipLFaDhbF0Nz7Uclzua2YNRL0AQYRfC82inrfgD/kqVp9O
o1KcZLN/GnfXuXACvrP7UEeSwmN1F7LF6vzhEWS6D42o7yXx0nh8xMCHpiQMNaYw
ztLvos5vf+AftrYNc75XJ5yhi3723Yqjg9PyT2NQNxU7x9DW2+tLGuP1sDJcFf0i
KHrsf6HFWxK5jgM7eGqMfGI/LBCATPspsFHq3gABiQL/3X0+RuN5YuxIRAg90QPL
gjwV6GRBLXtjEoVOS/eTtHZnK+kJA/9jbrcZ9gWOrjGPenCsEuBKO+EPMp1r+opw
y5fHKzkCTiaDyB5JfwcjNFw6LNjBdnkbhoUyfvssaePCVWJ01EIlVMB+nDn6unjc
/CgexrQbg9B1Z9wJvbL8HJnMwThHxRH/6dj5AUUZfKDN9KiBXFCCGp4liAApRR4s
+gjf+2yXQJf+6Jjei2x8W5+Uu5Ay/rUDGXtzBv0ZaokmXW7vehbDWZiguimtMloF
odynb4ZHtG1rMRMrDmDr7YpnyCUCJAtj1wO8VnpLCBL6YUYc1zO2t0B3o4j2bHM5
45+B+QLquaCZFeVeW6WrolNhXMz2zGPMlKOVxTrvazaQr8MWLLxeeW3+kKowttbC
bFI/Ba+WYVrsjJA5AgHW1JX/ft2Srf91RH11eSBXU4MiGcTUyZ62GGlpf+RL+8cP
bsWRCMN2AYJqhMRGKvxs7oQZVrfqmIec9kp2mUGaD4m2v3zGYhsvUDyByjmnE8r6
NkREOoKYi3vcQCUd05TospYwSfvy99v0H1Pl170i2DyRu84rvO0Hpvff8mTC99BO
JUVUh2+M19uBnww0Fmjg/JaW1Y9Tbh5QHs/ln/clSNEsHn6WWtzAzNGz97Mmtke+
aeqbtmqMEqcx6/y/8hvf4Sj93mryK3KuXPZ6Y0smwO3vqDqWP3aMx9ec73r3qCW0
NnKNmCUdDdvhELozDjvueHuFUB96R4h3vFl3R5nRdqmuYIG4muDMZ8ofOSJSYMFn
+6RdvPFVQw3WN75JEx7tVK8ZXCSRYv1mqviR/RrKh+cg/6T+TkIOSG5MkWiz4//3
ex0En1P2CcP/K8Q1NrdIn0Loa1Mgxmrlhqk4/esqxyPf8aABxqilD17aVGQaaiJd
WzD4iITYvx56QkxhD5b12Zv2W8XDn/YYQeI1KgrxFsoEXH1RgoS/nVHVVPm89jNw
neuD7lioF49KkV8Hdjq09CcaFMaFYq7TD8EPnDuifb+nuDwdfa6iC0fBLD1UuFFt
063Q/z+g2FXmMpCXlOnuOu7e+fOr5ppx+Q0TuEKkPOzsSJTntdbKCFoMbxhwLO+o
aHdAw6S/XI7bJQ/J56KK7DTACD6w2GjftANAid10nerMydaORQuU2CekmwrUQEu8
w4+PvApdcFD+k+OO9Cf0Z27we3AtyheSAqPadCpRani4fl13HE9gHCCQBlKOFPmZ
LvFGLopSGWLgqh6ZUfVLHyQSKZpiaXIGJexjsVpaVg3YsG/MadV/hIfElUS3CPYd
qxfSHqCWKmMuzVmw8o6cWJ5ZzC5MdCGD7OrB9mnZflc0+73Hgu0mqE/ZGyd/LRft
6b/y8wFUbKFLmnzKuvoXYCoJ6TTRUkwDO4FxenlaUwlw8AgTjuG/ugKg2b4qJlCJ
1ICKkOZyx3vzLIaWTUYl3McTPk1+kq+VIb2HX7LRiVbqFdkHUodGjHVPkK+NaeQM
8O7uK2YlPK0uKUz4BSHmky8emSbd4EcEitIS57u8xtbqmwF0wxQEr5YCuK6z4jBt
PdFBa2vwNte+IXIxDyQGlaqfkBvSpB4pJPiW5clpcQA0459ZTRxiUjWKAKvauFI8
+AJz89Y8c1QJSOUSaZ73kY8yABKu5GrZtusYL3/QMj984yYJVRfagPkfsRslpj8C
3RaWe46uech6vQIe1ty+leugN+6YFKR/uKFQBoCLvVRS/lhYJ8pCZsVsSW7zi8UF
mYIYqR8xrAvxU+iENiwounidUp1ro9vWiiL5X0YNprDHTy64AHC4KyPU8m+6dYy/
YWNOfFmQNx1yaR0k8PWxOrHo59F8f8aOx5g5KCKkaBHYWhx8xzJaclHjTWgaJfLW
lozeh2WbbxGGDmRjmf6OD4br/Hhv5ooX59NokEHM87nJ46K9V8XnpOSfv8b8N/Gd
yIbTHRblCImew7py83dzgshTok6i3jcCsphaUjgsVTvx5k3ZGhxezqlgr4VGsTfk
ui5/H5wp1vNqjQvH5Z6GLqurClvhqNhzFmNfdbj3YifFPUPihu5hzVKTlQopRniC
FEUFTXRzcznQsJxRXGdiUlOM2qmiA1MUXkKaH6EMYdIO1itzk39z3dchp8bafm2U
o+vSXb2vxXx2T4CMdXfNi+fLkgdN7Lrr44wZPgEpWDftcRTl3NO7HKbynoLruNtH
vFFBOqLbxT5z2rT3kOX4FWGPQK/82wr9fuom+VPJaCG+oxO+7iPgQLRsknzQA5VT
d/VpIyYWkNAcAHBaeCPu2xwezSAMHTBu+pkv+Rww/fFt5TgOoUHshO11AtvurQY+
/2HosiD2pyuEbD8m+9K07JQiAvrDuYfJHEErkX95uAc738x6ipglU6C6eDRU0xLk
nizT6QusNK26ZiRoP+K+9w9ZTtxHBbfe24Yw0M23db6DscP4avboQdeusJd1cSqR
8U7WnAx8W2Wg6bLovphUnZ9EqhNm4u7L6JIbI0VCS8XprKN09pr2btWymqT9OHdn
sRDf1hYZTuCh5Q1RpGFWlgWQxPSRc6w6qo5gzwi1jkDZ4tbnR3AeS2NlJEDPJpSK
8wCF64gaKpmaMrsbz1T+EkkjxouKC/DI+AKv08C3LxpREgDJRfxEq+GKjBlrN3be
QzA0E2BAbh+pS1bmkHGqh69Koizs8YZW0AX5ZKWqOLqzUAx10/RSguxO76LDhff3
pFR7D/qLWIbXKv0Z+61PU+EPE6B8XjB7Kx2Lj0Myc0O8ab0xPRlQhyXfE49VNDEi
TKgYHuinJv021KVrvBuovM+wgFttCfHOvEoi7ORyj4YGIC1GSuwppkuwmT9/+5iR
FMzBYsxnJpdW/uGR9hHCUCXIItB8TmuVFihX3yG99wd+dClfZ2e+HE9IJ/niiaha
4Q6chOTMxRxaFBfesUJUhVPILLhvd82jDV8IWx2nw1LiULuGF9Dv7Ygbr3a3L0ij
mdj1iyL2z0cT0TzyezUnYIzLn1B5uVC5wAx/+yonSMJc48O2FsmE5nOHxBx2MrTM
6rrl+PXpR+4ggQRuZsfln7uvvrI0cxkIoNa0kq4j5SD39a3gHfk/75XvxXeZv1Zr
JiD75iYj/gNzXETqK1V8SWbr8O5U2/7O6bS+l3qa1KKGVeCLEF/b7xjU8hq9w9Ow
W2QNt2r+BRYoT7mDc5gqoXWcKGeWo//ePeadEsDa9YDGF4sj3H4KwTl93YGrjxj1
YGRIlMVLLS1tBhfwnpRnxxqwKBNj/SnLKYPrsEwZ7BG/7AJeCNrrMCtk6LYA0a3g
7KaEZptgEiab3o2S7Z0VjN0aeWRYrj+qBoOJ/lpK+5/C/ilLQX5X1FO0T5N0mRi5
yiCbfs/FzVuOuzFRJABWR8poFW6OmSBMy+5VN0Zp14xNRPNBliKCl7lhtmb3tKLr
PKX1NqJKYxVvc2B89TAKTCfFn2+TeYfM0kDWdE9eam6leRwlIht3FNV32mkdkCxz
6T0CcWfl8pvk23D2aaOrVDfGEBOC0kstBc1b+gozk0NHJwOdlXpDIVMdC+Xiyi/y
9Jx7q17m2WjX9EJvEHrUudD+4peV7oTEma9yoRWHT/FMkpfyp6h3LGnZ46ObRQCx
xoaL903iTvShTa587UWJK9zjmKiTPxhZmt9kUd1nRzvNaAM6aexwddcidh43cNuE
QZJvlPHwwbd4025qbmU3SCRjRtDbn6setDwd6G3mhU2j5Ub+Sl3iB2128Vg7RRHv
n9eHQ+eUXyOfT0XgWdPmsTlkYsCdZ7M9auvjzkubCl3lXe+4neXvfT4QZYxs0/1p
Vl8Q+YEgdbatA8XBCEtrcb1/mG2rHOMJnZ3XvL3KeZWpzYfXJzX+oqiP2mDVBBaz
N0qNeONMAynBY0BXjnv3ErBhp9v2K4lbeuYKrE8GMn9nTc+ceOPhuoSfiEtR8Csb
VFt4hlA7nSpWd1pEmQQ1k4zvwXgc3j4vcDMqP2uUpuvlf+NkKsx5QCs6s29zJMe9
6UGHkH4iSJGawz7vIZhqzcjrJg+PKCh3ygN9+FOHxQSn2k0IjNTKv0lycck5EMdB
ylFwqchirgBcuCFvqVpZlU/BJmE0whSSRAAD9TZ+6a2HioCvlWH8K8XA36+Ae6w5
kwEpT9dLiDbYYxJEWUTRrActBX5qPa3lnIFkh49lQ58t8ttQzREVHHp2mRSVPIJj
NZ/Xw480cYFDs3Xysn8x2yiJ28PMzjU5TQApSuZdzGHdpNlzqVzSzYHYLMBxFWfr
zCissvpEtfUzG/ioM8XhcqqdLlG2i2Dr0RFMEQIQK+1lWyk9Qk7+mibZJ8WeMRhh
JiLiar/J1emi4Qmxk9vDyY9AkD3mCZqX2Cl0pwkSDivzrkI+lbVBa8h3qd6odLgw
nmklfo16F2eXAlF6zrep6tUdDi5kIxiTKT3lQX97OUIkepUNmaJ2lvX0DH0ygvD2
tLf717By76fXoP35L7wKr35xdKm01bfQd8fJwRaY8o3OH+O1abSkKhZTvTLiSzOr
EimYkHb/cRIO0vIzNyuPpNVy3xlRnpjzQTbDeIDzrOOQHOj81CiArmLndnuIjII0
a655NtGP3nXBOsyXbMDBy2+3mGdsmx+egZpOu+dO3slvZo5xnwyd5SPwDsSmjUnQ
KmMASPzldcfexAMzi7IrBhwJLNGL8pKX/XZx4KpSZDtSgRiFogVqd1gRmfREQMEW
sUd96JPWFMFOj1e+RdZAUZx2zvubay6mvZJ5H3RQceLbgEM0xJUDAR0cyeVfG1gH
0645BAFUImI1IQ0e+ZlnS9QMNJFXmSRQrPAFzOYeWbgz/zcZN1t0R9YxZtVQbPiY
9jAagP60OPvF284kvMkujBfBnfMcn5bPHITFoI21mbp+XdW6nddiG31I1E3d4yw9
m4i89+qBfwrgWNRwKpwRpwHgbuuKEw8ahxSlFH0yEqirN7KofGouBrPvZVnlsK4q
1O5Dsc5dJE8p0/X5beeKUKbgt/A/9jDQRuCE1YTI4HqJ13kMm6HvV3aX8+uHyjXp
XL3MY+1SrppOy0Qr4llyz0RbhTn8wP8tIiI4C72p65FN8aGvo5Zv8DkJH7150PFM
ALwJYIu4TPU2CxdOUOEx7UC3J/C3/Or0eGoPa1lWq7anUHyZGY+rw8xF6YiVpLPU
4lbqk8XNow7r2EXM6/dk5B+jZQKNA90XSYCUo1ydTIXerEIHtWL/xjA8cfQHxV7D
vF+lisRo0W00lPSJgyQcvX9Sm3OU/9BM9Y8QkKzLPPAndC7NOR2lxkOTuHKzZajM
bp1jhHi9AwX3bg749iRqR3xR/7DbPTOdZGa1fuSk0JhsYsCgGOB9EQjL0Z9hDFaP
6tWz2CNF2peNEQpOEXisbhKiD7gp/GyF3z8czO5/ibvAwE7DMtCoc3CY5gwkD3hg
rht0OpbTJqW2qlPRUSxcakKchRG1INJPklf6QvipE8WD48Q1h+arbMP5JmjjpiIx
JT7nblekCw4RfgN0H1vwC6Tma28TwzCSuWTvU0m1GZTg3lsCy10sR6ujDHiznLNE
T3fG9oSOqE0if1BpLy1//lBld/iT3DEu073tnH293LKNzSuLwGXvfnNDz3aX1GrL
SxNUAE+vWp9Y6HyS+HyBEV02sKycpmONZNCz1S5/FQLBWs/7cttHqW1K0+QJKTCF
IL2+OSvZw+b71DBaKYLuCB7OgD1ji/Gv8pGe1V/lGSR6OrK+ToXPShBbserjnIvF
9s+d8DArGROQe0flfO4yNR66LxIyeBG/kQ1jz9lBCfRxKlP+/ThF909lTB0TfpwR
bx3pe666G8m2FA5hNZWZg+PrvSzcbt14PKrE7SlM9M9LZVDzGc18QK9eknqEyIRg
uELkD18w2lM6kIPUqGen+i7prvU2ALD4y8TOphX9/a0=
`protect END_PROTECTED
