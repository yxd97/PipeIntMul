`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VkiQiJf/aLBkV620s70GNi+p9I9MYjSkG957xpHgnoiZAsFsRDnL10hEYCsgsEgq
EtPsDIg/Q5cxJpJLipeRRlk28hjY39/jBzNHw/M1QrQBbPfs/q0qbvKuI1LOiels
MUBSro5jOmYiEos5CqAWCi40zyyQSMe3WiJmrZmVjHqiqXF/dv9zSDyak/TrceNJ
BGpUi5oKKwMLG6wNkQTpzf4+jNNAhVfE4B2Jb/CjUtxqwQp4Vhs6ve+29tIJ+WJE
+vd/kDp7rrsEQh/OmoXqfh2H4GivgxvUh95LWX/cNqHok9OnQJ3hicXOd49dOsH1
KCfNap8GP081sfN/OJJw4eh1jB0bWG7rPR3x50xbnE0J7oVbYOuMxF+J8KPH+iM5
FA+cWKmLfJlAcZ96UoQUuA==
`protect END_PROTECTED
