`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cYhHx/wj2P8r8HFVhZCI1GfnDXldT0hz5QtkeQ9dAiPHEjW9BJpQkIFv/fvfe8Nq
xzPNnP7pKHmg39TD21QSrOCACNwnEJvmz/eLWUNx24zQWbqD2hwWpmr1xQQrUNeI
8VDsUf/qPK/nePBh6hg4CBq5RqPooqg9zgwn3iDgKxN3/1KNYoC2+1TX7rEAD4Oj
R8zviLkIVQlfOxvQKlKHXfFTodV/a1w++DnpVQS0IMsdpP6dJyed6QINN+/dRYHk
oP2SmRv8kxkCCtowPUwGZetSQhSvmmSd2hbp0Jf8ak5X6Je+pdfPwc7j2XKL/Fg3
QAD5RCXG0NQfvXPKnXPf/lJxvQvXyGjgSFvMAuTu1d5csHmx4tULKdsjtIePk6T9
xtMZQhII6PoN/tYqUJ/bYsD6OpydiZ4Qr0h9T97qHow=
`protect END_PROTECTED
