`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AYFa34VTtAlRzu0DtoIA0guZUDYHo6/KpNG2H0z59RVvStNtzd1PkMH4Zj+EMP43
3ULRWLD03NKszvBf609xOf2Se8SmOYkun4AYr7vkakST9YAjjRlgM3rURHIK/Jcv
9NGDNG+RwJdhtrafiItemkVS+qeqpJ8UvRn/m36LXyWvC72Tb6Ll2BvJ3QWEz8gB
juOF5o/KWGm7+eJipegrwvijMMv5iNsZ4T/J4DHpBAXA3HdmyOkSouEfPPCP1s6K
6GRQqqbuegaRXylNeuiSar0bszPePMjcavxvxU2YNs1CN+hTWI0Ff/Uef4UMLlse
cSqkF/jTymVXbOQpb9SK02hb2hTOw5NMRyqpquvBsZ7oUfapSUURvtjorohiZiqj
qgX5M2glAt0Txf7h64MbjIoVbOt5Dm3knO/uUXCxXgqIsdSwPQ+4unS3i0/N1s9J
`protect END_PROTECTED
