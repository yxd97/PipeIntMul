`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
felPcy+FzAK3McvYl1PtOT4B/+vGJ8nVT+oJ0EV7/zYtnn8DDIQnDSrbOtEYX8Wi
YGzycrTLn5WZ5jhG+fAy/Y/g8Rdn7rJUKUNWPe5FMTXLa55SALCDWW3zYrrKLwN/
RTEsOC6Qx2TfjZFJR8RNKbkzHlre3ym6Y7O37TaaTVKA03KdurL7cLSGm+LdXsRM
0kxluYx1VNAnxciU0L8QDyD4dUoIYvnSI0FEP4tV5b6KjfluyWJh5Gw3X3rdh76p
ASVvdGP/AR4o1iFpvqdgqphz462j7NE4j06as4bU/qV07H92xoUiSAeq/4e4Xvjl
9Wdpcv92WqIOv9jsxBePGgNffV3hBCUyA2Pqm18aj4Wc3ZHWaumKdx2YcM1/6Vfo
NwRiDuL1f+xLXSl81uG9X8/jrJ2ABGQIlMpHW+P+R9r8rEX4RT+p0OA67s+DOExY
b/PC3ImpofAN7zNt/ez8zve6VKtaHHUYVBrZxtb2azqTOf9wR/iuhVyUeH19kUXL
qJX82ozL99HUwQbMVUTDIGIQ0qTGQeQn7j4LVvEiNp35RuvH9geUxhtvQb340VI8
d8W/ztNGoh2ze+cOA+zW1MezQ17aKT/m1gkVIRSlT+n4zd3xmJQQyJTG6xb+vA62
vXJCiIyUHm/fnuvKnCxUSD4QK1lSlY2a55xltPJMmg4CmKxS3Urh4zEfg9PSWJrT
sFamNjLXMwG5lbWXB++XeYJThl0x5xkz4qfZUf/JSDcEncehRnG29ERszi7zfk4p
6VIMyy8JhwnJi2Df7WpWzWaUhhOdyWwg8ahJ2BeWvnmhED3hmCOJ68/ZUWsuHO/P
LYUEnE67wiwaxLQ5+XxuAjEICvfgf9ovVzh8OpSUgTZNPwKT0KrdA7NFcgaIvlhS
mj+bEKvMg3M8WkcCyRe49nDIwGBGuY3HQbXcbDliBLVZGIYgdQXDnDWa8OXr/aMB
hN4Zd1EQO0BHPvNbX/klARuCj6dyyczHFs/pkQDXwLQIpMeyKhpzaQdMbNSJA+kk
tpyj5LfZHCyaiw4yRdMsOmXNBSBwc6sHvVGutn6XgAeXSv0bEidieLXvYt3bSLiN
2+WzAvdIRKre+mkdQy4kG7rdZhl24PJIXmzM32HVU7Q9gtSZisR4TV7c+mhKCnmJ
2lKsT8mBf4lONxp4YaRVAb9JI1mJk7Eplunlt4ltryAAew431mQely8VuLIh0ghv
/Bc6ciHsrNg2QsJPH7U615lDdxT5P2bxVEzB5///mtklYj85c6loM6jUSqMzKMfv
tLhSZ74pAhOzaE6l8IVqXaqkR869AbN/bojKSHsiGsM7uxWHD5LE/nR+ArWRcHEC
pfYcBUcPXBdbGbuab6VOjyd6bq/U7j/iDi1Bo7oCxV5krXriYzVbFpk1WhZO6YBD
gwE095prHltZXvBoF2y0AClVtFPoveU8TWMCmRYdj/B809f0u/wdTVpfQcWRMG3O
8KJQA5Y9OB/Hq6RpTukjYwr9IFxNF57N4Fd4ww9NP1m0HDRuF2KXXwAlE7TipbNZ
npXJ6j2pgbM1PTc5PaQSFjUWKrtYXscrk6brwMJmm0Rj8Q1ZHpyD9qi5IiqAV4Tx
TfczROk2pTPLkyhT5jl6LZGsCVWBSso43n4vTY9XpEQvnVb5PZuzUfPibI4Ml/jA
9JetDTdF6Ooyjar3EhW9uOARzpLE8t6UKX+bzT/R3TxQUtG1N5kHJ3EZYtyMQ4mn
Fkg2YoUk5QEKj+TS3QM1mADSm2CNRLnuv/2cAqn5JU38Yd/IemQ0J50nCzSRLB1k
5CesITt/e0TMs0DF1qBC97xUIizVR9v5bGm4hNK5PmT+5lQ4xQT7Se5usCmdZWPf
+2lik+FEPbuCKK2mPAYpVsBWN0Uk2BLulCRraI00OrudTXP8Ytsp5J2Pe/+bohmy
+gZhrvA+QnEk2FrHfY6iAol93BrvIkJyLSUJreuLZvaj3hZC3SgnqIRRVNfG3XRJ
MCQLMKoakGhvDIbrO/Nn45SoO3IXnSXiJnTry0niRayl1/zbZw6t3FYcA32B4hSf
NaQXyun3gJ6QLnfTvLbhxDri21gsg8tj4WQ1WNq2/RRnSzbJ8jRsD2+oSFiKKIAh
LZGlkA6cOEOupybPGmY0iIn27awJ7xJ9Pi67rj33PKU5EsF0yLp738bgCxLMAlIF
3YPfWspWoC0as6gDtXHJkz+1x9AxrarS+S4sl96aVOTKk6ZIAGmKe8EDSeJiH2ID
hdlt3PJAbmVXHjw+C2okdho5HVxoBFPSO+7V0qke8fsKmqvCQrL314ln2qPvxqGv
7KELBF0q95sq+I3pLacg5IqktycR7NfzEqnJBWkkFKn9i+Xttbd+SNK+mFah3yz0
P6gqaURp9zmi4DFkymPw7TxEDepwMR+gKdLDdpEXW/zV0ENux4SOHnwmm//cwRKt
dZXOutupg6AbdK0zg856m8FXLJMCYfQwUc7KhyW2MKbBzJ6bIcYsxIz0nE+8NmV7
q+bhcxTyzgwk5L13wuPrSIYkKnL+e1+Gtpd+G+IpHSWHvhNSf8nNHT1JTPC2ksHv
6ValRBBOhR7NtMaubH7zIn0rI5SVAN+BCTZ1/sLpUcSZnEyJ0K+MmSoArGKa0HRz
qhSEue5wpo7IL08momF5N4IZNyPoE2rkMm8a71M4GhMdjlq9bBJZqvNnKCy2HeOV
TbB2WdWtiVq4Wjc2FRiG2xkpe/vXvrYP/HfMemgD1EflxNJs4QZD711diQLcsZ2p
41X6GKZY5pY6eLwSuROMb5fM45ByWjs7QpZsG/o24Mr3gSMAfSLn8xDzEWRC0Gv3
NRdgfia+eW0DeuON0zWwtoqd/9vfYKYkP9eVaCUGuL1R7jNBgzpklY/o6hXwWiRn
bn0mm7kftmw9PtURCYH3rjZ6ZgetWsp1ZaDRQRnHIU6zSlb74a7aYU9dA37lftIK
fG6aTxgdrX2uZxmN/n9Sd5ygyVLl/WwvP8I2nOtRwEG1VFiYpHBDOlv62juSNIfl
8cgQkTTiaJGAcbW9UjQy2N+fxZJHwWMyWB5qD1Eoq5D5Z6mpYHf6uRkSaBwZcw2c
PtwwygX9qIGKtm1nLQnt73cm0V4FKK5f0QTcM4EgEiYYQnr9AqR/ZpJCfYNtN9U9
12KNa1HO+Q+VmoOmB0GHQ9Dj6ktb4mxhMiSMhfB9/T6e1IUSsr/lhzi7cLYTBGuA
j2lmHKU5y5Sex6jZQ5lAfkuLjUR1fx+O+GvLIo9X6pmQP9A90r8TehADwXkTDkVt
RtqP6qcBz6aR/hijHOD4nschZIjRYots22EiCJqKdaV6o1/1M51ZZFUtXnkOVyTd
Hs+GdlMVx8vivOKMtLifI7EPPkE0Sa2gXs9ANfpUBvSDeFCyisoT+NjyvKKqh0BU
22OUHCx3WtTv0QTTvWYOCvgO6b10psJtSaEBSdU/W4GWlZsjIa/Dl6CdJhdS1gGX
60b8ettfgTTQpERWK4/rkwwqheYYw/+id99RLlZm/27JQh7nYvPDFrYeXzxaFpll
W6g10MCae8qxaBhJCRuomCLq3lyguokdm1gFVqXY8MNmAcO5KanTnFmtKFRi3Rmr
PaaHLfx+vuTfRPQaH3iZj8xiCiibBt6+8nMmd06dePcQCE4VePStPhY8XtmBYfCV
9FKk2GJEocChHpAxxSLkzGM2eAAW6l2IWCE4QHUyIgdA/DxsNY2TEPydFO+AdC0Z
UL/IsaJ3MKUVWB/y2LoAyweiCT4rXJUPWGPOn+7BqI3MYBHg3tv04rCfpn3d5e4k
Q8HAR48OZCeM937K3hPHjbuSBfZJVyOQifFgvqeeYosr7yfotg/CDvTAZJyp7bN7
vc06RTvgwVs9H2v/8JeiHfknofgn4switBZtITAN89NwQkzXs2ycCLRLuI1QcvqI
SDstBvywaeiqixMAs6k7v/7+yUND4k7cB2nD8u526E2rcoMk/4l17GNBAIIM/WJp
HTU9AN/oU4h8fvD9UkLMca32NfzBSRxGH1k5qz5IcF6rLSF6/FpogwQJjWJkEDyF
tDREhWjzerqxWKrbbvyIK2FoJg58M1wF1CXDy7kOEc4rOmXvzxAOA0N5SA0KZ2R0
7ypa+UzFbiXxvB7UfZoMXld3aiijEGJQB8O5esEn41aWeW+UmsFBvc4hqu0e77ky
mp7B/m9t1bYIuyEhLwayuIsoW7LThXuAIzGHNswPTtxFASbTj9crVNr9GbEHjG32
PI8yPpFOMVrNYl1gocorIGwOS+OKt7taiv4MxTlqTZRjYDMGWg5UP/4C+kvMRn20
cstta6y1K3hPenQO6/qkHdeKKN8xb0IhsduRdAnaAbX3vDRyUbU0S33lZ0/4U1ya
zkPV+mlpTcrJz6iW7UJTEjtFtKaROLkqYee84ucNzvIFPbsBUqTTboO8tfV1IfOh
J5pLVfXrfUDgxLIQfBQ6lc8xrRCP94aD4ZsO+Jxo05KVEh5n5ZoNUHgYYptnToLm
R+4L/QDxxJd4KisaNo51ZM1/GfIQd6uP2R86MtSk9cKl8ckhRYcWefTc995C1DZS
H3hWdbR0Vp8kKVwiLOvvkJTD0Hh3oXZbih3iPNitbwRfgep8qiufj+QXoBKod+ny
WJJK9deVuGaN5IXoRzO+UDFviyI6kIOoLMCYKeTngnp4ZmcRM1emGxtbvzzrQ3mG
vMBk4+P3TPwNVufNpBDUcNFkK8Sc7+hRYlWTnpRaqD0S99v/0rTY3Dvb6vunOAKH
yOkv+rk7c+F6MCAJdRGAw7ELHtC2BXgRWchSb1xPDC0kGenOZtVgeLAMePaMiXdx
tsW/LjUUuuPt/EFyykvx9bjwbbmWEekl+3OkkRt4oMROcgMArhfetqJrPmf416AO
00Sx2zkh7no1uI17qPGPeL+1/deIJSTC+JO85LJJjsVu39ngwdHPaacr/vVDl4Oa
i83HQyY/KYR/6tqnlc5tWUz/0f1+/S/nY4iKABGdZIwO8b34HHxTAA01jweLyN21
lfrzilrpungmvq2qCya5Uzwq3KWibX9LreaSezqWCx+fzjYhwy5z7aVN1MlBj3qc
miiUh3msqxTHNyuE9J1FMmwekRUaQIuBKo879lZrtvsJpUUMb7mLUz3cHJiPUKsc
BV3hek2jfAjX0xVEcUFPDZKKW+iPxC9UtB5VroLolWHV+dYgqSO/lm7h7hQNKj92
WZ4Oxy1uv61APVbbGAjKbgQE3BB+6i1vmsTT5fVMsIbNdl/LVMv6FwEO/J10xEIS
UkECnOfNQ1qq2Q5/fhoBgSgqIf1qU57JcOAdNmieGQ6RX6o6v7E2ticog+u9hmqm
J2YHTNYt7sm3oUYOuW8Wk9fOD7GlmURguHiwCz56QzrZDJ94DNYEgdjftw+LywSK
51Hpwa3lNkSKdabxch917Mkbh60oMTNQAKndPi2tGJNNoXAtXuN1Spgn7kby5wa/
A9U8xTfxm8pqNPLPUSR4JcCXj/yQJnsNJVbz805AVhfJk1zJQDjCv9kfhjl8NYd2
ejooDNsSUAdbTpnnle6FIN52GXOnW57W7A4GhBdI/MG1uNKkJDzKnSX0ZnPWl0K0
zdsEUyznJqKmRs0gH7ufNDMbAQ4C4r++hOlU+PK5uLMLYGNOSb3RvIPScZ0p6Huu
/HbFcPRN9Qej3hUT2Z5175jGax7fvv8D8eWG0ErIqJEvijGKADPwvDBivpPtGjoM
Bsl6DuRyXUJl7KaEWzF685fFBnecYE6SuHYVVDVo4jmSLIyZgJrMDVNXxW1eFef4
6dZjXy5HesWk31lyfpT20XlGXLICW7SNpulMA3YFBAteBFdhuW16K9EiXQS2yJTJ
iWMbHe8PycKvRkqmaBcTB1yFKf9WdqslY29ukMqODprp8tsprqUyPzx3G49vm3Xj
HN3Y/xClsUDWmPrWY+LlCSai2DjIUC0KBJMM1b4tBYFyhtp0KFCeJ0NbNuryM8lY
d8yjHG1j++QPnLQLElXbFW5vw1OKDyoPWcAqhjVeqJUe97VrvOFbTVIyyu57UhN2
uxvlHO9raCxsPrpS0in9VNgSlaOoTTTC6W9G0ShImyPRlcd67V1o0whApsJU7VWC
CN7GCLKgzV5Y2u0+Gx22FJBYgdXGzQ4QmwtNM9SlpP9QUPZBrKhf/VRcXYfMmcEj
X2FRux9MqzFgWA7CoU0D0yGMDLk16q66J/AltSnHif5sLRctuO/GbzlsbLJO9/qX
hGGA4xGSZ2LcuCKa98uMFaSCuUlYH8eEdEp3Hy9x6cWKUnS+A9UyBvG+edCAx+Tt
9lK0J59/maTI99uvzwVS0pyTJqPQPr8tWJ8+sUHJIa5Wfd/IlCXQDmxs1/4huNR4
vksAJaUr1zjrH1hrEwVtTxqUv23Ggx9JH9QfCUWNIoIu1OQQW+t9cBYHuqQsGiPp
Mu58wmICjXudDV1QiwPa9IOlONjEoLTfMe4AKx8ASzzvXHYVUFtujpAd6r45apOU
c1D8smuXurzTtf8Pkbm5D2P8JfunjOZk5NWZkkcHPJQGX+1ElKypRDUKrqxwg5jB
AEIvAUJ7rVDsjcwq4H9zPxet4Z1eC2DVtyDPjr3g6zcaS5qjsn7e0TcaS5MrtmQ5
QP+RmZWAF403WhR7kOKYBg/+oKEEyEVkeoHoRxNzea4PT+JrcA3FJm3qZNujBLGE
U2rILLZ98G/Z6sdSrT3oKBjofwDYHDmIImJoTymnDPKUS9w+0EDakzLeXM1jJA5O
+9v/1I3mjIJTnaQIN8YSl6u7junR1oKIdgCfJmNU6BorqTQ+7xoayZJpOO8VJdQm
6nVMlPEZzXgwrhQl0s5GLs5+VNLO26A+uYrXtmWr3F8iAT+1BNOrqlqP1uapj7cb
1Th2K+3COwTGfWFe26/tYt2SkJqPz/fUTNbQV0U0FuITDmppE5H2nkz0W0cUQKVl
GGeOpSdJfv1C8YUJzuQDirLlpBiYBOWy5sC6EeOpJL8eoIAEn8h9NO1NngJAjjIG
EBpQNzXOsrmLafjVSnoWG1kVvSiKYdnLZysp1MBhyTa3SQsNtLmFapVIx8l6RtTh
Aafx6ZieMJHVDsCigRLBNMxwCU38BgVq8PRaw7zuG23HPU9sFxBjcToMMoN2jp/e
S7H3f2S9YryiDCYpsFVDC0qt7f4onDm9+WtIrq9WWg+38jSmUAXSO57T5twIgTF0
G+qNdAMtohCZSbc6pOZFOcHnskRwAJilxe65HJZK/d42DOf74YW85F6Te3wl9npE
GVzA/t/DNxfhiAKkAdQQn2+GEW3FDMMdpSwZtf3fVep6dmcCGvPUKnRSEPctXcmN
Hlz70lXG2i+VYEq54hsxCLCWHNjIJQxmwitYaMQk4iH7W5gmmCQ5LHvglLdx8U6S
jNaKloNLiWdFrXEFivJtoUuxj0qELBgBvyJFty2FRgXgE++iY2Y7jAx9jPVO2Ttp
A9Lr8wuxBRaInd+TX5pRXKAhMVIbxYCQMlp1SuXK+vIuow9styYk+uci0iEJ1Eoe
giwGIxfnkR8xNPdNthxr1mW4dqrSdUOiiSnoKni6HtpX+5XXAkQ3gupAA7EZbe8n
6+VjhFpXy5VgSj8huxJUAhQpMDEoT4lH0Hydv2H//Vz9You78lO1tss5V8R2OLZu
SepGEKgReqhsUoRgpxATau0gilWIskT4ZRX2//ALoSsC2S0aCLwzgneAzLc+oQ+I
N5uGZPxBCNkCDlSxwTNSmklMOg/82BGL8WhNtiffy58V3S4sHU3s4yj4mTVmUZR9
QJW9ZMTCojzi3+uMBaRMy2JnFG3voLBOA+1boGv6hjoP30OYTOtpCabYiIrl6q0p
Y3mvo+x/plfMxnd3g7470GX6P4ib/rG2I1yx7b1ANIIt1GosYC4XdyhvPxddqIcN
oGO3D6U0Trtj+vdlqrMdlgGOMX+Dr9PlyWnTOamV/Ft4VlbP2ERqP33hd44DLeCH
aZG5+LUJWAselufSXQeMy/4q6PkTNESrrs/dcdopNxv0IqQgch5xL0PFLvFQ4miU
p949Jjpn0bfIoWzPw5VKRga3dBLa0yQdV7BK2W1pq3vgrQ4q1ABcY/D1eVf1wJd4
Zgk+sH35DIzJDWTbLwc/BVAziJrDvQOOsYci7GB5anlvRxVbyNJOGwS2Wb8HG2Bn
ctLJQ3/Fl5nSqSBJhnaglllMQqaseNuI7Kl/KKjq6no=
`protect END_PROTECTED
