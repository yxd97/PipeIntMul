`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F9a7QVT5812veiCJteak2LVfByjZl7yeCXTZ32N3VBW8l6jNAzXGiTRo2cyQTW/s
v2nfa1+Mbt5MVH5/BiTmzzmetzqwHeyu43xZJ+bEoPiYqlH1B8tB/5gbt4XbUALk
L8rkymqxBlGkzghPXr6hqMWg4crF4yA0oBWqgo6XhlcxCNbCi/WPlxiHx8Ux6/bD
UGVILJ8hoWZxxiVeo2d0P/35r6BnmscmsVsVJk/H3DaLEKsTu69Lw2ptET0G9lIx
wU9OCj8MPmMRqKkZASHphk7IVgItx/mmNf9CtizT8uvho3a23D0zEjCsEBZsUsSC
za9kgq3P59H19Ly9U5jBJC1nrdGYHYHyskwhQSLZVzMivGZv9yKncQp9vLyRUPNk
7qlkbKKVeQpkSZoNLx+R/keeeLA8P64JpEfMPKMkIfArbkkwT0GQ54p8PwFEb7+C
3qcMs4PBgim7p7Knzqjg8hUcI/Liw+I2XKGTeq8O4iRyDp6+eHCKAuBkjbMRQHAU
`protect END_PROTECTED
