`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Or5BOieEboQj3Q/rBbYTBOQBI3juE30Ty4IZvYyhnG2vZwN6Av8/9usaNl12i5yf
j0xaRIikwP5qbN2kLK1eRFfoq5inSW4C0FZaRLN/CX2WAC4+NvFb84E6oPf3BOzg
/a7OUTimoXH6lgchll3maWzrgonKtKVU/g6NI2rN7GMOVy8+E5Otjj0iikDVno8F
FeeskuzMUUdkADt0C1FRs4PlpG9pYqUUPhp1g5kZcs/4pyVTqrp3gVliUNLr0xG2
fxyVQkcto9zKuQK2RRsiFLz2xaoINpE5i+SnobFjYA/caV0VNYl38RPjFGCRVBr0
O4rnTpIj9TNugwxIDbnDPsH1S0WEkgNgAVYfV59ts6dWpNWcP7hYRIDW+BmqCNSO
TM1qld+LNyzmKss2+ZhqXOYfUyCQig6lk1Q1qV5oZlPYkkCfDFiLV5lfE1hlzSGO
R250zaV5WoP+qwVGRscxNYKIywtEqzkJtFWkQkLF+yjYj7IimYZ+H+U9U0TUdpPF
8RXq4nsSMFZ987wY7JMqDCq28ge/PxlPl/yZzZ7251mvrMBOAqJMtUt0KPWVoxht
7NwTpPW1gt/6lT9uOsl7dMDNP+Hatoz/++ZuCtC0hyYU0UvSOsU+4bBbXSzN2LFW
K+S4jj0gVtvhhzfLPN25APfBSrz4V8cvnMRXMqeoaukNvt9dxRas9EaWMO3fljlO
awlVv5fxr7WqcAm4F9/nUtPI/LJAzeXHhasE1l9SRUtMCTtI3yY1p80Y28+FMQSw
g/s4w73o+mih9G27Da+uq/97ETtlITgghRxWu4AgfwPdYJ8lss17NE1BH9c/Xequ
2ypIX5wbXihWQzsExnEeqURmdbEwoOo9Y0IPgmpA9+NnTWWfZtTNTaLWw2bSrTGY
MPMkFdfwqI/3KRzc/b1a4FdqfXhhLvKHYuj1hDAgvrb2UhD3D9gurmrcKZyyAEOH
`protect END_PROTECTED
