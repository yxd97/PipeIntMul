`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sgaUy4xHS1kit9RcnpxUC2wQGUWkEbCkGqZaFMaAvcwNyVMgx1X6uzE9o+PaWlp8
EOT43Boo1UtE6EgpPt+Xb77V8tpPgToGgzJmWwXZ2CQUpStSUwI1nJFXFPwRrELo
VE7nwk9UAumElsAHwLsU+SghOZRY+HfwfX3PUp6+BttjS1Jz7LbK+aZKnlwNgpUH
fHCoEbnAk968iY/lDfjjynI/6Yym4WUuRnXy9XV4xHKyo2d5bjoufm6oB0xzXWiP
MV3EPQ00VH2FQOoOvFh+PgbDywoueJNZP5ymCKNZRBXXk52a4TljJhDplzdwqR0s
ao0J96XIe4Q8j6E2rllhvjBSG3tOOBLoQy0ZxoDNFHoQYQvMy8OAStmr0Hjd4zDK
AZyeFXS2rHKVmboRJL2VOnIDK/j+RVmAW4lGT8SGjZC7lCtn/Up+6+j1FsB5X6Zy
3J4hKm3eYgAIs9UOx3cRpx8q+1Apga6WvKMNHcq39BO9ggNEw6kt3mRKsJsGLmvC
UHCYF8xLtcwFj74XHpYmP/s/zeWJp+di3hz4YWBmdIULgWw9jwFO8N4RhWJh2cmf
5V5FXTEE6HIO7h0OO1xkRAVKrw+4PNR0kP4394/rKn1snpkNQVatMbapw1Lw/Qtz
+KCoTR/Ix7rytYrBX7vfRIfVr1igQ0alVqIBeId8eiZ+83I7UT2qcZdiJrhKeFy4
GFYVoVLb2zQnthcGHormKglcUkbIeeaNOrPxLzj3wVtK21bhUO7lyObR/5quDE7k
XcOKONaKh7zlNeaSQ06DvS63aLn/QlbTgWTkT6zxDaFhu+b/7v+NQchQYrac3kKY
kVD8x1T5PekmaIfd36ZzzoxI53c/ch9eodDLfHXxqIzo90A5g/fNoWMJbfgiPQvy
6hrZpLBVILcqsDfA2VdSn1XYDMXVDONtju497GAy/DUxuom5ga83jSXIYIWoQgW4
Kc6XSSOyzEHyrkP7JJfd1c3shlCAIok1vVrRDlLnD56gAQstPr+CqwJ5QTYCOg3I
tBFD7vBFjlgWewOboozMJPMRaszqBKsKX+YwhD8BcwDxKBvk3ylrAw7lx7Rag97e
SCFHKLE4a2pjyKi+6PgyNrPV5uxnglbhbO7InVK5uaUQL86xNhfGTiEz443SGtfj
eERJvwOjVUhkqEPpd3USlA6KYC1mXO6ArruBeDQM5KFo3sHu2c1Lf2DADIHdmfH5
JHt0EqBUXXmNQIdf01BoMPR5kv26uScdci2Bp7mRZen5UkrCvjcI/HTq/wCQiFHe
7LxWBDOtwR3VUKXmkC3/hwRuyIctGV+B3ApeY0ZV4vRy5joUnLeRfoxJkTKMcCEO
hQHFyILfpkvmmCMDhiHhgc4bym1UdRbDLFttM23Qa4291fxfBVqKR4WgLZp7pm3U
Ij98xF0h6nttUM6BzCGkjpmuLI779Le8ZP5zGVu6i4d/GbkqeE5eRBu+2IW47den
INkS6qT2PxKyUePY+C3SCSP3EOsLT7iaoHFB//CSAADAxLi1LJxzGzrWb6vWWeIX
cwyMgVxzyLugREo3+HdJEFyYLU/3CqM15QOu5Xe0EGM0XbPaplODaS58jvFF+fbq
pqknyr8cbMR5DggXio0c+lUIgxkxr/9W2F/fwsRbMJdLB/BZ6JNjg7DWrxpqNgiV
zbgPAn59Hm+IvleHQkJSoesCADZxf/69zyWJXNEyQfMEO9g0/qTz5jDsvc+5gLpN
XoqQy2FxA0A7Wc2/9pQYF4Uw4wlb4OvgS1UKjtU899webaE8fQusPtVqSdYd2FFb
hJf4RzzxKbxTXFwIcGNYilkORDe4FSsQZhMfzj8Xk9BDhOcUrcWXfb0ErsQoQQ50
2uIloSvlm1IIWRqf3cNlZaqfUJMgPmeB/kh84YRuflxbyGEMGFtVPCrjWnpBorzz
3hnMYlhe+V5BsCPKQbt//bSH2QrhEq2C1Xv+tkpKaOJDCTjvBg9m/cg/sm8WwRvD
kW3NuryJCL6C3HmiPSqPUJk+7ua7DFkjvDZiVyh38S8dFE3pknamb2zj0+fOjr5G
OcJFJePc5uaFq8xZF30FmrzJHLCFG7mI1UWbGnNf3NP8+RM5k5AVkwom4yZP9fDO
gFyP/pGhP/AovarZwLKKtzLZO2px6BjKoehJeiAqZA0nDVijvmA+Kg5KxtRYv9c+
st+7GfMAe1K/xL1wxGpa369oh0K8fs2Kk7lOQlakl9Kf6Jik0YKe0If0eVTrL8ws
XB77P0LIBcx22bW+KUZzbfMj3AK8H7hXy8+ScitmrEo3/DzzsbnFn9/A18Xo1vYO
zVyobqf3jrfxOtvrlNogIJuyMIdBpT5RM1Qz/4dumqaSiEXTzTS0ZJfcb4zVWO/X
UOCYN1zYq3P7qhCyomUjMAXtpPc+JnApm1G7twKUANXZx4QTKNBtn6Z0/WjhvYwX
BlUAgmc9fyqvhX9M60iHfbus723LuBwP8aR2vqrGC3qy1/JkM8vRqz73RGXO3gFU
BW30mwAU+iH/MoNcoGhOY5ab1XZnEdYriE9jKLsQ/lJunTA5RmUpCxTBkMRnn0rh
sRhLfJjfWClOIIBJf9OctqL95aw+yIbAKdBRGCU7Y/Z7mGHEAcvc1jGAJA3uoeb4
ycvKHTlkPrG3RtjsH96ajJ8qG22G6AwHJpc4q7QKV+mlezvXELvY38t+vLEnibge
HrFxnekUZpnEABEMCRWC0/FWg6NbCvedqmq03dwqM+EV8923gtRh7Z3RAjb0vC5j
x9jw5GImSMGZFbPNy5NLXpFh4tmBbZ6Kc/QVxE7oKjUHO6EwTbf31PxRvARJUAfc
DBy5Rt8BiNuW+zPWgM5ZsjxjfaxVFgh6D6vHtp/1l+iS2yEEX9VC+5Oss4SxvwXA
fZrg9ANZOFH3PFZg3G9bkbJNxIE9/f8Pr9LutkqsGBu2nuSPUBiE8RODwHjOELWr
k7XCAhKchxHp+0AbgI4IbOjwlKqSPlxPU0q9uyYi/jeg4/ouX1HkySPvoRAKewAM
1Z54JHN3rrB3sRvbt3jSE0GVN2hCRrRTkCIdM1H8r1nDMERF7vL9n1UsXESDsbTo
hAIUmeYvyj2K0B0t+dwwkMxDuvbj/lXW6AqovT5Uk/CuD5pvkKL5Q216BBp8CT+c
OEZUKi276jX5lff5THWq5lDiWBZ/uxBoQ70D4mmdj6tkrzrGRNG6dzgEphhzvxsC
hyZgvVlC4lhcaZAbtWoHMapSlvyyRD2w2Dde1glA7M+qZ936yULvbGESO6+UupbQ
D1ziCENR4gY+UF8zWXrkecaylUMEmkq8wHNI+qJpcFG3FOsZ7HCkdNNhcRVNqv+t
75q5xbjCEv9LdTBoZtQLzmGMIANb10qn5bdW8B3X5yxBJDhOiDcj5RUVsQHVI2My
HmlL5YO0xRdKT5nQkl9h7FkF6d50VZnBnEqJDfFcpx4db4WdY44anZSlAQlNkCDA
Gdizxx2/luDot0o7p2nv/ts7aRkYTip49ym2g2kp9YW2dTIx5b9gblUxuREdbj8p
vAH9AquzIf+aorjYQQ3VUO8yBlYDkiSbhpFHTfGYLU9N+He+JKEjX0Oafj/aEdJZ
uP7IFkd+8aI94MZTDC19M9rP5aYybjOEWpIXJjjnL7PZ7crsPRd5b4+u0ALCkP8/
YdmMJ1BVenpfsJ3hysoHh3UCCuFPpFExjRkeVbG1aA26z6zeSzc/GOia7kG0D+qx
4lnu7JCWCMMj9aglSP4NCax+2TUIv8B8PVaknCxTmQ4mARCjISrQSrSTdF1k35ph
NF/ahljSZomMTr2AQ9cKgEAtNTwVhgh3/XqT9YJJWZGMfguQCqZgChp5ZNQCMHwr
PVJ/sl4V7z1zB3TmKmkFFjgfGFaqpnLCw7hZwXq6SIm6XmsoaQSn6XOyniOIkyu4
mec/TUUQ1tBN+w+8DdyxVKVS0xgUtnHOubi4s9cAplPoaEPm9przFx1Ip9akQ/er
a69TFid39OtMo/WpWeR3J2Cyc2avse55RPo/6FP0GUYB8McRIRkC/Xew/phRNHdB
oDbhgVnmX1opDgSh821xaZ6mW2tkhn1vONutbV5xnpnbFTlqdwlCuzmoyLeBgRWu
8oeo6NfzcdJyswOtLfqpcecFCNJF8sBMJyoqJl2AS3QgPhykN7ePMQktFEayWpdQ
3beDJHf3nh/CffDtLN4vUm3p3eGUJtHm3Ob7jI4S+Spa6C0k6UH7h1CUeg9p4x6b
Kt682HRRTkR264vNkLhte9GzS75vNgTuo47FTgidmAoej+mdjrEKBK93mONv6m7r
DzHEj3jSizD6ISUeqXhs4GBCnnunZ6sX3ULf2DNcHNnHu7NGmyhyVjY9r6ziW49R
fefPTNA88xCTPlXkCdyp0a4xLxcSDkwO6ksrSu74au/weK23zbVlqNYoraRkNyIv
ltHyy/BLlMW1mjL7AxQ6tYngW1rSGuJJYBugqOpSXSvGaqJCSV+CYx4LDsqGeGfq
/+pL+4Wc9UeKub3Ocb6po1WxI9LymRnXap8hrXc68HtpGhpBeoRDzvuZEv7jptnW
SR7uP1r+ceS8l8gi6h9YnJN3c0ZiqDc/rw5jwTzPhEQ+uZGrIP2448oxwE+ztryW
2eV2vvczx6BQiwsGmWrCNqKrrPYVu1DJ9cA8nqmmGpsGfXfNEWgHWGzezne/dETH
zypoi3RkLF/ASJbqNDxCQk/TbXuMKkQXlcB1Z8tM80josIU4tv5PY7x5oWz5GnDb
nofs0nr8Y6ILPVEljAc2htI1X96db5BHMsgqK1OsQ3Rz9ovp1qJ+CRaQDJLqC5f3
hQnSyOCqtZGwECRrnLMcZzBLppur2TZmXecZHKND5x9uCft4lsv6b2MS8SabjIGi
q7KEtU8kTCfQtnW9ZiKKFSFcllLJdU8QM5qXGmE0WqItDcXYAzpAtMbKrLJ/08mb
AweatRpfhswGW0NtJx+cY3AeEDytMyMsMs5hCzA3tRu2z94lO1W/mv1YuJMVrMdW
j/y5A+MUTV1wQ1kUgZR0AhsKxqSNn44xv751fgAy4o9DmNXVgQqHUAgyLRwfZQId
CKwbLh19g4q22pa8d2BvbwD1ua9/qrdcUvRt9amCtHeKofdqkRcwo+/+ynqn31VU
QghDT45h/x/KbwMt1sz3PutJL5yb/FZ2RG1rdT8MpMObGmS9u8AjJjU3SRxrlWJq
vncecTyoycRzDjerx85p28vnDHnDJepkwULDTTB7hVvR5TtcIMclY/sAeq+oNu4C
Qq2lKwE5grF453RjOZsBKLTAD1M1klnwVWvHXzdFbBTQbYh7CHcnPNUwrBBWacQ4
OVQMBeqOdLV/gZrp9w6ClbdUT03ZpmQJ9dlqJJQ1V7+D34GtbvSmr4EKE1gn+fgS
mkdv7TT41Eydtaf9vOgl+FoYQEQY7tN/o/kLaaGleNkGBiW/t4sMvDw25WqLz7Kw
aVAsovQYU2Uujj0W0mtvKPZl+NHQdxVTlFfAqLIEhgGYv3StzU/UHBsh6VX2cmIv
EQI6ovhdt8GfrGNHF74Hi1T6S0nziupSos/eD8rOKU++F3u0jEvDD0F4/c/cJbqx
YSUrf3CtId1ReU+j5WUFOCNi/LFC+bBjMqHogZG4y6bRunSOg6AHlONnEf7DIMPt
+x5BEcKT69A+VOs60bz56sVpHEAxj5GIUlmI89WavAOeTL6O0c4cZ0IvJTzrKfMa
61pMaIIZRTJgknrxReIKRDgXPgpzNhPqUBTkV2UxZYkqa3ffVPPFE3wup/n7VaRx
sAhA6GO2N5JTFr/PtgTRkK3LGAE4W56F9OHoxtLn0ZfimFeLmpJD8F48zOvt4tVm
ozh4XxbMRVp6nfSyal35r6Pe2V7c9OUUpUpd/ABbhZEt0U9eGqmQeUXhZfQ1vKid
UeBMLkBmj9O9SY/TxZiqInHb6psFvHxicSBANlrCXSSCu1gMz5TFQ+ymYeVW9hng
+CTo/d4NDxhag15jY1o+SFIbQlIYiRNK8DtHo4teH7sun7lWU/pRZM00THD77DwL
nCCRl48nx85oqbn3TFTJdg01GWXMK0kluRnHTCMU7fbOw9KS/88BbCo3VeMdRXRK
6x5nHTOY/sEsROkbYODt1CMazhWEqxuC3nAedePgB0c0Gr9xYSwmNhqfYAEoP8K7
CBU5RLppxEONVbGEPbnsb994Qk1js2ua3JjdH0fq0b31zpiyprNG3HFtWSgTJfZq
sm/X3Ov8oR+5/H5YTL36ZOv94t6zJOokFOucV20PdXHq3pYozkOp8FTRJNO5mtyV
IfuRj/ar2xswUQO99nFOU7zCxsQLSuHpW5C378YO2uiF1JysAG/xkS+KydAJuVGT
VU8O4l56Xa/PeVjuIoJWgWQ0K03qWjGmyleC04uyL66EoJuI4R38ebhJjc9ZWzvm
luaDr3AeMzdNrkLMOXdxUJc0uW9JqzxZN55+xqM3DcuM8FoEeYM+NYvKn6GkKu1y
rkJuTK960ak7+X0hpJJ70A4VzHhkvPIdiEr1Dae5zZ/JcbLmCPEq5qOE+ga3h21N
r2gpBFBQkAOcyDI6z+CgAMNQSQc1wKu8R74PFCgOtEG0ndQOAo/D5CN7z5VSG0QO
+gwng+ASSVE40wCtkKDsVno0GcFYarRXHsBjCwlHFe4f85SwTsNVpqQ6pC6h1inc
tUnnRjdZnLIf8XtIzZtd6yL6A2MPSb4FmV+5UctiSXGLpaU+q3RAncJq0wVq0rWO
QjCj7ZfuFEVBtUqUgnwellb7grxyj/6cUiFPswDT5175W2ETc4sxlhkoMQDQURRN
cl3Vc+HhzQVhi2oh8TGworoyiHnwdPk0g1Wd5xRdH4sMON4EAJjqhbhXdrmC/7GG
6im0SPCaFp6pjuLID3PksXaa7Qk6spPkpDJVnA8qshpXzy5vNNgib1JeNGfoVRqD
WewUXObTzq7JVeWuwVXOhaGbOBxeSCPFUAZ7WmsgAnf0upcBlo3fQKB2oS7U8hrK
Jo920BODhzNnup37U//fnKFgt6amHuvhaQk0D84wbcTA5YaREhXqrZJXSBzTNc3F
CNEjgZkrVvvnlKVHIZbu2meNul1X4VJl/6ObeC1vz3r8XdzxchcmXeb9yVbmb2YQ
ZmBJ2zGgMmEzyE4odLoo4ec8a+65/VSNFGm6jY4FuCDkSFDo7XeZfj0msbN056Ub
DqgwghmVEY0OWiE7epmQluCMqJaT1P1Ujh1pJRIl2TZS7GA2HxyCB3EVklKdsZJL
360JA87SyqkXDcnfPHQMbtgbnMtrRDFyQKb5hnZG7jonooIvMa+ffAC0AzrY1j8t
PlkLC5/38BCkigrRwSZOUdS1IzxIwxigElZS8eqnUZMPKfm2weKxXbJPW4up5r1D
iFTzSC+Q2H1VY7xzWJX0ElvcIk70MD5UxMxoFjGacqqzCbe5/3ds34mCvX+a9Lgg
yVj+aFMTHsJz5nEyFYwZ29TX6DtfqyXcmzX+Rv7r5MnXQHEsvhxcyTUd5nddmu4s
4rDd9RfKAbc1EPHyUu3tDu+8Ow3xrdgXhDRkN+VBF9DXBM12Ikf44nWb+qOLDSL3
T8YGUseWvgp4J7H69zw5h9HX2JcGeb2Trw4sn+OFeDCjeZCl+ZkDqWwvC7uaDWny
zn1UubAf0/nC9+NXCf2w9dMHfYrZ3aK0yE1ADWDI+f47WchsW8vSgyXDuPhnrD5N
qye0LSQpLvCPc9UIaCUWz18n43zk7WA9dLki3L97VHD9x39FrRg1treO2MImTroP
6k8aQTB25Mj9QhaAk9PUBl8Dw+ATl5K0JCRZUxdGrZMCYvPzmdDBDlK4thQieglF
5vQw3VYyE7HA+n60CsHXEJ5ROEUX/cw5Fae4+IsTy/fHgVWtjSYDozqmC0wQ43/a
QRu2dH90p4LwIL/eBWYcl3JJkHxKVxdGQ0nNC47BRkj6fyreN4Q4btwUh0cc2qUx
5jU+JncfAomFVM5y1vLoBV1luA2kxPIC/6N42AsKznPyM6QlqUi+a6TtiXch4FCR
DB4UXKds1IL8EbbjYlPDdgzvUqx6MigmdHpPm7bEQ9UEotNAZ9rGHGwf5JGCIWuV
23V4Bd3GUPlCOWdE1uqcAtZONmZBrxBZY6V5ecml4H5gB/50YFomWiISY/xWz4m4
UmcI3m+VCdhSCcRmIP+LvLg9n3Hud7L3B0RR77s1YSzj1IY7wmtsqI4g6SHy9us8
VAidotOVUG73MXgnda17ok7bkH/vCuSPEbIxYAiCIagSJmD0giRjRbK9AERIUHQj
oVhFxvvjGu6fMVt0azsFXeWgDc77dpJDQ2G3UYWc2p8F26/oRV0X3wIX8+buDMNs
igNjYl9ca/v7wROZaStZgOYF5mwHdDT8VAouMK4aExGNoISd8QOdKq7zSGTYO8u+
DV0vdnixhP7W2zZhPJQZYNPySoqsaMBLDrm83uwobIQ2MfAbKcIDbCT371LHKQbr
hlLiofL+nhZlOWffoq2aCkD8J1m10wP34ZJev3JZziCJ5eiQR57HA4+Tw20ZUyM7
n8nNNVo6GWnCZg7bItXC8iJXo7ClKHJEaEHm4jbU6SZ3Fjoex2oz4GnFafelL3h+
G4uzYoji5Y1baOJNgbiKIec3ITbnlmMbnRyBeC0tj5um90yVWPXiDavWq1yeQLmv
iNdIx81ZK5TQpoftrQa7QLvvO/y49FZgVB+IPb0jUemS8z4y95VDreXXg+90rESx
ONxa33AbGj/wyJUbcHDMkfgH44I0wi+391/wN+K6i5NnujlyDeIlIOan3b9uIt2j
Wvbe+SSXKReNV4kY9Gf0kxY1AchqZa2ku4ITggINPrnKf+BOPi3RQBR5NWTsNlcK
+dSRhynQZUqPSmZgmRLpYw7cBVqMl98CVP5ZE1QYmMlyil4RYUDC2FpBT24XOV2x
WghlnGIxbP79ds1Sc9ml/becFSUjtjrQurTfvjzsSRBfyRGwwhfV0+RWF0kbtnst
BGIP9D8AZF2JtWZRAXM5uoWhntCZjPjmwBJyO56TfY4Z/2UrBfKp8uOVzC3HUdPm
t4kCkt+M5iqi9RsRvGsx2jGtBG8q+1QFByBEBQ6GHNEElIbRu2qRNqw6affrrsnz
G5oKxta+k6IVnOLWYs7Ys8toqJNZm7tgS1yuzuicvww8b7MWpySP4FN8rVoD3K7V
stU8hlTHWzPcZ4EAKfCTlBVgl8jVgsgMp8EnYDdqghmgRnJHauV8JEPJM4y3AtDt
vmv7bQQQ8q03w6Aa+2fMDL98s6Z5rJJfqyS4Y34Rbx0D2dtWTs3qprQ52bKTBQ4f
l0tk0p8DdCJ/VpuVurzGth+WTlI0aE+5QDUoy3I5qQZGfL2gzYDCOiSwPFjYt2L3
UVi7n5YtxYK45XKvdxgc6I7X9IDJOaxdsxAVFmoIetxOQ17ZhJGGT4L5bkH/UYAs
WukRnOF+9o7V6kOKYfRmP4tPyuBjlt9IU2ZnHmq6eg7BV0A6MZl0h+m3vkKLc43M
hHUwOtDtuHwxH5AFlfRlnl9TzTSP0LnnpWE0hOIRwa4K2oR5IbXV55oBTGoLRIIT
efXkU9+Vls9d3sr/yHvXGUK7zSIU27mut1CY74sIPcmhNSrhvhUj8B8z9CU/Odzd
ROmi9N88MIcBqp2vp7kvFg08gdhZd12jnk7rDXadcOPCtUydFAjmL7b592L5rJdE
Yk3mlIXcEZztRKFwfpBkrieV2ZhWO9Unfyo2L+cza3ehkuh4lgAQmSUrg5C2DEZt
jAIWsbQKJJfgzAB+RjiI/iE5JZWUiXh6K/LTBbWx/6qP0J7dOrUhVbi8SUfsOlsf
vIosJGN/ccj7miPpKCMG20r2wdZ+VmVJ44R67yUbVIeCcqDPF+EPCPsl0URuQv15
tab630NthyGsqYzdMcqds7huS9RdWUSX2XnZbsBRnbS7sWujHvRLpj4EwQZpXx8I
Z/PIx1WXEKrz9ZLMH3nm0PbrHlc6LgkKgR2ipgHMqqxWpNt7lI7rujk5Eql+Frwr
R/ITRRXTr6IXu1A4Anq1HVGNptD2+b4mkhGOAaNKehSErSc8jArQ/e9Yhes0Nmn/
Voq+AsfQcwvIxLM0kWSQuLVw5y1hsaVhNb4DjGChblWulHz/7xWjkAFVHE6cHN7G
PSOgRGXfSH/ledRh/fs1dcgUO77uYQgxKBagbxDge0506CzUSxhNiH0gitnYoJ8/
bbsiaXcBSVwAbufGCPPzCQaaVd9Km4KFzRDOyFaqX4xb95oRc6Js3C3ijNdmx6iL
QES3fq5/IvgpUqUffTMVlPERt8CUOsj/C8awZV84KGQoXadBcGnpE6ju9rcw4uSc
aqQoY2ostYV1fLI+SRJKNtapGkoCnYVw8ljzZ65dhUu8edkpJnuOubNYPc1F3rL0
TjrsdSXb3fF2JBzN3IPe6UzRxeN3TYuPk/7n/8MHeWMR+vDdHu+SsnM+Pg0tqwrJ
K6NKQgUvkS46pOn56B8TQPoswQ0Q0+JvqdFShdVRTzwaCuTF1fHj1CIp5tXxSk62
2DOaTMwIm7W5Axg2Mza5cF9mGYPB2e7u0pWPm52509A0EVtMQYOeluELeAfckFwu
B4PQyWAJ1tPDFDuSGSj1yhxLa73UCUA7Lx1MOLCAvpAFAhUXHjHEzmAFKLywYQgL
WtcvUJLTrZOumeRRQby6SuS7Vho4UwJKIgQRZ904azHmBOGzJXJ4iaEwZBW6q4MZ
M0ttV9U1mCgrZZzVU6zGl57gf0oxNyHkOOlSioAOjhgNCP3K4AepaxUI2PNLBHsi
4Ux3juwPny1ltl7pziq2pCsYARD5+tsJrhy/5xIQUco/iXfopwdgfub3PXLZAUdT
gdfARxMxUCdxb1Z2MIZFWve2RIFoboKwIMiGNlC1Bg4A8HPYcELyxXGo/Vrasj6G
1iW4DlAak+KMRmlvMLTWlKbILdAghyu7kuT39YYzCb+QH5QeBYdTUSEywZ6A0PZe
tBhgLTuT8Ly0QFhhPXHIkxYVlVw77nnc/QUW+8NxR90UzC6KqN/+FTFXS2DbtbBU
FjVv9ApGfdP59IDyeiwAmYYvVrEhn4Jx625vrqQYFb3YRwQTRTI6Xiv559tnQWM3
VW8Iyg4sZlbC2Ja6izRbeMyHvOhwz0vKUztrfvDtolsCy+2EU9Or29UakHEw5MqY
4sVw7uuBuNDN6X+ftQuig5qzwD1el1s4l48XSS6oz0EAYvyAQtbxd8CW99UWFowo
ZoCLw/6AQaqO1itnYd1ssbZv0ofJ32aciwHaV70EZIeB8xcGAWCC/l6UBt+NpTEB
AFNHX3w9tiWvlVGCUT6zDsLynfiA7EJLxH0Jakf755UdaRuROveV/GWW9vvzaFTB
TickHfNizASPfb944vx+SkF3ALHaJ5BkB2EmP1zd4pLd2CFymT49d5xMtMxoRmri
No47qPUgysO3ldyozGLZtXzdv8QjkXLL/b+XDUKOstTh4/iqpDzZtxbtm6Ybbfor
0loim7fcX5V3fwtGTBIeK8RrCk6kwwMYBl2GmkFlfR1cOXW++i5TqjMqfjeQgQ7Q
6rTVzOsC8IyD38sIUL0p+NPCFyoNmkJY6vbz/0qQp5f1NJJbWe4MzI8I2kZzLw6n
Gt7EcSMT5ppFjA4yzrsvEijlIziR/yZJLKZk/BBbwcfzXUJbDPreWEOgOsEdLoGJ
ZbmyqnMCcOGTpKMrekkmPyJ8BydGlcdiKlyONyVZ9WRIPoWtCYHvDYFvCocHVCZp
Oe8v5fXlmABJP8sLuUrEj/wkyZXsikhPIDOQ5xH2gmNHuQ1mQl5zYnXy9Rsxrx+P
C5DVIQVTPltHTC7x3PrmWKx3jUGmdAWwdfVoAP9AZ8WjVqhjTcL100EbmyMn3Z9V
JB/789lQrbPrZjJ3Ru7WKzbkjmgvXAuMXQ/HXqwRYaNK5tk9q96ONv4V+UY75CqK
s1XljRi5aMkoPh4ax2iKMzpacpyZ7PyYoFbxn8OjGaVAqRlOdGy8hPR/tvekVxGv
5wDsPXz/8JV6RjvXmBAgxC7NU2H9zfFmEee5CBZL1mdwCN8XVSPFJGq5Gqh24lt4
BCOGoZrpYaxYXufCZNsGoKVNWOd+ZscmjzR8OX+Onj/FaoU2Jf3beCqg0i7quPed
/N+VXcJUL2OgNy2/XggEGO38G73YteFE+yTOZtsuPHKJHEmMzMNExWSMAQL2BF8Y
I/ulr+BaYRPPWuR1y74Qt/ySiVPlIb0Reg/3s4PXyUzye6uL4IoLdayPCmqiC0JX
7jBac2Vmsy19QJCvTqW4lWEaAKVc1+JnrUR3ptdqQyVdSAxDzyZwl+43VCsFk4be
mccpu01y/zRYgjlFa4CWpLCVM03PlzmgEjqnPsN2RKByZqfkMJ95ox6XMSyDDlNb
sFZ49sTiDU6WVSAy2hKKrv6AdN/UF7Wvj3clodbxyAfmwmd9ncbE6ECGcD5pBgLX
t4K6pl9o/jgtiAd3sSs4qwgEVHOuUEFMCQsConCMLTXLmrOSMQ4txGpy91Q8Npyl
6QQS1rjf/YgTUEZVPPxY2wUCWiEZtI9fMVcisp0MJPFEqChvBTB5ZIlTHZ5z7PPq
PG81Qy27j3n+rwykoGQMqtH/VpY2I4BDtiVo27BfHN+yCSMaPpnxUtCbzIrIh+ut
aJOW7ii4ZuMpN96YcW/Yu6uqqz3TNafuzuuShL7oN7rSi6WcdcJwD1x48okiEHXM
awzcGvndFucm9V3QPt2Zk1Smlh167ZzS2Q8caGLQfNv7eJsI4z3KNlqJplaqdH75
N4MtwY+XpbLcCjd0At8z9Bqfw2en0PthKGEOaGrZNsFvArDP26qr8GD73mkJDN6S
JUoz7zrJtn3yQ0twGpwVjlmEQopGTlODxNpDZvpeFJfgnVoFr0peBiumTrwEhRBK
3C/7O8mWUXOe6SzCKGwfuyru7KdEPpVXFjO3O4q5hqRGUw/q1OYt2lMeuGVfB1Bz
nfLnVfnQ5AIRErote3CUc5UzvIuLh05tXq2jWwIldk8gH9YqB33wxTSF8jSnqxBw
LMMbgAx4t5NqIbM218yZdHoHjd35btZjXbqaRqefCOoRIiOZgQkiNrQ73i3Uf7Tz
E7OcNZBzp2RIMQwzAMdk+Dkai7VO0H3391jH+8xGLfTtFEu9wttJIuk/Jg37drQG
KgQJ8DH6lJLNEptk8W6s0v+/0awS0sXKHsA8nZ9ZWjUaIzlx/pipFJijkLDSlRSa
A6MKjtoDrKE8jX5F+FM2K5CAfjuHZtyYPW7QJaQfFGfjgGlgDirGnDWF6V7FEyCE
1Gj7FSfhQD33SNJk+WOGDe3Bb3mR7Iap5Do8y0wn75+LpQ2bdoDHA3aj5y0AI+nA
nYIg/ohVlJTC+TJMo+GM+SOfHLuuxwpr0RdxBbgLFDPVPzoCXQwwNEoNbIBfn1+Z
pSsNW1anEHLPhOn7IilYCfxV60my5p4npW1OIjJ8541364/NcUKFjZYkWV4ZgRHX
4o6lvdd+eaUNwk4NViFkIQvc6iohmKY21OXU/dMTKsHrne7CRdt0DY0n5vRHZ+Kn
lutkUHZJFzmz45Sgicgm3+xpNXA18S5pmwMaAuuF65MZ18uCKgozVq5bK6og34dW
upScbmZKM+l2p9C+kT5IDyjpHoyWKI3Ut24bEBDt3AUNXWD94DN6fBcRtCIsFuLE
8Rra1FZAcPcdhVx/qZK+Itqfx1bLLKvsrVvMXRL47QpPFbbGHrv59GR6XLxHa+Ob
aMb3A3Rq7a18pt65enA9uQ==
`protect END_PROTECTED
