`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2yyUR65KS4X3b50yFw1Cs8vgsXBy5He8xOGo6xyHdeAtda/KcG3xeuye0Ly0DW6b
XGgJwt4iYM95TRo/nhEeS9hlNgcLsQ1IsUnU0VMC+zwxceJPI7WGuhotnF4srUxM
vr/ygzcaIebOq35OEd94ZfymAH9LVPf1H7JfJLo2yrkIEANtkNR0xLrpgQQr9G0h
6FCW4034MHk5hoxGbyMesdpAamD8W2faAgLAxugMxIp36CBr+WH/8WTEPXAPocAk
++hZ5PBfMfY/FOcL4/5QVmvb04YD8VNBulnb8bIttUv6tKHJSOKgqO9mdITG4gqv
WbFYmT17hMv219wKK5ZeC5ZGwdungFBYa9F8hnyHP7iylHtUWgHXHkXZayAb298U
cpjsIAI7LwT9lmxYAn5kycDBgrf4nvs0dLyQARdDOVk=
`protect END_PROTECTED
