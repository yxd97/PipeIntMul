`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ObSw4DF7Ots87aCnYH74K3gnVwtICbyVpcHntulfiNHkgKvcmtJ48xuV2JdWSt8+
KABsa7DN+KgkmZU87bWYhiInlMrn/3A1rBQajhXGC4BOH4n5VNg76mU6KYx6x+yT
UBMiZFn+6SgwQ+jHfPWFOFyZbSIvbnBywkUS+qY4QfhrYY9YSsfuT6lBo0qDe5NM
Mw1jfdPyP2fsqPk4n+cULvSmQsMojMPHXA8SwgIJZpVi8NaZFnlMuDzD/LYzpa/L
fdd8edx0/KwONWplLM+K3ELjdO/oKoQBrj7a3iL3/4lVT2kiLT5madcwz/o0heOX
IbuBNaPRwxr+6NUyIbUKxg==
`protect END_PROTECTED
