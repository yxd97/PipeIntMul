`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AiDYHAZ15oX9kM5m+j+qO1m8KJQ2E+iiDnjpuIVqW8CXPhB1FYB8U/FSiNWhQRn2
CCe0wbC3u0NR+A9qrOIpRdMy+I1AgDdMhoCiJ0sr8kgNznXKfi6HkAeTm3Of6QP1
ozFJnD6y6K63sWttUhYsmv44IEpG7IqYKf7J8jgrx+iZy0D4Uh4FYMifunYNnnWG
EAyVMvYubwl1svhc8qMQi0sOEeCP4WvMgJNO1Gxe6bloYwnl5NZ0mov3tHU3DkzW
lKFVAvp8L0j4QQ0i2mui8/ENlgY9a9+xhJNqmxjq7tnpt344CCTn49h9u8d8A+Kb
VU4hglh8mniwYl3UEKh1FUiToOCeEyKgoiGUEHcuBEvMJAlJd5VLOGjKmRATJCre
GNDmtsTe+uoVAkNvVCt7GXKA67dxBq08pqnYWiojv+F0BVWovG0/iBWFBsWnDLGG
FC9LNSiWsYhUo/s6n1FpxdQnSdMCrDwQYPGaSYX+qwFGyrpmspFkxxpti5NTy5bc
ZXnHoHjK6KrLX3Lw1HR0yr5uPP5jiF6BwRtPMFDut9uZQwSClF1nrOkrfNQ22RG3
L25TW17dSfLsuCKmfjxWOgY0GgZYl+DbsbgrfM7wmxp+G0X1aSENyTyPVWeCghF2
9+6s7RpAy8FnkjyMhEuhOOdEV7af6WCTFENh6Abk7bKobNJKKf7MxUc0jPKxGOYN
v0avLcymOKJ3qtsadNdv3ZW8l8HOIyrBya00iZ1EJhdPvUDQr65qQYPR7LXyCC8L
8b9HKKHln/xipPORJ5+SpIyeE1NJBUafgiovK4ZsNpqO4YgayecvrPwq2UlG6WC5
peU627cbdGZJoCAJUGLELewAtUwp4MR9kT+eln6O3szorh6y9uzH9J8lkFt4ov5F
kiB2EUXED4GdBlvuO6hc4n5Jk+xsN3WLtho3nb8CjwIYd81p746+mm5LfN11unP6
SK0rVKTK94l9dvDTpXKYwszuPsaZA7BGK/z8K5T4/wk+qTcaeSdElJgN+bGui07j
E0phSwcysaWpOE9kO+YNTU/YmF3mscsP8TvedzZt17s4/Z1Hk3ukn6dP1IxQ3e25
qxe6zIiUQgP1/2mP26iHbBq7fErHIGvJFFEfaHQ7iSwcoZiSJWJLHNPl57giFwU+
9G7gTODN5HIdkQbOqIUPPLmzw2zfF99artWJr0LoIC5Bdu6CtbCE+pYYzmdPKcQK
fU9OMql/EXfxPKbIFGZG/dIJp06YxsuEsuC50Vj0SwmTzeGttN6JY1sf0/CNEIZq
RyQxZMtE59XMHq1ch4+gz8qEKP1Geo0fM5RNWXudQihvW3lvJWxHMQt8LcU1imjh
gBYrfrJR3Wi2v6D/FZxjo0WpMulX6I3D5T+ZHZaB/wi0waV8zqBU6cHRTVmBAudX
dTby8Pc/8ZRmXHUuuCXnFvLcxLXkecrFppHm60kTIVzMC7/3Q89+crWCbbCuJzwK
luKopqSeqWsq9DHFk93mZLmyyycPpinOBUb8tOMz7OB7QNRCtly+XL9fv42sNzF0
EBGuNtLNa14HRHM16Pml9QHKbwG1TB1mOp/leLNWsBnQ9bIgXyd4JidlXtTW/PI4
1gUnNXLvsfEK2xwSoaESdEeilz9UQwmtSqe+wK3t0xzen/EFc9qiD+34MDiOYO/8
5ms0Rw5+gALssOTjc+sQ1Aw50vabbef58YPi36Qefpf5JdZ57GPVrrhj54/wWaFZ
MOBK/igaESfzo06ReEViPgdwPNZsRuT7uGIdnvKaRCwNFUfZnAhDsb/0WjmsApDO
GR28oNWB/A/IENTnedckl/OwxkwfUbOUQpVZTzIQIuBV4cJAfQFJkqVBLsF/Y1SZ
kd9QkZ5ufJQJaP6DHDmjky/5J7ey8yXHwbPl1QGAMFLlgCIhWCx3xbqAb7+bDI8c
ZifLhk4Pi22KrLUM10zqOoAg34xilAfMgyFFQ3jmGNmtez99o8hYH/o0WGxPI2yp
LYZYq9UPHV8GERoG2Rm0TpywW+0UtRMojZ8KB2cUnpAlMzeIS0LASjqmt/L578vZ
GAR8yh56kSWzMAuj077WDZJjERBE1MQpdRTqPry3sBrvzj1UQ+JG2sHV8VnZGaqS
GAj8zE3ozoINfLvfDxdHbZ04htuaxe/PkaMq2A7rjJ5rZAra30H/QH3+1ZDp5dZ6
j+NqSS2P5DGuxwb38zt+Tknpc8RGRZxybUYxVFhiXtOCyf4ijcDA96FMH2xiHdA6
woHQKr5MRPHpxAdGzfzOFvysFrtBuzjW+AFkqQG2oIsfzY6zv86KZlMuUMwaWrWk
nQUQ+qB8yL3yZlFwvMFLAEuUqWTvCdB/ON0oIX4x7IAEtuDTC5uTvbme7mf8vsW1
W5ruYXbIs33vuprw28ku79WDH/P8VJC7LiwhmBj5jzyNpypMPfZsSLeU/khTwxAb
9BLnuHFaoenL3vvmDRR9lGIJae0ZsbJotu6xOBYebwoDu+/8W2SnAeq8NMBQrRAT
zLPJbBzw9GYwZQHjreJAUOLoRwpu9eTkCsrz8XP1a1G39L+96m8V4w8d7bsWSIll
pcSis/+1czn3y1VH4NSy3+6SG5fyDs3OJOKuJBEiFCHRow2AR4yaKQGds3O6W/kj
qg8olWHwo3cym/rFiXmrWIJnGbP8lu0jIz+3T5EDKvaD7XFE3NBgDZJ8kfzKz7hq
5HVVASEEt6k/cq49sybQKGaMFwmZuUGC9XChQZ2nRlJ73EfsvBtbX0X1UUw7cHIT
T2s9H00cfNheA4v4QVeO2IfamYzFNTeQkfKVsRNCCehxJ43Z/DQnLyKuOXsa8k+x
JjCBi0Jr0SwkuXq0QqSnkDwl0/Dx6U/IsjBw11lN0ojZQhsQA1a6XGdoa9H0GtcV
mZASs+9SaU2u+oaEzGqNQ93CTmjBIrLMW5nWYtWZte3tBTqk8NhPuUdJWo3eKtR1
ozOUvqo0Wt0Nfy4VBHkEaE/+CKczvIjjCrzCNgu0ULPcHi4zAkbsEvcmC4j6Hg2K
BmEc77SCI1ZlIs1RnbvKuMf7s6rVpb8BL5O7hKFlG8PzPTqe2q7kMJa3by0MxW70
gDdYKnJzhjQTpumMTlaodWJVPKMT3gKlHNTWgk1C+GkwD24jTLpYY1XSsdbAYdeJ
ie84OWFmNa/6KGJi1H77Y66FZ8LRShpsgUe728kOiqTXioxLrJsXypELiwHtckON
xJ8dKy63wYs/OeLnxRhroqMlKZUR5GYxnLXOtgMaEugG/TKD3Qp8W4JJolGBHFFw
ZG4oK7auQY4HAsKSjhgj6KzvgNwKap8Ej31/a1V24BnaP7NdjH0p8yj30JI873XW
tC8QhmJxL+SmO7a3nNf7Zb6ObGINWxpBjrp9stJblVyX3FnhJ0WYGrv03L+HxmmK
H3fb6Tw0b18sAb6mMYAoFq6VIvQcorGxKgdTQLe4nz3dqVdalz/PCN5sAATOrqoY
lpY3pi9KgoQJv93SYu+iUcDfcS9CX8IbYMiRBQSNt050GukMmv2qCu9ZTLPA/qUc
F0IN0kemKO8tIpSjsm04YcNATzHlLS84aP+YRk6OezQo4X0Hwo1lic4VFss4DuAP
1vlC/exZfL2gasIgHsFiVyiOx7qTCKquDCLuVoQ3FqEU+b3zVB9U8LIcK9MBJW33
10OfGB+ds/mvLY5tD7n8q90sIWUVfLRpdMuZSeugu2ZqUlfSnRKD96FR49KuKYRR
aG/jlxZaJAOnsnXEokWpR2bX3hjl1o78/M+B2GwgQxqhmHfKHwedu1sVsSEU/iX3
OaLQWuq8oC5TgOQh7ovhBCQ6OEl67KLbH02zwRNd6bzMHkgZos0cha9R5aqZAAz3
trwOuUdOMsyGcouP0bh5gv7Lkd/vQooqI5JtmuZBy1JdY8tGv/xrHWGGKgp5gFaR
DD9ufGIBYioQ1o8qtz+d1LxxrOEv4IOnPkdTFv9PbRPt2pP6THIYh08dmn2KzHgL
FarEZn6oE32EF44XfEGKDRwkSJOqKuBaVNNo8Vtn46Q6vrcfMpw/lT4PXmAdqEy2
fjs+U27D93GSnoLKcC02C8Q2/ubbBE5fcuMMnXu3Qmzpnu7lLR0ueN69MUFQlhVw
XJO42CgxNtTOpz1JXkUG+/eeYSg040fO15CK+PNAi9a0C5A+pue/PlwtoNgvPvoz
klicGeb5vQepzFBkycJhtg1H2fhasZFQ21K6kO16goBCmKOexRiad/PMcHMvSb1S
IXcVVY6HYcPS3jM2qdLs3tZD7eiBvOmnwJejitT8EMt65QMwnJnwtHGazB6GaFjF
8bBO+K8Ay6X0Ekl4oTPwlT3IYhwFdE5A2/j7rstmopWs5sSkyqwhxquw86f7YBvc
Pgq67jVRTrS5HR8xuIvmrvbN7XKJ7VbVlC611/3ekzH2ANtpqmPw1Frb3XOg2vr6
s7gzViWLgkYVyKHE2f8XR4r4fSJRuagHJ3KnQkgW9F0x1+5vgMLxUtUUK6WN6/VH
iIrl9nCpGw3Hagp5Is+Vgx9vWVWBV8cGhtvcl7xvevR0juIyqBhqmVe5cUkbYzid
lUWzbP/nxFG8ZsIir/nz2yQvKho2CxhbQXlbG2hRpEDJyQiAGdn4UX8R5+PxL3df
dgdKqwYFd9d1jdPOjyDi1+xzRU4zVqszKr+vHu+xo3E8FsilU2jZxbdvXL6Y/xi+
zrQML8s4Lsm/lYPJ0z43lFcHphCGBdK/5NYyeNAJRgeFkaEhZYXcUSwSyenEWlXh
AAHSC3HR/rWQmV+gwSP/BuznV1yxcdayzxNZc6cPZxUf51kbbdZQmjz+NO+Y5G8j
oHe1c2vXxUZfHXhTAJvJe3Av+B1ScGTOKWD0gQY9APPYAPabk9V3PIamjiut9uby
zNpTOubLmOxs8C4w9y1dD9FqpNVK71mlg80wbfxGrUmvDmOVXczNF49zUELyHX5w
dt/Ivy16F0LQKi3FHQRZLHP6fZQ1w7ZW3/ifisgI2dNvjsvqK3+Jue7SuFQnQ60q
FrtMcqrETM866WHR6cuKAYxJOEnT14QaHddoO+Xof71luVdhHej/FThyWhIFwbYO
1FY6if0EjhGfaH6+Vt6GrjEucKOu4HOJSVeU0LQ9qfT70l4kC20TDyOthpeYPoGQ
Sv+uW2hbch1jjbVNeRj4sBNljOhzCqmqAnGcI5qCT9dflw1UpRLAX0e4Gz8XjWJc
4N+2hrum3iZkOXWwvxCTaCSrTJ8hzbCOkZRVcV/P5EIlcqN8Jb//YQrCWE+oT9TB
XjIVH9Tuaroj487iDvudmyL/I1FMCWgr0HgWZeyIOTKlkP4UcysFejIbeBrlu1hC
7uW9NV/dHClL4dsSl/7ckNax/m56A0MzYiTHs4aoLFn7eVs979cq5QcG8guT8pMD
SWXUij1cresmOfsPrzUVKhnoVet5MPh7Uiw9kKmoO4YNGMV0kDRf90VBMMBCtpfE
3AaR89P320RGfl2A8R15ee9+sdWBVHFiGnMpMdeaJ0LkNQPdxcglrJ25AC3ZAhlL
hQNQRHBns7en797x3q0MrlAQP1m5uNSIfmsZNnkOsWw070cz4CZLF00zV+K4H7s/
wqiDCiTf1AKyVxbTcICdDPJdcsP1iq6AKUtBJ5o4jBXzPdVsBARMl0sYahObnb5f
2HHT4sduPwnu4a9zkkPm8w9GegqP0qsUMFIE5wg+n6l9BYsIiW5UCf0BpGEjwG7+
nEaTyr0xXo9Uye12pveq4MJqfMJdAdUSuMs9xQF86JgddfuXbIonplt+JoNN3v+P
16LiXgvh3I93Fq1nTIed+7akUxeBRp8IxkLMexawKu5q8PUPLCFsPgN2Eprq3z0q
SkG5U9chZWFpAOjOPZ5puTEw9BIQ2kKCZSq+0wO8CH3UvfRLO4EOmIVc3BZbW61X
kiN4vmDU8dn3FtR0sBY8NMb8Z3WzfNBBvNC2tc1LHDFa7890Bffgxujwggn1u2iS
IFmlkzg9YsQ9CrqVuCzopArk+IG056amfmGpkGOSXB9N1ILUR3aZ+7/DO6+5ZzEd
TSxGxYtzyRzha7xxDogmFtA6JGBtq1YO2n3KD3Hh4moH09pplSe+jOOT8idkOaO6
dE2C9eoMQdnEerUF5akojaju9Bbyfl2oJ8p59Q6J08sUqWbY+hhmi9HPF4MMXmIR
qW4zI8Y8poXU04rprSKNYA2t4lvgbkNroMndmxZ/c3roH8Ifhii+OJONIC3x7mKL
1ma0yrLcTUJRmbDP80Q7X/M+SciaNrm+V+a8SyhmMAqQXxPM16WVcTQlwJ1ZV/2Q
pkN513iSC5QBqb4vUUB6g3gtTKyp1xDh5Cps/oWbRdN6ZhZp+E+pn15gXZZxP7EQ
pMeT4+kdud/a+6u8lIfON8TwngZOaGvPrzveFjLaoOizMHQzfKy4QtOWh4vUcLju
/jSrI5GoFBnLOOLNZ6u/iB6cqUSdpzp0fYmrha6BuRJjuEdz1szfBH0ZPNtvf0ov
3EyYi+7PdTHg3v03xe1jZnNOVPXyZm+5D8Re+cXVg7270XTEFj1qcumU80jVqEsw
k0jJpToEzntylWbSmpXbAClG9bpMt6HhRNkgi1Tj6+oVJyFnReuGmxxucSq14tEO
WzxfQ7S3cY9M2+xIllXXxGYMlA3c/BrzOhowU1fAwodolvgp1xUPy5JyxaYLvoUc
ydw0uc2dnP6LbN7E3leLp3sRpBwyloOimW+sPrGGuc0Wrb4OBbF9i0xVCZvJ4T6s
nJlKfdxInOi2y9v3Jg+F1NTIpyiR+k53Lzg26+BF+wTmUBepR5npeVBoQgNAcX6m
DA7SIMQITNMfc45R/Os53zmdKBpeqksp4e7BQ1aX+dFlX01MljcOIiOqR20fUtLv
pGI+QAs+iIlI+0J/K7osqqFXYbu/1cnbCtOUV83bvUXXrzUMjRogQR/SVcswaIG0
fQgfQKoJlV43lA8NTjZEfsXRDBPKicXWtxZEw3qs4hbj2iIOWE0M5VmbhagHN6Kt
SIQr45B04PWEMOkZIPnzDLjSK9npzQKeMyIJObVAuhRezQUG9aTX9FCFYPTXM8nZ
mMEdoICe7+hYoIUYRLcUg7c+jMDy6dv7ZKUU3ELB+j/hMmUdx7a6+tuH1o0i8rbU
JaaqvQ2SnXnq4lrDhVqjtiZBuoc4SQwt1ZBDp4o8O7fx1aM7nCe3AqOQWWP63Z1w
vKz2dVYfUVpmkSsw6LaX3blG7YsliWtNBKgHZUz0+U1DN7ZxstsYu/kvjUEgpPCW
KWcSKGFrp/geOW+tnpTobgkZPDUxaVmYctiMqLzwcyGXBGRKBH0P80sPC9geB/lZ
E+Tnz5u+qLbwjiOQuwWG0Q4VXKb7djJvnShvtSkQ/2yVKr47rbSY+Tk20q+vVOKE
hYVBS9QJgGRa3iKSYF5C52ENe5WDAG457mFk+9gk0v+HrSdQDu/kFwmt2IRAtzgQ
Nq/UMIBegQpq+4m7RGc9rgp7bHouivC2R5hbxb0xkzZSOsbngPCTnva668evFVCE
Dq6Nx9H+5+aqGLEjx5SZWha5qG/NK17JlzxmIvAxXYM0HENeFYGjZ7SAYDxpC3Om
rz4Mp0dSchPMjocDgHXU6HvenE16EjfLTZw8/WKAUL4HMSfUU0NNXPRm6qBI9ccT
Fi72IbDfMrYl/PB7xd0qbN752WWyf6Yl/3b8zdlpokRVHGA4hG9d/S62fvM4CW2i
w+SQ9Y0zb+hArNRrkCCNVYYr7q8apt2IqL0K/ZZK03cjq3/76g0eLgw1xGbuL4/A
4hi2HTxfOQycjQ4cObktf01VLT+y+IlW0Kf5e5fXDo3v6me4DPOxLMabsbQH382+
hG17OHhMa05s09DdHjKKMhkxOv6/ermHiEWOIn9jiGDknzI+iuKN5Nm6QBjoVgce
AlDwj3ZErFZnNZ3a785OE0GzH/pja670JdkM4yWwuxic16iydgt7IWqdIAJCFUls
L1PDua7zwAhuRI43Uqz8BAiHupgnHR9ViM5Sxvdgjo3mltC1f3ux6bBUsZ5bNQI4
abwni/2sf39W0zlQ6OIvCClosi/ntt3zGHAG6B0TKSEuoqYNLL9Ppv6NYP6vswY9
wgcU98h77s+OONOvhpCU+H5xwr9DbySPpEMP8gAUrZkbtGWNjEZoQvFTIHBCfMTh
J45K099ZVfrBe4PzjfYrn4RJDku7oE86zVOa+yuwY1lOOnQkgQ3n45WnXZeA3vSx
iOAZmV6NWlpaqlF9zsoXCgfml4rOQA4EppMnWzFNpr5gGUk2Q4z+A8AEzx9X0oOs
Xz+snEL3ZrL7PPCf+uoDs1d8KrWwYE/VQqKDmgohmfoY1D5zhXQrWyXJ5oDXow9X
/u+aSpC4qDw4OYAkmcihcmy//jEbtiJW8lcrq/fpkPRK4kkrJrzDBDk2jmGszcE2
FL08BngeAJnKo8fXsEtsT5f/LSNVj8hMx2JBEh+VWXgxNlLCGmSdxencGVddJRD7
SaHwXf/lP1yW0u+NHY98gef27v2LFMF2muamjWANJVEUzVoOHGCJ4lmrq8an+Bwl
HtLogiKE244b4xZqTfRAKVV7V0jQoJlEXvAHAwqzvTz0oEhOChARNRr/ZlM4nP0x
uvcD3HfqsvEMNT9hJS5zmx8tQ2EvLr+gMRydgYNO+ls0SRRGdIFS4Doz19VxK4XJ
48gC4Cc3j3ECs7PCx1WrXYcNaH1/UovqWMsTHhZc4wjyww57ypa9azaozmOQaB3H
XIRsAACvshOVoWt5p6Tg5u0krlud+0hVvdmfPi5uhzx+JsO/FN8G6hsEgV8/PyEH
sctq3eosSw3A4v9WVTDSfXWkScxOPmkJHSCTJ3sd9A8DeiEXQ16kepfFw6uNxEH2
jHYHuo3sHvZaMhEUg8u7Rhr/0sy8EWcxlxYVqLAANmd7D+rkNMmJwwkKiQpdg4IC
UT6MH1Ego1UAyI3PupPO3F2ZRQ+ZHwJvQr5M7S0n9Fgm5aKRo9i8/z60qZ3dP/CY
D0BFxbuwTrlXPzH5dU9T4TUcjX/aKcxy3CHrflXl/bpDpdRQ+VWe60Gx2XmjnJXZ
d/62GDjRiCPc2TuYBupts9Qff6bQmoMjIZSjwYDTsNpsNGAL0l5hHPhkQ99qRKfb
Qd5m8phW7oBzc9M0ulWdeIwcc2QHTxY+rC0sjg6EneE9STp/maCVVdjLdLnwN2n3
Aol/gHVVTfYey72O/6KWYR7I8tooRTDVQnW10xm58FwbghrfDVvr9LXvtaDFSW8X
m/8N7xmPwYlSQKA6QL+1mhff5NXGuPLeLWTSu7ZuW9q0xa7soERMBLW0XRPKYh8b
KnM7NMqFjj6sVTHqCMHBxdpW7XZxdlwt+9yvmnKEXSpZQlZjcPaVkN6+bf4WnHGu
sydyGnF3VRNXS/mSIGc/bcIPkGuKOvAxly15lKDE1IuxT8pqFUAQHukftxsVT//K
ler4B90UxDw8r6fQXmAYRvYf8VP22/2cq4OR52/naZ3po0NFZJUsca7A8t26TMkF
bFAV0q2kqt/gx5aZPKEBU+FRVIdA9+RcG8t+nBfoRFySPnutS5b6wu4FNm+med5C
88VjdmYDuHTGBF/RypoitZxjmZWCv9fOCOn8ZglXb7c7Pd4KuBTbBTDHeb/eB+lf
7MOSTjqZSsQjF9rlvWtgscQOPCKTCbHX/onMv2ZGe4IiWajp9YPJh8reBYyfqbss
KpvmesCh9lcj9fLPGdZQLSROl27EMpqsuEVybK0kigbw3r5MgXkbi0RN3G139ANg
ttltHCCwkktiZyl+oG6giFKai9URsE8h4Gvn5CEj6JNF8dJ/INQOOQREo2PxnWog
xwNbuWYpvU07z7ltrk++Y8ygH5JA2dX9OM0edfr8ce0zCVSrlkZKxq2hHl8NHnun
BKYe+XIxqodykqGXtI80QciLYyQ41Eu+kR8qzN/ddbZ++bOKZnTOZd8ajSCL9vlB
grsBaErM27v5lv5E9pAXbYpssKai/m1xofA3fsEHwKj+cnlnrNRqobjHlx55KiFW
CS4xZe+aKbG/+/sdxcYd/ozPH39I27bxKwyduVE9g4gLufRJdLdtHq0XH+f2pis5
uQDYVn4F0uV1uYjcRJZ3abYEyeMIdPxYO5LSuNkO1gK2xhCzhGbjDSN5+A1KDrTH
FVTtFrTZ8resa0uCAWmKXGChoL5SxglHL/eD9ACtMNeqpltDuP4+QY20jT4yKGox
OjjS8Nx8DxMw/cX4zqTXGMQvDHi66rplKn/JZY+vE5UUIyzEPWIghDP9XKd0oHck
JDKs3eRH4WOZP+Auub9Au90Z83cS5VyG5Kz7QP6rhLF/i1Sr2TTBiVHSBWYgrKCc
Kvr3HzcAfwQWoFIINbzHg5BAF6mpWPV5RJxfg0do0ZZi/XP38/nrYVkgCg+2OCwF
Bu0aUz5ltWaMPqwTOw3IUSAZ/mb0KO6nO+08ljyJzf/WJz8gpqZ3Fsm/iZAH4luG
2UNKyQMhHirsGC+xcX/NJaVdfIEluEa5nDaB56hfn4mr74LaCHGh/rrTOe8UiQAW
eYpOYmb28IJhIaCrXJ7NtYPYUpejMkelqaUbrvD2F8NCqK1iMjOBfKwV3ZlZbccR
4YREvxGMRpTn9Iesaf/VCoPT9svlFrYnF5FS5GaX+O7o0WKf6wZngEbFlaknFSAj
AsTqwcfLA+wZpaCVdu6nVqTaEudE/Rl4xcxvpm1qKTlz6FYUqWkoMvZwTKmYKJF7
2PP5zOgO7V8OcEODUSRMfQMfB6okqf5gWIMe9Dcj4gshJIkGscFdI/hGfrWFXzm5
RGGAdyQFP0f+qyHm1CbBMffm8UOkrlnrTqouydrBgcDLuzZ5b1SHS6p2mjpnM2uG
nXnd6VGEf2wCGGryzJkxdnEHl5hy7NzkTVEASypLNRZS/2Rc0bjrnL0mfVZFCqm8
bslxOneTY/uscgvyZidP2nmtBc0WImwEASKYgGzo95vdVOKxiSrLXAw60Ar8E9vh
OwwU05PCvgb3bABypkwIvN9rCDfW9WvLnIS0BfnkMmrtTwI4BFM/Fu5ENW6AsrrZ
xVnCV1a098zR0wxRNXG5YjjPoRwbrxiu4Jr9Y8JAYTGpZl7YLqM7nAgJE3DjQNT0
lrKpb0ejPnWWgetPOlSZvG0HZ8S095bQxJrDUn0ehyMGRK/484cnvuyPXZyUhl1E
idO4w/cAW9EgzmSfGzAQrJjg4QthjraWPePGNLTWa9nEyQARw60+oYmGDZVpDH3/
LSVQHvDcyn1MGP43Ic2D3tuSCM5lVw+bqpSGOa5Z+wJu2rD58UEuSrlvey4c2h7+
f9l3fojgfH33/T7LmsMORA0sO37ZCbx4HB7Rq6au6Nex9jh80yeIWMP1hitIss4Y
PrQ/6MmMsAQi0/GaPteMHk/XOVOMF0GuY0e3R4DNheF+dnO5o78jxYbNqceVMygx
7dKVODgbjGBkB33HzY0xkhhLK1oTrZH4kjsf3c7kqnIiZ3irWSwpy9CZ22g8ijj7
xBtKbIqRIlWc06RR5k68L3Y028R8XCGhqRrvcUFwMXj2W7sv2tSRs6BYaZ9QN8D2
sQHXPPR8ocmnuwS8MrdfbabNJXXXicrRE2EIWeQcz8V7S0iE/HYFSbpoZsQrP5+3
G34GQkOItKP+zUjmgW7LoD547GrxaCPrpv4cTw6cEPdIxK4v7BQq1C6ugUuMqEhn
mjHCrhN4Pgdsx3PQyo9lrX4BKGqYqGmdz5FmJB1gKT9rDJOOCCqM+tBQZY4DarkK
N9ei/zXYnWtIa4j/xzOMp1GMPBPAsU6AzmR0k4WLZf4f9PaR17Wh8B4c83hrRgQf
LZZJApyU2YOetmHmQRTjDKcHPiROGv7cf/RkIiDT6Ja3Ic4rZAHr605bRnH/3oCw
JaJCc7Y0Kyv/rRIK/641Ys65RODbDBNlGYew32rIkVIbxTW06OWVLYKZHkJm/jWk
mr99LQ5tEa6/Pp1367CSVHqsQechEsrk79BFfuMv6LaMzT5GC2xm+67Y59rwcdXs
JMPUR6gHWD9ReF2RwDxPWIPYLuMTOgd57yPU30z/jUXJShTYXLNSSl4JT7O20yQH
Vx1UxXVYprY+k8pITsTW8btG2k934/SdWS4rC5gpZLgyFxBTH8FyKiH2tDMTgUxX
X6K3f4w4WpEmNB/V6qIsXRyY7FDWV1dw+7BlbziEm27ee94Mvo3/8QBh4gVfT7oB
n6RLvX3esX7TpId1qC6pFZzZtVihNuXPL/ykfui2bJsdVD/RreYFnC4jW1MvIWlJ
bgl1rnkygkmIfQTyFWMFPv1vGsc7MQWfCkO64GJA8IzNuEiGc8xfyM09qlNK38Bs
hPdp7ndXiq2RTBcSh2C4MEn7JTI8+mU8uQXHZqjTl+7xBSqscq6WLB7u0sWJNphA
KarSahacjTuLJedy37vmU54z7YNrhV4dWpGuyjHKPJwyP8FJM+QuGGD1o1X2Y9x1
1dw85qZeHyNvf2EYpmhY+k6qugc+bkWrrdmGowtgjzDMSkFc6sDM1sS4fSGTbUi0
X9lmu8yTZqIjl9W49DeMEQCod6oKMaDVGnpqcNAT80RxYuvSfwmhB2pgypYg5GI9
Z8f9Hg7BshFf4NgiAjYdmE1ro2jmbU1nCj8mrh0LZ/qML3K8GApvPq87GmcXX/mV
4+3ymwe2eWObJSIQmHcXmduL09IcZdIILQJwe93a06+IHdw5kSd6ZMsbpHppzb+T
3sEgjL5gtU5rompM5FzM7od04bqIf5ibRNxDU6/mRzPlhA17EEIg4s3KJ/SrBJzG
aguhg+nSQVz7l7DUF2BDFm1fIB41nTWOVwWQGAKU3+1DBWqUpn0x69spiRXwDerL
bFuOWY8gpzX/6W3dtskAHsIL1rp231QbYyM1Pi1DhGrnkQshU/2z75MrD2cMILaV
sheCu6l/b7516O7lc0jjdtFa92KLLhOLroHazKHdf6HBL8FHkzllmm84CUQVnfQ7
4BHrG5px+tToEynfk0Jqdzw72lIDcGkJU28YssiIlJMTxUgMQthHrwfq8c6OLCsG
Lbv22whORmNw7bjmEKMx944KfKMUv3BnT9ryFpmTVRMtY6BSO+b2G11naaIm4Nxf
BxazfI4pXXdd4j+K+k/wothK+ubXaP61LfEk7JYbfXR8sh1lFMkPU5c2WjpoNuoB
cfcm3J4QFBFyWXWmhi7aiP8PoPDnOlL4QqnSidexanMrjjTeaEd4Oja2P76mXEM3
ZZTnP3EgsC6QxD4zNFRb4uQ/Pc8kuVSRKdwgcT7BDpQ7I1/2FaZvA9HbtKCXzEgu
a6l9od+0DBZ9MF5CF5hMr0R/yxzovwm82BNBdJNGkAzjFaeX6y1SOc9sEggMpBzA
eHqcOhvlSEjtBvhuFryD6udO0fDp8u7i3BvL6CK+RPqCNSDPPpf6ff+FeO4FVfeJ
IkuxBImHrxxrLl/YhFy9yLT7zrC57LuacGvhyvTPAnx1FmGXyjjkgua7S+6h8RC+
Qptteyw4/abwgSdTo0OmJW4yQkEFVrBgihc2jDaCEt/Kym/K9yS1JNf/yrEHGY4I
eOsunnLB9GJUBM89Re/CiYwjzfIS2m0lO6bqVWe/51kByWDEqbycQ0ZAZNUywm4L
xaVpc1LbgZfE9udKcXdaJfe2ucyxnDWJnGvBKvTBu5c6pWOn43SSozpGq/V3P2QR
eOsbSJtoNWmvpm06DD98rOXwDD3spNTWYyAQ8eUFaDs=
`protect END_PROTECTED
