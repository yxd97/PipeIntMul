`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TZij3i1+/IcIMMVR1bDMlRYgTEp9hF75QNlsN6/1WchLqsTMTCg73frISwhOqnqx
ZGEasNWKDWPBB9ttZ+e940tgkTOTR1TO0OuF9yTK5vuikaLVWr6BgQDnHHxHSGQM
BTo1+exTJKkY5FtBCmwjv6ttBG1Gzs7dF5hDPnh86KZCD3y8NkP8qQi1OScic3nm
udp1P3d2nvdjPCWCdrft6FCzdtWw+fKIyIjw/hu5TSpfhDNdHAUa935eabl7n+Im
aFk/lnfGzww0+3ZyuAgZisSkMMynOgImQ/MjTWbFdKTOO12c/xoEE/3pFTYmSDa8
ORkPwJqks2zIoYsb6OsUow==
`protect END_PROTECTED
