`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZMA3u1Lgez2nqNQ31VFQ8eH5Y4DOQfOM97EKqg1oZl1fC3zQIZGU4g5V84NZYji
OZx28SlfNblTUhx2y1Q+cCtCRmhbzU3LKYEUuF0uGa/v4T9OInCTIk/+r6VC5LZe
QtCIiRHsRLO6Qrcot+SEUKwxz7Qr8BnQwQpagqMX8ZUDazXQo66PBvb7sUwqcLj6
eb3dqpyolFf/rTu0p4CZmojw+Mk6i74pJ//+ABba9Ob/Ia5wsuD0bCv5BPIHtHve
2eLcDO1EOvWP/BXpP+040laOfwmwfIBcNwemJKfj9Lx6FFWHThM4M/JYuodrKolh
gaKDQy2vlMzygjkjUq6kkej6gHO9x84rJstk7QyKaISHTFl5QhqmyXRq6q/T/f7D
a6sOW3ou6yWVvdRa0ZBI4Hcnf3ru6Qax3/NE/EmpG4Lw22PWf38Txm+eQP320MMK
Ccxc+qnaVfkYn/E/E/HIoXHpvKXXMJbaKnCyEZnutws=
`protect END_PROTECTED
