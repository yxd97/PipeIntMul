`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NXo5wPMzHlevTW6xCfG3AwcGyVILk+xb782gWMAP0bovAn8KbeU1kx6AkpKdv7TY
zGhtZIBU5EpQGQplRQnAQ1IbNy3/LUmWEBNQl7pqyGCxlHwksNRKpwpP6E0a/iYC
gGMrreOkLhbcv8mQGhkbp3yqQTViwWWEpnbe98vFxBGKO5TEH8yQF5HDJJx1Mekz
WjHIUWiT6XQ++cDaDbQX7f+KoyDT2uNufFecY4PL9iVi73gFei9fUo9fU2wfrrxe
4CfbaS1I+wDeOhab2bkttFH++q99aTHgKY5xcspB5MP+U1muAmBaxQO0ojZyxyzs
qwh21jcWIzUWOg0ct72wjdX6PcFCSHAnO7P2WJZgPPI/KfD0C3THTqBQuy4zDUr3
aeNvgXxQF1dSusvEE65RIA==
`protect END_PROTECTED
