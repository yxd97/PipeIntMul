`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Khg7AN/M8lOgyAaY+q0FyTWjjcD527RTkXkJ28KCufxlmXi9CWGpsfLAsDn1kwBD
gX2YxFETuesbg4oQy+u+q3cf5B5ZjJGnGAjBWtdbi7jCarYMLiO5ecCeolBiLCuK
/xkYa5Fx9nbXRTnkceRbt693W5NtJ5REzLJu5l0+h+QTZtMzUCvwJRHqPvOx3VJX
c08aMDVto306DDNL/V66uhTMQVKRiJ5HiS0joT6jPM5sQx/4qNbf2oDKwPQkO8me
wlt3z68wu25UCcoVhha5xg==
`protect END_PROTECTED
