`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NphDRUqFtiavkjFhArqUPmXAKLFeZ0/ncB9zeOxiUzuDgmYNdWBo0qg1oTjBcsO5
+vdOPceFOhMSwaBlHiaMZZ+BBfInwcT/o1kXoMvDpmY3HYLKp3bm20/B6pha7E+E
KGptPSEjbQeC9p1v+/9injiVkYVb/muYf0tVp5e4fQOt74mNKKJwpw0LWAIY/zHJ
Hvq1HORf9lw0AqxMB2ou3duke/xXZAtaP9e7fpuPXr0Q9Sqn0xRLUKDiOLbYWu00
ru9jTjB7iUnwxjZTXK4hNV69LxwvNTZDysXc7KFziHkSgyutQ3IfOx9kfF4Dqzhh
BRQQ8h9yBxl1CleW9ymM341+5m9IUCco71ED36eaYR+LMt+COYBFzFzS4CGLuQ0I
tlWOiBxM0kpbQIGFsCPjcJ/OgzpwiNdTDs9yJ0Tbgcn0jryVAhVNj32WRybIoLdm
lc/vNfyFIGe+vgVX0IMNCRO8kIo1LlaTwiK+4Ogtz0MBGeuZWvVoj14fFo5Wha5k
lQhGnbg6KCcU4JGD8kQ//dhltNkshjTMIPU22qptUArLWyDMAUcAmrtS94INBSGg
VdLs4wxzRteKmeEuu7lsh+DGbXA38Tcydwy0nYJhMqQbP9aknQA4e7jaHVK4S2fz
WdRDiVxPhFQPezEieg8L2PLO1oD1kelcyiv5YLnlHl4TBWRIfVB9cMW8zluqkR7J
0JARYp4PLIXRYioxUcQRudcBmOwJfZbkRVaP4tVsUiuPgTi+U+CFGWC+7iAq9rXz
ECJ0A8xAa+8h3lU/0T4jITX+dDs6NvRw+EEbVHTx3K4Z8E2Wx4kA/TdmFmhCoQYx
IYlk/lA8eUmbfUhC0ehTnqzMnLgnA4JZebMoM63UE5ttFqQ3SOGSkg5KSr3akNFe
C9YpbtzNaXJPq2u3P0Mc9HgsuCGsW6bsKjAh1PoXVX+ZA4TeXrjWfR5oBpAtjRJ0
j8GRijJgSLIayqaH0GJj7Q==
`protect END_PROTECTED
