`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X/CSVDj6MyNto+k3TR+Z8TON7MinZAOWncepW9K4BuMpogKZtpbvTyuq2sIMogBY
YlxRUTLiIRWoRttBmGA6mpDZMNgkBKfpVEKw2Ih8mHA6+edPgRN8eid1eCrrQ7Gi
+W30ef1J2cycrGCGiEDgPTVJWs68QmcW4tgmFo6LE0R/WSQdm7wZgTbGQculsc0p
KZV9nffhU41GyJkWNzsrF9LvFMWA9LYViQZeXQxZQ9a/ziGTZmVJVtcVCOZ5RWNz
xXS1r0PNF+qFUqpSyPCr+brTTC8qsS292aOXGni3cLWaFmTiuF2Dad7sPBxXsBXQ
Bd2foIwu+r653lZCIHSvENYQPfqiXwi+67k86ObXnLkw2vnC4tlfh8NwVcc77IUr
ej503GnXlhfQf95QvwC2t9U3I5IfVtxybYf0VOPmN3/Ln5MXoxGCx07vZUVxfteQ
eFH7pyz90JanGuO7Kr0nDzO+sdoFfXj5OcXhRxVVN6NSgDQ5Z7wlsOguMpW6HWG5
OPfoLJ8tUNLTC/z12Y98rS/4PkwCUByNDYJ4WKt2E29EEjLU6IPGpJ324mpYDYM7
Ul4oPXkkBT0HlASBVhszrYHPnXe3pMjT0lU6wUxnKrTOEd9ODbHdAPQPwnoLWt+P
dd5Z1nRtRxDL9HM7lvejXA==
`protect END_PROTECTED
