`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rV2ZvBt9lFf/C8hLwQL1Nu/Pv380t1yYD8gpOha4t1lcRMdOYg4Vuz8F+tA3fiQ2
2Pe3nQzQAZ84ZZqOan1eGwjyKIe7bU2wE0W7ugl+ZF1xqPlZU2+2wfCaMNXgkwEI
0UykI3lqitnw2XaMvfGa5FpfnGsCJtOoiOk3j+nYYIdDdYWMBPQUVo/+fdyBYik4
EQsCc/im/emwK30pHs48E/FywGyN2dzc8jOkkNGLuCepdAwbpmV6VDQTXm1orzj3
wzFF+4eKlT0aaM23tYK7zSYlrYbJAXCddRQd7t0nYcwquvL3O/Gl7P7tIR2wzZCc
3ZYNtXyejrSxYScEV942gzcYyk1MwbwP2RiZL05/5dn4vHSMoSnuKWcNhMJrq1aM
3yJ1hVaZEmRLgpiyNeuYht/pWvadFXbivmFoQmjOk2YmfgEUzR6aWiwKQDlLT+mR
Wmbd4XmTj87mlKilIBQ6jur0jDorKfPQkMLOtoBmTTgzmJ0syUr/+R5Q232CfaRP
Z3kjLvc3uUog+ZXZwVPd8a2/1ruIUOa6VA0tN1LTXQrRjSlT9zmsqpXWT2D29W8u
jpZhN5ONCaUUQCkLxW+2r2XDpCrOelVCysmAmXckR5UsPuvZFZafZZItoU9wQkMd
JJfVBWiEK4VPe7krAaAR1oK28fskNMGVwL3BZbEorKdlmrwFvaQlM9v3l0DeORe3
CpBygJykVGIwQ1znanJcdciIM5haEBpw135CzbdqXLmITbcsjdj83fQs6un+VXM0
/50yu9SJgrpR1t0j7DV57g0RybCPb8lj70LjVcrHUUeIRNW+HyDnOkwSh/M/Uw2I
cp/YF/+0a93smHmb2hP2YHDB6m380A/nqw4BcF7+SkBpzmhj+blpMdqmiVGlUcCS
VmRoFH25rsig7daC5L/8O6KKyaUKGW2eCJpuwV7ObeXmLPw1oYDojuPY7XLYVGoU
N2edzbWhJf7/EWV0q53Oyv+Un1mPYcAtSB4qtVMpt0HT4kGl0uceuAamQQ6NLIU/
zw4LLNZO+FjEda0XNEANCbzpeaT6FR41stXDbAX/ctpJhMVdYzgvXzB8dHyS0oXT
A6aKoXjIVKZwbeiAUVITiw==
`protect END_PROTECTED
