`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LnUUJnO721RPUWCcVpyLP7J/Un7g7faU/RS1+QRTv/7tr5x+eZGyb2zR2ngdv2fT
aksyVkmPE+/aIP+zJc+u/r0OecZCffRcxhRnEMgjaOxxwpetUkBLMcCL+s9V5yc0
17ivOF6JiE8fxkwOygZpw/1s4Ll/PgQDgsoCiJzfsVP1KN9UJ6iuZjZ+Fr4NvzQr
nKRxguNs7UizxyMF199x53h/95/eqY0ufDM8p8/zuykybCUkCZPlSqnu7spBTr6E
KvxkBPxbJB9pJ3zHkJ8CuHkG2xcD1b1/FF6jKdzqO0UFeqPaX+19la6oBOQBn8aD
0rgbeT2Z/xNQ6Bu+yaXhiioP49sgX1YyEebbImnjxvF5pwoxZqkDTF3DGcOo1Vd2
uogcEMwVBzV0W7q6MkQvUg==
`protect END_PROTECTED
