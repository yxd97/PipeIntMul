`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xevVNIlzKBBZgPx3owxAmQeZY+VXtxT8kncFZmCRAgYe7ZkH6fdLljJANa7J89yB
rLl0DC4YAF4PE+fuEKmVhEiSMxbuL059k3kQjptwArZa0PXb/3FBCK3SgyxZiZRx
ftebavxmv1julDGK2MnI5ruXCBLQIKdbX+RNuIc3ME4vnlzOIvgzdfGG6aNdVbOW
NJ5QjWbQWBDEzvTaJAbQowkPkJunAMkrzAWnhaIWfAAzJFuS8evR9D+LbJN8OYwf
4ALmUjc41qE6ddLh4cFFvgXVi45uGT5edIfLu7hZHiK2DZUKbTxDEkKgyVy3NhUO
BJzkW74cVwtLC4UHvxk1C7jkKcFueIg5hSa6MK/9/acTZiy+Cyr9xB9lXKDKlhHW
xwOweduzb5Q4DCPpPbBNLcAQe3QxP40f7VKtKvP/589coAFoaaO69dggeSFuosh/
gLIVbG3VY7xNYeLUMAtPnoFVphbNDdPrjWs2EapCaiq0/bNKABs+Md4cjO1/3CHX
IZuM1evcLyjX28V32vcLArYSyICvdBQnuhOER/QrjoNpjZgS9bcM0pjTRwPJfMMr
dT6FHzExnO1UmYFxeXXYh+iVfTE4zdmV5Jlggmjq4Z8pnvdq+3DxY39gfG4TbysB
2Xs6xQ1cjv6wucypY/ouPV+LOZ9Z3sBZ1TXnFW/eYr7jT7o1L9B4vgI34UuErN9I
FnggECwmejZWR98sjJJE8oyupruWegU7bVnbUqbbqkfxYljBQ2CTFtfM92fU7Uui
3Ut5Ts03sYR0YNA0gyIcxcF7RHOU0OyifDyp2MDM2O+LeVYnlySrkW+ZRfLQIAhL
O4Sf+Tqd5YqDg+An6tLcnnkLRjJLZw10XdJyIZA3kfXzTj8Rp6fbcM8LmORtrrc1
mL+ekdgzWIXr2N9WUb6gZTXk+AMvMthhCoyBBY0TZCGmnplemzJOxcdjsusHvbMw
`protect END_PROTECTED
