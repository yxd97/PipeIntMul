`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CTst00f/Brlaj0AC9/nNQc1m0ISFpbjGzI1f4KwDswiJiMU9JdPtn8ytWivNYB+6
2ingbppuxqf5UnD5W5VFrzLcEXzKxbDmPPEnVYgMSCorhtNeeCPdd6++7rlZsRHY
triURVYZGxv5ZAHpH39sGXXvh/FGPpprm7Ark+NooBzMCTsVoWgJ2XQZxrsUNILa
XcJmB7oU/SdbP3/kpyCuupFQZkMmAE9OHwf8lQ/FlQYJlBNxx/1Q8ZMrx82FOr4/
vy5lPPeSfRQGSQqqHaPel01xQoCvf72y61a8O9J4sZ7jr0VWyBa0FGcehceXm5iO
E1ARnB7ZNpiNvZd8s6Z5F0Ruru508mJIQaYpmeWr0wSzT7jPtkZvoU8g82cX9H7s
PpPoYOk2Kj71uYSZnkgGGmcQyYfbooW7S/IC1vmVOgM4yAM9R1fZa9ripvNVYeZC
yemKTSIPvKRqJogUDgM5brp+sACdHxtF1c/T/uyRJED6wGaHsPnz6FMsOrM6a3SH
yBK3EVQK9YrCJtb4ApsqD3t2vS8T0VEa8IfqO2sLjOjnK87l31Zd8WgtItOPfDY+
xbbQhjqeYHc5YaIfkHS5zxPg0IkAuREoPhpnbK+hFbFxYTi1GiZHBex88K0VETsG
uTLp/pRhY9QpBRQnm9xFrHhCxMpdEZ7cYpU96ZvT6GJTiqTDUwcfyoROrmtmhiGZ
K86v6VdnknKO9nyHms/twkx93SriXBmUkFNMz0EkMBvqk+GsXVLjwlC2XNlqqdOW
sVnuxk6oL+PAnM/TdDcwekcx2qzaO/9RGP0lj8fFmhLXf4q5fRoNrKZe5va4SVo4
XX/65XODe8wSeO5+1Zc6i7qIO6rWh7fW7wkVg/L2wSVlYN0IvtCZ9xvuku05txoi
mbSS/5oEhaEZSiZ6Rawb/sbJ5AfqFQ4UA48GZ9tj7q7LQE+qZBWJKCqZFkdGUNde
L1wf/pe5u5OjWOmLIgpDC1rPj39zZBOeRq/hNX974+e3gAso9bBNDL3lZdiifIXI
o7iDjY1Vb2rO5Cw9tx3XwBUG4zbjfdPe5vCec0BGDr0NU0B//soiHAUEtIifXXFe
q6TbmsZwCV4L7/t8joU9/08EpwrAjeF2G/Peza/uOEulVlbwQr5T1CFsH4wXGQVC
RRlRz6a81rzsTAkLV0SIq0I7HKxhInySD5EtBC2327K96VG1/EdNSLISdjZMEbmC
Nr+oyFUxqjHaydjbqkjdta2M1IcRc/QLTGiLxyV7PF4FdMoFRwo8dmB19sAXa1l7
wfUqlZWklAgI8R22eNI1qvW+j6mJs+evwlZIOh2U9fKTNunP47bexKbzULHfG+Oz
zfLZomJCCiwwPUCvrQOO0DOrwLAJIzqZTtkDSlPoaXT8t0H7iWPPZ3kRxFf4WQGQ
UdvJRD8H/kpFEUot1uvDg117hYT4d5rIpp9PyvINWG9q6KqhrkPR/stVk+fBmQaY
IjvKIXYObZUnwJ4nHlezntUyzAwrdXj0XU9Qoi+jAzc5RZ/MDaNEqBYzANggzHtD
1H5uddpKSxsOiNSNQDkxbMgUa6cEDgXjOBMX2eLxOi8NNFpIqndSP9J8cWj69wpM
+iOkd2CCIBPWHtMBSYrRimGrROEP3mj+o5w4o1aJ4clxQwoYHT7b7p8RuQawoJZH
tnxgcMmAImyrI1q6o+Gd1E68n69EnIdTooIELhqoVVn8pP6sNslWEpPdx9PXdJtQ
8foiZrHjbnGkbh5Rvwys3Xsn4t7HSdUbe3op/GcdxugsLl3vAuXpJFK6hsrByBoH
x1lvB+OLJl1kBDd1iS2DVLPLakZcLhTyW5G+PgN3t85yIS4wdcUMTNO2T6fysrzO
mck7HsEejsccBJWsqGGQic2IwmOIyKRgH/U7IcJ38acpWGj3u8WMiGNO920AD5IH
ojZAz8mCfNgVfnywGieq6BN0obGa6Jmi0nHFhIeTG/irW3WdmlA/qyCZvdyoV4BB
FbkJKb3QhwEVWBCNrkDayf/bBJJQctHPqhHpzhjd7CmS8b2e+hqAjVHNqFpVWMGm
hj1D5vDJ9cCm7qYKY+KPXt0tINtK6gA2FOHTo3iO3j2c9UgMibBnvGK+bY61YpF0
bVVGUTBAWR0tWkJBs+BQpoZFA27nYrChtDrKdVOHNgHJZai3lkJqaoqjc8Q0jpHn
2mQWcubdgV5LRfo5MWeSqcHWeY0C7Fyn9FO60snnhDPYK46TvasjGMW9d26uRtT7
yROQPzk0OkPJvUtoCRLigVSrYV5rOXfllOPyjTij6Xwn7BVcqRoI9m1IL6pZhGvK
trWPjQaAXOp/TpaCd/YC6sjlBzANrecQbXPHKqnqNVkKcIkM1khVGGw3AzG8+S0h
mtMmbkxz6FkCugfa8oFu1fzemhKoff2h/wNcxmFc7ocvnwIw16ElDOZnfuIbyomL
lCLA/rC424po1iKqyU7a+3+wsGNpKJZiz+g0WASmZ2gIFce2+CzaNxjTa7V8twLF
YJSoWW1H9g6DMgIU2PM//dykbCspKp6hwhuxWj0VewzykdDCiZS/QAbwpfDnTENh
2YVl/iY+96APfEan9uzV9IKqPvQfr0P6GQx6qElvEiL5D+CoB4X+wJy9sWdpPW/P
sPpkZmLqfNA+FZK4N8pj8wx4AHFJ+7knRuE3D4RGo4wGgnZBRuaVSJ887kVer+pZ
OpEWV/4iCQFYf0CNa7cVDEgrRIDf2L+n29NQcJCFYmrdd9r1STiiCDfYHdwaTUv4
7P7fjCjE4Jw6E7i6tO/BvCqFcBf4rqpOSWUZPy98Fd21w1cJ4OBhxK6hxkUZ6CqP
ivmq4cNmYny3Mix/iuJe9QjxgVon5GhUmwQti91o8DkDRnGz/OapkrsDmDutLge+
bTJFOAplctxEKvmCFTZZwPXanqQISe4L7ucq7vL/+Qupg7pRusyMaiHUQ7WMS70w
eWdcZEN7laNnVzdvuJ/pIj5KCryqZgXkATo4pdBSMro39DyAwRA0NgpFd1vKkCyf
R83JCthwXDUOh7LCRyQwWdOj2GR++GaM8VqlDj/befyAsUyysYY8E6WaGjrqHHJ5
zToi7H5JwOBRm81HoiOc2h8BaXKoQ6bW9u+QfBnykyPLTDK7MjvSHceCWFDuKboO
a+lgZUC3Ikq12/xvHjCaIXeC8aWKapkzv2HVZq153Cdy8jy7Ze+Gk7lpTislogkK
rBdPDM0zHN4lykDw6KIjmC9wQQ0OBlbj2o7I5H47B815O3lG6xmfFDZxZBye1hZu
FAPsTOk8rnYX8+kHvjP+yvshnWzsBMClcJN23aTIKikqp/DOGnAjbaT8REV5X6A6
Gvca/dTGIeRRvFTYAfY73qFdAadyA16NU4LQ+i4bHF/cWdEyeh8XqMR+aPP9EJBO
oPecuW5RsviMA7WuEcZwdEm+YWpT/5jTvA7RuZfU9FI6mTu6eVJKawdJPju/Vht0
+f2rZJ5pgRAcEmYs8P/NWnDbBhNAv1B13b9ADdWvLGHasZG8zqckKZrcRwmT8ibJ
s8Kg25uEG9nczS2K2nxvc3uAWrbppbkPun4ksKl2KBEDdjy+l4vd6P5I9+zwSOeE
xRUBSbOjtarhgc2GOpupiEd1FpGq7l6LuswCNsHUSMBDzK98tAyghcLEP5YiICF8
/Oqt9x5VqkCPu38rBjfUiXkiCnwhXPq3YGIO6zW1I901y/Gvej4EotsLJvXKiVTB
zfcRCoHBCdRamerH4N5JzFbiD6ROLZA5ZwMYFlJSd+BfA6D3lcKI8q8Fy0KYyazM
ZHH5jPcr7AJUZEBFwBRbRUZ/zkq7L/wO0PN/KD7dr+ul9mPucI+QXPmrmb1nMNV0
v0iIZZansSRIS2WQh6TSDO6NKl1ZEeL0UNrHw3Fd20E6pbOGS97CqiALxKxLXZzc
6mcbUcs5KhlnqlcCfLe1refQZTfidR7wS4WrwRlzR3wV47xNS7nytuHI67Z03bG2
Rjm6a7ktJyEAaYBAx0e5AhGf8ZSSSkJCWWZ/6Sbig+Pv5BTXh4rcendDaVqTwpD0
bGVOR//31BU9m1BU2VU+ydE2NP9J9Fj7P+wtPZQPKkbSTyGGb76mKvw7N2rx7WQS
eqQzgz6QVEDEkw1sGZheUObQyY6YQwy0jZ6FL/ypO0PwNU0FisnvlTmz/MZG5/vq
c/X8lTsoO8mgByh2fsyYhHyED3kUR5zoQPtrBP4JX++N7O+V2CMwa/Zrn19QgeXC
C3KLQboiy1T/Uq4kKMPqVFiw8jNIfxJdpCoDn43z8nAnLzKxyC1jYCcH2a0h32FW
o4CCFPjClaY5KcRedpkHQPFggYFeHCeK63AxCJNNCu1O1+gwdzNUDPS6elmWfZ+L
t6wfHctCHdif/Faj3BxzUEcKWMBzNc7yevyOZt/Fd1SL0kn4S4fxOf96VEt0m4Id
yoxfCkRijXzWrJBFg3ay7wxRfUSvqqnTbsLltgUpTIuBdCGOyjk60CJSh3/59kkB
rqVUGVctImjhCEq/1spBudG85NYL1Z2biDNesNLIFM+eeVIB/2BLf1e/M8rach0E
hfZJbaRKQpfIJhLwTARxBlMN39auBoRSDgyQulDlCuhUq8kEFQ0cvksAUSl6/zsn
+dTnvOs1rpX8qVBUxJU2kyBreTHst5zrUYLbtUuYHBEzE2W9/u62K8LzpvPyjyUh
Y9JtEPz/TEwZM2TgGVivnxe9op84/a4rmGCQAGnyxO3Qu15WW7gjg0RNpkH1aojh
nH4ftK/TESKR8QD6GwcHrokLtkLmLewd8U37VADsK2Kh+7EEqnKipaWodLTK4mdO
SP6rU+rQsrNSz879V8j7nPFcUAW+PsggHl3F+vXgapC9VFAg3lIZgasm0X3O+8oQ
JChcp7jtXVDTt63R3thaniSg8CvcDdFglb+dxJd8Y5SOuF7V57MQNE+Oz8fJgd7Y
`protect END_PROTECTED
