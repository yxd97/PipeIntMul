`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ekgeq25rm0J3NEG/QwCj+YgcOcYa++CC44sDywq20HepgHpdj6YXr5iApE65EI25
wS3mkxTrxC+/kD+OS3YCOSuZz0HHbopx8DMo/EKOYtUsJism1QVJTngiP+7k71rV
gdECbiBm1OPG+rC6LN/toczVJN8nv/2PYdZD/tzbCsA01c1oQiFCR/viBpvwPlnp
kMg0VSYFcTs2X6RwyrRiszny3a1DbqaGrQtoy3sPRXn35QZj6PgbxtFmsa+laBOo
6Die/CkYbbjoHspM4HlF8KkpYV+jH0x4fWG/cY6Ar+qB+wGXagTIujadYTUXzIQ4
IbUXcg7XET/4tGRnEYxTtFbT82Bv2Ge6m2FVJK8qSDmtfeVAmHbeoO46HegMF1qH
TFJ2Nls/q9Jev9lWYfGQYoz8FnyVSGaSRCkPZQTtk1Vrq4sXvbV2FmN3qJNPZb3C
xCIZIzWhK+WE8JvRv76Hre0aXXGdZwZhuqGD/8AANTPpIsf+MAjuI+AUHkZfyr0O
`protect END_PROTECTED
