`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HV3DvlaT5l0HlIXams5GDjNmUfsQKC1LKcoxTf2cJiv9PERVis9GBCObVyxOP88T
Yb0j6GBF3T2+7xCUJWJe2LVq0GIXh/S7ND2AQ4VeDRw4P+enOBlmS5C69IgVbWlF
MHaEWLIQ7NkHWRL/OKW+kKZSQMcWY3HkB6sMXalGNzzDPqhOf3rB2XhQ/Mu22qYA
45igYTCjYAoMX4y8zc9F6H5VhFaomJKW/USa9hx/5dVHXdZG/cNzowPyyblijuiv
WEYufbGi/HIt6djj4GBSj5PWifJ/iAj/tz+2PhHlk+X0dhuKn7bIAHAB8tXmA3GV
7jB5CB9r88+GI+YKroDF3iMYlIUjTw8BmVylRqughN2nALjdkP8JghJmvTrHmbiU
1R4nxdznFW95yUyTfIOSFgx+NK6nBKiWI435WyHEVhAsHg6iUWtkg0/MlprR1Rhb
ao0QEcAZXzoNIKJSLxtLBhTgJzmOTyuAVIg2ZL7y/zWWwI9DQv88ACFrZejRBDuz
kLJaB1jYwCXNn5jYTqQ64Yqp8P/4WGtwLNqLF89hmELQ5onpiRLXV2fCyFmblrps
vPIGcRqEOHerDoWCP8tt+U2OfBifD+UqyBBUbyel9YuiMpUWxBlE3sOH8tLHL1jv
KcPK0ySMaWTdlpdA2TL0iOcOOc7euHKWGISPXkQnjhZeIzRD0BBrvUsDgh+gSRzg
JeepkEoJCVCSXR5lyE4r3WuA4T9U1IeYTer36QzOA7jL5qUz0QCpcgSb5Yzy4Unt
45Ej2x1F5v+vHSjxk/Yd5AiJS3J9YCNyyjfaboSJefEEyOSawPeFyxVmQ8A9gAgt
SpPSlSF4z9uaZLXKDeO6mhUxR/RXdjBoXXdtwIf1N9/x7sIEkG++Oxpfc+FSnxfD
9c2QxAjdcqrb2mItsMg371tL0K0QMcFmdYiNDteKhMfBGpLCB6X2R1kCV4/Bgdbv
yXy42UzY5EQ1QN6hsD9ofAcixxJnHOYqsaSHMk5IvZx7zCrc/TNsy8Kq7C49gxXY
YbcSoelc7EBHQ+5zYUZKmim12jizezjrW5Cgw7JnP/IdmX2ofCYarMVu7FhrWVzL
MtGUi97mTmcra8Y7Eyxm0z0w5GtviM26h+/mekk1DHSRUx3P5IcL28bpqALE4E3H
GYGdoX2G5B5Z8xcmRnMYBeCiPkaE11vVG0zu/t5JGMwSetRC/pDQZnoVlCX63IrB
st/tzBBK3VV5yrAlTNGmvA==
`protect END_PROTECTED
