`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RpR2UKbdsZnHNsELJJ1V2Gp/FKziqUcHnvLxenpcCMqLKSvJQB6rBwstUg0uizB6
//6oUpCyTMk9hhvVX8xlDkFSpynASHEMQ9AZ+rFGkofmXvncPMIMSbPgYPL6iXq9
n6hb17aBFeSm3YrEHuPUBMT6aSeYXbvoc+XkO7fRk9webnVhkx9lmCW4l1tfayL2
+4OfjWrUoFREcRvDn/NxI3VUxqSbmX2zb/C6kmOu0mzZCi+8xREWKLHK3RJaCnOL
ImFP4YE9UqQbPV1e8uaeZ33Oi442HXYf/gtv+G2M2FASkjRHGI4bbFYlOTBxPOSl
FRBhA9TGARu2ta50XFMYhTiM9xcQfvezspjPViTtoim3cdRtEBKxVFEiYbVaAXMS
LfOMMUWRoE2XZ5cSvcfSWqXaiY/Tde/kjGvvconqpuZu0gQTcD5BtQts9/YeRU14
6zhpfShHDLY84X/3/X33jyrvAuoPwaayxh4DWasf06MfejmZZUyK0S8av9pKEQF0
gjfJsreVvt8cutasK27jqgb9AalLZCsq6C4Ij73FvzY2ELUkn+e8xB4ZX1UKe6mB
Hjb8uIm8v2UcBMh/1DJHZGT+TKuHX2nNboOacxGt+XfGBDfZljVDurrPHw3CotBG
xyeKTGilxPvDeTF76Q2VdoX+EOxyy15d6t6e7RiHOAeBEtEHVxg6iHK5IpCMSJzw
tXw0LfxVayrID9gCv1wJQV0zileQs0xceiGhf9gRbWsc3L43Lo30q9ZFumlfGvSk
CDD/U2xheyUI1RLzYpjtJ7OHupWABorXE4+5aDKgq3ZVTcUr8ec/rL0t0X2g+Ugp
z0UEP8DFECGLI9U8KAWlUbe0Dsjry1m0P208TjvhpAU8o/JrXOdEKmCigmF10Jb2
VWUt30VvTlA4RANdae/Vu5eop3+E6UeCX3Z/DM51ZlUtTGiJDShoGKrIWa7PtI64
Ue119o/MsZhunIdRgl3jw1QOK4ZZFrik0lNMqOOwTmF3EtWfEqOwVM6Z3tFaYNiU
9MgQzY1Kg0xkMQSAJJ7SAgN71/5594EVdojbE12jrBpNEyLB8LPIrtCoOon/7Ok8
HWKnO0uuvOiy2k/4y012/NE6fl3lRWEseEKvHgqpaWh7oGcOz00h78nPC2elTMxA
OvYpXmKXsjGR+QaCGonYZhPMsz6in+LqHlZtelocV5bhpHuJROUmyf9P7T+6+BOj
2Sb+C1uBsMMhuQgpw1J13OBkLrp/qrVJXB9Rsy8qiExYs+M/HtqCNCiPJ+ZrPKal
u+mFwqYupTo+JGxQ4xQ2M05+UHM+BXAagKWviO35Q+KGKOiG5zX1dbeXhFrIQ3h+
vVQ3zAg597alkwQnWRFkiogBOlSpNFC1ViGziIbaiN3x0/9qtKHn6S7I8Ts8Es+j
FOV2qbhMccWeFtjSFwPjZZsOZoCF6dP/g6PNAL1F030lbUyTBw+q5f0/AHJyTC9X
oLyjxscqEb5r0EWp3Jmf2/GrgnEJ5CfckShzxnzIXBds/hzso2s4ZCwyC9wpYv4c
Gs2N/hW6+5/6GZgd3DnbrIeXx5Mrdx2cReImgmPKtvZqrO8oH/3w5rRvRVarWyh5
NKcYdyobmBugSHSxSGhXu4EXx0WFm3QQKcqbsHJMp9T64DVTBqjhmnWKUelCVaVZ
7ZMSx2bVXuwSIEFm1KEKjvZX0cjk9CWDovtrDKccI2lLUf3IXkBf543KNWk1K4gY
4oDesBVeuXvitdbn//7vcWcGNBB033Dp+HrKIMONr4yLweX1x+eUFVNgIE4x1JxG
mT1L1/etMM9wXie8V3zH1SVVx8C54IiGFHh+hz2hGYOYJuJaIe5xPVRlfPMSOQuo
n8t+uHjpDnKJWWIQpn8zN98TuLIX7yHl1QYgV3C9C6O1y+dVbVYDuqDUx3Z+mQjK
QckDYbQPkum4jWwUMHZvb2Zl+5ZiUy+nuoDI4/gtNHjY/3z7WXcOY06zsiPz6BeD
76A9wNcHZDY59VTodvchlH8shgwqsbdltIrhV+rBDwYdE7bSfOKogfdeWupMdfkz
fsd//gXYlzwevKmR4BiiMkI6Gahzj7mDpX8n2WJcjuyvAcKNR3qpT08jfsaAR6xW
0HZ8W8H/AFVqBzkwK5W+a0r3Sdzbu/K4RW374cXbbL7KjcmAQYTmhNumbRONrVEP
NfVALhzgHBmDqg2J9zB3pHc+wWXW4heY8k5r8poVpZPt2ozJJi5ztjEWaMptffm9
A0nGxi9MqTTYr7v3hAbelz6NPlGiagjAdwWpCiTeOrXU/Ff0dyaFTJuZT+9IgPZA
s21GSXF+/4n3C2LZo0kD7Q+cPJTP9TWeYq5xYcCrTjS6ixHj3c42iZGQiyq4ny8e
mStij0oBHVPldmY/RMSaDBjCCCrlhCGxMHHrRV39/Z33p6AQSIWzQC4ybc/Cwgzd
1dx6RaytQ03IthC6ov3LmnNQfNID2y8aSPI6TNO9GnpmT+eve6caD6gKTtQZ4Dat
a5c5nitFGX1hN+Z5DHwNWUyAEZsnm1j72ttYBHNXctW9nq+kdDORaMhnz00JhIW6
0D7Wj/Dy2fWZE+PtKBZLSxs4wtzE567vWOVjh3lSV2JqEXfxNqnjAA6wQavNRbCY
6fJ+ldgVsiZtLuicTUXm9F5alaQBNyeDLntuXsjJZMG1h+HwIjB8xtoPf6qQaLPI
QDfCeX0y3VHKXP1No0r+eIHkXo6YyVvwxhMLXlT+XZjtJPTbmp6fCEm2ViGNp57w
XClK9qJZIWufczUAH9jzNjhYdTyaI+HCWV9V3t9nnCzc1LrHE4oaV3MVw24ggI0S
0cJ1ge/bBwk/HG/jPx7nqA3c8rrLGPUidslAsjoD+GkSzQMglvP1LJGbPBcpb2TV
eqJXTYdT+pM8uHRx+iGTg+ngovS/hcUcyBa+uhzFp+nN1Oqgf2GEZCDv1cYOWtnu
YYSsdUCiqyHSnyDzufrJjg4IZVhcJKTNRaqxvWGcvZ/Lu5YMEJf+DzBuEfaGVoLs
iPyptDwN81K4VLLuXDki5whNVOzdCD+2ZbWa6LqbT+nhDg5Moxx/aieokAUvKSBp
iy80PvkaOqATKrGjZFDC97le9ogVog+wBEsC++yBJHuj5OtXKLXTrW4EhkwkTjD8
HvhgwdcHiDnk4mZVOo53kdf/GFxpJ2sBGoZDICd7yUYn6yIyZlehztFBw+KczXkd
Gv0qmXiY1PuxGj89u+qLZXr1w3VGw3Sc7nIwbwJ5DVlJIcSn2oaBcL8qM7xAFx1w
IGpXT++98Mc903x6otAB/FfTD0qmUra+CHFjt8cRMx68sM0YT4XEBN++1acRycVW
zENxcmUM/HjLchXgHqgw1Q4IAvxSUnpn1YEnQCKfuGmyMowxzttARkYoWFvAIZ9e
I8WTs2OBrWUgO5UAOud6Kgz0ds9Vc+zlcDINudEjk6+zhtcHt8jqhUH3Ux5odKIH
RlBYE0o5fKSyK30dR6lrlaFkib1Gt7rtLdRCjI8d0SX5LLF4ZBBribrGfCtCEd38
tHkGWAvOwapvAefs0oVs4oo1y/XpnrJagPV7+QeX++3+Laxm+avlDbpbR2dLTcgq
0yP1+GTUMI+A4mSrAAYXtKsl1Poeijr3ck25qsBkarvuNZ0en+PYbA3SmVnrZ9js
y3Ibl/zh9LBD8yydbhfjqdKq19ktnO3ZNg1vND58ZeCeY7lDAPJLn+iv1UCe0FWM
P6KK7e3D+3JvJGFCTegcOQCjxV1Fwxik1/aHrz/dY3ENxvpyPQzRSsuHSl/vdhjk
3rcLlNLs2swjFswk9QLaNALKlNNPqpKANXTbLkrP9UoPtsm3Fjk9JDgxWAEeitdx
U9mQAbS2tyaCimQBTewX3xYC4NK+fJW9HLSP6LEtQUeh3whK+Lyo1mopc4VP61UG
lqC6Q2CyFk8NFJHB7jYwlM7qhSYdGMQReI3OynWnUlgvldpv6fnpCPdgLOBMY70M
1qIZ7WCsmWtxbqmTBwAGsZcuR+MasirxVdQM1t1yvizrahE35owklwhkt3SADGyx
6pfPsW5EQCAf3vT2sYTgvB596H0UDZrjBSs7Ln8QqafeEXTIMOM/3dLmgnKip9PT
kqvMcqd1NXyM6wAxRhnAc2e3KrP4NVIhrjpoBXYvwbgntgbXa/a7u6o2Q7JOvk1e
BoRRBjhvGyCAWHeWVwkKLEwRoVWeaAW9rVeYNpryP8gcWPPq7yhGKkcDgbKe9rnl
q2TZvsH6Lgf3E56zZ3pOSbqREEcKUYfXuube5gwNmkM/TKMBtAKuq5+VhNL+Yt9f
Lu4KxX3eUYccZ/RjR+PGWHE5hYp/OkrV7pIGqGDtUklelqV19gUzjSNtjcCiXwsQ
fgzpSIG89t7EgzvdweW6IOrxfmOdsKdSiD3AgykJhxIVPUW+JGS1hx9tWRYWcM3w
joUKCk8sxkGWPreN94AsNQ==
`protect END_PROTECTED
