`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbVhCgcxtArXXt1HlS55dcBxxGX3g7HQkWGORX2eH6e6V7k7Q0DjFz3viAE7rJOH
9uPMmdq1OaStwgR5qvTXPr+lcOM4yVcT29thMK/0XE/Z/25DyXO24O+jRzoO3U0I
O3M8naC0ZDY8pQNjTfJmbFm1gMJaPxKCow5VkPfPANiRq4xgLGiNOy7pNYl8eM5m
T+eaXJ+kTLtbqaSvRPPR1E9kOqI1yuOuM6wvr352Ia3BQ5Anw+rxmgNpJvmsuvnN
j9DCOEiKwBwKe8D0SwMBxXxbymdjpO4WT6moNETJO5d4JQrOxXe5Lsb/w190jecC
ihJQ8p1RhPGjKh3iTkuGcj/+BRobkL9ymMVytCwWf6CaI2+faPFB1f3pIpKXzJUm
tHTWVd021iKUpLk3oHVQeaj7Xg9fHm1hf5IqE9nhntM=
`protect END_PROTECTED
