`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u7ygyN/iXzQWYGrTMeVXjeO9orgYd1UGDCem6S8HKZba/ggPLXlwra5sLVb886/j
O2DheZT7U4TMp/vwkSgkFYelz1oknrgANDptevpAMEyFcLbfAoObMLvW0qUmfokL
4LXqCsHvsLnVL39Bcoxeber+z5ub28kP1eZT+q2/rtzK8yJlcHCShwM42FPjt9Yi
TxNZsNm9K7Bzb63e5bZA3t9fE3KF7NG61pTTX6YFBgGuakdDyfMD+yeNBsjOGJZY
nEkYzrNgW2WP+OuIlAu44+3IuBtpmVYLhtC7M+fypv9Q+R8Vn9oaIKxWOzh/iQCS
x9dIWb11GUMXdLh6Wei+BihVKBJMLC95bxKUGFYatT1imSUADRPMjUQ1SsbImiHD
41E3d3ovRHqKrCijzOgyOIF6mamtTf3sHg9LVO0t9uFAHlBgiGYFfetxGiC6NShQ
5Ay+FCFkgjpuEiQsalqwFqOASlNhknpodluN1GBghzLBrEMwXdR1jCbGqQTmmoQt
GTV3RlKKyapdtHIDgf666lw9d0B0mRi7NTrwqJ3VZp5Z9+kYeeAQEHfRNvJ1MSjy
XLOPT33HS0emt8+xtPZsJ+7WfLWneUtcAby6qGy2BnvMtKK6scwea7bgTFAG0O4j
AwEvi6TMkitVv+Y8MbmnakjHeXcJD0iOnfjlP6DtDE2gWER/+0zi8QJRZnBpxXz4
XVGKk3mETNLMrnD3uD6SNHoYwOciIgp7kPQxEuuu38la/c0UwagVu8quqG26hhqV
5A/Q8czWkwQL8BgaS2/uNzEPdIU2M0vxBkFOd0/fjStf7Z4/AItHJSuifSDE4Pbd
plnDi50ccGjSQbHw6ZsKPaQj9HfMbQWmkNT3nLzc9B30nuNXlYLfDIY7mtV6PHiK
PVvtdQPc9Fp6OBBofwEMJ8GhoXI9YLbiWWCmINLa1To=
`protect END_PROTECTED
