`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NHvlO3/Dts7dIjdOMZNz6nmpTifeD5PluhZuaX9K+/rjAN6Q2l9O9JImvErLduI2
1xYLg/MG+YRCq+wgAjv7CJCHhefE/VtGmWiTpM3dzCe62JA9MMHS5XXlB7G6Rq3y
AVbYygYu709MqRsKNUEmXAb/sSp0ARsK9pfNCkfEAXz/C/Fk2pp4eXhBCpBcgUML
ucmznVDOezc0TLIg11txBffXBS/wUkrRnTqFt3uPs6RDXl9Z5/s0Qi5qPcqAJaL+
HM/Qm5sBJIPQp7pl2Ya9nYZxd/rhcuPBpYMUcBnyxM1yd/jnStRipdJxgGEtLZH5
jqaIOQ29RvEEO3pqJqIVIB0TtDi0Lkzg4jZtJpvU9lWg4/r742C8+4oLbMT3zdv/
FX6x9gzw/mgsbidvXD5T6whpr1IPVqv4QX9eduwW/6c=
`protect END_PROTECTED
