`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vbc5a0olD0RRbhgggZlogOlIMYJQGGTjkp95uEI48NT3Ti9SKSIKJVJi03GikS42
5uV7JQgv2BbHgqtk5QOxEByDMrNUF3wluorvpQRY3b3TTUtCyaAkrmDVJEIubbxq
V4wgKP6QY+w6eD1x9VeiTlMk8po1Cv0SF8Bwl5/cGLtL/6B+4VYO/oC2wAOfs0mP
qBz7qnwfHx8IyBJUzyGCBsxw6cIjPM0tGs+QZydO9U0XvnDJ0YIKggcuo8u96NHe
qfZ4yyFEQL8szITKt7lLhL35W2+h2sgQEVsejs8Np3tqUWBi69w66wHIm27twzbf
Nuo37UDXalXRyAxY3XC64jZYoz2WiIg5oJl5RPk0DctuqDAxeKgxqMMz0YlSFaas
SlmQp/CmRaZWW2asbnZ4WcroyNEl/JJtBumvcXY5WOGtLbjNv26ov5WvZHbKCEAk
CLfetoNnpmGeGbNmJB7YETv2ryjFyzNV8IMn8qeEab84ikE5dLpj85R/U3xgIQGV
qztcLq7SGevt48qa2i38+0dr1i+Ftn+0Qekd+bKKcQEqtrAiZ/ZxlSgl123J1IKO
j6i+25D8FCIcD7EozcRAZA0oP/ftZVp6AAbnSSM4ihfFGddZfHQ8xpmMH2cDFwgE
JcD2WRuC299YeEvfCE9I5V1E49Bk9ZmwLQykA5t2TQ8ZDHkVTKTOB6Ac1fbxqMVh
HwHRtMc3DFskc25R/tmJmM/dWZjvObXigAHUin2NZt73SStycS5o1oSHU6Lk/mtO
0dCsrenNaGkcVykdbYYl9yBixF7lmm9qQ0kV3qjhHWFhsIFkwbeu1Pv3WOLAgKb2
YZVjQz6vOhvb0lz5sURzBft2jUzLqty6+KjPjvc7ZyWyeHID6e/d4IlNCy0vvMIW
sOuR1xPLJbpMeN/GEaeGTovi2+r82dsbQzf3D+VuthZoGxteO9WAUv4dsKJukPBS
/lubnyKMK4tWdGje78nMZuLgBXvq0/Ja+3dFnKk6t14YQcrGOM1EegQqEOMaPA77
G2JLAdy+x8XEbfGBLY22nR41Q0ERjJLUHrNf9h27dSzQMcs9pCODFB0R+WHzHhBE
5VkQNjnSNUP0mLb0wG6WNNTjXqLJwxdYwOh9bJvz6leNkHxXzlzRFt7H5g2MFm8i
GtiTG5dDqsMpYf81vLOSyjUvTZA41qn6Oz48dt50h2opyUMLcpXqGV0318IYbjzc
nuKHnsgdY0VdNF51CcVJ3WqMnY8DpoCAsFZy3T5oZolUOqkpEYpCMxrYQ6COsC1M
yJioYE7r5sXvzfr4Ja74c5kqryNFVLE/BHhfG4Wg1qsNnAUQ8nO46vdeOcNYGM0o
fRcF+ghFxAGKnGVh2OYMyCJR9l/+4tLLYMzp/WoPdaK98aZTC8VjZZUkMksh9sKw
wpjO/n5kO9M8z8Vf/ZtIFJMYS0Hv3BX4+syRCn/f0creqhQ8IWKaUF7NdpSbtVn+
2fEMgxKNpe7Z9u1WXxNhhqmJK1CFUjcgXRWUXTyoog7U5QqWnOnNtWj4PCJA/z9v
TzRCTozTMl+MCDScVi+4yOS8OnZt/irYs3RCNTV5N2UAHiihFgGFUd1CyVhKOq5z
CY+ydZuDsHLBwj28FJKYVxLMqAW02GYps71LgssQLIZ84CbzJxD61F7pWg7GLuqG
q26h9UzQfZEHg9BTft8rOPTxFK2GUE3sx5Njh9xbm86CgkWAtrj8HJurbtlunnTm
swBqAzVDK8UksJqJQrjLakBaFhzk90cggo56VKDpf24N2gpPClcjI1VO+YfSNL1w
fLFGJQLJkY2hEn2TrqV11sxImB9FH7ASXKm2ywB/XS0N7nYWNku4VhnFjd01hz5i
5FanceC2tWVIXpOP/aHkW84aIdAHx+SzRvHe03LT6l452S7s3J0jdzu8tfRpXZ0B
hb5IJLI6W3qJWaDUFqIJJQYI6cS3LvlurnIIOU4h9gATNDWSYTRY1RAr8PBBp8Jl
loFGKZHv7PIC8BSyL2roLtwTGrhdYtofhwJtqJeWeSRmdhoP6PbLOqFBGmV/hebM
vSqyzKTw78nOGoJvgyrP4OB+nSIDkzbhU+EfixFoaYOu7E68s9FPwzCww171z8ku
HUnWoaNIMctppx9sKCBXWVj6+sD2VCNnsTHXKVoUUC5qWo+5TYYxInQZ1KGrOFIH
9Sybzvx9/KB/WiLIkHfORF+wHKwzwsK1qv4h+45E7dxkgJhgGBnjO0Ihly1VWooB
ZaZdDqoK4MxNv2tmdjT88Gvo6eFJ0Z73oaGvDqcwO2NQwfCvDjePOqMeCMIr4unQ
/FO5JkbIRnGZ9ML6bCjYIPyWC3+vOj7yJUO2pkRnyVrIoG7BUvTsfCKAn2yUNvXE
QCZDlM8OhUJJN21VYqKrDs8W7GVOnsxyHatdxZKxTQkoGbvpSw5upMlkyk0iSNMn
SlE/ycTJOhaw1qmRgD+KVwfjnpuT0gvvuhgus3PcQ5WVSxZdKnvO278hY5xmDT+l
RAXb/jcgxFY1avgHX7BHqCDjGUk4YtJxE/ekiHTH2sPxkdNPfWIstmK8cnDnggAV
riD1K56JfXBu0q1DzzF1RWKu3WTbbzDpYRjcA2gHPjac8JpL5vP4LnBl9AJGvUQO
Xki9ZnJP90QOU2Rd2ZFA9HXFxnYfdZsTBzLJVROvTLqvqWb8rSSKBCZ3t17Qbr3Z
9IsyQ8LNVU4Gudv9BP0CPltJ9vumnvULrTxI/WBG2dbvnwlQq2KqM3EXD6aWGJhw
JRpp/4/g6JuAZ/eQFyvxoP/d1ZhjdtIMszQk4VSlF0tZPxmA7ppg/kHQaeE2/W0G
qZqo2mxTZVUttWsYnu8jiKYvafWo557RMyNKCwpr5WZIMvbIZVD7sCu3G+sKTGZd
80swTtr7Q+NqTjdRgJ45R1ELbDD/XGe9yAbUKXUzGpSJVGA8kX8DegmFi3q4+MiP
3Av9ZOBWU5eycS4kJrjWsT5OE70X6/k1EtKcUU4HQc6UGaO+qvMpvXKfSCNnphdL
Q9YV64S4lOsrMAQenPVrypf39Sdfuq2oa0JithLsOUKLdCcnf2dcqeFZrhnnsdU0
UQsqOmmch8ROEkSZK9x7s+nul8YmyqmalkAaOCH8wCBFGK7dDv6V0av99lZbs31e
opAGOhtTy26cOLD0kzq8srUivHaVszUIrq2bxmOOZpvJl33N21Q6MrBqlzH596xE
6TN03eWhhGWDcg370Rnb5S2rOGiAD9Kr0zu/k6CB0M2FubxdmLiXLIg6ct8/lSE0
qFnKQ4r70XcFeYjYr85Q2mZ9xT9zEcCUtFEyZtS2WybiuifMIsoJ697p5vtLogvA
BLHIBHYHj2Yin/aoANSeuxSMO0LV2tQTGGki2grvo31nKi+hznnO4EZT4HIqP6zA
SIdAGHLiZNQFikJoUFCDEBR1vishZItXggB75Xi29v9fFKJ3Gr+p32Eh0TuYVzB7
a/QoJBq1ssZUgTIjHPuKznEGzQbrZqdJBfmha/ZLCq1evMHAmxo8zztCeRE7xFsO
/WEJS5yO5catIIdOczVB6GVqx0h/r3+MGPZ8NVEbfVk3JbsjXO0V5Y4BmAH6ufGx
gnqqJPhCjzoe0boUW3YLEVqMT4yq3eQvJ8vHDs5a1vklgHT/EXtADnrqff+OeuGU
O3P9V1U4Q5GmnMUPPJfIFPMrCaqZXoFM4V1GQGcUuVIgEf/7h4WEmI4Us/TsulWT
EtGQXHr/KOTovbdFSp8mWMbat3KZrqrrzfTCwCyDyikOHxJLwAtnE/eRfLRySBSw
QT5MiODn4vh/Dso3uptnggrS4Ibd7QR2y0lB12TV71Nohp2Rth7HyWt+IEws77rS
n5omiBoNaa62kKsBvN5ZHsl9U7+uHYmY4X4252qdA2WwhT0PuC714AnPOIHxPAxJ
HtdeOiqyptq4i7ImToyA51Ks0RKwcK8I3ojq9R5vWiO90FWq4naRr2sf3t2Ca2AH
/XSFcMBy8Pck+uw5bgeoRl3BehcEvf+mgMdvQuCvNZZSsI1cYPJa/uIFqEnvZK9R
BsEhIpBZkxApEBsLLxq8CSl636higfwlg8d3roTGEAuR49yyEHoY1XOsHlkahros
tDDnwP+uFBT3mUfcxDzp0cIaUJBlooDFhgZlPx7z5godZtxrP39CCVlGF8i6uuAg
YUFzAQdSIlZEXezeBc1MdwWMvJhACNTYAOOsdKchP8ewa+6c0AaAzpwKrmbZUj5a
VrDiCr330wW+jetECZ7jwFF9n1eXCXsdOE1O1rt7Dq4ZlX/PZO1ct9DVNcXpIUHT
5+aD+pc7fHMXkhusLk7MUeJLzt6YZXAoJG5eW0rxECemjCFmtKe6SUWsxvkwteNk
ZTHsNlx2m2y+yF7u6ySfFZqs1xBu06nl+s5qzrVatVyu4KbDblyrD6ZPU3G96b86
dKxWaSXoKPEp8GG4/ukh9UyN+Mf4HbUakx0XxPA690BE9MuViO85zPnMEbhOKGvX
7xVaAjBJmmKSJyYLKW6yQu+ZQDnl79PVYy7ZzTU+ftIDgtNmm2Xmbz4mzUlpfYxA
FzznrvjtP5dfsLleZawdKK3a3wImQLvPr1bhHxtiSAZ5s4ptvYqF/BT2PQGX7eRW
H7CGg0q1gTYZ4Ob5vOV7bP6s35+EVI0aFAAP5m5rl+C935ruazLwdlyVMKw0irTZ
83HijtzokhP63YlQPV+xPdQ6WE95dH4/jZ0hnQO0hjFKix330hCyebdMDrn+khF4
538LFraMBJyMvx84foIRUkk9re/JIJch2Rdphsf0gUcYqcNzICbx1bfZ4HhfffST
Mrv/FLTFod3GmJu4Rkg5yKisGo0DqrfRIwk9gSpTNBHIliG+ZnBRrCpMWSpeH6zk
PMlN9w80F37sIvVdLVdlJZ/750gfc7mcieuWTVaN9DimmwkGUIV+4yQxD8/9ruga
Pdp58WBSdjfSqeqJqe3dkfQKE4vDJNf3S7VAT3e+r9+Ow2Ng8vjZEs8OUETccbD8
sOeE9pZoVH6qCPca3rbIVF94jxulWZd/o78nFyUzhIC38ydFHXUDUWdPpSOZHf0r
rUSoxP1SeJxYzc0CW/ZZ7NrGMVoCnAIufsUW1llG9+XMF3SXQtINJO+qtWabPImj
RppEf7Q7/XDJoIvCKoqoo9sXkuJ6YZ2ui8ErtvYEhsywGQPB6Gzv1n7EoeH6fEn1
WLNBp6Tl543TxuBtLLU90/OFippR5QBBININ0uffpZr/2M3YsYumc2lS/CAPAfQD
pRd4JG2PZ0mC4v1MOPbNV8CXt880mVgGLaRrq7VIRp61ghc/Y5P5udMS4NNLAjiR
CsF1xH0nmnb+lK4uMxfMnAafnMvpEn2yu5GGJ1+2QCWqoQOok2gSFMJYmU59HbgE
22aJ4OqgQy4SEN+uwlyxCJB0krYq06ZeJRoLTUKKkVU3Jsy01xp2fljzznT7d7cJ
Xg/5NE+rBxMqS2xnIc4z7aGGI0cAHIkEdLacIjSKxoWMOGHvsB68oZ5aRCjWozGU
qhvPN+3FQN/TiXWG5ITiPQ2pFBfSwF2PUahaXxsAcrP64M4qlCYrqUI/DsqK18qN
0Zqemh5YcVSbRmEkEmyheh1b42FZGudyc6swPYHmuA9sSvqJbyROhHOXRyXvRGNA
H1+27MIUdXGJy0KeAG1qLfCMkszGd4oHSPLyNE1PfFCseZWGHpr+YQEyoEi73eP/
21vrMnzoZ+LrI3x31Bvq7wm1ryJqOU5CknKzByDiGWHvDVIdmtrdAZ+6wvARf575
3dAdBgOAkuirRLrKBH/6lHjBThxnmz4HpzxCf1rEA5LXzz0QvpNmEo7pkVF+Mujs
tT5NBXFJ22ZTa9626zqlQGPSq9RFQLEyfjXKP7OYI/42mz4+lL5VcUv0YOYkhVKa
fk+FcEykEsI9RIPPUEx8SW5nvpO1osxs9Uv3XoHAjfB2FeTQ5mBwDDMEXPeWk0QK
HejdPfAjxaYzkVRRLS4EkspK2m5cmsn/fn1asw0k4RfCal6H71WsVRnP3zRP7e3/
C2goaZj8YR9qqXKJKJAFQF7V6Ap14gvPE4ujb12NEO+HcCd4vXpIRr15Ck95UL5P
9HfoSIwTLe+7pDpnWv6JwGSHbZU1rz1Ff0AxtIQSuvBFx1VCe+llQXO9zjx8pQfc
y0L17wx67Gm4bKES8kW4utH7bEVDYughNcjdrg5sHh3cvW+ORADNvRLhU/1OVCvA
3ht4gIoDXkR5ZISXGsh3gTRj3GprnYY46BnID0mVHrsrUU10m3qbsvEL8z7tjoGW
WxavPNGKtb43TalJwFfeEr1lmj/I1/ezNRHs5vH/qpsDV9eEVX+RplMWeRLwm9e9
rHCDxVvWH1C1VT/U7EOonD6nzh/mmdKBKB+O1nPnS1qb46mGt/YvTB9ED1bm1mjI
lkchhef06bd08BZ0TBl3XiCm7Mdb/9YFNqWIK6ssjL7mPlUFvjr533zhYnCyH4UN
s2C7FDiwkWPxeRvKeZviqNSmrzV/MuQOUaNX/pLejNacDhM9KZxjGf5vP91O8jXt
jRsrOcFUBviJOgUeorAG7OeO6VYGugEHFGwZfPiTXgi3d+8+khw6yddn7JdFuD9e
JIfLGbBpMBukaXZoah5JnbHzKPdpxkok6HYyj8+3tDOypqaJ86a3qLwlsGNiP6xI
T0Ni1FFxpodvfJv2RmzBtflJKA8xN4eauPhVvm92gt7Pi9on694U/GcMMo68Ogp2
erE/qGKBV7wBbb4VdMGR2FBz/v8xZRINdMV7irMLYDAhjd3A7Mq3yHpfjTr+uUJW
8I9uVNgLmSf7f+HoRSmSjnGwvXh//lO3pXdCz8Y628/UXL1L4DopJUXaeh5fPOF6
cQcI3fnaHPpUznmmK7rT6IGQ5SKm9qdczK5qnRErQVhbpUfRE5Le/qGiMzRUJvt+
catp1mtoFXJwewDvUVI+j+M1DKru4+H4SWgljtUTdNDx3nhCSOYy0UfQTxBjq+oz
U4tl/1OImEgO8NoyoI/OIg2O8BkAwOJz5WivgZW23BUwgDQvhXFmRjOkxW/RHQSw
9x7qWa7zz7teJHHWQ8ezVMASLUBrWGM2B/t/EVeOMB7oEdLfg7EM3iITyLOZKzQN
fjjFJiaIWWSxYEhdU3d0evzHCyDlalz655xcSbCwlhIkAibn3xZUq2/kRzsUfJUC
1RDtQKgFbpM0BFuTTipQyPL32T26pO7akOWlNQQ2bZ89476rqqOgd4sG7yCJRaKO
VZldjZLLfZI6yYH39Ad+cApLrI7f0LA5yjlOc+1B9MAQL0PMwNyvAKIaIpY0Cyyz
zqeJJZY3Xxszqa6ZKJMDKqWuh1SUZ79CM1PbJUDbG30c3u4WB+tL1mfGRryt590+
9Q8cOsJ9GCl0Eiwbjsx9UjRyYQS83OQFAPE7vlsqQ4YVzMxWhsItVX8E//3egNwi
am+k0f7Q+pRo8mAjpdt1u0lkXBstjxq3rAy8WA6r42okWj35z7uOurxFYfsZx7aa
C8pjUqQz7lJaR7SMtgIgQUqZ9xV46GgVSIhMBWOdXRyTB9aVdBG0u0oM+RCbZqBc
qERrqgxmh/y0tGUjhUjc3wXXIDL7Fv3LhKQIMKbrVT5OHu7BwvJYDS8lHtF0sI7z
DlcMFQkOyd4biTlMhX9qsy7JklWA39s1irs5n6DrEsv3nJWFE5I+pzpZen28m/Gf
newgJ25+xTNAa4CEC2olV18jT0GBzU+kUeKc1IqjMYgPAnmUvf6OqfRWP+P9LSxp
DG6dKR2dueynwopz0C/veSGgpnjfNp2WRB4fAKdqbfs2X0l9i+hiTOxdKXMqaJsv
SQuWAvS1pX8IN6Hsq3Bhqr4C1aF2FNH3Es6GJrWhD4++xSDahtr1BWl/uPB9I3u5
zJxXdYqVN4qHNdZo6m0Je22BRAupP89yLPv8qrEAFBjQRaK36EatsUrvGFD+PJQy
ezVloGb2Q3dadB3cZehfzv9rBgV2jx1Gyn53gC3JKqJTEObbDDym5tt7rAGZGKA+
Ll/sZRrA8CX0km0TInFw7P7Z4lnLLmLTvqKmay4FYCjYIpKMmV2tA/im+OyEiUPu
AcoWYEDtheSl5Z5Lwc0ZcHhAKAuV4qYtSJvit079dvKA9Fv6nkT4vq5scUMWC0GT
jNXWSSlJZyMzb1hO+aG9AufGg2Bbmf6hbVeZJOz2Bphfi4zxQ2C4U1aTRWCIGqCV
HHRE2A1/E/Tn04RruZEVEbZLoRMYdjwaLC+FUtKRx8R3+yqXtchkMwAn3ikxKREo
ODuzRPD4CfWji13XzLaSe3VXKPQWmWGj0OlDKxiQKDLKhxhWlMPuHsCYpn/21n+u
G9F4fHkMaXIQmHxwz3lIGRahVxh90C1WZM4HUU5jNLgLfzQMbV6I7fKUOfykBShb
U/EJPIUCQJLmavUjlNa+okmAXiepbDPdUFPOp4Xj6FgPJSExUGtcuRh8CO0grS4n
kkKFDslsUwWL4ru4RN6qhh+JKH8u4sVVu8zbevAiSiUYZ9U1VL70G98e5mB4RHd/
nb39RJd33foWIyF7DY9r/2P9qrniAtglacBACECGFL/G8mbq5t3uc7nvefFMHfJQ
cMcKDgMEoT9GtpBrdbXSLYT5/FU6QFbyXoHMRo8oHyWy+u59ieBQwUQt2gvv9AFA
23JyAeIw0i+WwHcfx4/+yKTJdB8Ii6j0VcA5Qg4tg2OMm0oeN1DhAPJSvShFXoH3
J24MWL0EqyCOqd64y0b8uhAYTPWwj7Mve9Fsi/EueTg8zW8pP4gbLaBTXl4Plfdq
4MVnNJqNwVyNTSaMy3L/88o78sstaPlDHGCFhTl1BOuDTii2zAAwUt9wD4r1hZP/
xHMUSZ+bx+z9r6H0R/dOcMJ+GNXrG+TBEoRoNrtMT0p/C3QlPzfOvlIGHuEyUg/i
tuPRWtJHsQRaOZhQ48ZOVJnldfihBw4ahHt6hFSh+T6k4JQd5PccoxTuRq0QoTfr
CTw5K8ZL5jw9fI+eSSDbu1k3qUMLUJjT6G1yCZC1MH2dZ9WCrEoRUvNEPZgKW7K+
QB1hHvf2OyAPf2d4L3XKPcZJR+PMbXRsqvaRf2pCSwk/9pcS8icg6SnlZcyGpKj4
ldFogDrmgV3MGE7jlik8ROB05TgCegPcKQgwBO47EznxsBV0GF4WmvWZcYj2kXG7
C4wp6vYbNWL4Ux/dUUfRQ0WCHLrUO6WvJAQBx4LzEA7VbtdqcYCB8c9wEzoM/kGg
rZgJgpG+vrtoErFRqt6Hmf3kiUqlE4XHptcZPgeBexBnMiiui/J8bj9LeRuNRUsH
AM0c4MR4AMtM7hSOiv3blV2rmUcO2lCv//pbo2DuZhQlzsIRNFWKN/9ET1V0Kqe0
9gJzfAyo51yAIk8Fm90BtPgWA9WyAYGT3va5wgZtg/oqViTHoGI1cQ2Uk5At51F5
6lPqf4Pd/PQi04j/vn6xP9HwLFoh0x5AbvJ4r9wLomNJwSc9An+M+Zy0A3YJlMeJ
4YouyVtkk37cA3ldk2aS1mtLow1AP4Vu1Dgym9Ydf9+YICj2INZ/6eLQA9Ryk772
dxtC4s5BbAUulvWPY1ZlMD9yDpeNprPmLqf5scaBMGuZ9smthjPZnB+dR07r3oCU
AAG4G0QdBwMXbLowr37llOzoRQWW1igE9QQXUgGOLgbOEtkVaJFei/nJ5hx+UxgG
H/7QRiH0EvBjkoiLRYVPIi0TeHIX8AAggCuJ+5v+lqhk0RjGNbc6So7dRUvJ5nps
r3oEDBN++TtG2lxdIlwrumlpi91Bazs9UV7Dw45tqchevCCqVVRwrrcTi3bJpH3M
47NZzd0UQ8k5ie4XByG1wXoZ5FKUzr0Q57i89jOQvdyzy05U8lZuUOTbTXhDZAL4
qotEukkTxjcEI3zfj4LxWjXZG6yw02NJY5ACLpVZqgcqp/KZGaSQmZg8I4o/NvXk
qkRQj6x4eBOs6z7CDJaAmorb4RZZcltMkgPuoEHk/hcsgME+iRh+nXJas2xu4BZg
YjFa9iSEy69Tt1SFzIo8H5krBJ1fjnLBut2wj0WHSIQafI84wSmOvWKFOzictbYT
yXXmeC0FtBIke17xcRKKdbk5KhEBq6+R/f4O2ZfBi9gfaX+lNfg93UYS37X1cHhj
piRJ0g0fO8bL5hBjZkSz4uaZ0PlTROxBlPwGXtoxCuhGwXWy5wGYsscwR0HGnJER
gDfqguIW6CuUSEPV6quRUtjZWaFdDzMRFHsFG7PBoNJeMNgt3d1G0cKZRQ/Ue8o0
BoA3d1osvwRtoDNlTieW4nyXTiLpWOD5oapt34LlSbFMXo3W4+1VA7uvrZOnDMJZ
ii5cFc4GOhqJdqUmv8XQrXgztCY0Ta5vERyohMFXUtqKa5wqZgw7BwRXTZuQgOa2
A/mcm0mdqsmP9pHbDqKYvyNA/4OHdmTWNBwCRmaZjCKd1RmSUQxEaIAI689z/f/C
RAW8bxRNf70MRf7KHErFa+BtJpKd29MA6xGGszO7nE5Zn7P/i1B0saU/G3TQYr1q
2WWy2OQ4EvQJpGF8mBatwd0ksPjucmN6FrFrwDHjWRas6Y/7FVSLpS8In0kzHpsl
yIe25CuezTHOt6l8ZvvHXfhX/7jQ/TqL1u6WDBifg8XKd0VWHMJuGOIrZ69bR0Ru
reprf0lsOOlYbZlA0xAa69jHSfi7FMXl8kMJVpJjiez3Zjz5dVHg04FQ2skuMC4O
oK3Z26MgcdzfM0nrY4Sx9juJm/QFcai1bVzXbAFwIrmMbB2NT7zbMmyTNS0fqZH/
197KLrNzT8fMUulQqiuMuV4HNTMKq8d74AHVvX1BetR84rGJnLt4Y5sHMN8/mKU6
yIcLA/wRYvvpiw4SJk+38GcPLPHZLmPwV8dadBhHmNUiuPy1TpMmakBidSOthe7E
HNks5e1g3lFjEFwAzyvYNN371h4HI1SMiMoIyvYOsnXxRY5I01IU6m/PYctPd1Tk
jtPbA6DaNofksg/E3CqGJgMbYY5acwa4YOqFRcVgvCEBKqAsOmqClUWeESMUdsP6
VG5LC8BMnEJTCMPVOyKEiRJmwkn6bijgm733D4Ls3dVt+FLGUriz6ivmbPs+2sfO
0GejNlTu6/snZXxpfoYmtIa5oFU2MoUKP6Sx2phHo1g4R6tOJqnUsj7bFTMJ6WUz
E0NZWPJ0uvirtwRmoAniTM7Ym5feXlEAoAn/HXdTL+I5RdqK7CxjbtbVwufm/lEP
ACFq8bKHXWDLpYWweVvnSU5OYn2HpR3D8dudftrpj02n0MVaqESKiRQGIn9vX9/d
MZ/NLdp7/3D9c/biej2RNreFLo/07mWX/K8MnvCo3McluQ6qB3hwDZFjMV3daHi3
/BMFoj2S/rg2OAfD3le62A/LkeQF7ETOXNu+HHnfLLB7h3MaRbhpYGvECPM8nF+0
2V/0MgeOlYf+ncPFwvltL69yndforKzu57ZuX4/nkWaSQp+9diSLKCJ4qa9cQklD
oBLk3vx/O1nMEIMkWoglayrcFBxYUcAWz35VKx/9eXAHY7I3TcPWeUAy9LUjB/Zc
zNlrYp8EiRuPmvRKZkCVYk/MRt2IyD91qsYaOdbQEMa2ll0O3XUk+BPNHpiA8y7o
GKz6p/3dcq+v5lU0rc2VTV7uhblpo05ipCz+g4Hojxfch94Hd3rbZqh1i0QDn+be
4hlyN5p/LrXexFmq0AX4fyAEI0SecsjxkW1YaW9+TT/TdCfHlnOVSx58+PeZPXsE
hcQefGdPQls0qPS5rO97nIspIW5B1sTnXbboA6adT3qiM1ByqgsLKniiHtO20nWm
IN1B5ZufwgG2oNx7K8svSiXd5d4T4/eHxVdSvDKbTKVJ78IsvYP3IqTZ642/jXwx
6NbyMLzXAbBuPRy6/rbFlJaDrp0hgZKyGY8FPMQJXGqAmfxBXWcS8janp9eNpj1v
T2oiXbgOgzR8jr4syBXyk7kj7aF7jVAd+oHLfYvehFh4jDSYr1Bo/bOg2pk1/mHA
TYYP12/63PlxhBskQq+uQyURKZGQz5syjG0A6q0oG9oPlf8w7f3s8yjlVki3V/2Z
yA/kJHiPi0jLQxRFNesBssStjQ602/fge+g9HDnTa87MD1GUBrIGXpnzE7x5iewS
id1Ifarr3lADuzEanVCRwPVOoqlGyfZnMuocridzRbOeOpd40DDiMkc7/47Exxgj
c+sYrCtcCScIKXAHohh7GaCPUV7oYyEJj7iBvY3JFZCGZtWnHPu2/lMioWffH2Qd
T+klK19ih6zoRdg5tHRvOMrpooQt8mPryR2iHkOOjLCxfM4n/DwcIjAho9I1oSdq
UKMnEjXYrwiaMsAx8E8H86IYMgqP82mYIfpItuYWlr+ZdPl3V9O9STwtwHqJzGFs
zhlFlqT8gDJu8z2w5gTxJcF8CsT4HRxtv9gs8sN9kCYHZ1xO3PEnFtiCaFk7x7jd
T9aws7opMNzYIl17tW6vc//9Aeq7G6kHLda17qXtAQ8IOjJgoEi8PCjrwVFhMewS
kbwtqkACNesXhZ/vs09zk622BIVFK3R2f4PbDhxxWKrY6kFaA3iKApGmxQc6Y15Y
sohyt/YT31vH3x8xkgM79Nnple2QWHBp90lVwHGU7YqL2HC06IfNeSvp+16RzG3C
U8GcPluW45IZ0DJAOvvmUnklTirUl8WutmbZOCsT9hbtXzXg9djg+3QxSNFoirSS
BBjeGSQAFnS2ucN+Sv/sgnJSUBQvDxOkHVllRH9uVhTcfY5RtEdGvePOamZUb20n
lxND/XrBW5dFPN6k0uKC45To26lawIWquhGAeUoxvPzFugNfMLIZ3DdJuKwPaYE4
2hBfMHvbCLs4D2/uIKg7gzTQc3wMEhaoXijo71xjP4ljtTTUTd6WfFina6kOabRZ
jpDRKsFywPgsHm6xGi0yU+NPLrPHKIxiKO43n2hU5rLf6FHE3jZeuUZZit8SXVzW
G6N5NuKyujiibb/j5T9oRKD1C08aVg3VWVcZ8fUeyK9CV3fQzfLAobXxKJT5/QqQ
b6w01I1vjVY2NEGM02q0pXxtBwCBeE2kGled6lxSnRavm5Nog/VCEJCyAGH3Fsjn
c/+ca4vRXtA0GYhuow2HyYuYl4xF7bsVCotyYnH35TqOV+zArHdo3BpZ7dC4QLpk
KMm5nD6VVdK33q8lKxKFL2yJdIR+J1CFUQfcKO+iixdzbqYnZImcZWu+EG73I9bU
2NEaTySQnu9Wljgy8A3lxOobP16Pp2QKmAlMFxrODTHRo5jE1ST4KcUvoomDWdgx
V2Rlb1r9zjx+DahY1nYGm6oIzQEouRUSNueVXfgZP86h5rqenL+DBAw5N1h4rbEe
11T0TWAoNQolo6cUfLYMbZ8a+s+d98Jr1bzPdlOU79v02cVCQ7JM6LpXycVhv6Nh
CUfgA1gjXpuo0iv3lS0pHOpZe32RSFQyKSQodnOdCFu3rdOnmSaqkf0ZdqZHjlJN
OtDm0RaCLOf6YJbPSkO8EIs400aSO3/tbEKvRWWv3V+Y2QGuGPtCJz5ENJLgq/gh
gdgAMq/zXrSOMx+lz5iRghdxDXss2bppgqJ3LIt5NQWvTQkLkdk+LqWHRWZIo0/4
KzzVsBqW13Htr09gGaItRBgz48OGk52ZZ7Mnu4Pm9VmvN49lQuZiDqVvMhAv1kbo
0vqsAz2UTcjazlNfk20vCqQc7lfytegVaqj50lBxjMYxTl6AiZr4alsyRQ4zlo8p
58H/6pn73B4SvXnzZJlVJdSu5uJBRDB92BtW7REuc/oDyS8zjAbZB6qgoDOFTs+u
jbwJMpylFMn/DtVp20o/Pz3aJF6lT3Ve2//J5UA0J81ZYz7Gm4AGIFHcq/oXGviS
DuydHkSt2C7fjI9kYJbN9NKIaXQKZkMl98S7nJr+ggpjcxqBM3A4avSHzl5/EYYU
Y4y6FeyeXfxF/tAb2hvCPHZywudRmwRiYRjsHKNKPA+9yJCWfGc8i8ctR9VQTCIV
U4NxtSJWyoK159kaKLOVVyaI7C2QVKdLE2Y1Xi8eFmpqlyBgZHqeQO3+A7HJAUdw
QMxlLy5ua+rYv8qdIrj6yANNfarLgwZrdJ6nma63G72RRkORO1nPflj/Qa1VOzQk
67z0qLTvdJpR9LeUfOM6FB71SArkuBo+V5JJyLzCmfxwSpr+O1HjgybVqMuTEQPN
hput76mjpYJRSryYQOBReOz7UrW57ibfM9OvEL1g7uPJiHzhXSx/9b2dKbenqlSf
AanVa2n233IKGcnjoBNkGfzKTBnQnG23RMHnNQqVgRLb+0IvPGS9V9eSeDQjFE//
uIjSrWkd/5DDrncU+aSZeZZ81p228jal72lmkaSEuCPaNmnIvxRZk1EOY3dlpj6s
iUF/h/XNV7a98lGHQJy2k36SgZlK2taQ4wsNI7WBQVs/BII6PnhsQPwe3ixhLcox
NPBpYkx7vSaWC2qaS5NTwuZfP8Z110eP0hf+t/NCgl70ZrD8EfRnjRGeiV1LFHwg
mqeq6Myoxm4hu4uzyShlvD6moOcZc6o9vB1mmRVg5qgJFemL+pUHDFJ92UCv3U6x
mWA1SQvlhwQGcPLR08u3m9K0zXWqyNNQHNxSvULSsEZ2Xfu7HxIRBbRBGrhtPGWa
+LIpZY6GEqS/89bXfZP3SK07XITX4ckMwbcQEzeaflbDvAdRZRAcdS/X3C3clsUI
lFov9JuaZBZzkYjRXjtWKZOz/0weF2alMe1Iy6DkmiinXUc6uOkAASdScBKlTpSC
Cv8v1Nb/pf4HIJsgrMwkRoJCbpdV5M2hMBPbNbtgUGykUM22iXXVmNQJfEDU6vE1
BikIqpvaMRx0weiRHHUR1KC9lVHhwkRdOGXKw8mKhBWS9l/3DXf07VqH14y7YEmt
wzEVd6pLdBtYkFUIWmKtfhw/QLN+cuuT1hzTEl2CuTvsjxHVGZ1mibVIYdVdK3SG
vxfsWTQt9opTBQCcExnWxrClsOlkmMWUDGzdFUsVKXedTk+E+Jkgbj89kqUlko+A
yCNOHVX3ktRqzUEGVMDHBFSeOL2phGOYvgZk5htuBO0800ZMPNWzqBIoBHizddoe
42h6HiFC8X4pkZtD0sNAqC9luTcwbCE6JEuAU6hcLoIHQSb4tzmIfraXgvVFavn3
iPX7FaGgyCOCMRmciKFDANrxumaxOEoHJPN/GM6xUBW2Dg6I9peqI5mvXyPV/tLj
TpawDfKEjtK+4hBc2rskBpmRwL29wSbVhuRqywweSWTlookvN8QokIA1vnUNW1dN
bcs1c6Y8RQSZbiB8vjczeKYfFzOX9eRR0PEkRMuKNe9O8w9wds56pYNtagLoklxN
CsXCsIF1jvLVXNB3ncp/T8OldcDnjYTQIB71lkbQdhC4K1GOVKRY4pwyeqtHwIpA
V/nou8yhTU9jX2/jo4QMCgrUXtfJsP0waLg86aQF2hgCV+Rlm8pmJ7MvXDJq0zAd
wGdWpIiWkyivfKxeCO+82LKtj2O9yl2yhYKZuCfMyKZnOxUIDiQGN0nQLcr5os7k
D+CHD1VuGdohjJwhznPHB6Afh4vTA53UMuY2kIf4Hxh01dvFiPHy/XBiMEovgG2g
eoIXgRCj/aFCczLKDo/BeScie34tAtT9RT4YH9sLYfhUdg0wP2Ryd639PxWQ6pjb
n3LEarT0/ihT+laQakI3oBCuuvYsnMkZble35DKaUSCinSdl+H7XeN1fVG9Y85xz
R1CsXOUoNVn0ZCC2+G3SWkNbvzDWcnAcTAucNnnNQLDOpyZCytrnIz2D8Vs8ieam
wo4PdD3I9zQukvtjF3oxYHBrkrnfmbLR0SoRe+wVTfMzMOt4gFDnZlDOLA59O81h
ouHQoggCrPeXG6kff6YfWbeKRNKKz6+y9gFp8JxT5xQgVRDObQeVG0cx2fnxExsM
774Tlniv8biZBNg4PjBFFy3yYr69tFtm4nK8vR3rOVM/F9fFh/ZOq/B+jllfqs/9
qxjlCECYL0klyi8lWT6B3NWnklkDYWvqkDRXSBnoL0mNqncDw+W712p+1HatuguX
vTSedRLFkItCnes2MKAtYBKCj/3hWJD3MjeC9RxCOVlqkq9kIGVqsgP6mBK8qXJ6
WP3logTFQhntGX+fz0H7l8mRbudPyjPWiCspDV8/4Lb/RLDDCPv6Ix+2aQtnHbHW
aJiwJAmLPOE3UVo6qieIfelyB370rGhP4urZ8E24hedtAKX4C9WnNwyx2kgTTClX
D9EBoiE2Gerfu8IJilJ1LtQs1Pnvt5pLAAKAvTb4srtqbqjqSL6TgCqnJuBE/qlD
7UYdz4Pgm7/RMCAeSIljDcm9/HnxFL/+X1KHq41UtDuSUUbhcPL0MsTmpooSDzSP
OLb2HXNEPcv2UYzMPra+md69fBqHCKm59WD4IBGE+bv0Y7K1xP4IKAu2NOapBIoi
+QegLlzPiZ9yRdPTKIn2qFad2tVRtyfCOm1KLcuHJ/l0X31Ewsxi4+oVUgLhnVcH
CdB+mP9bPRNF97g577AdXgb6svj3Zl2V1s+b9Vq0zJxBc0BI2RKArcd+Qc+kVwG5
LWD6QfgJ9ERh6GLWOIdwwvtIlHiZN0pnH8q0xhmx902UvqHJDJmW8OH4ccQkaB0I
SMKfL6WOo1s1/qcQLkfBIImgy6ipYE4K9BYqFe7GVSCHOUxBqAsZORHW/3oG6INU
LC7ZaLq4PwK11oSK4AqtykgkER5k+hViC6ErQz+B9ODRxGJvQ5vo5YWtgooBNxEw
zxHD5UUCs9leiIvXHKIFePzYKUV7FHRYxJukHrwdTnrQux3IVFeYesj3DZHpf2qd
fum//Y1zT4eieR7EvhgcdrjvmA0zRV+sbc12CViQiAIiBqh/y+/SJ0Ad3KVHmyk+
Bx5AHJBaMRZ/t5aBv0rEPUkW/9wm8/UFc/3VjTJC1F9opguL2LzKcDdwETGNSVb6
BIK8CJBi/9jkSqXcBXPzcjYjy9U3Wnqk2yiZ2KhhqY5d4BjFydBWuTbKnTzQ8S3G
qHqwtHSx0nDTRDE9M5BCt5uRFRoEYgYktHlVVRSEobmJ22CJxjDKByfq8lmpS3ub
8KfLGgg2ppBQGj2x7au3T+1ow4t/Wk4VVauHS5GZV733ANXTB2xLDIbWcFMM0Anr
wD0BmG5QQOyzSh2/ukA0r3nUjEEzWQWFdnjFk6QqpO3Aelm6B6Jnd6qnMPzk/MWt
Uy29A8n4xIG6f5JIx2Vsfe5UOPAmo65mWXYXuKokdHPDiqsbDWhBN9gTnb/j4Pg9
UMiq/wJ3BTQecIe3Ixt+wcOnFJY6Vv4K+VwNFRjvQT0OSCNopSy/BoEwRMqm3B88
Ey9GbvYL7Ct+dP4X24RGudiJ0YxAlLt4xmyxliSMJXiL+Rm0EZ88cRbCH6mrDmVf
JhEfKB/7QX/CyEnLqJcuDadCa94b7c4/E3G6taWAoNXWXmtMI3efCu9f7EDdvmTO
hVQBF/8Mjize2GYLiemPMaLic92jEuIXQeAkypvHW90eDZsfA4pOaKFDLp3tlZon
yasKpfoi0whwiw7sibI7CpZ7D8v/usmx2UBI0Ix1/wHR6jvTm47AVBr8ZDkMVbYL
ES3NK85D+Xp293u5ErYN8NcwkRmsxHZoiShvXqES0IFuUfMouCsSkUFWeKGtrwBy
3E2FUpZHzVIlrxXaZgSBwxmoUscsyF1gN7vWnZDTvR1Dq7q0MDLYGP2WkJROtJva
H3NohOsu2W3fiIgf8fQcEt0B2pdyn+FpOiMuamEwvBVRydGovWQjjx/JbEwS+lFU
cJf+xmePF82hQYzZE/1ltgTnOQMeFEex6fRX+9kodYKEm5mBnVzfgEHpVQDQwmni
mqGcsLjbL+Ui/ZJDK+TbEg8CDNSBQDro6N84U+RIt05+JFSAwzZSI5X9HoYBm8NJ
SMxEWdttG07wHC9m++jIF3Tkjo35d6FefxGv34Q3leDaur4yhSqmqBB3jyqzk7z2
mmmN5JH/0aK94ZM5WWw9UBbdL31negV5Pdws/NcbfBRF+Cx+KFcLXRiLVy9C/OiU
Czi5fbSgkAow/VO+eFHeUGFHxzbJby1xvFb5vDFw/D+vBEZkO9vlbSsobqNP+HJP
syGYyCd32VlA0MwX5E4YAy7b1eeg7ejs9OXDUOYUeUCs8x/KS19SyvPuBmPEutC4
DhWuKQSiwopnJhGDWttUzfABPL5tyiVvMBfDEjrNpDLfDJxmZ3HTlZI/X4Lze1dL
RL7JYbIOqeXdyfr+G/1nKoXVkmgg85nVfEFOdyROvZdDISsMJqTS6RPsYP0n1nbT
y7kBZZ55gWAII/E/Oj2QxjFAuOMc7Rxdt7ykuLaHNr7QIUUYzhxP3woEwN7UStUp
45hf6tG0DjEC+kh9LhWsqXBH3Ze2ZF160P3BU9esMe0KXdWgcqpG5mCTou7kW3al
73AuzSS8qVDeyKaO26AcsO7LZNvGegHUR6QlTD1zjlRTb9izR//cOfLg7UVG9D1T
OxsM4+N3Ugf4EiN/ZvN1P52sr51UPyOsGGgsnr1+8ANhy2iW/LhF61VxY4DX0sIS
AokPeeeF/hllZpwPZOQBi3DVFqm1sauT6pCd28gVADtAaghxsqXUs0XkqIlJKyn4
ngfjfmidOwl+nkydn6mnCLu2hT0pMBzL1UTv8rAk9hg6LT4wcKLKzWuK2F4JfQv3
in8t4dmGbK4ESYv0CHxsHtp//xdyCdf2Ccz85N5DQ7mWh/k7MlmeAG97WXsbEVmt
uAAdCgEhRfZV2/d0Q5RkZIampb9xlPjuTk2kxcrKNqj3appE/cOwDhevqN0D+Xjq
Wn+8zcg6dnZ+nWxXxIXYwqjABdkeF660IlYLEd61jC6gWUZXsrSvPxzXPoQO6m/Y
u1UIeOKHNcv6ikkOYK/lFTUl0scF7TtqvSYxaI3ZxJzAhVlxeUmImoJfmyP/sP4K
MILCYZ6q6pNWUAOqWv1Cn3kgW7X8E7fZc9asdMXFQ8N29fdJtEl0Rv4ISkt7GOIg
Ld8b3lw/KdyhvsN2NRCldC61XzEyxeJRTqhvrX1/RzP4AisjNvxakUgJMSln3zQm
mmnl7EkCsYWQpSylMB2YNTanJwehL882wKiG2d0QMusFkcS78xVK9zKyvR8lisqH
WzbXkZi08Dc10kwA+C9M/fqoPoLoPxTFXT+3kygLjUf77DzqZ+OabwmaGhgRn9Hg
LRur26xqaCrkPWyhVAQN85faw76pEtvl3ftFS0NxoISp1oLusbHYfUIln7XfIp7j
wzTsmupXD2yTxXrY1ZePKuU8rQ3dLfu6onm8njO4GvsgZsYVe4549+09Ve3fdzmO
EzISnVl4jR4j4XsYJSr5zdY5h07Jd7qiFHEQcYhtxFF3nVn5Q020vaVvl5c6y2oq
dlkjaiz4oanfiWN+2tii0pjSUL5sTzLxZx6oJbw73pmXvHTKWAqDmwctayh0S2qc
KC+hJ2WsGQl/ttdbhbGbIo95bxZBkRVlM9D+cm6KBT+WwlEXPcXkpVyBBuzBTwry
fmpVv8PIUr1S1u4SmGOXWfAowk7Y0J5JAss5GWe9A/PDycVBzHNpOelDgcL3PiZP
W02OnyVzwvdVcYpqYCTDDrjXqeAN8GCu62Lvaetx2jhgwd+yJNn8/Q0k7YUAqGuB
HrBobIGGlsYCzpzl7+vZY+HXsNyrNJgZz+RJToRpelcAuNMTEa5PW5oqBwp6sY4h
clLLjoBhE3EZUoBi1cTC3qwGMn0FMteUWRT94CGob9Q73tj83gN82xaFup3TECh6
RQGCFjxLxlkGl0jr/Rjk4bmNdh/Dyqfcdtin5Sh/jeptNt8vbiu8oJt8W4RanlfZ
+xUizijP9J6znzj7liFFQCLKBejRwUIKpSc+OFzv/5VxOTOZzxZ+qOH5AjmDqLRs
34K4uUamkOV7C9VxtDrKgQjyEWnw/q+sq6Z9zk14RyQX3Qa5TDUD5i0hE3BBTDJ9
0+eP2oorm3Tf2HtfCCrmMn0w/WuiBKyo0rrErO70eJ/wTFdiKOPQiYDhtBynMnoV
34u7W4ltq41LXbUKJjuZH9PVXXkJIJ330MRPZ14Dg+me5hHDIZY7jIwkxI5XMEHb
WYdD2vviO7rUJdXnK20+KbqR2JKb9PRiE/S8qqolnjN/aZe7qgM/Ef9Lg5HCFCz/
6F6M0WJFkVwyAEgC5pZ98LT08rPYw8Lnc8Kt1F0bVcUuRIpHggme4cWYGEDFaylW
4jCni2cXEfgxSIvcAVZ1vo9ulCgbtSkjVof+Gw0FCA8bdO2/SAJrYIfO+b3aUq7a
yIT0kEQsr9jFV3DcYoOlirs9RaOAAoUwY9hWHTGeFIWp0lwLfXpvnNZ8TClQ0WR2
FjMV4kVsMqxCI0zpvOh++TJH5PTT80pv5YZBQRwQVrvOD2G1/67zYsYqmVfckoju
4Wi4mJKwb1Sm+u0gWM6uJorehcDo6X4BxR9si0lHzfAqX8LA7y9oXCE5Y9s5A7l3
5ywc6jhCEyKMuNXsEuchSkszckRKac0K4Q/rblN3A23gp8mNpnmJZohh8ck0EpJz
guap3TV9sQpASeRr0uViENHQN0KNoSxUNlhoqet+r32ZIlA2uElO3jUCED2xOSuz
iz5cFkwfwFEGAsTEwcCFWvxR6bl+oCheRc1iPG3PX2x0/1/7uCaR3wwMu6vSvpT9
y2YIp6b3B5E21YXj8GQZv5rVai06K7Zv5tNXuxr14YbANJoHmRtn4TjueBhjFL6W
7RIZk8Gy/eBSn5/BUnHQxXQ+LOFrk6CheSEA9gD55cwqYPyZNVqnAjKqmXZ9gwP8
8EOLS1eYFYf9FseT8FUSrpE6QwXc30wfDhzjQCJL5tf0uRtBt6M3RlXaUN5jIzzo
zwyczclNf8qhp7PTtS99AD4fahCyjK219/rovJc0QABOvCFTpOSaamjLvNG4XIbK
G2jPrmya9NRVJiyuOnIc1LPAVeKoqvE08RDIcWFqKD1oZTdM/ak1ybI+0Fxn/KFV
G9vp1O1mspVBeneND5CC0djEsxGcRK51k/VMGEPJl29lLdOD6UCF4vveGo9TkzsV
o4SidwToINe7H7/9u8E9F/RvbIDUQD0Ic2MjmicE2UhDOYJmkD69JR8qDuhTFAQ1
2sSMWOl/p1IAqawGU5u030LqwmEhcc22+5cgImrDORx3Bzy6X/+ytyxsiFNBn7fi
d+L4gMgCSCDNFQ88fvdmXQO4Ozsv5n1AfvGCh/LJfCoP8RFpEtKlXrnME3Ql44Fx
sYDLsEbEktZOT2X7jrcrfLghXGvldT0tNShd8EO3Opd50Vit7Fl4xFVJLROXx+Yx
kR1z2EpYeIX5/7Ca2jTyO7Nwsxby5YaQ1TJk+gfF4Di+C9CxazcYleTD73YlINEJ
WdjeXHD9VTfRyUgABIPE/sPb/bJ2TuLBjVwFHJIFbUVZyZR7yHaZwIUe0SW+jLZo
2k9T2CzQ8s+FYFrcBOIOT/VwfE1DhmBdE/ia69fvTcozwhxG2gN0Ux5EwMame2pO
NwylyqpFgOePirmlw7tJiBIn27kjOTXNsWQPFYrkzR4+m4HqeTEQTAEH1jueB0m9
r17GX1AZfW56AXCWgi0cVa2Sb+IbpJ4Wim1+Sor61prOXLYfNaWBVFCwTaNQM8ru
Rv087upCRo4u7q3CHX8uMiSsnmc+L9RX4gyJ7L20WPFcUIewaE0gkO0wmD2jBuC4
gGCAD0yPstOgAKnpaPoFDoHqG76WM37KfNRsOI7s/Fktk3rTAGQBEzyKTs1l5fk4
PJeckkPnJ0gg2VX06KTmLVlTfO4Xhu3DhUNCqHLuLbh+D9euoeZ7beklRML9+gNa
j59LmIruQZ/aqPz1wB0MIQZDcIl5k5W/SGBlNv+EAU3zgdR1/oya7118FiymBGcb
h9Q+31mrQlZwtyU3FEdGOPdAJh1oQh1TREh3jNsy6SK52PikG4P3ir9WCSe+pQmC
Ziy8a1krE2byMjOKw7SsFlOLVZCdyiLvPGn7BuQAS8pwB7cmMqBrv/36k2VWRuWd
kHcGbr0BAMy+knynLOqeM8G9nvnYu1kjoL5RpnaIoYh6FXvbEnl1o0rxzCnOqdu5
Ls6aGN9aAPn7gKl+7qlK5nHd2FLHEBbxG33KdhdvMd5e+sR9GCWzJnEf/z3uN0az
9q1mdQp2plepFBr7oT5j5MDxWfZM4uH4GkHDC3Z0LISCSdaabYNz4uL5v6aAW0M8
+GlARt1o3QZS/4oXkUS2jO0etRg469GSNlszwVtACLjy/ldl/uqn5LSdbQv7Ndma
C6t5/g6UegpIM2a/WBLo9zFaLCWRo62Yt/J64mJWDG1+WEqykx8KE+Ru9SFwMXTi
gqC9IEITuruR5nresL02Ah738zyPjYUFVzQTKhd8nOD+Pvdp5BAJSJRlnl/FcrXm
E7BNkS4BiY7o06HRjvsEqmQ8XBVHDDUIg/etCA+M3AmGNl5X1k8YO1GYHL9lEk1B
yWCNblirpB30nIwo4hRlfCooJEwE6P289rkG/rdzufxCEvdmC9CUK/NOclNLxPhe
NKOZKCGix+STFjDofwPcuulHWQAfIMKW1nns8venAWlRkthWK6dMtOsPgr0H3fjq
oUcLwWRJTYiZxCjuTfu4WcL7Rl2nOtxw4DfKpx8dl2KoGUAUhnPGELES6F7X85HC
j5xinmlHO8dyMIEPQ1X/TasZ+a1zoe+fNA4EtjjsXgre7UBtLEGol/ioIx05+e7O
Qla7bJtfQJQMdUQCtZdaVO6/yJypmdNNYl/hAttWPN8XeUNqSR0JcUhKoShd7q3x
tdhNd15DT5ugWlP+hBH+j4qawSubBSPlYBmNlvkTxJJnnBmy8QHYGAa0j2I+39k+
iHVOZgT/GG0JrGp0k71gPyc4hwDfy5HHvcdJFXhFbvK3lHIyL3eV4GUDV535Wbb6
Fcskpl+tj691pTpdyVR6gsIOcrh6KYUdV8CpqDlk3QEULV4RLGRqE99un8ENWpZ9
gBVa+c2cZd4TTZE2GpX8GMzPn0517HRgQCV2q4WrSaC+z6chyMgJ90psKiKYdPza
vTnlcP6L7jtAjH805fHxm2dsmZFKPjW7XurjySdgUdtsXbubvpKJyNW83Kn+V3EW
D7PS8gxSTv1EJDX4LbdTgKBk1DKz+4xLTgnVdHc//WheA7e+xh13iWVxGV4RDAWn
h5RvYHPc1E6rC3LMD7G79pUA2UsE43UQw9oKl9epCF1Vi6ELCbDSO/c9ABm7p3tn
Sl2EJvwIQw1ubOSx7+u2Th9PuGgj9OMPjvUevz6CfUK9i++o7A2A+v2N4QQGCuDv
4kmPXkeMOd+5i0xuVNkliOp916xPQeFOjn+lSsLjebPVIsb4+fjltsEXnUccrRmw
gJ3WO1bY1cIURf0n0hN1CcKreA0if7Wt8k6V6uRD2ctOyYCpHZ+LgSZH3X2FCf8V
BIFCBI5KO6njyw5dAKypzVM6G4C8e3QLo09DMY8R43ipVk9vD5+TEjvqIyPOZZ3+
hkTbxlZ9oqIvdrM4lmnFQzV1cEVlmqRAvF6oEXIaKRdY/0nT+pPL/OQhVp7IzfA0
Jydx5LCU9nnAoL17rRCnuMcclM+qT3oK0A+OQrbdlk6BH5PPaTLA1FGOPT6j1qt4
jPh0Y3dxhVCCI9AhP0uXkV0jgKU0l34VdQTr2iPxC6BaYF12HZo0jR8FETRLMhLJ
EdXQfiqH/AAq38aim7tK8FLvyjbvk/qifbkyyLhwkocIKtKSRDuQDT87Hynt3c5w
ggkpBikccm9n5PmiZRo0Prh5oL62FEaoEPyT8mCIO8h4Dhdikefr/Khfhr/lreAQ
0XuAPnoFe7svksrMWDp6C8onhIgTBoDjJX/Y6O+td9/8cns5SaPDP8qfnRG0voPT
oBozxYrgYqlUEFoqb63p33rjpDRT1qutzIXyi98olDcyDCh9c4lbeX9P+3EKf/Xq
pR/+G+MUU/Ew1ig29x8pGIWBc/L+f9HDpltxE3VI7IgryIYR073Bg2VUDQ0mODTa
9C/7/cucCnOQfR76bYQUJm0fZKK4MTyPIfqILDjPSCv21cF2eqMiC1di1PB4NzJl
nnSMjjL2C9OQxil7JPfVdY8DRf/onHkB/kw73DbFp89g/lm4Ak+KYRjGxqKFNSTO
jRwEupiO9QaCfTcSySSK4xW1aQWX4oRlc/FLFBlS+04BiRevMTXKlikBniRGXD4I
TxleWWX6/hZDokEW9gTg0Re9cGdaPnNt8uX4i/dHbzpThn2Sp/D8nZ4bI7xFXI+l
eQJSJWYnRmb1s5BWYYAE6DqY9a9UsjSYW63x3xdwMFisLwpWuzlefcBdy+R1UHDj
SxHszKLWm/i+b8mSKL2yrL7UGGmIybtuO/+LEFQqEtjoLVcCfHCDaR+gDYWztOkP
uwyB/mR1Q3SkakKAi5Lwsm1y+zWZeTzQM4g6WbF4GxzglSf/vEmzUVCuCluMlBas
0mFZmpd1SEMXQDjIjlI65+/wrVEwD46tmdVcRD6CfIaPuW5PTmTZttCt40LCM4bu
UX0RbkZ/YShe7vvFjr/vYF98+Iua0xEcENydcmluFdpFJaLdzYUFHWAVNe2YfXuq
yiFWAxJJ1lMUFLRJfU0NYkcNbG4M3lgk0O/OydBWwy5kAkfoUP2zQOY7BdYKNQxe
KxCafGKlDS5W6MJ7QVTK82lmk1OV1YUXRsv+xR8YkHRZEW7hVaIKKLJIoHJlL0DE
dhvRskNjC/EDJXYWY2uVZ+2NtS1CJe/SzOd92hcitkPGMwYuV37szXfd3Hzf2z2J
PU92K3c/qVz/uDRb4rVj+w2RRwZPgJBxPN5WXUzpbYs72tzVyYI1QTswh7bN7aVW
3xd603DnDVxcDEZKgp7kb9UVzeniuZ1yOwFzNzRYms/s770qJIb3onMFmLM05i2s
Es4nbAVYHQF+ZgXSVjdNuo+AGkARYqlES71A5EMUHRIfnwvfumMO5j96oapnkQwW
Pe/WmiD1oZARYa/pAZoimwpUupDornmDNl+F5/xIpV3s32Hfb1YHC6WB1JJHcEJW
WYJfIHI8jRPQ6kk3mB9Iq3hAu5cSRBpAQ901XdLC5EUfbU+GsPvOjx9osy3HLNqm
nQnz4cywESwfO+iBu8VuZpQFxvsFIWV+midYKJtT+k8+FJspkGvpuXBNzMcFuSab
4hgBoBf25Fg78pJDH2x53V0Pb4YUQmzo3f4UHjjd9F6psPFIbg4rPfWjJS+ITxVd
BYxZJR9Ss+/0FGDaqq9VxxmjuEY+wfes/u2GpnvoDykSdn6FkDxPB6/Bvh0Urgz6
9zxosEWKuB2ndYli2B+kGX+dcZ3hu0tjOv2HNF5uRJC8gEjdP5Kd0deplDhqqjn6
S7i9XpmJw81ioCVTSt43AfOF7o1lqUYwywiPCi7Nf7OkM9ppSM4duAx4xDF+DOQ3
tVNbRn7FbTn5y/OK+1Lp9oNPMRJGkKXRr0V099o82ZieU2zupidzJzO25rSbW+WT
YQnCZd+oxOvrBzajXXaOxrG/ZziwpCO/YULgu4A+fNr90/7juBSmWwRCSqvm36vP
1r7boPSel3oczXUkqmFvybzylEEevKJFnCswOJ4MIIiVA2szr6GzEJ8sx9MLMB2X
AMNCmS3bI8k7SKXNIkyp9Qsts3tFiJgUsVlqTxZZPdI/WWzKBwmEX2/xsZECwsHM
YAgAP/lNp1UMWb/ozTSsdUlhWDnNDAAsCUabdnAsPnDXODjpNbgiI3Kh2LOfwvXT
wy47sDyQ1p1Gn//nLipEkDuk5puKG9ISuU8SWMM7CnnSKRkgrOc184spPbhzm1Ip
lK/8nhNlf/lg8Lf2QZUMzifgnKdJvLndfEckaw+taw5lAvvKHgknsDwQKzyNRWFr
VCToZIQSkHISW499seShBZx5BMH1+kbpJdB7VD+hnUBtiH7xbrKtEI+8sEpMI05c
PRHE+y6eVQOOjvYvc6Yu7TglFxnI/LiBwhhd66rHS0WIqxI0iEo/erpCON7ZqfbP
APBfHCNMUDGZHFXEtrug4dG+ayO3dxtuJseTaeqdFmeWX8hTFofQyQKIg8oFRYfw
tD+Bj/b8UrVPgvvLY9orG2l4Ep1Z6/2AaBI1hl7qeamP6APTv68Xc/qAQ6/PB/4d
2JiG0wCgLPKryG+uhvYfHPD9t5JmzaJtpYKuvJj1BvLvzT9dFnic2yr0PJjNHdow
Xv9l8jer2025DdtJ1r9fivd0H0Q+/Plzc6Wg/XTYREWHnWoA6yNW+jjf3bykfY0g
NucTGOgLMkryL7oyB0bJlzRMfmcY/F00P7nqF69uzDOl9V6toAAMshG0rI1z3sOl
AarTd52dGWyGA5dLPxBLA1VN0IbO7Q/wgJiWlxs9TFfghHf8rNf4adudwgCWn1IT
s0K96X47clqWRuiUW2eojPKX7CQkfZ8daZUCJ5PcGAfRFyfGdpfm2XetjdRPdDe1
kl0S9K9o4xzbsb8aSd+QFMPK+LosRc1HWd46JQxhrQ5pSREaQcQB9WDRBGJuxwUc
UalqQTgPXOAPvewAlGCxlksZlFw7TQJnGBVdYl7pOh9Q2it0XAeQl4iGVse28d1z
ivqlwiapFcHisb5C/1IlNMywi2AuPv/RA5TNOGG0H5GLBhhNZD6Hy6MtjfEVaiL5
/kChjGhZYsvYzE9W9ZceYfEg6HAvP6gG1oZwG/3PIpQlwnkc4oVvrE8wSy86JfH3
+zW8MKbLTr1XnKMzWQVAKhOrme1Y+mx4k2OLMYACM6QcGaY155lvA/NJYR84ykin
xt20fwXBzMz0eUB+gZdYBr5M6ULfhTxT7dtY0x8ELRCHtYpEO3XPv8fb4pJnYTS+
3tN+/XZeV+F9IXt3IBx7RpK20Z7iu5iRIOiGrC3CcTewPHelPwM2z74IZCCo5VGG
3kImnuYFlEyRk6kpFWxLuS+77FDOZuM+36upxMhFrtSODr2Wos4UbCdCZmn1nRZh
G9VknnF772FdTVLu+n4HnbDW1wDqSROOCTsTRWEiKxnDv4uuaihahG7wFqmvJDG2
88FlfCeBu6FnJ0ADexs3+O5L10wcG+MKYZ27ODGcJgVV/D2AHEYMmx+PKUWa2CXF
2NuHtJ4eQVqzgjvCDptVM7tyL2Rm6w8DJLH7iyBHLSAGPJYrnT4u0oQhSjh0qod1
H2jRcd6yP1rRkU4LSWezofcYagZCRD0YTQv7CkG+HldVQR7bYYfjHXLZKcddSOWi
YZDHlWFKHeIzFL+Kyktd2s24YnPlphx1b9rEP3LH1CrIpyGq/25/B7a2zwej7Ijf
U2p6Vabh4qX3R2zdhnNxpplJYnC6TIJ0i3eDwyFeWRNnrp5mNjMnY5ZZBpX3Q+ip
zRTDELbC0BnMyKM3+UMrNGM84C+czhYAQbaF0jjOxFbkxkdM4wDuLRObQGysRGK9
JBtOGL2NNXD8S7mPn4dtMBj3+n/DePth7wJuvpZ7BBQl2Lo0VSVYneQtppvcK+Sa
v+1g7DN0dTmF+h1/kEUtu9pPU0P/Hesr7XriQYZqQExypXUPJQZyb8zxh7sOBd3P
Xx4BXuz8C1YGxOhJBJXp+olJV+35GkFQwU0iLG0t54FGQyqO10K1qD8IL7RQkkvj
kgHyUOVesiALTbK9lAu5O5eF2B5mUgMBraxXXze9M3kUGONCS1SD6vO/eRDoRexw
1NMQi9Fv/B+HGcT+mcFMPhX3G4LH1joC3ozEegNVm9ijGsWEWAKTV85qJOj8Eh3+
BKmsbzIQkT0Ve+6oarA6vFJnHKgnZ38V+r81U5+8NsgqFiAgjYp3jMK0aGB0cHtw
VABGJsmEZL550EeMnSGjkWS29AHxx5m9S+ru5jmnbe9T066yU57pdOofOc3XIQ/e
6ch1iliOWc8atMDLAi81Ia2bwwDLDx1tUgIFQm5xd+FwTW1pms4SEGpEJoRC4St4
PrwzQTkvG6jsWpbP95+a6tASze9AVbrsG3GNdl3XIOBIQT8dtQc2G+lg4qFLbY1e
qU4nCbjHmf9Qg4KB+m4A+hwBfAEEzBWc9D1eOCj24NyWbw783x6grv4NTDS1qzfQ
FlCiQUw4HP8LUIjinmyGQM3Fzf1MO3V52sRGtlQ1i3UpogTNRhJF0/0tTUsrVky4
jh0wR0oklYHGd5p8Xbv5bw/JXHz2VJVsPreaD9LmH71FwtIDPsjFNBEjAfg3SsDa
c1vJbk29qabZ8DOTDC5J1LEabcvDBfDE2uwJP1pFPIkj4GFZ8cTpj58w/y6hej10
Xh0F0p368j9706RLZjhmH7dmBdZ8oR1BB8hohbJ8eQHgc6H1PFxrrIT00GQd92Mv
fI7WZp5yy5jyKqJq58sl4LFVA6KCyN3AVgrNVNlcOf1fxAhJUvyAZdG2vCl7KOQO
S1oicDCxsPI6/U9Azo6ZsH8yjDR/JFTuL1dF14F/wM16szlagqlYJTCaZa19D3WB
F+u3vP92Oqf16n2sKqqv8ezoqB9Zpt4aR0seehI4fZ+wbMU1wHIwviHop/EhQ+jc
vctk7Zn1xVa4YPC4Hr5yFImpW7ZZ+SOigZaPJGrqBeU1HA6OTnJZ5pxjGEwKU/jD
8ftrkwQfoAhvp87RHZ9GNTRbZ8EI0VSH2Wymwf1/AOE2/rp5zyMbFavNRxJ6p82C
WsziBqYFmUUnY3JLO7hLy913r1mZGuacVyqIiMOq9FZGwjFRy7AKHy+5P5Ghp+Rl
OREFe3L9R85LzPGTHrnqYY1p8rDrEWKl0/VxHoca0wrFcp7VL6j6OHI3CwOPlp1c
QwB9bT0PvyT3n3MhzChhLW0hDfa8I+sQfIGsKleItEfwJXxN6uDADtLUg3wuEIGA
wjxZ7BT/J7kq1JurwuVWkj59lw+ash92RBr7lmc8ApNmn4zMKBk9bv24upa1hwPL
rOMHfBGtXnhNt+MzeEKbcPKj7XiMwzZNAi/n0LUu+OmV2XJJ1HBZxIBbOIyuolZa
5lmeToR5erQg9I9rPXS+dhcggZbNM8lB1NDQcZEcCnV3Ogh4ymApAh7+eMqWhTjx
8VF3lf4qcZfb/4UG8iNrJAl5vGaVLs4qn18mR0xXHkyPODMDVNrQnox25nD3wuHh
3bE/Qtw5TYZpEc0YOOIBxmFOJlrCy82gq37HOeRpJSfl434VEL0OQhAwOJhxAKFF
kRT01w7qoeqEsz5J5WhBSX1VfXPUXSipoNsBy0EM36RsHZhqIQymLy/XCLN5/QSS
sGT06Ajvundmx0CtV2zWD0rgEbndsiJkhd8zTiD+VWym5bjEVPP3KcNRGrqAhiHR
u2f9mmJ7HKYCHfNAlwvKrlMHC9BinSOtYVrYI1wd45VvUzuEh9mSFBc51uO+ayAC
WBHWwB1LFvIN8hzAPfkK1fHRJxv3k46dHtB13/NK5syeiYm50X2ykIV2Lc9w2Bgs
g5Zhr+JJ3REWLeKZwku5Crle8fKudl2uXhamG/UQxdb62HPeCEG0U1gDsUFIdqgy
aVHHgQjN6ffnairiEmb+iLjbI2PyY9PukyLL3iohp73+XNNni63OaU6i2xIlyZb2
9LI8Iim+wU+PiH36gGvNFTtDfoBvqdM8YDz1AthgEFA0e9PR37azuOV5SXFzXTlA
S+vYC5IaLhwiJFU1nOyU7nL7ByeO9EZSfOhpsaqYWz0ZZe8xf6p09mIzZfCza3Jh
IVWk5MOQV87/Zi9HgYFJq++5D70Sykpx48KmI15xUfhK4rpQ43G6ZWBUlq5vOiXA
JohlIhXiVhnX2TNkEgP2SMv7xSesdnzXpRji4sWqzB6cD3c26N0gnS6idd52PzxK
5QxnhWkAozPtu7g3/OYW4G7g8bwF34p5Adn/F6BwqbrNXuCvR5dEgHfJ7s7KENGk
3+UVhFrFNgd1Gih7vgg1NhU3TrSCSayTM3EFcgq164Y1beRWgyAvXXBDb3rGh8TS
jQvDz6kg2axc0ssxUasBX8IGUvXcDvpIAR9vhr6uwvDvN4Gp37ytUNGQVoGbtSy6
sxE6h9rcdLbeDmODl99g8DTn1rLK3oecjsE0pFpXAMuTwNPTENt76mgbfMZzWYUj
BhJ8wIHDtxlaQIaCRf5MNuW7BPLP+q1zoflwBytTAA8hga/5YAJrKQb7LqTywuyj
img7Xi9irknrIjd68/H6gEqtmZypdqNswzrIc5Rn9/RlJ+CgBmPqhzcpyUKPeVxd
EGTHACGVYnbgZB2gjF71xbT/hMs3LgGp7uLWEOw7IgJZVDhp4Ka2ZHWZcrhZd3NG
FkCBrSCJcMs/XgsVJwHf7GPkeA8j5JMcXgD5dpWQTXQypKJYGyGbQCCGt9nBmi0F
KIoBIm+vFz8jqlnaYXdrDNgdcuyPZ7FvhM4USVqCwseGYDDbqBKeJVvHdGUHl+BC
yWF3Q9BaVymE29UY0pgSU2ywXeRNR544YqGbKgOb/W6dtKV+Z0SAi5nqp65AQR6o
RSAgdJ+HAn4KVPV+SQbswZU4obuo6i1EOSQ8KRgB/Lo7/xxpjtYKvJZoiMXZUcfG
QITUMsvRWRyfZvsrl1a/GYkMQPR4pgyXh+zOHr70CXRfX+zp4mfc1zKrWjE49cph
gbnFvs8jPnGfWdueZaqtbH/OBla8f3Bl/S5aQWh2RENPPIVPc9Omm+dGaUt5iA5Y
N9XrsvQnTmYMX4+YZEd8w+dZdqyPqH5DttwSWaqS3JwKFKmL4IPVEOyB0m/Ds/cr
qN3olXS7eJzTNT0G+dBXoTHFIog3HZVULXzsYrpFCGP1FYl3KdY9FMSkVXaBqIqA
6rM0UhsD1ON3MllirscAES1k3sSOhOggye6uNJXwMUvYGe5ud3HnzJOoV/a2KP2Z
NWfMwrie+nZ0eTmG2POVyHAwSUmXOzNTDwTGeLrreCOMF2I3JFgTNK8kkchbaXjJ
f5evMjB4aA442Dxx/0bahS4yLrP25k5EmMT4J5oHegyWMsicDSKZFF3m0mPBa641
HkW4d4Fl5l0+KtEr8R8dhNxqJaUevBoinFjWGLpt/3Hrpdu6ZLI3hsVJ8CrbBURq
wpzjryTVetAQYHDAjgQmGL2I1VzSpnh2eFHT/OxGJcao1XIoNqIDyWAjwPqc2Zq0
xIUITjOamPOst3SsfRVFsAUfwXd7MLWX5gkz8AS6SDrzNnGP7pkU1tBprDl8k85q
ZZ71ORlMAFckt4iGUz/97nTylDKVPhMzEBnWcCLFBCeZId1cDJAau0sXn6PjduQs
DiPhHYpNp6dFn6P3aNeXNjZ5Bj8H4HoxnAvoNo46bJVX5YeUhnldK7a6av6Mqf/k
z2uuCVMxYV+tBb31QgRAnQ99SwuOvuN9cqwgco4l5/iKGDRL0RMRBq1hxcf706vb
g8XDwgcBEIlJ0Qomf1JUzrO4S2jW3DVUcc7TLWGi0PYVu+74fuZMR5EP133QsfOZ
TUXG32O2FjzgKNjgsiDD9Mh6DAgv93rMhYFGaFRMKq2pa1B14x62cq+VGQIBLKIE
V+Y76rUfqnZ4vdMufv1RYX/Vb4ZC1Vg2apHoqZSty1spdwXkvacxMxfV21ezzfWU
jRXDH5ukcRTJT8Ajcsk68iJNuNbMKr71B/VfI4BWBkbfYDyGMM+7mSkgqm2x8ez6
44PXsjmKrhF4sR9hYri88zbQpDoD/lNkHYR+SjclqTYyCwjj8wvn5tYrGBhCdQm0
86UakKskdevbc/9wjwN/n3M8IcMxk5EjiLeGBLDwwCN+SMdvfTDZpKmzjkTY22YD
T+CEzjqypQw+XLEOhUrRTbJg/7ETuL9U7hrGyXH5WnSR02sdhKFU/PRicHmYaUJf
VTERNBDV6UdqUG2qZa3+HLwZqkyPzTW4kojlTHdwEYyP4FajmPO9TOKMSyaNh7dG
Idej45m8H6ZI9OSEoQk1Ile9QekTGMVJo1ditLZPzwP26SpDRRTToU672WD5cR+L
hZjUWC97czbHPVqk+5qh0nRQgS1vLPc7QUlYnXxQazol68YZ1gNJTBUwCesIBH0h
gfE9salWma1jBY9IGKXfo2c3glrqEpuY3l+2P50r50kmXFm8FEg7noCBLoSKKspO
ffEDKkjKws8ZzNyWRloUU10ZTYcR9e/eawaD1DOqDumk/Hyy91Fvm3XRv79S3SJY
w7SjjczM4dI2fAtAG+pQklBQVXLnGyvi7VrCvhSa4aLHwcDnYhbWU+oSclre9diS
gmOJiPpumgfUX3SW18MgSrWbWc8ypFvEs2K/mjfDhEGfZdcIkJPJjEkk+XNl9E7g
vsZPqCpfOS41ibopvXlLaecJJuoYTbW36jYs95RHxz6k6T38ceZgb2HpZ5adtfoL
a3PxV0JvjTvKBjVdtUWZHlC30QMklxjvrVbGnVjzgmsI37oH6oIGg2HSdGCRGGIt
GhTTgMGaoh/88w5dUaEpxWyfY6zgLsQNlONYXoFHDMJ0fZ0ITbGRecAggUWnmWSX
eqCd86U1gyg5R3LlrR+uMX1etJMRq3HHTmRTc8hX+JiLIT6mL5T23DZPVXaJwyjp
m1bI6dLmvtv7cAUhPdTPzjkO3Bfayc3AJDu1OZyleELFNxg7Q/BI3VSwELtE5k+j
2MUUkd9bL6S3KyoFBW5uBHuH9rZ7qCYWstRkjvn2rz4CJ1B8qJI09grS8LB3otzt
0rtQdwN7vox1o/Zo4CI5agIB3rU6o40a3/8jmmJmPnKyqg+SP7cqGKFG8zFgZ3aO
0a1yHx3QMa+7LbUlXnR5LbzTpoTyQi460/HXFHLFF5Kp4yTM1o8CoyBgwffKF6j+
grpwGwB/FxaBpC/f+Uisi/QtRIzkmmC4PmpZYIx5Zgy3ZBpvEkB+y7xo6U5Zd+IO
WEV4kNa6Gkwaxnse7pjcGenGqOkShM3Pa0zU54DxITQ=
`protect END_PROTECTED
