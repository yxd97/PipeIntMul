`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3liw/WepysDoxl18fG4OY+sW2OpJqvjIV1lnCoBRqyf+v9+Coi9Y588MMBZcMJoy
bBPUswh6mmql1FVQykHndFHuoKPac54s1465NI+SuBLD5YwRzBAUAO/0x9tCqIEl
diVwetnJlbLt7onthq8YSWiM0us5K8wDhW64rczIupvv9XfodV4DiGOH059Hhawv
0wflnlrGcX4bHB5Xp3PFriM7paX/Kg7o5ZCOIiqRkL96k562pXwfuGW4KOKXoZkM
C/ePaFQiWXUeZnRgrsHdKICUstVxA0tqeDV0AVOGUR2aY5T2sF7NrmWHD9XpGU8J
ptcrrbO0D5aHafCklqFNwX1DigemBYPZRIXZxJz4/1qQmBJKIbHbxybORy0wf4KO
Pu/EdrWaqWK1S358LSQjKbUjTfiL8MJJ51dIblBHwhS30OjXL2n5dhOuEYAsviLQ
y/GrFRjkG02845KKPp080yJXOqZAL+9/m6tmnmQh9TI22o1wpmTuZcISLQ7K8z5+
`protect END_PROTECTED
