`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RaNlxVKygCxf5yDYpD4NM2P+t/WSzduwig3WI+edDiJpMDjXF39WhEwlEMCXzrlT
5FgkaSchA0TO5RANAdyf3cREMcmdxVQO2+maPNlMmOSbEZXxetnIO+14IdWVhA9X
QrHcRXE/5I5GI6nAHMd3Ih/KqzefcuhpGk/KPjt4/237yReOoahjjDQFx815ICtY
ihurmS/PlbqBpQbNIePITFFMoGKv6Psnl3AvZGoZJwb8sbMMXINn/LGjCv5Pe7Rv
9/BWPt4h/RXQWy9f1xsYMNIsYkZhIgr2h/lntQeTRl6d/fTXd6X4PLSq/9ssEhPm
RjTnozTCWbUTgCgEp5YqM9FVEwRSkX/KiPkSdQZz3BM/FYHnf3Vn0U7weRSvjSyA
i37pad7zWEf35oQZ0SWKiZiIBePPs5Y+8Fga9/MnxiEJ8w/D78tw0c7BHb1GE46/
9gktJSqap9KNEBLaniEIesAt7y+mfYvdMT8cMKpDxpSHqEVUAJp32QV8QiYKNlx2
0Q+UVyvdkXTClx6zcXamiyR9rg2qoEu2hgp3gZNy4EZG+rQYoVN0aBh/nMvzsZBZ
nwc2LR2MiTaN4Xu2kLY2AqyOd2GiIDBKOZUxH7ck5TA=
`protect END_PROTECTED
