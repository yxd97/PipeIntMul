`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wBxQHlu3qWTv98QhyQ+k1gZX9XmQtFY8CWksw9DxvB51kQaapS0IEb9goWnoWyVk
NpozayFdflaizedqdhX3IjL2D9xL6c+qjN9od45zs9IgSs3pCTWI2FWPmkwTopWg
q2K3URQeV8BCVP6XXPcHIIJpW/IxlgIc0xNPYwFJ6jPXmtPe70fWuYPub6j2GH+j
IcfzImi88Nk7ruhxdVcCc1etawDGa404+U12ebxhucldsD9gBoMbIzr9chlQUzZD
y+FGsI+k5iAssVAykHhkwZLIXWhk3eWAsafh0Ox8o7xucr54JUMIevaGkJnWhm6g
TmeeZxuNb4SVkGnEu6cKiQ==
`protect END_PROTECTED
