`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypwfpvdFJtGI1D7mhnNQ4Auq8jBCKhwDr/17Xc8Bh7hSKYRR4tIFJtkonoJ6e2tW
gPy8Jv6bDsGciVrOByN1W1PmmT569z7PQnL7HAHZb9WxoyzTKLmAeHgViR0IwKPs
1FLuRSJNbustO/QqVLX6IOpldzYikFTyyhC/h1DlmyzGn+7t4jQPpGfrNR81vxe9
hwktm/3F6lARjkaX6ngL8Tei/tcDrmt2r1/F24xiID+ENJdopTiwuJSR3wXnCzDH
TV7V9yWNVGi0U7aAHIPDt9ByYP1/kSpmnIwr0g9133BkDb5FIJzCQALRXpis0Wjz
EcXnZCSNhkv04jAZLyIFSWS6BCKbfNpXY48mIoRxkebqHddFtKsA32vLI8nUfPb1
4kb2VS76MvWXqYPHom29zxVO14NPdr/OBVRgtD94udw=
`protect END_PROTECTED
