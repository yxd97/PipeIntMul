`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zuwEhDUfB3mMUBpAw0admPhoYC4kuQQT8464XSMSBz43ZiMkfZNrx8/FlBLAqdcz
QSO08C92mbABYpA+Jc/unbr/a6fYIPccZHTdV2hWtRUQdtUBcWkRMqnxoHBe+eVi
nj9Jpl+n2zpUX0mJSrF82pBdYtFl1dAEUbCK6bqYSo8Hi/M+CcaQwv7mzwRbzMTH
1bkuzVfMrpVa/qtmLm/gdt+13L6paGB/tRhGuNkzsi9lMgO2I3yq7ou8KbLqCc4C
o4+kLr0FAq74ML/z8EncEuJ1NMhTU2bcDHWe7+LWwD2ZBP+U+hjRomOg1Cwaoqgn
klu72wNNhfmTc0KuI4Th3FsGRBhEkjwG9P/apwBcZT25DoA8uR8DqshCqQBKvgY6
mp7WD11O+mLNt6L2YhywNnQ2LLn4y0yeypqIggb4Xpo5zvS0VskDkMA+KmLKgdy5
pD4NOzxKeGAIHQnPCEfIdQ2DuLUph237TgBP6jrBEqNA/pgNz/pVuTJJin2OS1Y3
FN6iAraByj6eD1eNuDBuqTuDadioCWEiRim1+gpwByDdlR50Sxnsk/HFdlS6eAAs
nwhpK3ze3k426o1xHk/0DplU1nvskucXyOf28NAmqPuthSooZkT++X+fNpjCSY8q
ulki06cKYtbgmU0SHh7w8lkQXduDWEHpUm+pU7qXlc9Fg/X09aVenaCVdGsWHWsX
lO5u/lCnauGC9TzE39nRRT0QuRGE/lmASh1CJEfKUmni7Fy01HmBLOxRHspHyd1t
RUAJPCSwaWEGcqbuyNuS9YwCPj/9rd9a37UOKuG7VxTUFTsMOs5n1pDCtgkXKmkF
KqetIR3NGRxjMiGiWmxtrQKWqd4mryHFKuZyHocCV7ZUfQbd9poPk8JtMnSLZNqd
y/oviBk1NnZHbb4a+Cr9zZfo1etmpGfHqz9+Y9YLIjLPPWnF0kYdF501vefEBlHH
`protect END_PROTECTED
