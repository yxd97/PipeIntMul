`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U5BhDcSFxBZgPqe3Ir0j3ZjlL+r97NxHtsYhZb0t8Et0BFwvxO0f0eTIzbskCfvD
xHtXU0THE8P+wWrp/oNezszZhVhsYBH7usUz2WCWz/FLdwzP0h73u8LjHavHbfcN
BF6BoNIk3QUpQsDsPyLSUbswFcEyDEUuJ45EJMyXAA+BE5hYfE2FN1T920pEuOFq
HQP0+w7qJZoEi1HQcYOlGM8YuTpTJL0qQRJ2E2Far/We+riBw6Mbn9K5c8ngWUbd
Iupey/rTMFurHLkWLQ5wyVTP5i4u+vC3dRHTu+wvXjKiVxdsyk7+eAm92qirtbLJ
5lJS3oxRScKZlTmVR0ETgasrd3A+yqs5d0lguc/KeYZAhnrLgg3HcJ24jQDm3FBy
`protect END_PROTECTED
