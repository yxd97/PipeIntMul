`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e4M2NP+PQln9Uv4yTeL8GTeTpHMnxQM9iBxUFSyqVP5AxQGcSD9QBzYd3aYTnZlX
BAu5zPcuN9lTSafBGWfrUmKKYgZi3GmIK35L+of3+3jUm322YB1s4cYk/nPrp9GJ
TPTNAdN7IdvnIpfLQ8ML8BE2jieeTjVwGcEM4+2cPkFNWtcRP97Ok4NUkfq4pcHn
7Zr8FsQ8ewMQMzyLW8vvMyUp7amlOKfrhS7XQ4DPIj7yyaMpiyKr1YJ/rAuSTn3J
sdZcAn4njR1RBNKX1ESVB26HSYmXTxGP8nNhfHwVggtT18u2eR0Fyn0yWykCdYdQ
Ma8j9gagoiQZsMX8txM/ugmpsa3Zj+zlulhwB9hNWjfVTTObpzzIbpCb4Xhe3PHN
BKChMNpDpOXSBlRnQv1jrmFHtqtlySZuVZ2gTxOzPp16Iu/9r9HysSaJ0QKzPIZT
Bw7pvUBH9c7tmjPL5TzINyXzPrCq+dCzCcQxyzNjX5gQ8DOSudNKN/RyfA88gS2D
TL3mqRWWh2hLO0m5t7EtcadRKSFhCt9tuotBshn3dbsvW2YB+Vn5DDtXHTlTjp+v
dX/ViaLO/MLZZ5++bzAinA==
`protect END_PROTECTED
