`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t0nGqEn10Kf7t09Br/QGgH3+RmCOoKoL8XcH1JvZyf2KaDlAPRBEm14biQ291LR1
K4QbFmNNRMLX/m1nRXZL6BN/cQegUZW9Kni8J4mI4boowEUCq8rXntPchSvDxN5f
UiyVCSF5aCAtgqWhsLcdESaLuq73Ie/rh9yqI3EIuXEmGAh3bNOs6M4HWlO2bqzt
hsAZPxIaCu0GyvZb8CU47+KlVnn/vAST2xIlOJ0G5jXs/w5aq5zz6vbn+YVFx75z
mbsxzo/iasgBuETHJaccHxMAFHloEZUDY10ugGhe1Ckx7CHR+grFjmSeEs+YAT5W
jXby7pVshzYLCdY4C3y2yyL3xbmtkPpSpSYIZ4wS5JST6PTzlI/7aZji8iSPRSoP
NLDsG2aEVsR+P9Ue7CrmonmA86kdtGAWvHSLGD6STxtgdDs6+/M9oSy9qQuOo4DM
Vaut2Dzhd5YWw0c4Po7BP91H8QPyjEYdHmnOjGo3by5kKfjJwqVfs7uxS3PXnj0L
7uyE+3V7VCUlvF43tgCBpbmSNDDAppoAz15e9gVh3oop29x5NRLKlXcp70x+g0qr
E/cwRG3Daai7NFIB2u4+IDEv30YI9evYuMR7tFP5eNA=
`protect END_PROTECTED
