`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bPyq3tedYdW6Vf+FmE7Dr78y53ONRvG4KeuisSmsZZ/bJ2+UrfRVCKfMha6nJOC/
Zjb85tki9ccMn5cJ0mmMMyMJymlCGZknI9mnTFh1LmjmHBGCA+VMoVuGv27KbDTG
YObsUT9/taLj74jjYqQEf/VIeH1RiPWrcjUkR7neW5TDCGcsF1m6rEAmcDXlPH/R
n/qmr4h7YUcL6YvSDdcMpr6DAXCpqMLIWhMytJDgjyw+4X9ETXn1buG5ENxaD19A
yevPjDbq0n/EPD0p+es/LqHB8UOw83IY2y6lT0/C2lUQXxgnB01Zy5Gsa6YPTZMQ
op+FG+AiqchtX/e0qtHngG80S/IfXJuLucRW1lgLG2fM8skWvgeUW2Wmw3eDW1vB
St33Oxabs6pLTkdJlvQCr4XpL109AgnbFmyAlPvDhGV0LE1736dwzRqa8AC2QMrY
A/7qEoVSJLdp4CLu10mCmTEu/ro2bRa/NTMCG88EJZO8x4MR1HIoqPK7lT/TZGVM
TrWlkLQU0vRUPoHkWLVcX6xWCv+/xOrTWfNGrWm2iJO0IuFfHR2RGX9vZ2LgIb5S
K9jo4sDbMHaQxKNFFPLBEc4fVm58krmLOVrS23eToz0tzng1TNXKj5KueLPuj72L
gtF9zDFMz7Lcfc2Za6J4hwh4LWW+0bl/3nBik4k0aKIaBfXvWaRKxZ4Rc5UjZ5j2
eHmnjW5DHCaeLlOw/2NfttSDx/FnZBxu7o1kjKtGxjN/nDqM9U6+c8+thaMkmFqZ
frXUWrdga6vTiMhQDeCXo8UtJWBzlCp3ZlHL6F3Jgcfl95wI3odYe6iX67ct5pYQ
zSN4pTqAeEghn75OY0Ouy2JC4IMFZ9xZsPC6dZODt56p+gKEixCvCM7YqkZw9z3f
ARaN19gDSBLv20n7OiiOTxHdyyj8P2WgloICZ8mC122n9eNzrqFoiPG26WYXW1BZ
qDavcfVeJ4njyBrzaZINw88otFlxVEFTSk1nhkPO0Yl8ddphGYh6q5hIettP2++g
FAzuhEAbiSrSCrzoWxKyKBJ+PB2pQ5x7RQwFud+vPl99coBq1+O7FT/KRh7WqoBe
i2kbcEYa4iJlxuUMOmdNQZ2nLuOVoDpTqeE+SzDOGpbbrc4N/MjZ/C6hIGaNAywc
`protect END_PROTECTED
