`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mN/IEZCvxcMk2poXVL2ropwq2dQ580i948ZGhGuABLx5eY1+g/I1eAPtwlnW4yBS
egIxu+Htg0WTcYSeiEkET64eBOp5iq/v7MzcSYIAu5X2xYxmEulITQfMPzCNlDAc
UWfyzddv95jE8VgF4yHocYoqnp5begimEs3MJGI+B97im5911A9RCkdAPzKA98EU
adU5VQ8mvVd+a/jpvVA7qf/zSNdr7m36WTk+l+NuPgCdgMy7tV91HDAJR78i/reL
PEU67Kq9gZFc/vevPmc+dBz8i+SqHi4hvTfDMnGB4eK94enIVJsyAs1558zOT1Y3
WUojB6XY3t78zYWGEvvIyT4YWq1qgClcQK1i3aDgI+joZgd1ivLb8HlrdBMmwfTm
`protect END_PROTECTED
