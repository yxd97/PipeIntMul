`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ASw0RSg7gkIt+eE/ePqr2zu3nnEX/t/MonXpTELPiXmYOiqhw/fMW2TDemz7T+3r
1ssgRIA9C20BiL+WRdATl8cDqkXAxc35QK5e0eqYKuDTrnBvpxjzSqwumehzbIql
jQ6IoSu6iYBnd4EkiHEtp0KJsphr/I/ZK3QjeSgj8wivlAfHNMBpDzUWCa/8IiUu
m7ULGSmrCotpBmmIaZP0aQNMAEIn6ZxEZSwFzTJ9AvxQXRCzACR4GxVavJfgtsAo
QdfaanB9ZP9jlEjq7fIx+ZkF8FPZcuvVE6HxpDwKrgw=
`protect END_PROTECTED
