`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AbcnS+b6oO29SImw1dhzRO569hxxi6GLlxA/aqp5EWg0QuPpJJpbFrw7DCmT+rpu
gt0ulTDD/8p5pPE5CupHjDzBAt5DiJwCR5K7UcQHLUpd2sYoLc0wrKACu/WJQn0X
7prqt97wYR8mRxnD71q0F02Xm259ssfPWeDpC55KGHeaIVBAT6+AtQPzV53oK5Wa
jVWJamUxHlAQHA5PU4iCUfRErsnGxlt64V5hqmLW0dCPLIDAgWcn0DuUNNXCMc1p
3fUqRYTmlEfSo+gJ4i5653J+R7b3DrdMuENa+/OBDn/EVSzZYdEvRl9vV8dUq5I0
3lsU/JfO4A0pJTLjUvagMlyGIMfMag14zySzwWblXfoR3Ox33Jju5VbOw0+oXXgd
1M8x1Ly1dC3G2eCPOcc48drMJZfParZMrBHTsNgCI1x1sm8vh7zK1o803f5hny0Z
RrOsYMeplfkC11WsyQDDG3GMvroYVi+tEvCfXnMHPcNyu07kJsJ8nFcAdHCFWZNF
3Gy4615Op0fczeOIawC1V/94vHRkgTli4oghwBpTBj2KNLsqV/d7tO/jHvV/NqPK
ibWAEDSBK3eA2RzFJkbjk505y+kr5kOyHLWRMQ6pY5QSJrhPWv50AwdWqxq6IR/9
PtZcDU9/WLQmZ8f0v6bJJo0PoroaenmSOSoOnLI8tO3qWgwb/dtIRfgqmoqF5X/q
ipOOnmDRnsUpmt1iE2LIxdIa40mAgUnoJA8mdRi8T14qzxR9DgKPhYPHLjI6JKnm
Bty72B3fYWGam3zxRdLERk/LA57+jrk/eBbTPNXNaJUxK97kXeP+hkpIqrps7EtT
dfFo7YKVbyoNIkj+/wyrHKOAilB5cWG2UjgyhBtL2tBYUQv2jXjKej+GW8uXVRIR
8Uq2synRxxZPnYRAwXfRBpfBzJHPpFlIAcJ7lDkENezxQ9dY6xYDaVvAPKUsLjYt
G1p5lqnWZ1BbJSg70ZKERVlYjL4176SXne8TP1u8M0+aIM8YBXBN42C0AYXWVM2T
wTLVSoUNeikiWGXbzUC2rjVulQWcYhS3urCR1GuHzoyAyHjlJS0R2p5rpRd3zARR
guilhR8flmDNn+UI2oCuMmzHTbIWS0kYS8y/OiBbkbUngSxo0pfQRZMsqxsoNRHz
dx3xnRTU1G8vwG+V/mzbD92desLE2h3thv75K+LwrG+ttpOLTeDlOt15iiz4AxHN
EMm4uLD9dYrW8EKsKsuFTtm2M91yDtpdSwDmlHrc5LhP1HqLIkvxL48avnXbCC7f
0cfBw23vzTTUHm0EIAjriB6lnd4vrIvAAXTThr2S7y/L91nCIpo78L3T4UmrwbVv
EN07WaaiIAjHIcvUatisAYauIC08dFb+lx5L3ke9iz/fnmNofnsaVWg45ilOAW1w
LZtBwFu4S9wMwSp5mX+JJST/bVKAD5KgYxrQDNGQS9CKo7trQbR2GZ1RH/xLD84h
0g5xB6YiXr86t3+Tb6GNJzop+mrkoBMrMak+Q3WiGUNyO/s+4Z7Li50kiJ6p0erj
70g/it+SXpSpkAJ+8Aw+SykKpTh29CIvgL4hum4tqcJsswKKBOaX3SNbphUQyzfh
yC9cg5RZxQq+kb797gsFtfoaAQPzbtiJnWz2vsRHAMxthI+Kb84JvRyyCAprmmVB
Hh7FvGeR/cYZ65SVb/gUozPg0hm0aQY8g2HtON1SeLjZ6yvf9s2KE+L77gVLULxf
1vX1u0n7e2LH+2rJ+HKw2swMecGnDYsWYlTObHaNlnttgV/KufqRP18V3nQRaUPa
74WuHCm91UqjJmTptw9OKvLreI7FUXr7eEcV9dVUj0N1Fr9eVG0IB1VtaCBibIQI
KHe+giwCDH4ZY/6ymvfXiOwhBPfexePLxXj5sNc+g/qyG6xZxSlmyxJcMh8qjfiw
PeKzJQB8UKjKLBRP1BPTpdGLACauoflQj27a/BJrRSh/3rHDb8CyPy9CDZwIyM9Y
lIc+bW+I5n72UdBF2/0cM7xG3kCmrA36YDYh1F71xtBhOJtJGJ1eI5j4yi/Q6tW0
gaMJ+E3LpEd2IC4UkGvENIJjaOpAQCaDOuJhTtDCTScz7yIeIm1GOaBQ6kDqT6Gy
e7K2/KERLEsgGN0FnUUAxPoWQ0VVMGeNM2rAQAqjDhXrH1ASD9y5rVrDt2RcQjYT
+soiANCVzw6/1YjsoKO0rie/qi7f6VV2RMka4XPsZXHF9GgUFUt0DmgBRsrArQVM
6Ez36OHtVNMoIEwQejMXD5towot/IHZSkwoaNGRx9RptZtzPa22v4ekLu2rSR4Aq
EpigDSGOn5O8/NuatIIQWfjF+3M7ueDq7bj5Q7wdWkjmiFfq8pdxEK45vq/+r+Zg
jRzL0e1vqqBfPhZDRbBBvNNqD78UOU+qiPByuDJ1sK7SgQkTeF74ArOCnHDTXRcM
uY2+bP7GiAHlWFI/WPT9JXaEGiSIJwUJIBShHji8mNCyQk94p9en+41S8PHO26BT
80j1jx84yaYiSzXQd6cNy2L61/uB+FefmKEEN+LsHCNhAmS6gB/tbnk9gWK6YDEO
lL4/lcly/ZI2eXAGJoBP6ytD8bQp0J4b0MEHTsfoeOh1ePFfvwxVGudh2WrzJIrf
ZOGg0oxMKpDiyHTL8rdAr6ySds+DdgopRbPC+Z3pmkRf/sz+ihWTmTBANJcW9MoJ
/VhHNzfwPSNVCNjmNfT8jbXDC5Pihn2bgEyGSpVdkZYLlzxc/6PHlevAa7D9kU5p
iqkW2UvBRYCFp1G59TwI8S3I8rgo9CYJxocYxfNBOgo0qv8SEpfrkV3R2HOXi0qS
x3ozYE0rUmc58jpUW9KQi0s/Imu4s4D0glQdRD94EfAKxfa05sETwpLDOMB79G/I
LJNQAvYlZH2/x6Z4OwHuqQkQnI+RJdnU5CralOsQRs8xgb4hYYkKSr/WyPn1Fwv8
Za0hJ5bcDDdG/0Tg6JEnU346G13MQSraqhiTWDqJG1gLWyrz7UEzuiPypmE54jCP
G7pOoJSMD0Ui/xWBQHOPCqh19ohdLHw6OuBbvP4jcVQNjGdKh5estaK794cuUEi9
UFv268xtk2jHYpYJFXZkk9lPkBcsxoVj2ShpVQGiNxADJuwOteMBpEJ+gFeF+YOT
VNOpXpO33pD4VvJ0UPzVVpRmiRzBneBsOVYzkUJO/SHuIlwUzBAtF4xWhmesHGDn
tYBS/3s9cOUZGYI1TCcv5AGDyiQiHDL88YvuAuOV30V9DStQ3T10xDaPdmxKDwu/
U7oNhsDBJjgBmLq4odEoWWVNkmrRELivMH2LgzibrKEFbzPNOY/ljKPuhVIx0+Ug
G6TkKJKGuNgcbZSwfPM5Ze4fB95aZC9jUBrn5ipVlXb1K9OlGyLObghEnojZvI5n
JMhwmqT28JbJyvh0AlH/aFc414IMQtUqWPgfk4L0UftOzaa1DhR4sqYEXzl4MBzP
mt0Kd/3pWytPS6P6N15id/Rk46zHyQs6BApIgTpx4SBHQVY/jVDy8T/CiD2oIQuu
PvRZ1U5QBel3GzsCH6xA+KOFrw6dslrqWFxUM43+pIrzJdLq1KnuxzbeD5ad4enu
asi6RUtSAFxjm1MIrHkdi/Eb6Ebs/EpRYdiYYVzIpIIP8Q187xau2m9b8k5Fe9Eu
3MOQbduPGFJh3i273fYcCxuu/MEZC/VT2jWKszW7tUaPSwFPFlbb3wMs6/EqMi3p
OXyUsVHWejUipEavywa0nBowCJHnFaEdlFBCuuKED7wv+TTI+o2uDQYltTTvx6/5
x8BhKwWq91sK8goXA1rv8jrrzPo9TbJaLXsZ7xpfm8oE8Xt6hCz2nG65dfXh0OzK
rbR+AR4tNjY23hruFzAt+bZcdngc39Yb6bupaZ/ThrRkz0Cmjs6ePQyQE1hP2tep
shieVR4Fkcutk4ui26XKGpFw8/oe2RCilQdCB6o4kYeYZVs8Hn35Iu/8wv0MEfhA
lUdkPmUS9RYSMDHtMQgU5wI1YjHfOKTyiw9gMfGeLFbaPzNl9Be85OoUx5wXEhpv
2Iy2oyb7uSZIlWpYcTLh7HN8n2C5liz5cVKt362KDo9ALul+tCHfzN7erFcq0HaV
AmG1ejb8TtLZpXwofvOt4NR7yBVktVQb/R0VFFiG3fuicJpRGUHhNOsa8SW48f5O
6VtdP4/ppwXs+04eN2EOfee5RZkL4S9CJwan/2nZiCwFHwXxX25KhokuT1M58ZWz
YMpSAkmkCGPGEFsuuq8D2SSdthLeJIoiOn7OmFGn/4LOgjUeCb96dXW3Ugcg0kkn
ApRYxQ1IKuLkpHifQNliY5+RFrJvs433zfC6FORAHG2Jkpmi4wflZ5Wgh6Ntc2GQ
cKHDU44e0xTcqeilRSWx8viax5GaR12GNgMfAktxoot7XBPE4uuHQe+7lOhf+ffI
ZAaWaslUTsuOWu30iVbVUvmG0e7wwT0yZqyBLBjDC7R7mKXb5DvTHV/6nUTB7lUC
iVxtlqgnY/uu8XJKPCKoJq7AwCVqxMC2sh/gQNn+OxPaflzzC0r5xijmbXxM5nnj
/7ouTMumjLvXccZPurceJFH1nH7TpGl58o8xpCfoE7G0Os9K/LhMWsaPgJ7maWkN
XgRLRyC6YOOU/frnY73U8dVhOntkD6g/xZpsYIKsKcq85xQPhSH9BjYvUw17YTOM
v2tZFiFFH+Qgv37Q7Ik28ahCpi6ywbu/Q4h99i+ZHoN8g3pGeSsIpadJawj+BEAh
zzvWQIzzOL/GfTZ8gXmghG9Fvw7/czZHydNBOG56dmCnqBBQ+2RjalEhYVIuH/YP
gTtkBwujv8YDGBgsOM5kgQbPGzEmdc6Oz0N6DZL/bUJcUcTJ3qFi2DGBk0SVU7A5
g9XmSM2m1P3PyzbmGBhFCXac6TjniVHzaVJaPB5f33m/zJm6hlbaS6cmZsvP4PoL
ztpNZBRruppTTzzWR6Cnz7+R0hpkyIKvb2HmYr+HnMWMoRp3SlPDawTFmDxem7Ps
RgbvqLVoqgcnPSnOFyMFqv0gqjjHC+D4q9sBQKztxbQcJktO5iNPoyJFZOGB9k66
sm9JoHS2JEX5q/925l1FAnQl9XtSjJ5u/8M7QP1ZKYE2RwH3j7UhvqyDtzKUiFKW
sJiP2nrF2FglUUeH9+cMkzxjsR15lZFC9C9aLwH99aH7w7ffoDi8q4+3uiYOzd/3
oMxFUI77PyKP9X24QE5cApYfCaqphuGfYEVX+NXXj8Iopg4xfqEvoJvkwjgK0umK
IBv6uEFFOGQ7NPQMOs/t/jfwX7pu6tiMTneRYzGa9sQ9xljWRIF746/PgDuTSrW1
oSNFwRp4rAZOzE8ge5k801o1VIU3eDYXKqwUj9xoLQklw+hg0sFQyMdp8OkcZolW
lRTqmiiVH2BwzdQ0oLX60o0QJJVs5heRypx6oNmdnWv9i1nuDwI+7QbBGgBm4bNM
t2oUKs580sGVyjqx3jO4KG49q4IOFgd8KR9+pYZQWv+wUmqwaSCekScdnO0/mVMk
SndgkDUUNs+gB7EO3vw+40SH3y1vjYADnzILK8LyhaYKzfd/2erVBpBaTePrGpQj
fH16bITC37bIRDhDCSVlKlV8LP4HVKpvWj+UklQsl2gx466UGj8n/NzWueNo9YBZ
GiJgjWyBmUu6USZYCczyOMj0+OHx28sgYt2bBcWBf1Jt9Rvc0gIJxpOSxxyCq9M0
PZidd18ivPOJwrC+Qd7KcENf5W5Wd74ZzqayCJ0Q5lmr990S83Hk/2o6BdVPiFL+
xiIGmg0aRJfM5icUwKhbuWKn9nlj/UakQC9Qm8yNzkuiD5Aj91OOjNbd+nq3YVzt
s+sH5I25V4ze6THxpvEqejhIG014boNqLOsrmXpXaR+wiRSP00hI//+2EDx8TpJV
ThU37b/hweIgaAxcnJj8leSQbCH5cuC5Ww9QmP9wsEj9aOci6sicUVWkDr+mb1r9
8vMv/k8set10gBZrcylgDNYNyiJG0EDAraG3pX8GDEry4aUARZtcP1Dij6c9ZTLk
1DsKC79kbrc1Ldg+jfdYUOxO52IUxfsFr8jvnLcErXX5qxCjMAnk2chc9LdB7CnQ
abgnU09ws8fRrBtqrXjTPm0I7luLp1XzlWnba/dS/KclUQXgh/PN+xVeT2abo+5I
/YKGjggvVZ/HVpSWqiexa3PxAAmiprbXqbAEQj4IjRfmS9XoQ8tgghJhHtBay0e8
5KwXL9/wMWP6IaY7e2QFDwcNd4pnVEdqIxUfP7TyF3A/z0ST0LqKE2HjISWL/g5g
kcRV04+pnyr9VoKvBGtA8JO4srMWYw1w4GxP/90jdXS5glodgR4S++FfIIEtKE3s
`protect END_PROTECTED
