`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k+86NQfx1vhxhLo85ZiojcqDZuCTSahUJ4vVfZybdSi4tDFe9lU+Iut7xVo+HHlB
CttmPhgerHSvCRWGIBPIN1rr1tRAJljLmYcABMlyvSY8KmMpeCZzZ354QeUJnXph
bo+4e8itCwVYApo+B7qYpwOdUSU8Rq3Mq/AqLfb/vlo6IxVGGa1GaT/MbMsh9Zvn
oTRcysnxfg8wD9ODstzo8pg+JiK52cA2oG++XkCoFVfJmU/7gYL3ICKz8D5ucrfd
QV/QD/4fYqZQHIPryGCbSLg7/nX0UozHz2I14sO2VpB4K+PTzjOQhKzmtX6fp6EG
aZINmby4kKYl9r/2yyEAg0FFhZ49w9M9O56WEd5Avm3MOWrPE46jnV/xk3Q5qQUR
/QL0MSDS8wj+dRqbGnv/fpI8Yi4Hl5WoWrvmIRGG1sMXn2s4y4ZTasJb+ZC5spXz
4FnBuhfIM7xd6Or0h8McPRJOXvXGtFfz2tj2u8PUWcq8pQmwLQpaTo0DktH96ni3
lued4P8/iQCYPkBCWL2xM9BfRmxxCRpLxK1zGjM3CFqk/5bxMYy25CVQKxCDsQkK
3ud788y+CBgJAdfNfTCqan7m4rnDJOLexIktbbDTqwhgzJTQamJBYRXr8lE3q5s3
8iGpBIGQLvE4MYoPEHBZX1WHzZazE1mT2lCrPhNz4bF6lgvE67gyfXriX86mI9dn
QLHiGwqL9BXtP8mRuCYCJtgWR3MsFKAqxRd5Pb1dnweCdRzCnkxKPo2L+VeKhgZZ
R9kCL8MpHzCkNaN2UC8UgYuWVnw2/CV36yJJGoDvLm3dgauJwzEjMJKr/x4Acaqd
lMecuzAaBoKmUxYUWn1ndIqqVbHNrqLCVoyQN5AxeokEHiSVkRcma8W6LGd7TMm0
pRmilqUV567/QUFDvjxDJn5tTsYRwvuKZ2WUi8mdNiWR+I87jgc8AxnYq1iErAVX
X4DjwfPkxeUalPdJP0GfSOPb+FWNEzyjMVOdnu2wBew=
`protect END_PROTECTED
