`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ABsfbFXmnCI5o+cv1xE53tlKeQpqea2UAAgZZJRUiSKtkIOd/7v06mXyOwPOJBdo
wXWZw4PkasworZmPrRmc1ubuimE0JE0tM5GuMlNx29N1uz7J8Nq0KQx4ijwfBeJO
GXUfiociowRlPXnGNYhQWQyHfWCEoaddOPc6Oktu+RgSMdWvdUSF/pjxc5D98Cy2
SlQxdgbncCItYCw483iF31RBgQOg+R9bVNFR3i7VdGqiIJ9twW9JcdgidOIOUrH4
c/PBR4u0E+U3W22MJmZx6eismbKpzzrpFZuYGhvxZtrMTLBtRYAjaBQb2NuWy88X
GgDJsWtgDhiOsbuhYlX8KQpI0GTXjYF16RhYVnNaJstXzF0FrfsDLeODFOP2+TYz
LdmHbB3QDBEAXo6xvLk86HrdtdoUdJ0YZZH9UbP+HZeWhjVW53/hxCdTYAcuOSLf
K44eg3FtZYZbwHONiuAAKRa0r1iB2qYCNfX0GJqJU/cXFaNz1bLkXjl10BfCpIL6
mOTWD0DDmyva/QO/Hbse9lLyqjQ3/5znABWQha7BcqBYOFhD5Z9cMZlrJMDgLOEi
wAfZ/goA1iGHXZWp/Imhzq4lADFCYARmyixieTNmbMum2BuRmxnHdnhNEALL8BtL
99R+gafwLr8g7wVWc6OLBDhRod4vmHEeVePQ+fwxnWYZdP4RwIQ4jpGB9BciaahM
XKq1rng+b2SyOqNSknSBPYJ82pIZ26jBwwQEuoc6/IKXk+j4FvVlt5OK2+6VFsbj
j1JqQhAh4JJOlxeRXX1416yZWoDg0K1zqY7mM2sLivldcZxWuot/TG+4WxGFDQVw
YNn6J7GlHkiazAqk6c3Rb1QBHOgy8GI6M32RWqgeruSWlmQzIzYFv/h3lcnd5O6k
9+9LcAbJ1d2uB1lmu1mdSs9yt6lDMN0In4yT9dUP8BX8wo5UuNGBVVgBlKIENonI
hBBrhR7euqb3YaqvwhH6l/TMfbBeg+xucppB25wFdcF2ECCPgJG1toQ7g23LcfYA
eoO925bsOLP70qS/u7qg3J1FC6sTY3CN2pwM/9x9rBAGvKRN/fVwv16lblRt2Apx
9sqlI98iJw8uYTUKDW0ZFD3z4Kn1qF7iNMoPNOmnWXkJ05Weg5GLo/BkjwTi/3ys
27Y8a6eLO5xgvv5z66LXrogxWMFt6VnOKTqL6LamgqMGnTKbqxHDcaHokMD/FLYh
nsXknvIzq2ojnn6c/hav6Bj4KmUSVRdLCC6S9nVPd9m712XbKhQHUTzjyKnu+235
Fzb3lthJICfwO7dMaSX9v6uw88IRyPPS+r+h27nECg3mNg1QFGR2KKyJO7XB6Hrp
Z4zHAx9NyAqxSL7DLuGFUun9Nyqe2v2jVWjdjw9SOJMxoT34Se3ZNNTLmfzOoZMf
zS9WPcEWYKM+LwOU7ErR/8LrfsAQAhZp0zQ691CQ0QGDSNV603Q7Gko3VfTI3VCd
5m7mV72d3xetQdRwUBUwfwkULLrOSXNClT3LP6O6Cqf+m5JNVAUFyiWOtaM44o0l
LQIaPCe/xweAmYSMYJfMxHU/9rKh7LmS9Q9q6tCue/dUJYIcQVwrFR/aqFcpE9mp
C5Air1Iohlo1IEAq+ZJF8bdi0aRjaLsg5XIG/oIziXvdVRf/eSIRQWI66bKbpMHD
O6jtvDhDy0Mjq9jLZBMgSVvwvb5Ur/9wW+zJ3A9jol0=
`protect END_PROTECTED
