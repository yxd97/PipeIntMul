`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M9joAHmGqlEkeXHj26EY9MAFgCkEDY3prlYOF5EAq1N9Yto9KLWl6TbSLG5dbJ5Y
lmOBLS8mYTkX43To6TU0n5bcoVJNG5PU7NkTwMTvjgMaSn9vO6PNw++DesHkOL15
9/tCmOgZQrZdORNBzDjPUpowq/4cqeP/jDEIC6GneCiCrHvHYQnTQIW/s/CuYAdD
80sdt+5CGqAusIj994w+RijZlxrhKnkGsMAnM7SVPZP474eXv4uXm85TG2W6Et94
/aIHHTrQX91i0iZ9slNtuW6LqB7LP9VIHMCYYOl5kQNAmnFvmR1gkvnTce3ikvpG
TNFyRf7rh+L7+lMS7LxcLAv3mUzPhZMvcD4a4CShffvlqvus2v23lKBYPguWXfw/
/PvTPTI4vmUA5hGfBA4ILcXr2mmykoAxSbFN30Mbi2Dy+Gav1lUyBQ+eMP7q2yUU
I4KZNRsNZ67TUJ8HElF3c/CNmvKktHivB+V12pfc0FqMtopM6jao94YBzIcn6P5H
7OqwukJEGqrA3iwjhLU4c6MmsaL0xVkbdmeKYH4xNSTB/udM+b6rkxUj2f/e0Rx6
nQcEjik2LLhUSPHQemoEadPqzfbKZ2whwGAFqAKYtFIyvUGY5lwQxxRO5Fb9gd1z
ZVmEDrwYtY3pylGcENbICOh0ZbjBUcKSCeNyMXxd4zbA9fEAZiGAoLiLrAF42HUp
gwxzo+U/u8HG4pDB7F1+uIVxhrWO9oaZ2VbQJLnDZfIUW3bKy2+xZOMxddEc/1Yr
lL1EkUXB9BP5iriWltuZijYI8UBAPUT+kL3TrKblZ65vkSElnPeHDdv659LavoPz
O8okKF70KwXYrBilA/z1FG1wzuVu03HWTJcUvik5WQPihiK6KdVnW8JmsbeH5h5r
1RXkBIGREeA2oCcIx9d6zSpKaJ/ogBsSbI2fCHHc9LoftCOEr1mBb/Yn1f+1Xu67
SkG1ysZPsLkq9ZaqLCqYiSTVnk2KffD9x4r/tsdids0F2gbZ/uEvncoMdy9E6KZE
i41sRd0SIR++cTsQ4m6HOZqL2Yc18nyOYhC36AOJkn6coR3dG6/Z6xrmZXMoWDTj
OsqlcT348KX2dmMVru7Toy02cvlaBgd6lcLjJsiNSAg=
`protect END_PROTECTED
