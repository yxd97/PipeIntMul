`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H9mSFL1pykpjfQJmXLGnrKz/FoNLoOxzwqC45KkADAaT1Dabxa0g8Y6pkukjbVzu
xdude7wYREgNCnAhEmSXxUu3Q2evbXwPZVDS4xFDWesg3TtZfF5eb2R3TXAIN24c
tceoU/lVWAnIsmW7hywKq36i8KrjopCw7sscw8hXWYYbKXuBpsYJ2QbFTa6WGOz7
xWLJGDvaVhfgtvuEL1fHl8QmBxqsyfZ3RzgpUH/UEEPbaI+vCcBok6aRBkf5rstP
yFD5PGVVj3AsG6UvfOmu6y5Q1Js3eCJBVa9HumFKW1nMkArGf9Lxo5queIPKWPRP
s3tfRYjO7k3fV0Zx/neYC6/fFvODdZIvberDIqgEauSWVq39VaYhL8A9OpQbMB+y
ikrCn66PHv2IO3oT+hJJy2rz+iGMadBzzRgWRaho0Ems7Wrm1CN15RDRlA1cI4Fb
bGjpUWYCt3YOHjUOeaRg6XpkBz/OU0pfPpLlB14mph6tjlyo2IgWm8zHAKGBIhz7
aDs8dl4dyPZBEDNWHmyQtfuYZwlF33XZPz0nrjcoPRFK3VW5dHzrXAa33K59QLQG
cPGaFe2y/+mt5HUY17zgBsGo2Opq9PMuebrxkbI2JXf4EpwtdEVdy+RrVFHGaBeN
d7NTvRSJ/1AiOUXw2bqRbdBAiSR8VrNy3JHe7jjiW7R8YLLLhhwl359+n3N5o8K4
o5wABnJ9PUD8eJTad7j+rovl2U2gW2pJozRkWCSfxWorHPujEiR1g8o2CBPMKgEA
zLC9ILpXuztZzLdWqMGMfJaQ028FOYwt04i5xsIl4/8KjZqdGfdpn9hSSd+KmxLw
9HQAE1+LXHJKWsPOVQq12nFqw9Jj0hxzX6b6qCWzQYu+bgAzehZgAWSagH8pAM5r
KYiSMKBhYowJyqF8YKd4fDQ/r62iUgLjA4PGhwjTZZuKrlnlTaYrgozYFc2I9ESL
PlGE5vP+V2O6/0/9JwdUac3RVPslDohHvYka0wltJ57z43W01ba9b08BGiQA95UU
wL1ZBK6zkbanLsDiYxl8IHvwZAVYQdvQ3TUZmMH53JsozEZos3CqLBh0NTaHXs3l
flmmLjhiul/lozOFNgIwVtIUKPBH6ZCfjklJ1vM6CHKXTVQkgZjeunGvwRrK4tS9
5Ax9jAI7LgnGQRFmydTlYjfJ42GJEf4c11lgHA/NpzOqlkEbYZiMgadQSLHR4HF8
`protect END_PROTECTED
