`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OZowXpW62a1/bns4iZCnJ9ACkn1eo2fg7HMR+W++zY+thpVE0tHOoaQUgnFyPPs7
xsw/t969/NZxeSjgtgr60Fy1qqB+/+CiAyvlsa2XR51J1QuLuZQDxVG4+ggA0q/7
m4sj5CTM4Wf1La/Mg21aYcS4DXkZGguIovqHhFl8YvGsq+dru1bIRQhpzug5K1fH
SZN0gab8+aXCrGlKB+I8Bwu3Z/7GELK41YBv3S/vfq20QCAvH0ZDIksz9u4e+wY6
za+BO7h/koOYfT0oOTo6EccKkPiaGwIP5j7JZBBul/FJ9nVvoI4xI9TihdCCgpWK
FEeyibAO58k35iQ0M6TZXHi7kuk9zKu6F0EHrvKlYhv92XK0vsKINILj+PhvlakP
4ohmS00yr42/rhzfvqPDhGVydQIM7TwQdDel9QjquteYVVfe//y71rKRi/mzAKF9
CKSuMYPL92j6hmK9txTzxeI5iDLy3f3OWobjv8NZFDRnpa0UoRVyVxflHsC6018J
B0aSBmN8yT5CUYj6XAY9GtAHVOFJGk2FananYanbmwGJo9PwjASTCsvHEv6Hu8gc
UH0b8TsM3G5gEwYMvNUG0fvE1AAHl4Is2CrvVaidsivJivXEHQ77wyttN2I4MiJ0
Zo8CASmzoh3yJ6C/Mi9NK8MQhaU9IsBwbSusYV6riM/JZbiB4AjTHqff2PXbbw1x
4n7/rjzCkNWMgI9tNM4TVgrNBZxVNTlV2W0+YQRKEWeREOwYxdcXdwmym2zTddG1
suT+eRSGJIzFa2e9CF0+W4jyU0FJFGWCdhBQuO/suvX+q9wao6yb7X8YSnAc/dD0
8PhT/Fbvr8sQ3P2LmnLk2zThQPo94STvfoWOws+LZkXzJcDXT9+4sxHHazNS4SX0
G4FEcwi+BnvXghVx1ToM5INQeGcFLW8ehSqM+7W+We+gkQFHQtg82Rw0NIVhJ8wm
yKyj1cJQ71eEelBVbaZujLvliMbXzUBT1ehSVRt1RF1O3JRZFav2qooR9k8SX0aK
VBiiqHTWw/zOCyev/7m3OTb1ks/9F30fzbRlOh4g+PekBagPC7MMZDiJVlCO4yhF
Pqw7rh6PSMyuHJzHW7AdNlVPlPMF5fNQKkdBbZuEUoBhHQX20QMtcBag8F9u2dlp
Xab+BavCYX4Z343X204m+jLyBb9zyfCoEfTH0/YRp7lqRf8eUr+r0ShcrL96L4ho
/0wEg66igwxPkuCrlLgAtwITIYccErn5n7qVCingGZ48UVWcjdzZV7KP12wYJ3WI
R0aHGUVxtdHIimON3nXfL6+OOHeBo7bZ53Fe4mjbeKyE+p3b/MIT/MNUr+IM90Mm
i4R5Pn/4X68fQlLIjHcUISEY94Y13SC1Dk8d2B+cUbBsXTrcYOiYoBaLoTXJ29b8
rVDwEXjWiGNOBhjSHYlmurng9Fob37hHfXsBi0jnuIuik7fGY2IdZ6UKK8wcN9hb
yE2nqiIVduVJrfwO0XCewucuHqruXaWzuKe1yc/55zt3xFPbPA3VhlxrLpLonbqL
SbfbU97kbZbtY11brzCEN6e9ZIoBMsjE1u3ueQQ864deWzeCnfHPHBVqpI/pFFmJ
2sMou0rWwnNQ6bRjYtJUMLYLlWVRkGJ/IiKtv3lY8XZaYmJHLEhWP+IWOAne2GVs
skdeIeiKrFozM1xgNHiVZdE/iSSjDitjKH6X84rqE76+AqgIubwHQ36zMlWTc2NR
Hxh+k81NPTLOB1HxXlDZJZSnO9GJWt1hVEu5eeURGr89OAnnJ+yBs1i6b3fmejcd
DL1w+WavjMu1Ol8r3S2pBDEEeBoFBvNhdUKc+bHVf0eqAnTUtKvAJZEx1e/3uGLl
unBM18mvuKiEtdi8wYJlqLsDWk5PpquULWeOrq+t+t+vTryH6XO4knvPbMC8+bXm
0YF5IkyySN4LQLovl9oZN+/bN0IfmdSrc3EL9mb5INcCEJ6L74c/cQIZKwboS7E9
TXW97u30fEm8mSQK7YNW3XpSdrNHd8n2DXnMCb2lFzNrNQEOwM1ahZpxVVK2LeoP
FN6jvop172BegR+Biy7YMczV9qvhqezMWSxVnWNuEps=
`protect END_PROTECTED
