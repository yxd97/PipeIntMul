`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Cw2VN781UXMfl+Mozl2drDOVhVgjzVphvpyjY9Ay9BfLyXNYHd1LY6fZNvpG325R
OvHdwe1vHev66UmvIU4zJMusKihJeMlANZuHynS9EUCistGg/ftT7GgOxwTFPcDo
sFBfeRnls5bw4dNiXAKNS9Febs6k7XcKutcQgxNDW1iRZGPW5WPhM7p+6/0RDI/F
VAEEGrDDIqzLJ056tcPPjT1cxQbEC2kYQtrzwFkHIW/bStdYNejpkGpXFUUOSpmp
XQaQ9BUm/YoA6I3tKb5vYvWBVkHsZBfn2jHFk+t9L+zi33fKmAZTl9JMqf0INzJA
zOT9G7KiNvYlGfxrU+kmC87PLhOPtYFe72RlnSXWY/drShndfAAqxuppIuR3cC/6
VE/zQ/EYsk5q7PQURmaHQcZn3+rqrzkqT/uQS9HI+cA=
`protect END_PROTECTED
