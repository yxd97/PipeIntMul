`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GlKIxZ5VpLsegnFkPq2rwB9ymDLwQvmoyL3psxPs6+pXWwZWnKjouFpeTCpQKQgr
MaiWsvYyR3vKnQlVvgax4g3cPdfkWUm4GJvyINICKoXCeYfznH5YMeZPOPt/9/9A
rC4RKke4EkflvaVF+zJeknoRIBb0hCZOEkhYo8kS1//y/+JkSUfiww0LZvWrmH6K
KiuclmwAufLA3+k5dB/SjSdSN3ocnB9I6QBEjY2EbFk0deS5PkyDVZCtKBoT1foY
VlwtcxhTDIaBpTTODpTuwqqZOFHdB6eY+zKImjhhEF7FZdsPF5ua1CoJpYDB2B7z
A+HOlKkZ99Hv6Pq0sI9hrrb6kRK3NVrtS5TKo+z5VJSIIl7lhPgZwE5HZRII3byx
h77XTVum4y7UrkxqUT4uWjx4WzR3mONbObsOjDoMVm+VuiikZTh4gblkF+5+MWtP
Yk9RDpo1mZHjQY5AWHq/HcBQUvyH0taVaqUR4q9DcqgeANMSKpwWcbfQ2a04xanT
UtaUq5gnNaaY2SJx+YH8Dj3HygE/pWvfy8naFv4a9FFJn+fzw+/e6z2S4oKeG5Wk
0YTTdIXSCbsnHTQv9kSwxHw5W76s9kyei12c1lTQe/COyYCkGAzNw7b39m/JNkWO
nHrkcShdrsMbj/zs7ofbajkp+QvBydmHGEeV3MdPVHOnksGuWnfK0Jq7M803ZjBG
cMWTXiccWq15Li9H8eXUVX+og2TKb/wOjfYMjJ3Y0puEGEm9XoPKyIkStRayX3Fh
piKhVZf1ZG2Z/xGwUXxmn5raLOb7Ncn1T7DppCBcCKJdkJf0N+3ptctxgGHTUbSr
+fL5LMWnQCzG+i3iOYdNp0sCFJEp9Rcm+f/k70S/A+ArPo6cu8cW23pMh/+qcEob
DX98hYfqnecXeR+/E85I0jaiMzIBMKJ5kUUm7st8Zr8QhQcZCp9vATo/Z7/ezPAm
CnPtGdLCR3+zbfgb9KO3GGWsZYKZdZEiPhiTkIEB08VEdLJRy88jUmihdCA6j5iZ
R0ExR6qZJ6Sxu7CxknZvX8SbFBnZ+s2BW6A7tFeReQhFfI2f8PPZU/o0w+0d54d0
QBL50pJqiWJaWdhr8Jrp5Z2X8Ly2hxmlBWNkyDv0H/1ODt4i6B7keEVEwntDoWre
UBZtqqPEXm2D09Xa36AK7zdaE6TWOHbczRV089jHChdZ5zAAX4DEZvsIn35riD3v
uZY4LCL4ptiHWj8FL+agUZsIpOWC++dUnEpVyfS9sNMOQMGuOf65g15F08qjA2uY
RmWYoU19lyEF50d4GBrShqaNVA3f70e7oqd0KOszJUr7xvclEUeCxP7qoljBi6gF
i4YxnjE1Y/w4zzpOpHiPtJp9QESoLzHphizFpsKsRE0YIMsQ+X2tfYz+UXBJCPAv
Xi0WF1WozSXJiQyAHLVWA2gsmYEK+iou6clCNGOw3PlRXSS47us4dgKjbebFsMpE
2ksFSr7aeACMiM4gYIj7qGR6dmSwD/GtXzToh1wAVks8zU26Qx3YVd4ouUEPTBpc
JjzRvdE+Hd+thrVzaUFkrVAIWzN8t7snp73hRERBKkfeTaN8PD+zg9p22sWyHJR5
2zjVza7Am9Rv/ZMU4WaZ7vLx56MwuY37pHqfUxBY4BqxRjqsFxBPtd7ToJ/TrC6t
v88LbJbVkEQuBGAPhI4dqfjLq2hk/n2QKWTj2FhhQmhN8gPTX47BQ8JRnp/+IITE
DBGotujdOkVyCxI/JQXqvd5/yDUVkNVf4ag604kAla/UFK0i+3DByaB0GjX6d9ih
duWiWDfpPcRDBnEKPiJgPPHxuOr76A/+V3/JHQ0irdFX/7XXNpbJ+Ni2AaMTV10f
xGBKVLTSzTmhoX+Od0A4KVOavAlsVQcLPsZbZe6DWHs8lS4hEJOB8qu7oi6cX14i
Y5Mm44SlaNTXAbt+bd9sDp7TORECPpgaWYm4Qr2Cb0ZydJy/0rdAu1g3obaGHTfD
ceQvo0eVKA95lMpONaRYOQ6BRC4SgP/66KwzXbK1vMmKMBJJO4rm2QWNi3FR8+fJ
LvJiSxASkNPJweYhI+fvSJ+mmhWZqSp/km5iR/2w9oIfnN11bpGli9VN7T+UdEwx
OfW6JfVdOO0LkptY589GJP6DC6F9AkcXUyW80Z8TRXEhvLwUmeNQddjEMUwwLUsy
au3nT6MdtpDXGTn9YBhJ6GqMdns8wM/m3PXUiDsJwpwD0ur7h63f+TzH+GG2DHp3
5rPmmsdDX7fVgaST+AXVJ+QbMYBAyfHCiygNAyGtJafuT3WwA2sm/5HcpgShPWgN
`protect END_PROTECTED
