`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKC0h1z28+VDLpDKPQRE2V3Bz+npYWSOIqbWrmc9NM66x8hwu/eFrjPWhMNm+S1c
Wxqo4i5fCJSVxFOBiYBS2S1Hkr5CII7UI9UMp/ZoNcGNzjn1Ws1Fo7n0RwkYD2Iq
bJKyBy/pY5tJIMv9nz8MOLbJU6EVUlKGvR79BfVWnk6Neiqv+NbCmOlIDZSRh936
+aHA7kQg2ttqJTsfY/isvHw9Pr2pHzkJDRvbZHwEnpXuHryK7iQ+NIyJYmOF8zTE
/k4aTv7ecqC8JfG2c0M41M04EnvwmkWdNclMrx5UoroLCLIDdRZsjKwaQeKUJb2Y
rd1rjHqFxizG//XiAF+n7ukmnOwFrAyuPtskIC2zf6aniJh2iBSzLf73DNwlS43+
vpZU3plDcJ9sAkEPQLMzkcj99BrOlY+Z3ZjSduezh87GwcVC79Ypj9pCfItCr6to
82dPj5QdhB0sAlHTYDhXy38MC9dXgSWocr6XqC2peSZ4LA3oEBjK1QK0AvLNH709
2FRUWP9s1uktFrpewaaCIiqTNvO02oYF8jG8NLsZa7ED8h63i9lOijkFQIGgBBwM
m1hWlZTt6wtJwd5Gx9YwCpJ5m9llLN8O/OFhSJ4eIc9SRtofW5vjCo64liKJ6qXk
bMeoAHHebBd7JwLz5Cfd0peY+pay7sFc2/3aTv6SWLXUSnQ+Ye2Ggq/QfS8vMy/6
YvAgfHeLeAUx3FqhCVDRoHLHK3F0zP13fAQ2+noj8EXEUDj31Txkf4xzk9UTkmLZ
6dSDnqaRwJ0kSZo0JOTuUA==
`protect END_PROTECTED
