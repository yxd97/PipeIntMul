`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuNhu0DOYxOjsS0P6Yprt/d30GI63H1YRGJwJMEJ5wqb9pqlf2lrj0aNnaz+xhCs
6d0n4sMpAwUHBPaaGfLEppMNHAQvPu3oJhOLh308nGTfoh/EnBCYj4X1iEBSb0Ml
No5+giLZ9cGhSesSJkyeJnHw4PzFT06ZP3VBgBjIfj8WBjsP7MqMxwlhv8Nc3+TK
BPqEsAIzaUzfrZM+jmflkPt5pqyZuzltF0KnQjmBespv6kBvxA3IB5GFOB3BeE9H
WRH2qp5Ev6RBtDQBhgyo94HSeyEmGGq9XBHkHr0LNHF+uM/xomzNg2fHpWTGeZ4T
T3ocJ9FOWC4KVHQJZ9WDnFbyLhCjxrfx3m9DqUTAOHoCj7HJDR/Tiz1q0Ut74lM3
fgJ8zlheqnfdFHRu2uVTKFnsH8gGIdciqzITvg5mgYE=
`protect END_PROTECTED
