`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+PrDaMyRgatJxqERTbGWLyciupWvRVfgAwAViX/x1cE1wibA6K7GJPOH3ZI87pz
BjTmaT/LgAqaF0eJqPgaLwJqdqWzrs8X7UrsZbWVGcEAJfum/P0+ipYhZU1u7PVx
7AOjs8KQ0cRlaMb3Kl4/E2L7owrtiuPgI9DqDoyxQTg6B1yPe4okRzE4heG/3/nI
g7iLFHteHaTASg9DnCsCRodkSIOo8MEDq6rqbXNRDjMcyRiWHSFS7+ZoQ+6EH/uf
WEJ3YJhmFDUdJKmWzuxPwkPGHrhsIqQEhQFfHkLmPOsaErlJfr3GAfVt4VqdYJmO
KIMyvTRQICmXuOcYqE2UnKOtovXgxNM0Y7n1mxqj8Zv5MQUTldPsaaCHlC8CFQ/3
3VGdIXHv6wV2UMtLEyrhOQ==
`protect END_PROTECTED
