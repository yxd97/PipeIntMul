`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6gOkTowDmBqq4GofJyfKLdh/qa7p2aB+LIGF7XO5GVg1nIMJ0pXDI8X8DgNSyrx
5+y8DuarBJ7PoO9KzZuP2C0flmIdp45nUMTfkjSZxWwPF4ge2JbfWdy3BkGih02Q
dUJA1XSuTbokKzAFBwOfMrgVbyc+wdE06wUAneDS5ZrKkWJ7HvIJ1XmMAxoXsLKJ
2gRT+1ZbPagyVIhFyLi1E5TbJbEmaEZSlqD4trEHtUqKhl1jW5v3wznUY9vj8vTM
+BbtcKFSb7jhcwdrn7Cm5Nu6YQEJsw5MV7+AAbH61MoE/fFQZMlVz8oH7p1LRyL5
+ykIzHrRNzieqzPInNb97/1tAsPaod6i1aCOlZ/EZhea7p2Bht310N8qzrPm+4/0
q+bG/JOGPrugkgEApXuW+UURWsAzIq7/q8wg4I/ygZM7yLhTlh+UzN2X+i6/lflE
VE76RmOpI1kt4Lfhd3F2lZtYSjd5toCX/L/3dr/BbMR04ZxUK0jyjO2Beq3Rl1PN
Kas29yFFz0Zg6faU5efsLx0KdjvohP+4MA5fEAY8XGJ+fgSaBzFv5o1/QdWJKLnY
T2ag956koPRKGTl3kjOZ9tNI9njLxumuFbUmG1jYOqYBDP8yz+teKSoz10i7FJnM
DsO8VPdr3xo2TDSdQjzMV4/VHAptcxagY5HlMXJB9Gcs3IgJqrrnCoeHDltfJ4pc
TC2PZNzNGq5E6TPv9HLfVwQJu/4OUn4bkGak4GTTvuci4KAw1XX+B/LcXp4KJI26
q9yJXF7xYiJw7Z2Blbin3FYf9HUFI0AFBQXI9+SE9PBdpQbMO/6Ce5EoMEIjSa3e
qCr02F69w1f1v8idkgs0idAjXR5jG4E0lIAz4unQ2VinhrNZZWRF4SkfeP0y+Eay
SEAkbY4pSXAwYBGQkNBkrzzbqJe1vuS/KrBw/JHdjQLEecj6qHcJpVVndtiQbLCT
KuuZT+GIwsBt1ZsPwEyfHnpq+7oMDxJMMipNguNdI36dPigoa5jQHe/QPPnzWfE9
1izcw6g6DQpXd5uS68/AfnymAZz1EPjY0w0K6Mf6wYt7iBGI90bKkTgdI0JrCfs3
bsnacjXNv95yxTWSPUgQfaIjCKB/DlRzYQlJKY6PzCMBMCiGDyLIOYi7RETzIavd
WLuPPQOaVleuk3ARipOHv4Q0F0XqspIE7yWTiRAJ12f2EqCKMNOPODYAhx/r0AST
ogz1G5SdS7MyevfWvW22etUWiiFLFyp319KnlE+T2WU6xftVdK8gagLQrRse+Xol
`protect END_PROTECTED
