`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q1CjekLWo7zhqhnxdRYRI5m3FlxX3tPlg28H8LMCo2JuT+cwB6aNEp34yCbrzloN
CwYhthDYdb2+oPHCvcu+qVKqnIrUVPA7XWfAq3fSw/5ROn3UbUNKI02+7fknZTkP
/C7BLgGcDGgkt7JFjrMViZabJKXQ3U3y3dAcDXnO2gCksZc2IWm0mdhAql8ci3bK
WRA4ZfTAR/1DTEJlGL7V4aPh3UqKwv4i7crzdIzEejVS6QWB7pV9eaXya/GlFpRG
37Yu2H0yhoqWARzfeL+zFPoHUBhaFpSza6g2HlOZfX0AXUURXPCZHSygv22yumJa
DRzxkrAIEA8G74ZjgUylcjglVFY9lbnare1MtE1bFUrZENdJYjPfaRmRJhnaBb3X
Douybm75xn2LzMjZ825jwK3ygVsAfReq/JmXxsStfh02VVgLKp/jtv1jXLFtiAR0
UgitfHdHjOXpmhdnD7p2qcgfk0zIeBQ01XRy0ha2z4gOApjOY3za5WJWt2r3ISnG
e4bY7h7Vxj0LPFo4lxrKYZtTP5dOwGfMr5v9cDIoGCKy9qGiNlOMuQf77YhcOrfK
yrJ1CW4gigxb09NYFtcJ3VpY5eVSLXeSsW92Je23GzIEU/QA2fv/mY9MGMRLI+7S
VR3+FKxEd1ppzexMiX8nW9R4Z0Y9Y6SQ8uyozCqP6D3VqfOLp8j0mC+U0V1Vz5pM
W1Y5h+XcdjROHOcCXIJlD69p+f/JbkDc+Cd/82zhp6TFrJe+fcikzkWJ2pgiqxke
RhKTkH82mAslEv2B/v0m2COcf8REee0puUkTJOQ4GAjRoSanJgfClL0ctdxxg4QV
x2r62FBxkFj/ihLAeTsNJELFMOTg5IO3VRBQImSuRgON2fJ9C6suAxl3jaxxOdaN
A2IoBGbv3T1eqKoQhq5Kg3/Yk+0i2zhAAT3g1jMUeTwH42iQknkZcMk3YnLa/+FC
qEbVOGIcSXKdW6mfg0V5J3Dh4yodK6PQr9IaClBZJf1Ol0crncjGdxFe/0VJK3PD
TIFoLlyOz1OqYFXVeTUlrK1K3epLnguBVz5+ItzSKA4yI67B+NwdWRMkjV+OkuYu
+F3Pd9J/YHIVTHtqcMCFWnF/sMmnhoHgj60GLDBGruItpyVEcfoa+116rKOh/6eg
MZItYakOk9JO/ZKcnN6rV0bEVnjwwNT7/gEuEJMKjb5o4i/3gtYqn39gIeCRf2sf
Xsz16qZKUAZJerXxD696Yl7mVHDJuy5l2DF38SBhSHRL9RyurQrMh6nqRC3vdINx
QTR1I052jy8wc2Lxj7qCBV2QbwlbfJZbOM9ofnTZxCg472Bj2yaV6zFMppm4a+Yk
8US4YAnf6We2tn0Ttb4Xm3mgtVbnAdiK2xE0Ic5mR1fHW6vCB6cJpS6Nd3rVKscM
b9Rz384jByRnhdhZ2+uecWuw5A5DC+0fRTx0OugUjmcadRRmHxWdczFOOQhoMvMo
0uRgE6uI7vuG+kKtUzIu3I42FJ/XORpUYtbj8UQbBhrTIcOJYRwfShhVVqTxT/nL
5f8I+JdPeLFSDFpqQP9aeQS3R0xueHrh2pifKBq8BqZsfZKiCZOknxnoMKdaqwOv
XvoQIDlAewty1j/9BAHYPqPwrG8Zh5zTGSH+7r/zLa/x03GTGLwixq26YpPnIC+1
8Eobk/AmTYzzBoFCDg1WHT/zg/Rv2lw4SDr02gsznEBft6jEn7eLAsLsZsSQ77B+
Zs10Ll12cty7/OdFXR90m3wI1efNTDvfGpXyfIXbdATkMproS4zCdBNGCixDAe1X
DKvJr64iPiEud4/oWg5+S3NWdH3a0WlnHmlLr26UNmqWwtkpiEvWN5xakChtTCQ3
xGbYHtkNI940W00h42R4Ph34RI/k66Wbj5lwBZxtCVKY0IY3ozErpFvHeH32Z9rR
9Q51/Q++uxuCOHOp8fwr+m+sD+RdTiyeOBczTLVGjJsqvO/yxdXbSK2pdHYwcsYt
4kYErIo35XJvmUt4Ze5lyRt0CGtZgOTS06OP7okZfcE1l7ZAu0mKrl+lkZ/KuRD4
mot9CL+58raNtTYwKOaF65G+igGwVq/lGw76tORQi9QmVctutwJwG1G5TVKA7qMQ
GxosLzyjK7x8wfiM1xK6/lKIdk18QU3rC39bYR8OgrCAq1LJolRS7+plx6u80wkX
sTCiOf+4f0mo2o6+T9Gt9dVle0FP95c9lUOtrUrmo5fJBmEQUgd2lixNkFZHGWSX
vstuJxO7qSDWmR+Xba+/Tc72bEQFUQI6tKZjEZ5AX6C0M+s5pw13KWngvi7UOfi8
eh/rqMcsfgS9O1gArzI+Zg==
`protect END_PROTECTED
