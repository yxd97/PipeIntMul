`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgmyXcPoatJ4AGXD7hm096lASD61QTEX+eP9fDzSxrt7zkxhQlPDZJ3oqpM+OpqV
n47O24NaiXC1jKWgXOAUE0ssaZaWWwVsEwjRl1hmRI3aqAIPHfEfH3kqlI3AsIBe
/BddCoE3et05RuzQ0jp6v09gRSguSiOylk3Ebrvh30rFB5NMmQYUViMNVD+0LYgK
IoWWv2eBB4JRa8Rp6ttwRKeJd/IDPALl6TTJDuy7lx0jcE+c1JuESJ8OdnP5n4X+
6qzKdWxdsvXzTFKEeNIjxb1IwgU7C34pdXrGiAfdnIjDmFGz1Mp/yVY/VL9bZcef
JEA9y1njhQzd/kUxSqV6pVgTeX2ICRRi1Z8mDXSPpORAE/Dkvlya1vKfkEEYBbgF
PmLtRKPmphzUSETvQ3DVCJv6hgKilSF+wVUJLmW0am2NpIqUq0hmnzn1M1ZtdZ81
//5gAf3tjbVSJ7yS3jigbha1n+3MhEZs5Q5lgB6BJmk=
`protect END_PROTECTED
