`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aF4umsTYjLYMJYNYD5u+AMEval2kpHtosIg1yz/UwrV5MGOc5aWc0xdQ1gNyD+Cw
fVEo1Yp5iD+15xxzJJUwyl7E+BO6JPe/zskb5+huyRFJLZv6l/UVPTP+H/qlB9u8
VeeGOKK095xGl2uy9n81RhNohIbfBXS99uN32Gcce9CBj/6SJ+f2I5smGF+wqCTy
rVjKRzJBIo9rYAwbOBtmh+SScvTebFEAN/1+FLXSSG87o976RiqyRJRpvzzMhooQ
QhG4FtBlVu+oLUPZKoDJcTILKLEDoWouXwKInmKD0QohGA1CP+L11bGkJvo9xhFa
c0B12k9wEYU4M9cT5TlS9fAUtZj3tHS+6Cbrz3s7ZJIj8z4Qb02lVs+fu5Dpjy8L
9fUFcTfWURsmzIV/rLeB6sFoXGtL4at1LJouJGIrOsY=
`protect END_PROTECTED
