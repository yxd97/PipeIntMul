`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r0YlHdlAqOld69bkvh63s2tata4jG0N6nVGZPZ/+WeXNUCPg5lg6gZ2sRCNsWvI2
zNWJvcnEiG/mHIL+2EEb0xAcBDWk7FlhN78hNiYiyXzT4WwoNf7fC0lYHhrQTbiP
9T0HSvo+EEkTA6CgAUpL234eapnHYwUgKK4HDD3P/qk0Qc63XFPkN+jkEaFl4pOL
HiiLD3i80HVWrA0tocysXZKig7+UQSdeojGbmD1wiHOgx1eAZEO+xl589IBaBZ0c
JaM1Q/EDmy7W3NmnHj+V/p3gyKOMljn/T76IasjGN04UjUpUwHnjS8JMntvbAsx/
sxQ9ecFo1/RDphuvrtc1eQAnHOSjUJ6lLNGQk8venEqMSx8plBVCQ7kA2aaMK3N3
m83w0Z3fznhfAV3uQ2KUFiKujCgZNlFxVR0E7pnoXHctBw6tbPYIwqPsrJVTQog2
0Lsjv4cxJWw8WQTLou9RsddiWvvI/crCtW90ZG0SywI9EfAaDU2HRIKxuMvu1Aai
`protect END_PROTECTED
