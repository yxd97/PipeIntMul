`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCoNCof3Vqp/BDZYrH9ClQbDaYIgspps9uUF/0/lhMHZTYpLPK9kUXxk4LVNlotb
X1QZJDHRLxTv1cwLOUaWkV+zO9gUWHZFhc1lyPgRNuccBTSfMT1dV1q07gEScCgz
DLD0BAe1AXFgFtQ3lcZ7ww6ApltvJrAGaeJ4cPKX4jgDgoFxQAJo1aadq6wSsAZU
lTTA5JzJvBwljsL6MK1h6aEtQmR9s5Chq3OzbFj+dyDkEd+btT5hHVVzeyMfD3P6
XHrdxkkIppXU8T3xRw1P8kjvFBtLUucu2yJq7Zm2Io5a5fYfSvtrLtyLY25Yo5/O
DmFHU76Zs7Lzu9eCq/4FDONQHhbtfXc42oann1QVtTk4ru38EVl62IVKdiGVYQiX
Zs0lQcuHMWmiXSdvKcXJQTZQ89L5kZBKiol/M5TZMg7J1OQXRA+yrTsDd6FlN7Ds
KdhprO9k1orWqRGHMqygPJ+eloVd1mqMIi/O529y1ZU=
`protect END_PROTECTED
