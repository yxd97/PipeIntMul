`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zuSU5a+F8Ar/cAegp+iTCJgxRC39pBJFcg6uhORT+f128TEECM0nr+IiW/DqB6IS
B43xlmgeV5etNHvtxaWMYyr4b+v1y79RO45pV5XbxQ8HbKmfORBTqPr/KzAGwIeE
Nk/oWokh8vrrwS+5Reao3VAZQGXqE1hPbcrbH07rBYdHab7yoyCb3oXQsybWe0Ih
fSqQffnM4M/P2LbUgieipVy+fiXc8R1wYwC32CwfOMPGoobIiCuO6XjLK3+8owEA
NWvq56swKI2yaJuF1/HclLpaOXHSkQBWsoku26daYYV5y2A7/Xc4C98qDSak3YdZ
tbZQEYaKzBW+wtTmesP8bSQc0dY1ahzGW6/tFu/9eBs8nytYfNX2cE32u8nTYFmM
a1AhUF/cv2nd6dV1o66CVpX5BnVj2laT40vl1XkKpgAyv0HXWxISiIMbioNLi6YM
z86gjTzT93t3ApMWA250HOxMFfvQQYMda2utiWpFrGRajWFDsHtVENJpc2E+AjX9
vCoNh42C1tSlgy6cwz6yZVZvZwhpP3rADvjggeXRdjzcpF84G+OC5Jue9SWkCozg
xFTq12mr/XqRmqHd2gIPPT78kkyLEveCRvQ15DjZmUl4Vmpo+fHXO0m/UVgfXJNI
rfhSuNcrL7XB5aOzjvhheMlWLoJNOJtJUr18MncfcBI=
`protect END_PROTECTED
