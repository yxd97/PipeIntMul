`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ymwo5LCzWHeDleroUSakHgm4OfQ640/noKR/KO0JsgO93bz4pZ8pgZND9tiT7+A/
Teh/gDFr2AzcWn1dknOzM8RnPCJwR3Y0J+4d4vn6jXMQoxXsqbhkLwdAWv0eQKN+
v5rA8Rl+SWw+wUmfTKbD1eNfcStTCZdP0A6exP3Hdkojy1FbhmbiBZ7BeuCPQCHQ
PZbIqlI2utvJXM6gyedtFqDFe07BJJ3V4lTSHWBi7WL96PcqQejPW4fwr+YMPDB8
TR/tHGMVspF83PXzi57J/3e2li2IquXnQkQIJHaBae6L7Jj7HiTFDzf6vkoUymAe
SaxkRRPkWIzCC+tE2VR+Cnt9GaFfP0Bnlqko32Dm/cYnFxjNc6DDw36HrTw/Z+RF
L7YJkR9VXZScq6dIAzxxBqivBlFAOTpcXAo6bABpOaqALzjU4MLgCWb416EgQ5eP
AWiLxBhDNihuUJcj4esfGU9xmY/jKUURqRmKWT7YVebqr3Jui36pu4WZn8B/E9Nw
A6QcF+ufrBqxWPU9uLkQ8MMJMENkit6VvjK3MQJoHwPp+A14f+KITZgV1haSjUEv
in3zHp3cF92w+TK6jwGryR5To/MvTssT54Nk2vfioN0ZtMNTI1fuThvBXTK142G0
Um5sqmZbJEsXEPMvpLzIyyrqtWkIgbYvXsNuLABH7ZXZPCLd3JTeErzIfKVvgMjG
MOOubUGVtCticNHd5X5CGWUO31LGD2OK8IiOpo32ja/KgMKCxFKT+dctYV8Tm8wY
7R2Fm3nXweqOM69K+se0juM2WwmJICr8OHyyQmpmQUeBv+2M8kdjJN4lHHtTvuSc
1L3an2plCvBYhhzH4VaolS89kP7KbHSs14cVMopzruD/1lh/OwTzbUlVLtXORkHI
laGtZ8AWJkyneLeretzTbTdZR0a/gpuFWndgO/1cvyfk9BXdu1haR+avHyQZiwSy
j12eLk5UFxeAvecgYHoiIvNFxv88hG3OUDNmMIOQt2IhThE9eBG7Xc2j+Q0d4s0I
pOAmYXjd0MLL9v1deCUppMW/93Q1I9cGWojBB0B6Nsz/aCXmV396e20UeS3A0Dp4
WSuQUbz2s4rWcpL0H7N1LwGtEw27WvD0O/2rIpL028VW0ASFDvaBK3bbKWtWFS/s
EnCdoyK7KYOwCLbHCiG6KCCLx1c83xSmODtwD+xYI9dQwLGRXhVPPYnRl6eD9tUQ
/O4fXxeLJd7zxxKRDM5vraSNH6bup0OJdlH4evcpthEfEcBY2pdq0praNlkbrXti
cqqSOtkLaHGWABR+fd1qvyWp6+Od28jU7/loZFbT+QxMiRNHlkRFsel8q0ih6y8a
4fyp1Kht5k2OKYCtnwdcqxQBhPLN8yXHaielTRnV2H8tKAwfH48DqLaxj2sR94f4
jQsnG48OrCZejBkOENUUmHn7Ra/pYKp+57cFi/kzNrrNULUuP6/yQBzSHuTit8fN
HmEYyNlmlXe+7TqWoRYGzrshhu82jQDebE+jSQKcxClxErne8WJ7p0t06XAlQZw/
nyktYx9nlmiyPcwcyk4FFonBfoCFVE1piFcfyUye+3CFOlyhaYEvIFhR5Ia0NlGR
G3Dl2HomZoB/2G5JGT0uuu3i63FhZd9VOQGAWiqiSSI8SgrQPPoeT/8x3A8503aL
V37SA6Q0/gCvfQaRs9zrrvwZrIBhuYPUS/yBRsc615ucyfptVrPJLX3LBFv2N3qV
SwaZWVNBtXhZNhDSHs5+u1UFSmkwhi3WXqrLYbZ3QTYqzlXPY0BPi6W24juTSJeE
fPzMtKgJesolG2Kj85V+/uKlnHU8hbiDaJ5I0pizT/eAxv+ShQKXSOlAL8r2hCTq
wPOtaIc3Z14WDV2+H8ci1BlR4wkbpGv33gxzOLrfO51LP38X50Zbb/+rI6XLCpWR
oc/D1QUOrazSzj8sPB5u+3Cq3Snmm2S81JEAHcq4N/drbe0lzfEuKP4a2kiXuVNO
SwRm3Lgq0+EQ5qhu25HjxvLJsHfxPs1bK77OSkah9thx55uVNM6kvNxzCuzKMkSD
C6xQmNIcmHvL6cYjBZwYworNMNCg3ZDBKHyMewpWZinGBwsVNxfms9I3NttAyS1I
VJozoZ4NxEEvCmZ5wfblkU6G3ZspcMwEUEKuYqqzxvgeOKwyHNBOUHfrz2LboMF0
0sWGO50Cnj6OMN39wQ/W9d7KkyJLL1WPf2+h/TvIG+LKpxOVJX3dkqOJUOrB6WXa
dOkp5nZH20Nl7pmd7X0kmSgKF9SQUMJ8kpu8Eo719hNvNBZrdeF55zbtmR+uxXD+
dZXvjRwqUynJnCM0WNCiD7deZSxjawYgUdMPNKxQeR8s0JqSfkcvWH7qTai5rpJz
jOyRV6qFN2rflYoVslLAeFCKJbQP5lnTaY+bX2ezPKgnWxASKtKv8KvGMnxzVjl1
M5pxZEigBvSCvTi1gbDdQfQjtVq64OuuQWi9eyGgDVTR2GjNPGW/UAQT6H2HbAlR
xN/a/qhQZ6VaUUChpRpoqZyPCiu+3S9bn4tNlReIZYQ1UqGscN4Z3mLiymP3nV21
Alysu4ZIaUcsHHhn3N8Co22iXk1ASq3hxKD9LikjnK7Nc7W4s9YEgC5dXOUMHvaV
vc8xNOzMgNfJK8sEjH8tlaXSuDuuuKo7kgz5RWsgQFPtHaETa3aBqSMJsVNj1shQ
0LRnCtQ7qRjCGuBf3bpoq0rHuBxkigyLB4LR/K7vMrd0Zec5aTm/yJ8+fZYMNsDV
tFrIpQ8g8p06md167ZLUOg8qx9qmgAD6vU/yURckKgr6PAwtvA7QgzZv7Gy2bxdr
3vkeM6svYkqL8vudIni2ek1zIwkxCeHWtH4E0fGQL3ekMEBiZZYG/oziVQC5WVxY
NJI39JO8EHtpCleJlxYeEkKrNly3jfy+XR/9tkYWvTH1WPA0XD6p1lVZREqlr4iz
jpv/SnIcmk9/aYS510K4/Zek6k9GCoVtAIaBCAQ1OegBiDh/yt8V9njBLawR+y+v
zBahhGgvlW0W9/lULJLM3+dpPzup6qBRZnW3wG3JVRoaJox6leiohf6wNQ7fsPCx
Yt00fVlZFixV015AeYwuk72cicRi/UQd14DPGd0TWQw9ZF+AhLx4i4JAP+XoUP42
VGqxaKDdq4ToJEvctViPtvPRKLqxHMVK86dx+wxKRhfp6ua0QmApNINPm78tBYoC
xolcl88kVXthKGTFHH3fOhR2DmZhHq5qPOjmNMv8CykbGYw6+z/cEyNBm9Bor5V9
fSDYHIi9RSjBGmG94muByLbnkvYFSw8NQ9/tWnEkZImNykP7bs4K/evW0xQDQ/es
biU6spdn7hbusegzBzo8G4cyRuODhAmKfN6KyalmArtRpk0axd93F0nMj7/IxhLH
dkirteX4JVwdhydXkX3KiHP/V5DDoDdJvX7J3WNB0WzGh8aPxReK7jy7a23SmgWO
cI8S9OTAmtOkHTd4KsiDtM33LLqfBocWVUHalAQnLSVQ+y4D8aNv3uQH/KyfEfMC
g26hmBUs4qBum1CsjCkyYqgTH4YfGx3iZy9QosTTHBpsfqftRKXYLPmEAslPwSWO
edpLrpTbYsMSubfNkG6d2+DG0Puew+Vbm3zGVw+OCl868p0YXXUagzLCIsF1apKD
It7elmPOyzylQ5W0lMZM+1q9Av8lBpl64mKhohEomYtftijKPnB5DAnn7tuFJ0KN
/umb2dfnU/l7KBgr1U8keZYkWS9dNvtlrtEHGi4AHrAJTK4ZVAz4LxXGqoGxcH5u
3bsclQqkMkKzhJplC7F2xVPddYasVhOZVUFv1/SdHVWndnz673PgnIbVN67H4OQJ
Zcd7Ea2Xk3xpFrIhDfACnQrMP2yCVQkuj4fREzPO6FgMsyfz2TkM8IGxamYbQNmY
2WaumU4oQQHYrZjEjACTaAU5LJhe+IO2KxQis5wvmhiq0rbvKBS6vbvpuqlufuEG
+zjUBsidRCgWSSjCJpu+lsBLDq7bk4MYBch9NLrPVGeBmJZZiCWodYhTWshk99Ds
YlUbW34U4B/pQdLzTw0Z2d3KkeFlzUOghVUl8c3Lr3pNEiarMOz7RdmgJF9wnjVH
xF058gEN+XBA2wnhMS6+laeGwx0x845+U0pBvc43Q4uxzp5Tc02kjfYMf4G91NEn
fKv7NrE+4b22DOsgD564/U9uOXNK+WKDe1tr7Mm8XDM//U61MfkiZrKNMnJBJs4e
3tc7/piespTjYi+G9NOEeg8HgOOBT7YsXWoT3yL8V06TMef+Ed8Wut/llHsKBTPn
tfpvgWue6nIVtf9pr1u1bmGS2mpny7QCexSGOhkkZKdJ2Ip1WYPqVezdm4tUk4T7
+tzk3i/TBG6b0x/9qbDv9sdcoWMmq23YMr0Zdnwkd2hX1/QBptFIz3cE1Io3jdqb
1miw9ZF6YIykshVhar1jLP4Z/IXl80SU3LblvQod9l9rH+SmdDgYCo+bb1y1bORr
LoFB0IgLuHFblt95/gRXWzG6XLS6deJcivtizlqooMDY/MNwVUzNz5icdiOwDpri
dja1AUBce5Fg+Tr1PhVyeUVC+1Iv39AIJSYO+NV92d0qqujGgnfxFKMpBEcVeniA
fofSKlqbIQGgAuEVFoVCKph+qvPs8WNdUUTTTygI8koDXFMTXZCx80ASxHji9Pvs
6hmlq76u9yf35Pxr0KXFHlhF4WxKZ5vStrOSi+F9AyfES+X2l2IMGVnWM9WjrKJn
`protect END_PROTECTED
