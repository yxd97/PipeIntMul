`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DZsrQTg1Sqm/TdlQb1U8mdyJs2UV7pYoc2ZWUwBkZscepoW0fCC56ymzlibjuQnR
siQt6wtgrx4Kw7/hBgqcDSQMCzZHUwvriSFubL6CiC7zHhJiRHaVcBuhPYZjDVVR
sbekKoq+lS87YZ8I/WeYKO/AVKIRaNmUFi0QDWMcB/0wJHEtZvuT8Xt8GABmsupX
Ts7I0kDuRqnftxyZUZskZKwgVRrlBus0VPxcefN/RLG0Gk0/vrlGXJm95hchhqXM
edcnbR1idHvaPvXPHQKp1hVK9lsiicaHdWJsbQgQKDqaARlRLLfdro+9agsjgF2h
cJHFKFgpsExI/nCzp1dhGQnZejINryBcUVG4sKzo90ZVbBmtjfh4MvfABt0tSL5n
PrBYSFeF4PiyDstk9239uTy78QumceMr2E6tNSMPLIk=
`protect END_PROTECTED
