`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3v0FuUMkpZEGq5Sahl661L0ADJPcYeHjbFmyk1wMceOOmI9N2fuYuX98sgd0eTJW
cSxJ1Uswqb4tm4ax7BD2cRqtGhccOANIzkn/4nfyOSY9FxkcMISQLjqSPFLYPm/G
RELF3twnFMoG43s+bCZca4PJ2yqACO9MYpokTDaNbuac/sBKMI9l2FcRchu6Rf2C
8CBmIItzoptiiY/a2mTQFYpaKXRFqJ1E06LfuqGrsiNcPWXgMo0RS8Nn76Gf0u05
3p1O/iLP0MPDSuWMf77zEGg8SULCFFk2I0CzWNuc3Ic=
`protect END_PROTECTED
