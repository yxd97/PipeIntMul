`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bIiP1J6w3brXHGFMhZDRq7NnHPetx5nxjHY6TnFWK9GXAaKOJxKgWY0XIpNY4KRh
WbrJRmfdSBAOP1KRm0pYLdkv9x/Yaafg81+TNZ66pZXUVAU5UmDpQ17UD5Ab4ow8
9HoRqlMiqYCDE9Vd7W6mtcckyVb4NJhHCHCsZaHtDN48Jxj/x0sQu0SxBmq5p5Pe
N05XxqwybG6jpsTS6zxZAOeFKimNBqKR8Lv2yx1UJzi+TjOeSGaRvWPnPki1yvAd
Zn3qw/U7mYkPilm4mUnzkoIikp7T6v1S0UqbB0UBMnMzw2dPoAfogEATP82Bzcks
7mY2weHKNmkbTXoCyLn+lX46TcTCKivVqht5jrgXMp32+XIfLIvALkg36AQNZFq6
igv68i1iAGKrnmi5xMsCH1w9YbixI56R5/L2mj5MC6msUcLLCI0yvh3p7NQG4Fg9
bfJiaCAPuPSaXCa0bXUIb23xTa3hoL1k6svenneOKlU=
`protect END_PROTECTED
