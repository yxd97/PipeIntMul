`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
32l/QA6TTclkX7kbwzlgjFgpxrJSYkZo2u/QTPGjYB2PpcVtdthU2uuRx9FnIgW0
X8u3Y6Wp1RgDti4p3o2b3FS5EJCYweekTDnesWu2kwbB2mxTwbNbo1SiA0n2Rm3b
+LR6axX3AAxQbeVm7BgXUeY2lrgjEzKE2DPFfEgZyvpnfsxt/ZFx2lGgLtJELhIB
z2FyL61dV6Buownq6CcEPX7AWYPR3/LfsXG0gQ8DqcUMQJHs5QhyCzRCCsabZb+M
83De8frTvdoP5GXRMupQQH6NLDOSg94j+pcja9nDuKhkF4SG/B1piO7trixqxHLI
w6RaWQTFHF0SLjEexhpA3nghK+eOOpIl73+HVCsXpIF1RKFYeJWZGZgFgBRLebSk
KTUBojdUGmpuTG4XRPADK/RXQVpRtwcR0B0QQItjtSz+/eteou+N5xnS/J5qGcX1
`protect END_PROTECTED
