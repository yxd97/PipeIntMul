`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yHroeBA6rJNN9RqWRA4c4aNy1utrRKt2g928fk/4JR0wxEJLpcMwZvDV+FFF/7y
OD3bI79gGm3DRKOx1FgJ8+PWxX+8Vt+YDWWX7P5R1ThF/WTZ/0G4xkF4KYH/n8es
Lyq+vRtbLJSCU5Jmg3a625oFO0qBZGNGCpKJ8LEDh2TkSbzM8fmpNCA20KWTNP9H
IJC4kB/M1ey7m76HsDLo0tCspxfe5+Y3jIiv6xmJe/YS6f/K8ZZnR3uN4lpQdhjt
71tbDhz8UoAEHelwmAqnZOqh54AnqPPgGqkQyti/n+wnbgSdSIJwQsbp9QKaCeGI
596eWox+hFVeeS0eCWfBIoflAvEPyBGqSDIalDfZcZw5biKGjyYAtBymMorpo/FX
ishCOozh0Hr3ywBfEDjuzaeT/pMxAzMhuO/F1/moIUqR3MQnGu7RLlJFj3rFkLV0
Vu7UDxix9Offw7CynM47o/7cZriiRvSTocBr/RtckiyJPwhKvUgcCch5rSPLFwQ/
ygjgqLasziTjT+LcUeboYeMKxjKZ8G/K2aM1dS3GRi1f3lnqTp6SlLTkRzDg1liB
aCrE+agfYHS6hZtIl21QvxITFz1R5CfTchu5fWe8KW4sOggUl0I6ahvLOzVkOCBy
EN0pHy865l56SyXS8ecND/i53E0RZOC9Ac9SzoS3csiRnDz1SYCB7pAQ4tOeLIw5
7DzjMRE7uw6VXnJu+9XT6UqHIsErT/FYR7ffWx98eWY/mk2WL3kDOLL5WVSyVL9T
4ytKB4gHp/Y4WuY67Mvhi7IaVf3W6lKkEu07ae6gOP4hIA08hg0+7FCWSmJy9WlJ
47Ll/adDLREMpS/JMESCT+hRCWLJHcAbCAktr/wFjUJ9vhql5dhdcpymlwER8Ggn
Qky36FPKVEmOkz00QrCGByh6iqy+FbP/QpYmvMtD6Knwm6RxPoZj1hR7kkYnNHmN
4Cc6YDCl209lYuYLj/ehkBfIJP0mI0S+7bgPUOD0+XyyKHTIzZTm8Lou4KkC48a5
X/LXGeggCLOfLUT5U8Y26GYzNvwd3SAaTc1alcG4bXXLlCweodfhz97QB62+WV3z
9uE69EWRFsS+B8yyaMC9obyz7NctcJkoUC35ZuNfHW7zuPxAKAgm+QXpMKa1LCJa
lQCzZ9+HDXGhwiBSj2Cp6Q==
`protect END_PROTECTED
