`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mbvdhwHOaCJlro6jxsrk0Z//LxsiFDyDZOWVX6AiXsrbMA50K9TV3R2IeQw9CiCa
yCwwYs+6sQCEhiKYLjIX2pJP0tE2dsgCO71GT/SWjhBrQfHclVdYnZvNjJ1maoMH
PuYQglUnu53rN6ePKIZr32yIyBSR2IDidgE64ir5Gs2AYOBd8n9D3Kec+PB+7Ae7
WnH9Frd8cU9wSG5i7jOB5Pnst6t4g6191SW89YZEJD+oW3CkrCsmRm4MNJJ3bdn7
lOrX7YmA7aq7imHK17uVE9f4E3Yp7QhpKQIwXo+jlyJk/4e0QOhruTCvpXW5xDxN
OnmCsyuDRU2NTlhYImtpqNCKO3WRU350YrYCwU5ojU4=
`protect END_PROTECTED
