`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zb0IzbSd6e7+ybslQ8l1meV3epzSnbKfz5D93MQ8NllznKS82khUhFELxRgcRzZS
EmSDK0Gr0+jF7d0aC436Xf6+bvPU/RapewW2kWiu0cE3RaIoaGbWfTBUPWAAWbaj
lQHEswq8dd0I6lim9BMsjN4xEOq7iyzaQwhXHlpaNVGpdnpUdDYIJhXA4oj0krdO
g33oqr3hx+aTU7mtefbwXEpee6w17IMxuBESP6l8mSJURbsqSsFtPWQsgzOy93QJ
U2Uv35FOr+7T6BqG0HXAS4+YQG/CKb/SirPgEJtx+Z2cxCgeoX+26Hl4gKwPuRPs
m8WzOaiFWgplPlOT6NuECWSz8lyV7YDGzfGx+6TUaGfxM3rMA/ZtOex/wINLGECx
bcU6lTpNrKhO2Bt/oGIM1KoIcdZ5cTIFLBEPwDEKOfuPOG9iSB4lBIqYS8H9fyRF
CnQUsljKPgtzk67qkEXIZaVAintHxL6G1hLhT7twxyepijs1jMXFJIRUc6t9Blgk
L8Q8byvlDy2nP1G5Jf3lqtaLZT91Gapztwb4CTk5LcB3jZLdsAuPHjq2wFCuH4WJ
nv942TPxL0t2z8hsuLOcNSIjP7dN5BjhSe3fELqMXPkhah72lCceQglqdFpTEaRw
oFLegbqRvhAUVUg4+FLCIbC+5WbwTWVIBT+jqpunG9KjdaNMVwQGclFHE2ocVgiA
SGUEPVVIjoYsV5ep8P98bjpUGZ9IcsZ/8LOECnKw2iJvLSqGTFK72PJGWmnU7cZY
AWU6WDb6o9vC1g6XF199BcM6Z7uFWR3VWQVBiKRyZsEtkIuze3SAacHRGi9iXJD/
6QBnP6j80XV7Dgr2ty7OIdhaH58D6fkAZRG9QTURSbd6281AvIvFoiIkCN9CJw0/
XyI1K5Lpwpy8GqUe9n7HG8GeJnATSG2BuCaK8ef5wIVeoIFwsZbmhKXvzvSOdM8B
8PL0Sl1RoPWh5tyvbMF6qw5K6zmhNGiDqr3vZUvbJ1fmBWjBTcHfwvkWZ8Ze3nio
N2E/A4zwUzJU2suWKBWUYuYzz4sSJ/Qqh13izkgsXZRnIHXaBYOfi4gV2Dkcz4DK
f5To71tVb/+gydfBU+FbNkLdHrW7BOpVT9i2h0XwgBoeUHRzojr3VN0oIhx1KtpV
w8XgMqnA7SlSqbxGSKsyxNWFMdGVnLwhYm8ygmw0/6TOuZLmNjh8BzOjkwndIrqi
EW7Rz1CwWUBNhaB/18ksNhPjHQGFfPilZ6/A5T1jsebWZC+dRnRoiYRnev1L03rD
KBg6V6Fwba/t3kkHRo0loqlTuzFPHc9Z5cGjXIUKN/Nw3+ktCGJMrgLOcnK2cxJL
yK1aLujaC6eBqiOoW4zI1f/G4O71BUjNexDCMYeExO/iaQY/+jX5azAKD0l4KSQq
YKJ6FhhsdFP4Z23G85u48+VnUpiZjGmUBzVqnbWAW7X4K/THs9J7b4L+2mkx3YPb
I2s6zBfMnq4hMJ26ROSzOOdSwAk24/VgDElHlDcAUtFZ8tzMogJ+kOLpfOUtOpEi
qPq/TuLaV+CeIdAzU4afyy1aYkKq9nOp8r5UqYA0i0o4I3b99aMJ3KCoNMEOp4fn
HWHAwhUxX/sA/YcSzpGh6yotU3zPrszssftxgm7KU6FPAWEa9V2l944bKK9QmfdA
lvRwpXwZVPlBxk2hs3DH7IR/ZHLdcICYF84P7bjZAZThoeKcTEhbAUnsn9g/u/DR
7CaS6O8ITV6XlqDcs7CywS5FXUCoHb5wNVgzNndCCcQlcyGC9jvQTFeVwdfuBwE7
xmXBmcXUXHshvptPl3hnRdZ+ILX1kcmqcHzKCMxpgBUwqMsv1YzRKOk0nJhxoBSU
8lYhz7ZzE/Px1iWSfWkrfCyJfcd6Ub1oMr84/XYJcA96C+ycTMhL6J0TfMF57G75
i9MssFET9eL6QwfeU5slBIRxL7G/ho3TSf2ng5mlxm4eWfN9Br5Wmi8FiEPcvwzc
Cp8AFPIVXxsPCC3LxEC7bN3Buub75AScDSv1fKpFmd1Il+bVr7q/sXz9qo95wHdl
XqRJbFNT0WJ4PU88ojN1x/qPzSWAmmtCMEm2o/WoXQ8Bchd5qIYMvjtPHqivKp9x
Vn0uKy7wESHaHt8dw9tkaMGPO2lZdLQe7K6/WIOqcO18bEPedd+KmQM4gv/E6cK9
lVtxEBoQHMR7XTL0Oic6fDRUz+hYB8PfXU0hQ9bsMw6vLhNYsUkGnSnhWoVW8/KL
tDsnR0ya/D1icFz1+YB/HcZjLiunk00JUTIWn700hWGDQ11GqarrTDQQ+v7VqPXE
AnIPPcEbReX3mdUdZZn5Lehrk7v/OiXxFkCcndsCvsu0Eqx8Kmu0IhkhDyVaSHH2
U7L6GRfewMRFzNWjk69/Pudueyi0RGsKvuRnbc9bm95WDKS5PYvJ+lALoCDYeJhy
rs2fEMVH/kPqPXmvP9shaOmzziZDdwm+CIFlwma64jJHVUkpoabOANNI9aOqTSWj
+LJm6RfokTtKBW5/LT0X1hwP6FAeSlZ2VUkfUGLSbArWvUfQRgJkgFJ6+3hGRNVx
C3o8Iky3WgcOeVvHK/KRLrsqzc5n15CIlc01tO4hrhcuKQGtXIBCS/zk9CAlhNv/
EtvbYXsSIn3vmQdxKhN/MUl2MMr/Y1sEOlr1r7j54PK9vF638IQeqVRaMpRA2vpk
AfgvnDZVszJcGFY+cMUrUH9ilXcdBdiCBZbOslUq4l3yYCj/MmbzhpA20Z6Gi82M
0Dm7UM4gepWTGeSQpaS4mOqQfRXHtkePT06d3b/hy8dCj5DrDg1jo9c2SMDDvC1x
nj1klC/MnKdd4Hfd6FuhNX4d9WmkZWn4J/kbKdp0qmdsCQ7r+4nPGvshuW5lHp/a
AyX3c0L9xDLrU04IC0YRTilSrTRjYjkqSxF1PitQgtbc2JMSNYe8zircaAmoo+JZ
jpJp0aRmfpfhbCKb3hGJl8kgfWC3+AJv6pYwkrsh9bAdfSndpIy3Uf76cx3OK1qe
+rmO5UU1XeriP7FHvORhLxELmgSNgJ+NGa6RTB7TG+gueTi9NjTKIhKkETSrvZfg
N+z0SEio9JH/U2uu2n6NJTfwHAsfIy26Xfe+fVAMVq1YraFHF8OIFIzLBJHYL3J5
Wb1l+sgcAGsy3jriy/WCCIJnCvSLK+5FzvGCuOUbKZk0wkaHBeR0Wu7276Ua69BU
O/FIk/eM1bLX6mj0UT1ToYwp8LiDMVSBlVwqVDR4GQg3ud+FtOmtCNjN6hf+MG5a
s11gCsINHjfxG6AwBB32jkMgD+B6rIBK2BHkirKMc6xdoSNXzNd5O/BBptO8Qh7L
2fxNlgynMvx2bDOmEx7zJmctzORx4+v79R/TkWdcjgq0pmDxR2Pl76eR2EuHQ+GG
wEZWwgElUJ8RP2SQKC7LEW8axTAzkaxuXichLvMKQuPnCArynGcsoxlYq28/FYKk
mrH/G49pBcFcjnASXquUNv35KsRCX5SlBDdzhkdqkQM8WZX/9aCGgfsSCvhbliT9
JGPNY0HqJNkd1AjBX6AMHk8njZQuVg8G7l2Eq1slGMd4rNDcCWe+6G8UOcvOU2qw
9AegO9XlO5uMPxDJQcbAHqVcpfUhIMAEw1/9dIsWd6UAHcBuWfoibBn27+DZusLJ
SUedraVEU6TaR0lTpLT2kFTTYQE37LMdQAKcIo1ON/4TLlavkGokQI+zhknYismL
mvQiUn1RiPUh2ksj3pl0dKM0XoqlW+bX0MlX4nEYogW3lqbhM85SPOXPwgX9H62t
ZlP7Vl4evnbr82xEaCI41S7wIqU78buj663qud2WvUEg8t/JpcC+vgQU8WK1HRzM
LAaJUNt6E6itANDX88ajt+jQ73DHkJMsF73eFsR9WqvBIWyyrdzxMlb7a/+5R/xQ
T0N7LKZF2v2DzBJl0rh7fNC9BwTHumyTc9mk6xo1RFsIQHLSGulkOfRm6bAVyOfC
dZa0kh8pogwqCXxxt7yirz1axT0eYV2e/kDGVyqcNhP4JQeBNDXLIGvKifeVNOlQ
zkEN6b6k3YRZw7mRPcripHHYKXpr4KVgdAj5W6x1xBbcxGZ/n3eUt3XoVydN9C1G
+I8ENeSwP/ZS5a/Y0y5tb+lzq6gYk7ZFfz3Gt4TeGu5hGXedZXrUhbiNJGif1fwU
DwgGXCJ+KvkhctRfWc3xmOQwv9B5f2SNObceqEbgBdGhtC6oTCYI2NYX2EvUH0hg
ArLuoK1J2q0s2j0gxcHMH3SRbQDYfrn6FQ6mWPs9n4tCkKDENbLpYck1y7WFO43P
04L1qTWbhVNXvj35py37n2d6uk5T2EvRtCi35nv+OG4gikxF6HO/rXi2PSS98/AH
uVQtdVwapwc8v5/hoRv5obtMxApg0oh8sjxghZZ8gg//RHCR/sDzpOZl2yQS9HuW
U0biM+BRmT4AG5x6OYsMndapfqfgGmEyFQtqHLVAA/mpbQjOQ7I27QHWjhhSwZjG
nrOT9jGqc+wOutyqd7T6/PRs827vIomAPnCOeFs8EvgPs/cr/R1xhyKVgqdgVeTL
d0BBxvKL1800NIA7Dgif121lsBA3YpITt+1jfLlsIJhofExQlcdDrHbUue1OYjPA
RUf6ocV8RN7gdtENV4CLZ+m2zlp2pzmG6fvOLyatk8cNIhHUg8RN2y7FMXqMJK3S
Dc5k2XT8HH+L67+iov9jnSbvqg+eslE0LlDab6xeCvGMbC54yLNK5196u7cLk+ge
xPxwcAejh/XFHXEj/GirAX1471cS767YzQnVyMg6Cyyjvt5L5ybUFFfTKU59w803
Pr66Z+mMZ2Zi96vxTqeJ9HtP0KChO/+2vlvZ5BjIPVumPid6I4ttYKLan2CrbKkt
+o/nNVN8BKB+QmoaPTxXn93+o2rqwFSqxJYOxcAcsyhWJ79PbG/BRmGU1pVnDjjg
KShA9NdjOLvmYFja8Kxlsjv3kLpV/Q3EqFckJYLctS7ZLu8vXceinvxcjTEr7d8f
O7zUOBUopxcbrvg/+dO4Sy84AYuGABPZkjWMkrE0VtsGvYg4L5KcgSplF6nMlcyQ
skCAn191hJYjc5qRLOHXyo253VuK0gSZTA4SVuHYuXSrnjyjfoJE1GMZOOmNJUNK
gRX+XCAYGgXnqdZreRIxyjEVMJQ5hOZ3czBN0PhFVOo2pZsW7mR1VqgVQsEWUzkr
1oC7TDHFnAC4QTrgoKBmEaaqMTt/tRCT5tFtAaBt1OxyyXZRErOhLpCmpz652gqh
FKlM2I9Y7iGkNkdY2Ilt194auHKfy0eUstzJo9NcoIrARcPw10SK3MkDApbG9qHg
qJcg3pa73yybqCsqsT1jILL/fwihXgIWCDPAMARqCz1tkRTko9VfUsE/bioUYHLj
3lNAVVCnPDZq3hBN2IP+UOR4sd72dPUTGN3G3LCLCPWKbAI3yXI993KGq2sBWI4z
HLXfh7KkIytrZzP2pDFO/mZdHrMLWVbqeoKCEr0x+AR7+tqOcp71lkKqI13pe5Bt
x89dfIMEjzZbsA1xx2290bLUHy0LZb1XIE6SsG+yUINO4togAfiC0zw3uFp8M7Mx
eze85ioLphuWfY+dJ5qcf51OLWx6Palb3h55P3Elm1AaMNcL8KUQJP8z5ImydwEP
cRYPeJUB0Bo7gUhzNZ+Wu5VrHYAZRf36RhLgvEDfNVDDZW9DAkLh6XwIXq5BsJu4
Xo6Qz5mvOVWgTDcUYr60DEHtqFB0LLG66QgeNAi+rjGJ/gefw4CWIjFs2YQ5vfsf
O+UfGT3fQkBjYBRucFLDnmF1N32pF7bxjOxxvIRFJJARs5Nuzay9OL/jh4OJEchj
aoP5MDr6v7II+JThlwelc2CsD98br7QCJ05AMHKyXwqXeiU82H/B0yhcfl/pX0XB
hy7Ac66XNStMvyUqr/Et/0E1UDVPTj/zUDgDj/dBMazQ8sFZxtYfphvZTg6JUs76
L5S3kKiDohlY7u//uD+hEPE+Lqno8yLsXO38o5TRNREpAbjE7sAt4mfDqOQ7+ijj
CDpK1VhkUiAkZNkthqkDGNXtWszY16yhkbbufWj0WVvK3VepfI4CoL5n4RIN6pVo
FOyU0C1IxHtugDZfGZX24sbUo+RYeDr0Py7IjWOeC8P611n08gsP3c/BOkLH815l
ZnadwpMkrELCAmRsWcbsw2MPKH8daLBxEaRaR/ZAILaGqRAynzUUIBbsoZPr1QUN
/0AovGdBSw3zm0t1W5lgzhCTRqMmGVq3ORc8XB1QZ7mJ+vof6wXsD2Qyzcjm2SN/
8av3vCovqOQd6anPGI8h2DKqSfhVrj7mGHa9riQvFUc+Jif4mbGyfQ9uK9PgxG4p
luBSGwV0II5Jfi+Z2h1yoNw2LmipG9Vjkz6MaiAecQgVA0PIBOlQYWFOgft/bKge
TQninGZa2xMfgROxqEaEVFkcHA9XRcnMWfjXSQo5HqdsLj2Ulo+jflfgDW4rLVnF
M1a9QXF+vkm0f8wN1nxKMjgh9YT20BTYi6YgKbZsB0JD4Pa+A9J4e5g0U9H99uD5
Mu7Vpe5Jumb14wEULdudkhkPjDKt21VrL5BeJXEXsJ9EL6B8Dj7Ym6kHMfZ3398J
UKvuOsFl6a0LY1dPoF9vNZEpNJdENxsB0IjEf3NU/fvTvatNhQ7L2Spym7UX1qO8
T/1EEEJwn6fazQy1M9C7XpDr6oYYMcIz9LOYp466Ic0xKC1YJFnA+cgF++/TfNzt
bbfVnyNsZyU4lU/tXr4z9OKpd/ZgMbdizmTnPaH1H4TQDw4CZnHVSPzNRc5u8Cw3
fARjlLLy6MQ52MvXZMWZiP2GZkilWBbY84yTwxMgFz6btz6HuzzfONhW/PEyOhpv
hpmvFXk6HOGf0foS2Q16vRmAUua7T6rw2B6WexhgbD4vS75G23Qui5oMP0seQRpc
MASc5BX0wtZDheq1E71ZXUccngECx52q3TIoyn4fFbGRh6JrKKKd7GQN2Njpz5Z3
hk5QeKANv67wL4l6sQ+hkFj3xPDl+DG+Y2SqHG1wsDD8xkzn+DJeUZau/FHe4dqn
NBYzExZCzl/QsQLjPjiGTgyq45nmhhIKsg4Yzja9Cdt3OCYB9BidWpRlZreYQZKf
4o4cfspHXq98/Io0xTD1kwL9RCaXuFus0wXDaBNzwWgXdTWagzDb98u6iSfZoJ5j
UNgJRD9fegKsgqns/hD8etWLOmaN2KhDasDXEcDzqeZMIdRtWALDRaoKkVjP6a71
E161uC0Dfh3bAT2wFalqmwlXp9nJUYVw2upvsU6FqBmnt47mVt6dxaCVNkfFb0+R
gUr4ks12xe5prhWgcbti/4fzwp0HabiLNcsAkBbtbLmLcvM9NVLl8Bqp7PyCIQx9
dvU5M+mK1/XZiGwTq0KXTBsRs4LZOQWbirq7TQRQhOTmGKDeGqjbKAiC3/SlyxE6
rYvexcN++pB3wMPoXZUucA43SRDsmoMiATJtEuWtb9MaOZqMXSmAW8CXjPXuwuPv
7mXXt22cy48tGQ9L4FhG6dd8actJP1Yl/AAdiYOqS+ngkpUDkFYiZfglV7LddTgb
n+zvFDytec25eyJUVRlS2SxLOynvYRFZIqsRoCryzcomey+g6V8G9oReFf8pGlNv
U1MYq7ck8AkwziTpKLmkY6GJdZL5rCpS4jXdMkGL0wD/W0nPHkX3yrkIIrXIHtVz
fY7LA3SQFF1jcDp4r3d1N4ye6L6pJwJjpbanGTZ4d+gQAfo8pZtNEMNGOQUyGYFD
1hOS3EsDcCCdPX2KfZ9LmrMNwbGZ+kIsGjH//ho+VDznEhni3CRBsUM+0Bx3tRFY
KL2lwkrJ710+TGdm90WK+E/9UQxnZja8KJOGJYSRIr1U46t04IsQqzV1gixe5BcH
te50qdY+BIfCCFp9edgTUgyGJ7MnZLYK60h239NJ/BFA0O5IhXp7xnlNtqnh0JQA
JP+yIM8JSLIJNKSmfOf/8WHCQQqITuPxCurFA8w7Qcz0G9oyUcrlK/c1lOfKgcQ8
9IiqSAqi796pC2456BtGkAgQQKQQ44l1R7eU2EOOY/sNCJat7tC4TJO2z2trEpNg
OwkIU7mmGFb65HwoxjwfiCAXmya0ElpxGT5pMObVGPyZww4dTGYz5EUdj9JMDFag
cWtJrQcCBH/TFp+oFBCWpqlFSSdo+TozCRZALy5LwgaVEMlaYgMuS5Rq8KCUxd8d
pypnilPWgQOfrWvQmlF6748aJq21iq7WWpao8A8wAztOIEeyyRzVFZHPqLmodtTj
BAs4aLHxdw6+cq63+i1BUcVzgG6VNvT4DR7JwjVL2cZO5HojVPYUzXF9guST4uwp
svt8tlVRZ1Sz7Che49AL3oEcjMkx0tebaucIRsR8NQF9thFB3dPctCehmXK2xpxO
VAPT+nAH4UA9vv5HAaIC2G9HnNTfGlYiprjwVFDK/+/BWttDQzWPmo2E2uGiMWAz
tNtrqEJQzr0du/et9QVSRa2DJ6JbI8zj2ymZZ/C6/KB/heB8iV0G+oL6Z7Algp/8
7MavXS9z/QKXR8TrflkSIkPZbCV7FV1/S9oRHW0PPSnjiUY3JnmP50ojbj+jgpW7
wLO0bUxgfWOrpnvNIAHNZs2igAaSqQCM5Ir94ALwv9CZyde8u8MZM3e3BZRZ3PEd
93JtB8tAGr6UADN2mYdTvyqaCHn2V678hcvhXreKOjlM95ND9k0T7AoGSLXY7nS8
ZVXZtAWOPeOLn+ezMy2tKnwuk0lO13mAY4nmziu+U0e8/wEjV04lp6+lXatoAViE
JGf63tjao65vpzAXU6wc66pPTxBOgf7e2rj82shB3ZkUEJEVrqwKyPrsdZDvXneg
4bE0YLYbg57krl1PR0K0gFe6Z1rf7f9kweSW938iL4yDy4YiIh6tc+a6fsiQSLt7
WBxv1DsvQ2GOD5e6EPHoRzjZsBxyVdiwpUDdnbKT4T/nZyyCctuwQW/qxvzsjc/J
idjpRyW7rJN9U79TAFdeXmaXYiQ6pMJv3r9t9ynK9E7aI4+e5NW1jKKlj3qBdWkT
qJJU8qrzWCIyDxoMvlnd7uOUNYTuW+fV89Q4n7atYJ3Vy0dPHy8/vAXut4hs+uTd
g6QKPl6l09SOPx7FvDbmrRV40COwD/57auIJfi8aKbDmxaffTPtuUherBL/vgfaK
3mJv5ykbTTRr6AIIeMTVkJiX8weFW2lf1nWdZKxBVMSVgjN+JlYl98j/ajysAHav
i9KctVNYdZw6mFDmwbJ4tECbHZmReWi0f4POFedtSaiaxcW0E8k+sm5TahUcRdhM
s2dlv7s1lZtanm+gAjGDerqElOFd1ZBDAK6Arp6YyPj4gvpEjgCQbnB96tHHc0yu
8eKQOKCvy5b8y0i7v3mv77ua9qr3xjTqaL9Rb8FHAt9K9ONI7eJJ6b32/XA1aMZi
j6KVG7lI5AVNDGEmunlrWk/9leAGdpuG9+S2yAfpWJMNb68Y/qyhEqdMsWOqYCA8
Szv9W3JV56Szg1glk293YaCssa3baqsodtHLPJzOc1sow7mikDV+ndx0a+16LrI3
c15/mcSKBtxK+1V/q8csvaQ92BPEQUuAwXyrydjbDSWIMBP4PVCSZqyNWTmaWPYF
rLWlYv2BzQ7YqhW/Nzz5/2ddZ4S1deWWpyAWhJth9AA91ve2AuK1MfMvwp7s1+Du
Z1qG8fJX3n5NKJcYxW9WLPIlDakbxrqHlp6am5hjgGAIvNbUvmMOJ0We4Ro3hzZv
KWzmjUEqmatJe6lXGce4ONhDTiBxmKvfOkHWyjYR4Mj3AVS2OXm/9LJzDoy7IyEJ
lZ80fYN/hqyoYJ2YiTZo8UkqPRJdUml+aRoSosu2XyXAXw334eKMip3nYx52xtPh
izTQKImyipXR5DigdLbUFE7wCKqoA9jElDAq/+MPizoLu2mqIjB/kJG4DYlMlbav
0SEDzJt5vdPhzq+mdk8xQbmJ/t8fyivQg9JA4XY0gfPJ+jQ6LKhBDbn8NjA2U/Ex
dAkrHYx3oOH9zkPflGFdD9LC7f8Xfbm2DA8k452gQbe4Jioc+esTsmgshj9+SbNV
JNMqLaIAEmYCqZalTyqTJyqFG1PrtTKrkOQeelLa7XowItWxxTySdcHw94FQSpG2
OWEG6aaJiL1ascrGruBiJs6eV5ksryWolJG4bVmmOIBWSh2wsAVuQTCxHVb8whQO
ioD2hGGzZYrTKteulnk3Rbym03NnR0FBbHYeNPFT9k5Fsmcg8apiOIxKARX4WQYl
WCzjDfrPKtmhxEP+AaR8kHzJlT3shtV55gqb6QqC5Wac1Z+ZL4kyRtWcHgnre9OE
AbqHXHM2eBoEkJJxxD51DKK/t7Fne7lGj6uOYMF6lYv5w4OUnnQtYf7xUoC+OXMD
nKjClS2SegBblja0aEpT2sj0lJd6wWBoq0FlXOJ9yOslkVcZyYtc9Dp+zZUNlO7j
gSOPULyn9w2cNQWr91AMKjgxUGtoVLKOqyfMwG3vKHfSmJnT+KW3Lwm9baVLnmEt
/0rmFIXHjlKWPMh4Kt3e8SkbLIfb9LE/+i8nDVtRQjdzLIrYiZXvr5/UWJtiRHod
oSEVXqGqNjMb3V+UMq+xc/3iSW9Ka8djZWf48bSw/YoemeG6xBT7tO6v6JkFFHeO
ElOTtDHN/+TfH9SpYFOISrSi+U9NEKLkR3gbrJn9GjnqgtxIZ55mjbsQBF/RfvsT
vRs6TelZxXqOF7+pBxBvieOsD04AHUXRcL/010yPQwUNTsAIPOAkdpCIg9Oywk3Q
wj+yM1ar/yYVUTdb/xJqhRnq+NpG4cGjLklvAHvhz9Bd9rsSurWLAMv6/x0TVMvr
T5audmi1FI51dr1wNyMAXqT6Nrnnx6BenDbY2lGXYK6a0QXJDfZfxeg/ezqS6Yb8
hS1kyk3FoPgoRn1D/Y4eJBPK1oIA83E6i+XVGK9DwQwJM7F+koTl13qULa8hpQud
EQcYXfQcUupBICtYsYoc+Voch9PzZdSZyGoUkjxShrynHpr2ktUybUUbx8mkPyz9
nIvvtJ6X3dFfQ3ktsfT/8qvEeix0eV11eW3r720Hrns7OrLMIEvh4Pys52Hdxtcd
HM+BDaoIK7BKBhTXAB8wCrdAiXZviJ5Dv8mmDxj+XIAYx4nIx7SoHSWDRJuVPEXr
wa+V9ibOCcm+toFi/ERfCvh1MDjalIHVqV3B75EvPkqIPMeeykzoWRZptSGUaZTQ
Tm/36AihRqTtXzygukbzlDjnoFVtZU0ZRBwVsArSzfbxtQS0rlLlCTBS2H6Xka43
i7aLH5U/uiFPYyDfnv7HsVUwlLOcOzA9TFfLUXZhJrtggaPJci2DCCk8hB8VuW+Q
37C6pJaHkhhorXY6xUGs71Mn/v5XfGeVy1bhP4OYpHwxE5lgiJgeyn23EJlgZEFa
eKzIuzalWEaFEIRISb1Q+aOaqeXGKW4LJCS4Ox+aAsJmYNWoGYe+cWDFW1wh9G1L
4ucdEwWUMAd5/pxJB7dPWBgLZU76ktfB0Ua41to/M/oeivRf4d+2ZXWLAGsS5JSO
TYD3os6eZcxgGd8HKD+VnzsugKZINIgzGiRvoFh+iwMPVh1rzfW/HTNZbwPdkWv/
cz8InX/REb8RbjsuVukkBP4CF1rHYQ/hoviRGBDoo1us8OhqCjcxJulFmOybjbqa
3bGjE7lDbl9e60D8wHFEbVp/KR2oOyO33kpDYD/SEWwHGzdjGzWhMZZENEcJPq6e
zvqt9oAfQcUpAGztCDuhj0Epf33mDiuEN9hHuTS2Yh4EQaau9POiDeSKHt9iYNss
fXAZNzezjeEiSA3T6umonzwZD5iQKqmSmrmpW9F7FJDH3siYLBW5hqez6JwQFcNY
7YpAbO6BPXxQJO1j91kqcV1AlpGG17aPdAtdGNOuwPBAMHMm5kBRo5phy25z6D4E
N4uP/nZns3sdsY5NvPeHpdtJ2VLPlyjO2GVewk28frDLrXW07NaS/DqRFfHQxuPn
q3KkmOx711JgjPnMawwbO3lhD6jB56J8A1PSnJPfaL2uCFRoTAbxv4XGvNrAHEaq
AbVsIPqo1EI5vKPdWU7lYOUqGhb6yDajRdGXF1QOyBZrV5eGBKJM+FYOasrpBK9n
sMsjSRrNKa6m7FKJgdi6bh1QQst63IeqMULe3thf/1C8uAsVD1YwvriSMUjhSNmM
yLKvr9BVtKdnQVhFgqaDHkpJSLiuRuS2A703VK8YfWvd6Lku0Mk9NY5WprRbr9sh
xs8GCY1468xtVZiWiZeZ33FKNPHxtcywl6zBx1FSHxi18+LoehexSQJKkRyM5B5O
AR/AzyW6OBlM5dawPYxIcWF/ZKDmYUgPedEILNjSNknawKs6Oq7ep7j5ZfDiUav7
leKF0zpq6EUDobrpRMNfT1gWt9eW3w1iNm5JOHmpqnvLcnnzQ70I+ijn0fEoJNu9
cHANB3mhecIPhqMp0i9hlXNl8IH29QX3+uMl+fy/9VDQO2lh/VrtGa64sQXTvVy3
W5S4GFn9UrCGhGmBNBa33v1KP975equlF2Tmsxjq5Gubg8sJN2n1SFGWPqeN/9Ws
DpO0k0waVjRPYo2PhMmpTO6Gs+/P7c7AmTao5Eff5J/aVUEd+5Caf0rO8S+5TMd8
QRAFzWGlhmcD3zW15nyF3Hcp+Vrr73f47nv6XdL1gFYYouVoI/S9u9gSYTImhYIQ
obcKZjoeXsqwyyoJX9L3rCADGRrZ4BYZKln7zpSMfQB+hLrOi72lNoMqhk8EAtTJ
D4O475FwThzc7IFKA2rHoDNcBNT1t0fUT2t8jzuZhauQgnVf5h5pY0pSdGRQp7Y0
LX/pkxhsjGwQiCAx5aqXhRkTg63LU2MFJKr8MInPEURaixe+XxjTRXt8wawQR7P7
CkhdQedF3GDE5/kDWeB8y41FAobiNKUKCdZf0yV6ULBmmbtbJTomaHFOu4HjX1B9
Zywi4KntzsCVkq1I25ek43tHUebGEFN7ry9c/ZQRE5KCwY6oNu9W67balkLbFX/U
TCdumd8O1sCY7uAfls+1Q6KuLJ7ReQYK2YQAcQZy9GKLNpx1PUADqF6zB0OGe2jV
IsBX3zyERv37VhNppHXrVo+3IVVCUuD0mWBHmLFW0YjjoOPdfNR96+xVcmdIRTIq
uq+3KNIP5WZBbp20ws6vHTAkrIhgjsyV/z5jsN6TQuBL9hs8/rvfLAUkeDneFYHg
4fXwsCkMaS0bvBkCVTZnDHRxUP4PjpWcu5XlbpcdYMFpyANa8EFnYsgflwJvZf3X
sxh3cOCXQa1oGnMuAUd+PwG0oGISJp8M7S80YKRGtohepUz0Bv7C4/Fd5LBu7swI
V5T8ltDP7GFXqDTY8Fk/NX8Vt/4t2mY6blkJe+2lomukx+MZMIdeeCN9e19ZJ87j
mEIHe8Jgc9sbmfmG+kxFLzvDf+M7ed7UUjzZey7GeglpJeOdlnlAPgsrPW6jBH5y
zJpJeHpKOb103YxzooliFzTbEAUxmTyu8CTbvuPGtytY5N6nqkZYxfxDxFi5g0xR
gEGI/t814xrlhzhn4+k/eeD+SunSgOBrJLAyd2Ecka2h2mABZ2C83iqZqhM3LUzQ
o1sz18eL7+tdpA/Jg/YHsKpNHMEL6tAgAU205fHwmFPmIqwnk6p5zRCU7n8AyeS+
4n6hR3ujQK+5GBloTbeGRrirouqnukorcF3Ge4ESJiDG+lxcQH9lArdfd/OrCFl0
3tsVxCu3lX1JfQpywonBn+0Tv0h0EZqssALIQUT6iWb/VihAu/gYUpK/AcRASHfB
2Wa0Pnrd6x5L0TYEeHcjdL3pxBU8sol3tyXn8jjwR7fPy6u3SjgZ568vWWO9RgBH
Lb6V3y4lalUiMmrccYkkJWQP0iZ+dOu6XqJEhf0xRIAhFb6B2q+ptDYmQSOwHqxp
oEaBclNjJhRGoS4Ck6fQi5VdiBAX5lOlQek0Bg7Iai4EO/JzX8YxX6H+KVS5iK9y
MpHWu1Cl2AclNP2mFPCgUiK4e05Vd+YGBl6tyDiVrHwQ/WumuskeZODqiYqS0j5h
33UDDahIm/mcy1beVrGpAIfkzkFMgcCVRrAdE8idb5F3M9VH1U2BDokO/NOc/ZYB
K3PCssVAWQP4vTDbWkn1qV2g6N7n57gAvumyhwSfhNhCtK/cfid2XsmiPgpqKRJH
uGhfP4DfWfC/+xgOJ81GEADI/MI3xDp7YH/8fMP65YIhmQzz4I3mlUeklGU570so
yPkBcgeLFQ+mNQfBfEKX5wB2LVRRw0ddzzpyU6365KR2XPHQBijavw158PlHkRlw
ZlqDECH8/bwd13a9W9cOYwt28vye44N6OlAVUiPg5eFSrDNssVkeIcoIiTKs9Ry3
8iN/8cEiTQ2YiBqoFC6BKlCSHJ5dDqwDNiGjpU+p0feZfblgt/FlyPrxlBaerS0P
Oq9+d3VluAPvam8bGd8aIeXDoS1i6i8bOOozT1ZFqkDBxBicniUN+ZRACjUovzR9
ZqwmDbq2WZehPVhV9nW+XeJk8QmWovytfpsC5CVQV1vBKn+HW/0tx8DnOIdL0zZp
eflVkJDRhytjbJBpxA3f+UTBqV9EUcx+Y9xW0n1KytgOCH+YJvcjEr7/kEdILy1S
qS1QLQHQyXOpT8AIeSbYHidf1pABVlwvcAsyEXhoak6kGHX0UOoIGIUirmAoXlCS
nDl7mERLUovTr4iwTE7aigWwJ73qoktmCV0iDoNk0TA2eLDuxpLP37lkX5Qj8h8T
EpC09SYvdSQaWoBKDYSQc/YsPmkXn0jJ/AmjH8lGauAoUD9m/auM++w7vm4hnTG/
mqYiebIDv/DS/+R5qU3g1chKg3U1AWoJXN2/VLRuHbJSbMVg3uVqpeojTHb6NFHS
MyCD+qmNWyIiRXLMBFEEoK0j4LkuHfrO0pXTm2GTsRpbNnZ/6UcaFZAssVnGgg1g
I+mfN0WJO6rmsymIMVlszgQeSFF7VDIwZ5P7akNheggwKhICaC0U0ZQuJaj7UrxV
47mc5wpp1NRcjctglS8qXEKusa1DinfhOSXYzFSy4iTecRa8s9YU9YU+DFQmH94A
9xR9Qm9gaa95fjfnPVRNr6vZO4HwOr2T2pwhYeLf7E0uztvyBr80p9DtctEtLAEJ
kPz/oMqPPOr681YVCK2RvLt2WpVoz6IZQjmnKbLdagxv26Xda/omc7PttvdZF0YJ
N4YBrjQVMGitnDdwkTkLzzJCTjeJmr6tkhGkUrVjYf8=
`protect END_PROTECTED
