`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaAOP+VuIgP2FURMb+1KeGza+usIbB61lPtvp1UDLOdbhSkj0mihV/49LUFSvJrp
TdUP7eieVjpINdwKsTWI8tIT43gwbaE1WUu/dkm/eNEvFe2hV3FBEFJLbl4ffjwk
ColOjyX/t5Vh39KCO6OIvW22VQ/BlsmkwgkBIcRPeiZK8/NWJyD+z8wxZxbyJzN9
mFXRfi8rqz0rF3qYntzw114OHvelXIQDEzpgr6ho4+M3KSASk5s27Jk9OUBtmu2r
15fHCuDPDn04JcjnUyAeGZxGlNXSNLM1jtPYnpo0lwSxNndl08UfCev789oq/UlF
sJ90tMgRJxdAwTccJuzWxrXCT76c+LPbQXzBynkOky1DZXTN3RbNb+2Si2Bcfne+
`protect END_PROTECTED
