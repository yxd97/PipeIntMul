`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vv0NwgeLBYOUU2LtQ+sSG/2uNBC8Z6fUQf+rOXXQ1qapUQvsFHyAVgokTud4vK4L
UPZPgtCeBi1G/Ae5XV1+PN08ArlvcjUm/5sMfQJYDOy/rEjsVl4VMyWjxBaMr3gA
1FcMn/t3OI4LKigwZBKl66lVBP4th3wWQSPwTg6VLtjkyirwZLJFn/z660Yzdwn/
aoWS9K4frXSLnx3KmSvXI8FF+qjJPW5Uyrpg/YqMiNoUazFNKvdbxdOz2Lg+PnkO
r8iRCTvO9sCW4NvosL53C74+U5G6IdolLPQ9B8bN2X9kUx34IqVTlnsm0Sn8ph4U
eGgiTs+h9xpDaE3mTSspXp1cbPWVdCjF+xNtVQyO10g6YEtdaREmbAgMg+vBCr9E
7cj+UDzoU3F1XJCIFwC1L5lwT8euuRgKflRhGLfOOwYLZ08HyBarhSYLAhaUM4e+
nex8zVQEnnn0kWMfK00dVo8gDryCMt+SIeckmwPNYhhC/3zasb4t3bd3d7ey09Vd
1JrWU1p/Woa3J7lyWUuDcvcAhhg/BUk+HUwjc3Ws1SnP8GHvVTnK1zKjp4EqP8hN
codiGFHNTEIAjNK8hyPG2V3WCdInBwmizVQyS5d+sIQkPCPSvnHwN7uHSY5hKcny
BryV/96kEE0WzqAnrHXhMo/ctWMfSXm4bKm+QE/iKec=
`protect END_PROTECTED
