`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ncv/5xrMxwp8xVm8FQ+aA0nbofCkI0KzURpDeZb9iK9DS07Zctc5qPMGdnucYVLs
LpcJRjx8T2qBSXQ98Znzz+3pDSGOy7OFr/244P9AO3cngLlh56DVHfZX4WquGpLa
gQYJfiFy6AEtHPuxQqs8XubWTHuY2O2dywB3axrL88kdK/OxY/R2XJRlsaz94Vbu
AeKimGp/mrMdi9B9evKA2F7yvR48OO8odZrgVMZhGpzy5Nv2xiLS1ltIkCmA/nQC
xWbfyRo3unLQA13kOjToyONPJiJjgS0yMj2ta+av8jJ3upRgZc1PGXMT0wEhXI4X
c5e9SbESA+5fdIx/qZwYPYFK+7bnA+KQzXp6QN4w9wWU52Ng97OJ9pCwlgyrXkzQ
6tkbtzVvPZ8+IZECbNsbKikKagBKfKmb3HO4K4EKHIOPb4rICiI2NTEWQ1NH25se
AUavT/oRIF9DyTO5QQT11gMeA/XiG92TxeNwdtn0XAzBoNEB12WsMO6BkJDbx8sn
44K3pypdDfSr3++Em4QaoDVxyTJKzm7pRrys2FhuBznEkYFAGkQC8xbx9TwagsO6
ayHeMP7AwsBygNJmTS5QqqeslQjTccfBUr0XmZSz1m6Be++2bHUkNiIR2VipbmXQ
MUQf5+4O82vh8V7IiD51Zs19iD49dQ2Ui4DzDZlO8h0w5gOGTa/UcpkzCotibmU0
Kl7nDnuhZaVviXwxyUsfEdepwUuF2W+ql3IY0nNEgJWVb/hcqrcZTaDThTwixywV
xTt4xNe22HLWBRftY7Xu80R8lLr0LP/Lx1k5PV9XJnXDYmJ07f+dRe9zwuFQw24u
9dnMx0CQhCvb8KZ+5yUWtCcx/4zTw8S4B9LUfJpdmjZG312uXJCX8KoM0AJ5P1WJ
7SY3JJkOgQc+QHNf8yKFegrChYYW2kSmnc3d40d3uzw=
`protect END_PROTECTED
