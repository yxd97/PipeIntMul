`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7OeAdUWy4C72jZ1YJ9PxgZA5/HtCRn7+hr10sdI9J0otLx63+rw2t9X8czNr8jlF
u4WopBdRmbrbBZkGx3NhoVTYH10EWmM4PKFuvht7yDpYHxAclIFOhiTM68abTSrB
8ovfAmdlXynvcSXDmLTvrAu8N+qJXQfkfDkwxJ5tqETvsXjVfhspVqaDW6dNi9Bs
rpQq3zJFfS+1STI4hCQn5taNWiKHPIaU2fvedThBUvdG/lz3XHwL/YRYBTfHBQRd
ex+q/2JUpFVHsZiSqiT/5hAHeuO4bdGj0H+7Yf31MPlq80UjfY9dEHLvra9JZsVS
VphGRh7ahW5f32pP+3iPNpPXyzzxEsEhjjy6IX2VwZPHDIvUKm6/got3P0I7Z8Ne
7LulkPS79E6Z/4h41RJ+ufNU3O4NtpSPiA5adQYC6gWWKYuka4AbYAT7e4V5tAAY
2nM3GqgxceMRfSGAd1R69zJSMO6lfbHegBr8AfAk0aDAL90lFXbM+6UXgsxzK4JQ
56+4UDQoDpNcDHzS2Cz+AhajzT+3QGTGCI6MC16DsdoFvjLxbOa3afv0GHS8S/2u
Ekq9K/2PBz43sgtuXqEFAPDpsRhCfoNhYdsK8tUb2sze8GkCjHMctHifhuD+4H/S
jFVYIVzlWrKZMd7Cj5Y2MCMlkB9cUpAUOYbi494rCBp2dewXd1Dmz1HV1jy6I+QJ
3TB9r080HLJbqINU2uYbxmz2/Xs8AMr4rj8xOiCVzGY11I9ygTo1eFwADfsmF8jE
deI9OCi3LIrQRmrI45u+6uN7Xtj9rl5ToqJzIWc25Re3pGo0mSZi47SwZ4FrqpkZ
LPB5lhXWHBgFQGx3kJF2/0oSSQVFRUFj6ZyxC3oC8wUcgh3yCad5zBrPwqnevwJj
qwkQD2EQrY9aGSmDGXEnUn6koFCUy2BhpPEfvlVc0ssFSSX6gZ2BGSkmS4mGBcow
3MUSHypY3LhVflOkNlNtEQPGulwaH8euzHK0a2mtmrayQA/w2yV7dqmlvWtFSo7b
Xhj1rMuKUlC9Da+Wsfpf3V5yjy+DVnhQkI4BN5LVihUb6Tj1wvVupDDeyxiN+WcG
I69O42YPYUoLfCThiVkj1W4sVWEMBT3jJAB0VJrr2jeyAU4jQvyqkj3Y0heV2VYb
AxbdCTD2eN7kjN7Xue3vRVaSNhbL+p5MVVg9d7fiS7vDWcnKwHWC/a9sfFlp5w8p
cQYUk4pzhNT2rEAt1YYOZlvXdsysepQzNdm5PQtjrPXGYev9eMSk+3ZeW9dJXn8+
SZw+qHRHUk4++UvBym0YQ1btPIIFXLcovVge1TFVd3J1bZcLdGxx8jNSFKimLBWT
tnvFTnO43GBwXDgeQAIcfRRDuoPguVY/efam+nBVjIXek+eswRNEeNEx0I+uQy+i
jdByje9nx8s1DlUGJSx8hNQ38xPE0SOLrSzBfe0ET1OaVE9+m735CSMd9XfcgHyT
Y86xDjojFGMOval0qGTcoc7FdFHbZ+IZIJOth8qfUqxAZag1seL61CPPCPXtE86y
M/RzSapqo7hzrM9loa9foWCgVdIq4bqS/pBiqUS1VcGhj8zxwUGXGDSBmr/Z+8BR
qGb4dhjlbw68blygFiRPVyf6O5O033FQ7eD956/fzTM0bGCjr0IQAlHKywpkxnB2
0m7+MC5yxwWZszFMCbZN6cumAX9h6ul5rztqNR/jvfcMxDDgy8eL3GNVZI5sDni3
q2Re2uCizRQlCU59VkMmeu48zKZSa7BDmTR/lk7d05vHtluifyvTY0s/dGSK8V78
NnMLVm0r0PUV6QpWKeddWBxN/ol8uLnhGBCEoFTAxSmdfvaCTjFJ4n7a/8d+HQi9
taBl5ge83MZdahLy/Tdzv8Y0HTon17gRyndjNWp2vdTbR8R7HsmM1wwuAMTmJswn
8I2PJT50sNi4PviRapo9J55CG+NbVlfsF9sSleYkWb55OYVyVcQ1ZGQJhbCdfoo4
eS72nuaQC4XhOac6rZ0mHJNjwcJLYyvSxZAFC8Tym8Wcp87E/tBvbWIOaqayJVw4
krnvACCBe1+CaUoyjvu0HMeQGgBxJiiUKt0TjWiOFGEdmWjqDbCk6SKpmynvHXaz
05j2pgJjsqwE9zXQO84UeKf5cPS+nJggJ+lDo9VPT6QiG0cICN3IxgFNj/xdWFru
LQgdSD57t+E4+4r8bkFyq32hmVClC27F0BAJ7S2ACGEmwTlsAVlZYRguajldzwDu
2LgOJCINrKDoy/iTYVzbpmyE0sAWbqJ9m1aWviC++u4ZrpsDCyPFt8IgaZssx7Bh
WxPHsCPJtW3BJs9v+lDiA5eCPEtkoinOo7m/prcIKfORwroq+XbnwxjpdsLkWYVY
wq6OBXoKMSjszk8iC66srnfZhFiHj6Gv4PPZOIAEsH45hsihmpo8Q6wf1YBEVWzD
D2qPHu9MiuYxFOxJ4JBZachkqxGSXQ0CsYwYgjchMxzuBXvG8SdAF43dro3oswPM
RBV9QGtHkbNWCbiBeOn1w5JGLS0DHUxAx+mczoMoTDww8fmE5wZXpH5xz88NGyH/
JqfHQXXTSvjbtlFwG4GZtpbiOyWjQe9YmPjdIIbqTr+u6MA82ZqqCGnmo+qcDQQb
5gjDbGy4r88AZVq+bops+RC9Tth1/fLRmTGGYW7EVg1+f5DSQvi4xctVycoMEvzG
ENSbhc8Z7uAeELJv5DZ59GRNqhPJdgVW7QiWLTE58qazrE8fQTFdYqUlPQ/RRUw+
i151Znq5+SeGviWxvm/NfFFDMhlV0xHlL3sasJGvJ2aTEwD4Pf0WV3dZ5EEdYLkv
+sGFWF+NO2EI9PqrMuD2e0VtqK3zHseHuu7j1apgzB7AR55GUaCpaDCNQp8tHO9z
2XMF4vBKSU0Wu+ZoJd+0Lj9+pCvMqxT79/UwlLK4JW6XorL3xnRsI3cukg8r05B1
`protect END_PROTECTED
