`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IaG3vpYKYUtzNJjjedKPXrTTeyxrDEZPOr9oqPBMWcs9gdTYPOEDuQJxY9EPhRJI
z2UkSIY4gU+mO+htVV1oUH633KmcGyAz6DGBs0+dPcutwT3aI87QFdWh6p/5CtNz
gvTtCukPTtYklCIlOXDChTmg18XRiw20n6UF737V12Hpf8Ls0tlAKuvzwFiALhlN
cwYlbuBuaT2lkPxZENBqRTijW+FYDnmTwAk2UFzU/uNG23nUkE9+g+r965Ssj2v5
hzpcs4XDBCTWyGI+njOD+FgHwjftQDLuUEXW2GiQ7cntjAOLyGbeJirEC0QUuEJ+
P1jRRzCrYAB+wkxxE33Yh64HPvCeQSjz/cRZbsEru8WZB4pUz+S/5Wsw11doYtGl
fTl9IfGHehtllZKSHyLEoIqfhCT9INotcTYxGe8oUEXgCwmGsbG/VHQgqJ+ZCRTJ
r/zXNnEUtI94fPtiRdar2xT+S96zOo7yV9+jEaMeHumL0kQOSjwT+/+d5CZVdMW+
SngEh3MNkzr0GjN/00FlNHnNvTdrHerRphl8sMgZi3ANIXhafmX0UBHvDoKey9cR
khmrml7Y8tckCGMt2hpqusfM81lab6U6bxZmNz7MGEEAa4CefDDKEmvHlSseKYPf
0tEWjuucDPpMecqLKSttd8qvE3qTD882iXMcTLu+SHD9R2325vDjidc70XGWzjow
fl0LWRKnFxovmKNfniazLA==
`protect END_PROTECTED
