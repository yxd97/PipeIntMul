`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYanZG4ozxIRhRBYIAgiM3v6G4TweZDQwl7gHtzayZkr7ImRO/UpvI3Jcjwt/Luu
7f/VVLBhmXF/m4ZW6uCjk6e+C/KR84web9CI/mnRKOZ5dpTJcqRYkSrWtHTQIQ+o
kll0zCDOCJJ+0817hSuzWCyTqoyf7o6jfNMF3vCnYAm709Vo3W11WTCy5LV5cJCk
MhpL7XH57jxIZ/bfRd/0olpI7TnzgR21L+YQwJ4+xyrVIZOFR0NPtcVMSRrI0XMq
qiBqAtUHyQNqZrFq5ph9kj4nP38do6Fvj0uEPwbuBkJ+pgX61LCQdOIvd+eDG8Ky
b4qkn5CL7xQ84GTIFlT770B7qtMJ5CmtosAuu6dZ4xO0NlNBX9AS5WUn2so1l4UL
m/sZHLrnAgV+wqWRU9FVPPig/o81HpeAoO/+Il/n36eWzLIGfxenHMksqHzubTEu
J728SbBnFhplZ24ku4zZ3tFtnXXLyCwHOV+j+C5Ucn3O2OgwMhuopn8zxRIuHmY4
f6TlQI4+WWWfGjpxovrnyNPUsO9JxfLyezlVuPr+72gY8BdV0EOCpz1tZZwAMw5a
NQAKAnzYiEvURZJYmvH896M6M8Z2zEHkOechhDJuXsuWjwMA/S2Kbt7GWYBaXqpl
mATvKf+qUkP8gbwasvbZxOvWdii1/x7Opubb6TnBNtL+enM3ip4cuSceRh0Aex33
ZUFXLWqqvEkQGZK3U/U6BhNDtkAM31DFlIwLkt6khak+IMUilzvGNVokq1eD6biT
R7o1+6baHMXsjaTjQ6LSgJzQJX95MtLgsHoJA/IAHUgT8mCQIEnQ1kzh3P+BRYN4
nwoSR001b0aONsTfgQJKRlJg6zqvulr9FkQxl9CvPTqhDSZk/AWmmUUE4lMdOSFH
yRmwgr8egQcKEd187dETf2YUR5e4Oavh/Wj6xxz7TS5IZyxukO7sYcxf8jfoF76k
Xf89SnmgyqDeIhxutiA1Y4yvYR/84cs+SKJ7zBHqqN3tJ38ZdPD6wXrY/whv2EIl
8QLo5soi45MSIUpLhyah6SJtYCDT2x/RFBbq7qg210ag0VwJXG54HLbwzbHL04K1
8JaPB0v3yEJPnlV0vycYxxLGRgbGwv/nGMr/tt9Dv7nri/3x+zuO0yumacyfrK8t
IJmne312XYyf4LTVFZt6zytklql3g6cj2SuxX6wS2hikuIxTE8cFMIlwi4vIJuAT
HKRufRVboamNMeQ2KZodMsUZ3RPbYKIUD16kTdWnR15unuDYVGl3+odx9qDRm0f7
if1ysRTnGv4xfDeXxGONCRiOpZnD6wymG6Vxn+B57nC79TIvejIrt4cCkkJFGXPS
7L0nHyMUzTT5tyxuuW8vTBwwRMJkYBECshsnEvDO1Vb4KyfNG2yZmSEYtC2iw4ys
G29xrKHVIUO+ETp7WN4Cx2cfhsHrjIW2xpx+2ww5yRw9q+80BOKqDzk7LYOzF1wj
`protect END_PROTECTED
