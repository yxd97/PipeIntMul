`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/B3tZjO7YrTZoHFoG3mcSeGgXdSaBa+JELIjVIhLZVRRxpOVSzIwr7qbGVpNEaoj
IK+/3PJXVRNE27TVDDkql0zq+8DcIjZhZ5u3AViBdQVLULX6KpbW8Y+43/NUCg+I
LaVRV2FYHVbbKGWZrmKpxks9r5kFsCSmhYiuYX4/ojHCGJ4vYva6OUyZNVCzNyCv
BJpTmEm1C+ToLiGH0XEuIvvpaz5meTzGfLYRbGFacoRTvnIxqVLJNfT8D67/RExP
F0E13OXkxiN7MM3nII4oHZiFGFitBjrTRSvVeiaMQ+y1IGS3HQWJrTFzFiusNNTO
v3fdHPiiCPQMigiDxkuZR/ddtNRtesU8mLxHxAGezZY4LgEGNINTtdjqc7uUeJNQ
qmD2+xXDVaSgNXs1Q/5Yu3+v/qKPKjCX+Nr4QYF8V+hWkxUwQ/MK5fu8q49kmObG
jnfvQmNV8A8SpFOuEPJERz0xBiRgG/51gl9oR/Zbdd0/2mzmDpSMvzXcWsTAYBuv
5nFygGnyLOPgYHC0E6Wn8y+Z97UjNtgZoKHqLHAFpSlsub3da0Sof55LTQgYRh6K
FXcaVYV7cgxLpz8fSZKMiLa/4Pg5avj06gFMO3Ph4R4=
`protect END_PROTECTED
