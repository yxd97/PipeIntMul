`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OB6/IVEuXF1UHytTh9PqVQH/JH0NlcNaqU6b/QZeP89rjtWZNir9t9OC89BjoeD
Qu2wUCYqG7wVCRodXWU5j088BNuv7apFJr323XZyP8J+JsshmSGdtcAg0rvjP5gz
0Rq7CHoNB3+1IT9fwbChfLXXfyj5MePaq7xslosc3AS2J+VIT2cx0thH7THB96AI
JmvDwaIlZ57BSgoHlFgDYuZ8LgWTD/ojmqVQS29n8KAu57D7ievvSOTm6/17BFNA
Nl5R7LZj1i9qYOhNXYQY3l+KP7uN1dYyrCNz1xzKm7Q=
`protect END_PROTECTED
