`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NYfFzijt8V80FkIOFeXp2lD3R3VM19bPVuvLnfnPBpXHd4hbbiMDDUWStqFDyUYA
q0aWlQnM+4CM3gC2yocl/xIMA0jykZTihRHwKvJCASKyGn58Am+Za2ZxPDjzgJgf
QnpgAYJWx7mJyoNZjfCf+TE5VJNA0TBwZ0t9NIK7jsZTyfHZB5YEgSa7yzw1lMn/
Le6pqcGFn+81JCjpYpj8tDex911d+U2qnRSnuGL1jWhqKiKt2+MQjkWf8gA/pUTI
VDJ/gztRjKXj+agnvvAH7KPag7hXVMzZ6c11OuZ2WkHwwlvFN5Bk9V21wstrq3vo
rfIZ1jpqSmy+362kovqB5UIf0JTe8dqKmczcfrNP9tK5zLHOjdZnTNOjRoQa4IZK
RM54tV50SvRRByJeV13s9FD9hBtTKir1svLDu+Y3pO8=
`protect END_PROTECTED
