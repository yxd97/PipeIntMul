`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8l7DxyEUuDPNz4M+f8oti6ld/Vlk77bFQcv1xy2S59VOy/B2tGilRDXELHK42rZT
ySodNR1iZjbyK/bA7IisUeHlVw9LtnYwAHbVq0fatpFIu3a9K4/7x+Y9mGyI83r7
Ac55YIwSX6g25jSnX4V5xPao0LmjuTjoZmgk+AqvTsE2YzEvztij/E6riD3kGsmP
UeZjfSz9dag98vRY5O4Xwycqkl+j+jCyGWTLUWvz8W+66PeHgYm7nR+suFeXiKRa
W3b0Qm9EIcTpI1eeku0xwTcgi7Y0aVE+uZ/kAfXwgO6TuOlJaH+H3/S5R1VoTnBr
F3jvxYU0cthKBH/HFt9XcNBuI+jSGita2HhekY+wNqaltHQOTuc8Exgj/brFi9x+
b58dDBUrOb7ow3VmjU3QgnOawGi84cUr8uGOBPZZD1UDxsEaS+hWGUQOROxgpBIq
VBmOMuHePy2AVBvhqMR8t3ErQEPrVdziBxJtT2Ni2lkRx1F/O5iHKDnRKNqvMZRI
DCl/udKifRJE+3ahzK7Dd8nQEnVaAkKaHNtng7GJPLICea2/kdoiROLlbISOpljn
uQWXcs7+V/zs9bG12WzgdYvIYrEPA9Brr9u1SqWyMi93dzvWRwIFYAGkc8qa9wxH
K8t328Zsvmecm4+Ydj3xSZCyIwYXvRcbW3YobnwouYVgtOoO7pADXNd7HnDoRP1H
Hsz8grhaPzgkQNyuaNYMhv7UbPXvArTlGICe+dj2U1iUSpqvZ5Qj3gy1W28EaLxd
5RcpVDzkaCokpabeoLJqbQ==
`protect END_PROTECTED
