`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6ccUiO9TgX71ljLz3Gr845+iKhnAiwjp9/DjUzYN9AHCeqROulfdbeTTWXM0zuZb
s7NufBhj4WBXWgW2rA+bWi/mB9U/aiXH8A/XxIuTEvZWIVveXfEdHsP36nQ0tMMt
O2bUYkgt0jUnHjy081aZTg89lo7FDtaT74iN4omcHpap4rwVATE9OmMvACegcFmy
Shc6rJZvGqJNxRxWcAZodeFqtZg6QQTWFY8C5Uc5YZ0auFV/G/vWiOwC+afrIv04
phPvrmPbUQpgMKbHTGnQZkl4IrMg8ci/SRbC/1Qbbv7t9GZWOH+wsH6Fkxh1Nvkg
r7yUu0F3m5iPEOqClZYbs5y4HDyGmxNGJ/44m1Ysvv1lSczGBdpMcuVknwtDCKhb
d+gI3kSPfkSAGlPZzHqoSIfA6nvxnMZ1wVqZISYdiSiHXFIY28/nF2/bxnEXILnZ
`protect END_PROTECTED
