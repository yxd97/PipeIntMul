`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VSmmbeGRVrtt/MY3HuXMx6cQkjJGp540cYHvTK0zp4fmmRLgjm2SG5UaO6aoBRZ3
Rfc/NKp6+Oxqto7G1swb1bViAqN7R8LEMskpny3n/FMRSJcB2Z4uZXzNfvtHoZWP
XYAH6DX1XUWYqsVMXQYYepWdcAMrCvy8vQrJplX0h0ed+KyV/vkQQaybbDYzDwcX
zvrrO45CIkJZn2Hh9oteznhsVpqWJaeQLvRsSczgxu8Iy+pbBAEKD5shjS6EyjVg
/MVp4OpPShPnNyQ078kiTdQmz7sZu1IFUX0ATPmEr/xMdguSmKrQX6P2AonqZeUq
0Ro/7OnNm537wzZ3Fca13FTRs7FDyXI7cBQ5PUxI/xwr3UvJ48jXsbBC0vV/u29K
DZmvUFreNBhqUeT+NYDoI7X8+HMbHOP74yvNIxILajo=
`protect END_PROTECTED
