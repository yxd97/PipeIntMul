`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tMKqeRpU5xnyoThWjLXJPFWM9VJzhVfWLZHvk+PKIBKN9VfNRx6By08Ycj4+eHD5
t39n1NcFrgllc1dVw7iq4MbkYzJXvvFExHwIcyOqQyh/OZ86fZaLW/UN6wxggufp
BdJMrIKMt4z85sf7I3Lbr0m/Q0wdSUpWDW+7XO5p9jWt4QK/C1Rr5ySfQvDG4tS1
lWEOpTEP1sQ/J1sHeIJE6TvSmhaIjgK//nQopf6HDidwuayRClGoHs0HvJwggwmx
SCqnONLexbRxpb5tACqNDdFKIFeK/uYz8mLV+cfZHrIdN8xEwlBlGHg3/vKUkp9T
Y4DDc/CR9TR5n9Pv3G+wq3iAGrs7iYHiW0nYLMzcqAaq5pefju0Y3e0AHwqgZ7ZX
zMnNsH6sZ12D+UE8lgtfS/q4VdIsBz2WrvM5L1UFtDWPmF6YnJ6HuMFPBHM7oQ2p
ISvPCfrw315/7NJs441NUxRQHUmlpbVFIwI1EmV0wuxM2qI8qIcNrICLMXV3Ysuj
P7FPz8DJNLNeiFuma3hFoNx6tOYG/zx+0E8DsJURqeXebK4sDfu/kKpIv590nOxX
k6+niAMy+AB3Z4WkgftS4PmPmbPNAtgveKZb1Jwo3pHZqyB/pIG721m0GVNJ61Jh
Mf5uz8wNstjJ1LBQ06p0mPbwnhKPB5B5hRVWdv/zk2uJiZkAl3jWQrqjg+SJo+i0
rU2orTKHD2pThL3uiQvi5HLPhMr+z8uewUQKbi1qRM2GzHpeu6X2+s3fX86Rcufy
RBKAE6Yof2ReuMuaSvZwXEZ72l0CgHiRacQ+5FF+b45o9YnVLCtDyakJmmjh8Bqo
`protect END_PROTECTED
