`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dNfo0R1gFdQ8ocPIuj376uFhV+qQCxGfeh4FcAJEDU0N3rVsvhb2ZN8hATZQd/+V
y0xp9qw0Zo3YRGUonjjclj29lkkSdahbyusdDqY2Dz4EasUhNGpTHvlgzZsHNNzs
nzkW3TvKZotjXc2cW9+2xaKPDKXk6a3386g4hZwU518ecafl6HpiR2zEAgwOmguc
XbqSVPSASkb3rsN5FPJJ7Xg56Wvl/ucPhBplAwT7cSIYUWnfTMFiwITwNt8Od0ej
NY+IenyJZWO0BfywMWQmvnRPx0jNspilvKuHCfiu4fmd4bKZEcJ3g0AQ6aE0glHP
a+IzD38tzsLEufcYV9qnYlvedqYpkjkVmhFIV6Z3tp6RYWMGsOLsRi1mduXrXG2D
V3XZNnNK/gak2w4U2TYIWCWiNazHW3qZgTcE0MDSe7ZzWC3yvyUDFYZwQkfmOpuB
uX2W61JyUExjIpgfTSkJ44yHj0rin86Sl7nLKxOUBvcwRVS0Z6o09gzrWc7Gd+5E
XWWoqa6s3LHsf3Wf1Bnatm3fIimGZG4e8FUfLUBbLV8e8jdjP/OuH6YtxEVNqQS5
lnrCgzj4TPYmMxesSbnGG65iz0BH5w1Jp3tFFWE238QgzVIXrmHEOVVy7kCG82lD
7mrLkH0HicJ+JV2JazDiaw==
`protect END_PROTECTED
