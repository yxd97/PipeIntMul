`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4+hX3ebcAy7Hh1gWJAIaf857r4DphHRlCtVCOTak2mIx/rnNgHF/zDF0P4Dr6Mg5
jSF7U1s4MUxUDFy8zcohH3RxE49XEzcenXs9RYEKV+4yGXxjseKE4NENUSw1kXky
dBGuIpGvWEpjDFHNZciOgweAetnxLD4am8odk0rbf+wtVJFx/vzhiN6iGkcvCk9r
/ForzLao12H19ECvCt07bl2NTa4CyKRsLYbT+SEwjBsoxxg3yDhaqblRTpzIHCKY
8TvVB5uiz4FF1t9odiIANOWvbDcO91SDlg3SDc0aKjc0DsN7/3IgB6xKdVs+j2dD
4oXN8Jij4BYfJDzUnFgfjTztLb/s7VKUjaRd4q6qwMfru46Uno/vVvpGzpVYUYEx
ol+gzMjuoecpw77PzFczaUCFVmbPeXcYcQ6aAHrFGes=
`protect END_PROTECTED
