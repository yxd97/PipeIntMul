`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mnj+a1/2q2UcuIxfmUijbBeDv0tmvBe+qHtLYnG89T7w30MMCv1/NMmhgH4q9esf
nrTDUOM57PChYQo096lH3jCANtTF+wpLQS83xkIGLIKkXPn+tEK/8ejPLyO7StoS
Lmo1c5hxAa7VnJG5y5oTLRT0QXt84oZ7irKe1bLk88LnhR50PKI+JYYBwfWM55fJ
nylLIErgY25gS78xk2RQPT5HmGX1rQZuXWXOUj1ka0DqEkolDPNQxRFIxQ4XEdp+
dEjwz1LV4kCbSBIKDu5iIkh/XJ/RKCRz/MfF6UAFIWXH5h0OwkHj5PssUjBtP+/Q
hwN9bv4hDNME8rd2Tl/x7QQeCIvYLouyixuRkTzry+rO698EhRY+uYa9gVMDZCNP
SF+a4Xejn4CQPYRMf3ucWlEkzgJgTQZlXSybEiNNrtqfRbNRbDezeIR+MF6Hcur+
YLaN+dzi5kpOBw8SJP5xtDxgtuj8ebcuki3eMZLQ8H3EYTmSXllgL6/5uNKWn982
SjAY56PWkbkV8GBqF1ow0p33K/nC9F9R8T7ZjgLdQUsJkCQo4Osqw2GHmbBx5aCS
PwoMDFekjbGpkHITGKYxOMcugrmmDuKiGb38gBFVu0tLgTMFcyjbC1BACO8WtBCP
GA2U8NvnN/78nwXPaHiZFhbryJh8ke9N0kFc3/1/Xr3rM9v4lkEdPOO8jIFkpSV7
T4LEJ7ba5W8H32VhN4KeqBmkP2112aLa4L+rNPQIuF4bi01GFCPSLas9WUrMLYe0
QqZpCz3O8afpUdX+ZxXcLtjahkj+0HPkxFpO5CBcgzHrwaq4bwHw5LITyoV66qCU
scrQwMR2jH0qTC8nHYB1pXnnV5otm+ByM5OLs6xCB3EBmU4bAoqPV2GfM8zYcdjO
+v2l56L1LlmZdHW6iEyrRdJlKN6r9UtTXvKOpA+JUt0rhB+rY3fQ12kt0CCliboL
vLCsOJWa5+bUKre9tdBAsYOhXeytbyY/XZeg6BscRJrWoZobIw1qJAP9bK2mK1HD
1jFJjIfBPQ9ckMO8Mr74k3AJFENh2PAJx1phLMxCbs2qtyBe1Ginnhsx75V2oPBd
9C1chf6Lji9kuJZPHAOREgBb0O/Nhlm9f3L1WgcKdmzazOWJB6xobAqFHwH3wioa
s16uMyLj20QSie2UTJXnmAGM4DMvs5Tp3DuYJVxHwZ/Dyd7G0+jrtkoUF5vxK9Z1
zv05sfUBVouHSMORplgaQVt/DUoo4WRF67e/PR0BL78=
`protect END_PROTECTED
