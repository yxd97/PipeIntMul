`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yQ4RD5N0skB6AYw0xwEZXywzWyRM2y4AFo//4v6a6+czaXMmpXvDBq0uGayJgYIV
95tbeXS45yCiVOYD/uXee30PRSzRn9BPdfFrf83jZiHkPIyzG84f9e6YLZMtjpj/
eqIT6si5jejEONgCY/XMhiCIALRN8TZxdNdYeSqXR3o6jVv7gykA/jHp35b3HJyY
zwEwNWuNWYUQ/xVDU0QxXjpjTWigG2/+yuDdJQShQC2dmvbjtPGkxEpJ+k43n8qR
OoCIPBLEsUp5NEG6dsu04g==
`protect END_PROTECTED
