`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UPO2aSPWxis7Pbuoonoe8rJltReGHnFPqH0wqUBmN0WpTiROXh07W+X1mCm9f5iG
8RIcVpfFGy2FbrsUgeaSchv2VjaW4lABJGoTcan129cOKwIhm5dLYQS7GsU2DK1V
kYUI15wo+uaWxZk+vn8xM0bOjpVriVq8QmPmof/3P3xoot0Sj0m2m8tFQbePbDj/
1UN0HxDqTQi8/BOwH3DChJMWLJFPBJuJhaKp9xssxYjX5MiGG6ZRCfm5i5M3U/Y/
o1j/cfLsnJc5QaBHFWWegfFJ+OGiHX9XYY7eoS4vyRgdQi/z8e32qvHBSRub/0dq
QbWpXA/RZt1gbI1ETpVlmnyvDr2OtcBt8XMVu46/TwAQaZqquTG8/ZSfP/Eumc5y
f1bsn1CDbwXyAOEW8ITCLdq05fVMXNAjcCH6cqzPku1tQ7lkkExMdWoGyknhQlqd
`protect END_PROTECTED
