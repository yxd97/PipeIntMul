`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucBRTpuhZW5HkdHtbBRTKyx8sTd/SC5H++SAhjy6WzO9fUVlpW7cANDBWTP6vtr8
8AMUPQ3VoGi+Usb/OE/pn7IoAghN9F9XlmwgXAQtobhWL6Rxak9xr5WJyvWyZGxQ
JbpaAZSUo0B+bpsDEjg24V32rsOrXUvQRhmsf1Yy5VBOeqlObF/XCYx9IOms9mWv
7XKalDFeoxlI95+KiOpC6UFPenPCsUwdVrb7+4jcmJnjSlhwIh6ZCe11mhoeq358
H5qOPk31/0b7QnqNQYSkKi7MH+1wvECoH4hoqH6B2nNC5v3XF+v8EVpbbX7xYOAs
di4jQFOiJJ3yAbkQB/mm8cHURlm3Z9djCCR++QdEhP0=
`protect END_PROTECTED
