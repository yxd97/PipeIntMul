`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O1OLelK3U3011T7ORnTGogapeM5yjJDyjyjcvVKIMuivEvwABSxV9gv2SGamZFbD
z4joFsD/gOSCj4xKLtvdE2Rop4jqjlzn85sw+aPIyK8q3BU9PrhoR2+CDlwUjUfV
/FpMvTufwUz/smHIBnWol/8R8tpiyr3FC5PtqrxOq93A58iR9YBeiWEotJcvdJUI
nUDJHk0F9wC4wri3DtY9T4PG4blkt9tFdaWjp29lLdAQalblMTmOGm3RI3hb8s8b
vIE6stm7A3X1pBERtDQQBQcvx7qmJglK+uA+tcWali1wpcJ/jG6At+eJKXG+qTp+
4SQ9V0rUtAHswqxCodg5tl0zitfK+BuJ10z5VGy6s+o/Ssm6hruhPJtqGyKak/Ym
DOYxsEQ9fyqnKCF6NcG8sNd48zrePru75S5Ato3i6PakxD6kniKJ8bG9OLDRXpGs
ICbMLBZY2Z83a6IrEBfzCkfMzFPdqjTaD+MT1TrkH/qaq5TGTIHwLUrYohECkTzW
AKkjUC9jDAkHbaKqt9lh3/9rbJFxsJlS6imqMUIwTqQuMNr8Gsy0o7UsVZDqM+Ol
dxUg35zZpYcMEKaYx6IaGA==
`protect END_PROTECTED
