`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GiMeplh00slqcLDHp69c+YRpH13rK2u6iAy64Mff0hF6AKZMXJntkT+L3Sc/QXyP
EpNsbQQhhfFzvnhkbdopXtrT+4Tcad+PoxQcHdNk5wAiayr5cHQ6ZozVLtrAbxoS
1p2N7B4GUQDfEzc9iKo/QP9Pb+e2OkoHtFFIUR/mcek38ArWou8Lvn+b52Ik1BIO
aCImFFlx2JHDVtd5dx++I7vSf4mAcu798iO2tpZeYHYu9drqpCelT4J0xMhowLJ4
fKM0cnNDNFzsa+VUr9mU8WbS3QO4PkrgAHQN1avImy09c/5nkOt2LXhnDP29DeCg
0W0qvJ/yr0yIm7OC8oa1M26ZeAR/hZQ6Nq8fC8M0uRibLd3Ue5PgcIuEvdxpCRZn
MVILru/3pMSH+n4X0Z4sruXCD5/CUWsmCZlzPGWPD0KDt/GP8WAdGaBJCJ7c2Zf+
oYyw09R3Ix5sbI7+8yQfPlHZkrtj0KhqHns8Qhlv0UlC0s71ntfjKNAETOTWO2KC
462V9zcbwEqwW1iEFOyBk0QHITFzSmiDMuOJkgc2o1OnMi2M5UjeVpObDQSF2l77
CRmvNlFRbz2tDsleAjuZghfKwm3apXK9okorbWkGnB/uAAy4DJ44JUd2YR0+QEep
l2HuRFTX3/LhwBlvWMgxcA==
`protect END_PROTECTED
