`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1kP7Oe6+AIrFRG/uxbRLkNv88dWCFXR1U332S+4w+0V8GV3uNUdpW1A5QQAmMXkQ
zBdYJVmMI9waKby8mSFD/u8fousZCQqlBmSFVQztDtAIGy6MHrVRFfhNbsVXj3R5
SxYdVJoOWyYrPcBsYi1PA8br1GQ+/XxeJWbYHD32lijGRJZ2arPmVdPSxpmUqYgZ
/mvRsmN8xX1upt5SruWx2GfV9DHvCpfwjbWB29kY2LrvxfoDdFDLsiZUUhpoGixn
uZgpkiStAaD0Pik1NaQpnwWQRhVwQxUt7UfYpu0LO952Yezvy+OeBblQCOctUF58
21SfaTQJfKBnADkhblQoI38r7mO9g6n4PYLj1EkASSpesY8bhmuG1FL8ED8QuZq7
Zd76TmzNUlP7wRxwmwax5je/G+qc1lhvjzn4pzjWkBA2wUG2wSrYue+WuM0DPzbT
lyfFDvWorkafDlFddRqsdr3YTR5Pg6dNZFRUH5Jw8v7te6V507ce6CyrITcjknOQ
h1xOfS/mW4VnWcS0bIipjWbBIDIJs5IKyNVzqzzsyYNmBtfBfuKC6D5NpPMa5bFO
1du3nlG1yWI+UsiiyC47KVwrtq2A7jxxFJGMylrjTmLHsge2vCFmuhaIhWkJzc9c
OSwpBr+D1fIvS6vQ7JhVMmGm1XXHGEeyTxRf/jLFe1C4GI139Q4TTrbUwQPaeso6
JSiNn3yJnwJ0tdqPfBe9MvR6JP3pO5wQGzsJc0gTTj1srgkZerUIjHFreVoFm0CA
PJmoscfsbv60yGjMK0/Viv7Tg2MQwtHQWJp3S/DbZ6ogzkoMNtNc6V1XW8HRQ9P1
L6b5LBigdn+RxWaX1RwkXqeRFKevdJvf2VSCBsFLKJp2wQzPJ8qvomtz7/FJ6bPF
Ae4efn1XhQiKmFy1muaILr82mEBRA9izk+DUvCtBLAlWiOA1an67NKES7zQIVwpg
EK5BzwjXxnWrS63p0nVOq7kkO5SrsQnZ4d7N2VnktMC5n//uz9zO9HM7bON2TER6
RESnBsdbCQ+5ysXBACbhaaJl+daGJKiqShYW3+as2ZXuhP3wxA4FA1ihr1n6ISB8
3cHnIvESUUuTkB5M1INpN99tFaFb7OkvivVjqSVjPd99DrQ5I/NvD9kve5J2cbzx
OAmzVwlzhLGDxSV1zfx/AAJfoDqMQDd6cLqu9FiJzqmkcTK8+0NR4RGfc+Ko5lgl
vEj6ewokU9rganIsYdKYhTU3+AgXVFKgWEEpmYxmQTf+3Hm4Gar3tAONxGNghU0u
DL/C37qu4q1YIERLZmztKEAZBcekRqydZBXGQHCZJyndngfhFrQdAPMqa/q5ob12
Wy5/zsUKojmFaYaFql4s4IOQEG4ZvuigPhxD/d8lHaGaE04hOrM3VTLqnJBrhd1E
2wsSOeNKwB6U8lgbeRXs64C6MRCMbCH+QPQOgeIOvbJpiInXqmadG3uZr/xoTIG+
+THX2QALVLWywR83i8ftXSyRl+crKnfgOu7dMddKKifJ1MFfKR4em4IYhLh7FIwu
w+yxaDyPeyy4E22gAoAAXi9PhJIvD5kpkzIQ/QoulqoOmP5zrGTgtpbG1CTqQIra
NAyvbzwMaay0ojLiMQetS+dg9nBfQtzv45d9w+3bsYjcum8cVpZJhvzbSQA+ITlB
mKQpQXJKo2zs5bvFtBGBivakhQ1m2lSVbhnzt/N+bZBRWynTW71GrpDXYM02Q4Pt
o5XDdIow//uXsmuurKWygqfIbE5qOmwnSDf69Bzba8GI+5OdkzIYJhdt0YXqsCk+
gBVVzCNjMR0mzSGeeegDXB4eZRQvc9t1KrvLOSeiZeIxwsNLJ9qrad4x4LDVVbEF
Zs1picR7q2aYFYpkIaTGFlEaAHhetKaenPoWgXNyNe9IcSS1cd2kTzRhLE6uIeLp
bd2KpYhHwft9Yl59V0OI/T7mqjzXlbL0yvtoDNDL67apS6UjHK978FyoPjc2dyYR
XspxFXcIGI+mFf38gJMKBYu95yg1tMnFdTHw2b53/a4=
`protect END_PROTECTED
