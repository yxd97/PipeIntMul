`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pd6Pygv/HgaibSgIHvjgxfGk1PiMIT9ogLvQvZyS8N3OWatc6G4JRDTz6fAmiYqe
5ys5gHRMQJgWAlM1HALipXtBiqgNEsxfQPXfXOEc3R1/LwjvIuKKNRKrYz34A6Do
XmXJ+zlDVfeSK4kpXcRxxK7L2vXmlYZ5qdW4j0kxkjYsfo7pIdVE1Ar2OQn29VkO
bYHKc4NF0peOvvk5gRK2sc5WJ9iLmYZr0nkdUpm/RqBzpRb7eieqRoWZcE+9xRhG
Bdi3wEkxdQf9WzaumpML9QLyCKjHGguej2VLihKvWFF8htoQwFVKcj2xlEZpTEBh
vfAu2/0c8y7GydFoFS7G1w==
`protect END_PROTECTED
