`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e8Y2WJVEgpvDhZ1QlOZE4O4P55kErXcnUXOxS2eLjxJ8DcoW7tQ5tCJk3VfV0sV1
YDmfyvJWVab1P3xnHf4uIBIg68vdN7+brbmJGP7YAVnBHohI4FFYGKQ4DzncPb3c
cvPmeqoH/4GdRz52p/Po0q3aCmpgJyevT6buq7sjnYZvG0rjfgJJ0H9Y2YwjgEY2
gStKll3gk0oOc7ZqJnHD7GjYKM2MaJo2Acw0SV9dAQ2PMp0VlUHtfTQSHOAQRV7d
ieI1lEk0El4yCLuSnWSWV+ge/U7n44FVquoWTCDyRrXIv0eGE2JRFd1rmx+H2Qof
`protect END_PROTECTED
