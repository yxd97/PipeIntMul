`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WuRbxITILHRJJKYPNw6kNxab3jmFeiSXlotIFdU0DV5pKU38WeMF7ubAEUit56uu
ob9hj32bv57wFCv8KPDZmIScka1KF1K1sf8toO7IbIedpgcqs0ZgDSPWI6kzgqlj
eORH5a7SbtQQZLwGwgoPpocLmGXlHo/3LpljSKpgInnW7PSP4Ei2axpA85ZuZ2gV
cnz+OBXbPZ9L0N8qd1xrfjsmuopYsGKb9FeYuHfnClINdMBMpfK9FGSBnMnTNp5W
XTNLtI0+eQ/uJF/QTM6z63Y+/XjdWu46ovflHGSYBsZnj1L5VPBbQtA9u1XjVxOz
XtYQGzQ8Qkyo0iNec1A92ajRBItuSYJT2Hf/54+Z8IBvzjkz5C/G98VM1apOTKey
xDRIH5uDJ5V71hVfUMqPqQ==
`protect END_PROTECTED
