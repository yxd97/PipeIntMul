`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HLHb3VaXoqNZ9e8txfTirkCdMfvTc6Hx7BhRCFNryNQqops5U7RrW8yYBsZh4LkF
0K9B9eCs8yQt8hyAZt0ALY21XbBtbbtUuvYwHMsLkOZgOD74HjykTiC9jCcgmFJv
Tjt62ZHc/nJBVK11eUWXsu+XvP8jvfp0jIlQvosKJwI/tj/+dnHjtgTB37pl6QA8
XGd+YbR2RK8ElUv3guiQmQ==
`protect END_PROTECTED
