`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUgkdzd/F/CMOuFAk27JXFGTHRyGYKZJ/PpcFoiu+RBiINMv+mLL6rbwcF4df4/h
8gQmRedIu8nlTASqSltv5nf1L3HbyOtSaQ8MWvILENBKmFYZNfAzLYFRLYbW/wHf
0HsO9itnF3tLkJrKyw7FFHK0eBIqouNNZWgLEMVZkWUP4WBHeKq/wvjzYW1L4gAB
4iPNz5bnWLHN5Emc9gk+ZuZWBYWvlCnOsC7J3WLm4kh8Umb9qdNzHtLCzHRXIMfg
BD3QrGGEUs/PpnIPN4TAMHA0Zd3/KphceFtlNGi6YYW3Sp9ZWxkfWjkwdq7mlDkn
rGN9Y0Lsirp41TZCW2P7DhpFxWj6/nI5xrHjSF5tDdUcq8ZgZOymCvQ77uimCs2y
gx95lQiDxCc8pTVAFE5YiawmK3zLz12WFK+QJwEmNNUIHePPdHlhlTTbaq2K7+2X
6kIM9O2dDC1JWNS059zpv07GDYZOoL0ytSpYtGv2bywzT0iFmgn4BPqdUB7CaVjH
lZQqlNnB8y7XAx0/YhdTUzQ3hizShSuSgzcttOLV3CUUHcPlNkjvUH4DCvhL0UAC
cOq6qGqVRUY0YxwFewIwwFjYP0ZHcTh/5ifvvsgkqYFWM6+HgG1Jq/QwJglgBJW+
fnr/y/KLXNNV+ZGXgpFJCHCA11m1DpRctIZX5mRWkG5UDjPjlM9FFV8ZlXvOiqO4
wqg54MpDyCvUCv/b+7ROQzolgXbFrvk/N/j4nd5hQsQU/V6EJPJ28y24H0J3SLqp
X+yzmjqZniC77ywgYzooymXOc2TuGpIGTMeMYCKZbn+IGareP/has9UyQlbAaBkm
7weGZXstZW5Uss4tHA/elPr25We80DKMCvnGcSw7z5PY5tiJWeKVrLuet8XncUfc
tKeU8U5KgKoPY8KlEOyDglQ0g3I1mwDrzcWfADTwELMFsNjmkVzRxkrlU6MDGzqw
KLI3foWvAgxSgycNRICIqXKfGWIYsnnAvn/CTf1ayDInw4c0OXHgzh/C+c8c/1Al
izv1dycRskW8PQBiOJvzRuJ/9IQoeynQtY/AHcviWy8bf9yOr45HokPm7PnnXd3t
c73Z2nWsIc+Eq+f4DibjDuR7lg2O8eSQLid4XCo/Zdf53Q93lfiLWLg2qIT2q0VO
6mWXbEaVXFLk6y+fcGeDu0ycspWDqoqmscYFWBQKPlSTbPstWUpFiR8Ylcsl/IZy
Z2SvUuqIo54xlhbxcjvYQsx8ygE2ACxYXL4krNr0MGQyr2TarWMq7GqI+yCLE5F0
haoD0yZ955YacdiJNT9iCEzCdfqlLavTdMqifDXu1SHpzCIOO9qYtCIJs9/koEtZ
rLU+Et8fHcHDccTUWFLU1spBbR5ZdQrIbf07Jn9+YHGMcStrB5s5RgrndEt7/dcf
IX1HT24T+uZBDgMUsvs/4X8gI2XAP0fGpA8jfSsvFrGLPsy8aUSq4zLk+/mRXPzs
8MbrGowuCMEXL/fEOYPx0gK4yFqcD5yxOctYXEWTsmVp38bpVBmTMEdJCefYZhe/
vQ4i+bvgKmH7sNS4RgSU2D6yKwjEozafluVipriC9rVmKdm4peuz1EA+oRNsdcZc
yMmShQJYuqXUm25UTc2QvHofiVv9KkOJy8F0rzO3smLQX0CpISwYBNEEo0wWOHuy
hU3vIIsRsi/yooRm/gGLi1Ci2wXQbNrzh4d/38TVE9tk50wnagLJMTJJAUhuxnFm
epSWYGFQpyjGuc/f74TVwxCNnx6GzpUNHCsKwqXktSyCaMH28ir2aUTA1vm2jJYM
vkiP/NxYT+AjyzxW4i0/jRDSC/OjbDM4uFxWcOlI4+8okIYyNO0JbUSy294LQGT6
k4xSaKjjlhIPkZJQKtiSTcWun/0t6UTt06aHL1xYOQf3rPxT7P+b8zWdTmiSonQ0
`protect END_PROTECTED
