`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5QTb9XgABoMsBHE4lI4CAsLcwWX7QQ70iHn80oPgaib7u5aFnqA6iVgYIEpimsXI
BPAf/dgJFEVLS1YPEhuBY3S6H29/+rgQUhVzMhRJ9N4vgzvedok0JwEFnoSNyA3H
1am4gdziKEmx2jUUKguOsVvLwRJF4yM4RUTxKP++5sE7FviJy2WzU0QWJR2WqD6w
RLWVUSPS9TJHx6G9KQ5DXSR0HJHOxikZ55Dg7wVOaQzAYsqeG/Vpjlm+h9mDTJXG
rboOEi8O3kFDseuq57ITm/8Z76fJkAG3fjCRwt68HjYZgT9gWd8VIK08e9mWg4HN
Lu2YWbL+hnn+3Krp7i0/UugRl0CzZKv3/7R8WmyDtCN/ShDUeXrO8w0IbStyYPRz
d/rGCKYSFGLir3Sh/BvkNCOcw91SBX7sUHtwf9hvfMEW4Om1ESXfwWN4L/3UNLQC
fgJ/V5+I7yyISNXoJ7OdY0l7TEN+H82T5SiHmkoOZB1L4eOIMkHnXOufRMm3wNT+
Zbdm4ShCLSPRJCbxD1iUw2OTwKmUKe5y8JtTGL/B5MEpYjA40VubpKuFVu3MMAFv
0RhPO4ozifB+L9xBz3swR66bxuXnXzMw3pZFc7eq9TgSUfUI0blIeYEP+85EPnTM
tEvUzrxJkazPOUxppg4Jb+yGRsUQ2ggslGd9WzAqOmbvlarDK0l7gX7Rf13r6xAX
u86wWa5wFg9PsZatrarYFGL2vlze/Qfc3zkbs9QfhKemL6X4RJpQh2qRA4RlVmSw
hX/UOUTyiLgOLtMppoMKKBxr0Arn4fa7xLa8QB9iqPjDWi51yWVroDgza58psh0c
DgoyIZP3yy4dk2gjiXreAZiGDhLUIcDwAB0vTeY8tHxMdEx3z38kFOl4IetzG0L9
QMaKa8h3OkLkcnpBEwKYi+4yDM53IYae02rAtb+CdPSZ0vedtUnJ6MgNP6jV9zSm
mkKQ0N/UAhVSC2mHW0s0pWxv+km8enbu3hOwQE98mid4ZaTvTfg3TEX1t4GLWa6P
qRlf/q/imAwgvCtACgRIiQ==
`protect END_PROTECTED
