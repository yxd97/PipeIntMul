`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QgB0tmYX50+t5iRTb8Bk+LY+6OXPT6pY5ih8sY5fs/6VfxDj3UkZn8nmS3V6lUhJ
ax7Z+jWgtjqcg3o964c8Rd04YFEt+Ph9AP23v/7qX+g3umbDVn3Sh2qqNuasUzjP
hlKSeRr5U69J2FA+dK/YkNnWIB5keuC9uGcQEMuga5w6OJPfy4sh9ZVmvgqG5AOx
Qi+zNJky7RLsj/WwWyojX1hpkdKBQh2aNFdp2S80o66m3UmnZUptsWS5EiFnCIzw
dF/gz5+YZQI91l9QQHyxt+ccYs1ZMcOJ3M+ABio9Nf0rHv0zdibiLoo418muSZnN
hmzjoIVr5w0jXDhjMYTZAuB/MvzciZuj5vvOSjf+TraJWaXxYbWSzfQYsGH35xLS
MVtq11t13eX46XVmRhL5Jq4aRaOkKAoeFRZvtObBNSY=
`protect END_PROTECTED
