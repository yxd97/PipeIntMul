`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zX0IWvtzG67VW5iV1NHLZx6neonEqqPpLGb2nU2HrTSJbZNGTYYc2lx22lEQUdw9
N6pbedqNhCQ0auAIGwhZUsH93R4sRpqNcz0jeNnmn6i/f+SRVrNvEHuY5yENur1G
bD0gto2Mqh/sztezdR2jF1nVocwe1UDIroiEkocTdMkXCXRIsuG9eStDlpIfZfzb
W5SkdEzdBwdB/dWseKQUeiCSFpuXoFI8Jil4wOmLN/pP7eLcEb96bshOgzpL/gxy
Ryd92HZOeOxlGzp1Fh8gBGVxU5kK0FpcM0f0FvYLkjq7EOVyqdAkErttzHZQqfR3
gCZXKhvNCGvTeNM8FPOw/GuwI+wKPhvAL1y+2RMxOeGVlGXLpoNmf1ALhXhNTGMh
jTgBXUnXxzK3veTHIo7O7Dex9IoPz1kWP4bufyrNDPxI3pQ1c6bK3rI6gM7nmEMc
+bjKYRZHnxHJ2YVwtdvbOWYvwjrGAThldbvTVrnZwvYZHsCvRCoXeZ9G+wWXeugq
vffyhgJBDkWxSOkL/a27Krw7Ksu9fM2FrvSmMsylFr09tga5qQWX6QclDoPp9QJv
aFX6zfuB1hcMzSfqHUwGoBWi8+jlXx6/408mJwLRpk26wRKiL75ImmkWMubVRO5H
OPbthdee4Mc2dexbzStUUsRkc7KtTgER/eZykS4ZeLSHp9sSzaxrCW1yNoay6qT/
cy7tCAuLwMQq2z96+sXeXfUll1GWS02pIzD2ZXUucpG7jKyGr8s0Wyn9zGI7T8Uj
ORvdhNhrNU0RF1dJcjaVPEx+AL5cyb98/kiWXfT/hfbTxkviGagO9yNoyDeNuOne
soZqD1ZoZGPDXy7C+jQsIVSQDKWeW6JsTcE/vxo74eo1BIm4FjuVLf1Hk8Thq6lJ
RjsJ33f4ptjvrR0h0XA5cusBsG5qkPSTL4Bt1alDYezrF1b1LZUXJBnKys6VLpBs
9q+5vJqGPUgzwFggKlFK3Qt8ZCpeGPCWQg/GERTsAd9vPw/ia/RZP44OqbGOBVJX
RiybBFVPuedbqxqbgAR1erZCqRTctiS+P/GtdsTVNhjphFk9CkbgDGy3uqBCxx6l
2DPLsXRkHHcXjT9KE3gjmHbT4s9RK7WXOq0nc/B/2S2E3e/Z27/LyJ2I/SkDbv8E
kdwgIaVaRt2yyEJIw/U8yDAQ4MKnEvEv3Ucjrylqpezu4be7rKNdCI4PfHKJr+2O
mr5GqihkgNIHtI1nlISbjLrbWXRtlH4SotZ1JK7dOA+uv5zDv81py0+0uotSM7eP
rlTi3If/k6JLB+F5Sjwf/Kmx7pvBIzhCNicAtfZIUp2XjGmFP6yz79At0HhgEAZh
+TgM4orVqFMyeYB03cHn4MXOvscUNu9/ST3gWB8pkrP6rFyxPaoMRDyUTQVT2F5M
6jjGwrU8pWbuJyzEBcvkwPdmEHJBRBB2kQQNOFRbzy2RXaPvFFrQgCdafr3JgO1z
NEDF4psJ1uuWIQa6wbB0DY360PO+Kvtux0mb8ZRbaEGW++7DRPKO5QCHTH7iLJyQ
MPK/83XenphvqoRTiRrO1Q65wStCGM1MSQ4yT+IfoVPYL2kpiG9jBsn9cQMrJ7Og
J8WERT8wfsRlv5GzPRyAmW896nYUnx4odIkqr1u6D5j2qpfaWeZtKSOmIrswcuTV
Upax6Vu9eEGOebLoJk8AK6rvcDih4BGR5ebYBZ0n+494veI7PKx+OqGDBVfXW9WF
TgqIxNwDZGPCqdP0MnjyuPHTTaWAfNThd6e/xW4I+1a1Gf3LdmQDWUELp/bPSLUS
iKAM5Qq6/ezH2w0g7GxYeGur1a10dBCzqo4AaQDLizof+Ti9R53fDfnuR6hvIJ39
TGx6AKtoJcewxFjlyP+vj88CRjB91vTYC3I7z9+oJ3vTK/wYbKJwBByhKx/s+v9N
S7uCd9uj0u3hguZ3JGS8KI3dcuuZglCbIpBfkWgxayVkGp4jW4nCmQ14mKtIY697
JuRhCLeiKHihZ04Ds8Jx/tRiDHASCwmwy+VMEyXYLB3UTyEfvM4g1WDdTEdFWhJB
lZCVvRLBJfw32EUavFML+syb+oM4amJKxyTGE2Rc8OPZbvzBr0oUlImybjQYgaUv
IpsVdy1yK9aKfgcXKlc/ZfHz92vUEGGV5eCHpUf4zOHUkW6G5YSJRcWnHNp6hOnf
V1LlaIGhkOCX48NZ+Ke+J3WWzOlS+rkIYo7yKo9fktn2F4Y+pxPCl35yBy85OcXg
9n1lmqWDWU+0WVGe3cMcMzpdbqUJMqQo2u6Zgzp9WjVbAAtjZ5ozGrkxXffrZ0M1
QARlmFfaazM8LwfAruwTIUiSBXeqkyRDjjy6Fq0Z3YcSx2Ewc9MCUO6Wk6mILt09
lrbcq1w0xwAA0HyC0DEuBYd3cbnne4RB26/JxD6O9FfBFhWd3z7xeGHKp9Kh1bXv
l/dXvaE0/mLX+bTFXwhGIMtVGbb2HrNcbBSAaNmCNkolCmpucBtjKayJNCAus7IP
3sXZaUhpvETNIcQVsL9wWNsebpGd02xGvVOJxUaSNn2AmUGifUpouhCbRKwTp007
XBXOKgOhU1cxpXVMjxX+RLokS7t07CL/yM6Sg8Hh8V36vdpd3K82TxDf+pKUbe0M
efJuu0qH7d4bieq4XvGdMHBlSRBnvpspww32DaHexsmpNtDF24eDxBqflsuOiVnK
0g9Zass8Z/EZKvmCPuf0dWRtCuybExb5KA4v61BE7TWJGPVIWIlj28YMLkypOqpE
yNIEh5UWhAjS7/mDmcJ2zPr2tXGPhF57LZIIVEDMu/tVAKMRNuflvi62POgp8WoZ
NJpI0Hba2E6iCoc+7bjzlHIBzr4BaA+4xbqLqWcqaqqdPY23YlCeUeLXOs7qIFUX
6mGnt4P7xD6Vhv1PF2fl6b5paTV0a1Bv/h7m8bqmwCXE0rXci1xSHm+pnM46qAY7
PFcG3HXD9b3WQLfqaL1d1JFDywL5GLv3d2yX6sTN2vq6ZhqarVBwkHODPbV2Xu8K
vx8hYoXfNMFawWfBfy5qAzmMEj6l7Xl0hYVU9wBKIm+UP+awZft51axP0mhxqMyO
vXu8hUcUiZCZZsNHkQ7wqu0u/Y2qUmGIEw3gjqKtKGp+YlHkkwnEInK4vEaZbliu
SvxAfCCa1V/8OyDoPTCqU6PeTKG698fVNk8k77Lp3nlSiAOy6pd9061aUD8DjI16
DedFZODhbtAF4lZOfz/RuNKpMdkYOnleV8k7w1iTMYn1P22hRrBdRWNUH/ZDUHQi
6xl6gKOSOQ6qYAyXjHR3Atskkj89SPeBJ0mPcQYDRL5eeZsIAA4tf/PPJzq9ceXK
wXTg1enUymiH33Bkn4PO6EjL4YMbWUxfWz3O4eHiwxu3e433j1StASllO62DCzb8
h1V7/EXP43WR68vb+5tVBlyVWDzUHAPuimpE+fU2WGgSkjBHnyXi/8uoUCiginGp
77PuFLNHdf4LN0/Ajw9Y7d+MhgcxaWoCfpUW4pecRxV26Y84xx+jO+EV4GSKpTwi
u8InRs3nVYtfwoQFB3eTh/RFmvda7W4boYHmeQYsqmx+vXAMIfjRa3pj59770eyR
jGHIdpXnr7wHX0158xcQZwJdtWHnshV2UMeCY/iKYNX6xDFdRdankJrZMLonVSHu
2Xi1ATLzOOOsBxPOHZB+XADMpYWHvOr+URpe6K+kaGAUttoD7skVmRATCMxAoO4D
W/vz+cHZESdc35VJjIpBzd+L1j19bNoEa/LRXyd/16oDRE2veaLc4JxigRVR8/l3
bmnkP7HzOT7lqGQ2OKm6fd3qRaVaqgYF6f09naRVeLGgqKBv2eXACKurH/dCzvzP
A7w1WEeWQ/T+83Zp+1I+NeHCF/YVwBB6YnJd84skqVnPqY2vpQvmMYFhsIlBXSqU
nKtf7feROSqUTo/GaOrnVleLDNFHqZvYOge679Zt42efPaLB/S5ylPNy2kdSNSAl
D/n9BllAWNzamIzsVF1OkA6Pun92co+BJ9xAwY38bwei5cETplLmjCNNSzesslP7
u2IsOFsmlIC7T/10V1UwLLqUBI2aa13owG8oi7H1txbl4OAk1zDMNHCXlisdUaf5
d0rvGwIrxlabE8TKpZLGLj/cko5eJCO35o5KH9Dbqpg3X6DBaa3SsFiPnlQLNVep
Olpt9NO3mc7Cqg+/ObIi9q7w+ApdElroVI3U5wDQpui59luDb6vuWoGRcU647ERL
AwRDkJkYO6tsBX7UcJwIBr4En9OePLSyvVnzEt7gZ2dZVYoFvTyHTp/OkY6ABGXV
BkiCCxgyx48YGk4NCGKMVyOW12u6Up7FECjncpL5DcKmzP8Pp2AtE+ifxBoKcsAM
FMNCuFRdRuQBke7oB+Z8OGdXq+D8O3rDlNLpzTjGbnmYye4T2xUU9tH03ZpZkao+
FGRn3xv5b0MbWxJDQoKzMKgXMPK0WPVOobNzQja/rIyr802IvcMdmBMGEs4nsD7+
y7tHY38TO8mOPuOqkF79SreK70+RH7dNlGsfEoy8tnKcbEkaXVOV07eFw1VFCyvy
CHyue3mm1NcfREEvsnuVd4Hc1paQwpGnWBMYpmsBRCDfnOLf4p/Uzs15xtH9pcrf
pPfQS+TgxCowWEQjnkt7aC/5UaKqjSH9C1d3Wqm7ooHN8SaAk0QdMPQj1ddjxPsN
BJMoE+oOeD29S53MOLXXXlCYEyEXxN3ckYv1nWlGiw/bskZHTa0wqA1kfmA9m/aE
tTEdnS55sWKMqR8MOLNFPwu1UnVGdzeoPHZgSRrROJj5c9DZjLiGy2MuDVzTVjGw
UqPYRoN1znTHN4ybsvU7kXpLTbV2WOSxYmfn9ag53JrqG4//WaS2bzh4vGrhuV3o
X+FFwqWXIFQ1vONwTQsx0fQe8/N2S2rwYXF2cp9Zk5eew1MXpWoG8dzMzjS9ZXLr
e7GB08VQsA4ns9fyInNNCVs3DTExAAHFGbdeDw/AbSiYIpjTaHDnZ/lDNMsUMgD6
8GiOYl+t2v1AUzkqaShkowu6b+Kg3Hl3bBv6uolsswQqh3F5xbR62z9ecHFyckw3
8CETSAr/h0/nw95KfWRC/MuYP5vCr2KmQM2u4bfVkQG/cGWDHt0mtDzljnyeZei9
hqBK+Az2LoDfzaRbIS76vEuTAmJET2DQqiUr6jLEcDH/W+x/1KcJGDjZ0rSMMvpb
tmQDVllDvZ27eUkkMcfFhF2kwvQkTwAm/uIIfmAAO3Zv+E6ZmzUDMcvpDkv9nKrs
Rheost6TSyqBiMQk6qckECzdoAFboxejUyyAndRiTntKcpzFqGZuraANRb4kT5Qx
Wx6zJVHb9shGJ0x5pp2BGo995k9sioAik59vm5rX1+vahMNndUsRlyaRu8wdkUg8
d7HIE7ePbRZZnr6Me4QVewD/C1hKezEDep5lUKCCBb5hvcd8EOEd93UTK3oezV3d
TlcLv+ruOZiBZvOPP602l8faL+N2bQ+4W7pNT7mM/b3JHmhmUgzoKyAdHjPQexJc
33E6kJrX1tPV8Wo0A7hN1LBj0EdXmR21TFBbhmAZoNesRy/XUt6ZpeWqSPfp1twZ
3ClhKJS7AATq5CIPbx+Ld/fhZbSHHjBps7r+fGZ+rvecd9iluVFR8qgfJJlNa27Q
P+DDk65Nn7xytgjmpciV0+ZZbjJyCiUFCUidUyOhHqACFA62m2Y+/LPizx18f5/o
elsh3ME6jIyopToP9Tk8QPtkj35xfrhz8x/J8XGOoZo24fCJZ3ru2pxoBS6AhYT5
hZmzBIeINTPErbLorTZCm7qpXSaDsLoKe5V9kAhvwsiKa6avUgeahH7Qxhoplb1w
l1kPC1DJ0IG7PLx3XSkFolliL1cLvmPCGB8uTaEztsLYCx8VrlMxhAOh9wsOXEFp
5C6Xf5Qv/NFbLFA1lHJsyXoKKEYSbDEBE5HKPgx4YAayrr4kj+7Zv3qsZpoJ8iIQ
5VyWEVfeb6qCge6IdPCITRkQ1GRkB0NzOHgJYt4MEBS6crkINtgCBXwTE4AFhWVD
6ny0zVN1htyJo6vEXcL35gNZhjVomhXImLKfc2kSdNs1a0e0+ApiEXUuZ5Q2Y3+n
hsSZTEkflo4qg2uahwbo8qoxBRujK7dl4qOBH85p6sfj+zkgoR/QLy0rYD+swC2d
n6eChw5o3XkQPYBl1cbGsmYLG6s3rUGzkoDh0UxW2G0pQbTRKCuUStRLCXMZ4OVy
obRhH14Xf0QMXAFBIzb+Utol5KRzYWVT7cGKRFsK24P9Nze/g7PvXtQBwCJXPtXH
jYY6d72WrEiL4K+f6GGBiA==
`protect END_PROTECTED
