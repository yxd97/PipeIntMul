`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yeP0NrKSbAWFGu9C0pefPLHI6yXC5T8x8b/HTuxShv2jASTPpcvAYc5HYGR0iYSq
ptKn89bG+fNeikvVAfUQpkFwkCsAzonoAgDiyCYGw8w+hWJJYuxmd5Na/DLTHh2L
q87Efdbv0TtWCIolgsItysWu5cUs7gLsrAs8zdnkAVIO/sAF2HbQB0OOGgIDydjc
DIZcp41OC+dh5sDFjkwiQWEBbrvGlDe+TZYocxchOlMzDwa8Je/u/LJQ4cyGtO87
tV+R78VQ3tMqvp9LTHABz1S1sXVtI26pXt19fTi1eI5cdQ+63f4UulAo/WgH0SDQ
HySUsMhIxAfsuROMQQZyXjNczN70lIRL738jBxALuaqERaRdbrcLOiCLb4jZ+1gj
WuGKMYrdIJwQnyDxmZm1zg==
`protect END_PROTECTED
