`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7q5pXr0ekm/CrX1EtONEUBtRFL1+JL3HPQin6WMwA+M6tKmogOo1Mt+7pvwis7OO
OvvvOCcmSRdTpbc5tABWFfeNpFUzI9YukSr93aNX88Xy6dbnQvfbU8OL6sN+uvyL
E8erK7WMx12XR4cQrE/n5F73buYBbkAV6dqwdlcVpxtRAtMrHgwS/A/LZ4h8eXwB
vKtPIhq7frsMrrEa0NDESMhTdV3qLPt37hzETKX+fLxR9i/qaMFdX9eGpGk/RYFt
Y+7QaYlrcoSYTFpB0wmaqVnOI7DaFLhzyXBUSBEVsmheWzblj1Apy8gkjzWdrOCQ
lyltxELcL7usl2UEREJ2fx0PkqhleGgGXZ5Ep3UdrxYW+DjY065Sql67EKRVUQxh
OSLqyaS7Vtr9zL28DNz4ON+FV1PKHHSrOGLafHfK9D6qSvtqhdfIvLjd1bYLAAXv
`protect END_PROTECTED
