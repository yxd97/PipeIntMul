`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MTp+gL8+X9TpnDEb8eSogkPUWi1atfqlVQdQlF/OGaTvONq+NaB7ZqxbOpEbtGcX
lsGuGiKX/lVyo6gv0W0FWpjBydTOVggjwtnYEfaJ8jjknCzaOQRwo8EATGzq1OdB
R4BNECZ5fBtglHvah6uBXCmf8lBPPSmKal/oMw/K3Cm7a4CVdyze69CejxfCsq6c
2kInaOSSxeWZonvqMpCOQ0BGRICVK0ks7lYhE+0i9Dm38AcPo0CAG54qpc5nYOAg
b+sP6OtW2WvJuM9a1ucj66kJZP5vIV2CD8eCzYhMk2TETMLTxpV0eo+SigciFArM
SJ3sOHD26upYPmyIkjfNN6Zhv6r8wYdaYTnPGT8guuW+wfL0MbsnNAhJ3+MBL5zz
NG0Sr4Y4mThqGCEu4+2+4Wtl915/lWiq1QF+Wnuk8I3BQGxLXZDnq419LNV2TJOq
WTZ0ktmn3RfhHk/9PBkJu2ORn/KAllmHDQrJN5lPnLHPDlDs4rR3rZCTN6VRX9SO
BlRy5y3kjw9rSr4T3wT3CIFC9+kB1NqonlvT/XJ4v98hqk9Cr9ahpCAh1Ss5Tl8j
yu4d4vm2CT1MlV66cNtkmYH8gcicaXQG8pUn0QXDzLmFaJgbN00Klmv25NDOzARQ
p1T7Jo/o0xjMEL+LLz3CVhaqUrLEd0KlDGx+k5b17tlJSU+QBJczprH3G978MxHE
`protect END_PROTECTED
