`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0ebXnIcpjbfwcb1BZkD+iURN4TUgmCr7Ed42ZyvwGAdDfIy3itk7A2r8LnkDZlA
Kis+l8XcFcdSRRRpLF+p1l1/64H6QMKd5kV/6QmEcUtjxzSZhJI49nyE14euqLwX
vmkP1XUWs3H4CjNQcLWhxUw02b8FHMW+n0U51oVmJQVwlaUxQIEjSbkL2tt5RExR
r9wHMZs33sIXSjfzBWMl2LcOsXFFS9N2R/3zHFbZdO3XlE4p26u5baUWOynrBe4M
UF5Id0JB6r155yUeCZLQVb6KBgrg6/WamPgOSB2OUlklVaIerK4GBwAYYJ443ZCx
ZMNWARqwPyqp9Ty3+oZTAF7ko8hCHfOTQjY+iVrQ8Ifl+dAn3XdC62xCijUghyau
kdxhNVQeo34k7/83KOva/ChW21E5OwMg5WUhhOfoAvs2/uZlkbO0cIr12GEf8XLh
N7TnYlHNnT32t2Mcqj8FPCthOP9w6VZJ0mZKJui9tNE7f/o71tNux2bx+u5xk7yb
1UfIW02usB1jk/WRAuenGSjVcQyyneDVSu+UiOr7jbDSuXXkkX2hhB/ylRMJIAVX
VRGbkbU5nSsbd7A8jXuf7sSia3iZ0nwviZXzpqnEjYG/GsEOcoANgfr08BbPBBTE
eSjwg2CcQ9rjIjWMe4rrFRZyPto7dt24xBEhsVQneOo6t/df89aYmXTgYEg9hZqW
N9tF8K127PbDORiTcO6yuAp6q3s7PLukLvX8BzVeUVgbB0gAY9Sbm6Zk2gWeFCqi
fnDAdlpIWmT6CxJKSuBwsWO5/dYmwEaaqJMW8VunUVZ+sYBeVLDAVHSUdg6T6qOW
aksOWmuV/g03v+EwjOUiVg==
`protect END_PROTECTED
