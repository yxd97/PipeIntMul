`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5m5rGHW4UA4o8U2vnhH8yaws6WqXE0ezM7fw3ZVtlAjH2MwHf4qRV4X5ctrPx9C8
3TdgAbot+nXmuwzsvOgeIB8o8wYmFDRDM8ipB37WEfZW1+nPgiQk6TG2LRpEri1Z
s7545giAGwrGtajwU3rJG/k/x9vIecBKyuBJni7hg3bXO0u/tki5WMhLzMO9RGCI
2XpawhYBQvBZuZoKN6OYD71p8CYgWhJha0rnKq6dGfBDOSwVxqkS+i923WKtv2Ye
JrlGJHyidAUyYxD4cVgxAQp1E68lHRXJLiOxxNReMr7dtsHTJNM0VSd0lS9WStWK
Xa9mLhFTqtfgv2IAUbJw/C3+cV2qKTQ6kqB6hcLfkbJDjh7dUjUzWHDYLeB8uZBp
`protect END_PROTECTED
