`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+eW93UNVUb0qKOri6V7dHC73Lklotibo+Hmqwe9zFcVFbPgYdUMRsKAcF40WaEp
T0YYd+XxoQZnXGYtPRahlW1js+FwEzdtHwAWbT/wpCcS6HJsz7/lvNxG/XMBqd4t
dyu3CSigf2vSwGc3VeuwBAWy9M/SLAZjy8kKev7FCjcbu8tpSMboi6jRiSU+U34e
G9khY3n5A7pKuv6wlkEv7TwO1oWiutWNw9y1k7ACgfm07nKwYSnhf8gNJk5wSt3c
qeAKHSbZrb/+AAyE03pSkh4ZqRdPIsDMuO3aU9UZSx/G6dmNKreKMs6kf1M7a/qw
gJTo0mByJ2BZgiQqprVK1llpOzdhobTvnVJv4HNTnvsxS3UXe3UeRr3Tvi82QiWO
aCP0UWc4JpuCfuBx5HXkiiWvvnvKwzi6IgY5Hd9rgpX1KhHBk1qVD5JtkxGffCT5
6ZiyytAC1sHjP/DjX80lkGLVjjcFXuuj6eo++Q3qiY5lZgfKZgjuBKxWsFnrt1lu
iRpKds+TVwhSlBa0btvE8xi6JLwQmHJ0yPG91ybic2ZuabUZaXRL2bU5G7S66AOO
BCgKkoOlewLVfYyenyotGVgBqgX8aHRRri2vxikxbV/XPn1mkjT+i6/3KsanrxdE
14aK5zMK/uJvokyvnrKNs/KGfY3AiZPGGCjq8uIx6i0sNbm3NqL1SMeo3FQbtC+J
kiTim/DEr0N+u5k5ymRWSPJHpaB5r7gpMyhjLum4eQQyjIFTcOS3x6BPcu4VJKcS
3tj2MXYLTxaB8uMP2LVjaCB4EB70V84lDWng8w3HURmR30hA239ytfnV9SeosTNJ
Oi6VrFdzk7qaJJiEoDuFMsqbA5sVaOE/ULgMAkmphM2fPmlwe6HLGbyINfRl7GGz
BHxkLlv26u/xLkeGqMlxofQghdluI6avuIghXDwMD7p7uKVdiccNbV3LBj1qEPEG
SX/NmG3TqQA6KkZv4Xxl3sR4dIHJNVjBqheEugAwkCGDhHJdi2VYmXQlqkh5Nfdc
k0Z0VgdaKmniBQkbvUsDTJfhpsOWj0YV5sT9KJaAm0HKhLFFF8d1iL3qNt1XxlUx
L7GgaU+nMbgs1u/lkfm4wh4bTlmIx5HI/cdFjriT/LE0pwnYcZyn5526NlmemJyu
E+cHsNCyRPVUWJmFBgHqTnYt44ma0eo0S5yL9vtfvuc8K8lqxUw2EmFnJSqoxQVV
17niCQKpcb81fhbNjnTf47lvwDw4Q/lUUX5Z8QvTaeOhR8eu35OgUi5/tBeTVxzz
VahF6GyMUVr6q8cOKuADMROhnWQOGloO4QThVWBvC44Nl7t1pCSoMCN6wsqY9r+Y
T9a2ZNEE0jmojph8Yz/6I8Weyl7bw1T78wFyfHTukj9sX0mkxXGiloQjs89OolF3
mKhncBMYVw14XbwiCjt9CC7Yf2lb71iS3ZgXh45Rb9xQob7NcTv5A3Bt/eskfknT
UbvwMS7ptZPvuqC69uHtpvmK8nUSMDWVVzsXTFsIa5qj64ci++ePR9n9ZFVRQNGA
jvHN0a7GXbRMKTt8kuGPwaRaZbRxAzp3y0m0nlJdYNk3MrJjPxtnNNE6PV4j4rPg
AWGqyt30mgP0czCpkSBlBwuasXoz2WR23ghh4J5dkxnqgJ8+ttW7WPHqjos3RruW
lgk4Ik1Dvc3peJ7eWuScvbE9Ho4HwHO0Ax23l2Zcg+6RgIBkacSpT03IBXdpuzou
ukFKkr+WKaYmhY9/0z8qhCu2rz/Z4o1URv7+qVNhjBZme12Bnl7iOvEGmEYGsmVR
G+aT7c0t8i4nYpsrUaKADi+iRtwZCO1Z4smS6g6CzIhx7aE0B8gZjx6QKUJ+Qv1p
iYtStXrX+G52bxYrtNtUxRJPL0zaRqHmx12Yu6fQqOpvGz0WHNg5g7h1tPgaDCNc
yR0xdWyZYvkmJ7kqdDMal8N0pxCA5Xo81TzsUBTVkXqdhFi4lKCnsuHnazJsUP7E
`protect END_PROTECTED
