`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DGqLbEzX6LrRXilzFwuk6V4FlNb1H/DtwXnADZA0sh+hEjqICEyQhZ8Lna718qAq
DvjVT6YsAIO0v7DNarj0b/h0Nfw/9zTezHY3wBSGJt/zUuzlQ7S5kAKp1i28r927
Xf9+yxZLREgUkeOWaaqQHKPV/ZnKRTaxvKzD1hGEQP9R+YfLiaRMJ9tLnEuAVdyz
s57Nj/BgPW/spUvDBAniCilCpKrsMNk8E0PdGofB9gJsj5xVLE/+cqQoU2PaUOuC
FYUwoc48kLjNAUfqwmgquJjmD07UlsHUcR7Kl/yP8QJPH+1UH2S2EtOsFj99kjmq
wMvaAvKHLilg8Bd+RpURXg==
`protect END_PROTECTED
