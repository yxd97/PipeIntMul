`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tlDFMWxlQ9L0Vg6/tvkBxHhgmIhGN1tgda9J5NVEQNOakpb22mGiN7DsZngZJFVH
9eOC444h6EhkB3Spl5j15kOlwg+1gm+2daEEXaRQ/mkhr9t2LnaUou8RGx5PPMf6
ZNXOyWgz1hP9HsFi8iHUeqbMaiC6enSmP7TkSSovVyQDbk0XcPfKzgqVzKFwfRXN
YCp0NT9CerLN8Y248430GtMXWaOfBEeLIKbGSzNL7G85FSyfzCxhoI5e4E2PMOB/
xf/Vde5vFf/Jr2xTaAd1d5zZKTUgTEkBfeAYUfZzXFowgW0NKaFZjP+5tVotD6/M
dZg/hVMaWjFayIRUX7IPVg3A4KRqeikLL2E4SdMKyKWh0z52VpgDufBpx9qM5udx
7H/QW3Lb0ewHY4B6LIUvcjRuao8YJewsStarzQj9iMYSKxWifjiB4QrKOlgIDV6u
tdbVUaKaVnr84yPCKGVImY61Kp5yoZw9NMxWHXJvkRhHwHk0XY2SvToPUF59+zMm
D+cQQ9MFxIt6AG7igS8J9rV8Qfzfoqga0yMjAjvr3JU+jR3VvrbwJlb1O/154w+U
p7B0ieduY17Xyi8RqAyzOdTEBQ572BjfQShj93UsZqyt4eHqFVmvkvdIgWmhx0f8
TTqO3P70fJZKWam4GVXu4u2CkCwiKTUq4niLuXJJOpcvujE0UAq3XquGKNTGOd8l
RknINEJ4OsaNfC6Jfss/gaqCJdcDoCSyKJx5q+xNRxv7gdckUn8xerzzVMQDvNP0
K8MYw7z06c9RlVtD20hI0ZM+lahd1zV8XGY8eUyOk0lqtcsE8NH1XUEhFgSWUNGa
nZItW8yx5IgD/BOPB8z4hfLgCZu9+7Uu3Y0sb9k5QapDbzq/4kpd79HqXEDIqNyM
OirP6u6eYNWLmaCWFqfodz+rh8ZRYDvMJTuzqzC6SNgww9fF0AfPu44NsFkTMGdc
WgnU0fswTzQCKPNLlTvssnYHxVHCOc21lELvb7fRcbibKDhO2DkEpDmp+CPFL0ou
`protect END_PROTECTED
