`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nsUdmTfwp0ZU/6aedKIGK47+q5W7xsZKpLdHbZoyZ0kmRW/43aS3smzfqseCNL5E
VZvcIG6ZU1UBAnHX6rK30FMZD8YIBPnsQ2NSQDBOAYGGSp5kcEquG8as0gyNAbUe
/fl7FIjaQcXuK3ZWygQMEOoy3tiQHtXDS09N44r9sob3ykExeJ/Ne49kz1O3lvfo
sbD4jHltpDzC1Wr+v8QTpRXdrbnVNOFkjB0WzWt8AbZxyRpbnJDuij9X+0Z1EcGu
AEMoUcXlyjJFQr478qLKINdMyeBMuPGE9h08bYNsAdy/+tDKJaEMWZ2G6KSRDt4u
VB8yp3Jv7hortcfMCOLSMZLl2nMT1tANhhmVT516FsMlSGhs0wA9B1D1c+LD2clu
XB14SouzYnCPjHt78YxCFv8urXuIeVyj09hwjnQx15ZodllaVZwq3/4tEB4IHGyY
5C5J29lBFHoQVLS3TVRuBRvWTYsCvpSyqfOFLj2q9r9U9K1WvGA+8Ch5JhMBDNZ9
Qyy0Ip00QuumWSMBVHocD+K05fqe/TzmOQ91g+C4IHISNnl0QSe6ZQ2SBgrv1Q4Z
LRPdpS0WjUL6gSBoXswg/zffvqIVGYgXLBpkRvRbE/nVRUzkM7a6xYLh4KYiYT+8
k9+X196GV1Hg/Z422cJHZw5hciZ6uIxntVJRWWkPymZYqPiymW+++40yc0GPLI0h
xi7sCyFezyuxbqrOwAoBKMEHXqBbgRHz6CZAVV8hdV1HkZ+aH7bgI0PfLYDgyJqJ
ojssoVuJtSzsRL7FVi2uam4RJT5ScN+AE1P8AQD8+s2DqQ0BVulcrJu374yr8dP8
i1cUrE0JtQQMfF8oQNp8KhwDm9Aa/WnayO3TgEpU1u5X5tZmpNb+9MqoUyYi/JmV
OikqzquH7+koETfEGoDDJy/eh1J9/pfzO6XW7oPxBNYTL/n+8F5U+iBtDPpKU6mb
j5pG3a7e4PdqV6QGFVz9a6mypPw/9c7+indaTRs078lWFV6XPj2P8If+0sqxIwZZ
Ia8wqM01VPiiG+X0ciX45UR2CYDno49Kxte8zyslAuTDNxldW9kRx9rzWGYjUIns
klHGeyX8BAKEUc364wtsT0pD+vToo2F/6wv7R+SnfqFs2H0hiIICZG/gA/C0clnD
/ModUKDZWil0S+uTnz5/5NMVVwI8GgDWRUfvttrVSDfYRp2Xis1AAG1+wuxIMUAQ
xxm9RJMoORgbOIZcgfyVhz1kjr2z9TC6wQLanWfHEqpNi9GNIHSUkRquqvppqCor
61nqC1yHZ2joo8/oUYV5dz9TqsYKKT3vAvkANvs1vCyBxMNrw+SqeBQGFCttAgC7
9TsMlGjlR0Wi98wW3ojRPNEWGGhmI5GuzTNGth9vHPP1R7Bz6CbCPUR7HVzbBAKj
TwlVEf7pMdqoT5xZ8uMmYydxJHkGPHMffb/VNWlxFctabROXQHRZDbdM4ohsoLNB
j5Y2G48BJFSbj/zEnGuFLpvjenGs57dQbsHODZeOpC0FV+2783DXSJByLjyMaV7C
Hq0fEvCuN0TWIu/QyMtUb3xwt+Hy3CocEpmAezMoVdufKYkc72jims6QnvPUSQgU
DKYmW5AcUjd106d8yk9UK+QwbFocmFa0ewjGRoFVOTQnxDifJv4kImf0QA9PsAML
HDZ5Br6qOaJp+AA1tJtZ2NuZSU2/uIzX3tN2ARGuNz7K/Yh7LzRtujA0MV9MMG6T
G8g00jYi/mKPhyYL6JmY1Oy5g9tlVW9emNBsRmKiSj9KCkmZjnxV24GzUA/B4xls
UFSFmYCy4yrPmRhfYk3eG+1Jehh/FvmvVWbuWZalGVo=
`protect END_PROTECTED
