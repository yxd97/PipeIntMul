`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
78kKVEOyLvkxdz44aCaFyEUCKH3ewzSNyNgqY1V5h7jthFsna5NAW1TSgDIC4Nsw
IODxLrZ0ncLsJxf4u7d17k20JDLac/JapAfXO6ZjikD1EAhD6JxCVwllqXrgpqdP
yiRM5NycTpFDa98mie3is7MuC1CZYQA225KcBN0F+4dHEEBiChs/1PDEj5CTNfY8
I3eK7rY5+DSr501IS4g34znitLGLKX0nTjdiEx1ZZ9R/G+KELA9kYOeTvoN+NpHn
y+jMHB3Z1EZl44YXStYyx6+eB2vw+wEWQQGKzDOijD4r3CeTBxmAd0wN4vJO0QtT
K56v46NuNtivlXkRBB5BdqRtCdzp4zQ55ZTyHY6wf2IEj3hApwFcX9+Z6mhcxT0R
TQH+MLWl1iXLrq5p3mjeAm0c1/LiOY69dDtKNFk8K9MorCiu79DPf3h15tQr9Xqr
h4h8KIc8Q0ooVGHLp8lRtImgmvKqpDDyiFWj+/h+m837ZRg5f8vHoMi49MozhU/W
HruIxRiiaMkRabGdYICfbt1+H33/S9opl/wJAJooaycE/X9H/evkAfZuM+yJEHOx
FVK2vUYEj+BvtGyhrWuzi94ytRs+SJnVMXvOWfm/ChG+BSD+H714lp5qKjk41NhV
SjfqM/S8VYaTvo/g0xHnCby5SPD6dpnd5/aCW4OmO3WMD6gcZsBn55fTes710Gvl
sN0ksBmW0QzsO3x3k5piDfYhOEgdldy3ApA4lOh09vrS7KGTbhtPlCip9Fzu5UGp
`protect END_PROTECTED
