`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vuEwbqhVU9xMF+s+MX6vt26iFZy6Yx+2xAHf3YnhdTwmQz7zF7G4i9n1GWODCW6j
03GZvXbx+a4CwJLiyXSm35mzDDb8oBd41i+YaSzlbGOKQNOgdo02YcMEdULMdqG4
tOl5Ez43jT0aar88hjAiHPiOI80QSXODkMM9ErvPm8uQLRkqNLLUY+BKbvHM/u4d
vtGvs3JH8Dt95E/XVkrtSg+92RpM4uUvLN4KThyn2qw6EoE76mNk1YeYfzvtPFLI
CZM96Zy/iijGCyloDhyK97nC7rh5VugDP/HRqtJKKh90/q2m84WjQvZFHn2mCi/B
yWX9KIpC8BVWjYzrF2lUy/JlW99s6q+EWEjODhiKQfGJBiFcrYhpAK4fGJa8GkRb
PvTEc33ZazDkDR5rCvl9E1bH19nEPx8dRsRcZmTApCkGe0z106RCeisv7QsesDuJ
qeQiHGfDkrsQQFvQrf4R+pUXKW4ZRb/VR2a6fQJD9YXNt5JAD7NEL7jPC7vA5PuQ
JOsRt+AroZz8zzMAdo69UyzyiUOot3gU8GFktYvz+xe6pnN7F8Anj7F/pVlSBqhz
b5gPbblLv6doNXXhGPEJGuoMd94y+QvdR5JwYlRDPX4=
`protect END_PROTECTED
