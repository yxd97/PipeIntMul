`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GFGnVr6y/XG9JeBbbvaK9ldQvGjne6GAb9UxmMlvdnOv/RL99cR+TlR1HYmIhlID
c/BscYsgGDyILwEkguz+FSMLRWAYpMZx6DUw9sNMfxvryNdn/0K5NEBdKZ3CN46G
sKW42t2rg2GMc2nDDsXTOWMDgcLOcR7fDqIoQcvoBNSEl5Dbt+DI+k5yrxnpD7Uz
q6zICJvw/+LRPc6iTuw0wK6AMla/ukMmbSNBKetNvySloXXxeU0sKG+OcChJiqR+
75c4ICn4iqNdrRH4fxC5x5Yk5g3z6RoOuI9Lqpo2l0jzqKd9JEm502Rpsq9Ougpw
yGmySaamTjdDxiwobIGWWeKbrxlS2oD77SCuX/1ngFVJq0FiOnHr8dRPiqk3JDoV
mMEUsIWt6aFSTClUAyajiDsNo3mDiwkdVxfXYRDSKKhPS1kfMGSeJdLHqH3doiyh
8iPtlamdPtWL9Y9RQqePLssu7Q9zxvA7i7a79SkrbUid23YpPcekJrp6ACXL1BGc
t9Z+dl5BwXaHjEpSb1aNJSym/p3tGGrYvzAH3WS2ymaeTNDVf0+/rPLlJBKBUlm3
mDcS0xr1mB+fo0l63w/qK4lmkoYgLTlXUKgCONAEJNtIz0wlRj0P7SrRFzYxtN2n
1b7ypkn9OTMpWzKbjLyI9P2rkpUNZ8DipbNXUFrdMs3IZcSWnT1HdJFuKyJhq7/S
dQ5Eph9yG10p4B3DitB2WwNdJJhez+e4nsbjY7/juDoZXdO7rbOViTNU0tht6Nqm
7eq+ZzayamDp9qW+GnH54na2SJTe6dJWQ1X21qmPlfTw65sNr+ZzpVsAlumOVyGD
14CyyeTGVORZNv0CiP9S1IRlqY1wZrwDxeZjNsOLcTRW+aORI/9ZBHAx060ydKRD
+zY1LgVVq2oOh1/igI0fW6P51ANqsVh6sfUWUNwNmVXsZRNhIemfqwsUsXi33dHM
FOGfguvJj0LJI+HlbJiiMc06OJQlRtkDbqOZHu0n9S8qVNVdVxEvzjenjpeIEef9
/Se5UJ5iwAXU39q7dQNt0P+sy5Vzwdh4EJXZ1FY6UXaWkLcjy1had18/yAKVm1a4
BIck59+rXe+IDwMGS3oyTAmQbj7IVO4ndD8vLvkvizcMgr4fCGd/ENQbYGAAhsUU
uPHKfsSR1lnvKQf+FA80SQTMW3lqckxxsuaR/xwMJ34umZEIGEUjKYrXbLNIHfUv
WnZw0X+213BrBikSYssRgSf/Ys0gwnVdI9V/aTee7+IydX89aNbUQfbeaapDyMq8
bGLmaqDO0QnOM0jO1VgKi3Mdcm6/uIOrZnErHlxR1Bse6kvPytsyCOnZhvGs2Ju6
3+QG69oCA/LbiV/UUUK1mw4nt0uIHUh+C+NymEWDGvJOjDKiZkG95N3P1u+EyWeF
wXHpanbMmhgPwU2Kp4Q04ik06TwEwYAacXRAQNFTEwO3uocuSHDvRW3AqoeS3uBk
tuJ3qz2jsrb0o7l228Ct858+9EX1BnF9FCk/LBUF1TKgXuEYzHVAn8WCw+8uszIQ
G8FWplpA9/vud2OdqBV4PlJg1G61cDavlpB7Yoi/EnpKCeOjzHhMKZJ6W2a5Ky2j
VTp/1CjPxDRWqyF9fWnH8DeH+BT/Wy3qo8en2MxNSzx9HvZota8kdmegn2gPkLap
lWT71iqHJIb7F96Sfo1iCgLIW92x+xySdo8eQun+80khn574thCPEopYwgUSR//2
3UobojLVb6CYjY6432dJ81v4dr+Vua19kFXeQ7VZzDpECUIdU5jd+f3JhHNFbgVi
cIT1qt1nYdTuZMLikD2hNnCdfrfWWru8AJHanCNBz+HPYPVIJBq2/u8ZNu1Awj4P
yfKFfIOhY/hmYwvG4yLMLORB6kQmvIX4V6vs556z69Au8xeikZUOy5SpR75VHTrj
4ScIEsyqOiGK340jwsmXWTnr2dIF7WUyZ8Sd17o0FMjM/n7WzPoVytFjWyPU+Ic6
aVXvxGkXRZK1AfkVeUNzHnxnCIBa+/JypCxmW/SIH2JzrZNNqxyy59Lq9N/kkmOY
PqgYGFbnGjx69gNO7pVGlyBuNPdT74BtBoCrAEA7z5vjvfofiUVZv35BC2LIQRwI
r3pVkV+J0YxnaVT6vVNwSgnRqOgqhqgITerbNuKkavcidZa1rLbpNBtV29H6mwkq
jRzYRwFzpLUStRF+Fjo6k2Hk9v0r9pT/siWv1i7ap0QOY3aGfthixIEYsCqwTLxq
4IzgzUG0D7gnxsXB5ufBM6gUxCR861WwhnXM49CmiEey16QoO3A5OW7/aenIO3MI
CxID7rIZBCYy8vO2MsBVsmbg/XwtjHW3iusOi/Wm/EkwiL4C/Q3YyYXHlvOEQURm
vNyoCeNPIHBm/XgZ2XDItl1xd0LY2/qlZaBk9bMKtPu3x+vfBdGwaXcVzyX0Eb3p
myAxigOwm9LuTfPFLEWzRkyQYa/X1ZvJ2U68P+2zZzmYPASH0/7pz2Mr9eQ77Wlc
MGEbgQNPUvYByPWKKe/QnqCylTB/Znh+/UEbV/E/KJ7I4zCbPG6bgUCtoabFBiCt
O+jX6JWjoMkxed82HtICIjrH3PnMOoXSTEGvhx2rDqYTOEeWD3HoUPDSM/LduMNt
/HikSM8iJI8wD22nZJ1Jlf2MMm7fSCt7Xbid7pyxkgGNponfnIa9aAvHCmGpzaOq
Whj6+sHquQB/KCJUdfm22f3wB2JeH07QaJ/SOrzZDaiHKQdO66cX8X+qgYhJCDDr
IHtvRDVTNYWYDysDg4BvDDQGdFswzsHATwqWzP5kt06i953MMqyJr504TA+RCXii
k9lyHmL+ESiPn3nCrTKQDPUdglMQCTkR3NzzVcCxG4yeb7akaqyx8TKrn+rNTKS2
l/NHjr8wB+MsBaaU6gK3WGC+s6/o7rqQvtJqSOgcTghggEU1lxFlxVigo0HSRZVS
spqnVVjnaBnDsYOJ4UySiNIWUObYXPAl5MwxnJqQBuZDAM3x1xPNGC8yQaEvPnCI
0RBPhhtAcZgG48Rdgk0umljpZ+5kFjPujCPeCTM817uyFpBsnzneoSCrGIjHyGV8
Xyg2nqz/J0CcYr+Ft8gl/gcCUEDCTaWZCY2TvvH8QXNSKQzd2hUMAZzoRl80i4Ja
UrPuaGjuOJkdCFAc9AwzpWvNVsBVKdqFCkg+AL55TurU/T3N7V7kl8zrhHTQ9BtH
XV4/IsePZBNvyKfPbsL+nm6ryF1Oa1adyHIjROvXeOzpp8MANDPzaJr/aRbVyXVr
oA+48NP/Odj0F478LB2IXiBZaClOrsltRGmVHhYLWfTsG44010LNKx2kvBLO/GqT
WGJ4tXfmQ+pRIgT6IgHAN/ngaK7qToByhURSz06/Ohuix1hUVJxtanQzeNiP4qb6
iESCwREKvHCNUWdrdeFM4zTiFXhg3C6ufRNLJppdqWl+F1uzQYOlaEVIOtDBu8gx
rcVnu/1/MaQYDBtcdq0ppqEpHxVgOnaD/gVa37m4xeip7xbmQhIKaFI3Ph4lCbNS
SZ6VHMj0ZhNXmylkeg2JlS7aQDYdzJ/l3k1m3uX8f3fhHzZkcEs2dPfBP2mXIOaL
pkjlUZDmR4k9XNazISUBpjAUy30gErBHKXSidQ7p4TtQtkNun7Vln3nkN2/kGFUp
ZcTD2kZESByMmo64V4EnfrZJ6vWj/m7GM/8AlysitmhrkSGR2pyOagN+teqFyLlz
mYpGfIU2AAbWWBAuFfT/9iOMx0srK12FzjS5GggVLKPSRKYbDMnLSVUGZ7aI4D3L
uMZf3fedIyNUbUkQ1AYXfrbomz7WYNNxYxB+CfnftwXJCZeq4dnBX29k6p5bauSv
QGn8nNFWHekAuf9rzhRjqLODVd+iASVz6uWZlzqumdp2u2LUme80ayOM09eP5dEK
YZ+NmXEO28nBjSBLcXR+S11vctyUrFMjHMfOj5+fWj8b96u69Bz3gdR+g9+XIoxU
Q1RQYv3K+ojOWeG+jev+enLNODZz/XhoIAK8cpBfeTUE+NYbz/B6BukEnRftBQDt
QKIC8AlTlrwFvY4GSU21MjVWlt4HFtItKydVNWDUS03ud53sayi+U9RP85XVI1t/
C3SQdtlz5YWetQ/I8BDuAtrdj4vsKO21rUu8G+a4M/AwnicDVYNddnpBOP6KA7Sg
VBzifp0/ywncfJxFLEnR0R08RRlHIAoos62t8NlUIn7IyBErlUAu+EkVI53CyilA
I7pMdFG/GDZG8nfTGd1+XBNR1jip62jiesJho0zdOQOVbMpMy6d6TUvuoHcs8sVa
FEulvh62vrou9i12NFECN8/Q+g/HHw3Gf6T4c540e2hco53tmvIQu+inuHMkpOEs
TpPR+dfl5Ze6vLZRRrJWsWZOU8omYjq+AW5OmXgcCSDrt/aatSIJfd5ZY3GwDy9h
BrlxjLrJDI4OR4Cb1axPMR7BBm3a4qAxC3qXHT+ju74Rb9iqtxbmLVM82O/y0eDa
0CRbZPxRHA7OR22gw8XweTqzrjnLUwQJBYk8j/3EvEhG+K1BR/9Atfjxj5ffREU2
O9fgAeZdIgZ10xaQLgvgUfAqIJef6I55HKAy7wsbrQMxeJKEJDUm2p9Q2ddOf/T7
KaGlReVuuC+4ep2eoPDONTIGtoGypecTWUpq4vrXlejunk7QSPNyjSQfDXVikIFp
h0/nh5VKcOy2iYcgYxEpu4FhLcHzdG9prtryuBrxfecBR70EH2safzxtMX99UWRM
K2MO6Yx16Ztj2NWiOrov0oUHAJN3CQVPo+wGMvJoVVzvYB97ptb+iisTnWO2zuRS
wzW6XNu0AMLuJ4aJChbwKd+I5hYG+H4zX/laOed1PI5R9yLN4o80wYWEegqimyrn
M37K2m0ciW5Eou7fm37w6GreZklCgK9DzTakfnBGs6FydqSSG0p9R6CLJ5vq8bsX
fdganNDA9fnvcYLrL1lCm6560XeetI8N60B0z8C02yvn22l+MrclqnKyyNqQvR9i
P/6mgK4JVEWd+31YqcFPs1gtRyJMxh4JFagagp2JacU8g/4CjxPYVqRD7nOM7gbB
L/vuiTAb5OFMJUYV/XqcBIla5dKYBdo0x4Jn9vIqb80EMXtAodqkhtjzXbHYSwom
zwXb2A1+0OcJSa8/dYq5KD8BgoPeYBpk30/qeGDw0bjE40bJkJx6ztBB7L4WGcrS
GFjt2LyiDbUspiGR7to8KarDRBk2MYvuuPM08TYZpjNEtq1xlAp1xX6Waoc17R8d
fMcZx/lyiVGi2TwzmDIWV944ATxelewwxpMXGUYAafGQq0fIlD1zfnROum3z36Fn
FlZkumTsAgrt2wj+gPdXPPJVjhGXleBJqTVeEOdmP+zU3AimSKrg/s09oZysBpcD
4agKwDy3qVpY/ySD29eXDMZ6XY2QXjnxg6I9pB8bcOGIoVcDGmoVOGNhKj6nsSor
eAO+QwrjOp2B+J1BF0z9mV0vEwBnqC84y2mkJZHnWlY4jwyBgWh3/CKJk2W4gY8s
RShG0M5uy8YKZFRfeNl/FVrhXSbR5j1S8Qe5uun35abLhfWyyiWp7hmaYTWne3Yi
/g9kk/Rl8scX0nlMWM8XgHxNwKhKNld7IQYrWlw12qk9b76Gs/d1SA1UepROr4ix
O8a9Jzvzb4Uu36b3e7jzqEYQvB0g+KHwbabiFoT8AISi3WNz56L2EzidTw+4fTgb
mqs/TNumQ85U5o3X340HPqspSukssonguy5dOmCCarrOgxYc2JM2Q3BkoEyUEotq
1dHY9L93ZpFtbzVzoA7cdErsIYg3LGFJGX7VzIXQIr65+R3Lij+uLhQ/+AO70Q6s
OmAkQX5xuhP5mhf9pXBo1UeE/xuuStAIA7KEtB7cQO9MTxTlRozdgcfRWet0qshd
awDe3LiiUsQROgLh2katyQQOSWgxhBXvQeqzatUAqgZtEIRxTgXSKNJwS9Ox3f4B
VoDGoNPrU4Qh01VdpcGmN6BF/iNRGRp6M7NUEcDiNkuo99jFspdxsBYw0fgaQqiI
r76gGrpzPHcPV7ScrvkDuFuMaGEI/fZS63Gh/09EKrIhr7d84vXZEqQtb/ewWpov
e9PIqNkIyBJJ/BjcjlK9Pm3zYtcCEn4xyRyddvWeVzLMGwRXbghVhBn8VuaVMz0Q
QqW/5++9eHH7KVAP3N2C3ul9LHGJQC8+yRP7VqmmhbpR6F2zsELFU8bpOsWpnHvG
+/9ugjHXglg3gp+abdajjaIUjoh4427WA229gzPErySNYC6e+A1LbeAQgrrSBkFT
UCxZRrzrNNOgL42dOv9fY1upkjG7zDj5l9jeWcphUyeYdS/vRfeM4uHIFT1kmOk5
3ieU9eN0rHnp2mkf9Uf5QACMTP7QeuFu/s42gbjZ4T5WlQUAiSyY/VJyW//bIOVo
2rjM+R6YER13xsPnGLVLgUHlIL+gXegjmQqa2neLbvJ2mJWOrICv5E24Hqpd/tzv
H/b8T8KRD/dcRRbqNCmy2+XgdRJOe83prEx+Fg6ovZCSutiNIxcQRXaftv50DHu3
HO0hSUyC73XVsQqWUTPVLjWdvqLv7TUQ+7EL2yXZ0iSV7L2E2CSeh/Cqo3E97Y3x
htXCYqMQ44ZYnxuGGmpSmrbiYVyDJxLHO/Sjk6gUzbkVmAE4lXsmygwc4EdrU6yX
NtSu4hwl4evgMsVUQ9N5Tvg2H7TLsXn1Ump9aFGRgAzM7cEidQSXBgBxvSeWCS7U
b7HJotGqrmxDdRcuqzzwrY3K318A63M9RaStDgn2eIaTKl4RGC3nMFVwKjtynJkH
OEuJca0OSosnI0CwnXBa2GgdC+S8qi3TL+Lj15h4fP0fO60qWK0abG93lffLXaNk
e0cvPGiP5gM1DLgD3kTZ1AbcKBbpkSLauLQHRdUYj6OxBUUVFYvHOl5IYt7HVvFx
CzX508eMQ9ehzmcSmcNQINh6CwpfrSq+PvaVYxJ9KWDyDyodF+DvIbmKKb8NIzGX
H8pHI2cTT3Eio0q8XDm5RHcjH2ajN11Qouze+Rmg7HYEIB/GmVlt7X1bsqp2ncml
IV3fEgcmp21dSXLTJGFMRD7d6e1cLpi24YSc7FeZ54KKEyBcwtaHWcURmuxEdXOF
XLRneh/GqdY+hfF2zbkBOK3cF9I5jyE2HNTQSx47o72NTkw0XATnRfTe5NUZPzrQ
MJSoMPU/5IMbRUWXm80+gmfj9o9mD6Z4whrCqPp4aMtfCxbEDOHo4zh8SBhhSIXG
ZAkBNzhAX7Oi6sEcq73w+vzQRkj2YLdfqdbbjMf5t0TMHibTDYr+3w49rQOnhvVy
2sS8XMi1rSz+rI3a/UyG4MYPzbACuCFZEOldFU5HNuGYcl/TZtutFg8jl1A6m70N
KxGBsfDb8a1vUa7iHjACCoYHxn0hGFuzgiZcErdrkoO5Q3z6JHn/3l2am55I3QpQ
fz/VxoeWVnFgRZvo9tPhg393wrv1XmsihYFH+4QEsNqq4RcTEKwFH4NbH+oY8aWj
EPhRhoxPNh39JDBWL3KbxVRYSV4MCFURzqPBnMF/8bAkvWcuLbJZN+iR0dPu0ZsV
ibYyLpDGdKerb+FdKPUzOheeILAD/PMMOh4CtIzJ0oxzRey9R0mi61jyy5JEHWNq
lTpNj8B9vp0DaXr5L0EsTE330nvGlWjPeXO/6z4bIzuF78u0VGJufNLEPVYG09or
mKXgfVCEJErpeDI8Hk6t6os1VmMi762LRdcelXIt2n737hD5pBtDn5T3VOHp50IT
ya1NzZ6XrLJO1piSV0LtMc4It/SEySNjQdYbEv4oWYc=
`protect END_PROTECTED
