`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KEmPeNXDp0y8f7q//ZaOETANja+/kkEBCASI2MPGLvaGtkQXFMU88dAm0Q6vuODu
C2fMzxchJHPUvcV4le8TzOkz0ih4zt1W7fG+p31UFS28F2UP8s5WhDdrMhWiREfC
KAVr8rt7lIXZrwFeQMbFt9lf2zpcSRLuXL1e/oBsHmcNBy5EKOrnYWdjy5lMyKtu
INvwggvEt7lChlKPQ/ij2jcuPaOG8PobELLrcb6upF0FMFjY6+hNjhbQdov6bnyo
T0dkY5B1EST9XvEn2SYeUwUdMHvD3iDkQWPmj1B/HAADVZ13yLS1jFJPaXgYmxqx
j7V5SK8BF/psxL4PJLn8O37B3qZFt7No0HZu3hZYyQzeex4k3eq/VMNnqxTNrqo8
2L9l+Rvl1rk7SI7aaXF4xg==
`protect END_PROTECTED
