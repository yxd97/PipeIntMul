`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3f1JKl7LcHfoyF+u6ZDMLkmu8FPWVhLxE6oycVn9xHgeLIkAx/PqWMH5d/gBOXzN
XOzqOJZz0YQ9VjFNzvYX7BstVKYipYhvVZGR4SPSzBW27fo0Yzdl7NFIuqmywyut
62MY0f697GYEccsjqyAD5rwEEXv2U7M9K2tOOwshGx4gm3qBDakNg/HlwYnbWms4
uQroLZLHt/+mb1PbvQkG22+A+UJaS0CkeJhdPTSyaccRKm3oErDUqbFuyvs7AJjL
cy/EmJvYdjrSKjXPYOlNJPHy6uCSUqcM2/fc8I4Ji3mH8hmR/kl1dgVXnaGAPKql
4gBh/5oNqlhBfv/ZQOOrNiargcjSaEofH7PdtgLDNmgJY3MYL/zqwuhW47tlIjLe
/s6yI77vj/C6H57HsGHfcrKL+fXNVEoKjX995VTFjO3SZ9ih9tPv9FlhLIg78rkD
tZK9hlq1Lqof2uMo8+hVfhtQcAT2g9A3OxnoUkDto0h/HUFZpUNpTs+8P8mvXflZ
SJvraCV8Mog4kK9mOOFGSMw51jlkkNxIfwhhtK2Vm12904q0Wvk5CVNqn3/oTskV
Dc78TsneZgYzZqYHe942Kw==
`protect END_PROTECTED
