`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pzOUKhA3/k5Eg10X/RamO+pAY2naC/gJL/P3eUjjbfLOghY+sfNSOCv1JXb2IzP2
ENYB4kOOofyMIbr3rEGrBr2KJ9xeTVwufiWRPLxwvXMaYh7wI6/w1fN5/XtPyNcs
rs0hzC0FaqhyUfD5uS7JTBWALqcDkClU8IPLRTa4cIZE3AKAymH2bKcK1Ky+RzLB
f1TvohA6k1QJBr0ZrpoIila8jKxkIQkowKIROxB1gbroY3CiLKxtbvUMTFDWglK4
jUFS+T4gNnDlwA6e2ApNRna5rsSUvlWfnTiRqjeFcDioYtbiU6C3D7p9mlwlWNjc
UegSkMMTUN6wyW2zQTupWF/xpxZl2e2mWgpBTTJc7Axx/tVx8OB8nc9d9WZku46+
BMClTv/ST9Ee4g0oYmQLIj/jEkW6C4EOUujlUWpFkSU=
`protect END_PROTECTED
