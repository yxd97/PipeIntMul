`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Htp8cxZJjVvyPOD6+/VJ6Qe3vpgBN8XGuqZlM7nknOnvt3y1g7ZU+iQJWc4DRJNk
Qs/LyIli8ock31MNQBZVEAw6SzrLzaoplEYTtbdAxS1XSTBDoAjp7IqDmhVF5vQ4
a+siK0YB3zeKSl3GSwwHsTF+lzio8XTrGm9uOynn0fbPuXrQJefRa1U9xx3fSN5q
dTfsgdsj0LqNoNPD8WC9YHI1k3LIDLjyrKXzLJf9mRggxBaF3W6pDa6tVXoeR9x7
ZnDj+WTdAEhhl16XSsUVAbUJ5ZrqH1BaXwWL2AUBIi5bpD2+CqPN7ZfwJz9BLh+1
MRMI2ZDP5TdwW/rOrJVEHXcu5CIjB6uIQ/sROVzZKKeTgcoglIrv1qdOgoSOhYEq
Rrdd0y1gcj+ThmeAskpir+aczvhEX68cFFHgD6ktVt1buDQBZC+3yd/1Ua48Yzcy
rs8P1aAtDU8j/BlzHBaDNFgNyNZKl9elet/21dlLrktiVqs7vbZH8I2OWXWokcy4
G+Pm7rOWUcY6unlz1KN86czdV7kn5HfS4eJrnuw2jWSr2yz4BntHstMxbJju3gMU
CxV0Izq11M0tCmNPytpQdkozN2/PIyFRA2C/i2YZjMjE/5hyQZPtGE3Rgf4yIYTv
vLDmOhddbUl8PgJxTJKj03wZ1Xfq8s8zRXTVUX7rnmG6GBwOR6dxkWKigOKPp/PX
m6yxq3P5PNMdo/tag+PENoAHsU3Z3NUlCMMRcil25lXXt6XoYElDQEpMndVNwVzs
lxeEZY2D+Fo+NvfHUwbNi9KHCh8HesngwESWlP8OMO3Usl2tDnIm+UB5eA9NkBBq
rrn+N3or9tfP5jr0uxLVsmjRHv3YXOWLfgGwnz/zlvhWxgGw/ESfwIhtyvBzTdE3
y+QkkJhklz0cuOBxdfk1+6WyybhLsUqptTQaF9Fht4jn3utiXS10taM3rTLbHt4G
/ONz3ejQC3wgEMBLYlWrM4v8xPd48jJ+CFBayjed3CsLVCBv1pGlGr0Ic8ug/5in
8qfQKSixVwVoG2yuW0CSbqJ43FTVfrxaHkOq6C0XPRLfAOVVDnvaXVv9+GRIAhZl
g87uHJDV5o7koynrV3L64c70YANt58/UUn1n3jq9I9KG2OilWRzsZ5x/E7CoP3tR
`protect END_PROTECTED
