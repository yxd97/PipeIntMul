`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SmM25fMmxKfyVV+wHp5en3vdyJ10hYxJNqIsUbojNrHMBVOBtPb8unA3c/3fLmNh
LmNTEXh90WB6Dwx73NZugvhOBjmbaFvj0kolIy61cqfQV211zIcNfQj1ilV6/gT1
HUsuf8uZa/M8ciIqPidxHlC5i+zd5oxpVDtLVPTuDn6WP5siNh4vJdXVyHzKZFOT
5Faq672rE4xf5mlxNb3OkqYqwdj1h1S7+l80z8SIfM2HTgodJlZQmUaegxvWh25K
EMhvS/4QNcKWWGRB3wTCoBqlUXD+jtByvYMJoeHgHKjRlqBxzdmMyCUuT7+e5lyg
vOwQgv5O3YlPZAAdjlqzKpeEyzdFqM7bxgzEhk2JkhMiTWgHZ8KqUcMXoszJp8vz
w4+O70F5gHPrPDFS9eZX54C/LHThYyeIsIyDaPZeVGYs0qzknXqkWDvyYnugBTle
R/jRRSwQLODS71dZZv3RrcVd0CHHLLp5I1uXUwuGwj6URiy22MbhxI9PpjDWMoCH
cMriZbwLyFQBVWPjXRS3FHYc9jnWULVGzZykFCh58X2Fqslf76R6AErrFzFuzX4K
+RqsDzlslfWRv4uFkUs3PnZkgXFcxZbMgzm4R2njZ3izAlL0axbDPw3jJJ0pVgqm
NtZ/zmnAfHjJ6Xb9SNoN+0MoBYd1LfYqXRn1PuCSugFBA71+h6/CXb8AqRVwgM7c
j58Zpm8bPqXFGn92XAExwh9wKYN4iiekxc4hvNv2So88wkU1p2Ox/P2scs/Z41of
`protect END_PROTECTED
