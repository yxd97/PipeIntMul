`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MFX+DFkV5PzWQ8+H9ssc/ppVCJAL7gNrcqtvarS1dEy20yugUtg1VPLB9cvsiSG0
sdJ1lLFA/woU4KwoLsHWjrP6G0QQsD2Pa7RRDoIm1JGWz6DzAwK0AaK3O2Qyytc4
AK6rmKa7RXz9c/fATs5YFc0gcn7pSL1/MJQkVxms0JQeVHfM2jjrWx/zGm6sOZi7
MpLbHlJDzxCw8NuFLSw/VEoOCqj1EeJrnOeDAHZboS26lMONybjAPvhKQ1Bl+e+L
0ddCPzbUmY17lB6IntC9nlrazibEMFixUwgXnhokpYIG9zZYshMe6ZDEQaz5qhzL
wG3WD5KrZYit5lSba3BtXkYSes9y6GjiB5x3puwnWcInHRfz0+G5aMfRxDekDnm6
froyDsDsexOUugTV73++AB0YNiQTddr1/8F/odnYE5iZm533b8W7FScuQMiEM7fh
eSB7bsqRFhzlsNbvMabAJHbqhH3JIL7hkJadNpdyRCvCNZ4XLsXTtkQm+DPuAEXl
+9tW6chkR+qU6QJU/7uXbkpNrF2kJFqbZzSlEhg6NunGX6dS42i0I6OjqCcdhLv1
SnY6RlYQhgyLy2juPXn5Vve83FZvoYWLg4LBr6N15l24hON/llZ9aGc2sNkt0MKH
YATgEefjygru3QQ1837Ce8VtI3eCyAgc4cHVlhSAw8M=
`protect END_PROTECTED
