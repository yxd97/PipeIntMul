`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKcRUev7Qp8ZztkLAmbqIandN3JVTAYbO8lZtS9uME4Oo1PK866BIAiRdteMijRo
y/1lhRjJMS+eAadBeSCYOVQay9vBnBVe1+D8cWXId/IljdLw3nf6oAj15xE/mRLI
pu80MkWnPQ+/6MYlWa7c2Mm6Hn3K+lkfKu8OfgEh2W6Eu7PpJVJb1WzBlmudng9h
UTi7RGDid9qTYWvUEQGe9Und1kE6oWVDIe2DTK6nFP46cDrPYxye3xQIiUn6lGZa
hKJkAX9VKk0zzlxE8AB1KA==
`protect END_PROTECTED
