`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gbbvj/XxkpVJ8pKqzCGa0P5TFI0/6E2nKv9UEzfUP3prhY8svb0NnFb+v+qCc9n9
G+6eZc1V637M1mNjyMK+1Kd78v58ayKABHgogmA6Wu6TPwwBy3xnoceMhQFgydWO
8hgGvHBezoA46wU5cDy8Lh1e/p9HLNVR4vdh9lvMrK+YH62t4iISXXfsWpqbZLXr
gim4fT1eNP/HO16qzvPVtj+4bnPaef1v+AysDNoxvp8JdtRCDQrLL2ugSoyQFYQk
crPEjCvvbAv4aEyAo/fvBAyeDZ1hIGJwECcu9X/H2RkmF5GcoIBDoz1pNbIsBTHb
QTGn+SmpyEon5bQE91csDGsbc9VK9jpFw3gIl0w2c+Pebc4IE0ypizXcEL63BSuT
/iPZGqU3g1H5A2+CoW4l61xz5v1a0T56VKf4DG6x5awkNXYVodOrB0lc9mIUeyIO
`protect END_PROTECTED
