`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QnG3lkTWIUMEwmN1rHXx2ZMC88a4nRoMqIsk29ciGpFkMQ2t0uX24FOBSZQKPEQr
t49M8o8Ki4RldKZS4LWpaTrf78lbVu6tb70OdOV50lD/QkvUpjYEzeC3V6eUCzZp
d3DBN+dbfOBAfWdlqpuhlYPcr181t/fM6sTodffK+LN+WAZ3loftMLz+sE5HNv29
L2PL6/jHzu/K4+0DRoDtQGHi0GHPG9FPX5WbbxUKAD7MKruzpOc5pNHoQgrzwp4e
eCsArmo7a5b4d+RQ0AO2sVkrmWx1ZNnzX0VLvPMrniRfvzXyEMZJxLKnoIaviTXS
W/5NYfkYZZv2dOVsV0k76cX+xysPUOUobBWP8FPsQSXXGhQc30PxBjX8nTa/e/d+
K/CC5RZOjSVyUexR9uyh6gTTjZhT7BAcH/zbD52IpaY=
`protect END_PROTECTED
