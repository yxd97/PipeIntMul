`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
psR326xc82OqW1Xjv5w5WEOqWXketW6u9fun+AjjcW4qfjHInCbUu2kApDKd8Ef7
PX6Q4C8S8HaymA+PCEnk020Jy2NLI1yWbaCTymE5GakS/ipfwD0SQXSk7UBXWw0k
vU/Q6YjFoTagxg4b4ocCkk/A0fn0+mCiBmH/IvJPx12xD73EEGatOCHOHDMC79Yp
//VcmVlI89Due4cGcPYMfot1JrV1JHztl1fMi7xdbQ6tdjEtFFNQ9coo0761ehG7
cJLGPl9qu8CX+Onhi4tIqbsIJ9R5H3qJXUrkQMuMVWnQZnAwrISqrTzBJDKcMCi+
DGmsd5DtsOt5pc2VQarZdMZiw/fzY9ekCVcfHFGYVfv52SIGrxnfvLJdQE/hbet0
vgL51mztiptic38/YQiSC8WyxMPHVNgR6CF9yEw4DB1ydS8ebuvN73mwr5Of/vYN
0bkHho1d8VS1gM4rE6bcDRYBZnhA6Icb6Nx5tx+92pt9hhToEm4Hn7sujf2dV901
SNQm+MyOKBJ6b+WV7imt0l4OOIlpwMhdvCQHTruy6eZyH5ByYFXvl0k1uZHETA+Y
wnRKn9dsySQRb5/RqheJlJWsr84ONzzr0cuMl1HiINGUCUjukOuvzK5iZBf+TcLv
nytsYYZXobLlr5JAQUfKtrMeGobAjGN2N6rWlgyOEDPDkJZ/Y5y9YMEyUHRs4hEN
QLuNlcEzvjJ+amIAU5Gzpw==
`protect END_PROTECTED
