`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QGcre+fKKt5h+doCEBur1Tgu2SLjNME1nPRqUuFB1fVVwAIW3edv2GQFJdy3AeLR
hdxE14o8dysPGOGkFPsxyxN96+xmWr7v6kDH1EWtOAKFTB9tHOBkr2GWHn7Mfiyp
puTXKQP5EcXuumk/ALGpU+V0Y/s2bl5QSPhlYh7A1wG9blPmnOw6YB9uP10j7Cof
BFfGgwG/PJIf4iYDiW54PGslfMAP3IL9LeTxck6RWVDe/aKHNHsKD7VYxoTTqG2y
7P0eAgGmz2nkG4jPn8vfoeFpPK5jPrMuDTqTrgxHxM3zg7ZJ1eXgUSdtOkakOlci
dngGljtfN3d3MfoYpXGezuA/Sx5/5CIn3mArW67CGcwc4sjq11c7RKMPbyy8V3uU
xsB1QJJsVGdKdByGxPF6TXZPBcmUWqGrmLevIs1SAOkktoWO4LfZ73inQPPKjZ2c
+/U/jRAD0uux7uzvgfDtdg7hpte5AuJ1cTdDEY2h4Y9azH8CA2bzP7O1KvPvl0b3
RwGo72zNzbvkaXE9un/f0G98WVTojPJXBYb6lYVqF9eZAsidtpSJXSZATZxpZraq
MX/ZB8Cd9Gme5sY4Hve7UurVf3WCDqdqu396q6W8HUq61QoaYptSfe6uEYdOeLMm
mhne6Q8Y65a3iBu3oHBrDA==
`protect END_PROTECTED
