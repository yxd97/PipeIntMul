`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Undaddq0CGG1GXPcP5wZySaZIuc5DHYQRvd9qaBx+h95NabENOOzf9p5HHrnv/hj
Hc/elBVYRgsE30pING3OigzTEM1QAopilufFYr5fkeNGltuEi3TuM63GzkkanBw/
bX1OfdAR042PvMpKiCgfu/vLAvNXjptVH1SdlyQxZHaMGSo28nwWPHO5pfdXpubf
rAZBFpBvipt4U1DGGDiCeNpMYINc76o850RRLVGzgUzltit3YJhMYqOv6zVMRE4W
HXXza4ZJoPAn3r1P1ItznUnM3TJgDJV0PZQNU/UKSAedGaByqcQgSw1bNR9/IZ9/
JB0Z6mV9fOyPpDf4sogsZQ==
`protect END_PROTECTED
