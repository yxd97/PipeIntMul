`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZMfKcGe+Sw0qozswyUVb1TOceuWc7zwXBl0gHO5mF+fw6Dk6HBeG1vyGw0S0+Hww
xHaGxnVsRxe4Q8frKdjc9g90+XAN5pSSz7FlN2fkMs27mGi/g96PgyHCXXo9zq+c
WaYsk+5SM2+ZjEwCg2sIJqE9/5ssFstvIp4PJfoKY0GxFcfaAcptWpMbSx7x7NgR
wTxTHQGNVa+9gOmrWaqrIzvCkmAAnLtx5ssvBwStOGsdG6alDhBy9gMAJ5U2Or4n
fGz13LdYVHBu/eNpI6Cr5XEQNPnveFmcRakEpnhrb09pZtHZHN+26Wi0lfF4oM5X
oX+zuu2jgJRdKzOP1+XA4lj+6jCxi3lT6gURxjQqmhLvEhjPnGKTV4BaZQg2kJKN
sOuOEZnhxceON/LIsmlCV/W85QDfI1gEFJ6mIxn44Nssg3Sfw+KcaAyOdgejQPp6
x05+tjLq/59xH5paO/Er/mE4aTcIzqLqGy7wAi600Hs=
`protect END_PROTECTED
