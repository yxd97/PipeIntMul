`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
egmCuix+ySN+6vvXuPXWBrktT9FwM+1S/Ax1Xu5EzeSzdyLYPfDC5WIAl89Gpo54
9GOYaYHpjGAOTZP1CBbhnKcMQZmE77DkI9pEplsxyX2vgXqNamzNG44c1uysG0y5
4bTSLwY0peWkuQQ/ahaqlGlJk92e8/oLWM4EsU743ImlGjl5IkvdtZJVpP1ORWw+
8clqIUPbAJ4yg+TTm6woR1fEOXy03lUEGz2aEy1PSSAONSfbYXhbKnMvs6PyXz4G
cqxS9jeUBNuZSN8JLE0+t6rC3kqCYlWjcpHQQCLJ1RbpnMr8csryTr8NrTlM7Xtj
f1vk7Z7h2czqp5Q9r3+zkAlvvXE/MUyPobGM3fOo51kPm7tOl6W7u24CjhdltJM/
xXcoNLrWjX8+dxq2e0ggHuBz0v3pIQiYw8J2RBMkmSZg2bGBpJLcalJFlC+xd2H9
NIZhextjh4Xj4ffTpaGM7bdGlLGsAf5GVbur8RmbVGM=
`protect END_PROTECTED
