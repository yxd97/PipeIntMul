`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YaDfoS7oFhd4JMrtU8rO3Vbh9K64xf2y4AGOBrLJ+XTbG6r+VHVTPEqD1eBtULRN
ePyZtK6Gdg1s+uHGO3wYZmO7YuoKesrNjNhldvnMsosArmI2z51qySprHEyLxfTI
c0Ts0Aog0b8mw0TC0wK//rtyQAoqn23SIpmHrDC9WaRxjYlfG49QuSv006Gz+UAY
DmhJwger8XNRgqmydOpLdldvo1D3NZRqFO/aGMh0tp+3IW3XpZttzLcRZmSGTJy2
TfaQbzBOdbvMG4Xn8udZ/XBuLiVOP+OxmgOoz0MLwtmDGyFXkBufZgLaZBMQFt7F
sbazYsCzsGKONMkIcdq2Oyofcf4H80jVYO8MbkPLL98N+4YeVWgqYXOy+RWE+24t
cTZNVgSuB1tbfC5RFcSUcXxnbo/dMlwWcv4PQrBcMD0BUPfhXulOItAAFacB51YY
qE0oYRaf2iSXjfgWWxrS/X5udSKme8dp0g4PwFqnTte3MOTIifjl3QWq4/fUol7V
3dS+kY9ZMtmuHWkI5SkW21YCLBiwXDvrmKiT22nxcxcWegwYwUH381DpMYJRdDLw
iLxWxOheuBVwokZAxIORJVkVsZohL+2XApV7nzAPLhWi2V3DQrwOiaENgsKKcIjD
v0AttzpERZzKPDLbo8GGJGQ6f65wfhwUg8VruXRYjc7eeT9jtH0L+6BqKo6tCUq+
O5zBrCzRuvSdzCpebCvwMaSlyvYbg/SkAhmZrfX0EvkqhyzY+BLqTgdlzKYZzYWM
HFIipmE+zqsEfA1sNEiuY++CgYoBdpt1s3uNk7n3R+XuhkGL2eW1FPCHVIlyG6gd
QhrAgNHHpl98u+4cdI1+DlUcCcjTaeFcDaC2XElfORWB6XrhwLhckhEHJQFTsP3o
Vd6BW3Za4O3DQt5hmEHwJ8IgruUN/6ABAonlIP2YYHFsWVbUE3ifCZFeepBxnNKA
C8/Wa/2LxSvCaSjcptcXdQjl8swxRmQU0x08gUCJCWBOIjKAFpZADAid5tLtTMMb
gkBiz+yONncPp3DNPwhtKwh5kBLaGn2zLnBzTkvpNkALF/+woerUWL6dJ991VQv/
DrQ+GgBSJtc4ZbHYs8dwmlEOVEb7jSC8+r2eJYFadU0xY/9XAJNSZjqbaavSou+B
IALgzQa14qQiIjSU3KHQDAT4GU5L0p4glNBlh5Qzt3tKJysh/RcrA/fMhixYLoQK
mDdciG4AD+EENt2fI0dd+Uq18MjjOVBhGlaoW4YE+mTxxyCXwN0XRfURPAOic2K7
E7cw0QJN+37dRt+9Uqqib7pZqSZTkN5SKJC20q7gYxBok53uwOsi13yVZXcXkLfx
7ydrtzPbkHw9AHYBKpgVmmsF46bWGfWviSU3zEMiMUBoxIZbB0FS1YYAf6EQvkpF
v0vns7QJixk/jU5FgBGIPAs/TM+1FYbD2tJXkl/Fz9t4DZW4nxMaWfczdW3k9VbU
cNuhZBmybRegxdjli9nHzy8UiXpmlkJGKjHrIuWIZt8wUm7AXAk8DIANSW+laj+X
VBIZfv29QlFH/FqKQ4JSmi/+ucrOd1RLCyPxgkdGXLEVZpjVfDz8PgVht9ASGmcQ
EyTv3lo8BgSwfOwqVLolYkC4b1AdFNGjemnhwbP3OyxTqsAUacpImdJrLSItGE4Z
mCjCYDFhIfrQGXZZo6D2lcTAVexMyLaW4pgaZXLUNbRaUgYhdibsqbSn7gM2yKlm
ZUN/pd13bimFBwShPae4iXNFLulZ81OI1P7cMcClhEeQqxnxqr9tsN1tZLFxxpzi
1MN5IMLBkVKP1Djxv+f68vUdztIiSxBax/8sRrEJwBqQzFEyFy8+F17I4II0GQ/B
l62Zg5DE0UIZjSvvynaIYDq3Qs6vPtEBRInJ+Fc3XN+TVB06LwhMA3QP9iviyJGQ
HttGOQQGL522c0L4lNZs4IPfrME7zaI1c+6OV6+GyI/RC+ZRRFbBYmlMw9M7kkMV
JMTfGOkyOrPMTo2b0J7eew+kWz7R7ZudqFgRXP1D32QyJ8Q6zEOtQmLCRwwffGDY
D0P9InAj33O5BBfVeLWXfB+lyz80QH2+8JP80PNkcD4oM1b2a08txgQ9LioKDO/l
6kCKsKvVId8Y05ENBvs9+eYaPOT8Afk/oSIHEKdt3LwWqZKltiPo3DW4MhwLA3lU
Oqv6UFLAJ50efWT/crPQ98YBSxDFqYc4EAUHBHS99TBfKGZplwDjR4hY4N+DgE4D
Jn31JBDE189nqk0ziFL9/kOSk/R5vQkKR29WXRyqsfC5EG7iJdGnIS6vhbFnnFdh
krZiz1cFhi9Bm0US3khqdnDG5PSzhvg0V7seR7otUd8qFyqoJVQGZf11Ujit5va5
YGKspKPxeoJtQTabZq9ojFqfhAwOWnt5ZFwaaEeVVMi8TIFrAnOYfYu3PUtQiMDz
Wj8tMx1PzZ9FiJxHwNZawhTwTSPAkQ+aEhK/JgovMUoN7OU4Zcmi4r27O5LQcE+j
hEAdmbZDb22R+HWfRz4yIS++d3wLpKLJsRq8qLD5lbVpg+vpBDpE/94/87r8RAiE
vZqpMhbiz4yJE15DrWFYUqboAiQopTJV+3G1e8eZXlXXUG0mmEDcwX1cCIxuCSJa
XsQJ2fE+ykyEFSN+rEX61F4GTljkXLFVs+4ffVwFwTUEev6yB1/BgMjBihUH+Uem
RhJ/rYfTjWqEyaIXjGGiQ0Y8ndotuzbmi9nmbk02y8dmSOs4n6toXc8wl2rcSK4g
5dl3x2D9MpqB1jSjgxdopkisZcaRuC6uDc74wTVQx6N4XPOsFwNM84/wVaHHJEsx
NHy53egoM532ULtnowgVTrjZ+0yyMuNmvxWN7cmFmmagUpekNDuse0mM281ymDXF
nNhtE1v86rL/68OTVxH3eKnz5RJlxV/MrIjHONiAsyOOFGx08TkIt0aSHAtt2Dqj
O6IvCqwpynDKG+VlwhsEMza0RnLRhIty8hnRy+OKL4/2KpHwAlAfo+kTkaQsKcN5
A/EEUcf70+A84SGj0jqnIfuGOeBZgYCPNMi3vAlvgWsipkyko7/IaudOX4NLQRLN
mbK4wUDttOWWb8njp2W5dwpaUAEDzNUWm6EX2b8IwJ2dnQejWOublagAm6yqQA1U
f5IwVebGWEs3aQI5nDFuBTFjdriirMKgtE4xHV4d+Q2aWnqe7nanQlpWTVEj/f5Y
jBCfTEoPuvjXosemCYGD8ThJ/4FAOJOVE8iEWseCZGgMqpQQKflaITbXQUf92pWN
sMexKAghzEyLoOBGe4KzwtSqkv3x36RqGOtHZU5/2d0Ci0JKOTcexDFM+XF74sHw
RHfHAnNlm8p87lTRbwYUyXR9yujoda+GgocIRZAz6n0dJT52BAXJsMleAV0w10iC
8nDPjAHzZhev5mzabSWA2TixaaQvQ1VrEFF7zRSIzlE6sfJRe7YhXSU+DfJQPMSQ
iqgcHuFWTcB88g/oldAZ5t2f/7qnx8950sOYkOqWNA5VyqQwjI51lH1if6Ysxtp6
gjPBOTyEBw2nxFJO1/04hPVD1c/SoDyTwBZkUrWtustFrdKlF6lizwtezy4MMnEI
J4LyoWjTJ2OpDxecBFQUZ5VizPFNiSfSBWbNIZbjwd2uguMpYUozErFuALHJ9PSQ
ffJSilziIdPw21XjDrbmZkU6PGy53L3qrkXBhyO+JP5TAHIFlkrhlxucLwm1s5Mr
JLN0S6DZHhz07U3xfe3m4Dy8kFbMdR2sP9ZuDP29C/w9zosoBbfHgnT4Th99ZOQu
RHPZvzea1cirAdeRhkWMFW6ZAWMGKvUTKsWWRcDC78vEHsdlPyJh4Z+aH8+sYvJb
HVcW4UGjKd5HrwKuTPcQuwMznYVqbU/aNwjIGBmg1ru3gfuWZANWDtsDQloycX0a
JreXEDED0I44y26xBBGMscpVEGzb2PzAe0HSiJn9/PBGWkyYhPZdSep2TkLeJ2Sn
tW/XHZ7E4tdmmLd9aldUKKgCw9Dw/PzEaZe07TTM0RS+tld3By7LTI+0hcSuhNW0
hwpszQuVgz5G2HaVf9eD6ZSJXqAxIqnlDyRrkvMj1NblmqMit94VuLDXbe11eiMC
ffMq+bpOD6o1hXlZBYqx1LMQYLyMpjkFqGFLr5A7XTqqiZWXx7BJHrI9BAjxk/Te
gr9I3GhPgyv6+6rsoVgX/9xikJ6ndN2zoMszmzuVJn3qiKsaUblczoKkgHEIInXs
GLqXTVzcgRoE2AmCpr2w6Ucvg2V4nkR3hCxFfuyC6UIFUci9G3l/X4USDchM12N0
1L3XLlKTvRnObxV0VyjJ5Y0zQYArIV40PgU5G6ZmsiW+VK79PkF4LDSPxImO4Sy5
4kMmsvibvYRD1u7lRvUqlidYTWXjOCNfyvMvSu5AGNLNZmZ2Q+flsCLJZaX5WA/T
1cQ92wgD3t+ecbnjsNbuyRxg3Yle7a4hfUwkTbThXPVxa3HVoRK8LsqBJPXAl6hI
br5EK4g5V476qIebV0RfYVlwOOf7SnK+x/jf7Pq+uWkDvbpx/rZpqP2Vw1EcuX5H
e6HOqWYbIWQ3Pgv6HB3ZksbDUvtDsIr6WsDOsv2OAm8YQnZoOyRBgrQt1Ja5bKdV
yyLohJ6kDsF0/fqFEpJiRSb1ZjyuhH+5Ff7IwbqW7jYKA5f2yln5XiH+MAbblUMH
nFqQi4Lmb8Bf+a930ridGFLcfW3jDQ0kgzMDkznbk0RAFf5CacQwxzY9MdAtylRM
13Vdc+xq952halRenWcKS9cx8UWxCnEJBY+mSYUcA5Jh5SdV0C1yDHFK60C/poyw
bHCzLl83z3sDrkNHZCO96S4jLPeFgo1WFodsvawiG+DYI4BfUpLKoaUKAe8Tu96D
NRvufTYZB1CxamVjQBLVgJ46CejTv7QtDJIY6jOHG8gzPndyKB4NoIvwIRnmNfoe
TrXn/zkQM4JXDKKOMuQ10Z40wjyaeg0Ah2blQkiGl4iInj3GmwoJ/fKN1z80440S
ZmIUcMg+28rb4A0W/Qv/dKd/lzlv8Zuwdl3CywsVmyPNleey5CadHjhW5NcjDINj
h2H9IAk2iybxzN3hUjwjoqddd9UYQ+p43ldcUCHn1AIY7kyTtz6CgG3CrmAIWLWp
Agm9PPjPS2hZ1zGjvVwlTNnnIz95ZAkNylobew5CKvn0IWILX6KPw/PxYeonMajb
ACGyVP0Ow63k1JdnxDbXx8WYt43R6eGiE/DM02lFkwGjsALRtZJz5CH0tUu2LWxw
OkpJReEPAUJ9gCCP0HpicqwNuXap3WaK2FR3LZV11VUFWNP/jLNw9+3UVypZ0vQb
Laib6asC+nYb2tPU1Es53EFr788fviqd/1oqDPn6m6pT4+J+m1FoBsqQ1CWBAtcf
3nPtV1r5Y4vW6lvruSNDix9aG01yHme0mFK6+rDs7VbLpmcC1jgvzFlT2oydkMLL
q/ytPrqUW2cotkas6CuRXGwUaaKlFZ0uy3nEquaIfUn7WoGjzQH4VFB0OuIhrCsC
eHt91FMLRNd0rOGJ67BTirgEF0aHgjHJFehkIfieDZNuJyHr7LBp4aVxl/G1EcyL
juo2Ctw7U1yBJ9rzJt6bXJ7OkqQvGl1bdoK15lH1uRfXKJ+SU56BthWHoKEKPUNe
EFyAfaVmaTYETvAqqLP68p/KU5hcNSgF17td27VpBYjmkyLuSsCOVdBIcqNoHhrc
wpx+M/forzyeN5zsU3eUbBWqdKp4rVbhPPih3WGTFFHSD8Jk1q+OmPsCq6wKKCCu
dWvBi2wkp+S6GWs/pr8VxKu9uZyJ/ZEgAR6TemNEYBHtRkm2Et6N7fIdFA9iRUT+
D9rHmHHVaIDKhH5xs0weQMzo1e/pu6Xy/tA0RgM/2dHK8IYkKrtgLOj68MYDBqe4
U0BkU1Ls9V93tqRGJMMucJCi3DiGkaXv+9ZkT59KiRfTW9+zhPrNlBU2pSupNaI0
IRchjKXMr3HvGYsaqaQHaVFN8jCod/qJgzPvnWMdawmGHY9tSEkM2JY89mhDWePd
pGmuqQq46AWRdbHmjuK7DO8Vd/TKK4uXvVXLIQF4iiZOoEiHUURgvVkQ2/xAvMrE
z0bA1nW/1xrkQypVTi3tcm0/f6XNSn89Tjo3nJAtWyajgDeXqaSqwuw2upTHH5Ph
RTmAtEIsU/po7zD9J4+b3Zy6Zz81jjNUQncaRAmLfEJeABvR4l/unsSAIfbMsMVh
0+ZlJs4cseYMLv1/QoaLG1ya5BXo1Jxbd9Zn3WPNhlgtqcUJy6qAgKVjXc7Z8IAw
uXaXWyoslSgzIBBWP6E0lHBl71P/DsmeIKhqp4Y2/2c=
`protect END_PROTECTED
