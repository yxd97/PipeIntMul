`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
peLe9LSiK9n9DuHF3y0NTlZvBoHM41+H+E+laZzSUjwuS1eCWPB5q4+u3UOtWJgr
LX6RFTVQSIcs+b6R96PbX671AMdnXuD5r3meYdNsebfut1TGnD+MPDaKfMyyc5Al
WLLP3m1b7eqHBUq1FVqlYxHVJ5BWhZeYuS42hmTAzDDjeEGfUx/OwqjK8A9mXdZP
9Z7v7DBhyMiZSngYbnq23I6d4dfwm2O3RkyIlaARdZ8Gm+PKSNfgU+3npydAoOZA
yfidoREHMUL/Uff23UNIGLAK5p/iUy0KK6Lm5elkucv+Y3UtPumghUpuQIHXqqqr
ldRWNci+F7LgIS1vl21U6WF2GMID4CfPODzkWNCWOwRBizU9Qrx7Eq1/AU3X4A2i
wAdDC54y9xv1OLWGhqw/LRgUNaIhZxk19BfjpX7F4wzJeoLE9R5mc/CBelWc8yME
KmQ33oW9fNdYcCJate3vORZC3Fq4kSGCYOMqVM2iPN8W4QNzRgQ5/kZBHOvVQ1nP
`protect END_PROTECTED
