`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4VhtrVSUHZb8uoFRLcJiwa3xcNcPB1gMV/CjTW8S76vWU1BdrRXc6wOpmeE5OlxK
Ox0N9Q0PUfuOedrhzGpdLaVbBjANeAZ36hX6EQg98qNznc2SbLugm8ILWp8xeSxc
/SEU0AeUBC9NdvFNTDvB7ZASjJIx57aAcqLMwYTevkHpAbESxcihxHIJxWKnEs1z
NtqQaCYnpNZ04H4y3LobB2/0F/uOTxzLWofkfmtyqaXRuuBMYqjo2mdE4XmGKMPM
6r90szKAzERmV3Bv6QQMT4azc7VG1cmx+IgXEQkWDLpTm/CvT75L3d175fMKafMA
LdbwSiGyv++yFQEkCXFu1g==
`protect END_PROTECTED
