`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TV4GQb5H9da1Ye5WvbgFzzviMyPROQXoObv/SNSmxm95LGZbiwDQ6iukNp49Z0Rc
OyakFaHyhaPOmvvmiiSrtMSpd5hWMBFybBzEauStR4N1nsQMW5tqOx0bq1fKlbNF
O4gPYJ7LUziUqWXJ/tv7kepwevMucAnxlIlc4qQPuV+MAm4OHqN8GjMUTzCz7Gts
hf6v/m3z14VSr+5iVU2U6ZfXNldJDrrmcxDsqxG62/jq8RDep/52kzGxlUuKalGM
N06JOsN/FArQqAzU39b/B79rGXyy9hhR81gwC4ND6IU/qhviSwFyJv2g6/qT/2Yh
0v9J0MGQohyc15FzFTPka0Z/JMN00ladaPSDwIR4qUS414G9bHxhIDrVriJkx38o
0Sf6R6A35/EtCMJ5tPcIetF3Des9y4LPf3t+b7ehqbakdb+rVZYhFv3fcCEBfizS
r6WvnkP1/BUnrsN/9MHRTucA604+sjmHu5fJ3849Bw+ZQQYLPVKyhQ5F02H92t3h
XzZ3a/jqPMmyR5xu5BLaHIQtIwdMfSatYO5Egpo+3vk=
`protect END_PROTECTED
