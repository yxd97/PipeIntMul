`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lKLRKazyteIe6jV0vscl0yB3CBlgGpZxkRaqvOig8GET/KN9SZ1UYC1Vx5WZwu3x
rLzlUgKo/WGvW53LymthxzuQMittzEO4J/C8MfOKxvOWNARP3mf3h0D72E5Du9Nc
kBIvb4AKjX0EH05dWSWw7djLFsEyVFmsnMBO7QJC41CPyoau6w/tucNxyA1CDCTp
dG11HKG/E5uurep7sPI2jIgRhm0ac94mqKv1+W1NFQzB1p4NPfTqqsnK498cvIZ1
v7JI/3/rSGr47ZcazOpAn0P8qWPaby5OR41JPNRFU4CKbbjUlYDT29dSQihLq0a9
kGPxz3InErz9HHqXiMQ1c3geWlWCkXPHFwJHJR4V/R7dIj+leb3cs90sO7rP1Ylv
MegzqRb8id8AS5ID5AzbUQVE8YR/S/WPVnrC4E5b/+E7wrm9Cp6IPlicJTmzEmWy
NCHkyXeE3CwO4o4Fh5A+2x6YyFTQiXvcmfWKA9egSN0=
`protect END_PROTECTED
