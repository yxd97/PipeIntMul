`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNiJiJ4xmgfJ17aSNJP8qWRVKWIxzuWh80gHB3oAvUroej0aFZ4m9ooV5swHOvmO
X0YOEqa0Xh1Mzi5GYrIaSdMC9QOiN0W/8CtFL0ImVIu4bm5bIoAex688kGjfLvpN
PdIELAgco2TqnENd4wjhCV24O6vQTkmdIwr/Omnv+x2TtHFAHQf11s4f3VUqNUZg
edoR6uXgIT18fhbLUQmVoAlN0mQtReEVqMAj4RhIrt0ClvDv4TrS2gvf4eP6rdfj
HS/0zajWgtdgiGNTIPq/VE6M+1X+ExgeIRWRzxCNiqDiLYpR9ZQQdFiqD9g4RbX7
K84p0RvGNwKFcyrP6JV+jqve18wLcXHo3i5t23jbiX4jwMrFBo4+mqCa5QNCVJ0L
DtTplbD2loLku1wOSFaZaU3udlgsPRvGD4zMyVVanCBw8YppmjoEjPEUBaj28q+b
cja4B2wg1fdDr9F3XFt7SKo2COTG4V5eG2+I7iLlGXl15RESTE6kw1GY9rtxK1hZ
lXvVCV7He662Q2f3SgamBizw6bEF38OB1FEJlJ/aBUqit9VVXWky9vIYWJ2A2krP
s/YU+7s9ey42gym00ZTATQ==
`protect END_PROTECTED
