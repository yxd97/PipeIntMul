`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bYPRIuVIdWNVuhI+rqTsAbWeUNGzCrQrGXdbhdyPRzZI9SM97AwWT5euE6xVvk21
bH9kU0QD82+4xf0mQ9EgHkilD6Bhq5WNqgxLznfaHmLqsvbW+lchW8Zps4311aWQ
nVrvvJuJNHGmWeUz95m/1XBYJnEMX/+qIGWOQES9aDpMSTKgNclkteCZQZMBqWK6
/yO0rtFaBibfE2W+VCBVmz/6Fr3+81Pkwmg229/tO5ctRCrq61YZYur99TLCA2GO
MZ4on/1P0Het2fhYGhxPhXcRcz+HAhayKdNIW96pxvIPrrzqEyA4F8D+DXZxIwun
zpULFsa6k309Ip3orKKJfd54ZLiy3FrGuXlesNAGCFV5IfK27gbmfyU6+emBXuND
Gzk6hiHdgBC+NiwhW/uyyPyibGJGjbVNmMd+RmDDcgCoUyb0PygTtE1rzxSupkGN
Orzam2PjfqcVfy4DmjW8ikap6U7+bdRdBTZXxWx/YfMIMipukrk9eF98h0wlc5Wn
Kl725S86mmCEl5Vj9/UHWRjzzK4QaCc08+Gn9udh15Ak6vTZFmOc4/w5zNGzgSWQ
5/oDs/a0GwqScX3jl5j0CRpy1DkYiU3/IJhaggPXt4uV4G8HMp9NUnqlWM/YDhNO
xb/lyHTkscep4Zau95OEUJrfbYt6rOFt3yIv2/UeRAlnli5KaxPMIeqS05URNsTw
DMaB2IWUhzo55BIWeJYxRxUvBNOgEBX5TbqvelsLsgML8jjhscReiAaDUWf8SnBp
G0WEo1KAtLTp469qgZp2KjmodSHUlxGmBJpPTNWYtxp+72aSBU1wT9r0FhrVYLUI
4+PQDbdzcNfQJzZz3P0KxcYU+sVbyCywKyZdfuKzDIJbccjQ4DjmCyMQW9Bgzmtc
LzPNrWmG3S71mPeLR2uFYIl518hisjWFwyPYvZ2Pe3eGAYVmSBEVTZWaqiQZy1qH
9l3ERgMk7R7yZchcFMl28jPZnFLVH75zhgocGu4hgqrzFTegc9JwA+DrAlDd6snO
`protect END_PROTECTED
