`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JMzoPFDnlBqvhlxpubkuXiwoyHXpKJ69N4ZFoIKOCzR/2VbNAoKOgXWKvPUJHjEl
vJfNHHwWq28SGYC7N6ylbSvidzRfpIGPoVzBagHrHMdIsp1aQIiiv22SG197gJ2E
d8sZ/ihhpGRwMRACBpk5l3mgOTz5KfW5jjniuSSgnogMQeOj32XbvKjPwAl96oKy
fVCZSiwuiMpuJ8cMDQTwvkwEiWNsfjF448y90N7eGzvng3jozi2OVjbWJ7sa40K5
ZwiGRE+0CBWvJccx1/E7Sm98hvPgWa8FmewKKUthi6ccrZZ3fRHEJWn+uIytLiuh
U5J9X8VH01lZfPtB2zd80TIx/jEt4rGerHmtvj/WzdAZhwElkj1f7yiwOHRa9ygG
aXNyFIL63ZOIbD6FJZON579YY0mZneMjxyqOmbkAJKA7LSJgF6S8QuPRxnCe+yhC
q0RQlzSh9JyDLEyBhaMQ4yyO2bkFoB7xsLDUK/+QW+6ERHgrzRCpxzN0fympZplH
8C1cqBDUSn54bqSxHid73fO6mF4pW+S0rfELfYhGFeY=
`protect END_PROTECTED
