`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6wug18ukdy3a11sHQ1O9gX9eCgrGZqdOVYEsBa7lX6cIge58MIa8lssAWmPoDloq
0GH8KQvkLNnBpVoKyAYraQkm2ebbQlPFb03mlDCbMgF9HqI/90lGux5Iz4HRKZAg
J6sWEQbOGe2Z8RU0J4sKpzgTjd0oNWlM+cisjqKgiWE7JtYrDTJ/3BMtWAMUUF4l
ypj8y1UsPscsQ+oWYv8zCZEMq6ovFE5RS2zeoW4AZxwCcNdE066ntO3vYqewbLjv
Zx2rR4WxALmUml9PUyDfz+YdK6AIvaQhrAi9uUGAiIbTi1Eln/cqktBfVqDosZwI
M2PGxEjVmQppOjXT6qUByNpb9IaR2IAlDx7f0D2YUsTsbXZ/a9MbswX1BKwB+ruH
sritsYwBdT0hfWKwTMcnzLOcjcx45uUVca1PkzVwruCFRzGFo+8VQIisumSZNSut
qpkMAEpv+47CimBPMIbvA8mPo5aDHF/0VpPzzZMOhkKyf+WJwMZKnkViDkmsD5wy
CRFd4NqaYK8MikMdPzQd/OlnqunoWgi3jDPSQ1ZmUS/JTEoHYPS4JN8rIe3/bo/i
2zhPXfUaaRKvzPp84rHFsk/kGBwIIQHVzQdGLPcTOSSqbcr/stCkKQd/rnOFQp61
3zix26g1bnkuDRzdZk3vnxfX3jiwqptrt0AdRiVmxVblVlvq/TySVN9uY/LOMnue
ZAVEVvIb7HZZ2Y0IDTVoz8M80xdFqcXoes37XcLstYF8Sp2WsnxlpusRxn7LuVgz
f8DjSMQNoJlP7LD60hBu+Y4Y/dHKN2PHm0vKtyb2zEY79y+wymmKi///ZKKpT9KK
8KZJoCBJYrWH01FARlcUE465kYDDI5GDaVVxM4FeyP+JGLnvm+y9G7/GdvkfK+Wt
vL8OgI+rpn4L/2cfqhzFVIjjQDKdgWPuWLOba9GdkZfmyAt4i2A2suszk9uxX8Mv
w0XEyKStaZygDyjEcmC4OwAQCWOx9Ec0v8Z4f1TNpC43f/u1lHcKEWQjgKaAFB9w
3H5BSEB0bWFfFSiCDxrC34MKpwaF2A6VTjA3U1a/mtZCaU+b0/tWrcTqnoqzWaYp
3mjjWPzNjlISjIN/xnajpaW1Wf/a/Cqm+GCq9puEbJ2mI81ggRthebVtvDIIWiei
Hyjp/LrbHjCZ2TrYI0co1zU3/M1ofHLfD2ESR0XQv5AzM2GXOS+SORdoC1ijfi8d
e3Rzg9MavxQ78TyJ7BSyqFWTXJCsYaM6vnEL4W2kfdqjsy54K25bZ+y+70WHGXD6
g1w7ML/BsLfHVw+iYIotq40V/f0/Walqtpr7LOKhrpxZGMC/2lg2V6S4WVgQdTy9
6gsSjdjVdgQR0jF3mYu1kJmIdREtysEQBEzy3qnpvnklDLlZi7YRLpIF21DnjEWp
1wR+hsD6y4Dd2hmEcko0iKarHytLrODBrEAqhP5creurcJcHi6hHeU+JeBy++h1O
jbcIkGukL+sAA3oLL5ynQ+XU2hZIw74808k5P7cICXyC90inlfoq8mcpbD4cneNM
8mxd6ny8A1O0f21yyYl6/0ZPBnHYdEmJJgfGzj64ImIUBTWunVOEkW6jFbyPN/hD
7juBqW28ErIBKVRPmdy97e7lZyv7TubFVxilWrHlJSOfWeSYI2wTn1c7QuENV0tZ
QDxHsQOAmQhkQq4bSjfwVuKxMN8AXYml9EF2oU5mSpM=
`protect END_PROTECTED
