`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ifucrxFH5iMirRbk9uUdnc2otEeqQPn6gyhp1U/nx2Mel11/aoSJepBzRQEiO1xT
SLomUVcVklPVajZbdHNqxEgs23cX9smbN7uLbn6rBPPhR75BmaRqEhrnnRo8u7aI
8AlyY2av0rt3gCPCc0qqBuN7Ys22NfCPXiL/Ac9sq9tX4l8O4LDbLYfp9a17dq2Q
dRyDDDQbUsgs3Jd4vk5jvU4BGkQsDd/OHZFSDKw1wdeVDDjcM43MW1KpHMBbwIde
RQwl+4lyhARsgl2rhjHPOsLVxfwkbyZn3OYVBZXUtBeBOu7Z15fF4DraLVvSx+0k
F7WXWvv3B/ewcDzLyUxZ2+WSAfjCtELesdSTyJUXQxSrj9oms/XD2OgnYMLK9xmd
uGcDbdtZ2zyD18C1f+g2nY1CMOWKiNd3EcRuYNT1Z19ysfNQBGEFiLEYiHHAo/Av
roSwapPFLqZ2nef18KrBJq3n9601A+3rU6LPlzz5e7fq0MHl3eXYmjL+9u4OOHxz
drxPS464KasIkOpvhN92jTaTyV80k8a3ZowUbcnzl7A4WeKPq3v1I/Q8TOAdaQ+Q
3b7a4Bkn1rcJDlyGlv8n9Q==
`protect END_PROTECTED
