`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5npmXrO+jowalS0QGdOVQ/VKtGWFmfGBOh+C7q1wswJ/lyAqSLF2RkG+mc5TrmrU
N+Fhu/o4KA3fsRKSO1KQ+fyP9NO4C+xHlA4AJruKCTK0PArOVU1lzBxKP5DaR5GZ
xz9wnJvxIgncJEqHZV3kVFF8VizWbjqc2DXgyv4/fTT596BauB4a0VMqUGGpx4zY
D+MlI+qmpalev/Pj0TGajJO6vloNshH10UpT1Jha/MghPk5oAqWh+Q+n7rA9B05B
6sXRWO+5Y6jK7rLXkOsHV73JMEGKaniMg0AFq9V4bA504oHEiGIge2D3TZ5XwIO3
FrdVfSK0GXtu5jgwMsBqFYvAA2M5tLNEO5ZA68HVZUM7d4IkMwKYDvs0TVSLCsfD
boR/kRuabAe4oDER43uOWg==
`protect END_PROTECTED
