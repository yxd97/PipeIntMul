`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4n9cLuGqlDoQLF9hH9P0526ZqhVLc97mbNHtcjV4vnFmX1MKN3d+MA6E3rDiSvKJ
GXbEk2OHTosOFCFzBuXkR1JGUYJPmetPaHO0byV5Jdz45JAc6hZJycrQP5u8aiao
siIYQrs4VJOrM1GZr6bxW/OPrRtGPAvOz/D09svsfgVrS2+1Eee0zmUMtjDwjyue
2o/tR2iKd5XqgHALIrSBuyAWXa++5HFp+kTILAxKhrD2b7Dep5vcnnA/PM/QO/TM
vBe3Qb3Myftm6dEMXnsfmsK10qajxo4qD4NujleQn18nSB187yYwrS0HPRigmqn9
7OM4EbcLQbiAvcd40VfXjPGULql3jduGFnig5Yxxcwjo84Rd1cjpEut6K/LVdxtY
hgR4yKnz2TvLPb241ijrb6TDC5VOXP+iuwB3ZnC3v8RQ7UOO27O8/cKmLc72GVmj
xm2ZRINOGcMeS6vABg6C9uIkdnULmMYBhgwjbFN5qJl7bgBYhYAvWerKM2Uca9MS
NfsnkPCaQEcyz6TOD6WW5LDVnH5JZAPZMLBeHTR8c0EDnRqs7ZkVBGZC/S6KMXTT
nTbU1DC+ug5IlgHjLPf9+vZ2nQ5i68dsB+gbXZdVBkbzWo6KCOBkAaaQ522cm1mb
FU1WYy4juzlZBF5FF17Pj+QUVzOTf1wFdHorO0B9MdTSfX2hESg3CFYNh6yqQYzo
Q0pQ9YBFK8R5ylanS7FmhePhlu3i3982haGra8SuGKtmfBRTwFnQ+tY+vXtBJpJr
5ZuqE0w3QFgyrzgM36+02M5wZHRJnfnW3knT5bB63PqLi9Otay8LQy2jlyYCxDg7
qBdgWgNJtsRM0H2zAlSSaN1gTeL0h3o6tEuQYCVFoDdlLSqy8WzhutzOpa7E/uI5
GV2FJ4xmUKJv6Jp4mp0h7gfD4WkDJXZVwSq3vl047An32x8WzibUKKJ/2j/dR79l
dXhV6JRgGVpWRTbo/u4X5g==
`protect END_PROTECTED
