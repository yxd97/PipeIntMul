`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XJPgRyxSv8oE0zVWluYoP/sS7DgyDifsLGiwEReQzeeaiFMyDmYaZT2wdHvoJi6F
St5y2xY9VKq7JtLgxTL7NCoHWdvT0g9GXsZep1gXKD5rtS/GC6mpfmpWpZMVuPyl
M/0+XTbx6LQZyFztLZfNxwZpadats8Ri459psghbupnjUy/4E4dSlnETG9C5h03u
fhL8M7+jHrkZBIuMJn4hBbgJAwgiTpAiFWZw6XSH2iNGEbHfl0SsogYYZ0I9KQjM
cUA5iuqgUj8lAiwXCuccP1TLOwwiuNZKmSqkubDaMcxuwbMnVIe76g0z+8N8BS2t
zEW/uKXSuDpgdM80J5rMqjAEsSQMGy2/1IB82nvqmEvXzTYtFSP+Axg/JNO0sMVe
vQb/SViiGY7QC25j8oBO4j4dMrrPGMfkzMO8LZec/152+oqnO5LJkNCqLpBgrqg2
wiGUOpIepfpj/y135Vg62MNwcZOqrduU728kL+IRcdTWPzGSKhF+VjLqJik9C/uw
`protect END_PROTECTED
