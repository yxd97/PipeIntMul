`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UuUEoq9KnkdMlhuWNa0RFv1nZFSMVZGHE2fBGgB9nLcit+0p401iYMPRVBiQ+XGS
apcfUmGmHWU0ADm/QEw3Uz5QURqKohD8pBnSNK4QllGOu4xsz8vD/iNK4WB0t/GC
SzoHNCAPZCnMQOzhEhOxms+LaEUy4HLzEESLWYd/dbXauDlFUUo6h9jBcf0Gq9NT
UDNMZ1II6flbLlOy4gOLlVYInANaWHwFyGyXYc/QCnnyQl3s8dJWxEXu4ZTgRyjA
r2ORSfmrJaLgQj49I3eggPEMJk8eJvOe7OsEWu8EQedKCFhmDGrvI1/ivML5fZXR
P3+tp5FZ6G5uahnlYQY4RzIPudm/BbPahvsM+GvHp/k=
`protect END_PROTECTED
