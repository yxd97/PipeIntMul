`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ucTDIoomE+4AmDBrCyJAhyMz3zxZtvBdoDu7h5pv+MB1NcxZ6jFUtXW9m6oI5Xar
vOOxt0mjK/sJ+SL0qnrfACranGwJdHezk0RTxClcGTxcTnWxPchs3f4M9A34NqrE
FL7s1o2KkTi8wGqS9WnH7hFQHht+iwTBjJ45RA0L522REqRLO++cUPygJoUa1A14
fBr2zUquu5hkJMguNT4LeRPOAIGMHBBDbSmZkSRmsSSQEFuOMiySLEyRqkJkRH3N
4Kpwewl9YLHi5bhMO946epgfddSAuUjKcv+lneBZ3IAYY9rXgB1XpbAVW/u+oyqb
vQW3gOkviJgzLYEe53HPJryOLmlktIigS37vHhiFa0AxWt3rrVRhF1XmSzleLwXI
6Vva8QazCq+C54AtaqmNRA==
`protect END_PROTECTED
