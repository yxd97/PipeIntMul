`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cAg5MoFmRptn1+hyw8YCsCqGTkMHBhCJMdwo4IPtNqpOJC+pJX08zPj7n+EFXmVZ
1XWmat+y2e7fu7f0P8qdCL3WZ9FUobbH5xNFjoALZ7ncVaWArWUPPG2b25W8UjjY
64ACbczqLvmp3gzWU03hK0M6isWSDi+pQ1W29Vw6lnwb/AvVbOn3MNMX4Gx0V/ve
TDhiVjUX+g/KDjXefrT/UwzCFwqxFMm5kKfSk5ISCzVAJFTNNwQyiMqLyqnac3fT
`protect END_PROTECTED
