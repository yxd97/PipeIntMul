`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bh64TsLY85rBKl9j8gDMeaEGx9aDCyxYqmwlfzqgqmhwYutCLTYkcl/paKGZSZLV
o6od5Y+V6aF3pQUXtJIqZZJW63o7G7b7YzjFRGL8it8qoiPzh/VWL+kYGzDHpEKw
Jg6VO9BRortAlBqO8NuFSdJH3CPf+xsZFrw9ybab80Qumxyj8wdNoXbF0sk31633
u3XiT+agLjQIQV6emM37hHHnXnPRPhDVVzswLdzgTzRr7k02O9cPnRXSQlHY+hdg
ZSw9cCuV+KfRPLLmrAIVqRQIIsZg1BrQoHHYpst5r0wlooPtFT5IJfE0Iz8q/F5l
pxvSVd3K8Zr6FwwoM2BYtd6EnEiogaFuEUvmbKmlLw2QP7bM8Daq+s2HYwNlJpTo
/XQ7EEdDtaLL3Iresqx1p3kSfejKSrB/vr9eApAG9NrqSgoaIKvjpl2jqcCTKWm7
Xof81CpKMV4axv8hCdtmlonGz9nc7embnrZ2lcq1OT/iH0XsAt7y/3Y7CWdDDjid
xLT0AtuCyp9fuTg4qGwK9+0z4xQaeCd6G+0oouu/is3HU5diKwetJ6DjNC2dBWZ1
HPf8Go5et8orAoI588BaqvQD3EsiGZQtuv+iDRVe/R7dum4vQvYCbQjy5V03UQNF
5PqUtFG5fjVamSuMRjNQEd40ByZnKlKFtLq9WpplhEy2fWa0/wFhGZMg/XRV+6l1
LI8hvBZO9rpav6zfPzGPXXiLxC24bFP96KPZGiA0VC7B8XRvhhaT1uHI2ah4z4HC
fGeX8SIImTjzPli1CJI1m6ZQYZWRxEzRUmi8GszR86WGbK23v2OpdAQ4RcmLnMel
0hCqcvOm4Z9ZKATEi4ER/PQqF1jrhJMuTNoHyi5u9ISXAdqRNDGvhfeeJowo+TR/
MoUy9DeiXgnhBsi+yZ74ihteGiURJy48Vt65LVC5+S3FdM2z39kSFhMwOy88HmH+
GLAmIrGg44MHxSCPKuKFwQvz5opmtfwC/Lm6ej6gVMJLIv/iizxa/fumTpVk0QR6
DLyKldR0+fImH2LLUZ6r8gkUeWQcKoz6C/eg6ZXQxhTE2qJEqVYyA+GgSimVHSH3
eHXeYvbxiC/dDzUkwJMKNgybCbKE1C04TGl2pyiK9ULZsZtsT7ZOlxrytbA9Quya
GEED/Z2URamLcpM/OEWVOmT72ZgwDc8nPvi/H0EW5mrGtBQUPrhbbwo9P3qSi8MC
88vrYNZkkRWxUgi9D0E/zLgGCUp3OaNoNp227abIUkSmBTqO5wzUCLHKZvm4t3bR
nF9Y/3QvPbkO8E501W53SRgj0zbF2j0CciFbc0I1ft1k9XtZ/vxJjvUVIh6ZBPw8
AJSyMjna+ZlgL6b4037w2sPpxrokBLahfhvypuzdsPNiFpcsTGbRSo/V4YwhP81U
PEO5ts8RA890E/Cvb7ZWiob+X21m5ZCamkmNF46vi0ZXYPZBQqkmfGFohlhV/bK6
4dv1HQdSIquY39cVqN1Ol1WTmSWMBe351D1EIMHNaAAlcYWUC9IJcM2bizUtSv3c
JIvfz7x2PjoDwTzyLI2f2uz3ekHS9W2pIMYOfLEIqVZbwwoaGryIyZmCBpGCl3ZT
uT5QSmR2yJhMW1QzJS048d/WjsMMBJ67ntuyLGmNCZrj2oo2vUYRWtKXpsUHiEpg
/kQMXJzy3OFZHjDgAj7UGNMFIEHBTPcKw1lhuwElnxlxK0BKtsDjNi61EONQgwau
`protect END_PROTECTED
