`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SxiEvmW+YPSFi1UNeWDeF13jYmQ+A98kM9jb4nPBWshDKm/BY7sKg2bbg6vMdocI
W/pC95y3NtEyncvi0MPzdm1BV50eCQ43Gqvuqr3WHtZIFIwvVl2Url+z5i08be8G
AKxTEF72g5wxMufPKCOrqSIV20ssmlh7EVpv4d/wslM0TPYPGFintOmbGf53Y+S9
nyQF2x1Ct3XBqVGpspwLp39XpNFQv48giXdgDNyviKnu3dEfw03kD+ZXUH8LHeru
0OCs6q2mcuoeReadtAWe6lVp8mAAoUL3OZAQzkv9jiMvf0HJUJzfN47ImBLEeJOF
Y0BB5z3KNqeK0qDLjoVx4RDr1xlvBKp/PQvLH7PhfN1uDxUwlChE6PQCtmwvQh9Z
ST7sXa0tRToZTdWR6AWMiJjhxRvdfxU6MiSeZFeiosf4XfXwqZO+fOGerHwvFtJD
S/7AG/138r2lxOun7n7WUh9uQK70sna2JUExJDTPP++OlvOF6RpuEljcGPpgIBqb
8JsneduGSsQ1W+JPc+pyQ/KQ0CqNqbLoUM7eR9muSvS5SZqqtbOZ7IYHvAz78tc8
`protect END_PROTECTED
