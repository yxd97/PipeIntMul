`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Ok76/7vNp6GKMhtT4m190HYRB7UlQ1qBAA83kH74uGWG2JR+JOo8jzBbRRsYsG0
auSSrlxu56CcMIFPyTuih3HUXtppjeyjWWhKyJrZsjVzWydC/UyYLbragAeZteVn
nih/HPQCWhnqTnq5rPr0CUvxQAaNL5+qtKISBDtKzwE/CbrzHxSkeqry+Hgz7jmf
Ug4yNlgy2LUKN9teF5YtDSGwpIWNVpVJyB+aZM/jrhYv+r+hPoqxYDBxnXucvBqq
ASRIyBuu0fOkpBvz+KXtlF1KkRmkLggwRc7T4TP3leC6g0I0Z5pY+0wb3JoiZ5LK
JfEIRVxWchncKGOnvGihKjP49tq99JLW5G0UFTZeOptt/yPnGdE0KA/IOgENhDX9
xbAODE4/sbETcv1GWis+Hz3rfueiphH+N8Xx+pl5X2BAPUPpZlboXwg3B1G3i3KA
cRZTlbmbTfY+MuuB8rikd7/eNiUim5Fg58Ow5c4cMHdPqiblm1oB2l7jhWvMrXfo
ZZqfMt6lTfpPuJVEC/LRCOBMWjpypozoIQdfrBgZ4GM=
`protect END_PROTECTED
