`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bnuap+/T0jKptQfCgyM2R6loyW9Ok/CSoGA/a9VQwxrWLnUlOLk7j7Ts8Qsfgw4O
UGawQ3PeOhdyAujsAloLRGb/Dedzgcxfpm1GtFabiNGMQJ7FwJchTNBNVHwukgQV
5dCV0lNz3WeyRVJOaUVPUWCXfSoh9pIATylUXWQa62/ufV7Nb0CWVLe38Z6qjIYl
KxEjQ0mBfF09Raqm/5rhW9GLyvOPbPPjbMGisJYSFOS+jIUoKggQ/RDlWXYP3Adx
d65w8TLWUUhZXr3b1mlFUVZNm08sZmP3Nyz+KdN0sg6xIYT+LfytMLFW/qMjtU5c
dkrGDbN+kAh3iY2Z8F6a+1raLywFIuXGNlHaFTpbU5Lre1VTHiD5s//iRa/LtVlz
`protect END_PROTECTED
