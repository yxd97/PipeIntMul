`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YqHBSj9zBsc1hJ/29yROdtBUwX3rjNEA+Kgm2aveO023yWsudID/oKmV6LgSTqvs
la5YMAH7Fl3U8oSgHl0JFRaJ5tGzo4SkY6XAPrffH1CM1yK8ZebRH2LgDEoidJLd
oETIc/3ZbZQsAbb3ze7ONQNrGRJbr0ezl5oKlw3eaUN7obgvNY0SBcDNBgY7mWLO
l56tV/hzoSlsMGCy4XPkxp4QJw6CE4QQCjn7f8yPb9KCv0BPP1QquIpmKn4aDnMJ
kyrX+Rxr2ZiMT2/6H6eaBMcfj04IdUZmfJUFVGp5EnMz/BgBYZLPBshG/QuakZTt
TyHueOfKzP4z4UTJYFKL41zGqtw/g7KIlU5OZTxcWHMkzAywEgGNBSBAvOFnqEcd
ukjepVUkgPdI1hBzXCRp+HBZz5dnxbudNDqYW6mNyEXoiOE139xbusf3OZc1Sqbw
17p4jFqQDwlApf5jUAsRJrYoHjUwoEBAlJHlTcKQtJGaWGtPNCsL+MQzYqIRMX9e
bySsj3WR2Hd0Y8J3yvSd5Q3xYia2y7Hz8xIGfDp+b84FNbQB5coqRIEbC6zcbHV2
18IympJslRtOM0r0S/989rKlMsDrZ9jRirnZ1daZxY8+QOhYe1u7J6/T/PNwwU4Y
K0kbpO89QOyPsDfaXWLivzaS80PWvO/EfsFgnTwHjFLJl4JvsZmSt5HfaXJ1ph3R
JtffJjXDHmS/RlHcWhBGhrNH9/JC9mj3XpyMDrkyhrCtQwRScCHC7a0xX28sLltj
UjT93iOc44Msd3y9Sj6hdVSdb/jPUzgZQD6kmFGpR4+hKtZUfA7VsYvj6CvJxN/p
gnHGuqWBxXCrjsv0qJoH54FQ3f6TLHcWsl3+OF2oE4nhA9DgUqW3wb2gOtGrlFZW
keyTJzRE+MELphjqHtcDbK9CQP2K/XKEe4U2Ok0wyLOiKtK8JffI3zEyNLSBZOS5
YK2is5soaw0XMjgQg2/fycjzWsaIM5p6kEzJDswvPUSD2HIOvgyngyT2bzU+pSi9
hdY9hVrXJr1FsaP3wyzioqUtHN673NhgkDOG2uYQMf5OOYMAJVY4lM8MqAbqUImn
5kOGf5i66u7fGPYhwLdfspqK9gQMzX0yU+iFyxNeR/aWqPclGztRF8bx1i2uiluF
6YnSFKokLihVQLW9pM8z4uZs6zXtvlOuXsioOE+ymw9ABiPhhS5SRHCRSvz8EiEx
nZsA94kUe5PTil2kFJqSnk0NJMgIpaQUjYcHSxOHghzmnvgbDWa0WnKiS0OwtrUf
J97NmMXCH5W9soAmcI9ok1A89DZrXV+JjJWLJZUgKWpYrJgCytaeXowkmEu8bM1a
hhOx+BltrLjcdF9//JnMwXcLdrlzg9JKBhhp9MN/T5WkygGnY9jCAVVdUC0kPoL3
cOd+y2gUGB2VUpCeahWkaa91SmQCqeKFhGMrDcP8vtXmrXzhnYUj8quN2d5+4vKQ
tauUfEqlVF1Ojdoox6oFKCBaUBgQYPke+Ug7cl0hRqOd8Ls741pIW4N3Lwq7X9NL
dE9qf6djQZ2MGnyk95mTSAqGh41LJc03iPiTznYO253jvbsU4yydv4YLVqAB7VRu
ZjvXslD8tkXc/jMauiSN4NO8Xodk+NZYt7dpBxWvSx2EUY0dJmXjjS6jtJtE6C8v
cInqliJPk28cGIISHtUZ70Di4FyP0yaXfWQwcbri9/BwQAuTNyIrb9g+e3ndrpnc
+puJQ7Bto8gp6i9UgJmojy9yjkTK5qESr6YdVPjO3Cp1gKWkwLnCQLsZ0sDqXjgS
R90ETpxCB/A7KC3ygLbMyP8Fq0FbADSuI1tVyy+RunNoUlRcHjMlCZIkDpihx9Z2
HDzh9OaIbi29U6++/ng0Sbwww1WaWlodBIQJXRwMRi4ScXwGWIMcnhu9laOPWVuL
u9bPFmb8+mgNfVmmQsS2WabVLR2V3zQlM1EADJnBTU6Vz/EReVwwXKy592uAXEKh
ATR8ETJuc+eJTpYfxOYYNxdJ7GSkDIxo587dWxKuoJJEpO5aR8ejgJjKGikPHNJF
UrYlbsyULzB7GuH2VuzV+8BQ+bdLf6i1jMw1x7PVA7OoeMZp5evyIpTEPzgb1oTC
NbPLwIQuCj5tFzhvMqIeUE9reArbs4hvcflLXadnWCkKuc+S+CHGCb1nRmgIgOi9
lwmEz9XjHjTaw/JN/0IcZylbKt1uFgr/KTRm4RmIvV42PdJQPzX19mZNSlQ36wB5
H4zDx4iBPWjJg0pkTI6ZKERmI+mmbcTOfSDLFGQ2kRZeUb3HSX+F9rQAqAS0Nmya
fcckUIczby4OQhYjdidxjOCT5v9EaLqxcBzo1wKSgVgXXKH+1pYT1yul65Z1hZCh
9k9pjqBdIG852jDuel/9bD8NYGx9N7YlU196AgUle3TwB9kJ1DNciuzUgonVfN1O
GFVdq0ePUQxoaQIoceJvfBsdO2FWjgQvPIHNCrYBVIdBvP+FRDgAt8/fimfYVdx3
u/WvvpCCO1tWKnJ0WM9BjzV1t5rls9iSGtyghH9IwoUKTjRL7TvBZ27HHEUoZ+tp
gpV5evbrN+O0OpjO3sNEqPg3PG033P/+QmhBE0On3ofF8+H8Vb7R+zC0RXMS0zhl
P4ZzBLx4Hg0SNFbP1zGFJ9IDrq4Jjj+Rrz+ho+9qZM/xknz4QkM8nDkYZEpffwgh
wiHolaPmqQ5sTz2ogkWGyDWfYuHC8ORhZGaGuFL+Iz2fc+rI0kn2QLGBJ/2jwTHo
D96Ikkb2QXGlkZuc13vXq4T5pmxhsCjGPHn66sv+IR61ZUFMZ59PDH5bRuVVagBW
31yh9AsvneAx8DgUkZrOGkMh+IUb6n7SpKFx4ZwfYtYsnwqcAA+gsaOrKnpW1Z0u
EmEbjDiGP19o4l9PjCbFhC4c6Zg8u87H9tE2Kvhxs6wAt3Y8SYXcWO//Ntl8HDjq
HBZcG0gprSqFrW/pL1nVpjMyvEAyiYSe9N6jqbyWWPyFJoX7BMvzoBRNo3gIjRYC
wm71NlDDEiZH523pTU+9bSk97nKNIREssJ+pNsSqrPFsv+tEoAmq50SGJw+R1hfJ
DJ10zbRHF/Y8grfFyidl+iQ75YydpELKOBTJYqBH1DHQnh5/UgIzDKZrEC+0UDx/
EjEqRsz8W3TDuaeH5mXhgBUQfP6hUjXKAcsWtWt/AAXLQGBwKe7z3Towcvt0XS+D
Zu1z0JB2pu3M13sbNWh7wjqGMCp53REBwBWTm1OMfPwLJMJHPvs8rzLaoUQufeJb
nSw0pYQTN1Uk4E5XdDvMAP2Sg5EtADLZgju6pZjfhcg0HgG+Hv/UkhbOWXTeoTSK
HZjCKthS8gRWrk0uceOucv29ViTdD4ELCfoIIpuvesS5ONN3VN4GLoF7acnQmM9i
BpiIJX6jsPUu+zlloHUU9bf9SZHoG7swv8LdogjN5rZADh1kmf9OItlhd7q83BbG
5xV/6nOlpQ8ur1cAN73L0546p1wiXD57zdh3K9XmFO2fJSJi/1DNTwOcB0jioz76
NpkKpTpPUJhnBe2LlFXZsQfFeSjJRPDibsX3ndpZ4MZzurlOZqk0t+z3WaHtHUqB
ccDsEQUH7oNbmiyr+G1n/yJyNk4N6dxvYFOV4MvOOOquVqVbkEnlZgeI06cWndwX
JcMeliEOHTek4WI/BtmUShQflkmjrD6n+4zEW5tlJiQY6Sx5ozkduupz05iwK8tr
/0RXqXZzLP2sO0uE6rceWBrOwxGKvbGFcITJevmpzqisLTkxv9qejXt4uQABehwE
7mlG4D5vx0sLSOeD3proOu4fce/7/mgiNKktfR58wrYscGe9CAXt+lqE6c4PTysZ
afMMSI+1Q/nuJl+m46skODwneeGXLVR8Y3xfKn+r0/EHvUGF9owYezDWUS7PjZCf
34BumOW7sGmstMZpuCF+iB8O7T7VYTeMOltKZGLu+Tt9ijUs1mCi/Jv/KiWCSI/Q
6S06rChyJQDestZ/2w7i4R6UmGbirKz8ekl8YiErHZwIuR9YswfCXNPTPuTxcMJ2
Ncd4wbliqFy9XrqguxXfuL179JTEsxrFtj2bo4jXabPy8OQTSPkgX24A83Z3Y0AY
SFIgxjAJt5YCyy2QySIM8Se8p4ZGNYwA8i1MbqRX4O1u70p68Ed6ODJx2+4kK2jB
7xS7Lcwn7peLytbCaXIZ/TOa4N//3KmK/TF6EoaQvO75w/LrWiOWK/4b+ALf/1Lj
7vdrjebdTgUmX1iSbQSg6sJ+KhPyriAyyeBo86KKFiO22HaPYj3cmJUG/ZOgBfzx
Eh248ITjSq50zhDYCsyGZYcyAG/f6AuW9SuxD9em1+DJRLldJw6nGWLYcy5QvqFi
+wqEtAwWHXPiylRD/AmBlJgNZuQNXLyGtHYH3pwC9xuwOLpJTBvf4D0hJn4EQaQO
Doplbtn7TuXxgscLzZi8OvxyRTlh6LMplmn6Q9zwOKLsqgY570Y4e5B84tWdCmLI
7uhWb7cvUC3v5L2QID2DP8zqwbh7H/ZAKGJdzyE2O0l+3/ug48PRdUMb9snI2sGw
mI06Ia7tddDNUNziHxc4t7gfRdwtkVMi3+5D2N+XlBH9ypfhJcGdojgHm1K2PtEu
8sJXpvd51IPRKvTUxW/s7sM44dUAmFnNslWKyTAJtEOFgtFO3A6p34+qYrdJ4Xw+
GH8FoFCnDOnn7g/o3Nyhh16b3pXqQKJ3wTVsN63n4y9Le+dtslqpvs86LTJh11PY
e+37oaTBjvfOE91eNEFpSE/DI8B++cZt2n2zPtR3rexBIqCmBfa5r2kk6diYoJo9
2fqj9sxq1RR4NMvXHbWePwCB/11bLTZetPUXsmlIraXVi/bUKPhg4FLrMr9NpZaD
qIjASzohYkGcECxpjInRW2y9p6zf9Cg7OUyyrcOm6QJd3qnU8OuvH9OICIhQQTwZ
3hybtHOF34Z0N6PJZzKbEb/x9O7vim2qU1VcU+S7OyaYRU9ENnil5lKJLru6qgZe
mkm1qeqeEF2TPutcOmiUABfjg/QyuLg9jo0LvUBG9+vB2rOzoIZyra+ugMApabv/
n1YqI5bYtrmphUyOBwrZScwrRRHy+L/YjtQdRm4FmziaL7l4oQylOuBHrGVNa8Q9
ccCXLQfDtv7xx2ezyyeECAAq9NSMODefThQZS+yFUcFRu2lZUxgag6Zk1hYM1fF0
At8XCVdEBGZyRH2NIVqufshBzzXDGodJ9ie+RS/IgFYNrak+bphWp7Dd3Gl5JBXH
jaXNgHOSvomPEEedsOMnKuYTTQ7vGTk+fni5ojMA2hNXNd5umtJWcCRSFRkcCebo
VlhTX/pJTvlKh/P3L2HXlpMgajRIHU52ka7690NLblbiOwqu7xPzLKvRl16TdGab
0TcMxJazzmgzXwVRJEIZKYxvfsDwwHB0sFJAHn3mMhcbu9zins0FEZu7yWeZ5+qD
nYKWIWMaS+m6FYqqPo0655KgaE35lB0hvPQZ6JJNmWIkuKhJ5g7jge0QisxbaUJI
JFEhsUba4xsMVrogDBzm1MxWkJ+783FhjsLQTHH9BunUOtwQH3aBG6RMUcds8HYd
VQ9aSRnK0VFcMaR3nL2FAc6ewq9LxqeQuUTbfMcNnD9iyJ8ztJVdHsn2YaJ1YEhX
U3XXGZWpR3k3KZigbfICy4OySOcyI5UZtJ8a9HSCnxmUzxVAT1wY7CxKq21jvQ0u
fLHCJoneyiMZrErwUyjOzHiAGuthCgcfrRrgQToA4LaKvvty9kr/528g7Gem/BbU
zqy6JVO5w9/Jr0qoftg9TEJWHhbMkY1FKjmJPcP1V3SKzUjDtgUCYg8va18WVtVj
2arrYfsFYg+QtLN/lZKC2/YkkkbqllU1pSXVQXYGGjRTPAzHrr4YcOTMJR0CU5za
UPhls1ZVSOxI4reoEO/U7jfczYp5SdbZOfUxOgM79L80xw6T3lZBN7/yT/L1jbV5
f8EufM82CLororVRFW9vUwUtc7P2EW24YAnGdM5hxFduubGddba75MsmCuXoQfB0
XMNKhqixvIZ/iNiiIKqBBoS78BMDSVDYWdkW3qwxkjPkmq90blo819a5fqKWkkq2
HgQ/U693vVxU6fV5vwOvegpW/Y5SosTlUTq+BNzHJaDVrjDKHyDUmiHSMJy0AXLe
ZHYpIhMVGgh/rbsErtaIZBrUI3gu3lrufRNx8zzTu5c54WjDXKxjZYGllzg/LQro
ShfhNw8wY1hohD9xM6kXOHlSbVxlqQAmqBJWIOvVZrFPmJDyobncwGjCuekrgtkg
/bWouKUAUfbS952v/6PXpXc4EIuUTZIghLSyUxJnYn1PxEvGyy8Tua64chXNV0/h
iYSrP/S4s77pjgRxQsxx70P483874PHojCSlGYpWCTCmM9gLG4T+eqDJh7QUZs0d
mwcSpdd1nJRf47G16Xrw82rg8IGJF1wE9ZUMfc+bSmgbhCXnsd0+fLdVVxS61gnf
XRRlpHpx4DjaZeHIKJQIARjBrJJtZ710+no0HPYUJxk69T3ldqrJ0bbcR/vzHh+D
y1kgNrvz3WrJpZg2lvnP3xl7+gjy9LK/ChOUqdLpxPjERmMMiCb4cZyh5MjUp3UP
Wy/+aPxF0W8dnQt9376Stczm59usBFd1PIkcMVmrDpHna5bDdhTlR72exO8xA0qD
syoFHfkxeP/+4mJ/GKFIE2BTBt9dZSxolawg/o8+I9JgAmu1J2oz4XmXI3MnrtJg
WNVm2ygYgwFnNs6dnvnv172+A0JDdecIblSF8drml7DsgDSbN9zqVtcVVSszomXD
xZyv5xLeM2nNF3xmfdtSw2Bj2PibtL9OXhYk/l2eotz6itRkOSdWHle3Crk0v2nT
2xCMMjpTq4mCyqqvv8XHn2Pa5nmGGwuXuaGSvo743uIW9PwvgWWWP3APoTZqBVKt
NfXkMk4tBPDyv8r7fHs7/7W1M7HDMgxgaYhXeSC4Fq388JmtQimEcaOXw22/tFub
gSM3Ihp4HrNHYviiNk2SokPxMr9VhnSoFSclUzss4BoGeEa4mnBxEcExtHe5osdn
xUSSqLPxwdwrsM8wesLzWMJWI5/NfrWkdmQ8tM4KCb5E91xOcFvsRAzvImkoVof5
cyswZI4SfrtZISlk3djSR99apvNtHwSshOXEGw0cKK1/o5E3J0fmaWZZaZrpxuQx
W3vgL3SlDkVE0NOQh7p1+o+xHDWedaDSKSkvrpcWEA3ltx5RhZlW9eHvPSYs7SBT
MG3iEWZBQNYKiIc0yHYIjFhEQt/pC2E+u51kdKfTDHOywZDQEo2AJ7gST6N0p9VU
Bfa60CsBYnWFOPtesrne8SldInFAhZ+y57fWV6VTie9FMCWgOSeh1KliuvDIQru+
2BZIKXjyjQYjvTk5yDGYqT2Xh0GXi+xPklFX4KEuhqN6uYa+BM9Kjk7HGbmdG6pP
4MtGvV+E/KGWX8lwnEiiL3SLM8phxlhjF0X2C8fDfqdUQfd84Xskzoke3Y1DUe0a
71TqKqgiEMQV9vCTpR7zRtoqH3lJTo9i7LS9UxXFcGpNe1cdILbWp+SjQKGfi5Jh
XXHPMiknWecshEpW0Jyc0zseqlsC0J0l5Bqm2J/L3InWjqe5veX/rH0CvwtKXrbX
bJYprNOgJK8ipkeDsiwAtss7MI7aVom8BT9vHYI56JSkAQtYEwjUQWEtJNueXqaQ
xYgh8+WiowUwHPOUHIdPFg5rKEYZnD0kB8E6wwa7ZdfpWnih3yirG4R1TMJDzN1Y
A/olM9itpbsYr4pBVze5p+G1k+9CKNxPcngRl3czZ1kaFLt6+BtTLFw3WH7oUiNB
vjjeRxLNWODPp463VKtHyvdi2c2BZfJBjEuESihQfzB1F9czxiWrTpEE+y05udUh
HENGg5U0titedpWiJF6TmQyvc6zKu66YRJWAwxEpmuJXQpNqYcFV4c4ecuVaHM7r
/3S5MJj5jo0m8XeKdSUONQLA2S2wZ8aCRxHI1Ed3HXRq8XKud7eboMUNqyF6SR0O
96cutpiPul8M0mxuHC1pkFn5DJXurxC7PV+XI0jNQdmn5fXpjM5anbktQe/jEfdV
fxTEoQf9Rp2IU21OWdZv7CPP+VgoIdOLPhrhgQDbw/tLH5SvilUHM8Gd4zkUJQue
l9uh/c3Ju07DU2NkzSk2E3eyl+DCiyDu/kXY7WspebuTeDSsVruyzUDAwXvw7MZK
ns/I1898XusFlF0NPQOcFYeapJws2QWv+e+u5qFtWbcwdOP3YiIgf81E6SL8RQ/K
0fIZP98TUBnRnTPqGLNtn0bnJN0EvcFE2LRQSqlimUKPhivyFHHMR7rPHwcW8TXt
JxXFf9tgQu/vxOlvYcjkAg7Y16ZsFkuHZzYTy9fBcUw70mWHiggP/4tE4VnZYfTn
V1S8tAX6HUOcaTvnS6U5T372iOgwGQppAvkCpt3sNMoiUrhWkz2YNj2Ca/1sMWun
zkCK+fO5Y7/3yeWq7xZqDKeOQxCY4tWWnyTxgeyomtj+r34Ji2hpRpufgig9OJt1
OswHTYsxjwKhYIrVTZTC3aMLLz9lOe+QvRqP9j/CRPJjjp1OgIq07agQb1Gjo8kb
7eI5mqHvbZiSghlk88uUDLePvE2Sb7JPXXKCbZPOcySozo7X61ZtDYovewifru53
oPzkx5erG2hwDwRPNj7+5kya2rrU8NKfj/JMGmHPgbMgENYdJ4YudI2rOMXGSNAG
WjBz/ErCISkB1Pws62COKB/Ppcw9yvjlDIfPwlqe1FGl9v1KZjgA2wEOGIdjPt9z
qcBGKeEDAf4rOIPuOavEb8dpfzy0FWdm+Ls2MBdhCxE1gGNMS59nBU7PwqjcKPFI
/US6NStE5zScEwPQYuHu9r3mTnSPuNm8bMY8hPDrIl00Je4SNdXUH9635WMiLk59
mjFSYVstImxK+pzJC5Wz1Jrx4bl8PXm7NfIerPaukV0qJpJECx02YzUnJvltQh4H
t+QjjivTH415/iQWvR0fvpEixxD4Ma7bqgF3URMG3lo/Q/53lAqfSk7n8mpuDzG6
N622+zFQ6YQ8u11RGcAximzDJwvmn6I8Q7NWFK5iGlpaZm/wFoxR4HKcgxSkANmz
UKYn5DMuuyZrCL6ft6iKxPDYuZycjJnoZmw4h6NpSFCI+vaDuRRGOML8Hu0bF+Ek
crhDXnmMbsNOKmKRVLVhXLt854ITTLIMk2Hg1VoGKoweyz43+AEfAQCD5wrUKdOG
cs8+hOx54eMQ4Dz4kHlC0I+vaZfWkvjXVD6uU8IhYrQMyhUOhVClYKtAZl2cXFdN
GSevVY0N6Y6h1OSRpjoiczhKMOyIr9Sd4JL0OqqHcDZM6/dRq+MerakxA76SJt5Z
LU0bSD8Y31mhhWmM/oT9qtJbwP8q2n6HKNojLD/Vkw7LtiiUE+ZCYihIavRZIbTo
ebjoyFwNBCXXBtpyLYSE+abDHjGs5Pp34V8pA/jrMjNjGhB8QRvYm40IrWu9F4oh
7xiotYs5bgHUMamdOUCEW5n5cqAeSdIBeUTrkFVXJ/gzKSA4HA+mUhOsIEwuaNHI
dTa++GXjhDELou9BDPv9wn8ueSGNT1ZIryEQDffGnx6En88WhOwy0YOa9yQBx/of
1TKR5xnS3aHgGbntcm8RwK5Xlb3omGOP6qCEe0heOQ3iwrK6JRDrR56yjQFguZ+J
0MZwmDWvtWGyfppuolb42HDqmC1+DU1vqqPRdUx6DxmvCUWkjZcEt7KV/tDKFMrj
j1NMWYoo1hnF2rC7PNuszulQ5ksJ9hudB/3yg+SZTQggZnZMRMU2i7f98LDbj2kh
B9wUK2YpsxpjRmOuX1SJuHBNu2LgLSQh5Hgt4oCZXUEDr7kpgaGt2DA5AIdrexGo
gu8JlCug0qCXcDMA+2eXDSw5wCpjx2ct2oAZmSf0u99KHpIYSWljCWqAHPVZc/4D
MFjBD9Zg1Lh+8eI0NzmwpaWqtD+IBZCRQ5O3onaWc6bMQwl3hLfEK7kAo5hOrEEF
JJkhiSQjctMtxTbcNPijVwqVpS1KkfpYs4LVN6D1gFTGi/RsB9AEiG1/0OHZp+SP
t0weHhnjqnQ2YAVCoCiXbNzqui8u5LX3cFfW5USmnFd4tZJz0hfUgsVbo2w9lz55
7KepH12PeN5rAxcGKS/r9nmiSzY1gm6f2RxSrGvarLrdg3CFq9S6Y/Pwoy3ypMPV
eXmfw1uncz5oKRd1hIrv2JGh1CwwBPxsiEY0YTIYlvfSA3paMeHJNuqw7T3Yhc5R
3ajTsZYsGA3dVMezGDWvDPs8IVcSicpbxmLwujiS874HW2vu0+89/QtRHCnBae/5
UsBXTLe7T/rzcIp8PU7A1espNpbC9PoOCww/TvbBoyN1Il3uyN+ZsyAjdln1Qyu0
2cyA99w5VZBnXd7/4UAZPB18Bl7JuvGObvh5rHB7rWi0H7nO7OtBDVynIxerxLIo
zGCbWxYIy0SA9XSka5falBW8/a4fZJJr66752HLgaxNX6Qxduk+1UFfDAki8fG9g
QC/ioFuy+Fl0nMtx7i9yfmbq4A67YBeV1EZ7/sQbU8KnKWYjCPRG7mdcQAO2sjjs
l1ll9BLYQAyFmO+GpYIfgiywS4g/yECQ/9T+IXGszT83Pg/PlrMSV01n5L/EZRuM
yADtCKKWARiMP3XCU9GQXWKQB/o1gQMS5lO/kG/tLa84MViFruz9ldctWgYCqMSC
fVEMh5f/bGmsn1ejOEWuygO0OLI83T/rv62G0RWDfgkgwOH6VHX4DD86h6BSrCiL
+A9eibVKLieS/EH3CbXs1GPQiRZ6vGMiuo9abNB/DhQc4N63B0wG9t91CiRNzGt/
JAWNP+h3Dtgsk+FlTBEfOQZfEVHIsGP8Nn4ig3kouyOUCuxwSOhoUgYehasN6zgm
MGOw/eKF1gV3sazLpUPYV+c1qgsZK4mkU/LKzskQoGFZcfLOOZgI2cddFN3m+mfj
++QY6NIoyVSbRdJF0cg88hf99J5SK8Qo8Fz2HoCHSSvcp3h1KAATDpBMINFoO9JS
ad/9sY+H+3N72vnsRv9VngHLMM/yj+gHJEaM5Grmyd0mPocZyfUUadrE51OZLG6F
XHa4hQHaygDUN+BgtzJyUcPqHMAr+uu6V3Fq7BwVx7TU4zwBrGoPIG6Shr60Eht0
5lmmLsBi/Ik0O9ulA7J5xpdUrAc1V+UdnIHwG4F8rjXlh2QxjaCsCstqPlo2nbqC
1y4ZB54gS4kvSPAw7KZFA6/GLtHw4/RUtSp8EBar0px3fFB1/49rfDFqlI8Yr23x
laLSS1uZGzgKUsPqGOespOvNLj5B7Dhckxe5eqtEukmand0IWcJo+1SwLJy0eSvg
QNEDTAQwaUkej8IuMNgDDBsUcSaUbQkSevxh77jhjzL0MzAvBoNAIUBgp3Oq9Cap
BKsQGhxZUOtxz4/yskOaGvL0Xa6ueJrY7LIAv2bgCwSpNOU1Pyr2tSEonIBWCHkr
CLDezC1gdNRKjnCDZgbLt4IW+Xu0RV8bReVrBJwtOb2XrrAZ/IlJ+q/TjmtFZbr7
Nalxu4ZJjtPg84gCJ1I8YaeorpJXJm69QrVQkHfP/vi9iTmmdZ+849lKclI2i3W4
14vGqR4uWtX/CH9H22gl6Z71m8CQL4lRFMBixgRw5Bowv1FDGltqdxdJc1QqZLMv
oexKRqn7dkGXvjpHkYEBaMr/QwnssnvFvYwG3bxIB6C1JtYvSdzg5CeExLEPzB9f
UzV0YvZNp+0miQvKZhTsRZWn6l6IYCV2F8/L03Z/DfKr7yN6CBghtSuE/To8my5G
uA+zWieZ4OwsP1eLbfyhGO32FMomNBl54xAcrzWED1jVB8s1NZN4IpEiqki8CPfB
rynuJw9/+iPED+ars5beUkqWFlIHqyS1O1kiBHc2uYJaj3oo4w2l0LInytbc4FoH
JmzAzXLKvHZHO5A9KeKGOcYeDAQig0yH9e7eePTgttq+wEcyP7e9Psv91P5VFYHu
zTEGc0Teh6UxD0WLRYdVNCcPxUc6nGAzFKmSOu7468Rq3s5roDM2v6rFwrjLOGch
27cxkFB4zQqwJGIddZjYeCEPQ10kMWo0TisVTdmlS79cMihRjg39awIcx+s6vPmU
chxr3rVuY6vwmCIexwgKN6S8XKqOElfY+eJkR/gKGO7QA69HFXW7o1GUfvYOOZad
07d6tIgiHYT7mXwrsYcXe72isn9W2zskf7Ei3ARTEf/l5djIRDpYy4Ra4gsCZ9M0
oe237kVQv/CpqJ3XPD4IFYr7rduoOQlJAzD9zV6maTS/1tsV0hRHGc0A9sbd7BJi
Tbaw5joN7Xq0yD6KFVPDdNcSm5reXo4FvGb7j4QMH/NNp5UXGJG4rtFJATcHnN84
a2mmhQ5C7mA0yJaCw5ut3p2jSxfLGMc3OvabLz//ohTc56cXNgGzHb2Jou0o81FM
IbR/kzmKGTE7fpY1evzcq3jerlfK9ChRbAlEnMGDLqmvwM9G4BqNYLLYHpqiG3pc
3YF4mCgZ74N1NWlAjuEM/W6iUryAFHVByg8WxyeB5FNi0vWpsr6ArBYdmq4bAUyU
tQaYLA5/w2bAu1DUBQFMwobnbpyNx4N+djHlt8cb+gSVn8ReFJhciVmP9Iu4e4KR
rFsIXtzbm0JXdSmKPDWZVvVw3IYrrZcgsZ4c5VxSgNvDtNIA+/Q0utf8JUrNcmOr
F3Lhh5+4rsF7tF+x3o++JKUDMScn3PaQCMHfNW+/yOZDTPvJaIXd/EkbBCzFaks9
4S9g+wDf2GP3utRF5FfKUOtDltAOx2Dv+WmSCaql+L/ZZoWn3NGN23ZtJ2g93VbB
hL1Spr6Lh3puJWSgtlbkZYmNYENOmb7C/UGYhpcF81LFd2u/w1PqU1MwVDD2weVx
3PH3VFGw7kZkSsnm7FyoY39C+qKdlNKNOfzXJTavAEUyiYUkuyuonc8SrzM+HpOi
1lHfH1cxZDcVyXZBp7agarjwLXK6X9fYVpWYaq/+Oe+kv2RgLAzPQ+pwswvAGyq4
NJLhZQQltXWGfH339JHlSWy182L0e63iJY0gDORxUotOrVLzA1lYIX01L6bjCkBU
XtPqnJt4XBZZqdZeg5vDdU7A6NQqa8KXuKLIfB5alSSspJG0MFV2JG9QWtsIFat+
nmWYKo2hhMGmpjyF6RXYalQLGT1KuHiNc47wGMSWWeraCLolkrwOMt/wqnMco6BX
f6x9kNvPsA6tuFqO+seTqGSdNdMtfqDFpdjF0+PpCR3Jq7TF2BhG91z4tw5AC6mO
W9r2k1+Q9sjW3aEZPUXeKN+32ylj4+SdjYxN2wG332cm61bvYg6ID909O0bRqq/b
7yYWG6j/oUHsxfwcDu5iMD8XK9PXtsWe5+Ycx3YPLdllP/yCeJ1k1E7QoHdZV3LR
dMgAqDlRsJ22vsN4UO2OpxhJ5zEUF8oiM/I2p651LOKnaz6wlVuNFUHybdyLE2p6
pD4qlES0bV6kOQdFKBSiSm1VU+WLOlN3lLmnkPeIG+PKb69+QbysfjCBSMJ7fNH1
icckMPD5ZHoCcELdiQoih9tjsqFsNE/DEteNTfzW3ijrnMEx3uTd/SyhVE/jc946
WCDdWpN37hs9S+wiqlba+PMUtd3F+1JQuBk4ZemkdhPDrKMJTiyR1UOTaycRty+Q
V8LsLwGBURwUdpsggDKihlU9IMsLIQdcwCZLvF+mW9LsfkKyerjnm+vqH59btUUz
ux7ncNqOlwNXOfUNFXl5O6Jpml07swNdyrw5By/Gr00d2Kighkkf5Ol8qR+/GLbt
cgVLjUNiNDHa50IPbdgqyvhzmlQ9nVOxDpNl6LO4n2bSLP1VutVhun5JyAVRsOHK
Q4D8Gfpx9At+p9SnWuNeWJSXT7uVScjHOgnR5QlqICis3xDF1xKrpeiNIBRZJLOw
puGRccsJRc0sg+ohip8hfuuXC0wE2dfUBVnLl9pA+OUzcCzMysxBkGLViHbZwqWg
S9/PeYJUoDGA8JUws3hdKlAZi5DgDlEDL4QUHb+AtBXS/bUu4Xr77guoUt3BcTjF
OMBzETCLM4WdnJ9QrWJ5eGm155O1wW0Kyz1+S4mxs8VGpjcrW1no3+aJSGTUltvq
16szLWBLJn7D7aHZ6ZPvj2PFQSyWHDVdmyuYem3rEo8Yd2qUv3qQe4PWy8RQQzoA
H+uiHb4V7jf+2bhyyZyjmT57YuYztVLA4ov7sqNVYhjaVaxGpDBNa+mTDIFhKFbw
d/e2hNoJculzja2/OeDboPcZGi/iFY/GROUqQjNkK6omGJ+L2zHDSzsW7Dg6JkCU
p7Xb6Pu8rTkkr0FpSelsSNXqa1V3Gd0tu8H6XmYmu6K0VfBg48SRMDP3YV9SUFnS
LSUKl1+3UmzCSkEjBHx1bpjAxFURRrI02v5xmvP2kAc6iwYB+gXyq72ZNMr2mVo2
vlfJZwy0/3cwlpRLoS3+xjhYc66vsJQlXvh45wojiHM//yLac13srLPo3D+5Dxwo
Gy3a/z+z65gaef3EN2vABnjgsGTqbBZJs/k/FHGrYfuzJ/tZiS96oJFQfLOcbnSL
hbtu0etHamD7/Dt+mG9HN/ZiGh87Mptu7hn6bUcsZ7+ICgCuxXUgmRMWVrSxlS+R
wytf/ypck79zsBzEEHhZanPQwaLNqzvx70dVdisvEZnd2rzLQtyev0y2wRPg3FZ+
sSOS0BKE1ZFIg6Fy1ElXKsxYvT7kHImi/ChgsJVWeBN1rEslI4RkqhJ96KQy2cAq
YLRpHR0t/o6pdFkwvIVXhcqn5INPNBIFBx6zwcMEZicE5dJp3bj6YLd5grMn0A/m
26OlBpw8qmsuH2zWfJ9a5TEkta2N3tM1k9FYFXoWVqrDbTPic9Uapn2aWCHQPqIP
xPFtDIqvYmdWBA7/WvyaQqsjtdWj+yU8coe49Sw3+UH4eTEk/QQR9aGjDVlYBZlp
DfyY+eEJRzmfcQuceMdXhpe56d3bmf+GohmJ9cwcKaoCPDQeejeAFdcoqJ3zYe7Q
E+3Gx+7KPfHU+T3Lzo9Loyi2INBb1lN1StHy3wqe97uKZHCgsOSJW5AN6d9sW7vg
sW342QK+ewfG7vrO59xG2d4ekId0UtTZKPq3QIGPky4r02ZnkQF8t7N8eKo0WOng
82ohFSpHDVxJ/AjtrdtQ8U2rIVw3QND1qmW3hDVQk3C04zwnenXufb2cHYIRdrGk
Si9hU7TjHxZ+NiLMF+BFm+KISdb4+P0H7cIa/+RbnMStgDnZkHStYWzfxkLLNsjt
K8OqRP8IdYH+XNAhlLD6RQiqECflE6INrm1tFb6HM6NL1lGQGxAWGXHaS22OEl4E
pFvnaM/OF+3kRwx86SW9R69PKpljVif8Pc5b/o9Rkne3PtRIo1EB0dRRrFYpCcv3
lqHjMCMmBk/5f3nDC+HHEpESdxP5MtA89bY7aTmPMGO2zmbjlp7aab3/+ZcrdRrL
7rWiT4TOxqZEUTygf0jsxwZ4ySNkzp9PTS9izYkdJiOVBWz/kZGcEI/AFYuUJFIz
nocLpXp4y3ZtzpL8jVXDn43NaDN3Ah7ggOJTwqgdsL2UtVd3qflNFXS0e7nui/q5
zWT+ujcUXpyv8iqCY/p66V7f8Ur3YgGsfDhLCJIYIU1l38MYGy+42Zxn0PgqYea+
WF+HdTxUknrCN6MW6FRUXbrqGTQDI6EKkk0aMIcTRRp+5az/3mddu+0dTCmSngZ9
O9FrgKOerdkm4ooVMKctYYqA/YR4JJPPTgJPGhzQpfoqbuL6RdMPtNaXy76/e4d6
R1Z5T1fBCR3CYTybTO2pP2mz+uUyv1E5UC9CA5ArgPMAJJiNX5z6lQm4ag3FZAw9
t0vZoG2R5Blq8Ewu88ABgiqiftugV1kmyxqVPj7FwbVvC48Pfm32dWRKCBeTgX8y
XU2LPi/Df60V5/4cpqb4uv+Kh+wvTNOZ8V+eGTsmgnVDU0Y8a3U/ZxoP0w9OT1Tz
uloonF0DQM5SLUbN9EgOmz79ctwRdFOGpD1nA0BS93xhEVVMGdCfSgWjIdHTCjYY
H5lUypAkDBSDJ5H+Nl7b9HTLPehZXQp6R/QWp0kNiOrxpJuORVPRE/rbVEX6oT4s
EMZwdYjz0uuKyvZzAK8dqgMw5GFUt1BL+n1RwfLWUPOkV+uzWOywdIr1r3sBmkGY
mwxp83DYaVCrjclCrSai4T85r+uswFKvvipmfOdfSDDCw8FZWk9b3eSNX5HcjYpi
YKkMEtnEC2pD+KaXOZksR2/vMdO01UjUijzrwX3GYG1+vV0CZzFZIe62bqFDicKg
5Vg1eK5yuMTJQ3U/tX98hH2YI30NQsUYC794l4yItiMQIUyw+CrJ25PhZ0fxBYjY
h4cpZUDuZoPwAEmuwOpBtEaX0nMwhkYNmbjz8cbuoKdkqiJ/8iowdyefWni6ghzf
1EBZ0xtwAbRNqtTw99qe48TDtpSkkQ1m7uQ7RaTXUQHOY9qbEyPCu6yF6XNkVbIN
mRESQ1nfaeUZf0FYbLwSk129W/yFlsDBbZc5jffNQNNbZQg9qWC7BRR/ZaPDWcV9
L0C55gpF4SLm1fhJOeguQqj8CusZliXD07mfNM794Z9Vre2LR8GiXynmxEUQ04Un
+HnhZHMUAma+aRDtDHV6CBIC4Stser/qEGrlxf79pSliHiaIt9nGkqVsB3QYd02g
/WZh+lMZnetm3OR/XWetw4K32J9J2Rrx1tzvhFepGtdmVWFxz2uSTRSIP9I/OXvD
wfJ6cBuI26UoWGyWkX1AwcRMe4Bg4Jp0OEZrhOjb972LZhwPiV7cTa/NfU6RQBkN
gyjRQc4jGeIYnF5qBHD9nRLpB1OAb4uVCYMZFD+fjyhtrOsY+ttr4tsjj9ftygoj
kLceqgbikXB+gbs+qV5Ho1rZMuQ7ejikjTvQ1F2SCDh2es6z81CkoLuAIbRWYP78
ATL+lOkoTPbfJP7SZXywXUjAzNaxYJAS8eJtmbt46B7xiWGzSJiF+D/7PfWo2CdQ
xULVhLoTsGgpu/rMAqlPQzP4+iL/WON5m3OczjmvtI1vlfN+bX+fflJotIAnaAHG
Uhsxa4p4jUzWRnIBX+1ogYdYtq1Bbf1ig1PNeEDOZZpWlqe+D5yEf3IgUeYLKHs6
KylqZFRIlNKrkay6n2a51Lko7kv630tskbnBmhmIDYPzM08aXgCn45o6un4Cqlzi
dqdYsLbKdzwWikjSvBvCGimNc1Les0MXGW949tTFA5G3UIPANelddGZTilvd4pgN
nDTR4SMxyXxr7g5oc9MubGRyJaiObzage3roTD6qDjKHo2R0UFvMYH2cqYMkyVO5
vL1+qAyQWAhMYVokGTBBS7dF6PreOWI8xq3puZgWsO+FFf0K/nqcRCE+Pv95qr2f
vNBv88SVxCFg6/HEAbF0ism6Tc1rQ/wzuxEJt9RzNtggh/UtaJDxC0vhLFPGmxbJ
zroo+pIGHUri8LhvanxkTezkoMna2SwKR02wNzqwujW4yJbNv+odVYTH0xqrL6mu
NU7t4uZv39LCSjN30ydy/YZtNea9+yFuqlBVsS2onBsJdN7yXlR91Ehk3Oj59Nb3
7re1QioaL7Kr3GBGB0WjaIGvxoyAa4VyUgOnhPt9KTWI4fhZXR2idZL1kke8pMdL
A6sGNJAs1Wq9+brHf+ildOFbm8RzEGYNdHjUkVYD4ATSKmv0u3lxV+cjAdDAtwEM
VMAdBFxR2yeo1Kni/YQB4lIwIlo4iyR+pB32vrwUpxIhNNymIBstXCB2eIYqZVOM
BFFJKll5wJ4efal3+yDA0sAQ+STu6ZuH/oE8zTU+AzbauQH9IqfKVJhX0YHjltJt
MVkruyX0ZbzDQLpVbAtBlfwOAk7B429L4GIuWDl9QS4uXpz1vDsBKcbNJT8ZjCzM
yosSIxirwXgqx8uX1ni8Xg8ihoVvXjI0Y6E0HnU3cGizRRi2AITEvIqTfJwq8TwG
jMFVAeVreVLgSySZ5VfcgqxsiFjPwJI/zrx/G0M1p7/HkGU8JRQiVhtQLIxKXyU6
kbMlZl1gwMhm/gX7WpWZu/kJdbAEWUQSy6MQ/p324tRhKfQB2Nn424mKKrlYnqq/
mNwMhJ9oDE5N2CWHUq5x+pWoHxuZMB+nGWz310TGWkAYwPl6RnZmkAB5DfGBEAM2
20cMfEjMMavzYTDGDqEsReVDhcb7NS5JribJrKNZ1GuFK5p0ANNjgzmOtumh6aaw
8ovwkT23/SnogtgQjP8X83LPeuQ66mxqsWnC79H5gYWJpoSSFtjk9x1VYA2jPESI
7spYijQyiLnhj0h6RmByxsAaGCQzAoackMrakhyRWc52ufz2Q9FkrCXusWJiWFlf
IDPOpCpJRCBXmEcp2D0fUiBcw1KXGWwDuwWwQl0rJlKaGFG4fe64VleRDuCKUf7e
EYy3ljx/GYTVEDoXhlz2yLwAQvgFpQTpiVUGF5TqSFjL1TmssVvlZ3Nx9TmpIQej
enCGS7s+oEcNPvHJN+NlCS3zrSlfFL95W4Qz9v4h/zG6hjZ3uzOb09Q6oA54Kef7
p4xEDCWuavE8Sko6qCggBoAFVfNOVVxS0V5f5Jipk6njqUFS+mhmGQttK2gVBhCA
/WhqdoNgdeo8q0x+SnFRcUM2c33J/kiS7YkzRwziqpTbwGyOTdUx5Cz+wDR9fTA1
+XPb4E1Uj3FDM8fJWTaIWYc5o3I6ufdDYBArwAjZ93sneT8YK3+o5+Q51a99Ix1/
Kk8XvXMvKnnj5TWossLsDwfRwubPQlp9Pce4cjz3MgLtTVWrzHSgVPH+4w3wzT0f
UpVHz+UOMum3A41ptAvQ16rkGaxhuvEFeigAfdzFcwZHLP5OHWuXtsMGfcnDQq43
kTTysQAhbn4vWXPL3qQF+g5JHw8VO7+zVyjoFcPs6GSG1yPjW9x5WU2n3YpJKTvn
wW09sGCIDFFo17BtVcdxEZLgQvFbiqznqrlq2WJWU/kOqI88RQbsoIWvFf1qTYmb
ZyVLL99uCS0R3IWmjLGyErstNx+/TJluyS/27hjLRpUqyeY79Z0sq6AtUV/Wjiij
hNKZKRSHCSmcp/qb5b56hGeT34k6quKMNSZZhpQqsikMbsCdrp8eIjAdAj13Zs4j
v0knf0gmub2JpLMR1R/gtQyAkxpNnvUySmhWiMRC31sOcG8+Tp7Qnr+heYDAJ3q4
0eV+2ugkcCbVDRw4Tz4VBrIkFXUn+L2aumEibvzLLpB/L+CzrHtBkzJzJTcXTZq5
tZGNPn7aLRotLKEzgMT9dDHXK3tXJ56b0uAiryw/Dv0AK1qj0+4uU/sQLMRPMN8y
RI38vchDIaMwDIdrumP9Zbb6yCgNoBApVqR+erABZ5LBsXdTKv+AD6bwWBbGpIWi
5FyGn9APUwamfcj/6ZCWDMbhlSHjddtbSQOdHIUXJPpP24t4ryf70QYIfZTSSHC+
+2nkwXMy5l3GRYsH7zBAYmdtjyu8rlyzT6vmcYBUYrzYx+imMQSmQ/RxsityJAnC
T+7Dh4YdYVIyKmmN1trF1TAWeOE1NX5FKrddDbVyBOPKnll9hPhuo197cBMCHggA
+2xAzHEtBqgvgnnya9qhpoa8Z4HdzBz2JIIKBgshHUHx0DMcaMIhhN1zWdd8toW/
4P+bOMioxMnDmOVXLyhyKtHzYsrOI6ftn8Y1YwUnSeSvNZm6t49hbycn12ZboHdD
3OwqnPjLFvhIfxpGYiLgsdUA65CpqTNsgN0nEfX38B3460zfKEp394Kg1KpvhF47
k4zqpkBL4US9ecFVnjmChIQBzebaWhwXxljY3sUxqd2a4xHse0XpCZIjfUN+Gryy
KmmO9WGmfBRH6sBPXroO5fah+1GgGH3kHn/pkdKkKWk0UEti+J4XOcuMFI3B76Ua
Htbmhxw61ximxH2ZLlYCXP9Kj9iCNV9dXtEU0hnhDQqWP3TJK+xtz/VfkmqNB9gf
2PvvCAbLldDpvGHH2FZIoz8C6Jsa7IsQTcKR6rB4AWm7lJUrmTPodJK/uIvvW4DE
G94kXZ6qkkIakLo2yc5YWZZc07yo+LtB0Qg67zHPRWsJbp8e8MP2rSoYFfLxIieW
PR5Mza79wm3QSnxhzE6P0uSJcCIs7XaL9cYrDoFuX9m1VQ3uRJNSv5O1UUF+gc9g
WS0QTQJuvCexmhQlX/PkekbnRIrKfD2NaOOR4dLsCM8sKWomb37YUUHrW+7cq2fC
EuAoMVuhMZn9jb5oAMgObu4tAU77g+ZIXQvTJEB+I008Ih/cVH+LPCE4VKCH5VPG
YdDOu13XRt0T2wdrRoMyRjg52plZLHnfDWK/mwrbq0PeyJAdJah+u1zIgeQdEdoj
lmL1SWaioFr0QsYZ44MauLIX0m0MbElLF7w6HFpHvuvpKxu/ItxpPs0wPkm7fh8B
5PeIy5aoEiG9TqYk8AMER2ueemyywOfLqMqHi3fODDdmye2oDx24Ud3EXek1eQTc
2gKgoKok6ysffs2yFqoQCDdgNE3H35+t0tYHL2uQs2vJ0dSg+OD282i7PWVO2HKw
aNPSJCRSTJMR55E5MLnbAaTljoKsFvvmUJx079xsRTrmzunGaj9Ib7l834meedBT
m+ZMPuvHEkxV2y5k7QhGH+qVLynBRERd234VmskjN2QbsR9JkVduf5yjH+dqcUvQ
Od8Nn9QugbhvVTO7BaNc+B3TUGZvbvmGF1oAF0q9gcTA0ZCM7NbCG4PaVORK+y+h
/vL0aYF1S41dKn/ht94nON4wEtqkGBrrUHTklN3ZzwyKpRcaavlolzSRCj/xsx+i
a8Ky801p9+LXykyUiSK2juHe21ffQS/X0dfmQxJTi8QV98YH1eSWJAbwN//usI9Z
d9SpbtfX5lh5xjVObLVFEwPgM2PkeYtXZM9BIRYT39w1OzH3t677IqK2WfAhmOVK
Dxoi3Xf04qS57nLDK82v9jnuZjJaD79aJxeypSHsECEb+vBFzPHa0wiYEH4PSwmb
a+sI7Qx31NrHF5DsF6ojWVJuFmc5WjAv4zXxpfs91pvmj5iSsn7RPbZFdd7/6rEH
dUR8ID0T8AI5isRSnoH0O5Wx8ZyAfZ12c+TU82CE3aaYNcJAK59LOmlvClUPZz9x
z3aiLwC8PrsyMCbGS+nuzaGDIAE4Bu/0gjsWm++8iihyfLcP2qZpEBNnT+WLdu8M
2+sfQHRXY7sE1pjB74UDvqIdNof0ObYXkTt+caYXEzinBNhpVyXLuouYv/Qj5eQT
L7pNw0L5/YELRADwwNPpqL+fEtu/ytC51gf/4UkTdAQTXtNmXUdWk0tBpDG3jit3
zwz0WhZDEjTzAZy67FcUBU81aLtWRPw1Y9dL4qbTh+ss49zewyXfG8/DIMZAoUmF
QJNaQRK030rzluQPk1gV8zgqDKkDrGVgM3Frez8Ry+vPIAM9qb/O6eD7xAJ5bT4H
uCxDp/4Os13ZPoFApD1R5rnEqj+SdvoWd0Sqc7Gh3fdVVdzoV0xUk1rx2rVZMcQa
7NezZFwyn2NRsuVKxU9f/Xnpwb99Ot+pzBJQRlcomsyisBew6DqaD/KM6s+U/JvZ
gFoJ2hoTaZUl6aiKswxn86TiYl1uRo/Tb37pW8mKya2n3QlAdniO1PnxFIR9TzfW
OK6qtTe7mUIFWIWbD8HMO4439M7wace/ilPcZfXtn2qLmgWQuFKMs+FXj4LtaDox
KdJFsm5bAA6cTPLXlKpmJQBwtOO3CBp3RnoS2K23AxbCYKj1l51tyGxeMO0PSBXJ
BpIrkIaKeik8nzJm/K8P5cHtHwtW6FWxXKoCKTL6Rlu58HTGo8BvIdBmASsrIBzk
MV1VH7EgK/eH1/lybP2I7KYDnCgOkkyWRFuJwDMbjmbyzhGEIA9cP2s2VzGl7knl
PtaP05rhY0rGcYHw8SuUe53A5cJ5oqpvZuBz1QRGlin61phdAtbQJDqN2XgzyGds
E3pu5+CU7/aaISGOYvqi3c1TVrWxTKeHyqUU6LEIA3y9MjzUlSRpcbd9tHzxwHio
v/c/PWUI6G+gotkw906lycbvQfBq5i/yDmnQGt2D30ckTgKwGXRMmoTBg4X2QIho
CKtV1l2kSM0OhFb7uIDi8NyuW/vN9aBekiyQH7uSW4KYUtM0UgAlRDAAKgUMUqTO
Nt2IuiM8mqoOgkYafeeihPAGQwkmZrgBgCXxihjlQbQe+XUcWgfPZmmO88kG8vlJ
8JhaLAJ8DCGCtFMi96e2ZUoJk1qilJgfwcsIH3LS79u0cHdgZANyExTzpUnCyefI
GP+C1KPHhS8WmqhuHldDe485is29IZ87zVhaFb6wuZ7SMYE3Ze4s3534dbATAcro
5jggp4p+kThkviRF1DOvc82HhuXYfJqvVA7LPlCJvCkta3P+pv/XfutGDAiakWIv
p+72qn980jZ98SQLt5NV8F3oGq9bvKKhR9lkWjatgvXjmx/SK9G7VygSoUMa9YgU
R2ilwmA7Xa4EPMhQzkQs9IQaix+tL+RqdjhL3hvm+blWQAWuvyXi4WFRJkEy9+ww
6uwmsYAjsRriP4+5yQJ/vrAivyIAMl/5mU65Qn0zONvBhhYlC5CLKbhkMISCY8wK
C9biGezCSElxpwwQTmfjz21tqA6XzpzVeITE8n2JMdukEhmojjBZbzOC443uZpUg
0BzmOFs88HFXwXQHqTnIgbJBUaVvwf5SMcuEIdVFaQngiAkSajmdyBpQ9EItzVdW
zrCIotdhUXuy9+JVlcPSn3hK0sHZvPiXsf0ljuhFzuLJ0h1MdojWF/vqZQSl5edE
AN7+bdHPU+Hq9lcDFt3Sag7aDivNuG/L6qgo66LNvj3ovg0RwUZli3AFoNxhxBUC
G9XRDRMrdiTF34LL3LmjQhv4wBTUENzICSXK32nrSmuWlM9LtvrmsYL/KknOD8cb
Qbc+1pCCbN0Up7HfgbMo3SU7sB8HYvXWajHU3TBYaNlv/BOMjtizgs1ACFOY4zDs
Wo1l8Dn5RPSnsNPYrUgGQAZDvE1Z90pSzYbthHw2ZH4Y6xHGiFa3CX9RKokA8BPM
6CyeE1ETPn3LPPlB9h3STs+WattqFwo6qFuBIP8TUiVcPKzgvOZ8m1Y/3a1lPZyM
X9pi6FDEfgPOjyOFeWNtsdDJJhFFd6pd8Hq0JJnmrqYJS8pP27BLJqRRXACeuudh
RbIGl//uyfcVAzHvpLfKnpsbjntIKu8GjgI/fWJGPDLeXKW3l5vyw6YeuAxbR5qE
OTDJSVR5Sqwp/3H/y9QO1sNoU5lAhzlFFmnK4Qwkc8n27LelXPO8aUCpjqegedwy
pQbk8qWaNIX1+gJ0iJznR5RuKVWKqtzerf/BWfQWuPIeuM+UuB8bh6ReruFszmCR
beOk9dY8tWVA2Kqb2WH4X6kLUKdhbddDKLQE4NTe3b3FzLxyMDJNBvHfJRKah+0Z
3WpWxyQqdKYnzZ/CQl1LQ3OgT6pXpXo7BHf//1Js2+ORU2cOKIhGoSgZuqRx1apg
aOgM0NbE9IRTG3ev4XWxZsT5M8mp/SEvTodZare7E4CyVhQQMWzxR0HPXDTCboMT
A52lIrEmVJiJf4OVLgXwaWc1UhgABlkavUzJJnbrqhvcy6924gGfym8uP0lBA+V7
82hMEOhwQoVFiujYT+NnRGWjnh0oLeBAhMmqwWvFg58d/MEJMR6A95rM4Fazv6Wo
mTjFbe/gBLdMMkbyc0gPv1fGKXpbpbvBgdJ7EHrg1Lb8QLShQHe6hfJ1Ju5slC8/
n0FfVQwD23pAG5pWXmb4o00cBAt29f9Js2bmNSiflaxIDdET5sUg6J4G+K7vPjON
IypeG0OhrVH1d+72YWSbeoowyTJXEEB99cqmgF412qC1luhg+AjFkxUODxyrqBt0
bzfY5b3ZlJ48ibdNtzSWEhnRMrVTvWOTHt4h7ffkd8+y/+y9NgRJ4we8fLYtfBCO
YBY/l4/EUZiPXNMvKwnEnLW/Ac6ftVGkVkfKCCc+28k7an1d2kLqv6/NMD4x8yPe
pl3amt4U2tB0+d8ma99SeBvGh5te9GH7pjT4x9wLhfilng+RC32jRYWelp1bYgXw
1sPgf2Lbpjwa8tMXxKPEMrYn6IPmR66j+En45c9l8Gae1HY7VrlIa7hsLmW4tgQS
ifAUhOK5H0FHON2im1+5LZG3g4MWyaZ8netT9of2Y5zmJjPfJ+IlEbnlZF79b6xl
HB5KciMx4YhmjZn7P4sLi+8ftpXmiEbftQikU/P1Jt8Z23NPDO9Vp/9tfSSsK++x
ujUJ4XLRK78d6+MnRzzD30EmEEhIkZUgolnp+uYJACWK72Ggu0UcTl8ZWubysDrE
iMn9A10lBkLFYVQv4wtjwOx/JCZtZQXNHv3DG0aUQl1oyL9LmvS1XJa+Dub6C1pF
aepwi61RY0LNQfq5oWIozfCmIhOvuL7EBqTqHL3QDURbK9N+cPj4Y4RufVRZsWfc
yTe06FjSFvXfr7fHhnf9Vvf4MFX7NvCnhgMCYwivmRsOgBIMWgqBlMFmz6VukaXC
TeYnfPA4KVfIcP/gtdUAyzil6K4DQ5Hby7BjDU6aiOHb8xLibCBYvVyQ63VnQJtm
WfIWDebmpCFNcaFUDgzuWvRyK//X24p4O5lAn+0/8YS3nFtLFcUbBiOug7GMOR/q
94pYZcINXq64NqP5yoFXnSy7rBuiAul+BV/4SCbbr8gZ4jFyhnkVhmYEcJxWGRtL
qAJ4AmhYCuFIRKulCnBH/P0av9IX2I7Tks17rHDds6i6+psTSYxmmV7ut1EAtf9/
oygwSp+AmYqfU9suLFF+jCH+aMwC/B9cZlznZGmRjxqK/QXaENS4Wv10P1AYsA7j
mt+Dvq7CufqAUb/8U1aHTp3ir2pybMQ4nSBDf1i9YfPKoiwISRbbDIFUydpRBBGV
3Q4jAnN+mInfKTXGMpAsiLdDJLPF5Y/RVfUgtfXJcMjc9w1TxoMMS4Nt6g3Jgdsj
PMdVVbwdD74dCJb+6wsf54TjETSqurh4Q+T62OungKMQnrf6YjWBolyZPjCfViqw
074LIV84YmWOSznIEITqbrTpMRCT8/vESAfI+eqE/5lP6Oy1SGLV574G/nAHIIzA
aUvaac7PgLdB1jYF0GRvW11xI8aHP4wGyo+z8C825gsrleJk/oVdDfcq0YKGWrhd
VzMU8oKQtOefIZz8NEv8/D+sI9IigUCVBu8RAloHC9g65Mrma0xD/E0xn4kCdzDD
O6fX1xgxM67ECeE0N+xcBxmuH6A0ChZwyt3nYvBBnSfXAEj1Ih0tJARVIEHPSHWp
VkR7wvGFtyJueivLf+JKPSfZstHicUw9XangylSLMbrh2/S60kQ+98/LXlNvxpmm
9yoAOop1Et06xDyPRrfeaZDELzJdJ+57Bp1uJdd3fIM1qsi8Q2dK4SAMFoUpvRqJ
gtRR9bijl7J6VJhLnS48mCAvTWj1TcHr294Rl8HTkUC/tyOwGVfZaPyMHNy2aI43
laA2lZm9rZ+NONNT7j28DQDJC/OhlBclMkJPoZt4GsADt1wS+ffDf0bpw0g98u3K
Nq59dhfnoV5n52B2O/6Gsy2IBPcPnrGEp1WOxMPnTA94FKS/uZDmzyA3ES4S3a2A
sSrZIrr6g4A7un31iLqt5jNeDbb1cLmVTuuf0RgFq0TD/4dOa9mm1IXgtwB7cvCZ
x3xh2Sjm5VRIn8/JGW7oIiOgs6z/ooLDJmgq6/PeQgySPHHwPa+YN7nt8Z0uUIsZ
ZYjIMRXa/gmk4Cu2DNXu3SxvgrJiQlNpGoRe1uQz6vet7YDLkAUwJ+jfmtaKeg5Y
IrN56uxF0wDOgbY8lajH2UpGdI+E6iYqWLV+RsWD0HkSqg6V/shc7xQHPyKP8dHY
mGlhNFZFM1AOvQCrMLc4yXmxEULGvRlMD1cTD9FFLHkXIMOEJ5HFDrra0olSE/Ah
z7vNNSP9SzMpBwW+JYFOou5qmWz/658dlkqrndtPkIHKAEF8xf1VBuIfKetu68js
z03M7kOGdvQnr+BZ6a2uC6Bz/LRZ/akxu1emeZRfRNgHw2tzCR4v2hdNEeXiyKPf
lBwc4paHE2yxykRi4Lv7YcNbOY1z0qRACQQ1oFJTelHF+5tIWvw2Cd+Znm2wfM/+
ebpvP8//uFA/19oy/bivBHm+BPRzpwphFfjNBG8M3gojN+zDh2bG6lbUJY3wYtKr
4wrsdh8GES232yQfma0EAltJ3aUTjWYgD6BCI6xbPJCUsAQ8tqI3rTZoG5MOohGu
2Fc6h3gNOXkXW7AqOBcxWErOGcOiuKi0cp3REtDbBrxkimu4cC+mkHKf+DqQjwfm
6gzbW3hYZZxpsE2sZ5wKiW65SLyEQv04IpcVYJn7HD7ho+vwtWtvuGxrD3hRjOyV
f6MEGLp5C7TcRp6lwOaReHBbY8jdhjfWmgdzMmmQ0wGMt7lmx8zQ3t/V3AJ8raJw
lGDUy74ajCKtomm0jQPF82blArflQX32BnFrB6XCouNdLBQPot24L9XzVUqmmm1f
kajUtUXEKt3B3GMS1drdTVfzasc1JufNowBTBBUy0cCIpfj/ikUCJpQ0N9JL6EFQ
uxujKWXp2kAIWNTGE3HicCUqr/iXvxP08mbaC+8nmQkYCqwFQA8rSoEAOJvDg4sd
0nmJlVeJ6isnoJbTdc+/F90nwkXTKpz5E09cHYEajkcKU+w5zWYIvz9ipwSANJBN
HHW93pRzR3hLv3rl5BpAhJoo66lXEVxMDROxdG7ZinuDd3sh+XruyEe2uQpKYhjc
YRpHitKfFGZwbF4vhHtwauhOM+oI3LhvmmC1u4mr/Q8p9fGnI7Fde+FagVN8c0EP
9fB4YHKUITaGNIkoMRcchadeMddvr7T/pdfua5XTNkMP2sit9wH9HpgyuIokfyuI
zWYL93W+lhGmflMCe70UgZkMBy/ZDo9sjOfv6Om+stB31VVrOYM8wAkJFljeLqfh
KU3Zqo2t+w1gwiEKQ0Rcl3ZepogGuWDW5SphiM8h7Ka5i01kFIFkjXE/Bo6gZPJ+
AQKKWeYqlYzOrSNEeC9IRj6HKUdVvTP6QWCGawaaXJHJF51Tvdo4TweynggoitNo
5q3t0YHP252k44RGJq/TuYd1t3hTRprSUcNJFYWP0zh2nylouiXpQZQ3+PIoeYrz
EOFxSoTZoen5pEz3TsdqNYmLTUHNZpjDm2xKJnHgXFxxtUKCLI1VGX/4JWPXW3hv
A6dWd20uNY9kwNHsYz9AzjDZ2bnpmEScV7/DPlsCljUV43bSWWUvDjiUJpE8uqSi
DV+SdJ0KVyS+jUU1aCPjZUJirzaMspm/9kgKauVkXvAapzuYeAeloYVE/+JUoLh1
oLx1/9h6i9H17feTwZG9M0hfv69/ZB5lQvKaR8ECsHhyUWddc8/T5++DWqeIpvnQ
2iDQ65ymFS0OuMZVknYAqpAUjyhGwLd3Ax8qBPNkhIKqD1s+hJ211YJTzVYdLHfa
C8/IE+QQ5lNvGviCL3Ry0U1Njh99qSiIMFMoY76bnM8VLJbP4LB3MtibPZRSK39W
wjPqvw6wp/IkyEMr9yGRMdaPqZr7dyFp6UpUD8OX2K4Q3tDRl1iuZETLJQjoldoD
Ql52atLXYbLAqLFTKMwbB6+poUD0vSVQrq7BcZJrgM9j2Y3DGYdhxuLlN9HlNyeH
FCVZpmGxKb4W7qxxz50AUdYhUNqV4BpKKT6X+Hxe3tvjdn77SjyXFSxzJLhi/AbJ
KhMrXFtTTUY41EaxQaF2lHXGi/E9E6jYFw5z1/LvXSyjLT0Wllny8AEg6dLM1ob3
R0qPMDTI/9q71j9bzsV6CM7prYG5oa2i0fK2YBFoKB26D9TGu1GinN6RJUxpxBN+
rEIzLjWAGorLJy934npf0yyh7GuYLyDuLfx3W6OLnZrbbyS5kuJrl11Rqnsl8uH+
n4GtIzxBOzBLvroE/yVWaavTVDfYOY0RWj5PBaRST+Hy8c2VKR6sOJVME5V3w8zt
KFtcrzGrxP6cmoy+NCWRP9T5b+ntUvbw3wWZHxTl/Jdnv1g14ltx2jEjfInbEckU
fXZUiCeAGdHwkHZma/LibACKj3GEgDKu09mMcosTCyUJejkv4DgRSi1iiAHVIbJg
xb1ETGc0krPgTGL1RnmzgtIa9J9rug2hxXJ/G1OQWsFKVhpMInExVSSGECWHczOi
NDqdl6hRKIiJZPo3G5aV3bxE90LO5kXc5Fw6TGi28RTsRzTbV0OUZP2fs7XJ1JCQ
WnpwYykPh4eX1CMRYxltB/Zg0u7M37GWQDtmV75NimFmOrxsYjUnjOqAojy8ENq6
sYAKLKzaZ2rlMxa9RFubwECqtjBBJiX+xInP1SKT7Qk6H/irkDR5KfBzj6vP5JXU
OmbdweEDqgCG0Av6T0QHrsibHun86s0A3s1lmHqNAvKDFy6yKd9dvh6hnsCHC6fg
fgVyOKhF4cDRQzblgW38wDw3ET/cTVQb+TiOM4/oeevGcAemNJCHxo4z2BfJaj9R
xXJYC8nlSYv9FAzofy7nomvTXtDWOwdnqoF2AyX3FR4YjMHHVuzBoaBsQaDFlWZU
Vsrf3JQ68L+TIs3Ped93w0jwA1jE/7SDnRdVlVw/TcYvt96GqZuazGlkU7dg2ulc
o8JL7Yx8f7sLTFUPi76r5MSIc0eAtdPb8tv/ScjBj+v1bK3oCixJbATQBuhfANtT
ohXvrXbqD4nPgskXW7PkAcjub+TrD0qFi1283puTwBJdEIx0D73s7ZLSyXTlzvun
BY6PIa77rQN/Q/t1swdbUkmd39FfHp2za+imtKgVGYo690Ox/IzeJDSFiUICnuXm
AKHEf6BO/VXjvIrXbhkA4P8S6TycPlUrTmZliAzRDHXdIANtWRbDNB38kmMKCl7O
HbMVAs7/UBTeAWRX+6ATm6aVVRANMmj1Dyxqi/plBipCh3s4znP/6a+LsxXdpY5q
W/wGF8FLXAz6GxU9ZW6W4hprJvd9CjkWHHUWr4bG/HN8agC/rW7XnoJIuyyCq2RP
EepN4J+DWBXUXkAyVZ9LQtXeYsuiKyPXUFunga7SNE+0H2AMs3h99xfb6GQMpipv
1Tk50/oK3wxi48QZkAoncwI5ad7HAWC70qRpoWkrtsehxPtGg/bAv4n+TyGN6HPY
svpyzSPd0Zg6CwC/LKUKzL1z7v1nzU5i47Nov5SMvzJZ6jOoiifj3ZvEpszbk4nQ
INeSyJqpEpS5ramXEEulyFolJBnDTr9zlKHGT+Ex4bLZCfDq5bi8OaNngq5JSs4K
b+lMfEGiwh87DrQDNSvqxamJTakykh4FnSnfs9OOowIbvgF9IHVdByBlKp4IjSqe
QUq9tO5o/IS2dPozH2MNrR5Ohga7j02wCaJuDrHM1IsV2BAGY66ES7vmkq1ywRUs
EaH+6t9HI9btpFOIJOy34zL0IZsVDDMc1PtAX/w8UXBri1e32NAetLds7Vfg7BKF
LimHphACR77D+Lbl//ycZ2W5NVRX17VEdbHayYsb+5dQ5AqOTng5qL6OCuRbRWvJ
EilbabRYV58hsZfgoHIfVnk86hGZp89boW3a8xUxrTDJ4uLHv2BjTMKuxqqO+lct
1YwL67BWBOMnvh9FLXewsj3eSRxaqUrso8bJS1x1gTDTPVxYDYy0r7n3Du+JEpQA
7euNJhU0JiKW5SKdyYZSam3bih/9laHi14jqfw0Kp9ba40HLTWWLj81w84echHmJ
8DuzWHFzh03DmFQz3xCvGoYnVMRjz2RsPxzdgJG4FVPyldDRW2tkVTehEypRPDX2
L6pdU6qPSfTFyFqvTAIiSaWUaxyj4C9GXmppwCi98zlMn8jfn7BuRM8hLeK/02ru
xn164DnXDL0EE4SENmUfgn0sEryhFL0vMSmnfB4n2pMnOAq5Cl7iVRqnP6YSj0io
fbrM4+2i0AT+WnLchd1zTV1786QjkuyJmROgJe+b5e1SvlFDCnHIiL3IARmoV1/o
49l+JvgS5FSVarRJNKJStb0a6qnZUKXwQpm9p3q2YzZ0+9WKYd0ZrTqDZJQQIXAu
9gO30nQMrVolo2DlpbqV+Ezf9RwH0RrGugyqUl6G0+ZrYWk7jxfU/X/DWBL8dI9B
liaUCEo+dzbYkf1ReF70l2B3lE8X1tgRlSHiuAVa2XzEsbwM9+LS9xPrBKz0ceIw
CfJLgeq5TvHaFbhtIdW9ATCTxfGMOKjukTl4z3/hpt88TpIM4whjji2QyTt2nrur
IbdtrKtpP2jR/lZ5B/Rt6O2cQt0uY1LPG411Axxi7scuLjsvEsgbT5P2oEuRuo2P
LKluAm/N2iEYdBsvFyXLYclcFHzzv0E7HQrGQ3zEzg4UCIU4TZ7FkN5oHlhw3iyQ
vqWXtgpEPopgK38Xu+wOcq5L5nV8c/20ahhzLzVWqfdEdtNBuiMLip7e+v7O0PsG
HXA/FFqQgFHvCbpE+cplL3dHDDVKCq8JnT7zn0LFtU/kAJoikcPQny87UuCWPxq4
mYOk8eIBISVv69Hiy0JZrOsh5HHBSH1a5gJRahiQ3Jbd/N8k6tn1zvtxa1VQzFmr
1XsNZYuzbPCsqDlLpGr5jaNff7pJZ/6yiI45wpG8BIvtv81twLrhCpw2xyu/Vwsl
sf8ZS+BUO4ikvHelbuzd5nZE9poOn686myKSkpDQnRiRJvVonDZMlmqYciFtsdxU
FN3mSiqxCOcPLj0xXbF1QGDuhF4Kc0JiQDQG8vQhWsMbwuDNVHngvZRXS3cKbB/p
8sy88/2XHVG5bDMasBh4AYnV6dOj8MkC7ogN19gFKQUPeN4dJkmdovLXEqEy/+w4
bNSuXn5C1ErwVQ3lPgb4Wclk6z8wnWEPvUGgRxqBwJ6dDxstC9TR6F6eObvpa6hr
6Cjnm8PrLuwMqLKU/i5wde2PbZJZBCYHYxInhcxink9Hvsq1dsGggGL7Ic9+4ei8
knDpJysc37pRpb0BGtOPe1r4GeZKjp8P4HhEYnghTdkQnaq4FA/iLD1k/1KR8bxm
bvfs290zisHFD46newHR0ht42PCp8NVhloUr40AragrO39Ecx4rWITUYn+InGpOm
WSM1XvM0lmqoHn3q5t8x0uIJJvAw2VFze8DH+HWYTpB+9cDeyLFsQh+Z42Yzs1V/
+D+K5mg2R4RdxPWZMb/VlqXAKgKyEeb7j6zTqmXtK90GM3vBnO1tkaLwUqWpnYFR
N5HQ+K8oPCG+6wjdpNeNu8T7HeuIsJ1hiHTzzSqlWdRqAf4nV7Bua/UqB61D+kgn
OLLbG7xhHkwqbngAsZvSoIOF6+I3Qxkfm3RORHpV+BFQVpu5LdR3XtLM9DVFSsi9
qjm1FbWriX9PQ/g8Zfa6wlMZ9p6OlJIjfSJtP+k/nKydqMuIzViUFHzJ3gyqxH7z
guw0CwJ2I6DPO1J+wE8lbKZtkOQXR80rI7IGOOo4PBNmQtQoGbQQfxn3Do6j94BK
RNBp0e/3w/ZKnAVLP+z4xywZ75T2E+LX1axzY4Rm/BM1OSlsB4KoGlk+wd6TYzeL
a+bL3qZChJfERKfok2yrlcmz9bpWTOY0g0l1qwBLh9aXXMBiPVoRW4DKfxm2J7vh
LkilOVtLCrpCFdrC1diY3dT4tMwLwhfl+5/u+s2auPCyc3T2fIfX2WsuYEziCyg0
Gf01SxvIFFmDj9p5EuQBO8XBE7IpbEmI1djnAiUFnLv6l5jo9aZEEZGJ07VPQLS0
9RjWBgwPy64VSpo1kq5wjk47zMeZY5eH73BB192CfQIHHzYTMITeAVbANPuBBo4e
BR+siC8iavTw1f2cm1dh1Rr4aV8rFlYLLbbuxssy3Ph/qvAdTOjoJ3pH2C29XYf9
fCrOKtbthbWVqZAA6e0KVooTK10JY+SPpNB+9yfYKAV93WP7zw5JFM574FCJCu7g
JjrDG/vP9GVXckMc6hZvIvG39xO+UEEsTVGH9ay6sl+UdxpECzBaNSryIMBF+Dyz
cK4YggcZyMBTN2AX1bpaL3GQ3YboTOdvfdojDqYvLfrF72J3+PAaiBBlQx4d1Gjg
wN2h0XzRxROnGRRnRjPKx3i9u4B0iXYyHW8IoKaLMjYw6U5ghOgX1RUWpwxUNoKW
JFxmgFEAlTF9yEhGaSN/1XTJPndwv6vHXit0C7pF+gXB3fZPur0jwLMMdRMaS7Hw
HkApa1A9N1ZKx7krTZiDRDk0pfuT+CWZ9vei4ejfWvYqsk04p4p1GB6qDGZdvyhQ
YxEh9zlW71J4IKK5J8Coso/RFM4aSYqqdkQfTgbKhHf6Uq5Hid8lQD/O85/Js5Qx
/hjMlHWEz29dTdCGVMGIX4smKuCFxrc9NYAefl+2JYuDX9cBW2ruCrwI33qpbAFe
Awx3MAD+0x5GvTXcUbmLjIYc3THiWsj239GB0KAZaaC5Yw/qdvt0cv17O4DGpZky
872oV5BwDDZCamhC5fKgkPbu6EPlCcH9ry8uGoY/UlXsuVMEKkCscmCVbL3cLtz0
9rXBkTs4E59dnUXu8wsHpWPGVWl6jOlV9jeeEZCjoTPyZKmjrHTNGnae5Ae3jYSg
el4TF5QnX/WsiBU/O/o8QNEyn7KA50oHdOeqTpPxzGP2Lr0QCRW9vrvZAKMFmnJu
gUUzK5XGWx/syhoIuvUfz7JPrCHEdcd4VDl6wzAs7YGhO5PMZjZD3KKDD89+Oath
Z4QKOwkTpntZ1SfFtb7j2BwRslytUjvQvxM/8T5WVVf95EMMVI3Pocm/R4WBiOLq
M+yl+oQKrnfl66E8zaToVusUFi8S+9lgCQmcSkGJ13n/YrN/wpNqLCJNPkemGy8C
qKwEH+3WrosQRcn4j6i/IqjTG5zyQCkK2d68cp++UpRykInalpOQ+PK2Kro4FGAu
WKSARRdoRb4EG/WejHkJsNbPQbKzvjDjQsvtEzGe36uKUOtuLA0ikxk7fD3nRTc4
JMQdMtg+z74TvS9qRzUmHGdjY/BV4Ttk9XX2WprwLVgawUeULQKzVUZiyei9XMO+
9l5XA1ynegSusD3POZEg4A1YrvgBEc9WpJAJd6gpTonAeKDhlAxG+bVBfLXDaPKO
pZGq0+6yu4rf4MfIj8y245aMiM8kbIvhUF8lmr25vcCygwtZP9IHIh4PwJ0Szn8C
Ii17TWiwnPTsa6ytP6N9xurVoRozag+yzmrmf5Y/guWOyWpSY7FElu34dSeHmu6K
4eDIkbDErnQwYs3UtbkheJVKS42yu8Xhbz1x9cIz7Eo6F4pzmiv26+LiTBN36OMs
py0FThjN3aSgkeMHY8ViKQhNxeMRUCyEf8UAj4IckX8NonSuxyHZI/KvVWXCA8LW
+0gb4D6KQv84xQtv10krDesq8ZIey228d2MQv7yAZ7G4J9don6KiCQEV+qW9E5Ya
RTVnBgyZ/A0QlbFVllKikDSZ+flT83K7zgzFf3LFPO+JJ4extF4Qj3ZAsB+bdpwa
49jMEKWR3EWmP4p7eyFeQIOj0WFRfriRxszfKZ0+n+0izFQkGB4PEvpDazzjDcBg
N985vWvgPAoVeBfMwV4y5rrsI2o86eOPti+bl+HH6s9rHBNlMhJHwoXG8dT3FP5e
N1fTncOwU6Q00yW7Ls9HZA9Rtzul9GIyLKZYmD4loBKNM13dcE51YHBcfDIie/R5
lKKgy0FeGlWqyWQiB+L37aq3qxWjzq2hXDWja7PvhgwGWjih//5ykYCqq4DEyWpo
V5WHpDxsS1RceurhIR2igRuNJTFzcz/yUpNvVtxid6mvMUu+JSy9fpghnbOyOM/f
vt9/uuAYw6q/DbfGCttrQlN6Swar4a99K3eZ+f+os/3kPQWg3Q/tjx3Q/SfddTgS
R6a8rOJ3r4cZxvMwo43XRemeZozEzkho8kfivfmgJVL8h26FMEnG1UPhtWj7fQvD
mSz5o/O46n8mw/Y5pwIprBbH9ib7RwkbB3eaViSDkn62uNYKayMMDCKqDR9qONkw
V9NHESsFjG+FiIV8VY2YKdJJycjdyu3kS6k01PiW/tO6zmQfwLtGvgOgeV+mkW+w
dAWPWpf6GD/m1juFXJfGORFzv2DIReFDx9fYEIq6e8m6qj/kq+xWwxAIuQp7wOxx
z+WUByVKMCWSvFJIVPSO0VXz2jncPqF0cEnVybQdPeRhOK6H1rG5iAEwBE/COh+w
8Hp1GkRw9V0kfq9J9TvNr09DSgrqX5DFcHy7njfMaaAgxdU8Z0hJGl4WN/wE8wA+
mvMlNIkBLMW6pn56V9PDqAKCL3vIqKhzkih+E9aOML8/e+QmBW54LD2UOANpsYAr
HTiApkEgCJqdv8UesvATNKOcsjd4GY2lYdvOWP3IzzkbL5Hvr8XbihtsFqpy4J5b
r1a2l60rLjTJh3omO38iek4rsh3eXcAuVlRuWYBH0cARwOwVngU+96ba5GUAJ9h8
5IJZxEswfY7d1RX5DXUzY1Dyxfm+ky9cWOe87/+DvtRROKbAHymaAjIuCXdmpdoq
54Uvyvqw5AQ5df3lJPhjrBN47ayv/kWC0PGFCby87h5OADVfv9/jYHAw91DZrOy4
WPDOalstLMfFrIZ++ch1VwTlpSHOKvxzY1SiuBWKDMEAEtqdkBEji2s4apDsTGJ5
xMGLPw8G2vt85iDmazcgAY5FozjS55K8ohVPt2azEpy+hWNKMtLC8ry31oTECRDm
oWExjjTEIoMt2ctjfyusUa6cTGjwb5tmCkfpZq3lJ0f/npbIguKlse38DS+3SbG3
GLzSCUWexafBPie7fP00ZMM4J6BNq2t+Ay9QNF1EGFexX8Sr9L6TBWxJcqHllQCu
FWaaTA9LJgN63kr0ETuTD67oNP0u1+7WBawPXvY+McY4NejyoztpFIIOzv0FCRLT
wc8hl7/mG/655Zi6BV7STDLOek1F24y6HEAKaucoD1SBuFDf5IIZWxydE0SdUtZX
0QKjI9Mrn/OfmA5WeEjQaL8bDxXGeqm+VIGDEOqM6yF5ENn0whQHOrMdlXg9gLvW
/+m7WLS/jCydBWDz6LBsNn5h4mZmFRhhLQQLK7V06WsfXVnssOEn+J4x+10ltlhR
MyC4JpwJuQs8qkKslsFizGnaAEFtritTVdRU4ohSnAgKdll+ItL4ZiNhvzaJBzWE
ODZoyMJKiI8OF2lzad55nr5LpQ3wgnIsawkIe8CKwqMyo9UDR9at3Ic7rqbjK8Uh
bA5T/uSCJdB068MJ4gVzF5uJreIEo3i6nhVvJ3LNOM/gSgdJbztFWQUdvcDZWuES
P1aI7DKK96mhoy1q9KnBcIg2Rgu2gxM6ZLxPJOS6qogKvFoNvHr4iXs1edhDLhIi
4TDSDdC4f7tZ2Cbep2fxNoPFffp1BA2IHDj9t8at5e7cyG7t49xU7U3/EzoYU/Hf
nNbp92Tj8qKOWHlhqge7lzSKC/GdoBcWHTuMuy39ERps+J5KDEKx7vhj3m02gpKj
gfZ5NJMWwQ3B5nn//P2WXKmHPdkYJkXgC40zMG4UMqXESjLncqh1T4jGx0DzakIq
k9Aiox4albH7WfJvwQKkCodZRn4D7ENJy4R/YkPpMKCxO2cYFjttITS6xQJpDy5K
kRKQsOt4Yli9TldZJ+sLy9aKSmBv8wky9v4lSVMWFQaerw0jjRU+yTFBCqvUqxm8
gJlEbHS3zne3wbA3E6ZqTjcksTM0Nv7/2LSxnWWZEt0ND1TAYiLol8d3bq4BvlBC
78G+1HS2J+QmE49FIF0ok2/+7lYy9Tqsk7RovW+Xcf3aoTJ1ufFV1GoVdYN7D5aw
1v8whhWVnT0rNq6ios+VLMy6x7PvqD+bR1nWDsli3TgL0GTm5HVxg2r0qmfNueKL
Trx8F8zjFV0DJ3OsSRz5xVD1eTGTyYSELs1SmVXTepWszKlzE3kZUnkVc3k1jKGR
AyHGwhOxZj4VxJUExAN8kh2PKg7FceGcKyns3POKlaN/w+TtATKFE5dcBMFqtCzc
qQIBl5VZwZYrwpiqkmcnfPaJi+Ooir4LHZxehy+CRYF/6OvFKoba4lOptqG02nGn
ye6CD3d0GwkOzWMy4BeXhs23TEiSzzB0Sj8hdqdU4gYOUBbiup8FrKj1SE5XzRUT
e6lCc4Y+0Z7tutIGxAtGeCw59tHNrgGHIwL5YQXeQEuQHQquc2Jg/rgooiK4wqWf
M4Jcy0opwV6niOO2SxGUq82aB8mWbtj7TRK9yvUj//4FOiwZiSG90B5QkxNtFl2u
uXAnIHZH/IpSlTWeFsd2AHBOzQyhQv5RdUWXWsRG7Q6Crh0vuvoAqk3fjyOxw8Qg
ljqXMIWWo2KVKAfkZhqdCo/rRZ/cjkzXgZlH+qA81Ox+JReICuz0cyQFmmdduut4
ynyjjyTqU+9J5BgIgNew8zT5O+6/adKVNYQQrDI2ocbsqVLNVe7PuTZU3zx38lMr
RylTDkl/SNLsq5fIhBMmeI3sfqaPXNtL0BdLC3Xs0bt5C/9QcOpgygTDY2Yd9yOb
9Op9nKMSbF6wtNAX/P6B1Z5FmAF/MG+Sew834nKvaFQHUlIt4PVvNTA6+8hq4shz
y15FGGbixgVtianukipg9eAIswRPUYnKUMiQIjYeVl4cgvJplxLH5Xuf5gZDTeTM
I2vUdUwoVOKSYPrWPPIuYBCadR80LY7tNjdB1a4sTthhyD7iRgNE7YL0xMYTTuNk
PvcGM9T3m4G4KUjpdhAH5gBJC6hodyLHiG9Y5qsXCC8STwFqWvyknWHXOyyN1Bsj
+no7djVDIInqn/GvyeZr3UVym7o/BceY0SPh5sPBsFEXrrqyOhoyZPlhOxMb6RTn
oaYJXYE1Cu2eDqQmrPIaTyhnSRWS+KqJdILBabfGN+cPSY+aJy6lPVEe9ysYNJJJ
N9uojgoJufnar8wrTl+nkkGMKiYxHAhg7sNx6rKWqXN+/KQ0/Dedf5N0vR2BXKB2
3HKtoONywTNxNmhIB0cwmUtGtvpW1lQXLiKJPp1Zz/GcWKo5U3zH2L8cuv9u3A4a
UhsxrbXkqBzybF6ZsyIeyPLAdyPtIgWs+njMSwtnJSv1rXTBtWcwjRegomLCuIyf
7yiZjao2UXMTYI8iMv/YC6mfrwmOwLuLDXoF3DOyPiwmiNga9Uhj6KwCRwPfkQGL
w+8dBxCTRKqFjtfNLrO+5oxESI3ZZGHnh5cjO93/CdBPZiqCHgXW2tn80D6cPDpH
DNwY1CaDhwRwO9CHrtI4QIXA8wCFSsBx910wMsfedxzOPxEwyGIbhPDtPI6cfYHE
Y5uZz1wjojsD78YUYSU74niu5MQPL8xU3qwz8yQkhFMcN8rCh387TXSTaZC9gDKH
XpKHLnHW2cNbplAzRmnkjeqXxcRYG9sNnkIVGH7M4OAEg9OLZ1/HZGc6lNFM5S72
MKxi5a4hEcq3yqG7MH6Oh9AIwZpENuhQXddcKMpm6Unt/MwsgLuYV58LIc59G4hV
feiVpuvxYg4TJUpLfP4V18m5SswHk4Y3+HiHgFgW99Q2Z8c/BlHb3G1g2szxAWuh
WfgXcqKKL8rPhDRE4oxbls+XqdZ9XVSqAVNOR9lt2bRo9wL2MfQGtsATpOtXOFU2
xABjmarXNDoE4kLRKim7XngUjQnIDeURvLzJxpsN+nLR888zZeKp5jc77RmWti3k
ZPM1aesYmxQ8aWFgjtWhiOc0ifwEdnr8Q/AfT+FS+DfccSi3OM5OUHa4as8lDXlK
Fzye4a0vwTCiERk3wH68f36sNDeNeOVKc2eCe75KidiFyASQnq6U060XFwHb1r9z
nWsJ06ma5qiY7LwoKgz05kV90Qis4ObTMkcKodrxSr8sZ/XjdD01o/YbLCHZQZEx
DTJc/n/srcXrOVoTJzcdUJ3mhkttcSATjKYGZzDMEI/G/OcHv3LKcDAAELfaSA9Y
tGORc0LCHU9LaihAnhLhyraV5kNE1OivrCcrJae9Ny4Yi2X5tZKQkseSl6M9ETI/
PWlLE5QUeWdHcfYoQosb73YRqQRabuIXzcpnlmLGOubD2D7HtyBSA+n1IJrCZeme
XefoiJeA/taTQWNlP+/SNEpI1uJq0aUIYhqdkiRCRgHH+yfQRu/CUFIBHji73GSw
GqM9JcQ2dj2ocMO1d7GzhXq0UrrKLkEO8uRxuhfd+wICyqnyPrweZwW3H8ccAugy
wuCekpNmoeLVHhxPXOngmMFdIMTRhxP4Tl3HjaGkvNpAG3oG/TuxpiaZ5HMMUu8N
bqUkW1B5Wy+i2ffv7Z/Op1aKnmO7wWHNh4tleUHuCZ17YT0PX/7aEsPxYq069Wim
C/IhjPaAxxMgKKlXV5IVtU4oT7lZH41JTHlFCHwojVwOGDwh/7VG0jNxpkHmg2SE
Aswp8hODtHN5gtIxb7PV6i/aCznA+tYbZbEfN4dhA9cjeDfTTAjMyYoePKoOBVhl
jjRje+ishGNNpdTSIqxVtvSZUdu/9ec4Xi6qQS8+OORK63k63q4pcVjdPJ2dZDVX
Q7d7IEQs/MIttQiGaUfZymuEpmR6GcQCHg7iHKx7HVWrC0cG1XJZ62Rsg+qaNjru
FVMaNI26hTwEV3q4vybr5Rrnb/plK1/uHlrjPXVxxQC3WxigamrWhUgal7V+bz9S
gWXRis9GT2hWjUDXx0u7O3xY/C5AIAoM5SzmElUj/b0+PnP7A812DaZ9MJfrfkMt
6+NdRDdiPjJ+LcM4Tjcnn4qGJFaNIZ1jtu7gDddYVWLeeF9REUWz6/Fi8iXYgu0r
+ICdNKzb70WwKC9HOrx7jgO/hbnxB6idSHCdibIdgBBXB1h077Z/0ki9OzFAdiPQ
REd++crdGW5fcbl5zR8DP07HBFULKTeKKDsoQ/Z1yCkEksKISPDVO0H4tZb4NK7z
ASRlbphqPvn09WwZKlNiMEwAYJQ261TUsvOlV3MXBYDmYmuiJ2pRMNY1K+H/9QgC
XzxKdNJHooWdoYvdhl/ci0XKpjP+xnzoyRkfM1N5NbG+g8s5dCotoyGfsTUe4PyA
46/CwUKw3IMyE9Wb5ZEB3HBXDs4A7eKKEjsgDhXliLzamlhgp5FJi7YK6fkfIAFj
ORMbe0MG3QoPPE8SGWCbkq1KucHu5Ioh4CZVYtY3rzauAxdIDC8lGMRTeI8mFpAh
RGauuedLbgYZmtzCpLN/GQHcpnHdRCMH9mon/CyVAT+xr+vUoezTe0piMSrHq3KM
NxWbXEQHig35oUgXzibBR9QiGYLFpPlb5LyA+otIwT5MSzCnn2TYgMEZAnvngJG3
lhhsxhSmuzIv6phYkDV6HiwmoYf4kcEcl6RPNtMgim2EYdDFtunaQR5A0d8P/v66
RZFMYp4qlHfJuUunU8MB0y1kxF8wF5Iza4Iv7Lxk+1QRpZg4sAg9gWHzOSCYkJtj
BSJKtgA7QEdyRBR58hgVDeoKvplwy00qPqpzuat46bqYxFl6Fks0RvLBDbCHNgo7
cechQ0tn37xGuLRlpmBq47ep97x1brFd2JlmOXj0NM42gNoZ1b3ykHoF90UFkoVl
ZfRl9qtclgHpD1XQthZGbBeO82z4YVITGiatC2uZ37WjufmGqLDUPdgt5re3nln9
ZNsdwjpLhMYbqYPjWcToHcWZRpACbm5P6pEbFDCexLGHMDdkrJqNcH/kFYnXW6dD
b2WMoGZeqQv2UeSKi7WYnL+wjLnBgAz/qZI46IYI7njwqndPtKyPIvgjYaZnjKA8
QsG3XxzvguxolTdQKqReQflMUWaGAVDWv+qz0o2Ugi7l1dTslTQ2EtLItdR0N45/
E6th8mNfhFWY8e/kFpJtwPL62C4ON1gjahtMlnl1Z50XG2fVmvWvI3PyvPmDkV2f
vzMpWGBq1DbmKj1WBb0KJSXBDFthrpd1divtyAwiNaCn69LIiOPmCimc9jHdAE8P
hSyKAHikCMN5R+0BM32lqR9O1ADfKts2B6NhJQDqvhs4YIoLB59vlQv4l/RZlywQ
C9p8O+uJuN19KgiaM/oSZ9ojIQ5YX+imqL8Odlgk2wmfFDsH7TzeLCF2bfvaK8a2
+ycFBnSyIa5mxiGMr2/ADBRBM3nGT9XUfCAdVDdQYB/mLnKh+SJaCzHDhNOhHOuE
ECFiAU98nimafTu5Ie3KKfO6K4JpTowoPh3waqqcIVS/LlKX24fbiAM02HDdd+Ha
hiFQ9mN/8fQk6AT+4EaiOB93lyFlXK48wrFjC0Ejnm+VLOLOdE0odHmi51e8B/Cr
Yss5Ri/s0Z8PsMK4W5ceYQcJAHmspAZtaXKIQ+3iq3al2LapPWjs9DwkV3E3waoi
3wy9/Koyg1uM2YlkUl5HjzwKIfJbXuE/F8A9pQtk5/908Ztk0g51VobIy/9Q9d7v
pgyoTT7rKY7alGnsAwh+1rqI+b4cj2xyZFX8XS3phMlLuxf5wR+b9aZ3A7sINqeL
4a3D2oBOxwsbmk2bQ511RBAR0ilaUHAgOyuLn8kY2/rFBMesV7eHKwSWp0QQoDMI
xbVOcdqmGckrMuXjCwxuFUXpxufm/fk53ggCrJhW0dGWTD1TWiEyINTPoIVCZnsY
W+2LOf11jFSq3zJZY9Fg9iOzUHIeGTMApOh8B3VczYMPwOKHRTnrYd77GW9M+jNu
IntupLZcqjv3epp/ESMWkiSPCm5pG5ceHlR/UEy1aA9VHApYXwejrP4mvnauKbQy
9t64LrfHQvrtZAT8jLbKdihyEEoEhHKPLSquT1le9uiPd2bZHmClftdjEVILnJke
MlnHuyG1N7KNxaQ/GioBQH90AskhWWrBWlgINE0J89zNeOelw4ZetPugSSsJDvLL
K6iIDY1Al7JTXKR/fSWCIx1DsnDkjPi3zwS1nNuxJJHokltGxyw8TdYmA6XJUmsO
DoEhe7VVnUejKlSfxJSiXer2+lVo+aV4myPtyJm9r/N6qvERULZGAjPbJVyadwWZ
TBv42CvJZ+mPb+MVzye+I110cs4zz5yTQdyISj5ToVN/djDSQmn68SgQFDzd+7Wf
Q+hdU9vxhZOjo+TEgeol0PGpW88KNL4fRJNrEFutyqg/44rn2yvJBLfWhJaMXP1A
1dAZenhq/w+QL0LL7lRLg/ZwdQWCcezQVy1Y1pj3Dg2ap7Y1W+h8V5Uxz5HuMyi1
+I9yhyo5XybBkojAdzMCRnjbmhYdGXTk4YQxAcc0V8Nr69gs+z9hL4itx+52IOxA
OAJh3TjU4u7V7SWL5niiSEKdMub33zOB+pSQZUWy+ZlFGhaycjm7MnEiKGbT2ESI
0eZMfXTwf25d0N0mRhoF+vVnF2sRj2b+KDepV17q1TTkLdHmDUapV1P6NywLUywK
e6/yFxBk/xnaUOqDUgzkS1NkEDRYAEgNBJay6LYQZKplm2P5WM5BlUMyJK6CdFnv
UxPRbWIUGBqGWWO+vhIaXZqNEB+1a5LnRlOg34dxW2rndO4n/yU73X8/2atFpmfZ
gvvwUH0XOYS+SxHIeUaVy+K6+fABcb+dcjDcXOMN3CYsNT4z/dCSta+XVagFrPqm
EscbZ/RfoZ1y80UsOFfjV9VUe1tnYTfAA2ybQqi8vxjhSfBvoo97sSyBsvJzgtpH
yiUBoN+u1PzkqJIN0NJysb/h699vx1sSIPMEHNKWyIS7zdeBYur8Iq4GUCXenmp7
4DN3LD9uaGl19d00gx8AbkAsJuQds3oxdyCxmjFWj02dv3bS2h+LRlc8i0L5avie
zcMtQqs2GzjJkwiF6XsHB7y42yIK++6MM+WZoRbxYFv8s2Z8i4f8mv7YgImtS605
AUPnYUfoW1L5YgFumAqrZYEbBUTfjA1RT1bUT/j0RyHRqfk1/oUrRsnIfnWUPKXD
LSGZ74zsHxOwLC3VwnsZhj19PwZX+XYvPMQovt7nUeBJydA/1ys1PSAmqrelupV8
XqyTqEgRsPVWhYBRW1h+t/Qqey+kkIs5ni4G0fs9bJOB++35iH4omhBUK5V0D2ML
Z4b7NsdGpzDvaqmOZZjYW1VVTNs/RPNkkNIBhJClMzedVzY2rrl72UWFXL1KmawZ
+uHx41XrbzH2odJFO45YxE3S+PJQkeh1DaIQcHBd9aHMTiyICaB7HKnfhbVHBD13
Lp6ZTqBpk69OIDQRquKvA51PmAUuq3vZ7TxYgdwMwtJ44GWFR75gTNFeY/Kezlp7
Gtf1X78e/7ONRU/oUGaf1hhKyDMo4TYmL+Kwzzut0YXwSz0uSE7C46YnF/z5RDK/
hnUaa4Duc0raHulpjEVjWV037a0yA9DFH68Q+a/ENLXu36nO9ItGdhMOVDIpBSy9
OJe76WCGLerdxHVZba45ZcdlB/NeD/AVcti2bj5RRcf5fKvNzTDj5E25RqFrELHn
hENqNspSgGlAdrZ8AxhwA4WhkxGoYaIe7nwS4j925JvGoU48HhKtCRGDJQ1bVCIl
EgZzIorbhKjv8v9Q1ixVw9Vsg2Wry88a09lC5RiLBVESYHBejKE80rkXdX4ROOQC
GnWOb52B6RGK4dux13mUPQztjLShmfYiYQoBZrwOuKNb34V1HcJ6h309ZbRIUfuF
vW/Mesp0OsUUjzeeGZOeHDXLd9Lw9YzxMbOZIbhpDbiXqzNbuvqy+vl9VlAetEbG
vYroEsi7tmJWfYOzm99y3X1wQuZN+mz1BxdGay9rnrnOKIL8WHfOaozc84bKhC3B
RscqFqzJ7BK1UnFucg0IxVjCRNiBPcrS4500aLz3dd4Djl7lkfBnPnw1m+WWorBT
mS2N+iAm8o+O3snHZqQHeXvPb3GVF82OrYATn542FfeOuH8K4dts5Hpf9fJeI/am
HQYbDfVr2/Zv1Oj//ocPcy73q4cHPrw7GSnwLokpMkKP2EyiUh4Y1O8TaAmKTb/c
O5g4eJu//e9PdS5DxSQwRou68ejOjJ32NB67yxPxrWAkFErqOTvQb2gtKFiHrW6Q
BHsiFML31Wn89mSHcICyFJzNBGS267aP3i2QqfkS2/IJAYMNpntD8vLOp4dYEBWr
0SX2+7f3s8orn1Te8fTJh1MNATDULGq2R18aH6kPrzfbXr81/VvCwVLVhthfngKK
pMEccrORMLXVB6n4gsZg8R/0HrjMdk8LzL79+XiWP4/M7Kpln4zwk0qIsS9nnj6m
ixg4GAtuzW/m9pvZkiC5t+EXEYPHUVDzfBoYH+hktV8ypvlTiXIF5LSrwZ/FC0Kw
ktrZZ9DPsLnGhzXg/UheTzxl74+puXUdvxubsIbnBqek50/VF4kPJjZd4IS9kVlq
AgX6/2qusjXClt7psqviGf3IlUn848IBmL/R00Hw5GxOqvmnod/eoqJ9w4IwNZgj
tGwupcoxiDL7aWGFqzKhPh7K+SWQIPxM/RdgXsUKZDALoOMDJaD4LAtGObzWH2zG
+arhz41Xifniezi/2sxYgUqDugSYBqrRUd7UoxCtCh1kzVxQiBXUbAgMxjVtdL3r
FWuHa3/JHgO9r9utN8kr5//oxBEYUz2xG6MzKdP+xkUVYud7QquC4RqE5aTrNU+h
mvIgkUxUftS0Oovloe9n5jzuAql8RQg5pA72t2KqXdhjwIMH+4A1rL+pCXdgZOsb
hcSB3dE2dXcyoqGh/Vl/s7TOxaf2H3kkrLAqzxUjSetd6+J+wY0pOYPycMazYTmz
NYnRWGtserBovUO2mOzvEu4DAEmRQhzDWxWHkQ4/u8WN/dhCldzOW09QUwr4UXJq
vqRNlMiEgcva1ceiZQz1NU67TmwCFvuXaysSkn0UD3HpVE8uyXpI4t4Zj5K5Ohp2
+00P4eZwSuwy4Z5swHlYHUqm0hFfENGdA1XrGZAg31q/0AySiPsMnOTVIJgtphEf
SvdTzFdEg8R1L2qh1mcsDTrNxbADcE7cFjfAeB/0FSp1B1Y24ZmGgYmTUq66wZ3B
fpHMdfv/wcfPYFS68xc3+zshxRw8afuD0tV7/XOl6Y5R+YpmNSEAbUw2GsqSqMXq
HuAsqkH40iTWRlwFTdcrwA9rJFzCfOzq6pRjO5CSC+gfvBLNa6QBas9AZI4msixA
kkQWVv9o22T9a9pINU20HIWGE7QyMFtRtAcLmMIJ2z2NGsD4o1xnBO28dxHRGJfn
4bkwTLJID+LBJUiW10jg6mwJiwsCXyua8VwsJAA1BYNaTYGpJW0yPXXVRp64TFlG
Ypb9eilyu30NcMjoNWDrTSoUOg4Wp8I9S8akVtaLaNklQpjtbUoPMRhq0RUQi6eL
7gZy6pBMtWxxGIcJjAbPqIm3RhrU52HOXFrkLu/mqct3jWh5tp8Y3VVT1YrbamMW
j95Dfa025d/TCUHkMR7Xs1UNlRenkBUH2pOvHcKYO2KPhovHNPfByxx3gJ0eb2QF
i/+EWW6Vrq8tVASb75n63f5snq4moNF2MVngDGoFLq4iCp+msGRgtWN9iiQsXoct
Bez10JWBj3JwmZTzgAPNSD1Q1l3u2lRbss1a1crwWullN33u541qXfthfuNn+ExU
PEv2ya26GcJHDbY3xIcAo4+Mj5Ue0WWeCZ3W3MgbkoiAyZyCgZKmkP5nLu6ZbHFK
swFmntE9SUHNY1IkWoZUku9T9p9iJPecM1PoPb7kT9L0RWl184G0kCOTOQk/P5G0
WTFZ1U5/6cE+j4+mwC1h66phNm3EP/ePG4K9RRp37t9Nq+CoF7nejOABRXngtqdt
OnNRHSkgM9X+asNy4Yv7Cc3LRB7wXcftdNjJEnkWP4ri3dsgaJyFUEzaN1vFBuhF
tG62rHuxqnXdbn+x40NihSHMMt46SjPE9vBJEVKX+heoDtPRS7gxvXYUygXWMFxY
bxvyMvYD2b1scVwBHoBbBcWqGlCbCn65+54ZG1I0ck2A04d6wKFSIAjSXmL4ma8o
NvqwIeQQ4CDrfMZgKO7tA7JIo1C5OH9Pfh4N7sMUsNHEDB/GU35HSK4dq3fRGJlA
n1519iJBrcyeFefh11uCDmbwq96QUGMTKJfdQ+zCG+TWAOmQzaEtoTKh09x5+HnE
By5p7j8in+WbBnK76KEmvSPdG1U4PHQ97y1F+Lk7ZBzrZshVWToNvdz36GybOAl0
ZGxvAyXt2ZL5K5RwVRcHgl3JZCVAE227VQsDo6IVlfyaBF+kmY9se7w+tevV/j/W
OTgXlabUL0mk6K5lYW0VoAGLeqY1Q/OwdD9gd+ThOiOdIdMbGMnE0yy24hmpLFCr
fZlSfgRKf4bRNWkiBD597dAsG+43XVru0Wkm4qD0I8VBkXeHPXCr1F1DgkHGvcOo
5ngRNn6cO+L7uuNIrUmGw/J6oHzy3j+XAk8VauMluoPNHPBhg58o+CuSpgaTIjnc
NLqOwj1ym8M5mo0AcYcXhZUPrz1mQAAfo2rby3C5wRuv6RFeYDfO5bK0g8z8ehcF
G7h2uiZymUl96MYTmxLx1AGJA7U0LS+AHrmOfPJ37TisSsHmrPEesQ42h4HcTiAd
PA7oqw9meRXJXQRiiSa6Ee3wcoq0jSlPDlq5s8gWpkdJY6bILR1U1FCCgHB26MUW
tEwMcusZIUjEaTLb63okZjeVhnQDI5lH7Gx5DLKLUN5oZIHh/w13MHNC/8MybosH
FsipWWyCZH4HHbWG5sOS8CCv6NPB1S40uzkPI4IK/d8bS6nPyJOS9oE/uNmVnRdH
jt9QZDUIeAEcD9Qeq/ft3KnsBDWT+1W4oFhvb6nRV1KMIJhEGSTvLNeyxgn7h4ce
BtYLZ9FHBEKyojAFP/9QTKrf3gH+D6o4JEy/g5BK1YJ9LZLSzGnk8ZKKd3p3fS9d
yK0N2ymAD25l7AiX04xK0T4+Ut1+578SDp05akYsim2LCMJX7ScUXSVBsdw3B/iW
sT860FuzIxJtsM7k0us9cvrf4rjqIXvtObaIRESfgq0+WoGAX1DOeKJZ1Mvae7Ul
o1QIYr/mdPNOZWbMOllLOBsgjMD+3YPJhGcUkeQ2MjBON26vuRxB0OWIOmYN5PXD
TIcyuOC1deUH5uIvoYcKw6FgRGNkhqiMeQ9EqyvQyikL+aTMjbj2PUNFwhZZEmdO
j7XZm87jWmviCEGx0CgASQXHdEMfXVgWiLMLYEr2RS6TRliFUKY5sMdVdbqxIf94
Kc4bX7MVWdkfhzbvMl7bGEAiordZRDfUzpH4tYALv4yX8hlZ0fBdqtibbuIqKUvK
jI9nvJB5w8ISeyE2cfvbVCetguWKc7217PsltgViyw+R/MdZ3QJ5sYQ1yq868UWr
4HeBrF9ssl4EsTQ4VvPqj+1ZjRo4zweAmYIso7YKc/uE6K21/hc0s1ZZCnr9e0Xh
HqAEO34dExLpW4MHV9Oqe+K48Wo4rDVf7BlRPaudbJ18t6sLyuacjZsqTeo5LjeV
6Kj7//zjMx67hEnpOz4bV0p0xMFkunWhdsD2V1NZec1iPSg6JPTeWtCqmCt3optd
X7qY1t+o3uwGj0X1bmlh/p5UqtteoRvokVrc99aQvoWaqYQ/voydWZF64gctq0M/
hTotHd0ZU8dcQwrbZK/mIBMcHFX8EWoGCHaNtLQKkRyR5/surSLlbzzf2HPRiLm/
mgW/o/RIsbYUDEXwLscZG2isITjoS+uBr5innsYVcK+eyAonJ2PPqOiA7FP3A6PV
HCLxhLes0/Ryn+9CgnZr4YIQfK0Pdc57ZNvUlQ8F7E7o1+ljIu/8joi8dYrQRIJv
uOvyLpwh+IzoAcJu4cxxHD46jVVAqi6jFxqtjPdM5iSujxuO4ILB3I/FYz8BHa56
unnOBJnGi9axVbx2/PkNF7JySC9mBYwyxsuKjDpkEVxzOrAr6/21sOSeoT4xC+qo
CVIx4YLtxD4hdiCoEY5+zdjEmp863qZe9X2kaltaM7cfOFvwyRtue+4fSx8Il/Dc
ZO2bCsrJ7LPQs7ljspYUe1MN0vxf718Vmakl1D0C9jc0kEytpl9gT2HlcbIXa98r
STrXEBHilNv1/MbnWcIhEPF1lwg29pF5+vye3qdrZsPIxWwTWAPwWHn4uWzePkUe
rMIvWWvDDUq+9Pz16LyJY77x7jgwlRKWckxqsUnCVn/3KMVps3WVZz5Rhde04m3S
cG9XqhA7SWTs6dnhLOeswiOEUiYoLqMONxp2c6Nu0FkOrYjPTQrBzVz1f/KUdyRF
hBmpXqRPYM9aBb5OPRO0M3olvJbmQAlg/mWHcdaet2Eo8dPODLkmx2D0squ7Z1NB
7gQzyqm4vJg3YEOsfTw/KbkwHhRKeNvEeYLJsYMMbJ0rit2ZdpwffVo8aswpfNBk
vwSMWFgq8LoVEdBIv8uuOeYQWhFupT+OZjtlKi8coArvkJDSB1ajQYIJ5KnGdqHI
pW8c3o2nlvwETDS/VtBDvsYuI6cm/28EKcpz50nSUZhaN/ObJUWlHb//yZENW3LJ
4XjOEuy9jN8c00CXcBXiXd8NioZfiLaQ3eDMsfSP1NYYtNuNetOGzl3EjLKEZSKs
QJhL0yU60DwW1n0coIcV9Sge+sJqhTACWmVhPU1Ix1bTkIPqiLvm0DMd8FpnnTuI
LfxY39dObUu9lW0ogkl3iqZKZ/L+s+08fdGDyPh0P+OV5kL3UFGiz+BdiOfFNqA/
hVl++xTQOL303VYC3xqVSIL9W2znlBAUK/cMcl731BaBfocJAcq/wcXC+1uAdykb
r70GXkL+RmKe789XRBSRDiKhbFUrQ+552hRLto/hfI3KyopZFl1zM2WZnVDB1oGI
09fZb2vT6YDlK+LVraAiuycquhgEQUPY7YGC76Cq0XcPZXLHI9+dcRo4a1V/tUAW
FJurOf+hZ42pvWOyLE4vAEPeUsGVj0gxh3qdbntRKEz17PME/AaKACMGDXBV8GFz
cUhAbv08VgvdECnEv5hXKJtnr471lB+sYMjl95KtyDSFFYeUUP/gcrngxUB6619e
pqTiKDLN40G6Rb6lh7Ev9EjodC+LDOFdpMFGR8sXeDpN/PVozwhj/HUDkIIlLK4O
/Gdu2GnU0XajqP8ooyccLhRS4v9zI73X/17u2j0zokPf8KG7uqWaqp5oJJ8LMsh1
VlfuqtjTUhMZyJocMghI1cAFz5nSy0SGUXdfBhSssCrcO8nTQ0VfdYlegO2sZ5y7
XeA/bJTm75RJhtMdiwrfihFF23hKmV/39DNIMj+jetnCZ4r6JSIxSazidon34l9J
TlY5geOqoS5xWnNlw4Cq+DUluXej94EI2Xs0mxzJVR4/1QSHzWyIuJbHm4J5mS6S
78apxUHfzGGfXjXKFAAom5Ff0NaU7Ie/iqNBslg2XgaXwAxAOYValieasKQmJtq7
yCudzc8lBYG1weUddV0vMivXzA4V4MFEkweZs3jP38bMd+lvVTrq0N9H3OiZM9RC
VdLp0YsZJK/ScmDZdyQ36QX9T5pUae+n/rl6Y3CdsEdOZCEDhAqD+29y5STM8Fec
wcinw0kivMyrcml8ihBlxZzYMZWW1id2A6aLggScaYRL8YfNna5IXgwQ/lsAhu1N
KGBrnyz2r7JrekZuRl3z2Qgqktyo0xgZBc055CIZbTIXkogRQVhjdHPdj/Ua3Jo7
O4O79ZAE6WEgb+q6NLrGziUf8djFG/pjOXNA0VqxxtNDMAilmFlPq4Y0VZSaBKjQ
KgliGtehpCitUnBPeS6K5K/gz+h96BUb+e+OKZSgR4wweBY4J4yc5JUAIX/LO8pi
2nGnH6DibWWc1TgHJhXsOhqF9/BeTlBndLmKocbfMzjB4xsHPKsEmuB5lv0K8YSs
grPHI2rQwQmEwGJAyymuHwNoqxJaBaWHNycAD/ZSVK6LS7p08IfVL3OFzqfT3gWb
/doy/NWz4pvHVNzom/2HTQmQzyORdXIXZcWoOaogshhtlb6FLDlSarutpsLDvkcw
ZPtKEM48hOaIG1X6QDs8MvOhofcVosnOMM3lBKQTRFSOUC3UVUxxrVugbQMTJf5u
zultB+larcT3ZNoFP4Mwb/UWso87H3xnwE9fMiSgWgqh3dhjLVKW6AR4/QU4+6RQ
LPlltirz8ajLRKS3OWWcRGkGneINEGH0T4Z/Vhuqi/hZ1aFm7ZLKAlbq58XTteBl
jvArAp/QWzxwP6QaqNO0AEEc8v8SDaq3b7MUjSXeE7YXAuk+g8jGhnUvlxLqxyL5
PF/HF97BKNuvMOYJmM4ZTRRq9SmCzak3cY4ime8ZTZyoHP91Y9qjmxN+TlUqPqcD
qBqd6gSE1rFPGcBqQOPX39yOXJnPxipB4KQqdwA3TVDEoGdnFBb33GviNbmIMQ7p
9eLsRsvAEYv8BD3CUyu1wBcG9fy0IiDjCzBTOQzToh8TabkG8Vo94ujlPbMIKq1w
Oyobgb7CJg9hqDA1tZFpaDCFV8z02T4LpmVY0xZR/nZEVMzZM49zCMRLCepIuBtd
sEazQqSauJekWX6+HGsGCIQ+SW7NUahCxFu9nUZdvkQ3Aj18eQNVdwSG7YuCAzEQ
P8M+tNr29enGrA4Xw44RyQI1a6skXb8VkGbPHGUrOsXQc/oy/Tgt/tQ9jUP7AmrZ
S9VlnOVnlt4SECXwE1W0UlLn97xp26pgU8Toq9or0KDvWGozUABWfSqBpFtLeyo7
5GpVFWcPx8JyLx3KHmxhD8l+q91I/2yGjO/MqTNWlYlOyfMABAr8/QTTLW3eQN+D
8mKLIBLceyQMv1e86lR9tuGYiTGEF2kGnruo15fGLCDNXykuCWBBt/1P75VsOoxi
3dikDcebEfbt8N6X0UKoZ1kSJ1+U+uavhXWgU3W71VCBRCTmQvK1egv7hftme66H
FG0UrR3qCS3WuhVy/LYAMcfVNyFRjBRPTUbPwOgXlwpQzJ4YyQyIe83VwybPYbsx
uwARV7/NVpFRpP5ngh7xzDQloRj9E1pguwhyyW2To+CJcHOPOPCpkL62kBPrQXPJ
paYfso0DI5+8lTUTXWr1wdqli/RimQrF5G63qyIGpyLOphs2/oPVnw2ImJxv1H2w
B8+qqcoPxmkh/kAqqICTLM65KHcIbfmuEi7OXN6zVuaLZgqDvhw4NvwAMNTWZbFS
65QdXvOtDxCkpb/sYqlrxc+HYYWACuts4w7GiFSMhc6nJ3FvERPFD1QSmG4+JfPs
hwckc6IH1RGnq692iRGzjV3InFETxXk4DzDMoI4DBVckiIZ+iKhxSADtlMJ/hXYo
58eDM6YbtAOA+zusmexqxbTrQLmAyFMZPEFqOOi5RRnL4bf5bWdmN6c3sEX/D24z
8n14qfrb9L0o7nIQ5Mo3kFtP1SXvxnIKNHo70KGKDPKe0RHN03fwV1Eu6CU+sz24
t9jEL+liSbvFTqeF4w/WI0p53DpZJ0ANLeWROTD+qLQ3qv9/XXiP7x4cgliKlqIC
QCDZDNNkNJHEKCw44TRysMvsige85uGxJZB2WF7hOU9bTAZdr5DvAMBW42yHHF79
nopqvJ2wPTHG7++gmL90OItKWGz0iEPcM8dvWgZN12htX48TIYmQbDLdkSuQTxIG
oVHqDI2pp1/ehiI8nHutMrLlzBMoykFgNJSaIrO4lPG8N89p6jDxtoLXYun5+hGM
iwNnCQfF8d5kYdx/C1SbrMK3sttPwDEuqYo4Ja7ig1fnSZ/XdyFTht18+cgpF5qw
CD6uMZnMjguMDIwcoZls7uPArEScY9Vwg7gjq6N0ydTvrJ2cnHKPWxsuEpWRaoRz
R0u8y7C806BN//VWdUx2iMfxHyJENOrb5IjW45vX6w7x1mpucx6i5x/TIeG9Nqtd
N7Y+HB1Sn5BJG/7cpXgM2vjjSF74GroAa7RmJ3XgZU2tCyULhlmzY8SwWmleGerG
/fOpYAtNM9q4d+OWw2kZHkci8/45pWU46J6J9QgAYxiPSOZ06VfFnEZ76YI/skoB
tRssVpGPRWR69Jrv181/Np/ks6JQx+xTQy4M+dMLQDYFN+itdSJUQzNxyHXPshd8
ULa8idnOEgxK57qqZ3/nZVak8fYGVL6ajoAx4ZpJEh1vUzVUnUpXx6oYGsJLw1k/
klsXHw/fmNqBbH43DnKvlWdl2DeZowEqThLU3fXfIxmPhiHZsAWEOU4oqcg52gHR
ukmDOpuDIDnUe9z7Mwt/BP7UKTAvUsV504KayS4qXIiRH1uq9YGJN1C6y5EdILa8
XupAT9bTjXj4/5Y4KUKqLPOaRD8PNCZio1BjQ4NZz/r10IeT+4jbzjiSEn8K8ga+
quRbR10FAGQp6qBeKEvwnILsfTndjg7n4C6jqVN8WFFW6UzDy0iQICpyEEzDSHca
MBbEp/FIM6nYiWoqMM3Ex0KaK8LiCvLytBtT6kXyDWUcaBKhVkXIWJPRWEaT43nG
QcUD+ODvE5gAu9JOFPjICj/ayrtgYPaoZ4MROP80jserrjSo5tl/p2ie5SQqf0BX
O233HRQ/wugu3LkGt7CznjtCU1omySlqdGQrbIPuO6F/YUzY/ulYMO4bqnJbMgb2
yV7XgFawgUu+8KjzJDqfE2rSK51geGB99bhHjqPvEeViSAKE9Ftcj4ikye9S3HyH
QSO0nLJxS4F9i6SC0le8P5M1rFmEbqcxeX1y7Bm5JG/y1mcEVhd1DlhK9tuyKR6F
YEYjkVhchMpFNPvhLipRRzbZpJLlV43dN/x2yV8eO9UCMysr4Zvht5CyFITbn1lV
fJHzYOusi5JtfP0fKnjLtk7MbriflYJ0OzY9uef+pManlxvzzntyjrTUeiGJjtLK
FjEFy5rwXwnTHFrLKizhC7o6+KMAKrae5ExIvMUq2ZHaCZSBqIfdXyQiZ8euB32z
+PdVC3x4PvuE2P7ZvFdv5KvqldC+mRG0cG/Vl/OW2ibCPhlQp/eQu8sBC3je0ekM
/CQsHNrJIoIWj3W9YEMewK6TvDRe0i5pNh9rVeoG1+pUQG6Y86hho7Ev+dgDQH1q
Svg7EAgHCf14t9+J1LgZZNFRyKuY657Dn09FZzBZuCXKeF/Gynm6zSjxS4cKgKld
A5nEeWAJpSjYwmeigA4gJgwXXAq/nFjKz2meMyrs6fJuDe5anlsLt3fOf37ej3kC
Jfi11B8IdefXl41mzM6klxdBSgbHM0t0kw+xNGJyW/5zwcRePWHZ1cc/dV6Fus6v
uVfzzb6YSDasvT/JuIXQ2s/BpAKnonKuyTtRWZB0b6AtjK+flyc5OrgTFdWem2HB
4VVr+B4X4aLW0OFSYbMb0Bgw2edSSekgJFL5zLhv914RW5y6RfoR2ygVKPu6tUHM
YfHN+JjhsTwKbtcJ4AND13pAOwNJBxg3notjk9Kqh8qOamOtZm4RsMLdO/LxQA2L
W93iahaIh/9mDd0EGCpaddwx3zn+UgtA2afnwgTmMERh107A422pm8cp0DW1UD5W
8uMtAMUxCbk9CG3B0Tu6Ev6KB+VRD1pNJ4qFErRbRwGBHOCMZDL6ZKC+ipCjcPG+
sJxNoQC5DfHyoarCZZvDj039zoASVNUXfyfb4lsDPwWEqZv3AJHCDAKH+cwmSKhc
zhTM0l08sPvWdyvTemL3/HeRGXgQIYeUORJm20x2DQQ=
`protect END_PROTECTED
