`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jBt8ayAfKilbVO9cqhW059T+kOHNhbc6Z3Zd6UVgi/RzfMC1V3JR6ArwTLWwfiNK
KsJ1pDrAffuiZwJGkkLoNkkpcVFWP+h6wNX9NnduhA75LYGET38GENK/Z6vsQjP3
Iyx/FSOPONF7PNf7TWI+K0wc70NTKNzh2hq84cvq5MCUb5bcDhA6WpR7fEKdkSdR
NTRqn8TdkzRtFiJqPcMimcKrDbOLB/OBI4pq6yCslpz8eAfpxc6io/DCZtP/2N4D
5a1pMpyocXfCr3+DdcLG84zNO/ZbmK2vUUHaPBJ/Rvtrxj2oDSfTsBbihubw4kDW
`protect END_PROTECTED
