`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eEdQnc6F/msK8WSbFB/tn48Lao4AzqgOrGYARxxmtOCJV/h01zwuzfNo880P/P9E
rup9gtRsJueSgH5PF5oIfeqJ/eH/6TUVtvDUggQxrUCqQ4br8KPj39bsI/WV3vMq
A5h0fYKPK6W38q0CE03e07zinx+FglqA+/0/9FcMQi71eGeQ+GCRrXJa2TZ91ev9
dx+Wpn4rJpGODL6jLAQCOhO9NKFusQxc+nGx1X5LqGErcUk2oAsH3ff1lihcrs40
m0/nxDOyCEzIcq0ztpPSEujFHS1gGLfP9vSXcMkioWLxszwK/Ep3pQ1DazDUomUG
UT5L4tDZsFt5mybQDI/OHZqUiDEGa8ohAA/hMFqEQ4Q=
`protect END_PROTECTED
