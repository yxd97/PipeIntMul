`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eulUNllcLzAt+yrDdO4I7BoV6K5+Yh7hPJOmicUj7kD4x98yx1KlyQi1mMlcoLb7
cno7csSPxTzyVyJv2cx35F26keNz3mjr2oT1fX0oS/S441Vg5PSEWtH9DPSoj5mk
hr6Opl2ekKWX/2YrkirfaGwKuzIXx1YIhJI5zRDL6M9HFSTxNXPKvViToHVaHiUO
IE/e1GX21STEJOvITQQD3qbaH84p+DEsQJscSs23gT41+n55dPmUcXVmmf+KwnPJ
GmqEgkqlvArV9foVTL/fJt2CQeYVDx/SsK5WPoleewn0u7pIcP8EMOi+Sqdh8UQe
+gSdax53IKyU5oK/igIXV9kCJU95tc+C/vKXpzpztB0hWOy1rV1zKrJhGDf1e+bI
dy9RahXCXiOogeV16BXLp3gka9mZWDj/ygNUZFxxGFnMDU1Qoxo+JTFqY2ymA+Fc
jehn84+CEHNvXfEaDGeLodjlouL+AIJT+77zI20JJWwHZtpGCDRtOgTWf9Mxyk4h
wNLNZP+LXwyn/GLwks97x4TPLOWq1aUHq+pUEo6RHXSIsSjSQNt9oHyrdJspCy0V
0eqN2oTYj8iC7fLyAUBDa9NsafHfBO1CmOdNXrwAKbaAkev1CQvrv6ZqvuYnEAGP
yGulAUZIEoWK/P5YVqjsOvX+T0zSnuVK7M8GG+HyZfmoEXkqt1NtjAOdCbfc6G20
LZRE4OGnrNFzbCRqZehh9lEbzGaqcKMdhT8KLfYBvl5r+VIRIQZP4fpUCpj8D5kI
etBLfU4MdQ3iV2bagu2ETkXfQlDA0PrdJmyAy64aVE5eA3qNTPmm8FmcN9MJJOxz
eeYUAxSFkGighKrzcvB83ahb/nOoo7GMfA8bIU6VbH73beCemO6xIgjpHYKezQ1T
Lmv2AzzKJMtiTApnGQvurGkAXZ0Iu77CNoW+0bI7SUa0ENCl+1M9EGvmXuhISp0z
5cFyvxFHbLxcafQBYcFj5cZuKPY82bN3GwUhGACQ60PtSEK4WQi8kMTtK6duxrOo
m/j23i/RGB3MvCPGJFksirE9U8LTswCvM3Riow6tzEzOTjgR46oaxzAofiloGKyZ
YqEDxx//ZNbETXmXKnwRJT9617CljCPjLWcCpsjEDWiBj9aPew3epJEjKQEpzxJ1
1ddOqF4U98x/00+o3sbxGrCEGQTbauko+kMCHDTyDJKD0yVVY4zZaEvcmltCXm6S
fMri6ccb01nldbHWTPmeEuMHwFxnpVrGVms+mXtbDasl8YFXDxdHu9r9tt7rTaSs
IcaLJhlocH9K6AycuRJdbJZG7t1snIk4CEulhDBhzSJSjE4+9O/wf7Xfnz9LVja8
yO8/cUrObpZcFowrD9LYI8xiduy2T3kClFq76aWli7YBSVoHwVZjW9xy6W8kAy8h
1xIL2nPVTikMXApGt9bwI2A/RqIDYp7TFPfdl/Nb1rL0HvBGZsVZezFzbzDrYsV9
u+BruTEO8q70jzz+5x2gQC/MC902R+f/w/bxXRiNutxLB5w40eKyqho44ABevj5G
XoJXK41SUbtZpokCZPKNiWdVRaFpmF0Sd8wGjCZucU3Ymprr2mkOGMUozM+HHtoO
NiTDa4mdnSenM8HaQON74DDxRSZzosjNW3a5paPOQFbomXp+P8lWEd3mmkQJwceS
GWfOdzxpVG0cByLcZ2hmjjoVmriuW2itfoeG+PD/8YpBHXOhc7RgLADVAB1uKIQX
XPRjyHQGnXRS8yrXPcy23FWTKGqbGsmktjt1KNCgcTWje67daFeLCnGQzPXvL0IY
BhD+rlXw7T4lPRi0ErYohMPD4gr4ANUbcXqYJHIvl1JwjxUjjrUJmLgdlM+aYPh0
1YtdFLj0Gr9z1ViHkviuLk/OP8fBCtVtj0cWrThXSdRrP6S9dXzOh1uhcAH1FJFZ
hn+YTrjjkTf0qJjIpJ5qMuOaj1gVzGYkvATAfg8MadiQklaY5cjz0RASex24Ulr5
slEybMgT5pO3L8yo2zqNUZgOJJeL7aNvfgMCxXWVMiUhis3kv+1hpu7SfqtU3Fv7
vCYAuLRnuAgIRfVnjKiaGGuf1sB1+5U44atRzQX270cH/N/Jdeb8rvGKIFh20hy7
2xlgzSNSpjAGFp9OMNu21JsrPLHeUyVJ++6HHrN7oI4frC2CTnx7uzT6oRsJpRIt
02Zd2LNxiS1JLBuioo2Wz1nMOBZCJoq3pEawqcyXPnLfxzZ0UQ9eZ86bAL9/o4X4
5hnHoJEMiHaHj3j2nnLU7kvNWIfCdLfENpG8lElRheljr7+Vf1zCug8CuzRC5tkM
yE33Xnb6cVlL5Bxqd9S044xe/7TErUuBp4QE8KeZtPRTWYg4g2FMqu5OvmXRqGxi
//F5MMUIXhyCy+bTgCub+sy1uG0ccThx7d1G01nnCWk/M2PGKlB+FjNTjjMXv68L
E7Huq8CjnkFBMpOMWzKtv4fOlrUuNN0cUgAkuZb7PgPJ4gUW3ZDaDGMOdaIR9hh2
VwoUJQd9OC+LBFou+bBsZZ9ZlGa6aXVWZ9PWUiQiXQ1a6uf2VWU58XMcX1pMWjPa
6NVtuteXFrkWQB9wNkMd7JHyBTmERzyE7hN9lfTKp+WuTfgXhHWhcsvrzVfn9ENY
W8BMKlV25wmYs6G37hqoYSOr6nm40CGMiWYmbMk4biGIzOb0fMla+gl99QV9oX44
OQ2M+4eutx8RZPQyePI6iAq/SpLDfn3Ph/qMvf1Qob5pq8HYWCNdOzxhfHzS/GAw
K2nJjFSfNmweRNnU8Ro2VYJJA+iWq/fYvEfg/oZ0d7tgl6p+xHp/ByT1HhDmOjY4
2hrFVX5FYN0QGy1oU5BOnu6xpdWqJiZu/9YqTId8nfT9TA4s14mNMUqgd/qFWoRg
QupgPlZicoYZvHBDDWKHmdolCtxKioVKGXBVyBvOiKiVPtXB/bIsSSjIlZOORoz1
a860IClt5AQsMY9xd7OklAFoisP7Rd/6JmbPq39auReITsNwkF4tdEeoYSgoiTyF
HgV/QkgS5UkdNx4hnnslZXXW1zRUSbHeuOsd8CiDUR9Hzr8V36SEV0UX0a45bhnv
YOlN9yUR1P2tB3GmNJBkLWAI7Sw5kQ4PCw0CdU3+tdAku67We5rhr3BSFKhbcASS
WmIciBq6n/LvpbaIYWpWtqKAl8toSx1p0sABVAbHuf6Da/bUlKto33HWn5JDWu1+
rHhGibP9gIVZbKY/DmLoG3QMaokqHOHS0EWD6MS7W7Wk2dDxprTmEXiMWIhuajyX
go2sFbtjC3h7fTteBSpJNSM4TyqzaNePYEn+shOZK4uIvtHpejJh80i67K4uWT3k
XRjgDer5D3Gv7slz7B/xPoTldOAKBYr0clbQpBV7G55h4p4cDrxGXKfUY6a/O/Nu
f+S7zwFPUF0Sie/FF9OBf5x5Rn4x85fLPUQBJfJXzOIWgESIQ/8rt4VWHzTcU/d2
SUX7tWJRKJn5T9cMOlaUkN4BAIhBeWwfOzb/T3Kgwg2LZNfG+CnJ59W+Q49+zbju
/3pnhwxySwZxGYXE1Nls1VAGgLMu18FbFKxggReviNckxHg6KNUcCNLLpN2NPdJ/
5Jqj0DcEEhYolVgVI7JnoE0AkbgAeTaxX06jj/jzS0HZlt3DrVI36ne1yLWhm9q3
/TcX3Fav6aLV2+C0zpyrsaXrZF88MuDg+bS0xySO3DJxt8a4Q1sEulbW4aoDwuaf
irZIC5OpQ5DqXFHOVpKmOgREZwzTmo5WIb+hlP4+S0K8eTfTz6aChEzj8pyg+e5Q
IFdsbRf4PirLgBFYep2r0+jsrF5AccfzkKYt4g7hP3zWdVJTzJDpWy1OZ3dGrXIS
slgmfAQ5AYaSsNjtafEM/c/TKuxVDgi7R/7nAnIZw8wrhXxnk1QXoz5Nsgi6U0bq
u5nGFFCPqfhBw9bqwOuafUNhEfK9caPUe4XAqjTx38XYtoPmz0IbBlin9lpxkVSV
JVJOW+/8H6l7pRMW/Sfkf8wHR/VTO6B1HTXwxIKUIsazR7l9jGQWrQiWlidJaQoV
tc7tncLRJ4BlEejwTy16V0owq6T+oRE+MthT2cawf4WXdAqMXIWyEG/wM2glt3BY
843Au8tDSThUoIGr+5PfuQJF0fn503ojGBS/r+7sNjrj4CgjtLg1MBwqEjPCM+tC
tP/zUGHF7NTNlHIBSdQIFm7Z30sP/vW8Qhejg0LMZ9/zvkiYWqZfb1YacVPjzi8L
eBARzp3azkVFGXGKO9bPyj54IMoE1CFr6X5kuWwU5FhdGrk+8PJAWTbVOXY1FjzB
uzDS3696gTckSjvdS3O5yBsxj05FX+z8yfMV6owyLgxzI79GS2nXs48Nb2kux5/B
i4yeGNofPOKswbIvErmuGPKT+IsBQ+BAls+8fhi0gqZyucP1s8LFN2oQcQHb/hM/
fbbTCesaw3EfgxIcKWCVexdU79pl8iI+MTmQBFZs3x6ny/1JgVlRh5ogmO/ZZntg
lUTRMoxWolw+Icdn4diY0UucIIjSjgwUOn9ygFcFrdkvfZYRza5aG7f2zVyjvcRK
6hn6muCXYigfJcfeZ9YxP0WhMdeG4Ohqx1plY/ZUyWY4BVnBScMtroM6wwy62bIk
jtQkboUw4OB0aqdHQwNLrYgh8XSpEtih18Zvr+zbw7P/OkmC/CiKGyGreUc1hIDJ
E1RQrT+vvFGKF/uXHMheEw/2RzbS8mOc6xiDjEYEwAnMJCIT/bKbmFAPNVF/RaRM
w9zK6HL+oZaWXeYxgLY3HdcJLqUlkhfZgs82ZMWmFv07bJH8yTBNT+McbDvEKyLz
4Yks8ycZW9iUo6NO+aI8yN6MLBgGAhia4r2r6QJvst4y2Lhw/+4OBEWE5B06CQdO
rj/x5khyOcEg0XRw85HBQ3cd4HZXoLdEJ1D+3H4zenco37oVaKlX2H8Zk28qtgsS
9sV6iZYuItWOJE1tfE0/OxUjT2stYfhiveMhxm3aIq70dzV9T5R1RtaCECDDcFJJ
Qka+6jnziEhd2FH8KKnE+65x1XS4vk8/wQWdWRK2VekjvayX/hcY2TqIk6eYaZD4
QLMqmSsowLHkW6dGq7mc5BI1QL815+XrT8ff8faM+yHvSbHktg7GDPVLzmWYljOT
gr70irzOKw68qoXQORxsfwc8GLgMqRHCoMH36ScMuhWIPbDJHjkZZcuMvAmgvcRo
rBROKHSmR5tgwzzV4MiBrRbPidKgrC0C+kphHUeP02s6+17bTbQo6yUZmpPiox3g
ZU89cJ/Q6idgRtRV6dygKDtdbXc3vCusaWxiDao3PgiK//ctM/X4BljrFXld6hKO
/TZEpV3Hx9Rt44kPvWT2+oU/nK2igRlpNIYxY6Xq4yCzNRBWHvn4rI02RPuayDjb
XuEy7B1fOi2SsrBltfrjQ85DFJEUUUCD1zr8GEw5KlJdt4gn3LxCNZ+fjGTIgwvm
ZX/cRUbuowLI/rpjQbeszJ5aV2/tMJiwJZSsG/4bY8nv/JfsIdb+9hML+FAX7Aht
ZGlux+Y9adGxRjdMBE93pQkamsM3/K3jphVNsYG9YlGqj+HMIXX8FUMVIshveZJI
5n1KqeHN0d6gSWQJ/oo1cgDXPQcVX3kiX0qxMR0P0EoEr2oWUWU2aG+gupZqUU1q
lZ14XTi6QLTTNp/V68SEtbLZ3+AvVT8+vHUlU+HBpbJY+Z8wFOPBzqwZyo/XK63v
4lgjYeU16yrNLtrWjoKg4A/RuIIYff8gKQ3NYMbtaER/g5mtuuEqK6OyLZLLtOrm
gkIGilBEum1otm0S/BMmLUtS3703VOvepPFoGgNW0OZ2+kWQ4gMINeW6/4EMs2zg
kzM5RUR7NB/xdXg7qlX/Dw2U9XUGGtT22WzFBxbp/3939m9BL4jvsfGK1iFQme2P
kk34nr5tfRShAzhc0OMWxcKMVDTGXxDWzBcU+cW005oQJGn66D4qFSUsWPMomRzY
Vr0r8TEDrGahuLuOeBj/Rcv8MMS72m2PcmUiJFuW/4kejLkKmS2WXlEbrLY+lhFS
efOYwGeBmsKp7y1U4ekc4WxIHu/1hsYjW1R/xTGeL1j1Xns2P0VgbrkhyI7sIVTR
uxGBmI4kLP2eJO6di9bfZqVva4kbWTjFxDDrHtYdNX/+v/mfrkTVSLkQgcHbyuDT
sGOsLYCyBIRVf9veWO4fyRuCmKkcpMWlXgT5mbqoJQVBmFtReKcUQX0Y1Xu4OKme
gYMjKrvXxfjJNZSYK09LMh71OIXelWhhBa40HTA3m56NoWC3zPXA6ZnIWj0dANxI
g6vLtQOTogzGm9eCEYZBurRxo6atUpOFO4IvJpdNsPOA/POUSAfk/ZShylkCSWYl
LRwXISbwZ5i74IpDnjkkP54FGtR7xve8A7Anol9mEeurnR+AdqLUMqSKBB7/qhbq
lAR0DlLjb0CgpeN0tCJF2KjVDcseXz7DHerbpHvv42hIVcL7a/nn6dlW0NvYkgpO
jeuAQZ7WnXGQMjWTu5yaA1pvN+7Rltz9mJSLW5pPe+gLknh1VeGkHZawxi3Adi/o
sSrV4DV8/9yxRGhlvT5o42PyBdUaoj87tKXdtWSLhexGVEjBH5qFihU9++Nw7Kho
XQ0mEsW4bsne4z+I1FRL9sLI4VpmozLecfXMYCWvSr18I0gcZus93ZSMnC32JoMg
3ZRhZd+dtEDQsy/iN679F31EWQiCbv13wzF06CDbOcjB/iY2DDPwNLro63bWgQUu
TpkEBjsZ19psfizb2V3hQhzfiKzLsqeIlrjNGX9oh5Itcc7ne9COyQntpYL7lUH+
YwEcOpgwG+TC8ennMwEF2aYtntjRuaIOu0nLhqdn/6TmSa3UbOQmKkcdUmrDXjr8
HWOEP+Yhd7LVuYpGEyIsOkWWD0MVVE/kZhLenCVoTRmi3NQBZqNkJ/0kFX2z+5un
4hm3AgYJFwuLNT2c/nUO6g4CArDbzP6qljRpoI27RXL8WNRuBtKeUsIGqWD6FImj
a94OQ3y/kS7I/8gwsy16Q3D/kLfawGZ67r2D/OmwxwUQqSg5cF90y0VSDua+IaET
IuYAcRyxSTeceL3mFE3HJeJFrXfZcsdB7trR/5mnoqMcQBLFe/7nMAcKkYOy6Ruf
JEQEUfvl/G+sL0XdVJelMalqt/o5alIZtQj+j0fL4WmHK5R2FHV0PFipfBF4qikp
FzinPum+XMT57ddBPBfyXlnUKVY2bmJ6fRtyuAyxTa9WWLTaJIUAJG5GMmNJeYJ8
h1c6mvDstIxfdjcndjNLPflTdwmbVP/CMQd94+7rAI7JM1qtIAAA5I1BtHr+K3Zs
C2Id/ERZYFy5R2UU3bxsjuNv62tnR4uds8ic+yCCi25o7TNusB5orfPyEZTTNQ5e
j5jvNEHRUNpYlQv92zSS3BMMRO2CMIcnEESW4djPE9Jynf3/UCmMQFZ5IXhLJWGw
Y3vmSb7+9EzIEx5wQAjEYMGKJFwwwGoprLeQIfv8ufS11xZl72p8zXFTf89wEY+L
SIyM9r3twCqUUYrve5hNzu4RlworecclRclcx3OUc5NrWSrJWCKdxo2Ai+/wNar9
iwiQD48Xu8RTD3p+5g+Y/H/Ljekv/6rD88UdoSZdv2kh74/AMg9w0s5WqVdNtTb3
2m2Ap5hK02FOkIct5a2013rJimEgVCKYTcntx4TtFb3XLEQNmBvzls56iK5fJnlR
cj/WXQz32+FYRxBOWJofSs95HQtZ7o54PuYMYlXmSTV2LnjJgHQyJ5+nhKV27C3O
FPEx/MXEz7lipxpeyN+DoHxqT+gm4tYEyjdJihgUd5dGuYoCdHEZf0rQjzjA6Sp+
R/Jq5wHQExeU4AeEKJaBZG8y640AB4JIcHj/y40VVcmAYjV5uHlw6qu1UDjA5uek
d4A7YFC3bFIFG1E77+Fa8SPQDJDH3oLi1lIi/54z0qk5k35ViIVy7q4J+tFvdW4x
eh19fwFOQ3lj9QgyOStmT4SaTmg+qZZptKa38Z7dsDAloHRWYcgcUXfSaEL84L7c
/FqmrUBzRieI3qp7h+vc7M4cOEi3nsn82ngxK96fAKsEwg91jJ+pMZOpDrzBzBzv
z+rPvIjFA3D35yopftcCVMf59uQNXiGhqvdC0IU/Q1/eYHdDomc7QdOFpuYTRNEm
36FpN7oFbmNTlT9HxDuKzQhToKcf5UrLbo+wuvOKdOemn3BPY3QRHnIDX87V36+g
WOYkkAfPw1lQkHn803VOf8gm2IBi57fIjDMCToJN/m5MODUp+Cq5GSxYWPALflNc
XRWrJZkfqWOl5hYqem3tAXdR4lANV4yz9I+ej6uRUezcnwlq0HoK7pJAVaP/d5ZY
BYBwRsTUbLZVKtLmdCe41exF3y+jnO6IgDNBIgyLgqXpdMvbA24m/g+w1dPtfrwG
87WN77A8uX+aQID4VLw/WVjDWJJma5XseWcRHq4GRdDL7UKa7uGv9AMlLCCo1VwP
lzHtMLzDrTEmajvM4RFvFTbIMifaWOxFJkxQYcySjYcPkX316hHTx5cLEtdpCHlZ
62KnRPtmLFg/4zbtVDJyfH/Fp2jR3oDXe4p2+AgrTdnrpboj6edqapFzqEJAdWIz
U1UkvgL7311Rdj2KLEpvadXEHMQLOfb4+PpSmw6bedxiDnDavpBrs9sp7EI+LaZ8
vlpN7z6elh633kZ8n7sUdBhCOR1qPtBveTBflULbNN3uwMJpKSNiq+P4MtH1XKM7
FHlegw6rtIkaADVxKrtl+WdjU5iXd/TqcOwWpZ5rNrXbtg0F6m9UtGLpQd/6HudT
gdSIf8lDSdZRBGo0c57LlmTWcbqVHpE/+UcXajNqYL2qi3taO2NCACRezafxtV4Z
lTGj+DllpnMjruBvPPlMCDNwiBqs+91n1F14WrJQ02jC2y485Wof++EGZVSvieDg
hDtu7Yn22Qs5uxRIJ9PFbOBEAMxZnmDpfQO8gR+t8wuVx3bvxRVR0uf4OTAfnZ1P
FvhvnhonqVRcdgXBbJQGCABkim5R/ZcmRg6l78iZ0DVMblb5dGoy137lU7geK/bg
F25GAJYlBVXDsHAc8VNJupqNeZZ/zMjYKvLu42/dFu2D7PEh+4bwTCmXvQCCK4H1
W1I3Jsx5slinc6Cu+2V2c2Kkz+eh3Hgc/S/Zpgi4Zh8AIBeRjsCuJNQxgPx/LFEe
r4qOJEZd7ZlGW0DybPk+C0WPbpIerpJMr9jOb2DKOBLGfu9wiYGJvzB0dxyYnBmf
vmVWyUH2JNEidxovqLd8BBLl0lXw+qe/MxwHPl3JQmgXpCE+lHNb97b69VBO8fX6
FjObtIYImHu9+wYuW9duucr4JZz8LlyEXrkqSSOADr9JThTmmekfGLFZ/vOwvN0e
frYIQYJkLsRd/R1NY7svy6xrPSyLgeD7akVNxflCNVUSMS6YfHnB3meb6/8IExzu
Bl9uEO6uBZCFnESb+kv08T4c9FjBQLHSu1rAd7xkXlOIsAP4zmv3pVuV5gpNAHRa
YrwzSUFvjqlGaOrlrs3ZJn25y6RZLLHVcJftSPovVCKlGLJ8KEI6HfkjT+45sEuS
ca7eoYaCIzpdy+XYTY9Hx+aND5S7LLsGC8pdpmQRJwRKBiz8QotWb5vDcVet7n/o
dpMRxXTbKoQwGkR3A1Cm6aN/akwhwRYNywm5w5o2uLXoz8BaaTyS3aZy/3O44SDS
Ew14dzvuvXwBy0jLvD3Tuc5SGSwz2Tjy+npY1NNnXyDnRoLxY7toZb54vgCxyHyi
CMqm4ydGUQSmqgoChybrT/UGrr4iW22E5v/+3xm33lM4nbrn9sDpu+aZE6bUdkjo
D/CwLKseMkSVlbBcciA6gd17fcAcJmZ2GN9I2rjqvY1OmYYo/3b3w5/a31L7TVMD
DYcNOS0vX4pcWtZeTWvCBaimR8i5gOOXbS0UCsDHlT4l51amNvV3zA5nQCUVuEhm
0dc/h4XVyVRqfDqYYhuP9SE2u26dMfVDMNYMtg+NceErLcRPj5hnF4Igfcea0UHH
Q9OtjvbkkoPD6unBuiYac9N1VHydjcuRNQAYTgpjdum84DuSh9N07MppabBEsQXu
kRl70FHGMcLDkVh1RUdqie4V+FIwni9a2fOT60RVne2407SmAi20flui7gzT4kuH
E1GKVI953dNfMfoP7hAXBfH7EH1+GAkEN1wYfCxr65z9Qk+d1j2sDUyHdmSUKQrY
ipFnQx9yKqvDTbhN4BpdDankkXrbCBk0S7sJuHUIQT+XVeGJcAx4wZ7KVWPi2Wct
1jTN9mXCt2VgnLYD0QIbdh26OGWbQNWjcdgIJFXe0bdtvk0xJe5nN6pY2ECtBT7r
GzNY3Oo+Bl+LoXmPfYzvqpwKyLu9KsZARQZEVOL3ra7Yc7FLkCVm2U6PTWyvUFfV
pl/uK0CBdye9Boo6PdboBAhszk9taR+R4CPStvJAh04hzojpdkUgNNxlGy/Facns
xLouh5d4U0ZE5hXltbdRZtu+GDnV1LKz+VVn1he4l/KmPlah89Cm79U06ngWFJjB
+Uc0ztIQUCTV6LomAfjllCZIEUhZWLCJo+cE2QH4MNu+GMzRNWGGO+Awrh8ia3KN
8qg8isJAZ4Jss+WjU28MiOcwUrhmLu7HqJlkM3C7wmY8CZwcmlr6Or5nAdtuC64Q
UfAPppaqD9EgWUKcshYF6TQ1+Z3mlWoklB/s/+lKZOjLr74co5ECFYNpoIpFsU9a
6fHOmahYkpczOP5QtTsye2EIoxKMCf/+0Tw6WPObmXU7AFMOH/K68Wtf2VGa5Ll8
LkHbTmtLe+NiHDlFmLv4zY50MyE9bAxinY8nW3cyXz5yzm2DLdjgAdyDWnG9trzr
NaEjJE8QGTC3bjAFQwz06yOStXRpkz/8OKI6AttRZ8KzsM6GXUvyBSYy+fF3JfnE
gorPr8yi82eI5IuiiajCZm1ChH9w8yc0GWm2Ivp6KxjJXilsA+iCQlLZuqEDKvnJ
d/pYPkAYGGCyAZpuCWy/0bnJXAgbueqUAoZYZVDFvw91fFILXKJV61F5nWUtAus6
M7+OfMxjngBDnMJbgdEymqBqYksl8S49nX0OKAYUX47IwkxH4V3qKIBdXyN1yMtD
KdUvZq+/dlGwPBG05NFqZOdYLKdc5VXVzFQGFv9DM+KbfZ5rcK/ts00Ygf7upYpy
Rqr8RTnBcxi25poTpzyvXMmBK966NiBkWsEBmY3fBZeup9HX25B7/ZPGm+34CoRv
PF57Z1OjsRmssFue7/wXrbb0RZZlBphswZQDZigfwm1JvY5k034h9iQu3Zhp7BlZ
SM0n7YpaokFIDT9Jv+/zgfx9QLu1b58vLgQVZQS3mvSuaQVq4QcFEx+UVNpZtaDp
F6iExCAxEJXo1FGNwVca1d3iWhpCYqZkwLjDegJoEye4nnFloOWVgpDID9Sx/mnI
WkJeUR9TnupA4w/kB08eGZPtyWY7kI8Uftq3lX0vOkUExEq6HIfyT/HCW8cDT5Tw
q96GUJrDr0xFRyvDVLTdjUvWAXWOt1/mO9wpvdHjdDYielzPOFmDcN6PiXanyhFv
Mknpr05Re1mOCJj+TjkowTmmttsVlogdPT4xwmcVkthJKuF1cW3yvJQUn15Tx/0A
/TDAPxEZV4GZefuV5UATQoWbmxp1V4owytmrltk/09MVxBLVeEIU/9TGRcNr/Bo9
uA0pzTMRJUnkkoUcT5flQ2dJi+XRS+0HPNllXBcp+daBDOlOetwUQkXDfYywM9GC
JBTVjOwnwcnbtJSf0obMtOBsMEkigpMDa0YDlLaQDOyz1uYBww59T6gO/Tvd6/Pl
CRhtDLrqWUNgskpJiH0oDWwUkwsZGZ4vCTI8FZmtXY38ej6mUi9U+ry1NoVwZyBf
ZWgNyJn7ZEHrw0OaY8ZAuzEHtyD+tMv0Ekb+H4JRMkz/XYpaLOlvPDbFwYvVJCYp
coHcfe4Vj9IZbXIRxj6ZSpMqn4osQNjPXnhb/9CCd0jUcVOymcVlgiaNn6j0CLVM
vXirByT7u1273B9jdD3fUlrGBjMbRS03OOw/1uC8d2LB+LdYG1Htg8PqTawKJ1qC
bESMpVYcjLkUjIcy8d3QZz3cRIK3FG0SbGT8V+pqRSiIw3Zbolh2N2jruBKWqHEq
fYCwyFRXNHLbDsUDPDl2/YVRN3jfepm8Wg6sTN5rllowvmlB9nA4VqjIIJ1TlBC7
xVNYkoIa4DFZ0vosCnuO6c4F3fSJdf0G5Y+2avRJGQU8451+/23mMHLyKzNy/y7y
Hrk7pfBil+GbISNO1skfyoM1VjcuWDyGfMHFbnKpovZMfDx7Zaa0v101azI6dOeD
9JhjPoSurmjwnKYPJzUhkiMNqwP7iBl9OHHhfnmxycwWlqYOeU2h6XJou54BnJs7
wLPMO4QzPTtfIfYkDA+hItlxWyQ4Jf+ecxV8K4qIYHwSuRXG7p99xEliErWV4tq2
eu5TOHgiDMyqj9OUOPNfx0anJSvUhP2L5GWd5REhtNBXR+Z8K/rsSWfF80ch4y/M
kJMHhOhAi8N7n4Go8+gOTDuptDtlIzKY93fJE83R1dhudji0hiOuBKubiVadhqc8
YOdg6e/uymndedLewPqmeLzmR1CNA/UHINbHGrpT2dDyYrPoSI8IDqbJMcOGHMy2
QyI8g1l2lr/hypqpujcWY0pH5OYu0VzC8juQwbeZkNBY2duBl4pVHFQ+ZIcoMr5S
FZNdkymkc1DYW/2LwYkldxf8oKMoCIehkmbBbjbsogAj694SLe224GMl9TE1f5tr
4DZ2GS5CjrgnFJfco2NF7GJ3eryhbQvAFNTTbntQHoMwktlDERU2w1AKpHsi4rk5
US3sQ0GLEfogoxXFg9KLxLdw7dxUSIiq+5xoXbpGnMpWGc6Lyx0kP4tirTy/zmt8
z97Src0BCFPO9w/g4bN6VDjh9sFo1iVgaZB3u+x6VwCdZkKLJaM8yqvIOX3+LCfO
RNa5JrWMfkZSH9wDO716ZF7/81tNc3pfXIVWR9S7XLGV9zXRegn738zFql4aQ6gS
8NB+EqFnSspuPxIlBnW8SfqHAb7khICYVLzxa35slR1X+FHXqJDkGV/8SsYjDT6O
liHmxCKJCa/vSTMAUB3hv5GWloqMzusqVIN+FeYEvqFz+XAUY0UkgmrI4UQUKqEy
0HCHk0J2Wjrrae2a+jGtz9tlEHWCEBe3a91/5OfpjrhC5+3qmVmPpG1pF0x8uppr
3e0I7reYdjUJaMXAB/jWRyMg0kJU4VXQgLzGHUKzHFU5vRQXVBmg3TqBWIS7JV+b
t6ymtnR4y5iltt2+atiV1yXyxNJE2u4VPJk5gznLBb9RcA7vNPB815VUG5o1rNxS
KLqGSEz7wcH2M65gQDnRA+ZVIBJN3XN+lp+D6qqJiG6DKsfeCVT44Ww8LHA5m+mf
lCE8NDS425Hc8RYpXKiInHo/+f5ITF0F4g8bJ+4qj7tzweEjepuG5EFy6mOF8CcQ
mZLuPOoIndm2oYn3LY9Kku6SLw35mo13E3UkNbg0ZYgCoQ/Ah4lNxHOccI1+PFWF
1ZFcpLDOR9JI9GtlhoBEk9/XgLNVj74Ir7mA34pTIe/nzfMwJAvDyHA95I8DqdUh
dlf/y8SgJtRbgFtataISHJDWAGrzpE022R0+MBkP8vRtbNTjwn+4Ur5TrM8Pihvs
rdt68rDZM/MFiR6Sd1/swjvh5OyZ/a2L3sMsm1D6aLNFGr/d9PVTLU9jEIzRYheU
d1dN40Lo94wVLKYnb4UZdE8SVNBH+ANihtGOIBLwNc4yoAyEWaSFY2eSkgojePxJ
Dmm8SoUJ2eY6MTArda3TJsECf2MA7NzQa7JJJkWdQWkos2Pms3jZspyxQ4sW6ZSW
Wzf6Jn3wkKZay8CwaPDutSNYxUcYpxrXPH8UBevan1Y72OnJQMPIlxVkYWKOJZ15
aRQi3kEUKVqGnVJiMq8Viw0r51w4AkHD7TrmKzpztCWnUKnlRa9Z83PBY7IEuYfN
goDJ+LmXfYemFld2mS9QhxYPJRon/a8MjQ5dc4xN3Z62jkk9WjEaFe2iVVGLS2ez
0ZqkIHm7bUpXUHHTdy2ZCgKgF7INXFfaAS/L8i8va03+5J7beMRPVbZrV6Hgfrt1
GBiLsyCtSJrC+MJk1GmqHj+zqLwbOlqnkZykRvLknNT8XoNKVZcvKNdPZulTEaxR
zUoigKXitFAzvFIr51sJkQtg+zB2O0JeTSvLusHbAAJCeD4fK3g8ZGKLoqbJuPHM
5TdiWuI0/WnI51xgiDYrwkoZnybv3BxXDGx08pOOMU9mzpVCBXxwzgjH1Msjx0VC
ecoBD7pkiutuPKVxE0EMz/fxMlTmYmzlf3+o+7IdJ7JjU2ygTW1mXawE9q9RFFU/
XuWm0i4AECg6pcqEhXAhoeTbn0WGqija6J4jgppOz62zMezwWHA7oUoZOGz871KB
TdTVNKVUR9r3/BeVr7EG+xgwLKMmbZVjtZiDEpE61y0Rxv33DUBsRcCFyrb7r3H5
G4YbgcFz93QC+ZgjbMQ+L2jh2a6RmZQ4tBZEPDcawLwGqNS9f2OuDYFXc2cqqlk3
qoWiwdXjXPxw0mgdR/B5xC/vhHWQXdOaztOCZ8FI99q5NgSjInxi7K415Mceo6DG
eSTDjAKkRQJnItxaebRwJKxwmRpzHC68Oeo4OUaif8ugOd3HXebMTre23pjJPyg0
JFYf45+AAiPmFFjf3rN/ozRixjAHYl94iJ4Lg+U6glA88If9CXnS0rDwbcEfsX8Y
GDFxegw+QjPNJXem260lvnQylNQbfWcTe+U3Y7q5hiELIIJBZjspgbgjR4jGCeC5
b6eB1f1uNZj1D5/BpZYJQOj9ldjBhYjB9fnBFF8ETfHVh7bkJuM5ybR3n5L123Wj
s7T0MePYBWmb/FKAItCrlbnydc4Yckc1qIe85avTDkRpznqvdt0GAFqwy0aQ3DlI
p1F9+8SOzc0HviDprpt+VOYnmJNMh7f790Rv29qqRnibIzD/33ycgLzoxKEuKxqJ
3pwKwA3r4s9o61ZtTBXqptY3rOev0E3lTG/SbGH0fL8Hrgb+hMQAyaMUKE11JMMQ
L8shEmRWfOfF+SR0t6dsu+EIjmm0u07dqQiAmncumloNP52Y3OYBTLa+VKcLPuMm
eM47nuzxBkrMKPBhfpI+CFUxWRdk4j8LN3CUQt11vFoL96JtYRN+GrjPOeJpzSb0
CnR/l47al0JWiqDhlzzwvBiNitEO5NhDM4BMZB+LbEFmqpDWRxab/RkaAqCLp2uf
c8RCZyMzIkDjwOh9M9zLMmR7Pnj0kdL4nst/2fpnHgXmhBFSA+g21h/de9qNat6u
J5Jmzx7YCS31gJJEzWuMZIa4J7UzTl6EUxZu2h8mui/tGww1LFo11wVQEQpoUgA4
7D7RAz68zdykQyRTCED2kvmj/oW/co6ZSMapqi7EOBTMfzEMJZaV3hoJ9725dn0m
ZWzZ5jb62F8MpyDXrWqOaxg+bqgnXK51IfIVdebmgRbimNRweYk1DU/yDENVL/Me
MvD0zM9G/RYulCUbJjcaocD2LFbntyetlyePFzdRYhZb3aoo03CDd/yQoOVV/Apr
fEnEhOL1f4vO9QIFB1+991bx7xeRFwzoKPf3oiZN/qG4bxSVv65IrlaVvJvK+W2e
rxnvwGA+rS40dpaktuv8xrtDTg/uRs0cciNUqeQ/OwiFwDn7Pr54oznouTNS4dea
7UjDLbiBmorgxJuIbTmvbILo1tNSb0Be0BWQ2LTzke4zDMS02e3h78lZcAtb3PP7
lWxc65XCNrnGLLMpqkfTDcQ+6R2V0LjzK52ttl4svmq/Qbcx5wA2Eb2S/GNWPSIE
H1uN+FNb2ZZo5G8f6/TlAbrbTSoTyzrZ+KGQ3sNSw1Iet1iSIheXpbWGDz9H+C2V
WTujjVn1OWHUdsOhjC1LKi/wNtLwscP6/DVWe1j9Yi+pebUZig1NPbxH8K8xZMYB
nTaib1TKQsyjFOD41zDrMLyZGvxf7GJ/Zkt8olkSiHJzpIrUq7DTh0bVqXmo9yi/
4L7WRbCtSCbfR+ponuHN16H5hv+fR2ytJPDOMG79fQ9IGrFq1QIkHtzCsbkL2egf
XU5guCAUfd+o7GX7NPY9eMGr34HPG3fzuvdEcz3Iq5xMvqS+zTovcJ42soE/PeR7
I3nxuS+9dGKV8OwZEdJQsa42A2xHeaW/pNrXuWuFIWXkAhOnPUS5pEs5XABnoCH4
rP3pxV5TlSNbT8FiK4tzaQ1MggNf1Mo2ghZbzvcGdwRciNJzjTMJo70FW4f0YFQG
VZm3kUizeKmiIevXfUTKjs1qxSmpe5kNogGxq6Oe1/1G48s10/dxl7n1P5FKtIMt
sq22LXkK862jzzB4chHiMz+PutYrZF3/+fVNp4EdqjtNhc7+UdGLbaNRHqRlJvTd
qyhDu7AFc10aC+O99fE0FojWvS26LHYbdxWXThMryT7kpnv6H6FWC9afyJcO5iiP
EXp3gozlRjdraAXoZIJzD4N0UjWD5vJEsJsD+sLSW+i0qxVlx0LWa2QTl3rCKpS9
aJqZ35kbICIutdY4Rk+ZQbhbQ/Pu3tSltOFtgM7dgmdBz7sCmCxphLX8GRvYwDBK
qC9M7hOhfxI5FrGCAbLSqTwRbKDV2MkXsbApE3l8XJqyFIxW/xTMaRrqrTFrmEna
MuIXeM9nRW3g1OgeeWFSVk2fmjuL3UU4bDENn+4/lCUZGeSnNh6O+30RK+CNpj+C
zU/VS7XzVFSFPrSoVA/ZDmgYstKIkpsUPMoYWRX4/Fgh4/XWzyRjB0u6jCGYCk/b
xHgaqldxdX8RelHVd7UI3YJK1IU0KFyw77mSYVoNOkIS2bQOnlf320uYm8jyp9ea
TgXvWtRj3M4bn+fSGt30KVXfVQSqQsMR7dK+NnYDmoE0UgrLxtHi0GVsQaVVFUJA
M9l3qbOpZ/U8BA8wgzAzwq04Koqsrvq8YMlJ8rk/+spWLiGwhI3TrJ9TG11ygxXK
lQHSsr6tckR0XmNIzNC4OPoiMAzPzyxuVvQK/WXsbLl49l923pSER7K0viNwN1AD
E2E8O1P3z1cYJ+JOSlJvdAm14DNWYJfwKVQMulhuAFzPRSLV9mWE6v0Z2SuyIJOm
llZfYTEo0keGFQIdJbn8TJhqW8OcvEh8fm2Wq+AKDuraxEQW7RwVl09ufuN7JSJF
a2GytTknJ5YV06DClMqJNQeve9/bcw/p9sDaebZb17JA9QXgRp9BselAuJsM+Yak
7lsp55nQA1ZUcsUPEN7E6B2shAeNCiPysUcD2Mk7xKqtkiJmwJYfQ2M1k9yvborY
BDRSYXbiHQX2c5b3vBwPrYwui3pz6z6BB+IwNd3lbg3jO9zy/TE7VV3D1xjaXsb9
IPP3WSzgggGZtG2iuXxztGBl0BRmOXPRRiY9xp6QbQvuth4RXkyLnm/U2Qg4h+91
01B6I8+zu1hqFx3uHoGVRqVJvIIXDqvWSc18D0+QVYrIFBQtQCGhO/qXdfL2b0tJ
4ssBsc1XTB5OgToH2y8Gt793RxJWQ0b4CicleFhtfHT2PAjlr9kDw3yzzywvFgPI
gQXA6DbaCJHL40cgaQuTo7Eyqnjh57eb2NkO2aHzsr3Qvu/Nyu4lJxRat9Zon9iE
uLsVnLYKhIf+rSxDoEjRAmu80C2IEquDgnItzlUSOSm1a+Uln2G2B+e6z95SonZH
Ns9B5Bbfty/j819sKoKsyZowqfhTlt9tUyf+cOCCsGAa5OHcwp0o+j5LV081AehF
xAz6/6PBbplWEqqwvXqvIcMYz81I58K+4+pVzB3DXfLIqEGvMyLczMtwImOa3vQK
D83cRwSVY9H2Hv31SP6WPtSLiSBwPBksa0GpxZS25mR6YrkgiiyU56ht7plktu6C
ssIB0Hd3P8bnjwqlrr5K9t+1I2xxnsNbdkVsMz4l9HcvHw9QgZrXDTzHpgIJJVcM
3Gq8N2JMba5FCFwMym7xOahSyfmLRq0bNubRGVa4X2lNHuegpe/eim06rZoH36wN
6GK65LKWdcfaH4CpNPYf+KlULWLvhe5SSSYYSrSWBJpwk/sdraWKMc+ucPRBD1cp
+/6WH5jm3ipdlKY7a7hu4y0OD5SRaCDeal631auoFJf16oC2r4ZrQzSqsO1+t6Tu
m5VVK5Aopc/gFSGg4RPJRh8blkTKu2l2krsqHVqOx4T4mQ6hT6yAmCEkTGF2YLj1
sCBPh69rAN42hhHyOofSsJMSydh5EK5WfxmO13aHJCHLsLQJXQ3JE2v4wvxr47XX
PDB+S8pWl/DjUz0I049VJbfffv8F66l/fkIdK/S+GyoLJF+7vo+LW+5fzF9GPkoH
3rDNoPjPzu1Dp1ye7q6spSZdIayRFFTUXP2A4D8+x/+YyIazH4Mf9hQTen9FVP0m
okS9c1CXe+DRGsg1oaKuI1qz5zNI6hIPiN3qh2n522Ws3ivylY3wv4lwNIq3lDQU
HwWx4AGiKCxNIPQHc8+HTPMCmfBxXyZ/5DFAcqI0BdB0k8tgnlafYtC12WMCkWYq
J++y1ffdkTTIqbVZIRmk7d6oiBWd/hoDgSGgvNImmjmC41Px1abJvUvx3CO/YmF3
BASbycDUVCGoiutOKoNhP+iuNnokgjgwjGfa77jA8aU8Z191NfYNE5DSzMGtHPfn
1MKBQ65mIPocpAfoF1ZIqxphHA81dpstRfzSSZedGonD2KWkqUDFqOAy5ZIClRNB
awQi1gcESIfLk5IzSylyzowHEV6JC7wBs1uDw/2DvfqrHm6Nu45DKIBlF21dyTJo
VlYbzzyhXP1DTDLZgjyAameB6ITMntxNIQOfLjnOQj6m7Y8NLZIvJZC0wbYD5wiW
ZLr8XYNAVsp/BPd6E3WcpdUKapBTdAhXS0eVoIwrDx7H54UyDrvWVzSi2hbdl+81
V2hc1FilgQaPquPlGx1rBItamkmqbiXkwHgPLkjFRgLbmgUTjW4hVuACdyHl3DM1
A5hjv/KxeZ83H7T//zM9olpuKAVsmA9A4Nc3g1/HPG1+xcQTUhNFtqg4jBWu1P5M
Tc3Zp8UYkOBBYHmNah2mg4yBUFdu98TxrFcWbJzEAJj2z9O0NupEB5BS7yeqPt4k
2icTcQ/2MTQxjo+9LjwfKQRD3IHKNauGFxqDvIGPeaQ+pfSt9VZcAqbUEcpBw527
+OV1hPr9ljrZ0e4y6U7sWMiL2/G+zPeNpTqA3HoS8BMWqYiNpONAoghstt9swri9
h4KFwBFdsSgPgOtuuw3Yqavnmdp0zyyp4UF0RiOCMhAx23NqzItmAqqM59gxRnw4
pOU5IoHXom1Jw7Dyi/tS0m0kCJZBqlvjYQBf3RpmOgIy4a3dJOxlh0j05eSahxdu
LaqjhMF7GpQ3zn40jDbqycJxe+mhjE5xBoQd79Fpk3l27hRa3sNssS/kDFwQ2BVE
40FSHMeZ07vswvM4QwU47lw4gekbcWCYteMfpow7JPlV/s4MikuJJHUxsIKjojEF
pSTYohLrPmDt27KFM4rNAASFJRGbgD9vW6Q3pM2GUKFlaHxX6c6G0BTckwpT/Nm5
oNA2qxdVpczlRz79RNHvHt92Q6p8A1WieaWguDxw+eHoQHExTEdZyfnRCt5qHzh1
Qcw02uML5HipvvAAcjiqd4VBqt6QElcHwiQsRMmKqi78/7zluIa+ooZJL0pRol3C
5LYxolz5z0b2K+zoPK7oOuFmHzB5BMzKj0RVdG4D6PyAWMfoxy31I1gas/2PRnay
a7HQJm44UE8NM38GI2uR1bpGHZns6LiV/jRInIyws55Wiy7OAAmS+3uajglEAtbm
BoYmqalc26r7Y0qP/AR05EjqyFV8PJE36as4G+neOyE95DSUxAiOGb3Mts5K42hv
sHDs3XYBAOqvensHYafqjeb2fluwaeURlHQubdvWk3KSPfctmMLR7rAF+p7kX0eV
O+5OJcxlX0f42xpruJKomsDT5sd8P7geeQDjt7fmM60Scas6rEaT4z4ub5bZbXbF
U8tvsqdQxMbg9quIcrQMomYj6N6xC7kXw3XAInr9tctxjSa6Z5TGft91EFqmmBQd
zpmGM8x4haunAxeZz0LcaW+SkqagzwjxcYL8TpADMYQGd+D7yz5tUWurYr3EWK0j
nTawGsjhU1bkOkrEMebMZ68sjo8S8D6MC5ZgADxtUfH2zzifEGj0U1U183LmZE0T
9fpWL87W1pY18mTobC86CLlTqgTapKWNtF5Bh5IuuY8Yiq3Q/GKGB+Ggocl8GTeI
HBQZLHBM3bW5LdxjEbgdvbbaJE+dgxPjIwdm011gxS11I40ugHv5vDv2CRJKZfeb
ZabafoNzcjvt8POGG5COs6nRf/R/Pikt5Ijjwtq+LN4uFTHUpjWTkyCdXXdTTMnd
lqY8PNnYGbNQwDJnMBy+q18KTKzfKvGZi71P6fP7PFWcGflRwzQyCgQS5b6pPgjf
gRL9fkF35XWg40OkgZPykaCaGEsVr6G/ycFmJmJkWiQ1pPqvsF19ojbv0+/GOi1Q
+WUwfm2iheTjVn7LqvL1yr7FGjFXpyyW/L23GhkHEhbSy2bDYM1JHykbe0QAgTVa
QypTRg+uepAGSY/wsdOP1WVgE42MauU3dMkU3RzK2CaFCbS2jRA/PaDTVYpvkMW6
iPaF2vkoQUwN5vS9UZ1dCDhUsmrnaHcZQBsUBHvpF2QkczBkImphgfnAvh9Z3Oxt
0LGpyWJJsl1SbkmvaW71umt5PbDIBzXC/CUpP/mjIu2h9ZSYRjaL7MbZzRAfWj0v
d5JtTr+p+XzlhzniYzIPQClDf9QqMqUKR9wncmT+BZqfKufIPcLMoJcr6tY+msVB
d87trgUBBJj6cckeVeax1xDHdrmm/mBSxtrXHSiekPap+P1Wz5QRK5/hn0r/ceAJ
eTd3rk+OdtILcbdpSSSSmhv9ADOpbCsADpBCBj+JEyUmKqqa1OyMojamF6cB/BEZ
erKS20Dz4039q87mORJLSeQIorc9lTtDFlF74t0yfC9hMvyC4bNIJuA0N2wX2Owr
UUuCI9W0/Q3naJs5y1izdLYxfOsm7t+g4ogfNJd8P1oObSp+0QN014jPRbkdqX7O
3G4p1JmmK4Yy2FP0Yvc/76UqzZrIrMqMTba9nDT5iYc65D+4MflW7rgm94dZqN1M
t5XoYBwBq3DMkvvq741b4CVgVZ5hOvwYqhtGOG+HbiWsTM+a69ClSNy/swbcPnBO
YusbElRMyvi8KrPXZ23UZJFJz4UeOEEZ5FiOf/eKzBdMZnMHM2I+XFpvM5b0YxwN
h14wSmJm7OoAQLCFVeukgabqXqUXCJAnXjMXsJL62EwAWkK8SntBL0IBrtwqu2m7
5JGVH2XnrSMom8ui3AoPZPI6Vt0uzh4X7jbpGxWB/APFnEI1hcDg+M6COuGAsx5L
px96/QV95vfwi6wAjEVmPeYRmIWiQD2sCc07OWC+a5q0ptoBixxUiupbN/A448mC
BjaJGX+maoSrfJRL8AhnJnlRmgQflQhfuOfuh8MpVwKOkEj9s0vyJWvRLuT24rdb
nqtPl6V4Srk4Ve8Ka3sye01yUBhcK+PdhyUuB6rupOzuKBEKOvnmSKJMuZvSwbVJ
u1LNCHEpU8BCA7+DqfcH8rNQ53MSV6ccE/VGcnqEIlCcoqHJI8kRkhmB6ZeJ50Dc
5pURXVNty2zRUsNzNwwDuT2dESfoziO1YP3aCw0xZSsziGTsVtSzdWfawAjEJmpz
ADiV36mBqoUlrrIBm4Ir5QDXny3fWWzr0bVYD32qwhGgXppju1zvy7Ax3sHPS4HN
qPCx2br1PqktZ/7mBhtSKO/YqNGECc7+p9iwVGIop2PHzK7xH/vDQ9tK3lojcycr
3aa1PAlKf1i4vOLMAYBq+mDAXeIK7nrE9wfSobPpyHQNjKoR2Sw6j83ppIkzykJM
7r2GzGQBtOi7cIFiFFCvieG1Z4hRR/RleYl2M3GQC2nTa1CBwuw0rXZodNTcGugu
dtdDQ5suXKfwHe38pF/ozA/fHMk4JLavo6FOrJF4fDVn1udqMrYj/QrR/hgJ0/3u
yCgDPQL0JtVm0fOPNs7lYU4BklM9aKv/34sVJJVJI0vTx5mmTG4xmL1N+Ac323o0
wHzpWvSQNUVyqkxNTEOB8Uz+NfpqaD+orgjdcBnOPDUv36V1pi0OFBM6B2fDoZ5w
M4oK3LMmobaVU9MSS+IVWz79eBRn77HPOfskABlrRNDREtMRPBqYa4nddj34k6mh
w8FQM4Q61iQJoYJqWoeKaOqvYv5yB3lRfEqkUGjzSzhTNKBIF8ncsJ/uxVgcZl2F
EI6WDPhvaQl1jzHw+vapWdqWo43p+O4hu7xrPolGZOLx8VyHe7mSR4NQmfRxMj0p
INOY6xsnajlTgXwRiA2Lkmh4KObR61JfHZsNCuIjpROJ3AT+CTkbDpVnsdl6uQVU
C0/u8q9mMItdvlvwUMJGzpN2juyyWvLX/NItTIOrKusGVlw846qsTicfJhbXGzxC
pTAx5cEvosmQyFEz7nIJaoHhqDbdNsfyriQ9Q1RrPfJ5kEO9h1oTbdroZ0CqC1E7
a6FL68MYp1KRE+O6AR4KP9AZUw60idbyb6LXRrq/HgF5s17S/EY6F6Kkrzxd3B+m
LxlfJG9Hp/a9V7mA7o/FWsJdoBh45QdAJ2hvUp1qvySxA2ujGEIiYYBu2BPflO+T
cbxzpsdM3zhWNE25p35cLCxsSfeTs4u1OVapCv0iuvV0wZ4klEWeRwfGbshg9+7D
C0u3dHlWuQFmzcbet5CVdF0Fqb5GQaezpFSG187Pr/qo813YRSOblON6x6J3rH5/
HEZv92XK6PDqDInlEz6DgUpmAJAMiQ3RAlWbFmlgcCgk9CpSyH2nVWMvMDKxHodS
0ahwPxePMl6X++buw4r7Za5zgwgcmaNLYkIyUdnH9FriI9xmZK9mCCoWFMAHSuj+
aVLXKNLDm7U7ee3dZ+0WaKu5IyHBME5la7fldMN8dqLbWyT0HjNHOFNTBDjrjxYX
E2S3vPVtY876/UG80sJxjhLghsHlC/SvhiXMzrzJWCFXRUI7DmHz1QD6AA7MhHAD
pQqnGJb/EYSzSlkmjvMyz5XALB/vPVrFxxPpgQ32CPqwa7faAM5bUVRw4pAu3suv
8Ztj3lwOJs5Oiy+TR7dGMVDiEaQAeXRng4N6VWWz8ZTri6IQnr/pez/9u+6xh4yO
6otBHecx1OiyIurlrEuMrORraZgja+6eQA3lanmw7veo2FUQFCs4az74CMk892WM
QpeosD9wC4BjcHL9LY4xrnfN0YKxXQ7OXDS355TwJVTj/niTCxFq5WJCYjmdyitH
hapfyD4DQC+mDQ+5RNMNYE4maKIF7sW0KzrQ+nWpGFhS9aBqJw+LM8Wn8aYbqBS8
Wr75pXb42HUEtjh6yWab+uJrkJLr1Et57j+anJ85wY+fBF6FlCI1atG6NeEMZxJK
fLUdxYXnyKQX8IEmRZDxO58XWcxmU+XLQkraSUGMBRoNa3VJ3o+rwk/TeXqfExKd
I2O7nxNay3Ih+wAJfieynpo8bLJnbfEcgVx0zyorwYM27wyyFHk5xUBbK9MYX42+
OV/dxOuBUaCIKllfipWlEpvJIgeY7NbP3UtJT9Th7oCYsoMVgZWH3mT96qSdv3tj
nx0SKOH0J3WX2xjQDT0bIjMuq9ANLHJR+ugPwC4lU3yleTi0ekZs5e/oiX41pZa1
gzpywMPKqP1OFtoSuQfsOjkXjefrlv3KvMiAMGeMyH/qJ35giG6r641Bchw2W1yz
Uj9zIVR/jm57/n05VqhpRO4GgijBXgMM03FczHHti7lh9Y7ie+fcj4VTO1J10lId
OthjduYPTSNyAdO/scKPLW++JJ1wVG9IVbhU0iMveh/33drb/lQIdIgsTtscbAx+
DgyhRBd6Xo36pNcKTsAaNgzqz3TXteSU3RPcODyVnKxfA6ngYlo82bgtmbVGP756
O/X4SlgDIV3DoqnvVwEkF430ALJAAaDuffww9mF+VO1dwOqJ7ojslh4xADMUWcdE
GyoTzvxqDQL4iDMS1XzQ9dBX2ag3IipJVFK0qtLx8VgB/RjyprwPyBUn6kEQBgoj
XP99eQYCZlyWXHpQ+930fmUlg3NmiRaCCEQnb5uiFSr2nm8Z+xBWvN7QKlSuitnw
YzdhC5Y48wkUvTHVKZHNOpcUrCFEmvPFVWMPDIR6VqJf7yfO0SUkL/SEjV7iLe51
ff0RjIjk36kLzhIJkTRxo2etIQugPp9xY2iJcUXWb14InU1zG+0mNmUDr9zi4NcE
rqQrFOVHfXbZdSEKDdDHmj3fRlNPKNzkggLCIeLZWLlaH/D7NusGFy7AV0IlyhFm
NkP7z10YhMrztZ0MZvjQEw8YH1CKSMY0zYgoBkuXbz1pmEAtCx1osA7aqZfqHFaE
GRbyEQH50n3aYKJtlceJyUydiX8Jraenazk4mPrbaft99Ylroi3JwSfKtjHpkRyF
KwLpCRbVtBxXASwr+OzcW6LykoaEKXpou+6wL3MhJRFqXX98dfNaKUEqdoJC7Nym
I2EKLxcr6DnA4x39G19pVWpWc2fsKuFmPCaSvz93qB5ysAKJQLoannyHWyuhcQ4M
Fv5jm15Qhh3s/l/+DFA3Hrl7xDwFjqgaOEr3Cm24rMVW7DKU+niKEeIB2WzNJNil
kxQuAQuVTflJGhoKYrSmLGykBGDKPO8IidS3XdAsW6eMp+2d9knI3S9trQway6NT
3BsJOddEyDnBq241v2lV1EOfT5XK3lnSKjh5FFoxO6BZ1psH0ZyKFBVObb+iw/TI
uyzi2PJspYOsHr7xZbdWxf4145EtMk++07ysUXBuSiFvnsJ0NlPasOj95hpT0y5A
QsmYNSyCb3hmJQ+6ErOR+pnEURca5udDovptbMvCL4MJjwTVQuzd+C/HeMh18s+v
ZRCXbAU+YBWx2H4QTLxBzXCTOuBkS73e9/oFDfbLhW5/qzo4w3UjeTYZDifO7bLx
hkb/U7W5TYyX/tWa/4MCUUr4Cn+S8uUAd7KpBJe6/5JWu+bldYB4TiKF5D/jhGVO
oZ6qBi1kSSaxwM3CBhEaOhWLCXcz0vGs2UYXLf0VwKpgU2cXADHpX9fdH7/2kZ+m
aY1f1xa96fpTLd9aqhoB3r9iW91V5GHFWLuCjwRL6aiVBIvvXBse9t2Cm3tKNRph
qVeSvKbTLRuJtF/RgW6iVSYrFen+NPL4L49t81h8TC5JfUymj25zzaq9ey6ggto+
gXLNBaa1ZXLTBUch0H3WXUiW4QJNbq9UmGYs+s564Fuq5/7U5KdE/pUdCe6ACgDx
xKHlUhq9C5Wv9+pw/rerbQ4dC6AMNV2VEVFQruDAYtBHCHC7e+ZXLDzfIwp3ueKz
1EG4HnJTOaYbXsTUs2vueWfBonRxc1YgjtdX4kxJqqiKyDJs4D/enRyw9uxqcEpO
MJFnFR5H9+tr3zcvNx4giOB1YLD3EgC/ogQaTMPBgdPgYvPjw4doLqI2ZICd64NH
dY2KNy56nVZfR+Rhh5WK4m/OYJNmZJwrKh5D87zCdt5RaN1Hu0i2qYdJKMKEPzSe
d+Ao/52CxVbNadxV0g0OTdoM/kUch+hXLfrkjIsaciWyUno5EyxEaaE29KE4jlQa
h26v8wDsuRUyW+UzA58XoyWt7DQJ1NgGk7DK5P9GQBGoQqotBfJ4G/DvxGrCjVuj
N/Cy2o0gb/e/Aufpm6G9U7RsjSu1LZxEWO+1t5W58t0Iu1kIdWHK8SGT4wDHL/dD
poNLrcE1pK4l2wR2v7sN7Cvik63lwaGIs73RWQSfhMlKbAwxdU3+q6rBqvWSSLzo
WBFo2gJeK4ReTzoigYJTLnYl1gxXmDKhYHmF8LbAQYSOMitxD7qc8gHjdWu+/8+c
KSfrkVQVSjPUBfF7F6mRVMpuoL+Af34uqEVAMf51L31/O3PSvimM4uNYerNxw/6P
SUk5GzgvzhKHR+F6RI/s+Z9kTCabBgidrlmlBTO4HFsQf6uBWxjD5w3sIh5knBxz
25PdeT9hJsSMDCg4O4gq9VnihdveZAMqQBRELHrhruiBhEAPjTUUKnxSXHr4Sg3d
nbkUVGXkqzOtwia/26e4+k9df/0nWw5hNxS9UgPQuFseTiC1zjqsEotbeYnD8INl
JQ7LpIMwG9FU5PQmdOFdJWIHHq24UeuMi+uzTZzh99rQpPzbLAum5y1HuCCUnz2w
bqP4alW/lso8E8aZk5cqSf+rsHUhJKO301tGk9oDxZ6RnX3EpYxnK3PvqpXWMmo4
tqEeMEjW+07X9ltU9P+lnKXdLr77XGF1FreUA7fuIUOcUnA1WVjOJwwgZFtmDuIX
1orNxTOuBA9SI7es+pq3GlbWk/mBjCdvOdxMPa6m4Yq6ZW28gDusujeWxlcKDR/m
cWLbJQAiAWnyLT0uUY5J5IRHLgJD6o9aRc0tmviuwnAVP1vIYh6forqXkOostZFR
SyE7iKyxnCQxYcoMaJUeeVOHwLfEorGuFKxZrzDDGUouMQjWLwxBG6yW7PR0j8dp
hQDnwDMQcLlrxYJhjsIvb/bEM/7aY8eNGfpNf2tuSxpeNEnK+OJFJMIXDfXRSbjp
h309N3i4MKhNXIst9grv1lBijlocdvGAVAwS89M5n4bHNJcDM/XyEMD6ibpRtVsF
PVBBYJY28clpraGqJM78xQIXl2d/OnOQpk5pnoLHknBLUmk3MztqQTKVOz9WUT0b
YM0Y0yE5iSFCnEgsZRTynXX13LB+1i9HePhecCLZXCAIwhDZDkp/W984N4fkK+Wk
TeeitVeLnflA/o5aSofowSJSiTK76a35CI5xv0OUN/jmMWXZHymvwt97DJQfbN/M
4TNRaiaIuQE+RogKb0/Ma28Fgt3Vg1WblFIDadr03xYgRo4ch8Ohfe7brmGunS5I
HbWz2OJKwNfUGZvTpwixTxCp270Mzy9WMiD1/Alyka9UxekH2eOkdAP6wfNKCeHw
xDqcTNFnR/DAEKo8hR8yrkX5SvD30kSyUObaPbIwXTqzsvReXj0xNkMsTjsmLlFK
33y65jNyzobVeXutDEQgu7yHJkFMpoNaMsyVQSMVWdlBq3GC011ZxRCc94XAG+qO
2EvoUg7DlRoz7H4UMps2KXPLADJ12X7ewvV1rC/+5kAEk0Y9CsUcZgQEMJS4hF6d
6UUUU1XVk1yPWgNW/NqIFY+r3+g8bDXNgQWiJ90DDdP3ba5kRrNivluUE+JIijee
UMompYnbpUkIFQ0B5ZFq3HRCCoScL/OGbQWkiOVnBsk+/XaSonOhqusbno1JGV3M
cgqWitY7IDAnO4uOFSLfVuAn7xJZ+h1XR3NHFt/T+jZGpPgGbma9LVv5DiAXH2at
+mbH9E2FaSWiFaTR8MvCzhHsCGo/xQ3yeQByq1gzAWiILockZSU9W07K/0ml2qdJ
0X5gZZgdtQsZVmYJPTZfT/Zadba9b9H3IE52vQjXkZFXIYeUkJZ+mJLOoL+7JX99
uQXAy1fQ4QwzRX+3yI38hrWN4coWaIjQHrWdjcnNVCHI/N7NycnwzqiG6812taEF
KyoMv905bAS3LxlkBRz5vA96RdYYCi8DX8Iu6dlrhBHkOTWmioDFcb6wz2HNBp7d
9nZp9PcA2EHkJGUe4FW75AOaL3HSG9taEY1W7ogRYgUNQth5uyjEvVKxDskZxSdN
x/y9wbzGInpuwLEvavI3+rrjsKy6mZzLhbilSnOLpN4WJcMcDj5ZTh5eb9qpExdW
1tkNZJgXzQfWXKc100ZuU/PSfYmAlAU/d1qWsiZ6pHJqd/+YHILx8vG48bsMAv2Q
4bZ4AlipD1K4/enTdcD4/PkzprkUOug98pNkk9Burzb+dgwAGGGz73q0Shp3Cdg/
NHC/nlnjnLnMn+809JGyYvc/S3i914A8SWJ8ah6x4+jdnnX6ijel2wZauXrQ9Unp
22pa14/2ghlA2t99Yj3wRvnIZ+jazBMA+dFmpMDBNLtQHrtfh5o5tFVnCQrTgeBa
ItWKNlxT8K02jqPhx5iqNwA9YmgvVgJhhf0PiaQtRmo8UuS7NnjcqYPN6yQlIzfh
TFrQqaAag6leIShJs4dXhmy9CkYYV+fVPfW3+EkNPo/RStwYGUMokvLf/ezp9N3R
dRiVvnld85uWSlLvXOFPyydPlDJbX/an2MO3lUzViMTTYjr+6NZXxqh0071PO0+H
QfLzHdXHjDYhmZvOCtLhTfmFbDUvOmQj5ntlzDXBV+aPuPoOB8PZfZvRduqEUAee
SKQ6D152RzivtORCom6gAIeykRNcamC9ED+9/G1RPUncJm9JyKGtSYYMF8sE91W9
mJwWZ/J4iA+tI2yhtP12wCGaWIBzUUpUFm7/pEj6lrhb4ciyoukzcV7Fhd6ve1xw
9DJ/XcIxVjYV4tacjxehM7+9HxM3lZvouR1Vlhr6j7m0VcB7VfKil5ew01XjGCMP
d+l8/OFuf+du0Z05upec643RQBxxr7PyfNf3lo+r+RgpiNMocXOdQvSryvdi4hoE
aWMw3MYY6C3Xr6NHoPYKepAozVxQ4TTOrAYWmA7P708AXekRRBCwTQT5f6BHvCtT
GplvtaYL0dWFvD50mbyvk8fR6eTyXtnwjEUq774mCzE92/VpL3Bh6XDdFQqyBxR4
7q/MF0GCbcZgwjRud1Q8YaqCS0SLfQVdoo5IB+uORDZN6C09PWrXrLUdZ6FYf7tW
m2RtS3xLWyVOtkSlCt0qarhJlHdsd67FzemXZKCjTGPPLVI3pzP3J7hzH5nPET3S
thE7R55h8SG73A1JYYy/NTH+Nm4fU3fWo3IoWFWhbSMYxZXx5+pMd4IPNCvYKZvw
OnOdqHNnycbVXXDuPZxkiOLLVCRiHA3djHFjyPUEALV11ldodJ4ls1XjjoN7ST89
ZKh7FF5mQ+Du74KdF0rNV5EvH9/D/pcfsVxBfw+h/K+vIjBrLuHsrrK6odyZPAX8
SbMzK1fwZcS4Q7aqd+ozu+ag6iy1QPSPpA2ky6/IwFdMvGp9kvPCZQ2/KdTX8mt/
TIABEk/NhIgPuUHj0I9L4PhsnejsJN18FGLd3NuQP77CCf4usjUd4EYOXd00WFKL
fM5DJwEYscjjG8Q0/0qtA6txU6GVnBYKui6Ng6+8+Fi2HcBmRjg3SGG4wxI9L92K
TrrrB1vD6LT5OZV7mnHbF0nwI7n1xOxNpD4Ph2o0Jd6HFwWtCCUFlBC9K5+OpCC3
6mcnoqHMVG/4aKGIv25WmyqH8g9x1McciAJRDdmqsl0wUFxNzTbkH9usEgkHqwR/
67SqJlozIzA07GQfsEUQMc85zhUmabxUGj95tGNj0mBfpjljC7DzYzZY7Goad7Rf
M6QL22gOcrg5gAE3N1Q8gSzcMy+Tt0r4VdzlkqRppeXtQwhpYGVCMykEToxDoJhs
nJmdRJoQLvZI/zKToAtLIOngTB7f6GY7dmD/+Ic2sO4u1r9HUPBQAvwIdcip5UUa
76KSTx6eD0FxfWqVWYTNajXc6yycPaljeKoEI5XWc6+SoDOyyYhSeHDw+uA3FUcR
veqh3Vn2WYFjx3MFswdx90jl/L5mFTTpPedC13FX1CqbjhL8HSNRsx9vMeUwrgb/
LZUXZdPh0OlnJ0OlHKZOWIe32MsUBaihMFRaBN1ZnBWUZbSucF6DBf1rYYjdLjrY
DpoGJ8svFQR4edOkig5dZTgrzXAY44b4EH4O+xkwFgWGoeHZg+1qjHE9rATLv63v
0MoH9EEiHmUfFdm9gp37Sq7apB7CQMxRIXgFJy1OLmUA2XyDX39wFDXDoIowkw7y
RtcB8pN7HMyejs2cazQaA+d9qoGCGQxtmkTaK3mId9TrAlG/cnHMI0yDaxz27o6q
zn+b0WnMSduldmM5z/oXjVdZBXJSw7EQx9+j9K4P4eUXPCYtNuYhKvmIZi80lCNn
L6BDeth8KyDN/LIBm3wqUL++qXlcMtWGHKJKRc5C8K7EC1dttpPipKMEw9tJ7XJN
llB75i7MD7LZgbYJahsBRz6LNdGJEMd1yPmYxiJdtNA9NiAVt/vqfY3no+Nd+Tsz
dp5s9PxDlicp4EiBW0PLNHcessVeKxf6FIGSXvg9cv+UKlj7nk22zgOFLWEHNhnm
gIh+m6A0Y8M4eb448zt+ib69bk4+ntmwHbm/NUtvZ7xWcrIzk3nlHh1sy/CJX6BU
tVtQHS+gWGHBL5aR5EEssulYQE0dShIZVNzEFZL2pf1aGNZpSAS0/cjVdR/UaAK1
kYK2xu2/XbKDmKJXcJ7slnIopwriAqTb6cPwbFW9aUpNYpFwtUpv5DtoK3skwt8a
ZzfiypRq0NUqpiaFyUbmqAkG1eox9cQMbTjrzn0VxawVd6fFmoI2LJV4uGRcxGFB
GzHr53HkfWRy0lz4YfyKuB5o4jd9ujREmeUC/lfskm2ghvbqx3C/iND4QVsYgzBP
FVLLyE1su1j3uBgktrChWoeN4vWUBPHhO3SRC+6qRQKJvWOe+lPZpri9Z6gOzC3B
e3lKSnfQwiDbc7qzoE7hTOiI62HgQUwQpuENsdZc7Uk+BDSyS0lG8A4SsuHrwZT5
92J3RJMfpdTI4VRWsXwyNpnWNyXXkLd81XOd5zkgRmskNkW7yW17vGjL2STUHbut
0osWyeh6mS8vfBXYEzARrL6pc/9tn5LYA9sQODrZDYmLL/omKY3OBNySTcvHOE6Y
sjPAPjTr6q3KwNglgRECrfl/WZtAQozw65G/y+HNZZrSZIsrPgogpEE+eS9WXXbl
QZWLD8+NX78dJk7IPRSpiYYr5ttEycg5YT8p1ww04YpL5swB8Qe5OF2uIibSVOad
r3gkEN7qNPa3yrBw534SSp4IxP5B0oisZPIVrGyfaoG7qukowxnqP9FnBPrva5RT
tiUdx4eqxHzObqizJIaokIvmHkX06oOMQTfN3+XWxnabta3ysb1a8IZRlgb1owNa
G8BiqqBYZLGQBa+OdteNiA1fUis2Q0hYwCJoxBYkJEXCePk4xiPvvX090+flw7+d
sEGq1sswvCZNr1lK4CHqigcPMFUwpu0sGy7cYoudjqzIpcxlKbuz1rcUUIr7wzpF
oMJ1eqaKmZCFNo5Ym86hQQ6rYi2TEY1vzqxrz1/ua6XPMmdsqfJOXdRVtd1rSk+2
4uPdK7MYJvmi2Y+agswWXwGP0SSktUAotSZD5rbzSyuHkkQlHQbxMI7RmeXXCoFe
iCVvwCObL/Sx4zi4AXjPW7edFKXQqOg/jSG7KtM2ALLOcAEhbkn9ugsObUFAmqvS
C34X7glDxDGxJLVyoMGLD4h87sLfy2oyxy5GyolJ9ofJiSjPIdp9cGeJatdvQzJ9
WhDW0+Qk6P3GY+nesGl+AD+nKljVqRHIG6LQNRUy9eBI0YIZc+upUdjRj+W8f/2V
jSwIpnWqUw8bYDb6gtIS0gT7ZS8bO5gBLRB+Y5szZbLl5IjD+FnN7vYMBcdbsmmG
INFAzfYEFu8EjzdK7iBUo7jNEBQhcpObU+71u0Y+tcJj1fGCq3Gg8GI5z/zIvBDc
lypgDhkcABCcHPOy2PmTLyoen75lEZx+iYRpN72yUdjbi3OuJNskvvMmle8jgCyX
fJ/n+3sTQwnTizqW8BV+A7wMxN1A5S1YU8JLcRbdONVyzU0VB0ATtcnQ/OLLl4Zv
r3NXIOW+ylfs9htN8lWdsQWnT7OTMJ7UBDQtgT0YLzTMfuv9Lp+1UWvtCEiCcz0d
N456CucJILcITw+BFLIzNymnjOq7ONb5xUA/J2LBWwC1m35/s/ecLzQbxFrvL8a+
HJsap0+yuYWLDtjlVwflFumQA2ajxNQp9M6bTlJCANjhnCDcalFZQW5upA4Ih4WN
hppWLWb007Xh2d1cTT/ASHHVV68CdTfh7vc69sgxIbYczGRv0N1qZAEBl8gOpcRs
iBq7EslKHAeTS94Ad41bpFaHiTb6PxO5k89wmyOveT1SxWSTLYsrD8URmFQocTVt
I+Az9o64m/VcbPwfwZSkDTkG369bgEi2ZhWnere3VNUbj3nHDTsFoVF6W7tH+zpY
CxEIczJR9H5Z2vmywwRvqxBiss2R5hwfnKnXG5+iat9QOeLCiYDiwmdl6bUPws3L
IRkC757147tj5gjsK7zfHSKS+z75t7/OxK4TFRmXHWPDuQoj8VZBW2LRY1mwiffl
Qed/yBxwEG/+5t2NSpHoVKRHredfmVshwb4G8P6acfKjSgRIgAf8AIYykkxxyw5Q
AvMepEsHJHORSvNEOw8u7JkX/FzRaSZzEapfRsYctzxL6vkN+0aU/QxQjkP0u2RK
GUD30q4o6ieRNeXYdono/CsF/qR9L866P+RlKussOJhLI0+4GUHQHUzkrn+UCB2C
uqNrQF5NM/q6E+GenM8i1MxHBWoH1jR7BFnaqard0hETThWLbzfx0pfJZrfewt1o
gS6DKyAN34Qr4BVW9AHYtLiByP9hsEEMUb4UbETjDHxwCf8pA5IUiFYPvfDkqEOx
SDQiCZ16u+gGqZ238y01jI8GcrQwTvifAyrFmcsG2Gbvy+VOKK5xJu6kXx61/NcA
u9KdPfQrq0ekdmfCEl07XDrzw+ru+Sxk6pZwQ7xAAGM72/KyNs3fZpBk3DXLyagg
e3sKx/9cOJ6P1bnfsQp/fGxmg9/A4v7YuBp2EdVnY/NNARBzRJ/rQD+NMhB8YQ2w
8b2YNOv8WitfajYGxxfkOjMHPViHLT88zbBCkPpOrIHLw/TN+NBB6/8OgqHXqPwt
nHBfPbnyApEwPSAOAD9XFz47/8iWu3cD9TIK6wIWqnrPImnLIBEZezOBQRvdg5Ls
ljnVZ91TKNEY5QINWt2+5WYD0c6cNk1/TCzF2OqXarBezU25bTQV2u7ggnSsEy1N
zgduopMhHLc3k8e81IONqONGkDKVgZ5LjmwqnRoF64BPJfTsCyUlXqxpZhYQ3J5M
tQQL6BHM9Dz5LoDCdR8MtJBvVPeVkctrAfaAgRp4OON45m+a7OLRo12IxlkCFRVH
3m8KL0YTgXQvrYRxfFkLqOw0bJb0XQuqlARSIXYwVpYVWXlTHBXrLyrq21NTkfjQ
PzpXT5zZWOkVmKQBSjnkNPa/wHssRnyWWmuiVOUwYM9XpcD3k8vNgWLaQdpciZVI
1q2TZaTPffkv2PhqPad83vdKeFVZfq5GfexR6Dco1SQyvOIoOuYGNxCTgiG6L1d7
4N++NJGLtHK+WDFPDqmzIF4mFBmAZ/3OPgFZ376B74dn+UIVKKs41gBmXa7tM3hE
WJJSsYI4CE+L5d07r11AlDLqQNRtRZZy/5d/SQdlCMBTgdCeYX1B2jlRI7w0MbVc
Z2qdy2GYGKUInclB8PjUljkPBa0UjYZRO+CptkQax0cbnurAOfr6yCb0tISjGeFk
kNx6Qbg2EvSh0DTPczHKncuJsvsapgvh5oaf0WiKwfXUcxcdM30jYmehjKlDvUrI
vQ3WymeDyoUBdWSnFK7gvm5oGh21Kd79wSaKhMqMuab73ayaLRVGW4kvxsIQmddG
mEfXHFKMxM12atun0xjL0tT1s5zsGoY2ufQgoCUx5uwGoB9zsGNBMW6JOAmuyOEv
dONY0gb0xQGXFa/7l8xlCVkH4hveQCUpF+e3wKXdC9NvRH5EfYjf88Gcsiqc53na
ucgn6xgPQp+3uXm3z6+CGmiBaSwjtsEB2WeZ42E274Vyrpeu9HmTX/YRiekclHZ6
ohRxaNESy22sfqCrplHzfM5AR/gSyzKtuE8twsFLS4PzvePn4PNMEmVZICueB8ad
3TiRsCZLfVkOylxrr59OAaf5ONRzwrDDfBZwGrpDvalw/SKDnqvs9cPHu6o5x9D6
clJixVeUoaX++v1dQluLaML7X0RvwIoSM/BcSPtbOB9+O2LVsZl9rTVDvJuarfTp
n45W54Rg0Jr+213pVc0bAh6QfdG70KrZSu6RPeSiDVGe4wQ01wJBIBxWBBT8LM0z
oRqXjsis8MEObegAaeu2dmNnul6i7gzXuGE6vgigr7Gd5jTA8RhTCn4PLMwfw/dF
f+X/Y09Ok0lwh1qlaXpJe9+u/WifTHqpv7GhxJzHVytQBUiPS7+R4y9WgYaqoTBg
LOtwlBFMBfbmtGHwHrZmiAImgxLYlNN0aDJPbA1pDp6jQMEwtCO0KReBkEUSTH2Q
pd0btsq7++5ugogFdQP2Gh3x6LY4CqQUcUbqNs1G4jpJdhIUei9TykoHh0Ap28ml
W542f3FYOWKEvCePlpUDynZh1bc96Cky2puPwRD2gXUfx6rP2wgBibrHWaCJYwIi
QhBuS9UqtoDkNUIh+svsb9CymDDanNc0zOLKOYntGlyUYL+rrA9rcYBlOUcD+ara
skOk+h+7eQGojQzw4cI4P4AFO1UjdcnnXtX116mJlGRTOEQ4YCLdYT+fwOHssOwo
JoDjBQkEpSOBnGqu97uvo6b2g/JHp7DDLrIwCW/NV2s5jMWOPYBclOT+iC0ENuYP
37r9lasyEtJd7fE7bHVZDr44FkyTRBSIOb1rbmogqcpq2RMJzI2J21ijkAoR5RO9
yodwPMl1Sc91FitHgMptFU7Hcl35Z2Znmfb3GXjmS3XJ1iQnMG7j5PbIPQsq0M/k
KSBiP0dYpda7C9CyPHUKTji7zTTAPcVKotJnZdTuXcR3M9nnyVSm//Y/NeH0W05F
VnyKVQ8pT6c+NEw8J1OM/sxb4PSj953t+N2X/5fxtTKvRhTS30bSj6OzNPUN4spH
0eRIbwAm6as9FOqPMPOK2x3Y+yNHMhrQUHRzGcVWDaXy6kUs/v/blvG+cLb3nR1G
bj9k4AiwwR7ulvX7mmhRfRD6VFfxPZ8WQEq7u/SEqIhB00WXQsf8hdKqjg4OLMgA
/OQs2rm1NEgKP+ufCoCqicWkmajiQRqLTdJsFmDhGokmStyTqqLRDxllqo7HKpHm
v52qot/sOsQbWo1IuQDZA8QUktb80C5VyIKSE/gZzEWQHWwfXZj93ZSSXZQc3ySx
EzxvgcKnryyQMBTSConG6e+N/hHyILf2/fEgIOyqLcUMeoewfbA46iNrkHsiueRp
D/j9GfT8C35eR1AC9eI8wtQs2170r9/9aRfIetDvHHZBETRCIin1cJxnFZPYFnjx
3CyrGyPjcQWfTazWdCziCKcMTEuaha3bwoYBuEcDh6o3Qg6QPQBqyG6wxqAWIa1x
fsydCyMBsmtUiRjkv2D8HzmlIjcsIv25jrY3rVG+EvTFMKwLFINqqkBYMe+rCU4M
Lebb6X+LISVWUloIkKMjCFFJzg9Q5TYKLwDBdtGBxkmoagPTQuO+xO8606NHSM/M
AdWVDg8onwajEIMORISsVjQXndV3PZcw4MxQZUiacyApkmpzVk5BVFF/bORYD7dj
GA56CAhUrKxvXKdBwfU/0bhZWrCqa6WPpRaIy+7HnU1Z2dJ+D+6Y2ZiTEQuXzueI
xsyoI16rQ8n8+e/3q3qy3ONnQAAmAAL5UVDDodiopPhkq0hW708ZETDwnDFmcPHL
yoFDtX3ew+gaSMSWTaS2tA5Ga/Kmdbx+FG0vQbIjQ6hS09y0uQwofu9I4OZkme3k
/FRtl3tIJ8L2pJxTXOtqedToiv59q8yMXNnMSON8ZFLOyS/HdmA8uT/eI/uw0cjp
Wq67w9Pt0q2CJzN5ViWsD+z4nbsfOG8Hk8pttHh+PjxCd3AxOdSZdNSmLlIFDlMy
u/s/51TU04gQ2LEky76C3cU/Nkv3d8P5zGiYGTHwJ7W7Hkm6gPbAoNfvUTVvpwTD
cMXUAqMG874SfuAgUxNURTYMdQ1owP9ATjPP/kDGnIOBHiq+wFs5eOhTzGProXSs
5yHommgPMbseyoeyy63QSWAp68aIacJS7xnsdoNc4nWVy6P3hTiRZmd+w9HOFrRX
woVfup1u7ndgvBGkp1Q0/xqrBkEoTv1B6anCe/m+nMdFFJJV5w+qPqK75s4q0yTF
x0WtwX1eFpe/akpYv9m7e0/WqgknCcFMe5DL02rcQSz0x292Y8TLUc0e05YbVEA+
`protect END_PROTECTED
