`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CL0EJpVguuEqeQUq3PE/l9Vqx6pY2vJ0Q+X8jJUItVvFbWb4GbPRvwbiMNQ3I4pg
w/eFs+pGdsswyQEtzNYm1F1RxUaZ9/EHoenp5dV00Bj4CWELll9LcJ7Ic9oaIhkn
Uk25OMibzXyYhL4z+x0ll/ql/8QW5NxQ3X6xQsUPqWHcFHDl04WKiqzTBiQtQwuJ
cjg+U30/PPdcjwD3NuKj0Ysxeoc0E53D2rFyLNVXctFtITC4M0XymqI/mbNDIY91
0qWMiJi9xENRcIxryMxVdixaF2mwKAmBWUUTT0uTjyAgmSvYeLmtRrAIBVV985sK
N4roE0J/jONrJUGM02m2YggjIlcqi9jZeahvWNKO3CBEHDedqn3442Y/X9Acy4OG
xKVtZfHCGy700JnC/nyj407OXphJ0Oz2CAFx9NRyxg+xhVX+Vv37YOwSVZPKLfW0
s6/j6Dlip2JGznFvYcS7RIySrpfakn3R5SmCP0zWQB04PYECyerBvlE7m7yFxPCu
`protect END_PROTECTED
