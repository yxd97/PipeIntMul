`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LipNMloikOAcuDr7HacpijerBDmnIlrwpJ959KhDv+bRlnC9aNpCHf/oiXVYyFAQ
g1xD6asQzuuAEFY+Y18o1Rh544fDc/LQtnr4Luppte2VvrQBZJSB9OcMjsHo+3ia
dFLgLaJf3mOzzmf1BvwFP0JVdyNXTgYksmJAoq/6YDmfn+OeFCDvHzKv6gy1PpGy
kKJy2DeYZrMJ2jzKlWM9KIMjKw+3/XquBEfy/5OMEWILxWwb6HFNTISpl8yzD6ZV
QbG02hKBB8oA3sD2YbXofihJ+WcxalgqIGKpgYA0kajghF3fBHMe2ZXTHzD3bI4h
DftH88sEq3hO4O53HEi26OX+tBv9FIvczl9nZxvcViUGPgr3rXg86sPVgLjDwWiL
zv4pngA8fwDBBrHtN/4D1RfqRYKrp1ahUz/7z6ysMqfcdE2Xr0mnv/iO1kJlOj9s
SI0F5QBbm/KLk7tWlMkH3hm/rxx0xbg6pe14fT1jfdIWPNX9LeGtssYw/s9bVoSs
`protect END_PROTECTED
