`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YuKktwBa1tHgM1syccRltBhHbiE0m/u+yHMDxG1XYWcoPLKjyt2mogHawFqxIsRD
B+Grg+8G2Sd/qfkk/fXw03tyvlckVeiaKEYNCpMxp+UhTD+bU3/5/uYNx4FZp8BI
zezaZmyx1NdTaIqjkBpZz/XC2bq2hIyu0TsefhyhhI+W9qjwlg/BLl0wDIf7sufk
GA3JrkkAvbXklpKUk1FG55BaxKmMw3L1JYn+mvyC7jQPOrkX+XFAAfNdTYyvKA96
ZZbMTzEQSI/GBIay7MaN0WRe9Iww6UUzy79mQxyQIGrB5htdRN4VrbmU7Aif7dlR
Et/g/qvy5+EfwpqAx16v0fzwnkrCoO7feNMfCwt2SDdBybcEyZMFPmjON5yxal5Y
yls63rIzo61NxF5HNmbQPvFlcz4cW6AWSb7eU96DM0t/2166Fc6TlU9l3E0MFcwz
03F5P0VWSlUA7DIuSvF04m0/7UdVb85j1t8kUBL8D2+JQ2Pd7aaRm4mLC0scXFL2
KQ0fIw1mmts2gQZEFAcTXw==
`protect END_PROTECTED
