`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3dOW+iU8AGTSjBSiSGR4maQRSgpEXQhPlFDEc+3NPdy8mRaeZVpcrWZwSMXyfVif
xeXRXUKvcoUa2cLi+dIZS9Mrmw4GrKyPQpbDq+VHxbVSKasIfi0YOnbVht5q3e2I
yyU6KGMZNQTGdz704LAcBiumLuWxmY6tw4oqj7hqGArKHpQIcRcS0EwWz3VyG2gp
v1kmP1vbbzZ4cQoBP7QuqQzEpU3ZfjGeBAByhiuyDG81nCKpApIdN6jaDcHPo7i7
MIMsjUHESZZchBDrlI+BHHpWp9I8sBBB5BiF7ayKXVKiyfPJhl3Syl6Hb66mTA97
iqaDFS936nOKv0pXhe/ZyM6U2krNOWOlbSaBfwRahMfLZBkxH4hjcnUXHRlo7/aL
wSsRYZLfaMHJ9/juidtAFlD9BejcchXriQ4SSnOBtGXDg4N6n/dhyMNOKAUZt9Rj
spyk0j/FwdGrlzdjNpvGYmfahq65oUVW3CKEHwFaUfdnQkb9Pmlhu3riMUxvXvB9
Ui53vl6Ch7yC0g4jMKdRPwPAB1m2+JBFaK4vD43FTXRLNeY/46EZy4s57uJXWDBg
qaz09uTFU0N1+E7irzzvOr8uBpFQ6tW3MT3cLn2RrgyUPSq7FmSHjN7jXfYRYSST
HPNGDkjZXtR2puCFFlOBY+CkfG05k3tdPHzQs/yLxu3l/0DJoUDXBV07fzdqv166
+EMtWmEqEYOOppF2l9oaZLlIJ3ReeA9FMst1kaTmKQVnIkmvthx5Inxe+QRl6XnJ
Bl/4klLO1v3Ggh6rxQoH6X4WkJXkUpBurpDe6xsDbTLzwqHdl/23GPA/mOVJvyPM
nl2O1Gvz8KdgCraKvuFJWvTjiLc0UsUyVPEALVMLYf+7IpnS8mDnAGYF3Sz/lmr6
ZIiliLEa22ijvUaSaNdEI0ogIbLNEnbLPD+XGhZoKPx5tJZgcZa/h+IxIF69/jae
NB3IdPHho94Rpewr4bOI37Rrnjx2MiKjjuSWvDXF6CJwnouu7O57WjUdxfz4AXRL
Zqe1OF5zI9+VM0Fci6JG95W9fhIedoxDRcn9kyrt+HlS7eZDl9NTEGkuwumMUimy
JQh8UUrcAiJN5kfhhAeyetIGwXmxEZwgIvw02aRj/iDITIbJQ/nzYE1lcm2NUirX
njuMZY61I+tSO1Kd6lwEQEZAxgPtG51no2KG25MHJA0k/C9y22q3ym+M0hIFfuy9
+K4KolgDHchYbLNEJKN5j9I4weqsDx3ycWXud+TjOj/Zjz8I5Te48QPH6oaDosU3
FijNY22hwVU5dhqKkqY1PY6+ijI9BLaGp/aXETOEIR5RFAIVE0ARkQKN4zFJnofC
ORK1OOJMZ0GI3D32jEUGkYNl09Hekle/TuTHjtuSD2fPBNp1lIKXtegwCI799V6y
bOTURFB/vO2EYo+mkKCuem1ts6MI4FHL5iSzmxCTuvPSn4XkP5hgr8O/QeVrj1Ls
j9FsuyC8XIrCtJ4/AxRovmxs0oS0DYb/QVBqe+cncCbaQ9e/50L1EHdstdI2nR6K
XTk0hlvMs9PEdSmJ11nAjJjaAxAFjxJrKeBxiEtLBUZXAKRqx4g5DS5iS3PXLItJ
BqoRUbFAl8ZH90Ti7U0tEuSOD1OR1kD1hPd6fRTBIMzyBlrWn8z2ipwKcHLfOC1u
K/XUbX7gK93S0C9TGRYey9gx3OUc9xBwoY7afBHL1+65c/UlsO3U9+jfXtCm7ba/
lGSlAKZwXQVNQrNpRixupMKXB/nXZTmAyDA15uX1oiR2fv5F3WA7Sl1UkfuRcAPC
eQx/fcFJA1cLt/X8fYT3zHW3f41g/HQEY3DcCqd0VFY/hocV5CS2rmcqhnWBxB4a
44ocELDnRL2JwEeA/nN0/9FU4lqDO5Rc8lwKA7CWV50F1UEpnBGhhSW6KNDVhMmr
K8eKvaJJZz9T67G6gK6Xxs1jMF8nVzC0CY7d3X1aOc3sKHNI3AcQQDoshiRGEIwy
cF9qEZAWqRdVClsuDhLR3hsGYEiXLfUITkcG6OBTyFX8GeBKZPhlMDwCALk8AN96
f2+lmzPbitlKDAkpcH5727PtVktJLG3w5QIF3pLwyGUyPOk+xaD/sZBhYYONchad
5ZM9KnxTT536YtrR9hKGyADFE8yrMMnSVgq089hjl7qEUQBhugzYJJjIVO6EY/m7
KgWYzlowaHIHDjKqvMwBF/IGI7DIAXVFhcok8ASdGL/t1PvbBxrZsx+Scis3r8E5
R2rPQPYFj/ZozYt9qxTgGjJ1gBpdEoL6p0c5m9yYWW8FZsIK9W1jlm/9GXoZip+I
Z2b1k1BRsBUU58c3oX9Nac87FYm3RA+wSCCCiYiq0zG71hOioczcruCphjsuyyop
KODgxcjFkIXaETaTfEsbkBgeH8Cr5Ogae+iyqJbfilCefuSllrRgSFqN/V8O9TRv
FfjfmhLui7lD9IzQ5uEXfoZFNjegoDo6mflnJA8yITto7nYDJx7ag1G3p0r7DAAY
4IjpHAG3ZJRZ3T46tusyVt/hI6GOB8q43QOkZQmY3/5frhJjmIkJ2F1uKyXieSWI
EDWUet5jGtWBKLsoADLogjZd4grDV83cn67nunsPUycM6lJz+2PQtwoCw9249Yvh
XmlOikANycqfFYfwT9DtFRPN2GQTgbtRDXo2iDhytI/jRApxB/quNvMHu2cvsAHS
JPihW5PTqFNqH38uv/yG7mhIvtqREUm/CQ1bHBKiEPpwrdNODTQ6t6Rr4HnwUC/H
jvFalWtuZAqZV1Vo2aYASw9Cs31WiC1cnFlG6k3d5n4fur2XWdvo9SJiMjBYy/Fl
JWIT7BLQ9pN7H2vdqIqPiwKwxI9T/ZBKkCQp7EFOeA0awbLEbAyxaCFXhfTZ6TUA
fXOi+cGgj9bHLOGrTmtYL7pVerd9pDsi0nXl40SM4Q656rGhqhhwMJP4VbB2o1fu
A9uTRKVyJg/yj7cqh5O+F8EQs8aysIo7SuMhtJmQGK8d6rhlWUYcHxuhVpF0wwBm
`protect END_PROTECTED
