`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1LQQYBWl6rphWgFGYwDLj5B+pD2LS35KhUanAeuMYQjCUhzW/7xY7DSYba7CbyLK
/rNe2j64/qXbQcdrfrJV1ctpbVjBtaQ1LCVVFuJxf53eq6VkvP4msbE6WuAF13KR
nTRlCJgE7yUkxdjGM7O5TwciS0QpJuDpF5MtZwM+V9yDSyr0DHArWnPnhpFNVpp/
prsZERfWENPJ9Wp1gECUuG+nhvqzxz8o8RjxdutBp+q3nKNSFBR+mqSaShtN3aRC
NepzT7YjNsJyeUoaiS9JJLWfYLcavItRIyZNFFlLN4hg4kj0p12DcDGVr9w2htYn
i6IfTcRddBIuN5iGeRch/4p6ekH4A2sQ7qi7VFm6/yFEMHiKOtgXHVKYYRU5MuNC
leWvPbgCrfUIRschRA3epPmPpz2YS6sEbdoOgpc8+6sikEzjM7+r54QO4/JpQdVk
GLZQjyfhguVrQLLQ2Ru7DABVYtfElOg9kMwE+OFJKW0auhWGBJDI6y3+1rSpbbVR
0PKHpUXBe44DVrBLLqSEzUW5JM33tFVe1a2Bua3ZQ1lXXOcxgmTTx3VBFWhCJ0T+
VKeK7EJxcLqG11aROJm6tAglcL+5hrmz2wFPtDyr00ocZrRShstHrCMq7aHgCH9j
84Svl1m5MhUB8APaImLDgLym/sDMhlJb57oQAiSy1aniom+AksxpECB1cRPm6Atf
FGNyDG0uYFOrEC9CBRbbHILmtTB9sjjRhQC5pkzcbthjZlChVpyb/f9c5fO09cEu
hxgVsRGH1+lm0Ptawf0j9D+2CiKN3qsE4U5aRSCC0vAW+BVjL4PpZbwnztoKIlyB
wcPBeBjePCPbUX5bMmOMetauEoFt1nJzviIDYXw4U9bxrbnVlZcuIvXkqJORF5zx
8FRKgojz+/YFxy7vCWlT7QLMSx5K3eu7oMVJwaPYI02aEIygkU0W/KmxbELTk2Hx
XLamGZSXtcZ/BiFvPPVDFWgQar8e2P8Yn+zUuMpTqdIyIiEXOX/hkF7aKdm0qK/Y
VSH9jnbAHX6oSGq3i1ZVZ4e4YIut6Fj/kvIxpY6898HXQXlmZx6VPtcWGy9JWcHk
BTL66e+DCaKcTODLBX6zS3x3c17hoYWkpBbOO4ZZGu9ddIYZiJnTijwVO0lmkA4Q
cvvN2iQUseqNW2SwxCbcVxxhTV9IJnuCGlx7YjAUNpOYmDHMHj1bhCUfgbW7PMHw
Kt6TXx4sxonrjQY6P5qEc6J9DpWz1PL6KrPmkjwMp0QQE6KeRkzSc5NGVc3VBXlQ
7cggR/7m0w3H0T4c0RuCsdPIRQBHt7hIM/2/Y8otrpWzhuhRXItYP0DZRKQNOMcr
F/vdvvyC4jormbSj+fi8gV26f/HDX5dzWskUBjfkHIzGyg46Dr9ZCEUWaHNTAcgo
CwvBO8MogdKPU2D0XUgfoXQzGdLybBGVE2DPaF94krQDmWhVTLJ0AmgAdcjT7KU+
S1uUwJamzSq+uGG29JlkpGqLNr0kwVb7ZOGJ3PcV2tyQqMYZqK3bp2/hAK98mq5F
rTbPoFJrzN1c03QDYJoMJp0mvdmOPqS4cvvLYdxZzHNavVEOrU4ZfQZ5fTPyJ59T
okDQHsQA/zR/+VcpFfCCALANy4HWUYoAOyphJ8t6JYtgy431AMGUipiaMSj8Ogdm
/U7f7u/686ddu1BpFdtzEvWCqSarTtDXf0uJFOHFxWyqCUAYn0wqiTcWHsscf+hQ
hUDdsmr2vgxw/T2QjYKjK5+xVPRwg0LdT05r7UWp0k9ImNSeRcV4aAqYIAmuwimQ
8XLTmu8nAeHTxyK9vuI700BnQvXjGe2pO7lo2QY2rz29SNsC51X7h3Ai5c8IKXli
FN6LEdtw0UZziuff7A8FZfAQbnApACtwwg4Ak5BXTAgngIEgMHVrdZnGmsJ0VIN/
zqfkK6AOwzxI3ielJkuR7SSxAAVrZLCwwRn/7ts+Wuwv7t4A3kl2YRmu7FPZgIAc
uE48qVkFTPf7zUABODx80fJ9TSAgpGS/9D7NgeWrYyjaK8hwK9uHWWac7f8BVqd9
DabAS2tf0Nr3skaYMSZpRYN5FQaIRhsv8wd0teQgLcylXMDviqWHm1zihYwwz6p6
+MLKgbrmZa8kK9IA2Xd+wek8ynLDgE7DQLj0xmGbDqtkq0KDxoorJG2rriBB/GAe
NSijK26MYd01RiFNGV/1syjqrfd0EwQjfYbnSTOjOqmxrtGUFq53Ej1wg1wt3AX5
PLMlgMLG54ft58VSEdl0uxhjrKXnJ0gbJ7teG6CKIWiuXNWsD7GHyFwCVFvxMgb5
oV/qd1n7qe99u9HeC2vh41eppym67lx9l5LXu0KdmMVI4ps+7pRrv2vnpU1nqJue
0UdZAXrZhJBPEgeYzzAgMkctVeTBu3VftEHLNldMhL8Ze6vZRmNPJuiOnwZ+WZ82
lWfqGOm+c2WLOuf03QbowcrAHI+f8ADQROhz83rzcHeFmrD5vqZlMd6IuVLOD1Sg
f3CkbylS550FpeMFv1ARSAeQQ+9SY4IRmDyxTzHEdcP7QUsNovahV4uyv97wWoWv
99Hx7cyet8ij6bms4mxgqSJpak8LhafAD2ZRc4DsnfK55m9dqe7wKF0Z9PCCArvM
DZoGhUS8IAeWvTtpvjaUsYpyD7+83jnNzyN+LepqnN6CCLrUPmYQe4/i1lviCZ5+
tYo3JTJEEuru4WH85jsiren11zV+Q/2mG94MXn/i74REEsbseb8hJpG/PDbgRiQ7
3pJFsk5kHeRzsfA91EKhGoHeYIFx5fuOXbyhLj92VqLWLvb9Gieq2s0qh9AUK9Ej
SXv6kXl8fv/gjTEzFw+CMal+6c7nmUD5KTqsEhVTfiEv+GagED1UPh9vmvV9BmHN
1BmgEthhJofyOuJKz7uF9NyBXiS8rSop6T7gu+zCgN3YdpQqFwNRmEZb3rxSSOKc
waXemi+8IqxSb/PPEfAKvnnsOC/LefHrYTT3Pc6RwIuEOH08vjKyczeqU2BmkMBx
XdHMM3ezUUSIB/Vra4/jn0jcbIX3pNIoJwfbD1MsIsNkQzhU7sU0xl/qsMbBaXlo
2V6+qPF1HyVC6xFARBrFVWahJUqhf4EKtF2smGMmpRopVtjUpIigwcPxAdsnjzdd
WhRY61hrnzJBn6eaMoY4azkCC/k1iee5Bc8Ctd0Zfmz71FZoc+lCvvh1P+99HWHl
LFs+vwKenmcGbGonx8pg+OyMmF4zFFMOrwk6j1GodC5atp//hMCNWoneBRvXoC0F
GPqKzqhnwdDsvgBZZxOG61w0mhq8RRpxueGnS4ZiRs4vJzARTEAu2R0j9rSs84Cx
07mgFrpH4TtzYHcKN2JLk3tOdN9ghtWnsL0kLugYsGYiVFo7tNf5lPFys8DwvChD
oQsP3oAJIm/iQW0xOmO5yQ3bTlypxHOJQbdHRy/m8SMMzzvcR6fTJMdvUugIEcCV
COGEO2BjKFJSlTeTL4VAsJfKiSMgByPizn1KnBxx5uB4HrY/pkoFdS7EBhNDYoRx
I1WZokqbCWHpjbTkmanrFZDz2GgzIuA0XTROy5CjyoTGKAjcTrsHmmCISQkWyAjA
DDMxNnS51VU4TtZSmSY32MOwLavD7lMZi6i2kwo4/OVUvnF/Y7zvoNjh85UYWy9w
XBu1W5CpYoAYda6Aa2PvE4zgpnMi+l5mUeLFToTZj699dBslMVSkNT3c0z71BPLY
qC6A49/czkOaNC4CpKEa/h9F1LLhnTS/1Kvv820LfGL69pnNehiuJwp3kA5iwGVJ
Z3OwY47tco8Aahhk2gdw8PxEDxkUoC5vfgnvEPfR4+k2oEacHfoaVfaxjSOdOmEl
Zrgyibrj3KJjx9RWLWZFmau0z2ZdhQm3LyzqmVNCbBv8NHKOihKZXxtuJ417CnB9
zUVZETdoRqa/9PN09HnqbnDrwPxvCWzW/2+RsvlY/WKQGFlfW0Fga6x0uxQfUcpa
h7ymNhJOrGxJZt2HqGvLj827ycIVu/P9/0KFYu66CyO0VmNz6avvwiG5W+6IlJFe
cEs66iosZa9li8oDmQHWJbJu5i9c8yHpsVNeSJ0vLETck+wkRDiG+01bfFACwXxx
nlLeXPgNNrzkf66kVqB+31AeeyVunak3/du2Ty/ao1jeHlBfSmaMArFMLgxycNQW
uk4mVyeww4JzHjjSv5rhjs3+EWEpbEWy9CdBI7aTOv8fepULTEXrZWfcAyOWmXjS
ZiMU9L/ISXRPw1Wdy8QuO+cdIAjB6ttoeKgN3TLJYppwXaAIyPQGK+/NDBoO5j4S
ypiBtu/CFECuVuaOBA/lzf0W9BpiKipxxdGLjM7X7zaVqhwgT9yDvEHaZdcsRcz5
n9/qpkoaCPClG6neTkEcdTwCs/xuGn2RH4coxgMxuSo+CAAVY41uPIVD+Yx4qIc6
re/u/abCdC2NVly3l54sU0PrVjIJj060Zig48Ib8iGgttD3WINnOiD/EFS8hk2ja
G7vr28JhTh2X082EcJihLNHrB+1F5sc0lhoWPKfgsRWoNPDu3LuC59xgP8Zvdtdt
IT3U/+qe1YV5tQY1bbSm8lS6OJ/fIWJnFTtrCNmqnmwFQkoxSbSUFZ3NFhagBl+O
/dcqHG26z9P1sgajaafHDVqCUaaVZuorm41A2djSL3BLrDPD8y2XCBUokaf0Lvck
c4Y28128ulT1PDeoakvR80PVfzBbipl4XEgjRV+WeSVxLlJo7mD2DZmtzBbl4rCS
YOKWo/1mSH1Ktyt8EzB7YGlwQKa103Vm7B8H50lOJ6yMekmY05plwLbfnw090TA1
CZj4U6NJbJklN1T3xzg8Elj2Y+2ga6j8Yh+MPCt95NQc18yUmgffa2g7E0eJBw4R
oDniZeWcWMMkVl4/MCYZzb5WyiNE5v4w0uE/gxtqYqAIMyYtjkfFbhJxWYO6+yv6
If1CjGWXyQMLuIq4EbgzvqmPkMk4jcR/mTG8eIKCg85GwMk0gcbUNrU2ES4bwU/A
WdTEPjTDPgspqNC/s36HFycdaH4Gfq8bJh65WqzTpBtSakgfmvMpxICgHW25GfFz
IvRxXFyO9W+WEe9zFWeksKhNmW6hI8bcziGOhoQ0WzfGj2XjU8oKrkeZNOQ+tHSk
W1nOI1q0iGQKIK+mawM/t5FeYTvNmSvkh0SflCC/OCt252QDB9lji1CCHJ3p1RQ9
KOvYdxexYvwTCB0DxL0zGlb6zBwBEhvhcvHtdT7Kd1eP6EF6ROxE3+meHueXsdzL
RxKILLOH8RYHfUfm+GhCEaR5rrYVymAOsvtz47/1dhCB00nYpu01Y94C3Tu6CT17
0vDRF6l0gKHQCSbJQTUx9Dz4jQO8uI7JQpglBD25wjp6/coyKamylt7hRqjA8nvp
tiXhY1l28VYaj7E46s1GV1a544V6qIeJr8m1H/UMOEjWe5ofB/+HMr/uDdgv/YSy
FngGLjxoYgwG1NgIhGFYJX68GskEv6SpFTzZ/x61A06JU4LE/WZ7E2U/ZXFvjWH7
oQ0fvpcfcjelnLJOoNHbdpyrioi8ak9dT+eQhFLdjQgLE5VIRWpXHKF+gFbWyeYJ
e8MgoCKM4l/fBs7ubK0vvxbn++Q6hrsARzGmgqSpGShy9PONaK15elmd3uxe5T+/
txzwqT4Vq5Q603x5pgbNnE3EpXmKuyczpACgjGJ/9OrcQ0YkMy4jI6v21BqlWDvG
k5sZCQ3fe39HQbPILcS3/X6CdKyhz9H2nA9kMG35QpWJSzVaLA8y0P/rRR7jQFY5
nJeLNUgB36SaS0JqQmKYWc5eNsz42NXsTgwuzbG6F66dw9EZ5kjBZiTGE/mYcOrf
yRbZG/cotDg/8B7GFdYTKF6bsXcjSo9+SnWsw7ZCYnVEfta8ZGQEv9EGjGXowdkX
sx/c7FeSawXKRkgSEX3A+RLkK2EsoU8wkFifFofzLXqz7wuB4XPd0MjYeQPGfFjk
ASM5qKubROFCz00umzdlI4W0LsGK0iYNZDt6h6wukXQ+SIRwC1pQyNT1xgQRyYrj
yzrLhltSxAiBTxHs7GZUyIHaRUbOdNxXHN9ardmHeYrD4tPbRDq3q2gcWQYuepPg
gLSb3aYxUDLfFPANPN+GiUqBFvnLKDlWo7nx2K1FVCHeVbJ1WEBqJLPr6sB9WqEu
9hQC0YScePGL/dMfdry+7q50Kl2wBmrVgbXuVXPGI9j/7HVdmHK8sA3lhNRFggaw
8cmDO19cnxdhdLZGdAz93Viat478GpWPBBOhTXBI6Qkd/JeOSxL4wKFEdC2OLPrG
CVyELly9cJGtznckpDvnN5HHBrP4SzNKQPrRJ3idORazbFymUrgtcNLwiEYECg4r
vCsW6HdujFzvgyAOzSXWAQuC313bn2h3ibOSidokjWl21Ex+Bc64KW7BPDo01yd/
Z160ea8pLBINheLuJHGJyeNRCqgWWhNEhLwC3TeByj0SkwRIuwJpFqOqDmWaBuJZ
cQZwnuWoANb36MxMqgaMn6kF/UUl4Em2z7T3Qb3mAh32m4tF5xOid9zGLoTAYVil
0yZJCiIQBgm+IlsuN0P5xFctOFi+47INgDi0du8VZa9wK4Tbpz3hE2MUwYnSAEic
yvIDP9dlAObq0SuksbI+P7/miWHT3bkwe1PNE6wbmtodBcPtQ/092CzHySKqAZUI
Vsj7M2lt/zOOUgUvdYM/wYdvIBVV+4bzrgO/6LNQdM9XlE02phy3vby1Cd3yshHD
JQR6fFOBXsgGdBQkRJeB+ysc/lv3xpbxPkBvnK4D2cKesUCNm3Ou/Os7zFj8qNsa
gr0aDpbzUgQ90CvC2De5oZ2Svn8uDn7pbm4UCdIP0DLF4kk4T9CZDRYvcLcfgSXq
LWdYNPFWHQJ6ZqSyKXX4ZYyRZzIgyrQplahUisSBoom22wN/+FSt4i4ppCAukAJ0
fwZ1rbJfzXFs0jHIibedgPerKYj/t6/ajaq80FL7YKi/lfW3QkCSGs1GAQ478+Bt
+f3tmhHa2cHz3+rybRy/9/4uhAORURlwOVkPfMpNNpesKybWIB/eBf+XjG2hi69m
G3BU6zOVBPB0OddLMqA7i0APC9RLo+LxzRrfqUom0aeGvYg2up9hI1HNM/pjbsGn
1rfZwpfXz0nVL6IYmqXVD5ZsusF518T79QbqpYVzFxyNspvsm+BZA6kPlOnLpYvT
CmnMNcmXS0yrdCugd/DEvvyi8HlcUrPIR/JUNcIUS9xN+yd7INQOUr685EvZYRFT
2amkgcpFwFEBWmzqx8ECMAeP0Or1nSextlj+SJlwT7vej5ohGgOxEAWXD0GrnAi8
FZl2JeH3SzSa9xPKf+0adPQeLo5OX3mRzGh4qQ20qxepdqgKEQ+cEfgHPWZWjjKT
VzuukC7hwCkfhaQnCbeDKtUqH7qeQD0bO2imf5L3iyjINwZQL2wEt1Js9X5jzGvE
ro0hutJ1NZQAxDOZCD8/lSkFyTaSmmfD+nEy+XrNxfzF+5Y+Kswxch5q8db3viWC
K82+8Yh40LlXEi2WYdmwhigpofijNMSTy2VS9eZERQNnkCyNu5a8uFksdkvID8J+
yAUbFQpALR6u9mxbuBTg1RxUQUb/V84guqsnWnq94temcB2p5dxBY3ahQuPVsvGG
j/V17wv5RYaQ/bI2qxKQ+IGhVib4ryEufMB37Ll3kilFIZm1OFJgSCHBk42fYQ3K
2c8s5SRgFmxjzjtqTo+Ne23d7IV6bJTsdGbCHPni7kvigFWg5DbwFaf/3ykZX/zt
NacGbL0L83J1i+x4V4DKFA4Abmnm+cx0+5o65biYq0gH2xGa9G4CWdnwKgQzHumH
XdX+Bv/YgT7S4YWVWx98r7+i/NIyqdHxhAAruOzHDZ3xXBsHkrkB1Mt93YMe7Vou
NoS4UMJQzPKSqP/amSW4+ggQQy2FJpr/jbySW9nVEOTyTpapvgi3z11LkReaEXac
gDtaIwZior9EbocAG+MZl0PBD7IydPzo32sA6GO8/aez2A0rOhXGhok4rhHH/dP2
AzwplvXf2hOTzTOoZypjyqbEDFUaX0Wsjkt/9woYR6Vm72cRjiIahWB1+fhaR+JJ
mVq+SAijD1u1CWKu8rfwM2pdSUd3Sj7txpFigPfKCz5L8nUhlzRQgIXW9BUEFp1H
+djgtT7UlgsLE908HmBjBd5CjQ35VfcJh4OhsCCcgBJ5FZl/w9A1bkrQdMM4gD5A
cvGBahcZQ/FRinB9fa2z2xfqQrjYo0/hbkdv5RtBaDsSDcQoiOY2EIrAuzpp8Cmi
cDAmQeAkCPg8ifxEuBtUypxK23hUZuDPIyTWqqmWTnOnGXmjLbO9u6YBE9YM4y+b
6olh8uYLCBtlPICERqyTjHffRbcDbo+aPYAqWXGzCGKbXoxuc5WnWSnDAjIp+u+j
clolX5Vr6hWBLcz90Eu28SizTeS6gNebf7ujfLg3DgNhE39r+I+kIF21e/O57fBO
wIUg9D8SrOQaHLsEFEhIX17XvilHpWyxBE8KWxkXFvKlh5zGD1lVT7ciRSkc1pr9
dNbsEpQWh/oACeVLW7MP+yVdDfnGus9JfUpHPpMbeiHioQihZBt58ipKHRHiMEZl
j0YwkRJ+5zBTsPWbdpn8NyQb8nNNBuH9lMSnxJaTEfBpY1qBDS6xo2MP4kdvXvsw
iH9/EreVrwGga4YZmAoeiuk5Y4V5px3NOWcpxs8bFebFIpp2BS9Xqvo7QI63hUx1
di8SSP3J1H0DN6kgL3ivfnQ5evTN4ugio+9K1DSYHl6ag3C5PaT4nH+qQMrdThAO
CFxUvVZQZEvU9Dt5W+Zp3QIz71tjB6deuRrcKbILnZJzrvkYb1tWPISQOZ5IeGhT
Gj9JoTFBC2+wOedqdogXC4BrK3UHFm6jXg6MYKHp+yUjrAN6+sVj33vFjohNN8nM
4m/Qc1xGRf4Hp02WXLMV6RVEMsqv+YkkC7h/2H944xF1RiYLHz4MAnFD45eATZsl
ar+0B0UXRhSOQ0ynlfFd58kpsynTYuLjeOI0fKCK+lVlV/9k0oBv37ZMIzyKEDSA
GKqvQUI1zysiQOyD/uLOuU7Ne+KFMw4ZNcgFyTbtioqwKWmVhQWyu0kJ6tgpfNvr
m5+cOxE5Ukr1zFHMD3eZaP6IXeed7xgMiUxgEHSBYMLAGHuhLiZRNlT+NVVGhwmP
feG7ilgh6eHqX5ALP3F5z3pg8OIixJV/g+ZA/0iQcAYxPUG2f5N4q3dUfNLOyVo8
ZN+o49maro+/93t/ImUNPXeD/Xwu2iQa3MrLHOLL6WFcnfpqRzX0fX3nphcVj3zI
P7QaOEd1fbMtoYT+iizH8SWHgaj3KpW9y4ewk316BaXm+l2R22j5Lsh/544TFkzk
tdI+nQNBCYmejOtB17EHYGs9BzOJrhgcInqpcGpY8ATW97bQC2qEd0yRQ7oPOVcv
2hPB4Ycj8uC31zrN6f0spE9hY98yBzdWDWViGWajgTIWcAGCSxWTO3TnoF7dB8hB
eMf2ou7Q51ie5C94pMEVgYkHUusuoF2VE5AgS7Nx5Rn39Abgb0Sn09n+U9EfNsRo
WR/FNh2LOXU4/dBkM4Hjj5A57+iWUIdwZ3+zXCsCDxExdcQ2HeH0ZHw1ztQIKDVy
Zv25TfZOnXNuWugey+jXhbBpGk4HLrm3SFRmR8bXvDVtoZCUk4SLMs/FfTsTFXvR
1J8Gw8g/yA/aNQAlvgIVjsvcPoDzjSpbS4f4/OrvgmhOgNf8sTwrl/GcNlpXiBbJ
e06vdhom7FTLJciHelW0fPccZk21Q8QBGFE6fKclzQIlXqviT5NfxOnbIiKeGOyT
RWklGNvHbP+7aGkKXE6SHywSieMPSI5g44jNmRp2NJJO4016Jx+z2VWl2J2c/Ryd
/aNaGLPhzqVqi4ScVL5V68T2fBdGQ9/uwxp8JpNEpUuu4a7yNkVCnjqIS2mki0lb
f88kMQF9qwLhgbn3lkOw4j8/tGSWgtMJSLEReYYIcWqjMfSIM9s0Y2IvZKlvFgZb
0TlVEg7TAybivW0ZSUl+ybJIzbY0KCRnsX/MV033GtihpkDCL8seS2InQu380SCZ
ePxcr9XTrXOOFlOTarpB93m3gHooRmEx3b7jEn3kXYMib1sWLinYBlqyPlkf5eOl
QhuCp/OGU8c3pevI81kLZsKBsRoe1e/g39A8VkR04/WTpfbb29FWD7LrnQL0Wl7b
jaVXDtxvvE2NhaaNKznruawCJA+F3pW3hd/Sv4e8dHGU490EojOrByW2v+PcX9yX
lhTPI/oxQSDVOTu5oQyjwAMJ0Vi5h0JARrPp8naVITICWIL+kdl7B6YkV9umkXdQ
DbLEYV1ZAP7TtZhmTva+Ga5vvykapc/VPGqv0VnVW6AbCfLo4Dj6ZBzmlFJibwCs
hXLK7Edl3TFWWL+z/m6lSdcfdKT1gzRmFxDjhG97HOu/4BtJavXhxh59NXg/FIXz
TeRDPsWkPDRj8wVZ/9EObL7e+ccO6tcQvPTEnBw1QLl9wfpV5n6Q+zqfbBcaW9no
kx4fH7glK8DSjZpkJFMh+LGIGha4goWIl2kXRs8M4REIzuBdGh2oYYMqDEdv14Fw
BzJvObYlS84FQFdlDYRp/xC2eC6iHZCuwXq48/O88SKF2/xyiubDLaLjj4lqck8P
ugelueq65Nb2T3wl2FNC/z6JhxLeHB4DcUDIjzaTSbohHXssE1JOSR2mzZPDxU5P
M+JM3tMjGWmfX3PG8kVtcGVNMeac+oLn9k5ICu11ydkIT/RVceQ1awuUJUCebhBf
HOtX8JWBWvhM/5hCv6XGTWDkeyLI0qgC8ZT025ksac5FDOAYM/QoXd9dpRtW877/
iS8mZtE1ZMjL6worYmSh5NHRZXFkZyFyumlD0wpVpNhm1PRDDlIwuawaPKFMhm5y
G98HeKGzjiySt32e8mFq+dFRaYZb+/9IzekEdoE0e9B1NImy5cQ+zuuGHnd2rJ6D
dnpurrzVxLEm0xtxM653UlwNJ4KqwWEUw3o06ZlEqtKlR79X9Vfa0nFFMmoKvzhf
2m7SmZ2i/nSBJsr0zAZOCDxwbYkjFTwHeWvZly4C00suKUgba1FyiDxhbGNOKGYJ
MeyxtRLZUpIx67SAcrCXQPRIm8tzYQjRLAHwJsIjG4buzn6GRZxsecKpzPvRBvkM
K+z2tVZ1rPiAUaJOUcheNXjLQPM4wWNt3xMhXjBUzp50dlqBBbhMi0+IJRbblV3g
sz3cBShUQL5r+PBFNBbvg7F8pMnvOJcilYFIT+lB+OpdRTP8kQByjj9/k3QBkzZM
xrhQe+HnencYbLeVqXMEM/0WfNlfy2PLRdHuoHEe3XQ/7XwJxNHKyIrW2YOOvRgW
I0RVN7CsVbziA6YeiWSgSKZKNYcxdYm7VSpHyT6H+qMSq4zZ+KIMH3hoMowNTnSm
KKjqADDqgFTtOwWs1d26cYAUid70Mpa1KbfvZ41mk97C+OD7vtBAXT2l1NlYn2gN
iD3MFSoKuucgrJdybdnvb1bb7YBFUwYPzmO5sbxbBoA099MSU1cPEPp1/1BmHdU0
NxJ8fpNXFAj73H3Sn0MXl4S4KUpeMgmE0AHM0d8srLLPNCejcTKIxP/C7VrpVVqS
C441SeaiSq3E11V2EPCyF7zmLlWC8yMttWUPFMJWZSQ8ZfxJdBmbqv1F+PfWWa3y
1bykmgt/DdlPaCQzyitQOC1lMK83Ap5/DwZAUaf6ojOpN2LT9M1MnprFb7XXtRyp
uUMbs0YnNESYaECzRro0XWFE5P7VJfeBCoOug2lC/qquzpSy73RPp+C4CAUjxJgL
JmAX07bc/CVABN5fVxYI378idXQNINzs/blq8OumkPDwSsYDGLEaeb6dXApHpnFC
uj9IigdkUgwXcu0Er0JcOF+GoNvPt2jC7ErvpEsH9PAMNHIg4aHg0syUGqdDmaXo
O7Nbo/ozY1gNRSa7xv4lNqa2D7NCvipOQdm7CS9zQPdc0mHy5d0u/gk/DtXocayp
Z+h1zBaNZ9LFzmgtEKUVDfWKgC6jBYbus3FldsXn6VklwESKYktagicYWcW/YNJz
tSjkWXu0xzaeBV++KDzJaWJZC6bQdmoQAZAnD+VfYUcdbMcATzKQoKkzaum3gIOY
CV3bPt8oJn8ckOrn9n5TGTiU0tie0kUvZtopzZCZQg2sU1nSTr1QW3wh3EzCJfBn
CpNt21vddXkrk6u1kfXWyMRY+UP+gS5ifjOSyFT7ZAhw8c8meK0/HwFBXeONp+Dp
OTa7APn6ef8NFvrBHoTCA8FPjBJqWZbKZcEC/Yv8bNMaP//Jh41jnl5s5sssS/KR
p+ghZmS8wTJ6e0pGyzcL3iqPn3lWXBq8tMX7ns7AKTfJsIZQGLZD1m9UiWhiLiPp
P6p/xTYPhtluoemrker8ivbXGJbOdMCgNcaBcKivkMSbm/RzfGemWXgJABrLtpKX
OyaTzfFnOWqWlWSl5xHegYDpAzhUTr9j+AhQyk0NYu49ogX0NtgXb6LSUmsyYy8P
waeDKxuxun4E/jyCk4dPGZxGROwE3hBfwOFnyOXH3ImrgdZKYl7gLh/hGO8/iile
HiDeVmhcDqZkg7jJhPmxJ/4mc/agZt9YYsY0DRGI14pDdgcyUAhBbNlsInmQT64v
rx9wjJXHp2bz1bu6tpcoo4R6WpM2HjQew5j412vTUOOLfvyBcj0IWsI/L8LQoiy6
V0GFWNa9L7YpZMiiH0xr2cQVT2giBjlyAwTHXW2i8ces1UVMFTU1hUQBVGlcALX1
SWh6rTqZkLqhn/2xXqQuFTCT4siNQOqA1kL/IlyLKGe7Q7Q5DlQMF6cxTEhTsaqf
/z6mX/LFCqwxPZgYwRtp7nStlCtQSWyxLSAa6dahC2WnQjyDKiOXu40fjkeqAmsJ
s2W82hlOV0lLNtinqjkhS/dmXIF/MQMsSvvw6aGSjwKkl0xtX1t2M7WvyOZ0/U4t
JC+tMQOkd+BPTDpIAp/E1mE5Yqwh5jJOb5FyUrw4t5VPSNKE1SEH5DVduFyXnsmu
esaxnIvuXWaC7F/u1pqVsOyGyaXzcdxIdL+Ue8vwxhzIo/IksLdJaJHtf8SB/T23
PQVa9qgmTp22UO4tjCVcsBWqv+5YTmCSOLC+SY5jRl2sW8rO0JN7h8WJbxKb6BdL
tEGcEGRhR0y6qk2Rn4LzrM/bLMpyygZRb6Rwp0VuNwAINE/S8ZCNeZgRfQVnjtaf
+sElF5YqcAcNkG1cCdtycYIIzuar1QOQEt043tTlFnZW5n2P2UxaEwVrLNUJGLLa
NDdPJaCNVTyLXUhVgh3vnCLQzOrhkcNlVhHlj/BQIq126qWF2nt/mGsEuTMOdpx5
PSaYvMTIdUJVJBeJ4hkF/8BngsuIi2OE3sWen+iwjqEsZAuEt4OPi5WdjVxuDRo3
MH5PU7QtBuMGfal5OprnzGg5rrhSk00qboCOs+aERw/iDTDHquEhi5P6dqcWdf1n
O4m3pAwpe0TcqvXHP3ZmRpSCGuO94w5yJ60+UGq/t3WeCupk0Vbtq9iA5HLsvgkG
HdnbZJOtBaadYZhhVHUZZxL2Jomat3+dwCJmyyus4z3ik4z4vsVUBFKO45SCV/2o
/LdY03/hMVj4bmKk0ZKhlTTD2tCsli2+QPdGbRYOwEQXg8ungRFuPEypUiCBb9En
yVbRFMvk/VE5K1744UycJlEd8RV6iYJXd4XWPZ8LY3QB9r4RZHr6gQGezJPXEcbQ
MUhDOe1wJ/NDuqPksNbYUavBR0MUW9noOWvQB2wrdfQB8UHkgQphli8sCC+UcfGF
3EOnlu7LbX0dzaBFmhKaDTPGA5CBwkLyhTllU/cW9iPVqGZ+5c+SQ5Yd8NeU0FHL
YVse9jDctRN0c2MOo5vHSgJBERbevZe8Vx/XV2uKaXHo+swHaOLjrFSNZOi9AhKd
kFPQpxUTNr3Ft9u2HSqD+w9MYAmIZ45GDVME7tUd/lge/NDALZZvw44V2kpqs59m
xsBHHwOJs/joSUsrQ5X1dTyTr4whx6y2kRopJ0MDziDu9mzpL7ref5V5UAbntVz/
243vzN6WYAnj4CUmUf4O5UcaLaJtAnbj1q5YBAA4kBAchuJb+x7U1u5CwU/Qm1oL
eE2MagrwFbvHSi/u9POWcysTPd0G7+Q4p9U7uqW3KuPZ9cX/8SlOyEiY4ggnzcHa
1CZ3GPzB3AYBjPkMqv9QQr+9NxdYFHHA6JX0nsF2RfhQ8A+jgYPZ4kpjlWmVtmt7
uJEQSKnwCOGSwIsGf6RkbdGzyt2iPmyGi+rrnQ2NdNv1xLX/BnFhc5SviDPDpj9k
ECUWh1NO4sOym2OZywUysJymO47KRY9s32QhZhS2iSCY8Z0jaJ5WTWbRm4UHNhyf
2K7px3tuYEjpnkexkqCD7DXFSOVU+5MKvxEvPvAiwYs6cHoPb7wJ9BzwZzSOu87S
FfaWQjP/3KaD2lsIR7bJ9CFoEkauf+Lm0bK9fYwGbNZbDSxSlwwyDZ/b3defjNSm
zI5FiUXXRqHCUM48TAA+QlIGViUp5K2RS2YVWRPnlvGAZun673TF3XK2Bo8W+t/I
Dd+/mhJLMIY3LfHKVgAfW9qutmP2rcxCvHizzUkV1YeCTcBktZWXnPxWvZvNtkOa
U0mAboJfec3ElemBZykXF7yaWHKuamJVVeeZy7b8WSx5QnSxycfwIlaK8ASolKIg
O9tHxxqY1wbQ6WTu3u5wM7HNcELASfm00TEx/H5b0WW6u7DpT4ZQ4xe0vPiqi2tC
cjnOP6x0F29zw96mn54aGxtZv0h+0NHchRtIG06eG4OCkZWX4wPUzQuyPj7IijSW
zKASiArUqyBYepqRxVqobpw+TSxTvxFVMAwGXaZCGMHJT9ZszCUPKn6yR6TeYVO/
V4Ag5K8xrhC2bvZEnslXenMUu7IHJF6kYWsQYTte+CspVx99ffp3vUKeS5Z26ZIp
RyFfzVTapfS5eoP6t2ldkNgvP9S99vrZpTL7Cj+XQLKNxBfydEp/AFjZ8WNK3cRx
ALZyxNqvNPwhk/OsluoJ2U3tox34BI58abTI1PmStk0Pw0sXymFZY6imlgFrpCPb
zrcexIqCkDJlkLxjcoG3c1yCxDytA537shzeoCaucmip/HYZXhLgcgDlM8RuAhpm
LVLt4SG2GF3E/xviykYCmnwzSLGU2jNBokBoxIJOYsM6LlbBjKeope5cDDQhe3rz
OKEjAZryBUYeVBbyIeDQAt50LW1Z6Ohpm0EiuzTjlTBvi3S5gLHGUNd/liqANlUr
jXkW3igS7YKI9xIX2RxfXUPSIkeex9KZ/7kX/fNEiW/fIgQv/XUisr8BopwKZB5a
cA4jF2GxAE8zbEojRULxFeLTb3lM0A6iqui0+fhiqhZgN/14rp+OTYb8+0arJeTE
IDFFxBZI5uPxG6Zn1myboXd2yibrGa67l9PE2vUw3gshnYDiUU84PQbCk/T/7M+g
oVSrlO4hvmt0lElEJcw7mofXWnx6coiG9FAlLQow3tzrVJr9PxzUaOCF/oHpngqv
ZLEynUT7NslTlEBHlwCxXDsyDgEfTpgcTpnokFML7oV0TPBzKK6M8tC7rzqFsVx/
OEVoCUH1ks+hdCEjib4UAiRpzNj9T6Pse+gbuNyvVCJ8CNE56Rcd+isY+Hm0rOul
TAO0q3wudY4/wj/UVUjtvxmOxCCSuafvBNOJ/OGrnsfeMiX81wrUJts/qzfJFpCq
hqKtTwOZ5UKKC3M5nDkOUtHFcJibufAKyOSx3nQ2s3suk8GtACGUjEnLWdiOxeEL
CITSpPqmTp+qqEDm4n/Pb05ZHTY1gujAvS1KnWbqabqwN6CiQ1I3/AZziWffLWcb
CMB7ya7KEP02JiONaK32MtAdQ4HsFbYN6IW5ANQOF2TD5RB2c/DqnL+33wtIKq75
7fpIGEo2pH420PGzLpR66amCl2zuelrMwfneikI5Lkp5CXWFBEBp38g2lnVodzEB
HlWsY85OJbiB8HWMNHXgRaOk1XO8gdf3H/GkVS0FzAMsEUWst6YU4Qt8GEz8+l3T
BHHIRcHP9l2HcGJcUvDdIvjk+l3A+IWqxLJmUKlyVrD+cwuot1sVK+OzN2Ubh6Zj
Mnedn/z0qxXx+CmO0e3ReGp0i6u3CRlv/wFXcGYhLqxZ8LK3pbyb9zI7sv0iFNET
PEr9U1DbKKhv4dP6UzNDUeK0KCvU+EHrKL/gkbIQxPPier4smL0we0cCF1rZgrN1
J9wIaXsUvu+kVZYLb9B4QgGXKNsksJK1NZHPPx57/zFr4t6b91s6pBY2ftGrQliC
1aHbAEUuzRxfKV77pFLu/PXJwk+GogeNfr7PvZ+ZCY1ajQGI8WlVDL33BRYZDIAs
ePgBkcb+L3v7zaBTYrJDFKxV3ROmBD9Ws5AgLOEBNxS/xvmdG8PxvdN0Gy+xoiJc
VRFBdxs9vJjFKrd/dY+HSXYVRC4nn3HN8/jsV9V58TpeYFSqfAaMmZHx5OzmxMPa
6zbW1tmmQTa9DIh4YAi/4URzyxxdm05l8qGvOgXzR8HgvEDFUa6cspFus2HC1qkl
HY2/5WwVhyoPuo75nQgsXFlPGU7QeAUCLEnvGwSn3skr+I3y4viqzuQAzJpBohnQ
O8iNZj77qkIHkH6Xor0UkC1lcM82kPZok2X9+7LsV+rX3YOovBUjNlsuZYPBBlhV
IgsY9SHTlkIvNgUp2Yb36GSOfRWPkQQYPjcCEFEN/JR8r3Fry7W4FwjQHRhA4iL+
h7AsVNHpe9WEtMhSTbRn0OsTUX6frBqpBUxsYTK6yi3bOqfrK/k/4KdFjuIMytbI
AptX3U1Zo8htv3Q11ptS/TegzH5Td5iP1fKo6FftLwCjpkpLOyoFNTnBKfJu1Tc7
D4lockCHJqfPQ6f7dYnYyrAkb0G/XiN2H9FQ5CzvJ82U9WRF2pmCgXMsz2MpkL60
kmXE/DHCVSTOkt8/HXxTTUBI11CYe8XhxKBdSkw3eHy92wjZGq4vD1+dSBZUtZ6h
UjpGF4GwHvUWJEtofT9m/mBxjMhaZTZ9lc+KMW+9yZP8skzBbNsLGJPIAMyTF1PK
8JFfQbh/ekQ9wWJZWPP+Vz3VbZESFiG6IXd2z+Jc/yZGo3DM+VdUUNXvg2LOzlTL
0CuHjbVbUY2Y1tY+2/Z8xXUE53FWzlUXTOELeiSzEk9MAG2BB8Dmt5IUE1NBI3go
DF3ZIePMmQjnNdEUE7siFhyztBobkqsQ6V2r6P0GBB9rZe7DxiU9QD254f8c4olP
h+jJgx/p6UYMg9y4CsejmaQo4hya0nSY3pXDbGPl4K7CQQRfjfq41RmXIl3RPd1S
g1I3ZoDvV5tByaIHXhZLGTdtkGOIdS0N8S6kFk8gCfPn9zNR5QkEixxeLYXRIKzX
WrRkCf042eobb4zsDpidad44VtvRx5tDZR7qZw/uBk/u6rlf0+4AXSTZ67/iZBWi
OXVzaL+z+ntuNQwfWjKGiYg7x05ndmneBckwh8oQm5IGwjQSOqs2uGHNs6GakapL
yad4OfjOIT3IgIQu4s6GR7fVb9um/fXbG/FuSp1yKIopqpHbjhdJn913BCYQ65ZG
yLiKvVtMs0bHZJKneKcOwl5DxzXouXRkACDnqCKQbDoBF+Vwk5/Sif0BLe12Dip0
FVsAbvZSS0s4ENOHwfs86YyuBG3FpQ4Ty0ERk44gOYpumjPrfKKwI6kTklHIVGNt
FgOAytGIpV2oKabcIqEgw3X+IpTUaJ9W4jXnTbHcMPVAco5jQQgoJz7OjaGJyklC
EXOMz9L5cOCsF3IQN/UbGlR7wMUo7Ge8GiaCqyjKaxEh5S5F/7ZBW/q/69W9j3rA
Hn+y4N47qztXf9+Gsq1neZNe9YwZxFUm+FtHRw8vcXctTrtk19n9Zi1I2zrgPBZm
XXQ84+leAeO6ZygxBgj9boOjom+vDbJm/5NaBi/ChRN2OBLVMftQ3+BVonAne8YR
IMUQlYL3fM7hn78SdGZyWK90/4nfQH/GS+BaZePp/rCGZyTNQF7aTn0alps3v0GM
mcdTEs49RW4bxnahi+25X2i6ke/88le48OTdAoPKJjOWuHnw2szn6+AQbUDBE0JD
1w39Ee7EDKp/Zoc31r/nfYD1x6t79DOlhautAiBpGKdG3vqnPa6u1ljCHQEd4bSI
9rziDZkd+A+iqxY6r43/RCF0saVcV4QEK4BcZh7O9VIrm7FrwDFrHJYgFRinMa9B
WNMbdA0GugG0GNBXwOmWWOHRFDMHswwuFsNe+KtuykVdZ0Pj6wYXGbNmIyy2yyKs
WkMVF+gzYkUmd6wR9bpdxYNF+162FnJuF0Xn5p9SNJJHUxhdBdRXtFsEdzg64UKL
xueYIlVsnmZckUqJyvig24eQvFsaV7XyavknccZREuYKnuylbNePQpEkIz78JIh+
yVtXbzYWH4+zi9npeIorihbzGiSQUZUV4ySRGOq5mJgxyQ4bRGLtYh5x0wcK1Lfc
WG9D3sVaM3nDuoL+z/gmfhLBlPhvpuszKJbYLjntQZrQZ059fBOa/GslKOLnS8Cc
szbayMt4bPi5MGRRSA8NDyEc8G/PzX0PEBV69ORsD01UyYWn2HuIUb5ea2FbrvMo
KLrj8kngVRvhwEgiq9fRn2GX7e9yD5zWX9HoNTK4/yKmvLYZCSxVVtCYHdRIUByg
ac+OiOswGOAcAfu/gLIRnAjqMzuuQ/SO9jfUec7tCZxmWtPOC9j42emFNvHwP0jI
+5VD5BJz97QjWBpQMUeNW6E2wJ/bUjlSe5KKLKx57y6lVgg18ZDvrVbZRCQ8KKJR
2Qg4gx/vO1hLtcN56IqBYZ2z+2lPrMU2YCs627Ojuk1jp4ikv2wIaOY0kyHTqzmV
iVrnUs7a4oPPQyFMqpX6SDglQEJIw81Va4U8OvLjTPqE2SEA0tz8QsF9qMORFbRl
/87BDU4Al80xAGEs7c/rZLYZ1s7FwWfhBX5xoCFjN+zvK63yWQSxniXQZgMuv9sx
Qwe0AvgHay7rEBb3PFCOWBbcuKhZnjuDLKgk9ml2gFtMe/w5mRQzFVdQiwiVZ268
6g+wCYL7A5siCXkV2VrhJzPtEBrq5HL1Lgroi7DTWMIIItN4cKnnoAlgFnJvnuC+
7ZXok/0SoXBA+HsLkSBT7U3diWC3C+agIymFAAvJVTcYoX2ZrqzHeoKkatF8k+ZX
siplS8Ep0xrgG0BQlsJln/Jt2msRxGVRI9IrDuQR0gphB/3xKUVLgCeurKEoTzuv
JtJ+nGU1l3RoEDL0U1PWaQz5uWJLLc0HyRIh7KHl3vlbsZyb7/CpD94QjJ4skbNs
v9Ftgck40ebwy8hfBG3O84f1baG6S4u2tuQ0ms4kLbYIv29Dhi4xveO3f5zBj2lZ
j/vrit5sQTOXfo2Pf5cdRcsXElNCOSyloA/0/2IkX1R3YFAugXXTT1gdTvoC2H9E
VTypwloBu28JINrrgrHhgyehvidSWH82nbASaZNSwhtQUjdLbG4ZTK30FWkyr/PV
KTdByZMY9QiAS5vrKovS6jfcY/Tld6Pj1V/HJhJTQLZ+8TYZXONkSejuHQLj/BDN
IaqFzuUb+5RDqP8f9zf8z1w2suQ+lgcgm6xEdpcCdrAgkjtmgcjX9h0m1jEaZdLO
FomxrxHqXZsg25moqSQolIiR215hJpH2PRJatD6PNAWkXlBp5VBDZJsujuHVA9xD
GzL+rNUXWPShAbnnlXbVfQ8Yosf1o0hDNRSm7jwIE40vJ9PpwLkiE7TjkxKkV/O8
i45+zT7/Wg5H61aAgS4oXnqbR9YacUbNG4D/NTciue5nmQXX7HRTOSWSfuRxEVGH
dBysMQ1/Pqm9kBgNRd/M3GfVL+dM5c9oWqshjxRX1x/i3pVkuWqFejLTjyse2ZBe
z6sTORd0hKEkzGu7b7nmWUG/XKRdwxW9Id92ntoodRchu3RV7TViePWHkna2MwLU
X5x+/4+lQYyuKRGsxc/Nzc819l6yneRLF8mQHYxX6f5s7xmXN2PIyBZK6FSdA6Ko
Xry6fTZ88uZmUMmdAnHsp2b8zShCmfWxhZq40nRL9DtRrsG09JvkAeq8Wzjtxrji
A5CExgEx+K8lv6ocYM70C2L+ydG5blTxWdi/vxhaxbpV8l5K3wLrB4sPVBQsQG8F
JJT7UHF+lGWwEu7n0VDcupjDmQZ0WlLAjuZrlzXP7Xpc2DzjQbVL3980l+rMnq4C
RIQaSiO5S8Hcb6TXa6Tjhp2Qvm9z92iAlwbnTnA0qVlOH03qAG8IQNnFyjmfUQ/8
jAFADLoejuXbffVoLyrUctjC5NI0jvsrlYMl2r0Q0U0XkKM0rrk8fy9ehX5LFxY8
4sUk3SUoW3d5PH3aO8sBzKpfD02S/4ENvuguz3Q1XmWxwFcuMbbfNkSjeRpB+Lg9
Lm5tOf/sDHs0OFqh7lq+d7XaxZUu5uuV3If2WKFHfJMFWZYBoKq6w0zRWpjXh6Vr
AUr+y7BMmnqgmkc2FvCAeJkb5b5mL7A5IEBnBrS3cduU1VpueSlO6VvH4vgvZLS7
abL7vw0DkfzRebHtW/k99ECGRBDXzdVRAvHwnuXlfrUiIMhYreEQL/GHfko8TZI/
ZMKhu7VYqIyskeAhNxUc/USjPsOHaJ7fF4oXWVLRPIkUhSVmSjHZTLrJfxyjkRAh
UIQ2J8257X9Vc4gSb118oxE2aTTe2PNz+1cOkifAIhZHBhD/9sdbrjxxqpcVFqYj
xq/1BXG+HTwIxYPC7PKmUlZSQuEWaKIJK2pHySEoZkBvuQOVVWLzpl27HMZIJpFo
46RT84RY+5jPFnjJNb4SOcEsNBwGH1I7WZsE+sVULA018XJJCcAOTnU31PXh6qXl
yuY3YHWJxJ/rXGbSdFHNScXSxfrOS18edCuM9OHzRAVBlk3P/36aKViP0OOIwwwP
Bx9xZC22Z/2Yf/rclSEwROm/Qkpmd9S+uJZ7n0oMdAflNG067P0nsQEXR4I3lCyS
G5iTNDF0YVNuDGqy1Mv9VLKX1mVvam2uOSBHGOblVtBYs3auLIONzO34bsbLrmj3
3D1CGwbxUTKGI6L/INDc34fxPWB8Q/0PFMRk+XnHNQ19GRfxS6lS7qYHp/KHFe0A
suZHJaKqufoZqdWRh5cDMqb5tP3sowUPR2BsqE42xDh5MSiAXdKVD0hxegnlKLL3
5ip7VjwANIjpCIyGfMO5E2O83dZxr1tX/au4FXAuXpi/3Po7C91pyPOXVCjTsrkr
B99oZLZE4wUBihE0/al+Dwk2eQJQspgYltG8bWO+jPob5nV0debC4+UXBCxrElwq
KWGv6wGAuBCLkVeEuWvd1VWmfB2f9rYPaeHaAfSQu6DjybPqphG7iQbmG0JDt2tE
3RU1rTg0wXS9SJtPZKx+zRvCOjetH9oSkqV7eUUWAoF2Cyn3zJts3jRm0eAOb/hG
SpzUa4yMIzaGO5fmxOs1NUo9f0EH04tQNCrysZabIUCQih9/jvjv9EAx/Gpa3itl
FmKI9S7kL4La8UHNTyVJGAzhOSC8T2N9egt1OpH+T4T1PTpBEejSVzHZ8pL8W5qy
cwlfhho8aYHaWcDDLg9vVPAEK4v1DC9M5CF+pPEa7j9IQJvAqJqOlDP3JiX8eQfE
3ofOtIrAIWPQHGTsarLp8yEHsexCieKjCWqqqf+5tPS9LegMBOmckPOnXkoRSs97
F7nyII4iOa/ezITjI5tU1+JcqZkdNo7a0NXqvgfJT0izF0+OKjqXrmQSGiGPSRRQ
w9hZfdWvg7rCu2TIBMTGV+ghavQ18aF1d7Hd1eFJoJhYmhM35smIM19slFxywQJ0
LovGfB/kzQIGiy4FJE2EpKNbdJnp3ldyTWP9ZKjwc2TZl7HMCrpG2JKWQIDnf13u
XBUEiaoj6sfRxMvdoblAFr8lEj7aijVyczE8BkXHYWUuu+qALxT5v1mDJSodAwR1
4mMSRAZbZjn4QJGt2Ja9xrCGXe6/CqgqhmKa2k9O+/yRf4d1nZhQtvZMKjDMSsjK
DtECgQ2B08gxwGhA5WW1M7qhvhyFTTkJaTD0bRTw5jcQ5ZxlDZyzDMPt8WYcPhio
qwMUIO13gq4cT4hdfI28ugx3rObuSl4Xv3tNexf2kIS8Sse4jN3bc4XbfAc0wkIj
7lTL78wzJFXjifALUTiQOC9laD2gAxxsX2ShSN3clVuXhWuxREwMHNJR2qX/950B
P6o3PChjkKriRnfpWkVoEgD8FnvCr0v/RSatIw+tqEJPh38c5yz8uDGjr+i1710X
1cCOPQrpkoejMo2JXl9ihcwDnxJg6wx4tUBdsQzrpPh6U0H8pXwE/bRoTXk7lCCh
qtavudrtv9zNUpC0LknEncCY1dMhMn+wk4dmG6Q5z38L5gTZ0eFSLELFJez6lIvJ
YkC5tCeqFjhKl9+o2kHxGRO9LPBuXsl/74LC5cPh5dIe1kSFo0uWxRjcXwp4doq/
qNHXtJBR+NQ+j5ojpNx2GeK8QjDgHxWL6Z1eoZqV2tCHqcd6CEUE+QY33L8TPeQ5
/2cO2L632+zzxPkLV9KWW4gN2mMJRzgxiIHnrlPztSde/j8697qM5B6xhCHf2YzG
DhqTsjkPb7Bhvo/NkyUl+egij7U1zsbPCV21Y5VPmPCoor93UgDjPyS5Qap5lXE9
2z8SAcVYWz5M5+gMv/xf+IwKt+/lIAkVBfTuilpOhSGb3W24kyvTieSus1S++H1R
CMBdMwQvSB1wmVtNsQcpKFNSwZ93l7sogiu7xMxr4z8m40fuwncVBgIFw50fluyd
Zc/g9YuHddFzsEScsbXFb2/CXS9rOmjgqpLeQhqf1fi3Pu7YoIlo0z1g09tBS9yq
6tc1A0uj+CqjeFlPD5UjZNqipmceTTJfQ5Vjcx3tqcIs62VHrz2s12y+6sz7/kyr
/eYZcIhnqg6SgruXFKF7RXnk3v5yYlyAMlsF8C+PbExekgCTcap5kYGoPqfLMA2U
f7eS05yProLc/ahqsiqof4EI1IDUOchZOVVOEW++MuXOxdXfmph5y1s31xPSCF5F
mu7C6uL/NmYfH1USYPSbs2ppMKUZVrYoRUTy+mhNHnLk9FCeNhnDIfU5lVKnJU3G
R62YLjWOCRvNVpXezsYB0HreRlyxC371J83rOadrhzOLjRAnwYTfzu1FtzZX0Oj+
M7FUWB5NneqZEOlKKMAZng+aRcNe9fj2uSKiiqHSSCKr1EqIUBZ8ne9eqrS+Pj3A
zknERnW1P/Ee1QpaRAST1weJOhk700WrhxMnS1QCUsW77Lu+HFIwaPeCtZe7PfAJ
HgmzHB9mDD8wUFH1ooWTzBbkZBkR9ZKax5TVpz7LsFeZ0lVUIx2zUZDE9mc1aVEe
JzqGr3yMVwR005IcGLfzG5cuC/ot56DaQGtf1OysByWzFNt2EVh4mrG8uBLBFAJU
+WROOxVw2g46OOHNsyyP9wW61iR7I671a9gF6xyu3GauXgJO0GqNHa0ERJ/7AygG
caa1eirqAwRw4WIPcJyuSL3gQqkL3GN7oiBmHjhfQ3tnGqsE2BkYG8GEGZfS5GXb
QlW7dMJVuyVE5BRfveqhPnIKMrQCgXn1z1DdikhksWmeunerITdOmPBelQ9o3CFp
GvIhLJDXAnvWIfPnm9jb7M2y/RKINRqnPq99D195gkQi2JMOmzr57AwVxMJNwCrc
r9KXB2q+uV9adVcY8JfuTs00gzTjXdoJAxIvakvrmWuDD5IgjSfCfSs7NAcvZdaN
HqYK6x/LCO3xlv9LArUMo43SUyVDDH7PAKpm/ucjYNxXbE80nKLuYN5THXqdme4k
Xss3mwEACv6m0DehIt10PVzXFNLIa4bgF68oFV7BllR3FsBplNGkXdO5ZT64mMPh
JgOQcs+q687LUT4MwnLxegd4/4sa5TK7inbLhj83Zg+hBWo6eS0+rPUp9GtxavrF
YX9SeXgjw/9/AGvDYnAlKtq08XvUAvASR1GMt6sAifPZARFPwH05TUc+90XyXpX6
vTmioWwXYEEvUJ9cwBKuTCpjY3+Imvpk4Im/oePwLjrygbwVjBPR9oWNnwbRiNNs
w9ewWBrj2lI3T3auMqKblqn8bG6wwG7xNqthIaTX0EjVOTXnmzkP/SidcMdHfhWA
dtGoFQX7uBBFvPWZ+bT3KdBGmaB2fm4CGZdnDyNGYJ6Mz4dAr+sQk5nzhlg0slZx
42YrtLRr5lN0twJwNjins/h3DxkDiPzghJ7fEuj2YKGiXG+LyjDJAhvj0pNj0too
bPkRL94yv0XgJa8QBq0gYQkqe2r9lXIZUPUES0rVWVe4/yglwdTCIwijNyEDaeRF
gwczTeR5hDItXWSSrMAMzph7CrL2LVk5iCYb3eVNdqtdAAIPfP4z0coyauTci42D
p6CTLScHPkVhzp7EQl1T2B0d7Cm4gEGTDSRkmSRh5TswoGNNhVRPt0xQ7PAJyxI/
pmyo0KfbkoHnrLyX6J2HYfsUrBa2oBQfcYkhbMRcLZla6YBqrs4XJN5Qav8mlbcK
1PEiNSk7nIQFDpQG8GDUPz+dQKqO/abiQHdHNrtJxObBkOSFtGp7J+UMxX/bwoga
9N6XA0/aKqbSHAVlZdiD+3NMvuaaV+U4ShqqSnketivFECJMZrS2DHAGEK1X01V5
YFDabZfr6iFT0Z6S4/wNJk7nZD3SoLmRZJnwlXzqdCaNR3cSRIE3Vrtmjc5C/gJA
k1snIgHdgMQ2SQOm/mvJIXbt2E+zdPNzfcIBbLy/XlRXz1pQpFGyNQbmaMUxLe8m
/c4+IcPMOCyh3+mYzOAfaw0UnyRrmikCHuVtKHtXMeWoxEptk/sEZwDO0aTp+Y7c
kgsHG9kST/oHxAtfWB9dCSFIkl/uz+NI4Oap1oG7G5diye+PP5X/YRFNzG3M6EIp
0C8Eh+1fzSryWsbxgHIMj9Ub9Vqg7QXYZhr/Pj7rG470yqaYYXMpnlHhlq/wS/V7
+Jj6ytBOStri100R0fGvpF/f2Y8UBdme5XcU3z06Xii0iC5aTHZaODU2PZ/MR7mO
njK8ztHx14uE7m4+fHHenehXlg1Ye/B5+NpP28/p+mcr9B1dEyXhCPr56GnyA/3M
ORgl4jFOL7svrd96rfrE1Kx/XJXj7nFjM9PHn+Lt8Uyv2IILey4J60/c8XflcVvR
8FZRXOqfMQWMm2XzR7Gsk2cZnCFW0naaXfhGsNI5+vrzVID+i5PDAMJBhuZUbhmw
DML+jXXVr+0A59NddROuQp01mglsXr9Y5kfKXmr7itzjIm5GPzXAYTMKhB+cJS1k
q2GouQSycXRy1Ke7TVJQ5bBoDYKsx+Qh+jp/KnqDCQRdCXPBv4R6h5wvgFPIxRLc
D91f1MQ0mtPV29IRiJMTQ3zIRiYNV2KfpeF5acqfrRzoyLQ98DCLZM8r1rXweaF5
91SFPbYydG6Uh6r9HpC2b5DkDN/NrNO9ri2Hwj8UMDTdzGyYOIG+gDfZa9bW0KGs
Qcq/gWQPCAzMYrzJ8DXJVyXQy4u7qkbA7iWDq+i0fMLQ8nKlKI/uzjkbJky6DXx+
8TZiwwONPS0dmWam0eiHjrwQ8D2mCT/iOnyraXcgnA7Ze6sx2rJ/10rngDMS8ame
w6Mk05YM4gTXBxExxwcwu7zQeEFF4HeXXlkHxnsLmnIeK3N/9ZkEhCO35LhyiloU
Ks1HdCrVybaIlCMY+Ca02PHu7OiG/6B+up/2S8C95xGXaLGw8UeRc13kufnaZw48
AJLiH8yBeXGLN0VrE8MzBOVny1KRgeNjktzqTbGXxpuFHiWpYE+r+iCt8UxWG4D6
9FeZLYzYbbwHDxy34Of8/S9z2m8fwudzqAJm48mfjuNTPnBY8PymkpRX/aeNoqFN
4q8It7NrIGzjj3un+SU0+c7LXp5ggFfb8Q6+spuvppLG66X8OZ4/JTw4cf3+5hyK
MeZL7vuJpCinS0z62NVRCBZOZsbfay/k/nCi/BJxTdkxBJc2n7UYN1c5oaAtVHw9
4y6rykCIml2aAr9c5pXh7+abPNOwEBENfWBBfdecAx9WoAaj1ppJyeT+z4/Rh/Hd
vYIUQQBZ08t9E98GBBOGUNQxmS9viE5f/Qsf/15v5OoAUenAHikRIMWMQ+MUVlEA
GvMrRtP0QtBcy1bWWpJHeS042lbfPe+rYClgbXtjEui8/6JY5EhtNC08uezAQxFJ
aFIkPbRTtE5gBWmI8HalETy3yXyA2Ymwb+Ri9gJqdgue8DlzZgwpLvqFhkT7uGIu
uhh2j35gkFaThZiVHVlv9aYabilQY/RuuiVspEOpOWT/5Pr0fsNGhKJxzy0ejtiP
S+nyTieAYUJ3OSF22q3txXFcYFuxtZ9jii/5q0Kaf5+8nnaqXhECm2i3Wuuhe8nk
kZ1QhClLtbV2WJAZ9dNYNGhXQi+nDKhD+zK5LeyN1y/HWL1Ax6ZoXiJSq9aYqpgD
1SRpPTe/fI981sZqerAoBEof8SRen6EoIkQcvkAfcK4Nn03yEYuvHML5bjSBDyNt
NIoEP8Qffs0unlkDdiYxDGkwflCqSF3HD1AIJRGwFinaIxVx/l+Lgm9F4dDAP1yH
sz8KsRw5lSOVF3SdxNkV5DTfXV4x+oEXhQIIzbknxPw8Doi2aIx+y7zvs3HHBffr
Xis2uxE2oI3ojBbDoM4tc2h7amqiLr+Fxo/KzKxKCSz3ee92tyiZMfOPDQeqR8NO
djg6kuwAXon3V7/RiCKZfbAKoCUKvBaK0W8bwfzSAL0PW+V+6RtbmzLHeC0LMSQG
2LDHydmH47dxktPoE1PcNwBsEOxFmfnpMMN7P4mg/d7TCL4qo0UuDPyP6nHn9SGv
qkW5ScOSeZkz367AnaTG5xU0u67gijndjVt2y4/dwrL35hopLa/jlHKMJQPIK0u5
S9vMabOUHnYB1sPa0bf+0f3w8FOxpuHVU3Gv2zwCfe+BifHVctSmSzp6ESnNGoKL
pem8iNYgji7XRq4U0MFmoP9+Il4GBIj/TALW+ITW/zgWI4FgoNpflIx1VQiZ+o0z
iro0DPJzn7eSW0GW6w0MjvunGAc4VwguONfIHQtnOsN3I/BScjMgdf4Q9IhCNTt8
DBERpP6B0GpQgsQIHOdWO29ramT4FdvlJAhDzLSKVDewIrXA3xOS8qYhgFyGu+Ek
er9P3D1aP4zax0MJCRuUyFwLolGDTNESyl/+RsXIczo3ys7Py2dCUE57XdYi3J9c
d5JRRw9HXUPAqfb5nGfjPy7zKJpm5roePIWk/ztUBHAtzHdErj4l+LTgBC3aVlAo
aovmtyknBl0ghI3bryuevMgc3mEOA1nUz2n7mK39w1soIH6axp/RFR0Bk9Ph9Ab2
F5vAwKwa+86mBWVW8g6VNB/C7fa8KEQHqHRb0t0LZmN8hn6EjS9k/JBEG2SpPIw0
W+FROuxGkQn94HOVB8yy4w60vbrtJpt1494AuZuz6ZOOFQW3KBkIhLtn5te6Vmgm
MIUrWpWP26YoCB2W018nzl86nIjFFGH4tyNCvCe7Y5Hiuk1lR+jFNYwRnxsH5P07
oJoQ46dACpgfYb/RU/UPwrv4DsWFLOzgz39vbwYE+HKpd5Vx92ClGSBt9hUxLngr
pMaZHssTbB44i0pas0vLqWkBfhf+niOwzYBa6ptUu9eGwDF+MYQH9zUhN7dkKfIA
6M/EZLZlIxxJd7u86jCoyMgRRqcO42HIf1rCHWHfaQSJEEXsoUF0Okh55TspJNPe
3pPs9xVye7IIp4bUcLjg/mMEZK0HhWTOEdb68+FdP532VcY8srU9jLn+YXsgTZi9
r7h3DlI8DWu0LzHxnGAvsZQQMd1KX8l848r2PotlC1T7pExVtR7LtLf0ntdGJebg
RsJd2t8/Y/VhmppFAKJWtFXJcA5fytvUU4kt2IqXT2oTt2PdKJOJ75ltozIhMD0q
001jQgC8YPH+CIxhUuejIkqM1TrUl/SNwn/dDNnzL0gURi0AX1I8pQOrbaX0KVnf
hngjhC8boW95fQx4b7v9Yti7A3rOfpTyZPj1+W9V6/E++02j/uPTmLeAn/kT7PnN
4WFi81JWgvrQq7Q6ENEC5ur+Anr3O0P+55o74vtYp7mFCpfEtIQn3EqC/z/lOcy+
JRbhgQPonvGfuC4K0RimwnYdwFKtzNMW4cg8/2QR6XAV1L/H7zSqknPnLHkJxzsr
ce+aQq/EUiMG4u0vl7NYry++swURuchOxjrb3nQcx7/drkyGOVRN4+k5hVCwqGG4
hy7Cu10rJ0uWT0d97aXLVf6tUTkV0xO6CnY5TUZqJJSUwtTMEm/yQ34jZwphKWhz
BeX/g34MN3Khkv0lYF/FxJYFOHgeY64aODy/fgAdyhQzBYQyovT6StwZpEPJyupQ
2LEYkd+FDgqpX3cM7nNqiztsd7tiupgb3kd0UrbQNZ4r3yPr1RgguMOJ8wKNxNN3
CicqRcj89PuNgzTVoLCo6IeBJt9+hwnnFeofS2OxQA/JbRWSu4XcF5d2OqiTOush
70jeiRrgYrVCnbI9XusqiyafM+ApMgeI1w1UMbNb1IyqZbrl1pB4tFxE6/DXS/Vy
nMpZ3hhmWdyrCq77BE//IPIyNBYoSQthLyO2m+nAZSXg7kvY84q6VFvMYZoA+ETt
8810grYQoEVyStBgTMmYsqAeSl0pZXk/iQoiJzuBmLkOu2t0kygGRiUzK2PC+1bd
XGe3BFB7X3kebdwGWeyBAV5icmsTR6/bGN3qYagIYwe0XR/FYO2X6Cn3ORn0occI
kC2BGfye8bg9FgAvUdMfPTMUfR1K2PhYXdDPNfaxnaeKryPmxNzhiGQ0+ieKYtk3
w4BFHeR0/HFjG0e5AY+TtooMpDzW+7E8gBLcX3GQk6cC7AHrWOjMyTxB3YhIRZfn
e5hlHBcT8egFnYrC6593mUHhZM+Eh3Cdb9ni7he1/gJaEmy8aV/tOAwtbIGOCdWJ
pkwT/fY/ZJ3PK4Y5LmzkRgtLa6GuioaTFm4hFMKk42RHTQVa0K/kxF8TNgtNIqd6
MvcvNVeTSVAf3vGB8Ep2qJe6Y8YZd7tJu1Do0vBUFK4szroHLejSZnPUXrB56746
TIyAMDgmP+uD59kEAHORxT+GEr/+6bOjpKjkXzAHuIOO397nDXTO8lxBhtgxdHW4
olbJDosu47HzmoYwTETDriJYtfPaHDhRFUyeol7CArX6lJUdYmZCrJ6QNiFNxaqV
1Z6N6qYRF7MC/bMxIA6YJ8VaOCTobAu5XS2c9/cn2bXeWr8q5W2/WDTaSoiTD717
HvBnMBVWlKqsd3QWSdUz4/8S1FFS8zEC5c2KtsKVsni8wjYfgII/0Xdwj+aPW0vk
kr9uZ1rEp2txasWJnqbIcV5m2HOPf9ITUq/PXhqWhONEtTf7YboYOPCXnwc300/S
z+69oVSidGso60Pa+9N6CGo+CURUowRoHJZYQGaNmsnz/jEsLHWAtEcCfBVJATLB
K6uhOx1ijuYuOL5kArEes2eRdt+p9kbouGA06qKQYYMppCJ++u9FTAVLdQdMaWfq
mcK3qGipDkzii0Q4dhPFCkDwzzvBMRxXAw09+mzFhJ2xUDe1mlhqVgCPtpFTPuab
dOOiSA9nuLSTREpqp1eOUIsUfy5xquyedrFxTdG7J2kqn80x/QEbt4qEJoPhdb8o
rKHfhJ/5n5n4k9mtj/OhiTPMfajk+KDCImAHr8EKMlbpWGdvT0es4FKr4wEDNzNh
E/p16stkpucepMLJ689LdRCeUrWW15bLAGaGvkApByMsv164PSyml7RrZHuZ+WA0
06D72HeY5uRZzW/LrfbJ1U8yhr/1E5BYUoiTGrk89Bhy/sI1Y74twFAP8rBizi/D
cmQ2kjuKxjiOhUbNS9I36oW7oqJPEBSyPEYI9CNCexzyCB21dir/lqd97WQXeohM
N3/Vp69v1dXC9lYiVRb2TCSxYVgbygXOVf3ThuPfoPfVPM3XlKq49Zjwpo+uY3pW
5dIgYL62Vo11v11zKkh/RXPQC+9k9hlZwEyGyDuYQEJPNwEPm97Q5ft6XrTYDqh9
0cOtJH95VrTlCfpNOmlG0WLpU+B9MkkgahSaL9bmbaJSTEtyNs3tREwsZnD8DkEz
gNUhfUcLZ/9DXuVXC33eA2d7TE03ittFglqgmTe6WCiYD1zXmFVx7QrfEIHEs92w
STK6trpERu2gMheNdX5iLGd7oznLpDxKHhsokUWZoiOvt1qt0gqHp4Ytb7jm05gX
0vd1xG5nPf+ho8YOJtiKYzDCWXqivDVUh+uUbaXoedlSIy7PB/ZhGqpfzeWcoRFy
zRZIhhTdP742bE6L8iTiBjYAwTp342d/EJ5O5lfsxTa5R/hjaOu/jKWA9i/U+ckB
CJfsYd30ClVay3JQKsvolMD2KmeiBKGMswCKbjBYYC9cHK/A+LuFRNC1XqZ3PR22
RPp5t3Iv+PyP81yw+PRyVb+EuU50eyUcAfNN01w0PU8FJbZGANHQaqIDWid5NL/z
C1u++/z4H7Adg5ew/bdgQ8fx6rUk6tAaLE9oWK95nRe/RwfZ9mmOK3IjvcCI//Rl
00gVDrAX1xcEwyTd+K+5BqAQ/Lcwol2e4lpNUsMLdAWPupF5klN/EPA7eLhegqgX
HOOfvkOaQ0NJfoLHyIcCTqJ0Ipz4rD5NFexl5aJopqQbxB1AnhmEDcPWvaL0GkQb
r452jrV7swYUVPsP65YSUgC/mCYafYeEntQlWPgc7L1+D0+qAmxMMwqaS9tI6HjD
xI8fLq71bkDPGMxltv/3pYAoNJk5trO9/w1fvv8HkUx4sgfbpyVjW4ZDKckZZM8A
dePNaeCMJcThxgFdRxsMQGepBwG+NgkHzaQBGrzmjO8xrByiyQ3YB1Drdb08gqIU
ZX5lN3KwsZttCaU+tPN1GsYAF8gOWQpn4tVs1yBo9ID53sMxe8sfnPYlZTzlh7CH
BS6nM+rMMdcob3nUj7K4I6nEI95iiQbCQzNPpJ1/O/oIlCCB5Rw6FHLi/mjO7ysn
BVZqaKwFgIYTeQ3JNSUwUJVRG/LYAW8GO89Ym5FrWkt6uX7vuBFwKwGAzllNDwa6
oktliO8G/CSCyfaEuFXyAvwZIfb2yg1a9B/iw/CiNSQ0AAR/o2bD0ndl0wxTFBzS
qAGCrmf+PD8vpJZsqbkzCchYsB0/TrmmpNzc+RsvXOjXqPbrfcwvfHTggto9ezl9
IV7iuHpEDidgk501SVfyzlkSgCg3WrFB0TeQuU1GjOB5UTCKnbmi2E1/hUwiTdL3
ofWQUm9Z1T0Z3QWqxQenjr6TrLZ29D0TkbXTapmET+XrKAUBeE3jSgoYoE/mb1fu
ouYphqhPV+447Il0guI5m3WHotaKTf6xV9N9epy0Gboe4gn/WGaGwNombkOEiKES
tRSL4hWpzoDdSKEvvZm+kxXiRt3B6wuef10ujn3O5h72GD+cJ8jWogygJk8bKvRj
uwt759ywxkRuTMRvXwmy15Xs5aXzu9oM9BZf3z6RmauUPGD2dqedUEEViSy/kF3o
8z5fJY+vfr+fYOggArrm4FRrol411utyjTmAVo59Cz9BWSHcRPYOp8OnWfvsyeh6
nNtXuHNhtk1YzVdPh32zW0Q6G/QzX5Y/HFh7xLohiiQ+vDlaLr1+Gf2d9r3oHaRv
RwNI9JSlujKlajUUjZZYRJBaHIio4B0OSH7406aWIH0I1+AcCO/gHReBqtLKqNXT
6dgkKiB4liW5K84y+ee9zQ9QxrLwki9JM4hNWpBUODY6EWVAkBJf62LpsWbuj5LY
E7iLmof3Kixfg7Aer5KgvGtXQ15J1EJhIU5S+/75NBhY4rgnh4cUhgQrwjyr6m0o
0X8+DmYTHT9Z8Zf5mnDfqhqWKAIr8Jf5s7lp1scoeas2uLKkgxfd68ZI/lM8HomV
0ymxVWZEXGA+64DdqFdXOD+jWshEKelZ5z1yWpiXOs1/1/58XXvRnWEGLrSl6dCV
kftUMbvJLys4IbhhXs+9BRnKE7BIQGyXliOUpi1yaAIk1RC0hITw3vksIkrhj5LN
/v4Jn6O1BucKLnmPht7YCkjqNnmrehfTGhgVOTvp0JjYIgihX4Rh5oglFh47YSoy
Qdo2ISbhn7le34LC8cMA1gPDKfUws1A2AV8eo8FLy1WQh6YBdWt3N1Kt5ftKK9bh
nRiCxUze5F351i52mu+WIanuDKhsmssIHZ2Suq00UpXA5uDfMeI35UQ4eaGnLa90
4kYe0eFaxE1lvykUor+1HQW8vxC9dPUy9SRxUgFwBCf748DydNqbUGxite1RGfvg
R9EPGCk04e+vusdlOGuQgjcICsDG/RFf4Pd80BVpOkGJbzIzXPy20TyvhFzWkwXI
CtcEN7n3JK3RiuMsDXRi5tRt1Z/Wj6fgW8QgL0mVdZM6OEs4BobG01Uu71MwS72K
FDUaEShg5hXK80iODE25yFid5SszeqFuDKwdiSesA2g1hCcsVB/6YWBbx0/Yc/OU
YeOuLN0DfxaUY+u6FeVFmhLPs9OVlus1EZlNTAmqyohIgHzvafzw/k9SjdoacwNk
JyCmhYSl+Mnxtta4WcbbcM4vhZ30zfJjY39DpDsMVmyyn0GZDHbsMwhig5e4gKtk
w+DUe2bS/V7+7JYg5HAG0D+Wh59AVeFfEl+h52/h8/mcrgpdvW99ocmIlNii41B6
uX27EUK8nXaD4yDX6bf6t8iPKJNBiu+wDtTQvTNoCy6Xwly5H4HDmd9GJhZAhVtX
BrRpK30UE7MNX4adVUYgvTsWfpc1mFk0ZiPKhVtw6DuqbSusCB+0UMt15toBQeqz
YZ5p4dBYFfBnaMfpZVA4o93/YWl8qg1ScLDqRXEGgS6fi9IqkL6nPFeMG9/hvwyh
1VWnGAv++wliLDKOfLjYka+vHLcMvwfM/0Aw2mYjNUpnjGH1VhVqezuH3ONK8qcf
TuXFguuUSbcJsd4nVcZF7Hl8FVEQEnjej6njJQyLs0UPPKMOiuZQmhB+mPTxYtTt
dbLNW4cC7g+pC5QOvIc0Kxv9RaTO+kPMAvzhIfTlg192AowkRV/IVe0JBqPuPRFU
0cFTAX3rx14gOkxyl3hFjpGZi2VptHBI4tatOoKG0o989WUByrevbzR5/ZY6R/oS
GMoLPAy/q9XydYB0kb1f/n74ntNpS7hlOuuqJvJwUwRkQs/wIE0E65ou8DVXllGB
8Z9lMOroAs+oPT26WUgsqFWmwcKrD7x09dnoQ+/VkRxcN/gKvrk4OIn5ylm8NgAb
uA81uomu2yGvPEHlmCbTaYKmWZsmQBYnpFW4VB+d14KmevjSFINtnBuWE3mJrwVC
lBtCFCjaPOVlSDcisDpHPpTzZ7dSGRxv10JwtACDM5VeXEbjAhFO5nNvXcHAa7IR
e26h7U/tqTYT6vvxEZkUGZCuRrf+gxrkJxUM06fZmcW5yU9WSTqPg9jkXqaAFfj2
IjPiQdL3bxMS4v/TVbKJc9EVwEpO24cJRjbjaJAuc3P5w/PtdcFwVJE+wP9ffYIC
njepUmCAvyTx0mdgPzpvaDzlPhXcZR6VgG1rYFmjXKa2KYrVERaqmV90mwSzQ83X
A1KzRipHXCKPf80C6C7Xa0tzihx0MCN+v/avr7OaKZn0ixif5uJFoj8caFB+Vik2
Y2lYtSrVYqk4buI+28b30OM0oyWm1KkqVKkwu2qfhOsHbtU7pa8NHR+CYlXq787k
oGuUF+e3OR9aHq8eWbk8Pvc08tI5/aLfaNEJyDZFyWxsVe0oygj8ZeilJf1OAV9h
WnAxCg0F19DwnG2Cz3+ki4ZVlOMd8mbR8FkPz33D9GSGzKpWrvngy/2aU037AWGN
K+K9R6vggwd7RuDqQYhZYwJTCJHnaw7az2ACg/vH9jyEEctKBv6xwi9YFWuYZca+
+HQjGftEGsIvdHWVo5u6IC4S5+Tbb159RMhu7RjHVMWbS8BdHBDGxvLoY+26fl6p
K/pqT2HaZjn4XSzrUtXgi0WAS15DVm5NG6gwvMgCJdjxUkzj4WUJC4WUHCQIOsPG
nbSsXqh+EkEDBCOPC3Xm6SiTFESC3lJpRmcWct/4//S0NUo39Z6JUL+/OKxYXUts
VNev0Etw/EIiYS2yxuYLLurxpVfLLr6Gy2XYqXugosmFRB84f8mT/r1wOoWe7JJP
0Pv9uSS1dje5AWkM6iFJ++bDo1GA3NoOaxlv7+fYtk1IJ8OSiKoRuBSo8Rk54gXO
IaFH8B9B2/jj86QZq+97troDvBzKwTxN4eeov2/Q13BIWtAXjYFDybsaF4jQv5Qt
EWEn3SIJRoqgJKguDtkn0zoS2p30/r0h7DtL5IH8ssD23RF8vWzjCdKqB8y4Ublr
yL9EbhSpDLMxVH6vd+ehuuZF2SXwqefUMkVXjasLFtHXTO1o0NZZUp7UXIK+S1Zq
DGi4I8V57yEIcXWE1j9iVpwluK0vIjihP+FiELfper7/dlYBlNp0Qf48u+KQWOPJ
L0p45MQHDSS2eZb4eETI7yy1E+wfkZ8VaNZ0dj35kSrlamobJhpdS570sDoCA+qC
OktFNW47R0Y5FqeEdljMUSNdHaIeYNwxrbI3MdzU/duKAP0XGfX8iQCv1Eo0shoK
2XEuF1tsGFzPlHrQy/l848pfmtzwBX2JQ14jV72Dn9N4GZaNtJ0rDrCeu8u+xhtr
spuJUyAAiGuCWaFdhtNtL3ma49n9MQj8sVRS1V9UMF8ATCPqg2/i1c1OP9OApYpi
n+05lN3BwLJPBLZXEaJ7ulUdy7MqtH1q5BBQ91XW2wSDlvTXwYJ3RJ02v/g2m9wq
d42fr4Bs3sGWUt2/aMy9jv5wjBE42yGdIId72fSthfPajWf9+4a8E+BNlJZLqgkw
BUbQpzACKbBuG//M9o7Xi1bnr5E2IsubS2ABBCj+3LaoFNdxdqlWptGd3T7m0N+B
/eL7x3P+eDSu9IOCPuUJ9MfkFPp9JXb8/JcWzgovAYVhoL8CwwVAtS54LMKwYNiv
HuTbO+RPv9xD6MdwM/RkyNvEdPEFP110jFtAXFfWzRCywu4R4JJbyFG/TKnNxwvr
4ozFLsourluVrlde1LV16Pzsv2OOMVLTYyl4ID1zw8RW9QR61c75v1BhrIvSf9VO
jYCXKIWnvTAMWJeSGSfJ+jZJDsgJXVhSIw2I/mFKuqy3mtG4ucxSQ523MsR3fIw8
+1/uJD3UVYDyHkZbiPtLUfuZBdp/1cRCWPs+RU/GBKMILwWWQ2c2Bs8fXQ6iH65J
poCXjp685RIbu3ZNppYwRDAt+pDXOI0K3IBdUcXxIdGUcYVKQ4lmgX9WsZ/4jSmu
ByOPSo1L5TDi73iL8PjoW3tIGO2awC4hDz5cCEDJETpCvoau2Wfe9oN/ygcUrHXo
N3jb4E4ikizCEpg9G+u9dLmytAWCnfAS4L3y8qZqwZR2P8nWzzomhSRhCHMY1mki
1vJ2RfUdHYlugixxMr4oMG1o2Oa9xy71t0l6EQcKNS8UWe/jJ6VIP8bDuqnnAAc5
K8WydBSOEEN6PMI7+RUVh8ba5YoD5BwaSTpGAS9HjQ3ImgjxvCBtdQbL6fyxAeH1
9JJ2AOkfC6cxUqWIuN834Oz8BvAxWt/yFUd2KzUO/ErrbGhq9xl/J/zWmbZXrOHa
X4or7b01unjTUIOTlSS46idR3AkrSWjzktgdOD8+IxZyAvjyxyXwHiCDEell461H
Iz0zV9o8b7N7FmhJzp8di9L1KZCmi3EPqdmIny77zphs/VR2XLtDp+3rbrKVGlC4
2blxNxBc4P9CEZLdMF+eKFEBgAZVrjPKRIoXVMecE3aAeU9JX9MSJeKOaZiovQg3
lj3OqeYmmOBh3E1FWWQEnMLsJj8t6oucTw9r27xsP4hrAGTnKgNTK3+S39YB6/cF
poYg+BS2rpK4Ct70YpCdlmW5O4AhWxesiPgR5WP+mXQqfQNalS2nVQRmqWf8BmhB
RQqI7dZUmiiW9XxTxcNv3FohNwyqZHnJU3kkLwTYN9Z0fElLKRuE4UnYIhUTPPX5
RF3WJOtOH2I8jReCfgBovr/erjpPTf30fwL4OQ/PXFEO0nW67xISQumlf031rEQ/
11bsUNIMSvSNPazM/ndwtUV+joZxA7KY+qgW04SmNrj3abPSvIw4BymeRCeEH22N
qgmA7z+B6drG8pwiJH2uYpS3hrZ+mCBUiQkfyRoe7Yv0M5P/sGPqBeomBat+InjS
yNvZb0ix5VeYSy1MYH+vxm1guOGGaJKdZndMgG6YpsBTY403Vms8HLJEttnLJ6le
jGEY/BMaVE3d3+eK2X0waSgnxn/wFLNFE6baexTbhymYeRhN2iCzEeRFpoxcHD3p
bk4RyUkvsev3cX9jsp/fIK72JpM19LKqBJ2oXMomOGU3OeIAKfT7r+rTAzYCe9z3
PyjjJGUVpZYUF+9+Scbm8cDORxEOWghXjPrsK4QWy3pcI8QhykL06NgPJzeD6cRI
tu/I+0P3q9ANYdCCmzjgNazD2dP+YVw9yT/XrgCHmcljY3zd8tlE2MfSWkV3rMo1
gEJVd3lcgPeyHwetcvndj2+v7s/YX0uUBOTHMD3UHyRwpVOVXzWQbrp6OitpxNjz
wpiYs1V0qrQB6AsvfF/s3Si9TvuNmGKJj1BrlUgSzjAvmLHhQRjyLe630ZcaV9tg
6P/e+mvAklYUIUW0azfidULmiYmD6IBqke0uU3xv1P6w68ix/pJ86NO/Bmg0Z0Qb
AcHjZ7xsht+opjL7aQhRkWTbc5VijnS+iAYkGB5dB8ZSiGTjF0mYEcTDVALZD/HA
JGpYZRbirW5gGnMlzZqgqx/SebyWnJ19bzlnMaPjudmhRoEmbVpBSzpQhtpYb4Ue
IIyV0kvw6DOlQMklpIemx4Sc0RMJ1JwtFZxX5Yf9YTdK4mFHeCEvDAK3W/SoqEII
oVGORm9lDVCfydfS4uojyPJTbgxvFlOFAAdbyy4XgJqNVr93C1CpWyPdBqmoUoBp
WlCG0gKPGr6u49apCH1vN6NeM1hdVRhyrszB/Xao6FtaWJoM2aSa68CnJL/6VIiZ
xdvBFj5zrwOo/xIjTWn3n8tSjqq2YQA4SMA4BB9FSUR9AnaxkEt1cBfjapwwUFE+
sGt5BX44ZLdXg5LmOMaXxhPFGQTCjLFdYAEd1m6vy7dpGeQOCDXFj10mj3gXuiNF
ohKwUApl6M1YyblfXZ18pG7zo7ATHHHqK5kYGBJX+LsW9F4O/2RIt2F9A3SwLMZf
rT2W6MrXXYi5AENrGugsCKaVIM//qAfnh5yg2Nx48M9Bap/HI66/g+7yDnwWDCor
/s5cjQUYaaHjsdR8Thul2K6Xd6tzZH9lLiMCgng8K05Rl2tL7DyFvbx/vebmyP/+
h0HTFPnb1wA0jw837L+QfANRxbl8qnmjgvk1SJD8qjTrCtsiWfLyqq09FFATZFU/
9dNqHxgVB8kKjCSQq+8QyJLCEZ+QJH27K63leXx/WcMHx2bEYgS/V3VgAD+IJ/6x
ehwqHItL9S9GiwBCkLgbAon+khIGc2pSR4Y5o7Dfjac/mommbF6kX6ae6RChMSm4
2c3tbHRUlqH/4k2w8mwhFTJn5Xgkt7856CjrCxonLHxHI5uwCsUfxBrKX7Kdl/i4
EsXWaVN06xu2jThHiok2XuyeCnZXqwPU4lrjVV+lSlCgCsnNCsw8PRVYvWcTGyUv
1qB6oql8P/vcED0H/mA2mUBVpEo9R3+PlN+I4tE9Jb3gf24QV/IiNAyPtKgUl5nX
JN05SaGWc6PNYJRM0YIfW+lRPOdqvpHuoj3pdpPN20hCSqym9bVwZimfNbEFFZte
IqvbBIXU3xtUrubSPuGHqDNMZQrexSrJ4OzFDMmuJ3wP1lYr0BGDTzGx8oGrG4VZ
V9bg82vPg1ouAjkqWQdqfbsnqzajyAsa+usy4bWZO2BDMthM32DB8BKC3ZaG0oL3
hzaDH2CyIo5nwS9ax7jv4n7bXWAGW4CrImQdECEukI0T61jZ+YU2eaEYLTZiLfhG
LjEwndtRUtfniTZ4xs9JU9wIPjhwV+wA4Km4VYChS/S7F/xpmOl47/wjBjIfwknK
6JSYbG/7TonZdldze+kA5qTQSgpT7x3Y8q2mqc7GAR77duN3g0AKqtXIJ4rhq3CF
ZT2RbT/MlYz8l8fxiDV4mRbVRNXL0+OtMB+5dQQD/Gv5UzMCXxnq7aV33kAH13BY
oS9nH1VeucI4FouzB+RYPCB3gAHV8+zi30L+ZCeHALW4NZrkHxQMSRDWs0a66QNL
PYWdnHKjYrzXGAmayJ7Rs27JnMNhm55SFkJirJzoIqe6S0jVMZg1JJwEK3bGK8nA
6V4RpIsSTpBWV+3E7pT67kYTaD8j9wSktvlfzBxqi3oCUx+MZOvpo2U1YJDl0BFl
CXKCllVvEgV9/R3C79iFuBPD6S6xk0HtJjEs93K/NdVGbtFilYN8+A+wyAe7GMZu
6NV5ENOJoojHqX8iJ+SkREmMlmjZJ1TPZgtjHC647kxW4YVfAJVSyexOdKAzvPr0
4CyP3EwOulFUQKbgD40recJfvtjsBI+3IQzjfS5JFMETH43SiFXzmQbrIisjkIil
yd3JWy4XsSFVXrS6e9YPzl/0USNdbOpi9ixKsSvt0H5npWMdUayg4QF6Z52ujLCL
wZLeCmVeXrWP7fy8FlgOqZH7NDs9t5QG4YrGHfv/qaJ9aPLUVl+rmbJ/2x64QNLI
xqagSOK7iir0acgmR3CAbS4WsKDSwvg4eyNg16FwquGIoyrdMosUGY623d7i+zie
Sj0QM3BAV+wcHTJgU3JMj7bW0uHU6lfVTnc17Ls5y4u2NpsxXxf+s2BVlZ41a6vs
1ta5uRJ9pXtpfEZDmnp6SlPyLOJGUh75idE8OODXj5lZXko7vlHezDW27cwZoVZb
vXQYIRt9S0xm2NLOPdHAIGq4CW3G/eVuz53QAfexxHu8WJpUhrL2BqFV2CCOyisH
Txq4UWegEL8kErKPh4s45FOF5u2eaXD6tLHqA/7Vh2M6wNVClATh5rO3Jzrulsbs
os+ba+IffFVLLRJPVs3EWK3PqmNxHwhTFXfxGmER9h0Mj3Hivl+1Ied9CkdVLeJX
DT8SXBK3ddGfc6i63D2l1Mv+nz5YIfpPNOiqvJzR+YLAbrHPgmiyvqCk5lFJxqBs
VofuVhB0X8uCfpEoquR4g3q61IqbeeYkLOnznZb0EisZRtVbtbhFSOBdto+ynp/B
7MB48L/Izip+bzQQ+7L/e7f3X9VsAr3/gd6Hg6wdHBCmuHLGJJvbHVR/wRzl5SQG
10RLp/VHwA4m0IN0JbAS4Noniqs94CbAlQ8rbdkkZL5x+uJIOJjdgsV4ckumQldV
uNSMYjyMek6nqNcAI/id4Kt4qbVDm7V1JAm4Y0mS08ulNNCHcWk9MwojCOU98xrD
k80F/RcdRp3zFOBkjDE2UlamN81RLgV2QxeVm5zchymgzVlXzrtVeNbvAkbi8t8h
dzsPJ2R5vXP98mOE+QOCKT9mICvaZudbYZgWdeKLFbXfeUhsn8SZ8ReVZgL4zs8+
N1WYmK4CMSKV5ImRzAkPrINm1Vp42GCol9XRiDhjaHtmFikq29AnS1eGIByZNFPD
3e/p71BsmWbbkX9shY+DTIPogo9gDISqtfIQjazW+qDxKTPPW39ctbLoYy3ySiXc
GXImdARVh7OLqlPAMG8oXiwEsbHczMyey1MEE200MJzhSBpkGaiOhRerY9U375le
XeFOJIZl9yV3Bc4Ga0VjiNhdsRH5ZkT0Tv03cCeI2ATuUJoI9rUw6Og9C/nOSj/t
GDdhTe/5a657lzWApoZ8KN1UrJP/ZWQ3+N4hO7f6ziISZNTNJmc0AjReOz19wvDd
aA9yA+rN6/EbXbZK21YSMFbEvicsiHYPxyVBEozj75pXeuBmIedCahg2zF+391f8
1ZyitcX1046PtEbGLKMaGLvs2BPkj1Y+qPSkvgc4b8VqeoOsm1QIaYLMDFvngMnu
PPVGmw7cfw6GjRoSadgzASMiHUuuYJXEhfaCbQ4FFNQ6SI0ti96QjYLbkuXcpmzb
6OkN4ezK+JygzZkHJoRdkpdMfkr/HH4hTGb6I3K39Rlu22jAUMlCq6hfLfqV+bmN
l5lBUyXojzVm+l8j0BA4ey/T3k1aAFoyvXUqLF9Tx/LA0DjshoSrUZM1VDrMIsEi
8FN/vPNDwnDnzKzUD4ea2Yb2K/Jul16ER/L+TCDEFZAcg7Kqny+WzVCSbVlUvkq3
HhdL+MH+ZJY/4q0fIxzySY6TusZmB3ienKk3OfqLl2VHuz3MkUk5ZcKPvIidMY+5
QR7oQ6bbGWdq0Y//nohyTAyQdfbCDgchTrQgeHI1JO7U5y1NZWnP3gC+CQghMpjU
FzQuEZO4LqMmPwyqcSAAZ0em/ZSkAqS/pHyf+JiUWBEhfJlMpbQu4L3d5VJqshjW
3JOWUVFmlYqYvnkpGOCW+4NwPjEL4Hu0dBhXBlqfV0lLvCAfM6hp1Uc1ca8LLR+C
ZWh0uQRmPcwq1HcVV/ppgxLU4a4eFQGUNilea6KbsGzsa/XyLCZrEEln8L+/Fw58
mzGLEJzlUXRq4S6HFi7Bgie1YlHVIeYbKCJbOuyaJOgef0VtFMvlB8JjF3Ziqa4Y
RkKTrEdgfZ+u79RL8zTxG9439fFBVdku1Z5BRx/qduJ8wk/YQeiRfOnb8oh0Itmk
ZPVdXb0m5/cNvkLNKEVDtHeqDe5HYDbnIe3NGDDStXGJ3/y8/QaclNJp44nV3Iso
qKMcGjgtBjd4ob65C15N6sg9z5eWaPxHaseRYiRIdWUGvUQaa7/h6IP5oeqYuAky
kkZUNa6ju0eM1SEx13UoiZyLOSevYwcI1OYsxDIP8LulA1VLAI3Cbm4rLbMyQP5P
dSO0YYHeSY1S8cn+7EbfdYycGiJo1nxAIrzCCU321JWuAqDPvr+V3B8VHSEvtQ4X
7fFEGi64St1o2uuX4Tmihl8oF4L4E4eDe3AIGF0wr4eYDBxd9kVIirC0iO++7Q+7
Rhye2ShXZDCtHxVXPhGDrjC56l09OnDMcugi6ed51Q1F+VeOXxHg869TvCGCLLiU
+frbBkoqkmhoaDtcpvmN6ai92Vf5GbILedb1O62kdXsfyE8GsFSIuJkgyEwE+en1
Ij6n3cRxBjh2kA51BF8H9O7ZkAiCVn9HFaUBR3635F9x4Wju5O6AyU6diCWkDPco
tm3Pxw0jt9y1qO/mwrizy9B9CnevRUUi49TCZs1F8yABQXAT2nLWgzhK0CRGvQhP
IQiL0uhHJ5qHmC+AfyZEUptJ2WXAf6DTRkHuC1J4tBUDiOfVgwVznAzv3S6tYcdS
odfjyWNm/3FPK004MsTIjkHQnaSQ7V8Da07swmWg99hpeT1KOHhrb4Xa4Fqsx127
6Bfot+d55nUA+Is8iVCLM2ccZTSR1eLwdNAxQR1YvesRd9Jbg/8Ii2nAwy/dWY/n
6jKgUOePjV5jY71xDT5vjAEPo2usBeHqt5VZNbx+QR7LCA0XGln557YWAs/OaS0l
ySwd5D1BulF9t7n5GuAdrBK4sb5XZgsernF0giQfkv52vpmO5gLxTuC3PFnbMKbW
Owa0tiAGpS8qpmLr6vxwHtMfM3R1U4Fdp4wjaDUFv+BS+irIqEFHxkojhUYCRwuE
3EIUiV94xiH2dMpYJ3lVzwMaBIWEZ0yBVdN0TVYyvcKLB3dxJmdz3ZuQe1wq3faM
zM1Vdyw6uK5YB/XE8BzsjM2iDg1FQK5r5ZwprNRAYkwwIP22qyVNtMRGZEcrFi7y
Sc8RNHXGgbcbgsg1Hf/0s3EVheezSnGDdzWgsAD5hhzC1S6Gy7Tq9d/+lUxXymBr
Z160+FUPSik4L+YIQMs2/yzob3jzEZYMKilAhhYisoUoFkdDor0Lu3/FnfZDDR/e
GPgjkzFMzMSNNbnMIaHo2HyqU/LISB/aUtTC3/0KAatfQDPD6nQaqGXfgdzSk6xH
ccL+vrgXcgXHzqiEV4t2o90rAXdB+d3j1yHRcdcFLXxB836gbwMKG9xtf2xYY81M
nkyt5gmfnFmin8HB37o1JRT0jSjLgeJ+jqtmMEuYH9wyJYOxIMk/b5Pfq96b2vBd
YOc8k6tVzSBR8F8DHY9lmrNhAXpWcGLlcvabFea0H4I7xk6wmK/uzyeDHdyVf3oU
zp8AvS7RLxZ4oxkE3DP4MJGxNbgSSLJB1ZMGdWjJWwj8cjUnuYpAuaX1DS00qBh4
3TLU4DThsUPDRzWYc9Jda3BoVYRQDQKX6X/ZyQLdGftk07PVEru1pWrusps/pXlj
CVFfuNhJX1iMqJUUgdaG772rMjOw4KiWmSH3ZssSOcq1vODfEBXA/70RN0PX5It2
VB36SD9ede8XLmT9oDNw5KB+mQqMXawK6ICZfyMIyEK1bnIWpSOlmImJSf2xk3jp
dN2Yr/7SwQgt8b8CRDHJhA0y1qALTMi9zLjbw0XeHh4x9GMi7duP/COssUQ44ttW
WG6/Dy63a7tAwhybLr5tXhrO+yTWJvmzAJr8S9lXxstU/zNoM41sB6Bcf85tQ1z6
+BR8NBDPPZ3bIIxFqt4Q95iPV/phCiz2VlgBNkaY8ySpdR4+ZGSpCglxof7zmToQ
0YgLZ2iblrCywvWi5a/98nWEW/HR5cf1tKa1aBfVrA0bE5FC3qyHKuzxY5rnpJCG
W/A+WIiUH6abBzqUnnE+FetZREQT2VqEtNE+Zj978qTRE7L0W0NGzyyL8eAhMGwn
9+AU9ECYCraCNj78meNF1RGgc6UtarAY4uF75M/J2bZqMKR4HK751Ev3KKoJvFLU
eHjfo0w5MTqyYG2uziO3WRfBDgcMaE0w/jj52WCkxOJQ+QVPpC3ZykcboODnb5ZB
ptGwAijHfczlabK5S8HcdyLZnPU516XzE220Nts1eE47RC5szwhPj6/6zuGoZvMD
DI/5pZXtNRxzdLnJjxh+tqZVhT+cT/YPeYkkW1AbSWm1+Lfk0fyuaFbypV2Tdbaa
ammdkp0Uw1AqZGnjBOsZ3+p/YcTcytyVqYmGtajQGb9iurQldooi2jWg+DeCyaaX
XpnenanId24fVSbzRjqZ2YGB3dVrFN3P3/MEr6DfYxyfN4KjuQ60T1fE1sdvUN+W
yofjIyYqAt8jgss/gQeIEK91+buIUGFaiCfs1pVIcxAK1QQkqdCG8ortAWEYKhG5
QCfebu/Dj4ty3O8K7gsuqJiGR/z3OFlsOkguLqfvgd9htK0QcryDNd/GaKAY+yDb
C+W88yom6c8f1l8rtishVXBnCsOoNppSnDUWi6mSZb+T/vje0s/KZIFze5HKrmJg
wwLNEdaEex23wohAT+PFwfjzYiHDq2jnEcTa5zccmJ9t27EeE1mvhWnaBbCr0+kq
C/uugnujJ7ThOH+q0+g32ESnmfXnIm2A0Cwk0o8NO3Oeq6d12o88N1pJ44AfOEBZ
8174L4V98YM7ILe0TlTTICCIA0wSPn7FHaSrqL8v9Jq00wR3OQ6fxHV0jnl3DQ/D
52iVcGLMNZQ24XuSx7E5hxxpJZYKNflyP3YeOb68PLX0uVuWtxxz8SMhNTno8TQr
Te6UhwCuZ/RjNWv7kLKnwqVga+YDdlFdeSfCXDvCjoLSnO9ZMWJMKLCru+HoqTYO
/dc54/f+gonKayRc6OTOJs1Y+zkfb/PmVCq/JfwoOEyyfgDC+yu/zgrHTAm+tFSB
7m3m93l9aUGL0Q3WNpIVIrUo3Mi3/B+hEvLteZdhKn+TFDsnVauOZWV/WzPOB+Yv
Z01x/IfeS+by0MpLMIARz4roBvIlAbNCKAElncizgclgOdxmLmOV6WMC+KWX3rSN
bwvMk8hgRRARGDZ2Gu9kt7zPoJFREP8buzPbeq30mdw92bSL6lWa1uXAI4JZb+XJ
vR6Usfa4Qr6OB5ov1Ra2EEKE1AlAri7HbYdo1BO2P2Nw+xTebL3QW7k5OoSPLc4G
q7zQddO6aN08skgL6Y3T+E7eTDGB5LQTBTI9Wquy+uqCXldk9rWLwvhLvbLyDUls
w0npGe/fqzi5FKzNwceKmIcx+OI8847vmqwVedaddvFX3nrO6biRxhjEvFTt8B9A
RayMXlr1OTJ8bGRpSnVTdDWDrgbmcz+754vB+tMtYMjSRPAC3wdT/nYNeJB8ZXpz
Ll8bfLlUFql9GjX6b/pQgmoXTqPUdwrrIvJ2zqozNzQ2wzrGaXCp34zNqvmsmV5G
dllYt8cXdoxN72/1yy5Zkl42Xp7AeyKXtqpL6qeHJqmz9yV+PeSsHfZDjoyLO4bX
ZQZhzckQU+zElG/js3Wtxtp5nU9j7omxHeVWJJcU2dTLUuezdcAuks3m8BG32f4R
++UECPYNqB1zR9KkLJu9WxRiCD5llu3yZa1E37znMlY34t6QgK2MDGl8/npSmtVk
bFk0KZG1cqcTtI9oR7sm9WWNrj7J4lpucm0mDct+rY7HjRkN5yrzbQbSQbo+ALuH
fxgQII1w8659s2Si1pTpaPbc0RpSnzoiCzxZ1C5dViBtjuZGtERpUrN1nJbz4+cj
+atiW/jEvhUJOJVJNU03zXMQrqPZjHMsjaAgmnx5PbUZB9Jxi+X5T47ff2qSksXD
vL7UeB1WH1b7sypf+OGl2dDY8BuNLv3U6V6P0Q5PJ6bmpOsSPI6ErVGJagH5moBV
LJsfDYqjjmvJPXiZ5YsysV7qgCzYhkhsKLc0yuf6pTLZuWp2lsS8dG0UWa5cdIe/
PJqRfywTmtOR92wokYGrsJgps9LnRWVf5NfnINip3Ahx1dPhUb87OHd4cQvTbaO0
G4Ml67yXXCHd8R0+q8LwkAH2WFvjWfdfQCsL7rzD0+Ckaz5MwfhnxK1bWKVurIIO
a0mZyNJayluGn03zXWuC6FyD7WU21kkUCvXQzSLLiOHFOEhAlDXOBbao0JeKoe21
1OnIQ4pE9AciGrNuyh8yjJ0WhZpEThKKbmU/kZH8z34TVNT3k5ulfOlZb8nBVGlq
x0N0MUdM9/Ti/041DuGCabnaENbGHEmBKtxehLq70ieGhM1Dl3q2JOe0Xv8+YZoC
Urpy/FwSRrlmaBwPIpjI4sHh1KUBlT8RA3l7cyA3IFk+UjPl5Cu4HCLdRGVutZ1i
JtUIClFiHH5DK/KkIpxMjvZLFKd2Th8hDpwgEjimEg+w2I4eG9XBk4VBQb2ok6CS
oubJ2JjqgVZh6dy29T0fIi4n6kaKr4wRgTxD+dXnvS2du9mCLAcxLRG2h9nyAsMu
kNB0mDxZ9AQFYgLQqoTev53TNJlJenGxgTLviI+HyvtSdqfvHLV67GTuz+FKmAlJ
dtthwbrC9EGptR/h9GbOoyOlkBP9JzhyxNTgBpoHZXcek/Xgte0Sdh0CYwh7Uuf4
KjnVnT4++S9JI3kdLo60oRKwV1nsFory4ticaVsPiUsltDWghIFaAU2ibAwvfae1
KppwFxt7Als3G8/L8mtREixkA3SGDdpRLt7U57fysmchelqWA62dxSWHZUZYDfh9
G6rtzFG+g3fbS6AGsBf3m60cVCAftGOFl75t+m4DvH+f+AqhDG/lbrdjivNBx7Bh
btK3eJUchJEV0WX5KgWjIzyU94mOzK5VyBdIboo+UahdrdE+xIIBF1vY7Mzihx/z
FKDZYc8gbAekO6RmuZFi0EazrStvnHs/dk5oxfxN4r0V7fjqRjg1Y/iANdhsiFzZ
bhsTVZaY8iVQlzdzKTif+1dt+gkaFUVSTW67o1pzitk+nV1ONj/8/PX17KyeSjYU
8zf5TfIcETsLY1oGAGp+HfCt1q60dQQ9F6tK1goam55ZzjUHxymR+XQlcoe4tuBj
Tbyw4gXDbyvcKT89wRZ8pkwAzayeqxhVXfPRauzPl+1QRt1eaGyT3UK3nI1vsrCk
/m+4RQaPgFFDwNtkD4LdR/82Y1M29C5uMkRLGH17rNyv0Sjf69xcibfJhPyw53Nl
M5xr4JJEsUCK9Qhkm6L1eIIn67nE8WenvWdR465Jk5XqOcgs4kk2/rzEp+sbxN2B
2BgA9kVsCQyqw0BGZid6FHIW5Wlr4CWnCwmejE2qtBcLLejE23Gpqj0Q+3bxDt9B
cgo6QDMze1nAjydaTJvHKI8IjndqOual5vROe/Mm/W+nIdoq9F2P8zqP7dO1O38c
13FxoO4k9ctaKYYT8Q2hWyYCp6jjtFX+xScWYolJ1g1DluGk8der+3FtZqeZbvOb
rblDPB0BnEeF0okS5H7esxtrORSBACbPLEANtbzI0bBFv9Y+Y/L1oqWRe0IBKTmu
oT12r12VtJAaSJq3dj214RYYMTIcA8Qq8QMG3soIfh027O2CnZNn4l4oYreg4Cjy
rDXRMgno8vkYjCwWY82QnG+YpJqKRfkjiY9HOC7KOX5t9BlN0lTHqQpZQjH0KioR
CjJLxLckz3l6cya1H+KzcaKFLBVXoH+VwjJguKt0ppFeeit3WKfOlXk8nAg7wVVz
BRLL0GhzfhKNdh4cXYXxvml2QouMO9K0o+UxVKb1MHgYx1f93xxV46oIIYmqa97Z
T/j23qPcr9dq7eTFIsEiqsxufR/wblzfm8k+abRQTKeXngi+du8a2kXYPdlo7/oO
ZsES5rqYSv/C+U7AVefHpdTODET9Y5Pi3o41CxSXkfz0N0EU4xg/pB4whauMOBV5
JEVynKyaCAjkUml1QruZkhH0GYrsnOVRZDGOJYarp5vtw1gQu5oVjWKhEnu12jHr
3PN20uI6t83Qs+4CZIT71jx6Fv0ftZOMpew1kTTVdhpk4Ogx7T6u7u4bmhUAg6+k
5cKC2WzCbDR60CobMSeAYRr3vHvEt9EqqMkAkxMdKLELqWZczetLL0Rz/420aSYW
Zh9p76i9owV9KWp7ow22ayAAIl9NzhoJxsFepzwcjBWHxC98CU9HsDb5Nq5IUJ11
/dIUIgaDE+JZaqk3BUcxC7di37Vk5Q4ezDjbzcVPAUGisFZyNcvNmqEwg3PiX52W
gSmpO7tLowHa34yHBkxpug0r0XofRbsHewKTfavSJNYna+2y8mcyPyfjlvgHqsVd
3Rln2T+Oecx7LEOv6mjnJIYDZnIFTChXV5v4QXK6Zx4Q8wxH5VqckDTkjhchtLXI
p+q0gM4+lswDsPQnRBxcKyfUI7RhtBBJ/nmCqt3E9BcwXsq8X8BdRqRD6WhOL6JX
1u7UtTa56OTVtt9eWBFNsD/IcxIoMxiqNALRvKIVJR64Wq+EmiTpBJTQ1HFKHNa8
5p9c8DKZ+niO3CLxo0teQGli2V5hFo1Ot7V9oywUmodl3wLtuhNd/QoLpi1rfBa0
Akn9Uh6qIr4mu4SYNXuKN6ZBkw14ZH6i+Nf8EQ2uR5BgT1Gq1Fe4+LqaRlqNE6Ee
+2+8/p2vmEWp3f3aVERknLb4Yyd3pznb1IzBTqn6aCiscV+zAcpx3JguxXTIJjyW
YTsb6jGtIJF71VYYztrK8D41U3ttM/0znxud4PUV74Pe96R9yY8ZXIz64kPSWPgk
4vWDuJHXg46TpSXxo75cQdLTL3FRyfthi2EFr4Yveoj/NA01nWNSUUvrSexYz3E0
A07EVfEy1LoVFD8ENL/W9+6pndKstNOzwSjvPtqfEzRBShDxVKzk58HuRUzDP4VM
DtWY1Hp4P2bHc7eExMFVBN1nY64A9QFI+Lti48ijPEC7z37NJJc6h9uZSmjP5ZUv
ml83aesoHITxPRmu0o6tTn0iuSbn9YCzNIyWL3ID9m7I6iYzT/eBq9qwlxn4mgkW
iyrGqj3d7bJNXoJckhieWBhndQdymdudpQrKVYNxDfMrkEgDsGQbrOWP/Osr+Qiq
LBbN92DwEgLE488MddtisvMHDIlL7x+Q4K1PgVHDqkUYnf0g4oIpeXakj7iZJyfb
LQs6sydtU0lxdra0k0i0zyvdv0d2KaJtCXYoGpo4WzuNclW5SiHJtJB4l5Tt6BOq
vd37uIrPEhJ/PV9WKGPB8/GAzVusDJx/EP6Pp1NZcWcrwIwIRQVLWa14TcvnEwon
0YibBUZBGuUpN7HCoTn1L8pih/w20TdAft7cCimjO1J3otKjNw6KRDhLNylfWn28
87wCJVxnmJ9TlDSE6HgBUl41pMKdIET9a0lcyKKYbpr0HfyzuWYVu0VoxKJmYiY1
SmhbqAcZtBMd986VxYf0ugeFlMEYesUSl/+yohne3cLtrOw4lO0bRLmdRCICBobk
JCwA8N4iqq/keKuq7gHXB4bX5quAQ6fhaRbaRUWDFz4uu3nunVQWZvG4pEV2gWxF
txkj5Z+brEjVbHXq80UfLbeA8NVnxZ+Fy84+Q+7UTXqvZFnEHYAikYnF4Saie501
dUCZ096G0t4zfxcWey+RMhsaLlx+epaY4ltPvMN8fRNmnNpWPJyVyE/MjzG++Ajl
YBlStdCPNSMtrT+KQl6G4INbvVObXyDBsMpWll5vWwuoxDBS3bWthF5ZBQkgggIh
UPVSGusYLm4wjdBWQTzCioj4Z7S31Czjq4rr8pruIvLF61ebquaN/L91zgjCksAb
bo0ndWyYwT7KjA1sBCdm01eeBjBUuoop8F+domLP/dE5yoCUVDBaVh6VDXelyfrg
MXqR5rgtwLC9lauuVtzMI+ye3VRalw1+HXHtSbR31rBL6voinFrWGML3baG90THY
NcGX0BdglCRZIkR2Eg3H3n21Y0oLRtPkFxCJH+irjQQYxpp5LD7RSDyDacXvrxjV
Y6CyL0Lh5rNSZVENfmHSvhnIAGaFIFB6e/FhklLwXm7Obfh4x8kpnQW4PZCaQiv7
u0AbUugB9302wsjXJyMmOzBuJP85Bx7K7nanu2fhiXf09Kft4juXwc2BiFo5PHvj
CzzfME+vTzagesDzSj5LrgWNn1MDXGvAZp2Fue/Uuyhk6gwEsCOJ4QaBgC2gIitu
93nt48qh4wvnc8Gh1aDTFhtF94zEOi6/5ioDqEiZCmvnTsrw+cDIVHIBOkEZXxhQ
N1TY++RUhDQ4KUqBywlAFgpCgOR3zMXiEbIZ/+xiOPjEnBI/i1Lz5lAdgIOevKOp
IE63ZKSZ4NevXCC3BaI4l3NZ2AC4yzhSKSXONxLM2yJJTipfYYVbyx8goeqGBqi2
wxy9JhC0r3qbnB4XoBPFb5jOteehfO6NAdXzG7T7mvLpzxz82PcOQ7QMCaO22gez
rJGe40Gk03satBMpGnLDNcyqOZMbyKclSfuspcLfHcHZnm4rLZr7wvtJNzxzOTbs
i4ZYRXNrjVolSPTHBvE/7p+xqV03GWCe4VpeHLMQ7+1pBTJY/7zVuoyE9cVcYiUP
JdhIQJ2BVdCrx1vvNSJiF3WHuTxWCsrk8BjD2zbHfAhHbn+jQSph2YrFdTGSRdOZ
/cTWDQDGy0Gm3bnt2wH2z0bLW/3sRgihrRFJV1CpHnPTb5vV/+nRchFG8TiR4UXd
8cuKIONAN/LcTe2KpXrAzLeuZevb9YYalaO66I37xhzAssFUxsiYX8lt1+cK7rX6
hnrWViLcsGfaTMP4Wcn+Urnm3YBzprgR5JzIfQmY9gNHUkGsuzGdoeAAdXcA1DYl
kwnQEFacgX4sWWrLrp84Tzkh8Uhn98xnIBXaOQhk3lxALUMcug+l4Hso/Qy+wXBt
MqG7IQtM8XW6X9r5ruGAgi4+gYEj6jwDCF6p8UmrpOL/VB3Iq3rWBDNIX6whuDw7
iQyd3ImLOe0Y6WQjGMsF60u3Nix4qiIhQ6DUFFOCx+YBd3hTd+KT7A+WJX5wg/hl
Qz/vMa7oahPaph4NuweGfjlkGBJCqDnmXLhDJNDEA+zGxLsRuJkWR+ABYB+CHel/
5w/Lv2iLTTmekuaTXF+64olja16dR4VMbXrr7RxrAZfBzDiGG+C+mohOuJ1cevu4
hnezsZJjEklspaBfKdsR/UXp2pbhINxdAn5Ym55x3HL1SI/SZIGkX5x8cqRR+/o7
Lo7GOKqCl/KxeU42brT7QdJJYZLuk4pxqyMXTqVU2+zm+6AMv0EOVJHla6IfDZ78
G5sal9V6WNt3TrQvOUEAk7FafNQgVvJzGm0f3bBxgWWiR61ULK3aL0ll3nCnNHzv
mIuBpJXF/6X6/s6piW+zNN12uiRgeLmDYSSEhMdKKvQP7arrev/hdbq+NfmbrRwC
aNay7zVSrBK4vkiKPL/DqVjkThSDZTRevn3yF9D17ACfiLzNQIUK4z/hkmD6g5wg
60hA9/udgEvV2U0mRgJvrUq9AWoK4tkKXbrTA3kwiwSsWhq+53vHN+SDz2y9ABk4
0H9rJHywx74BsynzpySbGy00TLsS9mPa45IHaCKUCtsD/09nrzE/2Nx1HLrMCmSi
mCzUb30+d6Sh+CQ2SCb3WP8FV7llIIMk/ZK4PtuT5py5VooBX7m6BCQWJa7Y6gAW
Cn/tqlyfeC+m7XK67ZdSUSRcyrQB4fxaiM2CjvQ3JC+H28L06pAuEw/DBppd+kQh
4fcYKkOjZ/j4Ed5mD+s3cmDTW3vRCUghZCsibuYHwVc3VDJAg/nO1M3SMkUd+KTJ
cU5j6FkhTG8r6y+9orfW18d3TL1zhN6ragrhAWPJzXu5zsbnUJq2L0Fs0MDgEf+W
+NE+Z5K/yEoExa9dDKiNj2qlTf9bVfDA2aoRbgVei9pOj2YvdfsLYy5PV8RjxGhw
Lm2qnko0lAox9frbeBuZdt36D5mgR1rP1UljAGUZfdsmrxbBDKeezUIeJ7u5lRj0
JSexT9zICBBIesTqZaNFMM2AceV2B+mL7kCSD3XpWDe5EOzBONpisRQt9o/qc7Gb
kztrPfII625lkgCWdLWMvbZeM2ZQxhKg9QLO5wkkfL6HLUE4gMsN7UjUxP7cmysw
K6aMsx25zZW7nMiybiLbhGFejMoC2XDCEy4oOiUm294Usyb3nuEeb9uXvH1Q0mPr
KlgeJoWgWOGmYI07A970+1dhdWianGQfzZLzeDPPWgMXaNH/T63FdhRxprTpvTy/
kVSS+J/j2wkT0eNH3LPRc3f1inkQXwzxfKxTym2xLCf36mNuA+qS9z93RNCmizal
jqE6qsbaQp7e2dogS5jSTB9dlOcwvTOm6E1gXj3uvDKERWU81JU8PCyeixDrH6iO
SX7rQRb1ipfyDrM+Rc1279Fv1InozzCX3kMS8TU6txqUAw2YzEAI5Uj4sHTGf70W
oy6vOfA4MAJN+l9xbs1Jj1TJUxGOkvmLUbMua4QhlPG8ECe/2pvew/nJpqv+EP+/
SvbsFhMe4MNiS/USaNA31JkmmAE/5vXVb48FejOx7USAvxi24+/Jd9QQTxlEesiB
DdiMkq4ZLnL7YYK+wTcPM0PBHzl7tU/L2JKfUsQnPxGq5pT8JWm5Mojd3IeAaNN2
ES8UKFVrc9BfNEMsybJDRMhi9WPx9CFZnRSynkk7nJWgPL+JTQ7KOs0iiButyh3N
4MTb0FBfxcmVDIbNvIejJpPliiR6SRyd05brHLOwEbDr+lH8+TAUr64NwITnvxQr
TpigAxtTzF8CEJtS3LEDb4Bt7BILstsmcPWF+zy2PGiJFogGtG3yLgEnMbai0Soh
VUTT62vfYjbg4y1B/ji7MXSSzi/15g9c5g0UV9u6XlGu2FP5SHwSn08mvvB4WSH5
sK1n3Bv7WQCjD44fguckWM7NxEnWf3+EzHkLqQgyw6q1Dha0FrWDGt6IyDoUN7FI
0Jwl5klNFsXjGtjT9+2I8ZwURaSPrgSsOOADN/RFdA4C3uVsJMXlTcBeXlPplyno
FIOyoKgW1K5+RuMv1Ll4GTYb4QcgAT4TGapmjdmkeYKhIWu4OT1kxWzJ4+TndODK
EzEoYkMHvGw2XpX380OS78AxX9oXckCxpkappzP8mIKMVQG+wIhfTrfyZ4xVtCUk
+dIuVabLqdx4pdwy8ySZi0hWb77iKifFBN4Oawx4+ZbsSjyXDEqp3hgfCxa87o95
NsWkPKR/0nzke+cCHpHMUnH0lBC1Tm1UFMfKX4cSQ7qarX8GfDqSIA8HELPjqWqG
25RXHkq3S1rTqP/smcku8L0kPPNRbBxaWflr+G5OtfJj2J2GHB6zdpIdy97Izgmi
7Up3D99nvfZjURcISZcsEEq0D7H3S9aGasHWbkcjIm2yZEvGvlJHo71rqtUJf7CO
gAYlfnFBlpikhOj69YkmzbNtnOxMkt2a2R06Zoqkxg2SHK00SDYVI8HjDe2GYXDQ
4QweKyk9Bowic2Ex3/7V/sm6hPPvDJ182ugQ6tXesW5DZoCE8a/s3BlOxJy0+0Hy
5vjueZHLlaHJqafp9aPsIyy/Bhhx9DEcbsGIMiiouXreeBcSgGxGXjFt8+VizL0A
pIqibv+gMRLSgkSEZ46iu8FZSLPuiOao3rfZfPmFL5Yh4F0i+p7+H1IGWTVokP5Y
cnIcwp6ViziH5ooaxDmdjURg9WLBPCTf/r+kBylvvpXMYwxcNBuooBZmr+hYn74Z
bt/SUJleSqZcCC7fx4daxDVAd6Adb4r9/e9iKLH4pEMZlgSTLGD4Uy8erVtf+oxi
G2YQyvXGYJkm2m9jul8jptGbZJs3F1ecZ7ZbriXpX2E3XnnnoPfREBP1yVdw43Xd
DgelikGEe0UCM8JCMo7at11Je/5BQKtX2VnWvVAQNii4wyFfMWo82ix9HtLb/WQh
CAjoqP65G3CvQUNUyksZaoOm0nOLHt2MISaRcEbZlR4Db7yaWVeDwDGPSfKK5zYC
sv1tcwDjLkHt1LNwt7VprzEej6SGyU19RwMvWGq9nJpTQZA4vBgZb1o5dvDOK5fe
/jKWHszeudYGMSb+9Xt5pGwwWPH78cEGvom9dXrQdu0ChG25kphN5BOj+X0operG
9TBxGTvnfamVtNAPlcsAk66MMZvbL+/4vNJGhDWdQObY5KmnA30BBrgIRojrplFz
DmoUbZHV897SOOtMFRutLuZKOtz6X8JRziJFgtT/BmNJENsZXWkupbGzBGqBJgs/
l3OE16E4yp38vg0J82iFnmsiWEWxSJTFDCd2chd/FBKAvpiNjFk4LGWKiDxf8xZG
1+d8W9+omWYOVD6Q8LxopclguhO+CuQFtA5SrZ0HQYoc1gJzkkfkXZ4WMA4QjJJf
/mZz/eokGlgvtcGVuC719v/f0SUGGc+sKwxXsyCfjx5UL93byU/keoV59bpr4qtp
IJTlC7i9vojTGP8TLetg5ajrAAmMmlTne8dXCHJl70aIFsOHlNEj/bsnRQYFcFBJ
XY7DOBirPCpGALEGC+cG/alHv4FlwyvXAg6tW0enCsC13BWPTu8Y97/p1puYAfd8
qYd4uZ4lxmIazlKpCJc49sdu/KCgu930XbRYhagFhwAnULWGMgkuzRbXvEkI95MI
8Xk/fXGiFlIE/wyI6av0uFLVyzwmiPwa1kq9NDxtozZmHJqKGi+TzbkmG0E73HGU
c2lcoj4ANO4gnzqnQ/T6ll8qi6i0+AuU5Jo20c0oqLf0qHR/XRiIcuciwlLSsYzY
I8j9iO2M92BBJDWaZda8gcNJMc4d5VvvGvbXucasUQRRsRgnicKqcZQcd6lFSXmN
blAphxv37pdnZVa1yH+h2/uGFS2mPT9CUiGm7cpJMgF1Oj8XooPksV5oH52NhUYB
HmsO8f8p04+EEggFg8m27nsajycJ7/o9aKXfr5B5Y/EE7PE8+xIVz9Ke/Hb2g25g
yLW/2WQeARBO92WogMF6bCNrRYQX7Q1ItUaiD/4L/DpObPXOsbGrrpuKrTzdV/ac
JEYD5YCDUY7YbpQ4Nm4pX+zYjUo2RUehM6lBE1hr3WktXQr5R1/YaUg3qGmTowzk
bLimoZsDBwDvqULoy1YhjrtZKj1J6aBPLTTLK++LkWOj1br1nTwoJ3iDKwbe1Wa8
xGg6CxFy8f6sECpS92pUYowKMHL1hQt+5wZEJCSwrvT9vR6Ne4JzDx5C0plWk22Y
R7moInes7C/PhLOZ1mNA+nlu/V8gyBI5kWJHvklVEfmRO0WuKDGCQU8EBfWkRLxs
hKyaOH0wd19QV21gXusrNFYGqg+EnM/ZRDVzxGDf08pHsYTylWdFzZPPHRQA/aPo
HsVQ1N/wIljerPeLauRpOFAMxWxbAMmg5lYWRlV58fOg9ViovfZRe/mObvJ/6OrX
3jCJ3kuBiJkIQ2YLTUODY7t+NVRx6V/CCNIEpcNJBvpMIFnMxzU4XarRpxqZ51VD
bnnmOFxW5RL0es7uXuPMzFm/v0Ct4oQJTISM/YHQG/eOMT3K6rNbGmYW5VbpwNlH
9ycrT3A5vW4FxT/tJ4AIjQCfLJ4eMWf+QT15iN+hOZBIbw9GhQfhEhmwwBNd2CXq
t3Cr5plhMtZ/wbplSrOFc41Y9FWDZ4npQ2kuLVfD/3NYQxBphwQSr4YH6mgZ/DNB
QLhOwqZbnRN1ScXvURrJQbfXnJSNDPJ6Ap+G31LgvJ1cxiLZejmSHD1pTiu6kY8Q
w0aQnTqeBIjXgzK8x2sEAsYTTswYtOEdshAP/7Q+d4sJphjzNBFN1XFrLkOIVoFg
s9djNgfFT5Un2Gz5cCEzQXFAclQARuK82h70ZsJOC58dqMIl/mldGtSYRuepbVGS
3xqw50hZAnV/K+wFUrgDXz5fyXl8qOTGNvTAd7cTFaYNtOGJqoxb289Qn5SERgin
652ultMgmOo+i3IO0MlzNJM8myLaFighYsLAmBC36Uij6rTu0aWqsUSf1Civsl7D
XlgnQcEku+Y+nYaHJsWUXoqT+stIqVN8Je41qJ96C251ngwwToIQuHSh04nRdn9x
ORr7G25I7z73iXKN5VLXYBrQ5bGGIXxsacGFfIDhcF6ZfpgBPdvLph7r8KlM8YDU
0WVuFEhxI0kuSXzfdW3szCFpOwrbA1gA4pitlSZlhpiUp39Okc6FHCRyWVauxBlf
F9tF2R8/ifLrULN+ND7awI3u0gMiS164gTIuB/yc5AOfjAg1NyVK2WljTUSIy7Ol
r/h0w1NrsSavFRv1o1O2NSJKQ500wtaEQ6sxd7ztl4fs33p1MZoYpP9fxaq4V7YG
70aFmwDXVE60QeDEW8sgvt2kIaEg3M6q6GLvWtayoTU9cBze9SA1T5g8+cX8t+XX
oPXH0ZuVeB7g/e1Y6x7gKmHxqVOwqkBxRKY02HbKji9pbpfI4hA3kIFN5P4KPlgH
v118a2fdFFxRuWhjljbc9yFHSIaxbtyRvdlasDYqmZkDYNNPA62tiY+TosurD1tU
CfV4OJrJZYfGfQvHUzjXuDoUwg7IY2D+zkyrnsz2wgHRyBmtB6uz+kcIFngarUF5
+GabHo5jGE67IO+3+pZF+KY+SVdU7C8lPskyDM3x9kkmeWyae+LiOl+HYC2t+Mw8
hKxwaRdDfd5HzDpd9txSnJAqnRPfJTO4NQ8azv0VaVioRNs52tjli9ZmBqCokFu3
feipnGu83cPUASX57Adl+1MYpP1payBpnXhC+vgVFApMNrgvXsiVFe3S42Nh7MQl
O05DAXPn74d8dKwUZooVAq3o9V55AsHm5JuCWlfDQ2cGQc2yCFe+LKU5dy9REL0e
9KVyK5N9/Gq6d1IdIcQq3xazgCd52BZpWIBzTFeCwOcmx0W1TsKl+f5lhaKVZHpm
lYgZfR3m6y08NJWXREEz+v+2EHvKlkGQ0AoxHOg9ECqfMFRWeiAo/9Er7Q8r82iQ
65bLLRdFHV8INHe3kea5Uza3qTdm9jumoXIITaaDNmfnGt2hq4D9P45g+0OQmQpk
sQmbkTqVb1vR1S6P0U8ugYzNZvd9Ja53vWi2sCfhnTJD5yIflDGmiDYkTdQKwUAw
4/9oTsyTscI7kv+jtqQsYh7dvb50/KReMjo6+h1KEKdqTY2XsNpu4DZU4o7NmBRf
vGKM6SbyhjD8Oi1l4VCtruFRjZFHN6aXfqFBVEoOGIYiGgvrSa2dCgavEbDEiMoJ
MXjNEqrEiGITfhJ7xAxBM5EPzn/6/9Gu8nFwVbBHDgNrG5PVU6TTKsUR5SDkdzCz
oyJQqyX8ANmKrr19ZDM5m3z4yNSL5NmvE1u5ndv4z+vIkEJxG8AUxD9kOuG3sIH4
ia4EGMkfOtnLttKCQ9wp3LbAzGpSjN1xUZshOCBLw9SUOx6t1VWO41FBC3kzveir
kIHWEwc8QwOImcJgLRd5Mh/EFvGSnUJOigPU5TMHcFPOasG21IlA/66kqH7asTay
ZQyGx3kVi7mAfU9ci2ojmUco8KrM8+fHfwCP1iBC3M7EjoEgLBsoPVUL75JczB6M
FtW8t9t03gBKrEB1lkh6FNFR/s+z4uaNJi2rLBKx6OGJkWhq2n/MXiqBDWaHZM8o
3T7DPpmlmDoy5XhRggK7/B6KIcBubpdPes1zdH3DVkPzl7iKn9m87dLCz5cKGtCv
lO92FiI43vI1en35NaOSApRgTiQTAdki1kAQWQb13xdtoE8Ez4/YEPLkcgBNBbwl
AbKOfYRAnwMR3S2DdGdCIP0xvnVZBSn1VN2FKwJVSpXwidx2+cYspPX/7gaFqeJh
r1xKme17Ow0Os0qkVuIhvxdQ3A254Etd63apDYN5Ld5N5LAQ964/Fa7ObkaNUAAY
PEXiERrUaotMaos6VRkDRW+7rBlDnmN2gSQXqqs2xMziBwDWsor6s125qQhdeWtH
lWhijRAkqcnP8KSNga02WsUyuPm1V+0AdoY0tJ0GHxb+DKVsEQixx1G1MMgZ5nsH
`protect END_PROTECTED
