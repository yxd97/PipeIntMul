`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0A1ESf6LpJkOBrqaABFJD0uUoovUZP1Ax/caKBOTkexKy7b0bu932VnJC4PuiA7G
/F4xlam312hxIwVVVo8Kh6HMP8OcrS6iux4mFWrKgUEnc2G8cq0imaSgLZCoalTS
Nx8yyIg8E0EkNZG18FZWh7npU+CVKpj+KndI6eG7Wti8gdYwKoR64vqsSby1WBcK
s9F+YgCopXT6ODbGU3UZjYykEFrNBB1MSfhAYTxCTikkOQVch9FPpamWW/niyHSL
LHcgKVppo/zbxAkmaTaN/WoXLo2oeQHppEdxnv0HpgWLQp6Zf/uxk25weDxSRZbs
hl/JxBBMX1ZPQpPF2G9+r2wgeqUXdoUbz6c3wJ5uu0TCfvocUVgOjjUVRYZoT9C+
4Olq5toieiJB+ZXHi4AFHA==
`protect END_PROTECTED
