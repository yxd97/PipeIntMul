`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVPSYeJJsT9xlmUMckYVoHUgja6oQZd2jBEmqQZrvbjBNH5+77GDufy2CjS6nYTn
1F9zdurJUCOTtsqEDX1by5fet81mqmVaTD98q2g1p6GibZPjqkhlzlcA3NjE5xIm
u3MSk759J+H2httAAdEKhGT5Qtcf0hGcDAnkvIVokFKsfd/Wa2ERG0feSKYyDtF8
l/tVs+UL76H5cAV/78imazel57+mMOP+X45a+QjN3lFfe5LYr1BVUluHPY6/3aTj
VJirJ2rzwA5YFRZP0qsUoPWOYXaT93bvGzGxuuvon+LbnPEhWkxXVpVxVuZNKMVe
j94wUUi8uMoNGCcc59IAGUhYO5ZrMRv6dFMNn60z9pluzl2waKb9x4FE3JdCqJga
HyyEM4Qa2tambStbWgK92bkgOKc9J7Nm+QFs8q0/JnCL/Aof48aA4E/cdIN0GIXJ
aIH1q9Ayj3gd+l58qyleHiy3o2VUKNQRJt0H/ExlBTuSf80uqYsWgAer0XcaZusB
/dUHFsuZQ5ZtRgqXdPPE+xs6hQQE2eUFiBvNy2pVvuWx0vyOm2kqPne0TvA4iKGV
`protect END_PROTECTED
