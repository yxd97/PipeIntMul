`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r7+xjWY6iJ3fHoLuXuFwpupMgerbU27AX7kmHoLxtsX+3lHtJriVUlVpEzf0NAK+
b9Rj28jHbvDiC8rj6Khlg4JkOpv6vE9PmPDIlUR9bMtNAIXVGtT7c+cFU7IzjyBS
Kob5DojE/NEwym7HhHfHCvi4PTOJ0Ihq9NndjAX4ZtWrsyriV6z4n9qzJBo2btVf
jOYX3qRvsiPnLh6nb+Co1t21R0kAhXD0HUOGkEd8pYDij3Il1U4lu+YMt3soRNv+
i3maPAOnnxopSccpty+B9m+d8ZV8D4fmdTS/jU/poGm53rri1pEzwN+PIQAFSk6k
f0IYdNW8VfUewN3r8ghkRFBWskLlpGdxvXjnG+RsalM9oy7jH1Kj/m0mIwrFEhnh
091T96Am+/jKPwAzDb6gBpLZGNyRpqYxr0epPzB61S1Df3bAdp0tRZyg1VuJzv45
xuCr271FqNvEKgkArXvvgaxfgassqQhQ1dQsLjzLVbXljEqPuyX2iHU8nQWDMMo8
lZCf5Rk/CSGbHOv42lr9vaZFAWKt9ZKevefuZ45Pnz30XQLojsmmU82Mor+uA5U7
aFV7U6C0c/u1JYQsG/5oQACjk034+T/vjPAzQ0lJsleIkFgTGtVT2MlXQcyvOghQ
MDJ1oHMzBsvJega0WQ5OV0qlk+y1u49jfenzPQx35BAmKGDLIma8mOaJ4qHAxyj/
HeLeNZw6nFsVJLbZkN9VIQ4mE9xb6zzn2Pvd2+EuR/Qa3woLfij0NRA4jfOU449m
l9wmhVHSa98uB26tK3Xc0W1Bkbor6QseH06VogtKKkpUvVNakjkaK63HgqPSmuZ3
VyTNfOz+QiSH9a8rQxy0WovTUF9D+ZYLhjl1abdYoLP98JaHTy3VFMXScOiaM4DY
OmiVc/JnUQV4PWu86XNVqvD0f3its0/EUwYk3V2oxR61+3bUDgDpckQ+t6HF5hQa
IWyFnZvnro3TtiCuPeFdgvdKkSOgzAUccOoHPJ08x1byeZidN2y1U8Yx2U85wjmD
5XdjgOZPLWjjqtOmzLhzfnUoywyqzZE9RsjLdoLwKM9BPtPh1fIcK6/U/MCdJSd7
Zy8D5u/R38Atdl3Zc1ABTLgn0gt1ZHayrPjN4ac57VOE1eZfPSe1zCqAiUR9e0mk
C3JIRcZ8hZ5R7QnXu8fgAxxuSZDWA1NMJd0odNcuecZZGPtY8jmq22ksZtLMvfxx
LnUiN2ib4YqZ0+Sw+8xFIfu3XpU1NtnTKfmhizv2C5o6GBoqNp8RdcnPJAINPOLb
eE/Vi9NK/VLN/hdW093PKIwOHbT1j3zKIc5yP8rcl/TB8TwDCsrDYuVMyKeT2gxR
MtVyv4dx6OcCfysIl8QuY4IOqpRRbCtx+izFlOI3TnVHi/EXnXaGEoUxoQuUi1zE
hOMAgLnkczhRKb0iweNIX2wHiqc2STbctKi2AG+j0rbnzz5ldUCkStq4B90gJcIt
eylHnd400AeX9AzEXCmh+72H6se9tYZnw3xnjvXdpRgn95YA7I0/n+1aGaTeC8gj
rttREcMoWNTIb7Fjo68gc+sBHOaE/HK4sxy/Ly/JvRESLdGhemuuUgeAV+czSr34
aZXecHJtAgKlKrFxtwJQWBOL5YicFdMd3JVRoYCeJ1pQbf5JJm+K8rhGv4rUBkEM
Oyj0wJdTombNzjk0dHsVzZYpUEsXffeFjGVuSYSNTGbfyd9WF21TsNLVvj3Grlvr
DVIftcaYADcUOc3R3t/1zKUMHrkIY2Lwt1hVrSN196s=
`protect END_PROTECTED
