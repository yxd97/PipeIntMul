`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqEF98CYNwdKWeB6EaFoD6uBMu0z/kqbv+61fnx0LkhzWPQZZ4XmTlWR01FTtOoZ
UPYbUIIK+faAbvkHwHRTdeaHDujWkYUSdTdAL3z7fXkbB9eSKMTJviy8490ObhU6
BlVmNJVpAmyYbuWW3yVMAJRK/9bDEGfcmur0z4GSlrZb2wqOFmmvBPd8QbUxpzWs
vaj3HHxPr9uxavumkIZ9iDuhBoSc7XHIlnMqjL7f12nNnxcOSiu83hwdKHgKyacZ
BxV9gRJSqJ/fKxOOfWMVTRJHXny5gb6brEJhRAt2vPcbcbeiK4ZG1G5GAIOpzNvQ
kE+w5o0GLgT90+2PLAVy6Xibg63GI06Ac9J2OiMmI9xpHdqF7UPJkDbxDV7mpmUb
hfWJDFSw1YEevHFgqH8hfal8JKGOmS0FZrcPX1lqBPoicXF+oqNAfE1zsv/aMJ3e
Bu9mJcpoqJcTk154yyiXc+xFrEdQaKW16KMz0oFayxXn9X+RsJE/6JnEmPbGtTYE
YYgb2XvpmCJmR0ktcIyVIZqNi7IDAhodwiaIef6z67J1uJxWX713jg+v7eUaJRUQ
L3N/spkJVSLmjXd0lRhUCWkciER2VbvMySek0pLaq9hk11weh8QtplV98+22OKc1
pOj9kAhZZGXIfDqjbjmZ39nOivmfBjdl7lCVVx1YRRS7ehpXOWiN6tCuip8Tr8rI
sK6ON/KMWSA/6GIkmH/0SwAw3Mn9s5/9GWSitX1uP6WKhzGGL7WymFHjaolto26h
64VLlSVwCNFOTU8tRcqNoA1u1aTUEmispJKSfPb5KZzWNnqvwZnFb14XDb9Rnt8r
vePTyWbbkNqH7e5CSS62o8m2byY5xL6OjOeJD5kwrNlju9nkP1JcfcYTi/dB+KFX
2A/MAWVER84W85oGuKhGkvPgbf3NKVG6l5GCs69H8jQgbBaP2bCjAlO4Dk6W3AAh
`protect END_PROTECTED
