`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nrl4u2FB66rtvsgKXx1O873VrlofFudKK9VfdqdYRJ0hXgEjH2MJi0oIK6nEQcpI
VSrDg4Gff9TbJIcxGeIpOa4XPZ+rmhO2cfKGXOptVw2EMBLXEQX6mSRt0Bmv50xk
S79gzBANQkRK95A62OfX5McCX4wS6aU6BsL2SpyGBNrgkq0T28bNeimf2OJNZhh8
4Qg1OIh/MNexYuCwUIwl2vl/K0Rt5ovEOHApu8TOmn9mUOH2zSZSiMyK6OqO72Ko
PDPPVAgOT9LcaCQjS19DQY/Dl+hs2CXYEpX5vDgbukIaw29shQRgy2yClObMf5VX
vgS0LQGQUF6ZzFvxky0umOHrVM4NSKESv8uYSK8xkuP5rn3BqmbJ9EF5gfWQZa1L
08sa7w9koOgQFFQL3xCyhg8m7X/AqsO5kyhjqhZzksRQGCRUxe7szpEgrpLKWdzD
O3pAHB5mJHml/kskCB9jMWZvciewgSWx9AZCHeChsgoVlXn0sqtW3oDMIemXFCMg
dqoAOt1rKgr8R0hcDLAcBwd9We+R8AGNSZ0UdvWJG50rHHI05RTT6PXIrdkd4jtV
BdNbOWNvGcNQb2szCkGPeA2Q2O/bpKEAaNVkEg5uincvp+2DQWcF+LGzQKFM5Q6t
WiRTqVQtKG0YR1+H4aH3VAxnVZ+UhyuwBR1MNTHC5bEyF0XDsDktMam6/VYMItrk
OgS9kXD+U9jT/XhaakPnzA5zWxC9ZZrWCOZX/AgLKgRO8dqkaJlFoo0ZNbySlOU5
y7KvXRc6wQ84lH9dCONnRiVXDma5LkUUh0yUYsEg7D5rAvnwVk5AgoSaWXRaHHkr
d7OSB0igzRewk989q3v2GpldwGwFTjgJzxhtbgeIyyVYpEzimFiZbMT5jsqde4OH
iV0iTGVWiW3EfLGp+PVYohWFG6qWwVU6/3VSPVQVxzU=
`protect END_PROTECTED
