`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s29XY1U6XYOSI1E1uArb5ygnu/TfWADBIjAANonKsbvDsQTR/IIKnP9Ny9ygDfgx
0b2pkQ5LSjujLbaTYz81dftM8kMpBxOoV8L76Ta52/xAYsy+VUsVje2l3RyK05nM
Q1HJHri5EvvGpjk4WTjPBExKgQLpP2zxoomIMGVA0hLS79RyRk9QeHDp5XYw4Qvw
LV2n4qigimyGosNHni98mYwlFrddKgsGm5XiwH7fjlhW4huwV4Gk0vo/ued5vEC2
ol5bfmG0aRhWScScmHlysJQbyKZwZShhE4GBj665xjJ1XZnyR+bI9Oaxp9lV4ML/
oP37ajVB0qjBeHTROHPfWFk28QTpexQMUY1KkiPIAy9fqeFoQAn6/mbRP6wWTyV+
1oIrznCMoHn6qgnOf3sEjVHbiIW0+891oBkx38Ad6PIyZSrqkdUGxhMF8cj4Pf2T
KdKDz0SIJ7t41Z7dKtMAAlZf63gPLz+QrrNLBsg61mIopsYhDJlAHLkKZCJb3rM5
rev/YXfnI/95OOP7CeMAOytQYHClXYPm5Z1fCQ5mov3U0lLfVPepr6czG13Sddb1
S5CLsloSIFm0pYo8bXD1PNSup73a8woGziiPZHhrbEraFd4H4xrA5c4Y8LqFruNG
Nr87Y0EC+fGp9zLzTcY6jce7aO8fm6NM05RLM5WXDNiH/tQNb2grVuNaXnl9Gymj
ffia8R6S01w0qn0glvCpK6//DtsQ0QKBJciSTAuXZEChbTEpA2xoqgBqlZ/8itg6
h7ZdHkYZs+NsvUpO8lARcW4GYthmaE2IerZ8AO3TKwrX/AKMXnxA7H6lMdro8cAu
JSxAzAeJ3ivexv4DBoDnpC6t/racArHjT1llwt+WdK0HjxMyNG90xtEeVWLUNIRk
sNYoniNqJNQsoTt9Q4ygicl9wZfcFcWfrwb4LEM+AZH5RtSjkzgPv6vlGlppWJ1X
6qXXyMgECrEwdqIz5KeeAzGRdCw1uqoUyULottqVKmM=
`protect END_PROTECTED
