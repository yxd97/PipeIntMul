`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LUMCDa4hHMb8lXoNNKCFJ6mCzx+dBaroEyAcwXJJZdRna2XOxQLa/RARBt1H+I8D
O+UO7JTod1DS6c1su5Wicx/Mn1fQsZI1qkyq3rujFEhrD6IgSwG8zYMh+I0BKGoe
ZKijdAcmOXzIkLY2XaekmKcaSiM58D4Kc9WWeO7d6LX14/2/CRAW0/PVT0MFeujz
Xqt61xhzMp97tghWZiLFbIKeRWD6y0eNz7Wigx08RFxzvJfwg1lTRsEmhrmLsjcA
FTKq4tqZgFebCGZgqNq7U40ax1KpL5P1KlVSkwUffrUR8g1ReOlFhbEydq8TdZHJ
k9ek9R8ORee1FKef4mupScFd/Kcn5+lvuMcQeeBQPqBhbaGzry3MwW5g5JHqfJww
7q7OjDT2snzC/hc1+UUDAvBAC/qiZgHEN6dq1VIIsaN90kWwhk60gUSbIrrocKr4
`protect END_PROTECTED
