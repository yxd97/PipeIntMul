`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wpas8D5uaY7ELHseU91ZKaYXShs6G69x6m+Gd3Ky7nOrMLnhuTGrOOyEQc/4bpMA
0qyLYgaNWqhbCfAPsxc34Drtl4a0W4OTrMDGFeQGrQOX0+KM/v6o/Mvx3faMDnSo
2roelt4P00I47WX08HqmKrnAewgFrfWBuUqMJsHi99pWgO9yVnIqb5IAzxm+iTJy
hhMxNnEZMH1/HDWHG9PfkzjOtcZHONDTn0yuUilmushYKDdDqhj4H1oeTTRZ76N0
C+A7moFya+FiWwyoEC0rSZwOLg65AWDo+jW0g7vGi4pBdherlSN9Va5yL7bhVLVp
VrJaPFHS+4m47FaDp/zQC8xE3bLwmzu9YMGlkV2vspSf7afYJRi6vTTwOby2r2ji
NxqeJXJPtCtdhYBhZ1TBvrAZH13U6lVCeuqJV/xDca8Hb+ODCjoukFMtQEGyrwZ8
gp4Yv2C25JtDhMZRq+ckT7SKfJx/n1DLdEUgjw5soqIR8Yy0vyH76fPUZQnBMfsD
ozQBpl2jz8c4oGIOGLYRzJlcelLdX5F9Iuhi1HVEZM1hmaQfoIjPLLoe2IQMykg8
WD1ONBA6gRF9bF9VGPh3QoIBm99Vgy4dBWDUfBzsLZ0e7jMSdXeAk4/5wo1KfayT
O1/I3RA/jh0HBwfNpm8fnwx3XzrroMDob5XBLdLOcf/kGPWqy/jkFepIOd4MzVwM
QI9zPSpO3GcZpzQ62icxCdXjATtX4twYrC/HfnDXsJ+gRiNk9rgS7Id4YmOUBLll
43Xr+x+nnxBtRn9W9WU9M/X1eQKkz1ggvFvsn38jlZA+rKaiXTCAdku1n35FEvG5
4LJqeFR2cV3v7K3Crroixy49lofn0sBXdRfqy33P18cdwzkv/hPV48e503qKd09W
NdsWTodYQGdha/I3W2nn0QKuik9ov4Mugcg7lIFYDMS5hzLFLkxydC8XYLpHtMuZ
7E01bspASEhR741XzQV6QJfjp3ahBn7OoDi6rQv4rk1Xr+9+eWFDy0ZHF+NM57sR
kkZx9GBVCM/cLJiRjOa1OCaOMYmMHW375zNuQ3SH16wv0xMSri4MGrM85ByiZ7JF
mX/MoiqnymbMFsnMX89F1Ryexn5LFytUvB2r8IWQjNAydgcfmcVmgdNFIgMjG6yB
E4434llP00ER8szHVUlU0pGzxWlEi1BRsYbrkzwKuZZyjrCDXby+O0Ov84n4/yuY
Cf+Q4VXL6hlbobXtMlRks0Pjbkt/Mo8ZO1lQPKOjAf4z9d9DAIxR/DSiKUXBpB4Q
MEx8obW3cuNn5vyKMRTETkHk1GdMB76I9KMOgLBdXpl+0oi3PNPkB6cq2HbK9IeU
Q+Ri0ftv+e8G5LYVUhh1autw9BMWhVZpe/9HEMqEyZtteJCRgcanVOriv0ESki26
LFE4TQdqY969IH6qNM4IPEZ3R3m/hjbdhd+NqmQ6LpgME/4nzaXwaVwaRojJuwgT
tmI4xyQWderJVob6fEOCD4qbwvOUwTm4yD551n44923C9Wz/V8maPEFsUZk+mzI9
oGpyKn+Ag3dkKlzuy+jdJTv2hyE+Q6pVuHd7BXmcRxsmzKP4ihP4OObdVN8eVaP7
Ga2kAipEm6elDlut7GPV1HpE2gtUHjfRijh6HVmG/OdeMDQ+TXtY4aodQyRWs6+r
fge6bz+Ls+nitYxCSD52QNiNJTqTLoJvZRD7nybj9SCBimaoS7NBZLuEw+AIiO/Y
bvdrw1Fga4h3jM6GGUF4WXYesq/NvrXDaW1lX3f9Fy/6AgWdnO5lT/of/LMOAZPK
fYpYHy0rig8easvqrdM9b1YW1e901jGn6ghndWa+8x5hEwSMRIF7YDwMk/BK/8+B
15Rpgonxm+D4durCFHD+Zzx++qh4bdtE7t+Bq8IpC+oS1jMS1IbwFiyQF1QI9aCu
d7PJc+RtPcN1XxVZ0fYGAa07mRK0RB3AgxSW23iYWNBOnNFMYlo4Ajgb3iwSvMET
ZiEH8ZWEvQ81jZkqDbtYeyv5oDY8v8nPZAW3kPsOiFp5M+y18zaUudLtmdVyndRY
sTfpPPIIXpR7Gu7kzWnDoGjZh6B9Bn/Os1dhjrUy5I9U2P7Fo60D6dwlhVwfPInC
4c8suuqfLluwZOV8CKsZV3rx9HgUDfdokkdyAFHya6cerB9VHkUUA4uAz0BIs4w0
PVF1sugcFFJYASVvqnDjKUkQpNId++4wf8nUqhHwZVLuahdk9cFQ7s8jpE+ZYZud
2xHVTnlSGvVGGO4K/5wfMw99z4lVBnhQDFb4e1kw9eM/Xu8mCnAZF+g2enBR9PKq
x0kJ/tPe8sFldABixNywnqklXkrBcqeal0bkxHVrB5+KS1HOwAXY0UASvuNxeMdM
MlcW/vgVK27p8mhAo2NejQNqzI9jC9v2WsJgViVkl6rp6oW/PEgHLnJnB15KsxIG
skIXjks0MrNxqho7ieULb6DUsbIW2FiAVVRLxWhPJxXF7eWhxBI0ZtN9v7EWtsab
1ykght+7ug4xvnpYIhVJC9Bo50ggUcpvJR+gpPZ6hf5Z5/kHdfOaQVedYKsROS1p
RhvnRjFXnEbDq3OTWgrrHDL6CFMkNf1l0+jLBKRX5YESZt6Jx/oWscvJtSJNmsnu
ts+/tQWk8UDMBcLE75xMDQTsmNROJNsvshuCKmq4uxZyfeuOZvb3x8tNN1PYDv1g
SNFaIF5sxMFtaatsasJoXsojwNpJ3X5R9X9ML3o94y++QoBZEIXayz4hZ2VQLaog
g+4E8KodCdvg7MFo4kOa5LP3z6OcWt9T1YuwdETsuzXz/xar4Ld8n+GjUqpy2h7+
DsDTzJrhXBJTk5HARvgAGm5MQ2ChIxe+KOwnoUFHTPx/nIJ1NP+qVqvwmg5iwg2H
Z0FjdX/BFZR4Y7VcU8WL1lsJSF2uHhm1X0YoiA0fyXZAycYp9wPm4PzdkDXGNyAY
JEpYJ+EYRxU+uH2zkqGG/P4L0IPvHEXriNxP4PMTqf6ArH6MnDpCxPLqh8Qfiu8Y
sqsQm/c+sZjkzJkWMan08BvZlV3GMTjQ+V1w4RtxgTyrjgJVJHTDZth+4Qju9qqa
atn/X0XgNYXb0IoMDCrv7BhZHNpqX2NZ7gquo/XRJZJQLZ8PZ0TvvXGn8m9EYenF
I8hMR1yqibqxHfpahgg5FPFdOwQyugN7msfCrwydqAHUVrejrjGGHLCMGJj/7s72
RQ6WnEZlfBE19jRV5bNbDu4FBXaWwf/1ROkQsIEDQvbQJIizkfJrWzCUX3mOrQXv
X5Yq36C/J50q9hH/C43mvAPeNn0IO8PLnsww16ku3I0Y7TU7yUHbUKwMX9Jzfa9X
TcW8F3QvaP69bTWWWheHu+9fIYINfaexQXTStoXkvCF6+muEIJ4BNOtIkLDCJATp
qF24dXyM0tb56LgdKn+5bmq+KBvMlriAdXLJglyLTPjbYsaHrmUGPdlWXl8OHSIg
skW6QXHK4M20G0bkVvvpeH8hlb7cevZtKrECoWMbmPFHahLpMDBNpYLbJEF3OeXT
ToLy5tigLL3UHTf5DZ2RNPDhigo8upImsWykYtY0AhsuvgklzIpJ549r/BARLK6I
TJqkNydRe3AQhki+a8Na6bg6+vWwRY3Y6mxu5kUIXAtvtsQbOwMP4Tn8mc8N1Lti
8gbUtn4CNK1RfbgN91BhClxngiwN50xiotKdgdcXsRIIc3ZH/jRIVv3WMg3udvFH
XZCPtucSNAqnLIeBOaNUmA9JVRlcdMjRPvc4qOGHAir/Vu/EFkVN45rdWVXX4zsE
9jZ0APQH23sntGUsek1++hoMGqiRrILhcXgZcbquXEX9w3N/HVZ5RD5/s4I2Ek4z
7X0wEifS5tjNiOYANk52+7hHqL+msBlL/3VsrMfbOqpkk6iD9ngMTCluOmGsO44g
F0fx2KJj3Te03NzVfHZuveP99nsWRsvqEywA/w2rrmIB5/eEe1PClpzwHOgCEc0+
rb/482TMSA1hGbHMcvc5X78W0/O4hhQQjg21BaSbIngiRRKC9AzAD8Z2KkStd3WS
q/DScTrJ5ryY+IgACuzC1fqS+KKNaYGZieH+ONHHMQDsGNjJMyb/THGbdINb1Mac
IRjx9tRP8BxRbRrl7YKkzaO+dRbYzBQESAdTT3BKfLHr+U15qppI0P3LbRpcvGGX
ONWXHQ7MG63S23yGvqNY1+kUoFOAygVJoQw4siFB1orfYhglVdQtbr8mpwieHkNo
Eny+oHk3KJTikBQpZCWo2bpMMG2hC3R1kv/lO/yezIX0fTGDd47QcR2+QUi3UM47
CyEn8eleHnfYfwWRGew0rm6u0omWrsYMN+me0kIoNW74s7QFpP1FGSadmHp/Oz9h
hBEe2pZXZ5NIA9IsvYzGZO70yQK2xuUQ6W/nOW8BkwxUUqqOdVSzPnNr8+XrNygF
uFBnsgdeGOWu0HRaEh6e7Ya9uYM3Vwoewc1dzqbBcy4xqXmgkPWDxVO+G6rSFB8P
pmtWdh11PObRzKXkqWldnzOcs9+jPi/rHZ1tKMEgGoPUM6spRfcbSXninrQ+gFAn
oJOQNAm7gMC/iauhjmHqUAaxZ/6EQ3Q10ExA1RGkV9TJ2eS1sKyz+vv51VToXcUR
Da4VCEFem3QRV5L2acfdFrgK/k+oql0s42WARvgwSi675MX5zeO0nJlM9Nman5Fw
Ml1lBMDlOlvt2hDAoNNETrANZVVRbGWeUHRkOHAhkupz0glWt0Tb7c4psOgBt3Ih
2/JbkitWnWbQTroqZDOjUGhW9aTblTGqi/ebFbSjvzdEJbF4nq4wwUn60R4kWmrP
IQshG8oHq/zVtPIBhv/qQzJQwPeI8+1Mf78OWuyfX4r8jT8RqOiL5BCEhhPfFgdh
HuP22MUA+nBpz4vJ+IumuhCtV8xHexgKBfoN25ldKh3K/2U4t23F9WdJ4tj8M0uc
bcXjMxrd02LHCxmc0B/GpJOOD4fH62ODygC1EvI/pHmBDQkZ3Dwp4UuVIucf+dpH
p4Ejw/X3d61IRbIVNkiHrCe7nyPToebR0dS9rkZc8Aw6iQ/0zfSn5pVbNtw/gpwf
M4Me0evC4g/7jiA9MiipwfX18VFktw4DZ9Y+8ASpYGXqdOOivzAPccUsuxIbX2Pj
JFQcazrpNlYvoHBCJQkkKW6gfE/lqvy9YdrQ1X0kxF2h5yEVNY63dlnb1wAWZ2rV
ZGENDCOkm59KV3Zak+woI8mwaFiIF3VzwZSka0klST82YV0S7SqqBl5D8KQhcjt0
CbR8T/kJmulqQzzzc3QWtx32VXEefYhx860Mmd8KUeB8bNqmW0y/sg1NN627l3vY
PX/xuOJYSIC0Lnf1WiXZW6Qoyj5UGV/Ko8JFsECnOe5tFH5wtLjbp1AnbSxx70zW
779MInir+hydaoodzxhgxDs512Fjj1taG8/+BKYPRQTNzJC2tghQUxB4C21mozOj
0Optp/c80d6h8c8oMVbWdSAlUT1gklNyNG1mXFKZJYH2mGPd/Z1kyAmfkNo/I83J
ZE/FHsU5AxGpr+5ldK/ryxSkYQyFBaTS6IFf/5ACe93Sgstme54x2g0JC9smKkzY
aNhnRyhnsEwq2iEpIttjZNf8HZwD1inR/LtXvtv9kGX7J1mwcrwJcPbdR3rDp+qv
gy9xyMslhgLB9Qa8esaNJym1iDmeXMuq/ojPq4QS3Jh4hOJbm6Z5MkS5pFkkbmyR
JrM/R6bhe+b8IJ9ov98GYXuPO4yGF27SmBPn+nGE1eV9pDgpvEF3izbVjyyTiSec
xUEBzuISgQD9VrQLWgo55V34DOi8wV1ZRXqn47OSGpDKf/YwXZ/4S2950GSgBDGo
Yva9oEtcuFHD3WkGOvZZKpn1aEKHhFV5PcRsDp+O4cnR22FlbuTQulyK2PEVNVYI
BghTEgmQj6MCjrvKI0pLFiqEXWLjGg6picEUbPz5nWNTmj6ui88QL9ZLkwERRCLW
HN0Ji1wF19Is89mwI+VQuR5yipTO6UqvPOy9jFY3PbglmTekOZ47vvzx2yvJgPRY
JUerbNwWUcNAMQrLezbxvW4LQYRawo0jujACVFO7PlkqdhdswHweBXcwA25doh52
KV23p+PusAk9uproz3DUYk99tmMXYQTjh1z6RMPBxu0v7BACVj4yFR+U7YzzOa65
bI2UNxyN+cwrNfFmP5QjBkzgQcV6yfYdgx3ZDUshgralkslQFra/Tw9w962dUmkM
+sew6JZHOsOeYqcQX1/dLVpS7O6uBzQVuK1+GL44HrlHjM/pXiSlXVzJGUeIUBo/
N29+kW5TedB5u674L/UzyJ/uNkA0zac7g9oV9f6GUiPN8zo+cKXu7+RRmi28iehQ
5MKIsR5r5URDeRS+GNtILZrHTSUsCZ9In4FN2yCQBB8kC45wy9F5BZFLU8k0JAKN
r20F3gvLLQsYkpuFju9Z10zMyfWkcpR3UbhpKlZbhZVTbF/OE8OpGa68572Jrk65
PjH5tS9TL5WCPflfhsP1UOg+DeCqKetB8p6z5Cnc0iLc81J5/MKvLZPdB/VToll1
cMnAYTX/BM7Y1mDEI6XeiS3W48t36Nz1eAbC3xd+P/jO/Thz2cSYeeELNmAvB+iH
fjsA9gUv6Dn2w5+oynzx5kxGvNUADe4V/UpUTMpQke/RcsgG+yNLDw780YJgSpWB
6Hgz6gjh+Xzg4nkph0Tsih8h16wHq8T9hoQgj2ePN0PhotuPpHd6rRpon9T/4NKO
BPtZnYASwRufCwLU8y6HcFRNaH19BA1Hdm76yiy5iit1sdqChUgHBnGOUkpOpDBc
/acF5AKx/K/RYbueTFTDXefnnAy8k6cutvaaXQIKhmdYtJf5oT0snRFq5yVbwSzK
kWr4IUYNHgmE5quLUb0iwtFk4gmTvyGm/+EsG9KXxykF0DPOddpzAGX7Fc7OXoyo
K+vVLbphuq20vicHEFsawk8Es1Ap0Dd8Aq3PJslVcERKmfOA7FufuWQR7tPRI/yz
gvhDAT79LCly5TfEeP454N+ryenh1qpUFXOLMBIk14FeyEG7OWmbfqJlQKyHvC5C
petHrkP2GmUyoFbBTWvKUtoze8S+ZmKgASfbw3MadUINh3rB2YXeI4gcd06KPuB3
JrcWXmreuXcaN0rR0jow2ugIw31CA/Ddj6X0ys0gkYjoWjzW7AUSLE1sVS7/hHXs
+WhUkqfQF4hgXg3jM/HzLWcG1ny5IkpwPlkL2be0XKtRtum9n3tkdbrpk4J+2lIR
DCLFT4Shc/KbX7P0hxit/+1/sxoiyCoOB7BAkeiZ2N7SNjOAdx6LE/8Hst1cW/pk
Cfhw0qPGSVNP7m5h2f+XCZay5xfXOPzS1u6kraNWB+s+QGFbIVqqWqvbfRudwPeu
aKVOtvil7/ICm3gd50ugKRn7Rlfzr2G4LN0edkhdmTiPkA3fpOKvKFGJXuggfsUC
U4SnxICmXNdfsOj+gHLDlHHp8wi/FyrRa3UAekTzzjiR40ZxhWFfCQOA5VSoReAu
qv6gALSgboKwMQeq1KI/dT+VHronqPs6KzwQMIP1YhGwQ2wfZjcKtZEdC4jNkbe7
vQRheoaj71lIpuc79nPNHIzmS3vhRFRb8M9lI/pVZTA2kYq0ozeCBKbiBptNkpB1
pcxl+mswORevEzxrG7jT1THtKHJ/E0Uig202VO+HD+g43l2Q+NCgvDPtODs1Wbbp
O+cYOw5dO3sp/+t6FDwe9xchLX7ka/7R6H0yZNIEI/jHlXW50x9p/Z1oWgjwwZHQ
Frm/hAa4703FH90rgx4Zr8ojkZtNRey11IaySo5zwghDIc3PnRvfaCAAnJ2mqEZI
csPo0SNm9H6SUCHaYyd9gEiOpMhKHpuOwfrrtz3iVFPYoba0iwLxOwqamIDDPCkT
UedzLByHLGb4T90Cmqa99XxUZY7R2Ntn9EYvgzjCCbzWnYMap9jXIooTyqRgaSAx
L8HXivPAr/o3+qFttPoyts1NhV/BYvRhn8B08eqJO0ea5s6iK664M4j9iuR+x34X
zURNVjdY5i+ZAvOpWzzrjJZnb/8ozSUiTJ733lZ9HXNVZt3qeQBuzWg4KJJABuRm
OTSrPQU5xwr2izmi/psDODxE/DF/HJs+rY0shhO1tO5dVqjybUKgF0nYpDG3VBdM
ITaolfn8A+CC6ztVGAy9Oc7Kkc5F/CtxrPuGnUm8lo3GzT5WYi6sC39r5iUyonRE
kj9jnaMqwpXsPcpM3BaUDwu2FzyrcZLTWyTWgygvDvt71DZiDZy9TuTk+dGRRBt7
8xX0vUjpFl0q3CHkTtrFKlaRw/GnzXoCSDcbWdvdjSxfUJE/M58NqZ3Ggpeg1kdK
OloRFkmQ+wlNT04zHrxmYX4Vk22goos/BvH0EptcmLW/eqKwP4PHwN8gM2C5luIm
oWVDefB1JkuV6EUV7hNZGK6O3yA5UFXk7BGDTV6ZkWlktar4GXtu8lK+zHQ/5tqg
rAyRBUa/HHgFLNy9NhlMXYHEmdaIXYmYg79VrUNPT7443wd5s6QIcJT7kUIWNgeG
BDQriFO11VdZMHbs+vHYRxNzWqWtt6mQ44GlVhuoLitWou4YNyNxUwlEx5lv3m5Y
gwwRoD3K4XfzQHnoRibdfqFDXew2yB21KEmQw6U1++xIUE5Y/m1xSIiDLFVapkWy
Jn8lLN/HrjjJB0eHg2jXK2loVsMKFhTVl0a3rHUlkBCD2vBmQnFstOBYSXAya1KQ
NqO9ynsIVp7mbiyIsZlUs/P8yxkFL72YOM89AGWboZUmXh0f7wX4wSl/vDY77Nt5
qi2ard6vKxox81sGSpxZDdpcxuD8ZKX8YTDl9l4fFJTuY6aEZL7MITEzrzhSdZZu
2zjUFpWdjIYZtVrNgz03KAtRnnyIKa66xeSrijXPO+9Nl4OV8fEA6PtTf1K2ygsz
oUF+COwb5o1vvepp69qjoubpSG9690/1xUzFPDG/szAV2JZOxLhl+iNRNNV4t9eb
/JzwW48qcUAnwtFBSft/0EuZvX4vqGvlmhNx8XMJ9Jjrg2OMhKXU9gRzCWpoRHqt
GwUDxCzKr0GjVb//QXryvMaUF8VympQWdkRBpxeqWmm9yKXSSaXP4Ozpi82kohqM
TogGSN4MMJXz87q+XL7KYNEDWZGV5akjqlOAeNdbzUuYjQ7FEdx9MKBr6MIAzdvJ
nTgK0YttrA/K/TIMb11lGICtYP0AOp5Fn+Vkuwv6SPQX7c3sEQpOWZa5AdL5UWjw
RDhlfEx6hR4rYsaFUCcohAxnRYevt+X7tSwcB4YWC2obvsHe1ZrOdmd3Qk1GV6Xt
BDOvD7YcHhyEEv1y/IjgCborRdwLSb9LtcTL63LrmMSc2CFyoBsaRbaIEWzF9zHE
z8zwkFTGIJJDrPACiVjCFpPc54ArHn7aw6lDc8g1yRE4ijy5IfpC5MMyA30c4Gpf
x3Yh5VHTKJjbM5SEeX08B6jsX/4JVC8GFfR06ZjOpj5bReA7lhZtinZubiC4t5Fn
dkaSiBac6a6OMtwBl8YNm9pcGq+MNHSDPcz+8pnvyMG7vqwSsKceD2ii9BUYYe8Z
OJhEoB3ZYb/RKFOnd0WdBycNuB/hjW4oG7YC5AuOo9lO7MIazOHLnN3hhr/OGwii
v2YU/IOv1LYAkwgc88d4ZpVVxdBtiCcaNBYk6+Xr+cExb5XJPZvF8UIlE81qTs5i
ePRogbWYKOYKld6qhRaJjrWMyoGSO8w9lIq+juxTBwCk9BjskPuCN8x5ZqK1YiIP
yK1tOPDrgntjtwaQnNfgtF9wjr11HDyminbZTCQaHOJj39e5xpvUKHExjb/8gsXD
3tCyYY99Lj1PKcadwWKVHhaQR9v+9O09Nsy94Q2hg7vgBPZvp0PUg8tTYoErIcSD
rAAw08l+kzvW557JHTGes/tYzlFBdzRRTuC/k+p649HXq0WVEx9XVjLRCnwuKSuv
SgOQCg/2Hx54iUD4kKQ/YpfTbKcycvKX50z1mGtFFtD3+ZEyZPMzuHuVvzHLvVE/
YVUDHUeWNBp5zNbRu1OD+d5UgyV15dvINf8K2PA0pw6sDdcixTn3njUvQrKrfMaA
c7qad7vpTKlFRRivjNB/0+BbdqEICvt1Q6UQCLMgkRtds5eUPV8xVRGPr4P70Umw
GdERua25Sv9huUsd+L5Kugvp1dhkbaypfiLJ0IZaV1GosRG9B/Rj51sR8NAVCSoJ
WRabT4YpmlEvELXL4EO8UTD1VteVe7JIG2vg9YifuQevySaAuiYkkgw0pP0bhNBS
j8uELDac0ijTyyBZq/qWxVhFixz+N24K6lRrW0RRcVK2uZsfS5JU8U6G8HcQu3LZ
DSTFKvtpOCW5m1ZgNbIDwpZ9OBWh4U+PBiXyQfiityMUBtieNLLCBa7phVlmoreg
78FNVsW3oVG6iigNQJOuQEgookMWmXC2AhmbV1mKIwbg8pd/WpFXJThM5/JmvBuN
WySJEGN4HBIURbb42anlXS2ZHVjasJ1VEKdh68U5PWGWB2EOKpxkiAzqXgzcBS+d
sWI+3R9juhv84CxYlsXB37teWNTKSHskWC1Rx+g666a59u8NNEg6GLVGdPms6vtr
Wz+wBE+uQL6TkCKa1ns7S6yLl5GJwDsrJgDNMoSDOSwLy6h42FVCB5yAPS5dYMo/
Ou08acOjfg6sllVBZUxlQZQCIdrj9v/Mnk6UU3vlnyTmnXnU6M8EXWAq8pxjhajs
h0KGLd2r4oEn6ooD2SZ8wKTphtzd6Ab02lQwdbryiZsapgubxoMcQScn2HrEkZvG
7Xx80c8vfDUdFH/V4EU21tWQLb5bIDbpgBaFYcyDbk6JbuG+kMfc+xlqINVdh1ss
BpqNo6k0XLaRnnvC74ePsoUScFn2obHdkfRW1vXUdWqdxwjpkN1Kfy2jfq4DaAKK
JazmEoQpVwjVQkxSDD+0LRV4FRGFouytGzFVm7oAjHn1gGdh1Jnrp/B1xSSVeybD
qXuu5WBN0WMmTwH9gvmXBPU4xBKCEq59wfke47c2vGmjdyUmJ+tpvIlQj6youLSh
ebN4g0sehlEM2nY4IgfnLEEDUPogOPD4upJ4eK8S6bmxjbagdv+iuq4K8U3Tgk4n
nZ5XN/qtWpTy53ooKtS5eyJa21hbyGfzI7WWthxvBrvgyDZkZfcaDDEM6S9R66HH
7mFWX1eV2rTlhH+iumwyJL9zIgxKz8tzP97MTXx2Y9KKLefM+HbA7FqySbFmvlIU
lCzeZGKSkMOxmtslEkj2d2IYdJL4F7y/3HJAbGJF1JCKRAuThnYWgP4j8ZNEyIBb
Ac1KmH5PpIX/15VKmZjTpE5j2YG+yRz10eTev3puFjIJV3YJUeifiWaz/tiaRbd0
S8HUDVDOkkg7PEBkuP2Ln7mc7YLkHJMeIDdMxItmlVNe7tb63+pE37FaBa+O0DIE
RiRYkhCFTKEObZEsqKtpl1++hyBnqvmY3QjpRqqX3eq3zciB8DbNL7YZVZ4lCFy5
zVpyB34AAEaaBSp7DWJlBNKtXlf6tbFNFDSjQ6zyxxf+AIFZq+ofzSdIZOddb0D2
IGYUpTuPpuXFoM9gFr3nsnoBnF0CGx8+gNt5roEUrnV5UWtNNbaiA6SjF67aBxop
aPwzeVx9gyE15toE2eMY3iqNzlI1WyFtNZRua7GP7HdEgdRSe8D94zSmtLoExdEJ
4LEQZP5UKeoLlPSChIPfedzYYcHQZCJeAEaCZ6SrU4Uhf6WvulhgF0qIvce6tC1k
t96N1nZbxF2CugR0xTHBZiMFBpowZ7EJVRn9qs2lANucNU5hvOpyFXUInpHCNna+
FYwlhG7T4hmE38VvIXfYxgN0edu2g56YsGdDKKyHJYNp4OLvidArGS3jADPJaHJX
Xc+57PiSOcjJHIAIP84zEpR46k8e4vtYEkNwS7gGrwUFBTIqfiudF5gT1GBgpEPe
YjpZ1OPq3tc1SG5QEITL0Uvma9ni/Acql1ZhAsFRen2/9EoIk9i+ZcfRI+OhsIKn
+swheSfCg4mYfxfKRgENY7r/JfGeuxZE4f338AdVD2gYU1A74Je+aB/GMnxfHEbe
+2hLpGjA8EG/n33Q4w5i59YJ+UnLPnJcF61ONdLwHqj3PnQ7r1R9MliaqW8AZRvO
hpsPGEyKu/xqfVbALxYhU7mRz+a6zE1WcRMVr0CmH9On8FFtiM7bB/JKrhySv/qj
PsGFJvSbEHD47C/sXAZYHTMDQcWKqmNzV1NcvqTduL251kV32lrLRR7eVKLpRIwk
8c5tRJ3HUxm/1DaOC71kYgOqe5pm2K3Ka0cl06un8tiJhslDKnTgMaoecpVCNmcO
STl2KKWZ5jPpYLTof0ZSQswN68EY39Nuz93csHptEDabxSsNY3EhYrWtBSbkZ6dq
5x34BzKGiPY/U0UiCsCueKNdy20dzbrIgZhU8gn3ryp0yS+van7khGj2Nt1HShAk
eM0yK0BxI2NZwbb70uUYWIotfYmvHb5q/FpPh7kc5OkVCngYcvgsVm6YqzFQ7ZrD
Zql9XS1wG0BcM++uwNb3Sisrz3L8Jxk60qH3/f5JD0INzk+VD8g9fTIDGNHQG+2+
/W46ub25RUAikWNT2CGrn2vt5vn1NdlZnj26sDwy9efgOgld95zlAE8qxSt0jHrj
2fgY4tXEnA7Fy/hjuAFr+yroUpHDddj3xj0e5ygl9ryugSzwD1tSUcwqUd3Ukb/d
F6dNpyxwty4mfXqEK9W05k0fw46WjhU8pIohS9lrHLn/WD4U5qQdLayqyd7k5W0h
QnmIZsJC+8eC3veHoTmEHZL75zY9C7CZeOkx1X7HxQHJKwagz0IqJbiY9kyWYQTO
P9ywaXazjYopLJ3Fe9L/e+IIgVb3WjkPq8+I6hbtANTE4WWG2sDxxKbmurjrBadd
s7G865Wm6Gzzh6jYW3o7KnqVNm/Jug0BjIQFIn/K+bD4DDH7IEHbnAbSlDzDKmIv
gjVX9hHKymLJBBLVWg09Hzm3S6/gn30wHDNG8nOsYQmozAptWPT/DXfZopoUHpDT
bNlCNvhXd+vKxV+Ll62SgHvngyCmRCoF/xSPUnpehSq7OzXv/BN6dU9kGX1Yr3d6
KlLRXSbRSofCNLll5AJamOHaSs1yGoOtkCwlITnafqRWCJc/uFZfx5hoNau7gWms
RYxJcwcAYCDOSZBWr0yb3GVYM9K+NQ0nkdtMCarsdG1ql6k6RnO2vrWXG2dzhrsq
exOX10xOROb8P/Al+9INZqpjZQAa0P9YpVrlhcx9C6AvgBdMQlecA7Kqel0YT9MP
IMJjWxHXzVdxMOrdplfDqEhIk8YO55DfEAG+wzO1Hx1NrrF3wvxBlhZEwWLdYNzv
aVP+oj5RoH9WAXvU/NfsXwW3dN/WgfuMcLnGVH2TCwrektokPTg2nNkTCAaW/KXY
57MIEvG5T3tAPGpMeIBe4gOi9+jIySdZS+CdnblfQDoA9Gd5XpC/iuBXGppf2ybi
w9qTrctLWwvqjHGjvOK4nmwQR1zOCnDShnjx4yFLb44AmOCwA2E4l7GjL2S0+FJ9
oJYlMQOOj1TOpN0iC6D+WfFamzhDYbDVMiQnjewAvgD97t7PM2TcVR0oWC90sgcK
G0L9P9sDXo2som7fCtnAGgpP+aoWuEg16wsC1DuXrzNmSMPFyAzI6DkVTUnHBoGu
NfzKtRHWlzm4XeJuMvR2YokJ489FEkiW075U0tUSCH81OdvrR8eK8z7jZdC6wdKh
44AZlTWkyBziSRGFs+wxhhyXU5p9MOa3+QppLO/qkjEbtet+zYR67zNdIBeKjjYN
QwUQJfy08MfQtmP0OW1P6zwC5vVxartupkRwMSU3biKh2CFarGGGzDlGMRDi3N+M
YzXELyhot9pD9WGO0W8UaqOHNLc0uxrG5ELP69qux6Whec/fYoZ/CIb3s1uiCKS0
D9hM80FwXE/WT+y6K5HLz0Wqg1X2U1rqArUcp4Ln4GvKumrIRKAbx81YXcGzPCjw
CXMm/tlcZ46suW0iyGwE/C+URKBRb5N2hoqmwFi358ALOzrXDuOoS0x2y+yFZnsX
jnOxJ8nzbbWde/p6NIL5O9eGYWj7MQ48vY1kMN0RIqWNriAfhURPw57vArycrA1o
wtIz7dDI+eYqRC5sVyBxlCbsZssbV+mSEbKOssIb/770suJAlLPYQ7bi7kJIDy+D
2wkdhn6r+OPOQ8jAguyAylKTlMNspZL+qYiE+TzqAEvmPWDFyzaC6EpXSiKgesSt
YOmmM0vbC6imcmZOY92e1x+Gz57waJ7tRviWtAnCP5Yri7u9qAM/9xKxBAuJcjGD
Hn6j43wwOEJC6gZ6SHFKCc1s+Q8u1/rmcbempOnmufk/o2MkA+8kq/AeJnpjjvTz
4cJwFbfln30QDMo0BGYRhHn+1tRVq1zD0JMqLJWVhP2iFNMUA5nlYdJmFQL5XL+F
tmdKhV258HJ7xFySryp/mTINX129g9klnMKG+V4xYmq4qtMMX6G1JHQarz9VfRig
Se/ItlnRVqLbVRRXgaT0+O1ldsD6zFY3GamQyOlB5nBPRcz14Nf8fjdkdPbLDEmY
huJYEAvJJHjdZdHq/ngnLK2MECQxNnx6mn7SQtmiNt6J2wkAcyCbgdUIvj2J5uGH
O6djVlKx2kal/WWb/DvIE0cZJOdTScwb8rgYrxyMRg1fCx99FJpN4kOqWFLqEfx+
3pv3hgkXqJZf5lS1497ecGZUY1JC8W9967DglQ+Cl7/HMAQzVQXo3Rs412kxm12o
oS16h2T53hqiG8Bjwq2TjG4rLLv/dP+MNTk7N4Xy1oA8dbVV1gVmVOlHS+pH0FRX
Kz3Htv8Efc0twxIyS9s659ifDCAacw0UrwcKZZYRE83YCH/HoUVXz4fgcESsk7R0
BmhGznYLeQpw6Yi6+XDpkaHPPMlmlWi34XtvPqfp/ydcwpajeSoGlkyVpG52SPrM
yPz/IDiSjSr9uBN9jBG14SOjVI+grRTxk/VQeyGh8sKFXx2lHS/KAz6SqwuysHPP
xYMGibDQnfxZ2J6FAPjnCEw0IMjDNVAJ6w48ZJ4nVpKREjqoPpM7Vdwa3CVzQhMe
74S+WJn0DZoRMlzvFiXKKabV2zEP6bxe0/JvburEJcSbW0A7sDcYXQB3J06CDUyI
CVuBQNiqA0z14bM0FT8KINODvOkX+lPYrLq3Utck0aGGFvIqx9h0oaJYNDY9LWu1
Vs3u+iGPmO2uk8RjIcAu1SfOEKd5REphf2lRZcfdd13lenHALCccrYpLwhXyHjGA
J4+S8ZitmFsuA7qzvMfGMg1bt41SYWYxWAWCINTtvh+FK3vRomGR/ij/nq8/WE9R
6gR56TVN1xWdmLiL2MhGmzyEtTV8kCEWIL5Ij84jYEZIWKFMPrOv+oHorFHwOsWM
0DY0NFavsG8sQDIJ0BURJRERuLH6syzxSylIkHW2tFhuFZ0LnzP+TlIQZX1C/DCy
0DHaSxJmu52AqXeOFatgNOfPw8ErVhbK+/7L/jP9kSfnSMivYn+EOUflVlQ3oZ+4
DzkmIT1hCGwYRwTTD5vIpvpCZzlTX8RTEK6DxJdBmaQ/IjY2qu0Ptrk/0CBr1Yts
0YFySUWst0wq6JY5t5+4Etv0V0PdXMNYZFNV7Sj+jDDNSY6HmyjEAlcY/QzflAUo
32Dhs6H8JEkW2+HsEQxxFHVI/bxGiuGvxAFBh/bWf5BehkLcRoYVW81VFRJyvmau
/bK2sTbm/QaRxN/uRIW9jlX7I6sQzRKi717D0pZOMQf8Uz/R5vz4gc9nXAK6BGhp
oVq9S8f7qnIFRA/wFbBEozWiVdOaDkvx/7s8KnsIZIbcLeq0aYJWecp/Hj8uBdUl
xhYaMmA5fe243nEcx7ceSLmjamCJkU/GPAIXXN/+iJVgmE+X6Ve0vwczQJzmjeGk
4MOeXOLKFd5anJnI+9QKwkic/gFg0il7uPRoNoy1eCNs15F9eA+9xcHs8tB0Jt2K
SPY4HLxglzMTUAZspMR1VKQITNXP/wEJ7XiGi7I6UaWBVYbxQXRJtISKnF2VxSHc
EVNqj8Mstqp+e+Gz7o2zgeT/dVxhaRFqw8UF7OFRwuSuH1VrLV/rkW77uypNGfu+
9X0ePIUF5ickhe6PAOqZT70/JPMLN4fG0D6OStyAwiAaIlTIDLJcj+v1PWPUkEtQ
Q9B1vAYyelh762xsr5UKiWt45WsO6VVNsva1wkpplt+VhjqIi0HBP3Hz5EqpYbn4
FAo6uTKWbZ6vA4b/BL1lhxQtHSA9C/6Ge4E7K/Ekdw4YcFGDI3RPmd0xzwaw7dld
dA14il8F4gPrkMSbINy961G8277+I3IyYAR4quc+NyiL77QNiClj6mtzuolJfhcV
11ReQHHl2FbOc7SmM5ukgnfUfoRl2GuCbZAaIEfto+LY5pctgpq3wNT4yYAl+fla
PJ+GgZ5PXK09k4YKRZiiUGpozNksgapvmaqnXVh56bxbhjVBUEGM0p2L1loxp50U
MMxK593KdgfTh5HImiF6aK7DAnjWA6saOLtRrGbME28bhCU8O8x8vE3CAU+Bggtn
3FaX19k+Jd9Gqawe+MmZ4H0i8HMmxN8xS/I6N07luB14iIWG7ovcLLA3PmS6hY8s
XoErz3WsFCkuAE470xFYjBjVJ82t+TFt0WD7RDo94LvyENVrZFsfL3PYmZ4nL1JI
lh6kYRgxHwvRQitDVTNbbVDB7h/rOLKAVa9cLRL/dBGmur4DOeTRrGS4mMjqsgMb
0alb/tIQdt/+aCu008KhNQEG5z1qKOQhSXp+XXijUNT52Yn/zzGRc8eiPLAwN6yw
Ov5nUC4dKWfmQlZlFkX7X9uMA0/bJYFmzsrwj2+xmY1/e88r1mrN6AhFEZTPBvS+
Wr5tlDoGKB8e+86qmkZ+5NZpxRijUT3SFcGW+ETYz++3pmO2Cq4U2hXp3ZjPEmmL
d7UY7YfmCNZVZxYbj0Cy9PEGesLW1vjUc6u9vdo5UaL2EutuvlNMeQgAV6/5I9rP
lFmh5wkpXyBvvYDcv+iTqVBiEZUAvGqaKikWno/NBBtTkrjv6bKbFSeAtaLQgbT+
VhFBa53zMueDD32+7RaBxs4MTgsSQIxXxAwiaa371EOr+gXi2wOvwiHMAAC5qDQ+
uXz+P5r8CDZeCJJ6V84GwjNwwEwHAMp+wQG2BXEc5LGsIhZOiGztG5/qpyBLU+oY
IkEG4aYIpOSW66/I46UWU2WToapt65T8lpmkLnw26d8A16kLuQlRg9hrGiH5tLzJ
Wl0JS+Gjnc13Jc/D9+5hKkRNy6zzoVIQgsM2hBtfZxoolIjq6W7Oc3tY1rEpwU40
g1DdhvMWwJcGohqPG6y8F9wep9PN/C/Z2nuTflMmGCdPHr4ReasSNFMwuuA5DxEu
WTZKYbjNbGFusllEV2dS3iMVgZ51ohnIDCChCpM7onKvEWxFCXqXcoxWYoZCErwM
Ys/eHAsKPvZ5ZPZGkrNq8Pwj3IRBZOp3b6+WNH1u917rLvIh+iq0xEjRn2K380hW
iNXtpxdOvLRwm5untJcaGmP1XcdBiuK9rxYSTcp3jDNq1D+AMph71nmZmSkFx8l6
xOeKRHCJU6gB4Zs1aetenJZ1GGylvxKyViRoRIFkJUG6hXNAPHDAYbIB4vAJslzf
efB/Fl9dmI9NA2jEUsTxrZ7MUtavx3cU8tWfNH2hHaYjgpMCVjv3lBIo1PZmiLmo
UoD2njgQ+pQcH/sXAbpdLCqgstVb3TAgP3EQfcfIgMqOuZglm1ygzt9KXwqo1DbE
UphwZv1jqUJSrck3svPQhgcgOLyhU4bFT4/2gpjTIqYrbwnIl45S+FuG3+v0fbsm
GTdohmJUQGeeeDO0Ny0dqHjbXm3CCLTCcEeKDI7LI+UgczwFZRPnhG/Q0Y9yLu1j
+fxCeC7rXV0XV+jmFB3TBkbcfAfuogaz4/xsC8zFqfgZQU/zp0CiAeq7853YGXzg
dyVvr4yB6E5uevkjux9BeQvQryXK8bwPVDl1ec4g4iZSRs/snu45PFdJWJc8uKjM
QTW+ZYbUEDEzpoip0CN2pEwRdNjLc0huvpGVpPxP3DMzTB35wpUxazZnm68IXRZv
WWWDs3WiCZmK5QJhnbMh4X3ZOWVE1etyiUUYwcyjKXCW/MUZCMU6CNZ95ubu+B9y
vuGxXIc542pas70cQYUxvMgLVqJc2zk8BDAyZQoD5Gu0tSCl/LGEkBXUh9H94VBj
/YJwa8Yiax2zR9LOVw65ZG07Q9dhZEttH+pefxHmJiSIKQersbs6dGPyn9T7oR6C
cgPuPmIGmjbsQJt/O0/7J1CXh7M5rwgLemYOIgD8+O8=
`protect END_PROTECTED
