`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1xKSz/cU5z80xv4fPcmcrKKA684UOuLBsfNjjjG1P7bsY/WF+vGjT2dpdcNyX/Uz
2MheATKP9WArRRfAq7M+IlDyxw1el6bm3BGcG+ZrioRNqr3pff8YXfzFLaRbmJkP
OUXAMWCPhGuWeZHHpT4IFP/AlaPAP/VkJPbnFhzG8vTdwZzvrUZYjPmg12ZlC+/4
EaIcj1Ogh/SDxOtVucsdcW6THziAseCXEqRepA81IUk9gJGtNrH5bmW4LFwpNevH
5Uj7K0ufTwbcEpyC3EL2SvtX61Avnh9NH3HVgyGD8mn7XUkb2bX1lyAMqEVlwXDY
OZQ6wRZGt6gOylfCF+gWCsGiklAbiI7P+AABN+N4aWWudUFU0F1JvvhSU4pPjAYK
Me2yH8StgBrImUJa183Bp7qOnwJ2u9im06sPtjbtB28=
`protect END_PROTECTED
