`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nTTFuOVBUoLbbQ1kFa9zkogVJs4al0FbHNkWYlon0H98VxdaO2DANO8aMgfABHv2
UTiPqInnLJHXrz2i1+4yBiXrhqMZk57oD7oP+6qzetmW7XzDmQuUft2MBShqwiE6
Bvhks/i5Z3XuujYzVNL5zoObOmni8D5VxJuZ0Vn57fNdgnH9YLEexkQz/QTYqztg
SibtSooDS8XZ+bp7jIhDU4U4sAtkXSj/YDMaRDkgEZhn9DdNEkOUtJRuDlztqkEY
rrikRotldIr5IOpNC4uarv6JVlEMCkCqYz7efMu2/CvcMVnh5dYP9FIe2MI/f1QE
ktguPGBlAbcY9WwEjp8JI/jlfhQhhshKktzMHAd8cH/4T0mS1IXKYfkxBePgW3w+
9YHS/hiEX/mI38hl2qsCMyPpjnnWIFsRNUV2uq+FodzHj7Gu2d1ouTaiKxN5I5Mn
ZEwXOz+hyXTbQJRauSl/yDK2VHTUk4YqGgcguFeC9yGkdus2h3RMGPmzTH8ini3S
jECLVF1b3XuXhdL4g6EBFUF8a1NUPoJAIYNE4eiaKG8VZGFIaM7hcbrsfZfYzuEB
tRWU82U2t/AqDsk2znJ5qz2I0cezjLp75r5M6ruvVih3fsimWib9ovuVxzvNQ9gZ
Gmx8zS1pFPO94WxzNPuP/HTRcZ7P661xmwGm9ezSKT7eVr0Ui8fpHtXTj5mssRGM
ITOiSD+vXDyeDvi2MsffvrpF9wdE2q+T3zBrdDQgzm2Gp9m/tpEgLM32rwX1DAv2
YOyoVxyijeYuz6/6k9Ds90UR8kP6DR0p8hx6LMORrxfbPumB2UmftQ4dO/asqzn1
2OmK6DMRrX7fNIDPgqbOtu2FdYv0tw81Hn3/zCD+8nfx1gLz99hkMxXMXbgNy0HY
Zdap2RBqaRaBagN/qgfcyaLFYONbG78nXVQwUR+0LF1HaemstzrWM74Yxbe00mnD
Ffc6zdXRgGvYvduIxT+Kmq//6VPX1iF+X1/M415jYbZU/zEOj6CyCZRtrCeLYluL
jl1XaIH4MX4Vy5/QHMPhqY6rA9MrqExmwbKzwWFHJoC6C0pgyPRyiEvB3YDg85Hg
sOJHjT7to8XcT/MEUG0lAyEg1o5XXKsg9aMnVG3+mkUCHLB1N3/c8l7CiRLUvaKs
`protect END_PROTECTED
