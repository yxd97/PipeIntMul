`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1/MkCeFCnhWl2yF/ImdbEl4wY7yh+GWYtOwVqP3dRiTqUXloyk3rPJaEqnk3jDX
Hf8suwsiWv2hjKGNmmdEPd+oTzjnB8BRbWp0TuAwHGiIK1h0ldanO6TE5Y+rr6FQ
omdkm7aJQVQdZqk5LlRsDDbpw0V9xn+8pTz2qxTXT7qq6FNT6mgrCZ5a/B6751wG
vSnMNHGxgNOpJBw1OhCVTUYFnoBVR4OTF4HjAPBxdSJ75fQIriuZD3vQ9giwifpp
NEDToqu2ZlgIOGFPOkrgNQHlSvzFBotF/jRa96gLbDuwruDgDwdxVvuGgsQDeUjp
K0AIE4CmYXYwNdBDiv3oRzUfuVE/MDwnc3hOJ/heCZMB4w2iGff/0My6gzv0mP0u
ZDmlYi0KchLFxi2y2sX5bg9jM7FYbNlo8XMGI9H8JhDOiE5v3T0gMqulS5MZpDeC
J0/tS+jcMr+JcXwvqkklFyVzKWxjdfhjZSxHz+hgMoDihpITUNbo1+1EGouXMsux
wuuWlNaEXjuCs3f6Nq+gzaPiQHHZDJhKSVDxcnbDxX7GSCAfw5COxuw0X2CTJbI3
pn9Cd1g4OTSyXVMxDif3mNEFJMWuWwh4yBkUmwnai6be8eyY9jQ+SQXDePqvvEX8
ktKh8kfMhUsmWaVMrp2rtntuKCBmZhJ35yLGt/xJU/LW828Z3EmAxbt61dihvNQd
PFcCLLUUr8TxQEAXO8CMt30XSGI0IzD6vSuitCNV6Fph272IdNbTCnZPTQRSvNoB
nX2I2BtddW0g4PiuAqTJmuc8cRWDSh0QCM/2GXLevB4vk2+GUPR9XggQk8C0uFew
lFT9pGfU6ili5+wYJIqQg0mpLHDS3qR8A5B9ESqKKHsrJjMTFCeEewA7uSsz5RgJ
Xrq4lxzjnCpjw7ADBXHtWwajXlAOR+HmQm2vWxDW7o5Yu8wFHuVmIyK3/yure8vx
nguHggfGDYwntocV9OG+RzlpBcdwnlZbrAsOXUOlimswpGlYxpJ2Abcs1QiuGGvh
sKBbcE/n6tt4bvNW71vb0h1LRQMZ/qfEGz2XE+6idSRvJX4sMzCYZ53vwLGvnOPh
0obs7RjlgQldV7gV2ICbgEm/+i+ZIjTbi55QbyLO/uEsi9/xyA4SiqYMAHnKdj8U
Z+p86U6DuBbjGfS6ReNfB8pQB63e5I0PEmXXsDqL/qD9GylhIkNy6IUA+M8ep5FA
YhK72D9H56/Jm1lrPpoF14e79vuIGDJdHNtpX4yCjFeUTIi0PtkIjI7fDXQhIprx
80fprcTy1HLk4UAUvz6HC+Ox0kOo4bkrhkIrMMvajp8l8XrmWZOiVYwHOEm88+j8
iw2333WA33BQ2AjMboHnlmPPZ5IfwQkdPCPm7cN7e/CGdJM9jvI3muK3881cXHL+
WPc/TeKsZD0fTOOQijfc4Z7vlY+6Mb+YLhsdNaxVoUbhR/PsO4/IccLYgMOPYaAG
nTJrVjt+niZKVrmQkCP/Mkf65RU0mYnEF+8aTYbp7pk50lqKIf3oU/Ld2UdfEH4v
egHO2evUhBqaBgy9o6d7Q4d/eX7dNJ0KSsGXQ06gQQug8+QSaMXtiA7YXHrzs5sw
mKFi78qex+0Y++D0/EofcQtsx8lfdxgl2cFcdeJ1GV28reLs9d0Qtk6QNe9Yo57z
zJObfpinEFls1mTDZsjFaW2ZKJumFg1npyLgPebs6mHxDvU8O6d2cjopcEB+RziX
5Ha8UMEltPgHDirg4bDp+YbLvUBFd9T5T14RMD0alxd8pKcnx9/L/Gp9n9HWCYhJ
7ErPNObNoKcHwvYtnPZ1E7SzupLNX0CYqY9BkGOrAzkLWlKfQuNXGlKtQV/BFrmT
DZVJdR82GVLNYLEvflsw1wCE7JEEoLGxEMqjqmwRip1m9gajwWdhwAVG9ELStbU8
LZw6nCDoSDoe5+BMbnmNuUPDqS8nLEeYQM2SX4oa45kMi+spk65bHatKg1OXy2mG
6qFlcnd2F8LFThODfVPis/VGR+4tfP6eRG0Ib0TsqHrNYaQ4ie/EFjcMKGuoK7K6
btpSh9onQm4IPt7O4GyezAAkVQNDHDiQDfn+3iNG+suKp1HMZsZjREFlBC6IcPJy
ykCBPdJ0n/FayQYx1R9r5dg4UndVFTpL6/bhOn/2qEMOzNceEwyno0g9DKm1UUTZ
CxSF7c+vulfUC3kFdAFC8OyNtOT8yzMJrsHcksXECbWKGik1C12cpVIxcgsye4/p
aX2msFu2Zodpxnj9rSf9sA==
`protect END_PROTECTED
