`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TNxj+hppFVMFYsVoS7Qk3Lduxcu6MiNjiw5Lk2QcXG3YxCJUg/g+qUNQhSNw4YEF
R2ukNv7U09/JQBT5h+nIi+sUySqspkS/A0BFjpWYulhqOs8Q4A8B29cgPfgpS/mw
olIPGl2ZIcOFioJRqwxpgUs7G9qVZ6N0n/AW6RWiAADZ1uElph8yxrCVgaSj6KUV
nVKwP91GeohtXJBptvYMy5/oLHmX8jusnYlSqhhF7NRzFrcd+58XyUeKoHeWjQwH
KX4zjF+f1Ah+fGrn6RNYhyPq/uZ3QpQ/o02YXHtYYIXq6ueYDyjLwLib71IMHGNJ
+pdHZGSwC8YBGltYomizyNDDXbEzS/9bGag9Zej9ZNU4aaEZEWrE+4+qzIle5wHu
bEYW6p03kcbImK76vgd9zVu2baTX/gc7E8Z2HT3F8zY=
`protect END_PROTECTED
