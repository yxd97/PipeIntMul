`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgmPn8O5omJYnOtJM6QffoILHVAbS76oyCQzEfs2wOHETpr7e2tdUbmwEPKto8Gv
cQfjwF0YkowjhWAzWGMDRL7FvnkLq3nKTg030sfcoNs+bORnc8iqHGeCqXFTffuj
s4Tvxb3+TvU8nyJwxSMdX5GKYZLp+lZYlB/MuPTDfzbSSWuS68dttaUs6TZLZneo
9xdvo0gNyKFP2eHbl8Z329X8vlBMPW1aKmzaI3awABsnMUkyKcBjkYThoCGf0b9n
+DKPi7LlweKqxIwQvoJ9ezobH/3p6zVyOpXoESkvPCpqQCk28Cd0eTYvH1f1buS8
MxFZUWfNgmrFckMGo8UJb9Zs8oVj9dPKjqF+T1NkAO6b+HpXR2hILp6a+nINKpkm
8Zj5cp1t4d+GQ2aJzOyLZJtttoflqFS5ImnxoxU4k04tFRKerVvzJQklHwiqjnhb
+1abmJailVGfmLRkC+leV4/GATXBzovkYeHhD4qPUZRwu8UpZPs4JIACFIf/53Xs
B22eXxWtl3B+g3Ht3gsLWR1URltfeSFEtdkIIrUVtIwi3wtqAwuNu/+dptygr7ks
q0rzwpCl8mqyIYtmgBzgnNhOuj/vEAi+zrsE4e3LEvBInakLrWjKtw7QuWyrNJYE
n6QVWRVnv3arz7mezGfVeGG3sJcPxzJvlBzXc9i4l6R3gzz+EoZuHZwneF3MkBQA
riB35eusyvWwZrh5q6r7KBk5tpIpsApALhZQLlDDSXiakgx0t/aiown31IXSKlM7
dV5U/6m9ApdMRQNLC8JaezDUk+F6PuPwdsfaettvNSXTHt6QIN2w8SbDQEu7lhT/
khpuiciOdPji8eR0IDcvHvRh9T/ia9PfDwRnZtInsoHvspFdEWlNvlOuIzZvPL9g
Tqdw9biOY1Slpff0892qwMgUbYb4fLNK8MFjeJMPqXhIwcjELYQ5iexrIwmj98oL
2bGz6+cYQzWzg8gkjaEQJzMrXGeDBU3x2FNFxkSqUPkOR02YTG9Jn3XkHa19+gB4
ccmffcXsXiG7NswHjE5lFDViUm3dazxHt027/wKCvt5UaqN/i1HF0qnKAI3hj+Er
EjaX33F1Qdv2p7bvO45rzd2bZAn72DSD05x1e1+knihJJqcXve/YPBINnmjJqrsa
EN09dbawVjQTUBYq5nsFw0btN6wq/GZcVXy4lkStkM70c8dSRZBN47SHrQgIRoAp
BTvNi4N6P4Oe8wX5a/d7Joz12YuU1Duh7THE7sn/WdWs+VZLgiTIHZDz4Tkj7eUd
sSh9Q5bSOnRd/i7pLy7Sie63nUfaksifXXbdAby8kbA5fEjefiQXtd57yRF2ndmY
JDfjaXzM22lsjSAd4aXHJ0MSzLjRecsXpV6pk0cM4+c=
`protect END_PROTECTED
