`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/lN1U1U5yHMvVlRr4W8m+l5BOT18p+Liu+5lXmYXbjl2nvrEoKBrWSunrOlMbnY
Pet7ShqYEFDr+CrEHCKnEmDkxCR3+dKeDcnAXARgaJDeAhfREdDxtPH8pL8BV0ps
a467rxk6VsYiixRsDKPP++N6zqPkz087oE8lghJAwOzgy7mXRvFO2weY7iIP7W4s
M32l6YOyjwVUbTRyIgSfImgVMB9NMFrSg4p5PnewGXzmHxmcNIW3+nBiU1wZUA40
RcMR8GHsVrgU1oIZNFEvU8e6fPRYPw8+USd80nccwnCz4ETBQthRtCwzTUgwXXgZ
Si0Fn8V+IipoWhmW6HzW0wYEYtLVjNmdHeT2jfjM/9JxKOsqX9Dm0UyihLclrZBg
37BcEoX7W75PTHlHz5XkWjuNaQT5oOfYiGFBQrw4jkz39RBcZpv+KCTcNmRlyVgP
1k5PVxcV+nwYCy0E4kIHIyhe2HkMWwn9AfphRufYeIZu+cypL5q/K+tHKCrVgjNY
AHSRpz+x1XU9ABvaa5UKvLXHu1YqeY/ecJ5x+MWwFIWPGOOC4opNsYXZKQ9hqWt1
A4UlAbCY/uM/waE+lg12bbW1FlMAbh/T/2svpST0K/dDBwPYYbp14H1BvMefgYCG
0or0N6rSlzuATLy3W9FB9Sd3X+KhvJo1e2muObewObtDBBPRfCYgfQ2qK/9HavnI
WUQ33+CETuTetqup36ycWAje65im5aZL4/QN13T+t84bWzMZuudbRLzBLO3JiDtI
BgzmaL9Lu/K00I4ziHiRf+kbOwVfJlShZcccMc8Vkhs6W+2vLnYIwQ4m57OlGXyD
nKs46ryuRv4NGjgiCUkBdfXHIcNzlaoTf/qU+V0J0tbhhASs10gGAr1cV2QGGnHF
MkcUo5enjIjSJNYxmbuOHvqX9LfshqPybfmu2mnj8Sx1s/1lx8H4780z/Ywx7Q/+
jlQWYGNxphKeL80d5VbirJILnqdtbmko8P5FdqVr42WrgbnEbg36+Y4FvVbfkPEn
DNitUF0B8TgOmIZ/JPRqkS2CrB4pqtdCDaQJG2uM+vEQ0pC5+f9iLYlpFtYwDZxv
wmwBw7k5LfEjoR85F1ypo0UOxGE7K4YmbnUKB23b+1B+Mv32UHkIh2XL0LeL7t8U
2StR3UM6XL2INdN7vkkFWkFFchuoUejvElNbiff3W7Wlm6Rnajx9wtBOsE6Yk1q7
Mbtclm5d1ypeypNuH7T7HpmJCO5cNsAxmL8ccqTMLoI21REiKY9MXsIbGXUwj/yQ
Hm/0NI/KHUq/RHz0LBBnuj4b5k7fn5Cuou4pDkBfTIKU01rfEAJoUqeVdDsCKB6S
J/V67B9s00Dre1/4IiTLLwHtp72XF/gpbDF2SaJZ3+gHr59LfWmXV+0WvOkNHF/z
07vDhcG/RIirXscEp6Gy6o258St1Fu2a+jbyAsz/4cASpzxhc91ukYrPAphTi6o9
ZKl4D2vGqzBlrimRykIdCZ29oyKbaC9BHAA1eQfpX9onXB6jmkfZLLZzlnlJBrw7
de+zQx0jq4occdEfdsp2deZjE47Kp3LuFpdPYc9oxlOh2swdvMvgXdNxP9q8aU9N
dgWS4GHjDqNSJadmb8ytfDnDsO0+y3jAuIN2BcO1JLp1T3U6Kd8vR4zzzhZ4yVyF
ijQACI5QCBQ45MRptDtkx9J2PJINUv8IZb7SyDGoUt29+7e7ihEKfi82JRdTPKUM
EFDKveL95tYt18ToBuF44gmKdaDRT3jWgmQOYl9pOUACpurexv9tE+wp6lOIb8Br
`protect END_PROTECTED
