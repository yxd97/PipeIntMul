`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTsUbnBzxGD5Mr6d2kQ5KoexZxt7qMdHQiIa6nWP3MB24QtXpB86O1826VubmWlO
zyqM1qv4LM4xaNlS2ejoWh1yot+OqF+HQ+/BMxVZwWrs+g2oGuZcoB/CWi2q7rOl
m9k72xDvTX4pQSL68aR4aWEUXJV9ZBn6hUXBNtS9iu8bfaol1zsJN4TMgIFA1MEQ
48zSV1N/sfxtBzU89zpoOsTjL/FRYmTF8mgA420l0dfLCzqd26sbngkv8wWRLkPm
ARpsPRZ6VwHAQ0BrzmQZ86WE+94NNRxzAYMaLCaNmR9Yg5FYHCSVoag7v+e0Z4LT
cbzqL8ebM4GaiVxYHCav0SEbF5EEOYMo5p4XfMBlBr+a3Fs1ck+bwYO8tVRTh1IY
u/EBgDMLUuxBP2+PmU2Is+d/ngGfyjbkkQj+qMTCq8Q=
`protect END_PROTECTED
