`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NbifdpBYX8cIIC3XXL0ymab+6oazg81QdsUanxgMV+bPlPO1e4pnahc/qXvS9ijU
nCqGoP0TVtw5z0WHEFP9ArYUyDb68m4K54JnKV0wDHxnqImUWK4kwQYgt0aEzoAj
9WqXUKf8yISJQyUTBkuUkTQi6bw/rWoTFlw8pdr8Ti28u0/X4VnPmU2xSipyo2rW
GVdlde/TUwfavNCRpWDVwO9YrqmTf39+WwWLmD48+zi1bdt3w8msuYP8aH7gdNp/
IbUWs7rsA2aAzjfuLraQEAqq6pws6u7q1EPdPHDe7gOkIsz9NK6/VA4IViSt3jUa
5upx0eCVKA9VDaERpU7Oaq5/XH5YWKXW8Pxj82wTJ9YudiJY5PxQhO9LrXjTc9DH
56QAJ0UlWAdWjU5VwkD8W0111c9B+8MDT+2OV3QGJ0NCxi8k5brpR1dJtzS3XMml
5lknmmsT9koOBs8tNAvGipuOSvnDRqCazdbe+QnNsMhiiVnNiXIv/MEsMeFl+oBG
ED0Y5yaUBpZaz9nJRXiBMfZwpN9Dmd9GZpTfzizIJJMun040WLRCscEd1nyneM0R
n1kevEhTkPYwKuZqXYo1ZATExNCosEBRfxwCSeiLuU1NFFEO6JEaraNIVwcs0TeN
RaM35cR2/y0wEWmQMrGNtf8SuiEyQoxv7a8g03ww6JO9rXi/32MC/zzFNN3KYlV8
cCRWvYBSZROt+ARW91ugR6MEKh0/7hchgI+evcdGCqVSaG3UwSPhBTKG+GhyWmJ7
OA/xxKiHnweli1D48GlcSXI05Bf1mVBIBJRJlSJ6NpoCEcTW4Q0ZQUxV5/yq6jdu
iFVmP/T1nSk8DPk/OunyO8IUCdeaBaftqHapGFKM+AGEoc2lAPEfhNxjat0klfO6
bkEeRVYr/bWEvGDy20z0vZW/o0a7oc43PG9QZFoXkpxF8kpNX2P65jWrHGD/SJPs
4FkvFj4Pl7E3O+Sse3YkKeB/rKqCn447yyyZeUHETjZK6AcewImP426dftKraQl1
B/uECPJD34uFX/WwiZlVaqJIBzzdqELdWo4wAYCcI5IA7YbDNiSnCOVNYGaULpMJ
1s1Ayn1xmo+jVBP62chT5BVS2d/UBLAr9InTqxjadDARpaeHlfZCrSILZx84P97o
BDTs8n3MUJFl8KmZtYbZ2J1heHYq2oaBUlnGg5e5+0uq9uGRijY3whLsreTyscOD
O7lR1QTV8/dTzvQCA4AHQzk8y1dOiafG+SNGKXIRh/Z0Dada41OVUDceScee1lFq
LUaRKjRV+qsGhwlDUQiM4yL/fKMREfyIaH0RnC1zBgtj4KOJ7ajmj4HlDTEFPNcL
GdCbwNIWcuDt2CFTQRHhvMCXA/q/U0XZXZh5Iz2hWkM1gVMX0tNSUqpeHUHe2iHU
8jwxqTG2Fg+hNnMDSw698YjgEZzB+EzQYv6X8O139Pk4ulTHB4qR5SHRRTzK7bw2
DklLdR8Ji50mLVrJNdLY9qm/I/+/JBZuq2VnS4E284z3vyhHGbzI2u5EM0BL4HCA
WUufaOpWA05X9c1doMqpxPH5ccEG9oeut2FkXUDTbNfpSn6tsmJCJ93cz+eq1LRx
PQCGZjHshrj6EJq+k7hihp6THyrgtV8WVxF5V7ix4gEvPjORqPOepWyCXhdY0GHD
9TlH7rXE5CBpAh2Op8zQzlesj+73yDgWHmKCPKRKp5QDoy12M/fft8RIbZy8qFPt
19dETCO93JcopXg94QE3stlXB2DuYnK4r4mrSzjjfy56g++94JH0bw4CNamXRIRE
3BG7loh28uIURtzgF9hettNzdnzRm95kTFapU8DYSeG5U0vtkUN7WXGDuESQfv6u
cdIA02xy0VDOOsFvgJVi3xL9YSd8m8BfwIMLoe5unCa0tGMZ1welPYjAvtmFbd+f
yuYlqg6Taawcs418Cwoa1Cx9iLRFcaAQDAXotNQ7DGw5Hp4tUe5IFGMHg7AgAKAr
fJWWYkY23V7jEGz6Hvq/0s8K7d4O2YFwX1ZQyA+XgGNZ24g4X8K0Lt/M3K28Umam
Am7dVW018pthek5vYDgrGo2yiKjiVKAMqRBxqbocf2ksV/QzknqFOrDavb1JIhMr
CJJt+Dig0wA9Zd/gbZPCPNqXEExd8nRz5UWd5UT5e4LwCvpNpYZ6eJioITtUWrAW
UTzpw8h5khMNbLwlHKyEzADj3eCBSxKfeLNbaaHjwjpKzB/3m1ZX9EqOJNzWV8HD
nbZpDrAMdjbwEAYp7qRblAoT6c4wr1KYLa/okvZlE2zjDRBWQsj9tUemlFSbaXLa
23WrSPYcKFZ1K6QS6Wp7xoNc4yN7O0baUbh1pkXDvuKSNTQpgJbY/BjrMCljGz+B
P88npbkO/OjmtdTojN7zn2Ss4iFmGdS0d0MJ13XWt5ki7XULQj827EtD8M+K2Jsu
/Fu7gA4AIPThY7f7L0ecp+OC/DzKeOPhvXFjiWzx8gdvnCMLu7zkfW3OrYZwzpAB
hFflhA0amAqmVOYOtlTMvGXPII99KYquKwk5ZkT1fqTg83HBNzCrMrq7W3Wev5pb
Tqsafln1VJBz4YIYcq85gyg96NLX/P8McEjJ7fqOcVEU2AJgALMlrm1k2axY9XhV
9l8Rxb/5tcSF6Bel2EZ3pBV36GIh6nO5OSVlfBvNafw7vJWQZWegx2Jh6md1RiJk
iT8GrvjrGjX6nQvRLa7hgW8v5Weblcevt8roihrNq4J33YfZIlvgsxt24bzY5MfA
+BKfnny87KWFAv0VgHRR8q3ZUfVzziQTP3hQ8SXS3cu4i9bBo7hDvVc/sRa4e9pA
huWv9FxIRihKxFekRhSkWm9380eKJlVjznufVuPX0p/zZJec7YcWdeIaTDEONGaV
si5+LtsR3p8xcLJKJBut4WZ2XMf5Z0lGOVCyPUEU0sTeR4l0XKwqAcf+eCL2VcjY
HSwgcGPnWPekCRrRzwLsfdFVWOI7uhjNYwNHZiIyUUbciJr+gKjDr3LmOXSKkRye
BTDP1EfOZfwHiiDERVL+T78Ka+L3VzexLcrNObMULm0bHydRgJvWQ1Lve0gsAjro
3UCmDNvFg4X2h/sslhF81hrHNOOypxqYGX4su6PrSdd80K+gnHWxMFyszswc0aJ5
tLWxLz/vGl8e/J9ExlDn3PKF78V6VgUfph5/sj/P4b+Kxifqt2uTR2DU95+WaaoN
P6c5uw44Ri9K9in0CVJVoIIE9GoXRnYoFcuSkbqbtQB+NWjwyzPHdqp3kCuAcfkl
PZCEF5alloI9/gR5hEIgwdZ3dyjoK/IXzYVe5tY4N6z5qzmBums/Sd1SR1KSzTsR
4lwVwFT2vMta0Ht2uF3F5I86Y28gq0YLk63GkLnsucEEyfewtIOb8ZmM2qxfrMpx
QJc2N0IZy1dyd+3t0NrkJDabOxcrCFwqROA3DK/7/rIdExXFGGCjtPISuEeK6pyl
6rAbLvIMcRY69A6iFxppO5h7jMYCAGYY21FEzse1qu8BtX+rW33W3PAGG7VWUH2F
nB6ZYmSs4vkxRfQp4dJ3Vp5GM63UgGUBi7oHwEvEu8KwTfxhqdMMRQvydtK1fz3R
lF/dxeLNKouc6ZDfTfOtUcZ0Kzxi/2ZkWAOToun1am999NhN5BykzsTN/iOpfxkf
xNFFAkhMa7rxjuiiUTxMw5eO91QUE4HI+IIiq0TZKKy9wxMalKy2a30uNXww8g6y
wb50k2vhqVUddDLSMD2c3p8dVGxvIwC0yqtpjHKq8a9yXBzPnMzsFn8P90kdeZLq
WQJzwTA4rW+ARrD/oe0m4o207Q+nRExV9nctfrQBJ2hTONllEsRSTDvr+RpoQXeR
bqMqm3BSdiRoh7QTAA5/siLpRaAAAc9poOh6TTuRGaFOOn7UyOjNS/OtQKAS7dEd
/ggkXfKjRYLXtZhL8QcT3UPWxDtytkBSzuFl8IMn72Xiu6ZdN9rr7f6TpPoItWtA
wXnkdF0IScDHxTmbZL0yuFGn1HN5+8Bj9XeDB4Ssdll8/anHQgWog3XLbOKw6KTa
6XNG1IlFAXhqTsGNslNp1DMPBK0+qNGvHBd24blLdMdSjL4HL5+vCpCjC3r835P0
jxniUkfH3SIWOKX4aYLIWyXJ3CD2sDK64NXKbSJ6fmOFlVgMPe3ebLWA/OVaaJ0K
a2caRY4veN0HeepeINuRYjgkee/9x8oc6QV1knm0fn6mRqEw16mXtdVnGbNtBScM
ethSzI71z6HOhY3r7vjFTxoic6PqS9/turAwdbmFBf7peiG7qs9BrqikGS+KY02m
mEltZ5eHCggYtDA29VcSQBgbp/lY/aBcAOhsluQ2tYhhZYGogRR63uKZ9F5gqI+q
YfIwtAtgxjELz+kczDkE7ezViTYXHws0GJKCaH2fmBStv7+SI5iNmhT2MvziiJt7
CBR8cQ/XAhGaHqZVRQv2hRiidXDveTAJp252PJoBOZUW3hPMljfxa/jZax8KnaCr
jgp2UbNa9v/j83elvdpStkFb39JXdBz+/NDXtWUcP65EqGFhhQYV3Q8grKm5BjG8
6o1YfFQ0INsYVvANIFbY35zGDBY8PEinrq+CMwGTedgZxgXouBmGDdX7lPNpn1/B
c4s0IeeXd8m/EFV/yNbYexVdgHv6mIVlXmrOyzO9aQGF/zMYJ3i5hnPxil3R3JBh
LqP3F0Trc4CNuvxBslQqUdPfRHvWkSabtHbcclFlVwl3MgbMaq9xNGjfMUgK/RsF
X4jruA0p2NiW1r+SXyRzc3lYsm4uQ+Ae7VT88C7vCWPCwTepLL8O1S8dxA0DB2nh
Ff+hnqimB9cG3g0bUEjv9z3ki34P8bOHWKGUvBV99OJN/fqyWCKE7BV2eJUrEQVR
1V41bizqUOpKZHCjLMdVG7YBJcMgLpCC/6ubJrQ8Wim6LBjerXJkoe7YQwD35O74
RxY6AUg7tZ92QyRC4jd1gwKz34p1iZA0uBrnow0Oc94XNdiX6gz7id3AR/gGg9Iu
xLLk8npt6m244AT18teL+VLQvnwhjprLTQLoVNMgDJgHdkZeYZ9TzxE1s208KgKt
AAuowGUspZbbtSDcMHQg01z9+bpPGya3wkJRsy12gYrdtROGATtAhAYUUfBgjVsO
ZxhCItxsUrIoztxMmRSCK1C2NfjB9YCwtJApJoHcYEE8UVfVj8Q+rY8H1rRbpUYk
jp5k7+jMk0ZLfzYn8p0OP8LIs5rI8Gqy0gmLQ4WBN3LTM1YpNFaGMH/hy5e5PHOE
qmI+7/9iW/QFeQuuWBolj+X/n6+eJViBw3atKmnz3gJtlbyPiLg7wRhOvfLKm+na
I1s9wWzqNaDOaqZD8aMS/uTjPpPoVjaH/PVQ06OGbYKEG3WobP9/dKz32M8pbZsN
7eaDLCouB3GWSP8j9gFPkygffS/xca7PbessoScWbpWD38HFi2nklP4hqbmL3yGL
sqh7Ohh1/gMDQbn5qt87Jm1KO79J3iAvFSAiflODeaMBfBOFKeV+eRGf068Jm35b
rIW+eu9RetaqwE/yHl13lnqjWM8g6SygQ7GdsDuUMSj8pfUtlT17kW/9p57JqwYJ
5OsSplaUy26HR7k+PUZLSgjzYPIuxGQN1OKsH7yc2YI+rJ2e09FKbynewAISpre0
Op6VQu7RydbhJ4X5Wfdw691DYKZUx7u5qoHJOSIV0TNyZtF84qIN/W5Ge375Kx57
3vLjmw86omr8upKOs40nFl5J5glYdvPYBSlNn/lQ3MZEJRUy0mhR68L2NXvIoGfM
SlipbaBDx/nqNSE8cXee8Yle7Dl6ZT8n/z9wOdcLiDfTGpseJ+x6fBlANKsTvJ5c
cdVKYz4SKqHbzG7zP6PCYpvv/OtQ1Lpwx8aAfdUWG1HHzYWZNmIfSc1aNNUjQNIr
kg2WNT40wZD5p8IkLclfwDxmJFak1LK5O+i105mkqgDeOPamTWiQ0k/1GjFJgbqP
NFcWg0Ee4IwWR5eCJIPrF5Ml1kNgPOOuKIGVSAwaQH2UmHOGWl1bXPK7CtStMOL1
6g+HVPhg5nWY3VW6qZFG6gyTOtdKeK0zek3JLnGEG/T8Ol83z9LnCnopM8xPzODr
DLGsbWROA54licIUjMIsWLky4UgK482Op9CaoEp6nV4Q+JDwDTyK0NvvNRs+fyy1
F6fFGy/KABLWGmrmrMT1BB5fqg0MNHN2HlC8t/34nyt45wTldHIJJ67HFMdGLoez
KWvW6k6co/sQeyxutR8L2Zh0aZJp22GQ4Xw5qWJe06KLI/iD75vtfCrw76sKUveg
SDc+Ld/y26M9LK53hrMZlz9tE40izrE3SC7DYtbZOTk5Vc/c3DuYvzBdUWjk5L6e
GWafGyiwF1oz98oTR+nxBgJbtfxzTXHvQFiDHp7tofP57+y4yIfoD8r5jJBtixRg
qyXGpRVLQQzrzt7ntff5Egmvg0UFOIY7GAeEfk4KDVbLAx+lLVCTwsI9IuRR3E9/
zSa9qZQo5rqQGGiRI2AL8z3gKijWqmMXmhTGsWwKqXWkLoba5HDf0wWB/Q/Ol7d2
LX6R3y6mHNPkeh1U4z0ywJgb4MPMYyDnKsEDXBPC3sz4OE1Lge+Czci816w03cYj
zfdVz+356AlF9ofIMQbRTcd4kPMWYYqq62XqVkNXGZWYXiLjpzoUqcNajZFt8FFl
nFK8P+1isIEKT/MRFEVzV9RfMEJg74S4x18uURcuv/mkTiAXKc7TK4Sgyh10zvaG
FXvypo5XOJujfWnM12G/ol/i3HQ/2YN9pXgcuRaTCV8TORyF1+pYdr6pTzUQPT8P
Wm8/Gaqm7e3T9ZNscAQhDoaAlBwCXsnxwm4bza1VSoNkxL4YGLIA3663nh8Cbb6v
/qutUWq7tAz85xoW2t+TYDLGljaUOEp20uWDdLY+5B5+oUpaEvrd6DyrqfvRKXLW
Ht7JS8oROGLWShyzzN/gThoi7WA073Ulcok5V69VQ3uWijM4zTgsbId9kRhDHzWi
0RxcLustMbQesl00pD+xHONW2qfbxd9wSEBSM4tmZ0ra3TJ4+afTBEVwpbQeqq67
MaEZB0YI+Kvan76kIom6vbu76Hm8+FijM40j+nuOQUY3uSg39BRm6+q52VbN96aj
Z0EOphIA9WhJudH1JrZFZEAck+M+0l+V67Hi0lWxFx3GAeG056P/ErwGyHvYixpw
cJsc3oz4B0xBomFSwQwEhQq6rp82wTrZomUoqXV0LxAF+1byPW4C15tKMccwiHgo
d4dcKCEcmMo+BVuxumHE9ITc33EX2/8KR2+RwbNmN/JqjAwhu/TH59X/VTIjqAaB
x4FyqzHepBMN061bmvMU3NVXIX6FrLJLq9gURUhPdNvwhhYd6SqUzekn698KkbiT
6riDnSB0IOrc/VGs+2Kgu9RRRuO1Bg17NOWy8LY6c+7XmG1ko3/j3JtNfY7AumVK
JxKfh2n8wtgaIKNpVw42KZryZhTrLSFCLsPuNecoi2guDFKBFm4oLROfUTXIewD1
wIsM8vfMBj/+aHuu0Ms8lppM+LocX3421nd1yWhefMJc0A0MmO0yNiuGxhwvYGCP
/F8unq80hoKSCmo3P9xU7Bp6YYlwegbaQcHpToKVfqQFPQxx6hwDbBoO/cO9eIW8
IzsJlD5dxNxxf5gceWeHEsePAuOj87QZ3VDcOGUm2z+wiJYqG3Wkw4aUSUPD9ChG
aVCwnSLkqk+vH+psSmXUixg1UCk4zfzN6IlitZFtsaxU53KVaPDZuXjKjUDryG5v
NwHmB8wfiS/cBuvijjEOg5te/OIiqISo/b6VwSXXKLJlSiYxx7CtRQ1WmTVlgdQa
QQL8GXBZ8gD8QAIf2G+gwrJR3Ggyrg7amQxZDxEnV+ecF1K8cHIbEPUhbjjr7OEe
dBlAydYEBXLKArxlbZZ609hhVnosp1BcwunCziKKAfn2+JuxaSnjHZHuDiE1jFrA
NouhZxPSuInOC5mIxORrwdcAH4keyFeSemekXGRRkMofOM5XZk2Ln0LkfFFiem4C
9LaxzTcR0/ZrnYlGE37o+/nOHNHewpYQfvGxMMcepwQjeexeZdosEJ8Q+zQ2zDxC
foLlCSHz2UalqVjJwxLMasn+2a6/OAvd+fbFwFXIbuJvcam7F/mV18G7mSGW+PPs
cgBCj9QynNe/X5ESOKxLi8GvrUCgMRPUcYyU+Ba+U/2ZqIyThwZLcqw7cVef+U68
v98aNNHwWnUBRskZnl29LnWqCCQVewgTqUCw66UvMvWdaFfiiEhnNRCePaqZ8H8f
XWkn3Fp0KJUePsuxkeXdfRcOfLvGlierc62kVyyU3OR0b+2SQU3Xg0OFHgOVmtpE
BLQwk7kGQBvXaof7UoFRSp0uraK7cf3EwrxdQ9GnXJXJ0sFixpMPtn9gKNMIsxmZ
DwF/7dGCHHzjbW5ZUZiptZO8X42Hrld1WYpaFhhSB27oVS3kE5gOsMrZPpJEKxuZ
HWgZmxWZrh0lOl9y5LS0kGWJJUn73UadWMnXnQZIZgZfWbMkWHscHmaX3mDTxCXX
adj+ATFvcpLNs0yHKq72+Bl6JJMKuRuqd+L9QTKXAxX842xjPDb7VcRNzD6pRnq+
/W2oRlovEwB37QUG7y8OzrmP+uv0TGDr5jZE/Qn4TA1KlwaDiTWBQxKCa+EIoEbr
0CPUVwv5eM6gGQDE47HWGm3DFg363Ll1K/lUV+jpz48Gyi7O/g9zED8vu0xXCsNQ
a4dHLTd7sFGTIfiebSoxP9agkPWHKJnHBPpGCyv6G2XzRfQSbnQcWqlLZGRLC/h8
9VSL7xSahVAwjNJWdFQcNGhp+HxUEDAuKNB0c/TB7mwDQznvAioZqLiSbZen1IMX
4/xuObaxqup5jFcFp9nsNhZHax9ABqq2a1/H2DTp1U877KfUMxEX04I8bY6FekPX
ZdOCqj52J1p15i/ZaBgXc4/GQ+uReuNf2HvvpA7O2asGLIpuaOitM9CDDhjkjx25
3Cp+CdJw+NPmrkC7yoisbNKfPcby9QutXAvt8/9PIsdePqrVWppY5x1MGCbcOBFQ
lrjiWSbzQz1GslPDbivNzBtFo9bZS+r05rh9YJZuZPB5Es+OIuHmUeZ4l0MUcmGW
PoMb26BY8YXPVRyzXUQfmbZiCvuowCiKw3kCmIOgJtRj86kNW7rug0gKm+HUTb3L
4FEuHHRQRQWkd9WnyHOc9lHA3ffw/HB/IVDEPzSCDdIShKUkXCz1CSNaC1gWlvIw
O963ei71VSZ6cDsLLeaLqBRubTK/ZH6v+GDO6xVj8YL/iJpJ/2khbSLxStaybI5E
OBYkDZYg1FOdB1VDfW0XSkCwyGJcynYb4TMiG2ZDBGZrW4FFg90wGhkHIe8tnfHF
XrVSabg2dPparZK5Tjg4Eh2/gNVoLG0JlEyVsGRqbhjX/d3AYGsLirFY/BLbii+z
ZHN0073+7ce6MJJhEAZ/cGbvR0z3Xm+0tzIzSd6En3PpzpKWrVDyMInYCDAWJjJI
Knky99ulY9PL3wLvgMaaQoiz14gx/GGYQN5dntrvHS+fi2rDRtQIAEklN/u2v3uz
erLUBvtpy0RMEKpVvl0asY4LmyxZOYSYTGnB6E4ErYbJ4iBehVRHkgF0GOKjegNj
jPFobDFZ8aA08B4JkxgMMu2mmRqa1hQV2lFtRQEljwDkF+Fr11VOn3+g23DdG8n8
jcECTnsoQOW8VJXkFI2cr5nvA8KcrKmFj1CKvFTkcd4TQfUES6ZQnYGLOAp/nc+K
fRXodt9d3jcxNtr63cKzUL5BChYPQcXBzc9OaTtFJeybOSTo5MZd0h2Xo0Un1/wj
jhS3R9C835w50fwRfvIDh5VW/4xp9sxlQa75pA9XSWJ3U9ubw1HRWyCDrN1VJJNq
pLxMVScg2dYEeNvvD0Km6/aqR6W8vDvpOUe6HXWPjEwm6aNS6/ub4YcnX96j96yp
7Xq+7+77x29VakoVS2RVVhZQUMiJqXUsRaz/kvnFCLVjlXGuG66IVYM6Yafekd3k
iC+5N7E2+ZMIGpKROPRipovCQWEMcFQl1wGIALZQfQ/FdYoHNymCeVmQwhZXnzUK
oKt/cbXQqdJgQmXyRMAPTSHxjCK7urjGDLazSoKaGK1gtzTSstkjpB/iGCrbfcpj
yL3pdLsRWqiSLdYlqFc5RWJ8ixCws0m7ZmYK+9dFA7dEz+rbSv80GvvOV8DEODMe
TM3I40Hszid3ETdR56cB8sLQTbFIkbAuqQoOCEAyrbhhIy0yIn7VXZnMYziJRAyG
NG7ifTMF5mZIgarSEuni0GL/+kUcshhTFxlNfxtVB7n80N37h5FRFBEC/WCT7+Bp
AeA/Pf1aZ41DdnYqXQfR15hK7PDHFpM2hDxYaNe/4IIRzj0suUnNWTWxBg2zRGPf
LC9i0GzB/dzLheknR2fnvrxy19UZr1hxqAi75x9061FGSayEXig9/ZT68yvCD6g5
35qxJx5WKOO5rfdFcZ36A0EUneI4PBseRoR+KWpUF912yGdGk8WNAs/p1o2830yD
1t3Vzt2UK35y+gxp4jn414IdDKvewOUU6afOTPCbQ+86uFxDweJ1hgjRodcu+D9x
cgwjd/pMudD8fJM8hslFLf2xyfcV/c5jb2EilBukTMENJAKWPi6V5R3p9DUcDI2H
I6elOBmrvi4i1dxtAeOF5jHBQVGJUGSHoY2kwVxm4jVX0su0vxLrxFrP01YhIxj9
V344Rcds1JxH+rs8lxJ1YBs2Ea5Oyf1P83UiissITURrpIaR77Z1LbHWESkbfRUM
m9TQ+h4MS1xM1nsFpDwokH4soVAU/QjMVOX6c6VjTPf27ff9RpXwLCK80dqiQAqW
4fWlK9Axh+canOwQyddHc3P9Ugw/45uCxZv4zPQFMFNQyyPhtaO0qe+QAXRUpRVC
htlluzEgnUsO0fEfYudtntdx5Iq3IkMOJ8NTgBhmitEMnwPZrss/+59T0PEjW6ug
QlTDWFr2p5Xh5PvE3T5uBHM288CJft3nBx5DeqN4oE7l5Ya/iTRV4Ar0JrUHlwK5
U/09bUf91Et7fR7nOKMds8ulS+eB/inbaDOBkB+jl3YeanIAVjf1oCC+7O81dvvI
wi0uBboidhR3msg3oFrBUkApp6NwAJ3/CKBhfuyi/2xxQqQqTeGVF3CI2tBD+unq
oI+7XJCfyZSWrRRgXocOxKXTPVZV6+Nsxkzn9+N1Q8OEc2dTygBNQ/TrMFvcKUdQ
L3pxkokX1eCK+/L1Zi7W1wOvzJomh+sYpGeF6NRIprpSCQcmeEZC/JQ4R983kIPn
IlJMJFaGA2KH6aPL50oLZGPCiL6QlVLKGn7AOJ/SaKMsbngSksx98PxAWWwUc/1p
Ehm0b+4uk9Np2PIxS1IFW40ZurTqpqIUld5Z30edx+oTgmSOQf8ri/2n6M8mSYB6
e107g3kYBoKwaGVIIoV8k2CqLdaZoE9pWt2rJTFo1RfdhhiAMXfRibT4RsOuAwc5
npTbg5V+SQZynlL153IiljIf3BXcDgl7BKarbpGF5fR4JGP3GYnM8B/2ZZ4tpT1j
vVhaYRpumlzsfE//rgNcLrMuHms0fujapZ5xqEWGFKxN2cmDWuuvtZRgvfPjSIYk
XIKtGTkc3dzJC0evkNlUtrEK32gA57DBcZNDANMeR7CiMuLb1XbGajaVI254vMOU
UnE57919gyEjcvx/txW9JjydwT9aZVVFF63K4fKu2YyOlnsbwxaD/ET9Q1rexuK5
LF1CeZ2kFmVIB9d2FKiJZkYH82F0HC3jIA1J6D1/WrJud0l1m6+Fjw93+Yn8H85W
uQ677o6e+Mu8RUVw3VOdpq7zOkXoaapLiqNa5hGXMhr/FLmahSq/H/9nm9qmweMz
dUW6Cz5rtYq/Msn/xhuAk47gy2lAWt1HObiF/HJlWuGN/PTnzgKvzhaqGTs3/0D1
SZ2/PHC+BWdGexGXkzDUPWOfUuRktBjYUTRNZgCyLVOHT/CiyzwVhFLCB5m+ZYaI
vCX+Umgft/vD6+0yhQg/85rOpEI6GRSFfMPiFmtV9ORng9+3o3nqkpYba9XryGpN
NpScG5q978Q46fkWAkdm6XGa4v3KTqb7SjIHnHMqS6aX/x6+Crv7r4x3XxgSqNdJ
igGtYAwjGdFHSOhQLZBjWGDxIvhEW6ZvS95rM7ZQg6f7XTw9WqGBAlWUxDoIA3yI
fxciRYcgENNy+kn+kfJRFKFdMrLzwIZl8MXLxVTPk2VkAP6zGcsmgeIxGSw2vDXi
Yj9jpA+2iubY732u+TCRmsLFhsOMKnViyWw5tOcKTe8aAt0a6I6f91896PaDjFsc
5ojaYVDchW/FKG3t1CcJfLPOYGDKKG0MTOfzVjvbBsW59vbVYLuy5fc8kJ1tvjO3
2BcCkidt70470ueiaqEnnj8NRWNtZ3CC9RgzAX77Z1thb7t8fbSny5eFVt2DWnt/
RmwkMKDYAllSXbEz1DFh721NI9rqO2XXePweNiTW//IzcCr5YQBwAzSv4tsMg5y0
fSANhjYQ72N8pTEKVbn8UCNy64gfgU8Nmei832PKjFKoL57FlUflFOl34KrzHb9E
QF/GCUql65bX00ol7ixUtifLAgia4DQ/zCb9LvHxozz4wpRVyQYHt74gNPKRmA+w
q1kvArFW3Q3oz1ArW8ux3bFUasp7aPV5a511r+tfxz1qEfJsEIJGjBKnwrURsTvS
kEjhQY7Y1rgJYfZKBBvHPVFQeQonDO3K14EW19zt/QXFiMVCHoc9cOZaZ8s8YyNI
8dE5Kz3u+QhBLoQuHdWWwsqLiT7IpTdMyFHJ7OdCGrDUwhc5TqiwZepyZe2hgoxx
FrMjsYaaMnpWFn+UvW2pwW5SrGf6kiN3iCvNquSBVoiQjtpFN+07RbAD0ckQbarM
jlPNfw08qtWg5k+4+EuEY2PmSNwGCKUmfgBCWEH/TMRXNqlVxriNdn6yFIn3HI3H
7EzhmFsKucaeMGaGbUT1mCCDFHfFvg4ejdwaC26KMiBNGN7WvPmzsEfVUkliXkfq
kkQ0OzY3UPtpfkEYHacGWQntc9rL3tSlSeUh0CZc2rdfj7lrH4+RudKORCbWl1D2
yhnMxd8/E2tAQopG+jv3jxgkcfhWEfuHXxxbQCzg4tELkR1EM3/vgEnulJMTRADD
zdyygIEYr7sMQL04sWHLLrAHOIxR8AS+37ryW/gtIv/H7wONnvrNmNvMPHFnB6Uo
35OnljogM3pN/9wPJaoqUtPfKV/V2u+vNEeDrqBBUXh3Vo/rICpCwGTIPx8iSrA7
pJuX/n7+cJTEK5miSFh10DskK90ThrnnYwgRpCgmk0k6tXweKAxo2KCvI3gqdLyb
biVIPNEeB5oBvpZ6gVpwkWJmRaHhlpZG0OhVy25JDwPDKbMSYtpK5sOrwmIlLkyl
3CTbVxNIaVYBwg5XIkXKHJ7m71MR+03O9MSIKm0x3gSpbmdZGhdL/nqRqSq5ULFG
WV2dV5gFansNnLdAuoU6UcM/y/Mr7nLAgB8ixoXa7CivLp/PzP+68O058khp9EMy
A+mPdfjAOob2qpHmHPyrhh+Zp/RfPOlLsdamAAkr6tDPJv031tfUGP0PQps69fuN
Xc2B/EapcvzQAbOBVhLbTU19jTnVkf9F2XI4Br5lmSI6EHi+Ztl3lkNrA7Hiqugh
2eBp1LZl9/0JCiONEDhnoQ5cFO1jBb3cnwsUR9iwZvVJgMmTzZKRtpQsUJbrLOWT
edHRU8NMUqgww3pVae2np9DeknwVBAw6pkjsU9vEVGtsagGFZvRDf9MYpysQMJwd
stc8jrKCdk2I5RoMXV28fNznTXHHleD4ed1ynr2RpgwtYEuf6ZOUU2zOjMTGC3Ji
cBgIJsLd8rj4fa28a8x3MTT44M1I3GQlm3fvDVU40FS8CQBYcfq0KF0KeIghIakQ
4ub0HOMaiPNwnwUysJpnXw0jbcpdEcbHiGqn2hxPZMowXqTmag/sf1tlzAtju6sR
psskCrRxFNahdCUqeiypHiScwGlP34Z1RZ2gAtjFnVjSQS8brJ2WMfhjJf23izrg
FI1Vkxc7z53l+fbgFBYb1DvD0EObeDk/2ClaXzib08dFQQhKwEZpW0ARSoZ8gWsn
Fdjlrq0PUvAZdqK4tpJiMx7REuBYACXC/CIZIrqtnMWTg/bUx5HuSqnasqF7SuBY
YoZnbePxO6VWeEP1Vzz3n94BOg64DHcgPqL9xklxbzkvd3C6PvKGu1bGAvDVsWYz
PL0PxJziqMFyu2EQx4CSwH9FRIwFgBYOnYAej+MiyHIu8gyQyWgM3rPOw/4qenov
PsaXHFVyCylyNl2qFDjcZ8iMPyG86IEq6bin2ljwYrLFrl8mz+50XV60YsEpt42K
zy1wM0D8qiL4zcuuHKk6/VrgNmuVtaMRtcijWOD7a7i8VV1XrlvlpXpQgJlc4rfK
5E++Hm9DuTmOHw8HY9Zbv8uyEyAojDZXvB+tOf956G1B7l1gxm2shkez3dbWeRlp
sUCYtHwkPgD75yPUJ6zvUDaCjqhm7VEB96XWm7yFJLevTqtRLzBSLpEz18wF60JF
nkqdBED5He05agawJV2KetivJ9B93UfUbpQQiTmk7HXm3qNGls5+V2qzIlXhKAEe
S+cJOCIGGHYx3cwKsRbuAhDny8U697bdWaQjR1PBQxmCcwlI6CZYlWvFlkgScCt7
KvzVpCppMEFh3m1rKzhqQsXN035VjFdYUsGomr03/9qlUeDpwz4ZtKr/b9FCr8Ia
R8kxRK2pnY4LCj21TGVwgSF2FNA7GuxXN7P+UA29ybXDO3D1PiX4+99wwy59Aa05
+w37SNulYJnPnGQNC8hc0NwPndORZrG2u8Rr4bu/C6hQhpP6ua/xYBfhkPq8xafo
TT1uvx55qRocQEuBlt+HqqDJ+Pb438eKpxJrf/6WJ8dYYZvOxnYf0ajMcrmy/pYw
mIRUbez964h/J38K/zfra8SpHxN11J5e7co3KP++Ike7GfbQlmyxX2XWjgzkMIe/
fW2pAUi/yyJPs6bVbeDPVsqx0woKQmDihWOAIbF5+9hii8K57zQd0NofU9EL5XNm
0vc6wrpSJeVerVl1cLcy3Hniua7FWvHmgNlSRTjr6uSioXcKOKhu/x33d6c2mx59
dUbD5PwRQL1UKtnHUu6IL7xC9oO7bibJv6h6IUeWSclNziQCmQi3XG1NxrIUgwfE
ry0iRyBaIsk4fuAUnOgeZn3v7AAZPqurpu+UlPx4GA+XMN4t1tNJzb51jrA8y/zc
o+TA73p0RKi+bXb611Fs/ZQHFlIT3PxZSA4Sa4XdZe0ikebAsa5yrnXTMxqBPad2
UZ7WPtX3YW1VKeoS+EJZHF8MV9azEqIKZjsdcH/E6/1UmagBmsFxav7lqlXi6YAa
dsEX005V9eRI9l3bLBhp6rNBm/iz1xEFlS28uZoMwjgvbjY/Ol8qjFe1M+WDZOSl
5wlCOlLhchB09sGtIiamlFrCB1jIhlsSPKhPxe6RtLJtsvu/rtzkH7+GJfQmIrFl
W2y+H974YEWjtRRRmlbL6M/xO8hP9LcQO0NaHRp5O5xYxnkt8+cVzVsleqwFclwP
PJn8AvFI4Bk0E4dCn2/oDpzNDPjhWOG2sNKFYcvpmG7k1zPO8tKQ8JhTHSYgDZSL
2FDD4JWB6LaA2rRTNbyap+wVy5PXLwp5TH6n5wuLIOj7g62JjKp/XFfJm1tZ6Gkm
KcFy4rkYykAsqDFHSUR3XMKx/hzdGklbiSBNE8lvrJJ118tPu54XBrQzwdHOaEsw
Tku5rOP1VJJY955SnWYSJViWjU/PsbpeBu0LeGzfi2RVNs/LU0AtrUN1WznwehQr
b1cqG2iwaaHMbCWbAHN4aVGelLkX/yfyy88Tojyou4LAK2AWtqoBxymKo4cQ7myk
qhWnZWkB+P53FOI5NPDTZ2t8rxD/uIpNW3btUTWH0KseSP9iTs4OU+sPK77inQ82
Q1DijeCeeakFhRoh4sfNWzXKPy4uPYGwnjjrH7C3y6CsYe1OjogWH58z+uF3P9yF
5qdkOGDCJiw9tAlYsA/7WKK1zhDZxdGLRgeIk1TlHQkaH6ZbUdEISzx6n97IXFzN
1vJnS9a0P7+kOiirUzk7sygA7fXGKMmYcMT6hSDaZ487CgRmVcfdxORQV2O7KMzV
RgJJZh+ZIs/TIW6vT5wHRmk/0hdkeeRphdoQfVVjPkE9HYxmWd8lv+vET4bKjMkl
ces5F3rvKZgZAT0mLYLuxkJsGvp/LoYH4BQp8QsYajaFE+E8R/ES8nVu3kD/N9XJ
NGrgnWXVTiIzYN+r0xsRc4imlOrQ2v2nAx77yREU/2ReLYjviKEEpiDeiCdtUU+I
dx8L4J/ja3l2Knkr9f03OxpPIkStoQAmatsofxbwFrLtfh+amIq0LSmSLAlGIcnf
JpWQ6fR2yfNqxHxO8Rd+BtBXyHZWj+evU++kSlZUmg1tZ/SwWxfsVNIEW3BQabo2
3OSEP0yu8RN3vNJzNtkmxXsdjrAeiuFRp4+hOfdVUeYwz0pU/dYtqdoaKpYCB6n7
u2opYAhKWRAScVhCz/m3niAFK3Al9PFCEhUze49N9r4B9MlaCh5v8AXQRNBRfFaM
U1s8pDTmzmECS6LzooUO1+7u34aTERmwarg/RG5jAoqTHuKOyvKRoxExIUKRlLLR
CrJvus7Yer5B5Q5XTLfkgOagIj1FB44xjyamaZLCON9PoAIBcY7iWlAIqoo3P66o
bXDm3uHJ4jbjeji7n0SWSs9NbbYCRWlyS/CN67uKpDJOlS9TxUoj5XyNndh6GhFQ
7bgw2trWasXvUZKvf/0xM7ewsYH7M15j/9Ys0yzwYKfRaGj5WGsGJpAOkZXnm5hN
Jpo4OQ71FqvQAtdGPg1TR/pTlmdbREvSJ2mTKdJYvI5aQ+tG4r+8OwqmmT6sCcKk
zr/YA15p26bX9TzE5OB/eTQp99SExjEJMVVAUed3upys8cUrOqA5Qh79C1CaiJGy
ISaFbaEr5X6LhyxWM3DdmKl753vTlQKxnNrgNsbJs2r5ip5CUl/A5DQOg4hFSvuB
U/xGjAakbt+EUFB0A+M9Oqc0lGeaCWV7fojD4w2lh7x+P2vpZ7PObkFPKz5o5z03
ZR9HdH0oAbML24nD7K/21WQPVTevWJUgnGsS9x3oBYVUNS/OAdraO1bZvD/pdZfa
9RmuMtLglzMCjm8RV51hL5jLx1FRZvrD0Szeom6wyt/U49GOVU6HzA0udqYIEdoA
2hf3TMnlk0VL8sw3rwvxR9ljEYd1kOsA/8Tc3rgATGYcx8SJWbqLhkihHLaFCBfQ
XVuiRq6bU4bn2aRoVfHh55zfXj8qeUnibghxzygLttMNBHaxC1Ad2/mPb+6dri71
k6Z7++Ka29kdS7oz9LleQiHsd0VZTmocNv7vMO7wV6lR0lruXO0fDLUSsHBwnjyx
TCK12l0YLx8F7aXTU0K1Q38/eyiXKBTn79H6YT77dVLOQvp11Z1rOXmgmxyRo2KG
MFmI4fabVpHvEqjD5Vbh/A98mql0H/QWkHniJIuFXbzjrcyoKNZPIteKlj7Y+0X+
jz3ZbW+sEiVqjGAMCedW1ThV22PbVJ2tty4YG5lfoG7+cnTa4aP/IXPm0ih7zYV8
BOKbaQSKSq2fFcVq7iZ3fV0EKwSMt5uDOEsNEQa4x83/vdRi+H2zzFz9MevJGDPq
YxmM0Ale8CKs0i8jxkysO6/qIHzZkBYafHDgWPgQohUlNTW/XrMnkfVbvSnedT9a
cY9+G2MlcUgO5lvVhrwWprTc86UL9EnOUtZRBRHtD46HwhCVZpFXBFWO2UUiREE+
4yi/ruOsBxJ30dsaZKAmNZX9h2ErmjEU0tCBxjdu7LiyavTe8Ld2Qf39e/Izu7za
aPOqI4B589ffbO1taotKS8RGEBc5d5lfGTst5qVoKglYNpyRRiOeR606LspnfRj+
Li9jDwoJgLxqinEEIB313ZSf4Vr490s3yJwiBOYBJZ49tSyRbAyoBcHjvULm3UM5
rsYt/8MqXYTePiR8U+a6KM4elwnoV31OmfJ0vp2sPmFjVg9KhTwjJOt8tTbWidJf
wtsm+nVv2R2ba0ut7jrxYzbR3z7DAKixFb+YgXJlhwL766AOiarnrx4dq/gbqPVk
ET+U0Jkgb3fI943WUvsYWLuJg8a0qvrR6EbTou8554E5tk4jUDy+3sZig5tsyU+N
BNJGzJlxffZJ8L0vaUzczZBpif26eyD9o/oDF6qoeyIJDX3BQFUBTX1xoyUBWyoM
CCrEBbBaBEGF7PEg/v4LV55hP0F0OCT1bm97NCswvFxZo2vXT+FESIkDCyafEy2t
uLtHBoZShLeIoaWjhBGfUum8L/6tps0zxbVwtpCeA8oPeLI66RuoPhfZ/vNfauPO
+i5O0p9V1cqFRSPydG1em/JechAVGgXlPoQDi8yu/1P/mhLxwwzVOcnnmSHHhWF4
je4sjE8EnJSMP+L4Po49r8lgRtU4/jMwIN9/PRZicNlM5etqqh/84UvPKd1Aofoy
AB6xiF2QrEwGCk4qyMqKcDevs4iXRg2OA8GfSRySYQAColhFFMGReQRJfp1+87g8
mrGzWVeGrWsIfbL276PEnMaM7hOQJDIOxk5Z9AoP6CIc6OmMMtad/Nvtaf8Qj6W0
RNvGyScpMhfnYICg8njgjIUPdosBmaZQU4ARCDSW0VMHDoE/qmQljG1qxJYF9fkX
eUnD7L/oZ4CQVMaQngrywuvNSQkOcPoDIAAz9tamap5gQkN2iULdxRdSA7CDjXi/
Zno7kfR8rcB2kHIb6jZOq0BHr06iSR89m4FJuJwIm79gkcoomx8iDxrILBU7NITv
V6Tqoqaxd/twFqUl+3yYhryKefGfo+Dc+Zn7EoHXQauOJHJ7/zp4ZXCdZJ6AX72/
tk6d1G4cH1xICj1EaDu25AQlsUpycPu0mystE2SCecXCHuH32+AzgyB6ndonhMaa
ulupU05f9vEGwdM18p+wnHhvCEJITAqMMUHL/5N/c7tug0QENEoRs3G2PyQBR2uy
0pPWrE7MN+1lLrMDjmPj2WDGVpEhneYFjMVveWG/OFB0qoO+nmWlAOv9JJymlL7h
Tk0zQr4lVdXaopSWuihnrJz/eqKCzY5t24ViNayg+PeCIijhsvUKSE1rXLGvplXe
219f8u/X9R1/PdxgjN7A8zihm920OhxPHAoHFmVEUNBz2CDTN84aUy8hLz6C9/b8
nxQiNxOANxaHbgVHRCRq6acroYoQkYbtkIXiIvJ+JuM+Z+c2bpREs7aT8m7pifHp
UsCfyYOfm4QL2wiBnkyF8ox1mokdAnk0vxPcTA3/DfHfdlgkm8oyHmdbPT3M+/3L
1MpXg3jyqdMN2EatnKlp+FSVV21VMXtNhKttKSftWpqkcu9znsfuxINGRK8+Fo4Z
mG0ZCN0nCJlYSYDjI7k3F+JoTzp2r45c8OtA4T8/7IsEAefJg0cl+jTTaLdP6PAo
LgvAu93rOkSTJPV+0BdjRP076oTtPPD8w+EhLCzTwsD8kKFl0CguQKwCqVAPxO4J
6fHEyVRVnjp5MVZHZtaQg6g3X5r9gEDiZ3yd1qheX90fSID0qS+10/QaPPAz73J6
VBLh+/DRT7y9u7XwKo3Mbg8tjBPhGZ6GDMO3rlT8Op3emtwTKWnQgIPc/bUqixpa
Uy8e587KRj922Gn/Jh12ekAo649qPQS6plkrPZxPUWOj6/YCbtXKOnSlcTZYydk1
Qj+zH8xzDga17Te2IhbiqtdPseGheEbMlKr3A4ZUaazL8252jM2QjzUf/lwLbFHm
DuO7B0sWG6XFS1JkZpC5iIfv0HU5WIVb389lbYGAPX6dPQHp2pux8whnyO60Qq1d
DW4c0fWUUpLNVJCufd/mcqoZsIOYVFKdUs5VVIB2htkj/5snZo6iQ3ECeVMhvAl7
wi3eZ+pdZ58YdR4aHhkCjZbU9Teoh0NXa0ds0iRJ95x6ssDAoYie3lzdPIWdd1Ok
ymI0/f32DWdWZhhk+UAybqPfkHjAtj/Gbjfy52gKG09Sl/LE3MkcAzV87VtQ8qYf
XGk+p/UMpHufgJJA7pcPi97pbrblIxW13jao1+xBDrjE0lcw0cLu/ej4YVPMpUsE
CffnjJqW4cjptkkx8ZdxBTz2i3q2q+os5hjs5BUaST5Bj0yAo/JJ+9Ai8Du7Rk7R
QSY73AiIzcgmmrvX0h4SZI3LAepkLG0BBED+vFWEkyktWEiRt+b8Z5wQ/SNVgm3+
0wsT+RzAA/R/w0QMtxciy24cag5sLIEIml6NeOGtmfxqixW4L3eXZVQLfAIL3yeS
5XBAUtwuxl/ysMvyLxm/jgmV1KUhQR3TqcL07kACtkDlfZnw8UG8lOQZzWZb5UYo
nrJ9KAtAu+LcDDUaVBwlvPlYtsC/LT3kcYXtrLa31hC1z469Lm9KtkwAQvYqLReX
mipPbOVuJaYwdMQj9ZlORR/KbihRtDSB/+aXd9ddMwbeeBR8viLZqcZ72Rcofvgn
pdJi15HFKGi0ooD3MYpDpYNaplg61A47Mwv+1zoONLUKqnh9YTp6p7wlvKVDhPdb
N1tniLemVsy4dzG1uB85L/Gv91yzOULChjkDtoh19TKzfqvdOruBXB4PW6C1qHW6
s9TRbvbgNKUnm+UuzsMInHoy1wSD2/bLG/t7jYnx/Qrgu8eQ61Qy0UwaDa+iNB0e
6DE8mdgFu9aXbbRVTeK4K7T4xWyNPnZkOqxZRhAjuOsEmBWPN7kGyFtDsKYFPVIh
OsIntC0OXcVTlrVyWUtGOcXv8V988igd28LdsLazeiAmamYn3mifqpdx0KXCkDM1
xaUHUskBFPqFLiRQwHrq0NcvFg719JHzh1V0bBXv4aXByWeNdQz3BeDsuh75zLqs
XIynX5gkxsaipQHyNH04t2jm8mzTN7JM03eAqlELN9IbBh60MqwoOoQbvqYj7Dcl
iGK1cnyh4ytu2yK5PaM4oa20P0eNHGZuKP9jLIrlZov6fkJ9kZBZa3ADcf7u5hui
ItHc4IUXesQ2aqz8BTuY7biMh99tR7CRgcicoaKS3JdSaMPQxTvIG+3PBNMDF2Rj
JQLTAqetyQN8qhXZUs9Z5DiXXjglDEDjV2rJR/GxUovDQWAJsd6WlTCv0fXtFoGH
e1FuGtenGQeYSIpLTlSlN9x3cNLTtvn605fimVHfLDLssA1KoGe4awM+RaCU19ao
OHVW1G+KPS1NRH9pn8iwy8Rgoj4bQKHFmUaau5zPkXUk6f1hhO0vF5RdKfudDevo
Y9tM7CfnlWI46Fm1kZA9CgQbKvslAicEh86J/dc6HTEHWmE6hf4Oo+wDfKNhv3Ep
XW58Y7p02V53AI4O24KAFxQ2lNW3eZ3hfjCKk7PGjyNpMiKkn0AdwdJqHh4bbfG1
Et03nUnQygZJaCTEupemUTmPjgr6L2g2o4htuy7ugzGjX7WyUoFLuMBR9LqmOsyv
0JuK8KoQ+ys8zLxbXwBFtaOCLxmba6iANUr14S+KwlvAjMrh5HHsud1iFv0SdnED
/f/AivAfpCKiVuPWjguUg6xjLqIvKO7i11D2vU9uh7pw+9gPqz1pvSVvqPJmpgC+
4BYI/AGoMwh9+rqXS/1oRTAck9fFK1FqgWvnbjpxy6czi1PJVI8unZBEqSrHKgBu
jnDMiqT7DNEfJapFXxsWZ936NZUjO9IBYJACd9bbFspf+VDwXcBC0Yzp2nXaTjR7
ZoViLbxGIfCo08i/EH2+Eca+a3hUUPkNf/oGnxL/7VPM+SPKr3GB4Nb4aKOTnVNi
mKqPIstDOKdvVGJ6IxQQaZE1Y5T2xyIjpsJx4xN/QROLOeAWDgKMakZqqflKEM9f
Yb/awmpM4obbUQ0q1NeVaF4TgzwvnbXuJqCHeWmXNoLPwHSeSH7TLcqPp2TQWAQl
jd49U5zt8OL5v094zbWrtJP6fGaoCmijRtyPcBAwpSncoO5HQfQ5WXxkty94Yd/g
zMg0hb1baVHB+nmly8c6i94X4io7Mxv9uiwQaGoJsS2tauLrq6zFLBiuXlNruo0p
NGwdqxRTibm6ekGQBSkwKTjuX4ahHyzu9vMros0lZaZ1hWEIdLyoeQ+TI0joEciJ
mfxkXa14kDucI8ESgist0NbiLeEH5miRPgJNB2YXI8G99hZTXU+fOFdkdZmPDOGP
Jxk7Glr9bfYiGs1NQq06To6U1bftzVEwKmXr3VsFzi6xCRGvMA3nyE9X7G9XBYRu
aepWDuN/hog9BKv1M1uysEpjmk+K0vWehqDha7cvYb0/oZIK4/F85m+w2CiqGubg
WOrrpJxNqm5KxdgGT3qhfCKvvREopfH71YGnrlOuImiKVDKiEdkgPp6ImAsOQ84F
FSfKr9X2SsJ5ff+d2IbNB/W9BgprxhAXeUw1iq8pJX2N7OI3+RF5qm0GnpTJm/l/
RS8uj6i11r5hIPywU9Kr/iuYFYJnZgOWNoMY3scJfmLk2hJDjkb85PutIIRWZdcX
DiS0rodUS4RMMD4QfF/WWk2wM+2MO2dpz6TxiwadoaNWZFo1PuVhtqKRZQ93YmB4
TTTaq9P93isfSoTRHcnw+YoWszPkOYTgzLVPzODUu1qzattcQeD7BR13epcZL3S7
GBUKZdAhut6jxwjqqzdcll8gmMdN3ZnzWl8kXu2LVPOxyqd9jTk5ECXf5z2KwG3g
wlBcQCRdz8cXxaShqKGZY9zQE1vxrUuUYGKItnLxnkDMF991sb4cFD2ephwZ5It7
tXaS8f9tLD4GfarMHnwLEclqTmYiSEipIv+V1oL4ZWiLkodsMY52rlRlW62MHnQp
S/LIgUcH1UbREZ6ApOQ3YMSErqq3TWQQnzLFYIGKNiZqrvMomM2IzBVNnFH3xcpI
F4+ecT1k4j7NiYHFVxF5fRVxSc+IY+NBUtJQa37cd68SqxhZaaYzPFyThjep+82M
1yOUALjiFTF6HchcMV5IN0W1T4RoPizXIy7yK03OKi9HL1y2VCIJOKoXAu6sHuuK
TBJTvunU584ObzAjq3vTZ3E/h+b46ThFQp0TGldJ4K9A6kmP8l7mxfWp5mSn9SkP
/yukQ1SLWQsStWkqFnIJMV7cTqBWVD+5aHir2N731XXn14gs5JUBLDcvMPdK6u5l
T1+pAKUgDUR3qIKQfRxUYwE/OFFivrnj7ykp9MIAccRj0bMRREa87lhIdKruHNnD
xTos9Hn2ph3d9RcmGEBnqOOVAFiDG7LgKijB6uP/juvExk53PKM/OHVgAW6HfeWP
AJuYxJvDJNuIMmYtsTg0DHfSMyGhZXWllbifyLBx9c4DVCDNnyPx7dURVvjL6R0f
+trv6sa5KhsVYNOXtgzldBqtpR4TrmHdbOBnf8Tb+eRo1E/EpoTe9UASYWdVmRsI
vb5PCRKj0hP+ILHRLb7qo8y6ua9nhuA9a2D8SQxyV9wifRMD+bsuEbdIf6HVpgIy
s5erbbZIZZHkaImMVGhLEtUlpvg0j3g4cUrZKSKM3qJLfQ2v6xj39bJB2nIxs9C3
m0niKtn5ea7k8LY0w0IHjuG6jq1RrECgPVhu24rQKlMq/tHkzim0dYQe2c4tHdw/
w5BA+uv5LoRlXWK2Urn/9iFlbiEmtHyFVDnjpMI0pRWIQarM4pz7FfL8mZYyxsL5
kWy6P8SeYehw7Oy103ZRz+GWtlBUIL+zWEeq1wPnG42DYEquIGuoVqSC+3vhRSvA
CT26qpNar/Mym/0BqIlK1VUFmwaY5BwmyyKTmQsmo+Q1DeROJ1TvDyIjGwj5QSVV
Hk6xv5aj4mYBEfFLPc8stqIKiNopoE57hOgyqL7V+RwB/viej8scv06+aSYLCv0G
uLKO76uoSHd6Elc/24m5/t3f6ouVugH6Zxxc308slOWEB10ksmbS7eGC2WrtTDKK
2+/8KAhSlb1yS2maVmFBgCRnhFt5lJ1xqYVlWJRDz1iea3bkA0UoHc9CQP41tWt7
R4dI5yhAjlhz0BUIXS92HbvSS77bRUHB7l4WwjjVLiHbBw3U1n5b/Kvp2i5GMe0H
/voH7O2vzC/CmS3UBJUFBKytbXFnDvjSirQVbk1rWNiCk2/0uJJTU+fEUPzbSr03
Z/VpdXGmODsB8yFxkGcpUbDRWmMpd8lDJncIABGoXhFy3B4qJcVswG4wdrnXuNa+
2qc/9ZeO8WHV8VyTeMBN7dHjZ/q5VQxzMfJhyNHH2r3GumruJ+zinFyPZJwSYc+V
WoL6VSw1hlRh0TNFzPaMziEZeDfMjeHsfzzaJC4tQ1KN6EG9Ee9ijvWGQnFAklJ9
R6J9AFeBferF7f0J4VW+iFW+4csavtb9tGLByDzIaAOXtUbV/g2mCwfPtDaJqwon
aCVy489FOdEB0EPxUxkndn+x+q4GQd0biSDus+XsqzyI7+3R7l0jdflIP7Cj3C+i
1TAX1x2Ywp/SRxf6NXKeFQzBPNb5t3F3SovqPAic3kWctLjG7CLNR5PfR7+k5Hgk
8W4v5WXo+4Yik/H5QZzLqWLrB/8xgxYsfDzZjL4gnJN0WKKx6/c1AQAvsKDQDkUT
72HCpkrIh0C2IRsAj6Sb59FeGB6g4otzw79rThl69UbcFUTUjRUL5pOHXoGKMveA
ukww6TrvJolCyTYK3dT17nD1ZaYQ6vtTC73qdYHEmQoBvAubslMRnsmwtpVcxA6U
JwTyUjfNx+aFy8g/6NdDX3zHSw3QB7tlUfNQP4MB/yub5ZdejKWrLcA17z4EZB21
mfNILloKegso/2Z7sFNm4SaU7Zfm+vlykIwC2UMjTjFOrNF6El78SLufNhEoXbwt
ceA11IXhtxModLoJY+/GJWOOpyuqeB6x+VUv0Ni7vMOHhMYKmkxyg5W0HlvZR6zE
6JEKtgAOVoK2AyEKgLASojSl+iuxU8Z+UlKiLFWKdSPBHzczhzgjpZuZxctFIX2k
4PnRSKH1VptPXpUvQUQbkL8mRQeXZE+VOJngChgl+1RP25HeTwp7Il9wwaEx/SNl
SPOq52VZClVGO/2Zyx13Fy2fASm+nNsJsYkz+TIvK8yCRN1TeSyIMaCdMlDEoHQy
fOSk4FKLbphqq7lLHJ+lDAjygX9r+bnwkspyMf9U1alc5hkXcQQTMKuCi8h0JjZw
7WacFPNsmm+bAFoFzN9mXBUp41X2ZKLmGkUOW/uTOuDnc7ZL86eFoNCUcLPAPe1J
dqxGMi1f5siQbR1LlfHrhAQBG85MwjbsIkHBQ39hNQg6GCYdPQxwM5/+6iXUqUtj
EFILfOTHlL+849OAu7pF3o7Smmv+hLdBV9K1QAEBoaFkUP79TbQgSG5Op1bXr7jc
H3Y4zYf06WHYLyij6karji6QYdenIB31YKs4HJ8ouSezQEhsTpqWNe7G0q6b2llQ
w/hNuxQ0VIj77A1LAigZLvBuhI+1CTj7LPm/6i53/ex6c/kLM4f76BcS0oaEPkox
wXlBbyaio7j8b+FywG+OUFxxo6u1bgJJSLgX9l/O+4HHsvPAgSfqRoor1LL171rN
GXmA7fvZ2mdf8D9uAGvBIsOtlbGbBmQiiIxzW6iAYaqME/wnNy4Cr6fsRV7/3hQq
gSTu7MpY1JPNK97hywQk/2cMyA8WD2iiDrnQyeWHIjBnINDirgZhm1d6h0kBmiuc
SKkGGdx9bDMlZwnxb9KfpAay+uGQ1ZS9/jvDTOoXTNdM/rucIrE4zbbvH46f3041
ecPCY+uN9vuJUZIu9MsIRzMTjHhNZohQF2hDwReuMp3QWqD88fQ3O0SY6z7g+rZV
F4q6sK8iQ2Bke16X4qJnFlKgV2NPkrxr92ZfSh+Ov/DOSpUJVBRKOq8vSDWb6Bm+
Vwy0L3YQdNg1iuqamWEYf4tsQBNCqDT4zt8FnIOoK2QG3SkYiBKInkjAjFjNcfU+
JztJKyxy5jpDSigcj3AT3S9Hy6IXkW7F4IttyF8DkpsKGxUahxaAtHIkIm+qr9JS
2uoPTYjeleNQh0j2fACeToQYGCSPrC7g3R3DM0Y/v2w4nJb6QQVVmNrIcJyUY1D3
+Rk/VvGuPjVg4YVDDSMTCsyWlfEuMPUNg1cQ/iSrbPd/u5DrkVjBfcu4S5qIbz+Q
5TZwXFzhU+O9GlKCaGzerIw+JzwbHlQKIzAnEDYBW4JsU+4VeSw2Jz+kEwMwXDxV
Iw6Qh6G5+LytXTuYglQmndfTshbDVMFOreuZUD2+oCEpNYBY6HU2GBhmxyTFYiPd
pVr85iPZSxkOtHGO2hvQgxy4tdIjT3IwA1whbELOkpb/4hc9epIJ1BnfmeGUv4NW
P5sNuZqcmBzSPfhgn4zvrsfgyGhPcNu0saTcHqKGZ8zFpidmSHA2E0jx9PfDALDO
zfR/4SW7dRRqb85f9GK5qdPX47uU23EPxypTh8eCy04M2H4NY8FZEWoue710QcT9
NABse8rjpApdckUBAu1FupqRGvGARl0Xvg32nZDlRTY/WFxCZeRUgrXq5NtiEPmK
lWNRJq+7gCu1dQDZ9oYrgR01ExxkDIiTvxi0QcM1DrsPWZOuPR0+vSSstWx+aL40
Q/OTqXBwvMEyFYY53+blQUpoPfxQV4m/uLiZTIzjLu73pkjqMVMCheRt+uTYlkKl
SfJI1ybzq0OW7MLNfvkqn9zF0aIcrAgoOVRaiuP07v8ppy+B4t7Igc+vHtcIGcmW
++3pq/JgIxjoislY6o7vkkXXDHwMJSU0bc1635N1dkaloUuymnMnP9rw3+Zw14aM
ymyVyGPT1iFRYKU6KGbVaDjNBGz0LRMmliLkZ5ATMRX3qe0rLxtS8q55+GwBPH2A
eV1SknBZ0ghzW+/QmRgVTOSuTwojuccPiREDMNBWhdKquHEdvZLf6g0H7G0n8KXc
EH7qU6mf+vsN4pBHjOj/S7uW2x8TzlfSxEW4GWgAyo7yB3cG5URGs7PQ9ObbUzKa
h/MxliWMLAm06oYdZpLJyyu56qSwy8LseVEM2bNXfcpjFMwXBNNWKO19d2SN4WRz
dCDsjdlPGM+taVZF9Bm+sYfBvRDo7vxtge2IC9uajzqKd/AVxbGvJsXO6KWZgrEg
82bIC6rrrnqvfHRP2moztyKItrDO0qr6bPzMMs8uErnXg53YsB0n40zLnMTuQSw6
pfgKgNljQNwCkimdOPAaYOW1Rb1MAO/cloyfJtCZGas9jNj65rtYwcyNDjEvmlqU
MxR4KlZiagFO3AJBbGkJx9ucqMqt3c1BPi/56v/BoHde+smlnJ+dgEd5ZrstMXNP
1Xapu8GFHJiR92F11CfXZ6sGv4DPk7EUocJDobDG5sfNP/1mDjfAdHYTgu9vVDVj
PI6Z91yyQfArWiHfeBrBQA+e2NOStArflePe7pw9bxVs/NT0ey4Wu/2KzJd+aV/o
FDPzdBDhAk/1hh3QrV2ICYYltO3mWdo6lpXR3r0sdGvGyQKW/nzbsuNyrF9Bq1+/
sAcLXhTAr4w5FnPjVSLUID7NYfvtdcRtYe8RJCjalbnDEcDxvxs378MEpHuckGIV
3VSEdkxQnjDQhB3ErMmuOKtI4//BJJ7MZrgu+m4FAstzjGOmFEq4+XOIkCXl7ce9
aup3oYYpCI1j7oivCnubK9Ae7AZPzHbflnxDl6FyscmC5fyK1pP5fP3ZQQXH9APs
YcEV0oKb2D3BmN0EJBU8cThM6r4oqjLMZsFyJmQSZvRnpFsCp/miBVsJovKUq1U+
FR1e6Iw5E5Xe0eVrqp5v8grOacNKihDKUGu0rKNIRaEZ1jpPq3ezsEtnLO01WsDF
Arj8TKpaO1cb/QavzFnMLKgW0q6yVbE/KwIuEYIYaAj548tZGxIQBnxkLeA2uq0u
mlhEzawkY9fdsIn9nZ7t6ypnsa+n0uimY6IRxHtpGt9NiPvwBFjyyPOwCh3kIj0a
mSe20jZ3NPPIfjQQ84n4s1f/4+7jP6VERHlySRm85pKEWia6zjrWt20FGqb+T13O
zh12LKchJk2Nh/lPfdGl3Q0pWE8iyXLOQ940w+frNXV2Q6jArg6+jNltGMjW/Nbx
+GO1JhkhscZLqnDmM2KUZ06qGVyTAoX3AcDkcqdPrPmRjoxKJRRyk7pFU4ExFucu
zUsneVSEEp/m59BM+pxBaSoFtyK6s47n2wgJPxilvl6b0R0WmR0iGRslGrBmkoz4
sV01C0Cnobkl4qK6OVJZlzwVP4GhXc1KnlU5hrnUl+Y3YYtOxSGh6Oi8MX4jmN4K
efCh/rIWEY1L73xIqfgZJL0RH43NvvGqv4c46cDjT38GsPHZ8TFWL3AcuoHwuFKi
HxgPVXE+zuakZHbHiQTEZDqYBORAl4JMRQiOKAqZoDUcIzfe2Eks1lf858J+Xmtx
WMa80Tux/o09bG+qGsHsiGC7hXFndI/jIm++ddybLS7hTOfKHUge0UA4x9SxIzNu
xmS4QbGtco7qzCIuXVV/+6QIHPJJjOoEr5+5INrxmXiRJT0SO9HUpirVDff4e6Cf
5vX9qWOhv7IJ6Emoy90dUIarHEnyQ4/EPy2+3M48+70wAkWiukXfKDTlpRP6xDtJ
dGOpd+rDkolhwFDdIgHQrZ3wQOw8Y27Aqoh907V/WewGC8MXv5DYHXqYd3T1/LoC
5nz9yKqYVDDTQzg7d3HtoW0tteGG4P+rDve5mTT5CEdQAB7Xk4qMtGrZlFe5cnFc
zl63IY83qKr9tT0lvoHzDYKWl5Eh9qmOCjSMzVa3Z/33QdIg7VRprvo26e2XlN/H
4i98TMaz3jB/XtM27CCfJ+Q+tjdXv68QfWoh/aDeEf+EvfgHpeic5xbgkUl4rW+0
mCN7Ky1K2dWikbszcbV/fI4p2R5696tRVzezwNzmWtMtciVZbtCgWv9nX9n3oMi1
tbr1TSXfs/Ilx/UCcfCumLtG+dKYwL7kVwV53CqfopzZ3jBAJlEPArMGe8OY8ju4
O3/I0tQTGI/Da+GkJACn6WjBRANerRtPO11v5OoJXDSeuK5HaImjwfF7yuBq+7wd
xDlHPJlDpJT9AugSAUZNfuXCaApshiVXg3YF/PxuM22XxeylFYgITImnvXAQfiC2
Fu2hl2XwKxUpCc0ItJ5foicf4YMjfPNHe74qTTojlrGPAhaYNBJaQmBG1oau0Dex
UCjr9+xiP+jeUr/2BG7bc+5THGnKZtGVZjnRahQHN5agTHLkjfoSc5LOdQ4qpMF0
r6zqHoALHIt3+pxCnB3KUODM70uTIvz+MsIVX4b6U9XWbrJVnUeGDx6MO10SDjFS
c+xUTnSxwHuwdOVENSBrFuYqhFRNMtWh7LWBPxaGSJlikPsiRff8YzN+1qU7mQaV
xz8uNkJrAXJagqqRWUy63WBoeCgS5V2FcZUEEdQZDe33IL62D39BUJU9uOL+Q7vB
HeqoL6Uh9NeGKm8yHh7UUEThYDYfQql543tRAlJ900zG2z1+pjNoHmfKAyjiaKg4
DhMfiE9RgpYG1CNo/wPfuZwdB9a2UV6IE2rRU0rM/phJ0QyVuooHn1BGVyCraYwn
UasjY4P+foARUG9U6lPxviYhI/DSbxzLgnCW7rDr+UhqM62AmqT28ZDUSMaLR+Z8
paawUK954UlZ1H7gdDJJk+9BY8nuwqjvX8fnYa9JWDrpTO5Is9/7NgxislVkHn99
lvV0981r6TiOb2U5WChUgV6Q0ziid06XsQW6+PN3/76aL4kdF8qzRf9Wj2NbmB4s
uLsXvesENkUco3wvMCyd1QMT9l9R7hsOA5W9AaQk+vBrFavOBjNhRaC8rxapfjic
JfMBCpkbJL3Jbn/0FyhcbQM0klnia2fz8Ud/Il9S42FPB0qNEekxEBlsS/KwzFAz
FTATb73qSgGwAF+X/2x1Rwzbl6SYeXoH+1kLURyIk5IBTjTWOrqVU0TPhxyMk1Y/
fSNjbJCxnLEIm8PPHBkRwChPew7yzOf7SblWNmEBEJmnbKVjgy207OpEK9hF8t+Z
wB5PzVGXccAylvnyzlve2S4tHGga6t/mByz31KdSyuk9fnE4y1Q827nQI4Hw/JhM
VXQiz7ygjrSYm+qvY+rQTNzgRnWIKOMY9LQDcC0i/gcg8gt4FNibyqe2nrsRcB8s
+FVeoNsEf25Zt/hXROhQoMYlJST13XwqX0ZPT7uX0n2llDOPy1XdelmKGjyjvobb
O4KvjoCljPkwlLh+qWfj80qyNi5SDsHGhBqE/+YYECbE8+inFPUFRhvMz2hzD+k+
nw7fN5WSah/ChJb2QcGLPOBAr+j1E3cfSOIgb775+4h2l7R9eITpZMrjdANHAY/V
F2ZfOOYlmOcqLGeM6a8KvIfiFkhXz4CjWaX6lqH7KuC1/vVG3ayAKCMmTHdEtsK9
tWgPhl6V0gWfhTC9wam1W6KOtmBYUewYGdNkdk+NQ7JQPnTBl04s5ncn+TBX7/G4
nIeogrRI9PSrmlvtzVsI6qM66q8222q7Rjj2aloYH4nuV/3/hSwrE24IGaKoD8i0
PLHMaUki7JJn8RciEdsATFTuB2TIbU16XpK0zvw/GgoefgCcbK3PgIimNWqkbo/x
i0jNT33+nTKoL5dzV/IttSPOCq4q8bguv9IRUDF6Z6yG0rQCBZ1yslfysJW52QTC
/4NcjTKbSUBo1cgXvh6PBCTifq1hWyS3wUVlyBVanpj4Z/SSoxo55eDonpPiGd1x
ZHCNjIkg318xScTnxOvffCQsVzCXQj+Uo6ZHPLOVrafXLp9FIpOzyqLQOf3qvYBv
/sSlbdQYnOtGzpiDg62W1KSah0Y0z7pV2fJ4CPrtSKs+erYRs9w5G+Lvk2wEx97F
0bvaspMmCwaL772hLz/nhilfvyoKwerOwcBtQxXTdzP1SCLi/Sr2toRWriStSHEx
kv1SB76ry76We5/P+FnkU5Vurk7HFLWPnx+dyi4iCEg5KRgDfjQ87yjp/oXZPNy/
ZsX8LnF2Z3zjf0b+BDFs9CD+LbvZg39XQRp8VP/T1Q8a/01XKCrzFjq4yBfQ4dcY
ISby5XUenl6IX0ZVwoAkPmwt8X7vBGmoWcWz3w97XyEp/FsPsgv223tjopt9EPny
blJjVmZYIoM1e0rkh8cLJ+Ku2QCQq2YD2KorI4XAp103jq2EWfSlBHIg2wpsKHfS
6+hY+67VG3bgXIYLF9e5SWXw63wNNpI/DxvB4I+p7HWnWK6P6jjT0jTPJbSp3GB3
sHBOGouRvim0/B0EbuooBRzqa/HFqveOZWl6PCqFi7Bm/veGQbHWQJuL05QYTFds
m3pv6aKVXFwpaMf7hSTNnzUSRInGKrYhEkdnpeRzx2zciu5t1enpNbPTCr2B6Rqv
onEZz9u7yDUFs0vX06nUoyr4Lnc2aNi3egVfz72xw78zbdCI7bGSOhkz7/uopxKD
Bc3tMy5jE9QlhVWx2TDSq318uUFOI5BXF0cZpfFvTvR2badQ0avfD4+MxS4Y+oNo
3IYpDlx4vBaDnNr7PYSnh+JNx3WBIPF7ZfK5P8q0KOXziM2NLX15YsRWBFg061+p
F6uBBNIaGgRFoRxxl3I63ZLqZLlb+xFKzqUxmiaTpb2u7bksQ3/UpqiU9M9bbDtt
lc1rupk3irLTboeRUSDb/DCw+8xexs6Jd0c8fUdXvKyzYi0qCzSR0nZT0jtoIeaG
o4bvModD92phu9nQLcgeglx/CjIW+sd/nN292A50XznfEN6PQEYOy1KTiu+OcqfE
YveyF9zDemstYSjN93CNWEQvVanPV8gFPx502r80B2O8OwNz482zTQe5a9n17NBL
UkcH/BltLxDj02b7kdfQ1IfvH5F10SIBxbSPHWr3JGBdKRsDZmSzcarJAFLPu6f3
NP99JVVvizPZiM2kqR0/eH0IJPo8YqDif1lKFdEmLzSx2Dj9SBI3+70nHeiykfrp
kAjvxtLoo23jezrzFUrqrdhfpDWE4FXM41RkCI0BrcNeKGqEig63AsUvnifmKkdE
Y9kqFKLqsr5bmw3A4V0PKUFGDjZgNZKZ312642yq2UmFo7HoAayyrN2JyKY2yUij
Oi2c8TaLE+TZhAN0NioRIbaTC0x8b4p1GL8w0lxQ49El642NJsxrQJjwjtINOoaY
wz/nKZjIT6yS5Yma50KOs0gvv3bR3ii3UNmLXHGHTH4FmFExpjG+fsA3SUAyNfOw
r3IOY2gc7dxAfbjDz2dAa6Wjyym8v+izboiaeMKGmCZxrvRMpKy1BSpuQJzauyln
WcRkMBuaifHQa076NWQsJ9qbe2QYVH3cKhwwGm8gN2igiAH+klDSuy85WfLZ9UkF
xp99IZB4abyE9HiNReOrJ8NQ6khQ9cImSersU4HewTnNOcxzA1BJy/fxBv0+pOUu
EapsnlA7lZA8mX4RBuiQB6Z9LXAfSUAA9b3zep2flUqXpWiYVnNQqxRGlAXPHaN7
8KOwaLSdou6PkwPEh9Z8uFHGGUjueZctgSorL/v0inqlfKARzp7cCoVJY8vg1nCz
diFVnenxmnBj/st+IkASq+Y/Ruu4JfTK66+P5p26dfBdGtLE4vQ3d0Cg4Uqj6/GY
YpOrZ8G2u1YsnIBg/1sMWmjBDWbQYhRbpt4C4qQl40t3n+PfRZMZgOosn1BbpfIS
mLbS8z5wzcJcrZ4C74RxxogigU8N2VZWJzIuPPqQ+m3qAxvqu3qKNbGZXFcYgIPL
nDfM6MB9ng1zzkbyRHTL1ZWgpZjxr9bRHgm9gzj7bTpDDmsb+c4EHHr5KMC+DfSC
WtaSH2d++hGBxn4vWKJHYzTZPKhchT1IJJWW6iB91CUq7twttB7pBPLfJfvJtiVx
g2spTISkcYtTWIbgek/eZu4OBtfETK0fixWQK0vAbNCUKRDcUeAGPKeRewgExBr6
C2+PRL6ZJJgXjbxEm+cPRZEGM9dkeybEaZOuUpuf/ugBM/8xm+1SGuSGD+wdymmW
saDssJ8A1Xh1vcwCSpjPNIAUEGQSw9llcCh/BV8TO/0oHDtDIYivB6+uhkisBsS+
kgeOw/O0haNbH0/kpDBjrJYLz9lf40urHoaaESiUGmRXiHTIi4fdwjolHCNeRgbL
d3Yn1Jxt2h+6YPcjr8f3KQcih+w1ekrI/v3mDuBe0YkIlyVdPpkroAqVkdGNa0PG
Hdh5yjYFMZlcDS1bS6NhYgCJU6Q8UJcGu6GukHKGNqQmpEIWGbJSUpySje1V4wS1
U//cZ8Ax2MDX9r96V2PUOqIJWms5Wq+1nmUj7pL2gPPmsnkyVrQCw1DY/gmlzhTi
FbmzPAL6wi3cVbFfykOYCR/LxfqFUwEXt1pJ85ZXhfPmg266fru5ZKwh4j1maOqF
syfJplx6TbafUvHM/gMyyASrRpCD5epMqRBhhzcNDB6tz0KvW+z33lBKf2NWj1dq
TrES/BBSqFXbrYpwEZSwtSEoAhTOyanyYmf2PfuWd73bdYbRrhfohhD6C0FS2oUg
uTcH6azQuT0p2Lu6Ux5Aa59BaLXBs+1lc19+IJzax69T+RDdlC6QVAWg7q9AW+N8
Rp0jE3TpYBuqo+3UIUcsFoF2O1Wzgo+7NTI7NINA9ebX1B9YL2+M630+fk44dRvh
Kic4MnYWDwGUPnhdiNcwhzMszuR7ljshohNQXSqQpAA1HNRS0uWArmVneyZ+8863
hcoxYabNQ0WIM2USfgCKTls5V3bASlRZUdnNcwInfS3mK/PJzol6cxPz62yRNcbF
C1RYpLUXHgmRLXFnN8MwuhUooLrYVW38E0kfef/3stpD7y5yBXSpIZO9LkSd9VbZ
adOsPupKc7p6Xl46YvdJjM+yAjVl1wZtl8Vr0IECoWjnljiKR7/cYpZCKiib10Az
Dbau6HlDJ8RKtTxgIMCaNS8eAL4VCWmKUWJDaskyFtPc1Fvv15W3tmpB14s2HdsN
IV5/cXbg8P+JuzhdkSrxdgKA5Nk+h0v/x8f4jwERG6vpsHJt+5VShxYzv+suMgyu
5WRwnaI+OhjaTo8OFY/XWYB41FLrpj1qgIpmH7irhzPdmfhjEOnNd1xJKcalbUG4
vMldnvGES/ePmsO/iWC/aHGEGRiUHVBrWgnRqzqF/uoSNWAjv0YWwC1eeYiwteYb
Jwzm2eFiHUd8Q/v0tRxIfdN9vhLzpdnp8hEpY03pZ8P6lJcNFmu5/ZNHNgLRNs2F
upSNAUu1YOYWSUoCtseThVXwSIYCH40++kzJLagdcRth3n/apM8JMdWNPCUH8JfF
JLTSKt04arVm04IQk5lak89SsxrLR19yPEUjHhngB4PZj60BD2yz1DHvby2zMbIe
vXjVu8TcC+QFJcepctr4pLaoKpsJ7eGpR4Fj1TZUaogsG2PogdmlugrpVlwpkj3R
8hUecLUqYBcBMmH1MSddw6WKfEO9PIT7V+a7qjvI2N1uJ2bGZNy5ttWWpeBIUA9j
IDOqha9IhGZvRVhD3A5CqzDqTEbNvcHwOzDLJD3JRBwCffGRS9DXpLipeM6HiyKr
tjFkrY+N8fi+TVF79TiBNFMPornRIXu2YBp3xuIo7x1vaT56VVhDeX44TO9nZv09
YOz0ZyG/ac8DzZaeqqgIzMRkZQuagnEdEj4eiHoETBpTxrrPkt28WR3l6b4IZjqT
qDdp6voXAQFvPSzfmftDGSW6vxkm89lKBudezFxEycwgBci+vTkNkrsPkM4vE023
06/GU3dC3+DDWruOSdyrQFI48raRtjPP4rzO6dHspWgkq2icbwcp8oEpLA4kEUXz
yti4nXPV4DMB88PIBlHDLZPAcu4dQHYJjpCizIS1uGaY1DXnd+VhDX8CJnC5I2as
x784rc+5b9SubNSXCwU1hJ9GFEpFW5aUBwytH8lDmJfTGZ2h8n4Dw+rrr3Kv/d2O
fAQ0lBJVclDwRH0TrFhS4NSF/oOLxobnQDLrSdxrfdZ4cVuLrNn+XtmE3YOL3etM
wTo4nWzImAWeM98KmmXSiLWv6a45FvdagDf5QOLr4262Oi8s1e13j1dSJT2lcqIr
m3k/xBVtWGFGeHGOCVL7aMs9v9eR/HVoTunBmdVoVF2yvWGfbJJfmiaRvwFqBUMG
8vOQYLVg4vQDd8reTLndavimEVisRnRk26esgoQ6yZtPElYATyjEJGp3103rpAyx
xYwjVdG1OhX+1wEcFFJcDMzKeTILc5R0nsepaiAO4ExVA75zR5+V1USnCbjdJV/k
Qfpq9DX8bLYtAgZerNE8jEoH9F6q76yBUxd3+1UEjtX5NZBxi14dbRi3580T+PyO
1/Bc5SZe8X0gW+18Nhdd6tzRPFVlejZ1XFSmdyadKndSdZsCzAGNk+RdSteYZIW7
vtiVU4SO2Xj0S8iXALs0kVKkSx+Ui/E1cB4WjIMGTsfgoJ5lYWr3b2nHHpHfcWGj
dHECBpuWAtOgTo8L5x0PGvc4tAotLZgSYx7PsuLRDtijMLn41+Cs9eSOic3a1Pxj
Ns9QaiuDPE9Z9S2ZVyWYskhSkEyJTx1UKcAt8Ks1p2cJNyUwLgq4Mg/5ZqkkgYKn
A2oxmHa2MASCorGzkSU6w9O4GYJfO5DGkEodpkh+XMAxjEuzN/ZmpKzbhqQpyXqo
kHYXP8nG8SOhmuXKYTOEMjt67rbvVZdcfaBe27/pDeButsSMiYvhp0EC3V/H+PY2
VPyxIVqG+plSctsn8LjAUOvrzt43J15+7ESDA79Tacrg3CaJ/zBbr6yJLeUU80Oj
Xnr6tIHa4XJqgzY2k+jrWJDu+wyCEpjoP8t1+XvcYHNgtSJNBniOnEPIcg+1Oscj
60Ojp7Zy85quwezHTeJpziE6S5wlcwnprklCTw7nO7RBSKMhIyBSfrgkGZF11lPj
nsZDuPsx94zMUjOfBKB412vRUCZekFQKnIY2C6cvEMA04nx7MSs6oTQgWhwBnFmx
SRYVo+QL3rUip8R7GFZQDshGMDArRdgegih/FLisgmDmW/rFm3c4B6SI2z8qBXEI
M0RZuF03TUlO6CkJe11Oh0k5KJ65OXki4IvWBPMV41NMN/qfrlecT+sVWSiVPA+E
fu6G98RdD2OX+gfWulb4vc7H7Q06RpfboO9f30963k2yJDsEE1KaqaQM2PnVjcfg
P1vlVhr+akv6XHICG4PRO32Ni6H4KTJJdTTvEptH7kSJ1i/x6NoSYG98/DT224J2
Kb0jnZL8GK16Qi/fES8tg7ukjPFF+01YW5q2X/bLdGjhemwTGMOPADExw/QK60F7
oQdIPylftkKo3DF2teSXf5hF5UccZjAsyRz4q0irejIYdI5iAem3Dim37BELzlzp
qT93HPRF3niuPr8ZP79nll9C/1a3LIY0IuKTkOGMNUOdtE1O2pfdBDq788iejxgh
lo5po4vSU5IFdZErggKUk2IswGgsUo6xxjyVLb/6XTLZupry/KnaCTyR5S8kpgTJ
ij84+ti7AMvzCBIdXXeo6TPLjK98Nduw/uFXTeADIkATo8ZRPZWeqBNq/79ueird
N0HDqeAG1NcBfDXl2iPnEOuetWKj3QMa5SKm/dJ/c2rsrpk1ol5ddTub88zRAfa4
ZIQUElW4jYvVExa358RygZKRDknkWkmHkvjK29gEb2x8FAmxc0AELDxUsonzW+3S
1BorfY45eE9V1S99wXLUQj9tk42hvMh6qC0losKXDQpOnWx7AyQTAB4PyU+83DtP
9rTWgF4StndmB/5m8oP5woMVhfsmkUpqHfjiuEchiYkqNwIVEk1AhsJW3VH8hxXa
7+iGG9Am1aSqpNwypAAnAgLvPXyBRFX3jTDk4gfWvGYIGBidFqvziGuoPO2FFgbR
b396/0qdlxJC97X8MN0AcckMZgw11/rDQYBaoYvaYYp2DHnWQs7o3Xu7FCHB7PPO
LdymP37UUfM7TAtDLhmwckJzm/qhekTKXEkxIn7ylPJ5Q3j/rh5FyOUFbWz8HoUB
1NODJsk+CcNGHIZSvSyReniFLnna73ZAlVVP2e0OdHE/p6bolm7YFlNLDtMsEF14
kUPo6ogICnmGVUpG23FkZEtZvyTqeFLqXKCOxSMdeo3zX1WanhLxe/GSNi4mHjdH
oHEvPqPnJmLeo/ulLQJvfGvx2LeYIFk1OzhSuQ2jPapM9lqQ6ENNH/RBK20ZHdFF
oDZt95xohbtnx4FjQGlAq61zmN96NmjGKDeXl5MlnK0wA8PtN/RwNgWcc7zOeR9j
pgjK7YTZlXH6VLxMP9HPMiSsetfprofPqbRhPV5dDamOXRNRZBB+WNKygeoSLcPT
Ic95u+EuoFTQcxhmkrzJk+/+BoEPy1D2GjyZSPeOv8YauNW4ZoScjZ85A9aLdAPb
MPnthYowFRS489LXjNjHK62qE+3FZ6IXAu5eLb8AnmOf0Xcy/aI/pA5/RkOPIi4w
UaLYCJxRdk9SNEYEwgD6gY2rlFPHv+DOodbcxOo7SzXsex7zTtTo41N1OkhbIdqW
XMK5ui4FBeQ/RAJLUjaMPM2v7bRiF7CoOrjocU3jsI2ByxyV5t0lMRR7tX59Kzhk
S82uQRwvZVcJ5OxGZ9ZbAuTBllavNxIB3ipvvxAxoGJ9w2adfgdKKQIwmOX3T4bd
KeIK2HXMoeWYLPuRUUrkqDirBqpWUgbo8+yvUiw2+iElNMmDwQ9UiJiiUiREYPue
h3739RkUcYFCcIWsQ0blnDGsTCU4wRhamptjT+5QbVMDGXKKvv4xJYEenQfZ0+On
SkH1hSaMMUwYcMhubRj0V9oCCgUe5yplg+fAUGWr/2HnC6v+vHa8AIp04dNGO7iF
OEQmikSOIjvNOJOlnUp/RsJGfKTg1kBFLI79cv6IOsyZIY4dz/AX2ygiUH7pWZfL
ylVllZWA8Y3vk34XKJKS8Zsu3ZMmbTMmaKFcBpzys4buZsQj2DG4MBU+/8czPeae
JyKGQuMhsTz9Ldd5+/WdDyhWSP3RVojYl3D5iTatFaZQglsYCT1As38QbcyFVoaM
92lGyFjlNV3r+2EmOZ+EEaLXCoiVOu+JY/HjA/0OELjqdmcOHfEpAjTcAoy5slOH
PRrm2Gm7Z+WgxjfWN2lxYw7rE1hpmoYsbnuVR+gL5ezy4qv+EwSxYw4OSzNs52Zf
Wba/IYnv2BIw11mez/04NXc4BIJm4Vr6T85E0BuFPvXY7eOIc8dfU7evi/EDZJ4G
a06DfRV3u5pR4DXmpmqiGBJs6hm3gsEwzDIAFgPknSUp+8FpouLyzmqvVPJTvQ6n
BlZ86b9Hn/LlEzThI/VTPSj8sjAqid2pvcYqvAlh3MewXuC9oHF07N7LVqd71eOD
TPJYVE4X6lPI0qqKLdxM98/YQkRcHCFKtDZ1k+4Ltjf4naPkfWghoABCMNYiV5a6
DQtGgFnH3HNnRlXxtOc/96fTnyjNKBJf9poxuUr3aFqRH3mk6db52fbLARAn3NpS
Hk/jpIBDA6UOgwSRZWOMWcLFbDtnoGZNISUgZLjsbYtaJrO436sddCLGxJ8K4f9g
rhjgj2eObsXi0f7Kx+6YXtpxiLDhk8s9Uubp3zrBbdkvVLoc2Pq8AYbzvRMSfHKv
qu9ynA9Txingh0g4rzOqwYZKWvsrEYP2hTT1tp0yokeN0Q1DI2Y3YFWwNtEmLyXU
punFysvSUd2/hgLAXzzXz5uh2h8d6DuytAD8v2RtdW0EGIWQHo/dmDxVoZP/wtNz
eH6IzVrO6TgnSmmqEffSgjG+ZK0ek7aj9TQmylgyg0rFTtvQppYXOsqToeR+V3Wu
vbWhurS+Gmw0+/9xI4ApJOmF5/Srerf3POxUHA6bRHpt/55zYYW5gm00Zr/jPhW5
tSZGKO78ZjemogzLvrygOOLhc0YCAPORTFmWc6XGicGDahBGay5v2Lm+91/jOmoO
dTrdcZXkn95oNhU4jiJeX3/54+tPiFtROQP3apgc4My0GsLR31FgjNvIEjq4SUVP
M+9gtnjdp4XzyWc6cn22nZR3Y7VUoPuJ6pDXbg6TQOYzrvN0o28cGFiKmKx/vhhP
3hXJrYa2fSeihQPUrGec2f+MEOwcks5+45K2jUWVGmFynK2Tb1QGCOdAfl6pkA1A
Mnaxub7QVK/GCOCMnQHWZTHXQfBMH8QwxDsgJdT7JvzCU5BpMQbBGVNHwWbUt/h9
a9naJ/MbqebREtUw8pzuWWYjHKI0uMPmVXvwhQsJJf7NbPKJAKESYIX6YSMuza5j
AqeLMrrlhgE3USzWuuI+dO7JpqXOggHfH9xyWWndLkd1th6AxO8+FIhYmHagTquG
VqOQJ5EjxeVZVJbROrVeSa/YdaKZGoqyPZO9f6vEUumlnUzliQDfTHAQu0oySvKH
jec7lCZWCN8rsKMoMslLwnkJXpVMPVesUOin8oueyH9bNMaz/dSx6bNI6/v8fbby
VZKtS1TGk+zEYm2DS3gSblTlLaNDwrwTfkXMudDQta9jlEwYeVprOQwkykVCXt+8
rm2JLVt9yI0bpLvGan15IkZU1KTurQi+9vsP164r2YS49kzEZU9mo7LkP0gkttIl
2QTstVJJNeEJ265Twlxly2PySfAYi9yKsXo6JCfKVhDxxkjd846rXN/la0eiWBH2
OscpSj8NALAJrXo/1ISHwWBxZJ6jX2cHtXAj6VV669jZX4wFdIJMDTSTihOzUnPb
omS4D2d5QXN+Fms3Qpud2Bms7rj4RU1WFT4mj68BWx2jK8UqOxaEuO9fNFvltJGK
OghUsUOcEYCpJOeW49gkV7btfpJPAb7fQAE0OsD53GW+uIF2qSX3+JUDPW8sLYBr
vyHhcru1tW0bJiNXx0mMwXQIAFdoLe06D/u/lnG2TD5G06HK851/xv98LPYswDyh
vGMXZ+LOkjVEf5OZN0JHJmsAxfq1x2fT2bBRwiHM+6suHs6K86hSoyOj8gqH5EIv
CO4aL2pJn+MwW0ESj2DK+qNDei/cG1J1mTXaoDcIECBxI40IdWchh3dUM3Y/9GHf
sXiaUnBVl1um0Dcih8SK1nID2JQFbPdDMuiC26bT6ud2v0OG6HGwUOi7map2uEy9
Okg6Ef9VypF3EwY+IrAxGPdlxrLI+TKrhzPXKN+DD6pnxZTbVztRpjktIssJu9ml
AVpLW53pNAzyafGZoa6Y/qwswn1EoUto1MWzQYXXjdAq9mfXl7Sd6qFxAzDDzxvy
+5wfdWMKOASNzSXT5uhf6MGy+hNXwN9c5103lz+G+zRReSrugRk86SjHPMD8CvbU
a9BUh/uLlx3Vf4XL/sA5E8kBHRY1/KAoIGjWjHEGwH8OeWvNUKA9onDaKXOixU9b
12m8xI1w4BFl93AeocWqHIZtsNNmpWw6nrHLIepBCWSKJWw9UaCMZfsP8jul6MXR
VTAdkIUJY6tJcxu175hwT123yfXIimhNQ5b8T2dlgvMd6VWeazgOKKN2BMSb4gHZ
+3zQmK1D3/kYmmmQhVnWSfKL23UycnGGU/pYEF0C8VACR2zXp5qVnAAoKt38N0Bo
QcNPq/MUYAunBMKRpVTsu7FVv+Fs1bd9UAFUktuwLWiiAJNBSY3PPwvqkcFvsfl4
CeyNTYd9y2HEgRk/nYil806+frwODKxAPPlL8285j1Ms81ssBwfblvMvf68+V4e9
hJxrf1LfE9cXBuNslbXAa1svk5l1PDBANtyd8liQP02IW1vq/CaEZ95WpA4yITsX
EH1MPmjQFcwzPVB7V4IrrA+8F6OzHXAdhIWc2P2RAwQFscpYAlQnr1xrFZJd8kiz
7uboZ4Anl/nHFolD1E+tg/1bnN+C7UKYe/pb71HvDTO1vU3ICs/s1t/J2A2Zphon
OfFaojJlUo8h6yEcswEvSgJgcEenzAi3q2VmdSRS6FLK/j+JryH4Er4NSp3jo3qe
wgdSkOO2O5Up5sT1TMSrhk2+6Yw3UBoW1JKnWpWPkC1KqBbK76a1CInLm9SkT1j6
vGNOuNTYJ3h8tM4SKiqHqFtyvCHe0p5RNmvF5Xt1kZ1zM8ECZBPXae08iPBilzNI
K4dzzkpPiy1O9LYwxfIAtsE067gNRiCsPqIediLo5tFuT7ai+XJ2hlG415OQBGe+
eH8nAag1uDAvAimsZjakoKPxpCI5lNJXug1axTEmDJNvHv7s1U6kg5auwnl7PuZp
9nYaqUnkTd1EgAGpoaMy1XJBg3CVRVY/6seejvYcgEU1NBP5UACDglsrkvOQ+CYW
Hvx5mwOTC+2Aofjm+yac5NjnyVvNOBrVQXo2COUWvAyEvKUDg/kBKGD8kGkauZlT
vIwr5oiSNs+tgcolFCSdPzOV6A83gJrH77URLl0omY8ic+AFsKOY5jsZNjxQJbOC
lmVccj9vLyCBAjceR9cMCmdb1DT+2JJ7mP758LdKId2+FxGXPnABScflDuVRKdFH
uDb1BjHmbS5tUPxiz809cAVUXcCC3jgxYla2QQ6N5Cu9Nu0yATfSvDAaHX0gdfwx
gvyNorVEWJsFty8ciYdXosG6HZfZPgehlxOh4T2BaVYP9wnpq989JLcFpu1Ivrfa
WF9dIRoUvFK66m5p8ij6FcVle9X55uIz/u9qxfssyj5jEpZtWOW+5csqFyrBwsQv
RQYGl0+mm3wx6tdsk4VAU7DbuJorF4qE7dlitrAioeVqLMr4YRWeS6ZVv89yoA99
S2RWray7ZQbEkfDlqbg3jneXcQE8qR20DCH3W0i/zoVf1UILi+nDg5xYrBMctjAB
eSLxfHMFRdRljD0u1sFuPFNCapErXiG/s3P5vF0qadEHudtC17jaJpVd7lpfCgRU
fmwvv+lF8AjH4LlcJQl0af8Xg1HPy9Xs2gTim1qFLWvLm4dMOtM7gt97hysZ/YSj
qpvQtdF9npnDFIEn/gFmGEdYT+An0gHncgloCkU2i35Rx8J8RmGYbSKDyN/sRjoN
9QHKTNdCoMr9fQdaZ4bqFgtpiNQ3uXQ4TdB93fwi5aONX23k8CNEwqsD7Tl8+ipH
X0Ypg+Sbz3x418t84Zg/2AFizY+vBem0nt2fKkbnuI8J9NbRv2YM9QgM5suGHmCQ
Bu42FxfFBwEM28cxZnwPLl0sOJ6YO0mBnbYJnBxm8MHnvLID4c84ivsGLaA83zdO
EP4ig04ZTDYsAHjzTVkbxSVS0MI/i6cQrx11tf/oFp+UZDk5KzcGlv6foH8WKNyo
3/w8clxlSvkZHAq7S1qKPvI0kGaRBOsGP7VrL3Na1FxVOX0cHDk8tLMoy2zLJj+D
yUaZRHHdCmMADymZ7ie5u/7hSeenc2bdyWTao9NiFAV5wn+vvOLrsLPh4CtGbnNS
R84ACSPNKRhNEIsFNv+NFC8wIrO3QoX6Kb6hYaKLAz03hBI2hvZBzK2oL7Tstq0j
cawf5UAL7Mw/g34OwLDJzskIXE6tlMInMF9w67RYJ1YjeORqRCYV3blCViatQVj/
VXej0YrvmIg8ata03nKB6dbX3JzGOc66zTt1UM/EortBbeQ9lATkPb0Me/t/CbCR
/SHGGGOfNIzfRap8DXRrkJjh5SmvqCblzZ4C81xNz5fEywBJ1CmmT1PG3XoOazXy
+kAkHWkEBRMQwF4tUCc0kdE5Q8xBEnXLO8Hm+TVG9iHcbfFigPgv8Y07id4DEMdz
VDhGfiHP50ln9a3dybU4Y+0JIkXFRNLDVI+lKZFJTBGoMDzUH0vd+ZqAB6PnkzO0
rpyZSC/QfFgqUQSTgJ3x2mbOUEHBgwzApkTqIhUoT4tYoVocYPfP3PwqPazammt9
ijUk7PimGAVtamYnSx86ILYixPeHEFOSr9eDhnUj8ik6kwUe8UfvPmnlJ5JvwFUX
sYpvX3+yjEo3PwJAD9rB2XTQVj4YOqTwuFkoCSNSljfW8P+8BTQZ+RdgJpLQvzQ0
WsqyXdh+2iZunY8ubwGCKDtnS7IUr174mREnQJixGj8DRiJSNVK/VVrx9cj8BZnX
8wuQQ1s9JcZumhd75auBv34FWuwu7F0f8QgNc7iCCNtMKiu3NmkkK8GfeJpj71Ev
dCFIlemFiSka1ndH9Fb9kmi5MbzMMXSNOc/xiR1xV0xPFjSstMfuU7qGHiUhgOX3
WshMj9gVgRkR8QyWwpbrZ9qO6teXgs2DeKqn1z3jJCFEVqaWwv1bIcszsDO12xRW
vjKBSucotKbaKQEx4qM2R/A+4qbxYTD49djoXnukbROshIrPVxmM7BaDl7EcLkYY
OACGtQiBOo3rSwNmLhh8Boz+dtcIHtZxriSAhTt1/klN6k2BNITJeiPIDckQ+QIh
CCLKFadxR0An//dDvhihoBtZgRfG/smXKaMKibuidKKvQ9KRLcEgTKdThIoHekgr
p1WQ7OZlPnVuvPRJmL4h+ZMpGMXAusxXYOqT6m/2wR3qM9sNXLnU6vg/dnt/S0x8
w/cFnGJrjQdabkjEp3nmAQvZ/zDlvi4EyS0le1Kxng8uujWY5z5HORNtOvSSi1Zl
NRUInXbTgVW7GdcKmlXnPwkkHSPi08bvaUYv3sOO4a6v2yjbYWkiMb1xpkPvBMiJ
YAQdq/Lq/myrxl8LCNcDr8+Jnb8ZhXXi8x8M+TTE31blRGECIQ32HSY086zA16v4
ldtNLFfKN/PANXjMNX0eWExjtXMbhtY9v3KQeS0N0OZphOiPm5zY5dyGa4uDX5Xm
G4rpb6nHK9SHuvIxA0lnE31B/+A+FAb3BUw3j4sgHZ6Ki2qEVdys/wTI5oAFQzYU
auk1UCdB88w6QZJZAXx6EzepspLCzL5pz8O5Zp30YEozLeDnrBSXjBZeqKyjSyS/
u2SRYTd42LNe6h1N1QKbZdzxuTT9qB/G431sAPpscts4iV1MDV99i4/80sJuROgb
c/X817n+PI7Xr3Z6OzYfukJ72HIbvhXH1PWW23tDfAnseU5HEcq1vsSAsUTvQqR3
pKiDmlkbFBz7ydo2H99F9XKxz92k9uG3oArPgRFGPTE1ggXfcHL2ATqym2WKjpO7
5AsTendB7gP3ZVFObdng0b+38iGA4LLF1apqdme6UtzMUdnVzZdQ1XYmBvTxQICF
W9JCSa+3Xvqz6UnPOUfIKn1EM8YmTaL0ad5CpZ0I2KgsD2ne0cbqQYqxKjW2LzLi
Ov/2Hsew9HTqsbbCK2T2D6SVi+P7D7xaw9nm1uBvHL/ttA/hZZFbawHcXdQZCftZ
Ks81I4usrRwO9HGoOB43MpYwvq4Z5U8BYhnhMcT8amfrkF+BQjWv7JYVna+wA2z2
oncmrQo9AN7bwFmBM3fpcmloY/Vxm05f13igrit7Du5zRuMY1QcLGppBA7CXysgP
M9Dj0LwzHdVe5k5sJ+BafZjkcHjFpJye4lsVK7syeHj2oJANzcpm3ZHW8JK+ZZ2C
36kubq728vkc+6xfZrL7p7K3/l+9B+T8p9pZrLVQvCZoZIErG2Yo3eSP0Qf1upoL
+5hojX0GefV6Vt30d6SIr+J+8ZtKALYvCZen75cAjCw3YGmV0Qymsvf5HDeXw6Fe
rwVTKeqKOBUsl8/W2X9OK0ftXxm0INYNDWfQwTx2CY+pMVwAR/SRrr3cXlWhiRn3
fNJqd88o6bk/vuhiUThdjX/lxlv1kOkCqAIERMlEC6P7AyFKD8hC2+b47zdz9NiS
U0X5EFGuPBf9O34vZAm/RdpU16rD2vbGv/3e58oIR57v+FAhCqB2A1zTaGmcPej9
SrmnlEBU2LmZCgmwCcNCv3vRIx9xBJo4L+6HU1ficp/9nl5CCGeztAlFcuYR//Vr
7Hzv5dqTD2iCVR5/XlvRkRgGTq5gorCC7eY5doY2I6lrh9iNGCz8q/hTZqvaecNv
vtMUS8NEA1YEEw0BB7H9oPPBwji+IPRkC4pN2Vf+w8IsC2rA34oib7SVl7T8EMt1
ri+cSoGff/weRPq6qDrVKBMwryjU+jic0VUbL9zr7XiKRs+bBih226175n0YR6sh
y/l4WqPBj0NI202BnxVq9T6h+jeEdvNK+s/YdkcJ0/b0sNxMe50N78FlINx0kuOm
E/ym4L0zoKfQDEP8Wbte1A8OIRmUA49IA1Z3zznDqjSTZMxM/BQl3jBj8BJxMCXQ
W3+9AjlbHwOZ5Tq6lP9+3KPTpUf6L8U++oQcLN9OC298k9GGEXGTkrAC2YXUVTnJ
FYMO3xWV6B9NsHSwegP4tXMjyvYFabBezQjJCPuhTCS6hUTuT9mRqDuD/ubSh5Jq
3nobQGXhqEd+D863S5oL1qm2CVvAiyhOCAhVyD7fwuRcjhN7i/B9Y+RKGQPIrDm/
DWW/UCArmSdhuVxRcG3e2l20yAJF+B+Sf63j2K/OFjA3AODpil0f6YF9NF/bfaoB
OoTvPOBSMvO6byzMqOTavnhaELCezba9NE3abxzyNm19fLRvFKbgScO9tNNy/1pw
5gRfMdbh+2yygDuwIdFbUB0pxTh1ZCAmUni9BGS/rGBiPFtK4P1mj20m5rISAcJ+
TWtcchB7JUBkUekBCX+6LGy4sbR6p7l80l9FlCAVQvPejhmKNCzQsSsaFADusTv8
2kQ6rCTzD2mMu3EOTzak3HedypMdgS7IeueEQayXfUFUUbcltGX84FJ9gEcIv0i1
Ax+nyq69qRimAUn876G2uTq6S5rPcVNc6fI7JCfUd65XW/CNqodQ3tdpWsSbY+5e
/YekC2EIVT9NXxhRBFYfQE7PcbsefYHYNNxs0liS+xl6a6muHgFqdZuSXomzbiQC
O6EJUE/3eEvtuPyQJBS130EujFY9oG5h2jbK0fjll9u30H8PFrp4LWK59fyL/ePz
UyfxjKzDLt02LCTe3W6M0CMCBUP1byMC+EcwArad4Vgm8J3u5++4EaAASpN2CYHf
t4GLsKB6ibi8saFqCjFgHDGTzFZdAKnNv5IHI7QIVkvqNvwgCyxsGTS4sDQ/KmLM
IwgMw5uO5d5IFAAS1dr7cUzu0wWVkLb9+QOWEE8nFQgs0uEx3Zj/kjzFeGwz6M09
BD3QwlRal/a41JcrRzAOHjLDlYA/i6Z8gSWczB1LFBbi2yyR7laa82BuFKABAHfs
HCPxZ/ecJP+bPn84ATRU/TF8OIMP9h44UlRaGpZ5svgLIVXKs6kYD7qV6XhIkw7o
qMRs0mIBvjt8cmtGCwyQ2kIfEo58k4WXm6tpgi53XM0z37xkx6rvF+q2gGTHBIp4
WTvcs8vIMf+7fq587gFvhtWCdYqHbAZ+PtOcLVTvAWUXAZmaNJNshqRW9Ei5hpwP
XT4vSEOiYL8C18XfcTOcJyVjMlml4gP79yqV1Oo/ALWyDC3k9b1kKzzELtqD/rmp
nUgMZspkK5ztHjuMBgAoYW63w3jdCHH+ph4s1BPFG79YMVtNvEMIqNg4fn+yQEew
U0oEWWAffs4SW2lAmESDrX2LXYikFQLTORPaUBvU+QWXyi4J+rQBX1CdJGGANcH8
5uE35XSDeR6kvX422EPz9AmqJ2smR8sQPRW1UZc4ixH9ZyvmzWhmGhofprbkZpuC
kBjVFvGAdBWu2UdW5p6+2hbboJpOzLbznu5BWctVj9ZcCMHp6Bh72JK3+wF3WtnI
kQakCWrLCtWJhTLSKfpw7mv9r62SCjryWExbchPrOB2o4DFNIs9UVaUO6orpAftF
cfizsUs0BvMGAHDnjAnGS31P+XJ5bLlR6DnyJBan4Xo0mjBn47pqwsNoPHSIzfco
mDqWCVBLUPqlF1F7SWdmZJDVHuISK+M3WSZT395LigHe0WQeToy0XPtK4lgk/ZXK
5ONPLYY/GOzccr3EpacLyDeX0q9OBCjx3i0JjmxcIxmCllM3tXmkUoyQJ9DVP0bU
8EeMdBEDbNVEurkgS79VEFWEsVVr09aLhGdEPQn4o9gwzFL8ebRvBkR/fewf/SDg
urPNMXW1sUHX8azSWHlICiV5NlJ8/ubRsODmW2BwT7exEQliK+KOjwZV0MR79ooU
+1nSsamokpofGPAqlHY4vPQBAbKJXEPTv+JyQsY9hLBOmR1JVYjlMm6fsaQJ9WcL
9WrcyFoBltJb40NMTr8yU4668CYtX8iwxlR/EjdzS8Mpz1l1T1TpIYB89Gt9gwkO
QfVmmb3zL1aU91t+1plmTnHvBAr/jUja9iBAhHnf1/Ra3awfIXiUpPpfXCBaBkBJ
raa0opMiNoXHpIfUCQr7kJIhS+YueHA/oprQT2/AL8MxcD1i9/+uj1FHD7yG5SCw
njM1mK6SvtAX9pqO4VXj/ezqeA6wV/v/9QnHNf3moKAEjaivTxpi1zkmEMeWVZMG
OrW/6i8moT3bWuaFhzH0yhX2v95fO9Dv3VEHtR+YQPAfWv5DOiUqMDdc4IF6oCqr
n1U+2FUkEYV/b7cRc9xOkBmH4zb2L2myYd2MVGrk2HxoL37oop6aF4WzR2HEapmQ
Z5sNS7Cswq76p77adLJl6c5jDnGIrJHd3rOnARu3N/VC5qaixtvNOP8S2BtsJN+l
fo2eQ3G44OTfvbfR5+Uc0Z1mjIXQZ9lFvAZtPgfEkz1DbnR7AVuCaXNx0jraYoc/
wJA5XxwvmG7A+d4dFA4zpq00cTPs7/qOFaMiWUKOoOZ9LTH898c20b3fSfwaf28y
GSN4l1wteYXm3M3TbmnaI+ITQFS6HXeAXgbsT3orlI1+MlDq+1K+z7tVie4TQBEC
86J1lwX00EBcq1+3D3ob9lZFhKyUYzFOWih77y7G5PRDyHoX1FDgfQe/2uKacRjd
sZb+yHygSicLmOkV8jPp4GaeSUa2uVZzjRoTkXT97v1xFWXdbrCsODbkHpjTMDuD
eeg//SVTqVN5V8SlmCZW7uEmnlykU8i53MavIYyIMWzx8R776vySDsPTtM4FES5v
BKS+Hp8wqaOljLq0uGsnpceYHHHkGR9aZl3RGW3xtJvVfVHgfmJuegDNfA5WbQ3M
hBGxHna3bPXWsws+0Bp9WVepgr88fdUbDGHesnivhJqPHGNaHdSGhHujkyV+UGtl
O9FhIU08CEZT7nD2QOGrOV00eX9C+3TMfW8sAAIGrkECdNLvyK0dArAcSBqMDGxF
erbgggyZ/C/+EQLFzkillvgGHFKBxCYHaHfVnefpBA/VYNluoKU5sTuyRMXV2I1v
vqC55V7MPe1DsEKlLHz5RX/amoSap0ujm1YfGPz6gbq0BLWmwm5D+6yc98Mtic3u
wIm/D7LO8mlYzfwC8B0qPQxqVKFHY9bq071tWwWFytflR0S/0Ry/MLdOmXX8X2em
TRWo5wDHoXNx5/46un2TeITbhuLVR79gS27k/UESHylNi6xP8trgcgUwyoLE+tX4
8qA7muU4siUCmC33yAoLQDHWzxXEYxlRo5pCxyhgrHsmgTqODkNvLhEIstkIdC/R
w+9fN9gedCt4K4zTBDt0nWQkqwm98p0PG7DhT6ifdKVqKDVukmBa3aYZldRygG+k
o+dvZkS9K6fbabVdsqLjH3LStw8i65bUBk4XB36uk+C/V1n2weRczRhcBZkiYQ3y
V3bPs/QCtIB2Nc86wj2zOvwprViqGFTTyJ1hmxFDN/n+dLBmexEOR6onz8NxuVoG
9MnvAYiQBWBpCKgiojaezl2VKHHIeGwf401UGUV23Uqh6LDOhiFaN2xWGcSHP3+/
1JrRKGu8cXtTGKZ9NHIrOog+pAufrH1oIuNdtIBr3K0z6gJVOXMQ0SMigWRGL0Fs
3jdZum0wbQbUv92tfYZSf8fDKKN9KAbub4fTrTZVUVBl2Vqm3+2Gckv1q1DrdhXp
VdmuTZ7uTzpbwQCEjGwkCPmrFhZYhzP9Fq5/MRjjeCJmChQRZPUbGeXes3u/a9v0
ZaRp1Cr5bkFXbFfuSBBySiJ0jHwvzkBOSrlDcHzYHRJfvlUF+8Uszw22zbOKOzdZ
OvoZ1zQNKgDQ2B3JN9f3/nvZQHXMhO335iIaRfciKNkyhC8VffbFFg8cXOOnSwNn
CJwS5z4iz4E+VKRR6BO+hJzbegcnjgBU1f/Q5jb4gDxDCU44naaZqldEgUl9tvNo
c4QJ2Ze1qbA8FCVQByImTm0eGr5cbLtBgqIYBSsPKMdjD1Dg+xiiaUPmb4yXzU68
F5ckaN4OfBCXO4uX0bw2l6NS6bTuIkx8Xr5XnvTwGFcPMjv0zr0D30gtRFp9en9h
s8qBDSBA5n8gFwoum9lBlmHiQy29Ds4hixbksfbEMXGTeMgkopFW+AKiznyvzt3N
kYLH4oNirezzzyEikKhmKlsqJjLjCba8+jj8wkCC4cjwQ/uCEjA5q5eu8sogcofI
dWbFUQ4O+1pSryY0I1f4UTZ/7RPtyPX6BA7SUC++F3Wv3IakKxOG9KBG707fAfPH
uY4CiNEQYqKqgYzCAeWJF9QNUvNhTefut7UObpXzp4Yl46tkzZWQYq9hHjL6eS3+
SUm0xqkujhSknLFeKUrfa+JjZKuM3bP8JUDdST97KfAMWc/0auGDmu2Bmn0ASUNz
UPP8VPyp5Mf+tHgD/9oD83dPNEyTNtYakUhnunHe8FWg1FM6V6oAds3tsE+b3Sdz
Vo+3huPeZf+lHfRMLRmtD74IeKWp2PnxymWop/B+HP6df225bV/CfW5kWXPy/oup
iBOR5hyNX6OdtmEWRbdoRYJwDzo1sdm1qtygso6cPoNWG5fS5eRd/HawKJPib8SJ
BBlflsO6HS7qekpBe3rdLyw4u+ITIh2Mk1/LBbw9TDVwHHIoVN++pBG1Tnv1EDYD
mft9xnXg5mMAOivDEuo/uBMxTFrLhHR/z7CgaGz70PbAKiv9G/wCSF/M9kqMuWPo
fVGdMQ7QKpwMHCPiaT/+/wdKYVfXmH3vHYf0O2uFKWJibblj2Kx2nA819xuhWrWS
ZpkiLjMd7UH3oqmAaxLTsulSzK7CSfqryTp4Mh8pfpn0NHT3VeYiHRBiP0vQyTS4
41OG+ttM9jDZb9t6Q2BvVDTdDbJ404wV6QAvH2IX0AEYDctviox2dLQSncaDJt99
xTbxUsUBXc1fx1LtLRYPsiMumuBDjGUf0UcBpUatibpAyt4CaW0J6zjOK3YydjCS
XSMNhdRzrVbPoIidDnHN+GU7SCLisYN7zzC7Gdy773OodkgUmfBeCdoDNBHcKNj+
jeUygdkmdc2EgJBpikuMwEl8Ww5dMWGpodnFrWvkmaRIDQSHAFok3zmoDky1hbXY
QKdbU+YXr35IxodzR80R0dSl1Ukb/OIY+EKVFk0vin0Go+gICEqmYuDxwIbTCuDa
QqkUj5J4fJPuFhanuwBIZOGF27gOpCIuJg7e4iO93kKCAzrFXYHDMnRhXaZaEQb0
VMNV7Ug3wcqvterYXQK3M7uQUIfoXcCDxv33j7mi/GEcwdWBTnp2TKaHkOAZEofN
Ffx2aPoI6lh0mR1FugTy1fzgZAz5j1n3v6Uqio0Do/gdZDlLG7Z2gp/31GSnZMe7
pkTBYGCehDr0AtZUweGYowBAO+jRmIp8o1mqgFKOzk4HTHRlYFFTDHOExdgSuc/B
whyR1BZSj1wJ9e7ZDQzuf0Qi5Jpkb9QKV5R4I2Ud4FAAc/eIVwtmRIusZZYxFrJf
iOUYAKYw+Qeskn6iwBwqRbGtgmnbozTYbApv/NWk9dHY0O9Rvae5Vsw0VUEv7sNq
c5F3kvoVaraGdQOyl36DAxh1GL//hOnVz3xpLKqz1cnZrZhpf/QdBj9zooSaiPKz
pJcojjidOF7JCSLQ+t+5wHtmUomYhgr9Qcfm/tSJaL3447F+kYLWS1mD3pip2qZE
/ZFEIlLKHtdCPTDz141Vug2EApst89aJZpQhp3OptViDpYQkikD3p3SL01cYqS+2
82bJgMEPTSOUrpGqY5v1Y7yOf4ZiUp2QdbOCLQjQJZU1BTIYlI40YR6NPojKGj9q
OmtZFyD1mF/8o+J0PUp42gQdxvnkb8M20eXrSk476JBcErwUN0FbQmJN2xHXYV08
Eva7N5WH5xC9WZQJVDmydn8imFNArCMPZbEZljqtsB//jxeaRhMCxMs/pDXoMIFz
dtLfpoBmivpAmzehVKhuyTCoFy66XYD1NLoVlQGouXEDzGk1hIgjnw/3wE0eQ1Bi
ej/PGF8iX2RieW6fd3hKbCUEMvFDtQ/jhWBFOOWTgdiFRXdns/EcaaQUyn3QqOmK
eaNNGoKk1jpEy/BeN74T1lBH6VvcLvGfkPuUAA/kKJedTqVw+SYgQR34W+gQw6Al
FO/+MDMRpQglKlaoy0nwAGMqlbdR0h7C0XIhfglFB/e5Ks0Ra2zagA8XW8+sThtX
P2Nd2GcoCvy1ZQSRkvc21k2S3hFAc1BWy+0VRKBWKssmPkMsrKpF4pRj+em6lAHo
r31NEqf4faCbT4o5tPr5KKm8S+ebNAvK7To6D7nXyoMIrqx4Gg3TxT65ERY8KmxK
/kwnb24M3HHgZ4omo3FUfDMWVdUqVWxpdn/SNGwUFexjCXEjmu/XkyHJZ4hMn+rJ
U4tLszDZCcQ5rs0Xp63DraJGdmYFsWWGYC4wtfcMu8D1KtTtJEntj0g5EPJCsRwC
I1qO2jH9CfLEtrptlpbi9wz+HxnmXu0ZcfLZzjM7uq23m4dFFHqqK3Ewb2Or2jIq
+DjvRdZe8D+UQsdIokGm1BGVq5pHx2M5Nl35ERsiujXM6qRXHGRTvSzzSXQWgpKZ
8wd9Y9opu1YQ2CZ4VxVOpHECHPwRqrdD5r4rJTz/P6EGVJyAk4D1jLQWZxafWVUq
U7IiB/pYZN1s6G0Bq2qSqH8W58Lrg80Yw2Grdx5Kqmhd7kKuiAuDfsYr7UatOhdS
2vcunw7NDN7/nk7OEKT3V5bAtkKCvJ0LiCq1xHwTj8Wp9yHzSj7jIha4Og86CAQA
DgVQ166XsH40fUkFSc64dMZ/d7atiwWHMuuZznWtQZOaqtsp/MGaF5hmsICmxgej
eOjLtisx/lvwiNPq9bui6eV9LHM9jHgACUE2FPh80+XYQnBPwXTRJSSOe8vaokAb
eAG0mZK62+/R/Z6wrEMaoyqrWDIX6poE/W37zcOonvVwkHyZ7qaK/rRZrsorWomN
Z4Rmrn9YY4pgp9NUGKsGLTAcHMlC17o2X/PtOZo3hyDKcn68kTi0G/ZUdMw6f91E
DECMRkrO5AbunLxrbTLZKTePc9Yasv1gSka9ryquDDH64y/aBF5ngrkDOoS6EjVy
yS3p6+MasUfWmM/DxPuMnCz5nko0gSftMevP+/9ABXIPLWvQ99L6WRK0BOiiMPSZ
88D1JJ5yL1bglouH7dkmu6bG02S2O8LnUNXNDM0dPo7j/aAhFswyHHRxIwD3pE8L
8oteIBRu/GlQmE60sgAmGoo71QXaHI8dgErzg/SPV4e6s78uA0qZ+gCSDZKr0pkS
u5Myjxnn+rY/PX1n98PpW7HvtqJ/dV1qWmdPVnVEFdAGpiQuNd8DZiT1HtdRVcFw
ntMGZgSO9JLKemEZ62M5iXcP1cb/xx+ygN8Ah7ZoV8OMv0k8FQbtUsp5k3l5KWfb
aid9gw/akMFMxYKnQ/W51G1U4DNyoRvJZ3ef4AASUlnnybqIuwy7wgf6BfFq6a6m
6sbXISLZAqdjFqz6qR83vhl1n1QJWvfddQii1jSFNk709fYVbYB1Z2yVfl719H9e
bp6lhLNwIVfwCP/q0Xx5+bK3piqXAbCJpFOAnjNMkwTw7+HavGu+y4X/zePav3F1
IYtS9uJwmGcWN+cgkcKBB3YJfOJoHzrH1Hck+Ka28NRtWWwVlXyyhb6O1+YqhTA7
OZOeZ3j6JfLyXbUa+lsTTl6lUvHx+sGFvEzdcK1gdY9f7fcXvsui8oq0cHSzFPUw
KNyWzwA4VW/h/wvmOXQ+ATRzY2EfpivdCibSB0ZympGeLQjNhk5+AJZXtMz76fbL
qn+MOg9TXksb9E+H4/tgtJ+AgzF7ziy4M09zVFsDWnfDqvMxE4SaIHTzr1ZOhwVb
8B8IinDyCPdgs1+g5v44OppfqS8WGZFgyoWxGscRg1MlR+ZlpukQQNJT4ZAbrCmx
EyD+AXtCHbFf+Pw6q4FqF3jP1tLcI39M2QqxZ+6iFWgpq9UIQkTRb+hATmuaReDC
l7oechVioMtwdBqByP0FBXxU2jn15tv5grMSqSlP0SYoYEP3ZrQqa4S/rlfmmPf6
G+UukIVuImNqXzp1bsWVMGBnGgolZYiey8obN7Luc04l2pOQ/KEwuv1YS6sbnDoS
z4Vh9w/h5j/ARiOVw4d4aGZ/j28ZrSDoPu3DMFrVWYAvE3k/16sikLge1rgIaUse
ajkPj+d+6hvEw8Q02sLmvSJqPM1vB/nSGzztk0Vjx6PDzUp8cT2V6ZngOTDhel3S
TyMnt/FF5rOO3rF+0cbE/A0rAwrEyLlc+CihsQM0OH3MwGf2XxWSDmjBmUQjyHie
zLZ56oPtIDGgf3WdplLIxmPXM5Vxg7n5z0Ar8r23oZI+Ca5hSvgrktGaZxe/e+3w
MQCvrKYdnCFHa4U4U1sKIUUptYwwc/LLRSr9E8JYYHOWdiRKsKlrJdlXq7eodfkG
KizVBk4gxegItclGp8tHNjs4q1EVwKhjw5c4HCcKHYUO1kSgvjQuGh0F1gDUXSiY
1zy7dlXt25g4DCaOObQKncFQo4QoGtEBSeZYpBjZOV5F/R0cXJ5b96mRb5MbgK2R
1Or8mUrKq0VP01H4qZYHQ4hS3a0W3Zy8fnYuBo+uqPo5+BEamoaMfyc4Qr7RIAlT
ERyzym3pkLCSjThQAlltPXWlLh9hsySrh6eNKqZyP9H/fSEKQoQH6fLlZsS4Zu/+
X3aWmTB/SbcTdEOoZC4B0Tj7qtynXwFu0BXAtghHj+NBDDZrGm9wBx+wjiYn1RDq
cXnRn+gdivPT5/nkSbyusndoQjdGAZ8a2nVpVT2zFWzPN2T3PYfIpyTTB6Py/x+B
ZajlU3a+XKWAG/gHMCgJGPOix5zsojN8o5TAMLvx64qmW+WWKCTsMPX8YvwzBMQy
u4QFK69pYLkss69iuFSIpV3Hp3BGj9Lx3WL+ZeeXoq3OZ8WoXkHjMtTgJ4HXg950
4/r/2jWOBwcAmAjTAawaZS0kXU+x65ZPHx4cDh/9BjGa+HOBvjQANAqc4AUzah9Q
Q+JXBvGHlEMorXGJlY53yEKB23uEMYm64sI9vlGr2/6UJ2XpEwnjvHHD8KbwUzul
q7l33jazXaQhgwCR5MG2ddw8j/+UVQJYf+BkUmrs/WvEtvv1S0xNkvwI5leCboDY
pn8tBchhowdxOLNOc8wQGkw97YYiXs6HJb3pAo/R0ujQf6NiHaqFPd4nQOWrQuZX
KncCMoCmCBryk6QPnRmvAy+tbDj7nP17JWw6c956vtddGJoNvwxAdAbNENZUdT2q
5sYFqtWAkgTo91Qbb/5x9hTCCyl832SsvrScYKGnZVi3acpTS7Q7wHW9PJgJhbzG
ANHPXVFfIjLUvuCr56bBFA7OTZaluwRpLZmm4k0fIYL4wEu+WJJYZAclLjDRYCeG
MgFp4eGkNNBMHpc4uA9yGMDrL7S8n1kJLjdYd5ViYtsgvvtTyRTFX6qRaGTJyQsj
SU/xO5f1DWOBhQPWD/DjqM8QIzlLQLYCiKEBhZg4Ej5iv8yhy3ZgOcIw3u+USJ7z
BucUdpkUNAwfLLztixIsa1nG4SKLMAlTbdi56iv0BM3bD9yo47VTKQ3azkMlIryV
O8PoDp3f6kVlDH2wc0ngI2OsqkmSBhw33K4hHPcHDQSYCHejxawHu/LRxItK/WDv
QOjVwRfTS3n/BBm3wFElIdtdjErfAdhZU3RqnoW27skPFGs8pMR0iLuBV0r/+YuV
rgiBFDcTLdv0kSzftunb7iC3KN15D3in10x7ALFTA47kxMFDmuDxemNOZmg3TcnO
3ECdPWHpJrmHbVRB+zOVF5WHeQV4qO1W7cGbQ0AZO3ZGYgG8g3LbHBAfdOUV+rvI
761yypMy9MJ1AK8QPIq4HPtg4ESxstbWBOagljvEFhgPrf3Jxc+wvwztVTx85a58
6qhkjYQUUveD6JkTIERGdfs5awxxe7uE4SIAX6pwMFtmQIktbtR8Hk5q5KMgZSU2
ZVGP7vZFed6Cm3QLGaBkUBZAFR2HZ9Yx1amoVeQB1dLqciOEa9yDSb1NbMNStb8M
qbmOsVV88/kBbS6zFayhQniQz0h83/CYeekFPCM9xzqlWxRPJsD3ed5ZplwP6tC4
tk0zfmFVGW1hTtExSGbMPUrl00roircl0nv3EqElg8J6+li1z3BBLnA/7cyik2LT
cX8B6mz3gfKZUMOdxib7VSv2jgl7ZsC+Zs9EHKPiAEdgCFo6ilENzQNWGaRLsUuL
5wABf8Re8JQHPSVitunQzw0EfNxb+Vcnh5G4X9BuJ7uAaFwWhKUfpnAmKFMGbT0S
vL6yRljzDGiVsSXyGfBB32cFT3NVtrGI+OL88SNlKp4fUnzjc2u2M8NyB5kireFD
BNl7IbFF4RUrIfNjh9THtiv7SrRChjqUkPbTALSAE2E7Kwrv/Are23J/OriKK5py
ckv03ecKB2CxdSLoYvGisoZBhxaLAfNvrVq+EZzgjCJ+hYXemV7DzEC6guqU4prm
NT4G+EtHl9L9eysHw5k64H9BdMKkEPRWELBNQalNdQwizE6/+ZPlsBijTGJC3XCG
hJH8uOs4IFvVQihKIHMic8N0lIg6K9N5o72s44q5J9YDvO54P/k43L1lb2lCtcpc
B3P6ig9SZGqiQrtwaNf3GDCt/QMdsO+RXzPOdcfO6haTCKnBAxmF8fIxRGXGl5N+
hHAU1QoiKNdsyv3AETjJrpm1ORr3GWdGY3CfSkzZQwrvw+490dk5A6akqRiqylw9
ujGIaKG+j8JDsGQAo2j0uG41c9f3uuBBVJd20iIrIgKD9EIi0oGjtBefaXYTct3N
SnoVb8SaCaYgbKr9RPP3k7IP4vtgaeK4ppI/leStUWZa1sCSzincqfejOkYqcI88
VVqNooKPC1JIYYz+O9fwKn8YYxnX4o2nkY2K4zHSpuXJ8a29oS6wiK249dPMlQYC
2XTvTIrn9YBiHNoN1dF3VGCjvddhxidRzRJ74tMnlaoqWBI0G3kAFGIj38aTilcA
S18kv15xUVru+I9O3YJVGmaCZzRRT/axF95Nhu0Y86gSvPXrQWlO2FZ8KsqA2rFy
b3iERAU4lE/eG22MtYe1JXufr1EiqhmNTFkHbnDPFsrrOALOinp2WkCpwaxC/MN9
tNVFf2jTMhDW9vnJalvIRNOVMluIFxcktW3893KxKRY3kdiMWSGh6+VKk9DnumD5
XM9TORKdE076Q5TsuSMx1NLwV80J2RDYKLfoJ0Pc5zJG6pVkNOvTlx7A2RSb00jj
297p6vK1xmRET5VNDaRlbs60JSbZ8zvqiqe2W5AbYtO7uP3+NInUMUJNiylXRt21
6PC11xDiw5MyEaoC0ZuHfB0aZVYJk5pDqpZ142QxCOya2pvxQKxxSeseaQpdruJC
lIL+Cac2w2ArysoaMuO6vcxra3wPLd2kbyLspdBvgQut18En0OucIHQXBQW8GTCH
6OoosYkx2ds0GnH1wrjr19dfAmsTKVb5nN/ncgV1vrgf32zeupIWUHSCeT2UyEl9
eiSVLzP4nZPrpn4hqXvgW3ejMAN0Jb0Y7zDLTmG3ab45feGvfk5PBLN7ihIAppo2
kk4F9DZ1s0kvaN53/LDkxgAmVX/c97oXEsw0XYyGlD487w8yfA1iswB3kQkpz1TW
Bu1O4K1jV+BmFKp+bd79QsJGA4IUqWSecBjPRgLff5hat/KXaq0KDwQT7u3Sp0aY
1oXIRYq84ya0tRacTcHgVNJrN7h6K/8+f1BYbTy2AhBiiYvdScHAZ3dCJ2Y3sXAu
xgHBeKeQCTaMCBes1r7cJQ/0S/EcyQ2jO1MADiIPg9n9e6zOTlzjOIeUsN5FVJGp
bxDpJ6dL4PdHX/O7oAFTiIIGu+10SKPWTwSL3cCvjHSk1KkCxf6YUa+yxHws+0gR
Y5EQfXxvmA4+FiJBOSOWWsmiMPHkgBusL7+tOotFnkKDPP8VkU2hAnXD++TlFIFz
0/tAUcR3x2vW11Cz2dWaKSeEGmefE9vD/qFiagLnl7gnIHrLmENWAxx5gZtINEQ0
IuhZ968pyBMP2SAqDUT/uBakvsGrdAvAYRdp7UqtBbkYiKPqz50XXcUw3p5AwfoC
OnEYgCtXtVZRXsIIdk/uYjH5jY3cwJLbm0PZykJI3YhpjDJo8mxh16lEM5ie2eyM
uVvf6C3an3N4GRS7A+aTdLFfzEKH41Fsj4lojbqqXfiejX0MaUwEwJHGWqL0ExzK
TugmjkoqG1mKoLJcPEuFEUdtFYnypTyozis5Q7aCBEvTINIo+WUbx4r2Y9x4J+AI
hwQ6YJVZ6DRB1t5ciddZekLRXv+jYZf328+XyRMNhdMK9Zz2j+wp1Eod3XT8Al9V
P7nsScany4pfAldpzJwM4CjHJwVfPRMBJcGt7ZBMnK0zy8SPodQMdmQ7wJjPFJkw
aNr336jlyo0t3NFvJqx5BnZJYP4UVtGwqpUHzEVUZXf0tWJ8hZZDSkcGA/Z0zyBx
JRvtNQgQIQ36BZ/rqb8xp0/mY5YVzbHtVaveH5f+NlLO6bHk349j0CJsyMOOo/UR
Fyvgpk52cAyxGwYCI6qe4UQOtmP3FnSwKniiD4XENk4h1qtRWkM3oBnCDrWZrlmb
YGzCPsiDP7m1B1bVAjE/7ChGrdjKaksqrR3wHhwntKHSC3QmpN10ZKc0NZmtFB7H
ctIZ9x7AybTfT2tF7585S7DF3weWFxQAmJF1lNLEMJLMw1si2ECyDzqORnAt3lsS
Ydn2z99Y4mM/eCY2HOULOxInFaNN6x3N9+u3ecH95r9LU93vNDlFVP1YelsXaGUH
5AfL9RA5e6pT2Nd4SDvO83lr3HlfZRK0pozeX/YbU30sUun7Pqbbivc4K0QoyH9z
9sQP4TFxRHsYAxaAuoC9+Dv7/O5PDyAc1VD0jqSrWBs3dBMZeK9RD+SKi57K6zZJ
riYWVO92x3bzmL6O1InYbJEOuTW/d7dO+srY0cheWJ2Qdfz+766hds7jSlQo4Lky
z+TN7i3oSxD18XvcaoYAvu5sN1VGNP51AvaJvdGRfw29Ow2T86jvlRKPVAqkmD6U
7kJgyinnCHRaoVNV/7w8Yo0MV1PwxNptGjr0XqKh+8DRMS5xJXYmxRxdi5jr3uMq
dKj6rFjmyd4NG/5Dm2CnNrUWZkHGVVhTeHPCgb3ie/DWu9ZJAgbIJiULeN65N3p8
Ha2uQ8yNGxofNW3Fhk/GEzE1fN77haX7uPt3k65OcaD1OtYw0rBvRRVYsOPLO8Kt
bt/Nq5GXA1dy9wO9t1h07jPQvazFoHgWiME6smL9nl3wQPGeRXonlnj9QPxTUWaU
LDYrMgw6wRFrImYNRolKFBvQS7limpALnKe8Af6qzs+TGu+1CwrbF7ZCgVKVm8K/
`protect END_PROTECTED
