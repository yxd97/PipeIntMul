`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1WvY4ybrpJg9szPFj6bLcu+wdXhbu5Y4wNi2UiKNoi3seR1700ZTM0fNztrgbBbM
qvUaZ+vppewCuFwSEfwxlqalzLOYhne2FRF7wCj/gYKA5h1T26t2XfItHwhZuPpu
b0/Q7iFYq2RdovQlHpkUb5GpCH9sVcHOKFgKagfhO1cVFk2KjTwxj0/0FgZMTH9+
TYjkMOIaCsRXe7pMzDgDpSz/J+a7tJt9pBss6VQ1eN6yNqS+CkgmSgqo531wltik
h/+wYuq1m70uhmxYQYpM3c3+3WN2uhyzP2FKSqsLqLLT2b6fCknc5E7lFCfDuGBq
rl8QKdKTSWkjd/yz2PjYfjsbGq9aRE+RtBZSOTCI2Dem2pr7LTlVjh1hzaVkyT82
ewVV786GVxCUwCAKhu4JCpXgCuLPgSTglMP92siGZ1ZsASzKoqsfYObkEhGsS4b7
PegQ1yJ3KRLGYSPiRcC3r0De4/BLMJqoIv27Q15/1GHKlnvt2rYzE3FPZPoSN2kx
r4U8w/gCxL8F+qJSqQ1fHS13+CJM1BVXN9adXWoO84N3pYvQUd6adUOfung1QGvu
jWiad5TX3qmzgVy4KxDLecLyVJJuuR4D6aY6eEGiBtM+rJcjzHRnQIFxtBR828XU
oA31FPIaoYcUvLPAgakmy0plyktPjf/xODkxMacAqhOn8WNkm1q7CqWpctCW+VEg
gSIEl1+KJaJU2bk9IyPKbZ+rDXK9okwisIeEjrYEN5w=
`protect END_PROTECTED
