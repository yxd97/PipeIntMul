`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zs8R0dOTLF5noQGLDQmLxu0WrLOS2A4jSVBgFkCT18hj7jjI/9UocftpMRdj9hkZ
ueqxQYfQySRToS1bj/9hvTiZjgyk7cusp5YYEA5GOQvUdNxqyRmUKClWF7dWarSw
n0grm0Gsyrow2cKduU6RcDx7Dee6yv9yNrmbd39dM20TnnVel24nu5YwJrstbggf
gJ1IXebkDG0HOqS1O+JqrqoObIxiS9NgmrA8yp16OOePZZwSv1U+KVT/DcgQxSCC
qQT4olZnRMhW2lPWHftznL/+jbTYsPu25VgjmrvajWd0KvR+6VEuWeKGnCLyVt2f
siQ8qu5ZcUqoPTWCwSxzL/7Hbb2dLLG6ycbq3INlTrWCSc9/YwFzyRBf2KBBGN2y
Vf3K93edJ3+dt6EqRe2M1MVjxGCBbc10F13EIAIb2uvmApxtD/9cyeGuq3lsmZmQ
KpGvjSjOVCL1kUD2j+pbOHeZUpAQDfVu2Pcg2sk+JIOqZC/qshpgxP7/DAXAMydc
JfT2r9Br41XwSnHEe8letwsjZ2hG+U6CtQmufN7sezXjkU6TXQdtt8PSC5NkxAYm
40WRwivPL31f5IrxN8EySscDfmZwX+8CScjePuXWqF0i35EogPG517adK2TJ2XbY
+YzATymCi2pccVESpvoPJzD7csXtf1aK1PNJVSrQOKI3MklKVNfRGNUduFsEujQo
YqgJVOfxMbgLtU4c5u6r7k70Uaii4hP3pBqkGCUkVm9LZqLTuVQ/YjdHkRRZ6/jI
6mV8+dI0eAkziSiAK30/RXflbBExF44UYSGJvziUytwaJADpavAE9KB81fYd1eG9
SEANZorw4gxzaG4LQtcOKUckQmK9pZbj9ODYz3BZClZE6QOrdbIdH5mSMHkKCZss
9pUBN7UsnEcnKsQkYRuZ5+jcvwbXIMC2ILiM2TBaNjEZvbHIwxY2jbvxzelshxLb
qM0vVgQH0YVtfbKeiasROcsL/KN6siDf5+pYcp8SpYnFp1Moe739i4PAPTLTcOHt
wYEbNw3Kfqej/4lyjn/dSatxG2Dcwi2v44n495nkV7Ztcjt1Ndvu7VBh3bRsmlz5
cTk8HNzTJPuyk+q072r1blERlVqm0qN8g5KWFQu+Y/YwKgukdeLu93iP8PRFflb8
ArKAeLZWgQBtiQOtxtcv27tbMpsV0dOhflRfICLpFmybwVlDOfluymshLYQgXs3u
CZ1JQHZnGVrDP9lYO3rvxqV72VPcFJkVw3gBTpYdOR8B9lmCC/ybJrwrtoAbNoju
f/SgjbgtG7+M+yKHBFMsfTPHginrEFsSmS28yyjw3zRRRo8yTTHQrGhki+i/bn22
SwrhnZcobBruEv197AFyyTLZ5DtYSGtLeOhyb8Tgdb9rDZZD+Xd/jLNbTAOuUqGA
`protect END_PROTECTED
