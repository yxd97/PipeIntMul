`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CMow9deB0FjsSAEKmbvyvNiJ0rsDw3kMix5rTwxkA6xchsG4RZxMjum1r7GthE/x
bDHhRuJpl0n+b0I4Q1UbEFDtl2HUd2egYwQw5bYXXeQnxFjpLq0JSQN2NM0oKJVX
HPfb8Nd2OMeXZWohAN/cCewQQ9+UeXvwsrjT60ZCgtI/zLoGqgnLREOX+s/hd31E
sDKQPyrn+M+8CpW1N8o5iMRCHTrQg5+Om0Q/QId8g0BmVY+QR49LycBzxT0JI3Sc
dqnXLzZ3ZP+QmIS5uwS/Tme/Kx62WByaBlSKSS0d5hma+q6qjsMZVCshKs45+QT7
mRd/COL7OGQi7GkqwJcDvyH2wHLgvIicP/Yuu2hq5+OlU4fVl3SmmCNmE8UhYi72
MdtlmGCTkVu3wcmRaeAYcWaiVY0uhA8V3buugYhw4bIXj2B8AVyetYWMnU0lOsSX
3ZR/+smB0/2CwESb+24TaMSbpgP5bH0A3B9w3cGQQ12i8K/NeOrNoJB5IVi8ejeX
WAhFwwNGOqgxy+cpZ8qTaSszb2dUqL81EJrV62AYh1b2xeWVM8FlIfmCEtiyT6TI
4NoRmSrodMO3f4Xi6YWYGN1ueSUTJ4gWL2s0Yhit5n20amZkQjvBtKLFu223nkRW
gRUJX0Qqgykq1AKl/HWne1DiUdxz55/dAUts2p8iUWAHV2hPj9xUbukcffbEcnEM
MsR3LlqDXGPuHPlHl5XyJn8egbmi7ztTAxpso2gkNwzwTqbE95PcNJZ8XC7M8Kvj
Eet3LpHIlUkEwWl/RIajZbXU0mh1qkBeoSMF+NcRINrpNtjrry5iY5vmMM9nPA+D
sFDDlKCqg55yNbTWZJXUpwavGkj+MFSCpUPuf5Rf6Q5QUe9XPdWkREDSMpN63RIB
/wJlGVZ5FyFm24RwYe42qJgRX4jHXMD7nCSCQIlrp4YTlwfV9no8Ag1lwmp1fse9
Mte2Rr0TtKp+juJLzDeQKiRFsBymSBtKLQK3e/RlVQ1GZiqSxyQVTQmw/RA1Ukfs
6EJThMzrhVLvCeh7uZjThjPkAPL/XL4M8l8FFUf4HbU3zyZ8etrd0L/6H5bZPz1X
Q1hXeexgYPV+F/rl4ssiVKyPKFhbfWGS0wW2shXKyt6xZLiBiKMl5TFgtNAUSCD4
sux1LpSwn10sig9ltqALWt5T8F0ZSLUUXQNkZSo6vXrl5sFU3i6zhJd+j12XaxgW
BYihQGBXtZQYfkXVXLeTM16+1HWIgVivp/jDVRdeP68PChn+9T3oRINjUxHfaA0+
O/plVBPUzGvijZpRfkFGopQgr+24WEpgUtCnep9s+dDiP+nepNf1tlcfaJ+UzHhO
Ht8RUXkvrxY+HDAPfyhHdnBgQOwWdHSOYmY7glQKPt08sJtZQkF70hrHfLUS6eP5
m/GIlCiaGOlRu/NK+o7vhL4leEkHLs3HOrkNYtkyEC4hy2TL10zONNGSJTo7yAYY
5nenZHoHZCGeZ1nKCxuWSl403234zunWyPscuw/HNHNKim/rtVaRDb4KyP7PPKjJ
ST0TjC5B8YoNpghvwwT9qzjxYgMBoiuof90D9ZCXP5qHcfjRfxt6SltlFLiR5tTk
jCtmYvqN9QBKybsm7tspkIx+8Vieb6p38YqgfIy2vX922sl+lNye26eLUcfNtcdm
iDEDK/z+X3pIEhx/B5zPxbw2CCppcbhimi6pRg6L/xMNZhOoMNtqxXHAHFCv2y8X
1Rv6slKtMzS46V8ZKTUAW+rsUy75wcyCsP77ii9/Ktx2SmfPBUpI2F5BQXJ8PoUt
ot0NGg5tnhxDdNJhBumL08qCAAZgLhKqsvB6GasXnjMPdTTFqNi7dG8f2kB9I+OY
DdWa+9TdmMu001cfSzR9yFgDqV6DbeHxG8bacFSEQq7Tu2CHA3lJcAw1P2xNViYX
AK6CrG+OBkNAj0sCdCPDB9LM0dfCa/sN0SEbT0rT/fQtPRlRoxh7TiyolMuDjmTZ
tvdeVgGATh2TCczzAmAyY0epCm8++38cRDWt3exhK2tic85QXxEClfXzX+7Yat+P
jqcP3/mkiAZfLauaiSVdMaLyQZf9yU7/0WGAe+bM4UAAcD9WkgLfZfdD5+TMazbG
6W3su7sVyFEg/hU839bX3mi2oq2u+A6AfYK6K3sHW4WUJA7RYOqD/ie+o1ShWlHW
R5Sc5Bgv2iQ1Zsgby5X+wXkvLl13XvTdW84ebUwejy8lHPrayycNzKHdcpGCfL9G
WImWVKGY6GVYs5Jh4KIo+rQ/jcD4JdVIqF27hEpI3z7Fu23FJYlwvS1NZscqJb31
GSQlnldvDet4j8O8x8F1u0zdFqNOvbMdYiwPloIU5s7+2pc0D6jZzun+RAr2wnFx
Ik+WRQ7Mz+J3iyF9I3M8U7KmJGTTQmpRwjaMKsHmWYx0hdGINYSiso2JB7UGcVDY
BioUPI4aYhI12SefbDOnu3+UDCxN/f02VhFlES4Vp6A5CxaMFUPKBBAObRxs/3xX
0cHhad8DFoHjVKu3spebWsEXGRoeHH7TqKa0vHqDOnvMD3IEBFGT39dyHiphdV/J
G3jhEWx1MqBGmPyySSPUH9Hid2W4KfHWIw61tZt9WUnr8mIW1Jk5t6Xa8dsNO+Xu
k41dkC8X+mBg8/05X0A32AqJWgdTRr0FCXNGAdRwllReL56lPf2Iynlk3J/YhzPt
De/HMsZKzboRokwByJLBB7ITYlv5HAS1RZiNtFT+oWbsQ3TUqzg3LHRdNHnNw1q5
RAdRZgLhykDP9ayU/FMvHsLW+zZFnZmdPU0q7ZoYJ40k3Ozep5//FOQt9K+u15d+
nFIefjus9hQ08NUPySdHcvngtNh6M2gHbdXhdD+h3yTQk+AmxwGh/qFY1/UVfOxi
ZLnorPQOZ6LsyhZ1jpAYtl3aCi8FyVjRm3mWeYi+yES4zgrFmh2eh3SApa7+588x
eLvPRYSOGzWrQezvzdwYsmj/2H2tscnXiH13tTEQeJ3+UHL3+p158FaSnH1LLz7H
KbiQdNu5LU0CDVj4u2y/H0e0TD7CHrlGl2pmA1gRO/VmOg6SPaqko8bZzTDuv5oo
CKn1VF0f9rRttx/cXXUpWrN0NKpns/PURPH23Cu5Jr0Lz+UYOoBG4X9gDciJrk7A
8X9XoElMMmruMW7fd4lX3k4LGgghQh3Z6kyCs7SqKqINZM6PM5GyTuwjgQPlz1VC
RHj7vWf/Dm8g2BZte0qyqshN7haH8Bsfh2RLbhoVwhV/TNxpuxflSegkB3mt5nkX
aQ66NAXhGzHBoXPlIe/lO0lP2S77cJlHw19jlfXFW++jdB2NNvcIAUmwNVimidLi
oYqprJVyXJ7mGiUO1ooXFgN22WwHqDEOoz0gXPacGblu8MoyhxTwyQrD5PVbBRki
3lLuHdOOXwtqOSvIch5Sq8C5B1avr03L9wURXeoJvtPz/eyjd3zH2hBXB+sB96ZE
9E+OICWplfBCjTCfb6cTjcM+ldIKFtuaxSXKYwMB7+eR2wHAMlloh7/2HPWH63hV
8QeqCsgwOql0BEtQ8W1askDyqpe/y++Tk4ZsgZLjT0mqtrc9Rn4dYOvmcTgV8iBF
AAWWOBQos6Zmqc1591PBrTmxiOb3VSLjaWieOx1ehifEvavq59lmJA6yJq4smLLa
LjFsEUIIgEVPhZyhrXBZk58IQSktVFckhNhx6YAZ6JX6MQOmaZCnWdTnDsz1+KOf
5tKHjbtjpkENSLcN8t35OusxpO9e0Kstfw58LmbkV16BtKSE2bto6H0YTTgdjmcb
MXgv3nLyMiUpTbkOtLDZInuShuSCfEUaVJ4H7oRaTNrZeK8grjUuOsA2hPY1+e8d
CFjvsMgsbr5nf8TNSqf3pnFt0Kq6U2OYTSTQBAFjBK3wGdRCCAdy0mCk9WzGYW9u
FhO5oW0leJLmV9GSD6pzXq596GawrOFbCq/p0u4uVWBJ4UWAADvC37jlzjTKbcPj
ptm0n74YqfbwZhXk/zPzbXRAxjOWkOeZ+SXLuyZ7lQsnqfOwtpat0pRmV05Q+GI3
SHkzrrRpVRRn8iyjuHPVb1pDMWgbuU8Tzh9fQMX2WzB7W0WTgvRq3zvdt1hNASCb
dpaF2igEILEdn2CN80lWsZiyWjjwXfsXlz+w5NFJPrcuc541o+4vYHD4QKELYNL/
+4HsuZ43rqgeMhDHKA5bR+B0VC6yDHLYiNCs67G6sM+9V14XU1AuWnZ1LkSaGYlo
5dxIrc1gORZIKwNaqFNCpqfPc3hpGtLHQGlv3tZPe1lx67wU1P4OhCjyZOqz/E0a
Bn/x4JmWPKGuhKPL9+msdcE9A94gpxw1I4gGpXCEQs88F+EEWQKt9bp7xg47b7l+
FvVyYASItTUN9b9xqkWqgt/wGkpQCd+tKnRna1uK0WZ5ixZPv2xUF7WscYZBjALJ
qCT0290psSvOe6/GEF/bI6j29JcKDP9OXWgU3ttf0wOWCDwlBvx97jBDkRaDHJRu
KpmAm2YV70gOcPLwAJRxrYENduvisCrfa/vdAe52IREcb3wS6e3+IE3eEmMLlPNx
TvZJcKzdL8dMOh6EDslsIG6xDZ72nX4saoJ18puf9paZuzFkTVKuGotrSf3AGIqH
FXBV18GZTOYHIij908pIld0S2stbgAUCEx1De/yaaLHZr3RfMAZpJFxgDAWLMBCp
K07sD050ogpCBJwNPQFZOgmSlNYcSNGc5uPvHhwURg27byO5J1DoaP+gddQNGveu
BNr5YKPux4Ow2MlU7Nl+voIDWV7qJj8e0RjUd5ObnFTl1Kek3F8bNSoatDo/QK2Z
HguBGwAg68k8JyLeqJyTL9c82K5ZaZyx9w948jo0eKrVXjoaOMAipi09Qnet/Ega
RICEf9LMUnmtd8qHaV6fdsOZ8KfstMzKGkRvYilMhMAK8R/dZ4VB6lMe3T1KsyFK
tzCO35kx79GpCi+EwrYRDROD5oXOZxrwDq1FI7xrwnkTXBwlswFNBQDrxRJ3/IEE
qowg7QscDcXpUKu4X3RG3LpUwaCA4pUwIhMbWQyNKurg32RRbd0ubQ1c0ZuDEqBV
DgDwdLbTQxljZWEMcrq2VHZ1oZ5xCl12PFoFX5II47GiOCNAznqooVvkAf5Ucwp5
og39sSHRTBZbfoiHRNVyKkze6nM154YHAXznQu9qgMs9sYj/4mjaHizUgoxpGhSZ
iVfAQS0SQfwSAcjrzIw/BV8EGZbO+8G9e0cTdFWB9zgJvAT9/mOhxFiHt1DAJwOn
mHGF/4Z0kte3hSdfe/z/qrg1HZGLKMcY2kZUnPlHxUWh92WoTTuJl+v2x4IupKmv
e++uBLZ+GcHM6INTvMgXjYKWBYwqKhg21YuPYoVYqOg4SIXirKmBkZ4VE1JIsAJm
bQTViIVMuxEB5F6NyUxdLw4xBg2mKnOFDDJ61PJ0gSfLbGUHLNhSjgcKiGw6WJH9
7bufsy4LbRTVx23jo7hKD4oaxlWPB2wXa7GBQkY2XUmYgpU18f+rYzHKxwKT83hr
YR30wu3eEwYq9TGxGIwXfPEcQr+pjWuIAFNCyrR3y5poYxx7r4+E5gMjpO4soEOz
csLDNoAJ4oJ4Tm41iB0u91vKsumqjJbdFzUr1apDn+FfehJu2BxnzzuvcJySMftj
PPls0Mw6nd9Y9RLvA2pKRkGOCd7VYaogt1m/rqnaCE6Dqayfd6eveWxemsGwYQ/F
nMNLLN7rS9td5D3jKgnJG7ZTdnX4hrPamO1jD2lhO4Y+kzD4PlSGZopnZTanPnOD
vuOFPSiAkq+xPp1Z6JJTRLqIVKS0XGxUyFPQvipjc79FzC8b/VyTPK4Lxw+a6dbq
UhO5ozEg6vIsVn1vm18XEoy50VMQbR73QFXwxRSB4nYxaVp0GMyGWmRcYFLKdDPz
r0a6A7vPmGoAuPsMprP5rQCHNnnQuTr6fD7nd6aE4JsxprJricwAbE6GvvSOE6MX
Fwpie/oTjkiWb8KJN1bQWfe6lhSjrkUeEQL6Rsjbg2NCyKtEpyum3lRtKdXSa/Fb
Sn2hi808v2piKM+Ve1facHmS4cjYHdV2JE32F3+OxxFeLNQnB+Jypg+waaOQTqt2
O7RSaALUg7rW9h1Y17NVffZIVyJrUT6CqtHttS7hr3/gFnhsn1F3nb77Wz/ElSYq
HhLpBWE2eSmKl1z+PxxjZceIM4QXw+37l4Ju8Y2UeQ551hoD37HAYOf3JOwO6FB3
D3HDzJ2+8N4JuyuMX0RKwzwsrvifczoOhF0dsULz7rm5ivzujZIhdFxo05h1gEOy
ALeX3nnFMqgxJdza1p2AjwZQX1QIbvI4XCRigef3qA83VulTmyt1TpPFGUVsWB9F
SgFTziKFCjWsWyXNgCi0dhR7+8ZiEGIyr/Yhoh8SNo8wMCY2NYHkL90ey2GKdzo1
5iWH+sw2aTMqXChf7Aqj+JQXF3Bn362mRnZO0b4T7eBGBwmXGlZBlPWzYzlkp808
CFdgQMeLsfKR6nxznYIyBzN1cHfizNOuKE3+ikBFI8mcRfjl3sch/RUmgG1hftlM
mpzCn8QaEzN457i5+8raJuxAM3luQ1PlehpGE7tMFcUKUv62XI5sGm8RW2Yw5fCB
B3HDOxmS9pSTQ6T52VH2v4QXTH2idXEhoRScZ61dN/LAY64kLduyM9vUOM2GxrhC
VK/XpBQLpycrYc/VokQykFzSXG5CtpfmfYJ13sOjAD75HYAJ6R626+65qHqTM8Qu
Pa9UOFtMrJSNe71Hxofszohn1RlW4FNwMMrET+v05v+JfGPHNlFRPDHoDyd9ksbg
8b2lQM9oi+iqIP/k0OpbGRU1eCLwxjrfcGmtAPbURNUqwnz7Y6lcGXuRMb/cWiIJ
6sCu3uaBdgNAe1UC2Njt6OQrrPgYAi6CLpeOgpoE6ehi5jcB7uahQYqAw9cq5dZ+
trpcxaaD0BPe3TKf9zQaqe00gAYF7lis2jXQ9GaHrhTn90ArLHPH/xCUi55UsUHX
r+CrymgbAvG2l06zHcVvS4Fi2BfqxnsMIphUecJTiGaU9rml5TXVBU6Ws940u7iN
G2c/wVR9uU7UTSuI7dB0QLC4aWva7tWSS0rRjKH3u/BEZXQCdPttvEDNX8IhMe02
vV2HvrwJo4XdYOTqXBnsE7vD3BKRhNc3t/ni48mQv2HpaKEDJa2rVpKQvcKl7RWl
MVQYz/dl9waIkq+s2hfvs8CldOEShpNpV1W294MNh/i6W+8jo9CaWipC8YUVYTDL
rz6IPpntIJDRW+qoesToc5XSLzlp6fvGW8iW89I4Wg0sRi61uwPJeSvKYrVAP8DR
XM8l9a4n/lN3+2XzGX+wufHktOIA8MNXI2kaV1BWw6NIWeOnXhAYlrwEsNtW1osN
s9XBSvqPPY1z3+8CLUheSICA1mIeNCvO1Qk0FuWDH0Qn77deQfZYyE/MNXsshhSM
6/hlZL6Y6GuDhO3fBMEgJVNvdK5HiFkNKoX9z9bTbQqHk5VhLlcDGORinhjgZNUC
ranAqWP0NCH1VftSG3TKh1P9UiOcjeuJ0abdFUDB+8o7g0UjhI4oqwNYLCwOawnr
OULOhenlqxOkpayaXilkXjDn8DHh4UM1NC1BDWeHg/FPDO7yLHof/9hM5hp/qwGn
KLDcm7Qus9siSU5QLFROEy0bppuLATdfhKBUq8nnWgvH6/UvWHM0tvMf7N6zK5Vc
2eg7R6yJU21wAGCSEAzKAiFz8iEOK9KixSjXCwf+O7VTZ6U36Du3lTgEuKlbJiY/
9V4jgoNZf6s9cRROWjnZP8guomBb5CuidARLrbMVW7ycj00jN3lrIP4uWUH4PNYi
DQQiPIWk4J6MeVUxF6jUpO7TZrbKOrzSlvDqUDo47JbjbnULM1TR+ypCMs4DQ2id
i7+/hx0QEv7QPoHq3rI6xO/mrVyFSzFStpKUBsLCBuCIcSfCjrP9+IGpOK6/Ticj
yOfqSjLqpGqz3vwkoxAr9cM0oFpifSKV7TDnssaHXr8hQctl28MyvBj8zp0yuYFf
EJFkql7R4pPwlJ6QoIuPZY66s5DGtGN4SUAhfAlPSNvClqlwGiGihYJ3KGt9NXo2
Mx3RkifsTh8w4YamByNyFSVF2Pep6INbXbHL6lkn7SqQbbOybVDcdM8mkNYaP3zE
LDfauU5bY94hVoQS6mn6SAaKGF7TT0xxKbz/+NQcMk5JgE5bnK1vKzZ9pAfzSs1f
QaE+P8Eb4PtNLTNeO7aI4edEH1oykycNtaHhO6DaotlWZFamdiR/u0DGk01Itb+Q
oD/nsTBuBgKR9kFZeYfz1GJZBvC3IK2Dut6XBoZAMCWquJKUjMHSKXJ3m92qZxNB
GI/gMpE+h5N5EjqE3kkIyYXb1r5OV/CePUn6yuoziiZ8fWa24b8/Z0bv3sWxiaFb
lfKHlUxjEjZIxR0BRA/xXmqJuHLw1gz/kQX+ZTe38CbbZVWTvu1DqBZtE9kEN4n/
D8meVOdrMm1KWXkxz85sFuVSvSQJEQtpvdCnRwh9JoWFMckhzC6IqWvaiENZuusv
rnakcORJzWRjHR5l5rS26zpqSPgBCc2E/ypd+CNtGNCqtU80qLY9I6i97R76km/o
bIuNp3GGWC7zPA38JVLjW0uUX7m1BseYlQuaOTmUXpG3KfIiwtsQWrviv5wmXuJG
62xp7BIah7kkDQ7coDloi1JdtUFqrXnWzk9nf++E7YO1XenvNNO7zfMxmkcZNgYj
KdvFOLLG7J5ZrkX/4lPP8+ejRhq77kD1JFbr96e8nnlxfq4c+24KL1wj5BJ1C+vs
zWt6A4tCZbLfHRAdchS6vrX1/sNci07OojQw04dbalGLxY0IfDNQq+uD0spLX3Q4
0YKKJ/ubPXpDhk00Rg1LXB9Ih+mgXMGQCqKtALdWxY6yfC4z/VKpj2mbucTa+zvF
hY1EGt6lqNU9wS+FS1SVuQkLxK5prrMzEe29B+c4v366Ulx/5FxWOOLFGxgkG83o
L7Oojk+vw7IuIfO4ixhoOQAxPjzwLeIgWIswKzRDyFrrDtyTVZ1Qryl65aHoxeKI
tnIhgH/eKCtSocDho9jT1fga9Kz6m6xJtklwWNM4LZaZHUmw2pphiOK5FfjvsKoe
Dxj6zCCq57K/1qkWn3O/jrjXft9l/Zf1k4SSkioV1TYdUlaGpONen1j5BV5/GY56
d4iXR8inpVp4xrs/58MTmdGFgCHFgGedYC3qYJPeELFgN6Sf942VZfsJQYmVrOvq
1SLGigscwuzM0FYB4jfQtBkb5Y6PylCBZyx6GnRpAO+sn37nmELsYKoNTEwlbF7y
fydNv1h71k482lN6JGOI1ccP+4WENlt7OBtfeTC/UU+8Qubw9IQUvGuQ9SkzDunj
/SrmYgwUEd5QDNLHOHFMur0y73cH1ua+eQvGVuG4Wzf6n/Etqvb7T3h8kQDuLlBp
+ta6hjvJDSNsZsR6agOxc7yYu0rA0RXaY+lBpqDMGIQtd2lzKdEyqFWq3GY48vSc
uAA7wEuw81iYoMK6m/c6ye8rw2FTIfaMuqfY8JXMQCP3eDrBcRQVn/9Sfkxyp5Aa
imq/WIBoyutJ+l4KGejpsTHca49TEKsuP1ecbwMUdZ9ORSS2Ne+1RMcNFP8GWdEH
Nu1r/mQPTbxbKZ/DmZ2uyv6uhhW1UqfYyxR/Qwgc+jzdL7D15FAFPvkfugNssS0y
jYbHMj44N4mrXvDyHALX4AI4X0DQOU6yj83Sk1ngYmPoJprzhXz004zI8wOtkrtY
PLJhvzhlxkJxm+aCjgrSFBQEm9+acCKBgh189n7BkH8lCHt3I9s1aM821BmJUDxg
cmcQV/mtMAF9O1kyA1GSVTtjzT15ppWfLsXaOkqWwTRan+W7Z8N9gfiJksKajZou
1pQyfrWCYF6p8eSGJQv6e0V5Sao1XoVr0ZSivbE3/RYFteYNBPEX/kjzDrnt4mB5
tGNfuCFq2tNHInrjj5evHJn64PgvCydpPYo130f2GimUAUAkAj90HkhAI3JYZ9Tf
fcBh4cuxG5k9signcMB0oe0hgP6MXOqJ1wZGQMOmHXA7WOg1HuRntnzEdG63xFVN
PCsfoxg2E9rzImkKkIEcvuPgip4xohB4FfJqZ1BKWofYti+9PU27pMLoDPeZmFXX
BtjXySqq+J++I5B3cfaMJ1hl7/Cpdj+4DXyRDBzStWwY2c3Af1uLQvtVWF82tZaw
qzZ/U3HNUw6MzvWvJA76QHRESOJcVKYyVY3YxO7j5wzm47w7U2LN1Q/Wp2Ic8izd
HyzjQ5FHqeEBfZLPgE00u8Sh1OJeIlL/7TX2S16VUhxjM/1YRp1+mh9LlfInE7ah
IyJLYF9sTlAVtaqATnGj7fawHnB5p427yYnedP5kZlZTyWFF/QV6P+zY1f+X+eeB
uWrylh0lc9NLx6zZI4UdkDy8sjse5M8skK1u0f7uJUD9ufdEA1L9CiiW/+/k9PTj
/2RgeQKOs539daFZdrUcsUl2GkQw/qOePHFEs2O4BuDXU+7kND7lSp0v29LySQ4D
JDhsOdWl8vxJb0b4yj5BKEW9BftJeY3+4lgK+9zXxpxo+kK3nOZ7JqMCMouvYqrU
d/x6ZuAiO4RmdXH6rezanX5UgXcbZ6efBovYX9mC6wIEA3K2+jPWrtqtgVMpQ4te
KLlJ8+f/LqH2IBIzmXVk11iNKjWBiqimyZllrmE7zuU9xAw1lEde49cfkO/aLmdv
SUcqrAJwVv6UPr6u2h1uA7l03T3hBVOW2gJRmiAA+4qUzjJDAgp165OgQBlw2rKr
aRo9/+Ngr2LFJGwmtI5t1y+bLQ1P3s9NQwrCChbv3x9HPfXKDAUDqYcMxkMEL+Ro
ip7bykjNO3kmhP0okeWaNn85c9qb8VHNJ6MQw3niMjg8n0/B2e3A6lAsQpSsC82n
FT11HWPwjoZHqlyufswt3Zvev2sVejULmYis7BwUhAqZap4djBACmXBLEsaOGtgw
PU044R8dvxTzQolGkGNIvZKbQ3qCE26867qdYENCrigjsyN5ZSv6IBPQsuEqV3oy
FhKLDCgCE3l8Gs1ZbORkwSICyts/T4bcSeOirg4TfNXKZ8C2PrHTEjLVBb82X0yX
/gALBwAKinP1P7DexZciArzptB1ZF8+n5O8ycQDp7M1Gc5m47EEDnaJ3qmfyzjIO
V6v0xWyKFWCMjTfrUFJYPhSd1h0lLe842IJ4PpG3hnGRrN2qX7ePFRlXnj6IjfCt
nZFnJHs4yl7OcBzM8drZoBq/qf9pWoFb8md0An0TY5S08oYUnIjwdhPSJdvRjFtn
JbkN1+dEAjH23KntbbopmsoQPs1oeILTzFRkGuv0kFRzdXy6mzX0F9qmkCQwQS+v
j9tgut5bFPXBHsE1TasCG3fGlOFZQPUBABiYdmn6AtAcU556lxyT8PeaXyGnZWOx
33iw6hsPt5i0IuwEwhdCy7Kd6Bm+ICpeSatNykAsPTztSkmow4nvfr2ZImexR6gK
fN9EYeFvkUJ8/mIoe6NMLvGCE3QqaudPNgMM1Zl75QCaiGME2gB/rWTld07iU6VV
FJnyJ/ONHYbWuctdYIwdz+HWggwsCq7N6s1cp6Q7OFH2jdjr3d6NhF7+Moe4cMmi
fCB7OcUdn/tha7Bj0MMFkQUrfep0BU4uYC1BUbtIzlPdKmcsCyTBqOn01FGYPsh7
53h90fT+As4rgkS1A00EilUMHVpQALyDbbUNE/xjKlxjRcW7vemB77Yw1FTlrQ1p
CCaTQKdtR9PZvKERr4jwPbmV2o0bO1ltD2j745HM84/gU9UL+Zvj+swz70uTKIfB
Z6yV0bb9IXcBLzNVpcA/raUqIcEonkcdZxUy4eu0yXb5A6FpFSt8Fmf2dZEYT/Og
qWD0AbN3hvxFMx71Mew3GQkVjtQ8RGe8aJrRA/sxRYvQhbfm2DalVt3xAWYIkE7X
+/7TViTqDPRSW8CFwhJDEENDcH6oaVPxM9FXZoxqkPy7egoI2LS2SVz+RzF+tA3e
bXLC2OismKRQh+fDTZ5YwwQzkhZnQ6ZlsnXlNHbB4D/cYAyqdGzwvoGbqEyarg94
x6cygB+9rsxxBj99Xw2s8J92+r9tckOZj6r/r0UZK1IHfOEBo/UELJOYPEQwRaKn
0m9VmvMsTTtSYwwjUfc3FRovy+WBH51yj6QcoLAtdb0Xk818t6Hw57ptbQ+KWOV8
da6jm5zRBu6yDqOEfaKq9iahMu8VDWLZfOOLMG6UG873pGKPBZ9QKPjMGonRSz3Q
J1FaNHvzpyOXPAy9r/godKIq4SMROaIlVVX1up0M9WClcl2l6lSjQV9VoUpB0J1Y
92OmxCwEP8hMFl8BZT8O8C9/w1ULs/ZHlEmfE4NrRU6p0BdmpqHnTpkEymbNo3q5
do37ibmn5Ec4+tVd8L9FtFgWaWrQJcOMtJmbZpkGiw7HY2zzXv3bYuxQb8irEFdG
Kt+srMSFXU23y4TdndzIJdXoC801pu17EWacNtuM5DrHdc5rvYbMf3salevwxCFQ
RCKbTwQX0DfgSsFXOc3H/6+jcLhQDKBvNe1cU2GYBuwSJ70mMfrZr/SkdhOXmxQe
9USRtXxrh+coFLMTYMX9IuHIMCMQqOP/N/3+w7DpXENMucpFtIuedDOYYXafcPyw
B9/L/rix1VoclwNzykHfb9ZgY9RIcQZBcDuyQpKHgjPte6eYOdvG6EpVFQLQu0SQ
x6C3rsF30OLov6VEWSZBrMEISgQRRAGy1pNILkzTSH3llg1MiISp7tJrQ/MBdyXv
YSgXeWrHLTSaXkwe2QBDq4sfw0IUeo12jRZXRN7OWqmtP0VVXfR/OzP/PYIhKt9q
ID+xJiuqZdmsHPmktMjLDQKLgGNUFtDiK51w9kLqNr44DANDoYTw/63+WHsYsLNQ
3NGPIkmLCFURHwv+2mgc74Z583FCjfrr8JbC4Uf6Onk/LzUICrOT45Af4qJQVMXQ
v4V4gTxAh1Wm0WF7FROrXFuhs+EbeGxP/pLOmSWB3NNfOoBUBURc7PP06ZgjsZix
UYq82wT16u6/gQmvsuOaCQwLZDjuUohbQ33X1fKKZiDHMR/IqZT9pKVI2JVpGLOu
9/TxfPJOnGzeuNEnUhS+vSd1bea4McJroIgLW73yRcT31CkMgnjO/wrm0Cbk+XMX
c/eiSi6blALnNNVLIZj9/BEDNu4Bc/chP3fxaGDotpRfj+s2XzfVN6SNLQcZ/t5Y
/NRlcW0vnNR1PBKAiTSX21SBZzw8g6sFgOyloq2tJkyITbZiTTVtBChUDZlhaQBF
pR6TN8BxuJ8o366Ga5iisaBmmsi2naHDiCf5odPB8OUyvnSene8j5SKuM3ucV1So
mKhEnYTuBudvn1Q6dV0BVodvNkCh8uicjwLdq6c8KgLHdlRXvhSnppgNSgxWLsag
A6i8c8HjCPYXR4y0tWvbDueYElpQ/0kHMZSZnl9K44R0nxJBihW2c6vZf+GPv84k
ai83lxSuGONkrFda8EOqUEVxxcsdCJHOZZnVPOp793AxGcecGzh1Qw8rzZsCSoqw
IQWV481eFI6UrnIvqXbQ+G9n3QQ8g3LRK7HxuO5YJS0iZvC4rxvtlLZWVwN8tFgc
cmiUXe0AuNrDOxtWRtbpK/HkErVPGdPJA4qz5NMpHjtqYEcRfg3jSQMxlxApekdu
6w8Ag2/fuolj7jwYRvrvQSuUTWheQUcE6PTHXQAhPuRlxLQS/k8AGpf6g9DmTWAW
QQgI2IQ4raHZX5Dzl6W6HkT3z6/290/A5pZexBsdj+kpQbXmKoDlNy3svv+6eVuK
FSjgAPv4pxSKa+ok1OUAJaBhXl5MPv8GBeaeXE3innOO79JWcZpyGs/PtbjPSCJt
zc2HLDa4RsFSju4CkP+ukZMDca2NPt5Sh7+DjCQuiAz3jLbYAHzqt4+mI1SLIAw1
ROdvELXw+USsiB1tfiNr9T27ppPBSLmYDBfOWAUCqJJQVqdhEYB7w0pS1NNQiTyo
671SD4M5KLRusKWkxRZzoyllUpawRnuauNmPGQsl7nc4+tLnvK3VpDG1LhQ5KpwZ
d9PGzVIQIWH/Zd7hfWknk8/0UDPusKkEq0zlWiaK98F+05jwbbngokcGW5A8ErZj
IIw9McMRG9KitffxSOZPaZAMadXjSsPV3rVbOc4xp91M0mGTXrGpBnV82WIUEpVG
eN0vITT/L8lYXiPcTKeg0+3KnAv+Fgc2DrdI6PcAZVkf81NXZOs4rShvRp27liQB
s2gukMoT5Cjnv/KWpNyDexhi4nZZgiQvwKBl5ivXe7QUdEvPiqDMb8SPse/Ky7u6
OuZO2/NBd9A/4opBst4YGvFlBV17dJL6xLdjgvGvWxBxM9hpR7rtSxtSeBmFgTbo
jI6jR++CJlfE422OUx9QDriNw6zvNTSOrgJV7eWgBXHWHNdqK9wWkDSGi/GgOxTe
SMTxF08w5uW3kJDy7QljpDF1sskg31wjo8tMi9lMUUbdZxPDufTWws9Lmdn9VOr6
sdlgh5mg5YBdsMC8vPw+79A5e3/xbYApUWP3LIdGPI/CrmhXALH7zXXw5tlqVyhU
19X+J0He3uFxYyMPP0qfmCeAHFWIV+b1XbvOQ4svKG/RQnoo1MPKyzw9cOXESLB2
zWdb2N0rhZtU2fNwkaUbrEOwA0Hm0orNJLpDIXctce8f4r6YuQzzFPzKpKbIq5fj
LLE/Y4SrgWIeNibfumJouPdFhW8W2Lkz6g+U4vrZ9l8xoIwKfvW6gcDZQKXwyPLN
undCDydvR703SknYmSogvq4Dm8Ng4ndCHX5d46InKXJzATOJdSvp8wU8LZ6/2GGN
uLdewqlH1CdWTdJiqhNWG7zQTCCpOo9uhWTjIjcTzQHiBR/ARMQRaxuJuz9E744U
YitKGg/9QCR/FjR7X/AArg9Rf2VmnuA1LOYvqsAgNZ0oOxABvj6IHEk+kziIOFnD
/kA0bKL01EhVxj1COi0DXUTWdCed9lQyuK1xPp6eHGWnaijFSskYk1oJOcgdnqqe
btqHVWhF8yYlxhff6KhQ5Qi+197zcMJdZH0kCKzpoaf0ps8165SHrUtBz6PxSHpg
L8FHGrFFr1XPAx5Obslt7m0GLwv0X1epP9Af8fuZbbVKDRtjgYsZzi3MxOmmW9aq
QZ4DTHzOkKz6mpWWkwrx42V7xAIrWcEl7mrifj7xfXWnGdkePfYZS2kXwrkY2843
KBcwBJ/XmDk/YJum/h+w7slj5YgdQGITWPvpM4swstWoxRoOyckqYToba4C9Ghhi
RqMg1g01g/GqTtwtT19+S9a2AdmW7dDDtRhXL8dYdD6pmiViWt5Ada6+4/bC1g54
wuaWpB1O50Q3BG39RynIgsS/Lz9skR/uHbqVccwVG288m7IYAOniTxYzCQXH6zGV
tXAuvgCOO6IgCO8wRKX6NkpNxN8rznkbV6fyx21Khzmkg0q0J+WG9tZ+ifbVKNUT
5a1MKeNk2rMQUJL1g+xVl7Jc15GqDMN92O5HwvqatsCwIhvj2sGu3ryJuYgWY9y7
zduGMiDPgLFyxnzz6yIIx9b/gMqM2e0uZyImo0Ss4LsxJdJUm+qRMkE0NllbkOwk
YjSgChbDOF6S89e9N4SiHtI30Jb5PF/p9sL2MEVob+72kMVEifj2Oi/3kp9s4fEP
lZMftFic97yTfSgTjUP6OetdmCc49U55vyuBDSlks0AG3DztrDIMqZ+AgYd74BIY
dpPSEQXIvnqY+Fdl072BCu9JXUojHqr8R84geaYHW5WglYebmi8aXq4Dd0v59kgY
aUy8ThIBFzYxN6eQ1Wi7xUK8R3xgzKY6KYvdsd0WgwqIX1Ut0XlgPid8iQxl3UD4
zVvcG+oO33W8687vGqTtOKj850nmw77yIf9YCGcmRMmdzxFgjYbWhZ0cJUa3gh0p
bt1GCSET0HmCm0SF+AD8O0fR9GytGWbxiS3BZBfhK0hZikS80gBZo8XaChTGa/Fl
0G2KGUwkAohg6NOFlOadpCuRwsegl41Depw8Qm7MY3+Dwph5QISqCcObIlfgxHs+
aeBtcf5BfZAtGc351yBfr4JgUTnv4gbAoOK5832McL/7eSdMOOZG7qYHPA7hfzoS
Ji6tu8BNgi5mqhMxEnc5abtSbXbdM6mhxEp8havaOihd0v6jNmttxEDq1E68qwV/
6ScT2xWLekrndhzdng1usUCj4/qO7bbriGDF+A2bFv9/kVS3gVfRMW8qxC6Fqskx
jw/OxcWhDN7nnHkiL8ZPBfvCJ2zLswJpw7JD4HWGHVO337+FYG7dAQQLB17Y1nbj
PzB6NuEctjohDIBBuoPcVhOmLd7UtqnComR5Oi3CvMz7KFzkohm7KhrXFadNLKW0
jzvVYWsIY9P8G6PJYOrY+oPuHhp2WmwnyBqjo9CiNfy1x+19uweepWkfOiUSNmMQ
5Dc/tBkFd7uJDPqT+I2KiMc0ifJSxX65NpU6GCmfJvIJGgV1mYU538Rb+Of6UPFh
JZPEtSitlr/nSCph8s/aSpz1znHLzlN3aocmoO5Gvd2hx0CekUqLCd7WyYQWb3JU
eVgGRfDUy1Q6l1rOUWrITWUaxBmdv9/6rDVVcF3r6P9xNuNGYiXL95CGL+LHm3yr
igznAHkYm8GG9onBa/E37J/nzVXsDdMfVNq5XsCQyNPTVFx5deyzUwokt+WkuVBT
Tl3zwKQiLMq3ZdXF8wFY8+PdQtXqcu0uEc+B4R3A7h122F84mMsNhxk9l2HpM9zP
amuaf3dq9O3m4KsgxNKq3lDYUzDr8bk3Owaj/oRLBUwUi/N9/SOWv8SRQSoSdPgC
+A7mb5puqqgrIz6S5z3DIPuDgj8uACuhfK0r1mL/L11KUGVPoJPs7FPYGHkn8ToA
JwTSms3w63sBf4bakEvBBHSRGPFU28088W11hNfwrofWirsOA/iMwtsePPnZERlN
O7iC2PgO1xOQVRC/UjO9MqLeujolYKRVzirK6emMAkFfK3fCzEUjIROId/QRwWBN
RzB4/D2I+e8ZYmd+XH3sT0k0lMjGWo7beZowbNJkz+VjNLJcyOC8RzhacJCwpHOV
cY4S/ztcoySQ65zgmQqyenZtALpY55NM7U83RMjylIjis1de0sx4XQDF8r+9ihwl
U0GmgalmZ5Ob1rKDtFSO+6U6TgSV8eZLQEvt8zc2I2O4BqFafkRJQA9FMUO7h9j2
qFvjqwvRFGxyKQNZLhvU69HY0Xw4e5vmfCurNSElDOh9wldlDUPNXmKpN/z65eGs
5FINYsiKbPYFuPYYRayZGPZ+dPD6+72FAjf6P6+QBbtR2+DVhIR0+Clrozv1t29f
kWCqZGgj5kUYMGqXFgEX3HAHVIBryeoFbLKxBnhWGCJgjoZFZoX/VJJWxmNrDiva
/ynjyrrbKZFZNyRPA2h3MWUrPiqf8MeVpphN1SimAenLp4AWO7T6E6BLdUwG4yp7
A1A8N6OPgE4QNjsGYl1rmWIxHGJ3oqHuCyAAhBXL8F5NJW62vhkJLTkuLfrfaY2a
m2VKzaX+oR2T0AnVQZMRRTe5cwjrpg2sT865yw7v4NioVJ21f0QYNe7ADJgKzAFE
CsUUkwChdZl4kWkTXXAjvjerarRzN2s795blhYXyBUn1eN7QM/N0S6tr/l1Y/XHG
ps/IfC4xFJpOKkW9ooThmNuMk8FQaFJoIAB3Gsa2wGauc6hY5RQD72W0h1f907tk
+XOld9BbAyNR1ZuFUlgZSp96ut/nqt5oL5UVjXlTTWntgPkoauOQwOC+SjcKxypp
qkzp7NGyuF6bc7iEfCgKSgHdyl/TGEXcRQD9k9ovFry1WIcHGcE7SNOHzAfB2hxE
jzGHA8xQVVxhcMXX4C5zJEyasVJi2nOWOwXTDmAqFmMJBTVbpXQpWfl6sZBWzZ8u
GCtjmiFE8YD7g2mFZ/d0EHFQT4ok7nOfXBmS0GlXDBVpmfEJPqDGvDd+IOGgCKeU
pIpTmIX7LCpAg7cgvOVv3fBWwdREKc5lNlpZ1xUjMVKklECiC+IlmdJ88dMyh60u
Av80lbbS5jqT/U4sxjuxEyNVQdcevtMPyay912C8BJNl6/YRCTkpR45zVL8kOApJ
quJJob9fJiobDabgiCGpntQ98j1h6bNJ1lZgNBSK8t2xn8bmwph/yNuUrtvRPny0
fa/uFsAncITaZNAPvgvoY1fVN8oLDPJ2jHTn8YKXAuM8w3HUGiTB9NlSNANEKK65
0LhuluCETpeI+CqTO/5ka+WzLSRVljjngMaXIA6RWmNuJp74bmMfq8LzP0WwVV30
1ySsyEqsIc2fYjgPybInjfsIFrIqxVrrJ5kroeI9drSL8RDKDEnHqJhI9ilFyd4r
q2BK1wpzvY/TnRh5yRaS2+RTmWhmglTJ9ZVrgE+/SiyKpamZj2TGBVmuqAhb9iaN
6o47nd0yrYNsVX87xHk+8vV5uupL1vnQ25K6s70bSgj4ZfQvA33dotHZGw+0eTug
izUV7D6LoJ8xL76tBR2FQbApO+2HM/NcEoIKcNn4+G8J1/EzkgtPueEQeOKJWudg
oGwVd8Rw8Fs+1oe4hGqRw5MzlcaRFUMrn/xLkCORgkOQ5isYblcgRZDANagcDC2c
uFdoC1SQgHqwkWQr24p1CCKrRvt22TbBtbRrEiff9HAq0SbZ50Kzg4S0AjJmZUt4
/eXbNC3r/W5qUAfAlFZm9jgy3ZxyNWuKKNJBNNAkD3VsB37D4VUwXClLszqhL0wM
JDjBscNWLQ9JuqSZBoJns3RLEuyazS1BzWrxD7pdzS5VL6Y9iPKJ/4P6KWmKWfW9
xGLLRFdeIXFdIcP5lM/6b1XEaEBgms6KVmVCZzeVWzrBZ8arHkFvJ2JZDoY/NnFT
EMy8FN/6vsjdwEFhpUgT7K8buuSShe1fqnBE+EkQlSc/6AMSlHPGq7JP4LTftEkG
2KbZKGEmoXLuF5aEpT2Cu4PwRtmwqauGs+SaN4Xsb4bjiTchvgrD5bwrJeQ/Ow/S
pDLi37srr4d2IzxDByIzQXPN1CT1dFqv5n0pEzMyAAjVuOXe52FixVdpSiYvw8r/
AwKZCakKVxRWL3rTx2ws8QMoqASIdxy22FzJ12AGFeomlQgffk/m2XDoEYzwT55X
yuSh+AOubqbMYmfuDqyEoOHnkbOnvA0Q2yttUSdqGUhWWMcsyAhTst4by7nLwcbh
opvnpGLmOYBMObGFDHXeyZ4gguAGBs7Lu37M4anR/e928hSbI3PxmzhEe+IKqVya
6+OW/3G8UxCNwXy7k0lSrNPJmO4IUiefFsO9I04AfCD5xADGaNjoozBZVmGAA/1V
CF/JZFT0nYp6oyXQP1+FN7EsKg51juaZ/Ny7CucV4iq+W7HCIVi8mVy6lBHJ9MS/
48eT3eXeBQdTKXOycXPjC8/vc3rcaqjjwYAXseOKhhWWj2HR0nnvE2ZPTgTpje+e
glYepD3/2Kpn3aXT4sBP4RHMS2RYK/DkYieOcSgu+lFRlqVBOtcCf7avQDlE4R5/
EAEnOgjQfLO5EdQ8+xdUFDiSG/w7XiQGf6hlPVwvKmQNsX+JzLU7mM0sD8CJLt4D
VcrXzzg34bpgBdlBlv34iKaoUrzgw2+J1xK0avVS9Zff5dvHU2lC1sIL2EJZZ1eJ
SHZYU2DcEIkMnd4tT/rye1sYleTrXsChQrxl4Z0LpiLoNLa7cUwSXWNS5nyPUdSO
8oOmsbq7OAvzQO3kBIHl8ZqgoWE7wpohcdU5S2qqq63GsK+58tvFm0Cy3wZOY3IH
a0PdkwccPMslMg5CfM0Y1Fvk2fz+gG/1IWssJzY49bRBD9QgF5bJ/+hV76VJLvEy
qnig4NF+uQM90tZuIdzt/aCcFDxCBYbEkH3bZ9WIPQrJ/Mn2YdzNYJIPbxxsRfNL
SiAE+kETYaYn8r9AWadk9UUvZdHTe5JBUij6VuQPmm53Z2LpsyjslLatE3v0C01b
e08zRHGibIhmPEfgrWKBjpWL7Ut+Vj+S3fZ2fKdaze7Xj+WFhiTa33gJj93qmfR1
VGgyMLrJLdCbjbqgGRef0C4QXVLgEi6A60ICbDYg/a9//5VQkTuGzyote0lM/jqR
rWK+0UwORWNeajHHRV+75DTeLv3DE+QyLktQWEfbU8AJ2hgKjzcUNmyVeWt6rkLb
NRVGymoc71bPiC/dWTm8T/HFKVgDZLmUmhrpJcMkNCw/fCnoF2iCMeG+kD9dDLiQ
/7gYUT0dIVpIovMfTv1uktVF/JRFEcAIOJULMfxH4P0HhjgnXIvEkC+u0YvsW6Fl
kuWlj08oFPozB2DI0LlrDPFB3+pUShF5Qa+24J61nbVB1A1YvFGBNlKObcg/Uk5t
1S8Q5/tHi0amcHaB0jF0lLFIjBa/AG/OnRMdNhbQZaAz44iTBiNAIIfiUhOSMYsR
zoNa7agH4lBQLxMFglfjeJVDTvgn5S1vvThItidAgNaK0dsJdfMuxX1iXEcvNWXe
bcSl32lNlr6s/EHFl/2GosMwUBQEMRyFMjh6zyln3Wgrm7HNfqMoBAZMrR65OqBz
5Clo7YjMNFw3qFl2MIitSqrm322ZEJvdOHuZjMq7ZLBLoQCA60MbD+Ko+tXug8KV
I8Aov92UVzsu0Kii5CfgMKvVGIAqcdG40gkwphudb/HwAaFYTPDlbaYUhFuK1Pxh
j9uUwW+W80ffvJmig/NqRgMcAprfFQhtdcSXluCXlOURGEV1oixZ7h+CzqM24BGA
cRypSWRaGZQv7B38Wbmr7o+TpkzamgPNaj6Sk0+H9cdGMAThdc6SJ59vF3sAzcrS
qXITfm0gv1L7z0BE9ZukudUEc1vhWTu43nUhQjERIenw1yQ/ymPEV/ELz1GIWQJU
dWZRcRYy+6FjNJjeUZPwTdC1+9yhX21IjiotA/HGXdZAx/ZuJBNzo1sPv9NF8T1L
Z9x1JMamzCEeczQ6Fw7SH4/Iq+fiBTCNQW/mJsg/NKE47QIqn1SsBTiuOtbjjS2A
7BpgbR9KHbBg9IQ5tfpqXFBKd9wWbqUWOK1fYf4HNNNVV9RBpNVIKzLn4xY2h/gZ
fA2+8PIp5YGy/6YN1j9SqNCMThGj1S02qpFBeXZEJpTfoeTi+MBQlpYvdOFtNZhd
xjw/xI7RSsTVBDU6OMxftDMf1helPFRMYU0OVLxRIDxWm+F3XwF6KCV8Xrvi+W67
YsFQcnqRZgGDhxOLiazx5qGwsJJljeb8VisHOJPWRHr2vRSnwNV8CNWLl7+qKUCy
/uCkVvz3oiP/upMUBD0JEfd/6UNbbSkmJ9GKUmwsZGKmNTinhndUCFA/kp56ySTA
VCI0TBv44RujoEGSxU/e4oZOd0wIqWnROscwd560xlWtB5Lmp3DVSPzGM8RvkAPB
lC7lCLP4kb7sz8ufIUIr+UnaSS2sP2OiOZe9nzkcdJpPugMMK/cTe43MCWNT65MY
DBuDrchu2GqaVbE0RAQOPdrbQHTzpThkwV8B5KMYt4noPIcFactxdQCnksMAp2et
6cAcfs9a6gkO2RYyMg51neOTdyczcj/l1z/E0pHVcFf+YlBbBuiy8BNDx3E8a4YI
VFx53pxGvDHbbI55kgTq0fUmoo+Rq9ITvdEsL1egvJLl/eE0fvJM+gWGRRCq2kD6
Av7IH47QIqozu+8j0KP7HQ+APg44m/50ATGWo8fI6QuhJQjrdfWK31vESgV16OSi
VwujvY6VGF/cOpxpKJW+FV8xyiBnTxWrlg2LTu0BQog1nX6H2P2AHt3hMUVLGAdl
nD3Lzdhuspqkoa5VlwOos+5gSbWIoVcF8aGJHQIPw5pNyTK5kubu66COX+zbjR0z
A1Zjod8f+Kh0pyj1vJ4Thh9sWHx1+qBnpKAGaTdecwUDldqD/Xv0wXd2CTvCVLkc
amMlBb0q+Parx4Sup9CT7fZef/jPVkCsgfupJBHJtA0CXFMHFNNnp+x5kHqZZi1P
rTPLvaaLB4FiCf/Y/vZOO8iY869ND5yJKHMjo9pZUYL0HMRFHk3UMhtPBJPBRv/W
vwejOqNeCBQbM0afbbWm2wLYEu4utS0JLb8BDJEbRHHxxSgd7Sjvxdgw7NB807dm
7AbbYFN/VTuqlmaHfOJbek1JuVrpMdHxbMv1kCV+f7iDnjHUnmtVT6xUYYomDrrk
+1laAAd1jj34m2AYchJF5N+DkrnUzEP57N3iT2Fj536HXxEcGnpwh6h18aENa3hd
dt4U6PCdUox/r1glrYjp9Labn8Ud0FoJRXBiGhdoSMYJazJhQkd7VsbWkI9VBst9
6juW4Xk4PPKyNmv1J6SoEXl1Zgmtil2vGz4+QOoMlENpaJfUUBoxdGBuV33XXGUo
JRFzGobAI82+86Fl+D/4RFrcgb1UK8aCxy+nkTOQn1sygvPorDL0rJ2lTD3JMU+o
D1o7lGxJY9db3xkbuQdSHDT86o/6J2ZTIypkuyXL0x5XDr9MlpRBWam6ilg3Yrc5
UqkQHZIxOLeZFOLjVByecNIougUdGWEha0hgCNdlVFtSCTnlq5Rp9tONnWJLhSx4
hhOM4SzsUC//UJjSow2y3dtd2S5HMQSw0dtEcHao/t+B3n8r2Ts4KRcEezgZ8mmv
DsISKSsRV3KhtPzFpSz1Zzva1QUn7YF43yFBWQVNYGmnwmmvlmfNvued4841bOwS
+vEbx6JH9mAxi7NRngSvOW6mAHu9uhvI7D6aWTVtHoeGTrygI/ArgHk8RFNTfWJa
3TQYP5iziMcnbRkke8PfiqbKT15E1SfOIViLHniOf1mf9SaVT1PoL/0UvuSaxrik
0gpZN7TsQi8vRU1RCOGhOHCsXvYq2wzZr7sTUzGg2vcFboz0XV6HQVwLrM5lDC28
3GndicqspaXxEvexfzhcvK6E9Xcp4pDwan9io0QLLL9nWEbcNsf9AvFOA5+hRvzJ
QJtvBBJ+VzNTqvwaHZd7edsEO3VJKOgUgYPdRHdUFHNry291XqE5Z1uiUanNFYt3
c5fYVY/m+B6rh9BBOLY2c6o4+twqdtXTvX2gMve+TNscpxACQFsZ66xKNok584Zd
HfHgunSGpF4/DqIF6qycKJ8/fl/Jkjv0WOgBFfbAlP1pPDL0MygFiThdjcCamOrB
7JDH9qqIZlf/uHMmZZS7jh//jWNcEi5oaQ2k+Kso9OZ55rEKyO9Yt5Vjl+Uha6tr
YyItixN1yOrMgLVwWNLfxatJBRDerBxZupJcNN/Q+xVOPOb0UaEuGjSEbamRgRFR
V6fVBuAzMtzq0WMuwqilVf7RwNqr/qQMQO3lQdgBrjBvRk5UjPRHEeCdMMua2r0l
zIlU2inrRTv233TrTzwLzEihrtkLibkU4/dIgbNNaah0j7sWOnd1c/qC43hEIfWv
Kexah6L6OOcXA1owwJe4YmWHKTh3KDsv/umh5hInOeCgGipJrFiBtMFa+SiQSCXb
x4Lr0AjLMd8Nijq4lyoD0bVaV1sywiMl6xdFHacjvzoDtlo9UVuRQOsQewaT+7wC
GF041gGjT+1R3oS454j4KbnKneCdxFcF+BMRxaK8uDnshp0KG4HTjZp8cjihCRrF
IYI4VG+uTVq7T+rsk5CanD/H6J1mDR1JsKVFszv4CexrPnB2CfjU8yq41kr59iUz
xh8UjOnS/zkD9Ub/ZL7jRfcXmU+SCHoklzVIiwVwepwirfkTPq4jukZ+ZVLccsaZ
gkO7o7CwMT7Z5DYmb6KsgQx6v38ixY0SdWCxrn6uZO2WsoT/SoMOuRta4vqQ5S1t
li2z6DKF+/9bf+2gGMAxwWRtUjMV4zrKggf9fLfnkxD3MKzxrYdA3gdJLr+ObH2T
0180Rl/vqZpDDOQqLJg6GVHS2/aQidW6cQjtOvorjm6NWTdYqxJHZUS4pQ0rMeGH
VzgPc0IXRsLFy7Ghb1E8PbpnaI8n6nAoiczNSU1gcbwifjI8mFEQDG6b8G0a4ZnG
pOGGgiT/q78imQRtOGG0JvqOm3OBAhJNaLNLO7PgVpJupwpEuolgUExD7teONJ35
U3vT0ULaTXFt7L5s+fIj1VBMvar37zUuL7SOrx1zitixvTwnUpTWJkqYuu38e1GK
iHiCKiOGM86GIpZRXJ00jeFA0t1Tyjbvbg9nWTEimCHEL4nlI6riB+V3szEkjcUX
uRw0Y29l5QwqLsWfB3aoO5wwnGtUiQ1spMQ4qUg8R3jvihqpRCcWkI7SFcPKXdQz
NGP5e8zZWtBVD11KUCs1BbMY3ia6cZO5a2qMNjA8Nyyw9MQj7xySlKEk6dpDhE4S
C90PvLBozRsckWPDwHbJ4KZ2pzfIYHQ1TIO3S2jaiMGLPuTmTTjoSgDUkgQQYvdS
1Rq59J2mAGNDjn35UO/+koYcVLW0rY1exWTbKtFeBxB7QpgDjQT7duV4E0nssbNG
vBtzxThOnN0RLPW0la9mEssuekcyh0ecLimK4tLfe4hWIqX45+JAGqrXlQVcugW8
lGO7lI8TcuKzYbXFOg2mZMu6oJegbRpXH/a4jrGpL6w+cUKLp6IZafh696/eU42r
EC4EDBtIXa2n/cJU4gsm5yyWSJk2U97xMcTgeE+92nneX9s8rMoc/96c04N7pPh7
GrR9ysoXMf+PXRhKlml14OxUTCAEQpCFO3ZISw9vHxGKti76gQsnGsUpQkkunHcY
eWUg69PJCixUPl6AcaxhLCMNFbzVhlt5/KKbanRhGe9KE0UmawhWPd5Zt6SGN4D6
VbeN5ja2KD000l7spvfMyhtEPz+vQg2IcYv7pUxSD0UDdRZnFfHCQ6gf+2YYlsFm
AQFGqoFX1HnAGGiqQZXDgycG9IKuzqW76T4S4f/12tPN6kxtcYVC1qlWdDzfmV16
vOL1dabefcgZMNIfm0X2QxCtrXXF/7PN8J3cb7FUbC5ZTWM2d7xFqqYV57s100ab
UJVT7TB6/qTLfKKbu7wALEQVlwwAxynnBOsLHMxJz07JfNA+uOdS33HlIeV5dGNI
7iC+OPoxOCPA9LAdiAJTwpfXZP159GiE2B22pZHjOkopDMbNTH4KW/EsrdAcuWMz
QlAoIbEIuTtpq515fl7cT0Dozjmikr+m+v7SR9EDyVhx1UrRaF3Tw0NZAB79R4Wo
/75mqjWCQOMpMwjllt16GgGnvHCpbeqE2EOgwt3NCPHZvV2BgKoGD/Yx26s/IpB1
ysAFzJHTL+l4TbLB2REq5rcEQz+dtR04Lh05CsAm57e5SvV7BZrIgbRJHXMzD70Y
RTTQPeWyxraHi+LKHh5UqihjNR90FtCaDt1/PD6HM8djeo+mcLC2f3IzcK8VHLYd
P/5Zcf2ZlpGfU2uDrKDrKuf0KSzJDpuO0qKDLMi4w8gKcHZ7EO/Wesh9uBnJseJe
oDzT34BwSEvjQkeL1g8Nk+Xq25z/besOWYZ98EGhrWtFDctFfj4AnAlyA5WEF9ix
d3RpHOzM2fkqcBVzYpQ/xQndVY5Wvdo4s7CB4HM9AhmYjP3FTfNPZdQQCrbRF+PV
sTZURtwDab1x/U9pHiT5fyig22gJFuMr+mImjausGdiQP8Ahn8fjLibss5ugywFn
wxbj3KkvcVnRw1uDJC5LP3jxoYGL9hFaAQsH4oznsFMfBYRwMDpFHv0s581XVqvj
bfK7Wa0ilTRw8e4soX+bU+wZsDxwLuDnzsrsHyxsJa4MGKeVcO8OB3tpkyxgMwCS
RzZfBy9soSRsO+xkPXTkMVmvWzb063GwDYPhFtYRuvwMQGPVgnGCAg7GF+C0dIwn
j0y8bXJEhdnvQPO23gs+vE2vxIptVgoi7jsDTOqmxAWH+23XpHHLyddCF7o7xlQM
YXqRo2kEsFWO1Ov7OvVg3D0nu9D37kNA6WkeFcYGzEmPs+JeCvHjygftAkygUXcO
QfDgQb7fWGX0gf5PbhpS/bXKjeVwZcxGUy9zjfTn9Ikej8uT1X039Z9cDsv2Jg0r
sM1wfatQv+HDvAyvM2DVWW8vNqCvGfTNBMNn6VfpTWtP+UxRrhJqAV1C1gzGxqfu
Nzn2NGceXq+P3CbLiyIeWX+cg7NnaNa5tFUwPZaMbdN1D9kyl88Uy0+4SwCcgpGc
HaFZ+ypy58eCOogwhiL67mIuPfJZRJkTHWlDIPil8QLbZcR5Fqd/BAxuM77SvbNL
8vV7lO50na8g0OgBSn2ok0wjQTqmo5+Huiwka/K/Z1Btmn8BJTpQOrUoRr5VYZU1
yIXtGLINjgk3Qz0huMZnfwHkgMcLGVkO3jFslYy7J3eiW4kuwMul1MPXBI1wBML3
ASOliavgiY58O0Eu8TyHyHaNQ3T5HRjWRecJvXMHG5uXhEesJgYV6PqF0ADPBL/o
YIi1Qsh1E0YQWeR5iBpbQFMaLAURj9cTaV42knYuOM3++CAUN5bj8ww9vvXCahs0
QAH74eNpSuh/guf3q+wWeWmwV8Bgjayt0A1by+j0YMRtCh1gXkEccH5N9Wcvmn3R
FAOs6AJR9vVt3HHdzeBJEzMUU4gDHrPcoSuLmU9VgqZMnmPr+pKfBjIXqLe1jmnT
kLTvf8hmrtcor54gyFJrpOCTpSIcLMehG/ypNebLwMbMDaMgrVXbn/DphsCFZsVe
E/h6zc4YA17EiFsWmb71JxAwomOvNoDyM29CrOz5xqtbyQ9R5+XHgepbm679zd69
sGlQJorTfJCvhrcUMFq6LzreOn5yjUVRiYLmlaAeh+Fc/5aJ9gmFkmNxDQLejy0T
K1FLBYJos0uWPuH5Tb32V4h1XB7M+CG9fq2j9SYHWLpJKy+vsBb0g2mFxz7+62bD
qYAJZP09LGZSQ1Bju7GTpvmM0Xfqqcj+9CiqjkOQ+E8sDFuJaVD5ug7FNREWfZMY
S9JWiHp3brmoiJl4GlTFzVzs4kolSmSDC4wk4W7egG2vdnLmts/A5xOOfk9eSR8d
p2HguBFaBgjoHz0UyqJz7qZUe3mv/czc9hX/qsT7Gyrl7c1lh/B4r7FRYWtkPwAS
5y5f877W9kSVAe8md07YAFfBxJDFruT/L7T7mnv3ZHfrOFqkbK86tx8ajTeWzDHa
ARZlBy4xsE30SF1MZhFD9uak80e9dd5iRNXJ/kS7Ii1uaL19iZYggnYlnX0n+mze
FhEJhutF/S6YX7mF5yjqAWXGNMRgpvifj7ZDHwZGAB0sx6pWgOMx7H2fg3vDcoao
ELDnh/lVQ51Y7Z1f1xgXK2zYk9SdDXPHINT96de0LPaoE2GFzCzRf2fFV6/umWod
XCOoTwaUQcTywtQPXC8UNDyNWg+pQMPtFcfSZf9YFSXcExceKRMCZAJN9RzPDHsn
DIYSbsOc0Y6VEQ0jdkY/sl9kSnYRkt0d4hNJxVJ4WEjgBbUTS+/n3z0WCSy0yK+E
gRm+E8ClKgl215bA/zeWuJjSkQsmqFjiFmlTvrjN4dm2Hu2hB4VCaJfGTgPSw18r
wNdHc6W2EGfx0PWUq8hr1eJYYdgCsswpZX/fJkIbFoAQAV1lohHVc68MUIPdsP9y
XRH6NE0UeFVWwA4Eg/pel2ymEe5HC8nLFKQ5DaVXp6MRypBcXSsv0XLlHXKayYGR
RdFOpX5XF2aDYD5jT3yTe4+4c1gRxtk/dvd/IOU38rxY0lIeUg8UkM9PYxxWmHsC
e3qYZk32lBdmV6XkFG0DHh6VVfJ13MSnXtrvOmlgloxoNMDx8/j6a0QeA2oHbMIp
xSqaFF6N2UIOl4XzUOR/DFO7v4Do4uvZIEATRL+Xc46OYDkNEkRvJu+8uBEKTldR
Q/suEA7p4LS1wqlT433jAKxuNhoA5PfjbaD0SXnrqpLFWdJC56fXC7b2qpl6UIIL
jtdvXECsnRiBaBjZTT6wMAv376PzC7cnkyv7NgtA6ktnoej17u75Ta5ddXbMPutX
9+7tjK8GmTOGYgmYay4gugQYHmEIKIpFidsgxJe1oU/l9sStU5BRUOQ1J1+Y3o3K
JAh6OTeUwe0TCwTNpiVnM9VuCHPi7E5fyC2zfd160qaFyzefH/4ePnKBAP86aKea
+GyAY+IQn7d0nDLTO2Oi5QxSUbaed5DKRKl/xjuoaJ4=
`protect END_PROTECTED
