`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pBAd5Fgogme6pid+JJZhNlRaDfZEzUPPhY40nPSTBQvlvxXLVEhbn7GaqFJX94vG
lt+pC3ceTlxdEeTEtn2B/7qcLbBvvFW86/EXLeyXTsa6JlFnqhnimViDbvUDD3OI
DjBhBG5aDnl7jHY6okM5Viu/ggTqbE9pYZuChoeGPWUijAeT4ekduOECLCSxlPW0
ZpYADmRrx+jvlXRWJcBGySbqmGLNNAocVs14ZU+U4PxQCDaqMUzBnKWSUU0zzP95
pUE783pAWGPOtXvEQ6LdQM0XwKdKjIslWyvCOnmYOj7uSt6vHee7XfF+sJqpX5Zl
/NPQxI4KbFFzC/GBLh01j3Px1oph+rCxnnODfydy3EGNcJ1gouZO5z0IP1b2DAJT
wfd8jtVSRKv/TpCTwZQe/yzKN5JrLhF9/1UMjZFRTSWNmmXygrLRWEpbVKKlGqmW
DMq4B0zoWHFubuY8mUI8zg==
`protect END_PROTECTED
