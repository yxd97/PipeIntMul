`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bi/gBVMKdfPzqmbRlDKeKOu0PLGq2VOnvJoD7U8ktPEfSviy9yRn6cetGxCfFzTh
wcudaDbTpeYfeU/Bf3/vtw5slp/V3Zuf3XpJGQ147upWLY+xH6EpuG3LVxfQmhx5
sn6grFzWeaDHEnKw7I1hwnh8gB5K2MM7CS7HLktcY+B4eR2i9OmJzGFPQOxe0Hpn
X5mDe/wV0MSee2CUHwlxYV6BFkuNpJgto+YaI8AkKZL5m6TeftPItF5LeTWC9bba
Oqa5oIDyWwIkVWhooT0OXYGdsypFYAgG6BkzOQw5baoLSA11yX+b/4M4XEVAktzW
diLM7nO0rDZweLQL7DCMnkNO5XVflyTb1d/AEC1bLvJfOvIC1vEyQDoNVTM3wLZR
J63GfFEQ5V6j403+Nn1SOA==
`protect END_PROTECTED
