`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Am+fwZUqp6T3YHQiDVD/IlEP52h4Ku6/A5QM7Fq9ikUhOUMCWX88UgrEy4IW0jK
/SHCYWrn4nerxvNSAO5kKEbXyJZE0Y19QCLAO7wWTKnFY7KyqKdVqQTf//SlzioD
2GXxlLUkmsvmFLARYWxyMBmNwskz8xjVmsZlpQZA8fgJPzwOPzAgVc706lM0IybX
XqKoMku41JZ6ZMJVhB+BBkjonkQxmfxMumHQTkMKA8CjGUNNdo441ZGO+Zs+kWt0
+TW5O6tuNFDyoEC0PIgip5AsrYF7QQktH3kFUsG4WX6WFlO3Uy5dq7m7Ca518aSb
ua7QU43LzywPTUfu3krA3FoqXQlbyddtJYMHL9851BonNsBnGupRG/MAo1KVc3+O
OZUxNwUsT/wlBVfKRqPioxqV+PJanBSFXdjjDvxNxww=
`protect END_PROTECTED
