`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GNo/QkvZuRO7dVS3WzyHMI0ZdqqN2a0nZl2140CUUcBMyuRYcT+xpi0EG+jdCqIH
7H0iNj7MTNDPlJz0y2PSUXkt17GuC7cD7cJMlOJAf9eKEgNZ0qH2dKq1HLmYAVRm
hQZwbvG08G3uCjpCzne8xTfVA8XJoM6gtdbduDRVDRRsyxVfwFMyZIcRxzQeQEQp
S+cS4ExnWYYvyTOpYmt920AMiLwgunQkef13VBwsa9RQAKR0inMuWCpyZbbmTrx6
DT6wOc7IanOjGk/A9u1Wa4J1IArh8DbRvs0wTdoNyY2uYzGOZ/L2uIjeWBc71Ste
zjrhLIVujw5zfQ27/bFUDZL+BABFKEmj6Z/n+hLil2QhmKyTXnTAL3rxTsOTgfJQ
6LpIBrJqfnlXQ6CPEhBrW9TqLobMPBLdjg7/8iyikSw9DvjYPHVoYP0avdsjSigX
8ynKQF8dBtGVTRmxu37KGQLIFyQBaqu9MgkMZTgW7yWW9SHX0JHonP99/juWdU7n
RcePdOlQmMbKQKXtPzPtymaYCWUBIO9Ivn0zIIjecadx5hn+TltfXPJU61Sxbcsl
sCf3tZQzYIj/zcHU5/MRbmyNjBzv/1ccANL1clpVScKhn0sdZLSx7rpxGZPLOJ9i
XAcRGsAzjesxKswdm+lqDNjGt6rHCYyhXZzmcyMlR60=
`protect END_PROTECTED
