`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+rC4qK7UIeKaPKgkusX2ovgHGNfCYZDqReDzc2N8s5OUjbhMeVNxm/Ljvfkek36
JdrnnuskqWew2/yuEaFZZ5KD36lfjRntw1vubBgFz/MeTal/Zd5zgYag0I9SFXi9
bh0/lIW0/8nSXesFClyvfrkVxW+GHbgB9qNYxsdeVoc2+q9qTG1mj8yZyK71uzZ7
4NZIh7+2TD15SAlZnK03Fd1pOVNmamy6zO1nreWGEjazWl7lmEcb/qdtG0TavOnz
ogBHLH2SJpqfa64V4dG0/k6IAHSBhTYht05duuiMhy3WDPfC13ibS6qj9KOCk781
q02NKktYvWQfrv/1XPoz1pbxjiMZNz3nqxm6mQIzOIyyMGxXFb/Ulh8KZCcNE70M
Jf4d63BVfTLRVKlYJh8qBHTpA7v4HKHA0RGRSdSDqQGRKS7R1D1HSUvUzOvWG6gI
UAN8tpkmJbd3+vQqrpQoooutW7mKZAZMtZ33xdBUtdwhNRUgY+3tXR1I5YjyxHgC
ZyeR/yz7jBkYND7tm5tAcQ7ehvrpsSgqcM4LEGe7IW0/bBd6qOeI0CxCgM4MXQIi
1/pwtCZ6e7JBpGRJdC0v3g==
`protect END_PROTECTED
