`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JhFlFGOuO65xOMQ9JKyI9yvxaWL2jwT/eZ1fVqqL/uwELsO8aSay8dR07874qV1N
HbJjjuOA+xnFWhHyiSBpBKlOvYKKF8OgPvcIA0CgH2wFE9A4uEUmYXf9kfkrAsd+
KVqzkokSueesn8ieMTjrhQ6/F5fYM1g7WI86POki3T4bpbATNOaExfvxtesOt4Hl
ADarvinn0QWSwrCJf5B82EArShdj6EnEQLIjDkZvJb0jM4CoijHwXimSDldA6qiu
WSUlDKHCqgKH6CsN+m6M4Q9Z1o8RDZlGyi5JZwbN8/A=
`protect END_PROTECTED
