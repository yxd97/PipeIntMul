`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YrBnyzf6WT/OPD6mDua1GHPaYtMNIGKaRcsfl/a5KC5Wn+7lqEyk5MDsEIaVm5uU
XgF/u3XjfFce2NKIbS8Zd2pZcZYs6IwLNhPwcU8diYvtr2I6NgFGm2rh4NLU/sI9
vYFtzKUAOlo5qW2B2bFKuCWLGP+4tSLJw/N5OM5Qx2dAJciuo6Ew8QVorhCg4fqz
j2EIoseyNQgreBUydcSD3cv4WMilqH/Y9PODrp26VnA4TXEdizc36IbZzakRhuUg
Dlw+R04zZ1mgofRSqI0DsOne/q4/sMRN51ykLwsS7LgrQoduHaDwF1D2G7NZeC6O
5euVw0M/yRzhTZLqPyv3GocynwTUwIDypQKePFHCWJp2CzwpzNvW5PyQE6LKPWAs
u7pYFfx+K2sCEHFOLQS64XBBKCOOZs9mhRuhxy+wjFqWM9mr19sR8KTU9ZVgg99A
zQ4wovq+jAvmrIjyoqkAHK36DfmggGvOwnHjdK/hNt1e23XJ/9SWI2QML2jqkk6l
zR/Yrbe+IRq8hLha0ku58IkGRxex6DRHpMB1lyeRLiBUc62Cq2ydCM9WIzyamgR1
VGDFfNbiM8AS+uJE+p7L+Udz+UR6W70qkPamPHtsvrg8jiPrIls1PqxIyttxtzrq
LBBpUHIpTHogI23FdtM5w/NcRWsdJs4nxLQMzY/xfzoIchPtF1ZkBGWQXYo2zhOj
6WILZh2/R2mkzdRt0UCGXHcpfgyA9xCYd5QIF2/JzwqiYMJSZs789Ch3cjuSXOQk
boFcwSySPIKbwHNhja78mKeZFFl+rCwr6oXxA+1IAzmrjs9fA0yxMCavQWoq7orP
erlPFjh1mCuYMATFZSnaTpt+USjkvngiHEexwnp+dm/vultGx94RnGgn1IxQYBVW
NxK82PUBg+K2G8diGqbqg8OriyevvMGoU1kbvYjwZVOPvYXU91zzMBhgL46uxqXj
czV65esXJKUvngxOaGUjQCat3KgpFvXPNdsN9AEZzPCF8m1PmTL6XBUPs4hWNrCo
7z6thWrowJhzmzPYqZeVhEGLRqyJ0WUiEoEyUeCWWu/xIc8ZheVXfAsSNLQjTjPk
xJlv2W7l20VlY/AzrrP3iP4TRkFnL1deDcRCQrqXrD2e/1XrzdMjlPf1Goy7BLIY
DLCBsYbpR/4zcDLZ+LtEuVWFn0eaPwnQNo6JgyHZxPnkbGuFvJ+LUUyRuJVBbhhL
k/149ZcBJHLH4O6dBWlBqyHOEk5Klmx124aaIqohuHAYcxmxDAttxJvIdMj4uYDU
PE1r2l9Bs1lCHtMDmwj2+BULLc9qndZV+86eCW94mR958G6bJn9djgC65e/hrSW4
ojOYXoLyaJ0oYa4ZiFABf0Nk/x7f4NjObX9fekq92WUOvr/xOBUnzozIJrn+VB1x
6dO4IVhasXeaKmI5Px9oM5xV8mAeUEVcJ4V54HcU6+DgVOluKFTDZAHI5Wh/HcsM
OrpKaYgbTKkTskVEQeMa4I2FiRZQM/j3for2K5akj+QOZFJ9g22EMPo0eE5hYExs
vOktHJy8IKItytnRPswfW+IDg1oGuAd5lgbAvJOpf1WEkTiIdY0j28C8ZzlGbpiO
D1nTOzePGG+rDt7qs7lFuFNYHvQmwkteHmyLhe6qXyWwoWzIwC9KZdLEeZEfX/kW
ywirUeRjHyuBYUMYvyqppm+1IHSeCPh74ko98jR0viHfwVw/6rqaG+4tKeEqwfvS
vMtKLG36NrHpCNp6BqqRfAZzWFRlTVjB0tO7xhTjjXRPH8pW3d7gXFXZbHJv6sH+
h0IPVj4Wxz85WLIBD8djg9kemowJnbP0HFZcwyLUe0ZvuQ/jJr8/syuzPqiCt8wV
O0jEac4jcE6wY8T8cNJZMpn0QG6aUSmq502f9s2foIU4/0Fo4bWHMxs/835YIgIH
gGsYB9boii4ekm/wHivlTP7iP/G3Cj93Zg+PaSGpCJnj2k0meZwxq7/7aPy8ZXtp
gWDO6VI2fjRuqtbyW9K6ZcCiBn9D9r3Ro5f2sofkmxrLHIcPJ1V9grS+/ghQLyjq
v0KsFcqc1SftKjoQ6297yWorHi8Cqx7UsrklCyAoSE29+0dnrQLq93TOrdZnRU4t
bDAeF5MzVq6vnbDbI0S5VIwWg8CdH+JwBSELpMEUHNU1ubQTGLU3Fo4Egy7dWmOz
QWCuvmwsEqaBbVT13DYHXEKA8Xpu01XZgX/OQmDWWdBCkt0ezVzp5Is3Q9TrKcOB
LgYt/eih0JFf+SNZsyOXX7+9herbgvcRHhPhhubpcjXutmA72od+ProLifVB/x9f
UBXtwE8CItbUv4rqMxQgBTQ6lUrYrX2q173fr9OwjreU4cDaSFpZuBmMv02ybFgl
i3ycCaK3W2fVgVWXCfGKlgNnqLfDA5BZ3ZPH2WgFhQ8QpD/Z274z7lCq06IOL25W
o1Pm3uOYZ9q1H5ee2BH2NhHH1rSZxKMySA/2ezrkdLAMY/abnnz4O1PBdfWqZFll
1w7ngwC33q6cB6scf8A47nzB7iy/yojb6VVG28Mcp6nIn/sIvDFNBhmIUb4PWyEe
eKGrC7M1TSx6ALqpOavbMJvw6LnH91OwPsovB7gAorjH6CBdTDIKkyjb7H6jLbiQ
/nJbfnUlsyd9OEtSwZP0MTYJDBT5mHTBAD6iODZdb669kCHVPCmOljOCUXttggN5
ruOeKgHY6qNUqfaylSW+hwwFH1PXAqyYsvfLy8Q9Yue1StjRB6bPDQ0SHAXw0bn8
+prehSS1Sf/l29nmyxh0m4uRheHN1PuwFTftsnHpMMNBy45xFWd9vrXAIi+FAbUg
sc0NtHxhnHs2FGxIPBQ1bkTaz9yw33qOnNoMGMvJ5xx+IVGBNDFLh9wbCE/i/ga3
x6ucknaRwigRGJT0VdlmYV7gLRLb428WpndZCxoQvxuzDba4QBsK10XjkkqO+pHr
mrHXJUQXinQSGvKmkW+tIDwNCn7Xm08gD+5Zy9jb2yrZQvLOZ+I1RX48ButkIQnZ
hcdxeRTDxDMWWZo3tY9Y9x5p4xyfMfvn0rK6VCsHE3Wr9XELBSgg46puzNxOavss
Sg/I1tt39AQ8WMBDhZcDCkgG0+H3G6bYuXi4EllyxjiKZxuG8z/EnzeIjlbzpEbu
KtTcMolZGCG7tOnhoflTPjs77po79tRepjlhdm86uTdGYZvNL82EhN5/54C25W6O
k5EzdTPnsqJuW12RZFSHhJtFF3JG9Mysf9i/kojGkd9mNXE/jW7p8/+ipzcRado7
y/IUaOU4E8OryL6ynoJRpq8eZSn3PeRfudID3purtgdqW2o/NN8Rw5WJt2/FonjW
7Py1EZi4RAYncAA5qIQ3lkh7Sc6A4+Z0/YF4bIcu94SjKUNdIGczBxqVQsMFgKZN
qc6jOglgDOZbFubLbkv1TniUHpZUTeql9JDPPu9VHPRjsNxiOC8dQgnPSaa5nOBO
nGyxHPBvQUOrh7h0q7c2og0tawV58TIcGxT0chTS2O6e0l5o4VXGI92jOrVvxBI2
vx0zZ66lEiAEjv1NGAQO5M/vtJkUBGLqDmDCk5xLErSyJPyTWAFpCo2MIB9q/I0w
61RE8luIHSM4JTjSoMKW4/Z2DuWVuHB3i5pqZPsD6bMq6Sm8bMTdetkvJdLasMTt
tx9eo5D56v3ZlSJ9nOh4jjB36BsFN1X2X0BBvFzex0fphNj+kFSrC2h/+c5r1gs4
g+tvVQzrlGlURygZROpHFg7ClxPAx6I2bp9n3UGoPI9qquAm5V7ULpSbFgawG93/
Ig6lKBkLdLBM0s1W/7lzcrieOxpI3liBdFukNOCiQk6/z9EkHt/4uTVFabDxLhuS
eAVHRP8SQdnKgS0UtldxGbXtemkKhNKRLhrkgSlfjBws1UIpXTgcxRQ7lyODHoOt
UsdmlDrbXmFne+AldiNgwOCiiU2pbXEp1xyk3kIpzrVQ9QvstDDrA7fL9z+XuFU3
X/GZOp7oyb2T3YyRuOU3iR1XaaLvuO80cpfUvHtQ0zzryTHsNUzbHk+hyHM6lMj/
mjZMSKLQ2SNm1naQ5w4EZ9D/t12P01dXUgWXT8x1LbpNsBbF+hy4Qy8iW6xuDwmI
/ZOIJVztGnBS5DIgg1zfGyAYSP4OgZ8bn+qf5s0aGXzKiR1m3kdGin+e4N89mfWV
n36CMcwKnmURMIuCpCkLSmBgRQPnsiprhvD6XqBUUuWzozAcvVP4aPqIODGDB8aX
LzZER4BAvmNaw76x+Wi+qatym6UE/CfCXdLRk9PDWmKK8giD1DASufvTGoLfe4DL
c+ldnTLPLdVxRv5a07mn62lCExIDe/LP6cgMlpcwtk4thwPNTVfF2rNh13SQN1tL
EuCBMA1p0tfky+d9jAS8hlFR7S/fj5YZtE6PQeET3RO7MFLqHD//eLYxGj1N/wu7
ciCtQffMOhbIsDVFOKz5vuOX2o4/b7bSNOqrw3KApWo/Q8rCcFG1l6hgSB9ACxyY
KizncZ22vCEKvpeWQTJvFhmZfDvrDRXv6oxk2sC5nLPP+s1dPfgGJ1zXhkVJqNGj
YqCO0VJhqJl/KnTqsejNtXofefHOvpA7mhM4r2IGKECridKMHaY2lmx8majnaXYE
6l7qybSyQ3Y6vY/VWdYvJaCUz0UWlE8Bg/YgI8Z2bq3vhFKt+K114IZjeajovk/z
JfVq+m5OM1mt0z2dLFG67JcV9Dw0JD2vq8KYT7BxKOOzD7nmiSKMR6t4XEd+inq6
XP1JjoBzg0Sl86X32vZRs2YOWiz0C/LmWBXTakh0xkEjaOk8J3WCxritkf2EQJmm
K2gqkWau/99p9C67w3QELCLwy72iTTMzumuzOSsFUejGSXUPJs8SwFdZ0QLQM0ob
U26SHAnIFHbV2/vBKgmlFHmDTS0XkH/kWou9ZUF+UKytegAZYa2pqE/znDHJKm2r
MLKhYdFNuXNq5DHyn9H/xm1f2ovBs8yl5yAfO+GrFVWHEy2lhXpMVr4fICc22kOz
CY2Ktm4Tp4fhvqtiYSGAlTPOXjRGKqxcnNlYPqP8kFRd1BMSnRN8ZQFKWmE95Fc3
pu2D4vZt6cLjXGCV+YaEw7Lqtl7xxmiqH8V3WpA6u/Z5RV57ONtr+47QF+FUy78d
+7VD7WsHBt0UOlvdQBMvkKZFYXKhbS3ekyVT8HFtA2GXisHVra/r6/IiAd+PKpZ9
tFM4ZoGE1ULs+zc5gQUGiD7hZKIFlYiX6mMEcBoRmFRp/JBIeiEPRlNI3npbA0tP
I/Q5dTkrWhy/DNA2qx1d9qK0JtoOxwJhEnDzJzJfTivKQZbxmli9ozphzqHrV3N3
Z1XzRVmKjRcetVSNA4CPGepwW+1GAf7gO7R5X3z/Z4brjVEapUELL3CWyQ9G85xC
AcCl2uX4XeV/hKzl/G7FRx4DMz0efX77ledBKZDCsLmbLOX6EVIl/fEKr6LqrxC4
`protect END_PROTECTED
