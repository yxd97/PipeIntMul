`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H5MJEQB5ujS3T4k2MRJKwyPGIrjd/AEPlnnANkgkna1Qxb/FpYOopS8C+azbeOiP
vDPZAVStr0sLft8/xeHjo8twfhFV96KIxSTQusg0QoGdV5o03tZFyCtTQtdxi88J
xF4AGaWnBjUNJXJPDqlfyZOpjvjiaTpoGU+okVUXxyL9WiuhvRAfjQfCtNg14o5b
/6wZKTqVxyu4SUf+jacMyr4A8zGko7PcJcRjwTwmWq4wUSc06pwC3pCgqbZk2GP5
ARJhkXZPcJvb8MBIg9zYa6Io22GRnHsJakGnxze2JbSJNlySrDjGSjE/D/0OVT+l
r0xqzPmthuQwjk/CdFYuRUMQ4n4GIqrWLdagfcpZD73uEM5CavVH3ZxyNI+ryXt4
XPAZyzKJsgGiMj7LHbm46cwW5NiTt24gEa3c1QEpAdIWMpWJaBV3uiryly5pjDaH
ZSiLFkqunMpHuHl1UufyejdZ46XpnvYq6zY+O7OElX4UAa5XzfT3iBoOld3Vkxo6
TOoT49GgErcPfPvb8IRnnIUBcHap+pe8yM+5e+e8+wnI51SYXpOI7Dkq3wLzloSg
PjatHSkpRWft5T903m0aTGmRIZIKs+NnuTF0iOpxKONiNXMj01yB09tp35QJC8nd
e0Tr10BIn1Bolg61yqWEkHG5qzu9MM+IMMzSa3816pTZc3tvNiX+/ah3i/9lknw9
94ZxbE4T78eCsBfS/Nj2A//1Krn6DPS47ruzIm4+1BkCCK/IqmpmT5CU+In8iBdz
9aoJB+I+OkW8Q1nBQqOy7g==
`protect END_PROTECTED
