`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e0yyZmYtU4DrJaPzJbq5kBwFX8w6DK52KhTU4oBPxJhSdQTFXHZuzFQAexRcvHyJ
J5R2F4vSAXlzzcn2UoHTEL2Czuu1czbG5gwXDlBX38C26dQNX1kFG/miCHHuaoQA
wloPhtP4avjyJp0wcUdEtBV/DcIF6+yx5YMfeybZEIQduSjKBdQQqURWZYFw3c2T
GwhV8O6bPho1/uMubzFlcXxBZCwlMsGD1tTP3hm3oJJ5LBPqP75Qk2gBl7ZwUKKw
5kTF7tNN7WIG+7lpYWje4qM47/+BmIC7Mm4Y5C/KlCQa3x+xC+WqkDFjG3XbYmd3
JlijsMVeAz31QNQURo+8bw==
`protect END_PROTECTED
