`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X9X6OWoTrOgFP0MhQhDUWP+uR0+n7MuCN+zy6I9A9i+NYeYib9/kc6hKiOn0yw/q
mTCmD1Sbtb6nB8VBBrEK3i+P7QjUKxJhRs8IinbmBmxHDKENkHrrsa7acViNnrqn
4f7kgql1UvsgmLrkhNyoYShuvijgGGHYKkIcqRp+wCZHrjnyRCA6NDYPr0Bphm+/
LE3tFcBF4Bn+dTbPCo2GFcaieozAPZFPBQTndiYf63BtGqunl82m7G4xGDGETmpB
uHzgJPv7jDv+Yq5Ub8KmdsZZj16/4tZqUikylejLrmpZLHTBRoS8TGs6dkPKJStR
NMFMks/lgX8FNm1Jhpy9h6U893/L1QhQolLGfaWFSKk=
`protect END_PROTECTED
