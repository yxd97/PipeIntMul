`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6GS4plnTaHkyjdtG6Mm2b40qd8BuX/Lwbsp1lVTZvo/DxC1bFsEHMlpTP/Gy7ugA
y2AXa54He8b0HDgzzMw7lj21TADoR0hPnIfzi/69SH+D0BjnE5iJveUAoqIJvUh2
1HApjTVlMTPqYFz1ebBqUpeN5n3eW53K9yyAgLJIxHTPVzl6vsCIzDaR/FTdFY9Z
4blLjObTma2Qin2pluxHfpkPjo7BBi3fN5p/E72RWT1Jv3TyqidXXK3ea3MYWmyf
YAtOGrPZGb96y757rH434GgjzDXrP6MxKucrySov08zmiu9eoPeKW+uMTRAm8ybU
69C+20Z0x1AFemi8U+ZjKz+2WyXRnJfzYveXYI5zqLpfAPNxnwvsEgUcki6zvm8C
A3LMJ1d1gKZICRTMk0aq4DFQ7svct0LtdbuwD91VBdGpwJgmN91YqiL6YuaktrCt
xy96/4gisMfZfcLz+h3PpbZ4xToS6+yWe8mtJ4ni4UYqEOY8B0Jm530VAZrt+p+b
`protect END_PROTECTED
