`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TKgtJhp0ngVpjZXqC/OITds+XDTu0me1QeLwhWN2/NrEI0lv9FUHdgrixreacg+G
5jLYWZduiFusJkwBS6s1HJ+A4xAnGO7qH4gPlM8mf4QVQPIr4d5ZwsKxsXVpXXFT
ZKsdAuujxyMMexc3r7iuFfTfzTCAkqQSYlPdkpqSA+HNCqVstGWMOKJMCDqBTUUt
74YO26vHjUBtJ62mD4Kj6NHNRXzFS17A1cBLMP3BLaEVcvbaDEBX9OCG36ufgzFb
UXgFykqW0IeWjwdDgmA/vRpWE/ObuJ2UJStcfFV9mB7nvn+mpis94ieFa1dWfOAV
PaNkGFYCaEvXz29+UeO7kWORz+o1ptf9O7551LB9mHBdfldUg7faoNYHcHo7Ivcc
Ls152L4i+FOk8t5Q8IWqf6JP5zpTGwm8k+7P/zsDp5g=
`protect END_PROTECTED
