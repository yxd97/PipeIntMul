`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aPabBzrvUwz/W/uGcJTgSOyMa67ihWI4if3fVpxz38fYCBcdA3UvVl4g0r50Se5I
9xb8117Mb9XUG9VoZy9ry7kkPJQZ5xc9+8nxeyDF2UINXqxzU4XxAJnqEcPh5E60
rRqi3AvDgFML7GLK7+7OaxEdkxrjy10PRiON1eMMeFchZzHsjSkCnDoxM1oIVuVg
16uVVNds4f6EoEmQHY4XdlLRIkwcUAfgilc82W9Lhu/qQ9zoJEmJJzmeLoOTNeJQ
eMsBeqlKAi2drlWSzfpYqQVOy4SxNVItkcQV7/KAB/24nnT/9Il8My3d+DC8D90k
TLy30D/NXPqCeUDl/Y3kR9e4KFzKWEWBHn4eKaozxXZ1hMluflSPGCL6ZyjCYvjM
GI8rwoC11/UQOD5RiIYLlHkN85z+kQDfYUc130xDjjgtiXWytDUTRNTNMpRBDQOj
Hg4aFHCqkkgvlP0ZSoAbcWT08D2D+U0kqdAPnR/NBsH7lXC7MW9W2nYU0DsEGlx8
qu+FKou+w8zyUIv2P+KYs3ecsLRH4urhXhJvhWACbZ64am4a1QUMoJSb/mYAQbP/
A1QkiQhQ6+epO5NmYk6CRrV4QUhH+N5FSOiwylCxeigXDzsJNRJB/DVPMpEQH7SU
zcen612lrmRdcjeUk2Sp+yafvLc2XcVwRakk5fru2VW6wazpaXN9coViaTYCqQyF
8c0D5BYeQFR8I0ydkq6HfA/HToBo16qW1b1YJAOGEP1FI9Xf77XFZAfQH6zDkuWY
p4p0YZu4fdzWOWrBSwJUIfW/Wnqvx/A4umMamrPCAYV+Gz8exkmZ1lIoLguiNOHS
ALk27Q/cwtHhJ+x1edrLwpylyKeuiJPEO9wwdhq6RSion7EdpRUbRYg8it1NoFtQ
jEJbWDNZAT8TFAswK1LssnzO73+ZFvQ22ZJq4YSczlAB3uUBL0zZbNVuNysVi5YG
ERd+uf1zNj6JoWeZysIqkn2RfGCVvN6ispuoqydAw8y7jKHk6vy/BaUN02E+s8of
rXfzQP+NsPDrfR0W5t1n90S73Edr9mNTcwQn/ERSJXIRw907AaZDC8vmpWfXxUwm
+m5RyHu8XxH+PPDRDqa/oGXxOXSNrKeZBP0En7iDM2IdfL8CuX6V0Ig+BA79S+Qi
KXW7yIgFhWLRd7OqioBEECAw1wT5IsWwHkEMhQPIe3MkX0IB8z3RVdB9wrWuWPdm
Ah964wcoW8H4mo4yxRfPNfaecqM9YYVSAi2dTJLorvwma7wTYpytolbft7lxkoPt
BVt4BplP3FJ0oFRrlbGBYdgr5qqP9bjsoPK5dVtjGTUCRIg7tNvEwa8m90k+fE8J
x/o7BdUCgybZW0VB8Rd1SoJS276D+ui7NbIFc2K5f2FkHlVIj/Tru4Zw6WBuvxwB
3q8Rlg8vmWsJkcdJenGMq9hADKyAAVX0j4kD9Pklc5MFkKzoT1itfEzzt9I031z2
l0Nhb8d7klopF3QYdD3fB2ttj1l3ILs8EeO/TOh8VpVVzSAczJtRH0zkIpFVLUlj
soCSrfu+6uBh3RPAP3PirW4TRpn2kJcEcdZA+a8rDWYzf3x1Pkhtc/p7eXcpBbM4
OxqsNLjqYuSwfOX1xVtdXlw7KOnGC2aZ++s2CZmm9zd/Sm5i32bLPsN1BHecvEeH
xu5OrTKEtQKeGE0aD4PKdYdM1JAZqbB4jhUDngFVl601aOsMtl5WMQWQURHibdq8
g+vgs0YYL3ZHKuOrQfXNxON+lYejPaIgnhgKnLkrA0mmsLEi7yHX6QgJqM13+AMP
pHzaua8O1yTuLiLhCvaU9k96MlxgRtk2eRllDVsxarm+2+LWfwfukLstVI2HYk0g
k7o3ccOKcusU+E6XMxPij12YK3QdhPq5BNqz7f4No5F+w1q4jNaqGaAOKciM72sK
oNw5kRrT8mUJsCHPS2uCfZHwQFaygBhFgliAcnR7McNI7qAQmbM29vFRcKyqE9pv
qz3nSeC+Blu80m7EoCCPHslO4Bfjie0vht+6xj13De7aNdRL+tRSQ4iqWCHKwf7S
NSmYqybIXDlBSk6P/79ys0UpsO4jY32Fyxl8QcPzVdDWHwMw/MKE2gGOPXPzT4BL
x65AvUqYT6UqvSbRJNWnNaohRLyyRHP2gAH+Vl8nc84uI13tFvK3Paz0UsqMnN4v
PUcW6+tmvCWjG3C9VV+E1jsawlfWMVnzBejwLvStIDksdRcBMq7y4YWAoHg2jM4x
tjrlVVAeoSIV39hv9UyxT3lqimhC+eQlUbvkD17YPDRjt+/fNjPUdefQHf/sI6/E
78+6YlYaaU8Wm6Z9DzrKPaV4stNHDNGqOkTmQpY4KaYhrFEMffyVhBOHw9HxuzEH
0ZUw7TdE9vgeLlywnt6+YroCirWNZG1t5Fh4DyI/ndXcbMxr/HDoh+fCgZ5eiNPm
bAQ4fg201ppKwk6ahhLNQrh5gmqUE2ZQrw64SqUJ2V/Rrvm0BM/QiFos8582BZgm
xNuIzbW+W+eJ4PpnxkmmL7EqY5QZmJGr19I/Wkzs45JOlprOdmQU8EeP4QezYLSD
5LzOYyU2inwbMxCE7VwiG/b2/jm9i33nra/fNljHEl5fQKKTp716G6s7Fjxsd2J5
qY8oTj6HHhF3FIMwbxEpCWyvuRzEDiycxCjT4ak6ZDNqo1Tc6D+ljz+JYIPVghIA
UGFqudwmYFjYF9FGMgi3lsvsyfxy91layoTK6xYvTr4ZTo0xs7Lm42tLz+NRRF5e
Kg6XMPzJu6PqR3GBrdCBwaniXk9ubYXphFM2m619ZqDany/kAL66bgXpAdR4QGHT
NkHFAgzig9fLqxdi2IErCja7SHStVts3oUUwjSuPUDEuk1hSoC642XZqytMFhnu2
G5A09As1PPZlICYXZoiNqFu0pImyP0w3rMlx4G12r1OYGG5pju+eVecIAqa6O+2p
ocnTUuvKQ3DcBGkwClvhrE5pdxAOwgPte5Htfnx+zutH0hqFCmdUlJ2JyTR+muhN
LQHQXplzK36CoWxbMLhe4TF7o64RRqpoRIc37peIyL7rxUJyBM8KoXcbOgz7YGtZ
x39vKz4YbMjIkn8lZ2GicmZYS3D23msbkMPpeoHRXwlpmwLcCVsnNGp8/eSgCLzZ
x/8vxUHrItWZBfSalHIaZ5rMXiIJaLJ05qMolb3M54O8Z7rXpGCyeoUm51D1paCm
NJuC46g+Fz9mLYTfiMvhavOtZvjSdcJxJxj4krctPszLN1oEc2aBDE92hVVNfrBO
cMB0nCAM7U27kkk+SwlRVKNDTjNK/6TcEFKGx/qAwFi4/VAwKOtIHVvQrJG75Far
ddgjLPDzuYjDoUPlQB3t/ozjeG8FTzcRkhx8SRKCRSmBPqt6f2h4C040dVhE46ZH
JXEjMfO4kDlsS9TzxhkGeU5I2dgb13v3BjXhd4bVt2Rf2DjfcChslT6MHef9IE1o
mGUeHNecvvCj8skcHOhlPN7Sw6PWomHXAbUYGsMqtoGy14ubBX0YIawKLRcu8N0H
M+TH+KIHcMKesQAknWZI0tSqpqxqnnic4qrADWv1Mh4DMpqMand3oe7Xp3p9mEfX
EyxKwoHCdOlRsH9plgLdkqGHD5IaCqQXzmN5DyR2q932VauyOjouUQi6tahjjhYZ
HYikcioPtHDqL0XA9ZN1Bin/9HeKp/BNMhshZUFM5ryYGly5SJgT0OCL2mrrjzDl
5b9uuFaPnCgsvaMiIjEp0RKfCBA5PwN5QrLnzlaCrLlfYZbJhmGrr8W+f8rks7gx
MH90NqMgnHyScQCqz8SyMlkn1+khDb4mab6dU8uY2b4gm5x8cUwZqWdgrpwM/3UF
Sf2lgAnFoLfFH5GzUBLeOmZoF0BjJ7ZAF58XK5yi/CqaNDvayXsqe5J20YNGgsWU
W/uJFwlOqSLWTpQBINuxW5a/NzeP5lO7/BdnvbmKVhOAghAklDHO/eYR8DRkNvdX
RV+T34gw8gWg3U6z+Xn/JXeG3aT5a3E9QGdwvN7aptcUQsY2X57emDzABppcMJB/
3LSChkpIm0TWQXfal/L6qqTfdwbRYCb2WptPiOb3FNiyIfWm+eZtVkI+O1ykAF9Q
vcrBkNDiZ/RaVnZSkEghxl/CDhpHVFqUbyYtsCbjqshj1YsKbS/CTc7KGMdOqQaz
9rDhfnp68QlgktV0ufLrbSgEPpObBjvhUgB2uejZzAdzPnpyTKwWtUrLUCJptULa
ScGr41pMjGCh47zfP9qvWepyVf718gikO11NAA0r0fbtipc2UARfupt4Y4dqfKzv
mG5mz1mNrpocBLNfl4YRqF+N3w9QUaqdYqvhTb7q+2xno1zdL4DTjJngr6T9n/kA
4kMe5lulyAtgT0EFh745hMYTPCSjgWDi34nuKrMC1FNJgH/JyvYRyCpXqlsXFvDQ
BsZQo2sQ6hbXwxTI1n8bpWfUqkddfsVHJZiYbtHh+3QRYwF/xdoWbaJwZv78YcoD
Xf6W5oCNimtWB0eKZP7VBOmLsuEfB1ZQr85vkNCOsvtYWXsgK+2Yo25eRHxZLGX0
u1ZTq0Au5QbGKBkhQF51qBTEm6rWf9zhEyhM80REmBRkMpM87F85GD++uEZOZuTG
1+ajgBgZLEtXSk/5G6DOzifuxpcawY7xFLC/FhreyO9MgPJ2WhHZGo3Ke2XVoP7a
vRyOpu+rP228XhADTyeYNx2PvY230BQLL9ppoi+sERti3RZIz7/NFQ+QwS9Q+mdz
x/ygQsJnd9FrZXojM1XR0pzb1UviL0QpDt4U9ZOES1wLH7sD7kWLdg25pNm1kl6T
PLFaxMohCihDIo8NQcE8BCkyD0l6x5o66qNJQXUxFsbmitsQbUhrxanfQz/1ZRZt
lEFlC1a5upF2dcATXojkJwiYOhxYQt5ypmk845hrTzoj7lB3qFbVmHBUrYgzYr0i
RngiPH+rJhBuDk5ehKP12ZDyJ5vuEPo4HlFYltHF8l+4L07ZWdidfz/Otx98ZxAT
VHTQ1ZAomTsJbmfRUTr4xlxYuK6l8a1jzQo5vQGn5PiJnzEanSMg/jmSugJBtZa0
0PFiG12jMl/hUpiCkvyoj1IHeCtP747hPS9yZbxi7Mocvh0XVGWpIdOUvoxmqePT
knjQETK4pOg8557T+zeEejgDbAAd3cr8OzdOY1PSvESwWV/kzKxyHj14FHuidCM5
dmb3Y2DUML4W09aboNOZwSX0p0UgeRYUWGDBPAJQE1drH7ZT50L3LO1Uh/WXxN8f
FNh2Q2gWHM+iN0NASeksbJ5ztJKcXwS67t60k3ZDi74qzhedmXwGmZZa0hxmYgiv
ZdJRAQwRcoAWkFiGX3zgNFG+1C/lEpGhdYsavskIH4UEsaVpf0fE0/P+HRr/91mH
09mK5ggOqZuR0Pvf0yEAQN8jDGFRzScINGYuU2LkSdeoRDtWGxMH/d63Ew7JpeG7
dvHK6YMiBKio9N9zJxt717WEborQKAYOApfHWPta3CI3CxXxL67aRSdyvCacv9KH
Iz6PwOEnXC9lz0WlbwUhxxV+gqt2c4DdGakR65bmrdzIFMYWsfHjDnsEV13aNr1B
ysXopcHQrFr9UoSSQWcD/6EorNTN9sdv2nmy6aayeG9InkjYJhdUfWrPcI3nQkBT
smE6lVyBXSpk5KfKoGwK7Gkp7s6jbTJN3BHD5S9JaS6NXSoKRHdHRlG1Hz+cNZN8
W/AbFjGvMiqpwZ0h/VgCZ0Fgc3iGKTaJ4KhoILUpYRiDlob6lp6dxrYkJGX0PKm/
cLQSJpHiinK/GUhhCxEd9kPd1WY3W43Ld6yexbZloqRtrbUGHDQfHYnxJtzpdKwU
usrQbtOiNRZ8TzvIIE5dKJ+tyZZQ7VBj13e1XDeGTSmlDP5Cd9wbmhMm9f5rB/6i
hyEmogJVPFsQQdPZ4SXbhn/bZR37UmYIp7Wt7cmr0G/0YvleFEarKCvX//dYkg7Z
LTu4v9OEhvRTxhjkPUmamLY4UU8MQHeplT+RoQk3sGJlyiKqEHoxShcG8bdUhqoT
qAlL6IshJv+BWyeEAAGXy5Yf8Z0/cNm3cKORdXrExxlvrufuvbBnshEEes4Id1oz
G1Cltj8KabBURTFf+kGe/7uFlh0qWDD93CodUYDeQuo7dPNcHWAyQxZGbo+28Hqe
A689djT5MCPu53qPkpwL8hMIvg31YoYbEj14rCKPYMLQXCrzo/WWyCrccr8HAPeR
kYAw3ztsixVq5f19+UkvuroaBGYchKw1Z+AYEunaNYbgnuadUDpNREwpd+Z7CuIh
HDD1NmoRT2RHRvIYslcvbDnJCWop9oGnsykMYf8J7XREMiI4GsTuMgJ3YfAEV2PI
tDi2Hztg5m9IECtzhYT7lMtWKhgHS9+VvMmknVBrPuEwydNeq6ViYqZp2J1rfpgm
FjDcDoBQFyVGacer9DLmb3OKhFoKonoLODFGQqlHSc5OFimgr87JbGHEfnVlM7Wh
d3Cg4pSl7/CU8IbVU4CC3SP/tsIjNVzw5Ezxx1h31O5fuHAYLbeDIqDlkullCUqI
8WmOXa30P+V+Bbd3rBEye1zyysix+jQbFgvjL2izUW9BXQxmvZPSeMy75/nK+qJC
5B2XsawgN7/+81b9lTWRYvhAOjNpv/V758I8NSa+mzXOW/PWTZdxaJJZb25L3wAi
kSwtjxjXMRKwxo4eE4vThAvhTuK4DRWJqozN25gEJ0mDLawoHLqwPU9r3HZGuzYi
a/5lAIZHXwrCBGJRpTwwSH2ZPk94RDJaCcYP5G3zia5riBDrH6cCgPpNRplWVe7j
/GMLehAIP1Qo15iRDtz+3bWIAckBDrnSURqVO3FVIK/tEte4uXr9KpbPkwyyaLyw
0BhNGzwo1ZOklfHBeK/eOGEheWh8Bt6w40LzBmY5aEhqx/owBayfGjoeWRf1cRmZ
HY6Gi40PgjtNUgi/VwwbLGg6O4VSqoBMT40wlJh1fTVrNCvJIIRhHx1IUVJ5sl70
xXnlSN1rGSbhb2hFEwIN7CzZgJv9E8HLPPCV9XBjwNrxgenDsmGnlQSRApT0buy/
jgfb+PNXbGBp9D5WmwA1h/LQrBJhpvbtd7VytI9DSwQ2usA4M98/nvZI55qdWG+P
kejJrC+8E4kiQpnxJdkNhbf3ipkIe2ucWHIfcOpdlR9alG69dc9jcTtrEKkJmLYH
wWfpdnaUTsYLATfG8jrdyCQrWY5grRRlVbZbdIz6Afu/p/cbVGSdcNZmSeILDXEQ
cOgwDxLRNVCiGiZVDNyNqzHylqUirqipSge8a5DwlBA/l6WabrLQybFY77ihynCI
iCA0VT2tI7xxI8sRHU6uYD20Ivw/p5Vu5KwvaZob6Nk+t0BrPYfdepJ9jeAUL5nX
JiSB1uk4nXswxQ0nDhxXyjzm2AaWireudhdD+50hh2LHAbjfvuo3DZnvffIMgE6Q
lzRXVzNNt0GId2HyjBCAX7teVFwP4PdgBvYBAxJ2+mtFcC3Lo6rPrHjm8hzf6BSQ
addECdcVTFMAxh8NcluGvx5T9I/oraYPG0HY1sSI1QN7mXRoeoTX39Bgu2WIILXo
pth53R9n4nxrX6cACIQD3+yd9LKhvdoS6Jd8Hpgs98NKS7o2QoG8xX2jMmHTVo8f
eHA85UvDGy4rsJULSIFAti9n1VMY+e/tb6dB4rb2mWjAWETsT4tHtZcQzbHhoOUd
Vu6xnjR95lOuVkUTjgpVBxBOL/4rQ5gGeJ/JteeRy+dqLpsnfRxoP0PYfsLNCRYS
UL2RdegZUCeQ9Fbm5aPZmnNLEywYxRQbdwuXbJTfWiQ2l5fS6uPEC1FgfwKvOlbD
08YyVEY5H0OLMG8Uq4egqtAvszzfHGpoT/KjAOH9Iw+W1cUWzv8Q7ZxvQZeKeRUV
InPQhu4IoYVeSNsPNdRAtUuKkcsG6NXduK2GdTS+jdsAy6TRfLdwdBpHjhSFntHi
IaSzZhJ5J8XDE1e1ef6DWKTbVEAtPsG/QTJUQvj0lr/0qwggDBNWLD3llz+9KMtb
Zn3A8w25vAzABG1JCbHJrxfqojTORDyZ0HZ761nUzCkhCrZDupHkApkDaChmeGqd
48cJSdxmGjLPxz8HUjil4SQMbmYoRmoG3XBCal/p8tdCPv5AbUk3IgxTUypW5EQM
XOZVYn1yy9RvQjF39z6HVNSNSZwiLXxSvherKhkMTyHifhQpRHp2GWgCXz5WQxos
AFQZFxI/5wDMOGsamhnimNSz9W67Ku1Ive5nr/xIWGtUOshy0wg0JcMQtKFrKiJI
XY5PgQVjJBFuQxmbSiYcH1U37Cv3ooWtOnykRj7vmd2Y0p/HUM9ewIh9C86J0wZf
X40OrnFIxvEEkukKtTkIHaQplSa0JbdP+G8+e0dAODuNiM933vzoG2MPEAlJWFBH
MCAagdtk61v0GA/g/5tXRP3F1mCgSCJreghXzUGEgBM/4/fv3CJ1JJdQTtK6j7a2
h3QodywR1diVxmN9EUFp3Bs975NXOhXdB4/cNm4JNekbF+afhephDWUVauMba5FY
3YTVSZJ/ukpSUIwd7ZY8pdkNgxdhYhEq+GpAyT8UFSpuLmnkurRNri2CQY/h0kVV
MvvDvZj/EbzzCI3EKYna5+ggg+r1+318l3a+B6sKnLS4fnqGzAYDJHZPNp2Xn67b
oomrS+p7N1xx66LHXH95Xj+k7EQSiSrFTENdafJlYM/XVt5o4IeYFCypbpBzXDWF
b+up6BYY6CbhMaGmPVsRx5ealRPV+BXfB31J9rOl+WONswY6Vol11ZuMysZzgK+i
yuJ6xYGSq0iIwwo6w0X5CAQY1Zt+bNOTkrbwFA5dDzwYME7TOXAZv49OF9Bsz9Qq
IYl/0pkcTJTkG4JX0mcmHhOMY/jCJC/uJqwPJET8L4pxINIen7ScSNwisW4Cahsq
HcE8VyfxuZiDBuEyELAeDZF1z2IJ0M6pkXfgjAqK8pm8lkk6l6P3zxcG0A/nQ6jY
otsbvE8om7J86xHWkDcRa0Qpqovbk0nSO0m8R64gyl6UV80f5V7mUJEYoN/QKDPr
AeSwwH44Ve2QPmC9304OYixzOWJfGTBAeYf1U75Dk+ea2L95HqYipU5iUzAfWh4o
pJ9ILgRRQJb9N7sbgPzmujcLNEGF114+aLA8/WRfekLBccgak3vssjO7wNQwPDwj
sUSvgzUeRJWwz2GjIUU/+8dCDqulTjPTe7dX41aKerXND+wsfp0yuj3ve+bG2Q+8
N4TSOqLy3kiczUlUD1OfdJ6gltqZW1xo5pZSSeUdJHX5zphjmO269tZXMRIi8W0X
FKQtEOozbGnd7qinp1+2DiSCul75UZFC5YgChBeQrC2v1BJkqGmqfXf9bp10IrHp
6Gt2ngf7PFNks/KdICTLYGMEVjpaxBF2MmDi+NiQxRQIBWK4le4EzkwyDucTAyM4
HifraRKVZm5b1VbK4fD7vhvBn+8hK3sPviTT6PSYCdye/Bfu0H2b48+S0j0xm58R
QMGogzNxGAvUaDZMQdOyHyqhabSoAC3ypXtBXdSTeD8gUVHUD+2E3kdHz+2U8U6R
VaZBmr2n5P3/0+mW6LaUqerllD8uyXf5+6WJZuKOe5D9/vjd5ujQfAWxNcXpT9+t
RSUC1T6rfrqw7fWPqVhA9HWSMQNFKQ2ulK0xeKuphD+6mr8fW0/zna87vN7plNw/
KG6Q/IWyOcbSJkq0azY91XVKLkF2n4zFE+7naEV/rLfza24/ZBusFylqKLcNNpus
HxaRw6xwWBs4ADN6zSmTk4XM0+89TFCTPbLb1MTCixukUPHmEc+AGJg5NtjVvlPq
J1ThgjzAwRJuJcxX+ZanzhNbquG1AIitny0zjEsau33l+PInusbo86jNIibZ0TN4
SOz74vHQhTieNRvkWpv4DuyR1qnW808kS+UnHgghiUMi3HrpyA4dgEymRGrR+CwW
g8mbkRsHuYpRQSjlGlcD5yUin3VSz0u+/U9hNSyLfalKLEJ2I75GqoRCeQZzvPoq
slEr4ZT4Is5MQZb0U26nrGr8yPfwZxlrijUic205QmraBPb5p0MKYjTBt+QRbrEF
2waOeA2zGl7KiPp2lQ6x3ziCk84sIgOOljmMNdxU1sl7dChnuNcYf0bm5BxazuX9
ADHCB/7MYEcH1Dw01sU1oahbWr7+3/vSYU5Vq59wCDkxpQLZKfnNeAEiWIUFUbCn
yuKQ8U5i1ez2xWC+Wsnvye9dzYy3H7NerfLqYjUv99P4p6txLhztm1w424BmGFKZ
iQ8nIZcbk0Ba3HWtADkZNQ==
`protect END_PROTECTED
