`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85KLbUhd49iXS7TKASJby24SlO0bsChOrRNG1iKm4V5Gl0BcnmML2PsgHrd3uBWF
Zh21t0jNntZajt6uuWzjBUnE3oPC6rnlcZ/uwVgGmRTiR9rrYyE1dsRYpHtRe+zz
Kx0kXgt04eVWJXZsGqRJ9kNxz8v6k7EVDYpvo2136oD2I41f96n8SwVdLngVKbUz
W7f0AzJuZ8chwuYpIlE0fGk1JBkCFmCkMkFaagCXHQ4EmkDPyB67M4I4GV/2GIqT
ELkukQ5Ed1KFL/UhZa6Xp05cItef9a/Qayl1HK8TA/lgXDle+8sQltKq0ME60a87
LTWHrD5otibbJyqIlf720P8Uc94Pq+Tebu8C6VkYG8ggkJf4pskBxvyxCfKF29gI
NXovOs9A7+7dJDCCQkIcPtyPRRiLMgk8GhMZwniQIqbdK0cGl74RzjXYZOd3HKTK
RuV50HXSZrFFInH5tGXE0Cqdu+uqA9O+tjxkV8X1xoiC3ysSYCSR4Z94i76yiusA
`protect END_PROTECTED
