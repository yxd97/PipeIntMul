`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qhqEu97Ucc8xziKmMNfiwgad3j5Lq21LPYh6dqo+PlJ3nkaRxkSc7D93SKBXy8gA
Ydgi1cetcOuDAwjfZGkJBNhYREdjFP/za5x9A1FKfKA0AM4qDz9phejyVe7BnQev
KKqu3nez1aVIc41KskaVy+y193cUHu0rQqWxcyvvxzOzHWmxuuC6ah5DuLZYTqme
GfPUeGFWsNZcLg1rWDa6A4749mzgYaEuZPjBpuEa3z2hCgdP8Cm2UHLT6JygEwbn
u8ClaJmiItuPkjJUP2xQDvk5oz6mLN7aDYvMEHxUZ1PJ853ViLU/tBii7aHC6hjw
7ZAUXHJqe8BI9JyCNDS0W+vF0O1nqiB7i93NzSrVeNR9TrjyckwrlloDncOYgRVf
`protect END_PROTECTED
