`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/uL+vI6xbDbIajLTAqZ/OK9iPAZrsCOuxMDJ3dB8w1MVMJUi3o7JC8PISNvBGRKi
+wOff+cAyaCKBJjFo8DmPTKOCVib7p34ZM/5DYRyc+wU12zmtOv39kpt72Z/7rKj
2xTp3ok/n8zVx4yNS+4UguJGijzmQT/vLA0WGY2Xz4XaQanncYYvsHw9VC1/o2cz
xaqFtQutUpTf7sZYT7xFq8fwtwC5WXjl1Q4Pq5hagiy1glQlIWb0oaEx1thPD1Ss
niR2H+Dz5O+hAL0gLJf9SYEmmxD/cuRw31XTtQJYThTBICy6MwBnatPQ0Kzz9Zr+
iX6KWYlUbn2O7y4ycVqg6ig4SRqhDyTkCYKyW6EhK50Ii1Rdw9gsKo5PYNDR0Zam
`protect END_PROTECTED
