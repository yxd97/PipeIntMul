`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oDNXUowLf5vdrfe9gI1qdJVt2KzI75puxAqaWZhfHpb3neG0YICZwwuy6FY+VtIH
bulEFeaanaGgvKx3RBAGUJERIKpJI7aBFW4JOsP2HkyEisSfo+Yv8LM3YhraxvTc
kEAkbUnxq6948e/XN8mOFfcUPaAhJNQrDCuAe5g4mzvkNZpf/IorrTeoizPDMBZN
beff46xNLfG05hct6u6LTgs5SCUQClRsb3aM1/rOJ4BPI3N9bSJZmjWrxwbnP3wE
+qMwgnJmslqxLd/4N6dtJWzP2r46HfBNIO9AyShbbNsZu2Xl8v6wsFLhgnGj5YWM
4Sd4i5sh9dvfARmoO0c7X0vDC8xnwNmHfMz2EIxW2to9mO7G4Pnl27luNPgaNChl
CmaqglH/iRdbadYjHsIqeWCYWej7J/fGRhjq+UcUaw/a+kmoyfa0zTO7M0TkgKIm
EAdG7fmDfhNOWxJ8hNREHUm7xDKgS2VNZyy3f2e/vU8UFT0Q30wp1SPjBD3KQYop
5qbmEFPQjBIxQe/C31YBQr6LucHZSygsPDtWKFuCB4B4vngalSCzeHQAEPN2cWJM
ScqrAQjvYt+I40Bf3qPiADCLqNpUtKAIMo8+AXcUHEwyIlNLcsj8jYun8b67Msrx
DZiQjwINi/fnnW+HuSL7cvfeCFqAmZqLqk7EYlbG0X50uGUad42EmKkFcbnvSFnB
1W7vv9fyRPRJZ6SWj9cGR9J6vtnqchNeV9ehACS81ln8Qr9btBTjjuAcnsitmkY5
OZLGRovKNGepOSHtIiIA/4TZ7nuBjqKeaClJ0x0P1fiDvugZw7Bucg2JlsS/+1c4
CHSWEZkMZmtn5pQRSbV5z0ePrPkGs7D3Ib5xnSIAE5gc55lPJJjPzmWOs38wLmBn
y51sEj2MOkOJiPeEvJ4m4jeCJ0CYFoUW9wfk+CAB8iuJ8ozp5fXGVaInh2qJuh70
ctITYbe69W9rqi1Qs/QYHcEiFBFL7/2DbKoRZuXcWBJBmdvXXABEWb4sqPI4pAb4
`protect END_PROTECTED
