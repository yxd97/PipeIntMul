`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
evGxQ1Y3cdaac8PtODhIqH/4SM+1jPItYSiTdrWq6KIYbgfdwbLsVSvUq+zR8U4d
z3CA9QRrLSUGby+3ZQz5GQODvkw/Ha/3nl7/1gy+kjV2v/+mxes+r6NGHn/4lSJB
MtYb8GABJ5JOAEdXcqHagDyFkzqI7ZBAK5fc+SdDzE9G9SyGTGtLXU9CdkcPPpXR
2nQvmTPt+rgWo9XKjFa6MQlOzjVDBlR6B4nuILO8Q9GgP3tCRJaK8amMdvkI4GrH
qYeyU0p3rdP1/ZFJ9iLRHHTMX8A/y+ZRtaDd4iGyM6Viw7/r/OE9F14YsvVDzaJ0
4776xx5CqzLQVMpSOa1bbnmyTZPF0PCM/Dkk2LE00zGfx7ygzlUtRJTj20bruZUb
XLN8FwALfJZ/AbFfUllF2jf1DFxIe6WYt6+kMXpYVc4=
`protect END_PROTECTED
