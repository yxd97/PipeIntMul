`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Oze/8kURa7CUEJR+6LCssP6gJ56PwgMa0If6KzuDwAbghG6vhGDJ3BX9XDpucEiE
EOL8wrZU9fomBOPs6pVFh802+mpZQ3sKdkP4+ROpw/kdKQ+Ga4tV4nI+v5s767if
bFcoMLqoLB+SUkyLxnolU8L1HH5M5aCKUNur/0Gtwz9SabGsggFzyktE0HPP4x81
jwl4MzMfWnNKVg7H9/tEDKRWtkjEVGjwOSDT6zyNPnuNJ+ozRqSFoSb5Ud8KEgs+
K/Wc5OOxqS0TfeZhk9Je99B4tVrlqaPn3Svb6HZ+m0WiWd2RKZsyd4NgdruCrzOU
ADaMZKDsrJc7MSxZ4msTmnBpBQGAXJM7Zd3+Zjx8tf4QawLYPCPxE03KJiStATYQ
gTcUEYQhTO/X3n1Vgqytmf6K50qREPCUwgJ3Xi9jyQUBVIVSQUw7D/bk4Q/5OdBW
XIEElskce4AQajKWJ4h+UF5giT78S67hA0ljo+8JNlDxxTwtzz3y8eU9uw4knVs1
Px48LHcNQsGUtle75nJmAqro0V0CHczpohAEJXajnc5U+Hi6utHLPN1VYFwDVonn
iF5dDv8XFfqDiE1wvo+O4nz0DTkNb4VGhodps3N7GBjylr4yOjg785k5izDU8iH9
z1htux1NSIdciVRVYNScGTP5hPAjZP+yorGj+ekO8Hm1/Ie8d7kxlkWq3NGRInhC
r1vXmMEaDL9H1wug4E7FPRRO2kEExYsLDDLjFbsbPmloIOv8hY7Rp8cKAelhUDeQ
e5i7GS7zW8eNl82E3Bex9aJNLY5fRzg7C4WxWStkhNw2T7UjRKVEXphgOIYqkOEP
yln3ZHZirrFFrCEw1Zgiv5WugKGL8Pp9KMJhkjdd+e6LUQOu0zm9j2NHfe4hHdyG
1iWGF5k//ZpIE3GE8dLETl26mHaBfpDJJQFQBrEb90Vkod1rj7EZcA5H5wj1Zi85
`protect END_PROTECTED
