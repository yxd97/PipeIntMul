`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PIVLi6AjAFAkHnhF+/wjPsPMImHglAugNj9ZTK86O0GSmWaBbmPwlKTURzTI37Ux
f3QlSkzh3f7MJf8mVTRrlzDPfEJDNV9CFXcRU+Ex09QDdmn+xvRNy8ZeygHzGBLb
Xspr5Ho+IofqxXy1C20GlTnrnOCHGJf32j75CuBCAqHOK7ap+9PUM4rjZ7yWR9C3
w9jug0r8AVsEqkkXGR5Seg==
`protect END_PROTECTED
