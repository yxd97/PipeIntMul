`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGxhJoyCz08qdhUIiVod4A3mgnyTF72mnC+beTw8L8ksjhooYJNMhXT9TW4XT9Yz
QCWxeMsHUTzzKTOW8zMQ1HeSZ55+YJP49BfDQW0XdfhKlDOpQc1I8f5lca/U3cS8
FmoSolYXWp4bn9u8gRooAlfIsqo0erY8rIipwCnlU/MBxeQ1Yt49v4/Uz306L22V
BHort0OHr/1S9e5hlWZOk0MuiUB6kZwNRaKMhy1Zmbw5Om7zoM1vh4+18bs05eki
4wO7tiKSUUnB0tacY1wdbfWoWQIVv4ydPMPhU7hHaq5F34WpLRYvrfB7dgYey6Lg
nObrgfuiFHjNIr1Yeg4UQkjwA0UFgIbe4Yu54AscVpUZ45RnyrWGCWjcQvdG1yf1
vGKNLnRNX3jy/a1HMrGIZA==
`protect END_PROTECTED
