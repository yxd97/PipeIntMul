`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JrDvRv7CB9DbL15zmwhx9DFomaqOhfzWzjD4odIC1olSWPS528g9gSffR5Vg7cwG
LUawkif6iWSSRAjjLqp4BMCdShaCiYEB2Gyl8mPCLabp9pnB7taTvQB5f7HYiHdn
8G10u0Lex+k/zptYXe0tZQ2cnrgfBgx9duhAicyQT4Z3QKtnsPUt3ZYJmNhQxHS9
W6GlYFjH9C8vTdq0IORwRhQLcJ2VS1AkjZtqY3M/qA6JCwdGMLKgyF/A5zou45mf
rLSJ/g/IJvRH/r8lpon8F3WcIfsj5vMf2M7L3MG2VN+x1kfIOf877Sa022crqR64
j4A5XL0gXTmE2aK9BZ9EC9OA6073Jw2q3aCG6oETn4A=
`protect END_PROTECTED
