`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GGK6xsuy7+wB0w8+TVn4efgTJkmHVseRNdEH9bUazGnV2zdV+OJbKVhp+uJ3PpFx
lrSO2JaTO0mQ8+3Yot6AgUXLFgpEG4BRbgJ5nBMVjZXc6YWd6Ikih7UrPQjIc7be
hYnoZV9jX5Y+ujmbcvD4XYnOl4lJW/O8B3XC55NYuvxEJydu5TZnb4GiMd8zWJhr
tDgJdQMVC+aen3WeAQBDfnn1QKMucXa4gGL7WvapaGtgdWUNHmW6W/Rfq+Mxq+l3
tSBXNDY+0sj30+f+N7rJWCdaZwmQUXctAiYr1Nw3z6MORStsf70TqQ161p6u8ssB
B8kHxk0mbTo7U+CHm/VvUjs/OML1s+GJt/KP0ti5IK48Q3nVm9rEw6JaxuzD4Qoc
s35r6ar1H7NMQwZq8bMnKj14PR4VHmlg7Ju7oy3d9bP1S96lWv65rPz14ZPSvLxi
9ciTnWcV+rwE9FRhAe9eymMbA9I5wsVpu4aIkShBhhid8rIsUM59Q79bwppRaYNY
xNGzcqFc6UkyLD7H5u+3JB8FVIh/Pri9SwbWqOsWXrXuxk3UrP5zwhp7lF4aveaS
Vz8cD+MMrsdmIaa0yG3oyQh8WUSpt9kq23X9jU+s83X5Dl/TXcIcxmEwZnbFcnBt
AfAIcLnONEydoQHPBPNMhg==
`protect END_PROTECTED
