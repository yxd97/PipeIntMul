`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJz+jr5bYnDzPH+oCXUmyjNsz6xAAGqknpPCw6xWqs5+JsnVh1x1J7uYp4QIBGO/
lvwd3+6qs8xcE9VQlGhkCYDAw80YSd8ch/pdF/+vo7RojGcBI26LybnzVArMdu8x
6eCr0/qoYPSrEqfP+9zRuHNzL743SlnQjiQ4LMzxn6XFvBCX6mKPRF6834gSexZD
vTi8nkSjhGyUCVGUCs+94T1TE9ef69zkmjDxdfFouMUOM+FvnKujDHLDJFr9gOAR
/UMcQPnADV07FL/w0ZaKTjBpXvRjrQeGOJ3W3cMHgXHhcCrmWr3aoiQv0hkp7Rny
cQyF/xHaU03AOLnUHu8E+90/y22l5/RG1ZP4UyBSn4JCxKRxV1IOxnf0p6lr/2Jo
fJtPi05LQzCoATesIf4ie3cGl1WaWMLlzyH3oajmOxVUsIzmPEj9kmYuqpHNxa7r
TckOeHBGwQzGRwRIm2AGcFq7dyL8loPso+CuYRQ2VpZc/8Qxf3+5OBAO7Iw634Tq
GKEiJS1ysFWjb4Bpe8CNBmW9uoidQ2l/uqaAr1MkK9JePVkZMqU2UC0R9XO3VI6u
/hXjv1jqxs4ehJw4r7aA5YlMOSDB1lK4wHIR7J70jwU4YPtVsiAUKRodw/wOZTgV
lz+JIBcdoWSwyvXTk2/YMT7Hfg7PAgoXpZML//11FT6SegtPZ9LpzvjtBWS9skNa
M3PyvoXdTZxzwU/VHYPd1FCjb0U56MSKKh1HmA07CzS3eXdkKrXd4Hop63xiT8nV
V2Vrhf/TjOnLgn3gqMR4ABUG/zswJoJRlmmBWAvdJlY9l3J0Wh8zN6ViYTgELupT
0/07GYAQICVrzKxzCU3dvDLkBBUbHP3FNlVnbKlFLW0cFAfLnVIeD51GKwIJFmie
P2PlnwSI5NwBxIWt9RYBoHEHyQuAEfgcSxRIu0Do6JnUKErOEBhRBsKeXl1BSI7C
VKRBtCaDwwaLibq/mu1B3cqI9/XQYeiKAvtxsCDu8wZttKQYWdTpIapKplf9zKmT
1oerhGOV9ztj2laYIR3oeXAQ+Md4Rghj4fvDK4JEqaHwwVSdj/55/oAELHpWBA4/
Rpw8JEhE9MEWGw6uQRVrhucrmKFsKOXBvHDmUaCYK7tbnphEWf0IxSTjhfJ1ZWtR
wG1C1hU+MxXSSl083MIri695oNma2gJFvRyiUmW8mXf7HzGKzVfMBqxYgs/jX6pC
`protect END_PROTECTED
