`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbJw5xMm73ipdBZVh2oipzoReafdlhYzhl4HG6LL1flASuriBD/VShnF3/WK18XX
4yJqBk5QvNNlLzVVNZ3gXLEo/2mv8bVoQJiJk4fv6kvoYa0Z1bxXfSWrnICbLK0E
rJwOsS/g5qXuFG7w555h5fkD2sQjG6NFrvRJysYEH4NvZI7cd+msOCCiANStcVj0
DwmuLqM3yheYALYEF+z1An8KOiKjI2WN1BSkt6GEeDpTcHZwaqMooU52cfryjCkr
o3CA3nQ6S+G4t+lRhxfLfk60CAextdPftnW85R5CGKyI+2nV7BjtKj0Ns2nDnLbA
6WbmoP72RCvOIapayVCRumsckXvKqGXPPvaALG8aRhIPQBIGw0Rxb1ktsbeb3vY9
J1Ba26P21uRG3BADEIspWC6vSP+I1zOein0c/Ny5jvzfBSvCA8XMXryMqvAkFk7b
AZH2Z/NPgZAcFfmaQjod5ZeplE1n18/SZ4uFSHb/lLxYyHSIiMqE+FT9DmEtku5j
u1WseOYGhYE1NADsib+MqySCl6KYFYdqKOYS/v8NADaWDNDDTh1QQXC0t5cCX/p8
hiaeNm1O7gC5ogImucrFjSOhIr44reCqD3TG5Iu6ykMbrPja9nTYT5KRQp3nWsuE
UMUNBgVSbhVjjFWCcEDPXdhC2taxWUpjLVpKftgrOkL/7WF1l1O/4VJoLv8WAZol
biZZ8xOcQdw+1/rhx1opzG5IymPAeFrHhEMXM80nFlD+I9L14SO7INQOxsE8GKL+
X7AH6sx7+u0hcpNCAe7Gco4KVCmA1xU7BPAD8eu25YsMvqaDm5Z5+/Sjf77WflT6
XGrYrLVHYqiK3UVWXIdzUxH8vD/+6xOCrpJqENyc1a58SdBY2mvckYiwIIZ8GsCw
Xel/xm/gp9eA5zh0Z24rMHbDL5ZA5fg/sSlz8UKuJzr4GoAnEWKKanvSpfQTIVam
I3XTBdtaAzowPAB2T41mquIkfbjBxw3sNDPu8sD8Vr33lMpEabg0Nc5eov0Hou82
I5lzj9ln8HCnHijtwMiAh7yyP1asTwPy6Ufnbh+QwKk/RqcpdCVxMsgEE3MkUM8h
yQ/aQwWE1hkp45YpOL0qKnUHhHL6Y3LnHpay6cNh0mvu3ok0/qM2rfJw8uxhx2c5
avPMHhJ79Ll6qB3IdvjsWokEjOjsrrnk0CvqZcsPJaS1MSawv/FrDUChqVVzkVaZ
X0tQULnYifdoaviDN7evXXA94gvCy5sZoWeVfnQPLFerHbYvWXmp1kesiAJCOr06
+i6XHrO5RRLTaS3YBUY1hmPsfyIgKZr5sX1/sHglruDLT+c0AI7wmCYu/X/eV+FK
2jmm6bdLHimOxTvp69l6ASvaaOuHlVcrsJOx74Ii0EPOpBG5PG3hZo257T1Cz64J
LyIO6ntwKpjFog3a/7x4NNCAsif+4pyE0JXz5d1AbgqUqsOh5sXiTobH8rfAsBx8
Y5qDmiwXQm1sgXMC6mva+RfhkeipfYHYNJm+2ARNIHA1RoOXUtoxdKkEJYxo3QF+
1NbaoNeRWYMSxy6UDSwX8fiZ9imPxyCK1DHqjIXjT6dmptQ3lMCJo++WRe4cphcF
87vxUtFJBcTIlXOpBb1GCYu4jusSQAAvyBi5E78hurl/wx3kXiw3bMs206dxe8cx
buEQ2tMUTc+OLub8Sov9zU1dEpQZNk9O3ExGrjs+VsAzyYJQOF/jNBb7kNX9efaE
/C+coYyt1Sqrghb5j57NrPPI51F/U/rwTRcxWGvtbq5pIsKf+bJGJ2Ki8n0RN4Up
jW97ozxdKusW27bcqXc9Jv6fD8bR+Oa31sgNsJ1omfYOLA8Jsiuj0RBrVrVMGJBU
maeN8OOZ2ZRNSlB4S4QPVUGIasnbgJ8pPa6UaVcdk0QPHE5nNDmJeqikHXqUWUa8
IgPuss/e/MiYszYJ8QoKQfqFkrcJvXTvYITXynqP8cRhtoUmjfYxisPDIu2oYdUs
fpGJb+mcGwoqQ29YfNIxaqaBbKjU1JdGY4l3AVc/8ZyBQRyv7fDI4McgJsAcbpRq
Jn6thvsOQoYGsu9AHueOgsfEFZEb3JFg9aNQ4GelIpk2WgxGrQyaJIDt1+ETGx3w
oVWc90ZtIr77uUxi0vXrVRGps3rb4mzBFkhhOmjcL9VcWZjgSVWKz590hbycET74
QPgMaNvoJ68jSFvKCyJqNyC4UoOFPWf01mo0DbtY6Buj7nyFhEoghyybqI4qfWpB
0Ez1yGvM8nM3Hyvr1Nv1eOtGDex1aoEIwooFXVVnfSlnYd9miAkDdsCPDA+5h7eb
wVElPvppUYFDGKL59NiQx1QWqIES6SqC9ketpmnwAdPciJmHg0+uc2zoBCRTasJd
EMymL3xSUsYZVrV9b28dpUUesw5HSVtUBa80cNHjtGGrZgbFg55w9uZAohX2kpK5
yX+XQwq/cJn4vRjNPbT4ZV9ud/By2fRI+j0K2CwGcnGZFqc+7chuq3ez+AAbMfnc
6gwAQfalOpti/1PcWNMhHhTFayfzYcvys9uLWle7aZ9qORabemP0XS8qowMGtwAQ
s9DyUUyGvSVeJ0Ib3aE0osT5DovGQszGqobJnkr46y8zXvIFtb4kYvlOsTZU4+bA
gLVsC63D4adJUICHRQ5PXAW+OahPlUQ3IcdhKbiMA2gE5WdY4g73aNp35THWsXxM
Pe8tFIKY9bOq4FhFdeYbvoEo1Fv9S6H0oRIOw5/VksPtyAdemXm1Q02g3syiCTux
bsigm//ro5NRZ3QzVWM4iZR8ZpzZixLoViTS0fvpNimEWUV519xeDMuTuKXhi2n5
+Z954MeNAaVqTC8SKKiElEdXMfRSsy/5OMU7z3xhXVXkZJyeXdDMMgDvJOJg6A8o
haDHEzzR3uk3SJYq6opRpvIqlmIjYo2o1MQfyqYD+zAOa/PaVuubb/CpQMFbLeTr
LjgmBFh+/mt9UABbM54mQg==
`protect END_PROTECTED
