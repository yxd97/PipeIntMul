`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J2a2A6GZYOflB7xiDVwM5iexh2+bzspFThKTMuQgsGrdtI8CZsmMJljmsryWy63i
rglCTDoUixDPj0q0SBkNBxfCvvkMS7dt0YXAiqiio9M+ewqnbh60taqmh3zFrw8H
1yRvou2ALnOuPayuN08Af/JoO0tbKzScKvijfiEJ5EpVyfueMzfBphpjZlAbfpM4
fT5rC3zlXRx9b//UhQG1d3aRbidobdKibFND1YB9YJnPt8hwbbyj+oXxHd1X4aM6
8cQB+H5CjOPBPHmiPDM2Tv474Pt+YFdA0X5zaidCfIM3h0phf+VGYJFDoNeKtUfM
B0ZICLAEKA+RYepX3qHUcYqgeZ4H/JffOmMLnzFW55IAxJBNhsAGuK4eRyNfuT1Y
giJqV/Ku3omXrpPolvpz4PKgvpZ5wYJ0aPTA/FydDJywWK/15qDa/RLa1o1bhjNm
trwU7fp+0IWwSwoHRxjAoMsaC7FCTrUrb4OrP3JmiZ92nB3UgQ2Wdl9uu4D+zKYr
B7sykZHkozYX6F6+/8RAgCgA5lWhjgfeaY0nr9ROLRPvekP5orYyb3Nqk4vqZJ5f
`protect END_PROTECTED
