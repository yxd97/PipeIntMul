`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
58/GZinYTSeDjCEtu2jv1dxsirAVVwN/OD88Tw45EKrOtyg953tUrv1yIq3b9GzR
sOSq9NOnKOnQSo4GJRsFf0lnzvZLCHnFCHjOK6TUEFNNm4I5VOJ7mCP5xuBfZnvq
HUP+Gfz0ZFUSx3Mcp+YBUCUu3JriIOgR5gfqocdKRpQY4WKGCik9jyhl0Z+rXMyx
+KnFzMdsMWIQ/fdd/GIGMum9MpJz4fSxMaT7wKmdYHDQAERafm60b/ZckFkm5NSx
SEOe/XGL8nT14XD7DqE/u2ALa9P6qVcHsB7b/lvZwe/DXnVRPBlchkMAKe1wVLs0
aJYgcfoBZ+4UIzV7MHITL2+Zhjs9fCCkYhtinQhlMn+/NHNa30CCg4z8of4LYHSF
1d5O+htfkfjVtUrOVFDGeXjN6QNqQ+aB34CrTFOEpSs=
`protect END_PROTECTED
