`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URPwIsiIUKexdayeIp8Vme0lEWwLop6hCVa+D3tCZ+QaAf/rdXE38+gW7yoQ50ZK
VLBwoR4WfeMgaqMAAgRoU8FTb//2xtnKHugnPvaePY+7twVUPueVhj6rh+N9NZbW
NM7GKhl+kyowCGYq/eOOqQhletjsau8uokImPeOqdYqYcYbXD8cCo+5XvNlz5aI0
lz8OkrZi1BacMgFRvAw/XM3hwSZ3mBJuKg5kcvEfevfueDkJSKUAWow8wJwa+abA
NrX0Zs1W5tC3TgADFfdpFqG1+3R5YQGFVjqUV4iPbDh45SY3CU4HJGtKQPO3Aspv
9UxeWesXsUzNGK2PmzRAF+EhqngfK2rs6oWS6ltFgMBxzbEuMNJHyI0DBUarR+L0
PEAViScHFWuNZ/St6Ve5hmMQl+RVLLNGG8QT8yIlwYCbNlE70TyqGc72YywLWbEE
C2r692GB3SiBd6sl0AL/JCT+AfuV6sUpjUCfpS/fEqB1dyN7jL0vPifIiyeGMtZ5
kdrCzgPBkoiTLsheZsrTwB104i9J/6H43tH7Ud2Z4m6qndad5y32Ea9PcT7oKaYw
OlAXk6BABXtkTx7HoqOuFMW7/p2qB0P0gPnDpxE9Lv8W2yOFl97d9C4NrDWZhEfW
reoutbDY3STQdjSGWqPTzcHh5qH01mdmXI3ZYQgZUxvLExpyrNeMlMkFTLVOarjB
LdidCP0ImcmBAPnqWob+6etO2yyE/pRt1vnb6778xKOcEAKRa3SqD9tjizMPgfNW
plhmp9v7pPtZgBGtOSgnqcSlyFgYG5lAD4SuJcQZcjV1h5eiXdNOai2F1fWA4Rdu
`protect END_PROTECTED
