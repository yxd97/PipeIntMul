`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UEuKyUwsvvw1vEYVRQpIiwQKHYad9dUT3tZAt8LEW+wzpYYnA3pks/sQjpineVnU
EJiOEBaFrmVVPP3nZjutmYt2knAb5/NRAe5swCmYJXtoVUsccDpvQOMTD5kXQ186
G6OvrJDi/bo3+DQLpxtsFIxdxjjSglHvDEdN+UqRWGpgllQ2m4e5MSVVm+1R3nKL
cLCAR4AbucWkB8MD56T41qAfAyIB+0OS2iVQc3Ijmk5hlMpxO3azUDRs4XDrKd3m
NJjoUhRpPDLAGwiqc0GH8aa8WNrnhvOdBlKaEo+HbAU9PXM5Jp+20axSf03qKE2/
8WNi8/6hDljSw7IixS8smxJDPq3ChM6uk1OGrJhn2LRMSmNT+mX9oEClLA7ozaQi
eGJfFTO4kEXkYOwHI3Ia6WatXp67iMqsTbAG9Gkw64c=
`protect END_PROTECTED
