`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y2c5qqSMafRlHa7gamoI4ZCT13PKmwSEMQIY3E65SQvvGnuTmoXeSjwhRa0UxTr3
e8diN96eXEOhqEtO1N8wkQ2SP4GmaPA4jIYuscvVxCcBFINMLTmwY9MeMBeE7m5j
6U1Bbe2QqfdsXtKK+XHVAF8+jAAxMLSH0OP4eBoW0QSYb/qWRHm8b5DKi95DkiO1
wrnMv2TYIlLppC21d4uYCvYAMc/D9pEdHQR1NT9yFB514gOjTpQketCqZ/5PisFJ
7n2SBXU4iB0/Pcsk7wVV3g==
`protect END_PROTECTED
