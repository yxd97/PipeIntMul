`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOUpMyRuWTqqb8FxIzvNX9W2r+ASQ+LZX3ESkKfmbY3PcK4O6NaLXaGardLNJ7zV
s4EFrhTvKxu+LrZ0CUaZ20atOCpo14ThlvlviuMO6khRnaeiBzNkMAVRRn9YlYk3
2cuFLZA4tC1czxo8jsa8KICQY/4yZeNBP3tpct1a4AS+xl1oc55wA7SaD83pcFNk
bwWwvumgk2u5yz0NEzGC1kaopTfja1KaKJlKS4UQIPEG7XNd7CXo0JkbLQsPg6K1
sDonuzPzZHt8MvLLK01w1DPPra8seYhdGYyrr+VKP8AgjyfAkdYafrhWBZKWKXBj
ifgGU9En6xaf/R+DBEI8h29SLHwa6oe4i5dw+ym0Vw0FdSl8p8aZXsjfl/6T5y49
pYhW8HoO4e9PGitDqzVJ5pEzyHqaL3uaFwr9+3rFw/9SxpD9xPWUzM00oalp7By5
aGFNZ5k2H7EzlNOnRGL19iFcW7S9qyC5RSM9HvANmMYhgy91n60i3XeDtVgiI3Gj
pcK7RkgjtoQx2MnTVhe5swq3Mo6C6kOfd9MAJfDGQQNqN1ueMayFEVaj4XGlG1xu
bFeWYBBo5So8T0rBiXOaKxep41ZJ4VeUl2FedidE4US1bKiDxJiA/cgFIpyQuZsK
Wf78CoTfhGMnr8jJng4DZv3S+7yPScmfR3Yi5XyeX/qc3cZ4WGzUBFhbBbAADxCS
2SqUlYrFZ/Hs15KczDvjQMqZl254jfNl0GGXDyvWcPhN/ypOND0v3lJyYMssh8tt
GdvqTZarxMkwyKwoeMe9sYL+DwqGxta31KARwWvv+PPhDpAtFdDuXF5nbeai5u0E
RnhN9yDqN0GmLU3f1jKA5CVT0y5BpcYfAv/zFMSZ7sAsqLBN9O5Ab+nVHHsKoPWR
tCzeWobQTd43XevnQVqi6vB1mvzGWrCQPNlZHaoYZd9q3v7ghdhW8VfmFQC+Gw9W
Oq6rXpHXXEw6dd/PeqtV98mt6JoSnpTUXaeVzIy4v5mJiHVjHVtFjeDlU+N7lQI0
m5t5+sgGPFCTq7len0FAaK4gS4j+mt5EPKLgSPh/r/jyonlWdVugm+jMeyHVNNGr
41MjO4AG/smXPzpC07PdjW07IQbHz9b7TVBD8ZNvd5nzGHv98ei7xQnORbyynqsX
`protect END_PROTECTED
