`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
21ZWEB7Hyg/9EectJpUehnj7cKCAON2JH5G0yHuzN3UUhXxH51Irb1RIQNbvzXtB
tSAR2GpnTCfut+9AfSMQkQgpKlzr9m+qWOCzaBi38fdb+aod3S51lZd+HMyW+UBK
+Axsvsmn1CtzivYHRvRBxvjx1k6R6VdiXe2ctG123w+wpUZHS/xaBu/4gOEyEJjX
I5Gu/rDJu79h6rFpJuaAyFrd/YduO/dV8FN/tylnYm4NMkyO1bxviOveCyipcy3v
hUITVkUw8LJIhj1qHRd4Qh3c7GbNZj5Suz2eNyCXdAYhIe6eaXzbpvtkydRFsEiJ
D7uu6huzvEgs/LbnJWBHo+AnP0C153LGoWTpfumQqcSGlwzJBQFVYeJWvAQKlFpR
BwTpr0BX84WeTdzdHpAHzvlB6UUq0dQo/OSoI/+FjfcxBnav8PmPgRQcahp5XLFh
nxwCeQJO2FFBFYpRxMpMn6eoUYnWfMVuuiGeHDe0f2VkuMHz0SHBEecZw4dWSMnH
ECpyP64jxqzTN+qOl3+x+/8CpJNR66PMy4L4GeXMnlRUrrS7efpjnhuQlOha5rJ+
qKkmbIUghkSteyyDHo0jmIDhSuwKf/QjfrmiJysIr9ZEKti0xii7CGnhbtFZajIG
L5d/w5E1NbSj+3CUJIVbko6y1uTBvmljeLdxv8x4JT6Wh2XjCzOtHyFXucUk5LK6
76/O9LlDkQjufBWcUkGBPAvBYuTJTK1qaYMQrSLTwa01jsXSShzqpm1aEpiEVHZb
BfzAp36gWUfySQHDKFITpAe/zBM49JzAI7LG5NBLrDypdfCwjdSUCkuALxfGofgW
Qv8Re6TlAD5XRTGHkRsQALG7lozirBFqxO1QPdhRYFgxIIRN5Se1hbu0ybs9hjlt
4gz6fHtWZi5lZHkJ8fUGxQXCAZnrWGYA/b7KrjXUfNA=
`protect END_PROTECTED
