`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wbkuYAywKBOh5kQYLK2c3wRPwCwCoGSbsKyWZJdA7wTVu/ERitc2lRoeBgoppdfG
rrGIWLvHqdVvKPwUPsu/jJ6toOi1i0+uXkH3D/ZiSpzUrIlIUgTbWuzXKZIPdmfN
TvkYW9CHSx/EIary/j3/EuCKWiZWwSjFyZgDs7xnh7DHe7xIixBxmYHShYhTknJ1
pPiSH4D0wsK4u7qU/DvbhOoR45Dij4SWMKp5kSQZQ59HerDfycrjLAGKbsJ+WGLQ
gT85QEAgrLkMPv1YcAr3vE6I8NcZm3GidXvx1XxSuk0NNINwmdGwKjbKhnDIS5xN
LajiX/rUiUObxQ4f4x7VIA==
`protect END_PROTECTED
