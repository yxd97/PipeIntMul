`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B4TWD/juFbMaEpRrPtDjb0KxvLe4pPNmdsp1h4EYiZFWZxjle+/31OyDarul2qL4
wyyyqqaPSp5GiLf4hQKSijbG4sbnc3h9tzPl+XE3F22eH1qqHrujnXiKZHZxaZ+Q
7JbuZupStKVLqj6ZFwfXG+297qMRY33eMXGERDhLtfMX0n9OJVK085FZQzBxn2uQ
xKFGm5HX3hcl98DXHBAqm78OCBSFfzfb2izVqKBpkDAXK2v90hgw7JyoqQZpf6AG
PSwNuo3TVQ/UoFhnG7Lye6HPXSn6hfj2ecvW0o06TpVC0F/FH99/Gzc484utfEf/
PSltt34qW8AeQ6bZ7bHBnRqHW9SVJrKQzFUnlF1MOnBhCQomZb4PQO1IVxrtOKdN
6RfPCyjPmyEbrmZ3N8NZ37P1auQIYw5HnBJfOYYOvFr036FBHe8nDKa9fPru9usF
VfeyXa49iZ5euVVTZUcbHuZnHjZ8jVlWrO0+QhyN7/Y=
`protect END_PROTECTED
