`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W+ZgnQK/4t35wGmsvxOFXLkeLMd+ZXSRjByXiHbbBtulhWa8atFjpF08llhbeDCP
7J8F7siLmIRKu6D1AacjcFU9HjXINqUFZNodjEIyp9ZqJJjcU3jAfJTCQyRYBsNM
TDAWUIpwTQ0dUjIsUjnO+sV48/DGb4PMV616hwRbQHlXkgx0b+dJMgGomRvoKKNd
g8E4n+49jVtuuupvngiGjaxAPsVys//96qEnFzwwSGZWgAMjMAgceJxDTkvm/u8q
`protect END_PROTECTED
