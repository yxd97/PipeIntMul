`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lB1BPZy4LapmnYWa238jXmR8FN8iTVLRevF0k8dwPi11EeEWiYIseN5ZjhiWZwxi
JoCnhDJab9URlL6TRcUrIwKvCiRsL4PWB3KZ9pSt0nR+UwLaX8LKtwg3Ti3VsucJ
RJjXaNgowFontTVSNCWD6katgvVdrK73g5eYltOwTkPPmx2Le7a9hxMK1l9+uVQ1
YUZFR3SLctruKcr8xYp9cVCZEvAqP14ZnXYuZnA3gJ1P/L6m9sKOBWpTamV01iGB
5Kki6XgUJX94/49AXtlXMENRUp0kS6V933Z7I5V9wsvEJKtv6z7+WiGtX+y7Mu+U
mLOMervx2eQijZVJTaFGCrjJnai90w2AG/Nt5u58DwlbZMoql2iUFfgDMwN4OpWX
C7XuWDIwWO1mtPBC0yMRBtW0F7VqMHOq0uvdlBqs3PQ7TnoMK+jSBeMoONrAdt5q
x1OFjdbIpv44LYjvvs5ajOgEA1fpOoeXf8IUKm2RpQyGyzlv2KL5sdGPCNvsIFXK
0pDunKNRKzYut7xHJT5s0PA3XwSVEm1I5Ao2JmK29//pjKMNA/6RlrqL20MzO81d
j1UmllbdnA4VMNYbs0Qy2gLQxkOIcxG5fdHue8hRXHtAz/R65edbsGoW4SImOsBp
xBvyDoaDnXEzf3BdRHEoYg==
`protect END_PROTECTED
