`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K766kNxb604ZDajygW7CXPAugQyzOiciAGxFCT2UjaFs8kW7/wMiZciIySIuYjzT
7bTtSW2niS0QolkukUOhI8EoEYXS+4F7aK2RAk+KFNe3EHO2ry4R5cudaAA060LZ
diOXcedUwiioTrNp44wHhZNfnRTdtrmb5bDzaJ5jyuDV1YootyrFb14p/u1TyzgG
j96lw7zEGacih6U8i+4ARUpPSde5DilCcRHQWx84o0Taschs1cUUlefZzEKu18cF
hTQhkuwOhnwmjRqNee095oXs8yRSNancDEjCM2cr+ol4P8CnMFocxRq/Jwvo24Ek
eLX1UhQ5+X72wFy2DyZ30uKegcsRQtD0rqT1z9ISI4wU2C7QM37oQp509ApkXXBh
6IXJHsN+LjXBr9nhWiDJsbXAm9Etua6qVhXeZl71KXDGH7ONdtBxT23be9SgfUFp
74RXgKUZ0YvcXp4baO1UC6harcbV2t4aJDPG3HO5jSiQeqBrV2CwOg5YZCl72N7C
o9OeCsoqa/EQ/rIs/AE/qNw35x8rCUsBPSHhY3jyGGQLYTsYJE9iiegro8I9MCiU
`protect END_PROTECTED
