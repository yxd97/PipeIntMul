`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fnvSY4H9CoydKd3z8qLyWOC3JhyxLI3S2z0XFWpaG7JgmN/BaPkXUM1900NxU4c
bk5NvlrTyh2J5lhfSq9pmoZsk+E7flUK2pasORmahh355bVTg6QSzkC3rchcNxRy
uwlXWc4D2oJxw8Jt1qxqed9pBaOo0uF3gc8QfoaY4v6qHRZdiCQtbshEgYIaeS1R
Bbu0KYy61Q7sbzNYo4gFCt9oRTY/hjMosEJKAzaAORS5uhwVMj3a0WHafO/baVNr
8T6A7DK+1bFU/nMJx4icx7LJ0l2bAkuydB598QXnKWg1pOFGEqFWkOyoIQzh4IYj
MT/Y4PbTHn+zzIxBFee+9ugGd+nPWviHu97v8o2ArjaXQtSL1ICkV3XVx9zwq31R
gW5eyz/r83/NnBLfjWGj6tyBpv0eOEkGDOCO0GCT5ZAYurmIZccTEarIK5fY9H1Y
39GDZYeiUOikETG2rrKmclS4zCraO8hwEU2vgU2VO8tbNXtl83t8pfO6NYx2UBeu
pQkZaMzDbKCPB6up9OUUhMvExyHMSApre9upRJ5qY+ihJpcan8k7fSoeigSw8Qha
jsZ4IiDgk74O1yauRw/qrUrRarFATp0px2mZwVc6MNtr2zRwNoZxXz0UCOCjMLsr
SZefEmE2v6FEqteB3UHcWspenlKZ/gzEUPXV8Zrlvh0=
`protect END_PROTECTED
