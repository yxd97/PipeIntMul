`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/uRXxaH6HkrHk+YTBwfiXQlDxXWbi3UC89VeLKOYS7cccS1BeGvXZa5zREptwgNE
h5ibV+IaP1pEgP72vnlINIWFQ4msO6k3wHamkdoiRb9ZRGoNdzWzqZ80V63DP7Fh
Sv66N6/dACfpXrW+1e5UszC9trxyQkTlo9/N8MWYYZBctk6vkH42kZ4ylreI2I63
0w7f1/XIJCLQ94bB2fzniZq8P1suqmwAy/4SBJJG2NzoIrileipGcpMc6ONP8siM
FdOqZbEOY9FpL8Yp3gnMbw==
`protect END_PROTECTED
