`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cqVEf9/2b9zAvCIAAvJuNYmuDjUTPInzIaUrjGJYCty4NTlusX+gDPK46duWJ5K9
5aVfvfRpEqPS9+Z2FsNmDkV6mKzZEfOpALUhstIUldr+qqccCYkHpaByddzrx3X5
5c690Ao0GjPVWyPiEG04QUiH/EWg/PukLtMZJ+LaQ6/7OsqUwtxEFu+aGtNqrXu5
Vdk8Gx39yCDGLfehcnoD1B3H3FJCdc/EkJJShUfyPErsvxxuy38gotymUbnzwBIb
OEofQnK/nVrZP+DMshBDMwx0bwLNxUobOooxZWUjyP1srIcfdQhmXPfnZjA0VsXD
dIu+Rn9fQN3mPOWp7ND8lvM1cnT0imXqRtUFEjMY4sLnAc0dlR/fb/rXEeeQ4+3c
7sGYVv5RWBJxvZkzh0+oB6uD5uMP83n4HFrmBID/aAWwXdaygLDJbiG/eOxd8uwn
Z1CVlZiTh/nfsHrafn63kPpwUHLUL5qddtloqLH9a48=
`protect END_PROTECTED
