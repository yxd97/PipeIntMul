`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R0wzphcMoSwXrolASbsjReNBDu+uEUyFjgZGVPJsoQAZ11c//vCKV2ZjjD/r84SB
FQ5flKphvq0IP+fdHuCeKkoP1FZCgigUewNC0QuSGE4LkG5BTqMsUw2u3BoR2jvl
7K8llkMN0i30UCdrAlBm9U4lXd735rKc5XEnEXz7x6mdvoJyvu1920wlEjUwo9eN
iIwqCLs1aQtbA/Nzt6fP73L/vEGOqMDxMVGEePsGuFRkdZzCjqieJWdYk9ulRGRM
E/mGWBNtBHSqW38h90iFLL44URjEmH4rkumbc4YLTiCCqsOcYYf7h7KsKobJhMY0
KNos8wKcvpG8i1dARVqMyZJKCWFFlih/YWPm3a9rZ8OmCbp3MnFyWwGe+/NgPehh
fQEFpLfljtauGVK9G1PMNi3mnPihrBSzpeGuX3/aC1Ce7heyUrt9bNGkdv3r8/dP
jaJVGNH+ReL4aK9Q6TRbf8Mx1s5Kd+6hYVCx2Chk1sLggksY9IcRjIAyjI8kuiFT
qpeluOltIkma9Hr2iRMDln1GvqD29B5ZVGmLa6As7pNwRHnv1Jv0ay/5KsmkQcs3
UNg4JA3MPlQL9utIK8ZOd5bK/ovMfRZ8D9r/c1NqC1LPsQSNMK6aTa82jaLmj1ig
xRgT0jOQrMfj0Uz1x7i3jGPbuNMmYp6DsN1PFE+nannSgw8PC1dEv28VNfAlDTW5
VGM5LXLdAuYqIf9XeyIlREsuWQH0HSNWclAg2f+0Gh5SIv37BF+Gl7AHiiuZTIG5
7ycroE8qOG88tjZz7uWUmyW731oVlkh2bVKi+E5xsrQKuQx5Pf+ipXZt9jKwLRrB
1TXxvbpSatE48+wx22096gdwIBIaVhBuI1RPzOjXXTSwaLjFuYtONkxah++NxKtf
xmXYrP4SvTXqN7LwphB/njeNEEtsHv8eZh8V0V6p0iGy4UcxDUel/uO1jeSZLPxv
/PHINdV/ta/r0HGeIS+6B4t6CAblXyspmtxhpTnGTRhsuStsOJUVGEkbud8wyusJ
f2vnOTe7ls9SED+NukCNkvyrcIGKKvKYu+8LIqrJZNdcvGlY407hsoHEdWIl9dNQ
q924ieje5KOb6v2U80DIVoYyQluEA5HsNjitxPTkn4Y=
`protect END_PROTECTED
