`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ypyVAX0PjyubBo1pg1Xsa8HdtD4Zgy1BRq323+dPvv1G+pk782hat8Bc3DH9aNIy
5HrGmUZcllCZa+88KVQzCRYwVelK0tCYAjcYqKzKyBDGdY9nEhN/i2UjTzlsDZqc
L5iK8tsDPzcOLkOtriujhQeyePYHGHhDedcT779ni1iJAYAeeptDud3h1lwgFVPA
DNifoZa8/KqmDe71gW8iWMXBF4hCIOPhgosqaCyRe2ugyW9VHlbfVeyQnOXeJhd8
tClzDiIhDi5tMVqcT9G9tQ==
`protect END_PROTECTED
