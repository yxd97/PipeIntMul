`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jvvDIIQmqHFkjmid9ivizqetudBfZDBY3ifbUFIU/ZmTCGsApdrkVf30q49Rr/VS
cqsxZdiwGD5lLFfHZ2QNV7/fudiVOiowtMRbxIdBMQpGD8Gpuxa8VrA60fR40tGI
eQseVSun6gELPZcZG7QFXfH1qBN/Ix1f7tLOsfbjvyDt4yGjmqRhssmGIniDu82N
RVfjn7Y/KpbRvdkmnJSvDqJfti9CRPviLEBF6+2qwr7OyqGFverncrznZRy8qQWn
eP7cpicJWO205mJNVEPPJiJcyScbibUfevPVOU+juIJlI880IUTbyzYBG9YMprsw
5khLcMUyWJ7pc7xoFObrgA+1bVBI/xSeKMKpqT8kj631Debl4U0qkD07JAp/gIZO
NTQw8zfKgSkjFtggvndwfcfMgJbT3RMgspweYrrd1YUcOyYzhDA3nXn2JxzwGMeh
BggOrdAD2RGa6AV4qRHErTv0Fp6u6WGNxFgaOFFHr8ZdlEg0o3tSZWoXCyhwCn6c
Wd89ygEwlec4LQorNI9LlFXaLfoP0GdAImyffCXaQ1hdgAo73Iek6OidJgNo+whv
VG+ucXNMxhCDuOYTgrO0bAX3laEOGmxdUUYs7CCYZWS5Wh+blNr3tO24QtFZSXth
xXrFjjgbRJt2kmpM3+mpMO26Dvbjk4zOaJH/K32YCdZjYr3AvWf7Sopv4nYnTdHS
5Mf9c0AUCaMOnbSRt2fffkcULtxhJGuAqO+3aCr8pdyfezBOW5uQchlO+KvQ0B05
JlikjWKIkNm5M+bxzUt+lx+MyJolBsIph1vEbmVrpNho0qljeWk/vnE3M3gut8Vu
VZk8lx1V1ti8zOUF/oph5wnmWMG4y05PKayUW1iq60b9NnYNDBPWlO+TsVlCs/3M
Uvn7Fh/LP9hN1FgsPNxfx/v69EgjMuIkq4tM9xKpubochL8A2OMJQvLKY92zXdw7
`protect END_PROTECTED
