`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GCDRQVZYDeebLRUpdcA+JeLIm3cLzZQqDyfkkH9gUyH23qpyTkmwfZRdLS6zp2v5
Sc47mDfPfsLE2fksor9f8xh1r6GXsIMrFKzB2sWzw9tVdEfXx2EkH0gZuixcs4gG
IMyWpBgxbVpmwpXz0LEFUu1crpkvdp6GHfu/Wzfj4QkS5aTVudM+tAB1NoH5RA0U
G+FF0ZC7XN7asjDAZTZCknkoWh8gCJjAlIbS3uHIaAMVZrFh7SZO1rCkIEytBVIV
1M2on+TRV7x9auKiTK7EKLVFzCi51jzVm61z3kQGne1ZEIwWTADo05jfIDx4YkuI
DwwBV19KKJzyKXhZLGwo2A==
`protect END_PROTECTED
