`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmmjgfjOSrkjhbyVqusThyBnzNgCheavEAOWQzz5FO/Xdy/c1OlFjsFYEbNpQjZQ
+Tl8ZFHv1yqNu159lcXqc4j5IBSS+LulEEuiPWHe1cLpFIMTBs1IJTZ4O9FSrkS7
hDnlapqMNy4WIy8UExR5iyIhRfV/yNrDly0i9rZVyZ/IBqvSYLtQibl5sH1witY3
JpJQ1O/BKRjD4aCtYaWQnYJHUIDPdxcvYcB+ZNjlsOVT7wvkHO9T/4rlBUJK7iuN
NroK9AQ5y2ohjejLhq/L5d+i1H6F5sNGCXGCm1O6+DfZii6svvDkPot2cDHqOnAW
Gg1ppJGq7ZdbRF6dROiQdo6OMeN7eTvUyH1PVdzlmA10leRHae/TdiZ6PRaIRybn
51xb4mhqFYlwT4BOe9RAhRkzzbeK47J3f6/wHvKoiH/+0LIws22ZFJy/wpQLadq3
T/+7p2QABd8bZcDN9HtCtXki5TNhMLKcZxNbQyFYETpvpAlPvNeRDHNPXmb9ue59
3azDVVL3OElbDfZdSr0DJSuH29RVTw00x/I6ixy5o2p5X4/z6t236zF5eNx6xr9t
OvC1kuuf4gDRZFyr9qGOp1e/XFwWU9uLEKdUhWKNmKI=
`protect END_PROTECTED
