`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Nb/6wk13A0wttiMExKxhYltPwCqo64zBp1+8D6rU9cmKKVG9mUR5hMDqJgO94omZ
INeg0ryhyplYmpYquE2MKD9XQS20RcH3Jt91mzVRpal7urRP/p/y3/2MbeP2uqQL
4pjF7Zq6kgitdeKEikmA4oelGkfIhKRqBOF7b96BB5mBZtazQbQVku7enUGb3IQA
FLamilvioctnMnHYjzovw0fY0CD5I9w4P2vc09L+rxdDYEyybkBS74TQpnYeNCkL
eMJPr0dy/P0qma4Y//GYWA+yH/JE7efOOyEN24sM68fVLDsxwPuxorGAIJ+CpVhk
PifYQ4qIvhgHs5gJDzJI9fzPixik/1eQbTdLw5GXKiO4O+CSVu4anbOlh4lnFsA8
b1Gbg95Gv5jL0vzcs7KF/AdR4akbpz4cnedGuYAiGFIIk83GMGUQVxn66rLJhHYn
LOy76knM489QqWP/CniLKU0kaBUYe+iWTGiYgHuxbUAK/wpw7ZhnhswYhWrT29NU
IC1PEO95cnrEviYbpWGv6pex1xMB/8LQnJND/2rlKmWtEKoMkQFerPMg+k96+pRb
`protect END_PROTECTED
