`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8n/sPDRngKNljGbWRmGnmuJUUWmmUM6fDB3UIBrCgkzX0U0x0to8uDdrJYl7qUNi
ImCh1Dq9fouccFFLW76DDgk2Ep7bSbpfPzgiTRi8+QsUtJ1qpyHPFAuQZbME9pAg
li8ZyPwwu5yD6EjZgKpXA1+duomlyEMAXWYoo1YC6Isyt08zCA1CWGbRp+P1S9aW
REW70i4uP/CnMMau+VLzOVEF87zREJYwLZ5XjdLesUFsYA2nkK7wmJNcegWQf4r/
emz7ZqWsUoaw+rZhLnWNiHuRy5cseQqldrZdDgRoaAAcYIXpeQuncxGrfyB+Skyx
89VCvDn0G6sYP7unCdI/iQ==
`protect END_PROTECTED
