`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9H10DBIpQDjOM5ClA+gM2xM+Rd9HX5k0ooyQxz1odZgvhP4KUNyWaHTjibLhIQ63
rqfRBWaCz8wu8Nq+eC9EtQmKskrCxkINhcqhSU9ozqsmq94DOQIVtgjIq7AYt2K7
HhMVJLS2S7Mq/Uj+Zu7Q+qutSou+lPGis9CDI1HglQQm4ivyFtuHyFlSKRr9xBD0
4oJ/HdyQFlwy9qz8JClHW5vuDUyxdGQMBJnAU1Z0zGwG0ErqMR6n37tC8/tZe9zY
DQP32vS3E7jls8ovi2XGRx3M1llICeBlUDqWdl92no5aB0p9mbg5YSm5Ja+Otd2e
YZCG2o/vTEVGsKSeahLc6vE/5EN3MxAk3VR1WYzLIst98Xm0PNI9tJIjKnaME6Xk
dgUounRsksUZX1kyGSCN93ZsRieksEhC5Dhzk65uyVHJs/g8CvEZ0oTnhvI1Enwa
6Zwf97v3AHyKa/zS+DXrMXAwd+G9ZKqT+rjCGE7rpu23VU4hcBXx9gGKnVdUruLQ
iyLxa6pNB2a01DyGqL8xOcD+sKcxss358DXqCd0fxCDfeLhnIiD1WsSfGaKy8LfI
M5XmR8iS44ChzGGADqDbY2SXVeGy3e1p9u2t82qmfO9lmmjn/8+jr1MylsXHFEgC
LohSOyd7eZY+z3xj7EB255qwrg/csblgINHcABawYcR77ET+CZnfKUesTopsiCGC
ymLvEzx/dT01/VVQrsnXhPf92QXoAmzWAt9BuAbJehg7kJrYm0cvWK9KIReBBZpa
dei0yO6ECAkkFjAGBbjOvPMvItaA98BgTTZXPRgjJonfgc4GqRkqw0l2g8D1atF2
DsFc63/1KhIwp/b7M3bOd6QDZhlXS7YfPNAoHl0JTElWVeU8ivRRFmq00YSSrJPv
H3nHB8g4vDHjhQfdVH47uKE1iLYrNebDKRdqJ5xxO6Rz9Bcj+Q9B8Npta8rtsSmD
ZrvI1SMyhdRsGI0SagcllRTYuNZly2cJ3SaxBqdmc8zzKIkciORYF5PfM4SMdvOZ
n/3bvUHaFXgAWCMW887IfpGSZ7FQTC0cGGdMTD/OWd7nKsN21U/jLxBkWH7xZMgM
wa6hDx1pJwZvoetc76xL3G2K1I3owh6Ssti2vQ8G/5CElqdj6tl5odmFcHl0fUNb
ITwTGEJxF9+ILwsT6ERf26denuEUrAeNUXTkp1jEFk+sMbb2E/ojLJtZRmWzSkpq
dL9idAihN2KxIw72dMmrnnsWcDh471te8bjUPSNgHf5oO7xa0+NZul6h9Q+q3jnC
Xi1OylCvqG4OrKWG/28Rp26kTX/3g5VfQUFPsLXx2pvlpxt7JITjrdzP1FVhriJF
vWTLVLkADDt1n3UK06yU8qzK9YoQua3mwt09B5W74W3zKUgy0KGle7FDkc9YMgM9
wGGof1sHnH1ew0o+PTxwwKhrej3eaN6ieHnNxajUhne4rP4obuReCYVNIrBOlts8
OL1dtvGU78uSDB/Ho1U8oMStpk//iabPWu4gw0sTJBnxSXdNrUMh3w+LykRJYiqd
36lF3HPNvABt3Gs0gupGB/POK2LU3iY6m4LO17XiAcvhyV2fzCN4dAXtIMi8ZrdX
fozboKIOAbK3y6J65c9bmoZ+dFOOnMUUjbQERwByehrAJ9b3j6McGShOz31psCRT
awY+FU73doiaEdjCh8tBCnlhuackS41lo/UwWCSZTRxxWZhS89MnFpHPns2Jb8Kr
GU/CHq8JG+Y7zs5uLQNzrxAu1+VcP0OWC+s7ZjhkVc5ZoaIOqcNY6thiWhhlraFG
Nf6Md16GjuPPRyq0ZvVCf7WljBv92r+pdW+HwSuaV76nNxJ7BNZMGreQKelzEH2/
obn/r9m+0Oex+hoWwPksffSYU5BOMnYM+UH2Ib85xmK/FIrbSkhcvbRmmiA6tldp
KRVqovN4taNmkXVe6/LtfvFc/TkRuH/LkHD1yuMu8/iuZjq0819RJdugfWqmj7Qz
GnHyQQT0CCnT6+2RaNQoe2n+5DgVOPlbwrr7xVEuluvq44iwbLFR5NjXWeTo7FYZ
hZWzO9sni6wDF9sVSOYvKyh9V5oud/ZNwY/ihCA8rWJRU5Pb3MKYpykZFqgWe2KJ
E408200IPfCpx9oU858MDlxNOyixg46xoFC76YIxP4426AsHwaNv5kCZV7K0KYXI
reWjBnCP82LacHdndCvyptuq+OduwXBst65Tx/5jDKWhtWDt5ZqfMUgCxM5Szgrg
0ROwOwVzA5PCXCLEJV6mhZolQhVfZE0Xuembj4v1p0psQf4Smk5sJe7AI0wFfGtW
plJO36xLyJwYSZ5mupZ43dbiJdfMQPdGj7cKV/4Z6UVGxjIoRXJCx92isTYPjK3E
xqweCQ9K15lQBeLp3nXaxik0BT//GXsCarta5u6jGLQRSObr+3y7qNSsxgc3cXaa
DsT9v9+Z6LLkhWFCwusbI4GTxaJ9NMITCFYcCdfF4jPMVgkTDCqtarUJgF5B47np
BUCVdpYdEv25FBwYdVwEZqI5j9GhsQBvv88S2TS5mZWOeYW5ArFRbFoKEiG5xXaa
9bo75qJMCrkVdqTfxOIbypMYfoZzcHheCiE/+0qzAwvzU/2mKarko0/GFRLOPsxM
EFrkGAxZdlWSawVPoCQBOK6fA5sUG8Zk7MKc32WZ+i1Rya9fmEcphyjUTki9MaTY
hRqYgknOtKce8gKH7/dyeM+lMMWlyfzYQWwaEt5O5qux/t+Msa84Vfp+u04qUgCK
YGApJVy0kjXZS7+1s9KrgDwYIqZwoSbu3FpxbV8HytAUI8ChTxuElYTJle6TI2dl
40YE2bg0k4hWbfibsuREdmfNhKUOOuuwle4O96kIUNP2Xa+X5PoHSxwq33CrUqP/
yjq13hyHVUZZWQmxhMKQByKDYfI47WtzRwmvwN9IvRDBtKBZWxPW/bJb7ciGCB0e
Dk7YGxOTgNCbSh/JRcWKjk+YqzFX4Fef8Qa6aziLS+bFvXV/xfUAz3OxuAo9IlJf
XbSpafP786qexhJvtsBLIFI98vowYRNYi/hN8JVdTIzecZEHyu+WUIchFt2cJAhm
ffMJ+EZB+m2wsml6b8tYT2c/c0nHjAZzCq5IJgIOATK0OCi0l9pJzmxcGpVfCgww
NHQ6mL8IuZx4Jf8lZSKV4hWNaH9g/csrlJNzobAqlxVmTk3klRzfpkO7Ti3ToPcH
PiT6doZYUrWMEtGB3ny0VVZTdkzAsUDLK5ZrMfno0AtIwLQ0HAgCJg5BW2ZI1DZg
p8uFkL9YP4wZsxETAM+FPxSA93wjQHhzBLURVWz2JeUAI6JNKgkcB/Lmk9RT2qLI
bmnA8oR9/KOwbdgjXbJCQxA3JUF9l2ltfr6b3s2qGByqa+PWLA5hnNhBCz2V45aP
rSO18Sey547m7UKcyshCnW2QHibjDVAd89smCvFWSNCh1riJUJuJiDq9q24ttBlY
KjjPaUtwdNC9P4RcJdWBp+QYWbFXlpA6MB5R1zcqs7JPqS3/BV0im/rif+qdVr45
+P7AvXdVSofK+BFGqRDebnOg9Lo5mubT3mnujOs5e38YMSX1s5hHaFsAa4t7ITxv
dmyE15QVhNdQkI8GxI9TzncABcSpV50nuDa4tzQkpH+G1KTv5a49w4UV+bfmru84
3kUsq/ZZnB3Vk+QUfp4PwPHnWmiLMhTx8oI/iEblp1ICpK+YrbPurLHMI6beKQ+Z
W8tsppR958s2i0AbY/BLRTAlHxNn8x7Y7mofn7mDfIyrYmliPn36ZJ5xRKEF8nY8
RWoaKPLPrH0fzGSDMC0p+r2zJLqNllAKA/X88NSKLL+tFDhOf8Ah4ZpLFaC3nu81
KGTQO/zSV4Zq3YaraN1B7ufwC9OjZXbot62/o5tF3kTkBln/jD5DLBgwAHBDmo67
kdjI7O99YAuB4X6/TCL5MPO7qEBF2eHb0eGFMH70mg2zz5fsN9imIK6+WKaTr+Du
9lrdLkE2pAEmmoGYs/C1pZNsFpU071Nl1WvGrNNpJJ/3vcxjfRrEB1S/EXW8/N96
m6sL3nFmVk3CrT2Awq3IQju7+XNlMU5xsMGPGUcQbWw9iy70GtepN3OKltd4Iqiz
21vcLWvUPy8cZaz3uU2Flfjj+gUYfG6sE4YRrGOK97lphVFJyn9iWa0YqTJmT1Pa
CIeqV2+0gdFUpuRxKwy/3Db2K03scmjc5hO/CMvPDj9tLox5vt3lD1z/a7IFu/TE
aZ6ZXDCZLbvpBB4fPSXGnJ+Rak0RpUqAsRVp43Z+NgeDtYQDaginZZzo7Bh9zHht
QOG0D1hOr3wnZ9qU15AkJxqrf8LBqeZvDkN8qAC5x/XtoqHrcBfMM+10aaSSD9fL
tFBp8k8naJ73jNufaa3/Uv+jX2oY3QBGxi4MuyCZ82FOTaqK3r3guNwZl3L3dSXw
HCw64vXS2qHJd7DqHg1PPuVKn0uzgb4c5wcHQH9tkN6kIN54rH5dR4BNlzUcyTPT
7osO7mIPXLuaItJEDDQiibzwkXXzgafmaLVJnvNUwrR0zRz8GMumzLlw5SXz/xU9
veU/s7rTdwQRxE+TWINWObp2GjH9usZAcYtykb4CBsWu5BI1ilf6gJkcUHIASgQk
bHT0AauU0qlMm64tXVruviEjBaKMxgJX1FOxJMOBxcaVJAUTeFQWQymOTHDIeEpU
t+JhAcg5amg8AbGM0aUzJI4gWI4VnMMj6SDpmZps2xmVfA9ZsgoVeDPsCDOVkWZm
naZnAPrCrNIYiqMIzJR2v22HUambNIO22PxoXKIGULYAWKUv7ZT1cQKEAxjQ8jab
S0cKU8IQYd0sZcK0rKr9S2FmyIRO43UkkzjWGwSzWXsNCxerPhHp+5njn/0AoEjH
oRovQAYd1MTUCtw3/R7kpuQRVLvNymGbfR4jrgTGheioZ19J83+MswMgfd43pMJB
qCoPUSoFFnrPOQumZukiss6L34ZcLruL7ZOjk7nlsF0lryt/wRSKBU3tOtThKR8y
d5dT7PJL4zJUD9+xIQFZ2RdpbjLOV9bibBmC/fGrqfA=
`protect END_PROTECTED
