`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CPPne9Yz91OHiemeiXdkq631MfTUHimaN6/+gavF722+TCPXaMvMaIIx/PcaWvOM
wzYC1ioxiOxejKJ7cu9/0Bxq/fipt5dGKI20dLxFCcZC8LvX8TklHOXBHwyvOSpD
g41H3zJ00SPFe+eKoU/A5A1Ph1HDfBZtO81cG3aSNab/5CqpWTT7GczGckxq/l02
EAcXn7ww2ik3q6pPPQ6+dBC2FTjW8FfyDqIYAQAVtJ68KTexk0E/HpqZwrz60r01
sWTjpK7xkqDtnQg8y0y6bF/9YoKAd2Kay/Rd9N5PrCE/mIc4cxVsY6pGMr+Llk3J
5Qa87UeATibAMcwyR5zoAc+deBLPqxqmeksjKSeuEZXzpSp68sih8ZQF32VzoG2w
`protect END_PROTECTED
