`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rHczCvK0tJoQAmZSpJ6tkdxnkCkfDk/m0r9DlwljK+v9QSlt7GJBOudhXupNf3MN
/ULI5gMKG0qhsGah2az3xsBBk8N//Px96c/UptnTNWsrf3cJHwo9KnDRrGTQGUVf
K8fcMtvaBLxKzZu5Wgak+wxeQ8pAqjc+nhw5QNr6xySAGYjF0KU/C508+3CvpTg4
mR86shYNawtR9bB+GeSvf1w6mYyz6qw4ZhE89lSM8F5ZfOA719XHWw/9+dpW/0FH
FMwgSkxQ/rShhFT3zs6KBUS+sbhmpA1wtPFPWbamqb9I28aHvBDAwJ5o1nHeV0K7
shAq6g8blUfMl8slAcWWmA3sDc/yvCMgnu7j5wFQS8XYhal5HmjX6NVthHyTo6mh
2/IUsySNhIzXjtDP2gKW+koLP2PJGps/rKAbc4cgaiBAS7W84/KJ1o8cbo4SGVVS
0yP2/VU8MQUnXh59EJ0Rrm2WLso8zBOpbZikfjkimoR4V8uCX+FwIFtLgoHG0CQr
bP3cQmOLmvgfFlma6WK7DuoSppc9WEmmPkAD7CBlkqt9x0NQ9fRO2O1wXxMnhXqJ
P1FsjSmV3d6ag7+W4jwRvkkumvPRicgQh6doD1I2Ic6ntKo7RKTQuipGcjhAuv71
Vwo3EKrRnmVj03JyEZeLk9+bOPyyO+jdyCE+NdI77deGJMetK43xk1/uqh0qnQp4
4Cihq3HffTtnbR4j69tPqMvYYLWmoMqsHzFy1/mGmQ+21MZwMzkhce8fJP50l4X0
R+xVxTSmnTRCUoRWj2RcUhLUNaMfxAyas0npzqp7GehjSpw7Qsr+ew8ZVzaHk5nM
jZZTsFk+VWQKEI/nSVPYSTo8EdQ7dNsEbIAAMe9RDTojMmH+As6ttSkkZVHr518A
DOxoP1dnUgpKCEqpvbVNqIZb4qhFdtNgfyU+JAdEfTri+A/xSnk3SSgqmNW6NFHG
UXpg40OFCq7PN197agURgDQyQdOAH4j3jmRKZHh7nh/WKJkyPnuNjaGXYh2cykFQ
K8cIeWQgWtyWyHre36QQ7LjPw81mWjv6mFTjSpeY4HFCJn6eMHVpcp0xg7CEqWP0
rwtgjeABOBuf+xvWW91K9GA2zEjelnwxXBsWuEMTtQaxyV8tW6ilUayMCQG70OaG
zR/2jZtzPCspi5W7bWsBoo7z79hH1+RXlIQw6AaqUIzAzkkSM/pRQsWxVDQC2M88
U8nOKKHt5ReiXo60KWO0arLzGPXTUuhme2C0UImdRl0a7LU6lnMGlGU/d9CS/pM8
NbQnfK7hLXstJiOmY4fklDfVwBIgul014IsXkr+2KzlZStsA8+fLu1SjqoV+MXvX
zLPgFwBU8iDHjB+9pWp1OQ==
`protect END_PROTECTED
