`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ynHSUkDoXt91f5/WSkASdLQXoNctssFtE/56T9ZZux0/Dt56BTC1BbfGYNDnF+Hr
wpzTevo1znP0dpXupqseMUAadx+v3yiivqelBuWGCUQZvXtQMn8O+RbOgKGJ7veQ
7hvYiipLFLUS/o1qtX+sQFOSLqNItqiU8iA4g25BaU+3LLJZBx7aUlrW3URSmnQ1
yUU2lJKcWDq2bia7dZI/fHeC/Rhji4It1jiDeuwZQWq2qzzah+rM4N5gloUMmdPf
`protect END_PROTECTED
