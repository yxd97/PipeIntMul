`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Io4DvmLtOADDxhuv0dqQhKHTJUOhY7kjasN+mV9KE5MzML36eoMBz8we2QkZ49t
XXKkH7dQLBPd+zy2Lou1HoxJJhh7Ji2RGnwtKn5prALI61R+qPf263ELMqzKMuQT
A/UvMeDBdeJ3L4yvc6KAfQarAmfSO6ORHb1dtX1UhyI5FP38VfapIY6EyGoo12dF
11febVl886ZoEByhHVo4x8wkBBYPJ8BeFZTgXMHUXvDjvYPJhCDMyG+Db1GOC5SC
6uQKcCdpXUp/PpjQLXlcE5xzqARKSuVIIaFM3ZC9sA7wqXFaL/cZhZCF9DZBbYto
3iExXEDYFWXd8ba/TpCvxdGcSdgsTYmsVVQfWFGqy55+bqWgSdOvqze3gvy/9EQe
Wwq+DaIZgsjWgcaLdp7Wxqas0zh52/IVvxdCeeWzhQPcbFggeEBxqSlG+Cj8f5AK
B9wDoNVe6/6HGkIcFa2RIcpbuqVO5glJznfI4Lm9puFceeX+QQ5Eb/wxpwPZEO6p
`protect END_PROTECTED
