`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3c9JqHhZTmH0V9hcxEdro5auNxYvXp5Q96CUAJVMXGxQWbDlPhQV5dLt0X36s4XJ
T0sfqTzLO73AZveywD0H5qUxT4ZIr7d79HqLOnnTPDSby8WxkyATxZH23yiYch79
xj6zIAp/RrV/S6c5EDchOs7N0bS3Shr2JmxDzCHoPCQPjrxUS1sjeJYIWiG3K6VK
JNxfxFqWEB+4onHbUqo1NOSytPzJp6Rrb5J8b16qt8WNVCDomZSKWe3XkL9zGEhp
uG4RSTspGT0hltM/jG3nxYP680T8v6+xlYpVDxIDWaA2BI3igVXXvPhH7a4cuspt
Xx8LVcw35KQ4n3t1iVx/pufdSIx5K4ELUONX0OnjipjR+kZNlp2WzKNLuxmRdsV8
w3p5/SrS7pgbyjeCbd8XdguMGh5slgWXKksbhoseNcnJ/hjk5rl+eTiyuHZd+3E/
fGZJ141KZ2d0Inr0wIoES1EL9Z4J18VggBCmNdXMZdzbWrKcyl1UISQ9whAe5mAd
YT/MttTtsYgwU6D/g5ETZBfh2Uw6zJk0MS7oXhcWBoMUdkA/xEz62rR1VhBvCBJq
iQgmcnojPPGmeVuA9ySLijgCO3QHMBH4Sj4JB8gfgCKCWCoTY1FIHqJXcM82hL3l
e9OPmgIspQXaUZQz4GHuLMqb6kP6CwBMaRs7il7cXk2tXosUlfEVMohScYC6XLYO
nhwpSrMY4b/x2apyjjkNdA5YB3jJoT3iSVqHzerTErUdR6bzMAndaCym7apB45ap
TMVRLpIus9r/ZJQrM1TYeD+HCzIApTz3V724RmjgsZx0HioGbnfNGPzcdRga9Sru
Xp3Leqip6597m2TGOUaR5tx2cN1BDKbt4PSLxu6zBsxabgCMP6RxiqfhOmz60Q2E
26uw4HClAZHey0BN/KHp4qihgIE1G88vglTQowb7m01BIqwFrmEMO1Li6p1iEHVp
50R4EHQHSOcfBwB0LOrNR4ZG4Ok+xQ8J71s++/IZjJZMpWp90u3E8PXB2DRoZ+so
8xnvOwUINybBJ4o8gZSaK/KT7MEwfG/FiU9XEQDOG7z1rc7UyQ8XhYyhdEzxLi4n
LYMsbYsBy1u0r9d4XMu8PnEBsTJvZZwtDhMOdx2rE4gd1q8WFgygurojr3YgCgZ8
IAE/3h8Zf4x4Ii4RJYRtfvyRvplbuoqiW6Y1yRNp3EJeMuzaa1s6Y2GXZUVgtiY7
DJE50U7eFskYBODJDqH486J7eGGdQHtFmj9XvgwRoLjfm8LeDkBdb6eExO2ROqt/
`protect END_PROTECTED
