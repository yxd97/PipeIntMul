`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4B6pmdzvxuU9ZwqnflV7JQoKksYjfVJvNIexyIwPF+mOikmQiNFEpGQFAHiG+zUE
Ne2HuNwN7XiJDe+gyqyo+alfrTSwE9uz1DXwwOTKW+5kv9RPvQf6ZRIQgCrHHk6A
kFp7ChiKDtb4qK+Jj7TJg+echdEoyu5Tr3VP4oO5UbixWkbEIxSONm16+3YdhoDK
PcH/s40qB5MWrqKRfjgMdacPCVWgYVeT9xyyQZhWdiAQVOhBHfX/UHFSSfw+Ti9Y
xFSo5foMn5Anw+eiGnay+Qv4qK73XYrLqUO8WfpNWr2XVm/g/4Vwe8vhxgmF7Eil
C9tX2bJIysbDmQbWjMM6CzC7lcPWRf2Z63RdOSU5jpgkbUVdQx+9+JCEkWSU2cbm
8UUd8+9EFyv8lXhdFsMII63uM7XBppJj1Lo2cBsc5zu175AsPneeAJCUub1nw3+O
JyHhoG79LBSiizFVlJpnVzIZ5PzTeqR9/xyMBqcFV9oYjN0YC6aGa1tZjDy6+Oye
zGvcs898aI13q6u3HrDTfF1p/eqBquTITB7E4qRZi0C41NGtXifkHnSdnaH9XUU0
4rCRZUBwDLK9iR2EItQSaspWwv9Snt4NSDkZEyH2mqzNHRKzGOyUkBwzhbOCXCvH
aqjwTEGZJZ2jTZKdo6sqX2P98jQxljFAyTLswqL6Dtvlw0P0OcKIM4wmoGftoXXF
OgUIDw3D7CnxoMziw59woZ3beCNeTRjc7iSzSOfBwJt9nKAFxTYKHmgve0/Cn2ZF
LoeGhiJQN1xWu1Zri0ard3Fl1zAMR9Mtjggs69yKFv2afdN2gEIYE583U0iZaZw+
fPdQtk6TImNOq9+m42spuAnHqBus5XFlA661FWkvOt//EthRi4ITye4zi++0DTiM
XyCfrSNDaRb4YnvtpYVipCa1tWzO9fMwpMv42wVVampXpMVpc1rfV0wZ+xwHSFlG
6q/qBpVc5QFvyytJrWRYuflVWGhA1v1fjdtTguTBPeZmc5C0xIPViMSkc3bqA8UH
+EmaromzArNdgMCIVv2Vj5oun8V8MJoH4JuirFQTjJDjLtNhWhjDmtyK8rXlZN5h
ZEjW4PCUHX8Oqg0Esrpu/9q2qk/5Zbi+9bC17JOorAtApIC49rPB0G7ckjDjXgbh
fnL54CtUdzssCr1eE+J1oDjALoKahgJuNo7vd5iAWb8+YWB5clRrESCTF/0WNEpa
emU0yyaqgrJSycmU7zbOpLK99zKCvXVywZYpXxyGHFeZyK8aKQYHcX2O4hT+KWeV
yu+vksTTo9sIAtoXShRGW0r0ZS+0pFoVnRcxGYsMipwncBbUKKDgQZ2v/fCVQecY
rAYuCeOaD0kk1QjiMBxIF9AR9lCBs1jmLfkEiQ+SK0D0lcXWmthDsMc+nr0tNVVP
VFzAkF0n729c7UQzvWdLn5nN8dpfbM5xFPY7q1I3MCGKRIdp5A8gE3XAhissC0A3
sNYTeh/Cc/4w1xGGRtbWF8lns5ZTzCe7TNe3QQvkL3zAdsc3s2qQq7HtSn/biJ39
wpT0LchZV9mHc9KPdvtEOZW2dRm8mP88txXDkUWolywyW7OHAgxltIJ7PvwA7yBO
6a9Bbzc4ft/4FZKREc8FHw55Mu6pA8pHrzFBLe6t3IbftLtvQtoiiSaVKxvSleIj
R7mSgMu99Fpe78WUD1eeR+e+9rLP5n5z8GggBY76w/QgzuITiTYGSW1watqELz4U
100AwGkdqIy1pUHXVOlpnk1W8qfnPhnQUOl18cHF4jv+XxkbBYCdaMcjZEcLBYcG
TfckdeYaXgCyXn9U+zkSvhATUT96HauyYHPOuO4W/Voe7Vabv3jY69OVeNm3arWq
F53nJ5its8loVqTITACo2Yl7gOVkzO+XHYxYUvYqmgT2aI69OCrNSsQx9GT3bM4J
QRkxELVkdcZa98oJ65xkfIgFl5kldQh/hhsVjeCOp6TkIztC4NSWM4ZMJMLt1aZ4
YmLlBwVrdzd1zenKKo5Uxqkx/uxW8TRmzUEqzssBg9BYZXTOaaLbSwwgfOMvYxMg
n0ZLvlQkLkLAGuItCRgh0SLk56vxqm/0pSocJdg7TAKp6HKojWDw4OlzyPkc7yBk
kCKLXxlpDVLYJfr4XAZBUessRBJ9/B5DvvrMtlIMWbD0UPVkLgUbAfGvl9E6R5PJ
apmei2HhXkhiXU79+NLr2HK8hQ2GR1jgMbbX5PlLBhewd92H3pOXu4XZfEy32LVs
8HsqI7rfls51RxGaO9bJ3xkrZuQJRaTuDGFlaP1Mk85O8vdY41y8aI4s6iCdKrBa
UrNqTAQiCdeRrIKWk5auSS//OKnyWcrwoHxe/GB36S8E/rwcpPATMA0I7+8jTfS4
25XTUxPAXEG0qGARny+cPq385X+tQlq0/qRoOW+Lska6YiiKj8RfWa2HBFp4nKEl
2BDd5GceIOryxS9NiBdnH63GPZEo5/oceUd7aS61ir/T3NEmt43vxgLkwcoN/aFU
Y8LaJsuCGYARLj5V0/q10u1+wsDKwAuvIA1kblzqGVQvIjt04p44WquiDzmiArzG
FyIIt34SHr42WrcD4copGRJV/sf9Gg8UrsyKXoS6Fi+VFcH5dTP9BGPNmEPPrKZO
xzjSTJ0Kp/Cu4nP0+4gkPswa9vIo8sREUudZ6lJquiPyJEwo1iOkOfgoVARy9zaI
agt/lbNoOoHlP5uHLRUZlLPHlVkROIVwGiCEjn/dmMk0+2iYgIHDi0a0LO9dR/fz
aCLWWj/3nj167r7lZd6v4/UT5+PU3k+3FPbv9BjboaFBlNm809aQkuZSi9OWSGhM
SnTmoybFKQfjtlBvVh2oIlE2Ry0z4rkyPaRPg2937pSa+dYq8W8uSZ6iRa48XXi0
LtlCAuvGIT/6ZScVk56cYJoW+4hE7a56zthqNMjQb6ZphaOejEq3KJepDZUf0R2T
cpxoD7Of41kRxvNnFAFbP31qYDg+7mx1Q3xjXirh1TV5GFXjzk87xraC3E7DixTV
jNOLglN/9He6f7CTxBiU76R04SOwundEDRpALBVDtrq1b71Nuy4wM3I5r85drS8p
Mz38wyQ8E2PmwgL53wiYL3NRsvbcSg+04AuCfFszePeZx4i4z+PpENn/mtEmi/Ve
3AXcVQVt+TCKCRJegWYGldg5CaDrqLhmhZx65b2P5I7Ey9wImU2vEW55QCbq0Nzw
AfxU2aqx4qhLriUqscWiQp/+6OG3WMLe2RyHuX+abapyAQ+Wxrf3cdcKnIBLBqPe
zVvHeAjC0cz2zDuxRqeunEGCPVks6wZOg6y4DFxbcam+jAlfB0o1aAyOA2oMbOw+
+cwzJCxFeZ+ZxIvfUM+6wAlU0sq7vwpB275Qc8mvzb3nW0sAn4/0Chf4s5Bmd0ze
F7GDnPlRtjoC/tVGoum3PF52uYPBs3ZzRb2QZ5aVrqJ5P813sPWxiPHoGQj5EIWC
qVAkbav+PEDHOjFZvzn6uBbYK62cs6+4KOK0BOFNRsUOfqk885kG/s0/yHla/eWg
iQVqxHb1AVCoWc5+evNy7pvcBNwhUQ3eofVPIO1WYKGIToALZcNnzujUPb9356rh
z8x01FnAiaR2VkOPn7Z4475A8RbtAwGzmG7De/tZkHfU679ooEUDZdJUQrloQuK4
35l/pmsOAWXdH8orciik1DrFwi6RnaKJbtLBzl6ZpJwiG7Cy3sFG0XJ8M2JrkL/p
UTh49COcJ89pC4KfIIUOmm6L9+tUHTiDiPnASxcDTgdSgUlWf9IJ+KkYiOzvLEx4
cSjrpn4gW/OBZFcmawcqMdZAwHsy20p8JcGA9NRX0GXi64OOc1CBUKhXXpvEP2WP
4xusqX0bK34H13x5IRcmlcFUFQuPjPKvqr/zAfDuGaSlkj91ZLkYVj3OHpEPGPQu
/JCfczACCdBNow+EqlKgvGONEcwzkCpIC4Xp004BeuXS+GB/6Vb+A0B5tem5LdxR
Q+1bcJHBixJpNNAr7vNnA84XXjAWVmXRcnyq1CrYNiz+CqZ35JXtVTTuHrZYeHoe
Vf0Ay3HT7P1rOjhQtQtjI6O3GumtwRd9/ly+Zvm9iGvHlUUUA7+ILKwTkwaTg/9r
C6I5FnkDka00t00/68xCTDBQUIyuyh1nFCHAU/jNv5v6fCzlFYX2CIBgj+anRtmF
TLDv0hjagl3v5RZ1BuP2Mj33/n/koxMRlc6hcY69RNvuuO1MGXnlKxJ7Q+ylJx7g
yogxKiQWmeE0wVlsku1/hlucXQOEvvMAoKQdHWDHODRfNhxJaUTbbeHwj5rrVeNu
jgSlNIpLt9YC1ybauczjjguM58t4/Rv4lmHapHD9X6HkqBtHISbTdfZaWcyBeSof
0ih2X/zyEIdXKWg+CIFmz2bC10fIEN/axx5SCFGGpROl2MA2etyEIAIW9OL5LK8e
icipIlSFw5nt/fc2HL/6BcpPWIDG1BNEK7hdvokCuW0UfjflfELp+zicw0he1Vg6
mC8SnLiK4X9zkzEohpQR4GrihHmh/WILZ3yAvfPwNVyOL1D8LkZpoZrEeq7BUyIR
p1QAKXeSzUuIPbgFNwO0mCr1CAwYPrT5mkHW5kxnymWdv6JmzWkjp+T9VKzwBijW
Y/RO5dsCs2TRI6eKicO4jXzmR1BnBOj0tlQjaJTFZpnh+4hCW6Z9FfDuLE5WRopE
XSECPnM/DGDd8pM2uDAhVjBwAafsC8q8zGlf7RPlT6qnzFkS6wWCWBfSKO2yLX8e
gW0JgUuVIDIqw3LjNX9ond6gDSLi/0fv3An/AUwe6zlGk2tzxNSLteNHJMOplgvN
VGHgP9Y0X7UhU8tXRK+wGFEbAu7ktJaEvQUp5ISMmwAoPzi7+7s8ylfbK/sZWpR+
vI7bM5W0Z2VBwWsr188oeWdMAMOJ4dKdas6Ut57TW2Sqf/pMksxuAipKLwaqomy0
mW50tKu7GpfRTiNnl7WRlMto+Pv4Mie/loyPIPYJV6Idn5WZm1iGqh8vkU5x9HHR
xNTZ2MuEtGb6/dlSexxMCuhK/d+C/ezlG9q5Vsbx1P5UM0i9zQxIsUd+IamKLNkz
C5ZO90+WukeDT4tp47IsDJ06/JtfFmi2Nta7T8QbwPo70iOvvrsxkc2j8pOu0k4t
qghGtttIW8ySv3RWWQAZboVjfXTY0rNMVpO8djAG2QV1idkfwbCUeDkW8PjJVJEB
HR1VXjlfLnsxd7gsOWXtfX1R45v16+t9uMrTdFOmOVFOqHRVkw1OGFba/Gd4NfvX
LyYVBnmd2OFh5zaHjU0hD/wW3iHxS7eVCh41LR3f6YfQ+KHQt2n+kUeqEJdbU3T3
oSHTJTBURl0zcR//qLWd8zQIST4SGY2aHHrndlYLPwc/KAf1fLyHprTP36eQJkF5
Gtt8KPGq1jrgOy3bmkCyLPu2D9Pr8wjopE6Ppw5++6K6gTQV6k5q1J/wlhjZBzeA
Kk/oEc2JnpBmT1bQ7PCuHmRbMdPidzSgk7UF6FRUrAduv3sFImweKE+KxKG3WqBD
3tCRIfscdHnuzXvGgKj7rQ==
`protect END_PROTECTED
