`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVZ4d9K7I29og3x1UPEDaiSUqg/aiBoMg9WyCxeA53ha86RNSRPdYJcAIHvo79Dy
QtrJfIM7cuGgx853JWHbYe3AWl5ezQr0zCziMXZPhYOgSFoPnHOfdx5kn3Ab3wkr
YFNvKopp4Bc+n2dJlYxMmrn+fUzR0+hcDITYTIhIdp1x8rJqsEKSGNeOdaCxhvdy
rFG95Pu0ZdP5p9Q+plWbMmIxsWckPN0YA4PRsfEAwrn8Bk+mwbAuiJ+Khs7y4pQn
if3abiLJGAV+HWVvhcm4iNPTjutp5Dp0BIOWUppr/5aXpsRs8FqagxGJbpye+q4R
JgHR8DeWRE3qlS6/myCpgv0snI+IBU+PLPKCvbWtykkG5sLIt3Jbyj7wz7/atuji
cMAjWEPUaQbokPNO4ShTrswQUAUbQ154vn3FqWaHeJNlmWyWq6oAL3+UvwqWDY99
`protect END_PROTECTED
