`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yHPkDD4GdNVjQP0Vnuyuax+3CAexbpn+74Kd2MNpQsPIVAWdGAUMIv6kkxzkeABZ
CsGzav5Llg/RJKLHnaPyY7tU6/j7g/SsdargRiNvhl7di3HL/xOyIaE6cBJTe8XL
8FY3rTe0yqrTQY66NLtZvcwSQ4jNh8g/SA+3TkoOkudsXTUSv2a4ezvtqkqXNltu
QC1NFaPhDdh70tmmc8KNOEonWTtZMdHOcrBRxMebfYPJ/IhPeedaqfPGoetyNQR1
1jYHkcrlY/JfTdu0n0BwemKvKf0jLF0YndW7luyTSe5JsoBDGH2WpRuy3UCEW4OT
7+u1Ot0dijLLSjXqmOYL7ye5A2GG4+iyBWS4h5IseLgVeYh/comYzRhkvVgqThwc
o5YGnyvrbSh2uWZr3aowGDpqaRUCrgEuU/ieNFFBEb5iYVis/oUesMfvZoFl1mV9
aPaMhMbp8tE4+j1KRMArVPft+3qZIJ+ezM2O1YGDk6YFyuE0wAS8MINmJzSInjcw
FJ7R1Bce9falkNF2HfuuvV5waBGMIBMqpI+pfO9O244YTsMV7W1Hjf/PVYIb2p+A
+QyUFpHUHX/IWlyMKeVHup59m9Dhw5/JgkTtKi0YMiznpLS0Hejs1CJBb2HKj2M+
PV+ERrIqNQza1atgUo/rfrKXdcIcwTngQ02LTeTvgrcONRLWkVPhnoh7AOxOYKuk
MdJb2iNtLIOkWrYtoaMGXj2A7cQ4ai33gHjE/UyJGo4SoFwQ37UDAWQmoM+2yuc8
cCiHCS8NTwswR4ERwbGwfuiJiGXgvt1NQlhqc4LG1/gL8wUYLfL8wafs2J9mpLjJ
UJZQkruEa8dKHhXzLd1VzssYdvRAz8Mpu44+iFL0pGxFVyhpwwqNJDfdLiqEdG5L
AHOfd4p6b2fgU9KwlrVvDllYEwRFdLlbCGpBLmdgwyUEyG+P2JLZ7SR3vsC1Se30
URiyytnVyvRYiHjMx6tvIo1SaZWOy2wEHLjQJ5ZK3vN+4mDQBceu3ieb8hXiF7i4
7vGZPCiAr2gXn0NQpe5ezGOaH3kJcrwGXSC2pWnz5yy2PtEQtqA0P/91Ph8/KFxi
tP+H2jiZ6rsMhGNq5RvSapINMbJ+uL8s9TD4zHYnKP8tp4ycQEY5OEzfMaFOvdPa
mAAyM/U0GEHl9Ejuv7X8e8S/iiCYojVia6M82BOJD9OJh0na4xy8GZLlUYcPC60r
wgrfh3s+opXD7vlsQpJUMhiLc0IJ5nWcAi/leDtbMMjffMBvE/fb5XH//anxR9CA
N8wOf3MniQILFeRIyyl3W/Z0ZTkleYdYZAjFf08WoVQDZyDj/N/W+v0EEte/4A0M
lGlIQlZS28nati/6aD2rF6gP4FdlWZe9rdcILrIpIf+N3GPgLp+2Xx5QoPJD4fgz
tssDvmXTPKt95HgvBdv7Yf0b6stftQBT9E6cN7aPWdOJ4qhUAw5z9VcVl91+9YC1
oK5LxUq7l4kaca3dJttVmiHO0t2o1bIiPGF6xOvNP0E9cquMcnDEc50wayqOOpJT
fBIKcoi1BV+zFly0ii/HN3V9HpheICsNr5c6oA2/KkM=
`protect END_PROTECTED
