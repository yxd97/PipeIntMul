`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P6RX6Zzhsy/62/E0dkESirf7lwizdtsDuPTMHbatybI+zOF63TKNnTPWR21xdsrS
zGHntRYoQ2ZnORND+nJyVBbv82g1BXJ4tNZVN5hqbMXjLtM7E5eUjfy06q5LtSlf
xZ5uH1Nz+zqklrPo1Cj3jQGTaVW2bBlUuSRSuCNJWgPwK+XsJbet0cNnQcTpbtf0
B81jUMQGsPHqQH9ulUN3/+WxcbJuaOwimNYnk+EtTqHLdH9Ae3uVuPladDHcfgUo
p+iKuXEYlEAYsSnnA3BsX5cOadmbiNvoUpUpw51sBlDSZAI+3jd8LY99Ci2xOhZ0
9O33fFjAee3KK2jPR++XH7q3qQPJ6a8oBKWYphVhOVvGRz2iE6FsvyYAps+LcANR
6/wf4VVfJyWD+oiviVDyyEHWKN4B+Zv3E2dTuKjxySWucJUsavURfWA5oEjkyD6P
tAn2EfAHsMH1WXhnoFBvF20wSBNQaYZkMvZos5GnPor6fcQmtzDcs0m9IdcQAJ4y
MgbrmTrfE2xsCAJuLSb4MfTsr8fJrfL9/M4hpaBX+5uO41tGMHF4/c9dxhFAya8a
qlLXlS6hYoitnq9cWHa0Yd+jpyTTRTsg0q7T0/5tUheDZcGBrMXKh0UuSgLKKZUR
gRKSZy82Tj8hT/zOieVFtQ==
`protect END_PROTECTED
