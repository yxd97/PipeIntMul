`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6D/byWyen80iC6UVT/aPdUwkCzWQZqf5btoYPCOxtDasZrUGLHwedDda4xpyHT5
01IeNdmCFWdUaJwuNUMv/lB8m83lytSYCJbahQc7RSXWSDNIA5xKe+W8RGBWxGLx
unVs17DjLqhnWFTn8ZIkJZup0grs2oVYv6GB5qL7/FBaZUItD/1IjXx67jnmXzbo
k8Gk0ovP1wNjSVoPTX9f3TWZ+QpH+li9qKP5uYGyVNczsCNw58JEdfLLYkHSwc6b
XlzXCXhNbGn733scVv0NolJfCJ4EP+l3lLTctdmD1B0X2RUIbJXwSvqMAlJA32yc
PdKDnguVcSCVVfyxr0s2KK/eZINUFhSXGfqQjGJ15b9yz2gB70uRfr3XgpRQP1Ib
PR0FXw0BasYxXxxN3hs+PG6vHWjdO3Q218ZfIKOPqJFfjPFtOw7bMUbB9WCXE1Oi
yZZKAD5d0CpcgLiUTmrljduwRKTXON34M6NCwfJYKgqQxRCyNDrTPFJaLY9Sqpbg
hcKalROIk66R3lENZtKIgmjEdjjvpOD7vUYwQtl4zVzK57w1+Ej4WSOLyO5BwxLz
gJa5cAE1LFnc8gOTY3WjkNW5dZWtYBtmrNwteSBp44Gn0FbBAg0BcsIACWBtaDPg
dT7u1aZ2BPckLe2GBdXAPNEKRDrNth+h2jnJ4o7+FE+Pdqq20L3dOApUhFjDZc9C
VqXCWUl1CAGORJXnf7+w90GV8ch6jwAsamUeUyJKb05/KDgOf6yptdGKL+xsf8pz
I1mgnyKad/QOm+FdI1bJSndthEt9+M6LNr6dfQheN/MbebOqJMMTc45jWR1jxluI
34XzV7csfF8yjYGdNJKeSikVaktnKAMJAK+OZzRd1Flblmv83JXQDOkqiP2W+pg0
JiM//548usfeFcF3SbZuRWKust4FE6C1SmuXNyRJ7zIWab1myt16fT/gVgXhVgj0
m87TTQLaVaAm6zK24azjZiCtXtms/vGaWMKePGPJ9jyhcJAE8NGvosdGsiWlR3xi
D1UoibDs/4m/05LgtgkGioPSQL/Wu/ytGV0R6r6Z7VcAahvNrvrKND56u07NeEYA
6142LlVlkCyvUoWe/xLT7dIXGD9pL+kkzzFmvfg+bXFVVud67WiwDRtDxLOOVfze
3B++vc8GjRWE4qPmI5FeSGTkqk+U2o7E0ugn2CCmG48MeFb8k5WVQwKW/sg7Gyeg
g/4ppNNAw5RRlxxpLp0BBBONW6c2+b0I8AQweL552saBA2bp4tK+ho/U1UhSyzSS
JXamyvxRN+0EqWEkO11eSU4/NfVehjquyvg1BUsaXSbQ/ggZH7jmLyedwvO0ymFy
OUrcNSyYF6llmOQAuinL3Q4Apr7bdeQitctAVrY2blnqQ4KbFEu9nsA9O0z+3E3N
RaaszE2cFD/eal5bhKj3QZB5JXWeYB6zOIBw59uEi/HznfBeKUH7ZBKjAsOHVJPE
s2wr0dM1FQ2yXvyova+X4ZM5B/+Uz2+Ya5FHZhffbR7oJsg4TnDdBs2DX2Twg/ZC
9m5ClzYYFuqczKIsy8+c55jE6vlmTQySPqcMsY7Rf+uzPtzXAEJtwp+SYYexA8B1
bBCmkT+2xldXTSamisRH7nbdP7u95KPO2d9GAvlqdphMZcwXkNqIGmr/KIECuVyS
VwkJz4sFcszs57A9Z/Ze2cu9C2Forc4art6KJAw+gAHgjPd/lbX3vYKezNvGpTz7
zAlyzbfuJcqfLm6N9m77gcQaKCYKpm2wcivGLnWVVciBlCeGu7zmDCOxaPKx8/gO
EKKsP1lAHS4T9XhCwF7foCtkflbcHpEfQE/CqsHC7AZpC27glRG6qNs4ZnhbLdTV
BF4gQj0+7fnUJpwTJECMJbLUe2UQWvoHPxprUEflqO6GEefwd7TQ4Qdd4UObn+HZ
CA6Dcp8pdn5NtbKuZ6ZqNysBY02XPX2BxG1+2ajJSY0nMUrnlUFQ/kf7XW/xAf6G
DxOSo3fXnbgnGlfezpQW3aBmNxuqAjbqaiMxi7J2qoVRanEZjP3P4s6KOga8eAtH
z3wLnzZo3S/tYzahQ000lV4ADBxzDyHUHKh9ZCqv8dWnuebeR84a5gjvf6Yuh5tR
t1h6y3BvdVRoGeJ2JdcyaZ3ySHSpKRYVfcWTiyAzI5iTr10IemUDlNadT1GlDm05
qq3qTCwNosj95t3jjGjF1YkUD56kLKmWB9V1wzfRFfOntVMHMQFuIGfXjVPQp+yB
SeQWBf8cUc/GOCFWz6C3vaZRlp3sX2qo5oDZCf3eUGW1/XvIkomax6OTbuTZT3Aa
XkHAeQBywqK7i7P90K+AO7KX3Ur5YyzlOqQcipNR73YHgJ2u9PUX0IruzlYMoiP6
I8wN2CLQLlfXc1pOPRtkMVKkdec4/43/wJPt05Z+r4vD1q2qarpCotrU0UhHurZ0
ep8iHAdkIKwca/pADfvnyk+KVsy5IZ6IoIMxYICfvm//32vRXaUiPRWwoKHwIQNd
bFaHoLeXFULfbq9rearf/mtGXxasLQMOTGjPB3DpWtleb27WUqMag8G1dXpd8LrS
Rut/6gSKGlaGChRuofdwhXkT/mK2XnlR2z5Sh/pl2IGrjDB1e6ecCAp6JxriYWRy
KpqZepMI5vL7QjOwPar9yQ89oPV0jZkeI7dLdFZj6Oxj8fF2hDynEMDCktPkCQ5G
yENGWHoSwiNvI/T7mqC/0tpwq7TlAxdPTkbH1V/ah9V/0LLCMUCouRuLFEbkihFa
iHBJjY9hZBaEIWzyaIM2MYq7pZHKjnIY62sBGfz7FVQo1Tnu/CgjHY+cg1Axd0LQ
ZIVHuFUepi3bnkMwKJ+Hn/nf6xxqciNPR7pzzmCkFKl+fw+9Tct6rYR+QlNbsAcm
jwXz2QdOQL8jodohnZTF6scbSPAhVUNqNqs6W3qVWRz6+alp+hiQBalKHvNtDv58
tADF5dtwlld9XyQg+j4fqZqb1SGefF4x37kvNrHHCAmBZ7Q4zV2bZFl49kIE0TGx
HCfO86+G9rgh6ZgurEn0e+0rD69U5uYmb85XUd2dgwGTKZ9ad6+6JYnXVly2qTIi
EGeasjeNw+HQYcwTdaUnXEMXXUfqoxXibI8kHchkbJ+dvDYKCSWdScN3f9xBVuqK
YlR5c+NmL3QRce+Hgq83VoN9S7zGeyquz9sUOP4rEcdOiNRnmgtdDqMKNBEcfg4a
uoTmGfO1HHLOTCrsz8inYYwdc0zAvG4FT5DXI00RffvUM/eTtOmkkOnTM+Ec3tJ8
Xu39dHTkthPTLULssbkix68hghPGYJMUUzu7lPh92D5jg6xoqNY2mAjlCltlDm06
OPoWKpCvDlgKTc4THhaVHjMyWkB8obCiLHq1GwhbjFFVlnjXFweiVKkGFfVGdo9z
g+jUE1n0xklBYU7wmMvVpaBfJodqjZJdsLnoyxjZoXtxP66k2RP8H5j0Gf500NXN
UK3EiWG+xRDEWxkCv0PP17HDUq3JMD6DrbuRugeNs4lQ6sPFQawO0T0QOJZnQI8O
6zMS8s/cVdIKuiXu/aoxx02IVCb5S1xhhzwx6IGu3ZRiBpteUB0EDBaVyg8k6Dk3
1uovsPOJMkIqqJwdVJBfFSDowMosmoh1QGlh4pNC5RzMw9x5QV/3vQg/7XRVi9YB
WWolr2Y4shH/AVfIcFL5Ce+MdMMHJosjLeKPj5PTfwN31IL/kANIgI0Wpf/6LK6o
jscYCk17+7cCgxwJGMCzOUDHC9AsN4tgvrz2vG67dokg3HkiTsDa+jsN7+BUQsBR
4oxLDWMYjzbO2H667Av3wcQJxWyY/X/WcDhf8wwim93xR/CaEyU3+x/o/FIih4VN
`protect END_PROTECTED
