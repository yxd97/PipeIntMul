`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FdhunOb++Vqg+X1wJY6HUirsyuNubXlpeVmQseGUMfAY8phj4ZKW8tc/33RcV98D
gPz1Z5fYbD4tQHX2kgAUePK3gVBtoj7eJ75UlGMtnhr1VXXTaC/s3OIsQjoKBeko
dNvJIEEdv90Swu1qAgk+9mmu/7kIj2dw8W4TOrGNrf65VH6U0eoQ+kIuHhrSFCS7
kuxiHlgR7BQU9FuUhnyIPiQfuPhXye46EjWsQf3KE+3On8DCigY6LIImf/ZwW/Gs
Y2B0B3UzCTjojl6RujqmsvZSe3yX9WIKKa1NMzY02oWQnXYc39hOyMzPl5wdmsM/
2li7LXmF2jaLH5kh56X503ed/gCAanuHLdrJFGjy2c3F16MAg7z2i3Xa3IkmIs5n
`protect END_PROTECTED
