`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aHj8OrYWhtCPYZQb1Y+YYGDcPUUlD7TrmCN8AvbkIUwwX6vXiXhQxRG4GW2hnrtF
tvQss0d0PCyKnR55gZHkmukhF99Y9/bSBL67EYoe4/6WqOT4t7/VLzYZd6zd6Xu4
5yGG6MJhxYoculAR27Mqfsu8eGCoyL+khARshXDScvKXTJFSrVtToS1lLLPJCx1+
u8Zqfb28BlQuL/hDLaSmSbLzjr/fsxcX53x4OLGjJUdw/aJ1oDO6jBxCIEbTjJUh
3Myw7WiMovKoMj6cTfMCe4a3MEIIGpSPtAswV8uoV0q/DPqfqnOJkUOU8agF5SSx
aD29M13RtgyQvkjYLRQ/08R8j/gcXMF5f6wby+LCyz/Ssw3AFOxSAFqWa0JicNLV
XPo1WdeBJrSnoam4EjKu2+nz/WdkDDD7hjOJvS13jOXsXvxF8JZQk2OAH5vQbl9X
ZDgLDRf/7bGcJ7dQNQ9ozw==
`protect END_PROTECTED
