`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1qr2gzCrkEwzZBFxlz7jfcvQweLC5Rs0OpRko+XpS9LOmjtU/novqWeLNZiVbnGZ
aCKl1hCEy9r2fs8Q+cqbanxVrN2CWsOoHTzOQTAnnrJjvz/u7sNZNBEZF4xKdWmt
2makcuGrTMfbf/+Pr+YHHkGsfPGMdHanINYWEVf+8/twV2RT50rXQLKTbqYwhLdm
tb/Lx3dQL3YO8jnfY3vgCHqjQQN+LQsN3V7/K46Y1geqaVfE3UMGAHlaHt3TxrGk
wF9haF6+dkIFmVosdqFxHt2gGa7Xw8ON6sAxjvfE+yI4SHm9fZKoL/zZlZtT1xQw
6QwRaiYmSGNNg9letxBlv32pg7esqfzCIZ2VlIUQNCxQ5WtlQ2xR1AG8MvcV9rZ5
7mAcqgTi2eS5c3ScFyppq8NcIeomMAf6egA+iOMbZvepaqyhHeCDIyr5jx9Xmrir
jgMng5Tt85tx4I6T8EkF8uhLKLR+kpCD0Ll0/izx0Quv+1Pw2PXfcELIC/K1Mia5
gt7Hs2Kof7O4ISpg7QzTs5aGKmZdDWtikTWdIjc8ePCr4rrYyKZyZ4yzTwowl614
IMPSjmkSGtVA3YsHz1traws0+oZcN2UFym7idYQc6P4hQ5dczcx1k5dWLW/+9Roe
IWa5QYlTSANNI7dtxYQOHVOHLucdyfkOTFjWr+JUxieeQ+9RQdwGqvuu70o5mU70
rJgqpZ97jWJpU5JK5SF/X1x0naf022a7juF3dZLe7jdIzAzVKhk3JLC1sFDNrLV7
jf2EGLPrI4FaKsB6kaHXqinDobACwlnCThAW6QpqG+uDZ4tHmyudmH8bMiy7ntc9
5xnFl416mZHvrlCN6IYKkbHeXDONsLjBBY3NHGxzb78vBQBmZaNfLELv2+czNaB+
oGNANX69wXmtCYdy6L05ngJTQA9BBjo+mfGeU2pjX6aDlsaIi0gZmNDsyh+zROMA
/NTIOu/FzzYwUqhi9qYfWUlazyQN6tKpsncXitVMeVPP/G4zsa3c5c45bZ+pCxry
uv2Nmu63qgJCBnHTryGj7gvLHIdDejhBGQyr4GV5A/8YbrxBsynsR3egHRShvwEq
k87p/ZrVi2X3q4r7GTSsF2YdH8rJZd2heGy3KmOaEj4Yp7WaOz0cQl0rgidiSxk8
Vd7bDwUeQ2MqcpDTOnIUQMAMQu4hbQ4o9g+B5ADQprya4+rCFe/fRYWSw477lgfd
v3giDVDL+4/JypZuqUQIBm3weshEOWvidWruq0YrEEb6CrbxxlV483rXR4uhCzef
g8AlP21tb5Lhtz2Q+EIZdpwhEyNaocdL05r1P2QoCa2F29B2tKy6vaB4RSy6FZt3
bV14rcMv7M7vY+alqWWMo7BLnHBwDoSo+blA38sW+wGOin2koVJ8hwpC5pm9Op3k
LBvJYnw00+eN4e92UjuxX8wsWPVnTiQgSud77pIUvKlHgzmmLz6lZNThfFX6DMqX
b9RO0V8RoP2N0BfqW8eqNnMnsThWqIzcJ8JIamnTlZ//sVRr9AaDFdMo9hK/U8fb
OzXP2LsJYw/P6NQwMzBwOMuZ18alhxzEoLs2PAPWkBrT7hRG1+248H3Kl7ijQPOp
xE1PZefl7I+FGMMeptCFAcwGRRLI8fVqNkfgzTNFhQoxZ4ptgWqvHFwtvBed863X
8byyOpyDaVk3/IAuqFxTxqi7hnIpshOZg4QEX5QmL5taTc1gR/QpIjOE+3xESObG
VNg/ny/Td+R34V1QcVlmhNC3LXrNuXpd6ekQfvQHkRyLRMXrJeQoflSLX4qJx7h4
kLxm4ug4DagC+M+WvpFAdj3TaR4lv0t4QA5+wqQ0NwoAlVewzepy64Xl17PLm4zA
`protect END_PROTECTED
