`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTm+5m/NHDckm1fTFW+9YlTXy6OR545lrUFR/TMr3tc9CrVzpkbxKXGRiIIWeoWP
u0LK+JTj62ewMoGNn0rxRyTvbGWfnJEkhM/wJYlRJzLwOE3Yd9duXKNU2Csrrdv+
U0vAEgTqQlfEOk0Sk7DMMsPpRJ2sJU39cQKEZE1/ewfd2CFJre3AuDE0/00+nWe0
3UHiGRDejYo6gMe0AyjJqsTj/fzQ086WRa9RYPPnKa0zaRazPEdMHdujA7ive5f5
9NfkCpPD4lireJTwyjyrrXxIDkcdhJEH2G6uDGAn7y4ZSX+dET3IKsSDQlLz/AyY
wdLD3G0n2VzL+8SHz43T+MRO/Sza6I/l7qwl7HUQ+4bxXYgTR9o4pz82rLomjmKK
fDaskTw8IruvIL9u3fxWvCvnsZTnXJueOzbSdzClK43nWH8xMC0s0UHMcerNLoaI
zc3U+rXwU43w36vXFMYt9aupPqjKBxKReNb0iG8y/BkMPoiSs1ITZUjl4drSyfyC
Z4ckTRroIaoIHtvh3RrZrTZVEwv5mQ7kd9OETXMAt56wOBPghVVzkYmedfmeVf9Y
`protect END_PROTECTED
