`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ftZOdKj59HqNyGhTc3qwoDuVawZk+0H9wRDilUNqyiWPWmmgmpQoaw3cJqkNxsGi
mAJ5gVJwm6atWa+RQaXYRtum7s/iBiH+VqPVcbuEB6uLDR+k7XDcvRBRIt/MkZXe
+I7C61ItLFVxfnvzECTU5BU/x1fRya84B3uPJSx7EHZL4RbANHwyRTbbemHuYqct
gJPYr8Vb1fezRr9/odnU2378pZ2Wb1ZpTfwDA99o83wvVksuXt15Zq7zoinOtcxl
Sp8oOpJg2ZsrTdvuZjZ8rVt+vFVX6RMv++LPwZSFB9r+ElavI72x7NonSGL8Fsn+
1rIJrKqNIpbxkkxPDCHk6pvMZWlaYAIBfHgyTF5THT7erZ05yWBfh1KEcbAZo+B+
khFPIdddtpkDPjvK9fSnPQ==
`protect END_PROTECTED
