`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OYVPCsvRl4ixOVrEVNeqryN9jHxKKTsMtYJnVE6fYalloqWdg1oaxq7pHJwvG5oh
2UiAYFt4LKqOkfhk2vbG8qCWFzjWjx7FivW/fyOHd9nvU7ErktrHHuTdgKqHe2tS
5IegwJafkLnX1qvbqHFgMSFqjCbTy20QgGW901YjmGaRk2b4Tiioqdi2ErGV55ZH
PZ2YyuQKd7wC/W83y5acLotPBprtoiM4CDdtyUUvLdmK8pZsZj11HaPPFupicNLh
nKbb3m+VMvqe4ChE/oD/9oYsl2a887Z804bX3Oqmd2hhZL+/h0SB5mGgA/r4xbXL
g71HOEcYzFwtnYi8gl8444P/tQEKAkv90y1WzlKGS4Nr6tqWB2pFNF6YmnVUYrLE
KHbnlzdoY8u2mJ0g0FGgykLGdVz7L9ebj1gfpIAjn6sCcoML/jgPeMyRN5u6QZ0a
xHyPLupiCM+klTIc4K6eSgNE/8X3KKV4lzel5jKK4/zLwSlCXK6udt6l00/pdw5d
ZzeSN1qB4QW0evkd9Ni9lXu66cGYa7TFlEUDY2gG7N37kHG47tDEEuwYUlFyF+p4
EqHBg6REjr3Isu+nGRPoRouMYT+sghai3qyOhnCIjfk/VUmxhNthIeay/vMnl795
mCVNc5VI12POrOnoM8UgSR0ffmyI6hDYRsXaCdRFKekZc6Nlg+tIwskfL1V4cxS0
OL9B9gyGo8QXzTRhRx64Mp3/0GYjT4ZDan3VptR9hV52Jrc+NTUlbmpJbH9yTSJj
91YfmP57a0dIb9GLox6lBZrwAn5/oJirMgh0nCJYEMQsTAaKRcvglXoNn1z6T/+v
v9I8EqUhicQ/YJs1YGyVE1ARkhSnoubTBkdj95DMmqd3UGwr3/2F6w4Gks67IU7I
F6gQ0CreD8Fzh6kDEl+N2+J/Xo6spZZUhN+q5NxJApOJKJ/H16xLiX47kUPiiOAO
w81WB34t+wgwBD2qFwGvXxRSpndyO1hB5Wl7vCZ9F5ek5FKx2J5sFXdZVStv8GQr
ec0HNJLvTKzUzuBAvrFN2JijLhQYWgcApdc5nAOiQfTnVuSsswB6/Eeo1I/uJX9P
z+3s4xNSeLZSuzrf9SR4y7CrEZ3WRxXyWfIXFe68Wc1mIAcVcLYL4RXJTlTWYjHj
p5nTwzy+yQxmVGSP+GXihf6FZaROXyxNlcVJQ4p067VbNAKbFE1O3niQqOHL9/bD
5r98T8r23dFRnD7SLS9ohHJOZplAgtm8iZ1/acRw8py9SSe+Nqki77KB9+H2MCfB
0OSH43c0DJm5hRD+YZvAJemXUEoR7jxh+XrRpodQEBzv/4rYyVn2WfH2hCkrDLvI
fickbadHuwSKNLdI1vpd7T6AqOxaZKXdnJm3SQdxrUU0PWoUEPbV2k6Q9D75p9fU
lSje4ozLP+1j1tZwzOMRajBLod33lt9or84sTSmCV1ATH9Ju/p/4dgc6tChmR/nA
OqgxcLqlKSaRrqyPK80unhecdWGS4fZvcBT8S2uvPmCjobkARc8WE1moxVXo40NZ
fNESCj+GWUB5zaSyfR3dcA==
`protect END_PROTECTED
