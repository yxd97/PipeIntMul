`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4JJHfVLkwDrba42DXHHN6MJmQjmWRnTSWnwxXWlcNA9FLihubq9wQ5eNnxqoAf3k
9tQq5H28NhPDQSvkP53dJzXLDAuP88dzYARxIDnivYCQqe4tQr1qRPSMd21BAeS2
LPaEvWpMUt4mJt/6wU6Kcv8HzQihaK5wLbG226q3PgQQ7XYgLePLLLT+s0rFCGTk
G7XH6lZ3QzAhNtsiHv3aGlkVivN+xFjuFg65UuNGLfWG++iDUgB2GJRH6VlzJncj
QGXsGKrLjkWqviOmcHzfG7L8v8Kvip1oz4FptyG3Ld1djD/hMEUbMAKX63ysfvRg
E5Ye400okrwVVYszBSzEhe4cCVaT+s6E6udKCBwp62kvEXeI6L2p154i7X7AedXP
mYEAfJ9S/vTt5DJm6l8/rfOGJONb7Ea7p6EGP/G5NiTrMHyzyqN7pi8fZ2JEEIYk
quyk6Psu79ZL7osmpmqeWDfZsVKS0qeCickMGUr3xe6tOMW63C5xWmhn41G+GX0A
EwMHXupR48LZb9oXSinzT/969qw5KvDTGpkWdCgKMl87pYZwSdw/iUq+Hkjbr0EW
nNQIxDDEmIkhUdu5J50pRqyZLiJR5pLHTcZgNgOL1mZS2UYcvWV3LhHyc1O15OVm
zzshkbhY16fpITxWfBF9ZIN3N8npRZSepqYPV9DR2W5y5biAuFtgs9HW6SkGXekx
Wa+KKVYM+o24qD4TnXX+Hl4mDmfEtAOkr5Iy5gxn7KbNOepYe+eDSJ0zswJitZkP
zAWlJLq/ZrKGwAZtGhF+mZhNG2ujt1QsFg6ev5lr9yo4T+f5JSgdxppPLFEkUOSc
QzgG9CBJ67JKNGazyGgFCfd865TYz01M73KQacGSU8PfGInVBcPJhNHFmhZ1uwLV
ReAjba+VQp3XOfLTkPff2ivKaeeRR5HsW4yibrlZmZsd6m9ubS3Vuie27OMFnW8E
LAcHI/bjAomrESZu39SBpVAPuajrbc20vszyDwWxM7Mhuql+QaUZMqU6g01CpcqS
6Ro1sBfGuD/LHsR8vUFLNrtmdcqFoyEC7UhZI16sdve0MRUkpcor7tOy4Tfak+py
c/hU9EMjt4XTzV3nmvDjPdZkvBPx1wuORP6siDeEIZ1LbmhmzRUYcMTW2i1L0+GF
cvqh2N4ND3XajOM2ssYuS9z3XPwBVxC3r7Ar3e2vkYa91aV25sLkyDveKvA1hThz
Lyaw/vWmKCZpPJOa3HX7aoqmO4wGGd6ePb7GZuoGVlfbIr4o/8Bysyid9ktYgTr+
qD0QUDwKBSxrva7VfpTwLi6Umy+ywnjjrn5WX43H0Hcizk+zcmIOOJTbOwwuIG15
p9ts0+sDKHQK46U5OU+vtiwVYS6bvw1uTaCj7wOIPXPsHvOxXcoyUIgiNiOkiRH4
wSVoKjUPFPejy2Wf54JPkPSkxTL0xEMzKcNSgkT4ka1vSgWKwRuuf+lDeTt8744+
PDp7Toa+oyG/FOVIRJNOaAk+hdPl0cg5rWdsI/XovXj4EkgkSnnKiKk5qo0KY2Sh
lFjQFt9vYjqrkt7g9ld6tQ==
`protect END_PROTECTED
