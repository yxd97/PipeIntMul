`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cVkNnGhHrqpCevc79JnX3W7fzk/rcyEpyiJAGfynGqNA4q9tE6LxSXwV8gZdpfUJ
aeYHzBRx5+JtUDK3+NCDJR34c4ViXfVbUSK8qP2/i2ZYVwyv2ZIUvjjcm+5BMNfl
9d49HZsfLV5eosLeAMjY5vLk+KtWMn1OsVZiekBRUtOyVTRhqd8/YQC3yJ7/ahgA
nP3JHfAUYpxNBepyaeo3qDeQzxsvAyRJj0PpXcsfEmld5sMWL23UMMH75MhYOu6X
B47OkZS9pDyLrXLk/2pcE/nNDzfnehHfLXPJXNOqw7dF4oeeY9A7V/2kKVxfYJKG
fQAWAJ3AatB+xkpyzY80gBS1SNGWYliK4z1HffnHlvww+NcUxfeJupEQ97QvxDg+
6lHRVw6zKolFoKkULvr03bmZnb6PEtLLftTf4GR4XjlNl1hkWwEnQRKwolFidBTh
FXRrkh73fIkI9L7hQyABjhDTMF8YWFl276z5Tioq2NkVAi02AP0eXutEd6vA6AOb
`protect END_PROTECTED
