`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fkO0my5z0dGhA+g99eKik8kC/K449Gy+Sj2jiz4vLl/AChrcf1USqHrRiFD48t9P
QMzgk1iNr2oFzXgeuH1Giveu7kWcS/aTTr8/PNeTuxZ9yQwO7gV2yerxWJRvEzBj
BPQOlj/fM5mZgNSq7pOzBeWgfjRj24lKoaxcWGYE9loktoBqKzrykGMWe5wLEzMW
igy2UPlCQOcN1g+CJt5rJOGziCqzoWdx2m7WC8Bzjf/DIcIa8GQYstZ9ZriJq2XK
9tvY1mlef+YlVTH88+ROMt/6uD5rqmZAStomoThlpQcc8xUttCy+6P3TOFAvrRcH
BvrI9l1Anu+cfWLM/RiUEuaLmTsA/uXgC0abp+h1teZ35UuW19VuDUP8XnswIJm2
oSuwi/Oaxe2JWTqTha/nKzCRK3ncWLbL159+KZnzllc41qSLKOa8DHECpnfSHsaY
`protect END_PROTECTED
