`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9ZHXbGQzuV4fCIyfOY+41GJyqpt5Ik3+DeFZcrPYZ/o03fajNTo+HripWPmncgvc
4dh3XtgKEAY2q7aiGhhq6O3PJEfxTLLj4jpNrH3T/VYS0tIDEnmk3sOETseGpZ0T
owEkTIbZVnYdrXJ6KD002OpnSLfvJdOIpyBukVxrxvFEm3HQF257JLyOydLTrH8T
rXJkSAP4yIDYVAv828Zr58ZqNH6IbVaFsDcYL82c2X9V0xMia+pOX2RXR1us8oTz
sW74J8ugDmwMoC8d1Ky/RqfhTrqFQI9R0TLoKhcOxLCrvvbHFwRpdyX71ZINny0v
6tR/gwuZ8dTo9gtBFWP5g4wDBAXXPa0fb12WSNKo1p8=
`protect END_PROTECTED
