`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5MfuOPot5nZ5Evnrd4unsom2geUfN9v5vgGMcDAcX64n1BllhOl1139nei/q1JEj
hnjYkZaAnzeKrRF6AEPraXVHlboLDFoiok3oKgF/fdK3ksHPPFB5aq7toizd3rNN
1+wOw6SVL9aw1qAwhYbkBIuCFOtNKS167JK2mM7LswyjFUVGIgOKA3GaJqzVQPqy
j+O+veSAXBAb/nkQbVc1dupVMPuwm6Go81SGCjDMhpoyom5WO46ZIbR+01L6pF4F
bE8hdtE2+HaStRmva+D46qudt6Kn2Quzj8ElLZTabXMZMNHkyR4kAiGLf2Xjz1d5
rId2lqriZ/hLcAGfB6i8yze+dffXj1Fqvq6NHzlG3CbxD44WeOwE2JDXbBVIIUU7
m0hgmq7kbuYqONYSWlmbplSNYA7VB7SjEYKNrUpEPbzyZ87bI81IHXHfQi43cmSC
UeIMYuftwGxmiERRKtlOYu198nVozIPA5MwaydtQzvAWbPIA3z8ptAV6I79UteEo
jJYLu2ojhK7p2Lz1pcZW5MSTFZ90UNWdT8SXuWNdAQVCGyl/YDgBnFewo446yKe4
KQ5fH5daAuBZiLmFVbk/s6Ku2tqXmYJsbwK8nJZZM16u3+xFPJ90lVP+QoTg+KyR
AOjGi28kQ5wg+Lts0LmHUN5k6mqaxKCq/MEbphNqxAE/m1sIZkOE5+2q3zU6RyxS
vwgjg10hFG2/Inuc2XVQ0vive/IWKc2ONR0K46J+iY/Y87Lf595TTjj93BHKnzws
06ThQgx7gMHltjpu9ytzoB4H5zVhF5np7TvuU+ZEB9RdUz8/Ab0S6zVy7GaROUCc
A7b2TUorM873vxyKTPyN02YWCFpqHFuQjDetRb002WwrHoj7al0gEf8NrZ9hDa1J
vn3qhvqaB1CjOb/62eHrZ/iHUERGn5hqAq/WzBmJaAd7cd6kFRe4xprcBN3jtejb
7/CxSQ6o0QQNGWfCM3u6SSaUfciixQ0bz5jmor/4EwOX7zUdHGM/4bWAt07t2fiF
16rGEkD7+J4CJcBSZFo/qQ==
`protect END_PROTECTED
