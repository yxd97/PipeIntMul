`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hD/kXw8aMiIC35KMo6Or09oAHs8FoS91WxYPVeqsoVjx/EYs+yyO2eFeL+vy1kh0
IqoD/FjOyt0t8Tz9LWwbBJb4UsWxyi0jVo+cAzleCUS3hJF0nEyw/RE0fXWdwHAb
6Lnh5Fzz39yGb4hADZSGYco/yuKXRTcqKxpZGhiNL1igYquFGIEVH5ywOTNuRetp
h3Khw5rykSNYQgRQ0hlEzfGYX3RcG7aP5ILIYhJICmT3fsZT0ShWhl80enMJUQWi
pFRBrzJPKNo4284cwV8Qyx3VQHzvtc6FwTYP2gDezJhTcf/Xl2imIAwOBktjyShq
`protect END_PROTECTED
