`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qrvfAXWJrr1sxRIO1Zf+5dm/b2ecKkgG8mBzkft9R9E9iOgFAoAzZv8sy3UV9Tz4
rrMZUgQBnMTo7r8aaBaJKYLb3DTBUpuwW++rwlVwC/VU2u70KjktjEfKghzBrXgT
pJrBB/MhSwSLQOJYFcpUDY7LlddpLTG5JaTxfkJ+VD0R+YzJq4JCegbtIbnXeoPv
PKsP+IBdp+LqCVS5QFyqvuJ/kzXvg38uvWyq/sNCHH493x+hvUkaGkK4i46Opcqn
wihpZb7SqbyuCV2PcCN050CSRpm/gczZJKWAWBeHoP551d/Sifc+zFObK8yQpdIl
NgJePLRYGvjjMgFQL6FUbtv3IGFzJ4+ih3ri4bbS1PQ/4MpLooaOasMQyhTwDaDx
p43FTy0jT8ENFgBLZuqUtJLSRdizrkv7Z9fgxWG3vgtSUcmxSl06ZvTg/2IN3Djb
GERsLcKEzdeO5w+CiEVq0tWrrG7D64XIrNDBMhxhvJOUH6NkmilujiO024RpLziX
nSPNY5uwMuXHfJMG4cJ0OlZbitJXagJrLh8sI3GeefYGb6elRHVpovuG877Hw0Ol
CPCy3qXrlhF5A59E8TLuBjid3EdqnDD7l7WNUeBvIeuFiNdnAOq81yaDF9AvWTMp
gZJNxbffMlUMPGceXRLBtpcYLf1n5dafqtsbrstnoCAyxtsQqdMxzZ5r+BWDh68i
NbfUh8dSlxy/OZ+TxOEx94maIxT3u3zTkKU2ckZmTH31Gxn10ZOjVoHMxVamUZBP
xfRllpvjU4NyU1AX4FJQ2nrWQXRX16an17HJxeliXDrzZUY9/uReU8Ktl6/7CLoW
8OYJDsgp/zDIp4NwZdaVhg==
`protect END_PROTECTED
