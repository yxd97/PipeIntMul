`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
InmjFSxkm27xE60j0x+TLYqqZutTQiualDMPhe7X2r3vFK1m7ufYG4SklzeKBhoj
ZNI6kkyHSxPkpltpP/hxpiRliGgOhtm51v5IkHuiSbbSX39cIVOMAnVkyK6SJ0hb
1KKs7NryK0iePJQrUq51rVWp1TIZ3z1ElUDEaooGrwA9BE8hv+P+qprZHDnFeHQV
1oJ09NVwliofXCX7LMcSqVDa3gtxWYoqYUbP0TDHJyusPgNbBhUnOgYrJ+0TmIz7
+oB/Ap0Bk00tetCZ1D+qjOU8q42aN//5Z6X3UFy0vx+0Yg4xJGG0zJ2P27Keh3XV
oeqfl5bXmcArtDbxH2ew/A+L+js2cKgqyUHr1a6lHOfFXBO0Om7gXizHIoa26FfD
iFoJLU/kyH47z/F3VSCjxXAeN+dUt9i9rrqby6RQqhZl+TkPd7UyGfFwbsOmFWFv
`protect END_PROTECTED
