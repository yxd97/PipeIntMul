`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NZ0MkuM9bw9G/GaCZSRebjbWwtZSxZNtNUmdHI15SeSplpNnzR6Mtujkzk54YdLc
TeLm1IZzF3KFL+OgE9s473AKqoqfJrlNpSw2TpF/VvVevJk6veiVuZgJMsveF9FN
mSCoXZzj9IfRYypkNg+r6RtZkCFsCEACWUgmbIvazPjc2/I/RgFb41+GJurFrDxw
JalBmk/YqS/wG59A7J7vOuh3eiHIFQm48j6weEoyP1/Ol3xeJB6QkGhNm2AOTOtT
l9QU2JHUHsTcRGi7bqDr8xZDXnG6t3uIyPD+gvVGr2fbd+MTz0+8mBeLx9PCoTIv
7M2L2dpfsOmvsK5t74ySzFmAzLROGWJ1ndHyL5DhMtB/MTyKPq/AZLFmt27hUZD8
lFwr9BGzWuoDJAftPh/2SchvDdV3SX1SknrLdC9G2xfe98ExWI5Cp1U2t1GJFZ5s
iYczROyVdZggAdb0RLCSSIDquieCS4KHNifnjBCG3DYi5ccgboTDsbtcebmPFOtE
PNWh3kJW/tMFIk6+ILgHxvTtG+gXv7OusyGuL9UqO8AN7b7hePJ69T0vHsfOtr7v
xpvEnZPKvfqO0xBm48DknIkYYdFxIzFDM8uflJFd2RCFqkNoNTzg/eN5HJb7lhud
Z1DyJtDADstpNEhj5YxYAVQKhwbUB2kcdlYKzjm8Cdr9r9EMktMPwAPJmLPWDBwF
4g6TvAeG/ngzuAEqAU8+SJzVvhYHA4pbgJFlGIsjLrqJ24IQu1osjW6pRb0bD7oL
tTYZLMP8iSoyRGCOnFm0/eJMqbwSqRxGFiGufYNaue2umQjYJmu82yuzTePF43T1
zRVOriStzSSMGtU0chDSSJtsB55Tq5eunggYlBrfAoon8bjmm12XNfKjPwObIbsC
AgzwFevwkJg7muvSdEQagjdb7Q2CfjKml2+28I2yok3Oyw/Pc77mZTOP154I+t33
HVlvtU3FBfmD68qMp+PL8iYabOmGCiU4fqG4iHachAGpOzXlJXtXiRXQoRztIDW3
Jp95DWQOuzCLbdLcyUPaAttaG1l7mjpFUAQWc7dmi4Cf6psvMttp30PYxV4BEOv/
eOwYEd10lCIfu8HPUIlszrf+0XFsWKr3n9ZVh8Zdcqsnv+2y63gI6wFUsrQCuwyG
VnxQw6SpUNRz+uko6bTZka5x4nU+j7tDMzCJka+3YJbxr0aVWf9ksjPwc4B8jeWL
6QNBV7PD1BA0f+IcUH6T1cUlCMhkPLUN88VGzv3zNbmiNCgWtJwUx5RSDFmWgdy1
mmAUDbjCUl0tVkaTiPE14FZaQKXT4g0lNLEx4N2JkkUbB+N9AnTcuuM8Pc4s7/Sm
CmITy3Qeq0ti0SeN3sKkc+ziYEu7ofodtSQd7TK1cU+dMruywmrK6dW5RqHYagwb
yuwHS3ffnHD+5tAb7K4uWr9OuZexY6DBKXXmPaKLKvZZrc5Ippv7ISoBBEW+vKO8
3hK4UiVx0Vmw72dGXUTdjgTaT4CokZgdOD1/iVXx0ydV4Z6RI9VnR3i1b3oN93tn
Sk7ajbq+aXazWZ62QUA3OqyrLRksajLwrw751lEzkxnqHIFTlp4C0pdMzmLwjTgb
jU27KB1Ct6ijGNbLnLewup3/3wtTou7XH341M48ZKl58dgyPjUjd6cvwwVSuX2NG
oN0NHIcmOR+bJA8d3NzO8xGR9sW+5AQ+7TTpBQ3jbXDV89ELlJsIueMezAcR4Y2c
AsI1xDcevBi+4SRg/cQyt92FDdnUfhqnwtZ1zt5XavLkZquwnTgyx53fSTTMod33
IjITtA2/gleAOIvRxPNHJuVNs3NCJmTDzGTfUKvxpQ3sfwl0zou25XTltkpkAFv/
WSxrDOB7j0EMk1tdndeTmeObcYmRPz2Ntc9SEB3sKnySSPMyt67mDYDxGNV3K5dF
yATB3UUL8ZL1DKxL0/AK9SFGJl0TOpOgiKsPl5fNCsQbZ0DmIYCCDpJ3eV+Cbdfj
ZCes4TNfe+5hyhH4m2K0nzk/j6dc/hNleX4hkau0VS2mJlxCW+QqKwxtIRSTtwDL
30wBg5syRcajJHxqx5JLZMWY/YMDCaW8nzabdIHa+IfOGs8uITzR6QZ9BHhkBOwB
hszJWk0E5Zk2ZLBVNurAFxNJ81RRpJkcLw6dVVlkEiA5Hb2c5kuOx5u+GaAnRJke
0iQd1ILOPT/gHRQaGxs1oe/tY2I7bOUkPLoUUS30dYpph1T4tOfO/NfCFG3Ilvkt
/6ap0FzMGeK2KDjOnZLy/RkcWTJQUpxf//8lu5OG64eUcSxe2UFBRMDLP202Wb8o
sz0ANyeU8t0nw3G1j+w4CeG6tSXstKySGvUs03hSEbNFb9Fih0XLmuEEqgBcBeHu
hL6N4sly9Wers3yslrODxvqeUTce7zts2EYSwIk4S/DRvNJuDgJ8/fxsCBy+Idxq
USmcXuIOkfych6CQ+mw8HqM9PYSuYkz9FsTSbycW5pCHGk21hQ+fgI82IjxDKFHI
RDtGMc8AhJcLUs6XvDEqps3smev9/bvCo9OAsJePSkR5LU5wxS92sN1SWM1+IZu1
xzoBSZZT2YRYf42N1lLRnJsLxQsJPk9TgvcNhUb60yCBjVRFuY4hpQQg4rik5kpt
7Dn8dXVePftXFZb/FwzzGrHpXGqdNBgCWVJOo6HDgOFMuvIIjk7OTAMvVB2Vi3bW
Q/NyPq2PQxNgES26v5RCWF2c6xt5kIYbhZ81L+2bDkrk8r20PpbQ1LlLQE3aWYa7
MPSqBzwlv7+/exHad8euXvEAT4XSTSHXp6hyDJ2RvMYBOadB/y0kqEeIR4IB6hfH
IydMCYeq0qrj9JevJJLSeSZqFMNDhSOv4Qu7UVs+sOccp6SUDa8ADekhTzQxszGE
MiGH4gwQ/LQjkReT89KRLuBxj77JuSC1J0SLSUFVh43mK4e4KjMY+sMbseFD5d+U
FziQSnyL0UoEzQZHlc+SPFO0LSL5QUPxUlEIkB+utrpeQ6ocTEHf9KFLSn/MRrgx
3UcnoAujCda8HYIrBKIxfx262Y+skZNSzzGts3oOsggQPRkNJ/kGR0ePGlPd2RJJ
1IJ5kOkge7JB8FljAJhVRrVjmobWCSmIuEBJQP3oQaBUKaABqilAXW8YF0cLgUCX
cm5b4KWyqPfKB7ArcszfORMj9FzVLI5SsgoiS6QacM8AemwHCKYGt0AkDxCd3ivm
8snpgFL1g5T3VW0f6s26voGIeYgVgICilG/QKQETf2hXdurmUZ9Kpo+gP9ngJPFR
m9jtLG6x8Uc7oUXCJdFEsAJS10zATAMiLZND/lcT1ALVye2D+fTE4IH+S06llwwe
+PeaE6M6W5+3QmG9agIf4BzBqmcQtD2uaQbPS1mPg0YdwoxlkanhI8BlWUeomSzF
9bvPz5wRFNsHCHZy/yY5nNmH3a8yhk67PMT5Ojb+jg24aY4ycWq7+r15/O5Isip3
c83lTEfWsDFvXxb4WIve42Lm0QR+iVeUuV8r1z+sgq39qBLybDCfMGv6N/rljXA6
joYme72T5BUfkBbX2jaXoUo/FRx+/Uqc03OcYublcWZFH+p+SJSQ+jKD+d2fpFuA
zj5kfViXq5Zy5Fg4DYE2Su6lxjU92wxRfbCrKlwRwbkr8La2RgHHaf7bRKxGYE7i
CPgyUELKn/W/+u9jXmrRQSaIqLMKrUBDz/+zwJIyZR0JPyys8RnxcyLKv97O6uu/
p34jkYh1KynEfBVgnU5QkVlnxvxpP87Rl8tariOVKjMSoUapnfVLGOa1N73uHvGb
H1TBTTYz6cRCwFquXYBglSpxjTx4fk5CCYADtJc0zfDB1GBneOXfPohKsWWOMJg7
WvUk0b7AiGTO4LczbwMjbbdjHOfPRT4AJvVFiv3QCpDI6eoiFdwon/vfHq1Jj5PA
TZkNee3lunqjTflH+/VOgsQRJMaGV2KtxoZeyqIf0ukJMgRhe8+ibGa4stbnKYYt
xsW34uy02QQWJ04B86Quz+MRI/ocTn32d8VyYF3ukJ1+WSjmSFIPE5OvOc1UHOJE
Qc14FYlh8p/EG1R/f22qjnUDMjSHYcitrn38BLlvi6PlO+LnTCV7Z7+jkn0sN3pj
g5Sgf1Iso6N/s5Hl1tyxxPzshNU46Ky5ekGxsQTI8aMRVDxqGATP0q61owWg8uGO
MUHz/vIF4Z7pL5ZQuXw4bZdJG9cPy4rZ/CpnZqsnbAsE+sAWAj6pE3qgOWwWixPT
jClqwyocykSC+ekk9ANgmqFiGd3xQ0SNT+EkID51dZNdqE63Jd2fgnsPISSkySqa
awpKyqlUutNfBYMIftj0VHZehJdlhBqYIoZpa6pOHrf8AN2q4Xf9M3BywdQSSnQh
9K3WlU1WrRucgsptFlaGsFYTMiZupxttLFSk1PyVHo/9j8JUg8UePE7QNnLWW9u3
Ujp+MN1/PksVFzEfBiWBIoDRNKi68PVqKoFdyI5TlCveK2RgqjglS3ZBrOYpr2fD
UYQFMA+Zcnx3X0kezU2ePA+4AKKf9sf7BtpQCExAImLOwGFiq6NVA6tSgaOjmZP9
/NFHv/j2PGrTzY+QxwW7lNFkETxUMEG2yEFSEVNrOjsWDf2swL7rnHpqesUJqYMr
aX1p19di93adXtR64lWLhN6mCxIYOeMKBznaSyvKN0iYX5bAaJYrW6kfJFJjTjH3
ePeG2sIuB9GCaiE9df8+l3sTTiX+AclGGukoD634uE1DKyb5dCaoUsDc8RHXyy7H
1v/YPGVR5KH/wMtN4jrxNO2rVk65I+6nBpnAvO49BUjua6Ya+zZr88mzAydFINp+
kYE2yFA+8ewGz3lDGYGm4Oqt/AOmD7GPZgrQBTwTbrZRwWMTChTe6XNdXw2zfa31
cdK7C1WO07DabeJGMsaZpRWS5E3yvOa0V7xbfIMroSfWYe8ZfixHFjwl3HEhPbae
WJNV9achz9Kry+7qxM7gbfLL/zwfiCI+bgpGMieYvSFtltxx2mRZjCxiSm96labW
rKxL9gplRAmnhvFOrGSwhHbTKG0DI+tmONgtTIA6HuppPiljsUkYojaVXUt6Pl0a
Ubryr/kss7aUeHAPKGpK069lh9bG+Bg6RWZrVHFzGTqZlI52KaJwxSq73bZvohgz
wmMoHvwuFE2YfN38qrZDnclgfjYaq2uleeUx0sh5mxjXRNd3rJ7kC2p68DRS5to9
ojF4v9USPtkSbyx5n4DJdFQJu2a5FHoouPmmyp+iSH/FiUKWpZVyHCGWiPinL4Cu
RxlDPAcBAhEjf/K0ylDPPJIu52q1prq1oWvTygibatA2w/ssdIx9SSaYVLFmkPkC
lH5H3aK6Mlc5/2Bz1MSKjiii3NvjmUeWY/IR46NLEKILEATOOgcOqx8YJEq3y1Ke
dIiegc5chgctTbW/ON5nPkbj9o9bCdYb7xwQXgE5vG1xukob6UTEuou7jDwP41c/
`protect END_PROTECTED
