`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9OyfLopqbkYjXQGR/fdkTY/4lJLAE3ULmknh5eEQ6jSuD7pTPmV1rxIq6UqKE6vO
yvuO5jzPcgXnkh7aZ2wGix8X0TLchJExZhf+iBTQEipPXTTzq4d3RuXojCRRx+wD
waf0mHHMMvZF8u9C+Ya5pEuNlhes+gQ3Eqe/rTt0nC3aSwmp+RCTS4ASCdV22h0H
PD7G+qfO5f+od5ITZvycCK44q7FVALAgZHVUjX+W4ZrVePV1AIuFxNgua4rYH8TQ
6MICB5DctPjmLUwO1/tZFBy8BPGZfHYky+SaHd9UYffCu/5YAqX7Wd0fKSiz8rnU
tM5YUAUzNxJjKboRVRlnPBa+xOnBZw9QJ+tvpbWCrXQQ1KUg34qCA8oij5rY2iRe
a0D1DC7nVREr88nTckZRKk/GeUarMlKH5Uys3OENJ0u9YTnbKmE+K17Tk8DA/01V
AUm2006bCh+PpGmWwcYkzqUW2sIqd5WDc7dtPDRIcHqSoO3w3vXkAXV6/FnBTHwI
L9O/YHR5heyUavHIBMVn27n4Nx90HExVnJmYWW7be4ZRwP7haoq20o27PUsl2ylL
F1ldrYhhwzw2mhUas0qB5PBmR7ya4Dm7T5kBn5jrhNng94OXj8YPcka5W4jiCsLj
NVwKOXYImDclrqub4Ba+GUhEo+EpWyKWNasz97ZQGY9bQZaBKUHm+/Okqpdem720
XMah/zZtxv51dyQOH5xaVXEqJfxRm0orEe1f3UWMGeot5eACl0ynQzuM+saVh0cl
NYRa3lBI0cLhV/NIFyf8GznHtqA9y84h6a5oitf/tbQ=
`protect END_PROTECTED
