`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
46lh/Fxh+T9hredbQF/6Wi7OO+nywpVIzyVccRzsg+DmR+iNxwd1OEkRi5hky+l8
ws5tRkKZGWYvk9S2QvPMoqg7hLrj6wL6rx5h453vgQ1tmtHuR8ShddZ0DgArWbrX
8vIGHshzTQgCxNKPBAOVPCejbrEbIz02rTC+T8HY0dRzZaYSJYF1Xxkit5mG35ke
eNlDV5ZwlKdCaLkdXNGC0L+VBOqge/4R8slGsAWi/MYIC73h5M9VE3Nuqh1HvUkx
dr9DayEbKeIr8r2SjlCVNXiaTTr6kQRJxfzTU3AcctW7qe7J1AcVCyJBr+4i4lrM
j+KbvGK45y2ElF0sNQdQOA==
`protect END_PROTECTED
