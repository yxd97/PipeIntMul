`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mdNLR8GmF+ZQisxecjFzPUYYQNLpnryA75iVnMakGrou34dEo40y3/eqlKhpvuRN
3q1Qk8LCfYgeOHSX2kV2fqN1G5oKreBlKSGItU5yNhd5Jj1p2KMN+KDEyr4WpRG/
2i/DCaZB8S4pKW0SsiB/FTlOCguCqaM8v7CVeB34EcZUf+3ANXCeb7AHfAnlB6Hk
Yw4UZAHjnCinqJuuEQx4RuV5U0YG9E4L30GHTgPmyjX6vSLrSKW4aZxH9fcmBcFK
ULkVK0DU6f3p6GwL9l1TbmliI3tRc9hm7FdxdEGZ76ulIlThIbmhdP70SYD3jjg1
gBLOUqAUd42au9IZWTd44Q==
`protect END_PROTECTED
