`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZMmv6rOdWqYiQtIOyeyHGsJlIrfuhkNFON5XZEOo1iRtEeC1pkmVyMA9SyyY2/Y
xQ1QbZtaoYwNF0K4VlJMoj6ntcp7danmSYNdeZUahWFkfy6RJ/ULIK7tO1ZAYeL2
FxogyfJKo0EpqGOtVq70kGziPvohLEEpJFP2HH9VPnKa3U0dOV0qA8e5ZAKk59jD
+4VRmZIlztOCOgT3cGgJ7aqxTq02iT4eLaYKr/JNc2ktftBnTBdpLQVgPdYLEl47
7p5hBJ7uVlb412K9PK/2O0yrOhhMCw2bsEsdTYbJpmSsZ9N1QztCNsiHgIpWgJIn
YNyPTiWKZFxxJDKhRtT+3mFJahFZbq4H1GM6WIzf4DEgS90mODTbQqY431KLUzSS
+1q1OsxLlhkuuv800X72zA==
`protect END_PROTECTED
