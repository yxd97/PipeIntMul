`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LOs6SzakU79o4rcUmB4mdlxRwH7QMxRsJGy24YRjhnsfq1hG3UMdMycQO/9MsHE0
YyngZdWNeFPc3/0gEVVH//S2CCgHXKpmTMQqOiTvXqbRfBAmFLaNPjALzrSLhd5c
NTMIVYUv2eXGPrm9JMLrt4Is2wIUn/su0mokha1Tmkk05ZobujdX1KYUTaXp+tuI
K4Mgckdk8esXy+u1+ElemD2YLoFz/5Ko7kjeZHYDj8v3xfhPOY+PTZSLxuyY5rs/
kR2LDtGhfBXDfRAE/AJlO87r1ucw2rS1NiF5gCicUNWYU1Zw8pIXpzd6/Yruejgu
P8CW7CY4vtTSXieylggwW9DyDXExp8f/4abia+BbA0+zZSFQTe1cFiceDua0rLpp
sJgVFBWQg7V5q0tkaW5EwvqvzsdpWv59VNttYvmT1DuMLW7W07Ss1nWRjGpuASp8
`protect END_PROTECTED
