`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfRHKw9Oo2tvuG333aW5Lm7VlTo5UcHU+Qkt4ox1emhRKmZssNqNq+hpB90RS/by
0+APiRnjMvEU9l3zorwR8hHnECk2eb+odOiZo8zUQJKzaxzzF64X8Yx+OW9ZOVYU
d1wsOSyL76AS0o0r9y/5c4pH2NI4ukU7AMU50ug1SyPlo+EYf6P1TGHWvTlbtDKW
7d4xXa1y1T2SX3B9BPnY4M0EM2qTC0iEmWzICuolYLm3ICz5slcTmrrsjyUj79YP
xS73FLLttrwOonD/Qhn8BqQ0Mc6Nh80OX8rjMEwVBLfVKUASZLPhR1wnlDVEG1TJ
f5Qful+5H00GcKnOBg4y3V09+1feYpsUr3JDY0a30CXb7QUOc270lp2/hJf2HotU
lrW1IE49cd3RI56YcfdfiFiOw04Ff3FtjVJ90IRzeOE=
`protect END_PROTECTED
