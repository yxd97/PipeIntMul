`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qABs0zfTlMRV+OxQJfVWU9NfnukclGIaBmKpu3XHTjCss8+wo5BphmCX7jOt49Da
ww03phREEf7sQtlMsWV9VVii8oY+y9ncgMlFdmIpMufYe2UfWBn8glNicjwwhD2D
Y3S1WQTcQ0/nA+DZMy01rzLzxURdaeO66w1IWGcwI8jVa+OjYNDoU/Fk7xHe3QPE
vXLClJ9yvWW2of2idB3vOyvbJ06ShcYcs4n9Y4G3rDz/xyLUHhpeyh9x1/+Ma9O3
R8zYZwkjoQTF21bZ2OJo9Mf7azmqeZ/sPTR/NlmpmxhxfV6aiUoe2PE1P1p8u1yS
7hUGL6X0IqdreUamP5kcAh4+SdkpUrz+mh6eHIifgmJP8TmY66lLUu6Wkg53cOwN
TUmMe/IDy5ZyYiUpjv27Q4ZWI+Mvjt0V5YKl/lxKtOKWnsMKXEr32+W5fyrQDVbs
5s90xSB0udIBT1mVUtNTPy+Qu0QftxAfwlUX9v8BZ4BI1BwKyvncy8+kZvcWiHvD
aqazqIWYJ2WPKc/tT1a5Y5NsY0/LYQSOo2wEPy94U7javaSJaM4rkE9eHQ7p9rxy
cGYeAzfoB1zPV8xIpi5smJoD8CqwOqUes+OI41sSzemW2L3mYqC3ONytITSZ175o
FmtsASAZCl/hI4PsbL4xYg==
`protect END_PROTECTED
