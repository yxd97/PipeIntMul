`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pt6SyETuCglQH8sF0bvoAe8iCzcRn9GNRcVLjlGml1ueB8L0/yU3Fe1iRsaEPUbc
Z0lJUYAE2pWe80ZXLQn1VXwGmEDMELr6grycmNj+f1zu8XG213bXCidC4sbT/usr
RoCAuBFaYy+/8M99iLu1wqimc0sYd/HEM2jjfl/UZbY/dssCd5dejgIY0pXmhVDf
3K39v7Cz1nCsgaUhQrhZi2A1KWeXfDJPMWI7hpxRo1zKtPp6w+hfxaUApBPpqTYv
wbh8DjpHN6sOqW4pmoGiwZbzmqzeHuYX0Db77mIW+YXbMWQwwH1j8IhH+Qz7IhPA
EwIjy5CNHfdm1P2uQcD/Q9yfUgcUcv2gpS7cgP79KZMlTdJCDUs9D8T7FN5Hz4kl
FlAcVamPSZjHfTloToCbXxv7EtaZtRjW6BlnwneGIXNWepeHIk0/iLhZXUZFA8ya
WEoXA8diYN4OStJA9viJrGi0v9SQxMo4/VWaNH7waH4FT2jggFbG8t35xw5/5oR8
LW0o7+QV+bhorLPhQH2qwF378pxo8R8U9IkjRDuQSnKV0dE9zQxQBvSREDFKdfvr
mQfTv16/g2H4Pg7CSMaTLL9ItoJpvbU6JqWPUIEKz3vQhUxvuFMexkFt6NhSNpD2
v0ruhAqKlo7IrQC942gM+ESWLOR5uK7iQAjF8UPnIIbqyDb1kaavMGvJEtIgrJWp
zyqmZgIdBBBnHNQjD5dZ7F3YHcQD5rVIybMylL2f74p1HfFXyNtaaQHeUgtI1Q8a
xPDhLPW6dS2Y6TO9iL2nQxXnejn3ikmMQVoEUX3yUcriaaIWMaeXvb0/t92N+JSV
qq71Kb8T/m27NJ2uQGTxh414EoaRttO/zg3rnpbsd5MYWZJbUepNWzVPo6l7sr+a
5cSophWE4u1J6b52uF2t4Yjf9NxrvZ6SuM9AInovJ8KzFfwcmPU8keghM8Y1LQ3S
5DSIjcUGAP/u1xfHggEgocwdUVtalE4fV4Z36Cmi30yFRmtsNOuXfutV/pao4kUI
oKK+0ihrCag6hVcvbhueFYSc9HBQTJRc4IIsOJc8/QbDwh3oxIpgPCEs1e/R9oML
Q8Ky2juTQMiZkcFG166ffOM+icH1bcxyUWb1xJSXtoiGrWJfugsNIce3jOv+M+Bn
aypPt+I4y6KVh9Yzz9p1Yeqau23QK2aXshS23E/gy2NEFbh+hIiGm5AsQXh/ZYL+
n0WkzgHP/0A1Wpu7OOiUrdWKCbg24xn26jJJiv8cZqbnad+5Odj//lg8NWImBw8u
RBnSAB8bZeSWctuzvKuc8ZH+diBg/M73O5O2Py/7/KxlOHN7fyEPHNWyHiAsmGkU
M/+xnDxEOIx1pwKSkSXYIXbH92RHttXb3IBqnS9nnvujTfNh63K6HuovySgutrG7
nXh2IGGzT1/sgGzKTWT/lwezzm6hcFpFg+cOJH/adDZADJbLbmqK+GqMhGqAy48Q
24OH19EIDM1pa4BgdrUMiiS7+RPllTrFT/6hmMDM6je+Z739IOcBW96CtBTAj3K9
xhzEOgZ0fdm7I2FsAe/dr/knCglEurgXVlBR0KOh0Kdu47+BIgOUWyvg+8dgQuYJ
WlGYrPaNQ+ucFdEKyzkqAOWEFo/ZPkECAUzxtzcfW5OPBy3Ma/02BPF5ImD3sgoQ
esqa1o1TqmTu3KLAR27vGFPkuithRDuwDirfPOKcJwBWhQc9GkAhrBB8jGDCF3q9
HGXHYbPaQ9YqgdhePvy4teM6zqf+HdZPRQEFYJiTjBqZfn3pYGbElYAKF6S/Wv4v
aU0YtcUgGCaZVGECRUjtyayymp21ndaLg03cxsa5BaCPIYeciUtQbCYBcyemFEjU
W13bj/cahkOAbABMqlPP8CteWb8NqBykOIogb4kgITFS7tUexjIIN08tu6vbEvQs
iq0QqQPn+aDiSCJVbeeietVGzOATcNFFdJHtEp9P3UHrlWlDhInwwJpNpWPqgWtZ
ayROHUIM2fEaZ4CgupBTrtuYipgvbKRvHdAFpOl9uSaf1rKBbGp3nhiGiWOZ6v8H
aDBjGsuzZGYhf22We2QTet83ElRdhC3mA8yy6el+HXgdF3BEkQKfspWSV0ijQtzG
Nbk7rUuGFuIc0Txxw1VdmtWsG/h00OuSoBM9tRge1HFOopNvXO7tGQfr2vtdKGho
+/R8KZu6PNXGKaQohdFamFwDTfeRRDcaBN4kj3PXDHkgRnp8nSU4wOYVWirH68nN
Jm0QaZ8cZOWvbYEdLbOg4HKpV9HiaGzkcCIvcax2NjFlTkehYfBLWKFG+UCjoayW
HIZLdsGq/yIrAngaekBbP0aVbTwinPQ3L5RYy1FB29uMMkFaynuMHzLfU87D1Rtc
/8b9g/L8Drf/EvKKt+XEAg3JbPIJm8a43Z+lLYJ9pJ33a/DBlio9eBgH5e3tsjix
zM/krP0geJfccvpzm1/Tpg8xj1+JX22UIzLDcGtk3DY5FhluVO/SW5m7w3WgUy5P
8StZT4N2ZxCNYtyoQF4R+H435lkTVa4ZEvxlnD2TkwgiFigXARQOtIeaop5fEz61
7QZwwAx/Tvnb5YTQq+ba9YJTt51PPGvTr6nzYQOFGMBGUfhMblbg55Blh14i/cEE
L75pSfBCJuCSsDS5aYou5EANMcRxeezS6GaE9GU5CofQPLG5VZuS/IGjvtbd07GD
/mmWO0VWW5otNwExh0d4DurO4RbwvKqClChahvYwizOxrOjAbTPychwhDKBv6/In
bw4cBHQT1wBXHRSWvnWq6XX6WBp3MrxgS6PX+ccrzOAbwhu7wOJLPmjDzn3AOc6o
dPyW3hSxxopg09WN45OnZBrIQOFlW7JxC48vJBmUHhMLvN9K6ktmvVJyf4ZFMlgn
W+6Vj9a8fWpxUvDcyc/tcMbhpDq24S594ASarrGN8hRtPQLNd3Ll53tesPZVHGBV
TThF+iD/n8KvLeONTOjhs0OwLsL/KP7gNM1jZhbUo1NCHxTqD8KPgSkpfvnv/c+E
C3Fcl25vkvU1CEkluEFAz03IlYSGk/MJGvMYGlkKlhVZhlHoPKMBn8o7LymANl2z
YRe4/drDj8TzewnnaDKUMHCOyx9OG1NtQq/Qe5xtxVqXm9r1c4X017pLJGAPGkvC
GYJkm8crgr6aoyv0Bi3h5NnPcw4plgbGU88p6Xoza6/ymIBRFy4p3GdF9pdMBst6
5oYnxWVW6C4ZlhFp6MLE6MOjOjiu10hzRewZUUt4hvePs/wWerfBzP9MimSRsh6B
xet4c95sjit9Onf6kc2yu6MX+Y6XtCFP+sNn/yH8NkV7rgtcTxFNiAkTqm6UnTjL
PAOfX2gGvMUqlUXAPSA6cqKoUSMFR5vL5Vg3Wtcd3ePXDvd6c9sOqZ7X90/RbNV5
Lo7RO22u0tW7a4LcdfIJ0lVcKonrTKV7uKbP4wliPBqgegAQ57/3atFPGeIsxX1f
uRStHb+2XcxGb8pPvAiecktnnNqpv/fo7dOv7e75EuEI+f55brDip8dWqi/f6nLX
D2HprZgRvdSeGai+lUC+MVah3amqglDwPNPJuM252SrVg/ZfNAYyUpp3p1bt6dwo
mPWfx1JpdsVoAn02kWxHs4v2+IRQ03e0MDu49uHX1g3h+DkyWmIwCMPhX/2z0v9v
DgjCvOM6eAEEvwROF3UEfVGkQaFS5jvNuMwRfbk34xLmCThY0SzTM+lZ8+jkcmYy
J0RtwURV48WU+xngcnpjsvf/bPgpN+GrlrxiADRAzPPfPjAG6OHq6DQq3qdfFSIQ
Li7TRsRkfkGDguo6GTuHgDNSFExeCoMs++QhGge6xmzoW7d0ZXKcWKMQe4sO4NmO
bpu6kAA/wGOmoy5V0z2BcZe/49q8bK7py6Jfo4J/VwnK1fMWdERqAKyyuipRT3bF
gYvoXlZRNWU3lJB0wj6t2MHlnBcjSaFNBHPe1Qrk1vQvJNaNhpVLUhazDeGmXzta
MiXKg+mbzEHvH9wK0Ufp6a0ght+Rj+gaCOnxEzArU4s6qBvXDVTnkCX4ktPD9tv0
Ho8bPHiyEuVVh1UWfbe7w4m+iyV/s2VbU+zTw91/NaAs2T8RasbY9v4Tj/4aeFgw
0VoQupQJumct/ZsLeq5fUEJs4yDzTvEvMRhYuhX+Jo/W9Qoy0EnnaHZu8mYlSx3d
8JKw+woBU/dSyFvHTHXasXBpgy1Om5lLyh3Y34N6EPnz1GQdKpkAWpitglCijVve
mYvgUXx3x9ZVIgenXqtHabH/50ZnBjltFiRJ66eeIc5a/7HTbkUQwVASV2a/X1ju
KubnLKNlIl8b55jsvNm9EtqQ9i3/KdTE+5uVqCbN4kmcxq7MGlgQMXgZ6+kjXhSs
EwbuMylzBaY7hQ2rlAcCmriZvEG1gBJacOA0KS/SgUDr7/QnrHNvOY/ZSMuPDbaR
1W2cnHZtHcJQzKvybq/fc/84lUBPr0jNHxQe2F+lAwlfYyQXqL7YV9lRJAlI+dLX
39nE/X2NCl5SNPqXVFgC3sUDU9MUmi84Z5N/N2pm4Ylyl+npFltKFyPtHl77yJSS
zDJC3n+eY65yr0QrNCq7Ttg93l9f5OeJvoiMorQUYjSdgHeyR3lAeP91ELR+7VoN
bGpxUOjPQ1ez2q6Ca9btLpQgK6V/Xt4zUyAOs5FMojuQSu+CE3KPtvz5DtREC5zH
cg2MvzmoQs9qQcUkKdVi/Xk2kfsbS/9lG3LAAk1pEcBnhN4d+MwGC49E7Cmy8N7b
zn8QSkg4sqXNU73ZSjTgWyEwdmeE7xu3NRutLt0lLF7V/raZOPVzEz9M6uESSQ7I
6ks4vNVf5o3M97i1xwkXcZ7SRpcysX21n2TjPtMpNcIFJP5y2UcfFO3YePs48xbN
20iAHGKiiSrRqBEpcmRETbn1cmqzpKpl1y7ehB5dEzfSaodzdnDqlwx9PviBjjxy
jLas1WsRjs52DCW9MyhWKFQHNnoa7SVYuAbQfXvLTY1B5pcsOu2ctz95XM2qfXJc
J2Xqvcw+K2+TjtUAbuaHuz8TMaPlY7R22ZjexWu9tRSLiDOn9UbdOaxe1PI0G2cv
wRJMUdk9CBxftmXZnmZYQdXBWDKiBC61YzZTFMSQiM5HBe+NvrkHt14CgYXYZIun
W4M7c/W2cWPOiH0QCvpdH2uDXURxyYBU2sEiiz+6y1c/oMDMa6/4ZPtPP/6rUjBz
ExMPXW4yQShqIxD1eakraizc/1eagez8N5UbdUHp7XCyFLo894L3Xz/OXxfEBtBM
ljuzZyXFMB3hmJUODjxnmyBh8Yvaui7YBy8pv+uEw5FvRDNtJUg5lQlx/GsCukJz
3egTTYLQhC6x1J1a070uz3ZD4FDoUOKWU0sGTy2++uCURLKd9cT3FrRH+n2D+zyG
oXPI8orQZRPvWAH5ZCcUPv1KquJBXuELzT98wRTiL0vDd2JqxKHs9vPMX8cMxdMS
XVelgRtyFkrHCJjoIzpiEtdibbqnCA6iduMrRSCJP8nixKqGBydbU+rv02+vHxJz
EUz7C+fp5dLf5V/g8Y3NltI0oQn0Vek2Ss4GGo20ZLDemHtJWbwuKCn/gDq7SuHo
acaThBtfKDn3HeGydU2f09YIzkIVyPnO5RpoNrYsRli37uploQYbCcQW6er7u3Do
xfMu81VjPxH0CPL+OuVkOvVqo822cQPZOC96kCWiNG5tSe8XVozm6kHKJVB+KxHL
LBsEsuK/ThLb2tbL/mxn5+e38P9b9LNwkdfgPd/qsSeGXMqlwGAR+I3JX0K2XR29
W5/rg71NjmbAU4MHMZ266+ew5rmvYnLWr1vWfiaWehZly+ejU+/Z7SARf0ODc+hO
cymf3z+1aOEDyBVKQEb0vsBcfpxwgWxyrUprfyaV6YM=
`protect END_PROTECTED
