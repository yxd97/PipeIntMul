`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3pHieodgwctEOAA5O31hr4YKYx1OiiSEr2F/YRiKIguQZ5GkjZpXNmQsKTBskPU/
uLNxA9QJFPH7xmjaqdPGRrmo/qh30Wb/sm79B3pveap+mz5XvOLmZCNVGlRorrFT
LNgb4K79wfGKNKqEtaUsXF0YtNGRBDF/IyycaDzQy0Q47TDQ8BmhH2EINk3cZ0+I
NCxrSZMNHZHnFrM5W80ScwrjuXugVjCNQOOywX9N/qxsLCGmSnzFHgif76CJL6cL
yDrLp1tSGcm6zp39bcz2pWRzZoYMNja0E2CxVNFKD8XK7LCob1YABrJGKI44UmRr
NaNVdYzi1D2muu5B23l9/fMpSHEiIq7Znuwfmy2lt92zWN/xycysyo74fo/ie2jL
vTyi3kmCwlNmutyxunyspiyYn26umm0bv4MF/Nb7f8hUhw/nMNCuKgRtuJWkXOyF
ISQfK3K4UOTvkxM8tys5cQZ90H3aZGPbFJGZUkK63wf4QOIRy7IvPN6aYkpcziIy
DPMGy+bbYl4oTl0+v+4zX3SmzE6Af8dLn+8/wgiao68IdT2NaK4FLQrJTdVIyvck
dR3Zj2KSevDVGKjT3q//6kfx9OG9sLrsKggsLkWz6LQhKB/uf4dXDJDlYS/feoSB
cc72JNzdeUpZKhTAAQN9a3A0dSgsaOQwLJtJeiKFjfU59nUckVycGQfyh9/IImJm
wS7UfJhDk7JxU4jHX0BbD1iXWdZEsKnhuSRbBv/C3qeTsJefGSLfgnu7YXJmlqZt
Oit3R5VxMktj51EbQo0gKMf84PxDb1xOw68lpgQIgJTQkvnbQC77/QAsxlK+CAbw
6EXXOl0EIjkN3C5VPHqKluDRQPHkXce8bgfnuUdLm2CJy2t9bRjoD0I1rZs2p9+Z
yBv8U7TwvzstvkU+/89tjFzKU3+RU8LPCY8nPUZJlPidNCr06u6T5Oeumrb9s1Ug
yTskEs08dmqnlm6LpjoSk6ClotP3IU8UbpDbIwNvpelgCd7u0EzCXHHls253vH9M
mbJeMZVFDR8z2g0Ea9H5li49T9oQQ5l9+VS3Bpkqup4pXqNlYlssrNlfSYIm5gg1
7BR7mkPNzIy90pKbxi/vWxzOjqzhIq1i+D+5fHaaXnb/iBB7+t2bMd+8ek5AwOE4
MGAeejTm5haZ1nrbNqlqq8ny0HMhR4pkpelk7vYFPLl1/+oFSAmRCXDn9pucUGow
GHCaTyI/H1kXKcioFlOvt8v9h1OitDzLTYbsY4VfzpEsjbacS82PfX8u+DQ2bjtW
caEf9jqDX/CKlRaM/FdAk0Yv5dJjw4vWfBWYHaKNoinfTQjhp08SRzRk0AwB5oYa
a5A/bMvgfDQQVwnFil0z+tSLwKTO9dUBbmacQbTqdiVt3KLP/tbvwpvbGnLlhDVH
/iIbs+xFbNe56b5hT2OS49h/rAjy7EfOFsBAbN06NJMKPNXYFp4Svqxzz/qCybzC
XJkxzq3qprRkD1TxDJxNguyRcwUIjXDeOSvKA7XxnSA=
`protect END_PROTECTED
