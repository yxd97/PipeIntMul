`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqHFVNiLgriObL/8ElzZgyrKtMDWWZ0Jf3SK16AU1qJAl+2yb9kEwfo1E3rbr+vQ
lXVEk7zfyYcK7ZWf/SwkrUgHHWJGxWy8gd4x8W6UAdD9mRbMfShL8yhEGFouOMiK
vyk8iBrI1w53+qCZslubDXZ1cNVz7MCYT27el9aPIUZw2HhpoYQtoLmxw32UY0OM
DjhI9CixylKjTJrVTejyAN2a5wx4Yx6NvWGG0U7kmbdb97GKpbxQwBK/SZhNp6+n
IEtn80UD8sS7Fk+hqd4y47e2VFAVy1mE8zpdBIWx1w/7CbPxnjWFcWyJtlh1Yokj
iDyGIllHuzZUcatEcYTIc/JbjwSfRMB9bGclsE0gKLKibzfk8xFDVy6u6PUaFXOL
6CexLp9sogO/mAJLrIZugZxFc3ILHqX8s5NDzdgmk/iWFl0igUKUdwOSXA7d+ja5
WrQn4qi1Tx/Engrrwr0HqLk/crOuDe8eRtKOmFHGhfWIrLngkbot6+ssSuj7gG73
2M3ibTvsiRJWRXhvG/LWFg==
`protect END_PROTECTED
