`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kcunBQKbz/weupNq7BoxK/zMFqSE6EuUNjIT5J3T8u2/0tLFlwYroWtOq1HxLy0g
ZavcRPVLPTiuc3QsEjX2VtaD2bWw40XNyErX0D7Kf7O+UoslALpArVWnAomq+Flm
2VXLHtOJ6y8JruSU/auLFGjnEBTyKSm/U8ERa2Wwt1lC8nGJq4JYUdJ5YKQcessv
AJGZ+SftZ62xP0+uyXlouUUFV85+u1lGGxkM5C85SoPUmVQgQA7PRSgG1RtYByvF
rBTp8C1h25lsHuXNK59viXiqpufmmDOphppqU5AP5ri5DP4A+BHBYaqm9Nvn4q0h
+79fRocytVswTPS/AmOOMkSgaA2P+/kxmwGDaKxNNlHnQjOUBbaUWur/kmYVPmMc
pCHYIKUJT8JHPZ4UbCz6AVGyT8pNRdi2AW/znMGbK4jIlBUOLKvRwz79sBNdAw+g
P+ogOKRhBayeUWgzun5ypzZ0xmXqv1iUkFw6IA5QUQCu3O3vIAG81oIfRrYWRqIw
lBHyWYNSv9I7EJ+HZXMGErix+tKKSvZedG5g96lzT/qjjgiRI0H/eMimjraeJIGw
s5EXPQ1XBDbu8wr+sDtk036V3X5/qEcIZfFJOQBis6x412zguAgO+kIUuPek7Jyz
1Cog/qEYz6LcpE6/WYd48A==
`protect END_PROTECTED
