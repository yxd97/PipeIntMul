`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4yLMxhYA2dzDLeTkDq2WlPvig/F+JTVabowG/rK5gBwPzTW4tsnaE1b9TuYCIQ4W
fkwDO93HjC656KKOk87pTTDal9Ty0B8heSiA3e+k68UFl2wt048ScGoIhuZxXTN2
07UCFNYssDJlo9DkZTPylo99I8LQIA/CINNciAzeWGNLasYtqtKPzW5rAZFERQ4r
vdWZCh/SYfdsmcICIH5dTnYIahcZJ0YnjKk67t7WOF2egV7iB6DJ4AabNKh0MhKD
+KdEgn3iB1NNfczi4EcboSRUDnhiRCgyoktIxrXcWRoKX9Isoq8ptpkoI/7wJoii
1C5LdtWgzEVHkkba3V4+bZTeRwnxGKhKIsN6vUzIwytNAay+QN08vcsS2onN9NHN
QtqMUan7vuJXe0k+5F5wA7VRbGILHPpxHT/IFcAoe0EqLhElytg/IOYHYIMw+jEp
vE8nA/wSbhu5jNjShChZuCoIW/9cK6UMBZ0oIh+ZCJN6slUu4eyJfXxobdu/Berj
4+UEEUh8PfKYVZ+4E3Ur+C/cCXcTj6ALTkylIeby8vj40ZwKOos+PfxYv4RbTdCC
nUwGEmIy+cjQWH2dgxpQl7MsZ0xCW0YqO1DLRsXNhsQIfcwX5GYhqnhNL91yhbwa
GhCwWP9+dpPNi8uOEf/PQBPmNHdxlPX+8HKNkszKXa0FxOCW9Megfda2S1+CCP/c
t2/ARxA5Bk+qfQ6jGMtYs6xSPt5TtqSdyppmPgvNBC03Kf9fxGa+hvNUKpGs33+G
PUfqewy06PqVoFzoZJeJyPKVnUDd7a/N+tT3VLu/QVy5EewlTU57IdN6CT92AfQQ
dvbZAGwkio9kRuMH175g/+S/KJ83YTfzbmZDjIEJTfegGV55Qw5vSZdjuqMrHjGC
8Zaw8Ywgo0G7+6f43wedfA==
`protect END_PROTECTED
