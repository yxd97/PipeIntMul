`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bGSYFFxrfsxwGDD0DqW1/La/7b7/zGr2IlDlH4s1mbruHdKTvKbXG4Kzr9Zz3/L2
nyz1c9XHmKPy7ueNyLWiPiQm3TfGKMDfaY/dkhE5lBCxDvRf7ixszlzJxulqhyZP
pL80yMUBlqq2hT2B+I4fM1UZj4FvApGxVjmGiGjq3yD7pFBSgZ65qhAPyWCU7oaT
0rqZR3+SF9j7CmBTDPjSaQlQ4mcWrE/JVFH7hGDErerB4GeFORKeo4bJ7rdkHCQc
gitAVq7VrRU+AinM0cuWLMnnnfM0NH0wPt2hOaQjrfuGfx7wvwE4t0LI34N8EI+x
iC19Yg/LzTx88oDq3kAdy6OHuqjk7shzrUVAo3Dz7ChlgnXSvxB6KigEIk3ixtmL
FPOGLobHLf+mvLI4tlNe/S19YrHMpitkuB+bOeuh1TsOw+F9Pu/3dalZ3vxyQOXU
I8dYMWPirZMtLb1PIKyI9P6Ponu7oFms/s1TRyt07KP6vVZpoPqVfgPrlAU0W5KW
+XAAxeoMsgzlpFbA38PaxxLgrjC7LoWjUxAJk4r2h4ocIaqvvYO1PSY+sYQexAI3
k1+W6jLjro5JoX59m0W9RJrKGFtwuPGNLo3mjxkxC3zhuZWGbmCh/dF9BsHFn090
Y1nAjeTSn3F6LciTH1VLuIXEIRpNud2itFdAPbIN5W3PpuCqG6QFXMqNKtQfIPW2
qSOecc0qHeRwAcWNho9DxK0EWJeeo6Rf53FJOjKmx3uXss+Hc8JGp2Pk0CjpeqHn
ySnx/OrZQ+iuYS/fLdkpxoNLrsaNO5WBTd+mcsWLLOYHdp0j+PbqPe5fdjTOWove
oaWj7mPfvzq8i0Vr1BzpG6cboahvEL9cZhIknyLLU3dWYER40cCqVu8LAf3lONsy
cOEq4WAHOyWIUSP/wD1R8vzyX8PpumX9TSi5lLyLh0jE8YyBqrSlmH73tvgIFa+g
`protect END_PROTECTED
