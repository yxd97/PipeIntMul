`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wbf4lnwqGYjotqNlD2wLv9FUGP4vy/eeOfM0qVzjuRq/0yMJ9sgqxxseTfiRV1V/
ItZw3bOF96JnbvzS5Nqf/cSp31as7JX+P6nSFoKBgRnz2QWuhG1cHorZHoMNclRc
A36fGH5gJt2QHBoY6h7PWMVdyCvxvcKdugOFoxIyUUW789W7PxlP5tc+1ZUkz00K
vsLFVSARAfMQ2T4kRQ/CezFIg176cmkImToPNJHM+/IvohBWZs2F20OITsreJ2VG
EZMdr3rWNbDbslAinxDa5bqdeh3tyza/3LO9LlDWx5Q=
`protect END_PROTECTED
