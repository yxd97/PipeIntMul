`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uSqnwvp+Eie8I75w8PteyKyCPD93EL3gJ4WnMSM8i4LXTcOlqfGl/kwDLI05x6LF
rXz2/AmIJu9GGXZ35OKRovhh33UP18pQoILRrjEM7wBbE6bLPEg4L1DbIxO+vISR
QwjaRi2IlH/SIfIHbkSTcyWo3eTXMrGPnvOZFxm4SAV2sGYDHLtXkGMkN8ufTMGB
cFKsOjKhm0GTCymfGVwUCr3nn9UtbNA0Ik7Wy0d6AX/5lWRuhhbDsYpqW2FfDKt+
LTVl9ICdkB917RcVTaqDa7pnXYGU9BtKjN01F0FDxB45FzyfyK1Ix4F+T+3ceqMZ
sq48EHEhkBGsu+xXMm6SSfAUwvvUbj+ze3+icaM8fvrg36JdvvvqeaC0EI0mOECB
j4UxpXPqZfuoAE1okVCPTrZDxptBrJQKzRrs/EjTsreTUmc9Mkjw09Sg50qUH3sm
greqkFLHg49oQYngLzQ5gZLIVz7jjh7z6wDvA4FdQHtfCucvRnBlxzXuift4nH0s
`protect END_PROTECTED
