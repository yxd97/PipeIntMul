`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oYZcwokE6bRCrQup6YS/BprO6CRCdga/KfxTYexZLSGzyNqPN2l2r/i7FxmJs2kf
IOWwQPbewSz7BKIWIPp0KEFEEoFIiYn8ti4dOroMnOQkjs6ALow+yQcWDJqoazrp
so2UcYegADrYv1yFqHpoVX+Q2SGn35rRaXZgX1p+RaDbBREveK7X16UYRiNZX+GH
zcoN5ZJRpTOPISp92z+PyttnFoiF25J019YsfTurR04Nzdi6/rGFnRs0Kehv1jh0
nQvKxMGmY6LLVFeWDKyT3DkkLHxFbMRhUDO8Xm44l5rmRwcXRx4z2sn3VG+h0tJ8
QwoZXvKif6M8QIkuSiNndzRSmQPvaVzNPb45+36yxcF0UHtSZSD7OSfPkELLs6Hx
1GnYZGhsT6J4+VV4w2ViqyPzwtkhQJDMudzYDfH/dgQOYVxs0J11RtgJhooGwpBw
KYVZhI3KcNpH5zV4BWWodjT24p1WeNgw5Pt+krJ6VjuAi2+QwHV3Uss2SfkiqlXO
F/JWg1PkY1fH6P33tuZQsjHOEEMFezuJQI1x4j2vE1/Pg85FXIW4yf/i03lNA/Hc
`protect END_PROTECTED
