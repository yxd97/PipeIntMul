`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jpFz4gDOSOeq/AwI57Ur3TdQIo8eKC1Aq+oTni+U5DhY4NuIsI6E4uIKxzEjJtJi
wEGkLWvAJSfvFREkd2zU30lvjIRqRD2TuFrZWSvq4EBVPL5TrCxOfG/X0k0pSDB1
Fyn6EFqjCpUddJDw2I0sdBldCWLpBfo0pBrsQOlWSKmB1OfoXfJHAG2zTb1LtPbY
vB7yomN89taYgGJ+UiIog6PhrEzmwObeg3DMAaFLUuBQOxjYwhh57Y+PgKeeyJz2
31FRnQKZmqItN6gurd5okyoyu/4TVJHVC0L9og56amsTCNs8+mSahH20CDjPBApx
HDL423SSNTGV6YXx53ZRlQ5w05jp6DG/+oxaFInLQzgyB6JsRo45bokIt1dGN2RK
yFrxPXaZMQZIHR7ndN/1Z4tmd+CUpFSRwpbetGyMs5NrgD61TMRg1lw90+Iq6Pa3
JmiS/aKcYkXzFy0O7WaGCl77H5TZbG3iIvJxS0UlIAY=
`protect END_PROTECTED
