`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ctZdsIAgXzQfpjIl8n8R3hOd5OQvzhBYfLSIzUrSFmfTRlZVc59QpfDC0iYnMoB
jeH9wuUT+ukAKzK2q+yPYD+sSYipTZfDNMf8BmhJY1AmcbjykwDfLM/+pUY4s0hP
c7vSw0xH7R5Z2e2waGD6Yn84T+Z5Lm06lsJmS2DmBLHGscYml0sCxLAcj0kGlJ90
sMXJFgE784GZ4GX7MLB5Ox3mLNMJmP2iWK7TL3oEdz8IqDFXDnapTsCAyNtn1JKE
xx/GUkm2H21hcn5z5Hb+C3GPFD++ewRarTSZ5uytBUdpAnBGIAEujVpXtV+1Y0wI
hHYAkIQ0OrcaxmeR1SoZSaSJIpxLJAsP+yr+3MCgkR+/WomC3tN6BZUqybQK1I4d
0vG4g17ffimva6UrNh3+9pIwArCjCY+eC7QghJz9qTKcg412kTDr8zZwhFcyuOQt
o1QSPBv0av1A5vtUeWZLAw==
`protect END_PROTECTED
