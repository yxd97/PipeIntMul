`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pEgpoj21zW4LExpQlHk/vx8BUaVc/xzSADJXGaS0fQuxIhUKKzWkV2TXqCGBI5F/
DUfYVzOQPJCO8rkHapBsd6QwSfjzcBwEdg1GX8wSnYF8gNXlIAgdrHs5B/ruX2Wt
+8QbUbybk90X3rTFSyj2Kutu838psTKRdeWzDUuBqaTZ1QdkEUQ1SNSPU/gB2846
DvErMNJNtnU1BGUU+GXczCUWB8mym5JAHhjEQk6oiRV1t0nqMaPdWY6nPpSC4Qk2
M7p9aw36YyGsHRHoVyll57GPZJNvHb+qccCI7yeAJTTCuUq+zrmwF+rUZCgQeKUL
BIdb5ceWWoZNo9SKZLs7Rj4YoDGK88DplnqfC9mkbftoXtNZiU3KU3KxnWqdisM4
qo7Andx2lPQ16O3JyzoGRzgxhViKJf++ZeYqOQwwzMCVjBZbFcOVKGfdkl/6fiIg
/3at3ruMinGldx8f1s7CMiXQEBvGlXaJFT9010BAM3xdht15S0RqrRRxgYdlylAh
wX7mjAfb2GkIXQI+Z/568DZAGxvVUEUrFfxXeOUGg9Tc2s1dQylxJyg8sz2NqMSe
y6Q0j0ZpUnnBdTtcvhWFu2mDsBVe0c1dAQAld25Qy9lTdA+rkY2LP0VWI5HUMxAU
PH+JWoII/Z2OsXzzDK6zmyZzOQNOdcJnYIXK24HDgn0=
`protect END_PROTECTED
