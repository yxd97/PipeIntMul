`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I8agbVYuGTFJLTZMMVQYCix4VSAq0buA85g3MPALZfcYSHC0rgpLWHR0+L60ttfr
v6KTEMFM92s7OEzBrvzUrTvT4zOs/CQAe30zlzsC1q91rEwycGeHQzZYKwtDUjYG
iKA2Zctyi1hWY1Riehz4Z84VJ5Pu8haiSIoA/KnF207RqIlpqeiVgDLQozKhG+FY
uoJU3CU9vEOafQDnmJilb69gv6L0AwjkHaUq2Ic7oQPtLzPiGrpuuDJE3DKozx60
BMlDoTC3oAB1QHVuOlY6Y7V6UiQQ9/69ItaYPDaK/0fmq2dOCNoiH/pHcPmtcuXI
2BhFc+U7A1/vSA881BsawfYBY/p6gJqY7d1T2n1HpexnOVioX1WOugDvaRhlZukA
vebzQUkOo/uA2C7zAwxPJpbSc8Dr1ge4tC3IbUCHT7ndZ+EJUNZBXBrDlI4EhP8k
GzTjOs8d6c9sQ1CvLsAO4ssONgAXJSsjzQ3OU+Qz5asjBUwVaD+2fTbFJ91qjvqK
10nStCyrHJdjh5/Abxm7FFf2Le4mxia49D2DXsZ8p93iTXFCXUsVYvf9mzk88wJK
zXEllAWUZQ71pcO7j9zSmzRVHQNuK2Jg2c+wVn7arJvdF5ebscXGBa8gqcdveBuJ
vKLXlvXecLjyF98aWnvM4Fr0TEPmpJm5epNdXpfqUOIy+3y1rSfgQp33SY2r+Tbm
5rUVViHLP5q23+ywgnUiMBt0U3nYZbihXjuK2T+2v4UqIkT8cMAexz5KWq9bFea7
sPMaYMwU8yMu/oXd//114nroozsc39BdHwOtbuO09iiEbnlEN2pwPFpMvHjozrkZ
4FH/beYU0u7P+rzoTbP+IsO0VN7Q2++rgFdGIjwECNvFArNindqSt4oGdewXcpQP
c/TKjaxxd6yWL0UdRmVUKsTmNmKbhGAY3+bC6p8p8S7oXJRILXL2VqaHfikUNUTL
YUVTXR5hsGqHpkgu/wMO1SbP4cy/hlt1pc7ZTAG76pN2v6T0S0R8p9fSy7miaooy
ZG05eUwxbkYwCT4mjTqq3hDQkYRPbb/5NGkNTRNXPy6LOF4EHQNAd9c/U1lrffUy
`protect END_PROTECTED
