`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wqQhuh00rpk+ydnSqdzciZ6itYNTRPC3lIEKpdd1FUtUlBQFCuz9bAQj9+uRHZrZ
Pk42WGtOz9LOJTiyqzxgEM2DIWgKCpP0OpTfaft0zhJI3nJNQpuIHrn9O0wfaQWy
S0xx0PlewZclBiFPudG14GkCMIvbMZYSxV9g7kZte7k/t4WbC6GI9xBOBec7+O7B
GhM2kApBf62WmYOb076QYC//eP94szl/3kmNNRbxI9pTu1S2su5OJI8wBBSbOkz8
/6fxDOnZ/3fwcRaVzrlCSvpN1SvNUtUyoNIOQpzHCD2JbXh3NE/BIs/ASZas/1/1
14JaQjzptWVJhPUu+asGJQL3onW4swgnTFndn9OZo51Yb7rjvzx98fada6/0ewpx
+dCVZa6USq+89pFtaDHj7QFAJnlQlfmKNPJBFdJ6deo1LSRD7LkOMgBx1cDAkGXy
dVDXwgmJ0z54ltmFseixMYPK6nO6pFuBhKK0DANtrRXtWjq/FPDpTFFoMt0QsuC6
foIlAnuLo6vYArywDkuROeFBKAGKx4vvvOVOP8LWnONINPdJ8WP/peeI0HCRklcD
tmPPXDlTPl4DEIFyzYOezvV50LNGcINuawyPKAMMOFGlArLMSpREkMBTkCZgYQcp
hGs/4PoCts6HrSaIf3gMfA==
`protect END_PROTECTED
