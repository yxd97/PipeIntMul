`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WguBFS8I2XJmPn2/F6Ic14d2mT4hqeGAmPHOPKXpLZg4FhtescuepSpfB0NocxbV
tKoB3LbTiWm8mZm1aIoxNDLWNCQsGPgyO0Q/zoP7oroUOWcas+ZtqcHRBytx5Jh4
zJgbc+SBWSUsjWFOAAgIYoccsOvQ0SbSHhbULAZ26oZlsOKBctXIac5fyzRw8gYr
pBKNQMn2mSfyaaYZey4ur7cY7FxaE5QbmVGfJ+8bM6NAdehgZrXWOS7tTSiqOdKW
R2GFK6b3NlPo+MHgsTyQVEvG+jnlbyPSL3tGdWwKxi6oC2Dq7IXk0mRYnihtG5EE
XA2JQDidINFJ9GUjzGcuHQSucvGNGbkknhGAPGurNU9Fc3b1dd0ncmVTfvm5Z+IG
0hZkDNT01kbXThHSgAdf+5w79gNr+5SyhDyZJw/igVbnlsCTDX5ovDoHCMVDzCn6
y+5Gsk9xgmWfTTMIxgndvLhH+091/UogUB3ZD8Yi9USQmDk+d0bcOs10RzGkNZZl
LhFVPanD4oX7pIKiHuZNPjhbS9Jkwzr1e6I2dsUmzOAc6HUKAHKJ6HMWRjvVNqCg
RXAWvgykkCF9F8ASV7KS47SLcprv/MzrqMwJE9/qdCNk6npWOiJeIWEdCIQJo4Y6
NcXtJldluNDRcPjQ5NkgkMrZhKaWQnRNdWqMeQrViQgl97Naz5dSenKiVZfaJhca
PE9pYcpl4KmTOwovGqZ41QBxsS7jjD4AmhaxkLB4KlOWptR7TPxRsMOK2EjdmHBL
hxKwq8ZybPcCAobxjbpRnmIKwlmaAd6w5+p9WhrDiLpyOIuEdgIDK0rgH4W9dkqE
XZwksfKoaBqlqfxMT5ppfaNniTgGbXBkx3N77v3ACrdd4E11MoGRZcr9SkbswLcc
sx1dutqBhrbjXMIpOiRNWhHWilvgCEoyxFubPKyAPh4URzrXLOs9DoW/Mi70BfVh
z/uuOjOt6bgt/BZpTSuYscbSDk76LPeQQq9Ljiuxks8OFlEc7QVyZPv4aUx4SZ7F
+Tm5nkFXQng9xb9KKDF0ZSsEsPhBTeXSt6VaQVCHxkMXPZfeoRkU0zW3kwR83bkL
h1vyuCWPosVoyLjIZcOKgJtybmd6ulo8WeXA/GId0gyE64VqKS2a45u9KebhznIm
SeMTB5SdaA3PAY11s1fTkJN6dkWQyusb0fO6md2zG8LV1r9OwBtvPNuB3WpsD+QC
3Mqk0MhNu8j2AXBakk5isIc8/3hkDeuViJ2swyOj3bDwiIP8l7LuGIuhIHN4Tlcj
O8xEBZiI0XdHiDiz9gv7+A==
`protect END_PROTECTED
