`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/YZ2+nJ6HUsmrnsD9rwRp1uo5cGCpg/YTmGyb9mBEuKsf4+5QmJxn/700lZ2XcT4
tC6gvo6E0EwC9GuDc7sdP80KEkPl+Y7Shig80BU2u43dNh4owZcfwbb9G3yjIJWi
1mhJQfBlsJXCvKEy7K5i+bnA+tNXjjmyvjvU9MuPRauab0l7NW5Atx0FgNVA13KC
gkjMk50tlUPBS4HxYlHuvA6/t8gnHUIeKBb5nmtKBgj20QlKCD+VdKbDkYW4Xw69
h8XhxWZO3hPXYoi/KDTuST7Iea8aY9QUtK7nuq7dYLdChEBT1QXJpMQMR6wAq35A
G/81sV/j9LH+e3cO7n9zZr9ERyN/fYtSKgDFJksiGv7+XsQra184jOMLUvyYPBzz
oV2e3sfnxTm4GuvKQhm6Jg==
`protect END_PROTECTED
