library verilog;
use verilog.vl_types.all;
entity IBUFG_PCI33_5 is
    port(
        O               : out    vl_logic;
        I               : in     vl_logic
    );
end IBUFG_PCI33_5;
