`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g8g/9BNx7fwM5CCkriwVNibgDNLY9slAC1iJ0SWHWdZQlv5s7Wc7uXFGaXLUr0ws
WwT+PEB646W6vFVFqdHlb35RTpr07fEuA+I4Egj3jTBdOlZTx33az6X9pDfmVt2S
LQuNimLhnuPRP5hKJt9tXKo6XpgvMpTC39ATpzdIUwYnhNVd1nOiYFJNbXve/3Or
fviyylAm/1Ok3HoELihbD9mE0gubTZQtzqBbD3q/eark7MNBnQHEv7G7UFFTsHn+
hGJ6hiiGsExri+GWXUfmgxHbl5Lr3GjbBeNHkJmEcSlRNdDLYVyjlx/MOd7HbsQu
ACAux7EVQTynQeuZN4NHqQjFDzjCkcLoMMU+V4lTfRsLZT52XVjbqHSurBpT+CRI
`protect END_PROTECTED
