`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hpt5BxXdZpcOAWGfWU6glAddEdOqlWe2hUprnJxyZqp/jL9LAE9DceovcETVxv1+
4rRq6m8vPf8cUV2PELluYp30M4OxhgPdpEm/xtU6f3Vv1MMwhDoR3pCP28+ouGs0
pmPhEM6dFHS9eRxuvp8xgsJQDD2rzz51e5U1YLnSIm1nRb1pHhsgrMFEJ4k5Mjo1
kKnL0X/m4+LRsmPuTQF7l76jMlhchNNdgb1434tzydCx+w7ZjiYh7PQ+9uMdEyCr
7bZ2wdutFLIPGyXRi6EcIbRDn2MyDrSbNbNFog3R7zaq+s4XeV2NxmWv8BZ0bhPn
khPh0AqQARZ1eBBpekgX+9ItJqhKPcT6MizpBzrnngrk3Hi3YmqeTU/Vo2IIzCdJ
cnIOq7tjdsYRo7I3FouaYEfnNa/PR4wlOHq0uLQNmX0=
`protect END_PROTECTED
