`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGmaZOBAZHgQLZoP6szXuDr5oOLOAztU5yCh16eumuhOHAPGxiMPy8vb3Hwo1DZ6
f25pnfquPIUZa+A3GrvRxng10ZxGpsDGNSlHTvsEjLcIkalAMgzphu+iOnrkuiJr
zTz7y5Xv8hUKjMDkIrjKOjKOabLg4YMgIWwUqynrQ7EtJK8zEMMxJWpgh/IKeZe0
9ZyruhVeBwTPw3t/ohr/lJFJ0GU0taxzWgl2j+VssHPI4FANxohgCYIa7EE6iczo
z32ypBZlF3Si4jhY4gUvBSxDh9bbIABCOYkytAtvRODzA5Orzk8/z20z3TeeiCab
cRulj5b49LjvvLfVwZkci2rRPCObH4l4bRBo+7sNnbVY+H5oeiE/AFYNQ5coydJ9
HSW/30eJ44dIG9zAuZE4mLQdu+R0MDQoee73U/n5NSsTZeD5EbBC0LDTM2zcmrpj
T99ofK0FxaHNw/eMP9PF51q9hoYzAhNv+Vf+lUasDgYKwe6Rx1EK6oBR5nfP6XLF
m+FDplCpskv+9nAwI2SiykpokE/6YNc/wAF3XSNl/ck=
`protect END_PROTECTED
