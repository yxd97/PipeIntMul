`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkGZ47VAUo7ZucC5QherppThJja22IeI+lMD0GPcjekNoYU17PdIopxP6vVKmZH/
S9fhcWxm7s7BAB2gcQGTHXCRwASHh0+uMpUPe/GDzvbGfzDkZFZAAH6Vyj1RpSUi
5zq27u8cLB2YVGJH76UFzkku8s7aCiL0L9s5/qRANDhSZLXn9kLyBGvU9iAj9vl/
UDpQ1a2JlEyYk8L8lVhLy12wbWGl1ldmCyAA3qBWJZr4sCJx4xCSlsxDenb5LnCv
lmI7+DJd6ceM0LE4H4mFTA==
`protect END_PROTECTED
