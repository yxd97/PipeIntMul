`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8hZVSj+EkUQdv7nwcOAEspp258XAXg4S5sCEDyvVJQloPqOLJlWKntjOfJrd3Ykr
EmuEvp6t8Se6HLMThqdVRsrdYbBDIkaCxXwUJOaUhrPTu0fHuFzlGfq4PgvCcQal
weEjOSv2T4C1MyVOaLzADN5WreM3z5UD3cNxtEJuHKsy1Z5JYw+qj2lpBjXUUxlJ
qOXLP2FAgiEJFDAfOZ2yUJQLnwzAYUGqu5CO3eGhI07tisX932x0aDosigorg16g
/RNNcakebFIyqTeJu8dLBXxCmFlbCxZfSPCgYURUme/MV+bC36ZBrS/ThFFsKP0G
K+U48YIJAML+ScznssQ7+L/L9znQIWvK98HCJvEnaznrLrSfK8F3S9CxwKO7a8I5
LjjIBgGeD+TQuVSWRvxcSN2EEMyh21iFc9Kc6QHSA9fEKsu6VbbjWSuwzupMHjUu
AJrWi42/rvyp0C4AXm1Cor4Yg/8R7I9oMkSiYdTalh6aVbEVtigOjdqZ9q9Egc3Q
`protect END_PROTECTED
