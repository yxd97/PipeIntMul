`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixGza1SuGIDxcxRy7EzXVS9NnGtau1fItWxTv4RlMZWJAn6Xii5EawNeLcREZhQ+
B8RQK/Ond/0IijRpTWidYU+Cm0+h3ugzHA9UzM9a1Un+2vjCQhAx8a02CTz3vJoJ
/d8rBj2JcFqP6FDF6xTL9kc7indqcI6xpIkmRvyHHbU2YADcssqSk6C5E0OtmFIs
RVgbPnFLzDXFEHdFRCnNj6tVwU9DYF+K3QmfiKWAGgq4yJnI1bNubYp1l14824MG
1SMdWtmgGzk4NMsTvnUMC4kBKCPisE/l8kKjRv7lfC4XYuNu8OjgaPhUx9n6TXh/
Ugzv/BW4VUC7ht057Q5ZbHne2ODbp12klX94+/IIWcQlERyvyWwxCPa5OYzG6+1U
VrJz8H8t0AxjMAzrLRTzwtn6N7+g2wMVvJs9atyA9D/q9OteQGNC2LR5YqQQacab
`protect END_PROTECTED
