`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bwu32+iwhl5I5jlt2BGhHQKQ7WHmn1hjiK/NqY1asES/bCZJpJBAFGniWMdeDIlT
mciOdJshwf3Q2rAaaizlbEcCSnwt7DyAOXyMX1vfNGIc7l9ki80GydRtSBDrJiIF
ZcoMIsBXYumR6SVUKrUwKkpHwXIHSwMu13NKU7FikHJxxUaIr9wh76LKLS7PM/Bx
ii8AC+1tBNOj+jdEwlrM2BbSKs8PCJEtQhYFuG3Lge+o7Q165sP4x6xUjHWFSoNL
ga0OGNwzoEBw0GHEVK7tPpTXrSE3kBzY25h7XpfPJfpNVdnDhWnyDp8H6Jo4eC3x
9ur56lPxAJt9nRyf9UKdc5eW5Rm4j0Qk0urlyw/TOVE53pWRuVf1uPUtf+muj4Q5
XNIGK1ZS5PO0Pu2KJX405IWYAL0R4Pbs10iC8xwAy+dSrz/RdkEhXu9gsdnJepxp
TrAIUjjwvMBHbiRSuDa6+q4Zd+Q4ad90hK1nK77SD9fLU2DgAM9HvcccBJX7Ypqw
tSf9TaC0VBrHVdUrOxR+OUaz30LKi15JYmlClCBD+IagHeECCJybq+63Lx0XuOg2
2fpmaZnkxma50wyr+6WstGlCrWIicWk56luWpfp6qo+ehngK2bVJc6DlHltlDh67
`protect END_PROTECTED
