`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PfWzxBnKjyv22pAdZKQeRdB5uMsXiOh8Rg+qf+MvK8uho+EkJCiN103JpF2zprBy
NDxmnMQU+QIyZU4aWDYdGiexiTveYaxoBAS3Baga5mqhj9390xyeNkMXnpTDe5a9
gmLYlNB1FM+noKoYUXqqp71NveiBWiWLvEBswPLJYPvJDAlgv2MUV5qWybX3zFKG
rYAwjclaKFoXVRzUaO5vpSlq0ZFbTPFepwlLh/g4uih5MsCyxZ0jbeqOFboBIy2V
8Uc661zH5fLZEziHxNwXHA==
`protect END_PROTECTED
