`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PlJAm1JhjEiPPeWQXB2y+HqRDVVFDPYEIvQoqLP6prN/WcJbRXcmYXIfwYa/xYgm
rI2bAFcsV1waPMI86lrmc/hZx1whHivAO/bFy/oI96AIJCR1PC4ss6Gx6cyphkbv
QBMHHG5XRLikocfTTdJ3rKCht5I6UoMZbtxBXHXsFP3tmjub83qMNrkqcTE0e9Ag
VRILHo0L5MDG9NJGeZhmvLiUqF/Xr6C0YaXAhk46b8VjC7I+A/svGoOdIwUao3JV
oMEWVBGdLR62NrOghMufTXZWZSHgZVH5E9cXI1IbYQgZaVcl+sAFMGt3zk2EXLJp
YvMwIUn4cOphd/HO32HrSP9+aAe8ajCJOS4bZy3FH2L2TgsFYyRFrxI7GqM93F1B
W0PdGiiAT9xYJz3azHY6aqLGJ1QKSUzc2ApXtr8QT8bytUvNWnPFD7GPCB0ju6hK
lwvDMBoM49fUCaCKom2SRwd56XMfyN2rMmmr3L7w8DIFiUB+5pOpVuHmmpKCT+OL
TcBhCIxKPFMNE/B46oDgr9WTSjpV2GpZ46fNisdLb14ljL6f0uOFQEH6FLp2bNh3
aCl5HgRxqsMAeySI7BJ4QNxQ2lRusKnlkEwvAQJ1g5ZkgTWIyhp/h+IiH2DMTEx4
KJtid2/EAKieMPgfgK8brQ==
`protect END_PROTECTED
