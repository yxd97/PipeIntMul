`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLIBDydEqDRc0DTgaINEyrenEf9H2qlen4qhcgN21g8t9VbaqbJDfQo8Smlhcpto
gh0VJAQVq+EsidW5PGnHBYM3Sm5eipZLP+9UUwvmAUpJ1jkI7a79tg2h4+ue1sK7
zZdCFlp6yLsbRd+0kqFSM55sKkxRaImcDrLIUfrxKvWQkEdbSvNiBOtiOiU0MqPw
+MZtZRbL3/nfVXTAEAo1zOfRBG7nZ4P7aOtbutvOO+/UZDndtVWRKbAruUfQGX3T
pUCTOX5cIB6Lu6FHHl/XYI9NLgYjly13SSB27w0+JGCz+YTCDfQAs1NZFscTalHt
rauUNdrgyPN5jN346okt20+vSnZuftQEWzO9U7qWu9i+O7Ww3+ZkgPJpxmBcPQ6L
qh/z0MJZthz/PcfdD5hiscAbHUr6SLk9o5ugsAWx1WSoJ3su8hbmoQP45n158naY
ZVR6C4448ytsBN+XQNgFI8+/ndpw+5fe3UYsex6p5I8IbMm5ZfrxnYhg4KpJ9OrG
yaDVLxFO6R1Mjz2HJK+E5xUTW2GbIMqkdccdiDk6GneDRtzK99qHXxxCaJxTlHAk
kbWNWMj1n7NoqHDuwJf1cqko5WxjegFsj3+6zOwze6Ua9NIGTDE8q36he7C5u0nJ
aDtJmHGxQHpfZsAxsDh+KTVTAS/IBCCrl1ziexnB4rCaRM5bgtJ8Wo0qRhu14ChL
8k1ReL600pl938dH90ZOBg4UAgS4+TEFuLfr3diAG9YUrFLshv3b5UU2bvM37RPZ
Z11Mko4DLt95USR4ulh0C6bMbsb/Whuo+5iuNgD3UAuk6dbAopYGmwsbSF+Hn4wc
yb3yIRt3T9U/M6ECDV92yid6Hy911orm6EhB9n+uyUyXe/EodqWeui+a4UZdtth4
qjcp2ozip8qLaRpBoiVDWBkMgXDMa2yvDp8siWMwbra3X16X1vqxcni6usqGu9xL
bhXOxFUcxfb487XRob9KVE9jac/sTg7JyVVtPQyT7dkWss+KodTL/1vhNsja4QZ5
XK5wHD05XAQsNDDS7efAIOnHzNSu/mlJMRY5FgXuxm0oDSjutMQAk/uTVi1GPDaL
5rWlQFHQQlxn1EZuRJhsXFArvrJ7BZt2OjSjaHGMR0/+y5o8vckyI6IA1plebfsl
K5ADGLYllUDhXVRp8qR0qS+KgAZ8GumnY/MrbbtQqEOrNAkviQ74kN5LwvFdOgJ4
+psbWL/QRi9SzWXlJZ3xr0cmE9IeW9GsvoMiGQbsCLZNg5+M/tI8qUJZ6bTk+DgK
uV2WKel9yMI9iUph2y86cEqo27Gc1lrky7XMrI48BaKsVuE/aTPzHhB0xPzk7Vqe
cv67kRg5krJBx1uCJa0HhIxZyVL7hVhVKKiiRgeaXrlwnC3JlJDXxVoJ95+zIp+t
LfJ4TMMThzR0REGduG+xiiHum/UilcIetG3FZJQ4QShVTa3+MuP85aclkjx3Um8L
DnIe+GZZLtowurxQ3jnMxh2cmWIXjOW0cwyddgnCPM+CH3vjn8V7vtFgl0BrbdYt
4swbjvd89RRHyttx9cnbbIOu8XasTu5SUqeHaaGndg8m/MwzmARhLIxuseDDku4l
VPEmDoZPeGns2ixKrAUiRBPoQydBHeKujQmEIlkKiwrXxMonA9o4l6nFB1WnIv6E
`protect END_PROTECTED
