`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S+fOYyF4yTnyIOEIZWnhVixDJZrJhqcU9WF61K12E6DS+KhKyFLSE5MuCzDQJg/G
XGeME+RJBo9pRyeoGPes34LHiP+L3wiYLweSrxFkSR2DQoN+hxizBESt92/gGzyP
9d5kCque8bx35d5cY471S2qZ4Wb2143DbC4gc1CaC5h4M5Uk0WA/gIFzjTiRJ3Ve
vSABhoO9SUa+aonWhw9B9T4kwLGadOPmLd7dyf9r6JGVXOO0CjSnmJgCoCmF4Aam
8KT7yjcxy/xf8a7bENzvIfxY3OWOi1MjUr3BOp7nbmMjnC9+uw+CETLiZWp8k5AS
Bi20h5OWtQHknZliiGNLmkBCnsMycHMDGaK1G5G4QEpW/fs79Aw3NsE8xI48rGNf
iRUxBTMKOqltC2P54sBSfF1d+IsiIeBsSybchR7otMN3vq+ACNCLUArQ3NR9Xqsu
OYTD4Bay1d9DasNDXU4FxHN4Hei0p8XO+JCAiOY6Egc6pUDsODEa8uf0YyJSTr3H
`protect END_PROTECTED
