`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1OvQSoF5kZK5Po7uomZPTTB6himTLYq8L6JZ+xvwXr0RwZg/YcRTWtlMNxWSLdo0
XuwhOto90o9NfVVEMXLXXgIBTks88oTAQpMXJV0r1I9fwvQZqau5LxtV36HWVOHD
Sb+f6IRVemRKT9Z1ocUlon+Bl1xJvoVN3OuBRHbAadGn3bxfOb/sM8xxfyg+apR5
mtfydAleAKGwqUsyNyu8Nm/cYLRJnmbFU6LqlLxRbNhsRyDqxxa0oM3E27tlvbBH
ncgkP+I67bLYBUxM9X8gz1+11Zt6M6llF+Q/vx172M7XFZjR1vJ7yu6QmdIY0V6H
/fKQl28RusZkYL3+OOs+9IEi2SiXzz3xTX/zsj8kqMXT7XXMdjKLg/B3To8lsPRD
b2N3XRF5qEHYBtWBkBNXcF1qw293/z76IuzvVAVAetZaAhPW4Ac59GAMUqKid3RP
bYm6v8GTSMZs+pFZT8v2ukggR11J1tilr97kjyJZBR71MxprkJU9LRFhaQl9e/78
61iMa/eda5uv6ZzvMB6BhbggMKIkf9KTBcYi1+MyVmMCqlp6TmqSYhVV7B/Vn4UV
RXoqBWPz6JdyqSHRNmBa2Q==
`protect END_PROTECTED
