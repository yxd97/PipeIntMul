`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JdTCSh8+hhTglBdbMU8ArI8+g5do4+w4uEiDv4HWlgRNOwJBztZBC5NVW9RA0cCu
OhSppZsnUmOxI1eWgEdSHpnrMxL7TuOT+2Jix3PcNE4mea8jHAGnEkpL5MZ0yHsc
jzIQDgke7ncEsqcitaZys7oaR/oDwoVr8Fi4gxaF6s5UA+fNp3VN6MsceGSTHQHz
/GvZAnmx5pqLvHAkdjm5jOrR4ZHvgYSuSDBvI7mhOymFUWArXs60l525Fd4Ab9Av
pzj7/6YiryRv36QjdPimIjhOo+j/2UXG1OpUOnqlV02EbrcJJ9NsWvQ6vvswPQy+
mSQqjvDNXyL+UoeNiCK0GWSI3QZT3n1rVdR+cnclj3LyxCi81KDG2/PZTwYhU9zq
b6Lqf1g+hwnTdQCYbV9+eyQBnn8UGjmpN4H67XOKIsdGx+XLO3oDYhnoZDqlc3K3
JSdPOlH6GeKzOcg89cJoDnHSOf4LGkrP4th0odO5gHO3xiQJgjiN4d84LgeTVgX9
`protect END_PROTECTED
