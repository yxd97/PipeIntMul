`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxvFF3MunHrukssGaCd32DhIokIpQAZOm7sjsVQCwMA4t2CK7i7Uc9gS3j7Tiy/l
m5jdNG6ECR9bIVHe8jBojcRrmXX7u5+LFIPa7eo23DymZGbsIb6EVZQs2ldJ59+0
uuJ2FVtPIJv/P9kUDU8+f15n5OmO7ps4bqza+eCbgOuKWGQekZ/zx36G0hE3eWdT
T767rUMNaXDA8cCZcLTL9pZkML4SOGTi5zypKxhQQhRsnqHeIFdegTIsMMUtXJ+k
xEHYRMGo7ZmZbPJfmAXi2hJrc5b1DVn/POeT7Nnaz7hGhlLaV+DQti9s3Fb0RHCz
8vwpPcgu2qBH2zG19P2TQJfy5ltzJ6PikTYcEWGRKtdQWg1HTkqd9I0SOJm0rB0f
`protect END_PROTECTED
