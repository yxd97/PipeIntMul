`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w8cf5kv5/5qANErgWJA/yHjvXKjpCjEaRV6hZHq3Ut2S+pKJkOdLk/LSA4KDnUjd
nJJOf054QhpXwWeMOXsrPQB9lUu/t9DtAXe824EaEkgKn/pM7piKslF6ucoRbJIr
s+M+zddavIT8dm9E1PEh3JeLLxJT9nEOkEL328CUV1BKIxI2s8FdtwAuVZSMrv+U
qRBs827VQ1inmF+riCW3mFIj/AzACidO7g+1ltPrVhXVQCvlgHM5LtV3ZYCAMTiR
Y2X0S1pTvdkBUJL4VG6gb81zdWzoCBsMh/imfVZsNVD9zLJJbjLvyoE/W3uORlu1
8QrBxrqkRZThPI8SYLwBWJbUUF2WVcBUMPMvsb/B5Hiyxe23ESPovxNVA7EuT6BD
aCo+tK1+5/u8BXEWKb1DLcJEp3IF43swF7EKSmXwpjA=
`protect END_PROTECTED
