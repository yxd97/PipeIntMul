`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Osd6KUQ/5jC/1ryF9z89FQNy4IXSFVl4azosmPxPMDZTeyfsr6l0/jz5EM5xjEq3
6eFowUY0YKlcWzB+UoCdfxnDowFg0qtI+cmUQv37BDucAThB0QVbHBpYdxjBnRc3
On60kAmVR725/902d7TEIhXckr/AVULf67RGh3X3u7aEDUEc/9/PZeAsvKhfGyTh
1rJsL8TwYqTDgYUJ+vNn4nsUTiyOomSz4TpEB5GzGLDfjW0agAw1Hmw/uFubmA4+
Oeug/HfebRJaiYqt2D4FkbT9F8GKdUyJQXUVpbGL7wb+F8XO3Ud3EKG1lLn2shJc
IjYhNOpHbYkynLoPEA/dsfKsqMuLBZVw78WAEdLku8m66GEUULE6w8H2C9jPsh3u
Bi2BQJnpYA2QjGldxFVt66sz/ZIEu4Jnq0L0HnfdsV1Luzo+z2+Y1X4HQUTfyJmO
PccYh7F+9cjOtzdp0lbL/QxY12MMhCctFwGBEIRPuaddQbPVrsaDwlCkXosEhPp5
Xo/KfOa4yoJc4pqfZElTbVrax8YadjYqleTFZfC31FI=
`protect END_PROTECTED
