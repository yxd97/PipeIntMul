`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fn73VVqcOiz7RB1mSerBEfLl1UAb4YW2dLvZMhpEb1hYIyhy6H5mv9onaOdNFSVK
c6DthdPDS7s2HNiPde1lDQfA1aYz4i+5k0TUvEutfriz3xSR2/Tx2azQ6HRjH5M+
EQq1mgXBPwH+a6tZGbwMVtixuW91w+eoQY8vcrad7x1alvIvtmWIVu+j/+fPitzX
8SGaFkF1ocFM2qGmEJ4kJD6hkH5MAIxhOnJLdujrwP4uD/0gJ0VQPkJjAI4AAwBq
qDaYB0q8g/MpXc//uQYHPrRb+5EW4nSjCB0J0J4W3LLiBeTOXSrDcHwdY8s0/ByU
pLwHQRvSoklD9ruvYPTPE+zl1FJ28aQ5Fb+4bPxskhBLLLbDoAjnXf1UIGadfBz3
TnN/RcRGxq81Iuw0sI8JkC1Ru9vMy6VeFhwqdsYBIJsw+aPtWpwkB1yKu6LXyJ2n
1XWSVeizhee3eat1cHLAoWOxuyvMEZlsHiv1ccPHfyVUUiqYp+Lz7KOPce5qO5+H
g9RuUff0MQf13pambOe8tFUnsvBemBqv3Ig8N5sw2zi3deK1PLwrnjrbLKp9SGoE
7EwQcR1hMeal7YRCRaO4FOxF5/QpIcuDoaSsgaQSlML8dEk3Bh9A0JL+/yDrbUO9
SMN5eqt+v2uQKTCdNM75IMV/eAvKg5KZXMIKRFUIT+5FNAtLn6+kItySm4RA2Eqz
rBNYsII0Gp4E6NN/ERu0BF7vKqYYxHpxFZoTKng114HXdNyxckuKEpSvApEU6QAV
dJijfywTehBnUjb/5P8xiGTCyiy6OUMdNcuJDtL8kt8UwRcJkyjQ9Z6gqXyv7BNf
7OxyYfY4xkzsp9/7+Y9H9Rb/CIbcxdLC+x+9OS4+4a4NT2M1x+p7fZ7/61/M9ble
i49gKj2XRh6eIUvrNBa7IG5lYT+hW699ozAPhiR90AMTzD5XpugwZWU9E73gJnSY
UQOesO43oAndH1r0QFt+EfPp0dEjNiZVCu1m/lDOieJbbiCTfrTsCINzPgu+AwQw
KEnDDxsDiC31dhcfa07tiAICz5DmRA6L6qLQweA/rRpDL/EJiPuk1dQULmmFBHAG
Skb27z/PJ8RDMi3q7U3OeIrZiUkKS9W2pdF6G21GiHYwEw7px5FodPbGSff4J3YB
RVPadZXMD9n3p7YB7G5y8OEU0uxoTR3I70zm7ROGWqLrKX884gSgrbrJuybW3hf5
qILw9watndrZRqD+NDvy3xAcwS93nva7QCiJML2VsRdW59JEeqCxN+KdDyx484ez
fn6z8NJJ/sfhmSONlpXTMg==
`protect END_PROTECTED
