`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0vSC/xZ0Yt8CBG/LRvZwo/9h1F3OEcW6WeUzy3diRHtiaqptkJBFB5V47gDaaG7w
6eDDjmCylKzOPyix9BtYJUhcDIPUC8b+sRw1AMwZDCWKdoBEgZobCgq/AHqyg5OO
hM0WwhmTj6XR1ZrQvPYvgec/p+PPUElrFTWfSkTQuqKt+TxNKozl33LDEU0/LmEh
RXpcUb8Hvi4K8qLMLhZkmG87gp5XB0XygfveAVL/o9n1qwKL30k2etqDb3rVskWJ
3CW/R/nDYIrre73QTqGlwS9bgtKpH5g12E61hfZUYmNNi9kx5L1ovLR07r6N4laJ
`protect END_PROTECTED
