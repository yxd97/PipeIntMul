`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WN2Wio+OkCmtj9HgrKbd6P99Crysam8Cme0oGlqq68+nafiQRqQ7AmA3zEGvxDqk
W4O1ZO7yiccp3ybXABz+9Yt/6Q71dWoXdvHEYVJSBtDhiytX6QjgMCRO/YiIcvIU
Olb5/eebs2l+4JE+bWy7DyS/nDGpIitrOXkSTznzltS4FB+R1Xmm3ZUrHgLOGL9b
/1ANX2QoVi+U7nkg+JZkJ5jXXNrDEGFjw3knkxSWYyiSLysiiC1CElb5zm5fo0RF
YGbeEYBDcS0R4ikwnzPLhINV6fCfoVZMv7tYNwM1lx6PqQ1Du+pAqgdHPAKFvnfo
Lv7IuzCblNXfmqmJkt9cwpl+i3LqAZKLEulhCHshPePsJiSG3VoA8VAa0mLwxh9M
GvRu5cy9rpQSfDATJMD1PS0vSE+hZbksvD41NV8Sheq6RRfdVDXiXHvMuf1Fzkyu
M9M9GChrBcmZKict9aXwRMOHWuROtCC68dTYtY34E4nQl5bYcOopN9KqCCayFFwh
/AzIR6sGHcTBqeTYpRPtlI5Y8VuvGX/BxmMQxYzwgUBSFncfBpJfeOgrjcLGKJWL
bix2pdnPkTOtl0bZ6lzhpnK406p8rrhUrFh2OQAlGpqwQDU8zA0THL6fHV/QF0A3
M929Y6alM3qx1XP0UsWW05XKRBua4Vbfh5jUVrD58FRvY+eB5ie/WS5mlVisWxsR
L6VFx4jVMSqq0DGxIAExoALfL8o5Enm0RI/2ZvjUEXPiirN9deS58JQrZdcH+Zi5
Iuq6j2w2MG2fye89qCplqQuwre57hLR4YbzXiKpzBwZcUY3G2XjMzwcN7Ld8b2U8
ZY8S02pHbddpGk2zOn43x9Uh8xA+OBkMel7Tsdoxc2uw82WfksPaDyQmLawxyONm
LWSaLpa05lnJNPTqLa853F+vWS8T5oIuObRdtw61lWQr7MhygEmOWziFhICjZdry
qxIYLHS2Lqsfl9XLt4cNYM4EMmBKXsvgRZ22Q7XXXqZQL4EG9xZKeOpzqGkF8z96
nIqfyls9f+AHIcuu2hiMpw==
`protect END_PROTECTED
