`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V0YInYyoSZ/AMIcz/iJljD3Cbx7x/s7TZ+0O9mTFTrUUGNp9UF2PmTxZrrtu9HRZ
LE3O/TLO2uuCKwsEYn0Oa994qpCC7PZKaOfRoCh8dsQhWvJRX2BBf3JPsIhwiAdR
7iMEYflSg3Sr4DL2PPPoyKArJzNiEWBXViKK0eyPr78uhDKy44r5QQyD35HFccuR
XjwB0UBkgarfeRIrurS4yw8bjtW/q7dR0NCoxQ2tlno9mlXp59xwqrreeKEks0b2
p69Swg2B/LuW/8DfU8mBPu/S2e5J/QicbS9nljwgt1z8efI/NAlvjXKFvLeFItfk
+eWKEV07BjyQ6lZ2VY64biV9nmZ08aDD0nFbg53yeLJHz06edO8uRwbwrHNi9p09
G7u2ti4+zcBlBksHvBjtoWugnbM3Lo9/5FBgE5gcAfyWhOajb3hvKaGZRoelY7pP
WyKKX0zLheHK8SNrNMVBhDz4KXevlHVfoSqfIzbFjwK/648f9fKRgilDWTSyICti
Jr3JbCYr1TuhFtG4cuB4WETlOdyu8elB7F2R3dWXk7OTVEJsNs506bUbEZzU1ucV
YiXOSg0IUo6Z0zXmahaONKL0DkB5HkQRBq2z4evjFfgmgC0rzU4zobkHqoxsbady
FEHo4f4eERdI1KMlR0hWHAKjtScaNesakyE67eP4b1HncCWebFmHhjyB19KkLyaC
+ABTV6oeyZIicBUMj5+pGGcpGx8V73SvOivfd1M0gzzlL0AC2GaZHOjGxz8qemFB
/kF6TENoF+OEBNgT3hPwlywdMuDuy9T6c0Wh1XCBcC/aBuPBULHx2kw3ATG1UQLn
byosiuF2FN3WGyZlPt7LRUMCDAkeZZtdMhWqEvSKsYqJWwRGxwBS/DrZfQUXvPVE
nS4pkDTp0hj0mF3UH0kXg5tVcTzLtcgogIbCa1JE+e1ZNi6o7ul/a6N4fwD/Snmo
n2ePxZ2aGg7LefKzyM9FbReEMhkGYNdXjg2Po1r9HFnOO0uUrM3ed43Ah7YWd0uu
PxfzyCk/YRxh1qu1EvYpm9giwZ/yG+Bfk3kFDeyo8kA2xUEzTlZq81r6QwFt51Wc
mMIFvjhiHFqTO3wpyAF8Rsh07/zsEVTsXgKRAM3+G671OKyVjpCSq0d/13pMVyOy
LraSd8LzxFsyEYRBV9gP4miPYJKaGEtyZS5MT0cvrph582bkQiaV5NuQvlG/vC2h
LyPK3DOFKR1R2xucAlD7bulk20DGuZxmEPQGjHHiaK3UEpEWbq73fH41k21zwqv+
hrPgbqhtI+9GB9pJsBHEWSv1at6fJFGayIXKKCp6IwchDeugtSpNIuY6W/MwSmWS
R6TAw5o0QB1+D2Pt/S7L04PTkfGZ69A39ND9htBF2VshhW3xMUH2e8YZH/8qy90s
w5g+xiqM1qXwdSv3//dyKkH3FzG5VHT5aBGQkz0JG7mLjhcxHLISd4FKVWdltj6F
b6ItDqFKzm+uJuZ/ur7hMwHqsWMvlC0IVmwwIuYR0JiWymE9YSxqhkLnO1mJE0La
BSmgbYg4e20Pd+YUmS40zR7aUIzpc4hx9D9MonU1TIkpPt5SnKWaa2TxTaFhN8aw
82qk+TSgeiGltaZNztmveQnDEyrDXV5P7CrrgvJb5H7qgvEkY11Y6T/b+SgNbRxH
7zdNcW0+qOeYIUmeEvtiLZ00VPH6wJ1aHkvJsD3/m4binRCadho+b3R2VhqsQt34
mH2skVZjPSSFK+pWyWaVTlly5/dhO7L7MPak04hFPxuOCqcNdKnYrH7DrZuvsWKh
NqQ/ApMx6kXDd5O7X6Eie6z86Fp5l7sjtN8wkr9gKLv/DNPZijQFGJAq+qhCYK/l
kPcfptxgMkqPXnIDCzK4WIv0PFwCeHoIHXfUkpzuaqC2t7LNbabvK2NCBA8Enaw4
pJwf/S+Mhoev3NtHH9VTqISO30uZqq5CHqSh4C72uFpTyp9fJxzdIzQptlTUzbU+
l32m2TUDJGJXBWCi1gLge2z6v5gGwIIr96E++AzE2TP8dWBl/hLGPjAuhUtb69sE
K7p8QKObKdck2rNwS2xLRqZidHzndAAh5wLGLIqp3yFr/VRxEpNRq1v5RNcdok1z
YtvF+jY65sF2RqFYftQZ64zvJZqxFSh2tKfZiEEqjyv3BH86lCTlNkcQ3HEmr9bb
yhg/YwT3wuy0irnRJR0qmjmgRvB6oaoBOiMwzyszRdIDuJS21aaZav/pnR7yrZnH
5wI7/Y0O+MPvV716xcka/qTW+dM7xPbQfhK2gTCHsQyTcaeQ56e/GyawvcbKd47+
DWF7UEW5pRU2o2GRo0nWvFx7+jRPJ2pN5p0ua+8pqWM4hzqM40oQQf/8pCeREX4k
jJ3pH3qd+GfD66k0WJ7hm7LYrpIldZeVbnFMidY3BzTFWofjjfrjZXvVlOBasz7R
g3oXrHD3aCbDs1icRJSu0/vyb9Jz/9Y31HuDexBUdmKTOlZ7Qs7FN0WyoQO1hQxl
OAslAh+RNpvtcWB5VI09wjJ7PTjSkgbP4v5QcOso2OwQG/IlBgAfHfz5w/qKp4xY
AwCesWXip4ep6POMwVxBpA99CsZd1ZzgdrOdwJglcx4oKrEP0R1FIKO27tgSU6Qp
pMvhDE7epl0RTQfrYwWOteDfHsw1aZfnZL5fN3QRQJy1EdLetUXStncQXKgHXwdW
EtfWU36nzcZev/Nqz9nnuKClMltshSaWcjZpSDDfRYUFG+v+UN8Bk2tuWmmQqm2b
YsGuX+q8mdTB+eeP3DfprIn1IG8knhgQma7RT90NV1u1+sTUTpsFe+JXsbegzgQ3
RqjhxLLchATc85HaoPxB82yGqupzPeyowtEvtG+UF0Cv45o4/n//OjqZ+iSXZcD3
Ih3ovdDKqoqyPSAkHNjU9H1TwqyoMKWiqy/qTC60FgAmXxTi6a/nCsHNnYx+aQiV
Yr1Ga0PbxjXTiploj2p4XQVrGOCH/jpkshha5PfXzmwpkU+cgu/MZHXXYyQrQGNL
Xc1uoXlU1hFeVak4YPTL8nR8Dq8Dx8Hbpx9oSbgyFaTC+mnFB8ctWvDYXxmgUxs6
X5/Uyi3qvDvLCN2B613xqoSra8krhgs7uegrt82C1jo2oxHLy3TDfdy/v/vAjHwR
mLixaWW3H6lnzzqkm+aZl89o2kz9+e0dzqkUBUuFSgs3o9lssHcSd88Uua6/vhLn
1k74LWUZij3mAfMFb5R6BIvgLlCrlXZNyzPpzXv6R9vO32G6hB1el1W9JL4VGJh0
jkUJ+vHfi8Q8vq5XDSY+XwoKMMHD9g3b9WBQd9C2Di07jUROkf0Yvyb2ou+D43K4
9zAtS74fYMWn2yzSbCVu4hFfhSwvKVx9hoR3vAzimjhjqhgr5ZjCFK4XfcDVMkvQ
UpyC4/RTY1wRAWfnvxCHc2DeRvP1ffE8nraQD4K1aY4P9hTKBBEKwJYMDghIJqMr
QF13U63BT0xB2WwgNQiRwbo5+TzjUr9AEd+pNMPAbVaxZdeWhn7KbzbJXdSS0TWS
xmirzGw2JtkEGDrZwOBXT/ET3gQNnKzojVlWZPzgnyz1hTho5ktuyC6QWpD1XXyn
oR7qiT3CWdAXy4rSs3IafUaZEXEi9d17gCLUM/IJWVgfuR3g7SIyo41ADsmowkYM
gvvBYH30hhIOyRHRw1GGDxIxVac3MGsBKORCvc5XdPfvp+guG9fpE3GtDeEnS2JJ
PqKHBXJ23mfkc0VHPM4Bg30OJpJB1gidtR58GO+G8+19+BqQAQrvs+1pN4K/7m5u
o4fn+FmFsE6zRDUgmprxz8WYZWDDZ2mEmlv7pLWNwU78eR07XmGYr+dvGoTQ968I
DpsiUlAc0sylnjon6uakfb0mI8Lr6r16sTarBLa/zZpWWHtNFKS2t/QJtpAqZd7U
VjtyncmAv/YruhjPEvvG2Uaz3OFoaKLNBnuTGjGuhRIdeNhQdP/D5G0iyRDe286f
/iJroiBJWpqslhHQ8c/vxu2yNfw0GVqhOwO8riLkVtsOwN8eMD3LaiHyiPIMQlC8
aq3Hj3N6v+WPwUgb3ORf1AhPK8cDHCZM44RTvup0xsl6RcNwp0A3XOlQCNUF0ze8
uBHePuI5RIQwvt8xNHvTAp/ztNxeJZSgqQ/Xx8PWZLkA1cIpbnretYr13R6vEEUy
mKCzTpWFQWTxmKMXa5uPRzoIkfaC5to22jFZtUT6h/fUh6z78UQ1NL0tBTfd1Qvj
Aw/PM5UCtjPIi8//GQb2UHyBJMnF247rtBFG7UWTLX0m4E6mhNeySsfdZair/e7A
Ah3y88wr5lFXXzI0PoQhXEeO9Hta2bcCEUsUxv+7pDRfT7nQpK24QlTtLOekIFFG
PYgTxD2S3/6XZ3Q5DGAbFG4hQIjg7zyvooevMG5icolA4hvWbWbEKRTl11JKoRGs
/0M/5ofy4QAcMpIFYQZsOLDgRG8OpEpVJn9RnMQfDcdHA9rMTebyF3vPOAprcTBa
SwgfBOFheRwLTFuK8+/bVEXoDQQw1pzkXwx9PypDg/jstcWS9pL3EuYq3JfISFpj
O4bQHaDqTbuJuk31e56daxrLdY9xy386wUV851C7VMHwInkIwyjhPYK7ZNtf8xL3
YXnUY2lO9QwyC4Vh12P4tLwvGCWb0dxJLuEweLu6uBxGGWfwuQgYobacerpnnswi
E5dlklVtz+uK3OuV5bH7gYiB2FBbOBDQPIFcR4Ieqz2wckzDSeYMjPHRyVe2RHAU
0PHHORdh2r+KMjJpHwidi0GZB7kb9q1000RiLGYvn8dWvXWbPns81Y0fh60JkenW
/11LrYbyqwDkVzv20Btmue6fNOTufMfOf2mwuZZntr4YXYGkfoSNhwBDElNret71
oDftAdpQNG0nLwKr6EA/6Uo7k8IgnDcMyMIdSGjIwxT3KzscUYN4kTYFD2tuQ1vR
NEp/WPI5Eo5fO/Zz0RmOtL2tL8Zf9FPZZEfWMAfDds9oZjBIjN/aEJ/w/b5QsKsp
UwuYsnk3uInq2kk9zxYP8BFanF6B3P+/AINxlI1N++tsGzpkr/u/9aFL/dVY5nhZ
8o+cBkuvZzCT5EqVLPxeNY8DpD7yP2s9SnJUNp2FvkoWBAT4WHERx8HCt64lNjis
7O4I9zLvucBTF/Y5Kcvo//rmIsKWQpSouuxzYfUSQGgibDhftfZUzkuLMbmrq/n3
N0r7eJgeG/nCG6pDFsxlfX7lZri7KYqLL+0/5Xb26qPAzVWhk+IwX/Y0FNapZ4+k
4kJwiHJ0oCw5DopvKtRiUAg+PpNn7IOHAFoFZsQe8YLeGEOn0Q9ltCk4XsQ4jwcS
oylEY9/v4eyqw34DhF5EtTsjIhFmGIRePycUI5HizAilpRk2nSNfO1J5OZy1IjDp
0qEL3s0lzLEtCndWD9INNgLHYLdwkF/ogKrvkkZ8o8cXhcxtPZRpeMVVqZicmlm0
ekbJl0o2GYlvubLYSqSq8r49UULdtGkrVL2S0/xTHWLS+awixOQEQllBmi8GMwrX
FEHgcIOQzbibzE/f5M5ndUU8d60nn5coLjKJARoFCAM3fV2OzlzrvchQ/0/4pDlH
Rj28MtoB6OV2i6NjikNYUsANyTsxHJ2bowB+6G+SkdxKdUaT71rr1dNvAhdLaaVw
p205erXRlaixXo5mYDPfmwVoEAJ/Dq3Z0ehaazg5nLSvgqSyfOhFAU6kvDa56XP0
xr6WX9c/ZeqZS0afetGEzADBHWlS+HKcxvKCuWqfOQmdfE8ku8w5qRZgzye5vMo3
0m0ceaW0E5a6FK2TY+SSEWHex/DvgAV2EeZvLo1dPkPgRPw74Lmc1xrHVtMMKKwv
2XbO9vahppXoQOPQlymB5GZMnFhew1Vr4koxe6z7CzYBa/l0ITEll2AYmgLwH5uV
mpjxBQY0FXT4dK9ElaDF2g0gwJ+xKhw9VzD3eJf/82u/BBBgrQjYq1MpupyU9f6f
HK4sLj01dtl5X6zEMqklqi+DKKqDg8e3ri0tTVdkLnwk0Odh/l75v0jVV1tHhTnK
lmLkLhG6lTICyXN2qGkFoSjLQkDWTNmEr9/lGpCXJYzUow8KhCXlARxswFs0chib
F9L5W/VmmEeg77qSgsK/uYbkd/dcptGIUCKB8gWvnxumbmJtl4oHP5Z3KeI/tN4t
IcG7xycUGYJ3+c5WLX90EHzQJM19195CKL1rGrtEyE1AHNHGYSBHSRxrYLCkwAk6
UX4dSEiWwMimTShW6edWH/rk1u07ldGLZcLNAZ1H3xUlaHj0MGmh06UlaRI6q1Yz
stI0fuxRia/9COj48wxmlJEw8JRBFvtyWe97MVrq+U/+0ZtN3cMG3TlyCoGvjKel
Qp9jkoGUwR0Rr/P50euujvmzjve3pFW+OcOlXrnWQK8/6cmhgubXlmffCgg3l/uG
HAEQLpnU7sBDbOGmnwEsDAsXcHNVoU4WiTp4eF6txDmK5FXwqwvbxzV0+CsQSyc2
FGCDno7qdinGeeE8kJab4bs3hDzWMgz/nAbcr9lHfKe23sSxwzOTbK1Tbj6cmVUc
bQYkfB3oi0+wyUSMIMf3Pl4I44MrGBYJXm9o+uMbr1E7HXtZ/aMC0mSknF3RdUEY
Y5wS8nDJ/OlvN9l40/++iJj+cnXV2iKe30NYkYGsRdN50GL/XM0HjyETrUw+PCN4
IvOI174bihF3tFS34H/EyVCHp+1PmXq4YFctZIdWNeXb94UwqewvFFfhEEGSldUX
OLOGXkQA/LOIFWbQKyO0hbj2QIwX25gdkayvAtQUUBraoGxFW9LIXshQbmt3C3Bp
AU/2ep7f8L5rva+eLecNzWr5kjq/Cud1mC2IaVXoid1vt8ixno/xcayJpd78A7n9
GQvA8C1bJvqnJ550gzPR9VFRw2MvwPKSI+57JKO44pg6+yz/P/JJEyzaEzKrJAXF
7cvXgfZt3lwlniyJkpYRBoa67XIJCv62rfFDFkDa6qBq6HvhhNoE/CmklmUP87TM
ECb1EWbxPZL60fpeVxk6eHVUWxHWnih6pReWInghpAwnWAyolFgaPrNdVXn0/5Z4
G1j5KWfMEo6wG0zEdus/n+JpVYN2Ph/2CDdjN+rkqrRHHfJFyEerjMIK+XUgMVLE
+DupgwLWmYZut78ofjejanF6MwXeevj/gW3NpOzArBIGfUCBwamSZMt46ZUn5zfQ
fo91TOQEAqqWSkHSOq6j54I7vWhVyROSfRMTstpBW9zmEA3Bpd2h1RqB+VbgaM9J
O6TleSvbyDf2NRIqH6dxbJftAAddCOJCVFKP/6Pg2YdFA/R3KniddR6kWVhR1IaG
pn9GL5FDpu3ALhA8WW87I+y3l2rGwEGZmxfYFsno7QaehewNqlO4fR396/aw3j0F
862hjZOcE4/LCFwTHj/LYafOL5zejuUMhwcIWn8c8QiMLFDkg4nLLT/lL3xKi+K7
4J7oDmz7vn/ec/SmVpsIyEXpfWjT1cXw1kHX3kZIzlWKPBqqS7MFhT/GWwZUOYh1
zS4z2UkUDFMKlQIC3q1ARCTyjIA1Qe5JlN7LVebBhabHdrGHpoMYkeucUVeSnmjX
ZJT0gZo+pkflEfg95/wFAbnyIY7KxXql0w9wfBhyWv1pfZFNVC+uduSsmmSBWUaJ
w38w+LVOqRaAshLsjjPZDzepyRfTqOCIPqmXQv6BJoGMAR3LgL9615qKM2S8ymlh
nycn7nAx243VSNSv+ycVzc2zSK2IrjsqzTSq2NaBMr+BSJeHG1ogu7XD4ClyxoN9
ZIl5goHvkqk6NSeDVCBp8IsxJbfkTuFHtRqmuO2mVz1iCUaVUCzO2WDaOLfw7O5D
sYAuBUqe2v05Kzp+nJQrggTKBTqIiz7e0MOnQI4ppRCCGlGXcNn09CJxyDehaK0G
LzjYT5MJLyXDQIhN0M5YvWTjU6qyaxmoQrY8JA56JZ3cIIseymS9yIC6je86auhU
5jCukyOkTNTC5PI6iAtOStJeVjV7HbOjjPTqteGlJejYK2JVKePjBP4x5iVNwmRU
1F0UpGY83AwpjnXD0PlOD7MTGORnhRxmAnqlkCV0twj+Nz6KaqEpbhLzAMYk4hBG
K2rzCbl6XagMgRn/o5NzWwxcedYzZCxBk0oH/9WKoCl2FWRNSh5mw8NU1PGRsswn
tfZyv916KXJ7pgnAybF6WWNJWRWbFteh5Euz40WpVijfHjz1vl3cUDtNs4XEDsvR
UFWFFh7RoUSo5rPXj+rcHK5SV/ZDcqCHgVayPKKtbEjfm4nJLWkl/yGlOE752lAR
/8HGohlxB0BC8gZbkTw99MtSsGLwP8RdVUdv7J+ThjcWi0ZtCAs6PN+bzLPed+ve
2PsJx29MxwX1QabxxN7IzKO90gsicI7Hp0U3H8ly80Z/drlo7QRce9YxJmdKbxUw
2jt8pjU4bhYMGkAOecmJf4LSdWpOGDlRNevCD1nIFjAhPTTOp7IkK1CBcPDes9HY
cUf9j1S81trA5uv4S9UOey2zsmvmxmPTDng+t84/f1kCi2gmOv+prC78fjj6aScl
eg7MqyepB77xmlGB96/dmxpxbmiusbxBDg6S6lGK/PwybvBPgc8qBNr8sILv15gE
BiUu7E4CBcG6y88Gpnufkf1oYiKPhx/Tm6SshV+owCSQAgIRBbjKlUqKdtqjxZEA
F2L1VQLUszeK+FAza4L2N4wZQJMbkO0uL+O/IwoybuiHQjq3TrNsoOVC/LHl69zk
qI5wtcMTMqDtegUWoOym/+aMiZOPr4u4EzJYVBC3F4PT/3BGmtflEIDVeUbWCx1Q
hPJTKDhTwykB/yZg84DPba7zpprNPiP+V3oihdu7HnFRpytJgx6RyQ+vuv0/BrRR
eBiYgVaw38jVwvfKVQusWZua9mMgKfl5s/ypMZ95vTBvq7CiBqHBoP65OTumi87j
s9ZvWXFZxbNbaXDX2zY/At+AZYfpwaeAF4YhW5031TsJoguFwpmPwSqWA59AW7Rb
D1cgiYUWDRVf6mkPEVKSL2b04Wz6JGQHDUhc6Lvt3l8Xm88ebsxXFxHQmiJKouvY
BWlVVBkR8TK8EgvA6Do8YRbUHEqBx6Sd8z1d20XskuXpcKjHHZm4BjS5l8uUqFVf
d3b2A+9+B6DcFbEXsmoXybhjVNGPJ352+RwcNxnjL/8hKzyTbzpWDPkh3ZmrKLjg
XJHbD4Veugz+X+2D8hhV7YB52cuNdhY6Ihp9vLUjAcWq1Gv4SwphRsbZ/Tta8ZBu
GRpFa/2yYI6WAW/pncZbrepdqgdJZOU3nReIOMb/zWZpO+hASI9GpNcHHNdKEDOk
kxlUyIQdxZ+aTDXBvIQjv0g/DIBCaAMGx74UUbIf/2lLomuN/Gex/1eCxzi19L6R
XnybvgSkDkyX8sDJxlcYaQ6uY23J8IcW9POsO0NI4hU3+qMBqg+57eM6rH07Nmf6
7dCLnlh5WfxwdAXqgvh/6qE1nGBSIYsjCtNV00I4rJf4ze++iIeOar6k6NQTPMyf
TiFUqdv7UfALUbDt6s3IZmXsltAfLVZMUUSaVEqnDKkDj+LxxwSZ+poCQ5zNnzNO
awT0jj2vS6Semm71jau7/Droiqa8oiuIjb8BvNg5Vlh2i3KAh4k6XklfkAjue44F
yAa/4KJImnbbH8IfKahvk0RXLeujPsQTTuETfRbHN0Wx7UQkFBHO4qMkG84kiKFO
9vin7nJkeZZ7bYS/U5olTFw5TWu9PnWCvWmu1r8EFRZ1DQ6gTnVD6aq5xHSlcaiS
KFjz9vrD1Lf2JzsooKA8bSiWt14wncdGLHHuFSeZWu5UcQ4YEshiK0wwdGnSIcqQ
wks3l6rjQWNDenf4dYlQsJzHcntzXLfIgtOGeiJPwN1fWDwUjUl56KHYzkZDqVCH
oWN4jlEEMULiwP+jzusTEL1e+34eF1LrXGK0Ityk9/nthoyWhj4ub4+m4hlJBsdB
Xl47T0RCkOvOB7Poukzw78WV98mTBS5HEaidcKUHCBfkNBRrf9/C5ATBYd7MTPwJ
DKWqAbH5dyCoaC40oBvyI4KqodB3AGCojvns8ascKtHHFwb1YjDc7mvQzhdA5N8F
00lISOVCRBQwFFdB+euNhnxCKixrcT/SuUQWUzJvY97G0ia+sGd2nrCNoUziVnuL
OhrOkZE4ul+CDOJgVDbnPmzuvt+17lz/bdtj0e/5RlkcEHOBnCYdaRicGLX6iNUN
H2gKXMK+bRpfOAhnGJgoTMKzOwk8W3PgX2N13Hv7FhcPgOa2ZI+tpl97MoxWzwK8
G6JxFjOxuVVyOgwxNmMiRD+qYVGU/ZAbBgB2+JD8VsXQRi1oWNBjwaBz4E1TCFrb
mzt4ehRNz3eVaTcTzLs8Ul6nOvixuqNCyBw6SqV9dIVPe+OEAXsK0dYrJMP+Q/Eu
J/2WtVNqCVwLMyvTk0wWnio9yHP6UzVO/f8V/0b1s9qHEUaTeRMwxM+QnjAn8hUP
9V4IFrcYpfF0lLyNQ62Wo/fo6DnZRGQAUbCqWVs3BeHD64Msa4AevCgMlFkjxSvN
zuIkDqdgYXyGZM6B71Sxajx4ukTZ7DK61+lfU3x9iyd5yzNWAEHuIaUf8SGQZP/e
1SKQi+n69QxZp/5GuOvgHMVgQN1zYRZzHNWEeuZmUjcVeMrHkMQMpdGkGBkP1ZVe
ZgmWWsFXJN7j25Ow03SUByw854OrH/IIUWzOZHNhD/aUJ1TuQ+tzXeDzH/8WgcPu
LIVPBOEWw+huLNZsHCbrL40XQnZrDV5YTBfka97IztcpusEA3iO2ZeDnx5nEUTtB
6SBk6cM94evUwD9wdKc9Jqc4m4f8W/ncG4cp0Jw743SqoCb5zvUAqOTvDTIuNIsY
AQCzqR/I9otfQE+Q22/Imm7KNcPvyt+uIoysaCBnBPN7bPzcdKpvKBgUthviNOWe
llvCn7Aeow1+ryuUeNsrhPNirib5q/cvpfZ0IWJdGTGmOTmDcdGqJTSXzTh17ftQ
SwkpbtVuaXZnfSP63vZthj0GhrPu/uvRQqeiYkOxr8VuaIuF5FoffAewq6y5Xqee
SIK3Lf5cN173NoRjU8WgCjun3AAsUXRTQ1LxXkoNReVo2gkTXxTEjvC8/9D6Xzey
lKb8reIxNvFRddaCm/e4AVRgStfNX4KbMxbkBtJYO6CH5zm7EcstGFpulV887ESt
vvGrz3iVsterPFMD1PfFX7paOe7/jaVJH7JCNa9NaNbCB92lU8Z+qWqrbnwkK9cR
S9b8SqKnInwp2M5IM5kM9+TExh4aufVDbr95yNcXxgLn+rbeMNNe0HlWF3N4+kFc
TilvQpzEFfglfdFSJdMjNBw0QvMZcUdFWh8pRdf1qXrs/bSsyLEd5RCyYHETjPTj
QJhT/bg+mOQM6wxy+/cv3bMv0pl/Zxw8B1RMQk9BJuiyzl5EMoL9mel3GnD3h02K
LBmsG3q8N9D9K1dlRflRxsNfhRc+QmSHF/4ULA0EH5m5OvxovUmO0vv40Zt67rk1
A9YPfCtejbDxU7AvCsg6EhUBhE57kuUZ39L/C8eyXMhZVKLHU4o67qCEH+nHDOUz
px9CkusWxchtJTMGG+pekK5ZZpgNjzHT9d4fmOHnGFN1GFvdOdqk3MOkjE2ozLvZ
u7neWvxOhf+8bH6+poDZmF7qU4FLm9puICaPTd62DO2gi/s6xcSQiy2qx2Om4VtV
wbRrZ4RqJIjGgPyzqx7kaH5YZAHQezZTCABdqcdzhr2O8tEPKg+P7HCMAa1hD3lL
+yCGStXP0AjC0YZ1YbWWpVrOm6P9gsBtDfuLtcG1XnALpkSpAu3ZuTZJsZbWZfmh
HONg7SSdwES7az2MV9XIaSzj1LlxbNc7LmMqt3XJgsHLxPuwti4VdlaHr1cbCTnk
LpFKka7kXUlz27e9l5coCn4mp7jni9bu6bJq2KrNH3UV7F8pQ0iKYq7z1aAP5lnc
3NQ/YKbIoNeqkw44sypcaQ==
`protect END_PROTECTED
