`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AQY6FVhO6Nk7cmTTCatsQA2Qo3DMZl3c5ojkssLDUvXat4Z5Kt9g1RKRuebznXQE
6PAkFrldkxUwEQKI33wDOeKnCoZ5w+mXCUqTx0UpmtHAAsI9Jn5duFsgC8yU+ZRy
UOmCObTZZe1405rJ3PvowgcwZ8QCrbl3fr+cYS46iLl17UC7zO54JALbeLzUs9KA
qiX4cJFn/8giIbRMvlwDRzQf3QG/fe2JqTzTY7ckjwgLYCIpu1slUP1MhPmCLhfR
WSC1Py179mCVjJzQyyQ+yrbVqpiYkQoK23bg7MvqJr+hvX+U+m9qUI2HkzS2ljxt
BGb5ZShKimJ4CyHnQNRy3c8jj9cnHccazXBwsUffb2Bc/pPyb+UbZiml3673SozW
95OM+AtGLhpTdCTzUL7cD7TDIBcEidpBen+4DfVqGvu6oY6cmxYRn4CVYVg/Bdqg
FCBIkhOjGu8Ds6cj5za2psZaYPtpCm9lrQRy1++aCpoRETgL6rSxuWi2XvD6qehL
1kX2LxoaCAJLdMUCkJ+FboXJV3hBfTaQFR0ia3vCB+6XqQsoY5495rOhCj+Ko67M
iCX7bJMIHDlCzNLzw8HT6wsM8+fdUuYUkYclwgjwKO3hLHJJJTf7n96xYJO/3X4f
SG/gdE3Kkl569OnZ+klp6dqZEDPI6rF8U6lt/288kOSz7Ga2o94MLW1c+N22I1vR
dWYr6GWfbxUtuhvhv9DLwDIypjdZqCG08dM2wU00FAYAzntdyoU5fGxCWPwuzB63
wFwTLlqYVcxMbWO+pYQmtpMugQ9dJ+5K3Ah31WdD62B5F2AtPm1BkRXMDq7x5dbN
1YGWYsi+QaEBD7Rrr1HEvHCr3uqNOEf7EeitsqnAY+xALvNPdyr/3mzHOgRrlVAN
bbw/CE36L4JptAVeYMZed9SysdCNGbhVOl9gxhSdoLj1ML43etVFpXAqu4EywCBb
M184NpiuP8OmlJKJrHPuMp8TwqlV+cEIQb6k+foeENSd5DmcojgfLGDIwkSj0WGa
ybhjKeZZKnxNo2vOv3aeGNL8VzRKYHYoPjxg8huqUbnLS+DxB94fg9xSfB8djp3x
FhpjrF5JvPolFzVKfasJvYaKIqCNK5EMNzV5sgow3SCbhHfxobXnWrvy4iLmvYSJ
6y9UKhfsDiimMo1aDq6VJbzI6ruZBMQdgoRAteszYtSajJ38PNNt66FWbJZXejec
g3gXCFo4IP9TdsdQDB4UW4Yo4KRt1P2hCn4d1xPPZUEm2J0aAQ/XUFQo2Fj0dcuz
Impiuuo/E9k2t8ahkxsBK6xrIlBv2v70RT80cvK9BWkoH7cLKj0anDVCXhwCbd0o
0peorsK94hOeQAsm3NpOI6jVVN6jIVRDTAvzeALcL1bOLWgiir/101RuedhJsfgD
ZhY2MGdLp9Exrr04I0dkZc1X56QS4PsvzjxaROoRlxwbaRIX4AfEiWx2Ly9N9JrJ
YgLyLiG18alZjxH54hm11acI4UJfdxN9nTYa39uu1lyMmfiFf4mamu9+vdBXfPMQ
N4vLzUoBQGIJnzyb2H1bSMOD04+D4npmKBDoJkxBmZyad5OWsBFGlqc0NoyQ95Zw
mhlPmrWcaJ+wFxtI3Pb0j1jgXgeC/epso1oA6XuqGnJME+bssZ1z94rUCmFDgh0P
9gQimz/AFKVGRDmFPnjPNPUp/mmNmynup5dl30t0BRA98YWPW8ack90OxfTdDfyz
8aff3wT71s2X5WTIIioyNsnsXC/UryG8G+28SgIya8cHKQIpxPHcrZbi2kSqAe/U
q2oVqYHCPxX650dkyPAAfeqCE63ZEAarsBlzcMxu0K+DqoGqdoBMPkPtEbPRRB6F
ZnQtgI5Nc0pLn4vBvcC8NgO7Zk47yOR3+bQcuDdvEM+k/Xx2rcaE1LCokgduWRFo
0rKyS48oM+26/sCUhQIwHvQNexT99oOUVrR86wYfmtD1CrSxTVn5Wr5SXC+xKHih
zJTPbb7PQUVoh/QRwW/eS0ytfkgHxpQrstpoIRrBb8uOf4I6iHTlaLD0q6/v5fiF
k+9o5Eyn8knP03i6sIii4tpxbrQ7j3waeYMdNviRa7AXcxKJpxH3ck4zUefMbnf7
TSZ+td7W1OzpB3l2X4p0iIhEfwzbg8fGUq131SG9k+dHU/TUzVqE+ZiEIFLG33qo
Dl/V+0Z9rt1amFfdK8bj7aGZhvPnABh++72bQgUEX4HXw4N1w59UFXXJJxyUw9ey
Bqa+AZxk2eLnLUebCJv+iDX9aJt5wZ8G0H7nHSbutsFtVyo8FWy/tqQ56fNA/58M
ZRYYrF3ANYXtVTpC6GUWrSeWHD+De1R53uLSJl43i2buvhGv5JIq+7Z+exMCyTeo
K4c9x3stu98qlwz5CaEaTc/qv2SZnzInHpFhZ2Vap+lz1gGbG7JoTNhJ7n57/1Ks
vl/HZoaYF9Kfla0U2bTcjsrGxD9GZ8EzS2bmOylbwLs4LaBrzX1G2uavDi74QDpC
/H72G83OGXhVrZmLofXhZpYjLLyPx5bdapuEThxALOFf2r5E4uZQYSjo/2rQZ74w
BSZUSq8jP9RkxQ2O0hkD2qJheA1ktp5R2O6tZFcJF2DPMSIhzEDZ0pNEGv4/7cTh
IKj5h3hsx7p3u3g3B5e8gKs7YDgvJ12LWz+siwkn1TDOOPjqrW+r1rfvB5b5prJ9
Y2/ZuEDOE/83zAEZXfWATsy4kUd10Nnrn+U9+pxaeD2r9NaloRGFticpcv/AEAOr
a+cZCU8+9L+qilD/YGyref7kWge8sfRqJKZ/hf/gIH/nTyu3ofOgCLR6R6N36BBz
Y2oVUZ6JgV2S4cck7zPm+RuWUXXa66/xSzN6SdK944WNK3zNb/6FeMZEbYC8w/qZ
wvrl2NEhCAoJ8SYQxoN67Q0EGoi6GwYurT8P/ivPHO0/zVtTBCEB7NAf3HfKEGcR
OP7Yi9SPCT6J+YIyS/N4gX5o01c/uUHqL3WwWLLPQKL2XusHeWeGZogvvOKjQGV8
36bk/GbHNqSEr8k2KdBT3wHRiuaMZ8u0HhiO6wmyQrZ6pZkvj8ZpR8mJsblAn4Kf
KnGLviJyltwQMwrJloS/rMqR0puQ8TVH+rftQf5YG6T8HqHvbRitFOEfCpIAOY3V
yTqw9NpqG8Evtfes8GP6wCLOgiGqP8TGLuWULswPx4aOh5X/Hc1xlm92+J9vbqv9
IICSmRaosbmRbWMCK0uNLOVOp6NxL0xA7WtjU+P8IUF6+O6/iwu/m8Hfi4XrKzOH
VWSX9keDdI40iSfbwR86QxGz52qYbDGQjGckop1nJK66SXoTGNZxvYKkFve7lqkL
Eoih0zgsI/Vatc+XTat9Kic74FM8LQKOrP5cCrAdqzuRZtkyhif/wtT2Ia6043Af
LOVr/zvCKbD97YVU/wIsdT0hJRLjG3pr5C+fKhec9WHMu74QJxDPH5iAv1ISZ+vC
chKs0sEwS/PqTysUyEd8d48mCAG2z70F/Yh+1dYOuidbhygB0TFtCY35ZD95Jdvh
b5XpgSVovl9WvFV+v1BBiMmZ5LQx+kTOrT39z586PUtv31XdrX7i9PYHLnhjqsFH
/np9ZtAhLJpG8mMj7NLLfVTmGnvFXl/R79hasfjcVukciNB65+3Hr2i9I5dlRdRz
jTOj74L6wtWR31IqTqop7tjo223Xq2e381e0xGA40zdW0+mfvz2tJb2uCnmf3oF1
gXbJVQ5A66YpDp1/Dqv8+kkcF6gktKOXmz5/3AGJxMaKO93JdIKm30b6SO+hOQ1r
KdyQvxZ10Uz1mH3Zq1d3lE1eKfEFmqGSpE+jeoLL0+k+u8K6aIkTcbTFfb9avfZ8
D3skAwsZeoiHRtohdutqdH1Pt48Nmri4mSGcV7AlJ+PrM+5hKiNTpKVVBd1KFmBQ
GmYhEBUoWJgqTRU+7Wy8V/WKtt0+95xPH7ln4EJJ469XRbnEk/lDOWmjeADeCLHu
KXsCmw4lo5nK74Pf0cUJAIPghZrXeLzsO0KFena1//2WzPWHYFPH7ALB+spVXs1S
LUubiBxHvGWk3BS+oBtI1dxA17Beyy+aQmQUX8VM3eHyln4pvP6j4x82+y7d1+Za
fSgNiGWNTOs5xsfvk3Owx0RptHP01nQLS+XTOZc/t2cvA+ydZy36mgfULLRpkbLb
cE06D9SFvLZY8F3c4LafJ3DIcDS5MsNjmmMQAsha55zSo0kFcXBgkj4GYYjrkQay
oJG0Zlh+jkXXz5EuqaK62EdeQDMbFovNuhDUUmT8LHe8cWbuHuOjzSMPN/S/DDh7
hi/KeVFloxdY2Ft7Veq7msD+SRVbw3lPfeWy3OVXrqHS3vaxeamQbXalWvifQDXT
MP4npxusQddtR62p048tIERgGChbBNBcJTSAoKzwRTnEPXPaU5b/RTYQ7P5y6hnI
8p0wBsV1ql9gwr2hbA2sj2Bpetn4hkUHKUzrXH0teVLuXTMdVdhVroJ0rlUw0mFZ
Zdc7gnpQRAz/wLtdrtea1yfQOkP+M4fqDIYO5ok/A2NbqBZOqSxmc6Sto3PT7vA4
iFrZt4/EmSSA4RetzJETWplzIPnJNRWN2wKYKbllno8yaR1Id6T9F49QhJxYGy70
/QEh6HpGyS5P54OMipSuiYIQN91rZN7Np20ovNqLOTN0c7BL0SUYkG69LhHRs3oR
qCZBM6Qybtq7/zxN0S/dYxr1XkgULIjHgmJynvPEJQpMS43dVoKrm4JoO3wP2tKV
9LdP61T4MA/wBO9qUvhG/dMNBNvqqn1bVQHo8SHfmR78EUOXHZlo4XuaY9SruFQi
382mx2LN8ciC4eRTzxDy2nCte6fvBYzYq/E0tZPB5eDtMakMVE0aFiOLnHegewSL
ZaGvc7Xu3ael0arPDWJrZ0WkSGSbqlBk6W4eu3TR5FhSmjZuZBSr0ZJ+nG4GSaTj
q0wdski+bbmWMPMTVi72cS/wl0NarBjbJ/d/cakSZLbpgg57zBnnrXdcOApx770i
Fqhtn8uSjlnHzTOfTZrOtzfa7EZeKTcMqG2/DGTGWnPEwrhPuKsKmCrrqMOGU92f
ojin8APeFh4JsDL6/kUIhlUuVJovwUJZ8ual1blCkJq2JnC48rl+8B+EnTE9LDon
+gq4xr8GVEIijXfGpWYFFoz1Gjcluj/8aAQs08exsQy0I8IuhDOoijDaun3ft7yz
1mYfhlGlAm5SHPZXfVF2DMfqyhG0aVt54e4yJy2ne1eha4eCukURQ3acNlIrHo4O
SoAUdKPdazsWAKMd8wCBXU+HggWfWFyusQdgdK66aal0qinqViaXnSaeXcOap7YJ
qDw/23Fuwohkfg8qtGAfM/U1Py9a6P2VqEkGci00D3IfAvZodHHRO6ph68qDA2jT
ui4zPj5if5cEDfwuBKzM9nK75C37ALAgDEpxBxGLGyaJTuqCU+HGvZFUOwzcgkNi
6aoj/yH/NnYEVV3K44V3r4ntoMg+ar9IfEq+UffkmD0NhxerscPXJzqdebw+u/Aq
gFwWYAemHPxwy3NRqxrsyaEmILo8KPBHYrc4mZnFBKOm4wnmpnzdrNvwo5L3/R65
8jc0x1T4BlyNjEO6Xy41pAf7NIz9Pi8ae2wlVhuJIcrFRS3/+lYQwp2VnpI4fyj/
kVUIdVqs5xjSWn+XtTTSiHRRuwLyNOV7W7yWDOUlydPM9OdPMSqVUNDAkEjgsbr9
6puZr5QLATThA++1sOO1Z7BLJWQJ3T5WYP66Wp0PmP/RU4TIcWxe/gTNbMXDysWE
qmhsA1LS4MKFUTO/REKnZmLAe8pOufV3TXHcaOG2Q0G3Ku0ReKvtfujwTueDcwEx
tg0BNkRpxgdcY0yl+hxW3tC0VX9Mx+bNbX/NVaTU9uKLD28pP27Apq3+pGhkg3tC
GcyhnfS+QGA6TfQ4iUPKOUsC6/yFamGkjmTWR+PZ6iJU24xUgrgUZf28A7eCaGoe
R2vfMJ8IRcTAxp0/dRvyKgoTyEcQWYAsTrp3ndCBHVqaM9MbTx5OVn1Eb0tploeN
HDoj/KgjTexg1DX31g7hnGkjewZqjzNWxVWhgEqRS0ZrREZKlDdhLN+QEtNq70Zx
JrL1Feokjpfs/jenMDJV5e6qRE11tfMS0P7kujh/sR6NStR9sLdr9xihZERsew4w
7nKvpadQtgpBu3Ww0APz3VMrF9igZ9WZmtKFuyKS/YSkePokn4p+DIhr1pDooW44
DZye1o+McnfvCZmCKKBQbD+8qLQ/vzQm1m2pPm502NPIXUC9hw+Qa4WTtp2x4Hl7
Ru9GjDAHAsX2NwDuTP/Yyt+shVsp2WUaPTT2vuTdtyE+0dxNLVhH5kza5PdvxWo/
+0sVLO5fWrXv62Ekh2puj+K0MpXDNDQ/gQv3+Eohfy4Vv77C9eSR53R2nx4jaK2A
sVfyHfHmjSHIzOSYuj2Hvh4oQvVn8v3M3IgG1rKHIBWSFqyk4VwexxU/NlxyQMbk
5h98/ULzPr8HJZCUMM/ragMqL+OzUnNgbnkfdDc4eMvrpVjHg9SWADk7uogJHNAx
kkNJfOUFQ6DZiv9xf73MeaNp0eX5YzDv15dSsTUM8/O+naXi1lKog11+tXmffIur
YD31jrwREoLeZjUFgKHY2vLjfxOyjDCK504bs4aZiJgRUD2Lrj9xJ3CRC8ZW0vtO
NVd6Jzo7gmTXIhB5MchahhcZPOpPQq6Ilu9be4FpWBlIOQceOwhCbR3fHqjDDKp7
4YqZFeA0OecItUvWIvv2kJxSwWdN1CY6IA1X83mFcysq46Ha/jlHaObaopFXXqoY
04X2G6mfj5a+E+21/8kZyJp0RVZFPIv4TTaAaPKIQsGdAxBhDuQaw5WQTbn5gDJV
yT/EdZW/8r4S0+3A0Q68/PeQtDJnZXD1rDdwyVbGRz0Wdd+8yjKfKkDq5IFmaOfE
ViQXhtDacA+JPH5R4o1j9dyp1IOfZgiub519UIdj0nIZ1HIO3JHzxN3RMe3Lk6uc
vZDKqta6mBDxdlE9vQS2HBiAOtOyBeh7GYh+V9wBDmtATexEr/ZAvex5MmbPkWfN
VnK+FTMRrmYbQQd+bn6RucqgdasFWqvpUwE+1pVddK74lfKzoGdu7b6fzPRt3Opz
015trCu75yotuKGbKAtBlb0TdUHohnho/pztNiI2eCKr5c6DQSUuSUbPX3upxToC
EnUIJIOrHKlL5BAvEVhDIR13JWugoqjbU09rtJfqzeWqzbn9wM0PwZJFzokV86p2
cqA9N944uJaycDh/oWQKQKpZJNDJJKKmX0NYD+GGzxyxmrZR6xSeY3iDMAe/8Qbm
k07q024Rlm6kB5kSI83iuSP+pBcFnCrqhYwD4zhRWccIbUt8jo4p8V//QPfy2g/x
3jPQwChsFGjFEqbi/epVxbd9072G/hFKDLYBv7QHnrSi1u9qWlHpze+SUrOQ56Id
lr29pUv4qQ0uzdlehWunPD2P/hLWoX8PntsMCmaKYmginsp3VTkjkEjkkBTtdQAl
cr5c1Z1qtvv24Zp7IWklcl7l0bQ8N1wzeOyQIZeZjSEl2NtLjR47W5iXnnwMzX/B
3jcPNep2e/8IGC8VyUXTGLvviiOIBQY6awd0yT5u3q0/kgIwEtgKgVDGjGzqoP5x
VqcYTqos5jcs/ZNtKjgT2I75jU7ynh4gfLdP/JVDiD7STG4b0vCfkvvgWh/TA+E2
QdK08wHY/aJncCpWyTX2zmOqdWV0WzhY5asfimt4GgufFPz2VXfmUPoin1rc39QE
jAxf7vC19CxREd/xnAnei/T6nwL4f56GXTKq1Pfc/8WbKmTRYu80hNzngBjI6qu0
mj4u5UkrKLUbvZ+3qtLsECjkThLVGwGHzqThq5VBuc67zfg7ALCOnY7os8YlIr5/
CASAPU7ei7zRiD4FlEaPj8yK+BGC6XX/N3zSKmQZceZpycdmkb57ca+aupiEypIt
QBgG9ZxqJdXmmGo4dUMMGmO53aDllEcnG3PwtEH0AKmCNtpJj16m2J3XRo4zVoCy
nglRruwcUH5QOw4EA0yHPF6OWaUnIPZ2z9WyYEGLlxoWDT8qjmBrqau/RY6RVWRB
UhRLRDE4vqeeISK2HDyeGfrIj4PgrvfaVdBRH8OrLHw/Ml3b0MIuHQgnS1A0vUok
jDswCpsJosb17sOrw/62VgjLnomHV0vdnl1+Yw9NdzkRoEWYQ5ps2tNGlShKYZlH
NfUPCUDsMDNpb1X0OFBEyatsLSyYDaVo9pE5To8uAoeBnsc/C5dncC/KJ1qzRvOA
ocbZW4gxGfKJqVQbW4/MmyIRK0XK89aiRHZ68/oPsEOwUfOpNdwj7I7G5zleIZkB
0eMjKXT0nwyyfcyDLGsrRUA6l9plmbx94xsDB1xrrpXFKoL/BmfyNBhwQrPOP1TH
KHsUdhaiq/8v3GWdHZIXZ1EvrteHJMN6qXiXKqfeA/iMMipC2ti9eDiiEZ1XrW2L
jA8WlUE4qNhgBbQ2hNpqu2WmL5vfUloaV+QPKW+b17lFIQ9A/IeOr3FHOJvcVlZu
BV/K9b66H92GHTbtG1vVAK1J9Iz8ASY+4ZT72N/hRE7uKgd7FydcMjBgwRx8Dbaj
wiNIbELvqzfO4VgdyS17/BqdwVwn2iMiJ/LbqgzxAT16m4kBJHR24dH5TAFP/gj3
jea/n2KhlQ+fVGOH8Huk/G/X46JQ/F2Av7D6fyjwKCf16pvqHFemFHMVPPq3FZJT
EeDTSlaJgauHqyUqNCXDE47NSYoJONpwrYXM8NzPSmD+k3KrBa+99M8UNC+dRjhc
zB1fCja0yQgpSvRUihN8HxzvSxen+sGbnemd2Ed4MJfyc8jwrgZfaHiWm15+aOXR
wMscvbS9f/O4t0gU/ouhqwOVzvUmY/BpNFZFYc58OjzBBQd/v5hMVbEq/f0w8rOy
MRudOKKq6srsZ2tQeojPIZHv9DOX9T13Phlk1gpIrwOVX/v+eVZXBn4iS0BnwA+I
n8khAxOAvjEX5IMN6cf9ez6voW6wWYNWftRKXVMZWCHNj70DatxfmvaFSC2EW7ly
JjqKsIy51twiFgecVuvwh2sH/gmFFTbSsqhZqXFYpoyOarZJTHKOZIeuB1gIDhrz
xilS2XZSeJNHACVjZsAqrFdjKZF3ROVAiD1hiO9CSmxop9WjQ0PT2tt0Pt3bwOfi
2H0vb5AHHh8RmfttdZWWtjK08ymulDNgFKBzXvcrIlNHKzwnJ1yKbulSLd3R4g40
Pn3sV4Re/RwqnqlCGipYK3Jx5U/bZnHMzdShrs5r+774OOvJDkaKzG2EEG4t4gSE
QRhBO6ab1mB8Fi4b4zE976ax3AUKZfO/yT2k+2XtRAOc3ps6l+eylxr4TT4A22S+
Uaa/q2Y2OGrg9EFwghfV4Epb6sNgOAZQX+Fkttw4EUYw2LltIw28xsqt7MGv0vbj
IDZGPv8U0LL7CcU/RBjb7gJm19ieAMCOJ56sikflicF3vGRlsqpDi9oMXebXvF1W
eyvcMAYDuUdlA682QsDN+gCAf/3UsGLacFO6syNVC4KyoQDux3W9X3oJHvfYg23I
Y13dxyvDPDHf0bA47qJ3eazZdefd16GwhmG3r3fFdoED6Uz2gNLZytENREV3b2XF
pWENTN8XNwO+l7I2U4ig4nkj+c2NqnmWmMO3dh7zN5FdB7sRni1qWXl00VQdPTbL
qaBisQ2OUt2+EVNy70tqDzc5s31/f3bvqrgnib6Z96QWTK7xQd5Ixu7lQmkx1Qo5
Jv8y+hL0sWNIm+Sh2rHRuQMoa9+02FyElbtcqS4ZMorm/UpToTSdN86e8QUSJNU/
P0q0Wm9W9d0Li53b0rvQiBctmodJcl2Dx9MtK3paOW1dpvXsKEqG17uT7+wFx605
+ZCQbAHz8klbv3kadk4dlrYx+zhJoLACJLKcz5lHgbsDuGWZqp09Ll1DpWEBsSyv
EZBmt2vvrTbAbSOmbKhpHMZfn5nBgrZmQyZ1kzU8m5sBFmVjSXIMqa+JS18CuT1k
X89WKQlqeGwHD35ulVpQvrAFc1v2aWbbvL8CTavL4/7nmf1UYdN6aZSzMaWSnWlR
1vCDz7U5egKrYjrdXCE40N6iSxn/B8qUNFPqXlEy3TgGq0vjFuubAalVr7puHdJY
uh+Ymt6Vv4q88R2DjzDBJ2Q2VGw8UEtrPLzTlGlBU5jpEMS889F2e3c+oOqU3TbG
KmJBQp8ucuH+kqeQRE0Il26ehK5J6jLG2aZFm/GOufd+AcXGI3GrLG/8G4phwtai
BRgH1N9YDTy8nvniqj7z20EFL2OvnKTYGoEtYfDYfYIwzlmXZ2VhBL9mnyU/Ok4D
NuNPlmChu34QJrxH2EZF0Gw2+VvjISkhfsL+brtn1kQrGymYAsWH+yHKz9Z2Sc5l
Te8lHJaUyIOVo357q1F+Lh4iNW5A4g+JU95VKnAlc88PYzAdrU3rD528zVBEpmXl
G5xPd4pDZlbtNM/H/j8YaYpmjKSw2AOPy3s686h+ijRBT1Cly/u3P++UaT94n282
UU0A1xcyJozHvldXOBy6B+cPODKJ8ZyJFzigL6+fL+8QMt42kAX6n0qKrtZXibjU
4SOJAUG5YMSuo60j6VBFe9yz0cavoybmqd9VLQB2ANCcQOE1fNszWGscBsHymTxV
5S7666t/VCmD3sCsOup7ggSe2zFF1Y5g1ulLgEQMwyeV0lWDHhtBboNeKzo1tCbA
K9qhYcsjuqqiks4OA5gVoEh0XNl9iquoE4udx0S6k2xx609dLqJrRUb6FJIvUWKG
pNh76okNKDfQPKaA04SbZc3NjyUm6oatPACvD+vc5lf5OLdq1qhXNxFEHT7saPel
jdjLX23ySStRfFbQYix4gPUQJua07F1oP72RRsSu3DL+V30xuy8EwOzSq25KSfXM
MdpXrwSP8gLkeg1F+TTeXRWenqigzOI+FCWDm+f6pN8I0bGMwI2zUQdwYd/Ww6bj
Wy4cr/Fo0/TjFD8XeKRQF6KYpcPUqjkMfEqHaTRmZ7hiZOCq6DdRCZd+9VHciTXt
I1/JlxDBj/NxzP+z2pVS2+u4zFGc8Axco0uWoPntHYmdY38UWhY6o3qwW5OlbbyL
cXmNB2/Qa09tuFAGR6TYaZe5ZlvSNdpEkfsy7CrP+mUzF8EA90fDOWWfzt0j7bF6
OGQfGBZ9n82vYkWx1MwyL0PEfR2miDTp/WneIGo0s+8foWdybcVF4HUKrAFpUT8B
acJQnkdJBO8HrgPXdwTYoE6NzaohlVnx29w2ZFjlv7HktaF2dotOk6kQ4SF4XtDv
MzX/1Sp1jBt5K/dlRkeEff7fWvj1ImMeEhMscidMTFLrUkibbITc+qlgcojEO8PB
JlO/V0+cYlYq890q/UjCVQG1bMNDNMqf0kS4OOLjUpO7u45Q+IfnLiNoGUPpqAcm
mYvYtMHh2FAMUIMJyoRI0dU2Mb9stwAs4qXveAhq35i/QgOVrAMCnfk+DZomVwg2
5KuN9+ZmQmXStmIu8BOeqpoDp/bI+l62cbe0eSxXyKrgzXYmC1DHGID/Me7tOUJh
4Y4Z3ZQKqxyQoVsFgZLcNxw6iIrJNbIkdxqPLx+nt/Do5/9acniA+X6uN3eeCx/e
oUEFtOIpZeO4kDmeDKrGRyg+S8sKkcteF6i7DQe8pC1gz36vnsJz/1oxi8Fx8rsa
YMGhdkx3T3q41A6AlAroRjUizRtf/07gdZJUeecYBQRMDGg6rcn80+hFp99YG996
8kynNfGrN6CId1C+a6hZY5uqkpcHQZdIiChayl1++Qdbr2aFaJ+OBcP6Bb9og1Gk
baI3vTtre5KNPWE5v86yf1EN/k7zyR5G2Ebmb2DQE86Gu+mFXt6QtePfrV25oVUi
/FGFb+5VRxY1IrvaeLK1SgJFtHjrARu1PtwFShCp2F4I3SNzgk5xwjNOtzQqpRXT
oxUZFLAtSIj6fqEudX87nG4LqEdIaqnhqQVwkmoNNkavNhGR2gGBbL1pv4UHp845
y9dPJDS2H9GxDIoEq4h2SLxW2n2jzpv/TCUxv4l5IhqZatRC0AnjgfBcO1ouw0Ol
SGptnddJOsGDF2rsQM5XTQLgRx5kHNF5Jlnt3kgbPhIweH90XaNpab17ktO82Y0T
8QovkDDXfIrLaTbZzqxkBSwitKdePkjafvgAkNw36pUdlrNYZE0ppb4Ao92NocKQ
T2vAjBv/+fe/cnLqSuWXokQ7ckoDa0R5FbaGg9gqQ8tRLfFTtlNBGeoFjYfYqBJR
qMG0mW1Ek0Hj8Bgk0eYAE+5YpUoWzELSi0k3NoHORQqlC2IalQKMq4utvND/QKiX
4VsJiIrUmb8gsz0YuBA8c85sp5TYN05PKL5eH6J/RyzuEBYSbXftwo5zwIb69tfe
Pe6ax+0k5t+bH9u3xjNumP2aKtXrQBPklEbhUthNw71qUT/bg/+U2kJg0zqzkBWT
qPeYm9H1oTJK53je+dDSskm3RyKYtzelwp6Rxc59/iN0RxErNqO3U+TJeHgC+N6O
rYFzlRiPN7ghpBwcvjv9C0GD39IxTTbORhR5w5IcfM9sWNbrfvm/riaVN7AsIgvV
y9uZxZ8SHyO811b8Mj3WrLXPQIJDMi6N3uGB2TsX4LzXvOXvBbypiGXFfNrReZox
XU5NhO90RHxJhyiVRxTbHAmfWIiHZgKWvMp9Wbw7UOdRRQurIv4HPK6YbRlTEZfH
qrHfhTZyWJrS6mWfzev6ZFV07uykIyu7Q6t2TVaOjif4pPK473L4oOJx4xtlJnhu
GSnhXuPAMvN4xtj7/Mn55ySvZkz53BazuN7v7KaO/SZ5BiQs/H5PAsSIfr2TlR2e
v1SFK1N4pJ40kVVrlUgWYXeFXvn0071yr4dxIhRyxl6e87qmidiDJYjjPo6PNPL/
5kAwgIfSYSUrV/V0AL4XIiNHCp01kXzmphTwnTyFXhgr3d0qXdoMr9PPQmFMtGBx
+Xm/gEUKaDxcesP+Kg1X8ruVzPQXPUIrwfaLX3Waq9RlA4mvRRovtpYYeFkHPE9N
jXXNxynbqNQg9GgtYzEb/wNa6OlQNJKS0nW2uGYndfssn0i0FVM3j2yQS7ma9q7J
LtOTaj+WVUS7hHdDBqpHOJ6lcIkyE+T/tynAVfN1yGfdm34gmuTbTn0Bp6HMVO5b
zClUHnOFmO4gNxF1is4kcp65UTulGKUCwrBNLIlfdMDm0RdvexsV429ASzxH7llO
/NFRWo43LYcKT/Y7WMG7KL1QiqdNHbPqOE5ej0c+FkvLCK06DDSBE3KSTGuvOjfV
L6O3PI5Wu0Hau5sm6Piu/PUcaPjm8j35iaHwKHqC8vzaA6oYbIcLO4VYSHVSi+zU
SQpDGgfayoLtNgF4PKCE8R0LSok3GMoawcaIPXo0tOakR5BGmhnbl9/ldD/lVaJy
unh316nVwZtf5Ddy9vd520gecrkv3648oMllfIzQGFi0oAxF2X04FFv9ylQ5f9dl
yZa5H3DhKdJJVN/EeeIfnqj8I6nHHYmFtRskaQXbZh3b/GER0Qr1QU6hExgbGHiQ
LISbFXi6TpF0pndCXFRIjqp/xeQbPZjYx77d/zmzo4QzdxaDCOUdKGz5lwRFx4lw
C9TzJiHRB/sV9kK0n5vxxZaXhxB4dG0PJfbq0qCX4VQIgHOyA/ibk/h7wAEFfc3V
kplCkyO18oXLl5WFbLeGnA==
`protect END_PROTECTED
