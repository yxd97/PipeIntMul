`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4w49AhvKoZs68t531CYDXdcPURYKOeNt+5bbZgEwpY5wE3M3BGTbgMVvstWHgcxx
9uGSej7hQfobB70czg+gU21ywVN05GraxQ0hwnfepB8boZrEdc7/HDBFlZH16Idr
sa1gsogasTPFAq+DACRpmfK2i567mAIJp2kFa1fKmtAVt5VCsmVQHMh+iM8efiZ2
bjfiB9MM9e0IFNw7k1pgGHPmi1G8ipfp0D7YhjMeBPoz8i0xSR8bbVm2yGwfqENe
rVQxuMXeNav0qvNKWgV21NfZfeghVzKdXIiRf/OmQ+Tgfm0ZQGcvGeavVEQ7kc1P
2BCrTGbxZLqHh5dPALE3R1nQIoOpkbZ2f5j53ZZWEnIHGAYcAF/v1ttvQoEU0nBV
bu46Xi3+rzjDkE9QZdbl+SRlI+mlZteJ2N+5JeBhoVSnnBoti8gnK8liRbH5Oqs0
IYythDGjmK1xjAwOtxr1IJbPgeEQ0AE//IB7PLSdvZKGqpM12CJk0vmgJM4eGoUA
T48tieb9aCZy2Z8CnxdA6kM70uScIQE/cFYeR7ZoItm/w9XUi9KuqQ/RGkFetEK8
AJgqcWYrwx/AYdjpBpQrzZHJ6xeg/Mw1+Xy7dTK3vgse0R4pEdqQbzYLMxSXlIES
sl2bNukYYeWhNvYLKGUssHfBI2+8ytFOzsZzY11isPYovt1pOeowiBvJZ0kVBVjW
/b+Io5rkEWvgnPktJyPShQG14zqFJ/rZH787DMoVkLGut9uuL0IaWJVp93+fB6DP
ZP4kUFcYsYU7TS4JPelpk0CZ8OeY3+A29C8svbi+kFbbLjQKAxOdeRxfkTqImfSU
tXHVNi1/+0O6ulJd1/mlKEQ/xkKMyUaD2AIix2UlLJ8D4PMEhytJTvjOaj5dnUG9
LMbCu4My2Cf1xxcYtmtwLVk3k+RPK1Vx+JwuCNJI0sHpldqucdCk60QQZ7vAOZc8
+B/lrAzBS9sTBQB1MC9b1AsmiqyWoUHtwD6ks8Yl9yc6fiiuZZzvZbjgE/32I8ri
8WAL74XrckFgfA9sE0VAleqtQU+vURPrTDlYit+xF7ZGsRmOgwSqBbhqMsAPUkWs
0/OYgjyBVVp1AI4FlSfNYm0vFnHnwz7zGAq6pbP2JhqxzQuTSkW+XG2osYZANuLC
cIYJNBOnXev97A6TNLh/GSocIZOWa00UltGsi2ZuYh1LyHkxqcOROgc6/5Nf1SUQ
K/KON0VYiBFAR8bC15fBL3Z5OYUJAdmE0g4Q9+Iy5oP3Zppv+GIuDAuafHpG8pjg
n5mDs8tDGph3ItHVEbJKuR2B0xM2sjrNkIgjeKNNz8oH3b3pMqTIYsGr8LWp7/nO
AHm/UndkjjgHEuNJfo5Q2ft8RHuLEgOF9K1QTfp4oyzKOjyILFBzQOnsIQ7f1FB4
JIoSDLbNFUyuqn4LKKgbbLq9QKqWMZAVOPyW1hMGtJS7iO2sgvqjCUh2huqB9/ed
qFpV4rrrvH5QW6zLRnnCgP4NKZEeQGpBaKjby7M3amOmRrloOean26DFjCo72RAR
juFeri1WFmfXgJ8FcsI6VjbyH2SPm6NjPjqPtkXxmg3nUoxpMWaqhW1v1ue8L2+J
Gqf3uWvvenQb7yKEjeLqVZkzjwXBE1kl7wQpw5U4NWBY64Pscd+puEGIJn4sMtBZ
ctMNfDwblJhPDApfCdDJ/bvMEFJorbbLWku7k7tPCY1A19okJ4gt7mfZnbXaOOUo
RrZyGrpK3FNa8wBcUUpwtWYsnDzVvB+9MFGpHFeCux++hZ5h8OycG5Dm7kVy/7LO
uchP7i6XyYH1WorASAjMqsNGnFUyl6HDQ2FqW4M13SsAELSf5h0e1SZz4ZrsO4nD
muCBWPyzUYTBTUUqFfAHdQ==
`protect END_PROTECTED
