`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kp3A5I+aQe/b+PKV8FUMJ6riIZXHLgC45/cY/KmIX5osdFlZMQ5JuRhvnf0ILCSH
gSozsrH797CrJP0quF/l4n1vipTAUyv5Ljo6JiP2YNjYLXH/C4JB3RUMpmRLDsgQ
kxr7s7jbh6WKLs1yWM2MRjQn9YRyYaj+j8ZIgbLEptNOa4PjrlqyjNnKKKknDyW6
mpRXXojeO1ymDdRqCX0n4K9nkSNUx5DdXDMOcR2b1Cf5WNkGz9Po7kGKiu7FLbrD
`protect END_PROTECTED
