`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cDsWa5Gu5BZSHgvcJqyz0VyTRbqXU6agTSZIAFHHq54dOacto4piljXFRzxJtFqg
vbt/5ptBbZWU4Str7qU07hvywPFl3YZHBFou1r/ChPacmnxpR/kijxQqEcdzCvVu
c2lJ1yLYzGqv1kBrxEUA+d0fgqDrUbhga/B+8+p1NBvB8hAl7MRdyVibtG8X9rua
pczCjeT1Uo8O5Ito65E6jjMBniXH0tQGFRwtiAhaWru8zFwjxrikQayaYAjJ5uxU
`protect END_PROTECTED
