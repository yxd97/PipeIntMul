`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fB1pzD5yYmCQ/CYsky8GMCN7gY+gUFAy83byBzp77885CgRuXeaoef7Ikisx3zU+
gxlrKRYAHJmdEWay/mdBMvzK8Y02VZRScFuv6Ax9++0/qQtstOG+DjCdjDNuvR6c
lCpHZeuVZHWZ+gWVQD1MrbzebZuPV7C581TAbH8TiGGfsvebRFRftJ2ugnwGHPrw
jglMazD4AVhupFAIER5Wm2pimcqf1wDKvTIgHvKuAABkp/3VRPbn1e8otcVg8rtX
GUAlIgEfeh8N8X+M1U6Qx1NgC2miaSD9i/U6yAJ58jmgt1pBEqHUyFjWy0dzneuG
eYqdgMD2KNE+8mLE2IZaMJUuy9aH0auUzScM6RsJwljVBLoLDLAWJ2pLBGv/s+1x
dO0HghHMd5uGrd49mrmU+/Rxmez29+4aQvZ99Yempa0CEKfDiulILHft5KecGG7x
tVSXrbEuuBZrWNn71GeHN7XzorUk4Ly6mvy5pnUfX+FB5JparKlTzC/qPuV8u0Z0
Zruj0+8MhcB+vQJS0YLaYEjyCs1SKQMH2f1E0lz8udRIFivk91dCx206bvQ+ECiq
9MngET4jT0cnl64sOAGkKyDEjSgZ7qxpqxh244SMGCVliDyV/t1WEQuN4m+QCvGc
fIxugY1IRj0mZeV1FMuB+vnI04JfD4qzTxd8XA+PWY6ZW0Kq0Wbu2tLH1a9QEu19
YkLNFZNDq8eYFG8LFgDtmMR6LT6dPSGEywMcYPnXnwVABojlhsExKO+OinwXzH2c
MeXxThHlr+i06fCIM5dJzplc5ZqbjmiwLCCHK5zqH6Y73FxV6DSHrzxRknaGD6Yh
R8ds0yOWy8+fG67t3SYzaNX2E1tXew/i4y7D66Y8IqQngWHcKxDHg+rY5nh6+FCM
j5vfK+fVfHFET94h5dPXmA5LyZjtjOnTBZOLcpWtj2h8J7Okv9sokEmFaNBDHF0Y
fh2PtV7t65xXpE7NOoe84/EOqO8sgEwQn+6gqgwLCKLh6ge4XK5iSG8Jltfy3EGo
CnK6qdtUj7aQWR1yQeYzbuHyAv2xm/0fDaj74XYawRrSMoXjoY2Sd/ftui7DU9gM
xGhA8Nc7OKSORkPK5/HlXQUFLec3n1q8ukeibLnihu76MjgO4hpD6691WKsqXn4f
9LMfA6ldpLZVNYrXNjDBvg==
`protect END_PROTECTED
