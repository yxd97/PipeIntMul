`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pQWtGis3d7TSH0ikwggSZxK944/BPxhmKxszbT1iGICkVX0qNKMMHRSsaNtZsGcr
Z52jgtkGlMQmoH2S797SyLTnL9G8P1/R0UGqUrZD8NPhKCcJO4waYXqAYPjEPU45
8AozjsYEJzpxQeTX3ChK/Lh6dq9VThTD9ZADpVNDVlDfC/v1U/vQdgCZDdkcx4lj
ri/xdOX9g4KVamTEwTOQFHbkntwP2137GPC90lXlSZW1JsJvIxMPvSWOynjHEqmo
kh0UMqh2MvKCubvjXJI9GxBZA+9GWfholr7Ka44tqnzupAE4bm3/scW3cxUU35Cc
NDiAYK1WWx3cCeqmY4wlRtOBKhe7BpKKOVa03MU7MkJKjygMzomyfO6qYTeTbb3z
6TCqxQnGrm6Ee5opxceURK55SPYcs6QiPYVcWn1jE1HZcEJHr7MZIRAM1TLtbxkk
5HpT8SzLiDvqhlRSMzmPgRb0gqimovKbWKbshLR3RD0ja6/Ov4sp2aorUD4rNXYH
x2Mf9aRQf3trRphYXm3Iy/Sv4CLGbnxiitqSHfdXAVk1qU01+DCwr1EsQDmANJob
oKxj+pObiKVFelIMMCnX9w01y3laQxKbIC3pTQ0DWvuo0iMypEcKzR0OVlIYMEb3
/M4KZgTQ++K7lDYKDWH7thtrubRkp5BUy3VlExA9GL7CofOKeP8oL85poeqrIXy3
FAZ6baFnlqwySZFSeWnAweRXbBptTz9oMfTcZOxUnqQNAxXZbzniJYkNktLks/Sw
JTbMg9VN569/bhMFfQ7aZ1coWVLbIbIk9ysLw1RqEvW8d3TJqTuGCcdIWx+RIbLk
T2BSxAChbtDq9O0R/Enlhi03ur1tAZlwtPIRsmz4ailR/euDBteZY5rk1KA2PkJu
6ny0yWJKY0mq9wFod7Rs1RAZnNXa8TwqXG+mGiOZB7I=
`protect END_PROTECTED
