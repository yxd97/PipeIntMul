`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BwAjNBRk7fLh0rarlqdbcKuYRw3rc/Gu5z/3Gm5AQvUJ9U5gsI0zV7eXN0XM3Kze
ZVjZnELLfA0yT9+y7a+fa7hr+0ZJx+sGQXEPxBdXBkemNitynN1a8fgvbz9Qtmcr
d/eD3YlrbM5nivBk7OQQymQMLeBREf6eDE9X8xArv64N1T+FfQQo7lvxJYUqpAiv
vREeCvsQvDpKoIDShVMroWI2PKm1mI5bq2D+qX/ilpon1G8Hl+nOPuboOGobnE38
7QrnvYBLkDosVmqGDdoFAEPvuVZ0tDCdiVzsoJlCdqce270SZ30OTWV/nZAycnMU
Zn0aO4b7z9aQrbOn17tblCLZppNVo5Q6b0RjxIfyv1lFmaqEEZj8+ZBeue4Cox5L
z3L8ku0Lbg4LpRDUXyjHgIoJ7BDwYzbZTDUay7AZfyA=
`protect END_PROTECTED
