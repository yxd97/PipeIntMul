`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dh9+Ph8uhu9l+w/6GOVxHzhYLz+uhSF08U99AakbZk5GdJSffS/WguidVVv7LFqb
RpPawskzkg0XPnZB5kxvHImq6PXqpCIavT57c/Lm75XyakEoR3bmZR7fT1A1kYJ/
xI22u5vjVgrjzJNMDg2c3HfBFNTum5TfB3hHQrqF6/fOBWqPrmFbPDELOTwFPasu
i2DWpUzFrTNc0/7mNQK2Vw2v3YdOKxo0q1iFWjdOsrWmfG9fld+cqnL8qO2Ez+/1
J8k0Ao+172GT+71+dTs64BAT3GKBIqlhBt1rUOJE9H3g13idRF3ytOklVGqIilqS
N/mCcrzd2zCZDre1mZuu+ddg6Gq7+Nv0zw5G7Iwk8fD2KoZrk+cBfXdt/itb8wnw
`protect END_PROTECTED
