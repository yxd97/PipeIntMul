`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
orFuVk98xpYOY1JbmM3G3wi6hPMkmALW0d3ual8WO6vUAC/Gr8ZNzOITbJy0RtTG
URSw3Wt4MilyWMJI9mPSVM4V1+DoHKmIRzppW7/72RctCHkc0D7q5InI32mo1Uzi
KRMct223e3iYwe4wAUgUw+C7wg0pwqjr53VNK1olEbzgFiIYzGGEZfBaBKFVpT7d
Gd8PjwWSkPBRq90r6I48fWarylFP6GdyxpwYLQLcoUhARLFqNNi3gd4nn6fy89Z9
05auH8K0ZxOVRKuBD8vcicXvWcvO3s7ZWJoUeF4iOXx+Q8EozEA++6WVdL07OwoE
xVgUdEIZEmdIhkm4kSYLf443bf5oKtMVNSLD4/YATZKBsACibwaP5R59yREubS/H
YXOyk6ATwa1G7tdHIfxnH4jzljrkpf1q4PGeVuv1OC+gclCku8EGIzNHTkjUFmse
`protect END_PROTECTED
