`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LYwu6jIx4fcacXKLiUh+7EewrwH7MNO3/62Dnt6P5cg1dhp11yIZjLEsSSQjHRPf
ul2einq1GFFLQXloMYb2F5iwwd2NRDXalL2yjRDQ0wBc4q824fPka78YX+f+SnSO
PIx7Ta0YROFqI0yLuLJuuDN2GfezHuXv6HaSiFIthizXoevCLe6zbbYI4NQ6eFOi
Fs3eP8dzhIgQSFoww0I8sffCDKOWJp7xhCsJoEXv6+0RICmjGA43DDxFEC3+LO6t
K6J+WhdUtcljSMOnZORNb6BW1XyFhWHFcku0F/KQiPA=
`protect END_PROTECTED
