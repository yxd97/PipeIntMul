`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h92BHNH79M6KOy7wc124dx9Bk/zyg5sVb7B5kEjbY0kAkaiRMT94oHA4dS2eYvsR
qvOxN/1mjhI/QpdrFT5CGS9aGJ47vCJQrxoyWiQcQlQHXdOJa02Guh03/IQCHnxf
x/EJ8J4PS+h2hebGRc2uwtnHxEB/nqTKlld2QGpqrMnC8E/SbsvDxcAJ5weMukcr
sGHQ0kK7LKsSwtCqo5ql5/O450kn+Pu/HQ0Q9XbNweAOwNU2nmzbQRxJsx7oJsic
uqFRpicmW8QzyfFptOpKbohsKWZFhT7iFGVki9j6o9FeeCoFplIDFGfBRcgUe3WP
KFJclO/fvMA6GFYlpf2wTzv5uWrJUtCg8XUQjrv9C4uK6pGnM48qNGUWGw2/l61q
1R4Kc4qSRHtYrz6EA2IR+3D9Ul0NkfX70eFMflR+OKH5+3zzWl9SFa6bFT0Dumul
kJvjLWEaKTlhPictHBzllV8JYKm+0XKFYtCuT7WASqU0WD+ODKe4jywTkxTBW6N+
`protect END_PROTECTED
