`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c8nhJC286wBOZ0zkJ51s5wpxtk8HApXdE1J0jNrIamuS5PTuZj8MFAfZJdp2ZkbP
zrZltv470W0pUbU5RluH1pI0OFmJj2KAmlU7/8MAIpfG6KID8QrmxQDUEE6fpA1l
1fcnQoAWC1YVPXqETad45BzajOAtIUOC+Ouxe8O/m5qLr+w0pPV8bgoE06Hd+G//
nNyr03tA32CDVyWOBBCijQy3eV1XL6JTk5grkxZ7MFv8mYCRSXxV3jH+C1cdvVqk
WIV+YpNc4iikL3nPJaDh3866/Eu1p6JDxhO2KrrLffyLdVX+4KZlLVfmoRgRmJl8
rCxG88cw1sgiwyQhtxhw5rlbugrvZ/tTWHS77+LJY/dZQFdLd+1VGs8aO/ZbuqIm
O+ctrPpKZAXgxNumWwNJzy/GSZ0p9r5qHJ849a9T6v0bgyyFHL7R5CV25bAbv0fU
ny0XNRWsFyl86EqWEueW02tD99jTIC+7xyvHFIATCFiAAGet4PJJFgv61Ym2DLec
72zI5OEr0xcAoFWaUsQZu0oDhHGIxqjEp5fD063g+PAqsmppyZ0ALvJwjphoUFqt
iSJr7Z8dwWXeshc6IUyf0p6IYdU0QXBIADerDCnKkSE=
`protect END_PROTECTED
