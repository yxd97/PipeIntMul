`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Z3wmHr1uqNv6qK6B9TlZDg+lB+0HvB+lnKEY3t55hoinu3a71gl0Jv1/p2fIbpB
qbvCpdeSdTpeHjK7coFCTWrsubNyW4T0kH3lOIdn1wapqq2EBoiXbaU26BXHApHz
/V2bGAU8kTQ3DErpBXv7dpbb+TDDuo85itE3QxpwBnZtYNb4CYcTQzQ6SvEJ1DHY
Hup3xY3tsaAlcMsWdqKxbXNHEWKDry9P65M0Pkssfiep6B0PPhK/+M9dC7q0sFqM
JfFBrpxthToBsU+8b7zVltnEvyKChDTGIkt92simJ+545rcQwYWcWFngfpeb4Vr8
`protect END_PROTECTED
