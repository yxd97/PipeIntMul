`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jPyUN9cAPv1mDMWAud7YPnjCnbhm4n3wYOujBxSDbPs+xtgl9hszM7Li/Yp7qq9
O48yN5sY6sW7Z+nUaFT8Y1xOyVNUqafd3rwlIlfmNM1kYtRUmhSdqYSiGrwlrhro
YI/gGhWBap5h++haTkkS/Hx34hnYnHE2zXW4wLgR+5DUunNUV3MsJmPKlhAYJtaP
86/ag68a/+Ex06fm3TXqdztlzbpOYr4RzHXeWlRR+ReNoOAqIkUKE61/4wl1WMG9
d8VtXvq/gwDaLqdLPttlNdfbrRqWtsZ2Lnvu1/B+EUGUuZmZUxjeoY/X6M6E+dVY
C5btM9a9lGTXInCurfGMSzHj2uhkykgzFsPZt+YAQe4=
`protect END_PROTECTED
