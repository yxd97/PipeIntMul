`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HzT6dNSzUmFnNlGReZDouV7DpxoAMRt3kBdv8VA9ss4sBlbcVyPYED4vehoLb3t8
Du/KN6zRuhf/fdBV8kMVk273ZoCwy0kwUrEKcXiQDDsbjO6GivtFMYl9poai/no9
9eg01XIUxOf8GiOdgmpPxBQ7mCcyCUxBiPvwBYU3U0wo3c4+fz3wg29EjPg46Iwf
T6pj3Q6MoD5YBTBfEv5pVdegbRqOn+RjXbgzxEvkPZKEJVLe/4uCZxIRVJbWtLFi
XTJxqKwIHNV3FPuPqp1892gak/TaWOOtYAZR24anknw/Tjk/xKeKxZ08QtH5q1A0
8Rcrk8AaCjJBayyPs6l+j/i1R61+gNvX7qgYHQshuKbetMRBCZCCrk4NlA8EB+Oy
fmquTqAqmKYRig44sG2trr9emm5mwp2sRXvXE953jpnVc+NF8GdLWa11ZMQpubcq
LDUhqTChKx1kyAp1KN7IGj7pklJMdWpjsGpaeZ6W26ar8d66Np3GVmMxmWe1lYLI
uRpSb+jyWemITYNcoACgo7qIGdemVvhwtq0cWuBQHfKktwpn9KjcH/9GGFQjI1M+
idFqj2VY2Lc2fAJs6662Nxg4vJfN19RwC8RlqbANb2tpO8a7vm/ShLxi3erlGyNS
0wXKVfT0tTjymotV620W6rAJe2BSBTpAzhMP/gBxUTtEGCn6TtOezBZbsvpj8+5S
EXJjK0PCVYb/zsrAIB0pBg==
`protect END_PROTECTED
