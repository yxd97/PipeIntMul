`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nQFeJ5RooXlqIW3ybIdstm8dcligswiwD//xtDHIuMx3Vvv+At4KVpxPxpPUOQV+
GT+A9PCcWB24sUPfDFlX99n2BeMtO2jsIid2PrIWBAXFvQpRywgfxmmVsNDtR+vb
h3pTeZqn/yJ43nsdNyZI5mXrW3NBeBBNAijjeirnobnv6JKJu1acuzcTBtgzJy6P
ioxe0Lpyer6+z7ZD9jokBvmc6i5CqsWWcqQO3TSDlOIYPY5XaX05t8glI8gK/1zI
/6QnXFa+NzKSj6427mhtAwTtd2SFuBJnwON7sFXxAoNx5J4XFbB2yzNQKyxOXShZ
jSTe8uGFMgr1lGUiX0Vx7ohcZHk23u43FLwbYnUtaK+EYLeWZmeu36wqO+Mi8FcN
uc6fOrHkMpyTC4chPh30SgoxOp8sjeoOcsHNoqSZ4hZDPjGo+ZgVJY/jzveOSwFR
C4ceYLzOWFzgaJ2zuiBnkI3r6ZLrU/5Eh7/ntmXmELE=
`protect END_PROTECTED
