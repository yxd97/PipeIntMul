`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rR7O35aDpn3+v3Y/tJSMgxDMj2j8RQ4oUgVXcl4dOBRpi+bgEiG/ngFRZ1Reiv8A
bY3P+sfRQWOB7qGXZp4Y+UCQa9xgGyAiNFDrakn9+BUBSqzytcg7A3AGFtqBIyyY
Hqy3VuYgCbc4iC2X52Raj3+M/OrdUo4jT0was535y64v1Qt6+OfGQRKeNCJw6x7x
dUZ2fxNokhhprmn1NltUUIUjvrb28qbfIdJdwOFqRFH/SSIA6KABBKZxhNyOL7mL
VzkEK4xzgipbzkTB+HW4t+kdr7MFSf84pcLNHgK/APY=
`protect END_PROTECTED
