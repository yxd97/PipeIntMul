`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IfFKrv6zADPNSqtLzartgDPF2aXZvgYlHodLHHFgGVIqhg4i58/mbcw8a0gMZeg6
67mjiXRg5Bd+ncpTIMadGGD3rDYqCmSGcJtUrrS1EdOE32zgE7Nq/1kGbQkWjX6P
s5xQyTsGMfnXd0RQWqTnflzzudcfKwVpWIjOwCCNo5zsRTCrcPpjewIc92n1IKmF
hMKblkxuULrpC/kduL1E8UimEqbZzukiz7ca2XQI1kDlwmzRj50lw3GI1ZlHbzcD
Z2wroy5pu4cgo5WUMmFrSxrrW7Q56fOkZRfMhNup3tA=
`protect END_PROTECTED
