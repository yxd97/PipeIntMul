`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lt/rbAfOtORB5XXGe0W1L6bN9RcmR1mR9wZKj03qqQhR/gC60jCa+Paw7J7ljtQJ
POul/7wA2AwR4OpdIOlJmtjNEfe+MOpQTSKsJnN+G9oEp7vdWBztpmwmAytTy2fN
V/3t0N8kXa44vtiUvxDXJlqfXzgaQmB7Uu9GELWe/jV+gajAilN4wVGNwKrhRtbR
B5tGspfpkDnstesX2zg3IfM3zc6v1sD6fv4Ag6nErRLUSka5wHA5KIu00+md92rY
ANtxLHKWVbfb6rx4P5heDilSvqEyhfhCGMmFjuW7Bt8=
`protect END_PROTECTED
