`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RbYu1oQj2Ak1H78ZssfwOvXUXy0Mv+82S6+uzIOe3htTC0cX8bWSIb8n/R88cCFi
nR4EjufBXdA8LIiZdV0UK6zJ8RFrNOIhFOfwFI2XAmWirFSKYkDyqMGYyuHLJ+ib
LVeKD0XS/kSxAieETC01cw6Spb0w2UDxCHr3NivEoxQg+5Tgmn4HbmKNg0szSF99
vito6xmSxronkA+rYIWvSIynZD6USLngM67oAKc4B3r0j46tcy1unbn1lb9mBov9
VpHTCNWhpWXdhW4cfTAZW7JDkAw2kM2LJ1sSrSxy2I7q43PtHP49l8ROEiUAUXAE
fZXnZCep7ExWZ22mDdKO4a7Ufw7zwLXIvmRxxwKySeAyZSTuYz2SfySw5zFhStY9
a2Ln69lXvIcA80JNUtybpsMbyHn74THxQoZ5ziihG3z/ZGssyqKV/6FwFvffHjzw
aCSR3PJWZocsbVxxxtXIjw==
`protect END_PROTECTED
