`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X59XwK4S5qdHkms8JdNG11LyCpFtRpjTWaZ2X+Eois4dL4xB8dt+IF/9+2xXzg8b
Z3MBkHDFrxKkv7T3uM5G9OxWKQON5tAinRxzcOA3DIFAfEQNjmtvGcf9p98MZX+4
kpKCY26odsuuS/mIvliXYPGQVsh1PdrMU19M4LY9ijLKrnpjn0EuVgLlbY4M4FZg
De9011gT2oD1Zp7BiKj9rQPrK5Bt6132f4/m4DMkdWlA3EMpcjvYNjUDp3SDaN6l
RuFxPEIdUWHMS+ekZnlsM8P7p1amFgkmlf2zL0wKFy0Efj/H9rWC4O8sINI/k8a0
`protect END_PROTECTED
