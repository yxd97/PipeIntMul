`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pf/iFL+0WFzfdZxFVOxnEVMaulttNdNP+xOEef08WcobouN7Hn6u0liWIlLiFS2m
Lot2+SkEkaiLuP4wC39afe1UoFLAldrM3RuYU49mnsEhDARo/fC/WgStF4e5hSHV
uiNKljFBx2Op5VpkGVALuouAoubM3XAstT/0Mt4Spyuy7gmnWjXfTKdwsAEkO14K
4ng6J215PAg4owOHtMY6qfdK/1E4N/HB493Y27NEn966nwAC0+LPn1fbQvlG8PCo
zp3v03Rs3dkMsPoIC6Gft9mdqSWJSnkLy7vL6lyg7zPjbbOyBxPyqP5L18FhB3ue
SylJJB3bpI5XCMShk2oB9hqkHtWjM0+lijJ60Qgkk+mhIW8Qqg1tmpK4UFfCi297
k5Umpf91/uPRoRZbh00QHTmgPmptpZTZzAgcXfgooRskwm+PRRdTn/8yjR+r0vf8
x00lSIptSxy4iEyfhx77J5IBGHUqjCbErN9IJ1hnOd0e8iHTK4CdckA74fvqykdA
lRU7NqgqCC2NzMRMgsFjZKmoMLeI7Eh42Nnieun8x+A=
`protect END_PROTECTED
