`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixRgx4T3K3nz5VTYJUSi9PPtHdSk8WWkg2IdYGaJ4tBlVCaIiEimWmUs3RyywDaU
RHOFwvzeeQHRQnHGZD8Yi8fnL7mRN7iWiH07brNOpNJzKb0WXFUzyxyAhBwP2WeQ
JR29glaWEpFiAk0m0aoKHKNUzV/HlAgkLXSw/brpqdYTdNbRzwjowF+h6hyo0TAo
uXOq9VXQea2pfXsQ6tmT4remJ3ketLk5ZoY/M7PgebGTRj7J51obLTvFeyLyMz+b
MAwpPMFatDDgZjBE7+qzoVgZDxxRc2VNYxc0bs8qEKeOkJD6vyA02w4wN8VOU/qd
olJIHYMRaK/eC/acKlMtiJ/IYwlPUxwz/fqSCHnDAFWvSgqTTc5ewpHNmNzMKGRT
oF8zkBcLlCcRgg/AThD+0A==
`protect END_PROTECTED
