`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tejim9TDSEdv/z11BTB95OA4tM3T5YePIhIGGSxkBlaCesrYkGRtZL2v5ZqxUyxZ
9zS9Wfvl4WAYsXbweNKEXNrTX98amd8Oo+1YDdoj2ugFyBuqEVA4FylyXStbNgU1
V0PR7UO0kIyYy4OXBzTKCQ+fne5uE2nusWO8HycagDLU4lMgJ6Z8gbvvbSj3lSQZ
90FkSH1ThtqzVgFZTJlsosKSpPzdvHLBoKH/D4u1i9+hRsgQnElnfJgeyUL+VVB7
JCHFQwDu+8AXuBBsQyHi9ScbHrymPJ7kOiH0cMdr4IJ/gQ/Ht3tZE8Qi18UDB0rx
+o/g4uGr5gYzDz8aK9E2gstEJHmYVKBlc5FSvqEvkfklSjgyi8yC8zvbjoDHryJD
KO2+KhB04sl0+ogMOT9mUw==
`protect END_PROTECTED
