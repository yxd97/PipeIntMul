`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6bTs0/FNr0+4ZlyP7i59yvuV7TDi5m/l3RNTgpYuB/MUbXKQXmw4lVtKMqhL8TGg
eFnqDJeI/qG1IONrOXdT2oH3LXT83tRI2qL5CkR21aGmpnEJO6pADZdDGCEfKngz
ruDAkaE6DplZaMOtCMDxVoOQ07VOQzoExr7D+8yemS54xp5rLz1ENfMAsaZArAeC
KzX6MsorR2Q5cheqLqSFphkg01wVWDXdi06auWladYJcnqQ9LVlCLwL6XbsewALh
pJp3dBIW3IACqxP2jRgP8fipKwf8NixfNr45jjbC2zMmbrLfRKCTTNLXrK511PNW
4IWOLyPik+T/GAPMR2LdKCcdJlQaP1gg86U2CYgEhKlzVPL8u2mFe63cWR/7jOg9
HLKeljkRtwMJ6BSd0TOMV/3+N4pXCIzMrmzofceK41X5gRnl51NE+x5WT50gOh1Q
SJ55W8mwRoYsZgCTSm7F4xd93XWnLBTBmzb2lffe++YKhnGZrZdLAQ9PeQbyh1B9
90o23QAe1JB8IigvTQAY1JL0ZIOkVWNR+g/8wgm9Zs5hMAw90jF77AAk0a1KOY/b
`protect END_PROTECTED
