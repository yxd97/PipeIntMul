`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JY7TIuNTqSo8VBTf+2PYWuEfrqVEwLvPZhiZig6uA3i54jiF98zQdQTU+NzhxTdk
ZzkmIktsAGQIgbgEcFd8IMR6JHNN5ZBmGuGsiAT5XPeklWtpg5N7CuOwn+RvODT8
w0ibKG/tqJloCYjZlnj4LZ3v9M7ofxy24DyU/pYlrBb4PAoIbeuDBxsAIOI/NITW
85W9i2UfFG4vSicrD1BeOSB6WJPgA8LVBezrq4bfR153VqygatcwhwGIjle4eNyc
jrJS9rqVmCujcbOYWjrTklp0RbkfuM/Nfz8BHRVhrpT+JlJhyKqc9k23chVTdnBh
wWm3Rr4O5DDdcjNkveP6gA==
`protect END_PROTECTED
