`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZRGkh0ju/sqtFR9t/ctCIWuA9iDPVMMp5epvrarcoZnuiwBsM28KErvXk14KPHHa
C+ZrbKYHMcaVZAoIVvjaHWRS8wDYQtLZUlYXKACpR6OtYv7GMHWJgklqPqdcCjaW
/7xVzYXJgmgyKmPW/LuRl9+MXz9Awu39BAz8a3gsDjHYXt6HrqKKlElMwl23stX8
4Zq9PPhZyzwBj2rFBbR4adPVJrQ0OmhdWitc3s82ObHlj1r76CoqT3fJXVlowUpF
OrKEvxQmnLDv/PVjypD1KU896DGq/LltnlVOiKsEogyomY1W5T3qIKpMWpxJHCM4
vT8nlWoQsk2UMRwLuJvUHkUI5iBmPtPMOdC5RWX36QDPtmoBbm7hem4R4t3RNqty
ZiT/ULY6ZthR6z51WXGk2Q==
`protect END_PROTECTED
