`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tk95jka7NNX8Ak7GvVClRnP+gzPvUs3vBG14SOWcobjiPrkDNKFR1Dt2PebqSGqL
bO6mvKqtIWTFtV+wi/UBv0QUIf6AH64YJ1fyqm77EPq0O6vvUHnSwMqVCHw6gCkm
aBpjChKYJ6yczExq00qqTGBZk+Na991yIAw+R1BPkH7YdtSooQ/hVrMGwznfc95G
Vo/wz/K8qa2YyeM5DEpp4jBHfmMkYudTOIIVQ+WLsGdvxWbWA13YINZHbx6YBkp3
zCNGqXcDkI0jNkj9bo2amgYTI/W0ys3EqQXVG8XLTZOq6GMWjngZ4UjIh8Qk+O5n
XoNC57JZszkp7U+hwOnZPE+uzi9QYHEKbv0KZ0fM+LDgQaEs7mGzIJ5dSThBcSUL
Xo39BzbGkXFUAom7Le8ULB4C1QjBnY6od1gHGHAdFdaChTIw3/hxIbTUKbUoPkkX
J41vMB0LpiPiUwZnTy5fBVh2obMiXZw2AkNFPEYJEFIA5bFHjcFfxDXpAMXrJEzT
`protect END_PROTECTED
