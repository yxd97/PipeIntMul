`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zARorcKPWTEaGTlDUkyaX/D7Der1MTioY6mr4/jye1ZuTcib2FgGyhvjs0tlPohS
21ECFwOnnn/RuPJyM/RNaQ7krZ/t1qU1OVTKobtBYFove0kLMBmHY1wKSRxwNBUi
I4zX8k9VGce2Yshczg6HtMEoQswQu9bLvEVqNJqSZOwvTvKiW3cCV/wg1i1y4/tI
2hmQTXhaV6JzWDBO3OjQ/DE9qrkcmQ5NY0aclaYVL/EQTJUx9GWAbowHyskvt3Dr
LaVQtz9Vc5PFQ8OnZ610YzhHdPGYSYTI+kMIYsv5Zm47aQ5VxGNf+urhTRmkVyFy
Hc2/3X8DCetSjRfd/wmRc2owLJfG9mgaKID0Jk1dLW86gT5mmFW9yPHBSw6NdqgH
/BCaiPg9fAzD/MgABHPsQI2I6eNVFye2AxTNwDPjm7O7xypy3Jc5rcps2Q1stYOP
lqIE8S7mRij8uBWGqsoveNc/R/LSjO9zcOdDGodQ7eX0wdd7G+56e8YRc6vT5c8U
KdCTAtcQrvd/+3U7inshwZajVANbe4V0POCT12lqslIOHOcta33H9dp4UPhnsdsu
mskLQQVfBHV+FCHo8/Vw8/TW/jIvhGLKnsSizs517O5c/0PzT4OV+5FH6jfNVLJD
+NFF1a4uKJH01k7Oz8ZPlg==
`protect END_PROTECTED
