`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AxP6R7Z04Nqn5nN4e1nWh2U7Bq120qoqAp3To51y6UYqon3adrT3B75S5O7oR/Qd
TMSPlPRRU4T8S1prBHP+xKYcxcub46gKVDcqyX9NFZJ0t1/Ok8lQmpowNtSDB/3F
sBYOVEqdoLISnb6/Z8fN9VnYBuI2KV/uLLEhTVNG0uycPGXakMZGkBaHi3kLai9B
RztLoMyQZerHYcfQWK/f+QUb/CGQdxScYn8ELu2Vc+wwYcgznEQJE6otaGj59OE9
LJtXTrQQpU2eKsLQVA3/YvP5f3azukU5nhYofXvnvvtx7V50XAdfpgpAwKT+N6Dr
l+piUw2P4l1RV8zgFAnGLqJwBk1/jIwvBMzgWjKXBFTuSIUSgoEqWiKrJO5/4j/v
/MkX+VziEcKn1fxj7L+QLsdy/ehQfEfj4iewtF8f3qzOj7UQqPLt9+dUd7znbCo8
zPvQYXAG6ewXCAAWbWVs49gEOgrNQhQae4VWhJb5ObUZcByzxxcZo+AFao++C/KD
PuFSIABc/34h2kCbZsrJ3X7A6vKceDKGSUquApHAkAAWKiDWGLgMQ3wXzHqD4Alk
lxsYs0ds6eMNAK74qXExIY96d5XnRnqQP4cfOj2AflIJCr0SqV5gPrkScFaS72Lq
6zZb9zsGhclE6CD5aOljOpd3XGSDhFhAk9Eh9A2ZjXH48ov6rg/ZZ/szveuoz7fJ
pZfk+RsIqLjcuMoNyxsG9qkvkZheKWew0RqvPAd4bjDsSKIZRFrfbcpkoomA2mxK
Oq92XUJWDSoNGXxqxiynugFD0DVSPcroPxGjxL3gtYskrmnctL8/Us05S6xUm1QM
q0e/zsOodVej+3mOotQNQujgxIB3MgPthz+9v7Ge2KG4h30SbNISqj1cFPAEGqA0
pc+wnJpkROCX13OeG1qbXOc7mU32DBkDBr/4/Etpiq3Qugk8/M0ruf7tieR8/kj1
1TWMYZzgA8+BwmBibtIMY9RLMdik49shB3IlOXH0sCT73x3cuo740iOv5mRO8pQY
+Ss1mbLOF8hNNuTWXQZJ89ODtaTGsMrLLN/TNU+oBab3wvVWvmrNplYIKoAl2Ab1
eY6MjzfMHpHNfGFiW2+oeKIZtYtolmk4eHNwr3JQifIJ5KnOtc2vPC7uQAKvaeoB
eWYkdoeKTyIGfT/Wxgj73c74NqkP7SWYd9H4fJ4sngP1L/6Jp4zCJMCVEBz4VwqO
NQzlo7T55BwY3zBqRZCOHdbOkPDFavk5WJAvjMqEHp7Ql5HMuL013ynC37/Oq+es
YDKBeJ41WxtHylJuP2xL2XKWRnHY2XdcIn2yzrxXdBb9N0c7xCJXkN2AIU8LUrBK
Rp2Rosyj4llhIYTfEigknOJJJ6pzHkQFMuLXQgZAI4FUlGHHlv7GNyeizsuEURRR
Cr/sPa5RtpRMzmJpzp/9HIh33xcB9FHnPxCJqjCPL6eIEw2hvTfJUUwhjTBQEWHM
nIPUgm8x+QhucbduX7NOjB6SXMtO8DGaygbDydmBgsTi5jSmeNIShF4j7LRTH0bo
jCXwD53219lzsR1zPGJfj968uxnH1jR7cZludBM3HzrYbbDvCina1prDvdF96FF7
S0Z4juVdZrkZacYnnk2vy5ajP5KBWQodYCp71jSlXnWdWr98fTIFQBkj5UHsr5qh
0oWXT4fBZ1LUu3nJmf5Ot2YQMVH1HPQLnNrTPpCDHPrw7tYBbLQYknbREgC60cIb
ydSnik60Ta+5VHKEfMq3f2D/3PauM7UJi3T5sGJR5ncLq7GQ3/6iAGWQB2K+qszT
j5euv35ucu2heCA7YzBP87mFu0OYxOgJr0dBGj+r181L289hhMChHf5e7rIKWQa5
U1xekEoKlnkFMEx6Ab+JAW+Ulr7shqNTkQIJiDSxZ0A=
`protect END_PROTECTED
