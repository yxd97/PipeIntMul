`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29bfyDvR/IOew8Xik1KOgBUHbM14sbYtKdQxqY3O+2w3BEC2dkut6D9CpqB64OwO
ZrQzNMkuILSgc5MXxUcShVs87CZWgTy2np+nrO6v4OfmNt5h0ayrKF4WhbQAt6mD
aK7ZFBt6xXkD2ieiv3nYTQI/+fGGSx8KdH+bfCkmOErFuz+7D8Lcgm/fRxi/HTsa
3jQGyhGmy5QhYNZNMhEttVh/MH1ulP5p6XZHvU2hJsUl7QnOxd1EVs97s2hGbl4L
QNZyhmnm2dN0+qpy3eDl6SlfjgiW4uCmXVNGn+m2Fxvjp0H4xwmbAqHoljpdzkR1
0Tjuey+5avNhtt8Z+QMeNPN9Vrz/L5KmCoIYQnvZqJgowEk/1XaJNuQoo29lPqUR
l1QnWLc7H/zCthEqrETMtA==
`protect END_PROTECTED
