`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jt+nogkPU/nEMlpKvylPgKzqFC+LaTDIYR7kiyv/iQc9ZEI5yZK6F6xTcScHFOhh
m62OKkRZs+l9n7XC6ZNDc5l69Ft5pDUU1A0d/H1hwHxVSy/9C26bfg4Wc7ptJGSm
E5U5q6bdUY/bqA81DQhPuvVgVH4JxeIfS1oNJwQrLFNGmpb9hYoiic0xdKrJ0hYE
I443JsxiVQF50boaBL6SllbBNGLDY0GwlfR9R4bO291aqXO6JPa53msiQx/axZS0
sNBPemKM9rst1L9dhCtfeOtFhjDg+FeRMtQs4vNfpwqpM0wv61VJcPvhm8T8JfLf
zB12YT8cqqi28kZdsqzcbg==
`protect END_PROTECTED
