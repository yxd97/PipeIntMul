`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wOn9/+UxtelA7act/WNxGvqNN6nfCY69qWbvR8OFodTNbGrCLIkLDLDyWPxcfTOQ
UCfw5FQaId70RWR68dhYF+iZtsiQm2E2I9uawtObpB2p45ajEwaJEsI3RP7GzUYo
Xcnorwcq7OMqodyIiM3Lm4ScHDCo8b/jeFgCUXlCmWHd1XXuuOnGMxX6AdwA4I2P
Lkctrba1Doov/7ieApXbHOLfpokcJp2KLmybprI+XeGe/iTUgei6hSmaS9CGoVw5
ALPw1lKvsktcBEO/3u0g9HZhcQqBUWNPFDr5UG9tpuMt4ezRpcLxv5xG8GymB/sl
9Z76jhtJGJLxplBctfnFmmYlszNyEmvDAY3egq4qHB9+b6YOsse3kQv4+M0BuzEM
O/cpWd3tuu3wVSi8jQlEwg==
`protect END_PROTECTED
