`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aP+Tsy8gdRYLn4j29sxp+NcArmD213p0cp3WHrnwtIUESYsQNbR9rAEUybKOYIU1
Dp7GsKUJQPG6iRSIRibNgz+6PNttRFIA2rRHrrD9GET9VIA3P5RmIl4V5+XuJ0vf
YAi+5JO4rIA70KO0zO2bbatZdn9jskuJB6cbmhmNnQsKLpeC63R5Bju8yF+OX4xq
244Kc4DmeiPHvwRbmQEtaj9M7SKUily+Wsjz//bZoLFQ1t1F251josvtkMEUm23n
3XSxF80P9JQ+yUgBM6JUISDDHXmon1MIClwNcew1hFBck1Dnx2lpf229zmGQfk0s
64LDM9bDkLwDmIKVyErbQ5NRiPpGzL+OsT34ctFbhqZvJ4eLL4IkLAhe8SNxkZaf
IfezB7u4kTS6a0M6jAqjbb6KhzgmCbc6twTaa/wGeki/aWrCe7sZEr3b/CfMe7JO
ra2o7IGtXVJiEOEgFsy8+W4eihx9Cz01NLlwZk4x5CMj1KtqKl5OHP46Uyn2A9lG
89HIcwGeJ3mStdjX1QWaEWPcK7X3pTSa4aq4ydCglTMKDynnyAW2h+vzqmuyHqg0
pGjPTko4HiYPsqzBnGVuBbXFQ4Q9XlyCN4V6FzUnexv8O7NKauLJAUdFBaQUUO9E
Q7Tsrtc8efJhHVbTT8DQmSdTepMcVt5ZX+9Lf6zv5xPfCQ2Z5sSNZOx7JoVBJl1X
NPKtXRUxZXDvJ5+GPVd2aJwwo3AcIczBeeEW6zNnvMOkuqFlzo5PRf5sLLd7hNUR
fclw7fN+yXFsDRavAZJ0yei/RbIZbi1vWWG/hneHwgx+G71go26tAOqCSezOXvrm
5kgxT492LHMk+ORAJ87o8LcfjiXn7iqfk4pzXtND8X3XQJy1teH2cCSE6XWDyBSJ
sdtTCD8ZQE9UtglsY59y91boTrT33r2290g3MPr3PsUc7Eq55S9YurBPcp/KCmip
dYpyikrFK2x7m8EE6W9J38dXRLnTVkSslFqvnvz8NWyq6OISyt7S6GpQM0PUT9b8
7Q8PaQyqFlYtufivhmDCkyAyqjSrUB3F37HCIIS08v9LRXrUbhLbknBAzILFLYct
inZjhgpnaUMlrYPT4X7Kn+LrWxYFtHJpzkRgS6CcS6kR9nMjCAftL/QIuFFNoBnT
31QEn8hN2LViwbs3q9qF27SPu3NyHOOxWJ6KoQ2FCIK/urXIErN1gyE7Tz1ixXr3
7iuQrtebv0OKc63UGUPN6KlIIOfrQXfZUPEVyiYF5K2gBZYnfoAyGUgMOoDhsD4d
zvNWB/VFwG1Sb+qFYo0FsWjmG5yL0k22Jdo2kn4Qle6eNMK6g16z+zeT1K8f7kOd
mTH8it/VAGdqoDNM7fI+BtMQJAYF6hNiYupUkP8KWPP52OHJbgWu9Q1tipXaIA/n
XYOp4lEgi2zBsf4pEzmfjg==
`protect END_PROTECTED
