`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q4qqMTr7GrZaWXxSEwKLAf/OLaFrnDqOA5RZEDNPp5GM4FeKN30SO6TSnUXoKV78
Fx4rU44jjksztmmLtP3wQUu+Fp3SeBGYFCWsb04EVhtkLmdc+obCWsxhKQEZZfOz
UE1ZQ+ZEIZnABoloMvYE91QjPVtnk73HKm7kljWJBpg8SZ7yicqoEWjtCzAfzmcC
xxCkYGilB7LP++jnNX0qlOLuukvZg5ZqReGRKcWtP82V4ksoj4nUN4AcEw1c6l7v
9vw6NDJaGpJuII3wg0YuRlfiV+GYhvN3gzD6VdQPe3lWqBHk1tU8wjDBqkZvMHTj
0NucvZ7w2mVIZzfjALlK40eMR9PUZ5MTMM2JKCXepcvA7xwx1/R7npReLEZ0mekH
`protect END_PROTECTED
