`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5bh/DvzC4S9q8H2n5emRvfKkQkqRhSTBExpo872uPvdICf6eSDhDD+g8+zh0++P
1GyZ2aSjXbq0hzrhDUic8QG4r0zBbVy2huGlxWnRi64DI7iD3qJ7DxuWU5jfFyBz
29bkDeP0lXsvGetHQfJ6Xt2gb+wzQkb8gMUYnhedxBkssovUTOvyAG49WtQnbdF1
RC1cLvGt9hzCA1mNxeabujNDAQ9/1bUl+tyBjsUUPmu7VD/xNeNn1hHdAc0NS5LI
PftMlS56NMGhTPLy6S8fZZoDbGr9i7mtM3/0xVYpffSSi3C5LbP6gbh1XiG2BlhK
Z1z6KpZMFzuzXoRX4PN+U+2d3VeTgVSvgpiVHhj8kp1VamRF9hhD4o+hTEw+0BNM
`protect END_PROTECTED
