`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U+c8pdhDZ+rdEEJ6TcmBWqVJgzva+N09MBa4HoCVP5Gfoy29cj9xUkaaopKacCh1
cYhJ2bntg0jqRZXQoAXsu6lVwIvlhcYB2LVZ7BnkewQqz25KEUUOTD5bYQJHc58Y
/tuM8oe6q+7BethxBpoyO1FU5944275pPZ58pyDnKriPVz82Wagv79HBzlQIkOaL
aWJOAvVAt+UPLxXzSRbt/r4YiUiE3o5oMA2hG787wpMwtr7WFNOrtzAEkcOlX2nJ
U3oYjpNv5OLNpZV/TQk3I3UanJRhwihO1znbVB/JjZW8NFkcM3O3t0Z8AEatRKcN
O2K0TECu3UnoUbOMbRnzMvI5lQBjB3FKdLNI5w+CE1JOr2mEwBdkXsNI7P4I9AsV
wChnLIfXUDyPo+I+wr7rA+WszdbDSQE2xJ9ZKdym+zXuBwzRuQ3+q7oJacn9yBrz
0RCEXflVfuwGZzZPOQuACx7JSGCDaAxHRAHSy4FsXiJR52vXvY9l1LnXT4H0+7dc
`protect END_PROTECTED
