`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
akmXpB3O/KH8vysdfPlKpBqYm5ejUoGY6klqMQeWdoYlwgQNEY98R3dHDfeGUj3Y
ZsY8pETHraWN38BglFkBbaZfhO+AHzbsHZu5ZIDiw1mAAIlTp/lrKw2xhVanPy3J
ggT1hKQAn8O5EjaxHvmAAMYnfp1kpPRRywb2b74DMxygNytN8gjNiW/bNDvnGbBh
J/1RhvdC95PgWxE2hApaeB0c4bKOzlIqF7msGrKchMYYmmPBlFnY4naA347UUb5Z
SlxlN5m/EuocOvppawAwBSBE2Sq1zbY743T8VRyf5T7GQIfxDn1R0Bg8j0rJG5U3
YJ9eqePk5zfAFNzGO+ADNQt8viC4OdJLszRrvm6IZdGf3MeThuyey3rA3slj1Bad
Tv9MKcMqmshPYuuZ9sM7GMZsF+ArgFVJvgCxX+Cu17S6JyuMfLTK4E1qHx/8PZuE
`protect END_PROTECTED
