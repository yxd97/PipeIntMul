`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eMxzB1om5Gt3zn6YdwsglHYsERw/VXVAzGnuThGTL0Em7bSnskbJMyyjHj43hZPg
tDy/b7+49kax01EPVRixTIyCe7douhg5lDsGFZpA6OtMif82uwEw7LtUHS8TFPBN
RskFKS+CV62zpcrE6JOznnRid/yn/TNzQqKq7rAUBxr8Yf/ll81U2QTkCarGr75M
dWGJBv/cgna28wiaKvFs2tT0YWxy7qvBEmNhAbEiCT6c40NYelwvQI8GnU+ccSnL
XC0oGlYkeeNL6KJyRUuMJVKjrYiroedTZRLLAiLoo43TRg1Yq+qlMXwO/rbZQTA4
rzHs0pKVUqSS3hyIBxfBFlZGUTLlxcLDP/5y+XxycaYyMYJ/bnKCwqQ67hMc9JOH
QKFZdI4XC1EUL9drtSB0VFSOQBKqgUEkGDvnGvi09PrdmrebQfOy85cLYIRR0GNx
hRwMtPTVnm64z3xkGhrqh/fFd4k0079CgNA9BEz4hHqlUP9RDU3hHC2Ce51qLcvy
jP3KNf+nInwLhlCvKacFyZAbi2OujmFrg9eseIlpB4WS8xMFrrzeA/cJ4g9DAJZ2
dkKNshx8qWBw1qsSYXfd4VCXWKrFnQ2ZBz0ebVpxYY7H16W7zbawWrgMxBAIj4w9
GvIEpi2CM98+I94BaYTsuuPad5jYjviMlVmbi/TWBsgQvuiFLm5hv8J+qup2Z1T3
C5DNSkNpVSAwW/u/IKZhokHxh76qJI8x3aFHlVhNdwTibgEBqsM2QPc8sx/Rq+Kb
C7+HGbM8IZFkmlT7NvxcjDeK/KX7Ms3swZ2PAG/o9jbmvquU10Nt8IusnY0IJB8n
PKM8q+xJANEi2C+eSkDv203+lLOTmR89GFW5qmxnZBaJ78SsYdu8LOlROuwu723D
EqwNgaelURVoNYVz8Lim5q1KpJNDZsCQ2/UaOmCzx5oEIKq4z6fSL4KqzhuDjLH2
61u5Xup+5yhXxZ+H+LmzET87o43YVAfI23M6K2SsZfxHEKDtFVkaBSAoPmRBu/UO
Kek/O+Qxtk4MRuhzA7UkZsiVbG4PcmttUWzu3uSNNQuMkiD1BTdC9BTyzMQ0b8n7
HjQ0FaRSIl0YEkeLphyA9eqME1nU6YK2tn0N/FDxkfbXEf8GFAZFErwl/HFFVaZM
ZrisrxMJEFCJbQx599v2UXepRXyv47gx/2NS/q1sVsqpR7wK+Z3DYsGxASmywqqd
mVMjpe4EOlwrO5OWkgMcK1pJ9oqQUBbIi5uw34YX+pqLCE3HAn2F1i33ebVFr2+Z
oIHz6FnU2I/VXfFyZJdbiYAVDHlNlgkvwfdF4LfFbK6kich7E7f5Q1JliTmGjM+L
B/9aLF/j0Z1X2r3iPNA3jWf2wsqV4Y11l9oyhZNhSbw=
`protect END_PROTECTED
