`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S/omZBrEQMmeJTDy3Y3Ql/DVbDBVOwAbluH7XVcdOl2jUGl2jN9ihvUSeRN7j5t9
rlswleVS1xMyBiX2NIyYLmVn9XjNuHao6Io9CPwnZNi9PudPVrgk/qSkwDZufcs5
jPlmw0wt9kWuFmWy0r7lwpZWKRwzePmDZ08iWMrdsHm4feV2u+0U87RLZloginNg
+51amKou7olmtZlqRWDaZbWVFiQSSs504q7sqr/qfO1WLTuwmoYq7WJ+z/bfaHcC
lSApaulH6g4wu95HuvTa4sC5Vm6aq/Ws2Miti6PX6hM=
`protect END_PROTECTED
