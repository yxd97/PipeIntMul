`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z/+3EGkX881u7hbiHin7a7d3gjfK03X3Okdnunzj5uMI+EGvLFjpqDPonP/HJpBs
OwwhOkFTkSed6XEShk8UR6PdyjQN0mx7FhdMOiBHdCd+R/70xm5V6ajoJFYOcAfX
QoX/k7LD+eEiBxvITmB6qWQLF4SY3/MEnU/HMe/rURrdMgxeVfe4XUclHpBVo3tB
FTCtYMuuwTeIHL2IJGCgkeV4pl8mwCJlP+fhm94Oj6BCG/cCpc5mcqpmsuZGWax/
Pg3HbX3UmhqchVt7bk1KORKb6VeDYhlbm48OR38RPcjLZz5AZDN3o7DOOa+Ubzpl
pBrjVjzO+WmxGSm3To3Tod+QYMnNVZPrd+gF2w+uNWFN5oavwYnZA7nSyWDDiuem
y/uRgo1od9lCFFgF3Nu/lwhHAFiC6aSfB/QOHOXhjN/xBeqpixsUL6bdetbKU+dq
`protect END_PROTECTED
