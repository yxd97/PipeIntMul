`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Po5tJFmUWIFEd7iyC3usLgLuEpX3su3Vx3NW3/YS3ZsXe94UNcnx1269ZLcZlvDo
ExdUZKlQO/Df0RpFG2OKK6VDC65V0b9gkYJHHyAtVljXeUKqnK3Hn1XMDVL0eCh8
zp0ir13ptRoFUITJK8hrGXeECiAId5649KmaM3l4LS1aDz3LNpTCneRpOPFTnbmQ
b2lv7k0tv4/p6rDodyvMYC4oI1ffceE0p25VN4P6RttPcwoo+Uwjw///oupjC1YM
E1aIHcApVDtCFgqbraD7dABDfkEzJgKq58xlYYRCwx2CrEuhUKK8SSPe4/I29GDg
StGUR3XoEBCtL1uizNKq4ExXgBFvtWadSTiyKWZE170n4mtprUX0hGw2MkacJtvs
hOEwtDoF6NuCwxPuULCI7ihp4ovc/XAyOYpngQFGUV6txJApPwvsLuDsABKIT1qC
yhEOWxHdNCXv2r0th/5a5F2WXx1JbV4Z56kc+pCR+TQz7jCOr/KiQiIRU3U3oqJD
DTDOqESBcKAqNO6+QPUsmUDWciTdaqMfPCNopaD12gfglkUVpNC3BpL+W4KmH8Eg
Ew/fxKYpI0Xh5pWKlAxTPojY6wjVDxjHaBua7c+gTsMbeMaK+BatrOPEPl+tKLx3
M7frIhBSwY6WXTj1050mjANAUNlleG/Uo4Gd8CXMexf0JkZjgjQN9nm/yNJMeF1J
OawYruxOKJX01Ye7o+yB5+RvIcPxV4emPSY+nDYvDXwNrV6l72JKq/sTJnZmaPZr
OZ+uYabM8BfZ9Xft0TvHBJthrdQvpkKk/7egQq5q/74z5MBVY01fXZet6V+UOFYZ
8R4iA3Iz4RJj6bgWDYbijA==
`protect END_PROTECTED
