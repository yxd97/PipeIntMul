`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KTu9zd2T8WB+G0X0bkLWqVfwm+HgEofVnlW6FXtAuN06cTwrFGrPq5YiMfth61+o
JjG4aiWXSDs7w2XfYAZavFB7/H+6/MFjzraDwuIHKC9pHmAwy1aKFq01wmesVlEk
5v4N0vlALNd4n7v0DGFKVRxPe43dxKYv/F9M3/ehffDNQ5MjEPki4ynrTCbiYkjM
kfLLsc6J+1g7+es1Qe2fPNBfnK6dzcogdS3eaLzyunG2t4kOuWv5k4sECND03Plb
DF2uOhZEx78U/pYTBrToQtSRP3wZKE4P0khy3MARgzOrmsNjAfM3SIcH20Yyx0Xw
kLcy9BcUMgStmrgGPkzYqkYWYWvpl4U61WACSPfy7y7cDNJXSOdMKhrb8LJqHTnC
TfAWjZiQpmgiPSyKu5TMctl+hhxPSIoDz3+tXWobZK1HE0i9q3VMkSjoBDbUBFaE
RAcsRIIqkYzfmNtAXAE2/Cn+8DlSV6ij1wdEXVllA/p29zoV+882j0psQjIrlPwh
MDBgyqbX42mI8pruGPCBGMTPd5E8+bki5w0zZZhSqObZW+P7/lbL5ipY39FL908k
tnKnmHORR08tgFbyYYUfBs1naw1JqQOpRXUaASA/Nx+8Yqxejt0sBj4EbWAESZxO
7OCmjW0Gp7KZHJH/wKWQVFvv19ZIoJoJNLuhhpjp4T5HVTwrLfFXOmrZDECXXU1u
wTYRzbaXhZ3ZO00hyE0yDNGeTbG6eowZzBFAiakroVkzpSy/eHSmeAdrlljL1u0F
PCa+Wdcn3U1tTm2AML/fMA==
`protect END_PROTECTED
