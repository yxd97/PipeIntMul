`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sa2tZQE5JBN1/B7nJFWo4qcuM0sk+WR6PgCNSrcusiEHGnK7LOvXxDfOc/qBLidz
jOgvXi/qGznlDOA61u7nCATML2bn+I4vtlBjuvpFhUJM4JErVJ2lpTRYTGFlf9wG
YinuuBx3x8jmcn8GZtTPAl2MOk6s+/xeF1T1rw7gW9e3b0NevsNb1FC4D7L561Qi
f+yhsYEwz7uyXUA7SuwhnW83lZ0sDTsc071xEoDQ3PaYzq63XUzmgqx1tQx0pfHd
cO0XnMMX3mnHzNHflh3GHt8C8AsHsVJtzx6QsSUxbfF/h4slDe+gZ58PgkCcyTEo
fm4ErD3HS/y5IiWYDzPGSLfTUDqUcT98rmGl6wud8ckl+IJ/ipor9hqmj5SlYTZF
upqQiCQMLSDL7HrCQToNsB9VWhHnEIAT3I+KWDiSvN2b5juDa6/hgkykNcG7sOud
pjCKt376Th41HZXs67En4jMWYGwuoizFTcSYPfNmNoXYXxQfubOPXlPjcZvur5JL
Xcz4OCj/pX0/MvMrukgGV6cj67uHh7u5ciL/k6ofaZOotwU6ePoAEytiKUe9wi3e
aONm/QcGxm1WoHzc3z+o392xg+Lt0pNMQvZd20oI9oajANGsTBcoOqyKeJ8qwJG+
JcHI5Sn905zdWnIVPZExTp+U6O8TR/uo5d2CKOGv62XLAI7+4glpDoKxbriFTsqq
mhw55C6tA0wED2Fyuz2ItC3UckqTe0G8xmwFQ/vsBqTffek8ptkbPBzA8Wg+zYNy
lI6MWfx3jjsFJCN+LGtW8xI9Ehfo8rxvsEOAFwIq+NE0BuOkGjLNPPygq6dJuIiw
xI9z7S/QxJr2JI/aALDCoSW7G6HgGOxsWvKLTIwIq3LlzLmzgWuqrCPIhv5r2c7t
`protect END_PROTECTED
