`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Enhlh/+ryI4au6r6q+CuiSZXsxbDt28Wn5nkw/zUJPmy1RnXR7lpluqqAoN9ilD
pMfGsopcKHq6tbwMxNS+nQAeVubuxLh5zgPV3JFITWnZQ2lDf4mXekdQkKm3S7bT
TVpgDw5UaMzKlI6z+CFby/LzfKpMMy/fdDrjN/2gy5Pr79jYLiTDoTt1qoqgWGgL
C/gqf74/8Si9zA0Yw8HLjtIqaQMcf8yFgJ4Q+/x0ToU1xAFBTztxoOSyOyb18XbJ
fgs8sfvFKNkak76zIpLV4ZebN1coi6EU3xNzRsVIqr5F7ieBRxqqvz7dut3nPmfF
LN500P7bkbnXLQSEIL22LQyXcStPpI5syawzJ93uYTnG4BFoJ6U2hGxpOOj0VSU/
TVd/Ypoo+RtcMId95IshzzRAY33as1oBk9brNqM3z8OikXglDjKFDk3S7t6GFehf
BiAEYqUrcd9weviqV6A/4M9MbpvXSnu8+QAeelkUEe0SzV+bhWkOTzCCmDPx3/nq
JeoSom1iWHaCEYj/5Cef9kvWWMrD9UZmg4diyF/9/CEnK+L3AQQ4Qyd28Ywt5+Cf
AYZ+/FT1YyctILmbeYvPR2o4d8ob0N+K5XUXO8h6TrBcaRtQPoQGFl29SynconIv
ugjIBbZ8fVE28/9COnOPhC4VzWn5eFnTeebB9bBjrqp3mILSadYmzqthX1TDy8Q5
`protect END_PROTECTED
