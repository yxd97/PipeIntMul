`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/75iF5cShuhfzpoazLVQxI2VnSoSeQYEc9ylAx0uUuzwVctCjtYL7DkMV/GFCO8x
2GHT1RawW5RY3KnGG3xBAE1YGpE7SKj4cZ9LmpFEAeSDfQQM6q5rQiMS/TWeUzNq
amNAq4rGUcgloCvOcMjiKzP2RnITn8LoSlxYDdF840ZUAoZkeQGePurj4EqbYrUP
mky7nfb7oweC8s0ppWQYGBSWFrvpgZMs2e9rCaVNGNKZPPLqChAz07z3cfHOPd/U
d8F+/KZdungw1DmXA5/sC9Nl12qUm7irShtU3Yn22o+HbpUDHLz39kY1ohX6bSD2
rGs/nIUXGq+gUPxNHYY4FA==
`protect END_PROTECTED
