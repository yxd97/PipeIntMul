`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68lMlWLTPq/oN0LrxDXF816kPal8uj6XipfSJY1ZL8L7f7rskykI2fZ3R+s/X/Th
CEjxIuxukHo4OOYkvZ6iJfvh7Qk1QoFqSyyRURowTSfnDsSSslQLDcR3V0+jFH0+
9xmSL/nCz5yUIbDn2m1JuWEMFyoq3l40vQubWAi5OqiFgUVpND/9NsjMjUFlaaPl
6YoTvuMNgvhiYx1D5GbAisjHgkJgCb29IVaZt0s6enETQrK2w/4sVbfRzbbyDg3z
WFqRhV3pJhSv9DxQXwdacTvQCB6iSIR37J8+Sxn0PI4/NvUatA1TTJpiSJoz5AxI
BkWpRItcmyUclivgYvdUURn3qwahbxIZIpiXuh06Nbl7RR05lIo4quukuxLK1ci6
2jRldg6V8o3O3a/M4ZSiesuxx54/hO4eyewfgU87DI8FDNq8dSqyuhhEbaM+0EDm
`protect END_PROTECTED
