`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cafUDZ1wck4XDHnlODyjS4b1xVEPbLBTxkbTDo71cn054+qfWGL3LmWB55gVbFMa
30JlP2L5JqEq/Q/AUJ9HUcN/qqUewbOpJWoVYEfm/yPlAgScGKNTwdkvkAyAAl6X
EgL1/9YBKfQ5DZ6VHgwbPUAyTHUEBGjHGQ1Tgk21jvKaGs0LB40wtcrAuMejIBpn
UZ4CsLiwMEsyHAfHr8hIohWTgLrnKFa9mX1AEIx7+q9CNOLCNOSwsv31OH9U45Su
dYMG97Vg68j6Wm6hLJiK1xAV47QayHkX+IwfoPt7ATJ57ChOhP7wPmyFB4JkVOx7
mUnWYtzFRg1Ha8DrVzk0JzWwOtpo558PRjjQMzL/JJV8wdbtpjrxzLUoRXFNpycG
r/rGPEJ3/pEK0QrY0eh2gY3bOBeWwwBdoagObvwLDujONsK14R4CkEdCR/PVDmJO
0FC4avYk3b6P+fML2ESfSnn9YLbdAdr7QfOcMlEfGaKy5oM100u5IhQQUH1qZv6R
38Xa++EJvaYwkTH/dGOOJK1vDjsYaloEwmCz7pMwk9GuRwIry5oiUvsp0eFoWOmv
+1Z4p29tHvIrCbGF6u7ORVKaQOviUHPQWmVSFjypmgl237lHSW8eY6vH/KhruZ12
S3saVjdQWPjMKC+8qSfIN4bf38faL9rNuVL03FKRPc+GmniVXmJFWJdK7JgNMs85
iZKdO6nJ+VphJ52NYtOtaWQIUQaME7B3qqkJR3FCwb9IOGs86bQx4DcbsEUpROSv
t4UdEVyEYEE/XcG9OOlsfN2KikbZzMG+FAmmpATgau4XPJfLFYDa3GKAd+brLIvJ
/yYTC2M5sq7qWBeyqA0Anc8pbMZP2Dl30j8bx60qaikz0nTmsp1wmWVjg74RXSAv
kAAOLQ/Rf10OQHL7VNddoyRtR41zEAUDKojNSGX1SeuE6EVMQRSSMGtwMuKONfJn
plcFcP+KyKkabxHOD2ZJp2BdJxEprYxl7l4Zu1E0I/4cLTCyxs1VhD1A+RFyLS8W
wO6FwPmG5jPQJfYjf0HaMJGXD5lvsbwZ5Gr6DkVwyjsDB0v0ku+Lp8aJsTsiusqL
e89TA7F81gahLzReQ1YW7o1FJwD+u4Io+X200rl6AICdYifdnxR+PEjQbXiQUfCx
Uu+g4upt3GXx5ta9aguyA5/3wbLkCu587YIjz22S5+WYURe4bNojtBQ5hloNnst2
1fJHk4bUZVd4IuhEoY4CzJ4xfb5XwE/koHgvcLy9cSV8viwjx1bLQUE8Cn1y06hq
3RxnLIOgWPV0ajbZyGRcVlt0yAWl0syrkvEzPQBVicSCiLi+5Psn95aQerkPFk90
9blQcB0hsBYHON5tEw5MMyuumDbC/6ruqegjcadpKajsc4nVrhIvKmj7qi56llGH
tSlsunhD7uUBZFGPfNHDyIaNvaKV6fDAhwVTiDUdqJz+swvRmiwvKXILFjYhE8qo
q2nPhpsAAfSHnCvp1Xsjwi6kVIoRkHPMYmAwFb2kMigSAjevv9lmswTM1xGTbs8B
TkwdafyxzfgVsGIaNPFZzYBF6AR93Ez3Qo1gUikZFCBgYFTq6u7BsqHc99i7Ss+X
g+ZZkLSsAL6FA1W32X65bHhWoBWfeHIQj+AbuQ8LmuPg0lF3qPDJvywv/Sq6Xzvf
UproAwqgI6F4nXOt332dn/KI0uqmfiiOSedNAZcWzWRZ1zJClgsEtioM5/bSqRkb
+x37Vw092/j0/aoDHFUnmXjnxMhA3SQLGpWDLupcqffjDHm4VMH9G173OrB+AQJR
poxZE8JuPo28L389roK1+xA9I+gx8hlbvJnNpzLBqsIHn+spT3McpZ0mwNw2DYBD
k1peRIPJZk7gefQCDoNjF+MrAd/ktRLpkkLBq/C+p9F6StUjYs9CUKRaAnU17Xih
5jp30f/f+WhY4i0Rb5M9iyHlWpWUewAU7TZ0fxseFMC8gJTAHdY5BJy8l0JJ0Ai1
htgz2CPP+1q2hnq3n5maOgmNkCHj8pn2n8fjx2ksWH//1SBMrEZEg2Q54UnrqkHA
pQTFkTHbwgv49TPtQE4HbHj8a8XIGya2VDbaKap2bqkcfGVmdF/MhpTW2WgcnZYT
0Da78rdYhCkV+qdf2DwM0eRhS89WCk8L4cq44utKNkV6qCQiMCHL/iPE8S/ONKNM
5FWnfhMYvySQGxR7LbmDWSjrbv+0+n8x+CZe/aHid/+rxm8ynU7/JL+zj7ictKa/
q/rJwcvZYQ73UPxEhNS6U1ILaK0Rlh9L5Wg9Lud0Lq1knUgpXVAwou6J3xO+ZhOB
tPR6rVX6U2DzOY10bPXHEAEPuZWdeKDucwxUaVhLT015QaHWz2KmjrVNB7L4QDho
ScvzvjFymDIlIzF2/dR/J81oyyxjoOWr2KM7NMZhHiUW92KtCZDUqxIINtd3OPQY
km00P6md1A2USW9IizWDOFjnoaAGFh1wHWOLIpeWoykJnziNR+/TkaEGGbCVEVPt
ki1hcal41dUrLCNWrD38EoFalKwPn9blnNB4DeN++LsTKCOU8TNSV2rSfjAbZRrm
9jMDeUteCyC08HnKiSdKwNQRBse/vT0HKMG/ZpS0Ql/3mtRdpf4XkPXrDBfKQt4g
n2JN2Et8rsSp34Cgo6gDaBorPYSuBXWiMvX1w5un6VfdHQHVnhbV+ecLlnKLqHCM
HwrISGI+kfJEkr7l9sUnqaicLVluDvNy8ms9io/Jl/61l490XNMEMn6UdWssD5e9
13YHJeSwHASuyhYQXdjOCFGD7+3D/ZMttbQYY+6g6P0qoL7aBrK+2BKGNHPhfEJe
NPMZfmEnB2k0QtJNDU2qM/jefvAE3wLVGqF3cGNZYglA0p20up140Tt2YaKrxvJB
VXbrPR8yaC2IAdoOJ81Zq6LyI8cY8dH9iNcS1rP5d/MzyXdDMjdZK9TVnbpcozb5
z5dx9tvq/AfJyjjf/2+kkWSLX67yFtuRe30rVgC2wLdLaZq7SkpH6j4HqtAV/74u
NbhFkRPe2RIOYft8zml2LWjXQhPWrz944fktIFnVTW3XlNXV/dEDLhN3mp9NADSF
Ag/Ewh5Oko+EW2s2ylT+pcG3GBRi+BNkfJM0ESAqzOInajdbTKyUlfcySKST48OM
uYPvf6bXBlrFAniNp1RbrAxHH/Uu7ApOxrIOGG2Xw1gn6z5863CeU2uu/0n6pmQB
8XucAs4WsVd4xOsmaHod2cCiQLSVbvlkjtmer2oHA/7Tphj3hg4pDhsq9cQSS2YG
8BirMbORuuAuzpZ+R6znHcrIllmvF0twUO0sDU6a50xG/trz7CauyUqQUCVL82nf
IAdPQys5JA63CQPVcLKCL/DCdQURBPez4Z3UMCu6trdyf5+FI8Keezm/Kyuo6B5t
JZmhWK/Fx1kM1fmcqRsU8fbjAwexavcAzbUOzDo2lw+XZuuOAx7AuT0yw716egYK
BgWBbfLAXQ1Yw1cP/B4hhzZEZJdJljh1HcQEZDcTJM2pw2M06RmIEPFmIc7zbeUh
qf2clYURvDqG5gIViw7gBjSax6eKyJyk+ushn1WJL6vK2pjJwluv0S91e+U6Z4+R
KuhxDc0XEf4BGeonSFREDfPUHd3kXgnOz/gNkt7ozu2b7KeqFiacPgQOVZgva9Bx
9U+zGlfkdl/00bEVl3DhAvGq+Ex0aO2p1Jt+vXNR1q3sVc86FYE1S/yHHJSc49d9
fPzH3hrmM8TaGs/q3BzFqMcQgum9vXuaiePambvfB8r9ab2C7JFG5Nvb1hDb7Rdh
WFpek+Izc4/ZAerpv3UQV+30yTCJ0fxbr4Wp/aq7AU9rqBByPbAKgTdvO5Qnu5Jn
InyKjB+ktEr/GQNzjWhuKQuHTv3LEaa2I6mpyG7I3rE3LJiL950oHvBL5A9nQL5G
Gz/bmzyundxUotfGzIScrTqAG7uNc8tHCaEXozSj9JtZ/yafv8O1tCOV3QkfdF+R
gqX/eOKzAsun35A2SYxBwEUvzmZcb/JYGh4dVUR2huBnX2uyNsgg4EkU/q4/B1mq
bPWXP/xIkbQ8o+kZ/ZqAhtob3XUMxE93Urzd2KoOHntmpq4S73YQvwH2FME66R59
MCg58uqqaJ6hWRFlH+QLwuDybcqoTGjcUbE8+JBwWY4D3US7GMT5FZfTr06x2k6X
CFJK7YZBW0fDnlu5bTakDKsc0GF9qgFEuFEZ6qUEhyaKi2LyLHwtcKJ8d3vKHrNn
iCcf6EwMYk9NscfzW9c9G/sv4e84X5FU36YVKv3nJyY82NU1lnT847KtMbnEGNTn
nFiwmfDR09HiTaZ0dRM1TrMGgdcW7Pmmu0f5JpLkx2wWLNmcH9lk9hPw4BIhwtwJ
LBsp5QGMR+duDfTA3mX9T/C8GMuOKHTOEB+L/7+KjNnxNE+/p2zz+ppG3R+T1NVf
TNJmVLt32zA1pnEtTpPS5kekIcsti1TJZjJbbiXzsQ47ZVwDzspPsZFZfDUdAJ0K
X1AvdUUwzkNkOVZKabPCO4/3RY8AJw5my46iq4Cm8jrW/AjVP/1grAK7FazVqWBB
lkA0xASvHpALrtKEjTCtPFMbc1G/JV4vbesSCL4YDUjaX8vzuBFV+mfGD1xbUTEW
bKwGE6wCv/am606yw1lksNKJ14HhxF45Wl8MHfHAkUtdiLK6PUoXhrodmT9sxTaL
6bJLqQakCo3EWEVSGtRzQiBFDDZpfmyuC0ovuwAd6r1wzxRAiDjYzhUWAg1ahNeG
LuzjxEIO4FQlbXE4OjPLuus93i3ogDlpdGUt6pzMwp4GTR4ihu+JewOylPXpH/b/
6ukl1r99ruA8WgAbap29vmNE6X0IiZtwXWv6zrsRe07jryhIIM3waQfczHTUgaMw
jAMkR2vYjOBfJjNEfx1Q95velvtnapS9rAlNXzppHXemdf3trkktTm99gJA7hb3l
F7Gw+FxDbqhrI3Sk6GqKQs40NJq0C5SUu4bbfBoLTB1cTX6x8xZFGD5RRbO60Lkc
HH/44YLl+ttZ0csSTGPeCMgjGyfb51N5LUErUJI31AZr0LZCEo99aKAtb+BSBG5D
/lHvlIZS/iczrbTwYBHN1fMqWqniqM8HdcQNq5QmgB6uBsyIElqbyb+F81MdXrja
xF+S/EKSLXpyLCUDPKpEjulbjWlaEJXVxOUwk6W56QDc9KUO2Ie0tm2IgrD/q/Sk
Y/Qk86kYg++vj8rk9/3eLY/4ifdXx8gDMkbrXK6pDaRkaKP1rLu714eFP75gszIr
LraP6ZcGDTuQayV54nOkLuT3RmWHGoQo5qiroCDcijplyxLHKydSR3UwBHONsAF+
bxqYdn9OERS56ec8guwj7K9vntkUmokBVd8yTKawP1GFpJNJ7FktN/BuMbZ3HKVo
U0ydd2Ci0iOyPl7bFkQuLjXKryDLASwT4Wsi1HlgUVG7TSPMmHigj5n+a1E+FliD
qu40YrsqDwgSWZ0qQ3kHeGjKNfYT3gj5ZogprzXCGaHkO00ptW8qClyPQW9Lt1s9
YJFvmFNOlNxosBbPSzUudIULVhH0R2OLlZyhyk86a/fSgiDIf52lyMcilBRUV5fL
yUS9Oa9p7gMpMEenN41uWoeXtPxLFp54Htg3v9KbJ4gokEUfej1hZpPHfn4qWIW9
IVzybW7h72JiUYw3FKC2dFbCZMdmYqNcnIBLjmV5QebCIlY0WC3HxnCFSQusdxyQ
bwzcIivNejLasH7ifUi9RcInsW/LY9Tsd8XaNpcH9N77VVZONft+GzJAwKJ2lrGw
PwsEX3TyGCZvYaK2eQGG87Mp6qIi6cM2eJNNXRDuvJWYbRzk+mdciCT8CwViXf7y
pwidh5InQYiV8JKWCiePr/Da01fl3949jY6wqjYwNDIo0/qgSLaZ93gwspKkYxAv
pjiCZBAu4b7aD3/DlBsd+py2xeER0sGPP4kvTf/teE2XSLe7kuDcCLf5wNwNUPfi
mXUqJk4a9+IGc4d1A/PjGjWynQFZ4ztt/aZ0vyBY0qCNO4g5tv1gmEp/1jBMqY9h
J6Tuj+zTN7UikTGWn4b/iPsStzeIulJ8E/rh8xuR9siCP8UTtsxzDGxgQnThw8/l
B93nJ+Qwo4qPl4C08UteVinLmxYK3H0xk8MRrC55zh7iJY28f5MzmYfpt6E2t0Yv
HYTEbNQsYqQfNiMYtxaPzSHwu5rlghNkcfuSbGiK5icg5rjnKEL6bDo9bt39IHJC
`protect END_PROTECTED
