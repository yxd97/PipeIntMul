`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0wZnamUVnkum2EExCVBLv/neIwQtD4Rfc/jqi+5inMUPKJHTU+ND4HF5yOcqAwM
c/dIcmtLb2LlRtPISlM+E/Kbiz5k5XEQAKX3H/+DrMKWWhOW+JwcZfzD0dlmfdXt
iAqvM+ls/aQCS+9De4V3QfgFnIyOYAYmUxu1kTqZ5YXhS14BORDq+HK41Lva8zEq
8X7xtW2jzZPgN2GjZa+xRnN6rwvRSDasA17TKAsfPoMFTWDeI28NZIFRCKMuI/bc
JIVqrHX99lJWqyIBIT0M4ZznYyFEP+zj+BKCfH3nLmzC3NNj0JrWGsqXZbRBKUmt
Nit+e8A02wHvGBsczFg5SQB1s6s1FFAcRkPfl8UMNEaawdgkZJ5Lohnwf9kXWLqy
AmBG2R0JKOoXVPByDTSCBWg3iJFKqFTzYql0xY6boGHH/St0tsxzORQiMi+fkY+D
8TMH7KOrc4fLAJguBiXgThuYLqmqkgHMJDbtHlpBwfD8/LEz0SkvZ15fF8Zj4PcZ
qhlUI4D/J7XCH81Z3Lfzj1rM4RX/itvDAJ0+Vr+sTCy9scshK9BqtHHQkqFwznyP
2Bs8T7MwDMxvnSlkkblHsNAxmHSGaXjZuQIVvsSsuK5+AL/zGNxn0NJWSXfHlTJV
3SN0j9BUZUuwgiPpAWcItJSY4dzs7C7HWwyWocGNAe2Wneymyvzsk0szE8tnAdLH
hx/rEonNAcXMPp6e8LqP0W2NaTdJJbxPtdrsdLAlNZw/ECS0L6Vden43WzETdWBn
wNjajd42kNJ0WyYeeMuoteBT646H+vwCsGbeXrMHUHmnmaZ7u/QNfdNAcH2YjkmZ
UHHx/8tul918XE9smvLi673TPW2tIXDr6TSsdnpLJB1xzT3KDyXZrIu5M2Iaas39
OVfjgJre5BBazxJUIHuAXVZggcfKgWbtDBhlE/NBTS/h73z2Fw7FT+yBmcCfgeeq
U8rRIf0+U4PaM/V3SVCU3zoxPxB7tJjp0SI5+P0FRyqF5GzoZGZJt97wG793DjuX
`protect END_PROTECTED
