`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E8m35/FTan9w74sFREMz6HqrhCcsOZDGmRY+wfg4r+aNrew9WUKmUeCI6G9sVett
7QeilNKFnlrdbImKeJPusJ0yfMYMtsO6iklFeiU6mUo4iqMorZM5B/drhOns+syj
Jtv47Vd8tzR4ZcwudkS2vNEh9+hmcWB+UVZIQs1VldViKYUW9ubxp/4IszuX3YAj
i00sQhlHU23gWbT1jRsXpiyLm0YUgVWzLznBrW9PmmSakw80EaoBPnkNLdr8R8z6
EOhflBT5FJgq+90edxio4CRrK4lCOuVWwYM9NCB0+G5TorW57UnYJ5dHNfASqfAQ
hXUPUee2s/NcYDIYv/VUKbSI86Pa4lARgS9au+RWx260Q0q5zB8BmM0DaJsvzVvH
QU6UgiaaDjK1pUsICeE1Gi5Wsxcwijx4qRf0+GyPK7LD/63hXcR/gCmG2WiMx+s3
6XU+pl151MjTUW1+/dUufCFqxWt9ryazvtFRsitTr0wDq58Z55OK+DPPEdQ0zMpF
ggL59hLVvku6AuMdnP5BU0Yqva+MjGPUJ3c3BBS/G4DIwM9QIJ/E3ckpRmEOzVsa
`protect END_PROTECTED
