`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D/kVWlYFUsMjZwgRSEpvGnkh9rCZHTEg9lLWnEYw/dO6AU87fN13SDaHpT8Sx/il
9k5SI4fLmTBau7wMQozRmukgoaovjhFHMiUvZQF931pxAdTjvdI+S8bWKUVfKeqb
azCuyTd/Dxt5Kj+s+MDeP9AVBUrsLUpgLrRBWeUK6NNd4Fm0w3nuguErnbxDLZKT
9JU29EG8mJWHW0PXZ1/Zgiu2nWvsn8KuGZOMQmcoHKQE5//8b1sBEOt+oypehLTJ
xNq6p4Jb0n/vZLYlg934HPTS6kUpLv8h8s0XCvCa8y4Vs1gQWn/k73c2WdX3KBjq
lxjeia21jlergHQmcvBrLreo0ho7iz34+xbRxQWsMqULlLuL2r9SGArnH6iXHQ/O
SpCe8zzlVbdYtQQvYBkJ38ihiloJvDLtgQiLmTpRw2ykDUZTEiWw2UZzLESYWath
q5X26AeuGYHAUgvpR1YY52ICWXz4SVoAyqNydsoZYuINZC5m+QqIy5rG+TQPY7vL
CgEiKgDqALaNPv3hL0FVnBktr7XmS6GK3zAyxA3OD2WjtlRHDwFIhyGmn6TUbngO
7NxiI6lplWLjXmdDM+tUYg==
`protect END_PROTECTED
