`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
au9LGmk6PDA5pZZfaX/e+sxt8xD3fEjl3EbFjc6kESrCLcUzXbnQeNY3Jvd1G5d+
Jly3ZCpXhLSWHO8lOQcMHHRL/aFOmHB1yk4fn1kDbJk/1PDKyhoEyhDPaL9z8r5d
G26E+nilAyboOiliFd1hgfjUqCDE6FkDGJ8YO+RpW6fFh7dhPIDBNgDne/mG425H
sJ1/RizAljdFBhwYIBXnrjU4M4ztVdDZVCoRcUN0LRhhMbGyXVJCQR5bogMFvwhB
cA31LUq0YVVT9yjuI4f1+tBINhgdRxd+fleJfv77EnN8gfwICsqzKwF08lJREuHO
BmyL9U30c61IUlCNyuV4bcoTC8XjAk68mLh4g+qbqzAiwDjSBv72IJKplvTZx9fj
9wvhA1lW0gQGaDJSgp8dczspVVypjXnsFvSmx5dvgrU+ULw2NSY4HIaHgZmkJbLX
NIX4cVuSN67jsN6yH0B/sbc8HcQari3/YSguIiePn/YGPJPQS6BMydBr56qIcAlU
`protect END_PROTECTED
