`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XtCLg2vmWy4IeYP2OKiBV6Jl+yaqkOwFUAFPcJjH1wYclotLcNfO2r0hEJR2eLiQ
iAgll6js8mtUdKO29Hvz4D1g8PZj1dftcusmbzD/OiNG+0Bk/3+uSx9Z9/KbVvut
tsvFS7D6d63XwXPtB+fApHBVIBDn9mAxqZRO1PBHPrhb+Vkts5vHtN8eyth4f4bk
C+lUzFIcHKddFkW2SPoRtcl+cHTqq5EWmcgzGCE/BBQGfdA3+ZRGgIYcj3NHg51C
SpJfcKKNDV/HiHXSREO79Ph4hBnKlZzqMPPtkhujUeYCUP0sDkXk4LYvmlq3/dLW
e4XJ4WH6dhCYh82Hnp8IyO1VBc9h7lNF6iR3uZi1ib+yCMVAOyVqtFF2N1JbQuoh
cbfLSir/xLWzvuY8XZCGFEGGBMV1+XnJ+4a8/YP1dUaUbhS+vx55Rpwu/4IoyXul
mA5MSk1G10avG1Qr/+oU/aqFRaka9z18wRDij5V++/aHfj/2SwGHGTxF+5y//RnQ
M2v9x/nx6Uc27CgXIM9siK7aM7OaD5EJew0s/XFkaMYNtsShIM3pEWSV06H458Ih
lvqMA/MRNp/3OUHKxDkQJg==
`protect END_PROTECTED
