`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9dNgUFF2I6Zj0ejhtecVv2OPMkjsWgGt2GHd1iwAR8yi8R0uoFZW7BkfxEhTgvd
uLNd8nuQsz5Gv1vKuSVevOfkmNPkBzVqrxqqzlzlxGyHW1U6YyqyTYZ6SxV34t1c
my9tbHKxHDNymJqJIDKchZ8ooT8Hb5IcyVUPLOvJSECZJchXV/vSMLpY0X1FgGip
Ny3QM1j/bzjVl5eh5JPiAtfikOchSxfhVUDuk5Jky78yZHr/of0ge5vYYYoYAtyz
/TvSAnnCRbQYC4rjsi7tbKLtCwK+yrLOuSc3iqBfj7Us35nEup2NTAkPxE6/5prH
`protect END_PROTECTED
