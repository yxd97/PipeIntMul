`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nNGBWkSpXUKSZ8OhZ8U5gF6Ng+MWDhYnTyQgTBi7kXnWX9omgRkzfggITkm/iCzo
D+YJg/8QIi5+1itwQ12BAHVVt1GcEOWzjY7RhjtreYxRb2QuiUnK2WmjUBXoZHAh
fjNJ5/z7X19BdMrqRVVvUOkD3KGfGH4IsSOJ1kfhFjPHtTrP3+8qs7AYfINge1W6
9SHjdOMoqcV+KuQvbtvvGDkmCTiGdsm2ysZuI3e8/f7ya/o6brgH1cVVfVbtKCLi
Rv6Psqb3fQT4H63h2v4rQqn1qfYJG82ikQj7ltVilJ0GjMD3dehKEbr/X1J/RYPr
Sp9kC2ranx9W9zl3CUpuB6EVI6SNiBuc+RoD6g1ZQgrO8r7XlhzEiTRleUhStt+V
O5KRilwsMTMCp5mr+ecdmuLDKMLMO36Wlxp8t08MksEYCy7mEgVtMtSzWaPQCnLm
DiOx1gn/wbKrQzJigKnZu5KZyo+o4HfSN/hXlY98srGOKj58O4V3IX6mno+1vBJM
SyWpCZIwaqDXwjsbv0LJOHMH6QPLQZxj36q3L24SBu9jNY5uJPZhRqu8UyiBm192
v7Zt3N23DbwubFkTIfA3XfdDfgzSTP28NLSCqRTbvLziGMEHzqE67UfU53KETs6P
GSNvXu9YRAq7CWaxhwwZAnSoOx4g/24efQuQ9rc3SqS71Dy/88aaGFfAMo/lSUzo
G/b528lFL+ktYqq+co0o/Ymn9sg8DPoRDAGxtQgYoMcgVxaJK+ckanrMqfKwh7Sv
/vrrAEfIvIPpUFnM0NwMPy7EY9LYtxcvULts7YOW2o7nPo9e4SvfC97BLCMJaUXY
1fygrp7rLMZ+Dy99QLF9XxM7Q4vMTQw5wSklrdhHSeCC34S4J39B+YfwM/0s2jvn
0xRir68F8cSX84BnKTSM3Klz8U/T6iFLIkPosNT0zbb/4z4MMbGAS8WjszMt8uV5
bwI46VPCnOy/+V6k76wbF4ZG1O8zxhX2VDzMTW6wC0n21oUl6CBTwHd3bMMueGqm
4/arueALmLtigi+6vncRAybHhfMpdssxg09qkj3ist7Mv6WVA3tTTZvebFQ6/p4r
l6N76/rwmElmbIvEjjzLAa7NkCw9/S+kHSitYFvaHErcQe+9bZ4Ysvt5v3iQIYw7
7kfkD3YBPgWW7skxbEfHnKknYRcOlu2Ign1a2pr2DngbtEFT3IMRxtV3RnGK3MDR
x2CMr8YRlY45My+Qye9Upe8ZBTI9ZywjQYSVJlVKbDxYvvtbEeSZwub3SuIfNArN
t9Zg5e+LBHXWAbX9/aGN9mfZ48LKFEh49Mq6rYQiIj8u8pXZUfZzT/JR8fxLxMQO
4G+njiqDCoNTWpuf/21oEc6h5/VPvswLsL+tdvdyoPo1owCND1879SuF+6D4kEi2
C4yDoJuMGxeVbNDjSRx19EHsfETpNkOrxhfoaNSBDUzVGPvl1lz/ly3XTB7H9Z7N
sQjS0063h64i8bIglJvANJgF/c1adS4D+ZLruC93ltu/mLqXTUei+aZ2cDM9mfsD
1+5RYRrmW4G6TfK/Dcv6a7uPAiG5bBpbPaKzHJsvWRsoctZYu95OQQyHWP5IjMIB
4V2NpD0X29Jr0VzfBzCoe42ShM5AXRnc3YyhbPKiSYN7DItJx4ump0cvANEY5e0r
GAa3mf2DF1ojGKfaX0YBHVZlf9j7D0noEovwi2xEyYgN7+Eu8mpKgp2fJY2BaS3Y
Z5slml33zZtdEGdJDxY3dwP/YZXnNmb+GMo6vGY9SAGlmeI0iu0k8u3Si01Y3458
1dqi5D4XtZXrfI6+XaK7G4m/Rui7KM4d++AAL3899E6nPmfRYIxZSXOCuSZ2AQMK
VojA/EoyYQ2rZtDyf1/R3cgjcJi+bV2t2EGdb5cqatE=
`protect END_PROTECTED
