`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+FC3D6G961jRX7Upj1zeZydhYS2plapqIfTY/Sp2CGTLu6nKbouyKJYCMayRcjT
Rlo0R/CHgtAqfSQn2RFfcomUEAk4JrLC+OFrG8ECicQkUzW49kkLAg6D26KlY0fg
OkUon2IpjKn6LRz+JEnhIQZp/Tyll1lRGWXX4FLJOa5y2zFsz+4oYDlx7sOe3Vyd
hvE7CkhCxo2oZGseZySk3JMdN9dq5ExOvuUgOazlaFqUlU7Kho+TrSAkqfPMUHA+
xs6r4D9ORXr92/jtEplR1hVjXGGLJ3UkiO8eyy48K5bnDRLRPbnylgZhjYUa7nUW
qt0HCT3JPZrXAPwf12+DLQgF0e++bq80QLworOUJFZfgRNF2vzWGxfYZ8ymH5ieE
rLAFPuK4GRW05Jm2Im9i3RqZfbrWRlsP5eHgBLqKf9+ZbyqS1/E52pOffa5BbKKR
cjsHcWSUpKDqZ5c1IsZaGQ+rRtlFubJSvJ7VT1RKLRCx5U/eYp4xuafle/W7+5Ym
`protect END_PROTECTED
