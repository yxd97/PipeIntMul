`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Icmo6hNO/DOmdeJH7FQkZFHdUgqj+0/F80U8HC1RLMz0oPgC3E8eMktfiqHWp1yc
0hNWQJfubigRsr/rLPHXtqbPwYDVmzzf/J88k0/NK30wtL/I4zLQvcDHxggZyD5v
S5oobkGirmJMV4qMYivoIstjUMq780EK8ph2TvB5T2/UWa8ZGR0TBdj6N5+3Ekr3
VR7qedoG0oJ2SbNNdcXgWd+TMPKRJRJ37xuYNj0uwXbKXmn/iOYScJpwrg2YzP95
kCpKMnW/F4qNKBxTnMHEu0qKu2KfJiERi9IbI+aSJ0eyjDesJD1F1LAcgBCoAYcc
Oc5p2RQs7NRbzHAkW2BHnX0KlYnW+fX6ghrabkfiy7ESyQDFNW3NHU8xn4xDf52d
dld6ln6493B0UKlThG54qiOfEofj4ab8zPDGY+suVSmybpmWFEuU2dBDtEisDAJS
k8JG7bSlTeeHCWTKkssusrFjxGxLR6tplbDWXfMZdi5lYNelcKamfFyTiiCOH6L/
5sDfGt0Vw5O468mbc/r+BoLi/FknbaguKQrqaj3l2eVsCNEWTEETj8vyyi1Os6+I
eogw21cSrv28EADJQ0aOA6zvNgU0GTXFTLpqBNJhC0VODoarfjij30dK14UGNs3k
RVcRp192vO1XvmYaEcWmtUACMYApIyIxQns1zl1BWhY=
`protect END_PROTECTED
