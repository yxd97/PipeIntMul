`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kGSmO14RlaKECv4+iYCNdXQ3t7Yx8QxrIoonCvxqh3RWgJenT5BLkoUYX/12tfCN
mmXpo7b7HeiFryqMknZ5Bsxl+rdJCqH47/vN4VB9c4gVEAeyu64TL357Ok+YdEw/
v+AODlYlpvlRd5AlwvP2d6EUndZAq6DTYQo5wyOLtlqZdxDFIXvPcsIyCp3Ac0eu
XnNoy4mtEfH86HhtEI/MBbtaGzd/G6xucPFVzwhKrP38Ezw3kthPYDKPRlnaEBzw
kduuqU4cBDW16t+aQ8TOFpcpyhT7AUaSwdJ1/Iubd6Y5zb1UCLIxKjTIKkj62PL3
SlM7cfzfyBxcKQhhq0op4t8DOB976dN1LIZRXvdjZipytWr3iLYl3fD1MkSsMSlC
`protect END_PROTECTED
