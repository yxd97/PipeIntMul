`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9SPbv55Kwspt3aPUWTNCLRb1/Wk2L+egHJNvBHNmyto4F8vQN/1vBh+fJQYg8lI
8AmKwOQwSkasoaCxxCWhXxR7HfGoMk8qqmxQgSZ1Cf5zekskVRtbMy3EHwiZ9n6O
Q/JgyKuz7WjYed7/nbmxjzXU7C7pI8oDgCJryzdSxklGu2HY5ybJ/5i4bVY8H/rq
Il408wxpXgNBlBrCcePOdBof/2FObLHWwGB7GGPycGh/R27JYi6a/Ii9Va/sKo13
l7p2JY6CSGe6Po12/rgeF5rR2R+ioNH+ZcqeNzdLevvlGChbf6hchTrQLY0lDef6
Q0LGdlWNJPwJGNzAOfs9NXrqePqnZIJGUaV7MSi0CgVNtguvGceiQXxy6QHbUe8H
iHLG5GeU0mq7Yyd71E2XvfWVhWPRMEEDTapGI4h91l5qIam6/9Vr4a5QKjzmWQNo
yvkPH/iM1rGG0eUXI3OOBUmQGTeEMxtytQpf+1p4eEMFeJ4mHTzluKcWQUQVaa2r
MJy4rf2aM+qrdSVhhx6hDBzqYCEmJ9HuEYVbwIzZWcXJqppTUO4Z+Iu6Lu/CglUa
3AQw27/dwtMu0jQYzqPVWQ==
`protect END_PROTECTED
