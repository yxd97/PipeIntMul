`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Unxol52rAog77H4wrfPMGyixPMxWuAWnGRWPYV/E4F04RCyf+J81AlmpQicnFDAm
GY8OTtmn8BYKVR5qoFGcfrPXxe1yf8D2m8fZ3LFmJEJWKmH7IksYk2xGU2pa4H/m
MJKqjlgwzOarFjFJ0M/W1BMTIWWZNlud130DxsDKiHhTIdfB77lMEIE1WTXKF9Ii
Iugb63bMHo947DjUMrjy55LOSnwPP3CT3v3YD8u/OtlBQ7PNFfQCWegWIS+M2T4H
XRA0GdR/cfgxbKx1OY5tNvJjVMfiE354HmD7Ob5I1lBm1s9llriHHHAmiI1g3fCE
x8c6leeC2uiOrMclCF/mOaXozgqX1fBXpLQ0f8QWeGD74iO6RMSnqt6jsIIF4zLI
`protect END_PROTECTED
