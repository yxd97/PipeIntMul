`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cn90CwRusvi3k96wKoI72pQjHHm7rXiBbfKRvp5vRjX8SI48RpWJ9dQ5sBAN7Lga
vnFswBA84ElEqRUKomhisNK0+Rfz2FTbrD5vCBxbj3zVUBUAL1Rq/9KRtHhSxxOg
LJljUkVcV0izZJAU3kXVtoCklDiEfK5nQSac4I85Sr9b3I9Au/ZRK5Jw/NE11R8i
9gp98+MZypq+Li5KvkOFbDQAwLDkSuMnq6bQ5zGUYq+MIX3b+7stZ8sjDE1QyqNs
hfVLiDdghtobNBjKFUDxuG2GdCk9xuMiyfMrmOVpoKUH79VlWXAc9Gu6ekCu10JU
3kJYWjQVd9GD8P1+gfp7C6nUgZZgV115nXHV+OU5z4kO7EodFwFpXvdtlktCzkJj
GOmH4Lu2IPqREEyFsGiuHbrblGLF3T+vOVDuPh5RnwyO9pqa7Bjfl6l+DcHDaAlD
WbFlzPEuA3Je9lAxyOscoF2EuNvqyVJdpALMhmUFxpE=
`protect END_PROTECTED
