`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v0kDCf1h28tp8p/6q/w0goWQnPai23gEOI/FxLPbJ3nCxlkhj7fMWqerixx+1i28
LAWdX6XIyegW3A41cOKog/FJIQWidn2DXw2j2KHGMrZh8PKQokYTtmTjQ82Bcvnx
yq88Xavf0wWLP1Ho0xbvsFAK6Rks7Jg4bhlOsG6S7XLpncHOo9BgN+RtuJnZZKN5
ITnALePtYTBa9fKPwxyh6GZB3XDLWZ5iFhhf0u1djCCu7nGfxu1fiYqP2GS8gkiu
MeZrqkU2EpStpWhXAhKAWhBrmGFENDKgdU1x15hoMXh9stETsinV6p7l5sJw9O1H
weLe9XDbf9G1VQcjO3F1wzfBbkhrrH0k4a0Y2lKBbLa9g0R/KD4U/kPynEjDixvk
nYyLjsTuK6BYTS61Bbq0ZGTBOm6xndoIZGrTBAivqrDdNXvJFaToQs6xvuQdsaXg
Cr9WgTBKJ7GYDp+RBXBEsvTva5orvSAoaRMABxeAYMAcXqYRdR6aEgxRvko5+Dnr
E3euG37OcEbzC90QNEmBgYX4/JmViCVtPlixWEjpOTBzzFbrYbAc3fh5HUfJRG16
`protect END_PROTECTED
