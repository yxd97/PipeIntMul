`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahUHcKwDqCNbl/8l1izcdpYw1x6JfIukc4vVFhN7Gl4Sn+UZUZpSAylTRIfsvNox
L5dkZBKTAF9J5aVHqs7apAGqYgfEsFz8KbZsjMS7PUA7Bt2Q44ZRNU/0gGJnAymZ
h3dFHYm360s7ppbmFBA+ZYgnxa0mhRTQkP4WzC+VYdsNe5QPrDshh/Onj9GOBcWC
WyljjKMOrtQT1MIIaakg/q5vxc4R/4S/ofhXTBusMduqQClgRt5aVxdjIraX4DoX
yWz6D8m6OA4G3TOFihge7+osWZfQKizvUWnuW/jgWshCU01iOIne8PdZrGepQ5gu
FsFm90Mel9F08GikUA+Qi16Lq9FsXqWkwHNT6Az8Ewqc/03ooKodtUnv2pqyIaLz
dBQn9jiLZZN3wMBJt4hTaeL+AG8M3efgs5Zcn/chWCXTdTLpHZcAfKxH/lZubXn8
SyIAmBcmApHC9NJq1W/G7q9f56jsmtRmeFK/LQ6eyXDNdMwLzaaxj4f7eese0sPN
YbR6dA4hHaLean9J6xEjGrXIIAdHxphSN1gii8SMN91+h6f9J32cZ1ByGmg/v81i
PKryuGyyKg1ttVN/pJX7NsU6XphQtd36wjaM1ii/5VFsmMUwtjq1WJEu4u1m23nf
CiTalEYt1pJ3zwiX/AIHjSxn0sMUGs+W8Jq71zvcFqlSrQ37GGbSPIlOstkV0/eR
TVH34khQLI1mFAcgIsZ3PRQWRx/V93oC6wUPK9qsXwKRivNHgSYFM5MZ33FvA6GI
vCe+So6PqgNMhjjiGHCB6fb+muuHG4DVnF0iy4FB2WLMEtJ92sq0cBB1UvPxBZKA
Gqa07yW8DuOT7HxblN5UPnlos9wcv7gpfmCs3HFBr+LrnC8zfdTC84z2yNZgG1IV
YXDeipaz8BvIWPng3Es0rmIWx0RXMImun+QXiNbOnIZ3ZxQh52lXB4wrcw10K1OV
2qzWi4J75a0pC8/J2vK4Hh7dn2KNDTxPm2CsUw6DA9s7R/PNcs6IC0tACxrWaoF7
Jo6cgtWyhHxJUJdUxoqDWBIJnbGmpKR+P65G0P1o9w/Q4ghfzNLSs4cU+/isnAEH
LkffBLfjFVZQEzM5FdFsfe3POF3Q+NA53iOJqtTwhTerrx5MehxcuRlh4WAUIGjo
lhKWcas1oH7sefSi5LGXdlRMUAyCuDHq8hbDODBpU67Zv/dAV7PpBXT9aEQpRsAm
FEURiKw0Y4KDL2KYOScHD81RDCKM6T7yUXi8z7Ux2Uoaxh8QFA0qTl4jDa/Q7zGR
GcAk/YX0ILdBSEYKYVyDmKp8wWS2u8tPfAwENMKwvldw4bQbmIMOadVcYvL70a0Q
1zwN0yxc9QLKq2jYAQkgFEXOfCRXRxFN41T5zyEHn40c+MS7vOjDPCCpBQ0NJCkE
DquUBsq8Irw/gZAfaF3oAcU2VJRlcbEdwoe7HQe/BRdhbgJIe5xCdL7T4R6ycxvC
9qZoaUmGEqkupGVT5XkNieCVU8mHdfd3ZQkq4pjmBrW9zPn8cpUqEYKwdPwYHRYg
LOuQwYifZc+9P0yGuUsUIimYEvIq3zAUq4oKSJvOdMForTkIFzDCKQUEdlq8z9tW
Bq9Nv7ygbpup9p0Dg7SYehEj5zv7OQ1GiG3iqKGLSxm1zWU62xs8g7w11KJysV8l
NCsXJIu9yTpbKOozVHxR7sfrAjVO0T8Ob22YlPE6CdIycwK6x4Rja5rKS3KWO8EG
UgwoXc78Qh/8d4yMNx4NLhZZF2ycDwP76cuVzuNugANX6ZquBXUKP+TN3lbh7Egj
7YUy54Ey1NZ4Yu0vWTmeTPkYzCxt5HyFm3J7lZuONuRd52cyHAJdPf34zudLjj+S
ZXPvKZW5I1QW+18xDE5Hp6A69M8liF3rdwh1j1/cBTO3dgQmMkpL6hrke27tfsAT
PfzRAqWi5J2Mvi+YxnIyNiL2loNaEyWQEtcZ15RQCC2tS5xcLkDF/IHaELzQcus0
wJfmVw1nuUQMBzUlOujrAxnPVRx1bMQjwKqAU1uCFjNP5JNciPh7CUPANnCsYsv8
3OItgGMvxnEsKHudgmU/HrnpDeXXLJmWJaBxUEw8eo4SJFQBvWZqvcHf3FgYkgr2
vheiOX2zmptjfloOvWrD9c9vyoXTUDI/gi1aDzOVFKYVlxq1bdCPwlB/fyiTvAyJ
Ssm9vRXq8QIroD7Ywlo/8qmT1ft5ugW6i41lZ7eiuEiH4N7BxQM6txi0wcT9YKhr
QPLHfFp7rWeUZv6I6QEzJ1+bffOgEWijUSkOFYb0XgISoCYz2Wlb5Em3r0g2An7O
fdr3FxN75wyIbbJV3W5FffJsZalx9y0JmpAEyyrSEqCrHxlmT6qSp2dY4UUZbdM7
hwwkMUNPpJqkyB7DmAvEaqLHECi3+uPAmqclfczmu4wSg6t8r5tYXfnn2VyFOjqb
iOxgZ/kx6nHc6ImJ2c6h5IGLzzA5zT/dI4IpgcldJgNwmut73QFEIoHTTEfT1v/b
v0CHWHT/o9S5VgrE8hKf3VyR958c7fX579WVgHkUTKgQB+iR1nun5TOJY4LEjsN1
euetE+ZW9pBKWCqvYFRof+GI/GAq+I2LoiDoXQa8ldcy4Upfdb1fp2STvNvqTSqF
ktG8dn+JDIJ/QnqBru80DXZ071r+SRTsfa6WC1a4HW2leYs9vOVOmMegPMyWOsHI
gSItCfI7XikyeTKuhrb1FcQs28v/gE6iPlBo6pyfVSP07KCtDGCBSe16LsD/lflZ
EaWpcdYFegjfMrX4vfgssYWNlltyiAsC70NL9dckoepysfCiy2YaoIwGgCFQ60Kv
Nc9vNtOmVO/kvB38QCS8doTF5mLqIsX0RtiT7cXiwkv5VX94iDTG8RSV2FHZdjvS
TL08y/UklRSSHUsln+Gjf4aTrCAP/E3sr/1JSWMKTm/P2djYBmQBJ4HOGuHIPyvz
kekCAFI8r7TRp2Kj+3vK3thu5XG/y+Ilx8LC5KZLsNzmYDn19iPO5wlKD+33mSv7
KJwOsmtbCN6iVMB0K/zDLScUVVTnMrOrJsgJizvGlBf3rmVR8lKpytbqVLdGLPmj
IHhIQpugm2yahySIzL2JnQy2jqGIgYiLzoZ67eeeovCdncc5GY3g5R+XuxrzLa3M
CF9xlk3D0jcuEBY+n5jEfjmZtt2zfaqXEFJMPXQSqrnG4tWlyYFVkEiGEmIAK+FI
U6liuAFLUHsjP/d5cmJdMB+tvQOktIEJAVsBfobfPd5Lfzd7NjPCFtiMBBXkI/Cm
RZkm0r+5EQEymP6+hP4qKhgJiiL5Bjpgg/6pBXi+IirlWUSo3XFKSJPbhPhF9vuQ
rFVZFFBtJUIkvti6Jo20WcvfuQ76TqR3gW/2knTZfWXqdOV9JTLxOu5aJ2N3hUo1
8chQqARfYihRBnJxcMvBlw8ockRrEnT2NL5RG0AAYjuXbBLL6yUpqqEVaSE5oKz6
/UqhZew1NMeJ3GTJgPoxCsjvc/8HQZLYq5JtvYS5ucvnU+AkIeKd9GTh0ZiQeMB8
/v8/tPM5bKy+4tIKwiFh6dZtzbkqu8D36D3fUr/jmsh40awogv4px9PvxvnmHjNq
`protect END_PROTECTED
