`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5xE/yyDVCIQ3Gk/mPuhKx5He8rDs64DmFPc8/95hc1uFA1WOYgfmnKTl3PVbIfIL
ZxhibAu2lyzlupeQlf4VbtxDHzBDnM2RY5v6QiRYcSgDrbV9Ofl/Oerqi1zqGs+i
bnzkEcruEzvijMKmOzsXgGHGwodzjSLtuztGinLW01g+erIMsn6IkODU9gVedBzv
iqkVSMlwwuHLo/DUkoYGPzoDjqSEZvA/DPBT6Vgr7bap+NPaI5FbTvLq7CerA5Si
9SyX4OcH9hiHHXyhWZpfaw==
`protect END_PROTECTED
