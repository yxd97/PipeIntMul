`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rF/UeCxBVjMw+qwAwCMNedjwikktqSVhy2bRJOAyCT0mequ4PS239laSwjwzWVin
70bgvJ4+ucOwgOjr6sboDWRjakZS75gghcndLBm/1KtOAfyJwC0fohO4ivz20J8e
kRdmvS1gR6QYCSqhSxQJxVy7OW4+nsPplOaw1aSXg9FRv4FYzl0sczhyw6n7b8az
ni+GtUrGJAB5C47wWVJxphlN2MWphFp8Ys47ZPlAueLWdHBdROnjFDZiKYVt/JWv
2piolvyCEinxSa9cpoIko62vq9pYoIi+zRdf2EBi+4tlqF0ok6e6CzhPsll2Ir/8
J3YH9GCDgMCAX3M7XJ7C4j2tPU2MQQB/MTBg4FD/kKG2wwkNE/5T+tZGJH+ENNTp
HzzNZr4FIGlznjfqH/R2Akxdpx5mZYp0Le8EAIS1IwU=
`protect END_PROTECTED
