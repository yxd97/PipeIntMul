`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1l4Q5uZFcqNuXoLdSMIW7dYldUKDKt5DvhgAqvIZOofCLuxGccWsQlrElRQFRg7X
mb06L5QXTF5WEUvQ1Z8JJKqeoJTg3U+opVNVka7WrDoSYUAiJsUZlLPCREquzo9y
VN3m1yui6fImhnKO79EEJp5zDjcLBODn9GKDWcyz33Pvw/e4dakA+0B7mzAH1Ljc
+cZTp4vzCvgbveIahV3rQJsxKlZBMWC5//xXS8p72epjsGo4yDAB4mYTVyMdHhUI
2hguKhMJOIitbWhZy4Dp3BwLKZETTo+8mO7jsegBgKVRh48OGkRbjJtrpvh4sybY
F6SJ4nwa3++ejxi4lHmHX+lzNoNgYt3or06PBVr9VJw81Sd36nrk3mMrTKwvfCs4
AGTlFml8MhuLpN+3BE4NFNzbOOFyqm3VcLuz2ABzSnFqibxD7kri+11YrMC6lERq
`protect END_PROTECTED
