`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iae8xG+IBl/chBUpvueDCbUVQxIL3lZbfsmfawJbGw9DUQy2Ktot44K0edavwOv4
cXCFWrwvznETXsKmclMOoz1yetNhVcQlnx2Mcc1QyMaHihQygMHOCVXUCQG7bKkM
+auQQqZUylslM1M2xjTzLClIh+/Om7lOmEwcc/CZaDYK955ykXYloAHlMSTr21Qx
V8iEuQ95x0fNTWhDzh4mnJwwfNVgxwA5pxrVCO1f5FjvQktT6mHwr14/yzJ4vV2M
lVWsNRWG88z6OOHG+EKLYwjTQccjJckZvMP5ssWxvpgZ3fT7/nZRIhFHvBbCjSXg
RtSriQ+XveHDywF/gYZ8FRucGBXeuV/VACsLWe2jXqCUj6DmK0W8uXAxq//45JJz
seFvraD4244tB6cocyM+Uodnx6CnshQfdSZXkBwrkZ1uylpGTD4faZoBAoXYic+4
ocuLQSS3gAjB1XMqnE/XUI2K+B/Z6xsN+w8GC58mTgz8qb5zV9MEO2FIcOqAXVCd
A5y3/dRKd5rolt+L1LG6EaD6hjZvQqp0wmHiyfto5myJF2fK8YgZQIb5mKNim2eH
Lj1eNsRuEeEx3Y7po7NGHfbKjiwN+K2RaFwaZ4x3ErR/JT/nq5Ss+zRU32nhJflz
6bCFY1NtX+pHcAsHTawG+4oE7TcPRh5PTXEAkddYO8k8W0NKSJ53+pNcCAsqVFUC
QzcaTf/YaV5V6dBm6+6LPsWVgLd0JZO0b8hvqfcEuTlP7EPiwfygVUpmXl9CQhiF
w23W6KPOB5kf7n12uC7qPh302W0L6gE3+Z9+KzlgNSVLJYGNxdbjJOWpAZl2tnf4
fK+PBhcNf3JCUqNVRqE/S8YdomDVZIMTX7ZcN/9jJX6cCcvuTGz742kWSLtNX5B2
SlFBCUG6NiQWtFAzt9FggAm5txDW5VhcCWl60HhfsZ/v5aXpM13znt07v+XYWmA6
gA4JAUE6qPDP8e9Ttmb0WuUEqicyd0y+ENSY/r6iiawpI+waoBgTxRqQnT5cATyR
`protect END_PROTECTED
