`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8+FkM+uEDct/MKDQA55vovcM+HdNkeNaYyhWMn5NlAJobcMprYJYot7hxARqAhMZ
7UcVvhM65+LyeNQyZVk0uLzmuDPSjuy1jS/a+8w7OUseeEVDMTkAfMw4XUecMM0j
+g1M8rfpFssJcbplJfd5mA5QBirG+c772BFpGsKulMDYOz40HLn6qqfKj9zy2Anp
wUn5XozSVJvSkM8PvMm40Y8CHAnoV57nCjf+rlc+8bC1D0TAg9mGEHi8p5bnkMKV
GW4ucZRXHSzHJD8fvvczthSEugBUBiPFjmakNmC94KlVdmmtXjEuxOAUC0jlcHZx
/dtZtV6umcTKoGKqXC2Silb4oiH0HlbXDKgEYCXC+t42NVVpGWixQLK5UusmSo3T
nBlxToynQVzfn1wr6+XHrg==
`protect END_PROTECTED
