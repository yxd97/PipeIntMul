`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOrqeWMr88xbDI1zergzpJQOeFspuak3rLOTrZB194jfxz+MSCdUuGrCbpqyj8Mh
AtT8HVcnZF5+07wLSANFQVGrkkwfcrkAG7DWjP0XgcvOpjzE02i6wSKsMby9pMQA
vuTi1hrjX+Z5G07i6WxjAn6xxG6JO3vWoXI7Lt8+C1IqHmCo08hEbbk0121DyLez
wU9dKtLnsmt4cj+X4SEUm2ydcHihunj3XzWRtVVUM39gIfPIVBSbnpD++sk1aYgB
Ellbg0T+jroS0KRJgifhP6RcnxmzqIDj5H0k8pmvHGs=
`protect END_PROTECTED
