`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mk7DIFHlXDszXLeqjszj7q2nRnQora/1NGiFM8zZT8uPTeijslCl19PJtvwKa3uj
nh+iuc6lMW7ZZwp8jLDNi5b1TQiAmM2tZo9FzrD4V9yOPWeBrMtbPX5Qda/63WKy
h/Tt5Yd8r5hy0/SKLNiqn+jajjOqzee8K5S0AYeWd5gRkkp/TtedzHGMVh7C8/at
YkGjlffMZmxF/wSMzsW+XNZjOM86sRGb05tLb2hkYNqWZuQJStKNwjEld6PDuME3
GTQZD/vwC+rXWPulIAFTlsXtOFHhDHNbNPVrO/KW+IEZyq0gqv1zNlZ7wo54Lw94
WFlbSWQGMibcHVLT18+C89bvBUvx+FopuJE8NkZUGFQyOgZHjU3pQ5uTP2IULqyU
Ltja7uarr1Qy4Zbs0TDUWp0/ef3U0OPKt/tHclMstqt3ijUtW6n0UVSygvGRGxrY
luqlPnVTUTdsdal+vm/jgbthdlY/yE7s+XteqmicUPo+f6Mh2w04zXkDjeQba18k
gu8Tsth+wABQHU1Y+B3RXMVlZzdC37l9d15QhlO+Uyo/TsvEgouuz+g0bScQwHas
0EOyal81SUFrU6iEW0oFu0ovtViksSmp6wljTTKwShA=
`protect END_PROTECTED
