`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8w9ZE1H50BKlVh64tofSCCE1fGw1pZm0pJ4FGoeO9llHPTqovPGRzn04u8y4GEa6
Kh4p7DOPUDAdMoYlj1ExxtqbFHzK+LxArGtYPHbI4IYv/AEx6sAmM6IOnKOD8Amu
5MXBdoLDE2I/4pDCobvHDn7SLhe1Hn7/PU/YC4E+hcDBg3x9qK+e4aYTOz84J8js
/mqFPIwBPuEL0e143P6b8nOqUDYXSYyJLZrTdyxWDKI6UapkaRSppqDCMT09PydB
ilBAsRg6B+/LBngcw5gtrHs2RK/GgaFdf7O8k2NqgRrrQhBDAsirYjkabFOlFtX3
60cCumd2aWofL8qEwvPZX++0VqVX2PaYYjrG4sIKKCudrASLv0wFse87Kx7hF8Ru
Wq5Z2DmYbVxCnxY9zsy1pg+YawXkASbYXNE1B6EG6/LhyV02KIxH3c+h/ZnaptoS
NGMglesWWoZyb3J1nkjzjCFqS+jgc/0lWc+LfNjTZzcUJmFUxbGK6OQDcXtILvGt
O8MdlKCqUSY0kUN2R6YWOTWtnM2cZ1yzORp57Y1H7Yx5vDpYCV9sb7CdeIkE8gDC
n0aJmI1C1U9n49XYbe03GevH2tmHKiZ4ORJtYGNJRhkm5QOaRsLIre2OYUxOgH5a
9vHf+TjfMhR2aNwl2RlbebbaXe8BwsQQG6ntvWq6URjcj59GdpLqPqPGHd2oOcpO
RwXyepSg9jLw8NsGPVVtrjYEL0TsD0AmmcLDkd7a6H1N+TI6HpxL+bumrpgRo7vE
Pa8rl5MxqGBTsSaV8mJEpUVb32joUoBELhtwDsGgNJpfLyj8dCy+M1W4sJLSebHA
qmu88/YLk6xCWCvPbB5Uwsu3GIo8J6KOMcVoPIsEjX/7uoGXwIIVCbz8+D0y8uNZ
EWMWrn34l9KJP5k751VcBJV0xNHJ9Vc5aRuDFpHLkqhRkGEZehs0lsgnfyZaGMfu
GHnTj8XoumaChyVvnKbS/6C4jaLPm/hrDCSSMEkfyiUitzFiXQuYjZ/cf1vLOGum
w+cOyvsAa8D7FST5NuoI/fAweBPnRDfMerqenpllruRCtp50eqBJnYKFvu76ypyp
6Q231a0U2OXqBLh2gP+I138xBWeuH2I/Un9cTclLfEE4pRLm5N9tyjauuEYDP+yw
+a2rj2TDxtghiyapAISK4au2Cbt5R/KLNh7j68ZBxU7X59ZgqGKimTef5AZLiufI
RPiNN0ocYt0cdy3vQjrVq0P+ve51IzN5Hrsi5e+KX6DWWzR/IEb8X/PkKvaf9yrY
++pmGpcPWOGs2W2PlQRy2xNHSd111R2L6RzsALg/phvMyh9m9LZHpaJwxZyoGiAA
DmxVcxl41bE5+sz1PJT+fR0I3tljwAGvwIF0eLeMZ1zB5DEpgJN0Pxaj2so758s7
DEZm4uL9BPxQ8/L7AMK1mfXbXaHRvvizdWhlRwv14xZNog/FcthkTXoVcIydrCti
cW8AHiMQ/xb0tgafiUlipfFz03W1s5jaxqpCNCV6vLvQatNUmm3ETzu/+HFVlmUn
RjIyvIpWADKNa/0p69SP3AuZDlN9pv/c30RQxgH7yih+uePVNWP5cY6m1iTvFqlP
YYlwDCX2bH5Pfy+w0Wg+9Bx4Z/Q+1JnxMiVZ9s6ezV4RCKhfDZGn6Aw8J+SkLRsh
RUhwqRrk1rDdvmjim74CxX1fQIBO0Th9/uBEqCikykDCNj12UQi9GrAk05t3bfOK
WnTT2HeHkvNCTxvzGXcR/LhOw1/eIYDRJajPfeCmQ9jeApOm5iIc9RRHGjuIRCh2
bjMvUmolhNQ+73TXsKBHgpXi7FPikesuwwyojRPXziyo7RSurMkADvoaJved55+v
dnHLftWALWGD/6gOL0J0RBvUoqa8VqChCUaZ4Oi+1HGX9ownZBdNFzo4xECaNGGk
zgSB1uMKe0eIHl6cNgSlJacaa2x9hXDvHQZ6otdP46Lw/ZDeqdM/IUlmavD1a7GM
JUp74TTYM9PSuclTF9i1yJBKwiEGEwOSROG7RxzGIGVGATJQiGlfCKbcic6Z2vIp
X9aC+l6ZiQFo9fvhE4rJoGM1xE6zQjN1AAUFssbun7wfms9//0pgNzdH0G4ZXbPS
2Fznn+oW7l1Li83w6ItLu+p4UCa/cVdvxR8+3wzup8KcdeVPvBDkgJ1uGElc1DGj
G6lZVxjSs67H57U/k+FJ7FSCTZcY+QRD1RZU+7GGuDJnDwMesdFsoysd6gcqoizi
iYfZL+Oa47yTF9xNdFKrtHHZ745LSYE1HJtxE8KblHRmj4e5ED2XljOAiwci1dvy
Oq1eNHfijH0IDRPAsU2uONjazcXeAONYyTs3HhfpsUQWAVBS2QkUmEHLk6BZfnHR
pmJzD7RBUvR5meISS4/gezUZj5sMFLDHtLKzvujv46FX4+HZeA1rWbSUnp+KuAPZ
dVn2EKqTCJi7vGfxn0RuZtE5iL1V3LNa0mTVaLNTnSicvoLsCWNUJiRrREDXPeAY
18XbXZY/j9xBjEYk24XGEJZJIu9AvBqgm4ur8ijROQzSlVToMLAyHFr3Bg8bQ50O
wpPr6pirrdHRK5z7xqKt4SQDNndyMBcMR9gCHFxDWBIWlZ9Vip1eI8SEwQ//wbGy
oH7zLhljRwsyWtCR7wxjeYrXu2LF3hztTQc/eKaYD4fOV9GKo8ZgeEURFTL1f4tN
3pwvNiE4rG/XDkoX4+PxXU3mNi7aqMLKGraePM3fuPXc1Yw9hqiBaoaoDo96Vo/L
IeoppG4sq/NgdMBNs7bYNQ0D9mK79GD6sXUmyfv5M7clHuNfZhcrrd9dAMbcpiVN
egiCaWjiS8UJOeguQzkZoQvlpQxgkHsSgMh3MKm6AMiQ8xLPgtxzpQ6eIEc1xKdz
YFo37R65dCs8dsZs5s2GGDRqnM5oxaJh025DyZjOyB/lMaT5+CkzgYFOu5PSCS2O
0b3rh8LWlbz2lhF3NVP3qVxcM2rJ2igG1Z5YifvFE6f/0UQn8tetUlBVWSZCLX0S
gUBa5+9jgRi1s+CKq7u1RJVKtJ7Pmi09lCDUkKh+lMZUvPhHosuPX+e17r3120dw
3TLIpy1lcOIO9Sal4bq0ZhnCLae5v/5WeGc5GkZj6gu4ttPqckiQlmPBJ30NiLk/
lbbKD4CdamaZuuywyae6ihlo88WZL1NG7J3xvVP0NosXy/Yna058g2q4Wyi1x3Sj
IdyHHOUJlI4H0B8JFmpyP7oek0r5ThYvRKFnZXqKtTIW4x4uZybbRlgDfPnYh2Y6
kgGjot8OeLPY+Rr5gSwnvgaRdwbiqQwSqVdZefzrAuDnJ43LivDODRt9Ubfp0452
Ax01T7T6oK63B9/SjKAV/KEynpVK6ULrVqzx+BMq2cgM0aemeSuaa3ITmzB3GLOB
btcomGGr/4udLFNnY4CA8WA0XCKeQOYuI7jWKg1g7V+LuoLMvbcM3tifgfb98gtA
UBfTmrrs+lz4QwUduy4Q0YT55cMnhcQxBUTLnDAnnUjICp7LBKJqEcS3IwFyFoaX
GjjPqApkBUOxnBEUmnZ+39CzpnGIvjBzi8CePBtvx3fYK2LtiMUFOYSWbNRdf+mZ
jPfftSihos58pdgfyamiBG7EdDuPURLXBFDXP4eNGfujfhJIFD4/lDKUl40mK2AQ
uqG8Yn/hBMbYi98QLDd0Pn7vz1bkatRW1vK7r4Rm6E+DJLJKtJOO9yGnUOod82tC
qWMBj3w+T672ryCz3oPYDmVO9kwNUUFh80wBTz8dJQ2jN069Lg1cipeGuFi7bK+D
FKVL3wtnyq6nyAH9vWPCdxuIo8fS7a0hMt3UUJ2k0uwMEyWk8OtqIA+KFGX+ufSl
XmrPIhU9dD2m3TfmUcevApUBoSkqfc9eRFFh6bjPsDIPdQ2HaBy1VgnHXukUlaoe
YSq82sFT5PO2n0X9hCfzhmFmNzZ/EbqXUlqjme+HQSQGMztYdKURVprFxNN4hLK/
Zz0GHhYvl7H2cYOWNyYwou8fKnXGzce4ntAlQQp3ujsFeyKcVNz534R/5vVEEAIc
1o3+S9E7TNYangFiX4JugqF1FzWjS8ex0GMP8FY5drlrcuwX4Ph5/jKsMYrVevhR
CGSpyrk9+RlmJeL78jH+cN1XHplIM8VrE3Oar4pUgATQNdFzgil797q75MvhS9py
/bn0h2DK+SFHFU0NIn1GjMoTWd5REk64lypfyg6LINn2ckM44wo0jKRBop/FnI1i
YZRsaSjwDhJ+vzCXrVoni3jHrwqlN6mLnbaO2lXEJCAIAvCEanqqw16O7ummmvG9
EgQoqcTTKf0uh0hAsJY4eqSgLRgWsVVpZZGTvKLwbKWcqiIyWa5xOduRyKTYvui1
EPI3zndu6brpoqr2T7DjAsKrljx9hEDOQ4VOkQNFSPkckeXKI7MLu9Lr4VyV2H3J
PDbyxrEvIUCgCTTEvf16kivLxGirTJuIRVBv0u/dtfBEFxBfAXzW/nY8btFdVngQ
CsRlX5hDpTvBMLIppCtoQJLwcWNjSMpOAZmEjuPfWrxTwzDBqSZNWqGS481MLyed
cGPs8sQV5GyyEY6vsg6FGI0zkKSFZKbDGNkWbJSPqYbxRLCoaSs7qE/W4aVnvqIV
mCawXpHiGOTYv4633uOSBK5HP5MDNaWmNucCNF0bmoVRc+ADwEvWghpJguUTsgoD
WW1HFiWKepsMaALLcTPZOjnd6rlZOwdVQNzlwOTyQBlzIe8bHsg5tbc8Bv0Vlpva
xQFkYXDz1SnmwS5Gt4ZWZUI7cTecQwp+C876T6a/hGNC5oHOaCGllbrTXUxAChC4
Ky5xh+UgwoTmxln5Bc64zuso0NVoR3Hf+3hVR4x8YzWbPahNOP4p0sM+rTMeIEtM
FFHmeS5umvs/pvjpaqH4MnmVoRk5CPvKOXZVgKmVDRhQhrixYS0UifOUdKLeX10+
qXpd/nbmhFabmJo91FzZOzxeGcODmv+GbhwGgxGD/lmCMNHkzqjxPHN+bOC4ft5e
1x/M5TuOfI4W9+mGWHfuFJuS0H0mCz41oP923yO7ShWOJmiaTV/DsGsH/HkT1xD6
ny06dhRVQiiECQpkpFw6ZH/tPOZW5/VUqHeggwYPu6C4SzXaH0mz7UN8CJTZ5KGH
Jih5aXIaGBcpY3GqvKSUEzFfHtJVS2rk5aAOgUlQ8dVb4+KGFnQjBW/9+t6OoaYx
jCLdKImzll/QzlS59Jc4AiP+lDl+WjqFdhUY2bCsH1U53Kfx/XqU7BVKFhq+S6/k
4a6HHE+0ue4MobchaEnRSxfE2W/+cxCx31d2zAPwT01kX88e/qlGoiTJuS+TOFmK
rlNDDiN/q6B5fB30GaC1Y7d3rUzgFnhMEEInOk4aZwaG3hxhWDBsTchRSdh4Xk3t
qfv5LjfJSwadkpH/ejponk7W1EKugdpcQmP3h1P513PnOPrGq1+AnrWLpFXEP4Ct
Lujwp4pHNvStVCCwtVmqR7oriLjyQcUSAYjU2vPeBeo5n3sBDoSgLmIYKbG6cQ4e
cgP5bV8nwA6P5IysLXohfxPH7h0wFqRa0LmKPZMI/Dzd8QNttocK2iq+UJ+4+5+b
fI+Q5l1WDsKYHLI9mRAtl3GjdaiWhfIYoMaGOyPXM7Vws2tTPMediXIplIn7z46G
p8o5X3sylVg9KmobjQqHZfdq8wIxb/yXjxgmRVn4v4L7pNVZayBOmi3rSX32k4gY
80//GSGaflptBFEBSjLlLg4DrrJqnqdJK6wn09Bpxj5QPSWYSFtJ361WoVbkkoJE
1oVQWzfkVVpokaXDFvpV/aC+gZzKZKAotaQ0Pm/h/Wo9yVg1T6Nzxi2fLNlTimI0
/7nZkSAcHiXVwqfk5eB+UlvQKo6As1ocdDbMocu0xEwv12/uxiDQzYIbQQO/myyH
JjJkJeoSiJ/UZgSQHNZV7HFiEhhvR/sBgDyFzTL2v6TmFFVMuAbY6mDb13DQpYpw
815wWzePz+mP8bZ9n/DjXTKYcuIRyA3cZ2MpnNhSByFyuA45W51nmq9CFfDJ3W3I
PQhlsWjrgGx8sG3++gnzJfqiE+YrmoSYZQj2s3ErIZC41wwAK+iCYRuaryfUSpJR
zEz0RMBoQ3VYzfRxfU0Y8ntXYWpROIrP8QkfCBzKGx2MJYjZ5P/PTmBfWlzaxjFd
mW5DU61kA/7uzxvg0fa9xJeM80h4ss7Do8Zr1a/L7J0Nj19ZWWJKqz4JbQMpZUXu
7QgXHqeKwLNP+7J/W6kAzLrkjUn5Z1Ba0b0qOu35F7OzEv8zDeZyxbJ3pD/WLuWL
mDlJYRmbkBJcFEpQ1PgFEs/HunrQAGxnkvx17FOzJi/zv9bMPebZZBcUHo5Aj/Xs
bdic5UjVkdXN4ibQMq3/JQ5fLdWqyFbb5Qzop3FV/0+b3jE8ltJrVKZyeHl9Myzl
pOvoFE5gvslpO2vBLG41h8Xchxuk8vlkkcCkSrV9LAcgsFsM8HrzpiftshPDQnhA
l0wdIzdD28AwPmfqL8Zh6idJ2I6WQQaUSyrtnXLahtjHVekzrIgXdLcLD8lj8e+J
Obb0JIEt8lMEdnF9PYXSKjptMGGQL+hz0K7J3gn8d1bdIyLvnCcnk/WyikrFK9Ta
FIh05dbEvOtTZo+5TOA9GVDV/gK19juHK21p2bgIJDspP2lATIQKrKwo1uw89tiK
ioPbfVGgkc5xAor8U8JEBRBiGMT6ZmEMrLn827mZllgTZiMrWpWhMzdEmIsACHS/
u6CG7vuUbM0kFtm90trLXpHJRIxMQfQPDTklIPBD3GIPqvBmIeD7/kAYQD2Q9ymh
9OQqPd+SKxMCuVFrB3F6pVygYSZPGPN6Cx12Um7fLGUe49jL/TQqNuLkE4CoRdD8
VKTo28SAX0ww6G7hMMUyaBqenGgr9iGNZVjxecjBqmnualYzdTCd0B8PQzR5TQcV
zyEmATszTE3nLT9JFWkCr85DjSqNqeZlX/4sjf1+D/Gxfiu6IIK7KEb5aRBrkZ9O
S/sfGKr+T/83Lg6QYNkeCyUVO1Kw478bGtwqSK2xEWiCnXjIxC++fU3nO25bLJEM
raF56K556LYDtrVU5jnHpt/Z0uqhKI7hBkNvo4KT7sriUWDYu6zwHxndUa64CPg9
5dOu19kvZCLPoQ7H4dalfKYrHjV3ltV8iDp5cO55Av6MsShsB+qzGX665d7ropcd
eUnykJuq+WA1r4HGqrACoU3Ws7fA6FVkxen4SLJgpCVtalykaz3TS7lf+Jt2w5pm
mZMpHcLrqffYp5rMQjElQuG+hXR2cHr2uSh/7I6Psd8VLIhoH9upF4eU5wAeJEMq
JZbO3RKXFvLwsS3wvEkLY8v1C2OQtYGayvqpmIiMMFfJ0816jdsYaPIU4zjm/IDP
0CKjOGx5ryVeQhJSKVDbL9k8jyZFBmJpE999YfTCuKXWbD5DI27Yfz7A/nGbW87T
HBoCCVQeuhGBUek3iSNHN+w387fqKB+Pb605JJNZjhjR/ibcrOu+wlyWOOTSGylh
i/V//fJcs2i7rjIDrzXcXlfz9Ti/HfBTpyIE9SFed4FUtiBUx6bqWoOYQvp/6lQq
yqcmX68OuW6dSDIcDd7w6OT7OtjL7iGlEdKdkqxRTqeSfZU4xxIwL9aqTLvsRKPF
TYmxGWabpt8eViunzATwumJQwn/wRNEMxKjZBIlAm1ggN1lIgnwYpQYDXJm+qaDv
9VrTm+VzqCv0FS7iQE7YFrVwQSJQfk3knkrDOtSSzAp7PlHP7quJdeMNinorRH1U
fRkk/R0OxW/Bheq9SyOSo8B5Y4icPjGjFvVsM4E6iDVBRhgJ2mvOP/44pK3NK8D9
JKVpYmspKSDN4aHLiaoMv76QM8mgMYNmrqFTvsJ9b0fZxQTNHaDvRI1fcPgETn+s
z9msV4U4wCP9xyDu0jKQgeizO/uc+T/0qVEvwCtfUFdmCoPfLfQ8wqjUipiq5mPG
N7czIoq71AtNYUA1byqvQfgVcwxQKgAM5B1KquhHy6QXGXhXKLdRcjx+lgJ0+DSX
Y9Ax2gZbe4nnAWb09SZw0pPEvI54Uk1Og2T0wQ1wWJ3Sq9a6F/XIeKmvlNwFtlN3
u2N8LXWLryPmHlVVepC+cKRBSc7QSZIofWMp5nnLTfvRat7MLMk5vOsZneZOxUcD
qoK2t1wHAZbPwu8uZRavHt/SeTLHrryaw8QgAQvTTar1aHSoOoAVYYqapkt4XScP
9HYx4RNSrbiMEaRPvdotJC0gmkN8k1LQqqozXNU+LoHb3nCwCNWcyYx+H24Viq/b
6Q7lmj/wW2hxMC+FDY+5dW5ai8F7w049trsu34x4tdXCg+xYUYI9PDPDOoNi7ZVo
ueQH2ixsEPwS/eJRoVQ/hIIQLxKYu8xRzkAtAAu20WzvxC5yGz49JGDB+04pIQn8
xQHkXitTZHHHnjx8bP0S0UO4nqhUNNIsArntHOYLJYJr5KEennFnCchE/980L8oN
34mPrPnQb+k0ijBj/OHr1rk7vOKvq1pmra0as5pAUwHV3xgIu848TVqSOB4D0uUJ
GyGxdtQ1WGtgT6sXWAtglss7CMPiSpC+/LzU2Ij8oLn2hfPYmND9lPBZWGjw2EcP
pcU2MY2RBqxgLXT/NJdjeEqNt9xd2VqhxRNDloFnf/lN6gGUrAJM7Hc0BTp9LaJO
dgRtFz75ejO7nvAyjh8whmEuGbDkMqIfuzlEqDyuddDAApFKD18/vtxehXlZ9Hr9
X5sLt3qZKS0HDiE2G4PrQz4Lq1OjfB+yuzTFa1R/BZ65O/hCAi1EqStu0bbRnF0Z
T5dIw0NWedW7gYGO49kh5KSJDwBn46ml9wBsh3OB2NZWC9r1viNITcNk/QyJ2m2m
IUwPY7BMGU4b8ihJje4Qa6rKy6wizD33EJDPV/KOZ0E21oCXDS2q9HMneuCe9WiS
qj5zl/gUNNyr6TohSs35/LAj4p9iB3CcQ2zgQnxEpbBC3GdrEM+nA1E7rCmApxhC
5pWgLlW+3LZbZYdmmfyy3reSYa69sw7oBvlb7Xm+AC526YBmEgyFeAHc1cT9Va7G
ePKAsuOc3aT5y4RNC4jeLux/Cl1iKeCg4RMgBAxYulmSl94FYHUiigUUpTDy6iVY
tDRqrqIHID6imYN0+JVj8g4l71GYsnvz7NTTib7mH5CPNEEXlXH1+gKiHPwbT9C9
6SQ9iMD9kZxsmpBLvio79iWZYMxMQEYxkyTYzphJkCPS75MbBk5FUayjWzcTHbqJ
4JkdVHWBcjL006nXcXUXy8zMud2eEKaS9iNx0q9SPyZDnrRcrkPVtsO5YPdbSrHT
u/z9hvgLbsw3O+1RXCUxYIqNHET1MfIEDSbj+oTJc44oN4HL/oE4Ymr4yfbtkYlE
qPPNUlMZ4X9aRN4NH73WObSD7yysJSPou2Dg6/NLVcwVxCOqrPZfyE768kSpMEPV
P4IuQde8z9mAteifLge+r3K4luR99TDW8fdVKaA2Zp8cnonVhEsPVlFuYdJk7FY4
bkPDkPbOD3yxqymaMHF9rwyJTmyWC/vkoipuOuJiwgqLJhmDElExvHitySwiuY6C
7oLc82jt6ufgSIFayTkUY8sEwao+yNVeIfJcgKFqu8ZUsKbN86tOq0e+f/2zHbqQ
ae6sQAttWp3UzGYiSWypR/I3tP2xQZrbRc9VEnYOgN8Hj4pxtYtjj0YgsdSjy2HK
SIX35v2rFcrtuX8ACoWKxCO9lcWE4jre3D1x0gjSt6OlVSkkqQjVFWED0qNcNIQP
zECqe1l9GGiYcDft4oZbIpa/qWROvM/53ryqYxqxWg+Cmvz3slJ8df8xSWnez5fw
Q4C5ZYjaNQNK6o5sJXlc/y3RHsqPUZnEFOybBz9Gj6MPkqZBXR/VM+zgp+RpVHAv
2ncS7Np/n7eoPFMweVL0VQ5p8sj4GjaUHMzYC7I15TQsfYysfTAwjWHi20K4o+cP
safXgjCAIJUDEK9ij05QdvcegnzxtcUdQDuNbLFsu+kxhrFGnwvNXh9yofRfeew2
+s+RRAAuwkYj4uk1/txfuFm8zgAiJUJa388u0sTCvfJ0iyFMjV+D8LFunIbhp3oa
4d+PZqje6shvdX88AbAZNSQADoSevoFlZEiWRAS1dUuh9eU5+XxhKd7YyedzI/+B
2jUPARYkc+t2V6zx2EHo42f/pGu7gkOV8tdaFfOhCaUiWRCnf6Kuxxi2PTD5Ag0V
AJ3tHBpmSkv634Cuv8WWicV687fJCzY0RhbT7OpI0UiG7KpSi12Lx7A7kKDQwUOn
X/OT+6/vRBW4zK+oER9TCYXa3CeTLER5Ws2PFmseqX3u3vdB3aKlzH/EPeDWnq6S
M4nNh3b1FkKciUBK4mVdVPKkT1Bod1cvbff3PvpwJHqR+oAkQuVGRGcz/ZsD0N83
9cJjSXyV45c3DYZYHPcivGe9DidHxyWPO69PiFL+Jm9cyDgl7Blm+D8FRoRgVka2
EQ9sRLci1TG8pRF8JRvDZFEd68J+P6lPKe95X+Hczp07eVjHCVA/BW8OTxKxtRcX
JOqBRZpQSFGeFU88oKwK6gK2dI/MI9sFYvTJVLhoccGYgYRLhaVcIjehIxBcyeW2
AA1ktTRc4lWogaOTG55xS8FZBTfxRBKkL7QflDFDjVtwmRn8pVcMd9n3/rEjAuWS
3qY0GPDPfmNzFUE3GX73kwxHYV73rxskkbyqEvGE8hgc9bhLw71TUfZmWSg2+MAc
iKbhg99ukS+yA5uWKqM2SotOT3MfFYnM2vkZ8G6nKcZ6GHnpy8c9quzJzjhJrzKv
i9n+v9DFjFyj1WqZOHdC27osAhZPNLvArktJhLTw2+CRZyqogr4WrSnTuZQIW6cO
hoOLz6TWPk3h6v5Pl2YZtl4hs8bEz/XkRsCI/FJWVvsQGd4hQsdwt5pe/ti6qcOf
r1lnb9UExyyu3TNzZgBtekSG8SkkYjQvFb1kGeSRZro24l6vVZaYEek9lu9mJE8P
lDcDDZoTJMXj0vqbIw3wxRHNM1rDHALk/kpsrk1C2rxg1xdxP1zXk3VaNwgzuO7Y
8MVWYrT1YL0c90/9lZNNdBEMW8C3O08uraH1ab/adcG9lcYUcg6rFiDa5XnJQot0
RDHPeAf1lfGnYQlKW59mUhWEqm0Sp+mjd2C0M96VedD4Y5Bvi2WgTgvG07piNUY3
ujGoFZrH5uRx2tdJ5wtXXj/AvSdlHueNIb0IcZ6WjV+azupf1wX656wd2ieEHiMD
QyUlvHXFA7VdbI+Tt0OZDcJG8E8oMAQwPbJOesgUl0TozndBaxzfDvyVCrqdw5ZW
PxVuDpfsMcDih+azlJKXqJFtaaIr/7VcLnlySEuRdJw2tlJe1+oj0vybjxTaL61D
84RMrlEDf2ubNcprHn09bQRe7vcKwUyQvV0YBBJkaXKATGx+fjpworbwxgfnyEf5
MSWdCSN+vJCVvzzsD9ggofGhcL6yTMb/eHWxArRfHuqttob2Yj1CpwTtCYUS790z
NCxTdaGGaUMFV0o+uvduVym5HLL9WeIWid93ls712nRJlpqBZSnugSLcoqxsrtiE
ECEJkOV6P3KuVorjr2qivgiWd6b07m3FUxToJvXCnz0lpN93TrBWY2X/KBfP4U8e
wERKjzwSTtiz/ZFHO9VxXXjpJDf5AnodOzr+YIMB797qZtUFaaVmvDuiS8ObtbSm
bBG5PkgpeoJYseYxgxLee7mDKvqKe85fh1q2RaSRpsQRGzXw2nuY+PgefGVsYsw2
WypigOAhElVsMZ0QGqosJuCFHhsVFOPKXC3EMLog2tt/bEpJT9fmHXfECTfv3/6f
cjA0jvRzV3aiK+rFX9bltSqfRc8YwLdS1TLxpfssR1OZRhxbcAtCGpgDdUNkOXyR
5xRBMO1SB0gjEry9QqITV3gCvc/pzjEYf/47ktXwTE8YaP/NgD4qgWcz3MXGOrI/
s01dHG1Q+5MWukXGvMFZ9BRU4f93m/sxupiw/HU/dhbtkoTIQKEPkMNIWVyqOU3G
YVZkJJvskq+S50Nnq2B5gn84gcRdIS/owBs/9MPe8ocGmfKvEQYT4F//i73XFCGo
2b//Efz1JoMxWpFrB+2wkl3FwZTzBsxkvu9EEmkH0uDlhrgl3wMbHWOLCe04hEwk
a7wToDOnjU7uC5FyIWn5/o9l9L0MH1slHRTUx864sxqL5Ie2E+UZOOh7dqMxhy07
0YGid8DZO1S0lehYmZAnvh1nCyt6cejrJQGaO+jNwHF9UnKathnXubbleKkHORf/
dP7j3VYHfrgOG6muuD6hSGrwb4HIsWF+GKD6ondTXI23prd5jcpbyhHx0yShVrxf
QuN+ABNt6lRn+tcvRrjrMLIediJhEEXTfy7CFOhFv2OqDhRir+fliTT/axrzm28m
jkrnLuiZmdm2XbiBm5158oCIpY4zd3gk1deViRs2c8bDRWo1hwKv8mAgYv3WwZrd
SZSx6mW49IS5bgJ+0xIkjJkUM8tOOMN/tGk4Ta807fVemNbqIKulBV8YkCKR7+Zd
f3AyslNYHNXsl6tyudUiQZv6r9GyyuwTg5C9JBnEWMhzdDSxKoW5IW8304hcCg29
bbF5XUScj+RhUadMbmXxRjWPHCu11OSR8Hhi3kANxvMJ9ZkpgHzd5A3wQG4/UsEF
ZBR1Q2Pq1blxpi/ALHJmTEhYE22CJ5hzLkGflfQJt4q7A9+g3S0N2IcBwMoDPHUN
OwxKdiiZ77PX+/BnnUbHhcEb7CTudKQpbhlgYSUql2AnZD2Rn3DntlVVHs1jIAYp
oDDU7lehRlDOSDxXTLcCeDsBCpwC/90qOxZm09OLrreTeaOxcawtw8vkHDJxZC/+
OhG33QY/yejufxN91jJgdBzTFT0ww9RE55DXZlFZM+7LxudVBrJvuKvNkY0psGkW
F0gge/0qFQgBKYKCzouzrmSS65K8xDIQQrnKH3CGOAmaaDxSpcA6BRgsQDH+AEeR
XtWbbXFTYoaOpGM1ZGWMPG0WLvMcJ62wqJ5CGICrhXb+aTRk1pXcvUn2oA/Zg+qo
LSeVUslZ7G3WgZopO1Z0dPb3x3tS0yLD8eSb2ZyU/7qLtVxMYSjm1Vo5G71O/Nz2
YdM4h+EG6h9c6g+DMCilnU5uUhAQWb0wKC1w/2w2JIzly9/TaE/6Zp266ir6G/gd
HAXF8dOw6yH4A6akxSBPlgukmsTTl96UDGa9k//yjo0d63l3+RNIWm3yTA+o7NPr
nrx27P9T4t8t3bN40hih7ocsUx6agrW17cZZbOKkUktGe2kjK5uiA3aqMSgTPB6i
m8oO5THAq1f7V2ML5UjffDBqSClsjQVsyLvf3A/Gh9nWU4pX6Y4OCMnZUKiO0YWV
KtpzhG7f13obBeNSH25C8HyMmrBlwfpLKjNUnoFqQCmCzM4lzZNyPbqPnPRnEHuG
IKFhweWbnMQhlTi6G76+tdbkP4ZPy2LshWoSYXxjTgkRxsTZQzOU78CY0VY10Wuj
cP+7PqlveZjfOLt8JOYWDbsqkpNZFENB0TNzAuUUqRFwgG45n2lg7IfBE7cuz9oN
MSi36YzzYFezxNXMoRs3PJ+LVJ0wk4U6Fc2QYIAKiIQjoHqE6LuKt8tyJuDNFcMS
rTLnro7ZhOgN84ZRZ9aNHpSnud918ZyGUbftuq28ajZzdGtpHKoyhlPK1GskGH/0
6LYktB1omJK+0uaHTCZv0dM41IdxrKI12FTnGIB7KCHpwONGD2fk2E2FAjFnXuoN
fCqA6O8FYjA4HxurRRCHC7GO6sIPELN2CiXK4gIfqGc6ljJvxc0Ij1SOARqXtjIV
wYJ6du6WUTftg94GM6juVDH0xyHGjaw69PvDm/uUERE6nevgR8AkV71DebSnD0LH
A8IirWfNtvBA6D390ZEY0/SQRPTDHXZRFjhDnDVBGgeIclzXI84YXqDhqxe/Oyw0
mJDUkWmJrXId4dbz6ntP+86yQ5NN4LUgZlH+wVXfPbmCvJnsxKyEMwvHbRCrqE/a
5ujsBDvh8z0S+vnzGmF1H8eHbEcABe/IU+WyqW1YhAbt+bJUDL5nsCqURYSlp8MG
XtTbOatEk+Yc2Jy6P7lHXq0+bhmHvJgjUPOHMgujmPXxfcHzu0gnaa0/ZJp6Qzga
gcpBQ8FXrX+ki4ZzGmYINPRXYBVW/Y2c0zsQzInLan6utKflZZ0AOxsDDJIfTBDl
Rl70NL5xfRRCSe7Kt8xBHPl4AQLhbhyO8eVmfr+wHzb882zATeewSE/6V+FYHxSo
gvhyv+VGlkx5tZSju9pyRrNG7mMBVSvkMXVZiDWZnlOXdVdZBdpL/vsVkIKlq1rJ
eCCPzqQhHXLNY74RTU3SlN6+AsuY98H03zhSTvOvCZMGsnRDKcgZ4BKYRmzqRw4k
C5oqzrRMoYjFOLSw6SBtPQbPcnNJpQTZf70qkPIcCfrXTd3oipd5/gYvwvV3a5dk
QfAAIsvNX5N+YcOyppivgkMtcq1iAGcqj8ax6VbcBWnX2bA+6MWy9IdvfFjr6qDi
bQdxWQ3wdci62RPUwTZx8ebLX+fRLch6t8u2IW+MdpfcSw5ZGN72Y1bD/Q0aN+2F
7fN/oI7h8InXQTP5V5wfrERmN1GQtD42q9Dll0CXYD1bwKY82jTmwgjB/CG1py6d
UZjWNWMwhUIfXpnA82xzIzkVowOkDGVI4N5/mUyt6IEG3N548wlRUdjeAtvdyKgd
OxNq/dzJG68zglSo8eJWSDOWpAUDprJXAPMdvzvzmNV0uS5cZzsia8/KFPP6cyXH
2VvMV55DEkRULSluHJClW8LJDIZ8teoESMyhqM6Ggm201aiNy1Wyq5mB5Qt98I3w
6lbDCokkfINW2dq6FOTMfYy3VNLG/Kpq2UjVSsEzgsbgRC9jce3MJi5RvpkPSkwg
MYnpAz1b5/HAguSAAgx/Me/O69k3/BDHxEFDmVPf9s7rhKQvm5Bn7bLn34JX8RpA
DjUE22tY/ihMnwcc/5+Zww4kiOVAMG+6ihzb8sZ9HqdSwrSfCsP4nI7H36h8M4N4
FiAy9Zftutgs6oLiLTkDTm5DtBiMWNbZFOkoHcbMnQApCIbd+2yMm9zYFzhGIzeE
buJfcGaPNNUKsBkeUGBLJ9VV2LLbILckM/qZD3nd8R6aa6XDX1eqWrBCIQb8BvwO
OFy0DjB8b0VNwhPVSmgXfrKHJOqcJULXcgUpMvPMpQGQSFVzInm/HZGhWV22UFEP
10rrL78KrdSqDhD/+RykxT+rxE8/f8bZB4xkTTsgGGUNbJFOzsCy4jPodzIJ1y+M
7u8bdtu0ymamZwgYmcBJXPzBwaf2kvqXT7AEHWWkKAxrlP9/YrlV7luNSMikShPe
hBIOn/FM8uNRic5l5hdsyPE0KdoNw9D6WuU7623gey6GE6K+BclGC9Ew4t/L3FNr
8z9sqQM2lzEhjW+oKfGjD6b7x2RHUahXyD0KDfaU9hBysS7QWqDnRuCzTDB60BEv
HIrFVDLKDFidUjeqqzyBXGMYa972OkYhCIl+tN0NUG3Y6PwtvmuirzxzpuFReDgp
0KMuU6mGstgKjI9kHoPtDx9yp8XzC0PQgiDxq1QmH4FmF0YYksm4wjxQa+XjAOla
S1Fq5xhi+3Ecad5BPgbHvbsrAkF5x3RaHLkmsj6MKST2B6BStSpXtLcZPMsPQNmB
INC0o4aVFWUejC5WBKWB9jfepXGpQvPNjTWWDHjm3JQrhzAp1YS8Mmq7N4gckB3b
W2nnc5m/2UCJR8iEOgBn5Aa7vpBGIUVKbD3JrzxySznGVOP2nPR+S4t89qHKFKPd
cJ4OicL1P+tWcBEaGDbkA4QzXVfZVBkYlcasXOU8/NDO/fL7yzhO3i/cOM6F8TaV
UrZ8H/lx19CJstHhT2j6zgaAbUgcMRN0KG5Fun8FxilTjeACdQyqpNOrCcAW4iis
SvKQOmP0+QBskCXRUMyT0cndhhvapIQUYK2Il7z1Bn2yBDDP/sq2p2qCKC16KH9V
7Yr9Df5dsspQuRS9Uo/XqGFTvpqckXCKJeFaLVEOgSFSFAjHPZF8/2yoyp6Y/H/A
9wYdgIqBf4YBbVPEDOHYIlSnmk9ZRZ+3O4l6JzbjpuCcIe2qk+MlL99KoZqrWgBG
UzEnx2E9l9OhdgywuPL75T5T1VJu7MD2cJG3VX8apEpcngWfvHfXKVm7TbJFgaIK
74qgLBSL224sB4rpeAz1DH96K6qK1OVmvqzwo2hJjeiiHvBpfyrZQJLy8ReRBL8g
kHrqCMLNiAI8XRLfoc+iDBat2/MTZaaGJ8dyh3p7Sij/f+eafD9iZghibCA1vQdB
6GXbDFUqFfIOSLjeMzyZQUDLDlHo/pUqfjB9Xo3KBVbz0MKZM3cSUP+j9na6hvy6
pVXPejIghtOMKoWGiz7HMp9st6u7zdjFmGICFTv8cvkvVskuopr1O4pZmw0eLV7i
RRewthAPZ9pEvTiA/0IEoHVzZ/7bmBRHwyHy0hSUx14NpECBz3dr5Jh/4cHlRXrK
wplq9RVbHLX5xJuc8atIg7eQB23fh0pto0CqsVKcAg3ywXdvMTVfOMvOHh2pbqeN
RXvci+6dBX+oFLmL6iBhoYa0eZt1SesZUpocShp1EFWtQPZ9EF9d9bFL0vhODUL7
Yc7sUQPuCkD0cLp4YT5Z5+ndBjak6T/Sr8naa5rTsSJJ1J6d6NxEZoauP/SUo7/r
M9T8GUFAAnWe/Q+GyIbYQT3CGOdovFgBKjcwZnw+D8VeNEDEeXQe+18a6RT0RNtT
kZkItypcRpCbw43iFyZrxo1FKOSRiuY4AM6aWTGNF4JNCWccXFg2xpUx+KbEA8rn
qndMvP9Z/nag2ovtbB4eeSoKV3uTkbrw2XPQBlCX4CUZZ3JfYrfQ2SHBz4Fst9mF
eWKABZy/WhEh4Ya26iSDtLw1xW/VhnlN5aK6bp7VYwOE0IPf6zPkL/q3Z9ejmC2V
4FtWNYypd1g7NEGaOK8e1Rpp6hfCrGvcp5bFa8sAvj+71rv/7Lg6DuliSdO66Xf2
CUHhRPCFs2HA2KGhsJdijcROBY/0wfAe7dsY6iOtOQKqYIkP52H6ObH5w1lF0pQ4
DYj3XybXQBdveXqeiYbylLNQQ8TkseAonvS2jbOpaoL/2kK2l2FKlG9ngJ7P5xgF
VCfYx2o96/YXMs4CGq7gDovvhENiiR8J/kFibiRoR1T7hnXGRc0sbVv9Xtd6Zkhk
V4MHye+EKxnunc8+zdC4LLnqDAwZ5ILH6Lk3RrvzsUXKWQ6P7KmEPkx6cBlmPyfg
8E5lIk6YwP0AEtVPGHhexr4y0P3tq0yKSj2UT7I+5OkIHQxUJ0Ae8wVLKcFOJ1XR
0dfaTn1EMXi1PZKW8+qqdVMomZRZfMM2GenudnouavtxRUALWpoCz3yR1ekbxLdX
EiimB+SnMCVQEJf7nzHtksp2NBrirb2kgeIqrOTg80Ea8XmPJ5qI4VrEH+/3L/5n
Zw1yYjYegpKVdS7eF76MG6/0NgimKu91e9qFkVK0WGv7Qdwct/QUyrPniQTWKckL
gEhSP+lZYRpzpwwITZGDWtESQGfT+bvc8aJ2GIEhAOnJ++Z4F1zlupTUkwxyBakl
ulpoL3OwdceJQUeK4gfi5l+Ggjn35jRtPRXdbvyEFQLe6RHtIhM5963gLuxXglgI
RCSbxHh709ZxXF349CquYgRrIJzy6fW6XWrs2yktJWFua9CHyjg0g/dNHuhOzvB5
KrbIPsXq/RFAjL8ZPWrRsXcequWde6wjqQPDv8CCP+gqBR1426GpGatZQcVAdhcb
NjluasL1Msy2FMJ/nC0wEHvQW6xnxiGxJVombVUMs0XXNqt+SdL05W5qcnPYq6FN
dN/sSvzLr2qS0KgUlLvlRUAQR7tQqzb/wyFTlXs2jUL4kPIbha0QZaxw3bR3kBHU
EP7a0kRrpKgaWyWXnIwPvJRgC4yw7OEEb7H5vvErR/WvmskIyu+6wSRlpOoZnzgn
YR6VDQXNci+0U102sqAl4PQ4EBZrdJl4QPNFkL5Fhz7MdDsZLCU/aKb25DIJaRQG
jfDCu3mk10+5Uu2TrGL+LrJBBE91hClvkkhyE6Nak/suHpYbigLCXqXKmzcYhrWx
C4PkyJYwJcIt3tZOdelArWLal6seMZ13mYsLI18SYUqvLBXEdfIzj6VP2bz5+bOh
elgVbiNqApEI7wDin9KgfmqQXBM+LfOdy67TWq7nnIe+l1EV6qWCUpky7CyNNeBL
F+ff9gwzfwrdGHZrqKTxIB4ruqReEwpbAzDI/ZOzS2VEzGA/fiMwm9cbqIwwoX1q
nRD+uL0jB0enNXVG+PXurpCgZXbAfOceAFLgqKW41/FA6soBrA2uAn1d4siFw/Dm
9z5CroqtZ9zK4WUoRtmGizJVkZaMdtdfz0ykKE1p7DwGE9XC/Xy5+X8Z2vRDap4g
Mc2oe2N4tVlYrb1Jz8OtY7CxY5HW73pu3GOzDrxvw9z3VM0D/QlDcfOK3lO523tl
X331EvG9Zy0bfgScOd/qTKBPKgHmlgMG4otKp+JPa9Kal4yNurWSk6tKtfjrNG5X
Fru6fYn8Rd/xEHLxEEUeMFGi1Ln9+D/HhRGR8c5I34OwRKW2kWSgV6goaAIDYsDy
7RGUvUZnC7B4vYD/CykiMAt5dmLIklbSckesEvY496HACsutmbFCj1zqs0+6vbCZ
1KMfGT6D6WEfIVgFI2mbi7PDvR6xo0N6b7FOk73904RWQAiEl2+gxrfqD5YeKCx2
RGg5Memmx/iDN3PUlGS7fQYh4g58n91PfFiO+SJLt9XDJE+Z+vVc21tdd4+PsVFT
i+7CRIIus2ebM61q5s1iPv58ju4qMw0UV5hWXK9HWvU5oOPOI0w8OAd1e1jWitK0
OekFEm6LjZ7+vw5ZLM7QZ71NuX4WDylZ4ctj29HrDTbF/x0qGPww2hmzwYYIvxr4
n9yIFRNJsrXHVS601tnHo+nnJF7ll3vbmvN7EjQShJtknKbGd7o5af15Nnyvt3p7
GWz+wR0pSnPQ6cFwLF87cSUYMwNDUfjNKIfK2Gk00A78795GqY/bEVaFJZtswpI7
jJFhrqCFWbH5fyCOAfPLtbdAlfb9pOuH2Zt0GGSMIGEpa/acdI8UycAiFQIU5RcD
HIBmS6cDuTYZG8/jyYV7zat0+/jc3wBaPJQhYnTD8yPaoFPoLO0Ip9duWFXg6mST
XZKJi6Q+aP874rPOJnqL4DGyLBW7m9bEgHX/UpjdCWZfKkKKL1biBfuchcEyzMwY
G4GTAZTM7y0epLUqiqky+uAx2SijBVKJIF8yFTukHyqNrg7kH2yujiw2LglfzwsY
UJ/RApJZTEgoI/c/HqP5NGFeK3lCPSmVzZkKq6xwEK1E2Ug0aQSToaFuuRJpK2Pp
IJVJG+uayZEvak/tYVPpQRLK/LBCkUvuzfjIGMSaodG2KFpExGDv/LUcjDoh4RfI
BrHxhFNFe5kBBH0LSVbbEQFvVnowlM/yRNPaw2WaaWy6sGo0Hd7vIwyZQGVfmmlG
bA+8wuX9CdyuHM+UODo4SOQ2PV6g/knbkx62PJm41IkoRe2bwjc4qyzWOmoZKT7c
nIM9BQuePm6GT+DaoLdSc2HeFRJQlGujxW+Q+tmA6lvaaLMKkWnTprkV8QB3sJFS
bLL07DJBCZKHpQZU+Od+utthk6YH1bTYVlgSbuk2LNwUkfzN5LF9YrrefpcHsUbw
sipk6Y5FcL1rDHtJgZ6IWO8yMemVtp8CGTSx1pQdwe+vU+NMBLEUMrQLMrDEXciJ
FUC5cLbZN7fq2as5mjdBcYyYVzYZKQ/5x5LQ6TK0/irF7A4M3QMwh8sZm+b5Iyui
n9p/PBp/ANEE4Tq3i/mLyM0fEgWGj8vGeeOINIuxj4bnlsLKsZT3f1LUJJTpR6h1
Bjcbt3SekAzkgvOKRAtsP8FFy4FHcYmIW+ZqTYBcFhXHPA9VNSwRa7nll7PT2ex2
WCFNIVykcKKdphd3ByT0AD9dydlIxpQohvQTqkA7gtSxus/rGYuYHzPopWnSQHtg
hkxiNUWS/g3Ss+E+gZIo5gjXUi/qbiQcR3G88cPi7cbJZnHvNH9H21Mh1PxE3o/r
MPvqtJFGYTweLp3+GMznU6rx/JkwBZrWTwwu0+HgY24MGa0611RFLV7tzxfjcoT0
tpIj9XP85YV4MYgABdJ3mCpZcUs0y7NWlXUy51rtXZz7o/jcmzv/+ZeiyUZmR/hY
SYrQI3zaDkOmTrJkyVSwu9CAK7oAVaOL95XttDX1Ks62xOu+TGqc2vHDmROmawEV
HMnNxauc+S36jMGYFDj1rds06D+DRXCYlTQkhwr2WTJNWvnO3DyFPmejsNpKztvJ
pEF7u8LbwPd6dlFLWozRItEhRIiCUZW2clvJ6TvQJQlsrcJKmH7ZTgxKBvXRxAIv
xr0DZUItfNlTa4JzQQGxxeAaI62kydsemNRmJbIBfDAjw3B6Zw3sYU7klSSWQjRk
WqtCNkB+cT0diqydJcDAH8Zj2Vj8yAv08HjJYeEvFkXyktwd62Y5focnC+/lwTIc
zqoYss2B4cPDgcy+fc4OqzwJqn5zqAJDD4aq8QSuTe2GZ/B7DXd4si5yny7BnT6c
En2Ho9mV38jaJej1gNdW/woxVPGW4wuuxOKyIEEtuCKG0EXDhiQahyJo9LwoJJGO
nIbg7PJRDh6aYTferuxREtwJDOrffYe3FajeGLyCHkIoyH88oTK8PGpG2IfpT+1i
+EW1zSao4HnsiezQXiUrJyVm9jM1EtXJbU/HG09r9Fm+aTux9FkIM2mUoYqLMVgS
CfTXKYrTsfEwBBfx8vTWR8MZK4QXS3CM9jCPCBTTxUtmv8slorfZ8xg4J79kK/R6
joVUPSz3cYf5eS9s+pm2rfFuX4mAjbulPZzeQetrMqmQW8SU4oxiBkVZK8mAjV/f
/1hSV1y6pCITLvZ1Nh/IYOlzBgbQEzuoF++mohL8Wi5aCYNyWSFII5mDeok1RAQq
ZbuYpkcxR0Kq/5vZKfqo6y4nkKG5jNRfJPWFAd04wTXUdSvVBOpgYcVtPrmtz1qH
JTAflGOAgurzlAO3QJDGjZ0gmTPXg8eEv1GXbGIkhZ3tLqhQ5PKEorLIko/Xp9gb
TG3G2qiNnrhjPlwxyvR2hNof7Halsu9U0ELlfw+LidOj9EM6mrwfjsE1tqMMyre5
HjNsQk40OzEc03mQNFWOYSxD0CO7JO94fm9mDoNS0ievJzDUZ9cY1d88cNVViOgE
2bTeCWScMzGPrhWrlkdC03w1BJE1SA1pmtth4U5tizgVJXtic+vQM78+FnliUJ/5
M6zEBjqooWus6mAdcf5EVnYpDR3+0mbPU73ECW2AjCMJ97DcGWZ/UoBQHvsYfcrp
/jVX3kbCS6XulZ2qwX8/uUS7yAcjaqPuMlUlDM9lwqgAwcJx7m+/Fm91fGR2c25j
NxMculZVQ0IDy0AGdEAws2x2BtE0KE2cakBQwgmDTsxXvRIgfkCMWuS0knMOe42r
kV9m2+XRO/Dqd+SmFXBohEeE2LRJvQmA6SZRvS8xTjuH6yNrCSj8n8SFUgmTgv39
OhZcOQRvZLpVuZkCP/IO4Xg+xzYlvM4XEKN1337FfK6TSSCEQhs1/H2f7rrG73OU
whkiZcOmAqKTpL9//h0zLw6Xc7qusonlI2KO+DVH9gAeeKUBUKirAqX/ZrpDJy9u
cQ+NLemAalFEE3I+NyVHTkN1GLPQat21NS02/F/Rs2pzeyP+KyMiN9FFQgFK/Hc0
kMTswL1iQjTOflXcDfuQs5fEa6snnqLi6uIyfqHYoSdE6g6hhKXdo0srO7/5os5F
6AGJdAhcnnAKZe/ZERe+6UBeJwGJYtz8augJMMVLj/Z8nYCDLdAbRmecBlhcEo5o
Z732aRY+Np91j3laBNbE0MMt73ge6ZSjfdF5/ttKqJQwiAOJnYTDYL7+xadll8Fl
9jDgAs426IjkX3EQqcjnbBUn3Zw7Kazojyp/VRx8iPM/xcoUfYnbxDshCI4MHKV8
akaXYO97b+rQhp0uubMiGZcAa1j7EkUHWrIwhPH2yPh1gieQe7ge15bmnbOIPeCI
jfaGUxGYqYSsStW3csKox4ajVdonD+Hr9D7YmhQ5Hjh7lvg3Ejw6nyNPiFj/lBte
wj5/zs/28RTftk5WR34YpbXa0WX/DJ2NJxqe5xyHrpmo4IMgyqrbOz4PSqeXeFgb
BW430L69yVe43UjaSQYtESn3FWUgwBTohvsTgE0GQH9BOXUVnRqQdYkQdXZykPO2
Vj7sqvjwUNFreqqgFFlMluVbBC9np0LVDZG8RT/Fbw5lHkinceGxRhYoViaCPD+B
2HLYgV0pwKh97Pl8QBnTOGUL94bPGE43anWAQUsH+55S7JdAGfJD3CmGazpTzc8g
Pg7gGy+rQFXcbcDNnDDxegAr5ossd9zjxsu3V8dNSXn9UZhNU9merxyniiOUjfGk
gZXbr5h7wVS3S3aryS9pUHmlqQTqcZYa5wlCso9e5sAMtClT4nwp1aOHYT8qo7S2
sAL2LuO7CwNs5KCmwRgrZ0vZaRFvXILRSpspqEpPOT9KcM08sIgikh4IX9Bp1e09
UsyqlNW36eX0iiNN2xVRnXuIQ6PgynpV7Jm3Znk5vDyaac67I2/0IGcXBTsC3CS9
AFrKP/IZRjoCeXUSNnSHpdDaqq046IVYae7qhT5gndkIpyo9SrFRtMyq6u+r/O7F
YkfHIgjfQpw6+38FeN2DKBu4wQxwhnXJn2MbaJf8MaAJqN/xo+nBzX7+yGO9tV/3
aYZLlIYFWZaIA3nGESp0hYMe/anrKZiXvePcloA3oNogoa//wr64zjOKZhRPkT/B
DMsOppK2wEn2vmhFHqjn1QRmHQV6nSb1OjzyITVxWZbszooh3lLstAAP9XvyR3mC
tZo3DLfAntiNBhFl1RV2OQj3WHQlVYS0xyrs1fG/cN5tSCJXGtaVyNmn5xlRRpEI
R4tQWjivq/IB9/UrH/Y+SGQGuNUprOE73ADoSuC/SOVll8TLGQG2gpvSMcs/yK0f
ILMYDU4J5Sbx5ElsDjprVZHvgrOlDFFluoOR4lN8KWDEYrzGAdw8HAYqJD+jC38e
weKdpZSeA20b1cM4LO/LqjVQ5zuxfpddc8EbiXX2M0/N1VnMQeLKhHv4jqc17pbB
MLC1LoOfeMs42Xnf2Ri09svDajzb2/F8oOm+2HYpb2oSF9BawrqvlBDsfJXLvV3r
gOxRl6X/rAQELMuQBBSXAGQQJaaQc92467LhdAAp8i6SlC5xnIY/uENKhO5QLgZ/
y8279txi38axDpnR+78H2YbCeoKZGT8A+zV8neULl/0m3OGgC2kK5dk+HHaxAz8E
qEmPLURsGmS0urL0bAXO+TeELTrfVyCb4kH+CB85dn8wdtIcBNz8MfEs9By9tzVT
f9az7bd6th+HQ673Zj4pHYFWehPY8t6+FOL5vhvHHksjMhdLOVfhT6SLdOnYsSU6
8cOkQRYZsW/urh+2MkEKOeCVjv8MJngR0QPZ5Ml/xLSEs/PHr/cDSkmGT69aTkm9
XC16C6VsPdLkNKotkoEh9sPrqgbiUX3NyL6WrM5hrAvLf0+QWmnLu9Ib/fEJ8Lrh
o1qHkHDyaTJBKqyVYJpDg5lxtpqeuG3vdRqGamNbvRuqqJeXsq8N7BxhQNpH0aZ0
FIKTfOcT8G8r00dBval/VBuORk5N8xYdk6kUnOLXoT6avkh/tOUeLyXqvoRqVLx8
0VZzVE9YsiJF2UnB6km+zNl3lWdANHBKY5ZfcHqcmKbwaegVWOlX5d2mc61KRXRI
EBwaTQRhBVWBeAmyKY76abR+OmYk1RweI3CBmAQz6kbhd/tulF47eTFecUYwzA8u
7B3+R9v2w85JoTvUN/ZZAap8xZ/aqHNq5VxNO9yhe0U0UFHV1ZVbxYKGdWXtzrz/
HO9A+c0GdXppRVoo9LaLdn4CPgoXdR5CE6aizxL5s8+pQ1CIva+GRoODgfMThGLN
YvIeqDyjGd+Q3vYet1qUQiIp0Ht8VhP1dcq0vq43YefAZ1h/7xfHTqPgnH9zF8Zo
cuYCL4be8Xb6WLk7icIDvYNNnaB1zMlJVujlbSoh4e/W7HO1JQsIFBYSmhfem5eu
Qu00B1DfVC/QSV2EpG3an+lgKtLxNxJ+OSTDUgLC+sCuv/Q49JN6JBw4LzdOjUQi
uUqI/SX3FzoNFYByPvn59SoqBuU6EzlItwU3vTZmIwoM2xiWNu+CeLdO6W5yKWCB
EP+7sNAMXHwrH8rhxaKWoeDEowDt4maJLaw8oDyWEcOIpgjvLfz3OAU4TinndhrX
ylvIJ1zpiOi6pVpHJ1IPSqntt+udktLf2wiPQocTXsMpybvpMjocOMr6GiwWH035
ZmlCd8npxRuSQDnh1smLJfLYHRDl3KkyKDJxm9SgJq+Nclpvr1RUvQEH+AW8DYuZ
AWLvHhoTkjvwYmYDj0JaRpqdgSMx5fORGyaDLgkjdSTdfBqUR6k0VppfxqLJzbGp
8M0JDcqrn6D2iM/i0I5fd7mFrrUJke9vFzMlsICUs0qgwCPISFx9m6tqnH6eThGd
kjOy9RNEqFL649OkG66nCrWkFZGW4hamPkxewA3XKWBYn2GkRne6lDysj26TE3fL
JSp+J4h24yqSduI8ergSKONFaAuJ4I/Y3SzObJNeNBjQw52X43YeoDO399I65a2d
/m4xMu8kh/fw9rQ69kp6PzfEdLvwezlPq354QS/jdhvghJAbb9dAcs1/xw0+pbCW
xI5wnhMpt6Yv+l0RG++x85y7UbJYVCBbkpvNMB+AqMihm12XBstOs7orIrO8uumw
ySRcF4z+vycICx66h3K5PXdrMXE5qsapC3CwY4/RBSRxDV+HSYzxyzUDID9Y5iB+
U5OQhfYHJ3kLZmOt9HZ2d0UHki7Q7Tum/QnIyzhFCh5jTcW0vpJlEmz1tr+eHKvb
Wb9TakTd7nO+sTDJ5jq3q2A51OidnM6oimeP/e4pweVjFZIFwjAPRXLslOCgyMq4
cMGLf49Wui4T6dYtNr9glCOzQfKnwkWraglbKuPH4UIl6osp5ftpalhsMz0C/h6c
2TUxa71LkFFTwUiO9LsGAFvNR/BMrG7I2SVYnVCW6r/H9/1A8cXMURmNrR/Pmd8o
GyAcvuELej/hM75ko4xtH3tT72ghJZyjpMZ7EsgPNkZkeYvld6E28wnUgWlWA3LX
Bv9rx9R9AHmf6qsCYSuPnTopjHYvIqmEow52F23m3XoJH+pKcLXRKDQghb7BuhpS
MMChJTJytVjE3CX/uwPhx1Yerq5F/r2JPQorWtx8CNGBfBHFh3rRPam+05BXByoA
88MI4xJ4a2u9/gbXr6Y4VErDaQlpnclNCII/lImK7W5nQHcTSViIEiAO/Taj0DPI
mSN6z5utM3EfYsBWvTNc+1xwJD54wm3rsLLXIHaAc/dmp68xGQOKh2mnuBMs52Z+
MRnEK2XGA25QhTnrZWj4iWyeFtqVcpKqW1D4W2WA9CK6lJ1rVCzpHGBMa/4eHJ9B
PCrZd2lWTKghcS3y6UU6av1DvcxxINAuKuCATVMigjcZ4LYHMAu+IOMXz7ODQTjv
REBNzT0Dr0PJjg+fNba80hi8ePo5Gqjmmz2uXYIum/PBT7rpZfKWfX1KlsZFwzRl
qlNoBL5o8Fiekb8Mqk6uYuJTn4/BpJd+9Q2P3C9RRS4ZggOXhV2IaFL6NRy7pjQL
6prXWa/z0JhrcWOp/RJMVLJtE+sNfJlwe3hGvAxIOQ1IWrrnEyeLB/AlRoaJVxd2
qkC9jxU5gatn0lmezDLkSwBvzka9ikJcD/b1PcvrzVR/Qk0AjihL2I8osXJdr/O1
2UurWeM3mQ+8rbwrBGG3aFIvju8EAudD13rDLnsQYXmWwkaUwEUQwp41Atn5BjA+
v3bkCRjZDPqAG7moPuVmHq0B08Vq9qRHC2SlorZiMjHPojEQ2UtUkIWEsC0CB1jz
rHKlvO9K9Cj1ZqqL69wHBL0ug0eaXjjSc6ofBpcicv+bKetzh2nNVBknXJyXVkOO
wQ54dA2EEococ/SbnW2p1u0zv3B/PCLAGhJCY7omrJreqflDqUt3cYrfV3gvfxW8
bMtd8KW2Bv9d+nRVt47paROoDRPCBC7Jm00HFuqS0GJBmbmsgfMDlownv13NMEMm
6LFdgGk64l8Z+4CAYSCw1ddxNWSWguVR/FOSsgZoos7Ta7RlOo7/bsxlZsRGeNvu
xspZeherp8aseVpJoLbO9cpO1mJV7eMHqZRWXpMqCEsP/SyCyIFhAiOYxHPcUbJ+
KNBsrRJ7NlCBTq2tQn6q06+Tiw+u9wTl/RyvzfUZNGgod/CnErunjJEgF0l7X3Ft
C2JW5yFhhQGfPU1QaElW/1EDmYE2xRgt+LXHOt8J2uxbyFmpzDHB6KG2wP8a743I
EGIHKGXCbT/8Q1qeHLG8K+HeYL0R5ZdB1PlHvY3GMRZsTZjI18IdCMOGTyT2mGBh
EJH9tNZ/oMARN/8qlN1PeC3H2Uxlw6PpEs/NbZCV4mT5EQRflO4we+Z8QrHeNJEe
8h/xbBXzkqX4sfhuArKHUZv1sLnEJt8z4q/TSpmmatAjnW/xoD1FbiwoVzhTJ6xd
ySs/ubyHdrx75tAcHiaPrmQIOAR46khGlbLzFgjkK8g1+2YQb9hmtTrp5/U8iPuH
bjORXwB8vOoZTpYL75gp6dX9sAO/PHr+quaedMmHqoyyrXZwamjQycPxMrS+3VUB
xhxfSLgDJk6TIFs/E/A7ogIAwTyapdKfDYg3nf5mu3mcojFCrkOimBoA08xJR/ie
kuVaoLLUxvH4qxG6VqcPqgyDY8ZxiR65R0JIrFbNBdGhwh1+XI1fFPOIfUo1DQ7A
a54OvMJt7pRvxuJfemVHJaQ/MBmT0CcamERXb5C8CtedaQqsouNldzkam9lTFROq
2+x6HX4TZb9DgXYSXUMII3FFvuB0s3Fi6fxqAXSUGg0SwIknHnjI70++ld2oexv9
Jv5IyB5VTTGbHu+lBW9+2X4SY846j4zyT7PvKxZet2c1VH/NHmjogSx7bvoV3nuf
L58ffnTVRFdlF48Y6AO1lKVcG51l4qH/wzUOAD8ahAZWiNxdZWExXXba7uhsC9M/
MjxFa6nzbBP+F8OmTiFZaFQ+tPFBw5MWPAyJmwr8jdhoamo4e556kZbPksdh3adt
J2fAsx69tR7qCf+Iib3/a1huHMWyDQend1K3H1XzPeyskHgx1liGI2ldgyzrYvBg
pNjt0tE8n1KYAJ9xIZpwxz8IL4GxDG8J5NlJ5W2WMiiQPVp59D6LGwZZqTdJ8nIX
R7sQpDftaAy6tSqGuma+jTUEkkjN39Oq5LebuPUbr5i9qeG/eWotoX1bbdZNqNV3
46AOcyiNPlJPgDMxhZlao6fbpCKq/wH3oOduLJL3aFCs8OlHGq+gYuov7TMLUU+D
BIKQrEy3JqVFJgO/HrcwEPA2O5fWD3NQsRCwxGnL1EN8p88bxobrOfBMsxDdF3e6
PxfTOSsx0HZJR9bjC9eE8AVOoEl8dIYA70sHQtd2Map1jzi+hkmbz+1U8KqoTfKD
IR6XD/ytiiuz9Fann/yIn0BEuGuFU/Zix47lJM3vgWFIe468troAY2VSzr5g8Mq4
c8CUE3znm0V/oCNrTL1XomGMTuDOAlJlE9zAE4I2M33W11KVmkvkJoZtLwbkgXaH
UnaeLgUoW0lINZpJTrwYGkvLsnEYYOnjAENnIIAuLlRa+0A1f88YZBStTj8zOl+5
aEpPWUMXvatFPUxDyw56wCGiUkDVWX527P4zLc7Dnp964ewoVb6jYQ0Mc/cucIfQ
ozS4uDEtp7DWPSh9ph8o2jbZ4lNyGoT/gjZEnha87VHuBt8/lOGIwXUAejxQQmez
4qtWFAWNbSsYZQijm5WE2FDepOdm0kgYhUvDK8u4pQlaVb2KVWpdScEO8DkwAwOR
usx0e1bV4dPqh2Y1/sbAFesB5bw8APvKZj2H0zXr8hIPBrdBdx3Ksm7dMuFHXOLE
VdMfw3AjxUi6x3jPgYiY3cx3qgJBS0Z3dMg9gtLNm6cMqfmoLUNSKQF0iICzcd6I
H78cV2df4OQSoWIF9YE85n72HGwUvcpuS525RNP597gm8ii3iNvkjxWANEKwrVCR
c4g1sFwKYdB+qqtyUDWgCnkUbTPPwsdev/dFoe1/fXydDtIhhXilmZkp9hM2eIDx
I/sm7B6TNuSdM+ab1oDWA9suHklXBri5nwwGnDKtWZEWPmadcAgEvsnRAjwW78C8
P5Y0nxQuepA4BMOzHLxcW3jWjA1wC2OqhKZu5/P0PSoj4qFix6HMMElpeitK9xDe
f0re0R0aDG2k97RFVgLYECRXFBtegV0N7CJiFmi0vJU90EJcQ10LCevub7E3PCF1
x14WXPdkON3ebSlS5C+CXM34v4xROXOni/mbkkslHXO6JwFK0XxTQClB8bDHofn6
wrtR9t7EgCRdrzPDRwkr9HhKObK5c/6JmQkvXos2kYX1G3Hz705lK6+fkWLqlbiQ
3WYXQoKzJ8TzDc97BhdRBG6rWbjf/1shwuiPg9N+eJijAL42C2wiceU3jrj2UynG
LrwbvXk/wPGiISiWJHPA76lCH2eSOgtLuI5QqONvAg39VWUMIno6C9rON3Ty0UM/
p2pL8SsSRULVRMJsibbSDN0yI/Crn+yQRGTCHbBprMSS0fC4Er8rPfM88QJH5a2F
wnfpw6qNg8hRicjEYjgBsnLuUgTNb0E+Q6sI8Q4yznh/Yn9zKOAvs0evRkWJmwFT
4HB4DjhFCcTCsPn96r+sv7nRreOqlWikgxyJaxgrvt6BfHO0J1Kj03fnaE7FUb4n
RyAjUdF+rh+LVIlF58b2bBA3kvsndNNg0CEPX8zgCufQ4ZJy2+xZsr3PvSo1/qfJ
GLl8IwK6SaYK8O+vG49z/EgmyxgBG/o+N003uVTuKFYndBbgmLi9KYVh8UQHUVYA
lINWmEoa9vGEkrBDER8VdYe6MVpZe+14aD6qVtj5B/uo0ch2dLhHjbTqnEtay38C
uqIrEv8asy+Ram2ohUbcCBvGKW9Q3RPk2+nasWx4NqXzYWehLitEV4Jd5zpabv8C
Pxd+FMiLbTFy2s9IR7ZYHQkYrke7OflM6TXZ3Ld5N7EyzBjR06hkS++m+NOgJmmW
YVOn1xkdjeer2dIli3xECBSW16UJQtvwaMfw15iROBiTv23dTKOEYdHvf08tBFsO
iFFe7NKu+0YPGgrwduSCzN18TTKAiMlRBRgwTB0eraSVIYTOwQ4B9vxct2xBpF0C
UTEQW1fviuKpVRb/n5tTzDPekDV9/vN0/VKl6PC3Lvi5K91rn/Pi7568A1iGJiit
3qpqMLAGQZrC6O84aVOWpZLFjevNO7DDJhMlFdtCRFMgQArxWd49omEHAkoozXLt
cDRdnJMtllU1/2YbCRdlcd1gaAWDTbb2NMzQdbeqc5ZJg46Ug4AHr31ZbtCi9BKy
GTWYPEIBDDU7zn/pZGEWejSVlQPxOBZBCRiwh2Q4BNHRlLDyxFNl788UgnVjKZmh
JBV7vFJzPFWK6KEz9GDEeBe4Hkm6Jm1K/l+Cixjx0gvVvV7/r2mNxgoyxNLKzbHl
sEKFIThtkJ6tQEQfPTXJ/gnSLDDfwgAUzjKkKzoDXaJ74OpNq3XQgWHl+flIdeal
RFJe6hHwugVzqWXddyAVLJr3ylR5g6g5QkvYg9740SHTMKu+zbtNwBf490Mbv0xC
WBvVpJY7QG3QWQqLzLskpanEA6rODOC0Su+dsQrgqpC3OO2yQnTsCJY9PQ/Nd/ae
r/DNwE8AaCUMQfkwjrX8Bcf/xx8RCHITkpMNp3dnlHm2TnLBDrbkBV0fsa+I9fFU
FrL6G3FzyVPeBUkFFlAhvC5DHA5zd8fz5K8S6A6DhDbbObOfYAhvnsQuVJcr0/KB
Ps7zqFqIgkW/o/6R39JL5vdT/zKYZW/UAwY/cIv43aAxizuByRpjjPdQcOOiCceW
JaOzvI8cXz7vHNy+SnGKyCNaVSeWas5Tk6ZoMFXyw9ki0cOZj4Xz2QDa34QLHE0F
mCXzfOo963uFoQBkRbyEDIWqAInlCSiphL3S0x+FeVNWmv6JFXFdZnuu0DyNmXju
hk2yVTJUH13CSody9uXgiqxLUCmWiJYPRZQj21l6zcIN5B0Fznb4AYYRUaseafKg
M7hEEFMVQfYMJz0lROP8LAWvOuzlGMHJD5ro5PqopS8sYg2CEWWbHxduz5A/rrGO
XY+AbqW97UzaEr6CFGMS6zBb/qgORnvdFm+xuJJVIlQJBo3ROhHsbYjLF6L21a3n
EfZEeOkGKfAnDnk5SAVHs4Uj8CPi/0wabJ/B5FSzkXf+04Ll5nvWYCCW/XqOS9cw
jmQcFR81MDG5sWvZm70PEgMXWNkEWDWMbUMjZ9ThTWQ8QzFMirqSy4MqlzvWFEcC
cpG8sAoLkZfx+qXFc/pnR5Dz4wXOOueLiREwn6HYCLDmJl8otUXic+t2sznPBIZZ
rfTyGhXsa8cnKSVm/k8gCuWtrnsiWapSXiTH3uqZGL8mSSRn222MgeCAIscKWLp1
xzTiVw3y3m3ssRqlK8Jp7HUoEDRZZN8S6o8/vaPxsnhf7cgX2DzhGIRrh71wFLU6
VFGhOsDnhzgRIqFWLo810uhxaAWCL0ruH/AulAHlJDZsC7VH65bgPnOMSjd+hfD5
rZucoI/pywypKZsb8bnG72p8HL+6hEh3yzeTddHTuR5mG6Ii5tt5E994IK//22Im
36NqAeumM6km+EFnnxQ4FuB8ls5tXBADBdxtq32lYHbt+Tm4SQPb/aBCIsDi3Pic
ilHhuXjUcZDzdxtg5RkCKebw9ndFTDZ5GGOOTJSyroftUlA6tlbne48lvKOBMczx
MlFy1yfIyySPoziNwEW8WqXxmvi+6TM4CEsYSizpJMdw00Os894/ZDw3+z9L7EEI
6PbS1PsT2WRYeloenYbR+E63tM16SwH5waSitFNXtsUFZgqbC7gKRbAVCm4T+GKJ
mLi4yha6WbRI+jioquoF0+i0X0vC1Eic+NNadHgK+Dx4H+u5N/fB63KbABOK6lem
OZ6NfM4CYipNblkVYcpjHBVgv2EhYLJb86wbQ2OlQ/gYojnfeU3ipP1bHaPsrdVN
4VzjQ11eMY3AykZPjKYaTTR44amEIPBZURt86dDtMhwn/u35coZodb1pxy117JX1
+I/BIXibNnPk9SiZ4cmgorlCbmNlIZgvX8CyEHIH8+pMLdo182wetG0MS0MEqYv7
H08XvmMapD60A+vysgtGjQ87DnbkDL5VXg1MrdmlIOUhJFKuTrRK3tgSgsqSJk+G
I7zvNNIgeFdnk6Vb02991OWQHuYTkJY/rXXgRL0G8ms5PcMenDLSz5tWNXobC97/
4qDkQu1MgESteUVZ/KJlougILmoLrfO6QZwfqILi1LGuwvgOhqqH3xdOodhNfnmy
h7BUEDg75UIQqOk5GUhNXmRK6S8+IdL2DCsBGisshhOpgXSwyZO2pAzmaacuIPFT
74IrEOSwWoV0o2Kk71erampi/E/5u9KlKbNvMZXUKQI4o+Beq9/iFKA+P7cpMdrU
2mznveUQYBD5vFYXHuof56BsqYIf1KkhYFvXhvwuCBV91V60iEvQPNykL2ugN+DI
R6m9mqAVc4V+cRZa6cTFk6nLMsH4bKSbXeF7KrQ+5ySuSE1jEfXuwYnXXwYhxnHv
nDC850kKbFYfK+0VV6BIPX9pxoKHgHMfMO43nWGfIg0qycbnXfSnvzQKLKETubHr
VHgzyWghgziIkq+64cZt/VoAfdvwRTHG94GsM9BrdrCCBrIXqSLKTE6/06hb7O9H
A0q2BJsKZ5nCJDNji/bxWnpo5oG4kTsvGmTbF/fTzA/PGYZoK3mgV2oaZgX2S5Ey
mF+Yoi4kd2tbvjeDgg1wU1+9Mop4Epoxi0H2P84B7d8M051f/IqZgEqENuL0egK9
+j1v77iXzkmcQcJ1+X0NKFLoFVrhqV4tET8nNYBr8g+rbvaOCCmWZVkHGXfS4oq7
OMEtx5/i1mmvgcpjGy/PUisHoiJDrE0io2mmfKG/8RfNWBPh5AVSWkziGkv5vDWX
PZqP0Ek6zJYw/SSSgdsvvmk9Gh30CjKxZ2oG/PlKWkPn2wzX873Uq6r0Up0DyGkE
x1FLxdArwrDF7VDWM8eTVAgDxMClKOxk9yBqJvlDbW6YdXL9LLQODU+smiWUUwz9
ymd3JollpxlkE+56mbjMLvZbCdaP0vrQeI5W2HS2aLj1xeKg3DgWL9MidKDo/WQj
Y+GRR/nY9Eo0521RTxKVEJAyjK+mqGUdPBOPr27OHnw5YO8UUfFHWNO2kolpdrnY
MhOz/YXRZOdYEeuJBCDqm+jesA7O4pnuq4jBfCZbKF8h7IYQd6pV+swTvuzzB2Xf
vNdANZn/BWL084MoLda1CZ0yN7YnIJkllPweqIYVwtaqlH8U5lggbKmo3pJDMfk4
jiDhyFFlBXk2DY/wveS/BazB5OEhs7wtCCcybqacLuYyyH5bkjDGz6D2EnvyolHa
`protect END_PROTECTED
