`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IYWOfdhcGmZ5I4Adc6f9d4WcipTEFOOosRKLuizomOq4m+QUsSV4LirqL8bwOI7I
pj0FQUsplosglnpFxhTPgDbb0h7jUMW0tc8ry6olD3pSn7b1Van2A9LDXnEA0e6W
mgfbTe4+PSDCf/YcovmPZqyXyCJb/Hek/O9jePgT4GmfXkoFgYDnT+KPtSSotMyr
51Bu8nl8StjxW8bMendZhhCzLgorO5nLZKgqHXseSmCdhc/4QFKvLzlI65RdBZnE
lzmGj0qlgDrGF+UZLVnrf5JpWvyXfI9br9FPj1amIY1qRtAZJKXr6UKTa46GR8bR
q1Sh4wsCLLUzGOfFSqsNcPPjvG1oemJo0cfxBf/3MMv2wik2JbZCX/pUnkhTk4gN
4rWR854un6bWHpL9QX3sSrpCS4mjV+v+Hagkbfe+dq0=
`protect END_PROTECTED
