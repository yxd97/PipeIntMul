`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEB5lIKydP1Do47SNUQOfrZ7r4CN7lVELFPZdzzoMN07EMEG0y8l4Ge82Zz6f+pk
Q1p3pp97VaCi6XmC8BeOadKkgCzAAEW55dr/EWN+yt4hwAct1PUhCaS2wPeowHr8
+jHTqsKUi82cLRVcf1zltc5Y1HvCsr/HQJjpWLhe+6zV2r3txxmI68um3VSf3noo
nRb/F8a1KZqVTts/AnVBnE7EhxM77NfGI8pu7RkPC/cEepNj83mS22sf/sdZYCAt
/YwxTHZODdFuaP1ROT/3tnJMArwEM6f9ToBXPmAWtvPYNQ2JCNS+UFUR1rmSZw3U
/GkyW/wyDRiaMqX1QWUx8QF+pkPX4KW0ZGteUE8/BpcBE6l9Oi95rHLsbXtayA24
MnsLO77ewxl2XoYdYVpoTkUe/CBhAememWLJ4PJtpzBqmsjqFm4RCHjMHFCwYmaQ
Fi7/Jfysf4CDretp9qqnqH3BVoL9FzC1+DicyEyrh06Nqsq3oeiBXxZBzH2PpkyS
SbKu4gDQf7lDbF6fuLQv3QzDAiBqgo6sk9gAjn+z4yNG+uhXJb5xt+MXnYJgAVo0
ZVSlcUR1+JLChHkhtXz95VBSs06eHd/xFJWV1aVtixxS/ULB8E+ZTrM8PBucUPds
l/3Y6DQgjMsSkJOAHxc1N585BIMBJHeB0Vi90tmoBzmOepqsDpdyOdHfi7BWQkhM
qjZoXYMFqhXl43YWoLg891l/LdszrxJ2Ms893L3rymDqNlrcDDPXNVpjuD+34/Z7
TvTA77O5l8rJpqtTryfivALsfXtrrogKZTNH7w4WZHI=
`protect END_PROTECTED
