`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b2Bxg+6LiWdRpq9EKki27zwiU9Bdo7E6WbHGRehitTuaF8z++1sMcMX4663uHFfv
v1koOz7UZh+NIgKrnMxB1FA+rfR+AfAM8JjTKmAX/b0eUrYPwIkTQbkZEWOrNu9B
hyGFZLW71wcUsUwCY0hpsB4Z22qzbnbT054gxtxBWLN8TtnpFAB+9+wNQXM20mzu
fVP+1nqdzSISSo5mqumGJ+VQDCFhp9/aqDNkCvAg1albqNDXQUEy/dPx0yyjFwws
VUlgbr0CQBR4jU9A7eQjikZDmSroI9PQZhvMSHdKN9IRB11gkYoS5i8givhbhqEH
omzTn1tdGLWLKtGd5qdjd54mdTfTsDIoZySn3l3d8n+/tVLTT5wI4d8ht9dxde3h
RUFCGtdcSPeiDYCCq9zaD24aKxsxa0KYWRRopHehvsHtqEzELnT4m8BmguDFS6zq
aZmIIGwUDrTVW26yyB67RVt8+dwVafIt4Fe4WdBhBtJ0WYo802Q8nYqVfgsvDdqZ
mE5WECZQpEntptvNOxtCnOB/f5QTR8nuhzDUy2szg258AVRGTfp4zxLcXgdNQmDq
UohSBAZin8K0UxldYy1RPLJd/mvusp5UT9EmeE6LbZa4nBQ9+scLBv9vg+vvxyM+
+ePtawgbYA4W2vpk1Kt4UYRGIEYdOKSO1kpv+vlY69mtJ0RTOWJkFIevZWRwof6q
qsb5Y9Xz9gPogADeZLhGr0I0SX9B4+vcJ1HfcZTB4Qlj11LulPTUoIrtgr9RAmIx
m8waEdD4/EPU898sV0DEYJZaadI4xoUuV2uGY7yP8u/tc1kSY3bI7achNDPBR5jr
PslvCvoIJr5+I7oWVaX8XQgUjVE246p66iixzU4UjF72rhgGVjnL5opaZnUwKZUJ
2k9bu+isBWRsi6XVoDZXRIdfmLvP8Mm2jOzES5T61Vxtu0b2CNDPI/SCYjfhKJ9V
VhVvYTUlXBMXRfILsg8eQY95v5ZrWlJErxFAuinvSJWJcqallQlMNSHli6PlB9mj
DXAtFfQ8doodSKn2AWPKCIX4I1axetWYyBIXzgiTMmGuDVxBKdrzWWC6gYaAlbJW
hrTAlXcoyDENoVtLBtgDnYBk/5AqLPzmWuAOdztZIXxIind+wasidWF5ZaDgRR/1
5kR5qtvmEGZjIoqcFKpzHjWeItN7uAxZ8ArVykzKlwTQAmod2RV4WCmnLAJZfVA8
mzg4INjlw0+i65QMk18FJqf+GJFK0UIdeV2NoGO8sgmFIWJTaPF05rBVFr/5Ig6T
p7r3aQRt1/1JMSjne1jYaDS/CWSk7VWyAO7TUUD7L7g75Llf2lHSy1bnI7uA03j9
gppiWpqQAe++e38s+S7xQH7lsHtSgJ2dD6XorO7SOFa3Uwv8dD2AFIynt9ry9LXL
8vxCL9GfXC4ZknuIurd3ckA/wiE6Jj/7esPREJxwAGIB8vG2qMUr2bm5CSTYYD+h
RaZZnCf+5vPx/E2Lf9PvMGOuG0OGzhAPTikGQIhmxswjcA2GClKKEbTdi2B87x24
OpO5Kp2iznNt2JtTn5MIkzOpi7OtdJ1APBX29Dk7FwjuLWpOd5UX/9PSNVGjPgP/
WxbnS56MP+T680Kh0AktW1iYTXkohmd6zIw9QZzwTiueoV/Uto/WpNhh/PLLsEuU
u4bouzcWL5At6PjKdAi/wptnMqY+7UQwxs/32Js7ezxP0Bw0ypjZGZMwoL9HVZmS
VBFuYg8ocGOoQ9b+d89bdQ==
`protect END_PROTECTED
