`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CBH3NCdo7mBxkiMoUcT9czVOZ1hoDOta6p2LBoanEiWGietFZljnZSygc5IxnBGk
JE3MtdwGd6GZtqHjAUF6Xne2L8yiC+Wa9PO5NF2g/eYABc6RPTRlbB8Y8WyEgEzg
XbYcWNRuQzfrAzZbRnZE8VvnRSDD/BxsZ/HM5yHBGLcnEtTuUN68R75Z6PSeCQdO
ZG/YpBXZFO8qSb4E3Hch1zhauBiEAdyLAx6IL37RdP0EeZkooqm2FMUzd69ASggw
4y9qDK5beBiOg1AtaFvwlaa0bTTTzCx/vpniJwTxubu0xze2240vz0nF8wybI+wO
zHGB5LLkwTyAGB0TYZxQV/kdaGjAy+Bavyu3CE8SetZPo3vxTSpb997ivCBZpcS4
QZN6Toq1JJ/ME2gj31nVWQ==
`protect END_PROTECTED
