`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/m6YPRRR+y2U33P18rSBs420HWj1IqqeM1pv78k18jmq8Htdmqmvd0/iCfkf0UVu
z+BQQxN8TtY0ZzM33onVRuagVbePFbr/L1oOWk7qjExWan5K9wSleYOQZFvztWUV
FB4bup7sfzlH1yTGHZ42ZA1rgfclWvocrTJ+vgqnyggGP3LsLlPejcikpi/gXQa1
2zhOXqVtH4D6gfmo5PyXD5QXAu1V0ACb2XvFouFnI26CmmVLyBzUULZuispRSzRL
V98C0Akn+cYp3JS/2rv2d+LBsfPqN81H8wpc+wlBgGlNpzuX13KbCnJQpGj26Neb
jTv0YNEJp3tnufhoqSnslL4ND7TsVZ9Xfb11tuof8stauYyCOzzemBpjFv/+OFqg
TYAuUyt+Jdj1qFsTigntYcjB7u0rRqO2PZFE6Er4qbbGvnDptuzsGuETz0LHYnH+
8e1fxt/hFlKwrwUUI2xMoWPUyDbjE+vCF346G/sCKiI=
`protect END_PROTECTED
