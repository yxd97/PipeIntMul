`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsPXbBlMDEnfC8zHv5s6ZfMO88kCCacUfaIDaYhhWH3SgaJ0rV41ih9jhKyoirNS
7d4EAsQb2FOnqMo3h9S73TnSG6m3TUq2hodi+xCQiNeG2nGywHYORKmECDv17c9h
NTkHAlc0c6DA+I4xPXjEhfrsVnhATNl/HEyRn7dyPG5ilnVXXBvI9tbfd6N3e/hV
ncVwTJejl2fykTPq3GBKekrZQ+8DLZe8kkoAN8Cxx+OCGeHa+Yi4U4hmo1l1NLpo
8CHnLSRkC2rq17bBdHf1kLw4yefJW0Gb2M0FZu/K4X+61XdWVHRRKIszJrBVB7iz
`protect END_PROTECTED
