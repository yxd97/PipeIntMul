`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5FEqB6DK8jO3eM1Xrabu2pZfPct140ZNWKccUcUrvi2/UqyUNS0uVtAhSr5tCpqR
GPCLWmA1vUHUK1NTJULLM2cO9wsTin/UOEMm6+0gsQBKR9yf4U2o67G54sd8maov
xEpKOe4yZgCqb7wTj+/VTkRv3x9pnNB0EcEeIGGTCa/fjkwgAWQ5FGRHdDNY9XYC
BEGvvNMAwnRjdlyfhRsLU2anSKHoWqhsJaYa6dSoZnBojalDc47D/FrSoJqjTQgG
pDyk3Vaz7Jf2KOPA/5BRntGxLb1Fytwu0jWhMm0AjHo06oA2l5+V6tfYEF4bQ9GZ
sO9CAiJ8SKWhzRlC3F+Yp/btnWHBeEHiX/ax2IzkHa4tqmTROJaWFzYQq6zrsyE2
MVDVmVTMoTOWePXeiaDjLd2yOtzVwadwzH2QNocCdMBCLgG7xaIXtParR++PM1s2
R+3/4vcTx10y8oyM0EkTVr8kSCwMBBpnY93szbnWTlU4laDa0QhMTQ4yRbVx0C4t
D+eXS3zGR9I2aGw93jvbysdkR3A5wgYXIxdBD9z/A9jCLQXwOjtJN+0ViCT+R2fd
8z3hPOiO+3/lKoo3LrdZN0nHtnkXSy0Yno6Ryz4dFfY=
`protect END_PROTECTED
