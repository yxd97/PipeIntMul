`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gqmvManvKrBOEh7MSFec1K/xiKpfVGTMarL65Hpm0yomToOTN/ntTHGGNVeO7XzH
4aXJbfoH2up1Ea5/c0PSgTvTaaKoH42ZJGjVRw0JJaGSgsTAvffIneBgjvqYsD87
9ro0zZQBMer3KbqVJhD5o0OTn5pZTnibMeF9oXY5aTdu9lYHm6+ZJqqGNYjxK6jS
acetJGFQ519LXbdBgGoauu/IXIqlvi2XWv4+v2KvFjW2Gmv78T5PdYNoEYxmWKQw
VlYOzhja/NCOmvO9VxuVHMpNFn6GoEhdRl4CVJWgDU17x/O+VdjJqjN58mopjxO+
COw8+Nx5q72ECNaysG3fYhyojwYKZGCHIlD0YmypxOYNSYjul1zokoDIt+vtFX8Z
F/dJfZeQGgBgv0UqofrtiFA7Hj0FkIhTR2XzhfIJ4GBEYyBgMLgk7m4nZNPDUxDp
3ZgN3v8UQj3NIoeXap3eF4UYCSj4zUaTWRU98UZW95ioB91spLKRyThyvv20n1Hl
XnicuMkSlBh2lvBTq33+rqqnqHqPqFUsY5UDXrOuvwgWVG5wtgxdxvhLBE9v4//O
Sr4Lh98Mum+XCOQ+CXC/v6ZuXktW6AQn8RFW5F/mD3ZJAo67FGz7lb72qROsH+HP
2P5VR13pMD3Pcm0OfJ2MVTqcd7ZmiLsDVa75mqac6olBaCtMbNGmTAg8Xh+YDV2l
01fvHhOfiuo1A/cI5dCkzUkbF7hmX5sjC092h60BifxV2e4CzJk+h2E2k6TNjxmA
DpZfMmpUCvsgNGi6wY+nNbO2Pi6ng04A3IQF79UrDIYkZxGAnDnWLauUMYbs3Qs0
jGtlv8By+Nyk3o/a3dM1MQ/cEd9sWcbN5KfRk29VsnOO7tpVmVGLfpVdk22JMj9e
O3d+I7T6Zk6nIClAhz5Ewq5F6VSP4y+G0Dyvr1OL9APmARGYK8C/sISt3WVrbGpW
cvRrv4eJG84XYazYQqO+FzJbqzoRg8ODHl548kecRurGxHeqy80mK3z29WSSqo7+
KtYtvJzqX0QR1gApBcqy3Vz7OS5X4QgkI2Bl3I/0RjZJyx5o5ZPTrWAi/4uoYidg
BGmIQv+XcXcG86+NPCxFtQ5kttDlyWyRRLksQRwtdUM3FlyGcIsE8Pv1Gs2N6iNA
oS1hzuFF3aFh2BxJGYFPqQZm6iYqqPqlmidFMkoUnVB3KWpM/l4uBMkcthsJDfrc
UXl6RIrVOyJU3e5HKjjllSotHe4Eghl0BP/RXvXYqMyOYyY5BqJ6fDwN0T3TtN+Y
MKGsxoUKKx1S74RTt1SbLdUQ9oRfC7eOpbhYEVF9qieaX09Ci+p0FHYTS2og4Wgr
awIoGdCBJgK/pfmpTGvipTms5ItslDv83Q3T7qlfXPrjwRddQrMCFx1poE+HpEQW
IxxqapdDRpAseqscSGLUSQeJ2drGQpZKRcaq8BiMRkh6wB3aeBbuUDExA+yUrnCd
td1QZDrmpQObWnDG6AUrBfGavEpVo8Wx/MHAYCaoiIYs8PhyDuuksKuUBkh2tyHX
pLkvPgVmLRh00r1/iBxQwap7ZWOxXP6pruq0nUId8v+ga6XULd+HxM8n5H2XU994
rlSq0vCjf32O/E9nqTCVNtuGhwsdHSFddWJe/W4lwQfG48jn0bghHx9PRsIwExLo
9IyiXXpuQ1YYrWcLY7Fezw0N/sHpzhhD9p5TnRIovo55++wpQ6D9YnSuWTqt8D3M
mHzLJrwd6BqoA4Dn/yj96ZNwK19DXP9mQs1Ul6s4s4MGFGp+hanrgsGJ0/qRmmjZ
wmbjaaCIwwGzg2cByp3MHLQyySSjSWdMXpDvjQsPV1f4buQJUWkkAGTxZm6eMAtL
NOhtQOGEMO79fO7Uke/lqHHikDLHukG+V8jJfCOGe/Ad4UyRpJQmWQuZsg7bfZ1A
Val8F13RshLPmjbV40Lrg3ZSHpNiFtQGIsB2WwGIwz669UnxUVgiA020KMcvsXlc
mSB/tjuaPTVlRd+3Bv3B7KIohVhLnPmCLO/DU1fsFzq4ZScT5mGU0X6LthEZTWCC
HapTv4VeRmdMG19Q/m/Yy52h3MzCHc+QP3wEs1L29xuaPAdP7a8m3DNP93Kt6dX/
oXgVXH1oftq8ejk+DanOcIS31NfiO/bBQOMfmQwjW9/vjsF1fcYIx3ALmbc0NBDz
hcDR9XbFmAItWK+9crCONMJGThUQ5Tyl7L/I3+zaS4qynxKvi0LspNd22budgjz9
EYNiws+4W7p0ySmNf58I5oSYnbcTTwnIfpfC8tPHGemeQs8LO+1LoPXm4fgnk/zG
8kYzmpPLA0Tr3XkrmUCPeg42ygORlqFM+QGFZy3LaD+GrahwcWDDongiCWhQHhmt
R8Gveb82pmMK1E25V+EFBSI6wyxfm1BkST8KDBN8b8Wl0WdVONrMvwQhtJ7oWIpA
ByPtBrWgi2V7yEk42VNV/x/OllKK/KAy4ahXROJ+yo7omZf3H2shmo0hGtUJyXgI
an90v+mDFJX6MspfeOGc1E2OrSsBEoR5l0sLOLnB5ZrL7AsFIslw17lTjKGP/94o
tFppCD/UlvIMxxGBffgAW4DNNbfRctMgG4FFqZ3yaj7Q1eVNqz5pI0oGlJo4Tarq
l17aVYMUGknsDlNUkhCfue1ZlfPpg8xx15AS595zhRN3lLMNroB7ZNIQP0KEjz+c
nsa2UvuBJCkzboTrhc+hg2gtgdz6Hg3Ra+t+AuNp4crjcLAd5KgAgvSbkJQEs6lf
IHUelzJldpgZdncaQbecPvNgjkYH/PKu/h65zMXD3H91DQHwYUGQ7NtBBDe+jc7K
EZCnoEW+HcLl526FKs/RwNXuQD82fq1r2SRpo/+mIFeM4kCeMGrtCxw81fUzubX8
FS9PeobpYacZhwagui4oqQGqjbLD9OBcFSSLiMvZ61TKq9xXM4vbmbvaS93DhYHE
AW6ZpO8LxpG61Y+MfSQC41a2u56xe3PE3kw8/Wi8+eTVaF3PDfGTys+RMcuzxoMv
uOizJqcZXc2nOJSgr0NmCN/Tvbf6zxxhRTH/0kNQG7ebxeyqvjKPry14S8WNptu4
d+y/OjvmC4wJ+6MBfUo+mMajdONhTpQREalkqc5fsIOefk2Ih2AEwrNcln1DDQrP
ukPHmn5jyk0QePqOTn3ojx/IZnDb67VsMhe3Fe93mj2Kj3kVkgjm/PaN5aqlicgP
G1y0koPwmhljAys0VMC+NFn2T19VFO9RG2+qm30Wt1gQkWCNVRXBve4Oh5s0VOK6
AMcTy/kgbPA+Ag2TP2jWxCVN9WA1wwotauZxMRwR7sXaeDQqRUXC7/wZsw6xPZbq
SirDE3paWsr/jDRXXsd8ryPbK3UWzl/63/OHnyLPMFMOex9lt864irOKBu/Ztesm
162WG3niSCQBtlv21R+hWSFw17hLTtEwYeE9UHbEs5ABQvfRaonErH1z+PUjmeN7
jGi/is8nVS8/O66DfizCxD+AOtJlllEiIlfVp102i51ljQaLC941jeRgLySguXgU
V0qTF+BoVzYSuS39OpBUknc2VvWVxAe4oJkoXYX4TNsm06aS4F4qIviEGhcsPSS0
eIrwc+oXp6gTYrPsvIxpTd16HXWPKalZj3m+bLUNOykmDoWrL+6NxmivtTFLnV3d
vW1oYmgkeFYeePo4GDH9RQ==
`protect END_PROTECTED
