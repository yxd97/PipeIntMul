`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3PriyrI5v4pww5JI3PV1zRgEdCvgbSjoeOUenEFAxTb8uDromJCWlQi5hALvknM7
+k3pR2YRQqJMe6RhRvfL9+gA+oywU58xnsH9Ee4QCR5Om4BHgV3f9FstV0r1JFU/
dm1UN2JJRbcvfTbmrJuWzqlg1pA+K/SCtFBGACZFDdf+YKvh+WNsWGPN+CyTwULk
gNonnCT5XQaLx0m2AbOZPyBiYv1N5DYKS6Dklf1t04bh9HnPMqfMzkv7zMqv+d2+
HqigAb9lqNF8PkkXz07h8KnqfiypyUgKOi3xLL8ttZ2cHfVQSMoygVo5oRyqI1Ux
fd/ASr0oFQY3aEkYS6ILFGY6oG/yOdUoHFFgEMEXXeKelGr6fmBLYNaEgGU5FvO1
kYCFdWHwrJxwWa097cehAULOFLntwo7AJtBiIdCpl0qgF1igb2rfP3sO/GwUcd5z
FUzlRYu59m922fYAmgT/h/UhYhFRoONMvn1LI6Ma+uY7PM/uNRQLUjEEzUXlQnaM
Q6+KBpY6ugOYupHSgmjImNWyuV3H5KPeZTx0x/2GtwunDjB3u/SSJ6muO5YopD7C
duzIXWnar+MPvXfRpU5VCbDUk7R/cmBerY+hg0acrW1Utoj+0SggFlNGGM0GUWs/
13bWglFWkKUA++9J7AhurzLjKOa3AuMkQI6FodK0koiH6hTc3ajFUYlZnNFamyyn
L11V/j1QZwSWMXdrsJi3lucNC6CDCVhCZAA2ZM8w8UawMNr9gnXvcmBRf98MQHZI
bKrHSI3beobyemgajzsY5KwO8p9+9kyKdb5R9Ulhh+b5WKWFW/hoca1qLtyqxIlC
OSyqS9MG8zc6ROFLzaniPQEZxUaQFFOAi0o2lf5/7oSq+Js95pOPj82R24CpFqbr
MEXlrAmhCSFVy0+MsUtzKPsrBsw3rlcqax76R6hlBkQbObg2m+VbXbyXNH7FTDT2
Gk8BSKx1I9k9vFBnvYur90ultRRrnU90xsdvy/2uiivZ1r/B9jlq+MLIyaB6u6v1
`protect END_PROTECTED
