library verilog;
use verilog.vl_types.all;
entity GTHE2_CHANNEL is
    generic(
        ACJTAG_DEBUG_MODE: vl_logic_vector(0 downto 0) := (others => Hi0);
        ACJTAG_MODE     : vl_logic_vector(0 downto 0) := (others => Hi0);
        ACJTAG_RESET    : vl_logic_vector(0 downto 0) := (others => Hi0);
        ADAPT_CFG0      : vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        ALIGN_COMMA_DOUBLE: string  := "FALSE";
        ALIGN_COMMA_ENABLE: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        ALIGN_COMMA_WORD: integer := 1;
        ALIGN_MCOMMA_DET: string  := "TRUE";
        ALIGN_MCOMMA_VALUE: vl_logic_vector(9 downto 0) := (Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1);
        ALIGN_PCOMMA_DET: string  := "TRUE";
        ALIGN_PCOMMA_VALUE: vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        A_RXOSCALRESET  : vl_logic_vector(0 downto 0) := (others => Hi0);
        CBCC_DATA_SOURCE_SEL: string  := "DECODED";
        CFOK_CFG        : vl_logic_vector(41 downto 0) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CFOK_CFG2       : vl_logic_vector(5 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        CFOK_CFG3       : vl_logic_vector(5 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_KEEP_ALIGN: string  := "FALSE";
        CHAN_BOND_MAX_SKEW: integer := 7;
        CHAN_BOND_SEQ_1_1: vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        CHAN_BOND_SEQ_1_2: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_3: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_4: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_1_ENABLE: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        CHAN_BOND_SEQ_2_1: vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_2: vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_3: vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_4: vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CHAN_BOND_SEQ_2_ENABLE: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        CHAN_BOND_SEQ_2_USE: string  := "FALSE";
        CHAN_BOND_SEQ_LEN: integer := 1;
        CLK_CORRECT_USE : string  := "TRUE";
        CLK_COR_KEEP_IDLE: string  := "FALSE";
        CLK_COR_MAX_LAT : integer := 20;
        CLK_COR_MIN_LAT : integer := 18;
        CLK_COR_PRECEDENCE: string  := "TRUE";
        CLK_COR_REPEAT_WAIT: integer := 0;
        CLK_COR_SEQ_1_1 : vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        CLK_COR_SEQ_1_2 : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_3 : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_4 : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_1_ENABLE: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        CLK_COR_SEQ_2_1 : vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_2 : vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_3 : vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_4 : vl_logic_vector(9 downto 0) := (Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        CLK_COR_SEQ_2_ENABLE: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        CLK_COR_SEQ_2_USE: string  := "FALSE";
        CLK_COR_SEQ_LEN : integer := 1;
        CPLL_CFG        : vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        CPLL_FBDIV      : integer := 4;
        CPLL_FBDIV_45   : integer := 5;
        CPLL_INIT_CFG   : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0);
        CPLL_LOCK_CFG   : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        CPLL_REFCLK_DIV : integer := 1;
        DEC_MCOMMA_DETECT: string  := "TRUE";
        DEC_PCOMMA_DETECT: string  := "TRUE";
        DEC_VALID_COMMA_ONLY: string  := "TRUE";
        DMONITOR_CFG    : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_CLK_PHASE_SEL: vl_logic_vector(0 downto 0) := (others => Hi0);
        ES_CONTROL      : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_ERRDET_EN    : string  := "FALSE";
        ES_EYE_SCAN_EN  : string  := "TRUE";
        ES_HORZ_OFFSET  : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_PMA_CFG      : vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_PRESCALE     : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_QUALIFIER    : vl_logic_vector(79 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_QUAL_MASK    : vl_logic_vector(79 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_SDATA_MASK   : vl_logic_vector(79 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        ES_VERT_OFFSET  : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        FTS_DESKEW_SEQ_ENABLE: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        FTS_LANE_DESKEW_CFG: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        FTS_LANE_DESKEW_EN: string  := "FALSE";
        GEARBOX_MODE    : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        LOOPBACK_CFG    : vl_logic_vector(0 downto 0) := (others => Hi0);
        OUTREFCLK_SEL_INV: vl_logic_vector(1 downto 0) := (Hi1, Hi1);
        PCS_PCIE_EN     : string  := "FALSE";
        PCS_RSVD_ATTR   : vl_logic_vector(47 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PD_TRANS_TIME_FROM_P2: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0);
        PD_TRANS_TIME_NONE_P2: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1);
        PD_TRANS_TIME_TO_P2: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        PMA_RSV         : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PMA_RSV2        : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0);
        PMA_RSV3        : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PMA_RSV4        : vl_logic_vector(14 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0);
        PMA_RSV5        : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        RESET_POWERSAVE_DISABLE: vl_logic_vector(0 downto 0) := (others => Hi0);
        RXBUFRESET_TIME : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        RXBUF_ADDR_MODE : string  := "FULL";
        RXBUF_EIDLE_HI_CNT: vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        RXBUF_EIDLE_LO_CNT: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        RXBUF_EN        : string  := "TRUE";
        RXBUF_RESET_ON_CB_CHANGE: string  := "TRUE";
        RXBUF_RESET_ON_COMMAALIGN: string  := "FALSE";
        RXBUF_RESET_ON_EIDLE: string  := "FALSE";
        RXBUF_RESET_ON_RATE_CHANGE: string  := "TRUE";
        RXBUF_THRESH_OVFLW: integer := 61;
        RXBUF_THRESH_OVRD: string  := "FALSE";
        RXBUF_THRESH_UNDFLW: integer := 4;
        RXCDRFREQRESET_TIME: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        RXCDRPHRESET_TIME: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        RXCDR_CFG       : vl_logic_vector(82 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0);
        RXCDR_FR_RESET_ON_EIDLE: vl_logic_vector(0 downto 0) := (others => Hi0);
        RXCDR_HOLD_DURING_EIDLE: vl_logic_vector(0 downto 0) := (others => Hi0);
        RXCDR_LOCK_CFG  : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        RXCDR_PH_RESET_ON_EIDLE: vl_logic_vector(0 downto 0) := (others => Hi0);
        RXDFELPMRESET_TIME: vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1);
        RXDLY_CFG       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        RXDLY_LCFG      : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        RXDLY_TAP_CFG   : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXGEARBOX_EN    : string  := "FALSE";
        RXISCANRESET_TIME: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        RXLPM_HF_CFG    : vl_logic_vector(13 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXLPM_LF_CFG    : vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXOOB_CFG       : vl_logic_vector(6 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        RXOOB_CLK_CFG   : string  := "PMA";
        RXOSCALRESET_TIME: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        RXOSCALRESET_TIMEOUT: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        RXOUT_DIV       : integer := 2;
        RXPCSRESET_TIME : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        RXPHDLY_CFG     : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        RXPH_CFG        : vl_logic_vector(23 downto 0) := (Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        RXPH_MONITOR_SEL: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        RXPI_CFG0       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RXPI_CFG1       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RXPI_CFG2       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RXPI_CFG3       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RXPI_CFG4       : vl_logic_vector(0 downto 0) := (others => Hi0);
        RXPI_CFG5       : vl_logic_vector(0 downto 0) := (others => Hi0);
        RXPI_CFG6       : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        RXPMARESET_TIME : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        RXPRBS_ERR_LOOPBACK: vl_logic_vector(0 downto 0) := (others => Hi0);
        RXSLIDE_AUTO_WAIT: integer := 7;
        RXSLIDE_MODE    : string  := "OFF";
        RXSYNC_MULTILANE: vl_logic_vector(0 downto 0) := (others => Hi0);
        RXSYNC_OVRD     : vl_logic_vector(0 downto 0) := (others => Hi0);
        RXSYNC_SKIP_DA  : vl_logic_vector(0 downto 0) := (others => Hi0);
        RX_BIAS_CFG     : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        RX_BUFFER_CFG   : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_CLK25_DIV    : integer := 7;
        RX_CLKMUX_PD    : vl_logic_vector(0 downto 0) := (others => Hi1);
        RX_CM_SEL       : vl_logic_vector(1 downto 0) := (Hi1, Hi1);
        RX_CM_TRIM      : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi0, Hi0);
        RX_DATA_WIDTH   : integer := 20;
        RX_DDI_SEL      : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DEBUG_CFG    : vl_logic_vector(13 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DEFER_RESET_BUF_EN: string  := "TRUE";
        RX_DFELPM_CFG0  : vl_logic_vector(3 downto 0) := (Hi0, Hi1, Hi1, Hi0);
        RX_DFELPM_CFG1  : vl_logic_vector(0 downto 0) := (others => Hi0);
        RX_DFELPM_KLKH_AGC_STUP_EN: vl_logic_vector(0 downto 0) := (others => Hi1);
        RX_DFE_AGC_CFG0 : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        RX_DFE_AGC_CFG1 : vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        RX_DFE_AGC_CFG2 : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi0);
        RX_DFE_AGC_OVRDEN: vl_logic_vector(0 downto 0) := (others => Hi1);
        RX_DFE_GAIN_CFG : vl_logic_vector(22 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_H2_CFG   : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_H3_CFG   : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_H4_CFG   : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_H5_CFG   : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_H6_CFG   : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_H7_CFG   : vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_KL_CFG   : vl_logic_vector(32 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_KL_LPM_KH_CFG0: vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        RX_DFE_KL_LPM_KH_CFG1: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        RX_DFE_KL_LPM_KH_CFG2: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        RX_DFE_KL_LPM_KH_OVRDEN: vl_logic_vector(0 downto 0) := (others => Hi1);
        RX_DFE_KL_LPM_KL_CFG0: vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        RX_DFE_KL_LPM_KL_CFG1: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi0);
        RX_DFE_KL_LPM_KL_CFG2: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi1, Hi0);
        RX_DFE_KL_LPM_KL_OVRDEN: vl_logic_vector(0 downto 0) := (others => Hi1);
        RX_DFE_LPM_CFG  : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_LPM_HOLD_DURING_EIDLE: vl_logic_vector(0 downto 0) := (others => Hi0);
        RX_DFE_ST_CFG   : vl_logic_vector(53 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1);
        RX_DFE_UT_CFG   : vl_logic_vector(16 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_DFE_VP_CFG   : vl_logic_vector(16 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi1, Hi1);
        RX_DISPERR_SEQ_MATCH: string  := "TRUE";
        RX_INT_DATAWIDTH: integer := 0;
        RX_OS_CFG       : vl_logic_vector(12 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        RX_SIG_VALID_DLY: integer := 10;
        RX_XCLK_SEL     : string  := "RXREC";
        SAS_MAX_COM     : integer := 64;
        SAS_MIN_COM     : integer := 36;
        SATA_BURST_SEQ_LEN: vl_logic_vector(3 downto 0) := (Hi1, Hi1, Hi1, Hi1);
        SATA_BURST_VAL  : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        SATA_CPLL_CFG   : string  := "VCO_3000MHZ";
        SATA_EIDLE_VAL  : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        SATA_MAX_BURST  : integer := 8;
        SATA_MAX_INIT   : integer := 21;
        SATA_MAX_WAKE   : integer := 7;
        SATA_MIN_BURST  : integer := 4;
        SATA_MIN_INIT   : integer := 12;
        SATA_MIN_WAKE   : integer := 4;
        SHOW_REALIGN_COMMA: string  := "TRUE";
        SIM_CPLLREFCLK_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        SIM_RECEIVER_DETECT_PASS: string  := "TRUE";
        SIM_RESET_SPEEDUP: string  := "TRUE";
        SIM_TX_EIDLE_DRIVE_LEVEL: string  := "X";
        SIM_VERSION     : string  := "1.1";
        TERM_RCAL_CFG   : vl_logic_vector(14 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        TERM_RCAL_OVRD  : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        TRANS_TIME_RATE : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        TST_RSV         : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXBUF_EN        : string  := "TRUE";
        TXBUF_RESET_ON_RATE_CHANGE: string  := "FALSE";
        TXDLY_CFG       : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1);
        TXDLY_LCFG      : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0);
        TXDLY_TAP_CFG   : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXGEARBOX_EN    : string  := "FALSE";
        TXOOB_CFG       : vl_logic_vector(0 downto 0) := (others => Hi0);
        TXOUT_DIV       : integer := 2;
        TXPCSRESET_TIME : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        TXPHDLY_CFG     : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXPH_CFG        : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXPH_MONITOR_SEL: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        TXPI_CFG0       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        TXPI_CFG1       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        TXPI_CFG2       : vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        TXPI_CFG3       : vl_logic_vector(0 downto 0) := (others => Hi0);
        TXPI_CFG4       : vl_logic_vector(0 downto 0) := (others => Hi0);
        TXPI_CFG5       : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        TXPI_GREY_SEL   : vl_logic_vector(0 downto 0) := (others => Hi0);
        TXPI_INVSTROBE_SEL: vl_logic_vector(0 downto 0) := (others => Hi0);
        TXPI_PPMCLK_SEL : string  := "TXUSRCLK2";
        TXPI_PPM_CFG    : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TXPI_SYNFREQ_PPM: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        TXPMARESET_TIME : vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi1);
        TXSYNC_MULTILANE: vl_logic_vector(0 downto 0) := (others => Hi0);
        TXSYNC_OVRD     : vl_logic_vector(0 downto 0) := (others => Hi0);
        TXSYNC_SKIP_DA  : vl_logic_vector(0 downto 0) := (others => Hi0);
        TX_CLK25_DIV    : integer := 7;
        TX_CLKMUX_PD    : vl_logic_vector(0 downto 0) := (others => Hi1);
        TX_DATA_WIDTH   : integer := 20;
        TX_DEEMPH0      : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_DEEMPH1      : vl_logic_vector(5 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_DRIVE_MODE   : string  := "DIRECT";
        TX_EIDLE_ASSERT_DELAY: vl_logic_vector(2 downto 0) := (Hi1, Hi1, Hi0);
        TX_EIDLE_DEASSERT_DELAY: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        TX_INT_DATAWIDTH: integer := 0;
        TX_LOOPBACK_DRIVE_HIZ: string  := "FALSE";
        TX_MAINCURSOR_SEL: vl_logic_vector(0 downto 0) := (others => Hi0);
        TX_MARGIN_FULL_0: vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi1, Hi1, Hi1, Hi0);
        TX_MARGIN_FULL_1: vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi1, Hi0, Hi0, Hi1);
        TX_MARGIN_FULL_2: vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1);
        TX_MARGIN_FULL_3: vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        TX_MARGIN_FULL_4: vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_MARGIN_LOW_0 : vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0);
        TX_MARGIN_LOW_1 : vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0);
        TX_MARGIN_LOW_2 : vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0);
        TX_MARGIN_LOW_3 : vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_MARGIN_LOW_4 : vl_logic_vector(6 downto 0) := (Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_QPI_STATUS_EN: vl_logic_vector(0 downto 0) := (others => Hi0);
        TX_RXDETECT_CFG : vl_logic_vector(13 downto 0) := (Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0);
        TX_RXDETECT_PRECHARGE_TIME: vl_logic_vector(16 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TX_RXDETECT_REF : vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        TX_XCLK_SEL     : string  := "TXUSR";
        UCODEER_CLR     : vl_logic_vector(0 downto 0) := (others => Hi0);
        USE_PCS_CLK_PHASE_SEL: vl_logic_vector(0 downto 0) := (others => Hi0)
    );
    port(
        CPLLFBCLKLOST   : out    vl_logic;
        CPLLLOCK        : out    vl_logic;
        CPLLREFCLKLOST  : out    vl_logic;
        DMONITOROUT     : out    vl_logic_vector(14 downto 0);
        DRPDO           : out    vl_logic_vector(15 downto 0);
        DRPRDY          : out    vl_logic;
        EYESCANDATAERROR: out    vl_logic;
        GTHTXN          : out    vl_logic;
        GTHTXP          : out    vl_logic;
        GTREFCLKMONITOR : out    vl_logic;
        PCSRSVDOUT      : out    vl_logic_vector(15 downto 0);
        PHYSTATUS       : out    vl_logic;
        RSOSINTDONE     : out    vl_logic;
        RXBUFSTATUS     : out    vl_logic_vector(2 downto 0);
        RXBYTEISALIGNED : out    vl_logic;
        RXBYTEREALIGN   : out    vl_logic;
        RXCDRLOCK       : out    vl_logic;
        RXCHANBONDSEQ   : out    vl_logic;
        RXCHANISALIGNED : out    vl_logic;
        RXCHANREALIGN   : out    vl_logic;
        RXCHARISCOMMA   : out    vl_logic_vector(7 downto 0);
        RXCHARISK       : out    vl_logic_vector(7 downto 0);
        RXCHBONDO       : out    vl_logic_vector(4 downto 0);
        RXCLKCORCNT     : out    vl_logic_vector(1 downto 0);
        RXCOMINITDET    : out    vl_logic;
        RXCOMMADET      : out    vl_logic;
        RXCOMSASDET     : out    vl_logic;
        RXCOMWAKEDET    : out    vl_logic;
        RXDATA          : out    vl_logic_vector(63 downto 0);
        RXDATAVALID     : out    vl_logic_vector(1 downto 0);
        RXDFESLIDETAPSTARTED: out    vl_logic;
        RXDFESLIDETAPSTROBEDONE: out    vl_logic;
        RXDFESLIDETAPSTROBESTARTED: out    vl_logic;
        RXDFESTADAPTDONE: out    vl_logic;
        RXDISPERR       : out    vl_logic_vector(7 downto 0);
        RXDLYSRESETDONE : out    vl_logic;
        RXELECIDLE      : out    vl_logic;
        RXHEADER        : out    vl_logic_vector(5 downto 0);
        RXHEADERVALID   : out    vl_logic_vector(1 downto 0);
        RXMONITOROUT    : out    vl_logic_vector(6 downto 0);
        RXNOTINTABLE    : out    vl_logic_vector(7 downto 0);
        RXOSINTSTARTED  : out    vl_logic;
        RXOSINTSTROBEDONE: out    vl_logic;
        RXOSINTSTROBESTARTED: out    vl_logic;
        RXOUTCLK        : out    vl_logic;
        RXOUTCLKFABRIC  : out    vl_logic;
        RXOUTCLKPCS     : out    vl_logic;
        RXPHALIGNDONE   : out    vl_logic;
        RXPHMONITOR     : out    vl_logic_vector(4 downto 0);
        RXPHSLIPMONITOR : out    vl_logic_vector(4 downto 0);
        RXPMARESETDONE  : out    vl_logic;
        RXPRBSERR       : out    vl_logic;
        RXQPISENN       : out    vl_logic;
        RXQPISENP       : out    vl_logic;
        RXRATEDONE      : out    vl_logic;
        RXRESETDONE     : out    vl_logic;
        RXSTARTOFSEQ    : out    vl_logic_vector(1 downto 0);
        RXSTATUS        : out    vl_logic_vector(2 downto 0);
        RXSYNCDONE      : out    vl_logic;
        RXSYNCOUT       : out    vl_logic;
        RXVALID         : out    vl_logic;
        TXBUFSTATUS     : out    vl_logic_vector(1 downto 0);
        TXCOMFINISH     : out    vl_logic;
        TXDLYSRESETDONE : out    vl_logic;
        TXGEARBOXREADY  : out    vl_logic;
        TXOUTCLK        : out    vl_logic;
        TXOUTCLKFABRIC  : out    vl_logic;
        TXOUTCLKPCS     : out    vl_logic;
        TXPHALIGNDONE   : out    vl_logic;
        TXPHINITDONE    : out    vl_logic;
        TXPMARESETDONE  : out    vl_logic;
        TXQPISENN       : out    vl_logic;
        TXQPISENP       : out    vl_logic;
        TXRATEDONE      : out    vl_logic;
        TXRESETDONE     : out    vl_logic;
        TXSYNCDONE      : out    vl_logic;
        TXSYNCOUT       : out    vl_logic;
        CFGRESET        : in     vl_logic;
        CLKRSVD0        : in     vl_logic;
        CLKRSVD1        : in     vl_logic;
        CPLLLOCKDETCLK  : in     vl_logic;
        CPLLLOCKEN      : in     vl_logic;
        CPLLPD          : in     vl_logic;
        CPLLREFCLKSEL   : in     vl_logic_vector(2 downto 0);
        CPLLRESET       : in     vl_logic;
        DMONFIFORESET   : in     vl_logic;
        DMONITORCLK     : in     vl_logic;
        DRPADDR         : in     vl_logic_vector(8 downto 0);
        DRPCLK          : in     vl_logic;
        DRPDI           : in     vl_logic_vector(15 downto 0);
        DRPEN           : in     vl_logic;
        DRPWE           : in     vl_logic;
        EYESCANMODE     : in     vl_logic;
        EYESCANRESET    : in     vl_logic;
        EYESCANTRIGGER  : in     vl_logic;
        GTGREFCLK       : in     vl_logic;
        GTHRXN          : in     vl_logic;
        GTHRXP          : in     vl_logic;
        GTNORTHREFCLK0  : in     vl_logic;
        GTNORTHREFCLK1  : in     vl_logic;
        GTREFCLK0       : in     vl_logic;
        GTREFCLK1       : in     vl_logic;
        GTRESETSEL      : in     vl_logic;
        GTRSVD          : in     vl_logic_vector(15 downto 0);
        GTRXRESET       : in     vl_logic;
        GTSOUTHREFCLK0  : in     vl_logic;
        GTSOUTHREFCLK1  : in     vl_logic;
        GTTXRESET       : in     vl_logic;
        LOOPBACK        : in     vl_logic_vector(2 downto 0);
        PCSRSVDIN       : in     vl_logic_vector(15 downto 0);
        PCSRSVDIN2      : in     vl_logic_vector(4 downto 0);
        PMARSVDIN       : in     vl_logic_vector(4 downto 0);
        QPLLCLK         : in     vl_logic;
        QPLLREFCLK      : in     vl_logic;
        RESETOVRD       : in     vl_logic;
        RX8B10BEN       : in     vl_logic;
        RXADAPTSELTEST  : in     vl_logic_vector(13 downto 0);
        RXBUFRESET      : in     vl_logic;
        RXCDRFREQRESET  : in     vl_logic;
        RXCDRHOLD       : in     vl_logic;
        RXCDROVRDEN     : in     vl_logic;
        RXCDRRESET      : in     vl_logic;
        RXCDRRESETRSV   : in     vl_logic;
        RXCHBONDEN      : in     vl_logic;
        RXCHBONDI       : in     vl_logic_vector(4 downto 0);
        RXCHBONDLEVEL   : in     vl_logic_vector(2 downto 0);
        RXCHBONDMASTER  : in     vl_logic;
        RXCHBONDSLAVE   : in     vl_logic;
        RXCOMMADETEN    : in     vl_logic;
        RXDDIEN         : in     vl_logic;
        RXDFEAGCHOLD    : in     vl_logic;
        RXDFEAGCOVRDEN  : in     vl_logic;
        RXDFEAGCTRL     : in     vl_logic_vector(4 downto 0);
        RXDFECM1EN      : in     vl_logic;
        RXDFELFHOLD     : in     vl_logic;
        RXDFELFOVRDEN   : in     vl_logic;
        RXDFELPMRESET   : in     vl_logic;
        RXDFESLIDETAP   : in     vl_logic_vector(4 downto 0);
        RXDFESLIDETAPADAPTEN: in     vl_logic;
        RXDFESLIDETAPHOLD: in     vl_logic;
        RXDFESLIDETAPID : in     vl_logic_vector(5 downto 0);
        RXDFESLIDETAPINITOVRDEN: in     vl_logic;
        RXDFESLIDETAPONLYADAPTEN: in     vl_logic;
        RXDFESLIDETAPOVRDEN: in     vl_logic;
        RXDFESLIDETAPSTROBE: in     vl_logic;
        RXDFETAP2HOLD   : in     vl_logic;
        RXDFETAP2OVRDEN : in     vl_logic;
        RXDFETAP3HOLD   : in     vl_logic;
        RXDFETAP3OVRDEN : in     vl_logic;
        RXDFETAP4HOLD   : in     vl_logic;
        RXDFETAP4OVRDEN : in     vl_logic;
        RXDFETAP5HOLD   : in     vl_logic;
        RXDFETAP5OVRDEN : in     vl_logic;
        RXDFETAP6HOLD   : in     vl_logic;
        RXDFETAP6OVRDEN : in     vl_logic;
        RXDFETAP7HOLD   : in     vl_logic;
        RXDFETAP7OVRDEN : in     vl_logic;
        RXDFEUTHOLD     : in     vl_logic;
        RXDFEUTOVRDEN   : in     vl_logic;
        RXDFEVPHOLD     : in     vl_logic;
        RXDFEVPOVRDEN   : in     vl_logic;
        RXDFEVSEN       : in     vl_logic;
        RXDFEXYDEN      : in     vl_logic;
        RXDLYBYPASS     : in     vl_logic;
        RXDLYEN         : in     vl_logic;
        RXDLYOVRDEN     : in     vl_logic;
        RXDLYSRESET     : in     vl_logic;
        RXELECIDLEMODE  : in     vl_logic_vector(1 downto 0);
        RXGEARBOXSLIP   : in     vl_logic;
        RXLPMEN         : in     vl_logic;
        RXLPMHFHOLD     : in     vl_logic;
        RXLPMHFOVRDEN   : in     vl_logic;
        RXLPMLFHOLD     : in     vl_logic;
        RXLPMLFKLOVRDEN : in     vl_logic;
        RXMCOMMAALIGNEN : in     vl_logic;
        RXMONITORSEL    : in     vl_logic_vector(1 downto 0);
        RXOOBRESET      : in     vl_logic;
        RXOSCALRESET    : in     vl_logic;
        RXOSHOLD        : in     vl_logic;
        RXOSINTCFG      : in     vl_logic_vector(3 downto 0);
        RXOSINTEN       : in     vl_logic;
        RXOSINTHOLD     : in     vl_logic;
        RXOSINTID0      : in     vl_logic_vector(3 downto 0);
        RXOSINTNTRLEN   : in     vl_logic;
        RXOSINTOVRDEN   : in     vl_logic;
        RXOSINTSTROBE   : in     vl_logic;
        RXOSINTTESTOVRDEN: in     vl_logic;
        RXOSOVRDEN      : in     vl_logic;
        RXOUTCLKSEL     : in     vl_logic_vector(2 downto 0);
        RXPCOMMAALIGNEN : in     vl_logic;
        RXPCSRESET      : in     vl_logic;
        RXPD            : in     vl_logic_vector(1 downto 0);
        RXPHALIGN       : in     vl_logic;
        RXPHALIGNEN     : in     vl_logic;
        RXPHDLYPD       : in     vl_logic;
        RXPHDLYRESET    : in     vl_logic;
        RXPHOVRDEN      : in     vl_logic;
        RXPMARESET      : in     vl_logic;
        RXPOLARITY      : in     vl_logic;
        RXPRBSCNTRESET  : in     vl_logic;
        RXPRBSSEL       : in     vl_logic_vector(2 downto 0);
        RXQPIEN         : in     vl_logic;
        RXRATE          : in     vl_logic_vector(2 downto 0);
        RXRATEMODE      : in     vl_logic;
        RXSLIDE         : in     vl_logic;
        RXSYNCALLIN     : in     vl_logic;
        RXSYNCIN        : in     vl_logic;
        RXSYNCMODE      : in     vl_logic;
        RXSYSCLKSEL     : in     vl_logic_vector(1 downto 0);
        RXUSERRDY       : in     vl_logic;
        RXUSRCLK        : in     vl_logic;
        RXUSRCLK2       : in     vl_logic;
        SETERRSTATUS    : in     vl_logic;
        SIGVALIDCLK     : in     vl_logic;
        TSTIN           : in     vl_logic_vector(19 downto 0);
        TX8B10BBYPASS   : in     vl_logic_vector(7 downto 0);
        TX8B10BEN       : in     vl_logic;
        TXBUFDIFFCTRL   : in     vl_logic_vector(2 downto 0);
        TXCHARDISPMODE  : in     vl_logic_vector(7 downto 0);
        TXCHARDISPVAL   : in     vl_logic_vector(7 downto 0);
        TXCHARISK       : in     vl_logic_vector(7 downto 0);
        TXCOMINIT       : in     vl_logic;
        TXCOMSAS        : in     vl_logic;
        TXCOMWAKE       : in     vl_logic;
        TXDATA          : in     vl_logic_vector(63 downto 0);
        TXDEEMPH        : in     vl_logic;
        TXDETECTRX      : in     vl_logic;
        TXDIFFCTRL      : in     vl_logic_vector(3 downto 0);
        TXDIFFPD        : in     vl_logic;
        TXDLYBYPASS     : in     vl_logic;
        TXDLYEN         : in     vl_logic;
        TXDLYHOLD       : in     vl_logic;
        TXDLYOVRDEN     : in     vl_logic;
        TXDLYSRESET     : in     vl_logic;
        TXDLYUPDOWN     : in     vl_logic;
        TXELECIDLE      : in     vl_logic;
        TXHEADER        : in     vl_logic_vector(2 downto 0);
        TXINHIBIT       : in     vl_logic;
        TXMAINCURSOR    : in     vl_logic_vector(6 downto 0);
        TXMARGIN        : in     vl_logic_vector(2 downto 0);
        TXOUTCLKSEL     : in     vl_logic_vector(2 downto 0);
        TXPCSRESET      : in     vl_logic;
        TXPD            : in     vl_logic_vector(1 downto 0);
        TXPDELECIDLEMODE: in     vl_logic;
        TXPHALIGN       : in     vl_logic;
        TXPHALIGNEN     : in     vl_logic;
        TXPHDLYPD       : in     vl_logic;
        TXPHDLYRESET    : in     vl_logic;
        TXPHDLYTSTCLK   : in     vl_logic;
        TXPHINIT        : in     vl_logic;
        TXPHOVRDEN      : in     vl_logic;
        TXPIPPMEN       : in     vl_logic;
        TXPIPPMOVRDEN   : in     vl_logic;
        TXPIPPMPD       : in     vl_logic;
        TXPIPPMSEL      : in     vl_logic;
        TXPIPPMSTEPSIZE : in     vl_logic_vector(4 downto 0);
        TXPISOPD        : in     vl_logic;
        TXPMARESET      : in     vl_logic;
        TXPOLARITY      : in     vl_logic;
        TXPOSTCURSOR    : in     vl_logic_vector(4 downto 0);
        TXPOSTCURSORINV : in     vl_logic;
        TXPRBSFORCEERR  : in     vl_logic;
        TXPRBSSEL       : in     vl_logic_vector(2 downto 0);
        TXPRECURSOR     : in     vl_logic_vector(4 downto 0);
        TXPRECURSORINV  : in     vl_logic;
        TXQPIBIASEN     : in     vl_logic;
        TXQPISTRONGPDOWN: in     vl_logic;
        TXQPIWEAKPUP    : in     vl_logic;
        TXRATE          : in     vl_logic_vector(2 downto 0);
        TXRATEMODE      : in     vl_logic;
        TXSEQUENCE      : in     vl_logic_vector(6 downto 0);
        TXSTARTSEQ      : in     vl_logic;
        TXSWING         : in     vl_logic;
        TXSYNCALLIN     : in     vl_logic;
        TXSYNCIN        : in     vl_logic;
        TXSYNCMODE      : in     vl_logic;
        TXSYSCLKSEL     : in     vl_logic_vector(1 downto 0);
        TXUSERRDY       : in     vl_logic;
        TXUSRCLK        : in     vl_logic;
        TXUSRCLK2       : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of ACJTAG_DEBUG_MODE : constant is 2;
    attribute mti_svvh_generic_type of ACJTAG_MODE : constant is 2;
    attribute mti_svvh_generic_type of ACJTAG_RESET : constant is 2;
    attribute mti_svvh_generic_type of ADAPT_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of ALIGN_COMMA_DOUBLE : constant is 1;
    attribute mti_svvh_generic_type of ALIGN_COMMA_ENABLE : constant is 2;
    attribute mti_svvh_generic_type of ALIGN_COMMA_WORD : constant is 2;
    attribute mti_svvh_generic_type of ALIGN_MCOMMA_DET : constant is 1;
    attribute mti_svvh_generic_type of ALIGN_MCOMMA_VALUE : constant is 2;
    attribute mti_svvh_generic_type of ALIGN_PCOMMA_DET : constant is 1;
    attribute mti_svvh_generic_type of ALIGN_PCOMMA_VALUE : constant is 2;
    attribute mti_svvh_generic_type of A_RXOSCALRESET : constant is 2;
    attribute mti_svvh_generic_type of CBCC_DATA_SOURCE_SEL : constant is 1;
    attribute mti_svvh_generic_type of CFOK_CFG : constant is 2;
    attribute mti_svvh_generic_type of CFOK_CFG2 : constant is 2;
    attribute mti_svvh_generic_type of CFOK_CFG3 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_KEEP_ALIGN : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_MAX_SKEW : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_1 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_2 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_3 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_4 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_1_ENABLE : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_1 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_2 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_3 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_4 : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_ENABLE : constant is 2;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_2_USE : constant is 1;
    attribute mti_svvh_generic_type of CHAN_BOND_SEQ_LEN : constant is 2;
    attribute mti_svvh_generic_type of CLK_CORRECT_USE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_KEEP_IDLE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_MAX_LAT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_MIN_LAT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_PRECEDENCE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_REPEAT_WAIT : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_1 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_2 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_3 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_4 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_1_ENABLE : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_1 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_2 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_3 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_4 : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_ENABLE : constant is 2;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_2_USE : constant is 1;
    attribute mti_svvh_generic_type of CLK_COR_SEQ_LEN : constant is 2;
    attribute mti_svvh_generic_type of CPLL_CFG : constant is 2;
    attribute mti_svvh_generic_type of CPLL_FBDIV : constant is 2;
    attribute mti_svvh_generic_type of CPLL_FBDIV_45 : constant is 2;
    attribute mti_svvh_generic_type of CPLL_INIT_CFG : constant is 2;
    attribute mti_svvh_generic_type of CPLL_LOCK_CFG : constant is 2;
    attribute mti_svvh_generic_type of CPLL_REFCLK_DIV : constant is 2;
    attribute mti_svvh_generic_type of DEC_MCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of DEC_PCOMMA_DETECT : constant is 1;
    attribute mti_svvh_generic_type of DEC_VALID_COMMA_ONLY : constant is 1;
    attribute mti_svvh_generic_type of DMONITOR_CFG : constant is 2;
    attribute mti_svvh_generic_type of ES_CLK_PHASE_SEL : constant is 2;
    attribute mti_svvh_generic_type of ES_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of ES_ERRDET_EN : constant is 1;
    attribute mti_svvh_generic_type of ES_EYE_SCAN_EN : constant is 1;
    attribute mti_svvh_generic_type of ES_HORZ_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of ES_PMA_CFG : constant is 2;
    attribute mti_svvh_generic_type of ES_PRESCALE : constant is 2;
    attribute mti_svvh_generic_type of ES_QUALIFIER : constant is 2;
    attribute mti_svvh_generic_type of ES_QUAL_MASK : constant is 2;
    attribute mti_svvh_generic_type of ES_SDATA_MASK : constant is 2;
    attribute mti_svvh_generic_type of ES_VERT_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of FTS_DESKEW_SEQ_ENABLE : constant is 2;
    attribute mti_svvh_generic_type of FTS_LANE_DESKEW_CFG : constant is 2;
    attribute mti_svvh_generic_type of FTS_LANE_DESKEW_EN : constant is 1;
    attribute mti_svvh_generic_type of GEARBOX_MODE : constant is 2;
    attribute mti_svvh_generic_type of LOOPBACK_CFG : constant is 2;
    attribute mti_svvh_generic_type of OUTREFCLK_SEL_INV : constant is 2;
    attribute mti_svvh_generic_type of PCS_PCIE_EN : constant is 1;
    attribute mti_svvh_generic_type of PCS_RSVD_ATTR : constant is 2;
    attribute mti_svvh_generic_type of PD_TRANS_TIME_FROM_P2 : constant is 2;
    attribute mti_svvh_generic_type of PD_TRANS_TIME_NONE_P2 : constant is 2;
    attribute mti_svvh_generic_type of PD_TRANS_TIME_TO_P2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_RSV : constant is 2;
    attribute mti_svvh_generic_type of PMA_RSV2 : constant is 2;
    attribute mti_svvh_generic_type of PMA_RSV3 : constant is 2;
    attribute mti_svvh_generic_type of PMA_RSV4 : constant is 2;
    attribute mti_svvh_generic_type of PMA_RSV5 : constant is 2;
    attribute mti_svvh_generic_type of RESET_POWERSAVE_DISABLE : constant is 2;
    attribute mti_svvh_generic_type of RXBUFRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXBUF_ADDR_MODE : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_EIDLE_HI_CNT : constant is 2;
    attribute mti_svvh_generic_type of RXBUF_EIDLE_LO_CNT : constant is 2;
    attribute mti_svvh_generic_type of RXBUF_EN : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_RESET_ON_CB_CHANGE : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_RESET_ON_COMMAALIGN : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_RESET_ON_EIDLE : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_RESET_ON_RATE_CHANGE : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_THRESH_OVFLW : constant is 2;
    attribute mti_svvh_generic_type of RXBUF_THRESH_OVRD : constant is 1;
    attribute mti_svvh_generic_type of RXBUF_THRESH_UNDFLW : constant is 2;
    attribute mti_svvh_generic_type of RXCDRFREQRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXCDRPHRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXCDR_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXCDR_FR_RESET_ON_EIDLE : constant is 2;
    attribute mti_svvh_generic_type of RXCDR_HOLD_DURING_EIDLE : constant is 2;
    attribute mti_svvh_generic_type of RXCDR_LOCK_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXCDR_PH_RESET_ON_EIDLE : constant is 2;
    attribute mti_svvh_generic_type of RXDFELPMRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXDLY_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXDLY_LCFG : constant is 2;
    attribute mti_svvh_generic_type of RXDLY_TAP_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXGEARBOX_EN : constant is 1;
    attribute mti_svvh_generic_type of RXISCANRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXLPM_HF_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXLPM_LF_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXOOB_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXOOB_CLK_CFG : constant is 1;
    attribute mti_svvh_generic_type of RXOSCALRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXOSCALRESET_TIMEOUT : constant is 2;
    attribute mti_svvh_generic_type of RXOUT_DIV : constant is 2;
    attribute mti_svvh_generic_type of RXPCSRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXPHDLY_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXPH_CFG : constant is 2;
    attribute mti_svvh_generic_type of RXPH_MONITOR_SEL : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG1 : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG2 : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG3 : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG4 : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG5 : constant is 2;
    attribute mti_svvh_generic_type of RXPI_CFG6 : constant is 2;
    attribute mti_svvh_generic_type of RXPMARESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of RXPRBS_ERR_LOOPBACK : constant is 2;
    attribute mti_svvh_generic_type of RXSLIDE_AUTO_WAIT : constant is 2;
    attribute mti_svvh_generic_type of RXSLIDE_MODE : constant is 1;
    attribute mti_svvh_generic_type of RXSYNC_MULTILANE : constant is 2;
    attribute mti_svvh_generic_type of RXSYNC_OVRD : constant is 2;
    attribute mti_svvh_generic_type of RXSYNC_SKIP_DA : constant is 2;
    attribute mti_svvh_generic_type of RX_BIAS_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_BUFFER_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_CLK25_DIV : constant is 2;
    attribute mti_svvh_generic_type of RX_CLKMUX_PD : constant is 2;
    attribute mti_svvh_generic_type of RX_CM_SEL : constant is 2;
    attribute mti_svvh_generic_type of RX_CM_TRIM : constant is 2;
    attribute mti_svvh_generic_type of RX_DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of RX_DDI_SEL : constant is 2;
    attribute mti_svvh_generic_type of RX_DEBUG_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DEFER_RESET_BUF_EN : constant is 1;
    attribute mti_svvh_generic_type of RX_DFELPM_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFELPM_CFG1 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFELPM_KLKH_AGC_STUP_EN : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_AGC_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_AGC_CFG1 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_AGC_CFG2 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_AGC_OVRDEN : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_GAIN_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_H2_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_H3_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_H4_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_H5_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_H6_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_H7_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KH_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KH_CFG1 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KH_CFG2 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KH_OVRDEN : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KL_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KL_CFG1 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KL_CFG2 : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_KL_LPM_KL_OVRDEN : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_LPM_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_LPM_HOLD_DURING_EIDLE : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_ST_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_UT_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DFE_VP_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_DISPERR_SEQ_MATCH : constant is 1;
    attribute mti_svvh_generic_type of RX_INT_DATAWIDTH : constant is 2;
    attribute mti_svvh_generic_type of RX_OS_CFG : constant is 2;
    attribute mti_svvh_generic_type of RX_SIG_VALID_DLY : constant is 2;
    attribute mti_svvh_generic_type of RX_XCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of SAS_MAX_COM : constant is 2;
    attribute mti_svvh_generic_type of SAS_MIN_COM : constant is 2;
    attribute mti_svvh_generic_type of SATA_BURST_SEQ_LEN : constant is 2;
    attribute mti_svvh_generic_type of SATA_BURST_VAL : constant is 2;
    attribute mti_svvh_generic_type of SATA_CPLL_CFG : constant is 1;
    attribute mti_svvh_generic_type of SATA_EIDLE_VAL : constant is 2;
    attribute mti_svvh_generic_type of SATA_MAX_BURST : constant is 2;
    attribute mti_svvh_generic_type of SATA_MAX_INIT : constant is 2;
    attribute mti_svvh_generic_type of SATA_MAX_WAKE : constant is 2;
    attribute mti_svvh_generic_type of SATA_MIN_BURST : constant is 2;
    attribute mti_svvh_generic_type of SATA_MIN_INIT : constant is 2;
    attribute mti_svvh_generic_type of SATA_MIN_WAKE : constant is 2;
    attribute mti_svvh_generic_type of SHOW_REALIGN_COMMA : constant is 1;
    attribute mti_svvh_generic_type of SIM_CPLLREFCLK_SEL : constant is 2;
    attribute mti_svvh_generic_type of SIM_RECEIVER_DETECT_PASS : constant is 1;
    attribute mti_svvh_generic_type of SIM_RESET_SPEEDUP : constant is 1;
    attribute mti_svvh_generic_type of SIM_TX_EIDLE_DRIVE_LEVEL : constant is 1;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
    attribute mti_svvh_generic_type of TERM_RCAL_CFG : constant is 2;
    attribute mti_svvh_generic_type of TERM_RCAL_OVRD : constant is 2;
    attribute mti_svvh_generic_type of TRANS_TIME_RATE : constant is 2;
    attribute mti_svvh_generic_type of TST_RSV : constant is 2;
    attribute mti_svvh_generic_type of TXBUF_EN : constant is 1;
    attribute mti_svvh_generic_type of TXBUF_RESET_ON_RATE_CHANGE : constant is 1;
    attribute mti_svvh_generic_type of TXDLY_CFG : constant is 2;
    attribute mti_svvh_generic_type of TXDLY_LCFG : constant is 2;
    attribute mti_svvh_generic_type of TXDLY_TAP_CFG : constant is 2;
    attribute mti_svvh_generic_type of TXGEARBOX_EN : constant is 1;
    attribute mti_svvh_generic_type of TXOOB_CFG : constant is 2;
    attribute mti_svvh_generic_type of TXOUT_DIV : constant is 2;
    attribute mti_svvh_generic_type of TXPCSRESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of TXPHDLY_CFG : constant is 2;
    attribute mti_svvh_generic_type of TXPH_CFG : constant is 2;
    attribute mti_svvh_generic_type of TXPH_MONITOR_SEL : constant is 2;
    attribute mti_svvh_generic_type of TXPI_CFG0 : constant is 2;
    attribute mti_svvh_generic_type of TXPI_CFG1 : constant is 2;
    attribute mti_svvh_generic_type of TXPI_CFG2 : constant is 2;
    attribute mti_svvh_generic_type of TXPI_CFG3 : constant is 2;
    attribute mti_svvh_generic_type of TXPI_CFG4 : constant is 2;
    attribute mti_svvh_generic_type of TXPI_CFG5 : constant is 2;
    attribute mti_svvh_generic_type of TXPI_GREY_SEL : constant is 2;
    attribute mti_svvh_generic_type of TXPI_INVSTROBE_SEL : constant is 2;
    attribute mti_svvh_generic_type of TXPI_PPMCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of TXPI_PPM_CFG : constant is 2;
    attribute mti_svvh_generic_type of TXPI_SYNFREQ_PPM : constant is 2;
    attribute mti_svvh_generic_type of TXPMARESET_TIME : constant is 2;
    attribute mti_svvh_generic_type of TXSYNC_MULTILANE : constant is 2;
    attribute mti_svvh_generic_type of TXSYNC_OVRD : constant is 2;
    attribute mti_svvh_generic_type of TXSYNC_SKIP_DA : constant is 2;
    attribute mti_svvh_generic_type of TX_CLK25_DIV : constant is 2;
    attribute mti_svvh_generic_type of TX_CLKMUX_PD : constant is 2;
    attribute mti_svvh_generic_type of TX_DATA_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of TX_DEEMPH0 : constant is 2;
    attribute mti_svvh_generic_type of TX_DEEMPH1 : constant is 2;
    attribute mti_svvh_generic_type of TX_DRIVE_MODE : constant is 1;
    attribute mti_svvh_generic_type of TX_EIDLE_ASSERT_DELAY : constant is 2;
    attribute mti_svvh_generic_type of TX_EIDLE_DEASSERT_DELAY : constant is 2;
    attribute mti_svvh_generic_type of TX_INT_DATAWIDTH : constant is 2;
    attribute mti_svvh_generic_type of TX_LOOPBACK_DRIVE_HIZ : constant is 1;
    attribute mti_svvh_generic_type of TX_MAINCURSOR_SEL : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_0 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_1 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_2 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_3 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_FULL_4 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_0 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_1 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_2 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_3 : constant is 2;
    attribute mti_svvh_generic_type of TX_MARGIN_LOW_4 : constant is 2;
    attribute mti_svvh_generic_type of TX_QPI_STATUS_EN : constant is 2;
    attribute mti_svvh_generic_type of TX_RXDETECT_CFG : constant is 2;
    attribute mti_svvh_generic_type of TX_RXDETECT_PRECHARGE_TIME : constant is 2;
    attribute mti_svvh_generic_type of TX_RXDETECT_REF : constant is 2;
    attribute mti_svvh_generic_type of TX_XCLK_SEL : constant is 1;
    attribute mti_svvh_generic_type of UCODEER_CLR : constant is 2;
    attribute mti_svvh_generic_type of USE_PCS_CLK_PHASE_SEL : constant is 2;
end GTHE2_CHANNEL;
