`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CkfPgzQ4YXDY4sjDbv8ZweF2l0S26gwqnkYLksLck0wkhiPgnxNqGyhSExVj2joB
xmqXhuJ80gsaIJs1Ie0k9XtZ++kPqpVPSPybu3Lg1ItvBW4/Bz0vl16JvvypUR1y
ii/CWoReEhCPEOQipaTGlwDonAXxyHChl7vap4dwQtY8o6Dt+ZmKEmNIMpqyFsat
7iaXKWC7GgRvjNcf8xQGWGP2LwGKpxu+eNSUJGmA9sHNsXP+35g0DshMRczrMRDj
jlMYcK+kdfnzw37P0ZD8zP5Umdx0UxTKK6YG1HS46mYJAs7V7wjVnbzq/YJhNd0l
neIXx24xPL3CH5ObS6wBxWxMU4h2sEzJASVgOJ9Eit7scikygEzr4eyCBlqeQHlO
Li5PrB4nyeZ8v99BTmdLVze5OjbkQpVQeCrq1nwaQBZH6eWjQdnVL0GnQHYkEv3x
MT/knFWOeGJUGXuRbywmeBpvQ2rS/K72V2XcVa5LwCZIv9Z8DHy3tyWUxywJBrS0
vW6bXGwRQ3JjEFD0AMJD0gfgZWDkODPSkGtDnwOZeP08Rg+Nz16tXgvThinpX/CR
D6BU3tODD9hRDCrf1av0dw==
`protect END_PROTECTED
