`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7N177N4FVXjwtXeBRA2kt2lo+7Zq3UwztDV0vhMSJbiaSl6YpKPy5tpmRj7Znlz9
DGQUXJru9T2+Fqbp8cZnlxU3OnZaNm1uYs/s0Yy2Grggn85RMRKMOR5b2ZXr16NG
C1X+y4i5XhfItrVC17IicxaHliRL59aNjtAFMb+Xyc6cav00XDJYmENyRwtSpO/m
HTSkiCqb1r46XRfTW6pQiRlbPcVftp/A9COXPeXEFeklVf2xi7CLzjaHkwrTEk7a
pTFcGWpuMb9+Rq/7Ewhy+guJUR5rgk2iJwWjO4wx5ave1QP8MIh72+rX2/lH7mbI
aWW8j6EgIJ3BWH9yo7/mrz5CeZN93ZUmkolQgApuBG0GzITKYu4QB60UGYHkwJbc
DjDJhb5NaKqH+DHV/864Nc0IsqDO6TlCx9lvgMMCTnBHfRmA/F5HG4CFiWiEu1fE
`protect END_PROTECTED
