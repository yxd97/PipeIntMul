`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQSjlL2XgN2+Opa7nYxKjLleMBF2HlyktFPZchvXyus8dgkrxcyWXsS4WPlFOdNP
LVoXEx5Dm8OXuhFb5owd0HxQkVBhihK7GoTzAGfiFrVOcweDFKGA0VXVVLGntZt3
xAengAGTs0UFxExj+eiJY5y0pXkbnrlVDHmN3xTppfJhR8PDO9X7nAeiJugU+3RF
TVPxtqeV8xCLJ0iVf9s+8mfMpxa8fUNS0vfXt6whFThRQxzuUCXR4r0nvTFnW/Js
X+JAQsfIv6poQrYRJ+EgRgpjTy5xekx7RyCZuRX9kDgUCHtzaHaGH4YuFzwotXbu
hTjP9fvudTNWW1jRDrB/ABwGu8xBypZ0OjOWF9Zzau5igtoXXKX0i2hjAT3aougT
g6Tod+kyQeRaKkoCAEDG3A==
`protect END_PROTECTED
