`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Skwfz6sTC55hhoU0vpBb0tvU85UsHwb9hD7jisYXp9BrUMfZod7DQ7awWuqVlAGE
5Ro0+RfohZKp5eZ0jJ/pDoHMhIdUSYwuIDo7MQ9t30B00X2lmKTt0eMOSHVxBpod
pNaxogxK/hV5oWTlLbOSNh3A7UnQnBVESeD6uKIWOQIq1W7RkQ/RgdNR6D3WdgV9
E6onuv1X3ukQrvzW94bVxfs7P4DTw4E2wqsZmzmkQX070EYAhsUaE7yYZUGRScA/
UBIgvX8RfxSj7wK0ooimr0z77Wz8pmW1Jeg+ODvblx065Q94IN5nKG4WMKs65H5F
CJhtdrLtUpaJXRM2LcjF74XSbkome3V82dA3Q1Et04eXPYusBnK/5GhPhDJN9br8
hXtLbP/vxMF7KQTJC+pjZwkh0ynR7tiwm5iajcYEN77HZJbqXCLi9XBgAoMFMaL0
eNAh6M8or/1wsfOhJN/41xNWhsYBMXgsgcD+UQ5FePK2HKVo8fxr31qozWoq+ocV
+FigxVJs/I4JE5owLJFc0Wu3EtqKYDvDNMap952nhZTkECj1Kzt41saCUiWPhENT
CfpAunFdovxxc4hws+Q2Ni5K5OamVXhwtbpQfn0tIShHzlCdkhpiblTb7fwlK0pj
ap5AxxYsF9ICNGHGAb4+/Q9jCZeDQgZS8mOMqbM5LHEqf4Noyi9MwHt3p2wTZKx/
M751q4d4+W39BSfYIhvYEsfuWG7sNlSXYUEKfvBKaUDjUXX9NGhBjVduiGuLwxXE
7LThtGMgIFBf+BigYdXrI4jG3O68uYyTyl1gchcAX73VGu0VgAcsfYdfFYbPuKcB
VawKeg9ZmGTAQ5Y3dx7YnGlpn13dlKyR5lwVwwr3Wqre0lukg+E+/rz3S01ccrCN
e9EJ6Ru4bVubgCFpNRtpteXAHfw7OBgaERAWYObA1DKI5RZ0oX+fJV5CPCrhKu0X
OTWP2f88lbzS1VWsnLigKFYokuF0MC1oiB6aLjhk8rUzQrJG5lHkWj1sC4rNp4Ea
Mv4wYF/OoJTHwL9ny2JS+WSOrAEurUUaNTiJAJ8OpbLiLGu5gZUOsEkp7WuYG0zR
qp4fj0PCkg79F+APJ50YV/70AwuSKphFDdA04jZ2mVJzDWuzIqQTq1+Kw8Q49ZKX
qD7E0q7XCLkgC7yvrZ54f5rD3gpHsBKtv/gs6+eKMNi6L/0FVD6jTTl733NBpG6z
OVCNtAQ4aqcd+vfAEZH7adW4poCL3ZRcf2V+RnxAOEEXeVy61RtHkraAHBrv0tNb
32mr+7GqOALNujA/ZxAgaWsgawZ6Yu6RoUxz0Hu4Ov6nx4ZsihDs2KWFUbXorQl+
nTqL/BmCeUDnpZo/e8Vql7xZgY+8WHKTQ005v0x8vL8l3Ycw76zE9hHX+pcFYs2z
YC8LoIzba3nhbdKvG8Vv44YT5tJ1/6pbhb4Kqe9qa1MdSh/qzu5o5/GFlg5WUcYF
X79QfJQrT5WidQ1AWq5xoga2uFvC+S/8kS/6bXCikwQzVBJXhvIi2D5w3ftp4zLF
kFs84BYd8/EsWxeTav1xoJmdKn++tXjP1vZj6mWOBl11+Zf7J2YbT7+nPuiycwwW
K+YDHEVbK6eRi/gc8EQBsX1h9HM0eKOOZ0VmEBGkvMOFoRdgMEDwUg9r25fCA2ef
GlyLaM/51kviuIXx9Htm8CHc97X20DwFGmx2+B2BUk8f1UXxRTyssOlxxfFpFXYU
a/QpjzhZV8gcNbU4oyulxkw/PsEvwbdWHxak87dnG3F2EIZul3qtAFol2M7CA+sV
SqbDLvA2UBeW13lqfaRewKw/fSBykgakIcA7ZLW+JFqRy6mt7u0V9R4VvkTmGGol
lSIsft/wWxowvPG04I3tQ878Kmvll3ikUcv0vFGTENc5WA2HbjUmS4lPoRZr12Rz
NXsCdm7XDqI6Z5HWyAClrZ1G9TgbxXOEsUisgiesDO+Sj6FDvKjLLWiUig+U+Wtj
wO2/5YbDzr6Kmbokax8fGVobc9JlQMPYbkb1WxcKyYzwLufrEf1rBZk0Cj6KNDIc
AD/K7ACSkrIhsxOzSFzsYC7UHNAuyNTi8vdbrsoVijfJ+piiRAw30x2lLRfkEhH3
ZtSV6LUPSPTta4XNKy4Fis+ZQ2x+PK3dZ5BTkH0DxYdxqaBOWrd0882Mfwz2WXEX
JKYQt2ZgGIJEl4ZWkPQJRYrv/VUxi72ojtn2rECEMbDDJRBiiRXN8RCspm6pmwXy
gB5svwFpbPOuuQCxmTKoHwTMLkzUIaWZeNvtAwLWEPl+UVeYQLaBDgK44/S5ENlD
oi7Apoa7YYW4aA/ayHqC3X1XvaRezHkq0qP3qL5IykrU+F7C6BVvlCkuZodMIgqn
9tDkVs+vzhCDhQzIApyhWpGdOhmj2e/7x4t0lCzZAIlsbp4jkUgD4Kvng6ntJkit
WgcP9/RWDBamxOHB0flcWN4xbDgiOHfVc+2ZqTfYKM9d0aoGuowXsNyB+CEWSI61
HKWcfJfr0cogrO58Gsa29RJ4Met5YxIdTLH8U0u26AcAqd1zLCnKn1Wpi1KWqZzZ
YeZpJAvps3QDDExVo9QxAoe8mD7CbVFOXj6lHdw6IEG4quzOmFMDaCztHwhcYxUw
917NgTkWWW6vZR0uv7ffTgS66p/acAWPsDLkE07mTOz37wcOEV6SbWBtUMizyShy
QRZtbUZ6TGUqWHIOl22j257G7EoL56g8CSUakwI6mncumc+Aa1t2X4yAD4ZKLmln
Qec0gCtadnQO3vAnHMKjkGWwplB+icBq40GnXBrS5q/zvY8gtPsXNH0uMoU0y3JR
7fbeCp7VI1v0jEL7UrZkCz+6ehhZOOW9p1EvB1+ybFyWG5SogmN9KpiSNxDwxJUR
Tm/w5baSDR9LPf66T1N7Kr4JAYQuN3sb1S4QGnRx5utP/tyifUMiptVD36RoQsgX
ztambgyGy57IUQEVZeT3ep4SqWn0brbPsUGIHbhveiIh0F0I4DiMTOYEsxh61wzu
9kdNG5URQQ1QSDeXhEdY6VaQtQ4qCzGJbV5+5LRo7zeWBpkZcmCznO0gvHxTOQES
lq98m9qAGivcB5dZtB8vXDnqEnluuwmQPov5hfTQ+gBDtg1DrlQnaN7q8u4/62eq
aCEB6QwbCYN9/zt1mRD3rpCRYHDjDlviBbVyJB4cG8/w6s366WGPRFOTRRbIKeJm
cTWhk5yDeVw6hJyrxLL7wXXhFskQmrHQJBTcJ5zLqMeulOmpuO/+LwhsiRblK2iu
2twGviSkPTzRWHf/MKYLiZyu8pk42aOAXytSmjsVU8tuplHgjyvDVmGmRBd4rbuY
BBx4xFBmmj2KX/WUAvKgozUhu4ZjyAr8DTETnDj4leAlAoFYc8cEjH2fx5d41e2A
Ok0UKnJWtwp3gleMr4A39255OZrfiqW/lK6ZisGlaKc375RB1M/q7F5en5PzFZ4/
2JZdFVBArwe7hJ1avrkc6PI8wznSnzRPZnZsMgtNBEvqoVPM1gn+1XH2//vbsTWC
C6G2iXgRHnyIBKvaXNf79FkzNnNbqWFkTn97QH4vVe37CebE9OF3LXt6cV+j5dLd
71weMTa6rH4zDDv7OA1TBcelJwj0ZpST46/zxlpTQs/SLT5lIw5vE+VYsbLcgP7o
1BF0CoKX4SGKmBpVg2UgyDWt29PX5m7hOOGzAea4GXPTiqB1w5xj7o5ENVWKAXdM
VSSS4PdFoOC6aTUU9D25niND0j520UUJgn23eGU1S2DzrU+6pzOpYb3J6/tc0e75
r6MUi4J9sK2mUGDhyup4u5Xm6jw+Y1wR2Gq/eSl59K26q2A3LMX9iQG6OajZx2mo
APFa58hChEtof+Za3RYspRTpkXHhAZRnvILO3u1E1a8AIsVeXHnFKydleA1YzfgY
gUVEElr/EXK8s0WisZAqU+3S+oGeZTpKJBnOTaMRD3vToin/DeoZRZanpDPoUMFb
cxKUM3eJGX5wLi2/4NmbjNybgd9WleabBhOYsQL/xr4ixmaWaRZrsV1KT2mA+s5/
vPi8rQ9Voe7yNOn8Vwme2AYYb36YXBpdsEpYCnYfcdoPNnM3IRrZXsxPmZbOKF5c
PBZjPXW0Kbfbbd/mGAnfTlSgZd2CVY84wq7gfOrYEBQKDEbymWr3XOYOcT8UsfTU
XdWUuAcvgq6+MRqwLthoppCOcMTxhLS6qdRDOZgnDKnd+xHv3vIJ4ZrvJP58PEcs
mvvxmF3IEvegzrmgGX3bFd+8PVJg8Kxo9GwCy8mDwpoNaq6yNLzNt9SFPP46BpgW
Z9lVJFpx177RWnmZqxstNM2MkIwEESRsnTaAyuB7xzXcQzzFUFXXDgNB8+O3O4jy
D3YTSwPRjGlYFgYlXLw7OhLsLv52a19+TYYOlPirJ4uL+QeKGfr7hev1MaHrtw1O
zaVIEYkDEIGoI+MQ2I682qTQWyqcAan8gJVo+nA4igVe5lAMoEF7e6JPxOSYp/UA
ADvIfdZLs5oMnZUM7ixKOFAoQva8+4pt5VKQmlUbIIpA4ZAcjbTC/Les3Nzqx7n8
tK6jazgF0bhVpvp1FrlsyflNL3VWL9z16/VkGwsU3hF++Ncv9ZRCn2T74Kk85puI
3A9pTA8/D8xg8J/q+J7QhupLIGAkcP8MG2PzzP40TH8jQN9drJ2miiY8eu45Un8/
avYDb6Cl5+yeyh+xHDuiQO1L3o9ruzEMPrx6ZC0S+oQmUq5WdXnfUujkq+MVrgCW
rELb5C/x8mkpo2UadFgG2GnX++bQC6m+w2x4coHzN7oBUX3w/n+JfxaZ8q+tV+BD
gvTJrgiLjqTL5ORWPJhoVwK8GQKPOgr4acUfgGGAaE8dcR3zQFY4xJrgaWU0BG9O
0nARgInIUzPbf/TQ0IUnbclM+zC9SEpd3yh/a6s89kzO+QPouRGE6Ha5lwKaxRi4
aHAaWiJe88xEbTzyrzyIoqTqb7UvN25nher72wR2UebtYKoHE3562o7S5/mVsiPk
7vuYsKLuUJUK7M0B4mSB4X16DHRJDdI3kvFI1V5MRUoKTIAqDHcDU/kFv+B6GfYh
NOsQi9k4qSvuhf0zH8bSunWWHl6nZ4xYLLY6ezpx1jbQB88SWHKWiakwKu6oEvvL
CP4skKMts/VqP3/QgoFvVqIuNPyLagnukj9xPhG08Jo1GCQcrGa+KngVJngRl/uu
jKgPuW2nDnp/EpYiNgWexliFBvvtrRzsBUfCiVbGHRDLmyGowN0u+ZctC96V40bi
ld7pXnbgVIs/LTVx9TJHJ0DUMGjxO1gtGmghng+MnfxfyFfT6Gc+Riyh3JdeG9/P
XTqKvtAQXbMXUnncP+DtBB0op2WwdBJHjlZw9Js07TE45dnPOoW/k3oHr0nPwwRn
IfSKh+YUFuSFHze888VakYko58H3gtydAxJnujWmzU5xDzTHjPD+RPuQPQI+s2CL
edIdxsYN27PbwmHFIEb8xsP2RAFJ0LHC2iUj9FMyt+r/0TUcNJG1dviCiKoGh0Md
v9W+FT6mPFkcXyGTWH5Gk92FvPFwPvFzsBjDb3SV2Ax3NM8G8V+J5+gWxFGvz0n1
jy1cxqislakT536o7CPz6HI5DDfXfHijUP6Qy9MgFmunvwl+kP8mOrs8tU0TlXOF
7dmtPkWtTS8sv3BHkcPAuCqdEmGOdRIV1IVuRJVnGSRSKez6ufSnLu5/khaXnTfh
gnV5Hh53Hv9XfoGwHkXYzd0jqoyDIKyfaGdV700piMIXNDcg1h/wZ1midFGk15B/
b7JFiFOUUISDGvY2bLBSPpDaEQLNbCeXJg/s/vJcy9T5ko0/EYzpeOq2N6RvqMs6
sZZ4cZMz8RNvNuIIDRQo5ssUctFM4jN8Ml0g9Yts0rYSJCvIHFghOpFthLF34d5C
nWXJw7sjBbhoP2LkvcioTTpwKizyWD2A3DXj8o2SIv6LJGCX+nJ3fFWSbQlnbBMe
j+37I0aeABBb9q/aaIgPgcX1SFPLgVrCJ0Fqn/q6hczjOSx1EQrf+XffDejiMTCC
5N5gA6qtHfbO9rGa4d74jK6wls7w9l8ICYJ7tdDJ3vbxiQrAp/GHmFSj3ppT2RQx
OP3G9XeXGa4bHCJAyCS0oj8HCdOGgx4p/jeForvyVRPmno1ZyfP+d4bCOfh47jWp
eH7A/4O4homl7zer2hqXmEjh2byiiryrQTXwkWLnmwpw4+azrdw0qAMrWDawinun
eKmA9TXJcPGKpwWWNKJc/Torhk8VVRMF9zMmGXn3XX2uxOWjAppjHk92Sid/zcUE
E6iLCyUxr0f4I4QYQKTcgAh06r7s4MrHvKpejdGUyD07N9cBewn/yZw6Zs1S+4ke
EaUFJ9WNHUm7oXDowABJcCjeU7/5HLqJ+OT9SVgqe6EJtzYPzdHSJZzKUCSL5pOP
Zyzml8EEoaogcNDknisOxYxREZN/KV/shkyJpDbzH/JnDl915kU/nPlIErf9lgpA
+7/Y4aPJYF45Y2QxdvqhvI3/z+Cqds3K2XwLW4Z+WCxvvWibJqB4rrfnwfJStmqU
7c1hgk/lJFPzLjNXWhpGeo52Dm4IGB9VavolK21KkDM9dfhvdi9ue4GTSa+oTkzb
dP9Q4LSGU1jhHQOCUOthBI9W10m+KuPzFDiD9azzwVCP8Vhq/WvMUquDUWJf9BrI
bkqBiMzJENC0Vi93cQY8V/RQDA/UPhwLE9xnwg1AaPcMrYLiV2AXZPeNEJFHFnb0
vu7Pi91tWh+F8A+gRwSLPk/T5BUpq35N6txERjcqCgbxpHPGxR7vS21SNFrSt+C2
mTrav1IyKubORKmW+0tx/vyZRgn1nXmeHHSftBXOTJ00aGI/x4FtK4NGEb1aGsJw
UaG+I28qX+MlGu0jU9ifNpbsjAj+WDzIPXIZ8thGgoYs5WFTkTPzX76FioUPISUs
6svXYu/Wxw+5tkopp/uE0q+qIfbvLzsdzAdKCRADnLMQlmXNbmEklVqWDBfapw/y
6bZR/dnSQOZ5h/8Rj1tWjLQUYwkw2mIHnt+tHcAAMQFMwr1ZsTJn/JKW/zQ6TTjl
7Y0cQfqQp8U/CvbU1HpESR565cjZ1GqlQcmT/3BFeFSYYiV7U8fAVivfdYC7NJea
qv1Kk4I3MuDqcW9448KaFLvkrLY2eMlV6PniGZiypAXYlgAX34k0kmoEhC2Ox7yX
gj+2xqhxlYy/miHbnzqOJb/svSZZkMKs8vXUjW5pQvyt1TdiLZ5UA8tOOVV4xHhh
3IZWiLK8O++3FcJ8ti8tO4JltMPepdzgqwFfT8jq0ryCLhKDket2vHV5t6k9FCFV
c8js2Q1JKne5s+7G9u+iKoQs5LFVVVBlqX0nYW1+8AQ6xb7T8xVcvK+NBlIYaWnz
Ecivblyl41zCnE0IjL/zpy1T8m6J8P4+xIChlAqPxfutVLaUKTv/r2K/oQIJZStU
T23rY8nzzDjJsLdJT09GUCyYBR1MhEl62BMKI81Uar9/PTe9jmxfYQwMl/GWs8oZ
MhggLjH+qqGjocz73xahdV3Zgcr7tAlqAnDraWJrx3lp8Q96nS5jSbJDry5eHi0a
qGX2Oc/+e/R53Mbz1+NAONTyCLq8DZoFn2N9nwPCqgCxePtV78ez1UKEZPUZIkVx
Fiiuhe8Xj5hNEEuXfoBY0MdzaiNjKdeTBbLedG4bVuxzwj3xmF7l0Bv23uu8i8Qw
vjg7BFs9mkTrteB9rpmKdHp5eMw2lZoj0Y2g8SHEQ0LAl0ALuyVSCwk0rySdv+OM
5OXqB5aEYZIxBJqeB8Qv+PG9pz4KMHU1lGzMd0jm1/vX6qBM33vIw3ZUM0PU1V6L
dz0Ix/0lN5uYPOTB2c9vkGa7dG5dtM1ZGMqvZIXNmqK99jYIK50SKW1J2DFeQoCx
hvwAQNLL3D2zeu6LUYH/hPm7ofRVQrQIy9XKPO1hEiKRw1Ni0mJ+Afuo9TSf7EWI
gDgC6sj+h+69B4twlx8mP9cDTZko3jBFRXSkR4F0Z+QZY+tU6Nadv3N5P1Kbddht
1hsTBHM/gSCYNZQFgUyCZHDDssJ2BkeWZ5dFee/7AiawTLe2TJeZQS68YtmYTMUO
Qk7NYRvg8fo6QKWsz8yTEmx3dPX/m56Gc7+cS74rGx1rRqvph0cTdzEuq+N4V35h
VM52gbr4NqXwJiibqnQM4ZdPf6bmAXaVeXlkzdleXoKlMtWXlRKxUu0wMQoAjyQ6
oP0qZKyanLS8O3XfJgTuF9ILi9BFfi14IzZuvG+nwZwlFs17o+AKsigH1mJU+rp8
1Fx0rkXjlGFGAwDT2ANPl5UCXbtD+6OZunqm6fs5NSiG3dts8WWlKm/5azUTKR9i
kHZosxnl82dwiDfQPHbFH1298ODaEl0rNWUG1aO6/3ep6uPF9um85EiQOcMI0OrR
JogHSXMoDaJRo+A2YM+hoUWGGQqOk4xQttt2Yy9BaH+lvfBjhEhN3IvRe7S5BIIR
2hA+5z59p+SsdHLneDev3zvaV+O63Zfo4RyMBhHClGtXPlGvSzxvYgvZYxn5Xhc6
YK8EGmmUMVmokBcn3t0yF7xlRdwLr/ZYBMr37ar6GO6ReoTZg/HaYQ8V7jAiV0Cd
5I78ZH8AfEK0HTpDt4STeMHQ/1ZKrDS20nacld+3+bFDfYSEQGCTIOWAkX8jrd9y
5ZujsMs8NZonKzZgYADZSOeEgb0ezufANysjRBQOjCPu4L1+9bJTB85x7EtHpjWv
W6YMfCODbpDZqKgGo+d22mJQ30hKMqZqXSeXvNO0rbqIwfwojHHyI6lsv8JMsPUb
UkbGydDw70GWx3gE7TC9fODrCPlBRQptI2HriAAhBot5SB2yT+dyRMtJYJK2GRul
9WlS2Sq2HxobTOVipt8B0GgtHzEl2v8aczJ6LxC40u1gXeZtChoCF2BTO7D2gjTd
MFH5VxrR83kg9cCSRvcR6SM+ChG+zpkO+IRXH1TMJacT5t+t/iFJQqOGOKRr+5TR
sMmeZ63wyxBni/bZw8fLdtIklP/BeY2pLDPqL34vJzhZQBDEDz7RYUsNVBzI2s5T
lpmc+n6r0p4XH4jXov9vkP5cleS09WYi9/rK+Tb3dKgdFaE9ibhxblrPYx0pPR8C
FKDKea0DxIZUQShiTKhPM/Cb4AH5kVbvW/ZiCJoE25Xumzvf2RTnwqpVwmQpVGKw
VTgLGYd5WM2MsGLuJcBzjpKthoKWzsCC/wOMvBJI1TZbGouB5LbUVHJnzSeyocVv
QABqd2jAG+EArY8KR+ggyxSqX7Jop5x+Oz+U+SSYe0RihJJoeNNVnIP6O8jDbKiE
h/7gg98trbMA0+YkFyVqHfhtelS/xMsQm0aNK1bL7rKN5JpKcGvzATlxYe3zm8FS
P6U3JAMS3GIB4PT986v+Ubc6QjpfNLHFLQRvGiU01zxwmyqX6v/IjmCPVZHOZh8C
kQxrbcFiBzcwdtbeOsI9R48XbQydxcr8w2HsmrdZTO+V8jSZvRj491MwOq6P5aYL
yqJWbfdjx+0DEtcoCYD4NGFAU001bjFYxs3JN4JoiNg8l5LbQAj0JvcKUMjWyQzH
Ccb1vcBwS6fHVgieyb45CNp60rX+yu20xklfuDFcHOwVxMNP2yD5Am+gf14u03Tf
zqw+vrfJbcOcHRNxH611ByO+5HOxHrjE9JFrWfhItjW5plJKjhichi41Cy7EK59J
Z9CqcEsZ8Vui0BBlAMiaDyaABEBLXQV3mjg/tY3iwOheva+z457cXtWqGtCEwNbG
8NpB1e+3mt2xfyMcM6jDxUcBoUDkqePbcZBP3OFgubyftFUmIa/jj0u1L2kffFR4
92Cj+/kuwmqJW9/xtmzYoraxq9ujCGdaKEdDZ0XjEb003fr9oYJerY6nqOx3hSKl
OVlqqX/+LDkEWZgfRJ2Hmmb87UzsJMMRyD74lV9y5KlFJp9A1roxrERu9nUP9KjX
XQqg+3tfr6fBpaQt6Jo12a6GjDXPK0ZFNWhVul5nxrTNrXUTmC3ludBK2J/786h9
P/AFejXlCFcJzZ5RtEQsKV8j5o19NEs4AfYfqoEa0bed7RcTxt+3qIBF4ZWqh4VN
UfRlOjhifRxueVkb+/xK364CDazdMwQ7Ju5pSc5DFBMoEFBLwpB1AaSqzwDUJLXU
9NpV9O1yNrJHPdURieFn3NfFw3VmLtiwghL/AkniNd2F45u9CKCk2MIVSotHYaAU
A8klRdSnHUXMqqVMpGUymi5c1r04pqgVSlGiHYG10dJqJiTga94m9Pfm7MnQFv8x
K47yT7EHpB24MlImZP6y7utfcypZogGsmlLGCVpNl1SkOCla56IVwCQ1dlvmt9n2
0VBD5TwLa1rxJ+K8MbVK0uo/r23WxSy5yJSiiQtfOzWcj8lZaFhQojNqnDuwwHBI
mfg52Eyg/KqSWVXLW0CO50kIuiz0cFn7iPLQoMXTLo6m0DjsPB8BAarEmLKC80AV
P6CWD4seLizA47AOH6+vKUR+i0Neq9T52IOA5R8jYUX2m/vDmc2NGQ9KaKvbHU5v
l0/iVfp7ykdCvT3A1vcnPHwLCANx6nLgqJAjM9+OBG82FrqaVbRRiTtkgodvjVmE
f70GgWThlpXxg1e/gmzqk1sKN0halmY632S7SEACZkr+4AS5dGVE3XCvyG6Z4Nyn
LeAzq9UJH5E5I0AraoMNfjTxy2WhLUtW5aiKolTZJNS5i/y2xymDxIHx03Z+sJIL
YknYyNm8DMadv7Xwnu/Lq7bZF+siDDaBwgNDiIm/yrNFoBa7Mx+mtkNU3pjAtn8N
fmGcKiXucmTFHvxws8FbFkEJDdaIH08sdbWCCfhlfPy5SA+BJgNJT1/FHGmkULYX
Ta1PPrAitCow8SmCf7oxRBDs79X8cKwtnLk8H3T8ClM+HmztA8h1sMisbRRNnLax
wy3K903SoUxJtVcd6PpVE/rh0b/P3X3OmCd4agzANZhvcpyXrYfKhO2dXE+W0y9W
dUVXS5ZiV5JXMplmI+ZP+7o0N+2yuyckEFrVh7LdPT0FKHkul1EZt7qUwho1nwU4
NNoiLzvV01tRYvt0HqGIWDRve/QFigbKyqDoigXku3hC9OhYz8v4HVzKLtb7eCck
+C6NvcXzmgWfXpFQg9ixM0q01uNwDzVEQqzHlubVwB7YO7bgSIK89loYoIqeWBJn
YKG5Ez1ef+xbk80EBBQNhhGt6T0bCOT8zYmqhaL3O7ZZvbWA7AVEspbuj5trCW2q
e4Oump4xZeXCKofmcYG6a89kIH6nuIa8PUoIxkjQ+wnZQfPtSP+hTX84FS9fOoEJ
WGwVo8cnUToPl4OyNcDmZwC1oV6HxllnG+A2V53PhzbKgqBGldBKbL8Oz9kfPafY
OJtztA10dRNUcTUfaP2kxW45NnWIinBJjHgXTg0tuCm99sBio97l6aAimvDXfztk
va+4oyUaDCY+pHSrg+IyzuncYWaWnTx7qIFhk3sKauL7DzQx7a5xU3xLZ3vKl9Hl
w8xskILC3sx44QbjqVqWR4Gc0RilJxAeoeLpRSTkkVEHJv8TePPj7V06ShQb4Vul
ObWT9kD7d5eSPeswB3z6QJp5ueHC6KlqX9SeEwq0yWhw3AKUlj1Lyu5WgpH7ShWQ
eSWvQFbHd3VvBWjf0GGp3kUWEoxv6WsJmBQFUYLi1cSA6HL/VJebjrrq2mB/u8Lk
269gGEuwM9NxV+HEgdhMJfX1ATSDHlubuXeRl7LT20mtttmhnLdjq7c4poSwkQIt
N5gnMD7n9ZmgU9y7LikvVqoj8Au9zSsEAqugUxwKFdLVo8THKA/kXkZiIuW0jI8a
/vvXtfn2ObU3aoQ9iKoyFH/YO8eU9r0xqGvGbzGroAziE8dPN2e6NlWAsv7xv2Z/
b1n4ZXrzvtzBW9LAO3M4OHShBrbB72GxYlIQYnzlt6nAnN+N4RBc1MKo954JJ5ZR
+sSxsaZ7cW3Z4Ar/bxuLqOSyLESHpKilkEc3+zq9/12eLxgWG/OnTOEktDCKtqcl
VuN7nLcNuEHX5QUU6bSZys3XmTe7CLPKxqX+lF649D90fCqpCcTF3DjYHGa78YGI
JENGOUvVywLwasdeBuIVPkiU/Ibmlxm2uWEeILUKZ7bHbVZmWLOdep8u7vBEp00H
CWnuN+KKIDBZXn4X7SYfGwn+xPwt6OJ0VOxvtTsdO3hRCXNdbjUwaK2EQBOCoKkG
HDN0Gw6jraqEoP4ZIMrenHJpRYrhI2fWWNhhqcee6HbXpT44gu2Qc0XDGas3GTAa
Z9pcRuZe7gXbJv3Pn79ETuufnHcNZ9VPvhIBIVgEVkvak0REDs8a3lz+KE09MQ5K
oDSWx4ZjW0C/FhPW9simQnGdwdrWCojnFB2/SQRn1ORv3eGo4gP66PoIuNfu4Sa0
B05Qrgi04h+hGtU2L10MOxeLlNVPqzehKOMx6tLHuM0UBdGHlWTeh5+0h+gY87ln
0kBaXVl9KHReYj7RGQvw04ZiieEeJlCbHR+U1K9jdNp1r+tv2Qh6ftZ9OU079FRt
LMto9BXUwyhqLRCUscUFY1oLAbBnWCUhTRpgaJ+kif6AWFCzbisBY+0Ef2KRAgqB
1Wg/cKA0MUIayTzbMM0wiAPjcvnpNap4FSryyN9CfxsbM8q5lEQ4GOix0+98ODaX
+kGlObenodHOlAIZaC8FfPIrI3ZEI9bYABeFUIuhHsjylWVbOx1Mxa/My6HxxCCk
PltihrRoasyFRGmsyUbBjaWbXyQJ7lzc4sEpP0tcMoUuPOd9JO7n2SZkOPWocn/G
qyRFtwln9T9bxZbHxJHcvQ==
`protect END_PROTECTED
