`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Oohr8suyG4hiowV1snSlnSVv82QybN2lPKARxYlg7t3DDfshVyr0VBV2EFAxzDT
KjDc2ZmXJWYgfh6IgHyQTtEmXM1h33t3TtARqDvR+jeKvW2sXYTdqTa2u2+9NhTh
QQYT+wGwLxOXaNUa25M4HomP5goVAeyq+cFJl62HqMvBXnHU9XSN6V4yAsayJ/9h
oVYQis6mR6PJzGY4GzhEdozc6MS1MrfN0vrPPr+ob5Uc0y6ihOJuWzymJyA+bt46
31hdq6PMrXtUEijkRJixFw==
`protect END_PROTECTED
