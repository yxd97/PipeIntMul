`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
waOWileESThldM5MkZuv45aEeBhwlrOPhpkfdHwTF9QHh10VDTPfkSPRxkwQpFnm
j5ZyvKiK++xH4h2rS8CDSghI+bMHa6hTpTKzofhqHa3z53DNZO9HxBrjak9dGHTv
RdfxAxYvVALu55nyll9ZhmvyGz0gRzzBsYitoxSe18TE6CgfxJ2kBGyw5gc8EjZF
oe2BtTKSKVZlcubt2yc6Sam54L5itTUMjWjZHs6W2RpDkm+V4dY/JmkCKkOJzav1
M/4Fh8FS2Y3onC4L+EO/fyQ29SXxoC49FravxbzuPs/GfVDKqk5TmSXBeD3Umb9U
oxolj8i7p3KZyP05WBxSXQ==
`protect END_PROTECTED
