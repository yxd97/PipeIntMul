`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/CEb9pBefBS0AApEM1NgB/SNzR0Dv9P4AJTlVDgZTEuBLygGXonaYxxF9K+LS/zp
mPci5LYf6Q54p7O+7b9TYq25F7tUPpiA8WUZdG5w3BQOEedhtzZdUJQZf2s0SVCC
GDiws2pVEp+knaXf5fcQQ5A93YAdH+eXJCTEXM0bZwXGeKzfeA6ERri9rbVdjLl7
2gSaI9e0DK60vi3nYUaGV0W9U+ElSxGiuxCpxLOhUJ330UdsL4kcDX1rDTXa/RVE
sD9kPi5YZlxogZomP907cp1ttebygnn0dNIZ5WqKpdjy03rW5NT24BryC4YUn5yS
b9EJSUSnL9e58hDj0KSYgmUDO54ZTmmjo4FnwzRkNe8OYdsj1DELGKdld34f25kB
crRjjYoDwUJAZi5S1L86n56p0Kbb1j+FgsbOgFQGoJlxxT10TsLRqSoEwGftwBcd
xGWo9wZKIGjiXcclziAvk3+RMFkUyDITr2vBAkHYY/xLoqDHFKD9m6rk6qZvIgww
dMdp/BjoLVbyPaNjGTmEdqdX8gOTQMw9M9bH+9imesOsffS1oKBUyXYBY0neM5l7
1T/Nz7mngZIi+o+OQHWXGdiKbvVB5UYVVL1sYhxtaelTObuhooBQ5svj61OpKpn1
HQTC1mdVDmanfFhyJ7BWxzbVxYqbDPJHJ3w5j5ZioW15fg8Xm427iYV8ND6egn9e
GGMR69DSHStTpDOaHjPco9N0ccKXMuolldYV+lsbIF8UFPApP8Pv1ag2pthFkyp2
IEN3N7yt5be6fhilo3E21mcOBcS2vuveeCx1NQyrJRbPmMSX1VHesTLqjHPaTNE0
FguiTmN484KFJTcJvhUdqtiZ2JGZ9AeIxXH+LJSigKYRrPwFsxtGmqdZ8hsgWTrZ
24r5aF+gSoYcc1kmtHhdwQu7wbnXo84g4Xn7ebzCpLSZzDS58PGKrWO3PwET1Q4B
O56y4RDtAhfubErSiv30YyD6WKEHOxQSIg6Tl/f+icGr2kOnlVKpn53t0SGcW3YS
U8WLd5+llGNeO760pRLiscgv2u57uX4v8nEWehL8BB6UYIlVVSFGaRcnaYEFF7ML
rytF0/jwce23mCNJR1mBg3PbtMy091o8u4xdWuAsGTncTn5h9c6Uy+AJ8xUXrLAJ
iCm1z8yUhI0lMsCEvJnZqPuqCY2kwitPAOb3kBpXRifJH7cqpoF93lAqmIiN2hTr
3ys3NExqGZFv+TnwluKOMxmC4AJ3KdRpKmdIo+7ibqYksdk9WOJQU7kx08mluFaF
lSzK3LUxvEh27tDUaP3UOo76uIAlQsbufUU+bSu/WkPEzAuR/exB2QDapcT0c5ig
LS/KwZaCSKc6Nik/DAziqaDs4Kv/jT4O3+jvw2nOCRKeZdmP33RQnDerbDtoCSi7
7MByS5AGWQeFx+UZtYl9lWkBajq10wlpaC3EEtLm7Jy5pzZVPwUSN6g0Iktv4muR
vmQijspdAGpNCUCUkdVCvhDatVwwWL8k6HaOSCAsKprTv/w+yjLsHdAgudQFFe9o
U2uQF/KUXuZv5qR19EP+LD2EDjHQi4GTUjFAx6Pcaokv2w4lwD2rW/Q5ow0POU6D
AxPdgBabMGCWAYgQ5OQR7QDz4sPuyfJXXQ6vJopqNjIOgWOaYw7JTDpelZgXgVXF
rCHeblAl3WvJ5EDtrNl+R1Q/QNkR0czI8D64wbRnc00z4hDyLhSNwgGJk1s+8uaE
vvStuQP5bsvZLoxCWAkzVZ2WT6dbcrvHEo9K8d21K7ECgJnNbsKO0tniBLZFEisz
RZiaPFA/gd2IW0xborr4hJCxMtiXLEnbCGbTtfb5HSVLFxpsVqnkzvLXo4mXtS6z
jO812SSUUjDmoiMH9zwfNBGX0tMwxcogcY9l0g91hmoiKC5saMNLNfQSqpNJEbOV
JLyYGgxt/tWtXqMaVoEkc/4zoatbpLg4ddkM0luETqixBo3Dcux5IFKceyxwi2LI
aH0EYzxjjhyLOsj3I/XbaHKRrM00wnsX8I1ZHteK4VB7cOmNwItSnwYrvWgSdNNa
8zlNkHejuqmpqCEUJhq/DwhOUzcmUN6ijl+k7AHoAFpmW/MC2R1349HPN+MzxcY4
CpKUD0z3S1UIzCrBF3cvb6FHk1DMQwEUacUGwBxKP2I4sWBKEPMbtHwCIlDPXxk+
6dPrJ9gFjQlh552hGIYmC+3Kw8q2EJ1x/yaPcsvyy7jhMxu3FOxfE/k9NzxgF/kR
uHaC1wB4WoftDG8PJOquOxTY6gZ4lBZ7o+QIR8EAx7Qh2MhT/w5VGQa506B6CzfT
Cb+tQuSYUEmb0X6409qpFAbv2i6qC8JFXHBdmSxwKRQqZV/7khuaHPzbuPfDD3Gc
XiErxpFjy3K49ZzXZFrtMn+ANheFdpENv9bSEHlnitntRCL7wML+ON1kec1wLDTG
SCyyuxw1eY6aopjDE6k0Tu2kBbXImJTOhQHBaD3gJAt8lOl9uTZHIUHv+PNy35HZ
OLceMeIxxtaxHclSFvKf78QcNXgZ2lF7GsQMCEgRjJnLdAunj734+/6YYOpLpY1t
XxbrpzvMRZdctmJvgN+M+N6E1sOpl5hR3jSk50R+u9/ip/ZXgegUsX30XGEY2732
G9RKSzWPqEb5hql5ZnXfNXtFcf7EL7Y7qxTQk6SQgcT/B7hUL+7kMlemvZR6EmUl
IAsalDS2lpIiovOjPksYo1MtrSqS2DiSK8ZOUUh7Vat8Pt2Puy2ECOVgNX8SzF1S
AeyYGofy6133g3zG9Mr/41vBjSzpqetv6c7Et613BcUzjh5PnFscA7Y8X31Gb6US
bU0Ggw5pcEryeuu0TWP6J9K9sRNysGSCBN8q9P4szirsLz7wYRDA3nvOVkHeGs8L
NgntuEY5LLZBMcvYrnKy4sOd/OgKRwfjadRjIrWVuXqGYOUUvQ/+eFxAlGkoJwTc
P+9YuBRVMuURiUuNjzwMC1JGtKESljoTycAJOK1KNh/sAScWmoRizmHdsOPOGzs1
ywvn+ymIvcj2KYh69BVlPBJMM5eEGnQ0jIEps4oCFv4E/o2Tu0lQpkhqJcixfOn/
Mru3/HT+0JvsVyC3W4iUbclJnArxZ892+GNl9ThBtWgthiqWL+XxFLZykTTcL+NZ
y0ssdfufp/qegnG57jYWra2CfSngwh+7nEFFBJh7Kg0fVoV9BiiGT9Gdy8dl+Tjo
uDpbrHQF7V+usQdqkcUnOfD5fOQRnTkHFWFlTgVAKgPmSXk4MGPT6c2mwadY2xft
P96CRslHUHQf4Gh/GbETZBprSfGSx3EgjDi2wyT+v4agzd5KzgMhKamJKU4FzpWd
2c3DcE8c0Gnf88FaAgE1JBXGduXfGjBmFb7B/uxRAr6OxgUCGgaTM92OEX/MnKhy
KW8B/sChJ+uHy3HZ4OexVqrU/n1idjY3vRtuH2Lu5fiem+jp7UibQquGpRjWDBUV
Ik8MxHOcyGzxAdhtdo3hcgH6EtMSYabbO8SmNtiq3uwI4IWLjG+8UkSeILHcwPQs
PHK97xnEUY7+DU4abDzhLTx3DIYPX6ZihXNzEgbST+D8bDTDw41mxRQP6lkOFDCw
6se1WZiDA8wppt2Iteh8d1vjfYW1Ha+sl8zD24zCYjT9WZ3M10TJA4sqSlx8Y0T0
AVE/YzAPpPQaiqIrQ7C4Obevibp0EBlfm/WtwiKGizqdUQikkmlxiWGfsgQsYatX
sn7nE4tPcLMGgQ+FHHlbmFdzp4SzoOlhutHwTvNzcqEclKTMwAFmQWKRJ/ftuZXm
hZ+WxMnUgvLjPK90EBd4VyN/cRBP5ys/WMtBIkrSU0O6ksTVykOH5oUWy4PYeNGb
fbpgmTIvyArm+Y7hqf7RmHeqnyICUMxbPdz5o5ORf9YV7PbVtFACR545M1i8YSwG
ZsYfMNUQF51BM1s1WlCge/fN4pDCxqN2BeqgmqeyrNv2LhLE4gRrVQUV1HS0k1Uo
O5mFdNcu4s5FZpXNyiH7UvTcKx2EbNqXunc5jD7wmSvBd9ZjZJbtiQX8Uz40YU4t
fNqJzge6EPtpLJqQ3+A0AzFuKH4FgfpxX7iyKwC3kL+alxJgBLkAf8KF6yMMqkfM
YlF/WS+uc/vVoYQMAePRC0q5tVdeMxcdnUr9mq6H/6mJK3vsaqfk83bHFeHuyzg0
1/UP93EgSGP/85eMzzJfbKIKOENNofsZPAb/qVfMKSe5pJ+E6OPS1fzBA423Qeel
65s/YP24DSBL7n7Xe/AmcPOiXlW7sZA7kpiRA5oqZ+6eSXrxTDI9vdz7IIHO1gx6
SOXQ3POa1EbPlDCaVQ5Z6lw1sAjN6CZNvqq3QOreqWbVEXaB4hZNz32OIkbvbQU3
9g08euz6XXklfE7aMzSmG3iRmM1wOlRdXtidVaBNLttLhTgfPg6CPmOFhe0N9+c1
sTpQmrN+39O8fiwpU3OKa5psbLR5ncZcBcF5svmnp7Ig3r+ppInndqQ3MHI4jKGw
bHUj2AKkJ6IcTgGIaOgroJ3FMuX20mLzXs73lItBQ4bqpPxM5VE7thUmHdA0U25p
glcGYGImFRFfaUVmlvX7RDGwyJIC9TOs+RWkqW3STanjvGN6HarSV2B67LrtyMcc
lmMX9NT395CzeVTbFKNg/M6dPAL4Tf3j47xD6ojo/NUJiaBaPMk+FPEMrabYykgA
OjVSIhDavDQQK6ZH/4wTHBKA0VMFBMZwSWL4uwUEhScPMf0+1SEQiYdY8qQUESkq
/6cKQEqLpHIh7WViq6J56eY+kdGCyY7a8ibs8cNfni7q2tx4dF1UwsZT7jQCGFxi
w9neDkXLMevk0JFRu2cVcTfXI38YjyQeOM8XL3+vHp58Hw8bgGI9CM8v9ZXM8wNZ
3KcGyo5eXpsajbIjqr6/VAf4UAN0aLNj7s4h4fcmp2D2XdasKfHDDyqnFOj/8b/O
1WgQG7KZqr1nrsZVoRHStxpAc3NZbP29oacLFGZcI8COiW/R63BkjAkp08ZQa8NB
izE1Ce3pRRsVsNW4CpXgjfJ/lIasLPeXCRxJW7H9ZQF974arKxT8l+/hct7Vez2H
+setajUqs7WIBp/fabBVkI1NAQlsPRb6WZYOe1WazzoSHvPnctiLe8RecIH/vLrl
3+O024DZONDABsGgY7uTgAHKHhplTqlPeCXYY4Zo9A1XX2NenKAFPWgnV1iWwB4e
4qIjQuqrSTNePcFgcVZXPIcObZmGj5JjySj2brnIeoRUZqI0Ex0ErDOhmKUt42tj
XnbnmOfbLrKRiyeRTiU5EmsfCMgNeOWrjifwm0NYjW2eSPoR3neUNYrEjdi67M+3
XbKtrFmKR3kSIHJwdQiKtXxHt76IjUu9Fdg46mWuK/hO7T21ZhTkmAi4PiSXr1GC
/NAzxtv9spgBqHvfzUTf8Hf914ClAFJ9sZ80bCASrrti04rjlQFt3WOLKsXKUBEl
Rfrd2ZDD462MrTsB/0nnx4gaW+qZf/Zo3RwTd9E5y4O+07JbXU2PxHnflhck+7js
BuURSE0AEIeWrSvT1Tz5JntT8tqlgjSeWffUZJfOrG5ICBaFHrUCw+Q8CQzRmLR/
q8oL7AUotPz7D+lqGFQ8H5b0V2JqXK1w/w4ZJqEmrwUfHwADw8pucqVKsj8xu9oE
EFYWaIRC3TljgGX9P31vQCewj96mltTkjc7kFBtT7eZgXckXJn0HMiUHVVdEV5qg
RRebcy0NzZQ2zGpR4aiCJP++FSHZiQbTyCBM3TNzoW4tFJ1QKH9KfFSqCDJjJ7Gn
DXfRvFdvHTYpXnQDLv5KPcdeFyeC40UXrxkSZmhpuTeTKDIUK0C/iSkCIdBwUJao
255XFE+KjEDZnXOiR1vD7HIV3tcLtiJ8i0zy3z28F1DjxDtW4TkL2Ts094ZMD986
1T5Q7tU6Rs4LB7eaqgp9nc2iWneTv1No8Wbjtm3Kpg+1p2f6mDnNx0ZC85Vj1qwP
7/eZ835egI83f9yRwrk7cjeKwAVMIWtDIKm++GwdUbYpCNbjY79sUs4si0qnKUwL
aTuCyj8V/TsShGmFs4pgAXBEw9Oip3E/1GLYDMxoqHa9hCEBEf1yoJnSnIvodSes
qFp7iEmR/OAW6MijAjFSjYuBMySht9KhRrVl0oWTkNcviEzXgTOKi4oix6GRma/z
qroD+2ZRg5VpTTgfhLzJ+f2+1ErnwYWl1ZGasUPKSBMM4q7EDWBcC/XwQZr9ZhHB
XTXqoVo2CMpmbozENei5K+O8dbhvpPw70UzR89o2+8sEsxz0DWRiE1eanPUc9i/A
QA6mFBTY2bIxmOpASQL+qN8m6tVEw64WXMSJHyWfJrPV60Mnfln8xo6YVpgcWurF
Pr0DVCUS85ogKERXTW9BFZVMaleE85/gYX5Aqdw2TgZGrdBljM6LRLw+geR+1N2C
LJc1jtUzammOq/11maMfSgbAqbt3wexLVN33fFM2jJLUCiKfA6VHqxBA+LgEiBp/
fiErFMXjnjGjNbz9hzMRO+8Lxtf+udvAbOftutKYMiB++U0Rw7cM/l2T2bhGvJI4
0YxNiiY0qSpIpXtn4VgQSTltDcb9lgtsyHH9wU8Tce/2HKCVrlKF2+tP+kjQqnVs
0KOnLMqU4H371ol8DKYbH41eDqSpbRdRA6s1WHuwPpuFaBa6qg5LBaRY1yxNkOUi
6uBRsgBMt5QRE64fYOecW/yPiJeF9UyKDPd9LZ7tuY0U8ZFNzjYF81ETNCkqzU/2
yJIoUcdSnHk03dxUO8vOmbYFUXN3rktyF7QUvC4UOK5IyMFR417WbheH/WuW0O7o
DmJ5/okk76yOpedZbOLUsjXC687t6AWdnrvRhDqyWhTURcyxOoE+MtpHshY0F/ut
3Lt698DJqzNHZVv0E9LliJsC0XKpZf0HF4J9JCPiUubVjYdr8FgWuYwSrmYE4dXe
vDHznuH62GX/Xdv0AXW3q+M82nhyP71dZMuGW3wvcy7ltBXZXJSH3kGRJn8CaY7j
xH3B0psEhNF9fjCa0/DYaz3Gv9dqu0YA2bDC0xSAaJvynV14edaRbzRb3/t6oaMj
I7mh2bfW8/r8zTqHGoRJ6k8+vc2DC/k6QOXkKVIZzJkPK/sTlotANqkepQC1H3oU
24u/B6t6cksl04avIG85MoMf4hJXGtVNocl8TbGIxb7hFzPRL7s6AWW5jp1XidNo
OSc0DW1tltM+R4e0EPlIEb7POx9Yq2aakEs1L7F98FGaNSMT1j924FTf/cSlnR+A
wTnQ6VEeZEKX3nbYa7xZxo8MXYPgMTQB9bh50ScSR2bw/a9JKSxRhB5rjGEcQJQe
vhMoMKXHWii82CBL6LR6OyUYQUaJUrnSskcuwxX3aWpUbf98SfLV4ORhBGTE18F+
boXVhkFu69OtUu3bAfrZCtmZULQ8LOMQfvK7GwaGUCrPDEQmBqnV8ckw4UElvjih
HW8s955s2hvHBYIRPcw231vff5n6x3hD7uUklHu2mDlvSfO7YY1TY6Xme+d8t5Xe
jJ8HnXdayjaiyJx7XsD/fEROk0yWzdgESYaEmYji4POypUV4tcUNmAeK4aasGskL
jc6Y5uxIj9azNexKRYWepGHjKeMryWk3pvrxlhD5TAHq/bNzw5KKn9L2Ji7tZVGR
TxDFvCBWWF7v/a+HvPT+I6os0UwmUQsIWgSah6FfyCz3XTr22oYtwvlY3L4PZOFG
nA0IwU+IIxuelk/rG8yUZ6lRhbnNqhEG4JvpCpP69P0GU4rPqH9n7lpsnpjXLWDA
BhqlRpc9+UzsjyZB6l/WcU4gCKLD3ZCXKhW4PXw82n9emC5kNqVMNPUEz2NpDj+L
t2M6yDyolu08Zr8uQi5u2KPSXE3qLfPCh3mXPNoxFNUkwz6m2iN5bxKD0hf5bBBw
Yvr4S+p1pjvYYONF7yikOwJtREYoVG40A0hSnNSWF1mRVq/j3v/EbuSzwuw/Ue52
Qappy7XaFdT5boJ+IjkmfmOH+lsHPXgenY9D5kDC0mdzCCHxC/COx20pfgJY6wXa
CJubojJVdrrB/4JnVl7iMdVNMT4pNoQjTOlmf4q7BWjcF3C0aJNTeLVboxODJ7XO
QK52n+JJmvf01WBQxs5abgw7leSUmQRuuIZ/qYEZSapaUr11qzaBTwhWFGKtWKnJ
Nu2OEpJmDIAniSCzT4UM4fLJ13vDUsAKRtvvMRXtVsqQgM7svFWTsN/yl8O/S6M2
8jR8cmgb1AkkPzJWtaibK1frRhjPLbZSoSu+9XaSIEPrkZ9xkMXVNvFmIkyG6U+3
XOLUddh8AGFB/Mgw90SpB95AQ//qJLSyKF8pgeyK85kBuoHXYl0ylfNVy2n9Q4cg
H7ZtdGa+g+sWzNuYePJvFPBrpsXHioE5vfdvmerPYzJABpuE+yP2SIhc8fFgeZA3
uOjdfGTn6UB77iswTWLUc8PMXJo8D6ocqLLD/yozRoyBNja8zmtEMJkhbhTJQqII
yr6jiGhhWkY3vG8bMjYdPDeIAKM2kQ8uBlv1SuK0f0qsTqwNJQ2ugyrwdbd/CZyy
Y5M/R5SG3FBVyIv2vMgFoDoLwc7Tb0HsLm+bvSAaYD5Cjm/ZMTH98wRJXgs/bpHl
NW6WQJIerq76jktf+Sk32YRsx8SQMVvI3UN+qBCWeFWVFn3qrt328Ap8+ZHXqE1Z
O1SHdyeSwHKi4x4SGplWf4xueeoduSQx6i33W4aZNfbbBHwFLdF8XWIo9eAADYZT
tBsZLxC8YN5tfE/OQ7ZbofDs3Lk+anQ4/Go4comZzoHvJPJFwKf2Bp/NyyT/+f/c
jEZYkyoGFAiCw52PgMfRQZwNCdKGk3s95v5qveJuQGtzFaIM59Tn2ybgWccGHJTP
SMaIbWpj0qZD91oIgKD4436iHKveTCbH8pIRnYuTrlUKGa3csvfG0K8DeuhOBBxq
WLL4arDYK3RdgeNQ1+xY+/U1Lh2BGKx7BaHMgPzq1KXuwJ5zLbRHeJ7yAZ8PxTm8
mujRnl21LvnncNtiaDJ38dNuHT/smdiEmWMDCOEhrLWhunDxJxD+iu5BSygp331p
WdMs8+JVMmDeqnN0UwsX/FJnMoDwyhNBz/7YFqE9bqymEPrdhu/8OLhtcsEy62yT
wQbVAlKdesA54CJznPtfjA/Oq46bs4RaD/RPP0HHYLD+/JWpSfnyRJLMbjN5z+jN
PTI+EmO5ovecYCCho6BvmAO2ghgiiPXmAomZDLMITMllOt+JQ/eM8fLx+3WSP2nl
i7h82Uf8PpO5PmiflOUomyo4lk1tpfMOaAnIroPQUT1HeS1b90CfNMBxwpM+8w6e
Ua51qc0bJRVDve8lKZAruEC8OurA/NZfEO4On0TiDNncl/ywjTAtCvodFyw8sFl4
DrH9C7iM7nuI9FlBxx2VQ9Il9Ax9d4T6tsxuFZiI+rxDsFsFgZk2HZT+bKBg+g79
oq1PGFz04Cthv5jB+iGqT0griPeZ6xA69Y2H0srPyHu++6qBfnUAhNaqmXsR0pXn
yxy77waupe6WkEzu1aZZ9eu1QtV1H3TO1fKl4zKVUkqwJSow6AexNoAdV3L+tOlv
mFTcREP4LivzyucmXpCiyRgmDV7rZoh+iCqkVJ4vlIxZ0FX0MB4cQtz2kID17MwU
gQmbOeR8WmMJoeKceW3xXq5yRO9iwOZAaW8DmuORc8+QFXEKGR7OgrlPMy2CUTIW
g14DGJHBMIUwBCiPppAJ+YYzKpujQBUj7YucVzOvKKsHcsEGHYKSau/OAx7zLGsH
EsZVwQ8d0siB0kKxL7snSJbOT+HQpn23kR0+IuIrOnDGXMfTKqf0bL2u/5+hYh/l
+dewcJINMxcHZ5R+t4JeUzbgkYPzQQDQTkFAIQds8P8sU+L1gqBUvBIaMS3usBoE
JlhR4NYzQqB6HPqN3ZD5JiuAnlhM3M7syot+ng29v7iOAasSJ5iYQbc9xYkbqnxq
shcP+F9PtAYWNqrM5aI9JFQVhaxZKJ8wMkABHxyWX8zXXB3FRpzirP3izU1KbJXC
XfRhl+Mcpv+j42m3vlLDw6wNMSB1y2qCn+o1cktgy2ST7sGhTzxHud8Xt5UaSz29
Y8B8Ea6VRY/Ful5wdFpVKKB8whmL9QzG0mmluf2b28Tu6daspuuVa1+z4uZLAftQ
NoEZyp9Iwt8jf864WYzpoaJAwdSiSg1XMLStjyOA1NR0OnVadJTqkVr1RnXiyQU9
ymjkZxvsl+QKzCpDz9oiZnBL5Ti2ums+gBIBVf57wUmW9e8mtEFA2H9Ed5q26eYD
Ym9tVeAmR0pyv09nsZoU15SO+VqWcRl0kTnnXwa8B9rbof/d20N0ZvjlpcYChqbd
NDd8ML2S3ZY6ugJpR2KKDwEZJiNEUBHSzL7A2L0LaZCHbOA7b0cTJXOkigfV57no
O7chinU1VJ0FwMZ/vBF7E2ESmWtij9WEiZIuzriuYJU3T4nOJNXKXdcKQLQPdS6l
w7x7zbC9JB9bY9mZoZS56sGIlPlxkjGkCsgdnlVfkwZWK4u08ZzsXC+PnkNo0NW/
MZYCsaGXpjKuJklY4osId9MnIRzrFd8ZwC86UYyte6ywC/GjaniVvoW217Wmtv5J
SIbHVlap4nuyjk4nyltun2pPfdjllX9yRWL95qaOZm0N2Q1qv+u7zJxBO/uuRnqm
FtlwR9iy+RYHtDxujAyzxOv7KHEUyBwEVv+cuNcMpB3cRIAM5V0s1ZYf/LP5p5IU
5DiYIzBG3haH4rBtBX46dtlD4lzWlI3ZXVHR7fcEhVepDYZpZgoMyogvSCW7XktR
8XwPSS6buu78infiqF0VfUVM9nagZ6EmOY8W/NZfGprDnG+vyx2CStTomkYiaucL
dhsfQa8kwjseyEMAGyAwSmnZxO2hTPHOA7l1S0PB0SR+k8GT3Ue7hZJb7FOH5/qY
4K9xway4xi1uIcKamltnimgGipl/mUd3YJvdGqOsfEFOx04YjczQ9e4/MFUVr8LD
7oronwAFD/cEfX2My2wDMylhyW56FZJJF+i3rQLFUsxpxtzGObBhsCrADjVXNXzK
Pf9FuItDwE/lz8hjwDkfQO4QDKUFRKmyMtHbMp0DR44YSaWCXnCeQ5k1BWi0bOMb
vMLD83WMJdD6dCiDBsSdMdY7PpKL9US1PWSPVhrgQtjZICXT/5IooyXRoW6fboP9
DyEdENUNBpSJ4XclhTCIK/QBnJqCmQB+nfPIUzxFndP2Hl0zYw3UpNOgq/IcvGHS
edhAy2J09to5/MHcvWWQjwhKLiwxp/esHAYG/3ACh+ZvrGA53tZURn0+CBKM2c7y
iCCz8LDLdEHufLHx7Hbii70YsNspNSp0bsny14O+0Is5CUyHveEKMLlpTKcQcH6k
A0aocVCEB2wVcF7JYIfkkuRasepsje/WgIcvvJO3i0oFPXLg21rKrAK/OBk/yy6E
ZiGYfZDQ4135DGwQ+TPSJsQL1k4QtvY0vClD8BFDfQc+vfah6t3D7VNGw75k8LFh
Qxi2/uy3zKerqjGfhnIuVy8LsuL+nhhdDnv4QUAlsZnkzxdl8mNSDtzMWvPcuXwt
c8DWd0MshfIByCmqMLcmKlICHdP/iXElDfTakItPVFzebjta04WmrS11VNYwCj0M
LFjARwIWh3N5wZwooS1/RPTCpKRvn51Oqu3V4yrw22MIPQuS5i2WKEEoqChys2GG
pVIY6H2rWjQWTwPu+xeKnDcR0a16M6NkeUTEnn1IfMjeJvqe+lOpHLOfJT/fwdqM
aFyBNFZXDF+BhmLUKdc7omVKUlwJnFGj8XwaeuIkwNzH+ChqX1MH/XkMmFxdpK3e
Fwb91Cz6LibX/MsmcvHv9EWLByi6Fe5I8cbptNG1DnXn2FeJlco3+JQYMcOh1dR/
/J6hQHCa3ZcvW2H/Vdqy2KTme0P7liuhCRdarEdY9G5bsdVBCKS7tcRESTvR9BAb
/oVyk3rxNJqfTSfksp3GAeAxkR/0+xB2icIULQdkzI/jKDcq6w9jOS86u7HL34o2
igyNf18RhdgKEdW0M9yYADvjDTREFnMU7aq0Wc+R/fYyZR54LpbhZI858RI4ad++
MOb2kN3+4PLek3eVjRGkoalUXn9VzhLtUpg1ZnTGXoRlbLjr5rj3ytjX2Gw7+L0X
2Up01ck3TZfPkUNE9ELbFRB6PMYg42JjoenY29J0SkXrFGW5iTBzkNazrFhJB2Qd
SfT2RpTZ9BK9T43h9jXzx+39g0ePHWHUBgYfAsPHGV1O9K5osHzpgW7L/OTdsZVC
SpC8NAYm9UvyZb+qsYnm7e5WXwVuHUioju90L4iNX4JMFQneqBf1FLtgfVc5iJaR
2Hb2q+jeIi32PiVEuYzDO7xbzzN/Bknz+5nCnpH0mKXXnqaTBzRE6qT3oeW/9W11
rHzZdKndO7uCNB628S41/cv7FAu4viS8YfurPTx7gK1lOBmFKbSy0XUxdurOLXLm
m51JwFqGB9Gg7GfiFfYorj4a9zAHwIN1SVBJkrutoHtj98sT4XzQ27G75IerO1b1
jzCN80rwD99ovsaYleQNhSJM5d4fm0bmM0jcyaAFaUJMaQAf8R5fkSJrvDVRbI8y
/UdLontlZxG133ztuGftfPF8zWAIUoDICBmawJum3xVRpDbh7ANQuKYPsJtUn3P2
zCheG4El6n4w3bk1COvQBef1wRLp7jj4Poo5jIyj22tk660Zaq+KSyXPH/Yhhvw5
kmgQQyylG9coTrnmOaDZB4g3/8wH1glA23xXpmfSG1vxpZSPZQzfUfAojhdziHWC
uG+chuvVu97eaycwLTIt8raKLYMDG/lebOZHrVrPwI+43YY0Z86kWfVY//YONGjx
cIFhCaXRCnJdsDMjmUHZJmayGbAcbamB7Vc7rMdD6K8fBdO5HkSSVRlSGlPznRW3
4AYCAyywJrcJherLC6mEQh9+CkSgaHm0YODIpM5jazNBcJ9uFjjNda4SmzhiYqVq
vfiOLxhYECqfUPsP032e5YVLkssAJQ/Lju1T5eDPCkYygampOf9TS6DkJb+550f1
u9djvHdjewcebDctHOQT/4Zdq6jrsckK9myE7xy2gZ9dUt0bVb7y2b4ohepTJO0Z
Wv/9/cQtp262QwFHMhkNwjk1XiSbQK7NMK2UNj8wrarClkZzTzf1FRyuXm8pw5JS
WD8HGhQILAKTtcvhdMbvu2gV3DwbphXSd98IKhFJbQPoh8I7z+m99ab7A4fWOKIP
LlQbEqWxWgU2zv4mX9RBO5DbziFK7jrB4xkMguuHunydy1RVHsQYIBHCIeOnpxOh
REOiYjymXv75cCGy6lrFgHOl6Grmx5pR76JNn6PxnqVJoxBpPxeiY8C18bRRmjw3
cSyoKS6cxeniK0aLN68QgygvvG/fugx7bINHl+OdYJVPYDYRZsMTZvDK9u+JRKP3
7c/bOcAn4wBttp155BWU/rxh3UnCvvqIbGU7BwDt4UlkG1rZJdYkbmCHviR/Enzd
5TBrRIQepck0xaFgBbibS0DNtcpw6aYKMpd9RrxQ/OSerRleFYb2G+5XJcvfvLs/
xY7TtFqmGVZYg2bTJUpGmSlhnSMlTL4MnAz4nUbFHQ6vicOpge7Cgu1usK3iefom
QOVi16w2a1X2GI/CGLZVeupV5/N8q8hAjg+aRokGeZXI3638j+3fjeXofFPxbJe9
TEAdmW4XPsKeeNxNm2vK81L+SviNeGLD0zDfidruiYRutRmEhm6QSvQuUaJGIjjL
ejpjV9s8cIS378++YBl+1WpS1Vgm5jbrW9nsUzqvhGikiPXY2WnPWa24/lPrgbXt
jttciNbojCkzOtMRAOeN6aWaporQSlYt8JtzXI4lPI51UWO8BvrZbfS5XzocPRAz
9ZyBEJ/BNdX+QMhvxIdRun2aEFTNf3mwOwn3XnuGFM8J4ICQbHRawkhzdY58Cgjf
VPjUOo/KFwn3HeAARdAF1dnmEW0ffyWjLZv7RF4ji6ofWWfVzhDJtJVbhzNt+Rzn
pR+cuYydStWauLKKZmJUOgmA0JzAVVq+gyHg8kydshudgAlUVC0gbn7MQW78rQ9g
Huw6qddaGQgngC39sp7F8S62kqrn6qlVjydFOdGSbtZi/ExJCRkG/vfBCZV0QAuh
SsQ1daMHuAAmwGv7Q50luTtK+PZEckEb/y/lQ2Hveiq0tKL1V/Has/aBrOfQxnz4
P3MAwTHb7/0mMDc8myvAYz6GkfrCjK+izUOHhFB60q4Lderdd3/RVwoZrZV4Qh6c
3pG2wx6nbN++H+ZUqMEJfHCraqy/uXNcD4d/twQeghVhbzg/ifLZAq6OntPyNKdQ
lIWIOQDLxC6LkN5u/kAbo4xRwg9YjwQT7LOItoiEVdWczxRGxY9d49sKyF3DW+mH
d8wMrKHU7ONRzVRkiV8RqOgRJvKQvVqFOOwH9+0xsuSGw4w5EBBpJ13vXnaDD1Ud
oOWEdF/Sb1IgrCQArWjgnwqRxcFbPckInILNFOltYxcjHc8x615s+SFuI/ctez0n
a60b6oAJFAOJR3jHxorW1Q==
`protect END_PROTECTED
