`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/PxJQ+Bd45GLxWHqw2DxAOa1JnUo6nwRykL5ougWouBA3tbTXG5dFHLy9Zag7Koi
oVHtv75G7GPE0QIKm3pGBRIWOKlzkYbe8UGsaykgv2BdmMdcWA6c2nmFDBCMxiYi
j9a3xhS1clsHNsDLJxyNAz2JIxHfp1HpfZhELpUaer8t/Q2eqZ7tkbMlEeL1y0RE
CdJ6V0X4djB5vxVnlXCo9GxumFXB0M0WR4Pb2+mB2Bj8I/dHDYW3VMcmiBW8aNie
PRtfhIV5ema5Modv6yHkmm92mBkR7YUOravERAOyHRucTcXQj605M+ciw7ikrxiB
1EQGgjXM5ZJRcVdK6sFJiW7LSQytuGBMTFk+iPMWwz+JRfxPcCbLSZc0awtUMkes
w9eB62VM5yv2S+VcIiQ/8ktW0YIh3dYI0S7cINwAWQfp3mtXs2hskTMQegrDy811
yzR0UKalir4PgqSFBxoixuHMmZ0TDbquu5hcuCOkj1dQXHx3RLT11jCtucjLymyq
kKZb3A7S37W9UOLaS+j/h6v91j86Fi/98Z6fj3Tv9RxPiRsQYoV4hI2PBcBerM4S
guVZMNACa47ICqz2lJcwbOpyMXI/icqSom7GPitcdNydLfy7q8/B77nUzTrAFpLB
Dz6d8SxS2tY4XfGLDJsLzJqDp4ugGHOJN1RToSsufUGglNSpW8+QGXDqIL8fTbmM
TVUHTbPzaLPiPkh20kt59Ws3rpyjEFSkhAqMA8Z4p1tUY/vgmCUB/Qt4xohDN/qf
bJnjQzlokHn3VbCvR1bA9k5cKbaMK5+WstboW7UxP1/dA6n91JgOgJuChUrJGeFz
Zz8DzW9maDQe6davgrVUDmrR+MFGAZieWR0QfLMzaVjO6UjUAIhI0GoHHQ/9FnLg
3RmJwa1IyMiU+p6iKQNppOo9YByru+vMo/ORu96BxUFNUAAJLJpSGUBBFXJVUMgp
bDSiofU3cSJj5rs1C69OSr/jXEGvwc46YG6DwlZxdvipFiuU+6TcaaXT5BAF1CqG
4VQe/vu8d0m/xGITCNwGLKakj6OEa6y7CcqWvJZfHvXtL+FyZczX/rR527naQxEi
OczKEzsml3ebRLFWsjy63eoTmIoOjD8qQGqkCQSifjh7h7G0Rrpqs26cERLGfiXM
lia/d6aXs+hiYaW1xYAI469kGR7qCUxVP3p8qCA/WdtpGyAu8v6J7j9hp6MHQ8oJ
uw5qCZKmJk9SpQm5FqTLO4TRqDfQd0XvUXTTbR4PF/Mu+ld7oLQaNf8hjrM7PC6E
`protect END_PROTECTED
