`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XpdFucVXWUjuZRkzO+SErC7AQMsC/1T4nw2KZbjmwFcebL1oUR0mkRyyTEeEyLYh
Q0U00kTapyY6LRKbq535eYYZBCPDETIfhAkhcM+MQWAVQMEeNRePjDXblhakt8hU
vAxX6RB3NOCgLQMRsOGNMYKYP0Fp5rpmuSs2svQc3lj2kGz81vjLjoBhowB/E2zc
aj36HerXPH6ADsCh9O5pLpdZLmYOGzpvbJmLPf9yTuDjH6vDIdWA5iwyrX56bFgg
LVLfD+QaTne15NLewvMjG/wVzEPD04rpc+Gg6xLcLVv8SdVSVHmXIa08IdgqnFmj
gnpJxpLY3otevNALkEgXfzd5Wsx7HZe+94eQR5seX9mimUizBqEY0W0TjKurtuS0
5XSp+6xoLtAKuJD9cHs02JRnIoHNkOirFLXU/8Xn5tlfydF5qeE58E82SOp/gyOt
Hem787bd4Nnxi8vIfL9Z+EKV73Bs7S1TZ3zodC7FJwDp4LHQZl6ce9JreeaEI2qK
xSX7vWnTRoaNF/ayjH1F4lj9oQmWcsJH/Zr+xsInCzqLpReyzcS8B2ir1QHwUFGC
pAPSzHEj+J6dvw+3QdLbE4RTrsZB6aIsXo1OAMU8vXxvDiMUbF4k/a1S1WzfbU17
`protect END_PROTECTED
