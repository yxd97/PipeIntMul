`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbil9rSK0aqZIK2Be2aQ7xxIFiXgFGVLPZvzsh/RuJk68J8LdzCsJQuj6KlfzBmz
DjoIS4rqMj42gSPLERtx6pLr6TvgLxpMAJxC/wBfHHmeg2APPTYEM++yV/Z0jxA/
gE+gc0CYVLGWINfSLs9RNvjgL2ATJMCNSZ5Rbk8VYPjqrf+85GzBIFZy2N0UXleO
yW2MTeq5PyVUHmraFOdXAgaXHm3BHm5OKsUjx1YeCa2bPIDyySNrWN/Hz2P5yz7u
2J53u8q5IN/oCaLzsbDvMbcnMm4LrydzkuKUlU7JmhIwI7hBdi8wm/0ut69XhUwR
TebXhVmEQ6lgLHPfaYS7z06AEtF8Uu17zXML0S4aJvPqRnUJKcKzY/azp0+WIaBp
cPM6AzTr8uRKRyG9hm55E4BrrlBf6SSBChKjsMZ06NVBL3Vz+x0EDc1ykqFS6bn+
`protect END_PROTECTED
