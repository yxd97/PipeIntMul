`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FxkaUcuH+VgumG8Cy3EQ4ks9es/odDXOyLVSCh/cUPDeEqfnNLD7gmfYAsXSyKYO
5x2tRpjCGeOQQftAw21Md68ImEbFBfc6Lzoae0ngt7z8qH2CDEYPgkTlD7+OUXyD
prgcurtdr0Icgegv4nSoN1K1C8kaDrvZ28NV9SexTaniEsN3MeqiKsrVVPiDwbIp
XwwPIoJ9egpAGH5vuXpZcxRujL30NTbfjeSNH3ZOpUoI202fYNugo3UsiaquB2xV
CJZH5SN4Y9094kV/v7hhTzKng096BUdHMbr5+SHuIN+hERD74dzynZa17eBzx0WF
fz0GFfJ9gpn70exbvU3guqcWvVyEDL65/dOWc6q8MF5kMfT0nFcWwH1lVWzlllWJ
mOxGhOrbmlhNPhdozIOHhdOJ/z0YXyRIzihD4Hm2jB/jEJQGffTrUYPEMYgYntav
2jc3SytSyG8pZNhu3cgQfL4W25Jlz3nV/gBJkpNPMsiG37kUMZKLgxfPls//OsIH
HsOKCoj2Q38mnk/FSHA6YRXVZ38LT4Z49h/oiUiTTPTF+9OqMshoAhaftVdlL+RI
7X2QkUzlyh+UF02yfKMZ9U90YWRir6xDcDqjMeQZlmEpJdrW7DuRqPITT7ES5V69
ApnWbgkUkkpaomfG+5VX5w==
`protect END_PROTECTED
