`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rxgcpJ6zDoJAHnsUkWNgfQZlKqLg70rkYo5K7322pFxWcqKO9gVzORRQrApWfvd6
d11yChua6F5ZFZ+9hpp7Lyw4D2/z170f5zVKiqrdECkApo+wPwJk8sW7gJhjxyYZ
Rire3w0/A0hEd1XmTZhIk7mEa+uZg8qYens28SNY2JXZuYLA3ONeOWDtrS8g/hCP
PGxCjvQL+ehGK44QIk1A/DmSSVg1SQfpuBNyJk4GRNkSRfdhehcAf8dZdEoTHJy8
UvMNw9T6vg1qDca84HnC/I2/2g082mjtAcG06YBcqElZBvUqoWBdNVmOGtY0nyQg
T4tt6Bdln9orwWzTQKpdXcb2adssxMJnxA8ic1hqey8sQRlah561YN9e8ksXNK+G
PuE3xGG/AxB0t/etXZYrXtztM5QwsccBRuP17CHDJjsrPCUkvxRumn8Ule8SBoCJ
`protect END_PROTECTED
