`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J12QWYuYAnGeIRiRNGohxipIfmblfJwYBLQ2Sy5HKVMSrW7C7cGj+Sl5eTD10LPo
xafTOUE1R1Am4Jkxe0mngdCb4GeATiV7xIRsWlB6XTdJtaW1Xr55/zLR7+ucKdQW
ifwcKiJTEQHCKoZpClfpJfaB6oBxeJYlpu/JFN2k381Qm9QQaHZe+Tg/+6dQOhF1
JAmNA39sOciMzKvM7Hr9iUSYWCvRGR+L5H4prkWE3a1Pi6xE7kaZQGmgvOHuoMMG
GDiMNlIEZ4d9PpLvwCup3iqTzp6Ltd+zemeq8aO1sRwtIW6Oxdj5ibPbu00odd/5
cGdp95xWGXc6sw0NkUxfBGHBt97lKqG8ikHmyVyXC6hB03tlPfEStVrIvfYyShqp
TWr+22gkJZ/GcgYH2CvUTOMOf8I2pxUfUItGNtfdBM8WoVz4I2lCJm8RnQ7eqU/r
DZVIUU23zA/93m/l7W+Pi+go3nldZL3/CL7pslJv3LiSchEKhkkLdhsSwc1jmKt1
4e1xqgg5sPqdblLNp+IjGpJXx7+cYfEHEc5bYEF8eUCzyDMz4LofaNmGTofnp0vz
Al821njFoCZ/1j9cRSDL/eGHgLVO38kKHVV6q6Tod4ahQb9s9XANGe+7o4+z5c58
hcnTxL55q7mIV4nDDhe8xTv2f6Jr9m5wzuuoUQJ5IU5EHAAz5b2nJ7MN6OVgmmGE
FQCLcC6dHpjdLyTnvljejBPEKyJmi+D1LtFi+0pm8zTdrLY3OA9EDm58eNaSgaIk
8g/+ubi/NJTo6YA+ni2ziRa/TQJpTvB+Bbv3v/Og15uCUPPGDYW2Mvs2cPfanT5M
lITSUbutEabWGkVOLKkd4ZZgre6IpNbMeWCUSUTytI6oa8qrs7lSgupO30So5S0e
BhtGkmsOHKcwApx3eqZ2+osE9asxGU+uIN33MU6Xc2Cpv/cdycxG48NkdeZzO7IE
qCbQ7a/6ETSt84W5hsxJ0A7F3STGmb6Vjo1B2hBGjt2yIEELdwJplNSg9fGfmR6K
FPOs5rBgzHae8UaBiZT+/lJ6dBMF5J9sYv6pysmEABQGdewLQfYRnKmRU91dYvS7
+EoDnuS7P1EFp97wm2h7HhpFfVx3OZvWgFS/6WLMchmw7wAhp5ggdOCUtIddaAyN
LNvjKO2U/fjO3uza+GguSjPAMulqhHcq0g7WZ0zCjsUXBH7sGQOOtS6HTIC/bGwD
XOktojNxy/7DMRWshmEZ31ipU/Sfw+TNgsddfJ66xNL1CTWeKo0H3MlorVScGWUr
ZokS8WSfMLRdO7bGfdOT6rdTS5biGMZeyfhmRWca8aL3DjUeObiexUKaZ4GIt0//
ULIG8owJmso3fxYBzVBNQnSMkFKCzxVK2EGolFy57kfQoakaWJeK68UO4KyKROX/
GGTvUiHVNH/X85thD1vOFks6RGOxo570+wkB0waRlLJtAposBleNoi9Wu6+EMHlU
hUwR244B0i54xg2abDbPZQ4KvrjvOeIeoKHY54vAdQ7xE32+J9/kaNqcytbSjAAv
NgiLVzY3eF1M7WEPk2UfInd4sh32qCwDXoMldFiVNqTajXgGoh9Y9AjvF+9oAPF+
41nbWBNuCazMY8uG7if1rVQEqgHElh8f6I/PmZ5CVxTfXTK8708D1i7V17Ue9hs3
1ui0/bhVAU58E29D77lum8V/NnDidCFcdB0XnUalkBpNO2v8P5waDgfb0HhJlw5i
ObD5yNcI442Y2AfeDzAR6ojKjDyMAT1tK80dtu/anuFNYPUJ+82GanehrnY6ibIr
TmfOp0pn17b/vPqgeUrjudXL9NwFfBnRpsafg6HgT6VQ8G3fzo3i3oa0cM7y5gvx
XgZ9TO9iTj+XUh9aNbHOHCW3mBygRC/G7y1AXfob/g2G+Kt4D3vPPi/wgFr/s7/I
4xk6gPQJqKt1tZ+6CemMgfbvH5JXkZbPtzW7NSYolR6RDympx3CtAn049pMLDki+
LF0eawMcIJ1UTRr8XF0BZJGT47zDpmpxI+z/VwxENO6UQYYRv+P7vRd2Crxr90+j
fLewv5FPyPzgdv25d+nEl17jqkxck9/KWILjg3S2mH9L5Ve1yNDvQN/DK84G0k11
ryZr358QBlvXH7omlovvYbDjXYKNLSTfgYpJDGkGlFiz9FFutUEKQlmikI4E1xRw
GZSkxmXztvwZyk+6Un+BElJ2/JDobyZ7d8+4Il1ZoQNDFpbcb9sNLkEkl3xTWj11
nfPKCJ1rLWiJ4qxADurU/yp1oxnDqFkQtSyDX9o/h2qAx44fzXNrw4qaikQzjwlu
y7Ljp3pGCodCgSExfoSNzh6OmweXR961GSYca3XmPD06d1u6/rxoV+Bra3JOg0al
RBqJjsSuAdUHDZLUW5E/25hqDHEp0kI1i1SLfXAwOjF+L396/g8aVn16GpDP63/2
hDlq5mW78ZictO+HqVf4w+riqVuj/7trEMR1mxGtAaT2FOHVui9K+QwZZ4eYOv7z
/8Islk1lq6VnaxjXgiKg371F7BZYIFgZCowcqeHQT9xSuE/m6oSDrRRRW5F3Nu8b
qqoA3sXv5mIjmLknoLD03eeiRUa17lpvUJ+piB3v2bnCYd2fwD2wrYqR7h7gH/Io
ccX7s28zcZ0YmRRTg1EIu/tzrmI3/AA+8vU2E+C4Er46SHDzZft+BqkT2yIAF/Lt
TUM2AiJCZZvSD1TzIuEXj074cBZYLtgc3zI4uY5ejC2aDjeFbWmY9zyiB89ufdQI
/HkGmHD5y8Mlkrod3Hgl/rMuePiIdjvFi8IwDhb8b1/3KDeZXKE96xSkQ/vz0FJG
0+Q2JEkIoia1RRUko/ILDlRfzjrYat6Z24tv7GzkdUES+o0e0aolLdlb52ceb2xj
DauAPGBoD+8XRFiIDmL2qFu8dYYGxeu6gqBIj6JIXhAtcZUbpISS+KJGIkkQdNsE
euZounCAEX+bc73GcGltOgA5/lmhDWXnrfZ8hJIbHMi73znh8RPSD8j1QM3VHwu1
kKKhMcosguU3/0yTweb4DCqo3/CSaRoygk4HZnsKrn4AH9hu+TRTP4Cj2L/FBFtJ
oXz2djjO2ov4R7Nff2lPWgsKyoRRtKnyff+ZQsrETFYA+39/EGdf2G8cLblZ/5OQ
lcsynZLStwY1EKp14ChbkkXruIYd86Qr4AnrsTz/H1RvhRDBKYJhFgyBgmyslPRY
2SBtPMUz/JnNKza3YCVm8fTeLMy+KsKOXyW8ZaTrN3jQSAnl3AfngTvUuyHJ0AUy
T/rrNMzFk3u0jCNOm9vRfD9M+4LxBfQ4nDllrGJk8li1OLuppS5FFudgO1HZJs8h
4v1E8PU/JIJu4zNA3kPTOBSeIbPoKnrfoP90v2Gp8hWroO8kVqQ+dMptjcGjUu7O
kj+jZXPSxkoo8l70Fehtfjv7FMzYj/G5W7OuvLAb4yx7FxfYpIA2Zas00t2vl3zj
Bf+GjZBjRHLbNj9hP3/K+nycYu6eEWvx5x3uqTKsWgveWKnpH24vpGCuLW77bTIv
6mFlHIc6CTijG5Ncoc2rwmnSH8uInyTE9VAWiX3DU2I5eMyCVwioCy9cx4zzerIn
U4w9D1sSsPhCT2ZS3uwRzStC7mxta8ugPyFqb/6wAD5rVVjVufrdSn6Yv794UbcC
fBPKzg3RMEiHW5rZ1WbfKU9sin++mHsdcVL029k3Vvc4e1gvv0Q+cLdpl5AMszls
X6oAaVOwXScuEGIXUrodLXqzRdTe8TkKXr1maf+/gulYkcm05Gzj7+z6WxK7n4oe
jL3HwP0uh+s2miemqOSfpZ1PLYgFQeHVqFxs3dhlntx9tKFkiFYaGx+WQuG8abKP
Q+5+Ota5ItefcSYpR89iOHPsTjhbH5JykBSctCrz+RMY3Fg5Udbv21w/rrBnW/jS
8dWAC2ErFonGlgwEv3CFUn5yr7ZE+84OGWv7FxDlfU7/OIKwjWNpZDuAgQYRm14D
fsGIAzufx7qjuCyvKpHHDfU8oEoIlhlC4gk9KzXdPLiBF00G/uZw9nLfi/VekfNK
gZKQwbGHegRfUwrhSpfVZVGWlq+13LBaKTxQJNEDUR4JX85pTnYoy2II5sghG8rJ
3qM7RWdU4jLdNbXoQ7wrJ5kdvqnN2Wtf0z4gLqrDFU++pcjLP+1ucByrYXxMxcDe
gGayLYtF4UoNrQGin6VlXMHHwzAVZaokQ7O4cPRsrb9w/CQKaI8PMMHiL5WJcE97
MF3TikrlxTpgHLdcrzkC1MYW8Y5qAikk8/jps5UWUQhymLqIjABiUallzsXMQErN
lRKntIJYOoJvGtf7IDzD8aq/EH/L6dlpcBI8+x0OM/kflp2qzeaee1mWvl2IaUB/
aZ/CalKT7mI5l2LyxSdGWDZPg54yTLtvR6L8w18ikesx6AAdMgh23wfz+H0SBQxx
xz4Os6kKHTOSjtqv7XKZnuj2jf97FODRhqwX/kVbziWkM+K/MFP0fmmyT8mMra+i
4LeYS6ovLnQIN2U8A9B6kxERWxTq+GY0pxBBbOLT+HzfgBWCBSz6BKCqXU8QGY8s
1iVKDIFyPS75PM6cFf1Ke2H3BHSwDkGccwbD51VYl5368gNefybVV/ZLLmQrRsIA
D0lKjEBgM3SDVBzxVdT4IbT0kY/0/mkcEQWQPGCWTGrffDooEbsIiQtgktypDZts
Rcf+6kstu19PQ4Mba+h18WzbbhS11pT5MXfqp/ekC0Kug/uzAaL7k4i+QV7FEpz+
`protect END_PROTECTED
