`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c48x0yRkjZGWsjI8ImeIp4ltcdeBwtQf7zafm7hAxaIIUCaZrHmHp0dudfNDla57
b4objgeammn0RWrK73/1+L39+KbBC8s87Cxga15lg2lElQ0a1q61Ve1pYRWQQshE
jzecg7AP2XcmZfvFrVw7nWPqk+GLdHqaMjU+ku54JovOZQTxnr99foPv2ti+NujJ
eGxJUAl26IQDoehwUqAjgUzFyHSK1UMGaApcEfurh5uN+gLt6XltyK92y8N4gKut
bUvRu9GJlQbQzvkaiB2QMYbxZ5ATroZA/syNahIx0Ck3RlTfyjI3YEnrbFELNkyk
DOL3wLZl6ZKPEzht4jsxzPjI/st+tGQWvzuio5AdMlVm6TSGja1xJrjddkRqIHPe
wolElN8PnwLmNS4ijPes2hb0zWplgKU4SGokhgkDDwA7O3PRMvErGhb3FBB2pacG
JT5y4J/p0SABM+6pIyf3F79tsAScZbBRmKoYAv4492aBnsOvgexAKdxKTevBdU+e
/zXDilN9Lkux8cASpMfptkK78oXElK4GlsvNWQt8ZfA=
`protect END_PROTECTED
