`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p0StQ0nUxrALAeatMsv1QhJyXxSt3W9bFk4Xv+QFXJPoV4J4It+JJwn7Db/NqbzC
AEwP5+JnoTFd8qqTAgiYWRkwIiAneIpnJ+0WuG9k5RTejKVsyFY9m42m/WHUHJaF
gBCBIdzjOaUm+Ei5bm75BZen5/YXkBxYfvPZNSRHOs5XsgzpvUZW4i6vd4jPIo0F
EnizUSPcx8dAavEkMLSpOZeo8vbWfLnRCYnhu1Zio8MdJa/Sk+7JCHqFRKYCtNdn
FE1TqXCyCyT4IG4eLlWYWJNdxmGG6+Mp6Y/XvfyeDinYrPLGEQOdvSRmfvaYrc01
6BbShGax43Lyl9OZYvWM9kApwf7hEzZ6ERgLzY3+5XeTyRcM7caAW9bZussZxTUj
lr+8nyoP7pPFa4g2BJf3okOZx0yJGxFTfO1jrGQZkn/3DYF8B2e4xfC31YPMuOxw
9kTo65a8+SJD0Hvm2DKPH3pOmsxr39fSXup4NQ5JyvJ02kCVlVXUP8OVf0supaj3
hwRj4ORAlx/ZQj20BsMvu6gr2Df6U8CKmG3OYy5h9LD3OovTf0otbjlyEfCswx84
DM04B6uiaTLmmbhRY6oz1BkIlxrZzwXcsOWGfXyQkhWVMyCl7cts83E7PFwHW3pz
iyPKgnD/vEakNl0hB0wd+5l9PgHXxZJGZV+esdwuKvlMJkk5pCbFAXiNTzFn4nQU
JstcH0kpORDMgCmURN0O9fHk1W+2ZFsd6x01VudnhjPc0FaelNG4LJPKWXzyxsdN
RZstNl6/Ahn9VNJXNkkq1mWc5WdWz9QK4vsc/YFr7gWUl577txB7Be1S9K3xpJtt
MJOqMyjbBotPGxRME4mCriAzokcxbtU3gLYaeXCeGtVzZlYTYGuT8AdHY2AfAMSb
4u9ltS607wm0SeHpUzta7MXz3Je5rERLnx0/Ae+6zBBl+EgyBMnkPEom/VNXBHjH
YMxLg64jVYOwSJ1tgJJlLx6C7mE/eEwo9FnZV2YDEFlOsLaSGCxDN39xZwPxRtpU
ZGyoWyZFMtK/za3f7+gk9K5NSCovA9EjabJe4hisRwhTDdUOUFnRuNaBPZkllz09
L6LbiLr9eTBvaEO6V9LEEY/G0sqP9stvBxVU23TkX2u9SdLyo8f7zwoZ60bmLTSr
Gv0JerlTETUo/oOfwQs10Tzmr/rJZUloA+Hb3YWgudgQM4y8i97lFaKzCTl7q6r5
7z7kyMQyWEeTImm+LpkiAyz/aGQhLndjreHA4S3hg8n8Z2BhB55IblYzZe13w9OS
wLfQBPAPQ5EObPZBei4eMYJfup+T4p1r2cmWDki3in2O++qpOeTrD3XdLRm49SV3
IUGID6J0o92+cOCwg2bQtXVgHZrncUXhCe3QRn29tihScf94EohfiwhfvmmL7z/a
9QHFkD6ayE5OT3BtgcXcEXOptSVDfOA0p9laIl4UEy7IuLRM8LZrh7rifjFKePvm
mehn+sfvgQskw5ARXcDGkPfCRjP5fhz8RlMWuiHBOfkdSzyBken7kCy4+81pfzWv
LIlbi+8xsMo4h02hQOh6PiWcMG3yMJpk+pPMpBSE9u+uGAp17CrbkO+0rmZ+uVBJ
RulW4CCEi8ck/uYAnuKMdiiFe+v8gddikk93BGnTG/nnNxI3M/ww0O2AugoSbx2N
ru99zh7DvgfGw3DFVdY/u5O5ZcD9/qMwHOtMvqVn5uVW9E1Df2zjr8DJn6aMu0pZ
lSkFY9VJUnQqKXg2/ITTdWJWL5rTt+5NWk5nUWycVKwV6eCVspMlVmUTKR5HXZZh
q6Bs7evbVgz5oNZTwRvI55PbXEtUT/LQRpVBc2h4zWSGrwB7I0KRAJvRfoPNuYK7
dIELuM8Lc9Qp2yqImFLTeFo3xdABUtYW2yTBYOu/PueDDM7qlpVSJ6O1yOg23rYe
qOZhbFMZ/aG3Klzb73/JpWcqyYIZLX1gdw0hHDMHwmxCcarpjPHraQMbVfLimvgm
JVe88t3rr/45/vVqGVvS4dCubMlRRz6HSaCMQMtwnC2EQGP2wmws89X+MkMLGsaU
YC027UONY6pHltMvTm4sCqbZtVIjv37Q56ntXwkWRFPSgqxim7engsKIIyNSOSpY
RVXjeu1G8wiDSEwdjZyenWQf3+m6d/bVB/o28x/BvUgRQ20LzZL/h6Bm8HHXn4OM
XxciWzvJCx9CpElqU2QPcAiZoQWWX4v3MmcA0G+2X7esAXS8I00nNSbGIVc3xv1D
1uEeddhqX+J1ewmKOfRWz1WmS6EGqOOH9jNPAAqC7952lwTIYl378TfWiuh8saQM
PytVq3CrbTsqbaLkw2yBgxuA0nUMo/o99WAXpIUpu2ZrS2ZI4jxYLudbnepeh9XG
lFo8BEFQXoJizLiwmmk2kUn+iFy5yqeS5I/EAK3jwgKNzsHqg/51kbGltARkaEu6
dWkfOdf9C3TJNOA+ai5WAmX+MZbcTbTlqjKVAjMN4EG2OLnPigt2SUOKKtGORymR
zxLPHsbZMGYO2k/aSdlIQx+ighEIhDquTwcg1BHYcx0f2NyaXsqPD7XBz4qGdJAH
/oEKv6kPtVlsLK6mB21NloS+0uj/YeNnDZu30SnWIdjrsOSlV2WZhzWpAq6Jrs2F
4Xcvckkh+QJZD7AOx0qFcDP6gZQHcxCPO2s17NFhqJ4QvsSU7n+5pG5Lw2jJXobW
ZoQPozALaNcrRxCXT53ht8lHpngT4Bswgte38hisUWuJeBrqf3eB6UfqUziKkK/O
dE7+BEFdfI8JfLDxpYznDal2p/NIYJiB1LEn14fJ2R/smjNgXYku73Xa/zEEEAJF
i+a+I9ja6oymxKZ5GV0SPh5Ndx/F4M7yCJV6YiRJ+w478WZDXsGh9TuZDD/3iND5
TQEnszYVRzINrevQ1vnDPFLgzpdb/3+jGiBLEK+40gWQUVe3oVjaTqAKUZuh/GPP
Whqa+/Tz+fBR3xIV7v6ijZZ6ppNL3DCYcVudGnVWDB+5yhY/C9bOHDKzi5GNb2OQ
vji6n+8XfZjkbSxXLlT/yxsIDRP+40dNYYL80gjw0LhZRGIQTumdEJgJUXgOrjPg
wnwbrfc2Tqv6gwPr7CVGeW3rmdIH5g/HEMe4fT7yOGAL0ieZlzMF9YhgMu5GB/iV
bHCKXnMb/wqc6dsqd4OvJQRaFUpusuX9j7os1I1uCOBVng9xRIKxKqdTm6PGzAUY
Nv7SRC229dgArVkpWnjafOxBhfFJOQoRTn4BX9LvTz8j+6ASulE/ZtI+xIyuQOck
cB2g8MAMgGMTeFd0EXA3LlIMCX/UfYnbIps15T9UZSQinnbbTF2e6GkBqNhygnFF
aVUInhZLki93n0H17jWsG5Ke6m9td3RIloySua7Wip+71kuq3cPnNyHsu8TzvZKp
KWVwTPPlrp2ec4QkyAbZY2oj06rvNvarjl0XFIUlhCnBTFDwKcWIldOwGtMRjEJ1
DajeFJejfu8DeaK2ninoSdCZ7TWpdu/bnRp3Km9cmTbX//rj21A/ozqisvIaxqF2
VySAFzar7DLGKoe7vKsUPQLnGmp8mpMY/mx1UAAy9HMe0kFs0WsAKeCbFiUCN8X8
lqIATw4ZPA/969wkpbchu5Rmyn6DyKzDzJqjM/yi5bB4/6R8Zvhm/+BroCQRD1uw
sqSRkjo6jB4bIAnGdVh/QyTd7aTqEbVQnvB5Ueovbbn+9nmntaGQadGDghr6kZj2
CKmFyT7NnuTH5xbDpbGCvzO3grCD9PqXlZw578dtATrZEV0KdFOpYWCGy56V4zi1
erJQt5uyXxjgHe/4QPBXNLaYlawEM6DsOjCATcnDIiaMbwsmQjPN64/f0UrsI6el
bkalQeL0Dp0++mhv671+3DS5kxlGk/muh/CRNqgumYUeZDN40s8o8GNMz+5x66d6
ubvGvTa7WCARDe3xmXDBVflWJSncoFyC94mq1F5y+n6ghro2pBG/jRifNNCRKuPq
LQoKghcdru+JnxbltmkNrAIu7p8+Mvb8oU4QhmRw4uHFwxEB2chQ2vrPqpGzSS46
B3XdN1RqGNLP1l4XihBPxc+svFVtR/yutMBx3QoXBJIGxI0K6SrCABGoehpamkHx
/bnp7ok6h6w1LHpNuBaXVvWxu+pReSV/0UphbTKxsVQ6+ETQgeUuYZIiJtC9IBFn
2dvyshWcqJYUqtNla6SUZuebG4u2xpO4JMPn756+vwSnfEdCMNC54IbFaKDNWVvi
WEoYXfqi6CRHtR/lJObstPXFw9NxFbKUSjiFSKD0B+gDfiUpQJXj5QnBW3DXMAzA
WukmbeBQyuWYTwY4j7An2ondKCs2oSLHNGdq+5L7HiH2YzPV7s2E8EcV2KoFqckW
XErQdnqsL/vK0pekex0ug9oV4gU2AQKXyANbf9WF4e9qh4GGiMIYFZo03LPnSYWD
B7O6nw2uvT7oMFjPuJTGiqDupjGsJEmp9flmXyYO32vWm9vcRSGfQmn05P/88gJl
UtG95GhtGj3p0ylYhzz8iGPW5l1HJHK2ZrQFNz8JgEP1SDeimxGJSoiYhg7q5TQm
wJSd3cErBqO8CYA7KupcAFa7rFxA9RFzaFy8BE3MatDibWMZFEXpfNwnYzSy1e1s
oJPt+AAOQ//uQNOrkk2cyYEbXIY1Ngu9ojOWC6EIigXWEBlqWbKSPAXQgNpHtiVl
JszzVtdVLFQ11Q4dZJvPsCr/1wemm7y502CGVPUW6rXhun0m73Ux4HrS65kBB/6N
oQ1F49vtAJUXup2xn2XqXAVI6SPSmyFCPD6AbaK87XRFaZMw8x3Ih2wL34c/iWOu
0uKJSU2M1181PuOTaiGh/0vWfLdaM7TD2uUB2Xl7hGdNOZXEC7Cvgq9NVGi28pX8
Q4xXjm2oFbO3YCFM9n3NCwr26wqnwTCcOhEF+lGif0J7hN/uWZDOsaikhAHxq5+p
pOkzGamvFgETz+oS+RENz8CNQKxR6vOMEV2lWSCJttyqzEBk2L8Hg/hJkYltNfFZ
oHjUXutX9+KbVhCpTr33UiPHia3OgggakL37jj6G8fSHO+uyQKUbkguX98jQtYio
36WQiu+e+VoF4v8duh1qufVBxrBqI7hlkb6RWtlaO1JBPJ0LyQEtSP8x6mFfELZp
xaUOh1MspALCNv/aXZochPN7FjbxknHptwULYwUAdjDW5n6MZ2cvXih1SsHyiauF
Rj0UtvXK5114qMAQQ0tf1HK/HASPZaM42zAPJaZO0HTBeIH9L/2NMqxonfwJdhbG
w8UH1fgEqOZ8chYjYyLJEHUYkxOdfh9gVKKTr3CbvIc5vdOOLNUOs5KwjjLJBjz8
nL8UFNJjgXNZUY0A0HANxiU0DnKUiiVqSIYdmXS0n2hGknL43rSlFpR2JSUz13N7
OGHDbVgtsmBgRTcjOamTelEVnf9GljPzofDS7ntJy4eDExO+RRnNy4fd3SSZyzdy
TPR53niBu+yTf9Hz/esCCg==
`protect END_PROTECTED
