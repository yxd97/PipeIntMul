`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aVEZo+3jURw0KYXXoz01d8zw2Q0Dp/fEUqb8uW/Labeok2O3XX7GFc2bhFD4uZHN
RdKX5L0oUSmocglS807kKv4ZK4Hc4vKf/B8RZDs3eq54sE/WzognG6+B63od0Jk9
Ijgh4WkmTSiUA2W/aw1lluNQJq/51sQITvqCb8pRk6tiKckUuGvfbMjUNkkZ51St
dV6NnAtQwQ51WQ4eLls9MX/MZyqwtgCokVfPyIFjuZtRwbk45+h8NQDGn9i3BBNV
PNmoGsn4+7LShae4KqoEoUqw2OSss7yOjiE8ZvQkW8OwGIP91Ssdk2ekEFCThLKd
uabm5q3ddND9ctx57c6Aij5//XYCKLEbDILgnWUfiih4p+HmevNioybglsR29dO+
Em9/1SAFPtFY8IbgxJNqmkWDb52I7s3CUM4EUfvbusM=
`protect END_PROTECTED
