`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uLtn7EbXNZgvzqu7NlWsEgIPi69X+7kkU10nLbb/8FfrxkNCEmtSi8hfWbqw2WpP
015Hq5RIDDQYxGH0lEaCdXJfXHF0tb6LSHwvIxW9i0WTPxolrC13nWv11o/y0x1r
SuE4/nNH9Wr8MEAtGNdQFm2Gt52VVLjZu2YiZbTVFKJ5vb2OHDQCO552D1fDldo0
qhrY2lTVubS3x5Bq3ahwUECJctE3P8n2OksPc4AezrMLYHDTEMi8Akj5q5yEjbl2
m3Knnr9jyoIaXpuj0OXinpjKZQGXA6iL4PsuGN4ZvNTy2m9SCsH6E9S8ne8e8J4l
yDO3WBjgc23z7TtTN4In/ndAbp9KRPEkia367Ri7YoM/hIvy9I8IrFb7zO8xpgRc
4uqiYda0eEVKKN8Dwz+BYXcdBYYGs1lkT6LLMMksG78umeNCa4TJam6V76y+gEqA
KMUp/WUPjnfnMHG4kpjmblrBZQOXlLweVbKNRhMVVOZBUSUDSf/J/AG5fOdRObxY
sXykn6RsqgZC1a8rMVGKo5sWU5YqIyV6GKx1UyUvUYIENcrn4fdHtqjsW5ZLaSYk
HkdelLQFeMY4Ss0boGbxUw==
`protect END_PROTECTED
