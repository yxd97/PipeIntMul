`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ke/ZoZjmIALvO3vlBhFzVjZD9nLIAr+8HXPETJUEgbk/rdqzLBBVv8IGfzcdpCkr
rcBMu69pGqNGwK+7d023HxUjAxkh9TXb7r/CCaAqXfu+7VAv5GuHCqk/WV78C4M3
wGa8Kgs+Vq89lZZ2b4Wrp5eAVBIDAQ5SjNJDgQ/jnadyDTvg6OngW39ppnfathkE
I6sBSHH8WpA7I8rBO+C/QlXzvtNNCRm8zKTpv9tr/wxkkgr2+1SF+ymlw9UaK3yS
8W3DGhW8CmIYmM4YC9xc9A6KMEvsEZiiYW1rLeViAowNUVqN0u8/625VuQ7Tazfn
++JA/Df96mRXQiOSEjMWbKeg3UkJapJqm2zD0OyW4TxbeX9p97KGVEDb5pV2aqKJ
zYSyM/6i7e9mnOCMacaAxLpKCOPltirO+X7Ua+pCrtr6yN02bcMXcUJE3SYbVvYR
ZO2DuLqWzW064m2eL9tankqpwNdykaLOgs8kMOfKMmIMS10FeaFhaU1YO6GSbqI1
QxVTaYpyNSZ74vmgGD86W1txZaCrgi3balN3o0adJ3RNC5ijpdYH6IDoAmgnDhUH
3lMgPeiQ/COg31TIWTLHmvIHJEbtv9XQlHO0U3wQ4g2tcXpozmVJiPD4hC26PUt9
OEZzYJshI/j1ac184mjMCzBk1dkxBA8rS8+nRyoRkuWjI9DGa+1+ndYu8Jn5GhBf
aLjaiHYUyCXrChKupZuaNDA2+V0PItxvMwwuU+ne0uf/E+CX32NqQGNyyv6pvuoj
venOFh6WI8OOs2XWT1fqf1psRYPCsPBo8x3F5Ju7ujoGFo5NnpMfgxTwd3H4YNZU
eZeHInwWhHbf5j7P9yFrjrZ+/Fn1Z+qJxrN70PKn475ky841wVBHlMMVJpTShEqJ
g1wFp4B1QHHc+batakb1otnK4AvBFF2S8n4dHLJtyObEIb9Y6oBO1+GBNTiCVstx
uBnZOo03Vgetyh7439K65bdhlJixySE4ZgGadpRCbomivRl8/L+UqhBQGFmgd2IW
n1FhDjU9x21sbFhn3JytnxGpmysqg5/vrvtFbA7XstfVBYlvrDJ3/Ssp9F2kKCgy
1YIA33ZAIVsOxb3P/Cj+YzQ66+f+aYb4O/KFPgKH6asNgAKLIL/CmP8EVckBK35d
CMTa3q33e/+NTADP7sh7/FdjnxBc8U6QH5khTieNzvmGmiiiImHz9Xq8eqfulFy+
0EpMecN0h9BFWbMBDthiScMLCuuYizsJAX3zAnJoRC1Fnjh9EuVHWVlOW6LvIhZY
YmsR5UMgTIJ5K+YPkRyx/yLZmh2HyXDaC6troNJueoVlg7vi+HUTEyy7aNMqvklT
I7CQwXSjXtcQbgOABobCMy17ubDeSW6AwsPbIkoyRtDnkLfJuSMBeQl0SKDKSfe8
xpaZwr8+4bUToz2+p7tauVVtbv2EvOqaFyZDAz3FsD6E3LFImNtova17wjRBK45d
dO72vEUTrTFlPAYi7YWaH6InVUGoX/tSGZS8+bSokJ9hwzqmRxHd9fqTr1XJ4ztQ
+eQCmZ3l+qNfotrXtUP5EPMW1sIevAFiHR+bZ0ram9tfsHQ4IjlZ9amhfioV0pqw
sAa7H/aiCGoZHSvuoWkm9fd6O3tjMkPPIbmoOCJiGMqeTNI0dMU5xqZDweLafmLu
VqVZ+2CL21RD6GEclo5YRm58Xs1GzqMQG/LtdUb3rSomO+JaJeX5tZRESDqmXQV8
LC2oGkhueTIV2vP9fZQZxo5GPDzckAM8XVLSczccHw84iPRYyKz839nhjX2vKa5U
4pWB6okKMS8ABPsYxrSnWmgeI/w0iNsave5xGwffuG182j3g/MgQiSVAN9ZpwhzY
DSb1Mg5TGOO7FWfzP/J9YIye0OB5raSRH4Z8er67E6xATjLmMt47JvCXzoejej/P
UXiaNle9VqWAxFH3DSyiiyPJ9DPPxQslPhvHHVWUVtn2z3mmvIJqFdrIG0G4KmLL
uqaQk1BHqilLwPvlsd8cDlvbtKz5F7qq3GyJNKzkoIHbsaFmJGP0bWCl5Ic6oDus
Zn6FOXRHaIqQ3yoCqv0HNmgUfAkNefiKXsKJMf2Kn3Afrw15ohfkppof51ReBvAJ
pgL6j/sUil5wKfVpgz8UtS9mqCpty0F6Y1tv5m/kaqcbzHZWNhkfTuCaxkW/PTMi
fPFS04Cbs13RWJakgpDbA7BqRkBzi7r5a9p+cPHRojT66lwJSzEcgjuyysCXMfFf
aZEHwBTyFnzIPhZ69Q2ZoyTASYjXmwPqmeOHEflF2gVHLj+AmOLK2C7Ce/mKkVSh
+3Ue6g7Rj2xYy5u7xcI04WnfcgOP4xPol81LBd2gLnjQgbP/uurEy3VMIsTDdM3g
jdVKWgP2Hz94aGghvuhjvWtj3osBe5Konc0ON8ip+9p0EeWzvG9wK5GViNfCKQyE
mdbetyLYBU4eZcBOpgxjtvT7S0NpOgR/F845+o0992D4zSgdxder2lfzC17uuaSc
KMe4wpqAHnKB8Pn8MI6GQ6c756WizkTFRLRwnN/HgO0Co4VpHLFAIcTsgBAj2KIj
0QJMaxX3HC48p7e/szMPVxMPqmofWNCpij0iPGvvI0s3ktNQg5cuwUfw5nI/tEKL
RjMjwykXyCCFEVBhNk9CDQ2fysein/brfFSCetzhBrkOJcpBdjdN/Ug56CoNChBD
d+EnvQMr6qEnaJwHYiP168e8fz3wLYBDOJAjDkq+iS8Y4xjzgjbeWpw85Vk/qOih
ox2TdfP6cKCoDWHlE1L9ENfC/grzRilrv4g7uUXGtX82Skgne9MkUDreX+REM6T4
f4H28hIvIsfThXvY5NZ4OaqaJnzBZ3D8USx03reYC+Q5dp0k0mfrOznz1qhAw0ij
/6rHYEk/1nyNX/dMrdo1Bxl0fbtOCtIPR4LDFL2ctPHh1DYJHaeLft6DENJ8dg03
eR2c4Vjo0o3X2CqWQLIN3G344MdipcEg4pgyc1ngfUWKEavs08KqCARyBYuHoWoN
JUwWS4Jz9Me3z8VbXICNSYSj7fck8vYDOnL5gxNHGtKVGxhCXofZBxklnb6fqNL1
QnHdZe2BhQwF34VWqmy8D8kzhqoVVM+H7RUbBFRE/peCKkmjbIv3WAQHLZQW5pLJ
bbps0lddLLwoiPtRMfy4ZHxU06oA6DikmhuLSBG0i1kJ6byunt/FfHLGYugqunFl
ZrMUbArSTrNNT0x5eZOEm4JAhs9Bu18b95b9oH8mW8XwhSvIdB+VH6O0AxJJzLin
xlJgm40JLnHel0o2J/L6Fdt3+Q57Z1Ox9hxatmXf2Q3gXNbZPGR/1xhol9Tm9VS3
6jdre29xdbN3wqOMetvR3aVmgVcRMZL1MnMSV4evmEjG4/AiaeTlUifk+/WxC5ai
wWmvfe8CB2rzReANm/+Acol+8WqoMPP0Jda44U3xQj7ltHiZ2NDkrLHTjIlp1d93
7R0lmgjmTrpDG+/q5CvOdadLFPwAVBx6Mqq0aZY9N1/8YsKUSDesAnwnstp+ETcv
0ZZExJbxSFCIKWE+rNM99lcNBNnSb6tzUx3noGsVtp2FTwoMXGs7NLUJDZ/BWqao
nkcA1Cw32hxLmae/Vtmn2s/hEYzfCkDFqWM96oR0PEd8TNxlwtCmse+N0KIA0nXg
3eREXW/vtcQ4FijPtqvxSzeGahLXxfPYZcoPcSIXg5W15oJrQDW4UnE5v5hz+39d
Eu6HiIqmD9Eqv/09PxspIgXwsNv/iBs/fEgaQoSNBZLCA94ECr0sMoZr3zPgi+CA
JnlwYqCEsDb3BsCCv+rs4Zcw3/MiJGJ5QiqnPv1vRCqFcDqC7/Q04GGsFT00wcsQ
H8y0Lu54rgZ5Gj8FSrhhA1F86mu+FUtdlb8j1j8vJ7UsznioYKbK0pDLKG0nLGg0
WFiy2/9J+eaf1rJP/71uvdzUMnYcaQUS+PVqp+jizwdxF8iN63f5yPiqIbXx/lp4
57ki0/3ffFCYiWejKNrfMRnPiqArthmnEo364bapSFhCaWksnBIFQL1Nx25yBv5b
IaZqxxaoNhE1PwqBs7vu4Fph0s+/DzVSGsCmz69rXUMgi4XTlnoDotypCNngLZRm
CDBm1FM18DawMBE+YKxgJZSSZjVSZvUcUn/7sANGUK6g6xcfppcoSU0rCrc2DLJw
kXoBYSG3UgJptHMC7muOIMpYJ7NzXGgoPCuy9sajmJ/4SftSrevJ6QLjzRe18sEt
slifSGX0hv9oljfAf/wOJuFiF9+SGoWOj289MObGG4tItlUiLkZjWikmfQESypwp
4wnvC1XpMb7+9FF9QUMupYhgaFBp2cE7QFFXjFdNWnKVkYmzP0aLFAMrajv5FmJG
2zXVs4j4SPGi5KgaqocDWa8X/ScNnFtMr4IPPfPU2AWleq+CC5TZGY2abyxoO+Yw
283nj16vUiUr2BMJaVAsWzCk5wyN+IKaIJtjfdpsUfLMG1ZcOh8lKFydxwKgJKL2
ULg0VX4eJJ4CB5BDiZywMO7eMGsnRxzlbRetTfEulMlEmUnED9gfJD6jPOisEcWU
A1r/W6LukCin2wvoJjji1IbRzusWZdBtWvRIC4iWs8Pd2HgrALfhd31hEJj2JJu9
MPyOzPWIbfpUIK4XjtjzKXjY4wsMhXZwnjv7qCwnzLQ3a58pGTuh2aE/JmuHgdNS
UV8cNh8RqIR+DfqW8ff8Ez8hinZ4na/b71Lq8WxfZy5tJGIhmE/QaSzhXcMSXgcq
M0e/LU39478xk8wGwoPgOlgmEqd0RH4X3AfttJdQx2Tmcrb6ttbVpfIKV3q/MV14
TG44NQryY3cxyoWo7MS3dB5APlylOmeD6YothhwbhR7dr4O3GAG2396iyhOx28cs
fGEwVtY+3gdtMVmgPTMYF056WvoVss3KW3jvypYahR1Np8NR3zVdH1LeN8pPdaQ1
Tu3J4jvUFSuZPo+hX6YMR0wfq+pWP0R1ZbD5ARSMXnwFV6ODpZEZEpevbi5+WkZe
5AcXu6UlL1FNwxrDEMtOouN69Kv3VMEZig4NnkKOoMYmRSzSj4Y3pibVjYi083bu
p4KQ6yD8HFsDOT91sIhhzPVAAhj6cs6SX8dIWp2kTa1YbIqJsQCd12wehe/sS+Di
6nsvn43xIZH4LEtJSSvayGxXPwx4n/mtAar3OBQxAfl7rBw8B5pvQi4PRxFAXhn1
jiooGonbQKsOEqW3cwP3IMKvsuqdK6WNcouSDW6WpC4pjvHa+80KHWKZsxCVIc3u
XFvk/iTM08k170upue3FbJ4rGtrNUA5HgU7vsdwIICxiFRW+PCiWuGd5a4YNJXYz
F1edDMkiK5UbpFhh2Ao/pCzUf6mWfQ5wiD84dmdtYQVI23Weol1C8rLEosjbNSrW
0JKCBFCiHCVG7EsoXR7Xc8u987Nqeit1LJquGpZaQeH94QsQZREGCPEzCDx6E6p0
llQJbl10nak3vKUuWO9OmXjQ1lYoSIeM63RocUQ3UmCyYB2y8t9Ty8JPN19NCzMM
nD3hdBI8o+Pafr4QzZ2KaLVVuaHrhiOj0S2THMbkoR4PHU6CY89JsEsTwurxtZLw
YmyFnhu0/Z4ezSti8ed8Eg+4R3zBrx+yI+czl83rN1sb3e+cONkf+Rh5qv2Zm4GV
s4XKZzKXlWUWDDNdHxOV5oJAJ11Sfxnriv/IiPsF2BNm4OxaO/eXbWepu4j4x1/q
In9yUekpleaxlT38OwysUzqROAIfFYshuv39FPSMLp5MyPdmPWtjU2eiWIXhzuiX
QwFLFAYbbITxVC0WxHSv4/ec/UHEmuKl83VIn+nUZI0wRRsElAWEdRE81EIFHYrs
tQOKmfvnJ8YgX7hLOPkoYAsk526neJPvbn1v+tU9xnZQZXyx6WwdvZLYo1z53cIM
LvN3vd3vVVhsZZdmBYk2jjDbh5bxWE0lsW+wKrOVVHFNF0/ANjTwXDW4f5vi+HHn
Fs0muW388KW30wEYsg8f/Ii7Q51QBfwGkmOyHmPEA803LImpVWT+AuW2cWVcY6yN
lZA8h7LuNbVFuQYHL7v4oVeRAfvbVQqsx+VgmMZceeilCPU7YAVZlXR+GMk1x3cl
KhjSMqo5BWr9+qT5queKdZbB0ZHtw2ehT4WJCvzkhWCN4GkW5d6M0PnAUcAF3iFr
JqqBvp4rjgmfIIWyKKXtkqoFhOJfHAjSXbPcpH1dSmotRxQQXrzUW2v34Eir7/7i
MSL3h3vNOIjbGuSU6dS7SNXH0HHIJ35hBW/PR7FU4Khr32zuEMuJuGqCeBleM9Fw
eftIWIcxKmgjJvjcdQbaVj+Wq/r6jRdolNtTECsQRFvul1Ju/CUM1iDB8FiMBs5l
iWQTjM7s6neNZOZEZY9rMw0QF7b9B429Gb9fY4skKabnHeRekySSZCHFpH6c+Khv
s6hEKpqflhpI2S0ISK0Ciw8tZfJ2HwcAtztC4fURN4bYivQf8OVVF2MnVKtXvzkv
+H1cSmSy7YpgAJpCbALVht+xaT6mBhE+2YBP7Iz4RJtoOwtBQqWCGSnOgxtYaG/+
KNBidGdPm592sGHB1rtt4qYuwjinQYIz6BPl7pCIKQQ1rSOYiwIZHAk7gujAmLHr
vklIinXharyD80YHjEH059mS+9j2p67ZyXPsNJR5qHCeZ46gSBVRnvEmyaKSSjRO
NIpU3Gcn8nB8tbbnRfjzteoDvKmFhYQegz/OYme2sQkHwrNoyMedEvTa9m2/hy9O
Kgg20XFVj9H6V/zgMIv6n0XfTo74vG0+1DdUdlYy9+afSKiE89fko3KwClA9tU93
XR0b8RdGuVVbWE+yIk5AkE2U5WW4VXhpTMhsL5culdwoiJ4sqfjwYIVOC4Vv+w44
W1w7FJyAj455zYBrk5gxP/UwDRmQ9zm41TidWVGBRylyZqVo2g0gGYFoWx7TQzoJ
XWhrdu52n+OqYP1bROB5ok0OK5gFpqAoSx3CYT2TvdGvytT5WaPTJ0rYM2rQ4nVf
0MpUhF/HcVZQ7N9h691YG2xj6xJMZqqCvOSMDB0jZ9UB9wveJ5YTLzNw09sueRZr
2N5ApYVgIZ3NXRmrrWDhnCw8eyenzvovvHp8iyvCSDyT6NKIkPSHBzQjMdsblMF0
I33AFX1piOHDkwylaUzfLMSpcQ5mQYRbLt2+RageukcIWtM/a8hcDPap/AWtYdha
DE/yN97RQegzt6mzrWuujY3p7LurTBm2m4cBFM7dvEDr4vKT3Gpb6JSRPxUEgfK0
UyGqihRJdWV2ANPGZ+LF9tSXn3DrcYQVEJPtdgQC25ynANnIIdOa5XWGLHBAbI2c
2BDldklCTRYG2CzX9E7DmklL8IpZn8VAN6B4p+tvSGI1E9pmLBBezvJ3pnSN6FW2
7fVE+f1hzoP/4wQ6qBAwqTqwqeBRuhN17svPaZZRmsFD7rn8bxs3eGrNwtF5mkHq
oi3IvCTboKd3hiyfUgOQ910+RQeu70sCT2JE97IKaip01iragYhkHuSAHfcwshhT
oWtsTQJpqlRdPIKBDSaM41sVtGr8jBcNwfIrj9nFxS2/XWOvoKeRHIRUAaiGVqyA
vTKP4pN6wtLPCg4UUMiG8clc78CijLyJ8RvQy7nwoIveJitpUN8jn+ImgRQu8hPV
X7KRR9/oALiLhhodkzfR5UZJlncvEkz4dHE+HJbuIqwCcNX/hVMd7WhMdpbKr5dM
PegikVkTHZ4D8Dy/MQxENhnyj8nDjFKFhURaRLFaGO9i8efsLJOeV5CCUYAFq1Yf
BaaOivzvU4g9jI/MGhPw9HqcPOHprj8YjdpHVtkkmUFalQW9G460pAZWXL7Z7uO/
7Ta5Bf4R9Sri7kshSa8rLGrnn3K3u6sfJrPs4OAaTd5mo0urJtJ7kZZtfLUN+n9j
MiQ1ldn8D+o3v9BoUiRpwOBJbDNlt3LCMFzFK30539zkygE+lHeSUIvM2NdbijkJ
sp7Nmx8TO1KzWv91g8Ijv19WLO5aCzF6rhOtkVALmY0F87yeOBXq8ejYMORnS2z+
6MZ7WsgBEHqqQegNbCdvRygc3WtaGK74BCbSbsyde9BBvwTBHDYtWEO6oHMZ3GQk
iYhZjJmMUJ/i0Aj6pHGXvZRJQDG9dZiV9Byua4e7H5S+6Lnoz2Cu4AmdWlqN7DM7
TAdIgUi03UFjqBMAQF+FZGppwQ7gLICbUC3fAi9jQ5QxUheXfh1mjibEThL+Ckjp
dYQ65qziMKjXbDAhRpipI/Q0HXHF7A93lOdAgZ0KxhklxDSGaNrtp6+eJmOfyBU1
nUWsbqMamXnrv1TWQJsU7+JMXEvSE2B8m6BsoX0jGrbi+kFfSfGY2K07rPSEtG8M
uFy29Tk5BlpM7Z7STIaJmaD5IiaNGoZi7FaVWMPoBJjXNQchNlCE1JqW3SDvrcBs
CutI7VeTolhZJAfsIKv2N+M7bm0EmRa7B/dDTXCSA5HitG45q6Sj6PSHstj3WZYN
V6rgd/Hicu+NI+Wu/qncyzq9jL9xfzovPhhN2To7DUW8dYUe6wTQK48+/kkZ5akP
C2EDCoxpmb47MCXrWmzu2mna0R7t8PiWDDuT+r//u8ktJX948OiojMwaTy8zpm7M
MBxaRxLvhmLm7oQ3RPrJ3tR8JPvrKvQx/Xk76Z3e8bwml/WAQGkNXSUhQZ5trx36
HM0PyHgtPQgQ1t2dOtRoVxOXGQlqAY1Tk5Esi26gBcTzSvprKQab42i1vMmZBA3n
5kJ3cJlN8UkN5bGWKFRReh4ZCRKoV5CBeRuw4ias791oe/Z+EkBc4yjvQiBwVoVF
ZLe+9acTqHGfV3ylNGO9r7xwY4XjYoLMSuh/FpMW6jcpo41yvk+QU3TScNyUI2Uc
pd7GsXu8C67jNsZ4tbS3umunrKzQPog90ltDwO3Zo+h/CBvskuMwGR4cliFOxtR+
ggWqVuuwRB+FD+WgtsW+Btnejus47A7tARxdPh9N9vRBg2dmOi0bCvZNgMdwEqoS
Mn2eQl8rbycaEc7BUj6ohC7ejaG2n+Kh+EW57NYRI4onhw5qSNjz3f3tuJE1r6OB
KjQnqguGCXjC3IawVVN2NeLLtxjUKMCOKmspcgsrEuBxsw6y7gsPaX2Z8BT4uXaq
0yWYsel1Xa54d/iuuVIyw2leYfK9ROpVjrm+leZ5/gVRgagWwDXTbqK18O4Lz5oV
hayjBBdj8H+AemMxuecDjgUgX6vnkNHzR4CT9Z94XU1XPYzbCzcDI/t5AkzGj4Pk
ZOGqa4pFH9G76ciEm07jwV4BJeOkKngVUnADy/oaxCsYBbd57S8H83g9FXsSW56N
JKdVa0RaezQQJfFVYdLqZVTmCVH3cAA+efPGXLJYDgiFtUvp0Bz08I/Ha1g8/2pX
gyGk9sgkIR+JP/pPBbUBQAGUdjXqfQaetAQygGUsHRQwqQrH+VOqtRuO9cFxSr9S
vE8Cm4cFx+5/UcSmJ+IxxRCmic634PorC89d9258ktQcuZ/vllTYBfZZ/d9ZP+Jt
2TGTj75hgVFAKJ4htAOsi+REZcsP/a2pzM3VxBx7E1j1eEdOWkZRqla6Yec36vlV
nPEHEk8nzFZ+NG06kwc9miyf4LEjz/WX03sczgrobNtYdC2svCHU0S/8FjeLL8/R
aKp4xRrimd+BvNSraNB5Blw9HyTuuv66xaHr5/2tS15fkYqx5s0aCmswpGvQ3uGm
Sab8TCwe1r+ieBxL4kp8x5MPF+I544QYhnM+X/G6zJc7xxbMnVzNGkruQc/u8CD8
ZOaNX00qVgFb5TgcY4jaYRduMHkCIC8Tdz+miNCjkrbmU2A7mxDIeFM9xrqmF6+p
0/e0suKHm850hNYXw5Ehrsf13xMqpx7M4drUKtDp3wDPwgXv52+/Siv6TK+IOBPD
ZbLJMQ9sY6OEcW2QpLaeKPoyXMwqnY6w9hsHH01fdpgXBlKsuFocO7Bq8FP1POh3
vrjaxSqaRIBsneqZy00GhPALP3C1y3ER62v7HZ0S+ouptx3WQY/SIonHhVv44Yca
p47GtZQ/XKiZyVcrYJHOFKZKe+VOCg3cX+A9x7DVGEVGQjiM/EskKl045yePG+FU
iOF1J18Qi0mu7t6QQIFORiU5TwSBWocD+VZg22yxGejc2uq3zNefc7iLHMHiBy8Z
nqw1t20ILI4B3pQ5x7PzVag+WchqUeekAZLfHfqjkj5Cu9W7MYfEeYoHVdnbqw8a
ufqmLpJhVfAImTBwmVG9cuaw0d95tH4sYtQtLSOrpagC46tGW2kcXJyjKgoFXC8n
jU0ruHu3EiWpwb0DX2jewaNko8+pO8xMsSbKUfGyZxXkj2a6Tob/y++hBhSyEmkt
G+4BBYIfvmrrpfosZ/cf0gLBnVYFFkmG7yHn8XO5y7VkCiGWNr1NhA8VqXifhcwp
1QBQRpbykcwY/KB4RFZkFhpE6KgllaO9KGz7qMe7McWbj1d122ibfty68Gnr4q1y
ZheFTa9kiFzNyiBz0bLPjh2QhD9DJ/UtVUtoBlZ2kpvWJU8lLMZcrlv2+15FP54L
aVKdV+7Ew+UIi1MrqVabJQNFyNYi/HBQrRIXLeyBCiH5niWKNi0fI3fsj1v7wJ6d
uLhClC/rqeBGKsPBVDN62iMtIrKoQYnZF5b+2mN/gTVZf3VcrjIKtiW5f38YwGQ+
aho5zlzewA2mhbUlQhrwwjqJF17joGkEtDzXfZFiskbar3JMll/IdgatHFddsg37
xfW/VSEwiOiu/da7AQvl9cZRjM9U6dDKjY/Wt4uM8+J4SEPexXDYVZqNB8RMcA/f
nfZZHwJmG13rMnL/xl05MMDQNFofSTzb3MzdvZtCaXz5zxzQZTUMDYPbrSMIi3aT
Vwjps7NYqRFeQ26MK6znAjcP61Vc8Po2gVUeohbyYQblJeURd7QGCJcB7RFNoWNG
AI9i/GI6BCCoUEIPVK7QCQ==
`protect END_PROTECTED
