`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7qJVoZUCf/T7IcGLQj3H4beYvpJ2v3n56AWEHD5RO8okAnf91SyFgrCMwoI7On59
w+1O0CEM5ORYLNl9+z332NMWuc8V1epMJsCYADxgp7UvBI+6A6PIUdCF6715mAK3
KckcPxfq3dmQl5DKQHvBI8L/osrZ77EyVI0qwVsh1WcAgtAnZFCBEHHDJRy2KbMQ
HvR/KCORr4BWbIElbZ7jRGaP4hVrDwt/s7M9XdW+PBCUYUhb5da1IIaQHyA75OFK
rTCq5qLLaJAg7TBs38clN/4fd8tvPgp3V3H58HQds8SWzgj/jvIUCx7YC+YChRtC
s0K2fCJgLLUqVm6HDCV+TYxOjvlC3DtA29v4F2IELP+qpY/Ny+0JPSgAzLv+5Yk3
agfLdT+ilPI8W5tdkOvKTw==
`protect END_PROTECTED
