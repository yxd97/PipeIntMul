`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MBgTbC2HiF+ml4k27HEgz8Gu+NZX36AESlsDD7rClFd0pnbpI91jO1vQUKOD0qB
5EkLzD3BmKfi0+8SrmGQfidbhR5aYNJG/f52+cDh67YxYu1U6+Or2sO72EhZSHEt
PJ5zhBPfKkLZ4FuJ8RFel/A2QEZZ3HbCmM1pf5c6KsEi5yPnn2wtUd8jGpYNugd3
QM7cPKsBlDFMWnYEY8Cqk8tB52ItFSb2yCkrJWilaT3qcjix1UuZbiKIVID7VZHd
jCT+Q5kBbY3rS1go9JHA4aeARI0lRfkgD52tsXhMc1xUJCSFYI6bMS6XLl6fCfqP
42B70UcBrgkNpJ1gbztKe1RqSkDqzOQ8UJ4psycCETv61+EHvIFVxDhLqsep48eH
eaHDEZACI0XRsI2g8FGMcxRI+n4RLt3g8L4aoHq8r3kA41MRDfRw529lXsWvtgR3
WPZR7cggsSH3u0VmCkGCdDyPKihhBLpo7jwEl41rNxRqG/1aheJGUIZqQY0z8tw4
BK9Yv7jUGbdY03vlkKNeOadNlv4KkCpyD/IIy1Q3XINIEP11w+Ikn+iyBXaw83T6
3dROHL5tvyeJW1pjgZCKoceQA9atnnFD6K6TkxKnh0I6lglBTopkszlwERH1GAXn
k7LD7c6NaDr0oToqX9hsYPmmhr0UuFsClTOqGwJXJgq3KYNmN7RGFevubcDEpxV2
YKQHCgqTaTVo6zg9+GZZyF6Wk/1ve1w4qqlJoUovgGeSElYNucHE3Plh3Ft62PUd
aGbPSrDV2Srle927zAE4jtkuSeEBvoNx73GoBKKluI1P/pmlSOMNeCkhb7fbdDOK
M6RkN9UHZ1JbGm464UndkzecV8Ie0WgPRhUMApj/BWW4kDDfVxukWdQWW8NcDgB8
Y8qpCzGGM+TSKZoFUVNXpbIpqyZi9dnkpYVWMuhE11k4lGhNll+/cXYLr/5j7ir3
NWiJCXNMAFdQYwNC7+U9YqmmyJVNwMKKkvkv7fErA/wviNvMPaGW9dUCbMXkKIsF
rwzlsbXxtsO8OWTJ9MkmGh3rkmekP3emnCslb/JTJEsZKmdtlZ+ug/pRZMlPo+wq
1xT8/GdkA+L7oeJXktqUKfzhpCFseIvM/WeqKtCVCMKJH6e5n1pMILec4tX/ZKEq
HySHgibCrKnBSS4ReQ/VzmkMpOML720CDdDP4XkqPtV13BfOocGoio2WSBfJCB2L
D0H2tMKWJ0NkFH8gxRgXdOseX1rl6U6HWuySVkxgEFfDF/DrGwuAkw7dvPAn+VM9
lutKlGHU6miMPgGCC3IIAsbGnYKPihYCRDPxSmZAJ8UdXw3Nqxow2Q1SbqLiTO2g
jk+ucG5Nog325cAFGVupXpP/OID98t7edrS6hRrxz41iGuNFeuzE7q/XeZJ+sX3q
YoXRGw7iAxQfVTYRdzV2ED24fdSMr28qYfNFbfLytDp3bZjmkf688Y772oU0RIhc
RMNXqZ+GGVHq9xz1+hLvQg==
`protect END_PROTECTED
