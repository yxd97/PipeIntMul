`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvwO9VGpFLdgLt0bXQ10Avo9Qm/CuOGxLud35968qMUcKz0Rl6ALy46qbAJZWjhP
XSCucq2kDHk4ewBtRA/aNiwUGcfvD55b0qdPj+juedBvjCqYD8BfeCTrdCrn9XJx
rzvpiGfOWfaiSOKeOjrZiTJPcmGFMfeaw9RUh+/yPLuOQc41ShH0DklvADD6Krrv
id9EfHUBPOcdYhkDk5pOIK8aS5e0XWy/m8Ll/21xGVxnidU88lyC8WSUgypDRoUa
BKg8qWeofQi+gJv8uioMyjxzsjpExdNoGfYm7WiVlzB+0MvDh/ZtQKg8CpV9HeHM
QjpvjM6UFXv8K0aRApIvqKW69PEhEcPhuAouNkUN7jbztJnLqkFbahQNqpU2CnpT
MF02drVqXZJnQaldK+VRC4v3VYguGXMVR72skQTpVBBeGafAaOcVCP8772p2FG+d
RghF26s9I1DpTkHl6Nlc5IpWu3PIxBLC2/RbLHHVXrKC0QT6Umy9FeufwbsqUGKq
38XY9fwF0lvwTFvJ+ndVIlaH+j6aYJRQDu+pnuKmqZLl8TyK9oH6EABO+fbnnP6L
nJqm7gJxCRa3UI+uGLs/l1lrwnVl518f//PJ+FCV1x0=
`protect END_PROTECTED
