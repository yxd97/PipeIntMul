`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M+3A/qR8VkDMVvaftZKJTfh8lcKJ7o9uEpLye3SXaYUGB8FhnvacgQ53yb/5jSna
S5FwEXY7d9FlgKfetQ/odpAi+DB2JtQaYTTUm/c/BtxkGbhswp5c5CK+lbYz3WVU
qNsrrcripwzoxiImJCMsaDYP1i4mzF94EpQ0Tbseqw+VwMIJLxGNkaWrMs9woCiv
qC+cpzKVTLzrvb9o2sORUFBcv1q25nrJ/yLAPAy/Oo0SRmd4o+wTmXBdDarwPInd
BpW8j77S4vhxbrLC+4QJ7QzHYyED+h3MxhSUf4uZXlTCbBv9Gu6eL11S+WXr43q8
9XCgaNU4dzu19qqtZFjmq/ij6w2M8mFY+tDkZp6nExNpoEa88HNdGs+H3ylLZHsW
EN0HiBcvRuCqAbBrwYUv2enGv1zj3C5TamBN/td7nnXX5Urs04idzc+t8FvXQK+3
jku7ABtxwPlo2B5R1UmXPhyRXK/DTkOFi/kUsP4u5KcRwhw0sEcRg8lZMPYeFL1q
uqvydIiiHQPWw2q2IgbVV/uro1mzukA6jaha2ygLcZeibxJ4Qc1VT5AgxS3nA6C3
ntRbsyxenHBMrcDr7gXlnBaIiP121gwS2LMEvbkRxdiGlSNfNwi1xY0C9vkeMuiO
g7It61Cdj1k6OMVvNJ4fGhax+AFNA/l93BONXPUZDw7dIDOEJUYdN9tvkbKogwG2
zQm9wclK2ulIDMKVporWCyzAxpvRDlDqarWPnj0MIW7tvFoc9lS6f0KESVvJxvxr
icOPYXLwML1jEBUfU3U2SQ==
`protect END_PROTECTED
