`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4vxsrnYqbCENujUtwJizyW94fUs6Kw6LNs2h3Vmg56NY833uA4jI/2ve6PwuMmM3
ac6tOrMTMuAH7R+gbdktLd4wi9aZnwZoV3FJJ3qBSg/lAd1jIm6d3ISjiE+vV5fK
nPxltMbCcKBLpT8NRjYJNnBVi35QZyQ7J7BNQJB5EABUNkapQ6FNoHW0x15JyCTv
+X8NBDnljT7/6l/DBQqUKunnvcruzs75CGuKzrU4dVU0ryn700WVhui0O7F/xm0d
i1S6ZtTc71FNAX1eZRfU6jBCoqUsiCNE0/z4Zcufj9H/rmXhXINTlHL9dRGyMOR8
OPrKw3wkEId41bOOSFLOZDHrMwVm1A4gMj7RBkGkFNxPxMoAb8IqsHe8hVILBa29
fvmq+96kpbKRT3xQiJ+IlUMvsUFUR/tZnBbNIIIlOS0yDMXRQmbyFK/959w5yXOW
ujAzu+pZDHWAVm5dPF1nq6RdYKsfNYYwUEwPURRgnxGPpqFsW9YsRMcB4v0/OFpd
YmP2V+n8wzL2yIuk6Boy//Hc+sM1iuHu+lwLJ42dgioIUjwk4c40N5xGmZXcIi/t
IYJcTQ+v0rhIV5Tt6uDz/cjPjpOX0nTQVIOoRjU5H/pRk9AwPQ32/MIW8JXgARlP
TNJC6nqpDwdwXmR5uF1mo6Ovcg7Lm0rN3QFD935eDqXTWaN5ciNrVqLFiHy5bA5W
Rmq5+bqw9IQUZMf0nN+ZqRzHh3nP7cNP8xczn1Xlt55QBu6VnU6xL5WPueXGQQDR
hJaXIzgaUCA7J6lczPRfUAtVUORIHuTqEmIS1zWXnW7T3Q14vchV73BQ3EKg0NDI
USnez4+kRtUkQu7pG6tYLV+hdgbccXta6JB5ElDCHXOo1vEP959y/+ydBBoYsFMp
7FyiNPytmYgt0SH/M63e20L/Sj/7PcsTu8mZuSpjU2UzBTfvfzObJ835RoWnQbMl
i4p41wUUmIKvel7Vjxqp2g==
`protect END_PROTECTED
