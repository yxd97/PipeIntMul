`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VXPw89vGyLo21tT4LetxzU4kOWG+KQm8kW1Ygu3EfzX20EicqzCcn4TNAWgtS91t
hSGvQqudG7j/wK356HO+792BbdbbRFZb7iDHEl5/qg0kxw0GReU+jyubA6Bx1YWv
jc9BPBK1iQF7yHQsbAjditKrc9jeiBGdo2fv5Vhof1ikc051HhLLtGPxnoF55j1U
ffT2ynQ5aWLWOUainjHhXdLZ2bJam6XgRaQ7Bpe5rOnFDDLHsehTvhDg6FFQzpin
UnUusy+fhvITPG7NAXxXblB3eGTFobkOGeo5Va0qZ8ZlkqOxG1N1ouuWE6J/7o5g
T/UZ0+i8Qli4uT0VlsaiJ2MIp9A3878ckYviSGDhmBVokXJ8tCZf5IYwIfkxoJfZ
n5noSPQle2tPn+JGM1FqrwzmeSoDARemXNUexYIRXapWwC7VN6oCT6TSjRS5Z1Cz
d4wtkXAmyxkzfUhKdOPUKsybjEIpH1hnkPPBCGj9U4RsorC80uI9HXqX14vZSFEx
xyLDnqrBKUcx38gag1XBrUGfZxDKAjbg671rOVf4dciOKWqL1hRwQk7dgREUsaKq
a/gEkuObEoJWZ6w/vk7s/TWnWVZLh8Q4QOrzT3GwVlHJivqYGFYPnjyS8zbliv0e
2JYU5GnRXfZv6tcwr3RIBIzOxAk3GGpJKsZ6YfAVtw3wKgplwaoDrWpWqSO6Kaly
/6bG/9p36MUD5gy5TfN1yhSrDf+AciyxTEQiDU3FNPL+QtrWS50mgIqpVpqh6tDl
HHBQpaYqLNtEmp188CPjF4m4IYAJ3lT9fgvC5wY3SgfrqoTKo9kJIIrOFbpoXF2P
KdWEvhdIqJhRciH0jR3OytMxMYNNmWYWBuDIKp0X1sY=
`protect END_PROTECTED
