`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
75sgxljnQFkgue861Y1dXr7SsJcRi80AvOvUy0A/KRvgDncrLv06/AM6QmjpCSUD
/Gcg7qgehGFjSkYokTmRJdY1kLUWji9GZDvwPovB/0rrlDWC+IZ4BIGGHwfeNk/S
6mKKk6tFINmbKAjI+8PiTSSoF5/xG+Dx05sZ/UGXQ314ja0KmD1cssxrHqa23XcS
ii84o2CZnK3Y9A9zs0qX4sghadDSLoyYcvdj5bCrK1lL5fy/NEq6qM3OfPkLJpsB
//vYyqgZHGHXleI7C9qFlcV/GG/Z8L3qWhrHKiO81wWKQZBciqIEyv9GkLRO3Hc4
QrZhGGOWEREP/IKDIfcBKbuwkNvcVJ4vBToqwPWW7hkTeq4D0wEBHxuMeXcDEA5G
aFSVTqT0nCpqxrOx4Tme2oeaAL1cYsSZeRJvwnpSt3w2X+bUltn6JBgas0XjGO0I
IMe+qE116NFm3anCvHRR7+/sRXgBKtMEFIu6Bgb3a9ydz2sZdLmayInNvUiPTLbN
7eMqS+VMyItXQoFPsPyBgikIXUUrcxa2qVjpbSuo/knkHj6zdzYU5FD46C3xl/RU
8H+3UohW53wjNw6zcM1e3hq/Za1gKxQ32r4rQ1rVjnZkIEcJRGC/kVNTJwsfzzDQ
R+ikX9QPp/QPc9NT4vNqkyAaqeYNATZbFU4fnV/xmS7JATtMd1oAJ++F019Vk368
8hF6oHqWN6gql8Qu5mjU/XVT6OisnVkPgsZPxUlhvwTWifg/wrivhit05k5a3vY5
rTOqConInq8b0uD9NuNOb7oom72V/KtG+VRaZdasEy/iX87nlFrIjMoCv1en+oya
n7RZLubD19HSv7C7E4MmgIh3B++xNflybfkjP7z3q4wSBKghJH+wy+DYrn1IWENS
CJCchgLo7NG7D8WKkzPgecs8glzAoxzDEmg02PrCKl0jQbnWeYUeo5G9co5kR6/D
EqraoRqqjWJ7A7uBMln088JKUIuOvkDBR7p0j9hxJfxSSlqz7SB3lTfVAoGq0wqv
c0hUoXgCJSiaM+B7KJoE3wEMw9+91JDMtf8FUPPTUuf3xLRD7/Z9tSYsvvlFVpGk
5xayODRgYfHVRk1fknz6lxAqb7AFgPOW0xAKocd/9ZR8cpLo97ppmthfNA6t6bhF
/LSpuoZ9HeUXggbpAttcMkddnIlbUXHTu3fhjg4M0c6cX82U3eFERLcURnjUYErt
P3RNWc54+a6Cfv6mX3vEM+6hKUd8egLvMBj/SCT5+vH3sL4Do+tTgCrRe51nUhHL
zT5nvx9EyWuoRgr9FjzRZ4yKl9ogrFbMQpzQOKqJmn8Ga88UZZ9s6EdEXpFyWKSS
wXZ23TVebf1gGIoVrQZZXkaCekKqZpuVwo/Ut3dhG6XSuB0aYES+ABN642eOEzCR
E/0K07yXNnpIvq01jRGWdp5B0qG0v5I+QZ60Cl2cEiFCspsJfBHJCX9m7BmpLaZK
XosvAuObHXypfh5FdvdsqO21iTRgXiw228wBdxGoHGJxd46mDd7kQdPvTiCuxT59
+//Y3idq/1LydJQ4ApZuLfU5FSdxNmQjufVBKn6XHyu2ArMEUP2ZuX0l+h7ZDu41
V00PfM28fSkMzP1PBbXO+6jnoN4HuTUh04v9YOxSLCXjcjQ185wVjAhJz64luk7E
Gdg34ZFBLc2bGFC6VHHm6ItUEZryuHyeSXIbI3b9zsFDM84KQ7ylWRkeJ+Prkum5
WMGRUOUt18yrtErhCPFpF/42FhCWDxHC9JYNDJMIP+mZqiRhq1hAoeR/FSqi1dtU
cotHcE0tyS26A1kMCZlvLWMdv9CMAWb6HyuTrBmZtaNWW/O5GEVfeMm+mKlGhYKK
GYuCgjIgp730sk7dKCZHkjb5ETF0gG3/lb/4S89qhOfSiHhhmEJicQCqn8gofnuh
tbxB3hEfiIs4oeVbDEfFYlS1iYbZYDMOr7t1aEB7q7VcFkUBRZslz1bzoObTKr8L
tAg2n+o1cClKSQJw+hjracx/ixJ7SqJwLa6rPyKxjc89LrM77YasOeEfBkUC4RvG
e9/gMcqm29IgU6WA3DpNsaOy9cWuAQ0CzX+wYIdSepRV33A4jf9uVtuLeT6xekt4
nSylC54ch6d29fyfrR7ffvhn9jpPuJfsz7LQyzMVv90M4JPB5m+H1F1Qw1+lcUD4
WWvIaPfCVZDAdM6/bkVgyrEicwhh+aMmqsnCUDOaOHJL8rdWh/uX/nmckESiXeY+
Se9t1hCv273j4GT1HYOO4gZ4nROz+YOvo+zRgHZzYg8AX7gjc4jXyA0OZkWCb13D
UXw5wo5Fb3P63YARi8oa684UcG0epj/bZh+1yDmyOlZJf1+AsA2/CFu319wRGEIc
Xnkc0gXMJjXTtoVUsUl6G9EMo4INj4L3+8wNEs3nTkBO57omxG7kZoWjApLMzl7b
QbU2P40YTwIOSbGU/yJHKErJkQ5phxNOqdASfNy0nVO2LInjDUfCp8pW3ef4JbE2
eFLo7NeOMsiIInMjHilgp5kEX9GiR5MQz0b7Hjbs+4ZQSIbzuAAwcVLgVuBg6Hfz
4OpC7tWYG6lQUoLglIsK/a37ksOApwkRAwc2cEZrovZH8ONojuvGsNel4aJ57PXA
DauaGQhieyd4TbY2VuwYTWWTZcJ4rUBeYLKAby1VOoqWtNgQ//JlErtFe123AdQj
lK+l+e0SMHSZteIBec35WhqDxA99MzMAjGnIxxMz/e4SSyio5G6jW370CFCOrxZJ
wSjWBuMxjebZ2nlZxNQeTp6ZUa0q47F6WELZXJbpr9gKDkjwpya5FK+Ah05Nc2Uw
SmtO6uLH6JSF4olKOub17GX38dJMDD2Dh6kf3r7qzDLFiHNqQaPQnT6ehiedXAM3
RjsJ8Iwm6xhgAmOqtF9EK9q7Lzs0VDom5d3QMr3b6aoD7n7neaxP0CawuVQCajne
6Pcqd9Co1hsTJuggbeopvCmf52NIs8A6LbiUBIgUqZOmNh+fEhh+E1XR5hLKmMNK
cAg22NeRiQWw+bD9L4fwAmnOl+HA1DEkKJZb2zRr2xahWtTBgpI8KZiU9u8awxuW
lA+ByZk7X9SMqeJRVVVFMHmAjRd+hCYMHs0SS4Kev3IY2M3vpR24ASc8MAmF8KXy
M2tc1gh/8t5ZHY+kr/J6rtHtbtvz5IExkhu0a9y8QK/VNgjx7BWuWARsiPkpc4/X
0mg59JJ533fH5eV1TgvQJEFtdEJERkQ/388ioVfkHJm0rRF9Cy1DsD/BMFDl7DNy
MbREPsJjoLn27vCiULnkfUIlJvTgWlA/waICMl/mqxJRVXvKoHzgnpGtAzU4E66u
yL3tN/KLUr2138LwMLZyTd55k7Z1S9Y2KDTMt9XIiYMKQbLV/TypNhCrasBNzC81
LlgUsER/X2ZVebr1qW3UNndzdub/AR1zJpOoR/tkoWeXkJv2WnmausyW4SykV6vA
mOmvsgD3pU6kr4JnUlF1mXHMLi7fOJ4xvruSD6CFokKTycZl2JL3JiSjr2kX35qb
hR0nuon4Fn/kRgEhuAYjnDAkjWpYzVuUQhB2wiCDOgM6se1sXX0/QfEnHDTjagg+
2RosveDgnHiRGEH5UdF3tb/RW7wWKhiltgM6kSEQqijwxZQeZNdM10LbpdkooQRc
QM27M64BwbGg6bRTxxW3dLRw9YDL7dyydr7X/LRFqRDQqqnBI7K+GkT99qjWBmmw
O0iRfCf4ZilPfW9BLrWXMMSMwp5Yj4vgIza2OcWK6a/9vOyKa8qKoxv3/RgN8mNf
FvBsczQ9eB7NTMULPA8MwiyK9osXwBj1pHEAlrpczoT1SIy6rQiDE4adT8RqwX7c
VqM9U7dvP+4vf0AwOT+mk1JgI5bITS/8fhkfwXlxdDuBotDFsVNsfD5CrxM7zI57
m3U49AK5dYlB1NXMVF0mIvkAiy8zQFnd50Y6myZa3qQQiKfIMQ06WhgWqKn/lB7K
KNCUO4CDuOLNR2/XZ96DamncwERgNREprJZwCe2sCwNQtJyqgMSgflsZTZwV+H7S
syLWE83XpyRy8h1lw3mrPW8sUZ3F6fh+YQhnd38heg/Tzd2swhiXsel6YzxXwjRV
JOy6spcF+uxWjuewiliVuyhGRbmyKL4LLKHAdAuuRUHSl3CYYdikpipfOCxkpU6D
4DgRRVACx7t/04tBm+LGbx4oqlKZekRdFFzumXpk9CLHBxayTxRTgGJM3EM7XcFF
+kW7Gyw6NtqQzrQl4n/ABq1mqa8KpyGEzwsClMnn0VjBluemDqATpkOz5gMkbxGy
mmEt0BEtaNDf8K8c+js/LBtlV3I9PSWi60D8pMbdB3ivgnS4rLhh/ly/MUilOExg
pKvZVAtDjdyaTAUY0kTgLRgm6o27rroIc6TJsyuAVEyPI1nF3MtVdGNqFVkjzpE6
0m9TKhzjkuBQHNHjM+HU9p8lbQquM2sWT+MIcgivPpdMxmKlRLi+Q5+BCO37YXom
hmzYefxguoSMq4S5jsvbuy3EFHsMttFQSwp+Kc+L6r1Xovjs4mEXw0Azvjw0gxwO
nAtkcFUJI4f1DB+NQUeao3eNuEO7BQo0KrNbZ8UVQUN+E4cxebK56GnBnRxqmvKk
nXev4SlW188wc0Fr8sniwch0NXgAGzDvQIN1OwEgr+/1eBg8D3j2W8FX5CTwlEv3
tift9NG9k0PDbRpxvQKUb7t3onh4qODr7+KfwJ54LH72b3e6SiD/QIr20lioRUG5
P60UfFx85ZPFG/8/VxTcFCnvf1wxlw9xsHuobE6yVfN9QEWSYGvJYrsiFY4a3YII
n+H6i20BcfrJm5HlbvO0le5s9jIwoQO3OSoo7qAlsN2MfdQkjYhiZLCjhVTWfC5x
ylZrOBRexjah3CeoftrOTxPu6p1PmYfG5AP5lmBK4noxIgUixbd8rZQ/fxqy6RyN
1aGQB4zS78Nd9V9Npi05kPROxEaOBGQ2i5QpQf0MLe8iq1AlPJWAYD6SZjebmZSa
3QuN1AHriKwxfWl7ie+hlylwhRqLmxmOu78k1Vr2sNszn9dLQNRQe5T0fYFnSoxe
kplmw3LVEDiGbuFQ5wwqXbfmGFjReDYj1tZFQe15WtzsBPA+1VXJO2yY/o9SbkMS
efnSOu3CeLKvHdTynIO+ATyIvC/wIDUoRDhH9hs2CIH16lSqnsfddZ8X/rDAdrql
T8bT6x8EDmikNZI+Dj+DhtdoOLYoUFJ3OjKPsFXk4ap4gkA6YCyoTsHnvstbE11Z
31oEYdDYZwcezNu65DzKiaDP50fb7i6xcJNYrGNgQb4Bn2aX4AYUrodg2kF/6jIB
62/OUIWcBNcilCtgtW2mcHW6PcaRm2V2urg4igdwSHiJz78U+MGg3O7uuI8Vmpfe
zH9xhAgVVySNWtzPdDBbhasYRK1c4qDX/5aTmu3fbmy7TZiBPw0jq0S3sdMQOxSY
iWVcXkh0Fx85/FHhbWpZnmf9VvsKoV4ZQMmQzZYBEaCW+7o/Jpz3AIIh0ywiRnIg
LTLV7KpfTwIoTzJVbNliBHiSvHWU2SlzRWkRaKO7O+GUctE7j+pF6Mc/buIhFDSz
KVkZ3CsI074SuM5JtYZz7y/R/99Deqb4EydQMpBaXwaZhuE1xyB4onCxUyqJ4VdZ
/D2eYAvBN5b1zyy7XHe9NpdEfAst7yKMxdZB6CLn4nH9sImzdy4/8ntFUd6duF6L
TiSeye4Fc7KWsIlhxYyf89F68EWfm7HLayZQL9bucO4rdkHjd3/H+Dwo5cHVNEYj
hiAD3eLoXxBhMv8+/KYQ7OBcM//7rdnEACtqK47zbLDw0o14jm6fnM1jhmiAxIl9
5ctBcQFrND5gGc1hbLzbbiR2hZYRebWKj31TFnAXiBzDg7D6gwJzNSwpVKuHJBw3
8lpgrF/qoUkkObfEnNJbq1HhnV7B7YQjWg1xdfaPioZCFtw4FEQ2Vh3i2kG0t3cZ
LIsjmSdOOsc+vzcC+8DRcBLihX3c6gkhsgByJXb+qt9hXTNlS6/MocSGQaBmy7xd
IaId/Ymb0zdGFBaohb+6VvEIhSiz3QQpcCPpZamMflRtLoYf6FqTJFiQ6uwwxPQn
iLhZ1IIjWjAaIBfLpdAIuOwWBqk+BGVJ1n/NZcuvpx8PJH9X304MOKwI9bBn11+e
QFSbVL+e6KGbgyOrMmv+os1xN+vlYT/WdEBkpINsldHA403+hYCzoFR0nz4fjqm1
XVFems0ArKyn5vWJt8CABgejEHsHmIhHxDI9iTnW1wtqqG/zeX+WhX6jv2VoMU1T
2qi7jchP8/vTs8a8a2XywTyJSiXdqh0tHTC5MwhK54zgyzDkAhi9TO3bCsxPdVsS
dMJaNkKeBeSgLF5XbnDuSazg6ROrBV1yBzcAL4gUewASJQUWLQzzzTpt5A2qvoiq
BHd1SBVYMbaHerCCQI8jYGxXRKJZssIT75cDELtSIIgkWQXJQI2MKhunQLXTzzXg
zaXxPeQf+20vKd7DZp1VxNo2uto43a0pAO6kGLJJEZVbQNOd3JPurxK+DHFxbBQp
Te+xeR6tZhhXVCJxESX5yL4dc0cmlEUOw/kCcmO8ziSemWFS4RDaBiZiDao4+jv/
+tICH9DFEmfxo016PAdIO5Cl0pluPWvHVPQ54TtHxbwV7hnGgs1KN5NenMI7zFyl
CW35GL+ffn+aftQY7hlJVcydQ1WtZ+Ul83nsRMKbQohO1nCdv8ZNe45zs1IweT0M
mpfl82yqGlEI9LhZ4MaAdWdJOmlFwG/vMnAqZ2c4gS43CxpVdlnrnZY06fdX9NHs
BOftSu5K5UzRIG098GSL1TF5UhRjG8xOJ0N2uA82ydR+XLtRzq8FsDg+O/n5EDPz
l60kpfWIvGTS6gcSgyozWlbQBnX0dFS5SV8uhDvh2ngvz60mLAptMtDBd6PrzIVB
dav5cvxdYacBZRDOnUvN5EICrHjhZ23tlrISDh/mmbQrQAW9FmkW51u2F7GBwVVP
LD8szKOdm5Le/XAiN4l3cueH2fL70aQ0YY6myo5ualEGepEP8bA8F9gRI8rzg3D+
QjF6woBYYXYVWLQ8x1l6JKkfpwwRIbglYS2nUpRz/e3nkkyK1EmJWfZpiavdP3bT
X/3qc7xJbJ9DBfNU8gkcdf3yi3sDSOL9aZC7kGD6om1gkBcPDX0fMe0MmMpmLle5
sMbMRjrqlYNVGZrAEDjJb9TiGxqZbTtsQrzvNeKunyugWRE4S/gz6eL/jTEC6d7J
S3qTM0Y779vzg4MlUFGRBHOcKM2eryaMLhZESyV0Flr9dwxKBWxi1oIWTnc08Enz
2PskFmAlLJ1GHbXECPBb0t+c9PQ9y+5ReFE8HC/J5avTBRJAJGx3IRbQZ0t+IwEZ
ZOuzJpe+EjEw7OdwBt0APRU9j2XLcMdmzshRr8FXycGP9S2KrWDQam5v7bKTLkiX
8w4Yr2mI7nO67atVWfIaMBurqgQ8cQmJtx5qM6R1qG2+EYFR79/Irbl1PjDUMqFz
dRbbI4MOrIb5iY5zWoSqLqYcNYC0TP+5OjM5zXifCitMFV5Pw9FXrw2qWVme0H+W
BZQ9+7yIzbgXl53uEzywugXO5jj8vzyfWbXB1JSoOw3w/4PACXU43euEC5eqbmPM
jo+3JgSqQ60xBkXPWg74IZxxcwaovYNvTnkE+Nrw6oRMJgeq9nxIvdtXjt81p++N
lJD0Sn2S+MRYIJ+EEtqUAimSKCdYaExhZddfjNJOYccBmtTvZfBt/Ho4ZkmDoe8k
6fEf+ZXMogJoDUo2PsvPCz7vphag6MEpGTU86RlI/8VyQf8Ob4LSYdPciERSMsmh
psgQW/w8g3KfLCdUqY30X9PtndLqIo+ZXa25/gB06R0fofzoxcjXRPMovCBl+VoQ
8g/mqD8s4Q01zozrbhrEuKktHVwLZ6ELUShmH1niVw3O+VUrtqqyZ0gZdo3SZgz4
Wnrdo8UthosHTclw9fwMhksiv43oFd+g3+DGwlf2XftpB4d17XhtHFndcRSu34M4
+J0eC7q14HvnV3MpsM1td/itO0OVfwH1aIIhnAlVjLHglIPZ0NhZHLCdwejlb+9h
iNjEjnpkoTHRI+k1fbNiZF7gTeSm5rPDbSmXq61TxoSr1ag725DplnO4vvWY5kPP
Bk14BFRbFXIH21HwTX1/E1KFdcRNusLVsLlpiuuie7fp983nIqzhL4KbjrfXEQle
pY8KliBj1NyyI93/J+LLM5CbSba2NUYGhbf10GWpg7MQzBDr4swZLHnoGYZQZt6a
pCSzi0/uQXyPrx5H1C7wj3yj9Zb1JHz8lm5iOokOaqMvUgmAdVyW/OB0bmiVHLNC
iN41Mm4fD36ShX0k0wVPF1b7uSqW1Bo6n5arWAJwKniacp6QbYjKYTTWhZCJWjOk
Er4yB61p8OykLiDSgkuCP3P9rSqwPPv+jZsGYlZvvKLEjGxUM8Mx+sDjpQF3p6YX
UwWVh3EInS9DdsjnG4JFse6kXliEAlmheQRX2aLCkdCjzVpvRfi6NMNJvvUpARvZ
CHWSYIyoyG9PfcoOFFf8VaGYintWli5kn9x64R3Z0/buPHApMifgKTFIjN4AdK5O
xd0fm8jcQCGJCqIifg+/aIXXj8i175fxLjAmK1LBwa8jrjpCmsLDy0cFac6QnTWv
tQYnhBUzCGGacDEbwS8DrfhCWaI0h2pmMbgINUuZqgoXgCSFwLxeWSEkt04QJLLE
4Hvdbu8gVLctaF/FTkSsqLv//4v2b9hRnRAi0rb52OM/WNiGmoOR8XRaTEyT9Jnt
d1v+9JdbT+HOUP0QxkXWxIUNy0V7Sl5LmYW8Lq5Q6oU8bQqBCBRlabG3ZoGZDbcP
CNtoV1VeHOTwOoT/m28NpTeanLms8GX+tHCFigD4/rg6GtuI21lzwPhxSN90ZrA0
y97v2R+OsSXatTlPPsUTb1ib83yRM8GTL8m8jChvAroZrO3zCGxbQiG7xzjTG0W6
upZNpmKZJYmckgEOw6MwBJHsSq0zgBkRlMJLdekCfUT8J1fjIhbOCyvBwmj2T80D
+ChC9CbOuL8UmJDfu13ByYrpV8k5vAutho0PXEak7MCA/P483xoUs37UFtNSaFoi
Ktlm52h0D8NYWxC1mrKjwqgwI0cBGiy3agTkrszmIrkgFayQwMAs6dE8uPJXoWGp
GsxYeYK4RETT7FRpSwzSgYF0kQVO8CSnWBeQGyyGrIx+1JH7/G4He/R9050h0IWo
H8WbbxR73dK2MgKyZh3Ovli0tWUsmvJ13ueBS3bFtn7nfiiiRHNPFoNK1/w0n2jE
4FsMbh/UN14XScGA7+vs6cSmGrpfIl4+aU+h9biBy5K30K1FNjYdXSRORzO1HmJW
6NFUfp5FUx1b5S420Dq5lNzxI+ZwDIA7wusmyE12wo2dx09IhpK4e9jO5mVM7RWJ
/5GXgs7zVq5MpZ00ZS/eNsegKYdEHfk38jtOEgJlh3pQtj7ouDAX8uD84ibmb2Xx
Z+JQ0DBm+TtCuG2f1hdDfQNSlisd0nlGUt2iDFsfSadl1MrxMV1IKsZy7aRPo0Lv
KI60B7LB+sLMjBGWQat2H9HpvQPTC4kO6GpSCiO93MET8EAIEA7HBcuR/DULiBV3
ubt1HesFrPOjLGZ5dlBFvgQXbAPhcFF9OlxQVrlX/JOmsaRExVHWDw3rAz4NlB+y
S83+tClj3enGX+d0mmcqRYiiifQFCBca6HtHPVuvu6DRB34dXKS+zEJpNgCQLM+S
APme+jCesm4WaAv0q+sw/w2sCGP4ovK5jMgZ1isONKu9cRfNGdiyBYLzWacx4Ijt
p1Z+24MHftBJQPTKqYXZnKukEAVhxrcggDadhXVlzun0sFMvmfcdEOnvPbCxwO/f
eElG9T4W9UNmxhvemM5hKIsrX2+LhPDg2XWEA2sQNC+PV7qTzLYFkGxRk9S9u1i5
dxomIFgcGE/dEpk1YoZolLhCGp01tSxsDqXP+BPendFLRuTn454MYA0Ilvf4vJjR
MR9AtpSBI/9GLFG6myZ9zPDC33TII5I3+3qdxu/X0UkINYnj4VM+zX2sfBioZ5cW
8r59XXkP2MnikiLRrbdg++q5VOXQ05GBfe7Rg/JJ0XxCYAwsGJ0ODLV8+tNjSsMc
clqZPc96cxJhqoSYtyGUBIlI1azdBWB1xUr/Ug8XBtkvr1w2Y8Bb5h9/hm64CxQZ
1IllY2NjbvXsudrB6jFudfQxtIO1zI5FT7Xvrb2v6LswuOSDjXsmvUuJ9hZ9bmgJ
TbNVWJjGVMvm7/AEte+yy6Od+92fId7dgeyeZv6ewJCs2K6wolFY9IE74s07GuYs
hpfmLPyssima8FBKt77y0Oz8AmO+w0GkRIPV9lqa3l0TKMmQ42WsZu1MRU8KPqQM
XYyYjMpIMx8FjWHyBgAm+BnicoXphygVXfeIse7+sYMpl4p2mIW//2CeeGxfLI1V
eADzCZt6SXn99SsfFZKt0eW8CHomITzu7Ki3GHPMM2uVbrvXZI/JukhondEADzh/
Cz3YXtvc04106gHRel8iRAsZXVi2u77A0w5hDNny0mk7+OAqPO3lXzpSQ+FhbJXs
xqQPV1d4RnyFPtgabPRyVzhkJMDZB/maSyXpreOCVC70v9JlFxUlPLhqk8QOmzac
FK2OLRZkRuspVK7dGs5n93xIA8aHIge681dOqUJ0U8QEFIWA9Wc7oSCQfrAtDIh4
maGteKrajgkRPjz14WJRhnxg4EWMl6j0SnWPPpQAVGtUaJCvghXQ52Z3nlArdco6
VbMiqlZ8QzUxu9ju+qnt/m4uzOycn6PXJxlEQldVTzs=
`protect END_PROTECTED
