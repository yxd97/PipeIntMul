`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fjytMGhVOfRtFF59gN46/yIqx/+MVMKMDIWP75rL6EiHKq4XsCieLs2zZI+ektI1
HMekb47OPwIIudwGfHqPpYjEwEwTvHkAHhTA3q+shDfWFM0J6PYxMVw4I4rsFKLL
ozl8UP8LkBwRJ3710lv3UsxlKu83c2FVlBmQjsJpDN/3OnSVOXEgOBXjjtxFgxM1
7dY6OMvBzC3Bt/LKEF+arwCG868vUQFSCFOcaODX7FOa6rT5DOOh0Svoi6D1ZNXc
kZA6IVSLienZto75YLNGFvZYELZxooGIVkkmwqVSc4UFyuQvynF0sW2WlKthJ9vm
QZYcgPJWeZW2hL5O+LcppddPotn6IgwNhVEurteAj037K7tRjWQsUtKMMf7SoeM1
o1oknnRFR4nclsFNTkv69FXW7mkXnCa6AHcmrrFZ8xKhAt+PMmK3FcV74Pmk1pyS
ICRaS5rJIIhGjJSWV7CbtBXpA9JRyqH+oeWIIa7E0cE1pw5HYwpKsD789cqUiHb3
jScGJjvRjEy4ZHXxJ8tjI0M7G/dn+BFsRPS36qfBhddsKl2OV45ZDo3sjfBWPiSc
ouOGRseug9M/HknkWITVmoElUlaGmKWPH4DRhKO1kkYjNeSSuHbMzerRNIvpXCOc
hsrUDGz7EnYmAomwViOlpyVN36afIpu6AHygWTcIrQ5DP4CgjVvF9xny4HVDifsP
akyLCzTaaxZe2akCt3XRUO89/944rhCOzJaH61q52dUPGXpBHHAhQgry9dXq1mjr
C+3TGKG6fY9lldoAmw+i5oDd45H1bA6m9CMTzTBgWLDgq4iBQ6tGAbl3P+S6OTRP
enm7qsoQAREhdVT6RJqoIr/phnahY4Iwmj0nKv5Qtgzj2xsID7ExwSS9C7JcSTcJ
DeoFQDfdc7O+Kvcvvsxp3Of0xEHdxkeFVGh0rblP0O9vAi0psqd6GXPo6yAXsigH
wBoxG1Rzcs/DGfQ6+swGNkmIS1n9IbUbs6EEaxdsZ/bufKKq+SqD1C+W3wRxdlXD
nPfDEzlj3h7m1GGQ46ilHDVt5djrAK3AzPtqfcAkLRI7qJET9aYfaVUE/fiS1CfZ
QkBhX7cVnjlNm8NyvvW0u6dSpu6NgZcPFPZytKsI21n3AAw4Vt41/2djI4CvA+tk
1haVXwiP9br2iiV6r3vQ3hi0vBqCnY10uNy82WbjqUqHmmyG3tmVD7HZnqBdZqxP
laXeakN4iZZALCStdBUmWgZ9dz1M90kHMTaB4P91R8mgLEB+XUNvqWlX2M0t1VD1
PRqZ6QHWxrJpVok/nOgSBOivS6wiSQWrXaVKG/GVwx1lAe0KRD/RNSeU3m9zY5iZ
f5pvBIs/HmVM9uzQEY2+AZUkDpw5h6ft4joDYHPG99AxVuET43N+EKDGl4ohh0Ga
Fjl/+LQ0KqKPk7hIKv3ZgNzZEuqfY31oFznRNCfU3vqdP7Fa/HoxGep9Iki5lVsG
s/ODmkEe/PEM9kjxZ0aFi+Yr5vyoWGkf7dE05pXeUiycPc/NlsCF/7P7vUdCmQiO
kEK69MbSo80N0E9zIx9dE7IePtCqoCqBM8rjgsIqSHFZEzCb2KuKYU2cgNh6YpD6
MrtRijfCP/Ep2ttG8Tm0sChgKyehXuBQSyYcOqzqELo4/axinDcodf8xsTlCrhjH
S82IL5UyaprAnaIaqgcuqdnhRq8eCM9jdDr+lWmo5d4GgA/rSB7U6IIC2OnBK3w4
7/7GMMdLHN31EP71149qSzz21Ubgs08DgtRMs+9657Q+ZL1Hf0nLeTuHgcyq81ru
UwpHre0Rsko00s1yah7bcrkKRNaf7l9azfXrgHHf+KUK7e/03AL4N4j4YlaMjV2e
vfhaQsnZfItduVaYAlInOA==
`protect END_PROTECTED
