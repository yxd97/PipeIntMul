`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C19qKKhoirzrRAgS9h6Z8fQhVtk902IcTVcgMJ4BWevAhFM6Da52v/+PZ1w+deIr
uTmHg6mH5fAA/vz84gxPeFMSUGlIVjzkRSN08fDzn0r5lk4PEM1S4J/L9WyF+A2z
OAkc7lUPMURwURwckr2KxaqQHKotlHgeU75ZQ127EE8MNO150qMS24QryrNc4FmG
+kwBRlOrDuMXVoYd/7Hip8UKAzA6WJz4D73oFlE2xUFmndW/AzL4uOs8IsBQdMz2
/nyGLvKLVFuEl8dmCzKqJ5LEQ1C5OWnLAAx0d+rznajPLc291lBTCj1yg45ds5wI
uklVKCzQu8av35dmDXFhBAcTg9MPVPhHTxQkyrmfm62oUBXHoPUSlfCo+MYNLeBF
nxAZZZ+ttA42IVWhFiKcckXXu1Z9ZzodY0F09u0ils+tDVNAGaIoF0P2e6ei2knl
NdeS2CHbai4iB1Flf/sKJj0aKjt3SP5mrqTdtxJUolLo7O39i61KCTEkp+DlVKR0
Q1wnSGrWG6VSNgm3RqWIW+Mfi6GNBGw3uRfMSAfWN743nyAH3TJY++euBq5JlelK
iZxhk4TF3LcjahxpoJH4aNazVw9/7m3CMwV70ZgAVHVyexHhQ8oVf8HNyneErnpu
dTcMA722+NZogHnud/O+17EDMWum/oE84ZwaQIqoJ9u4vV++QL8mQYflEiHSMY+5
vIiK5Pd+8xrmwut5P3OvUbcqCG/dEDHF7FRpUtcvQf61MGqFpZnvssV7Mi+xuRey
2rtf+gXTQW/caRioZ6sgllAUTg44UMws/vdeFtR5B2kXIVms4/G3w9sMv2yDNeTU
v2CeM3sVKhI6Hue/trCj3isa244fJ2ScyfdjlabZXAvWZtrU9KBAAXQBvMHLjA54
JJ059gTMNU4QwdbWPSZkvjBMHKnVAeS0UxVQdVSZftMgIiyK4kNqIuimAEMZoHzq
sZUpaH5BRICwFuPO5W9dQnG1QvR/NcXb/Z8SPURjUUh7RA81BZs8LUQkeYcn45Sf
1NsLWp46gtTwFINq+vnzxb+cOVlemCBeOi1tpxfv+/cYDIfQ2uFI+iVZEcCBGuWC
Yzy2/lvGs3auqt7Itq5lpL7Z57geud43UMSel3NSgZpXnSBC8t5+rg30MDOAA2M4
fCuaKTuMBky1OVRzPpR/+UxwJ2fwVqogsuXtxyoOx17rl7iOUFfjGemTfz9oRFZr
dGW7kPYuH/wWbTmy8YsBN8QuaDEIMoR6VDZydNNZP+sb/XNzd7Z8V5yYFGRuOPdJ
a/u7jR62aIBIGBjE+6rNPYUktKUUnawNn1xGUJfgKplMr1jopdLFKW9/dpFxa0vC
NIHEh18Rw9imebJkhAGI8rvTkSBzrGVJAYVkRBKc1M+xLM7QgCqDYENFwWIbG08w
4opG0eOWCKlozVOpC9Dyb85+q+KPG2Hef9aJSoCs7b4MzgV7TIciwpM7bzySE1h0
bWZoMOWCNbKJnShK1N2xWvgpV6mIcDfi35WuGGKgFrbLTIF9MENizVCgr3eHAQRw
1SCCIiHChd5fQwSeC7Hb0GlX4YZONWni1zaAJB0IAC2ZC5Ppf8WoDk4N1+IpZHBr
Fytlfkai4+5+bs2CHcxWehPWA+r4439GH9BFgaQi15KWozmGqV364tYhnS3DyI2t
Q6MDpM9ejG41+qLoDZs9z4QlPm3y2EYrlp1FJ3CzBqAfV+izZWmIdK2i7ZqW2VyM
FBVMgihpV+zTEhWdQYlwDnTVl50RD5ejHDniX2gQM+s8pa+4aHK7ij7zfppHrJTR
GxWFZvJETX03pxaHSr0afkfJNvHVdaHrStbJ5rGq/PzI9SikC+v29wP55Xm6Xcdg
jw83ysFXJDm2Wm7xd8iW422PYx+/tcgTO2Klf4exCynj6HHsFRNETO+vCVH5tHAL
2dSlP2+nhIC1PbgT2o3yQZWWoDiuA0CjT8u1lcwq3olZmrxzP1OV65wVp39kWVD7
n3kQdhMouHKQepL2XBQb3+nTX4Wf8j0usJWX8Ys2tionY24OtzW6bYyKWoJKgMbj
Ryu/0RDMeTJf9DAPM2pfmcM4WtG91bW8tYJHJwovitTQoQMCwALzgr6fliBpBx10
x7MZWAfrPGMLyDB0OyKjyOECD1TSfIX7eO5CNz2HrOS/EQhwMLtBt5GT9VoIQvFa
O3Y4prx8WLek5pWdS8nOTrnfx2wIqfzzw/MwubRarWFc3GFGiB6P47rk01vuA/Uz
cCa7rvYjMHBE2i13BabWknFSWiHk1QWgPqy7RpF55LAQ9WaNzQPagQH1OrbG574o
+YcqQXe6ECGWdwBZ69GeocKXUuDaQ7lA0e0NIA0ezy8s3bC/6bpdpzu42njYAmHv
9nIH86ufo0dka7jTTPSL3YElgw5arPKYfC1B9gVjz06IhVTOElHZpheUcesaJh9a
XkvzPYeIHSdB/oKiGrqwPiOqoxcQQYzbj9iQMnxtufccoQ3/unS4b+Xgd5kBNCPH
H2xMVOABnYvJ4pjMikIksQ==
`protect END_PROTECTED
