`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DrRhtkMeu/qDQ7kpuIxbli+1Jnk17rV+QyE7hd7pqwe7EXveCHl8pvXYNVy0kFdX
+9WrhiGFStKGYMrD8Tj5NwnYYS8p5ZYm780BBEupq4NZu/UcVt0yA2nMjeq99Yal
NV+82Zmpmtq3xrJk9j4xeAtKyASY5d47YT8zW7R98LUvYFSd9izawhteZs3CV86s
tkwVBkIak5PkMVlt1SEjVUpQW2Bu+oxI6/48KbKDz3yAd8rF5UVYw0CP+vv9ze5q
PFf5dopxlmoAnzcYywuh3yUcabXuQ3QywL7hHHRcw0b/3hnuydEuUFmSc2fTKHV8
Hvm47dE7yEWeQ5GQl5JtApWfnZIuBU613+ctLNCTcamaY8ZwJA9QVMgQZglRDnDN
aep8QvwE2y8cs34myxQH9ww3eRHQodm4+wRd5w9P5RR0SG1B3g964JQ+lhpkhjMa
0oqLeGBidRX1UGKowLAYeZIS0C0Mu65bwc9amC+iWP8OwznSQeXXsNuGigz9qIvE
u+0fpu13Kn7qzU371LUGxheQdrgJNZY+aCOukwTI8D+L1QMLmXk2QyQ6sN76H3+i
HuKYkS0ZVtB1FJFBRfLyPitoOVviqT7kva1/EpjFaLsaswi/pod5LAovep3JHvNh
xup81POUfQ3gw1VtSgF9DjWuXF5FmKYXazG754EPrFp/lmX/w42I2l+okbNU330L
C8nzT+wmM8ho8c+PZ4P8KRSoMxSEOyPvaV2KdPF3yAY3/SyxbUk+DtLpLyIvYA/f
w87rh8Ygx2jglRoPu4clKGK8o0N0GOdFdwTWYbta4Pjts0CajSv+UPFxvKpFfjjI
ubST3tPYncdk3BMTOW77XQ==
`protect END_PROTECTED
