`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2C5lFN9hLd5Y6mqcH1fPfkhgM1f7sh2SUWO9hng+ot+zLlfcNDdnI9+REKmMWLmu
EXkJ1LEOhvu1fuNTvWltxBVovkUy9YyBrY39jZ/oo5cKDfW/JXtyiCZRgmKgxDtI
FW25fM6DI8zPrOz3XGu2UjgxE+ooozoJ2cekcHE1OZ1zsCyVsUJUCMfg3DOIeoyg
XUTz7KGM73cQqKwQk+7OvBnETdMHhCHaZ9RRo/zK7x1cJuln4HJN21ZW3XUB9xt5
8/YkNZMlnpcOdPLb6OXPCSZUpu1SW4jUJmBdE79SL6/qpddP57VEslGJoljdEzjC
1A+PhtZrGhGEtlp9nLNx3w5dx99LjVfEjPGRjuw47Xiyd9bqXcU0F/KidiZMmgrp
kAVrVyzP6QcJgBl42L0TKvsJN9+uS/1Q7144l1fh8eyC9xSDpLUm7qmrAz/LHk21
k+sJhV8V5CVMu5SkzLnIVdR5J6cVncdCIZkvVvPwtXOlv9dguTeXSP4SzotxUmGd
LZ6zkxoSpQWCqOuYSkvhnThe42bEjtGMdAJvqKRmjmVNeTWJoWjXq3KSkGqNEx/d
jwEvvMHN9d1KVXIOgizlyMgklvIUnKSbg6Vh+PcLejOwjnH9tCn+PPHHlqGgmZBv
FuRBB6z6QFeSBGyP216xJON3cGDbcthxT22dxEGDsonrm11GoO5p706XI/yjwr5j
oB4TgS2GtFOJFPy4x4nHwJnoWSULGiPxCpcFdzGrQjVmtu4zAVDspgZH/TjOh1Sf
O0HKn458cObGgpyPX+e1MGnA7YPFG6IbaQt520kbdTVthuaILddg3SbiAuqDtU5n
y8r27BZlG8rZN7dt9R1UJ2QQpzCE+92WZ+d59uub+xzyv4turE/EgJdtiug9YIzk
aYPj5Hik7Hw/tYkInlY9OmUVn6eCg4PxJPlMTZHK35F4eLn6KGr8jCDW9TncCJM8
KhzSZkUzNjbJgm8X3rgP1gLTpQn7StfsTFBnqeKx398OizzqOtm43Ft5LAVyrikD
wN5wCiNoPpJsYJh9MdJ642aXlvJe+50Sn/VjAg92T1FvcT5373kNPV8Od4B5Oj9j
5IZlVlkwGZTlC2FWJviT1AsOp7ghpVZqebdkUcRTfShbihGS0aVJozGdYAFxW8Gv
AtPzKLi526krVTb43drBmUhkxOqcbwCf2lhf9SEUPvquGd64mtcMSzx7yW17ry3P
rXZraC2fyP3JRjHctquw2S8ZI9guj8wL8RW0xIgBs3N0RssBQ5eO1MBm+MLnr5Zq
C7eMKvII9+0nW1W9dmVspxydDXfJfszBaa2vPRh+M6F2icrKrHQd/TOP1WGge46+
6xYBJXwN3UVXYrWo53gyivWVyiMD6P5EpijAfC7zTBeoAJl+Sz88vwo/AuYg87zI
QCsZrmGgnu4Z5SVqS59gU+TPfm6BuV+1k+u7D2dfniEFxGGNzt5mMnKj1k+Ysbe+
bzwNCWcxbPX8U8X/Aung34ZrhQEQVHxym9b14Ld55uAvvkp/roRQBPWRKX1fK3N7
tCrly9UXc8g80ZqY/LxsNNwFNTfqgYJYTFC/W6/OyPP2GLC0dr3Cr2YzaptOgHQF
yBfGHn1gRcA5Sdg+LQ3flcBTQeGRF99npeq7yssEAvAJf7QMBWUe+jMMx0yUhkOM
zNS7N8BPc2QjT3IvNeFawEyUj0LBQGUS7+x5aMUeS0tmZjDQ7PjdayLoo3AfP6M3
r7KPOqqPnIvY72eFWf7FFYOG86crN5vLo1PI6iLJ/yJ1VfpJ+OdZJMNiDIm7sCSi
WOwMoaiLHKZPjawJiOHAhrzZT/YyJdvrJHclgJgmF3onjel1IgJaJm95pUPNROfZ
hMUt520S06aOhSyjCxQLSo7KRPbqzNGIwOc6oFhn281Rv2ooaBefRWQ5tFlMQ6PA
2XiytOJEkWravQzOMBetV4iNNZL8TFLSR+fSvxuJdDrhYUrZS4AYaDnSnKGlz0Pt
no+THPZzxSbZe3rONU3GJHb9Erg9bypHWRZtQiWAYVq7d0jnplttF+E/nBZGFPFh
ttJ8hX3AX8TLfg4DtKZstYPUjpDYC6JAk8HHG2imH+qTJssc0REks2CD2HomTodJ
khiwZuLW/6kL+O+jNut/DDkh4vdlLsKNZV0g5GiCW7c=
`protect END_PROTECTED
