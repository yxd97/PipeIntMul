`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f7zW6FbbtfSgd+fqWwLDvY/W2SZZyThaA5qTZcq8jBE//opv6b8g23HYFVRaqpiN
5Jqt3lUr034BjlzBybacjpcgT3s+G0SGDPOC493pyT3VHMfZLbJhoExjdDbfkCM3
tlgN2qUdaGKel5Lf3zpU3NCAXIim9nAaORSZegsfXChh7xzr6kZ2fU7o/36h+svS
bM64Schb8yY7oribuYmsb3y7jS3UDoshGNK7zVxNzWmVrxCwcG7CzTGf84zGFUfp
sJ86g1QeLvwkAvoAOShLVyF3OKQvmoFDUCbNhKNbVlelSeKjtdGGB9dZTGehEx6v
ofTVDC25zAMIw+fIJ+fHauyzlc9Ea1ZeO3BvnpHM9ztj6rfRJ++49nMnnWIK6QuU
dAObIbiz+EaBvjRG1ZbZKQxSraI45NG7gP3dRKl4aCupy8u5Oa11ys4ggkfxlLyi
`protect END_PROTECTED
