`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XXpMuGN01OhWw1exZr6JFRNSaPqdTLMYgTRs85wXG/GrnqxwBfnVlIeB3yqW1+KG
oBexI1heE77cfTK7qUYNk013uGwFlaDnc7E+ju+P9v6lkvo4lUt8jd+IEmtKtf4O
BkLcfc+UsDRApPCKHKtV0Kvyhh0ZAk+4QF9VEawc91hvGGKsEa3jX6hiH4Hu6WmJ
qstxiC77goHfRuxQx4Z0MSO/0cgO2sWErTPgXQw2qU832RJVx69RJbZgNIMSious
VmIJvVPq796jI6tJk5Vb/X7zpTIC6a4TISp6KvGiFcoj/0luamRV7os3I5vqeipK
aNDnMkafRd0Kul6LXIP3xchA4obfxPD0eBBCrmZ2SNxA1m+Lg4obllNFdQ8TQdAu
atvtJiLd4Cgky+MQ4pjLtsKPEb7VhXgAIwg+8lmDaXxVIdOFKPzXfC/QTAJn4le5
iduztR8pS3YFsEpSciDjaek6l+Arzh+eUtnxoGKwGQgN2YauKFtF8IfXQc2NAxG+
4GiExAdRdDts2/7s+G+WcxRuw6oS0RJmatnFGfO/KDo+nYKSViWvEWVkddZhWwSt
/W5eHKJXtNYz3Xo0QN0sveqDFaePnglFQ85iQMgCcBHNLJWX/zeKmYJqC54aBUB0
43mx6TmRtcUTJkQSLPGv/rfAApWeVgilR+rtpJVHqCjMFFCjUqJ3FJbVHXA+zd7u
pm4YTF8aiy0urkBCRyKSm+Su1RbgIrEkTsFCT4hvQQmoHyIG7eDAS71u47Q3Fyqc
3BLUGZstT1p3mFae/ypqFaA2jgS5MZiG6Bx5OiyV3DkH4jbMqL4Q7QTHApKa2/fU
B5ywEhnPmaoVhzP46dOFZ2QDIpqvfWwESocSmfLHHJn0oAx3k4unFqIcbWvvq/Xw
kZLbhTBzoAeiTN5KXc5aSlbWVl5Fm5h7/RNibunlHpMBJipLUcrZYdiNy89b3ZVQ
u5hMDfZ2Ze9qSo0+bS54lLCNlqsbkO5Z8ARqL3kDnCgrCPl8LK4A4mnaMz0IsMZP
Ca59YseI5sYvsm7k1HtgzsFdIN7+cy0Wwu655wEm1pyIUc6W7kTE17ekMjWjV0/7
WLf9P/hBzv5N2/z5OCt9FAIXjScLX8eX2VGZzT0TuJRQpnrda70byF0nIo1gfFo3
bbEZ6iBn17jY6f/x4vbXtK86pkfpWRUbAOib96Rp2F6vWvaQf68Nv18WW9ZWlRHI
+Hg0E7k0wfFQxEcZ7Pnkgy+at8bxxbIOgNjOjzwQlOFLwWwB5zDPKAq0ut4qJ+yB
FsrLLcsL9n+URrXT/BGrKxbF0mXfgKPCXjoUsUBRutyyqk8IW/g9icthnhby11fO
Xvsiv1u/+zYtNTdFC33CM9Rg3cf18KE3LRESC4MBX8zmAxkCp5EVkB4EhbUfIDTj
zRa2+bDoO/vLWM+/CYheGfeoS12rkBhv7sW+6IyzwOMHj0L/tZSNsS5fv9KUfFEw
Mpa01BGVxkuOBerfVoOpWow4YEf6iVIDxDMoWysje7+/L7/KJSCgkU9Zwuyn5TPf
C+59abuLlQZ9R238glTwvE4D3GlR1I5ZfsQ8zxnBJa8bzWw6LsUKMh4DIapPj5mx
nA9I9/8hWjry9CW+leCfaUYEacTHSU0DqcMqDlRez5T4und9ITlVIDTwCu3GIBRL
jXN3xyf5jNrkvbvzddK36qE8BCy9g/5g5Djx3pbcsOoV0lpbthM74c9uifzWgRH7
R3m5j8R22od1oWY76aFrtiNR96dJSCo4VDh+TPG+FrRZrsD0H6p+IZDTlH0zUfgx
N1qTQeR369MtCxqTwtMfm8lmFpPvxDbagIg6q/u2D26mVHnFlvUA4+6liOlNSE8T
/Ixi0cnX2nm1W/u4EXaQV5+D81F3ZPFK+7Etp8UV1+5XNq95sZ/mn0sX+F9lKnOy
PUhNfdA5noXWLULIJe5mR5RSOT2fkGya2aIXrWTTFEMIjUCjz/OmGcNfEMymyO8a
9kVugKWPhqvgTKWsaBlIkjXze7Ez3ZyUbv0VwZrRixVXxv9wgd3xjelO6e+1+9tq
6G1qkovQ3/OClv/y21RQiXgFSeIrmrTHSxcviFeXOlY8n3U7+yMxuu/Cn+Kgg5rt
LlLTc3cQbCIdK9a49Rzh3QquU54rw1FksHMDXSqj9jahh5u8xXamLVXMGaVythh6
CBthrW4e/0NI7WV2tBBjUyA/byb58HGnPJH+HXdteXKtXftsq7uOMArtuWemYg+B
GT+ITVJ3D3gsRC1mVH6NoMfWTbjBbsB/NjmsCWHfl4GdXtD2egTw+8nllDCcwhZn
iPEsXOU9KCfsbPP6Z1F0P08YhTTfqRESK3dGc7GiNgZhDZ0/pdJEqN6oT3Wkjafr
2YH6Ry5bjptcyD7xHSMRD30sPrjaSyxd9nsG2xaVbIkqX5S/3BCN/FA1Fe4IqQQa
3od1xbpO3BT8vEW252AYlpiIMLqn5OOyZg5fMwK4pzGLTO5BrS5AUoPNa5VaRaHw
M4BHHNczOS8hJ7C4S2MplnStfnMZToosJPVdYwZkiofEbV92QZ+iDUm2Oz0W2XJo
YcDdiIUCNz63qN3tFlzn52yhs++ex5l8iYYDkqCS2btdlwGyJ28Lqe2VIzF/BJV0
ZukIAUqtSIWt62skh4cdcHCyBbtaKXDgVN0pG363ibxdWMZ5eXN5/uVF/cEaiLIK
kgnx9VflSOipEG4X223vWYLVZFbGLiEgxLaB9kibKxP66HhSOnn8Pubh6CtXVYHx
oTDV52gvQpqO1+e9MfW9mwWW//PI4umiY1lhnUAnxnTCYxwyYz7+gPH1h0UBTcVh
K/0bHM2dh7/PE26JVT+fhfnd5BUH0VtR1TyXYemiPmwd63o3anJ5laZ4M72ZTymz
ysKkvOV9kP3BjyWAmKh9v3GjrMWTIbl6jYttZB6P6+CSSbiqhib0XXAhmy9iksdz
f/zTeviLD7h56aOiat8iTxa+Znu+hYTrtIvE0bfEyuzFqFkgWtsKUtr23VECk7+y
1gZQGDdL7zr2rXURNDmAeKPU5aXRoXE/J6nz2rBqyO28nzgvUEwftRTSq4pwRjLF
iWRYrTU1HBig+aNFBeyixDm0dXVo5zagvjpIQRss5Fp8Y4guem+tOV5Owtd9NeLa
BI/hAJY+4LV9ML+Dx9BPaOpm2U+hzQdiXMxDy7wUiD2kPj31n1JDj5KD/7vF4V/v
YDd4tbrSldW8hBJnCWQo80qOgBSOmKL7v739Qk6waeczkwyCTq0LzdZeavWTtTOv
0nu17sZvOv50viLDKf6dsGYazObLgn2ho3X7UjhGylRQlo2j5wYSOacn9gCNvQaj
02S8Q9bUBGCTYqjDla2pRyvXv7tyFBUr3r1BVtm47bQi1W3i2lqAD7SSbUuu3uuh
8ejhlQ71p04y6y7EKSBskmerscEJTCmwHF1GyR8JLV8gO4uyHzTJ5EqG+SS95QG6
xmhiomMxunJh7iMrItXnez+2qSREahDmaLZIdg6a1U9zfEc6SxGVzan4ogKTohlR
HPTmfLBVvPkeek2veiuSI3iNrq+RK6CA6fZXRjNWf+jVeeB6qIH0B/LMo0y7DEZF
mHioHFaEsU09s44x8gg3RvLurOmFM5Sn71SenyiLRLLxH8Y0FBRp5C8/dN3VKqMV
eycWXJ5Pfsr7Jt277P0wilSy/JkNRuQoVy3kTWg0ZDk/eqNQ1F1ARub5aX2nqHG8
1D71LmygZEvbNMqrxJMUnE/bqAViibV1odMzb0PrcE89Ku14BYi7n58yPeVG+qcZ
k+xsfkT0gIE0QRtf1xBhU20D1cyzbUACcVchbEbtyQByUminv19Suw2CcU3wgA4W
gxu4TJJeIHtxIWuo8UpXbK5wKkPNKnqXW8BJ8JNirEuCbwzN06snnSWN2b/Ml/fj
q9rdmSOhEvBfbkeC8i12kwXpJCRWeRb84iKG6Ed2kax/qSPCt7CfYf+wuTDXJA07
yllZM7Y2eflSkLiInxZ/vLSpuP4MYYntUZXy32Me0Z72MSliWRGztbAkAoTn9Yqo
LItni/y9iejK9LiGJGdtMtc1EM0qLqpcr8hvMASVD2A4UbM2swJcROKGm26Pq4fF
TmWZkO9ONoZwbIHvey6tS3Z8XkxOBAwYxD+PHuAyHqdcfTN7GOLfT4nIzbBag67Y
UQor+dQmQArH9Hu7MF9zmNxnnaO8ooN3SmAiddfFFLKiWdkSt6M1x3ONyiTXuHv2
3bMr4+d9F0zDp1jEv9oR6/c/H4UyxTFIZDWrQ3rE6lzVmav9/RpUObq0Pp+AFSSZ
ShOve+MPB4nhrjJsuQPT9lYz7DBH8gCUqWQbNxZobF+DqHwyhuXppX6gOoL/XnIW
WnC4v1KFKNXfCEZZHUfDxoYHcM14oqN/kt41LZ17VyUQsNxk8MW/agGBO1qNJq4T
c6HL+QP6ScUIvjMr4TYYq7cefk9n6RpPl/+YOhmXmfFcX7hfzsY1i+eD4vFKZ1LM
rQQPZwYauXvLK+1/yzjNi+t7xn0cqM6gFdiZ1al5go5ip3oKhc17y/camAUh/+TZ
1M/qQwiZUoRdYDNYBweEmaLaK+ASzYsNq/q6zsZZADuLX1UNhbQa05e5hmtgHtXr
nGruC4wLjRWv+oPzNeEx3JfGosG8rQsGD+YzsWmYTyST5A8VjjhuhBeE5+GQhPe7
5FlQ35KZswaKtnv83l68vwk6FLxKjylbwhBI1ZBUo6A3DTGcqAO/PAWYYCHcy85f
k4XG4R7Ra025bE48nF7bzFtatgP8vvnd0MqrJNX5ZS4bUIFsEQlz3R/B7pw9omC7
B044kdIu/fayomQJLHN7lyv/G6OTcNr1ExPi4qe3vIceDxN+NhsjEmkUahLwdgDO
TnlhYc8/wfqxz/VvPYSOAW6HtxRm4unix/+vkNmO2vZLmqKqHCBHcWQnt/hJ9sli
GlAP3Zjn5eKBQ051aBcgkhuVWZtXeEdXFj9aX+bIopMbD36pNVrQNUahbl1atrz1
fCFE355r7q7KBU4EQODaDDAQk1yC8tWrXlfWs9xKr5g04CN4QOY+m5G4a9PX3mFb
evVhg5hg96AB85lM+VDh1R1q8ca2RQgwB+kq97rRp0oHdAOf8opK8o69Im00XDpG
FbF2fBo6TWspm65GIT87vOZpF8AYfDYIGFbmdc4+7eOEJ8nBUusVDwlJl1n0H/fM
E9xCkozh+eRGMepq7qn/YtmGipxjrRC300EfKtxnW+rYfQzYKGNsRNZKDzQ64Sec
YvVEyycvlkKxl8ppzxVns4NE3pa5VK+QUlYW/92fqFCUG4Q40soSc4IifZSJmJLD
BNuDBXPygItnntZGScVVjO2edZd/ZhB14lWpSMHZr8HCzOMRdCM4FX5GPG1+Oqtl
z3QVqa/k9ua3OkVHujUw1ThN2TwjkQeFlVjDDJyCtBY7RF5O+eqc9E+3FovSOSpM
/7ZTzCZy1J2MAxbrxwkiC3tMcX4VNSnW0w6ZPbhPR3fb77VJ2E55sv0yEUbYlgEd
cLOj5dEPXZXQq9xXPLOs3E+YFhL62oGd1Ab9Kf301rOHpmX9tJZL9Hq/2Pqf50BM
fnU/Awa9PAEO1i0/1JPVNLJbfhAyqGFirEfdLaM+RppY5kBFI3cwo6/kWjWOQSk9
xWOsDy8a1pDko/dmEAGes6r0KVxZ/7hnz84rEY5JJXJHIYE9gRK6uPOxkPAsopyt
ljR8nO6WWAtzRPJw8f2or5wN5b/G7O49q4vx2rHY8fTy9KmGblhSFjb0UZI67aQt
kRp+QEM4CwqqMBOqg5SJ/2vTPAoK2jxErZFDLoZDwbKVTgwEMeEpFp3xdviiG+UV
ogVNO05q8bDVsMMSSH98aVbQZVDgVNSp5hUvg+iKi4bCtYSTQ2FuSAv/RjG5f9jN
PHq5uEdiInAO2aRYFo4ciuxH2mSuLaA2BjEJJqiJrRtuZfvI8uc12SdXAv+9SI/I
haeedWzvGdQ0LvbcjR3D/kJ+hq76K780yAcYOROtl+6zs1X3OJpX+yNazdhrs0ef
TNNond9wXBTlf2Rw07yK13s4v292qP9YIgsWLYxUoOpf78S9duv5Qh5dlCt/8Kxy
J6eXCWxUAKnB6CRE8wMA3+fuxD9jHnY6Xh749i3Dmn0ZobfMH3eoYxDPGvy0fm9d
mTV2jfeWqsQdyAU27NaD7ld8ct+6i4osepqtrIgRQUh9Lgky8RFrfcHq6QUiLz20
RjAeQNCdr+g/89fjnh1Q6rrV3VwqnkWQ1/R0/ufZbUuTFT0dh6RzL5iq9dMwVIR7
IzHRN1rIPTuPmaPrVDcOHqcopfvQMfh2c9R5LzBNNhS+OHLQgltYzUdyKTUSeKgV
sLS0jSzj4wqWg08rWjEHRvr4HIT+LqsgmI1DKDNJbulWIixsmxTMrgcZ1bEaMt0B
yPsPkvkzBU0jlYFUP7Wi7CJ2c47Ae3dTDJXhD7IKhkjAyymMTog/1/mEczIiNj5w
DZiLofLzN2wNoK6HkB/BlacIP/agEwwucCGOh3wvXFnLd9ph/Eyxp4C/P1wskAt/
2WU8660I+LLeUswMOl1zApHyJ4xEMOZydY5A6dR/eBJqXc1/j+4G2cvCZwCao3yR
7/AWf2RaYcWsQLwRsyvO/ZCcqmHg+YYHwJe9XqWbjAX0mCtWEbwCSV0RqhAdKlx4
HXZPB73KL8gmNswjmYT9pAJnSAcVnfBO6tlM2OLKIGMS3XbVz9NQ+yaraJckEcD5
rXIVGUAj2arsyBWtO1F8PbBtvTQUVVeb1aUcq5qZutj0lEJsHuRFFkNRpLO8vu8v
bdNj/wGz2UiMdK8njv20rPCiFv7taNw0pVyI4BDP2pT/Qmc6AuS84X6oJtDOtSRE
BCMVno9EbCJspiAyGmC4AtNkPvTdZu25ISdX967h3PqXaExaEcr1FLYMREIuuJpp
voFDtLTyL9fxlDZTYECTVA4tN7FLPluQtLckpaqBz5jZVY3Cl95Wc1FUrC2qeUzR
wnByeL+rhJKiL45vlllRKTF4LWioPcpRWGN68R0wm0ZfR7KZWWtljERIN6tiTQec
ge/6yU6r3tvVk22JlgvAi4dRvxqeqRFp1Q6yhgbPXb8sGRniBrN0ZlkZ32QZf1S+
OyOEQZF6dJvh7MapnKQxCo3TxdhC4bPaafoc3XdGe3eZVeWduab4BeDxHIvzOO1/
6hfJfJaXVTgWgEARDvb2OCwteNwYF5+SQJFA0E3/9X9NqD/BApznqthjDHJZnyq3
MQ3qE04oOJUV7s/nV+foZUh3eTmiXqhY7Uv50YlJCxsFtOs6L11Kd2/FAAnJ2Cpq
Ga7PUxz4/fySfFOWYKVO+POTq6hE4XEidZRoa4cevP4JCBf6W5+7h3auF1dCI5qq
aSuFzMDKVfraEg6NFazPCtg1r94OMxXCNA0Euq/XCln25BxRp7FRb94hr09y4Bn3
ukMSi8Ofv649d6HOvrGmn7cDjVw/sKFuVy0mY1o5NLmdLRqGnoK4WkCH0X8mAO1R
FEM6rO1XGbH7FYvLrTYbonvfIeKMA7I24UsYeSQ2hyphvsbwc5/zlozfsTJUfZ3j
Is22pDvgh5kqSQ9w6IXZcjJOcBroYepmztkqi9S0x6DNMLDIhc1cbSenk+FGZcyV
m1VBXSDxbQX6WrXDVvrnY/Thl6fXS8UMZpwGlqbSckwTxrfJlc7sV4isRI+9M328
BFCVju4AjN/Nhh10aijmmDnskwcuh9wj7MuBUgDEMXoMmjMAgopdFvLewb+ij2aG
cuJvtl/bB9UhY22KrmLwQJSZTJyr2dBTaDqOJc+hLJZhxYbgYmSUDTLHO59Bi7xj
i5lFx/6owCIhpOQD4O4dpxDg+ThPSnlDYynp+aJTHegHWbUohldxFoZYa4AM4IVa
ipp8y4N1lC4GhyvlSISbs66PgS05uDIqzLiwlsy6H69Gqq63/v+UjFjFYMHqo2Ng
r9IQInEgh6EKRPQq8fjoWYV3EPUQy+6BNZ/wTVN3ic+h0qdODNCBFJI1gksHnpS6
zQzLV54WB0c5hWfwX+CSmoH5+mvM9p2Hw0Y6Wbp6vvBN8gfu2oUTJXB9IW3s8TaO
qQ9GWaedA86mdmfgy56YIE0YpvRc2GgMk8x+KGj4HBgffL7LhkWq9lCAV+ueteWZ
Jpeh2B8qufVfOdnDlK0ODfBswKaCz2bYBqPUuBwYtAqNKpREZTLaJJXpGNS7mhlA
0G+cgXB54lrLdrsWNE46UDogr/l4rWy3lmE9S57Gqoxr41pEUhnKBk/JYij1ftND
Gdpbb9siwV1uJaukj38x4VibRwhAVtjnZ7Gs3zWj51xKc9aVaonbviFJC7iC4Ce9
pnNTLbLQSB5onXT0FDCJ/CPDYd0HvAlBsk7Wi52+M2Xk1ttiF7QBdPAHfjh7MMQf
9uL9lCyLviHzRwJ+HiecEYhWMqAPH5j4D8UwCcxoCBO87AfD52RPoepDcsVaLpct
hYBi5IAne0FDCVqesrsE3vseOsyRZ/06GKRTB4r0tIz9ad4OdTQ7EdAyo0bIB1Yp
+tGSnJ7MQEx4aiITNAEEqUgtWYfH2RJMQaRjrawh5BRcuTFb34QC9ZJb1ga0vnzN
JRPwCbMGh2MVZLEE8zPjq2EPXS5qucXJleSR6wvCny02TVWej/SUhQuLdZMQcVGw
GMGQWsSvKJqxb0IPTuGBI4GC/TEUomLMvj3sx5ZL9rNOKcK33TwcOEo6+acB5v4L
1FMh4HcgdAkuViB6D0gAj1pTfE+a/VS9S485fhHC2XNJt5lEaeC0Wo8UsAfzU+qg
35hzdE6KQAq5vEuDcXumyZGmmc8mCp48TwLppM3dBWbYDalcmA0/RqlK8FcxDUOM
6OLcy57ThZTxYp10TCR55QB+O9L1qW8SkmmAjOi8Io/S7mv65nvQedbIDCve5N77
m7hnaYMFOgbgyenNqG7R5XfncbchhDDJyLq95jivNkKMguo/0J/WPusChV9+Ojsx
Sv7HIsiKWFeu6nU1yFPmTuN3nMzeHuxNvOMdSBVcCrOxgYzpMGRpn5esEjOHs6H5
cjcDvacnMpvvuZNtqDVLeZpU4yO+/h2rn3zzRy015hjMQDW9skUoJqZ1tB4nf/WK
XrVk4C2vsPTENg/fwUjKg8CMe6WJcQuwtYk9MfOAHb3MBhLwgGrsqTlcBlMezy8G
18993Qo8bO0GO6hpZAoAfudf7K/LR8eFjR/1/3WxQBQc2oG9X1NLuAz1xOpRY1cC
YJJZBgeWHSTnyLFgCjIq08LONIuFTwBspz3f8SnvfXfbf/ip8hinQV/7Pytbm1K1
YyJGJGpCsAsbPDgJxUQ1CeyTCaPWIBZ85bB+C3MfPvU8Kp+/2B76EjF92n339zzk
vI9vWaWKHRgUpXEtra7myD8H3rMxF2mDKeaM7HCE6MsKdm3e683C0+8a0NOTuwX1
LgoNVqvu418doMh38B+IydOMSeWbgvLQgGFTBYMt07jYuMVE3haCFGDzk/u0vrXS
zHryePaM6QbKgLa47Yuj66xUkY/m8YZqSV6FDX5lZflwKzgeKHNfq4ch6PWv4iwh
8e5RwnJ9iMTGN3XXjU/YvGhqAhJxNKm0WMnIp3uwB+ZN35KcXajzdQEBrhlj2E2W
YtXUU8h3E5zWRJfEH/KTorArluM8IyTZ48PR45UlYXCi5/voXCEnzZEm4Ak/VbP6
wmf7OvAaHmjkufPb2WmxxKdcFEo2a2nb5f2XZhLJe0ShIkI9wzGGd9IlPAPKL6Jw
GQ13GH1bGrJbI0W5SXRhwTcH+vTy8FOF/B781zSni7U4p+mtgmO0Yka5KfbLXnrU
xr6W9p8qVJTktsrfvpzq58p2rMVL0XdgpYdTFqjSPUctK6ViHTmxUqH4Odz4NV9l
bsFOGcVlwkOHaej8Scp8Xvq47EU6iim12TCPFh4W0aVbxOKZQGc78Fft8c43O+y5
ylU0ZOtNcGW2jxWKrhVfyVbSDh9/jbVwiQhwe63N4Uf7tA4F+Ac+d8Kz7YjoWFRY
/XWCD7yPzupZZymYffdtrjsHY2MuH7iBpujoNaGZvtYxJwDRXeAgx5fo7zUemsEi
Txv78fmb/IfZDnCrowqCEQez2rGNcAtaEAojAXoSoeTuYVRRaB96bbqDT41cuv7K
l+ZCw0q+cMZ0uywljIoe3VaT5cCHVosAoYkBmQ9FjJHeld2rMPw4aOtkkEAkoK4I
g1jqpavthGkNVkjc0FwPE9DD5UbYwhdhshjOx8Hb3w8uTlANjlI1IGwoMazyTJl2
hyAj0TZPXswmjfH7GWEr+fSaOFY0A61XVS1l+d5rE9+lIv+z8xU23jG2CJlSFMKe
NZzw52cfJbOaFDXeS8R8QXgRBfKXvDIM15dZq4/26KJHnl5jSuoBCMK/qKmVM9nl
QTAz9VxcPfKHwkjbye5PvSahDM94DTuqys+WrnodhU8/ub7kuVZEQgW2je6A5PED
vhKp6c+/sgLY754YJs7CCK99bvpUyef5EPPyOuyRBEmlLvvIgaX22YrSe3yvmocz
VlZ4lWcOVFR5SJEkHc943K09yUqpZM25CdaTwwkbHlQGmCQNSXM0akFi83S53rhJ
4H318PWl863KGwWkH6YTWFek0qR5qSy6n1WT+pWof+6UsPf+3zIm2/pK2XUtMtt7
TvbLXlMHy+RQhYlg9LwQ4a3v17C8f6sVig04rVvTcg84DOtB82W0pqQZ/lwX4FGw
XkXC6E9HNOV/mYmz8X39fyGuzrR9JUw558120ZZkmTISMBrHxmBqxpgvto+Y51Ja
1vqwxLMvCtNV2uqcXjKX/35K3av6bdsOZ55sU1Z2EJIp76I7Ukz0quodD89FK/10
ahgL0cNp2OkadzxKtKBeYwfRGgENxOug4vPUFuVo4CwQP8zWoLVC+tV3uO5Rdf+8
0DRijcOLDPmZZykkdrrOMFSkd+BSI+IcTpHe+SdY8QkGikMUzEu4siecRxOVM/ar
AbK3KkLyS7iuDazetYeH2DApVXYeYNl7PfklrBW9vRIBgwSDnHGSNvj6n0veRS51
HYsWBnsRCPIfrvL09KlFZwc472aprKYL2IJaoYVpzunxcrCxts8jRaML7Pqqu6X2
3xFjJCzDCY7lXb9Lt71sHpLq3KEOar6WtkpTGisja3TLpYlllPPjOJGL+DXvEn4J
AA3hz9s3bWPWqyr8RI/qqjFW7RYcAst2s0oPhDWQqWmiCrScBtwT0fEQ4LG21cA8
DiXhpk32fl5kzVmUAEsijB+MEmK8TYY85AbfxGgIVja3c8tZGgAktByiLvaspPL7
TG/WS+5uE/7OIWM/e6RO2NMsMe0bc6iSHqB3Adz3l/zwZOvl8xZZr/7bw7FwiqFg
Y5jgD3eGaQu9kNgukQCxkDBAbaqHvItuKwPfFh5brHxoZE2lZ9W3oeM7h2q0Z0AX
kzW8f8aIqJkB3mSd9vPE2Bx+lC3bpnpP8o+VUXtmMZHKO0SoAScAystvoNvy4h0+
WB6wFT1F2km6eVuH7O8+F2zo2NM9807mfLhaPgRrK5wCQb5wMm/LcFYgTUeytfR4
1Ac9Gga0EZvMLVugtrbzcXoC81GJci5k3Wyj33EPJywUZhRDna/lSGbDQjtcv8Cp
gwIiYbhAMfCB3O/inSAr1pRupYqo3gAlmxEJEiMi383KXi3jhwvSq9spYnqjdcWq
BtEkXFyz37ZGiIa7+v8VsK8GHsLOfgs3v1fAZwb9jfE1DWUksqBjmQ1fwRAaO5Qr
TvxNU59p4PIe5SxHYRiqzqsrHJ7LHBDSIursym32AM2ZEmsmCEb+yYdj6CPHT6nw
RM+6fLV1NAMeIG0T2XpAqN2rMzZHy9bBXSx+8QBW7ikr2r7flbeLL5reEmHrOpFG
S5E4hBGp4MjsHDy02E2Oy5/rbwLe7iz89CYl8lKLqiL4NcK7OXrqk2SuA5I54uSs
z7L44spAJFLfXS0HSROuBq1Rqm/kbVzcjRB20d/FzgDoJRb5XHK/ujaeu21JeAV5
CBA9TnqS/fCmi8sMKEehfpkJDhjmK79Ns0Y3tln7nbzv4Q/w4OsnT5TjBLkX1h29
RzLmW/YBcaNWKGzOmeGPHvuBNDQAMF0KmypRKKg3VennDyWJSqv5D+VCgWGbGrPV
qRBsG6aaDG5C8l/prrqlrdqbigMjzDQK5iM4wlFLtvQthkrfY5f3N2aufVANppor
wJbRthDykkeZRmMeOT8fTpwhsTYG8xoawS1gJqwtEGxS60DBm5AS2xs2ZB+Me4fo
f7BwLKZw2el4kciTbzbGOPTlZYCAMHdIP9A9qh6gGOyTPYt39SpiJuzjmCoOf6Q2
10p8disHCArnLs9nF7CErTx6o6gO2TfqWBxnJLZ9CQkubpc27rtWTMZEmqC07AaG
mGGaCH1m+kQKWBd269172aGRVlVe9FafzvxQIcvWE+8/+BSEnSIuT72YhMoY7YZ5
D6B+yTSSo7/wkS5ytAZ/+O+++Yw1SQwIMao2J6wFCQPSuH83m4GCyWZVzV+7HFFU
Zd6z4gn/0XB/qbcfQQtSaVbwHxfJ46iowD+rJFbBd+6hyjzFBIDgPmw4nFnSwKro
gFfWqBeOBeTxEgmExp0sSbd6PpqUnF+2eF6J1Zrg3duP/3s18S6IjP/3iG2SoJWZ
VyImW+ywuB0cL9LPF7o18t4ZweOCHN4HaWe316DQDGpt4lJGE52zA+z50v+s3dUS
MaVP6rMVUqOcKimKknFD60rqklu5jjlRDMpdszVTerAein2FbFM+d31rDt7D0XAt
mkVXNitYBf2slpb7cJ29E61bTowT6N6CLntrs+drnmZr5WXoTO8qCQ2sWlathgxI
q91D0j0ETIHAzcxjtD7IATWnE26gk+ud6RpiBhK7QNVJms+P4eR2R49BpMZLNA9S
6y+Xpe3SnkJDawX7jfcqkC1X4sl/CY5bHJbxNB5RdPMgOhtUzujmdTu0LtIpVP8n
WbKe0VHhXwEkvmcrC9kqQgGo8310YEjY2TOczTb/3p3hQTrm0ePZADPlj944RzWz
Rh9sQoyLF7nAi0aiugPwB0H31J2mxPX1msx7ZJKUfW6cvUBSKVj/Ce+clLWRofno
9yA13sXsuhPf0HjE8vRkT3yp4PZEuRZMvNOZ/qG3yanYVUeQ6jH+UoKj3ssJGmF1
AMKazvywGo98QPANiPgFBCuVjxpVOj1va1jh/3Luf4iI6DD+HoKVVGz4yYKI9tOf
MaLe8PM7rNeaEFaO4CL8SZR4D9x5q6R3UfYOILcLDXJ06auWgsmA5jaJQ8kv9XYS
wcgKZNyYL8bjbPMixc1FlZB7X2IcL5eXGpOhoAIj3YkS7Ux8zQXIOXlrL3tA56j6
V3uIofAOWfRqKVH1eMDvcHO7VxENdrV+H7zCenejzUan1j4xoinp/VOHDfbEhi1C
mPs0MtwSUuS5eLTd5dzTPxKZz+D4H4vuu4ySLY/1wq4KGN88Yor87+zODNGla2s1
Deh7uvn0MSh3pIgNWrc6wvQy1sDX0IsQwZZllCK/GtKa1TOZfYHubl9JP3JUuJz1
3SNodwKlD2D1Y+jq4zCJUtEBcFVf9bC+z+DqM0ZOABWpUAU0Xwuf5mr4jyeIdz3m
8cay9l7fZXtPhFM/EsUeZRGaDy/UHSyRZ5RH38Ds9LwU+6pHgj+6SQTEk/LSWvwN
Di2turPhOiP8bwVF8kktZLtmu9z7ctx6DextK0OQPmEO7Lt28tTgzKiRDjrmhfdY
R2jA376ADLzX1WEpLWCk2j2GrxmvOBR2cWTENgIGkr9kRX8r22i7eKFlb17dRzSA
6i292iLa7iqKjG+YyfYD2ay7ogLsuoUXOTUhXYe88p/Jll03PJ3r7i6YDJIy3l4L
zA+ObbGoReTxgdnK1AF0T1HWrkWXwQzSgs66917526rVBPKK8HwssTEDhMaP6zak
rZQ6+twt1l8XAZ9aOhwSJBsCN3a5EvEs50N9kHNlUtDGIULwTQMgyksdPxIxIKB5
2uej7qYxmy/M10P91uisVxUp1VAifnebbJFJ+bXudIksi3nFYLa4pKOUHW5FKLij
HcqObL2NTE5YWVHVXKpUvSCZLGayammtsMJDSjYxMehcAnv3PK/zSdI5w9YNdlmp
Kfr/QfOlOJqadz8iDp2jmRLPDk+/jluW/cIEWR+Z/ZxvMLnfg7UXYEbPcS7W+kRb
M3SVTDqwRCnMJ9RXbexgLCMPian6EMzoRrFsz14VAM/Re7wtekpnSpzjufVj42v4
sL4/oK2mhg4+BB2OToToRcPUnqyohK2d459vBv/41Zv65kvdlBwVtWlb2mAreb18
SEXueN+G9CoW7jYpUuG7ndcHmQOszhc6yWap0LQTJXur1Br1PdY5Z5JHJ02KIsxg
HJGDrTjUTO4+muPQEB0RJjrKg+0AlIIZOSX5PerVE93ByNXhgLnFh7BuE9mICy2N
no06usczQU9joY+c5Tu53PpfVNKImmdFeQZGUtFFdHBe03DWaZUNPuk2yZ8nVvT8
LEBWi5oqtQ8yHYuc5lOacv7O7m+8A5fjOxNEHFZlr/u7zbKUYyDLoCdQLmzhNJRJ
+k19TdJrUaV1yUIGwEQ/juMMaa6AD6Y4C+EIWvdb22bL5wbiN5/6SIffdDuoBAsV
FbMpovRpjmTp6akbt57COS4uxRoCsKe/E1fI4h14sQq5/haTaMef2UOPqkhHEXt7
JLClyLFotiJoctN8AMFa3yWy3PvSduPAZ3d9eEu46TiDwjahg/ybZRoWfSJlu1mE
1qZgzTugRtMCG2bq+/DvotMH68HaCcsQUMIA1jKy8Jsev0ZKsSyVI+h9YSLu1IhK
kcM+esY7ZEFOcztaX6WVmNfADHgzk4aTt5O5XTUQvLrSbJqy7EiJJYkLr5EAgscJ
f9J7tpkmT5GJ7XlxcTsgyxe/SDQw/632dkbaiEUwK2+abdMCCKmLqFyz95a4dXWO
MsECnxYdwkMEPM5o73HATMKDIWMBCQbcklOL2Vyfirzd87rntjUhdoyqtL0vxqoU
epzEFvb7R4MNIHcRvxviwXkw5jrEeVQStyry1X8ffD+OUtqmSTo5wZo0AYZs55la
3fT0F6424GRfeeJlioXwLN79/LlvKZEePw5UObrcZPLveG02lNoSUS7eK6DMuxur
bAZMQiXR1AcLQ94/yw4PZLwyXfBxjFJgCJrE7VzMZGjdktAAZSRkEeazYcrVYkLZ
f7KZKpeflm21Pg8/Ke3u0plKwJKS2swAby8QEZQOtzbs+lKz8nto0/Y8ewgb4teD
4gt0rwMHTgFXjqvlVF7DAvN8LSXovS6+ifMsoikBzTfSrPVL3eFSLwrWZe+m91mI
W+ZySE53QrfXWvXQ7sXkp5TXgJPD2kV/PcjXpCL5eybRLu7WCI3OIsAJvUV4gClQ
6rEPy5/vYCyipnwmsdgMgK7hp/2uB45GcCFC/ykm5TkDW9QEpMM6x6PhTLuM1y8Y
phxbos/cXSuQDlUm1LoBBpqe2Vd0QWcJl+ZZ6YqUV2LICklfEs7XAxEc1GG99E9+
IvEyk6Ha0Kgiu9mkjScUtEEGBRWzUPQPGeOTSNna0YOVvrJauxxvXiH0SIvPign5
1ziA4XyshQB2w1wJ3P3yuE4WSGS7qtIRP7NgunO0IP9zxTYx1yAi45ITF9V+E6xR
6ByP4cCO2SsvOPqUt9unPRAvft/R3aO6Lpg4rd4oCBXS91xZgCrtMvo4Q4vNzTA2
9vqHBgt4sRVRaTEseI6MLVTBVXPle3DNZESMwMXSnbD0baAKmcZsP15AUR4CcDNq
7m6tsJxr73gXmdMleDxn0XoBYNuL9qMUeTMnohmUokHEOpHk4GqIuGjkBJB4vGuL
CjpBt7nVRi7GdrgN6Lh0v/z3ZgF4tkb4ekuJh4LNhZGdcqjAt2bAM41JWbRiQV8A
XAu7UsnsRYqt3HC3N6moMljU/65DOX2D9Y+IrGpwf7hPLmMhB+xTiNcQcQhZAQ2M
W+t+J+XcSSmPZ71MPjrro80LeXRTA64oh84YwkpacbHUcPkWoTcPWlzWIl9v5lNN
SYFtd0h+CWihDv+Lre9n/piBTdSWSTmzCgKhj1Zj3tpU8lHClu4G/QxKexXrAt71
olDAdc72roA1ldtPyPKGW1b2Fy6ydxlHVMdv+nI9HsjAhTM9oq+j3/NgJ8i75jFQ
aQk2a9PLgNYrGfxRJU3RXfZ67a2dmz3VNBp4d2hn8hb+imrTY+lzC0WGsUSw5qfn
0eiVuGV5YpjLaB85M/+jy1acWC/90yA8Iz115BP2/6/FFQGxQMHdF0Lzio+3x89W
ew0Jsv5moqPNz65ohIuZC4XZOCOB0fvj04GMb+gJ77FeFaAXiozUQ+gohpjqgFMb
irgnr2SnHFb7a9UHcG36kTXLfwHDbWzOoO9X2sYURK0dJiQQo/yAFpGzkz6i6+JY
YhUXTLIz0xkpyxBxqx3+Lsaz61oHJaMZdAt2AzWfFAZMS/QXJPX+S/TVOHl8xh8M
XlWtHHSRzrJ9u9zW3t66EsPAOykNrKLSnf+KGAdVhVjw7oufiyXwGCnWlpgMzKaN
aWQPpgLWT3nmp2LvY6riXbd/ulX8E/VusUIYzsVhAFUgA0UdclEWwV4hq9MY6SuF
+g98MzxO6rBNRYZW9R65uW6T0ySUSmQ9vdMMV3cS+S83dh1UR/9HH56aZGcAl4ON
zy46oc3n1yfBfrMfS5MpkKnM+tl081oIrfznS7OAR1PwnoXt/f9P3XEcjGUe3QqR
XE05uuuQLwoqxrJVU95Cq4tw4y6+w+0TCKOIlBvAq45ZEvRHd6xUGLuGMrmFwm8e
OkQa/9E7ngNuf5ED//inEo0u5880jxeOTcj1GbsQ8wNslBIsHfhZDhcZxWnMo5Qz
K8N+SUEow+hZWS6oNPreTvfXF+9yi7nPJOvfdcdIsuR5J/7NhzvDkTKdyn8m2z59
pkvNWhtfJnoJpARVJcZXu/ndcKqY0G2l6ZjgGYqkXg21P4zYrsfovP/EpHLMXFS4
wzqsUtPWMvh7TRDl3mvT464hM18ivnc3Obkn43SZYLYmhxN37yBDno/LEhq+3VPv
DRkePYbqkp6jWxOW23fYcsBcWDSgv0ixpLMXIts/M0Mc9XA0ctujqZa7uwSFDpyh
Alla7QKFxMQMF3FKYOeJehKck+mDhdPgqakTvPlYZhlBMK4eR9sD8THS06tBKiLM
jLZKSlRmvCDht+W0jGXaOZBEU3xZA7XTYdY75KUSESuTVWVEQZzQAO/gBtC8Gsc/
sXA/rQ0NFx1cwohagEb4UsZf2oP0oCVVA/EQS2r4IeeSAxAVFpW4endnGyPYSRHd
mzRbCpGmgVWq0unvVdoVMZECMgb8b8y0RvAPsYXMw2s8pSu0x/t36Dh25GCG7sOb
2Tdq+opiQq3LjuoedcEQ0aBGGgbfsUFOt3eadZdoJYyO81WOozsgQNA2omGcYI9G
02v4dAmKWIjKqH67dJCm9EqSeOlubfrE4OexhR4syLNnDEbaPfE+0480SPf0dZqE
fmk2tmt7IV25Jooumsor4ELPCRk9M8IfaAK0ht3f/fI6XD1bpJyCXzYlXY9sWL6c
r/USMeFEXmwbYyQ7t8AGtuiOAE2CLHWx2/kDOzgJUTkFUBFhnQHrJkta7A0s0Y8x
4Jx/uU2e7mMROwjdv7eH4bCEnAhpddhKwoJfyqc0DD6N0qAovpIJu7TPu80MHcTD
8PMJETBQ/LiGF8WGqrAflfV3Cdfu5BDHIMtDVEyxd8MfSKvelVkBHx5fWB/717YU
uRcrbtSvnjq/UUCVkFtJQ1ai1rF0rJ0gyqEngRQIcOWaACAO+3TaYimz4Fw9V3+4
6GIWDaBDwEls+JHm7OPIvV5ZmB61X9+aduI/NYSdV/ABHRhC7/vEvAg3x0bFF0lO
VlEjdhH3N+wuqBJWOprIyhOIbvmWLasMbQNCImJw1elrdb/TJWm6qFPhcYeS3R7J
9KCfs7htzyCWt4G+57m2fJ0bOHO3D6+L6wBo8gwEoZ9jB3/77iqRxhUoeUWXV58f
zaKF3d+deh2xMC0B3d005u2lI7bBolF1g3yEC88RivdFGijL2zmFwEXAJTJkfspk
U2/zjOu/E934nI9lSBcvEcTmFDPVgajb50HmhHkgVZ0Fovn9RNp0spqNz9AlI3iD
3fzPc5DcxyETGxTwxoNvPTAWEUAFCpakMPDB0iDtDw2hCeUKfW9pVYaAkIVwAO5a
GxE93KiexKuuUe3gk5gzmth52VXVADel3Iutp4rQ3AYe6ys1P8ovTjkkaJbzfjVF
f2Y5GxNiB5lcKuk9LuAmhYjdc2Bzo+U2+FmfnxBNgHvF/XGUhixwW41D9lykmwKc
ZP/D6n3r7mlmG/E9nbKrxtobBhIMXgr0BriShztpBSY/KSHw/coFrLg8c2pnDPta
Mp7z7rh4oiZdA2zPsJFeVjGpPJZpMA+HJzujksiQwfbEvzIHxWmpGBYcrSlQl6RK
Q0ZXThX9RERYlA9rYbTaM181lsI/c744fdlDtBBtGsYQMudB+CRi9H/TD4vraTi6
tqGNmAIj/wm5S6ruxTFeJTb95PLdbW7/6m8qt5SvEZMbjsQRsKxMOWJHWXzfU3nY
arBIE08KqegFdmOja0W89Kndkl9iPrsgr6a5KiNuyTpb50Ao8dPPSVLncbIP/LQ8
CP8/DzhQcAAA+DOoDoPkirsVNa+SzOjSLiz9b9/3ej70Q64iKegaB/eR7mNRQNZM
d2IP99E279diY0mKyaF3GxHq0AqExG/VZ6YEk4dCcCTnOeaK9xhrjmxQWnsnpjio
FY0v3ynb+XaCi0/tAavd7o3PELlAUVJdBNcd9LSicECzndPCrSlSwDJ41FmkEHL8
xmgHpNewn14PJxjufy/1dkV+gEAxaJELxFZI+naDZscVEo65Burkbfz+gYI8tR40
jtyKfokJqizGwFccHV8W3JGZ+V0hIHoA7wP4SziQhJQFOYzNIg/kuf9Z0v71RLFG
luX8INcsKXPdlXiUoUG3H7lZ6giRrPm8rG5/A5e7QYDf9uay7t/48y+47ZvqldZB
FtyrSg7BWKVhYI2RW1rXWju1SOBzNuPm4icn0EMUFWoUyeIaaxSHYHF4uNJm6jJO
eCRy0ope9sJWYTqoUGBDE+SscaKDSIhFp4FG9lYzC0Eo6tYNUJCp59rfDqBHfUxs
7nk0RhaTMIvzyv/yNvf9+i4uX3Ccsg2KlKx81MI8DT9XhROpeu57qg4kkD2dPvKO
l5yUBlhJxniA/+7Uv85u0Lm2hda1mtD89TpXMUVIrN/5+0tXx2uE+gZWoyU3Yue7
1SZTL1Ftxu3LqD6uEkBuS2/uF/Ndu+kZqNGjicTIelTwKGVwyt7jgrJAFVfqgSXF
tOOWQrbzdDQoZ7PUF9HLKrZaMV65d/QGiTGVSyQO5Xaiwl7ofGkJdo9XFV0GfDjF
AljMpiLlF1g+NlH99YMK1EGksgYv6mM4CqzOlG/4YfwT8A+0Qa3t6tr7tpJYQDOt
AUk9SN1jmoxdTHzcyFWX13ebtfonNQwT1W/MsZd6Gb+ntonZ2CP/nyjxeLbSVAGj
VlcUA6eeB19ND6uf6ab0x4SoB7RRqwBtsX+UJYL3q7rZerGSdHaj04zF65wvqKub
APbfSB4Xbl8rGyM6V8QdWthldOyay2/L1M7JmJSdn2xPJOXvqg0kvz/x3tTlnoDN
TGG1tk5t1dOkDKciAcJKEKtva/YUNoe21LgYi/VDPKtbid6wVgiqNU1hZ3s2zNSf
+89UeKEoQkKlU2itJw15T+OGM1wbpgUM0j4op7XQFNED3aqSzY25kaUGpTz1Xfcx
cQGK6nKJv9jFxboNwHA1uPneRp2cGHMkeuMtselWnl2AnrSO75jnqtZsTzn+0L62
AQMEmd0f15bqri+64zEhCTdxADFS0O15bmvZhge9l3VJ5cJJUY/1GV0HtSslG8kD
uBZuQbsyRWZdlZCb0bqSShEQKU1Ft7hSduW753FDwgtqgvtGqttBfg2f/D5pI1Qu
sJuyVYNDktsVItDuxDdFjXA2nSC5/TCosEvytNoEFK83UN5cuLcRvR4A+gfRi4Wg
dQZEwpZEIDvzZo7iH0+8nVWVA414PhT/DexE79zzHfoVwMzM2cCxt4trdD6It6R5
AI72MpYnl/soSOCixY7dqB8pt1++zWi11/jjeFNyvm+80GAm/DTz40ZI/N8SrVBs
xoHGaeJwF2CVe4TbT9twmQJ0h7YJaRc591Z+ZN2ADjDx+jR4BOyEQO96Cd10yXWx
SCkb0er7lk5j/sm4GFP+RElqJX26GqQRsus/J7MUKdLG4jr1Dc/is5NSJwEZPm7w
ZDe1ZB4NmNKfKa52fMtD7YZGthr3ZmoL6g14fEPg2Y5b52RqBB1QBERfC+Q35gER
xa4ORgSSWJ5UaFuIiIkjn6/ORZjiWVcQpvWMmn/ZSai3r9oMMDnQnbEO5yiSB1rp
X9uI4P1L3LohmG1tk9cWXTWFomvFGsBqbnAUR16+hij8WFWJf6TdAXD7Aqe8lHGj
ZJ1mXswPcjXabSXYqsI3wBqu63BsszcRH4lIJnlzHnDs1KqIvFKN+9uS5nYEZRXh
KIW/rTPCUhElCJUz1hywgL8wxi4QHzwFZjNlgu7wyAKSe4ufUhsOTlGWgbQmPIfg
3mFurN7GyI79x6zFDll+xUkx5AFvhHSU4nxnSvbAAa4hNeQLdm5IEOzwOMNd+8Ky
X1oYN9p2XMZUdlj1GZMueqDJqv5NICYNSEZH99wOYGghbokWXudnDflCWdtO2Vz/
BqEqlJzLprsi2b8wgyWfWV+XG2vhEVObSPl1EmgURDcB2/RGobFIRGaxgh4Ja0SM
xz5ks3EKSdNwSY9gO6kOflr99ZmoASPkkWCq9Jc5MPfoLHEMBtOHfUcHpLf2/M5o
KdY1o6a3v3jiB84TUA3xUGbR42pWRlKT9kdlgqkIezCY6FiN1gPOaOHnUYQTA/Gd
uSWdlU7nOLZ4al2tr9nvctQcGUc9YyNLmM1wwB87JnG8IECbWOmDpvdx0WkBSNgs
ukX0ZILj9WptirKK51M46VEozASNsZOUhZOwJ5hF4/k5te+YYUIwxAYyewtBp+XM
Cy4lAoSQB/X8lrwU/ForeW8eAxGFEhIHFCCEYAOVUtMEGbd/fpsPtPiId0XnyzTu
A7RWeKZABnCA3lm2OkVklkAZNiMHKYf5JhrdXe388z+VdCgJJc3RifRxrbOxIMlV
Epotsm7ZfxBqZUqwNhuxj4hd+7vrrY8UqxvNP5ict3eWj8qVP64FZ9VrSW1OufMr
9A3orL2T+vIA6+kmgKI30771UtbTIG60A33TX254vL4hnek1uzer37l1ruJznwWx
0oe3x29W7tGn59qgpNU8664WkTeGOP0Vk+7u4Sz3dL57u/QwKbaI/mSSFdnAdf/Q
VmLk+RKukt5WzILBiRxybi4d6RAPE3XGa+Jz1eVYnM9WJFep3uJJkDNo6B+srGa7
Mq9q4WvLK42wT7e9UY7zRX4m6ByM7FtEH3mTmRKKSlK//If5FnqC8JGIzvEpz8ki
NeD92LhJkjGx1ALE1eJnhNV2++zucAbyvUCx2YIl2HJar6NY4eODjZOCbxKTQSxO
9WQ4p0nHNTVbCGsyQaHNyo9V+64XEFpUm+OkQYDLTJWBUpeQoWmWCeoVwV2W+eYp
J6RoYvgGR51UKlLO03hPqiHm0QIs1GCF4wmx71QGf23Z5c+YqDZNDG5clZkZNh2G
r6nZuV2cHLCF9+Ew1kVsSijVAywrN+ayC4lOJEqMsetevNtKQlZYYdoItI9yX57k
2PNG7IHdJbieTrLCd12TfLYO60TQ3Y3GCC023q0zqJHO5Q89OruqKT4/93ADJgSH
lNFVlLzfItXIJiiBgo8p3YZJzHCbnB4fVeBrBEp5KE99NDqFgipcEtXdhMp9w5WB
LboLGQEYbJYI/ZwHPjaVALSag3JG279kW/cbcO7nGu98XGhPazjUeLL4x+7NtJqz
wXs5AC4v2hjLjhCcAFOHDuP7UBzItDDICKRk+sUycJjvtrPFzHhP4KVQJIvtSo6A
eMQwEoLT3YttvEFSpvK47FErbs8LIN5IXSIjKvnBKZFKO0qvr+fezNWyfsrBpc0r
++jmTHJR3NsbZmB8YXqZJGvLmfTO8oSzBwOY3eDHencBa2n9lNkd34/oNweFByU4
0xOSVwBXE2qX8fWLKtk9PIs79XkeDlhNFm1E/eBOD6IhpElV4ylSi3UOZQTSOtFt
PJ9l5dCKIp2WkHOcNNT1FuS8t+3JAv7gsjR2F4P4KzAfmE1lFRahu5HsAq1rzNff
GnY1Ts90b47ugu2EAE4PtxqKigYdPev1p7GprUgimj/AI/soWinZILP2m5dkUx/8
kfHhjMHprM3LzRR/TOmFOzG6mO9XTrflC/mK2ykoZEuQgDSIPzlUCN/w077K2Ezu
rNaTQ5mvSZIwyTyvbGe8Sza/crpfXzsc1SOt71EsfLHl9zOzGSXoWfziLGB0nf3l
Hg8ZfHFwzo4wTFtfwFIv+8urlvWJliwqw1ONzDHgYLMIN6PuBbeT5QtAy7Toz3l1
+qujPJklIh9rD2vTBJSLe6UYWGsjeBe5jfU+jrsXLggnOJHkOU3e8pmhpHSEn/sv
Ipj1THKrPTOqa2p5Fb1xXNKpwno6MLZ+ta3ertAaTQdZsqHEZpTTfYzzHfQ3o8ra
qdoUbSG/lj10yp5D/d94xu8v4P9hFhvbws8Bzt7n76kskof6eUxezLFl9DjMLXjJ
vooJSH+3989xo9Ix0qYcpQwkLMdRK75I7tF1uknYoIeMh3xeQaXUGPtFIMDesWu8
wMlS88LvY2XSYAX+4cAlIPVAnW8NwVBvYmOlysavdDOuM7RtMh6vfOeafG9LmrDt
y3NqrUj/J75x2Bmp+UY5DYJtcm3jXh0lBY0IaP+fi+Cp6KJOPix7hJR/jFYqYeKJ
Em8eV/b4zKO15B5lsQan269p35jk6qRVzPcTvr88jrT+duyq3Q3Tcge6qR72Xd0h
gOdYE6mTTe19G3V7vEhs9iHhZJrhwuztZssVH5q93ew+naV/IExTRtMnabEKMG+J
fbLi8pIRIJYDmQZJH81PDqHKiQK4EaAM1GVbKRHWMvpnZMJLR9cBc9DoZrTg/do2
tj5f0wCWVLri00wnuXuDnc2RK5U7K5ZyIJHwDwKRV94PCrBuncscpeFnv2EG8En2
q9huvMElnVgC3kGgt3j7hiIHuaVleYKbCZCo6Ops16sSY9f0Dx5XUs64DmtRKQfK
Z7f8nMTFnwDiuSUjHCcr4rbQ3/5w5vwgYqc9g/gvlOPt4bYdi34EcwAIhoMvUp1r
SSZoOYRRoIjJqRrz5OlhuzspxAaj8dXosIUF1gle8sqmiW7P/8vC7+e9RlJmmCh2
sHVuQjX8dz5CzSEHZuTed0aj7Q7izKTG/aDSeKesYJu2LWE+J/K1IPBSQ6nnVCw9
042mr6pQ30j8BFRRPe2OJXTqq59mLyAMjvrPn05wl93fgtIGVH7OKs2hXGyG7VKB
urtfSEQiecpkpKry+1rSTgwoe1m/onN+CzD1YbyPIaX9QNblL5G1Ajy6pZh5Kqs8
4L+hhv6jTy0sLkI9CVl0QHwB6Oeot6XQnJ4u40XohYu02cyIWDu0CTxOywbmm05z
9DyXFGd4IfToWqJ5hadSqYngN/br/gH/hC71bmxK4u8MfEMEb1SaZeaP4igtrBJN
pIHod+nccF661yqs21xHxSjaWGTFrODMN7Jktx9JZ0bv15WHo31VlDzNWb1Ozn8P
w1O76hQiQSvzyo8bPX1BtE7/e220DiqfCWPL85JJm027iCu5wvZ1YTZWRB0sPO2L
5jDzLY6j90OgzSKJWanvkcZ7bh0nbzrSES1xS3nYYO3jOoEd7YB1YhvsZoRq/SEd
hVKerVXuOqb7ucI8UUXzNUVFYj3yiDgxbCk5RNxHqpJT1lSNPA5V46d00WYH8SGW
sTg6trcDJ/kLUvTD+cRkMIlVPcE2Dv9yDvet9lypZGBz/qZLO7YiLMxF4eu16EIp
UiLMUU188YdXHuD3/dnzrMY/ECfY5dZdcXrKmgWKkBT/wAebX5aq5Y/t+n9kETTr
IPXxBE0UVp3voaoipw1oebHzH9kqCm/Hbgg8kR3zHZoFmEG0sU5Y0JdNFDuNiAOV
3bHBbgeMJotsRzGX86EUIzj3jGbMPCEk0WD7FWdmQM0JkDNgLzVSEPYCXNVMuWqd
AzmsPEWbuR11NK6iPl8rcQcUsZJqis5V9UX9woEuMNQLm9Vg/FVJpnZQaxs5ttN8
SMa5c1j2DZXpA8bfDmxFRd5zC0rKBba+DshnEX7uFq4h5XvRMO22dlzzcTNd/uTZ
lxfgnywh9hJQBEswWPi+X4yg+ywTBthNDhJx6SKp8FPzS0Pcb24qcbDgi3xn33ii
8DxElFVwW7GGnohYwD25EqypnD74g+eO/+v+D35Axl0at2TiXmNMV8flibphsewj
DJeop5dX7GTNaKzrtAquuUsGXQRbF4PCRMU5ZKmFtLYH5kg+p/yJ1t4sed7bvzJx
/13C02oVDpny1BorwfVWiM0zdOn/Y0ySDB4K/BfRtYqHX1yy9/9LYqunfy4A5tRB
ncWccmh56U8u0iQqbV/Y+fag4N3yahXt5N0m6IgtweBGEkgJ9bDMjUZpOZsflpa/
UcgKvv+C4MTIUj5Ius+JrXcu4dnBZjet0WKFR0Zv1VUpQAut49u9T4+pHVfw4hVg
1oYLu4p0OBm2IDqS3JNGYsSpTX3u//hxbTdKzbE0ul9vtj5aziZOaxLlAc9ukIjg
fLEupBkmzhsbumwnx1J1sUSOcVIbl2q+Vcf5+WCdPowcIBiUkB9741aC37GFw1Bw
JYoQwwXFQ6D8navakM3H9ySs/On020AiI1POtG4tUCgIDDlUu4ybJFLb/5seo2mA
RRw8dgb+/BPuXrQVKjn5ClHVBtij2pHu+QImccj1MV7wlcBUluFJDmnzhc9QvxWY
B8Zv63sD2gMdV0yOt4epbPjIfQqTzM/UOSd/ipC9WaNwFYW3kLjr2OjcQBYUQOxg
GaoSLQ7+MjGCia+V5dFGjI92dJ/+o1Icpjz+isyU5edpXuEBWSJBTypFHKcdAI9v
L7h1+sqhMZEgwfUiF9CSvNg4zSizq9fIeUYBTd8MwX4yYVgJAQUc/k7k+EOGwKEq
8joyd1c/I4GwipiUesLy4nARTn2t6AmRxpuZPUeb+JzG2GAah8GwUNI1Jz7/QicD
Hjm1KCETiu204TnJP8aRRD1qZojTKeILHte+h+0BKb7K8Dbjtf8haq3SWOIE3+w8
k1yUIfKIouAnKC0V+/eKbKOiuiuGOQZUz1HAnJksJkDm+Gd8Rwxcyjrx+5jLiZCi
G9WgEnQ2ApubFv8AgdQE/f25vrFB+DRxmJ2GvpFKgpjaKjcLYghfUpavWNp0Kmg7
X4+chMtWVsF2MW9k8Xo3IKXAaOdoP0nHEqJi5TzRguvgGLzuLtfzXLzuazLVyouV
C3HEEf4bVhNHngLtQl/DsOzcfk6nQKiHcDS4rq/cZOgzXrIcEr5eRNMpdLrQoYmN
56srgkKKBHZrmVkAgd/bGESk9czuP0kGWYjz37g7iMUqyiTqC/6XZqezJ0Gvt276
w1JsolgH3cN+4hlt71zwCel9Mf7YKjghHVqORJ90HFfzbEfnFvqAIQtEV/ZqVPgL
m0CRFflmuBmvb3aInG3nFDkhF5DOscsgbpecIXc/YEfXwjl8cLmQXPDK1HjR8if2
b9Dtjh1DI3dtDOWasJ+H/lrOBynf5/ORw2v8Dd6YITnKks/2gWNd8xbq3m2Ui29I
ol4MlBVwBPOVyRO7FaFR5NKISuZslwuTow7Eu4XB44iSntvBZYafGyzTQ6a0NnYl
9xJxGknofSjyNbcqWTCzhrT6KPcOh0w57CsKR7bVhMzfOCPjzywFwkqqrqI1EPQI
wtlrR8uP9eBJxjJRlfSpWTlClknOMedql3kIILjhaQL/QyhCeOJEWsQIVUAtUU03
nasBBzcSVgjiaoSoDc4ByJZVexZBiaz/+rotMVCKhAmPoAqcmAZoos0ZRUxIasAU
`protect END_PROTECTED
