`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2LwS5wD6M3Lan5nP2osbFST2ZYqaTXch6drconeTZV7FztlZgVrfcGa7xKXNKh68
zv+9ai2E18r+iijFt1+fv9fcygCnQpZPcpO/P7DJHu/xUCqbHs1DfJO5O6gSAPwS
3ktAkk1nuY0KJuxiA/fe372x30TWHBlRHkLrBKLjJYOffZA+Mtxtl3BsFmFB3RNT
nMSiZAkB51s7pT58SMf43HsPxi8QRm0BcIMgr+YMdp9pAiDydNT4puOqCBGkPumv
yk0XqWtwKVNjebkCLRlQFQ==
`protect END_PROTECTED
