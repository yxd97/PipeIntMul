`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/MVv0fP2R53u8g8/6Hq3KkRFosbwhNE/jQsxmcbeZelzQSkhuDa6szpQl6fbnS1v
tpkX4kqOYvT0wJAUk0tHU45J/0V8FPZoNST5Eahl7FqxZSaYu3mBMWIfQKC9vf19
i5H77/BSsPV9Z9BlRupp9XktBPPFzx4jgFrQWXu1jZjI+CKiurubkUA6d8b4wn3g
IjfzsWEMx+1vfMG9MpaSxlIQzVaEmWOSswHvi6t8Crl8ZDMsnMPBzWQPR8WfuAE0
SQFKjkr6aRiay2EG2hpe5ELTIAQxhoN3/+6nElH3Am2ZtrA8FfwM0SMiT6y3Eeay
jPfMduMUs1hASY2FpE/DdydfhdJK+JhwREAC6q9DhhdJ+zBAfut0pS7rzGxvFPds
tPemJuCidFHZ6gyMG79RwajTktjx7Y+w5eW28PilQhWw5DxgY0uct224kX+7p6w8
dZZRneguytzeTPPFlOXdvYdWhTG3BHh5ul0PgjpA8qZQhzowIfcdqjfh8in0+liA
rdRF0VX2YQ4zDvn1ls9lpLQAF0sIL3zWraRvql1yjnl9VTx0Gip0ks0Rg5mE6357
t2cuMmv9vLP1Sv3ZtHffh82ySqwvLPyvncu1Pd5zmQmyKh5kJqtbgvtHTHO3wkbs
V6ZxvF3mIzPy1wRocM7YDwsRnqh0SV4GvmjYckAiSRKnB3QDM+DQKxlE59PU75l/
2niG7vst/XtiHogeyhFMLOLKxmorNLfTONC3DG7fLOepvWydHFtdWNdYCIarCmoD
PlpZl2To1jGfNAK0x5IxUeLCtyxGKX8DdROSAT2ClfySu27eJMVqqlvUO3dnNqjb
tkeELOIKjNlH9rvjKLGGo/fSJDb3IAHgBC4yi2ygtXXyAo58rqiiPG6w6ER95Vtr
dYsxqJ+Gc62PvkcNjRYUDRcsik2Sl2KbFAiNuZZuJzVyPV1demmWi7GI/qcaqOKj
ILnqNjUBC7J3tSWO8lBHYBvK/QL5BHGShclbx0xEkmbpaJsBvmq51g3Cz8S1lns4
h44PzVt7p78VrBU09lHaVSLVSZzJilWCAjAVylMI/F0nfzSEIL6YrR7dlDMdlxxR
8kfcg66Jc6Rf+SHv9ReElqq3+cebP95cqE6m5EhkgA0M/FrD8am2ZtU4f5jGpMiU
x549QI7ajVQxclJ+DplapvsUdm70/0k3VP/fWD10Yrh+iFoq71UQQWlIj7o+Q9dd
e9UEtWS9vTW1iB+8NesWK0TnBGY+oVd4sA6oQpgtdhLYZCPgWJZLhuYXMXIuXWDA
g+kWH8D0q8zDTPNIvsy4/Nda67TRWIveTdsupDilC5G4i4kGvtmwEhqudR+wbtTA
4enbqj21LvKaGIPdlwUtq2eyy/KRIRFUzGUExdNkzKNoCHNxsRKlAtcwP0b9te7b
K6OCMUv/FqF3XT3uuH9fiNHStWJkFEQbqYJ7T7lopLqi9NbrkWIQ02TxZkfy4k5F
Z4xxR45UAKTJiA+sVDfjHiKT0iHAqZKV4rqiijrE6qzuBqNV4q/69N1Ct8axpLer
gcmDTsBjgi9NecM2EWsFwbTODfH3q3zp3yh5dxt4pt4lOZweD7k+I3o52GixhrR1
pwmv++JO+K/I9yQ/WBd3Na44J3m75+mCAAsBXwz7Fodcu4UlrFh7pnxj+NoC5zBL
ZIbaosHtmt5hcphSgap+y60dT+XXe2TQHq/0c6jj2v0t8EL7tjGyWzaKhBTGxyem
lpoudKOW9h1vwmsktDpKMAQLBnEDM1aJYaX4sW2leiaZER0N6QRhbmhz7tUqUoOP
DjhDHMmtCh9CcOaaGfB+/9/uIzbONU5hIdAhljSFOuBe6LLzN5/0UG26PXkQLh73
BG2hJxb23gNQCOIRY8/ZPJmYlYz5YUMusYfYI40uurJs3Bgw0wdLphGsn7kNkKDf
Dj72JaDnZOejyyiauomJ/orvbcQUrAQr0lD2oxEwBe0idiOHWIiiU2UYnmSX9x18
6/14/D6P9lPUl3sgyrvN5tpLSfhxxC3l4/Z62A5agtLOfDv4rdiysSd9jUuFC1JW
m26rBe3pUT3r+kp7DlS21beYIAKlAcwM3nBT3PmQFzyfe5nsd0n3qdmVR/JlIqYd
ebe1rIhGwaT+2KLn18DLVffcXKuRlqpnpYE0iGGUBD1EapxUiIb/ggLAfu8mrXjT
PmcOZhqhnskqWLlBo8P1ixsSRpOlyjpeoudLnzYdyyIhLtdsiieitPTvY1LppXY8
GIklsIXoWH6M+1QIPRZ9DyCgRvhzKLEtRsIQAsNH58e6nYZfqV8K76TtrASoJo3H
cauiB+3Waq1jqtwMazqjNwxG/TzoT3TkR+2xK+GnMeNEsinDVXU2DtozjilEI6Mx
HEy5o4N1CM66Ev/VgzPBaoSmGr6IjVPOFOyL7SJshu6RSASqznJwr1ZxplxRevA6
5zSiDbFk0mrWKhVAsGDyzN/qgnHv+TmPj4VJC96cTiF544smD6UTS9lwMgsNArKq
hWAiYZk+iaXqirdzVH1ZPxUPFTJ+vrUXV3ydsszr78vsb2AjZU+zHwmUfSLMb/Z8
r81QCxtC3NEwO5OGj7acHZ24ImJzKkoA6W+HzEgiY/UjSwDaTPZeo9upO9wNGWQr
tV3SP7WFcO0thxCSjnCX23pRukpPt/09buhvKwP7fJ9LdeHzaxmNxrRw7MeogJeM
814Q0On7UQBUHcOkWolQLQy2OXPxwIyom2q2NC3J53VEhXKnAt0HK9uUtIGCdVhy
K/GQ4+6KelhfGZkK+TnR50janYA0RaE37XnBsHMgQ4UuwKK7o081yMcX6Ar6+mVL
XLGt/ZagSaJgnor3sULbvA9JcEoCdVo1Pa/qQN4ZefEusJN76emQwi1pf8UnU9Vh
BpPbhHO2oqw2tYLNZCF/4smJ47UBqp4MwztB6xL9hk9KEyub6+OL4kgJk5qZmqkg
z66yzZOOUB9XsNi0ZtXzraTG7M3sdMHVbut+mLSN+flYb89M5w1iojVOqiCKiUgW
+QjMFw7yhX4HRnk295x9nrSjjnMzHBIdFn76c5qBATnELhez2WEjJNtAVyFA4boy
zcDYbyg/TC3oHgmOyzflS/zmWAiZdoBvBrIMGduN/6n5ESQPDxCmpDM/zFNilDNC
r2+YVEDgyiGhyuxeVnx/I6ULXrlueKmZXZLA7ztBvXvhm69E8HRnA5NFehueQFUm
m2cdITMxgkzF08hlGtzytWMhtfH4uDQ9bZTnUe6CixzLqZIFX90me+LIgLgv/ziH
STjSw+F48sc5EYw/ISnptXiiEOr1+8k4B4R5PwExRkvMEaMzNJtiG8yJLvBKtv2q
uQnfll9MqzFgNjqYZwwVcq3VLIPT9+X9jrEYdSfVc2oLX1E7MAPyDlV688eGAELE
aIoBk7VmzRaHv7ApA0SamL/MmCWD0EVIoqNm5tv1X1RGGX249o78GioKxCWDkFwq
vQRPxrJFC232ERDPnNcySmHf5VKXo9yBQGrD2OEXB0iT19DINjgrYi5MWG04aZHS
klz+H95B5KBZzJgnplXebE7i3h+1ht9/KE57z+MsIkk2TSxI/rwwEcAyzuWGGZN5
wIjSEu25tJPwRAvcOwwMjvfn97sutzxKTfJe7KqyJQfclFDDnhrc6SEZcKvUJK+L
awhc0crG2mXJoTz3vdiadQRrgMMwi0EtL59RhBtfYDCGnGLQoGnm/ougVB7euskm
WL1YM6pZFC+QwCeSG/x6vAgOu/r672vgqf9zDESzZaOBI5MZxbv8hSeKraE72jhE
t4gsv5DMM9z3hKjOgzs0hfgXhG6couKSEc1YK/gCAfJgS0q/7y4UasFvpokE8NIk
0uuL0p31ik4DWyj3lnQDSkoFDsKm0RMcJCGavv9DsAAOGXuz5ZcWZShtctrYsdBD
J65fy9AOWAEmkxQZAf7xGPjtQq6TdLu4/dnB7wDOQCDyOe0SRJ6KqDkXoYb8cQhw
Spm2XmQpTi+l6ti/B+Jz2BQdYoQ3VKfeGsTLLIg9mc1MSJ5timvwWyBjlduyUbt/
EZsSIlUed4/QGVqebCjaHixPcTkWlljrQiV9gWCJIAqu7bsNesVg9mVLWqHLBxSz
2WbsBxQw2CmeupdOp62aQO/D/u4mShVhtjBClaoZd8cXAIEHw0CaiGaJvvQ24HpZ
1E1Btwi4sQUakDwUKUQDk9by9ILN2Oiyta0Ko4rNscxgfrnAsDUub4yp5m5SPtbn
E0T+yqzyCOceGQU0LiGeR5MqrU5zjqBXguphVFdnj+hd/WwThZ7FOMIZ7wERUbkJ
mK1dQTL4wkRLDPCMDk/ud9xf9qkBPXToYl3SbKNB3Hm6NmaKk7DXyih70O96WUK5
/EcAdrVWBEA9lwA63LjGC6gkJHSjqibu9ZcrdrzQjmt0ua3efzHoNj9Mlll198ac
AHN50L60rMatiziSeqlgE2OSc45ArZ+f3RU4yfrGCIg4x5it37z1tNcokh5QIFeo
hIrLDcDr2Xd32KqItUVLq01i+jXo0VNJ0FkeWAT2doV7V71E2AYRnVjoAgInaGWO
WVN+qMfKl11fZaoiIIHq/tbmnChyXaSByOEONypIxVdGyr2+RS+mpOB1taGkiDqC
eDgvwQ261xQYSJkC6ojRbF29AunfnARX5/E6DsDa0YzIy218SPjJY/GXIBrttddw
zznqVZdWDbnBZ3k3wgE7PTS5P6q42AdS53mvZKg5mpIlm+EWpIcqpmVWv1fDpH+k
mo2FnBrsTqSUexHTNIWyXLoRR5VdGaWdWH/93U6taX6RKTTuHouZFBKnwQyGVqtY
oCGyQ0dSIP9IEz+57mfyvFvxp2N6z16yCg4W+3b5IjIr+uL5Q/nVaeDkd4pvHYZ2
UmRfW+Vr/jnE64RpIrwp61NMXuLDa/UoUF0RciE9cWx6FH2JUjt+XGZ+vnJyKw3T
QTZPUhs67q96BGp4ni+u5bn0bJiC5ShEtHePoigIaBIPOudnBXkXgbUWcjWVAwmm
mZNV+vDKtaxgT//pKHA17N1yer9dfC0lSnZx+erghObdKfQMEBnT2lxVpc0EsqZe
la1SEMJvCD3tUa4uVdfwSiLbFYyJZze2oWOlm8jQU6chWO+N1BEBwhYIj+y+8zfA
9O9Fb9VPOShWXCcDMLG7sHQDBSQuE/LgI37J7fIaGhI3+Ucfwr+BcCWCcD8UbC+g
DPaqJ5brk2waCbBJexWCzFIDDqGCF3iZlqsiI1Atdb/+SNfEMy+a66LvSzpA0Dnc
nugQFQUmt+Q6ZBJl9B41+r3uTbi7cWWgVjCVD7hS4bkd2jPbTVecEiW1hr2a+Ucq
xhfaGR+8TH8aaUSmO5X2ndYAxmMnlHsM5g5qXDVCdZO5AfL76G12MFeQUJ7M6Rp1
dHf3X82xGI/bQMTor395JKCLva3VRbTrLqzT+t47dd8TyW3o37L9lmyHlIbtGBdh
h68EMnKob+ZylbrQIaSkXWe2uRwmnHglO47Qn8meBmb21Y+5dHKN47cNykZ/pnmh
n0KuIW3SbKaPux3rgAbq84cVRpDKkhIl/XVSMFu488bmwdV81C37xFUR1e2iXeWx
pr2+18L6fFdlaFsJkO2RS5dsJMhrLwzpOX5QrwJjtuvwxAmbsKAno6Ootg7A1DLy
GV558IxCEr8c26rr7P3foWIu94rY6t0/dA7wQjHftcpSpjtg2aV4IIsDm3bh4Ep9
etdIeHKQA4e5s8ZH9wLC6y+iNaGyBf4/P5cHXUMMGuVDvWxMyd2TURDF0nACRh6w
w90QlTDkk1TFKVODGIkQOLdXZ8ifgeHTem8O2GoYu3MBT6UEyggErYOtk5yNNd1z
/ba1c3RpdtTDK6lUzhBsAyaXTmgl6W392SoRll0r8PYNu6uXb7Q/xLhfGqWqnWSr
rUbjrXvWMqR16UA58bDD8uFphgY2IsKEQuL5zAo+3FkFNXYW9T04dcg3nPUZXAOT
lPINdWqgeohYSgp2zY/ebF0x4Vgp7ctQX5I/EfBa3LUCib8tO1+Y8CbAze4wlpv/
hAvePFT9d2L5PfX7Q0VHdQo9DKe5GLSEb/7bGmK+Uk7Kor0d8svACedUpxgZMaa2
6MRWNFfGSelh3jLe78MEpYQpGjeRa/uB3fHwBn67Tt+U9tawNIpA4jgYEfk8ddY+
u+IArXJFFCPnFD9HvPgVgQ1sr2BFmJBHNz6iENKJbx0lIEJacjdFmtEp0YVXh3Rp
eeg+MtIwii46f+FwrwASfwBk733JsGWmynpUstm9e9IbxVf1sZdNE31fj48PwWhK
pQiqJ4pM0Yqfsi8hpBR7F8Pm88VJgxNFHv8VJxo5hbV0L3ZVlylND27YLDwMGC72
X3ZyPCczfd4R9LoLs9vb0iU/Q51VrE2Jbry1P5uSgbChJ3V7oKqpDcbAIKkGNayb
vCrBQHlrndl+j6BUcOfGhviXShpiXUZIJq/U0qbFpvTLoYiBVs2W6RUaaImVDR2D
FQQfrW/yFMfdVf1eUnrs3OtwX3kEzsJTwx32KlsWTdQ9j7SjQzC+E5ETSh/CxQE4
rl/wKIBL3JixRiHTJehnSOkJbbUezXyJY0kFahwZ9iS9Ym8Ou3bRcCoQANy40fcG
vcIAFcKiQS7N311k6Lus6FLw+F4LrTI5W3mtz3c/3eyOhRfjlg0vwi/Sd+hrxTHY
rJ29qBIqba3GUhl3jDea/tQdXJi1Xz/pyAP3HxbXl4km+QkBtIqvMNv9Vr4I0fQ9
9A8QByPstDwZawb30JAqha32OcY5/Bw/OIzG+QKB1Uh3ZXpU1zp4bjiE6j1IsByZ
fZf6MGK7m6peOdWB4Jl2zyMTqafDMKgUB8N4Zh8NxiC6dkDGmfVZiXOXHcZhaThq
hAfxfO3k5K2P6Ay4EnUwFuw2b1lITuAQkZa89wxQ2YWeTJnSQrsNt1iMgOzisflg
8Wy6REqHwJLzgoLwwjWdkKLPMBcwFJ52rPnN8LbxxHzvTActrHXfJXlaO5lgtt8q
icveq53fZtGD0CZJKCgWU9JsSe+lnCDUICEAqXSDgnseTW78AQaivPpd3SZ62uIR
XL93yr7W+kiG4bwY0gXVOw0g/nPx34JzL/slmiiUBWBPmPI3Cs2PZ4Q6rKWEdYYm
LZ8kop+Ez9TX1D3jD/mGm4/4xUdk2C5mdps8oBcKw9cxA8lPS5uS0SWhIWu2bqQT
On5YdBn9Ip0YP4ch1kZWNqLPhwwUIb0m9YWMns72hYNej3jqwyT1z8LY38kHyY+N
d0GLIj+sHvZPHFy0nd2ISrk8Nb9gSpj2CRZ9w1L1G3AX9Q1CRxt6A6pozwedv9yv
YHwiuTgvfvtY1pawVY39NW0o1EmUipFWZBt3Ptxk3k8IQDZqeUr/o6eTBSlrK0Tr
DPquiGNtYYNTHzzTkqNU9eynpajLwJqeNLYwsegC9qmHBrwRMNJUH4sakmTTgylp
9IA19/uZTBAxkkOjv8tCZx4PRb7xKV+O6yzYERakvMqEJB5lHnscpF0EzcM/zGs1
8tsyLdInaq4wxgWvV37dPIw61IXHckOHb6KYThVecIDnkcwkvpG9gdMZ9IVxaokO
R0CzjLY+/EekjL4/33jI809/8sa+xqsL99Exf49+9Wd0NAhi5KNL/uyDJOVzG1jV
7dEJKOqZebuSDvQ1EMkSi1gPl58hG6VOfaTO8PhjG/IC2tsWLg/jGXFpcVlw8cAW
hpYxtdsxi28osSUyS/NiC3dd1c0np7JgJ97zFqi5uhgx5T43e5IcynTiDXcbztg7
7IU7m4rrlWW22ENIXeitue0rHzFTOrmWBEKsmCG0frZ/Vfi3vi/OIBwlFQ2z7cEg
NM6iuj2aTJj4LlJzp13lIfM4mwCVBCsE1Yyot8J2I3oOGwPKnB1zMSOA36w21SEx
7SMJqVHcPk4QrQanBuo3iVdwu6mHnrWGZjzQ8hV6v/77zR7l/zmcvSAb306A9j2Y
Alj7iyLQpddBbNYeFAV1MhHo3yp/CKOeaYZ3IpAG0zPb/p/6eXE6xrxGENS4Hk6o
SNcOseH8X28dhT/ZWBnxscSOzx84FYuBS0Xt1Bq5xpUqP+QUyFmRAdsbvjcuCBIh
HFTJLH8557wSsvHfnnxlfE8b9HnMUgctdiGZIiv7dcySdYB4Bz6t1wn2rK6H2MCL
4fXskIew7DBTbdZ8a1bw6sXZNs1kPRLyozLVla0C1SIURLzEpQ24RwQFOOBQAV2K
xNwYFsG2A72EJxJQkIWFuDZ27t5KHAOomAPZwYOlQ0WR96Bs//zf9en91YM+r2Xj
Pj2z8jvihnOSC/aDssHd1L+FGuuLbqzjVzNsemggi5YzpFVgP4JBJ6YHAMlbi1nY
4JYVbSzs42KA6wbHvqpcM1P5bcjIT3cSQsOaer7zi1IG0EW70dSgF+6z2q89Wm1S
CXNsfIAm7hwSxpj5Q+ja5aTNqToobNJwECvIaR9VZwGgMj7JEG9vZBROx4R6rOLd
GBtzM4szAwOcuQHle0e5jrdg8THLj4IDXlpgZjVnvZd6N2hz/tYOq9iGpIR/Mih0
Vsa5S24j7Xu+NwejdQOh6E0Doqh/yrfSJXSUKaRrCPciae170Hqsy2pWWnmeDigI
KTmTCDX7G9JxJo9qoL4+vJZGkYczB4BFYj+95lmLD2+emq89yHsjg46nyPLiZd1+
TQkewJiNaudIFsQx2i1vZgEm6nNXAbgJ/8hydVSao79QFhAWcDJC5RWpS0PATmiR
nOje0hz/yZUihJ33WDjoc3/E6vdtS4Asq++ynxmrMTpHwRkNn3dECFapp0lPLLmN
4skLb8hS9TnWe6PlunGp5rzN+u6FsrQ7J5BSTiV54HmIdl7Vw17sUZ85Aq63PAXq
eBLvWdXIOZQF6VFXTfU1IwXU+21n7BA/QaWZTetW7dbK3XNG3Ji26GjsEEpes76q
UP/TIMKVSsrgBM29V/L+GEEpqXSLxb9YCY3sF54DFcIueQc6gGNKnFV4AREPRNCP
OJi2Ja65XhaU5HFvnGTIT8JF57yyk5Zb/He3P4f8qqUp7vfs0H+5KUCzICV2qNCU
O3V5r4go9aclH9Hd/WDLaVQshzW/NY5zZGNoJfNrmqoJhYLF2Ne6JBv6oILhTiFW
7k2qMe1SAZ7yoQcc6pu3E1+hCSaUGR4mI6Qu/ppd7rikXPVxktsxY1tSlv3Q1GKi
0asM79SHqobqIqkxduCUvG6ipeH1KUILrS8zNME9ALqDFW2QeJFCma0V+RUlrwTM
ICqpbtEPpUiBpykadgLhtVSIOjmf82putL+4oDDK5LzVPxk3Mh8HwdoGeht4Qd6m
++OBH7fvDgDDKOmdRvYjlDM/UFuoB2e6Q4GLoi0OjRTN25nDwQeBP2CxJQ28X+wQ
ABiTRj/jzV+i4KxS0PxFRhNunCak0X59L0aPKPiOfjuDeIbTuNZrDmBLWyGjbAdP
7mXLPpgWffyzQcBjSI5cLW4EsrwqyZ1SsCObei9ffdxxSH51dv2xPPIlVsmD78qo
fJwlpW4oNMJScVVheV3Vi2tCotsquF1smrvecubWx/Fdc0yKaN/2jc2X058bc4GZ
mAmo4m9f0HhTu1ZK7c/GkHKVVWvhEAqGgxx0WbZ8FaFInMnAfnjvlAk7gqBDPHtx
DURiCMec8AdjUrwiRP2Sc3Z9J3zMJ31a3vz6DDjkV/4slmY8pES8y/teJ2MPyteV
AH9CFeZokvwjXt/GwhPUci5bjxSOjrHSbUI0WpA3GyFBPVz/zn7R7D+3H9XooKhl
xeyLqDxgFgE+woNWNdEfi4u8YYdFKV77BOP/MPkTGJrQ/vcKXCOadS7MSNoeOfak
sVDjc9XnSUok5wwHZ4jRuCTXac7ua6KTOaXLpe/y5M+fHCYC2qtR5VCYemUdnsK2
bEGg6F6CXyywsvqwqT7lwb88QfFYPldaD9bff6Ot+BjgDxgND/oBm02VEU54prlu
ZYFrvcS+4AfHHbjAff2LsGryYfk3ByYZiyYdHKftvnysAMA8ff6l4WneLG0Fg3Bg
NStxekRdPlFeU+sZ6jxDDHg+8ccE98V2Tp00GTwcQRisHswJezb/kONBdMjApV+5
1AU0bS1vZ14O2kftx8RbCGfBfbCyT58P8KdRNSAnovOcx18JnwUjVQ7zrUgwx4z/
1JcI3wMcedB8cUrmoR07sXnLVCC3ZxYoV4lvRg3h8u7gtJiPcgnFDyt/Ew+4Z5mJ
IxXv7KmbLJjeQSAwgCWprxBbo77X4+FD4AFEoKJGTJM8gUTWc1jIvyf1lVJNaENY
zFTXmYrt4HwSa0qvYCZ71rMFmU6DWrydaCwXN2/tFJZUf9EhTVoaAGXb/4efVEA4
OXqDKU7tmKBoeozy3sZSmxRTFNPwM/SPFJ0CunHdbEdn4G4p1vaEMU6hCNTIz86L
EGz0R9dHriCPlJlep17ejBpHdGscLKhYAEnafhIBlv3+a6TGmIZvPSaZOwh6klg+
lBzlOGK1mu5xhQ4cLFt2/z5N2lsxf6VwGwHtPxsSLWePzbIQyU2aO4Egi2c6Nruj
WrPt3k2ZvbW9gl2ltFKj/Gytex/1ARQTxIjjrSrGRJ3dLitzNJm+HpP5qzwpeKFR
cCxd1Lg5UW1U/a+7Zi0rl/4M/mI1h/5e/TQA2r8Lrpn0aUkpIuyvOUw4bsuZbEK2
Y1bxVCRoZROw2xd9e8ff4bRFadggpbzpZQjC00X5Xi3UhMq76k8jCJ9j/UX5wv08
D2zGrI+Wx6L9anIBxHOnR8DzZbx/g1LmmuLt+6U6zFIKX4iZMXqzd1wU0iR5fkSZ
XFi1+L+tBGKVY5OO+KU4uW9j/bszIh5E1tMIUbEFKnbLd62p6LguTkN0aSp7dcG9
eucmLM506R+wcIMoMQ6bVWiNsLmj3UcjMl3BOVYAxUamxMy063qSj1rZ61pEwr/h
QsH5bGb5oT6RfPaGvqVdLdOfVqI5rPnauum1TvFDpMIEyDz74VKPdUFZA6N8J+hy
OWW79giGxVgFZb+BdszU7aht9TwOa3MHeyJqFH63+A4RXJtSGubmgv2mf1Q5u+O6
KKTjCNgNWO0A7T96MjdEYYcWsRtdUPyYLNlzmYn40JSVXactPU6mTFzMSx2hZAFB
qKj6Xe3yC1Fy8u8FFaEqtb5CBqgKav/oe64qQdqtjGQOXhkyKJGKCINmbbNY1oZf
CgbSk9aHY8yt3039/AfpY+eci3jhaHlj0hPL+/ECgDSwatxFSfbo73P4ViJsuAQD
PqsFHB9vyVm4oC4OOVyHXFYtLaQKbd6XhY/Tvo/vBBNy2cT43KMeJqtdi0MbV83v
q2Eh9ITCuemC5FCAiNNH3tGug8DwgUh4+0AthKAFWwKs+m+7Qt4egE0/+re4Ac6y
Aa7h316jBr7oS7QkKzMSs9r6iEh27PK8QTAu/Q5kqqK7WYlwjkqqRoEZ4icX/K29
cKutL+QpL2kk6vwTAKZRBI+ycHbB7cgdeV+bA32NRBhSHuXgj3h5gJRZ3i/m6ehX
6iePQe3JcIl88lh/HVklkeMdI/gf7r8sBUqEn8KJmFAIt++s6IIC0ER0bMnVXFB3
7GogU+rY3uA1mXf2Ewbwz1urvLvjm3XMVgfFdu+wV+XXwUG1uhAyX54wj/5fRFLq
+shY4+5g6aOHUp7g7CN/RSwviTo8cPmw9rH1osO1DO6kdmGIkZnDHA+arEQPJqmR
3KxPHgvCfREis88jKyOpCeLassi/zgadXZrtRrGp3eN8XbPfAz354g5KuypPFPBt
e6XGNcFhQm/QlIyIkXshuDJqufhRC2TUAjyHzFHq3IFyvMQlgUB320qXaREcCqNF
HFSW3Tj2KgJjlvuVtsVc3e/wtlmteOiQwQTQE/Mm6+qkzkqlicnRBh8VQlIgOJYu
+7KbmD0ATLV2ZmxEAG3mbLp/osQ3r3e/IxZFXbNhkZJdTEb8Sl+hp9NICTTW+4/M
EWF0ODrisM/prcuX9Y4P6KPLKmaVU36Fng7dRFJPNVvQlOT8c1gswX5Iz0SQw9XT
g0F+o+YjWpUM7NJocQDUK458u6wAh0KoyK5L5JlgObxKRZ1pNpljJHwAlMpM4SDE
MrH1SPW/+YKiJWs9hE3Rot19G88u7rBsYeizyM2pj4eslz5kuUTNLT3oFT4KVm6u
GVOEpCV21vadJjLyVh/SAeckNVxlQB++Y/+KR/mmB0MjObyxf212psK8rFSETUAH
IRGhvmmd+RWlA8kGV/a/d048Ey0gvd2ssyvKr4V9HNPNNdIYE3rEKdlI0MmC4WIP
o/FF7VI/s7P3OGW1/vutnfHQWvADTuQ6TEWw5zQpQl+fMH89RHAxPRRd3sfDaacM
kBMPA4XNdyMiQ0TPGe+gsdZ8zlogyfnTw5Q7YDVF0ZedMatSn6h0PUVgrDUayIXb
BbcoV7VE915MS3R+Ro8eIGP/4dxkBW/A78EB6ONhrwsCgmG/hOffh/KZZx3zv6q1
fFvNkorpUoLOeXipdf8LBFlg6v3bWleq/EHsIb968sxAWFEcGgng62uIOHIpzd0m
d9sIULo/aKhW5hYHJsV8O3/uW7leOaNPURY30i1n+5ijh/JBgFLnVfPGLl88pSAZ
63xZCk9JeTENn421KQLwvvziFzcpra+jbdKbwSkV7zn2haFNxXr9gwNdKD9SSbds
jqjtF/hYLUP2iEwtFtEekbGN2Qxwwz8g0UGBtwDbW/g0yrwhpGaBWmydtUZvD+Mo
UOOv1Z1/KIOaM2y+n1DbCC1jQOYkFs0opVFYcwEtb2fPeilIQNnEM2ajgUbRr/YF
qa5QJe0ukJVon9AYUvKJBnInYfN19J70yYWalq7TBzfIOp7DTMMAVwqwu9eLMD4Y
UXs1+TzbaHt/rdNs5rrKkd5v8pg8PACXVlfav7iN9NdJPvRlcsJW0YUCdrgnRTIl
gquMCacxRRdNnYV+0XIDUm2L5Aqi4Amdn3baQc+BduOcvTIgEJjjk8uUY72EqcTb
VORV3fq0gKxlf22H57XsAN8gT6HnqwB18+lPkY81mpgUJWbgUxZf3v2Cve9k4Gsh
LKVI1VvLqmvhmj02FhKq3Mi0cGOl0tQlp9BkX1SXyP6VWVcNRyT89CFOHg7lqjLC
9uIacoRtbqGOhOfZOIazb+dyL2BbfVcA0gXb0OwQa4G/UDm9I+VHTRTmO+AVA4ui
JJUj7E1tkKmbCCIzuOz4TrMwEIhpMQ5kg0lXGXMOSTdFOCXnuVaSsaK1BnmB7hWp
c6riDQ3rczXl190SQSWvdCbbMQlHd27ygQX0mShdQUtzZbaWk8KjNdKE10s0df7Q
sK7mASaU4Qux7ULqX4L3WwJXzIRlBou7v41lRpJK74gkE1Pthc4AObvX22/vrla5
UZR9mp2v+vjrnpaHVhZcMxHgiy6elAJ0jBX7NfV2XDhG4LR+OQ8abMPK1lvojBVt
YuoL67dKRsOZDEKqVU5cqiZ3xr61FjwKwPTKBysHObDw7jc1sn5PM8SJV3Zu3fOf
/Ewd22n4XtrqoqQ2shtiJoXC6M90YVg6PMwxg+V2D6lziWzCgmYRv9P3Nil0GTjQ
47RrXeBjLFoTvXQ+916u69wfGObelc3+SPzet4mMBydCCLHvbZiKsbMTky8rHEBW
W2iN4HwrZs5+8TmMWCWAKd4pLKcp0S1367A9mSp7qclrtkm7gwyDsUtjLev2Jvj8
qVfoJM33pI3nN9BmYz9ZKii3jjIHiQmJSm6m/uozUJKO37dLe20d4605dwMzud93
5qQYUL3BbF6FphFZ8YJvS6W/RlnYM34YlwmE5bTIm1ZASLQ4NbObzxAujI3whrtL
5zlBqCxTbHpcqoVBPWuhZHEDZywcaq7V+2QZGP+iQV2i9LgrYEQiuEs9orcJrWZZ
bnkwuQywitb8lB44yTlHXo8XcIXXNQWa1HGcron/gUsXCY3pJkHhvGlWPgtvEpI7
eO3p4A6eUzRfwE5HWH3yW83SXCGVXJoiWOPg6RXXg2T8pIIdwWI66ni9q6L8EciK
Nu/MbJChFaEOOLICDPM8Z03ocF2yxZlY2iXGU9zaamn9C7VUsdDCJPU+30Sjy6zs
7tctT3hTYzTpYxv/7YeT+D9rb3xKnWJGtxBht1vHHq0e0A/1NRwQgfnACwT3XgwP
Zi1lPCo0TjUD4S4rGKCxzKDxhW+gN472EswP3/lOcLuQXhqxCeaF2Is6QRGL9sU1
6c3o+MOo70ryRXQTfQKJb2pxCX0B1RLtZT24wgcMeQrKM7z1JqrEPyKEUi0S7Dj4
hYreMTYjFtUUSyYiVMANCYG6rSE7aT613FlFkf6wLeS76Vg2nqRXGK90Z4XONRpP
15QVEUBFGcf+W9uoSgfG6Pign9olvUlQdh2FWivCgBvzvGF0/qi4TYgt5jaoc1zb
5i6yyY4bTGnWSoN+GdWmzGkhhzmlOP+CZ2Hlq63WVjCtC6/0wtNeEq+KeJ4blSSR
DjMjf30cQd/OBR0TWXHap1+kXrD8wlIDz+qXQTi3rZbJp7JMYfKWfcw9DHD50wKP
kTSbYqjgDelebghD5pGC/z/8KyrGndDT9Zkp5KqPDJJHgkrLZUTqvel0lx8/8Nft
4Zhd7R0IwX2HW0Bg8ooc0I+Oat4VxwGhhaYENm+5jaSq1GUUhSKwy6Cta+zJ8puH
iFBuX5s3W3LcKYb2rj0ioQmYWTzdIlL6OJlMWjlQGPp1kg0bM2CI+KVxJiagRW4Y
lQmYud3z5V0DCeZZIHJeqLiENcXm6jdsdSlEw0dT9jezB7JiZoyRGYap1OHo6tFQ
MinM7mTfMAlZgjuJgM2xa3gqLGhTXQHX6N/TQV/YSaGa2aK/UuXXDCk7JkxYtR4/
W+El5yTb3wDpwxDjurRr7xhUW8RPH0B7xdnggnw7NleHMkhqCIBBN+7XyZSTV7U5
soA8Pwnnm5ACJMoj2aFXzJGoiwWYVqNbG/Qiz5OKOqbj/qaGqhmQg7TsGqtdXoCb
tBXNfz2i3P5kXMrKqINnHEuCvbuPk/aF3HXxW/9I5KC56NP+BD5jnsvdcXWEezhz
lxTsOdrEekBOi5UrES0PggZHWe5Ty1AdwtLciMG3f1G2INCkrsLjQVPWidAPk3Lj
WletNfXtPS0Uiky9cOU2/Qo5VvK5mHOiOu33wVmpOy8EQaAJCmFmJtjwKgUhQ1gq
eFfaqXJsl8b0xgVSv0XDqWCp9gRnJXKadZo/F5QSW1626eSzQH+qPwwYGmg+t7Sr
hMAQGDWY4G5/KRG7ZsMFRyeDxEKTcwKFF96eHVA/Pu2Tbilq9TKZUmD8Dwq4+eOW
Qqadk/OExjg1N0V3SeSSZd78M73ZBl6SGzfGJ/+c3eHFF+9Tpoftjgh5n321lISf
s9YpDXqQA9P7C8ZQ/TsiNlo2TaumZ3/tC0o4MlRuZDXrJl5mSGfCcxoZDv0BUhkZ
DZACnJMoV1Sy3rOt4VT9FKD8xNpbtVMWquI26I9DviUHxCAmdwhVL7pKVlnZVVxS
ohyU1MjG8YS2+S+Jp2Ras1AwXUiQx1EIzTaJsKZLSMWkIeTqCyyn2JnharviFxXi
lNadw12zJBLh6sDhF8zS68SMUYtLVAFDDPKUmz4dQaQ3BIdT12mHgZWu5JZ+GQz5
PcmcUhgIU0Err70QvLXZKyQVznnXmBR2wPmv9u0mqytD3LkB5kunTh8+uhQZaUOm
oq8AtO0yEtm8x7Y34QrW05kVjPfAL47Gx4pysolFv3LL8T3ATyA/qi86qU2kh3jh
ZYLYSVNQ/rrUqKrGc91Qltik1fJHE6H5OwSPiIxRYnGgD3yapCvo3oImgdpqntTG
V5+OecxYTbsQc0GhhHl7EuukzJ9HW7Fj1ykPAc7oJZvicWHA1uch7YQiaee2/6uy
VT0Amh5TAmocMdIVtSpaPhnogQELxV/Lxb4N7Rs/iTobqsLvdAaqu+BuL5/ZteYW
UPUBm/z7KsFRt8wyJUVNQ7jQKE1h3vHyWiQoMHqRZnTvj55oBebbxGUPd4y6sf7b
rfvaDvRE7rpJV3Gqs96dgooAqOiNL3MsOPWqOy3OcEi4p7AeQNoy/uMPjNnBbLt3
YqcDoGJlv6b5yAeQ7NxR8U1rf4sY8f4URMCValkO2hRftrnXzzLAZstOWawprFvh
JVPC8s6J9ld6CO05LRtUOj6E6r7D6BcYLeH6Gl0kyIFNnwJujG6XIuBP99kcxuNp
2o8BxRUc/t3CIf0WtPiinzd5nqjl+DO6o/POmvusJ2rTrIxZUtYEY7v7OLm8/hwC
hCQAHSfLSSM1qmUFT8fJIyViHK7w31Hr5sXAWFnGPH+yhfqV1GB4s6Kd/5ZqsZmX
M4tmW6L89qytLhgP6uzXZ9xb9DR8HwjvwF96ErZUaGgWNA/FfIaLlJ2GBU5Ix7hn
OyI9CCvqKPt1MhkvshaEYu2oX6b6QfeBjkV8FQnW/A4//kCap0O6GhUktJ+/Ml0v
7UgfC2OyFZwxGufCCQxqsqcqcCUbzmn0IU8GOWysdl5LHnQ00/4ElgCT4gOTmnDr
jBeVT1WbrNeSDkoyPaxfs9AhahxbhN2dHk+5OhAh0pKdcNzTaAIVAg2TVBbcR09z
B2cIXyJfPOxrPeM5BF7ItO8GZFuRuI8DxgrYvQs+wnmUV1n2e33F0Nhit+iKKZqj
+ZZ8PsAzCjeg5eALyEAPHZay5o46RvgVlvjU0n5hxGTWvaCWKKnLEvfb+vaR5zzR
pt5ARBP3ye2rf8FFMy5fCHFqXTgCKVPszOdZKuTYfiBttymVbQE+3f+4mLsR2vzW
YRnfFCTxPzGKfcIrzK/AtUnD+OxYVvxoMX2gFIc08GdRd0l+wPiJV/zF8g4t5pGn
A8oLvXOsF1/QBfIFtkJvLy7kiI9wmu3tdqaqww2oz3XW8HGssFnIkhKWch/Lub8a
eYOr06UeabQld3UNGYpybjNDYH66BFYbTFICJwuAtMaiOdTfGHehVKnJS0V58hIh
Fev7cfNKM6u2k7DZfVKgqtAQvM9PzjRfblKnsYGR3ku+pJ6wWANcUI9xt4PTO7/k
jvIAQ+rqyqNg6E+gYqnBjKEuMwbPAZpVr0+JXyoit3d39Le00QqgvB4gM9BJ+vRG
2QCY93LVNV/8oGNkKLMJcWnqnVWPSVDA7mBI05Vu+wCSstS39XWfmLGO8arCll4K
CHmlhHWkn3cCxeXaKgMNz/4FYtrLPDf9HHwv0tOjxOvprWOYlijmVV9OQAVNbTSm
1mjkh0Twqnr10FFWnZkiIG245xEkGIgRaxTnG/0El9c2qYMuUb1DZaHKm4kjMsrb
EJo3YgjI4LmEM5ox9KSAcPVlUinjYcJ9kI2XJ/GpU+pUMkViwSvC9+dr7WW6E9dm
/DrkwtAS8eH+OxDiaZf7rNY/hxDKgt81xpu/lby+JIb94fnUA11W9pRch5leAUd2
NLGNjOtCE6C0Z3hg2kJPYKCPqPvHBZHSyQzKebkbAJgC2Wpz0VOOfF3xJWGtjL/l
TZ9dZog/PVI2OfTlWs3RWfs7sdRlEDZpF1eoA2Mmlf4QNkc5Yb3W81k0sPRH/6yI
tSa98Z6O/IJAubjm3ZfmtEbCR2GVuVYyWisczYpCdmXUa0lelWNCXfvAPZcRxYzj
rzLE2vh+nRJNhBWBed0Hfox0Q2yC8DK/xZTcpsDWx8OHm0KeiG1OWeAeg4V/7BZK
4siwZgk2rdHh9y/naWOYsxduCV4WRaxtu4o+/GOa6lBU0ffwNw+N6+RR4y+vX+RZ
2USnG0bIyTUq97JC610eXTsgg/B19nZXkXk4m84O0/co/0bv8o57NqMyeldp0Asb
ycVYkUb7Kw91W70MrzNePQBPhi8nLRRLLUOBViM03d66hVmwG+BXONYTXX/Xbjqb
DF0by1X/4MLkPVlfMQ3xoB60m2rRVscwAI/Ca7+3EisUGY7786a+vA12qivFZ62H
OHWSkKFw1OUKEZe+58MBGn5QORduK9KKmJ+pci8SpYLPGwLHWmbvmdWY7u11775J
mZcYFzY8ntRgD7KH3QGPnkQmpOb4w5BrTHTXBQC1HkwIRYd4C3/hLffYAqgrY1XU
5Qui/r8Raaxp3AtcaL22QPu+jOgvGSMkjae9flTTLIO8DeXChqcOLTra58841oOv
5A0wsbgttzQnVq7L6bKxY31ea2HAC7sNBeNlvZegKv9yO4CwIEcdqf6bL0z3t0ds
C4pRAC+NpfxWjLVYwkffM8RiGhvMlldwXRr+P4PgQShvdbmfPut1QhpUkuLpOd5y
mfGxo5guLgG+IigLAcX0Ng5ULzCvfSjGvIfpiVoKC5+DQ11pM2k9XK1yGhJGxcpz
PD67dYgREfsBR2jLLoBh1uZ5wml9m9GmPMkXlLi3kqYMU+hxQa9QQegqSq0m1XX9
RMo3YrBkvFLEuToW01wvRPoo1ibF6baYgwihu/0CXjyFt1+VxzipTcU9YOPmDrOD
6W70/b0h6ZzNDwoByEXBRMLUFUuFO5zndcvuA/ES9tpiq4IIGRe9rcotf02wQJU4
GiYFgFtBFBhjA3MnhrNBk5X7D6GhXuiW0J/p2dCG38fZ9QWWoYSob7/lKz0MCz3x
InNqVmOWL9baavEvam2+EepyYL/SlsA3jwME36xKnZpcRymyveDOdxY/WS3xUqUr
mNF/3WIHt36VEzb9VLQmE8dK1qAt5rCfY/CfE3w7rAN12iazqzZsxrlLZayEGxyi
itLq7PzlinTDXHaPNim0fDgjl0BKay546shKbGzA4Q2pBChi8JnL47NOP+ApXQyI
V+67KwGUud6PvxzTPTuyrmSciB+K5x3c0zZ/uKt3/7xZZjiADKyLs1e4CjM4cv+P
2i54ZWwXoG1hAzV+e3+IKCF5IWofqa60aLdvC1nv+vBNwPuGlFfHn+XKPcihXzoY
TBtpUK2k2dVc8rVU8btbv42HYt6eZCRo5oUl6MvKkKJm9yVIQ/FFuammI9XXr/e4
YsslSmWpEQz2G4kk6GCYd8G3E39Jb9d6Vd7uDS+3c1Gosn+1paUP/7hei4lIo927
gs9Vf6mPxi3P0dzAf0SEBSE+Sxi5zreldcJiln91lm0yHmqPAQkMBT8NM70np9TC
3gui9K0LkjBQdbb4x/6pQSI0PZy59cCmA+6jp7gQUCq7o/XJ0yMEMllOJDY2+uTN
gOnGhkuCuTMocUPQC4vgwlkw2XQ1gJbJmOBogpf9ODFlT7ycc6XpWAzuX/oPPTaj
wAy+3pp00snr0iCGX80OHe5WQAQDuNwnez6JlzSkdQeTEwLkg162ouYmr5fgoH6V
I5F/bkYPmLEQbuRrVGwcEopO1iRVQm9HypXpSFlvNt+sFlIn3pLeW08TbJD3VU3F
0zBgkCCB4bI6B3Eu1VKGrk8eG6b4xTTVcLJqN3CiaBCspiuytnhME++CWJtCs40U
KYBUh5uwoekQt/9qtGd8coFrmUARIeY9va7WUyHyZgAvDcL9uiK/m/xD71V9JN1U
7ds0fymzl9itk1zf61LEIxVmChTXkIFKYCynVf5VZ3U2FYwTrkVrjCIZUt0tNdJl
u8Mv6Dul/meCGWDMM87Vpy+hiIAFXQjD2N9TV/2nVkDJBh8QAlPWGK/SWq+nlkVb
09wP5F6+42sbsN+n7524sNYhWsIAB1+MrrMNauOrDi6LvtdIqJaIhDX2OGWm/285
w96Qpu92Nvlah6xHsUAEg//S2TyHN/5tIMhDu+JAw2pv/qrndi6zAZSNF6uvzHiG
kl6oi9k7LTdqb87h5FTc5WpOWkTJH37di+1dutUJXAY2uile/GC9nuUcSDPhldN2
LtIrTZGs0E3zvWJ8TKTzugOvX3725mn0pM1R9frdChIRqZkAyXiLBx7S2zMc0dm1
nOzS3PbI5ASSzPBtW9FTQw1Na3Bc1NzQ2NR3CfZkcH0cPecFmn9kecf1HmJEk315
gn02AF6AXj87ERJItZHeE3piYReYo0gkjp5fYwnD5vY/10JKL75SBhpJLR4WoG5o
090VuYiOhx9/mKpcJ3l+0NPsC8xAnnD/jrlW/MJRQDuIWz1EgiqL5fKEh23E2vfR
vz75MO6Dyciu/Z8Sg4L469YgSf1tV70ia8ZbK1+jxpZCL/nfT8eJa8PVJWVmuNLD
QCRZi+MLIGL+DceRWekr8Vd7XgzFGM5td0gpHqWK6miE1lq/nqaQit4QF/XoWxBq
1ItiqSMZUqJsGl6adyGqlkDrOpzW+lnIUP4fQPpnkPQQtnr6Eh5bqNJLqqF/AM8O
/nISIE1I6urI0rd4rfUh5jy4pDIU96UIehVJRDU7f6PkgGesGvDtZn2MNOr7WfTI
OG/Y2UYLiZyA62H+nOLi7fX8gRWA9jyVEhPEt9eq9aZpYysrPxLrzC66I+3q8mUm
CMVln5RrOx+Rn7+0bm60SmHkplZtgBiRLGx6WCiEwgWNifOydNYNMnAd6qeqHV8c
2YrdIuY+4d/rd/m54pIQ4gvR7JAe51GT6KfL+JkKvFwq50d4hs7oA43ynY5H11/v
bz/Q319XtRnhAvnODsE6igjlj8CDCiyyvQhceOPTDILyTDuGGWSKps94NhSsLv6e
s0jWR5DgHN/1UVpgc42yNkm0EXZsUo3k3BtVUuJki/3XQPfe/33Xh8N5WmMhkHNG
5930XGTNZW10lT5wzUg304EO7nhaaepJDcj+/G6Vh6iZXK5L79tO2YFZdVISTV/G
mTft8rvy81h92QltAn3G9vCJ+SIf/jlMoLk+2l1w4AF4ZrZ5jm/hCNCUuRsqIQ6c
WZxX8d4DN+Q3CzBeEc69xGvSR1M3QypU/xRuaL7tkNQkr/Gs+MeKYV3yBxqSM/Aj
tObbHpHl3fPVUwdE/2c9I4x5RS7cSdZBxgTcCv9pWjYv2mK6i7y6mb/TZINJHIpw
Pb+A1Ip0bEnvC2fl62nRdNRKMSDeLCoSJNgalc9Kd01XM1mvy9R/AgesnMXUBrDV
MejDrt3raXGwvWjBwA91yT3KZy1ly6jD3tDJ0zQHdrPv848TB9OAXwIHttQX7mg2
selQtrJD2vL0/t29fd4+wgYCEWSRpfAhDUD5XiFQl4XFrUhIX+MH/qOwxs/qGWhg
BkoT5t2oCcNKrnwY1r7HI4GT/7RzpvcZhwQ/VhhMDw7T79Z7CyeL9utkrJgWg1ID
SjRV8zj1yyWj7eTxV0ZiSqPvNVXEUD2oXGyLpfj3+XIfmYdzIHi48cFzlVX6P8ZD
Rui/r8LYUcvUwOkQopOJ2WdM0LkiGkPH26h/Qna3VPKjLHxBgYYS1RLZ3db37Ckk
oGmsYoc+TA9sZfX3i/ffaGtnv1xmIUtgfDvT9GzHmed4qA6vC7tLoxu7wYixsXJL
j7FEaXzN7gFeEh6KZxdeXsr08DLJxHOzUXA+cIiFlr3dohPnPHA3PdJDUCw2SFL4
ri/Ne+bwPs+XoKPr13u4C5NgAfiy6k7uC2XH4WarWBm0FUCidY7nd0akyJ2w7GiI
nELyifcI2HYUUG+8wfxC/s2BVKkPEk9tfNnO0bwN3CCPtHWNpJZYYwFw2m9zUwRv
pio60TY7jSWA7bhSzaU6RWxp5aR5xMBWsMctv9bcizUho78PFNZX/b4YEiPQyJ/7
sS8kZK111I8/+qsHIV+XOIu6IDCSfUchE1bqd+WbVWSouSvwLALbXeHWWt5mfP5R
G0vCjlwu2t3hSwIujm0al7QZgvmYiUFYXN91NC4NSMHrGP3yS/lbl8ntu5nLqLlQ
INsAMGhhLcJk/oAEJDRchrYn5R1qDaaIzN+enbJTB7mu5EsG/HctrI+N7eVZOxOv
aYdCEPM9WkytGlaSOFOsUUBULEJNx7kAPXRkThW+SlmyNOBlXtwKgaqIaEHjvnJA
FO2ysXUnHozJkjMF3ct7RvFsFG5A+jc+YhZS/A7rJ81fVx3nPOS5U2VTMOKGRzRs
172z+heoHANwNB8kvIkoEWpgQKF3XFPWPL7IdN8ls2/83y+6l5b6XX4v5QUAn++m
wgA9seN7iDG+d+lKdb62HghNS8EPrF0w14PTaivN8ZbE2SPm5Qyhrbe0lNLuzbTY
oMxcRt0eRaDGWRUM79HRSYwdvfayFTrvGtyjhp7+D4nHdxg+VmTMDyPnGH6PCk/3
O4+lJ9rQmyqS9z8uzfaxDTLVNuM3/ocNtBOsnu/DLeKYoD7Z6arosdDcY4Zr+fhu
ksq0B7X8coFG6EBVj15eaaFLkcUKFZBE4/fXBxLduRBU6gDbkibdc200e3qa70xI
EFH0Emq+09CTqnJi8ywVsiE2XSxvwVGSHa61lnKMezsxc/qyDZoxngXzpkvej4Ja
mzMkc01FqQZ8E2bT8HbdbWuMKdxqm53TVjTMULXEXdl+uZkAyls+rGPesKvjllWw
MUxNWbHLwelipp2ruESOHvPmLBLxAxVZXpdHARI2ED7Koer2v+AIogmkBSGOFX8q
QRpsd/qKUNaqyzsLE8Qz768HbkQShwKOJBfKWH9DWGRdyvilGeN42hT/BWkM7AAP
puq7ktGVBvqIkMEAB3ruYeyJsMZI1StOAKiTKyLTYuuozt/LcEojHGC9vAL3qyiD
VKg3SfxnOVSVPapsB8PbAawwIj14AcBCwJ8KUcvx2tSP0iiYPnSDN3spMOoOpBWF
yUVaSFbJRHN5VL14uTKFZIl0N40QKyYMyGyru0TO/Hm166p3zkmi87lYv6yQbZS3
iw4XJBZj8lrfSCQyYf0LSeEDTa7xN2Uslw52UhFJvbrA7ePQK7tPlNH2casFrVJ8
aFibPnEMY9WItV5iiRtEZdASi5MCgBNW6WsAGCLifYhQJXD47+T96PSn0/FARJ6B
XvsBnyAHrgMH8qM0Q/Tpv+WHuWW2yDUzAZVtY8XwY44jsRd04Aa44KA8eJunifJo
HKryv2eAbtjmT5Xa6CPpYL98ds1xpTMXwD75OrQAqsLvma4mmNI9Z3fqZKyrFQNW
2wMmnSdoORMkopiK7E2HGY6+ahooPUKG+SRGUMMOqXf8sIoPSrBbJ2Zm1K/a7xh/
vTefNN2u7ezU7dx6MXFTMyXsP200r0YoBQIuRJIblv6WMXDBh/dL/ntIMUsbL8yT
gfbAUGN2PAUIiSv3qm11FmhDb+o/xkCguU3vt8a2eQAQBs5vds+5z5irsHNOeYcs
7nII+jnhUXKS4nQ3KymLzsIpPACG2kUxqqIzW3vm10JUmsNzzWHN1skHL/oJtIZ2
yeOdyND0hFmmRVJjPsvVkpjgqlAqEVzoxc8ruCxBT2xX5AZIuQ/Q+5VpwWDc234v
GO7yGiuv3euzb+6cy5lHrBq+armJVj4goyMdHIUDwwMToS/dxdV0KHJo7K8M7orR
jI4d9c8204Nw6C41KMT7surkjZdqnwn/LpmKDiiOnBJoFzWVL/Ef/yqUpLAHlr6I
ZEpgCwAeFrgASutfcylgzvWyIfwuCymRb2GsaZtsqhOnPHzacuIdqowvidRRVBT4
qI2WCvJPUia8t3qz7hxFIsz7dCn4CQ/utDZbD+XzC9X+DThfZxJtk/L/KdWyCEzy
hqWetRWNX/RvvUpJS0V4F8Npd4Kfk9c2QJLAnt2jmFn2L7rAqj9LUrLEYSGErtKX
0sLAAXMvS5r9RpS2amG34c6SZAWEz9H9CsAPENNKr5SKQEMvq0MvPgFS0n/wWFcK
Q7bIY0zBn0a8cBOLhgacpRXmQcPi7XiL7oznO9T0y7ZrXwJb2lYvj9fPLV3+36Qk
0h7ZJ0bvWQA0rq5y/0DUiyUdvY/kgkNU8vd24r/I6O72AuNWlKOWeFsPLBkGtbir
fccF/UPP953j12jQf6glb8cBFS3FhPQEaLAMZERpOarMyefghiG1bQqgxC/okG6K
j3cDrx0uWoev0fwonhHASVKapmlH1uZBcVxi3iQM7u6so7RZiyxnKYCHuFh0neIS
km7lAKgRQbP9gYURYaMEJDPjXfuhkX9xVo7Ho3ajJCLTLVU75hzmzavGASMOwijA
p/BkMIaTMOzx6W3b+hg21ZSEbLPwsi46/SzW4IO7wKYECtKchItyVMeYHSNtYGZ4
sC1FTDGO2mc39PEYvMdTzrcuSuXqgAB0MgoNfUy1Y56tbxpUFts7yBbqNlw0ZKZV
QHY92Ma+8vLvixpLcgkVHcSjFQMYj8Ac8x4eEsv4HkYsAS9ubdaZ7JAqDeweHFSK
onpUOt+Vf//XQ8ORU4HnlIOsrCk5witzkF/5hZovb90yxbAErIC3DSKmmwhukVDm
SaZDilAkCdFVJGpuum3py7+EhvmUSAZe8K1AK+tDsFD633eR61SdEQE8XGfo7qlS
kqpFTL2bSPX4D5wpfxYeTy0NUSWfLkAVYs/6KS2QCyzovEKph3JVQJJburZmXrJs
Z3VUkFTzj7MVL9htzO5LhvvZoAYiaqMFxGcOY2/e6J9MNsxhTyXnzAltuLrOAWew
6GTEuNO02xO/WeZet3aI2K4ggyXKCb3+UbynJa1SKhbNqjb5JBPPggNo0CIwqRvg
VJBx3I6qZQ0WNTjpHQNZ0GI0um+WaeaL5fooLvoDq553Hr6fClUCk6GXLbQlUhZm
GJaAhsUYl+/4083BTVT61MFUj/WIeTeXfxgdLI+Rq1u+JV9VhUE1TeKpr5Z99u6P
GUXrvsxdV3T2znBs3r58/urNyMy/vZa7PofvN6PmuQjZbDtdC2PYfgO6P2RODLgP
6KNYK6gcQTxKkzG4obqbrWKb/Ioxh064r+P6xKL+JuAqTXFVxsk2ewfXVuakwVno
m9CpdnJ9RI27pP6NIfiwTUv8bmT4aSeQBSbQa2kZyosLYO8gUw+spBV7l9F9NXse
EuwrXQAUJfYuAiJjFLAxtktcJS9wDejiDyXf+8JZ8mcQFS4uSFlnWIJkZ7dP3jz0
BZ7oMXG/zbFwAwCTAeTdMcC+l9d2+0r7Z0SB1fp3Yzrp3Q3kWeccVVrWtwbBuivO
Hm0IOvqlFm2xUk8XGnuJTQTcoppUaP2/0Q36jRPR8cWcX7q7Rq8a08pP1+zdRNPm
Wda7hmNeV5H1XqeTY1414WrMWFh9mBcBaOPK6od0t3lrPTgcCgRCEes+/5YDlnHx
5/CSxZRRKwlFdvF75YltYinLiWJBkpru1kYiLaCbKDZn/A/0/otfJYfTC8zTGDet
YlkCd3lTmlkCpZkAZ5HD7kJYm5GYVnbgDLMoq55SNsp0g+r1bpQAQq2xr7sC4hxT
Y7kMTBe6KJn7xjGuYnPBlRfyWbBAuUZzpqWRdd0QqANmIN1we8dCiwGEJWi/1OhU
QCrMgvDn2b2IJuy9JJupeoYDOOzS1tvmawBE6ASfvFCMUTl9hqfvFJkDyXp0YAuQ
dV2GNJs9fNttCYi0bgoJZaSHWCd6J3LJDwsM/ivodMTHG1/ghGlu3TSBf6E34HFQ
bO0hcW9UXq9pAOfRcJOVHeAk9tXsuK4TK3bZZtOd2JIzqderUDWNWoorp0tPJ5eJ
0H828JF5bWAXKxMCsXQS91D7YOSbWFkG7NDK3HSs6GxgPRfkJ34bzbHytl4KuI8d
9+YlmOcFIJbsND9ju5dvpIQ6SnSwH+tIp5YcpMMiTogd7Oo0nATFMejeQbVexH5S
CEqh9H6XOdROoJOP6BXAeKhxJu7wwO6DKIrJX2b/R/Vk51ZTq9FO3LAr5u8T0oV5
4uzAp7yGZAkfPEbvrEnCjgOCjYCLlhGOmw7gg0e5OPXWzRh5K42TBcih76Wd2QNg
UBXsgFP1UhAm9Etq8X4NfQKSRp0WBMWTcznrJcLYN3kErDt8wN2ay/9eW1FKuHYY
YwYwO+acATFCiVoE2wjZGU1ATooS62mtHneai3KURKHtxSln4wsQ3WJQNZ6NhU2H
esidDGF+topUaLitCJwH9DegtNgF6N4+O0dNdcIiQGTWCeucdYGYnKCyAs2Rg2Ii
jwzXola2qdT15IIayOZpYg0FfTiH+Jr6HSZ2xKaKki1a81ZIB1Imq+RXRiLYpyIR
KFqbsibB7KWj1oD4vgpAeTK9WKqObL+4NljBT6f4hjLwH6JyUe2aMVZLYLnXfIO8
EV+/f2850h9eYXIpLHAe/7CUedEEucjLCeJNvxmqnUK6ccs+K7dCxl6r48w7C/68
A86OgvCSxVupCI+d9i4EalKIvYAJDF+uYoVrisbI/mYDRmRzywVY7Mxr4t+Pr1UT
zb6jraV3lrzKXFEfMJPROdbZ85YKZV3wn3AL6q6V7r9L/pd8cxNwQPgEYzi8GUdx
8UbQMTFY90PFYPlHsIXmAeMrJYX2Hb5zGR6Mjwnnoz4a8dPIu6jbbWBOpipog81S
Y+hqeeWNBh+2APXhpPEDRFBey03BaVnKJh5TVExoWMNKAkqnk1cRyCOnYz5xULB3
EbDGj6SGPzCIV/S8SNCr0OIPLpn7aFeiIlmYKME/sIs+n+U4zXuJRwRKUhwlw/Al
ILmqpF6iZU7Sfj/+o8SttutWZic/KKx133bqRQ7MhKTjUSFEhH5wKIgMyBW8OFC2
ufzEls5a+Wew23g3TbuDq9pORp8gDWFQaIRcJPyRixlMPz0HQ+mYUzvaxS/wz0c1
izS60WfhDk0vNv2C0ffqBe6NcnJkIDVYWP1Flo07EAz77S8cZIq2sIhs4KcAdLIA
pm12rIgRx0QXWt4jXgtokH2lJdEVZ2pTXlVg5SaDiDCvG6B8EgZY91sqxfxhzeVT
p1QYeVTsCp/MrbromlmEYRGT7KuR1Bzz9ULyrQyUoC9SQ9Qo8UZBM2/vE+GAO8VD
xhz+0knoCaCEIjXpNz+sHHIRXs33v2eN9Y71qwEeko8qOLVyAMs7q2Vyz/3uABFR
J1qnmq7lnAgaBDHkRrTc+acLkgi494ISNVR7RAz7SQX/24rd24E4zxTC2lKMQt4s
k9M12VD8wh00UtyPKS2WJRS+nNPvWAg2/YdhsMaoYteAna93NFM80ESibNWveUsw
QmymjqwOMejCipK3BHA80RnwV6sb1vUW9rsCmqJzU8YIoQ8CBns31nxqfYXEMklx
pKYiZTwAARxaZX/aZDKW31RTwC16qkHOpeEppVKAtp29NCTlckz0t1H3D8uUhiFI
VWx3c4j94cwHAHS4McnEASQpf1v41XLa7FSUJOl7mqv+2i24GVMNI5DzKSZpL6oq
dPZI9Smav+f69yvNSaGWMl75zh5bYp7D8JpWWPz03M4NnvMS9BCBNNWAkll3T6Xb
kboj23ZHmpGJgzAXq5+QJWkXVQqN+vGp9SYXGBfQwNu8XNCO0SkRWg++/xeI1vCk
39voSLz14DMPrWtAbiAJwbebsYE0FoiFWiD8MoLvpb0mKKSxuIlMW3ZW920f1fEC
2GXI2fjZiaksAlmP6QI3+Q4s09N/LtdMZvAfz9oK8yt/xtMCFIR83ggu2D42g/RM
gqggBo+PnKjPpd8BEOwvEVSuFzc1j4lnRT9cyvkbEhVF4hGZJCWc2FAvTK70J2oT
GFQyHJGG6K1Efm7RcAH1YDFYpaPp4335IvZJBH1V3qTzx5Q43drXD6ch5Aw0PRqj
7TgXttlAQWKw7bvrKDpkVsYpxlC9xR+Jryzq8zffbmf0a1g7H8CRUj+fObuOyHvI
nrsY0N89UTPiafFonJo5kfsVYXREejGHWLMV/2Xy4zbawptPcVPpYFz+T0InMLTA
Z2IgwKoD/H7gFCPS8QA6dXjy4YXlppKcsTDNFnCWOf29edskw+Wb1keDnDhWZ9oR
RgciFbJFc+s4JUi+hQsAPm/uQQ/sC2dMD7BsAARrDYJTFpvi8nHdHnjGt10214V+
Vv2cyELlRS0OYQnMAOvQds4+SLhb73OK1SAKTiUWtonbWumtiIQTUef5n4vXNqou
4O4pnBqQ1HNqZCuf/SQtlTuN0IXSRDQfxsVKHw7DhW9/oznfw+4R1FSrJZ8tex6K
xRrGGqYdYRN0MJ9Dw0GSa9pO7R9d6ZpTmbf/Ka/MYKlGBBwwvtPF3liNzb9eyRvr
lFp2qg1siaTTGwQzTKE+Smjfgs0cbJFaGiEsGwgr/MIw2ABUyoZj7q5nDELE1lgu
zYzq6fcsgGEEy+8C24pNpWqLU4RImH44c49OqxNbNGnSAW0REtz0gcPmq6eu+fMe
L4NwhQHekSFyDA0yIl2cc8pJlpbZDTMy7pn/3Iz/0VvLmrVXwxIlaBJd3k2RtiUm
zeYRszuiUnfwlzpu+V/8k320NzdHOoOqMwwywc/9ykxfiJm9eCbpaxlLD/HGGKty
M0T4d7UJhbTjm6e7RL/9BDaHqo8ouv3qSWy1Wfmn5sPQXHdCd7i/cauufrQIM2iI
3cexUleNH+y7pJR/WMg5DywkSLmUPgiJufK4s6R7TBiabpjNc6h1oeTj/NK7G6k8
VJrgoj8ALzC9YkOFM3NsR6NGTjZYQGNA8QFHzCtKd8rP1I7z1GXp912LxdrpPfl2
togkbdOo67XW2FRyJu/ntiE8gyVS2wLFN18m/HL7EsRUMuoU2JlZPFL9AI7fLl/s
sX8HVM7m+CzIdjgz8eqRkKY7PRlKPi5OTr4GZwscCpxSlUZu4o9aHoI8KISuoNgs
L4j84gYyQiBh8XttNsG3k7qjtKCGQIjrptTUvQhs3fUehXeQHoNSBM1f2XMDnhUS
u7VckzGZBrRJF/kW1VF36P65dbaYFJcFfDoMpRbagcZs+kxPFCNaa8+cHdao5XIc
VBtNsh4RUAkIB6Eeo5YM3UqwfgC0bkyp2vIeQ2En79ys8XjKwB87EDnQiDsXxvPu
sxJ8Wri8yYoR0qwfTjsUl4k540HetXTqwFe7RPnBM1iu2PiTg/YOooFWJCbtFLJO
iiWEoH1xYSMJ/NSF1BIe7begPqGMSRHrddyHRq4yWXKuXO+UPXJzrU/O/XPFA5Kh
xVJBY8HK8lJLsidI8ToF3BZqeVNiNY2wrsENJUswYrWxH9vNufmw1xlhrYerMNut
g1W6R06cP1sl0ncDwF7qZkumdJ374D0VTIn6Dw1dSILFOD+z/CdcF4A3NWtHLuAY
qYqFpy1J8j76HM0eH3ZpRPWFNfmIf1T0KuzzOFXXUUReifqK7/l7vcTMyfurbUMh
LBIDpH+06iG+xe1G74chnxqJMpQNVdHMnzpU3MNKrCMu573sMjXQkZMcGbLNJ1Rz
4xmZ93E1Rl1JsqQSroXXUPiuYJcjUAr3BEAqN6aHyeWdVDoGldbZvIBRn8apbEP5
DkRsbN2lXZx8ojQB/Q9+WMy1mjpn4kmfghmuEF9GqzsB0Bd91ugws47lCkf29+Ed
rWIKzVXpqWvT9h9zmkLU3DqvySzzYpYXKwnk+vTYDpcRNSNo8k7XU/d+4Zc1kABS
Lq33FaxrcFRi+ko7mdgBBaFEeP1KGXmxpbNnBo7tQwo0B+MeOTepUNSZ/Z91Wpi5
q6VZv/2A1dpfLh8XFXzDwX+nbT+yo7U0guRIBA2K6UFOEMu1XejlQdkUIbsDrZ5R
oFnQZau5j22N37cS3PntRWHbVmXqBKukkfP5KlDsg9PBzTztF64a9qWtASOvhOof
vcDC75FW/FxaoeXWwBxV/j+nuBJYRKcA7/q26BkaP8RdzoF9Rvoqnl+jPmiWqxth
0DMcjB5QksJDjFeaFg38dKxU5ztst60hUGcOSO1LHjI2+Wwg4fUWynuTvbrcdCF+
qj4gjmThtk/XaLvyECPL1B0cZO3hVvfmEIIDwboyZhonNN+rITBQ4gyfb+SQsKbu
8aL6Chfr+3suBl/SFMUcI7M7U3Ls/KOSgQ9hizbOYtQw/fvIAFtMwnwsqT1mnWSl
gDua8Fa7LvqGH+3eYtIBjl5BbrWHEPg3pBaw77GK2MXwGrSxztuR14BoKjlO7TMA
Zb3Bx/iAeERcFbOuHS49EF3pCgWGHSTokVdsYLwZfU1kelShHZ8mvmOfucm0yynu
/3dPWODfwZnNd1iGWsd7vedhA6MSUxbj9LBlOfRxQV7OkByXmP2COQnD+uWiiTTd
Gii5qc8hfgSNzNeT6U0iRWntT4AUH22cvT+t6+MjIgG87tOJllSKePuedlioXMhZ
e+gU7gJqWVoRQa0H521LyjM6oizOfriX78HaimkpDjsNTM1uzK09SVu9Yk/1IGQd
HZOS9DvTOG/TjKSDbvanGpJrWCCHGwESgrTo+lU+YbbBN0k+/zQM/aRZ73Uqv5U2
aipSClOrAFGz0eEvQX9Yz5DAp1pQORCrcxKkLZD1if3MY5U32UORGE3W41OJ0K56
9mVdNaJsUPC7oM7irJzfh7W40wpZfqmpTLxEksGxhbNKinVM65XBFr1+nfBW58uH
8WnGfdS4gl3x6yYWgBGe2vgUEoKH7sn+bc8yAmCZtZPMvOrtZiqHRbC0VLeCL9D/
AeiYbMwUC+Xr2GfSnJm3VbdBxlC1YrvLRH02JHEMpaObHEfTvDrz2/Ad0SajVmxA
E99oBnE90ce1BkTbqsFYoktwDGljlX3XVDTBnj+oWGDVZjzctaU+N/FHU4es0Pel
d2Yp+8FGlq82P/0zklEPJy9670w8tu0vknMJMj80n/lpFlh3Jw13v7ILzfdQgmqt
QQyU63zcp0V+FOjaJ7dSl5gScF5kgc6LmNcKGS4pFOtTrWfwJ1kET+6CWSwUEtkA
dSdrI7n4x+Kb5ntHz3OE7wgcPmWMqIaTGVvXFWDMSzQKyvgEjY1pFMcczg7dyxao
Q4vr7EYman77szDNZYZjmCuzhRnoj0CMD/WtPuZaomBF5/imDXeBqSjemCSy+7VM
QFNpy0LYZhIOfAbm1k82GNHfjWow2HXIhtRj23GRgofl71vTkEIEgE4krhilIJhW
P+YcG6wZ5SeTV/tD5zsQM1Iv+k3IvW1dXHmbzjwBmiSa+UvFxUbc5m52uEG2ZVlS
1/o9BkAse9YDkBqDl6GH/aqDiI5yuMBCId/WHgo+rtQF729fHOopzS/qgxNJSDLl
ksL15fghQfVJHbGfRVk0KfRNz8JfVMHHL+HnUIqoUHIgAwYfpZ7WgeBHtB77tsKL
yF5ijSvaXXKOY7iyXk0cSh2AqjUvN5XyfgQSSj1qYgcnFpbWfp3AuIyLwvKvzsfh
VtCgTZS5oqCB8R4KKDBPW/9vP8ZBqYy0cI/uN50/NuaC/ILkJf1+AdLeFkwYRfBe
HU0ty+EE5bLgMXHBY1Ku221bHE10HxN8jjDlXcLZtHWGwTW1S82bT9EGcGd2OjmN
VCIFmynUZr3YVi+IoBNgnQG2HnQgeog2aVVIuUPkx/bed28zl8WFg1KjO3Z++uDF
Ugf+y6gyMNCzR76GPJmNJo+eCmR6dZLhSNozuA6TRBWXR8eA6Swns1RaUZi8gpNR
9e+g+wnF4HFEyNckaNt4RjJZe0Yac+mcQlvCdLG0UnAyMSfSpP5xdPbsXhzGc5tZ
mHfxYr0C2BpTEY8fHJhb4YT4XZCc/ZprLh931MbW+hPjc+ku0kIwq3F8Ckhla+3p
b2/cQCdGmzZM3IE8xZB/jiZF83V5ezSt59frHXrP79cvJVIC40n1C572g18yXEZV
1T1OS03iShO0wxzvQKnGZBsFFqCaEn1SuWFTY7VvrNoap9736PFKBWIlzgFYk3dx
p3AlHBPGVvvCgF9BHJaNS3mhUBSeBSM8IxVbVBmZWzfq/tBLvTEn67WXzxfN0fLY
oZpP03YUk7glCREAupK48UnJlfNfGbf0D0wzVXoB2pVW2eEyAYBpDEYM43ukf2M0
IK5R1IHTzJGwGbB9XLBTvpkRq5yw3b8BRYYGh8Xuf9p1m7IGWIBdg0pCgWHuq4U5
CStsKbIwKofmZa3jE8tO98G5vHpVcExK7j2bdeSgIBHuzl06NCmeveIA8gr2S+sA
tniMitXEy/KlmKIyrkO13GJfh53hfWgIQpQkHQP/WC8v/POeNzsc4mmv2SNpICRK
BQudrMXT6OAwAQc/peJ6+e+aVeNpIVqRzG0/bu9HaTeDMuWI/eUHsNM3Y5/DZfuK
0sEcAkwFJSPMMgAda3QILKOYUag2FJZGHET90qOrCgs6RWTJnDkisvGG+/8b4ZKX
6Lm9nzDqkmNp78YtUJmMrbcjaA/cl8/SD/qmP/Jdzls5MrzJpGTKkAbNo6UOb3AP
LNbPmrv3QxNFQS0I+AvBQyRZgpxYdoqOQpYCS5kv5ZWpZKpKtrfZe+ekju70g3HI
N+zZlVqS9t838aOSBv4Ler7vDnehZTZLjSjqzUYkaBIzb6pJDYUCyb489kF0irDO
6D4oVt0UZP8xv3YfiRJMnHYotnGmnh5Nx6p4hOf7uilKE39mTL+L/7GZdkRInEmm
DPEa7uEQebJc3xGV0N9MLwI4UX7hFvW1SgTcpKYjZQEEDxIfWy7pCa5EkjQgSMno
iLTGsHuqzyQpScRZtQ8H8JHDt3p2YdToBofzjtpbvQKS+kHkt9YzXqCOkAPbWOLQ
nm3L8HEtKXcUXbYXTx9x+Zzc7dBSpCKoRTX/BJ5u6JJC2HXzVU6GtlEu3wOorj3H
HuOCRN8BwvllZPe5jyOeFdTpdiNWmEHbPP9+9h0x4tVAjdxA0i9X381XkMpcuRVM
7ADoS0nDDeVfgyTbY32iFXahAt5VI096NeljceI+JVrIaTcPo9yjFHiIdQUUSQm5
MtjgwHYxwobsVmbLCFV8ATeCp7QeLAgfA1DCzuxdkr54/kID8anTG8t10luVK//B
NL1ZuKV+M1096oZgQrx0UnU+AlBKsIWJVDqd0GFipeCHSGHTqFVjBhUshTDCcyly
Gg4oyLu/E0PIf1PjWVpcDHdTF1kiiy+waqqcz3Xo6PZA+C/jxrGG2nFnfko0NdOr
/6VjzLFslM56jY4hHBtB7aSkzxJIsYTfX865Cdaoyuy7kmDHFx7zR3YS1U8snjGH
Ba/I6Q/rNzbtlsaJQtJl3mf8elATtNDptp/GQufV8jt93GmvJKMW56A6VituJ4yn
gp19xlPygnNdJJcJL96eJ5rqce7cAYv6+Q3FKXn2ivcUh6RIe00JtSRM00dCFYzw
wPzibIuNXE7xA3/cPWMQpX0+cG5Kj2jIul9/S/SCdtHOIZ892ohXPbHWMOgnQ+sp
k47pA0jWah2DUoVMYjTlMFk8ETv7Yf7nVJNQ7dj8gxColjsQOC6axxkcNWvndQ2v
WhPu88pOruv9V5WfkPAYWOaZT8YWMxfm8fLP97Nw8SEg1GdzqdC8oSLlU/MOg6w2
UNhP8980+4FeU4FYX2CFqfdmiDAyP6HcxPgWiaKhPcrsGk8dLfesUOei2Nji3hYo
l2Ugm4k6+Z+wxq+nFIhqD+37x5LXpBKM6tkRD3gH0mQWkVhNR/3j+wj7ZOvA5tTn
GuCYulnNTXBXcK+cCda7HKKIqdRLY9MjfwWxPetKKXKU/t1CO/vhZ/nP0cSyM/dW
cFtFoyR6LWR5oRD1N80ngo1RzzFtNfSkG22hSpMW7wY6CqvUhBFwhs+hHjyuMQ1e
LfmLnMHTcpfUlO2IROaCND5Jus/dX6lSh0Ds8ukUiLJ8vpoAKlxjmf99IMHadfGR
E8qLiYVNwCdScFZGPp+J7Z9WnbKerZnfVrHP9l2DIJl9m6wvDzBQ2z5U6J/pQPgf
Sfj2YVruRRyRNY3kLabo3Ou8xeZbsOSk5BIE5HxwC22Nn2GisnPVo7/Wnb/73Kzv
m1Otp9b8QJyJ64opcSWeG/aAGpaRM5Odxh3wqcZtoZkNVNQVrPX1wXU8jC9hZlb9
3FU/ar6wLxKrKNeZg1oA0/i5bBE0PxsSH7tGmJ6nZiKEtUPK+ObP3/0Xvp5VMCyI
1WHKd/6UgFD0QxaXuD4/Dtj3RMNJK0EIOLe8pgucW9rPJpP/y15xcfRz7DM3RZff
ebaOS7FmOkwkQN9S9QnhXYHy3P31SDgiJDA4SzzOSLl30lW2SxweqmCmT+PC5Npe
9v3X5SmRwEWc9TtDGZ1VljcRNSvlJHmyUjLX0Vp95b7Umen/Wv+lKTTqvaFsgRSG
Abv6cuDhoS+rtzFcs5EnKz8iGfszvjUcHYVCZS0r0473OWOMEl1ofgFdi94XSGRa
1R6fUK9l3x7wqxLrznl8lxcMVyWfHMJ2IzF3Bx0syy+q5XURHAzEaEiqgnJ9J35q
9yT/M9LiF/8DJeStrFCeDjiR9G8CJSv7b9b2fEPeGSgKuceKiy2u1nIl+opCbYKm
mYL4OnuEMLZUHjvRQvqe8cYHHt9ZT1sZhTD6u7u7OTBks5N0TAfxX869Jd3IfztV
yLhI143Sh0JOMfrGnXVMkAO79PirMm+tSeWKUPuqtYKaBXdacOJOfyVlCpRXRa+E
QGBcrXcb/N9v0t630nu9vJmRRODfuKqdwE0U3Oq5XJ0SzYpOlq/74JXkg/1omou6
WbYOLPDiRfqtCFTGacDTHiYO8bQxXcnaSno8IXicUTkEbYfnCznJWQJO6yOO7yhR
lIg/kWX4U4UydgMSjNaxzWGjcE9A3beC0RpXQIuPwyxJE2fnA7oy0VWPGklvoPGJ
sLlh0dJdvA7kC5GvqIggkZqnIUvlhXwJ62OuC8Hg13vnfL1KiOZh7qb0jOMEhfNO
Bf5ujFBE+/LWl5551fQwBBOZj6InZ8Mkq4FDi7jEdfZRU4Ajf6Qh05ZWFX1mUhZS
PfonuQz9+/ZXiyyqudxTMvpEza+T3yIhdFbRzKPXXe224F3UQ2aH6gR0+nSvQhOy
MN69FYqwNw4CYSs1WzrXBKkH8nV1Ssc2DPZTMksXBPTeSSSuUHOS8DHnpNajmlKY
wEza4tfj6e8Kwqr9H1MxR7Tcso8HNUMMJYWdJhv4LkOqOVfKyiEiDBeJitZeEO/n
hkfydcVmk8iMX8lEwKxnHYblyFYVyFTpaYq3C8Pdu7bkwsNbXpT6idxO8M0y7eE7
M2PSj717A98UkbaS0DOoR64ehViP3Cb30tEUSEzk5iDtKMX3HUwf//zcyRKqt1Qn
ezAZROSyWhTOakKqKr+GOYmGfBHM6qR7AWEsHymePpO/4gnW6zx95eMUgQ25QuLj
8PaXwF34Pa5JWVa8g9LR5s9MCbhpQP9qn0AA/6+4ILqRQJn5WY4rIOoZzUXFioaf
HWhXEf8tsEQNdIAzy7B8DSy3yowup6mzgrQk4iRmw0ZwzAjkD9Lq50kPGxknzgWf
EyEGhuALf4ttOa40/so4T2l2XgFgMkZWK2Ggkbpygz3cNM0M+NlLcs8cPOz5Facj
Gqsb6ozL8lSvcFTRpPYdVF+Q19+JDRmroMz3M5Bh3KnEILFWTu/yz/nVF00zW990
NKmDzjWGnp46yEqYaj7yc5abrASgG5/gQXuHPxzU6KI2sDbxKjCwlwgQT6aad10g
pyhF3zD7k4azzOu+1JQqJXz7bScmDr54bxj7jR5AJhYH7DFRoVdLXnt3/wUAyCO0
wWaigYi4J4b6Sh9bxaAYC7xRD3oq2S6BiQi9FOdpKDgeeAS9O0WJisV1yJ0QY9B2
j42evliptfA+qmPIOM864I428wQBVDl8AnzUcC7wLTu12ydOckoGfTj2sSC7tgCu
JbFU30EZkQFR4h2DkRtyj9lKJ7UeE/5nWd9609oHes/Ym9X+j36WZxASHpj8SYRI
fTmWKzX8terXB1gRDecPntN4gphtdSjIv4wNUW9ZnTZ+ZI6vGx8/+KVONArpqQW4
IrmR3OkpaEpiC33KgY9nNXXOjWNfR6ee4nxicBxvlBBACey/idIEuor5VZjzIgj9
DMz1ogmDdPMNsn5PpjUeqsP60u6YNIpKHdTTutfkwtuYk/RbQ0hijcspn81nY2VO
GSKsOj6rUr3Ai0Wc5RW3u6LZ0g9fs34fB63ZnoU5VDUvGj1GrI+m/PocXlb+anDQ
urC1GaX+EixIvpxbIcWb6MC/l0A9lqksXDuuQNraZALk91qMHfl3UVaU/LwenBcN
nWCe0k4e/pvTHgLTG/TQdr3DT8udHIZk1rAIu7ErYP6or6bslxTp4l22fyuSRkiv
lVo+Jo8+fjRvG9nCXeib7M+SaeFTZV/vau3HawWPpgpgFl31wRmjG+pArzLl0Ysa
m5ChgTOP3KVYniJf1m2xRLA/oy7Cs3wCQhYI3rbd2hRhb7nRfvdM5g7aAhz/oE9Y
vY9VFlDHvL7JUPtOqfTO0nze2L9k+yMfRh3H7aCTk83EF63MPW3s+ItVnxq4oKB8
qJZ6XfBkFXqu9R5EFTQpIJ4UTFnfVcKL/l4vQVq3TyrOgCIPPne6f8wObGN7rDy0
bmbx8UobYFEHXFodJ2STkUPLOepa2Dlx//ec60r1Dk3OoubwmhAAFO340BiGpkTD
7+mkV+cbJ+1up5688ZJPdGPgWdCRCVUwjfXsjL7pzQbnmL+n/mQGdNaCBH/38lLy
pttst50CSDiekRDaBuO7k16U+5zc5yNW3B2a+8qy+zyQqbl5yTpTgZivRiGsnbTO
VQS5a21rCYw1N0yR2AFMWnb1Z1OTTjuwr3TuJGBPqfcZHPdN7C2AmakL4hk+gbmx
djn28eNO03cZlShOKN18oxJ+vYc1Wz0bo9p/vMPi5vXtUbMagLoAKmNo7XWKMgDV
MAGbQ467qBvwAMF20F+jZRS04nXfkcCbdlikz1hCvSO3o2z8FMt91Q+o1lNahkfC
GVK1/iwF8MFOq+Ke8g5SmWIlx97iMzxdbDAvLeIIewnMu8eCUiQvh5nSN2rAvlaR
XTCdrHpRZYqlUGrmVLnP8iV9h4lCSDQfLRKgVcA5f3Ba4IEWR+m7mztsS1eTfpcp
spjR5mQhx3VouodpstUh/AKPr9jli94JawMjclhfdC6yBwj7R6e+49RkGwY9lgU4
PseNXm+5+RU9gE/DQNdxB/awyyK1GdVDaGuEH+U3CPnCSM4zEW9MrR77BDr1Zfbt
S8b18UBHmUfXLBrhtFLiTRxkd+xucsBnwHAqHL3BFI8DL9hOn4m2B0XV3RJw0N6n
5QURjQOllBWPox9OqLzCQQoSO8V9RCwmSkgWOdnfSMWnq+jgR5GC/18hVD2SLcMW
Iqg4ObmggHEru2FUzXWOZhNWJEalXxRUqYsV52MYuFRIvEuM8J3jMeMj3i7pwl+u
WFfNWjcvOUJ8Jc4NLbQ2+qAOJF93pwPUB5d3Tm1vBEFirdgKuexuyTZs02OIAIdP
O58LN9VZVQ88761j2qnr7CxvPm6GS7ILNbwL729VKQ43t+Bo4B3X79XuSRIRYk0B
qCMk26dvH1kTfvZEFNkgXun7RjWTQgkoweQN96h5IbASJf2Y3vxjn84av3o4D45C
srHlwhtG6vN08uV6hLttYCOCdSSU8Yi+JeSyo2wivcdHj5psdoVWQuyLzaVPNbA+
7pQIWz39CTI/yFE3tNHfsX0cvGCN2PJOiYQJOTNCxOgzjl7cp+y1BB7zC3S7+28d
a+x5o3rcgPiiqFM/dzWuj9Qm/1bkRnMPswGPY3iVIxB14cbzHSWfVEXfAIMOa54m
lSbeL+rMGobWC1WgunGwHPoHMilTCs7GxYywqVqZDIZhUIsJJMco+OqZsGkLnix8
pbdwTQB6mvH4WWY/6/jg6QZXVguiEQrMYMq6ETWaMYKnErJjksxc2idJPKumwJs2
VXXu6qU1jZNhZU+jmiS3SmAhABe5ss26fMpb2OG+bbewpengJ/6e5SPRAMwZWi6n
5AXFRfJMir0nmfhxzyYLb3PU+7q8zVvsJEfErRFaSHqHUw3M71z0gdLX0lWTal5/
eQWb9ZouJbK3c53VqxvwKT6FVeYldRe3J0ZerzMsAbuLlNeT7YI7s3l/IvuKcbx7
EBhwDJlu5yprOpsgVC2wweogJVyUf82M+nAJt6cQRML0j1jjIHtWB4ZbT+j55/VB
gK+YJbWoEv7mmZZ6MSxb1+GBXmwVPI2MroU9c0zuAELNh448L6X/2DpmqLwnHoW2
HQku5hFR6jD7XxLe3gZ5HNFgCIacVphEapKjzVaYQQwvCTGMqbIVZkrmCfKtFzEi
34scQVvRlZ5UUWKwD5HtAhsYcEhxMQioH/ktcOo+HvmBarpyM65yA1k5+STSKl6M
FlG0Y27eD0CC9Z4PUlzYfk7M5sVifpSkerKcwOh3KUOeEoxklecRNbJ+9aKxoMxy
+OhVj4bRfeqZxb5uNw54jdBeALsb/9uZ9xTzvlDRJmDu3vhazATulIkfTXgZWH4q
qsdchoT/ZX2YuGJNPTCPTawShB307Wa7hTNp8Fhd2M3Nda+y38NL4QlD/n4IH9L/
7tdwJcsdTDSn3TOzJAFCjFi/MNuIjaLSyNQXXScHFiIHGctAJGHcjQgoT/fMZpxQ
DxISbgtNzLwrVkdkAmvJ1tkLsGSGr3OTQBDbNbF4apA0fk/uyn3JERt4ZZPJZVHI
E4r/W6FkIQOg7J3vMA4OkyqTh90X0sBha28U/hfj5VE5SQgy8w/xE3xyMBXe8yrF
L+9dLGOWzFouCDoDSHlhVhjosujVKMbXmts1VLWstF3+6Tzvza3b1EKLGY3gBhZA
Cr9u0y4NE0YEBTRrOuHJU6TsFdA9tSdiZu9SzE9Fn0nPnNw1of9QHWDiag1PFWfS
BDKWzJXKQJsG7kR9MdSBxqKS2cT6477E8+mwqMGviS9j32HdE7wyI/DQALv36nde
riuI56BKsqNY9Qgkpc7rsOdXdU83CClSBwMBRp4G9S4GWsk9P983r8FwwY2udC0t
bZRN50dmCQeV5ifIX9kElKHemTQqgUtVzMsBPdMMY1M49urMInc2K9saBKTdk+bY
C6/Ej/EAbFWk8DCH63350xyK6qI4psThW+fuNy1oEWoNGp9TpGH5QcpiQlniBfcZ
Qi3N2JCddpeaPAXZCEK8ANtq0efWQd1aP29NEAVqxxubqtJxfWRbG9onYBTGRXT3
Kp2ZfGt/xE48GmxopszUsA3FxWeY9VkDCnDMyD+S2BEpQ9SIMSyp1pap/m3Pxchv
euPycBjuHS/sV/0gIHL/ur3g5zUR9kxJVPYDeXoLULEYZlPFgGYozijjvrXgYzbp
OrTajBD/g/X6CUOfwvU6dK6B4io5eNByEWPVkr+OBmUMx5VpGzcjxV4WkPMEA2qk
2wYqeYaTGKQJUuuyin0X14UHqVGTOJh8Fp766qwPyPbMzz3Bhv9deKrEw22Wd+2K
Y7UPSSfxazn3cKL2WnUlVCPw5MSyxPG+/NUgv7ZGeTQjkgufWpjAL6sjo6wu1bgi
tW18x1jAaLLy1ymwN7mvMU1YNlQE5X3Ctlvm66Tb3Qx+l+6kRJW2fu6qtz6M5N6H
VyqFdqeBV1UHjPtqdcdxos9vNues+HYr/aAXjP8EJRgf35EYbbhChhiMzfzKn1Kx
4IbjXmjQSoBh0+wAgedc62IUgJdqHUqDmp3RYRevNfWCxM4dT1xeTLrpAV7D7PL3
CkFP7AHHL7Vh095FuGhnx6TLAVyfyEzJD5bxy7y5dX/mn+A7nRJHlgf72Lsu5UWb
IBZRzn39zjTv9CIVnqJLO0Ej9IS54eGDYyGHFfTn3Seb8oMV7yIuIyewe2VhfuJR
x4MsW+DoiUZOJ9GDKs+EjhXns3o20EJpUnItPeDt1RORCb9/tvC5dfW/2zDDkYF4
q6GdYYJPHGDtT1KMoRj3OfSYTpLEE05d9a/eotxJ7LegHW26TdSt9tGsJpxsLk85
fpeYzXBvlIeVvaDDwfRL7HIytdXSI5OzmFNHT3VTivojnyG2P/I0uCEbycxdzonq
qxzEICGxs/aD5ZEJbA8W8JF5cDZK7m7wtMy/RtgaDRu9jP4jNTbpoG54P57twgnO
EvU/smQFgokzZBnQUtdtA0KT94sjc5neEjw3uK8NgS5H4wNMiACGT9EoLlxWcqoJ
1/4VDaxFmpNhDJe3DbyF/aU86rWcJkL+5ORVhwKOftU4jP75mZTu8Oa6fWoPLN0p
phQ/GDMPPYyhd/rdTos1vFP8+N+EKpvNkPjBfRyaBFNafKxA65U6E/odLt9QffYj
Di1y3yS3dAEMHoLEyhDlEJkCFl6eBDfs/UD3gh/LeR3xEp/ONH7y1e1LIMwMCxX/
W7AzG6AtfgRHAUCgtxKdIsLLiHp8u60hF6C83vgCKSxKuR35bLuD0+Wap8GgV7o6
JH7GKvHJOuGJmnUuGRY3v+LzQSwRuqPSqqxpsZuSNFqh9AXRpCfuJWQRRITM1x2i
O1HhGTGf3pMeMDQOTPlk07ukcc/zYIgxxDAYwjTpNSboK573pS7wQ60WrOJAT2rF
a5B1pIXFEIbNUgu8jX9XMN2M76ZPee68Uz2V1m62ryFJ2coQFWdfoAnagk5z3iCD
PuORSqi6Vethdy5d+0D2yA1tkdsnUi6qIbH0jJlPA+zRWe5moeOZ1Qb4mU7mCfb7
8jffI1zV9YKF+GYotqnf4avgv3ep9Rnkz2KRL1rjR0IgKtipTXZr8kPfE+fJ8Zul
llILAtJOv5T3+eC00XFl/g9uEJvEdJqE9fuA/2EdV2bQt1ziCiVluv0O+QepZy5q
N44UzoxTR6KdXLm1mbHDsThtEnbDCrf04qL7U+F661J+rANnzGmiryboQHoVseeK
5JrfxH446/FuxV2aUOlwPmqOMkaakRq52l4HDvuCvY6ERJ27fHH1WYMDm3ypeIxx
Qq1GwncDw/axGTIoIftMiNIGFZ3Szi8l6pC0mZZVFVIVLmEW788wq0k9dwjP15W3
umzyToexOeX3vm2QDTOEERG9Qlrpb/skgOJwS36lL/kwQPnDyyy8LghMUgizJQ9t
pLZL2MfHU4HtRABOK25+yvYnUZ+cRZgbEIlNumUn96d/1BQ3Vdrr0JxfLZQIpTYq
LtAETXxv9NHjRNI4/zhDkIDSwETluCow1GfkS6O7Q5pgaSkYDkkpHlGi2ryWU4iX
K6yp/i3+VecX/m3XmN7vzGikeTdniFw8nPsmcFjl1MReNMa4cInjd8e8KFA+x4ZY
bPs06mjgwUwZTgc44M0OT/1CSUukFpz5F5gCeGXE6xwe2OazM3ALON1L/Qqyuxac
K1PJH6HkJmzy1HCkSQSFGDEGLytoec3k1oP/ofKB73G83oIBXsaTMwbBOTGT8VDB
AEncLq49eMy+rYFHtaePJm2uw7NBguCC7RDN1Ud08My0aZGyJU2eJfdbonZpEDwp
8EW0OEfPmVSAp65kpMldumc8pZZ+5y/ONuSIjIS2D5AKUO4meUjrdCKVYVB+8UAd
+gEAiIKyy3CpNaKNHbK87PQ3Ge3jzKjBkAQ/ki24MYxnA+ttIx85Y+p0a2FCuFYd
eLi3wY+gE2+aYITk0KHX5lMHbNycs4PJuVbSv6PjMD16rShPWk2hfUlmLNxqwmVe
kd+pgLJesidLHygxUxE9eyQOvL5F8XyQOssCopu03fl9XR4ppNXIyJUBeoI8cnTY
bPYFRsvLZ9oA4TUkERRdVSy5urm+eL4uXFKZhLDkhT2PI+24OxziiWFRyrFeuFbp
TFAbJqCMirMDHSMZSvTtdgTjmpWEz4ATuUydi0u5dFemYih5yguiH6HR+cMC8NfZ
Ma1t0YlKnax7ey6tO2zLoXw2S9vS7YWx7/Cq8zkkj2cHI7NYCSHbRqw+tlj/rg0r
9ZJrksfB4weOWg1Da1/Z2o57lyb3dDEIEYKuItW5oI+ynsFRz/GpF5oz/4mUqNK9
5sNuL65mbXX4+1W4ISmQ2QUmi5hvbyDjWkaX77cBOxMWQqsSQ5wk/ReVZ6HyzFpe
8//TPefpwX9zSUXHgzlI+MTozst27HiLBASP7eyG96Rdv6oe1j4wwZv6MSeVZvle
omVIeAEeWl4PIp+Kb1+D2zYhxou1fkkxxOsb0qaGMJpuNFlHIJ9/5M7XpWDb2X9m
pBU8p/GVSyoKZiukLEN3iuYQIpV1A1jY7NumVvmCpC8Ulq3gTgOlsGCVA5U0QrIK
PF3GNqaMLIWlgfqXK1VXp4SyNUIItzxRM4YT28RKovvPNs64eiUTBOy1rrjlhAiM
IIFN7zqa4Sp/0xkNOk4y0sx3fP0d5IAXFevquqVyilWZPqUgHmP7hNUN59r9KqPU
JuA736MhSC0su+j3ptbM7d5RAP+UFjT09rITSGFkfmBCA49jqsjobMGG5kluZiV/
8AL6douR32Jgy2Zf3OSF18HqspY0MJpW+clVxX6ojqtE2S5CehknKT7yP3ZWt+g9
zB/DUbCAvrZOznDe4cTmVojVAQ8inHU5LrmOE2JawSIR38XhEMBDAxO1m2xm52CO
prfT+dlG76EZAPu240W97eZbKwAV+Y/pM+Z/y3T5IPp6ozvSPqz2gokeszWBqlG6
RPCism1cEz0s4sxWrtM+dq9QBQEH3v3OhEFPb9Juds1nXWZ9865sTF9h+Q9XA0/b
JjO2LoywqudPKVSvTTh9dUcGMqw+TVKy6ijrTttgAXDbChQrx0rCDamQYOykxtkM
ByH6P5I/uIWYQeIInqV4iFK+mxoshu6auOsCACGmYw/GdodEb5i2hcv6m2LmMPtw
UbHIPruJ9jahHciivHP5MBZ1ftea2i6cz14cK3cCWZpRJH5Iyqr95oaTm7x2aQY5
+ovzRItigLZUp2iKSd5XdSMNCASJxAWhhgWZMtPu0GZus7nMQdpilq8/laPc8xym
RFQHQIqpwRQie/ptzgucnpvsOk6HEK0W9P0QfSVMjlSEIB9RbXsYiTMD15u7S0W0
z4miFJhibHqd89anUaWmNkoar2K/ftJdCYqG2EzyPrqhNCmrP7MqEmH/uaTkM2Uc
+ETxbTjftMCFsWlc685mN7yOQUP1eLUpbgRnKzPhv3MJzUfBjPMLb5BwpXXJv65Z
++OAToJLhNSVG6Igno+gpPKp7v+roZhvuL/zB3QsPq3ZkUMszyLXBWts8e7Fl6qO
mziPFTzQOgk6mzQd/KEKaLc82btlfMW2DJp0QJ+kXyJp73O0k84VCIHJ0T2r0Ysz
RVmPQYqK9bpj2cKRw1W6/2z7aKiCd+fz3bXVcy1MHcgHFeb7eKoiDJFLMOo8MaoI
qWqUr1f5XIwsEXx4QJd0Hr227AKfUBxULJf2jXt4z4vXRjNUdDgGXTrrMXky6Xjt
dg3uE6zPyD515kGYD1S9y7U3UJUEk4Ligsk9wmTlug//1ubyiOyLuM5JuKdZpLyz
oEtot8GvBWtUDtAsHZt/RFL+4nI7gvQCjYEL6rYA88EGt0hxqcnGhaSt0l1ZVSFZ
Xipb1FaS7CJj1HjwsvqcqkdWymSJJtSN44Sqstko6sd677hY+o+2WXIVY6fU7kdH
a4QspRDSz3jqyVlbyzx0ivIs2vtOs9pMaub5p0CyydXCbro6XkFe9wOCrmfdzXmD
HzhW2Ovxhur52pqOuqRYaG2/dpuwo9uk+P9pdZEhSvO93gW8G495/nnqaolFXBWn
t+Yem8nahftp8MBoZ8L7suCqKMg58ZYxhkKkM641Gm+lrqUZrLIOFZ1kDmejpC4Z
1d+fgyh/FPTgZ6QF4isdd2OGRWVabqnjAusPEKBdZyesgx69g+ojSnDNDYFyfxGY
0OQQpnah7xDPxtKCaB9OekCsKHii1Fu2J8PwETJTgR+XAr554oFXvz4BX+lU3c38
ZkCXdCdqMrSDLSH346e5cwe7v4OX+n9wuRb0ZHoDQLVXnIFl5QIpJefvY8RU8Z96
0FRhc5yVgbkWhOtRzYAENZJ2GrbFJWOgZ7+iYCqSwOFwDpToEwCSLe8rOK489lHO
bnwhQnbHVG8mw5Awt3LLGtOXy/yIs5dbbERrh4+eZ5hxOtGhkdapDR9uJu7DV59a
YMqh/uxsRpafq2SU+OKe1xpedC4STAFgTpH1sgBwFQUfIP6LaZTPWTWmMcnCsoES
ewsd9zqt7C/miLUkGnwv7HAF08I2wlyhbRztzszDrS1arYXXtGc7H36s7s1HK4TK
aZ0rwSwofaB64j/yIhYY6CWFS2fpEgp8jMpPcsLkwYcujKjcnXkTCJu5o70pMqIq
B06kNK/cwNBIeJ27g4b348bbQ24hX+GrLfMytsl+1csqSJ0l66u9M1qor6VrA/xB
NqwSPqWwNg5GEjFgJk9RD/gfgChPGknhd7r/y7eITOBqlt36RY4rfbz957AdV3PU
Dt7WUqSkS4u2MC1FjLcLdKbAjLGQIPw8P/TuTRzY4bWIhD7HOmAh85f0f6oDhOMo
oLm5NODhznJvWZZYBwm70yrl5a0GLaC+stqXiilyEitJiOdyX2ez5QtnTj5o0xrC
dT3CQQCqAzJy4q7ENzY33oKLnzeLwN8TxM44yOA78ZAEkBBWMB1ekKmRtrhE5rH2
ZNLGayOUlSWxjQsuDaxUeNekTh9tGIaFQhT2Ccao+vAHrqVii5bYrolwZ50apFPZ
0LRWVVFqRUXNzs+4fLyRdJReBPQo3V1xhs5OedxjFY7eLahACVldyBLbsijkKdb/
yIk/cHBy7DsvTFQaWijQvK+p4a2UyljYPpAV/Y2yIc2vpBetVssdYFaeEE94hLRL
AzUIfnpnhWU8pK0DcwIFyXhj2YFM1aWDEquk69cqeHuuBF/ZySsAskssXcr1fdDb
CuLSc82VI/ris2xEqelwfLrYB1pExdM5wDm11BElF12XIcFq/TQWYI2mt/qjV068
/a2JUDtvxPVTDVyRhoHLhjztNQtw/YR3HlwqV6YST6GLvp7gNfzKsemD+LvqWPKz
EL9D5XOCRSx3O76nYRWkcIpqn1ZKJClxHR8TXWpSgLfP9sptwrSjaaLuGXmMQYyP
bAIZRn2Iv4mP3mtzK9G7oX0njx8UykdORk4oyQjKVNHlj3ng4RmCrJsa1ZEpP1kI
KhFp0lncuxWnMYBWFlJh+WvS6uEDpNqNM3OGaAH2BA6JkAfAAUq7yxX/0DT0ohsU
OMvyw47nJ5qE6UVfrhYT2UwczbweW+jmiGH5SGJTcXxVXA5wdNR4FzL0FwAUwhAR
OtxnDEVccNCHqZBcEk6PSZrCuK+PogUAnxMo1mcKbmJzwbCxlvpgSh4f9k+MME09
Lo+T7JBFsJ4QjYAFko9zqb8xR6cuKuu32Qkp/HsPtaex1jLNySNXRczyXTFmlQQE
V5WyRspIwzwydzwN82OU5YsOcO+e0zicfsMkzTv9f63eESUXIGWenJXIZVTMjzaS
1GwE7SSAVP622GKAMNRwlm8L5k5UfOrVKeWyjMuZBKiudQvPt/pJeGjBydNX7jR3
n8wdiP0mKBMW4qMZjl0MUEhDFU4M/fwlZWUY8HRR69bCaiEIWGOTw6cPfxtYp23R
jrSQ7/jTznIoUgeyeFMe6C+ldEb2BuYlsSf3zL68R8cbbUtFmV5bu63ORpJ6kCH9
hl6UCFuNLuNnrjmC0PoshN5nhgKAuyMjLT4EZjYYcsbzsA8bBJDrSqDXi2YJq7eL
FlFM4rOxEeFmnodw/7dhiP+HMydjeZNn9/RJhGxIBXhzU5FHpCmyyD5urjOg33d2
G11pgeFwHH4nYgr+XsaZUejHFFoI2h/bWlzOkHobK/VQQM6gyjLPwSHrLtmO+vET
C61h9SYCVmC1lt7195vmfFqrf8JYFrLDNxzqSDIJBeCWM2oO1veIYSUwx3UmEJBk
rIzOCP0Kl1hM+37/cW7L8MFKZgWjXY4EDEZPOg8yE3a8y/n8z8Z2fSZWcZuCnVvP
wKo1WI+Py3hnoZZbIKCBD0No8xepxDiwNhO/HgvrHAKziUJkv1Qxh2XwjZvINPF7
948F0jo/fl+AqgOgqb2frMsY7Wwy3EBIGC2qXD8QRwXSnpwbVTYe4PgJN6lUEmJx
goAyXgQYUDov5SiwkcXvtk7q+V+PT01z2CcPYDy6ifirBNYQ84435sosq75MtM7a
FvbLkDXZhy7rmhlo3MepQJdIOvKpkJ5SQt/zBUkl7XyCsjEUsspW6hMxAC2V08ho
SQTf2LkWntyFU7gPbNs7hGyrAjd0SgBGmDUytIoSHhcRMujHAbnHjlxOAWIDCbok
sGs+kLOr+WBCu9WJRAy5m6kvjzYUxcqFUslGLc3b6+xmgkw9DlIVVPKpsuh6/mRh
qOxlG5/xp2WdKVNbdmkcmkTPTUv1FEYr149aEH7aPRDkoH+k7RK3bJn64aZtHrao
Nn2OpwQqZQJRpc2z1KsowNcJvqy44DOpK++48R86OAXzLdOUA5ZnRCPbFxxXgbTQ
id3sROXdzZyKAhn8uUe+QxoqeOF7+wTe04+2ofB6Xf+UqHIsgU2lejCT7vKPcY/L
Hp4/jf05aTNWXbwJgxkTmKntsdNVt3S2ZoqXwAUsfxQtHHYukoxrtp/vYkOwW5Df
ygH1MsuXZOK9sS8IsMEABA2CWLM+ObsSOXxoHe5yxtXSVCpNOgMMhqt8Ck2kY81w
9SBayn3xZL2V/orJIr1ldaI1JIQCpKq72ld9XgiCb+O9rKG0sFPV1hV4+BsNdxnE
krNUdoqR/PF8BQnHod0Q0rC1FAWdMkabSe8jBTq7F9MlYRp2ijqV0QjIyAnwNBsD
sMaHnV0enas20nIoJjzbAeXui34hniJXczWaUy1AuVoef+lCYSfDRR68H9u+UFMq
nMI80uSmLHIYv68CLR0VD9vlnsH8ycwMAK0rQpG9PSnZ3yb13x4iqTw5pR/nDyQx
lE7R2LrPw5ydc3L5WFrps3m0a5LRaG98dYeKsJNehw2WyyyzMYyC3DjDXPiPQ1NN
sPZCLk/841E31JzvSXeo5M8kMK33IovLRF005gY6QTQiQ8qHi1WUWUlV1t+yEy8d
A/LIw9txo6AzRqolbVcN98z9XD8pXBaNMIW8HCnzUWr6QuIbWWrZAan0Gd9DuJfQ
8TjSb2yXaPsiqw42Yi+DslRdM7ESIZWx8BxynRpvICYdWupdd6+NO6qAsv/qQg9O
dhkQBRVmgeUI3DXrXAQDYDhd2M8aAsR/RybIAYC/mBKN8z6yIWtWmJsIL4agu7Di
YwDb/8QapcJZn9H59rWet3ov7DT/6flSktyHXPydtsQhr9lqXqp46dOJyWyekzMk
HpKv6axRjuWKmb3udYn9tyFNuvMS2H5TAy8p1SssbKYc5o3K1kxW3zwMHuFLMnVM
T+eRkbP+90oM5I/dA01DmJYiRX7oI5LUkM1yBsHEOa+uJDteGdJ1oX/GOBhfdhN6
ap3/HSuu69J8bWUw4p4v/i3ggecebNJUlHneUnzkn9X62tXixYJQD0Y7ycK7d56k
VpZ0yOTOWxiqvUW7ETtr/09lEnirOZ/eY7h2i7MMaRNN4RHT3w65azzXVAdpYVlj
6srXHKOp/NDed/MKLatu9FF5DrEg3OA/9l8U3u05TgkWaLJLMqXNXLhK5+Dh1O1B
wZ5+QlrDN4TehRrtsIjSCy42APvQrsqM65GWaqHRbGS7wIQRuLFNSB5pYVMsbil5
Io3jz5/N1IDh8p/53YJcRUcYLwtB3bc3yfbPd6tzxUFw6OiJRCx4gVUV7lt/iat0
ILbsIJaF0CHhC9KQlUbGcNPrCLqYNeQ46SYW3IGqaZHYW4QeRN7vafPdHUHGNMhm
LCTxGnayYF2e7u/CNemFRt87ahMWqV8XKyUlLblrDv8Sy3xdKiSY6AEtcxrAdFDR
QmPrsyiAZSSC8pb2VV3ouiMLkcaOb6JBoX/f6nt+CE5YhQ0s0Tmd3BhVJsTVXkqB
vBHIxJJQ95uYLg/8O+6DztJkXxYt2xTTTAYwiRjuS7guN+3dYO2RfPE/09Pfsp+R
5oBXRsNgQcr8WIGkLkj+fx5rLx9MES7ZFvFDQMM//cgdlhsazje+1cFS9Tg64hPt
XIcixuxYRNlEW4Kf6TIjLFCI/ZZvp8BfqK65KxLipRoVBtvAmitH+p+PMlUCT5Ex
zEnfxca0qHG3AluTlXkoKe5DNf369R9W7TUuAz0ag2AcJSqaqqyiSDcK63PNZCF1
8So57zDnfhcQmw2DAeEmj1cO0tlncbv6ZyoxV8KvLw+CCR6mPYXOMDLATTJJ4Hj/
NhcnzrT4Ylq6wHarm+chBQ21d2IdQfiOI0W4xZCBWj0+RATh2mODlB5BOn4F5URa
TXyGnFlr6+gmRChUyrOjWSzASfV8P2siUzp8D7bcFAUsN6sZL8wRdzMgJSsYtJVd
jYUjxHJg4CJwKxBSf7FcqUbNRdAXrSfaJQlnDTQ8se1JF0aEfVDuea17jqOiXo5n
OY+W62TzOk7nMM0crTNqKcGjhQGN1knWPBd3MisEd/cmE+8D4xLh053m50N9FqnS
Oj1zKDqUOPgi9WfVg/HZ2Zc7OiBo4vbmuPjKDf1+CBDRKMbQbXm0PaXMzSJiUrUv
eK0x5JWKB1YuYshAG4YpmXEjTGA23y+WEEBjXG3aOMkCbTelHCR6kIEsZ1242RtC
jtjAQ6Jv0TrAVQ4PS2wzKtDmj3j77szebeSsKe6imOCXdIYbElqP60RTpp6G5BCL
+CelTga7cFn2WHxevGI4x8sOMRG9D0ZpAAU+KKyUXq3Nwh4MocTDyO8IVgdINUm4
IuZL5KF3XNyQZhlFeoRT8WQmLBF7AX/krDxeZXHrsQSS8kPdxRvNyDwvAPsQ1HWv
7+JE7CfEmhAgchOmlW1DgQBW7YaVHwow7VheIuJsK+a1FWLzZ4xwsxjUKymuUKI/
omSsXlC8Lq3t+1kHRrnJoKHsfCakjaKfjdHF2v8R1P93AjuqEp+xAYfTI/GxGYy2
u8mTMfUYscnew4KhSWLqK8RvWRhmIehzr8SOVmbt1mHlnKZQ8rRhdVtwJrUyHbE9
ekHXL/c5Nzis9zoPiEm0ihdEQZNwH7FqW1YhE1pV3deBX5wYPTFV5ChuT3tV2XjO
OjCJE7ItURQSo7+ht2EyaB53zT0wUCeYv6IFOuo7pojJY9vgh96+28g9Ro6yr6QJ
8QN+PPTPMmqCY6bp64vX0CJnJKxEplGqEoZlB7D6Pp53WCyoZdU39VMgHVl4SUq/
N1rd2nCGCzsF7BluqUMuEtOliMJXod3qJ3PADDnw2dGInG2/2pdxncPZCMjBum+L
ECRUNe1hXiLbnnWIDkhJ/6Lx9hVUzOrfGrBANdIUZnSgWi+s9Ba/hOg/ALAviJ7P
bHm0t0M2y+gRuvMsQQU+6UPySmcoNRdq9dwA3rFDQt8uA8DW5wjxlu1014wIHz2r
wfiDYRl7rHVkIXTrR4AuZ0vvWRGYmNL2prcWe3/j8hTaln8J97wwwDuom3DBqUWw
aKJeDCu/LgBh05PfO6srfA4zcckPVOyCWUK9NbjMtL9y/DbGChFLjD2m1Eahe3qj
yDcpD8pEF/Iprr1Qi1vjFFNX/NfhRZfQr9PF4ly277Z4FqPsBQy6sjFqF39OYqBN
UG9bs9eKf6sA0sToVycskqRPMBVtV9oV1orVXyII0MDlPw8RzODZ1X8gIl4mrktk
Xmef0Xk870uz5caBB5hJMBVBG91JrutjMmk03Pok9PajvgsyFc7YSIk0y2tvrEFm
1dc8VByG6QP7/P74FCS71nP3cmd4s1O6NISe/mNKxO5aPBXrR0AzBqDmL7TAYO9a
7+l9qDv2lEkyWQKldmXO3HW8Sy5DldR1kEtGaj5c28/Isk9sYEaIeEu38lOXdq4K
BwRgdVwxGgUcEjZYBKlb3mapsNe4aTtebma3yms1zuVdIpKlMs8oCZ+cJH/h26i9
zUuskJzkYNB+X1AJDIQKsokoIwuFUd4e/E1VNM32Hu168f7wHi0XhleJkaa7jmTs
/MpisPECauzqiWhM6ss0Fg6sposSFo20Rsxat0tL5EBLTjDEiMbKW1Og7ND6W7/3
eagnsPw4Nr5Wz0rTCTqOOSirDeDW1DWB8rUnKCgYMK3ZWrNT1qK9oQrUDlVgdW7p
aS4In0Zoku1r+r+2Vaw0sy9B0RApTVn22XryAshY4iMNRipUblaHvxhtUbQ9rg2/
VN3m5WTI+dizcNHq4hzFZBsw2ploSuGQ9JutgvTpMDZT98lqzv+tBdlHqgSsDMZR
LKRgoO2+oQchZsWR3k54ftzQhuo550NYIosy5A72jc6i5Hyex/0vO2rW573nGd0G
wvoyH5hw8TYfXAwgle5ASwMyxXz+x2wPYTZ3sFFBpiseucFyg995zs7r7GKlMVyE
ITOQ22lpuS4Tsk9vJfbRvhXSPCrsIA12FsD7dMClCoIM6Oi3Hl8TCrf/TRzFWqCT
AMNtYY7lgDckjJ4gs6RakCdfrB0lIxAv2c//o6v4sQErRVwwCJLcixr+RwpSeoa5
P5pezCVrgHjSAKS83xLzcm+dDnAdQssMCouq1N0uAfSmTkPMJc8Te+M+X59fGfEf
7aLeRR9Z5XxByW4ubXPXCcm2eApes2HJQZ3JwK2C/GgMKv/AirkiWFqzhFVNpGJN
vyMopIIRCJXlq4QXYvod77pMiPjejN0WJr2QiGfN66IDIPL1LQVtmQJ3ciH+a1sP
pl2oaIMU3egxKojXuSvc5r3sCJRL4DzcSevFzx9aA0/Nzn6DeZoGv1hoJxWAJ9JI
vVtwZnzeRwzjPhL3m0hf3usJLJVc+xZYIB2Y+JczS2rWK1a2eF18Yt/jfL1mRfb6
NDERd03BQabBdOZHUSwpMt+aahTEzAUj8NoN2XzHCGMOnPPgDXlQGkZYgOokXSFs
U3x29LAtN/sfaxbt8WzTyi4Xji0YAK/VRzuAaWX3pD/tNoz4U0mRhMXX/gq24Oxj
1DrkNvJhAyihUgdFVtxTJbWUf0g/mHol37JofuWBo/nDtGWlnqIqUE19mOYIDUn+
P8LyHPS2nNDXJUOVTkXQjTTxyMPl21bpvlppXXFNrIeveOKhWwFHnjCfbEifnNVq
urR7t3ZOJ/K7N/rcG+GSyNlbCnNFwbzrscnfTskZaXdZP8P06oUQ0Vhr3qoZJDEw
NfHYlbQUVMmVoCsAd8R6qT/yNwU40YjeZ8nsS+khdOYFk/HlbyrMqvIBpIpz26wr
7PSiZZWMfNzZV7ygYKUEZwFV09qwpkubAFKQACIyEdTzi2kNEeWlruhOUMQgzaaD
OuQVd3IJPGcZh/C4NYM8XHsqukEeUYzwoWcu5ORc+UjBErYcxsnJ630+fQcGunfq
fjHHTu1sOKDpVX0/3YS1oGD9jSHJaokUPadhT3IkknauIkpje29busvFXamff53V
Zo7AnFNbZ+8cK8CPOYjr4jpk8iLxJseLOL8ki7KF3IhIhEqOxdoyERLzQhXMeE4s
ryDBrbkFUGry3+lqWlVSDLw4kNJyhNsIVhF796lTdK7kP9KhtnFvjHnWh31auYKH
yXMmm5ZDI26F6fUzhTCVMD4vCH/OXIK14P6ycGAjFAAZtOevaoaIxZAXk+F4C9c5
oWeVHDAFXLCZUXE0+X7qbDT+cfCpcY7ZAUBcOccdgR3HPQWB8FHZcvOF4Z+3alxT
poq3aczqDiqBjvFwyIVwXbzSX+C97ni219c/7UBkVXjKMvYGPYvHmb4r7VRdSiDo
hd+lex5JeQOtELL6aX1OGOi0+4IsIvtGLp1BvTytVll7/zxMr7DojWqegaUak7A/
NsQsSSfeRMl7ShdFI16ekSUcqgO/h04xE1bgPCISUJwIOqrywHQzGNM6AeJr85u9
f2HDGmQMHKpf+e5Pciz4/K6C5gjnnpE4BNOuDcmJv6LX6tmgGb55LjYi8XCnOq4e
XVBI8VEbDfe2oODO6p0pRTm3XiRr1K6PGCJVfH9nOstNjppH09W3cJ1p2R+gXGEY
pEkayiexMOl5IV258PzFMxRCfxadAXEf+WknKtkLYWwOKDmziH8nsb6wGGqzbchL
cN3y/rlYcDBRk2vQvQBsBkPl8WMscaI3CtYxQEimCAQwGSNc92plgjbctSlmw5uC
hQNwlD6ZF0KLoWzK7X/Px/XPeUtX1+8Nyc/RR8iDsf/GPM5YclCm9XkURQABYelC
ntzlwv67RRzEMnatMd6ABfnvw2rnStIIjQlERZxhNfKrTMnVuYspzFIewdSsjMjM
0Yllzx1ezZ7TP/qySq3z6ka0NqWTU88jtOlpVVoQYplw88zXTXtMC/y9PhUpjHa2
AhWrDzkAW67pGnjKBde6q+XjT033IGBf6huPOt9bTao1ekIczbSMcEqhFi94ZPQW
ZXQJ0h5leUf+mrSXZDaBMClrsxYUTOkBeUjtPrK/VySKMWQ7nX0DhWvikffsoY39
ORGbwHD3FyuyZHR02lar8qd3/UcSSypYq/OrwTTAuvxIBBQpasCP5osDlgg9r9Lq
a5ToGqIUnxZKDIrcP/sSfWHwphkM6CGCHSZKFpNOLDBYfPgeiXs8NHVuRyk7wzuz
AQHvb97e/MpJYjTl9xF/fQsFlGm1YZlTDrIGO2ISOpaEavKD5H+4NNrTBN8YYU/z
+Rx3sMj52RPIkbB0suDIcjV7AF7g6htR2v1N4TND7jvXmP/pQaM7hcLQItAZjoHP
cLNHP7/NPGPS43ki+8dXh4eEshnkgkHFY8qTWqvPQ+ZdzCkFG3ytkvaSO+ZkWS9q
5yD5msjOH+1R6yB5RVvkFgPJCyY4wcGKcz2RZTm6sBAQZW8PYjkRhY+0TSQfj+wY
l2QCkKQyFUDpu7FkRt6ZJvUIa5Kn+L3cDBhVT+KETUBjewCPMIYhWku0Ko26Dsjm
BpEx4Mp94G/0xPzSjihM9YsmqqNXOdlIcWW+2E9lUC/2cNbqyeoeMH78KpvQGNjq
k+sM4zWI7yJOv9M8UON6CPRture+BT4EAeQik+eicf8V8EVzSdNkwDXxqZZZc8sN
KrniuPSAquop16GP8qG1FN3ffjAZ+HQSvUze8ouvUIblNi1NBaF+mXYwP4+Mu+Ua
Wdhel7sA2ThspbqFI0oVyLFgiKxlzgJay5+8TxXUlx4GAELjI10hR+h5Vhg51eTR
oCcl7zRVnhp/SMsE70Cxxp2wruymM6KFvFrzVYqA/3c4xaVt6mBtSPgjNyVapdVI
aFVLShIpwMEA+ubhm3OBvmQ/JTfS6HBzzpHOPu8QOV4toHtLL/3zwYzJMoRioQZg
gqB50NB3OOgLDwA8tYgTh0mr2noKda/gMVT7IThl0R0vn39/6yuLzcHaVsFZUIPA
EeShj2hY1aqygBCT7DxBa+MsfE26h8NxMUkJqP0+B7RlvNMZrTGTdybioRiwdkna
qaORLRzPwiviZEx+axVnjFY30zLUzYbUMiFAbQch1y3dhLFMQ2/G6FNnOKAm21WC
yUGlPDLXYZgCTLE38tywT4JbWw8lTzIUW5BBSGWdTht/kQkj+CsIUIATdSdVATbc
aDUPyBhA8AZ4YS9eAQCV6iffJHtn646QphEyOV7vwAg3LN88Oq9JBcw7xgQvI3Pu
+lfyEu6WVJXC6r7KqEgk04o/L5tDDoJw0qnW/2zJ0tQHpVBH9bR4dOnAinQw+dl7
kuikryOM7QVBjyrX+2hspCg1GpvEU2PUaK5H4711RlNFxwFko4n2GuIsZsXddZMH
PboYVFE9cDEgKTgFOZalPDbd4Iq2p8Lz+OLJxoJVpqPyoH1jsmmpkXxeUKSuh5QD
Sk45oAe9X80txBNr67eEIsd1+v2xKtsHrZ64EGkbH54mY8H74Tjb96og7YveDHvV
Q8yh4QUVKQ5tbAS5nTle0tQkB9ny8PeRaQ1/I4CwoVZz2qzSjRRQ42Ryvmf5vvbX
+/5r6/Y2xZR/VnwMhbF0IvxKczaKqunJLYGm+BvG3WFbp9vmEOu9EaiuSIN9d2fB
Ojv4rKrP52sK3fnLEh8sL08A0C8bsHSCep0XD+aUlYXP9sf4Deys6WdDsk497RC8
wndpT4OPZYBN0suOjIukNofPuLjQLqOa2VQWbDTeXVyCE5vQWr7VMzrbO1NHVZfm
qWdujq3y+6x4QT8jGr1Vp92uLwhkX4YrYfFkOH8SCnRON/5Y2+g7xlbtail6Z7eJ
dLf2qbK3afY0/EEg9pl3W+XdGBamzeLKbIqc4wDSvBMHw2kcsOLuLt4sKiyz40Nb
W0h45wp/x3QpnSQzzHMBJEygP+QPaxjJSIhJ4mSxawwzKESDSfuIvVWP/m043kSt
fCCIriuD9V+ePjDB7uvY5WZQ2UDlbMOZ/xpHidaOmX92v07GR9gqyEG78GCwOFs9
N0bpFldqpLAVBs0ADpqd9FmolEbKugkQzqj3WjWhKb2N/j2fb0aB/esn2AEIerbW
QUlfZdBq8WwBYxqoFBfLkDHZitf81sRpY0itHbmwAl4EqqzR3LdJOUmrnQR35L5Q
v6yEwWd9EMKuoGou4totjAy7EcN8QDO8aMHtdTdy2jN06bZ4b0z1NuvZKlLDTJQQ
f0f7Czkah9Y7AsMJeU2hBgpu1LFx+eGfVA8A6k+Xp6rjvLmfPuYAtf7bE4Oo6iCh
g8Jfps/AcwGbylKTjNH/zDaJ4bGiyqmBBK9RknluynhYMskLML58QPgNqpMBytEq
XgICG0qzkMn797RNQFXhl5FgQc0yoLJadTIslJC0qwcoa1cpdz/2VMuWsoryUJrX
0m5sQW+ppIlIe14jgl51nn+FtA9NDctiKiDWU4nk1G34XWDb+TYc84H60d4+NJiH
4UMkl8shFl4+UsqF+CS8vJAXCRul5DuZgDnKzGfUshnQeYJHZlI6DZpK0bhf3xQX
7es6NJLLt8vBmRrRrk5QvqLVR6WqVZ2rTh59FnhLwhmyWu9BNYSylBFRFDKqhCQ3
xYs92VmvZfxbCe/VQVGgHTwZAHlSXBAz6v44QpAWMB1tsEPbeafq4o/M4f2q59ZK
egmW9R3+dC4WV2KYJDscU2+nfZdkNaA+rSGi4SVY64QX3V9Z957FD9XjrmOkc8jI
zi/KlJANik+kuvLmLl0CgRmRuu4kw5SQizRLUEDOjbx81R1rgH5JcXXlr8xfgutR
9WcTN4pK4LyNG+wVowT8Y/h/TYM4quwFzZdIRpBNj0lhgRQkuKe+5g28CTOACkiw
kuPDwhTF6/Hie7lBKd6LirS7h80rwwoFdcVEdimCyP5lrs3vlxoB8FlKT93grOya
eNraDhqrzLsqdomehCtdhCFzE0E+HNM0PL4XFgKTPspeV1e5doo+wV1I8TlE1fjE
eGM6aAJsmaS6Qten7bL0sZecYgg1kN8Vznoi36Z2MA4cAxperfAMjt+Ng5+91RzP
UWY0q+D85XWGz+ITrfzeUikp74d/+tpmjw+DueEZp32V5zMkXXi3hEvMskHfJO7S
hi4HduIBh+JHyladHvs7t0JXPOJbBpNecsUgH+yLnTacTUJx/7EiEaNbNyyJ5zki
QmBsIvJUj0NvmvI8WKkvJkVch3yS85drJo/A/T+kdJG/qaJtcmCVNnFPx+BYV07c
JBt4WXdKVE0I1Lq0XfbXmOs432/ZaHlapmUC5FHFa7thQ70h3fWBDIPcsoLkfqoz
Dg/hUwmkuYL7v54eYOk4jLFHRWDDpoG01kQaH9WLQzYopUp7lADizCLc87cd8TKV
07Vhxubfn97tQksSjRJGrIotu0jpGJBJF3ILaiq/K2ulu9A5ecvU8+Exy6v8nhVw
oG4gZ20YZD9V8jtU6RfHymlFOut2s7pAi9v9wNdUJ5tm551FksXg1PaOlCmAfuiH
9M6skhUOspNJLGYzb2JHU+fZx0qphyUogwtLqLdAe5OGGI3s+7/puPHhqXwf4NlX
6Ivr/QR3hN2ZrUd0ZxakJydfWsLLjJB6MSICZNckU2ur+ptOsvJeOv9JAQ0NErE9
idTm3MXXA2lKgZExAcaIvTaKl55Eyr7iL9a6NqiEIXnu866OFJymimpu1E34UlYQ
ySWD1VGoFQtaG09OKjfjTmKpKdlCxToVZ4RfKCvjyhXwwHT396RPeRMnhGm2edFA
XZPV9Cy/NSe8zhRJd2dY6cP1GFPoNur84sm9E6LVJpjUfj7k9bpKYswbOtGwKrzQ
mE0bX4nskxYeVM08YmNi/Xtyo+XsnDbahRIiGroA6qat0YyG1F4PxhPSO5j84AIJ
YheywvtuGfx8caleWGtc8kPPbnLTaKcBMa0M/Oysx75aQZ/BW4LjY2KHAXoRr9EO
ZRZGKkVfq9cpUJqqdOFNsFrTqgA3UytvwrmVt3dWaR7ZFvVfU2peZRvvWtZJ3mkw
EhMLH1IT4iODtvrqGZ9bZfblNe+umhpZl5O5KDwsdZZUoQVkNCpL7idD44M1OaUK
zCu3fbDZOmXLZLNXe61SbdzOhKVxTJ7Vz480DM6GhUL/sm0u5EXoV7b+lym2cMTj
IZ/+jIIlYg5H3gjS9I7new3gR11W3mp5wc1aTsqczqvtf2ZBppLQuSb6BqwNfeCA
Kk2NFo+vC9Tqn8I7hd35Fm3jqErNkpQNHtqtp0oWQqsWyEFIg5NjDZpdxNPnchCI
xauQuhCLm0wnpaMTlWAEaxA9+lPtC7r6MupR92Z9FFe5EZxa3FEF5gUAggd4af9n
hLPxhNU5AYQWad6z+gT7gsNGXrrkOXmQdTcqqAKZYiIa78haHRsWmKVrBbfz2jNX
eIJPOBugzz3i1/dNubXCqXxymmeY80JqGOL7T/GWsZLEa7obA0xcylt+aHshpiOM
bLQ8C2b1t7T/652shIr+2ylORPDRewuZmw/A4irx0AA0Z8dSVr2RoLw6OiwuHmKS
glKN+42vVe9/GUWUkA5Gk4NQzVm/+BaTayDIesJ7v8FnvkZc89MXt6qvgC0epw/s
J6YGdtBKVP6GgbZjtTGrDflu9Co9Bv/d5T7N2C2WJGdyp5YYFvwWIc2TIUWxjuyw
WE9rRLZRl5o2Ts2XMoSMUvM/QTzmXYLzz17nNbTkDXd+zDQBRLvSvBVFU2WdMYIo
QcK/zxM7iIXM38c+2LRSrn78W8OrigRy97JNKdmNrA3CTugvaiVRiPFk8mF6NC8P
wfKAfMcqszlyq1l26ygLFIzmzFdwfrt/ZC0ED3HKPp8mxeUFpHtYMCB4BvSBNLkH
m3FUJ35IaNQD9wmMb48gCqqHRP3PaKapTBykVkmqItdcPB1Mkax9dFji/MgQw4a7
pdErbS8EBppztPbs/IhyToVa0/Hk8MwCHsLq+5WPwTJoiNw1Jf0SDY+G6+U+3GlC
M9yze71HCeEQ+dQlxs/dBkj4hUvK8XIvf1hjhkPq5eHgmhLSqLYWugtk2KSYP6va
troBxcI5ZelC/nx5FHTL7W6SWJOPFk6OlV4ax81x2f41bzBpjKx9X2SNXt8UiqAT
ai7gx/hx96eoey5nXq4bG4//C6kS7ilY0YEk1p5zS+lJb4J1LAyr3yv+DKm7JuH9
6smH4Yq4tgRN29YHxJ5Z965TEirDEkRtVUpFofLQClSVO2oW6ihrBj2NgG54ix0P
gB1WulOgSFfNUSpsTt88RvYoI2YtJJxutgFxAPltmgAexTa2bM/CvTOfyK1W6xxT
bIeRgsRViGUymPY4IyX19UbugxBOfDw38aIHzDR4tik18jXXf1AFTdkh7+QmXJeP
1UyKccwMSI8+GA/Q0wKJp9UnNIPKnBkHb5B+xrVJe4qJhmB6oZqK7TM2GodFvY17
4SapnLOAzU3s5FHfn4sI8Obg8ZYapqew7E4EQ2axhQHcHYdB0GxpgZ2zSjRpCrbS
ZDKw/kKOesSJYFxz20W57rMjNXuze9u8xeUlbTcOkeMoN/hE8xwGWDjn2dhTH6ft
P5yNvS9E1VfT0+md7OlofmG6xUZf5IMrBMP2P1RXQr9v1MhoaCucepMnGGEnY2Yf
TNWGmrVdQxmKHNPsFNLBvp+fgRerng40AqZI8zcIMrKDk6zYhBDlj9cck6PCaH99
uIwor58dNXyOljgWzbTyYyZ3O7NZ9GkU9HLosY7h6REMl9ObWShzlXrY/T50SGNs
K4YSvKjBSlcS/G6vVwC4Z36xAepjXtgQVY26xxVRY7VYCXtgmXOGu6fb2hzoFSKc
JYM/BpmaPxXP5dC6a11MOSS3oo55eJAcTrz++GeC1T+NTlmLajpbmzUNXVy7EDtf
fg2YpTP5btNYg5lL5VO1wCgMbNxNyAWiLZ/i/xucrxATCfI+PdQ7ivLEqHUaHpM5
kEEcGkJ6d05zaMmibuyDtLCNg06TeldvPCbLKxveGIRvdL4kPcm3EB8OEXm7gvxq
auYudsWG+X4Q9KPeW2os7RVx9kZye1pKlu6nSvs5sljkSpcgT90/KsZiTouqrJxn
Qlco+6Mv9m9g5HBUHxnUkUiNKKVBvqpBWcHStn9nbHhTryIjqJjwAf7BbBYrc7IJ
gUp/uw+QyUo+fHAQ9ln6wr+Upc4bP7HbHLNpYmWVZzykm1CaCWH6P1gCNEuXcZle
K6hMxRCWaKEtomVM7Z2Os4VQPznoVqSUIagNGPWhj2kVJg4KWDEdEaQOCL46l9Hq
wk6eW/V8NVD9LqA5jrdUO+zqQH2HvT2UgeBu2Sb3v2am+Tmb1yCrk8P4hQVWX5gv
mQwbLyth+GEu/OQIdwi1hJsRlIDFPoxXtK6G3lwLNFkXPQwIGFSWZBLfvLjZJeLy
kmw5a2LSAQimsUc+bw3CohKODYsXwI0yiSsVujz2cAu/YlVali1QoJ4crpKwkRZr
TjjwQwD4CuKs9w3fHURVDC467jabMEJBxKSd7n9vehLsy21ixeXxZamQNbIJDrbi
GzcZYNgEv+2ddUVHtH5KzWxY7qM8Az6RBYYrKuw+uHpMBmtl28iSG+rF4kRA3Yun
+C+F6+IN9xpRy6ZF4sdNte9ZuhFPdLEV9FI71i1nyyDuMlwpSBVyGd7Cph5nAwOI
E8ycW1jAInb8faDlQjZfKtZEAqUzf2hhz6EPS6np1Fxk2R6SjNn1FCpIryclW1ux
6OhpsLuyHFaOcE4N2u1DEzuvqOfTsI8iVGhIae1lKHfATPeuh6ASkBYAGPf4bCDq
mvoeKg7BaW2lKcWytZjbdvCvG0H7ydcPbpnKsoNVG/MUs9ioWZzuGHs6Qmayh7xi
G9W3OoTBsW+VpoSmOON4R3rWp0l6E0rcdZECyXg5CxCMzQfJOh2TkWGvFQPoIdRn
0j0WPWe9VYEhQQtqC6J12ZAWOgUc/1sfPbSvflu/HnyQcdarpQ2QO0nZUMhl9BcC
BoW0Q7g3lKFMdpuaS6b0Q5uvBp0odPYi7nwLWNlfsuAjpyeN/0hDkFhKAedPg4rv
zG182Oki8Yw8Ijhw/fz+Mqy+P6Np7cG7sNm8vWP0p3RjhWzcEKo2DdkwzuflOvC7
lvt4+wbZbgTAjAmWONeSEFBTAssaFDj1D2dAfx2OS/eYUzXAgNIzT8JbS+4TgUh0
6QQ/DQmJSE28kc9A5PdmQGPyk0zlnGLlVQwRi/KiRecYAM1ZPn1Lsd4ZPJwcK8a1
I1tMyAHD+oPB59DMvWNnFs4voqJSjY+v3u0fdm5DMc6PUoburru9VaAlAFwGo45u
05rFhCjsaqxr7JFprXA2fN6div4c4RAlGn58gM+azsgV9z3YGAn0en2L6/uwafU1
1IYfk+0XoC4ztN1vk5muIWUWdZycfEcvO1a0pjZ4VLFYtWfGoFa/u5o1r8du/sN/
M2om0o02MEa1IKSXUv2RMgzVY6wlNTQEhe1NEKcfa8X3TWIcDNdKdYKNG/JUwlXD
KgrTb7yQ4JnAUJ2teKQ8/6Agjw6oZwatUZOY2yZhIwfGzWFGTmWgfAkvk/la54/0
aNg1lDSdTaZ42GsfzIrQuvI8Qthmmu6a2aT54uiHmQXnG6pDhlT/y1ftDlGlDBLS
tdrcRZK12Vxx85lxbXJ3t6kSMtLuaWoOoDyGfGavzKAPiYKFwZsB+ICHvOZun3La
dvQXvixDlteKkAFgKPamk63uwuh0M6HP/cUKx9Z1GfWLpFjPTdbhapKODEt5MXv1
3bjx4SZ1FSSs6S1CXNSkjYeE/GY35KG/Un7NvXymjFhi2zQ4AyTTIYBkvEY4HTId
6rgV5xlXxXZMzwDhomAEMdJHwvX+/IKc4CgEVg4OSIB264BVh6mAVGJiKh544JGj
O/q1ySZoKoqAZc2HlztoKQQ4BUC4CWrLU5hsTnWq66Rq1hhH93qpri881WubZ2c+
Gx4l6XvZgswI0p615czQfX/zVd11xEP7kYSCaw/q6lZXY9C4z9b3/aoMtq19oHiA
lcmAPhcZem2Xt4YpPWcTqmGEVqqRpqorFBr7+I3ci7O1hzF3S85jSSBH7hEtX9Xj
sarNwsZ8iFEkz4EHf8sc2zkC6ynwHH043SuYNl6PzQxu6EHhopNqjEIkg7h2L7hV
RU0CpldZeNWorAGcKxloeFHyEpfjwHZxcKk6sybnXt9oc24suF7cfNQ1JyC8c/O/
CH5Kug7YL4YHYpsEhbMVUJgJvvveRZoiWkkHG5LbspkmS+KF1hDlYlIc4xdOQI2v
7liewgUkwHBM8LWnqPh+9re5dm7F+3i/3M5B5Z0OPpA/YITuha476lsSi+U2BWxZ
APOFT7h7qwZxwz/c2JWOXXJpb9sACz+Cjkka1LWZThp7lZHq40FsMNusAUjeZIZn
XExS/8uf/lF6dBK01lU40nH4j6zWEAHRibp7/FMXeaPG8Vvjl2zyP+ltJ4O6JglU
mKWWZni7KC/3bvDFfsLcbom68fn/uE2jn0PLzIVmsQz01moYoy7sjkkjRwr/TF++
mca9FwvwungXLb3WxCkbBA7GVN1njZEYlOzCNRlpAGIIrgowO8CyaZyfrSzwFvsz
j3rnfH7g8FE832NMLCHpOd8PLdbpe8STUeWZccnyko7xlWgYyioeu30iu+IZ19DM
0YjaaNyUtz3s1H3bl43BwrA9itTtC96u1qhsrPVLIh6a0/LnXAxld1ATetR+v9bK
FwV2LwG8EA9jnKHFH3gUcjI55CECQX8IRGfrIuida6EoUeJa9elyjXFUN4q3Mz4h
Znyvc0odCAX+4AHT4VxARzqWOfg1/eCjCeUpYbEEw2IEqkqFX2H7OoRNYkIjXuJv
nCUZrvoIfq5GYkCttIrgW4VPX3JY8ZCTQPUvPuKUB6TL5TiWXtdbYwCXaBKJ6uY+
XqUgkgJworTulnxtAu3nIs/RsXH7PZNevaIykpc939wFwpMrLD4/IzdnSesJyhl7
HFQju36Lg0E1cLG3iINibhGsUE42/k6soAtuvFINdNIbB5Hamz93FQ/aKWwMVi4m
Hp/IqreZ6ePlKv86jeb2rH9jaYZR+UTJab5JadR2e/bRdPqk7WVCtI9aY3xIYl6T
UF4JlvSDrdw0wqEWC6nmpIYsZwQhPEovQO5hueyoSBud6C1/aybFQVUXsCJzbcV7
/EUmrHcKAs+W4xArkDT8mmt4iQ9hFa3wZRt5v2bIgAdR9EUyW/DlGBptTHome/K2
EH4OZYXrIrxqwZcP2xmCf1b001tk0S4+NfUuwYm8prjZS5JNG7Eq/vzRSJLOxxGa
Hh+nVnl09m7v2mo8TXBsHE4iJyYw+isIlF7BiYtKBe5yHVfSLS2TyY5WMSJnEn6+
j72d1Y6H4+6eAjYTjIlbRWCR0cE+XPYGl0MEVb2nOsNoJxwY2qrWNxNnL2OoDyyK
rTgzVH17EWrTjo+7QDcEl4/pw157rLZ0hxlChj8xTs46oDw9mxNzR8Lfth6L8ClY
NbgWYEAUCtLB+23gXhDyvgsozEU0isURjMIm+eTlaXw1q91g6mr2NcBQcroVUfqj
fg0O8Oj1NOnnxrPUa7ixycBoN9MQKSPDiHY4kYsJNVd3+5tvVgnpOvR+DUybNttM
Bt2SY1kmLJqtKEntFwHF/I+kGrw4xz51o8A2TUX+e768bfbyBzscuSFi5enVfj3t
xcLXaidehdnbXj/pLB7Lh9jcvYuL69yarEt+srvaeRTeAxd0UkeSJKp8Q2yjR3Vx
DclK4CqJXFDVAAKs5ebE25sIYu3MUf10mStdYEwRryedv4NiZlSX6zhnoWEiSFmV
tm9zCPbAv4I5+3VnwiKXBdv7t0m+sZttllgWBH9F8lBXuy2W6AYhDlzxdbR/P0d+
qXokMIrn6IbwuXFdhtHSep2YRaKqRZoHnTLSKP9u+7MoEaJt/d/1gZvFf+cwW8G4
8I6+HtBI5g88NMVuGc3VMW4RTaJkrYHPkjaxWC9NYaDOzEY9KXbmKqPuy53v8gI0
3w9qUrfnNKonzyMRr2uQxqFmL/b5F9XrPRUzMLV/GBY5Y+mAbIuNqzA2lqp6GKIV
nc+MhIcCbys4QDo8H1IRTU6hMG8lGKy0DLOoU/pKZ+7qOvH8qSbmMt0BMCG6MIb2
a4Zv/pm0sLflJcsj3NDxDiuDW2mjPhnYaoRkhWk3daOHQyFI2WrnseJvgutRJYRv
UgkJYVmGqxU8bRwt4DnLAJBEac1+Gc9sOrIWB8vmVqgAyY/Wq/1C0CuEfH88GtMc
yfIPltOv2Az3rC44CcxIxAB6+5cj9ZNbnyLDFdLfZN02XVCZ/Kj4DNolDYqZgzre
XMdIcwpUHnN+WxJm7lGjYoSU4YMHiTgqkpCYvNRoCf2/xiy3My7nYa5w9dNcB7dg
ggWaYJ7boLbLqYKGzQU0x29kR4IPg7OI9iYfWh2c+wYFRdRFMiDetxSfJFQrsUgj
lb/7br7ckwG2829pt91l00uuvNM+xEcBxzkvP6GA38kJhF55eX66rBgd5O4OIhno
6yCuOf7z7YW6EMnY3lASdgkGNlBB6nbmpKCpNYypK2VP8tZtNGvFXZ0zgRYWYL+r
XCHy39sssBGSy52Z0bSaWGaBvmX6J5EsXVoaW2bMSxf5zuCPMFQuBs+zONQ554Ez
5fqG2NHDV6p1R0Ha+C0Ay6GGRfR4CYYUueR3727A8V23P1OAJW3hWcMuEfSXTOHW
4wCcV2t2uxG7ot1ql+r+FDaf8usKs0pTzc4Jo0SjHtuH4stDcyngDS1wRlO6wAbg
tjTMVbO2qnHNHoI27yOwKG5KY4jnXGxgt4IXZYgZ3e6C3A/om4n/DYSMIUQsBlup
e3dc8hmm+sFFbGEnHKHF10eR90e01jAtxvMs3WGYf3P4kKyc3qmIk1DO1QmNNc9S
nqZ720+kI+/6ZYKuUIWu5z9LtAorGzVyOCbvuW5roOgbkxpw6cOM3mCKpDn0eGBD
rfG7T/KMrkh77gkLjNP0DmRqBIi1Om/e9GKMsraLrVxKr9FUIVpm6C6MXSWwzJCS
qIaObHNSIbE4+t1Ivm5t3BNF0ZlThgffS6Lr7QQNQpyhA47IjOXyugw1Q1ADVaev
T0Ue0kxlLHa9tVRYwos4k4NJsLHpUZC5m8cWtKCis9CEJPsleZ27c03HWph1teB9
/MT0E/WZoTiY0HBejZ7CnfYK1gfyMICTDk5XDTZG53J4UOehZGfxsjFT/nQRt//k
fsObrpxw/GAdLCAU8vHYAejUoEmLYyX+S/sj5ie1pKmLQD9BJm9IDizaFcBftLAY
u7dBQiXDfAWwKPjvvB6Oa1cM2u2QahGWy8cyBgQQPIJq96z2ZadGHdSr01Ntjjda
AhM+NpoFsFABidt6UhB+LnPLnVGElUAO69T7gd8cXjdjlVQGYPQLsQofUWeFDxwG
zIKjWYWWru8go/IZsb96YNG8OmpzK+kbAOH1WiVjzUR87DSpH5N+D7tQFu/0qNJ+
pnNgmq0L8ecmThs+64bYPad8FdazHIJK5MUlkwdQtUt/9mQGwcMChaJsfiqqcYDL
s/IsfouqcgTEMeb1dxtc8s0DcVjAxH1sFJGWaVo7SIaVK+79S82G+kWmexDpHAJX
WSdPQtqmCDiXNZY6UOMKfRPRyOuE55lsMiVMemw9sPSgu3jVm00zzK/MNQHlC/fJ
4KQDBwOQ70jspeObAU0ghs2BI1yccKBYbUzot8rgVFF4PBf1vhZfhKTxRtxmHFNN
cU8taQYaN6H9gCSrfuEO5A2nwpyzbXaNxfWDb5aGQWXamRX3HCdRD1q5Ca2YteCl
+IvAVcJVYw8U3ma78wJB/WKsqRcFkbB7mwC4bpGkWxluBfuse9f9huK3aEUzDZtu
khFo6HRlJct8sXTK3K6++UPdWQC+Q+7fWxW+uDcAnpb05qNstYT4GD2ExpkBDMCk
givUgeFs8zS/FC0dXFS6x3oMoPsQu9hOMHoNEFx3wZfXMtRvZoFhdqvPczbC0Mdl
49Y34t7dP5Y44wWsBnXcpsI4pIwHgP3l/XFUuKTWf9snGYnClHewonJmNsMpSjGA
m9Jnrn4MD8wVKCyx9AZVqw5COtmujgboM7E2XAcjoiuT9Q5OXhxC1VIfrnpEXUOu
WubZvW2cbOo9GtscXFjq7gE496fIGIwlLI0KCkdFAVKl8cwUG/L/VFXeSl7fRJki
WvQDNlGwnQ6aBolGLxdFD69VCnSVLikHJPtfoIqDebhQ0FVRWXx+alpgpqTXjKdF
bqs2cmm082spA1vK1BsDf/qufk7q/jIeKF7bSbSFJ/eInkbfT7eMPx+Fh/uxZfwj
YuCEJ1fZeqx93PhtKJPvw+ZaJsj3fS0X9/blZOE8bD5LxBztx18K24O0Rx0i55th
Zt+LAadagQD4whfyqCwqjfnnwp0WoBtPqY9Nteo0ORSjzXEQzcYv5yj58xCV0jfU
kQiiJuXh3rEw6wElikgEGbVdMRkQn9nJ+pj+8y+S2c4zGgLDmghQKwdJ6nhyKGl/
wYD60kNSrgidsFjI+AmXVgLuC0L4lGiJ8VyNjp8xi3GtfSMQYnxa+amy3S7kAAuN
4pKgefeLP9sPtbByIw86Z9tuQvyQ12svNNdPHjCL78zZT05QNGyACwH0zi2Q6+1K
MLVF6PbRF6q55KPVXbIXnYvNfnnhTk4bYN1gsdig0zX0fUzksx2/7215TVYNiUjO
20xxaAvkAHJXTwV+pqfhylIVvto/Kgh0j0QsTpRn/dOiUo8rtNDhmp4rtGRfdm6p
6I8iC5GfPwHCOJ3Aypc1UDCRFWOzIsq6vhk+FXO45sjr4TDWY33x/HingXz8726r
AGfuF5aGozzRKaH0yBQZLPjhAjKD675Ak+12+IQokzNeERnGeE9px6VNj66N2DoV
MIumcNEckaPIoPqc4NgC4DnD1R8AsI6TzNNQiFGBTyFNfRiY21jawGsv0nBACt7A
BpaOLzAYQnAmOpgQUkNxB5T1TUO8Nfu7rmU1VtNVodpDUJRv7MvrvrteSeHKKLgs
zBhGQTHToABW9Jyj04VWkWh6YWQ1R3aGmixh0FstYaBnW+1jCu/lL8hilfxXzZ0p
ydNDpbfhKe07hwIBxpJdpkNpHQvSRljToBBrbOYFmcYeAwn6BektnoVR+alHM+h5
9yKWeT0bAuXGNZLLoQcxXRt3/dQGc+lwO2wXyOjlmxN1CnoOul9PX94xlTo1OwZt
xiLsVP+YHAUBLYFDi0Am2ThP1/EegkduJIA6be8GXC+Vxs+8DOFg6p1pu6lK1X6y
1F49QFNoRP+VOF3gRIQ+yzmOldw19ONzALHX/cn1bbbxUUQvJIN5ZtVQpdwcIKBX
t1h6BeiKIO6a/LvscBb+lt1EvbD858dsfyEhg8xvkHvqsKa8vKKr8OwEN2LYr663
PM7l/kTWikM3RwxVFEsB6IUFYJo9kRuNHPPYHSlBZCwp2tB78FIFgeVlE5iXhKA0
1dV3zMjLZynfevhmBAQUXAQ0FTr5mF5Vl/2FH7IBt26Ot15/dK1h3fpo0PIrNho5
7n6UCOLsvnaPGpLxXlgXwN/GPxSRTi15V2lQd9LJKFZpdtE0oktb1JEJlUYshtAU
K4ipl+LMqYz16YGhM/oFWMWyH+neykHSf850ZIZiqzP5fp9tgvoV6AFHLL8dO4ZM
P4pssSOyPuTAQd/wyV4wEzrvDXP12pfn79uQzdFFnSvxX3zWCypBBIZVrj95DBoz
gBRZaELRp9SV+fJRnCyO7+p+i9R6m0cZphWaqDaQa9zcdcVO5xsFEz2LxXQib2pa
+H2hRPhXClQ+CBOnIcl5w74iorag8WsOxnDb/25vdjCSVfuEvLvAoMXqZaGNZSTd
mwqQ3ZeJ8qeah0p8fUjtk14gby4CqbJydDwQBFdluunJYbyKF2xzSKJv2ll2aJzz
qPXllfNPiSOfcEmqpd9Wc1JAkXBphVo7VYmTu5fOAcrWwoJu5M6PX8RfBVOI0H0s
I7erv8G4mtvJBeXEr6f7JnRiOi9pYcPO1cs3PYv1Ug97AMnzdtJdxyGm16qGyID5
8t82yiPhuDa5eR8ITPQ5XPE1sTsFQzxRtqIN4vHpy68AvYMXuxo+6koXRwrws6zz
C1GaMYFh+GVGLjEkIhohR5d4p6cT0XMJtesnDqQym989jrRb5IAFq/+XzQuRTvC/
xymxhOaOuRLBOyHBaNqufxBCBDmkWGapjE3Ytq3/DquL48wAlM3HG/UFz2nekgHS
YEx2456MvsN+Wtmw9cuTU1FhdMfna6SxtT6wiErou6liW9ppMYfLjgXLxSQasFyA
Rfcew+l2nyF/D/ZLHoalI2aHSpu6NwbS0Dj2o+x7u30YAzbVG/NpEv6y4jr6t+Ui
uUMTyr3kDBQsbiv5+wKp4mbScm+U5dzvOqJfaboljumya3r4NlR1BzWFeM9dDRAQ
VcBmvxfFwhezLbnC0O4fnWTapRqSK1uQR6v8RHE48Ye0rTrSOOwL8tHeIwydYlNC
Vpuim7IFWdn8XZPE3EygGaXolPDcjFvEKhXlB7G1IS42uPImNNMEixQxPG0Bb9v+
iMBtOsAsB6ofLO9901/9owOnI/he3z+4Vcv5txayOzAUudRqqilgFnomGTiuFRZ4
ulJuxI+BLekHT/pHwym36iiAglSeK/fpx7XeTlnj9AbzmKJPYviC6tehFHIBxHz5
sJsuCX9GyerkfKOB4XkK9qLkGjcJBmveTDB/bNEat15qXNkgEFjS5CfPyqiKgW4r
naX7zeiLaFdcY+w5f9R3Ungrqbr9SEnfe346ciX5UrFzo6F7bPJk7/Be5mPAjDC+
EnaP66sa8R3Xl8QZRuGRvyRF+Q/QPzil6NvteCSdXVvUV11sLc7qEodveUK9/4pJ
KBclk5b6f4q0uWf7OS7J9M+CGHLlIpcnpnF7ELiAeXyZ4P9oIrV4BPLcuBQ4yKch
cDzU0PbIS6stlxwQlJLi8NBnJ04yJSVcwZ6nVD9SgKP4o+vO8sXY2im4c8lIt5N1
6YCfbtOYmIK+PC9dRb69e65ZaK2kig/oqTPq7jmlGAIw3BFR9EzH0H0crKEAtDKJ
PL0w6G/+UCrbSCSCzTsBpnXd6Brl8Nh4TM23KjXqeosTThLs2CnrNYZ2WfRPLdDr
V/iLcGgWAdBdpnnqAe84m/VumTjUNsvQ4AnNq6abyVxSIz20VffHM53F3KYWAu2U
o6Jou3Apj7uWC0SO6kHe+3zbL8E4GxV8TW38b58opcw2gFak8Fm92ir9ls4eLqyE
iv7LAsWYlVO14zbAkBfWabUzXoHERJ2NtpapxS0T9Qvdyl4ngeJ5msa8z7Cjbpj6
RkhpQRz+TeqBs5x90LmfkQy/uH69e96IbSfj/9Gwkr1ueRsAKeu1+RyEaqYjIFeu
heYjbNpPznIupw/emx0sygsMfxnnD6BeUZ5KzIDLb7FxW9V73mu/hFkDMhYKnC2p
Mw7Dnz3MaZmZfFiuj/dvKqyR1nTw4TvVR+TJlXRI+05mrT+rdaixG60WiUu1w5OU
TWdZqiIW+ZUc0qxuv1t0E88qkgsSFU20fd9zRi/RK0FBa2s1yhsjOCSJ/MaDU1nZ
O/IHyqF7BZrbBB9TnW1gCCnqmz6gHlTIcco4QSUjOvPQXpiI19hrFXBf6YXi4NO8
cfsf9nw4qCUzShzEOCTSgNpeLAh+/Tejk5vOdHX7jU6gLKe7arzxuh6D4Dj2qWEt
u4BPOhRzL+zzEHPewPh8bQ3BPXxFWUDkj3QJDqYhlKhhfXyARIEbvyLobtRAJAKF
2NF7CfMBcUmtXEF6+dUL15a0C7xYl+EMAksT1ljLWcNExJO7Od2Wx0/O6XrJP9qX
J55g55oBeI+fAtZbbIMNv2PfSnBi4BAnEJYlopr5mdWDRlE6jHt8pQ2+PUyOwbS2
xICcKUrVFSx4fFsRTeoWiECJkrwZ1vo6qNq6SBzQMmgmsNZiGSArVftbvgB/uPBA
hP7A7EUhOqE770iRvFsV6vJCuhh7/hkUALopBYUA7djNfoBabn/5m3dzofBg6zg/
tHt7zp2Rq0/P8ST3A5v8xr3I4x/Gn4C+XjQhcDDNuAKgI8D8SjNU5wyes5/gfksB
2e8j/UB0pTxNHgd8/MRdTXyvVjBkhPYrxpv2tabcjScsggHqcA6svLz7Z4w3/ezg
NdQjC2MHYGQScB+TVt1VoGjYYD4VBvPZFr0Buaf6gDGT3NIxicYfnWh60/OKa58J
oGgHYAJpuvGZmUoMaXp0NmSrtOtYy+Ig+405lfolRXJrTKOaHyrLhvuxIG0Dtpqe
ZJsZk7NqQHbGhwHENqbP1Wq/swcH4lQi/PmgMRPabxt0ot/B+1/mUEpGIraR0Xza
qXglW7elN0cIxZ+B5RM/faphRf826jrzWl2UULEERlFI9yf+Gsgse0mPLaLz+nJG
vrpUU9aaOvCE3J/+kMv6AfRWXewno0nrQ63w4496SO93F42dWt2/mJsLtHtlZqm1
RT+6HmJcFHIp4pxbYtFryauPwlub/tpRL3GkbilUQFN12V9NxnjfiMZ43RBZ592F
wW8nggORopyqTKI8tPYbYnDUIDtQ5X527xpsTh9uNrVA4I3sC0XBaPUpJ0LzUqpz
NPfxr8oWlVfAGqv8qpgp8dbJvyEptPpBz3GG9hNc1dIzG1hKe//UwrBpfn+QIjBK
S3lnozIePj3pZJ5m30xsSONWcBuOZxGkIje70FzJBAF4+KEAkI0bsko6VfMikBnv
5O+PeMmhqJlExXTxS0Dw5RAdlto/A9ki+hXRd9xKkI3ZDMIiZ2BPD07iw13qkiBz
S6EgpRjpRx1p9JNM9MRAZYJoZmU8WAXtfIQwPWtCv+W44hK3q+Pte046O2b6c6Id
60OStBGp9AA9CXiPaLvgHH+IVWDsJ0z0P4yayCmuGKYZWGuvansk6t0DnuETdSjz
Xxq5oet/Dt+NjgMpWZZPG/DQzVAhfLvE1xrgmAcrSC1itdy7TGOfAfOBMlvakNqQ
wy6WLeeuphTb2ksvwj1cCecSfkdyA3SAA5ZenSM5xdjqcXxQ3XbNx+CzUGjb6OE0
bj2i7TMsN1nhV6tmzvxEO7evGPqSRRkeKxl+WAjOTSgOV1meNZpY4Mhu5wcRmhcd
FISKUGvzg97rcQxDtjMpLjva67DbEmW0r9vAJ9zXgGFVHQERicHGXj/jsCNUgxQ/
+onf/JeE6Kgtepa13ePzkcC4/e31ownfIgj8AudMnJ2PRRnBL3vL/LLDUmqeck70
ibJ95jRL8PqoHy7b2Ftkai3O23W06/d1fSLFAp9cnalq4HewrF+G58ivhiecf5r+
Zmjt7z4Uk3YGPz52LRg3XFlvyf3gPFYzuUbsVuoOesQdaOu2n5j2vb3to9yhbjXT
RpXVnnW6hbk1nyxGiHsHG08mMOTHPI+ewsoPLIs/0kA4uyejrn5LoYmJWdHjdS9W
o8bUGDVJGviMHJju8Rf9mTlHV5k254IS+Ule/AyWzdU7VfmKnAZ4tzQTKjfWCWN0
MNyC9lPfH/SeHIIOgzOtr0VK5y6owUdfxBXdSJFc4z2Ylqxw7GPIDVSkjjWxY6Js
WPhriZFftYzVFV8vtf7aC2knQwt6g5yd2BFb+77BU+yd71MmoWetwoRHFV6l2hUI
q/BzZ7FqeJ7TF5jQeEBW2RMFVunFigCtNwvKXWhznWPzY3nNQAGo2nSX5sbXI3nO
p4au17NRDhzAm6Sl2c5UIncc7vvkr11yCG1mUdjXG/uR8diX26wP/kmPUcclM5Dk
u0lNYSO98fUGHrhf6VJCRSP6C2FLJLUBLvCxnXqjjVEbBAWOpBgUTdY6nUHKTi08
Wi5X86M/6zT9ERF+otQuZlEhRdoO9odKmlObPWhJTclP7CbhB05VPiCxrM0hDn/r
qr7OhRRLuDIfkw+nwUc5hacs66a0Fiq++Hd0pYYYUyBJhnxfSIig45xrhGlxzHPM
rqHQH+koVIARSVbOchFFEUrXn1wJSIxrwLRd1XK2nPzl4UCu8PoQOqNY/Bi+nvb7
aO9WK0Lm5MHGhi08on4xMYN/GQO42YLevWsXgc/mgBtwhkv0kONyTg6PJKNHqVXM
Map2myufuSaTv8Zp6KA8f4TdO3P5t1h2Z6Alkhve1Vc1p3M1RJH7+K2HkUZk4KGO
9UxQ7Hfv/2iL14bE5rVQhvEnqjpw0f89tFNhi1r8GMkXrDCr8AClRDSKOAu8elaq
T7Oz/KzJUB4Luj818kV0IuJLH2z9W3amR32wX7frS+lpBKfFlbGfoc7qKCdhsv67
yE/GrnI39/p1ztdX7xCDFqt2VJ/ywPWxnkOo+ngYVw5HOM4OSv4Za4XH+pzf9faV
9oUqPQ9x/n8SHz9Pxp9xoNwb6gbWQNNz5KI/vCZZ1KM7z//mb5eksJRjGiYU4PCq
E2DfZb1myhs1+Tf9QZ3/2c02rECE/X9+p+Sw3uGzygRMYWtNZ9xpgtOzEA04YqyA
1FpqOh65Ch0btZUxH/R4uclEhq9QAez9O09gT2Ri8S/R1yELrs3Xf73jDYNDTuAm
QtaJ01HllaeUibzobxt6tvVQXxwPni5drJE236EejvNVBHK7ZklhtsUwEXmF/s3H
DYG62QtgcYeCONEr2Q4JO33pW+DgRDQZ5dX8KeFaESxqwSVZBVPUHOOe5y3qMfw+
ZNYeuHrK/fKE2VqU0RhYgyFH1EWbikcjIH66R2H+X8FU3JohhsdL35HxUu5kMG9R
uyuFB7Fv2u/I9XbCMGeUFALmJyaPAdPvGNgl2jm1z/VwSXjSc9XCKCntHPUgntJ7
dupsl0kAEI1xGRcKuvQiVYdsTlhgsCw4Q3W+VMbJ2OLb9vYyYJPsNZXoMf8urwcf
qIH3mON1k0cPV2ob6dNjCug6E/aooh5BBRnZCb3youEhdx7dO9ub1qU091kInsf3
iNKXxCREqSwW97Fch6lXUlH044QLc6GxK8hNeUt1zcKyuxlXLcIz0SM7J4pB3d1x
OAFiJRs31V63Osh/IprB9zik4wVfXh1/nZG43HV7hrchfKujrY/s8dvYxSBfwURR
BT45YB/IwdU8Mwgk/GqxDNcljLZlhxKf/L+9amNfiX+XkrhiQBDMRl8pffqOJpYd
qARlRfVZz8R9RxV5jMKk7E7aVYzqgpvKiz7tQZ44Tph3MMJh9vUgfl5IuiYlWCM4
+9I43WN5NUAQXE9P0XYp/nl2srDQMWnNtizj1lm7EdGAoMvL1C30+xdMC6kNW97T
BpwdebQT2QkVxNOQvJ+QlOeK4jE/iEOORYcLgC1/XgN3PjGkbtz3h3S7VDQh62Tn
MS0BPuD1JgctF8AV3xiYkC4S6uKryVgDXIn4P+cmvfua2DRsxkG/yle7tCbf23yd
2YSsxQoxmyQK2hYeI/xgIriykkAVb93hiPGVr+Tx2uJarcdwoox6eKOdjAfdPyMc
LBa8p2UK1eyXK7bsND9ZRFm+RZDV6XQa8IqXz9WMxKkD8uQ7pwvcgtEN5qxI/9+Y
zOS7zj0oeuFmOiQ3pp7DedpRL1MfmndMLLC7GrASiZr5dmZpislydjr4HlNnXyNN
WhK8U1xnMe8502vrtiTxwuwg7951zgQt1fJMIaN8uAkjFwtlQ4JpxbQ/04csKGMz
NnlmbqRM38SuGL5vk+dcGpIIMWpxFsFflM4f4T+TK9fwwtD9G12qaaWTACQyi5FR
/tbmAKmcZ/KLk8SfCYWbIkGoKnWP1BggN/ZobfmGtGWcmiL7scesRb2Q80o8Qkt7
irTiiFmVw0CyDmuqWwLutoE1G/QOOqajdjvsqjMTwQm4/dy/5+HV0+jqdKgX46R9
LVE92cib/VISm392VwhAfzaKQpK3G6cw7hTEGb+BZq5J3LiB1tYKfZOu14Vj57ik
6vmo6gCK/yAateLreSHcw+091ymXwTtTL6XBDQ3NRfuj5An3Pj8/KVsyq3M1rZiS
Fh+f67sJC6jVikrAiEjK6WhVTjDQ7D/VMCIPgPC0N0AtXcDn5G5VpviwnCfV7BQ4
MKqhcdtLVmlGhwiPUPtCBptzSxzGXo/Ojv5MW4dMv9waHRY2UzWibLI3lyWvOK0V
aV6vy/qoF0xeJH+7if3vKWm8Bu2iPw2PYV2DMK3SAWMC369vKFgCVMCONA5bOidB
Or/8/jjw2w6UHCFUwowV0o9lE21SnPdZWod7SGlNgGyxtNH9Ek1eF8+gi4IlDbD1
cTXj52fOsT/dbLHsEeKUy+48Zh7dnfZXql2k+g8skvZ8sx7f9cbaaCubHdcADYaX
R87TzIpTDNBA4k8esqQFhYnY/lqSCMI/8RvMfA8fHgQqt/xXw3jt9BaimelmmyZn
47m933sY6ShdD0fN/1CWjjbFLh3yZgR7XQ2sxATZbv0LNTnIZ63M/KSAfdTeuULf
wkD9ncBFmUVo7+Fe/6VVuPdXBH9CK1c28+V5dYeI8XjDa2AaQ/P8an378d4rQ8/M
VoN4M0M3UqcqLHpGKvRkpGUpH62uXHtCyVKehUaMQgAqaihfUHP+Namrza8yqDKT
UqJGHXRHaoz1BFseVGHb1vlezI1DTprfkhPIUTZbg3E/y4HZq6g0nA0qie5RsAQF
acEKF8+fW/nAUI8FEJhaqltJhnH7RDbJYgeignZINUae1ytGBomlkDuTWXs75khK
sCwglEC/3p8EKsJybFJpYZ7Q7W8CnTMJh6meH/802OYEr9CwGzO8OHLgnZkr8W08
/nXil9+yzzyJEdc0a37QsUALqsWGLl9Ijhyb87yBKjFfV8cvrolJXPytHgiEEBTa
KnVyhBZhq54ey3M8AdFm6j+NuSlux93kA8iTp/38523ovJtwaBg6AYJv3Fs4yIfs
1ESp6mIWCa3YUkj0JFSqn5ogPCl2pZRZcWFJ9eqRCxuW4v9+atdAo1lk3x7I05Y3
yNIAColBQrPafsNnfGPowe6z4KSFdFOamwb+vr5zlWajJeO7OE85qq4KMYfRVTEA
FKLWXpJwrdMytGp3DGeFF2kDc4tRijEfH+lzahBq0WotJxGy+psb1low6V1lZvkV
dC9R4658FsoajfHi0G2LkrpMP/0T8ZMCa4nyxjLZTiKs+nxng7v7AL1KW+td6o1i
oXKrld0QiED7QHqDgusPt9S3NhY3FdheUAqGkBOnkKX2KrCq4BMA6WgmcIk5qtT9
tNDL+fOGrpUR8z3qrnDl01acFgUEjAxwd1N7mXgCGYJeTiqhhLMT5ULNerV74WW5
ELZ4w5X21eJNcmcRCYgMSyRT3SbxKKjAAaKfnveXdlPBsupLaiSSDjEvokrAcVVK
T90Uh4La/4YeL40Tny6kbytEsASmKp3k/RmGzsRoupWJaenyde8MI1tkz20wx3jA
u+EEX18ikYIRYCwOLEh0PfxOv09SQKxBLpU7KKwB+eTQ2m+IzF8bJD5Rdn03lwEz
1TR7+i1HYyhHgEATwtWLejJDWWLB2poBCCaoQZrJ698pnxusqq8ev6Kt2v+B8rc5
P3AqvswgymDgo/XZn8cbWA1ckkU63FXCO2IqCS7nSXfWCCzvsmQmzi9Vi7eDi07X
GPk+jcpy+yqafykb9F38EURa8zKblPyh0hk0tr+YmC/gZDNUZaAYq/WwtY3THwsl
OIPnJdHXh+IeOgcI/lbp2i2w8XozClmlPBP3vXtPgTDpFbkxyHYh8IMzPIhM0jDB
N5p2W431r9TwYlmAlq5Jkmre3BijOJd0ngbg2ZkqschfAPfpExu/f9BntbIqheeU
LR915Gj0qzkNtYJcbiEitygGxXUK49+bXy+j2cnxAzlapLN0RHyi7DH1CQ5vIVgj
Q1nxO/yYTu39Lz9gFWSvxB3+uAGStMQjtZlm/sdq1cKxz+1B4sDP2Lt5uFqxZwL3
PusW01CHVXhrwqIQfBwKz+QF71s8a7Sl+Wr3hrv94YO5J6FaYDEDAhVGC5EHMvuQ
kllIpgS6Ir+/WgBMbLUbkghU11/EQLYNw26NdbOOVogNUGa/h6f8D+LZSI+Rq73z
GhQjssoaXSPP/A7OCUbZ+3qwx0Ls7UDuYoJNHy9Gjd1NY6VcGrR6O5ObiQ3ps97L
rZExo6b0ZrYa5pi7kWNppA8bgnk5iGr5mUzZ54D1wwB6zGlDOfMEkG0Fv8B9fp33
jtDDZKlJfoyVk+K7ks7s8SF8SLjYTBD1hRuLAxyPBpU6uz4mw3KkOyTc0Ho0i00D
HkN95+sbtZ+lUEcucSZPukF/GM2TYx1Rm5p4hzzSJv9ulyGaIZ6djQJ2/XXhp4TU
s8OqzrBgNeLTFGct49H99gu552YwAHJnSvZVvgoE4hrxvUDHqIWFne47e5WA4nVa
xoowReOT9b7Kli+nXA8gbVuCH9vpyUpFfWLhBRYWMy/7lX5EhK4eXCTxR/PR9/1j
PfS/Fn3O1RHH93igoroxCxWr7cd9BZtx3EBYX/mRaUSKczxrQsuAIPC5dwp0qmn4
2VtKLncaTgswNDY7FzsmQwbWDpYEIE07z8wSzIeNwT6BZk+HwxIvBtY3B55+1oUi
3XpAceXH9QaJBg6L/QkCrYy4QnXklHIyBJi5cfuorLTNfE740P7YD9g6GbffW1yI
lbf3fRKhwjfPgI038RyhJFaIujfa0L+wWza1pw/pO6mr/KizGqM6tM5UrvCWuF0V
7yVnHoHJx2XviZkdZJhPNXxAldnNxWizFwSQhrl+bJ5pGJBL9gxITEzGnV5M8DCe
F75+35vcNo7pNDE8UgHWyYeNcEXW5vb4wlHaey0mzXz3p7MEuh/bzpsg+b9nNJod
hrm09WCckZRMlI9EVSGaGlrwruIX5EkGJcdqvBt4argEGGemwIEUwBMI6YF+fCjR
eCI6il693eCyVN5OY9NKgecgxNjAEkKOYRyslQLaTHJjxn+1ELYep3ZIoe5xJfA/
Sm1d+s5RiTC/TvMTqO2UoiMWL9MtlHeHHm5orFSLmcMhzT/yogE+XNMD+r4T6uFF
k5VD5eMVPvH/SBWMyjMKlJqpA6aDusIFJW5ZXfpAoyU1JOIWvzSUs0wHsPDhsX/Y
9FoBBL+EQyYVZqz8P0HuX6r9qrF+ws7Pn9sORbw/g/z2C4AEEOkTsUT7vytJu7JD
cDpIJS7RiMfxyRfA1KebLHz7nj8ODA8Vk5jUTxdC+oYt7xMJDe+0rID0zh4fYQGV
+4U3GkdQuvv5IohCtPNdbogVQvbrKCsc1AFgGqdRNqDkJJFpCOhUgb4sIcTcm5Lh
FsZrlzrgjdayuOFnm6WcjFpZ4rIIuYSRi74+49spuvmFJ7bWV8xVHsIu9Nz7OHWN
DaKaAA/AR/h4nvfUDXgFkZ2LRfw3zbk0xZqiyD52HF4VUrbNsTNxu/lCJM2rjOEP
D4TKsspq9l99uaI/MfZ2dm3MUZyka8+E2pBIiyqOH5hToVP3p0miYuYQrFaK1F4U
heRCa+o5ZNv1z+oOulRfR91F++ZWHYdi5zt9kS4nB9HpsHQqJtibyR6/BlQeC+vD
SnyWMhYouMZZu0SEEvUds0tVDr4Ic3KekE3H3J4oHQciRVkXHJAcd4tGpkGTBYfX
mcHtVFDeagtQAYxgCTKi+sFce3aNLBuJ0JteBHicrUP1zJwftOTJpcFhaPkEWh4P
0aa4dYOLs7DxpK850RIxc5mcEGuj/PR61hmNKTPVmvmHcZ1SH/xit4DvhFcC428+
fyr8ayGUMxBE2MIVSjk1ntyqwAreaTl0j96nzp5bJC53V4BMk5rA0ov2UQnhpPT0
yTGlNhO8DNhFJWO7Dqkl27kuJxRcA/6Sgi1nLj/g/IUbNzDVQrIJ/QX0Tylx4SbQ
YaYPSxxI5cSBZ/6C+ylxqXfTNB6nygFXW4/5W2Fanbp0sgSYA4hqiWcJ406X1fpa
5ZHO/OoHJPo2uuVGeQBoGp0TcVhg/ZRKMTfe2nhra+b+/aWaYsPeXJJkRV/ETJ/Z
w0aXIbshb+MDRd1p/KcTVsyroCO5Zhw1jaoW2o7DRV0krTUyLqX5CEdea0oZ6u/I
w6PJYkfiOn5gO9cZMuTvwKs3ODg/lzZTLhlfzbTXqulPGW8+99Wfuy4L5uM94BVk
gZsf8UjfBysw8s61bxmYwL4rWd55R+g0DJRRLuzfH4h2cDxyONgiKzEpBVA5tJzb
ACP/3+xs+13YpT2zA7LcuoHfWRfDw1WMnNPauurqMdwFQkNg7B9qN9N06rnSNerG
AeJhI7DtuTAhpga8+tbxxz1IIhlnaU9T9RuuJOsEV5liHZNFYV5rfmy308Pjuyd+
8jjBBQRiI7tUVEew+CCWq/m7bfadPwwe7wSqpaKGkl6cUA0KAAdxraaDyC/Mq6di
2YsCf/F/M5yW77JTEwqbej9RXmsRymLM7WzyeqTDNiTrv9JCk7VONWeW2Vmynl+q
aRC07QLpOTTX6vkeh1yfauB3kpPyZO7x05GB7gSQEVMZI5Io9YVyUKgAxK+LDNKb
csU8LkfOSkZRI0mJ4e6U/Pd38FzYKllx2VVtVV2Sy6chxsb2LcrmNuTb71TOo+d4
xMRWEfwng/WXePrFh5JSkQPsp9m/HHT1PtYXoNRi0GWJHKVilY4+CmolH5+eqNPh
O33Kp9KBJY/AUs4nEdzKQrs4QA5QHKWkSq6VWSVmAquXN4L1PhVSOIBIXfZ2Uqwj
m9QvTk90WBtwokMeR0zZYtv5mhBN75K08Bo2O7JB9IjqQIO3zOTsk+IRzpCnqZlY
y/YfgJD0C9vh4vTzzN80lBivEyZcVZfOFZNI/H9hEXMYQN41qboqRBKXs5NMtqqr
B6+HP/DcmflzxmruSKKNyrcfaJsEfufWkYIGu33h9+C2+/4ANPSBfI/yT11tez5q
uvPR3csJVMtl/Oi/KwNuYJFXcQWXL8xzWFtkDvm8fZkoMJcYuzdgjeIiAsS4bVRN
yp59No9jx+g2AXthY1iks5Fruq+SmY7KsLDiKGZfS8KwNLjsqAdei+ocMORUvq8Z
K7IvXGC64es2aeW/UnmlzfYRcOnv5UeJMLwhLgyijzHs6YYJxq40oyOctg29GEc2
NHBJfIGlh4+dJS48DqZ8KM03CaeDxxDf9xVJzwwd6d5fnxhDyKCWZJz/nQ3J+2gi
EwM1UV0sCyE+K6iKX9KpYJA2NLcVDcizO2mVcKRvhE/T17AmaXFGi9J959kcnYYY
sAe697huhHX4Kyb1muvVsDzHDuUtkFJfXFMjpJ798peIzILXln0DlWDJbPeAr5GT
qwC7AdR7CXOJG3bt1B4UnINQ+Q9WOvpqM2VXFY4ro2zsmVHfbIG/GHJMudRVsy/h
p7xOUUvWdNskLluTH/ImOvHbLTwYGv5cNaS9OLAexe8Wnpuj9tjyi+kTZGL5cpcn
8MPsULCbHbkZvCji3RTyXNE4jH4112JRqshQ4l8Xoc93SDR9LnGAJNZhJnuI1UE7
9sjpNRiGOW0zlv5zoQVBnIQWv4AXzwFcEo/I4BHb8yGCSbmp+FfFyfAGpB4x8v3u
AzaVEeAHa+nudc0umlggGr1X0nqugePSIQomMHOJg1ymAe1uwDIDsgxGf7LYfDwN
kGSgKmnDVvEjvmMepcRsfNRDaNGAHcT/IY96T087sw6VRJYE5OGsRtEBxuPoRjW9
+ZECE42TPP7aqXgVDImQOCaM+XuiovEcJPutTjgZAP0/zPi9UgdsYnmzU2HLnKFg
gTdRDTBoxUZzxFQGqgdRjJGw3E3C4Sy6cqRjwlLXJ+aVRr0mzIPuukkOVz5OWTCv
QeXb+zGrv5425JxH7CXj9nWgkrfz90GBfNUJ8NsVB7/oUnzl0/JkVQss0F6sGYyo
xM/iLV56cE2xdw48H9Fs8ynqnLL0/QCego/0+fp2paAXqpu1Zd1GiFGpNl2/etyr
hlC1FIHRRouAX99/kvlmxs9meWzpqVxcI4oEa5P3Elae3xjNlnQmNuZC3Us9q4X+
6vET92icOTMhlX3HAqWkmCukeJqxK82mUywkHkrIyhrI1vgbWccQ9/PeWJ+Cgvi1
KrT3+Equ+QuC/59/JMW867cQsCMv9SlwMmcDMPmsUwccs8TNnSOaLHio+jwJrLgF
03GXGdokM1wyKf4U2QAvCJURT00rPVSpQB0iPq83/AnDVfA/fSUiloWxmIoZdaBY
hNBotiKZ8SXy0U8IE5O6hOkb3+j/Ju2Ijd1uvp+6zK0bhw6hTiQaq8B+GIkLdrN/
6HV/Tl5+ZzFzQr9hWCQFdB1/poJJ78tQ0pZuw9z2TvuFJqSWp+oxw8//uzRvAXq/
XSRd4aLe9mWy2JhbgE/UZv9e6buchDIl7rPUINSANn0J0BYMD2lytyMD0ZmcfHmr
FNNPIM/4a32JPHOhlm9Rfin0Z9mTLV6wr3oGblUjdBaV/Za7mLRzoEiHds56SEb6
OKAIhvJI3Icxnvc74vxU8f1IggfVLoASu3UQr/ymsj/05OvD1mOuM1zBeeLOvfv0
RNN3EcVANVHB4uNxOlul0h3VDXj9lUTApfupnJW/D+Pi6d6ka80IrZsWn2XHCzji
0JK221wDDsLhnKp0wjlAvgwjJ1cmpy7XSFmK7PdRy8TSUK8aucWOZcdyOOhSysxj
XNXnfBu7Y2Fcd20ndNxBn1Zb8j0/04+NS0LHd87qeC8Z/CM/R5Y5yyHooM5Be8y8
1+4WqlQfvvCBdzsS6pn1vsALrL/+06BrivX3McJ90oqIVIP6AVFVykTXV+xtjUUE
PxJa0Ke7+gySLeEAg0LyX50nGG18uUXHoi1EyuAeVqYXxs4pxmewM8bmbMKX1QYI
tJga6FJcZqROez0dhBN/CrKwU7uFMSbftbv9mvUmgLKf/6GPIXVZLYAX3HD5Bhly
XhQB4EjbSlS1LkC6s96QZSfb46sbjbEA3kgDftt/hU7ZUCSiGpK9N1Qwzn/UA3LU
14YK/fEh4p1WQLPZ/UkHc0oS79njFZ4vG/PTDDFBrUPnQWvLBLA32MnB7hHzoxoo
zQ8jnaC/UMU21wHhyw9IzZissYLi4p/020wkjc4Myc9A4w/2wrUyh90IObBBZJUk
ujwtNt8EcmLP4LA2TENp8Ufvy8d/BRzwppxeXkmfneRYRHe7GMRqkq/PxNioDldW
RAkf+QnPX9fwZ2bn7LuxdVMdkr4tMSkkGd2apo09mWbGZNoYVpo0SlfhmbFd633X
0dy5vC+lcTEO2xVG0UqAjFi6cxMgEsPV5Os+yWDU0Aljx7V2/spo+6qEnEuwqprD
DQ1BnZ5Dxs3J4DepvvcfskMlQqmLzMO3B9y9QGhc3aDMe7yPyLiMG7MJJdmrsveI
20xdMTLF7zI6echtaEt+A9fhmr5JYNiPRy1CzXwrM4cgxf1XxYZCgLLIYGpxzYNM
9MDCrkdEDVD7l+lEl7h+HvtIiZONqTYNNQ6CbjCWyyRJIB5nhsVLDtB8pvbxTfla
d9PsPT06BDsKdDiBwAcysAngwwrzgcXQ0yclf7X5l6DwJeEXBt4scvqsqRR6Ztol
EK1PcGV3o5hto0a5OZ3POtqvnHztk7FSHLFUJ9eEiy7RDkkwn19q8ieQhYAuKpuA
w7tK7FboRqZANmQnPtYtXK4Ae1VKoc8SvIUDASm+Qi+KYnjv908Hxnk2WZ3P6djU
9Jmzbnzr1/WQDCu+e+WfO+270UEv54I+MFNtM1FOa+hX04SoUrhqJ6IW+JB+I4hM
qgx4JUuyfkXXQTkknNSwCkkJdO+Cu58hd2NxDqO13QGlT5Ezf/aDWg/EtC+szFmG
GwK0II8weM63/i9OjtwdG/fzUq8ZY9HXQ8Oz0eRGzhguN455M7+AdJGbakyUulF+
CdQDP0qJutuV5o63vUPr2u4bHjdjldTm5eO8f0O/Wbx51Tyw+2BcxG4JWm/RmCLZ
MH1rPChqQEdp7axtGPlHB7/rMxBKF18pHScqdhC9dqLtzkvYGrtbH+vUYtSO7cYC
7oDs3eWrixu0uLKpCoLPRklDMGAtYzohwxOdYSjQZjiRj/jeTlWcLSmR6P7KLgoJ
1QSg91zLNNcFP7KNN1eyOLoMPjct4R+wlm7QdS951t9IFwrZhH4o1JLO51rkTBnA
Z0Y/vwDTPIFimu8jv0Vnl6J6rHXy9efAylVCh/OVOBbuK0XF48nuXxixw+voBnqr
jiMueVkyaSXYAVWuD95B+iKdARHs97Xyhf5ODIgqT6n0MR8NK7fdOgmOOcszccLE
RUsKd5+R8LBniy0DPFtzsRjhOEe81eb2iXCX/pzqSodsNneH5Lv2HP6kDI49GpRd
a+BJijos81cSgBC4UwdOmxoXMojIrwc7JlZK1WuKxUZsET5mU4+6KL0RaoDuAITi
TsgMo7FZyj43f3UilDWTMceUar3r8BHNwr2eSvHFgJ7MjkzRnFeXXoVsewxP3VE5
UshtJ4Y6LJCfsZ1s0Zw5JnmR3j+8LyKzQCfZ6ZRSdzWHya4byF1QEqUw5FaEF/dr
Kydvwj8MrFugamx8kwGKyqMLCe6FSvzZZMtRx1F4nNIk/fB6Qq3dRdkjK/VSyB5v
lztndllggWe0H3v67kWmbe7UuGusR8QWqfYu83hvMYjQL8J/U1MKDBmIJjVnBQC7
pzYab/rrFsAMwszogk7B6Diu8axteM1dwHaW+DYE6epC51xJk0bRNR+BwMRB/rid
PRItYE7B/wJQmM3nsUO8Kd91wDQDxfa9WNp3aZzIkWuaFKCSVMMlOcA/AabWqg1k
QtT1gdVCpoqiX6AUQGbpheD+uFGVpVLhvtvjYPg0C1CyYpGJcdJBNUvrtZa5qKWn
C7AdX6vbqn77QyfGy7/yzI75lX7eZKZJbUFqV6m5wwOE7d9uUye2guEKj8wcM1YA
G2O6kTj07dsKkRrt/xwWfFpL4rpUsZOG/+88RmiMVpxVgZ4Aspi543KPZphm34gG
dy/4yTLNf+tbuBmF0SNZA4iwVxqZGD3oKXQlgTYPQ5+VlGPBQi5M+S93SVmtdBs4
qjtSXVJa2VpVYKyaDPB6ZPma1jPiC3ZQePRfP6oFJbz9YE/YNQDSoMlYfgsUSMwP
8atZOFR+LjSZu1iwoNQmLZS//fO/B+xpCiy7gcaIJWMpO3I2n8h1cwTxK7z50yGC
gIlzqurgVgRns/OBoio5z8/CjxBYjzdFroIpMhLOsuh8j6JXRDNSsoVWFRIM166g
HUqdHP7DWSc4Vl36TPBZi3XSP9exNJE7D/RPhXcyksrb6TDqzc3qQv1X+6GaVoul
BfCHXeR4BMU7XomB7J343mFifDJTLVCwTeEQFSvXMqITLsrsGdS2CipZ1bBllTkL
n6k1U8NjShhk45h0XOnUyZWjo2T8BZWbwwhBn9L6kH0LajoLBNoSNcKigRZ16eqA
bqutDeWDU7vQbjZ7oYe2Hbd3mJH7aLzMd5NtjczPR8xomq1rvLBJ8LWe3XsWZWau
2SCZdrvR6EKefRmhB3Ry0v408HHfKiNWni1ugviW2PBxA2epgbAsNst8IhX+ua5H
9pn9gMfQmbUTPi+GVQOfRIDepYUUDsboBNJuP1C7yOaQ17HYehVuZ/5jjCXguy+n
GIr+Ap1n7Eunodj+RBHb5HwuLPSp2/97BmpytW8WTMG/lxmXAwEnGcTMS/0zUKyo
a/1B/5otfU3DNkMNlyMp729T7JNE/D7ltAkEOR8d2osBtGVZjorTLidlqpZeHXq/
eZgnambSRQ++uG60sac8c2nYuaboRU6eDy/k4XpAiJtgVrOwR2r8MsndYrFiIOIC
BjiTAMgDJaVAzDo4Akewrozx2J3yy4oX2laH0AjSh8BE1mWRmlARGmIPzihXc45U
3ApJn9/OKtgAzeO+kEbfIqd20UfmIq8CuqJ0Tl4W4unypKFPX6vT4WRgVS+cG+Zb
MCI7MwOqFBvAO5W1I5nVidReZE3rp9BeFLqJw4xwMwRJwPA1HG7eij/hNQriXGgt
I34N6p1PRXrFPVdZaQgBr70Z9CJQPMeAm8gSL5xqLxKGV4Qv4aLIQ1UY5DuumgkU
BZhOzMeKmHKRQ8OMq2R63Mny2G0JYPkpU5FMiQkPB558CLg2pvi3GGAyNMQ1KHi9
CkvWE15Xvd2iZzxrRKgCe85tp/CcYUf4Hv/ltbnGqxact7jMYxj6/9PUbseD6yfE
l7sp7TqYsAQ9INYSpGZ0WWYCuwqrj76hFT6tUNCDnY0I05VS9ZLED5XKJxPlscGo
0waHnwvXTKgS5tN8TAM2AQvF/70YqkG0VxVAR/8wyaWc7KO4U1wuGxH4wDwxG6QF
eqY6/BC+2iQT9mA+uEas/WKU391Erp+xaxC8yUtnY9NkGRN18lxyA4veKt7aRcon
H8vzrs55I1tpSPAvjthZKo+4YSSx1U/ZzOMrsOB0vxFJ2RVElueC84z50Kt/uMBG
DqL9ODDjBfaHrA6h/KK/dCQtyrayd0EVyNZ/gYdMbZg8hN9nm2YOQcJDXZ8aKbtv
8wJ821uB3PQWDll5WhI98AaskhJCQ9oeEZfZTW8B6OcAe258CQSA35LMkYvAC+aT
wR+aYSzh7ow7kqoQDW8C0xUjuBTq7QoCJ+Dl/pjTe8YYtdy5EycrFExTwJmLwBxW
552S2fLy6vNAa/SiaMcQiWvIu5TJd9Hs/asUsoM1FiG1RH//TyBSC2AeHnyzb91n
kh3V/U4K7DKE0iFepS3/6UfwYOv+CD1L6mwsUi9Ea67dCKv6ZLdZDlC23ETu0wLM
XwAgkFOxndCdEpPBVsYJxGnnbPpFgQExjJ72W5Hd1DBQuoCl7NWACOaSMlSQisoq
yuA2yjVMv2LGtx83sCG18ybjTDUkPZ80vZ3jCLR4mr8U7XtUAU/h7+pfZkIQY5UJ
8sbCR6uW3Hq7R6oPN4/ArSfzOIxX2GyD5EGt3bifpPHGBagit6Z4/MOqSW8RA2Ei
rd/3ZDde501sXevg2Rd9qWsP9h+XMY8NVI5652Zh7QJgEWp4STGfA/YR1HOc7dxI
qDAW+50opTGykj9S5NRNXxDLM4twgN+RrbTudJdy3zmxCpZfH8d0QZATTUO3kxqX
dnj3uQ2CoZrto2DyCtbwPgIIb2Z1Qm+WnbbQn5Va1BV34XKBx38IwIiAHnCZKzwt
4waAEIGeTmRKN+I+X4rDwR/APF+uoPkJZRRIb35eIs+KAisSBJ/mdmSj1oBhWb2n
4zo5PnCl7d6LD4JAksBxtwqYiDpYhyD86pby45Ecjs6L0MZQHE3InYg9kzQ/ahSS
LtA37/HQmiLRRQRpNBueBkrHCbtLsaE+kFZbxwvqtB1Tqm/WGxAK09RWftsaIoxa
IL740QT52hwJUNssWkQxJYtEHyVIJN9RsbAgLavsXLnbfmo32skkXPBkux0qmz71
Mzdn+MGYG3LWSoettuwR6/bqh6nidtI48CwbLAZba2o8RpbjH6ELoXlelfJHynIm
dKyENq5T6kT8f4rHJIFio/ezCHsF/6VkTQelB8oORjdQ+tucfPoQwdJyZAL4rgXi
dFsagGgfHSLm4gXD156M8TyKzdBL57ILhDXdMdl5JhF7f0WRnnPEgDcv2Qt3gxVS
1wjEvpGzPIgpNge2qvaIuJC1ltMNDO/U71ORW7UMTFJOu04402OkJKs/xh2HV0qk
aJXXHbvcnuvLlWdl3utGlV7fNdKehplfvz6Urog57NljjEDJBducX+V1J/34YqRw
uP5evGoinC5AcOWDfVHWTgvKh1Dt9QrqNhXJnQylP6Z7xoDpsRD0NNgQ7CuHR7K/
CvwWBT7KVXPS9oso6Efga1HMD7Bl/eNhPQoN15g3r/dRXl3l5bKP208/QBVO+Fje
R3QYSVX2ZFx3KCZNF9w5XWtV9BHfpHXglvoAB7v/1pXx3xoCeXgOBe6o9nehrA0Z
I9ZhUPtWjk0XD8CleUeh3wJG+gwA0B9hs1e8TKBDxD6zAl6nc3luU8tGXeDT441d
L1jR097ywWWeTFlaeEB/M3ZanZdgefJOV/WjA8VbsKnn49sHVA+aejSgJYpMWJUZ
QdoEZNThveQYpULFUucSBquUgVDg/cg7wXrVQ58jDwAavos4i5vzDEUT3msn31Ee
Sk89U7M6yV+kQy7egnDFvccmYTBXJdkdMxlW4LJX1+t+zXC/Uega/iga4hyjUXzL
sGXaTUqKkRws31+pqL0Knm74R4a1cAh4QxsN+PX6MHOb0nhKwkiyKJEtpiMb68fS
6t9QoeNKVRB3AvvgqqBTyl5RK0ZABptoog16A1QLp2pZZjkWYR6wIM/ka3vMHRlq
Zp/x8AofDfwNPXLhNxrVXcbK9igtf+HpkI0jJ0uehdQxxtNwmsA4Q6T1LKyMYWC5
FrmNIwiEuy46NVgTa1cG+VtVChUI3hrFWrfDV9eUv4X6MiazWqlmWmTz0/ZLXZ5J
F5gFLLLidjFDMSQGToEmpPCRilHwiHy0oRR67f+5wirfKVL8Gy+84VMMHlZoG3G+
Jc3wxo1bDlmIqABZmmW/w25AYrV1QJgedeY5zR3UuZFXhsr7ac9ArP0siEDk2bhi
XfGhn4uduY08RGXJxBMGfifi5NZjY7FCAlPkggIe3Tk0C/bT5GAp5wdSMQSnsXkO
2HUaf2n+10ZCee+FGoyrmEh45Tz5zLnVA12HZMrDOBg3RxHboXU0CFNffRGEVZbE
OTCv6l8MzBdkHnjfN7LCMQwBtdak3r2zC1hiSsSOS/JEZISSJKCseT7wQRQTof4C
+e32PcPDbn1/vF+jhy7aziOhHHBzHrfuz/2Nke8hhCSwRtycFy2m13qbTGLzRWRy
G/QDHaXwSOqRQLnd6h43WIgIr5u3wibe0cphIrBhly/+dhz/Ezly+0XXOY4+deyB
Ihn7/iwyJ5DglH7WW814DzLRLaLORGm8aHs/wL/92WWKhNPlZjTKkoByMxPyWfqF
PZltfCDoWKBUMEEVmI9uwE/AeZd8cfnqekF1bhyTJOGosVzDwAxNxRxFxiuDiJRP
n32QkQ6lO+9ff0tjN3hJi/NrGF6zezRqOWp93gZjCid2ZpO6flPZxlEbYlaq/bs1
GldACyUANv/BaBsXgnjRwcIotImIYLGjEkkADFI1jncBzBYrqYM2Eb09Amhb5EU1
2bs+VA5dxY6vEaph5Ojz+VGOn6ZsSYVjPAhhRCDtVe12fU5YcovIQCSapC3QbU0v
z4NiBeYLk6jpMaKgX1OuVK2OQkmxgj2qOTHX4JcmAL1zMO7KfJYwVL3Qv5G94swP
ay4WA2SoJp63S8FkZmg2X7D4MSV/94JhHspZEnloKj8rQBECKPf/vNPjx9ImRi1k
opWP6e9tlILxCbyLAT9t35Cf5FjG3zhvYRtgx3zr0zhIc9yhUT5obccBQ0YwR0N0
IjQ06xMb6MYLd99us4INMXtSJpVqpKKk7w53demDpGnbyAmOLWCKcY8/SmK+Xkof
pO4O+U2hn2TNPXfYnbWTB+LKTEUWAsSz76qytrxYTAv3kOm+fDXzGDcpfyZi24xV
1TC7iGt3/N3kTu+v+Cg4L36MzzI3hfR2ZbBqnhx7ePPI/vExd0wMvCwklVzB1BU4
pzPbzDYX7BVoyN/omNzf3YNQVtaI45gpKNpmgjJMbLXS6deYFxbzopSm2olZmmY6
eH23OOmXLr7QlZzym3bRZrDsAXZDSHwwrsB4Wp+ew4AS9OPg67Wb6pXhrppsNEjc
VM15cRZQg6SaRNVp/NStaM/WXChNDEsQHQJt36Q9t2afLAVioLsu+X/6JJbswocV
KmNzFqTuVRE1CR+8umEBf5h93z0grG9k+4l5KmPyCkTBuILB9yW91KnI5c7xclGB
r8r2T2Vz/0AqMa7Jw3V83cqkqB0kv7MwRkTn8fPMKyoUZZ0ekklT0R7ylnC8kW6u
eSTDtx8rNcHe/srTLBy3X7SVmDq0zr0IpGiMpe5Lx6N66MpJ2gPGWgEHyRy3WiHM
zGiwSk962K3pj7PN5z423N1qzPRjH8vo4Fp8inEdkwKXphWDfPTRGsISNHW5OHeQ
oJgfKjMHpokowVN2etKnvELOZMEZAZpMJ2ZtbW7XCDCW6BPJ+JAmnHO/EBnfcwpi
ihZsDuvtIOqV/KXldbB0+hFmxgPK5RT2fIVUERjHuyz4TGrH7o+5ufV+XmNi57bo
jd6Po8HZSD02poyK8S3qCbR6zBFkX2blP9blRB1CqZPLvqko4biGdIzGUJT1tv6g
Mv5PRA67JMXPo7DNTt0yjBxsEFNVg604UU3x8ayx4MjU6aO9YlDasVFXhE/JpCsZ
RbJr0DlokNIhT2Cz/EpoLfqf8qQ7gT+HU0cZKHPnsomfqMk9pLii66f6AoXrSCXB
14sEF8zDQYRoQw3TzCMOOYeWRfMcBUE2rY0lkKdoUx3lJX3b2z/X1NbDyzk3oq/x
pGNO4uV8AfNnSi4pXkX3ynYHtoOlkE53Py/1hN4KT3VlWazdZjd4uknwMLd0jwgz
Eon9CkrAvKQcxyVfu7TCKo0VG85ArdZpQMrBng8+pGqy2+Com6AgweAxNV+WpTfT
ZiImf/9k/5U6VdxIVc2AIRYtIt+ufp9GjSCKITe5sv4HZVLPJFgbu/F4nSiLkVpG
/zewYmzh+6VulDj36HT+Vs8XTwHFsIwENK04iT/Ova2RrXHwN7klTmcEFtsPfRbq
2aSWG8e+BSCBfGFRSiUHI28+EcGefJPWGvHRZVc9fRHj5U9ikuuj0jxwgVJoHGAr
O27cF3a2jtcs6nVVgzRSpo4UxoO1H2Jt085AOER9O2ZGcPejGFxvDyD5guo2THCa
eW7z4xxqgebdarrBSy4vPhE0OzJwEkHOTC3EpRG0hyoYdkT73fqzLerKacY1NVjc
dyl++RN/XA3BT36Ypt5GMB1XHSyUxC3+vmB5NTaw3OCzTrX+KhwNRQOdC8yqnKyZ
XBLLoMjrhzq2x8z4iYYvaCXLZhj29O5H1xJFhQJxVsRCjBrvYyqix8ZE7dGTeobz
9FJiHntuUa8VhWbQp2BPEfXgpJozDO6o1znnS2Uf0Oei2CNTp/nM38m7l3PvyV8p
MwMQ6lWyXrgp8Daxz1QF37IqoTMcnTjaf3qXpUtA0z1Dy0Z7T/TrWOnaC/8s7yYZ
56fjAUUfA9mh557u/VFVxlFFSePFNLQ08YRoO6WOU7Fk0MIIPyCPZ5JM76pFzZMY
ex2BgIDedszucNRbcXUGgl8nsmkodR+t88ddyovgl0K60GO7aSOgeYZvKUu9wQrj
Uwl97JurUeKE5iwAau2zrQj8uLMK/8MzY2MtMOlTOIYtedzS839eFICHY5Ld9nMT
cOVFGgZrxpXVQS5GfushRvKm1nkiY5ce3dZ3SWT/djYh0n83bFMiVQ4I173W4CIR
WkwiAnMWBeNGXA9wgsRUkNL1GP+ZvhidiKMCoJ+uPdqTJ9i3pQbNMxeqqyJnUgJh
vl7qpQ+m10Yi/GBqJImiwJjbM+lHhhj/+e/KdaIQCf5vp6bx0RIuo04iKIRss/Si
XfiTJ7GNi6U0WErvsUIiDpKCO69/ttqORqqGVCeLvJZiamrfP+D7hYTtxd9DV7N8
FmlZCIaavVkHd3WKO2szrEuXMROGAJnywWbMw1e4z1MuyeM6uiRYQiAhmYyLX5fW
wQFwTHCmGVoM9h6xUpcTwX+es1d6SBVD2a5Y6vwcj/811X1O7C7hikh1Vt+y9K19
sV+JwFsRnyqM2Gff3C0Ha6oAYO09/xorugdZBhZ0sWdht4OpWCYGVl/g9g/vmhII
WTkMlzoua65F3ON6t4I6AiVO82KDrlx8BoMSPezLW+Maddx+zGeNyeq+uKoLHZsa
W+McX5FK2L3Q2mv0D2vKQ4d3ccKIhKkd8ff/VMMBwQzydCYSG+lc31pmVqdlBNf9
HpDIvoNmLGjJdPF6B23oKNgh+CwrnLOWySSfecI0aaDVH7wW+Q+XTBhzqhNmGl0p
Rd/II1Lj5rVk52Xbp3gPMz4JSOiqcjIflYInuauF4xD1WzcRjO2QNEscbd6NNE3K
fwPgd3yTJ4DiaA38oQhebhUyufm3z38p9/XpKfx/Aam7Z01zbAhwpfz6o0E/o1TO
ihTdcRlPjStuOvvxMCJTzil/0rqTFEtiCCblW8Lo9eVZPTZaCYlzWUrW2+sNFIiE
6pNpmsV5pNx0y47XBKlazSent1IbIqrfeZv5+6DNkh1m9EuiiSG0YF49BUYrQE7Z
jfSqSnXPXUvwNsPwacaEdSOfK8YPr/7yCqkQKuiuzP7FU2a6We6qQ5+O0gZPd2ny
3NkMTdCDhvK6moI45CkQOOj2OXZPUpCiuABTEjGsULgjU7HTau6ATocbgX2gwbYi
QExNl32aE8w0Q0eQVbLzpW+Q9UB/1TCMaWYoH7sXnd87PN1yWiSAMWI9IiwxLlR3
13rk4laqzWd5ABbYxf7mjjd7dNvp5qlsjrMexdsu0oO2e+RGuWK+Py6g5FCbSjPz
D7m9vXvUKkBCabm4c/q8b0y0yp+LBzTzjIjt45cp2jek+OnNhD401a5YYJuC19E/
pNpoUHjukiHqWpspC94oNftpDeH1oT3wVw2QR7vRueCgIOTxRHMQ9uT6FW9AU1Fg
6ZLSeIS2kCb/ccayLmRnXHPqi+TXZc7cQ5Dg8WCgD0SM7H1u4d1QVtlTN4hIROCh
UkYr3ZBzYO9qT1z+uIjuGQOEX4Tr1QjxovYTBcZ2Tpu7wa4GRHEQZDE+NiXWZzGB
pJguz86eEHzGUMG8A4gaidtP/SxARZVH8RclXbE1CKzRIYG7jkPzFpjsXS+kbuxX
RZX8R9De49LklQ0VUAU05F7/IXPs0Dpe8qKVSYySPa6xZW9FJwt6pGCv6Zh4XAB7
8GipVDoYoYAJ65y5GvXz6pehdxZW5/icPgepUezFTtvHNyCoKlOAp9OvLwsHKOu8
bLvq69Jdx4tXZR3UfHyU7q4/ZShGqMB37I1wtOGoA9M+BN2ILAA4dAQ4+sjfNOe5
sGosyFDBJ3TgZStEsmSjn4iE1fIQhjMnbkWMleMx0WpLlSjQ6FWzAjVae2Jwc2H4
BbzgHO3H709OFHPB+d+el8bXYvwHIn/B9xD0akYvS8N6XPOLAPuKZ9ufQj/wq2B7
RxwsMvguNuWUu45kQbxGeqoJcL4QUlelB47KY5Erj3U8hrSPV7wYgWCMwsvWAY1Y
fwS2ohiU4sR1WKx74Tq2kBV9A0TlOpv1L6j9+Ic399WvEStspXG5ZJyJOeytAxDQ
9V2bGAHHoOp1ChJrLsqYLxlc21mvZhiaH7qdJL5gZuYCabxQKUG1fgVhVUCB+Pc+
doLNvAUFwiS2+bCqwWkCSsbk7qJOmqnB8sfe978ukGq9kaxMRIeUNkol/4rfGyvI
dAJ0SxNBUU5owy97jEcM47PRLMRTWaZ5LUvAJK6Uk9aHyJDwKIxfSbgQP5IR3zBv
D/g5fnV08Ph4OFjFyMBkLVgCb+BK/7FgQ1872HH+kq7aHcgfjHg4IqiF7g5NDHI+
XmYzn6C98rfy6fz7VJzJvNSyF0aljQ0Yo9uFDM7Lmh16W6huKGr1sPEH2kmknwbd
iokrVhNU0mFDavMow3NnQEdL0myoMtEYd1IQ92JOAphfQzlhzo6NJ41dma6VHGaN
CN1n6Jb1iAXXszsUup6/K3hI/AyrKQdDz17wC+gf61O+5FeV3NKz637fLnSrrArr
HnxyH5Px7gn9bXKp7KcZw9fwcpdGW5B2dL0tYFgPkSwZtLCe4NmbZNFwJzSCZnEL
OMkqsYI+u4mJ5H52s53xrUnqJ3JXoN/vxuGfSy3iGUcwpEevzqIQlJ+dS0hsYU6o
2JO5E/5896fkCGxMQoTI81GAAV+5lsuiCrMmiJOALTodO+uglVFpRFq/q7YIe7nY
IUyHSwKv+hiMXasTPsJgbmH3Sk8FDtSCA5+2iP/lccOMSdp7sShARvsihMd/OO/Y
Bcj3Be4SMu76WbJgxh+k/l3MDut/vuMHiDohVbczCn26BdSraTgwTOBPt0iS6wUs
zuFA28ynL+g5HqbNCJ/i5Y5wTtbIbFef2M5+qeje2+XkpGaqqWO+Iki88x42LsRm
I4NOCWeDtwzgIQBU7Pl1Z1zeZdRdIIgD3UnTKTybEtGvujmqWxEXVgrDOg344gaQ
fMGhNBCbO7XmjbFIzCzOtfbV0OnAaaEJAY/7zbACUcbcz2RXOzCC5P3ZJ801JcPD
KtfmYNOdamHff4o9kFkU747wGIsAoOk+7nu21goOnphBAaUE2CZIpnm5YdAXkfHU
rzDRL2FHmwAPfZvekuxBSdr5jp0i7GNt/6e5jqYkUejDFoQISKIlX7516qdEJWqF
QR9ItDKtCg6V0MJdhZxOTbOhKXTdmCmkx3jZuWjRb677q8Ls6GmjTLIQinSvKge6
nHv9UFaGwZe0OnhpSet1sJnr35B/CNUOfMUz/WS9YIHqXGQPEyQ3mDo0uVSqBCkE
orK6TI84bGr948pFrQuIciG22DZ9wVs0kcHUBIsxNOHmtAsLptmu1QkBQVEx7lPM
Kgfz9kpH6NYVtA7DYRufvFUgSMurdn/YspauQco9c+sS+4GVl8HG487xsVfnChFU
8SVldvVopXJPg4+pj2qaGkgOnFh1rLGgavXBsINPcVTUTCjHT+RVZNElA7Ruw2sB
BuStJOM9uWUFZ5QsmtF1nrOTG8Jc2NojPGce7QkqP0e8+yi+hqGLXnjcbqLZe2o2
fJEsFOblrz3HT+5/x5lH3NlGZTrk9pDtpfWAHP5KJMQCzjdCdVTIQuRS8L0VHFtg
idS72xIPn7qW+oF51Y3LPck6vEQSq4kz6FBYDiDV/WOJ+GRmLwIEzXwrMLAICBuj
80WUACVYKm8+QhDjrTpuci97074HnEOU1xpsnY/NhQOaImOpL98MY3G98tgKqGHw
eU5mgcdmXtdDAsjtj3ZXSjoIYH+Y0hjCMT4tXC4muF35aYuCbsjVGiuydXUWHEOa
kMiFw6t1Y7+8p6pE8Uj0mB/9WiJIix4Yu2gOQoDEmKnh2lXNo4LFOdTyd+l0COe5
xTB7ybChGBguEbxoz1Xmrnk9mCssySpJZM8Qlz82wl20dAhZOs49cq/rcVLPfBsk
HZ/zrqrhQC067HU73NbU65OzRagUYrYlSTnGv7qwDXHZA5Xc7eBu1KIUmDKEg9kJ
/mIKAhl08TrxpZXZa4rYqxY7EP4Xaiv7fHOPKEL5GeZk6bgoYRLY79Rc0Xw8pwZg
qbSy9gsYDehpTd5dAvYEk5R9iDtH2SrZE9+5NuTyr1U7Ex5VHTw2OjhTIK7fBkoi
nLu02TZV2Fk3zHEKUHvHZSpPWkcYEkC7PDEEOnnPBguolJzmucz7+ifaxj0iWO4h
VXhwZIp+KmtcvC8J0A24xFsEPvi5ShsO3wHlodgc9IuYobFDb2CeEwICBx0NEj9U
4WSYd9OZIkOqio9CZlQ4e4hYBQAmg7bbJgG2MqkWJG1vfPrzWiXakYqydGPK+yv8
vuSQB3CMj62Ujf18vOHZBm2dIaEcNSz7I+MJXNwH7lpzgQwOcq1xecslvG2TPCpH
ouoCEnOzmCy9N3/rlZTKw23m2W9B/XTgauY0tkqljImc20J0/KXpg/lNKWzYsz1x
okJy9MN7Et9e86LfJWhPoqqdtjuksYiqzNCWO9IXmFxmP0GxMxjF48nNg/Ox7Lvr
hJyWgKtQnqLH6w2LFnfWOkIu+Dgvt8ylPxvLnycc4K4NBGg5Vu8YECoocCn6ETcl
F5npG8jJaOP9TJmhVQJDHq5LIIh2/lS9IKDRSr4g1G7kFEsCjUF9lgKJC6y3GQy0
J5fMTXxUhj3p734xg2ivZcw+7FHN/NyJ7QTH2VlSpwbczwTfwMzOmpL3yRvlQ14b
O7bVKOsd4OgHBTTjLQaTXlPiGvpez2uOEA0A+DAackX4oPuqbCm2zh4ZLFAz3IZi
RCioqsW+3hijjLGwsHhlPSs+SWwtU66Lg2fKh8lGqS/UyGEs4BmfN26p7BhAzUeC
okyDLEpABkML7jlawuYpbOxcxn9OrccUEIwz4KWSAOyf1dTDXwsn3dh4zy4amYbW
dONhHxMUwuNz9uCzSWjOgHIQkJEcaG4VL+VO7W+jpqgkv86OW2N9XapowjpfMPwJ
D1GVDzpwb4VG/dcjzoFHb/kgRSSYB6A/xOk7JnaiozFBWpMG9HUdjG1Qb+FIvpz+
uv8LXQEikBRjxLPtZX5yr8yDykIvqdsxDwt1j+Zf375M3kTb9Esh+x5c8jKrRMI4
X6utP1Zj24poTHoM42Wo27zeF91vWIs1nQlpr9hUA1OaaTwC5MsoI7sfn2rk8KdQ
AsJcxPZgS0wihggARtSoao3HkyVSe/N51+wbUyFVxKKjZLJyoPkDyRsRRqoeplrD
EhXLuD2uAu2mhXBcq7/JmTQMe5sTP6EfhifGg+GH1ZBuymNdJCoFfGFQnXDZclCe
JPghHipHCUjv6hM/wcDfuxrZn9YXIewwbsVCEfujGvouP7ulAZ58nrv0vKsA3Lq0
l0f5s0HGUBXCH608DlxbHVnTq6CmOl3qZXxyF/oJxKJFshjyM0oPxl06PUduh/4p
6HGQL7epkKCHG6igA3cfmV1A/gcs9FDVrUCngRqlRdfrW07NMlOjS/6LEhbOJccx
ppaFICGyOyesOUcLKmJiavPWz7kbmg8T02tcV2cfT7RX35Th56eqzhrLln0dDTdV
ZUfyaVAIsGUHbSiIAJN8t1Q8pkyircxlLlApDAuTiXjzMEOcm2RZPD2mNvAGyB3T
eaZDiRAFeCvrcpKa1ViSZFtAGjpwJmFwDEpdNJn8FgLTM1pLk7Vdz+oecaA8p4t+
NPg3ED95ffPt5ooFuHw3M4B4/pSib7Ejk2oN0jNENTD0QyKYzDzt8PHagdSOmrgq
JEVOLFhfJL30JvM6N9iz0dwggdVMD5XUQKK6oXspQx1xT/A8pa0AWtn1hnVRW2sG
fBO8Zqjp9mjo2lq5ntzF9TNK715XOwRIqWC+G/n8/DE+GQNahA7gC/K8hU09ma84
C52MR739U/joEdYpgt/xH8sefGA3UUPYna7Vy8jFsBW9GGFfHxu5ZJmemAFL5Zm8
aTuQ91A5l0z9z0Kl6+MhRnaGqbKxAyuXr/LyGlZ0waO+VVHxpCZDTN3QMkrkHBvZ
g5ZN3iO3TrmmCCrj4X4leTOwKNwR/4Hz41dleHx/Itj4OsdiWWf5Ranp+NGfGmRz
bCtagyNEArL+kqqKW75RAct8PMd0lX7PFgBIconkHFFNdcu0Gs9rTTH9ne7hC8Rf
RAZxP8uxcqV6IAiCYiUmiXSGHc7Aj4yx5x61ETrk/AqZgwFbTZ8Qryrt16gvf5vZ
/MZ4wFD/1OoplFnv+DG9r3jkWaOFkGQTm8cM1iiyAnsKU2acnXT7HY/FWRdMBYff
mMGlECim2eiRfI4l7oQV015b7cigPSaVuJ1v3n0iMIln8/uB64+k6EeeRySTHsJ/
1LkEiW/CcLt8NQ0qgjCX+1MF3toCgoqjCyIsVZYCCAk4NpIzPHW7EI2/CnR3OLEb
B+12DoBto4H38jwzpIWZn8o3csVxkmGvCSJ2RI5bAj1VjMRLWaz1X1lwPKGz90Ie
hmqBinW0mm2Q8dxxQ5a6ggnT/p3AwCURx4Uc0eTmN7OHI3zvYHfANYBeIx4C0Fcc
/hH30K6+Ip0e99N+sLw0DjfWBpzG9bEwFtRvNGx5TYMonb0VqQ9NTtJ3IzG1/+xw
kcTVRWGhiUlbyXuHiND3iv/HDJlWfirt9r9QgIOwoZxz9rm5lJyMxBJ5fTvidRAp
cnEB8MmTjpzByTAMZ4vTSpb8ck/n/A4zsZ0DVcFm2LCdPapUFcsNYoIDgIZfoArm
HAh70acFxMo5ZzFsju3vzf79AHWV4y3r4Vt96Hd2bXwoZgBvThB701NDUSUA/lSN
XKTS3bQQiTVSsYoak4mFSqTqTD9VQfspQUIPWOR5asQZlxs1TzVMf323ob7IsJ61
U4juQ8DDt4eLgTkQa4cEHPQEuntQiKkvDcN4sGLiQ5uBb9o2ngrvBrIsq1VH0Lgg
VwPF3uOUDlDjCZ1BRHr+e/xixpkI4hCW7Cv4/mjOKYFvq54JMMdq7ocMCpgHub9A
fenYQ5Xc9DYHN0AHfqnFqe41MLuTJC3gW/WBTjqF2gAt2aNc13nQEhuPvSegKont
yfaVDjKSjuvD4OOoLb9j/wHm6BDRs3KoIq4E3PhXz1OA3MR0I4FqFuJOF4J5pYBU
vYJt7r9aWKu8Qp2rUozW7KXlSXFuhR14QM73UJ5PDqfcPL3Fm7muv3cO2rg27FHo
zW8aKwq8VF71AvXpKT2+elM1/W1Et9d7QGlCjQojf/fa+oJEHGYTPdsROrSA/x5W
6OSiqf0/hrn3w2OvgFI1u2Q5kFp5ZrncHn6R3k6fMdc5Mv45vBEZGIk9kYU2IWXD
p67rQZD6aLCZF5V09VsosBxZWR06B2dVkP5xuCihEXvZ5wBI7yZLaafROrS5edCm
Kq8R8nbJIkn+5tja3qdICI74Z84f4N9gBXQ2k3goTSWvhXrYTeOnroiNCAjpYDXd
Fa5DMXB8LvSIk+b/uqGTtDY5KlRVejlaYyVZyJVNjoZyIaFPyjEbc5Ehx6o+W+ZJ
bK29XWTnRsKA96DZ4fCpBvkku3sM4dwRHCNKuP+ILwWEzEtVLFeoYG3DZoSkY44L
lWS/f5zi1ujZ/5VdTJgFaYFpr7vCRsA/nhXlOgPfsf8Qc/P8R33oPq+qEmoVUZDV
YDYRdRHrbAhdWxZ8hToQHAk/muKmj164wYKKfUS2LwN3MpI9P38fOKLcuX3gM5Lh
AWoUdkeFFMUiBcUh+G175a1AfA2b0XwNao2p/1EBHh9BjvPqjEw1Jt0OaMQgd2BW
B+/qIUtqZMUbZ2Z8yLPVNdUUzkiFpC5Ff5dh5PCv83zK8XR3yDiu9xu5tu+GiGBS
Pm4JRs+VqYGFkS6KoEoqZRhuEs9p2+XuT0yamUszLfcShiodYswxYNB+KB9+VNZY
CDxgmbp+k6hcIJaOr/bL0exD7HTC3w6bZu23SYj+2pMx8YwnlAOaqWlgBzlp9/zY
ANmx01+U/gC6+2lS6OLQwy+66h82mZDVRO7BNupAsYBWMweNCqXchC2+KXl6jFfw
UvZ9zLj3pPIDlqRYhMksxJEvStBJrqj0MKZjC+bIjWJu/P6/N9lpRt4TRxOsl4aX
y8/uhGqE0YWDaff8gFGY7I9kTMNJnDY5gqb1L/5BR3TZn0wT1g3L7fVox2/TCVDt
fLE3t6yTng95gjFX/5LMtsH2d+KycxilSy7+mKQ2IEgYEDXDXOzzkEwquMyvLyeZ
q35G0LOpdt17c576cv3zaR6/OfJLgn06y3KIm3UQ9UETMo9smabRiHKvrJxd6Vt4
Rr7mbwZ/oZAmbFVVIlWgYDROylzqgtNIbEPK3dbJCVWqXphsbh9WjfdV6ayipycu
TZkoIqd+j9ZX1KJ9SPSK2+AL21oP/F/e/qIsYdgiCSVmQhxIwBNGQiBHyt4NxkGC
OtTIKcJmSE6IvK0DmKU7CqFqHHborl9UhfK0LSeF6TX0amp4HFBNrfjl38MKLygH
VNQU70BsqZJDft1VuvoEK3EJLMfQEKuRSGjbs8NUSDTqH78Thjoezofu3IeqaHPM
T7iz7QNg/bloUBf9t/86pEX5ZzhA5awJT2o1sR5zk/+xFdSg/u7xXR2MObYErLGr
VrWowPehi3yRFwY9wZZnuzadb8KbsZ30KgJe0FKYP2RV6wBYUf8hckkPpf0Fx5oo
1wfzCGhMl4zhP49ylaswo23mYn2mbd5rxM8z1FnRAzp1blx+It2J72+WLmtBb136
Tf+Cidnv3ZECATrmFurkFf8qUStS8EAmwLibf4YBlMEseaTKdXPA7m7v+IkhLE14
6XlTGLbpCYp2RNV3GisbplOH3JPDryS+bOXCIXMLgF610+87zucYypIfZCefUh4r
u7B1ms6XHNF/QikLClmEzFlr39XPqq4noainCOBVSPTcoxX1sh8Wt/ROag+rrixB
d584Nvgfi1lR1n7LqhwPkCsQ6r/H2ymZMV6dcrywpwUzYK/R/Jyk18tR2zaUs97u
A86p8FHyBJyrHe9JPQ5n8YR4sBHh77x8b4Fos+9NpxLc/Z6wcRnbrQQpRzfU+9mL
MWUaVlnYNtsbjlnLQjyRZ6ndOCslFpYJVKIyWFyOPLnwEbKpXZ5ksfVQnBHpheIG
MfK2LaD2XFOs+/4K4msNBhfgdsTxsXbbBw12lolVu4e4X8s32SNz9jpCT9p6iZRF
BSF8x5cUox0uCtF9g/kHegxMnP3pnTX6uhENM6PHIlcLrHoeEtHQXJInQks4Z8Im
COewpAqHLu9CdAs6D/3PyrB1M9woJe0WX8C5+zUg3EUyc9jYrR6a9Ca/2ZVYkmet
Pu5mibEDn2io5xNyk/KDy/RKDILIjMGhfXxozWpnYo4yEGWLlXy5cTQYIlj/zU/+
NA9HCxR44Z8YTAluYVRf8KPsO4cu/qOwtppIFrHyV0q+MyaAcyGtkBqpRT23d+N8
/E3SzYDS5/3I8nQtEMS4jgvUc/sb+NljHKL1DkhrQOzc1eyJ0KsDNX1qCmCY9tpE
PyBbLHf3/3lwTKhP/qK1zJhAFkjRXrSuJMJuyM0qunWtMPgIAGmMOg3gKGYgVME8
DJG2s5AUIH4h29WEvxsRj6OzRRI6Ojo652Oer9KLbi3XwkXGpIjloZUMr5W5tBSJ
PqcQf+f0GTSxiO+Yj7oETT7/JuRrlIhX2HAAQACNRtxq5lWA48JZ+Sep/E3gqJ6v
cY9B3DBYzrozV3v+UvgEONHPCNLvq3/et5o2wDtltUvRqG40t/cKAxl2IQkr36V6
QE9ouGuLSbdp3A1x52juYYhM6HwJ9KjDe37EB1FWw1iz9bUFJfdlGq2qz8czmbGg
gYKEdmd3PhNv4x2ead9oXmGmA5KvtfG32nGyA3Ppm+smtJ4CQll2yWZGbUj3cfx2
udnkOgb8rsSI82vnv0CviMimRvAuthqx9pEFU7WdpLxqTHaQOFbfhPNsNHCmvWBl
LcKVas7psCAs1TUMCEMphlPyjLC0Qnj+TT7/JmOFWHcWf9FHVAF9Rq1QPNXOxutO
O0asRClO/CaGdR7pBNwcs42dfdA0mhPy1R3YK+Ra/43Luxw/oUXCiBU5yK58Cw7l
P4JyV1mCP8F/iVWP3b2KyXBcFvFl/OWfUgmhzyRySMK5oFH/1Zj2XCcmuTKVBsZC
haV79JJXOh5NqfaBg5/mxC9qfkLNm56ouJ8lVAeGfEtB6HMjKwuq/0dYgZnollvK
V5+FeflptPS/E4tVkojLzK+UiY5eIsC7F+tAq6/KhptrHgQsJfMtXoYMndgNBF0j
ruBuZGTt5kBVq2xL9dzDwQTSPjEeHijl1EI0qD9v5MjbnU6Wkw+GWMpleNR/o1Hi
sXNi3iTrLSwxnsfMYH3F7fC8tT70gKmglyV88/SJFFmN4QYQV/6GvOChhn5pwLzC
g/06QI2mAIJVKgaZ3ALsNOx7voYysGFByZEC5FIaDP9xUx/i64Dhl1L5Ukm0GDjY
x3kFBfa+r+HDqoqOEcTsb2aGSQfVzNvMpj+ABPApDoycqeyS0Ws9UuK/C3MxFbja
qnG9fVZBNvrx3EiROnybJt+rrtKsKRwKLTnpS4GPs+HQRD+g1r5+b8CsP/xn0sqV
tjErZaeX+yshKmPmq3nAQUl6LXZpSueHHVDLu2Opb2pKR1XyYRaniWXuZ5ju0N5J
QnzpqD4q/51llNxeRWhilpFaKUU5JKJB0Eq5+RakDhPGZLi69L9OTnuazTQOSxnH
kSxLjkJvl7aJReB8iMeJWG35c3gDo5vA4YeqSgRI5z4ikHi3J0/uh6RmfLp7PFjr
CsxrsjlgAo8pTEwPLBgHhNGXIya3AnbbOIgC1BI3S2z+U9Sdl/0+elxiDabIbS5d
2AxcS6fIDc3GUuqyVkrR9PeD03jqkz8mu6oXz4txmo2KqsgWUH7IHU5mkxA5loe4
LYWpu9GCnUm45RUCzj2wRSS9jMGKJX6JOBcHM5uQ4eS+n2o4yNnZPwZAmjeAd75O
iAh7aSEI39wht/8QV99orsH50kBHb78b7OIVzXVzNcRkOoRaZ/TYFNHvZTbAYc0U
qaw1cTc+eOe0U3ovKpNw3y44XvwXd+4RxIK64I7wChFVi1lQHDldwhXeVuHyysqq
ECcrt7Agp3qmLTvbmWs7lb6eANPr7cKusuMhcxXytzlXcCX3k0Z4vHgaGC6nUgDw
xqde1ZKIt7bKOZeFv0zi8AR/S/T9VOYWSJwIPU4JoI6Au2mICG0a/2X2Qav2ik6q
1zloH4qvphPD1deSoruk5QYt3OxSdPRLhUpiI63gywdZAW6ut7VN9+kitJx6piZL
pcBELGxtYZ6R4mDIKzIta/vxEN732oo/ChuBHVtR8JIDVYMpBe2OOaWjBDFGHj79
f1lNqgEqJ1mvBVOzxp3CNw==
`protect END_PROTECTED
