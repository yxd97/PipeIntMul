`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwV7JNuyBuMFksiyDHTPLNwKQrq8oBSaHn1NIWtIgDoOM4xupmdnqF7kbFfSzFsZ
24Rew7S8CweSpflzvJPD3dxtwvg+Ww35wnZeW8w8+MOLXlZjFm2NSTM+2z/vstmP
p5/6atv2xTOHVKfpxs8ltR9ZTtLO4qH9M/syIBcngbEOhz4+1nv1FD0uq4VSV9Yf
t1w1G9np2gCfOm1ZgB8AAs/KZhGB+YI2zdVgmRWbe6EUWxJInVmoxUycOrXWYlOg
R+QCx5J8+oZvQhVkD4yHPeokGtHia4fgoScnyxNJpUIfoPO4QWulvg2B5/+z/KyA
oyCEhT18C+1M4QET9KGD65dCcw/TnsKOAgeE+akSxaqZowEzCUskZLrWtJ8LYIum
5pWk302LSoImnvbfYqU1nw==
`protect END_PROTECTED
