`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sdNU7tUB63TABlsRkHcfkBL3RpnCzCjQlWxZLnV7RrUqk+fTerEGXi8hiA8/+7wA
4GqIbk8sS6GX8SG3CsqYnMY/xk/60/1go22EVYxJJmuJp8dWtwTtqgXVkMEqTUXp
WjMTvnkQNiuTh/wU/3z47XEjC6ZiVFfg+e/pmlfq65bABEXoMI8ar2InzhmdVpQI
xyoYAjJ2uoKSrriYojN5vdUwfYNaqSpHAFVA1Qa99+YoZtbyp9NLzOzGusNz6O7j
9GHjuQlYcsddchLU6aYKs/fDM0SWw2Qkb1JjuKssSxFS62nVRjR3dgmmgnMDfy87
g7uljcWPXIgMLAThB+AdKOYQ6pxvb03Uefm3odha4qk0l0bcFVBRrUumMKxUIN1V
gshdiK5OV5Afc4EHmzeTSnbNQcalmlOITGhe2XJD1FjBKNmR20pia3bpAo3+hUUu
EgFE0v1aG1ZKHtGl46Aw5xigRhAxwDfbQ719m11PvLg=
`protect END_PROTECTED
