`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OjjF6JzDNXDSnYQ6WypPshVzwrjA56sRn1p/Z3AWmPheUhzEeZpbCgrRToMqIIJp
LRRcAGnEc4FBzKp2UV7zgOejNgDHwiq4Gp5UN90dUD7I37vLU+z+GWqIz8//O7VC
xUBpvdV5mGbdyCL+PovdwOjeFzAruh1S8LYHNCeVoBIfpn7kbxcxtgS8TtApVA4P
vyjtiIEGHqRL0+X2PAS7pVubusLhXixxnnD3ntfiS8uSga1EQVT79tKatgw/bOh5
w+MZga/ZeFmk1kpDttnFViWv1cq6aK2PVpZZsvWzCUfBMRJn9yxieUh/lXFCzDmS
Me9umWaiBa1xwdbF1shFeRT71rx75RU05oJsm1kiRh4hiahR6q9/AViQ7oAgc86W
oUFHE9ihVjcs74sbVRMO51puy5TJ5kxbVHUPjCA8VA6QfY9i4xZSn6uReYN5LJY1
4KY0D+aJw5vBTjQ036IwDKqSmbA7DxYgmlzaSxVjzyU5+4oW2mKZOYyMnzMS4/yI
+dXiGdyQ4zpcTGyE/qa9Pd/NjYq6A6egOZO8HlWkTS7gfmp2Tus8FYXfHcniFEnl
J366BvL6i2j6RGCL3vTR9wrQjH6EjWg5HSJ9S7mcUqwBu7JS4vRdEzPG44QhfGWi
UEcggB3kFGa7hdVevFXDUCrN4aG2D5K54CM3ItSOggh3f2Wt9QF1F6mEFfSpq372
sIFT6h0TCyc2CPdqP/lwe0vW+SZvFF/BsHYsGDeYIxB+Tmm2ixQwAXkcYnwkf2DA
WWFHwl6dp7P9GjQodhFNukSVF+hmg+51QEjAaLmm0M+kPZik0g0LZVUsKJJT1z3Z
bYaTO9qpU7dLq844kE2oLu65x8qnRp71nmt+ZPd+hts1cwcLk5ox0r7pEifQM7mj
N8h59gl2K8WQhk+ZFKYah7C3JuwnXtlSowQ1vmWdNpKVigx9wcxrtXV4UUGUsBwp
`protect END_PROTECTED
