`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X3tRM9ZI8ni53rdBod//1tT/CQ0aSOq+KssKAKABwI2V5DG/7P27DAf2jGBCBR6e
1d+0NstslmeejU+lFExebaHCyTFymOc0iZVL1/PMyYPaL2H1papd2kaIbfo8Y64P
jqXfhZJvMJ/VdRlFYjpyM2BfpgKVQITpYG3vAV7vFFA5F4jYi3cnAl3fNsKMugUa
WG9qZRU2/bFELdohKUz8ADzi89OpmhVXNLXmfDo4Gldm3y3Na9dDDroSoXMfRyiZ
z/rpSN95b31ygi4AQrURyARPd8jBpHAXqw34TBEn64RMUpGhxaLWKYV6nP4qb6d4
wVgCD85rO0VtXx+nztdpoyOA7NqnNI1y4Rc/zpC/rjvnUyyvuS4TYSvBD/gE6gRR
vw7iSIsPounQWIdA7Hj6ydV9zEWrdenPVBGSz+5NnGRRcvR88uxZfqfAOu8EkoiA
K9npmld9GuCANtsHZ6d7l5zMi3L9qFpHoCOpbHM2cc1pmIe/d7gS+vv6dSL0BlC0
V82EYBFAUVejdXrTSDAYGrdgTs1eHOXTgJWCXez3bF+t5ZUbYg+nLxTv51NC/5Si
NDKTeSJDhr0LNuIUYLl7hf+K3hM8zDGyjbBCEw7PmQzKt9gL3SyosiFLlDAaMEvT
fK2NRWSwBYIiYlU2DSBqm2yVG6VdHxsyH0TNrJgWxgMkvXHWU0o2KN7YLUlgPngB
BLjfSLAGZfZRwQerSNgCCljdyV3hc5FfsjAUXA54LEhH3kWS6TKJieQB/prBXHNj
y3gJcbYKYv5vu8JMrVRwKZAd7x2zHBCNoM78ClvWuqiRW7PmMXTxf3PfuaLHKNtU
RHFThVNM6tZF4NpiP8quiFBV7FfG2Uk2oz7EUgsF1vrK7zSNQomvhITU9rVufNFh
tKHGx0pPNktEy8qUVu0cQ+ikKJ6OsDOQSOfNZIOBR4/DSE/G/giSJv4FLtWMbdqS
AcNELcMhROqwBIxxVx9JwFIafFCAVlazFQQv9DDg1q4i5sU2l+G5QicxKOu2LOYY
EI7cufhIu6iD7jAOLGaOnxKnrlAWac+kYxb80ib/6GWUCAWnruxKz37Lvbr0mOeF
4duEVTAQXVaeU0+L44mGrg==
`protect END_PROTECTED
