`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jGhFe8yVQDviRNI79mGlxeOpVLUTLqLbIjfVqGxNQd1ppRw0u6igP5e9xEFKTy6l
3JyRJYVBNTf4pqtEtrp/wBPe1wIilzlUI3hGRR6+HizzlDJKNXE7Pdv9DiEL1R8l
LNL4U51JgL6AntkBMPY/FnxJWRkOh2wAytmmFGt3FLEgqh0ApcO1tduF7sTAPZY1
+bqhd/PrajNqw5DLeqs+EIAG2L7hExt/J1B9c4UbOqFlUBu+tX78p2fno+WcQNyv
xcUuBg9NWNRR2Vr8fh6QNIhM1daDJ03NjqYrAxheBSsfFuvrGLIz8MX7yJTI7uLX
hKdMOPkgIydsHAztB0nFllXwZvvMairHClbWSRuBSVep8u5e9kI1de2SxOHeC93+
tiEeHny7Z47R9azF/DhoY5gE0URw1FcMgKY6bcJUl5bl/Hw5LKnsGkK0Rr+kIL/G
YtCVYpVB0g+6A3SrMMARi+6BoczEOIO7cnaTRAmmlePFfpJwHAOJRauOcMK9HsYj
hddvFdthA4Cvg8JGZ2V5U8iJHJJWZmKhNVaIkUVOIKSUWqnJTNGf3eot3HH/XYhd
lqRnGOi8wWV5cBhTU3e9O2XWYUpXPGxgtoB/bPzLwOiBIRENF0cx95yTWVolB8RT
+MYEkMBdl7ZOGqUeFzRZdjkazX5D7OZ7LifHIrnwPgV6caPIFujlMi5JoGvjMzuG
Ze3v/lKHbHCdLKF8l2RS4OsEcIZhHK17eljUCkb+KPDY/IwuyldJoIsZXsxZR3Xs
0GvDYab+llHCaM+kXaJnrIWJctUiu2QV0Osas5FXJltIa/r2gNMZdG4F3kvwWKP1
Xwx79uIm8oLDzWpfIGWHKL716xf+jGNPSFTgFlV4pOgDrj71H2ewrI1pIiUzvN2M
rreyosxcBGFWMT6yOxeDqLpY2JZt/OEra8iLEZpw89jHp/MJxEoaYdxrUe1u8kn8
JHAkiFgzV0IwIWgIqce8NsxF5N5Qb9dthpVZ3oCFboZe7P+3eeE0eo1pEodQm+wv
wTHBtqnPYVikqCERSTU4iCkRpfPU2lrTmYT02SrbFf5gsVPWzdRaYNgFpXWh7l9S
U5HmKVqRa4eX+UbFlBk6XJSMlz2rTb+h+C6enWqCW1jTQK6s8fIrPaaDNU42ljW9
HuVuE8PpRbwSNvKFqfMg0JWKi6cEe4mx/DbNiuJzpl9rFMWcYJIt7b3vYLztwX1F
M5b6ANcfNPHWq/yDZgXIK8ed+73WLt1kr64l4pIhopsN9HVB4MVwVMLU4YhL8DOq
dV8d+SyMjlzKUaELRB9AeftFcdBqNWEQJHD98IGvshM=
`protect END_PROTECTED
