`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T2jdocASzXflTegjZliiy2u+43AKfiIHFXaaZfq1y9Nj4UfPgsV17+YZZojx1/1A
cSaTVgY1cN8BmiaO6u51IVcMPz2mVh2qF8T6MZmZH6ChRM57oATGDBW4yQZXKiEN
38Qgyl2uCoADXiT+ROEMWBvwKo4VFieOYB07H9vMW/Eqyou1sTEWhtHJXUjJvnj6
BcH32CjaCry8U/xQGDn+rEUFhNecKaTtybbzBPVOVSdAg8BZBo84wCsQFLvDvxLb
foQrB1ALQgYOJndNKMY6XfSA6GWhgNeVG73OAIv7dOetXlmpsUGEVVrwYyCaPEzJ
BGFdR+ALATYrqe1Xf5vJXZAqzh0LrB7R4Nmiw9B+V0zG7FXoX1DteLZ49zdd5D2q
F7uUD/Zwo4jDFkXOqH3cOM4tGvWX49EexTeXc4FRxmS68SQoD+6iH7sGV7NBsiia
`protect END_PROTECTED
