`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aDcWCETSIQWhZ+pr43x0QNwUZWERetRrweFbap5au7sp5QEla5Hs1ESi1LmLOGmo
FXZQtJbm1zLJcnUTu9B71a35TL59OW729IAseSV2/l7psnfw7LBCgdNUPW7/R2ZX
zHd4FATkerQrATzAQuudmNzQVpFmI5WGUiHkGEO03s9q7iAGmrfo9+kSDKYO3Tgb
UpR/PzkY0tYfuxMhvVKTOQ8vT5cPCxB370BWCU8bdcyyrH4JFVjx/DnXS3uxoD/W
axJuaao4ZRwZylE3JaS5mkEvJPnMGFkMzl2gXHj7RyOtW+9HGUFq/5JiBBfOYr49
tx7QDumSGt+QeVLF4QB8ACJ0wko6qtauTKAJe0PZAEh2kH5mYiCCti62Vvs1FwVz
dGW3qn2Sr3KFQt1K16mRJGgPIwV20gFv28Bevdp2gx6ZT8CNBsAAqVxcxa6p8hAr
SptJFAq8HP8HATlBuasg1qjIEOpdsG3amfPhLr1rPJ5jczHWR3XXOqOMRF6N4Xw2
of8XNgMhc+4c1r6rupWC4CjEgxvaJteNdM5PmAyLY8qHja3i7lSsjvAdK7lsckoA
dKM6b2taUCw/mQr/agEzdJ9choI33dsc36/LFDLDcBDNL6vCXzZk5O0TRbuMDASf
PuNcFhGvpjJQRbm+JwwLby1g5srvnRl4o3wpO4ZCYDdBbWC5vj4lTSZ0i+RN48IT
WR6An0hyng02+IaHW8ggKVTGmq47AuBVs1T26YS9ESd750inOGrXALYEDNA9c9Wc
WspMGzj/fFyaaWA/V/1+fQLr1sqUKI6f6rEd77EgbzAOkSNDQxvU0cL7X3/wUvTs
9lFDfsQqXjwECGRSdmGl5DZ1XYIfZdjd567NePJkYvzgZM1ZR6uFYwwYImfElwsl
Q3CkAN1H3g0+TDBzBf4GIO1U3tMjC7v7mjpFqNwV49nWajSofwtGSmmmmAeQGjkD
TpU3BMVU9nhxTLDkJkxYyUXj9NZ/dUTdLQ6poVSSYDf6TZGPe+LDxLCnwpDLMn7W
IKYy99D8x7nVCIhl6gbHXKpJbgzGEIxGwxWaK0q+GnHx1BQakGnfEZFCouTbhZYu
tT/hWnl2c1q/ruFPa9TKRiOeCgSysjCGuVQ525n5DX3suQjFrOD1XfiOyUbNlSM+
8awmpYbL3uqOmqZRYkdLY0j2QbPvI60ezM8tbbX5LTvrZ2RuWCtdlAHlvRO0EzbS
na8PKy1F2RQ2m76ssHhWyzjnKkf+j8SgxQkOuYCQ7yRGcSTe49xhHJ3hPCaK6jnd
2VirOGi2Pdx3mQi/ML9dV/yNoev4GtLagg7UdvvY/uk=
`protect END_PROTECTED
