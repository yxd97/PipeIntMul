`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wzDNWy9w5hhDXyaSJCn6fpG9pUFzGtADHYf13R4wXz+I/wF3w9ltTVfX/w4xPvzM
xRlLGtUjN4g0/wbEw+zHv6VcUsLiHGRevt22VbTDqbB1E1P//M633+9RNdf/vfYv
63tQmIC71z9NLluDP4pK0mdfguquMzgONgac5kQZrj7L2DmvwCySYmhNyitCZFky
ZUQQLJMVrLqm1RZxzElTI7dNiuMg0AkjekTZ2t1dwmIk0hLGJKJeaM8jB7cwWPdH
QSm1GqmygqBcjecS9bvtuB4QKbxaq1l+wYzxrLD42raw2bF6SOfu9YfLM0s77/ql
JKTsvoPvZi+SqD4DCDHtGokB+9ycdWpskT8nhmO2hO0TyQ3AGmSeB7m1kUCyuXVI
kya+yn4uqoxCASGTMn5xlHTne0Y4RmzJj/klwjq5sh09yVxGrTAJOrRC8Hb2hHhI
vqMeSnCX356rXAhbAPA3nZMNRkaT9CUa9hkr13euk/Bdvd40AZyG5BuXmW71H3YG
sTH9j3J0+x9ViHQdtebxjGCYPJO2ZSHCC4ei6TwEoGA1XWbcw8UtWy+/uYaRqMhL
44CSd9xKr9M/iC6DF76AB8RHpb7PFPxpnBltEqqChrICfnLY2NzoqSvQtKa2B0lQ
`protect END_PROTECTED
