`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sRn6arL9rbN8kxUmU+ZwTkekLV4WmyGcteMuuRIuedyXpzSi0H6FRAtOjN7Igjyf
fRauySmrCGXOuBdHq+jd+YBJ/0rbPDqBiETtG95J4lZm9H2jgaNpT9h77vxQr3iP
8SBASABbrfUvK9fal1yFaI5BhFJq8vMUKYVZSQbHZovnNsnwY/Vvqj32cMQ/CS2R
b/QlRYdPfD6UUhPDzbtKWSg6760yhAhbQTbxGmjmDNvx+shgjD+SxocezHbiiV67
l4Sj2NKMtlVqi5ZUfm/vtr0E2lK6C9sYnyrh1S78ABoHbiH5VrTIbOWtjE1g04GE
qlfk5pt/9cZ2ZiMIaD9u44/P8GfQC4WNFv9I3nj5LekiE37VlmT7YwNT3msFSWWS
IeMl8Ue10kGay/h1/EhcWoiNq0YFrNzlWM6TcA+Cv30=
`protect END_PROTECTED
