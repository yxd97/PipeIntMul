`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWy6kWgd773mZUTJ+0EL/BdZSkgrLia2JqYRa5Z2INX3RP3Um5uDvf67YpQVC8Rw
HtZkEhB4WXdAhTLQEXvYUlDSBTcDESEf8wS14E6rqGSglx9vtcWuTNoThuBn2Ag+
pWjNNiY3HXe0hVTTBvOX5RW9NdQGR55Ks4SEJmsi9PaafEYJICvSV3xgMWughFAi
Jpbto6YQfzmwJmB6LtrsKW+OnyU/qg9S4OM5wObdvsEOgYQU9H2GuP0+JBhXMbrm
QjNyZJNt1jy8CxzqB7ZSj+OWoUiVniIHbbKjYJXljHAAxre1Ey9T/i5cqKaUYv4F
KIU7vxV1Q+6ok6ykEPYpcTMNOMEcdna0zc3uaws/zcdukrviZ77cD9xN5JMeYMYk
lWAvzOPbHZeYjHBFksxDxN4kV9dpLh5VMENug/94DSo=
`protect END_PROTECTED
