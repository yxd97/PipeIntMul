`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eQ+yQwUT8J3Wm2U6v6n3+z/Xly4q7z3lkZJCb5kRsrZpedBbcDoIibT0p+ZhrUhK
QWQ4h+l10GTrCTcgtLUU1bTBVtCcrVUUXUOcKiqADHG5kuFgPKNdK6HKxLYn5ZCB
FHpp8dOa7sV5oCQBarcenBBs98SzQ/o2qbuB1DPTHwa7scPmeEpf98xA0mlcjo8o
C4ratyGCykDN+eAVQp9CvDz9NNxTBrFHjcHOGxV+igsOxIvtDlwxCzWXGVyOrCkL
VUGVVBFJ6RxdwP/wfmM3gr0obwMQc4ovzHBCY5AV3q+Uld3GacSEDglIR7Di03wL
LO8xkLcCnnZSZ+Qs1DkPbbI+cjImddIAzzSe0XmffW5ElUjbSbrSCuL+0AYTxF3r
SQ5S9joNehIuIMihhXr4h3NNfhYiGuS9AIkjOW18yQoIKDLNhpJXZ9eVQVipBE8z
XPz4venkS4iafgUiz1cG2j60JX2A8nYxjalkZE9VOGT/n3GjLP8xxdEVu7tcR/W/
8EncHFlApMZ4zxhbySwEG2wp0bZyyT9XUlcXsS9WD0cuJYThNiVUam+VD86ACVOL
i6fmF5x9T4epwxK/snWxaWsiXGMHhHWhmMV3LLhOkD5Z1Ql8ofLP+Ze/69B7w47b
vnVuOigoNBt36P/y9ZZH68R31KRzDK/lBQEh4jdUTraQC+pfEBVE7v4T+dpxqZnR
FS1IATYrPkT7Is+nrakgWXDlTLibrE4Ks79+cvL2lURIkTcHDCo9r31Z6Ne17pXq
hdq4V0fQG11wX8IN2QluYGAwF0QhGyRgeE2YcYDLirPIyFIur6XWBa90XcQ1zllz
80OYjOpGTYP/FrYdr/7w99hSjUfmntActXRd54k9nvKN8iGU2srsGRIF+wxZ6Xkd
22PVvy/MG5GpiY9XoIVKEaVrFux46ECOPFVecZ5GkGIZRyPK4uBYspGjYBvDCI3M
91Dtnxe/0x4g5ipM4+LfCZXWXW4KajSpxiuban2RwfZlATFXOEM1HXWAv9NpoKzr
zVUiWlEXoqPWqJH6X0v4MCSrkxVIYo7XQQ3Bm9kB6wNXhV8ozG+KInZOOYSDnf+k
5Y3UjrwBqe5c5in8XI3Zn5yeHQfETIyGQ/TeAD66Ii4JfvXa4a3VYQL671TZSBPl
yWYvPisBDPeXhI6iKDe3bnJ+kMRWWKTzew46bWwTbgY0rIa4dNWtaXozgKybyqo7
3Rm7FwN4QWfej26FRKR59ypmwxSi0vZ3JcF19oeEzQnawvLiXsp1zdpgcfUgyWTQ
dYea9Qi/Ef9nXltmFmEwvBqv3h+oj7b8BQp6RARyn9o=
`protect END_PROTECTED
