`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLCEZGyJeUjPCkP6Im2/YOHdit29+GcIcC8LI4/ikPdCEDGTDJgUXb4h5CtSadqR
/k1OqCqNgzwkvUsG0XotCBbTN6MHVhbKywJtuzalpJp53LChkUtLNbmdLBGqniec
yHQRbrlz+wrUb74yIPOn7FZsQGzoNe2BxJ2IBppjEyFjPUQ++VtWVOj0RVbWpazK
fcgsZmSkdH8Xsb1A19wn4nDBGXnRSd8Jn6zCGoUeXaVN0EwMBe63dWU62CKIVZmY
jXmD9oCWMLj6rkQGOrOWNHJhK3x+Vncar2RYdBU74GPKV97czhqi1O6Lgdkl5Xwx
tn50mqGGsEvGD5MUe93bfWLCOD9Xyp1Vy9FLkHyH/swvK1PRQ3THdNWtZzpek2Os
pywGmurIlC8RhsWK4J6LMTRRKtbgrI5HHLpm/wDc7WJphuEQl0Z+wajVNUhsm4h1
oQVV2t8pwI+HPOtJcAuDw5si5+mpXGcrSOVuCNRa78Q=
`protect END_PROTECTED
