`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XLUMADLqpW3YPof2+6opMQE9+kJF6DPIhXmBmg2o635tkt9JVIYiAC9yFDUkUEVz
z28bwI1+bHlF6gm5eJlAy7gLgT3cS0+2jjAlWzUu0IuSNxMqumsVB0AIQs6UIhug
e1K/Dt+v+z2vo1AOf/3f8os+T6RX+B/tu+ZZRHQGBTsh26Lyl5izWV1UWuWg2Knt
2v24YreOhEyAmFjUaGeJ4+Mz4ykjSp/S8vGUCFxKladjZpZC80I1g10nrj3UTZ4+
8zHDtVAvUjM2pm0sPa/n4EJSLX5yAEnIshh3RXlNGGQRz/ZaAg34as4SwRrB6mNZ
J3ub40FB9peET10tTg7gmeP5kzSUA7bCLNebLtDhy4mRRcPycg2eUlZb1JVbPlSl
8FA4mWUk2RW/juIIqgfI8dm0cAF7RZZz4RAPk+5zMvBHug6i8S0xFHyPLghp+dnr
`protect END_PROTECTED
