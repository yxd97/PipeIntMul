`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CU/2gpTqreIUoHJy/FElaMyigIYRWm33ySjRdt20qQHtF5kSeo+m3v/rATtWXb0y
56mtcIlE37S7WAvUH8U1JJ5ohvdB1hohwjktZuCofSiBnXdH0hXOHq/Ueb0g2wi1
HiXc5p/aNJSe6GklpUim2D8UG9vwXrZzLtY6v+wUx8ycb/0BPox6O694KtP53VM4
bk5hR/o1XOxBoYctoyVOZgH+SOccpV9LW2PGv7CBVrYcJhIZhZp8HmNdMiPmSSUb
Ha4l45ZSqQcoBpuRbJUFAqijSMLiYUb4kVHLTVQTDb3JgNpfKZMwuM62WnkCwKaB
/Yeky3BfoqRb0zlACyzjOtF2zrv8vr7r8yLI55C9tl3uDuAa1e+EUfE1DRel04ME
VO8YBT5wZPUuAX/C5uWQqq9jCPxxvtbBXJjd9wuFBjgYV04XkoiPOCsGtmk9ZLH3
`protect END_PROTECTED
