`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LgzeWCulF1hVdNP98+Te9pHOIyDW84pNo0CY/YLgSfbIxWaM1az3vV9uwy/xbDKh
OEXtXyk1N+v7ql/7Jklq9op/BBsMMfgXGpb7Lzt15YUJwbNfv4l7R0k/MCmzeg7+
ntEJ6Fu7TU8tTOy1CvfytNP1/tbvuIjL+fnIQ0jZjr6MHA0dujvyxz/ug63JJ/yW
u9rO8Q33ZsbW9Cl5SA5IGUeQw31SJ6HPpCXHe/+G/GpKR9eSmy9jKGcxvRCgCxa7
+ie1gs12jsPyYY42gBiAWLbSOTQV10xVIMoKGgLxNhZ6uFTFUS7dmZjONCqGR/k+
ztYfQJ9zMcaDtXAPUp4+WaB6tiJj3NKKM4bflfCNo2STKpYalRrEjH6OrcRFp/fW
TLtAmp/jStTI5XfNn6ZecOG5N4ZVXeQysHHV8DekcyewqW4ic9qjXFl+DRhxv+Yx
+SwQhpVOH+WHa3vjTo2Q22Mz87JkLK7euYHflCcicpZ7q2DngIaS/22iEOCTpnbd
Iq0Dhj+4LWgIVNKVPNgDeVSOc57LSjts3vdyCcHcAYdSYh13P+k/T9L4ce/ylu5t
cnkGah/JVPi8fP4LIFBqdPEfro7x5uNId1wOlaOw+RyJ2E4bp9NlCG1NixnCa1lI
yB+YhMwUbv2KQPCit02eXl4tYIrO0I6hm6dKluTAget+F70ItjFRvgQym+u/k0yL
GfcbaibZjwZtR92zY0mtng==
`protect END_PROTECTED
