`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1vvJIj8cr6SfKCcYG470CYmSctjagplQ0mt23gdCThXInjUGmhtbb1RtogZBJUet
Rcs7N8hE4CsIT6BIG2TimnhuDTHYa0uKY1LccjJAOKEO3KWhMQ+kWKd5CBTKDVXz
DTwei7BDCknHBnzuXuc0ZEcLj8rofWG5YvnvRmQ6DckU6pr29rOtOr3LiBePmdCN
mVFBYOgWJ9PZMvFks6rbpMiKthZGLiSmoQM2IHZ6BQ1UabpB46rNH+J/9eR8QDTC
qtwAx84TIRhhcWClxw/ODEfZRTN8E+ASR9oC8ZCfY166nkNnu9C0Yq1SdjbffQCz
U2lGZWCOB05c6Y/WqICtoMW0rf4zdkHJtGfesCRHm/Z9apJmvAOS71QOtQdMySPM
B8ivRII0OJAev7/J5HqM0vqtdaaHtZrROhn4T4oY/uq2luuNaq7xybELaoHr0DF4
Cz2oU4/KK5AgFJxIk1fz00dPMup8q4T2W1Efomtr5cbtaIU0aAkaSVS+KIX48MxQ
iQXWOIMRHcvTRSdDze9NJIzVKYXTETLuWQUdgqiTLqKVHoM2rOgCRa3UShRGNd6K
qrnYgKtKDfWvgU4/fLVqEQ+NDGPFOs0HL4Mjs+11840FvnhDssbr06gWcdl/QxVS
l4UYLAmkFM/7TwCEujdiRrp+n/rZo8UOCiiIGNmJYqtYrOxPXTAqsWrjNlVOWJSZ
jh+atlq5f9Ny4OC54RpBKM/OjWloTss+AJEcQAhX3MuWo4l48q69OFjLeuw4vu5v
ICUs/4H2H1l/L0Yfx6Saj6PYpfJR0tID7TAI1oXN41FnuLMXQWWNFR2e7H+ATBBm
Y4j5tbKe+RcHdG+csPRqRfLgH+3GmaNKCad8zGRDxuhDpqIMIq2BWudQ2wdaYLgi
OWxq35TUxzvDA9HDEfJA9TGmFoQrVT6vUhux/B4cF8mgT8c//K08lIuk8FGd1tr6
KPdClN1YIt4u7weOQyoa9PbWcEZ4Tf8xQfndhVsRyf3IRP0zy+MuuCiWwhwX+vXu
TiscVRUs+CpnFd5XECDEbQv7JIUC3nwggPxULrsdvq6maG8/YC2RO8hn/N8el3gg
KJB0WJkkMCkZxvkHxywv+nb9XYRow3XEhgwlXGehjnU2rCKrLiq1fJOmiwu4H5Jk
wM5ivvVbHB74M/aOuLs3asMyxgVk2m1OFikWpPbuyoyUqAOEDQIiztcC4C5W4Pk8
OEE5gXFwc40hk3OQN6e7DPWD6504TAhdvtEB0nHYKbjjYkUwAsexMNfPWbxnt/rh
/NcP83pM11RvP1BEgoFn9thzY10FFER6qHA4xR5oJ6i0paiEGNQcjFOl+rUDeK7Z
1rGHd8WLz8HrII78KoE1oGg7AkyLIKi/t5dmpUjk4fE9tj5hoofz1D1J4d+EsItX
blVc3XwjEWy5lc0ZY0f6PSNhrd2LfAMllIC60r30GpSF3gc8UF1F9bVVqLHrjI/4
83juTVpQxESwr/Y6VVVFGVL4yR6uRqtGIW4w0ktue96Esa4pGB0/ESy+ZuUP3qIk
RV6wBRBRolTKPo/5BEnNOzURZsKqG3FDcoLr+tLwPVyGYHccPP0Px8+At9pzDsEL
hgQJXI8wihEWE6WH18tti8NW2QK/J4WUNFRJTFVXVq4s9jXzaTJMJLeF0BL+Orx6
FpEM/slaCptZcyIP0voUVTevdo2XN4pK2MXrQIWlz4wtdU3hLQjSqYT1itx7lWKy
xgU5e1KMxlks386X5EYyfdFgUtncpP31qNiBRdcTYG6hkMpeiEgybir1UlVTYjxN
Hb5r95JOEZQx2oHzgELPRCv34vpXMotjB3iH9ShGEbq2N4/+LatOgphH8GR6LBe0
jikmaSd/O2cRV1TJZoSxuwZ+kzJykmcBRNgZz8mrwpKy6zE8tic01fKjOrvugp8I
06arwpvuCRAp0jpbrXXHdr2Y2vaycHobnCPxxVeqgiHjIgYdhk1lmGaJigr/nd5B
/vHFnbKLrxGOJrXWbkOziZyN1x+JVkAcp9F5nxyqPmzY2hIjAntWOwlMz0rMemDU
h4YzUkvBeaV+XpQq5OFN77Ubnk4CU7IgxN+FI5tIVqFicS3PulWH9LCc9v8akgGU
OsZJ8GYYg6AhEAMHSP01CbKV/LFp+qfR7+iKYwSbMcJuJ9KFCsnBaHKaoYoo1xu6
ThQAbZBEWVPeO4S4ME7spSvaVEk77FqE6O/VKxEJGJ1LWFXLmxp4gnqHMsE/wYF+
52O8sCCh0dFABkSbesAAfl8r+XgbWDN209NNQpikV0nhkh6pDawj5pcZjmq+wvj/
eaBJuvXbZFo9XYbiZgiVrP3OwGD7mYeH8LFvxW7f4Mc8Jwr7ZSNGD2ZObCBl/zu9
UgwIF52XTVReW1NsxOnEjn56nuvIAh55gDdvpTYkaJI+P+068Fmd6jdk/w94n6Uf
619y/p0xpNR7LLPkzBivaPFD/X62cwgll8A0U5Gy63xgsNmjCt7QeqotqDg5JCkY
hEFzX/EIQtdSG7HUIFmmPoKheCqVPmIRPd4Uw4h+lTXkYuWAUqP5+bHGqkcw2wac
XqFR9BZWglbxCNT/nM7n21WmYMoz7NhvUOQIO+KYq7Xd9lSfG9LcioHRVjS1+RFS
b8xJ54I3Mi3GJhkAfJU82bbanlf2siohzURSxhXtKiKXpIOCh+NDhdNjn6HAWGBW
ptevRVsIm19yh+2hy5D2G+ltErLoVFzrDUJiWafaKmKPzPc6DULL/iY3a8IgtbWr
EyHxXzpTYiEeVZHKV/J+8MEYnxV2Way2vDozjW+SBDzmdQF3eXb0Xt0+gejVU2go
fieJXJ2EpWZBTetNU7tOoFeUUWTA0qm5jCwdGNd3PJwQngOKC60t7wMIoOodfaeo
cO/B9sB8vj7HhdnRL9VOf4n7vBNmruURSrQZ+hyelteMpztAwnp72A9SuOwKON8D
b/aJswwCqvzW7bEP0lUu6ZJw3Ceb+JpTDuIyzwdcqfGvNAyJTE0iw+TsMZa6q3G3
smTjqszqgklumc8ZLMQME0VpFJuQcATfs4U4SIlQQ751iUqs/x6PqmRXc0R9o9Q1
WuaSMOf+Xd6u9m3OblauMeoLAhKRvu2/40c2SDmuaKw8ZZ+XAdQpM8AMJ3IQA35+
uDt1wGfjnKjBTPVElln8SJfH6F4XegvZRL0JwhXZJA+427tW8OgyLN0dlB6s1cu2
PNHKxVR0YKhIsUWgT9C+AHZArFMqvZ3Fe/isPloaZQ12hDNL/XSvWu/c8WUkhsaK
vxA5BnaYz/LJZHS8/WhBsqlKL7FhPvqhPsWgNncP9DhNWOs+435b/xdFGDWlfG5R
ygnQV7R33P2LQkQv93JemqNRUF9yczDgtnYycoESx6W65MpG8eK31epkzXcNz3jV
Muz3cPxe3r8c7xaagwR+lTDCQ4pY5DUwrWHyvtpxpj/zuYpOLJA2PAoHhtKZBwsb
02NLQGYUXZkCpfm3Kah1FXTYXH0D8GQ0TiJ0Xqmv/3TrFGgHhgKUo91uA/e/Cm//
67q+sFvjlXUVVflU2t67CO8VRrYaGzGT73VusIvl2A2Y+aow+NNpU+J7osNT2jCM
QJQos76ceap6mqaDeMtf1OKHWzNRFviGVsFh6j7WCI7eYtTvweJpIUxrYnaoSrc5
RUtpf5NEYnvsXeGAS/bLItYaHJh57Iu3mxQPDyETranaXYRgFVnJOQ9JDgnB/z5q
u6TY955vIjaFjlmc9eXOWVEPDu3UhIeIfwPkYrMov0U1JPqzn4z69HWuCH29XkEZ
4ydouADQYxkz1MG05rscK86UEDkgpUMTkiPs2L5X4kUVt0fC+AnRIiyG8M1Cy16F
o6wJZ4r/ufb8JluaYZuoCCOsuLLIgvFwDQHikhVvh7YXgbXgUg+xhfKzepe+w46q
eXnqGf4BXJ46+b25H65L8AaERq04v/nNTG5L464d8EnHWSe8l0V2yFMjRsaSd++8
hGqap9qTG9KSjwPc8yGAJbomoMYoerRSbtH7v01zCH+1IUBw6STkjkBxGZJvTHVP
7YfSwjAC7pF9vFOdEs+obRyLtU9h0sUVPnUzunbp48edfs0ya4bBl5EX//WaK1Bf
6ZgfHaq7GvOc3+iO+oomdiiVCWjt0/LBeX+9791YnsVuablBOzSxvKYdFkY1Nloy
uhT800CkoJiMQhTk5MhrAbek68d7ZyZtj26D2df9AuOFlTVTnRKbG+3QFhzk/Vn+
grBRAQ5K4Bu/jIIN/ccUVsqHTnh8oh8Wt5V3FW083tSH1k46THZFQnZXPq8emLR7
9f67SadllV/amnPlHONX4VlCMUa/yKGSMFkN2uHrfalze56/jCSF7jXEwFLA5sMJ
auIgNvpfMk8mIAiKRIUFWZPvbdH9EVQIoY4K0ji2ZHWgUFsZQ/tUBZbTUb4elGr7
iUjgJXgSMOBbe2dekEIbQ5PXDtd6w8wxCM8jdppz2dviq9tm39MXNBOcTvULQkpn
0TtiWOayZ+e5dHzdIlP+o5BSZPODITOObRabcxdQTEvQAnnpVLlv56/lAUl2ipx8
vFPcd01SRT1Cc6ijfBkTYObhgFMpl6m2qxLGtt0emzac2v40S76tgN4ycJU5A2Ob
fx+bNbB3Kf6q9DWgj6tEaLNfkxLHNDxbYu0gubZQc1qcwb90IIDRVqMZ6820CX3n
fBsfylBiAuhZ8syxZpBxUu6UnN7icjeXVJ8IZYTVOJdV1RuCD/SKR8M2TMA8kgfO
/BNr1N0NvMVa6BgrgCtZCVejDOyo632gJrWPi6Xve4OGIkCBwaiLvQA2RyGTbTxs
gR7UaMHF7c5JQwAct/fQtqP+xRBG/E8OfLBus73G/yJDzVjGL8O7FujSeUSOaILf
9RG/ZBhF3CnxuKiQDaWfxcSJjml/4LMg6vWlH6P0jyvRnKyLZh1RdqAxKafzM+QM
rHvYiDXAZ5B4AkGXMVzUh68Yrj0/8JBpOFSUJ3sxvsoObSiUUXVa325gwr1PjeqC
sBLqZzLf/j24cmSZWm7P/YqxwJKM4nTq+AosgxsxtdQjIWo7dgB0QXCeP6txgLiC
Q2EcnNw9gOU/Feln1fbFK0ERSAFxW8IPOq1aCfOv/TVVmqbXLABbOT/1cPBwJ50r
xNpS8Q5Oib470pRHl+1CKli9cXgqobBBS/ma2lWNhyyBzp1flqoX8LR20Og377i3
dDRzafrmf2nifNZ+CMebOgwBocZHigGdlh1vghp5D3JEt5dDpWtsCLfPQKNek5RT
m/2N+2Udu3J+XHcSBIHBQmH+9kdj0aGeG23sp2OYhiAa3mwLAF3imQvKsyFx+gWI
LkslqmHFhxQ7OcVFCEfHsVIU/4nJut98cs4uYosJ+Q9ZlUHOr08Jqhz3X0eBcDO5
qLu2kLCvLFzvh6bl4+8NiqKy4lpeaIP3W2iogz6lGCJa6KXAvVRpR3wCZXr73xdX
XDQ2xOkItJXQMlVj8njkjBSIbND8l2xOBMugSaafvxYXVeHts9Hrs/vQgbDo12b5
6Ojsb36Q/qnNRBK9nUiUFBHKZsELeUginyNA6IcRf+jBBGtDH3QkHMPX37ynIIZD
FntHtVhWklVkKJ0+sXyEdjWQG6vqZ+Ei3Vajc/NQVhmoPAzf++5FX8xD/CGO2OPT
5BwG7z3EgMzjTg8pLyERQcvFvzXF1mnL0scFvxTEYBFKkH1pdO+gmwDmps1H83zv
drLdMf+7xQm6htkpgMCmEOFnWDKL3fKO7DGCGxWyDB6EjvsHqoY+o1BV+tmiwvdL
hCWllTFFFWpN0jbQeE489GxOcYZQOcyW4rDtg62iic4=
`protect END_PROTECTED
