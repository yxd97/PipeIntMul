`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9oJRDDn3af6QLC+l3piBVRuNp5RhkHbe2cYyP0OGeh2IwttqY9CVH5SWrD+R9Kq1
am/VkRHtv9M/HZUPsycEILlwqPIwmDcMKh7PgxUFW5MA6woLdBnoHki6Miqf510H
VFCkN6CY4pvPQgVFa39UslXr4jGYG1wpVCiirl/L+I4fpsq0kHWhjQ2hwm5xWVzN
AtCvh0chkU4zy5WfbiVQWtfAu2FJhgSbT7dExOc3qujK3R9JBYLq/7Wp5u/O9DS9
u0jBdQ0q+7Zngt/xwILk4hjFG2pQ+pcLWBoCkvzzdby7g4uLXriYcJ9mQ+qhjNXI
Au/bVY/dXqAXe3MgBH3Z7G6P9ct1shIMAbwuI3Lx1Q+Lew9nlHuycpDEJjrwnPoI
O3Ay4+0J4kSXw/ZGsiJuOOkwu6G8PhgjUGGR23KWx3/xK9pjRuzBY36JkavopUa8
QwmFGFjBtMJj89b56af3Rl6UOyJjO2zx5xzJSlr4KGb0f/1hflERdZPwBJPkgb5r
YX2XhUkOLmhlepfbL9KNsihy7boJnd1lcxKu3fuAqZqSHQI1y1yrzXhboBW6TxoG
qT4xB3LqMKjPwxfjlRH6CDE+5g15X9xJeMova7DDb4yzPB6XTgF3ZnzywPvvpUhY
JhThy2ufOvkHiJdK29vpRlXd1RRNnrq2V5CWy4bLl4MV1iIxwCoJdN0Al32Tm/Ms
3+KXCquUHdCNhNM/QGKznoxG4jls1+DgItonnUJkbmN86dn4w6CBr4BtemoKQcO6
50KoXF3CtmnrlvZByuDq2rUYpjOZ/8hfZNcUIPSbPifBwl3XwHVKFK8YUaPZA3bV
`protect END_PROTECTED
