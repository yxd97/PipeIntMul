`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
97hCgTIZk6USytM8QjDsionIC1cWyMiNDkR/RDesvkzfM76pSxRY+/dR05WT1l3q
UWZBHmZ3YHVhAfq+0HOIVsZ0LQnYyDxKy4W56ydACAA4IfOgJyztiJ2qf5JmalqV
wFF6JOtWEHbAx7shAyYvHJe2A1Gdex8e02v3yTmAozN6Hm05QAaj932Rf/XPGpHT
2IaOkP3dwE8x4lDZZY2m4zUMyX+fuxyDbjvYBhNKfOH1I+fTfVMOSms5HEX2jUAU
LInNZdXCy8tFvfasXH0vUx80CuV1dlriQFmnj/LlsI1qCwLDddoW8K0Cknnlo3hW
m8C+C3mt+IVl8dFVXFs70BxN+LqEPzJsmAUJhUZeoaPm0/wK2pKE/W/mSGTKDjvy
1S3kSKdogzByv5lzqVU073Ct3QG/bW0TUQO3HYgy0bwv26DfZnW3dqqYtn3zozNB
klchWB2nmrZNqCTMAixfjD7+BXpsDETidSYsY9u0NFi0TtONdhzsm/KQtOUloWKB
/tb0WRECaMVE+4o4Ca7hfkebXMGUv43aRrQsQiyZLLmTa3cI+WsQbLtEBwZgrejg
BupOvPhza4Irpmv2HEshHp413DjjdIEikYQLUxvt3lNBGCZ8cUETxNJVGVm0ckPE
q2LzWlOLdJaMy+4vD8cSxqyeze0TecECTulVZ1J2vzTRx+db8ov3Gc/XmaWgU+g5
yigCaU34UgKBBr5kVHR4IB7RMzw1tHcpgYNsMN52N/DWp+co0/QhYVAF0UnbEvm1
jD7drm2qpYp07jJO22sKUE7i3OSU0xmpT9VC0L6wsFJCeQBQb1zuJJ3GSJ+UzYtW
yBnM6DXCTxMLADKaC9Ln7470XyuqRvElcY5QwSP1ETnXSC0QsbtbU68i7FbJMOSK
71IzVM9nVryfnMRaSvoXtBI9nrIzBhb6c2L5NJLSbLK39FydISiiBjTklcZ+t+Sy
q3uCzL4e7a+OknZeWV0qPGjlt2pq0r+RBWqKQD/kUaTWH3DdTgiQeUjAge5coTyt
PXAmvZTGBrn+ZwFuQvj8k+K4nlBYDLD9obD1Xgz1IXPVFQ26UwmGB6TD5DPQaiCl
XJK/9pMICTnriUn7EdimXS+Gq2op5/LY+6LIjP7Dw6Hbqp/8epE0x1B1VLt4kjCa
E05Q8YUjZX43IbiITXgqdft23FCNWwLDfYdnJOxYCbjqDemSGbZKOXegnK2eMw3O
d1+qmPEy1MKEg5jMqgD9hSb9+bVpCMSleGYar8Gs+Cj42HUgeyk/McjZ9oX+h9aV
CwGTzABS+ezt3D7D73KsnNvfWQjt9e9Wzq2AUHyxR1kAtmqaSuxdbErwTWrC06z3
`protect END_PROTECTED
