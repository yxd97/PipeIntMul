`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U4ugYwcAfhiDZd63yai1elLNBygDbJwDEP8pgay1cexFSH6vVf54yIezW06a+ME1
TEYjHva1lnlKMFHVwph0OAcn8piyYjOTPPjRSgEpuVBEM0HWxiVaKbA5puhrW4BA
6Wbq8EHiK+YfEbiZyYlH50m5K0bnql+Bh+4jG0mLjDX9pgLLPcCmuraJMl2WbkJP
f8IFx9sZ9CLXho2FDhLWO6axMXZbpzFe2PLDSLHDK7ynwcF4eXgRAzE8iJ8eSV9M
P84J7pmjSycdjaQCiF6lrc3lGrKrkXqcmfKd46M7d/q8LY960YMoBT9HMaHL6Q51
xg5KJQrEqOfRbWvCGPQrNLqfI2CGA+hntk8r+TvAQX0Gd/JhPyFQG/mfAI+L0D2t
kboavl7bXhEmsASzb0e5hKFqw1/dwUiZ0xwMg+aqXPgWJWeWWU9eA9V61gYRUx/e
6V+VVYDE0CsTk/UFGiTWFYQ1VC/NZsKZmZAX1lOFdpmEKgcfJRNi1HGIC+2Yx6lU
MQ2f/q078jYAjrQ4oa+bTf4npa+vfwZQOj3/CoP/ZMozULpi635VmwY0O42xkFDP
tXpcO/xszEeNuLe/bNjBx5GlTePGjlZRuxCMWQOijPrIa+z/0DS26n976qS1Cpo2
7S50SgV0uCQcPdk+2vazKWkW37PpevHlpxSkfOt+Xe/U3YX6yfzjslsK19ch6/64
tk8GeXMl0MXDH644EvloQEDnKC9Mmc32IHnb4i9olsMYJLEROKC20+4XXhyAzGUl
NExsNKpXaZXkE8x7Imo01Io9QTiqyDE47rrWFnTqnZah+gTow0kfg6mPNwUl1bqU
DfcX11oxErlGc7R6qC4CKE4IuNVxPj8qDmSTTfLbQ63GGqWZujM90JEMO55KBjC3
q/T7QWPQNlKmg62i+ZoEekXaicsBae5izRJ/mIzOpWo0m+hTrHgUgOGRCgDuZP6n
pmI225u50BkPbAH6ZfgHV5I7VpVBy7SsAHoq8wgTsePMHd6dGFKuxnlPzU4PcLV/
IW8T8r08rMbTqwzPmrtP3KWPpQ4QtbLFBiYhnE1MaP6jTFz6BQJvLvqHrZpF5ws0
7X8iaclWk1uy9XkfjrFSvDnpYRIZw1ddnF4ZbAyL7BCgg9/2K9WaTAP+cTFOIYR3
KetN3Yl6s0glIleAXDKt7kHIH1pomzgIPTn99Y6rDiWjmKhZPxexbM+8EDhhXTZl
72tmWrotZDNMI2AVF0cyeY2v1uiinJJztRX5m/zymFWt5KKCs3edbcGgJsQ4k8vh
34TN9fIzDVZj+xExRj/YoTj71vdcOgPdnnHn1jbAAfcBb06YtTpiVee6T+EOulHj
7R7430jcaTrvDLxUXRB+zMBOk1h4YVvrn78FGtbqN3Q+p1OKjU00/Wl0Kinsu0zf
rlHSlenBHUcSkQvO6ZmEoXSWImuy9bCrhJnCxQ+qZoiZ6KWs91HfLNkX61t9PZIi
XihWDzgw2Jzoy8LgN7Uap7nxMhK0kzUVsxTMg5IAiLLRO53UWLb+JH6awovysKoN
MzDgD4ZwYxKYI9Q51WmPB2EhuVrsfZQPb+qYAT6PzqONci8ypce5YTkoTWgZtZq7
/7yhbeur92lQfa7w8fBu8naOkBG5K6d9IyYOVXzlHqWfBScoQAh0Niqudkhax/EB
gmWKC72SxSXOgGJAQlGVRgAtsMMc/EawAONllE9m8cSC8oPktCM3njPqTYqRXQF9
1Y3Orn7qwwubbj0NJrUGlokGg0usxcVDx/PQ5C2nfAfoFoBHtpq06rn0J6wcpJFy
zDZ0Zk6RcwuoqgsIxU2tZVU8csJzL/l+JAO+VmbTlccvNVNPmdVeof/99QhTeTQn
6zfYvQ4YRbZcpbtiU7I1gJEn6j0EIeC+uVkViMRVNxTJek3x3TBLUz5ahjgmw4c1
wv3BPmbuqSo60NzgswxibEAMqGxV8vYzcIR0DmdO6dc53UOQ1zk/Eq2L5IPmV8Qk
87GthICmsy/wl9Y4CyA2BEdhBNgvymMfFQkwqGrgjrkWLn6Ji8/rTRJmdw53Rn9F
BW2D6Lsptx7eWiWZg3RkduUDUXTs1xPlZdTGGZN6EjQpyEUn4BKx35Phbgp0Vrn4
vHBMuL1xQxjUHJAwUwOE2lT4rYY10uwEK74EoEmMkrizwIL4xzAemyUpeW8Hkxpz
p1pnz+Pzx3E665s+lGPLqQ5m9+ziM6F//7Fu3SGL2+nJFlhw8EbN1fSPr/F5N+RH
gfWDxraky6XLLbYjSxy1vHGWhTiCnFlLTovJsx+RBYXikZGNGzOQGQC038eSADLq
WqHbbKd+5brs2w8JSKnGiysd36Z+gn0ithpqwRt4yxwIc6nDApPnlrozYUSZSAn2
OQI2P9HAS/medvzBoEi41INTylb0H50L4B0IbdN0sXRiFjw7DV9tcqtpwXiYLeIs
TKc1FuKEWdUzR27ds0Lr2dPnIMwlL0t/cPuO+fDXYjY99cddEphL1en+Q1JvBJ/c
ModsANALaozQ6WlQRFxqGkavW4iChF7qvD7sx5qXrCd3wlRDfAVuEWC7bp7FDELc
dG22DWpIUWQ+nyLzA3/wO+I5g2Qtyiyxr4bOlfs7G8ss6yzMbcuSVwiKkdgLo6t0
vJ39H1GZDyijnQ07yLbtUWxH8bOOYYtyDKbCwoJ/H6cXcEYMiuFMqTd5W8ezox0X
ZNm/pDjX9JIBuJDElyhg/FfUhByKCJxuyL7xUEsVKCE4WjfPA6t4VjcZ0WAxPZau
8ycnFhd7S73C6+XLmQFHaIMjhqSG3OpBITsFjkRdL/56S8ELXBGU+LSflMdRuD3U
82ML2bisDiVDHHGOSr0aLj/XeMivofo2VjISfxi5WNaRt/AYt4BNGOZGqp6JpBoa
oW3GbwHcO6qpepFKgYj54O2bNvCQc71VcPSmcC39aB89Mv98pA7J2qV9Tj9QJlR2
noH0A1uDZ7pOycIuKMgdRQ+GQCrgg7bWkF7poqVwRKvNe1MUEj8ejqigC8qP5zGW
zS6XqMXr4TFyDd72vG58msgVTIcvpKDicrFrtjF0cP79sxRrqlMdkS9Uc96RHQLU
A1935t05EQ2zwrA6oHMItw3N0Q7+EeIs5j9Z87+teW5P/0pDPvAOxulI0x5exNN+
lmwa4Ud/HuWrpWVa28fnC+Dr5k3oSYGzQqBQSP1CFODx/ESOUlpD3dxf8Lf2NOyg
gP8CtCJ4fhM88LW4FTzpZzo01aF+mwaob5rp89JWGF1yb8LqRw/FvmVQ15T6b9M4
Fe0EmwzHQXCSgNM7t1m+fnKKNJppJPaseM2ZmcB22Dm8/83PmdjGy8+SfGO+a3sb
d0+Cl/I/1oyEqQWYKWykcf6wbVkIG6BKdYqPazy3KgnBc4b3BlvwAfIq4pE3vVlK
iXQ4jGhNoG09BbjMhg6XZNOHWhmm0BHjMPPURJtoaP/R+cCNLyBpLuO/ZssEa4FX
8ky8UxezH3fzIHF0aaL8Q57I90MF4NBIv52qdGCCbDXS5ulUTI2nS354e+Pjpm/N
KqEttIqEGdUzkSyyh+Jyp0LQDsIu27SYE0F65PrQkmIwXECN+O5+DL1seBxv5kfQ
wpUjXAES9erapJqSjV6kg6AKIo+tKyAX2mePhXsQI+qORwxpa7RQuWHX95vgydHN
i8g/eVxQ4/MR7RHaLiylGw3TYr0r76FaYPsR3U0oKJnfCmzHbScJTHPj6ScVgLGf
15OtmiMlmqlyDUxM93ym3HUdAaYQ0R/PShf1/WE9YorBdNDQFwU2eaj5EPah6MNy
9j6K3CIeXLnS80/x8d/biBlUxoyyylMUMlztuwiXpNx+0lCdOjz0X3Jcyi66EfNL
Wgt/pH1/yEFVGP3lEkfUqUvrviAP4m1iQYEFRQ9e0ySxkwh5LO6y7Ww9Q+JCMzS9
A8A4EuNA8Eeji0hyYt93IsAVTJm+2sTyl/FeAbcb+ffINj0c6TghLZrRFXjqaIJX
PYnr5MjcNTL21+ZFrwphPqh3bhWTWNyTTwZQZDmz5PDAgCq8MjobSZ3pFnjLeOXH
OShnQrpzhRh2Jh4bfgrYuT0iH8bv9jelNLxy/VNiXOR3q3m0iVRuIyQXmuflJs7S
CZwH+hZGBnNX1RD1wsfKKjJZ7E295dvbysnlZOeJPAw+kxXRubr14sD2T8KWLs0U
n1eJL7YJ9ReK0a8JAlOBxa132jyT7NMUhSNBLm5knkSEHFcRrxuBXdVdl4fqwc8E
PILo4HKGw9R/M8tCy2gvP91EPIbsNhGGijouxVUqNZLR1R8aiExHAcwx+OyRw4Jq
DcNr18XNnkruIqoXcMBe8WSqn5EMNc1hlyOVJteDXK1TPBxs02gM/0GdlW6mJ0f+
F8953HQeuviYMWXQF3MHGNptlmCpM+tA4wdlATzIkauTvym3vUvr3iYMFoa783tT
X5WYT4qKjnR/ZilRAPzQu8oADnVsKSZh/ycHf+250On9gF+7EK6D7ztpI8MFToD+
db192p9esREZfkQmxgClU2LAkKz9PkLuR4vwqGLRJb93qPSVNO+S4pm3L8Ef66t8
xd9/rYFcwHg/nyaWhGgUfU4oXkH1wtodEykCiw3Ey9ZyO7sO4xJr+tRnXoDm7IC1
mQbcv+bYd50bBhBYyqARz590JM3IQxkWtQ9YHW8sk0h1Am6TzczZY7c6DGkuXkfp
gafbQqNDdjaISEX4FzFaV53FgRCQfgxoD5SPuKrApbwXs0dgKpmeeGqc83nCTdyG
SLGzDxwN/dOJ3R8BigAQxCCLG1mM1Y3rtiHmRENdgUf2JFkjC0jKmFugsXPiEoQC
47XQAgbJUDns1OafUzv08aDACjqzDuOowk1eSg//OHFrSKImplxhzYP/j0WHy0mF
Jn/i3P46DrpN74tfyEo41HmJ0uJ8OEeODR98lkAlG7VhkKqX/fvWBAQK41k/CfEK
v4z/e/EM1Necohu6lmXbwJ67HebuSnXPGrNvdixpLyl38JePj6enHEW/xRtLwZDS
xNSjc0Y4GWF9otBOjAdZZSPk+YmtSVN0snOSBMFwkx+VatsQQoTHc0qbnEYKhmH8
u1DwM9RkMv5QTe3ZpvPLXAJog9EWRZTQO80QSDgO9cWKGtZk+W/WSNP64onjuq/e
rfkbsCzimN4XbM1w+ognaSXPSEwTeJDIigWkD4df02CUzr+vJLoJObZWyJOym1gr
Rt1zmKwQKyRBvvOYqq8+lKhyIsqZIIVwUpT5ht0j3MOYkX89JCtC+ZxTd81x/MGF
sIe3eMZyOdbdgmeCQNhDXLYpgKdeou62dX++6zbcQ2BB+EtE+C4BHB6dg7HQbuLx
+ZdWouWh1UaYB/yRssTB6KyPrkv2lqZDEvVvFB/C/MAlz1sRtUAuwaicmULWj0ET
X6iy6lSDCIEDw5/bbDHexJM6DAmJQISms8w4zx56+5Xe+M8UbSQ+/MM98F4UE1hG
1BkUbUXcOwPVYgFOIdstYKRZgWCCOv95Rauzqjl7BELOfLw3WYwQFSNiyjJ30yN6
xhOVvYoCHPoXQ56Qj7JyZSD4PNP3kTuchToXhQZHLSIX/vVsjEuIo0TOG6JJ0Hgx
F+G210BkvHNp27gbCZP/oiOmN22c4Qu34xxU5gn8p/9rRqyrZXt9HbEeA/4B4p1f
mcj+nnpGDwFcyD2+JUuln3UruBtsYiuQXOZPNWfXzxezYJFc/TNgx2XVwpsW91BD
pEZArv1aTOnODOT8KE/T399x0rYiUIcUnEqmaPz2ZpBgR8Q6e0PX4XVbmPK5YSWF
IF6TgzQ5ONEhH+dXhTGa4V3ZCr84f4OnhGrTF7bAdqE7guP1zdboz88OEG/dWIU0
Bp1NW8mpSlk/AnwkvYzKQj9DGDuq3M0dOhj0cTtRR9R/c5cF1Rndp83Z3TeILguF
9Y7CkhmQml6AB6PVtTJBpNjMWZgly1KhB/cHxR0GKIdSo1uDcDV+90/8o5IK5tEy
X0Z8buuvvBoPqZz5jTwJQGOUSrjU67JIqcIQ2L5t19Z/ghwquZMNSGdVqaNQedst
y/Nt5S4xoWykDQXNk57M0YN9WTJYn8VVc+DGHvoQBD/WKBg4npsLGzP/yKvIzKwo
Uy9U03WltTg9cia0AVFIPtr4ZxXFyY5cu/Oc5VVi3aGYHgswBHwzzJ063JueQndE
52BIHW3VM2B4nvkAYxF3sH3EH7oQ39G6Sm+euo0lqQ2fzDl8wzgXVaAbq4IeEtek
N126uJ6sR44UGHN+VIkV5RlwB39kd4ltgrwxKPtHSKmJ6s4bPFXUsmjMTW9icvxE
0ztO1haG/cXi4e4TZSVq9RPnCQFpJfuQU7qWAIYXYFpW+FB/mU+rNJ1aespZPdhF
96qgsDOgfE1+53MD7ZMYw2FL7lENZ+mL8W8vL2GPJN9eU8bv5o/jfCjxeyCn8YCM
qragIPY454/8FZxr/ieAyRQ5JjwqFcagWRLZXLdZcFypuVvhn07eQ74+Bz1GogSF
VtaMkL5adpnJ2ZXBJz/QLvcuw5U9+qvBN02afz3aq4tM1tOzPYiNYzXDv/ZBUNRy
4O4MZrJdmE/lKgaWu4Agmj2EaHXA1tdO9z7R56wOnJVn6JUjlXrZv/uG/boe6o11
HPjEulbadNz9NpltFMp21Vap1ORI+VWePzl76pY3zlKR8e6DgKg0KYihm2Q0Cntj
p8hYULIDPuhby4K1Nqw4hCn7RhmJ7NyutYd7Hy7V/ba9iTVWheH6xSnN+tIHH1lG
wDtgNSa/N2TcHNqjbb2DL2xuSNF1M1kId07uLHBd/8bvIAjO7ATXwKahSrTiJ+Zn
CLcTp6gSUJXhWiARSvIdvZTHcPeC5Z2SKlYn7E05I/W//Zy1yWVB1FN9IOPuBpjI
xkscqV16VbvthpS/RHKfnHcPolRzgl+1SNWKsZKphJ+IdCHb4/XGVB1NW/337jH5
vp1xojPoLBU6geAwQTP6kN2k/PFg5pQmP3sdTmv6NToamFybgMtIWLg1UNDLfNk3
hNWNEbD8DGfyX+uYuzi2R/FRz+6F4qb55eTxLoCslFjwNqHh7dXS44adXw3uVgjN
+ZToxAMB+u6skPHTR6gMPHcokS1Z8IPNvGjNYksaBAq9f8pHr46RuI1skW8wxQ4l
J/832xEQIlxUZMvUKNiE6suWmVa2cP7b1FiUGuJX4jRmopjAl4T3i5+Zmdd1FKe4
ecQ5uagFY3V0o4SsZUrUjRb3+pCde2O0X4SzMdZUTJrUOxQGUMFJFvI+kQGm+ohZ
SVOCC+Hkv9JhjQmNMEs8U903hYGh8TIHNHJGV8V9ihhYXIjIQOAcs6HmW9H++koM
YmWFGstBMs4ZVYtie/mBYLHVVjjH8jI1OYiT1tGs56f4QYWZkRYya+UDlJhczDeR
stRUxoSDLu1CqXsJ6VRADmxqr3nj1ooELCiI6sPkmQxDff677+a5139Yq2FUDrxm
pqTQaYJzlU7Mp6A5OYLdPQKgaD+90Mtg5SugW5hhfo0s8Bw6sHOYC2kgu+Eeas8r
kcpb4Gp+iNEyTMh/pY1XmVQ+dhAFX28MoxG9pTSpb80xcIgwEREgWFt3xhsBi19P
AWXxwv1Jueb42WiimdFmRDaOaK9HoT/F83x7haN19IbDSK35fTO1atrGKYPj83K8
M5vMfVwoQ1pc7OGqDTgdY6Gmqwnmb2dqNyWnJWi3ZHIGd70ue7mGFyEdoXWsa9pk
ZDFVpjlMJDYKd41asp/EmL3l93TMycl2yl23zeDamtFKTSpNbrzZw49ZiqbrQywW
zAjgdisKSiTFVaxBHEJ7CeFFeh2h13HNdCuf+RE4Ihr0OnxrcdSBztAa0d9B4ThW
n0tJCMihBF8fiHGSjQVBUj2PcckYdQzY0CFdfc09ULCjQG7p50YljCHqOHcmwp+Q
aHLd5E5OrRYONzaerAvcOt9zSmTSvqkl261rfP+OlojoeraV5xN0NJmUS441xCOc
VflPkydsA8IcMzRfW/uIY4gR0wi+DdTM+FJ8aZEJHy8Hncehm6O3QlkJHESQjBMN
LyvdDG+/g6BsIclzS15Nf480uC81IXitjAYXDV6z6yLuDEU1Xmp+VZpgr5+LqHJW
CpIemstEJbHkzQ9OjX4UBDJd94KSEvdUbw24Klpf82AyCIKT3U0Qk4cB++mMqvh8
v5fTjzanSFNO2hCLEJvWqMUo2D7/h82PyO3jIMqlA0Z1yyW0GkS0ueJ3Vos9oX+Y
cibWQiN+D7muKeGhLSWyDbzG+8JTN84tnZs4gKcPoum2Eo6o8Fb1D77e+ba7y+DX
QubLa4LQs1o8FZ26ViCUNgzmrch+RM23NICIfQfneDiTuDfD7qWAc73lx9mkQV/H
5ZVICqdu9dghId+sZzrYMH0xaSMDN4NUz8sIRUq8HsViqd+7+b6ZfjfoECtas5io
S/ll6Y8HTp+izaeZ+iuxNgEihcpTO4/6ByU+3u62Z8N26vSwC1YqUWSAXgaV4q2z
5jq0+scrigpb11R9TJfg3RFxQaKfF1Zhr+cgfa/gzhxEgdcd6EamPMmIRhptB7JJ
+C6twxC5b3/DIKqfcUYQ5minmJBUuIMLCuETgXJK8Ne2jRzxrfrd1EC/600Om1kS
FAXASs3yGNMo8kk7gglny4fkBefUr3Gzh+trcYrFbHJ6ink7WXtNXvggDIDfovcT
Kk3kVWJYoxn+DX1iRBSDFUsXxa6Z9icnLdnMtBlsZsb4SmF1KaUCnTWOAjmAYjk/
IpTEBqdZsDAtv1b/Pvlj/NLA6IerOFvqHXsSkc2kNSrDnK8sgmcs154E8NBBB/Tz
82GVs761jjp7CZ6EqTJx47z3y4k1gVzSLHfvTY8E8eBHvJeSVWikOsgxKtqp8qXa
1LoZ2QDcXEtb/AJ5SuMQXKAd7Idf5/Lb0peQhw28Ng8ke4OIMiDJTRtxcZapRnkQ
P8ekvQcr0/QrCdNChpMxrvTTNdJ8OsSK8sTa9JuL8h+h1EcMf/rT26qtN/iAUOLL
nEUooGWVXoLuheVOIngYLX0LRGqiD8dLciImoQDecB4U2JHAtqgv5nw7Xuj3k3Du
W46QNXBj2TPmGg6XIwJ2ImadP6n1+eRYhdeHNjaj5Z4GjEAFc762irAhztW9A7y5
02bHFcOAXzl4Bhkw7seDm6+5qqX4QIaJx2eyPHCHXL85xIoxDI+WvpLFXLD5Llmp
ZDEB0In1krAaXwjvRqNIdLhpbe1mmX+XELPl0TIDyVGW+nXdo26kXNjvOalk0tOK
EglaeoMGMr+vD2GRIgup9J35f0lKJAgAAop1lHtBDltvou9cN0alRRTn0EqxhISH
KawvEUd8ZUcN7YVIJ8Pr6tf+NAe/NdYn4CL1HIqHQpuAkzFf5ba0UNVczeh9SeZx
oY35PToyFA1lMKYWfoAcN1WQ2Qe5QkrO9bg4uuq/EE9e7AJEYoqOJ5229OhICznw
gUdKAiLqfQRqub6owP7f38yn72tQhAXo7eekUBUc5l+S8Bkmx3w0CuGvXxbrmQl4
i2MMz7Bb9JYUygYEQs5MpSi+G7JC0LuvKyJUXmGYQRopJjGeQnY/8Cq97r3yc9MA
r0HvnN1Y96WZ1Sp2am6hT/px5xTl53VuAvnPQzd4yc7VsNjBePUitoTFZKTzPDhE
hF63AiMXCY/Z5fq1lvlCn1cQmXY4z+SDBa8gUDwCoZDjF7g23ukRfJxEnvbmbzeP
ggaOjIgfWopCOzEq8sjFomPkLS20kWCsukixsmIJxL2oUwXovmJLQPTy1dC6PuEK
mkeceW7rRgyzYxzv+oiBASmk9gu+XfeQBTALPj5IR57In4gOO5tU/SWRtHWdKCqQ
cVvq20iSsuLgDPIniq72f0PW+QnaxRKWrVMnT5LKvi5coPCJmkNYdonJO8r0fvNN
NLRM5o2a0lfZ5fKJfFM4Qvxddx7QYaCnd/pQs+bqEDsZUUc1dN3D3wEWArjXJI2U
fpXZG9i5W3Cr+/XkgY0UYciaeJ+oVHibCuJ04Iu3r8/CFsWIOwQU9sVn6bIdPS+E
RMUj7NqSonZC1wcnniEVlaBXT7gaR8gRPT329ELNPJWCRnnreQgBQ0xFIu5u5R/3
RS2MSnKeOEgpSbQGyz0SmmO7yYM+XoWlGPpy7tfWRPqzZLiy7aAO0PFcN0pQUDxQ
UOwVpMcNrp22cQtPrug6YCGRD9umHNAdc9ykYqZ7uUkwYkp5p68xOfsPNtFyn5/E
83NSdC/XGIhwJp3Qb4MUwXTYLcjPR2ABYDVdsFnl0Gl6eBmX3BQHzBcaGQnRxdXh
1OE7Tctm2NOxOoG33BxRf9ZldMwZr1QBRQSrDidqHi8MHA5fZIGTlUA1XsyF5xFW
LzBk3gfzuujOocydoz7XkF03wl7cjHqK/pVGB4+GpqiM5vaaQHM2+cja4WMSzNAY
uPLQR0kgUiFJskJPBA9xQ4/9xXzAYJOj56Y+z/YHxF/Yfvd9I4MIx10JqL2DsIVH
4GfhdQ4J3eefwrZhs8tvPFwvIvCDMARL+32fkIngmGfK1hsb1/9TvDKOsgj0cx7N
qmu4obycA09T6zLgy3nBrk+3Emx/HOzBbKwxaWl19GQOQImx0h4q0g31WGz/PQyc
rtHX9m0ZTS/P3r+2WYHX6mOCFCQmGmpE6kNWGSmiQpKNxlDY1AQpKPrNiqBZxJu2
EgXK3aY0PSzJWFoGOeCAmhnEI5qgnYdwAFijL0bNL+Y81UtIO0HgKGUYcZsbM3ha
uaJ7bIdafVcVcxTyBVhOEMGM98oSIpiRjErGC45omGOewwcJ4Q5S+F/HuAudIJ09
V4omOp3CT9jVxgWVSz4tBttt7Oeza83IfuzKT/aYU18OTzRbMlgI4Yyd2ywRtWfS
d0tIJBPPkJHaQGzzXlgLHbOdOSBK/5k22vh+36i8YECNThvQRiaGT/fRo3VnhHFm
6myayA8gQ4SfbqVqIAQlJQYqJCKQTdBgSvFnhOikSlGv0PKkLA8h68ylEEKsLNwA
Bjumq1roJgibbvqYKO2UuLN9xZbUwDVWGcXYCVZphaEoBKgVbLJj8YXSExlFtfLD
c7mmNL5jL0fUD8WJ5heMTP76dsTKWfueYP6QQRg5SsdLpevEgsyx1lEz4FdZ0VKE
8v2sB4KBeyo7hTGfTgpBgu3xClAeQg9tjKEgJk20Lc3Zsvi2ga/aeffo8w+BmlW+
11eyt6F05E9Ynvj9GD3iOLRxNi0LUDILSFHZTxMHHOtd4sNSL/DfcCHBOTYgt8aH
32+FWS3ExcCs9TFISTipDFOTkAbz9huICd4tt3LtSgljaqd5aoHhibV5IDWF4Wrj
dWYk3MY9435AEMcc40pKP+4ddssS7xVp+E1ba4ZhzMisYUgwRYuP1nyTiE2opwV+
5X4pmLz+XjCO41ISKTS/wZ3l0mjPm70NDIFRHBCLIoHFFJeJiG/A7yXbEkDQtfl0
bENulcDQSRrf/ZjDz0qURTMgU8O6mydI09zORovo7yEy+7WHZXYupspFMynxh+gG
VShe40L2RgFirRDtY8Is8foNbcdyInnjiYBKSWzinL+2hj01kIg+FmIm3MdEvJvt
px9hr5rQsEvaCmT/vL6zuDeFwGa2ojf02n/naLLbnj2Sm5NJViaXuH8AjBgktaH7
PlDPPLyNnI179UUa0iwh3y5da3g+l3BKOlQ2zKkGx5kgEkNrd2j0qSSciG5AKMLK
ppYH5VGBNTqL4u0Ain6CyqYqHVJAfAqcjIALfsPyWaqo9NRQ3MUg5qw+OoW0x0+P
f2+Zum8XPVBXaCcc671UxOgXQ6XRgb4fv7nq97cALSeb4K8yILInbPny/clX9FeW
jssdSzoqFy66oSSoWTs9U/kCwkw59+TPmcqC+5DR9INAISiE6X7yajUhfTRqTdEl
REiqbHU5epOUgn7c45XWjpUs3ItS7+PWKFTDp59GusM6iTdKL988ye4l6ZmVopuz
UCcGii8RR707Zz0W8OmJOlqd80jLflwRC63qi6zrlxhMCDVB5TKWEz5wfBL+raqO
vVOqmcTOnlJAIw6vJLN4q8w9FYFIGgmFyUgQhScAtZ3PKwtpwxn5a2QwlVvHdSjO
fe79Mg1hEZ+SjLAcOA+Vh5zXbxY+mu9WP1A067micDgVTbXOrx0urQiQZ8zDkpfY
KumKWMi/UbrdfJXe2oRbsFVOoxOu5r/hhWj/x4HN44+atUrdlXMskW1u23E7UVaC
PFYymEfnGKw8+KOqSvrf+FZWgD6M49TpDzbGUASWPc6wLQq8pO433wjiV8SEbh0N
cKsjVFkmCD5AdnBFqdQbXsilLslLoUa4Kqmttget3cVia6GPI6aNUOMNO+qCg/8o
YZAESO4LcYkAnOZs95Z3muq/Cn5iYpF/qvxstWmtq+tKvl9CxNovGa/tcTSOQDU0
wcMctSA4ab3er+z58wApiRwy6wQNxwDj7EmEUB2B2k44Pug+ChdzQQ71K+Yd/R9m
utl+JJ5dTV5bdr5ao8wz9yN7TdWGiKvFqWNHCHWqZfuXomlb5tvZCNi93NUjqBeK
nNMq5+aRdepxMezNFdKtwBsTjn24TNN8QDKX2zAQFn3L4UqwXhxRroYgdMKB8N7N
uh0eL0AADHRTeua+jxYX7aA9mdyymPHp3e/jiFS1TSjYxuVvZqpHTxUVz0AL/RO2
YCzzUIIHH5SPSJX92Dtm7IK23SvMM8jlcI/h1bj4n0ZysDEDSxnNT1LeLXGY/+2z
qJ0KWAvUcv5blLQcvutKHyjHySQnREdSJyHMaZW30gClJHJurb9dmAqZXf7TpvU3
U/AogCkVqfgPeq0LqaYJOmJElfe2hGbMQwS7tyzuiX/hhZM/fPm4m7r8MbGLJhTp
hoOxXq1gvB+3iYOStegXEMPEfZFFdvyDgsRM+G+3uG1Js/FGOYZh/jCecV+g7Oyz
6yLeAC1TkVuT1rOqx87BNGMTXl9fXH9qcnoRr56nyNUwD2KGwdpsjan3oGcrDgiw
E6OjiCdC2WRuI6Hs+GtAftP9bx4f+naCFNUvplpfxf0mtTnlIdM4XLAPPzBT2OGE
iqwF9prPe2xz879lZE65eHUBVSVtzebP4Q/SRxSauux4fAERsiaExpsGhlvCPUuM
G8+E83d4grBB8vHKORR1DwVOPIowUDp+q4HR58/+4BClAhtfesJxzYJfktuFzL3c
nG4elHzp0mtmapddIeDBtnJJWdUv3LmD3uJsrkvnL6bSn+TEq1guA9O8rktNT3VT
OEVevHVqCsR+FwV6qSpXbzj0QXeFA7jw53JQaRaCEdqYYMDbzGweV5OQOvqKIVk3
XWUjXrcVtPmPTPH88ymTO6L/Jf/XSalBmlQrnPWHuK/biKOvdqJOxgzzz1HpFSUF
jPvuhvVPNscDdzjvjrM6Qks2jrpr8ELX7WwI1vKzH1W+95ZzSZU3ow1Sa1bUCYOg
n96fMr5tSYbVOwsYLBJWhqMpgaunY9aeweUoUSnpuoORutS1ROhDAAPQSX+QiYq8
EWQA+aWaJxybBYL22c0iEHPLnr/5CmLe6PKOwNsY/M6kCnGS7h2p0GJ8H0GEx3Eg
C35aC9cGdwh/03gzZArVEmtx+p60nPCO5JpyqDIc2VavLrw1x2YTYxSRSs9aadSZ
qhHbYdVwv2zE5Hhk4clUxf2shlQUgLPX4CaBeLPVNm/38TGwTGhqhoF9f3pmcsd/
u8f2UfD9V++1c7KPSA/xoWOl3e6HeI9oOg3StTOf5VaDQRk0UNs+jAW9+roxaG8J
iQuNC9aNei+cIQrKcsexhfABr2o/8khhRX3LGMzMXaPQ721hIPKtUooIKss/6Xry
aDcxnyfBkcr2wArhgqyIZvGm6XchkFzP6/LTeOmocl/NbuZuJL1OT/jIq76YUaTV
aByhRV6YWYAH9RgXvgLx2B6UK/KNFTBO6eFjWzrRy1WdxWIcZee4I5U9XH7DsMHf
ZkflGSphyQ8mm0ViI3nW8H7lPYBDIw5Xl4qOGhhbb9AtGcbMMyvZ5CT7ZPEFwllJ
6jiCykSR8D1GQhq3YyaRQrCojf0ygcSpXgg3Q5Prarsv3gTUTFl9qEWCezaBuDwO
tcKZBinAesxwsQ0DuSHiWJg7ludrcEKTtvI8Ripu7LLQgo1pH7o6s77P4rQM65B9
yOAMmuzbdqpSOPuwiQ6F3Ihdt948xnoJjGlrvIKfKSqdwKSnU0Ui862uMW+9GJFm
mz+HvmAFpNvcwIfosBa+RJ6QFPnT1fBh2rkX+w5+rTcKAvdfSgqhWSM10DSSOcs6
KWB3WIWZVnwgrGBpEJKPXjQeIX9o3Di0iIR4ktyd/KmGR0WEvkHu3BOs0ZacwSwG
hlJj1RpzyW81yLHWff/PjXoyUDhD1nJV7D8PnWkW65OpNYzLNXzUe0xq7vpeeCqP
0DBXUQNvkJ2W64CKPIdf1OtMN9IspuDVjzlkiGrG4xqesq6XR5pVVW/mbxony7yK
Z2idE/mJH6eges3MmZ21nSFm/D23jdzV1OIVS33dkPw4kQWT6Hj6Azr7V/d0897S
wm2qE6OSS1i5XsUaWeMMnUBGn/7BFHeFHFAGtWduSqipq5MNA9G/V7ZVcz/K8BVE
MvC0igmdBN0E7pkWYLmDtWk1B+kmiroRgLcd0RZN4fj2nB4pdl9dB8cKj3DwrIFh
sRuput5GxGOS0m25FAbBhr6Cz8MpgvL2qwwwQxczcm358AKhFSEwT/FvrXTUMrPa
juXA1OaYAAw2V/u+q1/FmFCB7WxZ4nCKgk6KxIl7J5NmoJdzgVhD+A9IEtSQ0/n5
3Vb3sNnVyj5pN3qQPZ58y73iV+OJeW9Kg7M17vJjMH7gGrk+oYZhivAxEcfCnoWi
wq/bjSfQ6h8L0pC6IN504H4LkC0UbtnWFSlqg0Hh9K9a+GO4lcfxpxjU//n9OdDg
NKqDFrxKuQq6MNm1NN0eRY5hPG425ydbS1BOEs0ahKne0cTRojDH7Spra0ybbhza
YiqUJ+l/CUMeGzwrnPPiH6H5nIi1iNBrkHNWRy5aABnUrHTghN1YoyjcmEjZOX/s
gxDWTk4LTVNPPUnzY2PlYJa9UNGSc+v2eVZUQ81wU0AyBgR+gF5EQw1mdENrhHyQ
rYFhx2W9vD+v+r4zto2h59bghqRZj3qs04rAJn4m+2xRGlM5PtT68GYSMyOe4U5W
2OVgcbDzbkrsj6CtBv0MWG5FIXofppDe44E1wpKzAXBFhrMoqYBqrovYomnGXQct
P5KqEL0wwm+F2H3uMlpYF54C418jJ1u3WM529oMPPovKEEgc+CBAX07kk+xwDHkl
tLkxQjuIduAut35aMz0PK9d0cfGABTdIUGO9LQjyUtwmgzAZYgkFi2UaFXso/TxS
3UFRUHYgu4RhlcPTxnyspFqASizmtGlwh+PgkSK42qi9yr8q7TWnecEmIY6x8tAp
pcXTdRJ1cCw73MmpI2YIFBRTvHMguezfxSwxJUn1I1qG5o7kpsINfHmnKgUFeV1D
G8G+UvyZNdNpPQS0EmvhJXPHNNRSEXjoT0PqzchDgj8bV941nm9zC21ULo+zcKfr
2VIXT5o9YOO+JA5CSjmPI6JRVCxQuzcVX6wTlCGezLezh3V2lyiUpAEVgciJZv8G
w/NHFGDr4NeMchpNS8rPqPJeM92hO4bNSjjMdPHE1TssiH6Xz45d9dQ/OPDqVblg
CrZvvHo+rxLSXexpoN0ePgpdVpwx5F5NM9OSz0J78QP/K61akWS5jKpNihcufNCe
tN60ve6hRhoLmWDrv3hjUvLpCe1g3I1SPTcEK8XyhHfA/fPQ9mUYCBotzo4t3R1p
GItXyCnkcCOV+X9Q8R4+UmjQrKgu3Onp7G/kfz4/zF4mV50dKaqbrDCSwph7h2SK
eaumzzH1I0gVqBWycJPdTuxmmvgnG9FnAmFxBm9vUDsOU1kd4JgNCJU/iOiwF8zs
lSaTiVzrC76Oo6naAEErUGuZ/7CV/HvKa1cvsyhTNFWJl7cPxB/zMdXZsN8UC7hM
vMyCadqtCVTopMJickEYrOVCXoj3uYZz2OP/iFS03UBN0kBuSPG1Gqm0v0zRyC8O
c0lF7lTjphhTtBWHuL6hmeKKkZ3PMpGVu6j6uxjEb8ZkcVYhaxa77weg96qUslOU
0IABue1DCHcXRmad3B/T9lYvALhp6IBrXnNWLilAiKHoS6pblldHnCfBXyoagRcZ
dIO8xZEo9NNt3D66wk9+N/41qi0IV5XMKHV8tT+S4vrQV/yoP3p3Li/hTl0oH4Rg
dKcJdx714vw471yJaeWJetmi83cRwt8MncNoDEHVBzeZqFgATp3LBeJLxWq47maJ
axoZMfAclbN2axpS0nBLVaXDxWqEShcx6r9T36xFbDlBHKP0Ap3yU/MZs1UPxu81
kGvSdi5PQMwdfiBYpZAjDt2fHXogDMwbZg1n/aEVpbt1I8DYj9SZoLveKWOpMNas
Vn25VwPsCSL+Baiuic8LvUbZKz9ziZHXSqqg9kcdv+iHrcournAvl/DOo81EhCNm
yu05bzvPq9BFto6TTYUzgJScUGwj+JqiDpBXFK9pxG0paYgU5Oym+3dnLTcJB+hg
dhX0oapOVuYZWmr7UuIixS5GVAg2yTNhzTflA2jyFxlftdnti6rryUwA8VLO6xue
PZ0N3cgS9/m6IWjMAwObHwio5gnr6Y6vZDxDxNUXni2ROMxJ2xP9xcF6Ziybw24U
5ShpwjMhYLaNEO/WiHa6udrhqFkx599yNQ/2J3GxYWD1WKQSNYLYt/w2RFYTtTw9
ocU9Y6l8v+rgNsWSp2EneC9yqvCsEechJwW1dIWepC3o4WSMbith8KyBADeCxICt
B2+GEhrQOInrqwGzILHS9sxcLjDqhJ23+RUkvjFb1/0vnxjDbhzqPEMnHDOhQMaY
qSN666omGtVu1NOF0byLDRn8Lj+BMXLQWFTMh64jdlyzMN8pDjUmTiiJvMugCbq9
wHQSl0aB/8ODlZ8VWMalCJUi5JeV9ri0cgSyb81qRcSi05I09Uxdx9GXXQaGAEPh
c/CypehiwrILzxn8EQHOtgLJTs1cJisld+QAhoVYJ1eLvImzXrVrqFlOZZ8up19g
0TaLfj5wbkszQl4EsP9MbYMJGN60lGg2dJmsdYpuG2ssvnspAfp78Jshm0CIE1S7
UcO+zywix0gnE8oefgpkI/CKOUBwjCSWVwan0WaxZS23UkmtBSgyBzNhAW54m8j2
vppMxP2Q9Cqj24rKAg2u65/6vhbLp26Nzyz67DFmRSga1bTc4saGruN0tucXC1ep
2RaJcxnzZvEjDwXV2HGqMCIksvCpssrBlCvjKGpuIhEpAFdVw6b+mdQQP+JQJ2mR
dZrX8K2tt0GNsaMtNk1WJ1ZMoy6z/OW2ohbz/jlLu923//dJIPcBz1v+28J7DgoU
JAbupovRGQS3eEH0SDCoaxKZZBNDFa+DPaIU916QOUws6s+/M0av2idP9ZIi3ntt
caY8Wg4PLnOC+1cAaso2dxXejrlTu9ZAN+m2qX7Jo75hMzHw+Mlyft3DfMQu915u
27ZTx7Zns0cTsGlOpWd7mjXv4akvs9Dhcf7WmIfoTqyv7kI9B5+YOcG4aWBOinIt
erNWSt7ZQBrz8NYqWawcvtcCtAoq52KoHDpnxeiPh8bfYQrGJWn/VDBBOUZcdjQN
U3GLvK9mRntfXHwxt6YT3XhL37BYCaIWzsus0PGOn0Q0KUBWrjAZO2S3l4GURCFK
ZLaQERZmerhGCmD+O92akqFvfT72Lz2GHDuR73BIn+ryv5wCHkAfm3CfubMJjA66
Z1Co3jeah6CTm15b6nKstCTE7+cD6irkInSqxIehTTpvMj9LVp8avif/RypY/zcP
dp3+uRQhTLKBp5z5oGkmPE54K7pf4Jz4w4YiGZmJ+6pRFbvVTTYEbla21LuRQgQK
VJ4N+TLbL5BWw1EkbxyWqFXXTPliuP0cd7nuNfyb01jPh3Qy4yjrU1v29E2M7+gO
a0RVkA2D5iiSZR7ujviCeASHnDRk+LiVxgaxcLt6eMjCmXCUjkN82tO4oUgwyE3O
idZmKoMdCgw8JW3vt8uca6gXr+KoTE/EcgTlq8F5+Kteyo/HrjnhsEOXdYpnt9xQ
U7bClLh6THbO1muE9UkNpS9Ln5PR0WxfVugWi8iR4zKC3eZVuxtDeTHNkb5qOMWo
XU0keVcdPdrjA9mNw5wxHTCGGZAnWR2Eer+JtX7zqJQ1RnCQ3x+J040VWGF5teVj
V/jYRnH+m6MEvn2vdqLVXv/Xw1KIu1mAyjnNDOU3uRYo61hYWtyw5qKrkEC3Er7t
47ZIpLPSLGGgDFfFiQkN7KP98JHi5Cj2gLMbOHMLh+1ot3vPkAqRPTV5BtnVpKJs
apA0BG4YqnqY24wPgSBmLYGkBhUUsSDjIW1gRWzckm1aKIIB1z+zIgrv5Jh9s+kC
nh5ZKRAyd7iYi79F1pKAz0OZzuF/vUQ5JdOEmfDKzuQs9NJqzNnr7LDX2q5k11bU
iBNgOi/qnNQUsgBIVxfEU/gSpGshB2FtTLDsphd96sHfSIbAZlVHSvEhDLkalHtH
r5ccyHOcVtYBe15NhrYMteQMDXwR65BhpGRNh5ISQ1YkbtGPKFo0dM6BcpCPou6f
CmLoVlWgkofJBmclzjWsqLRaXSmYxzknaMyXedVQuxGyTNVDVd6wpE0YUwAOOBaR
rJAz1b5WG0Ek0lX8kXj9bDdPLBtnWzdZpKYHzcuQFJAZEgn+9Wk+0Ko3IKAK5TK/
ipNKmF9eULjW6OFvdCS99qfaa0DObVKS1jDAcEqMzTcZU3joCgstoniyLdbo6zaK
9panp+1LZ3lka1MPtMM0jo/ZTzvgEMh0NiyiqFD8NLrtrFU+JhgDoAl647EetG6k
z4ZpbslWe/UfkVaOI2Bv3fg1l346GLjo4E0h/PRwbqk2UCMa7Hx1KTyYCsOQf0gh
CwbjcQo4P96A5xPJIzAy6uHChqxwFru5LifcypYbqc8ck5pcUl+b7eMPm4xD4lQO
/xNtEREup06IzxrZAtZivfXu/B8YCHZPgL521Dx13j2weNeNWV8+CFlgzpc2d02N
GXsum3bhRV8IMeTDFVskVhca3JncNwsxNSxinFgelphkHftGAF8gGy69AXEbhpnB
kSaieqWzQ0AfDKF8ki1j05FsVfL1C59+N4m3YF6glzoRXSXsPBXoastA8vfsobvR
j2ohfp5fDYs51+j2AaLtY5aaD4cMkEsjnBYclrqK/zIG/2yfGhAhg0PVNw+3qx/S
PatPvcqPg+wGeIzh7d48PhQus9nNFSnmwPxO75jpYCUHi3kuuebsZRngQABpeC9E
AEp//sHdyo/VRssIKlOsq7fxcqCuv8ZQAHVCoRd6fUGta+sOj1kdxBMbUq+SVrvv
cOpcebXzr4CzB6lONYJHY1Zis/jio4G2p3aJXzOujgKaw4fc7fXyjB3cwpNho9II
4jTn3hlp/sQQfPV1T0UjHsrzcHL4kdJfwD0lBmm1Q3Ye4F4Ybfqh27EOVLVQjsNO
vpHyUbWMDommKAWmpQZYrS2s/HixEKHAhzxoJ1DKAZkbR0WcSx77Zsp5Sk8YXnb7
6rMhrTv0Rpu2/jOwmDsQ8XVoLYspWyrXDn3fGrYhZ9Ybu6AYFpsLifLNS8mWUA/G
zvMZwy3ceoHwPkjCQhSSL3PZmxLc81i0KIl0F271oe5K9j40DzpdQ7nWlL+7VXmq
iyySUjXDzVwQ16nrL8BDk05q5w20crlR9eErAQJ6QKyitlq4zZ1BP3ITu3cIRyMi
Fx9EaB3eQrCvy0NDKtuUC/xyCKpBBcsnv/usZKD8GkwOfvkDNmEHesSd/dbfYoLj
UEpyNw3oRa8T/nuiNP9lRPfLtHo1G3vBax0oYkg5INHPNn7DdX3Bf688XQNlEYiT
omoZ5FLlEm5yTfVFFC5EHEJRUkE9ijxaYSTa3AAzX84bOcLIdt6jRUHkw9bgrCp0
sPvRFY9leJcjYwdTk5bNHFjoVtoG5Q2SNNhnBFzLjXP3hEgX7+Wx+6Nap1tF/Rm8
rlnyA4xttseKkw1oG0xN/0rTgBKTfDhFpGbCtb8KVMAHvJ0/UyRroM7N9BcNoDWg
yk7R/hoHm1MXdr/he0e9vGcu4SxIcNW6f2gj01Qtjs07qqLUJzPHH4LD3dSWu0t3
vu4EkII+a8ujpweNUDyWO+eMNlFWQA9Q1Slf+A8b7d8KLoc6fYCMP6A2+8ildPd+
9EvP/8jgue6z4rx0ynlPpKd8+aI0l0xRWqTCM+986g6xZbLGnERGR92yDQGOMuSo
6QTrVXIhnC6utF6UGWF/00tojWBybAFzQs+CLMt/3PyaWQyPkz0rnwKPd7AkZGju
JnU3cFCC1NkyzBJ6t+ULe2sDZA1NagFUOCewrO71NhDarkouyeI93ZAOZkGPntT7
hjPgb/bKKA/mu8zvEaylz0/89QNkbkXfmJbR6u5BixZAv21huhNOffcskAXBEAlx
shadKzkqkpz6baBsFQ1sjRv7Hb8PLih2RkwwtiQZEyV4QdZ40GO8MxVIejyXtYcU
Vx9AtP4J0X+acpO2KtPtsCs9nkM1eD2YUQiD10x3XcufbXuSrXGBsR3UPp/rv6eR
TTXoJb2+xGyBGinYpnWRDSts6J2pa4H+gGUuZ0HlKhQno3S72DDkA92i9XBYljHE
xMT5GEJ4bwfq+5Z1vlpuiDMEpnTy7xCLUr9HEbk9Kl0owdD0XO+oT5oP1Q1t0hlk
jIz41YLQW6DMwhNcmt/szE5717JgFj7g9ODjnFt+ipef8kZ0gV3XWUmEmdFD37UV
8+6i6mEna401ZV+U6/S/QPc+UD3HPsc+0IYiSp/cKLdMy0QVQ07ZZhJL9fjb9hVL
PWLav/RCekn9obkHK1KAfwNgkaW05z0CO6iGCIvT5Y0oRVU5CBByk8btdXZk/uqg
cASXFA4/6GuprOudp95mtC6EPthSWvhzNpN8mZ4Hrg/LwixpL/xPxqvhuTp8/aSN
ZZc4lV6oZ9bxWdgjlZ4/AZavUFJyR/CasxmjI69ohHwfFAAQtDX10Bz/1v9jeY+f
RLmtI6AU6b/dOsyWtcAaPTeTPviJORWUqOXwiBuqirFbzwnDONIYqb/6ZnTn13/B
InAXJ6ebhFR0iPRWeCdL6rfFq51fRXSSUtuCHfok+j8yfX1SXrfWzmmQd8ZHdxIF
zzu1/Qsvf65g9950M6TJW/skNjWekVNKsD3VE6vqz8DS6X8xkKaivanFMw31ch1V
GfZGkUNBqlSYLWfV+JxRn8MBoe4nYdlMJ56TrmWX8t9x7yM8r5Js3Ul7s6ygAK/p
/EGiIVmtCfvl70Ic0nPv1Usk8T4fmkem3/py10LcFxWnFx4pNTRqFoKLy/ZwKX0d
XS7GUkEWMnbgdPIqWHRFEbf2TNxp/63upXpxeZOzjOv9CVZbxfVH6r5SP55jWLlU
0W5la0BRVBjy1IHujw/BMk2VuY3Ze2Em1rLGmMNo9rO+Z+9JwJNzgTB9lIp8Y3pz
D9/9Lt9T81JA4mmJRmwWRXR87X8pc9XqJFxryvL4HaMoDejBEyOnwjT15W2A6t8j
mHVt+Uygequ0zdZXz7NnI85JoNuWa7t8IREPC1CrWWxSnCEZkA+7NifHihzFv541
8NtsealsBrsox/nn0fklHdcW8q5rCs2Wjfe2baSnDuBX6qHygyFCSDU8llFZ1Zpp
ngY6rpTc/2arV0PVeSX+/fcRrje4cFkxosSMxBpfER9wEOXet7GsT3qIoLETpRee
WUsuIRbYOywqsQzOcPYJdPAHKdEqg9OYQDqrSDwSa77JQFmpGyCzlhFGu4iLVRiu
8km0nlc4o5FjVzLGRPOApT9iXpOsga0nPcr62VHEC0O076HLOsvGFQ+OUVAx4Re8
kAk96LS6rYlRrtip4PnBZTaH9EOri7XjuXpxiFDziehj6dGuHJtSZtAVihTBbMoT
TqbgFTjSgraSVhFDdTpcW4GKIcka8BDXUVVA+dZaIHxeoieLhbSflhqOPHvsUegJ
sdtduDa7iCFW2NJdw65+Sw5+v6rdCTPrrJMcu9+0YKZXZmmujAaDoJ9E+obDeuzF
7wj3k1bguQBMAiHv7Hr/YP1m5ATX49Z+PIcjPHhUxRXqfnEIn5Ggdia2nyHqgZ6z
1niLOh6JGR4AFBpqOWsKRTB+rbV+6mkA6bJ3cbeVxjlIyPBuwmRTnTHfhW6+gFtW
UOniG8JeIHQcp5nPVk9ghnnOgx1XfBKugPagLg28na643hKU5P9GmEt0zH8QYf1K
5221CUMeoyhS9+nj70AVUIeiEkMSFzZyMfgorjbTYWJF7NP82Dr16+ZH9Eym31I1
KEPg5tEXm8IXnrDMdmSvoMkD6ccnxs9iww8WUB3VhAYJFmwEZPmAvNLJ9e0sGPbk
F28GRkHR1VYDHNrGqyQIaOt1uOsUt+cNGxStWmqRtd6EDrtqMmcyVWf4fL9fzuTU
DSSGqkYC1Jh1Tcze+wP8um4zmCRzawVCDXknGwCUia06YWzqcmFrBBVWtxu/VbV8
EITC33AUft5/Mvkvo8IKU8Bir0s9cY4vCndnRFASybfQ/9tMXiTmbO/8sxlsz/HH
dVuvOmDWEZQtbyZ/bJIKHPrpl7/sFjMxGxDBlW/rqbzxOnfgdC4T+DeOxtQ6mSsy
wG2brZppR8I73ezytCqVWOjODn27sNY9m+v9DhfvtzgYwsJJuJj3rQVNzimqJ1uV
TtWZgpBDdILvCqZ8vBEhfkeVPaq5A9hlpgkCDmxy89Z7tu2z1l0KBmUNon2i7zOo
PzutFxYJnGayev7Rc6gMQ6sSnDUdNW/IXbJjNDv/cM/z8CCINGQfgIMzD+kg4yxg
jYFA3WzJ8B5R3LZjlVdmdTO0/0Q7dAf/y+VMVf/50cihiaxZ4btbolaEQvpYd3+B
EGhFNLbtt+Cs/wckEPehMZQIuMS2pUkdHr2hyF7O/uTYwLAgEGLGeL42XGpunSKL
G3E6DTlpTB0jUmMPwz85NJUh6Z5m9F4MpoomYL17BcnelwTf8lGc9+X/RX8WeAjl
pO7BqRpYczb6TnIchwVhB1nB7Yi/OmmK2L5vi/bp73l5lYcPzqdBPwr7YYu5418K
NgeYiHP1hTeRBAAGeB1BPpqM3omKQk1r7BjAdmSChSMEIaRhL9dz8q9tBeu7PERO
noE6coJnPtsUUOsCHuv11hSoUIMfmaNsYaSugRcfjYMtPhOEEoM9wiQKgq/uz4Nj
DOOkpD2I3hJKbRfddQwlxLMKYQTN78xizGZ79CuBpFCh//5ux+QCeUMxsjmxOCkH
+VS76dl23oF4O0zsFvemVl99aqjMo1eYaYzKUVUmpPRjsKa1/47nF0XmYOkY/sT6
xH8O+si6vtZTZwlx4ujNttNGSGagVF9FsjNpkWI7ohliRpXaOiVJMhRiUpccth4K
JiL+xcSp5RMxWgJ3fWCXH7sYpSeSY5u9cwNNT9AYzkSzFMiXzeRb7sehYoq2tpKL
bApweAeUS9c+tfKMo7ZcOtITJ/UloCCdnmH6Jbw9Ad6swIn+YqIOJaKcaXRFDFED
jePbybzWyWvtoMJT+t7y980pC6g97mc9GEKvOTqa9vRYl+Xf+33mcGczAvRAp33t
PXCH9vp1msMLGzrksLJEl5ncWXYJFKaEhP923xkFj4Feb+u2Q8khXqcRf7/MDikw
P+rSkys4+ojK8MVFRK7EMuNouAckvu8OqJ4xCHMsZlGwxXLW2SNHr5mToRim1k2u
/mW0rYEyLqhkI/RfnKS3y8Eg7jZfehTPpGizBzJr3yfLOToW5XAwm7RqpmdzxZqX
O1sWFcWqs7F+uUFiFon+OJ5BeSuIjUjS2Bs7U4o99MRebEL64VIPtZJtGuMW5v3G
b9GqM+131MJqFOidVWQ2OHrBvreSgeTjVIDqfm8w9HnKw2Pj/qpVoTM778Fjm/mP
0baAbdNB1hSjHTkQdmVcV28/kVbr7ubbzKFiAhgRkjmSFC3JhLs76GTi+LcCef6J
y/1RLenStkMjJnOXUNna8fB1cYvN/7mXMicuWc88KkIhYK3GWEgRzAk9W27rzulI
Qi6vmH26SrAsbdlS4jMfLckqYobtWsJOKuvkbiHAwtiW8nMxMD9T2mt0Ha3BXd4Q
O9vQM2FPGDcRMokQVIXiIbcL+lF35k715AEvANbkK86KatxUvgbRU9XYwwfxqY5v
bzGZ+iKwDKoRApz0KiyMCIlvxQR2DyzgA7jz/GzTBi1b2g3HpuRH3G5BCMKKmwep
411PgDUw1wxQU9QTB3rljlZv2refpLnZ1ujMm6H1PfOgAh6nEkmCZV9uf9t0XpzE
OdgRANTZ+eGKTjOcuTMSV2vD7KqMsgZlCG4voRzluxaNY7ar1nFX2m/uS182m73F
4e/8NAfyu1fEYLe/RubDlLKf/ZP79nF7f4pBExhwy7UXaWSWqTLAuqEcLs0WZJVF
YvFNrUCJTn5bCEHj7ZeNDftnkeYlWAL9Q91Zcgs0nrywWuGHs7Xewq/gsl9alLP8
SguNrk27cBaZqqYmZjEbms5zS/bfJgeOnFjWz0eJb8Qh4Ea5VqoLhGdxslI2ePRK
YwdpqO6pticlgzusOcPyeZzd95hfe/W8nCdXxKESuHS1m6ZGaRAqcz51g7J1a+i1
k5aSGc3AS6BJDz60/8f2EH/ob2/A3CKdHQfzSJtmyod8k/cIPnl3DOU9nhXEyKDC
BpRZeP7NNuP6leIisnY5wdNsq4pN1JxfeYDXcE5CjqjfMNgdIkjgdeyrtlssQF55
2Ac0viaWWqyF0XxV5bzLWtQ01LSKZloV8J2FwwvqDFm6Aadvpz1wt3QoZftX7Rag
ZhTzD2+B/5SuQ5jeWqkwxcTv+M6UrxxZAY65L+PTK/KZWp1gYMXmPwJ2RoB+Y08E
Q0yvj1cKa4MKvz2EUHsUbDmwOoIzrB/xj0rk8QdCFNbspJD/1Dr7hEJD8mOUvypb
8rHzEc7cGSVLgX4PHlWEvEbssGcIamGIuos7Eh1RwjYRSuXq9XTI85AuH89LearS
utow7aR2TlM1Ef9zEDGwEWu/BLD6ZqjoqmWKZ9PtRBZjFLAA+r7kbYg5chK4ao+W
VI3Qt1Y7hiFCNnRbYIkH1ngCUYW8uOG91sAdD7aXY115RcSGopccYm5JgW4aKFIE
amt1je/JMlmq209GjHN4lIQLloqVgrsbU/huTxdGmzKRKpIBA9LyyO047Nd7VuUp
5qryiBRkFfAEYPCFgI1EM1NLb9MieUKCmHYo5eg2XEoamXH0ZGZZsbFMOxhrAChN
nZEUE0xsN1AlJH4YGZnBH0T65Duq5//mwlvZrnhP4bMqZjzfPbRwqnJLYkD83+YF
9C3SLzRjfq80dcWy70SUJgCiAE3atd//6u99zeVfUqvp5o5t2hnbbdC8qFJAUlgS
iEhEy2zPXe4NEhqqEiWbw2l6UhTO8p/5QS7rv0vxNQt2T21Sz+q2niz8bN+Jfe9t
0kxU/Mb2pmXtkEvn4yXTSAHrX9FyOdq3WAafxfAX4/A+47JdWYd5V8hHnAKDlFx6
iLyYCuKHoD30N+qZzxXipsSpm3r6wP5mI62PPjE+UJshejoXfIBe5KWqujo39NW8
SF2OXwWL7HwD4VkowrbaQb3iT7Jsi12jWFrM7eQkIMqML4mIQbEjvY7VFnpuOYof
6ujAHauk85pI48uwAMtaImiNFlo5n3WXqLkWenMkjN8qnkZX0OoRMsuHBJeMPxo5
DK4uLJzjLI94pZUg+N7/cCnMtQWNL3lw5X1cgLF0/Ci1jhp0h5fksqljIwU8Iln4
GJ+Uj1x4tEEDzDu7QOKPBWAqLYTImbi2VfPuWgmh0kpjD9M8guOOlKlOHRb7j2C1
IlmiZCKnPNf5hovpqogca6471nbHw7BVrvkcrWaia3844VpAc/gYQrjNnHMPNebT
TAmbFS69sYrnMK21E1co323+5tk6pC3Mxhmo6/0xVT+hAMdJFB0hdbwjjTfRwQHd
N6reBIrY4dV01EmgsBCM179BJ/6tcw7SCHIAE4NJhBES1Nelo6OUepgbPFf+kwaN
cQ0GNHsSb2Wcxv14TdHuaA76IqgXAf/NzPK0LqI5JbfycVBuAK1D7yj3VG9vQ6d/
9QTLUYw588w4jB9bs/4hMKxfSUOZUtCurApOwc3HAGEEn4uqCvBu3LrQxunnMyYT
kk63av7MFzWGVjPqQBe5RRnrFMydQSjOasoj1M9yovQfttTiw81/VYf8xF51o108
xBDRlbApACZkuC8uPsb0l33vTseHHzZTvJLetZVsFIfUYv3M2eymcBdYrlSbI/AC
JRLTVGiyDTGHL8lxJ7MIlds28Ra/2WqevxJ4ZdGdIGPOTA8qgPYReCoN54bQCsIo
t3mkl8+VXr06PTp40wy5LmP2mzjYSoA9hkCnrmLh+EtvF051lk/hNZeTC5SoitfS
hnpWzgGXq1O2q/LTKYHTN2NKFjitjpCziQz8r39OenLm2FPI2Mp/iWr+iPA8fhpu
cu6U65e3yFVazNS7pisMn8bfIREB1HVx0LoAbbYyNPNPMN3vmj3YMIgBmJP9flyZ
/rRTFkPsa3WaMagRL9FZX6kzBBbWovUX8WyYkA2IIQi7muEBndcCHf8HMLdXNfbq
owdHiI760f0bDZRzL2//UU21ycQap12N20NnKCW/7AqJlz0ES5Nj8evUAPGGzehr
oWwb0ZrB+Wn6Nu/I+ZFU9q0bm2O7C8H1Hw1wN29mx8a5woscsvJy3Kv+Fd+/du+Z
PE+cjWsMwa/qXdZ6vJw7uK8XbHVt9/x8YIK47VFv86f8yNPhrnl8E5X/vLCBk36N
Dm4d7gA6B0pLOO2mf/VYaU/GVC6wh43tOeLxkr45pDcYvlDLMqbCTzbUpTJActtD
z1ypm1vqc5v3bsAZF7aJlBuXVTQy8EgL0pXRw54z3/Yc7RgWpv3qN6dLDBqWDBf9
jsKjKe2jZwBQ2LKW54cDRIEOHjDVM1YqdrWsKvpvuUdjgE+supE6U7IZ3KRLQGYh
gQFB1oWXmZX94ETb1C/u1EmKFIa+X2ebv9D7aU/ZonTWPuv/KbmclU8q0pXXZoFl
HrY5ntrgnrdQrE7A+/hPMqNBYiX8K4KvoMVtQlHcJw+5LBK58R+lKas8JhxMns2P
OLyzIxmpHhh+VcpKq0Ya01a1IPRYp0MNDC08gaMDG/Z5m8dOBpoBi/D3XBFTL8wE
fRmUVQbGUatgvlsqI9Suajf5UgdXTjHb7Xh3R4xBvXKf3n9DXyxtw/fx+W0MQRJ9
U0Fg3N1QYtRBH1Gw8YdflHgDp6Ngk4Iz6hbRN4Sj/D3STAFa4vlRuutkJdWqT42I
Ap0aEsi2go9sDy0+SaLUX0rSBstIEO9yrmIUnJqanYKxr4NpgaTP1eqTa1WMw8MQ
3Lu2s5p89CtEttpTMQ+m7o9ljxLzctobFQrHDCo3lI+NZx5mnBV+sqS4yY2OgKVA
w9nPKcalsn2lv+cZDrcfyr/0GPxG41K48qUSVRQ7XvmDrFaigXUTECEMczXduxOY
58gI3WNq5eug2McT05OtCk+du+JScFQW5a8dbtz83pzD6iy7IAr4wye16P4JIhwz
X0bSnOAGFeCxSm2EMJR6fDX5e8YmdKjntW/J1mElUTJgiThrlJTxtjZb1udoEO43
10eKCspeLHBBPe8rppIUB7Ytw6Z0bT5nHYaECMK5scYYdm+mAhpz69gr26Ov72E2
DWTkqVaGTQFlaYwdlr4f9fMD244sEVyn1/eJq8WMW0WDTFJDjYByrHjpVH7m3Mkk
Cf67eJseoT9er2KKqSTcIvpK0YqtxBMajWLlsva1gk6WTbwa9s2Om6mkkKQQvNO/
zxMTBY/3JfIJJSDUmsqvPgigKYc7VL1w8ffU0XGth3Dn0FpqGRtXeJwuMdIZ4hKE
vOLjF4c0rXChHxaDF0L3WGwYEFQtosE/c0Vm0CbFDjoZjbWt5qh0kXL2foN3RNPD
0Nz9vZPBd2vj3osTSWYXL5+dyxzXpL1i/9ul5Oq75Z/tQ76u8DLGXjFf8Yf61ZUd
lRMm59hb8Y5ARZSw6EgbbE8leIlfeHw6ULmoCaCcwS788fTcROebPd1bWkDABbJM
EzvNRep0+lzENzMMDUqypKM6ClJ0aMTSJy074H7iMZ1oC36GDFOCkwXPs8UXJVT/
T1pws1+GujXa3yxdRj6Z/wMJQfGD1DYMTmufczBRifEk80rhsj4SUlIxiH4940l5
ZawL1wVun/UDlUETDDyfzu+Rc3JmhX+qHThBXH3JAI/d0Ggk9TB00l/bBg9QREg0
Les1Cur2T5aJMs7xbxfu0+cL4NPdLwY7ruLdjUqjuO7ziHFFsPEvvTNNhzXHPGZq
QFGf/k2Ith3u4+PWC6lJWoFt0hsWwTnV6y7TN0tO3EyZOSdq+/q6fBe1TZ+IeQH8
PmWZzObxhp6ZOtllnuuB+Y0zPMohQCFPMzJ2jjt9mrcXZElLM+3xxhpKoyH7kZ0o
FFvVc8J5uV1dbEOlnZv8l6D0kRqW8Y2hMG3Et9Cop+6aA755FeFTwQdACOur4zzH
cFeJiY9mATnX6vZVuRsUKnduVsepT/sc4XFOx5qe5iLW7jC/TKZE8w8mK5XF1hgs
5mQ/2Lht0Elh7nAIQuhiY6DRS7qX8W5XFhmP1Qtpk4k87BxrXHbcqNNw5Pwbl3+q
fTKk+9iyBId8HrTpclC2A1UVsNp3SirjntAa8R+H5Zc+guxO8e+Dt7yW4Owt77rR
H18upzncJuefI5a6SYO207LDkVjuBIn6aLzATqfBq4lAMvyTmL8ijYDIOYVGIYpL
WKoDKuVmemO6FeCra3NO62ne2PBN9gvm7lx6VDPdLVRQgJFk9roN5gmGOAQwxmnJ
9iBySi1c4nWj1KRstQFqF1yUlL/OaVGjoXPQ/8Abcqu6UTY+Q1X1d7BukVi+3Fqo
AAW22ACkghFMbNcJEFJTT4NadNcqDZ6Mb+89R2pfOIzwl0WM/N9S86z7W9c8NDDJ
uCKkg8OI+ojPn3+TQeDkNX+JwKJrfEB9DjAhGZjtUqGL1UpZFrpgkd5Hi+2V9E9d
SfQOTGmPnWzSa6pTghbkACLH+UOb6s+pHA8xrDrZtedQz4BCevSuE8UjKwdPQ4iP
9LeHM4lrPsXmFND24UqHSi+RTIK6YBkRKx65/ck4YHvuLwaQD8N5Deil/geJ+iFB
6fLpCxpGurZ7n67ObSLkK5sIZ71QnsimONmXzQluU5cROjN4IRfv2OAVeVwajNHf
6jjXG9hN5yAvlD1bWn2svaHFhKDhTrbxEncLGBHl5QWoufHRkHOqz09kMw9LeHTe
J80tMF3sq/lQXKEARibWU79suWHupLBs4QgInYAAejQEU6+Q88asoMlaywnz7usl
RhBtKenupBYklQv0Ur+MsOZ/tfzNbOS4oh8podyUTdOuzYelXZTl01MQ6wRWTIa5
Ai/IygjNYLIl41PJNid3QiAPA9KdoL6CKWVKbK1NybN2FXDWJ6mwaSVzqRhqabgz
sWqReCG8TmvOMBCVdDpnI6Dbtg56gC453ca0WuBpwB6IpQm95t8V/iELnyf4Vka0
c2PrFxweWQxTq7CT003lf6ldsDnDgQs+9CYgmCGl+xw2Eqb5i3TmNcdnaWfaHUow
c0Rq6fldpotrgZYUbl7hnpQpRTWfHLaZJ2z+7wK+VbVrEoujxTEgmiiz4iuT4G5M
dcgHRizQ8v/l5aV/ItbnCZVTC59jrkCgSmEEoDCbUgqBdSvWXX8VeLNzfZZtY9Qc
pEyt6IgjpweuxnaptM4aZ+tCuK9G7pNKop6/GloDLHFWqbOQpmYrcNqGsQDcoxcB
+/BkBMrHqfYg7/Pxf/Mn5bd2zaF0G3Az1lCVE+1iRdyjMdZyQUQYh6433EqkfvOx
8t/zfoLCkOLYAboMvqIJYJFkm5VVqgDZ2XGOVZN4DX1dCCRFCD63ys1hofTI4xcF
fZsCukcrLy3P1+4Nn45N4rM1T/8zkVM3qUrYojDaooQgtwFTgo1Lg04jiTQcQ/XT
1CZUpuCdVhCsKmHOdMZ8mueubVSSeXMeL6YQoRbC1hYdbBbLoocXRkDJyjXxC4Vm
w4aH1kNkI3HQFkN3ifthNvoLNXghE2pnMfkJdqyoR9jZho+yPg6XbV4ZXdf1xZX/
mER/wBexRX4NC5MEdeweSbfyMzdvrq/4GcTlOvfLDCEGLXWeP2EEy/xLlynPuLJL
aD1SQi66fJuG/ZuzhLzrDlOv0FCy1Vvo3jnivMmZi8zAzHMbfl+AN6ZEsmWc/D/X
GKajW35VgCaG4Fr9r1PUJduI5nEC5vERBpEn2uwQD5MqkDTsEqHcymLjebStuUEH
v6FvLNOJaISCAkPxwnuCC8Dh9HASM5lWGHgOWy0a+8U0AUe0Z67ZP3405JAzuP5t
tkM+6RFzrq11BKOnRc6ws0bmBpArUzP0kTNRZ4xExgM0f0+fpDjMcJQleMmQUNfY
6Qg82c/Sh2AM1qdwlTr93KMWBgRfbbff/8HsDS/gQcuCakhC7O6+nDeAddK/dHDS
3klQRvte9m7CYhwUhKShisGpDBxJtHcPSRXLi61Kn+TK0PgejMg6vvv709x+zzbQ
CvxlVWTUtbweTV+i9OU1j1zVFjijYdQ66bJ7rfCaw90TepzeKcS5MUGIS5G5iZ+i
Dvb5INtqzY+N1S57qT6C/wHuw7k3nIPxAiOMn3KoKyVKqmX/AO1V3LuXaU1LLdBs
2yL0hgRx9nfQoTsdaqe3zXiUflCfieCT6NBOqtsMPNwJ/Y1K2KSLJKlJIFhXxXHt
VupeMvosSdTUL3aHgkzdQljyoauOBsDy6Kb/NERNjBpEfNoqW8/HpqOChA12D81e
0XkheyKh7ObjkoMu35fPJPTD4oyma2vZAr9H6zPjPDGElhalCpC5OXnwhehfS/Qi
LbajvLfROrKiLDOgv5s/vieTqCVu7FT+OaWtwmKXmf9vgrpoGS1eC6dadsPsVE0W
ZDM9+60YDkH7H4sRRJd7nJlT+YJPdE+hPH1m1FZQyflqGUwgWYyt0U/u9eSdSt7F
Cl3+G5CMxCOZRlxKucEWWh6gxlZK0RrFiqvhFHBcaGYCbsfcnzBI19YJv2E+n7Km
XT3ZqKCMS7Vd73A9BV6h/Ynv4YbvGGXklZ5MD4kSOIDKHSaFfqAg/f1o4YSnHgrf
Th9VVCySe/hk070qaYPXuANIvCsb7empTTsIIh7qgYhj9XU4BCJ8ZlSnexLIqn92
2h8GRD7A3WJCEstOyAQqLxnv2MStOur38NzvHy9ziOWIkS/tFSaybnP/U2T1VfbS
9fo9NVbcCa7Ebwss0cOGHHauh/TPftvaxzs4zdYtfgCjFHoXRIH/8Z149x4A+ik3
bxSRphxzEZ1ik4iZdOs+mTm9Glo1GjbUfZrYiAeiiDJsp7K9epZvBeE3wbPERdhA
rhahhllPwY/yvOaDG4b3AxyCPiwFSoPbR/qZxqyhoP8wj6boNmiPPgQfCRvCb9Dk
R0rqFNFBkdiiqFVyRWJWNFYbPkyRdlN57/WNTL/33al9QRreDlhLYx/eZxn/w72K
Sc2wxGRgEwKTJbTHgeXoeFxK5h2CyFjNs8tnDFXbZ9DfJjVs1rjqZf6iEd5ZY9L6
gIv5IpdL1iZLFl5MMA1+cJfUSuFUm+dTX8AMD9tnamABy8GzMpHEuFsKkSRIslbP
UxUWbXjAJpZIphTPGDo4LF9qpuR2uzTDx/+Kn6oGXeX+aqsmrXSr1lxO1+ziZXTc
M2GH3nsqkxIen7tXOeg4zkhSREdulCQOOjlalEeB+rBD5fPPGM77nfO6qdAHs9YP
OXAlutvyt2t9SEW+fEWucuJYIJRlZ/htniM6Kq3kl7Kd7VIi1acULHPK88r3R3I7
rrnro/TCvAQ0vX9VFYXFBqF/jbJ7ztUFx0fI+H735SIye2Ez6iEV1UmwqPuXPN2j
W7fZQ0FUVsJUBpuN6FfhlRDF8u7W5Lot9gkzwKEAsxAQ2e8Pyl5ekaYaRZISb6Av
IHmfXUKmToL3YCIxnz3o11/Xg8cYV6ReqbsWIuOAW7xKmI3VgOmDVQlgHbF29VYx
LkJYp+AGRHlTJJpl0teCu/MY3xz4TV+saMsf5uPIgnme8I/0zpUc386KLOcyi/e+
2SYjZqtvU6ufMs8AUWs3bU3S8mDMul4KV3jkcZzsPulIcchjq/DYuEKFam8NUEcQ
eo4+bdE4TtG/8ryY8zwICDKjzPWvrHqajV9mTwnPp16LuPzPyB7ILrVMpRGoUA6U
O/lT2OHNWD12CMX3zX+NxvWMcNHYPo2FJXCQo4zlsFTcXceRBGPuZiBG2fSChnDj
vflOLyOAL4QxhMY+eCHW1APchmi+EZPB08LtiQ4v92di+CW+uc2bVUyAi2taaWDy
UfeJpP3xgAzMpCh0aBRdkWDzs4cgh9eEYbl9Wl+wanvwv7MQs9TMyh6gvSSiI8L3
ioFm/lQS3viOo+3RC7S3HOy7UCf4kaGa6Kttv5vYrqBh+yjbuMgHu7d7pCgeitVV
Nvf4xurE5OaH2w8bYsOIfgyLNIpOu2o1mlZ5g93SSq8AQhQHWottPQ3ECUqld4hB
QC9x4Inf/OU5uzfQKUT4ZfiU9cQdNV5jyZq4lGR/kYmL0DKYtyF/6cByk8b4fs96
icBwY07rFpYxBqfxmuzNCJ4BKXbXXf6pngiuO9ZYNq+WuclPXVL+o7hlU54coC+9
KTDTaBQlPsGnmgFhy7bE8AoOzMGSC6Zwa14VrFGf05MpP4fTmue8sTDFgCyg7NPm
sBCUvMFzy/PWG7M5iUuEG2/jKKG1JvTamvtAIhq+Q6fWwZDJKykINdm8vwvdycwI
xW83nZhjvaXU2XeIeEHHsz3kFvJZhB5j8whh2hJi3+oUoLKdP/XnwGn0wvzu0mM8
1XlA3Ut499WI+x/Xom7GwLqog7AnDFPChChTEhj5QCgchLYVMREIpNxUh7/wECIs
QnC+fR3EMhSFlkg/+a2ylnoTQFSqy7VYz3K5LYYznTi+t5cUtzcdytzLB4VbHcC4
JlVCxiDi4WXLpQCN9cAkByROIaGESsJffbYCBCyU8v/h7NmdQOEZDJZV9e9f/Kjl
gc5Xnv1UAikF0jSv5xNFvpP/5EOjf7DfOBMiZGRHXkVsPVA3HaLfbrVDbC0Lokvj
70wgmYUNk9QevBQRd/QLG5A99CU2PNPiHl4+IKBgchvDazI2uJ6lrTLq951eyqjC
vGDPvTLIHftBwBM0riekppEA0bsPzALDZX3yeCbx7YdBcLixfoPm9o2df1L129qu
n4s3m9f618oEVkVzSHEUN2wqru4CNMlGDn6AGjyPmfuJx2LEDOT9iKW/G9Olw9fy
lmBOhYxxrail4HBemjbusMmVZIXLn91Ap0g6lbBEny2REpvFeBC/ew0VfMYuT3Xm
N12dJ21UQcMlbxTwFPV8Jmg2xInm/LAXWkXhoZmYwMpbDCmfhVJ11hQLkMncpcMv
DSfUlk7wmvBks6flKxLyjnVZ8vLC2FjpUXqrf/688PGZ1wFyMIQ0jphblJWjAo7Z
Gfai/rccYyjkXlIxqnHlSErJSz/a7L8hY12iLxXIARlUVXyy+GE1XYtNsUpS9Cyr
yO5KB+W6vqFfoKtrNUOLGZ0/mSLg/GRloeJuvsW6jPdpuD/W4bJUDtxOCiZDdnxB
oM/kLgDvmR0P95NhbhTMpjEbOEvaq1HMHz1l8mwEWR9m06nBecoJ7Ir4nq95F5m3
2RlvgqHOkiOldDCL834Gc4WdvNZ2NzCU7Z5Rw2W9ABF7d0cEk7lUnT5KAU23uX9W
FvBw4U93PHBBbpujIslSEl7mlFjEWAoGOsv/1c9nDoHZziYhtDcdyKnjzvK1oRVF
olSUg0KFmJ/OU62EbXNqlWiWxarqvGxkmIbv7B0CbWIkgZ6XG4QRJlSid6oD5HTl
VCuRkmKZhwvqWjw6IedfYdTr+t0pXAzfNaDVe2WTSwOgwZ95LPr0770YxKoWF//f
TxjfZAb47h33vKZMb81siyuf9b+MgE8gwFbyVOJK8JEKV6ipJ/eby+ve02RUcPgX
GD8Rp/gHFafOIs7OOfIejtzZnpyHCKc9XlHZWTfAhbYLjhaoo09kgFfwXgG1QDC7
aTWuyk9Mg0Gxt9JhCtAs/ugwyqc5oZGhXICNiv1vOd7wS1yWlX4+FdRu/QfuA/kC
p8MHmVgoqEoXlUoPfstLVtYW8v+wbLErBiwYd2gu4c9NzmQMT4ZwJZ951uf2SJXd
vZX7ZMu+fahB4MFV5mfe5FbDABf5DKEvY5/D0V3EvB118YwDC63UospiWx99x6EN
6kOBDAEMIqhK5bTZgCMjjpXbgf2DynR1B24BPkt2gBZniKjdrrUdbhzw1Qx1dPbz
N4hnt4NDnNlH+vyEb9kDaSRBVFQOHVokwoVtVN2nYmQF12fhAFDW4imFrUl77BPX
eCX/JfXIlNUiKh8FcEq6RL75BQkSlQRA+ofKjT75bJCFcPa2HRAdmqDbeC8dnbxf
MhWNBjJHVTfiqOaORYIrNcuwSNzwwmwdXXuY30KThRSi4gP5mYRpJSv+Q2hZ5sNL
l9d9oVenlWDl/XxtJ4v498nctZVb7hRrNDBCiOwo9bX6iaoP72kpq4pAgbLN6k9L
3OmLG4BRQP8uZW4LbPS8srnhMJwJ5HHOJ83hFFuYy/zJkS6UvFeOT5Bz337u9DYa
t45kNBKkpdZB0rOiiPqP1D5mYexN8v+0K3c1KYkLvuHMSQJTRXx8nSe0UbDmJAmZ
WrU/kfa0v8YcqmiRZdlmUq92m+/IabRBPT032EPSyRwUcD7UDISBaJFNrmYud38g
L7KxSz0WBIOfZOkTYLVV2kD6wMbxAgFkr9RjJQrobq4PsSDgUC2VZftZ6YZpbKFv
lCP4JP09Ve+CqzTfT25x9PvY06M9+ZVEhKfYBPk6ypq3tBqMjNsX8ud0m16V0Yjd
H6D18B73jhRfQSLCf5op5ix2/mvj95dtIMzuzion6NtF1AggIDb+nNhoGrGwEUc7
77xP6nqEciWFYqxkfMeLHR5/20GA4CZE7ckmD33qHwVG3TGG98okkCbIXnAgpiDl
/pzJJJJYRKosj6ieCj1qu44Je+WvH5TyJ4EJw6hi4u3AKptXTDHmkSuWFlkdM1KX
4PzJYDqILuk/4r5wm+vJQtpz+4yIbyg4xg//9sSVDiUyxwDqBk+kyfzf0AyWJSZR
w8B8i4P21yN/tF2I8jGmIcxzVpJX4hZXhZ0Z8OqmrWpN+B69yv5vr+L21AO157ri
zT1dRR76sae2inRJv/P8ZeefXKjiuyuL6QbXuq5LGVQ/jV01d6NZBGf220LDmis1
bZBzj6aViBXRhaPeHFWhZ9jAelb7NWqwhEv6wawJip/xFf96R4MO/M6MJ73OTHoZ
Vhwn2B6o57c5WlHumz4xp+cj/y6YlkW7S5AFU9rYYxKBCKsxo1jc9oSXKXM7Iq9r
THLoT630NRXdnpgBOSyorKiBGUG6IGwW/Hoxen1DUDxDEC+NPlTss8+gotie0gEt
g2TwYW8r9D3VOyEzb+AsQGJobDCdBnDPL/qDKs2iVDpMbHwQG+y4m5ClRmFJsk2A
RGlm8dBvzm5gm3I2Ljk0oJN4d30qMKt3sByp9vc3muDOEPTew710MH/59axKlIpK
HVw1SJkY2PNibs74qOMMzjG7XkueEHOJq97eb2zgxjTI+kIqgGRvJPbJh+QdqNV7
jIYnYJdj2bhDuUXRJB8+BcbTMNlcwRFsp8FDlom0QdZe/mDgNSgFhSjIS5l9yuqt
LhO/QdbRq2nBVy93EVVV5pqp/6N9QjGtjWCZby/mQM1ac46TX4IrV2pMv0TToEWN
JVcL/FqimMz+OVZUherrIxERXt8oe+ktSkaxpX7Mm47cVfZpurvcAVDY84LkEoS4
p3e1zF7tEKillCyP10JGTcGDTOw6eAMRjgkrHvnPRuXJ72cxy+zMHkCj6vFlu0dn
MzDrSIEOiYtDy0fpGGV4zsppkuBvKxVSndRGFaN8mgAjcpg1wMcYSCfGn5nDkPK4
Js+EkC+FkUetm1Hi/lNE3fimtsSoA/E6fJzJUnHD0hhyTBPYKX0nj/DR9sPv2J/4
DxepLvnXBbX4kZOcN1QI7pTglHjD1okKHVjEdpuMOZZLGHVIbRuAvp+8dI8C6kK/
8zn7MqF3EGVH358Xs2Bez8voSG1fcz7/sWXrwG2UaGCmdmiBmiHAnt4L1lqDQ1Qr
YRUzAHg+EaAYsa66QTLaw6tNN2AXU+dPncxX+4T9/yz70o3sJMtpwZwnz4XVRrSK
s5X1tk03dzKPOU8Oztu11TtIoj3lPPW8K265ymST72euSNqKCTTI1CG+9qcXLwrM
+rk/uHgZJ9vyV8ijz7TLYq7OVkLh3lLGomp6Cxzdx1344j2+IJHubENFQNWiXlTh
JbR2Z44fIXRjO3dhbGFdft1hqJmvxc2DXjwTXh8tbonnSpniLS9olsw4Jui4euMc
qR/GYZW6p4sMzeh9Bv7XBSo8vlf4Scj25YVX2JZUaFDqJUUybS1Akxy8MrSEVvZW
6wNnwwhw44V0DLLZWup9Xr9yXhwBfHjtj6HIYknAGrfT9l8kbrNrx89+FEHXjoHw
+rPUvYZi7n7XEleocvS42+ouQ9EgAnQTTIORuOKc65gPKgVSx8qd9Xq6I3YriyKL
Y5PrpyUm9R75XKemZmjH+sL3B6r9YRTD4YNTQcCEdtEQY7yjcetzTGTra8PSu1un
bugRizbacdwabVoTq6heizZQ0EMdHe0NjP2bSCoRV9IV0vSi+YUJjwtJlQltQx1M
Od/zyTTvxSTZTobl+aQRWK0rmWXJzezxm1E5AW+RHSOESBuillQxaCzqIqoLQwFx
4ErJG6vJo7qo6ZWKcpu9Jskb2sNK4Ng3q7HqWSbouLc0mAOYp9K9F7IaMR77c775
+GfrxAE3D4QHPW28M1GRGIu3pMARc+LNt/gffw4qDDIUmQzl/iMZNo8DFLrSAWa1
VljBfXJd3sfAr6/1aSeFaixI1R4fgRq6+cPhf2EnKyglBA9iInmMjqn0Q/6vOcwH
JR99h1par+2QjAf+7k69zqYNgXKyAVq29TXpV2vk6Jql/G8bO23CkPGgM3mx0oKJ
2P46hB6UT21DebKXszbAQxc559YLn0fj2wIbkfOAa5dzZFbccfOGmJ/zw436i7vK
ZVcc0yfDjVcpGYHAzjiH8fUQs0P05TbyikV8MXjSJyXZ2TK+21FFp2hNbtaxV/ca
IQpxv/hZC62eTvH74c9/rD+NH//2qe4PMWZB4XhVseW+D4X/N+hi6yV8zK717Hgn
Uj5PGLmSzw1wpl97XImB2toaf+5aLm6FQDvPXNiws+r+65TG34wvQC7B/AKU+h57
uluzkPZWaNp2FKqaQo8rsp0VFi+ZFF8Z6r2n6eKBgImDlCitA0XHTByhvtoPiiXu
0GPEmLRU9FMUdHvFV7Ajgsk2wbuLotg81Uwm7OA6qBHSEK7w6XEfbDe2OGULdX2S
m60d8gBMGDXomgmEQh0lupZhUxe8kEjBoqFG9eBtHVxxIE7FpTylJ/DU1Bt+Av7k
Rqj640HdgLmnnO31CW6liSzUtttk3d0ox2dcsGuS6TpqBfS7GhteYhW77/cvyLbI
ODD/I2QRvdMmUM1ac4XCdneUoifq9eT53y8l4yIiJv8LG7DOKhez67NPD2x1GaK7
mAK+UG/+V/OAuzkjlKsde9ILpv8mSysatrqH5lsAxU9BtlaR+1iZlcX0VZBhpNPc
cqEaDjYRa1M2sQ3NFnANuauzCb2vbHtsdr60Wgqe/BN1+QV5YXbMSJTTmZN61DyP
USHmOmSRUGMDSJwXphEz6ARv033iwmQYEiyINmWomjHskRK/yyZvAwjq/1iAHFCv
EUADWwpuxKw92vnWyWjBAdwDw2FLSlbXKWT3eXGc5meXar13Pkm5HiAzW40dugoG
d30nZYgOh+oYvaX3UDVix5oGU6doxkUhNC2zFaHskT5+PZ4vekbH66CkBWIV4Ii7
mveoq6L68KLGXQbNyRdl5os1MKLGpx8e6LrFBrUOxw5qszEOfjTmaSo1KrxR4tBq
MyykjVUSxpq5ANHC6E5iS3SR9bX8mZMhwjwKbenG8ypl4VVW/zEe7RbIe2r+sW5M
NwPbBxO6fh0YcuG9zc5ktgVSAe7P7+WbiDymbSrL61yB1j2GSPGwgzD5hgPlkPci
DjS54P7STZiMl0Muo4SG5gOxVMz5kuyr7oqo88q2oHxamYAHFP6qiRsihJlrkuFG
Pi1rKX3p3XBWRncxGQVH5/3N+wDVxg841wqbxbAraub5MrQKqToE9crdpwcvDX3w
BNwWRk98Viu7vXNOSslCZ6ACeg/BVlC+QiDHsCmC/3tOrkgapQbNTh7FoxL8xcdF
q1ZKDV9xTQ5CONiGu8M1q8NP6IVmXxyD7FrktdmshcLTOx+ZGODnzezaRKHVz9WG
qocTCYp1niTGsx6vhKWDuUmatjeJN1H4QTYMouURSnUsGdxK4gWZxseXnT4ljFF7
PbeKUbbEcuyzf5NpnvfFiNlECqnfvsUKybzb27UnqiuWLK21rRA6gHS1hGiBsBHJ
xds3VJJT0qpILDYKc8WzRvrGr0I1wK+mD6188gLBzpGJe3nTDZirEcBG/ZMgJcs4
uySP0z6P32pTW2in7hBRAXU8IPyx8616CIthlliz5FJJk+KTDnuASwcScdCeHohq
xwLnLaGGTAqbsqrg3KSrNDYeA/2qYT2gmM1KlKrSiVoLtt9iJLXapN3YxXKGc5r7
ZeARe8bwl2GzgPCs8+bqAWsKynolo5bCKcSU8mbhy2gOI07LViaoIjijDnm/nlhX
tkuHO1mamvlCaC3DLXI9848m7FWA3REbpULPDXuOnfrQQ3GlLuoIMT4cAZBtkU2a
EytIUd6aIIAT6HZ8QSOp3Nq8i9ZmT9X12cfFjaiQCIGDNC8tNu/iVXX2FnqPE9tx
Qv5lM8uBQAY3hXAFYutqbgAcBeBan86b0qWpTB4hDLErG2CJwG85wmDAyhQItWMf
QVMsE0vsrdD5wbvugVqAswKDGNUFIpWz9c2cOfd3plGNo2zywCaEkKigrWP8SavI
asVohyELljpB6knJTxG47u3zEK0xRxeeERj5lbGs0eicsiz4P+OZ5hiArz6BDlbB
9LoX62HwDZ4O0ycSvapHP3Z+3L3qjXs6mi9wAyhaQz2RyCFmj+ysA2sgg4Z+EfwW
R+N0/DgjshLJdvdj45D/5+3CI4wFBTjFfjNdNAlXboYE+NnuS6JfWFfIxIrHUq5r
5Df0fvbGz1TNNF1KLEbDkSbdgrpnZZ53yyY3Sh6DGKg6Jk1S0feaOcKJcl1dFJ+h
zNOHtNrwbpJEQU8D/gGweK9O/ZC39MdDL2UcDbvqPRUDeYe6N90lA0PQp8w3drOS
6GxS39Kd6QDlKQf17d5aXvvMXZNtYsK7JWrZlSPrZQ5RzQSIJWdDJj9ud6UXMG/x
AzgIjuAqCTEMRtpaMbZnlOn/7DNxUsSlUI8mbZf9/1ZjwZZFANfQf89+7DHjWoqH
Bm+AA0I+DnDKYJ9zpcc544o7CXKb83yoC6CYH4HhCF0W+gd5wqidQc2viWBnl/t9
wHbCQ5VQebKZcRlTrk8ysQFECc/tnqczKPxs2wGE6BOov6aD2uQXanA/VutQTyUW
7XIrtu8j0OpR5hJQ90Sc+KgLD3bvAlLQa4rGlUbwdOapdVPVZiGJ9dtluL317WV5
d1xoJVLQh7poCCHlHUVP2H7X27wv0MifT5UZYEKNysrZ7pXpsQdnP5J0EqiPgdpk
L1lwmh09dYXPvnp/uxnJj+2hHR7lcWZqF1K6gIer48EVFVXUnAtTkEkvTjUx/PJz
v2im/qWIVqDLrYnWE2SpVNi676iF9GWR5WyzCNbqJPIVNgVj8zLBgRo0u25yFnsb
wPeLqqMOR9cW+8GFm7EpWb48f2Had1eRmGD/wqi/RPG+P9mTjRROUr93lN19AMI0
lR3TAHcOiAjFV0LF8YAyuEh8YI8Y+fFKjlizJnjqenu4lSRZ0Uiloh3yDYrQiJv2
Axyrwffe4DrBVEErAshcIz88aX72oRIdq1x+vilwBoopH5CUoAXOGHV2gQY5ZQIX
RMksoYm+6LSGCvlVK/7iVjTLB11d0p9+d5FHb4bNiwGP1yWMn5qvcXn7crVezf1b
UwM99q/TRFzeTArT7aplkzjnSVyWUhbXh9ottWRyaHmbk7BC1UCRycotMe3GnyTI
Jd9s9XHW89yiG286zh4/HH8gA6Lf4P2d7o/c5CZ/RgT7WZF3EWgTlpmrhx624HyH
T6S3az7ESrBPz2YBcGqYrE3+O9kd8JUZSjVHCWRXXS87RMHJwIVCVo3MoMBPAvSv
Pb/Xu+Mth2SxufiG66gUaVIwUrzpEpatQoeb1DU+iotvCvWXi0G66/2+ywlm6wdm
rWEVCU8ggnCmRi+we+D/Dq0Ev7fcN8bjkQzrdyToPvvKxTRO6356WvO0nvH2k0KS
ovI3UuLjA6EpsFBFQWj3wff45McFaBUjWA3/+iITJ9IBavHbk7uHudM0PbTAlyL1
ZTtGL4lWDKdjL5/n90hrr/tjIz9IDahvyjOnvFD8YwIHC2SBcY7L/l4Do4BkxQkp
LbJgMK4uYUuNxA1I8jW39RvgorNhYwQs8euQV4bA24iyQz55sKCKXQG8GfPpjF2l
uf55+glLs5SyZg6HZnqOvKI0hCTLgh71vXRTZ3e7RnwesUAppMrieqZ2uCHyPcyq
NgD0F49P5bmSmF4bzcP41jRZ1h8yku8C6U6JWu3wXK20czj82pwAI5s91WWyhmOH
DlwDP3KfOIFrFR1CALxeBGcpz/y86WACcXn60m1V8u17N7R5RaatTEcyNoa/9+Zq
acGTNhSdLV4P9m5y0biVQTf9bBdwjOPQvi3zOslxG08kLqGsGrdc6aI8swriLUl0
MT0LJHNPQpxxJTsldIw4HMILbZ2hdlTZXEAv6c5d74L7+82RZpPfjUJ6Fx4Sm5qy
V3YxY9us/MIUNdWU54TO4Tr43yIpM5apOmVhhey2RHzDWWNjyV+5yZFdNLfF395Y
2OkMPfZgNsUBA4kDHQn/mzuEOTI85XN6Aac9J9/yzDTrgMx6Wd29M3lCCjEtSqGT
xpduZSiz6XFt3iMsMjuwLQ5BXgEOIKRv6mEXzWvas3BNnPgPbPAt0eUwrJC6FKPI
ITnDlr/H+gkUXKXXBue3pcJkGs8hRIzhAXAv72u/nzMTKouhFAFKqahleYS3PeiI
ziugKDYZJ+aizKQ4TxFxZwlJJPfF0XPFPelgJp5bET0LLz+44gb1Xvyq9bUTjVsJ
8z7JzS5LwKcS9i2uAfoyLcb7wLsZyeMfW1z3QwiLy17EDrYgplvgz25YsbP0YCDV
5XGrt81p/ka/U6KlT4lVIMyEk7wihIIY05adS7A6g406JDPvw2vfg8oV6ybWDHNL
Mc02hhgKuH9MeTfRWRHEGxbPwXW1RI6G2waRpnRNDJpiyUfXmPStB5vZnB9uO8yO
N1nnQteYbsPke4eVDWMBJj40VUYJrFuJhO7ItvxwH1uyVq0nTqXy/vTmKVZFdpJF
4DYg/Oz1vICFhMs5jRTOPDQ/GyVATuokF6M6DFS0sg9vGBSD2C50EkjpKESWkqTU
7Nyv22jnG7gfshtZewNO0gJqDgD6Hz1DX7CBqUk1LrQze/LlzkNzBFmHkh07k1gv
EAbyUlFAmp39mkPhWXeYx28M9NiGfi/9xHagP9OEbPXKxLxTS1LdrLjPRai3veg+
g9LxkCNZ6GEfr9YtnxCWpE5HnNefOz8vDc8Pmh/o3LjmKeH7Jz3l9iTwymDMsEzl
vMl5m7Jt3D0wU73xo6epT8jgibwKuq2r9ofHXI6s8X/xadHfutTFqi/buYff183O
RIpWxdA8O1+J1dowlBcZ4swb9HRVRmgLkqeoAiNrIZEkmF1GY+n6LUQOy2v3kD/z
q+tMrWl+RskVL1LrW5PGUolIPiORinKMskpqYGzCRNIZFw6c1iar5/RzQAXYx11s
m0OL9KjMR9m8eSbV+/LzhREPTFMt2xL4Vbg+zP0W4EPlwhFiUqvMuPkZ+An/eHjr
ZasWnt+RaOn3xwPK/UaPJcPwlExbWOfc7/CsR6NLv0444ZUEVe85S1i2oO+hn8yk
JMPy9WxRyTOITFFXQs390e6q7onsSrl1JU1NHpVw6S+nSMsl7mdWvvX0/hzwwp2A
NHqjLt554J7ItcVQ0SFWdX20PRHrz8iQPPWcmUL4vWPZoKAWHamY+bRP8mZaIR2w
1nbSfiEcEALDdrrFlth7+G0vW5ZYb0f9EGb9oZApfVq1lN6eNec5rURUKxZDSKZp
Ap5fO55flZa2lYRkQTKarNqU5m+HanAVoANco7Wc5oYW45iKbaZflwuFmOvGkdCj
lo91oVEY2KvTMJHOaiXwfWCCNoxqTsmOayUVTNQb7QuLrMIuOk1khf3+yP3csxda
uyeNb2jZ2wDNCiMOWjo3w5vmiNzJ3bZBo7HosyNXFJaRXxJxJJ3NP7wNH1+OsccT
hFMAoPoUKAQI/hAvh3zHmEFgpJ3r3SJqaAhD5EMV9kCs6mANGVBB8GN1jHVzNjS2
Ae69oBJTBQnnyIeZzPZrqf4U3VFQtQROnYPwf2cR0e5o4solvj6ltV/lojt+hix1
gNfaMjbYgn4qHv+iiarWBNieKY4DByzDXKGtR6sqLFoD63isoFMvKM/i70SgVmYr
k1r3vUI5zsh3uObUTpYyucWXMFRD127cpoIlCFAML9sdThPFMykLW25QqsXJ4JWg
/MJFyTcRGO1WezB3VRf0/JR/+HADJzQgQoqirnIBUwU3MyWw4M8/hOoA2abfHLIw
e+hVbfWcC0Hm0bUrKRWy1wX5nL0YlBcGE3n9sIRq7ScL4ZpoRZ6/6GtSI/lzf24d
QUJ1fLWamwtyBVBQVKV3vDSoiHXy7KNRKvbbS6fBZq/jvkzmX7fD4v97BAw9TTFf
DaZ/q3xfoY29onJ1ryrIR1Ss2RE0AcAY0czej4pyvdND4PrIi9WHZgdeQOkUQ1FG
dQOoj1Zpg3+QJsmAcXV/7AQUgtUDZzOvyNudPYGNAno67qC96KRycFa5EriABvJq
wKOPTzf2UmgajxkNNxaEMwE2Wo5+rxG2Dep1DGJxAwYh6DkhGO6wq62EJfpqi9Q/
c/ObtoVq4wKSap8eQtTcz/jph3U0lPtXZAonCAYykGsFFfTHLeWgjr5uUVxrTJTQ
EzxL662hUfOUCC8EU7ScBblJZmri2EZJpb9K6cuJcD9KwRhicKNlWXAERYtNeL6m
UbRuejXfSPM9b2YJxDgk2W9xlYcUa22tQ8jvYIWo8Fqeq6NpwNrdrkLnE+xfE82a
shv0jDAkbWnG984UIKB/ZZH6raXVppHSMrUAHG7N24m+vOxYVwYu6wMVOSuY/D0g
j+0uAdqKq79Q2EVp1qgptvFNOv/ko17ISdnrCynvH6Kulqz9gqJs7ToPFPPvSzKv
BjO8fCWRRRGGN/LjjFaiLZFD3eAKZpuvt2flMxDGrkqG3NKYLAhUEVlxkzMHqHzc
+K7CaRil6m9OeM/t5AHuxmmcSO4XcbPY+XugqOg0maWHiV4CfNVTC6YKGdzIe5F6
ysjwLgf3sXcouSrIgOhvXM28lkgl1ZeVnp982Qt/IlVYiuUZ9s9if1zIEXBV1o+a
gAumL+S0mfVOJn2z0yW9ZJ7Ey653b0s12UJZ0c3Z3/Bw3sXyMLTsZNI+xwhLaYmU
ymMu70+h64BHfOTAacmdCYJ1f5/OJc1pCTRmHZqopIpBpwuYHRtB1trJ5cSK6C1D
1yBEHdstCYCrFL8n/YkA7XYtLqzN76Wp918XuLa2vdYk539Jh/jp3ChaYKh5jzuX
XnAuU030qQL4CYEPBiuVxPHtZ8M8acslJAR3P+5EB8i2uArx0WOvQCkyQiHBStej
OZaXhyYeo7ad/ET+EDkOIQNBjQzkggeoJNwAzxz2Wct03xwSKskpt5Ihx2kM2tar
UrHQ7ZpUPbYzgZBfnrxHj1LrKhTfDhy/MAm+8EvAT8tgWSlOo5GReRPZX15UKgND
P9swlHyXuLrJGfHgrteGMRY4csgsUjiItQDwgazdS4hlJ+m7syQjhW7OzYns6LEB
Pi3p2/jEqBd5yAulTrv8Bo1h0KYpTTOXlNHHAm5txUkNWXZuHel8PMDwpcjUmsSB
6OOnqOObCiSC6OlfuBJ5lbkW8ED7XT21jawoRq8gWhce9mq/yeBJfH3yT6BxyMKJ
2wZyfXQ8GFI4k+xQUilVaSFOZ+wPb2ZzW0d2F+mjSxVEVOTCMtI/5dUFNvbTqjJ1
Iu1SkVSP9w6thHdE772v1dInm6gjWY6M+wxSJUb93P5tULLTuf3AWjcAP3piUWY3
9EKJLmDJjlpj/VGh7aZfa0W1wqLoblcEMLWXbN++5UaTsio2WS3FrT/JcsK5uZ0w
jNSlHSb558LEI7gUWDn0+iMpB5hlb393Ka3fTTQHJaCUKCSu9WWESC0fe0jn0lBx
55SbhDjfzM2iAls1lXvKX984ktIiW4YuGEvF6jwYomF3SFzxUSobi6ZQQYNInIQB
Skch96Jtii+6oepreq9g9DnddAxK2e6bnYmvEFC9L7xOkUzm5jKQxajDB8XKtzBf
LZSPKAkuLu4sdwHQQ/G04dxLyU/QrsbWv/vh4HU/UXn8FbWIM6Rqtb4bejsqNDYC
NAMYQJ1eL56+81IQQfHRmsnf1ijV7X2B+LiPXIuxBprGehVpdgH+/duRA2dMLjsG
E+/ZPZmNq9EcAEq5INF3eP41AxrmmvQyKACpiBB5DlRuLarWT5c7K8woDc+ymelp
LhYa94Xgc6z+z6ScdRQlNL/+Uzc3dAlb+4Dm98NjMAnX9xCkjXFdudCIp/w0b3rj
hn7RqB5Hc3jp+Z+Kq/pSMEnqxhgVE6s6/tCd8Ou4ydvKI8TT4RR5UYA90/2drjBo
KuLvHeV14wwcBViLSc25TEOu1IaS4QK5bH5fl2d3R9PATDOdtGNYfWKNlmkEi0Zt
KEyt8k3BzaWwxmBw2O7hZb1puXSqG9xJVL0ohFmoQm23WYhObz4FqniYaqVf1c52
RUU7WQMjpBkIXM0ISg3oj/cTtdQXZN+3+05pEXxR49QAxSFOtN9SJnz9Mc+Mk0MY
UEMr1zBJg+3429ZQWTJ9ah96WMsj1Qy0woAsDwsCadfjwKU1yLIuwd/5bKdynpk4
YV2hQFM/C1ChoAb+1pByFyWVtg2I3aIuUpPsWjJ3Kbd7A5Tyoev9zyRNoppmwD7+
nI8ZUPVt0u9dcH+Phr4pWRWlLvMNmosuw/fTmWdlaP83iKO19XnYDWoMMHXBJdjV
nPqp+nUZnDdHHJvkOngzH6s2I79rrdFDu1ox5q1Z+Iri+HZXPcCCt1rPWXBE1twg
AHMLpNeje1IxEvkJ4dTdGLg/XmS1MTE70dAdISnK2EqzzJa3yrnQr7fWawL/eMlF
B6Xj0c9uc4BubdqtlIMjhpkp/3FxYdrScUpa+HKh+BmtkuAe/auQ03PQZ36mkQmc
jCChN5RgG/U/uTUc7fjbLz+uqcOIKDibzRoTHcd5hXR9pHaQTQICXvpjtsyRU3nX
3m/ShEf+81Bu6q/jkF7PeI103h1jxykvY0nAeUesufHXiXR8QhtFWen15yUyvJnp
LLDYBrnzXGCJ1GPqh9et7D8ZW7Lg9/VmY8eG6QjeFx9nOuy+RjN1cpICSsaUrtCX
Nm2MUXBvbnXQq+ZRXJw2Zq8opMH5K7FYC/Tm0SeRClrJw75KQJQsp/rX4wfqTKy7
RbTgNFZBdnw8vtsGOt5/GjO8gMRZphv5NcRoJCnya+q1fsh40CXZCg1tjTrngeuj
cua4KSdxWszHvE6nZQsFwC4qHcS/PDMeTTiaEDOHI2Mvp73P6Fn7JTLeNJP1llWh
Sgme+cZ8tk+v3Fzwqz8femgNU1IuqtRk1mmuV5uxPbPHH3g1uab1lx58oUaKKb0A
0K7TwsBeU6VMJxxcW0Ymd/Qo2FxwgrjFbcXG5x+DcLW1v/KgLSEQnZar59iPhjEA
B1922cc9HzKTuHpH9FIJSvilOTVckVQH5d3wLYHeGXOyZQgEgSNE4k3S7K5z0871
1zfgXEIR3BmCV/R14JcXRLXrtjDbO9dJNhSp11hOBwkDDtp6e0e/kSKSOvYDksZ3
OoGV/5r6KNDDNxhM5y077DVtS8EyF8mi+fs0vzyKS4DiWXKbPKL7cWqfn7T9MSf1
q5+cShZ7YoGoAoLSKwlt4TBwSQS/HKfLLa3ibCBVI8jUVaZtS7KJ0r1HK4OA2e8R
NZB2BGFceKwDpzQ9NbJuNTBPcPe6aeYSwvsPu8uKKDd3IkFjn5G29nkBuAfTUO7S
qyNAE4jgYCB5+A0SH3vP/1s4ZBDhdeYDlMilnm6F971kLQ4tA7leTFGqD88a02RC
e9nShQ6Z9Nk5XOKM6A2Dt3exDYUBP4HT4YjGSQP0OC8oBf4n0IFLpAH0gD5Q7PT1
KjmocswZ+V9xMXzGIq2Ns88B6gljmDV1127YCClRsWvcphbImvoFKGM2GUOtIsI6
d/qxU30h5Xh9FxouSjCjNWtJFs6xpgP7AfxD9Pd6RCvOCZ9SrBWeYxxeuaPQfdrU
/ksvg4OL4Dlz4sRaPTAMfXEUf0iSwyPHxp6fz66hjytdBVzoFc+h/bnJHdfEUP5J
T2ZmpbC02ZHGXaJDvMtdKV/lCsT8+nrqcQyLIQ6dMkrh8ssWE9HE2hK+RdnwRDin
u+Jx0lTdQsm8korFo7ksZw4wKUlNmRn0o63wvVPCeVshPGNDDD0k/tFqmFX3sYgq
UyLsJ2pEyX7O6mmaeloiHw/VyRKBPFpwA1K467CqLYtrdzjJUlGVY1sQY4ok+Jez
O7VmrRTOHvxBvAMUFOgSxaX3Cv4JvTb0KUL4yKWuy3dqYMMpQ9T/n9GTY8vCJGa1
Ed+nglajGXYD4gK9KlNHZCOpkqV3E+ml72F4GnxoacZjUGSJQvZoX7veorOCpo0R
J2y2M8V4H2V/zrNQUcUcEOThd663Gk+1bN1Br1+dgMWBfOAGjcV/gLfTdvLbcii3
x/hb89p/ybsbdyY4D7Hui1SQchNfNLtUzJ88w9bUCHMJbtwklLTSpNTgIk0uK5MC
LIXS36jY2JxddsuSIWPGRRyFY3Wijrj8NUkD5iUSDLfRRY10J16ShVMUtC3cGewQ
C7fDl4oWMe6+h4eSGnE2DQzcERfJncvaKeK3IUba9dO0T9lxdFWX7YIUrIHxGji3
NVRfCyLXCvWvnx92FQbbN3WoB+qUb7+OVAOJPDEp8gB/S7q/SQT2AB2CCBjz30OW
1xkpK8pR0TePKFdFCDrLQOjZFf7yGCVVledLpAzJes/cz2GdullqatOoy6JITBtK
jhdmmVtW8TjJQGW5YxcrbXOI+BmIARY/EBlFDo1eCShg2PBsuz2D75NLLBQsHgAY
RWw3tjm8Dzs10wn0IljWZwOVyyQb1bQZs4aUWyC2FNNvgnJIRldcpEj73E7JObMz
HbqGzC2FtYLl1WhzBD1GqkCfjIW9na2CbhRRDYIOW5BLcwqpJjYt2/s4ODh+OkJ2
QDt5mkt4xlhak2CLGzC+Qxu7D58S5+TDhNZbbKT0xK3/1osw+MPM0RSFCeUHiGR6
7BEU3C2Se7hNGkel232O4nmJa9UxXfk5XPzf+jd6AS+6wTf04A2tQdyIwkeTaPzt
fuQe3MD70e8Bhy3kUwlbo7D7ha+hJh9LVecK459XcY9A3ALZ3BKTerWGk/Mw5634
280dWlYT1hQKJBekysaPS/BAmBjYhID4GGyqxDdWIrgeeUDSFvIBGuF6C4BKgnE5
4vzMpq27TGcXDEF4Bux8JZAcWNTH3uMNhMX3XEjLeseyHa4XQzi0PYQcT0QFT7pl
ayAJw8Pl9zXoKRwiuoejIN1JOHhTvKr2AZsScE63vq+wzr+Saz3wwknsw7+emIJn
dk2+WoPjPYGHENnErUn7Gc2wcBEDjN7jFxag1wzTBsr0I7/GPWiMJUMZFQsaO8ns
`protect END_PROTECTED
