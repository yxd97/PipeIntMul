`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nf/Aj3rAqzytdYnRl+CCzxCc4BCeHTr+2Z0sAwzyeVdtLicpITuGJ3cWTTkJq5iJ
IxHblnWxXKJK4oIFt9vogFlF9/o6Tp7xbX4EFNt6/fQVtiNgKd7UXmGsN93/qusW
iGE0r/mAmikFBRAJst0nZxxcgsq+nLNIX5eUwV02+4OCr8vcrlA63I9lkRzr/8iG
H+ERocqxijDiB1gAhwfvg3hI/wRq3QxIL6qJBLLlnYMu2e3LmO9gmkpRIgfuLYZe
b3NOXadY6k/NjEuCLOd5gRtMeJglx7TlYzy9dGZ4VDIs4in0TPYTyoZFvHcgTbEe
7Hj1LemgkqjqjSA/ep0z58q9KuShGY5X6nkqrS5AW6QDkouSq8+TsSmjM6fCqkZl
`protect END_PROTECTED
