`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
te6n0RTEFlkCgazePv4buG1awYqi47jFxzbFZmZbTFL1cF1MgDZG365zeO7fcQH5
EcTSVPbtxLUWdf/7KWm75CmJvKlZzk7RG+DPuKQNC0MdXlVOU6Qaxgb/N4kKqNqj
fgE59uK+M2SKWMEQXq80l0a2pVXp/InOb408h5NMbFnTGJNCH21horHol2OulzFL
zacdmI68O07SH96JQUPea2KAh1l1xpcL/M+1TfREgtaBRnVD3tyUwDmVlju7FTMa
yKupr3IFi3YJ47lgl54D9mV8/6QKakJaeIwVU7yEs5SioDqa/xby+v+mLZkj6k13
oco3cmEkwWJ26A4UawBlBw1vXTK7P+Q5gKyXcvbTcll/kZsO0x8m3zaNKIbwHOes
lEnD193auBeCT7pK4UfDK7IKPIQ6c3E2CD5y++usPYplTWYEdWcbpmzEoRMmVHgt
ZzAdBWYFpZ4iJV459LECb7Zoi4zSkk57j7VFe+g/pmzR1cq6oEmuXuC1jY2maxEv
cf+1MtAuaap9NJ/f9UWxLLsxAMyTedD4JqsUAj6foMJCVsILI6qIUtKGto/7foRI
QnPpQhEzEWV4DX/kI9G7f4K4+6SFXdT7ECBA4ar2zgTjfttQuhH7f5Uoytd5cJ3C
+nU4+q6RldCuD8wICTbcWun6GrJ7xUzugezuCk3iicIOgl1J0PhbwVWCi/MV5hLj
TBv0LFBKYxhyzEWH3KdrpA==
`protect END_PROTECTED
