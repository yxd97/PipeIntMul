`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J0HT0ti7+bdLwS9HTSqCWAqdpXTqBBzqfC5hKROMTTf8spZ6j9Mm7DiyG/NMhOZb
t1Fh6N9owR3jZeVhCLllx6+PFdgagkd3X1mGgiSl132JHXkJsHW6tx7EgV/AICD/
RXf/31Q0g8thTREPhaNzVCc2qNNznK6y6cV8lU2pwvaKgmh76f9rw2I1VE2dZ4f+
oKkuf2S7DPerS2TzzkuNgF/51DXVHZRwdsobEPQw48LDMt3pXIQL1w1FKAgP+TUJ
MX//y7xlf2WecjWlOSjkgk6UtDZgulKb4ZfchC9ZAccgpCzCNndNRG4n1vmEjnBT
aZDf5XKVOe4Wt1RtxxUg/5Qn0B/IHyXb589oX6wgH7XsBlA/BvkWAEqMch9ASBTM
XOeX/9FQcvJwyMSObPwNgw3NVoKmgyDizUZB2o7YljdIQNhZwmroLXM+Qrq+1py7
`protect END_PROTECTED
