`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZLYUMiBpVH4PBDM5q4YgfZUZCsz1RW7FLorMcPK3Ff3mcoFwN4GuMfILnjDHS7z
RTrYmjVnjg0rfofrDUPiAFL7dYahnNZLl8cCSxRbSc5+xOMKE35nxtc0AtzAxf/F
whGLyVlhM0Rc3nIbD8AXTGwnQGbQ/1hIa7jWU7SvjoAVnLiEWI6lhym9/dyqehkt
ecN+As0sW8fdUKEMNTZjfj34d05tdmkj0b6Yvkvh94BtBNEUdmLF2Eusnz4mUL3s
7+qYeFCO3hH7SPF4j0ILJghYfXq/NOZKv6WikNIiGqbpOyHCPoW1NVQe5nLV0Vbw
DQnCGbAdCRDgBOhz3JermPd+ZIklyTx30iOY6jJvkMZnQ94qzu1uPgtJ7KcBckgs
gGRozT+YVn4/q013eNKPyJL+uXx8mjh/8ViIwLW1hc8pDem403kuHrmbOnHHchdK
`protect END_PROTECTED
