`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n9twkkd5II9+ErDjDaXaClsOdufq5VodKOnQPkic2J2njpVjEJvMpiCaVpoSX5ze
2/r1VOplHdR6NrCj1r8kz2rrTbN1sKqaerpvT5jHAU0cajXYw2Bp0i5PmZ2kdjY+
Lb5hUw3Ikwf0DmP4/ir765QcyUYY30cqDx8hJZhy8GZiNEzgZKLCwHaUmOrSg/C9
tnyvPZOi3lxv7JWstwu5JddgMRtZFS9GloSwS7LDmxWpC2pr3ZYDoMiQpt1eZvS8
8tX8CUcjKL7hVrG1BT8PZFpT1J+Q9zWNNkpcvaQhFi/+DWTGPxA+1KsHtbc/ok+a
R4ciCULVAeOx9IwHIDNNq2X4STjVni4wldr33Rs3wndAaDi89k/ftypv/dCUXm6k
`protect END_PROTECTED
