`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NeNJZul1pzrxu1u3Ld8U0QI1M13WIoxrJiJSgbPaBytMqk1AuSjIwQ+FRrDezg8R
Ipd7Z9Duuz/34b70n+i8BpHXOOWXlKaU58nJ1cc3mNyXuYhA0FVCZwor16iuaWRW
eZV0dNRKYnwB6vYGqGrVdMS85F+km1Ot1XHyDxVZJqvX38UZRQag+ESWr29JXiUz
ZL1b7hVlAN43vhgBseltwbRwWcrkVWrxeFs9Uz+7bcuZoQFSVZA8az/ipBlK0GsD
IlGOa4YFrFgrsfsWWohwtkXndfvdiI9lfJHoHao8asEz1u3TFjsXsfwnZlY6szsx
oyKtivKd8ABPC16D4xHGiuQo9L9Fb/+1Nssh75GG0NBu9ChpbCGdmazzVoZhOstO
nY5KcV6kYwpObHh+TVrLXA2OzRt/jNWbH8Eg//jqgo7f53YTrmdo7H6mKHjqOIA6
UOCu/L4sb5OA7OW1cWAAkzh/zhTH9qlDB1Zxl7J7e7g=
`protect END_PROTECTED
