`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
otrtIH7cB01RSkXJEbqt25pj2DN/DUrxb96DGzIgXAnZ6Vlv/lrPdBJkfO1HIPB5
OIFIcXeC10cVcKYoX4ikZBePCoDwkqVb0W/6nJC6K2GCVdde1IeYuC57N6HCyu0C
eHfCLxGqTJF1NraGE7+dvpLFErw2iqiQrKXgJ0/H+BUaNOjkKZX7+m0SuogylhmS
rSnumusHWvyEhqgbKnej5IaNxC+NFQuGaLH+0maQ/yBOY0KzzA5kMq+tM1oegjxC
rHF61k3SIiXVFiO+itVX62RkEHEiNxd3cis22/qU8pcCHDzy1E8zu6sk2rqY8sR7
DT0sTo9jTen2BV+W5fwY+fQb+4slCJsRA+VCc4DLRLNOVtNicTJFGdjumZVO/7gn
Dzy0Dg5MhzbLaQFuM/GXpCSrKYDdbCnguE8eO4j0Ctd5Zg39h4MAcDNsxhcqZZKR
WndcIFNHh2PAD0UOJAAEXytVaFDsBHv3A/xB15asKUVN6faWz5kk0StJ5f5Gkp8t
Ef5qXPn3RTD80IB0kQzqdN7H3Gg/ps3PWXOZS3JSf11qmzljaPKUUrrkz3GwYgqX
SRymSkzhrwXYFzb5y+dDIqn5yIRgTfFmnCq/s8fltQnh7tmFhlY7UAV+y5LBWpLi
0YfTgUyaPtR9d4VrB1KJbQVyqqR1lUu9/6xERv+qNg1f54cJDvs/zRz3XJDnfM92
D0ydvPXA1c+BFYMv2DENu/ONqF1a3iEfgWVFDaA8EosJT4ItnnoPRj6IpCNjnkc0
+1ebsTyvh8zq2ej1XddtzjrYg9gs8ZY/c09oVER4CTYb81n7hGop6XsYP/vnG8He
Os9axN3Fk6A13Eq5hYr8HaumfCxIe37+P177wXebAQUgTf3148Q3mSPUI9v8SkKE
XLemSJhYePbA/xePpgy8MscoePa1trM7uR9XqjEiXJXrSJYw6zmIe5Zti0f6GfMb
lSsw8UvIWYvrxfk8WF4uF0qx4dsXjf7n/3WHflx+O2mj1J+fIjnGU8RkQuAmzEQz
liS2PpbKqyZ9eYqNxgq/bXhK2tqJ/AmXRmiXR4zm4NAnLtRYH2+ZdrqYERYQ6Lih
HFQZTl/JXGmV3l/HnieiYSU2rJg2y5Vxk79rVn/B5SoZUzlhRGJuGICUYLhOBM/3
6IIVNJzTUzfBvjLTIMENFu7+fcTyKM+7+fSXBhIySUziRMHPTdTgJJhUyubwVhRH
KfrAy6OV6GVCzJeSETFUpP+dawlERblsWRxYTDPYsqQIRBh0cA9Pyouz49/tkABC
XAW2SDNNVwESY2Yc0+T5Z87cEY91s0/4qgcf6UQ3GMIu0gBMxDtP/20t+DvA2CsT
BNHq+iu12e6NVAjdabxv5QqpIDsS8eVWdfVS02SyDSljKBI/ibOntNATI7NcG7se
FirBrlIdjAf0OaM8O/Ct9jtSTyI2B/XH0qME161aOREJPsOLrcbO5e8d11zoAD3R
7C8RnTZPMg9l5ALKC2d0VeYSXJ+ow0wX/TehgLKehj4jnPgkGtbNNt7pjNzHOzs0
c3CPQ3vLkvo9iWeqrGcNw6FkCIcEP39gTdzPMnk6I1aQuzU6gW9c9h6N9DokVejX
qmPBm2Zkw/2PAAzvB7B2V9tbpPVqsW938gdYkb8Mq5Z6nyGbmx3+glkELnndRrxj
P3Qnn82Y8kso4zl0yjwfIUoJPrHSKBaod3aXtjQXbMPxokAstcglMeuZIciZGI44
1sSygTDzSjbkzBaVaHjetOahbRMWW4hdQajSDiG/rQCH/d5x3OANG7pT+yqyTe5q
ULLVLg2xxv+Yn9VH6dJdOYVtsR8qJQYhmROHUfgcAo9cFETAkIhyFhWUxwm35oKf
5pxiCVi+auLUKrajvd7QgRRQpxan1BFOGFeFTjX1lmbGybyOhntHZk0EcsOiUxRk
H7UZ5w2sDAUuaGBn06HRz1c2fQxjOGtc/kZ+TFYVgaFJ4oE8IymeU8k64RuAp3k1
BTRkmil92o8n8RNvJ09INNQx73naAEsDqH2948+oMjpqijgePmVf9+ad8G+a5SG7
BRA4MD5Jq1/ThNrWUwWdV7YZK7JbEBe6cErbCXTL0Qyo1sW6mt8ctRPnTmrowezX
dldS7oXSsSnDKhZINnlskARyIfucuYv11hrgUIDdtRB0Bp+74ADfsOmalZY5KVxa
92PeFSunPPgHpq5uMSCm8mWHecgJRsI0IlJ3PE8CelbI0wArl+0tdS5ExvUkfD4Z
zIuDlzLW2naUw3PqUt7+yyTBVsRkp8AAGR0OJ65hwBksUI4y2Sdo5sUx0+1oFia4
Lp6xSTURpBrEqPexActo8BskQd6iWki91SzN8nF1LQ6P0EAsC1juvJIWJrGHnUlT
wp0i4z9C6tsnhnAHTnB+YItuPp7Uvk8Hppg4cuf6zflgFj+jeOjp5nBJLOi1B193
YAQyU4hMaSWjZmZx/nSGJmjv8msurX5ocx1Byg6Vn/sSziheSGpa+nIwhchUTUcv
qUFBk6493ntX4dYHiSFIdtw6jZmhGdpFAJr1LA+08G//3AddrpsUuFaXPWBKiqNy
Ihd188SerPwelgB+8Jym4h78ToJzSRMrkzRe+UG7CdfbTzBo6hrUXxHgfemiRlL8
K3uq56SojMfo83MtkxTkZ0zF/j94HcnoS8LYO7Wj/vH0ToaEamhTSXHALWVj9EHi
f8rdM3s+eydC8RcaZKoH2AtAWp0dh1mIqMK1eBiISbs0hPspvuNjfuOvbJCK1Mie
/X54pzICEYUm2bMS/TLSgESdjDRjIAnGoiikatgBMDwzTAwMjlWIPNM0PKRbq2xj
gkRyZCcGxuv6q6pD2VARpnw9In48U5LVIpNiJZWLta6FJinVorU4xsC8pzz3NgqH
XDCR5t9DqFa1+Z7w3MiJoE3dMM/e5fTDEc2YZYuUx0EpTUYz0nMGOR9xD9Z/Sv+0
kijycJFdwYPFWwqRrlAMJdhAGLnOdIVt+ZKos8xVyzq6h348DZ8QfKe1ZQWEKIsQ
np/2OvoGwfbdUQbQAANPvSU8fBM+Ef9aXBxmypENN58rYY95Z8aiyMyE+4L5hIxu
SjMPZSIEBmQiclJZYyJ3IxxvmdfRKI0sSMIKJN77Oi9u7b9PWzEYD50mUngzsCd6
ddlVY7seldyonRvpa50Y3JQ6U2fAtocBT1dfKWsFin87zMyY04Mi9hldWuz8NIrG
Vqc9bwHTWYU9s7WBflUmOCgoJjKA470Dp1MQndsKohdDPOwVkhtQynadSl+xRwj1
M/sKmGhnpfp9b4G6//zS2hfUXvbRrEI/qQ55RUT6xouisv8BmnN2UABh9asTv3gC
LqezqKfjLyxZVG9FdG7EjCKD3qskNl3t6WVUsj68aAYHLww2ADfZ8SkFeYfOMAsN
v/dqCpEXC12F91hKIh9Dj4igpbFM/x+QVz1sxO656IsKUO5QzJKXJV4votFq8vrJ
xyasV/dK9vQm8wb7K/dRfadVes7mJ9d6Loc/li6xJSyEZA0PdI1XU/GsBhShTXLW
OAzC0hKA5pcHvuZYRNBQ93LKHULmatQob/jEzMEEUgydZAyZKBOO8MHdDgu+ig1Y
Um/9Zkge5CySqsLybfiAKMT8ROoFsxOiRIKbtcQiL6z/7w1heQQT+Ouj61ylIIkE
QykKNvBYBb5LA1zhsGEC9n4qg8YRpXpYV11R8fzJ7qjHz7nM0njP6bmnBmVC15fZ
xXAIZK8rZQgDntM7J5Dk/e92wzKBv5U91vpMrcqRaae99V9QM0qn7pC0dFRAgE5o
iE2pZZyWmZZC9W+xCMkbpF8qwa4TbMxDpb3roMPKtPC/O9F4I6fPIldDrGmVphLX
DEoUhZ/qcFyxRn6HEhh3RGlXTCvN8GUomLoknQvgFdDFc0rzPAL2U3DJqHPZ0uVc
7rDV5Ej5fogTtldA4HFcckQn08caFNA9Rsh/hGVnVBL6WN+Kt9TFaqMLy57MR7JT
SVm4WxmOQOyt+XM/WptssZJlV0/8M+j+2c9Kvudjv5mPuf7pNzWknPPeflG0PuJe
qY7DRhmnSkKNDw30KJMSFdLheJGe6EHoXretyU1g8/VMOCVZdZwFzVIps6ft4oCY
51pUFWumaC353XxoyrzeDUn7ReFcwTsDQ+UxauIaGEaJdFa5aD5r/Xe44XQBco87
tV6sFq7BMr4j4EkBw+JvLIhhzFY2+Sbhh5ZB7/8xkelQLJjQ3z3U1U2m/7xtPRlW
MVTHwU+7b+c+SE1iVA9fVhcgrcKfK75W3dli7R409PygHG927OCiLqceapHXXr5O
HwqHeF/S7DwkkbViEPYNQxnp17UsaHHNOg1HraDpJWU=
`protect END_PROTECTED
