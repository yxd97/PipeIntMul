`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LM9BzSPYJDIAr0e9iNMyRWo3YzCPkI3W1Gi138CC2qqld1ei+OBgEiuvdcmcQ2EW
Hy87lek12nTHMDbG1QF/TalgRNt8nTmCVpG40/10k6txIxXcln6bOB6QOKYeg/2i
kpSytezRleZrSarNZuqBhfHHDwCSQ7ILRfF0SqM+aStBRpw6rv8Imv8pFIV61YRb
qcWcU/iunXATNjpwkxia0gDA0A9m589l/VA67Len/A4knJHRu8q5Ib+SiPodqBOZ
ITGYZ9p7+MElSEi+HlydIIvg0wByeueIhNJ6QyyWF6MiNfgWY+Q+tOSy4JxvLVaf
ySxDObOiDLRQlamrcxTlYdAeTFn3R3zPoJqcK7XR1DW+1FCdK+neTYRdldhF1mLE
+A6aWyzWFSMqBj5dN2cTQdI0ho/SN7Ue3COCGSpHtWnSpQdezxgYoSCfS28vHTEU
sR7GkwtUJqewojsULU4VmPVj5rsKEwmqlxjoapmTHnLPklKoR6t5Zm1J2pvk0a+q
ZMiMjWkWMyMYhuZ8mUiPP9ZOkbuUB82dMusTXMVfATEH2pRqrXBkPSwzBKa7N/Cm
+VPEWjP4aOLXJwIM0fLCrCYWU+W+p0H0dnAAhdp2L3iKi/q/EvOcwuMPJ93IzbEN
BpAdZuALe4fvWmspiygyl20vs0GwMd8lrkIMkPxV+hzqdx+AdVSEoeHEqcrioxzJ
bfJLaRvGet6Xi63624rCluQ/wuRXBO9RZjrp79NmycIv47AkvbXn4o9Gac51vr6D
4aiI9pxxTG+V51Wu7hHRmuvvNsppm+j226aZ1npaAza1PXkyb0uvtIMvxeVjmhk9
ZMoLa5xQndzkpFE87j1K6BlQ9zy7/I7lFj8U0YZHL2d0//kX5UEPKdlM+E9LF0CF
nwIKFcaoxDeAxWpTCCaOU9mJCepSgEACvyAy6Ugf3bga5zKv6X/4xOczzyRJL24L
ax6UvrSVooNK1uJ0VupENeZ9R+oiitGLOZuieOMFBrg3E1y0bLQbrGyaR1JtLI41
YHEvTH0O+fTzFovtR0EfwyV29poPh0Z2s7J3rdxVMW59r0JJGKl1pUlcYCkEQDnT
oj5542oGP3siibAEViTcNn3HhdWuRZJinsQePhEz/N6mZI0oDoCvNQ00Brk5cnPL
R6h3C4hKtZVr88+NV3tppXjX3+mhBAwvkn402l/WKPftkVGGyWu2BOIqDhz6FHUj
15P5qE/F1ZFnrnnsA8ymNJj5gyWB8XqsnWQnQrboqUPBMFYZgI5kkp2HbnTbYddh
hSiNMKHQtZrDWG7dI2LMKSl+zVNkl+F5WlWQ7wKgft5aCdX+bp0OswXiKyh+3zFI
8cTbbCikBhWfP3ljX9h7R1UWfG2QgJOcYzKL45zLb9xnnnHaunMCfsYmpzVGgyNU
aFEWZv9sGh0wErrrIKFurzjdTG/vl4Aqe1nZVYuHUym1da0mzNgPue06X1Sdd1Q4
ZWdIKBo/7zfVBZsE4ks8DzFKmtOmuDmBw+pdUvgG8234PpzO6PEqTjelsF99fES1
HAg0V4se9A3cW78nJq9Pz9dwiubORV3XNaBiKTYy7v0P2J9vTAivRKKNQuF8NIHS
6AKJwW6q42cTuLz69lAefn/sthJ1m48DXn3WVxei1FFx2SWIIezBsXRvEt313TYP
EzmTWkqQQDyszlyLpnkMsnec4yV6OqYZL63+GF6Zp0ablOLOBGqcQosrcwZS5/dz
P3dwpIKYi1UOXE+z7nQbhN2J3Hv0oGLD4tiuUdcuCtvHhzMhYkI5xKGxFSiG4u72
OBunkLkJr6WwnuMxzgAvp34CZFWBqXouyIEuW+mfqlyJGs1PnPqb/HbRynql2d09
eSCUBYhxvqaBGdvARcspgAy5nvJ08MeLIItmg9ulMI65as74n1MrIgn1jmSFc7ub
`protect END_PROTECTED
