`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nL6NUPeKQ2SyCdcMns0fx+g4KDcnnWTUeG0B9lp6JhMJF8ipEFVRyxx9A2Epj7jo
7J5rdJOoZ68KjfOKj8fNDf3/W6q5WTlFyxMnncrmKsnwxpnu1LJMPae1mdrgCQKZ
K6CFOMZAJNNrFYT+ssu8PMbCT2RCve1OZLL5rqFjb2cMLaoVcicN65TK2XL2P5tp
Vpa0sITNjdQ2fsYVDMYapN6AFkZVuo7Qbx832tvFx++Fjlk4/HxVEJ6vGOF87HtH
kNtD2VhGtjDp1fxEhdpkOIYRmgwhWbE/N0AU+4Wyw9rz47QXnBcaHdZnenal/3aw
VpSLaZ0a8haicKREcwxjgj0VrHoSJ0YtGjWd6/72d7M/7jJCt3cRQ5UwqzQIENPg
dr/g6WVdu/esnW28X62Bj3JXh9mQHe/Z59oG1VPPLqo8HBNnXSAHrRyQtaiDk6iI
KCd4WAk8A4BNovT0dQByTArEBHmtUOzk0Wxwpz8ZFLjGHOSukahd185ZOi4uHes0
aGPzP/LPc7t9bY5HuNd9+o6y1aKhSfTfvvbRYZ+INbFp5hvbmlkOxwHrARgeaZlq
Vsps7cO4VXDNPdOu+mmP3khHi3SQhi61cexW2KQAr/36h4U6a1x0yKyxSKUhtQDi
gCI2EwzRECixiDTSLHxr4KfqpZj7zNhtGxNsD+cDrks5YgmpMYxE5eC5If77xcHz
S270NqOaRc+aijdOFCAHx5WCmP5nqdlemdC01qTnU/u+1n0OFnfdSCAA5NdFd2Ob
XNRUSJs6gWy7hvptW0xvePLzGg92NK1OxnA6X2aFegsGxEYzKM0ofxygbFZhcU/+
/QJdlZeRJxhwdZhN7gd63S7S6id8LLS+iem4OpLH2Ybls7Z2yJ1YZt/irdsN64x4
IXIz4liGwmYtluIn98iF5eu8qdd5aVg/UOA7+6Xrf0Y4cmzODDN1PE2cgDqBmt3U
knfcpu80VDKX63D0+JaGJKtT+yz3DJHKX4qiUjZx9BTJ35uwblda49Zlyr8ziuSr
RYGnFkYPTLUlAWE3PIFZMLw7/uSmLFfB5Qbv096iFNv2gGB8AZ+ilbpaZk7/SMo9
TXMn0Bphtjc1QPWrobNmPbMExy8HK5H5G77aPqS8N28g4U+YChexylfCoTzEahlc
5/Ehh0xLTD8GayBtEBHMdr66BVtKPZOJe0jIB24qDIJPN8Q6UGgjWr+iyUSM5OXA
e7Gb25YlZI78zhiYOK+D0A==
`protect END_PROTECTED
