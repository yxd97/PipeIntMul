`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5qbNJIZYHAM5oMysbNRSoZSl+UMAFVxjPhfY0ogxT+XvM/JnREXzOYJpIwaj8og
YtICIKtFI02k13upqV/EP8W6c6rf60bkRuSAIKpP5FZVCBK5DWqqMsNQ5RG1CUDb
kYsyV98Hw3wXQ5vkmylX6ovrU+87P3XP7NrezDFiaqbYdFoIW/iLUto7GZBEfkhk
9U/a8O7Irn4vXE94xN0dRObd6dt+HRTnrYKi4x1poAzS+SA+NrV7oiAClTN2lypf
usJOe4rSYwn3vszGxCo17Uor5mqXfG3nsvfozNlf/x6v9nP1d4Ngs9SuUCX/S7xi
z8fMtMP/mmSjpi6mHoOj3bBmec0yaFPzT4XU5gd50nsMINwhfh4sV+yNMraXc7w5
gZTTDB8/0nBKQhUzQJ+lejt6b8nJvEYdgBjbtNJJjvWPt5zwKKuxnCMM+2kambg6
2UzXqk/buEq1Yo3gS9KMTDb2pGZtVl9L02mDZlmbkWezhVcB7RAbTnbzS5CU5oK/
qv9mJ1rWAbL7AUfc5kH3OxeNztfy9f3NhTFqHo17ejjgkmfar9cq2SI7ZlKMe4XI
kX5NSX+ucZIzRMU2fdXdvKzgDV52BuWMC4zODzPKaofo/+PdIstC5Nh05VZfUuy1
FrKKNPiavY4aQDQ4Moyc3gNUduB0PzQFxQ34jIxfO4ViGHb9jE+sdlYORmpuQysx
uSBCoF3ZU4szXGX7y89IcPRH2H6krVM5ffpmIWKFpOD34ikLMDdTrzT/bGiM0sZ0
GVLzfW7xSboGBOwcZ7V+/2mHLbKd3VUrI9i/cNaXD95xD7hAMlgM9CZkwiRC/XMK
sOfv2KTXMAcf7aEiv1KXSPD9V11fv90oQRxH0stc4H5//6GC5/WQ38I2uEhipW6G
N//6BO1m9ZWzUREUEd3l/orOYeDNFPAzguAT70kwngr0JcwY5xowXr/spL9OJzZp
9Zy9w+ETfNziDAhW0nsvale0dTbT2bTQ5aJiPLm87ZCmYvUjQFrq9+e3hwZxpfkB
e2DewD8+Ix0dyTb7cNrX4IOlzNJOsaRgDp2VUpEfs/fMInCtCmSFLZaWNn4peHoW
skOQSDoazOGIsY20zNs5xh0ZsTgUkvehikTk5lEAt2Cz9DV9ea4t+I9Ab80hTaV3
ZqrAuguAh64aGNUzUl/ZzevAj034jyyMv+//H5/2keiOjCX8SyQhq3wyAxrtvDsq
/LDj9AFkyCqoDLdGJrSpHwHE7G1/lQ2YI9JOkpDRKc/EjKA4fwDQjoJvzFd/QUY6
QGfEM/lz/Jl5U4DEXgqimzTUPQ9zU0ziyzIJztAtmreiSocg96r8ZooW/8dXlrxY
pRaUhMHn5+6MfrfbVouwHC9Mrt2dMx6l/KD3mbvTCLfu/ixuldUxT1LUvAPu4QR0
u3Ap9XIXyAkbyo2Ly/ykjBHyTgWNBWM3OQN+SwZxiG8yRjocyfl9lJyGuJc9dyPb
uHAlaqr8f81iLgkv0MrMwg3TUsdKmfTJ4pIgzQBdlRnQBoZSNEXRZsWQ2oVydLbq
cA/5HeOBtFcRag4VyiOaOY4dvNnIw7pom3U6jbvTr5FzoHBXZls1EkHufVbX9A45
+02oc5oz7IBAvoKcN1o7SXDL5zVtK9WRMKjamLk17NR+JfEGtVRgnuWwHqsY7OSD
XLLgKSGdf9wgj6vvz/oVqkOSpiWB10r9V0IxydMMEnp4AdgBXq57u0S5p02e3l0h
T9KkSRAg5z1PKCZxacwUxMId4RdXpQQGoovNf5Ry5oRCa5IXSY8TNS8u3dAWwehU
B5q+T2PAhnMk5J3QRXuLWO9+f3xAGrCazOd9UldT07iQT66RLxXKj50tC4dFrZQ8
Qx1m2ylfpGAW5z2SMGh299gcB9dyKt06nyMvkKpvXX8XaFrmRYdAzGJAFzW8vxLi
dWia2avvwo5ixmFQbQeuwjOMfxbKQlMHDwNnNs3Nohg9rvbJaPwD+KHgI9gPU9wu
UsX7s7yWHFDY1DvqnINBeyGZVGg7uOC0J7NX/qaNCog+wi209Idb1OSV1ekeJYZI
Br3X72lz5a57SOL3HyT/qKwPhYleu7kz8HXD23esxb9c8S5VGr926doGVltpXJCL
qcYRY1tvr043BDhT2ZkNnc1ZMBnlGOvdz9gy0DdK5hv/gZLdCkxjjK6Otega7e/u
zxvjY/t8gfhALOIdk+mx61doxIdOaJxIAtgOen3VqvNiqDOVdjNBMXgF2dJqvpKU
w0V23+ZUMsK488CwtJp0z4J6CV97EfiduXk+PPSUUcEjWV6Zn2J303FAQRpSzHnr
8l9xKqjo3WzqMJUChEMjjAtX8GokozbpZNb1ByZOsqkpGhzmkDS2OoFHgCHkxMx3
qKBFpnYlIABfD5YUwg7un2U7m6td/Lg6MeASRxyOaTr15Le+x47/RzMYgJi5u3ep
0XUh+nblPin4wBDCHpjlzaPZpGa+v2b0Emvgsc7c7YrAsGXTniSajYXWXJ+VhZdS
MqWckGfvjbKw0I72uiXZ82Z4kSszp+2Skq75M7W8YCNGzHT/36HOzQtOxm9mrAMx
u5v31T3xWFnLkwEdXfGLdf5OfLrEwh6aJBXruO9WYKrOUlpxIezzr/OhOo5IqJIo
H4fN+6BS3aojkKjs0/OVspsuF/DG4znZLUo09Gp6iCevYEOaez/RGKRnxyNf7ndP
nm27p+r5i+6f7c+JziOOmiSgUC6OMZcpJpWgj6lSREqxApEdTaWjXtCZlCL5sved
RhAjxNvJBg5/1tx2uqxPQHj73X8npIhHCYPIgZNml4EgQYu6aT10WAq9EhY1biqH
oubLPZPdXPdNg7NQWflREYkYwfOOi4bMYgjbprcV6CyeTuA9FhpP26g+sYq2UGDs
lEfGh296kFMnPl6Ai39Avv2nZVVSYexi0i1gVz6UU5DCSSldKU32bdPCYlxPkAGu
ZqNqbZ32slVf4bR0PfqOkvR965Sono10pH0g4bRJELUu6kv4YZ3gVSqC043cu8bU
0hCK9XfdNQROlrtwaoZzA+BpUwz/xgzd2zPAaBvRxf4vBfyArclVJh1ByXYlhsg6
WnLc1gbGr+gyARxXjS2a19QCYsmDLni10ZONglvtivE06X6hEwwm9kvczYlHF2BH
a4Ke9ncCmCiHSJZ54YS9GGd/VV7kOBNA9PnN/bB1YGJyvTIcl6ABqq0ny3HSGLY6
/EzXtDbckbX1qa0hr2zKk9ZImnJnqQ4VnYzkashSE1CfFI68y7YrG1zwODkRde0V
mijhBsSD29RVSCe4vWzBQ98TI9C4XODZkBMzvute5p+WEY6E+efzcdFVUPmLuaTW
p3PGkipLMwL70MRV4olJ0lm1s5NEiGGuUy3FNeL75rlZoxRYwW1lt1FVqQLYwXUY
96fzUr26dpLm1UHm+RHPbpb9rvuosX+ThvAW4Mqv+YsmfVERb/q3AkqL2q/kODy9
H3FtKPZLdCmNCrkCFHs10brSCEmNt+aOUakgs25teryTyQocv1z9JNmFHUJyHRfL
qBi0ypy6K9IPA/HoC6l7JgVT2VrqmhIMCBqcRaNccTS2tVuzmW3ghHLC63WX7imS
DahIaslGDtZDfue1PXKvGuyOpu0K9fionjjCnwL6GQ12dsNbyKtfszjZwAyQYFpC
VrVlwNGguZb9CXgB+l5f8ci4wBo8lcRZQkOPx6hBsPXOUonGVqOChiTVu6rKHZuX
zGwMf/2a6vPrflbEz3d5YU30Wkdb87sYySMevOcpQJ55whx1ghxEXxVjLwSMl77U
VtUS056Gr9LPZtuJdJEedzamUfVYQ9HBt2xmzfgzzf4omAWnP96qiPtyuPZ0L7PN
tiZ6r3h2zaO75XaD1ER2skdtyNK529Q03e8AxoCJcDlZNZbShNx7RbwOZPzgTzUS
5wmoC33tWo9HOrPz4W7HFlfzfV2oPx31HMSywGb1uuoMCFMSFqYPGVEn/i2Q4Tfr
bl/xnjSA1WBbXNtGWbyJ/TyA/5fF/Uv4W+oWEnt3hdm7Lt38SDcxWrY9O54OeXoP
iBSJtuRtBrdtziivJBoyxTjbRlHDilJGK5duIa1xWR3uJ5FS22D4XPgioQqNc78c
Dm0x6cLUKw0KuAmDVVHzJ06MisWfDgPDGEo1JiEndr/L6FJ4OP9jeLFM1NRVAN59
atROFD7Q8RQE8ESc4wKx3nqWkx97opO6rVWPuHS/A2vltHIN8/Hesz0mykvxakhU
ZcsoGiDdygdQW4swNhqzcyAqFu389OEcu7OPeC3/6MUDElN73MBEwErQe7LtL0tJ
H0j3dFajZqaqcZvE2q7AhSAEjPTU+IKLwo8F/IOcB9lbxsQPQ0dVbU+TOW/fw8Ie
gZwAVUDpkDEV4yEWDdKX/856qCiiY32tkGCODiu/V0hbtFxrbxvxJHD1Jon+3RJM
uwi+zcOlPhKENnGLyNPLoYY3eOwAwfLDRjhz7cR3C4z/87OKdwae8nAUc+OeK96u
nh9Ey4NnQ3P5Q16gW+qGHNxsBpY08ckkPUT9W6K+qK/NWKOkP52Gdgth9KyI2PBD
eZenSeb0gsf0KzmzvFXZm+lrzUiZuE6uvBBIMNjvd7WSXKZDzJrRMmtDIebZk08c
WgZYhj/JaUR4maCesJwhjeOXatf+Ci9afv3AiOBMppxgd00PS3smr5Xg90T3PN0b
SbcE36xKG4g1SGnA46wfvlQk4zQAZ0OSm3Wd0opRKqXyYM3VRHamzySWLvMyPV95
c+JHCdrD0/VBY43BFn+mDt8qwJu9YHS9yUanKByE8uGGn33BWjnXtdJTYu7r5hAo
bFw1oIiOSeEWBVVlKyO5E5eiIbIIq4BY2mu0hZLwC8fg/fNDNCpbRma2zRAgTb2h
E4y6zvnNugsYrMnCP4CtlPzPtUcPxja9+Zkme2lWCaIc8J1md++2Cfa0REq+TjhY
Leli2ZVgvrD8k2fMEV/uHNGNiGsQupj7OUZZuy8jJXer8ym0oVdZ7intNr9tHSZc
vxL+Bi0+pPOn18HuPIRyijrzTFZuTRZckZFSUQCNXZsDEmFhEGr7NRQicc1woMBP
vJREKOAjeoLzSWMgnbM/i7fK5rtpZIfyblYhZcuuf366I/eNvQIsxxG3JcFjnYHI
u/DxDubheLS6x46j1J0Nkz+T2pvKLDXlBWrYZKGXDxXJGHGaW6+z4+/P5ukig9tH
kUdmJH5ujGim91gGTk7erL6YWcIk74h8hUGk+rIAh2JW+i7VAZt32AvOi+w0GelH
AA8oeRwdHZoaWgobU/F59Vwe8g+dKP/QvZKZpP+PL81M6MjvfQEZOe57yxaZ2gYM
jtX/H71pGQXr5iQ9YpK4YxNwAiReZSXIATP0r6S2ZpozOTpcg/n7kJCJkYHUKasR
xwvV3vNJeD9EcgW9NohqFQq3mi/jvFxOfB/Vswz76YIMNVImjBu5yzOw8jmVG14D
EMyY50VD18ILPOoTr3X4BgCHb/iv/v9pjmmX+wM2MshRFhJilQy18rUV8k7o0N5P
JMlv82OE8eBYdkZ2KqMSyw==
`protect END_PROTECTED
