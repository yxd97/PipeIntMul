`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1VwKdxnp4ULhyrp24HSH3BSXCsMgH8UtTaKjPUxr8o6J97GZYi/Iz7fQEDo/VRPf
bLbWGWdkp6fCB3yabQTb+aOlByYq/6hryZfbKYmdecOGPybHvdy2pW7SdeZ/ssgk
RYZTi9DSYVXhxtjXAZxjCI6ElR89MTru/KFGSwqaKp9s6kcq4yUBO6alTY5CTCqp
1Gq0x6BaaSVeMynywRxyR48F+sQjgzjnHZMOWtGmlZbPHoXe6R+uIVhntHPHWpxp
gIrUBLUSiHpO1wUeO2nqzA==
`protect END_PROTECTED
