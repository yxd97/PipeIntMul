`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DxuY3zF5kvZj58PLH+l5G7qI6zQgaUYktU1SWSldTaUhzn8UsxUpSU/sgTeW7nTr
8J9EJmotqCuUn7Dyrqwh/xngwOm0cBlQuJSI36X9WpouMLKp0FHjj/kt7ZT4zmGq
+zYgvTkzqtMdpYZ2muqV3upXCKo6Xw08rdpspVstyzyF82Zr2sCeb4Rs6x6p/LAk
kFnGtF1LDujTuDeFUSAf4mre1ot8/gEM7GROTgiZv4Cb2GJH7lWGBgXW+8rCaOp1
D/jkUUWJFhi11s/lqV2qxg==
`protect END_PROTECTED
