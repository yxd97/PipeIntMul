`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oYqjoTTZjFzgraoCEw4jkcPaQ8O+EQYjFW7Krq1kXt34KszjUagl/8foWCD+PQOA
InxRucIXUAVKap0YgPWoUmpOtLkIezLZfFK++7G+wwlHJGAk/8w26LiVfqVgnLHU
HwKYlor49h3XHouVXguHI1OslqE+uhiEZ+rHUaThAFToFYFbRZspEv1z2aYLKcZE
wZ8Vf9G1c8+wIvgUBLPMRxHhVbRUpx17g0SAVNgcllyP92M4iZwRF+C37jWJ9Eou
vh97M2xnfsYce+XRCI5h1zyyiV15NH3NgYUUDjZULhg=
`protect END_PROTECTED
