`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qt8kMbQxQtvTonQFNsTUwbM+RXAI7U18HzidWMjCJIskf6lMPdg/YA7hrwrLmZ2F
JILQ3B4bnHlvSOunYreVaF6q4gj8saOEQh9QJTKp4+85wrC6dh2S1l1lMc6JtxSG
gzpdRdC0S2pNBO/7UVCvzA3BpvhJ32Sq1PLISIphbzn4dilDwm+5XKlxgEoaYaYQ
t+wcLeBix3o/WjJ8sX/3MWitvoCGYOE5Zb3r8eLF8R7qBsHOKSCDgFuOTt3Dx4xa
QpfOVElJZKmKDRi2Ue6da0zu7W+EnnmYzHZz4Rrhs+USTGVOBzj3p7MoB74p5Mzq
MuTmulcO7Xoiek/U0dQL/EeIEHgExipFviC8lT+x+uo6I9bwWnPdxAUM2irGiSwj
lu7T1l3rItvlQEw+Dz5KXku3hk8Bm8CMlpQWLAdnaexXecci0OUXPmst7fxOuRwO
fCGjj1uhZp2TN00EJuauRu0drVpzi8yMhZv8yoS6GoqC9oBgQee1Xgq9852TwAXd
x+Z6LLOQ/Po3h+OjzMVewTYOVbpGfDgxL/ogDz/PwQUC3s1u6CZfmP+kSC/379l0
J5CWwfWzc/4DGE9u5e98dPiT+i2KescctPE7gqRdL87ebfHSg3+e2L9A1II6e+OS
`protect END_PROTECTED
