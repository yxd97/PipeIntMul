`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yDlybecAstg/xXpHufaBcVq1R1xC3ufU9YU0fq+WSVQJVa/jSWEsJtF0hcJC99+M
wY2g9kjy/LaDh4GhGAD4I3+IdRjopd6c1dAgy1Cb8Sx4WI7z8MIdiGvW3P/sKxWl
+cMTcQUUBI6KxcppCuGy1ftLeSyz77+RnFMskHR0Y2HgzNa7UKB3QNVRcCteG/eV
99GOp78TB5Zs32jB03M80J00hGOaulWBGovO9h1ywjfG2T9uNIpGvmE3NRq33WUb
eR3i8HZ0IrLtdw2ChAD2bbbzu08lwa5SCJJzq3zHkHI1gCIntJx95oDV519c93Qf
ZbIKKflUC/43hbuVWxP/7wA1YS1MY70rmYXZDqIW2/loVHMJVasb5QPHzRrg6a7V
toRWsDoBh+n3XpoKxGMa7L3NubbBxGm1RFyzNC3CEj8TAXRbsSo+FJ8ZbuDNzN9C
eNCu+4xR72O5oTC2YocABPQq/O4j/7UfRp4Pcb75Ax6rL9LBlxi9UsnTXrlByXNA
FCGiVAXAUAZH9WeivMzU/Eh/Hzdk892XwBurI5yaZDIuEmEzHxI5tkdLrXNWLOlx
`protect END_PROTECTED
