`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zbv4yT7g2pLnimcKKddf4toMlDt38KvQxYqVjfiskHB+x6DMKgEDGkztUbUYHYah
M896el/MB98as6EXFyyybDZn7LTXLhYpj9SzxzWH+6y81597D3me7VBIXyviOr3h
om7juYEbB4bUOKw9wQ+qsaGEMRLzmffQdOCRGP2Px/83cZrPaYtAIznyW2zxHMqJ
4sF8YniiSRjsIfHtRuQqBfhecU2OXD64ECc8u/YXg1J+gumN1IzvMyDrtu3cavZ+
6/GJIdkG/QHlAl3GAun7KJkOIbW/vAn34odeTB5eXpGhfcSD8dt1NK+NiSY/uqQE
ICxWsNfwPeyfqlqrOJd2/vuwVn7INGsRxt9QxB7uS7b1384kn0K8fFAM61Ieq0fe
MY0fbzIvGR0USXBYTFdNLtoK5H7HQR0Sx4p1kXVVpAcdBUEk1gflA3QuUwoZCkLr
q46JzLgDBklYGJoithQoecNwTTUSD776Fjw7yY1WS6k7HBNjO/lQCGd6JuWJwgCU
7zhESIEXrnMuupezZKOooaCbnmaPzN0khJrLM4oByk4IRISAfjxTTDVTRKQlXtwt
siwnw7ZCknC1SRHzBR91TQ==
`protect END_PROTECTED
