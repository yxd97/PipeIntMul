`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hkGqHOGEXNGRA1t1P3oc9dhMNJMbg2iEu1vLlsGSttSeWS0hT3x+K0j/boTKLFac
N+oVQd24z2kUSKFwBohMt7bDCyj6P2bIA6WdRxKbI+2ZxvK+NBXd3jMq+dSbv11c
wEFtpcpZki9WJ2+8rt707nqfXvw771IuqvPGUjHm2a5stvFHzYg+xE0wnlguC1HJ
uP1+456+wqa3Iq1PagSPMVAg83TqwHa34DzWMynvgXF9E5gvHRLqOiYX1cByim9h
M450U34/v/D5IVizhah7pspq8dBuf1slCkRD8RAoZ7J3CmfA2jOv2MdQRNWYExq9
GDC1hfys4V9UxBZs4Mh8Ko9ujgwuYj0msXFu2ifhdQNKrqc+LAYeitLAU2k3jHa8
+PJOBZg1j//1TOap1l2OwK0t0SfMK2B3LCV58u95IDP6B76qYBMOfOIAyhZfqr9B
qTemNMp47ZFsY1Du4Pp/yK2+8sqXkPwI4q9OjiUMhS7O6HQm3UV0TSNZmBl0vXXh
aFjiT4cflpeX+gXaPgRl25hKo5j63iwfLlf++wgeFwHhTzbZTRqi4tfV9r2g4Z2z
JKgfeW+Orl+AoRqds4CWG24loprcwbgjRrmDZ6/ltzaeK6y/jv+vuldsSXRfJ1t7
Cge5+GTKtvEzx/jU27FD7DXDy8emUpxrWkCK4zRu5svLsOM+oydV/NZrNmbAXgXp
PXK266KSWSJeoVouptZlblLa3wPMOjaxHD+cCAe0+1yHTW/AZxNz0Xrz8OWdMrIC
Imx/yZ/05kXhbMvZPQOnPRaUKtKasdEwNv9i/W0bTJDp/nC2Fj6RAaPwnZDh4NgQ
j1CBwiw91KE6sco3HZG12IXT3Q8KcVUgmp7si0nzN2myK0WEPFogGL6hwJrCvS1K
/HqTjy59WfeegEiVJ27uEfLLywrju5xN2XqKyP+NnmcjrASJd4e6LHb5sBGPwwba
ARRHBGv8Ou+J9nUc02ZYuw9bkuwtatrmzdx9n5R0mVj1ZrbpBkV236xH21Y8KsBc
9DsMhbLK66p9hcQmIwKvnoqUaIcmrRH9BEpdM8j1+sRkrrZaWPnK/wmUIBwqdaa5
HldVql+fCZ+nDOlCVy1vXIUvRtCucpLsi/ftEratGH+XMhdwMdaefBvPRUqjeDqG
QJumuBbh/fTcnYve4r90FlsDgezWswWBVVYISBO0KetY8Jur57JcSzr8E//rxQwO
CnBBkfVEDfP4WYhc+Qu0zj1c7FseL55e7QRjOYqhUayFGedFNBGg8WeYYZ1kSV4f
3n9R46WuJuV+CVyhhzCuLDb/S80YvVTYrypCMADH0nS3EjUmcwSDed0flu1HKY/1
E7crGVDoKBzi6aRStvUh1flKzzV+xaSYb6/R5J0rbv2SpQmCWizxt1doRVeaG5+x
09xGJsxcGorKu4m7ThixUHfrDnF9w+wQ3fVAprLnlhgfWMYElTqdSHRq3Z8xmBSd
vSUIg6/7Alv87v9Ldhozc99rEvyMvZ3kU75qTIbQ8s+15HaExJPr+AJnW2v7WXjN
9kp4qAhUrlRgwHS9R/ivCm8LqOkIic74gOmSo8BvCwZySDqrNeTdoXUjKec+/F1W
gbvR7EhFi4mK9jDTm3NOi4qyTaf8I5X6AnC26U+ld75ccwp7JzQoB5JkxhbLiSi5
z+lE01OOeQqjKkb6TWFwHoCwO+o/pKlJfBV+jqtJ3hw7HX+4xNAzSnHhu+NpUDLn
2Tsl97qg/FSMOjcaKVVvLm/VBfsH80kknLGg+W5X+GmHUYrm6ouctp/S/yvzDL4g
lQ91Fr6r2824ExaWELIc8c66ua5eq/RBRE+Y/ZkWVtLmVpQfIkGlF+i40wTJA8ru
CbF3sDoWIA5g7rTKVExVoP+sEwxYbry6PSlRV4oRaB4mRI0dQkXMtKO7bQmpexyB
xPoaqgHFCCtY9OCeDwzNkDrzHiDlKZIyQ0mm5Vx+KWAgnEOgY/EQsfjwWX5oafgy
HcUC3KUJAETezA8iGEdknMIXnIrlIOUTDRolsKR6hxoQsnnh4ee5RkbFFxPQ0fN6
/k3H/mpIaM8RtOVwrkEWrSVM5XJRIJIlYMtwhYeV+ezb89fN7qLBFrB6QuJLrSmD
e1j9aIZrO80ogfWKn/TR8eqsbt1n4LoAM7im1KtY8Rf4CHnlPhNmTV4b15QjUUWK
X/zq1a3pAz2hZa6MbknmxOcO1imjSofwmYGGkGFHKOTLugQxDnw71Iy2Wv0KsEGf
C9flNgOGca3SP60wNvp9r9af6lyicnRuE+muNaOadZJXxivB98VM59Wn0Pf6MTph
yB9PniGydY08nofejvTlX9p43jeURgJRhKGl2mVkflmHb5ksFpuKHC/fp2ccGtZh
sH2LrdzW/l30/x6EriEKVzZGR9g40YjfQzCPXCmP7Lqe/RRewKNNh6B9eiE9A4qN
tNG4dAdiqOASnEfSaGCNtrxMuQSDOqhNRMjKafH99c5ttNSEToXDR8zuJF9qKK+f
/o7/RJbU+GiWe4bNc+iXcqRwCsX5IWZxg8aI6Xh+z1/cYqB+e6Uj7uMS98pjOVfD
dGrC8vTudYCethGh6TU3qMqFpD0LX/8LmwapJbvJqMqDiMGcmBVzMqULWC80/jaT
jruKDQRgk7SKmr8BpnBI9twCURcmp40mWBqmo1BK3UhncyVBmnJb/zMY4BYJ3Mip
L4nz2m3VwGPlmCZor6sp9LzsTplRgASw61dA/1vbt7vIbniUGKqgFkmqSs1twtNu
+QLX6TPEF3itn5u3ApTTEajPL3yXk1MVLdIGdvZot+vZaMw+rK4maS1jf3Q9xOCM
7GZWUtICvuEjOqwXfTjxpCOtos2I1vKr3as3L3k5i35VgL2tWGtiI9Up3doQRPEZ
Mrfsx0ebQla6oMlUlV255E+JXsFUUjWTLGNjaqbNrDj7pPZyTZ0LUTkOOlA8/3bL
GL0w5NvtJFc1XJSBqvINcM/wkoFu/qI3csg51qe/wisoN61qlfipmI0reBJsW/eW
/tqGJM7qvnuVhdn8mLrX31eKY8KAjSo18/KmRjXgR2KLhm9fpG+eLmdChTYbCRBu
Ng67rN/hIPE0ok8dAtwnlKjI0QpHSbAYEVSjmaLbUt5KeDATxggrz64imEMSkALF
WalVWeke3L3rhDqEnyc+p4ODtwhN3BzhpEfy0YAZ9oocdrq1v9IKfKoS8vLWFdRH
pD96ss5dhn0l15XVMKhHTjrxIGHKHOk91Lhzq4097SVu5k2CzOhunG5AAb8k/AF1
XHPsxPABlyjpOFK5P/cdOP1JCtKBOAOiSQ3MkliQt/hnRihk0lRZNxdeQNglCJj7
EEuxqA3wWTcX6prEoqQRMr5jXlmaoDVoDTiKjlq5H24tTph5J5QBJP0ekgSU0bxl
+9eCXa9iezusaXyLIndOEq9kb+OUMGs1TpkzWdY+MJrGEi5ViHRuGyJKUiBvHLKX
Ekb2O7r4QQsp9NG+vpBtYo2FA3bthzGf28qZLz4p0QJWkovJGC3DlxN/0bnWshH3
IkkVaxLYOfoImU6vqpY22Vr7UOqigqVS6dXkZfpYdRYZQoLznXnWPmj7E9i60z/1
jHbqHHfw0mKH5FfgOo1ZpJI3DfPIubiNzuUm6V1I406dKsk9xw82j9mRuTINHWU5
scXghoXECGQ+3t8JSnWuAmM7WKxTWzKDQM5ARNnnQ4zWLGK+JCQIGV4OEJVtxoBg
WcMhIdD/YWUA1Gq/Bc9L1TAjySMo2d2oSuzjlKYHJRvH+D/Bx5r+Hw4Aopt9WHnG
zDRKqPlJdek45tcYCrwDOt3et5Ww1qiB7OGTjluRUilLPw51j9UP4+dFEBfIOFa/
TR70GBMQwtFF3+QylL5NROSABhcyg6VEVr67kOA4wQwvxPPq6BveReBjp7kJH3N5
J3/sCQXE7fDOxLPTkWS6Vu/3NyKseScB+mX8WsvhxtpsjKcRMSdwxTL7TODfUvoj
`protect END_PROTECTED
