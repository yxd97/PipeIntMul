`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5aMXOiIrBm/ptHxPZNj8hOeXMrNI/AEvIAYu2FHsH4E3cYQ5j5MZpvnJdTStMGyP
POntYK3RhxSYV0vfqTvgPcy1z4qms5VK9+8i8xu1RsRR882IbbQWsNJk5i1jr2+V
fDHQ+1OaFKIk/LgeAIoBO7RDDtn8CKFlc37Lwutl+MJeyvtN6tUHLxu7KIAtkL9J
bgzQAIFIdOzMbSYOexqE2/LzIEeysBHIBzSOD8PJ+AifyABq/rTqWcSS1LiBSo1P
SjH8thqeENC1voM+fqAuGq0kg1YHCapdIy1ZVdIDAfWx0ambndgmsgpjgdpfJFR3
LXn7u69+eSzaFGCBIHlrxI6I6lu+XM/jtzAX+jFpCDXPFgiCZKJPtfM5CNtqgUzo
IZyprcdaBriQdh4XYNWEgQ+7eUgxj4t/YtNR+nZMEOg845q5tYbT4aWuo+II4NsE
Nb2ErqHous5j/ZhRCUd8cb2sFFvozWAvNJwQ/S9Y4YE+f0JaYESG1ri3l9aRusvj
PLzdbw7yQ2bBU0+VRfi8ImQI5ICSst1beSodLHqD2EZnUKMmEKaahlGpyhoiky2r
`protect END_PROTECTED
