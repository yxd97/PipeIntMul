`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d03iQX9eayIt5aYszLke/yk308TKBssahTiuZ6pP/QTc3qwKbsPSABp8gh0GN7Fu
sTGvS0gQMT8fLjIcFWcwHc9+/HWsEpHu/98uhC6ovS1zToclsl9AnxlHMa5obhTM
K5ZEH/a12f8LOWHbO8l9ReahmPR39sE/rcVmQ9m+l0xFKv0a0boJr9a/9X7FU5Nh
5Y0nZcRjdM12DKY6AzKj6W9thdURqNwJg9OYRozjrVTnPn7Aalx5aALY/T90iiJV
4KxFlA7mhwpT+AO4OrIOApbLZCfRAScH6oJztsuyt1jDi/6kLuVNbyzbSSosZ96z
SZGwSbJWz/44ZEeCxUHgDr6dWOGfpmvjathBaG2iAL9uarKosaiazLVqQBSabCw6
BzUySwMKug0g3CyCqEDfReAH/pRd61X8VgSaQQgO7yF1vyl/itSN7uMAOyH1My3y
s6mV0ZYzNhPFIVmSAjBVv0yFUu64G7LdmKk1ZlBbB/JaWpq8EfiQ7YzqerfLzo5d
JiY/BqEwTpHixekLLI9OfeQFricyXa/N7bqjTz2YeF/Xugy3HSqnlSNBtxoU5bmp
c3aebAgEXlr34uELnLoHYeoS/+uaNXyKzenYlb1u+4hoNx8TQfbbp1vUkmgPH9ZM
mUUEsRPPuoodfOOpHnF0wnHehABQoCKzgjYcUagHf8cCgnbhyq7+3QRkCU6xo1It
7CKrXYq5d8u7Anw7Ef1SL/904KmDJvhS5jR0ZydHZpbsTiFjJEPclMlmf6fZyw1k
GKk47xkueX0XLQ4ScNrx/qDEoDhnk2I0M5mL5rDODYOvD+qYsr1n5FSzvrqIBknb
r6OjCVluDLHeHkA7OrXkcBZTJmYMiy7CUy6tqZ2p8hIzH130rzspySNge1xOR+Eb
9EUylcHGOA+oMyCkmjElhqVVEc2aUWgjymc5iK/0UwTsqn6yhqlMBZjxg/ie6Hm2
PXuWYyafghAoJ79oA4ii6XegdsXVKvhBeJHqAzpD924nHxaqOxqanObOGUA7xx/r
HYGxQ6Is26f0+Ruu3xyiPU8JCQjgcnYhC86GJ9i3OQpx5B6+exHMrs2+PLMGzuut
TQdQY/kuZuUyQcz44u5TyYJaGCsmLhs/U6hagzOEqvZugQtmEn1DM78jafTPab7f
YGqBlf8PI+3zbnfEpUoPl2WWW1njoQt67zdLOZxJn1ORHac7LPfm4LRLikVkUEHW
PNZdE50p/vBuXytWtoVHdWzybPdREyQTN4Vfn2WSCIwtaOAYwSr2c627cTNMT8xw
oNd1E1xnBLVOKqFVrctQf2674ilLo+BqWwd9CzUIX78SDlJyPlc+taEulycanRs8
494onsuBg/q4bRgP7Kq2/IMZWe3PM2Mq6QsoNV5pkB1PvzgSPW7QYdBpfo2WPfhr
3yUG3N6gzuTp9Pyo+xZUuhJ2BEQorMjsKQ2CTyZX70HlNisvmGidNh0QPY964hTs
jGHdXHhOy93d0M5jOoz4SOO1OWUtlA+0IvrdUPMXznZyg9zq6vBl5/47zUHqWEMv
EzEC6CWNBkNHYjUPwQItBc0ql0tagh0EZD2Sh5nNHXpIddY9ejoDY20EisWBeG7B
1Gp3W1109eSFmhb+D0v+u3lSzAsA4x3YfcpZ5pzCL7Ga/mpH952r+Ze3fUaZKb4l
to1EuwcGg2l839tN8tjVgHMcg4mxxldcfLmC1ntELVjax8MU5ZqeA2folpSluRtS
EfYRuCQSuUsLcQ1nf8I7F2PkeqHUNHTv48u9ZDtTcKMJqlNWVG4DAZaliQ1dP6r5
c4ILzsy5e7pA/kkMSJUtDTGsMQP9OG7nJ5DrGfefD70ytFbqUrcL/dZBWtxHXgaU
y3IrOtvoPJFHhnG/AoxK52Uv34riu7Kjp1GpLyGmEIoLXolB13Qgig82ChbbsItr
BOsMPHC/aIOxr3aa4wfExliods1JknsAnjMcFW3Uw7gS4Uwd1y9deCr6OMm/j6T/
r9icYx6UxY49ThZn64bTjzaQmrDVoLczOrU77fKi7MXg+tZFAqLmpsvZdNB34Hu6
+vVErDuYuBOM5Zb/Tx5mi6sgDuRCCSF8K2MSObRJm37HFTKvhcUEgCjPOC9+1VYn
wspmjEWWTEln/l12rcWedqnSD5MDb+ddo0CzPLQvUY1fo/QKUKuO8DZurHctGz5x
fTMidTRmpl6unsSJj+eTWZ8nfEpCYR9ZImSwWiwQnygz/EPaFRmPWBZ1Y9bgrous
5mnmUSoZ1OSVWoLuQjsSEcr2xu91rF12WF5QvzmyHUzMaCpMFW9cjmefJBnlLTOl
I1ZFwCM1Dw4yfSVk7f93rmwryagVR8BYEQm45y3+hoOVQUK5i1gJWMqazsmpz8pB
hJ1lNKKeli/YjN4sxQZURc7K7PcYdKEZItbaKxq7NAWPactub00WEU9KOvegT1uL
BTvAb+XyaB22z+ijXoCebV73F5GsqJvLXeb6XaM4pzc1sp4E/NitaKhrNKZ2+2AE
R2DIPDRjrCZJ2i9zSHMWUFVeESYjLuJ0dpBSqz0gOz+Clw/JOm2sc8O2IlV0q6UG
Ll3lkul+Yei7Bam8XWDts7WHbOwgwISV/uS4tedMyxjvd0Un6/bRwp/TqCAnsM2g
Nj4o/fI+Q3GfFiUb4CtonPfWSy/XjWIHRZNmlfvfH7hUxCpEGLN+1ZVlT4pMeED/
Qz09XQmtz6Nm0H7TgjvCdh/X8a9Kn3Jn/qZ9dKvJKbPuqT5AYPUsUc/3prEPzXJV
XCoEiitKU9lsKfe7wkt8ObEYsPUg5tox18qdnxcrdBBvKn7hYfK1x8GDrhblrNyr
sDiYxwDCCdbeCrqUyw8A9/SGs21ntf0DpkO9jEYya5MzAlCAx1j4iOj001BQIb7s
1DQ01OQv4H8TtjUzohKXnPCcdQ8mxgkdv6cU8rAZNETm5xGTID7Z02kYcqenWxLD
OskA2UeRsIxC08tb/ZOscRXr5okta/IMdPbI6k8G1qgu5EtHnAAx3zDe09BVOkWR
R800U3uuDApbW/G5MC5JeiOG2Mikc7IO4zpTw6BswRSuievA/l8JbOQFK92jznSK
dGW7yS2x3Z0Cpvbm5A1c9h/PqF7hOnjmFmQbWuxYSaWoFhsYUO72mw4n1VO/EbvM
krvkw5nkoIHFY8mvV5XKpBjV1GvATvexBZYbrl7hX54IUNwv9PzELzqjQUvfTJ9O
nxKYGlxFLTipeWtinJBQ1hPTZplzFKDL2BA03aCFSbcqRWiKHuRkj/X7YaDFMkrA
1ELsu/PfpneKllTK/VTH2OlcYcb6xsLoUcEFqRHbkni5XHRbocL24EERWEEz/ixh
YtZ/ky54TN70e2onUkbTaFJoIoyZtaGOniw+x5azhqQt42Jf+5Zg33tB8SpNpT5m
n3tLZUsWUUXLSwBD9fDTyDya+ZulgrQCJy73XM5u0ubU6sEBHwi5Gb4cU3fEEEw/
5zpNgO4oChwRlq7F8VnGRx9UmoAs7qMKDVqXpBqZUOYqaEtbQfFO4zhN0nIoXRYs
BbdSWnb6phA9G40phcwj4dfOpQE3oI0JsfIB7XiylhtIHz9grnQLS+Aey/3voMjU
VxWtVRDwjNOi3T5PaMcuML4nU2lX6lbHbPhUSbgTB/Bc68tUpHtapkcwYlVn6FFV
iPoA3BkdcKlumsaq2xsuD8wbKwEQbJDzsI2vkELSnzTWlL64vsXaOhypqIN3ot/i
3/hzsZIHw8+fSOjbK1dpiaT7ppwg5NzqP0LrzsS7wYN65t0O/SrH7vF2J689OU/+
RGd9XvW1RcdqVPXOtMIGv9cX3p9Q1VWPOoEI+phhButljyqspjktI6JLXRiXU1TC
EajXbWSKJxvhiLeR2ichyxNpE/50zJ6VXFegFiZXsna1w+Z/YZ8WPtR5qiAPvufV
RIl6+vX3df4mqs0801O50fXawViP0uoEfVj9NlE4W6pqQq8/Zv9kOsJPahDc63BK
rnKk1qL5WQBZgXyFcPAahEnoSe2SyRqIDkuaecAq6hYSHdRjcRWn+y7Dpcg36fLb
l6yXeJsGcIm03FCskOrSqwn8CnY7aEf9T3FLl0DvI3vDjPWvdUvLhHard2yqqPrY
pdACuDDZVohE2A9L5T5E59w1qu7kKok1cWjxm5TY/8d2vkObo2lYsO8h4PkMlKs6
FVHgA41Xxtk2X7jI6MEygmrau8V8PA08dyTU7ptgYXOn1ffF0NwV9DKF9Um0NxPA
OB/SdD7SikRp0ulqohz+ethbEYzUC6Hz0Zip24keEZpWEinB016200/DVjwFoc1I
L+pKKFiOpgQ54rT9A9pr8RBi3N07HF3foXsaYZ+zwZ9h3/g2HXiRmUh4/rrV0Huc
jgcJuqby+5PTlDUkQoJSrm5I167ShgpdiNNsOvAw3WnqGLml5NMi0ps33xPWaiXS
MbnO1KPBbVmD/WONQmATDk2vaKn9X6ViCr/LZCIvbFG+rRhSafmSuQ2lhDKgt9Ty
ZTH4Qljc4NHCe3CPTLDF8/n3I6smQbH/chP9/JKElh6Ba84saSIcY13uT1mMytUd
OHz0yIyA+nH8Uh8mFatk5JyZpFOpbDqjB0te6iSD7YOIJKBZymN604eEyOswHPgq
SSPVj9AZcYm6E6/CVI3ON82v4ewpNMi+yV+p63KYekmP8ht/uoPZn7y1hvD3DG4X
L6ceQ3sGqrSgbnAVXoedv/+/PDREcUhhT+iDOhDw7zbVsEiw88BoQxbFZh5itu2z
ym0yoHr2kv88TcIqT80j0IicnQmhY5RQIcYFPFqCBDF5YnA1oZpPKllQdILKZPfR
VQsB1EDqxbKZiQFGz8OZvYTo6Bz7y4RdLMOf85DobNzg+NXObrhYoiuRVPh4dCWQ
q3K4eN8bszdJQJVCJu91MbSSgzC/vqtuhRqheCH20WF5DzT1xlxQ2GemeDySPxHi
lppcZPbSq4NvAjL8xTyAM+V7zaxOaioZ43nGI4uXDEKPd7KhA9pZOcgdiOa40hgM
ZHyoPQ5pD1P07nl5aFgryYZ4fBaGTfJzHpsITczqKdpFhd3aDTfuYGzO3cBL+LO4
x/IDTmSIYns8ndwEscS4dDDtex4oSISOS1z7JpJBv8IqIZJB5rYbNB9yDIT4xd2f
IcUPRjGis0XM5qfjtH68LT1M4dBKLIiQK4fVPi8nw/FbsBUWrw2+jDN2JXe0VtiJ
BoI1QW90nC0r92mDcU527lEM1D96jNqvXWHsf/KnznEtOUsJbw42BZmN4s23+1+3
xMcvuiR0s8nPreZxwu1C1ERQs78aQLJbNqaN83WV112DWTCCl/DlwivML0U6qw9E
QLTKXMJX0szRaWkJcwUErWlE8/M9pnXO5tKhPcqVbO7Pz/IdYhuwYNuakNw6XOW0
BEL0B+xvhdU8g6u0H2p892XunLpEj9CZiRzsUBhmpyfp0ofy5IZzIRxL+8GlzURG
e9F7KRGFrX0BbN1kxRMz1N1BRhu9qkOYYD+JXPWtXm/ljmY0ZYb6cCjDbo10ah1D
ci7EeUwl1p7rl/QRinIzBTs2RY/Squ/hWlbXS9fBjz1b25pic3rgiuJ+hhQciTQN
2VqsIiwvi+6Rt53WfLw356dg/DRgjNh0+9ofavkhyBliX339+aQ/0yPZbBL3alvO
4qj3f+lzZGKEnFMPA0sxt3ZBw7hMYH4KN/SFtRx/nk6gxkoMrVSxbcQe21O98s3Y
HEGz1y2MCmdcTHbXyXW0RGc6lgr9jjBU0DHEGOwENmDv14BVODFR8OIJ2ENqP4AY
0sN1BE/bZDxQpAy4j++7QL2lAMNpxE1bXOA8FN7Dzn8e2Taxrg9xat5gDfyu3AVt
/8cin4u8AGK7GW6ug9oDUCV75QYOvX+AD6M0QZmavRJgaCYw1ogpkOGfOQQHo5g+
52x6V8UnOyQ9hgtJj6UCUz8bSR4ZyYK8TjRoECvt7a0JyywJVmxaGMDigXi7q4OF
kNuKSqC+ufu4uqVe0U0Eev2ahUOPsDmzx16oMcn9t81w3L9M7DfQP+aXNedPdbq4
PXxejZ8+I+k4hL5UzEQANlm5FZVEz4qpvWn8++ioXocrucWwfca7Z/6d4ZT7kPZm
MFBBFpN2C7/FPO/WmWe/i3apZaRPL8owDlhqku+NGRrwQP5MIkQOhtfIT8CA9ZaK
k4IFLCZIncmRwhB3rFMsTfndkx9S6KDsAWRhrZEFBlh4ZPj1I8VirrIK+z+/Vtw1
6qbuXH92saJcEvbEde/9BrtJMwYuuEhyzZMEFRKorsAWXuxQNrEP7+TuasLkGLEp
WK9LUrM2mkfW4sh/EZWk1c6ONnU8hqrWA9svJFYaby8Mz0/yreU+zkD6aqY7PVpC
7334L0jgvev9f3+sNkg62O6/p+7Hf88gUbct8lZrduPEfH94kDJMqBdZlJQjTcCX
ViySENcWU7vS9ITV0V3oz3KsQMIdCLczt5KxemKbUvHYdNR0brM/Ye6bZL3D6Jw1
r1X3p3pXIn5NPBNuii3z+JtBkmqVB+Y3QNdujnvtEJC7RzeuklvdMQI1WYcSzOLG
wK+vuTOQTbYQNFg0AIynOqlEsrYX9vS84UWBbOLmZEe5t4Nbs2OvrVDufAABXjc0
vRnv1nblWgcZGTzMc7j5LcbOHor/rV4SN7+89osoxbJpBifnzmAj3kOPXzCsGr4W
Nook9QF6h/Z2on4QPL46N8EcRwhVlV0XYsXOtWjN2ICAAu3pJIVLu9be803GW2bL
X6ZzHMsVlO+n4ycatvI1JWm50cRrJPvdPy+3QjBBNiVIP7KJOQqAQuvyaEMCXQ0z
Jwl9q61NK6dBea5jQleojho4tCQkov8LpIJ/HLKiqRMq0Ksu7Mc82kpvZUwo5c/i
MzaEysyL+O7myWN4HkAhUPuEg/uCSL4jaUqNBZDSJkERMOgdQiHfZidxNPhWwJ7Z
/RWj2hlROPSmmITX0/GFFVpG6MNwRtPVKCXIc4cZv6gUneqV2LT62Dk89bMTUZpm
0xYOOsYF+w9jZh741JL/vFPqBYvMI7FPt+TPJ9vcJpWsvpCL4sb1BctBuixQ2kPF
H/9TOaqub1FG8Eb1EMJK2URSj/BoPcHB3aVX86hTNZ9nu8lEjlrS1dXcUp/V3jlU
K/uhHOnw2WvZKhwO/a6JverY0F4N1WIXLhtCDNSafvTsOg4IhJTP8lttYynI861z
DF/p1NzHATRHmYWSCD2gYW4k+/CPCI/30hNuHAhRc7lY0M7rPoHJF4TjeG2MMrhF
HSBUk+Y0jLdC3pmLoirMZE1LJWe5/BgRs9xia6pLtWjr4Bhdak44yFeyaiLN6Wyh
E9ufvrsSlVZgn7vn4Tw3aLULbtVyVxY3wu6S28UGssHYA3Yv/VQ7n2YmPv5UQIz0
Idz2wmPvNCaQe4ZSjhRjZFs+Ehy94HrWMOT6SUk0OgV01Gpa1hI0+OR+tst5w2lQ
3RNWfGi+6YvZWp4aY+MYtrcdR23jZfoTSV2Vpe4XxI7mLOlaiBteOHQP4ntsF6Hl
Kre/+YX7tVtWAdik3EqK0hkxgHvfUYMcmvEnQvjsao7nRCpvf4pN2j5tc0KkhMmh
ZTAeG/X1xegfq7s0wvWGgQH5mRhb8nUFA6/NQyH2i48JnM2RoXyUtGIjirStzrvm
A7cOIcfTGwZgxCD5WjQCqxfEGB9d0vIHYv2HSZ1F9haMyL+mPyuAndioHW+7snfu
zAFPEM/8C4fj/5SwIsrvsAwhZuJkuowbZwpYHNCeUGMEiwYzOU7EmwkzpO85AVOl
3Szg99Dmu0wRnUVNs7yG5g==
`protect END_PROTECTED
