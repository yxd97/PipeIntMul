`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aqR6z8Z/9L8enx48D9szToklNi/IBr1zuI9RSqTNJwTZ0zh0BvUSoDLQJ0Vq0QgN
KzIkO9KFUSxxPritwQNit+bipx5TafrKTDDQ5fv4Pi33TJLrJLn9l47VuhXEGzNY
FSGp0+Sw7QOFJ5oCNe5HFFYsH9ZsL8CeI3SIdNoDQhDArd7LawFWimYJNhYmdjG4
yNhMKWjBOKrTWdbx9i2CXrWQNOW0A0vF5KSDC6nsbzVbge8uqZ2BMnrjU+6AKbpt
BPQkLSsxCXC3rIa7TiGFG/A6DFdzCtxqZIUY5JNQh8foXAa+mHDP2BLTEdM9Dpcd
exYvcvHbqv75bJVABELwvA==
`protect END_PROTECTED
