`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qGNwMnPkBXPs5+/mf5PbAJ1r6OL1PXkgXeY815En+x7sAkoKjKom2qFQnPK+jeYa
Dp6QfPEmmay+gbyVZnemIo3j+MUR9fZAWmJgvvggoW3M3euMDX9XQQ3bPLVW0QMC
xqxsdnTM8O+rP9YBynCsGMNjWrxDOl/9/btZ1kKSwwmeMoaR7HJOuRe511EJl+wX
7GendVGyuh4LkM3nxi+2noKCeCicAtGCSzf13luDYxwHzoR5sLoCSWs0c94zR+lA
FqW8DoNPXOvCMJqmfHTqfgog5yiVSXOjQtmU1LgXam+WoRDpNJG06Ky3diD4/XgB
lS450XpfhE23hBVQKqBxDo2K4TfNTPzx1LJn56iXhDebOlcWCqOk3BpXLiUBmbNb
SHN+29t14UnJ2VTC2AsYLyN6bHcueYf1N490BofqfeeoSiVQs4AZEUDhanvyMCrJ
ecOQloeRRiPkwVanx97WbSEzfMS8M2vW3PvLbqbqzVCJBN9nd1LEeKCIlUF9fue4
B/0jFJhUkZrn+kTcvsaedvR7Zl7OY0xGD/sE4tahhyESHOQnhgsx91fXOOLmS+NT
g47TwmGLnABLOWz0NWlPmUI5In+5rYmBuGZ7VPZDCNpR8k2bcgZlC/QZd8hjkags
Q1BJCXI8Y/TzMCNLb+6Vfj1VH4QadkWZTTJmFN/3MxaILNLIF+Dw/ZWRJgSnjCnh
jyFqXMtX2BjZYU2A4NIuaoXsudEpQcg21OvZtKODFD5qCv0dQUGmkFPkvDcZhWr4
Zbf8zAb3tOEZlzNzBCRT8Htxw9b447I71zMHhRoWolRp48zK898a5dyjwq5lvv7J
67xXCI4uBOekDwjfQsRS0rQkUpWdftB0HLfqhFNmg9GNZAMCxVXDVwiIX5X73e7K
PVms9Gc/QIPI4VTCbFmVZIOqvD9TlGWhDaqHT9oN47LSJh0U37Td13KKpjtpJ7AM
K5kULv15wwqMgOfg1mSZfpR3MwkZiA37seeW5dK51vq4XksXnXE7rjjgH1GGBWUA
BzlnRbBYy/HM9HQrlZ9xiRe9igy84998CbNW87e5l1MTXIybylmEG45KZ1nyywN3
iQebTn3mHlPloZedN0BSpr8xoqeUaSVwozNjQe1wmourCfKIuzMXBpfSQdlhMDex
tG6yjWln/FBWok3D9UAAGgAH6HDEAKmBngwJ+/9iiw3iABjsGexUcG7/tRdgDmH1
ki174uBg0bjoE7Dl2cuutwSafeAXDdG/sIAcwSIbZgYxhMAWBH6oytVnd7FA0bu1
/zvC+wF9zdY99JJ8eDL5tTy1Gvk85sqoVNReBuGXSoBh9VDzJS9r+v/Hb+5GZmXV
JZFMIOVx9OSwbmf1Rxdhsadvz21+A9Xf5BwzGWJGHVB0ngvbxRSG5WAAC1OAHZcM
XKJvGjCqWOQpB5CMteIrwNcqzPQ5iP7dUNLMv/4THlgoIqcesROCm4a59DnjAZGn
XJN9fyvS+guFe/vfRcIU1/cxkyjtOb+WsbA3hmHokpqMK1pNWzh6wigeZTI/oHGw
n0XHoaPNAOBr+iTgTVqjpP/SOaknteCH5OZlHFXjms7p99537YfQItnQ6xjKffPo
3hXjZXdNEvDJd8zCD7geU5iiFbVZ6m7hzoBfRZ1Ct8Wa3b7twrZiB/qEpntMcUwG
pEZdpzEzkyumfnPmmRj/NGvfTEaxMYXoSdirSRiLJccv+cliHdo1WId8+r32KB8G
pP1llGnSmoliEtRjjsXskmE4SUbNKiUOVguGeTqPbUL1C8L+Wrds5jf3tQuUgMPl
ISXmBU8i0hEHbjxXmBUyuIeBm1gkygjg7mu9HII3Xad9BZLGNR9AnCol/xKxwpYR
5rFdPspCYjjUc/Rczb5YBmtYVD6ds4qky3klL3PzO/huKFCfFjxztAkFMPxS9BzU
S2YF+RvPBGxE+FTqCw/1KOvXpXHggDO0IjbfyXQaE0F041Cww2Da4wvfEXNamjkQ
ZEfQ3vOWFouHZTs/xtPJh0FMJ9wCvhM2d2xVeuE8mtmVvcaDdpgQFJbV5QX+jJvA
eKGCUK5KVGY8kwPGoy5CJm4P9acBkj0Rp2p/PbnF/bjjJ7qaeXKJUjuHwYSNQ38G
NSmB2EZjtSFE4aD7NesXuCKMKNu1jIt3F5fCK6Bdg8JAl3XaRgsp2N5ksd0fl4bT
xefWYS8z6AbCAxMeT9US8Fp0eMh6ZFcG59ZeXPVJ9dxqFJECOWTdikqs4y0IE6KX
1TUGgsENCZF0TMWftRlSb3RZJVHY1wWm8Qr9CXYkYpIride3L2RZdgjXGf7JsFR/
2dWqOH5qbdbYwXnl6kX+xOgeb/o1hlr/WzHvGQvY6j4Bb2H2HY7QVnA92c9cVTcB
Ll+ziW4pNj98XdLl6SIZGONFs6kBc1Jt9KiKnSPjwXbr0TFLAR626UoczOJuJXca
0WWDJp1pV4jK/XVgW7kT7nqeRXBewyV0VmYGa67PUS+G9yNZKHpiIwfu4+LikgYK
1b4DIYl3foYQ11F6yg6dLc7JtRIEDbPN9rsOE9blb5Zk3O9Dbmk48fd1cvVipI6a
91ERtPbhxxqPftL4J9YS2gLfDUr2/fKPuVJmxeNqEzGqnfQF4IiRyU7KR8WtUQd8
5Bc/xsl5fCK1vRsVtDr6dbmNKziBO2q5USvCUjJyMAmAnpFreMk/N/Q7pyNu1X1g
vaFpFeiAvmG3Q8X72HtHlNZfCDGQn3QNYJwqBS7Ua4KqTx95+Q+PaOTYiubLKhQc
Mi0G8/oKu9mNhnAXOfFq7Yykdx7q7OjA2BBoo1V2zWGNqSepzCbHZbUXOtXbjmgX
Gtxv15lztDxvkmKMvtuDvV77st55evqY0L2vdlhCXvG+lyZ7aUt3r7YWEyBaeNn2
8ZaB9ciD2GC/2Mfffp2RoA==
`protect END_PROTECTED
