`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6fKNrbNfUQZaL72ltRausm1LJLrvwj54tlMy3CqTVSAxlW57P2GfWJ1BNUqh/CpX
VD5fn2XjeHe7RFSRsxN5uhuoRhKlhE3wLvUraaL0ZWtFPcZcl27BKf9IEv4Suh7K
JRLithhvQ8AoO1kx6sbZn7G/LggBcB7jnKvZtn9ZJWyJ3Sc5LWtWP/qGlfr3xvMj
NMtEv+B4LjzrbCfhpvXOEnvIyZ4gWT8YrVY3zdno4lA8X2Juy9M2HivnAVOcS7Fp
vbFknjpg2oWECcrurJ7f/S4LFSl7vP+Gh3mlTAJPpQot1FptwCs7+yYSXgIivqXW
2V7coQ75OzGqWnBAMddd+TX1N2keasAj0RzWLCvapDnwnycLAbqOoJzmELqP5KBv
D5BSZVE8qFZAEIdMvUwP/K/sDh633IrlaOTGkuNAR/ENEfO3UcsKY1Gp3PO4+sqQ
OlZjiha3YyD9U91dN4usQ0II8MpzU/CJ6fsCoD1YtnMkp/MtvgVK4FAuN1TsKnzK
L0gDvFgDpiFOdycwvemq23T1+KjrVpGdHgn1MxmNzk7ddNcWw9tb3O/PeiJGAU+U
s6XY3+abHYb/EW9mQqnpvg==
`protect END_PROTECTED
