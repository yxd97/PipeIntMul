`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5eJ89HZZtxbk6FLXTs2IrG2HjvPTk8EJwNSe6575NV3wHmjgY0d7HADmpnsAJj+6
7gvP9/VRPQl++y4UqE1RQPWLhm6AD91ty3PT/2GymleEEayW2w3Cn/nzTEk6r7qB
Eqjid49QX2ixYdTp7JHnlBpkG+cPYAc81j9cABkDhBkbBrnwjk6gsOdq+sHOYeho
sg3JdWAEUz+TDau7gOhWKQKeVlktl+uvXY2LLrGs4qNbkmT6NgiGc7EjZXfA940J
v0vPmDBiEK3xqtmjwOQbqDZNENmRnwCNE9fAP0yCr+tvLBiNnaZONaVMTy3QfUfo
qoUQRg9OMmreV6u9YJcBvoFHQHUN+dRO4IyXs227IKHmMxFIoMIPY+EhIga7nvm1
+hByz8JhQIJLg7yYyI5FLHSEXy8HV+8eKEx6EZ9v3GIuOAtZNeooK0MNp87fPBRz
36P6Z+kWTvADyaGpVVXpX5WlpCr7fPYsVnB9P5oeAkzd5HXQSjLS2ZE58lvnTCSa
KHzE4NqQ1HGO5ham678J3PXFYRsC9XJWGVbUlqNkgX+5ceRULNFdRyXuFVnw8qOn
YNJ1LNPA6ttRSDsqpm4AWnYiKIhIK4uV6mAwDZ1QXaSr58kOrQwRtlaoSv3YMeMG
ysg5jNy31XTQ0Y4Go2Y/arwaBplMybcYZou5kOCJ0NYgkHuZt3OxYjH2TxD+rCV6
j7HMDIbIaK4bmCMGfJiTGKhZlzCAA/XLnvaP3uossltaxqxrm2sLXIzR6P8Carti
/5UM1bLfppECBxny7a+lsSt5XYtDckNMzdFqPLjbns/t8kATT98+H6WMXQE4WkeE
o+Ao5SdXM6sKUyMlv5QvndnC0k4Yh/rtUV+8Hy7czD+YhC9cua6hXTH9zyAHAdfs
jk+ZicAC5vNgYD2m4nhZlUxyV4dow6Gct50Wx0hYRPVS2C7Fbx+RKZxT2satVSGk
RxnpCb+cLOdwgEuqc/IgFlzJ57zRiUDXKjeLCyEx0Q39iA2YeWHRVSO3Eu7zGfcd
x30irtMhXh7xjbEkJa4LGMfJYfFMqK0RDolti3wAvisSGS8Zcstm6YTqiqgC13NL
TeEUsu08AJj6XQMf78o87FKAPIvDFxahw2AZU4K94HAX3EJ/jyGpn4aya0j7j9FQ
E8wvQ4F3b94g7cabVwxszFI+QaY9XMzNqgsJwOYHDrRXj4KEEE1LNGH42SbVqpzN
YkpheC08M/Kndg/8GGDLiWbsCh2x6WYktOB6p138ZNOlXu/4tYmOqrxd4EDaO494
museSIOQXs+qFrvWX75tAzNRBXXfTi5MtVd2SegQ4qjLjf70+XmiE3bZnpaB6yRh
7wBddclbG5zIktFgYD2yvrR2D0rSQfXMLWUNL2E7OWYCMYky/vSViriOTwKynkFm
08LDsCjkNf2EcaTJG/KlqA8ubafQy6K+WFu7myd7SFQErNQJf+4Dg4iFL/R5U3in
/I7/8hOEZQltCSzOr6KZRZR2rnmaoIGvHgQ6qwqcNZXUwXYACeJu+jNZFeu34tnP
V2srsWKdUDW4gJFA1ZCpybYJcNDqVHS1HBq/wqiM6xSzgsoobEiJuUHvOdeXwUdV
1QVL5mUy7y/g+EW0TMXZlCA6jAxWFkb9jQ+HaO3mYmrqno4qPy0DRatrrs67HaAB
qTfMd8LLkTVH+raLr07aKllHsthoKkygdzFO1VdRV8F7SULC/2SPlDSp22iZyk8f
bSdS2tAEU0eQUDg94MLDBIjjCtzorafEcu0z7EnDUnV0Pga+UeU5AqLSza0CQEgr
l0alT5j1bmIU13dhKNEcbZGw6qx5/AQxE8q6SKkiACXkWsA88Axdzrx6xvITM/ac
Rsp/fvujY/iOvvTTDhtnMdZfAWnYYUXmi7AUIYuChF4ClnZDxPa7Gh2pt2srFElN
3ENbNerSKggB7p6dkrVPbX2ePzVT9lJI4ux4+DZOLNXutGqTkLOx4/Mtr2ynQQ0N
HKHfRHxl+wvxl7phgKYQ/Ea1bScduHAYJfsnuSl3o2XmEcaWQvL2pg+b71AutUlR
nM5jyspjd0sia9jcld08y50cDj0ywNjnKxitwWZVuLa+LQNBda1M/eXAkkTfCB3r
NCmNrhXqf1BxElHLpFvAcS4OruUGLijG76gNzJO2rw1G7ksdjABTMq7j2trA8QRB
G3B16Dhw/oRnlDbmfhGfFvGr2dK8Nm4jIRrWhkUAhUm5cz+dKI5+nulis1DEPACA
KXkSRFGEql3nUHv/6PTGKip0n3yhICCDOODg/JbQYcU=
`protect END_PROTECTED
