`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPTYrdbXYuzRI/rWVa7i4zjQdq/Tjxb3wZBaMUzbKk9/01VRaQ2Uo6iL28mdYmC1
T6KnD7Uk90ro1SqZlz5p5VAO3PrdKCttXbIg+9bZWaP4jupjFdSPKpWL2lPbSifg
RAooFe8Wd3yjIEtMcDnmwTHQX6H+xKGOP7m4Z+q1gP+5ttSisM9G8g9u1kXSAJ8+
NkToZq28Jn+J6465NUq3ULhmdbQdbZNbjm7vcB1+AgQHJ31KF1+Yvb/qK7U1+GKy
o/6N03RTB9MtCpNudLxfTEotr89M4Adrk0xnTg/8w5fGu/llgRivSeS3DV7hMU0N
e3FoNVni4cHkJ4OJiXX7Swll6K7J4n5k4gxDZP1eil2z4mjAoWc9uclnPkYXk2IG
vjC1+fmB+UyxDNlSfoCRjbjz13YSXDp7EFBfPxGhWY0=
`protect END_PROTECTED
