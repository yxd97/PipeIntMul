`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afxAk6Yk2XN98VOU58tG9VYTZpk8DbVW0A4t+1lXss1iWnkU23UtYcExDCLAoGTP
1lJ2Bo0WiE4n7BLrf47dJdnnJ3c+vML5OoFBRR8jJJvAE4d4BkjojECNCgoQARN3
RuAPTybExplk8i9y3G7tSTynshdMXjm2G9XTK3EWjUcWy1cm5pwDV82Y/WEq59r0
UkUEYVvtXevfe7g+wIFFGyRqc9QUVPMdQscK9tISDAW04ISzLzVPZh9d5sXZsb1h
vt7C4RucdGfR8fgbnAKEykfg/dVKu87aik3AYoAmyR74LQF0mEjveEM2pQ1AOUXx
3tAeJg06jtMrA2fLyGzPOk+jK1FuPHNXiWPw0Y6kPGZiXIBTmNphuLPObDkrxJZi
zpi2eLq70BTPVMH/VfkXwoCQQjDBuAMyngcJRSo50Zs8F2nS+1f6JvLCTHdY0QNr
`protect END_PROTECTED
