`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
faSgsrPAycI0+FCpiJgX/IEeRj29GMIDN8NU7huS2RnIeruRkOxKyvcIZEqENMYk
HKtR1yWOc/9YviyGXE5iDxqykYZ/N5yULP1uKP4qxw+6uWDulUea5SjQkI5xx9xj
Lu0HQgVrVtS1w3FTlM220kyppgpKF17Uu7i6U4E834+dRdxJG7innNpvUcT5/1NP
kVonOpqmc042+ZC2MR3wVE5ivIMUVdY86cv6BPTB2kM0NAQG17DvfAGoClyR0Ejh
9IkJonKeYw+4OPWgGD9a9tC0uw048WB8Ht23UxrMdPva4CEp/wZ8ygRB7c4EFAOw
stE8V6D2qxq9WIrVUvXgf0C4lsQzXq5ugaRjLcyyBe4ksHNuiEYF65sBtHpOlpI2
NZ3hb7vigxf1m3ZjR2qy2oaClSm1YB1qhpMpOqaQ7PWy73FAS9swrcNqMJcn9JKy
a/hVAeLFfJ6+s06WZflH08ukm3S80bkMHMBhgjpJF02YDKLxP8edgPByGDT4WgaR
Q7zzrYF33UrSp0p9nFcY313p+vZZRsNyLI5hUpeEU8fq3S66vyAMWHmEqZxCmoUe
7nEFuKVuTWkyBDSfUrxu/2U794yqSFsWJShCFVGwF3H5tn2AL/ivj8A1yLeI1wJz
FfX0cnY36r3owFVOdbNQWKBuVGwoKmwXHE03NqdycO94eAk1RUY519cnO8r1n6ry
AViNJk5NAzg/9oym1O38Tb8zt6B6hFzOlDiw4hHZwLY=
`protect END_PROTECTED
