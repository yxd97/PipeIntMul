`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
24IPEf7IW46eL7RKnjPPP+vlIh4LXJJkeJ62a+HE3b0ZCD1g0DRpmnLdkGxfB4+C
xkxZFMlpuYo0mNsbBGg54V5bOkxH/zmZfPikQQOmM4XuqawqHaFMzr4Ev78T/w0M
6W4KNwI61Er3fDhsvcaaa4klQqkUPEHRyFg/L8hYo2OGiO7jdB1yywy5kINApbhB
y5xm+EwUtV5UzwDVt9394vlseq9xQaeiGYIjQExZEj9H64mw7PCE0vPeJBeeawOJ
mmUqORAGC7pMS/RjOKUKFvTJscKIrOv+5e9CkRTYq/P81kOBLyFC4WATmmnF3EKu
0X3zoabcY6MEs7lEKxWq7OLT5FexC0Y1JdlNy6C/R119LbePHiINKD2AdaR0hVlm
pfOGxsUr5DE/E+pp7lOZe3xA3JyQfwGYZGUEdYyAs71Uh76gxteWxmBBxOIAvEyE
AiSO5qGlwNhRqst75ep58ILks0CH3nyAcHnl/u4UNMMibTFmOQ7K8SplmK7h7ltq
zeYV0gNA2dchSslU4OjyJwCvqGHQ0PsJLwc2vSdhCREJIDE+icujTl1TgOZQd23X
oDS6whBXCyOXAgMpG8tOtH7vzcXHFR91ggIzBuLv9qfOPiubpAQtam+WL9LjPT3C
508FpaIHzfzkMZaZGPhD+Q==
`protect END_PROTECTED
