`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jkm8K6fyMnwsI+1CEgEK0S2FBj1bl2MjBAikD9WNlajWdjqk79D1CRq+B16CUfCH
GCoMm8sFJmiBJDan8V5y56twgEi47az+WVtnrTfCdlcFNI8Vqf040saGF169ZJYg
+65GzefxsNAKBd5HcE86m6FrC8KkbHeKOilP7XpjdHuhX+YLjCBd++uU0MYb0qOn
IoRfVTBW5I5lOtzGxe0vC/k6p1F3V+EpSZQRH3KLh/r8QKCXhTeyR/v9afF/sOha
Eb70kZUZef+QVso1BACJ+fHqrtM536/55WGhVeAbp1X3NOjxywZsPrglIt1t9gj2
ZFNKuJ++1bEHzeUGyBj8tP//XDlXvhb9zeTNfeaIZWU2R/YnyjIUoF8KuM60zyLt
5QgmIpCQR/p9tLiP/rTRulDfwVVyygyx6lr2cxJ3Li/98tY6D5tvNFsrbR5CbXfx
6FWkynQEwHYBUpkRSBd9cOpcU5HPPYGW1MEG4J/JwKKVOkc7lgSVeMGseLREQhJ1
grUitmj2J0qj1ekH916cDSNtNtxDQAao/ZOvo82/auk=
`protect END_PROTECTED
