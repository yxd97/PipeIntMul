`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h7FJsDJJd7Pfg4/+RfPwJPeAtCqHk9MmdtrUj036DNMO1l+FQZts2FogywjUJL+8
QJULbgwsaq9WvWlY/j76dyESqV02tdJ6F9wTVYsfd/wF7cBRaNU/IaA6a4UZUkPC
uyL08rbuP2rPesceP6ofv2btQ3u5sWj6z+KvtOa8vL9eK/NsIKwSrz3frIhTlJVU
vUARdhM5v1dTSv0Z0Svjk2iN1j7p97slu5WexauaZMHTkGwHjuGMyx7Ix6AJ9ML9
o/Qjf8rgDZfH56jADefVQw==
`protect END_PROTECTED
