`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n5pAp7vX0N7nICRDWxmhpFvRVlbF/090scEca9Wd3NcqNJGUvAyTEbAtuZzhVs7X
QH1kRrXnmIKi564XyGi5HPaM2Qy96oS0+pgvKf4piOH5LPHIlvidCfOJpdf9hJJp
zeGxOhdyqhFo1JxMnewoi1F03o03DaiwSIvwnLuElQIL8JhbVif9+v/MaCQXYZ4S
Jrx/8DxcH9UXMXXGGl/2CMkQr5C4xQjMion8TonflZGVkhrCdXIQoERVgQ7dzErM
VaKAGsUAQc3h5BsebZQs/xzOogvLQhq1nUButETV7TfWgtolJNqNWaZZvsUbxv9E
D6sw6XwSEhaAHq+hM5BXDFZrzWT8vipVQLwPC6IgbYINxqOXHs55p9IbI08C7Iqx
qxgGwNGsjL1yESSe0qaJaA==
`protect END_PROTECTED
