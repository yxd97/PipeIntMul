`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5yj5o4aedN0L+Zkw9kP3+T0kldW9Mtsbyb0G+wa6K159QIQq7bIq9DjsAXRrBHJu
+kx2O4jrXmkzZBEKuSLP+JMz5MynUbfOFiHFnJBYGBt1iLQaUtMRySaXWWWaCgz3
9/EiBTYLEBt3IwxbKyWXmB9BihLTopwF3DU8vheUmE7e30sXmGzcUc1Jb3pNq26D
Ep2Vn+6nIDM/zZx2Y2MgPSezvNqbVRC3EnNcvpcelwKDBhHVYw0B7IvmmGdzPvqV
bExPnlRvIAmdUpTRkXP9lJhNTi4g1CQUT2UjOcT5Bkgh9M2nbBAdRv/m0gGRF7hF
7sPU0IDuj1f2S6Qg20uHu50yknZMTmbTCqZnuSfFHNckQ8rA/BinJJZXb+Wt9IWN
GoiTEknHehmQj8ZBJnO7wA==
`protect END_PROTECTED
