`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8EXyM3a7yUWT3rjLL1Xdq/34gIVFmEIFRllYqTuV5lN18jIF00fnPYr1l/TiNdSs
X2285AcfxCV89Mfb3qy/cuKU1r0xySU3BomcF5LZJFVW7AoSBHe/ZB8bm7OKnIW/
poUeLv2OH4yenaRODtKgiG2APsJzvfhI3aig7TcELX9kBpG3ybm+cF6EyovcAsdQ
gaofkY0gKV1KKpMvgfpsCa71mOMbLt3pWd/Hp7Vxnu9jY9HnoIVdkCiXYjYHOJ/+
lKfATi0n8NQutR3RI+HvfYL/nZf8pNLiLrKiBFZz7OPrVfxNtOA95oLe4dc+fpTN
pTdnjA5cyU8ZJPJ3b3Qc8oaCaMPUGvPZD7zpeR+Rdk5HZWU5SuPpocqR48HZ44qk
Xredbbjv5KUq3jNAMFKWGKnLD5mUjhih119V96UQOMXPK+lvAG4F4qodnhkSbtXN
hiqGhvP5by5KpvgMFrNwV3ICrT27VY4BLA21u0lftnwiwYbIbR5nFtczGYACQkLf
lddjTI6nT/ew6Z1uUjiwvZh5SiJy7+fQnxluSRLKGSedjpLoGqgqUEFXrS6lIFsw
pli7k0kLZgcsE05vXVnwkwn9xpQeiXd2LS1EjVe/BXtvl/TXfxhTUCql4tZkR22A
5Uy5a/J2QRQSGwofg92VOCbw45wKGg2e5+uhX8AxSiKWtrFxJJCn39uQrE2AT8Ty
G6yE3VDo7+odqXtMJ9j0KL5AKRWZ5x/PmkUAr2eyzbHqdjPkWEb/bP4Xd+jdr0Hl
ludnoLIOP4Bb0wE09291xIuic5lsXkFJ2tV5NWGo9WKzcs4BU/+O868h8P3oxHmS
Ckh0S2j1x6hvbwBoGlWW4zywnGkSzAE56YXhI+Xv9ciQakFGZs6FjiqiHy2qMrPA
+lruJuDAOAr7+tssY5tiGvdQYvLyuHPVaxj3pXNmW5Fev2IE7hnelIZuUn78CG13
0rMV4BsC/+v118OXDzqJaI5zFbrN73T2ghwXOHErz6+69gxNVzK3ShIxSSwt9C9P
eFYabFeJdebuV+P7gvR6O2CUK2eiQQ+sNIRyzoNPEZcYrCW2BAlIJatZT2ZxsG3M
nqeSumGT+KaGK8ncrq07U+wjMjg2H6Oc1nZ72m1cOCVjBSlFhBUTPEcG7G7mNECs
8vjIjlxj/fentKS+1WothBKQCsaACbXcdaFBxf3bE1k=
`protect END_PROTECTED
