`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Co+TqTmvxs0ythNTonlrdayU9+DSNUYipezYpMD9mWg4CqchTV1FOibCg+uNaA8O
XGxygV9g+6ZfXeQLny+2icvyoo0ZhhVJ39QWYFmAD7AvRBV4YwYDNu/VkoKbm2H6
Omf5x+pfzpXb//cjXyMa5x1oYOiL7nSZ+ai95c1ra1Ed1rJG9glFvjm16ixv5nFq
/qnBq28UpS0+yZFEiJ1G8FxgLNChjzLFdKm/CKOndxSARKCpYLYgB4OoxMk+3A6c
LQLEre/SW8mX+7lNgZPoSDQen49Spox6x/+Vebr9eTiifiWWQlWF1COX0JnXAa7e
cmbCO/odg4UgWpxKxyRLGRoC/SzihpMowQ5xC9kCPKrLzpOpwekoWOcsPLSx5vLd
037kW3XPQW+duFXFyGOCcwwSXjwRzfaUvoicd6UH2giYEYarj62Kmxs5IseP5lS0
glsOawZkrgP0GuvQJ0Qc85k8INWkqNim2KQyLNs/FrwqmHrmBx2myTphZmT+TnGt
PtSvLvGmSKBtvs2s92NGOuOxR/GlfEQrhd4NSm3JIgux7F1B5pVvFXtIUrMZHWoP
qFfXLdlq91Boi8jnR1d4HqmZ73++cWHeLJepg36eJ1ynOdOuxdpv0cZpd/C9eQsj
DxIzwB9dQsgrYVmbNKXXxK1SuDL8Zy6EJQL1qvm31PZVvVF2LSoL9gH1k52RvNn9
/R8Iu5ZKvKHGVUwzBgV9WxLGFDgD+W3pdqh5AIxZA2G7aSMdzukL6UotIViqMiAx
j0qjnCl24ocOtG0RA+wJA85gXeHF+KzDfs1hhobOl5nIDwdR0rPxw+kbdiO3TO41
tYCDd2aSR40Gam9xGu3ef7zIbVLmjV9mjS3oGvM1aor4y+Hlj00SyfquZPvB3fwZ
N2tVZyD43qD3ftmFE3HCNC1XkSJMdHhHJ/8JlpDM9h8qRco36XQA/HPL/TfJrIfZ
fjiLr+SG59asYp6LFkqRePo+ltPEx/s3HwJQGj7O8ZH359tnCkXdHJ9zelvUhlfC
`protect END_PROTECTED
