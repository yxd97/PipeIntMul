`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gLV2HvKGMmFzISTNwW6TTu6gVLEepND/bkULUE8DorqwCZhoIguEUY72hgK9pniT
WzEdqnO3VbIWQUxk83o8fOcxt83VtIroW9vGiCxRVQPKqxVWZF02vgckWZTTw9tD
TxKDlv5SxuJcfwPmaQc/X2ltvJBOM1P3N/G7iFOaObzOQDIllxALWxzZiP1FY8kN
6V5xjNPEVcXZDRFhaOGuz/TaRWcQDt0RC+3PwBe8mEYQ1cOG5I+My3mC+L/9vog2
`protect END_PROTECTED
