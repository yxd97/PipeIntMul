`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BeKzH3bM9+D6+hhwpc1GG4ZbkUXkvoDyoKGAkKkeMLwfaDWELZlhVuehKw7wWVEJ
7zoL1SElGvJw69kDpET1Oe7ZOD1xP2fN4tZvzF7eXewGfEJy4ZDsZxB+d/6tq5Tb
QTh+lR7cJ4TkumiLWRNRl1Zdfz4K+AOhBFWL9eBxb9o6Ie+m99BIGfUSsfgJsRi2
t1RKk2v3s6tsccO4N+cshSHmS/9SuURrAzyrezT367NhmkOl/lOn7S8NJVwxg3hc
+PhGl8lluLGOAD2+6NFDzFpZfUPpWHeSXSCLFjhfjYN2vY1JOGZ4YGd9xemvpnhZ
zK0YIo9UnaMhrcZLtolqeW8n6NBs66LY8qJWjVCH4ivWsKaq4tVvbvyLhQh0gjgr
lAjzj5OHLngyyPtupULrmJPouWQzSmXbvHbllmSqWTs=
`protect END_PROTECTED
