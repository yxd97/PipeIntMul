`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Ig+0lgtdWVS2WnZ0nIhQpfFn6cQ7GSVc3nEEv3IYQ4scDS0oYwGIeJ1/7OQtzf0
9yhkxqSJNXxSKyChxM9hRCv9I2UcPplQ6fiEuCC15dNuH87/VF98wEau7/NMhVht
9mjehSEyO2+uZe9RtWm1pBoqGNg2Qu/L+1If0BsRQ7UwtxwM+ldc74aakpPGEcU0
NcBgvzLpBOx9emU4/BM2/7SUx8RR/bgiOMv2959nRB+DB/OTFVoFWa6c6S0cer9j
zLJ3+Koyb05Qtovf5/tEVJ5SXv50SCm/Slozjn/wJqi14sx+HaB2WfN9mRTpgVwi
DUjsSBwzeVs3aJXUSuhg5E/mnIqTUTSpKnm6HnJsLX+3AmyzFMIl2Q5dcBbvOKHj
0T+N5GEzeNFVyJf6R3SU4oppvXMSxuyvcyf0JxIYbws=
`protect END_PROTECTED
