`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VQZ9vLjOnGPhhp1I51khwQtZt0+7+4J3siulel8ubvIaGYRekd1ytdhJg29FFv2Y
hxW/Qz/NIKCtREpxHFh2Qxjm9AwqlFIq8FgnOmlz6NM4F6HanlLQ7AtGabsOQuMC
dAoNOPegFTgqcK14Swsop2EwWwuv65IMmq1U3ecBmBnTqI7m5ghcYmuiaZWE1HK7
sDsCfuDYUji12yMEBeF4Oxo8vuceShwivXZeVBxn4ThPqyU0uOEmN8OcpXipy7Zp
L7w7k8K6Dy8hFVLxiboZhQnZgfLa0oW3YVBvmHNcIU8I7Sh4HovWWQPYo4jtgu6V
Hj6Bc/FKri4qCiZGpY8KnIJhe5IBgsBG4Q9+8x4I0y6zSKLWwFcZGLAunLTIrV6b
kTHf80BtkOCmnVbql2ZI4EthJDsdbEUCze2yTaHD1nUWUWqYkHOr2cE3WNPxaZXF
Fd5LzZFscH8D7Z5aTgzYuE1DiVRrOwhkHY5NDS+T0NpjGank4h03S9MAS9Qoudvu
fS+Q6/FQpusxEGmxCNen2qg6bI/9koPgcYC3tqi47MTXofcDFDxcZ2We5Q4IjtSv
V4oghm86sJ9w+7sZDUYjiB5TLurybS5qryO+XE57NoM=
`protect END_PROTECTED
