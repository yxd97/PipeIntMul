`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrcPZ9LCd1srRfgKtUi/PFT8d1lYMYNHQOhmELASJ8ZuLorbG+bNZrMEnY8cUWZm
XbD6yDUEwDJgozH1ZV/GxxqdiKhUdByq3ss+dn3iApAVYgO6CHQjxZ4zgJ1rBl+f
D7ahjBBZ2YmxwQQ4XBX+9f1MlAmIDOd1BqfZuiHXRCHU+9aS/Dy0krWeFZ05dbrW
/MxxboFLa7yP6xcX6SPAc+kD5bKy2+SWOa3Ox+ALImkHXLvVdYKW5GMicIUAZAD5
jnKV7Ld7lXx0W7lbRZxaJh5kO75Lmz8kPle16w9Izc9daISaL4J6hdA57Phy/fU+
Uu1mWMHDNrNyuyv/xVEZeTiuRpSJoeCTrMA1G+rXND71ZbaKaSzzC8eqWbgSDFMP
M95L9AqLDt5I4Z+x4kY0ZwPceMxOjVM4VN7C6yT3cmY4+uTmnVFp2q7WLdvj8tK4
HjEc0VGpAP4nM4YhV3KYyxe98ZEeBrwNTYKiV3dRrQ7HdttD4q/9xjMW5XxmJ0cK
ZnkCsdKZArTMyNNb+98dy+IsEL83kMOAuhmm/logMq0wKdB0hMmwV7hT6A9i4QLP
xewwqFIvqI3GiusVevBzupjq67buoQerSXIca+8RrcLFLIQ/WhebJiC+Gl/IMeS0
x2HZGWapOUUEvxP2zbaNDflfX7URXNIVezOA9QuPUl1lIFp43bqXZxuX8BfHVDJq
j/D19YJE1zL3Ieqe2PvwuDoR5mYKk8gP+TtLLOcgq3AmHtBiGQSlXgkJzUN7zDTB
MDXGuQdmApgsRGlyUfF2iJl+c4S8jxZXLlFlKseXugQJC7nj4Pu9c6zZVvHZFjSI
QEB1VEv0knmtvsaI/+BVakPBPBbYKgLPmF7Qvncd4+MV8H7jl0E9geW709jG2v7Z
EVa5q/XrxBW11zccX6PtBc9LUCSx0r6NDXRlNTDOkG99OT10NWqvb/hRFACXtowx
XgxNc3+dRo/W7rCTfJZ+NgoKv1cGun8LcgidDqia00guQvjGsmbh101Pbw4m9GKw
DNEhEDZO7tUPskbUBSjdj4HXRD9hHrPHvbWE/i+/pnMSpQMMN0jq8TtFVV5+qdR9
68uZfn3rkZt/ldjqHt5YafY0XpQ7SYRgHc5l1FLFWvEQSZoUsc13hZe+XNB1tugJ
C44epst2cKm4h1hHQy6gR0yd3gY4aVOcdGzTdC6Urei7O00FeXSAVluVAQPiPvNf
g72IaOB3e32RgAd4H/V8IAJtRoCxYWHimX7gg2IEbLpYpG2dIO2pOr0jpDelqz8o
BCnoXIN4tQAmE3qu5a4TW/ZNrePUImJCj12BkJoguR1dh+PAas0CtfxApfk6fJa+
8WQCKdndATnlCOCdu00t5kLRPzwZ3zP3XkmuVSwflXZA+t2MbM2RL0jhSDG/YX4V
/0g/SV64CzZw/vUrc8WX0lrbf8EOlwdGKkVoMbtkxLRip/Sa2YerBUIFsA6IUKgb
aNyEx1AnXHux2y5EWQCMvcziXmQIU3rGCU9ZHuAMObb6DR7/X/Rs5EyT20HYT+6J
KZj1gRF56D3YZbImYQ+7NmrJV4JCyLIuZn7w2AlMpvcb3js4PE8HQZqFdgIdTwrd
4UDKsUQp3yO1SCTWog6B5k7QSrqzIj+ijaektCOVToN/8LNzeBfqjo1ax/jcKgbX
58txSipikPIr1GC7BANXBJBYX8eN2Z98z2zmN7sEAK4jZudpkZSZec4HDKR2eATl
YdejCo3DxC4Q4jV/NrPS8vgE2yhSso5gO7kJkR4XQ9Msk1bm1ZIJ70QYod2Wy9bg
IT5F6UkyjSUb7QkxMjHXecLkoKVyBshfAxRbys7jjxljGiucnZGwYJdHZDPlR4YM
CIoAQ4NV2SR8jKC3KLt4Q9mJjcL1x9D5peJslsIUcibKQfQJ8NJ5guK7xceomSxE
T/2OcTGCfMxC9R7DX18h3yd7vuISJGK0wyaU+KhP6ulHf/bdm5DJeztMguXvkP4f
/J81t/Bi2/x0c0vbGL5waTdvbnoA2XGltZT+N0hKAnYNISeM9+9dGJ4JBziQUOZq
q/Qn8gyM8+up9jqoC+gCuY8zz8cBLZo7JgrXl+f867gN5zehUCFst5Y2bqY+llqX
0XJh8lBhA/KMsZTEZMUOC65R9upHxcS3gqJ425BTFjoP0TeMROoUt7gyR+ZZDZRu
XLPEfPzCWI/Srr/KXzKvAW7uPWHod7dmGJ0QepMwAWcnJ6NcZENvnwzpN9F7x9je
pmABnLWtFPFkFaJlctv7Xtde7zVsoLEZsVlXNqpBKwPYyN1oz+TQb4n0NdaBNeSH
V7QHX8OduU+GGGFRS8m2CJ100muev25v686KfsLhSikTVNTuTAaPQSN5PeAaFsIq
DUQpsbc36dPxjoNp63THCh8MCjR+ItIFmb3SUemTdGYFrXCLbrVV3YHfgk1O8oJZ
HwqjfPYroCkN3mxvVGyv00XqMF6bvQVa9prDDi5NQ9U8QB6DfUX2aVGIESZ0GVZV
wr0APmeLOWBdrEdL2JLxc5hHmVTGfxBGa552n9TK4ULtyszM2Yu29cDGWmirz0PP
4FKw7tiWQkgEFW8EPrZNLbwBK3d8+sWvBTxfs7ztAMlMZDLgk1nRS/u+in75eBXD
rno/3oXHxVfVXUi/yPNpdypS798FLFVh7Wb+flMLHwhbacujaBs1s+Cntz0A08h+
oeX8Q83J63+fByiKORcDejxjUwvKdCFx7d05NYNZTQZ9/uJmuGrV/GtUgKTPGAdR
5u88WEsiJunL/fbopyDAOSbl9QB+opeSlbpjg2Xcih0uCuLxhpTwH6Kt4XfAW+/7
45OrHCH5FLVRdiNY4q/9ovVebzglWFVCF41d6psh4xeGVm1VpvyqForJk290yqM0
iQS+GcTeGDO+5o5CdsAgLPO3pM2JFab0a5dHBaI4b3DsdzEBeTHAecpY95l0U1NC
naX5RIwYXclgmnZ8RF/D4+BzxrWV8ZD3d6box02r2l+e5zlGydFuhOAYk6myNEDd
qYmbracbaXceHtrMP1lhCI7ojC9ZWJZ/UydvFQdc+No+2ezDez30/KNN/sn+FbHi
LJI2YRxQwu1phE9NlNCWP9ipq9NBq4Bh7HhkdW8WKKO0t/a/ri4LmUzcfHPaDQJR
amOPtbOA+8pqwMrNLzwRQ+eJDGfjvBa9d2jD8yGKSsVcssAqyoJmDTJqlSzmxNRj
h/9ZAh0r5Xvvi6vnx4aNUisiBo5kI9pRHwR8F5jxzT+lZ5iPI9Z/uQeXpqgtVqmo
IUSquLkQwmNJB8+JPl0gd6Xmkhp87qel2d11v8kSrGRhG9RRalAPr0/m/4fZvM2E
Ak+KsKpdDPFwUO4YehV6eXIHN3Sa32JqejRQtonB+XCtg64vSb9jCWPiJr7H6zOo
CGX1fJk0kGEnH/i0OJZDArWpSh3dMBRUtSLyKgwlJUcuZfeUIu7itKczd2+J9o4i
UlgTp7Nrz9EIMjzAE05kb1gNKVFD+99RkcFav0JBjzdU52ZgZW9Hc1Qdw3wOgDGq
2/yu4tOouD5X94oRSHUBwcPTdBC9kuOl8gbYz/JbU6/nx1IVvvuxJZg/4wP5va67
3ixAld+OGmdqCERmdByF3BrYQbEGV5Sv2BvJCREvc6uqN9VAz7xBdVtziBlC+bop
a0KLd7dTU81gZgjToPwRVHbqK3Iv8IbaX2t7ZisvUtWhZPTHJT2eZ8sqenK8madp
HmXjX87k/I/0X12A7u+GaIHmcv1JvtihyJy9pWmajNR2yv5pLI2S3KvuMtsiYC+3
QIpLLGIGxgfyUzmFkliQjGiYYJihg2rrpc6vRlNv5moxV60DsmOnnIZyx+yQxf3C
eB2TC5LN7zUaSm1qkhIYGfdySJSwmjKtluWOKUW7QkfXroWNr3yUAm3zVuGWD5gv
Q84E5vlF4HlPo9wDIFljyRdoqlBuYS5oRM85J2+dt6Kw2l4p+5pRSQW+gLfWQkSO
OnFwbeD72+kmyonNaRCQsiuZWFXXj3bAJ+A/R1Eqg3TGQjW02NENJ3Zxv3modNaT
Ca7bCL2LzgzpA8GyECB2ifgsxdtE9UgRwPZMprPDoIIz4/3FCEIQ90GQU/aSR+RX
FXi8DCNmhNz4+sSvtyZnSawG2r8LxXGceS2kHxOQBLeU8NAyGVP0VFEIzd8aX/Sc
QM/Qa7qyDfQzVX2IYKoe+TP1LjWMzuEvI9pJ1BFrUsyOhkzBa8rqP2pZ+g3CBKfG
emcTXMpFLB2kaN20DxkM7hqv4jfrOJL6LMsdI2qPxzjX71eVoeVNvuIp0FnOwNDu
/SuABxVJDNiOIuKIJRAZRS7JUhEe0EZvydVHE99Ze5sFvBCuJ5PzTONPb05kRjd8
aZrfJzu2/vwAbHmqG0AX/wKuq1CKMmCplmzLCArMR/2PNWBNj6YCmmiIAQxKafEJ
SA78TGWZHeiYWO5V/cyiLP7nru3+vXRCXZIGX3/VYJnBSkg/GTXF3QczT4MthQh6
Gn582CkFCWp36TQuSy18f/xND7wOGs1OmW8mhJQmPzcnhhle1fU5El+u3Zo2pEUI
fUljnBkmai5pZsPxW9Lb1smDvG5DWSJ+uDwieTFIdWQZQA7LWEztokvqdHlfCJLJ
obmUexdat+kqyI6o0O86lt6kp/LJ+MgsvuSr3gJwiV1g4wlWnpM7bP21Y8ld2Yla
WpDV4CDWZzSD182RQPfd2uFC/yOPPp7VyKUkS7F5ziGfD2QRB92ezN2bQd9IeVZe
lLWjx8SIjffSoyUA+TT4r+WbyVZAinMDRthWTfDTfMlw6Aye9yTzHvUl0ehjtA6/
Nh8ZruuIdt7XhiibntOqqeoXbG0ZtcD55qBmHztPsuZiQohfPZOipWkBuZc3MfZi
609kCUQz0jxN7lm3YhgrijoBR4gE+3wd4C5NMboHoYBSz1IQVA/gDSXwEJQs6SGJ
IAHRgw3f/UOAInNwmG55Q127aWFwXCJVltElma+FHLuFt9Z4i34LS7Oi0MlC3erQ
3Aey40f9cjkTMAHKaV6Rqe21O0OtusDOWF/rHMIXsFaqMcNd6mTn2NYPzq9zDrby
nD9W5u4sbY6GmdOXsR9g7Jrwb3NNCLfhe8dIZY7qAt6XEfXj3eqmKLMmC54zHc+Y
3M/8hbIJD+4BcleIYE+OhSyVFHmAPwjz3aa7+g8idfjyk5rqIjNv0XvUxdsBkJsV
RCjHsc8BO05W9aPDD8C4a4EQSUm9KmjqmSN59E/YUiv0L5QfMfwhlI7Ylua5rcsO
A8sTEyFY+/Abr0H+8OnIfpIIlREMqBmX1yc2FGuPcGwWkzG22l6sbvHHRK+wwQe2
73YZfYe2xhElZ1fhDDQz1Iy1ym8Apb4pvxf4O+5b6Uw1oprZnYQ+pAi1JRcmQlRb
Q1wS4PW6VkW9Uz4zntv6S/52/SHl8ytm1dIDQdQGCQ0qfClKSUflAqqgD2BL1hTD
6j4ozsj809LxJwQQREF0iZCI2or5Tyf+fvT3TxUFBJYWyYqwvr5FDDmY0wtreNoC
jPLvefOcc7+E9JCxG+po4NaPYsJhDnESFU2BKDEGHKUibG5o2ok6Q2AchToX7mZU
0BwPkpWfb0760bm0SH5G+uPUEImXBCTWMV69OOjVb3mK9PbMj4/EB5jo8pttVF64
Jhz/uzASVG33PPo7AwSDFcyv5n1Lnxfj46erbSzC/CcAtNze4pah+f0mMaMGowFK
V/ngOimZSKrx30Y1dmu9cSZ19l+qCHtD+T4ngGuJf/PAhURoAy7dUFsIwQVMSHLS
qvqw+MKMzsGbjniIntehj1MXh/w5FNPSZYTolOP0LVtdlDGU6SAg0v4+5zwWFM5k
vhSCQc8gJ76Bvy3mi4h/kpbVWginK2Bs6Qqpya+V8AFBTGODzN2YIWgtIB6OHkBX
TY5a6e4IY0Gi8JJwzNhlzs5MxysnVXCiH77ITqlJUe6QV1AcCh5aofUGIF91nHYp
tpSyBAnF9UD5znICi+atRzAbcYzk5zeoZFx0JDEpCrutCc9zQHm3DV76zaeDnm+D
QmIg+EIeH2RntcJl90apxoe+kOTKTrMruUsj6ihO+J6qafkFTlehlumcDrMS6aco
A8UK9FtZFDq8ZE9PrDz2QrVB+DOqalOchfa7nYiTDe1c38XNCpN5qrGQz44Yf8Bd
0/UkEi+wr72/nYpF8KCc/Zx4SAclEBXd7CfwIMH7J3xfYc9CXwp6wBTfbkUDcV7N
b+c8CFimArSXS74V+s5R6nAFqX0NolBXbrg9J4ncc0RlT6adKXXvzc1W7LM+/9O+
Ve6Au4KEgBuUzuFLPwYQQkaYKwzPdqbGU7v0qdIIwhFpMLGI1iZxAZDIqXPpxduo
mzqJkUCOHxyUJe4MCskMnFnZ2eOi5TZurSoR3vPGFBwS70fMdzYmNPVh+McBHe8E
IMrhC2FLVKItQ9TJcncmKf4WVhK5imQAgUJpmAxqoS2sYzBDJ66JwG5mD+9io5gc
Sihtyu5oCVGCbSjby6NAfkUoxigSh7tSJ0+QOz2mVSRl/6+wr58zQNLzLe7DWjX9
m4zqWTQwyd4HwQX/lVVM1tsS5BYMcxudFbUOIAZwnp9swN6VunADKjh3TGs38ZtQ
SlXrTYsFVPx4Eo4NJ2DVyx1ikzYv4ktoGa8a2k3vdUgTD5AvG0tqcq6UOmPIB9iF
2RGTuPmEBYGKSlt2ynJDlY2CVA8dpPU6aTcKyprCWd3wKiQOrC87oCdhr2Zo8007
mXBGo2kubGvWE5HCSW0MKBaIZ5SDpvKEqlDLoAOKxwOd9NFKA1VzOg7EEzCJg4Mq
46RBQ/eQIdLDhJru6xcngaif737iwOansxMvND2ggKJFxs0MzqSLZ8foKKw3qs8R
IjQ8WOv8Mw06iD6A2GvSqNaE9jBgojPCtl29EY2QQVyNxgPUNfkWQmPQ/4Zn+lNu
5NcaKSVGzcAwvOC61WeXe1FwfrP8L3eJlBMRIKBX+y0GH7CuYVuBfRYnhr9vQnGj
t5FrKHlrpbH6YJEQpufs2v06s1CXQ3Ck8Y7op51rC7QK0Nr8ijoDLRLPPKbsqrlv
ccw6K5pdM5K4OWNbQTMQG+aeJON36MHgg4jfjJj4Ho+7V0VCRJn99bROuCYJaCKC
W2uFbpcMrkmzr7QGRR1CbSjTuugdvrcOubyM4tc0UhUDgsO6ICcHWEXVW/XM78lb
RRO/KUPhHnznsF4D8tjED+FACYLvnP/wjexx+oTAGvGjdz2JKT1ab6nx4SV6Wo5P
1MoYA5jGV/0WmrUg906hLd78BOmvHuHhiDL0eZK4lgvQc2WAS0FmjOfdH7jeXNV3
Yxu+sA6PiQrUmNBfqFtlpzpBeJ34AiUD09oTI/mBJBE7m+CG8wpvet6KyIkBLqyM
p798WN94aN6zVV/P00S0SX60Zao9N+Vi71yTtcsFtyfgoK3qMGVCXINQ2q+CUsVe
alxOqDlCv7hTnBilmCq2uZ/HMKIUNEWVBp1JHxW2i+0/C+dx0pozxWu6ynRvaiEU
BtOtmrX2Xg+PrwC3gTus9d68fe326pRwOevjnkK4SeRgWWh25Y8IdF5WVq+5xq4Q
vOQby+btzIgldJEqWf+DYpK0zanETdlZMF6byUvawvmYLulFeXq4LLjNMai6fJW/
t1eFiJAnmmyt1BjSlqY2wAwHLnSn2GM5iaATJm9ZqtyfwKg93DBYrclP3SfTeFtc
mavnADElY1tb7Y7TP9yobyY2YP39iq2G1zouTelxVIxnQtRBn3R5E50yjqsUxA/F
dBopONq6KxxKcsDKrehgIQauVMKDfJCMHvLavJ7rLEfvKint5fbob1o3UZ7qnkuM
VTSNTsOhgYKGivBvfFkzex7npGkVKA/thbTZ5nYqQDyh9n0FG6ZdabzikMjv513X
0X4BhrnqLp0k1a1BYEa+4a8Y/KAQdjO8foqEh7R9BGYEGYcRLJwzZJsYXefvkr+k
5fQoq4LzE+ettxwL0VwePArLeShtMMTqbgUflLKRgti2IuoBGbMbyJ/cKeYi8a3V
ANQIUL4emoKA1vX3hoWLpiNN0qjzS9Hz39AzqomSKaBh8aXcN7sGw+2gWCOOrp4D
ZAPS9jRH4i+6pFmM66r11hOLN3J50wpHoYFN7nKl70fcAE2/aoGHF0MP4V0lIv1U
6CyMJYG0Gd8QYrqIq86SoTwAz3H4DWyJHycwbhwQU7BiWgDAPh5T0noh01sk0TnR
FlAANiGEstTked6OBZtAvCy9+8DuQlhCl0+wV9xKQJqscJm6Gty/8mgRb42l09SY
qK0Qzr3QSVZgCifAnQyz/cK2JNXEl5/vTa+E75tcmBf/OM3koZP+dny8rW22KBT8
HINP6/pWCh+eewHDj2envnxdLE2F68ZLYZT6NvW0p8o5Qcdt1T5/027sOOmSkVzq
lZ+Q2VwHRTMa1GDSOBT4yxIRme4u0zQLpFL/rr+tISZGQabR+nsci9TmwDWlKT/V
/g1+1R2asmnMGqoWT2rTAziqONXA8BKozEWekV7Gc513xSPd91r0AOk9ck8La4Mh
KxETXDGuFw2Syqw0ArVih8JAZH8EMoHDN8rlUxadhUFftpTDVC8FYJWteJJo5pEY
SfpHYkdqm9Ff0T++ybgQaC2B+OVdzOnvpwofK7I8teb43X6rO5OqlRpqgpoGmLlS
+g99gwzInrPzGOey/Tce5qoUpfjovqF4JTgScvwD0SeoC5PvKij5q/ZdyLbc9dsM
lvcKldmsB5lsWi6lmvy6/d5384iulx9DlvsMsgEk3yGdxPCP9KD4RUYa2YvVTMBo
r0vH4inoCzWbHjhCAwhdDcnKEYNUKEbAxOTOhgHRoeUlGUKwLoyFmBVT8+vmWSm3
6W8+sFSBSFVpo5H4CPMJvFpfFlFBli9L4Rsdd3+3F7f4bqgf1U9dQwGD9Gi9SXVh
BIbGOmdmmg3V5vzAXnzq/9NA8Ddlkgrohjva0KTfm9TYE8za+3JpUu3cpv8/1gyw
p8e0vI3NqsIKjGwz3WYGSPhofKlZkZhw5CcBUSlDmBbfGzjkUOEdvCq9d/sa7Bnz
OwUJAyvTp9PdwGKZW575/SFhByxMh2cyvtTPhkFnBrmMyBw1659PGcS3GBMXXyOj
2ZNH/UYtZLRYAV3KzukUiDyWqbsAOt7tEG/lB6zRDODn6rzo4hlxerxZvB72uZnq
54Gkiem3v1YEEZ1qqiq1Wvv6LvXHbz4wJypu8Qxo6/j0lw6to9GvrQJvjlWLB3jE
WDzFcfxn+F5Y/nYuk1FfF6pml6WZDUZhRoTtw1uQ4u5JU/r8vDG3vsSRXCoY+qcK
n38EzCjAv6ZYw+slBf7FKMIbmwy1+9sMm0UlWUCIJRSKWIgAwxb8II3VlsYS3fNy
8o8uT5aHeXaqKPRII2bMJuXc7x0qVyxGtBN+tVnNK8XvuUmhexB7sRwQdpEMTKzg
W6mqFoOUB4UwsCGtNUOZOAd4lqhxR1XR+XqgaebfnzuxslDG3b0OCjcBUNK37B0p
G2S32IN/pj5arhhU1skV8i5uvGLcpNJFhtZqOgOcDlBBrSyDuZ5Fb8vxETl95haY
qdNnB63nd7x8ucEBxhI6wxTsSG7/r+X7aVJz+aRIovdl8m2aUBzqCIY2y1jHa1MV
mk55Y1kp8uq/t6V0B9gejkwDH43XgqVYYmymfXRxH9Vvr/yTlsx9HoHMMFKL5Jor
bMkd5EwI6xQUIzR7kGKcfeHCldP4XvlOuoQeByb6iPvro3o77nI7vdV4J+qOFLTv
thaP8lXzv4fwOBkfpphf7WQKSLzhGrkbAdx5kYYUqISdB2PweiiGSV53Z8wdlEGH
3MeCZnoGEBDuiZ52IyqOQhZ6MOeerOkU67bk/kthrIBkSoNktqyqqDqhgrgL16Ev
2Pp6bonohmAtLZo9dIFfyfmrc5qVyGg2BtKruhCo2ycFbCVdTbUZfuHn3W587x9+
3v/ZR1Y0Cl388hp+zYs+C8PXW4vHLadXC8Kcg2sK/A4bOMET57LyYXG7R5t2hF7X
9cLiDQAlbwwDYNFO+R1A1xMiGX/PLO97QjDMpDR3ycfVWsV/MQRS4qIsiFpCScqA
9vBURf7PRcvhLj2qlvliJHNIn6d1zyrkqmHrBqJ/YOGcfegexFHwKYH3AyFp9Rie
STAJ8wABwWbSlMYk+WmdN0A3do3IeVK7O4sZzUDWGZW+7aQlL51qWPE2JpX20S/8
FM2i2CMEfS6jUEqDsIm6t1IZ0l3FNHpvw0g0pwR5RuOhl/8t3fUJKn4mKBcYZOPH
6xvevR4JoUdIRj8bCqNHpmjZjdgxnGNTKPcfAwroJ2eg0lMoETj+wPSbrRhGJ1Sj
dQzciIhi0+FrcTDVg3buupQaJRrRK2tisbFqb7zgpZ/8BzMWxFe6JFshhNSY93hZ
88HoVgzgQA1lUYIXNtw1N13WxPm2+uOIyW6HhgxFVrz26C4FBaL4/X20/PFAVT+s
3ZAAE3+qdDp+N6gSOVfoG1w7XWFsEPAHdNC8nq0tblg0VENPu0CYTTxp3P5+Z4Fe
1MkXuFADmM4dOeOWKY1H+CdBMtoJA7dSE0HEfz3z1d3eax88aEfIW9HYKJq5DIEM
tXUhkSv82hWxpcGWvctmbpzEoKqP3JZNdablUeK+AI9JCjPA5cy+bsAcs+jFqwiS
V8R5D+pD6fk05RWDE/U+ANPONBl0nG1v3BtFia7FaM75lhd/Q0WafNbHDlStG22H
I2YIfwIU+WVE7ExlojqTcKL1fdL4PI89Xm8F4Jy3Kwdkyc9diiMMJWcange+RgG1
yiSNueO7wpIX4DCVU0WQVyj0tkhcVmDUF4zkUKqW1jComxO2xy5xiPB4XCwybfEN
cysKvhigypPFoTCJ1XSvgd60Eg4C77zur7bV3yuAvgA+05MQH0m0SBBLKpdIUQat
dcZLiiGXogy2oyqF1bUIAxHR41oy96ef99A194qBX93udrfj7RLqY388Jc8Nw6YH
4H7QFCo+tqcLitxguBF7UxqeO2SswPbnlPioR/8H15J0pwaubN5OGlMRkqDHyZIm
znzfI3/N5uWE5Fd2I9UO27YI3658Jpx8OrwF76rK5GHkGmtfCv7cDRPmsyx7Xf7N
Q5HlW03xyGyWbRXlZSvy8mrnrHqzosAs/3hi1XUmts0hXowA3iFq/VFtN+kJI0cM
c22RIdNpT7PfVSG1NRlcfvN0nU1pht9IQ6ZtI/RvB8GMBpzE7mlmMBHpyJcJsVGS
1o5g0onEBSs/5D2gfpUc/8wVp5G6PXG0pwU9AIUT3E5gmpUxY1Z4ErUh7LljkjwK
MDoyYB5jF9Pc4uDN00ZoDub4Pe6i7rExrBtaYawYorbhXjNHrRNTrJpqMXFkmNIc
Tt/4sUP5/SQrE0SHSnnE9nOqUVmsXTAa1nMOqklZq1fCG2y8lvuq+82VF9YIjhSx
4uKzyu/LdZMyvAUwYoSJdfFLxo2/17oVSivK4o31LP8SRG6YC0MHctn8xIsAZy62
VD1jrqOmu59laUR2rEsHFQlTq+pd+6/BgnBxP/wC5I3biN4OB/Vn4kE++4a7/FCv
1fw2SgnxCfR0iU0dioMavU30sgs6Mfk07dGdlbQlrIa41BWHOObP/zebGmRuDJM2
P6BrgDZF6aBv0OWPTvrA1qLeWtGCkrOTFAYnQWK+5Zhw87ZeTC4tTubQ4IxR1lKw
jf1TvZK6g9IWdv+bNORM7cN1dIPUjzZYS84nSAqH6ZNoGOW2R8NioO1RpqDlyg1q
uVljW86RkB2KE7wSwOKnkOYN9NJgKeeq+D0yTUDbmudOV/tNJr+cT7HKJKaKeNEU
2A41DzIwJpCq7feznQGJGLdEvg78mpsVMdsZsLiHOO1A/zD9/NB1Q/Jlgzva2vKQ
2s35aTDG0mbHx8FgOB1PmFlgST5dzZlzkHaRdRgXsLqFvvzAahx3We+xog5zNg8s
DNcYJzZWT3CJsGNbn95eiDTy94ctVbpEC84enk97T+dBIekyKIk8afF5qiFjgGa9
v62b3GTgadgwEDAUyVj2nt8g4pvU5FD6Joclop00Emm83LNcjP0UoinQLvgU/nft
5fyC9ZJbS+eTwfnU9LBg7Jq73EZudqOVngDRxscfSofrKXqDoMRWaIqXBJwSepyC
zioztB0PFedX7NsUh42t04GYjGV2rtDNR68Oodov0Aj533+2KqNFeH67MXDnssu9
HWu7HXkhP+t3BFwXfGj/fA==
`protect END_PROTECTED
