`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VciPJzGDi/zm1ZPhD2VB/aMaBCyYnAuWFF3b0PXq+hQdy3gZBpGeO8N1+JM41Lbm
w1UladP6/njpQrhe2JjVoFTSqbDZPney2bz5FxeaWzV4kXqEYyfypD2qF8iTcfX2
9mZbgE/DCzf0MQLh3DCyoQWI5VlHOhiVGkohDpMBbBe1yYnqpgtJeSFgBPFWVFGp
+JkvME2iH5G8k0HxjcjjGRD3z6ctHIOoej/uYOETbzqvwIaTm3NMwThg72OWFipp
eGnVCFsnfaXQLFwQJwtF+LqYG10pjsWeNnAIfQyXTBzwCia8zFVrxg8nqp32IyEK
SEs8bFjawvZJ/fyS6ObKi6nMpHb5ZmrnqYYsZH+nC8/JwdtJ9U4bPvY9dbUhTW3i
L/YkqCcrF7W4PBojpdqwSckORPbgHCP+qDcHHEbvZWxGTrYL25g97do2ojvZidAB
`protect END_PROTECTED
