`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vhcR4N0WWgOT7cwcXoycuUdY9CNXeuR5Oqt7tHKxzmEeeLdtPjocyN2EsZm86/SX
fpj125eHGBviJVrasYz8h43LiYPdq7baxKGkqo3fmhb1gndLvpmzWMrXBuzc4Q/b
cba+fRUI/Qqh7F1a7Cb8rjUojfY05bdPnC6uo1sxjPa8c/okSa0f8ifXswKRXg9y
id6VR+3M9tiHs8i/3caoLzWwn7nt/8klCboK3Y5Czx5pHzdadvlOQ27e6AZ1+Aw5
oPi1yOjQ68++u2rMiSKv5xLHs9bxOLWAQzJSDkMyyHD1QEmcHt2fzksRYHilueVP
zK5/XHbbGcjQRBgWWim5bsepMyirv0tyXravSWS7sfdgNjgtL2oL9R6qGEQvbxUQ
Erjiaz515L22aT6FtsvKtXzrDo8PCPpMaVe85kbNfys+Ortqkc8ai/hXK7BJIAYP
`protect END_PROTECTED
