`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BJDYmGLLWN5+WD9/D3OTqehhxrupH12ZELQzTKVVzK9OxrvHmhw/9S544UC8vVHi
PZxa7MHB7Zn1cLHrpYjwOUL+O+kvFv13aNZCFWjLbZ3aUjnNGQK0LJ9XSU2Xedy+
lw4HY1k3rGyJK9UJizMoru6dab3rhL5kxuT504DfScoZ83o2DETbatm5VcVqRutO
Fsdr37sl1rAA2HT3x26uUcxoa+DVsOUkb6wcIiQMIGbKBKkgeKzeppNSytuE7jF7
ZIdpCS1DreCmcVLBn4+qglCW+xMbBLSvTGok1RaDOZ42wrkJwKQmJCur45P3V0LX
NWJezMZJWKckDcwoaRM5OfuzfF6hA993EplAebPGPp77H5leIkCNDcfywCyeZWEY
LVsawCpJSUEgrkV9T0i3vpQQ7986jL6/vLYcrLVdmImKXWCMDRVAIlGjfITiyhZP
pBsUP/dwQ2xRLdzLoqiEFk2ni9pyhpEn4BW2Yz4IsuHmeEv97rnPZunL8vXGShQ8
1ihTlhTl18IebaRL1GIGGRPVTqlEpvKKSML7WN92FhBboV1sjkb0mN1WyRRoN7DD
IuNdqmnIZ7P4a56eaW6tdWARdZ/winB3lTXM2mKCxnHIT3/n4fQWKZ9PeCgv585y
YZeXsNoftB7EXNAPTjk4h7JopsYhPFpV3hXcJxfw8Wsfi2+vpxkXcszXTA/6nwAq
tPD4StMf4uY9+IEIPGHFvxFKh2xTt3ICKsX83er3CGUlvgamKlpWouO+NLQb6dE6
wAC5/Nt3vV/yYO9ng4rGENYApZHKrX2JWLm2kimgWTY8uDDMgoeBn2akuPKZUT8u
J8O3P8mVFbHYFAjUCY7unT/ElK/GuEOtVa9ABawj/7UlZH5d/Au4KL2Wt9JGqHej
MFctDWF528HdC5MgxqAdjQ==
`protect END_PROTECTED
