`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2fCpulgaQrlsKJxqHDpvty5Ofp6kJcOfdJi26VeyeDT1PZgsK31LA4tjctcly9E7
o0W+JdIL5FUeLf4h7BcpHo/eOquvr4xs8i+/uKzWDkQZGHqOUS3NV1KecLntnbhd
P9mDE9CkDK+p4/SABarYdZqdblET6ySmFWX689QeSNCGXQwkI8zzsz3G+1Elqp+r
ggU/bKH/7WQ6apnlFDqBFi4WSRdSw7nanNrmlHnpwa9qgvgr9sRwQ+a1Y4SSZS2W
EOfF1AdZO0R57f7ziwIA4A==
`protect END_PROTECTED
