`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M0ZLPns+75feGINaAdT2aOwer6RXxYCdy5Fy41OsH1D0n0YwIoiA/ni3QY6Y/whr
d/QP1eT6/b/sZC9zt7xmXqrUFxvVmSq0tG36SnXD0YBgVHsRSLiGpGRiDuceemZr
HlpqK5n5MqAMBfeWrDOUlTNnvl8qgSP29RalMd265ntureG9Y0L4VHOi2J5yKYPS
QF5dhFNTrsI6NJsC7S3mdlVYGcA0dNvAtdiVwrGef4MZzi6SQKXu3gEV+4RsHVLK
IDyU0nKb8cmAPzpBCfLgp3Qt7HK2UPLirLPQBHxbJCtvfGd5Uw1Z9ZFjoH+pBCwe
G0/97ay9C5bb6WamHPNsf1uMgYYWLiXAGIv2EHR1oH6rRHGJStw59JIAoMExbnrS
ew1A7LNrTIYdG6dD88ud0RjX/3b0wqWBr8AV5b6tAeRKhGlXa9meijTkvx2eiBCF
imbCUwjBehx3XQ7JND6kpzc/Diz3CUdGs9B6nyBQoq8WJXVXe1Pwfhw+JN01FQ12
`protect END_PROTECTED
