`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k5eOn/sRLfKrN7EcM5RdNDwX731M0xXh+5oPkVu5EXZ3B6e5EopjiK2qWqgb8YgG
iTYhL4iD1/ihDMMFRZj4WPEfCRTQRToXt4pS1fcw7I4n48PbrDfshwX3sMVIncaN
z+XvEznr5Qcj6NNOXb6JbmPHHuwpT8913V5jRd/4VCUB5VgGIRQEOrPZ4SluoqV7
uO0MSjQ4Tby29VerSmhC+QWarsp3dZoNwhIUapc0HwUSDTXJfHmrb74oynbdiJp3
ZmTnwkqdkjqcX7rhvYUyOfyMZJuwLGSmgJLwGxbxxmWtu4qOHRMCXwyQ6qSaMKBi
WmP1zNNE3WbH9xX+LR6ZxNWUzvzFOmalpGDQUY80+tedMf1UWurBbqm9/lPOA+XV
FyJTs9+IFCB7XHt3/yu+fi/ad3hzQUlIJ9TFAaFVOdVlwOi5cFn1g76aILl7CB2D
E/vvZzYEaB0qee+OvUVAlRZJkWzFhw6S1gahMdVOCLxFRNnUW+pMGCP6tnMzCBcY
`protect END_PROTECTED
