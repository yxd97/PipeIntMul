`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q3BI5+oiNy+jEdkseYaYkWHpJnXbD+oaFHDHw5wySXpGXUH+w19GfVvwsPJRgydX
giZ4E/e+2B8ZrMhd5nQd5umU6hV9eaJ7odRjT7btEH+jqnHP/WPbksrRhd/q092C
nr0oqlecel1GRTUsIrwGy0UZxJGKZj0MesWw16pDC7VlJMBpDFvWySAx+6GVkolF
xEVHrxJXhuRGNJY4Kd3DFSBfOaheSdI5fSlUEFjPDD+/a1KyznMf1gRZdSHmLDRm
cttGGVyMuWaFgmHI30atUlBJvVm4luQsE/tabayRgdOh2DcDHL05Vzccrqu58bL/
k8wL3y0Ze6ojQjGWQZmhNw4yDV1TSRxVSpQgb1vZaN0+hSCJkT0tBj1vBpkgT0Hj
WPb7DqoSe4CytXi+oTNI7qrapriXelS7tJMyGuVsUkbCIlARQbySrCA2stI7z5TZ
A7Hj7egm/4h3CQzlJMRXVU81PrLHmDaGrqn5UPGOr3SeeUon6P3Zu12BEfPAHame
eSxysVT1pPk6Yh/5HKQxjHkPtF3dxH34egn4d6q0tPrdxHK1wFu+h/PneFYtTr/s
WBy57+9DnWgBoZEG/Fc5c7lb8yXD6G7Nax/366wIItwaINIUlrT+uAImLmL/V0kb
6obpK7CdR/y2MrfR7YB8j1fQRwChd5RR21op7yzc8VtsM6pv1IllZvqBPXNPDGDB
uqKWw0Fw35Qes4pd9/3IbW2DIBa7ZFfnkFp1MjhZbFeVuZpN7UHIFmEYDEn+vDFc
YLdQfu878QUdT0aJ++OMBKPu4PWv9br+3IVkNKz9ekS+gKD8M0nSmQGjzs7pvSXm
5S1IzcuxiQ4mp+JNkMSY3Pg4MM/pEW4eJW0hdW9fx1y3nJXlfje0VfTmucmGozx7
KPy901yVxQWAXCe768W6XHP+umvz+yNuftSsvt5KuelC40n109EdoEHTZX6gPLe5
OqWdSLKHMiL3Isrf8O/Rm3m7PGhqgWCMQjD04b8HWKJBBJXojANjOVDdiDovstcJ
rLmrcEn1RxJOeF5GLOih/fNFi9c2M92YJUvKeALO+bnO+G6K2IhCHKgVx/dW0MuY
ajVeX9F5hJbQu5EUCAU/CPl2P8eoET4egpnG35BrVtSwwtXLJcfZp193w0wCzAea
uqoXzut4YyySGBMN7GASFNrehdDoBcLjRdTQSA1KUZ0TgVI9tzFmtSwTpsL3OvXC
RTM9ALrdjZuUIvZvvEvH6Q==
`protect END_PROTECTED
