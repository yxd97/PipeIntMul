`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FgzSc6cnzhoP4fZta/MVjyTiwQRQfXoUFV2dDqXCGE7Rytuh6uczMkaNRzG1c4vu
l9+cBdqoMi650FvJ3q91+pgNznWO/a0uszUOmQXCCNXt3xUtSm8GqKTbNfjiU/fO
KSbRcsCjAuRJ5ckqPFBJW8nd4g24SwxDPC1jClZJ1JjkxFzYxNrIRmx/U3b5vDez
aBzMIlXlccsRj8jIZRKP0q5ICSVFhhX37cYggmATNSxVGQ0m1kgcMo0/qbQpyDMN
KLK6NQmfWsTa9WfAqAQAOdzKCZnlJIztZ/C0EXKcte/BVWR09XLkfLoscmFq8p/X
BNz37IY7t9/po7AJYR/wMZWBoWBtcRZCwL5+fJPiw4THjgAt1WeodZmqMV0nrg3X
weGTvzDnZoAG4m/3NyDAzecEdQaKZipi7eWpYqLMUgw=
`protect END_PROTECTED
