`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufVAi1PxAmfetR/q0/r2enZ/tKkPZPKtp9EWq0xBLHOCgh02XK26sKUEzfVnL9OW
TXhIJyo2+yUQm6s7ABYyCkqZJMTb+fAwi/erj4/uQqfn+2qWAhV+Tqhv7BGkkaZm
loVWxXXJuVeXasmv40m6L0gLrrrA2IBt2bEZdUWCGSDTrEG6sNXKLjOsa01DQf5C
nH3O0KcwvLw937jc3SFWwLirgh0lhJqRLdCKrsR6hPA8zcSD6VqZECOubAMSXy64
lJ/D+umf2+Kwt641vfsySSRyb8Un+1U5b3eYIyLi53r1u46wKV02WE8LuCLD6P28
SpIbnBWibXnA4ATfB4d4KyoD2uDRpdiztf/bALCxweFE68HDsW+uLglMhzgI9J7N
5JYvhcblHyRQ+1WK0LjAMx7nvvDhXhKmkoAA2SXLwDYmx9VktZKyFVAyqMyQoM0G
8s0zNv+iSzJ46o7xundoF2gMYrAVq6z+U+PZB+kZ69YkscdeKQHcoKRqwU0/R3UL
ugKLqEC6jBpGV6vesLnzBJZiGJ3qMSHYO+PeK+XW+vvRT9pmw8asnKJQwad7XZsJ
CVcvRSZeuwCHAqWqcUGFIaUHiGwwwnFYT42V5FkfgaJIPiLJEn8LVXOjTjS8UzAL
Q9b62xLyv85ofPskM0cpvzADDf4gVFWgo6auUWpi13T1/d58z9vBnEhaJaQ0JNW+
8ATnIsYJvvO4TkP+5T7ljNZ3ZPvQPStnvqaZVpbVhndB9901MigpVlKPKpLFhsY0
Uh2pvU6i+eHsbjTks05NTNWWQZH8Frr+7qdvmnx1/kwstvorLZuYNFMOkqc7hOgH
GmrZjsA6LbTn8f0HK1ecdbC9/U/OkDk0+QlWghBZnbrJVUpAIl7gAgsi8z7cDhhU
cpnUn/Zgxezxx0aSPeINyHKC8rCLWYD7O486lbkwS2KX52U7K1tlfe7O9+hZa227
ruaaj7ZjxMMAwCzcn1rzHPkYoYh/FvOibP1iuCv5UKAbGomZlIIo6tlSXVZgLvrb
Kk42GMhWvCb/uo2BNyWgQJkohQipnS7Ir1DCo1we3vfPR6WGfl66AMfduWlXquIh
D9UFktoqIHInBqihuIhAzo2/9dT+Q3qI2piZt1wuFcYAqBvEaNRCClnq2I0nrfpD
QT+npv+AdvLGVAoguoReJJwS06H9xtMCztbyZ59K8nZ1EcgxXV4FDdQUWL/+NEv3
7wpNqdgHzEM/DqifDnNtuul/D3TRxAY6l5BMr7WdvWIpV2d2YZp71rJ5T9L3UiPE
DoVV2vTscE4pe1Pt1S1yV+OqgDXnwNQQadbyXelM+ISRU/7F3gEA3sbAYgu0EhbG
LZS9Xw6c6001xjGrkK/7y3u26uJ1prqh9de63Ycl0+f57pMxFTgZzYJPXcCs/x7n
VQEcBipsVSffTiSKpIj7XU71e2zJxsF//2ig9Ai37ntJe5VhS+bxnLa36BMUKcbR
nUJ3yM2qsBJEWrZka/ckYCAzT7lRg+mdOeppT5/UXmwD6djjSypp8Js7ZdgeM2xL
C6gZZ2pJQPZoN+TLhF+CEDoV3gSJ89MXTpV3M2sSeoi2Oagtfsou0o9dtaKn9xkM
+PoztI/KKrJb26BQr8OwKPFlBFbEqWYg5nWUnEtR5He3ShmCUw6M6eTOCm8DwKDF
kHI2P8l+oRf8yGYvlsZ7r9WVSMEEiREBs2MnVPJlBzacXTKOOXraLT1qJFsmNtjs
qbWRoh8ne3pVYjmuY8qONyY/lVH07DRTBne6QAQOiZ6w76bwCfAxVIc/z5TaxI/Z
9cNhZBMjxjbI2v0z9PdpYiEvpC8IOXN7IsZL/0/4kvp0flxaHi3ysFJMwiZxxtmU
uzikf3LOrCZp5VxaPV7kjZPAPqyk0dybPkDF6n1XOnp/zMeT0wxxrnOFrClQ1Cdm
FlS60uaQK9WuIw19WFjIxDUhm7oMcfBYrtBEa7NIqnlvY9uA/Ymb2ZJ9PV1wkqK9
sgCQIvWsGqdg7l/Tx6EIIpoYhlJfcKKue3uzU2yGDW/YG8nmBIh9i5K2vRArPyz1
WSVtsfrpyz53dIRQ/sq/uURWO7cdv5z2TQbTelARJxNxJN2r98GRJhKFSryF6rBC
cicgyeWXFLvMFh5UqqBlSkf/4G8GK1T538o90Wg2eo1zg7ZYjfIecUuPN+OWz/gt
dldn2bmhkRNCFBIwc0OQOGdwS8BrOQND1DCGcCOwzRethAtSrKQOYj1djBOOEz1f
53VoFBGbV9ERfkQZARVcO14wVCknBSWifpVRwf3HBbufzvV3/diC10LgdMJB/bFw
aAgzWH9JxLhmGqiYsRFoKoXTmtoPe5y4cy8X1JZ2uf66m4gl/wbeBMU2DV4psk/Y
HpTx1KJuEOhCls4No/kqihiD4daE8dJqV4/eIHOpborIwdSIv1nW2X/dgjcRLYBI
afOgpYjNoD6R7FD1Hp2s5glFuSaSWV8VDapWjubyRWU=
`protect END_PROTECTED
