`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O9CQXj+753EoQ1nYKoioNjG9hVtz+dFCMqLBgsdVy2rJ7F6L4uuo7vVo9ehBr3zC
3rzkwUCmACpDgOFNBt8mxsMcIC5Lrej5/m6Kjrzyj5K3NeuSF/wkkQTJObQ1jvUJ
q201yhSu12fPT9QISdr09t66p0vUNORYtbF78ndpqpBEPmyDX0mrF9VPIGeTfsJs
S1nWZSbs0xIUEjx+8xSxxC4f+txnQaiGz+StVOb9xHDh7BqQx5SFxbfoJGyXAlxP
nzCz2RK8TqBDL8Hvk1vtCQ2/jSxdcUZb9ErMusbh6sotE5BTNjjMLX+OT8qf6q8/
5m39n1AvZxkADj+mQaNbRHMcQ9v3WlR0FSrwzRkAdxGvrH/aum2iRr81WKJWZ0PT
w+chDE9geBxGIR8FZXXs5bhhSAfDGS8mjQeCawEVUOvwB3ZdmzuKrUFjNVUCNQ9f
Bt0YNErnVZxy1kQwBL7Wmj8nAAkFz5f0r7gAGhsigWpuoDTBSgkyRajdXrRx66nP
`protect END_PROTECTED
