`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8AJG3NY5uY/guYQcK+AjU1jDJt3hWKSjgGrq+LIOx1B+N7lEVvnlIh1ixcaCMIi2
XCIeKhCs/T9yBXheicgeXQybZBg1oAKTAFcfr8Pcbg2qg+6i7Qa1QLZmmNOVeBHZ
TJ+DRC6fADv+8qBMRyDizuchBsfvoCSh7kci5FJlXjwS/V1ErC6LvYXPFjMX44sq
0h4iSpYbaROYqXDUH4VYA75iTkMPWuaniJ5PZqMt8aQxzyLlZmTlv4//HyT/5gnZ
Cjqi1CQ1RE4SYO0qCfSvAnpFZeEpYfSFLlW2+U0u62g61blbEh0zv4BddMvN0AxV
BhKlcSj0nuO+/l0btCu/r85x/cr2M+YJMYqDXqv+xEn6UmpbZhEPJ7xvbe4RuXr3
mtBdB5gFDJTR1NScawassAKRb6XdLrt/9f9hcTcaJq2LdLZE5AcBVDeiX47NPFBW
vSP/uktak4WqSIEz2ydtKkP+/qHP8FNhkgSQEthmQYnYz6l6ocA4bycw45IDr3fy
JApHqswKOfdO6WYcArEw9r+YfJk/zPanKlnS6bVlzxANrf15yKwZKGqAXOyM1uGj
kQhMPAgDzdHuqvnEdrXha7NGVosFm6YqHlw2dhdWqFNlRPtO/JD2t3HH22EV+MyF
k2RDgvO5Ot/PggFf7ec8/tgepAy9PGCuBo5U0qEg1l57rbCCRxWJs2rC14S4PR29
XJJC9pVyTIZv4I1nuWvYRioNa8CIVxkPkGaql4Ry4rS8UG/ff2FbQyTRQQTudb8z
RiDrWsjfY/s5w1KSPesPSVQI5mVcwz+/Zlxx2q0tJ7Q3puEjW82xPtMLnxkHONSB
ex2E1Z5/ZVvCYPyCJxe802EJwqzvQWGf9/Np4rKTgGOe4LAGryKcIBs/kxu1YCCR
mDcnqs3W/g7sZcpzSkNVbEkVoiVAoC5nfjfPVwSjzt5aJ0vGxvkq8aaIbCYPeqgY
r85SEVb/1SkG5t/U1AaUISJ5JUpWtUg1QXKhC4z73/609AurserE6G5FbCmBrufw
IoqPgMpcYIgokVrngyOVOATZ2uFv/vGC/BrpRdOdcWQJ3MGDQsx3gst1/2qqxD6v
lAg1GR9qZ8Gm5hfjCdYaVw==
`protect END_PROTECTED
