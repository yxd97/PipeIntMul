`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2GSAXyNKAtZmQd+653FUDoUIjZyUkz2BOAc5cMybmn4JSuOtT0R9kTghniiTZyf
jQe7ra0yl37HqbUXJ8eJwLsQtgkPuHNHi2sHx2XA/2EyYelASW+JB02y+8EeC55E
CHeYRJdzOg2lVJaxhIWAUDf9fbDHLlBAqbmn1GBOa2gaFyUt2WiS2xxm4RyPhdgj
LtV3RZejbD55TXX+3KdCwF49f35OgYmM6K0Xh9jsfej7/AnXirwjHl9SdrSCi+AR
e9prd5PL32PYt5UlUhr6L2O3THTsZJTBOD1QTlD2496Bq//+HTs3jogNLQqF6xQQ
3SjaFPJ7/PKQTom2/L3zdVbW3+Olp1oPyT1MOYbRpaoxo652ADWf4NNZLQ9oQTsp
+DY/Um5lWgcE3ktcDwHYmNvm5zIxGU2oq6fHb3t0Lt9VPaHApT0HGlECPp7AIbmb
ZsR17qwVdAYzgliJz6siOcv9+sWuBD2gblBvkfswJzqfJHuCHg4uhyV69/Ss3Y0T
hemZ1vLfFMayhUU/Gmrbl6klnVg4dGQOpafGUusHiFl/PR/Yd3ymLK4u7AKdkHuy
qPFlBhGnWlKR470xapigf4sWSL6uTz1NKIdFXzESjzPQg/lDXDybPEZXUGygJDVL
HgAcY7+n6S5EncW6rvGEkG1uzd72Wy29edTAwwvOtQikGsEI7M/VvQUrKzf1mimV
1LZWb3D/W05nYbRUt1uoBbDbIzNhbe36r+wqnCUk6o9NEo9a2ZciNqLm4nqykl96
difDZo3/HT/lklF6/2aqNpUuRunqItsTYxcvGWxBzHJMgZyxgkYf9esAbb4GxIiS
qwH6sufY80ZT+yZCDkyJ8b5MMlAOvXq+CJDGNoCpkZdpFrG9XpYBzfz1z6ftwaL+
T1Q6BtgHIlG6wRj8WipN5sOuqATM8YH5vylX+5e/MF0dTEO3wsBfGWioGekF/Lzp
SBcCZWemRFW6wHK/3OzPf0gpIAS/V8AQjkBmJoMjQibXZ/IVUZgr1XS8h2T1X0Z3
`protect END_PROTECTED
