`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0lxSZYtF+TiewGiUUmbV6ftZ0KFiS1jO+VvNPRitQRAw1Q8iN0uwC5pUK+TapgXZ
EA7S53HEwjIieaLMzcBErkErstkfPfLL+XDTZkHSYlajXtR/uv6drasnGud3phy4
PRBiFW24JHnhE/OEHz/RCszRUezY8nq2peaefskEpFpFPySYC9MmTPVlQm7O4nJZ
wqHJWFbz6xR18QzBnbN11CUYHLpKYaAKH/nGuBpSql2xA99G5C6T9K/Z6WPvH21q
qh97bYA7OsylRGWLJ3YCZYtdPBTbtkbNgm4ldTuILDSD/licSjIRPlDGOiXfxJiM
bk+JzGi6yUG3QmbFZwNtSoSFCOaZu2xTKNMnRuW2+PexOjRHj0Lv+OLuk6vEmupJ
`protect END_PROTECTED
