`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fQaoziDxOwtHPQx0zktWeZgXc1qaViIHKQhavrS3lxVU++vrPYyb+qTGrSJPh/B/
4s7FiBQJ80Y5M/4oHlqDYnAzCjNpJvkKLHl9v5kYPFyCzRVUwhH8f28Vo0s8ji+d
IquFHiWXj1SepHhj2xRw47h1TPh2c18nacpUt8me7oaLicNLrvH0dPAukOTouPmm
j+tBzueSDNhhLvySLZmPIECmRH5QO8OEa2+HelcSiHhUf5TVuxKzv5TveqnlmdGO
MckyD87b86OtgNRuJS7KGJUdYJHnFwzlp4EtQQCDS7Rdj2cREU4BPNUWqko3hSoH
zaZ7jqnimbZr8qd8B+8BvR0Vvl4tFUJTdZhCdRSvwQJcKA3RmNt7t+xX3x9dSTGH
xACr8R7RWXgCLViAUakK3ZSQb/xOoPyGKmAjRVVhYuc=
`protect END_PROTECTED
