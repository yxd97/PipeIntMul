`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+yldr5vzCWPzvgYsigrIDhap8/XBz+vTdJtev0vh/+Q2HqUWNFof/eW6uILNMp2K
RXKk9qxfyqvoLooYOgUUk4JRtEK0YjbfU827r8EUYzxTtgEv9whW2EBuemvuuDYZ
nVd+C8IoanHL5h350X410bQQDXbK6FWxVfrDla2lQroZMmwgazSvi1x2K/jBrVuH
aM2SZU4sOPFcVEm8dZP9fzYwjq45xQnAVfdLDOkxS+Lrrga3lwc6ba2pomDUM2dt
EaMqOHGFIt73l/lNw0c4Hytasr86j3bpTv/xpMP238iFFo4/qrz3cNa8//GMRwEm
NIA00/Dnb3W+5bOWIx0os4kpWuFj5/M5E0WkBrBFPSNhQVhl557Y3D11a1Dw6Hdu
LFxDRd26VQ0O03a3ji1V1k1a/rF3Rx7kZ3v7T3hM93EMZP3p9Gwo7VdsN7QurI+n
`protect END_PROTECTED
