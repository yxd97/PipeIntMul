`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WFslvtqy37swm297EcPHA8Yx+SlI78+r0WS3bExxP1dfMDwJw3cHnOYkinecauLq
hR9yPbVI0Ygl1efFXnywtmuzccaG4kZ6vlOtGb5UP0GYhuYMsBik7bal8Wm1bx1f
qZhBp6Nne7KNArFQu7jNDHuqoJuZwgDDACh/UcYHbDdFA1mZj9qZwpPmDQKqfUOQ
tmPK6jerc1ydFMGfFr2+1efrvIz4MHYkPbnQGRMEzIAfoGO/Fu6vEn2S54+3/TEs
AoGhKw52ovKB0yU9qokZIcecrwrX7Ug5IzZ9/MPmJMi3yUaAiXgVpiC6I0RYscmy
W4ZgJAxE1AIxtkm28oaGsbB6UxMHrnBOhDXnPLsUZUW6565SbX0eaMhKb30/bo9n
8VIMHjnjQAqK+ewsHx+7JGNqNs96jTXBexlVxW2qTYC+YNc1X6FE+40VcDYOlY6N
`protect END_PROTECTED
