`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vmR5r1MRatqqBdWn/40f2iiIYJ17HsSkOlltQzJIBKVPHK3+mx3DhIPH8210idWa
ywkcNnDmX3pC9/rksHrYCZQiNYEzAcP4jdxPrswViO08nWWxhPGIF+FWZCqKf+uz
twLutrs2Vitq3/XPtlIb9BMGplhUFrPO6nsMGJ2a0aKN1MbqxwEU2CwlpDIZVXfM
d6WQpTKL2L6YKfAibrhFx3rO1qKgZL+aPzXekEqJAuvUndYe2si4Gj2x3AX/MB38
AG02MJWjV2+r7puPtGlLnRWgph9d9yNSmK5aEjEttHTTGIdzK98NvvwS5NHGB6b4
phnOtCdcBvRvua3rEq3uVqhTzWV+AEx2Y+oyh7UwkRfDCheU76Zn3C1JzIh7c9TX
GT1LgeGKxG9qE9QNqjHHyoPGMuFzCwvgUxASBaTzfYYfOdelr9QP1vQr+D6rp6yp
fXGXVrB1bu1/svS77I3mavZvjPn3VtWsnZMKnrV1xwozVfolUPrCj+yesnHsgsEJ
Zp8QaOJuAwrKKVbGMvP6omzLzdVHPcmjvUUpcctSl77Z08PZImd7LonAwP3QDgsa
qGBgJMHR0qzd50yOrWh1DCPlofcu7/RZby2edTVSksY=
`protect END_PROTECTED
