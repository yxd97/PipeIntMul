`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAknvx1RMaJ0SDI5/CCrGyroz0ZaIP3ulW2ekFk5uxNYo4VxScoeOwEnTFY5lXbs
lsFV4yBvh5OYX7iaHNQ8OYWTrS2iR0sAMzph7nVVk4kztoah0rD676rppqBexYrA
MjxtdKRxdzhEyO46JhAT0wy55Sdg9cpIjktsg0KifXHQl+XbLgDOU46aQwmvebLG
uxoeBfuH9AIgEBj0Iss0Qw==
`protect END_PROTECTED
