`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ScTJlDL5DToy1bQaN3c3AX7uVIAy4uRxAmV57EtM7gAOej2j2k1bXCObLYR9GD1v
Og9Nev8JH5+ETToskh2MsWggUSzQZWXe88t1cYcGCH0ASM7SqAUqFk0cdbGVTzpn
lliu+5PXidbhyK1uLDy25JsDh8mWoAMKjsCh4nJsz57ckV/0M3pNgrQB19v8bK+t
Dwo8weetgkKpVLrkqERdb96O9Hrp5dqsXoK3yj9fX1EFCf93yk4cnvNiT0gugvAi
lLM8qxuCsaKj1go7eXrv95CgjcGJc6hLIvVYVw4haLzjqYppZ0zRvwgLEFej1OR+
msLLwiPhgP3GEi9kH25VlqYsVphHzZNIzgjfDuoaN7dlWmE2HvaGlglthGouwJ2N
yyJUBmfiQj8LY/Ah4g5HbjTAKCoiQbYm5ktBuSET4Wl+H95r9BzLJOAjD7fES/NT
TH1Qbr8p0qPb6oBaDcLuE9g/ZwqaPyT6zqrVb6gNs8b+5PXVBu+bEiVB7fA4dEm5
BduX8YKTcOG0jz1nlttDP/7PSbQvPzSAYqQhGBpM4FNL+49VKc5Y8zcZwN+8d2Qq
MUu1Q/O8Y2/pc+v4bFLexg==
`protect END_PROTECTED
