`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
83xPjmVdhz0gEPv9FrXZoVgtLqh7ToEqAN2nX+PzxwmTPz+7mdAecMNpnxoMyVoM
vgay3KP1fHD+LafYw+s83bGWNUgWwycE6VEjLTnCda9E2sVFwZwcnId9vP7fpgyX
KEdHFkGOC7AP3drSjODjNUwb7j6AXAArARmGw4Y3ENMozvBbZipuEmJU0MMh3DLl
2QjimrkebY3me+XOvD2JnngXz+69OGH2RE8Pm7uHBo3wasIgz4azQK+eYS802qoS
j9xwKDTnqYW6irzbD/ZBCnrtVfnimwa6mjl3EZULCXulPMwb/1tsGMzDf/o9IxYZ
wAPPYrK3A7byHR/Z5mAtkqbmBHCdIO+ma1PNaStlcTYgPLYG+Wc4fUzdwNYDcZ35
2u0A2JWgTfx3wmnDpXQwqd18iw8fLl97nkMUCZvRhFB0VybrsoJKg5ZXWwGSCh3N
dW75OUm39Xg44qlRxGsNnyntZ/YDSRFIPNLHqwcHxm9s6PN2+MsbQH3+AvK1oI7X
vYeuFHGyir4kA1bd5DZP/n1wVRw2dfyituMPKP80xHYbw3jwdAlLigXPf6rdMQMh
GAbBUzdUaZzzGs2kJBJJUWuD5AJPMpKfcVfSR3M9XyT/uDNsofbWNNCJQhKJMi48
MYoo8hISmiHQjiKCMqWgYQSBZNe4N7PXtwibzImFoxUueqrdVeEy6c/Jhykm6oVu
CF1TYRDVSHgwdEbtrS+VObS76+OY7KdYD07HCNVLkbc8RJ7wsjLOSp1JoK7R1Aor
7mGK3LWmm9OojtXbsvyFVyV9/dX8AnW/58HJkhjH24H1dj9w3lJkXlTwKaeLqWq8
VZXOoRcniZtkwmqvphyLYml6wt+w3GZF1eNFgHCbefc/USPVDvWYwW6qkDp3zNdI
+bzwezU2tooC0I6UeCsGrH+FL1mp4WYk+LNKIXEO8yA=
`protect END_PROTECTED
