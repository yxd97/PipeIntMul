`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBRvYM1vtikZI92R/bkcECpn/kv4z0SWZFuEWPrvrOa2w/A8UcP9nIxTglkXCS81
pPtUYB+4hLK7q+Sq3xMhtINav06TEUEEiTqvMrg9gzlysQQpvCK/2z6zuzWj7OQH
nPPIsQ5mgWWkEwEDV2d+SnJJMDLHd7VQmZYwn8ezlNZ2R1qIdiS2nc+wOWFPHRRX
EOHUxuUxQ6V5gCq3yncVnG4CZlgy+7Mc8Yqp4zN9TAgkc5/SJfv05RrpDRcSml+P
SldngBke7tEAlzxZSXofjwEq+cRv4lYpq5CeS541KlUa0al3wfveVaaUBiuhse2c
hzATZt+odG+oZh2ni/vgZA==
`protect END_PROTECTED
