`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RB0Ouw0ECbpIO5yXZsAoG5caoBVBl23/mAIfNMMnIh9egDAtHw8/eAbsRtrwZxhH
0KbthTf5i92ZXzuUDjAts0dpPM6HoYcEF0useRtCyXPq5UA7liMeH6mZXPa/I2Nq
7DXB5eXU3dIARwbcPpKK2E20tWgYN84RXCMswIf0WReCCmoNTuhHSE6413wGibPT
JxahpTkpSDXfBGC1mKJEHwW9p1/S7Niqr3Q/ED3ZA7b/j7Xo/mwowgcfp9MewrmD
QUJemcfCdCsn5ZsgaWsvbA==
`protect END_PROTECTED
