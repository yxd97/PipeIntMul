`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqLAd05saDqf4vmD4kv1uMGMoSWGpQBJDlifTYFNvU4nWHxPbajKEreg22wAzrDC
36iL+MXGnBk/je3q//cHIGY3sTf4hDQEFsfJj+eyMOpg3+yyqcJzD/DQnPT+bh7e
5FSG18g+HmsFkMzoHyg88OaZNF7T92I7U6TSrO5YRl+yhSyXotDQt9HWYyNQl6fg
dp/K62tVKRMm3Wc3cGSfNk/ntMQxMEh8gzsiueQgyZbT6nXf2QxVoSYXq6sTnyL9
Imi202P/1wb84lhMNCBhx+h0DWO74MQba2JEvsmt1lx9aCMwBTKlkazygiB6J6S0
40ZNBmanRVbnf83HdWqLGnlp42ZIR+p59tqhZV4G4sYTKYhAnDRx83pxT2WGtsE2
`protect END_PROTECTED
