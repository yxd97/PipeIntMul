`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eh6oRgQvhgtPC1tBWyzBoFZT66WCYf5Ca2+knG2wOdrzMVvmeKjnEMGxuZQ/uh2+
6L2OXUQ14MD8UhNccXjbeTbWWjvXy88rg4lOby+ww94qatffpYrC871pE0vQrSAJ
9RZzUEQg0SHgH8QUcyJhCCP8MCy44f4fnWWzdBaP1vlAdyDD/EA2yseUJ8to+rCh
lTt6RTSKqqp/YqzOWe9S9WyAE6yzN1VZwyG4ibag2zmAuGWizYALR0ctTQa8JqMu
tu0qZtDoizhSex27fMcfGjKULke5fU7cr4iI/yb/UiFBpBfoVVsNPAFRkZ+MIymU
937vPwczHxWDryjgaXuumIgybxENtFilPjs8yGqb727UbswXiNMjgHUfBP0jS9I7
OgoAZz5s0cgTXK8wpB/vyzIdN1bSsny1UG0w0qu/9piQ2pDWZSBT4hGgwpgHf0GE
2lAzymkVmE5jgptnknnxBYSDQpRCf33PqkA/EMAFZFjV2Ep0eMGWjcbe4kNGeR03
gpBHrGEf3nk6EuLAOykIou+MqdGSU4rLtl5QAa40bQ0=
`protect END_PROTECTED
