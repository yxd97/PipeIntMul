`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vmx8CuW/hj43CMLoVAHghSOZoOfQ1sSUkf9CgGn7KVsCBMsnooTsQ0Smlt1l78z7
mMbpr5PI9lGzU+N35OkRctYQeToZOMG/P2TduVnve827eQ+SEuByclwzbnHy2Qcx
K2NxJ07E/l0hf0efK1FpztE+v79r6LwwaZP4J2gKAZni5QIAqBeGFbR82xTHJdGP
ZFVo8VolF/eNIl4wsX2s+rPIdO3lMJRu7FrpQDeEhkXNBq7r33rXS9e5GT3/DRQ5
bkr3mUFHgFWvaS55rEZpVc+WFBR/KQu2f9RoOjWwQ2BTn0L2gN9h31ztJ2FpicPm
dsnBefymOP+L43rSBvvItQ==
`protect END_PROTECTED
