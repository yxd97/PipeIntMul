`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ot0mGBbO/RZbK512GVw0m72ZG9e8ZijeCQH4tqs+vjVC1Y7M10IPYWXF+YhDAYep
gWZeXlU5q7k0wVZg8XD8MlrwLxraWAHcUwn1OLb76iU7pwo5XvJ1jSZ8oDGITlVd
0X2Vo6UIbImdbqLQYdGsKTu2g8I8lXI6bah4y8hm2atS9OFW/HPdllTv9Xf1h5WQ
baoFaBhFZe4zXlH4AZvj9AX2xp0H+tvMrSq8FOcXAUaPDeGtkLJd6ri5k3ozNuw7
y2c9DtKYosFJvL3r+BsYgw==
`protect END_PROTECTED
