`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5zwTN1tmVpeTqmYAocPY0wT2/Yh0iLXBMJBOQnLdyQJBdO2rtnYpBQHI1RRjh+Ab
+hmsgSvGAZTt9Z/9VzBkbozLAuf+D+R9zBTjzjubGbLSX4qFycmodGmC1FOUWDAH
CNEeFUAFm5D/fi3muPzqeeNIGMf90YDIQ1pTeq5xRKN81yGb+Ced5GlVYyi2nHo9
pQkT0wH4I43QSwYMl3aKOwLUwq+m11YJlTORNjj+iPOKQSLvGTb3jnmndoqJOfF4
67OreoKGE+waSKevi0XoZ3efdjfJGwlNsRtdztBARFuFHFhg0fPep0D6MY8ZsTCK
y+RKM7N7yG7rLqwT0/7VZn2aRQATvkUVGLcSLNJg/nhS3BTxEQbXAVLheBMVzD1f
o/rk1YICPzh0e34UfWEjco53sTtmWFsYuKVofxF6Vlh40swidYaRL1oeP3bWsdhM
T3fWJ3ag5wLTv3IliqLShcfHTxJ921tzZdI8mG4B+etlGdpQtd7iJ/ohMGYlCPfo
bdh4ra3w6mHQGeaJsKFdkf8sN9EFeHAQIdwo3oSqt7U=
`protect END_PROTECTED
