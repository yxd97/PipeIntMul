`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sCJXEud0yf6vVnbN9I6aJTl7QGDnp6LZJrdtV4axmWxU2q1dn3uBKm3qlyc9Nd1f
EBOldD6ROUGVjTj+2qYINmE30rGUsO9hab1xhUY9AERlNfUFl7O67z4ebhHPMuWP
N8sIQlw/V6BCD+PlLFaULM45EtHTmB/ogwoaJtbYu21kf7SMW2AqJFBeCBQxNLZh
9ITqRTLfziJl42csLlbuGkXwOUPnQ/lrvjTH/fuCw2NwS7cFrlNqfoCSTiERLWIa
9+YC4UApkEimi10gX6R8TzyJfEZiSUnMeUI1Q4X591UwIWQb1Tz6ComkfLD34Xyc
8gp4lkxCV0h+LegzA/5YH6LmlNC75lsWazRBHJrKasfdw9HnzqLu4ijmHj7ylnDX
TQaq1VpAbiaQ/iS3BdSD3+P5zCROJ8hr2wCpgvnj+MY27fdiaWcsnqyQLZm2+Ah7
zALGuk4YjyDUTSFi0iJI6kCFzvBkkRMtK78uMV86iyiopeIDYGxPFLtVw0oIVu5c
JnEv0vyCwgVlDMoe00i9Ih0Bc7qX5wYU8A4aro/U5smroZGYVjp//Roq8AO+gXvY
xTX0p/hHGObPkU7TP77NmlvlJnetrF2UdXPoztX9GB21ac8sPCBh5nVTfk+4WtII
VFYua9lI8A99O5UWOKhib6jn4HCY+52FHj77S9dFFufcQRKqVVTPSG7QPe43YDkO
W1fGczb3FwTjsb2JILtdx6XRZq9BXd/nR4R8eTDNlnOgZgGcLCCdaPmw/1j+oY8Z
zdCMZwXZLRNnu+MQ2n5DxPMALWazsIaO7+Ld/cmPWEC/vy+UObkbYEbKNjQnHzx8
1QoCrbU49jB69Owb5+M3rCgf8c59ynjTR9JSYlQ7Vx90/NvpExZ5n4R9mFl+/KTM
DcsTiOURZcVJaKl6yBPCk3TIXtn3zSathSVKT8JeUbck3zJbDd9TFUKp3nzCVfnb
WWKOogHN9J0MxKa6xHsh6ljrxaGXOED+A4lNqPACHhk+QE4EQD3lAGmBaYS1mOKA
kj/PXyX/pF8PsEyJqBP7j66GIzWG14CPeXi9bQMfCIEcaBZur9BGpWMyQ/Iz1PdM
mfECoklUt5n7vYnjzdsL1hmOtcLmIxDtm3FEDm1BSxq/RSNypj/a9s+VSePbA3wW
7ZKT9QPrC0jEOs5fQraxSL5Amxp4W5zTV9STMFdBUwujzP2ZL2RilOy17UnLp9Rg
ALBB1/6aKC5ZiX7jJDo/kqyPZnjetwtagAHPIS/pNnY0cxwva/yZct6QMP+ZbMVq
XsARqcw8mcKrpOmRSO9SYgQ4yQA1ouf9whBTxY5K43GXReisRYCtgaD1sCWBm9pD
DrhLO4uiL4Up87rQSF1asT8Ax2myfh+7nQ/CxafDqAT5a0aoWDEskBH2aZ06kNaJ
GSjWgVFu0GXkFSG4ilWQKVRjB0K67WHvE2F2DqYmK0hM6vFzdI4GYZwKmtXYwgaS
gsAaC4fstrtrVNyklyYhW0xe6BmirEvn86qogv2jWhH3U2IAEixrleK7WG59PnlO
G8YDSumJv0n/Ml8FHW5HxXS0jxLJrNav2otRR9wuusrtp5yu3RxQpXuls9EvzuvS
NN+Iod4PmoY+qeupCqLfltlE7oyqSGXO8osZi31/FQdmHKVnC1Qw/rLrMibUHn4g
bUwFHZOoSw5L0OYEYkEVnlIswTNAn/6tlyCYOVNg6sLihpcxJ5uFFpNuJ5VxtsBp
jdKLL6zLvAimUHXOaLF/4B1iDpMc1CWX+f/TBz0maD36f3yDxBlxYicPiWba2pcE
Xq2DnpCv0jSk1ZDIXGVpOASmY0ZimkhE4ib9iccwe5ko+3EWuK8/FQFXvak3buxJ
IYGw7FiStCX4fFtFoNpBySx9Q9xYzhP+ZQSnM7PVSCZDYx0HN/0VA1d1zIVYjCig
jYD+oq+baXSqU8H8HWFvxOusrg1wp1epDaCq3X9Vvzpul15FWguyPIPxD1PJZqbN
jUOwMxrwRw07snyqwodjVUVHxnTU5Y/+3FQz7jX1i4lgHhZLT2KTuc1Q9lTwpBx8
hs3BXc7/yXLj/wFmWr1W1AIY52G0/esBt+ECJDEr81hEzfEuh1YdjQRmUlSM7ZOv
ORGJIQKj3Ywy+me7vTfyZ6z/TRb7AinTPOEzUeC+bxyfgRE6ZpC/k3xcMPuE2Kk3
AWLWayIx6rwEjNTNpYZMlnzkBwjh8/NCWP7U/Gn6KTSikBSokhUZ+VIqAhpMbAu6
Th2lq7PjqFkNbZzzCDVZ8BJiCtTQmLtVUR2ez7zTRgIHEzpKusrPCBDNo+HaySuI
vCZddq+ulRO5m4cuA0P2vkz2JYaqgpunar+eYmSr16+AQDHhKaNJvl+TzFdaXYpG
gM0LCVt/CbQ345bb5Q4V4whriwZp7HwwyLXcSMVAhQzya4SgN8JwGa6gRURBQTeN
uuJtCZx6f7dI7lGhY7YOJWjC1sSMlYQZkSXJKCmJOQOzUhwHSK2gdSbmVVko3uAv
ZIybWBHQuiTvNu5ajLL4lKpViH5zKJvFCssK1ZbUG9fFThp89bA2Fep1hjP+agVw
TEu560Q9nzz+DMMm7i94YkePgshOYP4Ngs30rESVk5R5ILx/4jqqaWZvF4dnVf+/
9DlDGoJN9c2mLRD06BrZIpqDV+sviBVZ48WJICD1dwycpoA6okGdJk9byXIL8DK4
Pc8TuU3PwiEXsqqGdlUtQVoMPI6BViYdj4mSL43yOXpcyy6ly/Ve/5AmPaXJmhe5
N5sOpafXQ3lDZID7E/lYRVFhYxkHsdAHiFEQ+1Agf83vQi6b7s8A3ZC7MMf+3VF2
x/5tQxMjqnEqkhC+fifphrXibd56QhX2m6w9tQKr+cHy3HH00+PAmz51/BreTTKJ
M7U99cOHLA2Ekm7TfhNNPQN4eDjtog/J6qR4Rq2rxjg=
`protect END_PROTECTED
