`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2jaOW7PNQbR0ckdm+Uj4ZbYKu2ZbBhSKrovlSUlkebAoCMIyNWObSnnjMq8+iA69
Qk00ziKTaVcFkhB9zuzR+v17E1bX+O35Uk6SeA04BehaaFHQH/tZROwawD4jmw1g
b0ZfRUmJ5TXgJ2K679AtWQ8URwKeuK4bJQCIkNspNEuF2vW4R5KAjr29myuYFXoX
lz/DCua/c0VuFHWz0tT1cxMuCK4wRfIvdZBjAHlsJV2TWN4fmAfg350d1LeIsMst
8TT4uFXZ5RKUTuB28dRFIw==
`protect END_PROTECTED
