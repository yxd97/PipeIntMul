`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3Egyg7kvEX+0WCdujvczBbLNotRdmrVSTFZdjTIQsN/sp82dTStZDFXYcbvKnG9
RqKJQLJEIdtMgr5CSDbQ7psr3Vff9kyvgxdJZqq1mz5yp/ZL6SP5yhpX3RaigAYX
c91eUzG7xfdJg1j9GEz7K/ox6Rw1YDtCUMYArpc/OIzbP3rXmZek+ydxbIZwXOPm
RvMN03oB+q9CxpsyMqxyxXIUsr+vKhWmuvSa99bw73id+CTZdlTB7shFO3g65YKO
TI4jfVAbz/1nyFktlZO7yyhk+LOciechRXv1fppuzvhbyN0reB2gmqDWBWHXXZW6
NeUdAY03TA+TZ9y8Oc1bE+5IJzpNrtA/p0wRol+kAd0VtPfsR1OJYIGQez31OuPE
NXm4OSpWVY0vFsFbs1yZih53u1wjC2DKzOgPz/3nVbsAejrO6B/Ks/nqMhZhqbZJ
epkjT78ewG91E80V3Go1I5v92zBQgxg2cz58/EliwzCgdd2T178v3thoG5wuzb2p
JMuLyaUYg776IxXA++2cd842/OxHQ/3BghVm+Qoe9dXcDHDiWq59JmmhWmIIUqZC
mnerSDvJF44IYYmVErCBlV+5Qjt6vwS69D22AhHqSX3Q4yfF3UGLMccnF8QBohLJ
P6SgpNUaNNPimJcsdaGTDQ4Cw1NqCztDE5fxyswRAPkzwYpAlVTFze5NVHTKBkY+
5J5RO/mN9S4ogSzoIAW+p/nO4Q6p+i8+zABucRRmYDLOEex/6/O2QLR8hODNTmU8
Jpwryqte9nFJt5uU2uUtYzNaMRYOgnMOKPkcGU5S4Dx8I9d47CzYLn9YDwsO6Kcg
O5jJkdr/8cq3ZZkjapbiXmv6HVDJkN3PHnpjn65kR7J4tNMdqQ+K4Wl6TOMCjTZP
usV8Iqsifwju8QbGQiZibidpdHDQWOWY2WujujY6cVIS22R0amKR2/s0QEzAhYnJ
sAePnyuUX4w30b6fiNAHMgO+cV4HMB2t9J+XdSjKQxEdr3mbsQeWZXt7k5PI1m9e
2vrpfNfUCr3+hzogME0DjJQnGLfOvorl/qvnZnEWuKV6KJwcchPIl9VGM42euD3g
Bf3/yhGthqMRYKk/5Kn6FfntPaqfLCmMDLYwjgi/jxLFE6KwARB38AT2jKDoHLM7
zwm4JluQWPbk4JIgWIJuEvgWLCC2lLvP+XzLrbhSb3V0C+uNq6KcMsNnFjp9CpzX
`protect END_PROTECTED
