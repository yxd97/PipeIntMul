`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2HFeCCUw4IdrcWX+Qgs7HUqszstHu6gX2icTdtbEJyh4iS/LkbBB22188vdZotE
liyzOrZIPhNmPWDUNiiiSLiybmENNrvt1JXCHIu+Sc/AcUMYYiJralfqV1SiDNCV
nxSrxA0dRwcsTF4md/+5cvIOaaOSoDxlJq4gxzxm77lV6fqeBlzUNLyLnitlxW7Q
xKhKmU3Lsm4qyti8Beg+iHe0w2zKg7Oz8yuHn69mEX19Jvdyt5n7d/zzLvUdz3OX
1nqEm+6rRVurE/gYUvtHeQwItJRzDjhV62xNSVWAT39u+pj7RPYCZCxS8HSgzdzz
v0vh3aXyAioonPQIuLviUksIhEsuPfiDyxwAw6PlJy8A+hYs9IeyiVE8DtGnDbqy
rT1eqJYwlRBYdHAbuii2R8lJUrn6G9jGEdPRl9sQQBc=
`protect END_PROTECTED
