`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PIAk4ecEmGFOPPLwDgf3LoBtyghneS0xDMIweH7bGhJv519l58o+P25IWucDkdLU
Rv1TtFY/gOCYqlG47Mi9FuKDWF1ldxxz56mnQmXeqEgnAnMUBJwrEMb7xVNs5WGW
3fco3SZ5BrOAEDlQc3+pFp0zJK/qhzzNmk5HRHySmBvhETmzmwqYaBcWJwCWEZhu
wt2hs070Hilo21C9Z0hFxS6847eW5ggoiwDGxmSFzRizqpZhqF4k9cynn8MP+bcl
VGx3UOV4heSBJD5pGv0+/eZAYH9CAn0D3TJkwL8JwQLVXZmSWcexzmQBb+wGX9BW
ZKZq25IuaA1QTqYBKhF6c65IaKYnrEgTEPyFAx8Gz2G0Pk65xNikd12b9oBF/TAD
+L7DX5/EYUOrEqCdQ8NQCZP0L4J4+8s1V1R0bRCEfn8ju2TTsBeV3Mbfzckhnm2u
Q8RX9jY2gCj3Luza+7Ettdy64QlqUqVGpzBS0NrA3pw=
`protect END_PROTECTED
