`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjotObpiJcxLxCrFKewUU6I38Nqk8ZOmftGhqLULrmbwRv06HXNZi21DEjzoj4zO
1j5TELhyRVYQaCjJcaZJ9a7wt75ebmDa3Eqe+esjpExlEk0+svmhkhghsjIjhDwe
BFtPOHxV0B7oHBA/WXK8NmKQeOAbXW/X1w0zRgC2J1TJO+Qf60zFO3zs07OzWhi6
ojE3UYhy+sbwhmtDRZNjH7+FzXT5rEWIcVc4sUDUeZqb/DY+gaFdttHEEjOFjgsw
4iOoCsPe4lj8lkqbFJqlWv3Masa8DRMSeI9jglpMXE0Zq5n5FsFrXOivKRUkEznJ
SqHs2MyFEULNnNz5x5H5uxZz4JUtbt9XVWsx6YjEKDwOGvadH1sL01LynkudefG/
HRsADcgJ5PiSxepz0Q5Dsg==
`protect END_PROTECTED
