`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4HvDNTHWGi5mq5R6aXkT7SMBaIlYJdmdjaH1/jxx0V20b/GxcLOIAReJhSpjG0FF
TnlhAjnl5myXgW5iyT1Sw9zrehYKhq2Ft/0yBy4hWcytf9cFIPWX5aYmkHQ71Ol6
MoO7WEJ38BX2NnADi3BD2/DXe+iKdfBe/fBCliSjBNYfvZicfNDVaoJc1A18z7Iy
9+qSQcQj+FuAIicDeM+yA/Z+8zcpkKNoAH8E8mqUoy9mhw3eO2nKSoogDxbwXhl2
RAnwABnlOmqeIY7WRAKJ2Q==
`protect END_PROTECTED
