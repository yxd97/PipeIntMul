`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IZiz/LEN0idaOD4ciUOLpR71ZE9ahWXMc6yTADz9qPrL15SN+FB7YEkjX3Wpa97h
IgLEDAGaVf5f7Jg1eA74ZNX26FsozjhPDzh7PbIZa17jafeur1Hl0xNhCkm8hmjJ
pzXsMR1PrDy4Pxv+25emI+nnYVRmdUmDRFZRJldO3c0MYjTd7pr0da34ijX5o7/V
FMr+tl6zkuslxPY7+RkSO7wIC8y2trTGiG4paFLBS86UIHKRM5GdJZiqvht3YZDQ
diQ13MXX3J+w6ja/pE3FWsoIjrL5BPp4gdcBM3i73UKzxLydLiMXPE+hb7dbS96C
xTTJBdd+2cPnEgc418D2SVpplx1kOFxX4OtYCHaBJLzm2gVBl5pPhHyCbZjlAwYV
nkeIoctSCIUs8xx6ldNvovA48xShDv+U5EHdgcqoIwBb1mrjkW5Y3pqKsUc9ExSe
C0o4KIlc7ioKSRpCiPGQ2HmKZXyEdUmIMeZtMEAq6B27U+Z6pzIn0qyXBnuU/Fkw
484r8ipfcHy4vvtJp8p7+KkLmhJLKpayq518/UvL6YhWeKwu606tx0WNdEv2z41J
Vg0hL4EM3Ng5YSgYJ4Xuhw==
`protect END_PROTECTED
