`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9KG+sYgd5iYHIv2rxyCbLT2LNgy2ESRu4FvbdaUDiHBoXlSwbZG4tIHLuWIy2hJB
Ed7Cc0zdbPy335eW/fwymCXhy94u8PcZ09IXNweMlyJWzIfpcI+vQY16GvGFVH4Z
tT7RsInv/INxMJr4QQMpXCfBWHUKVCP9yZJ+NHOBB80eNdajFU7+wtgXrBZzHeLV
y3ZtpcpUoVCpEVzEO2I1XQeBegIu4mOYGGR1+FPfQa58UmYLqIZ/6oj2H6xgHywG
GFNjDjDwZmOBdKm7TFhelGHNUiUimylFki7zRk/qX1FmERn0YkVSQvL7NH7nGDrq
KrySRFW2za9Bce4sqBjqjEylYxyFaoJ+pBFmSaKAtU+a+kfWhDQTCusPBasd8cut
`protect END_PROTECTED
