`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZWHk6U2xvodcSPJGZMT0VLRWif4SZSF7U0bQ2CHygRyAgleEgFSP/ZlBw6ixVv81
uRjsVh0gtVGao0ebWrEfSs8nCtOVadeuhdzVcCJdZBHHCA9LS8F3Kbwmq8SbjeJT
khMgRuD7hAQ5uhjJ1YKgW1iy7WTZopfgMC09G0Vn+nsCmk/VC+2s3plolvo5+ivU
yQVbr4pXAflJuxVL6IdEmyVeVMQfl7K1T/Z20NAQlFNpjElkIxXlBjzTPEb4oHNC
JeAqltG79NP59pp4nuz9JA==
`protect END_PROTECTED
