`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DBjaLpqSTTy690VKi6lClxiHAFxwWY4yEAwNSw1jfXcE0DaIf3UZ1qgofenmqpSX
gnzmOMUlsufrYxMxEMcMkG3OnGTRrXpbtdSBn6VI1bYtM+Xktt/yjoucHBJ+YTMS
dGGSUnZGFwbif6+wxDa3feV59gKLi1TOeSVQKOUwEQvhR7OkzQYU3XTp6AmNbV5Y
SB+cV9th5E8xiZIVQs3SxYnnNNmGM5t/vNoTHX046d1dWHxY/kcBXzEHxaLObOqo
OBW7Zw3hHBGP243NJY77JCPy1zgNrSfd87W+9IgPSF+2krMh51M25ITogcYpoP69
kKQbhruuSDp9zj66sAp2Q2H0+yUHS0QBsUd7vioYZKHxpSkjpapthP4iFoibnffZ
J3W7HMS6DgBt2NE6dzjYfuOmL4ftGtxxyW3tmyVvtE0KVvShKBcQ991dDIIaIShx
5oBa5FU0+zjwwHL5LTirC7twxfPtoYjo0+3RXVEGXiOLvieuNolxw5mbL9HGMoJL
o1+oAkdxJRiyjCDZMjeA/GEwcjQ1RFUlnnKfhpYcs1FQ84ELR8WW3JwD9aeeToe/
`protect END_PROTECTED
