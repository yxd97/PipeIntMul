`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nPpVjHdZPNrdE+lLulmPRYDYsWZcAuGrBRbcKMDFizje8Lyk4iR3ZQjjdTAO+9w/
pkUESYG0nTptzT6e0d9WYxdg6VDualobQJDKuUYQAPj1x/w7zVfHB0am9g1j/rJW
/U3d8vcjpSYp6BxzFqPFBRxgMV3SNwppC9UqZJes1zy2i8YZOKKzeIcQWN0weuor
5TOKqM01U4BIpQuptFFhrZOu4iNJwxlKTHETbL35aS7N0u1rf0IGb5YCmJ0rf31Y
z1EWAktqG4Sv2KRPlXt9+g3746WPinVaF+49NvSNGArJxvr18Nf9TwWKcYVs8rf+
0oEOlRNqWMA0xBv7j2N4i+cPhxUt4YcwZWTj5rmnpJe17Ms5szEMZHZCBDMO1kLK
y+4X1jHj6RZNjTT/tJBVYGdB8wT4abnyot3awlW1jKfcWU+66mouEvDbw9UgH0uI
TmwONA43p3b3Eb1MarlOZC7rR9AIzK7xx5LhWnjf+bgpQ96Y2MjKzTWIPqAg6M0q
Zp6qmd4FO2r2cc/2Mh1/IQQzpfJPCzD+d/RYS3Ln+hhBWEi6CZOpA39mtUdTV1vW
5E+3lVYEDheZEPFjrt5sfpAFO48ZF6h6cA4K2JM0QAM5Fk8EAewKEIL4a6qdSg6p
YGtFAvkRb+TzfGooFjCKTg==
`protect END_PROTECTED
