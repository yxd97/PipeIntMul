`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hz6ZRUgngx9U1JQUmFt20wkXqo2HC1Hptd/XeRXRoC3Ii7GZEIJVB3+nrVTtX4+1
Ja0utYqplFrOOw9NKw9m29mltqSDLVSW1tDGlk8QnSkvS5h+NM7u3oM5BmAOqPME
k65rIJWCYSXLJCLoRS+Bs/f01KrIVgkQX6C/xf1MzFVussEBvnC8GJb5s0EaQMYj
6IOKOSeINQn7JBhG5ZeaFj/voWb4Xv1FKUwS9Qy2pZA+wYO0+rNd+Tb38TP5xOHJ
483RIkmUYJo3dwN/VPu0B2xAgxlhy+YrxbdOgF3k2oqjOZPs+Af0/yXnOxOvbRPg
/SLVHEAwzdlrE/rwMW6XHWjCMTRyvusCrlIxuNTthzH+uBpSrLyhPaBig5L0rz49
8QdJ48y927rGFMPHXrQx9tlU0hiPiPSnbj8Fg1cMGPLWoIjO97MljOcyUpdpv+lV
NKzKrid/IvteZCor2ESc7xcRr1RcI8fV9FwTO5vlbhM84RJMb2rk0SdyN0WNulgz
lrqAoTjSHyWh4k2HV1Zvc8Zfr+x9bHo0JZyeXQ1fj+yN/PRHbXr84ofAasGH6D8X
Xmi2BVHTBCze88Vm9I1A95dZLkGUMlGLvziPXyxlBO/CmnSGVPCD0HPiQWWztS7X
SnS6YMaGPRXdNlKdYosyk6DOrJiZP9+93TjfJANQWQvf95BYA+6muqkFu1C/hwzt
RYs/aThyKADtb4rtPk/tCy/8lY8U3h9CB33iHUbAdfuCDCCFO854yn5XpTUp6uas
BZShSR0F8hb7Z+cQ/T84lOldi/p9IWSJE3xqJmduaFGX7eXaLzx3nXzFFF1XQVOh
IyLoILXbYo7abTZ6dIYjumCCJI32bmAIDoCDdxsMTwbt2eSj5rD0NKrkoZt8WOkn
T17OxJ55N/bqvBDYHj9QWNKilDpKEcsxS/5CpZ7JNsvxIxSJgeL5tGX1o78I30dK
A8dGTP9032DW4rox0ssyo1DG0pLWrqAso3SBJF0OFnwAZegqMG9t02WcZTPjMjbZ
LD4f6jRSFm9o5VqhttwlZZxwoORp7swG7nWt+9tEWY1E5YzXVfOVjAcvao5rX+Xc
tFfabr0mF8LMPB/2ziuLvbrKMK6bMXu2JK4pwKEgS0D6XkT+oo5CyBFyVTeMNMpq
fMDDV/FD/dpXaupkghzxh7FHJ3+U9SiDoXMHYz4HFWDJSyK8sTjs2VkSjYykjuKM
sWyWq0YcCs4tqcu+PmTTDxaA8slRLGo+dPL4NMuN4PA/tCL1qSjsN6VstsTGgiyx
1a4lAcoMBaiSr74S3XiDMVFui9lJPG8+SCloYiZGbccPiiIsOUlbGnLDI3BSW2JZ
+vIsuATFf9utoC/mXmPpXVkBU9Rd8cHNI41Q3ue516okvJBXGShLfRjeQj/KddMK
AtMKpFl2U4wFMsq8M7r1e9W9LCpC5n7G9zxcC5AP6RKD4gAcTb2T36GmgFhy66cN
SjMiNP3/tMAN8LY5qaSjaSimnLzVWBy046CPa28B+2Ft8kaGFCwcNr9wstP+0hWE
qL4JwNvDYy0qL488mX+jU24eYLnK0IC8cIsgc7BsWUCUxCs/TR4fgD339trIp9kZ
RCKQ1gby2QZ3IaQfsLEO8vOW/ESUJIs+FpJS58nN9c0fyobLaQC4j9UrAfKVvPKK
r7oQRrfVc3ugIrZ312sBE6NiremZJEK6jzKadmMieYIowPCz3YBZ4xrKDAcYkp4H
NANmzxwh1C5qYTL4rUG42K9dw+W4PaAZ2PClxzyqszqQ1HFPHQlE2ViBqvRhpcK9
I6rxwfehN/aTb3OhtzEpTRyvka6+GUzkAu5b14mYzfXjptqKCKz6uXbxpGJ0xdUs
mybtoKv6Ee/75aZtU5AMnolj3I5xpwkDHIoyiMqG0VI5AQJ6BhluBZ4u5sNWaa9Q
NbgvWWA80uqJmWWrQmA47g==
`protect END_PROTECTED
