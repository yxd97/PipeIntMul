`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/ByPi+q52/7YZ2dBLVPtTwdcU42YZI7N+wn0XHi/3X07MrVAblKj9NEWeK3FNz2T
UD47SFCZmoYuxO9oAnZKlVRuV6AH4niR5lGHLZA4Oi4oY1rCANCxfm2/WR7+8ITp
YK7OsX6h2VjgYsosLptm0IXlpPpdIGw0Kw2yieHmNjzpJaHSrjw5bo+NragWoghk
B9RhLKcflV+mUiqHqM4kB/NxroXVbXaZE4PZ0qi8UGz4rM1k0vfAANp5yV/ypD2j
3MJXrkhV85CwlIQ7npuGMs4AOT+nhJYlAj+JF4qKPG7u6sXRySlPRuUrPP1cXtQt
cPH+gN96IagRIBLndeYTmRC2htuQuwNBwi73aHTeesPKk9AEg5zmGgoSCgxsYSu8
BMYVK915j/RijgPNl45MDBUOtdspxn4cz3ENkVsnB5YMoIdU1E8RoI+/Nt2b41Ab
JV4odW5Rq4rk3bgqHLyPQCvxlyfyUzv1xZR7Lw9kFWGiI6XG/w2ffHDYvRtc0Q7C
VfuRiWlC0l3CMSCVnnskil0W5JCm9icDMXh+2qcxw4alGPL8hwp8ddTulGIV0b6D
GUslrS7n7RrSFBVTHUSXUg==
`protect END_PROTECTED
