`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x7j7h1zN11f0a0Wwju9/wsfrxh/zRHqAl8NBdo+U0VfawMSq+byrFe0AOvTzoQX5
lUScDymtNDPQ5sIXS8TyDKq1mDwNcEgbSDLWH9+0+BsPl8nWRmE7WJj4wHizYC3G
DaWpOKLUy8Vbblj4bgoPmnmU0XJ1CK0bZ9BENeR5r8OOLor3KL9bjnVJ8TnZ4TS3
e1kb5m6p25p/4OiN1B7nUd4EbaBCcaOE/jGTmq36gV7OnKasAAv6vOZusCWwVpee
/Idy4xAcdclSDqw//Hie4g/kt9PudjMSHvlR1XrspGk8NKYkGhzH7aGI4TiSSFCl
hp4cFFUBpDreVG9pEJ4yw/NcYFlElFyF8J9al7Zc2G2GaXLOW3nSEq1GNHZ87dtz
B51+fB4PVnJ8iQoFTaEisSa4zvjcJ11hjw/JvZCF6BT6nsYD502ZrNFqsGd1UR3t
FSa+sKIgWyUx88jJCe2/2J1F0QlwKng1GxyH+ucwutxT/qyhCPlEvI3CQbjZrxFC
`protect END_PROTECTED
