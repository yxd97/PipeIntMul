`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HEFk7IyyRSamwcw3A6NOtftqjqDBve6e0Du1WBsVmX3HCzXKdd0bDItCv0y0gI9w
mZWR9g5EnA+soW/8/WGjxOlaKRvmv4fF9sfgy/TJ/GhqnqZz+LRMONCVM0qJHOjn
CY3kbf1nksqRrc4xYWIDU2JzYlUohCE18xBPQ54YzHn1hguOyEyXhsYnFxlD1O8m
m1l78dAcK9YHdh9diny7nHaBdU5ZLe9TM2tw4sHQZGV1YDwFx4FS03WCj7u3mMnA
8ylBypYmCRddFsG6LGWgBjGEVqlHTPSUBbRXPkP/v4RhKp6Rvp1Bj9Cwwm5xFE7M
hgiwBA2A6UPwjzE5/QiYVXZtO9A1kFPhRujx4yst5f6iKilKB9jqKvNtA/vVaeid
Ck9L+d7lgKE33Idq181oDsHYop5xjd4nM3q1p4ikJ2XryvH/XJt5P0tEf0yhSmPa
dM8ykc7yGmsrQ0C/cunkb4RQ9ElL5hr6fTy8JlzDtnzZK+BZTJHIM2H+cvkuleks
YhFvQlqmtVEnOBRIjquhWo9ydB+cTs7sJxCJ5VZn7z/Z6B9Pd7qsuwQgVvsaWD/E
P1r12LhLsDOWursh7iU2+G40T/H/hLw6UhI4ggOhhS8=
`protect END_PROTECTED
