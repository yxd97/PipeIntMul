`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xE2w4wnKU/W9AlO1/mqXBReZdk7K3RFPLaKG5UMp2h2ecwpem2cvVEtnDUjOFBzK
sZZdkY5nu6H+WHFXqtwhqyEZeVT0ZmuZ5XovkhGaWtx2V0ms9DH5kuFNoQLF4zUt
VbhQD3YjHdiXSVzSoEwarZyfkg3wifwmVN+M7Vj3Bms0MnonLjujzuPlsifzkqim
3bLdiqY6kpg9OvQhjr2SVR3PEX5DhYpUEXS+Xes+Wl3KF2/zsrwc+1qp14R/Jr4N
Xy/hhNUvgJgfdvCckpDcvMuo0FgKJru9Gt/8GguHCD33OFRyedxYg+VeMQ3BtJuY
5qficrYLp167m+7LmQ7cmowUvUAwdmwZYFUWfZ6opb3nCtH9qwXcBfXd2CwEWUQj
qaNlOAHPpKZcB+pvvev1x64xTm3U53RAzAeVFHSnvxxEBuKeoT5kFoOE1IHYmRCR
Qq5hIAGKej2VJgXfymWyvjKDutwYEN8/brIG7bhPHYMgfPKHnkn1d5eqWTHUacVf
WMagfIzhM2DdffD53aXfx9ktKaipRGoUwTKy0IjPxxXkSlF7MyC5EXNZjr9DcaCk
/r4hkVE0Gn+tItrUnnPYNp+c7zrXYDRyx29pCweTDXE2yXkyB5+YzNh/SLmxQ7fU
qDE64jCBionnXQUT6EHH2YZDnq0zftMw7wTdbASX3bU1Aigul99LcPNZUCQsqtDf
5vTX6md1Y5FQPTKCko81Vk1RubXmHldYYU1ADZgbwd8=
`protect END_PROTECTED
