`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TVHslhGTqr3KUjUGM144+tL2OvuzsNe1TMy8PTDTtyRPKxALPZ8q9AodkUSM+IBH
RZZKFR1K2Y+IHxBYGgu1Nm+wOJ1DjXl8KrgaVeYfy9zfDa2ke2Ox/resDI7SPLMI
RIetD0wFe1gMkjabdeUYHZ7qctz+Xkeo4JeUxkBgYlEYO7K9VFmo+DTy7Po9bt8N
Zh04YBPWgpQTEYvA49IEZpBSW9xrieOyveCfGfeYgJrGPFyK/kmxopNOH+t43N4E
9x4QFMP1CQnnzwLYzqtGHTM672jcls6Y+hm75XreODcfduElXHrpuN8GP6WaZDKs
OrtQGKyev2undriQQXdYJvuqDCzwSjsLmhrtUqqa0YsfIy6wjBNMbG3e6liK6nCg
usa9v/rcCYOBYHIU6+hnCBfAiSF28u3n9AGtde2JO8INOmYtdGOg1HglSfnhydI9
8U+ZGVsk4cvQC9i34wL+9U9Bh9XRrkZRNDc1bAmqvUC2KwaYA6PMTPkOBgMkLj/L
4YnW9/pLRZh2VdxhHqHFytW7POzekrypTTrhwi6geO/Zv30ekpo3x9HNbLdqa+lW
kS+ZVjmD52DFdkPm8pCm6S4nkmjrMh1iHOh8DzxQoGmGCtOWKzaK9QaGWLtnSOIw
3z1PCYJgmI3lZt+L0unBbg==
`protect END_PROTECTED
