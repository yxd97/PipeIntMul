`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j7QM8gh5LFMEDJ+eYajBWAwLDsc2K0cnCaq3SgntWifu1AIPRZU4Ev1i/RJt1TvB
JKtJ5eLGEnjWKWZSnj9s8q0eYukcpFRQddncg+uQ8fICHTsVbt1/DfKM5GYoo/qZ
Vq6Ff3C/4eC1x83ypwgCFw1UVE1YVLJuJaGw5IV8pcwwp+QnVKzg4ffY2743bNsu
FTUBYFpGzQgbDBw/JALeMhxvvCo6oWnPE9LPQsh/rVSRL1Q8VzGwvqd6RNQyOuix
OCw7FlJH/aPmEfjcesQK4TjcA7qcHvDvowliWyKgC7kwMahDo45Pd0kZ0X326NTk
yOn+HhzLFxyerFzhy6uAOvsjQPBhgxlMygX2MB7nu0IMJlUxMmyujHjGQ53PU5D/
wYkd6oLuhtgF9BBI2mFQbw/ZHEEn2mwDB6qSh/sKXf2cNKqfBMP1EU1G77VWYJfd
Tp15zZaIIRxdxjYZ+NgyF9DlEeCNpusXvoEJIOr7GNDLGB072F1lHopxUK5w6D+G
t7xHDcQRBtIDgSAeXVwW4SpRdfFxYk0FmiOC1OaW6vb+rWKiUygNcf/rWrwdJ8Di
ce+fO9GasEBeekg3o+oRu+06wCvh4uYe+gZL1kKLF+Ul9w+/NeehN7ecqBvyvunJ
QCpjWIJz16x/dOXUOHKlbgwrnTNZgA6Hxfxb39nbFDKLz/OjcXdmW2lxxYADHJNx
uOCkiUuXPDO9+RKaJ6Nib/uGU2z39S1p271l20ZsPYWZ/kJdwuMIIwUABkCe5aaC
tYLG67kzL8QTMaibjHWaeV+05+cPcsipkFJyJh03OoBB6zqoNFk4w/jvxP6KMOPE
`protect END_PROTECTED
