`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/WBfLLVI0RSUpjU0zMtcmgaEDLTv0Unw3RhxfS26xBuWR3nqgASiuF7W+hzyrIS9
5u+Q5nTizglsmxitUItqkaefEhVfYqG0HYO/xS2Us2RjVTvhHTJbL3cuskWJB3BD
J9SvGZ5ngCxjv2nnierY3b491hXj3de0JnjMIKlOCJLta6iqVWiPD2qBVnnVZFDM
0OsgXv+0xAu7+LfmD5igMW1UT5q5Pv6rMApJY8N8g7wbQ8DA0Phubz0+sNONtwVQ
X6pmCgbwV9ymw6zt9lmhb93p/Sk7ge4YQPVXeiuz+G/2Tva9tmrBaoOGPM3HIfnJ
wpuILwkL8W1tauLDM7MnQQmJ799F11x6yCXSOcan6b2+fWsZZ3k/bgw7B1Ea0gzl
88w0NQgGCRIkn/BJ4MsXtKkOqArd7+HzAqmpKuN42UuaqsTmkscShyhAJTmGXgAq
IjEo10KKIIKnW7jxClTeK+gioLCmXCQpNckp0YKcSDkttWmo704zMYVsfp/t+rpk
JNWd5xhe/wrtuAjdfPf7EvyLW0lQeQJf5tSm+bqnYathKARjGJkB2zx46mo8mC9r
HqqbA+Ktamys6eVLPc/H463eOpJBFHbDBTeczqdByFhoYsmpNJXlog5gYjR15kXT
qWVEOg24Wjf/6ATEXEkZt8SFXf56Uw3gOJDXV5LDQZ/H89cx+/IBI+JCeho8hcb0
jXX5byqv4aM+WXD4rrmmGI28tsb5wZQXLeP008p/D5AfTowelKbtAMatwK+7t7CZ
+mvgt8hENUZ/Hd7m1Eb+AB/ybHjFKE/V+hqLbi9V+d2QcaRYQv+H1uHTgrG4Gmnw
e5QN06QaTBvp78fygR/K2QgPVIpr/c+y7NrAYPJrbYCqKtTtilZZ3VyLyu3rSenO
qQYfVP0V94t7n/BVlKM74gZ0CrM7Ct6xgIMmkFwt6lufz16KC1uVFW/rSum/8Ty3
kYjNbSrx2x90iV/grtjYp5lS3zny2uDGELcLqU6PuaTimLZKtPZ7B+8B1L/d8X+C
aoVnzkr/nG3XNG65AQ0vu+iDaGP+TmKxQoy3jTYyxGSzQ6TJgtkyUh8Ohr9fwwEq
9GYBMJebdhmYpILg+RPv1SxufvfZV3ZPEFbjzKu6L8X6TmnZoybKdO4hzHjCFB2k
wTbfmg8H4Nh8Zna84jP8/+kNkTIRvkCFi8+tMlVhWxV4nzrcbJ48rhTAqZmlVtvo
P2gcYnfR5I2vh1eQk+bXLV1m2GEGjraLOUVADl4KytB3oNlBwI9DUAE25F1ZXJJZ
ub6estsSVCGgTfJbv/TQBiR7hCZiAHyUftQGqkypRbhAfwfiiZLxirse2OWH24JE
AtP0ZhSFfGGgGw8CcWFu1WhPsjDGNtqyn/dSnlPQBM+Cs0i41EidVNBBrTguzGwJ
6D8nnFlNw49RrFwXTvbgw8KWlbhEQt5MI6L8oCm02j2SOl42cjBVfZR8ciA4x3lb
T4bT6subTbCLcnzjg5f8QiNS+BlxKIYjHgxmBwENQu/NMAuolewDMcGeqHkxOPDu
KBexgdBz6C870SVpn14ceLDLcIK5frVUnVnTbhR2zvkOH9HqQhQHdaSZ46/K7VUK
i8ll4VdVRLAfHnT0ajFc5tEED402J28UpQaLeDceytYij9hne7gF9cd1kYlHV9T6
/PKDVoP6UT0IlDYwhZbyVvuO8mzgokr9lyMrqnaGl9UcxETLfcsoCDyjTVk9VHZK
nv/ZbQ1O+wQtnmXpifV7ZjflzXC/kiuWJDccWCTuB8PMd5e12LM6Hw9ug0EtSRRF
3zZ73SrZFp2Mw0tJMG2kl93L8LWjEBqECR4vWdlqmzMRFDOHL16U6PU0Zkkq2zxC
Pd1i4XvJKduEk9ctPIUwAUwuSeDpEZHG++Jh5kTR2252ABoREhtTXrLt4qdWsPjo
gIlM3eUoaI6HAD4TTHXkoDnJS9RYWlm6LvhHQmgmuUVUyhPWpg5NHVyjRMUbKTF6
wF1IApHjMQhvM+8EE08tENI60vetdLIHINe+V/v7kCr/pT2GrsRUZftFU5S5g2Dn
VN/mKqLMfT2D6VFszGB9X4iZCtgDa4SN6hgib9Viz3QL+hCdIsFeIpQz8Mdi0qwL
3dXHWbrxQCkz0bOBuvpYvWQHF2r5B+qX5QuFEQ9VBlkppMa7jzn2IPlRqXj04QpE
B6vvMe+gja08WwztL8r7dcj46qm41vCLzEpSmCVY6r20DHihh3RcJKGqnMdNA7n8
x+vNQqMH1ExO0iKeMF0b2DIDd2Ia20znNkcQVxZ5u+LrEaYLiI8Y17roTFdwTDw6
eC5l6Ikq1L4rGkaUbZ5qbGwbje93BdIsRBS4hszhX2fX9va7rb9Jvzr/7JoF8wQK
Ffq7nI9T2P8H+vnw9hbaiJiQcMeG+jloG00vPKO6o/GnbaEyK0WpHXBok8UVufPw
KkgRC5iAdwmi8zrNijcLoo7lYZtJlTyazMJ8Q/YS9ZHLZpbVcNeUMdrDqKKuqozL
V2V0XIKrJUuyWb3ZQOnct1U8eWtcXaGLQZ6sYZsU2kDcK1oFG9Ckg3Z+AFgrHqlb
Ws5X5fRLmDRALHQO7LQxe37rB4C+Pb912cC70N1UbSitPQ3NYtYHx6/nvc9RRPPZ
`protect END_PROTECTED
