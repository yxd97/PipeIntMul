`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CiSAm7k1a1BGSDizW2PsBqrP/j85R1yFnmYFbpNL7JkilPDjnNfzCBX8fVhiOfDF
7skr8AJcMSlYXvV0uC//tixdjazvJTZwB8SDWiN9NuwJa4jSPDCEStqGxM7Rimd5
AUCIADwsu/WeK4RTfuXtMGWHSqjRKhD4v+wS/j7YtThEcajFppIu9iQw8VShWd4l
S5yEAOdS1SiwB5IfJB2TrHKY1JOWjgsPAO2iw4x0WxBGFzyPZCyBUJkCDB+/wDS8
ff67x3r7kSpAuioL+FS/XFGGEO6sRkHs33/Epc4Q4HUTKGQXGuMmCcdlWP9hIMJe
5gn8T6aWdlD7Z1WYBaO0aFZ/meQlvRbfw2Ksg3qLpDT//thttu83HpQQI2S4BMSL
aE3dQGLQoOFu5gsKJL0Ats/hRM3xw8kV9ZL/rn4ygOT9Yl3ipGLRWlBpwAMiDxWi
rNLUV31XwZHfoc/RW/8BaPgZqI/eErnmo69jWkEKRA4Aekfvwrwj7Q03xfsQ6xQ6
QLCcbyEa5eNJ5DfzAWUKQxJ0xKp8YQ2WJQ96HoHfGfhIJJIkXBCQb6CreT9AydmH
rlcHZiBBSRYVBaGUeu0nHWBq8hQZ+YeicVLEnHSJGje6Ne1PRAshDLk8J4gyK6X0
Deemr7YuSXnMUs2HlbO7Mdis6vp9mlJdWqZGjGNub4QFgOD9sNaFBsclYRsCJ+Fh
`protect END_PROTECTED
