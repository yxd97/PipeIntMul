`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5LwTTzqyek7yP/Y3/YKiQDZRlEu4kQ4Xv9iRwPQA2+n/KMaDlDiUQ78Nd+qZX2j
wN9ED0J0Y5B5cMtDxrYdjkmgj1qe7x1ESZn2yBB/Rug8x+xkmQu8GpjIOu9WkKva
s3w5244QBo67JJkZjEfESUfYh/TPUkzvWcjRldBvFJq24sv/ZpHLj9gXVfhfvhB9
FRHNi+qNHItwJMDEC4SWxi+gFiyjUtiSeWYf9tz2N7Q3K8Kz+z1Ap7AwD7oF1JJX
iis6PYnf3JUajZs60V3335FEWoDrkFgp/dZ9Bbkwr3pT0iJUWPY31Rt3Xizc1dwR
GBgR3ijMytgaJRXmGvS4y6dlp39aUXyJQGYsoOp4yj4mPzsFbNG23M9Oyu7B1QQJ
`protect END_PROTECTED
