`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+eyAavJ7QMLiUUUduCaXsw5BL/F7hoRC+oppYAY7zikWjIwhq5DqS514fwEauixU
5bGCsMv30HuH0EpK99lHlgwT1BCnFn/B2qRSRwESlrJOgPl2LMdUsUyQoLWJdEMH
sVv3unYKZdAbMg7HubjyYTbbXiq165q77BRpFSJ+RdsQ50KOlX63QYQBDTgn4wpY
Wuowatu8FU6WyWNh4n573wC9SQDlc6q0OqWWyUs1/wkpd0CUMeY00FUnfw09v0md
WFjJIAwzzaZONyFv6XOeuQOrfKaNKghE0kryUSbh5OBw4DZYA+JHT/zhKFYD1QkE
Psg8aVEH76IB0UrXyeMHcv9TYyH2vBCEawdWWhoUt0aFmY9bvMncg9a6yBcSa8u4
1hVTyKO5zV7coqHZsEixTDY8Hwz7eGOCQlM+gR2HKbN+p6d7eH7xIIrjlg4n7s3j
0xhdBsodNBaSnPudoMWOxf2NRmEJAPwFGOfhQFLsCTgd6azPM/+Uxpa0lU6g+64C
8JsMK19o3cz2ZV5E0Z1GjiOruQc91oDQaoAUjmfPt1pW3dTQQNZOMZejlRthUVRU
2izU+AXhPIT9OZXH3Jc+Rw4QaeQVSXpiYsQdJcmznQUaMyZlQ+nioEYoUVOFcbhB
+JMRPWN+zzOEVsLV5RmU+Q==
`protect END_PROTECTED
