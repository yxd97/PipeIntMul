`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S1QDKhwY2k3UHmoodMHrZQgwZKO7WD1P+gJCldSGo8SZnsCGDlN0bB1Yrfyo1iWy
X7AwUmDIq3zYcWHIO2U7J/MBKhQNvftdZyKXqEuf/XxC2LU9b4NHdbMdcV1+H+AR
OqTtItTfXN+2cDAISfEouNc+dXAD82GA2uBooXDhUCFzfC0gUyKqV4GSveufdO2C
xjPD66jLrpM0GGnpe6CZQScijr8h+UaN4eQkGDj8GVrIoMwkZFYueWAZlxls0UtK
sBdLxD7CmHBDXNjPhetQQNOvHjq2VGg9N1aVGbf9Mgs+nny5EuVP3El0SWH7I90l
iqapw+iVsN4gm3QY+F3rdCRID/oCuUg6IiOWnlL4aCoZdrhWlP0P9W3oHo5cF3Nz
HgHxtDyrSadxYMgG1AyU/b6qRNFeRE00EOO5LFNQg/1eCxJxrw5l6Qy4ydDPCHWH
z7k88uD7GBOdK9ZwaeQuCUZNOMMetHKfmrwfANYbUZvEIK5wjNJpHHjA6ryCzhN3
LEuSCj7H8p0Fb5LLizBLPA8Tx10G8hhd0e+urBDe04yGxV3W2B1YtsK8f93Bdbob
8S3B8RRunx0eGYFctIfOgkKpAXnfvX2UqNS9oJL765JM7VFV004gBRJb/rBT4cIb
vnJ3R2Anyy3VaIHaGwA03qCUuklBjaeaTE2WqoH4NLcwfeh4AnAa9jhS25KoDFIK
OeqQxpZZs+1kTAnRD3+htu3fL7dUwgocQRBgA/Ojc2bLlXZAhW4wHvy0B47EJ9uh
EJfrCtJKG00X0AOFRMYVZcEdKqYxhWPEwN+QxvexVznAA7sQgOhXc/0B67ilgbWV
HnNlKFmmM0/4YohcQE0T4OJ7b24MMx0BxXxGpU+k9Cl0Jn8ueEkEH0nw7h29LM4U
2sz8Pz382xUyh6qKixqgr17h5/skWNuHsMmkBEHWLNkEKTEI7wEgOLOA+Ka7o+Qv
ZQs2ER+3u9JLBkaH5vl+5SQRRYr1zF82oRhVnLy+EawF8Ki+MqgGU7hQquANQP/2
jQLlTplDUFBp5kkNofiBDNctaDnvWt9yzx9BqpLQmLz2k34EMQd887WHE312Qinp
iuUHB2Y0fR4FxBRPB75BgWRBXB57pxAqrJP5fdMd824Et2pVeLkyPYNR2WKdPs7m
If5+XT+daT7Plbcbg+Cjulp3FCQeOM0+aZdTk5ldbg5pDLiH8ICjfPqbA0iV0Wm9
EToBe0BIMmUsx1rKEYSmn0tkaUujvzH88+Z3Ag1Vbp66JDqkovA7/VXlOzCNfFlw
oOvYGEC8Ujf2xiYzgxDRGiH5z56tMzoLGu1LEP4OxxgFoDsth65tlHUpac0XF9yX
oJpqYYGflFe4iUNqZt0l4W6+mV1ebAL9IGOrDbM786Ou0xgXxuPaaNJzKANEceJ0
z4RsQSkxknjMmWKZuX8OYukx2CgywGPVkS2OuYTOCLbazM8XtSixnnup7U6tpPfX
uo0S5KH0ZdXA6OgtxW6SpgHTOmn8KG0MwBgN/1Z/XgL1qKAU+A4fn/O2yg4OuY0O
AxvWtP3NGdUKk/Oxvmn//BvVUXtV9adQoszymVvnJhjDe4jT5bppx3j5dVpft88V
Oft5BB1t0+BIiiSswLFK0tm0sdY/6JWCecqQ+WyqcaeK8WbqxlC6WCveuHEkPaGu
XYgDQrPCqOE4M9ge5u7uBZ1hNS46x1yaUehoR3Ba+cNtESUsSv5+zzZcv4FAQAYc
LHbhWlMHTh4yby/66sjObRQy9THLC9yHFBYdZjhm9qx5g8kvI4tJv1ihcE/w3iGZ
H7UrdcNMvvrogLzoNqavXAq4+R+BuPeZl5bL2bQ6QWDkMJwhrHJdEl1wLB+oeOGn
LLmJ3NpoXLGBJCi7yEiqkSn41LYmSGsPgPS+qde0TiH7/bOr7OKtaBruQeW3ziDQ
r64T4UnKiOG4gjfbPJzyPObOikKktA5mvcDQFWBpuXhyv0TD5wc403a4LlvFcyhX
1mUzWxrN/M2gTSwr7K1JLcD+00umdcfeaXobMd0pcD9YiC1QNb/Mp36l7pNe34wZ
CwINTbvTOFlD0Xsta7Fe/kFoD5CUy0BviVgB0b1Fy4wMSJcSyrZWH46dhpux6l4y
1jlnK4JJcr8/rhtpRmgWJsygFIZpUBmvOHcVh+CI2IHbXAuRar73jmS1JRXr6+0N
WVZ+3lRfGOQLI5f4SmN4/SZ1s03XSjdaqSEVcIPvQl5KPtbQDImdT5bJaVmvCGe7
VuHrNPHopbm8n+3vKCAlLbBJbuVc4TbCV+TgGqjWxLZeHmR/YpJmP31oYQtLcR7Q
ibYf9dxHw0r4DTSBVowFfBeftFnSJE0WSLFgOb0CMdGfY3kGxv3rtmf4Jfwl3fpQ
WW1Bzrh/ugm5frAr8R4/pFR/dnO5GgjzPJDMjSePjekeFU/6kfQb3fXSEr7ERwxH
pLiEx5jxbfilrVZZCQvO3JqDm8XYg1XTnk1tJQG71gFZERcItK14TcOIkJULW0mL
G8hVEDHBEGtcULKq9ITWHIOZNqXV9znvPKHGVPuhIyDuWJj79mFVG/As7+diHibV
/VNCJ/nUp4f8p9FjcDWoRMzCQ16wpzQB06sKeAeOASmbtRV10LuNsC89Vo0SRE8v
yHdbAbP4imfWP2Nf/rilmH/i+rhciiW0O/ai5IffVtuAHJODqk+DrAoDREwPj9CZ
O72gtaxsPpfpwUjqID9xdodwAwnsGuHwiZmj9MjOPJbQ4Sj6R1/31wEm788sy8hK
PFnVvgiBcxbWX+ewhN5hTdHFV44ts7IQ9Fx1FRqjSMCVyixiGCyTJo4l03tGmUQz
MZmko5+ln1KlF1sg/U6voV/uT8fZ/i07Mb0RkBU8Wlz2RzzCFaNck6DzeHctGrbo
ba+yiNjqEcJP0mko7SQTracpHxtLduk9j9WnAVDOP9CZsm6lLcyYSZGetIL3UbHE
LOk7cgyrJkkJ7oPrG5a/wPa77cMfhp+o+/1jE8qcDzx4jLvVzFe00UTWH+WZ2YkP
MSxKRpVv2QXCsBn7dvYxOj2RlcZUYmMhD3RupYBW3qlFluuIzND0WllhXTzPKJqc
kpmd/60641SvrVdAiVOui6YhRh6mJR6a083bXoCRLB+dzEMC5stRPanDDIVkjt1a
1n3vbdoo1yQbAhA1mGPgeOXIXfXkTkfc/gVQYZvMPQoMy+ACu+erU3jeE1rjYz92
dsDhcE/MfyIH5zRXJzXlUP7Bl8L+hUhk4Zh4P5ZBZ+dEgVDiQddhp1/vLK4GOFqM
WF+IwBhn/7m/5M4VMLQgrIFvW6PSSBB2PFBueDq4VlLww0mNjCcaWteK6Rr1iGV4
Fu4fIPwXxEiVMoNDwsWKQR/Q9LEP+nvcBBPPU9DRoC4kv45Ce0aNnXsbaRO5vkRj
gFzYMDLs8hlQg6xwF7pT1UM3Daa46YR/fc5W1zzc5OjeViQVJhGBaujjE2qabkkk
GgE0uXx5omSAR3HE0QUBANXJlvSFweD1lLHpcK+5IOa1a1/MQToe2yYWXJPUe0bE
M8DCgm+kckIjZrZNCjn6dssg95MtNJP+n8ZGVA7y8L1yqWhjQxYRXOXYPhx9VkTX
ebUm+jAuJa47Pq0vYzFHaYvFmBnctJ9NXIiVIdWZDG690xFSzzqFEOqbhXlH0g5r
ztlBwSukCFtNYNfxXYn/4woPA9F7pCfhMkL9fTmEPU3anN6QP5ru7K93PRWyrcy9
EjuMfErCju6pOw4S0fStMwWOU1QDloLF/flL8QxSuWRpibcRmL6dmizlVvl0Clqp
pOX6hYbqUf3BLQxndtU4xa3HmF9e3DKuOg0ffizpMpBeM/Z3n2frQg2LvqHhDPdz
I8/QhACv5ToumTGh0ukEDc7LW49DaDQ+qponrbaPWXmm3OtCWUvMclGgBKr39AMZ
UbG34S7sUspleet6yW5JxC8e4WG4d37ge96mZXO6QVDhqHxdrvfA4voJbJCO15z8
9EyL0jfd9AqMLbm1AhlavZH00j7HsJGMXcaQbvc66ncu0HVT9g6WZHokECVEEksE
+qmLvAfxk57t9gfcdRNFtuqCD7WF5pbZa1bu4Ky9JPsBNRi1PZRw5+4x9Q0hd770
llU95j6Xp352Y3wqjLG3z3KMORblUb86TizV6nc3rOl7LhHugdNv3m2EEtd5nRSb
CFooq2nuwUmPLPgIou/RBi8IYxaPKmqBj17duD25BlfB1TyhEP/rMGJkdADQMgvH
hAY+UvxyRpvPbxR7TIWT+4SRziDZatanHyroflrvHDIBQkQH8ytG0kA74N7hY3qG
T6QTiXI+RUd/3GLTVwWHaKt70CCXTuLuPRBRiO6EwMQbDHDzLHWlH5uHFp65KOIg
K7CgMvx3PcC7/vdNvYzEmtxyzidrn1y/QtmdFK9k8rQzs3SPKdZ6OIxQjBE8fake
F84F72qZvtLEA2Hfr4o9H9YowuBzRnkMmUyiqZ4PiMBjilgudeJOLBTZjmkzQyZJ
Nu57sAzbk7FDQrcck4dyjxLs0tB8ZcUoUIzDy46PvdQyaazFRzMpSl3jFzZT+yF+
+2YT6b0VYmTUnEoDgExiW0S8YriiI6E3z1MNCi4o8bzTcLFFUnG7QKkqgcf223m5
2A0oy5UJ2ZfsC8A2TYDtz5FqofE0iTCgIRN6nXYF7ryuJuu00jEXZjQuP+ie53ra
ciPL1cygsnHiNtapaOr7/T1PSFdMJc799rh5FGDcyyItYpOhHkwS7ysY/fV5070p
JddF4wWMt+/qE5vpAcfv+o8+ER6v+hr3J7TdtzVi85BSfR5uyZ3MMw7VwwrCkvTI
Rl/QbACBtgIl5lCd+JW7n+qUOe6bcvSN1PbrHFP+aZ6unv41CS90QW5wbRHKafGn
U6vCdRfzzCR2D7uFgyT2UjjGDnu/kA7cSpkaCJtkrWB7QNeTsNxW3JjkmtDEeSgt
wj6uPsH+Dn6X14LPOaaYa9HBqKkcnrBR5pxZ5xr/QSsof9wRshNZh5OSmNbMmb8w
RF3esDdAExk7ZgHpIa2Q3pn9vMMo3NLjJguydakjY4vzj1vQXtXTaDS06jsFUCca
DD1zbJpKEdNipi065Fp3FdmdDQWlKZQU2L1+K0BubWeSeu4ugTTEDVv2QojiguZA
y5As7D1yfyW0FmLP2wyFMXqpMQATmb4dX60UY5suZYFdnmfULloc40aLNgLgtKzq
3nrz3VjCpGc3bilOy+m3ortXdoGZoE45D9xjGohGSUxVxcHXd/La4PIBJiqvp1zB
HHQvi1LpanFJaiSWO5TTRko8YwLJ7m8bcFlR34qB1UayCnnMfEWIeoYpJrZrExDU
PovIxVcPnpHL9q7EErFd3h9qF7SfMfYdonkEj21NRC5o/DjTfoNd4SojRwrJscSM
wY4uAW9Co1QgYTLJj18huWwZ1YdNgl/IYK/O6sGYKTc=
`protect END_PROTECTED
