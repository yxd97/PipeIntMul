`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rh+ZcYvzO3KPyi4n1DlEbLyLVjRCw4QcKMT/4bIwd6hCZBs23qK93OnrL4O7Ef+v
Oh7/+0lqn+GDrhpE13JbhDZG+mgt49+sGTMoZkecbfG9JqQKNIkvCtgn3X1FUeC6
kyUeaD2mG77/L+67j3tr9dNXA3A3g9Epa3mW1r8bQ1SgmgbaBHHzPcZq2saufm2I
dDk9B4nPULL5dBYCJmAzaFue8c4yJef9MaKIZVmuTo/J3JIfRPUfX9Mgi+rYuQlE
19HBOR4043TxpD4eC9NBbEPzoLz01TW0vZhepi/EfX4=
`protect END_PROTECTED
