`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DqI73TLRUKKQQ1dbiW+DZunA1P/Mi/AhjuMa+AdmUhxU+bQ6nNMhSlolX902zdvq
2NkvM+8LtuedMmqsihGamaR+g9/0VDX4q/aWnL+yQCaBpolBjETfFUt5z/SzSX08
FfseYeKFIsZfr5gUscFA+Cb6vc50PvUqKV93gtjmR4F+hMxUvVnvJnJRkVcTz1JY
ovzexhOrxi2FYnFk7BT62zx/zgbYarz1tMGES7H7Rg7dQRrG1bn8dbfihloDEm0K
9qSh7JWYHDQn+k8jvyB3ssApbxK3qm6hEcPu2lS8f7YGyLu6/urxMRA7L+LuoLmF
kc+oTSEet9uy6MEv+deKSlwisw71SF7pygsAfyZx9aavh8yiwGRY3cdq7iJ507fD
hR+0VMMpg64AsiWuyyqbxupKhFtWzzTMA7ShsDA6JQ/GcV4CzQvzHVGqxDt/EREX
XzEy2k71dE8OQqwjylKKcvsXTIWiNfWzelJGDgYx7rp7myuxbLrM+5fG0zOfv9Sb
9tzmMn5sCnm4AbF6+ELco0NCiiqIOYA6N4pWCpCiSKQfDrfoEr8I/hjzTYZk0v4+
D573+64QrJ9YXHxgekEX17RpEGuGMe2xrR2l9NAHn2LW5cBs+tXztU0vPPEVXgoS
8B8+AXcsTzlHL+XQF5WQENzVe8I6jzJRE9sQnZ7DEuE=
`protect END_PROTECTED
