`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+xwbU7qyQmHhPrRRNNYLf3ycIZ012HwJD4TN4PU9FEKVIr8088kQqJyS/Iy3aXE2
tIxERXEETgTi/mUS2kozQWfwmnFvEhnQqBxy7XY2IvfTCOYdDbXrNmdnJv9soKvp
JKDobRXvhlrPTsFUvzwIzxwGG/VSCqb/lYxrgy5bhZ0iyJcns/q+YpLjhggoC2S0
+raG6vgPd2lhdz9CoDudBMFkcUJ0s6GrrRSrXSeECiVkU19X5YBIB3WNQWhxwglk
Ejht7LOFCqFd3ARhdm9Jmyce4U5W+w4SvJUJ9pQ2/Aw9gIbFjD4r+5Sfwtn8reTm
lAMCQFnarYzD5B0ncKe+l+yrHObWmWrJAmIX7M6uLhnyw/0hADWuhqPe4421yCEu
fGeySQR5KYQCOuwD5dK4XLcFlgh93to4uMW4zv85Gqi21z5+wQ22hH6fSXZuTXRQ
LbBX8SiCEEha1LM7e32PWZoEVgYGRtoTm0Y0AYzm7APYo1PAA4gTGxCHr2ooQlB9
whZMUdU1sWxLygwvSnByZj44U0+SoC77JfEfXe6rmJC9N2MOAhQYeGPi3kPrWGbJ
3uT0Hq3uW/Gq9mEbf1qaVeLy8LZTedIOnIa8WULS/GCFo7y1OPOptDfuZ8Rmaq6M
URjmYd5V9Q4Iss5PmU2Gxa/ActDaRyZqlfnT6ymXAzE=
`protect END_PROTECTED
