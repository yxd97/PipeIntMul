`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DPfQYPJrH9ifFOKp3d2kJQtBNT8dpDf5ighB/bPXxfEgIRnSoSgzYq4ar/kLQdZq
dP6TVVPgpsh16cWJwtHIRTN8p+jFB7uCRpumqNojqrViHW3UArmjwKkmv5oigAWg
ZyntU2x3h4NC108GggJUkIzdZfaFImFme88MXLtylUVyEt+G5kAsx9IUq/kys5/F
x3BOqQxcdTi5g4BPxZdrmyqK48uGsT/fq9A3QT7ATR3tE7Kd1D7CVaHfiHOaDMsD
7VzADVTpuZYqnUxpUUA5TQHkYIf+AH7jtk6jnlOD7gbRWOHrhH9P/XD1m13RtCXk
XE8HYAvbXbdjJB558NPlz40bjyhZ3FmvEX6Kf/6oVMHS3J9R8eisFn19ZOImPpI4
/Ov3apHMaJx1GGZmQNuPtp6KDr8lvLFcTLod3cJIVGYI0ENAe/6XoZexT1ZMUR83
vlaql2tOQSIFqIBDmWgE5ZfJMkO6hYvmc+ZUJ98veJJkHJqJ9Xu0Y1OrBFugqasA
`protect END_PROTECTED
