`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PuHZ+/YCDlBdLRP+xIz6g/48nc7eDk864KYmuYcO7NPhB7af2jmM2V4Ej8YsyYHm
QkKEqU1OMFDgZd9W4TSUoYOFiGYdVQAh6jbfYX75Ya/8/l205THeArbR37jRBydA
LUqClWBO4rkx9ebLOAWI1Uv2tcfe4fPObh8AGPKaPiIMZpMNHiw4w9wicZOt6rbf
X+/agQSzauHGhFKUfvpivFVgfZG/jZhf59Mb5hrCjsSx/qJlgM2Fkx4n/dY6WH+v
wK4CvGdzL/smQsrin9cLVAkskQUR6t4tMqwITxTfL3ihbvVWAEyDKf0trZadPtl8
Hkdb5nju4vaeGXwGaFn8Po+33RsjzG1emcOaIplR6HknQ+hmzW78qnaCXXd+urjD
glmEalvRc1q1+FLhJm64If5PKuVFiP8ITuddmDVFDxTkRUzrT9qAX01cbGYMMgnM
s09to0gQISi3LvufqcHAo/SEKFX9qz2vYgHG+fx0k6319i9Xz++v6jW7nA2FlcZa
Z+oBfjkfYUZhm+v0IjzP3dZ/w0czOdVqajX7Yc47T/tOrbGV2/beHkXOd4prKNj5
jgh/mcxv6VkLOxDYNk3X7RS9DXHbkzlPC/6AOloYqiQ=
`protect END_PROTECTED
