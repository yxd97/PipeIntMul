`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yv/SZO4YBv8KcuZh4X/D8/2qyyt4gV2CMb9J3vWWbcCck4qUb35FyFvjNXAHnKFG
mW1yqnPO/F0vRT6rRgN4AvyVMRQx/eLZkJrTO5Mjz9MFeaPakZKoBEnJGyPtPXqT
/+5EgcZbW21ORIUG2pyCxXZk1JlX8Dkn0d2/vos2dqCK1d2+vA3atT3cJyh7JWVx
QpJpzIzRF1W9aXP9I/Fm+PnxvI2PGx8VHijDmku+obR7NwJeQZgNg9o6N1lUWraU
325Kptqm4YKeo3ihGRv3JDDzAQPTxfyJHRPj1E/t9KYxbnZOppKirCRTPrWiZMzJ
xFLC2L+kaYo26Gsb4e33a9eJiUJknH/3OKFdsp30vYPhBmwCWldJZeqWpQjxcIg8
1jeYQgHO9oApwP1O4wzCEShFndZw4DFXoYYSNghoPFI=
`protect END_PROTECTED
