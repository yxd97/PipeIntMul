`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NNO7uhmTSwwC7KVMuCj6ARw5kOih64WwBlJqsgZW9X4vz32TaWL83GRcLuHhDyBU
bcKBSz6X01Ccs1W4r/L6Pu4S24I8lYCZUsPSao3sK+kXGrKW3nPDAtoakHk1vvlB
m18ZmpU9pLSRFB7jCPWOLJtK7FsxeE+W3S0RTcEpMXN611/Ey9EOJ5lrXLGkcXpe
Ufu5H6lSKUTu0c4s72zIQbcKB902NdYEpeumrXRaIyz/tdxVk80KauRi93R0YObT
QJGxq1L7PHuQE7Bw7HBVz2HUAVKSlKioQDQ6Nb3XHUAW1d6M54LTNe+v5mzvDuK7
1XEbBZJ1QpJ8DXEwlUfcj40OCOKxqpF0fr7vPg9Ih9+/mXJPPRrsvanH30ekfots
nMsiZYCmJ5qY4ClSjUd/l39W9CqooeszRmNVY9unvNPMvT8SSibmP8GyaY9ACJj7
8RM3MIaeXeOtxD61+T0p4Im+IsNnGmhojL1pLlrQ+QSFdC0dRvcun86C5c2BAeXv
hBoVH1zzom+eV2Uf5RU7OA==
`protect END_PROTECTED
