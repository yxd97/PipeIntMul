`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0+4g+oSlx29Lprx+Igv2MEiztSB24jMhgkwwf93Sh67NtAVbbaNJJ/pKcD7bhWqF
HjSdVf1LGGW9v0Yx7M7VgvcuQ6R4abnKZlXFvfAftEu8GQdQcaYOHI+ZAYavDHV2
rSqsUNf5E0JtDgoPHrzA7731PZkZAEF92EfPJdUyLy7lv7LtylxvXRJKhL+L7jLc
gF+alGs+jykbldjS5aDG2PJOtJNjofhvT/lcBCjzktfkEOkH30g1avFD/WkjNq5t
aVcBm/vxNUvnp46M+82wswbNOkEdjWFKIAXbr7Dy2+h/2jEWkcBbIrgMbDMs5UMw
XGQ5W2NJd5va29BNFeel6OJMx0n7ascrCFSAAt/pR+t3FlEKqrdhOmkcWFbtWLzf
HamVRydUAm4SzKyFn5t/vtcZpfNdc2KW6BJyHprn0Uzl63fQeecHXlT9QTbnfa00
J1t0jlj+zUZsnKt1qxfEY6WhcK+SjnfPyd82fdNw+FKu5h9S3GdJ/u5HJpco83sD
hCsQ8i0nBA+15fwcFhBHMrWntu6Wzk7QyYikd8j5izFOZtfVjsPnJ43KvlZ1vGIW
4EsLxyZzaoS94nNjX7TffRUYgx2wPSg/UU6dF8uSbLaIscsPCauDFXRZp26sYeLb
wn/97MjSq1ZvBMycX/sK7xU38lXnLkCjTviMjPAJi3bEeyTpL7Y9mQEwg48YDHw9
Con0uTRUAMOkvAti8W59stQ/dMnXvkIxgWiJhLxNbJksrRH/sZPPab9nkuuIkvQY
KCW3jOzob//qCnjcq6nZhJB0blfqOgJdt7BndLMTuz4WfPhbx8zFb/XzkTQD8/Rb
YiTDQNvHX0PenE9h7aFg9g11DlEIoUqn+aOnx1Uei7WzYnwmuV4nvPDdzj+AUKxK
7bzpbMs02CdYmE3gvzzh7tiaQL1f8oQaSPkizTgjLRswO0NZqb8Q1463bKI3RHP9
oSj07kWdwxgWwx9gDno1+VA+au2dKep0IYZvkXGypFRpbVXigKD6cY1Snt/76wmg
ygIinsvPZQwJcNSaa51bBkW8xvzMm7bfHPc04mNTQZQgX5Z34nEC81IoDoRjJkdS
CYKeYdMuZp/AGOkJsGaugzxJWTnIqOLWZHQMp6jAhUiUwZq4sGlmk3lrlpTE4I7a
EMeLhIUvgjfNU83QAd6JlD43ZAW7m3pyweJz60zjSj9yIvvsEJ6Qlu78/EnBtVcO
2YHtiaKrMj9nhk4BbDItU3cS+0qUNXfoeWXBOckdZzg9KCXDJRs9UM13Eup1fp2i
Tm95TAvYUwST6kXWXw+1RjHNSQ3xZLsOjrDEbJUBnBoVrxPAdTsHFOB8XJlDMERE
XY3xd6GQs63Bj+hRDGnr9Qwn+ZlR00UZ0l2BHrKdEJPEnB3Gwn8kF0Zs8LKpXZlN
u8EAJKYdmiTNkw2gX/I/TRxoFhfN0AN5i4t3y4fyHWwfpi/1v4NrAwXIVz09aZJb
xa77HTEuUQ8+tIOiq096m9fpPQBCzxjgQThos6wKzfrYF5y2tlXZdeDjk7LYEKCI
ZIB2EYk5c3/jVARBB1n269IWr7tnL7kvc9AwyZ+MXeLw61C24ouK4ylUATBj9KOj
6hbIUQUYObWM6Im6WZG0gpitkHZaT15rztJzEotxLP2cPo5l9jcSWSuod9+ZD+XC
Vq4kvFuTV9GKSI1ODo/eTvlStlUzQLfS26lg+S7LV0cxrmp/thqqHXKkN0dRZZ06
`protect END_PROTECTED
