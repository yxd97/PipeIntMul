`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/FTDAnX8jMiP8edb7xJBSnD2kTuEVm9gdIJ/jekwitRwx3005dD/0+1rDwC4Vp4A
zv5qKtYy7koUXHSWrBRC5UJ4c89GHXVmQVEXlS+OeSS3ygRK9IL2NXQrx7Tu+64k
9/3Ev6AE1K1J6MdQLSwBgsbJYKDCGpb/XS0uk7tIFIEtLC1YPwrbSZ7SqOumjd69
KDA+wKBf+q6WgpWvt1ttavxK1n2KhGZQdtDXExXTO1zfcYHHYCJ2Sx4op7pDQ/4l
BVhTmisb00Fhkip+YK70GARQBZ7M2hTvb49qdtSz/4rwgSj7/BtU65AZJcT+BJT5
hg8vKsz4DaGRP4P17L5uK0PzEjodz0QxErkuVOOubM0EsQyKr3ShSGfHYWiAYHzx
Iuoh/Tku/vO66L8i/5/MdWUG4wq8BFXsWtR2uSxzLjdbNyBYuIS9S6+L3PzEMHd2
`protect END_PROTECTED
