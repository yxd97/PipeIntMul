`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IEYt3KkNV+Ppr6cIVbJyVr3JhDT+IRTdZV4VnJ08sMZU/tJS2/CtioJo1caSUka
V4wofJ+1kWUUWXCROGjYLcYl48FUXReIQfL5C+t3OOawF1wg75O7WxbRVZRiY5zG
CQI7Cqyp8R3dvuIh9/gpDdKViLT2tHNxBmuICYDKGHootYukTdITbgRm9eQ9ZtaT
gGnj+Oh8JA7fwqXhgXt7oWUqfF0jcpvKOnvdj42SD0lxWAoKheiEx8jMUVGpngME
a6SdIqrvVuxx75IfY+gssfcH1mo9PhpVSl7RRa7WHYNzg1O+MMQJkfIccqGSSt7m
0s5a8Y9aax5FtCb0ZViSvtSN2RMGLPpabKiHymNHgiULcVtzJfA3/Mw3g9x2bv5R
sAPfBKRiKwcRb6gnokkUoqfUPFhos5j++ZqVefzdUClrDlPB7Q9EBVA78Ms6ATdK
4f1dvfFyLe66wrTamsU8tMYM3W/wxZvyfeZcqP6asuGnEE6B8dyTKzgUr0i1w5YN
wq2ZlcGfIk9plSicTMlt7GTELVb8wCzlA2YMR16z1ORsWXVzmnGBeQI4bjfFwWCO
Vidat0sWdVDshRc2/kPyjEogntR0q+L9IkAZ9Y/HIWiCyXOqgxoSBiFebykg1UuW
TP2/xogbHvxtikQur3YPOMzGH4vlDD5Wrzo1/s3GGApQB6bfnibnu6nbMZ5wcVgk
qpBo9qwbPRbvQ1T7xgarL6Yn0Z7oUaRMh0/T2P/bToI84snC6b+uJOZRvWkiJEro
L6LJgAq/sFlyLHzxY49iuAhExhdb33YP5moEsXrbivEdhG3Nz75+Fx9Q+VSiciYS
`protect END_PROTECTED
