`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lX8JjD9jtuK2EYvw76A6Z+59/aVbSjV6rLBzpppZfdFZCHcFcXgkjdJ167G90CWG
EDivauH/nM7m/WbImUxsTIVT/NKSL5nIjMNMlEqjnr8QKAsxgNsrYUYOALQdi//e
iuL03U5UETewX94xKIq7yMXz4q+jToqK2B+JdEuVGJ9NFR4h2nfPOByWxgrMIRNQ
s/WXo0UAsXL0dqe2vG2gQgDAJa+4ObGzCOsRVthJhL3HbqWu3mpF8IcZ/AhmVflZ
E4F3k5oDlx36+VXN9p05X/tAmhigSeJjuCAJNrDxO3d63JgkZ3x5JFdDfL9u7o69
Q31AYVav+f8apJt1lY/AUmtbkeYYTjT8YPkKRoK0U3qKy/gbMMw1LsJRub85HzjO
kyLFqXv3R7ujWgqqHutAnfGM/bRm7WLgi/rYkSQB7yMog/VflSRpGmdm64dJnb5P
+1cQe21qflXS2U1JO1PMWw==
`protect END_PROTECTED
