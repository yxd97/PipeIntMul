`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tLu8FMDSJwUpkdyp19elThz8jDQTn/Ry3ZjlycZu7D/sNEaUW807EU/f8guxx0fM
Zi2wCI4dsGsn4AzxzCExPa7/CuJef9iszOdAPcet3LmbuYAK9t4BEveRNIstfLxI
j3o0E1hPrFxLlEUVkJdVqqYJKj3cHyHGA+wHUjrkHzIeBfc5EKYxu2OdGYsSg5E2
v5Vcj9qAsTrdJnqyJ7HfoQVvz+xi/r/xP+2Pqe184F2irz/m/zT+Hg+Mp1x6itdS
CIs8fGvwd1919ADtq2PK/uK5sR2Eiwfs5p+hvevbkI1rNc+HaUq5hlnq5+oAZLcQ
9JdXaw3UYiITIM0B235B4a0cD1isJBvue7L29wgPMUm385aDZN1zV3Nogv+IzmxD
UtiIHRJq1EAEtR1iXRPe9oQgSseZ766wedLKOj+pJ+f9Ie9v++GzM6JOn42q1AJj
lCd9b2SF8FJL4ozw95YDcx94ASw8ZNn4GXWMuKqJ6/3139hzHHS2HXlca+7VrKT0
`protect END_PROTECTED
