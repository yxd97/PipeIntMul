`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mFZZyAdmbj5u9vlZXvcwjJ6lgvSWEkYJKCBhGyCdEmMQbrWCEmNUSuurx+IbrH4i
YhdnnqZsAyjgKA3qgwM4lpKlS+mmRT0+3Zf2+1es+lf5mHm2+tNcd0UlWnksGSBO
kA4rAqa/sB1jpDDqzfzosZa+NVQjFkKtT3rKS87lynnI8Ir6mwkeO+3sSPgNv7+n
wkPndyGMb7Cg6wncDVE90L3hyfEYX3v5ncpYKlizQM8qPyzEe27zRdZi1WrO26vg
zW9NFSaJXsGKb8yYd2rBRhDI4zrz3KoyAgqXVfX/OoIbVodz+gXUcfpzHy8gJmzm
ccyYQyNTma5v3/qT7bcd+h1JVIGzjaEaz1AJkgFFP20Vqm4aTxFEBQKVPUpLV46S
G0wL4ifz+sqiehCoUmy5yApldfKeDCDzSGqpSedzvycct4I48wLamiv1Qy8Su4pf
1z/KgKqzrGJwaktVf/ATtK7jpR3SgseaDQ2RPEgKzgAnRX+JYinC+elrH02aTvzp
`protect END_PROTECTED
