`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WqSJXxyNFTNZwCCgIBAHW71iXJTF/WtRKn54BwREsO57ANHtg1kZO/V3G+W9e3SY
lxeSjc6ebpPqjJWCIfQS1E0GgpIJSFtrTJwSlPnp0c7eg0wg6MOPaRRJf26n4otz
iVLNnJ3FzVloSVJQunmkTr778WFmTDESixF5I1oJ9knYkowRez15/HhTYzl0b8au
L3q26dZ/lgHqMP1Nx+5fZtNx9ZaOBpJRvsTga8TOCC5WCCGTkerBmoISgWISrOnW
ieZspV5HqSyqQh/ufgL3AbhtbyY54ZA9z0XHZSTXzD7xb30xqaQeU3IvMW05kKuY
UAZn4K4Hk7b7NQpiDQJ2maJLPEqSQDYWPVQJN7N5Sx5BK+SloXFigz/1tKPP/Dn1
rubPyNgrGpCnNGyn+oXyXeEv4Ag7QSi0VTvL+iCbP8yEc3IddWPN9XQ+q5zP0ibW
sMbFU4EmUzv/wKEzNujJFeAx9Dt6p95TWMGFCeHQ3/myMo8WhSQPLEQVL54efn4N
Lx3FZDlADH2IeJqEoNzAVxKp2J7tYo3vTeLdZIrcU0ZOpsqyHMu6R/DWJLpJAcJ2
VAK+HMCfypgxgTt0/w4vsbr76TXWPQwybgB3ZWUSjjzhk0Bq81Mr30B76yllVF8T
pLR7cajB9vzv7dTr3SUkZg==
`protect END_PROTECTED
