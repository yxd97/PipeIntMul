`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
67OsFlE8Ve/Bug1RNPRW3o8j7r/PMWJEn1wI2+KgH2DLkzjBxCylDeNp15Oq2m2/
0QlGOBkTlynaNGCCmA5DIPboJoDivCWTUHmQPmx0B7OlbbudelCv6IEHoQMI00qq
HHjsHhIrfmeJzAr+uWIoeFjb9Mg+mq3lMMyPoP2/XAuNwQP1BmGROD33NXrs3qpB
eee79cB+jtukik+64MHTmIEj+7j1c+Mo6bV9xJA3MYeUEVEfQ2HYMPpbzw/ZOB9R
p0CMviZ6CiQlIdHOxMfdMKGDiC3nyQOMw2Ym5YG/6jzTUE5krEupFbmjhUAUPrre
jhyuRJtiYv4HRkxvMf1FobImWV+nuKQdUulNRNbsVLZxbaFhpWICR1IFVEhLi4e7
iKjmz73a8ZltuRuPAM63Q6xbXf/1bIqmAe1UGDgpMMSVbfBsgJO1Iv+m2z9H4uWV
bTjZaDTOWLuLnsIvRvzGs8suibmilcmUsOGkNqjgspjZ8J7NF2q+g678fd1U7Nkm
SbvaL5ZpnYS/2Dnf1EzWFrvP5m9RM1LA2VYD0wPVcQ5Dzuvy1uX2Ly8EKq5Pmeu5
Tj+NR5rzs6p/xIdu9XqMjAwoncoqfsX3hcA9xZInQu94vrX/XSMOehx1cBAkYowN
i9qW1CE1wSF/5uDRGFUHxjr42CO8ABUMHaqTE7ALrc2LygrQMWzm7NnDQFfOg69S
WbwVOi/FzI5Xjh3APEROXDX2ik8l9rBDtLWo5F8Ng8Q5bZp0WFt8tdOnUSPLrMIe
HEUMah8cS/e4PGMcACA7/1uFga0bIhr825HmrJ1rvfNqImojkiBs2sebu+sWmp1B
yg+NpkUi1Vs/bsJZkgCJGd96k2TWD84Gq4Yp6DbqD++LqHx/VIQ5zppEj561wfB6
zkl03Qimi+Ul4GGBDdpQg8oTZyhEuaLzAlmLRBzzku7SHCFFZ9waxL/E25IX65Vj
`protect END_PROTECTED
