`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tqzBv5GwGlCoZQXrzrwiqzuEtq038NMXNiNxmUAF0IRdqRdPrNGaVC3bWpFpFbBX
jvUc00jLkdTEQU/I12DATcfv5pF+wXytU25rISGelT83vK1lv63gijiuyu4p4keG
mR1VBt0zmskdj8xJmR18ZPP3eUeE/5GQuO+ZqrJtGBwTjxw4PvX/IHHD0nKTtMBf
KERGG4NmZVkxNrnoCNbeYxdca1oo/9JK6gQTmePFO2PN4xXtsbmsuPDGh8CfqG6i
eZdC0KyiYBtpzxBgGxxOecXIMr7oPiVcu0OaTedKQ58tjZ1paKWTfApLX1ps+WzF
VZSDzvePcp47hDDmWdHg5k7Hx2G896RC6vn7LLfX2v59fUJ9lUdZlK7T+Q6TCKOP
IYXNidTa1g+G1nQpBGOFjmPcIHVNK/DxwcY0mj+Xu7oeXcw40OoGzgKe67CAtD1x
BSHaJw7aylReBqldt1EW+yVpPEzegLdO7B9zNkOUNi4=
`protect END_PROTECTED
