`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
017U6Xp3XdTC4RFjpgkGEIaiOpDlWYax6CTdpbDR49/2oQJpXn8sa2aSyLe2LaUw
hDZxRn4hcgJVcvLNMyPsmvCe6dghyLOZiPgu2lhnUEmRvA+RKTqLYYYVxsk/vhQL
l4nOAwc88z794o+3wFJYVTdEl0kpS1bmgTwgJ/NmPGEKSWXUX2Xd/rJK+gkzkHOX
bxdNkeawYogj8GroK4SrK0L4kVoT054VkCrCzom8s9WU0f+F2bq7szXElg4WhwUi
An0FThMFKpDHQ+k/eN+fGA==
`protect END_PROTECTED
