`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uiyicBj8vCA3PGdDjQy37k0vg4BdpMiynOtedODfZklLrk2Lvtv3tQxLeOrY9lJD
POj4V+0BjnvaD7WPB1JghTGHManRvpTqnOCN1ukgkyn9Rr4hJ01+hwtmLmDTnGOS
2DQccGW9CSTu0NF34heaSsAgqm5HcTSXVE3F12eICzHIhc1dg6c48yQlyuT7UvPP
skzyj7nqYEp8BqlL49K7dzwWprds9fFyk5uMvs4zWjyjbTTXl/wpB37+Ko1FfOri
ZTmOJW2Kovqnw+vmij7dT+o7WMJOQGkCna2NyVm9SgANFFigfPIgPmP2MZ1c3yRe
/NiL9w8TPlxBJRKiwWkE8foq/jy04ulkBxeHiv5MmZ+2A0Bm/C6NGLg5vnN8ag1Y
1ECM0hkoe6domBYooTBONg==
`protect END_PROTECTED
