`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K9lWX2TK4r9mClXuc/G26VJkJZbnvKTjp0NKAbyx7lD0F2YLEoBGmyZWm+41pEwZ
PgcWGfWVX5qvSbU82/iyD0awKRZsORNI/J22deFk3V7XJX644yZlovjc+6hxGj0b
pUY44Dand0w8r5TpSfAaZlK6FD/8IhdA6r0O7GfidFkT3PtRZPcystFics/QFbND
8uo6owv0mEkRpB3Wg8ToXz3iHv+lDUeDw+Z/ojjtMoye3dKQ+cz1iBnwIIH5QG1L
NR6RTs9XcQDrgkdzSc0H4sPRuCS5rYQJAb+7xxa5J/5Vr5JLeTeTTsKuU4Fc8UnV
SyBa3QPkzB4ahayHi7cwHSWjmads73TdU6RvSIjXEXpW1FZ+gDbmGXl5nnawA0gD
`protect END_PROTECTED
