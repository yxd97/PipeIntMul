`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UgznmsUZ9MwhBgodHP0PArYYUI+39qh2fTQ3KfSSaOh3RN5Ltm5YwXcCZ+/8+J/8
4M+E+h0Xj6ljtCLggkdLcXYRLRjY4EUTBQMJzeqjILtib/OUqXZYbaStqIerLc/b
F2PqbtT/wZBX81vgi2vOXFf6HE3yzhrttsFDAY57wZ3VbzEZpwyJA6TwJcFNw6In
C+qGAUrCeOYbUau2UbPq+HQiidQaYM2Woh3nFY9DEGEp0DshexLPo8hMmkaa/qQn
YTruie9xIaKqtZ8j7Ihq1VckY2F/x/CITNsCLxDKe9t/cFcgsKcd6lnZYgACo/Z9
AgjwbwrW1uPMbPpxCl99AksjwOx1EKdx43a2fzJrB0XmmdO6JIV7GQs2b5DEKDDw
SnQymY3DeHskdLuOxn3OQXlj2wDV+YYObi8JU8LZZXXprtROirFNdNl0hNZzjJrC
S5G8QZ4sweNJhEubAgR0oRPbpQV/zou1hz3RVprqRIF0M1d0z0mNgMRjWkz8mFzZ
gcTDYFHXJ7g6bva43VIOaGXKMLq8DtCAGSY6MagrOM8aAd3BW2PJE25Hp8Flz1R+
pUlseVr95QjAWeOrs7QcnJOUXw7bo9Aor9Z5DbXxR/m+Wb83I4aluO9NKQxlSt+v
ggXxOYakJuCOZ+QTCGxtEDIA5q5iBVnC7AXHEZm65mO0aDkTgzPGXUumTozy6Bv0
YH1xVGPrB0B19HIiDnOXGywS2z/ZYfWvcMup9jXi/fn2kLyq/3XTTl4yHRchU9fd
NutD93fn7/MOEJG5tT8/cCLm5xjRHal7OLdaze0VW7gcA20zQrQdm5k8/PwZ/MQO
uVy5btLRXwRLQjpSQvcdj02NbZPjjPx71vGx35OYAa2Hwd5HTSg6ly+YFa6ileXQ
um9/h47TqEQn53Gl34CmLRXeo46PVxyV3RSKiLR5CV7AsB8VwrNWtEEE0i2A82jN
2crWDjsl0cSdrm7KCVJzig==
`protect END_PROTECTED
