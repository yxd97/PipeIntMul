`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WPcNAqt2+9dX3HohF9h1B3a3wXWyevKx1D3YaDw6CJjAQKm9k6hH9dMne/N6zCD4
cSYwal4i+VNtXm1Rh5lsR1eUUXPTFnneMRA4lTBYwJA+8lKGjEge0qjUIblunAuy
TFi/+EXPkv/gYO/nAa2pAyixzJVM4sJxEL7sCz0A1kBZWeFKOdh+UizquwbB2WrO
rfsnh0q9+bvLQREAOkaKIYq+pj5sSiJFV4Akm4GD2m11VjV4F05VENI5jNtucimu
vP6Nbzr3fbUNjhd3wl2/IEiXYdZKOGEyzuHpcWQ4q4li7GFmd4acQfovej9g9AvB
8DtqZgcF+97KXt4D3YhNS4nZ56+hEd9CkP3/TLBu7B8HIgvPlBNqe9yrT7Js/5MI
2tI1LNYjTA9nnI7vRftK1j3P0ZIzY4F4M0jullOaAATgeoJce5y/8HqksOrr27d9
R66szGdEZkRIwOhX4pqyxd+Y2qsRraH1CJno57T6MIymGnQaoYrEZX18RuZh65RT
X5QwHMFQU0YBOaRqq0TzsElu7K98VMvBXYF20WXl4bvdBqxATDcLFK88Npv1Ii2M
mP3Mu4HVSTYpSb++sIgs9dH9hJKXkG+goSg9KLVMwqG50sq0VyhCuLvzrsz6FuCa
LLLkTwo5b3hFSzq66WGQgD9mH8i7s7KlaJAKZ3clQzY3pOsJcrwYsqcGvUpOCuNF
P+ZppgvT+Wv6n2492LoeIZU0K8N4tqTw3aN5TiqTmJfaAn6drSvoyAfrEq/hFzLY
3mHEjBEmq6YfM+LN/Tjfuqxh98e6tHimNIFkvGlgFkBLjjL0PoAJFxC/3DVoMfAX
vuw13yUbk0km2fmBuEaAjfRUEVMLbuLLRAw7exEbh2rGgn8Krq6RQMc1+5J9PgEM
V0GqIGhUnSnNo7SiKjXLLAh1s5LQzMz6cd8lN3M3QhY9AIqjvod2tzJZKmPpF0ee
RnXdDoByi7nA30gM9YLVsQ==
`protect END_PROTECTED
