`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SYhE9oLIpitJ/IU38QhFqo/F8spqHgNHYDdcwq1sEGlG9xulnCExmGQe7Xu+HvfH
jdzzOyW0VJ98TBCj5Ge+tXjAY0vpq7kpIjHvkFzmR7FCm/WdJcrRlC+RU2vOW2as
vc7EMfeU25f/FVpCgy+Ln6NVnWrj9QYpVBhKapSmodTB8Xv7QuExNZav1SFh0bGy
Kl9HRfm7DCdZTCRJF7yXvbxo4iwxeP3UwZeIZQu2sNiZccYe3dxNAsPmWA08i850
EJmCV0dd/nIkjHbWA7v0tNtaOwOeNqN+VriSZ0iK1RK9TXnEMBocdpsJcUNFVJrX
pl7834oY1qsxGMDd8cbeDrj+hLNWVYCTmqarS9be+8q+olEDyhgSFhpnfpjla54I
AEb7jt9SyzbIblZjQkPuGNYvVI6kR5/tI0HlcDX1geGThwTtjQqfimtY1bmP+fE8
LkQyook+NTGOmIPpik6dauQLOkhEsH0Vu4fKm4KfCEe9qwcEPLXehNwpsu6xIKNC
693PCNnctJZIGlGrHnWX0PvohRHpA2DfFFAqiL9LlQz6Ftfe2ppmkn70wCThnxpq
MBqspKBae7XaOpqeVwQ54nIlg6cF0Xi28zwEYuwJtrKpeIWth54divPueCFYP7Os
RkSar6ZyAFSNtph+d4WYXQ==
`protect END_PROTECTED
