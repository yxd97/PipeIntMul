`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ETKJufN+tqE1B40bZk22866AbuBklhwapnnpo2GuIs6AqfKmuiD7pBnvSOoOEJLS
errq0szzb/Q+H7BRQpqHNAYYeL9vzEXdpQpJX9jdOP1VBqgKIpscnptaFGmGCXDv
cWE6wsnj4J/cNtRViu0YOjPkKwjFexYVH0nSaPSuR5FvJBf5bK32LDRzqhLlaffy
aJFZaeJjwTST1eyVCJlgpMvIRtPgXuVloyhys8mUlJhidxqeZe3G+h0uc5Gv8b5o
NCOo3kICMILmoZazIZ1cAE3pEAozbu6OnQZL9vsqZCht//lIUBePbf1amMKugFas
PoK+HARxZ+ZxfK0yhOIMJQ==
`protect END_PROTECTED
