`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xu9kfmNRdGyet+B752mxKq8xchQTfcFI5EHSoM8oEp1ke8k/UccQndr+e69IhtfD
1+c3A72+4IztR619qw9CVA67D8nmUxJ0fb8rgS3Z+jwMPthqaipd8wp0RvwZRmjW
6LFT47fYb2F2RnLNSlFWZ2xf38lUV4ly3nKI0FsbjNUaWQIxGmBi6nH+aerKBWjj
BoaRorpAxkN7RM2XSsEjUK+10WLkE2eEh0P+xYYu2iWAi4ugGsCxrUpQRaawCDiw
Avox3gc/Y/y4lzyMkn//jVkhMV8XQzh2aaSO5g6W/kaTblYY6yCpGmHQiD8ahBg9
Ghgh7ps4loa6TM7j//VSiye7/Yccm3BvBrfFA43/M6DdeCgIa6pLw2ljYA4++UOY
eemmJUtZDgPcyyvSqsIvyb/cxhYfxU7goVHnc3Hd9id2QqzNTS76/fBxVVFNTu63
APWXHWG80pDFLMMEhT7uEUBM5GQI5dBljZH7DM5nlps9cTgQ0/vSvCm5/vgWqDUs
`protect END_PROTECTED
