`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wnkNIpRbJvoOjjSNl8bn1QJJLU5k2P5hiDPAWEgJe/5xsjRA8A1OD805meuyJ8u
opw8wQbHr3JD9WO7gGEKgDKVbXpuv6Ok/GvP3mrL/xA9B/oyID5eSOv9hiC/AMd+
u9AIPEtf6nacjp84DLMibg/Z0Q6CCCs98y0eXgAuri7wYH1EwB5i84IlKNXZTdL+
eAKZk1aMv/kQoQ/svU0MpUUSIbhMTEbiiAf0RwoIgj+e3zszuLcp8YbKNLIrCJng
HeYOfwGVjDHGQo28hI/lANlDasz3bzautYZea3IceaGZP2RVRUy8f4ompoM+/Cke
8PEVO4b/5mGkgQROMFKNLlIqwHMpE6iS9+m2x7CU1zmBrEoFriwvxJzZLCRpEJNT
J1QAqWLdBiakN+WLsnCc2q5MEn5kdKlQ5FPOTwvcq324qDyWlEK75zN/NiX1ik0w
GPRCRqwbKF7TmZ96D8m7VjgZ3MND9Yfe2fKjq03KQoi705WVW2+buVAm6/LPsYWR
0mn4zM2ojRnGJG0rIAgQYzVt/voq70qwmopmZWkrUwhHU8T065G5ckd0e+Ca0dKf
skIbPE8rS8tmMDzLMCZvkg+cUSl+yACU/nepXjJG1CmgEDAx7BycKCZdRprOzSeX
tMlNv6izdxcdxWgOL01Pv1pw08za8hDfzg6tXVpqZ3nLdbcuKmTry4JXYYZ+/xEm
OhVil5WSlT1hVSs/N+8vqifVkpGJSXiimwEZeUNM4TtkkL9A3xj5fKP2DHUDOgPU
47/KTC2bM9GPsbl+ActCByEruemV4V/gOf4lMmdsI7bRBd+PTMMHXMiUrhIBs83n
3+Zg8bbngynbDJYez3fFSplv74wOm3F7P+8XSWSP6TD1+hiPO9+3/G2lxpxjlbdO
9LLkEotlii4sm3Yqq9MtwBuB7QQD/lr/gTm720RrZF5BXA65/6fCplpAXHTg6Tbl
M9cmhycRocfES5HcAvwlLHGLp+R2K2I0bxvqGzcqD8DG+fAA07nDuMp6RKDOjSoD
raeDoa6ksx6BPjqm23i33pvXlaGXN2nQHfzEXZU3UfM=
`protect END_PROTECTED
