`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nlAjufibQnQzcX186I1jC3JCwzWbBJ/WnIz9E3rHlqwpXhET9h3QLWCqcD66bbM0
wmymBvyoKpVBUO0av6bub0SFadY9l3fCcUwcqiOEW5ZE5V3Ilw0K6AcKEDn2I/VX
bXj7RiV4hhzJUZTqf+f4DVdDbLFiS/FhYz06W5YZn/JK/aUFvHC1Ddsx1K58sS0C
rsXiZPD4Sw/9eVQWICelgN4BSeWKiWWq4Xi+FLVW103HD0lsoMtBrp/x1B1EBt/D
9EvfrjLfOSEvVBZ/ULn4rMu0Tkw1GbNAn1cVeMWnckxz3aHuDtRqZXHRAcq9D5La
xoydfIT4Vb9+0OPt4IriWb/7wwtc0ynJLAGFk1Dpz5VAON4JoNVC1eaffzXSuVRP
lPssyIarwGZpVy4rNWJbLwi0l3xQurrVbyhsFkPB103TMCgMBdTtO7qvxW5ixUIb
H7nEHRD1zJ9OoZb7YelHcwxc3rBVj97BzzpDTfgleUn2ZwoXmhyP65R3vkHKN6T4
uJZn5eReljEIcnTzxcimpDJTHEpOnTScPZv5c1CtAbya1U9TsSaPVp3KUs4ukZFC
wq+DTNRPlP7z1mV6+uUbTVkPQNeVAWUiT+fUQTu8Pk5mClyNZ43+NRSdrOceX+Xn
VMGb4Ss5bvEn9PuIowhgSkkxTLn+XMuQz6gERRkSlcL/L3qhKmHq7gVB7M25eLkV
`protect END_PROTECTED
