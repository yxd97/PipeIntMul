`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XfTDJH4a9g1RWn3G4WTxWbmMIOZds9cfEf30O4eWiUYk72bG6wz7GcREpInJs7Tv
kbsgp1XqkgrY4340bZw3bEALp43whLChgFjgyPI0YTBuc7Gr8TBqNKsTkTiaXNoc
h7tx4JrC7DtOREPid85s6/5+G1U34fIyEtBpfn/9yuhXiPDbUBdAPeSDG3DS2mJM
2RgIQLk+9/8Gf0EZiYCQqD57y60a4oxSCxc7nL9o31HopvB38iDONugEN82RKZOC
4JlCVMj1D4qh1+U8ZpTzKzjlE8X7tTvCUCE7Obdrf5DC5xiuOB8S69WtlJ4gUAB7
w6zFrG+CP+2KrUMMf5zmaZpQNiPIppBauxyLT/zOIl2aUgUs/8KZt2R9o7Ptjy/B
No5cK8oM7238p5Z86RgicKiLL9wD2SGMEp8wkCfo8xu06Poh1W5LEyzK7uqWBqVY
0I5nInfOV/T7YZmw0aDLGfI1t75W+rTTZTntZfcPAHJeRYVAVsmvVtQ7NQLYhQsQ
dA16z3JmoCSD9r3rEKI8MccwloA0fTGPipwZm2Ky96VGpgj2urcpCS9KJMElfvxT
ScBAM+4gTDpKaxjKk1IRcpHXtTyYEE8NpN1pjdH+Rc/PE27jv/IZM4Aa0mJjJ45D
htyb7LhZ5DbnBreXesmP9xWhwBxrnIyV2Zjz5QM7UCE=
`protect END_PROTECTED
