`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JIbBeUNyFJsXwYg1OIW8nGdXF75GZHWBwhrevhBFs7zWv0x+F6QTlkKXD+Z7HOV+
oeTyGYHqR5g5TTtow6qtpIn1Pd5I7YQLU9R7FT2uX3vWTo8UJYVAPDq4YAY6HS5u
sOnPT3LKO/nv9sr/ggohubASMRTcdIbsgDk2Gpv42If99FZD91lUMGoLBgzMZJl6
Oaw+2lp1m1dtkHgrxnQ4hxwelNjFHO7a0mpLWPJfIUd07z0xcuWjGdg3vWjuJ22i
TX4DEcfcKScBPCS7c3ghNSLietptS0k6li0aejz28yLqh40UAzSszrq6DJ2364yQ
ouTrPngf9XDeYmbhVHgj1Abi7KrSL2iHecTEeuh+Ynq9G9ubU/jx0aNAxY+w33pz
QIIAtQc6XECaM+Wp+B87ChyjURHJYVcREwbv64+ngn759wWazq/XDA8VZWxzi1dB
eD279kLJafQ7xE0rTdEIqgQgKRi5sWshoJ6uFzjLnLFzNVRC5LDfIlTe6AxZOWQG
Y267DRmasBXHQsXIDmh9bqwb8EJ4fIS8ZY1sC4xDac6Up0sVW8EVwSaC8Ooq69H8
X45vNM6zLJgXrskIGa2UO0iV8qUm+uaKl7r1+y7vAFfzmwvQkiMnaDqJ+uQo/SE7
eEobyoC0O4/4QR3NVoR8BSL5Eajhd7VGpzUHW0mqrJ8OQ3UCW9aG89P+YN3wlTaV
T+EzkilU5rI2uXUBcQQ99FWXJ7lDrth6NruntwnAXhdAv8xMKSGtACfxKW+J0p+Y
thapaJWyxVEDRNmQ67UF0HMGjuuBedLI2VcC4JxRjM6K/I/CyQSMd9m7LUX2xu6y
QCUZsyoUKJlkZ3odGn+rjcaHCHd3FuyJ1z4P2YPvxS5SDFkLoD/faq5mnVPbQPpR
v6AH/ROqLDXB3exxyCna7D6OnTntB0dYlc6IF63gHxZq0+yBLO8ROJvU96cYmKBl
U0MhZwgBQpJ5sEE5jY6l9vHreyLwfu83+MGxr6GC2HKEVaiHQDDvEm12dCOg3l0c
RKKJMWVIVOAZlW0SVyx0oPDkvlmlealqKdSUfxQPC8VB1g/yGzI8hvAkQ/HQN/oK
Unzz7MqaYmRFfPmQp35IbdqevFO39UPKV4gnOhlqVnwacpvYJNeY6P9OYFONV1IR
WEC/ZCEGkzOOo6qjs9hv2Boll6IftvdPJ6845matKudFIkYFzNAgLoWwhOPRZh7v
BpEhSLuGTYD25gCGMiDr/7EC3lyKlyrhMU9E0XB39FeLqqRYTpjdC20FeyJbqK2z
bWFZp8iEx5VmVW4PRv8kM13faSFOlVyRrjfNPiM0TOlBnbRBAM0teGIveMl4jzLc
JmEohMuJz2g/3hhQ3fl3MJhmIK//my71eselnNGeEdcDUKPawO+U2Eklt0M4qpBK
fQIPd6K+IiyHZtE/NTjx0VSNR6kX3MNI0Fw+8dX/4pGscos1QMOyr7pVf6YUuPfv
qAE72p3QGDM197Ql22wS0RBZga0b6upCK/2C521PeDoKTkoJZmCda7fMZ0gZ7nmB
ohWu/K6j+XFijyOgJ+Dko28cCZOHEk3VlU+pOYpeVAof8yyn+kAQ+F7MsaEoTmNC
0OMXPULoaBg3Na69D+t21eGRvHrTbol4wtubpUZhi58aYxfzlm03pVlPDMUqTeW+
QM7xuaM4A+I2qWJZ0GdN2UqCKu+uF/o2Dg1eSS4JrO3OWCo3Qxsin9xYMI1nHku8
tqbCjNjZAXoD94KXuMY/Hz1IjhEMp8D7HGujkchM5CXVaiGmO9/TtvSwNJ/N+8y5
XZXLPn/R1bmtexu0/sCgJ6tIvY4x6FPiLJX4XiMjlbOG8ubCfHMqBpbSKrPTQUgM
0g2FwSXGXITopUwEeEkn9cvHNps+uXxlmabXsj68EOLvfOeUm3yQ2BAJHA7tyRoK
/YH3Z5tBVCTb+j8zITE+2dVBlYfrB7URLjyO9phQHnO7bHoUw0Wwcvkr6/+SkpzS
+/goN9fV4wHnZSltlX5VhCTTzDLLiYUHxBogKtBy1Dj2lwAxiTAC6muacoWJ159I
ttMdH8L9J7UPC/wSpVCQpk/poSXCS916ur5OMy9rPkStmLrgLzwa6kuQkZP+9rir
X7mQI+1Qya+CXgxCXGgj7dn1gg369gKzy+rl8B6Z7QltqFn6jLyVWEkORNu7GBcw
zbg5Zn+IgNPU052DJKpjEKa4dV33PKfcAnkNB+r4bcmIGXPbe2zFXfk7irGQoeyR
IP0FNRyZ8PxcfoF30Ab27xNRUXIfSntkIeN9J9Lwa0xB1xx/dfBlfUM3IoGTxeOh
pmhmPyy1lcpLL9FUFJXlbBBExts4tQn04E52zAmmEKdEVue5pLnao2he8ExZ1jTg
V6nCJXBWq4O0qRB/Lf/uO9S1CPcIn7Iv5xB9/syZdG9isUQVcORylKJnBK+dM61y
FPCNHujO9VVmYG/tk2fBxoq8GSSmwMZzkaUG+k/rEWVv6mZLafJk50wJgh1iuTK9
NfgpPuTi3KYXuh/JHE8ph8NwckNgZ5dLGWDhczhjkkPQJC/aw/29H+pT04yy/P8e
Crgn0ut65OwtMSeK9k4ZwTLSH2Mj5GBhvfraWlIT4ZT8U1ZDQcFhHmzubTaHN3lp
aUTBv068RUNCLTJJ05lSNV++YnM/uDUYuRiaIgIl3MLoMbuB3wjv+n8RanmkErCB
ux1JRJhEJX8BjsKTNLY0mX8DbE6OlZVoGS3MirXDo1xAB5QsXq1ptcYteckMkCiE
pnv8X7aea3Ld3Y8+0CrE/ZO3mg1uUfxB49K6H/zeUHEicDuQlSe+YLUVbdV5F9vs
IqZlViJAQs82rUs/NOT13KlRASIarfM8tl24YyrSAoZymjv4LZVNxQ+IVdCRmyr9
HmAC2FZf2etsOoSEcdcgzZrg0iH69AhCPMr7+b3w3lOL3tONQUp5H2xxcDMy4uIz
NP4sWyKn2uWWBtvx+rK1RRmWbalDEtI1JCaMef3WejHdJPpsVroYZlf/Rhvhzk14
yUxg9xTkNpBWvTkeG8dzWdJvKuSSM2U5kr8bVj86yJaVHp4kXeDAYuvavbEeUG6C
hshXTRx4I5KsMxpG6eQe+GBAd5zoI0XSyoddpkwV3gPBWmnx3QFabQkKKDPADuwp
UZOflzwkYqcPCD8e5boH8jamV4PR8te2dE4SNCDzb2mbVMRQZAzDBRA8Vrj7VFTg
Mvr+Rkf0tdImZJQc6VbO6r+yCfIn8OmyHT9IYtRI07EcPzyU7v8Riqjyiv/SLZsG
sTxzhfmzNeFd9KH9hQYBKyTQKAgsMglsdbB82aeri51hQp63qIao8t1llvCKYNKh
yPXMFZoKYhrnhxy7W88v+BnKgMevtMR18xdSA0LSRhq+h+PTa7mijg9GykbGY2ns
y4gHdvX8dMANsPtYCfUUN+H0dcRK7K2K68jRU/u0hRpCGVroASUvpB1qFD4hKLCI
7xtWhoQfc0s1/IhaOBzsgDbjCIlelYFJ+oQQEX5R6QMj2h3iIQa9mKbaGtmFHMy/
AxcGxUT7p9oM5ObLwL0elH3lGYA49tUHxPpuv09onk/lYaj7jQnREUIbiZgYGSfj
lZNZuxfWMEYdspZP//Azs98p6RKjpdcTjQyGK3BpHTOlGMzMCorpAHh4LGaJHNxC
FakLSMUhvYXbi9RAe+UjRrooaAVkKMTGCRRsST1iyGoNsOsOcHro1gRhhVPqx8AM
GunFdFzZ3UkC0VlX4P7yTx4BB7oFFnioLC5bmSJl696DQyfnhIVd3ElG34f4u6Nr
WVXw3UcebyCHkne7IzxO/uiHMhgvxsmJRFOZ2/XAcDANZLEi1U8LYZRDCnvVvs8t
UGu/SDCq2wFsKcTPormSlhmElhZOXn9G5bquhVeITYPjANoSol2jhkPH/h4v5lgZ
xuwjwdjttobxGcxs0WSeDv6pyID1L3vUJaXnQRZZ1KmjuY+W3BuPb6Kau3/knmh+
LASM4PhUaGpwHadK9AvlLrlTXLTQvM7Qy0vEhIEZRqKysbtx5UyOJElFGlBYZ397
bB9P0A8ZwsIl4ANS9TRzEnW4+a5ikEfO5eqpNjKZAQqszpjS4rHd42zkBnL4zxKf
YzhOzFtjcceWFtYqaYvU9hQ3p/G0blACwXqnjDHE9qNFj9MpEbmfAo+51AtfF5R3
`protect END_PROTECTED
