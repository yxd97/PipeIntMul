`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RXPzBsnKl6k6YzMWYGONADV6fCkQx8o32czFuSfDc2kNOrs1BtlBvwBPirRx517n
mLU05ApLnfAkZ/fo6p9R4fAOpz+G8zCL+tLbDPBZVYiETlaMvGs026aTLSaVdEhd
1YVtS3CEhbqvK59U6OwQ/QFNlZtts/zaIUFz8xHMn9owK/cLTlbdJGCvwJt+4eng
qtMzPImIwlzAqPCPWr7x1As0QCaRBdmCTOnuzCrWJ/+DNkBD11phVIYq+km5hxSC
KJL5CregolBf+NS4YcSkWytnZyuPXlEHZpGjkrk5EqC5R4rQ6XTowG8eLgraJVNz
fGB05rUkJyNFQur4Ju3AqURpM/1cecqBgPjj8hgz12brwRwEbnRfj5Tv9ac7yh+H
tixl4bMnZC2yisGAvzRlCE4ruEd+ZAANM9u1elW7+vofma8FXHANNJQUNpzRHG7t
4GziKolMyVZGMQKABBVFvOOLZ40nl9tH1m4G3c/Yha5tCY5tSBTWQF94mB/Ysbw9
`protect END_PROTECTED
