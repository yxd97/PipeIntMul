`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZTLYW2G3wf9SZyOItof0b8QATxkP5/6k84Yt3qS/g770semr/UOqIdjDvZ2NYLWO
hmLeEwahQ9BQ8Jp5zWN84GXlLzyUiat7XzY3pattk3kgnfKgCiBJ5vSJA4YVR8I3
oODOnPfrFvOuHROcRKNNf00UOIbovMCWzs7xV2GxyRiEejBryokle4/n++OXE12Q
sKIQOVfNNgnOgfSFxUOEi9ea3RevHCbWlvFoDemXZt7n8xImv7+nTd/fHjEyiGu5
YhP+11CiX74uHJkeCZQPWSL9Y340k296Ilj+tNvO5Fwa3Yl1A6Tr4hXlikmjRcYz
xqA9E4j1UUJqv/9ns6hSRIcunqbvQG7IzQ13toycF2E8PHmMiIw0cxlLdzSW2bVX
QJ5yQXA1XGsNuNz0hSXp4Q==
`protect END_PROTECTED
