`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvoKFj143J4W4Vopqc2PjY0SNZy5qOAaxtjaknjQniZ3SXlfYAhqK1LkDAHxbIwd
ve2siA+6jOtdSCk1mYlvnwQCpi/RfvmDPenx2FCuzJrfN2WKuD+fh/BF+nIq51Mx
ZNq7DCnRaRYXWNUEbRDqtkHOGSqRDKEuRcJ3NOiYV3HrNRYYelS12yh+xMrHmfT+
eDnAY+KGy8r3ouZhKvnOVC/8cEDgvWHvkToaLw7ufeo+jtNuzScChtRfkUpKX3NI
7KF37HONvSvqDnWRnpu6JcJPJ4sDjHNCcdhr8pNPSJfhKO79H2J3H1TBil4iBlY5
Lli6PwaN7p0CZvuGLFUqlkWKYGzhdakrv7EUgCtZkExETTAul2Zm3+n7Rz9m+LBA
mIsqHTzjXQZI5vO/MX4dZFxV05U4W71aOehWBuLwLDSjttwuGam/EVoUUb+3THzw
Dx+R3zrg2aKDJukadYgj2j/QeDfF6CsfUAzCeEbkfnM++H2eAlxXe4zIZjUNC4Zk
Q00FDcpVNnfy/+UsNd0QNHcKxGzk/oOr7YxJ2odm7zf6vItx2HWZunHS4ELLg/9c
dYqcLa1jYuFEWYHjqWuUwoO/uQ8zjvGG3TgH4HJ4cdPnP3AzzA3nyMWY1fhRBUn1
3kR68/iI8VTTq5JNcVcFXXr0GxBAkAZdFOkHXMggwe9nBiwC5veqHa68VPx89cHC
`protect END_PROTECTED
