`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xuEH4mqC9GP/8r+JGdohpj92rjvEka4I7dBeXr5kB0HULvN0WgYh/kr6gHmJWMVi
DJSQn8eBpVbmAItidB+61VMpLeasSxqHO1bVR3R8ERGLisevTasSiEFZI8QL8+If
t86yIitnr7tmJP3lYMH8qir3S9jIyBOmfI2LwEfy9bKz7YS1Glud6Sp1NzgtRZnd
UFEq3keFs4g033GFNcYhmGy1kDOfknsG4hmEua5qcamZIcatjYepJMHVnC2n16L8
sgpEFtD+F+lBNaIHanK8mZs000ftrPJSmLWgseQL2+c=
`protect END_PROTECTED
