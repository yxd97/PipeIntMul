`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Gl/2MNFtcsHMteFJ2splo3HekpuFWZ7qLSvGTYogP95C6So3j6T2shOp+qKhGmPu
O5XArsJuauyLJoiDB0fk6FAwLc9dOxCnHAsOu09KTWe5hjOw5fcq9F7gXat6I8ih
sdSshNVPSUAkgGzahZrv2IJEzvmL6tz0qBl8sYKQWgBpqiNgHJf88bXWzVMuRgLM
hXp4DWyxdV1CP5wq8G8meyctqJLpyjnt5CE5CAWNffRQHlTsoBMQsBmqQNcHKiQB
a7XS0yF9NEmCbuVxBtNZtlJV2sDQODZ2285h6KzTWQZon7KR455wS202TPWNkC9F
lxkglBu1jIxLGe/AdrvK2QVerXUukX5EzKbZAuRLziP3BeRqYI7PTGu3bP0JV3Iv
4yD10gbbGG46ma4rewgjJavdXpxGeajIyPbvRGquGAXTKzWuDhnpgBCR9FT1V3GL
MeLfZZvGZRw264mvwdVLw5UgJj0xsd0ni17kzvJDykrPYb+zz7Y9Xcra96d1nFd+
`protect END_PROTECTED
