`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r5Y1WYt6n8UCPbMfz6aAmpageGXH2JBnr9Zptmi9r/L2QewiET3dE6OKg07u5XuJ
cg7pyXCNsoG2k4pqyp5LDUPGAQvTC4lFf8lHm0fhPTILO5JQWJ7eRHCzPMz073Jq
639QqccAh7oVfOv/L+T0krTSePEIYUn33rdNJmGJoXS80zYgsna1uAVaInFslYmb
3gdD5jDxyDPsaVrwePHHkkRwVCd1xWjmR+DXPeWlDFMALAtkJbEXqxd6ljDLQnmj
1yd1RIRSFqsZQrJxPyHjUf5DF+peVOY2j2fj2qMUQs5ou8zEzEG5CfaVzIJ0RhEx
cS764r3vb/X38Nc2enDDguxRqeSqZdKDf4VNHXrFV1a275e0OLMrjj/DP80qAZkw
yuJmkZR+EILZPL6S7+TcIwkFTdUruyP1seDTixlG2ozrrfNuC58qfrNW1Dii/WfJ
gKG2H75qRY+vbw9oRyvP7tDvDdf9CuAG3ZlDPwpemhTL3s4PG/CKRJX2ERRA2MkF
7eyOaoHlH7nETGGUbPv9x6kGjSYZtBThNIfkmGCHeEtqVic8+lMoFiwGZvoRLrRA
ofP6VqbzvxjeCgAln1G91vcUsPQdzE327LgPveUK+1ODvQoIIGTEWB9/5aZTUIpD
zEsH2NvDvd6eWFVIa+HVwPWlmypHMh+Wei+UEVRrRKXTTKUOYFpG/zEfDRwNKcfO
fqhrbGWCdz6YUp4BpW9MjtU1Gt0I0wEY/0W/KrOAw38Df+5G2UYAJGxQP2mkiU2s
vy76hkSJAN8j7HVzuXrCqVA6cVQa4FVJSyJJ+6o4E40NgoobWox49s9I0ilRbkHi
Gg4xRBFEfWKNMOT2cV6EBOAv7d4iBgIh6VkAduQUp9+XDegvv10Fsla6go3jpdc6
`protect END_PROTECTED
