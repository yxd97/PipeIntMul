`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ns2baLfM5AnLQm9F36y/+zCVQSUKiZVE88K8UmId4S43Srxn01B3ETZY6c/DBwBq
a1ezOZNQ83ZKaDu5+uvAPK5KcqnEvtfarjBCSXuqdkO5XLFRqYjerAf64MF+gk7X
dJtjFLEi/p8/cakYxVZSeUVaxshy0ZwdHpMJUV5xLExc5MEXXsAXSxhWyIcPbRWJ
h3RO1Qrwz+YZl2GIjnGchgYzCrpgM6FeoKU+xAcYHqU/VpWZt+re29em3aYW3yhR
pOm8+SRyxHa9DA7958KKVblkJ3SxrER7NPlquWlqHR7rFBlY8DkMwWj94mECbGec
38KbF4ItgzQZ0VnNWJn5d5xbuL1GlGRqDztSqQ+4VNcUAL31LeHkvxquT7XLOd5s
j/0bdhcpuQwfsfJqONHqsEHQgRWBDTLdy3dPMAqu4FFuzf9kyNc8yXgPpxSCh5bH
mmDinpWMYC3YAeLsvCicyswfmwalC6amUJsfmbZsIS4yW1NntJx5TpF5/QjXftwP
YSUVTQL7DI+c3iOG/hdKdFEgSXx7LyloxlwbHksJ6k/zb3s3BQNhfzEDUZhktwPz
jFLDzw79SJuRPubJcMUveyMcZgy+aMVxfhkm7v2AIqcdYrcJlQDiHqCkJXriMO1z
QfkBVxSZHZjjYN/MSqYMFWp/PCd4e7kbCYZM1FfT5ZR2Oyo5tkHYZEm1ePxfMiCo
s5bi3hDFWaFllc72/alHEThCJ+o4dP7dwaCNRElyGA3SzfmKryBJ3KqSw/iyNbHG
XI7NibjRa63dapqfWRz216CkSg8nrhfJfaFzO8ADNUEdhtSIdHVk2VX5RlS/XxX/
i7k1rmJCS7Uwj+qFhYToQEn/UTrbNFiZu6bCVPN7R/d4zx802q6QkAJ7aiOucppq
DLHF9529nYL76mzGQfap8H00ymF4CYOnu7n594uLRaBYEGo57seLBo0qgSP/iwZY
HHrKlyX0Zv19N5ypWvHgHeeWpbQqjDcPBpuxQQrEGk6T8eW0A/39ijpIijgFsfNW
xea0s/5EOu/TeVMH/3ZH0LYB9HA0E1PVYgBeHwVG+WvnQBgMflkL++Q79UuMcmKD
a9XTu8csJEtVxxMfZak0bZpeXn4w05qhNEZdMDDwxuS9j0hk50Jcw7PRXag35d8l
LbVFVkudIO4ygtQ0QlvhNk17ui9+HO7+E61wf7po6uRPv2Q9312J2rtT5gtfss/d
3t0p0XTE8r4X0a0XS2Vjh9wN8IVlXMw74E4IxFr0cFJIBjAQZqXkgW2czdlgId1f
/8dL1uEM/bKNjPDsBcDyQnPXqstkeEUKlHwFSk9jyvlUe1y0vNiVcnn6YFtTKo5O
7DUsZkrCCCQF8ZTe4aEI7/TYPsuE2OHXgQMFF2xSzitf43jGhAnda5tIX2qsYO+6
LBAvjCLOB6E9kwS+i6YUSNoaKbHkSgcZb9WH6xgEBjPYWu6nrcg/PlLeTfMl7zeC
Q/deiSB0rcMlZlXgCR2lt0Jr0wMo2KpjstYnwW+XNH0oLyiTVzNKPlDJaQBaXrSP
jz4WZaIfubY53wd2JpMWUxzykT7xFong6ruSs3+AOTie8CCwMzFND+oWpL2b32wc
Qy7lXuS3jhpkgk/sTzGzonf3HOxIPO3pTOshq5JfRaSuVHFbU67ARboxQNCFHzEQ
OczZ+906INB7oqKbN0Y3j4d2CLWz9tZVm9saNWh26jMXk96ruuNHjT7ApMUHDi9s
ABGvmKeWDZA3CcCENkw/vVRNNt8Cg93bY/Yg6KL68Nf+Uuuj5umGjSMgde1f/MZZ
NNZQF1NVExReXHMhh8TwFmNzzh9vU8zX5IZ4PvcMEl54bxGd1AeZuaoMGZQB/MEB
+QUYWAlDJY8DXyOJBMLAEEo4chvvNEluuYJby67OQkG99FWIPsR8v1stLwBoOtDK
Xt/LrqPn7ox2FCXwj0DfBM1otbH8NfZLdPQhWOe81FAsd/FX4ELs+DP3SARVIM+9
dKjZIly81Lk3fbe8ZC8dVT4olDkHoBRUxqnAgKBvFEl8N8UVyGZ/F4teikPa/A+r
oJnqy9KjtV2mZN4/yeCrxbdNXXGI6BJ8IwC19R3wvqv7lFMzSH/UaHJla3mVqclP
wn73K8Pf8cp21elzu+U9FiX+bsB+sFtGITFRWaqgitC/DKaUrW9ntI4RmFojoWFf
V8PeE6qpAuSQzSqB4REJhW17VZ8wwZf/No+1k4bIy+4XPrwNOUu0C+nsHsKCDtOE
2vS6hcFHeI6iQlA5lRorfnGwiACC8Kng9KCT0Qjd+LPUiP0w+fnRKQPG7oAJZEwo
17mRyS9gBn/Cr9JWJh4c+SYGOiHnHHT4x6OMtOVZh34nqHpNQjDPy5qeHiZ/U2rZ
t5r9SrkV7iPCJoUsqZihCd1AqVWM7iHygRKCcXPlC+7Wer2sCkT/g3S48RNROFNm
Pf0ScR4o4eCTlXPnb6ehGMKLa9+/UFPyoSONu8SuqQSW2hUpRPSOLVzWxcWF5UJO
uJcomkla8SwMxlYYpcz3ce+LInpRdQhg2YH3wzjJHq2o7jZnN4MXvxxRiBPcSF7l
1dAK5fI+f0o9T7b/UmQWUs8iDWKFmSxUUnqAqvOlldk+hT/t24dZKQEv+pzKd9s2
hi+rzTPS7lh80UCE2MJ+zgUa83sHOiybazOvCGUURuNIR7t4qOy2WKD/NOftLAaM
x8iCR6TKBDaIN0/iKajtE7ETaDGdbhn+YchkYDhBYj/49EEuyetzMGsMmL/EfJJq
GhRQdknQLGsTAu0CoTLFmnkNjHZZq6LQuVVcRC/0MtpYuvBGVRUPaZLSocGeL5Nd
0eMezfAt62AEDMrkpvtbqw6mVUG7/mPcSS/dxqzwUcdlZHS7BLTwohAa7NJKBYa0
j8EsWdF910XPVZjGry/d6pDdehaeZlStiOmGPfIYc5y3vMTCN6CuiaD7R5d3udsY
UYBjRPthEC9U5t3jVhgzSWLdHm6PtVcpcas+sVQmuMacbIYUGNFa/pUlyqN2tl1z
sva6iXDDGMlrBN6IkYx3LhCeFNGeozv3ovI3sRoZdGBh4aEnrQr9ikvK/rDkIHwH
360KFz5FMYaRe4N+fN4S0+T4zLdmhVGns7uS00DOxjEhEH/qzufw4/WnrSZTAYZx
BGxpEp5gkn9vaLOdKTY6+Tn/i9AuSk0r9QSlL4KTPHcEHECaureylP+e5qHhTYRf
ruGCuL7Krtg2la7Kldc7xw1S9vXaKL1jZHpMpSNR+UXCdITAFRAxSsWDH9CFE4UE
obGhoj3jCyTPg8R9GBVGbx4oCbwiEXyrBJA+hq+SyY+xTBpM8LvI3szb9tM0Tf3g
64kxaLFvZSLivS5P/7Kkf15J/WD75qWFWP1NCzi5w69xzBVXOrLq3xU/2ANvjOml
iN9VOTP9uspK4Z95v/29bFoeFGQ4tBIayNOUURUrRCVVc4iUIHcbBC7dtHb7SyXi
AncVzHc88E7/3Rgf01J3jQnNpiTwwQMxQcfu4H1ZpiKUvzCh4hXE95m1YJxrXlpm
M916jLavZ5+iSqpgr/6p0blpsErxftw4xuLRqXYf0i62P+fHlrBOiv3LI2wxw159
grbNQbv/TIEKld2ei0CxpNCp78hkllk6DWthEqf6TlZzGs4V2NGJIIl/0ZKs0Ekb
yyeYBV0Acw1P+5A21OmoByWfW5XMSrs6GDwa9L0cbb+GWrK75Sy81mr8MuhZC0DF
uSsI+wL5gFScTvCCl+Bg0osJlSmVlomATJcKcTZkT5TE015/W4wjeZA/kglbZ3ka
xHawiaFtRhYob/VsCimK2w3sVpmwl9VWady9hIjfZ4wsTkLgio5YdkgqytZVI/Ni
BlOsb3Qay/vIoK2ZUZ/RguW/4eifyXQjkNdf9fkbVuPGpDcCN1wMhNpBmsmgSGQQ
sb5VmH20ww3TQvWo75VDPmTS863PksqpvF7yx3b2a0Z1F3rMhZGQ7tF6/2mRuY1B
bTQx4eIkxtl7egSqQ3Lo2AlKd5Y6lvZOktbI3sQzaVL7Dw+OKRres1nuxCQABQLQ
4pPdSv4LD3hRWoLlM9e0IK4mMlUuut1xdPebNuquSWYOCs1Da3BzIlsI/UY692HF
kVICO26U4116BMvwp3bnVLszbVOe0xH4eVTge/9mvna5XQmDzFJyZ33JwWsC3le7
SdDTlMc1POQ67QzPMyrs67K4tIx+rLi8OterEObXOZnuVS8g+4xCyIBKOa2rehYO
0NBkS4wzUlFNz5wcqJkb7NZ7TiFwecaVHXp1+07Fmov95fyZdG4uV40celQ/HkdZ
hyKCzU+3hE2RUggc4src+sO5pHHTFAkiAaw2LMlBtxJFYim1kyQ/ill/yZa3uWKk
uxVnkoE6QOxi+Yt93nhTpPT56neIZMsC6Fn4GSxTX7g5tmMX0uUKmn0cOQ9+XHm0
xMz9c3beAGQu8ihBmdNXiPQ2T8IdfZMKMYTAQEx9jGshwV3VjB61tppwg0X/7kuZ
GMZdurTyXMHifNl3kQvHamFLybBtucCjubk4zyADyrKjYu0SVXj2yyAEkR+RrknU
krfFIn3a1exqZiCwA4OeZNbldscfSzDeE9+2CifHAcLehc4aB/Q9F8w/RMLQGZnM
uoKvKXIixFRUOei7OmcDZu94BRqtGu2qVxf3SIsWwGmYb9pLCEqmKB9XMG+3kmkz
O+wizsXMqTAksf/Xaa2IdJ0ZXN7fwc5X2t5+0lOuqpO6iW7DY/CTR5nDnO6PzSJn
RhLWXy6i1UHWv2J+b9QJrFHFOrkMQirYELb4E6jYLs6Dtl+V+Us+nsWCM6O2JGlG
V+lM6OKdZ8dG2Bks7bQi0u25OyeGzr5Z36dfta5NmMq4uEeVHQy+SEUDtJEBEmB1
84rtoWpP0zloGyGO+pYLCWwXAL/V+gHir9bysUywIr8I9YFZNu4Hh8/rZxpfTEoR
dbk3hJwGt3KobbSR4d0XobfeEJnMKit6ADgeIuRiKLX1LtqaSuuGHRidccwj2+Y5
ihcgMvlrTB7uqOnajXkW771RuqcrQclZ0eMCpAZrgyWDyhJyOGfYilbKP4GwjWlx
ZMRX2GN07dihn90ln6AsC+0kpSg7a8WlvAlWHLDG6+jwj01Wqizdt5qqtxamPDI8
ITylais3Xxt2HbxpOgIdSq8SC07G27sYAw5WpnlJDiWMNlfF7yoI7B6lIhSWoxbU
lRA+tYavo7SKL+E5B9qBeaYnXPFgFZJFEMTVoPQm55ruix93WSRu5G3nYNfuHGbZ
r6NnxdKbgPVb+rdguQfxr3V6ZF0m9yEcSokHi3LfvJzUwJHA8jm4dwYMi9+Kq0XJ
HTS08qiddikav+F1siySduaBQnH65nZ5pYt++mSkAT4fPFrpgmLlTViQ3h6Cy0Ov
rgBUGrNX2ySeQUZZvNPbX2215DkELxfTRwubMekD41aVg/7XQigv7MmWeMP5e8V2
L2F5JxjtwHz2AIrneyegGha3s+6/vzd0pdSE59lGiXj54YoWFBONDu0D7fHDsUpI
uVAt94NBc3744B8/WMcYt1VUzGCUOpnS8O9NzUPijqlEvFz0qTlE6enZlrl/EGX4
mMtlEazzkS1obKxkhFX2mpJ+8u0lDMpM3lBPmzvTVuL2dbECCgPXUGPIN9uL08aq
QVlypaSiJ4EUzlLQxmwevEK6zehZ6WRSSzBdrK+j4QPK/z6VXn6xLBD67aLyO5+s
xJAeL2uyW/dNRNvImFTCDBhNMKcQY3gfbNNq0WOMw834ebSe/Va1eFsfooFc3u+L
JeFJH/4zFyImhsTMvvXlZGJnX2yObO4Jm34g/FUjYAr/kx901OBNYoBFx1rJBQOl
yoZnF7V4EGJ5evFQENXkpkMp2Q+OA4e1gELnXMfa83CH5uJf6eRBs/fqcsU9eqJi
k5riD9NWHOMIUvkprHRz2lfrDeM7kkP9Cc2q37syZrT1/3RgmQqily+9q0x+mmLI
LzCXIAc+8yPprKxyMGu3lK4+xr33eKRI1TB94ZXfSvWFWLgfRRBZ0H7bp374zTaQ
oe+38k0wjLMZkSE7mytrxF2BvdGxsES9Gk8sSn95dP74kcaBsQ9rm3589ZVGU72A
oofMS6jcgbhwhFIZ4pgr/qo5/Auf5UphoOeWgkTyIkM092NjJVyk3PSRguWzh8KN
YvtXrDjtpkut9PggQ7Ab3XOPgHRCCZ2X3pu7H2BywSYoZwNPVCiZbtjpxP+So6Qu
+kiO0YF1yUSznhtxxPENkvFtU5To/K5J8R/tb6Wf9E4fH8wnjObUXC9UEl0dySo9
+5pATHHVnVw08xuejPGMLobV/MCs1AIaow2/Ou7n/QHW6HDTTaRBbDYTJmdUdLen
JBvt7+2xsYpXcWzKYl6IDig+pEf/R7m0SOWUE+PPUUl9UwAD5bIqzrwnT4/3IMEG
fuAIP0JsrQkxj6UMM4m1S0P8eB9M8ea1awk4eX+7tv5K3GfU492p5www4lEq1QpB
ohB1Peafaf2pfonXx9i1t2C0U0wv5P8omcaQKpv9fBNoMFzXulyZzIuHjkJRawmo
vCzVQfRVpBhQ6O4M6FY+RISh40XbJwKHpeS80Vcy3qEcUv007wAr8x5mphKYA2cg
W5SmCT27jIoVoLZ/B2wgBaudIqo5e3Cqa2UUYQVZZPTq9DegIrsJQuIJ/MPKG+mh
oaOccxB63reQsmcUDfxBfggpQJWidhZeejIOjuqDoN8abbEpcSUGiNF6BwyVEl9I
wGVKNRdyKmxgp5JuCeEeg6RDvcYojxDXLRsBKZDfNZbI073flkUeafqG0/VgMQXL
c5/CY6TTxH1qwGCmYkHrLyewCzSXPzoJqJzJaUffpAs67zRcFdsAS1R9ETZx319O
MrlwsoLSv9HEZ1SjxDU8mxu5aznnvRITUrX2C0XOxlGmcwFs9Qu/H9OtbfUAnK1v
+JYG3DwjcrCcTyQeZFK1BliO77ihldJhMkratynIXcKGdRknHkcH8RV8MEr05Vvw
u7+4bxpFqKn6Z9K8SIJ5Xob0RqHYJGaLXPYgEOQJxHdyxGzCWFJ65ePGb170gPTI
QRRxvyZn2XBhX5u/MKAQ3mB4KYIKKNGERtLMHVDPp9ok3TvRHcKiwwGsAGzfl8AQ
ZbuY7nYRRf/BrvUUKygyC5gNT3gZDG1rv/g1xPGLLJu3aOozsxe/ad3KDJBL/oPE
xZC3b4QsJrizO8zKdPZMWVx3pJQgkwvageRN3QiNF1s4ZP2kNlnnkBz17lYbJ5Au
Ul1FVjEZrZuX8mvtTtt5qNWOKwipEtCaioChWhsB50sAGqY5UEJKSngsPCXu9/Mi
BiGOFGw6GRfRDK2O/NE6xx5t1MraKJ+gcDjupsgSpH0=
`protect END_PROTECTED
