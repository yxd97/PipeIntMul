`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iAJCRhaNfuCYruesrLTUc42DWcxnjLU8aV3bUNtUoCxlGyWVXK77O9/vHzK8uPeJ
mpeDUJ87idlgZJLrbfH9E2U3Fl1Ph6p/0akV8fWe/dFali10GSZAUlGY7Q0tFzI+
rZGxGQp/wBzC71SMFtVbP7SW6JePDd52lVfrOznGKTMv4QoWtrMd0B+arEVLt1Lf
4eUPKQIacyXGdd+Bd9XI8yhJ3lIelUBw9BBCe94lmGzrERygFPt//h94bgR7NGHe
tCaQqoQAjL0qBe2eHAP0Xgm94oD6om6fRoinDLXR2otXhNowA5cR6xJlrhJD6CiJ
O57vxKvEuIWzFpnB9JRHduFCDnDup4ovBVe/9d8UL6To0xt9nnd7Cc5tD4Q7mSV4
L4wut4oGqWRd0yeGpgPMExetZH+zL97PCbw+pLYdr8dexpPpu+m9EC9h9t/njUiE
O1u3XUTHAI5wYRWZJ8llSt2Xt2f9NzCQF4yQMq0pWuYWQsM9GYi09+1vSggg2u2q
BoOYS4yd+x+iFLtP/kqhPze+Q8jfX5W0HTrb+x6AmaI3dttts1gBjqMm5/yGSSVG
HZp/J6WQDO/nyS0dwIGHSfiCBYWCxYIvkK/thD6XvELRv0aBMnRksdMac3VQp13E
po/AWX34k9yY1aFTV4YqZa6C0U+ox23q7QsrHXgfWny0Zfdj1pQoH1AmKZLcHY8W
JXUYizmaiEiM5EVvIMXV7x1+qoRWVCz+62Y7PdPcn5v3szYZUDneZDd6Qo2mZi4p
`protect END_PROTECTED
