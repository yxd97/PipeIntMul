`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xouGP1Jtm+loOCXBzDhEOHMscTfr9oettAZ6LzL0ZGWzLJ5JTPDAHsZHzJt/1m04
Flh3bwpJVS6mfoMdVwgIMXFb4Cu9YRStTbmzE33K2C+j5jSqQEJqlHNPxVZNahij
isZ5WHj1KiA1sIbwJMyAno1rLSh8yhYBSGz3MUPJVQ4Yj5oQpoy3lurhZa1n/VNm
Uti1nJuvyDi5sOIBEXzhdRocv870n4T3WRuUvQlFSvRXp09Sg/yIqt0reBEgY2ny
QTB19MhkV048iH3eAX9l3CRx3Dx/7jrqVrb8ArFT/0j5BM1FAPGLschvCrzimaD7
pRRCGkjZCBISnvpSewVsGKuJ8lz3b44gGIeOMBtYj4YZSuLYOCjPjNC/AjbcASdz
fxpQcabooDFiZ+Lw5/8nxLOkCjKMUU2XwMzcc4c6wscaOgqjRkPIliO9odVD2xo1
92WUPxzBIP4ZTUxXzQGSW2QYGAwcaQqUmtUyspAxy/BNORBDYVRNDinKBmKVNh8E
04HXdRASQZJADBPzqjGGOM0UuPlp9CzRRQmPgGSKaInZVTOVFOhTrELFm42lBwyw
N7noN7GDNNNO/Lf+wAUI3zBfvk6FnbBeEEUru/yIXFLKj/cKjoEGW1FctqXcgrck
seOyD3IaNr/pYOfoygw4MZpvTnMHhWqSM3B5rVvv4Is37l9M83dZrvewmrMYG+di
Wy3jAAd+RFsDhxVGENVZ7Vl78R617vD68MhrHJaFUO+q75qw2Mw5Q9j/byiXsWhj
66k2KD1r/27aZWlCKCJyesscw0iv6wQiedzQqKqVBygoO7f2yHaHIl+pmTzKBk1W
ke6enoWbqTqQaXSfL6tXVYPSsVUBBuk+1VZdIw7sHxe2XXxNXKghY6I+3fghzE3m
WkzfQSBlKfJ33poOzv4jPdspnE1j2g8hGpFhfFP1MvOl6z1FRSHessosEmyoANT9
EoV+dTUrWaMOhFkCGhj52jSMU9nL3dcKAxsz07qFN54JlcX0LcKE7V7JiAQOIYJ2
`protect END_PROTECTED
