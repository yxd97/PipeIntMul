`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6tRrRkiM0SujEXf60F+NfKAxN35seaDu111s0cQmLyIfP7RD3npTLieB4qejtQwq
PpzXp+IlgRCpfePeO/58TQhi898W37oyokerySyrqIsbYWIU4yWhRXbHVEEth8Q+
z3vfE/qJlVPuhENjCQbV89ATTj/ge/GfctlzvZgCeQjfjonQZCEvT1NTH//g1+v/
YsOSHN3sgMk0oVwvmlPGB6A90fa3g3RDEZvv1TTfLDqcou8EHDyeXBF6hIvGZsMp
BicvoWTXhcdLku2C2aonko1iAcTbVWNi3THVtAH9sjd+OIuZdrM94lwD6aLoXoXA
Y78Db0bqNUIJ80W36As+qg==
`protect END_PROTECTED
