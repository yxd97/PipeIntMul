`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
52vEpvNjnlnxw0DGT/yRdXPgsX3+36z4K+pZGBaMzawrveKwhSFS5TvpvsIZZhMB
5ypdv1XXuhZzQEj7OXxgowAfNlLKASAwaIMfRJkZsrhSUY/NmUB/eRcxZgGkz/Ky
XcCIv0+Xgw3y5TPHY/IDJJEBFAs038NejuVey/fLrsvy21w2aOXf4SXX8b4C8zJ0
y6vNWn992Gohb+OOLwT7hdOr+xLMT5eMLbdLGe6JvPCc2/0bZpfTkc9bzTaMBNde
CVoA3kMRqO7DI0+byYBqRJTjnZCXKkoeu/14IvE1ZrTeAAL105aRfwQx6cjIfi2A
lhsXgWXq2tGKzg6iP/95HUv3u3bvJnQIbI8zIqR0qyjB6KxC0q0Uv43aS9TRRspH
OUIRTCOfPC7c5lmA5cffFJMOhG1nCyGxtN/j8dx1dkP5YPWHipI1DhIxe0rxorgg
k7XYUxOtCNh3D7gwxrqaaNSgixqD++BwlxCzus8KBteZdk5w00VTgbRJ9ZxKLW6C
54huNjkM6aq+LtGw6KJyUk+GG0bFEdnaus5XK5C8/HF6punwrNRxfqeLvfYdMxJ3
rGHOZTeSgf5+v5Ipr2CYsL8ttEAkm7jwBtTmMsJ4SNGoQzIlVUcZN+MFxW6iDbYg
QIExCenEytYTAfwNLPUshP7Jt2H+F70we9HCzDJFNa/9wkf4eH8fYEgcJh9Q27Oo
E/HKsS0h/4jTxrnaEpeAuON3XgbM3TlOUA2aJ2TpFVU3xRmJUEkXHot36Q/jyhWK
3gcH/uspfpMQO61O8WMUb7Jug/E5fNw6qHXtjIzSIaZcBDsyNii7M0zv8Xy9Y180
R2bTSKqRS/xbDP0YnhagAUKDFaBz682DTG2REMjYin84OkfMCjbxap28XEPAj2vA
9Gz5k9tq77KwEqP2IR4kEaaKrW8xfVGbUSqo6ckKkigvmlhqR520b8v6VKR4fh7Q
eYOtBBhqCqMIqGNoGSbEo+ondbHAAXxYV0TThBX33sXzA2HDCR3w3RMkCynfBU7q
TRr2DlRUF0vS/i/gvMq7e/ZID5eauhgNePl1m0qRgjF88Cy1fdeuMoMvspqyPXwp
IaZQmHN3N5b9NCcEM3DI9/iz1/tYKoc70LNfU5mcoh8fHdF18jWuNC6Fd9fbagps
NlQU2AfLnglSg1nakf0yXIDA5pNAHCZMt54yBQfW6Wfg9U9E/fkEsBwg/25dK9Hh
I0jqNj33rf9UkTwDXrUcnDG7CxbaL/TxQ8klPhXy7eAOd6UNsw15O7ez0MeHR7qa
YpYnzvoLCNA8POHzCu6ZaW23+sjDZB1fr8qfD8QfUQLnfEDBx0wX/IaZjxf5/TR+
K07qiaqYvYrpITBFkyiGN4p4sP8s8BavG819uU+jcxpyUouBaaedLI5IY+yetijc
fS9WOUWClLxrvZXhARtKj+xppK3r33Oq2/+eh8QGqTIhafK7kHQ6F4wE7eBImwMt
0hiZtDqw0BI31hvydHbAg09zyjdY6AxJ96nQLDS6KTYuFNjulVGtEByQ+gC17WQi
3V61pAH8weQNdjxqVkFyt5pAawRpqba0rGMY+9m9cynjLnsh/jbwU2dB2LCJMhL1
/SAQKRhX/ZBGz824umlsVgkVoUWgWj38KsumOwlFx4TesIKjb2jF2vPejiqaPdLa
1cvUlRXXiXM0yhu+ghPvlsEtsRO9mPcFqa6TVhg2pc8dVRlCswT8tOjYTUm6wPq/
3H6Wpv1L7CW/OBo40tPyjNvOqPhaDCZezeAW0mpX2EF7k5XLyfwxEswJDnypUMk4
IuM7x7Hj16m4yUKIyBnEmvBo6coZZEV3+6Lafk1Jq7bDtr4n1eV+3KFOa1ZoGmkV
YZmeUKA0+CE3Fqfm3vE2twW+kNz1apcNHUtZp8lD7IX4JpfbhB8BObgF+PbCjuZh
9VnFGvfq7F50+f2N0IWi/VPwpu207NdgaMxuQ+eQEpZkS+d8VXHyRMGrhzlu5UD3
wo70FQIhf0slT169W/ug5Awop+orEgWUvk2Wc8Lo28JPaYw4ftUt+XXp5Ic0Sg8P
pED4cpBwvorivP3XyjBrWdNl3p4s6blfCBlYL+uZk+6AArDbClSfYql1oZRQulRz
MBnnPTXRb5kTSnP3RyJJmIAUQpzILe6yCBYEIcWEqtvQhdw+RHEZzL0p/ZYNS/N9
R73NPt0BZraMMoXSfxCeOS7zqbMsGMwvk0Mu5vwxSZZeAAkCrd1LpYQILJceeAlL
uc9U+Blg2oRh6FkXnZtDV1z/ghqpLo233wZI+hPVfA4C0IvotCHg8B/593IIhfLw
lK4w8Mb3bJj5+X3UTihEyqj0rpbBBqULye4Ljo2bFluv0hMwE2Lq70MblRZCeVNj
WCjN/MbO0QaEzsJSc2fcE/WREh4+dSYvOh12+6Qps4obwcDD75QGrrgWKBPtTaLG
c6hMKSgIjbY9n1x1nAhcJtBjecvhIwJ3ga/cNg5jWVfZNnkLcuzpIA7YMJEJP1Bm
h2D8DH9zrImBV9CjRpXEN/phpEtUVA8bymiI6rFGBz9foAKg+W19fOF2b5mSJoDz
npX2c3BAanpl4kG0DccHYfODfZeUwq6DciW3kFmphPx+wIdOLvxFN2JGjImLGVF6
hyTMXbHOpEMRDPaxmM0mULKdOaJPJUaYeX7y9cta327tx4qY8MQShIPtHNAWTbf1
uxwMZ5wpTEie7LmIcnhFwwt1fOCMBGc+Msmsh2+PFftFyqOoFruCjcQQ9iM0cAdT
2FdwYcIX4oAncBgvcVV6EzN2BN/I0WOPxje6oMYdmWYIYY3ATak1AnGzE3xHNlbs
X8ZPJMDySjLt1+4ZDh3r4229Z5BvxdjpnGkuhIcPif543uEVHBtgt5boYvHiiYWU
Hoj1WZsrSPRnaAJQozdE1va5GASQ8xM+s6p7Jnlo2waOiCVmtNeiLYKFlpOc8Avm
iTVJdMMXTKr6VI0Zh/0gR5GiupYYbC6LIeTnvNwOLYbcHvRD44mHvS4AJM1QCCHH
uLE1FgLC/lbcZlxb6l6BB6LPZJPtwIy5QSPnS9PaXuDQ4TlunsiXueKP1GSQjCzL
STtuPALNFkxm4uzgHMLqAfeXeK2UGqbrDe+19cek6Q4q8RPM1wrhAHdPqzw31pzn
OFCj7GQQu+59PiYW2G91AAL/jDlDWoCQMTV2E/X4Paw=
`protect END_PROTECTED
