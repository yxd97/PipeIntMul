`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1E45wtXmH0tMx1cflVXeUjxA1kFBCcL86Vhs/TOxLIRL0B4bYGCLefKGA6LR5pYT
HiajZ57LcOvZ2Y9vQlpLrVp6q0wMn9aFRz7iqsP884I90qGTnEs+Qp9/gAzhHpQ+
IyczSlx3PYfpRLvhzBvV1578nB75qnDFk4LePgOxHUR1YBh2JK/slpEXpZvobSpv
n3JnHTCQ6qUFJkNNWz/y7CzBuE4gV0FPBaVXFzP6gCgqli3cexD2obp5z4sawNnq
VFApnUX0xtlmXSDSa4kLBrTftcbflwNoEEh/5ITURp6PETRQ6I0EVsRdkzZn30mo
C8eTHV0P6DL1E2a3GtYzGoMK/bDWDmnjvLfH3wvAuEWt663Y5Pv+HUxJhHLO2NyN
t2XRdfO8YbFBXx5JJ+zM1ARlna3KLTEqnhhxykZQMClHKud05Wn+gB7XZgp4CUCD
Ih3Hkrij+8IpbphmALhR0q9J3w0V0Qatuqshke4ZBb1KpS06MTmofnbbM4owNlzR
zu81/zAgo5cyyusmn5e5wer9bElFAVbBeEsuPDGEraA0ahuZmT6N9R2ukTHQ0DkS
dV95uA2Coj9DBwQzdsDtE1WAjk13QQY7WxHyk561NHCGAqV6bIzD6C7lMvzNDDLs
tNykMsqVf00MHZ7k59IUQROg5ADM/k0wWMdMYgA2+H8=
`protect END_PROTECTED
