`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oggsfuMEZB5NCmUj7bh9xhLJXLcUWnaBDjtbai2zMzm+e453kyPAnigc/l9I0zzk
1YW6lRvC9XMegwXp4HON8Dwi4WmdA7MO1Wt4zBNbFCiT13urgzEI5/moUhwxyS9r
qhNi5pOErbJExDAYHQHd6t8Q6Ud7m1SePKgWPkFQRQW4CeANCN4VTWmZskvFhVhC
wS86kyIJDV3TwRh4KXPy2cyUfjIqm4YSivsM4y6J+rF8YR50rtDD+1Dnu04wxrxj
IcWuFoKZpXVwt+i/8JwSW7TMVgm2wZ9nQFnRgujiAugFITRq5bSKQ9ZILW64AuGk
xzPf+BjTdDf1OUED36TQDIewB9YhVl3XJSzA9rwBzyN6Ks5SC33tiBvgcCQIYkRx
ahXySoNj1XNehleAfKxf7GbMdUOYxJRcxWNC9mErnA1tQO6gieXFGh2LMPfe3wuD
TCjDEmEls3rh6am8fh4qovsViDfa8XGsF6ZM5FUZPQaYwg+jnYvr2RqTQjn2j4GP
vdQeApc1hhPV1TVcgZrQJ/WEfIz0HVV9hpjSF/9Qo1qjkwJS6TOggh+ke8ihdnfv
SLvpNMyK0NYNkTLKWN8NjRzcySkGlIVTDP+tgn1ZeC7RXwrZc9JlkzQlfQFG6MeS
L6FVY8aA6RGelBwQkUpyItZ/Fo6C5hb19lguo3Emv5SIYyXfk0KU3qVSsW16LvwI
e1ht3l+wX+YR8jr4dLbQNLjDww6iuBthaGfg2mp+CmJjiSSXnWAw6Q4vl1CcBupY
ROObEJs5+WSkLa9xQCxbV5ehawfaoHsaUR5ZKV5k9P5OX8FpNiOfyoyirZTpuQI0
Te/AjUg+EcO5/7jgBHxxIFLQ2xonKLJ8dBv9hGDnNbLtjxbJgYdVBCWLrCcINfVl
w458oUxjFh3tr7VBTZHcfbOzD0COWgEWR8qF3YH6Om72Kx5fcKhC5dVeK4efi5+N
KOabBULgPBhP8dEchJFQi1hvE91jq/SKi+2PRzcUdftG3CN6zQc6E7pp5oGC0k9H
HRAiQ2JjhVMtyZHfYVsH39ToCmNRssr5HeMygr+ST/r5c48H3oORQYG008FmqIF4
PjS8UbqW6keBimJnTgeDUQ/3U2Fc3Cz7601hGenXhUeIbzm1jjkQKvtOC0hNX29w
ZnQBSTvJczk83J/zEC20xltCjmAg393SEHDtza4R+yhqtAMvDtN5MLzi/Q6Z5my7
78yJ5D12BSrBO4mQ7qcTP3cBSE7FDEoAPBbGCGANReXiDbZpbHdAtwkT/j1CBi7Y
Uh45ZQp9CN6p75nBM/m2pXwl+GD3KJQCmqixFNOaVg8iVb2qrPE9lEBBGcKG0ck4
ybSAyLznZ+NXORhsYYjP3sKojamCpJIeTERxwKlcSANOZqjt3f5KsN+UTvb2c8o8
PUcM6pDBCXCiq9ppl5rLmaaEU0sUPR6M5WWTpM204tA3qoSRbTjYq/q8fJzHGCjL
LPKIguVinSLF7nWmVZtpZthoWi/wIA4giUYAe2i/scwapeUYGDvs4X2r42S+VJxu
fTl424joVcjlTbBEk7mU8+Him58FfO44a3TD21NVIYwNZUnzArHqkI6qQva6GNtO
tz4YzeLJ8LwiqM7G3V3cRk4NhGJcwZ5rBv6XiXYl6+s=
`protect END_PROTECTED
