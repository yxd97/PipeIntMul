`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c38QJE1KRxzlvEswPMsF1F0q/RFXXQ1sAEqJSbEtJmSDL82BwT5L+uslT6ng+P1k
AQKvCC+qG9YsAQWPn8DzQfe8CHVv8N4pWRCse5MDmA+banvAFy7MHMLtfdxhWcXP
4PGwHMHG3SDcWN1HYihKxHj2gdfm88/1Ltugq/a0PwF851g7h5Ooah2WZnbKa4MV
KQE7jtV95kNnla5sjX3jSL7zwerK/t4dKAqiUouLdRwGcsSqVx/Q/QqQl3glkX9/
eQql9U0b2nTGLv+TsAnodwGCLVXpY8FFpLjGJXPm38+5hTaMAmOOWv1d5X76gFbX
7qVvnrNx7R31EKO5ad3sykewP1ZI+g6vEgEh538yQ/X5ROWhEHXDAlU+lhLUPNKu
D9/CiOVQpjOgYC6X15U6JOuCmxhH0JcJYOMHZ0MgD2M=
`protect END_PROTECTED
