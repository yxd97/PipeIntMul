`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KD+R+0FjBkhv8jfOGLGNcy/RlS0M3x5SBJD9YQ8MRYe4U42NNlb1NpJDHds1FCAe
SAGl2DnEjMROAp6A5+bCWq1XCT4Ge2X/mpW9jULZ8ZtpmcYCcGmibiMLPY1NRsRd
Uv3jPlpBUZ0WfnFGL+qv3wQ3Hcr1H5k9vRuvZY8+neGdEgK10uffcFOWl06EUUBV
Xa7jGvr2ztKdJN0plN8t+2XS7bSG8VEsWSpj+Wn94WPBoI/zuasfwF3UizNzjS1i
C2K0gZoJ44Qj0nhEFYZiCnpbxSXCnHFJWCdLSaqJ4kgTbsJgB9zFT2NtgYqA3VZg
hb235pfQX8U/T0JymCEWyRUmR7R1dTUvtR14O7jqCK4J1YcCkFGQabbIYBHA937D
eohPCZlhtQFqIbjcf1IoyO7CnKGe/JmsSLtfM2FSpifwpSlQRngzZwrG99Wvo5wW
q2wSlF20yL76fwTFvCsNL8JGKCOQ08ObD+OyUugAQoE4bWoxqa2+fdgFV0zku9Zp
qhvWPeDHaIfqu0xfihB8fg==
`protect END_PROTECTED
