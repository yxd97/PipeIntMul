`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XoMoD/Qj6tk0+HQBhRj/xZW8TlpIE/nWf6jKUAYSxX++rZIcCVYfYQyHMPuCEUgr
VM7Wq/gJfDXtfVBGYTfI7MhcDDxPK9bmSx2NDS9K9GNncTg+80g+YlDq74RSWq7r
Vjivc4IstACWNvnQClSVF09sGJD9+ZzMFn9/p9LMI0b7SvuuQQGywXgNqb5ZWxq6
D99Xlq1jAyvDiuf5uWGQNGueRBRFFtYw62bFUe6dxuz/zDHTmM7Sg9nFeqjwEvew
PcBKJ/3TWAA40Qx1gPACNDS7xveiRvDQOUg89HibpEO0EY1BQLYxr+CPm00bdqSi
CECuFG1o2iHgOn/q+KsjDvGp8iQSNJT9jjuGRVy0LV2I8fc00Ny27NnrOhcRVWq5
37o60bz3TYq/O1nKdycvOgYLwSMpMdEuNmj04UvhSK2S1CVnWt5OqWKZrMQcJzFu
lPnSM6noHMzSRxJpdrFPu0R5uSeTleP02IqcdvW7dvNnQhk+SLy5iYaePh51NVNt
aoQsSrmyY/m9vfIW6xEov636Es2lsBVtimUZ17rXTqA=
`protect END_PROTECTED
