`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EbJsKHXwzUY26oHPc/ucoorWR0CZgDf/q8N+dt/hQtMEIXiOeoIenKbdfkq4RIIk
xjSsOSFxEv5tf+FqSjgnTxs2vvejgtI0Lbcs1yLuecOuXJWn3xPkQdluGaDn7y11
oeJkYLW7Qsbedf79JT1f6dkqDk4IhMZlEN+ad/cYTx1bp2ggh7B5rNrC6cvFhDYj
clBzJrlqdomMGptY/n7wOunyVMWv6a3hZyF1r7pPa/KTPrv6V+Jb7P78tXoGdcq3
C8p3ZiZ2I7K0QePpg4rg0A==
`protect END_PROTECTED
