`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3MEseCCvki01A2SilDtQd0JjRaeiTsLTx/DZmkE4y/QgO0m7HUQA6tudiSTeqls
S2oBbMyAZQvbHa21uCv6VNxHqzaQ+PmnfUUrIDblnlYN+j0fSz2XgpxKCTe9+MXk
Mf6kshmNRgyCSB6sNKLjpBNP+fgCiD587/islzjQtzjY6pnTUJQ6cvuDSeYiwu/S
UTnKetJ9QUT5dHlpmMIGwVIvkJMzlWcWMp/DKDFsH95JPQhZSRjRCChZc88pwW0R
ozy70qOG9RbKey6EwFssz8z/w7HvdjMbSdyZQZHPLZ/z0qxOs4naLbxTLWdW5qP4
pD6r2b2HUx+JGKz7euaA1YwsVQq/Q5EGMc+YSXKQ+dfeI40Mox4N+1pfZgEd0NJH
CUyOTA6OD5rAkV8XbJxP1A==
`protect END_PROTECTED
