`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bvtMYruC3xVSIV97ENukK/fgsnl7/vbUI/WXo+O9S9vi3MMU8MasmwESRYuiyhQd
35unsYsHM8xLdTSdb54zuY5zM6Md+x/VSs5LN9IdaPvSzNokBfc5WNzltPZNOY7V
kuhD0FOcRy18jIQJ1y4/TwGDZMrDp8O0UZFS+LgsmQq3SUQ1uLGX+x7KDSI1lwCq
ZvgLP2gnvTHvu9Rc4PvVKid7Xivb97eC6/Xr4bFQTOiRyYJnClcc8TzxsnE6u23X
Gl61O0rwb+WVbgFwiCZWZ17Egv+HCw9Jegl+Eiaxlt32RhEg9f88ijujiypLrtbH
53MgAFiP2qocdAXBwp41xDF+GZZAMtc89A+LNuMNF4DRZDeG6CeSMO5ak/BU6jY3
F2/l+C4z7T9pz6jLlDMnNg==
`protect END_PROTECTED
