`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jwmZ9aV5tnohKEO7Xsrgp/460e9L1ij3gByqw5hPc2As63B1EP8Ki9pWP+U7oOpV
PIA7HJXlPXtfEp6t8DaCzg+/h9vZvx5D78lD4anfMFWVUQ9QE4shM8pr1mqXUcbE
3+OxLc9r4c6Sw9DfrLjAwYKzR9m0piSE7QnMtGmzVVbszEMZLREHNEClziFXYAVv
s2VZ8owVmMlYfetqmS2ZgytJu035CMAFlvARKcFWhz4nHNUVdo+N+pWf1wTG3zcT
/QIRk8iXGSScqQSvXghZGg==
`protect END_PROTECTED
