`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGxvFwED5sTAvsmX/2iNPRIL7tlGmc0vMo+22MG1LecsuGzY6R0INju+hRBmt2ZP
cr9626BGE/ErMPVQWwCPD3X5Qf1yfWz9TxjreX7VvnknfMLmHhBWwjIGK0b0t11J
qsnwSjllTkZMOxIVeQvfs3SnJUpvjSxF4jviN0dzhBsZ9e8OOoowiChFWY2XxZOy
UN33cJWw3MoGdvXb5ixAFAtnP2FjvHU33CtzOl70fmnZzKu5RrcYktFM00Xqj2BZ
blLF8AkFuS74GIIwGbAExxqo+IVL+mqCZ7AWqTgGzWAfCsqzr7lfLgBrGDAnStHq
PTKeR4f9H43SjF1cgIz6MYEG8P8uDbXL2RujSEIBUVTDQikIGL+QAFhF5Ei/NY5A
xb4wnpWMGyFBAwDDqrt58DPl9/g/vRP2mgiBvVlOjlTJKO8Zf3hqHnqo/1dZtXk8
0aQMWZNU6yY4SPq9hoFdfUfgAHeErM4kbUDzt769zAw=
`protect END_PROTECTED
