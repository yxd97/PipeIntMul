`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h1rR9bv2Z1g01olM6Vg4kqEFVQYrxXpJLVomY5Rj3oXT3BGzP8KTvJ/ZnJ4KrxgK
hqLbt69y5dV/kfigLLrNObD0jOOI+e/8d/Hhi5uQwzeN6LA6fcVFD2PPZ8KIwVbC
qR/DU8TsznnuFu39/769LIqPggMgDQwB9gxMl/VyVQNxiJv+v6QMZiQ2V8Ubo3H6
gBOfv1n23Mqh9Bm77U/jQByH8mC0iYOhCHgp4eyszgWS6CyJ3GZf1umn3xAkF4Vp
HbQoIe/e2xR6PRNmhM9riDCYD8xiYGjz8iJJ6m+EKnmRAzHwxF89kc/xUOXXeih4
Au0IV8HQ1B5tuNp+2LJBCl+1Nsmme0TshBblrso8JC85g9D5+HhJuD6DlsPOAFmK
eM+6Rx/t50gttq3cqRsM1A==
`protect END_PROTECTED
