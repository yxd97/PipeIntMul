`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVqu39JleZEZHJaUe1nCy0PhmJyz+pzqbbXbFvpwT/4fEHwj5SEdk2W7cy8W7Rof
l18ngdPkU7KynHmPTd2y1m+P4cey64tS+8keftWBeJ52QUSl413TFEV2c0XZ4wUk
b/WJgar6+ewHKe6xNZ1p3kiP83MV/NjIL0Qk0+wVhjepilKyNYbxfrVsrtozqSgy
G3/UjF98L0XIUc+z90RxpY7QUCKLIQIH7v54HDdlrh+cqvXfUjCdLmYLaNZPpk59
ZiJmzEg/X77aQdLzWaN3LZ8Z3RqciGgMKRHDMKZ3eN6W6qwh1Nw5n50Mzm6E8wIB
BIKA+FPkyTqvw6+Y7pxdo8vcvLf4uT9l07Vcwhr+1ie+ks2RPl1PHyCBvA7m/A+e
Tfn330b9wBhH0pP6TDDuqNVjmRlweQDtL6dnXxUHzn3WoH8lsn2oXUhxMiulH61U
`protect END_PROTECTED
