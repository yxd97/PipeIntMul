`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tzkibzLgbyD9wLwblNz2Cu+kzZtdoJ/apIctmt48j7kZvFrt4Uv2dBp0FEzMJnyM
Vowwf/verdnUixuAvGO1VS041Qf2TSBq8dGcGkRxZ6kviPB4RmLk381ycj3BmIEB
ut6QrFlgDiCwEDnWSJRmKAmt7XMFmMiH8BqbUgNknxscrXurP2OUhxLvV3562Jnm
uZuytet5suZxSwJqBCR9R+UL9wCQu+TQtxeCd2eYGw43ipgLHHEXNJ4U0SGNG+BA
S3ycz5a9v1+UWX27XWjW9+hbD9T7WHoxOXWYA3DT1QQRsgPx2vHIqlT2uZT9HAnt
JiPA0l0rihWwQmv8K84fSPNdF0pkmFHwt4tjnqGYGfodbi/rZIQtYHAmUUyfdR5D
cD/YKSndHvjkAawQxm/fIatMvF2JrVp6ikZGCRVvdobTjgMkV2LzLt/6WB8NuTAr
N9h181LQI7fLaE5bZBY3oozRR1qb/jWxz4XVEHifsnR9ObAKnZxl/iEIYwSRnOUL
hT9kx9x19sVqSP5duP2nRGQTdXOzOrYcsyYB2hZ0pPvcw4soxj6WimfGAEN5s5io
am7XIXWI67MmX+R+bv34EeCwL/aD+F/T3Yz94wCmxCFcGTPN5bKkIy6FVZttsL/W
+heS1u4SAOMerajTLzCHhrDqoDO1cks9rTIYBpYq3Mz+HgRw2drVKqak+NMsFMg9
/jvEiSVPL/BIpxSIEsINQ+gCPDA8IUss0mKrM7/f5ov14s54hpqwIEWoLAZ/xV63
HDGuxQUWlA3ynP6+w9eZQpcMton1uLyNaf9bXrar9lql5rP8H+LiFcuN3afPzBH8
UFO/ahtcH6L51O+UckOl8ZSjXKs5qGloYTwfy++NzisnlWDJjk0js5lkUFrw64Yi
AoWbnSizXQhZNbdg4CT4huED0h5vWNL0+3zWX8uLpHXD7XbcK3hWQdKYy0qo15Br
`protect END_PROTECTED
