`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O2ZknrNJCTRS3ilha3TX6/mzdWNVeiHTACbWeYsFg9sOZFjn32tf40GKoYu3Qr2F
AHPJrvifcyl7qNpAhF0IYGeh1iSGR9ACX8nydLSYYbFqZPa/o+5JNQKbevXlwNHG
30LZ6ZXIB/XU/mqif4IqbvUOv1wEfUWF+OZCPC6nQlMAbQdID0wCD75pK2c46q/T
8HduL6uHZAe5M34nD8xDsyScXT2gwQQYXanjuL46rzP+y30V/EnzKvrm9FAmA2bX
cjmIZCaxY8moVs174kB8IIRYl6P0y8JnDUlRGZUQVVtL4kW+ppUZuJdIRN29ncvb
29xt72LWGcB+qQqcodoKOSCNiCWyqWnlK4rROz/Bnl+P6SCyZW0W1incHf050Q8x
kvUQDMFC7fD++tvfYuyXkDEz8Ld9Qr+Jb+kbCXw5nIF35LsPGYQc7NlN5HTQ4QCg
OEr4RSvTyNXKsfQzjK9fHN09lvnAmAS8xHRvoJ+oUuvckLgtoTzI41vdP94JfS90
GozItxmfmXDkthqAD5k3b67gCOPWlV45rzUvpE5/GpeZ4z9fieN3Ocoh5AXFy78W
u1Zu10wC8KaVOON1SXPWZAGLFWBeN7CJENkwa1ioRCLLyHcXfvyJGnbdkPA8LM2E
wO7IomZF8DsTAuNPztvbr3NZzK1M0zxAK24vP2UyZs8LrTd64AQzLhGAnJ+tSnpb
gRkVFCZaYcPzGVc57VQJT4myxRz1w1SAMAqqIcyYFaNye1pJceAo7tvLIIEnlvms
/eJjuC5PXV5XVeUQCbh39j6tJHComtfic8cG6nJ9vPfxy/sz6Tb9NHLHuIMPx2wU
0PPB2oMy1bzTxcNFsSvIE+ESgp0KyKWD5yA04qY+CO+nC0kmGx+2e3E+zDmsPY5b
e0HbQbgFDXovvjkxP2mkaLPuycpSSgICT8hv1tKQxoXO6M9/LE1ZN8LQKg8XnIGo
mv2DQvOwIN6TMovtTQqlk3XLuN8XE/EQ/QvkjI4w7b1F+/nn5daOCp6N7m0AF5WQ
qlhrB4pnFhkrxUlNG85kSSeDnBLt8qIg+dgNlw7zyA3icKJP3odtNa32tDMTShNF
SNCwsq3A2GNG3EXEnfLZP03VzPUIEezzIwobf6LRdyU0RAwgRANoIpUEEK5GjkPm
JGEvmcroJAg6weoaXXisGkUqlsBtVyrD/GJlU2bMs7uZPAZ1pTT/X9FobEaemWh6
Cd+meYAq/oxe5XPz+WD2hA==
`protect END_PROTECTED
