`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h33dx3xSHQeoin4b/NnmT2iIhIgu/Xh5bbsl3VX/XNlFY/QcPjfEy3IpAVPqBizT
Gn+jdv+5re2OHV/tkbPbz1xdXw/kUYzvrd2TRXjQh8vq6H1U9W+aD34FfK5mZqYb
6qp4sHpK3VwBfEl67EHQ6Tpn9G8SY4hYuhmD7BtbnJ6jhabyydyRffNj1NM61wAz
o04i4dRdecHgyKkLkUVuRDlA+BlaGfe5FBk4yDpoqVEeeTjfVMFNZAhVFtfIhMPV
xBv1yfvB77pF2l6MBlCdn78DNonXKiGD0BV0Yr0LCq09jp3/PjF0rYJwewHhRGge
SO4ndcDTxb6lM/0qiaH3BInikyRqevsJtlERjwrE09MS3orgMN8JqmHzZDhhpSjJ
+mUbh6EdcFBb9TMBy/VFhRHcMW94WFhZEe0QTxdTSPe1rAJ+yL6ghb1A9oTRfi28
YseRxeYUr2MrYVyXFzSO6YwjYvnne3w6yfiKQtwxk1KkKWPRox0oqWs8/+oJBatp
QmcVogJOFPTVMKJQrHFC6NSFIlmNarG0B/jhNcmpqkDaLapTsU889+I0sV1QYiGc
UxQWGRDlCLLtsPBA3fwTozTtWRr+cpj8RWKCZQeh/zmOFboyJnFfEZmg5097amrX
BVrA1foD6rqVx6O73nfbDi9UHhXtMQ6yZDAqwOHWx5WiqlMB/Z2oCS2rlR2F/aU0
Piai+9So8RuOhKbdWcaI9RWhEOuKT+H1z2mWkcyULhBwtENnTMNcEjRwiDljIxWs
eqSN02n2HoWa24jxo58eRvwz63ZUnA0QePaZjVU8YAiyKkUEw5j9H5t7t1TfEigy
ICgbE1WT2uhCkpOe7ypbU36Sk8MRWiTtm4H3tpbyvqYIp95jEKRmzcbUXZ+147a/
UiJAmAjQwGHrDWmcZr/ROYHItXBvN921rxPNUss5gOyhghDvF8DmTRJsPp8Jjo5m
rM/xUKpL8GEeWZ7oAIwcY67gIFjyI8QEzpoMwmvoynHa6AqtU/slaXANt57rny9R
9qKTM1DUBNXIBdYldwB1su7oJF/tNQOZOqZRIWyMApVGfA6+Tlq9Fnpp30BXp4KD
9mG/Yd/rErfyqlmUnIrOg/8zV8+FZwrNr+tjc8dbQ8HNbQLmpuoreTdT172eEKUZ
Lv6oODXb86+t39Afd5v5ma0DzK0+tQ7S8MUy+V4lctydiuZdBYGruafjcET3s4Pm
wQJoYk6CwkSoEp2Yrjzu2pNWxZe/i3OB1FP9ijDYSaEMFJ+hZfepFPwqslhvV7KV
NTOaG4tuMV89uzZKViaz4+tYM32L2fmpqAWO0X7IUYNB0rFGPimvxmr8xzJSVjcy
Nkg0Hma2cqJoDYB7Ock/s6yVmNTlFGsawYWmCoPQOF6IU4YOHA8L04BToOo8N4c5
MKQcRbx1y518se4Hpn6jm7BMEmtWTIyDqsNqZZhWHFT/iga6UCug1jS5xmSuj+Pi
8Yb+EraGR1r+lAWtBSBQXygS9K0LHuZzjqapLv2QbwNw7EspI7n+CzydtHnJ8nU/
7+vHZQ0GOEeXwPuL+WwwBBFsVXpOXJRTcuoxEssCV/A03gcg4sNbJs1P1lKEEmW6
7xEv4lc61mA/3wzU5GUPtp0XnqZtMUpCE/iay2A6mgrVAfE23UwYD2n17N9Lj8kL
04p0e2JYzkURO8wRDsE7jsVZXM98Er4IRaAWfDzpEqnNnNQAW/qaCxpOEdPbYNRj
LO1ErXwOThSMpQ2FRdS8hVzkOi28TF0z6os6pwiVAgRr1MKXiP0rrLIpv+qEX+Iu
3mLPxFm+LmgmGMK8j3GaK28Cbn9XtN0HzXRO3TuCtLbJYD7jInK+CoxadKXG5F2D
Y/4mnz6hDwB/uoE11BWymruCsm/DL4S7+24dAnA5q67EsZM60oj02ZgK5ldnix2+
3zY6eioDIMEBuHq0HLcZc07QdjaVrhNLm3RLzWVgoX7Cb8mvdMFcZTKwpgbfAWlS
Y9UhQDt+TWCxcbRqLDBvNSLjc4QU/ACtquoOlwGUvmHkjd/FvkoWRgl8wUyEylPM
R5ghztrdV0uq7ULXLpGsZUdw1sHJgKLX21Oh/bA/9XG/KXfxlKr9gAgk7Sixcaa7
iomtRMLy+e8wENqdCFS/Vc9YLIg20yGPbN7PM45Ib+mqWnvdYHdB+k1YDNBAWupU
RPMSfraZ4Xh9SKeAN9xyPumnBTTC2gEVjO56/TJjRXL+zebavjaoO7BH262wo754
TTih0RUFLrS32ono1uFBPu21GkprlSOgta2k84aZipflbkFU/MTO+p0+9VxLqW8d
IhP6krm2C4gKNiwhad00DObFwf/jKVbM81CeIZyd1vlJWTuE1T3rR83zErw+nXJ1
ZZIi0TPB2nEuGLA7KVFNI0M5U9IMmDbtxrJR0PNkZTJjDlFhaw4S99jg1ZqVvtVH
ndCj8VSiWRU4LPtQomlmQMHfwrVby+Wp/i9640fvC8lJ9R0fgJgHrrBRUW/ZJCzm
DkiXMrFSrJ7k2EQi/2zI5gHclchtD57ew1jt3pc9FK4SBU9XC8+Ciy+YOS1NIVpN
eNzpUqtgk+yXqhZjUViBZ+LFqHuNShpJuX7fsQ3zBYC2uZnzRJP3iwNmhu4oeh2U
eu28N+zzmSHUnzqhaszY0eB1AoaAGtXHyy9YjHDY4TfDfMjM4SeXKzMgH80scCgL
cPMIcuPjyr9h6RT9FtxOcnllnnog+HLTuV6G2iM/CC8iMOEwi4rjhykY1H9r048T
4bRBXyMLg/7uY3LPyk0p8HIMPkwtlWnLQd/dPGMbMJq7hEu2I5Z9G2/+Jo3YH182
gaGY20QusmC2QM067IXXb3aytovGTVQsh1YDvGl8Z+fHdQNSzRp5wwSHJle729Z/
EBbiVAg6Ate5PLgMj293dZ32MKI0tQYSAKZyQQ3C41mAF9igYg0Va0sNRlZju8zY
0nbIPSiPJQ2FJqgkBMExzYZMAHJUJVoeWBpaDr3xCu92RViDjb45WtWP5xf8HRS/
1Xytx6bSlCRIgEoJv3zLC4yCsiUdHB4/SLFTs2xIpCgytJ8r1CU0kbBLrTi5zf/u
h0XilZgK8RoDkDo+OMaMlcNux2pAOfzdm1vr59yp3Fdw0yWkar/fw7Rbb6bqGrYd
JnqYhGxspmSKxbkF+X61Lpcc0RbnTVC0cKVY2ZxYJ/ADU7AapUSLhBAQ136+qP59
msxnfk+nB3HgTO5o7DXyGlt1QGKC9XHo31UEP5MZD8oNSHacDnBG2h6P9Thd+Me9
mxC+TNclQqcQgrQa3mw9PVt4pPdzielPO2I6c63gpgkuMEPbZU6+wW7ZqQYesPBI
htzQmT9molj0znQEsXWd2wh7uz6OgC8bX8PxHjlxPYlp3Ui5Q8R93ZQ73en785xa
yAvN6rSMdYp85Fz+ewYZKuytlH9Ns87zMa8x+KieX2lxrzUIQREnq07a3NfbzLf7
nG4AkPX2T/fPJRw5cl1DEqTU4Ta8vVsH3CB5B51XVMDqeihKBDoE1V+XrU/EJOZy
JauHwrFskqaJ6xAsinDHx5Ojw1un1K/5NDFji0yr1kJDi7pjc+9FQ079LafkTmfB
vz0jeKNO9p/vshkJ0kDGNRl0gGA+jr5gygQVwILAwKs6gGtRzmOYya5A8Vkkhx0L
awfrDubDd439p1mw+MJiF5lVGFQJikoN/iU5W3e2r/m5UGuYZ6ndggTu7UcLOKAb
qwn3bLfxG5KrRBx7yqx/Sm7VOBBxue5EAP8ss2BYgS7dROZgjyXUg+NDQPsGpVMS
2EUNd5e7hGkUGCF0+Bo2rK8D/rBMB6Ehyq8iO3gt7Bc7cJ9dkFHyG6y7E4NU2IvU
evkPDBrXsYl38QhfY3Nxwsi+ra3ObsOgZvplC4mUcXK3IUYV3JucT/19RQ9oxvYj
ukgjvl7lKcPZObhqxsxPuBgIQZTQuZHt9RSLN/23sVbnp94q6qKHk9ISnIjvX0yc
vNYtnz+OmaYhQizm0qDlBDdhXgP+y6so8ydCW7yFpFMPBtaED0d6BMLJ/qohSl1n
y0PEqRAbgUDEPRBGNj31/nCTSfR2QC4oQN/Jb4M9P0jaiRk8XfGNj2ZhPZkluAVg
4/w0XdSTuu+UT3aPf1hq+6Wowg5Kp0oo4TvaPLTXnJSH7PJW+Zt9JgqeDtwkhn+m
yMwVG4GO6qQFSUwVhphc5MXIvvMoZGpJkp5xdDg0Mdr5wAzNuUgIDjNCILTzI7sY
Du2OIK2Nv321TYyzD69JlXi4baRk+Ij3y7E8+s81p3XYaU9Zb2ny/KgEuO4vAqBw
hsPkjUhFmiSU/VjLiadWOBCdr/PNK3VfNH4ugAoxdFxhC+sM7BRHkVs5wBudS/6N
2fDwvPE+gdBBlu6cbJfxW+E4FT0+UP8fZDc2QnuCaJD4bbsn++psCZI/YzrIj9F5
gdI4V/9iTSV271rhXK4PmSc3FH1KKT/MVjrjHYe4Ul93mFAeAXmOX+h6jTNisWR7
3Ysv1FuVcOqC9zWe8uyGu9Ki+ITF2SvIVEzCeLtAaqmHVBa+lNwBQTn19u4/o6Qd
VIzQ6n7wONLUG9l4m7DpImj6l+h472cqnDs+3txAjXFIdInnGK76otR6aEOajzZr
29PTivXOmeAheZIVvjxC+TYspCy1awKsPWEBIvUO9BRQXCBEs10dYFtxNPpn1X7b
SYCLE8RMS9/WLOm+CZIRd2rVTow2V5irsqT5gN7DEcpcUPbq1nDioCNWoe6hgBcU
fovmEUi42Rwh8bVK8HJ250qSa1YwFOoBpaYdnMc8YNMqYqGpCTLtt8vUjvc4+nl+
K2liklHcFHK2ZryoktH6for4elwghziJKNwU6Oaem66uj7yoDV3mYwYtmmWT160U
bmJ0jNL9dNtklIgpqROe+vZuTbCNmYkSdRNMe9jhSB0nNTn0ADaeN5DvMFuNhIWm
uuWc0J5akwmPmmv7mggLfMpu9j4/yyJ7+wbfWFUJ29B/vUxdm3u8HrHbNpk7MH+5
K7b4upz+L6OSUFkCfOGhKgW9nn2iiH6EMs3JafagEAaP41WJApYIq9YAfNxtABiy
8imMTolJ91Vgwfwpq2Yi5JwjJs0kaqDDC7s3v031kaXXabOm0zMUHyU4kxPxKO+3
dWuRW8nBmVUSWQ5D15Dubg4OVRZc5sSkeK3sP12l8ZYKjU1TBsWrXd+1WUd+4b12
ZSdgbgXyEgGrDz3m6WDvxZW6/WzrUulzpc4F/gykb3iKDxxzSE2E8S4vhIOt0Osh
JudJ4w1mKvF9qUYlJdT+G8TyoHwDaOR2nPmSSguy+4netCYk5PPnkAZeSsFYedwe
QmaXjzlbMCTqlmOhTj62YYdrDGCLcbuS6rJMybWEYEy3kDDRgba+hoRPJKs0C7aY
nr2XTsnCt2naP1EbZ9CK+x41hgptLyRNK5gatq+S+Z4PGz2HDaaLnXYNkxnL3wB4
7OlHS+hKanyrjLtDeACBtUT5nhwx7OVNpbayCc/g0Gfk259O8Y9PsimfBevE3oSw
rTPfzAu5t3qeUe9BnPXYYSpwMApXtok0yrOhC112JzDbazu0pH5ND8Wk+OWhOJih
CIIiEA6uJT8WJ4DPk9eKdmetJlgcO5eWzKuoiczSnjTTrm+a2B7LJ2U0EAjgRBnL
1XwI07YYglNgdifGOywuINvNE0FUWp8yX2wt665RcQ3qKyP4VAjw65vEwvZ88Z/i
IeeC2VP1vZmZWTeNYdoujUhwnr+0bn3M7TLAtnDs5qpptXiAtCXMXY+tMJlxiGBD
sABkrlt65nnycIlQRcX0eURnE1iJ5za7FaSWpi1+j8VC7qQXaU4dmGhnDvSwoox6
0SsSBDToaDkkixwesV0FtDp8HpOfSZA3TkSirsuPPJ3a/SKC9q/YUn6fQRPuCtu9
RqZ3cLuJXYEUbFjr0Xhgly0MmplkRwlqp9objG10QaRWPBb3s30OkN1fT00fltJc
iLDhK5f6AiSHRn6/IQTaSmY/h4tFxpfIhIUbNcBybaKcEOgyDYWX5E9UdopWcSTR
9kVZg7mCdNYGhiMqD7DvDMCQCeDCutX0otDxT5D9A7l3QHAHJD+yLNsExku0gOi+
uTYeoHtJe2lvELKvIlfcueuw2CAzteNIRohu7KqB+udHebm5CieR9RefZZ3ritPz
nOC1SJ34Xuq4X/xveBF4UOWTuJVtBaI/yixJvupqlRfX3Lc8bMWIt+l/24jetqtF
8UtdmoN+htKGu9g34v3VHAcdsjB7G4aOZJ4yLz4zdTyDLQlGI3Q/5lUXwWkLkFK4
o5TBuMa/791y3ekE4tffgXTsNdxWw0dv+y4ltJwJlMrSmH7qpjqYBtIQqkSDK3cX
nZHaMVtq54N/2asgzl14pJWYo+D/SBXLaK16BmDDXbje4lWHoHIfkpdOMWdxvog/
n4tHFjR2PK5NRyBUYjmWIyRidKCw+VYe7weP6asfqChbqet9NKca9w8fPwrgh7Ib
zT9eJ4Fn5zxR/95ghBnK7F5g384K/LWd1l8dY0KsrvY/L3ejly3qqXSheCRdb7vt
II5dgWC0ixun88rhhLNDKPKnF/cy7+H+oEhHcAKLlxobn10+ES3RswWB/S1kfcph
/jcikZmcECb89EGSsHyxYkasuCo4DoUx8Fb6kH0gaMP/a8YcW5to10cnFV0ZiejO
Pw1maHSMqYcjjdem+YT9kOAP5Ah8UsieRb/dEBTVBLeT/CqPUv9FK26yWbZjJ2Z6
Tzhf2hYI2RFAOa+EnILvb3UV4hTxJpupi91H5aBKoOdDtvBynoBhGmQpbqKm3r0X
BXMK/gtCkNEYgJRoUj9vQENLpT700KLBd9CldFn/mhtJbQhziEhO1MXosxhcZo2V
BtxVeZ7f1u/1yXcGeITRb2hRYlWCVogKL5bQ1dxdIEGIarfbSJDiv88N7gvhDy2t
Blp1qDuiv0dZemsnpdwQOEhKyR/B0nM3iPGpRZwNo1bz7dgR7tIeEPx3cwgJG/j5
9/eNJS2o6SS9NoGQdMce2sz21mOJZk/fImm2/EDcFBzl8v5d5lrnutUV/WDVnUHh
RYVq/2YmS8KHUKKNcilYXWYvVTJxRZAmERnHoEN3IUW9ozt1MH3Wcr3aDu6bgVad
d1ZPwCc0OkQNGioeCA6KCc0wk/oZC3RjgctyIJxzIAHLIrgbsezs3AWlRPeJScEN
uwv6nZjisdiKC69Vcj5A+AEZ3jkhM23e7Er7h8wVVICtaG5QPACL68pCYwa6Fomn
XtNNgPIjBi5jSSp3Y1vcg7Az+36vPn+o1OF/W9IUoDcd37OaVVo66zjJgLLzdOXr
O97xHlVCtumA/Jl5KI4KkyYYOzZg3yhMzNRbg0/dMFwe7/SEAqH1YHD8tME88wXs
JfkoSuubTFlHi+T/l4SJKGpHYAegOFDMkW3+BAyXlZS0Zmoc9InrxLvQqXgoeslE
M5D2a9IAoRFCddjNzVbuhh9+P2pTv6+tQUFMi6rd6tTMQvhKZ1R/Vd4ceMHmRNrn
0gqbqCmuMrW7FpvbBuzJOupWjwE1/WLMJbThwn6Pfh1uGvYy9KygVzcPA0BBy36f
81YnPH2qfvba01RMOyD8qTLpIVCU6VOPuhYHFIdWghSLfUUdkY7xsKieZSR6/A7C
M5srdIQoTq9tAaAeUNqJNw1QsctYWO6fmU1Wjk/TUZuBWyKCriFraV2EGpS1RRZ2
NCpNPVGNlKpFQYa8umbMvNrd00qtbyVTPRsHnH8NfXYTWTUIrcj37XytGAdEBfoe
Q0FYINYhqjSOKY3argyIXovrurnexCLST9QAlj1DCTczLuyn0YwedYb+7SgY8EEX
lkYSnF1izdL51pOPyAiLGfuW/mUSDUBdxPS3cWZts2aU54z7FU/XvQywIdwScgDe
CFEv+24ai4J3Dz4jpP9NHqf/7s3zbTfPs9THs+HE8T/AIKlNGa2eloRCPsuijGeS
SD4ArotWuujPfLwqZJd+kO3on+GteJ5mgn2efvY0EsU9m7y/65LI2yzQXtvlifXE
vV5QuSOoP2Mswh6edbU6x/oC6d3EBVJgUU5blM43Jf/eX6SPUfnDnibAfQBu4DyF
9A7ai/AxJWvnzXiIpYXihYmcB4VVr44JFGLo8GOCxhID5uWFdHCq0IudV3VRY7vN
nqg8cx574JNZDUoIBxKYu+fEk2ykEqBqLc6DY+bqoexeM7lNIZ8a+kRU+FbsKHLl
rKdT2HE3RE8YNbmV8ndjbrVtBzveBYmZkUC55D5l91Ke/mHb32JqYJNWSbbe0Lc3
RBjCHYsHmn2vbp92gbbhWlkaU9Vpxs3oMmSm8OlhoOEWGxgGfqPJoY8t58kZZASG
ffcaEK7dCNfLJqbY8CTk5fFbNWH0RGCIpiO72HxLf8lE/jsX/xqXerhjNGzQdeQ9
7nuEdEQkLY93u1hB2IMXPQWQO6lnb1sKBJ+/m51cPx/ggPEK7lKy69jaRjP1vJwl
vh1WOOej3LFspOnfebd+U3go/MCSsNIbsYFCSOMC3v/gJliTMAxPiDuii4CGTqqL
VYaQro1H8Ds4ckNJaQSvUkWqaVpxb/EirdotG3BAXzEgSHkBrV6PcblL11xvui04
qIZWo+LKVOZ+9yUvnKaS2QwMF4b7QnS4gP8KGWkcUXB03SxewnltkPkcbrEkhgss
W5Zepvv+QSSlwId3TBzSFLGXtibjMvYzK82nGsNZgA+1WWTWm3WtvCG8jnFGrj0Q
8stYwAPEarrdYIiRFLbTja6D5e8FEY3LJfiKA+mu8SL1OpRzbSs+hgB1e+TDgrIQ
PskyHYD2XMt/oLHkVqe7XUeUCADkMrhu43ISco5587nAtBgYCuFPlSVBioHcVXA4
Rs10WqI5jSQ5DLZNIgL/Txhp53a0OigyxmFlFk3g7x1GVp+i/Bxwv5maAvefWElR
rXdWknnDE+zJKr2+QlM65QrCv/nZODjE7SYosPywyVl41c71Pndz5OKIuQDWvP2N
Rsly1irD5tLdG7haSVm1sBDVBKvC4k7eEyHiYbi14OpT/Mu3g9tKsf/CdeGiFhK8
tR1OfeAXQDQirY76vWhffaFrbf0ZDGSRn/sOb77eBjwXiYHdCuyg7jZsXr4UII4b
0QoPx/4Zk2SFOJN7poyY4H8G+6IRYDriMsBXPmgbuCSYSwCk9Xn/kjUCQoapmfya
6IttX/csXAYm/HSWVyOEFMEKgJy5BgHOfLnojQIugORYQh5gCLVZNSgMCDOtk9z5
EWI9pqz7vW5Ivqzw5pPlvXUvA/hUt1E5HrFFUSPI6CtBb/uQwUiNqs4qtoTxkagI
FgLMAoPsdX8oHzf76Kxz0G1h10JC3UzgVSC9O8VDko1+z0g8Kbk9TGnmUVNK09UG
uQrKun3HP7aZjOi15DLBAG6NqdD+PH3H9c07nZ+fWIDHtpfI33lnIqoeZj3aYgyv
wZRZb5JNJJfPqkoQ4DLRKQKC3aAVmQYtXeewaRgWIsWL4wGpm0IlKJvvjZFVfrmR
s0Y6NCVZ9/HWv0RJcmjf2WoeUDYQMZrpb9Gxd/1jU80MpU44OjZPkZiSS21D6fLp
A7HK52Rs1bwu152vygkIixTtJ50g9IjThhUNTxE2CC/GMnbPcKyvVv/0Y3hlfs7w
zNW0vdUar0uq4JAp9FHwM7J/DzUfI12lQG2RMkMjVDRl+VG8wJPkBx8+ezn87/d4
sJseQQakXW1hN0cCquCFNxzuHR5P/ESP6gDzbC/NSG3LOJrDsFVyQiWGCMT7/quz
PGdr8XaywoN9GQ90zUNpqz0SLkjzgooR+wGQsV2ezywS01fcGSNJGclqpG1Wnd4i
ksnkUXdCntbVzOTrsrxKUgWc4mxGPxPxbAzHfv9c1HkLEMr3XyTJ1C1vkk/VD7pW
LVPKjI0FY8Def6gXXa76AOO65GYbu4YvrrlNqgTq1ar6A/bDb6Z+4wjPjRp7iU5j
5WGrl54pJuHBrpCN41TzKJZaMXBmL25VD5zdspDB2PwBS5d/AlxcqsN/zXGa8dgw
Gqf3l4cHHWMFpF5NQcj9sAoeq3I93ZnWSewXWtlo4bZQ42tPilZUmQKSb6kSgplT
cQYcqZzW0Zr3kUOMfsQD4wJTP7d38/ztlSoGhnbbhc0Z7Y1639shq4d4Oa1EBULl
uRX7DaJkUH2o0ud9A5DMWwCNeCQD1ldvIwpgMaxlK2PmG/YVnmS75jdBAQVcRV2B
ah7LScltzpZm8wlCRIRxAHsSgTt+015u1sRBylRrhIULIqNRavfiqAGO+hSVdWMu
99dTELsUc4oB18MqTaH0GpY3jXOrbczjpwRGAPKM/EaK/qzrgIW8WSzH9c2K1Qtr
R9Trd+wtgZ1Sv/t/6+ayE8k0eunTiO4xnQoleaAcUQLw5p36EF1aH9puKueZXUPN
StOSaD1h4OtVnMoZKeCPbofb9deq5jKN1GURoGTP/mkHK9k8aBOPh9oiMiZN50nN
bQUBYrqS6Af9Dh411kYOtkYOXmLp9Q0mvfL1Gtx1Zcp5FCdoq25QvcTIQcUjH4jU
GNUk4JCqwJrnnOO4XfnAhVN6XtIFSWCph6nn6yxaRCN378ELqd36HuL3Ml8j9BSi
v5jy2569WEDGUKOx/fQr6cuGn5cUnIKWzmMAeCXJ9ZrYuMfuFo0ENlvtV0l3mKVn
F2UGwazETIXYPqbMPdGGpFML9Yv+FbguHLWWO1EfeW0krsSLJ7KO0vjkFlya2Zo3
fSzc1T0PCkVDexZwA8njaSTrjNrZEZhM/clxrDP6ExVH+F2OYq+Sg8G+fj4inc9p
xy2munKhDNPbnAzDIN4yAQJs1Dcbi/cUbAz29T+S5wrXTGopkwucb55YQ0ewZgzS
JpnsfguEIKo2cqONclpAWmhQ2d1gWqbOxhllQjBCgkgujTDYIXLqgzumjRN1eDqK
sOYMnTY+nakWOpHeY1CLfes3yQmSfA+P+Um7IIfj1xMSI+2uU6qNTUD2knH9nlAm
zJ1tJi4CX1PBjkoUOVMJy0DU2ICgIEuV0VbxzhenwMM3RlWi4tRyScjZ3A8doOX0
sW9J3QOalPttYvdenM2kMgjnohG0YxXLcY2qhGQRTmWonWHHhVzR+JibG3WwCnkT
af+vbzTp6eEo3gZj8XZVp+iUziO1bQED7vWfjsciMztXRYX0sXmVkjjD9YuGY/M5
vFprDbd6dVEztP17SqwpjrGYq5jrds/RFD/C5uQZmCU3t5d2DMytiZ59Sfquutja
4E1t+4AJmwPRb2poUWZxX77vc5mKfCk5bc5YWJ6lo1cKkX95cpNhl+d80MIP3vc1
xg9V2ltYnwckWMH9jtRVZP2uUcxhdSufhlIj38Z/HHcrOhOQzbxy+1Nqnr11tpPM
YZyWzAltM8Cp7dao1ed9jiMK8ZceCbg5kNRpmhQ+wCjN4U/NoTYSaTj1eX9DN0wL
8fcq5rfo4LDwLMVwDf6x7uXXwfI1xbzjpR6uKYBw6foCQBBdlY2zyIvmFziG5P86
gDWNn0XFk1mG/hXmfkBkwsIn30D/wPt4oX4lo9JWmdlzgcJjwN20KZUDxoA5cauc
als/ZwWcwTf8OK9rT80OOY7qiY9lrV6llC++fh+1HK/9fTuMrism0Amtzi8J3vcO
dwhism4Q4OzCzDifVvLhIsdQpw8r0ewnr4v5pxv+00XBDCcdOn8AJnyfkYealv00
sCbo0tWDK7LTNqNQ2m58KMGqc/zgh/re8mePnCBhDQx53nMi9M8o+D3ahIDI3sJF
hASiUY35ncbwlUmR1VEZ8aJksaQwpXOQSvVXU1MS/EKLfCSkVPJZu3aOKTe03t7P
v0bRKqo+JGQTsGb8SMOYYjiOcjUtbG5nFcQSp+ad+sCmOnZdDDeQmtGjm261mg0x
9GUK+MdLTlviwa5MtIQII6qgsvdeEjs2GncTHZLXtc7Mf9bBcO4NlvZ1uVXNuDtz
bMS236WpaVzdBrcTbaUVa2oYj/1WRTM/FC2GUgDvKAGypEw2QgpP/m6zwNvlMg3w
uSTnaZmK4QEjARKI/zIa5KvlMRO5MrThmuLjQXrUHpJto+8vkpOo8ovPVbDpK2pO
iyMgDncBENVXKyt43XWvZye/mXHekxOjr9yN/SJxAvk94DkxJ1i7CSSQymY6du3R
PS/5qJcJ4O5XHuN/N3Do1naRO56IWQSSMQnzK2g8Vfv2hpDM8dpjBp8i4//vsPMy
6kHxkFm2jOqjB+tZuoyGVe7wFdNhqp8maETbB3pyFxdjFjUf5YgaFriMTpuOhGvg
yDmcIb5LK8VFmZOwrDpWyDrNlQ9uf1OXibLtDO4kdC5cquD31Yg+CIBRSeA1zvE/
Su7DufS+IdzgjLoXnJjqXPel6uPCqI+aWveavoiTTkx3yw9BwUnaTXr6xGCijMNI
MqlRqjpZT8rj6HxbVDiH0D3UV8x7ew5rGYD1YWQ2yq+O7/uINJ8nGBjv0gYCYLQ/
YY5GWEeugQbCsjR+w0a0ypg07GzdT/hg3BjIo8Gk5qLxoSyFhAw8CupTcPyP4T4z
vp9MeuyzxmEvmvOWh91r5/zYwM8Dm5mcoHPt9/YJ3iFz1fYr6pzf8YBl1psnl+Si
DiJgY3iHe6F32vlupZISrDUl+BHhHWV+XXrFoAqn2ysr3fb+15lQFczRXLscT65/
DJ0R4yca/AVyO/OGBnZrrWM3t/F8gfwfPcNagfUOXBS2F8U0mYimSe/W/talYub4
ysKRxeA9gBywUg+Wh1+45ysXgyxbv0FuqDVOKCgRkrm8z/apJKpXXOyQhYfR4bBL
z/dUSPioykZ471SqN75YquPtnEpnJ6pJXYqLsauq2skZaNVRyQ/RxTl+IPdyFaPs
c8LJeqmbBLgcEKFbtuxz7jNljP96bB31dKSVKmPSrzCa79iuzPfy/mZ71dRUJvjK
5cFaj7qX0p5p1l8XPw7DZ5H97zfBH6061WjB8h4aJJz3LafXT9r7ZX2NQL8tm/Uu
AbwD7Wh3dqNWZzcUxlj8yle3SodZRSzIzaeiF8yKKQRmeQKFeBeXYmkuzkxQQQrN
+mLnDviYbqXUGvgMViCCZV/WIgFo2ZobX/J9i35RIkkKH7MQ8jU1QPa8+6nfhws3
wW4SATRX7UCMTaHC373zIv5hfkKLUSP0RAFvQ3u+RrmJTt+1yChIpIvEW3Ekv2Kp
BptrrT/VA9aG3KWvnmK6I2AKVPY/wCPgontJO4OO1VH655v1K0K5liK4hqug8LFY
NFRr1e1zh7+6pMP3+ESVWmBli4n7smFlwknn+z3FefGmwub4IeavzA/EORz6u+Wb
wsWzHrnai61tLgjnU47PyyzvnX5ZlCM2WgL/zjvTi4+NJaVUA5NdkUnRq4wcoC3y
bXmwEe/6F2JNzsWsN8BZe6CKXtR2FF//cQvqSoOxgaxTyTVgVcSlGvQ7Mcf+ohkE
pjWu/eD1e+75Z8TPrvA2oMeEzW4zJHxZEvNL2LRGaFotdG2EKKM/A91uVCaNBlMr
DEU4TaqPVFPLWXM1f6ULrAktLgaogWGozfmkIbxc9z+3/4+BUtM0uS+E9B8DLKdD
+ixaYjKGVNI/5VgYqrk1dzwx12BoTLsUUwzk4MOa/EfDP7autRIXqHuzTTzPp1nk
Hu0b260YAQvjpsb/XiKTpOQ70B+BBYPZnivkqwRok8BhuiI70wcNB5GUjP6+gmAA
CeulLPM4EEkiQiTaiAZvxixg7J4rN1ir5nKQgkVsScqpsjHy3SP0XemOtgDcs9lP
n/7B/7XZhas1dRKIYaLD66WXvkW224sPoOuOYbAZcmPn5hTDDz6CIzH1XolMFQyq
izFGroWB2U/MYQwUllKAQbb5coRKVwYN+HvOtpOtoVgEr5bgM8Yvw1MosetJimXW
pXuGOh+CQJ9fWhOOeVGar5G5uoQVJIYmmrc0bClrk8GlDL1icuiGmAjIN1LQoQqs
kqfMwR2l8qwIZgN2GyEsE/cn1Tmo+A6dF7m1nWm7fgsb2dmILjHuGifKcZ2ih23Q
U1iVZVbbZsuYyX+O3HiAfNVktc7ySe588/Y/0mTJFyHucqhRTgl5702bSTWts8vY
cd3a7+jR2Is4GS9BMdkEM0JY9Fu6XlTULGK9XtO3P1kzrvoXeHFOKWB3MpGeVo6R
pAXfpsCnCulAqjsJpd/6PuvGkzQVsZogO5Lhmbog01ZRWyK6NsMTxqqadPH0Cosy
kzn9+S+pFrVabfl/TXlPz16B/qiilcgN+Pa5NI9frcKc0feDULiat2wh2cPZ5BUd
CWyLiP9+dU64hf0/JkWA7DAwVoguigEysgkyJ2UK3ztuySb8sFCsRt+VIsc+6xg1
zd0v+pvK8+wCynzDH+zVEMqzOUO14O+fpAbNMCR8eLg8x3dqTJHIQ1bJejhzS+ST
Lqp4i4tZElKNPyvXuFDd8LrXz3+S7wab+7gvNURO1tYdNlF/Jpedl+hrPpB3WhDg
Up6gjnHfF6DyEYglmgLQ2o2ySj3VauaGMGQSHm34zbeDSZXyh/fWV5jxvDopVO8U
QxNqH7FHbZWFRFhqfOT/Zg5GGk1QTvtAUlYTtPi3+o5vi+l4z8I1lP/CdnMcEXLv
m2jMOkiHAFWq6XyfTmmM/pr3ZpTWSlzxAM3BMNAYojQMW3wLC7TCOjBdmKlIqYbS
0SZrcPkdvjiiKUnjBaHDX1nWZeEGwp1B/6V5CltvphdU2IHifXFYIBOfYmRavU/U
EasyXWPa6gXZGmtotXrQAJ5QttkCCkh9RGnWzAl6aFub7gLF5XLAzfOpjuO+FlJ6
C4ZFsVh1BGsOW2MyCkJgNlrN8gdJnX0JxfG+bwuf9sR7wKDHW7UeqWtnEffTiefA
lAMO9c5OpukQAxAITmsdYXKEHXoEP/Zu3NhksGH4w4bO/s5DyxG+fEYnITZloNp5
vdS5D+0AL8q74buZH4Z728jcTKyTtJiBMFuFYTLeNyuGcKEjPr1gskn6TPGS0k6e
+Z9zWMM/QvultPkXnu9wlKyFyrok2E1ACYkPNSrNZ39jQz2EfrpXjWlsye/jpYKs
ysqgk/SqjM7WhVByKzk89Ywv4/5wJFdEjVR/HBgdd4buG146q4z/zA0ucUm3XkZw
wIGSksD+qUrLFp5foz00s2EZrnKoUiyF2Bd3DyYWT3rbGmy1gX1d9vP9aiZ6zL3p
bglatXHhhHgET35MPU5byP0tLfWS6aAQPr95aAM5RENJ0zInbz5OE0Qa9Q9hcO6c
/tBtwU+KdvAfO3C4z3q7aTTQAAnrt53HEkZG15Ej32xILQir/HKNXsw6NnH+X4s2
TjRgvEJb8MgaEAMWrpmDLikx4rwecScVMyhG56dfcZSqlJKjDn7f5Wi5h/Abpfnj
LSUuKXC1AnCBaTpp5G9pNCna2RApdki26f1M1BwmWkBvsp0NByCMrlOY82HLHhxN
n2HllHOz1fg7Pfq+Hz/RoV4iUnjGdUl8J08fGb3ZgZKLTjWQSbiQOHS6Chn7fiGp
EZaW34moMLqyrf9AOCw6vDxIP3U/e+YAP8U24JLGBgRj59dc6K74pCBrN2TVTRqL
WmDOybDhhVKKYo8UFXo33rIZEV1K4EAvbwjno1GJcf0i4UNApdZbP4gSDfQtTohy
h92BWewvTh3dBnqBLdzfY5EQb4oXny8k1tO2oSu9wOULnsT1dq5mjv5XV6r7qgP/
KO/gMNEBrX14EH/NehzEX2Dcy+Y5tMjoGEyXb3vY2jVbwP+6QQCKbR3KetTPXw5F
fQQ6sYbWN8Jc1xtDcMCRPPyr5dMxDPvXhMXB2Ce32eOOf90/P9/50Z4tKCrLBsBN
n1Zm3pp1WMmPk/+iUcq/F9JoTWkKhmup+479DjRi5c+LahXFI5Aa72HCTCeYYrmU
ToM/eqcmK304ZrCmTagXbL0Pk3nKCcI6hqt2dqltee4ddzTV5E4z2kRtlQVRIB/b
yQRyH37M8/imjdhHAp/zea//FVtuIGV+3eUUSHYANhK+NRfF5ua9CDQc8FRtBwZZ
HsPai3XcAgYUGyON/2YWU543gSEyYPerZA6LNQcCmPU3Fr3k7W3V3itXlp/u4D6v
10MW7AslUJqmUYfqzvcyjEt2EVpDX/PjuNNnS8+ZehvxUjRO4RY3qTw4B8j2REL3
WdjqJ/06qEqihclEaOw6K/zWUKoMSV61KXt4eAjfk4d63HLjael6aOGe81TUMxOe
GYsLnTtayH/Edlj3TtnXqlSYc2NO/Azd1qBlgxZTobnkfS1M3g3DxVk+9cSasfc8
j2F9Lkg5pKApQ/0gNeKDf8jIQfGu3xFdaq0wlWC80XJlE4vTbS0a7ezaUNI/OEtQ
KOu5pMOrB9ZeiAOQPHjIMq7z9hueyUhaqy/4+qk0mL0+gb+/QqdzEQQDEom0xjF5
TL+kQMbi1t8Tj5ls/6NPet+S3brdrgDOPB1PdJYXKHKjUy1OSIDs+1cO1dshc6hV
UI9IcLF2hxlfIcv1/LZa3kFJb6GF9hxDwfh7jb+1r5W8ijpmMvuqbzgx4pGyFl+i
anrqnjUNpzjp8nGugyTdNrzoaFSeqkc1d25L2iUORBfijsDbFYI1p/HVQREDuxnK
4aRjpWdTj+iU03kJduPotbnwWaIdj6xUndCVNlJNY2HMlCyjXYw12xYOUo3kV4Jl
cyl1gEP75OWzHMe5dY5TrOGeYLNumH9nuGDDZo0OCqdNZd6WKt59LwaDAmnUKdJ9
/ULalkrfHrc+yVz5UQY5xdE5z5y3CtIA2wh8bvUXDbfjSe/9hkqhIWBy40CreklH
HVyGjtMzaWfToAs/9BCCs0fdLyILnpGDwuKLycDnQfdcQ38pWQSV+YJ+S0Y+VlTR
1ZLNUZlRBvNOHVgLDwDI5iCkn7TPOofNBXPk9fZnW44Q70/VSWLjt3nwrFHLi7/M
4ahhn4Q/o2L1oPlPIG0bq5rjme1swHXhIvUNaXh2BLN2zEuOE9JFJ077UFtoGwDK
p7q3nUH7fCXP7LHKKnOvrH7b+VkvxsTBB6o1pommVzUBuzmGyQ1LPQiV9lKptIQ6
Jme2BrxIdpUXNa5jAj8Xy4KEBXJrv88UEsmb0pX7FaaOQnAUQ1ix8lWW8RAC4AFF
VvPaCh8f2hgwz6/mmNw1cJx6XERosJpy4RhhoX8aeAiqEXjZHGJA2w3Iv+6KazI8
qOLWiv7YKdxkAy2td8tkrAXlv/nDW2Z/BTdwF73uu9dMy2W2QpDH5Cp1YpKaUvr/
m73qxLK+KOOqlGE+MPaN4KXBkdmI2ik5YFUBI8dFg7rdn08AQwBqtFiNeAa5oToI
XHII0VprPGHTeLFIt/SQG4okj4T35TsMFIZJ1b9A8E75g14hGZpMQVLJrTLI4khN
aDR/4Ton7nOIw8WZTH97jaavUgjC947SCJuNICHhWh38zIUCO5l51xQh8ydB/i7w
fBeSujmR5OVybd7OqCuc+qXO++JKXBAlRil7mYd3KydGPv0x+Jp/YHoMkbwL3Nsj
j3v7MsWCHSQDQKiXrgYV0YU376P22Yr5RL+xfP9+dweoz5cIMGPTP+PN7UCKqFVJ
Cdt9YDNJ9uP6NEnuQYXj9V1Qfawy9qTwE5KaWoq3WDe2VmNE6gIJHHSnoxMVRj8a
lUOHZX9RYLxY8hhNLy0inGA/TNhdbk0UiYAqdGIoi/N8PfaeKV8r9XIaI9UHnf1p
sKIeMm63pfVBNCnl2BptaEHOQbVzix1Bt4JfUKSLkp29VQp7poAQmnv4qDanzVlD
Z0OQ3sVM2k0cPxyB0Pum9Z5bz90NKKl+V+m9YX6Swb3hfTUQYm0VE2MdlkWgKPcM
gUuFPwnahhEiIUTsddShrwR6p5swEcn3mv1BriB2pTVs0SUXSigqRdZqj7tFGIjC
wFQ22aTZY1GIvX7ef6OI6UQiy/kTAjV7unWarV1bE7XlWkd7doH1+RtTUKiAMV+N
bpjrr7bjO6T2xlncQdddxHPugYVBwoNUeRHauG3rFceR/6nj9U7Ncs3Y1ftd0zlX
m1uxUh2kKK2vWkOSsldJAsqEcu9R+Rl0/37urraAd+2UCBxzar7CKMqrpUh5qkbg
uQAfpEcbS/YjCHXfyvgAKWng1+IAsdeXINbDf/h8aDv27ClC1lrOORsfhlBA7mN+
uyk9+XJAqc2ARN5nk8iMzmOUejm/M2ADwpGVU1Y+i6UV34+ucqI2UADqgXpRNNny
lm/KhIN/YlgHh6oxhu/fg+Qqn/sCD9P8rnNloDc+UOA5NQHxFPb8nmPSNf3uX5X0
EhqWwAjlE1gmbxQulZeaYBaiZUJgyV0VH86SbdCC1GU=
`protect END_PROTECTED
