`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NxUuqzUvh/5o7YZQJHlPnWjX9tfnhY79wX028Ig5caMRbyow08iFpSNueOYgyQo9
d0OjyoyOqqHlO2XtQPh6fUlt0HNK6HH+FloIZnZpevIVKADEDJcvQWlP+jsGD9Zn
l6UvaLhJ5zlYdCg/bHggV6aYmAXF7nZnmZyluQq5FPZ9Ul1FtABEz02z1z0NOEtH
DnXEgbtsGAdCqiu1mrrKXdHvlN1hKSyS/bt8ehjPoS8aNhE6nmMLndgzOCm1kRj1
0bp790VdxSnc0MZObXDICCk0KUG03JqHadXhR158nGOQhzISrTjDzGOtIBHak5FJ
gCCrP1BZHzeyo8nCgtfkShm76t7CuUusQ/mmGfbmrr5ZoxErswPjyL4nm5e3Zkph
Q+Nh9jroCVso5GPm/kQo6jN2+Rmwspka4Am1KJQyxJPgE7HajZT6gc/ujCG+jQq1
j5TeEYkouqPUmUvwCAJFdLmyY2c6lll46LEKnE6WfazFHyvgw/N6lKNMCzYBzSz1
3oNWvokRtUDWHqzFy4zpfrDuAQitDVDKZDZHHuZavsxVsqfMG3txM7U58i4sMq+n
88cyEnV3HP2TiQ6QBPenAFKhnFWxyMvfmZqHy5fODareCUOa1wMbnPue/TmUdH/3
om6luDNrnl2/yfRVD47OPhtgNB5HKkfb/zJs5aLkapGeg0BQUZmA44sKkzDoXPAE
rzTNWoL5GemZBliB4C3sEM14Cf/GMQMd7/EZkU/zn5qIsYrGhQNmRb2ZeOn65cCJ
hYJN0/xcPOv2YT6O3G/sD/m+Fw6ctD5xnbhD/xm7OuzCZ9jmOkyecFziL72qNdiE
g/lljQhlMVkhwp0+qG5RcGo0zlpcniL6JwVZA/3IUJKv7LL14oTlrzgbw3SsDQ+n
oYePFo0AY8mjI5BKwd9a0PBolO25x7j2FdV2cLrGfmQ++3pcjg+0Atr4TMuzt8Qg
RkE29wGecr49qlkThxoknOLnBNzPlvUk6OBbp6zF4egNwE14r2mDBQ+sMj1p2/Hj
9JbWnRkm3OBICDb/0j3ENmMz8gQlF6FGOLjtn4bJ1ZNWr9HZdby9S+Lbw1shnP/R
2p/iVs88Qv7qa4S59qAo0EUixhSMokz5W9ALsTXuEmXGPSEquG+oiNhbs9gZaBcE
osDLCO9i2diD+dIX3vqaMN6Dtjrd8sVnwbwXuJzPFxus4JN7nryTApnFWz5h3RMO
d8+HfQ1ndBpTrBvqqQ9KrmulSeXqxCSHk0W6SNe7P+Mpid5Br6lBiDkQV42eZy2z
RmLGsn0rgRLkNVwJXyNQDOX4Jg5nIYStAamYLqujOjZ67M8ITDs9woiKpg9aPHZT
Himz9HM/ied6YBtmdlHO3VFWR2E6F/Ez3YXeymw5jIuOaeeCd+pa4LJBdsTVV5k3
J01I0h9799qJhR2UKTuSQJP23QxdDoxjThLpsi82CiZvmQ9dSSK050MB231Myg7e
eUV9IUsgOuw2NMKa9yc6RHpBa9SM4LS8tRWcCJRXhlOjm2dUCH1dZGARtJj27Bjh
`protect END_PROTECTED
