`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xm9u8Op0rLs+3VdHE7IqMpuBwPh3feA16NMjQYpnxbi2EyLgTdpoLm1Zfa7XDZ6o
y2ISXVViRjbUlS47TuVsDFK6DAP3nvQAAkI85aLUxUoApCJ77EvKU5e6hKxjZXU4
MOSBXtAIgL5Ygl/rA2xJJF47vGFfJECsHcVJWD4EQgLlXh0nLWtunSMDsQ8iwJUc
G/J/6IyQW+ktP1+LCKbETYdu+ROyQVbbOeZ1B42oLlpjkX1kCTjMaH0gdPipHx8N
pCALIyGcbwPfaLHqkGOBxoFEfAqQuxeLGeBsaEhnhnCgdO5Jg5l56GbxAoYPtSxr
zpcDiL/ygCAZ2hrpOZSKIL+WvHE3TIVZwxTF5KC/JqmFcqIRGMgZhp+71p+M4wdb
mxIR2fd73M2sQaE9AWy3X2y5x/AcGy3DdCc0CO/ZdUSV8eLtgfx5E2zvmJmbZnwd
ZRs4Pk3eQHBt0Hx7ns9OVnHpeuB8lMj5Z+OKm7ZCK6YaSotDw66O7i+rAY+PjVfs
aR/Z/zIFw+o4xwQy5bF7pmysVLtr6NkJff4kh/xfZmz7o/SFH2VSCeVNC9dcuLlp
U8c56EikF8rmOdlRUmtRyM1FsQY2g04P1K1wAD63bz93Afn6Pp/J5eWznau885z0
7paPoosfOkrW1wk/JbIE7+6S24aAf8366PEIhxpVPVgRhKZR4ctWB9iXVV82m8pI
x40AelGpEpgIAJ/exDKYwRLlVQu95eShYot5BC3voUieIOk56fw+07/XXJqqCH7+
fbRmlK5MUsBSDwU1gnPHZl2Pe0gez8P2jSDWCGBOy91+a5A13si7uXnCsyJlpkc9
4/aZrf+vYv6e8N7JzW1B9ISYoUeU6f6yWcGjlBzorb5cbIyowrijptUJHJtm0+WN
lQS0YfcevqqJYG/guGFRhy0qPdBaWcVTbWzXTqFSGf4OIWJ1GilfPEziUU1jwhBG
MqOlAyOo2ylry4RtsQSi6NjV9aT7ZaWtUH9upeZrGLrOtq7XBwfu5qzw4Drk3dkj
tiAfw4RZK9LCpM4hEuz/MU72cDCvGeLLzvURaDpRT5XxlEUNzmErPj8Q/bQLk3jW
iP9frKjR57q8MY2Mx9TysaFv+MiMWQ1SlHItDsgtR8Lhddm7pQg1fRC37TjuqxHq
9QV+OWL9v3x1hydeqlBl+NqA2PvxyX5HIilIPmC0OgfBql9vTAw6xktGc/4LY029
eDd61Xx0OjHqiIJ0ChVv2IYWgBE1P+fNy2H9+5SeUOugFyaIJTpvSmwN/BQrTWg2
cAuPKNHVp2D0g5O7gNz2dhO6aXtKQRYq9F/vIoBLUU8i9BYpq/9mJCpQObOB/kJE
6oPN0eaNeskeFQZ5JqESDOQ6/l0WNWWU+xZzdE0BOcowZhVQaoKqHy4K0A4x+Yp2
nagBG8yykMCw+D3n1EoUk5/Q2HV94fxQytlRguwt/NahS7gjMfV/7JbNLHTo7TtV
BcEpnhD9VTUcTV8uQYKcKO6WUW+a5dYSO5miSJd0XixAarWedKJKDYFN4Xj7IucQ
Qw36/xrWVdVj8vd5872tbKGrkFX6Z+VWp3Tr350BZOvmbIJFVgrpGKkrl03kOOBD
J11fICMwDoTiL58LrYdz6e9PbmFYsKgyUlq07XwTKH+h6V/jBBs7uvzZkbWJp079
j0RhB+jB8K61o26/FPlCx7lkKXPViBrFceNQ7Bqiu1VomDnjNYdR6x/BuVY35S3V
fhbHd7MJliwLH60E4sSYTfpN4c7yDJ9lMXitfSxQY7uzh0LU/LAdGS67JybwEDvX
9hPcMbG45sl+4JsK/KRLx73SSvPbUGYzhwDiHbxTY729oJjIgi4zUaniTEUNhBpq
1I0PSpGl/GaFiv0e5LsVUNm0yPzP3187l+twOMqk6TfWBAaUpu3MAJIQ3AZapkb8
+Eq3GcfZ3gz0xfByo3fHjxE8QWLEr4CaBPBDstxHvy3goAoXYondQlahDyInFrQp
4HINVry3ZqGyR22oN7PdJtyvFRLFYE2KbzeOb+iZdPYhNDhwiQ0AK9EjMBf6IImi
4GiJeHDEe/2DMIJ9YhkUyLQpUDdpfcQg70WLFAKY7/H8dVCRDA9GF2gmihYVB8hr
QEpaPabEg3YG3crgw0Y/QkMKkkzSoC0E5o4DPfaQArkPfXfaW0Xy+KXFSj2YiDZ+
bE1Nxrrx4Rv5gkk8HSy6BukMpRr53c49GAMQe9Ba4MDwyNNxeTpZExNS7RJvwdaT
YX0c5RZfXTpPQS/m4zyovNs4bokWl342J77qTxs0G0aLKGtrkZyc8BdhEAq3QXRJ
BDVT1EAz44REWblQ66f2INd68XTdSQdquFB/FwQfKSEMcFik6T6G5513H9eNuaJh
KCPEnlY23LScT/8V55BnxUwDU81zS2XEbfzssCxP3iePJA8WxbtHYJ90hxG/vWp5
qQKqcEzlcpkHZAtWCCLmmxyoZifuTRJ61e1Enxw7HbdDYAazb1gfX/H65S2vt7oC
vzI5lvgynmL+82R2Xc/POTJjWuHAVhlqJ3xfbjS9722CI6Wit8TJ+R1/kTAVcoBG
`protect END_PROTECTED
