`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ki/ExBwagPLR6Al37iIvbC2kCnG9h5zI8/R45NZjIicVHk1guJVkttuHxvb56hw
9lLoYlf26paX85aBP6Op/le4MJYGDkKtW4hEwJoEbz0pHJLq81jTHgLAZ2BCooC6
9TbcSJ9vcMUcqxq9whSzc1oSkEsmKaKFawTpjSFjTJsdr/IBedhIZxi3yxqvObRQ
wEA0YaZXujvUSvNubqNvXnH0EOuInWq+gp6Y5rwqEZ5+0bZCFYU9I+niURXN9w3x
32bkAefKYKNtV/1Dj24MKLS6ScIDvM0RFrDtBCOx6THrp3q+JPTD7Ij7maN9q/SD
/5KpIhciFRKij2iUwo28lNGIYG0XJ14HwpTgmTS1Kg7xmAvjx3dMjy2JOD1bcYLK
`protect END_PROTECTED
