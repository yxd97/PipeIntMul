`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G60VjcHfbTQB86f0idVvG3+TFwdez9EC822uJe3TA37kEjxJW36LSXv3KYiN+J/+
5iQoLPfJGVnqMHio8rKoKGhs2m/0Jo6I2zsSKqAXIaN/0Dqk0hydvmpTUqOxLmnf
bSMz9XhlQSRLQnY+Kv1hky1Xrz6eAef2LUieVAo7bVJ2px4o5fodtmpe1kvkb5t1
AE68XiELdL4z+gq4vSaVunEQl/Kn7SyAL/c8K7PHKJjObSncSGGdWR6uGhTWeF/J
mBIH576CtsVy9ENdFETjq1v/7G7TqUlkft3Nj8cIvQmiiqfGAKmTmOWD8D5+B9DA
MDOb0pyQzFnPf3LzvKNotr87UWH0Ij46ePlUnl2xAzAtmEYfii7h9wsCiULlvvll
bQ0Q5+WZil9SzIhBZHlQs4Q8kKpmVcYVnHMlMZQZxO3fSH926X3hkbb07uASeopH
j4U/XZu6++B45BMI31o5UGjqQZOpXXqxuePWSZL0y9elPEFxfDqky049DjI1H/mq
dZZOkJaElsciHklhYF+fO7QKBipDY2C1Fbd3cMwU3mTxDNUyyY6A8X8r2FhUK4XJ
alnc6UQMELDTq9/5mkgxl0c92wEefjHP6ogWHoLhVnr/xJbc+Kw0Mpy0wauvepNy
OPqSs9R6Z5GtvyadQkLp+0cNZjzoXnjuFMnkOyKRmH24iOs/nE4kEo5HvOJPt+cv
wG0NKOCMsz1wtr+t1bZhT2KZM2e+34gOyao19DrB7n0lztzN3LU7mJxJ1YyPSy5F
fRwQC9eoSeAuFJ4kZ/EXdOyCuOYTOwaiqI2ZVXU8XjMxZFdEXRm1TaUhgaoJkN9q
bX8MUAu9BlC56LFTV+NjqgiTK/tbz/GkkYxRXbmOrZELvQjGnUXb7mkMJ/nF23WQ
HZPNYe/Roqwnrd192ddOZLGgLjaFp8oNNKJxXoUcpK4k2VvOfBfaVMDu4keYF5Sz
m9xDA1MFA/bOKST4SuIJTLhG7Tb02WH2gyIz3TtP3TH7TpCIqtupe9k923v+VzMi
J8W7SeJpOuU2WkCrbNeyIY1ChzxT8f+UTUIhP7S9sL7i/V2OASuFkrUCo8RyczEE
IjRNPAKNo/+s4qkbkXmczwTGeA1Ea94oDtFtUCo/afdn447bpqycJrCC3jR/Z9eO
3y/hEmotlgqvpe0ijLTkcMyeSJBXFSetHqz7EWS3sm1HzNI+v2qUluwu5urMt1me
c94hEPp2/DLMsDWWXbjkQaY8gaoEiLOtnnpE2px7GECrOA99otQ6ulHbheM4bk+l
7jWQz97L3VvgU9qcDFeua0qpXoxFahd3eFwRPazNNazAP+La3Yj8Sz5WlDkEwAlL
id0NnTddK20130EbwCk5/V1JElGXS7dCU2Kww7qQMzV/+CqQI5wJiBJNooMI5VKS
NfRznbqBe2q3GbgZbXzFaMUxxCAEhlARlT41BHDgKYDX+NDWTueIpJM45KNuI7C5
Xa5bd0aIkQIDR83Qnv4NU6o4bbVoEmFFSOvPk0YhqLGztuJnHjgdTMCGGUsm4QTm
0s5du7XPPKBEd9AST2M4jbg7jDkoJD0kzvqyg9bt7gG4GcN0vsPVZ8hsXRS6t+K9
bvFTCIZ0vDXxfX+SCJclwahGiOsrSwpYUZ5HQUhdcHh8cLMSbmTZseXKy/ndMpHV
HGBJJSy5Wyo8vqX3qnd0yOFa5tdACivITqxvSHGIxzJWrweRTtbBAzecV7DOue6g
fd6AzQvyxfiLaZoGocqMQnstX+UrrfVCKIkEptoxX+b9SEXCUdV+xyhOrKiPSpxr
WpLx6EKGiXxqwAwWDdpY4YtY4M0W/AF6NwXx9JOshMhNl1cYoNdjR6x2BSPVwgyI
AQKKX3pv4MT0GX4g1ipmBgLt7P0qtqtxE8tb5HJ3TvkrN1qOrP/SckhSVchXRD0Z
a/qp6Jr8F6S1dIB/CQDh0SZ23VRdibnghS09Vwz+icbcI7yOoFPCx/AiKZr4zwz9
N0YTzAAz7ywwKCVYzRhOjpYWEL8RDnP4O08ZAl+OyyZltuc/Watn9uPxR7nsXBgP
rpd845Umy3XFd0jZ7dX2tDx591bAJ1UoI2auzr2VebRlKVOxaFtmGGF9cIjj/QCW
jCpBotPT3re34UnQ+T5cOFZ0SoOxfq9ssMWLFnrCAY/XnOyq44E0PfPkN03E/Eac
1QKKsi55dq/uPJWchaGx14mSvWkZF1VPqmVNRCzHNziEUCeC2pz933jYh+TPuTxO
lmOATy/hPmcZQLiWTi925+Mc/0LoxXFLsKyInXhKJBAyUB5bV04yW+AsoURk73zj
453o4Bbi8NKY/ehlmkwyjLrZmOTMoSLHYlHucp8d1mgSxVeWRmiNX/dAkWUQaNCt
pTiJ4J0xfRjPwcFajzl/luH2yiZO3iukTHno2homXZbWpgnTbO0KJJPLMspKDhXI
29QLhgZcmtxY3xA+wZ5STY0EBa2mI9X5KerFVsCj05Y0T9FV0J6go4JQk6R6xiV+
xLzpR7JlopBZTkuh5+rrt2KpD6VlgfGAjQ4QcX6PkrGevbxfbzZ2kulXuqulDfWo
i0xWUX+xbHXwNIMTo8P8tOBBLIEw+vkJ8fZMvPsFSbg03mKnt1jr+rUWMFKB4m4Z
Pl0aQ9leDLR2bzK8fJmb3+4rfyFdNEuq2t4GFwi+78H5iAuU4kpJrdmcVsakaXN9
ghxRTNCSbmp2yWipmoIly6Kj9sR5tQgRmlowwKfIrWP0KK1j0UimF5bPue/eyhwD
acSkJBHtqxpTPZmYXw5h0Icz5SNNxIAO3k7wJgzxoyRf8LirD2PgJx9jDfhlW+Ld
Xbtm00Q5WrEVkeJe5GmO2DPjtx0J1yE6otIz/8U1LegS7hj09VVXSg74zCJSVkE3
0PdpwKhILCZUAmjysijaImtldx8QYUgS+hn2+YgeCjB7ag/4Ph3fbv0Z3MLWiKwD
H3pvtyd68wNUVpupXInFR7iyKjjIr/Cgb/8dTsJqNytbxrsZk1Ml6EEAeE4TLjyc
UvCwsQ/VNpW0/XVrN3VYhYG19nkiAo9Ql9oZmKMbc9r3OZBwU/U359uX7Gm4o1BT
0I6zwDecJ9Sbyp4T+OxG/vn3+K7Qz2ZdkDj7X02UReMJwAizcoW9UhNawG0AmH6E
4RGqNFJuPtSJ7oxSOO5oGKLTlbXa824iC+lzZ0vBL8JXXM3oGDvk9mFRxBhnayZX
5CZLHYhFucrvX7UawJQ1cKwPcItLH+kZHDsxw0wSHaE62nP1q5IHHbudpH/T1HXy
dSuB7Jaq11XjXOwwRbvJYQWwGsWewxO8P+sI6aLsDz6AsNsWQUA6TAW+m6hZuf80
4sHYEFNfLLuYUTyT/t8Uc3qG1Pj3GHHA1tKacArmtuIt5SxzClfjHG/WK0VqMu4e
5FqVAJrAIhFwZ45euKavI/bXNRQyCm4rq+DG7bsKwKKUx3pThPl62k+gT80jwUCe
Iu/P9GcpnNJYPbtAlRPHiVGsCXgN8WVwhHWCrn23xpnJx0q4cAUiM/8KsqUXTwrA
AoL2OPewUBTrI8JtaY/z32aDcSCrMYx54GSSHyr2ybe3G7Tu/K6HHvGZiPO+qdWZ
4jl92Kqy0AlxKh5w4BN+KLmjtf9++uhOWEXUs55C+pZscVWhyxiNukimxxrqyATQ
9Rs4KnN3xaNeQiT9AjarAwq8x7yAEJme2QNBMxGvp2sIWr8SIwA4/A0Asp6bw3+/
2j0m85WTDHi8/qyc98DHDaIIKK1Trnil+3WwIxbGDTA6atuDhBBfIDIu4gZmd7By
LSREM1TSpialbcqOflXYkmUVgQD0RoYGu0lb5pJk/RBNGtVA52mBqg5z+rBC7EJv
LQPkx78ymIqkdt1ZPejkAFHnK7j3jHEn8OO69YBggR+DWUjs2qfC3EfXh+yjT6rT
uTHCXbWKiIWnG4muwh3rgRt+Odnp2FiTmXfdd6hEt3r9OJCnqRLY2Jsf7BMeCcCv
IhNZ6eviCgFn4Fl9r/WuVU6sSoND95s4TdoBmxr2BXlm5KY30sIhlwwsOujHVPva
2QF5Di58ApPr2bV4RBcuMznYMZ1U4OKczUcCfqvbu38v8IPGDyPdqNJJz2RNQUXG
R2uqJWR31SFmLYGisgHlAXn4rWnrnsQ8IGgbx9kr8X5cJkPtobk2Is5PH56ykzbE
AZnX2/reF/cOvHclTtA+FvFrdeiar9e6NK/EGLSmO3xgNV9k/MdXH5H0l/Q9n2Jn
TRKZpb6WCYgnKxmZ0wIsCy5CdrrDLYaWuf13KHUeD1/cTTGtAvUFNeGo9F8Jm2FV
iCM+tqrIa+3+y9GMnmGDGsZN7Jg9MgyOFR8hTQ32e5+EGa/rB20HWREl1g6IdKLB
x7a6H1iIMGtxlwb1jlbt/bmr8kJYZKnaMi/NGNucCowKMGY32vJGArrlQTePKCUg
BLRzXzk8dsMGf9mWolf3swE2Lva6l8b5snK7gmSlV2IHc5oEncZYY2PXOKSfkAyg
sFtt5yLKYQf0ZMbynT2q6MFO2Q7MjUyhRudgvg53jyvj+GrbiM7AzS6JJ0sL833G
xV5xDrqofBBK9e34uz44k/8psSKrX3pcD6Eb0YwYav/gFN5DVLq1j5BxQ/kCQA/3
YQRgyMvDVeJtiRn07yAVJIehWBwSmoBTQ+72UeJktFn/SQ2JjsknrlC5bUFC5ga9
dFoBDB4BoW0nkWGT5f0OSQ/CWO0M3fIrjbEtfJFEJ9K7/xj7BtRDHsXN9L7Fakvh
+2Nm6f6nZCgrL7rPwhFf3n6UMF0jESeZrYa3hFbDDUefWfmKJVQb79HH7HCzoG4e
lg+rH0cgGGUEVHi+neXjC6jDF8P9t3jcHF6d8H3EK4L7PrsKDBxSEXh0tccgzZl0
P0C7gvB49jNERBL+JoY9bLgpJhNnbeUQzG1XG4vAVjz3WKnAAroXHIxcrlmySxJ2
qv8q8JR+mg1tAWG2lN/crihD8p+CltfMelZ4rrb7HCP3LTHQ47AZ9bXi3z/4V9DB
rgpulUqUpQDsqXDH+P8bhitc61e1//NGaF3UrACDTWwVFN4omwVbHVzZGJ/5jPm8
eey9T6h4gKS+s3CKTc6A0MD7F8hTAi40DZUXkDrR3DDH/d+Lm9413S+fQGSmIXAa
`protect END_PROTECTED
