`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lc91qsNM29DxuEckkZ5MiUICE92RrGmHWnxOYEDi0tK0uSZ0Bbyj8dutdfXmdY0o
rNBBUE+AA2qFy/lkfSRj6DqBop8ULStpxz18xPtIZKRF/9DkT8Gnb6DselbxjBPg
B3AQOYaT1ki7Bfv4YRdrgDp+XT8oLCs0lgbj4UUNSD/ljEnuWheJCaZNlwrimWhR
Iy0ghuq+4uWhc/boIrOWaA704AyrD4I7vdom4s5bqPJs0UbWYoZKaHBk8absXa4l
FDe6D58Dfuq2F/ntPLwKumEHEZ7w3CDFS0Rk6U3b8eQtWE6STHoORJJ3Ty1xDfEZ
mlZISH8/kWFSPzILZb6PEdQEGShTGQZvcpzCXfmoncTqmaLYI6kc+98GEgd4JhQk
FcxSMrOe39rPCv2tIcFDdEXZdRevy+NZHInxkXS1crcFzp22Zmw6fXvMqLt7+Hfg
`protect END_PROTECTED
