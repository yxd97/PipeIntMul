`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdtMpxGytIa5ilPZE3gVEGmAHQCbiveDLiwe1M1f6MXpbJH4SZX2km58JEuHXbt6
CzBXOJ2WmuNPgttBWgw3Dn39ckL3M6YnxH/dZopNrdsn0RFjCq31PhMxk6RCJnrm
hBZLI2nyUx5WJ8WZVZq69GJIVxOhRm8deCPWTJw709tkJp9UkLOwevZxRZNti2Eg
K+EvE2nsnWSF+dKFPMDi81YvKAmwJ8tbe9ylXhNyiemszQHghfjkAYtHUBsDsisZ
0fkWP8DpRNlMwY57EVp6JNMwFvt6UmsAXI0KxrulEzgjG7fD0j+yTSpRKuI0fO0h
uPIRLa/QHcb466t/KUwPCtV0xghR/fGuL396v7uPkwXO731q7RPaF+z+Fwn1o/Ro
gboV6BK4k1hzV4jd0kKJyRXTi5US9VepubAwneto3n07AvRKWo3xNpdMdexqZdBe
CWZmPjwMouafdh0wuk8y4p8aOGgm5WxoXgLCDkLPJnkUIoEqOZ5ffRlxKmJmKs0z
HjftyhX3w9MP1KN768eWI0fePZwWLsczC66hYf/FnLcK8ZluWtWe0byGqm8QGtxt
32kiRUu82DlfWuW8P4OporbbsgRNJIaJngOgk+2fU39HtSFUKlaJHqGV/IG7HKYg
QWrAMd0dkfswRBDoJo8vydFBNpVRyPDpBiDQIsPDuSd11Sag7TVen9Va8Y9booXI
py/Hn22+jpBaqzGdHRx2FqYDqu9b2T3jk4RoNXdRtok=
`protect END_PROTECTED
