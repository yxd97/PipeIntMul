`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dMREweglVLTH+kappVakDhYdku+GukFP3F7p0BFeCxzF6a1pZezrZrgY9sxsqrcg
Cj8uHuwhrHJDqclNpmWX8dOz9fl9DhcabBkh89Ybd9WTYRGQKH5ZRveKQKvGH27e
sD9NQB0Ym6zpkzNOxqsLkD9WFYydznedQRMkn99K25/xbqt13dvf19Ndjqi+eVsj
es+i1YaeLN+DXAsrbYATQmJQEoxNB+tmFhZlKZB5uuBeo0sQ4XQoq5VAa/ZDFU5b
ks2tupYV6iz44VwsARhJk+WytBp/kTOxpPNHg4ZZoUEiFXntv4GmnXo8ezUiXE+F
+aQXRVpbaz3n5vtQpx/cz/rjv1/ighWx1mPjKfqGpWRpx0n4/nauFB/4CFBoOY3t
AFQLRMdQ/vkEoBY1082dLEvREroTbgfEb17nWOO+7J75HmvSHk/dlhVDYKVqQmOz
YYoKJW3MR/qMHvAtR2swUMHNUg8Yb7KctE997oNOwG0dw5XKCkJRKXOQfCDXRXt4
`protect END_PROTECTED
