`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rPKhOPJwuKZxwXls6vv1qkoEZ3mJP/+oad6uf3qEgp4opUG0jmzJoz4gr2yelhzO
4FR/tYuk25+tKLCWvcFQeGfUdv2lsGMkotnojSFpBW16NcnX10MK3wZdMKNjXvl5
iOSHTsFRWeHQSie07Jmy+/6e/zAn8gfGkYdpszp45H4bDa6RzSa0opAPYlgrxH3t
PCRKZPxWFIwSa4fh8MmV0yA1uJ3f+qbDUZ0XCFT3/X/V3E+s57Kqw0+1LGUSaR4Z
ONb/L0WcpDiCFvtO1+q7uWJXsgETVN5HXXn52kdtrqAjcBjK2+p0fuG1lrTqSxQH
YlA07xiWZv4BtRnYznd0I4FPs0YyBRbQTTKU6elD1axRpFBp+ZpN61bZU6K1u/1t
/3wWuW6Jm1Fou3Amg4Y12g==
`protect END_PROTECTED
