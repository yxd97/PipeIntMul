library verilog;
use verilog.vl_types.all;
entity X_PHASER_OUT is
    generic(
        LOC             : string  := "UNPLACED";
        CLKOUT_DIV      : integer := 4;
        COARSE_BYPASS   : string  := "FALSE";
        COARSE_DELAY    : integer := 0;
        EN_OSERDES_RST  : string  := "FALSE";
        FINE_DELAY      : integer := 0;
        MEMREFCLK_PERIOD: real    := 0.000000e+000;
        OCLKDELAY_INV   : string  := "FALSE";
        OCLK_DELAY      : integer := 0;
        OUTPUT_CLK_SRC  : string  := "PHASE_REF";
        PHASEREFCLK_PERIOD: real    := 0.000000e+000;
        PO              : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        REFCLK_PERIOD   : real    := 0.000000e+000;
        SYNC_IN_DIV_RST : string  := "FALSE"
    );
    port(
        COARSEOVERFLOW  : out    vl_logic;
        COUNTERREADVAL  : out    vl_logic_vector(8 downto 0);
        FINEOVERFLOW    : out    vl_logic;
        OCLK            : out    vl_logic;
        OCLKDELAYED     : out    vl_logic;
        OCLKDIV         : out    vl_logic;
        OSERDESRST      : out    vl_logic;
        COARSEENABLE    : in     vl_logic;
        COARSEINC       : in     vl_logic;
        COUNTERLOADEN   : in     vl_logic;
        COUNTERLOADVAL  : in     vl_logic_vector(8 downto 0);
        COUNTERREADEN   : in     vl_logic;
        DIVIDERST       : in     vl_logic;
        EDGEADV         : in     vl_logic;
        FINEENABLE      : in     vl_logic;
        FINEINC         : in     vl_logic;
        FREQREFCLK      : in     vl_logic;
        MEMREFCLK       : in     vl_logic;
        PHASEREFCLK     : in     vl_logic;
        RST             : in     vl_logic;
        SELFINEOCLKDELAY: in     vl_logic;
        SYNCIN          : in     vl_logic;
        SYSCLK          : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of CLKOUT_DIV : constant is 2;
    attribute mti_svvh_generic_type of COARSE_BYPASS : constant is 1;
    attribute mti_svvh_generic_type of COARSE_DELAY : constant is 2;
    attribute mti_svvh_generic_type of EN_OSERDES_RST : constant is 1;
    attribute mti_svvh_generic_type of FINE_DELAY : constant is 2;
    attribute mti_svvh_generic_type of MEMREFCLK_PERIOD : constant is 2;
    attribute mti_svvh_generic_type of OCLKDELAY_INV : constant is 1;
    attribute mti_svvh_generic_type of OCLK_DELAY : constant is 2;
    attribute mti_svvh_generic_type of OUTPUT_CLK_SRC : constant is 1;
    attribute mti_svvh_generic_type of PHASEREFCLK_PERIOD : constant is 2;
    attribute mti_svvh_generic_type of PO : constant is 2;
    attribute mti_svvh_generic_type of REFCLK_PERIOD : constant is 2;
    attribute mti_svvh_generic_type of SYNC_IN_DIV_RST : constant is 1;
end X_PHASER_OUT;
