`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UOWFUB+tCtIrpFpUeDTpsGmAGswDQtSd5CfugxpkSVrMsMp4OcTP61uyAQZrfRr+
E2gJhX8PeYWCwyyoGwrjhNiggr+hGx0nwFW4aEqmA/UCLzyuWEJq7leCqlu5uf1y
/1OQqm9FXJO8sXy4cSJl7mXyKrf9QpX/5mQcFxQxLkIx/OKbVbrkNBwtkOFWi1IW
igKfTKFuSRK3gAiInMbD2zCa0CcyR60LIPw3stOBVehwkWaR1dlmbaMeLOESrkto
3mmxd5eAUFVJIXuGy5b+tIdLEaKjtTtKFI0nBk0AoiAcT00NRXJas0++/BDYW93S
H37lmCCp4RhuzM7SZdr6Vsnj12ZsHNOE96RLTAQYGmZKgfbq92CMbgIC/GjpPQZD
fHQ9va6/jhy6ui0NAelNkg==
`protect END_PROTECTED
