`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IFQvbim69TxSAZ9kqZEviWCpYb1iUcp2KRtCWd+Fr8EMIGxfnER4N8uYfCU0MDsc
3ZQWaGFMPJ5YA4kp1DfPt2gXjHIWuIM2D7JQOofM/KvOduPfE8N7LmNy5GVpKq0X
HyhaGhw0LsrNdtSSAFJvLsdNLRWGhQBtnMOWCEWZbxoS84eqCpXIXO3xo6bZr6Pi
DeSczVOqqUBOBzYTlJoVlAbVNRNQSJ0/2ZtEs6Z2ugpXcHGbJfFlMD05qMNAViFz
lpQiyNZxBOjEJ3HlOaOzRNnl3Ek6x5lp+TBE+y1cohaI72cH0YfIT/qbq9+plfq6
8SANKj3+BEdtqGnB5pjZ2CJQoymbWwoMuXBk/tjiQ3GmhtkVUJghhrx64QV5Wuqw
zoc9yliffUeobUlB3EoSpW400mxI2EEXYKGmI9RRePYs/2Rga9It438UH2iT8tU5
iF8gUe7MqrKnMNVREuUGdHUq36HUJVR4FCTPqI4gp2K8FufonGIkWPOFWWaU3NGc
D8vATnt52FZj1NKP7VrQbqhcBUJ+CGn6LWBzzcESCY0HpWUvuVZO1yk20GgGtrMB
PZVKKM/lb5kFCQjEFmoyrK2GW19NLsqE3XFkdryn/0nB2LF/zUSa5EnVacCu0N3e
hf1bdGsQhGt7PjCtzY9MiE73Aq6DlV34EJqmFck4ZQ+rHDfRBsLwfmfxdDyTM2je
4F6H2B50vN5XcfjrtR53ZHegTPH/p8z1ZnaNW+DivMPuarzE93kPV9plVJP9HPLQ
4my9cRrls5EBqZpirMieCduQ95uT9gWFywSnu/fzYNaD/+tLLAEi2ZUjVzqac392
VI3QtulPjHHZBwdOFl/1fdIy1ZF+pjplVrsuHOabItOWnBQdUnzB1NChI0i5Dr5W
S4sUs5voeHOLSJF/QjHambFEByEoa4RqDp+2LQBVNP/UHhk4uWo0mAS3NiO3+dSw
mP3M2IWkiub+LAkSzKJmCrC6v8AGqih7z2YI0rGIwyeyO7ZyM4/AuYrNrSRUZJAO
bQ4Uz0dStwohmhud9mjCMVnNPoGHrWnwK47+PqJUK49Shd9BChzWvyGsHOMcsuFP
U4bWaP9KFU5VinRmliE7wz2DS9+DdncYbDe97x7zhuGdpns6grM5EXN5xcDJh9vV
/ryBoBGznj682IGReIPJYQz55E6uz4XWmCP6JxjmHrH2tmtQj8iTvR9aJmT7DryH
6IvzTfyGXU2ZaV5Tq55HV1+QfNN9AFfjdhioT+E4r67HB605LCsTepHiUosf2Er8
LKe0u1wHYzgwome/8UQ144hDws9C/Nl3fwTX1PTazGWCAJYJYLTXlFSC3+lZ5SGP
vo0Q80cdxmydxFDKB49X7LBMxOOM0BU/KO8AYYS+SjZVUpn7brD5DRl51m2BRBdF
qZsEF0S5KNo5f6c3xMe5CdN4B0ztl51cWfNJ7Yp1hlD0b8+Lejolq+sLQ4mA7J49
TgjUjPB54uHPXErpz+RLHOpNDhlyjxvOS2e+pmYfA+IJVMga8Nz2SF3jYZKb0nLU
fEtgD8n9xiCaY2TBwmYQ9ruJFNQ359e5nRQj91PV9HdGy9NScDYNmYPlvPiY0ZuE
/3N913mTur8Qi52/uk5n5vpV80E6JWRw2CHmf/IHea9cvGguvjJez6Ujej6d2vM+
hwPTCZqxmTuIa77egL9pwfBee1VTIYEBDf36AngKzXx9LzCOEMUdVr/eNUhhgvwG
q9SDqWLAHTYZzI6QqpNvcCrqciaI1um7K+dOhz91J2X3bRiDyf/NBJZKHp4p/Zao
EAAnnqZaCVwuzyt1vFaCRoAHXKBtKBx0UIRDSh+d0frEI4nuuRkSQ30Ktte0xrdu
9WPQiqBJGbDiVAdYHwQVZZ12TH+v1YU79eUbgS0COFasvMBCOZ20cW34gXJn3okK
QMfrB1voiZSfqIM8rd6aD5Qm9Vk76LQ31HQueAvQb1CcD9Ru6aPx0Zkwy2J7/Bi8
xnxQkeiDB1g6NIpnaEDDS0GckEM0Tz2IV1GwFbekYMtoEQKwR+05o+24eVBrtxZa
u6S0CQ6rBxl4fO7IV/mQGRsrmrbUI6Zm5sLVNVyfKIZsG8bnzhcjcueykPWZh/fc
9SWr3XQEF+cm09fTQ7H7PmZcUVUKnlr6Tn4Twot8klY5GsbxVQIdZXbMXyRzulil
Dtah9q0W48iZ7XtDj5mgqAi/875GOZibFqWg4IZXIGZ/UJUMkLkWVk2lVVjFLfo3
I3sOdx/aHIq8lBCn7GhN3b6kPdd43kK9+P2/e+rOf2vO/6w7ZEtGKoi8EUfn9Nfz
HTZFQSmEYNzKOnGaqqRBm3NgM0w9qJX6EnzcXkgalkSM6D7EBIFWDOvaACdvlJ+D
w9q/j37JGqJ6yMjnxgv1sgzn6+VaNYApUXfwSzetH9hLrzaOjBaISJXTMd/4/uN6
AweGj0CLXqY29RqWIU3fq74szB9H10Cgo4zwiFgJA+U89IcXKtXoBDHFO7TNXpYF
oBdxZur/6bB0EEjBGUx/1Bcc369Shb4HCyLJdM+Qjk/KVlRpGnnLrB1DE+0K2Fv+
zQYFOXm8Au+WdoosfbWNve7Vj2IafAOGVJx+aAjd3/46IY0zGMqzSnZYaCVqfYBF
EgkU7P2Fo3Rg7Kxe8Qj31ViuCr+ZFG7Ze8pEtnu3kNUNcwcI+3Vx4ZeNguBJ1IZ3
GQ2trOSK4MYdjl6QSrgJeMyXxMXtmt+O6QmtV4ZZ+pZa5FpCfG7pIpo3ylpjmll3
QA8W9Y8mOx14B0G7ovFmooLDSNGKYD10Jb0QM0TPbXpLkuM4Mw39hFla6d7Cg36w
3Ge8SzueFGWjH//Vz419ADc+N3QGiBWwDTXb3iXwCopkswSWUy4AWjM2o41n9bx7
B+T1cKeB7lfQg5WZcmvMo9ybdw+61UY6KgUMUEU6kirXaomq7CpV2WsYHxEh4+fY
nUj9GT+Vn8lZgLBnVXCCiaNZIn3Qd1TtuMb2Nexn6vQ=
`protect END_PROTECTED
