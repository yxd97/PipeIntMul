`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ngoh2HTOqy2PdZdqbqKhkl5dJAghNTvcNB3IDinorHsENJC08Z/0PSO7QxvlpEd7
wkB5lMIZSjzAUy8XlKJQZH8p1qDGCI9DZBp2gxWWxueTP/V5UAfEWXAGixq8JWdk
U7ONuy1LoVZvfmrWj0Q2+JX1DJ3oMETF47yuS2XOMpa/8vdT+K++glJ3jGF0d2P8
uzPCdzx0jD/icgwENvIrGTgcP100B9NuwN6gMVTOlWlqn2bj0BXCN83UfDZpeAx7
hKVZ0hsfkV9HzjsTut76QvZZ2z/oSsGRjjdZ1aaBuFUfPIUyEzdETtbVMo3S5fyk
jbuCoAIqozMLSuFokRtReOAlnV7U1AnyyVOHelOKOzDOviJZiGrUq1SJiagG7l/n
N9CSuK1R4iGIOli/VYmr37HdAyhPqmPPqLuW5w6Exuz5bqEhxYf8KONjU3s3bef1
p6G8Pal7qOqDxYK9MfZhAD13aNBEm2cgeRijUgkTk/Cxnbz/zKFAiQ11cp+Wp0Oj
hh2ZttNLcVYonnkcB8ouPWnzdnJmy2MaQRe33DEl1Q8=
`protect END_PROTECTED
