`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pVMXglNoEHh2YnKlLMPN7OZCkOri4Pb+nzdOfoP9EfUxhQpDPceEmPl8UJoAR+TA
YBn2KXxya8iTrxElrnHgNdzf7aY5YtFt8eLBwFx4EK4Vl/p26kThZeIep2fPTCes
dNarLSZdrgjYAR/dvClTIiPkdEdu4nqHXZ6V1B7BZyZyZQ0aQaXm0Hm+vlAXG3lt
l9w6wf3hjEbys+/Vd5PJPXc73338DT80uekvjk1JQ6n53v8pVdhaNMl/z3PCPJjj
/HJX72rTa+/mp/HQuyyApZZLGSePGJEJ+afH6bH/gBT9jK4dO+VjU5VCbBK0bKko
qUoylXiD0TAXqlmVc5CjRG+myGysIp2N65o3DhwIoX5hsbSGvsuwjVsBP15U98Jc
KDMR9gn+pJ20eilQ322BmCTUalDMrqg2OPR1i/yO6egUBHywn/Fk3dyHKycc66YV
MkzkvPQh7FJM3SeiBTZYXZ21TVD/umz67/lTybOXwLJdG03gBBx2gQ3YbR3JJJpH
lVquWUQd0rclV9c7lYD2gSJcDzA2fnrTaTkIFhlX4S7H6TfEsRSYhjBi2UDzgQpr
nEysOojiPRZRgTdvO7KCnWsaYG0u5xB+IY2N9+lzZj0c0gOBNg/hywHptN0vTcN9
Xijry4h0KLFeS6mm9qHaFwjTA4mr1mwUPPRShDJ6QVBFxj3pVgLGvpNE2quBNLQI
waeaAdfRop4Q3WiqaAQjU/fKdycssBuYGRGvDIf2klibmWj5KxGvw4tMkO9iPc39
ue1KaAhDPUq4C+xL7wIl2P8bsmYfj2Nhms2G12gyKOAYV2RqJyMG/l5MJHgkI1ky
MkCz8xiZ8BBM+keOV/2y70M1Y++tZzc35XXpWfBuWYbbW00Rdqxz7gp0nObDBpuv
inmv0NgHlXllE5L38KVW0pRxorjy+8Jw7BoawkoYB9lMSooQpYeQYFTtNJtPIKsv
r5VFlesETNFVi7DIxzVKo6Ime4CSNL/44R2I3WV1M1aRfsOQRV814/a8Y1H03bGw
ixQ4VSLTAMIkWCYxuGv8nOmV3rS8zl+cx5IpN86cn6v6YtV+El905loWGV+9c6Xm
fFBQkby/Z+xQvAHXolDULXEiB4FfqiB9nBxNI0MiH+Jx4yAeIGsFJih9XSz8ghZu
4CNJ3EgAZ7luBlca4Cn8OCvT/HLm+V2DkuIzKnLUcUc=
`protect END_PROTECTED
