`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
74qmdwDW20NDcHCHD1q28arUblKHTZJiOlodbIz+r04lHQ8rQXds3vLqYNADPAsP
HvV1UFiLilKjApwuJlBBhBQw2eRICxkPmVV0+FwsRzuDsOfsvVQstUjYHADvngQC
QdiXmyIU1FSLNE+clvXKXUi+aRmRWXry81Ekdh2qkEOj6yoZf+bYVK2lTIfPHk12
X9A7XAfZTVcJbtS322P6rYlP8oOlDI0CR4Yah4VKPBvAFm5YNRI3tPNYT4+VxZut
+2uLb5ap7V7wTHYMZ3wvvrRjv6oKWiiSfTACMAkvcd23o/xB5ZrIilwJJxslTsNC
ejIhCqK2Juo+bmuchYIN5HcD+jHQ38F9/WHi+Z0h2hLLdUrWBFKHuSJvV7oZBRH5
vvo26H4lcTpC4xxOIwJEpnlCgVMUBme0z0oJJcby1YqGjXdHXfaFQS8W70kKOkef
uJu34xbg592mJQdTwXqoTcad0Eikk5doorMLQ0+ueWvNC2Ny432sO3T5KPhpFjuR
m7T2Melcxjo36VFugUlq8cBd8nF+Ro8sT5mq6GFqDybh8g1rx27VSBbZDWWblx4t
cAOAFksP0PyZ6M6TiJClty4yGNUKtkm9KqDcESIPW1Y8TICfEKYDCD0sV4q2DCsR
m02iEQhdYQKIt9LQwpPY2saKbDaeMu/LmQ7w5McRcoSx8uEIOlzGv6lszGpAGHlN
1VDxGPXmKr2qoln5XoFZkfn+o1O9TyIne82Xdtq3icxkW6vYBZi8uFABliRvtVXX
DWCKRB9axM1kRiT7h5a0Qyxv0O8f0JW0zlSQLhpKFgqKmUpUflq/qL66+zEl8ucn
jPI6XvAdtq1+a7j2haM62W96GTZb7cIS8TB5OmfX/xQgflSaEEhw++dEPXP0Egqz
XDOKo+RZyoNzZnu0d+FClLdDarH7Da718gFT7mq7Kv9m7GkUglRVg/FmoIq3TlCC
ZpG57cRQNQP5cV2CcZ+qcK7xYWLvSACvZec6Kx01+E7b8DP1TwVlVCwL08ZQ5B6w
hpPO0+kPff7xsn4CT1lHHkacBsai1HFYSoqwzenoTXyuLW7hzLhuS4WXK/udsvdM
tRZco3Dbv02cyK1nmakyEZN+IPJqVSOcLDzFd4Py2gOz76iMiqNUI/KN969EPbEh
dVFaMVI+qKm6xghXf621IZqredQPWI9p8LMA1lLbdrU5fjgUW1njbLizemquRA+D
ToYeg5RoV/sUY54FlI/KIiUUYVwB23OjdAIZctbvuD4xIpHwhsh0sEmJTiPwAVuf
7rLSaYRcvBG9pETRReD1jOSOLxaG+leUHbYYmUWEJfnShk36cR2vLM4PFWrkTGz2
zbX79EUBjX6qVqO637R6ANZwIO9SkCUrVRb5AmoiEeRQQUIvCFRrL5p+H02QgFgD
+4vIQ1qRB68fwDPbThoU8JeMY9vmHpVt58TB2lAUlzmiX8zhOy5dClkMyXdZrySc
qldNScRXIxvgbXjMJ2zJX7pNjn2oK5tJ4D+GudM2htLzBS4RTAUlAIQY7IQ/6v2L
AuTSHckiTy9Qz4T9kTwGTWTwklA+9U1rTCQoBd4bdvwJ5H4y9M6WF7cqKoZXtEy6
A89fQSIuHieVb0bfFe6g3/lwzsRd6YHhxVpYfv9bNn8x7AUg17CAzPID8/B+Qlte
w8WFJm/cqh60aDMsUDgyNF/IHv5IjPT5eoOHBsKiCGvVZoOKVM9WIak2+eNXwPrE
6hPBK5AofCQe0NfKsAuUWiMMro6afpTsD/zvRnkYDAYHfcmWHpA0bUXZnmslWfT7
BVegUIyYNPaIivh5us4jv2a1XcqZsP219QtYSHvRxSnanWerN0CNZ5yPN93XPfa8
xJghANmeOdBWvYj0P/TdqLgGCgUGDoUqXkcOTFtDww3A856eI5tjvTj4ua26qFz8
ARCGymYoQDApfu4POVmmF+zpWjPeVYgg3jLxgRlHNomLWsJhw0grGv8U+39miBDP
WSOECdO79jlgl3Xo6wMJrFwj9oXpaNVmzXtebtG0ZfBoqam4kngHTiIIZuRv4OFi
2f5Qf1/GsdpbFMP35VPnOHJvgLTPTLjj0aStTsZgBXzOxVI8jonx8ySQHSz2dWIf
6iL5wNVxUNiQCq10/StXIktqodhi6rSi4+0Z11gr+SIVOVUy1BbTU4XbOrHFqoZ2
Ws/OYE4+WxdeSbuI40XjoYBGy/85C4+2fl+Sdh5fa/Ap/9Ao7w3Xz8nlf3Ie0sRH
OZ2e3XnZ+/XLNEY+ZXUjo1mfr6/0mI0uGdLhaOp02JaxAD5zGbE0MBfZsejTK4YX
`protect END_PROTECTED
