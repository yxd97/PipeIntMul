`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xqUXRJFQ5+40IPVYf5juKV81QtimYIk+mmw5L26QNaPyR6Hhfqm8q83xx/JxYBdG
q7xPgiHhTNtY8bddlmeHmdhVF5LQ5jbAV+ACtlKF2FBkjq8S0a3byVPGorWjkwga
m+gdhKhD9GwuMmZfYbLnmtV/jvgbPF1t1F02ayPaxKQazTB5uOxMuJQNkj091Knb
AlqEtIH+gZfaE1hdGz+q9tGqzJDQwUpFy424LrPp2c3d/PIDQt/gHOC3Q2uvEVDC
5K6ArNKEdKTY1dCQtVGzoP9grzC5FjVd5svFNZ5OWu9ZRVmDBg1DWG6mz0cqGP6Q
EcC+fpFbdwT4mOCH0hen18Qy3zV3uI9yG6YZSJbVYFvUPltppsgaCBYJ/iDzCpmr
wkxaanpaQlGrnqz+Iz3ZfMBRygtZ7XLCz2AqI/CyZAhDWYDRZz71FLX4OYipmUZT
/mQZBgMdsiycRYbjqlRVXfHKt5z2PUQU6Xn4eYX36BL78Hdafh8lPyTq+EgakeWL
UTdJnYsDnCofCl4N9+tvCsVSt4y5aoDqqXfDvFHcfgt8RhSGUlJ+2hV1dOh3qcVT
vRsSUbxTp+djZJ6wPlGX5ZkmqDWQ6gD4m0EzYx7kVag=
`protect END_PROTECTED
