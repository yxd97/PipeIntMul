`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HbB2grFGkbdiUAeH9i9+jaD79kbXtUQYHJICtwVTm365JatdjQqybglLg3N6F3pZ
F/iUarMkQUApT1nLwIiCNHsxk/pNHrempHiMh5z5BtFj8AssIIyU08I2gUmFjeoA
7HZsdVoB/cjcf+XOrItzSwOGVBK6G6zf3q/GGSItmvRczga6sPH5XmPcyYIdO8nj
kqF9IFdcxDS/cEv/xMy0ie0Q4N6Hzo/DlDls8c3R7W/QyF8Do0mLVzW7v+DFa748
s8kB1gURba8AbC2kpB9MKzhgkCS+pyMFae9/egJdAwLPHZhGkPwBxKbr8pMLidRY
qSB1lN6GpSRFXg+b1EaYSOSwJ7jjkxF0mqYAKnLh4oqQ0v7isFSxlXgpoUcqJsDM
otBgdctoaM+5bmARuogUyw+3ieJYlXRrASlnk34+G3wGBXfRj3s5VedaHyMlAKro
3sQsJXCAS0UklVMdvcPaNvML6kfiB4ekhz2/ym0/mpw9pZXujRn8nDFsIaytmLvs
qMmANNMazTjEGbRhamGVkUSl0Wqv9p3EdCqbkkzts+PIOFLXylMihS84ltApppmQ
igDc3JQvl2D7+v9YgtPoAAQ40VC0qvYywXv0PlIREds7/Zce4MZf7PTuvz+itBJc
MY6pb9ARSf+mJZSZ8irl0ekvZv6XBu/h2XVLnYAV1ebi5/PoMyqMrtS7Sd7Dx0SJ
CZLFMgU7IQROacxLUXwvHqONxkX1AO6DbkDBUYPGJpSCheeB/iZfsbZKyI54VoG1
8SJYd3di4Cx8YaMoPdVX4rln2+JmwTHWSVoquxT18okxZrcctWtT4EqpU7yBeORW
gCo0zXONGjkOokwi5yHF89yt/Jal9kKjcmRh6x9UH/fmuIPTnJLxjo02SD0GPAEF
rgM8CktlrZXblooLEsS6R0QSLsCCeDsPevlsYm3SGvjgcvEXNatLij1t4Bt9bRT3
onhuhy2i3EgPFn6DcRy0sM9g4nieS2PC/fFT+ebGZ8dhzLVyswPrurHVdG8xuQ2Q
AVg/nazqO6b1BLiz2R4Un15/0WCfJrPfhbNHRKTz8R5QOoNdsNP1U6Wj9Ws3gbeK
O8JhM71Wpd34cxM4pEUH8SetHe/jOxbRTplyH+hRHkENfi8O3klcCUdGobUDkbRA
re3n7fHdQR2/78akr0/pILZxywq5XZMyOBYChMgi8luhEB9ExXAWGeh8shV7fDnX
V+uj2gPd0cR+7UICq4s+z1nWxUPdPm53OLR0RuCUsfEJuYYSi5EvoNRoVyNS1a0o
AOBZfo4D/SpJHlxNLuZ7o1Vt5O13RU7xDwYyvEOeEepE9+Y76ncx/pB+X9nHrhKX
XBL0LV+Gxu0Wz/0jH8brehZg/j3JZSmIyOnp/9sQ2yy88ky+gTVrbjpKv5J5k5MJ
INwLqejhLkmFCb4thH/caS5geAXvp52KOd1szdwa3jo4GZwzapEJM+zcfkEnUO4R
JxBtK2/XBwFn+CJ0cQnylUA5h2L6M5ZcXkWfRlHjFZxEel1jpemF7mI1Ol2+1W60
9Ivt60tRaprxn1/k42/uBxdtRjmRMJs5pf8YPhVOb5GGJqeHBPn/jAtgkRcLA2tv
aoE7aE2u7RdE0fjXKew3jUGC1tGF/JPvtsqa8boPFo+4y2HyFBqbKuUOuFPfWvJP
4RcKvz1l8atG1SvRdnawquFBdyAB+VDt5oI13O3KDYm+9DVwP6t7dn0ti9Dyhr2L
YIk0vnpbsJUr5iXRWgFeT0i2bTrIYednmJYCPNhXOqkHzKJFK4/hTr6X21b4jCl0
r0qva9BNIu+WMvN+Gz5DF6AfdXyv1f+BQwtyZzmlPN5IAbQpgcElkbVdstXCLIie
4bUawz5rDUobuzrbfOtrHsCkTDk79FlAkrgZxEr3s3C/Vd/vUNZFNAX7CWkxPl0U
H49PG2Vvuqfa/PwfAU2J6wwhMguMdtsnqlbtFB+aTBo26ykC3iDjjv4BbGHm4jXx
LqkegJ9KkFl+DaS7Xi6+rU0CoO8DnbB/erfGvFyiS9/Gu+m8gykgWpwG7ptqB8xj
0N2dRwzfunVAsUKDdQoUwM63YgJJ61Ql/T2S2mnzquhuNC8yCoWyRBfuobl/hOAu
8goUxz9/8yg6ektKDQDU2xp5urdQnz9joBPKqx/nFtIpX5EMCMV+G3Flb4T2Egc1
RxnqvrqLAQqZDwpKtla18xw6eNtsCZD+ckLE5s+bPRvO06Mic4cQqDGjeJI4frAO
BuO/gF1rSgPKRewFpi6xLYvdiT57nEmzZB7py3GBo0ohdzP7TWroAU76umB63ULf
daLOcLeD4B9o8f2tfVZ/jAmehpl++4wQP07aQz+aMU25CCXpiLCUfJxl0HbSSe7Z
MqTGNe1q+FYwde5mD1wFjcCutwXqUx8vcz8ntD8ao+xiKs853bByLFbKh9PgvIeg
lRCv4voQY3qf1G3jQAgeEl4ZdNE31i8XWEDYGvMQMcqkqU2JejydlKTFQ9GgC2Mj
LiKtQzOI1Ce19fwhyCc/laXkR0fnzXIds1H8e0HEeWSL6biDOjhGJYjdrD7L+qsz
XSgpimxTscs0HZeHbTxfJgx5a/8vZ9G+CASr1BTJEAQAczfLz/hpwM435f74ZmFX
Z3cnQMl4NtQLNt1QTIVR2A7q9rmJIoiQJlWKTHO2IgBWLvz2FfU4oixpGKI9o6pF
6IClqLm8cweDgwyhPyqhAo3EOw9Z2hvMQxMNxPYP0H2dpN8UkKHTWa1JTYTeNS9Z
XSj8/1LVZP6UiXruI6WFJZZBYAwj1ZJ1X+gpv77JZqinUpwQPxx/eSTBS57Yppmo
vS/4Si2yRMbE8r/V2uxrrsuVcRO0L+e5uac+HAyYq4XNVGoFKfFNhr5/utk2DCaH
WaOy2Za08KE39tm+HtIlWUVbkutr+1Rliy4yzZiM7LjCQNON8E7hdZ86RFbcht71
xC2VjuMMSJ1rwaOPbV7CpuGCO3ONB1gxl2pCfn+VG8otEk9OpLdCMayNAISBX9p9
bNROm6a8bFuJb+J/+mceRnxODOa7lf9lAZuGK0kmOWLjSXrCbHsqBT48t9Zs0pWb
G4sf1vs+XmlwRtq9w2NN94gPmCDFvbL8m17EdUonjbr8Gj+z2TkYa8hJeSlt4pGZ
g1H8AjPqUQ2AKLT0EAC0IEaNqToDCnb5sRS1oQ2mHchwdONEteA/SUys2l26ZyKV
qorMX9F6FoCEO4OsIfx7F8hKiPiQYokThH2eefjN4n1QvoCUoQa6RVonXMBfCycP
HV1We7trYv8ORGjC/JxYEiW7mYjxe+QUAJfmqHJsdn05q7qfNwrYe5EduTyXVyQI
9/5j2/oGmvxxw4Ddtan0cCyDwPMMrii70MtUriaVOOqKYsWZHZ3wyPZsDazPKeFl
HNw1Il7ArDZtoP/ExEh7osRnnpFbI71wMN+Hro3eUmSe2SGv8sSX9VTqtkKWzZ8O
wttY+NYv0FrMbjnqXESg0y0jDv5u/P7hZc7KaaUkpJf1o2PZOn9rZ1AV7NciFaMT
6tbDgPgd1N09CqqyezAnppfST0gkpanBnLxmvNvwAkGSk1pmslR918v4G1gRfrFQ
ZtBj8T2nGORa6IT0Tf6h/QH1/cOFGkh0DiDmS4fakYT/iUNwPmH1m7FE7G8nu4OZ
M13pgpEIJ2RDLixi/J+cSjGCM38P2830CtMOpYYxaX6G4LSFsr7dCdQHAkwxH5A0
2hxw0omdWhkRZou8d/RQfTwxy9LRhhVFCZKnXLFv2hY0SGMK6Pf9FMz5pfuXVvgk
Brnh7zCVRMVhCov7EU5RHxOIIWNnuczAOwBj2Uy4ZJsLEBh/JLhYV62DlSlCtEpS
JcvfXd/c0dWb4WrmfnjrhTOuIb8fUu6VLoG/buEh0iltr3DCSAVopPEkTwGNQE2A
nDMbu3K8Kd9MbI8cg84xxQTOfDR843oO83sVhgB0APoyOXQEzm8H12Zyx2H0R5xR
McOLTVcPYVo8YWm6fpFDs78fN6YmD7+1fpgAbhiizQjI+F4NShTV597hhRN+4Le7
yDH2E6O7w0221paoZ8yI7AEKypvJg10KEdIOBYRoo/0reH4QRreKD4POrasDCh+o
5ITwIO1NPKR95gSwtBKvQKidOmIm7P+2tCUsjlDPg62TCWBNQGpm1hmgOjQuANVA
nv3TdkBqLcXnZmsy1ktPxtWyUcmHPct88sl453yNMSz7oEc5uR1ohYG+1cJdWZUY
vAE/1y4SAznNRzKDaD6UQTPlIKNoQqxHx08BMG9LXWIbWtyBRBTOZXqEAk0DGCKi
oZ9BMyGY+6VNNFRpzoteqHFWor7DtKs0KnfXnruUFAczw7pS/CY5jfdlf2Tu3Ayx
IHVDAIhK0O0YQ9F09ZAsshapD3OXb5FF5LMi2+WJLuTKjb+0QsL6PBvQMYdCi98k
CzKsT2u4e3vDa4IB3BCwHDE6xhBFUxNC9VD1UVz1MIlf7E1SAi0tV9iw+m4Mh3Rg
bpxQIgG9eywYtv+1ag8qaNYGYbxwcGaWEfbC3ahvYPJX4RjmS3tCw4+fyPn1bdEf
PDDnuIrhsrSZ77hhkkbmYQ==
`protect END_PROTECTED
