`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAWsR/fTVjAfOHhL3Fbr+WuCkm5SLQP8eLnjtuEBvmE/w3F9uOxIV6T/SlPNKTwe
ahXE/x+lTUw+gsZJg47Mem19X0NGofSjlcJfJnXw0MGAgjdnCkfiC/vVdJHzJE1r
9l5Ux1XHiPmb7PKa0k0yszUE2ojAgpyZ4acRbQS+0RJbelz5x2UTpQqiHtuf2avg
J12MLHWpYLcLTfb8ykRHu8HKotYX7YOTQg80Y0bBNKiDk01EQETILvmaDDdZJcNH
zZhraGIz7MHDpw/bNrCxOlMiokm/N6NSPSz3kb3UMDOtdDQ8J8yxgsFMSqq93y0C
LxwyYCCo7rhyrAQkI/D5SwA7YpsInXZROrcVEjVYumBs7nQrrRSPKhcBE/D22kMS
t1+XRTXq4FVNVEVweZLoS5aaKt21zBnPEalBSH/8cgyV48eyxc3fZTM2O/x+ul8G
4Mcr7cQTlmfDGqrNVEk+el5uLUw9TOATdQC1z8UoJMxVM7MZNwUI6U1jpxiN1gxu
OCPr2KjwdiOuS36AsL/orbsNWBACTCxcnMWzQX2rzuk1tJPaC3IyvmvisJRuGm6+
EWQlyC4O8VOAIut+lpiu0N54z9L+mToh4JmC6VbN/TzGyZ83eoEPMJBIpb+bEwhD
IkOhqrv1bM0fvpGfJlVYsFtyT0Y5SCBp+KsUl5KHLC2bVxiIFQs6UvLG3IKsKqG1
UTx270S7TxJ3hAdhU9dEhRmup4cuzZPiR5LiTXW2g9cDQ43Qk+dNHIhFKAyy+71x
hZlaZU3Wnk+KobqkQZf2CFIyqh9gYaOwBRZDM0aSjDSGvWpOd/1lNSA/fejn3Ny2
uRYk0DJ21njBi4ozvBUbKSXIQKdhM49vmi5jLmwOD0mnKdd/iDGd0wjkUM2UyDXX
JzmtCvkg1SSInb3qbpOvUZxoykybtBWWxMmcc1DvOAPK+3AmuIh8HqCZWWIkZcdU
UfTtRLIg5is8h7FEqp8BHR/IZb+nRla5c11K+aFM+69RU9kw2/lRjGk+67sLFNpj
F0YdYSj6QmNngbLq/0uTsALzDbk+wgmH/scjVNDiG4G8cmUjowc3cWlkTjXTpo5u
caBHJCxeqQoY46ZzDxWLpwDtgBXXZ1N/P0EYnkrg2ENVUGAv80f56O3FaFkekAK/
mv6/GR3QM6vKGa9ksgBAssyo7mlmTf74ZQjVvoYJCsWKaewFpysSv9J5AO6eGCc7
08YHAyaGZIgUQ/xEu6zS1o3rwsmlkWVDy9+1Fj7upPSODj4flwqM/EMDDETzo31R
MpueGh6o8WCa9h+qqPPi0tu8asF+gSQP7jTyklnwZ1YfvJ2JTTiCLSqx8RWibciq
qNWMeAlxeMlhvHtgcBwblA526LxE6KL6b9EW7auS+4K6kDwp+O3nNZmRwG42wtUB
GXqxdRowm3LxGIyFYcM9rUjEl9DxiIhvPtj/8MYD2TFHhqXbKy5sIxHpFGOZUJvJ
LQyzjRUDn2dTymyqQe8e4SsCnlHG83pduF+IVjyCxvjCkllmQ0g6I3s8AZHP7rok
zqX3kKfAWvFgo+c4VXK7Gx+pu9U6PYoHcmTrU6oaCtdOwr6Ymu22wE/jDfLNX3Ms
UUi4rbdrLxvkueguShZL6CNeHkbh+1wC/SxIkPjtYvBl2kn7eXTAI2V8biPhzSqG
Ps74jbueFTHITwEODTApvxC0ODR0BmLxrZJEKrox9hLpYrHGMwCUgB4hUt7X5jAB
lfXaPrmDoPLDKSemIYedvYD0kwd8dic8sZAvNqbmzFhD2QzUiqLvn1LEhagU2XU4
T6zwS1QYbvvk/arPuDXy0mtGdFgXExwdk/vSy16UGgih5B7oo4PPdErv6rsuKQCQ
RMKIG0CRxZg/OXll1Xp2PNx2YqsxnYc6rHYDmVLBmsiiZZZMTtx5hfk4fWzRo+tA
dsqxW8tB8waz16pwDyNLKZfIMF6jBSsWECGfByuIcsmYzzn7v/6FGCZapxdHPsZS
KMNbtX2/GNEiciPUAGnZJQHS9AUZZXWO0uctMLZNl0WHl1nKCaCw381PInyHZe9m
9QyW26DE2SoUUiOts36U4hmIEAdHRkI9Lk/4emOG40opcSpCHl9ADWqQbu49op0L
22D2D8tYPyCyQCY2TmbwpQncrmrxfdnDMnrFeQdI/cCBDCJxSxzTPPQ5jZgeuVKy
pjYQj7qGxZeA7Mnyvu8NhLFH8zrPakqyJ/vTR9pg9zq4tFDzNqu1jhxCevJ05a78
eeIa1ykzKLtjA9HUhR+GtjmUNywPJZ1yGamRseFtr8O5VbDDhThz+ZW1LyD6JHIH
3pzS4LjRGdRo52ITTJ/SlIsMJnc+LwHfatLeMQXsHF1h9KblDdIlL+nqTHRjzMdx
wWRw8pU112XwsR8OAS6zjiUoOwHVoidBghrna0JctEXxOBGuHhxTttddV8oijHIP
DuygegYeGsl4flEcAaVrGZX2nr4JXDab3zPSaJayLeXNKYVkjGWhDCF5UIP5qE8X
FiAeCg+WM9y9XSxorINiYNTpHGwN53NTXYPZM1JsNODWSE2EcRAPWc0SfOlBD2SQ
B4Y6Ei9l8ZnC8/EbrBgfS5Tv1lBBTfIpwzTRP+rDXQCDzv/uuWYputhsnnrcd6FT
iEhrmsgbzgVXScc3C7BwhRSQJ5E1g6B/ifYymCP6n8jRKAuQReUavaHsvgX7hLmI
wcy0AeVQfKSsnpgdjQJKei3zRlNgGXTSlJrwKCE/ys45xrL22wfB9wR9vVb3bNnv
c2ay8EiB7xAqRHYUYnth7K5q7HlstqHItMPyGQCoNPvdiQfOLoTgFgNhkdbpFwnj
DUICbBV3pQVh4ev40w2kp9J4QAqfp5yIaYefWc7erL7opfUCkfkQ2TdKQqRG6RRQ
50b17pPQkD7gD1if0R4ORm37WJdF/8r8xzaBun5rMh+SzfEdxfvNEHoFCNK4BZAt
AOsjiWLA1tguXvGZyCPpiLJws/iw4S8OG+PW1a2aC2OlnblsSicoBZy3kUcuKxPt
arfmTkf2ZqAcSjhQwF9qg7117yKLRhNG2K8BlPpyIJ9tEfclMITTEO/fa739a1+/
CYDhuHfNs2VzubFSzyIfG/hrpd5chwjJEfFldmGCMFrWuLOQzvHXmyWzP0gBGQuE
CmHjDDv8IMVcmexBTruNmSb/qzrq2euAI1y00yDESnP9t7XmNNtjqzr+fPPISu7O
Qh1PmzhDqCqMM5lCMlavcDNyf68ekkACMqSNmM4oPcwnUz6OAN2B7t/kpbLl8N5b
ipfTjRpZR0/hhuirEa26lcwMqJi+9hWTnMhsI5nY5LUtCx11MDGm+xs85ivSaZZ9
PatsVTX8x8ZA1y1zDY4gtnt0O7Okt+cvN5oxc4Xzv+7J9dkshZwqyhyvAELTC3Rs
blXT1eOCHmlQadUuDejR/jFo0esiLjXlXli7BqP2aI7IY2kXMrjXiHsz6+vr64KW
9gTBKnlz2KYr6p36bkymSkLSoKdkQr5+jqYGVue5dZIlBKcSSTx0lpG8IThL0g4T
EULgqS8ofJghAtR4/YHKoA+UhguV9CeFw274iQU9U2aFnFIgXuyHsKoWmuOkmgjy
7Y1annm55Qzxx3AIa92yJd4gCl2ZYXj5oeCRdTlveQv0jmjpzwXFNWyxBD2JKVGc
zb6YYykXYjVCEgzkd7HKhSFv2GrcqhbFCNSvo0PfdteNAsOY8ErOGzYMPhtIF8t8
QxaLbRxe6oV+MVbNEBHRz93zJfNztRYFjprzPs4wQnAcYys201cfjmY3HxVO1Lbd
7pqvgnrrDbwPMbO/e4pjsdrfkS2xx4dF0ANWzqSZ/qtDNSfaC5RvphRIf/nSox0/
AgGMUeB6Z9s4OIZc11P0AxCmJpbsWihvMqm1Q9OtGFUJ9uH8cOL8z2/yiBp+lKOH
79nsLRa+6lmbH2GyLHPB10AUnL0XDHW/O/4wi8Z03gsR8zbpGcnVX+iXFbPcT97S
XD0j0p+A5lGAdxTO7IkY/aNtI9+CNY1SYVwU1n5i5xmAvRsOmHKmKLGfz5NCPggI
d/bSH5oMIxYdM6LZ1h/ohvzvysrLIlrvwzxc8rII7HnnhjLoj0Kb3yyilqZAi5sC
saQOwTqgvMHHmtSNlVJTZEVmWIn9YZ8dCKDxtWNjZ/iErlMjsnKjPb7umUT1EHs+
WoiKT8GjDNwyn0M5hSNaZdULOjwaIDOz5jrI/t4r390YPDRfwvvWAr7YPyzrKzic
xsh/4CUE/PavqRTLEYlxddUyiLdR2QClzO+bpNaefZQYwx6kgkULr/FWkdv+oVnF
WjNrvFOvZx6mgUX9VPyr+GkxXNkfCgOEdzF6eY1QkpnogMVnGskMpHkT1qR2JIs8
expywBGqL3qDrFO3oUXvv+SVXgMHmei25XMqGBuExPRbpvbiDzDorqpV3DjUWlXo
l4bRXT+vD3O8QGqFJvryhZM/hrV3Il/sCEeOd3owsjTCnDCOpXuql6XrXLSpz8Vh
FYn57D5zPfzerzsgl/Ifmo+Zs/Mtjq7cDkKyne26hwlX/+DAQsilJQrymXom0qQ4
jbe0oRAqfdQFRbdX1SKEGj3eAw0xYNOtGu4DPj4Redz94l4E3y2LB0jKPL+yaxyL
Yt8RD+spl6mJO7Hgwdww1WgN/IW9/8kKlXW2L7hmylTtAzrQqqoGnDcs4a/rmTX5
HgwX0r9I4oDARJJe/GILXngGXEOuBH3QZiO29GEQHjz0PkLXoL1q2FXvO9e3tWBa
A83ZLMSBkSuOaL8KES9hc4Cakf1HYbo9gHeVsYoQhktS3BXpYTx6+sSNKUiGwS2e
896pPYXCD91SM9/jy+7mq2qG5CBXZWd6mKXA0T1CCznS86HEQwLZfcEjK4nqO83o
C4P+D8Zcz0OPTYmDsDsarwQTPKnZ7lmbdmBAOXCBFCfSBGwKvK9lmCZOBSycOUpt
3mt8iY4wNmsi4VZIsLkX3vEKv7TRuHGcE52iNwLNXrVOr9gJ5ol8xP6PntDyU5Yq
B3PG3Syc6wXJaGCxFPyiVfAVEGnsYib+RXwZ2y3JnBpmI7ac3XhEEoM9llCMXEsb
OhdlxJ2nDWPyyI0+fTP4kKMswkAP2thfo8KMd1okN6R0DjqObb8giYV4YuCJHwYx
PUnnrBpRmUQNwBMCfW1toIHzP53UrcUb56dzec0D9ZA7Vie5WRYoII59wS7vwAg+
SJr8WKQUHG+5U79YANl48ric4H579suMSNhnoltrK2ZI4oim8yBtQZYgh8xQCy/7
1rJBp/pru0qfEOQbnYLXn75Xcq78HxKOcsLYYUP8zbScu7kg75mXAj6rmGhxgcnM
Us0SSybiZRUHLFAGhfn9XmMTxcF5nHbR3Pu3bpQjQzQ5F/aXJ5cWARm7CCySBaQV
5OZYsXdsQwwFA4VMPAmFiw8SgOOXXvoWsvR5y2DAwZbSw2SDFmu0mMcyv1UckFkM
BanzyoaYGrnJepMnMwv5Krepwhgrxhg+XGs7oGur4HbJTJvG6E2S3DqtZLzphgNE
lgDMMfusgmFVO+ZaZYCWRgNcxZk659zpF5+fN3irh0srPCdvhkS8zd57QlWRwKlv
Kw9lngg7xAFO5WNp5u5+ltDAzYa9nSHJcFzTjqMBbWd8s2FROlRAEn/+KR1Yiw64
OULHdXY7Z8dbnQd33IJxNmdJ5gmLEl9MUKM23UAfSqQln8ddQFqCVDnYCcmtu1rd
lD4Qb5SgLrkchApadyVcCwJxmqCx33qOArfiOCLiC9K7OIuwO1mFsZ4qRixNtqir
Wdi/4pLBd79TLVXT2AC8MBNM+6X/Vfs3catNIpvRzuuha/0eOQNlTzNOS/K1EU2T
u/VbtUQlgY6N1nALZEhwA27YZ4nIgAq0sLtNm8LMCjLSYVlhp2iSJU2Wumhkn3Se
LK01G7hte4HTZIg1IuW7OCxN1LyeEMDzmg3LsK7jc89FzomRHUQpudzXC2ud5+/w
stcG4hFT6HaeVl9OyQwVGWv9qtWe8JDpuL2aQDU3RDaJSf0xjTarhG3t2OycmQcb
cjVWhHqKpeSUWmqOThbZXflswIKgoKJFDn8kpmjealhp3wdSPhSXvSF1B42nd5/I
5eVMrS3ur15NBG09RgFI6qVSPSJX23REtbz06AXsxfhtZ3nlBS4r8Bg4U6sx7esc
u8mAJNWFjt4+LTYMcbnnEa1w7oeEEFK55RZeq6U7aHf5JuIFqRpUTeqQTaBo/t4o
CXphDJZ1yq6AIt9AuplJdgarqri4bX9myrFj8MEyoyUtAVFALDW0BQMCk83zteWP
JxdB0DGZ7avnfedSWWNANSEi6jmzJAwJdYrj0QTd9kjviQ59u3UGpfPYPNceY3/O
AUEhCF/pEVm3JW0Hg8lUpR2Bqd2sWjrEKY85dWqDR8uNDOv6gifxwLc8a9xEsATd
NoAMjgrK4LpWo+JlqtSIEHqOhpIqnAnvU1wP6MkerLtkgmEkZ8eOK8MY5RmqtxP4
kNa1A7fSG0TfdZAUoV3aYP9aqy9G8Hc4sasCShT3zu8wStrW+izTRhk1mekzOCLm
FusmWdbyTFTJSJbPPe+WNgGtcxnLDGfNSax/BBu5bTuKw2551YewQdGgEYiYZmPM
yyg/4+OwwFrcCCPu3DPzh6qHN/V+SMaRLY8sy7b0tht0e90662xgCOrE4LAxi7OL
6uYw8K9ng3qxq7jfK+iuQMSOqJ8VQthmHkVGvZoACz4qUzg5usVR0m89vhwszrke
Lv/3MNrrU0tYw4nj9mcMRbHWJxBt8cwH80bwVCia/fdOyUtq+0h3vp1hRVodtfjx
+2UIxrs62b+4JvGT4eNedPrI0bKs1FICceKLIQGT3sd0pOEqN5P8kude+AIQLwVS
P12IYxy94qDZwTxG3jGou6ml2CTMA/19z0CT+9B22bkJW0iCE+G7R7u1HW3wbAW1
+cuXIvgM4MJLXPxLMqZEH5+UPsWQPnUmuj/kuk9CXip3gvXgY94uDT/WRuQlfldE
OroeEPXLkPW9tNrV1WyEw4oVxAa6R+c30jIJ4HcwuB2iNupyOAhrHwaITEkBeR8D
nqTDxV6NPtBvsIKMi1WHUnvfSCHr+My6WbWu2WOogDaGhKrNuO/CJQcVeEyK4CPk
OWYqvikO9lERI7Xc1YacjKveswQ+Ghhuh0PMJY0nn26JyqFffJwBOoGZUifRS1Wn
yhUuKKX0FnG36paa065of87Wu7nQdShh9NeJaUuruDo95Xfb2ZG1no7B7vv6cz+c
wUIcPHe+Eiyo/nODXcpbCu9p+iwcxZ5hheLIdDAt721n2knMQkZI3RyPf9HdZWNu
qv2u/aYYhu86FHTVBUwo2frIHmA9tVj6I0kAWdvlQEV+mQnSfrnHGWpQiIfhvqqo
uBI3dlmW0haUdG+Dtk+ZzMgCOjvVn0sveQ0g7jrR7kQ3ZZ8gLzbFI5bKiJDtZamE
BsAKIa+f1ptsNDZLUMBo3RCmYoWjs/hXNOst3HPYjUNAnNSyPuIXQEeWkzIvJ9xQ
bL6Ddi36F3xjNz3hSVCt30yiu/B2mX5OLnVqjzJyoUjaoRPPHKMkkPBZ98hmHTRC
6F5T23IkyTqrnPf5Kwd5+G6Nn7zQ4z3QPd4/D5PhXM9Y9xcZm/g0hESUy2AHHZhJ
ZQVI5Y9P1CpbI8SQ2Zk69stIVehur4zG3XNeVO51CQerfmMHWIXI83n+9MretnZj
WNoh1xmRfZzRBnVuClaHfpuC6WFPs+OBNzwl2O7/EnNe67zUfaSjCeC8DcOlQxdo
7RQCZIicpYt5rOPSpX+SJmuI1aYSgk1XgE554gb0+WFbbfEBJdaFP3WXaeef5ZOX
DHxpANDOUhGEcEBFjF4sX8P3DUHVS58bF7lSJI0gNRxLVvTOS14AoRPByDvODkJe
AnbWa9Qe3z3nV307lbwtXrH9TvCGoLVfpcnN/cwF11eSjeIIDnI+piFJj3mP2mK1
AmEV3DobQ6OTUxE/MtuSHmD1LOAeK1qrWXUMjZimILA1DhIIiJ3hfQ63Y8+gEcen
1AmT4yPiERettpr9D7lv66tA7pAGkm339o/bK/NAutK6SgfOCL1kJzLcB62IB+mb
9bWeSnQPaeILAdVcSx0oO+bK7U/R/khtiTNu1jbzsBSzbWk2ojADs2skydTBSRqG
D3qbWL6Mp0LKt3uGGk1j/z8MrWzZsjYWjJMq1FxoA4ZNHNo73YkrQzc6SqxyAqf0
gKbJPhi5kzwtMqkiZB77y1NJa3GjGBBT73mrNmGXy9EC61SpttaiA1pUVtDJnyRd
+o4NDIYOHIXSsYJ/Pcy7n58OLuFgZvMZjZWrmoK6PGCdv2hS9Q4uNtBsh6XrS5qN
LDeT1HRO4Jp7hc4h+PP15HPj6WfT00opzig0GYMSl2aNXUZE+SMjrlfLs6H8wtIO
9FiIfabXqNdSRz6vApbdgG3pOcW7sG2feMZLaCit2hWWCc8GwDfmQTqjwmGuir9r
jTkdRGg+cWgAjtj4yjEqrttKeg0CX6jb+kbFlq2k62uUQD8CXHIHzOaXHIZ5Ik8d
mlWMgC/avPXIf1we8d9m7ZR7YJRu3w5yRZX+NHabrVOtctijuUtS8Puw+jpS3oN8
CADT989qRSsMyVyvCmMyvAyo0dk9+QOp1Ged4hvbw8Apx8KfCi56ptMi7qYzgNGG
+RBrckXiWzbGPDj8x7sWMTl9mdoCwCcnx44+D7uU80WPICu0MUdLhmfRb/ubIa7i
H+wgj3z/CNVqSsKEH0TDOYKeWtXlkGYQ5eSCdODOr655U+vjTFTn9gZNN18t+zQF
ge4ZsYHkKy6SBfAPVKDLVBmtQFYQ5SO6T9K9R4WZ2gerjEcTIwjeCjMzT3y3Bkh8
3xsyWEBU8XVX+VsKSF0XN1k0386q8nn08DQSRKSX1q1ASZmDHO9mrN5l5vxRfyMR
/I8a8pCH0jGU/DSOm3IEoyV2nsPzIzw+AuqyEIEbvsx4LcKu15N3No83pauCLjFj
s6zb79GTR4IZi6kiBztCp02FIt/72e1qBbxo5GB0G+F55tw+bv5pmU6oyf0r+eNg
dxXY5PXV3OoMUv/VrD+a/SdkKqYAqXX7ob2ApyR6XC+MGC/ySI3wg/Ln7ZCglAfJ
Sz4fxCBgnsqQL5dG0RgWSdMtZUOXYCth7clZuLsGjw382XNbqffe6V5/bvGPWeW3
S82xBqWoHVYSUCjUawTA5D9eHH5oJxMYucifFey7SqAyIOy5dgvpLd0JSeznwtpZ
cuOzwSM51nmU6BOaqK4YoM9SlZvSDrsz0R5fd2lp1LoNjRN26UiLUnqOwRN9gATI
+ne44lErrew/J1JAdVWuxaNRogtpxe9op5gudLB2R634DAY8sSLvIfvFcOZk5/Sa
5lY8ot3qlDU+0m6ErHIekQIiM43XaPQfKFfocy6xYO9H4Vg/Pjn855BNtpmPhbbL
zFrVRvfQyaeMGq13wpFV8bZqWf4VY8ArOoxCZiVEQqQ9emsxC6LvEUwCkBj5kDxI
2eIbAcrScIPGLtdW7jTumGKl+UhL6noAc1Mf5NFuOuOWE2XgcDAkTRhEwUSIvLmL
HVFkfB5UNoKZ8A0ImUruOcBq395s9Ysb8nDlllIXbzZ0FHCXCAnvkRIn2UealCgM
HZRtCKbdR2Ym+1Ypotz3es92rz630Yxm2gW/C4KONcQ9RqgvCYsEPznnqm++gt93
mZioakuONG+Yv4J0MCk7y9k84XQ9kF12ESSa4nOHkg7OW4s3pIBqdxwj1HDGrXLs
z1ikYAjEiqimZcyjN43uv0Dr9kGxKy9WyddP4cgbIWCy3VRO+1bTErU5iV1b5F+s
t8rBGo1t672tinIMFVf8rtj4130PBD/gg0Ml381iNFlCErZT5thon4dCZZSB50H6
l2nEyAwozmRqrJvF7f9ED57Acg8kktBTBAVX9UAnpO+nKk76KSc9nZghvym2H8+Y
AG7OfzVkB19IS7+zixKHOF4cjDZAiuA8RTBS7x8peUrQ1CcUEpROHnzvBHV72VHo
GM0AIrINyKyUNz0T2zV0FHlJnfWijD9dSotttse/WF04sJOxzWuPFrsbpspZWinN
VpQelrTt9NuAQVnTSNZJ44qtBbGptNUoMOvXaR687v98G7Mm0TUY+koNQIHoO1u/
2C/SzbnQw6yZiKisZpXuzHbZEI3f1C+ylddBFuZos4w5eu8OGufdKwsuLGXXjH0L
97nZcmxL0yjZDW3/TMqsAq7Q1bOIC8jYc1F7arvdjJ8RrlDs0cuvWF5xPLiU1GYF
La6z2CqJsPE5U+KEh9VW4MW/RqRs4+Q3PyLjsX2cMF7eWJJTymaFU726Wm1OYIOH
2lDyavtckYChf6JGS6Vr+5219kGp+3I9FtFJmyp4HWqBpUudbag1FAriaLX/do1M
Ml8LHq5sw8BzDQz2CczW3xR4antUwepJfOdPUIVHaJB9hXsFUSqtlqpEv4BWJ7Zs
td7TceTjhs9Ze4nImfGv65LlUI6RRRqALt4S1X3CyQMR/h94kacq22ZdvNFz/c/S
oJNWbRWLSJTF/T03uXxezIZYOGvmTC07vbvsJY7UWSbB86jxBm+RAdvXOswsfzJm
wfzNE/1wA1p26yb/3ff9WCv8qjrm7ed39SR32QoM4Ix6uvQlmuLSS6o1ow0nSecI
5DiAvQNeRtormn7PzROqRphH2V8eL9Glfr1Myehp5OWCJjycyMTw8L1yw7G0XFIy
oPPGTRAgcb5PWzeoZN+s7jqVQ17PTR/fK7Q2R2wx3gs87IiekB3Jt6pr0UQWVrLM
78wji2tnOWF3wIE7fXJemrhZFopunF7MnMBx7aJGnrkRK0dvF6AnDDX8Xv9u4n/U
Ao9eEyZnGjbyLN+ihlB4NE60KL2s0Hwrkf1QJq19cyzcJ7EFDUz2L9lDBCza7zxJ
W3OodD5ocQsYjhDZgSb/1pn4sxKwew0ndDdqBv9tn9oOAiW8x9v73H15Se8V5VjV
ZRws5fYXDz3p91JGOjkLtGG0jwPkT9iWPtist3cU52CimMe37xw6vBR2i66o2v0K
ykNqitlnO2kMKcR2oDYUKCv2eIIQ4vS1q2rM0yK/l0XHjOmPFrvLfiU5oEsilrZv
pHRUp70tbUT8CxCHxbAKibzzbjG7KwbOPh07ejsx63nXSUne+OJrVr/1M0Mj/dNo
7mTVNy+VHrxRWqQvyPBMT6t5JqboDOKQXSh7chzjcr0vGQITAstQb7WBQi1+0aSf
tckVhNQB/wKmWq5T4o28CIcNa176pYIu/GHwCgD+SD7uS9RO0XpPxeUfa/xeR9Sh
5rQfJq31ekXyLAp0IcIad4I2KpbFN2i4x0rJdxNkhUHed8WBgkir4/zQt715LT6P
wj0SUL8U0+QIQt/kz/p4oJZr04xXn2yl/Ig6+MNU/6ogzt4HQbY8jpn2sgDUtNxB
mI0QoW3/8nJ0tKaL8etyO0AGCfGSOCEEiyHeMEBxI0UAdrHw5cEUrQOvIlKbXLIr
jKzdhSTIAs4+7jT22rsB+VZcxrQ/5z7QismiVTNxgXWlRV8aN8pYePfLdfnwRyAm
amGepxWu+LuE/c9subvnD9KXahiwwzSMRLloXs1hyLm1bq8ggh8o/i1BsuqhiWwf
2XEi/khpROGEqVHSmLD8AGmKvDIf1QyFrkDyTPTVp2T/JuzaB/7CsM0T4UTwC59l
lE5vmjsU3+sBhkf3ClJOntfIR3yzOeSO51PTsaPMkzUUgRJBxjW17GfBWunAeTi9
uQUvU/bmiPgZIrZa7khP+9R5C9HxNCm4qhUDnDSoeOzscySBzzFBRdxqq38ms8Zl
wQ5QD3mpgjsbMSPCWv9wuqrF6JRFn0wXjoUAPtwkVCpeNjvGAJA02ZzSc8/Cy1UC
acg2KS1oxtfF7O6rY0p9Jl9e310tPkxzEYl6eB7OYAa926kZOJGt3+mRi7tnyXk1
op/UuZP3gJi/9t1f0MgvEa/mKA0W/VsF/wR3s30xipJNlLX393iWT+NSOnBh/qVP
q4EZRrf1vT9iOSF/F4CBp/bYz4DU8TBtHp6QuLmddWbgksYfKrFD2gG4q4YaRBAb
o9uAJaCuFFbhtFGilgnaufvOA5UuL+3AcOuY3COeBWLgAWU2TEtwIDd+Ac1F+ViC
VU/GDHdqrb6QBJQLX8Sb9OIXviXaXQledkGopduiHnpNo+YpaoxdeQDhBgwt8fcj
b7uk32+iw0fLOhaDa2zam7YFVapo3zE/n8B7rFid5kj6vS76oN1whzTY5+kArNbA
hKhJJMNrBI+hDjGUps0mEWJ1GBjVHQl140Xxvbk7ABjCgGIMdaBEDGXpjIKIefQh
T1SkwPT4mQABvM88FfRQBVL8SHFsBrMJNncXy5SXJkX22odYvGuJPg1PazwVacbn
vR+/cBuoa/TwTRySlBu/Qb6G4Cd/mi0em7f5I88YXkaS0KTLwEJVCP2aVVKc8a+a
wGEY0Tmkn6BvM/RBW6b7cGwB4RWIDprCUE/1280Q9LlnNmSfv7VuccaA4tCd2Zqs
lNRG7oiAQ8Ut8+eAfQ78RRwZ54xSiyRzBq3RkT3S2ACtOCMxWtgTZ8qvbzHLsNcQ
WeZIvsEsymap1FwQT1Q/JoMZXrwQ+QyiwYU19YCB9VD5XeNvwYa7Ry1StEzGQN6o
h+mnV2QmQIzXoLz5TF5QVWHmQfgdKDERDR0UeZYazK4nduy7aG9ht0R+tU3uFl2u
Q2VbdzdiH5m9gyawTaDRz//MWhniqFDu4nZ1E9cqqPPuLOBrRFUPcCbzEdCwGmBW
LfT+qEElIPAw04uT3xMuIPgbHLKwsh/0K1NUmaECPMk764gh96dzHnsR+jeRjGqs
HRFLjX5lozfKYhb8rfXEiwq2Hwuf6QkoCBNITFsN/6ucm/OMbLsIpsd6dBP3Ympg
aAEnVEvgp/tR2ugEb0WXJQ2hw9jRANv/Z16BFmiD4BUeK3jQbpz69TxQtm7UkayM
9hRTVlZLY7SUdRdIVxur8dtQuUKjc+jfAfpBYV/EbRTnp5uFmV+16nvk2doBmbE7
/R3a6v6xeT1zeiTBCjYffwTqeli4bXXNJuBq4XN+syfgtTI8Bt+0N634NgfjLQO5
7A49PmCE0n9ulw3t81WYiBHnnZbNVXku+AWLZTZnoQgYm+eJIiVjJ7oXxzDBKu4X
IfvWQQAQoyEiIbaW759mHHZQ3xVXKPR50SKBR0fszSnCRX4A3Dtrhzek3n9xYVH8
K9mWCff29MDMHvEKbyFr2VbbSqWlyJpncsHdEm5pmBGUc9VoTyMFA3GDAeLFFUI1
EeX4+8yblc9p53/KEh8i3+Fy8w6X7B7iiQoYHEGiC1oilqlrp0K3HP3YZ8Lfb8Wc
lX3uH1AsX1uv2jIkBJOszTCTQ3aeb6YU67UaGiD3p/2aOvEOmbu/1zmUEQjKswyx
g3YemDZA4cdqnWTx17oVcJBwdIAMlMhasvRjptDqqpqPK1aFUJDts5nIeI/F2yc0
t6M+UClq/E8vdys6U6xMdwA9UjIOVB6qAD/sDmB/M4YQYj9G0oBALuUQQOHYtOBB
hX1z9UtJIv/DboC0ctXEgGxH2dJLfqivKpv89lEJvzxXf5STu2o1QPwtG1J7Ma/7
aLliTbJ6uIcMtbBEtFEswSN8zD3vO9l5lP1XxnDGEeTv/6fKmfxFQdTg0iELITvk
R09zy7YmWWILbbjRXISHO2aTnRRvdxfWPaxm+LtrtWW/OVlTqZIzL/xA1LgA0eDh
MTdAPE9wHe7ayjquLV/ujmBErADvf/F/rduWSNltVl7OeB3wS3hmS3ukdjy5DLQT
qINwG3WROSEDF+zTmqcuc1Ei9SGPmv72TLfSOibaPDIkPoqtuKCr20EMLTQnH/iL
aQes0v3kSinkmmCjK4cFE3rBLmjXsf4FNvLUcmlf19U=
`protect END_PROTECTED
