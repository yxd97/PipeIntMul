`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZSKPzSOkCXuRKvkBxZQUHdhouj/6YbKBHcjPH/ZsO/9mDi4zqNz0l3FMOrUmIJY
PGgoWi3n8vuncIKcCcZJswUzm6R5XNxxwVu9TwEHpN0dcJnwtt3oWCc1BPiBXJE7
rQ25s33xkm4/cXDXEi1keiupNJZ8PGXg6VToYq0nsX/OLQ7TDG13u75/raPbYS6g
IiO1TUdQyCPTfGGRvOD5/etnmrZd/UILR+waM17T214LSUJl+lHvyO3OCXMCrvUv
O/Rm9WxjjBVS+5IChLuL1uX7gHrJnF4Vkqb0/y0nRwkzBo4GY8xmpzgtIDfkwAZb
RKB1GPlzjBRNLT9i4zLwGHkFXB9zaDxRqT1Or1+n+8q00L1w3MPHrx5eA6hZgRM0
nfLXuTpxVDIMwNBs07uPTiwL2Ad4G3HMcQ9NsiTv8ZerPFFGCP/WqrYXsfY/18g9
YESmsZNvaDEsi7OcJjHvkvL6z9oQo0IjX1EEQeJQR54o33qpXSo7ONJPtM/LKMJU
YimmBkuVi9zPNJPE4i8nCFO1i/xu2XpBVwg1qK48CAcqXKnQMVIP6TbBvEluaykb
p2XCsfkLWmCvuPicCx4rOwjN70dwddZrOOYVJ2leMtyavFb00W8cTC8LgT82/fRt
w1KE5UXQaOd6uYEd4pBCrvD0laTJuwHgpRCaVHTkRw6S0ksojT9smfP5cPQMSfd5
tZ1OMmDEkmaf3fGyPTNPfRk7T1i2Fgjw86X2yPzKhW8TkrL6+2vBR47KQt7nmlVe
bX6i3MIPSC8qQRxU3gVT2FCSJ1jQvPqeMUPW3WJ/AgPXtwCYGFD5wk+e9oObDChK
R1boGxihuP5JWEZdoFK+g2qYwds0NURoEJhgHU4YcQ9RMWrWSPVcenhngI7cxiNk
SoWQCWGZgJEkB7Q30ihyX2mbYAytbaBo3tnbt5Orw/cYWHK1bNG9zXHvftp9iohO
sNx2wUv0zhXc1xkqpR7GgSsNJ3+aoHrxIuDnoF3iTL96pXsNITcVLLkX7cF/imif
/6tUYjXOqiGzuJ1gzZ3rQoHhb0k0fKgDwdtIUKNejRtD5sH2ed9CPU9J1Y3dV+ZB
SMMC6oWyd6/w7AeOm9EWLOf1ErjCRIf+tsdjEAVMLTx7Pn+/nPQy5uBf6QPGSHZl
xGvvOqYES1t9u/mFCD13FipaySDcguQqB5eEW46Xnm58cnMQSKDGY0qUIXDJR6Pp
e6InUsuN7ZKDhN81VRA9tP1OKV1QPSmEGfVZZy6R0KSVgxo/4Cb1upcQ/dFuRddi
o0Uv7jCaULQm1X5z4R2ut/oK4OzAbxb5LcFXldCeJyLj1y97efvxwYd8ZM8HWVQl
x0AOwx9CJVGZBB15hN3c1Nf32lt8b13/QK5By/5yTXKBbHTKcfA38hBgNvs7wRwk
AyQaMihaGQS7xu2FYjwZr4ua0UisjnODp+jdd2PhXKA46lSKMMQ3Jl0oSsreGo7N
Uiw8lC+FOohYOoCWy8UXEl6GrItbAN9xw6c/ChCc+6lL+eIIzvBjwD5venDWjKro
ak73kWgTrHBNHQ+o2IwQ17tc/IZD9701dyPlxWx3w2IRYsYiancjvgAnqA79r6Gk
Gy5NDCjS6apcZRUkqIhoNtk7zJRg2MWZVL3wKTbNzuArAO6Zhg/KyVC7Byjcd5C8
bhemN0bUQTMspUULqN4Lxhtdv3OM8oH1oZy9UA8Wj9zS0PWS5aovnJOI6XjG2kyF
c89AjhYEhkLT5JyxKQfd9mcOiBLFxXZ9lk/zj3jmK0YB7yuVGxqMQex3f3P80Bcr
7cOS4MbV/FXVjN80TmWevdxuqS0P50ulJPrn3rPCuke2p0gRJEqEMIW3pJbmYn0f
MLHxKBBkvaR6HiSiBKeqmR9lJBS/0pXiYLXIveZAZ9mCT8iT9sv25Xkv3Hyr+M8W
Cn2Q5CrwmEuBMklZOrRMISdngrsiehhMoBExvLc8DGLD/Apm83HbkYqwuCIVdkey
Faw092Xk3+pOaA02qvahqr7T90ydzhbMVo+zRhX8tKagZo1mB2ynyKMsXTGx3we4
BmBB06lk4HY2Erg8XczzQkh5RTdz42mk2t5QtIwR6mp10DBNwSHvgThQsTU6hIxS
HkgtGzgKdjZQZcgXIWe3R6ofH1ZbmeFzI3kvXmHcPogfdiSoIkUbeKGUDKFjSF27
3QPNyJL/kE49HqSgNpeXHf4sw6WL89mAGfLheCpzMGsDDnaTr7+ZQrSJ0YadlYiG
5TK1zMDbd+1+HxESCm9FubzKwNjlpSADjWT8Fe+zjyfieiQt5HfBslYqQxglEWX4
3lb9TPt4I/7jH1m445VcqoFcb4SrbzA2B8opWje44JGj0FWIDqzyZBEz1Fti6fAQ
81X+8SRKDR8tRULig+A14r4MptsT/d1baWScmasjzavClEF/doJMp2trhemF0ETv
H5UPjhlzMNg79SFTcQ6n1EV1hiseORe0W4pIxucxnQHyriziwano/09CoBVA0GDE
jumGvh8Lv0ncI0pmcEWstkkNNYScJvX3T3Pdok/Qr+2/wYNMpyZxorLyuVep3xWS
X5efVEXDnukiW0HWQaXQa6YDkmhSPQ/TlVBITFVMtut/+t0sdS/022e59/JHWAvo
I6WcQ0vh1MYtQ5Q2iPexLjWEdShxbuaGAQhohTiLdTF8NrLb3wKcGQaDT8th94af
NV1xZrrKTzwkDICn5mVn4jNLSdikJqH1RZDrF7oWM4QpzV50Eb5O1mkzUc9oD7me
tRpTT71LZdONtYoJ6ogZ4gv5EczsPzdWzNvSx+YexXfQCI77PfVuW8NWrXstEKak
wdLCZbgwZSdU9mBXBruwWRHXfpLiI06RkQ1HZb5Td9rxXhiJ4nvlE4r4+riyNk5l
EBwypnK0wFz8Yky64hEB/QuoL9KugPScVtJpAk6bKivLuAkjwpsldCB9k1pbHdYm
brL7KbO9Nb45NklruJvCvfaM9QD85BNpeL+Thy2xu9h3cNj4K14BQSsv/7SMyT86
7BeST6smADh0Grn9iWQmG9woZQE5ExGJ4vIqiCsSkZ8HQibxIW+G/4aNGvgnkFVs
LK+0QlL7utW5ToJ7NFvMM/iMIerj+/GDS8WfSfxVmOd8YzfgVoeKzvVujk8/iSXs
jI02/WZhY3JOKN71vRycamGw43wbykjth5cDPOuWmXSmYUWoQ0wcA5GoeKCuBQ8K
OejcFKcQDoBoef1kSO5fHnvNaNyRnTQGmKwKik9+/ZCcPE9CDFXNXJ/2HfRNxguy
UMaoOZp7/4hPJPq3ZJqXGyc8b5tKq2SGlT/soXrd1/BN3ct4zPGS765JmbfrkmJj
NlzSF57ChRTrtiQcLP7Gr7YADy0/wDEkFqFzEQU57UXaBFLn2nrP4Gt6U0qiE3Kf
9YueAgV7Amq9rNEPPesTl639NsWEeoDwJsbmMfRhDnkX8TkoM/gxTKmVrFVmDQwh
5arcbfciI/Zp17RHUa68llR2fw5q2t6twUtuISRuosgDeJ2ze8Ig1BWOsr0M0xr0
AJIOfZOYyRzjtWgO2QtlxAZvP3NxeAOHdPN+2+ywD7su0pFtCO2XIm/la3grf9Jb
q4i1LSxoMoCIpptelY75lTOKcdktVG9/gm1qS6xu6WeZaOVy87Wz50UBxeBjExba
CggzmwJxKH0zS3miyINfWjchUtAURSpaLwKbv2WSIwV+JaigXqh7MEG2XCP9EDHg
DqXkzucbbyvEDH3otuwrb8DYh5Wu2Dt4riXvKv+K9avbVde6Fc8FzOXanl2wzW0O
IYpCagwIwlcN9umsOO6nqDiZ7XbmiLIpScmTpQL//Twea+jWHFr0BHjYNw7UtRPb
oI8+HktXP07AMyYCrtY8b3JtYuZmOgTR7AwKUcqCqdt1ojTMt94jANG4NOgyfnu/
E+tfAHx48KwyDV3av+rRFlxvvRxhlMBpnNbAT1rxdYCHUfh016VQL1NdkttOOv0T
erH+/Krh1UGezhM+N7rdAkMrYoLX0mNmGVVhPIC0zjq6eP7zZBQ6M9iMsBOw8c37
TItCQ+QluMs2bRpqBmYVTFC9uUY0AcuzPfBf5muMyKpKDnEHBDV2rihydbc7N5Rc
rwDVoUYZSjrU/Yvqfr+z0qCUDF31sLQj2zu6zsBKkKhPxj0GB3tf+AYHQ2P1NAhp
pxl7Vo1gveIsiuysvnFf95FjlH4xbIsJduESCc3K7oRsG7SYWJDmgj1+e907q589
YwhvCEpSqkSIhglsoLr7gXt/BTFqF5orq2URxiwGXWBnveFxA13nG8bvVsukW7cO
qKIjmvVtaq1/OJN6DU64hK/vWRy9J2rpYpcwliaq+X4TaSe6kxQudtWY9vkp39nF
PFg0ME7ckY7oqmYitKhgvQb55pyV2zl+TlBFLOMVmGOKFX8F9/QLsakI20B1gDCA
mJVA6ZrMw71h2M1Qg2VggsVTxdq5/VbGP9oplXt+7LjoUWcRM7z4P1pMOeFvn7I6
NLe2RwmN2qw+ng9RBB459Tny2nDFttKhryNTlu28OHVnTYxYdURQKCf87RgLuznG
B47DZkO3+juGY7ZG3zREKHIIy+W3G2zZlxuNL9EvuXZ1e2H6m18s4YkuVwjp81Hg
qF6FaiQRamWu9l635fRYqn1diCwjoqGvPP1USQJbY0h9CoMkRMyGJDMcH4LDbwH0
irfpfLde6Wfg7afNKzHCDIvipbkSfgjxQP1icxOpPmr+Bk90bNWpZrPPXP9LEl+b
zpH3wYcwJNVuVhy4BpGrRcG2zxZb3bdfsHHP98rTtb23NK1wYnc3lrweBaiAbj2X
2wdoXWaAEYsYjcebHGTlc2/4+K33GzHIa8v+DstTs9jOL+i1qvE4gM54mscmlmpP
GVbXWUl1UEaufAGZxPN8LQWz7HdAHNdo7bvrYSvPqy4Llhb4KQiC9dVFbGpVEfE5
HnRmfva1eO0AqkcqfaKDDo9P2NWsICdEqBMJnk64ZpLDjWREnpd+X6gzedJVX4dB
JogdAKREZI+lFpi2o05iGJ4wTIs6UGg4+PkvV2IgVWgxcIDRkn2i2m24mruPp19q
vGmUGLRfGHFMIO0LpDxdnlH1Hke65vgvbAz5q0aqmHZy8Ek6O7XxOjM4jv/R/Qqf
EjBIUtC4X5e+gyU2ll6pHzdshmI+fc5GY0NHFC4ut04tYXWnC6W3OASuVej2FgpN
hgA62+NbwjJ9d3Moz8N5ofqiAjK39SOd8fIEb6zCpto+Z0tTCmfB6VmvEUZaHvCl
N8AfQ84zGnYrgppZzqqBOz6oJvD1cux/T40Tsfql6aWOl41z4sXEQNPRwgFpSp/l
caZogD5YCZKcC+vQqT79fdNdO3FNGeMh3Rg+44g/Byx+e7KnLzBJgjPFu1HXM8pw
U/cr2S9yiWD/L5bIqXH7g9DI6YN5qXC3Xf7ob2f29Jekdr8FHJl0s4Nuv7115YV2
90jr6aUYChNHwvPnYoQivu5N4XbY9fnpg3nNK3bEcauempchP2Ek1QQZqZSuCLQm
CtwdZVsfnkA3Rwv8V04HJWc0Oz8aD9cy4oMjqWWCbBO+MO2cN2RxxQC+XVjsIQ3H
ozW3Lljh+8IhpA/RKBsE7uMW0Xvg7lVZwQ8w36NUeXb9gEwbPaA8T5MyI6f6Swaf
PPUR1EINrMatZLWcKClHK0Kq9jTc8dxqGK3HCnZawUPMqFnycC6XlakeidBzp1UK
++0i4lCUC6RAzMm3ntvXOJAaEF5mr/+nJOnG7SIloGcFuqgCl9Zxn9DMFTIkIFPC
xUlYbjRTb2RtKwsavI/INjeDAIcFlS3TxCzQwMNyDlFzGwfgWMfojHbM3C9Y5Tsq
fAKZGh1/dGynmS/eGAZOgTZ4qnw5o4wPyc9N5kZ/vaj+WriQDUvRbIbpbU2A77IX
jlPZZxtDlJgToYPx6qxmTTDmxjJ50YhjfvD5mXb7dbCLnLYH/6dwhTOSvibicthW
ITkZUt+1hyhEjLR09hCcx63avNQBiumR3yqpC1oWfgdt5HraMSiMY/aELeB5pGrN
+bcqYNdHG6aWRF8HmaQURzAtpLwPWyduXoOki9x4TyPRZmoivX19/BCxQRtfeF/s
bvul+NZYXNr5G2MO0oyxq6PD95l6M8tBKtnB7hwEV5QBne/BNU6R0Pga+NjH/qo8
kVIASUJfn2MM8EpJ63w2ohKcO4Epz+aQabM4Ex6kMXF1vz1q16TI6YC5cYjrx7YF
TtP54S1o4FupdkMuEa7GIh9Fz2kdol4Q4F2ESYojpWALZJ77ldDAQQ79CxvmbCsg
fNAOBIChQTC0/PdNEatSWo60MPfwLkBy94IDurdlVwgNYz2W5BaZ5XhSbdXBU4T/
XEUywS0qIMuzAJMsLH3oc59AhtumvcslpmXgUhiEcINEl+c015iLU5mvpZxex512
SgxfLZodlbwfAHMwgOzW/9hV8ClqgmmGP9nXDxyHaGDEd5PscVya6c9N/EVGZ2TK
vZS2qBAHoWsejJKFtYx7Zdq0UsPBjfdDiKuC/ynKVQPwr3saM78p0fmqpmuNfsr/
/6n7muyQdqr/SCkYcLDcHLA3KZlZDPubXZOCSXWnk1u+K52OWQuLk8DAI1i4mH0V
ujY44SXQ9Bd9UFTtqOcfbuG3BlBHpO4FaVWFswpe2V5TBiU3Gkih+f6kzDUeZlzh
4rRANcWfNhyU5Bfg6X+3Derbb2Rp0ZmsXiFFHLqjrDJIv+yloX+yUsa6Ig69MsBN
yO1xnteOlyPy0SegARlMExjVFhX7ur98w9Nn3qy5oVeDvXXt/HJVWFagjUYZU0uu
IRHtZtJjZXxU+usQVO4luKuw689JfB6iOQiEcdbzXBYuYD/mRUMG0YQKFLBr0r5F
YP7mXm8V48ZzAl4GWBwibHV1hr2WeYlXxiDr/j+XGPtllZmSpl64nbsEBeRtGlKq
kxohJHy2DrnGKCM4pWSt3MgYuLMYz8KpkbXcIPBeCaF+hy+P6ZHutGgavbLDFmRb
R6vS6cE6jwSPtoGX8Wb7pIIURNIIJI31QopEQkA1pnMvcfS7qwVLcy4+9gs9HZ/T
uihlMPfSxjVPDJFw72uIz9675yn5CeWBFSI7DLGwAgBYug2GYNQywT4Tw3c7OC2S
VuCy21PJ75E3o5QwX8To9gb8SooU3M64ayx4RV6LD6tEQxWzgi6fmjXC7hpC0ypH
a3RJ+or9RGR/Pe6IX6AH7Ugu3tUJh0gSKumLMl5ZwnogV+3mxP/VBDV1UoMm3Cbz
PmPfH+E6m0x9kiB1TbIuHiLJ7ZsSa/+qiQ/OE6SKAAvWTfNSPx0oPf9Uh9qpQ1aY
VXf0KI1NyG+hsgcgh551RXHHCMwW/zCju3qxWs0d1Eib90DysMIE7GRyXL8TFFz0
eEoJbdjPmbxwa+ZaBXf5jl2cAYY3nzhAJtnF+dJq2h6x4UZ67Zhir7g5QpEBwcB+
6pZSsGJu55HYxS+PeqXhLMjYRAaCFwnvz/AdNXinAB60YkHm1sGJmlu3nGbYwcK4
Mn/W6mUsMXQeu/hp4Cgndtje1SBFDpaxaipyd7dGdhWjtpJMTBx13VW7PPVBW5vz
uHy3GLwsqSxlr+/HjqaFW05vxo691yPWMlGl8YJQE1kpSqmUk/0dfuQLeDpFAH+q
dUF3BrAhquG4F5oRfTR/vhoc3YPwmcdOSv9jsxEoe1qfXvize6f8l9URKZJtjy0F
n9mn7vX4B24xYLRHGfPiP3UQLh/4FY6sI/rKH4rurAwDVoeawA2UXpdnDD7U9rzl
D25201fPL3+ZebWKUiFcXWFPjSrDORS1U8PXVW6jhFJu++inMCNLkxKMvCfEtQhL
isH/XyFctYiOaiI6Pliq8mpu/u6RGx1Af3z/+jJcoe9t77vf5KROQousVZ3mIrAh
HuGKN6MkFJKEiwsIspEr0IV3MvNfxkAHp/jLCHAl8ZahDnGx69DGVmC8+BrqoI/t
obOg9rat+FdOrTjzN8QN4AQIWFHEED/f5mKRHwHQ0x6PIHqeJ0I3RP9/9Jgod8Nw
m5O1iZOkcbx+DZe4VsmfNAN51U5pbEoqdmhDko/dQMAwGBjW027si0jmOOPwzhyz
pZMjooA8760jHS85Y0QIC8uN0mYuOhcT204UrjvM9ZIC1iI/AaztExLmuZR/bNWp
CUomKJznFc7MeTvJARmvxdS6KM56i4XG4zYN42unmqfSSPVNQlwao9y4AC9JkW/j
nX6KdKv8yX13Mk55MuiDLQQCgYyQuJk1+svge9MhxY938FfBi8SsRkEQxHg15aEz
VNY6crWubYjG0DMCVmWkF/TL6U78xvdUjU2PQ9Cz6pT83L8aohTB1i2xaQ1yrVWo
246i09UjdsXFIH1GKhjjERDBeMg1JZ3ZmTTClyglESmJUbN/Gj99ZS6yWMGV7Rrr
zTcJKA+olmP+b+wQO5IOh1LNkaMfdGhgF310vtvdcVrucEGny16TKIOgg90pPi9U
6FZ0oHfdWI681xaHpaGCnoaxv7JK/bO446+hnOV9tKi+niBvnR46LlH8cqTqD/+8
SbpDgcYNDRoVQTi14g6n6UH1qcLNfc9hJQ93Rtse64/h8SxCprDG+aI6K9BDq/LU
akt75FNswk11Skyb45aWXMD3NU4zzRXumnnbDlEqx8hjyGSmbIxKMXMoRLy9hWV4
V60LRoBcnBmS9t52CQb5lzXPb53W6lmbwqb6kG3HKwQyRCMdyy/0NSyNqQAwXwic
CfgpWpsHKwzctHXxjaybIhEdnF3pNAWDcS9bhvOVjnjiURBKdT7RhF80nIneirqI
iyqTMURWcpmKNy0QeIHvZrYFCJcS5TaAGh1fDibPkPKOLKXdOrGI0b+66lhqDPd9
TtqOebht6i+3oQhLJrL/HrBnUUBfq3DfXW1AGAXIvN0ZQu+lMMA4hmdDFYmaYAIi
nR4YWpFKrfRiCOnZj2XRKruVJsoVeGqrFcwMRXv1+1/yHPDRnRK6xJFDfGnqYROh
NwV5lHbzJi8BMSkaEn1GeeEdOsi/67mhxGyOhr6wucjC9FXAtsxAGKO56r6NJe1y
xnuj0lg68Un7yxBgfa0D97qGCaMl6iSY0lRKe1MHOEHmuENw8JC3NAwN6SoC9cOK
Xbk9i6K2nJvh4NQW5W9Rht2WknoXLFxeoAZvMEK46ii2w9NTqHvGet8c+eaXD3He
4Ocw3f7MxnHSlNZ/u1tJfbPkxvzm1nW4Y7/PnlW0luapHCneBqCiUnJf10/D8qaj
zXfTLhoGdVOGv8UfevGw7w+oIPN7YezsyltEPwOUWKEOGWx1FSXE7aySgUNVlS+G
5+nF39RWP2j4QX090rQQEmkcrI9tDGKWu9st9pvJYQ11Cxf9FCOF5u3jr/KTTHvT
vyzuuA8d575JgECqwmHKgCORMHGNd4WcaBT2lXCtSNLp+30KB+EBvkDO8gtkBEby
FsDa+Hy/IhXmHSypYULnj8Fh4CgpFQqTPhUxaSPSdG999VeyRihLxC5ci+0UZsTa
wOQlLNNoyNHQODFNol0DwOYTq3v5crpA8wC6M4aZsM2wNuOqhQHW3QYsczq0FVEM
N/XtWtCgZ/u2F8LxHzJxHLyF2NBXApXGX1hRdQ239G9iE3ATIpm/dXY1G6YPHGpr
5nRci5QGwVpruvbgANAjz3oqe4Cfr6b4dCC0UjFGCNjvCDv3o0+jGYz+AMnoPjmY
d87XCdOI7iNHJDpYyNhkqlk7peAaEWUNMqASJEwGUIFvldJW911O/u5l0+QR/GZY
WErFopbdtO9pusVx/d5R2gIzHHMKdbDVyzIjPR+GW9L6AD07wuWOd4y03mQn+Mcz
wj8xp+/p2fji2T6OIlMCC16zNUJUwIOiSis+iywUoP8IQuhijvsqw7ToK/oAf+iE
iuprrZEkGzoQpxmACiLSdJv0gV21uFGaUFUi4niWL9awsPaRBi6CeUaMCDLEndGN
xc6WF8nrAvcabhZdjJoF3Oj462SqeT+A+LzeIC3qdLA2lNgFIgJC+fpbQVB7cWQ5
/nj7kkTSH6vDfKGlifqrpzYmIfaysDDM5t2lkz2d6uReSQpT0YxzhHgq8/Y6BRgo
oieXTo01+VAlF6XwkUt8f16D+b5MEirk7a1t79ubNH7PdLttMxVtZvPa9p1q8Mhu
vc/BtK4jzf7KrEnsrdbA5tGtQdrmK57mmk5joMp6CWybtLBwLHpUFdlNYaWuvPFK
4h1/vS0KpyncCvnecyNEgvpYPyS6fIWXd5ki9M5Xj3pTnY14w1CgfU/Dq/lnHrBd
pvVeCR7hljU91VVtk/YgvPGqT7iTlag9ozhdQAESvI4DAmjrk1nkkUtsK3+Ksd/v
h6fBKqdYxIGlmiK2Pgvb0OLLKvArqpDW2+UZwzJGKVJBYOvFDS6fsyzaidsF7bJ7
tMGNVBAprsUJ28fb8Ujl9aHs2UQJZOvgcBFiwVrtw7FNrE4iMjR9uvJpfi4/WSSt
j1UTysyLDiDtROYmptdlUzsQ2w3315GKhiapxiBCJ2sjfydg6ldBsMibMlEkpaaU
gRN4G4F4F8jxvkPTTFQvuW7DDYq5wPWtnAyK/JohYPnvIl1iRSLEfZ3fZdctdT0h
GAX56eEkqpS9SJ9f/VI/P8rpa4PBEXF2mUzQMNlsSK3urGs+7/Ckz/+HrZxSSQpO
LhUAhDUEL/7W14hP6yaKH8Bip+GzKSiWOVmDf1ijaIaT4XHCSuxfH3YTVZ0W3/5g
ZIkKoHv2QOrsZZRTNp3niYJKPj5F8oLNKFS7f4swN3n4HLENd4wBgJiixgIVWOTP
V0vgoDI79vc30rJmvfUOmlbgPnHPZfNQtvwkZmThdqH62tQ73MW1yV/uhAGR3Tkw
yACooMJ0FbrauSNnAwnFxArsJ/M1xrDi2UH0/fki8WETG7zoGxyRmRes40YHe/wc
VHuAM1Lpx4oqwHwtvqemOGiVHplfks5W3+bUrfOOR6U3izmdDnCerWM2thJk5u65
GXJuxwdjYcYkX9pvZtF9dSeIIk5S/d9OY3J4edoVH4t30KgQu8l0iz8GammZeUo3
nW1I03da+gpdi2by1WUmcn/nEXaS1hHaUtINxzA64O2nesiibvYxclLn2tSFpzte
S0hMCJj0ie04eqdk3McmoUj9HxaLgM9UpVA+rOqJJq9Q3FBbV/Oo0UgNPj1Uw29d
t2yMZBsfpo//P1DctHMNXAnymoZwk/OnhzCJGcpAOlxGOWUxiPXvU/NbKc/bv7Mf
m2AlUwLjxQAVHJv2Xvrqky1oK+Z/pDgtdYLl74LuDSrl9w4KGtQgygDg8YBo8XS5
DgFuDLgd61GdgY02DF1N3ksjPMKm/4/wxfXAd9tU8dvQvR36mqlDyC/JHU4H5e3A
8Zm/spOwWR2mQBcvsfODku/bJn4Kt6JxuPwFi7N0rLDtbSAm8xnj9oCLXP2sw/b2
O8Thzn28OyFlYfnoIfnzcOMbz8qLCJXRPliiM4DSuV61ue87scYtdmLamg4z/ziv
sU8DvePF+/9X/sXg6lhb4m8mIS97vNIsGLLBEdCTbSpW1Itsx7ptvToJ5Ve+OwyX
Muwy+OIyaNn6ec96gWyfGEZ0zP+ReheBYWZOQeabgxb0+DQNdoDQWQrDBreB1vQK
3GEmWQnHFlxqX4yV7I+0O0EzM76V7Xl0Nx2Y6muDS5ekJlvkEauykqab2Ol4BHUr
i9+hdYPZwS333O/WRHeQIG4sMfu+L3SSQ7jTGdi7TWDW9QWjTPtaTX15HNpFIP9k
09nqYqNYCBEkHxQiWeIgIQ5qq3KFKsNwswL7eDKsi3rKeIwyJb4SRUAyM96Dxb/U
qKNWHDOODZO5VbH96g/K4EUs0NNv43KJU0diN6FE9zbTZbun1aUXBbffjxyTHV5S
fp1+9hEwb2YXZOeyWVMBSxGf8NTYa/VZitjFlFkeX22NpG/W6X/QnmsS8UBZ4UqA
dhEakpLW13ihZMvRnKPjdZ6kkwPTArUoK0gy5xRI14pOYgfZRCaIJqoRg1zZEBF3
IKlh/Oz/KmK1U9/7KKUZ3uoj9YBrinGskZEPvxmkiNDj8MMd0gM7E2zzBzxTifBW
ehvI+c1vjAN6C0dShKhFIZP6+K4R7pDI+24r8GSTfZrc+2pfwEI8x6n37C2up7wp
tiotqJ32hwXhdicG6jZjTb0AyHvybn34gts3ZdVBdsAvSMrfkwX33wa7cNXlVkQ/
PncuggSBeBruWgbP9/g2RFnEatbX6mEpZ9KRIHXTXDLWIMJW9l3j+kSpmTEhR4Z2
uHbQaEJLyPdeU6aPoidf94TSCMUNrDIqO8N8iuBgyUrdFgs7k/Xaqv8bjxZjhTQI
EgvMX7d1KI09AjCCu7nzoGIC7AuiMq43x9RbIv4DshAAdBkXeTTk0A5HHu+H6jBM
xtS7xWlFBlsMUu0X5RBxlSVeb6sbTF/GrvoAaCpNWRfq4WVWxqZ/70IAxF+/qVOJ
AdNnAQY+QMZzdIpc0DQ58CmGa5ljZ/9p1kfujUoK0a2KFqupkLtXysWDEXnrFn1f
LQwTgmzuXb10ZwEBNCWTaaNVJ10Ran8baJFWQtcFtksuzoyZu72kglfOmttxYm/e
NtuVmJd8mkeLg7vMkrjZr6nhnwFZS2cyGY3CLQbb5VZg1icvUV9MjFp+njRc4Vbk
8uo0wJIsTRP6Bbz2PuiNmWKFUYutPwNhZHslfv3IeXMxlbpRI2Z6PB++shDVC2eg
QJsMhifVYa8ghZP8EAHmGz9w5BboseHMjmq2dUPxZFcRLTZRLYJBH7JvQ1kdLDFQ
dbxdEaM11c1QF06pyC0E1pEMKd/pWLmzC6jLFPjIrJQR71CYJLW/md7v+V85jpZ0
nH8VhIyMnEleuBE/zW7AYUjROaLNTTf2PzhdCHdCxtF+amW/m5XXztSFdGp1FeMj
77+wJmvRZat+ALaYDG0022Pb/BjpYk7tKoc4KGBCvKTnL6d3WITmDkaQIHhtfQZi
1ju9mTlX0/QOahmm8aI3KU/+2/aacrPcYN9YpQXZykVzmAKHq3JHVoItr4cJ0+7S
KdpvxwQhQ8CvCHnUGj4+NFiO5Qo5jA+ebXAwG7XZcTNMZwfxaP7rb+SQDrv7IYbt
bqilcTZ+8dQTRjR1+1lNvnCbYx4/C+iu/p/gyAwNnRSxVro7uygAUr1ALBYFDY41
LTnGhQqQMnU7AEo0ddy/C4NKAduGr8ZfOomH6ddYC7FyPsH1ayeB7d36FwZ5pGK+
dZ40qWF/fq14LaJH+BdkM/4YcC1ejx0jrl50v31qp7tDCIx7O8aZlFEVH9tJ56tK
yLJ1CzT8Y7xKzyQxuvGqT0POVUodn3gM6xWpuiDCM9t+CawSbkDKjYVLSzbl/DLn
6Vv1x66dCh0aVMOmiP6vhMDkIOPnYEOKBxY94cbqZSW3EMeqvEe8fLT2WjfWjy+x
QhooXIY3fz7jPI32Hk+Id2wyx27vn+1n/cqnXDVFTu2XU1AQ2u22CbqqpHCOA/cv
Nq0YQjIOXg6SIqrQwH7jecDvcVQektXQXdcil6Yqre2p9BC2EypLstJv+cME9XGX
YabtvNqvTN2g37WNNNei1ic4zgoY5Cu8gCmqXJTpU0KBpvzwQ7rhJd+sPggEaE9C
oiECT858SCGmVVnlK8Fpj2xfpXBtRog00iPSfydCGdLuVImBdgf8LURz7pRfeFwQ
Ilh3Q24ElnJ++rEyL5Obz3ObuddtKDUsr70joX2+CiS9M1xt41atGNUCutr1N9Bv
So7K0nbjddM03ZzvQAA31v2Cje82JWS5uHX3wSUHFQHl4mKINo4FgNVG7yfS8c3+
G4vnOrm5IVEI6juT1bARsAVNpAtOxaULMM1Wi41OChI2mXm7M6A9WpBTadbld65Z
ng/I+qctRDjIMSFPALJ2FRllVvPFrS2AWsRIa8V5i2K+T9ylX3aS0QzyoRdiI9Dr
THVz1f+zs8iBuncxLQ3u1z2iGBgYQ3zTeKqqcQPkjS8sJbWHYfJBNbIXqQsJqiak
ECJ5TRHn61wb0i33ANC/fVFTHA3pCtfApyJa5PX2BN2lgibSCZSEe94KGzpQLXYP
LUHAJW2LsVxLKJZTCXr422ARcJ7aHw8upqgg9Xe03+4u3tDo/zRM0bMr7oskVymX
sjcN6tnMPR+q9KnS7KsFGlYLWvWUzIeKBktahqPsjj3Cae32xCvYYoy5H0uMrUP7
QpEvWNUy4Qpgkj2oSKtzI1UuuKYeRPxMhQJq9RIQGlSxLwRjdo0ub6DOsGBrVj5D
5u4QvBLvKSRnrSVjnbEUXpl62223JzDv8f8FMSBh+ICHjSRRtinE1/A3q9hlYngF
oAGVk+LxevAjL03VRHeolzvSyjfFm2E64kPTjhZLGAkmXUezwaTkNL9AVSipUy3i
Xyn+CtymyCLQrrfyuSJ6dzJo6Xiy8C3UIoL2S+RgDIVLlT4xyXGcriSBSM2plgkJ
YBcabyu71/OAugrW/xfRAdGCpZ8ugDE6eMIw1Ih7RNnw9MrYpIR91/+V9mNCFflM
tOozp6BYt8SqoWZxnJpgVkiV6IqCieFRg8OkTFF0wBILnyQKuQEbxlosYd9xBEqW
xZcsLkHkx8cVad/1sl+/gFHIBkApLS0J14bPXplPDd/zIbnfStUX0aI1VimyLsZv
+e+giXW3nUXrNoCyohXu0bBwDbSZzkP1wo3GShPFygrbk+pkVlN0jslQmcj5RirH
+yuYOXhWZXbQvZ/Lqp8rh/AJOQQj+U9+VQZaoMdvB26xn/HYy9D5TCrHN/ZbIFA0
90Tv1sr3I447KBQHKcJrG95RWjIrZPWMG2tAfA2CMq/+OtY46SWVnKWo1rAe2aM3
oa0wlRljjowIfbvspaloZ+SVZroPf7UD5IMByRVGnxmmOxavzttGYxTCT+oIMlKE
cQkWqoJgiWQa8pUSBUM+Nto787ccGv3/k2CQynQHX+FXNmi7Y7Z4vvFlteV5M96/
B0A0Bcib5eCm28V2wuVymL24fg195WvEQdHWeBI/IXOlBR5jrfeSSuOgAEzyRS38
P+iWXMuKTL+VciwWaE0p+7jKUgADQe3+qwTXP1tZb60f6g/CY8HsAeT3ktrxhZLB
IyRG83j8V4SFwzjkDmJGNjLwyuy7HVAiJt0/susvpGtRR3PKb3x9hIYvSVEAuQ9O
eFtHUb703c92WW8bP7uFLnJfTciK+7hZUekjLb0AZKpS+4cgPNbul32QuheWuTR9
jOJuBeMD1BSUTDJyuuy20T1BhyiQzEKYuD9u1CpI68lHhkuCfBKL2QSlP4u+dGa6
JYIGwU/vKaqe1DSnNLYGMQFZR8gYzAQClKlCcBg3udhSogf7xmFfVJ0lazPTBx3R
6fK71HgSmfawMVJJTrLjmEuxnIEp6b6dIL24mVklU5+ZTCpqQsVIjmBNxPK9zM+O
riZlEToQhM6Z6jX0xNTx7G961kdiBcgyuDzZuP3ik0VEjsO4ZpVHS1LOcxpKdYBt
MJVU2ATESxK+V6p5Lo7zoPp2WPwfgvrGeVS2rCsGpcqwA37ZPs3sNM4NmXyFbAjw
NktOo1gpl1QoAhwuorGulwKeZOPbLYXMWdGG9U5SISjfcjlKBfEgxHutKvpHnCth
QJYy5nNY0BCtAbaN7qUEVjLSekaSXMl+4oTQ2KVjX6FeCfBL8WweDSbU0y2l+GyM
Cqdc2K/WaZBE5qlyjUDPtyuSd7cuQAoC6buoRGE4MrkhwLD2ANVDWqGvhT4V70Hv
zPrgWrnbUOjWfZmXhIuhJSF362PwvUQJe28gxGi8oxjdj0rj0s8P1UEhX9N52zd4
PQXGQhOsOV45fhMY0vt/PvQpSoW0l7bBizOnp9m7Yyb/KrbbOC/o38rFDe3OzbnR
5XMri+nu4Eghszd4xRhZLHBL/Awm2ugT5wEYyeB43b+q7mdndfrA9SLNJg4yk9gM
wcSYVOEDAaHZgHFGZKL5wMF2Q4Nnj67vtfjusD64P7jMB6gwW1BGrizqO5OSaLAg
ZLBueDQW8n6ZjWR9xB1N33rEkSRyBEIj5FlHgt1v5rxV50vE3zlLhHi9IAe4rkFj
dE5kWDa9NknvNTlr/4BkOelNPI0U9501ezeHLrLZkvWNdCN3N6yWISDwwRzaTwrr
sAxc4kQ7qQpXEFeGtTODoRKuemIaJ3LhQYoNEsHc5ZvYSq5G9uw8KShUjn/FwWiV
wTLvnowzK8ChWRY2NHH/6YlVaR+Kja0Ucs/0dS3EvFLj4pBRK3F+JhnXVctykm96
ZCyXdChN1CH1XUv27Yl6/HFRKVPo7d0h3PrGkmT8Nq0yVFURxvebnwJE7bPuKUc6
jw+dfkptFnPUBf0nkb/AAGpWcJLC1rIm8RI4gU/fedm9dM8dhGjkeGsC1WX5VIKK
xUhtDc+TdPEmnO7IeJgxyDjTD5Mrtlj4IUba2gAvp1RcAjSpRd7NeGR60SRrjvue
1Csooy2DF8BRM3TgooPpru3f4SH/Z2oFKysikwz7PnRckxmEsRJRcznnB1BbMWf0
OPJpg31JKSPIE9hn2PG401LwAvYnOAU8eUpU6QG6n2N8S1jeownAs1cqKSLvpjjR
cDVOiq1YVrWVby4sZ3jQVl4AoDj1yiuPUrM3pibqQFRPQymBplYfBrU3SDfrH3Jk
STQgtO8JJA2rtYp2aIHd6/idQrIP3oJ3q/Mk1juBkFjNIFTJOefqlomsMzBehfas
8XNoD+mRVYKp2X94z/lpv54WzRqoGofqMwVwDopupoOWtallOe0DxhN+YK5fGD5s
gxp8xMxy3WGcDalGADzl3KZe0pytWra7+gdH7E99GAfUrZG1kD26k+oVg3Laxg2y
gRRJj48XVOpEbwifFEWZqSYTP6gAN/ZWYzZCF07/b+eOZhv38ePh3741z4KoSmTu
juU7eEkWZNXIsNNgqLCeIPdAkGE2lD85TC2wInxlf3LNvr1GkvPS3Gf70vehBgZh
ENZxdiFhym9b6/LgI9+K7nSwWTYAvPMfS2BWXzMlklujXNZreX8IPUJAQ2+b6LyA
lFbDm5U9sBlQCm988eda5lerE3kNwmMVgOV69LhXIA6rEdd2rGW4TW4DNvCVeaGK
52buyjrkxwdlF3W4z2Mw0a9r/rme2m9G206oMTCfWdPbmObKvv5rRhc8WRg3fNsy
nL2Gf3rTBOsZl55cbQYcsiL1N1ajZ+C2uLeBRfkV6MCNiXwex8oQ/FImIbXrM6B4
goNaYfyBCavUHf7lkCLzPb5l6oxkdI/6psHm5N1JpZyJWNi4awBXw1N7WRsLjb8k
RkAzuWLePPl7WMhPXvxOUNPQb45rqET5BqGdYi0FejVPtlIFkF+u66M2QbAKpFnp
K7w382yu3/K+FZf8I+mBoDySGiuIVRfgNo2BzqDoVehv8il8UV2BLUrIKHljtw3z
Q8J7FqqKuxq94E3YsNoaXXI9nvzVi7KFgOOB4VrGdNt+k9ngRaOrtDPMb/Z7kme9
RPBqsuWzwkXgJ77PpLSjXeyaR199TfU1pLl58iTXMZst+HbJrSk9gdu6V87/0OAK
woQPh/F3zo1qwqWqcz3NwmBW4Mrl8UOI4u4p4K2R/KTBS9/2T1wegGCYZr8+oAoT
5NMaGktoxvYOYdSbIDE8zWz2KKnoPPGY0xqqanM5iK5naDiiaNiEae4lrgwxZBN7
dcqjKx8zbQ1yBYMWMW7iPFUhL5PW0LaTOzOzVtyd2evSAyoJtX6vBC9LMeFAn2ko
tehugE5O+k+5LHvJE9FajGgvT0esSSddSv2tHqG6SQp0nQphjcmws6nL2RgOPz2I
Ni1bMo/nMNvWaH41MgR1sRx1zMeIP9x8/DMqVpWr3e8Q9Xaxod4u93FKgCt3izR2
ags9zXJuQgABkvmUL2dFQwRaRsR8mVtrT/1PplFLHKTOxvOBOfc6B9k0JQIt6wD8
fC47K3Z7GdmqC0NM+o8KblNKV/1mY/fnUjF14A0r2SDexadL4rsTSIM5Htdipzgc
oYn4fPp7/6YC32TpR+0fhCer0QQg2qwaf8hNSkkCW+FlAYIFpelfcVf4Mf9ZouSo
4UHrf0/tfk36OCWgD6zpomPvxbdNBkdqbqkWwf3PvsqZovGQhefgqiJXcZsNpf3R
3RjBwEdo6GGRAWkP5aK7SVT44krzCYjpP9lgJdNF5L0FAHNANbbHX6F6x3V/Fmpt
1weKW9XMpQ9WNAGQykg1nw6MARxNgdviyrFcpdD3dBwx8w9u5ABJJYWx9jQnB9Ln
6lyhGWdA0zqsglhZU5XBuRe/3lSXf/6tCo0jhjbTA8hQZqgBi1ueYGHNYb3V1awo
B/4/jRiw+4XbRfUjnR2cuc4AYJySUr9KEuFtmSxDPFEreq2JSvD99hYxHV1QXybj
/AcwYByZzVCADtteKG5eeE421H+kU1JEyK/EWzt+QnUvi44xwhZUacLgocvlG0VL
efV3EngggeEJ7WE9oXsr9uT6VdrAa+ZZfbXUbGtq5LwrOHgGs+BL/BPaJzx7btfU
y4h4gpJ9huTsR5jZlPQeQVPyGGIt1sC9qm8dXVxU2t/7sKyG/VTJBxFJ2Vr8daem
gsTeNHEg6ZqINum2mlq4WjSwEjVmPRHYr00gVZxzK0B6uvDt9OMVD5iPLogMkGjs
PQzFODEBnk+cJn4BUiWfJKbJovN3KNKYo5Vyox7V2epei/Po1aPSp2Y64NSw40fj
SqCs4ejLs1UJtOpAx9Zgb1b+FYTenUHPdMFMGhchsqw3TVInbhoy9v3Gn8tr2TfE
PjEYx7nyppy44TlvNtTqESvyqCS67bw9uJBR2xiUAP9n0tc+4o6i6DTvsJ1HgnCV
/m7yiuwExhuiUnjlH7vrCJxVlM/qQ9lT4X6NqxATsr6jcPMiG6+IaOc7PzQkqy+h
PGi025ptRm3IT2oKHj9KpzSFxFxFy0blqPFmar4u93kdRU5LNuofDj3RNOj0LDZr
Ji2RV1AqjryO0CnrlTvlc06Hw98vUreiSLemgj44C+MIYfjihu4/a9qtwZ2zXtv1
Gg0tR7nx+RMaPTAQ/TAlAELjpP/q2UwDEDNJQZICjEKh8zf1aC2D0dNE68Pd+h/f
V/3xXT7z5dTZlJ55qgOENgMpf0sJ9mDEG8I6GzvmpBmQ2C3NIttkG75gkiUEZg49
2sWUQWsxdqhlZS2n/p6X7gL0Je1YprkENP1nV1UhrwVRuGlX7PM7hLWwZfq57ybg
YCgXnCobD6quo8a/w0BXkTYyjd9zJdmsEI1dfnfeu5qGmF836+UXtmmGtAIjEQrj
sz3eki5YrXqKA8VlTP4r7grATlHssxUP09kN96OPScr9qzju88dEUmaEQNoU4OjL
zrWEhI1qz7g/pMlfxuiBMayyqRU8EpuzkV3PqvftaniAXhXs9MBv6WvEOCUe9VDq
h2Ao99mCexwl7MXdIzw5I5wvQx4/ZKCaOZhoTTmSwenvCL2008jaxvhPMuN5D3Zm
zQ1X0bQqIV8KtxPLMcqfbkCRGYDpOCC9sn4b5If4xzSe8GtR7uGGV9ah3rD4QT41
4hl2HMeBJuvXmYPmYMFUvsNMrQD1ih5qFBMnkZTI9T3BzLdS5Kun6a9O14QiNM6n
NgYlqinRTB1b3DbZgExicBJ+ksCkEuIzVhBdifGLpzH16JVSFyfsqihlqoN2XvQE
4/znZZwqUP4jy/CrDHxX96woQdUou39Z0UU3WwwPADHr0af2uw/HdII7GZEIsrMZ
iNmNs4pzh0ce/OtCna51QJOIw7MWEfdX8LDmh34vxeX5rN9B2i3ZEcdLo98YHzWE
cy4nwg9HqkrmuZOInkRKgqxdjKsdzmwK8TdcIx83uihR5jMo7qhWApsCeSlZTTK8
lmhdldEtbPdIBqZz7D6ovupWDLYxXZE0rj48IujQ9ytn8mXJmEY4tJAKOUloVRac
DMk3AmVzTCRgdPLmt1Gb/a5xKIt9WLoDNpZsxn4jNq1ruXrGgOhUk9sTTCVMR98D
enthIW8kGjTvHtQKpzcNy97LXiTL2cFmb7z+GAVwlNVZlyCbt+Rc1XMYcGHjAK0J
KGsj5UxdXiD/jSiFrFysX7vFq4qvHp8asTwtZLVLn9UUDUvXtBhmHDmJpASJrwM1
9ggqLsI8Kb1x8+GvJRjY9OROOU2IWxwoT+idAkzTO/V0z5d2k4F++IqJxwWEtfF9
u8jJqyxMXsK3Wk8lNf3foIW4JrLh3b9o/0d6lLi9fYTxQ0CrEF7jdeMOggNHq06y
eTfoWa+yGqFx6Ulp/KvJiup2UasE3Hgv1L2/386vuE9RCScVkUOWOuzacSN6H5nW
JY+/pSiWobStyAkUs4XTm2qb6Jd382qYrPfCnrX1ITf02JO3i3Jya4aGmE4kBFRa
pZqEmHr0hkh5NTMRmC2pGlFX8fvhIe3dDclp8dZKyi/AXufpcwCGVuCiZUCwAJdy
oDzIslyxlG1e3fNkp7ooKttwpaI0tPQe1H+QSqZGzvxtgX/UqRgkZIGdT6Xf+74L
IY74f/WtxUrZF9GpGgnu/bFmM8AsSo7yz4pr5Cs7ZJYZbpelkt8/3Qt8X78xTgDb
qFly8P7p2pWldnxfyHHMsmQMcG1DB6IR7nQSX1gZ7F17C9Z5U8lUW1C26gJqez/7
l7Cujp2QIV10QwrfD8mXGBsSg1EETbrlNEZaURt1s1QuCl7oQ7tWNsa04ie0bC9q
uZr7YHYLYCujiU/cP4ovRN+TKeYczGA35Rt0MEpFxdeU1RujTe02Tqn0atqo/EJE
lErWy/+dVVX8Cci8i5ix4CnO9c1sQNvbDASh5ZOhM8IppefVZQY6IRrEZ/RW69pL
TivlVNWcl/Ku/dSauN3mpEgI4im66gHKY73TuOAIKHPhAgb6a6btUnu3FXHZlUNr
889zDcwC9gtzMB17A7VhLvS4QL8dTLs39I2qz1RwM0GMjUcmeAOXRQ5z9nmUzlx5
4BKBaDGeVG/IrFeEsyzErmylnBiw3/9r6to6P7IvUiwdxmB4GWmNYuVAZ4oXMm9P
ojqGRsgJ8P8aEAEmXLDR5nv//Yqr5nVy2xtD63oYVgG0tO6Tq3zGAAzh8nrJnAmG
di7HT7gQT/6VDtNAuY/sC+8ZOcO4Gm1ur7m49MVaEnPIIltudIe1zZohrBkusSxK
zvK6C8v/Ru8cFUDSl25Zt/gUhFU+UmoKnPoQQmL76aFRpkXcfBvSDwXLF8i//44d
5OzBxTzQlDUT9VrymvXgzubKbPJZLfEEL1scQwt6UXbKpR2Rjbxt67slrOz+vu5n
RzCNPK0zSySE1KYL6jUWmIn67Q/hl7x9bIqnkMCnLYA1pr+ThcW/6i3nCcc3NXfd
8Z9o4NwxXwLDVijyG3JQKMVUG1JCzCeqh+eVUkpeYuLkyHjKDGeKRawKykaYa2IO
zC6BO4yIzH1hP9da7hlQ7oIKp8ZCzCSa2c3VU0El6fKWEKm5m5Aemc083BABiRvv
OdaM76Dgx3I8pcQoCRl584q0dwf/mXCLC6cbq03b87xehJs2SUdbp7NDDKyD8jcv
GAhpv3QhVlU8OLRezU0OjMtVCHyhu2jIIa5xrCOULq0kiDfzxJ88AWZj3dyceQ3I
+CqWP3Q7ZC7FyveeLiYKKjXMfHSP+YF2KNT0JtewruUH/AWPUQsbiYXxENSXkeeb
ARkt9xyTMhSCL1roxW9n8W5r+ASkOixsyUhISKcrtOw=
`protect END_PROTECTED
