`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YkCF/Q2To7BvbCDXlyrjpGA6uZjwAi3jTwrn5GBmBxtI4M3ArBhUtF8r9OuRYvkw
Rj3/ztrI7FzrJRLm/UZV53MdaAFacrGu8MxcV6S/TJ3Xgic0hzvei5gGzsRJjhMq
a12DqG7pt5f0JAvZ7hDEBV3zDxEggWSc6XNzw0+G+XRWLHHvYmAKc3wrm8CDsZE9
/VZws+VlUZTfte0h18RaBu10ptgjur24WGYMtTzv5M6gU0B6/ztFTGc97hlUXk0q
r/OcaXfqUeVfo9MEjHbD+JIf7mW5ZmyWxpa02Ogqix4ZiJidQ+vcfAPSIYVlCMmB
YH8+KFl1nFdsJIOCetdbVv5QD2H4nOWuujeG1IR70ELskL8ZJGqA3Tf9bZkzTDs1
Ct05bvZ1kxNYXU9zPpSZTiatoESZcoveJGlUNXx9hUY=
`protect END_PROTECTED
