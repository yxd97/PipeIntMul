`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbZ9tKr83LRojdG9aFF8yd2ttE6yZPtw+NmfvTu59cGU1tV41mNyVFk1MEQiMGS4
aF2iJxP+TP+CX202wblLZtWZKI3VvAuVyEzXKD+y16ZPtNQmmsv3ryTxrg0GHXxX
DOC7/3S3V3AqGC5KhHhokHPICL3y2gmQrMz1iz0GYhpjILQ4wSC4LQkfpJW0ZLe5
BSn9ceOAXvCS0pkfZLeY3t3EXK7k0Z2DnpEKRcIS+SVqr+6Fu8kmWpI8HXWq9M6Y
NwJ7GplEl54zPIEDJZLhnT0Rxn/4uuH9WQqChxee0SHGpHTz3aOiQ/kxmxmh4QkW
PN+7w43QIMu8rLTLpRub3XUkRst4U6JaUuANEHfFUXTL1tVHiF4/w3CQ3B8K5K0K
evjkEI2A+0JCibWW4LCgZQ==
`protect END_PROTECTED
