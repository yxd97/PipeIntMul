`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/VD6A8xsnL6CP1ofRZAzgNuV/QPh7/sDJ6WujLvarTX6i89NGtYWOfk1wROi5Lr
qhqJCcDIKEbLzfG09lCUrnmXDEx1O9MzlO8q+2w58PcwWnSUhL1MGpOOvqKq5j80
+Z/5T3ht4RLC/00BUiZOTYfPuT5v87Rq9Vhr2MtuCAqz93k7QywlTwyLTtxwWuJ6
gG1iWQLu+zIuyZPmTGpUUeMZrL36MwMjZXCSfl2XVdVkZZ9+UTK1OWxRHwl6+p1G
5X1GZlaIIp5/FURqrr4uO77kO0B+QAVsCUZdKrR1J1IBF/r+BDIcbzOlob17Zqxy
vvXWFEWKnutPVy0GpiJlRBZl6XTooRwjde0KxXpVy9f+P6QKNn+/jhYfvKzfq8D4
M2iujfozWfYeUR670dedSk17WpPjCQiE8bguz0dmeX/NujjVtSZBpWUoqkK26jGF
VAMmu3eWnhEWv5Tl8DCFK1UKhMcKqZMfiWXrMjmXrLbhh6wUfat1HkdYh2YpOLo5
DT7BhmggLnn0r+blOKuz3xnteNUO5xB+lrs1j0O9VgBqjZZSXAfnpcNqZu+0qcDh
n59Qr1bJb24lOiqflttXniCcFax8sup/o1cknFuERWGgstnWIikXrdCO0HBmLBIN
GtxtwLdgzAh0+8bKeAxjig==
`protect END_PROTECTED
