`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aEMFP6Od6BGDluxU///FTq3SL+iJn3FFWGPapnyPcSs2dpdJK+sKNPHh4tMlJzWs
SiZFubqr4lotAaIyeOz1D9ZsUfZc2E3kATEkSIxrTpOYOvbfj6esigsa7WZ45HMU
g+AkAUbjC/UivabIksdtNyM93e0lkvuMwB5t0vOa5+IOpqFKU9R07UZE3gV6T9Wv
8TQrXSPqf3h7FCtwZylndt53bCJ8M9kC5uaLuUE1XFPTBQjCSsQp3aeIBHWN0XDF
1vTRcS622jPv9ri2encCinPxG5MYJ0GgRmCjqdNG6/g=
`protect END_PROTECTED
