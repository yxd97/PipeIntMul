`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ky+w1mw75XqmVFCI9dJJGKoYf5NkrlweK4rltIdhzsdk28mMfTTN2oYxuF+pDcnw
Q802FStmHRKYd+k3ejq1tYOWtf9GozIwpwET63fSkqibG2sEJLJo2/ZhsWuyoWgi
/AOQ0HT7k0cJgPYmnmGK/NjVTSI9fVVBQvi0wbQJw3EnphZVm12WMb/GqM9GT+bb
YlY5tT9CQ4aApzFXiu8vd0WFntINN4u4Y0knIDth5xufVqfTpHdyzFiXbIGpSxII
6twZoVJECCu0BEZkAmryZSwxcqpcLmSqGU9uVXGtU5qOD/AkSSeOetUKpDd34WZX
XKJFupYcJa8FFcec/WHhkMOVy1drSdE5ybmSepYHJZ0E0j+cWH/laaHEgcu3j48/
Cx5SrCLJ7h5XuxNQ3Rq5Ugro8/J/9Gre4VbDtbcggMtfZft2R0gTbPb6jaD4+Bb0
Wb4WWnrRhTkG2TRqo65N2HKfaApfmPS5ITAnQOnntjEt8S66qruWiZQZPO+mg4Rs
JzFZt90r5DWSqVHO9+ZdON21GnVMNidXm0RbgHaioDe3qt68yggXw65qLuwDt2Go
97EC2Vpai71bmpbiS/fENPvZ3+GXEJ7AK4SpEF8QEXp1TWUeY2odu/Wo7PPFajYl
q2x1yO9F38Z2onx9zZg7EFxAW4nZLVKuI5UIAUiA8SoYJw1PRAZeoRJM0+AYkPKZ
lnAg9A4+RSKhgJJSQuvEjd64FUropnCx7+9Y6fspyYWXp5M2uywD3mnTnsAQJ5RE
8g4c2esrVwwq9Rr4KUwj9R4+jywha9NwfWTq58mC+m4/0eoL3iglJcH89nvhypOt
Ftd2ZqcoCEe7RqU3A7fQxUYpLoEzMV9NDh7kihmR+5SKxLAxqms6QW+ioag8tvMi
J080rJ5looNCR1WIcJ02OEN9Va4CL3ORbKxdEe2ZjuPwXd47Xv+AvnlenEIb8XnI
/0BklGWlwf4JINHIs9MzJcubU3fkK8awc1eQBnSY/jS/93aen6XAIUJJv+z0nD/4
paU9cZsKJ+n6kL3xQ/H0eycwaaP/gPKwXnppbaBL+Nhpb32Pp2HZt7D0Xc1p2yk7
m86b1qchWufVkPOiA0Qv7m+8c8bGHR/4LdUEV3FAzHRY7Jq/utXCCeCz4+seL0jF
v18Vi8C5IM/HqgypXbycvabN6YwA24fvPIaMfdu0cGlUlUqYMRHKSSqN24RyBdCG
sEMW+90LVKXG6U3R9qWKC1cp0hP0Yllff3w1TDuW08mr4uPN441vJKXOhuJzoBu5
vrk6oynDkND+Os5m7r7fljLY9OgR6G8t7fuORhsyyxXtSuXmCXyPijv/ixD8kUSZ
OMNNXlBdJlKpB7uWM2rxjkKWShQmNxTFCMrcYZPHJLfsIlZgf5NOkt0vmTIxZCtS
A2pxnHg1bPAxXHsQFIdk8ztzf+T1YzbnN5XhruSc5wijTJ0LHPHMBlLW/Olavqh+
7bVlK8nG6lVxTBMlJnwgbWs7D2jQBlzlo6OF4eOFMFujlpYFiL2eF2Vg0qYynZub
amv1M5XBQgTPVV96SXduvCa3yyP/tLinPVxk/iufktS23aciKa3m/xQt5qF4WQJA
RgAlM+TI9zC9+6RYMvm718Nen5ZWSx8/LLK4TdUBTA/kI+0m617F/BAJgsNJcPKx
w3g0oOhZoEO1I+biMbYZ8sT+E7mYFM4+HN9iBvXkU4mk4sDRgJEuFm6waYCkLG3V
IA2Q5Y6Ef/9wPhj3sLt9p5hpHS3Go81PLqt34T7dPPYqaGbx5YDp+t4hikBtHry9
LSYP75VYMQDCldMSlY1xuHF9NBjxIWAoRm9rv4L6mWllAobwKXg7Rvtydl4zbkyK
aUI1AGBppFDX42UahFKpZ7l4bwhr0hvEO2/4fbaDCcKwqyCi1fSSXEguJBSV2FNF
2D0M8QaAnhyooH5FzlQvP2UQpeigOR1o3AZMmxwjQP8uP1s0pku9OqCKB9UVZhON
634op7XGF1eW13sLvRpIwgm3M76QUr0vQSKfpgbt3t6lcPGKYLT9W2p3fA19HCJa
aZSZJMTLfbU21aQUF3RD6AtA7PdNUOdOdcRwZtSHbXl89ROCpd3+EE3dXsN2i+Bw
BBZVA0ubAhanDaQjXlFg5K8hp+w1Z7ZuM00ajyKwc3PSpWunoNT+A7DQIyQbMP16
jH9t3v6bPUgDvcZzLIkKvphkUk703yNuqwy9cl5iL5dR3dIEoBw1/AVpvJR28c0O
DsQ+jmoUYR/3/CW518lBz7Ioa6R6txtY1hMcHCLTXf4GH3mPlmQIbq9zlziFAHp5
Eg37M8JeyzTuPrkSZbobtVE2TjS1ka93DuYL2umPTTqkPELCcDTMbifjpEPfTiYe
6muommKpIoT8b0SP0x3hgz+YJBPn4INtXolauBd0VBgE+y+ptNvDxBA4MFvDGRV6
GRxLKeWLIIT59kq78pbQow407gQuFLMaGcm64eMwaK6BcUPGLjvechhDNk3tdHfj
CQrXMxUHZzXHOdbLJWjSTNEQ1gVoGjLZqEZSqeYhhClbRh/91qRuvf3NCMRoExjP
hm2ZNMIT2eyaPKmQvb6I1Aqxt8pR0bImGvOwnh1awadA5pToi3J3fPBFIQroNKIX
TZ5MOn2bhUZF8U+8sRBdYUU2ueW1PmIqh8P7mnlblnwB29jYoMYfnKlkbSqWh7rl
2BCJbbLQ75425VD5/uECcrvXXoDcEvPbzdTSoU2ZQKFJnDO04sFQ7MrmYBkugzaI
2wFk28apJiy/s7f3I52FoPPLQ3nxEc6ZxR0Y959SD/QA38YDjXYDjB/FAGe8BiN+
v/OJychPYKo3z87pQ/1iS7Fl5SqHH9HPwkoeOIwGNMLF/+/hCa+qrAdz34DUk5/b
nCiEgj6cOFP5e57rH/Qw09GSnES/1+1DHFsGfGYkZiloHtaKfdunaTsWoIQe5ba/
jM/RsDMiX+ye2K39WUqQaZYHBdLBSdoDL3un9x5sKnYHDYhMHoJq41XPrG23/vfE
lh7+urnjdramHayyfrdkGchYRWkqVLCDuZjtDOocK/unOdIF/vcLhGmh16wKT2kQ
akcvsOMGXbthiyZ7uHs1PQ+oM5vDsa0uW6epNdgVpmjenwjRMphJePzPK8n+t1en
7XHU/z/1H+ir1UZNva96aqfKkNwAUJfPty6SB/JX75Q913L+5OYKiTxr+3u2BKaG
x3nbutLsnOQf5kCv+aY3qS9v+CQFe3fPjoeQz3SBwVfQtGQzm3waMpNd2httT+RW
uls5ZChDJ+LFuOtjeP4sC1ZXh5qq3qd4tZnf7PkmcWglkgMsBYVDL0zaMEsLp8l7
dsdIkVCt8uHlVjBiUV/FGR5VLPGiM8D3qDSSg1NxrQXxotlDpy1U4G8p2pc/4o9k
wDsizqrvDToEbsFxPyVz7mJoS35VqzVudj1k0GBSNbnttihMC2nZJw+fPh3pejtw
XBOjIG9KZDjgqxPnpj2AG4phapOtBGB2YXDg1pNV/u6pmllH1C90jwVh69t0rcJB
bDSilfi3eU9Lt6A37w787YQuTpGFAhi6CYMbad0THqUsp7vVgZ5HEeHUXq8jMdMZ
MHFx227ARhfB13uz8wAKlkqknEYVn7+vR6cKmo4k2K/YOmGfCgMKeNi/BNHo9tru
24qgwEtFDksWDPAfQ9CdsSkGUp0XEodnfP6MyTDzarbd4imON+ZXMt4jehfGv+/0
IeErl1mpUqU1x63p7xujotmj6evtIAOK1ei5sQz12wkgAmMziivu/fhIrVuJYF2t
a5icDbI6Le/S476NQ91SR0GWshxKVtNGpmita9nRmsTK0vbyzUxltFadg9JiUnW7
vD4kvjBt/f1otTq8+lk/DR4fTSX7vLcgtWkX9Bukf+Q=
`protect END_PROTECTED
