`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOEFJTmS77X4F+JNkmtYxNZi2uCC5TkVmYXg1K/l6BVczIezYYFDAgT6Lyee5yZW
Y80SvxaKgQwwHj9ovaKWoaY2LejrobP8q0KtXGPrarikQBHZHt1PzEGWHrhwNRC+
fJNiXByrlbTNLxDY4BSviotGTJTYoWpT4KrKPOpz4mwhPKT8JbEwGSuFrMiGYjN3
3ORtnpz/w0/wyjQF+g3URF97vS03ABW88+4pLTZOlw3QV+O7TsYJm0MOeFuzelEi
TANtE4r6ElbBRzKCBzWZi7JNmwdCrsznFcOaSYjpLFh4d774CGhLNI+wMUkJkuHI
UYLQ21q2INChGcRUHPpI3a62qObkkEXlFc7XdovCWKWhuZRsEy6hgKcstbLSbHlB
9tW7c9mI/IF4/28N3krYZl5uulL+vJ62lRQbt/ZoiMQjDYBck98h7616znVpKoNp
ywS/2aOCcUeZ+prT2NUYbroasdYR4zGqeRPTy+e8aR2b+QE8/ZjkbbzqtXxGc6wJ
b7vb1QZAlus7yxm8egf1hSySteRg5Nv1ZEcyu1QuOEKifG3OiPKetLanABmKFh60
sDG0A9EwHRU4uwirY1v1K/l/EAAIuG/h5n9RrBvz91fcxoqeCzzCN8ziXv4wGHZd
WEFRqXXWwjY3viutsj7SnA==
`protect END_PROTECTED
