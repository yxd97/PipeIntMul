`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHROyR8GKzsbhbCo/wGXkonRz/WKksJeKqty4tD8ryRvg3xmxIn4r1krP7l1OIyr
ODlbehADflmo7gJCDlQgfuoh3jjmeBJEOm94QkdVmLgfDETeKdjF/RsWVUGqMYVb
15OV1kG5RoydJQb7K6OfGjC/21k7NxsfKfJkVCYHYb9Lfa7xyOYVAbcuvdPftdNq
LJr7+a2U91Uld8ZHw1espXvVB3o8mfh2jMnPzx8f1IKfly1YmJnXb+lvqSBsZaoG
GfNJ27qZwaZWG4NXg3IEzpZQphDQlyPcxaZxNOxJylk=
`protect END_PROTECTED
