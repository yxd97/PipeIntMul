`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+480Pz34uKQh6xAnOeAup+F8+whIQIwG9iuLmv4T4wDkv7esgjTZR08mslX6h6ha
x5YKj7QVZGLytkhy/I0lJ6lY8XJ2XXzpynlQDTH0i9iWxs9u1yV7q9bVsQTeBtf/
EqFZbasSxffr/bluZYij0VaLiVSgznPSV7hNy/Zyrar7GL1WhD5Yv9T/WXisvwfj
gr8/3m5hXzxt918dieWKfmVh1CQ+jzsN2/Se1MQXDIjCZDm7oU5J9o896vL9u7Gv
U4iToPVUFSvd9p0yj15Tew==
`protect END_PROTECTED
