`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X6JItLlmOKilHAoq/YjuvcPvkclJ7zt0d9Whl36Aay69KIF4i5zNmixIlh5M4U73
hakrDrZ9IImE5lJmhT59/V3E3AVpfd7JNpIj2ZaP3dt2N8oKuPGuWoezmAX5vXGP
N1KXppsEEvBX4FvNrYtEYWUHTSJ1ZAUNyauJ39lF092U88EfkntjNb9JfQR4Rih+
GZwgpgKOB9wrncBZaxSwVtMKp7rI+KPjlCfWoK8/RFXRZjPAakQ7jTm2iMeE5+qB
w0g1lGzDbQU8vcsp6P6s+u+pIB55GGR0U3FpC3xD7yleu5PisAZnzCi3CWdeMul1
k/SUrPfkpoK3qpeYeatIa2rLD4WqsRWliQG4VZrLhGywR+PpP1Js8NWQs1CH+s6d
FhX9qOAVQltPswsxJQtK2bJRzL9DMw50pNjOuYeemOP++yg0WGY+3OyVkt1tFnET
BYY457vH10IIEkwoM5CUHt99IR3GjBOpuN2bRFK2JmE57OErgs7NbDqytXW2fDUW
OIpE9UPJ6neInhIjGzrJN+R5i0DslrS5jXzonpZjUVXxQMk+7xxD2wnNqcXlqWZH
`protect END_PROTECTED
