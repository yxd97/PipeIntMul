`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GrXMZxLOpoLfUT4iJwCNx+qML+NRJSSb83lS6yJb4zwVSkgb5TvP9a5ipXRAA5Rd
p/eL+VYu4zH/jeOVWSL1Yb659ocHR5108j4RbzAiadTWEfG/7F85BI4no3hG8l/D
eONlrfhsqVgkFLJimeWkRkDgUg5AzCdx+6xH4WIMAtLf7NgR2Cs7VNREC4+Wq9We
KTA6q5SEvRAUUcJJczNXbzPHtx27GgVK2DQVkF8tPK82M94sEDdIuZ7DVf6OIQae
rRG4bRzNaDfsnLV0DlDRkYed5RwpKn98eociQ6/oLjgAQ6B8CTHx0uEnnCiuFTlr
oGXZRXtUoR27g5mHwHCWJh/YtMLZrUhYjlxsgY/5o49955wqGkGPJl7uEbwYpoWC
VGK990SEmHlznBreitscCmOLVuxJErzQ06SepTReSuz6KcdBAq5Ud39e1eCU7Bjv
XixwEwYri7jEMUt23tQ/46I5pxXj2Mr+4hNgFu/cd1n7HlCegJF2o72f36hPOOQi
bv9YAQ1NIi1mpXlIaId9Gd62bfypxTE0DaC7miSiWxBl0UCGdqF7A18q2AFQQfGv
Hyg2KxoSrjZRTK10qiY3Of+bO6OJCI6y8y/nEOdwuIF8rTmO0itJTFbT3YDk95y2
foGVKBv15Sk3SL+il2TSY6ML51xAEm72/b4nNgNkBs4=
`protect END_PROTECTED
