`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1yoinSoB4cd4vAzvsIoqVzDehvlfgvzjsf2AMZQ7NFvQJa63PL2Eoaz2RNscDmEi
CMbTz/+eS4IGJ9AvD45ejF6CllTvgTPKjIugMk3QW1Nd1f8Mf6Y5FD0rg91czw0N
jCfoOmbKWQortUk5s1eGRFAYxrcl2kuQo9kh2TLm1TTrYKALo8+hVIqbtWWRafzL
nbZ6z+wYEtaaASSyJ9J8qDvmJ2eSI42A9D3wnHstrZYO0cdvNYZMdsVMszNeJNEO
bL8aqqSBCfUBcdkdyyBCo32jxiSUPswtZK5F+ss2c/EcGTTtWKy+wZ1KHGMq5s9j
7isz585gQ/+YB1Ul1t1U+zXY1A4/VfVHfXNLcx3ZO2zhaWyCHx96coVFpF1iYOZo
kKI0frRwFKORV/VY/Dzv0AyZ/myzpvmyuCSVHBN+xF11gCc7o/6/T0x7SO0QPEaf
0DcDGWXli+w4elXWx8qS2S3PxelI9gq33HVxcol+L2JFPimm8zKlmT5M8OnZaNMi
AAzVH1dN2H2WWCX8PMbkZX6gjjm9PIWmYIliH/D6T51LqoNGIlXsuk5IMYOmF7dE
pjFZMP/kI5YeyRZ776w5E+2UIupYoNEWSUt78Gkw6FAUmlCyibX2zcW6hbTQ8JWS
lFUadOjXu1PrJusFTNOm79Uj2EyRugWv2MxlSHscyZd+REyq2eiF3M8jvcu1Rk1k
jrXIqWi+3wWOiRCD1zYQEvujKPOVeF9YKK58UnJvz4qIsd1WWAdmBVgMSdZLqbyW
jkXPQy3L8cCymtooKBLOUBAGBIv4+5x8sZVjRhjMSfaJcaF/y1NSCdmq39JG7kBG
7j0ldbaCDp/4F3DSYz5nNL/73iDv3iz+T+avkficgCizb73wz5KZMvQulVQnBUjX
TNEesYFe25Yh69FN3/FOLkrHys+1x7Cco93RAx1ud6C4ZtKCyLT5NcFFLLTMOXRZ
8JxejG6hNbj49JOvHuJsj3INJbW6cm6whjF3jf00tOQj/NaveSbeiFrsgXX+3l3q
Vf0bferK7HV1vu3N4kS/haTgHlzWuYUTQY9WCEmzb0+fB3iIclbQlgYUwV1KYvPM
Qbk0+CC0o+xE+OoGemYLS1gjcInWPKW0AQE0hjyn/0kilo2ctZpn/XRl0ueHBynj
Fp4vC8pTPLPPiNXf5GoL+rcleJrsyCV82zevEORQFN5RAFbGXfR3g0H1cDFQQ0Vh
E8uTjhWuTM6fI3zUdWQpq6W4AMlwBq4xJEDH0DxDUHgKZJyjUqC8oJgQzJ3bFcET
Nt2U2x9ll13ZCjAN//+n+/j91QNUEREBIFBmr0sITxJLxkDlwFHZu4Pn5YeIlFlC
ZfL4qgUL3Duk9TAdmoFoLXw3Y3n+N4LOlRuXuh+MXED1Blp1lq1ZhxqzzHDna2uA
xzgDp/UVOPaN54ftWrFDGynOJvoxTJhca+Y7zpSkG3z/Ip4u1B7QM/i2H6H34Bj8
AkcwOLlDBKnw19ScQmfABFTPdARQcDwYesI/40ffilIhtXORZXtB04aYkODgKBxD
PcyFYPiAygzuvKZzeAMQBuX/0s5mBmRDmt1y6eqIlbRhv13WCzhm3d45LcDLaLYz
LTsNOca5TP7dzWq0jBd4lvkFDqlF2+fI5b9YHC2FYzzOmCUq/O9bWlstHIKskRtZ
1zWRwcangmpfEB9o154/o8gaxjVGiELggLLmE4aegnWxxjZ2oQpx9VOVrpW4WPSX
wwIQZGousQTTGx22BrLsG1+adH1kVdweoj+SYkqngvPpc0LAThpuOQ/hY6GSLJrf
a0oWKKzO7w4hvtbreJo1NgH1DYA1Ncm/X1x9Tl5FkhyWQLU/jAEM/31MYQno4OVa
XRWvmQCGKUeEkt3GVFljvYQE5RWpvrRkFQbDC13/F1zgMfzPJWGocM7iNGZcEXm1
jp5XatcDzqeXhq/tYHq0r237HJaaPwnAG4g251MklTjVvU9U11eTKCp6y2p/8f8z
+BIW/sMgDHnF4642b4ML/V600wSofuylYpjCzICpYI+X1YqNiYdawg8/xCp5Ky8E
ykSOz1mY3hhfvpsRkZSdvZ6eJyuePHIT5dEMVOkAW/RMWHnI/TSOCLrGLkp/CS1K
UlMrUbByfwXRFGdynRsogHo8lOIQ3/HvTxfRquaYqLhmcjd66hw04WocYEo+qtl9
ExPHRaxckp+I7Za7+DMC1CtBz0/BxipF7ZDi0yTPluGacr0SCaGvY8gCzIUnPEO1
roi7qaVA/apgiy2sTvuyID2LZZYUT0L1LwiIg2ACUGi9P1O+jQ6a6zaO5IX7mbqY
mkzcDfhhA+K5XRTGCtjeaedNKKnW/03UYdTVXn4vv2e+k9zd0CsVr0OyWdHbX+PA
dvufc3IpbCQ4NE5Sx9GG96K+TO8PH8pNCNyG7/9CGvq4Y22gu/dtb9nPLLVhsYb1
kA5DSO5fk4ML3I3737OZVpy+dzTXdRE9lonTWXvfT7fspZYGzWG+/XxxTQvGVgDl
z3UeVDKJb93b2KYIfuh+jt+poomuCx09+tm660jsWDiHbhzPU8Qzk9rmMOI11Pdf
Eum6VCLnrQzrv4TL077m4J44SQy/L8/6cVU3MP7jOXePnrhbvVBpS9csS5VgC9vu
+uBBXeMibG0yrv1v0DitV2IlR92rf2OWi3KoJAxUdK8YvPJgzHJd/dq9n5oMd466
E91QWsOZtJ0hvWD8iBHG/8CV/tde5ITJbqaKXgSuCE6gFX0tvI4dmqd+b5b1R5gc
h8cSYFG4VDIkXNclFVTueI0nJ62eWiBZxVfsAzqEe9fRZlCKzOkBar3eo1XqUHKf
vD/K8oaC/PLe0WAQhH2L6ViA4tn11tXR9ShLNsG88CnXbN68Bo6hflrLlNrJa2aK
ai5gIApyROLLHU4JyZYR5dQF+Xqz04BLqoDzToSua18=
`protect END_PROTECTED
