`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JLdUfWi7l6CSFF16ogoY3K1VZvRYN25THXfqZGM8aSE06RRuHXwVVFnL7RsUHPTm
XmnuFYiJnOlYKzJX8bmlgmG0OHtA7yDjhPaVOmQcz8SOpwevTo8NyEpp6QttT6rq
2TOSFVOl2V59gQ006pwZXm7kUX/g4Smc8uTB6iJ94FMBECEdefP/QumyF5Ke2WMy
FEcs3sP5x3hf2BHzuD+mlJmAnak6lKXqWlgnPzXUeBU10EL8eNzj5xsLr0x2JWAd
0kIiumk2Vg+CEnksrYBbNw==
`protect END_PROTECTED
