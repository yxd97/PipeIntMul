`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KR8YPGTh6Rug+ShaNMkufH5Jk4hoNDea6v3xHLqX+X8RMUdKLzwMTVT0QPHkH0dq
SH6fiwvuV65PszZ9uHwg17hCgl96ldl1Rmmvu0fOdflX8EmmYfHxGm4tfu/NFXUG
cil1YRx5oA9QKMoPFm2Bv9JAGntpPZH1frBlUODYGtq8hvehswh+e9XC7GGjO7yT
Z8aloyMkXbZeZRO+Nf9MoHeAaY7APBxiWwqgTk0OkrMn08oIgSA68PP/aSWwjsd8
W9709h0Tnh3MgE3NYjn/f8Gubc90OSKeFKTfCAY6pTHpYi/P+M0LZGXwIDxdQVdw
T2YNVubQDWVXEB7r4kh1xkLs548slo9MrXK3yv6HAr34g1rzueMH+rcky7mtSwZW
PyGHnFqgIVayXHsmILIJi0BipGYLeEF/ZGEj4joDyb0/QosHid79vqdprmS+70yS
MPyzMD4idhcRmQ2mgHpB3rIPT2pOFnw4o/KV6CaDUchObntUxxGPPW3tbph3yAiJ
fUIfFWw3UQtFE4/ZQbxj+wp10WJ+60GJHmVFEDRUIwZuwH7n+lf6btfo0lSVm1F6
KJg3UGtUBIUqoEFe/nUry2Dk+w/3bYx4DxY8Er7rzoX8CbbmBEmPDNaPRPHL/akp
vhyY87hra8TCkjsGgaK+KJiWbhlmw5fNPCYA4Axgf+W9jFs6aYh32b6r+J00vDyR
QHvRjS5vhslLhvXwr4ZoB2XZR9sie025Op3tNow8rYUekQR1N82ivfn2ei0Dm0Bh
otDkSREfVkvk+LwAsckX3JWgfneH+n08hO8vD9c3v1/Q86X5QXtbenYfv6jPHk+s
pKvE8VRW4s6X2J4unFEGhGeP56c0sqoCzO6H1w9dtzFfOhLZ7PUC1iKYSoltFKHl
TABLTGVBcVx2nx6nrya23SIQTAn5J96Elg6mwHECnHQyQYNYqtPmTAHipa9nIl0e
5/mhhw/TVG1g+qmZN8NWbQBHPfJpvENyDB8oopYeel18nE+WDyeG0LbEN26QtmaP
rgBbmeD0W1nUcytOGgIc1sj+IGH3GrKUSE4uGPwwtVupkzfs9oGIu3MRlV9PjTeO
7i8YzYdjtTvdHL+d66om4E01P2JUy115cHcyxRMXPuMwyjXEycBrOoJ+aqOSUmU+
NU33MKq4xLD4uhNYuUDS8JGfj44Afo/i5s2YhDpKvphkZbWf2A9d8tbRRMBsGVm8
AuNgbRuIktvek5kUlbN1AEfcLi3TSXQGuqlu/oYO1byGgcNc5ZHtMl7LSAwMSElp
DkquA1tctug7sqqml3giZxaP8FAjyyCPNuq2eD+OL1j35EtVgzZzCPVmIY1mA2oJ
FvSnW5vJgmn1h4Vncbyq/DbGjVBxv3bNyWoXQk1QtNA6is69y5xXwLrTfYdboLIx
AYnhINtBrn0pMRK5buLwO4Emt3GQ4aFT1Uy1ea/PeTeM5YaA4Z88j//jb/XWgoIb
Mmjh4hxyC7MaUTpr+3BPVTX0M91K8lC/oTg2V9dvg1e9nTBmsL2zREFTJbDY+ujF
MsqEKebkFwObrafyfylNEZ88qeeuLCRdsSvl6gMeIkFstFy5YsNSTjNBntOQ1Y1B
4XR0wFmWC0gYeJxZJUZlSVayFEsAsyO3CslXOVNDy200EUuXNjDVZNURbV4XUeXz
WuW/OKOaZEgfSo+rN3GkMtKuoJvLqZErrWgaUXymdtNCyHADjdwdsqCm+Z5AZgsp
Ej0jmZ09kwXhtS13a74ZP9JknWLVdvcB/JEaqggu8FiNKXhJTnPmQHOFX75htNtr
Re2CEDqCbFEUIrB8q0spNVcTkICjgc65P4RpY5ad2mAjeg9s2jxA1bsP0u1rSgse
/35LU1fXUV+IovSTWaquZa2Ob7+tCCv/Lol7gj/NsWOGchP72WseqHuYE337CnJu
gKsS/yckkiJ4BYaGJ3gwO4SiShXm/jSCt7De+DhbSjfqMb3vInM3hrEHXjEd7pLH
h3ba//uQNrjZj34nCHuv7LlMmzIWuVq2Q2/juKSU86yqHD2XI2nr0v61v7ws4Wlz
BQCkroUgFzDgjWOqkGE3m4bdv+IdaQMyfKT3yBD8BmqJNV+Iif9t1B38nzGInNrp
iJ6qhyOAdqkXXo5bKsWbQPDC6hULbpMTQV1zKCrYhztWkk7KqpLjt9hlDbcOXHZh
WmkM7Rca/r8c8Gxv51PBPEKzyJscXDSMZfoR3eEjn5RiXX21F4ZVD3mz/X8GH9hE
W7FgsQ66gqzNNyoOTYQ845W0LElmDOtsc9aH9/wmg4n3hgIz8WHiAvWeU5MJ61L5
Q2v3yHwB9yrT15Ne3FtgthIF7y8BF6RzsBO6QAUHxzl3L0iaUolLWWLT68U4iL19
7yv2XpUUN/JjRgT/kJtzOG+WBbFRjD4YhmwXtY/D+3CHVjcEuGaE6gq+7LAcKQiZ
IGoqLWhe/TZhGY2MHTBKYkuXEKy6NdCI5Bc9iX05ahyNRftBpnrFufKa0L2FpJv8
V9kwh7zsYQE6w8/m4u4W3tgX1qNWh6amRHG0AE0TwyyHtRW4TKs4jYfm6av7tQYD
lU8UkoaiH1eBac5dFWKx1VczTijgqBQ6+hShDLesJvErc4bkd8iWKy2a4pA7t9AA
PxyC+a84/JScW778HZH9x/hcDMflQCOwfkSzQgaHhpB4hq6LL7lqUtQ32idZXZ1U
Bo87CPycyRAIANtD2QTRGZEL7zcW7P47JPHpw48kcxszzB1T5X7OZ3HqcPPCAgov
JXOZfzeskyHbIWxkOc1vrnJwoNtm83dyW5txdk4Un+8eitIHorc0jtFqxuHltNSe
bw4d48aEE5/YDm8BGZuSJjemxuttgfYlJyLgHEnv/v+ldRf2rTRYX42KVTG29ooi
9y7o1w74+o10TKromvJIEACvXLThrOZqgvLV3VG6XjTwGWf+mbDGAJmVrzPj82aq
jAAqWkSZ36qzJwb4VcdYEjNufXLFJuk+Bmj6EnTAOa8NAs43IcgY1ZbTNb+Tg6Yo
zHIkK+IbXgI7MEwDPgTom0KqYN/2TePs8iUaFEAaCjhDRg6L6w01s0bybUUNqcgf
NdhIScbNYLWzd79q2JnPuS94SPSK9C5ndZ8YsINvKsiZOZIMUL4oQCtr1kRUa5+F
T8aY0ULK2P8mUaEYYeBUfuqDf5Mr2dySL/N48MxdhmAfWAoXN9rz2caCtkCL+6El
UWnVqGr7Wdyi3MRkd8xFBaVxIWFNqMyxWao9OLvLKJGpQX4UgKKCblXpjw0vTzCx
jK1tc2a6yHaa9Y+E7xsZo4lwZv44/fxOl1OOlAoDjGK3FBVV/M0VmdcnrDfmB5LO
xuXUxn8+a/93q3qVQv9IWWpDmp6Re4j1YAya75jLFPopWqSTup3IgiK4ZgSadX5l
Q+aWZ2pKKBEm/HK652JXujLxTpIzvHAso+tHku4QB6dXJd18X+63zYgVBcgtb4LX
YJRkx4oqLDFjt4RIOoG9324SDjXobxpmyq7tS7FyHXyluIeK3evSQXxKxeOF0mqN
zdIn9C28HMxHJb7k/syDeTJfyHWzYnZwqZg4i6rLBefgayxCWc81CldYwM8uAWMM
efxgqBCQZzGWWoEpNQ/OXtxnPzT32IrLCJFnNHDjekwqy6mNaloQjk6hE2hY0bq5
LJjNV9yDrUe3ZYrpFmBXkGQR3a34HteabaU6xyHpHjM/M4qtDX73DjCx8sWr3leN
/lO88FhWdQoSRlbbHhTyTSILqrDeHXuk0RFplTqiqrAWZDIiOQGPIeDsOb81p557
PtVA+oD5bk/sLeJqtH8YxeQUkaAhOlifFlGxs6ZaAJOHugE92TqFZTs/+TMmp15O
VF6dSZ7SMFOonXxr849lU4IP0WtOPOqFhIGjyysEJTyQIKH8zWtwxvmlagUlKWti
476Ore/PK32sH8HuS7p7uPGX8xk6IiHk05xzoYnKkDlII7CpLVv7t2myGnnnptnx
fmAvhU/VlBDRkKWlvytEpX6TLu1WfZpn/pIU5776Lr1jYqiJl52G42dvcBRokLya
+xB1bpRgGI6dAl99sZc4tLKk3nlMT7rzUl0JpkcIMOQ2oTBULhU8bxCus+yZ0MgF
OHRe/8cOpoxvqag6RBgXi5EvRYX/71FBWi6J+hro+Q7CYA/TSlSkpmJubqLdhOg5
lj7YYfALYwNq1nOvMpVxCOnSFOcRZT50KqoE6Ba46eugotfOhdNjEBi5AbnJZTGj
88ooih8AerF0h8j3NgjonnI/5g2iCu0tSHV5wpDOK2k3ESDkZ+hMoRKnJpgJ2xVo
bWRUKbHb4KT0XkqnOh+xW+sgvcdbu4cb+MItqh9MtNJN+Rpllm1XkuI0+pff9Zyf
XodOewMveMDMhywAEfcVgFj5wQc5HUYoq0O4CuqdEH6IBjme4ejsiHO31g15jVYK
B4fzam9CSPUwcnMjJsrccu4OngHt0b+umaSdst2T23WTFW9XNkEDNokEKJLsD9I4
49cy7aL3+gGl126XSuZv3nS25ob279B3JtYEoJ0ieDC62y0JyVmEnHT8rJO3DrfN
6xltnVgnndG8jRaEtiL002h8nP5yyQ5Mfm35LPe/Rp7x7u4kifNUjDyeV4ZQcTR7
/wew3G/K1m2hjTb52Y3k+K5FaRLCMLncj30a1I0+Tgf0O9KZTxDdZr9qYsOb0QEC
KTizGNsR41QJwx0UWr0pco16WlvmwyykMN4ctJLgIlw9Rmec+aiqeuQpitQ6BNqs
boLP3iywq3E4Es+fhH/bQqDcISiPhBU/WOxTzwoMpJTQ+dFrBaH9EJTPyVkvi4mi
/W7Y13RPKOf0M5yquHXY50ZJBe+mMDaR3OFO9skfIWU8lk70H0aq3bOvBXK9WraR
a8OKxnrzbjapm3MF+S+yfhIHtY1viTHaZKgkV6fz+tTX1htaFNSerP8jgx8zOU1R
O+snXKkz5Z/OKqIDTLPmau73wMxV1MUC19+gHhcP5TyUL01Lrg7bMelG3xs6+Jfm
R6Bz29aOFgQMQ6j7z387I00lLAvsbPPod+wglaCch+XO0XQEoPqBEtEe++Zm4eZ0
6E9+OyLB7NUflFz1PsApFEno4CQNagQCVhDpODL8/hTR9X1q773eTbakCfyPkdxL
dos7uIPWKoX2+shZ5KUfr6n0CmhLvzW81Lq2mnhSEb5h5ao/XKjeki3IxFZkTBUV
CRlsopDe3bOtImj6HPPPOzaXp9gr3fVPh/iTiNGvLO+l2d0fZlwBZPnahDjQPD8n
M5mJspks8Lui9QUErZno1BL93zKlPiN+Dsfaev6kQJsQ5ffpdwPSdUY54od9QrI6
ui6PUTAEk4Jfv/IzWver/MTsjE28q2a0513MkX50IVsycZIZ1ubvMAiqQg7hRrmY
0FUbCnUYwmswiAOWOuS2+9v8me2vmbhnQljPZL7wlaijxP/eagpDyKEwk6hdsZZG
yf40C7/H5NrvUgcf4jnv4r2+zBbWHXAcIUuQFUpv3CoF3UHIBSrtX6CqNpIAS3Es
Tduj0CeywE0dDU6+W8QZtWRMGJUDM8stv84jmYtAsbxMR5qiJs0xbE8r/SNWngY1
wEUAcj0YapnJPOaPMN0nLWDYyO2rEUc9QQ1JjtJ902c8iYs07A/K41fgBtlXNn/z
rZng6wAKpVMwYRjyRKaE+B+sbGGTIORSI9ii6r3B++nnYg9Fr75Q+HfkMS0ovzqq
cdsqAQdUIhkD7nXyF7mPNxyKVOwqyevCmBM58PN6s7GtVdo3EIN6vTRL1WcWz5za
gyA/jr/gjymqXJRSisDngjJwa2g7dZ1/WqGHj8P+5wOb4J6TCVSuakGgwXcnYagR
iM+ZSO2PDrqrDGp4SxzPw+d2cPC9ydi3z69MjrK0JCjB2/uYgOH7sS0CkMe7zYvJ
s/nShO+Al2Nk2y5dn/DdrI3zgXgod33aD+1ijw4hmkFNLHwz2srIvsN8MuTSOIZa
XXtBVEy/KQqhSw4LC+SQbosnN1YWO1B2ZJnAPjSXipXpNi8xkY38tUw65wyObTu5
4C2j3h3MBkeORiz26OFxB177TtP2yfMXqo9TDrQYRrCi+ZCwCUpfV19JG5Zcydm0
SXuGTySISp/+0zF41WK/zYiK0YW5gsJf1DKt8kOveto8uWlCyLtGzUBRX6HGOtYo
7bN3jmu01LDXiJTF5OCe+rwYo2rWDcCWXkGDW2QgB+Z0mHGhOlkl2Xsq4jlRa6mD
yoOrA2owXHPRuHraq7WGChA7EZ1SbVmGff9nfOTfW4cXgKvWnu7iSDDZkP2wnOm2
0WWqoACpl5AxRCWZLG+ve2HdqKcM50ujAdElM9vvxldw3/iPbDybHiBXZ4B1jgZA
7YBsKAmBSzKShW7Z+Pkvg6pbplcvCsLDz/xSpJgGzVucR9HzodOJqX9uDFihVkH0
caPHJAWhSr9+5bk0hrhZbD75AwqfhyarXJf4VI3WVW/tfBaUuhCIbcKHemzNywRU
LYkch5LTzUs0OLwDKxnRuOJIk0KN2KQQ5uaF3NhZf7peDuwbbBRGmPBkBKT46aE7
5acdUievo62BzrD+Jd5YpVUGGM+RbGmpNVGP1e0+2VkxhiXq07wvQl0ZsY7kD//D
hdorOcmfEdmLTt0JyuwtxQb+rB9K4uQgBQQdugw8P9cvWe57uF4H3ae5Yj25U52V
wSlGjVKVO4khFHcj1L6ad9vhnpUxoSfT2BAp/kwn9/1SerQApvVd8BqpVo9t70zI
W/WnZU0ofgluA51r6e9mHK0dS9TP2FxZsCQBp9N6t/pUrawVXFzWnjnCFACi4Vg/
eSMNPdWyyVFgU0lqG6P6iPmoUDTXkJSDLFKHK8BORpuakRjdjhDLxsZAP2NO5IXr
N9kiUOVX1+GgPXTd5LBmhxPf2U/yI+lNhw4a2QbxjBeB0JFht81FaPXiN8HvX6Cy
0OXKMZUsm8dmrBz4pEq7ypAENSnIhUr3NoP3s+FsI+dFKiJ6ksmD9oqrTkIdWfXk
wDsawkH6jLOepbnel8b6VA5TAPTPUZF6tbdNW7f+wRum//MyflDwqi90Pdx1hJUd
g3FZ8GYWd/m5UETlHHs4nJXgJ+MSY8lH/Gt8mNY3ky9OI0VL4qm9r2MpfgQ/AWdD
AXV3vY7xdPpGN3PdJrTAaIsgrWiNcyQAEQFS1HFoONRknTn1fUEOgJzWoNFqPrtn
H03U1MIpsEy/XM+obh7AvSEwNbHjelLti+PwEbUg3DnPuqkUU234/8mRsMrzhkAO
2xqWwWyHg7QvQVcZWMNEGsin5EEikIUVg8GEMTViM9TZ+aeY4WfTkyCNZh9NU0ei
r77EoEDGEQIPT3C2sIN3E0M47xXs1ZIhpHM0uWs8fcOgzs6kKXJcLQ/bbshYAUUY
QEagGuwu6GLqNOYFpkUAs67CpjFC2P1LWem61lhil5/q3OQpuK7ziVmWtJwRL+ae
ItEu0wYITOMKiUzRyPi7MqmbxLlngWdmGXuMxzGF/7WntfSN1u2ACDsYPRAHJ7XQ
PZjLLDx58hAQVAYTXuYJzQGT1SRIrdA2nKPwihhvidPqX3yIX568kKDRPUQNJhuK
lTa5U+Du1vO9OyCwEv7zN735ZdLVWrMzR4ownTMB1mbmGDo/4A9/5NFf0OxhHH/g
sOmMq2D+VyNpXGM4VHWmhTAFVDWhZb/YMGawEe4IXOZU/xlHIAlDx1Opk3erev2p
gS3mB2rskYJW/2CA9SSALfCA04BJSk8OQ6racxRI8MaQe/RUuMyabonw7zrQB7Vy
K/W9SBUUJ2csdh+5hxEzmmDa9dVoJtGw2D72VGRN/+GwtplUVTUAr5AI+BQdGhoV
pL5CfS8p/ykOI9Qu49AvXUr1GSAt9VQeWxpcjq7Xb2VGHS6BleKZfoe8ku0ujEVg
LSYFAU8lY64Qy2DOot9DnPO//9fwR9aAmoz7i0HGA6dcx1V/rA2VglbGCSIk4nUG
aW3Qdelp9pnPdiixuYXgXk/DL5euYKdqXD6UfOcoqMOAmkWREbVWGXWjgBX5DZz2
q34S13Dq+qMY1N1II4KljzaAhqsEKXbpAhM1+Zq/HsJf8jUb0LkuD/IqvbgV7EB6
EI2AU+gZA9HWyFErbXT3Of9fgzIC9wqiontBjK8vaJY4KzjPAFWKtBpVlkON11XO
McABTp9wmrr2PQSZ3Qd1fVcTcRZ9LlgMv16eo0KG9uCf/9OrQnv4QkMB9upx6y0u
3BHW0ZnuvYKOgeX8oMyy/nfGmiTc/oq31kbU5N5X8Lfk3EvY+bAHP9FdQ5ghgJxI
ntCOEcjwgCSFLmK1sWd8zY6DyvH3FujAfvby0EawOEHtwNEFAJWYF8RSevMYz52+
QHcZ4qow8nB00OVAPcSc+kDHZWu8+3roaj55MY5V5zJZfQqEjdNA+BbH6FneComr
Dh5Pqu5dtzdvEuMqPI5rKhKW1OWvDnNNh1vNW21uYUZ4rDAGf3pz0rjgzr1pI3JU
JpoRP4w/S1zKQWbhT+0REzjImx3nkSAKG6YHKDcgOkJ7/nuHRxA+Kwa0JCNx0E8l
3BbG4I2tChTj+9IRzgS8FIovemy8I8BLrMahquJGJ9voe1H9Q4VOh+tFcA2H0Yep
CBTQAGFLb8zfoCUzLLdhkyCCsyQGeGBKDgdVwXhOqoNq47ZYI8ur5ROtVOclXJB7
Q5220qnWSUbE9315f3PDRRD7BtIbEsmk8GxvjnGR64Pyaiy5zZ02B9JSj3s5xSqz
IxFH4zVIVrtk/J3Gg1E4GcESNVhqZk+aBWrajvcTpDrFXjvfEy08Z4ZaTJPL/eaX
JR7SrJnWJ8+8d7HNhB0hmc9L1pa7gxbgqhvbsZefPHPKkTt9N/8lIasHgWHFFb3N
bTZPGwho2UGGjTl6k2EkfNxnk74eq6sCIeuhFn7ykgFZ4IOr13cRpva5TOOOTCVx
OxCuJrDkzq5eKVQaAQ1HDB1wgL068FaBed657ISdAatjw/aqzDLNsHxYVYGDOINK
4bR1DlzszYJn8F/TcX+vPDqdM9jBV8SfRLTe3J7exIXyncrw+Ei4RgHMkgxEzdhk
uwXIk6JarNRvunJ1+nMAaQc4pq/WKjudwoNgdJ1Bh4WpbPHluGTL7XytvlEHjiGT
Fms13/y7tV+ydJwoXc4Uq6T52JnnG6XmsnWb7/R3iPQ86+Gz65lU2RhaUr95jtIw
uYOb4S1oYZfrVVP4N593yBEVh5y6JvFzdoRwGHuP36eYIh6rUZPXou4DsMKZXNau
GfyTn13s0hhWuDlxrKLApg3ZYlcUdjWG48WNZw4BvGKk5l87LapeiBu+Xf/ZmhLl
sEpTDOP+yt/hqOOjm+o5QZdA/6nylf5tTe/Xo7szo1Id16iwWWxl/i904SHgH0uy
TOamIqYR7z8ES7j0GepY1TgiidTHAUmgwVDNSqCVpUpJHi4sYv4XaWs0EDQCxx/V
uuWJimF4l6DOYqzTWk0bvcRrJxvxP1raBlMppvgaQ3OSQ+kFkZlQ76Cw+pxqLXut
sK2/8BzTP3Rer+n+JKQH7NlSDIqqr2kSxeeW9FztAT/n+Ofc+bMPq+E2G9bBN9FF
cMIa3FY800qDdvX3AdV4Go07H6AALlzY5CqLlFYtZmO5b3iFqN483ku1hgfmRx2E
8Tc/wVB+dVpTrdFP15sjVGG0ADZgW28Nf78RdUbZ9nAzb9P8V3ftDsdB6u6W+nVt
awCQ8khj69MiJVslEqdLitpmgv3VZXaTV8ud1/GWpcOXiPyndfzxBkEFGZ4p91Rh
H+AotMgKWItd+qmV2FA5bcutsCzVc68keDXTCoXYs1EnG5RNyX5/+7HYoOGeu5l/
QTdYVZ+DyCrK+wAdXk/NfOlw49IxXg8C1HH2+qBOKBzYCc7CN+9JumvUTd3qY06k
9k2o8LhFDRnZ/zFmsLftbXXpJ/qdJxrcutOaJDBQoA3al+a49a6/Mepg2IUm4040
U6ejDGmrqVRz8dtBDJmpa4blp1T50Wepak7R6GbpW+9ZaaqfsCBaHfG2LRKVc+E6
rlHKXtrWy1GHspC88eYixD6yMzCiSqhYzmZSvQPIfGS44DWvHptWv6MkGdoexqug
6u6J1lc5QhU27fQUGFYSTP5WOk50OttULlbQPPRfdShLEIGyD9pxoOX8FGbZVBGH
9pxSfWyp8glo0rDUUHzoT+HQ/Hvv4ihfAZOKCRYJdEHDnX0AoOoWuKR/afbtSha3
efLyRkqcHOwurDizy4gvNK/bjCrIryYsB40YmNIunLhUH3sJvdIIhUHsNVZrA5hf
dxQCh0Pn4ay5YOqwSGszs/9pL8kZiAQkp5D5S/+wLUlU21+aS3kCpiFHFtObKZhk
05RC+8lU0RHcSvT698xjHSOs5Rm5Umh7Vr9EcHo7XOF/WIRWDGlKUgFiQB7oZ0S/
WlNtdBGuZmjABI0DGpYQMaFefDwA469inA4MHkPdY7FcffrSZhz7datDHCoy2H56
VmPqK1vu67dUjHAjrI9g+QooIcQKxvZbHBAflmVERD6lJAcvDXpgeF0+VAXc4CK6
eoFI+M/D+MvEzhPBuAMdutGM5Ugq1RMhp/90oyM3NPd+jPgoXNvoCxYlme9DIvjy
7mjn//hxvoBu89O6zAtq5a/nmabLrq42KE0LYW8r2ebZh9jFaPkWiS23hp5YIATy
cKZRiWzTkk25cyXpJQppIVdcZbaPNkC5IesZCIDW6z95/kIE0W0XqrYzF9hnSfLz
8fskQ3/fZIsGHNz6n0xy6fvmCUIYhvF+tIw9/aCoaNOM538003vox14FzNTjrUK5
WdbzPc5P1taOUyHbrGiBeIzaNhk3iRB+xOappjzefLNuTaeUqbX4rqNbzLo0xaT1
HeckyssEUfWSJFfPRn86cEHne6vzI0mf1JIpH3jngQH1E6VsIZgQG+Q1F0m10cPo
ucyIBlhTYAc2nv6AkR9dJgctBjcy9VlioUXk68S3yleUZ72FyrD9oDc8xfUesC1E
nGTuczV8xpdAequItSUPKzBRNaNj+WEopm8VhcYsj3pa38LMDLE/8uIRwfkqsFQi
yDz/8x+4BSVrkYxH2RslrAuEO85wTF9bm/g/8ydoh0MZewySDBMJx7PdvSvSeZ9D
do/ZBxYmoVwFhxGHm3L0CnMphKmo9XJScanuD+L8Jsacabo4YsfmWMluYYRfz2+H
K8IWv+r8ZoyNQ/6jKrNY8T1NTnwHETaig+m1Yqq0AFaGEHYJzeegY5V4M6khtA9E
YZtYc4n6fIrhGWt9IMbrqo06KiktkiLt6iQ2eC7tMxaHZ+y5HPgrWRp9IIQXkYpO
4vzAjXea/tfGuVVRV7Mwfl+77OWiHGW02cRFqouEqN+3GF+JQ0JS/eJJ+bFb92nc
pb0p3qW100IhghbO2VY/mqO/ALUl+dW4KmON9fR+s7DpgvoBMDs6MSmUsaaDj2nC
Or0f60UTwZjJTz/Po5AK1WQxatG8T9PhwR5MrHb/VvmQWF6QpIqqmZTrMC4IBp+5
UPj9SFWdhyd6pRK3vfrl857gFmQMqddte0nrha93rZe4zVfSd4RVzSqo6fQIr5IJ
F75/5NG8LS2ls1spweMdeMzB3Qxs8RRpMwdPKw9baSPejHcB303df3skpE9RX8dq
a49T/uOz2sVmqsAKKtR7h5ar+SHedHe8o7ytBzlg5NK2ejy8XD/9b3LpKkofVpbs
by/SmJyun99lwY2WZTlbP3tUmM1c1IjJs+x6r9uCcTR7QROGW/JVK+6vdMRqlfDU
vZesJq5BBV1W2WBPoOE6ctSqhM6KDBBx74x9fermo+Ivue9akJwWyRbqP2O1INKF
glybq5SwNKS7PBinGoPtpXLDmvZb2zphKm2opHlEU7hyhLEL8k5sLZRHJuaxQ1YO
7h3kgvOS7gEq0mJfFDg1lJtLVcJLwICs9hnLYXTB2xE/ZQbFgxBYMxtK2vkgztt5
rHMkovYMMK+HEnuh/ha43BumYdVDaYK++NAOIepmfftannbRQ6WQui/+3OZX8834
hXuoIwK3UhmCHTnC96JoxdYSyvtNGlVOvbBX/6sFqbGZ5pafUqFaQ1k32t6xPhtd
/7geoDSiboTEtQFnp2FryRGNHFjvgyFYEF8VIA+ar5mIdbj8LHEhlkbStB5mpKSS
feO+xP+u/U5/MzBXYvA8rQEAXzoAnVLJfLP4J2MeGD/bVNoc/rTvIUrCgAU8/odX
cTD2wdkwNOtDkt9woFaMjkv3xZufe+o8kdrG2ArxMGHqdmG4Rx1KYoG+pS3id2Nw
3wPsMhiB/as21+VSTpARLkMCjkhs5J9XB2CGtv+wHKYD3ERAGOdHnPU88o2/vaGl
hOEDQPenzziRPg2/XAhiTMGL/Rmh3suY2X1819Ps9QMVRmRsWliyX5loBIl0CwKW
eKjRcBN9ZyzUcK3dpoAoTuytmL4QbkDHrpn7gTrceaKAhPeQx+7B/HpjPfraDlJb
7K1wBArIAw7iifgDNd/dEskO2+OliaKrQkKqbqBKEsEbOuGRXkNCNsY8i0JZ+O8+
fHjo14wpzCKsxuWYwuFz/bzwNMeif7J31VtldSk0anK/q7K23HLs/sRFJ6ueAOCZ
BfmRCFHUZ51+O7kcwYMqpPVUDyPvnjJaJw1X72n9QNogIE6C6BmDsJunNtTPfeAj
+C/aM+o+EYP/zFZyiq/mpMr6s/PcemLyb6bZhVr/E/5fDP7YG9Lins+XfsAB05GO
VN84+T5C5wjAlHe0jK4eJakhdqRxOlkr15Y81ybihbPoKL8Kvvm5i03AeMqoAo8g
ji8p8VZWBpdEJsTo3zmb9YJ1TWEutLCrJZ9N2kBcp95m9+BpjeTT6tybQCO3Bdrq
7HM2aS5pud+Gvv3CKN1f5I3kXsU/A/PxPdT2y0bMF/oBRnLNA5fReIfUDpovolus
gY359U1mSmYgYP7yRXXwxYi4afKPAlFXfw35i01SaWN8PS2/RuGHOgkYBRCXRc4+
u9s2KzpEFLJgtQF92nj8OdkFj1vJDsQuYLAFc6kiFr/XHzlqX2IKAN0ARsQ1Un2K
ExRoZA2QIa4bFkij9zM+5tTL9S9l2sYhU26Pp2ebvBAr/+Bahr1jShBxGa1YcTas
pw/fh1omTM5P7b8Y+xyJUZIuEIez/PFXLvTOrfLuFraMA0RHprRW9xsqkPQIpnMh
E0vTvGvUkPv2p5JWjhhTzWwwz+/cM4ukiEN6l1ploBb3IdUCGkl6o5tepMBWFcIJ
uitm0LLXDvuOrSq7oTs/V839m3gxog4Gn3gmGr9/of6u9jBs1BECERClgQKBn+HV
08emWTYFSJG1S9vXbiGMbdrPklgW+1dzOiTTOEeUZ0tyoSwxnB9avjvVkMYSwTp7
6jKJc+NeMfO22jLtgMDcPlwkaF5Mi0ff9+lDl6gzlfkRaOTAT0DfEEJbb5eAozL1
9PS2uSSwQL6vrRmwLnpGGsc+2/Al++td5HgngeCSLMmn0CU/hDlZQqJ/qR670cpz
yZbYSokE8zzVTY+cmv0Csjw0vfdH5t6w30eEfxX04ef4dwNOukMZJ7Aw3LKh/WvU
PU1fIBRmcNFt8vJqwj4s3fmn0JOa6inj7+1+mb12D67DEhv329QRuWe3pzIzb1OH
WLtvkCYMgHHgiQmvaY+1c0QwyVqGHAgsLLnw+okfc6wsIEs6jZBZmURsXec6cXFc
8WvjoNWlsTstnzNuJc2CQP9t/gbmcXd78iYFarrB0HEn8y3eNmsG/UL71Q52oMxR
q7IjmNZap8oXuPHT7yyjn07RHlNkdtx5N1KRIfQeeJikvxesjRC2hZywqUdz7vFa
BfkgZUdjfzIOS17EXjNsvO8Jo65xkeY7TIzuLJ/4sah4S5eiqAfOroSetZrq9/oT
xxT9kBrkHV+lkkqihs6nVBdseM/h2g6arqLI4fvxyKqm555648Yj7yzgARmjGZhg
0L0eWRnWAg4CHsuE1BTMG4H6LJnVxC1jsdK1/GKCkr6oObQJGEyNADZlK1iy1jKz
sREHF1VgFAlJZxIMrx5YxnN0EGH7ZyWYkzkAqh1miXtT56qi+FuRh7PL3BpTWqWY
rN7X5Zq//3GRlo6RzO1JSshoh5wbzY/bkxCvWqN1jpeNd9FTohRHre4mvZ2+qP9/
tC3J5XMAtVMukUKnySJBJg2fEL+AAukt0PxV3Ogo6XHXnK35ig1fIerDDsZE9mRo
oLbRwzYyH4WqwNecpEd3pQzhjgQ1h2oriBUxcmeAZN58gHcLOc7lU+D3SaiXggBc
IED19qrlUZ09/jaQ6kf36JBQOHOglnEoqNPoX0tU2EGu/nhkgW0rg0kK83D4OtEr
5zy4r49dKW3aSoAtjaarXvyQq6d6TyJHN6pXdUfxezES7jIcLT0Rs2h1lGWA8m8f
g4ioAlSSThAfoaKTw50Zfi2mY8LdbraxN6tTLi7o6XYW/xvFtptxvzfxh6aE/27s
R+ySCf8C0OdJQcCaqSn9IWhAo9ji2YyNazRu4JoqdqiXJotsOQ88ghz15VPjZLxz
mZNfzJiSQgT+DSHT1DX3YetN/h1Yz8thEkMPQRmZE9a2MHGNJKQSeyzOu4KqbRp/
AdEoDDLYLJoJ+uHKeIhTjwIWTSSOpw4stB/gzMGx3+jvCSJwPk0yJE85OCeh9vwb
Qqdw4QcHWQ4YTnIUpY3Py1OHhn5OPqEuu++DlZWWA3ADZRJNqlV1xpTFi/W+12lb
fNq2jbBmV7ulI80MIxnwMOVjIO/gkgD5kb4ucl+sgJ+VVqn/cs2sNx7HjqC18FWB
DCuLmkL9v/nFKwT3rUPyboUAjO/pvGcE9IdpK+4vvOKolYJOTCosd8OIp0Hw0ebh
d4/KitoA8TqWFcmleAgVA/elUHP0+gz4YyZZEvzE3K9T1zLYVnAB8DtIvWNgpt1D
ZcQqdsLyIAZ3bcLgBltEgYNEsiUdgV22K5q4t6Dt2U3kr3wr5lesHQpW7ZQf87nR
F6f+z/wNMMlGREDHaLDe4y2fVEJieqNzE94yUWXrnPPHUUtWKyq/n0fUOsfD6WSy
tbkBnzj64zNDgdULDsabEaG3q+PznTXb5zjjApsBkUIe+wltwFgTlVS78FCQ22HO
+3l30aOxd4BA5azrpLaHyAeUyY6iv33EEXQhsyhmeyBFLpxEU9HglUT7atS3rDwC
ILNf8WEhgUP+rBxcMtKS8b6dlLpyeesnYdNTufMXQ/PFiS7f/fKkIOJBZweec1i8
0z7vxc9l5mwAPduzYMGYFJEhYoOX+307NvPbx089vm1u2/h16NCy2qUH0JiG+VwV
Nfad0SMCzwj3Iyn+SHInuZovLy9vPE3cKAF3lpvkyCA7t2wqHqkqjOr4udWEkPla
zjyZK9DNMp/W5MrQ7t5jbQ9WHVEeumDIeTollzPJ6sAeDmhviDVwT4BruzK3ZiUT
MomCra0achY483ztwH8JpUKlwAMSs3bAKWQp/7ediuqKc4p0u5SPZG6rwZqzIwwO
+uhKJxYV7rncSqLIQLOaIvPJpNixS/JcZQVTcIf/rnNIa4iLDDDHr4TcMb7BlmGl
y7oA9SVPNveG/e3VBbaJMazqzjwDbP5u2sHczTw3DTRjiCDFdzC0x3BSTHt6rNHC
FQys9FXDwIx4wprtG0iwUt+LAm6B9AsluzwJgduawfZubZzMjPXjX9yWZQXjwPae
OvLf8gHIkjIqMsRi0zpb+5t4im6DpMNCYp+TL5JPCN5wI57zA71O4Umu4MCNcEnP
Q+6uYvtG1aAkgCdrrbTNAzfne48dcAPrhF8K8CQyxezOpCtScL/y2PCg5yRo+PPR
X1A28YS+bEefZsfasPoIKYxRJXTYF5BxZNLF06n4Op8jxxNUIpnQLqGmI/00Lc9O
TZmAvPcZKiMhXAQhvqkTBzy4p9naBFHtjFyMUYHD5HltvRslNio/wvtSc2tD2bEg
GEF+yReQRIKJWcC7O4mnUa1Vo1fNYNVDoB2Wbw9qoJ+UpWWoZCT3ztHNtNX0l2yo
xWtWb1+p7Va8N+CUCAs7m2dkwd2tIirCmWzMw+IIJVRCQ4JSufOG+TwaYGvdktI1
523Z7CeP0vim5YjY2jiPMiMICBt5HfNyJq4/ehgGYa+NM7sj8km5SMc6ErXQpYKg
ZutpLjnrPJkWEk+nn98PYpk2XauCqdlUdDj1dG4kVMh8cFvOmrAMhWeLXj1a0TLh
nN2IO/3EcMmsMp9soMAntWIVHidRfZaOYJ1MlewbwOEUXWTlbl2pK+er15g0CwpX
JcAcBTVRMZBqzHXfCc+nr4TbuOeR38GLyO28kZz+6RWzrA2MKOG+U3tTytyokN8u
7QM0dEM1reWKYh8HFjgaXxMikPS7nKe2GzWQ+tUWDvrnIoxuZ4FE+UR4Sa/OUFTp
ZvPsOl53XzIN+z5E7LC3p685CkzVHd9B2pGkN1of0d6EUilnJlCOZp40/VXHOmWY
l19VOZdXiaw0KBxhLWPbtE1HEL63t2Y0VY9xW/uUHYM4M9WpI2M7u6itvfm3JdPO
pA/wy8iFv579RK3Bwr8SfrxTBSSdMjSGuHPH8js64B9m/BIIFd4n9nwfPAY6i6gJ
mhNmi9llMpbp3o8ikUk7AhX2YGce/iXzS1u9jacMwTMmzwJrq/nKfRF6M5/vHAz7
il+4HGK39nuMIXHE5O+J6fBfy3+1jf/wqzYv/V4xOUpZaEUjV9nNwMSbE9ChEydS
VQ+GpdS75m1tfju7hJDsVzPecuVUhi8bWvfHplppHLPQZpAy2G9sjmkk0bd5wX3z
JZizNY+r25t/pjCwRPZRwlCfhk953S6ltD368qqp0/+3H9XvoT96n6ooXUCXdfTU
3487UBub8v6Tjp1OaOAH8ehZnmmeKPjkrkKDZ79GkzUxlwHJBjXOb+KkhoZsUuQY
Xn097heFW8XsXuEAUq30moQRK5IUG3hucxpbL5N30KpAsdXOkh27snQyugYfjcc9
D3kIwpjemYvtpnf95zsN1zdwN9LiWas1yzMwf+QUnn5swmR17/B4nk+kmRA00q2a
mkweafMtcZbv/NUUJaObq1cAPGMMaKSyuxUSyrN77rutS8jB7EJx3eGUtvStFcED
TlrrDl+y3AGabd30PEPtTqf8q3e78Yqcyk3/HptFckjtcAJeYgnWv5yJJs593qg9
KOCifnTxsmDvtjG3wFMVCn8ePK9qudxy4FmD3VqLaPEfgOx16Wgb6xQZIAVuJ45f
CB8CvhniIhiz8q7Z2Ywp4Viyj1AvflsseyAlJV75iHGyBFF6UvPcPg0MzlXW/ndP
VF7KMfoMKXBNQ1If3haLS+qEmiOIFFGR/GInCsa0mSBAZ15LIKIl6G1arUSBlb7Q
p/GvL2PU1MTC5V8E4GdWqoACBu4eX+0AEaY/+KjRxWplDJnDdNau6Mt90lYP2/iT
vJQDyMZDM5QJQrEvq+T70K7r/FDyYcc2+ABnFuOwnOy23gHqNzqV5PMG1R6YkGpm
Rj9xlrNlA/u9JcAjnDD4yNmZPagxGbouamPVFLqI5R0bKXeSdx6A/CKMJP3Q8YVK
+wY6amdSI2zLpgKoqjWsrwEThDfkxJgvEnxhDNsBNSvw03g1H0J15kBGwI4NlKXW
Qyr2AbsAfzg+cFvkTfJ8naCjGeuzCXZO3VeI2Urod4bweMlQ+1hh809EIvz51+xC
GTBwfeWnKzFL3X/oVfOTCT64aeZRnSrQtAwPWaKWqMmzgCTEG7cnnpPoZWNsBrOF
EeJrCSl9qsO7OotDxr8dLrZVDEa3j1h0knyBIO2lU+1cbrWDF0VQUQmE0g+ccZkI
DhuCa8mqZOEkUFzNsvzcyM1zgXGyUqXbMlTRU7v3PQROILTv/hPmeD8Gh303S+0o
CxrraI+LJBXm2gb5djdWKqnuZmqwaMB51cIlmcxIZAgbWTof/opt0pYMSgnGtXCt
RUQD7i7C4rxySulPb/Jg+zY1y7HhAUcxpltscbnJF+TaOjSyhujsXvov0Y0uKhPx
GZsbWySPU77JujbomjUuimgIfF39FZEojlLHTGLlaPIZGrYYp3Yiq+BDmzJPmMXO
hQ2SO5k9fLTV3Z0CHr22BIbuI/nDs2xizDUdGb52IzNVrfjsbLFF/c1LxMRwPsZO
+mhnHCBdSYE3cHXSzt7IAerICPwaDsaDOTz9etPldsYzJqJqx/NWdpPsjadkFhf3
f4pciFHPmV5TQKZJdm0y50P5D7A8BGD/JI9WXnJCM7ySnTX4sh1npgR/+Fo2Y4c9
gtIn3wnobMh+gdoN3jt6uNFoHaWgLVG9HGHRIJh3VSLGo5zjQWirDRM9cyOJdF0A
zoDSEvcXVDHv3ZEZe1tv9Th6inA4LTu40JBOoz9m+6Lb8Ldd7aE+n3mDlvfS7a0g
bgUh72P/6Xs4CaXZ7/ZcKPwCLUbuCXPOAA/7bBMb9U0oFUol+ZXBP2dUGf9HPwx5
qBpfmJ1bEAWoHSD/WKy4IMogyCYm59gmSterr11OHyw+4+OvhyLJ0gsuH7i61POF
JoFY3upI5nDtD+KmxJg38zT0+MQHKmDCYkWQyvup845vYYDJYbJ0gedXSGdFzxzD
yyL5tAOqlogyWDjeR3b9uOgyPf6DoEm9lgs5/15VdImwTycr6p2j9OYibiLs0HdG
s63KSpWZXWHvpAILNBortadQS97QGG9VeLNXevHvcCwxF508oxCUGZqZP63gWeRq
N8PsnQu+dRzRLOSK/w9jzmhYq2X80eN4j3fILk9wQINaFykzE9zYuHsOYfrd8oRj
r9UhndVefz5YYpyu44cs8rq11+/PbDh2HxwTSDPd9hJGrChZNzaLURfPqOkQuCnA
Mf1Y5G9xAUoubXU9W1KBl3pDYhKi0TQFDGXBIDbaxFOuhAWmuSO13hn94Ro3FlmB
VNWVRmywWNlWchu75ln84dnOxcbQMG8BJt9RfiilN/5PuJLSht/RESxlc5tzQehM
MK1ql03HGMsHwlmNrK7jk8cLhwSOIq3vpgDhX5t+p9cKxFfrtoW2m9vT/V6Z/ABQ
2/FO+ONWlz1vWNO/0rqJInqisPbCsanFBXLeiAuDw4Nhzf+ufXAL/2SiBB0jW9Tc
QzEG3dgAEL8xnrxkKrfJomaqumzt9AwHSMOdS13pk1bmCPU6a+fT1RmfEXjc+xgQ
4UMV1FwIDEzDl/kuZcWU56CZZyh4gLrsC1+rsHNvi8v01H+KIwtbPI57igxICcGu
68ECTlYgwMAWdjYfIDj3VRnrTJSB3S+wS7sr0YRVeJWo4hJaAAwbM54RmDrY4QnS
+A40enpFvhqCWFFEMSaDDILAo7flP05Q7FmhWNGGj3ndPtfb83Njjh7HKMRiE/Me
rAUVV17FWcFk22nzGxUweopitXXi3NsuGZAn4qVa3K4QTqDGlDBgnm+U0vQeeVKX
vslO1CbF88HY8hIJnyPD5sCi7pYfiQIXREgfR1ysuWlgVhiTUibS8YA2FkqOmn5r
ODNbdytVRpG2yiUn7wAgzKFBIwMQmEDQM8Ga41cTKPKQDDa6855+JDAJMB8qq1OZ
YZlbSp6wxioE24NdsB5S+J19m4M+dgKzGrAR4f1iN2Rx7aa30heVWJVOlicxpaRT
Kyj8BESFbDEbymVNrDcZRg91L30a/HhaDQOtaqo14ZRgNQcc1G+MJGNKL0KXSkMl
rrRiBcw4tlQ7NK18GKTcMu2WncGYPTRSvZDL87ccsC0tW9CzrCC4e3N9BFeHzqNh
qG2Mdayf5Lxxn73bZzAwdbKVqjWyRNDEHG+xDq19rMc3CpNE6xpMiP40bbfO9uAL
CF+T9rcYgRkZd0QWmD8aG/2e0kFIyeRfOWBUpnHhIVf49oKJpFEkMioCAqjXvO4n
X9GAWYwj4JVULJxdZjkyG7et56PLWtELfkACkzlR83ur6qzBYdEcP1QKZ3pZrtIf
CIjAmaJFdx0kcXf7J8t/dbIF257NTmCIo8/bfnDJycVjkQ3x/2arrTj7oqJ6QrHC
mvYLKU4sY+4CtE7Y1MeTzDh5NkSDL+tEFVBuRz3dEjLhm2ATxrUvsdadmy0aZMO4
jqFtbIbUmE29kpa35P5HF4tf0/Sp5hK7NnD4F+wUVkYm2+w+NXYeCZ4rsFEKkHDG
7XtX0GGPZQNt/bjgAPDxWG+Lu3+fP94r88Os3tYKPXOq9RAeMmrG4dGfq5D6PK+w
zQx160xIwTAKnBaEjwZOS+fZmrBiSVzzKFhm5zsccXOMEup7AUvQ27ixzjqeIQZR
KT7QCISXNFSygQs64+5s9kLywIYkpc3GzXcbtVpomdilzMuH1SJ+keSkUqPCNWJR
/0rfv1Dn3T/Zgkkq4CodAT8gkYc0Qy8fgB7eBjAbNEpO9kNzIUaLRFPVzALcdq/t
39k3heDZE7FV+ufgyoG4SFNSoKy22WDhAPDXLJRdqvhHgNixXcwzFFvRvtnfqIR5
w9kejfF0G7gCslXiwja7e29qrzT9wp3kQeGAXJiPztzN0wV00Tm2kH6c8VIBaaKn
Kjp6AH6Mt1IPRZFoSx1zA/R1D/J8eHmDkJgKgV0tBuWbmazw4q5kqewYfE0orONT
gZkZwrT/yuVb7FcNY+r9uwXVSWEeVXB2FKwTvYQmxqov17zbJwIillTgVR/7Izmi
K1R+FgXPUiTs2eYuJdufGn4EhQyeQu5zK+gQs5DJsbNerg3dQTFSyqVBlgRy+y52
aMvd6ystmdNuOMq1KrddZwNmLdw0xOZsb0Qn+FvRbuP3pscokXxFK+RW0+Hd7jFT
DRJaQIgXlibfm3PeyWB4Xt8HRod4Cqk/mAt6E55FgMSzaijIziWFoC4+I/O/IhWB
xVlYKWqSLdS3VoLzYgNIkIdKargG9yGP6Uof1SznMtsaup1jTJACkIfT+0WPwayb
p8ZlRHT+n1FJfhaSKCUC8LgBtv3rWsXTA1uDckp6jjOOS+SjXZrmyz6tnShFsSTy
ecfLZ14C5mSz2VMpMO23Gtr/Cf5C7uL/kIprC+nvGhQNFLeA6f6pmhG6uRHr65ge
gA38i5StV5CSt3A9V19xIqB0LqWC7huCah5rqkQXz2Wl+8IqVnDeBDvpQHvJGIsB
ScARk8K0mHaCU/WN4tqRKuhrKeFYauDCn+/+6jN4Imj1f6c7PrBbKRoaqVP6t+BC
+mt0yjRn0O7R0tzIGj7WN+jA3dyG0ocmc9vK6L9kLL+cwOMhNcQYbob5424tNaG7
PbS64mWDYNVOVB11iPCDemUdXvBxFd1kzr1IgnpT596l7RjqAJsOCE6jCiTzeucc
u5d3epjy7slqQJwEu4nagxOE9VSnk/+sJCB/tggN76QJ40xOqehAbnmpq2g7T5px
A5fBUbpkKLInQ9RnL7rmGMp0OprnfW5pZovOJVDwCU1uM2eKDiN1vlnkBquZ4azX
AI+6nCal7+2BU2Zh3zPlt+ltzsnauWlodx55IPc+tw4=
`protect END_PROTECTED
