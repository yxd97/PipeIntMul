`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BNiXPYt5pt72M9kbk29kIZPh/5fIyxFT82/StR4cecBlA141HrZoRcORTW3nmKyn
a7jDHQH4yM1OR0R0XNz5/PM+Zuj4kDG+WVaSFWSRO4KicAz9X9UnEo3wePzDc1an
kMwSajZOk+/S1l3XSHs7VOqHAraSDVUlw/61Ake2YK218dTYeIX+mqUt1HI+hpO0
3Nab3QQdAN5GvuBs62kvhgXAaA63muTmT4f3Wqg6c53gaU54a4BCr/1+FbiL8zTE
FsH8jzWuNCzS2UrYnURQc79MFnE41cssUHlhdLmpsKNiffKZfjlQaA0oYQMbNClb
Rt6rPaw3lRXvRferzDuKeJum1bpvZdxx5GhadXHTIRpCDfewigEWKyXxNGLg5Lu/
5ISTX9Na6jG5rQOtxbcpIv1rtU/lvzBDOk+DI8VqkvIQCwSnxz2lapiWKSisUAJh
alHGS2E3as//42AWC7+tP+VcVP1gY61bhLb9Q/RDWEbcDpUJsUSJx1smZf2oywgY
`protect END_PROTECTED
