`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rb6FHzX2Ysbj2QG++rEH4h10mxnGPIGdqAtXnDxo73ts6aKxemrDA3anCOLm1uWQ
fANXQdmcuM0XCbITmsrPgcBpPN+a9+reIoXmJ/QlXCITuq0ooCGWbuiNlwzKXZAK
hBmbUm4q9n0y0P3KhNBBgxDU+CZkdNcKAf54a57xc6a12Y2HAtjinb1p0X1nO0ZA
uuhCTyh+rN8n+4Tbz3TjBNN9MmM985QjnOHrSiCj71QVhbYpcfK6/silvAyTlVV3
wBjsvIcILYLzSM6fNh29RK3CtHOXxe292Grifuk62gkmhS6IXRf0wBnj2eh7RApA
skqhshc7cUkOPt9w9sVOB9QLrBXzqWlcF80VCyenUqsieR/NYnaaRtVoM4SKTmpd
j4XVwRdfM8sGExvG+1AC/bKGahMRWSiK1a5W517BESGkXxvYY02dI3PXyeoTt3Ah
KR0ZsWhB1fwaPpjH9HKa25d1QNsywMqbLK0lgkTtNaNkNTXvOxDi4VbLciByOLoy
xfm+RUdgYLSR1AcmE9DhoYk6bjruN8uDlGNaT1qjWrsatTaRV3NfX/O3qdUec76X
35BDc5lJOXXvDLkO+N9P7LQTAkHE5Eb55Wfyejq35L+0sv4wvgCsm1YjL8byYW9r
Ldb8n3JwKhOdX5leaf/NKA==
`protect END_PROTECTED
