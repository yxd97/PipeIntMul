`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WrpbiBDSxBvFcJzT/ESTHmKN63qtwd9XACmuYd62Pd18P8gQQC2bZarRXskKcQbj
FHHJBDJ+p8i7UPtj+aJnJ5wPXvSjb9jSOineJXVpb1az4TBVJy4Gqf1v17n2K/u1
P6jZHZgJgz7NJS2fwoZ6vBgXDn2zPuOu5CH28AZdO0G8Zg83eEDnVI/BqX4NFBmo
hspPqDeTvsJ7CPrJ3BKl5/JM4N7nA+MBcecpjgtAFTAaLcM5odJh5tbZhbTcOVam
OMVmTaPV8uW5nD5iyK/sejL1aRlRAJ3xtNgizJK2u03QNh+Gc1OHaoKMdIoDVWgk
25MQINs3kxzvh3xr6RVMLwWOJ9oYH3WIjiPnE73VUmkaZCW5I8jOQExqvQy3cmlV
CmVqVoBcKZSW1farPHlL/aG38F7GhKnG+yKRAhDbQ4vx7Tp1u55JKc42xJELeiW0
o4cvEEBOReyszSwNW4nBtPQ/vjaTRGGkcCgW4nx+HX0=
`protect END_PROTECTED
