`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a43TYuEUpVrbBQqVtokJEo5Qsrisygv059o4dWSYOK/8WduMAXV7+fFKNQhTq80k
3XzDV2s5kBGz5XewXlxXDOY50vyfImM5lHP7+GM1bRb6he9qvoWqj8FE5+/Wkq+n
wm1XRkeK9BxmVUFK8IzxfaVx1y6ysCaEZ+tAnIaRkB15XtJLWzXRNjLO2U70Cj1m
4pHSoPnl3KS3sZs9TVWmxuGPLur+EvdGT+9uEbuFQgmsj9L7KeL+JUDJ6CCgDbBH
sXUrGdcowGpRjm/w/zkG1/D4yoW2zTNrxzpiFYVG5mvpSAZadXn1L8OpsttUWHCy
PSAp/PeGWdf5oAbcvpht+qY5qmy05QKjn8HkojpVHHUGuRyePDVmEjPkWaiWG0TF
e7QaS1GJiHfqaUVaak+Njx6dbOVVeX/WyE+XckaKJ0bS5MopVx0J+cubiKkr4dAC
XfhOqJtWal7Xeh8XjutLuL+a4BgrLV22GVTj56TqheO6XOfmkodUgA7r0UeLhjKA
jwIc5bTh80ziOAyJ9xnpqU4qiMxnLfW+gajTqMAFNXvNZQ/daFRzS7YqdN8k/CY3
lTTGORpVGXbYzqtlVLPbTxznseKZyham83Pxm8174zRBL0HxIvQdNbws+6Sbq4GP
nHz4JmQ1mFnf2UxCMfaxENUjJKYXA9gWo6rTWiF2tGdHecsWF4e+riZyGs6Z4JNk
M+ym2Qvy/ix/s3lUkq2z2uT1oZPTCwU0/lzhJMQ13MfbS5KpsEQ+SJg6EAg2lYI4
2kS0kidbDOt18KHUQVFSQiirkFrNkIY+fuTrnuEEVrqLrLDSzyGQbIujEz1HVf7P
cZrOr4GlLstanpO/q2B8kUdQkaCjdeekkNDhpwknOidlCkPv1IQmeB4LlMpNkIo/
G1L5AD4mtp1qst0f0NVd8ZzzB7LlrQI+1K0E/pafgl//K6N8Ve+6ufTasZcg0zZF
qJJuAlctLhq7H3ScqJCDS/HvL/c6KEXa4uqaATjdNChNVigFgYQ44AB+2SDSVotj
TETMIUSax8AEs1EMFp+jjwCTccv0TgMwc3V8hYWDfaB6Wj8i6t1cjLeDMQvlG6xl
Ju/n1s1g8xBg87y96fPZX3obyyxpzTw0g0U1atlMFF51zdeVebfvDMRllCSmmpdq
IwiQF7/WzWHlAHaP7Czz7uSvOPnLfirViU+j3q9CCG3yxrPPs/X7tAk5MCQDYwkw
2u0EoLTSK+DijOiMTlr1gyiX4e5ZWOWUh5WSw/sOD7iOWNkiFvF53BpdeifFI3Fc
fHWlID3+AxcviwUWie2x3Bq53x9POF8qlqph+8kk1H+wn2o4dL5xZJfBdVrte3tI
jUU5lBoSANoSzz+LKbfGhVbnpK7dHkCb/ezszEpwaDPjb4sybaQULPwMWzMGADhT
baX6dGKN45kx9ycGmnZdNnicFvsxJ9q0JhWASf4uBfvGx4vn4niok1dZEL2fGety
Ea4CSgwRvjndpX9XiDZrIx7fQ4Vq/fRTf76zm8BgUR566bU67k3QEvhBGfrXb3UN
BCFdvk66McvRB2ETOnD+iQYCVBFBdb902/4N6cNLJQ2qSizWVtW1op4iKijIeMkP
2VeBK9rxIznCesodp3f7CtBmR/NwkAexGuaqiCPDHy/ll25XmEZufU2N3FkDYNpR
7yFSVw5JumspiqVVKN/WiqfkQWoJMUVr+N0IV7T2fJTAgE8VfmM6xTGwgxb9Z0UB
xKX351bowSbSMSzXTMFca2h0Aor/qfiHptsIb7y7VOOgfq6b8/lCGaT9kkosZLzy
8UJ+aHqchKO8/iqVkM8rYpZ92WJ1JM9ryPPmR6kKCzJiSHSsAv4NnwadfwEixvjx
yz+1mejNg340uNmEQ2B7LzWdLi8REm7E+Wp95Qv82BuxS3L5sa0b3oM215ijXE+F
eUIqF8Wz+Sh52XXFEZSxb44nX5tDAWLuDygk6T2EALYN+2CkiNBzp0kXT1mEn2dt
ar/J+sV130Ijs3tkpbYdbc6hdDGJreYocC+CIp9N+PDirXbIil7df1CUDCiLVthE
`protect END_PROTECTED
