`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLjN5vXkKBO9ZNxRHntDukYnQKBfNhqCDjIGhSABSC/bRrdBzc/nahBMghz/FxrE
gX8XQnf8wz+amnA+Iyor1duUuE7vCkxHdcOSeBHPzM9NbS7qz/5U/4QvNrbGpisJ
nBqklLGdAMflE+DSThQznQO8XRJ0OKW3xDbgKIHDc/J1QMouMgMZ5Dj3L17vBgkg
q/hF0JWFvoJLwwQrh7s2BaA6PtONSUnvT52Pq9GLNTuF08+zbOgla3QM0NHzk3sK
b1LXDLd5EpfNt7SMSI7L2Lde2jyjMZ32znw+gPUpHx7QRaeD0U18aS1XD6chPf3O
QWMxOWFGNjXkEh65SOI9v9Nafw8+JF04/qcciCm8hFT/R/706b0jmW8SyPeUgt0J
PZLizyRJoK52mVifrcJoS5JRNqs5w9Rn9RB24gSa+mZ8vaqRKWQwM/RZ2H7TZAVl
di5d5jeIVtN7B6N+m9rFcuTheiwtYuio4ddTCSiVsPZNIcu8shhOLxEKwi1WUxxP
d+ts4+CloAEzEpjN89hFk4jjFh+YzigSxX8OIS4tD8cY1iG/MzDJBEdy8SzJ5LG7
9fx9zplzGkZs5wfDCaFCezqbVjxmj61mjY5wkJVaIB/3ek8KPHU+F0dgnaQdx+fY
4S1480ek1aN7SuLK2LIkMxf64+jpZtIxVNcDqFnml0zo9ZICtBuiUyHE05foHa+u
kq78bsp9O68k82ODPGV0YODQd5QOFsuWR1B06hHUNkuiB3nkORhM22UMaJ3m47cZ
ur990U/tRU0WPeAkQQ3g9LhRCLGaJcSUvf/qmvYcRluqYkmCAaVjrHqvWpkIGbJ+
xRkRRE/3br2S24occgTmnQLKOh3Jbofjxv5xmzAUz6xb2jg5bcfEyq9dwvx92uMx
+PGyQ6pGpK4Zrgvp0Hwb48FU6/K/d0JR9z3grgOPv4NykdqeZMNUO+3iIuIeB36N
`protect END_PROTECTED
