`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lB9Y7gWKfbcfcShyukQjpCBsyK5d9BFyeJgjjvY8KID2iyntxuGT4P1vkZJDNvs8
Gd2lxX8BrFFqGqkw6ZhHP3z9WmMz36bs97BkaHLoIxXwedMEhJjqmtx8ityVY4hL
F/RtfcAI8vH2ZBg288+1ZEwArgp5Mioy2t6cgKWSO5kqVxa9MlIwo7xgei3D1PY3
UvR5i6j1AJESc+Nao7kpV22OSeHwIczmET0WUvu237mMJtaRzdfBWV/JPZdgzNX+
PEh56u/7SZ2ct+G7Qkngn2LGnbSNGlhKTYeF6JT5aoG6EZK21Dr1nBJYCjJ5/owm
s3dtxZwRPGLDaniWFibkQvu5vpXuRPONvIIcCxc9bEXDMizbl4vInthx6cEfQYuV
21L13LCZKk2ncQhWS2KF3/AECnH0hC/l0y+yn778Jmc=
`protect END_PROTECTED
