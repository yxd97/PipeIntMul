`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uOuuYNZmeM5vg3k7OY/PURR0G5d82yE/T18Tt6l++s9Sm718tzw5Wm0Qs1mpykny
gk2HJcbMN/iKJ46ImNtVIwqigoxkS6hgyHna7PuLQzz6Fl8oGExK+gaN7Z81W6wm
svDsf8j3iQxC8N0vT5TbAH8ycXnJrEfKGA/H//xTcNhL5eT/3kIYGtefBxYmx8DV
vA/uvjCj3f3PNK9xn6UIQgNVoFdSOiRhgEQsGvHMZaHRYyz4lI8/+44uPfg4x6FG
+LgDEo9giM+IFMsEo3ijOM/0w8GFAr7nc1j2cSTE11Ng/bOICnLtxLAwKIJG8OjI
VEKU5NMsS7qYel4LmRiyoanzvB34MOsctLgcFt3hDRUZlJmBMpZd/4PG6eTUjQpd
fpxc/kr9DB7G9RM/yIF0y2FOVzOlFZ0u1XloFgyfO6TvJxvywAeELb/kJYZb/k80
L0GhNhi5xQ+HJZZ39VZTnNkLNcYQdSiflDsTfFvPdq6bllhKiNnKZr876kx9uGpA
bZzL7A7DMB3miZb9uL0wqwi/aXY0/2ciHDdTGpaU0DcTwLNi4jTp8csrmcHsNqi/
AK1HHU73H1owNEY9BzcFjmrffJkr2ESlwDgHRccaGKocMabArs9mu3MmHkfMeGAK
lbtLMZYUMSo6TKXMKPhWt+qvxKfhgNc5S2AJ13YgvTz3SHchY0Zo4C0iAOoRnRP/
sdk5dzN4gJffkOhDOmP9Lb8Stlash5LhjF6LDBP2XwpW4YmOr1JL4OnahqrXoFUX
YkxFgPm5aSYJTAlFtOUF3QjLtCWq9Q0cqf9/1pJ3vBv+lcklspyMHfrcjTjNw5I3
pdWqQlrYc/0Okpytie2TGp/WdMDGOK30r4lZbBl5957egLC5VNuAtcXRcDT6fGJV
QupvHxqL8JggMWyXC6m2AzATeban1KbeqTspXAVhjv1U253Jl6VbZ4vZlc/MxZLW
TEkG4FZkP0ADsg2VST1fdX5aR4r2qPBdwig3UjY5cDCR4O9WEaUVlKpUl6oA2FOd
VzY8d0Nh2mzoN9BLXeukaJdWOw/aps2/BbtHqrYlb3T0FieXFUbXoS/Rd2L9GDZ4
aY+iSMVbBEZogJpYJMP8PPDNztZmziQffNKqMpi41iNIliIFmPZM6aOuI0/XKevA
7tUMWdCqIo5zFadQ9tvRmxfgQ5TjPSUMs9Fma7LMGMtjPGIwih3W4gBXXu7aeuCl
Z3ipNj5YJtedVhUZCXkfWEWNM05FhiVd/ApCLAtoRZUFGFMaqoXonnfs1ChnR/4s
`protect END_PROTECTED
