`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eS/fgp/iWvCut6qsi6bhG/kg4axOsrs/TQ8998Sd4F8nZilo3LchnLTl+8dwoxRC
/MWncpPv9pmjqRSr3547dtWVKYawPP9TdXcVWu2xNW1gZ5Rk+oohV7N33avF9iH2
YDmJmTt3pt5GxHQX3OuK7BYzbAl5WVJf6e8+ECB7sYvl8S7F2UTkbOsnW3QMMPhx
u3X9qnwBuynp2DS6u2uBQ8Ci8oLQdxvwDKLEzcU98sSWabkcK/1sPn5j0UNB2Esv
hcWJCfFz85cCwjeDKFDdCLArx9vEC4wVgyxMljVAOE9swRaspqBzIae2QX+nGQUv
9BT77WuFdoE4nn/R5gbPQy8mH+SH4N7xqhvIW9moiRy0MFeR0knQF5lGWb8+zYbH
G8g8XmjgcyevzKr8l7wW2Uzh5epSGtWfIi3kSvAuWabc8e4DNne2nIIguMzqpSUU
2Kti2uHbj3NPmkyxnFM+qKBNhYSer1dZDjQlEmk3Yzdt8E7QBaL7TxMh/w4eNTb3
pJcBMVFFHiHBMwjqOV1dPaadZzbEIrtpcsgvHAAWzq/w+6uUv8bD6OeXmnRScY7b
s1SA5cK1Mfa+AJY+K3mroctKZDdepfLcLJWgONWwthGwUYTE3tvQJcTFrc7mPHXR
pz9Oxqnt9FqhwBVPr4ofSwpmH5QcIOykNHy/Q8LytVMBniJN6A6aA114jHabvZxa
4lNbcpzT/rDOaxHGhQeckInx55804tZxIPPsvDIXQHDJpvz4aheC8BXInpIBSI/h
S+kyb+FKk8MJIWF1TwXnvsEelrj7sOqHw8KcQj8OMSwD0ccD0AIbAzA7R2xLIZBn
UdZx1lZQ4nejtskzmNbJMO/69P8BM+v4OgP36Z83utTmZf1gbCd0ATsig0PgDeXF
7KFMjCWe7y1qf16AjKb+xKoKUt3j1fSoMSJfwB8L0HlNgnilBmccgVMKDswCMPJQ
O5+Bo9W99nz5lMVZfRjxJjvuljmBJsBPTqm2wk7uxE/Urgj6o42ubd3jXlABI39l
u4aBGBJbYGTN+Dh2rOixAQerBLkLm8KWFmBB1zYHrjyI82GQFoSasMavj6KlvnIZ
oWwW4nz+NfrSQnHeaOFtjwVyGrBbl/jWNNbN3tpDopwRr1T8IKCPuPH42vHM/oas
zWJKVXHro9TC6NkRBhJ0Hgl5iAoa9MJlj+q9naJeQf7hwzlBi8qpquJFPpxVP8BE
Lq38FIC5qon7JOj10jrbhP9gKRJeikBJ2i3tbNpZowl3K3sphTpdH+1XYrtSd6aT
gZKHWC+2a6t0nxv2Ttw2DYPUZvzLWUxaLUMhh8FirsGT4kSfWOoQ1ww/WJ+w5WZX
Con12fxjcjjB+Lne5lawb5114fKkeJDbV2wliFu4+DebPjhS6zmH6GDQ6l/WBkOS
H6ZkVCTWS7yaV9ZQylujwQ==
`protect END_PROTECTED
