`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qSqsKrxrM08Czyab+9QwvZpH6gupmr6KegSBy/dlogZLLn06vMpPyayE5iBz3B9J
ZOdIs6Qb+/5qzPTSom0joSx0BoCi2UPIshEvsP+ISTlrRFrQUrJ7Z9L2FifZFdk+
Ai7bkOQFixv36Wf9TqY5VeCY+0fr9cNUegc8TY2cqq/ctLpdWlbex8OAMrEXhL9n
w93a1KI+bAeIGGqOCTZN7LwwNIVpSPIynPohsXg+h3VDwAWmzvV/LsoHe5JjS2c0
EdQ8CGz4OuNX365q5Ksz3y/a9Z3/sSTrb9qARjZ0jI/NmEMkgvroeU39onN+yte5
fa2hFZWy9KVyKVTfG8tdm0GSH/PiojDPE9iOrX2qN39j20EkZsd/NAe5a9t94gKH
uY9El8NPbvjY67P9TWrOh1QVVfmBD447KqqkXkGW1ucxp2oY4MFKM/OceE6ASHWX
zj0ZuHZRqtoF3zdFdInOnV5izMMxFUQeTUMHRbZo0BbPWqFk+7Ac2d7GCdJmwFUB
mi4agGih9mmdenhlKYdcMKenOdwQLf2LYgXVsh/UYw8XI0ZZg55YJg71VX5JQ0Bc
HeKGDF8jA5VRUns4LPKFrD4L+2ZYOO+kWpFuTpF0+rHlF83yUIJ12Q7933Vz3OYn
sbOISZ5fa6fh+27HwpiJiPkX4WqT1D8pgLXeji+OgDhDdkxCq1EeVlYKldDd7p1E
pNYNF40r6tqCNKTF9KJDktQl0P7Yt+SR44CTjDOtdgny3om9wsnee2GuuRkyITwN
+W8ZMszBX2jzrl3qy3Rsg5/3MpJjsVzyJCbR49X/qdD11lLFQtLG1FCqbYk21dRw
IoFT5iwFoP8mILQBo+AJpOT1cMDlEpmbHpUyCp4Qswpw4i+USy19lqOZQewq/csg
IIRb+DG1pB9xxX+2jjUOeF9YAOXQsTQmRQrwnuA6MAOjgQZXwy/mljTsf0WMvtWs
PFk5DXKnlWmN1UKvem0MQDWLQuJPijv+u+wmhKe5b9/s9s9TCOouCFp+rsGfBXfO
Vn+KAJsdJrwW8lBV4Y6Rom4DXgWpIj1azfehBe6/ApH7UUcBFdG7QLRDAb0yjEn5
iAdwiEtS0xMbzXV2P4MKGJoOBObMgu7rxX6UxO8a0GtZawUinPK88+laDSaUdYaJ
tsijTOvJDCsoCcz2ZJdHdsLX0y9mNKloGfqocHQpdqIdSM1k/g6K5R8G2ioIg2XK
vOgMjYU74BhPn1sdOp6EUENA3amafrZ6YnE3j51ul1WufqRwcdmmhI2FX2RRRE6S
sDmumzDEnOlVx6J5JbLTWPOLoKPWIOrZkV+ln4cGI+yfYbyTYUWM8Y1QIIGquc8z
CP+ukfBMvRtKBLmxhWrirYsFwJ6G0eTaVPM7zUQhFrFCqh4RlBg5TMk3fqGYBGTx
gSiCnkIYHvzYdHI+U4pXGwP8unHkYopsXl8mM4+g2U9DIcNy9euLZTxZE98ouqJB
+FGOqQkYlg9DhMpiky7gpOeFsawT02LTTqmBA1vDscoo+XX0HcwKv96O+w+ROiCl
vTJQvh52zTh1HQRL8aFo98ayw7VNjWpi+hJqEusJAFDTvLa0zgwh7lO6P7zeZgVT
/Yvk8kMapvaipZB/VzYRY8okvlCIcW59hjf18+E6omBQBT9MDCV11mq4rO766i2O
hfrSJXwEgROdFR8Yhvl88AqW6qhmscv3BJL+LwxuZ3EwCzFkKn0rSF9MJAQHWrow
5UGzoIhEm7wRxghUbILPbqC+UIDvE4YYMuZ9YRNXkII7S2To3bxy0wgN21Lg/wvi
e+uw5cMCpJo3dW/woMz17UvEz9c95OGGwEBFFOH++4KPgSBagberaNRHPuTaQLuD
JKdBIXagHzFLMQYtk2aeiiG3J/YwT4HZmlDuRKmn4DD1iYIQnFNGqzfavJ7X/g1i
M7V03Wx9lVmg1+itt6TmxEqHyPVQiV8DStH2A7wDJzxPq/McbRbqxaHfM31wbk1L
VI1iM+hjpzuD9oeA+/EyTjwIA+CpERNBulq3q3Pdfvw8SXYPkEnfbCp6yB+69Xcz
3m/v6UMjmS3SP451V/BVkrCgG9GqX5/ryiWcI2N4ED8ltyN0+Ai1zOBBwDKcAALL
cqSm4yVJe5djU2oK2EopXvTHlvDCv1DT97nQOAcva5swdRoMrRzm54Sgnd5cjjQO
P0nXk8mHj61WuEG7Yo0MWxCT3n1up+xglPoOPVIQ+HtYCpje1HDEzcQYqcR5trtA
v0mLzeqvd0ZTCfgYqifoq2k9hgq9lhQEPkk8LD2T03ir3HOxVAArtCcC8GnsQrYR
vCVaOuTgZs3hoy/BjV8YVDBh6i21wl7zNW0NU2eh+zNwOkScP/DgedTWNxAuLgEn
VdnnK59jMAIChQqRBb0XLEQYdwOAgQUGw3GU3EKXyhn9OzPAFdlEn79SJtl/cgzL
JNmGPydaNZxyBks90w1MOopL93A4vAtPoliRw3JyNOgM4JpuElWMSjNupUOoMyH7
iujHrayIic0cAEEoc3APiKNrmfQmDqSzlGOXAfZwJnhknzWA3f23ogKxGylxJtql
FJIlFK470Y7dZKsBNAevvnwUM47uaxZkT9Naphfq3vwqTje0CC1lsgylcGnOITDz
qHqds41EQ6LPrZhg+ms5dmc7f8AndiV3LQD0Ymyab95tqOsMyytPhVLiqEFu+7nC
8zjpl1xET+smfUS8mmKbm8aSHz9Rk1OCF7zxWjxSvHwVa4DvOazAyeOlGd9dTpru
9qGh7RPvwT9wkT/6wP7KTeX8PU3Iz0s+eIQKQk8h8YKxQY2/yHueM6skYhCvf+G9
JN2Y04gy2jx4VhUxy/abU7ymTFjJKmu67VNX6i/WXBY6b/xBQt7ln49giKh+hOt+
WoeNkehbWGnbiY6o6Po1dxvE0HbBEnTMQQYpdbFjjAJLz3jh5wW7ix+nLMLCCCrC
hRgA5cWDGXYdAR34VTTocYnqUtbSSpxmO991xW9CMhSkK47nvy8piU0IVTU9MGLK
zxcW4eWs9cLaWLtDECOIJeWz7VFE3n5kDuzNH3YMv1cY7i3enG/rR8o4Lq0D1puD
Mlzj6VRvB5Cs6pxM8/OYkxEJhuQWeGOc3dK4n0E7WorcY10fUDB3fxnzfhFO4Yd+
0e4img9g22a2sym94JD6p1ctqHKHgBnwWyPLYuTiptzCqBwSMqIEr6HjaUlZEMcO
kdgajEUYPSFlxJW/ZLb8OuvvTp7lZ5AN0EN80CjgYj6qIQR+FoJ6Y6E7y9/xofP4
q84cIsh8KcZPEnvpmdWFrk1lTYhp/XsuHJXvjEMwdQTBdryOYfxTSza08kQYZoXe
yO1mA0RAY0GZ8RHUoMy6XOt4+uNyhwUgmRS4XxWAgXmONvncRjjBTylWRVX8o8YJ
ipmoRP2SVcMvAdaDFBrW7OguoumBKEhYa5LYSbYb+PQuzebpGKWIGBRAPmdO+sJi
xs1M17iaUEPI592nHR6mInGzcwZHExnUYQnqCcLEBhPhfCIAUELTZNLrHpHjX1JZ
MQWjG4TlBpCUWgM9Ar8s5uolQpI+9jXyvV8yijeeRL1y/ohQYqYag5U/gSMqA+95
KYHR006zUP3jyWxrG5HtP7U8Fo7h2VxymNb4Rbp3u6Q0KS79eV71ncr4mfbORJeE
dUYE5XsQDjLyKraEusDu8vsD7XCNhlIUzjYaHEX1hogxlbpShSn5EA72SrxgbYUU
z4+hBpsEwRfNNqNsfwYsSARFAS5BShSsXE0hQCV4iNWlYh6iPWsrYCMlhnyCbOmz
kKstbQLkvRMLc48kmkyUP400JIrUi7r+4IfqKw2Q1ukLwMAg+VelLOtLH+f2O+et
y2IgkFyZi3OLLoDSr3D7LnbjnNQqH5xsnHh7+JLoRM7+x2/8Rk8XKDJwvM2rr+LZ
7bqqfm86G2LFwCcnbgeOzA4CNHAFno0i3eKSSRkCDhy9O48aHV72c5p3A8VnZGzs
1Ia2wRJhzgoEGWnXpsmTvVhnMhCqNnXqiBYwmfO0pB3AvKohukajVQuazOgNWi3Y
wh1rXd7KVbj7E1cfTp6269dBm85WdIDAic5hCp0VVwD2kwRx+7pwlNpScRr+qGQD
fqai+JDguhSqHEchdUmZ+yj6dl45WMjdnZeLnlGUcjyKwfOGtJIwB58M/ZqVyoq7
23SgiYKyUwhaDSKXoQwEzV6K75ISuQ/61y31X3Hu9/sPThs/s1EvVEDQo+8DQ4iC
axcREnEilEOQ/RUKaWcL8NvcMyC47HyZ492fy31vNIDf8bQbknrRPLP4wHU18qLm
HYhMsshKM6pg7K2UIso9HstlZU1u2wcvQ8LWK7sXjS0sRcipuMgXP0DwYzbZYpHs
ot4gzuk8hZFBcNXT58O+iWqMlUg8mQkWS9QTgOJjcaEL9gHeTo6+PqvUbAhIpW5h
NQ80yz6daQIn5EPi3B2s1OQQJKQ2YmQ88T8FCwGq39ygk6onYj/jvMoBM2kXR8sT
T3uVyvgLK+PaS04fuf/vzHNDFqVUSl484fpM/1gCUf9MAhMiNlrX2bio/4fzpXcf
v53Or+lXp9INM5OB/OpY83H4MLP6g0u7ZSiWJ4ZGwF0AUr6DK8x+pGSFc5YLAx+r
DEpCqTs0hOwYyC9ZuQ35C/yygd1o0jPUNB+SYmHWJjepVU7mDpTL3eykPsf7MXUe
PXO5Lqn4tnai8/nE5ov1cng8ZgtnqdCDxzi3s/FXjn76xnHpPBeEKgtXW2sNqZwu
gkJS9X6eWgtlAkEF3diLe/TOAwsxgR2pVT+is3cv+aqqtrn0DWSHV6TFYFLzFZ9e
FkcmHRo3zuvi0luPd3McyA==
`protect END_PROTECTED
