`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aYcx6e/qx68D9WEt1pr18aAqzNlBNF2WM6/qiot+whAYAzsWYXe3qSEpJTdZtt73
Yzj2arMwbr3oNIW56xyJoKadd2Ucjc4KO2rBE1tO5Ru4O9fnrpsOW2WPmx5+w/ua
O88M46gv5Fi8kTkYYZL1A3nhD+jN2A8eFzR+gOiOt9RXFlZ9rbuKyIUHz411SJz2
y6soV5xRuLxy3P2DM1jO4bEsu9o71V0AdaqlAncxHGDiuB1o7YUwsJef0v+a9jsN
x1Yk6ykQANCWMCcaFscOfgKM/pDlv2JsJ4sOosnaXiY9kj7KUh/USUl9gI71MMKb
`protect END_PROTECTED
