`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MvLGzZK0fTEUED6dYbKCKyKjrc3JCKi2QiUAcARbNOy245eDLdh5ucSMJU+IDPM1
06kvFhnHVTUgAdVxyYG+Bk8iZGgKQveZRs3MnVTUXC6pxC8Vqb4pn+9NEIWiSOXJ
BaD4GMjNWBFha1beRHHTFZRQF5OMB/lWblsaXWT/sRGEP8i+htuSqGGbq6s7Q0ix
9jAZmbVE28WLwtS/naieutmLe7of2r5nTzcf+27rM03EhkiuUrcfXME1tn3+Co52
U06IE8t3n1mlSY4yYORZokLwvVzhUrL9o4AA7UFJdbDdwqrDhHtg/adiilKrlXKF
DWQPKVN4y1/Bfx1/EdfnmuS28LRc6QIrDvQTObHX7HM612aBG6gXyBwWGW+us9QD
bEeKTxPXkAGKVC9LczRVDRB8OnK6h0/lo4YcRibEfzs+9CvSLGiXtiFE1mCbqEHO
0i9CAqi+bpVTCvZUz6QLBmr4/v+uFX6A6sLTk7tvfxeymZDPfyzyABOo3Qmezn7R
HUR6C0X08H48fCty4/486j5qoY4PyhQHoxuMGoVigOgX4vjXdHdn8CzI5XSLjPpm
P0yWV3fCWXlRxwTP4UBj+T2PGYSP34+OsStewI1vuGSucBB9P2TEyfR+Znf0kS+b
GSuoDcePrKRvikPMR60ZSTXTDiDWORAjayH7jWNvF7zuKVHOh+Dbm6VTvzoxRtrW
u2ynOZrlPQ7B71Yx07fl7oeaExMl9Iisqwt1y3IruFTOrD+Dt9G3oIMHhWKsfMB0
QTGxw0zGm1uoo5fBOb5zMpI2xNdyEvuZIebqYErmfFj5MEQp22DcNyfnSpqAclDu
62UeGwPLEaj/Q5fMLHauSDuEZK3MY7Ws00zvIJRUQkyruns/oKEh4ACxVCXu2PnG
NSrNcqZ0FZ7OJ1SrRiHdlCv1R794qpFOy5jO918nEEhUhMeAlIFGAGKhj0SUvXQI
wrpnqFyVVjgMvem5yVt2TwGm8bythO/TrfmMkhNznvAoGWMyhExEijo6mEWteJqy
LgD4zt3G7F1c07K5vfAnWiAxgCJQeFkdsj5Ra2nfSU6qTwJxI6tiSTqzew1QPfE6
OmqcqjlSt9pv8dX8829Bm0VKuG0TjQ8jKtyRhCQA4Dtl5vjDxlkaSTO3Oqan6v5p
B3ffHeQ94OjAPyPd+4Uw4A==
`protect END_PROTECTED
