`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MzIdgJuyRRGR2yKzNO3sAYBsBRycP2dO0EXLS8IWTsRjTmQb3jHXcnTrajhnyEHr
bFvGJk1HfKjwp+ubnVnRlEnc4ar0+Khtdf8rkVZN2DGvuuyZpd+11RjOooc30p55
wCTwwX200tn3ouWcvsnRgmfF1MKmtsKDLiEVUhtPjdrSEsMF6jh6sW2zNEOHeJDp
qi/HXfAagfG5gF0MwbiKdzrBPJFsC1wAh6TNW0K/AZ+mzY1wYnibeo1i+PEJXkx2
0RZ4dmwreqlzELPz4337F6j1bddlkoiBoq2jVaffWyVEJvoLSMYUApeliG26sVqf
D1KWacu0KV2HUm0jRNWGYnPC6hADv3M5G8mIuwTwpuzeZE00fFaShAl2axZKTm3S
OPTp7EA8D3fzvoq6OEXKB5DdArB9i6y5D1IJL3npqjBc8yS+Ja+VyeJUyA0ve9LN
SQvI47azESGt3VWX3YYdMw==
`protect END_PROTECTED
