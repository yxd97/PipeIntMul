`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uqYgQ5tWucgdV9z5Bk6wmrkdqHfv1LkxWiyu05OlaON8HxvB4d8i8UhPtVrc+WN5
R3QXQSmLNqF0NfNCO8iiQ01t3MLb3wVhUuXvo98hVikUydzTMO3zzKDrR2p+HiZU
uxbGwRHajuIIJW67Smh8GHwN8VVG66Prmu+3gXxNNgu15ZwXeOQmmmIrHgqCLPmd
w7MG9jP8auCTJIz6s/ARUIi2N3VLTuPxHRjAglPItQj0H+Vp2+Jw5VBhjOKRvMjA
Q0uV6lYBt/FSt6hiFFM7RAyDZWNmYLARPjEUu0zMsZFc+nkbr4E49KWMX6MVtoxd
CZD+blFezgMu4Wl4q+w7XiPX/N4IYwZHeUUd/DFdmOAKiS9kZrWGBrVBHDb3Uyim
fwDlhnTEAkgIchWI+qICU1VHgl10xuxhm0UMQwz/m/RWLobmxH3DA3LfkVCHpUst
`protect END_PROTECTED
