`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cwUTJEsPrz2jdbUsk5b91auRrKbqdWvOICS6Owjg0IjYxqtC8mKgcRieJWp926J
bImzzmvo5nXX5gX+Zk7518Xu6N67GfHZwW9U8YBTOGiTeV/GgrXBbg7v5u+0hZ36
WvSx/SvRQX/zoqglS8kYRglppw4izu71a6XAiaK3b5SpPyHS3hq9QtDQ2JdQBGOH
Mc8WcEpXK9mFCeJ5fvKwK42axx9gDJDJZDy09GcfXA0y45PlUw918d/qbg4KCbcV
fWvyau87CWwsauA7++lkgtYxskehWWiFEyhxCObjyHGYQKJkg8+yR5FuskZh0NgM
4XCdciHN6w6kvfhhjfXONqHyzqnJJQ8edldupLR7UnpDS5rgjqDsso3h0Oqn0CrL
tqSX53VNUpeoYf4yvdTk1wb4ONL6MsUOz922gapGwt4=
`protect END_PROTECTED
