`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IBsFQzgTx0zdeFKbugAIdp8If0DTsqT8tcKDrfxTedRHOtXGMyGHgVvMBm4xfZoc
RzgfCQfJFUN++rWVMviYtXg61XwU7kBBj7cvRyR1BhYwN88G2w4+U8VYQ0Nm3CZI
C7E7zjyleSoCKBcQ90TMkCnBN3V3jjRh2taajZ82cdR77Iws8Rz8FhNspm2JzsOY
+JcUTxEOuX4cze6qoiL1CkIclEg9t6aeNgR3MK/8fLaSV9qVSsTj8XB//ztBjBVx
XL6BqjtN9oui4mymZOCh2Pk7gv3KyVVuFQXMUOmg19lFf0u85qFK1zEtfKhDv5on
Dia8rQWgoD1Svaz8vN7FUwiNNduxmXoeiZBFlxVTg116zNjoxtRgw2DakCgfjzxt
mOV2NeNw7a1dAW3fhLcYOQmKgpLa5ANRCF9IhRo+/Y1+SpqX9SGSDQ8Ht32ybZSv
m6+kjppU5gfRtOJ/PJrq/NI8xRSup0UdxT/bo3LWwbf4lTXAhz2DU8q7IoGnRYxc
+Ml/59UFzq+6EM87i/u9+3Z5f+S1k8gwMbBPTn6lwDk=
`protect END_PROTECTED
