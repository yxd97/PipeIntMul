`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FpNE4jZ/esfbJs1z4XYl0zyYZ9neKjC3M9glskXkpbZre5KPD2bfYqZZBz4aSfVi
kiNcr9bVG42Z9AS1hdM45MSnBasMSE4lH8MM/bXibSnDHhyDwery0JxQpt4HSxsK
TcUSP8IEnopzN5P0if30x4toj3y0/lNSbbtRBt4845akQxdqelmcqF9rgq3sdh8Y
01ATGaU86NczFuwo/Ka/mhAo9t5RcUPBWlJ8rOkrHZ4+myX3emszgfX+RTXJIBGq
BFlLE4R5RAprHmkyHHu4La9sP7JjrLdnYYcjkWC5xSKpbF5qHjKto3pgAJuSfE3/
rAzJUWuzClRJlq/RwYuqFXHdUOZ2nl9tvCkVSt1q5h8EgPvUx02VxH8BoTJQu6r4
wCNqx9lbBh8fAULdPrJFgFbjGR4UTsbvmWkmk5jWCOTwm29wlPEy9Ei837Ut9Ysg
2mHOPb+J8zigSGKotZ4CMZ4+xHwkSFV/tg4yZm2Bbzsqff+p1/flPtZ48fbcfUew
Vp021aH8Jjzq5Al/PjsTFL7GUAi02L2/FdoWjhuui7wSZzWtzjCAsqz7HQaLi3LF
uPsI5ygbwHziGJSR+M7oLjkUkAbaMLlJSQa77Oj0TfV59MrEn36AnAxFBjIW9r4w
WjKsqPRBQREfNH/OSeMsl+nlt0IoR0eSp0euPf7Dv0HUgABYkf5ngLVah7UDvC78
eeV4f2BupDYJ08M08tB8PmRXB5/M6Fk6zv9G3jsrn5g7zmO9yhg3dl0Up7f4UJ6t
kdIASRRTjEutBKGALfn3ojGasxGMpy229lFI3Pm4ikKvau5y9R8Ok2TDKu9T162V
b0Eh7wjuTvM4I8nEiOBMCrEm9W5JYndj8rJ/1UQiFNL5n26NDVEXEQLDuXWMhEOl
NhopLGlhNwMI+giMZoFX3cun7vqcoUsPB/48VebSRO2ui7Kn/zFG9P/kcvcNDm4T
`protect END_PROTECTED
