`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UCsQRJsFmWsAQ06Hyk6LHMwFYxLBW9fdyXWBY+PBtM0fX9gX2vl6Zn/yHNBkTOz8
+IJaJSgJQ7fsZxSBWNujXWa2tKPTQtBfOsHut+fG0LH1guIiQE/Ox/8jxqT6Lbvc
zJn7DJ9urTUpJB1bGXN9BEWke8KzFIGoX38FxJxDhAsw9w+o8OoIH+zm84cnfIUL
KWtTaEsk5MOHP8JSLvAVc24uHtJWZvOAXbfOrkKlZYs0QYm0ZTlJePPsi5yQ0C6I
LYVugY+e7Ui288GKtfjTCZGTap8Li/tHKczcF34+0YKjVkDD6mkh2xI19k1E52D2
reCyuov0XwIu1T1dnyC0qwCt00RtxJcrz+FuF+6QcImibhqnkWdJY4Aka1Pn5+Aq
tqXmIvFodfGJoUIQNuSsRcYnLWVjVjI9rxU1eXbxubgT789EIJvaB50QMGyUY65H
43eP7KsI77Jnw45P8vYLYZpMbRS+1B87Z+k80kQ0yxk0Rd8B+TwSb2aedq61Kge9
9EhKYP2Qq1bicdFp1wx0/MotIQ0JfsGr1IjgUOUNEd/KeCHP9yE73IEvRa22Uu0/
SJ0ZkLFu41fhwx/OSlLQHkD1iirG/8MxIjHDp+zVqMtOLPIOX2vyLl9M19rMqGDx
9s7qcxPTDRxJ8D9LjO4Do6N4ZOIOiwBsNPaqQh5PzvS73Wc2jA2EXDmcd4j7iiR0
QUfRtn8loYivRVawiaSTSCevXRkodKizw8s8FyKER7DSnjYQ/Dj66lFsiGiMzw0L
kvzGIIq9ceYs7vT8eF/f6psBZPC/MW4jYhAhgCSwG9WmgMKhq9TyYjxNGMNtXLD5
ZYOROAE6MbvWNpo/tdIQCPHU2/T4z8QWO4Hp6bAdO+VyPBlzOOJko9UxzMl7Yw1v
l+p9DtpReNXN5xrYnyjP2Vcs8aZDligmo3gEFbGsKnQ7A0lirkWzOFt7+LkOldZE
BV5dcPc6Ni54WJ2d7z5GjySbNmERPTICrv+OMWOeGPcHVIZLqGB2GlrnTQx+NADk
62gPOTRMWT9oIipLoZXtjWSxCbNi1fu/qtcaXqjNAZiTQT8qnvzumMTWZL+OGCyR
nqukxvnu2fnKm7531mnvGzXCRBmOK/AykUGDz53q5LCsyzGgAr/hEeAtOq00HGN/
V24WHK7ekyMPG8QglgcapqaIarwW+d4Uqj3NYIdalUPLtb4URMUfOhaK8hTMI5JZ
Hu5Fqp8DS8XwXVgSzM9XQp7ldR2+HAyiyZsQ4iL7pm16K+bGDixqED0rB32oLXK9
YM/OEZTNNYsPH4cN2HVb090E+PscaokJfbUXi0AgVFR3Jwfqz7E/PdoGxxZuvTp7
6qOvHWNrmBI7OPq/H4kWTDhbYwd3y+ZN04gqjTsWGXisBFUQ8fILWwOVipL797mR
RY35lJsBmHmdTErrLsWDEzImm2sy9RLh0cLF028qTNAonDuWowS1RTSezlxIsQ0q
GOUghg0P+vzs3R5SVjco0OYka7lUJEYwVzbLZOaCucBkq5t6ZwUssYYhdWAA4Nxf
xXTZbLncfP2LurslKOYaltQaC8mBP4LaxHNSA6CcusmQJ89c03cGtSQrqlFsBCQ8
/AwUGbe1BSFnkdcA+ZJjme5crHS1+OJCyqN1UihtPzwR4i6tzT3MA4GiwgrX8erI
pKEmNIkQmoAI5O9EAZl2bNIQhIxFPgkl5Bor5TDIDmCovMdAHgPG1v9a46LBnVOi
QnV8gWGEkyMwAme8SadpR528DVJweQwzyH5eS3wqkUCQeGmtdR6WGBZ495wTTAVw
`protect END_PROTECTED
