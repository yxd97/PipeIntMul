`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RqpR960i9fCxE8vm68EZ9EOMcWX42fqN0eGW1JOpMARdV4UDSV3kiVE+SFLoGRNJ
fdHEQHQlNJsk41C2o8Ha8DNeHFGuLrPqnNorV7PRIQgaAQ8IB8qXx5OCKZs/E54/
Y6lZjN1KbtFCP+NTc9USHENQxQZp8fu24VQDcO8d/dooGWgWysyhGCGZmQM8MK26
xlMfye/ut2/UhWGvLVzaJw12Rxk4+g7+o/U7lmvxbY/oxNTnQEvAix+fwY3DMcD9
JD9IvvHVV8Vt2WSzkF2/FuEs6t39wBSNZb+GcWBqC0s5KW8cH+WMFIyaB7TGB0kG
Ab/YXMYndWGqVgNPisAqB3Wv/Trb/4Hss1klMSwRefIefVj4oZU9xUCKMq39Lq5b
WMe1qz74uc9xVxQGBYBJdMHrY/O60FVxKqBcQ76G3ndh5WFEy4RRHbIvESQSu8Je
kSkX1h2TFQErJVNIAvjvXvN/BS2ILqEhhIjwLPTcOlDrhMqY4B6JDH55gfLkG1pv
uBRdjNw8MLATVhzRtY3gpo4qfcYTp2nKmBL1XPiVhJ4TmCijUoRxmIEUTsHqihX0
H0HoyDrxrtAC+rCgyaszGkhdCUylrLCqm/D76S3LXIOe/VsRIAZOAC1DEqWNRpNI
yM6foICRem9Em+Jj6KagTH2T4i8L1rAbVTJz5x3MZvDyoFvmBhHYrKBoCzcsL5H8
rJMkOdUKDH5vGDJIJnA4IvA4AKRp2tbDPZ1mfICtkB/XMQOUypU5TMp3Vu3YVjhH
MqYsg9KrxBVV+gF+CFprALSf/yViz3C05l3djBTLHJk4UYsVI1TVh1JcXFJMR082
X7XUWkyDPHcj0PRX9ikWbXfsF+I0QszMaKt5O8p2kMNbKevyhBIIX6HkqJwRf/Sr
Bj7Lz9IE2qk8SoscFjhv9q/nW9zUMVbF0059siRhdLRr340F3QHSRCKQn8j+sO7K
n0bXPWQoveM83d5QWI6xzZ8J/NA+h2vb1096Ea3r/wqUcubr4UICPh55WDS3k/0H
fWIvoAdiWLK1UcgkOgDnXkHTW3zdPSsHWXGj0cHU9Fv/Qgel/DoxJfSQEjR0kAOu
Re8ldvUJYkHaLSBUMCj9IB35WsmJWGXcG9mJsJHihhBPMuJkPqymLGhSXw+AKKvU
IV1X7gGijgVNLj1PCK+OMoFToDqdhqdxZM4MHwhCN0zJnR/QulIJt59OQ9w30NGq
FTVxVB0ls8N0Y/XjbMaQ5D9qORwhFWETpHJdzTCta/IZPyg1pCTjA4U6XJcoXZwE
23lC/tUZcF45+I542BTqmowsxTSUx7Yezx2z+wf8ptb7ePjTX++Jz/Im+PvU/SB3
Tuez6iuNVmLtnVzJUyrljsZYJIZrkLKSjBMlmiyGP7Hra3zBmNXlSVBflVUG8LBW
oa8p64C3kSgWmcI7E3AFUBntGqmeFqrRCaB2mVPB0MdfrCBuuIJjCwIc+t2wdPMV
7Qn1In/mQFYAfLZSBCBpDl+GGZppUPzGtoWxGOsrvEZB2/tc6Fuah/J1W2Y4qDzb
0zIoSNHoeGYSer6dZBufzucDu6l2mGiVYlnZvpjUTTzLXevTJqq+EJWvixmvOnhd
+ugub47t4rHlfRk3fSg7tWW3vac7ip+sjnnmJ9flzJzbYouWMrnUqi39malymfND
DAqo54H3xHc1OqceO+aL9cBCTh1PtjSicxV4MsAVmNxxUaZ5qU5uslCaBn2E+qIf
Es6vXYmyl1+V4FviIaLU0Xzv+XDxVLNG0iQXSSsguoUbM/Bkr5rR45EsUTFSPiss
veOMl37wFXu4kwFjARB8WIaopDCU1z92Af1WY2+JuSNLMf8sNXuuHb4bOs7HlSq2
UZq5iyX5bR8LdRAQApNUIEk4eosnGdYOBfjq69p7EbgNRzLXbGGKTcqVnIvZowWC
yz6SYr+SGPiZJ8SL12qPv9pvjL/8MYqNHsCuZyr50PG+prjwH1LHZFnj189olrMr
vYjPgK5tOXXbsvEhLiNB4rjzvE9F4YOimDyMW38g1NPa6iiaF5ElhsfWn9317E9k
tTxMzlegr9fMvca+FN+OY6x/xjUlgFF83Ln6YBFAo5mYAviQ9iKLyTFOFL4iBm+E
F2328hl11l0Ks4LSyDC7t33511H3au8HvxqmersEyJQm1fQQ0q0/wgv52WX2gn47
ZRNSjcP3XzYjv8/t8mlUfKqUa91PQ22isedRk/0f2sKe1FWr2TY7tT9QC9KHnoSp
yr/ibBEoZY/JvTbpUarAe23TlMHiYSNeugIC9Cu+MXHmahCW3KCD4Ha7OkbVK4kl
3yflhgc7pOxEnRuBDiHs9yMZm/i2UtBJNu9qPIndQqLaJgtSxawdV+yR2xw9Pzvu
Cr1DwH2qIw5HXoOnXe25yCG0qNOvYzi5AQz/H8gPPK6F3Gox3JuWU4r5LsogbUc3
vhN4yZ4UnEwpW4aKj8Db5siG6eiAn7MqdWiwGNnQdrMHXjrTWoVZTEcRXPEkF4nJ
U/NcczjK3YULweMcGfOAKQDZCyHuxdTUnvD1A0tePYB99ypKepIlrrkJ9pOjgYB4
9rTRcs/qKWobIWIdx0TX7gI6RIT9LgynHbYfE59/8FKhPYDhQIu/ANP5L/2bvHCF
AwdMvtAMQTFY0kK4yX5z7dpdKAUb3G28Zhm6wyWz2ZwQAPn3JPtSeqKw/3CT/OmT
huRdPcsg5aEdAd1YFTnGxfZh5DaX8hDcLVob2mZyV3DE+MHHCrqmTenCna/nGq+w
zpAtAjAQaz08mt2SGxwGJ444a+y0MPAr6FIGPx9/dhAJebqWY/JdY6ZLRzoWLG5e
EKl17o7VIqmgb2F45ne/3RoVjq+hwp4/RsNm0FBgUPvJQFZvNo+UfbLKRyhu8FoZ
h96vpc1JVnWdgccxTWxLEXJkiSTs2n84XYBhz69Efx+Twn9LCfpEqISyrfcUjC/l
GB8rhW1rpyPU/3ur91RVHROX9zEOZ+KgRvnCcBJlMK5ZOF7+NchNjQyGmws/8Av7
kY5Yo3JjCNra2rjqwS+vkZmipW/hhuxq82+v3TbbWXQalMg4QwzEyKFiruLIUo2V
nBy+Z5OQ1Daw9JMNKheOunG9DV6GRmODz5AYGbu0CririgZIpOt943YMvmhpZzpp
9BdoW3KPK/ZI/n7RZVrlRrDRQYnh6oyYgcvd0D6AbrLviraymaGsmOmmNWWxggp9
g6q5Siix1rdF4iTdOSnmpQBlP9lhIes7W6bQx2QV1LaOxXczbQV0jg2cVS2VX/Lq
fK/RUsa0UHvdNrtw1Ajv4hkvbOOIasefDE4Wti34ovyfAKUpjcRgiGS6jZt1aIez
SoIlu93v7Sy3iRqXpgIwOZ0erR1KSV/REeUQhM0PJMfMlv0yKMlYwwxXZP4RJH6U
xJu3pZBiYbAtq4KCcfprydIfx1Q8s2knDzIHiiLErj1cNtCivz7ROVBeWr/9gaiY
R4P8tyxTKoaHvcXDrcD25Q89D39kj718e78jFm8qrMveljr73YX8xUrkozoabB6G
kggcBTZ5In2ydq7MSfCKagYrvh9yjJznEutfKH4KIBu1qPfacQGOSxNyMl8aV/FU
TDF7kUAn0MhF4CUdZ6gqv2JcoLckqZOfUTKyEhbbBnByxb/FUWRc/MsHl0NzKsfu
e+7q95JSPiz9zLLnpgZOVtjZXvz24BMhXWHyClpd9jh+0hdS+iVW7l+DBpSF7KAC
0GwT/9CSa8gXXsSEtP0uKnAbGjsr8ENTSBWy9Co2AqWQexS+3l3+XErruNcFbpIk
uTkj2XV5g6FwQ9jJJnt9Jh8yUidW8HuLvzDV/qW4861n6WrahSsa3n/VSb2poeaa
+po6e1ynG2J+2wCZlwOsRFgNGq8Bc7ll8obx/S6oJ8WOZjNSKc464Bo5AA4tO+N3
IqWafGuJ8ersotourzIJBVjpYMZXv13Mb0Ls9CDGGihBULcnO9+VO4KTjYKReXM1
7HcqIzMtSJaJZbyyCKZgWnV5myubR1OzpfBMC7PYwOIToAA4asH3vC+bqxh9/kUv
nqYygM1F0bEaBCF97oh+ezu3v6fqO4lGUoSlP7kG11wW5j9nPcFxBxsgMdiTUmw7
zDZuKBk/ujGSPEUvW/GfppthaB79ZHLgTDq2m6qyLzl9LQhnpXoV4P3wh1gMHo02
1WYIKjxbM4fb35Sf/FFpvSpYki9eSzUkFM5pfPlhW+lq8r2omm5cMimGhGpcqQcm
ZvsRmTzgutdldyXDFhkpfLYFA+3C4w8f9yyHO0itvtW76DleiFWKPvyg+irp3eTK
UPHNfCIfKW2UoTw+mLbNMt+JBM/TtiQS6bEJb5c6wvuLRcjVer+L/iVX48mzDzrs
2cj6dYGavDlNOtog0QMT7fLGF4EE1kTLMGpWCZl0jpKqgFDfj6g0zXAOc0t/PCmr
h2TzxlghzBFPv6xKaUVdymjHIh866ejIQ5B8DS5STSeA3dG9Rt3ra4JpuWU1l5Bm
c1z2aHUbGaVSg4OBDyY1mJn9r7/bBx8tJvUDQhEOb3a0RVKmJQ1s0YrI9Ol4RvRb
`protect END_PROTECTED
