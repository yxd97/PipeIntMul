`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
deECHWKCNIZ97mpLHavjDLLLaU3+NKuI/5Sq4EJ8JcYTeHCGmj4xxWnAuTf4cxRf
cFnyX8B4V46iHOz9yaIcNT6gm0SMjWtnN5wS/dUCto4xRxM3Sg+uyDTBb9UsjAEf
vsBFcWXE5tzn7KszGauzJdnhtH1euExhVk+8Qlxgqd8gmH2eBM9Hry82y76MsECf
0bQrCdkKs8jB/uvBuhCIuYLq4NhBBYA/sAmS9g9fQOph+y9YOuXQMqTSvMUzQgLh
S0EitRYXZ+a+q883BFW8JZfQ0ThWwOkkRZWrPbpRP7c9+Sk7DemPwQpB+MTClnhq
cI8lkm4aBVbF/ZmpWB7PD6N5BYmyYpysmkwN+2c/tJXzA3OvgJJ/OKA57dkMXLC+
d7QbkM6p/ioazViF5S7gTWSBTm8d9cgWnXOjN0beeh1xwm4XSk17Ru8B5BAcCiwU
`protect END_PROTECTED
