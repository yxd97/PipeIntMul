`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWfeStiVKRk+fA29vjgTak0dez0ZQ74XHAcG/jY6zcfFPB68+UNRbg5Vcxqd5zrY
7LlsSiINVCIPQgmqoEyrdHZqIH7Y4YKPYM8LNoQUQSP/oTcYN4xig26GrUfkR9Zn
ei8nljyaFdWBgYRfbSaQdIA51jc/vROX9gccCO3oZPTrOIqER+2QhH23Q4B3ZXjq
NbBTKBCXz0dm/gzr/1V37gBLI5TRke3GydQa5D2VDpvNi+XYldXVSsUgjra5zD7U
vMxj9fJGgNtiEj0aUlPHPyq2IYimnHcCbw2Aktykbwk+yQTz55pTfGaPfTOx7dKP
G/FDY1mX9qhPxfSS1Qe7RJPDx5dH2Ieel6qeOkHj/msn+1ryM7qHM7uivccpxzio
vPqACHk3lSLhzKqY2gGmyMC2LnnVDefPtTlDhu/OzZJ3FARWEHUfgrpbKbMnwe5E
7NN+e0NfXrmQ8c18jB1ZQlTRNR9G/oAVYaOWHxIHMEScS96PYA7rjbefWIWUpYfw
LuwYPpC4HX0rJIo2Br8fiP/+3msKucMUCbao002iAS4=
`protect END_PROTECTED
