`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s5rcERXJhzWXoxseJBRO4VgAHvf2A7DG608NNInTMIOGk+mItECNq1F3OOQd5Wq2
AgUsLn7EcYcJAgES1j8m0LDnVYGha7Vghtqj9zln6hFeMHHl/HFYmhKLJ7hWIygt
XKCPox0uYYs0rr869PmQZFjyRROWYrfXtQQlNX2M7IYhiDaJLn+OuCH/0QBQqt1N
WsDQ5X/TiHfnU1zDHfUrsQjLwnMrXv0j4DKCXKuURRpJdwVkGs4CYZXCVlX2R5qT
0LgXVgAaK8STeAZnQbKH/98HALFSnMX84detLZ/fsRhmCqyiEP2EJLmsem0AmXAA
WgYpNB14mtqWwICkVyZJkkpbyVfhlqOungHChBlVmOlA4eqUvVRSogs03ppLZ+a1
QHs+2Gx2Dl3GRa32ye1NWU8/u0gjgMY5/H5K5JYcAIVrJzKnGRvQM+d6p45XdS+1
zV1jbahLKLvi8Mq5PB039xX1A3PRiHrESp/klZuHjuIonNsCyPxx7AgwXu8AZhpt
afBd7UYkQFeycFodGHPqYXrZkHyKucOjWkuVTVaQojr4hQ+57hhj4C/oReoMu2lz
qMMyDEIuO2N/DlftZFS1QxZ9nSfo2m0SujHpJoj//Gj4bUx8yUHY8Te0f9wmZrkX
SZa02ptvPU0kSs7pOwC4TmR2paVD2UiJ5V0k2vtOH4o=
`protect END_PROTECTED
