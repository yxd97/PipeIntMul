`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9IqJnD6YjaAEMbxhIhDmC7HcVmBsfBpkqHHLkLsBSB8tAEvJdycidZm28ypDHECF
0MiJWRF7qM6tCpu+ZKJPxs2UqrRTU0kGEf9JGZVYzIwtbYsYC5/Fwt44BwfanLtq
IlTvudXJQIgKT21iLou/kbN/KCRjKy3G678IqPtGhKgzVGyl7287ZJDbAP3zN2qn
rCf875eemxYBIfWnpwxE9o4CVYQ3Supdkz7euUgybXrTw4P1t/AZg+dqQn1j//rQ
TpxKpOGsSVqzf1jqrqNBMEkBf1UxyvQgkDfieieFnW2BDhEv20SzH+6TxAb99jsu
zCcqC3XVH+n2uhDz4WMMBCZT4UPGxyYVh0BP3EMz2YlpX3tTnKcb95MHOcIy4FyS
QnhS+Zz6LUAvS+M+VAJRdndSlcWVmMdhBS3/0WX3ZFNVVxTSe7KgT3ixxmnhe2lZ
`protect END_PROTECTED
