`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VrwOWY1SAiaPNl7Nvt/y6palrWxgKDfj1FGHeJaTo/lrKI+PZAVXHuKTQ+8JQoST
pUlsNz4ZWQQ/omb8dVvPl4QIt4l01I6NsuGLi3N2aFuBbqsWWIx/gZ04ckn5Ek7C
eeoie5+HnbJx+14K+m6rKcf+tv5sHQjQCmRz8G6tKM0EnZ/L7Iz1fyRbsxRd3Er8
Y77JO5km5ROLqE8RA6J86yKhTuTYDeWLjiaEIsX09jVJJyJPl7Jg3Ikx0UUrLcHU
anP7Y4QDA8F5Cw3I8bFLas4Mvz9vSEH1J+nokuIBH2dL2CiDSEW0mCBPHO02mKb3
GLa2APhiFuAMYWqS+V20mhFLO0a96nTmC7onO5YGoj9NIUl0LFM6CYxmQEmXgMfI
ApD4Hj6IKSpfa7mU4Vt/YBc2veNYJi2Y5VXPNM3qQCwdylJYydbJ4aPi63QhNLIh
yCRSpNaqVopRb/kzWBiJ7cnLEySJhELGGWtAIOGAn3+WI39uSYkWfurPYYDK5xv+
3/Gsi9s5HzkSve4czxqwP+gBvv3FyloVQbqjIsav3QjhXrJ0ePgWZzoQaMGBIBiM
fWa/ikYWTZ+XRJmNP9a9KOAMXaYK2UpF4hTUZP15ESJNh92t8wVHl92YLwThQ4gY
1JQdB7XjBQdkIApdOtx5D2HjKKhoRzEUD0FR6Crm9yClZbmdsJni96PxU3MCZrdV
ZceSk5uZ3Esc7A665qDKqokCDAm8s4ratAUBCAF3ZoQyiHvzuIKivVYqEII8+09t
8lz0/l251RbU1q0Kr/1jKa//ljjyxGfYw3E1EuaaWoVQ0+UA5vVX0AfDYMwXhhkP
12bPLUzph9PUluP/abvchSlJxPsqJ81P69DxghqBdzDZ40zU7XtNgMaxX5AhvWFH
Orm+B98FOwe8DiYzgsIf7Jg2srhAmVjVoP96MdohsXvRLGtf9IrtvK8vt4Wo6zcM
astbfWJwxNs+fPTfqqDZXaOQRa1c9cKm8j8/mPYpCvqi9mD++uW3QH8e7hiREDca
MZty99ZTfMzzsLwtgjl4SS7AVOfp49whpNx/dJhvXY9pGhkAM0wKHs21w0XIQINE
ci5+uw/SVKLJuQrP2fbuNi68Cnhjl73GQn7jyvzyiQdFRpxZAIBB83tfKl4bJV4g
wMDdZ/T3TMFsBUNYPKOh7NF5jIawau83djyEA8cv9hQADfKz8+vQbZ5DOEM+4PFl
dK6JtVSpV6nQ/SAWc3/WDUd9inkIbe+a3eiwx1PsQeCm+rclVHRZUhRCqgCTTq8U
cIToYMARfJv4P8fi6rcd9TghoEy6VcJ2QiO+wqgmT4/c42BmBnHxXJNwGL3eYpLl
LW3jAin48rUY3KZciSZmRwz9a2U8nicjoxYhTLe9c+rlnhyCERoFHGxhk2CLJgfJ
k87HrZuyCwLb5IUJEAdWTzTl4UppcLNut/YGfDNQE3mtFfp8dhhn/cN/Uu+EN7yd
lv9aVB6I7ls2UDT/srKuxkTLTXVe5DhfTCTSoZfp7qz0YGix4pjUDEw4GFM/S/G8
iyQwR9Zclt6fqAo1MniNS4Pg5XKcb6XhcF0dqXA/aWy3CRv6ls/YbfzxC9CjG1tg
6yGIAlD4Iu8sA1c4j1XFfc41XC4BlzU5vHZrPV1ige4paBoaCK2Ek3N4deZ+A6XC
tk9HMiHeZ5ZkaZu6cDSEcXUEPM8AWfbPkPNRS1yJStPiI5xEZxVf9xpbnkYZn5N6
L8/6GzXtD6nMQsF35uEghPP4tx4lBlIJs9eMdC76MxJue1EjZcC6Ns/ZKV5vY1fu
16aOf1mddSGYzW2gik22xVXY5NYIcdYNBSMLBmactE4zMRLphw8EbGQZZi6qg8K3
yhMWXhENEe5DGoNn+riPsnOpmG2pvF2GiSLEeIBqr5KaLZSTU0WiwGMocXz9LODi
wvbepdEL9B6mP+q6Xm8J7tsNZrMxRvOWXe4iVQmmYRJQmBl/Ypyk2EOxRFZsnCzm
FAc4zimp5i/vnc7Eu21l0iUctS6Rik6xBbcMxqOGs9SCKa9jXQJHVnVBBf+AtAp0
7eVDEsAtXCiSUkHvGiaewboOb+4xY7zjg7aaTtUj/F/JW2mhlm9giK0rPGeR9gdl
0uZTXw1sKFN8VpUGmfKCxEI2WbQ/KlyzRBA1F4xytdQqwUj7a12LBWq4tAslzwJ+
4J/61Kg03Ve1Abx/oLZ3RkuH7oqoZGBPMWVRibw2Jx+xf2wIDRS+tmSuNwXdcDNJ
Ov34DHYzHjIBAfVe9OR710lRlZgbeCcOlP+wFlIXe6VuUnS7u15kKnfSrGnMHkU1
GVDtKHeQUS11rn/hyNk3rFhq1dFLu46sq9Qyc4rt3Nw48WAQ5K9wKoZ2Arv3f4YJ
TJbnvxEuuVCYN/zKk5ob4vfhUr1WKXcEJzkR84QZ5tL6TGKhs4sdEQVPhPVnhZYo
0DFL09KQJ1yrNI8Rx8s39DwsXYPor1sw7k327eVy7Yt4MYiF69S6qq7+Uv5eHUn3
aWwCCDpi5IG0eGey9uuh9ogEhvrRArAMhccef7E3zQ0RJE8GWYbu4+GC1NjbtIIB
wCkQVQQWMWEAZgzHi49hoplCuavDUiV/F8R7puSWaXtHhqlfQQcAtprOTAhp/m7J
Xhd0DhClC+Xs9OxkKeGkvdTSVrId1bkAxpmUZyqHvMtvN4k/YlUrkI9RebB/8m3+
fRz1DOUC6PrDwCAvbngjquDekXI78z6nWkgdbQoBM8YCB2rUx5tSHttS4fJ3/BN6
ZzzzZgnW0eJeRb7vdaNH5ItsgTvzAC2fx9DVI5OS2iwf92MzxAZVX2LESpyWCeEN
N7guxdUPK0JW9Qp8DAFIS2WzfQX6fXNyKaN2GycUgLBJqyJjThfsFFLqHFGYS41h
W+rAAH9+n7b7RJWVwNU+wz9tnf2F9UpGtdzxEmqwQa8xzWqqgIqjw1UBqfnNorm3
XPch+kTr5B1S0fbfWR2yc2oy4HPwRRtNbNUId8VFDxL59P6Mqx0v+uyAH+X7yNKf
WBFM2RM89m1Rdf0okV4sKNovDU2IPv3F2Mg/hJZRymdla+WAP937JZ4zbPIgTbsm
mV7cZKZQwVCNlwOrvhAK5NJ1PZofAmDxRTHkKRV1aBFkbBTY5EFNA9i73RlNcNoY
e2zenhFF2ZsbjKAj7PWe2kuCi978gclFZKjJhoJjGqjjz6vVRChVk0UEnXv5Lupo
dHlS9JaogWIW/MrYQmPXkDyaN0WbH2bpDs1pmpX3nYrP7D6QhlAfGwiEM3OhsY49
sAokloCP+bOJwkDFxq6DWL7fdS0R3Nw1bvxxaZGwG+6XJjo7v5CX0+LmvKzdmRQq
3a0ph9cka6qTnxScr/6/ATijMJQvJ+op2IxPKc5+0pzoY3UaVEl3AVND9Lmm6UjR
RKaET110V4yLvTUPc9iOBMgNPolSFqQX2I+hw0yxTUubactsmnYSGgSqB93zQZ/B
ojCL6Ct9obGA2lOMeRdaehBIXeZZ5qNTVb4uyRutZ4wD3uQi7XSHu/TkSAdP+w7q
aOynQ0FS6gp4MuXKUFirph+7Xk45iZkWksbmntaqdzamzdeI6gS/rOkp5jqwyI7Q
YGOk9HzjmkE4eDn4XRrp6IPOtiSUuqbFT4a3nFAQsrF5FmPvaG7sLM8mg4+1sa2f
uUpCJtF2rmLBpoZ8iZJVHYLSRsseoiWkmw0Emm2lX1uhhzhTriw8t/35jZnWEwxT
2ZxJtfxkvQXfI7csx6a4T7/uACObxdqS1Hogz3R7Z9A0bP/V56k3Lmf9YpHOCsED
Ghzirz0vvHgj8g1bzfDJrT2ugw/+PARhsToQdalrNfB/sOQUNxyn59gEchAuQvP3
LNlWn51pOHkMCJP4w+H1ndA+WyW12UWps4inbF+NfNYaCS+B8RnLOJrgRJhiH+Wd
8Rw7AClLG1TLn0KOhR5BohHvg5kIu8kHv2QbDNOzzhvffsBtiCvFOT5EQMy+FjJC
Na9B1umN3FlRA01myA/Dk7PeXrrZpm+h9KSUTQTp+R7I+HSRAbQu0SBJTrM3CGH0
AOE2KFQIfyeq74IJ8Tqs0wH6Ds51+aP28lj/u1Kt3PLHUSrhFeOFwH94VSjAhoRB
3g1VHEKjF6oyknIATPMCaKWGjkMyWIcGDo7slot8yg4AEhwXEq2Dk3jzDr8b+svR
ZcQjfjrlE3urLr2lMMrxAP3zT9jftFPEKwDcOAVs3bM+y36k83dnUELrJzWPyoQc
hIO/V7rCrlVfFHwQ/gNfpCZTCB6mZ3lXKtYD9cYmiWQBsAeYGaw36VXyrUTcULsD
fxvo4kWZy4O/vEK2ZasnDKG22nayCkv4yKi10D8GveHsElHE8gOF/0ZYxUqDXt5P
z/AA/ilBBCjUMeuLWVwyaLyTJc6NgsKjtqw0q8Zmd0ErugYSQKGxMoagP7DtM89k
M5Kc8i1sMm7eKZBzBjFntdVEHCfVcSd2MMCKSOQvDTvPtstZzy77+jJOsMRh4z4L
jrmOmxQHc4D4I5wTDMFl75dUwcra+p+pJ3BRBxKi3kvvpeWmGzPadz77BJvdLg77
t5sTg/dRX59SKXZZ5B2vopDuNjpkx7AHi6XKO2yHU64jUcze/vY/seAJEx5OeHM4
GX0BebjUGwBYkDuoIpEC3KdfpGNfQEf309AiaX8qXNz0e/1iwRFb064Eyca4P+ia
1bE0wyKYGc54EMYNMBxhb0EMRYMWe+zVTS7xtt0xSSXnDX1fZeaJ2idWxtN69fKu
OMi1ADEv8rHlJmRTyygQpLNY9uZeSWa3t2UxcO83Emf8gqWHoU7MofHCgc40yfaY
7RNCnqB8k9vM24qs+BE3JcUvsosGpd3uaAw8TNcXvR5LCh8+OAFJ1TdEPhV67oEy
taXKEDPRxe2G35Z7CE1FkX7ep8sB2dtUirV53uhNLo4ovo4MDs6ixUoU2TVetOeg
xTWFGYMg89HsGoNoDJHgbr78ak3l41kCRjbqTaBA/dHqVJuQzm7Uz8epCQLs4ds1
0WTiGlwKU6uBWU6mYc3PKjo8pQB51E5hQ0ihOlEckl2gmVmzvYpkLwNfE7pAz1zT
FgQ/28kaccaKshaj8/FLHJOD/FW1oA2jZW9Y1ZAWtU1wwuRGVtnUIfE0Zx0ntkLv
NsKb9DCNMCn/ee+Wi9Cq28uiwWiVvcPfKsjoQ4V25F13KTThavrYsAuvWvJY4gXm
kBNeOGyDLdecef1h42pBSxh7iOT9aIK7SkivnaWXQ97BjvkXEPJ2zBdykxie+Kd2
mQHHgzz3YLWHBurEl03+owC7EcXuIb/HpRLR1iHRGppoqI8T8mo2pWeApb5nv0fn
4f59iK/bIdrtUO5Gua4XOmbv3wqS2hqAxWoH8qUpm00n5+Ca1QfIA6A5n9jF4sKF
FowNaioyfYR0maZdiAO38Vr8xC2ij5GLkdlpLmezO0fmvhJ8iOz77bBlJLcPpf9Y
JJpau4Nr8l2Ndx5omLgD1H9k+gFfoCXKKbxNz/llEmx4Hqq4SmrrcGUv4QuNMLND
C6SJsAvuxRGDQFY5pX+M2R4RHnnTlt9VlV60tqZqxclEgej2PO32iXMNVggPSaNS
5fg2zTk9AslIfcwmiy/DP7U9DrkdmjSmAC+pikuOUNALHAhnbS+dtiBViPIhgwhn
QnoAK79UxT6tlEfINjv1GjsEm+HHARQX5JPz66h4rYHZ5eqnymT0goP7YR4sR65T
PTrY+85EMyau5As+7KM3wcYUb2kw3+uZhR6fkedgTgVmUJI+Ph6UTrWxtWxfqUnK
h3xbyYc+yoliBHcMiLECIiOPQw7oN0WQfXq3RrotWABwXrwGLaIKmjMM7gYSir2h
Q1hlbn0fDSxfkCnm/c6atGn6/CD5FC6fVgc1wOYbrLSjCcd3UDHLN9MpnbiWtSkC
7QY1SQ3MTSmB99VjEi6GI1Ulcc3SzIRgbgp8aDN2FW0hRLKIbJJkLX4djgRIIz2F
iCGarpMTOMHfeDc5t8ooCMDQ1Nhr0ys7f/eEI29ngpGOd5zZWjdS9PnwUuja66yg
1VoLWD/6/5he4/ZMaPMHFzcTWn9TKs1KUDKpXQwCIoR7f4oQ1E2/NcqNI8fUBVt0
s80MR1HEdjH6NfyG5qLq0E6VCOC54MK4eQCMVp4UwldxXY9nG6ODWJoPKp6HL2FD
CPe+RuFeUoF1d2KMpev5DXPxX4SWJ+8yeHiRcHcBYQpz1QoKaqXTh5Ik4J+B3AAq
+NZvk1oKr89RmyDRuGTyaBiIi+I5D1bF3QJCIW8NluZ7Jb9r2rUCaRxzvmHLdDx3
4+uixHMAkaWN+Cb6daKCwiwFSOHeH4rSeJ2/HN78vF/ly41BaqIpcuRQU47l8vkK
Dt57vFol0GvVsqVt+DKsJu+lTAqdmzlbVGoPERGg1RWJ0TF3HXBZnFFBTBjxtg1t
rYEobl4DTIO2s1hDYUMiVRUVo0aBaqgjFUscWbdsUnjEQhlAedCoGRTGF2OS7lo3
UMr7yFQlF8UvPw7704x0zN5z6EA2XUKZZTGn4ga1Pi6FSHtkmDjftpurCJxqF1ix
dIH4FJMec3J4Hv5eRZoPNstHiug3KG1WL182i5yZAKrNsJwq7+iSNOcsk9Wr9Vnq
TfJJ1LB9UggvVB8QGYjgB0+Im+/qYmNbFaoat6wPZQ7ojjwj62azPMMT+eibQBKh
jWdqaMF0UdW1PUapX5Vs49OKQL6CBgc0g6OfQJv8gyc6WPsGC3Dni1vq0Z3ZUeF7
ZbwOjd1vQJCGxGFWnmFHxQD7kg3Ia2DRaDGEGO5Jnr7lgKn8shYpm7J2wEk+yKW8
2IJlVMKzxV3bpmiESocdHAUNAlurut9Gmxp4ZMdrWjGFxbyOAUBzD9kufeq6UuLM
2NvHCC8ShQ5Jb0CAEJZxEq0xqbRWp51hy5W4C1FnrqnKRBEcEp+HkE3Edt/81Y5c
mK+fk8dkfr575OAOHVGWppBZCOPXquxEFW3GxrjUEXuYwsEAPIdyxm9WQ8Jp27/f
8Y9f4JzCY/SJ5jz5Qo86e1JW/qFCzM6j2Y73bJW0qLqNZ1OV78Djc4AV6ixc/Zi+
cHZyQRAOB/2C/YquDzOHS7XLD5qkKqla/NtekN87aSFgj32rHcEfbrli1oNwtZ0Q
tGvW0Irg1InHUtZfGDLZzfnMvs5LXYdp0GijeCnVUm88e39Iam6EwOogeb4SHNU2
Daq3lOUJ2PZI8cimaJJVI4h7JMFbJzNikU6G81lv2xbWX6+aBXR7Qnqh4dDdquFS
PAybdS1+MjauMOSHP2g9H4ubttjv6USjbtyF1yTjpsKFANw4H0/sjIFq8ND9d81w
dpQUpMvzJEOEs8FlKCNFppN9tCegDiIqg7nU3ZIkz1ZfVwzeNe1ijJ44WCDH0uab
buP8luoBwj+oQ/hmRoHap/0pdtsbs3LFcCofVX9KKesXrdQ2AfxE98lZXpAgnM99
0P2lqcuq4a41qmUO+hRnEgQEHUjvTpcBYdF2oU8tnHfzmKUeOurR0sxdM5zKnnW3
DehRi09XkUcbpm6VlN3rSlKgEtmnCpz6Z/U58XySI+TnacgrKrMn5GLeAX2BqnH0
1Hprug7xcpCV6KaNjfyeu8IVM1mnRHghJg27jbm8NxRcC/glCfDesygEt6Jx4EIt
utewVM6nQ5qocPIKS74cK+O+NvHU+FtV/yA5kq9QIeD4Dc9LOpyq8kZwtE6BeVcm
cdM0ek3zk+wmuerE45jCQyqmnt9kZXAnKaJxHXVyru8Joa9042s0g4sCwVL0Mggs
3/6clviOt+T8QynxPwwmdFmQIX/ooSKfC2tYguoMRbixYCxxg58G7HNn+c4NQOGJ
cQ2NgEx06PCOys7HexgxxET2T1ThsBmeEnW3ZmRtsqDUDPDNA0oJuAjXlfHx4q23
KLmPUhKRWIpQ/26vfUcyMkZpe+o+8NDkiCLOiu0e7y+27kHCoJQTJkM4xNlLv+8k
NSZndK7JCQvoxXIK7TirXtbOrAGPgw9f0hoDkop6wi/XaDwLPE5PpduiDLHsPsxM
BIRuxnrgGRS0wy466F8qqGlQ4Ri3Ly2U+RVyWiiXfiUt5AdF/G3knjE08L2nOK0N
QVvUJAXpD+Hi06IccHPl18fVHbLX7FyXyqKLh7dBXz6wGtMr7FCVs4CUAONVzW2r
HlUW25CuRHX31ZRfPdQ1TEQxnIx9m31Mot8TmllZpLlMMKfkNPzL59aBEOwIyARC
a3DbIoGe1YSWs/ISvQaCIUwyhawLKO+Cgex30mpdluFquyoSe2dIIEAjFKyoNtBz
BcbkmOnbhzbzjH2nYMtKGXkIkODKNjUtfnE1L8N8YQqssIALc7z3wU+h6+1y440m
RHHzB+kiJPPWQPuDPA4jIz2J161INr9pCGbNvf32yLbD1xCoMjLLD8IARQS0EVE/
S8L3/+9aBx0BN/Uug9OdOQQNHIT2vRQeYfuKv9ePI2iRw5AsjImGpkJzepB/29KK
TFmHUIMZQmSnzV9mpthyXUhZmcNM5f3vD2ZNJ76Y7d+o4U2afchDDKIq//9EV8Pj
GZ9Y8nJsxuMP1rYXm+gU8fNxsPeS4UfuJN8H2TrCsQOqugL+GUT5f0bYDB70LTLg
slGd0R8G5bRQRcnzqubXWjRCBg+IlqFwsdGGIlQqoe2Zbw16EkiOfTfn8qTjmcym
J1PH/D8ohTHlm5NuHREZYE6fbJCJ/2HUi8RFyXli5MT14xZX7t7M2RzB37aenPpc
33Ocle57+OUPrr/wLOg5s/Fu+hI1+ii9VVsCDu+ZAOZRHqsES0zBlwsJZxBt5CxP
8RXJ5fHkM70tcLfXhi2oKQXvTrNB6Lsenk5gPW0nwGLQ1s0UngOeXiIgOYAYDBSr
EO7pY3mkNQySbH+aHHVf+9UMDzVZl4r7aWKy/tUqK2hYn03YPj8hVX3TeM98ypLI
aRrlxFI2QsH63sBIN9LJ1TzADJYxb4rm2858yXP1ks1m+og2ujHd3qpAorLtQGiN
nb13pIzEM5gvew8HP4hiDUuUNeMRBOq9yaH3sgtMjKR7l9YwZmrHakMvfYGVSe6N
zR4yRTpI1fHKYSZMbJ9ubaDeJ2P7QSAczLzLlCTIbnhxYVCVS7OfRV4oWBdtIWnV
5EBG9Q2mtuACf0jRehwDLPU+Rl5tukFzC6pQUxLDJwCeUmJtnEoCcR9FNm5YTuC5
AHv0jhYzSFpkPuvTiU/E+yTb4GeZewc2QpdjKD09v2BvV8wsrP0vxfNjM3L8CtWy
1BpkBdqQWkPro9Gojlq2ufWKzO5oF540x0kFbfFDDABnjhMpyYEjymkslHtEis0s
cqrLd4AiHFEyt/uQXW/9XpDX6iX8bqAfFv/ZTkjBtx1Tp7CTGh+evcHSXqf7oTjH
c5KifcGS7bHWgXpuu8iLfxiSonWql9FQAtNdm1+lPqbYPft1qhpIxyaADVZya5fN
Zrm7KQrJBUKp4ZSYC7DGCewzYkr5VJjVC4qUEgjgN+I+sfDA0I+4fQbDW3+2pxf9
JYMoHN0nfszlQFFcf8PCQMk8huH1Jm2XAWay62hEhkmwF+d452ViwWO6EUs4wc+H
EjTo9gN0ZjwfSrBD1R15wfWDt4eaL8Ep7I43F52WlASvxRlOS7U/qUkrwo+KPO3/
mVUWAFxtCPuhhlQ6vO3sRVhZkKR8j9CiCQMXPRQUtJ83wIa/Tv97cmg/vdWWavfH
sW9T9GpfKvN8aXcD9rnjje+LMinMiIMTBKf1P78ib9RvSGLVdlUgcY8EGJaxyYaz
fk8IlzoLRDQu7CtNS4UUjKyvK73NIMEwcWtFm7W4OgzpL+YAZXw7KM4Txb2BYVpJ
HiWfHRiRtjoQgMbbHw4Hkapi/dGVpJwem+varr/URfK+dCBe9ApfzZyqr1y9ny5T
FdyVTL44cuDOXkyyUeFhD+kufy7+LDAjDvlk0t49dT6kIcpLNEQShiMgXtyO5B/L
6U8S7O9y00TjZiQlBnap3mrh9aVT6sLqQlW8sYR2mygWvqhjwKUjvbVClDkQin+R
7gfZYvSa50U6mCgNPIoNqciFGXkBNKIGJOUFY4LfVLxp7DLf0BXvkxhiSQzBUzpv
bt2WLN3t9RYHT/P0H3rmd7c19477EmJ5jn4IsuvaxFyb5l9Ha9nH2UyznydgKrpi
nbB6beR6Jm85PgAa3DZi8oV1CRh2f5PA2vyP1d/G2pJ/mzAdKwJfBa21ab3jWj0S
ZIxb6Q7FiqoXaEWCK+9+d9LquxTme7sBCkt34EnKNyrXjPxglfOaRkAW5go2B60R
UH7MA01drkPasNLx6VEvcSpfa5awpytAlB7GLG5XpNdL6CtHYfVDmKThJGk8Ki3Y
vAcmgD5U2CoqPAUMx98zpvXu7D3dUV/fmytM3rbf33eWajLng5RNJabCav9UK8JI
ep33b1SzHCpxPOe6bA2WoiBFqNE7UzDHgMGMcQlF5ZjMsTXn8DC5cXOp3RPJeVJH
Uhh1Duf7LGWlTXZyf52Iq8wwRO8kSXzB2hIRFTHfNug8n10s/oqfIWud/D4JXI0l
C3+iYhzP67bO1F/kc/+YBWZWr4T1ftPX8rNGmQHQFrUVGAtcQn3XvJbc2EyFb6uT
gAcRx6FUiS2+O8iggjBTuUe8FggUHER6hwikSUEuufnBJm89UMOmKSdtHooEmv7f
6H9pBhH8T6tC/EUbT2okEi6ZaW7ydpJyrjUnzf2qjTN9EssBovnzUe/z149z4Bwu
guJDtXP+9DFJyLnSq/IsxlKM93Nw+a4+g+gYI/XOz0hT/9n52wm64RBV2DtbSoEH
A3cwg7D6qKudvMByZ/qDr3TT4PGjzK1zS3+kQS/aXqp8pKj7YXCtRBBG74kzMex+
tkj5kxjb6TNI5RZ6XQN7QpsBK+gg9DTI8nRCN/csgeSXrbc5vX9vUFh8749gJb60
p3JePa8+LZO+k8zu1IrPsAjU2M/EX1IVYzMs6tSNpPLGo/jhCxftC74ZsE7x5Zpx
9Ob9PvzeZ7tveF7u6dtSbJhzU7m+OyjZCRLh6dzasIMtwtQelNq//xG17EXu9WH/
C8Tv3yWfL1erwRn0zSZbZHHUVlayOkZBmvcUnGHkot67sbZdmULllvAbhLAKKx8N
hWFe+01nYnAxIMf+mqiFQ61NmUPwtVBNZrz/1MWggpIn0o+aFZ+x5sKHRRsNHlMu
6ufVlbRWUUjL6jLaKXh5ZtjEWn9YZHiK0EFsX0dbWmB3t448uz9h4wD+Vd5fS+DR
t6eecLtvIooAul5sUpbX+JBk0exFn13yE1/cv0Hct81yVhXHZJ21rKhASpKm1lmo
2z5gpFJOK9BNxPPSuaZXQ9i8xrrdFw5rGvXPXKTWH9DhCNJ0paTeubWmNyt3CF9U
y1lB9wv39JZjqqF5HGYMFzZGYQxAEuYslTyWDJ+BZutZYnCU5dTP2czKrFmKfbZ1
XQZ9Koi/Y7IqktxaGobfEkqEp16eGhGigLQOSQQQXcI1Hi+QzWqmXqbYdlpPhrKH
gfkBNdWvXsW6E9yivG/b7UFa1Bqt+NeA3NQupU4yp/ageMNsY3cmqoMtgw1waC7f
tu05b060kDY/oDO6vk/ctYJYHFzLetvUHuDoGn0wk49n2E9cnb5TXGQ7bdHjotAX
dpm/RhZlyD0UdBXTCTI93Q9okqWMUhSXKmM8Wzb7voP9pUWtmJkSv+/mlEQ5gqr7
TeKUWAqF0Ibk0e7r2EW9lCSttV0Nq0aXhL22xsTQGGbMlm5c38MZ8xxS8Vvu3fsE
f3Yx499F6Ztu+9/s7yzSCVhquH4uIfnfw8NTSb+eq6AWb302lFMeVdTB9cGCj3so
t7qbheE0dWSzGtGVZ6gn6qbH8pr8bs9Qm2HXvPqr8yoy8CXmz9qlXc6FDfXqSF4m
/HNu0GK6U5SlWsnEPSqJdF4FfWpOiIZ3kdUq0ho7nIIxBH0VGoVTBaDFFBOAlp64
Epr2d4iWe7aQfZUnrrFm99t5A/IIDTCQqTlcQEJQB/+B6F2dVTo2jPQrjFAeDb9o
d6nB4PYFbTNn9jXST45E+OTkoWsCn0tKNI3W5u5brr7OmXY8cRBqBgrm24vJrERm
PkWgUBUPi7INjxXNHSYdz6P/Z8InprxF3a1NtgjghMrR+qXWcxB5kKDMbSmgZBqk
08eQ+kDzigerogrdb2SM0dtMypZxOfw5BwQ4PY88ujlejFVFQRbI4F7/BNPc02Tv
8XGQBMieVPBF9eHYQbgeVA6ZJNcruUCikWKLvu287khq9XaTfw8HuxZCnbcm9JfZ
EBkQviZztM8CcMnHzkzbDt1zM1EvofOQnG26gbpBM/1avxZDPDBGzbCwj+Acz/yq
3DJcUo46rsddU2iJT41h1xMr0woX8z6VUUsDW61LN+YhAK6XA511EBThgAHSBHoT
ne/e6gqCULG8hP0+XmXb111K5DNQc+7Bm5HbMYcMSgRfh/+HrdOSoAAmiTNqA4H6
Gwv4oP/uGo+mRD7qnPdv9XUHWy14bWesDPrdMksol852wtNLebab1EyrFQptg6m1
YkGxMYLSyo6Kbw3roOtKWRff9cgXO0zjHJCi76SlM8z3y1l+QatnK5/g9ly2SSjt
anlECwtn09ERsm1mqV6hWtyyWmp59YdsTP3WrAp7R/m9IZaQpZ4LcIR++4P1BtCA
qcrUKpj97HC6jDtG/HDMU3sNRJk59fM5flDKmCbVSGzeWjGR8AlyCcX6E+9skcHa
Y2nltAKOYlPax+S2McOOWLKCZ0wqdRKGZz/qwRlB75lCCOl3hCg7oH5QOtM/e2CH
NLX/VlAweKRMatH4ZxgcFiUTT8qrWvXrEIB/NzTAZ6CiSmHIXAcFP3tUIYkC+AFa
YTDYBtcC3otF/srGRYv64P835+cqTFcSmqUcLAvDNsW8Tfzqpw5cMipsHxSv3n6L
PFVgIIjDAcNIGIq8YHoXL7HbLAIXa4b5E1f8S/1YrSP/sr07OJ5r7nIFRiprtZbr
`protect END_PROTECTED
