`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mu3d+kj8K/WmIR1YpWD7keB3UOy18arV6TAsucTgVOMGvy8ccYARTX0ziIWxYH7m
2tNQBDka93gtPUmendOJtqDgaQpi4iDBieEfJG9S6EsvfE8FI8qoMXXymESzinvQ
afc0ZiUWlCbyvonrbNUrlOwspYxrW30sC+hJderKZJs4MOrAYM9pIf7PrC6JFp2I
93RBWl/MArS9EdD+h8Evy/Pmj1/sWTB5Hc4yL7vVxv+zNo6YFnLRXlAd+gZa6W4s
aNcZrv2u9BNb/z1/cpVwSEmnCbHwzwImD6Qlw5Udmm3wDM9L4Q6fWkzWYeupRnPI
gD0Afl9NZVW0Ro7Pi5G/K2FsycTad/tvNcOcVMK+dDUD9SDBfDvAkFZrZa7WrIWc
8CxojCF7C1BfiJ5eZ38J3D13GZ08lctt5LH8/IRrmk4hoQ0CsxRL2/dyHTncIDzg
FPOrKJYQRBBvRl1tBCVSePK2eLI42l9ud754CqyJQC9V0Hw43tqejzOYjXjbDzJz
M6jhdCh6dSsTyaccodprMqDNFlUQ0hQc//BWS8Z/BaBJgK/qzsD5rOl827SI9EW2
ArvfHEqObEBjKjCYCYszQXURUhlm0t+NWRHBFD5kf0zDol5QX9/H9nZYjATwUrax
4R0+84gnRmludl7VhJA8ajhL8anTxKgFmjkv2wBSPOIYMvKowfeG8q5CSqXLV/TB
BcaDK0ALB8GX6ET8XxfM2DHQ2a92Cz15B7tMxmGWCE/4Mhw94VwzXD77aAJ4R5YF
U/hvvlAD/BMU0pDFOQ5i8TIoX/WgjpFMRamj7rfNOat0WwN+UH9V3tgmm9ezmpmc
Ipa2eGVeFhpOzkdgoiiJmM+XGmvsztN1cbXJ48m7cpxrmeH1WJgIGlMHsuEkUeVr
wUhQrlhFpbhCJFV3hxeNMLJucjzt4JHYxmtGdFxzLHybNnWHH25eUqVs2Oa0RjHF
M2c3B5d/KQiFPTE5Tg2HBO64rTt0F68IvqjDahzhq78dC0CplGiQiXu2Hojahn4w
LcLOPa9hSAwmOJLrKki7XQzxhHAFp3YLh2jazDAXgrg=
`protect END_PROTECTED
