`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ybtJQserz8EsaoqCOaTTpJ1aVTBD+hdwKXUQcaSuvXx7tTXATsF4I9Y1LBk9mXxZ
O+mel0ruUU3VEEqBkeV4AzNXANiFk0OvYhynfKpJ/cQCidb14XC5A2iuSPj1+yXY
gh4zAaJSYptIIv8pcabTI+Ys4JwlqmxOXzw2ytr75r0lzD4u5ZeGZZcedu/M+4B8
Fk1Gms7jXjCD7YbB3ewybOtzHfVjwMRsar4f+q+C8G8Ol5GIU/njJDUgeTSFTkSH
PnrqPSIf0tGmWPfG+7yBtNqry7W7kWSKlfqv+BTcUWAHb9hyjX/MpmKxS5kXdz9V
Dfns5ttpN8YcivA8ptTnHA==
`protect END_PROTECTED
