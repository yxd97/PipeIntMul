`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbUSLlphTgXGT3GsU1ylDkXVRC5Djy4bgyg3rKKESUgODUrYwDm2lzx6nk6Sp+Pj
SzxpWZNSH3ABVomXeytyUu8UZz/fMShv2hWIqxFk9/DccDCnWWH4bH3Wwn8x1fYz
yoLj7JALo/6vLmcimTAWa4G2XG8oJNL2Y19edpBBU1BTbzX6twbUt94s8OOIOTO9
EdNxLf8rh+HP/rpE6yCnZzwuE2WtPeErT7i9Crga4y0lmMDBwdvs4cDexHlsbvAO
BoD0SfWgFngdqTt8ORVJ4pivbaBLeQS/3bn8Lca7Lr+t8UwH5RsAmDCLT7l6btNJ
yYRWKS+ZlclrCZMfQuuhCjP6mAg3c9GpHy2QRZ79oS7ezeQONgKd+OIoN/6NlFEf
Jyg9gkKKXt6iEv7ej4HvSG3A5ScnXxrwE5A1HmBDucOS3PtEot3pnXPvJafHvALo
GFsnCoO5eW4hZr9WOplGJGeqUr9l1WWxswro+6n+22bvs1yvvQOUv6B6NDINC82P
Wxv/peFxgTHHzfJTfHUMtXtnLwqMMuNb3TYo+aYIVV2MNDUSvYkoLApOvzTUHikC
S6mSrttacPvBLnLtDk1AtqxkVTXMm7Neq+q0ZgQhVVsEkMjVh1SKvf3ptmKDn/dh
uutn7IKX53N0XAjDNoZ8Qw==
`protect END_PROTECTED
