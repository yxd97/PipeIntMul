`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh08X9YLMk+3FfGWFiGBNqdnRBm12WRr4ePEwRyf+w+83UW0YGdch571mQP2DTym
o+hi3qNcWUyZxzFt3eb+nlIThD0j5r+7k9VPxcK9rzcsITS+DJwwyz3KS5Nmj5eO
gPoaE33bmXBCinxiZ0uI2a2utfl2wNMfzJKHF/FbfsjcOJ5TgCh0etQwAnOP2FPm
n0l9xdzyCBX9/RkKWiQcSgkt3ZIySwoAl4OEAtMw+I10Tad82/CsBZVVz/Vecuim
LnO/lGWliSgf6J3WF0zUZTqzJ+neof1Ov3ek6YAquE8kHoXty8Hh0IZL3eUI9bPZ
WvR8hZ4sgl/sdnEgzza9IlcWJvC36eZZUJU7SUyNXvugJAUmid1x5TXqfrvROWWG
kYDQKlAbBcobDXrFJVf69x9npMMJRoHFwEbFhXh++Ja8QkUMuskXLIpnm5n0enpF
XNf8JuukkLiitIngsFk13oKFIdyL9G8vjjDt3FypZ+Xck5NDdSBqrECn7ziPcwWg
JKV9iwEplON0DzalbbgcqDcZXD/SdwARGCPZSToukWNE33noUgrDSRjq05UNtecQ
B0J84daYIzi/YLeEy+zdCJzC/wFNLO/zK42Eu8UIL1gvk+hiRk0Rl8T2Zly5pkxW
W49dJQZeU9y+sfYmdCXt21apYL7dihVWruKPk/VB6NgV2rfwn3rhGDdkPm4Bj+vS
CS7/Qt3xcQH2koaMlm9HK3P2NNdQX47sgNqwRzC8BVbwmddtJ8k6Uvq9bD59ysh2
O0wLEGwRU8chUQ7Xk0O4DhGqbUKkbsVhSA+owouzi24+VQqVl6Dvhk/PUl2bnG2W
`protect END_PROTECTED
