`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LfXdnSKdbM1kNZxgYG3nCv7T3enPvJ9AZVQSi8YxNAateqDzS1PJuvY7QiE4f4tk
CB9swvnvt3sWQU98LsTk16ArXy8CxLyiNf4i28dE6/Qc6BE/ARQNz9mv5pm7pC6b
+h9JNQzNMUUEkap6EUwKwPp6Bmp31rAOIJAGMuy+zD+ejDCbapLLufFs1ZKE304E
aNLgKcqHfTnkGRg4l08wMB2bIp20BMFOSBOZxKxeHQHa5minCL2bK0xEJhVwq0Vt
3Y3sEKhNdJ5Mj0firzFA/xtnaKw0TA8pY+UkipDPj05nPXRKSmlg/ZWimNAXG3sK
Qi0r0TRuV7+JlGKYlg75jGwfVtwO3WnBy/qlp5u7fgbkRgCuQeNLXpN8dd9liD0v
7MRe6zlvAeuZ0oSo9+e6/6gcIRur3JneT211DLwrijkFaStzAhY/igqZzUDCH1F4
H25DvVENPeFeB9LWQi64OAuq2eT03QiPEjpryzQoXWns4vX1OS78GUUy9yIcvPbE
qJqlpSKFLdhySB0zg3FMzfbR6Wjx5S4oDOQU0zlrq6cCQH/HPu7czi2oOxqtWVLy
6qh3l3H4siII51xfyLFuOB+nUWJ8ieXiLJsR4mVdZHXNh2QzjDxVoaZQFWulN4dl
WXkOj4Z49VALdA4OSaiLwh5X9tEFY7O7M0zYuh21v2F8oWENc/PxaF5cYWWjrwTx
`protect END_PROTECTED
