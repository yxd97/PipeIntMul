`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHxBML6TJoFvc1z3513GSDAjRvEToAEGrj7F08vrsBS24+bGJEsM/AlUf5jcPbOU
bWp0Sx5In0RoqfC+T2QVjTLg4bTFuup+Ic7ecEIHGJ8lfysdnezx4WDkxKMxM7z+
+oGrtjRetrf/lw7UfBZjIlBPe6xOTQdXX3zDS2XHa9wywRJD//o+jic0Pj2E8hOo
twd01tRfNDJKJSzsP42CPDmLP29zNySFcUVeqqg8C8rst4nypibDHMLL0BVU5adJ
`protect END_PROTECTED
