`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7v7BxJT1KT+3Qg7SUMAgDy436fHrEloIc2eVD9f3EDXV6Azwt7wZdXrEIRdt0pFg
qsHooJs8oGAaFP/OWCuIXDlzasgBXWaQs+2Bcy3SpfFZjlolhV1yMkOrKW98fPCX
4s3dDF3yo4P5Lnedocf5qfeC8TtPKJtVPRn1Qn+/tKrwc7oe/mDsRPbJ4x/y19HU
9nzBCpSyiYoyoIHNK7ZqZ27Y/9X9T9d+H6qJHsQlWFqm+JAUkXou8+Zw5sbqAq3F
2ouvqZLEDhpCii8ofLEzJrZAX/WUwHMz5OxQEv42nzgA5DqBmRZPaHaQblq05g45
CSLzaLwO1AwVrrtaykBeGlOI0iw1VS7Pde/HYU+qPUIz9VcT3UlJ+MJizJUsJ/Sf
pzq/+n0B1bE+uaaERwq4vn/QzwouPoxBMD8Aui8q7TIwloCib1MlVtd/s8oL8Iqt
P8DbHZQTTMimVtZD/HBlWU73H/yP9h6dWRdQgfV6fM3bfKduDTyrfgOXbSZMHm8s
fwJbgjzibMrDYeJfrkCK5KPOlj8bzTd4ZOo7tjbgZp1WY3m8ahRN0inSLrybrU0B
sm6MZ6woFKH0Oto1yybAldheEYOLjZNBoFNIiPA3TJJrew1R6OefgpVKVcw2diFa
lvZOvN6udsgGhuY0jfIL/ZFwVOWtvfdhfu/DGSS+cy6IgRRBf7duL5ib8gzWMbuC
WydadrPhoT4vGf+QGM7g9Harj1862H0H/bV4lq6jFrjxl1MMNLqZyAWsPOYExg4m
TY5Cs/y9ZeCAYl8rbtP3UFP+GDxE1+Mz2B4PFG7fy6ebQM8tUGGjonbnuQgQbkhr
RVWoYk1YgtjP7AlRkcA5w+RossF/ML7eGYh2Jh0opnneStWzrch9MAAtKX8whmSd
TVkgCHJQ+fBRH1CcSXiho369J3rX/A0gaoNw8EsFVFffpviKOz46Ixulfo9fUdsP
iGi5MtvYSaNPb316CoMI46VciCLGNgYV/aRwEIQG6DEeaaLj7NeBpg2HDwFxBbG/
YbIKKjGHilqT3KrdJF/uiqw++/CUEJyCY/X17FIXoU1KWO8qPuZgOj5PE7Pe+X+o
DD+LFoTtIBD1VWdEpmk+xf505PpRyWf2gb5TdWTEFlqwEfUKrdndq/IIEfdb6hWd
hQWhxRn3Mwz1EIaO41LGAxtqEA4bts6sT2xlJpbtACUeQhrO/F4U6yv8wtpQK4dA
c+I2f5Hlr+VN8XuuXOBtgRNl6r7XFZKwIk+u7dPWQeVHAmdfGOOVvk0ENRexIU8g
29bd667Mp35GezMLBL5ad22EYw04gsGEtAOU6XeIRIYe/iy0Nd/Lgm8ukIPPgqna
85ztNO2cGOG8c2eBN7AHYbuRLe6RIZepXcwNHDKAzInsIK0HGdNRmAS9CyMu+dwd
nDNS0rMHLrZKvFpaTE3cT8gXd8Ntzni/hEfXZpUMzMsi8EKVNJsVVlweJo6AgVOG
Z/RavvTfJ3oYbxlGeAnWiljQzfcPPz155p8tXijsyKy0mOzvdtw2KS72ul7v/V1P
IUexe4aDAHzxRSYK37SedwNSQ6JRLybAD7Ce+U1DE3oUk9/GR7tBXBhVuosTA3ZC
2EcfCLY6zOJ3+YHn0mX8GHyvE76Fpora/olsYq3QS4yF5qVMU3Xa1SVz9cLx3gea
647tq+TZHT5ka8UIitkQCJbbih4BR5Eq6rgD9aI8SxdTzqYAoGqGHu+L/BAw35PQ
CVpHG3p5eNrjNTqfyNMnzRyIROPJJDTDjraJlDfZkjAhRJNiv9znkXAeQpwebIcE
rPHqhKruX2P9m0O0joHtBbl062BvVY1zv8vo4ixiuLP3OC/HW+LKN/zKr6T6jElj
yqicgDy3QmrX0HFTjBcA9Dj74d8xXLhq4tgSDKwTTTefkQ27/j3GYFRe+MiTcuo9
cpyAhQjEOPBpwC/NHJV4gSPQZLvIHV2zWWahpX7v1iDMagyPLHRzoQTxiSInGEaS
wD+Fnm8UHwDWaOatwPMPf6kvht3v64mcdZVw+VJ+gWRs7nBAvs4HG67S6M+bltT2
gbGmKrq3nLejm2rL1ggX5f7ulUZ+jDYoKsx9TdtiyGr3EeeIGV/hFykg7UWQgOB0
eq+sK6XxKGWjDAnS3YyL+VcX9D0BQVSdMatRbXTXFzV5RgE6JNPcUmOn1V/l9Vog
ifuyWr29sys5Tfz/m3Pdg+RcsTAkqxD4egr3it9TfSB23m7o3ySHeg4FSLuVMs6H
MbdDUhYYRZyiWVaWkQ6T4chPW4uODsllzlS1d+EXCrIYP3pyVCmgyZbdq/TbwoTY
g74LOZd/SdwpCky9ojiRm6os9MAGyPFPnqRHMf8G5rKNdU46TlNSseOAvZpGhEIj
JDM/qzo9ub/pdRIfDQaqdrnRD8k3qkeWyDsBn1fmw+0mnHjn2lB3Pn+yJLvMDSKa
eKRfGsulJmPz6CTDBYi1hbGG4zblA681Su2hyLo+VoNm2Jg/B411xm11TojK0qW0
hREJOHNJzP1Fv+I0YQNzm6Mqo9i9JkCF/CXsN5bAjzO+W8NBCr2dQVtzrb1kBYOz
smdZ75kBNRj9wX7VyCfNcu6d2NZ5wrZyRZ5Q+p4jj7grwN88C3a+e7XafISa+7Ue
zarc/8ZcSfQ9B4PAFLr4uHjPNc+u6Q+6YvrJm28BGroBnvrezv96aTPESL8YEyIS
I/rvvvB0o6gd9+ofPgooSEtFsJltbdSJcy8ev5kbAPj1itP4sKMs9mH4YP9g7pvT
8hA5rbHNjzOMI/mwwrvBGKoUolAu5BmEWK3WkF48rfHZzhjRohNrMAjzKm/geT7F
6LKRTQJVvxdbMpie0IGG17fhhp+QvYXilq3OA/s0YcdTy05ILBKjAJqjwsT2Lnxu
bdQX1/AHN+x5qg6JQYSnLyU8mpWd6CKL73UOrjetaNaH6NJhc80JV/wzDPrJlpIq
VucIvZ6lIbEkyWy883H+a+htoLktoyT2VRgcesKZb45qlUXVspOAiLjSksA++aAZ
/NE0as3jPs5cJKvYZrbWCxtTgFfruXdIorZGVHJKZ9vzvkB5l4olSvcrWvyFGvK5
Zv/vFEglRIpGBHs4FT7GrVQH2OrjbeH5o9ISjcRSesuB4omtIVY8OlKsfHT+mylv
6l73HP6dqZJ121JalB1kW7ZdcXTDzaa/0kbE4z4KSGEhmFKQKVDbhYDUCkKE2Kqf
LN5speDbT8Q3Ph807F+JM58mFo1NiGbYhKZW3tq9/uueJwHJe7/W0Du4kp05qTDz
52cnDflgggywJyao+UQ91rxDwO8t25ybOiMm9bb00JcWMU0O7oPwkPZ7qPHkj7T6
kKrg4hxLJt4OZSNIkSJwgl4jZWcwyDcoPC1SjGg7U2NQ5cjCOG8er6UusQKBu1+D
ia6sEvEM3BG9i2O3MM8xd6caEErEW4/a2Jcb331rpgmz143O+Nvjaym1BpMLffHD
VRzEtECfgYgNkkeSg0rVD7KiKOgDMs8ZkaWm4kMcIs1cC6FcfFRbdrvEYSgvVgcw
zqDwqN5bWtOGAIz9NfzOLtuFyimVG0Q2VYhyyTDpI+vv5V1VxRF9zYHEPH0c8Nnt
+lfWH+MTdCstqxLV1PTgPaJ2LkrM3DV+Robbp9Qb9ag0KKoEJ9/kxjb9mSKacyJ9
zECFtvWtRvSlJCkmOGdos7zpREYaVzwhWWrjnIM/tBHjqdV6nxtIK6yfIePgvQ02
6gNk+VW/7frrHmocX/yH9y4hCfJPbtB3+VvU2FdEzSpVXAtvBrqh2fKvqQCobvYa
p+J/p/5vvht1DHvEEIBEkjS3mJm/NnXNWDdkNwpTNJehlpLNUGAGtxkNaDq00Yji
ayiZ3zM9P3wtQjn7aGOcJLfyC4q7BoJNPCNajV9IAb1kOpTujuIX4w7Hd8ykGxY1
EjiH5VwGBIUpeXLyHJ7YiYJsMAVOd2Nur1gToKNmTrhZxOxPEpQHWJGcKRTfAqiJ
oCOQGBLimkp98LuUT9YpL098ofJLmqnlg7jfQyJrrdkYFL73Aa6/xpz2DVOC009/
40RZcZmO6FHG46ZoXnhgt8y07JDKRXBucmDsb7HVpqmhYqIG+N+kWS5w4C3hg80U
qGUBLgheA2Wy4hfd+ua/CXeLCghek1p8nxj5gYw1/cVXsHBVDfeezNbZtlxO1d+W
JhJJrESbzsNvHpGFZc61Y+W5ibv3jGIYvM7J/dlKS+ZjQrLudDqAU5TA9Do6ZN6r
gofWfFMejLZwGdW9d49fE58gZgZGZGswgaBoq+YE40k5m3lFsU1YUs35ofn3w/zH
1jVvBeNTfSF3qBdT9mqbTy9/Sz/+OQxtWLRI6A/oDBuAvnnDjDr1vt22IaHW4Cf3
4r3nXh9VqJ8Wq3kedvmNK93RRyKZ+TRKQnV7FjnM72o6Afbc58E9WLsPulNjB+OA
wPE1XC+UGd/Bhc7R6f2mPIUlu4VUUoC+ExvmU9+mAiqj9n2Gg3s4i5XsOUf0HQGN
/JuWkOKE6RZV43i9YYQsGdiI0JXLPftu7nMd+V/xuIwW7unfguyyz/KbD6NOjvzL
SUO52FX5mXyiGFXSlOlUpmZiRwwmefguk0E1lVGAq6KYqN9dG3cIBFJRPrJFKJRB
p8SFcMnRF3iI0Fy2o54fG9Ob5b3ONIaNdmj/VNe7sRhBNhhYYXbBAPnwQk9h50Id
QiF+kqi6l7lReQcRUYFiTJQ0CZzdPI2KpT9JXNEqpelWpOgr5O3CDU2jV17rFa2V
dXoQjwSNbjBqkiaCbkl4/WI5XfgylAVWOMTbOh6U5CbwC+I8QcQQyhaK8eGiU8yg
Juhhrq7GrJ0sT1K1VeAO0eIhQw3kco/8zNNYcgFGzgPjhIxNR9q9ZUxW57QlMb2v
j7pJ5gpHGQx/1g1/8Ft5HBtgpoPyx5rIk3P+7AXeonkYPJhpsqlRxAUlktedyeRp
wj2BgFXSCatE85KoJcdpZz4Ui3E+q7rSbYCZg9gP/ghNfhgxgQUQ9NSVgv+2Sc6C
usLoaWDLbGGkz8WXykQF3CuwUGYA9TmvCYHNgohO8xx3mPaVWbdQr9MHckKyg44q
XhWG+LqqyGog10uhRXJdBPi4lGKp/kSAByDz9XgGJ3zdX6P9UVjBUCTWdNPVSrfA
aK41SXYyZp8PtlQMpVJWn4RmAUlQgO/MLU1YRvGvYuy6E3Ght7BL1r1pAediFqpW
udLlF8cvXQB/bWuEQsD8yQ3D7OikVCy7aPXj6a+KmTg2+PK42WXMKDBfEBybnCl8
mRVGjlyqenbvpcL8NP3+wpt3WJ0R0DMs8KAE9HvFF0U4UjxZ67PmDbyYGE2GMGsy
5m6rpk/O39cz0IrBSlxdWoxtvo0xc1IfXVPPOvYG/AtF6LCU54n40+j6LB+EOhdS
e86svuvHgEfbrBnRnUxwIjZgqquYVOAeWiKICzB4QQqoENkssPSr6VTAyv5L4//7
wYA84jUl8fIaAnyQPiKZZs8oRENnTsJJFBri72jMrSWhllr6WtlmFiABpty3r9bY
eAlPDoLD4uhn4zRMSgTj/vMCVrWjDOqdLosPhxhPkC2D3Wx77bWwXdvPt1uFi3iD
Vyo7k58EyOZb0E/Qo/oGJxb1OZy7ypawFJjVA2VXZRsQwDYdyBtOvl2kxo1vC9df
eh6dY9KRLFL1ypwX4F8O7LCFY6FoRhYm/Ecmg4SExsNXseKryIMx6RefZt2zxv4Z
HCkd8pICVL4gQEgA3Lbgs7/6oMGKVMJfTU/pPGKM1g7npkUJJIyJpVkuNSwS1uBo
1pDc0KNpeQGiLc/w+Tpeb5ibL40DuysnCF0NYJWH4mrOhmG3ibnd8VspVQv+426B
msLa2B7MRVg++qQmJsN3144NxLafAxpzwkjx79Qrve78mfEBPFfusrHgI+y/F2LZ
8aBC+/qqNV5f197swD65G1DInjDaLlpAT8lpf94O5YcvwGoxeAWUyDx2EYfgDjnW
niAMlgmPMJoNnXFaEBMxDSj/3mqAn0XjIPoFDQUm+EmZ1JLJfrEDnGlqGQfka6Tt
AFv8jvvrWWyuy3T5piSFptuxfw7mseOF6HqF1rZSfzIIjzcDXBy4pj/uBFf97aCH
H9ziRSjhFKapWGIc+yFWulJBaBkREXaqvRdlCJDLDjOl9DKWGi3Z13fgVInP6p5s
z1IZjiZUY5KvGNFTq0iB3CCNyrPMRXy8krTJoLLnSpwoi6RJMm0aTXWRObEDwGzg
kyqEaZybSjdSkc1GUdTPP6xsAUGQRDLsSNyC2/ja46lxd09kbfZgNvl1mdxjMNPn
wr1T0CEYjrV83bwws8CwB7U4pTH9kfFd7RPy6uAw0YEYyWNU+YaZJSR6gg/0ATZT
a6YBDEyOb29FhK/fr/6dQynxRfttPyKJqwkuxAXoelLrfmKhpIxjb8JWdoanWFbO
S76a+7sOVynuEklgQDra5rOiAEqp5eTmXIE2m6S6ExyXlRRnVOBq68QzSCyUfKd1
KYzbHHNW2W47oLuADL4t9BL4OKqRoPKRy4GSjftAHBBQGWpg2zu0OS0a1KCWJq9v
FQfG4FWp+UcmgpIvCKA6FOcLrF3m5bX7oqSvYSNqQKuVARmQOmWwZUAb1sHSLjGx
3Es1LYUDorjZ2f+TcO848kt4F43HBLh2v8lm8yx7CooFGlt4P6Ynw19ZciB9/wjW
b+rwzljG5hJ6zKBFuQoNlfxDN1CKgLoS7jdQ7Y8zapOe4y+xAx4PPhtImATI76lv
vE0sGkzgT0/Q3W+1+iUSq/SJ0qthU3YfSHqCcOHCQhwFiSKcsthQnW7o655SrXnF
w7B6Q3zFA7hWZcJpvdOZ/DTfEEeCcuxWTlvt2b4IuLGA9NmTpK0iR74sW3syRsSo
JwTRDZn2yIdC0hA+3bUfbAs0w1lh12ECF+tSekai/GNr90OljTqFcZnx/GnHH5fM
Uy2h98MHbTRjppDs6ZFjhQl8iK2AJcTn3qrXHEwymv4COUtEJFq6QiwNCrJGvkxd
tjkh6aakoyYYWcWBHJE9T/Iubf+bnDSDyE4CjkUzOIfCM0FOqFwmG8xgt1yDPPhN
7Bf+BVpHsEGpWPVNanz1CRXbuQjdAFpV87FSfjynjmP1hCncM8wX03FgZ4Dty0vg
jX3P3hrlD9I7yyth3gzvq+N0FigZOe2NQ1gjmJv6xPIygMQPiBjih6YPuCcLm5uL
W8hsiOgu0B6hitce9OdMJ4+hN8L8azfeP8yKDyYKgPxFVyioHheP55eNnXP/x2nZ
ESLVg82wEIx3myowhvxiGCzzKq14pu+1aPMgzDPZBidMbxuztt3bbaEp9NBcP7Ty
O3P0qJ4X3lfrk5JSDsYQuUujXGy6O2XpFGX1GATNxJV+0g8N5esmgHc8ZJNWjt1A
NAhomLfHLF30UpRABvyKBvKs6P5pMeibWt9FDeSkG95Zi0jBB2GmOV1rHs6EEcVG
byFmcqaGAvF7Scn9si8Ev0oX/QNrKoqGGKw+ZQ3VCM7zPMWmqX4XjEo3LzCPBqqX
Sz5c/LVv0Rai6A/IBnjq10fCj6K1Zb2OcNbdn9EE5T7EjHFYxXxmVTvKLI8j9X3U
ir/DP1J9qS2RRf23UtGepuIi4Z9j2HqgECIOQG5kMeohfr9uF2HeW0AANxz1pGrp
CLQtJw1I0ZiuaFOQ1/6/2Jwbi2GbtjmHk0o03tDj3dR47Qej6ARFrSZmj3pzrqza
M6N6C54/Eczhv+6vaXJi5Amh8fJujK6VzFNkZ8v2ZlFM/YcoVD5LgDXaLO6EGN8o
/fmgjaTchuwyZyeHlLwnhArXx4B/GDy1qvG1oOSwyJIkkenUGfeTX16f8zxaNydr
iXfHM9XuibFdcEwudskF7YlZ3rmnYubTSuT+XzJG2JNKkQa0j/bhqAe3KaY2POM4
1PxSFiO/g9p3yMRk4Zve6jbtYVis9UfXr393sShGPn61dULfVKVR+i/XGdoSV4//
SzPJVGD+qSvnuGDtXbKsENyt7BQYoMjozhWPIYYD9Rt+cTz057HtStwu/j85vd5+
hl4eZOJS9hGJ+UenAYLZMLjNU6SV6mtOvcBca8rbJAvZ/Oc0vY3jN/AR+Z/aFd+e
9lRstVnoeUzdrUmU51OL39fLOs0Qo3P4tu6LsjsOaMd4ANaOz+A9TJ1WpaSBdiJI
hj58YyEmydBLdMsoMzXI3S9r4xf88qe3chwjwL7tIIOs7CXqW7VM8eFN0Yy1Wkki
xk1jx5EBmfsGu7idCO68TM+6MMamHf4LhggvpCt3xVXYgKxuVymgrYm4dGnQoNKe
1omr7XnXQYaOyf0kWTmJk3UXybDcL6DiWSGzmtYKOLSAu6DBAjnVQR0FZWfpLCVO
vAda48MN7NEehuXp2zqaPqCPJo4xxc+L15qTTz/rc5KVFPvt7zhExf6A+O1ukzm7
ofVs58x2NDz0N8t0XtIO0m1QENL98fNor7FxwVS5s91/yF4ez1oYXC/uHO9/x6A6
8sh4TDRORaEFKlieRRLFH974ZbqC7FoasLDd+lhNnIgO34zNVeXSo51QmfnBL3YT
9McqN96jPbWFSuVKhhlokIzAklzHNXfz2/N9a026q/PNBrMp3TVO2wFcHdIURRSN
ktPNenny+ii76qspH5ONkdReYEAW0Qixt9Kaf18cWsNb/iWT+9lMxtlnymTJqCEq
QgDHGNvYVKWjo7TrBQGjEuVAVJfhpzRIPag8ktrz3pNTMkukJ8UBlmx2OhjaWmay
1VSqsMrw87bOGK1QZ1hs0BA59gl+7vxDcnu8yT94tRRFnGnpNiKlE8e81ttFNNDB
g7NkYDq6pxvANYKfsd6ypj6zS5v1KhJhZdjv+BbM2uk9Bbcak+sK98/YDo/P853X
4+g/ubThy5dZKFOSEHfaRYgcsEjGyTRTMTuQbGZvvG7gIGZsu7QV3ni6aL1ZAr09
DU5d/UDRLFCGkdrYLe9OBQgW3JY/KyZkwSfoOyNCWNZRA0KNgZuioFP5smg7RhgG
K6899mHPG918+tPgZazH2AvGdgoHTnMt3WEqlyzIY3gr3EOoWp1mpG53f6fVc+ZW
m0tMc/IGUnUyBdEIt86xE1pwr3x7V+xe0MUuzagHUI6B8JGFBMfEZjZivE31EHFn
qmqV/WKCDv4akpIZzRq6/M3EhLVuSbPpJbrA0GxSVS9wtCMZtxwNEA5tQ9N2dWPL
qyJalkQegY8xH2NJPRCyXoDn9fF84EIjVjkBbs1mXD10WNcOaEUJAhAHQeFqNTC4
igMOWsAxjOIFzJ+U3lkiJw+yLUOLIEAxk+VuEVEY3r7APE2RZmlbORNx2xvGCtHW
wph2sIULfaPwd3Mva9MNWckbiwQQ0nIRG+FiBLW+N1lGh4UA697hbzflhLmF8HHI
wzBEp2ooDXPR8vUiyIj3e/OWhrt5rv06WSI5NBY6HXdoOxOXpRS0tQSZ566bD7dY
Bk+qKaYMqwaJOfHC3LE5Hz2EPSa+VVX0t9igGcId6+N86ynHZJJj/OnwJXtPTP5P
Ah8d6q5aUPZnQuyuCBIFeVlDMn7RI1Vc64hX9fJv+v6vbRjkFtSRgX0Fz20S9wgh
yyw4HceRuOODe7V3/Z9VMmWCiKzbak0YmRtP3pIGBF7RJ/dYuZdBeY6lxXKEKJJR
JQ6+kFxC4rC5z6HbZrlA8ReI8We1t94y9qx9kz5EIziCK1zfMQk0K2tW/N+SuOqW
mPAaC0xISWp1h3oX/t9FLM9ZyeFcbOJ9aev9fHQqYqpgbkN2/1m/bDauCJ63+J/C
DJQjFa+1aXIWrLGJ+295F+fua9M78Onc+yqmHzAuF1w7iszKBFwfl5l5PRAZHW9O
z/D0Fi877xkRXUS8LAcom4isTwrjtT4KHGf6GbIXp48s9QB/gG1GuEaTvtfLSXlz
FGtFW+F7X+vxZgq5NbgmgDwppDpAQ8YpHnnDT3NI/AlIHz7mTzhrgpa+SlB7Dzif
qrq9KQBmQOIgGLs25QT6svGQlW8YOIgo0htXbbnUBX2j4C5EYBXxcm61I5vUwjN/
AOnBfv9LYAh5+9PnYNAmwI963lGAptWwsBf2HdRjW0q5FLgmpEyvUFOwaK7/eBaU
D1IvHdki2oxLqr2y218SB7+wPC7Epziej7nZhIW3IBIAzueIOubGksO1+2yp185j
kDRqdIuS9XvYEpRqRwLIZkeCx0AGKq+vJ/91P5EVXO2ZZKVdTOzFi7ZGcV4+VZvB
mge/nLX4oc58OpTA3cYkNk+r7IyIWYLmUcKf244Wzdp0gl0g7Ht9BVN2hBxL/Vu7
GHMmajCFlauIOmzDHgaWgp76ksulTKwrTHJ+6EQpXBO9X40N1Cpk7gwVpLaciSUq
x6Nzb6Sf1P+ffmXNAxp2Kuoebf/JGEeJc1clBzH4B6Gaog34nyaKZ6tMDM/hp3Ro
bs/F9G+KBznwAq5m229seVLAmngVBKIDnt5HwwjUwtUKcQOsWEPG+KfuapsGh05V
ddEBanRgpRYH4RtWZUaus375aEnnucQ+WuGdcEtASTleYmrqnXvPIPevSstRqmdy
RC3eEdA7sSJC96sC5pm3JTU/glcC2bw+xfFsRQkIW4JIUaIO0WXB+TJCHR+Uo11h
Awp6/o5jo/Oh8cyV+tripcNfqgZ3ZT3mtARSNTKCBiUrw34ItpLThplxkDbmEOLu
BlINzDMQXnuW6qiKg2UpQdTCmDFOF1p+di5KhvJhz+Lf44ZUXw9UULAGYMDx7MT6
BAMPhg9Ie7UlylmuxgHLVLfuyrPnNryCVqXBTs/ao6Ts/owhuIWaMSYUm5qpZNMN
fcUSoWz9YUnS8g6zS98PaZdbj9saB8UX19sbuRDC9CpOv6HjD0nJgtGMsAo8Cc8l
SgixWB5bnpyZxmtsqEM40zMXyjATqwCDxOx656Zj9BuAPZMKtWL9bxlEpXYo4A7R
Rd8fEaYl/dBItqgAo5gCtxNZd/k4w4ec9xYVTFzjPnSxiV0nfqJwbHebcxFF8TZC
MuvJ/d0AoMAkhQpGmBDLSOwgm4n0zBtUYjSs8CsENgXct+nkWFwNQg0t/Eb6Z68Y
rJlnkjBcjiQaCAOD1v/qKzlzFsxSoLMhsYb263Z+j1nfq5410MHDH0FHec+4RjyX
WrNeaFNbATz+w16j5ETMQixtkrMPzSZdAUZAx/PikzpKCEaCwyZwsp6/Zs4YXhMU
tcOykllM3julAFVlVnBWqAyOGgeFyWQ4Hh8SDCa3mAsJ9eLf9s/sQGLO7IPBYJY8
xMhfFsnpMsEMgc/+6JUS1O8RXQ0B/hu7xrHpvHJmjMlkPwEg3HopN5ALkW02ZQhE
3mnZnb4aXV5W3whPG+TT6RsWXLQk7JaLSpnydPcyKL0HVFy9278cd8WMrCk/9/ju
m6xGkc5FPOn2Z8Ck1IgAbvDkcRiqn9xRP/0gmvJJFibXV/13/bkU0Sl7EidDNAVV
ThGOWzndo7TBNHx/A38HGU34AofMsgUf4R3olacrmt7hyWzDO6SRtMBFMYBjhmsH
v8IfLj8uSuJll1mnggdBSkVsYig4OHii1XZ1GXYk18GVjrrc6BIlIeP1xdYm35HP
mn3hKqQK/3T5OvbNbrxddhaot5LiMBVIiMnwF91mZXwx+x4ZNwN1j5DJFzvdVmI/
0S5Fpbk2gdicohdqNEPKWe1gyUj1E6m94gX0xe0uob5yMK+58o0QQ5KsQV1odSyQ
ctcUZWc8jxtXOTJp776Do0Eu8D9usJHAnMULh4MA5IC8eyHegfha0D+uDLRfN7xN
KttmXd+Mr0lGhIQxlMmbrQJk0y2THjpIcusuKS+qLfB7pZ59ne0JuDM05G38xk8q
8Dy2Sh1z6715iB40ZUATu++I8b3Jc6gJChDpWuGg+IALrUiMqrdbSmAlmzbtXvrA
IZ5IxE1/wxwTTy7Elb2HNxXloAppFxt7Ny/+fpPZqqeQBINxyTOIFDvQHzaMj17h
v1lzz60L6QXQGDzY0NvLZ7YDzuvK1JHWHwxYC/kniqEKn2L5e9O4w7FCFTb4sx0v
CnKhRCFjkTfu1pBiAf6MNVGa79JST8o4eZiaXm3oCTDt71n4V6dnsOg7964L4IuS
ewfIknRammVMIwHdVH23y+FWw/JWwfKZZdv3y+LjiqPVYWlRBjpKFnwG5pU9JwrD
lcD4PkWe5N14MyIt4r6smtWta3E96eoz0ai09OkVTOIyn74R570hS0PUiyAiuwMe
OIU1MgFipJw++p3f/5iFMTPJZRYpH7bHX9iouSkWNNTOEJ3NV7FlpXjHiBHcHo/c
M3GFSYkyqQv6295UAqWBHTlNjH+2bApb/urOYIdj+s0rIetVjud3RUYx/BWCKi9k
ttGsKG0YUT6vxp/lFxakHTo6F3Wh68oms5gOiNorTAWaCvxx4NW+JKdrMM/1fYFV
lTRSaRKJ0gU8l4oe5Rreh7WmMopY0EGYEXc3hUjaHnAQsvn5J9GvW9WFBmjyfRB4
AATqy27XrhP6d5ws9l9NRjrYBmb0p7sl8ebDxhNsdHq0f7wXT6QtNzgpoq2Iq/gs
pQ0Ww1BGBVWJg/i7hQPnSGhBlasP7kiSMIxTWmhNWL5QASoKAPZVZJRLOvYAXHGS
TG+OnExOrn+ta1O1lu7B4TBkWpJnO4mJj3e8q2GC9Ncijb8Zc+xXSJNJX4A+8dli
O5fVcZhOQrBQ2AbnO9J9ZPLDQ74hYgWGb4wS3J18NrwzgrIqEbOrvjMVyu2Kt0Bf
Z6eYC/+QCNsvntK7RyEM2qpLYyCLtvFLZQfVToGNUC6VWd6pH6x03F+DYapyHHSS
LJnHz3uvCsINFj8X1UUHjKPiEF9HzU0IGT8K5QACe1vTVbG8wHYnQUWJPZMELFIa
f/auCgBIHl1z+WrE1HKgZlPSBGhmiKlT5sYDkNi+g3G6NaeIs3rcetdgi2bGQnRw
/7pb9kBjlGHOHWR5Q4Mda1iwbZRSFz8JYPrkKznOO09BnY6NrASHuE8Lw8q7YT/M
rnAUxAuwxvvY2WufVZe31CBBC+iTDc6kMHGrPl9A5b2ENsxOB4PQZ7yaBD4OztXT
qC9XH9CeMR4fbKbpxXfwiVGTp26aYKjAG008lwr75Cdpgo9LcJrCcMT37wl0OKv4
LuFVPwSd6S0NQqDOe5+YRDkOuv9opzoRRCRXsn439eFHtB/QNNQOKqpadIDknu2S
y9Lym2s23Du9JiVUylgoTSOQTi90wXWISeC93hB6P7Uid+guouk00XllAdC/Mv4h
l/HCxh7wO5/SrV4bfwZDFJMAvD/HzcpcHrpYbhtVV/9Ly+eJh64Bt+f0D/aLBtsO
wW3H/TgZLbIQ6PI9u8YaV5aD7SJrnqbOrGfd9YBbIU8SXZFK5EexP1bf3mBD96TG
1pLADYnfRT3w/LnYJS6MI2Rm/mjfz0u2GoYn3dSTH/xafgce13YIsssuq1VpDM1h
t0rvgP9LaoFlnyCBsupdosyuqytqzACNOLpo9pyTRXeYWmcFNeTc89W5qLbm+KSn
l3sEnKi1hbiw1MvNrGcL/unjQIrkC+mEus3qKvqpHtHPox1omvkCaKcb30B2tpSv
W1LBjIuwM2ahqCTW0qG0Iv/t0cpLf/IEIewbwSFfdxhhZOxYs+MPRiVojlC9PD1l
3smyQYP6jGrmU9/FYZMHSaaq4KmVxz+ZUq8G8bF2k6sU6UO9HFJxO6Yr6FnSu9vZ
OG1BJRenMxtvw0clTfYVxSfn+KDzvabVFtsiAK4bBMjBUEN9EktAThQOPwAKSL40
zp0UzPSQvQ9O09/ocZk7FQiBhp4F4zrn/x8c4ebaVCERZVEDAeDUY6RkWS+LJLDR
iesSgxHK7oITyTvIsLlwZxaEOKOu68Z1oxkGXdcPQ2xLpskT6IlYQfk0nVV2tf5P
PuejYa9+jhRUqGGBzKV+R9a2aa93fHTZfKTFCpp1DTPL0AOy2Fso7w+EAl83nQ34
/S5cdQU3HHbHz8Wq4ZRnZM/CUtF/ctsURH1bi45LYW7pRMLSh6C/SawzG2LN2hyZ
0nncTXGKS39aKetNSHGScfgdKTFbjFuJKHcTv3aJaWZ0DGzF99l/2kKbJqDWeIzn
/sRrjJzhQXVPAT+2UyW9ZweibTF34WouZksaQZgRIOgcoW74VnDB6+hmXpbnuN9X
5Rsvmx2Mx+pwduJc334GBugHoKk6ZU2VeN9+/6EQZ1ZE6jTHIX4DRCxWTbvhqb7F
AlYriizaD1ICz5N8NORJ16q5xRNUFODLZQ72qydAMpKU6Myx+jQrurSuPJzNyVY4
n4TYo4T39MB1uOipWSCRz1KVvXtol+j+/UsZ7OC7qN/PAk+kYxWZfCzwcP4opQdV
SdL6LM391lhMza+n/NWsQwljHcDbTm3aQkYEloSbbKGfY2I/eO/cQCcT8a0GvbOz
0fpYKl1941jgBPiydeCEkFouGygLxUox5ZHzpFSsB9GyVQReha9eATzn/ZOJG5Ku
o+5R9m+wB8V/5XqI00JlnrYr810l37VOfqf+XUfE1giENBQX2/jqzZ0+525KwN4L
cxdZbtJOy6xQdUeAPysajYe8OyrkwOMDIxHAgWw/O+F0ebJENilLhYfi3u6igjL8
NfwdXEx4etDdfcUeuE7slK1hTt9Q2vu8icnreEGo1NF/qshu1kZCcsFSfC1Kt7Qo
caGAMFPaKIXAGo9ONKAtKvdqXpZ0YGulKUEFxBhXwZhulvR97fwnbtyAkdhiq9vw
Q5k1+fQKASdn6KBS6aX5zCq0CPB3y7uJz/Lz2Klj0lzfRJRgA64bMIlXkTvaEMQL
d6gT7YWFmASUIoRItdaNWI0XMIDaYmfJUWkRXoMpKwnnlaBvf32wb0SSR8o5pydr
ZvCiqtvVifpKfiyq4xvAczuIEn17dox1GBcDlvBm/3upJ77LRUM0zVqNM/pDeQcH
BAmYCdT3srGSvybpaysYrsj9ls+8dIvwILWeThKWuddsAIbHkiUCfz60q9rlue1F
rb4LvHNjB1u1Wyycg56oSpN/xDYyGOYbDxV9StRGhALmmOG4L+A+S0XN3k74g+K6
7mrxj6dpZqWp4GQ+Vseogok+wUlpg6nDeeDIy1S6+72//wGQMHH3lvu9LqrZvOxb
yszYFAP9uFl/1YSYofJcD4dChceV6RPV+lSEeQrLs0O7FeCPxZQ/LHQVatQI3El/
aVj4AcQbeariliNnmvvCM0Q2+b9zRc0qtAvjKtXEjQnTTG25zG0bfSHwKMCz4T81
QSLkAqH8/aXBnpNezhf6lfXpkDeHCn+4mzQXzaFDDwEm/vKJCA5G+E6RkqlOxWD6
+QFt87tAZgx0TNiAl1PmPrBlyq9WbZdkmqoR7MUGA484cmsKzLF02VYcQEUGopg3
XhL+SrNOZSZz07g0dixPfoLl0aLiXDWp3Q/+ordNwHX/BKKhnXV2kmUIRK5ViKnf
xg5i4tKcC+uClQd97MSdLJ3HG/K+z+G/atdzDBXtSh+gphpxVd0ITzunL3G6aB00
rAe4Vi7jr9bJ3Y9zd3dm0FwNM04JOb+TPVk4T7YW5codTGo+B7LWGmRt4w+59clc
2+OkqNovbul6CdFFcoazAT8KkvKvrpnfBas1qQAAgnLGj4hfq7gnCqDwTjzgmhkQ
Opv5/t3uF5MksDWRBiOKWNuwY7ypo7bdmt2OZxoHkPJkFGJETTILPriipyF0ZULk
x/N6vJE/igpg8wvk4PJdp5kSGvDSGmpeWHI5sMP0+lcUcNgBg9mv1TeT/hhmAuwS
7aNKkvav3rPuknguYboLkSrqlZVO/giCOnYjPKC03sv5TZTIXm33wofVWLVmfRIH
f/QxLhucU+E66JH+09hbc/C6NaiUV8Oq7WXopGFCId/loHQeranHMVmlT4JgVUpy
5mpHFKwFq1yUtGkcBhg1RzI26J4N2pYmZq4fJ35LNMXx5TVJ11UI0Iv/XwIJOSAw
AfEtgYkTar9/T9Kc3rLKDYoVAwJ7BPON71tVALohBz6MqEzOG7C6irwZC6KsARIo
YA478sCPlDx0pUljYyUynjvQZ4H/vqs5sPskAxJztIX7J4SilsHofBiFIpePVA7T
tYLuQ3fs5teIEQjlE1B56/5SR2rWovEUd/oJkACrBsXWKHXrZAfXBT1nl+c97OCo
n3bQcX734hBoTC/bFM2RyzO7mwURIKdsSjycCoIquhSInLUbX1kKNoI0J+/6DkAd
hLUM2x81l1mh5dApBnaJMqa/1+NL1qvtsTppmgNSkNA/a9ksg90A4UsBIBSlHPR5
ciPFYTMki09ld55VXxR8mdnAgbXKGATx6D8c4ZoLNyFIGGsfzYfq+L5xFX3T6obJ
Hoe/lIsKvuJbgX9q5uCuxaShKvcM1Xxm5HWE1S7M4xSA2UCA+1sXLfDSHHHeZr7d
AbmpmCw0SoRm287FEAVJBzAtPxVlHUUVVPhxag2KH47Mwr9ncW9GJSMmIPi99zzP
X3Fo6C9qmThp9jsg4mUUzRxhq7lOD224Mwjcas2rOXevJ8A0PHwuxRhYijRPYQip
gM1J/oRMiAL5rY8OhHDyLOhy4s/BwE6muo4D93mBTf/kbr1Ltsg/bZZmXfW4KO8l
j9fDcXKJWGwg5fd0zzbf0dcfklc7iF42m3hn/pRryBHkEG9yPqz/2WfoMtxLNb0R
gCCRlUDNNke5d8DIYlaNHh3tijQunCf6ZopFte5qLTC06ww/YAhMti0U+mY2J3CH
P7GkB7d+LtzQEYQirh5vlzNO4dYs1fe6JCyoH96nzLaFgk1WYtLKSSDEFwzP32nj
bXPfXAtCuqnlifup51+XMm1p1e59PSQhlYpB0JlJr2oTGZCOIFW/fj0v7F3n27gB
qtH2tl55z7YS4b0vv3wKazJIpHByg3Uyh1reTDpA8/kNCGVwXW4mHwb0qEaLnZbR
vGY1HML+rzY5UCwoQO5o/1vVEiUTyoYoveRntip9kgsVyRa50bnTavbh8sEsRjRl
eZWfZyecpcbirn2gaQ9Tzd24CGnxxJJbWGIlBn4UsZRT1935vKLF7lcU/7qh0BzB
vP98IeHuLthzLYUYNpq1CjS/0FSCziXWfKZT8zb25aOePIxJjhtJpJ7GwVNyUW6d
Eq5/wzcXzUpLGZrDkMSOfeimBLHNqevXOeXWUXnfr0IN3coHWKkI87f97hHGZx8R
hEsgJe+LYQG7rqolU49OztSX2BqILZmVX/4InA8dK7EqDrD9kR7rZdORgBpUoC9L
RmoRAb2jOAzWzk5C0upMG/AUBZFlh7S0rSsZehKYCZbhwN7m7x4p5xNxCr0Rm50L
oywGiu2q/F5rGaITj95GL9fdEg3NSBUCI2FrlaqL8aVvxy/3RfyThChsjifUoOGW
AiIVhthkB4yjyRSHdx7bKYxG5blq4ZWz9WdmpjOhdYTo3btCqjI3dwuhT5y15i6t
z+ggN1euqlziChyyNESyif1I04wgz0nKIPx9pJshWKbAWw6fRPNKIhAgTAAI4sYe
LsM5fXZg05DrGcDTxTQF7FUJCN4QPUYKcgZ9JbvRGv1Yk3DaPPD6KkK8yInwBAMW
iXv7kKi06FXJFPQXYR6waagw6mhrvtstX30RphObNmGvoePBYmxibJG6qqQ/rErh
7q8X8tbXwv7xK4MxeFTH7+LWcXk5jxDbRNYrdeYzRgfu9ZPmpUlEd3e4tdzqF6qq
DdvJ/Wi7yXxwyjZPXEpQA34KE5vUVAH5mZRZaHbm3lfHGVcbtqFPChwNgjFv6gRK
m6WubdpIYZJ/8lDMqeBPbNzrypzLnn16gxVKZS5dxlUp2vx0goWjY8tO6qex/Q7T
ZTXzJ4vPZnu0ZT6cm5RUgM2ljHHJg+UTJ2mEXryFuJgEfjgDvekKy7jZ+lLClzFG
Ke1mKwpC2xl5GdDiaN6Ao9XdC4hPt/aZ53HN0LRO0WLBJollASJ/jYWo9CN48sjX
mtp/u9P6+V8SG9KaiWvvQW9jke67Q966nqfO7CnXUkzgm5udC+W1xFHs23bro0zS
Wc6PL0a4ndejYMrNQlbI+57C2WmgGUqWgjBn1IrA1nFmrVj6r+jOqeyJeuZ/FDs2
PzGQe7zcQTEHQBsIvlBooPjWtiOemOSNsXOXEBtLFkSFHtZvE42PZKQgSkXEm7As
uQ8SmreFUm8h5/MPY+t50wzItz6AFJspMGEEFjzT2lGm1hIJbrBYyHL5MCa9ZG1c
+IzK1zN5B5BHVFp5HlsGhlY/Z68OwEzb1EjamByRllg72i8PWp3HGMzLQV0mqocD
51zRmvwmOFNiEbYLQOugI+I5DDaXvbpHASRxTaaH9vGIdHe5gNXB819bf24fZxoa
CI6FIoJL8Bt2etagqtD94yCFwUfyhXvTenRJB8fFGuer4tZRZZR9caGxHPH/IDxA
tCWaFax4PUVhHHvt82P1PHk30iqyU9SNpX0K4c3iJTK0+z/wShHcdNOjSjqQ8f1p
BOQaci7yxDPPXGZH62IOmeBcDrLk/3Dg6yHXE6hZcKQj0Gjq0/Q6QMV9c02J9XL/
ZGZIMmHkTFirs9mtSAS5NiVw1iNc+Vdtpydpold/h9JJFOOOuK5bKrQNFzUkwyfo
724IUbWW3266Q4AQkFxC8QmijsltNnFvEEcQ8+gkaT/rBk/ZCw/9cOjyw/UHvbkH
KmuvwAGSFv5XEE8rGhdJ72JAt/W2Puhzxae+eJ4Uf+RmYchMjpt79A75xEPNuAXz
yq0VfB8byro40J9GJmREqCUEkrk+VFi/uxoJ4PllhHkTuVe2leDRVHy4QjeUpaeU
UwEV15q/TzgtcWiE4oG18JVflxqUlpLXqmGBODrNVQLG896K+gGpCIglGlrwojZf
kgvQN2PgCyG7vHr22tII5dlzA8HpKfeGINRcxgBsFJDDKfn+cuyZ9UtRhxt+cOt9
0zzvXKBK2K8yz2r19nQAupVtWYSejUzWZOxynVtfFWc0WmCFA31dUmUMLVaRNFo5
Ro3N7xnqpsBtdZ8xyF+stBWl+3ID8pvYAjMd3f5HgnZAwBs91eAzDakZqB2SXJ8N
no/w9g6F3VUBxI4l0YPOhoh6uDPmFxjxZtoq7qkGYWD6jCnCFgd3bZeZsO1/MJZ/
BkrTcaONi12Rb7KQ4RVL5os+nwyPNdaUT0VQOBl+HbN8QGlz5yLEeRFILx4UlwCT
7nKDoh6KmtpIF5BKjySfyXs8a0Ddj5oxmb+pXAydJJ/uKu3HDrNJVlZy3MnK/0l1
EVrMnZqPqQohPxOVYn8/pPt0BtGTZONNCk/1A+Uwp+qyg7R8h3GJPrV5mAr2kGRc
E2Uu7ZppWGpSSGwQ2h0Jq/Q96PuwDC9R+Cbh8aeBTuB4k4nuldNJFoqpsVJXE1uX
17It7lgqFXo39cnv2A49WKCqYLtdR6a/lsY+wCDP0ADDTo36zTLC93xyFs8/kak7
ijSZ+wb1pUs7Nfpgx+YuuTL/oz6ddcmWof1m8Z/vvoqPZFz3Rc4koDmg9teBdlLs
UV5D3KdQHgGDSxw0bEW6Sqf1YwdSxVpMDh+zLPi4tkikV5s7JQM0KChr403Z79tG
zYPbMf3efmZwcMVNE3D/greITpYACG4F51oRj0OZZXXByclUmzVGtsZ3NGXtWvRh
Ujeu45raATsdyjVlFNGilYjYfzPSybNKkn9hMSmDQZfEUSn/QTI8vENGdFLP4JnH
7MmMgwtLMsb5MJZHT/y7XADOZYb5e8XsvrnUF7mfehxUYVhSgs9oSAZ+uDTKSqHB
q1zFT1nF3UKDwjXnwJ75rKKajA8b/x3boRg6nEhsU8nEs/FpAma2yjXZuMjJlkDc
b2I2HRYjLAzlWjcECI14yfZPpjnjs7NHQtgi1rWvSGL3KVma07m/5rNilFOkoo/q
AvaTq68NHSL5+Rqi7Qvm3grKe68e2hbiZkEN7sfd7Wvj8wfK9ldRYKx32Q3fZ60m
5ZQNPjBJqeCTJ5kLPVgjzqGgOTCH5bybOSiVHv+wRYVW6B30lKIEcnzwE8ethEjq
kb19gGmR5VAA/mIlSnrHi3Lapz9AeV6vIuyO7mnE9MxPHlvVi8SyhC51eHkeCw4J
ysjwQtcbXRAD6tkM4ndCwPRoxNapr6sW3GMXF6kMeDCZglsaioOtcPMT/ZVuNDnN
Tzimu4ll5NCFOXWwH3yYGcG0rOytWSjSEA98iYzWI5eJ7YrbgW++jX3ktwSGVYU2
rD6ghErBUcx6Z5e94vlEOTE8RczCipoiSr+u6GhAxoA3JTEUGxukHvIOUrR35LU/
sbW2Ngq77C/lTLuCCjaRN4KoL1svjqzj/xhxl27EoPOnyyQf4RQTlDJHsQuGL8hR
n69FCKE2WW+nHp4hOaJhHiv+i3JedVHLrBPeF6r3CeLvw+Kq8KyQeOJF1/p9OFdE
MCTBI3zxWWaoPoorJBeRfD0qpsvLtsc4JLSvWwnaulu85SUCoaX3nOslI0LTFRqG
PuLdsUxOwgUyvTB+FbrJWlR2oKNybVDj7uerDRd+imNnO+6U6hby1GifRmMio6kV
Va0jxDm7a2ocjvWyCyAUQDjCWA4kffKJjGAgqw4cPG+cYeDeCg4dwN0wNE+VkTh2
+B+vbd0takFZahdZFmS0BVkVD9/Df9wK73cRr/EVjcEFyhwyQb6+DzVkJIgifdld
LaF/xurFT1ev2Ci90MQ3SLgGE+7EDApXoU+bW1y92lRtjz33XeGF80ZxEcWKTKcH
KkMTRyEhmwykI30NdAj8WpmZ96Z5Bh/fQNTaHoDZewl3qYAY07SlzcOF+Orvplbc
oYX2U10oYrIBVguCXg8N+NGrDwQCltOKGNpPdM9/pYkwyE4BaphWGA0z4bqYmQk6
GELQbCaBA+tCcS1u8uj9DbnuFSvj2pyCycrkDEWEaOh3gXEJUdnkTAVUovRiMuwU
LZa+7IraeI5OqGSg1F1wG/xeJMhxJUXEJJQeGNwWRmGZ6sfkOOK9NsLEUA0z0JRG
Jd4KPInnRtoi/4rnvVfBZ/DLjweSZmJ0ek68dtSIyZieQD5MYif2AaIEIH3DENJ0
aiO1zbC4oXko3STtNNf6uziRpvThqDQOAKR60T2JA886SxuqYFCiMpMYlnHN43iZ
Ruq2SQDa6OjM+zJIBAbZTEQRcBt10dMUQQ38clENaGXj//D6FdGo+FEMwnCB0Zm7
mxTDXC9PP82EdLM2WXi2PUxeyZNfB6x/0ZtvitAH4MQVzIz3ZdMnfuv7+yhkWV+E
C0+42XbC/IwIwe3noKPhXiTSkRbraiMXblRkDZPGvapke0+xKeQASoznWbVy0vcz
dSYUrv9NmAl6RpY4Wsr4nApVulMarx94RWznihpjkDrzHp1R0UYkZz2mA/TJ0ywP
kPe0uKZdv4UblY/jALQfMJ0F1iNfnd3QuIzIQlH59qM8wBCT/0ahj9EHwCBElFPF
Oe5xWNdqTx+7PQl5WI9mBaqJ+A9P3gDCK1meegKxKfc8hFl4TRAAPw3NaPmtyVXS
1XqxjlNmptl7hYlp0tfN2nlBWt3SfczPZ3ogX/x0sAbMzzGmavdCrjGTOdx/pkr4
mi9gh3Wfke022c5BipjquHr9RHRXa6Wvk+2mRR8FAfC9Gl9AlOINJLWYLQDOZcbB
PFzKPV1M67V2qRrVjomrBb6q4CVUjvcmLEG/Kw+07Te9xrO6BixszNl0DreE04Jw
YFxJEHVqWEvHdpgDtaISnFeVZzwe1fNHyKyXhFE1ukAt3GYELK9xY5JZIaZ0lyLU
yECIvSuMq4txs579zq1tkOGgyzWnOXQYPSNcxDBrOtUgBS6NHJm0jB79NIUhJWZL
wWup2oh5vmeSMpMZLHNjEiEDrxRoopKY6/zBjBKMc0tjYdUwgQBqhl4O0x04ARC7
0HrGFWdOQh9oKrRAUZq9kfRDnVojcn5ADGKe2TUQonI1D8erMogYUpEl1Z7uQhDy
pT4qFp7TAPbXG0gs0Lu3F7wg4Aqmv3d8FgUTFa/6fngHIdCYW4IRRqVWVBfnlZao
MNdRhov49C8h+FkGckq2FY2jX85KVwbAgX4FUXDt9VoWIwt9Q1ZssslmszsPzAfP
ARsNWDFVE3PNzTRrCjy5agZqiQaAUb/0gyAM7RiCluEFGv0QIo0wk0vsov+iE2aE
wAdL3+cwihwRr/U5mDbXf8ltXftjJ8EyZzl296J9YGnRs/0pi16UXdZO8ESSg22B
eqCWMcUm4xsAIqV3eyNdUL3PYWqum52p6DOdS0sAobIDN1mbZtoXGkAZTUhGXOfS
D6RGRuINYM+kNdHIpAG5yLZuDxRD3eTKfpXImMHTLIcE5xqK9LzNgY/+DSXgoSdg
qw2jD1aLpq62iHXc4O6UvjKeVYzwGd4jqxUBenz92YhGetFSrsP14AY7aGLejIbl
njJHG4WQoMtfjPt6e8NmuJXuT4f8NItSoTk3C1wmiHt1ssrkiNLU+en4L+yWRGfV
ZP1vRzb9i8OID5Pawq9O9yJhDhaY1HqiIz1SZ7WKbhDCf6f4R1/yB5Mi+5gWzCqN
DwQ6WMlFkvbFYcnZ/Vj/DWN1rpxEK2QAIEvm3AyIJyOXu6BcZUa+Y8ZwsMiizKsz
1DAUs7ORSvZ+v91S67BL0lcHxtIc0OyEJ2e+ikZY6GdSYdIklB0To7WGMdCxV90g
oqdIf2Ak8YJAtwXZ9GywrVVPKsS1xjDe8VNp4JkzH+WGN4zQpoJqJYZYwfszvgxG
1ohp2PRB3KKE4scKI3/6Stxt7kRxp1ZfSq+UB93WECVcvwFJSA3A0Sbt8h1CSe4L
XG0EBPEELpMPtHA6a8vJCAvC0tSoGo31iW2PGwU89qmTLGUUbl0wDLq32HNgwLIy
FK/z6nOpwzHT7ljSWpoHzS0KysTR9mma/i5fYnkhEo9HQiVhuhRB4ic55dcLcori
103qSftc1LsAkLPn4FSJzhxuTQDxbI2aTXLkMpp5lxMuxxtgDqAbKGoInic1UVMa
9wehzA1lbLUDWRQ65HCOBi9hdSna4rjSUdljHvsuQvG4j/W/SJtbGOfycND/tF/E
NwNh6cfclBPog/KCi5cu0DxTKluyQZzF93fIQt70O+qvL+URM1JtQ97fnOi4NmJv
qXrBc3PE302RUdABDXatMrSXtxkc5hCLkv5KMs1MpAXQVpSl2ZxOZjZqbtKKO+Sf
GqosIGwHHBrjZiV0KZHSnHaB/03FRYvFKfu5uO5Ne9B523n/WPQDL93NDlz1CjIL
1Y0RFwxqRv+FVG98VoRdp1DdeMRsP1mHO15AN6mMeeKUeDsmxLRoCp+yUNWvYaJx
X5JUEgD01GLkIkraxBa8jUu4FMmS6rWdwHBxYXJce+Pn4nKnfahMIe9ZzyRSlRGp
LVPJnPXUoqTm6FF0QFvG7GjxiQrh9rDcZOMtR4T3yQqG9F85gv+ngEeKJ5UGN9mm
87jGgaku6NP1bWC5O5C99l/KZg0DmbFWORRyo8VPKBzSZpPfZl+63fLVX9VAgSJO
7UA3SULgRZ7Syo2yKa+T1Sn/WdVQcF+AFbUvjit/HeWC09FwQJLH1x5HMyJi8vlq
rY1r3WaIxpllSTtIcLkfEo5Acy0UojrVdYUEbjsEu6M08oa5sOKU9l83smx2ivDS
AeaZ1ZXG6/Iw7uWzY19+JiavhvVnAjXlv4Rs2n+Hik4IfRMaSAso6Hy8/sGlZKT6
ThGyLN9ho02px0g8Q4xFuAWCb9McvRCYldRj3nCv06HnFeMA7inJtxnAojdR5pqN
plaxIdl/iqXXZDaVHfDm8xAVx5jyWz0Ap63feXCfPY5UQGEbBSTPgo/A5nTXPh/Z
UuH+tEYBz5w64scD1S786vchi4Ch7PQc0WoSEZeIVdWx9KYl1UR9Tdse/CrM74XC
oosOExoc6xA9fNiP5cEPWr1hZND6k9idjZBSw/ej6RBZkziXgeSqpdWRED/QKNCk
5tHVlkK3ZmCZpp3sazevhmoWs+WFTOq1ph/S9s5XFTh38ierumuG92by6H51UGUy
Sa8BSVhkdWXm8NQ0DgK4SJZ+FFoN8VxLj5YH1VS+Qlw+yWM0hELH7HWwAKfRB1UH
Sq+YAc3FzwOcV3/E6LGm64E7sQ3P7B95QEPhSaytsgQr3V9rb0JIThHxXipC6R4R
au0nP7IWIQLqrfOjqf8UNpcbzgs5G+twz0ombL4IfpXJ8sNFHg0K3Ne1RoY0R2H+
u8yL7vy4pjiRkKn5w3ztiyspdSalXA4EzWlUSBt/3HW4Ahviiw8BXR6RJFjLr4DC
MChvM5T2gtCbzJHdiUR2Xo6dljKpVxE3aGCxw9qOcF1gb//bAh1bGy267Ale5o6/
ecyjY48sEE9SyKpkqLBfdcP5HpJq5kREniB2whc1mgtSmB7+Gnp4vbUWwCtHb6Tl
24N8Hg3JdiqKKojzjKxwcIi5ZluqWV6wDQxBBlJkBh/BvUyOLur3xp3niVwE6v4N
39o0nyqLyzV3SqFhoWqVq4FNuzB9FtEvNYt6yKxkFHn8IuoYUT70CYTHtgo70wb+
ag0PEIpJWGXzXQxlsCbgW62kPQSf9FA6QwZemS0cjks68Vbj1Kh7uIYbDHdEsD1A
9X88kuPVEoHqhAzRxtRG1mw+CSFpm/h1VWGu/1O9ZkUmWMP996O2QRUQ3vPfSxKD
K0rCMMImHx/y1ypNCnFRPvJLVYpfkEiwgQV5K3Y4p41nhOiQaDNNq34yOPXKecQw
wUdwkWRut6c51abRojptzWaCvTkYVN4xbfxuPxSB+khyxclnaoMFgEYtJ/4UQ4Dk
JoclDs+H6CXuDLOLuUX8NTOFeV1xpev4VxPP+3b9DEehZ3e3K5lmWFnGMoDIJvGZ
wSwt/onWVdGoZd9qpF/AF4unc1v6x6ohSLisMjzimYFZEfOJDdcWiK5qNYVsVoT1
7V560bGvwCGQg0uEUmbQ7UkzGt+ctF6JM/ESJBh15khlLht8HLxdzYD0H4zHCI67
q44mLWUvfu8MGxqpDm8S+v2e3MMrhpojqVNmAcoNOToVyC//QVWlK+Xg4V/1p0mL
exdc7l6Ngi6n+XGhSxZImrfrdoRZ1PHT8mSyF33bi8ql3Y4m9sM9qZYI6GNPq7MR
C/7CD4GjizZhVEXp+L5Qe5W9yUoJkZMyADl/fIvsA+jWj0XHRfnG0Lhx9GNW2t2B
XQysJy36xjQ1eYS3sgE/F6hGHY2yA5wS+13vWiRJBYgMX1N2Jwp8YEa28vNYDrqE
B9Jk8hN9nxsvT5tLsamZDUXdyya8ut09A3adKfm+4q95BPotSgE791Ak7wipHp5M
hqW2Pb8fr5LDhOf0yVivtPI3gJb3PUOINX3krZTouSHrbr856kgNHcJW4JFvM0U/
Kudt1zPKGb4CvkT20sPYIWMIT+tGvtqNySM7SKAfy5kzMZYvo/KqCsXMzBcs8PFy
v81hBgjQxuYeO7jFLYiZalu+ht2zChr+vUi2VT/LaUe0Z2LbNMVbQTrKdYh0YmtK
GT/hEmNSIWZXZO8JmuAOI6lRGT85R/0moB57O5c+Ov+7DiRznVPTf90tvoddd3ac
TF5wCZlTm42fGPn+6YTWaLsBbSc+WoT6G8X5hqamy/f2+pZGq6uBWE6cKixqrezD
28+dN49NoNo1GegjV9l5zb6NKdFl00bI2vF205AudLu6LJdKCmSpytqw7j86H09W
EaL0NQOwnqyPaIoMVTFPWKTlR8YuTOtlPSW7N+XzO8/599KHSkh5hcqofICqIZZX
MANer5uMvnM6xV9Ln511xb0GG75M2Uawyf6IAw4DUocFaFSU+3XFlPxP/PBKxL4X
XR8bHTzSPptFToNSv5ldkylkvABMzilBY2WoUAur7CbimaOWXWvMZK5WFATJzBGL
j8YPGdZFLVZsakRjiAHW+59NufLXdvBnEmJ9jTbqoTP/W6Y1oDV5GxnDvhIZtuZw
c1CrxU6uWIRTNRA9b3qaSTXshb5eokx95M3VJgciBUx2pDtP6skLBoRDBoq4nS5N
z1HA3SvHQJM4NyaiVEGZUXjXJVZLPfNOpoWeFH6VNdYShZV++Pbuw1kPQzxLY5Vh
A+SBlXfFtTyubfqAwhF78Ym3G72bi0iWUXoZN8hp5Bj199biae0ryxPScwlgrime
g987z0cUg1lgJeAjrlS181hPcOaSOaeBJ5m5Cuv3QN1rkX3cH0O2VEWf5LGr8Ze1
5qj73WRcMgUbNgZoVv8dX+pxHxLVpXSU59FFQTkMnMpMlU/H6xLZmW44HYW7ilYm
vkeE+cIs6X9/+iJDQOxKJg621R0EdjXSEofk1HZnZ9S/qR+KkvAly0QC1cdSqEi3
6XN5Zc3i7xXZoGYAI0PE/XqlgyEdKlvyAQuKzxeQWXcXepGjryEn2Zl/tE91t49+
8VYCjsKPAikjHUxYTbUWzUAATWw87+Kj9aDcs2LAh1rW6p0q2zenBXtvRZ2sT/0l
84baP3To1gphoPabIsZCtRbqXdbn3WC5A99H9QEzbryVwf3uIkBSXaUhXpJxAvuT
Qn3abJ/3VxBI+sTjHANhw/HA+pTnWCMKYaqPSQwrKcitqeXz7zaNis8KSQZJ1UW+
1piIumaTAo4th3M1tU1/hPNMTvSR9LeDNk3C0RucxG7dAT4RFLTqB61TLkDy5S6P
c9CmvsxhWEAxMHdPg/o1H4El+kORx/w3QQHOugFkt4una5vsxce0Be+FHEAI43ka
ObJJJobFQBw0XVUs+We9Wh8HDNCkjwYt/aIM2dcnNf+40aRo82k6HqNf0Gp7qza3
44JPQ5ONn1SRdPHujlSRI6THxMN+s8fm73bbZ6slsMAKTKyC/xKNo39yb5tYFt1V
CtifFSoTna6bZZsvF3W/ki8MzNz3rAp6MsHu2vlh/0MHFbTVCnMp/hwfuE6x9Z5V
8L2jmgrDRTQ9mJ9Bep6oPPRRqFnLkvbixc9MBf/lrvCDMCDSSf+yHJcUbutBPFEh
naWSf0fBLB6dr2R85ygsnfNVHKIW/Gfu4LKp8d81ZjhO3KE0WWyoVZOH0BQx/mek
TrVoMAPLgz+swkbN6y7hHkIq4LaxkIzzUA0pYvMJw5NPnrhk8DizrrCXohn5mtFG
Gqb0F1G0TczZxVvY7la/0MuSbkv/KllOwNmOnenRC0QrZcA4lgdCSlmB4aISkZEU
w1WliL3ifdqKVCroqLSX+HGqWIcBlrq8FYnhM98pAZyBmhmqBhBmtImC/Vezz2+Y
JQrtXZSj/iwUZH+H0jXB0KCOJsqdDNYnwyvtOsm1vMggEj2YNu9YDmEYOBcyhcIi
duAi4AdWRuQpgUMvcTk+vKuK7aYTTuFprAm6se1bcy2y4aTsudzVuQfDUNsRvuYa
/G6kJYlDww5GW8uf96PHjbBCCWODseyZi4ZY69K0x7+YeOSpn7hUOhGKyWUMCx3x
2GnXHoVyMoyzTvd2itDUy2Eiexy3Kj76rBAQ86dkMR26zxBbw24NxvK8GunOBrQY
mJbm6YZXib7ovHH12k7dmeUGKtdQF0k054f1MmXwiU5xoB7kzuZnFjJQqiABDGKE
AGh4Gfs4juXQg2vllElEsn4XDN8rXU27A/CneMO9R38JkxU1COFLG7siBqjXdqcm
AmxhTH0NS7rPEbEDdR90otxX8ck2MvOH79/Qkeswby7291fWbaJjt0UuXspkWtTq
TaGatmOHZ7UbSJaFiuqW2MWltCt6I184Qt05+dK8noi8Zn3n8n5+l0ntapUD8HsM
HRe7mSni2yGDhnxBXH/BGYeiYoFl9+x+eG3VENdXSlHSeywZFp+jnJxx8uNQxxSR
zGfRScODP/3c7DXvZIAcGx4PcjMM4vI5B4xKQsy8lGyrtHK/GtmYdonvXehXXXhv
b/YSpvbpzxqe5vsfqq0FvZH5+UG11ilIF+JTPCzn24S4D7V1vAd4UfBjP3OZ9aLD
Fql3lStFxe23MOmjJT1TEab8qykQj/m3vLW0GbYhfqZJSVIJMdcUOm6ZRSXfrqox
ZR8IR4iX3ilCM/aQN9KgyDMfMdZop8HWK3Bdu3HqYhbvBZuTpvG1024K4MRoCw+k
Wbm7AMikWqqt43VPQeRzOON9vXOkMXoRdhbySHgipHY1krDMSF1dAFTX7VfmMYmt
yIjavFGKtPD/WgOyWU85dn+Y0prXqAGqU3PdgQC/MwoXhCPENh8aScmDltCixmTC
rhYOUqozeZfoOnAhFNxdCvC0BfL6sGirSwIR2m22gE6iw9S4fLjm9sm+ieMqT3hg
1gXOuwTu+LBvqniiuY/zHABe9KdFKtrPeYt06UEamLpOA9njwrtZ7FmE0A7DrLSw
64LAWKTNGonnW3VTQUdTRi2cWRRJj/eVSy7GSrXkz0o20x9nhZ1RBPhDMWxvw5zc
Jfc/RN0dCy3GXmfcLicLsdbA7d2Y6Ywhfql2n39FueX1jKZev7rGNWblJkTWH+u4
xFpXAnNfxD+YnVqRO9Q5zRGfPsS4/vOHlOZ2UTtJZMPI9yc00xgOIbmg0P+k8CQw
K2R69ipNqRTOc8b2rjfKQf+bI8owD6xusfy/YgGrMURfqsXTwSmvgsrpU1UpizWU
j5bhCaTLur7/OQ0b4kLZLLXip4HJQZ15PzOhuV6rEU2bUjGZcxPN3InhRilNaxqp
SuJ6uBVUhmSx5ss9s8anzFceGHc88W/5M2Bm1TxNK400+mwfqjXV4oIFEjuf9UJq
KXIQ0AIuhWRgaSFidK+DYYkzf7kmzZ1DzxG79edJ6m3x3gMBx8gc6es9DiVktfQd
ttPcq03VTyj9TvqD0952nKwol18vSnXLaKYJ43ibloU3i9XdTPDp27OqYA6UiJGY
Zw5tLB7u+D0Sm9skWz0EhqrCBaeA+bflaB86lq9NmT2y12fiSraDhrkSbvOTLzWE
x+WR6xoIDqI107gvt/ti++1eQbfdMX2/RDw4kRLz7kiWALtrfeV3eGtCIqFWqj30
0lRLyQKS3XyorDWHvWIFALAsA7XHpxBN4nbgaPWm+kuygudz0t5TnowLOw3Zrllp
FSPZh8BzCTuaq401WAD6sPwHFnadJWFJdsPq0lrB3nV20O/KcspFO6l36qjzdNPl
0fHvhnesI6bTH/lx1Ht8ohtCSdSoaVbnZZWuTwWW/+Zts3oYOZH2rqKlJbEviSZH
0HxRNSaLY/S7xakQZ3P0RjPEEg1n40xjGXieqFsv7yteY5tzK+JSYVlVn5z52pL0
rqCMsUeiOK3N+eZvp9myB0hpm9zzIN3QpTerK9vwq5bR+ShWuJPMc2vBpuH61TrR
Te7bT/UZA2kpMY4WyOZUDdZdUBSuF1+bFigE1QYjvAHaYj/aJtDqbGxmq7vfshO5
UUZ0yhca8DlSyoVuhIFyZn2NJbGP1haLaZM38AkRE4AsQMMcETkLjB1uZ5wzrBvW
+nwVmZa05/b9gtDoh9h+0wwo1dRy+Q0YM0yrjC+1vmONb5m9gOTErqhsxQnji1v0
GEV866b8dn17bUSfVi8m8Dd11giUxO/lNmFOz/zc/E9VYit1apoXyUZyEr25vlIM
iz9/WHFeY8PCXM4fOYuKNTKKrz5BVmqjOl49yE27sMS43wfw2Cgs6nDgJwjA1ykA
e5Z+B3RjpJdx1x5ZgWC81GzdG8J2dBxqSB25fqaAnaP08RUrA9mZjOcrXe8tlTzk
kc7H2iy/Dq8qEXO6sFUSWtC5QiK+WXCOsmL1mywSQt0wIT5x4dGKLcoyXmxPdwzi
sKikCD0rJQx1Qktlt3SzWyvzcnfMVqZ7nD7MOdsBc7/DzC9PX16ZDbKZKsSzolQ4
U2Q7w3Nz4QSpsJusg7PYgVkzJKR7guWX+/Xu1imp+/PYqQ5u+o0uFlnqZqKx6fcB
95la2GeQB8+NY3u0r8oSvJYtyBQg+zGvYzdISV8U1afsmugvy1Li5Kn1Zl/pz9aQ
Y8G9oIyHOXoNW3bua3urM1K2WWzxdY0Ag67PWoTTfMqxsDTWoYV6E5I/xQWmFTp6
6udjSeHwWFr411zymHRHL8MP7nqFIqsageRPxBvP6c/G1yEoNqhHTh4FuRmbKCTf
d9QQkiHivxOthpIBkqji+XNOvBCh0Il0E6uaRwfYid2iRrE450Q0pVds3a6f2WAG
eTsnY3c/55T/0YZ5uCuh6EQXfPrG4IvR7GYgSr7D1Xt3NE0TqlTrsEBnak2TAdKd
8bAnH5atwo8O/83IGeYuEMLN9wj0At1rsTbJG2rG3sKPbi9eLV2to6Fps6YmQtpl
kq2Qeu2XYB+ldZhm03Fsl7N63Pz8lqxJelwpUa3x1no4esicllm7sdTJ7XeChLo6
ZTD/7V0hiMDGMTchZ4r7o2De+LKKHskrZ7kCkZvFleEMbB2sXYDUDahgF/2tFQW+
L/oZgKrklSY4zdTjkGY5afiaWQBkium6q9KEvBQ8iT4nT8kpH3Yx1xXtlqGzDhkL
jRgPIeiUqhIeuCQTCvN0lVfauyYCdhIrcpTWmvcv9Mt5sptJe4IXLTywuZrcYy/9
0ZaqzTYA83NC3IE5ZFPQKLVipYygiYkyrUETmTkRsQk36VX/PJMq7hayGmyF9ZxB
M2Npy1H5HIml9pqOAdCQqCBOydVceNPCTwCWpFT2ykmfsJ3dW8NWHYy36yMnZzc5
J+55O9FY5oPbtGtGV9di8BnQqw64oofkHxqvR1n1JfTulZsVTKIXzxsPHBUjGXkI
5zT8mS2iQpWr+0F0pxhKFZZGegMHXB1KPvlyIOZDoK/+UDrzHIRFik4bZfMYdb4A
Q1uUI52sVCByuA3s2pTw7ziiALkhgC2NJnulBFxs71p0GiNISA5LN2ZgkYlU/sCu
03F4VMfO/GpCrjLLSBqYwOzeGuxXm8Pf3CzG4sEoUdDSwnvk0arNaYSZHszPzBsS
EH7uLM5FPgaTx8by9dFctcub2Vqfc/QqhH1ban+PFQWrRgJniHUN4M64mBo01N4D
fRjFR3EvsGEIw5JE3VBW/T239eO1K6IiM5DOY9bIgsNK7lAK0CDLW+fpFbTxzEZH
RM6o5CY3/gemMEfu7xp6lqkThfl2HPdtQy/MoeIS0NdGzOUS5LoWs5kU4Ec54iZ2
Y99AdZtTwELUdUAZV0Cyl2aB0CJMfRoeluNJuvu7EGtRBACTiKUE8BO33+y5ZVyg
LZ3I0zixzK/G0oL+E0+V7jhjS1+IYckDI3agWMVlUYkzsRWoRP20qcKWoZ8HjksB
uiuwc6SKDS/vJyiEyBQMZrGD5gBsvi8u9KDNl2hjysnOZuRXlHAYezfguSI52MVd
c0zCxRPo2WMHq9gJihNFy7GR8hokWmFWtTKLrU9Td8/HPn9UB5EQO45N0eIie+oy
uwtqbAqwvDGQuTzPo8C45EnnqK1t4JAN/3KbP4XoBnJARh9U3CDuth6NfRq2Zbz+
13lHzk4YGiRsBNfP/hojoka/hDDe9LUHeC9odvLo/5rUAryX685UwM01jmBwMwrA
FSJtDvfZoeekAAz2pcvZQLt9JkNVh2GhI8onrssDwutL0aXgQq8qM25LqC3VP6/6
mKIvOQPa5P65PLVyy5GiD1QIdxm0O+LC9VAdkUPlpF87QoZ4fYVNzXKIbsQMauuD
JysaCk6Qyx+iapG2XW0D4Fg3rbgTkJFctIRsAyPxFbWIwffKr1vchu/3Y9kxIjuy
UCMVL3mpsClUBUb1Xv7+ftHw+WBLSk8h/GZtHv+sXCEalq015ztQiNlcCCy+tjFe
SN2ysDd2FAeWsHtOavzrDkiUX473XfIpgc9+po+Uvr+aYUltcdc/HZPNmxhHIqUU
ZN0GtEFKJaFzQjyHjcJYagFaWKcPnkG+uJcHMCeFFuLh3Zk6AH6nxlTxi/Gyw85a
3Es4cNsXMQpTai8sVc4DfaltS/ZbYfTJdQkOSf1T81qA3WhLcn0MIVXjf3DYfJ/A
42tonUHqhSugrSQYIyDwFyGpVCEkC9HZ0BEgMwRwzBBsZiHmi74EoWvlMftFJ5Ao
EMLNkcFrXAhdHjHfI9C+5WBLSsnz+UfXldKkeJS/92FCoQQu+6Ymwb+F900eq2yT
PXvXZdKPviuyl76O/fMZUnQKFVF7RfiiJ39bTAelwlkxOKb/ffMjzzR4xCKTx4K9
mNq+syeBI+b5rdvYaoJa+lnpDiFO3cNWz54Uke4azQ2qQMHAHSnSLfUhqrg7ga3d
OsUK6rSNurriYSCuNgGF8GgDF/T4gmS44mZD7peu1UMSgrICv1Ubk0eCG91O2JPT
ZtAx8UXSDPehF9JhYa0FS7zZKlhJQw+1Ki6r2QDpl1TwfsG9DjnxYxPG6NLbZCMt
vmNnEBr1cP5DzqVbq1XGhwt/Lul0iWFOwCcm3dOkTNc68NMOg+ZAnXmE2o1irPce
G0/S7YkWCJlQ83NYwnUus4bRxCYsnf0nKOifsp/yzMRVyrm7fiXaKvB8uorZhcfW
InAlX2NLjShcNlKS0uwwSYtGaXIhxcBOA8AxCbCkJsSzjF6f+6xsPls1FNt2/gAG
vq4OptGdNeRQg06WUFgwobCCSmHTNmmyrb01LOu9xZF4koFSbvu0DUueDvUjyJwd
mHwLdTHtsKf9f4OXZaqs1w6hvq/dh2ESec6nTCj3caODI2oHh4QTtEcw7qyEr+F5
ytKgQw1jaotXTvSUYaZ/QNhyce1sIKsGjkbM7Cqss3Nia2v7yobWIjVGuEe0gy0Y
z1HhmjTpwDD1oirp49Orw7K5nvtYX+3TO7yWrYVEQx9JBDK/DlrOsNGdcs/qeY8R
jcicpgnfnk7Eafa/BV/0EnErvBbX7i5rpRkwO3ncH9AQpKYMJ+KsX5lIE9ge9HCZ
JdgafgB9ZZdEb4J/bQBnnuneZwfkU0kzMFw19Zp/91JQfkNal360saFjO9VpXiyv
2DIbg1bK99yr2E+BKEFPUrlg3u3DHNS/4GmbNUTFcw7CPbaz8Jt9IBHzdaJuAE//
4TK4lW99UrQoBwl3xkmWlRMvcTZp9GIcuOs1WIy2RZfiJxwK7I2Z7HxLAPacUQ7j
OhthCj2FjfPhPLNSTOfnOKCGULC4oiOQAHU+WDHmGD02rWU3pGU9H0FIyNSgGaL8
PpyVZ2bdSOUqKWERxivA++mx21iLOMsqzzINPY387A07yNUFEXOBmoKcd4YRkutL
As/u8iInSgEg22BHZ2QQu7JiatdfBXfqTIFr+XVJzEwcdbb4f77ZEJjUtu7enpyz
A1qFoWPSMh7wjG4YOr3fs825Ov4eA5meDByQD81DualJuYqgq2LS/uzP0uWlQgi4
huq3NsfJzOvWMEfdxDZQxjdwF8OBP6SITnmnPZx/LscUZ+mkWBQEzv7H9ZDb2Nuw
XBes8+3s8o+nV/0FbwarGc/gOOC2EC8WR1Ggkv0nCRP4I/SnyEgnLCLZnTQbXO0M
RdHpCHq7AOvg6gKPeVIP61K6gqvhK4KcqD8fpk/EyHYg2onSkduLSOK4uutIa3lQ
9zNymCJWZiurBNnODdVFSI/Fc1ZFMM527YZw5/KtArY7b2qKhf3jDoejSmmUFhVk
MRC2KxI90SYxNbn2FCj0skT5C3Dc9jq5c9NvrW01vHdAVq7n3kXcc+tdaLUjjnLb
frJaPK6UNYr9IgYNUxNzpPVgE+qHmvSwOQLm0zVrJsFslzIgC4Qy6DsFnc+JILyd
EYmmYm+Uk6klwSCAiUrkAXWjOroQfxokzqczXOB0GtkSzcXVIZn4nqumWPmZbJu2
lK6cVOzkAD7PV+Lz9vTkTmQ83cSaPSSe+A3y8E251HaHlUMmRQD9j+wEjMXMBAMj
7nt1xQ8kWiHd/poTbIzPYQnHaqMBNxyoO4fg+7Abx70rhu8/Xw/OGlKR4qqjrC4N
L1Wqtp6iKBRuRUK6JUbkJU/jtD4z4ntvql+HvOSNX15tLiMkBFIBLeocYdC6GGgY
K1pEbj17xB5On4nnm1Ixt3nsEsFZHvulpKAG4E3yRNTYwTaz3IsAep0YRA8IIRNh
wxrXmQoGv6Z5cFhT+vEnPP4WIyldSVM72iKJsy1tuuRfq4mz4Z1kEPmCTl1hIajp
5q7OtzNhuQolGF0kvkPpxldeYqTzSw+8ABTB15fdJWgKfiMTg9fmnR05vcqL/HIY
iSx9lSOeVLcvMHY/ur2UOA/Ho9sW7GHLr+8izN3Df1wmTwDRlJEU2bZVgysb0w2j
g2eYjyta205LskVZhT/2et49CPo4GOceI1xQVz/ZSn8TEEp+NFRN5IPQgwik8+75
oh0AeAg//mdjIoM9ThXKACrQ4BsxkSKnq3byMSjR2ssWESz+rELm32jJdpk6Pwn2
S1qWmmbyzYVy9kb3w/gp678NrtvnO5B58VlYsRO/oJdOuSmYkBJmqOX0sv8RGOgQ
Lu5CKnImebAKtOjC6Y7unkhb0J1ckNLCx4wc1mC4WK7kSjQ4dCRvvdabNwX63ixI
qIv2gBbkDymPQS42JwSkZoPbfCe7TQjR1a21zM5aG4H7Q91PfFkPz2Sig8/OOo/w
X5GlwWXDryt11OzlL90BhIf28yrXUfex3KPBkmtz3WBHKk3nvNTqiYTv6PxkUCuP
dy0iQXKp4A0SFdRTANoHZvgSoiEU0kfSS/QPLt6PHnWPDLWiCZQSXsH/zXUzLaN9
cJCAKSkHRyu4xvwoEGcwKhU6DxS6uYPaDpOK64VggVt0oGZDURJWnZj+3hAxOa/u
hoTzDNZL+p9mRqqQNH7sFjCT10sjANPX51APzCL+0xFunr3A7bhKJSDKMAeVJcFR
StDfeTOu/Ivmb+oKx6WhnOEf7R5AD08rS+vpgucvWR2snLQfL/iKR6JnDUPriKWJ
0Qct7UTv/FBk7dyVOrlE8NEJfV77n/vw3FUq6MhdtkxVTGH26gONg1J5jW3iaOF9
Jne6xafe7AhU20jRK61dQINF3IobECL6clFbEP8+bV2oTgC0bIR9FoDqkEXedeZI
maisfnVsBv01Qoiu+BF3hN1xNypN3qNmoDxd09ctpOAapbrj18UisyMxaK3pt6Xc
u32ixdjoOU266pk2rQ6LUcQAAR8N+lGbRtooT+DrCvXY24dn0cydDOjFWJZOPQsS
Txfqwl195to0XGQSmn0MkQwm03FEFnI822S3iAXs19+ELImoZyO664YNsWCjnEck
y/AAN8h9HEHztAO0gRECJQrEJoPso57/ZojBcMvLIMMw10OstlolMo/rYGzHy+V+
9QF9pEKJe0tK1uA1YKKFUKwrawqpgt+JrPVpB7/BPt/XSEvlj/nVKcvOqRfUfd+d
D+DCG3cURepRn8ascgUUTxndlG35znHL+b0dPKnvuRLFwalQci6Kzmj5xvDkGFX3
IyUTgxz6H0m7c3opib4DhCZQo2hKHWqe3h5kreEqKOSZZZ08OZOBLi3Mwybbgs/q
gx9iI9bAuXVt3+Hi8cwKMZNQy+wVL3x8oyiwJBaxZ6C8Ab2H/p+I8Vhnnb7dZKy3
6WskjYlqHFM4URclcEwcoCFiP4lOQCA06t72CYKIpiKajGdxlsIOEcJLM+gi3w5S
z6z0VAzSolcS2W2CSNQFJLZtBaO6mxOLXyyQzSBOwyN/GxTWMKu2eyIc9vNHQdSO
AimdFTq5d1c+6d/v2HTUgJCb0DDfMXVtfsXhcfp1B8q5UWQqWgiqAfWQPwLuIgg4
qM5d3QhyFll0lERGfMuQNZF/FTMa0IONCXswz9eKAvED/J4Qyswvq6Q/vtHFefgJ
HOLw2WijVgwqJa6U95v7p1lFzEJGMBbRgO56+2K/QpDp1CX07+6gw2tr/FSjj/sK
vyT/jsxCQCwE2ze8Ysi5sG37s7tuXC2r1QBMjl5MJwvUSWQhoipY6kHBV/RXsQUV
goPDvY7qcyyMP1l11aqW2mkCe9J8mXveOUxVmlG7nYlitP9E77lSZZSvvsoC5sub
BbfpKG9xsQivARV8KOkHokffMYv2Xa9b+VqdpWLpo9433mLI4N+1Pl7l/2HaueHC
Ar0Axe9uPS3TYPGdGqI4niAKVjeRV/ivV03AJmxvDo+/T1/nYhbIqSfJ8J1nUcb0
EVDiYSVKv9zw870/8HvAhEvN0qlWMPr0y+y2nfXWSUUuYnxD4zR+K6n+WtWTtdG9
L6IjzxtbLVkdXX9kDC0sug1CkyAbHW5tHuLYMBCNQqeUd6vUBWN5szwpoklcjN9Y
sHvvzmUZQQjE4lfdHagSLsqYhtesf6mDRqmzdIkoLdqp3A22eaS2YPAw1th7RTyP
X+fALsBusD4uNmpzqmmO7n+PoD3HKd+V3sBArrL+hMICYfH9CuAVOYtX6fIJf1sm
9I/C8zg46NrsPZRE3i2/dOQMkKtxMzM3OUcPNYoIBgAU7hmfPMng+FEN3DRvvK9X
J0frVOAGd5OakrIWFZp03N4CdTZWHuG8BQFx60MEeT5OutcUrw9uX6Cs/Y7QZahJ
P+ye2yTYl4brAn2W6VxfjIm3iNxWlUhk24ovyNq5rODVHj/XZftjZNXzPP2fWiC/
kpani5bDecixX1ura2c2QDC8Bfg13pu+1xeVxIIxkeokfRRC597Yd0pgOEvcrBKm
g8cVHVhHiNbn0iDS1lPzUV+BPCwSJNEXf19NW7sQrgMI4PKjQl/RTk7PkqFO36S7
S6n62RXqxUdmO2jmovb60yk0ww6SJ4Om2YVLdKgK35AtXhZpvE7W1fQjgi5i3Ag5
YQKPpZDWI8v1Nei6AHuZuSkhaVqsP22LWGJmhAnPH3sCJXo9K9zJDuqfbSQcMJZc
i3sfnWgYzJbWXaY6fBmfeYrdw5AG3B4T3oudDpcn71DlNFDAQqe15ecEee0jbdLL
+onLOOxSB0ioEcB8MyTK+bP+Qq9I135wGZXuATtfx/JaO7kRqwcA+cyo1QgHWbek
QDxQLIKzHj4QwsnMqOy869ezdQ+a/TQtTrjS7MFEr+40pAwXkhljbYdc+N3nEF5X
opkUNBrRTAbXEWEB0wyWtXQ1p7GfhhZLDguUma12vbwT0xuCSqhTIsycCVcPoxml
paT3LaZOqAqWmMunkoxMuvuSlt89Uad1Qt0uQ8Qbw6tRQq+DWV+38771Px6PAnP4
JY8u/qQJUd8sax0QKs7lp1nAAA1SQZ/PiWjyfR1fslUDoE5KHZNCwUuU2v0ZGleX
hOpNn+GjYJodPunxKSgQ1GAJ/ANPpCkgfLPAusU7Lytzj9z9pia53BNaQAirz2JQ
ShSt1K3NPluYjWD12A47f3K8FxRt37cH0gWh5xXimlkfsMptaXimOGP9H5AIxiBL
afG96n0yuMGCek2nM1rhS2A6q2Zopnli/iAt6VsCUQ17mjClswQ4CWmzHttH9d30
2CCwqLqqJAgak7/zJegNI+rR3DDHywNK04M8BJM8l2C7VdCUEpActgnhzo4zLcSL
xvzAP0UA0lMFUJOu/I9J4YNLYvYfsJ0bAWM4bjhS7m30qE91kZd6pzA+fHHmgA5d
BHEpcEHV39J6XIAZIxn0/nZelayg/MLyI0qxDKCzzsO67j0xTted84Tn3/zqeVE+
r0/AE0MH8fcV0ChjwIh26YaSoexAorMnMnqPqMme50NmJWmFaT2JaQ0wqEaUEHyg
EC2p1WEZUfIkM76cNFKdCfJ7WjQfVnZv2xydvpYBUpmWOn1uFLMOEh1umqBWHbuN
alIswMmZRIn4U37DPAYAPjz7N+KivGn49Uj6yfNrmwXyF7ykvc77yIA15EaRbrU/
BpZn7Il2QEn5tRsQPe5gPv5XLuGaJrFKsfIn2l52wtVRRh9OmXH8H0okNshtRsK8
QPEJgteZ/sB+ZurQ4mMFx4GccGlXHCw9UUo29UQC8VLdkC7Bk2qtcvrHFHp6t/LV
VQncTnNwSge8FOB3h4fyoFhuGbMbDSFCrmyI1N4m+usdbkVcKe8hrA3jXGXWAY8l
IHcfoi+o0eq1JfalLntrUr2aLhnUOJAtvKQwNym1T1Ao3/HT8tMSq5JR2pYQuHw5
LX4uMUGsiVIHzLwAfRfBDw7MROi7O6NqyTuD2rg8i8ERximRpNV0w3nhft96NaCg
lzu8gGIYIo+hpWgLx3zb/mnuXzwGyAx7md9j5eM7zwyuRkAvAXYlbmslNv+OAbVJ
D+eqCM6Ik7pA3wwwkUaur3zItCab/Es7xlKSuLH6KacIPIIieZlvuLewtdYuMZFl
PBQIS1cO+MpLxK7cMDXo/oTFiXCCboYWiz8xkRHT3FsL2sgJ7HQzukHBWhI52ENb
iKy0qgwH89Itq2YXH+SL2U4c6ABGhuAaTdARmkFfbN0C1S1ayA5NLUNlOUNIUQHu
yRqKvcgLUnHLp7tvo9z+OIE4FZLfMOx77Oqntab+3kca8oorb1phbSHx4PKSD1Rh
+28uNGXGl5eoRn0hdcz+6zzOZ/p8cainOmbN1/ScIS568uWHElgc1P879g/m/onM
jFeJCW9dz5bEnDCD5y4Q5ai/KHVUB+r3jSRjhX27djfLI8Rw8W/5IoXMfFWuOawR
QmkjReB3QYD5CMGawh06LBuOrLs5WrK8FgeYnX0hJyhDXysyanO0mgutT2ixkqLE
BmjbHYyU3L/sHn94s7iCtHH4aqU1Az4bzsVc5ZnsCt3xdnJ4bcMRiTHkHjXnW5Q1
mw67qrKlvPjPnbXFB6rL3n1uOsS0dJFC5+f3H67s1tI9FLpJ7UIZmpaN52HWXozw
yeqxN6wAAwJXWbrr81HTT4rm6X3DX61pb6KP+/mCByzvAzsSuP3tahGiox8z0gYb
9TcAhpN+QEKGWfU3KY7xV8OvyfbSMAmJ26ZjrsFDJOd8F37Y/j+t7Kku1zc6fDBX
08LvVkj6ufqOO44VxKJ5yh71MFsztVopJ+EhaFyBeMuGzPgG7P25I3am7qwkDAZ5
ZKM0wZ26HmwhnP1DeZ6n9iE+RmkJDuWwdyiTZ9xlaCdCnLBQT+25OHOnmL3x03iU
NGSSTug9/1ls/sg4SpM56gjTHs6Z54eZjbPl27v2+61WlBJYT0giuTnLnhSQO2jT
NqChEUyDXvtXzp6gM7vJsRqpWBPDo6nKAprmotV68JX2JBdp6fC1ajSyM6jDFera
o9R8TdET8+EQgoBp3aqUuFVmkS4JKBOsoaeU8hNLo0WLR64stcUpijp91yk9mQZT
EBeiEKVHbFdwR6ebejg0IbPT1+IeWy8k/qXsI5nj/n3RGIuXrzutsm3GFLf2gdpe
7Ta3/lcX/z7e3qNF8ZfgbkPDmdTVWqq7W7ElaYFJbW8vYcSnFPGT553S2zN79Niy
sKNjxBb4OqD9YMIMTkwaaVYDqDYHmoe4UkGcGeqTA23E01xyL5BJ1/IGrMsNK5St
MhRInAr6Qwb+YsWv+2LngYLndOX7zBPkFtlAXml0pbAUi0Q7CLG3ovj+Hr7Fwxvn
Fw8S63HucPrJo0p6JulzvlarhZoXSZ3mTdCeOQlUbecjMBH+x/aWwQFES4l+QiRF
hfvzQgy8kv6JYOW8KP6jpRgd8qnQZA7ZVsM2CMsh8SFZvCS9OHYrqVLF5dfdgmmu
cxveKZfZLMo+O3rEjiIrlmvQ2hZk1R20yjW0gSoNyI8UUC8elJwkPBTasFNoe6NI
1LXk36axQBTXik8ldQ0gxxRkZaFsDzVSgJjbhL+4P7V6iUusgJ3MABdar7/tZcxf
HiQdmSUw7ff7tilH2klXPYuE/v1KmciEU2Bo2goJlJyTER8OZEnC8i4+fms+D1u8
DKN4goRvdx3GjDY/iwLObPauBoG9aw+a1VRoAfjzjShkp5r4z3dx9IypuQofdB7t
zU2hidwb7zs0BtrWiFsIhRDiW0A4sdVk7S9w+miVyWLT6cUuEOePQV00wrCuDNEg
J5Rg84EOA8ZVJ0WijvxOOxcSu415HtQaXSKaFkbZqr7atC9hegW5MaF5qW3v/T51
t+2RVI1Ya3b4NaRQWrEkssXjimQQPqc+GVEKhzGiHapzy2350vKGKQiG2ylGaOcj
M8t/dh33kw2F/YJ2FGC+wxrAhDr69NCVVF2kUX5bQi9P2ii/AdGpJ9XRyuaT+jyG
SPR4JFg0vvQOh6VZfVCIzGGSu+Vpifd3mwW014a6BGxmpdB6vkjGWaYmKtxsrAhE
kpmLjAGZwMDF9SVrDg357WsekQtTdNVSs1Y4fwGo8fufkP1d+ndfk/HmjxWqNEvM
1rw9njv3XyDvPdZRu7bEvzflXyxeh9xqUo+7hzGKzc4NXCHWDCQc78MggCpN2ucl
5bisRTX/f/orhRAdgIkoPsRHj89CKcFXQGZN93M8H90n51uvO/7wMW/BE4gdkuxf
0/AcvH8uspReBnmtrPWZUAsRLZlWI90u6q73pA8SNiJGIXaC1+wTR2gFzKiSCYeQ
X3S9dhUqdoihuakFYZ6NcjTkW7KC/UHPiOnV4tcf1+htkZmtglV8WBYCRaILorYz
OmJTUiY6Z+ZTucdu0wkfeHMq52a1P8Ie+NLPVxSboE8li4XYDk7Qg/U6dTX90N0i
uDpsU+cWWPLJx+Y+qHbQ6rCfKXtTvdeC+jPlciq6V2chflvAkDuuaeoNX+iKLvAC
gTC6g+/OmKQ8tUSKCXKdkZ6GY/8OMzZYX0IRrX1Jl69kYoLQR09jW+TmkFjb9fnR
DmpDSV21jFpzgnZIYKn1racXTa8ybv1fKOB2E1EA2Ot4uXcggUaxowvAStBwikOx
uv7Q7M65n7JZ79cSroGRtd3lyUb+cHkmWe7eAtCaLDJR5o3ylqTdBhTLNbI1BESZ
26wSYyPW/HLvn4eVHi62cVx0CuH8zfWAstkv+ZZ7dkfD7np8y5VqRyLizRtlbwgO
Bqk3e40RCZ8J0pKtah5/wqrEGpreUwvUlhOieGJw0a4FGuSh0t4yqbQkMsBp8NP2
Nv90/fQgf1fULlmrFUMMuttQ0ADCr5A0PucokzA29lsgZlTz1JY1uxcxKcNcpVJC
x0PRcUKgBOjbjFT5dFs+qYCZWclZBYvWas6F17kUugTj4qyKklB9zGzQDSOXN1Bl
EmhR3TUIDg4tVDElPbADpnopUHAplMBwfiKL5shHSooaaqR1Q7m6fGyn6OQBlcSA
psGVW5KO2A+P1XcpIPZDuFBmj1Ut9kScCjprjgV9kanonjYa44qn4jvTNg2bO3Tm
DrKx4ju122tEYlS7sEXqiUG/ZLeHSNwqC/+31C9nkuO8+Ac3Ab/4FuGxlOJkwtcz
+psuMYLiBj74mN/RNa+MPG//nNnJ/2p5watSF+Mn5jeKHviYLdF7ONFiFsqJWalm
DnZRmENrNLQ9QTW3BjYu9FhlkV10nPlBUWyQh6JV363L/NNhxm0UzBqeEff91OmI
r1FTuN+dDGvV9+eED0uTgDvsp9QWNs7tLPjILlaTM33LZlwQMUMKHEoZEeAFSXHg
EWCjECR2wELCphitGuRrigAmoWFIp0LLAdEMyC+t69TlEqnMZpjHLaXGAgyGG96V
vmzR6EpZ4Wt9BWZeLIOCwCCF9qOW3PyoneLw8DIdFE17arOTLw3VR7eAushDpul2
KaJXh/2OHXtzXlJ4iL+yPJS276chDyIBjqFBp1vLN2G1ii5Nrmr9b/iElEbZUzkY
9k/2dVbOJelGkmjCJdOAU7d3f6XQF4a927tGnf19907d8zt9L75OHZEWC9Ptsyqg
kQ7pWUVzOvi7r+PLc7fzqwmowSDbR3ePfqTBNOYiV7mqRSBClnr/WhuvZVT7VTtP
LyKS0RWr3OoNL0xGDOhn1xiyebTZAC2CmV+ShV7UWamIAekwmY34cVJjZkBks4Ov
Kl9CxZ33ITqDLQDoNthIf2ROkM8RQLhiyqoE4a+flGR8dawVnK1gjGH5g1QgJpFa
D3OC890W4gcL/gBxFEdG6XCHZwB59IekmbAw7gSm0fPZsAyayE0cIzyJdC3njbnF
/j99bpLxzXzS/oAGft76p0u4cJWqPR8BYkSX5zaARXpjmzGYb/ovO7PgX2ULl99g
kmQ96vUjB+gfivzPg4hM+IB7zDlFqJ2/snUy69Gw6IOvVYvF6qpYYh+ddW5b9cfI
wjbiEs3hJ6tG5XNzEvuPqnHn8UM1B6sG8dHPIw0uyZuyIDudkpLSaJC1o5HrPwu7
nU43ayF5now9r4DcrtWutdhbh7u6VDN0TOVT2FGjuPHqb6BBc813uGXXuYzhvOXN
qmPkSGvS8TqXO7UJcW3vl3rpY6YBexJ74NOJ9dp8Y04gkmUiyi4jYoyAULYsTRq6
FH236xKJJNxoGKiQOuV6rzyJ8aR1+hDdUD3xcMQKGZN0NtScbK+LJhQr2rH5nxvz
cidXyHbiKTYTb+Pujc10UAr6p+dYBsB4R6PpQ3OOBau/Jy+zPmgfaq097y2fnnsQ
fHUPmtlD3lwsr6069zuMlPPTZOTtSzurTzMz0xFVJ3nwgZygDIvAV8jNw8t4lKdI
Oim6kAJps789Luhh59rDrE8SnjhO06RwifNLg0U5WWZ8tFPFq70M3URJaXj3M30R
qbwL+bnor1jVRmEQMQQikG8kcSPa+aHKXtMfDbYThmvYWcMruBfzB0CFGoqII+QM
HLqIqAnQineNmigAHQ5ViYip1GCqRaTWQDEPDquQCH1TsNNXBodcijTOSCUx8P3N
fHLsNfRaVOdC3j20En66WUyBhd8GBMD8kyVCfKocYXLuvPICeMCdgfAeUY3aaOD2
Ei4hVnFx5vYETAK9/FZcTqOhD3btyjdTHbbbbOptooun2lYehXKqqWGgUQnggjVi
wBDHbCaW9l8cos2baNltTlr24N4c2fRbU+vFBTpfcag7yHE+gnObfe5DcU5Ur2Vz
Id0VMDeAh++dOFl1DA+TPIY26Ty3jado/lVYfdcYJVRkF2foShtkpOT/8OXkhzA3
9jjxMUfwHSIaOuh07GcESg1sf7boVyTJ7uS4tGobAK2bs6mHpS5vXx9YjWJWPhss
6NfpUkppYbOS55+ksSEgytGtUwGM6BIz4NV/xR2WF6wDEDHpBW/tbt+sTyz6VIPv
mOysixYSHYuvuMBatNWmrmmMwYsp1rGTFOcDFVKWqlRZ99XBIQS/2tq+NWhv9Mrg
pdDLBaRs5erJu2YOjweQ36DleI8LCwT6IjX5rOrHObTdLqcGt5Lk1x9bRroQ+r6l
UqR2FpeaudMafvL5DNy6IST+hJxPZTq9VxUSyjr2cPWmr1w7ObKZGJswfYdTZ44C
tcW7cOow0QifEZxKxojg+7B8SsgxnowvS14emwjsSUE6uokDtuutjAMDqICAJq5t
f+jbDDSl/qPXOjiAt5L9L6vTA4VNXyjYgcfDeVGoCh8QpoNLRJ4hCqhxRR2ZrqjA
ZGwr2vMT0Vt78t/dFgOoPD+cSTM4GXsUH5gcYhGi5aD8YU6TtLhkHx7VNsAZyHYT
q+5MweiJhz7o2sG15JiRZKpscY3ULkLw6I0/TTAKB1luoQDndB6GO+Th5lOszuWh
UF1wEkF8lJeSmlclYqdM2eMXPOFw5JZO8PLGDP30fadjlKpTYSm51tBn8gi2n08P
Q193aCdUXT2MmL6K+a0OBuIYBtTWTjv5JX+pt5eEqt05cuSRFOx+2vTjwo448wwA
y6ODzklsgkR0/wZoJBay8y43Ah7sZcfYwc3aHuboQ9jD4AYo/SvkbVAucSSV3WzV
z4O0VRcY1A+BMJPViFRIfXvlS37j/W61kw7hpbm7DOCspZJWBPEMX9574pMhwejE
ytT7sfzqdF2dDRvRKHt07dssC3vy6fA2UBpyK2uks0YNBhKBK1FhPeqU4GLwTyoI
dSEJ1Ymp/AYUvumP+U37qhIHJUgGMzwduhm6ECh1QursXTLrbtqx46mVbSZoJ7d5
+MfBVWTu2KMbN0Ow9QAT7hrkVO1m+EGsyLhwdmF2RLCdQQbPEkB35RL10p/zEtrL
AMIp5QoA49RTuSpnD8aUxrHDgiP2q+0cx7YKxtP04fZ8ZvYIuIMimZ1M4EIv+Rvj
lO1rnhLPjF8m4GiRi8BFYDEwPFRqsn7qrxcZIhJW4vJGfwYs0WRuxKAucAywPCWd
yFOM5yju16Lu8XjOvHV12WcMnEmVgQz7y+ij/7oJk9arsOx+tRuR+q8jppvXs25+
AXMLHjLpPhu6Jc9hKys0sNw4ny2vzrZEc/GehBScXzaSl2TjntmKOebqcG4D8ct4
ckwJGPNqeK+3b+NM1AZwuWsypdqy5xE/RCLA16Lt7is3duNXuuUK+SdTbeQ4BspX
k0VqHfyGKAdz+d/6SpQ82QNOk6Dfc+TXXDBd15CRtGWxa6/CmbpLH+OiC+t+e/pS
qN6/c5u7d3qLh3DECq36ywaPIiVXnc5a/zlbFNxWnHWOMiJfH0LjJJJqE58SeSk4
30WAmqN1htuQ5+q4X8Ydnn9KyqoexLXEZ35V1LFAbpxaeDevBk2/iuBUyc2ofbKn
bFfcIXbo+Ocs3Of7kHhNSKBfEJQMXJM3J951hgxEfJpHZmkE3EOaVLRA6H2pCwA5
4RUfjBNsGZSNfZgwH673YK+HXlGtdIlS/M9Gzi5FW+I0qtcNSCm4a3RNKEuWmJaA
EOcOeA1x8MEnj1qR9rXgqdfPhAL7Te16d3+xnT1ujImi5yvQ2X2jb9xZ+WgwS/Yd
lDfoULIJnTgcOA+/IRMOk7CDbjLP+7GryuoUjuNRR+BezC9nGDRPVqQUZh3nT72S
fBIX9V37J4+7jI623A6ScjesFRsNgskhllh2/l7EfaUo+BsJ3Q02l4mZdfaBG8Pc
IcPOrgwr9pggqDQz/F4dGgyp0DvnooQgFNv4ibcN17WCCWvqAPjGGwocdmIIGi/c
zIwc2hi71YnKhF19UdblkHGW3hqsqQlvaExQ8ZO8UNAc+Klicb7hEJBBJFST8fAY
qdt+ZLd3INq2d7Z4OdRa8p3u1OxIALfbV4SZhOxmtPjW9ecbDwFEdZ6aJYtBrbLV
+M6b3eGus62uRxVvSWMezpp0nlh5N4B8vmcfaM8rcbyztXNysgg8Sd7dB1t5tbbY
TrjPQjZetJcL9sz/mzb6KvijJhACdva412RNg7h8RF31rRBIQtIObMkZxQzYSyz9
mOIz+aVQo7QO1rPgS6VXHkxV88Y6F1wxn2VbLhtKFJ2TbUdhmPe0ZNLWPU9VzUpm
0lNoDC6GB3e28xebtQkAWfPY/cVOOLYTIqZVZgmQPd8oxztQ7rouXMqm4eWGwdh5
pIKAcrNKHQE8gmKG5Y3xcG5izLM3fi2BscbPHuazFxCslLzo1mo273EzUtUNwKY/
+92J0uEFy6UfCUs1yTVCXfwTIt4uEgQUjIoiik8EkZv6nBJZDr1NDTRxATNeYH7q
DIWjIaaSG0FnpcXynj8DuX6RFIpyAiEkGlraRcwy4wUnBq3tJjtX4rJXV674uAo6
BplErzYavgsOh+bhz2SWXcVdeN+/dItkAFoFerrNi0lTI/4V9UyVYM9dhWbqvjwv
ygQTWt8FJ34kmrp4iLQP59ssDAY/WfrG8Pe3Rtwh+zsSXJZZmNto9KVjhCZLLBXF
qLB1M8e6InPuyC47Dbb+LFHCRobAmNF4oYtDNrwA+Bbzzt6cfqr11yhmjFPSuP5r
f9mEX6gBQl3ZtR+zYSOvBvf0wVd+azQLVj/QBfxd9HpuM823rUJgAYubhE+PX9Nf
P7B9YloqbBygRcQ4udrmPizoBFGF3zypJMvksJUZmF7F4FjEaIRa3N5iPeuONXYk
wDhMpKZ6oi0wERB0uLDIM0L292j9FS5Nnog4pPljJtHGo+fdKSTZSDKuDyrTawrK
824FREwYCEL+358OSEYTkbPzpqNmBiKc9c6a9/hXpO/23UaC6ZZtMlHB/es2J2A7
Jaev6u/KZpw5Yjg5at6ePSTHpvmiiw4pg/3F9biwhgRAtdwWWvh72Ty+iZdzVOup
UfwkmxlK145WilpeJNoCZ9GsjQ4mMSozVH1+Ueksi/8hnu4ZaKUgFCnIdyKpRBVv
uJH49Ko4MdPbRylJH+naHe5HLkVLbo9WeecpFhOzlcZID0OfCDWIVRp/M5kVVPHB
IYudmmJJ/r1rnaL7HPEiby3Ggul2USy1ZYoA3kaBtmxzKTXnL3py7FL9ujdGKbOx
Ub2xdmcfyqbMiTPlbDOuhXHspF8NMyY8skJaw+PBqLN4m6drcAgHUMEvmqJIsqvn
1iZGdGsroh4j9dyn5zZsJmVadhh8wivsCC9eUkQJcLIkIyKHaXj/0gAxD773S74B
1gGm49fRufz1nIW3D5IGFmwyQ+vdFS0IaLEjm3GUDgUdW+aCAoduGySEPegn0dMF
DRxcSVR72HUpspLHPwNGXur/MWkfj0jAZAmIwbMdhwbe6b/kyBYIIxQDuQ0oaJog
lD2eg9PoEuwsFunieCdj9AsfhVDxFgqGGoOzsTlmjDUBROzpwtoOaAO8xt6nv4FK
6BGZWqlBUROuTlMobxdfI1c3EwlUU5S/qUkFQWKIQVLM4Eh3SbVmohxuyr8+byky
6N9x/6fpmg3JIGuyuQaIuYOV53+s26CauOvTIA60Glafylq0ADWKmU1j/WAf4EXS
Ncy0nVYwuC5eo9LSQMGAJs5nAPh/DJtz20gB+BXc5mtFgYa+w54oBhcHxSOJ5XYs
aj0lCHeTXDPtzEWSWu5Wl7motZM4nnLp4m60rGqN9Kk6CaGcPO+YtAEVJKT/EyN+
ZcO6SukVDxicSgNv7EURZ5/xaAXM6W8wTS6zBvboAN73yZ+wljexhPrC0V1QqBaC
d413EOi01OfVdEhti548QLHvVdTtK2JA1/UKWZvecnDu7y+0/hPyO0suDkG7jVN5
chIUggC6tcn7mUxT8kx4fXrbum3cUcNYmakQ4NWog9ylh+Qm9y3biGTj/ECLJPpf
+BwE3mz03AlGmnQN1xezcFcRkfSfKw2wQdciO1BAWFD69KsgZX+r9LZS8jVQBgYU
fAmsB+y/vzn/ueTt6rI2uC3OwfxviTnIBw+hEo3XsByG/BrFRIY8PVmRVF8+Ee3m
gvOcp67KLuK6F0z5Ds+5wtxN30l6Uetek/hG6xopmTmZVAXLSoFEmLQC6hAxZov6
14IqLabNI+aN94/F669pyqceX/C3vbs2BN5mohkubZ6VtLmSFZ4pbrm5pcii9cep
h9oWmZOwnPIKhZy3vrINKfX3MA+Ok5NHuNGoefJEe39v2M6udO4HphUcSCuAM5Tp
FZVpJAII1EMo/hlpyJorSh/zvWudeMrTt0WT/lDKhauy8TuuHBM5O9DzOxFm5TMd
b871Sjo23YYxgo2tggOmNQ==
`protect END_PROTECTED
