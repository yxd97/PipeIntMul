`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mjaEVe2hxDZHTYqXVt4vhT9Otu9Jidum0Mad6uex7P66evdnFcgz7q5ekFtCnX88
Fzl/LwssIatzy5o8k2pewbt+ge8rgrw7c/uE7Z6hT2tichrhGgrQuYOnRY6g+fzA
8p3LLDiprEmLJjdWaoaX6EjG9SvIMJvLsatf5Fuwf0M6ip5mck3djAG7+QYDPq6g
iIqGZuaHhKe/JvZ5UOlNWmGnmQ5adGu0KpOUCoYRWbbpFTM2Dw70P04MM2TDqxoN
/fQgApUdvoHtsInG2v8Ra0A/mzJuDs1C9ef+nDJ6BmwOs2nFt1TKBMicXPBp0AaQ
TgGQk1cWCvOKKUbxWrsrVBclCGRi1RhjYsSapdHW8RDcd75ILQosWzyDB/9GhuxW
jqljJpAdzPvcyaoWVMRvWZTbGY2hiyjPwzrp3QsgFrBuZuUlkegG0E76zzVsvkL5
GDiQ18T584zQvtKTZ8zloFBRRfOHven57H9ht75tcbyM9k93GoAiMQBKv17mkVsi
RRGznOnkD1Or4WYCZSay+AAbsgMMLbcCB3VnLlu17CgMPyNurSkXFia7TDRe0W1S
ciwtK1OTHV7gDLMC8J2J29ZmBT6idohPzotGyAROgBAbWrVmp3uz2pBZDpoWtjup
0O0dUALE8IhpNEPzDu6xJp7ww9fJJm+y6RqfUQcLJPxGi4LnDA3lL78ZyzlLZTde
a1ReRQXr3RRFfeE9Ijh4E6Yo4MXNsxbLCdNZ9UKakpcGrb1P3WI4IcaJ7x0M3JvO
0dXxxs5Xv/HecLo/unYGA5vcKNlLVq+cjYUWhxJ6PD0qMj8FahjLefx1WKzMRfrn
5QNEt3aLcVMTjWdAfci8IAiKVLQv5J9mKe5yDWT5cB/1gRI4DG8f0KsnJbCWVzbz
bvz5odHHJ+VBlKI5BoqDvJbbcAPQdlbfhOkVRfHkgx+BEBrbxFeRoFu971hUolsP
NK1C/mzTJhDtUTTSjwJO9g7CVEsV6ki3Pg8rLG+8ME9f6tCx5fVE8I7muOR1MC0k
iph1UowbOzNb6H5Ir4WrogGSUmIpPpOgjXRGWceORh3D7b7TyWxa4AAlWu6E7AYr
m75n/jIBBaklKVSPImnTszAvvyRcql3L9CrbbnFVTl14ZIutTSJHypacFhY64VFc
z4/m/zHoR8ZnqYmmwjZBDA9mFOC8SXoiz1QhVLsTEEJfNTfg4ejnaDI56b/HLt9H
yNpndNa8u54RAm9i8yO41O7b3SivzQE0Xw4O43twoElOhWQHEUAIA2ljwkp/9M47
Z85GGz5RSQrx2XQgtQiP+0V2q1aSa6871FLFtjfFSSv3unq1+siyl3QFiWQzIZkz
0ocBslXO0EYt7i1qPqWJWkMrqf/phXjUGLnAmwE8rbJUenJmZmIYJvNJjNNIrA09
tZ8C11W+3rob+skw/a2WDrJYLua/dVTEA/ncygf7ubkkD5gxAEH1umgzjYMMpYR/
2/t/sCBUEirZUAUrs6sSvjKj94rMdlvBUoznF9aVcbjzP421k5khR9bRH9pgCrP5
APtbd3kVACK+kjoDO/LlsI6g1ERd5bkQq/xYjJ4rlI3XbR8eBwZlGWJ/MIEcY3Vl
bpAWqQLCd42DXeOqA5kxu+9vbMCbAZBTKryteLstMi10q4ejipaLnDm3hVwAEX5d
dbWC6Kr1x3lNVLM6lnCltgvkeLCYFErWCDNVZK5H8qUYAZaDOlkVso02n/oc6goK
9FnJxIfXReQHKoxndnExm6Kuhq5/tLFrjMssy05uBqdY6LGl41V0qBlT5MwwBz+6
/RfHgIb7cFGzv1xBmRb+mQsUTxWk9YDZRznlWC0qfKIRyvsoYlOUGcKAYj0Xj7Cm
iW2LM3nkdUPbjtiMdmT3aNuvG8sKzdd8f88piPaSszq49ONjamXjZie1GDkU4SKg
KUSXhpuZ/zxFyPyhso6AbXLxVjgUtjdkONhXXHA3cmqTS1U8K4cDJdnvknjvTpLD
gpBNPlkn26Zk6DOuk5neWy60Xn9ftezwMlEamp8ngjZ5XwRAM4eoGO3U8c+CbrV4
f7W8EPxy8nr4le0spJ2gupxiKHL4a8SgEf02xhCT8MQqGa17gQBlCfVbe7CKDcou
Jl8CEUHU9OX+o0dHeD2PxQLjnm+qwnVAo28i263Q1pq6EN70HWYxAXgIj7Vt5S6U
DHnFidMKN1E0TQ4WE7HJXTm3LSTHzOHMPxfJYFm0bSpohPoJTBLNcElKJAc5oe5y
xdTwGjOcNQ0IvvVtJ9bIFImUiRwAqM8M2j8b1eDIHGZidIhaFToygmWF1QqOG9lO
Ni2tBZOOPTDzV00+zLofa+gvKua/0xGily58nTRe/OshbAc+FKll8+KIWBvx6bQs
p0ytfkDtRy2rx9JS++b0zAlLjUFeZ9GZFC6GC2RG7rAoUYGjildQTDzy+/2JMwkt
rzNxQWXCROhfG5iu07f8vlGeWWYQ/ddfMGy47P+8E3UBuTDdWRTbkQhouWjXS/yP
BxU47WA8E0xwz1M8fyvBcIJHXVaiv8Dm2OYTZlvpettDZc5alu/jIlKo5KrxXSoC
8vdi0nwrdBaSlkCXb8LSIXyH61PBxYnK3cIakbvfl0Tz1fCYGVeanE3p11VINcEK
ubhjceJpfS3ixy5X0FyJshYL0MtHi3gQvbN+x1oSrAKtK4/YlD00FjQrqEkbuMIP
pp0IdKLY0W2x4r0ahPl9aG6HT9N4ExcRITe1SfLYbf0XkfU8jz1Vru+zVsiJSHh1
S9ttLnlnbJKuXU7q3b05MV6Aco05YrQQgTAqmzRM8R/lvRaNTX/iP4SDapO5V22R
GaaR1SaI8QDzLga6fjqn/zKoahGHjtl8WgvA0+HCW1IB2J1d1VK7pfcyq+WHYWPV
9qVPhFWFvEWE5LI2tcndPQbA1JoVPWO1r+HSTkQQEyKucOO2U4u3cb56BuCWIV0y
7P9gfnqCGdNlDLK+UansV88rmRlJgNniQ+/7UhdcwwmVk6E37ZBER4Xxk8GBIMQW
sJwk6iIQG/2AA6+2Fbkdun92mivSxEoTFUmixxVxsw/W6qCY6Oacybc79egHCFTI
uAbYYVvDq3SYK1VSe7dZJXtWq2OKKo2zxNBqVpnFX/RtsQ/mQEzuIQh+rGCIZdYn
vhcdR4cZPZ7Uibext0C6rqPRWNIk84s8UnIBz/2pXq2j4Sl+WS3A7Yr75YdKfZQz
XD/HdWv4VmK0QJ1HIdMsTag208S8IVwKSXunMg3kYFzJWpil2EQiZ3ENs8n0S1T8
PvWed3bJDCIfaPP6p9iS6YmLKW57svqJnBeeQsZTU/tNYEoA9pqN3QRu9veUjutR
Qvk0N6bOzGt26BAAzVpdQD4InQQzNTKb+dGakacWSc1DnCQNxlUzIwo7EohjnExO
5NBJmmCSsSedAD8R6Jxrz8rAZazpILkfrGxaoNfVRZ33FA4CcX+wJXu5CeWGIyN7
a/VJnr6kTtG6Ek3zxE7DDeiHP6T/gyldJ2gRJ0T9PcbQ/4c6up3KotwBZfATk6CV
ptA9bhE9/8r4Kd2caM5JNplWnvt/DjB9keg5xA8DZ67HpTXS7lrWjYa7qnSG0mTh
1qvmQ4bV4pnWmfIL0Svg0HawqZX5K5Xa0B8p4ESY59G/3m07bkwd+3XT/V9WjRqf
nboQmJM7BK1gg0zNxRakVSp/BibcexLizXK4EGoEn8ZoTQBLNMcucjrWj089ZWWE
RF3K0yWMABWxkIXy5fm4P/QMLvvJsiVGw/PWFt1+HfNSGQroBn/fsGVqDV69Dsoi
3sCHLfYwB5paCgMmRBy/19I175MoZvxmbfosbHbLqMeSxhWwCaDFazSC1ODBSR2b
WNlcW/X1tNlKoqTtmkLVeFB71WRinmxxNJaWINecBD9/o8fHMgFG6jNDnF/p6+pQ
X+EPqoacFXUR77RV/fnkebRHlUWQVujPZ2RFnqmUGgFIwVax3mxbP4CR56CMDU2C
JsddxKxZoduy2sI5Xa3TP0aL8WQq4AYUMRQsSY+aF0v1rvxfH2mweLd+Pd62t/wK
z85FsytEemh3BBiw7UnP0nEzD6JG/0vGsIAm7am2bmxIt5bpvR1n4a+YeyssbNVw
nk/BuBkfQJTdxYZ+xMAT3HtAund6izuBNXC143uzBIRCgNRrzVFHs1kvbdUe7HLK
p5VqREse10W8NeITlyUUuBY0SmklreO//KERCRBqcIKqPUBWsDDjmmRTD/Ev/ayL
tADc8MviNK/DJ1c1x7MFVJnR8rx19qDJDrP74CDrSjFlhnw96rlzdCfsfRXrU0cW
iyLOS2xQECbTmP7h0eKGYQlZQI2LzBRp80HV+WtKtd4ZW5Zgueaxerd7yhRZahq2
rgRySA8BmIOkHUm10K1k+oWaBzrMhKgbX71PLzeViclzBMkCnN1zZAb/IJQD1huz
opBNV0cLu4orf77BxfYHN0oP32n2xGO8iCgHMy63Trx8JjvAiBc6xvUkiXGmfir0
I8D4KWMFh5oSU0ZquhATr2IY8zz2Q9d8bWv8SqYfUb9PoxOOzKdm8keGA4eI9dAI
9yQYOEFjTtq3e3g8fB9tv/tqS43f/Obyz8xR7oWx8OwzUNNnHnlFhgWqEadU9F02
F1OCrRbtQv0jy/TIIeyEZBBug+suEwf5PzVO+ggloNauQ8+x6i6gvhjD+ODYhvt0
xqmf9sJEYAyGL2FzSzsY5d/zrIkT31LelM+6cteUedg1UwRvxu3FDihnTdgDnNEC
izheHicjTmo0HZP/58RpfOO9AbX434ku1dEu4ar56J0JKKqEhDZ5Hp1hlpoji0KC
eaKAs/NiHAaW7hKIjawjvnNLNNRTLEfrnzPlLEdS/J8=
`protect END_PROTECTED
