`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g07WhgdxHd9Aq+LQRz30CPnlkJfpHcLXTLJ35+VSsiPhYvJ/sf8VH1WQupfLrQ1M
C2zO5ZskLRmgPXzaoWIRqYVxPn82yZTx3VHDJup2SGsLWojy15wmlbZGrMx+J9ED
s7q+Nwonp6kfVoGgBBIT33/AcICDAYxVqUKecwA5DOuqYUq5b6SSu+xmguEY8mCk
AOY5k010UTfE8YopO0SdMVPFcm6zDbnxL/tZLpiQO24pTQz8cGRJJqKQL/Bu2hHg
FMIJlZrxQ/d0Z+KFevSJpEx1bvMDO2BJaV93GS1UttZDN37vJCqNLmeYUERaw6xN
P/OoSdnC6x5lY1nz7nqUoci1kQ4TFJ6yfX0hgaPYeePjpkioRDXL501wGjwVjOlh
plIxhW8o1QFifF/sbx37p5Gpc/o1C6i1pmm16ru/dSvYAmudpvDX+h951C8kGWiL
6aVrHWzxrg2fBxfRasOHVghdxBUh54KF86hVWEcx4vUQ5X4vC21Eizt9NnB9LNho
6wxpIUxHdyGFBT8rPveUsws2L2XUS1cPV+2n8PlIJ0d3DNO+U+1LwkptZsYkaAeA
oNP2m3raaAKJ1I1lhcr3CQquOALIyLUjwVyeDC5rqRM=
`protect END_PROTECTED
