`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aSui8G+ajOrMypGIt2DAYmbxa41TrULEDXrRaYPs8pLv+dJscZxD8b2jLFBKp4rq
AAE9pXnSsQ3/yMkyB9qIlw4d0bJ6NIiuYibsI4EaCGBMUmToEWt/O/60RRQmLtbV
dQWHMbWgJ1IuAgm+Hk1+R0JfeQlpywCaA2a+Hktkt7+BNpiU34Z0jKcyJgOZwcMU
fAgPAUXpteyYDuYr1dGIrgjs2POAk9ngl+iI3zifmIF0j+2EN6DycW4ITIznxgQ/
K8gs45YEc759fSiO6TcR3B28fW8uFtDLLM16Zx2zthQPAqs2YlfrIf6Ld6yq2d/P
C4K8D+4cVxIQqnPEZM31fb3HRUjkx7nM8Q5d1k0d1nLGUf+dpIp+qkWstCpjDk0c
5Lr4phizZJsqQ/bbabkqtV3nxu278Y5J0cOsgH+sSzw6f0PIPIpTuKIL2SuuONmO
Ynn1j2K/PBcUQPcPHclKuoT1EaKVY6qrTQwu67k3+haiyKTYadLetmKrzC05YiYL
`protect END_PROTECTED
