`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
koD0/rzENoQH0+vQHyxy5P1mmxQsTpN3LxpnCW89jKuYxN7UssMj0r64KJvB56uV
58uNC+v7DQecLSj9UQtVJYVe5mGzzUjUqR39lmApEs/rRb9XUTkF/MdBlWPeBKeT
RI3bPXQcX/d/wfDbvRg1AOAVv9WH+DQbccLbKTG+GHAi92SYeQajOQBaaz2IPkvz
9xHxlz2Lz2ie4f5i0t/qxnLI57DrQ922a6nkl3XrUeZP4mBJmJTIDmYkfzlFtT7s
/wH3rK+TnrochlsDxKYCsmKcvCqoiNVuh2pBCNrjiT6VbTe7smh0AG9H2LdMSFD4
biRzY++i4NhM+ZVyQ5+gHlWp3O8OqJiV5UfOsFuayxwLtfsfEacfPBuMN9d47Bet
+6FLpfFc8Gsc+d1vXvG1soWZgI/Ru+mmcjVUJC3eKQnwF/6zPEHPz/yu6u+wjVqE
SC3BMb4z1ONFDcS4opbrraD7BZlgVKb8exHqPGY9MGzWoCYrb8P6UiUpWR//HI88
0qJd4KuqCvIkOYJpw/Ka5Jo6V4pyjdnMD5eR0uyCAb824eacVynQUePOPMKYHPXC
MGeWAOqOM86PE1f/1Eh+FVBU/sZi4RO5S+mVR7N3qLC4cG7J0/ggi2eCwOJRNyyI
DeptN+9f3eOC8leqdcAI96jng0sIf3aWa+Kx6ISnbTKkHoSh4TrbQFaVdVMaaq2I
wDZKBFjRppRKUMuyE8olF0MTEgrLOfhNlkkgs/G9mOrsiqUY1JVctu7INlX/Iru7
1+lgUjUBe1ViEoeHtSQmpUToyhGP0M4tsM4YyNbBTRVio18BfMy3rzOekUYPmhsd
euwU+lVakh/YDOpfMetgMe6MoIJO5wU9TU/RhwrPzn7bXijQdwmX3L6iOmVVf3Ng
67OoXvy7SCUg9pCI4rJ0AcuDkIOCT3sgj4+ZAdfbbkKVyb6NBzF19ID3VQT18XJU
bIXU6igf+PEJUOv/fx16lD7DoqMsmnoIe261bxBG/AjnF1tlv3Y6mOspW2Pxu8/R
XM1vmKuTDGHeRKMSKUyNdPYKDezWHoWW9ALrtFfLteIOkHLSu/371LIfULjKMjnt
kNb+7RX2lfTB5zQCBJuWHfBWwFjAGr35KWLerGMIB4MB5p2piEGLe1WroXH/QMkX
DuMqHJFMbDEKs6PTg+L0sVPLAuhm9yTURIOeUYkaysTxT0yIB1YgGDOZ+VsyjnfJ
suYKh3xhi5IZ/8+wRXWDQGJQ/1Zdo7vfdqVijcF550F7wFOwtt6hS6PqIlZ6sLSl
M4bCSJVv0nE+Ud0DQRoyLAxVmtB13W73PmQ5g6O1b/9sqKwisSlCK3/RPXOGK4b7
t2EJCuEQQJIlmBq8vs5r2pU9cRD8XpUK/coNv3d7QQH7UTmrTlf83QV5OO5zQIhz
C1DXWyfPFPBy6zjmTtc4fXlSye8S6pdgRfRuoe6cHlz2ZvC/TiKBOUngBencJCJz
/qcwq3I71z/adM5wKHG7mKq5XyjDDlJEQtMArqL36h4g3Z6TJYWd8o6BB8aJFJfS
MssRYZQq/204I29poiehiJ6ACxNscgBA/neZnwFNX1enGy2KT+mQVHCv76CzfVZX
fWJrZjFTN4dssVScNIAdbyRYvQxNXbdJWqChQNjIsxwqTHVlIdbFA1uG+bOvjImo
H5izsJJsB3ocgh2vcbXOkb3uOP24AGw3oFLAUlkWLnIDaVhSZQdHmGnQfisgo9jS
MKoCG83D6F3MxgJIVxH0ASwl8srCVOUsHsHqaWeY0aZflaKpF1U7F9IU9SRkhN9H
GSbU+k40Yw8YPc9vWGlpFaPKQ50Hohlak2BOFIqxHXP7RyoBhwfNDNwktQ0+AsVH
idmyy39HsRTCJ1S541gxeTzYVCbjFP/bvMGVTjH0YIMJ1A29I0+aYL4oMydSnfat
KHjyiPi5Mkdm+BTQDSTcjYlZA6Su1+pTROZJxNb7rBHUIABqMALbFHbIgRKf1FYd
e4vnipbntwMNbI7mkyTtB83+c7l6UvOpMuRubzVOYmViPUCmuxHdwWmEICFVp6YV
6fnp58dJkUm3mWCT2C2gaNnc/0hUAsgd6q3/zCcUFtjg2qof6CKsPGJLUvS4TwMi
Vy3z5U0STGM+AzIAeZLlcEsMSP1lSYTERFaLqJgjcMNIjzkJ/h0ex/EAH0n6UwEr
qPZhGv+umAu0EEkEnbANWHaEUCxhhJY0ROCZ+cTHRH1sAx5FUgYU7R46A0TR28kP
dN/5YBMvX6OmwPR2FW524eqQxNJRBgLHyfPE7WGCJcIvK69sKxrY9Xdvwqdr0UGM
bMvcs3F31uSFWawE0oHpUo0w4r0TNJJgfvdz4FYyyP48WM3Zx+vxhjWwUGGnlO88
rKIfJliv/tSg5Wt+k+bwbeUTIHREHbZP0Csp/rPSGjb4WFcSRYTMzbHAf7gEBXgk
wK1NmORCp1eLgfpXh9LQz6XFS9zGArxBJ55K/slsnXOt8fnMLYP/ugb3eYFJnMHj
WdNxQWIX+k0EvfKXuU3XCk0lfLyVepjVEyRBTr3d1ZH1UMfER10hgGR2yDU6eEKZ
mA52XFh+qPp//73IwhEfDByGcHQYKdaYeqpEoqFKuo2uFohGiR5potjxLLdmiXwF
/Yfc2p8CAQH32aeiqr0NO3a2jekmipLnb0Gy+04+766XYhRoX4YvA1KiugIByyoW
XKtLuFPGjPG4sP3NMXQWovNPOGnL3ojyOup5y3OlW0A5PJQkUVxyxguG2zPy5I08
REArVov8RILwliH1vhdTeGSprp4EJPIMhR/LXFDaXVByLBTlIx9w6JHwzuqycz/B
wiKpyuteykGwtVq7AsMv/WDTYF6XWCqo6nVkqJkXu7EUhXkHHypNwzDyBYH4NfAf
WkVg91O7nSfMCElbtzi9k0o0/VhEFz1wfulQMC0cZhIDNnuJeVJHuyPiVg0l/jaN
mGg+fJOXKDDXVjA4zU6QXm8VHb370r1tN8AdYWJjXxDIZgbrewTxKJ8dp9tuRImZ
OOXvdiboMFOORzUSs+KNsl4rm2BiornecZpkm57jUwDugPBh4z9+WpxNdFMQjn+Q
QQX+G7oF028undvqMWkvNqm3IXcKcTkOz3WZ3ZFRxqnlxfY86E9LGjNxqZmJv1UQ
InquhDpimIkM9zP4GPxXoSonD9+pP3k/9WSZjX+OBlqNK+kZAELqDVVnAQht5QOA
Rw/JcTqoEGNsnTTTbwkCWndSYW0FUXkbLWMLb2ihhl/ZV0PzU0D3gGs3t2jp1AmA
xRcLM1oAbkRLnEDzZqcfErxSo35pMypw1kodVwV6DxAowaP2ZdPAbFokE4pwjNme
K/M7xcLdk7mkEBntHssW6J5Vd8tp6NYq11Uc1zXF1OJkuuwGjqkXJf481Lq0Dmyb
UnROld/wfsZMcGHPXXPluXm9sjtc9/zazqPF29MnT7Lg1viFhcu1h8h+PQNPIyTy
gZSnnMF2HGu9F8H+PLRZ7NuVxkyIPrarbfAaEhGRy+SCtf9tRb3x3VtY5p4sMzpT
DIS0jl3Hk4+BC6OeWv/P5DQF9QzF3QlvYXk0efES9FoqnUr82xzQcsbuQys4KmAU
iCqrDWvyiPfDvPrMZGWu65Ipqhyw6o2iWbVJJWtBDczd5msdcFmX1GvQMwtWGDip
aX2zxHPQV9W6xvspwIi9WWK53389hoJcwG3Xpura5Pk4mhML+i/uC+hxqyO6N60R
wqn4TZFn+0p/0WrfjkEUgIj6oOi/BePjZpW2C+ML1Y4EPmplMkrgju6/GTSOFGI2
mXwU9Bd/Dlk3JDFQ0I51X1gTvRqzi9EgBWQtZuj0XdBtOFTUL8KpBJnBomYNPCrS
XVf5ZMzUmucFaw/6ZRo3KmWAlZN0JW/y8ut0ZLAR1CWNhP+Lnx7qq83St1niCvK8
HyuItVX5LODuGydbgibZvE9/aRqwhoSLIneQssTsa0KxMI+kMpzwzcTNKwNdFC2P
wR7z3xGlrsTwBZg2xXh6pEZ+lmfwzTJrXlY7sTLsFkRWj8vdD81Yom5QM2UragqC
eU+QTtEI623EHRkfRO3kxJ2bJ58nPbbxtnzTVOL0kwDNhpr909imFgm9APFu1ucy
eAkO+NNFxUrWk7yyJtqpheIbgwxLZSjMb3kzHXgyWAlXdf0zj/AHhrrNEdg0RaD2
jjxttokyUZhtEiv/IO1jZ5HCSNTHAPbJWEJo2rk+f34faV2PEPg4iYfuI9LLr7oP
AtqemXcwA7jd0KE5fNNFGdkLb9H3pA5Pc89kRRHvnqXyoZF7KoOqnEXU7SoX9TXi
swD7eJE4gwGSKryF1CMaSkxDt7OUhLoGMCxSbWA4iiWCwOySBbzaFwxLI25/mn1K
y6u4+KpZCsGW4Qv4WqAw9bsRnj84nk45uCjsZNcLCuf4mHCZdv+J8ikbTe9fu51L
GeyQ3YjVlg/tbDtF50pyBDSSRwOKUWjPfBFkcCKPCp/dS5+ikX1rVAqjBFs0NOgC
c2mSoqqjCBCPt5MrgNiYJd//Q+BCJc49dp0EgTaWXvSmG6+XQXl8x2XxIIdMkfeC
oy8sePmUnKg0VtqFiBJFz//RbZP6bzi+QYHhGx4gXHnqCSQF2n6gChqBb6JRmitq
CoUC1RNzf5lxMCPQHOvmrdQj+HJXaMab3Lc+cNrIZ6H5ox04cRdh78/STvBQGX5U
Hhpu/wVDO+MP06UnOhQWtRw4ilcNLaqE+VPmHOflNnwujn6J0079isPGoOyJ1KtG
KvBup22km0nePg74s5LoIcDMY37JklHcualqA3c1JtjDHmARrVTnX8G/R6zZXXjh
6OwwJQwxLGi0L5rUi9ubJln+oFbngApOPtX6jlzuZ3RLjTNiTfbpHMeJjlM1jfXU
v4Buj2Bmfs6OPvfRMrxVZtQRV0bvbme6eFxPVCQU3XjezEUa5F34yOHgKvgINuZt
Wbfu9PizPlGjkW2m9r9lWXi5f8OJxI75cz48UGWcnUIBOhLXU14iw7GmCNUWM6e7
qMBLCbeWIuKbu1Zh7mfzAR9eASL7wSFAd2QGraehEFVciENuCPyGDR3I5WaHB7Vv
OFDk1vOqlemuRCA/GrL0rGaEvZXVn3KxnEaXig0SIbF1V/dZeRMdXzecnD85bIJt
Q9CPDMT3bxYVdC3iEINq4YSgOiotdFDm0PpawJjMlD5c/9C9dFnE1YPcliSao4YP
UL1oCQ7h1L1m5ZBPxxf90P0ODb46DV04Si2hoYaxKvSDfvXIbMe5FJ5EbiPcjROk
bU/dBv8yBLomE1pYyZaRPLT1Dfw5zcYIDFVT1WwhxQwVyNuAmyr7lXwciildXjOU
+uUyz5OLhxuFJo+V9BqU36y/STWBWQI70dmJ5OuYQMj7YKj60hvXarpoXmv9XJ5U
KkQf0VffQiTRUM9N8NKd2FaTqwgA/23rISU2K3/YiCPyYCVp5I/SkgkmyUaUnaW3
PpZwPza/3YJ62O0/x2qrR5FAHdcQHwDmzQ0jL+kHqYCCbkoe7SAAhgYEyjUu0dPr
Wa4eja2IDzFxkdXpcAlOI9Pu74R8Mb2yXEeUq1uaDXwcuAJwIQ72vy/bf4TBrum7
joQmYwj5NvmY56cb2EIEzCZNKxODt2ugsGWmJ9i/hq07cBmTY9VZ99fas5N428Tz
CLDvrq7T8kofjWuTlp/UjOASgYmNO0Y5exbNBaRI5CTR3pUytwpre6zhDZF8bo+E
X2OAR+r0W/SVT52WujF38YQ6W0hbqyOV6AMVYBpC+RT1gwDowziSRJeqo3aE7lJl
aNqgTdJA4yP7D3/rpSu6J6hcemPCpZ0oDXuiHZ6Q9ZEqDPTjd+I3IGAZ2O1BbZOy
fw8MvXCrN6ml1SWYTUeX4yCOiEsj91JBnsEbY1+p3JKwHVFw4L5xsHexWjqcQRCM
E5KdsQtL6/XCNry9IKE7Hl6EuROjT7iMePL8X4yN7KvMALF09wo5ZlSE653fVBjv
3eKp/LTb2fOmuDt8sQRb7HMjogXg85hS/YIKNBAc10hjECo8YT0Fz6X7udzQ1G34
YHNiuY/HCBskGuox9T97XRbW5td4OVoLzeQq7uMAiuvp2LA9pFHSvXxkSZQvgOPn
Hp4sKmmFJZlcISsQ47vCS3HyJmR8/UjUFQ+L0rjt6rSTMqsXgCkQAB0OYkAekVYE
CPbqW4Aa6Cz0ec0KN1rIdnoqkn1K8vgncSV1cqwkc66oVNMlIJKRc2yPqNe9mOWH
jn/dOqp6n/1QQgxjjARDgYKK3nWsHHa6rJH3WkUoQ5zaweAaLukhD0n/GPpOpNnq
qWZSR5idynJTLiQ1jE9ej0N1e7DfDDQ/EmvCfv3L2fHnGh0cM82V63PL3SGC/FeM
7peHjQ4X9TH7zwdEHgwXbGblyWrb5lCMPt/t+DJjDti+q/jUlZ1wvTdjKwPsLsd2
8pV/Of+WWXbmiBJtDUHz7mxNPzTUZw7RVTOQHAYykwhl2QQ/3nQ+MQjLCOUvz5Dg
qOJIak1RSrn+yGicTlq6A0MRh/zDrM+1MzI0QPtfGCFCAq1sl7kmBsgx/iKYliVR
eg3dQjD2GlLV2Hsl1OFMJG8/NE8LYN5H+epHpAbPYB6KbNHuFp7QsrlIcS/Cf4mj
YYOlfqox8sT1WWOgygF1mfXZscwvvR/gsADJ5Ty17USQfH5HZ385+hdwzpcGlhhr
OMgs/JS+e9bEKZs4RfhGadSNPB9oeMo6RORLNEiWx0+0Qh6YTpJzznwGFtFHc+1S
0dpAy3OsPqkXJ64pQ8POZABzqMmNXMYXNEPynBCIR8NbikGd4x9N2ycaHH30bdnB
fKp401X+M+r03YI7v13AZX74xBMuUYK39HNf+N1dAo2ttKXGTNVcdiY7xHausHQO
vQDPm6czCFijqf2eCoBcuq/2iTugKXjy/kd8gl8W2uQxrPCkNbpTFYu1Z3O+g5Ha
ynnEb7az4YDpNIEcKDrxJ0+N2WZNlQ2Vpmi9Rx5zLCxgw0cfhczlwZMcFCN6ilzD
S9tpJgZ+n1U/+8dmoWXCEl0GAdVZ08p9kgBrt2g3XvbmFQwhkO3vYS2mNsBCKuz+
cc8TRsXhCfmI+HOHAmC8Nlk96uSO3/2RkAHT+CyKNGLKvp3WW4zAnmKQPI/lmJM1
`protect END_PROTECTED
