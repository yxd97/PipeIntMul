`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mScKR8rUKUqRyUQAT5M0TwdmOwrOgilux9Asvu8oCqdAnhusNAFGpR8AzCxktcbs
L77g7k/pq8bu6Lfp5oP1VrbZaeS4ttd7vNTOqAJQquMvUJMy9p9TLHO1hVMEtqaY
rAVnICRgrk+bdROyNGhB7nIXLPR40RjtSlHYQicCyIaLt8pzmFch/bJWsZrLV2Xr
/DC0cQYeELPeVZdzXlu680cGMAqu+skdiCljA3Ah78KIsJhXltslCkl+gL3BEDCG
HG6W3UbNBMb+eSxfUzr6tsCaG4KSWsL6D6p1GDpFbA3l8O2R58H+PHCX7Vhuc/a/
6VkSTQ6BjO0T+KVwA/U/gqca5s81cKC425hyH+phwUcMr7tbuiN+qrsE6f912lSM
5c1A3k1CpJKRvPYbTCbMcWzgIXH5smfDoShjfOv48ao=
`protect END_PROTECTED
