`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jf2197n4Md1ORfvwrQzvO8QF3ojoFMbqmnm+AZJuIgUp25FgeF0ySdYBio0fit0I
wAbpPdGY0wzTSB1gwGRTFc+1t0DXEvSswPAYieZxcO7ZokcS0Uy895PS5Zo13DfU
tDFmz1v6L8jj6OSSWt4xnOGM4DA3niuHYQxjmYrbsWOcO4IVSVywBxqfgwdP1erI
ICDyzzxVD2jUFbhLQqzz1PTT/wRJjWk8MOjHS4A+VynAR887vhpmdku36Jveh5Kc
o2/7S1jRKtDfNjgI4FNVI9JZ9PcWQpmBtc6faJogE7oLiJ9sy6xUdvjFDn5i4oi+
mJMi+Bmm3uTh4D5lLPEY7GQbhtrBNl73lwnTX6xyKRMpxxwDQZ3r4Xw0oLzfvnPD
TT+nrid6XsEVSBs9zjYvSwopiHY4v9pl53k/qrxRMwhMrKpjyEgn39Z9q6UuUhk3
xFJW4CtET6OiyXfzSJ9ebWRjsuaL67T0vpBoqh0u6ERmEqPIuzbcQnM0zeDUlzq5
k77JgOFFhfR5zysGZ8azRCJj5YyKGMdoQf7lqX+62eH1CmIOCutMWI5ozbK8M6KL
l4nypequqSAlwYydYzhelYgL5EdX4msuR0P25TfnuuPct36gw7yrf2SMpRNwTsSV
RZ3MKnzbXgGv1s9XnJkJy5hceuUGwCWiFWnBE5/A0Mz/1Ni5iotP6/pXeUfzLYFb
erszXXyvc+yi62HaLCEdjWL9uFOrG9Issr4gtKT2EjV31eFIYn92u0LTCAwUAfUM
hmUSnAg0EGnB2O98iVROKirvt7xLzZBudYGXfqbvt93QMHNiFymrBSLtw6LBZ1Kt
qqlcdW2rVUWEpHg8LR+JWbxfbURx3ULxuDrrPkZvD6/IA9QYJ+3w/eUAwwlpsJGE
V5Hp9TpTJJG6pDit2pzCYd3Jfv4HW8f4knA2F/oJb9Uk8cDw1AOuDaeHZLYtA9VM
U5H+CrpG2PzuE6kJa/LnmN2USojS9+5LoDXgSZ18WAwE/0wTdCM4ruaWNltvbreb
rRSvXzjrZPOgsJjnxWNKwncIHR4F9/eJcVI/E1TWClh6hRWMVqEiqtIVcy49Zack
`protect END_PROTECTED
