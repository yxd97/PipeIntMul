`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XcDGPutG9StzOEif7eqdiqkCo7KnDt03MNVIW0Fx8NvEk1H7xyDdDx2oi2UoSsdT
rPPC8aWkyg3uWft23MqYpzLUYRj0Q/wPT9z2IT1RUXmnDSS8Y0O7L0Tg7GuASbXA
xtnlwa2I7m4q0Fjl34EG0hi4qI3Dhg9PY2dfxXLbuAKPBVLnVijQ867kRumbTizY
KGyERIXkww5ffTAeOU4LHKMF3Sjtd6DL+prI/qdVxANa2oXh0rE/bU3XQBUtpZD/
uDHky2L+1H65phFZNWS46rIc5cjw5n2JgIN7NKTYDvgS89D/paE1euaD672WwsfB
S9e0NOeIgLIu1m+d7/Ha2UbhXN7v/yfQFav8x1l0i5c4HtX+tCNELJTJ67bvYXlx
`protect END_PROTECTED
