`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tBpLYWfJdOemTsYz5c70UftTzmQkeQVsZG34dmERI2ueYEG5yxwOTrsWV16tL04P
67LU2fh21K3ZuUkk9wXaPc8CW3ZzRYXVlSfRx7GCF7Kfj+GF3x2qEjlZRJBnedGq
oX3AEHPKfbK9G5QAKvrLS5t9jJWJrxUglL2UbyvB0yWduXFxNCs6QWO+6qhkEk0W
hkbPP79mUFD7GFrRqv+hBEI5HuPI0czdAUQHtQfsXCP+Bt3lhMkJTQ03jZbDaW/s
8GMotDe6L+kn9oJggM3ouBrBz0usVfMBZbXdL5jUw2U=
`protect END_PROTECTED
