`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
B9RALL3DYmh5QrAsARx0vVKT1h32dAjk7HgRitjNOek9JoOsDCDn1X+kkB/JUMq2
2gtFNktSrXSUz9bqo6aVRgRWWE7WQrvZyUqzxoJucfHWXrvgKw3tWrpfBcJgGMs7
adYQuaJRw7DXYZdo/rH7054aIpPR305lFXR8+N57nPJgCQ/y8KhBojRQw6A9mkdh
gkhvXZr+opb/dhG0CrebLBenLm5OMLuIHkqPBL5rrP3FICp0flxNeuTumrJmHu3+
FOs4VcLl4f1s2K+XKlcJVQM4Oqg7mlXYC25siE56XJQd89WPxtfoR0EkZsf5IpEj
NXLmAy1mhRv7IPzhxfbJaQ==
`protect END_PROTECTED
