`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+rINCSHdFgJsKaw7v6dF/A8Y36v9jLr5EWPtWoHIXXSJ1NfTnuRlaE1+RVjYM3Si
TaoOaEdIN4B8NPhXs+cTQQRYCvxMbzcpdfwRUiVSUVxrPTOM/wew5RVr8OjDJC/T
Xo4hfbR3Loog7v8F1qdDt61W20RYl+7A/7tcsAGlka2QR4LsuPSZd916BP3i1i1n
DUBaA6NzUqILNM7KKuwKs41v3AbNgmiSKqJOcqBMGbyj3pv0N4qRFzif/3dVbPzM
MBQ8zizYfoKirBHE6vVaPimg4rHM186pCTxNAnCLkra6HEgwiA/cWABfPEMbvb24
epivW2gDdUkqkPcjn46Agg==
`protect END_PROTECTED
