`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0HS4S6MviYx3T8KZajAd056oq+NO5cIHi+8nCpS46R+nv48+4qpqIlBP1DWvIfqq
h+86eTCzv/M6UXQ81x36bumci0jHQIP96Zz2tW8ryTYH5R6nJpyIJ/jkyrVehTlr
Qed6mTEKs3GqptkG+B8kpCru1bSZCT7fjro5GI4HKgM94+PbI4GtKZKO76rSH0TC
9ytArRvvcQHiXVMsrdADiCkonPlKOph68lk+IXAyJafErB0I6kl/HIC0CAp95ebt
A1goThm2muVXH+4n9gGFf1WnGX4leoKbe24fqcbO1aoFJwev1yIOG+oOZ6ee3Ric
Az24YgswGx/kWW/do8M+3o5rRRCtnF93v4cU5K/nL9a2nPBHSYKvbamE+KCM6Zdt
sW/akXYBnI6/SoZmPd6Nk7uOdxJAhnScGunzFk7HzUg=
`protect END_PROTECTED
