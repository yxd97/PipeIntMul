`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dvEeiBLcHjY2Leby5XqFBlbLUaSYM26haVWvPpigpCtPTEvcSuqzg/1fZlzdVCTn
yuuB49nSfH95+A09Yud30WfbLTa3CKa708Mnz+jFc/s3HKECG9X/baGo4zzydV4a
/xfbXwFo2wvQyDPVyzvNOMy7D5Nkt/wVo4TtH8FSr2aVDpffTDt8t+k0LB9cp7hb
HJgRf6inyKBVnjRvxz6Ie8A/mYfbhguJMejMOwDO0OknKWNiFUItqgukKdlU9Qhq
vqRNka4AlqiZR5vq/EnG5P3PrDa/dswf7/thj4xAunbzxMydU4sbbYdRPoXTfsXW
YnFEpA0kZtuL1RjVy8SPkxMdgDtPVvdCC1+AVK8gIHOIbEtaSqL+URc55GNxTkT8
EyjlQ5Sk/rr2u9+C93XLUS/tdk51crqCDlfgRJzCtwtNr43ZOkhPcboiQMem+PzH
hiEiLs4atduv155J7qTjejcAQfkhc2g1MVBckGfy0YyEwsaEy/eW0FechQvjF08d
8fMGErgTs7ivkc+ibeGenv636n++lHmiDwiyYIEs2GtGZIrUmoJmJ48WcUy6mdTm
GDgEccPBNl8RbkYX1WV743+IhMD2zTVml784T1pxYqSupkulpMg3hQAE9SxGXv0l
JFabCJrBiVEJ4J/aZ8zLE9CQmk6n8sL8pNVClIQjgzNnqzCd01xz+Di/zbKqjMrE
`protect END_PROTECTED
