`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IhxogYZmRyzO59Tew8ZuMn5N/ylgGOtEtIMCc90tFOKt25lrldtodLnhGZRUm5l6
n+jaagZ2QJUDizPdJ5REWeWY4j9iM3RJkx9Y4DTdpggj2ZWR+QV26M1ZztAHz58o
L8kNa14kzxb6IgOZNaUlddBRjUkP8VY/1163R0iZV+5gL2yjCWy5MIirbVjnaUMU
UyIvouvfO7/+tQopUFwg2bfypzvC/oSiylkD3KTzReiuahQ6xmg1cDgFfxEGGbyc
9zjGgUkbWcpytA0fcEWYPIJECHNOtgz6RB09zDuz46i2kALYGgu/eJeyHKNujsEF
QiMOc9KZqjv608xsgID1BEiPfHYrjzLsxcZ6KI04REUQnhN1zHPP2oZGaFP0BARM
toNLAqRyoTUaXmiGr6ulnClknIQX9PM77+DRFIP1jVqvaUv3VLX08kneqwUT0GYp
e22bWym4pmIKvOqL5ekn01wdr8gTmxfoU/aRN/uCLd8Qg5Muw7ONgjEPzjo8RhBq
rRvnnJYs4lNElN5oFVF6ptx2rl97sxQMlYZ97PA45byjx/VMMjs8bTtSI89nVHzK
y9IUxxVpNI8fFC/gSyf1Gve8ONh14jJ7cUAkpjSFbpFeU9njIYfWaOQCw4UPHJDS
+KwHZt3pPH/b/RTYbAzcKqDEbGLsHwOTuav73bO+FXgnmzuQVjo+Lhjy934NRUYl
H6Y6kXfteK5BlA9Yqy4E65UKjGwN2Oi/94I7/pLfom2E1JtTELRChlLM33v0hm9A
nGX4SlN1xp8IC8Zz5DDDHYl3HAMk3CScNB8PtQ2E1UsVqoQIWmp2v5u0tr8+FC+3
YDxqwsheuG6ucA17bQCgtr0042MDERAwX/3Mc7xe0kl53rvnR+JcY8tAY7ChXd1O
6lPp5+4CpBRXzyqZrCHKxJYlrSsmOmmRmTE+5c1RpbY=
`protect END_PROTECTED
