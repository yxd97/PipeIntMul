`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WnqDq9WiZfqQXY+b67FyzTWpgoGZuk4FFbOwAP6OJNVuBUK9nf0a7q5yLoPQH/XD
rHHe+tBEq1N01ExXN2b4a4101HssGYdil5A/I2koSxUDcSJwm8z0vH0hvcZm7eVU
NmISomjHpEu3FGpmzCeQpaGjxG8GRh422+EKgsaPS2CvRaseRA0AzILR4/4K67fW
C6z6yL6CAu/IaF+zr0prwLJvMHq8/aAuSJHyK64/JKUrPfUgnuVKBWGZqakdkf1G
Ao1jjpBJDpwwPntmXCowLXLnIDXwAHQ00RGDyjMbBbHpdqTy4z9zFIlvXx+kBy3s
K7aUPAa7rga4F2yo57w19KHP64XPAraoZdxxsZ4V8rKgjJcn22Lpm+WiIZ5MEDyt
QWMt6+R7XqW1OzhLAa9p04eekZ0t8nl6v7HqzqKxc55JFjB1zC9qKZnppyJqqil6
cQSp/JCSa2ckFonNnBdA22nRC1GK5hLT9zf3Y18pJ0HT3fothRd1n+omqwDvxDgh
xRSegF0v8Pb+VEpJCZTvuC6XS/CuV/cOzF44nGBbVjD16MDhdGAFWoJ1OcloYD6F
k1QKmAWxJOJwG3I2N9avHR2DcvZb7eO1qbkKK+fDgkIg8ppKcareKcRMo8xgH4sn
w40l3Z5jc3QXLJ5PhED6U0c7/gYXwpqJ85KuImZt7UsGczteJ1Vi+8opp4YjWPuM
Elv5SGxJ9okGV6d1/i/n4ika2klpoFTMA0r/Bq+IrxE44+qavMi+QsdcPPQm6Us1
O1ODz+bKXz2/ic6HWVNRkQ==
`protect END_PROTECTED
