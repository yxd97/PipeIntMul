`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TLlR8cUVHKBKQTMs6kZM47XOeYT/MUtOtN/P6747SoYVJcF4CnSHt7/zW4RNrw2h
TMvtAMn0o3pc7np6D9VieR48omDmQ4Xa+SXMzpesFsVlH+ky6rbePxevlIy3B9Po
4bLMuX4Yro57/CZje7LIITARTF0Sw+yM4AhWlO3/8DnF5F/PXas+Nq4q7BDlNetu
GQwn2I9i8+IvJvAmLhALJqACosDPv5BxxCUYT5Rl1+CAKXtcE6RcjnR0sKgrwn5G
z6AW5t0qIxVNu6QslQC3vQu3SCh1Cl8tSQ3/FViNrhYcD/Z2Cweb3L1Gk0DaXHo4
xRllVRP7R5Vc0dHZkvKhr9c4HYceWWHmHysbipUlBPrRePblWs+DkXY2+MEdeooB
8ivVrQ5dDJ1x8u5hpRcUrBCGADITkgC59SfnE0L7iYfjKmJtX+GgCUNkpxAgoZ+g
LdtwM60r2iuyy2NPVYPxdln+4BHdrVR0Fj3LqyBSiuKUopgEeYkpl3paJ4n6W+dp
7wyFxUONKorL6NN5aaK1JaS9zQvLRIG1zAf1J5tmlZL1JFkZHFXryeA375ksSeRZ
kIdVupakcQ7VCG3aJCnzxs+HZpL4a4qBDAc4VOVkTx0=
`protect END_PROTECTED
