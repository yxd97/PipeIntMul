`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39/BWBiB4oZhluKVZMeEJdze24U6PeCi3CIhUSCkhvl3V19HKRyRhsY9dxA2Nm2H
mn4LJl1eSsHoO8WCFsCSrbdcigpJv6ZT9qpJ+kb3zev736BwF2HC+7EA0COuq+3y
NzvwkWbOHBbsu5oV5JkfTWfkIU5fIvM5eZkivcfFRDnRC5VZ+w+6seuITEMpLP1a
ze3xV5LCNsKxeCdc0wna/j3dOjex8rdNal4Wqs4KUX20ABZjEe+WGPcmuVzxEnTD
MBLGA1GHze3nvGdp2oh/xlNSwrQM9ku5FnGYodwJnT2jxUyp5PStrLSc6BrJUAkg
FvcfI506xB/wfoZ/mRg++D83gNSgJwnb5a6oUZJhTn+cu4jxT6Wn5ePCRgxNBDQZ
hwLgOSA9GNRZdvwXRjwCitKgHLvXqNgnyYl88FidKLAjenrt7rmBA9dVmLpx0pbj
u4ze7K61oMNeC9P6ftt4HipeKKNJh5aqLHjyeGbPAEweOTlrszK0ALlZTerQ37//
`protect END_PROTECTED
