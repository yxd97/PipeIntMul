`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mvy4uPXXEoNQe9ne0jU9mjnpoWxtD9RhHrXYiQb87cpefLnX/Ap2xKnphv7Noerv
lW/WpzhbsF7kfdqLNOfCEssMxhTn5VhxV3HyTnHm0WcVjPolu/s0wSfhJfPceCby
83Z+wghVFfKG2i9cT5Br56XV44IsZBHHA/4M4c1jlUd1KzeRAOzLZuwSMtZcWojw
DPmT+Yoht4Q87BnK6lUqoB6GvM+IrG7zdJA0AC2yOEQMwfZI7rmF0BQ4JkUyoP+v
`protect END_PROTECTED
