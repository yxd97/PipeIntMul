`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wkT+Eq0pLCMejb0WXiV5CcH8JgttIl+NpKonV+G4RrODuN5QHQFB5MyOEXS4HRuf
GtP/Ho9t17G+UdxpQEtpNGcq6pGtLGh6srOBbu5FOffsyiIW0V/8dUJAbjs9Jcrf
ZmU0rS6sUHZDZBOFyEU7mgZOmE5HbEhm8gcf0gN247L1F32dW5T34gIKXA+aUNQ4
RVhkUxIBvJpdwqiJeA4sBKni6YvhjW/qm4rIlks7wXoq91J8swOpuVXvrPaVjA5l
Ik+zQDVnKQTLiof+Ca9waiphFG7icGajloCvOHd9mA/wxt5sMiVGfkE91DlDJTHY
4zf/HWba37yw60ypVe7RycKfn6TT4fc/gomJa7UV4mdcOYOc67D0xkfu9XsKCsvV
zQv/3VxeVs1J1Qm443kq4O6FhJJBClQbxIHdaKt9d5yIHti0RXMV7Ehn6qgqBxba
Mh+Or799ym4dyOsvhCG65ELYK1Fhu11ORTtjkyaeNEkiHxh6qylfV6cYBBJd0B57
k7ztFBgtfc46gOFMvrWShQ==
`protect END_PROTECTED
