`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GHNZN2BNw7oE6QCOGb1nEzl6MkRpRj1P/bjN7mSsZekjoz8KfOoGxIKK5BZTGJC6
DJLJ5F9Fm0ULIjNsAIXh3xpvNZ8e0kVSr3tURmUxYKxoRk9t4l4lB5sh0ilXIE+s
fevPDUD6cYbNiGzNSHrCbAB2bVHrPRw0d4bosIMjlIlmAICTNT1qp/jI4O0cf1Mu
A2YZJDOmrfVhAkL0fpmOOoapAQWtXSuA3TJefyxEND51e5lo/yAJmdfaXlkxD686
vYYfUyJqnNK06wffNoUmUQTkA41N+M1WEG2NaSesYEGwM+VMSRzrXh7s/gtSNHTN
aPLxU9F47wCEauZ+XDC0Pqw9JL02r02cN89ee+Mi1EaY7SoC+bBpcgQJn4+mvwR2
cTZ4kjm52RH/EP8HOw/IHQ==
`protect END_PROTECTED
