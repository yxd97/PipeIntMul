`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7RB0ousXYDzTKHzjl8czlUwHJlf/CoXLcaXBGQw8cIDaPTbr1iyZYZnzp3oJmW2c
P4NdskZ0Hsniru26G7V4QitoaNirI1POqOS9636O8wU1sD2a+DJElcPH5YjTLo+5
C1rWFlmixZ+3AsZP7HMWMpSucdeHNSidE5qXexbGvKKJzholy7rQqlUOWt5dCNmZ
rkqSCRaBAAL2zGVJOrxVY9EtYHw9qiz3uTikDg8FoV5T5EThd/3nOYQtTeI6/4Su
gwGKGjgkZEQ9bW8XEmoAbRLv9+hrA2al+pJvo3gfmBnKsE6LLRz2AASCYTd7CLmE
YTxQQlS21WqSjt+NkotrnkhH5BlPkLfYPnRUjkLWtPNPpu/Ds5ihKjWCWzBzF6d5
sU25F7CE6UeUWKCPE/o9sg==
`protect END_PROTECTED
