`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E10wcneYTRzEO+ogvsMxtLHSq3QrY1qOleDlLkEbo5XwLNFQG5FMxQSEJDK/ps8c
LEIm9R9sP9tHMoMbgbgfGCDp7/8x1bS06U97KW8JhICfnZ6DbG1JlM6pCRD9kE00
LQqvBOS6O4UW/cD4MhE6NBQ80ZnmBrG1lQyxxzWJBGy5FlQiWPBcFN0iy3VFVa2n
EK5xYr7Ilj2ttxjypYSlqcM4tcAeNlHI4cKfDlAqlsREbCoxx3R9yGoQHVOcYO7s
AHyE36VlbiNG7TuYNCtJ5Ktd35CP5E9K9m87ZkVkTxlaFgezKbFQjP5xKk8DH4W2
uKOrqBsK4IhkxuCDmcfZPYPlicBv7piWhf2Ee3DEx/GivkVkw5zZTVgVpFlT9KHY
RNd0VWXuN8djxvflnJ5izZXvtCiGhY6uW0Dcn/6uPwxiYyxegvebCW/wGq1737VC
c2FhPcz2q0PcpBH4haA/m68KV3ZV/EYwRAv6OM8New6RtWerVoid/tibhd3H5kyL
IbwiVOrFyfjJ21a6vbf9c7I9nuQlOEuOh4PZgnVIgxOQCcIaJjGMcvdNG9mpUox0
mv+S/w0WCfe2ku0hSR8NU6nrhe06UuuYmei74OWajRgqrusLkQywzOm5+VqIFCsH
R42Tg56ZBuH7zeLjDXfr9w53CoGeBFaqa+PJNPNO5so=
`protect END_PROTECTED
