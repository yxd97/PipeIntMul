`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l7lMlso4cQUOOTd4l8a4QfMrxbRxrTff1Cy1E71+MtJvIaQhgJHWKn4PUh+YfFN+
kFNLXaZg/OyOuTD0nmgS63+7zJNeeLx+oE1Yn5IgiC544DWhXXhSQZGxPwHPux/2
NIEg6eqGOeLmem5KIFCFppMi2x/vo7UeEwwsDjAQB0Pz+WjJEb64ModCMsgQ+gAV
FyrvwIRtT991BtO4eO32ijpDON1/sdpkdCB/J65GlMtJwYtptUZImHk471dnpifT
iYLGQOxBmER3e/+I1lZcGwumbIbt2r9bvGZhqC1f0ol3z3pXwWL/KQYzC/UE/9VM
`protect END_PROTECTED
