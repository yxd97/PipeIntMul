`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rdp7UqXdDREqpMNt7nbyTEPQ00Cqe5OPAT2fkTQMf9EIkvlD3Nf4INERvAZsrkeE
9jl/fbQXWuBWx8M+rhe+FnLsf4cABy1gyeGZmIu4orsq59b6fzenlspisfUuSV0u
w+ZjUznI2etLGlOUsraJy365PPNpD9kyR6Y3vzsmV9Nc3MM5bMoCPkFgJlEiJmGP
/7z0FL+MAvWZgos1QDxqdK7cFuDbM7EzfGAOiJSND4E18JrctV1/VoBeq/qqvYCI
esvfRf523y8Kcy8XikWC8X7V42GBDP6AU8ouLOfoP7NcMQseet7EvxOQHKKUrVEe
H10q9OwzrxzLdHqWZ8pQ+mj3jVbC0zqz9oLOgrcazO3ijcRRoD46G+cQa/AU/CXb
GxiSZGmCeQ9p2m0tD+rAo3vusd8w4gGMYIpiMPQANpA=
`protect END_PROTECTED
