`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EMuL8YwL3DRboPd5X1SKr/N4Q/WL3kiQ2H7O6zF6zA455X1iAZESyLRZOB6+TRbd
WAD2rqIHvDW24HBVGIysUTrRxoDVr+UF6JQq/IxrmOSvP5IMLrh6rTaGM/ocY0RW
9wSeYXBBsvJJSNjnNkjuvXGs2AWfp8AqSZw/4le3+W4PCd0eYXdTKzWs+H5wLmEY
qx4hRmapJw16kMhCvRhpDCSJlD/bqKFrK0KtgB8xYE5uyeG2UWARBeUK7nbimtc5
gz2VxScmk+JlnN046Sljwzm+f/ndD/zp2Xi2Oh/TKA9R3joUvSxVI9mw6uwlv/F4
+9iriF5v3wCA4O7sBL6YGj0q9+1Bo8tTgFQPp0FEQbMIfTS7959k8Cl6jOvFqSJ3
+hrT2gMBgARqc4kPO9yuyq6YIWeXeuiFLVYU8HzdvF0=
`protect END_PROTECTED
