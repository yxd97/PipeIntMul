`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjdOQRwcQ6urjl3xIpU+G06UXzp1hfsrzY52f/vy/ktefRh2qdn7by3JxBc3j92Z
TQiBGSgvU9wPU51DhuwJbSqk3TadESKZdfJ8dxNso7wbL8QdPpbTXrzpr3o1I0mQ
bkfw9QsweXRLdeXM9AlU0eHx7rrUG5WmI156Z7T6i2SqJHyo4YRw8H/zxd2eNtOg
bakhh35Em8yZFjzOxvwizn20zplrNxYXKJSrd7a8OM9L7Gv12ASHhE1LvybowrLK
XHjMHTxj+FILx9BvB0RDk3k2t0Ud+g2Q7HxBEz8+NjAW3Fi0KCP2bM7YIfjjTxIO
N4SXxA2svJ1HDzR31QJ7zDNX8JLuO9Uw2tXIMxOVVC6E+hpAQdIl2o8HxqGa3GYy
tlFW9FnKznfGytF3zdZb9JF3JGObyEmKkB7DOpsGx3vdEzdz4EjLecUuev7SdKGU
CjJxgmSCYW1MIDp7W+Mkt1sV338Q5gt+p5CEWZaMRUtW3+bmCRy8sx10mOmDv/bI
8/u5nA4eSSz4kiVEytzJgl0z8DpEcpFLlVP0nMfbX82X0hUZPhEEYf3lWJuSgDdY
hI7+2O7Q5y1NT7ifPG7mn8R6f3tkk3eGDNXlEiRuLnoy4Dvufa11iJo6nRDUMTKp
bUhHaDrW6EUgs4DAdGFs+d7/BVMrGcYYgIaaO82ULhWyQG+3k8LzkSOBzhXlYFqZ
SmYyI3BBuQHoh9oamO1zVC/vDxvZpbf1414yvdkRhHcK/yfBRfVeTeFVwpOFp4+L
6wqbUAiZsDp7F1AVVOzqc8pcOaZKmuSYC0CTnhODQJHmizAANDaSH8T/xOkEK7Uu
x7cYxhxpAIvWEg5L8VNpVw2jyQM6GWSV3w/bLPNmhDACAClB6ipfklUrbkOTuN6A
e8LlAFf5eit6TBx2RmSRcZQmO9zRwEjEU6eE5qJglGcTGxfQXDex5UD+6safSaYX
LZYRyuYD/w5KNdC7wQDIyE5b3STdPX7uelKkWU8ESAMpGWPx0pgaZ7Ybt3Mcmul2
Ues0wCaIW1bz05vdYspYZV4y2e8D+43QnL3YGMaNYLX2dOtafPwJFRaJ36nbmnW/
EvwRoagQd2/uBOxW9a2zoORZH0GSGiM63YvEePktFjmggZWBGXz/9du6AVPrFCp9
o6ujtz+uAjeCyCzsW84DZkB1dQ0I7vuA0odhpQK8CvuURg0kDc37cxaqhR01ysLn
jRgv9r/dnFOakXzBEa4xQYVJb3xyig2EaCJZlR2i8/NMk3z21UXjJB2EpKx8+yxm
W9VVrn7AetWudKnNROi3X/XEHh0wijVPE9RyA8xmMRBhu6i7Br45rqunZ5SjoWpF
GMv/NAn/kTD+jAR0M3Z3LwjCB5Z49VPFKRiPxrZn/vGYNNy2+Ak9JR0hH6j0/Wiz
/Oswt+XIuZrA9W0Yg+o4FIvPApVJN6KnK88L/n55x70Z8YXANinmOe3MB6Hl6CPd
2abOTyckwTCXfFyVHF3TstEAf28OikONjkqY2SARznhjUztzVzZWAL/A7vuT7Hna
fRt3tcLGOwI+warPV8mjJ6uQgGdxWlOkXmhIlL0hj/5e3QFBM2Vzrz+3AiPsIMA0
GDMYC8Z2kwrvItROe9R+GnweCcxgS7vNO5jqQIipBXuKVzhdb3djln2VYSBLW5+c
iRoEYkDFRTddLT1Jwqs0x0IxbSJnX8GpGffgFfj8pai+S5YiZMcXBSlRrQetUmq8
bSgzC5bPoCs5LrDqY3JdEYbt0K/W40LwNXn8QOaHgePC/nvBNRpDHzy1xYp8zQYA
I0NlDVW0vX+ZJoGbwiI9NEpq7Kj6g0bG6qtaUNJoUaHTGvvs7Eu1h90YDIsV6k2a
VhrZaMM7Xfre2VyDUTbAkfYme1Dkr3Z0iQ/Ob4YhysqgUQhG6QUXLFPk6ssTkbKC
6YUTNjumQ6TmL1I41E65fKMC6OZlGSjkjXi3RWj/dvrkyjxhoXpw8xSnQv57elRN
CAO+fgctWvDdmGw7eKo08OLJbhplf0mhKV46YT1kCk3zILXGwZfQN6JP6zK8p7hz
1yo/KDfg6r8WMM23K9z3ZyUW3ghfrDiw1uiegYydLNQOKtL4/uBal/R8n8Rcfo6O
BQBLIIlz9VMXy6O9HXpZpV+npaU7FQq6rijcbDhF7y8eAVzk2L21SxwLasNdYK81
4freu3gLJ5QaVcOsGiTtks6DheOH12az0Nx1N5fcKIVk5eUdof+E3o3TwIdmmck6
+BEvjssiRbt15/AT6h5snBTJJUeTAfZkccmL5NCBmdMoiVH7bj3wmC3OYdPnXLTb
9rovn31n7u31RQW9ETg58rrZYurC75HXIyXGS2fLy0JIwGr1yBiTsMJQmO+jqGI2
9c7/RWVoVPeBHGevYc0VSt3RY0sshTKbKRg3Wa64GLzgGLqzqmo1WoF8Vw0u2pSA
mL9SRtOjZR6hoxorcf6oxqrdCZbaZBvsxaHrMz8bRpCsT9+GU8W9z5c1bgvQoq0C
MdpqMNj1mmvFKLD3aXkgmotJNe58HbDjpv0ZhcY8ndtq6ELALPHXbIRGNvaOLBrw
usbgz61whNMvvSAr2WFf+q6BWx97lt4/+0MBYGbQSq+yiv2yf6Hyn95VJnXiQfAY
11704UKpdeqxt0BwduD5vfJxy8OHOXPjgSeQgXV8AGZsyd11N6o/BsHDiW3zdydI
80ar22aKzW5xaQixG0xxY+3reICp+glWuhtP42G+v3k5efFfw1qkqfxLYwtK5hEC
T9xXHWTA2ZLzwKUmVtcSKBW/F93GCRW+Tch0sjeAVQkHHyOJN/M+DwLChVCblO4B
Y5oxM/jOMRL56gSpNXhhqrzjtgJ5D3p24bHrC6yXwmv1rENM94hkDM9zEkYcJbxQ
L1nppYgAfYddI7MrwBfko60ZRZFLPhpv3aZkD/WtKNqNd8n8i4K6NdEid6aoxzfw
iuGRaLGiv7U97/I4PqBGF4fLptAQJ2G78xaSkzjC1WGH1wg7yFJIdykoqzpA5Ut6
`protect END_PROTECTED
