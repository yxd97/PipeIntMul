`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZ97njP2RXfD+8MKjCgTquexazuSyIEU1K/9whUo0fTy8mXgry1W3tTxmdfNmBFf
X65GPdh24fV3Pl2hZeoxRmNjNu7+Jz3A4jmFRohdvesC9rSUONPE91nrMzBDAokc
0jU1YTfVTwA3Q7hZ1cwa+Au7xmbiN5uWISjzEFnQl686ZjU99fxywAbjPd9iOvuj
JMc1oAf5XaJGXcT03ORVe879UEeasxhdTx2CziiDc7SDvVXH9MSrOPKhKQxUZzAx
0bkUP1FVCOhlFZrLPnBUKwEAxzDMwA0VPshsDmdV6HiXnGfV18OPmjY3jefIuwtP
cOT4td0z0+UHJsQnHFjgUMVAfrMZoto66qeDJLE+gPkdkoKJJACo9irN1S/PgpSy
JFpfapU6qIY1651j8112jStffLtnN0ifEPvodMPeUIKQ2UCpORvWVeGyGUlGiRfB
SKBqRCTDxdtK6La4lcoqfHjV4aTg2pu5Gnkcp+OGEQ1/KNWC/CamejZ2O+4m6UuR
s0Jf47ynD2VAkZ5/f9/QdQCfFxHZZE133EKyOYL7MjMF11j9BjL6KwSItcpyJomB
EzwgL68jsgjJvD61tLXHi2Spe/5Cwa82SpBMGR86Azthr4YeDBfBFG9r67MWujTW
2OxZcDv6aHo6Xbh9W1F/B+LPYzFVyXDm+IShe/uR798=
`protect END_PROTECTED
