`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DFo5OGJT8Yn85ErsKdXDsbyHVAGLJTQinhD4GibABJPJ9eSY2f/WtFqIMeV5Z9Hd
q0/rO0DcgF/Y8tB4iRJKbJtDqS/6W6/BLkDWWRUUSm0pOMkp2mh4x+WxJ+yky7AH
of+Cn/CubgbphGbOv43wZhXVvoA2DfYRkyrBHxKIDjay/Q9/7n1sEqgOb9dU6R6l
miHEfq8kvK64dH+jaI3VJGz50f4l+8MbFHAA9UwSmmqPFkBi2QFWWnlADxDsIhu3
rejs2veIyKoV+EoqeK89A5aGytVzjj6aU9nIwptsNOz5HPC/5WMoXq/mBh4S73mF
kM0FNXpkQQ2bVbFzwPK1syhwoF8b3IdiqC7f5KMVzV7iJoTof3IEhKOQ4EbrPX7V
0nRJGuFNQAQNRhxeAPLkERYM8xNpX6Mj/cljSnKXC1UIHdXmzqQeWNQCikjSCVnU
ZPYzu6ECdtCsexXVIdRIcZothFWmmyDhDx2AdjPAxE4=
`protect END_PROTECTED
