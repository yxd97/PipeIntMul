`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KcR1oboNChalT/uVzB5STF7YfSQBvxVMPR4xhLnHYD1yEnR8ZPA4spxS+QO9epXM
4e65FFYxSUk3xloTy7vfuEOZLzu8Kz2MlI/1I+rr7PvgcUxkeqoWfL6v29wkhBQ0
vO6jJ6+wPjs1I7g3t5bHuQiyVNt/I2UdwlqZSpipaMQACBpZXPzSkv6Qu3g5CvAN
t5MVpuhJvIALUOiRrUGlibHmkgiF7F7bcu/HL5fFheG6nQPRGB1WeG2MYr44TQHB
NA/XMLgoqsOLV3BIKUTBaNTRwwTzJG4Gv6ytWGvLQI1Db/mDaVmWPyxuvkK9k9C6
/mvl9ZSAlCq1Ev+cdasPCQ9GzX9StfjyA282/J0ogQZx4BzTfqzUePb7iB1cVLdJ
NqkEVaJdbdlEDM99zuzhwE07nwCHb1gVKmRltuXdRPVRx9TY/4STkp5DTPHv5K6T
8uyjXFvuVpPcecf8fZnyn+g8zMLUOnwDv+3bF1Lfbqqo0ek7dLdz34qL8l5YdjDD
`protect END_PROTECTED
