`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y8mrPeK8wgyQBFiJQwvrZ8oL+AdpGHXMo0WgOSKHkFFXL6x4+NF9IaJ07vndu69r
Obz6hjpylVgHgJVDphKHsEVyTvMl0/1ILbqLxsrosry28BdOE7UhjZL6ju+wUqQe
XB6QAtcLUJug5sFf5k+0ioGKTHCdXhsDhV3dM7ESUmdQafQRF3c+zotvYnAp7qYl
k+aDiKdXo+fcL8+5xSUHB7toEGWs+e0Y1R2322xmyWZpJIwTAXVgUzauGs2f3LDS
P5YUdwpvp8HlMxor0oycvlMKAwTRuCi4cVK72sB7coF1EvPQlSLu4m7/Ux/xvtNO
Pv2HiWpvF6UNgBVfrcIgamE3FMsn0yMv1DKP17ghLi1x2RyPZ1hDhO9GO62iAayR
5aT9jdzEXk9Q1/lmxR/b1Q==
`protect END_PROTECTED
