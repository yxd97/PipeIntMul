`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
35L3j792oJA98X2iMmscnbI8kPGGTpkMkhLPP8UwFrWYbF+2QB2Bpsp/xu/kI6ho
b8yo73Lr0p0jEvz6+b3bNjTJDXOFUea7wPOjfu0NWah9Ab1PU1yloVVMPQrxOxs9
96MSyn3P+aeZV2v1tQOCdnM/OlCMV8Dm33AB+AE5OLzn6/122ydvVYPly1/Fwn+u
SmGL542KWJTA6B4Zpr64vYOF+cQzpGVyd+BYA9qGiAhYBCrCRhMQ4CL+CR6CbQm7
aHsjb5YJEsrPxxt612i22umIH/Ie8eVqOkEgIcq15UKycTPLat3fNMrIw8eSq1Wx
QDOzpr84lSXhv+G+Shn1pP7kG2draOD1RB5v0LaxzomQgiqj5d2gAhS3/qyZyy6m
DhMAt+OppFLf+MeBsRV3+F+bDq0/23LgLvzcvIdM6b/fz/s5gLo2lzyVyg+LhQqR
Yvyb+w8WBhC23WARiBON+lqTN+DsdxCB0SIq8kL/JEIPdY/yWNPsCJKaMQUyBWdQ
EEfXgdLKEbIruiuXPI7L9eLfTSVlsEDj/pda7bLOiIOZPeKUAP7M1HqDn5kT/2W1
zUY/L0vVHw4WqezPFA6woDzcU49ZDiSftm/AXgqpGmLHLQ5HhGnEjiGfkJCMhlJH
EQM3PRTU5I7I7Ls3w70KHIC42xREpISEymFC4BapmYfJ0TsdTjDssJYrJniC6M7D
rfo4xXwDETVlZFfis5EFgqVccH3GV1diH9OvWjdAccOCPXq9B4jz7L1WnsaLe2Ik
GxuYp/22UHVaqWMnsHHruQrsLqKZJ4x6DmGI5pfgSaT1UiN7XlKxDpuy4Qs8uqQ5
5eO1UNQWH9T7UUd2KQNH8g==
`protect END_PROTECTED
