`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KQq6WynPPkXzw69cfFABj9y/V+1+svEzP7/waT4LOTblAz1XGEwZv4slRrLOKpGr
PDONdzogsBgrw4y8T+wdtr2LXOUJzkPMf99/Ax5ACwlhBU9Y9q2v6g7UIiHmsjEt
qiVlnj6io3TnfxODkcL4BOa3wBbxL6XPyKYaSMC2FM3R0vmne1qw1k+eLZFX2IlC
cD9jsH91gKz6NT/mkcnTFkpfakkqCbGqZAhGDNVERFhIWs3GjfAv9oC+g1OZ275A
/NiFmuAoF3azWSNyEQ1hnnLmGFUU/q5VXw1mf7VbovG0C2woO+RY/nl6QqnmByMc
aQGkrVxzwuMgFfH+SY4WCOFF7qxaCseh0GG5jBnUW/M=
`protect END_PROTECTED
