`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6OgX0XtQz5/My+E7VxmPxHNq+COiNbkpbi4LJWtP/Xq0mwmWIi1sofPVP6oOD1b7
AEt0QSF2kirxPb2SYJ8ctsuDo7BgrLUdkXFrCStUmGJmdx2gdi1Bv7EzmX5XdeD/
OceqzffC+/7bLzoC/0s/H96iwe52bbmhvSMg97cE6kmCa5x1MAlhIHotSam3iFIZ
3R0behQyveVREq/k5Se1aif9CxzQqZCAaURV1J2hDndiPFZyk4Xx+Lz7DDQd4QRN
ZM8wmWIWSEzG57MDrDMkfoqe9sD727vMa7Hn2oAugYQ=
`protect END_PROTECTED
