`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q8i4iByoSHWkGKMbVnYOeZ5e/ecT2cmRPqpxVZ+wPP7vHvvvziJwRaE6it9Jxk5Y
6oi4fPra6U+Sj3YHmc2Eqe3SVGPdSVqWHK3YSSTDfLN/KlUBjo1ZSfm/29TrCEQ5
3lILKBJku4pvpg7ZceVp3jiSxuZnFacG8hUhn0vkpE9BsQCZEDKUZmo1cckpvbFt
GzsNQib18fzy89z0HZ+Z3suXPtO1yffx+AyJRrmbZvTQqLG4IqgbHI9U9cohVwl8
cPGRS4VoEs67krOkH8JvXQlI9BmCuPus4vpC8GGEfnJpyaPEaoGspWtEhnzTnX/1
F4nnDyg7FTTfEmxygv+MJGhbM+7WWO7Rz3C4PbviTFS35eIxRzba0nW5H7ptvRHx
sy1E/fh4nXwcDlWP/GrewyKh3EeHVVM1zM4wI6wr0A3kTu2ltcpdPfO6fnQd6WtH
Wm30Blpq1sKaH1wdFFzQsuOc4oYiB9txUasDy6qa5S1YRFfmgBkcUIkcfrEP+XvU
sGof+7wb7uQrcszWrNCRRyiMIQt1I5Jrqc/lQ9EMLeoc+WoZksfDJXBfIT2Isgwt
XaD1xMiqmUCAHJVJNA362fbAf3wgMO1oaoLXIcTJ1izZMqKRcS/qe+P4oSpLIwlL
o5APplzQx2PpFiT54wV8MnTZVoue+GGj+i4IzRsbact14VCFwHDKzcrNTWCufYDe
PoP46CnTUnfb97UoyGQgyydxYoP4UwKZYx5ww0XGEu5EB20ai62qoDaKyUonuD1i
J3PskTudQs2QJjZ9NoMvrfk+RRF8QkpltNv6Sp3cP3e7J5uKJ8jI2HchpHZpftuw
EpVhGJSrjgY9p8Zd9bb+FDUnOxvUyJhaJY2+kQ7q0xsZXf6o06dIxR1YSgBX2qH3
ha4fDRhdFSmuUXwYuKywJJk2Uj40JO//6hJJZrzgnuZ/Ha3UF5WBqgD0I5J4ybew
ZJOftwQrJnlBt87xPEZhwmqkzMkv9Cza2NtAgDSmeg68ms3oodIP9A3vpW1jzbPY
nYDzsgmG3YqXgbYXjhdY7QHWkqvTGAbqHs/VGmwk7nWfeMmO3M/2Jfb7UnS6xV32
AtG2s8BfWxHQr+7Slrn5JMDKuw78ik0k6SKuapk4sYXWLSoyaFpQdbz2z0jzGG6z
IrqCJsgI45uCf4scla5dhlM2K3fWFoYhYSkymzhf5SDPQWqd4luid9aj+LMqKdaI
gz3gBmtvi5edBJqnz94J53YEHgIQJtGhad8+XcpXE8fR0V7alf3lEbJeQ7nuEPZU
O6+bm5XYb/nxBomATs3m+Z5hdeIKa2nN4NmxISbCGDILGWCfFxxpbA27SlTMlg/R
G2qRXOvnmImVS1Op8IvEWzJlF1nAnwbELKCV2+J/mJTlxuHwi5d9EtmGWUnnqGJ5
TdKgJK/Xyrh/a3bALG3aybWlePeTRdSKMS8INCSXQL3nKR++3PRbP32ldl5dTVgQ
tV22nhES3WQFuj12EjGaNvHBjCTjZFc2TpjGLlm9Fzs6FgEQ1sIZmyrLmGQFV44x
hj98f3OEW/0KwAjqc2uTRbOPuTTYszNAet6IH9fBl176Qh1jUyvpe1HiZ3WWE9HK
9dYgjaUMngxhpbmsfN490aX4ATX7rbmd3fvZHPXaEyqzmlLF+rWHgea2zHI2Oi+X
d8kbqgY7kM+48THqBPDYEEDu+n4iWVEcX6pmvU7oxHEFdeMTspayHPiAxDDQBoWv
YlrdV+ElFR2ipCFDAvWLV4k9WEJfDPH0W1LRaWqqgF9hYVX9Es6YDDBLtFnI71ly
Lb7bMyPuyaPBTS8NyAmYBLtIEkyuXtSg3+OBFSsHFBRfmSprKXGOOPNc7W36T549
RF4+k7k0L8Bp4hnVPeq3T2ruC5TNorUdV3eaG+pt5U+xFFl7tQZXc+Zj/j70E9rw
SCaHWddwvt+Tz6jafFwdTE3F1RPo1ed8VqeTN/lqq/wNIf+gEB78UAVCgwFcP4aZ
TyjIbJqUHIgEOs9rlkkhApItsKonXod2aqR3C95sVeGHPf2N46z3WSEeFCSQvHFK
7DT1lPjyWTJQJD5MxzE/NsNXXC8AMKdW27ZCPQCLeLnnlLcVf1Yttt2xhgYORCBD
9K8DvaWLVH5OpmrWruSmL6fwuTaJtgYzgv73TBaLN4pRIp3MLa4FHcNdcbgmOdbe
`protect END_PROTECTED
