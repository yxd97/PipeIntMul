`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bzwM9r3+2McjN4xeNlVetPwnlkBT+h9Nv6/HM/wH6IpigvwRg/BrJQGgSG3HUtXf
SM2A3fn4tE83OhrJYehci9WuAUf8ZbxDSyUwa2fhruvg7DSpgg8eubXrpSGUSOGd
nffwAJ/3HsEclVIaqVTZ1hgRbWz1SNqi2UFx2KdA9XTPaCGKmk/Zcxm8s+z8TqUB
7pRvoY7j0blYkiERVQXndnlUdkUuTxirXKlpEp9Ltcz4v583oe63XKCtE6+mOtSv
`protect END_PROTECTED
