`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wcc6f4ks4G3QY3IbN4mmQufCO6pJOEy2Hb9fJ8DQhYmeTwWRKJS6thrc1UemHtjT
7RUpsowlDs3nLaBvHdTJuIt7VYHjUvkWzvX8ipBi3CQ+GRJTjExh4hh85Iq7H2CE
UyTOhNdBbyyvroi7FTmqdsxxfWbv8RnOGrEY3ETU0GrftKFKQjExi/OItS7j3A+T
RDWkb65uH/u+Xh/DU6cei4wS081SrHGwUCj7fxlPBWjrIXXQ/JCltcd9u3WJBEVL
dkVyMFs5vzfDqg9SAjxMiu8jBuSs12ZcO5LGLHZTw0MdJB1ZuqS+E2Ro+t+p/Lmf
zUNNKh6lJucFrDWZQg1L08vDTgT7kJ7ncDP7tIJuXwZtRq91Dsq9mQ7E6lq2ONPX
ISmX6XBHtapdOH2ewQC+ggm+J17BaCodQyCaqmlhCGZhstIxKykigt3idyIhPGhi
8nZ6MO5OlmnMAt5Fsl9siASwuOQhpX1US8ywYV+AFNbCPcXT78/BxCvYabuTyVbT
`protect END_PROTECTED
