`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q2NegPYaK2zY/jtZYoY8mbyG20HLuJhepLRw8bWKPGIh2h04rAImFIW7KSr9KCXn
ixTulaov0BhJrEVBUIwnKwnJiATRX2IDK1xPmcaII4WKRaMa5t5ztFobXiSTGQyx
Su0DwVVDn2tSYB4LQyWwP3ziv4VRMqkONlju3JbccpLZgLftHhXAF52iw3hGzuCB
sSgVtl0+CozPMfCPDEBy+V1RVoCStxpEZXOUEGPOXbM88p09y90nNb9b4Xykj2SQ
cas9pIu8yhQIR9eWCc7g0oDQVmQ8hoeRA13a2hsm8zXqCVgsKx2f4xPhXiS+Ch+g
`protect END_PROTECTED
