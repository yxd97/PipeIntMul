`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rGWTKYOduaAgJLjJCM9K46GPNbvK/AdoydBEBwNw9C2iR7wAhavDV7n/PSGdssNa
fEYZNpt5ev7RXtiSgD+ljjCyNSl+JyPfykihF4HDRPnYEBKkRCEhjrJ5j9nnk7Sp
I1dS5GtAMTufDcZ8JsOi9+6Y/HTCgkTVhhazDQvS8vUOqglP8wGYw7dFTW2f+paF
b+44pMTZHJTGP20vZV0OaOARAXjBv1jRwHaNMIjRS7KlINQc7SafWwejIw17/V3m
PS7ZE2ZEy2slbuO3x4l0EpootyvdQOrLE9v6ctIGVOBTYFLwX6nY5isAbrsv00wc
voSZOzFc4kJg9jA9gXmGn3Hjyq50a4fh8lMS5MnZ4SdK2vUBRq/t64NF5FBVX2RX
xPDQyb7rldpbDvChP9ONjFK8jWtoSfzc/h8vTuUXUw+mQT6q3DGWnSVrk7qDDeHK
g+CqQix2vj5sfVOWN5wN4kRRpMQH3PtbHOh2hSf7mb+/5z5WHeD8tjoi8KJ9/3oO
ckvzyqZ97GJ54fcGmHYvYB90tNYzBHU7SWvdxR8S8AlZoMKeDIQgHC9sOn7IeRQ0
ov0Vk7te9NC3XBP8G+uJkPAR7jM7BkOlwS5i5KhI2GnnY39lLu9S9hm+R4NvOmFA
hGjVOR2WGinXy09kD1Pi8B6PheG2rAU1mvymTT116utkFQiyBgut97lyo2VtgiAx
il7wLUN838RLgxzeNFTe2V9LWh0aoGVcqZg3dw6RPQwIA3tEp6V9t1lc/Z+Wh8cm
d46Lrl+MIF8fo+NhftnZTycCG8surh9fxM5P/9vyhJc7cOeeYidtq72sa04uRNoa
5/Fcg7i+VJasIuNXMqT93vnuGTQ8LRbC+APT41yg8idz0KEu/nrto4iDmHCC9CNs
JDj9cnT6JxWM9PwfliuCk3EqgOdTchVvW7s/PkPTvTH3O5v8HhQ+qJSqzsMIKzw0
pVeJWKcl5b4dSzrPN07r0dlXjdwq5RFoCyientT9mMF4YgKeZ+2S5s8lXLALNqZv
3aJXgZ5RPGNRN1ywNdzJs7ePfZh7FgVAZxXiuh59KOPYoDg/Fbj9N1UGi+uTHjWY
`protect END_PROTECTED
