`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TGICBFzPpnZI3Du/AYZ2MsnPQX+5DC3TA+zlSUiiLqmAqEHujwIIontWMi5wtq/z
iSJNIRmYq0V9AQORdY9jg8i/c2aNLl1AIydbPl1CnBGciTLQdfZIViDEEcPIiSpu
sVp+Uxp5z7/Xfsao9wkeioeLUnn674a1KDyWA5gTAnedZsPqS1GeG29hLIdocMZx
cKVyxIbI4bJkvCSfp8kUkb3fgFdP20+fw9Pg0NjkJDiwcMmaPbiOEoYUIiiqdEvO
Nwq86C2YDeAs0pkBKufET502TQPz9dewDY4YpluOcRkCv+WDmCddyOno0xTpno8Z
scmNstB7Lkp05VSxgBmYMcExVER8OtKTiXkTZJ8nMF7ED36wiBDGG8qqLCghbKNH
GnBJQLsdM6t7hA5O4PJUeGmZmqcve8lAhCqTu5EthXlbYOXcTtJWiE+EvA8lD8zY
ceHYD1CaMWz+fCk5EJT3cs62UXk7PlmqS9YoUnTGzTIL3Z/HFlNsGqXm/jVPGU4i
LcFVN6C85gvDApy48fuRquHAdoT4VcWypq5pWBu6OOyyZjfsDizenQJCsOUn3rNq
cBG8LwJfmg7TpPzHiip4HknJhaxJ2CEvp4mLA4orScNWF1u39ZxEFiFbFVzCMLrG
O03Z0InVVG0ZhNUhy/DYMfAqrXZXhnv5TqQwsb52bLjbXZrpoFrc7HuyHH/zqkVn
OTSY3Ke/te9mZCqaffQOCddnLqiPigtg9qI/v/pQl9rT4XHKa5dKx+tNJ2awHqJX
Tz7GpHHa81n6D9Su5SOH+MnjQlLTOiIiDYSJDLXALXcT9egbBK9sgy4sSfzzU6WJ
ibNBl4iAKFCrY2VptJd95cPlFB5GdMQWAkWMBnItxbn2Ufbivldlo08/4ya/nog9
R8aCVoz4gqgIDacZccWk5A9iVarU8Sx1O9tAxyOiYYJTn49rzgjLGjvKH/XRNw5y
9GfaoZ6ymSEDl37BZDFjfehHqPMtN7u/AEG3lcqUGkV0tGJRc9mLzAXJ2InYc36X
W44dzD6IztAEbF2Wuyk0IifGHpy6fgMZaAfv4N4plQTzs4S4xGGnUCvv+dftGHSQ
sXnSZny2s1u7yqp/y4U/CiFOijc8A+KHSyX08JgeNLYKi51QwkPEl6/7BVoWiiLu
l5pwC/ggZvnJllWO4Vz5Wjz6Nil2E17gKamV6V+YW+FjAU7n3IvNgWhC80BAJUdO
TedGngky9jYqNCt7zorJBmm9d3Jkg7mz00mfjgPwKa1bhxX/JFUbqJkRpebjv2v/
x9XsOLFHGpqVsxqr256t1wqpyJp/etAVF2/fZ7hvGcqjT/2YGCDLQ/tJkvdMgudh
nmTzBHxELGjKF7g5yBDTgoZX9xR+ETRkjEP2JrjXbbMteeOZ96vCBRR08lvrEZyE
59qUzlORQKaO8XPcCHHiXsAsxYqGKM6psCOaL9kT4SFzC4yK/gIMee1xhvk2pXWv
12ogFpHtHp771QhzTKL9DFOgsxXKZDE3EbWpgvJWiof/2ECwatVSiFuivZcK/ZnU
q8XJI7/Re0PwmM2gfwKWU0tVPOLaLGt/7OijtUvANbcXY5KfHqeygoIpMSHbiZp6
l07K0ArH8qff+8w1cKcti7q9c/clwSQvBUhB6UzGHbHL780SHRRkxVuf36Eco/hg
I3N76H5U+d2q4/qT/S5rxXzBctDAe5vgGhUh7GlvQTOJCtT4vhGFNwgc/ELQp/Ue
mRR6omVgsxPQwpIBy7xkHUGwB/RzgVEawb+jNOUM73SMzGmAfj2u/gf+yKFsUWjO
38C09OXT9A2Kzn+5Np3Lkh65x8VF6Ql+bSVUrGRfULku6/w4DajJxqwqLDovDZGU
2yGGNbXcn29MA/z+pg9O0u05pX2xAsmBUH80COg+EC6rHcN4CldE5t8klvNRiE6H
6qugoffwsDY0t9pkF2yi1agBWX+aoHTmr8UNXKQLb45ZDQYSrzMxeN8pmJCG72Lb
ZHbGfGeJt4+oPBs4mQ7anPCpaLYYWW6NOL4AJ1amaAMgNLM9lBnEaLZEK1b2eHl5
Nxj/nd520glzVZplCMV8NRoTCpwJ38UTIPGTrxALl/G40o8ZfATZ8qWmZjWOZjV/
jz6zb1lH8LTnhFseQDr/zyJCXQHeguS6Ttw0/C7uwK6aqR/v734kMLaiBaJKvERY
Og7MqYHDxhyLFYMOjNLQ6y+4mUubJN/ZP3nMxyaVq/ZXRSvp8jkekPZAhcs4yiGA
g4tXz8cTZHjdn5zzcdra1U3XhwGEMvjFRy6t1Fonb9bxJU1qEMXrVw2FzNPF2xg3
iQcekxwQ574TmCy3vPUwVe81tgRF2u8kRaGwkOCw1BxQeOPDBw7/wt9JS+E1GjAi
NjEvL/3L9nUP7Gj0V/ItjAlgEYGYJEfQE+TWNyQgX8raXeDl4EDdhGh3lEPfoN5E
bOfBe6y6FOxcycG/GPoqsTfMIrLHkkeLVkrCqn8vmuxPE/+iwuBogVlcDZ6Nqb6U
VFpXEiptZDuxtrejFbBUanof47TugmydFwucdIrw1Op1yyzhceA5lJ6TVqqXJUst
ELcbxYrcMZ9+OPZsLQE987vf7nBUMg7lw5GDZmqWxOOGZ5lLR9C1GpkTRDyPManc
q/Xu6aSXQPLsnrop5SYj3Y71MQ/J4bdbwytSZ7ScLaWOxAwVV3VjjpGWG90atWsC
DK5nINjZYmQo8mNQH/KNnNm8t49aAjvQlJBVsMJU6iK2FGSKDPqAtUYzKlMucsoo
N+CBus8H5aQVb3AzHScdKABFzGsgbduGGYpeWKs6FsMljh/rziorBuy7Iq7NT7CO
AGF6xP/YA0Enze+l0C4h35Rix4FWDijEBmBDiQo+TIjNWpwcS5kL9va9BT4etUWo
tjs7YB6EfuqFU+dLt6vV7MqJ/ULDv0hQDC0xwRZwCxsftOVtV5aNGAx9GO5B3OGI
MqTmATishrOfX7mzSYCO5etTJJWBJ93HVhbHGiTogpfxFq3aMYIo4OnkvJ3mpiZD
FzkXcqfn7+OBwrGCIPjTFuk3Op7cAs6DJgD2ZhbAoTLakpg0YieBrghXyyJ53gSu
WWIY+jSrPxLLCZmg1xSdJLZP5XHc8H8F4e6ag7l24ypGa4alvDvjxmTTj4k/d3S/
2BnWjjT4mqxE2+Yj67xCsYL4vg9a9Gz/SOajYxI51ywxmzrbzhbtdYLiBXOERM47
JdeE/+uDF2NdA/u5/IxPQyz4nHHWYMNuYdZ3R8M1IN1qt9lh+dhAJtBzR3V0AtF3
q8mHDK3t4p6O79TjfzH3SHzwk83xuY6Lq4OAUoSMKMavZhRBLDzR1Gh96Y9pCCMQ
WBUZDYbaJkGnspc8NcFDuVTXDKqikad3fZypD8PGxb326+a9MB4by+36g1imUmw9
60vkMqAeC7WTTyNbuxs7dLqSfVdRn9dJkJYIudwTLVeSb5xXQ8tiwOSHA8enOIQL
QNIV+JW5Iz5y71ilJ0j2oiyRe/6Cer7XDqkjKxTxVXaic78OK+K1tobYnIfhMcJK
DhEVMcilaydDuwzUHIhBtI8Srf8v3ebbnHJJZHQEWJjS6zcqOdJDW6APbC2NbGBj
S/SyxVBtpuNKb7O+9y3ltZzMmSwt6UOyaxiw+UgjQobOv+NCz/souOLWZXoKeWfR
7wMyoL1hdebWIqhspxxqubHcwWe3YuQ4YTYyg3PiK5PQH/0yiiuFZS6WoDOY6JEM
CRe5S8m2TIT5DkUQKErAapWxpLgxsNSrDXL/pienmkllm+mIlXpCG8IXVy4arJsu
x292QQvDer1mldHbe/ZSz6F/XUDpXcdUtz2UR8CRxBse5SCymHhVE5IvEsgADQNh
7hlIA+xBwR0OXIYyV9BvcQRhBk7GK47hx9xsPzTAAlbt7te+HIsIx1Jqb99nKTeF
AjOSX6aD0QkgQShfWjD69Vet1K8/tx57pA6r2UML20lqyPjjo9VMKKOpEnJZs5El
q00qjCPGtR08rjpiSnT8Ut3A7mi7fpxvnzrkPi4S1AS1Z75N8s4Aakz0hNQgC8Dn
XLdOL4LB9vHd5e8VHGlw4yVn8t5r2TF23qzXE5FnHwNX/Z+6N+V1LIgaGYdBt4dT
6WyDPOBJU/tkoti0Fc7O/1YExRfK3DpO7SOlZ4zFvt6uavF8EUxSiC94wKLZoNvS
wSnqytShCgSxD+EaqWPHnr7g4tSCh6vqM7ZWLhQc6QKvXZuooxfKG+Rbd5TcLHHZ
csbgcseJ6ZzQtgdi57Y8Cjs6JcefmTdn90CUIpWDvE/Fs3slt5drqVu1JWeBQ4w/
jP+GL/e2txLBo7yo9OQs3UtsifI0E6c/eEhhLadwnqS4lwsXfPbpNLZqFkvp0IBI
zhBLI0XiURAF7qs3sHG0eHidQhxPPks+tc60KhrFvEAYuxIuXVE5hMow6zmkhEWG
pMe85zIugbshHsAsWhd2fvVGcBjCulH2tqdx55SPqhtTsEzy2G9XZOGuxN7+JCPK
1oXRiYsy62dErR6UZQsj56b0qArYAov48rJJoQAV4wKZFWxmagjgcBEAYOoU+gej
q0IrMYatzVKjYQ9+9bRCOFSRyApmRGIeEPtJSJdqPQ7FaLPrXUWIcjaTerE9valz
dZNup9hDvBhG/P+EmnuWCiQo2tuVJ04CXCfNKzsnjGixuGrnoNUYJZ5OcLoezczG
QLHmEWdHIqcfgdOBDQsoLyO20hBqmhsYDw3zAEPzRVFbYSBmnimrvYkWuZ8th7t0
QnU0eIPhpO2qulkAtPjPEALeblfj3AOsYwwBKNSF3gNssPBvecrcTcTtM1p9Ap/m
ID33h+nOH5THxhjcE/OYQO9J706K1qaRqKUVb1A4lb5txYF7RJl+U4I+PIowJYg4
OJgQR8MUwOhRnLGMnZeoHOO+RzDL5GUNhbKu1QnaaGpwwZvefLcVlz8Z4iHly654
r8xAWrXStCjQsiFSIjlYdTWXFtiRspvE7dLUuPhgc0V+qNsPN5j7LhW/rM8aP5Ct
z9kHviiaNYKaVz4sC1IdI9ICIXS0ADODh/hOiJS6Y3CGmJ9q7qAEGnAjO/qNZl3c
13PFxD22tQ+gSqOL2uK8k4ge+/Nk0ZaEbeUbHo/7WUh7LAJckzldOOJiq9BOZNXd
EwLxNtNJaOllQ2dkUr5Akj0IZ8u8goB35B7+BzFp4FM59krqGU3XQpoB0Ww9ppJJ
OLkVZpBf5VXnJETsl11JXiT/7LMWcSozR3kPZ1z432MFCj258BJE6AjMSqREF5CC
g3np398lajXtF1BmksmEYDw9TKtdJ3ruoEsn0thEFRvldrq9Rdj26vPS0AbBFPeh
UoTVsyVkRP6XAIK8j9fsWoHi8P9XVks+sgKv49vbjhfo3qMu2gmJuO5/ajYDFqN3
B/P27r0sWuYfGSfMNEFUCQC8Vd3DVOH/JN0A4ZiVWdFk3Xrmnesqk0SV7H1enJCN
bdgFQEl8iKOzlqa2w00N7KMSN0WjD0Mk27n5FpQneQk+aF4cuwJUojDs6u9eFYy9
YtVigT+WHZZFo6uBY8upZLPRy9ylZx+eC9GA63XMaNoCHNz/MdBbBd7aooVZw1Oq
0oSu2LunFOZW9QTjUDSph6aYeNNi3AnKJVe9ZXOU4NcNp078K8aL3wxBZ0g4sadQ
79upSqWPH77910SUaREkhu/pkgZWP9rmlw4tQ7fRvZQARQpTj1IslaWJn27CWcJ5
Wv7C7rgW4BcTtFvuuJBHyuZO9Og6IMn6nBeXNNjrzPZveWheHIE/JU1wKdh3H1TQ
V2L7HObZ5I2g7pf2o3jP6FOGnhkH83McilFdSVr6eOos6oZtksSn3eF8uRruiOG4
aRuioXhPH/e50A683WHQfb8juwlMtiLBWBPxpVp+pml98ALC0DxJ5EIRccSD+vyM
1AzGJ+btt00FE1hW4tQV95rgbtCEIbKwc0NRYncs/CoG7K4L5V/iPZ5WIW4i9k/I
5on+OMNWphMzc6HR1APWDRIy+XquYQFKKmUAC7CC3r/0zzLoDL3im4mSZQWH0MHI
34nuQr8EQ240dTFGzyRfXis6zZNNI0RUfkL5hy21xHJhNIIqA7qUEZCCkQg4n9kd
3lAheQ1E9sRY6zyd/vpIjGlcpjjFYXFnngtMb1ROhy4o5EJRvY3xBQARrvjM19h3
q/M+0h3DQ+Nsn4jdsUY7PMo4gCcuDwer85YtY484iVmkFR0a2VZUk5MldVQoGUFB
omKezRKjJE3kkDyom1uteLTAK0OAtJ64oHppfJ+faO9e27JV4CBSmAOViaUdT42x
6u0i6Sv8RauC3vPQa1FNPAkoEjeUOIUY7xEQYy7ztdtR4lYG1qHMUsfAuOI2nWEO
kT1G0+Qboh+MptuPzEuoIR2eLMFYs2MSBxFFeTHeReIdleeOXDE9B2LjWGc6c2Dm
PyXJNlhq3iCkxso3tzdgNNp+o9FJQNBWG5Lf1l9RpavRL9VL2Q/WjB9ZWnCd868D
73iqi8jx3/fyTVPLQ2KqH489zRvFU/dTNr1Cd/PGTXTjUve8o7lkkGKR9YpYK28d
W4T79RBrpDpgAcW4Yv7aFCfXuOmxuW8eNEIwt6pVF28aYGlz50Qo+HiKjZiNKPDr
gAQfbdxTAsLDD+pY4bz1clW/LhCj0CsNmQ3KlWFKiNE=
`protect END_PROTECTED
