`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TIFBuhNdfM9/ITKtLFsJrQ3nj6mIypYzItgIbpRF45GFoYKSYqzXhLnMInybyjDp
nas2/+MmgjOKwlei5AZWBdWZeb5IJJCQw42+E7XIZJ+TQq0G/YWmX5IZUoqs5ZG0
LDEIokV7Dq+w5gGtLFdlxWAx92minqholv4OM+5K+kWoc89d4Wx6f2qYrVvSMh/b
LO3+11Qfntw2z3p/erDKNi+vCfWb0nMwOjwCJVDuwZCRWhnjbvMlewxiCnZ2irta
RN/T7SxclkklNIArtmfhO7hGRIWHFGQQQt/7p9t7xJ4WrsUUgq2wQm3n5CmPVYLF
C794UOs6IudsB7cFYGYELe1awZpTJkvKQxFFY5HD0T++40aY09bipmWGKVLl8wkO
NUbHCRma14VIQmmYO7oVGoN0/Nr1OV8HEc8YLFpEeyZmMkeIqT9qw72o0NIQpRNg
I/V6pgk5JaH98+PaZELzm7ohdIiUmz/+RxZZQI7z8qQYz1AU6DE7PAjTULk1M7zW
7k1/BYp/6iYHTvHF+uzLzJL+1pmb6Ekxc6rYcyZbqa61MTqF9YdyUUU+a8gzu+yF
Jo8AeftFA050uyXEHQzMn0B1shCgQE5oJJKUa5piAIz68SLb1wUHTE6ze1av3m20
AbpZylawQrDYZ8xCqeF7GHaS0LinQEN1MTw/yEc24wfmn+kQegxjHPtqJgVKaDGg
+D3gLvZ1j2a7tvx6ZRH5i69Swp9iNKB4NNn3ehmFZFwPSwlmkNIR409tBlkThywg
Wfc2bIwJ6UspsOCxt7xYeJo3lSTkPCCEnT2IwND+qmQzm0ouyWEkYF1wVAu7D/W9
oV0q0TDuGGqNA48AXte/LspgDrgyB5SHpry0uWfamFXj6Qmj4J2WcIJ6T6PEZifw
gGfVU4nyxEpm+KXV2HFwBPpwKECc82HmpXDHmW4oRgYBBl3IEWCQcZlCHOMv8XeX
5mi2xWwETx5OMnX4ZW8kB7o1qyiAGKt4QCxQWXLNmq+ColrRAsAnn7FIDahEjBmv
mn2eds5W0W4Dm3agPZgV3I0AoSSZLkYYWs1vSBuYjxeB/mv34hPHNhG2hrC7sm9m
YzwYdaikxPFmZTlZ8m30K02x34MExrbKPfKNcHAMpT47u+WsBrhFjOZz+o+PDRYL
1on7wxTTsTGZAtIn+1dwXkCP8LABLNEtGbo7X1r8eU8SLSNYG6pCdQaytihe2+N6
iDeoU51o74AvBe+IfGN3sx2ht0X4dIIcE3uRbMc8sLLFSEv2ScrqNZd6kxqVOVEF
F46TITQIdtoloGhdT6sEYNj6PevqkIstPjx5axcjU9+HgRRzQ3sd0o043bXDgAz/
4U8i/BsAuUwpn4FRPEFIuVxK8gfNcylEPIxKDZdY3nUKTs0FFTM5lzQj1Bl7UpZK
hTv6irWIafQnpasCFcA3uGimuE9HEsRgPnYmg5Ep8/osUzLVsu0k2S4T/HPihKi+
TebonbJ6FnEbIof6Jx2zgtRk6+qZD7mfOcyeSb6SdQ1pdtkQjtuTZKIMALvFGu3e
uV6gL7vC4HUloTlJXBdwHZkKmgysUoYbw/Pgas9BXZhMqyaAsA+o/JT+EaNT7TW+
ZFagrs9mCvd0r2g9QdUgXQayZ1kK2kzYjoNhQCtaRu+qUMo893vOIKWgO1Gy4XKV
OdMCg/IO2agFESj1e8bB9BYtEfbi/1Btgg9SKU9TpIW6utgx9XaV89iDlebnA5Dt
X2y5gZix5oZdyZcCyFttfd8ASSJXA1N2PetXmUKMaUhutn70DPWTloKRHqa8ep6b
Dbe3HqFNag44pRa8no2X4i26fqZve17N7yrdSzm9tq7DXp17kUZQyKKtXscfeUFA
zEVjRNITMLnOpoM8quOh6lKyEsTz3SOIFlXtyWWTKAml3laJjTKpQI1OCrA6NCkW
hwH6G+SXi6ATpl3HjOFLf+yLQfRKC7pH8r00+BN59bIiny2WFMnjvfAzhZclYcdT
xzzoCmuVtLIEpVBzl7FJ4m0mw7t6t12B5Pc681rgRuEcy/YrjhdAQrzzbd3QK76n
A9K6RsXKU9xLwYgqUeJz15kwDq7X4EBg/GPtfy8uRFBFyXWOIw91jTBUeXBK0rHC
QW737mc+poyspWNxLH3tudsxr5EHx17B3EWKjGy/RNNV8dTQsreQw+0x7mbusZHF
r59k4dUB1cCz7KD7YQ0ICwz6JTDql8Ua9qbG3ntXzrIFrsUAOUeSwN/Cb5xICsAH
FffSe9t9rq0/pUwWIQ1HwBhpXo1aCjNgeJIsjgXcenrvDfkP7/qAC9vr5Ep4AZHt
E9qEK5N5ksl0SE2lNdaP+3tuEAtaWh0xjF8IqCg4ahLlw1OIDGSKsZVcqW8TxThG
e1S+3ONqEwh0URr+7NRXqlO8zlFywI2Np2ptQ2FL44q9ZxHQTYz7DQTwKQTxMSCv
jYIwgMHhipOGrBGpfOonfgj/Ld2lWRKUPYpXPTf6F3AUcbH3VymSmQw2Vafx3fCI
8jOxPpe+jiF/vlEmTM92dC0+tPR3B8eqqXVosExDN2Aya5zGHKtaOrzJMI5Tk40b
McjOu6jGNMrLssbTR+t5YhZcbsObyaXrojiMssUvwj6jbI9WjF8G6yyMHWP0k/Vk
zZ5P3I2m631TWTw6G2p18R9U3AYWfJVkD/eJynFtbS/zpVVbtL0yMqjNKq7VK+Xq
03JK/qjRV55d6sdtP2WRKVEsYr0zQICEL0ZhBgPogeCIcyUu7zSIUzS7RvQJqcGQ
ofpIzHGq0F+ZWW1HbVr6twT8F23dSxznNCwg87tFgBr6u0+yQGDaPlZTOEVROU5p
MK5CJ0pNEuPakxvbnLFhjGNmCBwGDprUqqrwrhCaWrFEMECvHasqTUmi0fjL+Tsb
Voc6WhnPmC/+Ay+d392bstrq8T6s7czW1xKt6iwrVNlMG0ZejxdGOAhA+kF7DKNT
jEIEVElc1LKWUb91AVUl0KyuNDXf2iwTRhKvEdGTMlCBM8KvwXvwcQ9cnoiTGVCL
M6SPYZGomTg6BHJGizQJGdSXXV+l75sufOjDaI9l22k7b5BBvGO6AKYbNPzSqGuX
n/1gwm9oV1WKtJ/25GWNHntY9xL0HWLqS9FTJOOJr6OKlI8D4diSOqVfvXPXCQsE
8Ar1KfyDhKq3LVJMCs01d2jNOuOAnJ6iIDhXGpNRKVV3402oDJCL09VtVzPZZWUG
YH7sRa/OmyoVe9fUlrUZQyKYDUFjivOUxTIEv8zESytHmAoUTisAmbTeW8vVTQ+H
cQQlYKCFxnhmSDlzRcQEa1GCdXSWREgkLqP9WEeu/nBsQqwwhX9EvwOKCAm8UwMA
lZgzhUWuY3RGAEEOa966e0mMmxjT1ByZwXBY8NOnLHjx+zX9dsLB0KREGldQgw3n
0CIF6RgJO6ITJHTdNp5Dgt16EsJFUBekutpOdpaHeZdxUQFCBGvfiOhpn+c35fIW
/uQIk9/f+SxJSHNSiaLtzFIuldcVdS5knUEfswIhgRrk3CB5aJLSqcexhU1FX7uo
2EYht9Y0zvIx/ctQxqtgHSHkMLU9xOw7xPOx/efTyJBUXY9HscJt9/Q1sGjHQrMz
v6Uq3pPp9/RhCXvSNUplXNDWT7a4h4dpvM4F7Nk52HVMX1Vhnb2qmDXBaI10rJrz
wJuYuiOJZNsESIPKt9DEg+b5BpDuedH1dnd8VKVHeKHXytGbH7u8io/4H4BjBvgx
NRiekOODvYLW39bvD0AvdIQe806VdiMC6j63D79Fh7hjESlW5MzPi30t6gDu6Ek/
3IZLhMc8L8CIXuSP4jsum+1d1YHO364JLrH7iXfJSyXZVblAIz4dYp1YhCJRvyoe
zX4HlzZz3KqXiRC+k5zwcpW3DT4R8F+q1k/frGfpgsv0JMu9KMxqtY7r62aRLFqK
gIvQC62Snhjt/cFP5kCnT0W0JKgywyAb6U4QP1boE8g8WlfpEdhbF/ZHVkfnyD6j
d7W8BAah9fXZ+y3YMPMvMGEMEND2V+CIRiuGRGkeituTQPLUEKfkrY45Obq9c9eI
utYDdLeRLFWeBXVd+sLPmAvxpeoTSD9+fp5UqKEvWouKMLQX0oOlEkxRt4PfO7lv
9njI2iHZV6f/M46YVdynbG+n3IJtzkzI3omGOmjhRJ4zSI+PoSVQzIsW0A9dCgWE
kSx5wqEoIn/0nPW248K6u+k7PAGJw78Oc2XVKCD4Yxj2omdvU3hnQQ33GjIqq9Qp
HO7uLcI7SfwoEEML4GRBAdLtDwgfMU9+HL25bVSQZrrmNfJPOwx6GcZtMALMLV9J
cswltkUc1vGIoHfjqkv2Z2vMYA5bReYh1V4PXc1Jf+tpduB6cR3gidxIs8YNXJMR
g2Il1DvTK6kgqGbk3UHdUksHsgaHFwbIPiobtoIduziOP1378SNjZvPcZwIEnjYD
D24n8u5POZrtG1hBrt9pN/ceSC6GOccyD+9oiAgOAGlOWWDQXnICVY4CeNjOEq8u
HQ36iojxve84qHwjpqCRzzO5ErvuXiWzwBTmfUseKg7qElRXeEVJtYehh79QX1y0
7RK0ocCU/wE8z6Ling4y56wKkc2F6sT7lsatdozfHDE1sgkxdJVTE0eHz0akQYqJ
+Zy/J/LUXfDTL7hzAoiyDsInzw0rarWIv5XBEEhSJlg5g5WP2zHfQzCTjECXH328
asdkI6iHzvI+Q837BJGQUi6yMgmVrGEcCjXyXj21SY8O1fawVwakCv/+r0zeh+BT
lVdDl5xwkx/gdJXk/Q6WYGArjpRrtTMYZuhh++Jv9pooi59DiKO9oyOQC09G7Q9B
y+XixWl0qj8ILGMocQogT7QYV8bWhkYPR8JTAyKlrRahHKSOY62C9SL6d54RyDCd
jkLCMsUkGHHluodmkyvEDIfaSL1+G69fx/o278JsIWER7cG7cYniYQG33qAlHUfq
SBps8ZUqz9wIQosWIpyjd0oR8Dc/OYyRybZHTiDtPSIlnIG7UrM/6axW4uFGBq0/
7RBenANVWtBLlZ3jrPIgLrRqzYCDN4E7ForY47wcLXXL0JI/pOqAx5l/F+xKTY6I
8A0DohTUuy9cC3K5G7EH5LIC0y/eRlOz0rR97rqLcylFN2JxCqGwPj3WgViHqoJc
nkmCO8g9Ejr0JJf7YTzkhGQVR+l88nxtGohscogXSbvoa6/akOJPwIBgyPLIIn6I
96LATF9y1DGlE9yA5vXcGBWM6lFz9LowpfP1tZjJb2lrdAfYjOd/WV+Zm/1DCt7Q
bb/i3/Sjn9vrUWeQhxwHD7Q4szW3AGI+MnLTkwhXlCf6UEx1HZlF895P0jJq26lA
PaCFmlbd/XePwZX7QUr5qP71TOc7Tg57pScgChlD/vNKL0Po/5/T/dK8gU30m71l
kByODjF+MFkN/6T3cazfnOGv3ABPFs4tzu4w2gmKPbYLShQ8v9EtjQ+1imTOEQPY
2+RRcglZuZGU7qqbb2IvlcLvQdsS1R0auxX0EQATTBBgBZNEz2VqNNwM2E0kuVtr
l0K+FfFkLpqgmsbHX1pchc2ep2c6c5THe8n4Ac4enrXmXww3BBDy02CLbZNu3XEW
uE7lrMqaBVx8aGkg3dS1gDJ5TnrofZTVVtH/Rr1zeB9WE8zCoyq8ajsfFTLX++vs
xgR7m0059N2wIclphh94ogyEuUE/h42fDRrQgHoxcdVn/HGWlJMt8QAOTsSFPoGO
2tQkxXLDwDJ5+iSYLGbwNSdSqTwLEJ9+cOozi25qQ3VzQgdTx6uWnnJT5AayNiJ6
Fn5+nguyci39BEqqQg0rrKKVcxlkeDxf41b+lpyrSmL96LH8bpORQ8KmS/5KXsgX
PkogfGKhS0AXtHrgsCxVLFRR3+19sGvWrC7aLdC90oJRK7FSphtQSpIAU95yo7UP
rklnWjYcKnEA8LRwiyDicQeo1ueQlWx2zfpGhjR9S4lTeUfuQZd84HWn4rqL4dQc
nalgRwyTHicczT88iymppiHAgekk1YZ/+8CTOmHFHmIHSflcHE/HuOTNTklN2G5s
KIttowNxrg9jhO9l8qKSQMo4RC65IEZx9QwxTTlOwlUc9l5VVOj6NNICYa4UHXpx
bYmSMMNXGkRmiZkpT/5gJo+lWC7f2gJUmr1YbNwbN3QIEMmZwNcKINfaSVgmY787
j6YZypAhuIsVYGqQndxf8Kbyp5rCL9k91D4Xid3noVjDmmuGRYvJ8Ccq5ZBuQrtQ
tKoLRw0174YsI1NE2sNYYbj/Cf54NfK23mTFz/h+o4uEU2CY08oyAaYnhAPTmgcX
mqTVdRa2HI+ZbY+WHVO47x7JCSTIbFUXanTGE2SleN8glP32SBg9jVdkhQLZMrlt
BjXwCi8ABKKgIKW010FxWqjmF8nJ1Duhb9pVm7iC7wswzatAgsxwo0t5T222xqgj
xDgSm6XKofy9XqN1ulmLRC5HdJ65uEorR5AF32tIHNFRH01UHmqA4WTo6W+shyY7
3mxS6w5PEFt0FEQP2B0zNbUGgtn9TwAqGMQFduLloBkGcR5lgQ8uz1eVCRU+Ia/6
6HX8Fk+0tPzYSw2qowVSxWlirAYTcYOEhomtxVoKjrDdVCkf6wA0wDnjIYJEH9Fh
chxkFz33awtuNvItFSR8ZWoPj/YQrObSAbJfdpbicvrS/lNqmPZMQn2uhfHegCjr
V/lj1PPd4lmd2g0p55ptVs4qzKfdF/IFWEVnkiKDOi//lE07OKbHt+MeDLbQ+dWK
4qJ1sjVJIfIS4suyANN+irtgRIKj37jkS9lllp1v8MnRZ4dZJKWBofQuF90khkqr
bYcnnVnF7YFE611Y3baZxIJ2Yu7vgK1Y62NyWydFFowgKZ9D+vLDrAR6XHF2wh7t
kn3A9pXmC2nOFkAKgLZjNZc0g2uS4FR/7te9E/I8G9D5WJ7SAMJeX0+9yuXCY/0V
vlM+/3Hw6GhJH7RJWwogPV5lJCI8/iTJ6B4I9kAQV/91RmyN2Eqpt9XD0al8jx3Z
sHDKl9p/Cw+vvbrggyY1tWB2UcAFk6uwwUCeJKwbMNC32skxi1OWkzYb/w5QVw/Q
VPkSZEiU7EFOumdUhJM66S4tuQSJgaKH6jdFAjaTs1qjyWkxuoYquVWC/AssRLdg
jJ6K36TfYdtE/U7jiqAMwihVWFi3Md6VVbq8G56yejqlPx8ICX2L1lN0s/UMqr5t
4pwqq2kjB+jEzSqAuGS+n/QL5XkX7fsXkJa+H0SdYRGYtqB/yxdX5Eecsa5AW9a/
4BwZdRHdvZ7mSW1tHjlWCYFXU0zeG2JDhTZd5uX2bR7RIQEJKB0ziH+yztISKf1S
wfyiy0PGAb41t2rPHSlqwbS+Zt5K8P3rjbDUMrQ1Ujm2WFDIixueADEPl10Ppq6n
NepaSR3HK9Crb63sUSHfASmM43ZU3rDhaxZcETO+NWbiL5/VpHFG9JugoWthqMhZ
3sr4SBs5aQF5yNW18xRXwO/VA6S5FbYd9WTThV9+8aOIUI8dxf0Km4CQLlKZp67y
HsblQX/bsL0FMRYVPvLdx9zRrKz92OPpjM7a9h6nuDIW3kW3eWmjPvgwC60gHK57
efPvqXW+xFX3fQjrlaB2M8Atc2EwoT7jDfK+3YyK79W2cMiT9IAmmbeGSXtLqjhe
NXoUhqZhmtp+pP3dwQbJvOKxv1uHXclQyc5A0Clk25e7A4yhc4zOkCOyiaLStZ9b
jRWEc5c1pyD76ekoS4RrMXzrPhcLi0prNqAaA1HJ8cfEJp4AwEeqU3dZg0JCWWqN
LRnjhymXpR1VMcEiLnHFO9AClXGUDT+ZDV/dRgh6Ro0QtdUPO96BkIn5xjUoQmfE
iNhcDMtTALpewWTjhlXgOqqfI6SlXZp0aGuOouz0KNEhPHE1o8Z8SQBwN4N83C38
ch8qvgnQQ9uhUEaatQq7LFIwikilIWSnPxVKM1cRbOEy4mwHhiVq3wjktYXfozRZ
zlP5RoMGDunXxAbcjm0nBPratet0XLkMZpnEDIdS8k46uJ3HCCTSCiKIFsKBa1h6
9el9X1fnotAaoWOcCKuEt8f8qaUI699MEitM+fXMqv8LEFf1I6KTEDm7zMIucLkd
0vO9MG72bri81EnwnwZMV/LnFhm+7bLYdIHdOaookBxAUINilhNMaM4RiPqf27qM
dESXEAwJ1wfn6PA4VwCt3lfyKTCctTCKpprFCT/YY8luw1kW+E+fZTRjAV/VYo3c
mN46LInJ10cRCWdzMQbEGQS34PsdwJNAbwl4I9m4CZK/f3JFg908tT7uH+1Urd3p
tR2jKZIsKVafxtnaFOXZZoR+4iuS1SI+RNEBodvaa9KPI9song/F+tqZEXMYAn79
LO1zIjUFj4IkDDeSGIFxZJMg/WpzXHGTiznRiUiij+t5DLQiFOiEm5WukyDmeBux
CSOtjJwiFgr3mvwM0mi2RiqcjlFJFEepLQ93iNvm06FTdzD+NeOdS61NSccw4a5K
dIvZCYsVEOPGBk+Q0HbzXvOxKZkZeT4Y0hcxJIPk6wWeUF7MZK1zFn2qSfcYl1Iq
FYKMRdaiIIzpIitdThXpDaz/T0pAbYvt7ahqdA/fOp9dZtxacwFAyvh+k/GCFgKb
D1cF/cUIu7vtVk36RPgPcOwLKPRL/jbxkEstedvD6UWIaGVhRcJ5bCJlvOJt7BN5
kffwRWajKjoEJQbT3vXMWHu8mHeufBG45vBqJkzXWTFOGkNnrX8zDfKxBm4pYVvQ
22/7Ht9cI3s6eIco3eJOhqW/he69mlx26SjP+TeXB1tjJFFy8IlAC5y09glCcL3t
0GFLVh8VK8DQd8iQLyXMe+dp5/U+AKmdn0ABSp6Jcp7GlMMAS0W6FPuc1Zm8YmY5
0KrFz16wk42gdH/CFihzQqTLGBgGMI1teshlcOKD58FnNrjf+/dT1s8oIBhDKO4L
InmrM3pSwU5DZbsF0cSLhSbq61yTBMPzZoqNyDLdrZGvW01lQa6ipMNudJXPPKxy
EjqiLb4N4lFpVyu3ZAojYS4fcp1mmVIDt0cnpaxXHFGRpBjiDLVFkA8itkSB5Fyx
vd0WyY9nKW7yeq17ZSkG70gjN7B36gMp5y+ALZ1phLdAtlDQMw2Obh05ff2ZJmiF
/E0wR1IZaagGwp65sqn25wbWFFsTTi0xP5fdgfgUW+jDdY5DCo9FNOaZnASBNK5u
pvYRfyqRxpItUYN2hlgAljco/Q1KiY6XkxCxyCO9gVe6GaKA6QpN8AuAGiqfkcu3
WNl3n3ZtU8d+j32qTo3/Hq3JPY0fYMQ/u+NHg37R94ox+WN6M6vj5dhxPgx3ymVU
gcMe5q5CbUGv9csYlxELD6iNk6WxaPn/p4G7HdEfSHVMwFdqmGYySzNS5MaV/K+m
dOsnyapOyEYwVqzlVD1vm/Ymc5/I5xpa3y0Ayi6Hqi87plSWJUjCWcu1iypN+Eed
IOTYODfqacFwdrSCfTv0VPnqcrj3gRa8prChqrAK0SXXBKRj2La4xK3AamZn0oxr
iW8Zh9SnOvt/rMSqxTFvKgqlDL6qBBxGRb3FX8Jr5dN0LqwAp4n0c6kuWi88dADj
0XokPHzJxfxsDyM1UnyK2w2ZXxUIVOQ5+4eYpQ5OMdtxwFoAJi0wg2PxH7DsH5E3
i1jhjKHvpGTe3ecwHoX+Xv7jNTamj0NKXKBJ7sdcq/Yh4xlfGfnzOIUtYvi4a1AQ
Kpl1B861g+OUNDmsh7HuR6pgEIuJe7jz66WVXi19PZxvgQH4bvA3c+wRsQqgxVx2
IKTw1kVATEkW59mJiFLgCQ2Szmp/hKcemC0tHKT5Mc3mhTgiwRECzDbSJFw708X4
1Zk/KLAqs+w106oBbz0iwWKFivwX7o9Hy5Kblo6ZGfxCreojJlQH2uWPzS4qWoVA
W3XpKfIVEVpYKVa9kyBr+lf79N3/b2vQBUcom3RL/OHqTN/ndh7VdPnQYZRKVRVC
ke+OgFiF1EEy65XAoHdBbBVo5JArAL1n85hxsAD36fRGOnojVQnVZ8U1KIpKauU0
Hxu1sL3fOneKX8l4RpsDHMhtykH2q6Y8wDKhDu74NfmOii2zTGCp36WwRQvNasJd
NG9yuVALdMhLhjtL4PUS6KLqNSwbcX3xTuevNxFjCuEmclW/LcaIwMvmvu5nyh5y
9ym0RJgU8x9ZE3FlEo5vbVprvs5QvxRKIURw4YHiPPCCAzkPX0cGutJLte515hYv
sp/0wZVK7shEE94Iy62urypoH/c2jmp8j00j0WjckswgGdgOc6x8AEmXOvVTDkxT
OnwZ4pZlyz/A9hFcoVgchvL5mC+eYCqcGgqdNjnPJaaWJjCI2tNM3ED/q2SRMrPZ
ouToefjNHig5LzaBveU67m5Mtd4eURI5zhEAb4q1lzSJi/NNHdhAa4muGPCP2XPC
+2y2nD3CvaZ4rTLeLVAh57JIhbAwhEK42bFrP1oFkqgUngHDtDE8ZbZHR/mC3ZYc
FLeyoid5VBgFWmcB5l4E8R1RjJJJQ0aMv1vuGOIKpfcyhUNX8u/7vMMsnvfB+S2A
BGaBAw5aF4JieYbS+R1XCyjXiV7R5Xvh2kXw/2HR/uSzYaTtji7VAWgnUFHlQWN9
ZNjuJ6qBMQw5dvHgoJDVyXYrILclzMJ2Zj+vtYKnhMCl9iQC11aURl32BLhUlkMm
5NpoMZ4qSc5+/ayuuhLCUGJI87U0RQOlpqVlmdDF4JSuYCc6cm0ctNFKzFvgQVY+
J85tGRw+g32xsA2RpNA1lbDe41+SAasMd4DyVu60UQgYLefc1kcxc5w34nFbvK+A
3jWONDH4I7Y7j73WbOjRV1vifkZ6QY+5qfKJ+smhf8lrBfEbnPtNnlp8KOeePgJG
fo7SWeHTqKxn4xUMYy+Brn+7hCY5oKizBqXlkl2HS6spoEiLHAgeziJtcxK5iedc
u6wixEwC4FLTHxswBiDKCPTH8sdrR+dIa8r8TVGS8H04wQGGgw23mJb3rW4PEkO5
1xb3h3CocN6O2XYVfTPEm1pR5xt1mLjDNZ9z0+palTYKx2yRUTBXmU/WPjcIVFNH
F0QN5bm7DPv674VSHMS8yolmoC4poqb0rTRU9qW3+fc3WOVcm4lsvqmwpfs9Xo2Z
re6IOQgB/7M2wtDQUuVwsb4K1HJ3U0sgDtsbc+eWS3TWAn5jYD2eBdqX4MiqZ5ag
46Hlprxmiabc15kdoI9iJf54K6I1O3R5TAr9EyXPZ8bMqbZSrUKLwVFFmNT3TREZ
ZdyjM+s2BXmEGB3hnKwx92LBxga8bLV2s13apONHwzD1NST+b00bH0vR1P7KAg6M
tEoukErbu0WSleX2M+0rsrXkSlf2a8EP93+DrNUcIR5rrA9kzZOeT1CtdCFKwC2T
a4X275hPfUKHVaQvv5xir32BjQigrjrZcOlrJIrzjVO1Jm8MlDuMGcWXL1ule9np
WyMAK6e43baUp56hqV7orOFsiZ99936AKzWWwkwDs3laFXF8z0k2M1LepfspYuJF
iqw3eOWzih1ZPE3yISwrRKR6RDrgxtPWnV3Of7/7qNOZ6mzMCBvtahSUX85gFX+o
TUi8X/Sg7VM+5ze0m43tBwzz9pD/eJmAd3Rn/rSnKpZH28yDonw7M61abo0TecmO
dF3enIiyebLIqtTfB2sJDR/xN6hP0SR7bzEKBwL/9ubjy2uLeg/6tqS5smTBjdWs
UkyB/vh1GHyY+t3ObtX0BthuvTNdRFROYCQQOvHyQ3X4X8rBofHEnq1+V+6lbFGR
FdGitlLQydksQXQO1YDFYXtV4+gUnJFpX6K2a9Yf3i+vETET7e3+8SvZVRW1c8Vd
XCTML5C16SKEYRFUaDC34S9IlmR0ksw4DrhGi/LgR0bpW5wEG+PTuwyMtrcYlzIy
F70W/aj9g7JgiQUM6L8qMTdtmAYd3r+LLvxAk9wxIstGxqMJg+cZDhptdT7/yI1V
1mxb4Pt1+KDZ/aQDDB9sWgq8qNea7Hv5JBmSynfg66X+zdF0EHLpWl1GiNKQV+s+
vp3QCppihEp/P2EX0gAUSLKL6WAvidydgERn42i4Rf/1/mIIOEhxVe27/gwr7FjN
oKPTWqSDIZRlJ6J4f4TkDWJwXKBe7QpNIbZK+octPn7/T8TxcJSGRV0hujfKhBWY
6A4RCy5fO0iuWYwBElSmF8Ya82LIkiVja1VgQhsXkrcQGgI+qcjV+hZwCetc8ehz
PUVokU+gsXxGfvTwa/lsIldSFfnBjThrO438nnzerX0CiuY33GA893AuUx2tyshd
EgwRKTEnmkGPuMhmIg7DdXz7s69GsJcIJ48BKRM8Me7ylI7gKt5qR8Hln1AxwTMM
hqmML0eskXbZX+2ZBFBBppplBzb9JRIetYI02CHqn1bsj/VnfSnDLsI6NkZgEsgX
KuwhOIb7ch0fHNLGRSoB8Aw2NSahKfxetpdCCZeI+zOi10AIIRIxjEb7uDxCl4Uc
P63H6AxljItZSCQko7Md7x0QyeuQlpc4FMAw+QspulRw32EKqd/MaXoHTeCnhUj4
1MVX18Zme++Tl4y9zRbQb6G+FTHUpSPKeFpxpXHmbCELd62zgh+CVMCYuzdbQt4I
oNQlduPPb5bRZaHSnUtYgBzftDDbNsF7kEMNqS/+ryj3jaL4DfakhwZxbAtvdHTQ
vCjKcr1IkMYRvcmCHHoV+MmyTIKhddW6EggnlSzj+ZrTFcjsYCBi0u6NKIM9giGt
H2K3cm9FZLZ+drgew+udqDcDjpB0rvvpjVR+KiTaZmFQTKRZfopbVe3BZF8ML98c
jvjsHOOiiOjCgLNAbImRbjZuE56uR6Eu77fVkS85YLeH0N+OC6MpZQa9k1Mic/A/
3bGBM04LRfJjKnkEK1NaPOlc7xIPoOh4Mqq7PF6nCfsH5yYNFyI6uxSh/v9NpuwD
2vRkaI1IkayQsPhi9WBZwYthQUWyvbXSsoF9zUj3N6WDrzXVVQS1VMCp+KBl+x/c
6uWh5lAwCyzLD00voveGiG7JuseuWWwWebVU6gw81aDXJqlScHl2wDMXMCAhoY3V
Oz0ljDkwcU/am5RSzpux49K+RKOy3i0gtPkkwHuWfGde1cXfJHKqxGUKz9fn2kml
f+7zHp9AtCbXlMaKCkeza8If7zWUDrgfb7T9zWU4zSEDWU2agVY4rXnIXmZ5G5f4
l+xWhoz3mGwS353kacL7ApShGlP5CYul0nsR0C/N4BQybIUKpvCifUlcYv5dhuf+
Vr4LTST+aLcWUSL5m2kF/uGs4WOcYxEBLcOriLBsALLvohlvp38xpKOuZ09AEe1n
IbaD0Sy56HGC8Nt3S4kQoFS1HRCulD1xTO2GRwdXIL6zEQdLFTyE6lfqoMrmslVP
xmRmgUyeffXtmpqBnMeEWf5qZpOtpqroCcbilTrW5FrTJMWwwgYBlQTLHhYakHNd
K7NoU3R7yAumyb9BBZOIpR9QPhRFE0sylPfug8NZX+qfM9ay/V/QhtL3BYijHesY
QqU97cCT942EYkZb8/GVo6qXZC3WgN8Yhp8vUOWZNoAiq+Xq3FFFv83gmjoXfuyo
Np7R6x94DbEvzahIhz9W5Ftnz037i8GBrnWQu5bvLRPvMqDEOVnIBNnDDQFopGit
kI0+MV7PgtK5FNQZZmg/adpFh3E43Qu126MKD/FxA+zhU1jUh3sDQ4cAtAEWKPiO
5cBfXU2dtiAXvmj/NHhxWiMlLcyZdF5lqbk3kWmaL+vwfL4cOjq4z0Sv92Wi++2V
Grk9ekml5NCki2EiyY+6AuQ+OfvE9HvuPeTPdwMmLrPpkszJ7hXuJU82LSs4qct4
WEzSAD0jLQBsZUBFG0HPZG9qHXoQcCX8+UcI6YJ/GZp1ehtMV5vtZjpxBRhjPOfO
50FAMWGqAL0lAy4ZtxO4CS9xIzviYta0t+qrvm2MW30GJAMtunDpczo2hHk/erMY
vj0s6UDEPNx5ZWMebLWJjN8iHWepjYR5cFBuq2qZxMQEcSIU8oHdqhZncwK3MYYv
GGBnz8lBJDErejL2T3CVr3UoBSSv1djpECVei+u5GMGs503rO4yzi4Qdj5UGzqvj
wzPbPnR4L91WR0d7RGeNvhBYlfcEeVqcqib5vDTtgrSZB408y/tV63V98/XVhS5B
y4qAwZXwpIRese81yY05NDvmQQjF1ku1N0v49+Hl3Z8wPiK6Y9QHhRUexaE5JfMs
eW3J04JSw/YFUqWDepoc2S1r3Ulk5yFStzuvSJdXJ//uHbl0DY5l4YdE4ndTXz5f
aa+/cW7cSrblDw6OY795QV7t6NWlWoeZpe89U6RzNpwwWjsnbLmHK/WOXUNPIFyU
TWA7wLVeSi2iNXFOa2TQJ0s4+uA9hy1kekBJLc0aCoCf5K+0aL3mdP1psE/ifbOZ
PQJQRuqHNIIlvcXxh6v/lA8jV3UMF/8J9RZjwSNuAmknrInat+xRv9LCcws8xPsi
shBgnT0EyINqYKflqPLtyVSOQhO2qEf5BsL2qS6HM1vFzHMknZO0Cf9Q7fX6IpYv
unC7bIsxLI32n5/ipPBfTWQOrbGgNZ6S/qecH3QdMA0UKUbxBbjB9tB0P8rTDn0d
sbEL3m8G3Q7HtW7yLlfJi+FHyj6uHTgVnmAFuTGb4BK0JutfL6gx4NU9MHJMFmcE
nG+5WCen3zf9lviy8oMtrvH3/t0GsV0qf5GNYbdbDV8V1ddAGEU9G8jJ5Qaw0uid
9S2vCv+nQSTuXQDHw939eNWHX5WXH08M5rlNsnZVPrbJHLQBoZUWqIcSQNGP9FuP
5JQ1zmTECekalAIAlWz6zdC+BAwTDKyGpGFTyEzTeibV2Utvpzv4mh4XbBFu4LJl
w/Q8UzbmjGSjA/FEP1jvac6AeUwIrN/9nxWcih9ccvULH71Cey0wGp44id97bfKU
Uo7HjmTdiKJjzOkNlATcidY01p51/DeTepKuy/YNhqiv8dN2xEVciqjGLoiDHFSG
YcwbkX202t0/2PKtuVsVNacQ7iF+0O04oqxRaVUAAz7FC5bDyUfxFPxgg1XoYXsH
XcSKu75fzSMRQHY5yjUdX6ugdY7aROcWstQw8mJLhlLAG9NaW0GajJoD4VatUsgw
l54pilqORAOtt9Gxw1ZDOb+GkYXtYXz4/G1k3OqpSDTM7vdWQZKbBDjbQ5VRojEy
pUCVEB4LrjJrWKJkHMkYGnRNQGNHtBUUTeqnSCHEblAWVOY1tv291vdzfv/g4x4Y
QgJeNQtVAoZxqR1IqPPDd994j9JT8tx9+nCS/Z8+UCGpLgROFSfY4bY82YFyFYu4
Se+SxQxlCAmgR89HIyw3nQL+eOXxTxXU8DTCZA9J5uTZo6wo5+0fxNW27H2ET8Ut
DUdItoSxUo272+F00tk4Tj9GSXfUixEE2+tpGTvcsNycgCnDOzvJpMcmG5jxTjob
8kvfPcclS9CyO9NpFtd+gRbEm3XTkt3nCQvBe+D1bYCdXvHv+WGJdbiEJtOELveS
n/38Ife7Ok1GpvrbYew0nMqb0Tz33/rb8GkaBzRVXRBqjfvt2ZmCKLLMNzO7i07h
5REJFiuVrlcIJv/NSGcj8gz3VIugBXYqWABjMBlweDAn02PvnvNK9KG+lxiEPkiF
CKJyS8ikJI1K+ta/b5Nys90Pfs/gKCCA2ThG+dm4lqYczPoi1M12WUHO0DdkW3NA
hBgcXFkD6eFapLzVZ/GI9m5u+gK10PVT9meY9aF4YL7m0CdA95xBha+pKRXM1HY/
7oGj7PqhcxSIZETW8SmJpmjzXCGp2ivTJ7HJOlbszrnTJgeDuiUTda9wDfAYn58L
bDgHIShKUSZB9u8rIhFvMzGc72Pb4hv/XEk1ziGOCIV2FV2Ld9/i401mTTo8ytSV
MWmFGDrbyvROs0YIZYgp5bNNBoiXmU0B3g0g3zdK6qGnCiZB6W/MX4gxrENHfg+v
AuMTq7JM3MmepdWrA3I02/gHt1vqOEV4WoF/uyTjZ1/xdnRlM251rG+66YvTrHVk
Nxq2b8rpzRVSyshaGrdCv+HQRWm3thWNt24jv59zErq2rX6mA7XZU//oCKNRrDhl
DmPDiqEWCzUJNEllO0Xv4qjxdYJ/OBNPSG31wwHdzFHfUshp4sg5NJ96ygO2jDBQ
PGJkXI1wcFE/NWyAntaevqjIJ79c+WgE5cDsP3kL9qh6ijO7rZ6REFiA7zMM/n6z
q9m5/Pi78OHUjUDcCLCyVPWon0b4kn3tjeUlLmHd04iWJT33M9H2BgRvD4UD7ydW
yR0Lpi+NNhRGdJ4u05UDfa1vb0kGlwzzwzjQraZ9F0RCEAGF5I9jJlQN+UvZ6LFN
pZbWYxJ6LdTv1NVLYBb7CzKDzWiwUWzaZ7WkzCzXT0Dm1CRwK1wArFJ6psU5nK6f
qWqUqeOHSt1CNJqLZzTymso4DJx/ccffE82aJktL6HxGbTkzfOnkikK2PGVLngDs
QjzzDZHcAhwnXrZ494Rm+zH3Upz67fYfKtsqRk6DUFMkUcD6871ei7sXwDB/FoDu
GKW2LdD0Hp6A347uTGAwTJGsvOsbFOu7d24hikiAedrHIdiecrC1pn83fyDNKmJt
8HBmoCQz99m/7BnPwm0h8y/xzwc1UEU34DYhoIeiRKbTz3qLHTRBkKmWaBFucGN6
IerAC2Fht1Eg0M4i1nvrb/NEqcS5f34Wb138XBGT8wQq1lzyMsGAVOeOsn/LPPBf
mFgef/NV7189WBRDPZuKgkhEbIsHJ2K4mZTVZkL4h3rHLUoAHTAmePJOeTmG7uzp
ev+ViqK5mieeqpnHIju24TQ9EsBey3xcKdfBA3iiZCXGTdarn4ZXkOfkhRRe2ZF+
0DIXOx4LoAxWpgZD/4kQIqiQlbbI7oXhL7QW10rtSKuVhJBsbnA88joqr7PHDBIn
smkG4KfSHAQNwhSOKMcDerQRjJ3xOaoD9HMmqVDkJ5LUsM1gfT+lmuzdLS3ngHbl
laVyVIp4oLZGrRExpl1xOE40NZPbZ6PJd+92RIEygXLa+svWwznZzZXEI4/TPZP/
r6rOnFIwutruV1Js8UETetz+4OlZrHh9zihMbl6H4EFr3s9hURQ6ghXz8mQcsDhj
0j1Q2gVKvfN2nn1DlAYHQXN9djX+S2bcUE/ozjMWQM/10ynGK0/kZGBff2f7sTZU
oEN3+FlFjR9CLhnWPXg+J+2JARNNbFnZm7dwe/RmuFWQi2I8BlGokHlolU+AYD9t
FFBbbVfz9yiXhIBYiwAuKuB0haVBGI4PJ3WMPUwjxW0/t0G9sI9ruCNn87/EhRl/
+hgmAjB/25iDKPI5UbNhJZelOYcipK1uYOxdsN82JpLoDiXT2vyXgRFkyAdBkuh7
MZdmNRKKDbd0ODrKwYNV+yY64KL7MyFfKkDhrV7Q2iAZOjik3rL+9PpQtIWEF6rb
icyahJANCNCaYADpJIs/WXX7b4A7GzfdJr9CnFrWSUXvvjdFBjbTwlPFyuWrchak
EKif81SNO9TcP7E5yPhXgtl5nIwBQK+dwPcIhbzDhyQLHRNzgXhF/9CgAmsplIlW
kk7R9XSLRSUIxzbbKi+ymvKvHbWV1kH7MOxTP0zEcnuTC9FeK6NFnogUP1tQD1kF
aBvoldtm/xhjVikzne9ez8wD8iL0EX4emSXHKiVKgCJ/+tJViqW6ZY+HSumn0ReF
s/3lPBgoDA7jcu85F2U5TLG+rj/W0U+gJHMDZ7EKH5fDMgZkscgu+FUo7tUbXgs9
+/Lud63s+9iEfpIyqVJ63UBC4Za1fHmxQ30Ya/Amf87Is8OIIznR1HfYEmbxFprk
fRVYIorhtkbwjVWJE/fcKkgSHMO/wMN0olXJHFzp+NIMjm40r9RpcFEwCKusb0g2
bi3Xr1lYWpkX+655wEnj/s3zy1MxZ0UTYDr/GOFiswCQkVvUSAgdjRa/IJ1DBbBR
np0tHlv8Bb9YzHdwcRMnsnZQtY+P2eNbl4EYfnY5gX1UQjDJssXv8AsMOT10uJO2
FRAr6GWYA0etoIjx1MvxfiDLx/mA1SwE3fGNJuAmF1BXj+lx4lcH8pxBnAEl3GzI
jMMoiLiOwYdL/VNtiXuM60NRKTg2GZs5sGAotrOM7cffOG1mPJLVxzIPLPdRk3DE
Hxj8uClMgyRCbb62nHuqryUjC/Le2beIoUdsbRcRX5z+a1upAJBoZRMhlht61T+R
NSVHdTzCKiJLfWuGc68ZpQ6z4Rl7A+j1NNctmcAU9SYe4BUXc3Bd7f1WZm3OAQ8Q
011nZOmJ1N7Gms9bjfPZwoQRsYki1pNK8lzjNZAU3eFA7TPCetiEY/IiOb2SsrE/
Xk8DgVFQqovm9ObnH/hPE+oc4/J525LcwzUw4V+2ZjturzGAsrJ/A3g+rjl399LY
SGOGw8Iq5WD/c1crF4Jv1yOBwInowR4gYVxf492iANpwnAGgmgzsFCARHnHMUXEj
MtwtIWpzPwxru6tlJqw1YuT9WBlNV4mNJFW1g2b6ye7/A7zii1G/CzDVskt30MnR
UTL6NlFDHA4EFtzZEl+WU7E6a1EPQdv/E0H2pRamidF9T/j1glJCudUevNzuC5kg
f8Nd46mA73DeTxrdNug7xxWGP1sgxIScO/AOsc9nwbAsfOuqtDVgDN8pn0m6hFJ5
r5jtgqnvkKzVqQffSAiNaMG5XSBGtKDk2J/aeZvdHDIHWhv4Def3PEc7IFd36tH1
rVrYH7vf/NqJjyEFRPtT+WDlPuNYRftdYeVecxIbSbylEJ8+i9S7Wqz+eLU1iCj5
/M/dmuEF3XZ92Cnmu3r8Eeck5lMASsb6mD5fil+VXFoju1URu4/SrcyoVuPJ/sEM
kCbQvvPF3WlWMfv76CjgNzgSj/H/aVD05f2Z1OIooTeTM8aw2Cq73ebDeLGeP/1S
7EPauUaHP9hnw6VrTbv/IeZq1w6vGbymuRAfKtccWwT+C9jK6lpNzXwF/3GOcIW6
IEOu09Y4U2ckecDIiguIbdecpE9GnY22GRKnPLJZxOdm3vf9UJBnXbd1Qp3uA9/0
PJEA8JHEtz+N4j9WpBNneXGPghFbHo02v3Wv4eVIfjrOr7vIDhT+5+dKgwKZ7m/W
tURmPa72ZM2zbQO/H0wpb8Q0OpQP7Smy1PX5fJBdw0xYF+Nqlet3gpGI+IXo4Qhj
PHQv9+JnVeHocISJu2MnYWSEqJTZqw5wOHG/hbjLl6R2e8055sRpFxRrsySgPo2d
3fLd0YOuQn9+H9wwIolEmo8Af6W3056elCAHk+sS8O1jQbYCtZFq8J3haMBd0m7R
T2iYZFTvDuiYXJQCQFylDdmRlz6gPo64dGvGSG1tPtuTC6vqSXtgFM9cv/nMwA08
sDZzB63t1Icm7n92J7TBrDzd7nhC5UgkW9/ZZCyGFx/9RFOFJ+EzHcLhF4Q+aoEm
D4RnRSt/IlHo7KEDrb5LKCAf3EAwP4B7+6+qOQO6cIeHYseoh8E381GwD5XfPlaA
Zdv6qBD2xp+ojaLEJDEtDXd5yoeGD9dMVoWu2xcr2lTvaA3xYUIPpH9Vk8Mqh6PU
CSviIpbxCL6TLoARJJVLzq1rcx+7HghJWQKAx1UsTzx8/BT7u20iCUFGR5NJtuUH
ipcSa8XWivDfZfuA5aaLKPy8WoWHr+3PlgQN0CxwleHO53lA5GR71l80Y0AN+ZUq
JH9ByZSY0DT85UppsUkMqUZOV/p4t8oKDilAaUW90Uwi0Sm7jZU5aMJ0emkUWhZp
nHENFkC1TgB7/0vGUL6tk+Ndjf+mcvIIEdv8FeD+NWbUOCJJLWjKEoxzrxEWnPrn
d7sG5yn8lUMnPIiEVtY9YeMy4r//2HkA9yqxw2Q60tvLDCo1kmKJmCUfp6kp7TLR
e3lavClX+kldUVh7UeVWXmqCczSX3p1KtWZwLfcts29/jOMnhBIllUTiPfPPsIGs
Morz2iW2Ypubgf1/7VKwxVJdnsBP3VYjzxaBCwNOFdAD1Vc3zPMz6DZcNDB4CGhu
4FmT7K4720lv5zugl+WCHpOCCyDQqwaML1kJ6N3LXP6PmdY8EFMLBxYVHy/fvaDz
2sQOjrr5vGsw6OGscuhEcNanUZUNK6Y8Ks5P7GL47lVW+QPSEJ//4QPmp/sLWFDm
3vPVSJ4MuPp+i7NN24bHkG3rSDqw7+1yzkiUbVUzlo8mM2FczcrWU2qDziG+kZxS
W2FEorgg1Zr2EbN2gZ0zucgEvUKquMd6odDg0rWPSD+i5Mvu7eLMrloYAHgsbuhu
BgAaZZA56LxwXZNGis+QiQhPoilX188vvYvv/FPcf25/KbAdNaSPYC+x9CiiWRIi
btnO0SKzpGH+F0dp3Ct0NZl/lwmzjdH+Mhv/+pEFUfaazGXbr+0MXcKzEXCV08Z7
6gAGFn5k7ahELfyqDChXXRCJz0UNTl3abLs6VLqt079QtVIRD+3TFGmpYZi0SqaT
vJH5UrsYNnM/pJ+XvYuK9sLiiuUs/KyfVfNbcvUnfMeCadHBF0jobrUgbXKB57RA
kpUDXqxpO56JafaU5ZUuKlIanwJ7q62v2sPtQh8+EQUwnPkGu5hz7MY2+Ee2aRk7
jK2ppTjfqyzGTFKLyiQep6r/U82KnI1SqjUBAcOJ5zmuGHnnYcNLId4+C/JHUT7q
XVIotzXDzwwqKOIqZ/Rl0YnMrqraWiNkh2XaIufGri66IEoTJ3uW7N57syRRw4Od
uXXWMit0jhnwtCq2u5/hcq3FuINbcycQiuAor93CJCirPr57eixv/3n5yfdX1KNa
42YOWtA26TUwF4um+YT6p1yDKBDzpgQMgE50FePZgmW0zkkpOzwfVohuBlU/5MFT
/fSehsAJ5hfW1RJxormByHwSF/KN1to3Llm4QVyC5UvM1YgtT3RjKMS4rMvlXRNI
VbVLaiKDhiH9Rxznh+LMUTo2Q5FQOSg1Sl77TwlABE1IM/r4ontrY+SEZCa5z1w7
HAJtNRMKIgnPNyAb/a7wARtqGg7KG9UWb5aN7vFxSXFMVJUzFm4jRDRFpXSlmBQE
6IHnj9GhBX726C4Ah7X7uCIZSsTmaVnfK/fYK2AUatU7Nyk6JsVSNh7jYAOuHx0i
WlRpD+fnpPkfXstG9tM6uoq75WHiJY60B01sTmd4LsVLC8AMAa6jSFKHrPHsSaod
9m5DCifLFUajesrZO4FdLJD0d4HPs8VJGV5i1FK7FFY3AWj3sLhLnZxE8hy7YPTf
IVvsrGqjUfZepfh/POs2LpVE0xIQvLKkpGLV+31AkF/UTuQFOPXDSWOFNU5QGAKF
tl4xBpqM0sas6OlOq5zMeeiKeJtokaFniXJ2rmlcg+UdH+Eu2FG5jyr0NdVSozw4
xtmatP08hNBP21TiZAxbe+oXMZ195kNPPMR/+7RgLBd4yqSfMUOHn/aSn6zJ/1Zq
l6O4Zm/WVOETtoMw9uLgftcv9mkAUnFDB9Iekfqz4CHISle0W2ddVe22zfU3t8GF
YFGs0i8YfMOR5gSXAyJu0bxMNOIN6bnt3nNCXAWODzYKsGeU8BS0EfEtEdvK3JxI
SHZcLWwh/EiQi6948qnokTgXAr5CMEPJgsj5JjIxt9G7kkvVKq79vyiN+2cZz8LD
WvTVZjEN762IBahcL8w2/05l8pXpSSqJorW1+Yii8jnIRwNsd7Bm2w6NdYkVii0L
hN3USXEVzSVJn0DgjtV7UR97jGqeMb8xtO19bRfl4mHbPlePsk0t6Uc6zMUtEFEK
wMOWC+naIwtlSkyJTFZP936G8Zx61p3s2WqnZvLc+G6uy5LHVx0a9Q5t2T1TmkD3
zFyiRSIg5XqouA4LsQJGBCLVlF/sVJknSBup/fcq919eFjWM0s2FBht/CquS3uwn
5rkVxIyV6WdfYPfLjUn1D8ltAeL5+XcZl/F8bDXN1/zni78xwFPG+rbGpqJijnNV
PLttj8H7H4eEH9+UliLSL9vZK17YAoav/aOMbR76nNp7oh8tN0c9nsaClii0SGsz
dpDpatKGh67270dtqxG2grfUFwjtfxp/BD//2GdF+O1m0lLJLmjN3VfVaUOXSYpG
STx8ZKIrBnOTnxxGofnQKdFqmoWSvyrPa1OorcruFE0S++zThQY1DmA3R8WEvT64
0655ffTD6pnm9umv1Y+0PJ0+GBbQgu56JABkvHtbcu8IEhjInvpXZUu+c9CfDkZh
rcQIv7/oGKhvrdd12dta77nnGyRpHjUnisfm/IaVBAhTnwz8NrDJHbvJ2T/m7bLr
s59wAWzIuxX0xv3THsOTNhYhCPFHHMEp045qp/sLRQsgjII5SX1a7MGJ/zkJmhdP
L+6pjclwe32LgGWhwlVxdmi0xkGumd4ALiBXssVE5AgxQbsCUpQzod/onbsTdLS6
q0y3/KRIjSi/ls6RAFI8cwGKunqM4P+bXz+2QRzyYjdn0QCBk9z3anS4bEQVb9HO
uUQyluDpU29jDWlcS7hdqjJJMMDrNraPjc5XeQ+cmNCk3cMwBcvk6bIO28UTEfdE
QsiMJoQp1s4/uah4wPwiCKpClWjBb7iUz6dA+6T64W9U1kmPMa0gYyudBIJoEtm0
89SRtjq7cPkdVYvL1ac+Tm5aMoRr79kQsSFVwilj0nWMBZKiozRgiW/dDYomyfj2
f9+LC53FKDojD2vk8NdH2DITREL4XJ4gFuGNMAcXdqcfynIDJUJr9M3B7Fdqi2gN
/raeMIfk8SYBmjxN/aaIS1caOsa4bYO6TmY1KFlK0qbioiHpOJkVOAODBZNxwI4I
2/wLiWw8pu0Qft3iawjfVSNKwyB0/uTDjp+dWmtZvXi24wzVsxoR7Wr6Lg460qWt
iJNNX46E/fZsrdguN0vZPtEnI+32epwD+Ab6n2AzcckhYrriVM1Ofu6dUwlpU41W
1JgbcFfRyJ0aFwQcmjoaUQZ05Wjq28rQrPv8ytNsZ3FhffuqkhG2iHiDMFKiQaTa
qNgeEsdTOYGJ409GYZovbJdOSsLRUypQg3ALtJdype6gWZkPNrBusmMUeg4E5ado
cZy6Z8QEw6A3KeXUJBPbGEa+2Ydb0ADgAztEwsopD/V2fPqIOsawoUk3M1HnPdsE
JElXhz0YBFIOzvJ6KpU/xLIRxA2Y1WDhr+3h6ZZGkOk9oMzeSoMAAngbJMMeLueX
uhxFx/Gkq6cq54Fng3sK4ycGbLj3Lrwmt8JPagSe1MUShWUO4KmSlndxLXrXEq8z
r7aA6d5gZHTe21poRwXwDvriAt78sqkFjshQp5WG5zVDn4aFCFTF530W9AvANg9d
gc+XuhvIDHMWwowAGIzfFk42HPu09PFvCFddygF+fAfBis95smEnYwbFBmRr3G5/
+3f5FHIwvtnE7PACbor9KfdWCcPP+Rx8AMETOnUUxd05nr2/+U8fWk2xrsu6VcYM
uVzHCOYYHeR7hxon/T3co0NkjJhXOW92BqGspIwlPoBdclVVEHZzodWIDG1TWcjl
5wacseoilXoGZVOmlI+xh4qRWYSYy7j6r6vvl+D/yeMFXDKbHkdoTrBox15l8bcY
NmzxiBWVBcfJ6z/NWcnftVGmve+OoypmiZZs/iiW/zjcHa3ieh4cshq9GKpOO3gu
bWeZScam79mNbrxBOLLxIXQyFNNj5JF+DyL9E+JC0mWv7Yiz6L68AbovGMSDSbdo
66RH9OTblnhZQdSRIT7MzCH12mGZ0wNB3I1ygLjw6DUviZOvFULJ0VrTn3iP6NYz
8u9dTVXqRSPXC7C9ufyAspgbKWO01KsSfF+xklTGnmZFH8zsTyxgCv9zy1U6ZQi5
pT5YMubKXcH2yZSUK6/hhitYrpvUY33jf7NYFwQdz1Cvx/jnzLUnz0sNnQ8h0CzX
TV0B2eJgbrtvr6f6zZIM6Vmv+as5w7AIluNIO8fWMjyH+FxGKPrqiW038/0RJQvD
c5RLdi3NIjGPmC22fFm4xDDm681kumXh1duHhOezmcsvFPndN/4WV9t6VitUQMvo
wHtZVP6MpcL5jMvVw2Ce6RDJ2OoT1Bk5TDaOKPM85/a9+UqUTDIabL680s+C1sb4
QSIPSO72IiotDkxOySNOGZkF/HEVYJleLkGGtCEaHcsfosppa1MN6BB7WA9kCKgn
kNUKW+qvqsq9kBL8Cu9edFFhSr1fFV4NDtbTuhvkbq/udLJcsOeich8Y+3rYQDmf
otzxe2cWIbHQz4U0pUie3acQPLBGHSi5VCe99PTUacHg64vniXgnWqxX15bF8Yqq
ci66kxY5wM7ysEydDt0//PF7pP5q4K52YXARW3k1N+PtMcljTSDgrOQKouJXlCa9
jpnGgEJgkqEHfA6XXfuEA7i5v/IoQAUXryZW4KNqxFvOGin2VHgLqpipab2l/ngW
M8o35LxcnNyMpGknNVprz7sA4B4ExbcVkyGLx562rRP8y1uxgeMFAqMakquzErHI
WEWdkNr1i9L6JOX4yTs3L2Osl6haajEw445/84lrbuPwVuHubHjt0aWXJhdgxyla
xPAMkzGnFKfd66O/vJNp2VHymWGa+nZeI30U87HhQfMmcwP6Qk901deQHubqYL8Y
WxcPzwnc8SdXsAdtGUEY8wvsiwFfaEw//lSPWgEBu/RbBBvlhszebZ/ggDfnDwJP
Lwag/ZYNvH0OF6wzXAeUatimRRdoXFUlGHZ90d6+VRf1eMmW2Pu3T9VujltyjjT6
T0VFGaZ00u7enxkLivxYLT4mAu31YJZ1TAQFnEpbU6zB1WrZ2fOXCh024IfOatuN
p/c/fJ0TjR/4ZSojycFuXfTCDzIrPspPZcPbj4h776YNeSs60GaZZ26OoYKNK18/
2AzAsUiPE2aGAeS59KEJxrxZGh1XY4Xlg1+aifGP2MnH8zCCUBxhJ0cfshHd+bXX
eEmfSTYN0i8zF7Cmjp1Y+AdJ6N7ArNGTYLc1QAgtxbg6sEXFP+m0Qf4w+yCmOd3e
GNYpq4GJx4lFDmdXWSnRespafkUMs/2W4jHDG064S+GBLWMx6101rGkLqL14Sf8I
GXRnYATm2js+W9XolIRxYMIIspAv/AgRg1xfCxkkKei6Q0g1rzmc3PGoJVM4GqjL
GJH5NN80InIm9aM5aRwUoQAOT61onp5BXCqSja+mAe02QphWR/sLe5ogemXyyJ7+
C/4AYEDKH+dw/ggkNxKddYAEVvHA2PzkobhSFDF89w0AB0YzGoBpiw96IHAosOMp
HZz8A3r+rt+MetffnxjBIOiR0eQhm1XZrK8FjJKE9FxTzMTsPBR/fn+L7UR/v0WI
iUX6uvRSVA4tPb4U2KerzdAuSZg3yiF+DMc15Vb76FnGBQIGLqZT/TqjvV7aBSuk
HdjveQ+u1i/kx5KrigwtkrhOtxQ5m0cQ7X2in5LRbtzDRafaFsfi5pwA33fBsnaB
zM76UGfRMogoPKi3VdYjmAOruTviwu2WEtsNprwl/+8aw2XF1TyASR8p2Z/xkRW7
WfLQ0O0ZgUJ6zVx/h/cRj74i8bP7Z1hAdkFeamicYoj3seoqN1qf9eTV6yc5KzJ9
zTKVpGBj9G0sHkmYEdAAc/G9O7856SD2ppBf1/ZscWQ6D9aLPtOQnJEa70sdFCSW
Rw5oQpjFLIFXiWCtm5dh7iMsitWLrxuKcFbjDwnNswx8A4C3uivXLb/0tnDKgT9r
ama29uJQg7lZiQFx5+pyo83A6QsUd2aP1vrJT5ZX4lPdVENj3k5Vpf4LbJOY7+AG
NONO3IKItVENu4vpRb7g5ajpqk+uXtrGAlM0nfHgri8uBvkyMnqvwSDzpuykw+bG
49Q4dpgfnzBIdUc7G3H7y8g/NI1ZNkLq6K2hJs0CJfGRbpJHxXeRfmyL0MQuE6F5
GdQPQhet5EcQdpg+27RPgEfgAfItDi2tlfKu4kwAU27CLBYnpC1EnOBIajTr9E8s
NHLtMVOsYGurQCjFTSSqlvX4hlqaFaS9QO6pHGiO4LWxbjgWDb5yQvNomiBHB657
mc48I3A9JbtoSJwrGcVZVuOq2FFslRbgQXukaHCfWekebCFbaaHCNt3uZc6zIVaj
CkQkquTZVyTEx09WbsE9rAmBKOK03eqhGNy0CDpKaLWktB9m/eO70SqR3uubtdq7
iRjVf9VDrMwTpGz+fdD33JIHoohS34fEB2r01ufw/qeOHzDeFR/DFHqQbev15nVa
gygEx31uwmaG1wH7mkSEcsOeRF7FYe/c99o8lyZ3oFL4aVorGO1r34K1EEbHV+dQ
Ob8YEcVk1YqVaE8r1nOKP7L6hy1FOdg46/FAcztn6KXE890eNUWZi9mtwl4Zw8/g
IM81LfBpsxtbxpoCEqc/NPc/Idx/PJd1XdWrigXutALJRqH9tJyYpR8Ww6Yso/M5
URNcB1jDTiYUZC0AzoUzjns+RDy3ilemdbK/nm/xcX+rvEm3OjAG2fxGKSHRUAdi
uaTRZ+yemI3U3LRWT1lm7Y6LzATtRZ7rNOj4lgshs6/m2G4jyX5AoVrhMcLcRwVV
7QrJRUDA5QaWJhlEdbeavMBzyTKs1zkjXWslP+Skr4baLCk+mY4CVaWTJ1zhNZ1O
8QrxeJkgw82Zqob2i7Sor1TTz/gngwtdPK3sX3y+oWT2LZGeHgs+sFimBWDaD/HV
Eg/gJIjntFXA7u/+UDF/7DWQh5ICcBjDop1md5sdywM1BSm7HxDkH+zIOXWdGtZB
rHrtTo5nPIM1+ZvS0714mKhznlvGkh36GmucN8bK/m5n5ydDIpat8lkjwB1awUpb
RGkEUpkzWFwh1QLELKeaCtrY8PNe2i2cz7PV2INfPCPy3RYlSyGuietCHGHBqQXI
BkWXPRgB5qFn+2PqfKsotcnzBIkdsuXxXWnyj7BtXqpBHbl0yZe7de28aMUz7FaL
8styC/O6+FRi4dJH4pCf+jgET7eRpG0fReQPOHE/8eXXlSurdxhCq8b6OGReV/GR
GIkFiNOKyyO3Z5jaZlDLo2UrQhABBLy4rZ7yQgWwv+szaUMwC3QiXRUSMdZapFSG
zvKMUELvmIlrJcaPRLPdNwDzLlcZhDtXhqcRcD/AHVEGyORV67f4eoNgH6Lpwh4R
Asg4ekXA7jAWJB3BxkRq3IB8MSI6tkVTy13+COHToS9ESlW/Rv2QK4z4HETVWBJW
VCrVvWtADKwce5Fi0/q+YQk5D1ajXo1fiDW4APydZihXMoM4XORDCfqBJkmGSadZ
76rYDTEcwyrChf2ZRLNX9vijmQhLwtN12/hT0NwFmey2VbTqx0GrLUFqoBl+lbEh
v3LKDsEHBaHndsg/T4xvS9nHMl4UwohC+wnBq8/Mc9nHa3D8GwdegwlM+i5GDwXI
FwM2SM9gt02ea4MycoeZlrcFuNGSr9zBIzgh5mmR7RUx8xelvUkWMipd3NdJKEqu
gkN8yWyBzOzLNDyPN534XUZsUjB5wdOjXt7TGDImRjjKisxRbBiRUVQ/FMDRaG5z
8hqfKxBQVeh16m4e/moX/67B6pNnTiwfSQNKpfVPJgW2Er2jbcAZS/DcenkDSR/O
VVhaMqK7MHFPAikTopoDLX7zYLEmL5aj3HqzJAjDWNZvHWyMKHzZayDto+FUKQLD
po78Js/Et9nxyUNe+IA0m0lFZQKy9B8tBqITqJjHxWsXvVOpOJ7GRqfhk1QjUMB3
i81ZaQTL4GUr4z+5gz3Wb6EUI+Hfn16xU9ylgf8SEqo0fWmFyzB1ajiXbyD0OaG9
Yt0do0cpunQxB7DuQbiTZuIoN71Uu3tv624m6vAQy/pxqGGL7RtOcllh/xgXZh66
DNF/OQk1khwLnYtd57TKpC+rfEVC4DqF/y4D4PNHPkbVEmugATdkPmlBYFd1Qz+M
+9nQRKffkUAhYsiR8RilYNUVhDA6ywDAZa8C9P1cnTXUh0JJsDlNjd0vWjUStO2d
sH80bDKjwlG3PBR0SO/y/fgjtnz7FPEU7UCQd4E/NhWn0tg1OzncpDvbNT9fhaca
YlBdjMguycqbKefQhPpj0gWxQ6jUxglkoIxqPpJPhw3sLRa8C7SNs/Aho0Qngue0
FAR4CWDuvp6jYIQWtWzN+sS5kL1xk/uU1r6DIyOXnqxlgAQsFzi+EBux++K6kHzC
tm6MPwd87/5ielA00xNLKqJnKf/l4jKlQWHNpmo8MeYhqa+TrvhLuxWage2t7QH2
m8rjtzrg2kacbSrGwm9Bub4QMoNPLYYcSccvj2zktGTXySPierwxgiaw2rCdpUMN
MpjxJ4//3INV8OWtBtjCWIKkXFWBmCaKxjBj1QjZWiTVdQyq+tbhm7J5LfLo0PZ2
iAJELo6+wFcvcBnoBPWcPSL67lbONYY/ki0yI888YWT0MOcB55TBmU7c+UvBvaR/
kVAs8i6Hd1zzpHKE34m5cd5CJl0z5YoLsY0FGXSB85w4tTUmz9YRDdFvHYGC9bci
Ervk+0frphw4MzlCiPBs3jg5UnFpWHoFTnAqqYkOPAqyuIAYSXtlVdM3TOJo+Pc+
D83t9AhH6jl57I7AGsifp1CkEyxOBx3TX5SsJcZPSQmbWO45sI6rqwTe/Uu8l6F4
XlZLhTzJR25JRnOz9uMz8GI3Mzv5RrWGavLHn7ElSaF3rFlk0TPW24y4bhS0+hTI
pUS7hoO75M2deyD/zdXg/a7n4Ws9JKUIPVpIO4txvVx99bcoNhYcrS1FwohN2qU4
IXc6d5H2vhdw+4Xn2Qw6UQJyF2i7k4ZdHChVSZff4sjvsL2c64ZGv6+bgZ/T0lJl
6V0mDvjzV0FKumCCOx6pdLBYs4UmcEdZThIzZCCfxK4znEv7C/BoDFeq37f45klC
Vs0nCf+Yi0G9HYg6gi+oIcvdXk/6HBNDpJ7GONCPaQvUp095fZB286XweG3+AUdN
THJrhv+Jl08AQErhnQZud3uTn91N1FLvcmiuRjVKybLHaFR5cHZThDqHKcd/TGdO
CHk7jv+M+gxNz/48nJ3kvLyhk5Z4BiobBjxiBSosV4xymOLWVO0CZKPfh67cJmPb
wnpq7ePcPjY3XrJ2p+aI/Im6azCIcflAK9Zw25Fv0clS0OUJkslONzNzzJcqMbw5
L685nuSE4z1SeZEPdjOP16Ge9Z0zVQZV4r8yAfjwcFEgfb4SAe6BsT2jc75j6qtN
DvuKZkbvRFnh5Y9X1x1CROnDqW1jbxAaC5PCwLiPk2GDBXz6HvIl8zBDSGPoQ3c8
A261KRPFnLKvk1j+Jc+TEPN7jQJBwsXW/dM9nPKHioSewERd9fvgYzIGJZlSCfdZ
SmkMjYU7/mWTOUplHJ53JeOOmSAmPFe5pK6tg9SEX6AZ5mhfMIa+0N+tG7W/fSUI
26BCkMdPN37GVRsK8pSFXY+3r4G5dHwTtdmm4npYzrWZ97WFasqPMMklDy5XnDbT
+l+QBOp18N207oWm+vHJn6m0rOyZ1wLzbsDyNMEm/ThL5fcaGuZi/6qfSXz4kOHf
OWN37uSAWnSNn2jr+nDEfZYeOVtLoyyU0LDoyo6sR7q94tQv/1Spel6QXo23XIxr
q0H6GOqIzvkBo//bb8mlVYwDoFHxk3Cm8RsTfgsjKkD4K1j4C3Q83OO7p7K5xTVU
Plwnp2lTAYUTHkB5CPCiqauMl53K6t5VxvC3o8G4qN8SIUV/SGtVcYGz8UOA1MA3
acboavPz3yYNJJ9mcziGWdOYn5XkFlkjZgJOt9SbksmNrEVa/26gbNF4I7iDtqlo
dMT75zaPQP+GJ+NR4cSdWXkms/Jn0BD7VvhHmQ8KtzK4ROHsWt3pqHsMfpJJ+Dtz
5+rLZi1XHxlLlwaz3W1gaHDg7zylvIEJ07hkWNd89ADvlg7G4vsCBNkLt/lKzk4x
aBw/9+D6YQLsPEJ9tAUd3V59hOeQw/BtE1wL9hPx2uOMZ6jhcSrAUXd6SI1sgg/7
qY4iCfM3dWml89OvD9vTZaURhqQtz7RvDw/mzYeiGsRJTwmVm51KZmqIwPoxNv3d
qWFHn7L/J5aa3WC3W6RxwuKDiuiJGifTuQkZBRpPfuQ5l4bEQD+gHO/4UIEbBZwf
U+yKKtUxonWgXsswG63oUYLFADyVNEbh2onTzHYnp5DpdI2xhIq5WtMx0fh5B4HW
tlMKlyq2BM7HF4aoD8zSNBASdnJOyVFK1h3cmfHN+u0qKmMRhTNR5kNKjSXLqwa2
zXnVESHL5Omj4UBfPifBhK88jecDvxEnXe14GEJwaQAf7rFGAPm3fOKpH3RIzePs
xo/8UrfbdLF772+HfGek0gt8LmTpmFVpmp34sl3KYyXrqq1M+y9hIw0ZAR8c0/MH
jOeTA8xfdOMbx0qL0WpTiHpjZ6q8CeGq9v+aa4NUD2s1HzoteZ/JjpVf3wfMnDC8
/7QT/P/J43uPrjJzQCLk52ru2wvam2tr1sB6kj2gDREAwKFkTqtllgUNdhfOPAUE
n/pkiPorCJz5d2LJ1FK+6+OdnvI91v6K5wDvducHF/wm7MbyIQnDGrl3lFfbGDpi
94d1adQ5i1cwYwCZi2vYjApm3rOPnFd23+GUr5NKd5yyRdNiRiWhmRPIP55cejBk
Yevo+RMFZs0geszuiwEscqmFZCGWpD60vNdaKUL6IsHNHPst262+33Qx9JglPpsr
dqP4S8v43HHLbUyCMbvec7x8rPCo02+alyVYsnIoyZMkglpjo+kIHw30CI1O9c1U
EmF/4/QH0TYCbXBhnmBY+rqo4zNP+OzxI27zx5w2fB7hulZOraQmElv5u9qMmfLw
NRtYhYIJvPHPmgOupn1zwazkmehS5/YqAs05wfEgvjtYGFjkwiF+OJVCgoyUVN5u
KU3cI5adzrwoy/B1tIp0aGtUfLA7UMoM4h+W/qlrgg0gfop434E4aq4Npx3+ckaH
wFNfaRhoKg6QM4GKmjXlDvTmBvhbfrMqnZ6FhHO9pbTI5el4G5UU9P2p3aBZGu8q
AqiexTAFWKpE3Eep4/VkP/ef5RmfMbZXc1O8qHdXX18GKn3C5oolt//dWxbOKnpw
ZWvbfeZ4kgRybj/tpWlY1aMyDRt00Z4Y5OvHGi0rpBjSuzYvH3qY911x6cbDxf1V
/fGY7PtiZ3SZ8OAzq63aQEHRHjbwo4PxZKextm19amzb/honZbqi7inYiAuGBz7a
pWs/j3ZMsjIJbP4jWmnFMP60neOrMx2Px9cC4WceWfgLbKA5CXqcTIFfV6A2JW6n
ZLJkPWgrzEf1xbrD6lLhXp3QTtMlWaod4ypSp2kU6TWDHNAvbYJo5NxZsccK21Hx
0xKA8y9g7Jxz02YZZ+DEufmqXBQeMV9U7RWA5kGb28a9ORr7Yt+H0Y+5JqJ6NTbf
UOjYeLdD1NbOSF7X5TzSbu2op/JdjEMCyrODSZFVy9RM/ZqEPX49bvXvU7rmE1SD
D6lBomSE8OhQYCvPgZswXuXB+yJEN+zF42ggClCRCGimfl6E2/wnTWgtr4cl/Joi
JnO1jet18ET7T9aT+aPaVtUwA71AxJGLECOqb2iCLuYs/ot9wxo//UZW+KUCE9Ne
yBn613n+Q1SSWHU1FCETzYPigMAfugfNlIYwcTDcSX6zm3FMZAMVELjDFbZEiA9J
w1Kk7qa2tflmHJGo90nciINx4JKxq1W/9tNHn7wOGPVM9vp1l1AHE6Y8IYPul6zG
mJXCxErdQCvAl/3yfMJQtJH7MU0vZcrf68Blyr7NbkqYDVyRJR93wfM+B4hgzS+g
2rHxXYtFUDvnRHXzGYtPhM/VTtnxy4N3UPLxXSqDpTbZZXG/keuArXGbJwijXbXN
VqojbDAgSR6vshNvKeDb/lVAe23yGqEXzgIoCUCJE6pTulG/mWCJaaZMtoUJxDkc
eWfLKLFNWBbVG+aVJes567WkSuc2+iEdE8QroLjmGh56rM/OEx5N9aZYeCBG/tdM
QJCPGueWdawTDnCQ89yh6vLDmRHuJvI5J/WN+zVX6iniSzWVHD6Tt+Wsa2JKQBrL
UnslcOnmFVXT7P5VE/wvO+fXqWI+NoJVqgGbv7Wkj6m+y0O3arT0pmE21sc7MzR7
zoanlAupT09Zv806nZrocXzMKZNdNVm+oNP/i9LOdKOwnjZxO+qyezeMABOKNtVU
t2DuPNu9NCX1s+6fFmrrmMeSIyvbqUGX14Sk1ddDOCCi8+a0PUYakiBPYm/ivBTs
UDh5ofIFsY0xH4pMIrK/umqPVpk+K6yTLPsALFBTvw/ox0Y31SrWCC6QsA/yX3wC
SP80zQ8cb2LB4Us97Wj3Ak85MHwueRIodIU0wiZSRJMuPD5Jz8F6CbU0s1/raqUa
F11c0gbOk5fVSLzbYxtuBvm3bkO6cE7T1TI6QlMItjjZwcgVKfVUzoxenrRaS283
3MBYGRXRdP3vBdFWDiQk4MgsfOo7BTj4GV74xRFcVU06JcI0gEKCRaA6878mH5Xu
KyKOUv/rxgjix+xKg7RpaFI9UJtHeyjyUZcMJq7J4UO9Wro5lQOuDoTlapf/6h7Q
5DgbqcyysAbDGNo9eBVjeZVajHWDWyjyOg0tyeh3Iu414V4KYPvcD4kldD05DtmC
0WncjhyTTfzutOhzngzcM8bW3KcLu0oOh0Bhf5CQjXYerRiLMuiDT6vJUGQ6/3/Q
sD+dqDa4uWN0YNzuFPzb1bmLw2qIB0OA88oy7oBhKXjEr09C5wQjYwbE9zhQLTVn
7fhitNL8GdS+8f0FedmIjVEG5FuBlBcO9vkMVBWv+D7TEF6DW862kJjZTdaiP1I/
6W+s7vJQm86PBhjP6QSOvFMtkf81U2MGWmhWh8dDDUzNucRebwc9dB+VHOURJNt8
Xklv25S9TW1LhHAPsr7y6Wdk//VHdKDt2RvjMp2Ma9xRDICiRd0tuM7XYFA+tKVj
EAnWcn3YGErtTwDJY9JMmUaHcLTSje0h0h7IPyNZ+tHRqk7i7FXDlyiOwggVqnh2
bu+0rCYPSfkG7KYXT9IDPyoZQSTrywUA2fOyeOvzkh6a7E8Z7JMyeN3z9G3NGAfT
L4dLhQixEkdH4H4oZnEBYzPsuDwu07Fp6kBKtb9H9MCUfLYRVDzOxmuiZFZ17lF/
A0wsLOFe7TNFntJh+6IhGi1PgxHDH39Lv6sXQfo0pkNL65jFCx8sjG3f/Uv94Yxg
HXfWKeSYS1NxHXetXhVbYOx6XsrUl5pNJTttFm2eul4cL6w1TW/Rd7a+F7udaKYG
Mmcp2+pyphfUMWqbw76aw5Q629shXKQr8KWnhr6gl3FnSoPIRSoCd2H1FD0+x1JU
rYWcYkKQGiZqujrYcW6TQMWkQnEZAQMVon+4KdV7PFUACu7ZMc9ve9bJhvsbkClg
Wi24nXp4BPxi9wAgTtijuimgpZVBwvSDhUG/aguaH9mpgzQCFOh+VjP6VL2HnwdH
vELpm/lUdp5PmNkoyr79Q3AvWAOcW61cNeD2LVUJppwSvvti3TlQiXO3BP7PxV7a
RRAq1Zi4GlZe+IAVaHwTVXOfr9M+sHVbbbXZChjaFImZziWVc+SWdkUnolGDv+ZJ
hRcZR3/5q9heNPDu3jnXWrLck0IFJnC4QSrCyCLgsizOE8eptkJo4Yw1L8+ymGbH
jWuAA0yxR9bYK6QJ8WfgLW5wO3BbajAsc/XWFuT4vgVBzXpK5RHXdzVm+zYHaVHY
wFPa1ZKApTE20bxRz3Ri12/ssX+y2VOHY+RmPoFKITZ678G0FWALy8HQLXMBPkwa
715Mu6hwyTtNB0upJ8iVQ5cL7C+Ba90/+g+CBWYCSwGJcry5s9p8s20OlON+W06G
f3jPtFiaoM0FpdN7B63IhPmbWq0sw47oi+S/N1zjirv6mpM+r3l8fy275MKtyMrE
/oRO/LW81x+zosdNBIjinHU//jDQKyvf5RjcZ3+SCGMl1XzAAISS1zsXzo+eOtov
Z6j1BxgDXWBATrauz3lGWp1/mJhzpOFno/p9V248pXGLpAyOzVSRihRgqdGyR56X
lNaHLaxtG+hQKmnXXnZcOyRsER9z+vmsm40ye6rAle6LyF4Ge51Pn2oG7dT0SVJF
XRr1R4K1r/KYL660t0W9/VucKXVWYQgi9TXC2C74dAJb6mDrVrFX40sYQyLBGLnc
tAmU+SaFLU3gmnS1PBLUczvQxJ9kSiRfCFlGq9S7eoVYs+OqjoCKvQzP3Xua2fYZ
VK1JZNuU2nah4Su+whFwpcP7O37MBLLiThAIy72F6ULxptB8p0QCTwcVh69iJ4ex
dEbGcmnQ4ODv8QpU/6iVbEPsEUsC7M9/4q4N9yX5eHiwpjnU/3sYKX/meexYQUHg
zYBuJtlPf8/bl905WTjyIKBnHmTsm8H+EeEJPJE16z6bVG7VYMOPyOAPkNYONe6B
jKQlFYCi0EVRdFViDoYsq67TQwtYduZUwKtuzqp6n0zY1t581f5KPKSLv2bI8Kcu
/7EwhHrGqaoTmk/2Z+9WB94E79zFI1Ko3/7JsZ9/ooB7HmJrDakntpkrDC8hkj7W
cKrOVAtOQ8543R5ZOCc2yAkUZZ7hAJ6nzfzmEBrTNYub9+oaA2Ace9N+kkWDm4CG
NtuyYGpyBWuMyz0UrzRxcdCJGt5h1W0hHkRM43kROjPdx/45iR475WhVRZjDOfIF
6jFt66OwG4GW6ILF2zi/Nxi7nMF9zmGiltrNQdkIIrxXqxq9RvXwoCJRFCQB9fcJ
CWQg/zIse1eIQ+Y1+lXyKbyFG6vhOAmULWwaiShcvyi36OgHomWuCVQNa446NiSi
F/WqUPvIVM5gogdeNIZhLXyL+eXFFp0Tcvl9T+Ml5Wx2dDsPeFSmq34Vx3JtLrsN
ekFs3TxxWAySMn3YDX9Ol/e9ad7qTo9ZA6ceiHEoQPuhOzAOv1D0Ifabk23ItGEZ
OeNnQEwKVFcOwmCwlGkSVWg9s5ff5yN/wkCd4j5wv717ycVHntH4IU2/o+1bYg3F
fHz9hx9GWreiiOk6UAPBuXSGWlh9ldQ3S+N+uW2B+tdfaAS3xP9S1TDp+KBPjPbw
9FritnwEySOO/p96HjelniLwj4ZfOFTxFRyuJzsie5UWqEzQgz7NDs6M5ttyofBG
L0MZPwRQ/IjTIVMuRt0XCmRngBpA+tAeKZcq6yRp7jlWBYx4WW+fKjTqE/qv6u7e
pFh7dsFYXLZc9+FXTkBFi9vRuJFCAfHV5roMmgBel64Id5Uo53zzTUrL6EixliNr
h2Kf2kfngi/9tz4TCYqU9SyBU1w7yq5Y2Gdo+nE0tgWlSiVwGn3XOOdTQ4eeUoZN
oo8T9yY3hDl6PdXqEJvEkoaT5c8fVy8qobXHNfLDd4g2elwkFxojKt36ND47pP4R
umCTreusF15h2DpnBgGEqUqxZLm/oRSbkrWWk2q8+iHylF/pOFCnIhMzmICtOZkf
b825xEadi0xTW9V/fLCVuhE9WTT3EoDEyfyRPa1QRSAfoNH5PpgjknPlV8sgnIhy
4+py5PoDUkWvgF1/O0y74veyQFVRtlEwRRwAbw4e6S82fyxlgoVtKxGbdCbvLP6i
hlTLPabbF7kaqdPj0rtoqs8a5nKzuU+PIJH8Km65kkf4QJLhmHPvj3XIvVSRPT9g
p51F+MGF9i6IHz0maeJe6zYIKJq9rDQGAmnrb/sKAjt21TAI/LR6MDjGOoZFBucX
k+jI8h64wcMjtJb7Kn5LzfZJKN9yXNM5/JM/Ld9TyRzluLkpeOinEm0wbK/iSqDv
qIsuRYQbJ0dC6dyBxh1VhB8GrISQ2/0yN7Qx+9SNA436HANAXfNTSkWXDOMW1V7B
qCUx847g3Cf5J4xD3Dk+uFV0y52XwlkcOrdG0QqgSQHl1lvrnx4l3BXUvT9F6oKY
jiqqiP3kCUAzEaJowK4PEXa1lYOfh74Jo1qctMXRMzAMLTJukquDFv48Iab/hRQq
5A0sm9h+UM9iB6I0WVDREdKigLvDFIcYs/T1xh8lPlci6oDKAIj+sBDqg3vIKik3
KrB6HW4HwskvyGPqJVM/rNJ/7gqLPa4Mb2y34poe6P9i81stCDeSYseWztI7xZI/
sT1maToI8sRmJXJ3qt5HB5Ld4931PxlY3lfXBZ/2lYGseSFORxlt5UCITEnYUdsK
ezmmHs+/wq3PNL5B/WcgpgZuQuVnG6aMONPwfccXmizRxvpFyMNz72afxxRhLWwW
KBgp5acXrP/ykRQNsiW+nXZMuFu0uvguEdPaReSui8wB1BYprMfRKhI3mpxLtmRb
E5xeHdgsG9mOmiMjpQA9IjpDKJZNpM7m6wX6F2A5XMpUBR78mMvav0TeF9guiWfs
ddHKZSikoAW+XpzXzhRcsT8Wjbhx21jcnQQJLcx+z917Y9R/Hzfv3HB+xKz3Fblj
bDzw/rP6rt3VY1Qgo3my8UowKcLFoaryft9ozf9W9CxdYMnOPPqxaauzIylTE7mv
9PNLpP4hP64mQCT8aLWDojxL/KK+cckfHm+fFhyCbASyNPv+4gsmR/euuuqhOGaq
EFSRwHCERqVAVX/wmMajhG8XKKebTiiTztdy4D3I6q1GrxuQuGD605FedRPPXMub
5ZVOX38v3Qk0FFsk44uRBKjtCqHwF1/GT44gDMuYSB9AdmEMUljxfc83AGV1vcto
Ej35WUih3/hu2TaAgE7Q8dxSMJw2W6Stb9BN3ZNwigKHdc/S2Tzm/L97pUzKXJMN
uhcgknAviJCH97sN7KNfAhAclxfqOdJw6PIgBq5eYXqTfvFWTNWE3tAktkvCGHzp
omkCWpsotbOMTzSQvCl9Iwcp6xqkvBs3oLBxDHspxKD547ikrG/Pkuh7KqTjg/6H
PTaMaul+yglR56LbMtfrsECdSp23+AfWCB2Cgu/TjA/GX/xUC2fyp9tSxiZV7HHE
noYW0xqcRUC8G57MVv8T/tccz3rLi2Us+szLXUOMETMGlp9AJ7N9deTWlNazxRQa
SaqabNO6Vkuc9Ww8QXpElXV7n5yOf4L5EVIMSSnNwSoileokuziD+j0rramB0mLC
9enV4pVHC8CJH7IAJmXrH1XnDCs3Kg8sA5AVR134gGG1jp7O+wK8VSI/qSQYUZTp
9xANNBJvJhcvku5HOWJPwLeX1biVlyRQbcXxMHpremTG8Q6ngcayxc4JBjfBWNcc
SWF8meOeD9Vy4uDc/GupTZSzUijgVbCHje5j4CVf/3lqK5p2gLFf3jrXA0cBEhzg
uCnVOMLLI7GGppQluTplk1usQ+QgVv/EUKsprZYSqRF+2qXuKwON9nV8UPxGJf0d
dQX2kR3JcTWX9/TMHQgU4P8x4NhNcpn1Vh51cedhaHDPP+975/xqvdzzupYKdl3i
fMxzMxgXruir/5Xt0gLZpb1gwjpmRJj7P+RdZXIkP8VDkS/7TYw9bnGsrIcIUaRP
hmQALrSOzptSQsrvj7xjeznZD5Er6jjF5898Ohtjq0muvZGFE91NJokTntfRsThx
DktCwuKN6wpt27CC1RFwzv2JzoDFqqoh1PFkaFkxuZlRYWMA43DUAxZSTfBa+Lpl
RZbKKgtmHSXVmci+drgVoIVdntYQerWikpm1qoS4FKaF1D5VxQLYN7NkWuekFpCI
Z4JgpkG0Z8lZp5DhuLb8WWX3SulU5F9Yfpuo4wMMhEk1AgZdDLzfzxgI4aC0HCAh
kbJgd7SSJJtOVvGeLsb0iW2rqwX03m/XC5131j28C24KbXiXP+Esgk2PrBMZi4wX
dSs00EKLmLDNJsXs095pMy2mMPrIYcGpouqDUZRvXVVgOVa/BiDF8cyqhQ8JLBLk
VrPJPub75/3O7NcJGkioVhagMLvNDn7dFhCquZGXzf6sNT2lV7FExhLW1r7FeOQk
qLsIKO2dLq5v4LK1cV5uBTJZ5EvfjabtfsGzgPYCqcEMfqvw9SQGMVEqH/OZB6vf
SY7eO7GCfxlYK7qwH+j1vl2Do+BwlpwRIFJbttFyOyEl0gueu+w+stjEgWMGe/ps
s81yQsF8m5ufklvl4HvJ/EH9bRLcEeSwLa5uPKdAE0gH7XSdh6t73QKGLAXFRbJI
SwNKdwsvv2UGUsQuBQVyPS/lTGg6uciIORXBkTRuw3kTJ22FHmqX0gzn2IIn7l6D
3me4JUeT8WKy6nxkMe6EM4NG+yvA7fnZ7O9/zbwGIQ9gnX9/nO6LnjC+gnoMO8Su
kNkfXesWc0YipsvKAg6hQEVKCGPxhaoBrBeHrttf6EHOiO/ZnAghQLQ9kc1km/um
fGtcz7HiTll996NI/yPp+2Zgs9KqluETe/BmH0/AOG1v/WlJHs1BgFFy47yYIh/K
3B4kwJU7om+XCudqTHfEzqh23i22IuqScijmlkPazboJ/QgqfrfSeHVVWUGboT7T
TZi1aHFZ60x1dcSSBxlga+dvoUdgFpauI+xVcLt7/JxvFKFl73ncVbG8MAoSKWnk
+zH8p69Zi3xawU59UuHYAwqdVEfNOkcPkpY8IHrkus8HdrYULfvwEpK8ynwR20XO
Buz4aarz1AimBUZgUkMXoWccU803xV1mfxumyMSVkSgKtVEpep02JMXdVQ0BK2LD
ZAJkfT6k4jMNbLiMjtzzK2leArbp9dZLufOj/bcQZ8CzIdfE4JKZLDVvAWBCTiRx
kyhaQDybWwPFQFcsAF0JLrE7oweqjUFfDJrC6DnxKYtCUen2HD785FRZ7FPkwAvq
q6lDNGI292EAYvwvKk4VsBT/L/0qN5pDCdzUp1xPSF9uLEjlrDF9pNDS/u6hf3ZE
yN+8yZxQBB1olhB87L8GV+5f10sIZ32SRnpQpaziHboZyBAvrVRC0cLVUDdFFUrB
6pm8tGP9FLrz8TWVQ5+WJUA39k06E6/nOx56dB4QVycoyl61ozkw5asfxxss6XWE
2UCv4VWUrLJrS/qW8fJeYjoSRBSBNfS6lyEYQypKFjMeVRY/yr1n+kbibG9w4X/y
iX/j5eaDmLUooEW7Z5WYsE4jevdXlflJGHQlH+/ap6ON34WjZvGIZqHNnKwVY4x/
flHkEcX0IcalFqw/jcP84eVAWZaq+w8/HhzQmrkWrVGuvXTWC6zZJB7ktiD8RDpq
60niFBr1So81EeezZsQTjnb9v+CCT0K36pmw7LqJxd5vm98I+/a85uYuREoRLch7
Mzbryf8x/yQvzQ4byJ0uMOKlv7GdTICvYcym8Q6jzW0k7mFHALdmTJIBy594JYmO
yTQIey1/WoQv6sV94AeX48rIt6GQUobUgCg/96oTYitOMHcOnBdoDE5rJOCgiSTY
/MOfFlNM41BzoACiZg58Vqn+7WyuFx7o9WHa8eP8gjDGRznEh4D99ht9DM9Jm+lj
EEG8+HYCQq479t9aqyT6eJud00Sz0uIbfXAeKU8HqQM/pw0AKnXdNXEWCDibdBrS
I3p8hdG99x4EfrYKKHv8ZjAOMdaw79bdovkvb3Aoo7/L4mRG3kVLL98QCobVvhXj
UMwC/U43oPmifBYAoEohZH4J2a2MEspsER34VdiKEfET/1S/udEnpDJkrfG8c9xZ
MsM8KFvea6Y05trLwFJtrI3Za2XCbBEVV0IZp5p8mxnx9opdt+yIxEOW/UFS61jw
qJTzlvGmAM1PMPQzObvp3NsDQxTRe26x7jd0uljbOMapeGxdbezmQws2TQhdB82h
gEEO9C1LniEDKOwWYicS7eTPYvg1oma+YRNiFQJQULxouu4CyxJJ/+W9v1/2N2Y+
7VI/5L4HC9/eQ1GTz0Ol/m3EKG6WOyQILG9YqQiyxiBBcwNP5KCw7GYnn9H5ao/w
PjAWxhLbkvsEiYPW0BV7lw7FlzhBCPAmRkyfv1pypfDj5tDfjPskceotMKi/6lct
xsW4oQ6MXWB7zCU1j/Puz+1Kt0NjUa278cw5mgif+uID7uuUSteVEcG+dqPqhcKN
VR8qnYg1BPJBiQ7157mC1bpBW3nc1uHok7Nch0aTPbuwYPXjxJAqBEWpu4Ti9k+R
E4XYDthhpg8bG0sV+yAtwMcRIMbFdXU/02eESAusDqQFrO9IbsTANzfIAR4Z8Hb1
NboM+g6ldqP8UOV9c6ZNS5v8mkAX0TNI8aUT9HNklXl917DIiDP0LwtKQ65iTaqV
QCncOjK1dDRrLv4X9W7veyTn3iD8oWwMY17VIWJorF0FqUlC8R8/G719jXqpwj9r
tWogr5c6Q+cfWgZI53rE20goZYAxu6q3YcE9fjR+Ws+iIQEcL2R6jAUPXKzI+uv+
oxbeybrYIslw4iL9jdflUJbApRzIZkYx6pJodllaQe316FbpTJOQpjovNDcfuC7K
UWVJuH0+LnX7ulvgR2oAOhCUYlsKxPLyUDrihlvxklSO3Sbi+Sqcw5C20zawLIS6
JGOQiHD/j2IA4xPcdPipTHvCEJyLZLkEKTBAQP1XMEKwuF7Z31yltlAIrwXR6fGa
mdln4MyVZZUwajGCOjZy1Wdc8UysKg+jwS+qtGO9Ppm1knz7oDKi8SVk/Y9B2bxA
pHh9rynaAiL2N5GdmrigXt6HCHdeXpLC8xYMMA4RyC3SxwYM6BU/r0dt2LLkh2pP
KI2eSc4OU5GBqW1l22gIo44+gJK5ya+uu1eEsdeuiiOBUKDjQaexXuEXWEU6AHiN
Lf4cJILBBBXLHHmz0eFV2RCBVGJZye1budp0csuxLIPd4Bv7e4ki3nS367jHlwxK
WKeZUG4B01Ovy0Y48kNUyps+Hcf891QIkPeNg/nDw639b41oXKjIajWnLjGdoahy
qfa8mC25WzQbyfAV+AGwZMQ6w3lIpFitzlTgQ3kuAyPa8WF2mSxLBZp6c4gnSRhs
iBeTByFeZ/8X886ZWTHUNBneNfjPSotHGkNcgEkr5W6ytg33Gd0Gmsd97JoWMahr
sNUBVPFn7OeIYn5kl+JFFrVQLxeYVyb0YUU2E8qFIBqBgIPswIv5fI2Q/btWViXy
L2SWHf33qCRbYTPgA0OXC0zCH7OUrA5SwAO/S+uZRsEmkwFuMwBXSj4UpTsab6v8
EWFFIvseuS83lvgYS2sRUTNC5PjC9Pb5YPmuYsQpy16vvM3YTaOfmr0eqQiAKcnm
vnYrKbhg3pbqH53BZGFO4qmQJPehKh4qIcuBIBgQCfpYkuTrlq5fw1s3Zv62TfOB
mFQHsszhovUlx3/YyqzVSn4DxRXbofIMUOR6SeT576WHXH2+NZCQIbddzbBOR/x+
llFv6+mXjkkwnrtEUGKQAYj0NU3R/PwDVmoPaLVr12U1Rfv87qDIjT99cm2kYh2r
OTwPb5tXjeYeP1ED5dsS9opBdhN+kxbRE3qtx9JGBfDaIU2fc7zICkdfTodBg8/A
raI2MI3nTPYUiUu9ZySXOjxOvkmYKB9i9XblmQblGEVRTuKjmKjJf4Vkqsl/3SY6
EVu+sa6eWJpGygsrb0av5GiJ4a/+KvGvAQd+CmFNVRXXHp1D3zhj78SaQ2DDmraS
F/Q4eWt1YCgudNTUhIOwlJreVITAo6UVEjX8iHNToAThs2EhpCFcsRnr7q9/RG3l
9kO0tpFKvd0fZ0woDUEBJyxrTDR1wytKIES8g6fZXCmR00gF4G8XR+rVkQV7+m1G
4Q7lr/GlONPfSFGX7LsV7acfrt+2MJsk81jU3qE2aFUOFNVlZR6X2uicyAtzAJLN
z6LqOtCmhiezVkjU5rechJx2ZpNClTbJ+0B5pgHIxc4M/G3fdP99NDHKv3sCY4+t
CvqME5Lv3tXF6PDSMPkGLR95mUqe6MPm6J5JhKN8GBRthkIOUKrOW7OSewDweRQY
8HtaNWlCkaAhKnIu6bad8sXEL0Bj9zhv0wj2mYRfFdYdkj4N9MqQRuW8S7k5MzAP
RwprzHD7YXEoinHnDislJBU1QkSOtg73igks6ygFXgroc60hUIbcSABlT39elRSy
X0PO61L+pkpByMrF0QIsSTVZQApHoDlKtg71UKyQvGb7Z1Y0FAVIX3U8HghAE+dd
tLDizV9pMlQCh9Z5Pz6/D1y6VWlOr2T69oZbvxx+jOsB8rIH+1AJJ73LULG9mYEq
evK4GEIDYQ6S2HtUOhSKP+3R9zZ3flDkkWz6eG0j3AThCa2RciIoOvoF5e1ruiT8
wpGMjmIj+Y5sbdJMdcarSlwp9qbnvV/Lyj1Rtismhb3xGul5JMKTJ8O1YRf6ug2d
IYQYPFAng8LsURAM+ptRgjq94+Oj+AhgU+Uc082jgULXhxUmbl+6z9i650XmwwKT
U3tjhB+YCiE0JeqxRsjnkKEgVqM8uH3Hg29q4W1cihZCFtXN+JuguRnAtLLbzyzQ
o7oX7sfqrK/RCxXNeTMEIUmx7ejdqyRejbexLd3hL6tis4ZVyb77HKHG6yYvjbMo
5LJ7Zopp8bSPkDmal/FJz1xOD2u5vrpd5xVrq8WhpS/x8bjsInol2ouC9q+xdQzh
AVYeWo3Sd8PDCbN+lb5j3JzRPPfBErxoBBEbRFbW4lBogXmmSHyn/qQRUijiGrzJ
WLAiXvluW4l9NCayP1OpPKfl1oY6nrXmxZUMyOBfZmYi4aVD+p/0uRRLtQhHTtlp
YGdg9fdzcfofgEB4NGgEtJOX3w2DbxtfWS4bBFUS/yLHvPtmld1L+U7ckYAXaL54
rF9UqX6hjiY4lz/ALZhazf6yPFAGCpqun0P4IiQE4k8bmZhdDvGsP0MwTj3HBq7q
5UMTeycCP1pPxUC9NADIb3FSuA6cfcQlZbeg+MaEKFwUtozmglq0o9UJDcphMk0t
nlSsFTnX0uoHSX3rZ3js9lvkXkNmrrzBjG6Kyz3dxgxhGSinusggV4Iu9eVaCbe5
m7ZPtOt1PLxmdW8EIfGQwAgySRU5x8R43UoYtBOPUp8S2p75iXLVQ904+r9SSwlJ
3C1JrbzSRVr0oxdR7lA/ikZUanR7rGh42b5vZb0S/kQiLeAKFPTOkgOSGevu1KLw
21+T7TfG9Jzrq1kr+EO+UT2bdgEFgqBgQWY+vGkQqCXui5kDVG00q7GKJ9gDVHQ7
edCQnZQWTlqeWcb8y2EysIbLcfX5Zqn/k+dWJr+4PoB9v9HiGRpyZRRGxE5bp3vK
oIq9JhqFG7cfFJXXrUII0uQ9V6plbDohifiBMowb+XMXAoLKLvKxx+FE/1S4csAD
3NCdu/flcM5oD5cFqdV5rU6w4ijpT0z9ty1jlxBhxEg=
`protect END_PROTECTED
