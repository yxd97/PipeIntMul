`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sOl3pVZCdFtyxw8cqjHAXS2CqItrUbT2B0ClGFbKYVyMHWE2rt2phLcMhge0Zt4N
SavYRXF5Gt3E4qZ0dCopL/4VVj+LKydjfz1nC1zaIy0gzp+bu9objeWpgDUWL3ws
XZRPj50tyw42Fe2NgUta2Xv07HclCYiDaMKkM5o5bzyyhV9pdJVm+a118OazO4Ra
/0jkD4acV2f0VrqF8E4DfLbvlqXUcFSVKdE2SIz82JnVGreVvvs2TZ5b3Eq3m3xV
ovWMm7t1XzvYdB/NoGB9bw==
`protect END_PROTECTED
