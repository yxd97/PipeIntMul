`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QZ/PqHH2daH+Gc8XeVprnutFDsSflHhtwg2x7LIlZ+NYNlifSXM7frNJS2NghvA7
jh1LuXnkaOGoelokXVRhY6FvS/e3eiXkeEbkb+MjQduRkzjDl+IMCFYDLo6uFOak
3eb6gnZv3R6FzwBjQN4f5PjKRpo88Pg9+UvcivzYeyEtAVmeAQnmWi22Se9EMJ2R
YZauGXiQ1N7Vl9yumgU2LA+83mKf2HVK3Kmhv8jEFYq3mV9/WNgWRf9kDQxmX2Xa
0TXg6nZ97G6MOowSHE4UWr7DYXvkfgV/35LxyOq1Og9ZrXjtZKvbzAMSKhJk342D
bK8BWFWFhm81KfERJFESIGUChsuHxt9ui+M6BYEy+lQzHV6FWIVvk65SGsjBnvm1
RPk0Yxy3AnPXaodW3t/+ImcKeTe8dYPjm3/XhBmw/WQNT/v2liu+7eq5pdB7S05A
1XWzOwm0m6SqPb6S2z7fAHHkcVvSbtpRZOYlmFCv2l08xEo91M5NOiSUOJCByHzq
pNvJJ3vPoVFFizVHYVcc7jFSeNkuvsiVd62U+fLnGtASUI4rSfGkOD83p7HcUUqO
`protect END_PROTECTED
