`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0LHwr6lO4XPeCCZMJi52jP7OmEuVitfHrj7ZV4iXvhn8Sp/1GCr9SHLxCvHOX2e2
66HTEVBBOKRtbgAf2KRGjCZPo6EgfcM59qbuAEWQoeflLIWNmEFU+eJTnstZiesq
pgmmLTNpxrtXvHRE8YZoQlNYbZW9RaBBQxDHVsFazZjkelw1uZbyjT4meuAuL02x
Yg0u/lA4K3oqwlltiiG/Sc1Q+SWeR/ECrLzXMIigxD3MK7Tspk8YGvkTUC31QGvO
gFyuEubeMZlf6MSq+J/rrv+6R2mZjFB6T5yRr5elAVLo4XtfMIrKm/YgXqw8Sq0i
ySW6JC0P6gex4qsBwPztZrBNNYhHxY2c/3vfWHfKBcfCy+She5nBOONPOpUYoxxm
smiBm43I6Vav6Dt6jeQwklu3GH4IkRc/UycjYSHoeUV2lU0nY+ux6ZAP61OenE9W
GPePxv2CZfP5fUQsrAVo1JP8J9Kz3LXqlAMalkHOCF2LNPmcN8nBSG8527SB2R62
QkTnZa0TE1jpnOsuECLu15BKewcS2qYBJpLMfgKSKK1JVqY1r/JHIei+lsoYf2UH
bvgpFuYx3iMSi/adj37anQYGrdojDdJY7fRPLrwhde7Y0+jl38MKix54HZvAKTTh
h6WlCSdQ938rAk62rHnmmjmyD5YFSGB+4Rw4YMBofWciV43w8dIVSsxQe1MEG1A5
ZyUjfo896dVP8GqtwO+0MzJi2p+4fsfYxHXeI/1Ww9xWvxEQONCidSUtQA/L814C
oSPUWznykqp7iHnB3qTEH1JS1fm1u2lSpnjWHG+V0idHPxQQ/Lt2u0q/RDJZWlpK
Nfx2iayLZytLScB9jLZ2jL4PltQ/traOS9rEFqGHx0cGMD3Yl0dQhocEmntbjApE
CkGlh86AftCt+vDdSTDd8yb3TSnAtmqmHQ6EBp2QFpll1t83VnCiKU7vD2LvokG/
RJqanNr096Aw6xG3QMgYi9jeItH1cudTGpDWswD1sAnl2fVM4UnYYA1UJUdLHAth
PveQim3HCyX5ZT4nwYyYczhVtjbRAri5o+XH5+CRHik36ukY4TRkUdUkMTzzb5/o
qXd9nTrtncljigIXJUM/3rzHUvRpNYGyvOk38vpBCLa5fLdwyZcq81VK4xzyBuAL
hM2RQOibmuQqrJuJKH+bowIQ876n6Z+/y9UjtKaBX/bShDTbOLNS8gGOvX6nu322
sByyFFD51tNEOox4fsIsQVudso+HSCodt+9krZdpXi0rz8cIW79hwSpPGh+2q5s7
VnF/fZL0/XR2BNsTJf1K4uAij//Ygg3Ht2A9yOSTw+obh9+0V4dUyi4r+MWRtlTB
DY01UHO8gzxMaceNKvhQPWACm7WmwF+HBDQSAjVcoSRAUcQZGUfZd5U3zk/HYGsZ
kPjlr0jd4AHJwEV4fWZu+YWyhFTeqZLkXBDZ+CJJ3KJ+6+AJnOZr9EmXPVQksA/0
HXYV54TBAsJiVZ7x7p0D4ub+gLPz9hvqOgzcU8i9XjU2Jd6gmgqpS64ODpjs/pow
MCV13En11IWR2u4WGAzGPsnNkhcms12Zs9Q4ZxbS1Xf74TvCbgbaVsB+PwZlSatm
8jY+Q7LHpScahdt3LH4M6+dO6LtS6Hkm8f14hYts0OeQpIapnUmCkwB0iclZTzKy
TUYOKt1XcM8rg97IMBqd6ybHtrfoFtvlD51xSh2k57EBp5xtADEtRzGrBLVdnjpc
Znsbk5Vrl+GqpkoBdrmd4y56weBb+JZEuEM1Fj5cWfWz09QBEWc3LMVF+H2xfypd
bF+DfTrElytakuPlmrQBzs6P5UWydm7F9z5dAfD7QydrCRES7/caqdiwdDbP14AG
xxohisOTaJE7sTa3c/egSw/7md2ZxkdOEZCgz9MRFFnKtahcBEXzKOvOyl+psC+/
aqSfv3ZeDMPTTAd60iOwgHm0qLrXMICP937UraHGzvMW9zkchmwdZYCJ43SPG+ZN
Qwg2WfQCcoqBvxm4axIJ0MxoVAqxT417q62T1AuJj16nz6s8lY0PS7HSeWUwGDeD
kPNjyxvZcgRZggOY0gPEap+SbHRF4Jv6qe8WmEykbgrQ7oyK2Rs/af5gZ7AUhNnw
S7gqDHy8+15QiDBw5Cs13aNMNl/Vvhhy4NnEtnwygFgpCkYlX22z83PAoLwf8xTU
fC4apNqnfv2xKJTtPRUw4y7vvi1RQN0wCaQkolc96eFBSnOxCn4//bw0t4qQQQ3i
ftHuil63bg52DBAnUolZg3/jGele1BwkAwVMze6E6amBCE2Z77kTXngckLTQTEU3
uqdSEYq0zEpZjBOrjeMA7bDdlCUvsXP93Rk2ETTXwfIY6SRTPA/GzK6c+CvTDu/u
4beRd4qjvkEQW7U0iMx6xVPFNuKM5kkAorotHaPKAJa4M8DL+sOwSFuVnw/vIELq
qOzSXiy+l/JbhCZyU/eTBtB4uTwtY5Qrq3axZ3Uupv03ZVT7eDBfOY2ad5pX0FSg
89NsApVzac9W4kbRRX4ycOQptoJL0qDTeczsxSdMdt9q42auC7Va0wyNwz0x6n7z
WZFSBZcFyqWvL+2mWPbQttuDURtKDNviTRP45sjP7G5xElmeSOQmgrAmHa+SKIbi
s1eVhUO2nInwGG2hJy4pX9Ua1zqbKpqAkbN8RfNYhE/2kcNahjxii3kCnJx/Wu2k
exRTyeebst8h1YDK6MeYdM/E+PDJjHZjiKwUoC4tKWS+vTKDfSNMS/Dpwb9E6Yma
i4dtdg6q4NcWAEsHMeir4Jes3xNn99DRAUUoZyg1cugk3KGKG2rxQCtcmk9o6auG
5PoQ8eOzZqfDK/batpdRyg==
`protect END_PROTECTED
