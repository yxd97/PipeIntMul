`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
365uH6rH7m12BwxCBHdYsq1BuB4ABWVLQ+Dvxw4SD1hGQY8H5pnq8pU/ei60GTRR
G5wAvlc1BtwScKg2GnNKowD1xJAYGJiRvI4o6eCCvpfsqIk79bE8KndAiK42c6qy
RDm42sDgSnQXiLYxAj2DhO0dePgj7y5CLdEcPVpydk0Odyip3+fNyWEK+z6Fz1As
/rV0cqNakYFIyFDY6C+2ba6bv2sD4bPgA4lwIqJRDUgODUGxumfpy/Akb0Q4ZoEL
Lx6CCKX6xsupaXRGJyK8Dk8392zPrgzXjAecDZe483NNg78H9XVM9dhh967UIJOb
lNMSAKaVrbj5XWbtIGbhhx8FUtIcVCcRzKZqrY1iievYw81zH87A4JWnL01b4asV
blCgoVXkXO65qEBn5F3oT22xSavqhP//cE6YKBmf+a9hbGjR3sjb/j22bDK1ECL4
b0aQd1RN90Cnq5zgWakk23tvuUy64aMQTjr9LU/57T2I81KItwA7PY+feFPKVbQr
C8XF8U6Dw8IEGtBursb4SYeeN+wCX7Rpr+tqZ/cOD+fCjt/LStXgEBet3R9/+hn2
sRSLgmWb6RUPop3Aq3xDSsvWX4vvk/qeCk6q+p8+MzaFOivqMkz5OULGxavN0PAl
vLS89hu4y+XeD9gnf8dNvARoz5R9Vz7L71a0WnrZWieGtspRo9vJv9J8RPw36okk
UrFmu0ty3qJAX5ylQjBKYggElLqwKYd23RuqsCt5/f+xSqFlZGQvULv0quOHVl3P
0Qu+7/HxkgQvPL5Foy8y5LP7eJm/4bsIyowGsHWIHWTw+8MeNinqRXE14KNf+TpA
AS9TVyXk1kL4keP8UzIvBRjMLW5pfvBgLbQ4y0hAfYZNRDpP8rZIzQi69dPbK59t
AnreDGrLlSepy1UjhMix6r3EdR55EeIwsElppSjtp+95hPrvewfF50eXNd7yaXd9
`protect END_PROTECTED
