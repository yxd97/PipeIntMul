`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyTnGWb4mIAPazMRkHFDk2xISXeDTXDzDrqui77UrBvwRjkgaMjTLfQt84PKwRXH
zBf8wrDedu9ZzLWPL83jgix2lAVn6ftzlOpiNc7Wd//oHUuoiDmGXoodgClUmqJ+
DtwZ95JB/civy60DUbomBzNexix1ZBqAVxyR3TregHOxAfsSnWCfREk3w/3Y/wRK
5apW7vONuIqOuftjmqi8gQe+sGg9G2G/kMNAhNSfagrrIeOQK81oiVv9+qVGdcr/
LNlAt5syp+4KfjvQUQdGUInfhAxP3dR61jpYq2PP4rUE/wXFm/eCOxLeqyrcvP2d
ymF/EKTEhuvIA/HNa7k9vhp2ttywLSYYV1gP1nEX5ThaIFe7u1Xw4fTOl0OTlJUa
xtGU2zY6cZWMHmaJZS+IPK9Gyl6zinpKpSwozuExPXoRiVkAs6Usv8HjoHKgySsR
x0WOQjWerA36H5KVYNJIurZAEDKKgpes1Mi/WYDGY7Q=
`protect END_PROTECTED
