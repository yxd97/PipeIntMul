`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xaGXC64Bxu6ulVy54XhHNT4DfC4BzWMzIffbq0jYhUDW5CGrKbt0bDGavTdMlqfx
amEQQ7vEegpkZS5BQjDiXmo1VXiPGXqvdA06rKUzpLJ+hY7kJgYGUWbI+KHt/R1j
GVmmg5v+yqh050mcf0H373IZFTBf+TRni5Eq4+5RRCoGmAnWmPhe6k1QrcGEALsh
XsolBl4SN3QgmEwQoYpNsASOAcA9gghWmixigytLJdBPcqZfpJgIsnGmsiVlckpC
TwQM6RC/j7wbaS5YBFlDKspubwPcpsz8PxtuVBHtr2udUXZ6X4jWdbVZZRmLFpQZ
okEzYwkLO/js6IG8uBvTJiSDkcu3Nfy9oI2xKtmWVtqgX9KGCdsI0iEbtWMURsi4
PVRakDpZT3rdIlTJ+20KKG0MW13+1MCz2Kd7UJTxe7T9szb2M+sibqAvG6lcKXk1
IyWeRlIiGJ5GBQeg+DVd1+o/p6eJniefXJoTwX2bLm6KD1mMPRR9VjB4Aj/c/BQ0
iiu56DijmYDWHAkftBvP0LUodXFozV3IMsCxfVr4MXJCikE7J4IdScZTKASykh7U
j5/frVGGR62UUmOUHTxy95Ei7Fms0tchfU+mBW5Olt8XD14EDQYtp9dXez6K1TyP
`protect END_PROTECTED
