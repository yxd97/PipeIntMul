`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EGzNg6QdsXDscuNwav3I5qWGe5qmWHEZ3TAEHJoDYLanzz+rYN99BGdTBCN7aYZ4
rSMD0j+Gbdjq+wbdkk1Yc18hcOrERaWfO1UcjWZWwHoteuqQQ/esZHgbNecsMTGU
5yX8Gb4rWyNwc8K00w0wZRO4eukATRuFso5pWrKoH/AQeuKaIrgDoQUEGdqh2gaT
AjwSt/Gp0yt8JgN73qLborIWkUS+wTL8tAU07pz/R/SnhKrMzXVzdueYCYQ7WeiV
NLlGHkUGYuiVr/tXPcFbRHprcUiIuTknpEvpynOEeOV8C/ely0lDo9S7c5hY/B8T
4OsscGLkcM7+cRXU815IU6l/ykA7H7U6kpmboEIl3QHUTKPRVr2Y68r8Z5kV/5ng
6jPrWMMxafl1pCGJwY49iykZQnvZ9I8ofX4ITFiWntm1F8FEW2NBpgvILLOxEvT+
FCDNw5+iNDQGOMTwI+wpT5xX+D8XV94nCGBZ5ZWTY8zVCuDyNDgejlLMKtnQcyCa
Cfe9M+8VYScTmGu3l4XZBAdNkY7MI5XguVFE5nOqLsEV+VYjjL3IYIo9SxreO2k/
`protect END_PROTECTED
