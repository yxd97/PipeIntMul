`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fqlow8l6ZKz+iUKTfduM4HmLm2quIsaiGo8wYPhuGyW9mFORARIQKxMqJdVUDWqQ
CJmiGnq8d73ZOJi1n6hATEgAzWMK4SmnuYBY2EK84Yg0BwaEY/lYhlATzJZIZWEa
roTPkbL5byXjX6zeaoFqbpT9ENo9hK39V3kGbRDG6FTScvoYYBZAo0RpR3A2c98g
9xagzaJgmg8I4EXpjNyqd9yQOuTVDi0oxE6FRZHIZNbZ/CZ5MoKMYBRweg1QY6KB
PnkbEMQSLom8ysi8uZkduPlohSLXS5UicJS4u9IWH5zrSEUEDZUMnANv1lbCU5Sz
yy6ZS9aVMnuonBVgmt+S2rqf2d9/cKeJ11TRrjmNKILr84NefOGh1BE/9MTYSl22
M3QMVzYK2SIHOv67Xlfc+Rcf8SNg1vKEopr9SnYsbAqqvCSjE3TvozpsBT66H5Ak
52RsJMIt6M+i4pK83YbIuZqXM/hBLi1/uIj1Eg93sVOMjswRvjixfYIDrplMUHcJ
E/HG4VioehBQ3fzNZay9U76g1CtJXrJ/jgJZpYhnDOud9CMWZO34eT7/YzHpGQc3
hfP/81hjE4qaY4AbdX8Di8GKiuyelWhFFyaU4FUbWV1E2JRr26aYxWwPsSssH9Cm
trdj9H634lm2D4/Ky4W5tLlANqS7WUgI6WTX2B1QLaKZlEeQhAU2sJneVGd5T25U
QlZXQv/6qpNMovNdZLPHNHfQYrQ3gJw2NbTYAucTY6yV9NsaEMxWFW45geOEBaO3
7QtnT+UBTi0Zg7yLgMDI8Sflyr2pMHJ8C4o/sx7vuNfgZ79ETnqx9MNxpgo9ZrYr
ZXvoaY/MszYLUQ3zKGG71S+P54EKZwgQDXhT7XveUq+mUS2Tk59xPGsERzVYFPAz
CcH45Fi87ZLDoTd3siRt2zRr4MmUfOJzlpD8t6gPug9jWOnhnKO8XYpiRTEi35s8
tEpSiG0IEsFAMNUXl0bYnviVI67gq2nfA8HR7lUCM2KL/6Qu6kO4EJM1KrLKdhRK
AW8mMcKHmyqSNb5khDGMLqCCtE1kGrft9v9+r16Bp1fHC4PjSl3owW5h5AqnpH9/
RdFdBYnQxmX9vMOqmbWPnzKD717spmGtNxFuypjdAHh9LXbrQUKEvixEFY5rz1e/
/qW8kFhOySJO/4YlMPWt09rDfkJiGEZJ08OT3fLgNkdsTehuJo1V2U05TJQdy3bY
zvTKo9bSYD35gJ80Vryh8wZSwXknuP7lJ8kmXleInAI2n4JN7F8FXxJ2cMJUsIoT
`protect END_PROTECTED
