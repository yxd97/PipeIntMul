`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lOwAnv1i6NGAdRYzwAfVklt4T8a2bmPFXt39AqyfMD4CrOhg/SPLWIaGrM0QpKN2
i6Ajgs33o+eiR4Iaq2V9nb+HmaI2n7eDQylYRnZ9u/OL9BSU6X4js/d+5BZ5VXr7
YcLA48CpGnxV4lkaMMTm2BaBAnOcT2OeU1sRJGqHDUQmY9Yh5OwiKzPLS2d4D8xq
Q0nFmrhLRzOTO3EcmA9tr3zCRxIEaWNgCGmNbcb2EEtV43gUgOZzLWUjeebSuLYT
xigK6fJXgaqc91zMRzQkh0kK7ApI8QKinS7/32WgNUJM+Ozk7Wb47TqkUt7Ai13S
9CblW4VUldsf+MZgb/M9KEf/J5N4ON84K9da1JSRIAbvkWZDFIm43UotjyD+Ed44
HfWojB228tQJHJJF8/mQQ6EsdYYphf0niSe7W+t8Lxb1OoqocS3io9znx8KuYETu
SyKKk0sdKwHnbQQCrOX7Yn6oQn+SoEBZniaL2Iw1D6RHeCuiIudQs0Cp9LhiuPWa
emmEMNycAP+ib4sF8S9G2CsZcUdZYBqp7QaBNLVpWgTPWFqvud4UbTzz/h0G95uG
rCDr2rVNdHkGXQ4Uwf0ivz7rLuZ/iRj5frYq9WoPUhyVgWdP84e3qs0g8UmZd5aT
xzQ99O8tw6VlmPreAECeHA==
`protect END_PROTECTED
