`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k3O7kcwFldSPwxZ3YwUNDMXz87gLlSswf+9UrELd+/SVrJ/Fu3iKjn3b+UMcNO1s
x5swRMvB38n6X2oPfR4+slH9cmWCsXP6+syVVKoqJZ6lt4pZyuYzRgwSsssJ6D38
P64R5a+xmzVJXxeTCllNwjHcArs2U/aZ37iYLT4/ITIcnZE6FGoAutwC1WsWBogj
tMBDmVAMwt1nTmkAF2wYGU75POUcBM7lPMlGz8eP7T05e9HwR+i0RfcxdV92sgNO
+bWc1lQed52C47QSfpxfku8ffioPQ7Viw4YY5t5g5idHhouaxnH1EFAV8bAfuZa/
jconcHy374kmjlHvy9KECY/l65HXZu6bVr2QGHuF48b/dL6JNMcBr6NbrEY1Litk
KaEBoZsaMF58XfCSxvdhoZr/VJImm4zkjptKsK9WXqMdR8CkX6rU+lhfA86OC3Yh
HBt0pB8C3zPe7u3o64qQcNUq248t7EulADO0vemfSdVODWQefaPJDBI0ihCLQaCU
sayxf0/0hUfIkSC1OTenLh7W978uE3uRP32UCdKMH1AgyfNuVh2Reuqake+LCcJf
2UL5gnzIz4tl8Gxl2Fc9wsuU8s8DfaLctBiwx3PfrSskeA7KXuJChDJVoO/YfNAR
Fa/zIFoAKRvxrA18J9QGeRY1s4PbSxTK790eMdPUn9ovjGXuAQ/8gJjadgjelL8B
ya3AkUYVvW8mgkOmLCAhNECfp6xlpjW4OrhVAFfgnXwcApNQz3tVRMmrsnODWceT
iVk0TSsjdj1qkP+oBKnFb+qtJRYG+JPPNBv016XoI/SB41z75ukdWc8Lh7rm7vk/
+JBC/FB5YbZz+4d3b2LSL92zfOAO6SoMh+2JNFERAbAvuCv3oeoHfGVMPR0OLTxu
rvm0mMR9voiAJuKA3Ae7dAK8vuQ+erOjgC9m9GhWQaDBU6IiTgWtZN2pHRigg5Jc
8o1ROZz6/W05OQwL8EvCu2uWO//I0RTBLEfPJXnfDgwJZQDhGnExVl5AasvmcNQg
0oRJBYgmdCOqes2O8MoYNbq7gOKrZe6Tds8CYUosG6LJ8qTytVsu944WT36wFgWG
sWXKBg+gpgYe11M/cHW6mmCYPFhpCQbFVa+fo8hd/C5q32HVtGcN6VaVzoAKrVDa
WzTl57MAqsCOlWk5AfE8GK5l8Rzj9Q76rgfT6aHZkWDRXPJQuS20tVZT73NUJCWB
s1R9ib0qhrJv5QhwtWl9SoVoePGyqy5ig1fieaX5aq+z78dyCU5RZRX3B0a5mxbY
FE6NqEXPkktcOxTQdVVVlvhVu892mpSsh9hZMt/IzOKG35p/5KuRDH6yZtSyIGLQ
2LWlhMroKrTY0tSdlMgJDlERy2IyIR7DM84BSKW5/sKIFbpopKNZsE+BTAcdzR+Y
AeDwcZSPo9URqRNtVukDToY8Hk9XWoh9aziSaGSxLa7klKbL8eWvSyBSleieUp2V
uHHtNQGPf1gcV4SvXwiNKzXXSuAxQefXsVAPPskIrBCkl3dRAUZplpALdqHWRPzR
VrHXto07dztw4Sf5NIn/3aF84CzcPZ/5gnNAvUzIssrsrA9PioeShIYZ7jtvtwu1
eZh33z7Ea0inHFGKHTkL7Ue/uAGg/d0t4XEgYRIlH1b02TthROdWKMw7M0sTo6bm
Kr88pl+RZLK7nXpe8m6mdFJXQDTshYQGPV5ZfOUk0IYa1WcmuEvlwY8lSZwZQzco
4yWPvqAfWax0LSxSWv08FjJQF090H40jSYoYPLQCJ+gm+/vGZ5PAWSVMWQggCTwe
R+jlNaxS0TS6kWyDj7347H20Qa5qfB6W1EHQI6nx3bXIhxMuplkz6tdj5QS1HvrY
pPk6rXmsV68LqDtOts0dxvARqa3eW4dv3cfCwxEMdqtpohCpLA+Nx6oThGt7fkp1
ebYN71iDbVJ/8VZTIk/tJeIMecN5R8Bu8wreNcQUULMFJKZRutB97gG3cwjcxqDY
sipzy8wnaJchtELCdE6Fu1nrcqpR1vH3jM00RrAh6XvzbE/hciWEbsRn0WDugS2b
8cz7JowxzNhGGkbsQ0taiPTrs5Pg0pnBJLiURek0FgjPwaiSqgYX+0absdyp9m1K
PvAiBogmscV+Oj9SOoDVufqBw3oZWsGmABP0yQ2coMiejhd72B3h1tuPoD0hl0WM
UH4UQ/KoSA8/XNWa/22Om1NUjZFubQs51HItOw5udpfTecavApV06nMnePtpoEVB
ro9cFmku51uadfsqbG2OC4+zy8J+smqClsaabubq1auz8Js1Q/PPg5EoWGxjS+iV
ebo/AhxISmvFb3UwMfZdOLkPPNGcmiqmwFwXTW8oc/2wCDQ6h2hzWmxENw0iq+pT
z/+n7rtQlsrt2BaXrYg0cJmM9PLKAtBjoqN8k49Es95wftWr7vqNiJ7N3DulaWKS
cTwAWfkSeFzv13LAW47xrqxCCSr9adlX7md1k0PXdCL5bcpWwM81ncwu9RXowDWQ
jWVQV/SsKhwgnThUtnERY/f2QdKDub5vuCT276fsrUND6H3rRlG68wFJ+PJYWRrp
SKN6eKLzTq+Js2s9MGFGDZHBLRimXox0CDfq9YknozTGNJq+zRPz1o0SUz4lNU1q
d7+vTzuR6MA4Pn6F/9jz6UFKfKJT3LYnpzCWNkJ0EsNQf9aiWvGq/mGOHaAF9J7g
kI6FdbGsYeHiq8OQKqVsJkQsTkmy6gwCxXAi1UOkRXhNyy8SGiL6x5CCKpNODX1N
m4yt7CpE7pvryRlCaJIYMLc0w/ibM2FlO2uffmYwGFCfwRkU6Njz4kRA6xt4xAwn
0Kjo2lhA+oYQJVyoLPlB/G8BOoGTmgxHm5DLLvKl0d74LbAW2jqqsWLFf809R/l7
JuMzhU09m3e8byUiuM24qanDza4S1DBY5Jrh4I5SnhmnSxnAwtw4Nq2ND4MGsk9T
T/D7AteL+0KSwPq2PUokJSdC/fM9pRuOatlUvJHgEzkx6P8+58Zt3Lg5K880ezjy
Xvk89uoymMp2HwH+/yT0mJVGyTOKk6Op58hyiC45a1slSmKFivgHAii8d45NscK2
zc2ydTI5eNTqemUe9p5NpCTga9VSbOY0JGQ7IYePcqSIucEROZDhCt6psaArQAYT
s6oeYgb8Fo7CQEb7MBVgIMNgxPl4Xy9fn+Qu+NrbNaY+Y4Gj1NQjqkMIuOJmuOCg
2qFCakKSYdO9nL/+M90/i/v6BM6fMuH2a8oIaR1CWgZYsCwM8YvGPXrH0g4E0902
jhGsPd9ZQKOj1DZwaXT86BgnQV9wH7eNaFGkBBqm0pdC+o5uUzjE3lre7h98q97t
4X+jNtj4IzWv/VqyfLlqBkrAASgLUQlowEwML5RKehaoArelFri4cZRZ+EbDFTb0
Kv0AGyE8qslESa8WAd6enXXvWqlehtdA8m423g0oNZJvDDFPAxINM75NxmFyDaF9
8+x2uP3jvjXCpNIPJMhjCKmev6cQg6dajw+qpTQKNHDgNGAwU1KTnw0ZPDZ2m68Z
XOPoe4zvUmrHA8ELBcmJwF0Gr2XsgXTExaiZs0JEysEFS5Z2lH3gOMnUBQqoGhjY
keAYMrt4UmnfX08nzQuKcoCm5Nse2GkedBs/azBeKY2o2Pw0+yELl7A4c5UzOwU4
+3Sor8dqxyeO8kFMIk8MC9RPuBVFWgK2vFcFtFkPOLodP2krxDUQc+0zTX5NXL0v
sooeY2mUxDdZe0KLr3mega2G+VQZ3P4BaJICpxZoOV11/zqdiGWO3Vh5yBqFrsDK
LRWkJm7AdICOmPbhAovm1HCz17dSjRvuCaoz7MBcOgVStr7kUipt2VnM40e7cYmf
Kt6g+1RLvLViQyJbqXvk3xv2Fjt6wgrg9/NtiCbgID/BCBzmhZXZQSWWuWpUEHf4
vzCHKNxCGqlRlM+swU6N6js3lhZsJDnCp6OsMfDWK8pFpZ8ufVTkximVGPtrpGav
dCRYkHKyZdflj5JbBaImEEnZqnZ+cpDNJUGw45L5SAtN1xyIgpDK4rAa0sKClaFe
vj4KTBKIy5jHLHjiA5tHqo0hkSRmFZJe2Y11iQBPnPF3zcX126DA3U2/r0wyKw1J
vk2TNwhj3Rf8TKJAsH20RdcnhCv/KAsd4Fc+3n4GdiP5/ifFSEJUH5cLSwT3IhHk
UrRfquVhhmXMvRKR2pjm7gQeGDmYjqXSqA9MJtDA1HJzt9VaGjzjHnFUOZOdhU6p
i5wb5o1kZafTaBteMnv4pXnYCRwAQ3vwjrR12+T9uvfkC9PBiW8hbPIQPnnU/jtn
B0hsVXAC3/YOJJXyQ+BCoP2IIM+B6ifs4TPKh1BiwYb3159eMUYR3yxA57bA1u27
MUA4XRDZd8uz+7Y+F24jkWVpVTfEUedYrXU3nWcpFSTln8WL/JsK1xJvfu0wFAft
OBozGvKE8fxWIa/b/6R6eKAH/9eHSQvPtX9HrFbslt9In6NTS1qT4dyOrJR1dFQE
Wag7/dwZKkXQCBm3SQRMOs72yZMnczzv17pMkS0z8Rm8prJPf8zk2arnqXi/4HVo
qeSKgyhj+gJGntIBCxIz5zZrtSyYPIlGtMu1Tt5I9uTA36uoNCRDrTcw/OJ2r0ij
RX8o65nODOsnVe9M27b1+nD9qtEBKmJTo0U3KSVqPzgV+V/4mSU7TDxy1YI0Q41I
5cHVHtKFIImM8jFMUPW2bSIjaDqZp7HvT5XDw+Y3JTOMEwZNLIorhZj03PljWa3d
QCYUT0X8emmeRC3YGpdRi16ArhM7b/IuBJZd6905FaJvthbDglYoqWz10+HGXEgq
HJDAKxAzCW/OAyXSJJN2/Dum/41wB+W9V7JcumcM/o76PdvceedUKCSOdvNsMSIR
TPaEHA1WV6D12WLPzKM2fDjgTeiRaGrg40f+qKUTtYU5Jn8u5xBGyE2SUy8Znblj
tJe9dez16ALkC0ty2UVzx0OhkmkzQEE1AwrWOidu7muPlxn0bxVO1yFeCyh8qBbd
MUn5uZP6wT6OWF2L3LjYmXDq40gdzIxqfg6i+QR+AppTHp+B4g36xhA/4e35oT0q
F3WRXUg6iZhZGQdoupKqvooNhm4zd+Hl+PSlU8AdbBYkraIQbMtoYjrbQAhw/ou5
LMoMJJVconEXWFpXMTEtD2Sg+jujyWXkGODjkVIM+uJkkWYLN/qfU6S6lyM1ye22
FwRTDHrlxx9wix+pKayMCYScGipIOaVkTZsDsGEcPFj/o3aTwrgHFCfpySwUiYJ6
ZjTsQjgumd4ZY2kYD6CEGTK0x/7ge8bHAkTlJx6g09SRT6wKqXofPq1nGF1zIyXY
7mFuD7XVfjAFQ8DEXVvQdWEQN2Cdy0Ss03S6FmoilmJujH1n68cZTDjO8ONll8TV
xnQ4+XU8oZvsxFdINnQ7sQ/L76tKsROkSustB3/jcwetE3LiQ5Q8dA9AifRnKuvX
p2DRGG2yUpOwpHtOwVvRHkJxGugN2U1q16HuW0l7sz4XHNpnOOkFmkwzA9oYUd/B
F/B6GupK31ZEvV5XJqgfbEfZEiNZrFbWrR69KaZilb1M9QbWVgI/a0hmfEz3xTFO
B0znwz1BVkpFp7Z6jD2FaePwRrgfqhI1CwHVTPjViocNk8kSFXFcAWI4giq3mpH4
H6ji9PlKo0L0n6MGir9XqBO0/JrLUV31z8r6d5sETKVJDNdzaB9q7k+Od2ADli8D
3at6xq03InqxHb+WkBSBJ5B01MtEJOLDI9xoFzj6SVRWOoeLBsKN4pqa8xJ6piSR
i/CCN7SqVBibJ71ETVDawIRnUzZO2Ao6DYYhjVoTgG8ruGuj/FXspGOrEzYrZK6R
uaVUD/S46Oal470kGFg1NW/FxYyJPB9mGTfSr8UuiK7CQEuf6u4yC2Nctp8WPo/V
+dhPBfb/rTPkAriOHwbeFrsFc+TfLEuTeVXzzsLH8H7no2iUlQ0pGVxoKZOjbqWB
gTsKu1RJZWmDldkg6TRzQdtx1PWhz9e2ws2QzBwv5Q3IamFSOwezlRK9FowmqVBj
Mm0/iAjVv9SQnFIqZ5KD2n0zUM9u63hw0k8EbNm35uMxE1V0S9Uwz98/LKfuKEjQ
Rnq9h+1f55m/TcNXBg99LJpgRDHNoYw7POCFxsv9XWkc2TZHpoUrEqxt2qtbyrfg
Yj3nEVSmSCpPcHmh7W/3pyMYtWzaB6TLSxpdwXO2IMSp73kDL+a7LMx2h2L9w7oS
1j50JxA3fXhi8zYSFHdHJEdn/DjkNYD4RUZWBbkumeyvFJ/v18GzH5T+qEO/8C1e
tHYoVNT4qABAG8aFyWMRZtt3OclaEJIoSs23Lm5ZvLenVW2qAPIyGt1VB9lrJ11n
I1NUT4fIZRQpcrw9HlRFA4Di7dXayU1r3uRXNl0Pei3C9LURk1j9nsXrpgFlsrBG
3bEEmlqkeBm7A7k/xS2jtvfRvHEvpn+X2dzOOdoOxXmHT82m5OTI8T3Bfq55H7UQ
FI4EbUHhquD8cBYVoLVLnZ+mEV/iSQDb5G5/CiXE8G0Qp37apXOW/tCocNY5nXNY
H1zb+OD4oXmBHXrrRM0121nCiSSwfwzVaAwa9zgqCPXdcVl63a6pX3gi5NzdieNr
mMH7OJZ8CwfL8PWkszve1BNKTpaav/dQUbBA0HYBgWEYl7e+AXYv+7YSAzrIgLCj
UuNdyHjDQGA3Yu0g/82cPtSbTHSiKtRurQxLqnKU8w6qJi91jWkmGGFlJfuTVfWv
dNqlqFoc8cDu5L++FpiLN+2WvWfPtZ2uImqffWQFKwhG+0jK0aHnRFEAq4gkOzox
kAXvK3xk7U2pH0OTleYp4xo42Bz4iXtqsSRbooX8oDvWaaet4LBuO89wBb9kEOsX
8j+76ARBVYSIGX7sKWKOMgW5kIfUq99hHtU6fXycWuY48kzWQ9oppcKrR61oZOIP
AAqlHaFvQ+WuNxcnAnwKGjVXxGGp3J4+F4md4I+cwFaMwB8wjzE/IRwDoXp8FIS1
BqAyO39JZTu6r5nFV1OcEuR7ohIFwQd3+w6A6lufYkwJi8t2p6Y59ybhCAJikXQ1
d5q5iD1uYLvzJT3+qW7a38Lx6idag2ZBWn4RvBc0W5yTttOZowZMCcSOfSklf3Tf
lFeALgywpDmF3oqtMDhq+WsqFoka0j2DSR9Ikt/jyIaBJvEt+0hcop0trCjuTLAW
W0ivt9lU0ImscWNMp1xUztUGtnd2fDAMwF/lOKAuM8qUvWXqjB70+imIWDphWiB6
0TpjgFK0hTnVo8O5Dz2vuUoO4SvRy4KO6NeoOgQ1eG0aS2lQ+OAAesnCRw+hDRY0
LTOy2qC/+tT0h08657WgWa/smrdevJttKr2P8EP5NkO+1OiI5DWqzg9TFNDDLzuy
M0a9Ldim568794CxZnUqM/J6DS8vG/JeAJci6Z2WROgYcQ17+iI0UMvH+3ukpVr4
uZmy85kFFwTVktYKSvDQWLIEde8fRfwSGwNaNfhdI+Li4ytM8ljWbv6pi/W7hHqW
lLR/fkGrstHQVIGFoLQjD2X61fBKugG61EurK1KGp3WGNGMDOIDAOt8OeS/Fu2L2
W8wEabuaBFLxoMLh1BukC4uYVoa5QDh33MvNAf8NrA1uYMsMBpKdNV+DJwcb3r97
MYJ/2FW9S+OI8D5/DarPxoRdtWTi+WLRJITlOei9zC5VTBz9OCN8DPIYhVcI41lR
CoUbtCs31a2K3uhtgQ/A1M1dpSbF8kwln9/AsPeoRfT6oL6O2N/fjus4VYFzy8+j
AsTIZVfJ8gpiKnFOf1xQcKX+qZ9UzbpZdMElVgq8WHU8sAsxFifsTyQE2SPHzTap
lYymNmX6MaM9daKKs3Ar9xzdyws8mUfp1zMXnfeAXfR1wGmlC3ezIyAX5WRHK/t0
ey/Hd5FTZYKY1IQWfAjm4IOy49fIRgkVOdLty9K5rgTvz3lhnByEgUmMwUymmbz3
xBdb8qaqyxn1D9ZLIQjxA024ZYXV1qKYGlC5YQugR1DHQiauvSQ2q3txI7Cu6EK+
H5t+lR6kgqf69lWzgNXfOz/9q7BExUysp/MmhIbbH51GWtMA7BT/EEBXXmF7MfLR
dW8R695lKwft9xLLcz2QypeuFRpFUNCrjLlclfaJ7S3Syvz7/GulW2KTYvMDz23e
N+smQJij1qlJcoqhX9hJQi/itZtkXA3NnXM8iTWD9LqyjiJuvVyneQ0rd0LsoSOi
2axPnN4OWph1mlR77czL2pO1QxGEJrFfovFdo9UYUgW2Y4QcaRxB9bWSKXW531VI
h+/nCT05HZz5XHnDO4qXWTsvxw3GcKTdEoxF7YwW+CO1yRU4Tixw0gkS1CBNG8sk
Jgk3bSVNWnQarbvk4TvbBjZ1A1s4MLZV9jk+rdc4axTuTrnxRL8re+HN2DhzE/lb
XoVItVD/EUFS/ZYKKnlvh0dMYUvPYJHNu+vC2SXAQLznIvxlZ2pAX/WczQSaW8AO
wghhico+MHVsQ72tiCzdFVkHO+Q16q859ic/Fea9W04Oir3f7yBqS2crrYg7TDma
MIakthwAlAOKOFqiZwT8HyR+wGvYxyAuu+c+3xCuEGqdJlMD85fEY7aciEuH7l2H
FBzg/nkqTDF7YbWAWBRKN7d0FieXJXRtMRJg8bKXvYszR9coNhPXTybe8ngVrfyN
nBZmZXAnCu0Is0U2yZRnqjh38nwKTsYKZgfMeuAp6A3GOe+bD0B5qTY8S1bzO9h0
3bH1oBpvFSwUkCdzeETw6h2epv5dV3vGh9llXvgaTBKkrc/RIRPYv8JyNEqDSsLX
+RMPg/ceOq3+g1LD8jCNXthvVGgTOsWUi+8IYRMlXd5NenJGCTfJ5Q4y9TDTM1DD
Lv6saeOnaruSmL04jvj65Wk68a3XBlINhLiJHy+F36Sbp78bz8WfB5ImPXwoDWEw
XpgRBDwk9shrYQsDvY1pp+J1x6T27jBIV4CkHRRgRTYruukwjN4pKaoWXwGnCnr3
Bl11k6OCcWQdfVdziP/oexYPdMZkJEJTUSi0gLsHHUIdeQYwRQi+6vowGubUtkX2
E6kEKZvp+9AWDH+tItSCuJ4OxNfZvwpOZmun8Rydm/FPCGYpENcckIG+YvZomzxj
8mpaIetCKnByQ02+B/6FoFTHSixMpN9BPuGJTwYVGqxculmqwBNdoQhjniPzhXaN
hSbmnnPfGeJsQI1hE4DAMvcaB7qirLGKrMwW8tm8zB7SQMeLNviG8PoJw7x5YnqA
cqA9lIHmeBGF20lOrwwX3eJAGf4VuhAt19B2uEGULrI+m+xZk+h8XepUmGeTVaFw
SAH6UJ8o+NpHezSXTluQksKYtl9f9xEITxnoKmDutbaUWnPGxNoe0i6ab0f/kBf8
fElbZQhjIvlFuz1jxSUozQ6ioi2ghZvaAS7dvsix0+JjIeBI9rnHc8bAZG5axKns
dsH48uP0o1t/Y8COkBwuq6ADN9Dj/hh4WfCmCppVVKadr4W7QDOZA+2aeZH2Ml9P
gd+GEh9T3AoYkKvTs3SkayyWTLbh6rqz+TxVAYCSBspRHiPQTea9k4NNK2/rvJfq
g0MkmqJ7NwyIkSmA6S6pszuTxU7Rv018nTYdUfni18B9zKumDvWuA8lypDPm828K
Sd6uJeRumS2OLA6KYM7bfYWROz9xAdluQN5xFL5tV/YmbrI7djDq8Am6oDhHqLNu
4X8GPVdXnfmlP2HONtmp2qRupwO6SArIM3CFbATrG8uW6zn34/V7fqlbqXKxWbQJ
Lda4qSFVh7JJw10fjJLVXSSQgDWZbvDaj9T8c2ld3xQ/Xhw/jypvZ6Brw+s2V3g+
nHrJ1aGPiaKOeUl5v1X1j4U+awAtDe97QqZofdxJgdZ5gMl1vpKKNSTLCpzVaAmw
iwd8vxb9ciPbqFse3STby+ZXIIb/R8Soctbnw2u+LTzm9kCcZx4m0RTv1I9VPMDD
h68qAHEj8hZChul8FXwKRR95VEvJC6ETXeDMCyVRotXlqKIZ9Cje7hek8F4buZ+T
/7gbzOI6BBRHX6OUKKou28FyJXK4QsT71fI4v1d0RETch4MjdXLxwJ7Y+zBaKgek
RXdLN2JnLrRonbQO1bbqf7pMD2r0a54eEmZfZB7LbZSPa5yeJ6Fjsp0H5n32LsLn
pw5X3cpOjgT+xvNcJuuTstYa/dIiSXi3wZ/Zm1YRRKjjuSanynFcy3QxE56uPkQK
7A8RX9d9YWOg42v8SZiSsQyem5lrOKVYfR4RkQ+5v5R3ORcB3w6+m+bLQLFfiAA/
6BJWPrWCxCEQZSG9nu5+ZZsCquMcFOThtuhOyrQMjgOk3NKjCubUWcQTKKhIMx9w
oerMVTERVdDVaxYKrKfnvpGM6ESQuzlrxgy+v1jHVW4UUheDqEIys39iqSz4B6UT
SZvlMbn+0ihX7OqebBHjIXMd7p+OMTLR2zd0JduI0IoDr9Vw/LxS5QEvMln2bxQJ
6K3cJO3X1/Yd00v3qC6Lena5zAvBGOpj1WBOx259PTBKqcQTxJnG98g8zKcxujwS
o7dlsj0XUqjmyyVuK36b9RFnkKmSIeRH6PyGm2YAez6rQutYmgfXsOdhh/D6LppQ
h/79rSlji5nCu/9K/6K3XZUu5L1vSxSSf8XdmpKcYVFc4NQma3mzCh0m1mcFzfwy
0FJubRJPUG0d8l8RaEo2bvxTZVc7iTiMZ+ARoa5qavBctcp9/DsHbWVxhHbjQ7dF
DuzcCVEMiY7Ka+lfeSbNFLFHlnfgiQy9mMcG+tugKpdO57vCMHyAneV8c0+1EDO0
uyvGO9LBu/NylH0qKYVtI9gzOP0uirteJpEtG3UJghpux6egaw4scw+J+bAGcxSt
2jUjnXKmxndcw6/saE86BvYGVQ2BkY0qVYJmMZKhbEoGqN30xzDA/c4AJtcG5KjY
gGkh/kcVnaSJTe+N04TNliH1gfvOgcJw+6hKA6beG0oysHk44JdNkCW42AVFNZPF
f+Ooa8XKolKnowIz/nFyq6WXCpv9PFAbd82dxohJPVCBxCK0WKBuvzicj2Nt+NfR
KdfYLN5WhvtkEdcFhHjtQDARR7B4Aihi3ojGT5dWYX1xDRH4Ptort0eKI2/CNSi9
n++TdjKwyJP76BEUKit7/pPRsVE1Xc6Ep81NhLFpFDE70mibik8XYzf7eTVzgwKZ
pcF2k6IS8EhShYAH7k+RDow2HibtqaimCdPHKad8dJDSMZ7Zrg6Hnyd26Mvx9y1/
EQEnQKTn3Z2AjhCYjq7p8gBC9SL66WQVdEbvidJ2n7v3Iuj0I+mmyBfayzYa8soh
MtJYaloR5RnwOH5eUTFrUv0cl64tpV3Dhfamo+C0q+d2DszL0JpyhTPZFSXx/EA3
w2cGWx9/cOUwh4iRO5voJwZSqqp6zaZrhGS/C6WigLpa3eHehMqJylILUOCvCSei
mmKmVvZQQr8ee7GmgsJdHzKY45MBVk1obdvxpAs4OhwTVoKVcHIDquETmoZIiBoV
KrMEmE2hIVZWhTM1rdY8rDUdyHMaXwR7+SHlp7SLWF+owM8FngiLR7Kv+QcBeIxw
IZBDfPPJGRuMORQG16qztAonTQgGMxjZ/d3CJ284wfFFQ4F1GgUTm3H85dclP/kC
LvxEFyp8WUPZnPd143OK6TApm5lICBWQHKwEjjwZtUQtsdDbwa8NdUWADN569C7X
bpoquPUeBZ+0aheJNPw4vsGRdQp05z/IGijiIOjOk2dr6YT8xF8yX6nYh8w/6wQ5
1880q+rt9uHFljgkeKGM3mgNHs8Mp1V3NSpRpP+tI5gPR2fRpTxBTJhWg043pKuw
5q5etDuWJDMbNDA/QarNAdQfqS5wLMvMwVzmC/0fajIwTUxx4TD8wbUGsHXufbmE
rlW4/Pb6YNkw0CU+d41Mrq41ZFcQ5piy3lWgrpSJZZQLjZeRuCNtyE+wgBXyeMj+
EtFZr6tcJrKWYAa+lalM1yJp4YdVVNYjfguyA2WnhUfvPk004laUb6desr7qhYbA
WqSPCY8OfR9vEKZHsi+9ElRJxGv1RBvPcMbYyMi5UMg76NP/ra0Jy2vKNzu7ua6I
39p9TJvlbBCPBwvXXz1DjDej/VXXA49PrwEx/dilbglzKBGYlxqFWfkOHbq5M/QQ
MBBMIFV9j1NC4CC7PCwhBBIwn7DftMxLp0/0/U8umlUvVVXmsYVqhf6Uahl2/QQJ
XdlL/LV5YxnyESX7eDhxk7bknxwRJ+TL+WSnaa8PuEG3IIcy32APl9bCrcJ9s//C
fDhmMHEM2veMTmTJWSSw+z6UNdUjWXPLzg+FoyEZUpI3T0G9e/CGzl5mp2sQuNrR
R2YRXtl6isX6tf6aP6Z8TZhEYoL2FP+vMyHiOexEkAt+jn8AYD7AbrkPMslk0RHY
SHvjws5WMHR5+8hY5Akq8AeryyxApeBi7JweSl/EY4H+TkBvrfSamgDIb0aU+AWJ
2G/nfzrkVb6bu8UzjdeK3Zy2FQTQ5sB7AbWTM3DU7Ctj8iOgrsBAN+71E4uaUgYs
CFZtYkHS7GboVfQqznaihv9jrN6qUkgkFq3oDLkYNMkGbsdAXDtNNkvIA9JTxyun
bzGAwkP7I3U6GMc+anP0wI2RJrxx1p2dYuUn4HrrTXbd+tAbEn5zzUHp1eoBMP/7
IBen2x4wpL6OsaVmuL3+uDrFcXsKso7At4ehTyE0DeZaU8wUZk41NX+akxmanFh8
tRP6tr6MYogSOMypPtjoIdXR3qL2qJ5ChnnAkMBS+PHdPzvfSDn1T/kymPINOdCi
eRGXEnuBungAFZ8kIq8M0geRjA0ou0+4ZFNykvYjM45Gsvv4jFfLO7sMXVfhN9mi
4d32RH0REbXTsGB79FqD5r6Uyuqxko6zYiNRJmvuAopQhfhpmpfltYYNNwjolUXm
TSkPjnYwGpWhiIjMVGRmIzH2fVeRC+tQn4hO9Tt2HWR+ya0aPPH/BEk6oK/LTTKR
2m/Jj5R3MuWJwY4LcUnRVcP1dU7WF1vbkprOawhTuoi5LuLooF5ztR56IGpG8QLO
s/0MYTLoAy5HwSho+xsSss5Nx1C25EeDfrLKMV2NDIXQwXfwLzWK5SDh1itLS631
VA9LkY7/FXabygFptz5btX3vjfUTdQGcD8diE/qpGALFH30S6JKmLrjvCfHLPAOu
gXHyNGggftJBQFLSicnargLNzCj3ky/m6iZAs2VPg8CZmGYPQap3ASn3IeTtUHO2
bg9k1WJWmkqlSqCMwqN1AS1flidYc5FUlDEDehfAQwbw2NqRHi3AU4wiq9vL5Utw
130AdzK0Z2btAi57NZG4YZOGS48QRX+HElJrims0Dube9NcWqcx7AneUmNAQk8aO
ufshdlwo+Su21+w+afo8enNfjEzOb2fKmyKfzpDGy0s/RHdq280M+wPcN2Yp1UoQ
NweJrTOddjX+nEUheaEnR6pNzjmNZkQNUzOiJyk/kJ/w5yct4Tp88zWumpUfuxXv
M/pAsPVnBHpYLYjvD0itXZKZX5yascr8BH+AiFQOahuGKsjx94aoauDLmofJ4tIG
2pVtkHtnSZjxlgqNbksOFwrDVmyprZLsIKupAzf+ncO+q1pTp5NMII0RMiqyuz82
e5Yzf380oCO3RnbilqmPiRyqKs+IJcxOE4oNObZ+r5ZzuxLek8YGY/blRuT67tW/
ba01o/cn6DCO0T/FRUaaPTCk2vIxPlX0egvK28bve6DJ7E1xeF1RxY7ujOFkuDhe
F97fI/WpecQXYIs0K1swwmF5vBT9i4bgfRTKpXPxKlI5c6oeD6jV0Ovu1vp2o+Vi
0IqZ55BWHU7PUd8a+jKVCsZtWM6qRwTTtjXVk17LlXLlvUHSNCf2nJPKR5LTI25i
VTJjK3HSX4H4zzSx6DUpmLNhs1Sgp9sN9wHVYGtZpkZGt/2U+9kUkHyG2M+aLRAY
92Gg0I6ztUuI/OriFrzGTLgAVV2edDFmCOMz5emAAUjBEYWJZKLvWuJ2sax8Af1I
oX1DjVDnkF7pR+d1y/ZR+VFZA6tCwHhtGdd44yyWAVQiIav70ZLKFtfkbOuU5db1
L38xVBwW7xbXQlVWLJ1ABSxwufBfeR6FcoiCl3JT0qIuySjSIF4F1wwA/PDpo79F
ZzU503xauh2Q559+P8U2UOxqLdb+/9s0bI9/xCsWtaGTIi/FiHa/6+f1V2pZczxt
Z19xTUYbDZpE9d+n51L6XN+fA9CBlRYcSOjsqFwQ30tPcqdycJD/nIrxAgxx17pp
mZUjoXoZdj/xo5JllobuoGEiKZ4Phx8llghipOMDJ6EhblaLHS4JjLK6GTE82Wou
HiWUkosRXTKGaax++WUwNEO3kwkxK4APoyQVQOLSkABnWAHAetd78zMgxIx0Wjic
+FFAs6w9hiLXJjNXxqXivh4a9leNnW22zT036SRlU0FYhjnMKFAIz8TGLV53Ct4v
mR8v7RppovjJi0BsHOXONaqoVcATeVYyqHPkP0VQ0wIubotorqIc4ZyeO3C2tCWe
voemznTYamnACHG7lsNhCsYH+CGTOU2ZNXs1YhdWam681dWoOlCQdYPABx4oln7M
xhCNjAsr7ZCyNxfHK92iQt47VU/B/sE4DAoCDjcse5bTFbheoaVESI1MqHdsgtmK
FupldyUBGY0eN8TkMe9TmAsUB2UhNZKpSKOGkuhCMuYcQNjM3q2wposK/aAPIKj1
cPA+Fk4LDoH/aoUcEjX+DYiqIHtBd7pHRUu+1hs66jwbEE0h4kCD3baS2XP+5KWe
o+KQy5cnEORn5aWbdPmua3O6sKPE35hijNpRwP/tNfSp+GH8eBT58oYbI3ajD0fj
ipS+ohXoVEOZmkD+9kDkBG1zetEfV4Bclh8RdhzdC5CkA1chqWNNJzgZq2BHf7Or
cfVu+G0j/LQTvRZcFczYSusuF7jpCrBVt0si+YG6PH+cPmsygZviwelMI9gvaQEh
5AAvhmn9AZozqnbsdp9MUg8Qtt38VL9h38dQdntcSpO8upeSOYMCg/uNUywRIHi2
Yk+EepDhm7WtZMtO/yg+PwMbR+Bka4KcfA07GN3j2SD+sMvIirhYsewSshnjprjz
uPJ01nI37AJUBROi5+W0qoxaEfEnE+422FLVx93d5svpCHwIDtQ1RQQVIA+DhFF3
IT7GQZENa8d3NVZdKwW4tav/fC8NK7HBxXrAjD0N0oqr8ApA1GVeL+Pdwf2GlNif
f8YH/z39fXx2iP0ZFQQnhcsljZqxg7i0oNHTKdmWIhJWJoRzxyhVEYgHAz2P8FEQ
WvEeeUg6b/mitIXmGNcisLQ5701xbionfAi4vYwQfpp6+QGdBCnM+KuUCDGI/I3Y
qskQ79zx+6AQrFMGaHHVQUn3HUliykHtbzY25iOYX6vsXkVbUWcU2ItnhmHpsAxX
ZJHyxwURTwLEiX7tHpfEYXt64miDUa0VZdn1FTdDvf11mG6ZCQRR5RlR4hPYHWT5
FkPF1MRjXK1So0Um7ZyEWiMi5CRJ4GJtaiJPxty0y3ICSxUnBE9rSOF2khYsocH+
tx38kxBYFKp7Sr8rHMoGiIrmqhJYS6WhfoXd5n/MMb40AZwk6lvSXYWYS8Xv5gMY
hDDxVuOmqoJeS7f19RVYqgrSaxs72hBN6Ns5eZI1l2hTbhV4fDUty94cycRPzRxW
oreWHaqryNamfygMrYlTeoaA3NO5g9TBK2a4oQq5CquhGVqFGsBkXzTAd5vyStPO
BsidjpLoGDsjJnRUSqd1vDWf6gezT1hAUQTuUNWt+gJUwj1RYkV0IC4X9aRHRvZf
5RWAvBy/ZIfdGidf3jgaOCJ3/+6AbzylaYVGi9nZLdavz5TwqScUDOX9dEU5taSu
bwHVbqDw00J374ZNOga87N6Q+AnVHyRvk13Ydpe+BrD7RMqHNwMBa4H3UxbPdZ0V
AbxCY7bQhMf3NV9g0hoDeC1bXoMDpdyLXQSIjrTgepOUqvelcm6qGvm0PsVVKP//
iObU/7oikPtrIeFsvRfM/eV6q6Tf6dJUseBkydnOEy2L6LI73ycTaZCGgtEW3dsp
KYj1M4F5yCDgtS0UyClorqRp9J2va1GYyISJJ8W089jThntHnYGg0MAnqc3xZ+vV
qENKZvjBCWTHrToZnCse9PeTFHucokCFsD6onRlZ3NTzamSOJGox+sygKaQz3jE9
2j2LjZo0+uGe7pXMYvbsQrHNje4k5/0y2KovIX/t4KYpvrSWdcbnvY8ce7dxpXFb
Tn0vLvhth2F3VkJ6cFFJIa2/0w1W3JjWM7aYZo72jB1qheKFyZB0kuu6VVVuRLsS
SG3bbmUx5zbzRpCYTL8E7WY+493/hjMFcwkMbBCqwSDkeKL6dh9pfcEXzxfISKBp
OeI5tFIgcfVTHhnrtpfg0LNq+mlQxa2uXfnhBG8r7ng1FKipdlvu8eWdcMGwXiiH
x98dYmBEFZrhIo2QDoGKUwP93n3XsE3iQcDiGTw6Q/GkjELQPszaWW/oWqYIX3qD
fJHjsNWWAtZk/XX24BjeqcmAjCLEcJriI9FoPgZhBnPSOcpBwpkK6HK6lxVcY4C6
3a7LDcMtKi1DtKDmvRp3okLNO0FDKdcLUJA39jjaOVqdG6LcrBPm5y363eBfZ+H9
c9p3IYmfI7vVKMMqfNfUEbUgoXH5NpxNwrBAMWtLw5qmGtXNjJf/C/YD11D68Xfs
is4+mc9TT4+F8gmNPhrfZcqK2PJNfuB42FiPYZgVAwsFgt98okr1FubkQCiDpZ1S
+iyIGFVjn1EdkL/0ceVFPCkDRGbFgGTdd+T93BIw+Igz8DGOmVcwK9Vtz5cYlIvk
dmqfUEXgxu70aAXXtTKaKG9g8C8jq5yPf7izSQabHjb9ep/CvvSepEDU8maMjSAE
q/Xiwyvdmi22rIAdAELa0wSunddNzlY9IFS+f2Zz0ujz3/5okCzK5N2UlpPZZ3HH
z3BOiE8NAM7FOVlGY+fnw7EmUaSEZd6b8iwQbMqWfOkR4OBRYDgqEUG8bp68evmH
bCOxm/5SoK+EMK/Fnp7rCM3n+CfCySBIzEWSA9jm0JY86zQ7n+v+536c/5+0YtRS
zNnLUY1WSJhepwfFTWULiesfUDjjsqzFyU1PcGHVJr6HU7fFpUPNJE+SOmWWC9Q9
PGt6swMpResnDAgFRzdLFq4zlLDiA181F7azT3vFfh93BLV9KsQyH7Jr6PH4m/AK
GSdqaiGhqS99d3P3cif6BzI5eufil4mLcGnzRUGk9nDt4R2MxzjxBXaNh3g5BjMv
X5mlYPxLhsr8KhqcVmO0V2UYL88+SYOg4ZQgZ6EWkoJa4rymFvZ5zTiTom2tarS0
sywjWEV9HNdX0+/zCiO7QM7YMq1jWw+ukosJirMQGZ/8Jf9aBFfszfQso/BHctMw
I0HJJ/N5nBN0mTf7HO4phCkrco6O4YGkuiSkd5L3n8x6LRHHVZn87o8pWfl72Vta
J3Cs5nxsKCT9jPj6qRQxJhR1ZYeE0Z0TES4qdcrfsALY3U8u5M66yTHS2q6vcbrh
PFVb2c/CNssVWgvoDkNJPXoA7IobPED2cx6OybGxmIqdKjmZmRtkHyziwkMIxuTn
TTYI3g2Q45uUs6YM//J0GZcgzv7uhJwgjjbF6WsiEQ0XN8nsYmD5pkDz/YoseP6+
BTxBDic+0uXNgvtYIjrsQN7lK8p7Hb9tjice3flbhzr8j9lWaX4yFocxleRNl+3S
2txp5t7th0jdm0Zf7H7LteVw99reuLMfo42rs9uaMtCoRqArVwUuGcvmRXxYlrbv
CauY6sqjimuFYdCaCSkWONmzDkErbo+BnLHlKLlFK9gyRklwy+KVPw3bSY2vC4ms
K4Nu0aWF2QtkDRe6xib4Z5rg6jojpyQN33+qVJVzGmcd5oitGEvBefgZhbB9l9WV
pFceE+l1LolDWcyNAFl5KjKQ7uC2lhQrSqc2+1f/1zfwdhBAl4vJFn+JmC962lxc
Af8+oPV0CB6IXEvtUxLyIXeqRhRE42ztjVy9x/fOIvwB0SfSQhT6tB0DRmconoCg
1NL+oYrJCQNBoNHGeHVAOczCIKawIS+LyRH1Bh4jCBRWpdqKG8sUvvhUV6bv/1i4
VHTRR1rLvMSAIlC62jryE95NHlqb5IwUSZBS2MScuctWHqeBQrs1xvx1XrXO4YLX
1CZ0oNmpP7wOXXZ2NYoZ6fRT0bcVoDfx1y4H3pp6GDtKrpbcYkdUiQVIeXon83v6
Bga0oInfJQUIp7exnoDs8EpJM/GV8nB+IdqmqtXPkhLLkhPWWtsiYnUyPgL7t2fI
fs/5sa8D7Kq+8a9M/KzZEjzx2t6RmcKDjMWNGL6PKemwDnuqVc0Wyi5sntW65cVv
5ZdsSc4xPik97PIHp9JjNhmxXoZMhlFNVQsa83EjNi0WeeDhU98OaEgOy23DH0TU
jqlO/orDAKf+2YPWVP7eDRiFBW2QAXGObt09vz1xtQbN0ygg5sK0ZACXXjsJl1kD
U2+2WTqZbw8TvYPHzUxtuwxKdvTM5ZyrkHf+zKbf49xqUB63wi20aexKvB2roOmt
r614+P2PVGM4VaFtwtTouUBs4VaRcSUh9OSANiNQ+/ckSC83cr5h2YvyyJ3Zf42d
zDWboYH87zhV8oibuB9rVFjzGmKc+t4palmLQDDHSmZq7iyF7jYw7F4IMLMGBubp
GWB8LQ9aWfdzzx4z8Z0OfQVjZcEAc8MvvbD5SXPCYGIG0ii1VPBBGc28Ex/ATEg3
PfhKxqxl4+VyCZXpT2aa4QET4eVgihVFGevZ+EyPdRO/DhocyQphb7mnJNZAMh0c
sSjKgcJB6ZVzaf3ps5LaMYv6pSt+h3s+RW4kiUnW2+QYWj2FunHlDb/Rf789R2l9
UX5z39j1kWb4frVJYemLL2z8H4CY4IFW3myyMsI5jw5MShpcpC7FOdCErQ+d675k
Wy+4YmnP6PYbZbBNtDKk2191WHzhnBk8EuvDLpyQqO7b3mgaOCw0IunmwhPdPRwo
hbEL2+KGHVnI/PZdFvC6wSzzIfEdiPXX4fA+UVj5dIDgvxSslZ9ChpRHseqPt3Uy
oVuB1JwkoWc1Js1uI2p+n1PswKr7kokqI4LiyTrz978nMSZK9nMmPYNOkM5oDzPn
+D83CWafr2/eikuVVQK5IgCZ1SIL1WUwPKcqAcMIMrMq6AtmmjHQHtxnABm05YDm
MV+Wi1Ff0m7ZPe3NJdN2bwAU1rt3z1XHqMUld0ZbNLfvcAwpvFl5Pdq7ndVaCzma
LLjrTydSdTCcD+9YVxWHynabJ267w2wVflTKVlgt6h5R71z/jrut8Lv3VU1EMCud
vQ9q+xIGjr1voY5bfmw/CxFCQjF8ooWDdZIb1yW4aCICUCuWoo0UlauCbjzu6cEX
XdOG5nFBB67IfXqOlojFHzSWAA50+qIyJtZrsVJQvmWA5s/WWMUtkQeuKO0b6pn/
BmUFJldYSzC23MrJDo+KsAGO33xZww4YSWRewiXEtYsSAkfbcLptf480Y1bk6WK0
AgTMw9gWlCvQlDRl1xEjWGYT0QU84TJAaHZqgvI/4/H9PnvFmA4NqDJ5YJVzjdsu
M9YGmlMFJ5Qcs9OXlNeE5IUpg9jtKuh09y+MdmM2Mha7klinD0KHCZYpNNYQoEQ+
3q9u66Hfa8tL9HR1Htp0FxZzt+AeNMEj8pQZLl4jztQCqFBhWnjqwgHQn3w1LqPW
SQ3bHLndbfl3MXGOuXa46nWvV1MXZPtqHiyFAsHYvM4u1dsdDL7RA6AKEe/VoHA7
kYHbnAEaSe3OcjwiKgQl71JTTOtBds0sB4/IRm8QBjFUfw49lmRhdq4rYFDZGvPh
oLJANJzYa29NQ8QHKFH9w2zqkmpLMdx8rQLp8XRzurMAS4/OsfEyuvZHWxAPFlK5
7AFwdYbpJvPdT+f55trzi2p2EbufDb8eaUHOg1T5NXtBOa/KaMjPfn2rivxLEQFA
OawXt2sw2o69ti7HlZL9BypvBnE3XeygNXh5azwbOg65iAXDV62YPQMXBwYZK0ia
RZlTPawrOb/XICLvPrHNZNlajwtevhZC4h2Qzlp9x+dwukmq8S6aRpM9yTCAEmqe
cR9BX1GawcrFbKrx/Kedyb0JxrXPBWM3cdmtZPfKCElCowPSIZ/UX1BPmvis+0LQ
czn5gYmLN3W0qB7Gc3oOiKDcg60lDRkIa3QpJd5cFEjXNHgzzQua2gyRkNOkmSpN
rgKQYOWXm3fc4zPl1j5WEl1VruLIcmUSfekeQoHZ8MTl6mG39uJLrUpTgF613+ha
BcBJCjwrQmzXXZGsxFa/I73lkryfTWh4b6ALj8rStEmym6KaGWTmO5O0KOriZEKL
+pyuQ1HRdG4sFnoRyqK8377GUGhWjdCjw9wLxM6cDSp/lpha0s5JJjWQ5kcjIcui
R0hndPQznUJgODm7vSDX/4dT1DY00DDbLOmqCxO+EFGpA8u8AZvSSUCNUCpCxr40
z5U4xKIUYfv9xgtEfoMBTCoiY0DBUfeGd1ZHaA3jxKEfWfciHk/ezjjCU8H68wIG
AlZU0X+bfmbdK5yyHHbXhgCNaNs9E3d8u7KvXXyfsKEhW4Ckrdgm3n/Ty34M24VU
k7hSbcjDZOXSEKNhgKY28W6Mbdh5pwL3OcQVd+HyciufUuYrDK/jSQxV4kHhSr7V
T+4lG6jH8ejKVSt3PrgZMSnfbpOMxaYSg+XEgQINOzscEkUukF0+clsRutNkqtre
dfuNpqgTJ8iCvYLM7eBWQ4vJv/R6VDFtK2E7GfiVBPcpUYAOezHPZUIULIbnq4Qp
kiLh9UvkiM0gaES5cDtYy73ec0ajW7fhmSRbQ1q0zfX1jpqRjH686rAJFqQAF+Qp
UXf+kQ7l+spi/yFCmGMWc2VGG6MC6WfEMTzIrNs0/yDZwt75ViyUXZFfOzgCY1Sp
lQJvVnxyZmUNK9pl7EVtCZz1Hzq2rxS2xOQV6X19RtAnZAW3Gs+nNM7eYFUEZz9t
3KK4D+MulubbW3yxGjMkYC/i2e4IVjq4MY3pvoMd0hcr2M8QtbYDpo/nYpd7oEDm
1RhrWR8oAhakmUYfCMu4oAOwGYVb6Er5wYdUVGXeV/avruKcN2dXeBFAWDJgO+dU
kCw9xf06o5Tb0jYHVKUWdWylPvac7FD3Cmw/hdHTCrVcq//dHU1GG5ZLaVvQd0UQ
Q+BeEMtJkNFKp08aPO1+GJJzrrAfYc0mrIAXV4irCxLi3okfy2r8n2pGTI2dD6SW
ITV5f/PXLKtlCpZi/eK7DLd+aNS2NNEdU/nfvPlFjYRjdw5ofx5bxo3+gB0UtI+4
1Y+UZvvv3Pg++xEHbnY2pu19RMScYLEYKTur3+ZmblT6JiCerUvwfu8/SH5S+kRY
EmdHUM6vBkB3zu6MpMWwsoKkPE+fpsyi+jYY+baox0ASk5p9Oeip24hIjzSfXgXI
AFMtBFjDeWIP2CQt1bGPo1WQr8m/9DDUqJd3Ku9Nv8jceLUUpUpj/E6oc5fswPT7
6rWa8atYOVeoRuB4ZG/T5vdyF6nDzegk7HBCFxLeMS8MRWzMVbUP+xaLOA5VxNd4
os+RB++TLfO1Nfr+kUVyEh2UdnWgPBIdVunlg3yl/ysQCWf/mSokolex0pYdzEpo
BMgx4ag/1xCQs3Y3BJHXUVfhdt7nYEEYKL2fxhxtkHQssuHqjDJreQG7EfPFUNLp
8pb4qRB11/8Yp7nLWr1W+vL0BVkFuoPFSPvlk0G2l8dWHfIdqx87AUNdMEc/YihG
7CaVRi19FHkkviLRXtPIIFf45T3kKre+7+XP/fQ+qweMMwRqLLaW/kxn84AnZgw4
UkuLUlyQsAHldrpmAP71gq6sFvZkdOyptmd0wVKOPpzhGaP9oL+QOLL8myt9Ce/3
nZ+LHirJCaZ8/fFvKnxD5xyLc4T4NZrA/Ui+nkcqWu27I9qnkm8Xy8R2YYXsvv0t
Q+KVnwllhUxYMTFiXkjk7Bjj9ShCC1Ua6c20/Z/l9TdSAeeSjIFSkl7VFi8PXIHg
aDacM2DgUNfYxJOgLQCvEYi5lortAirisQhR676ungTQv3BxCWYZeV/oYphUdXdJ
8YQuNEUkNW3hME7bMT6Ce4/lqGooqyZjsTGVXjBGZRFbd+RtM+RO9FeJtRw43//P
yiz006IxFJyYEQMd/ZX/Q8IRIfRuOWD2EzqUB6VXKRP9Csb3+6Kf2Cuz9sXYJQUg
iq2Kgw9cxyjAfCN8p2RKdBocLGmN8tGwZ11JYElplvPP3MWx8S1Ki4Xi1UxJYhMx
lbMWnkn2s4539A0OpxzR9DUCh6bHMchRBlOSepMcG24fadn50kQqN/LyQ/9vMkQv
4qja8b8Jzr06LbB3Au38+o/LyjfdpAmRmMFF52sYfvrDcVMjv1atTwr1bfT/3frU
KfM18kRK4CWsI+G/oGbhvGtkyQu0/6iy7NnEuvLozS5CcVEulQUjLixFyKp3enPI
w7ZPOnMhJvR2c6yz7QEUbdExZ3hiIgRgB5ABQAoVmRD2xLOUKW+K4d9tijzfgdd7
PLzR2RgZjL7s0pRLQ0JTuI3kB/qgnAYwUUEN+Cb5Y7/3OFcZxzcREBr2ZzwS56GC
5W1I6JWsdFJngG6OhB87Z65tQ/6XlmfoRWWIqhT86exT+NOREeBf6pyfIkOR71cZ
k7W49QKZJOsy99jxIrVx/h8vALYsQH9rkpnSLoyU2adp3HOQ9DR1Xpib3SvSqI0l
zRs9I6LHg3ACT5kGuLXAxKFFqA5h3gK5vfZ+3UeU8v4LsTt6jFAvLu6ihx98uTeO
4YIxEWDGiKE2SGc4fAyHiw74cR+m+D2sqoFFuLttrEdAef7HCMwed9FaHpXxBy2b
C21Da9nY4f2N5TG7+3OeUXJzmhDK0x0XLuWr2aOmCGj8hYehKGjIxVGkolqWJWRR
XFos5leB3udV+PLC7D1vLPb6H6yZzKcxkzZOqNxxQmu8YoV+oMwRm3SWRPAORqFw
CffR/+QJ/Vud4qOd0kZY/AcTUuMqwRE9ttRnYEyq+VulDZj2vW2QP+3JLKlTe80c
70YO3zSoF5pNRdiKWdYmP/Deq5Tf5i36rhnrPVukIQxwqta1mg/Sd9oj17c41OJq
U+lfWHAd8qOljTMg8E2VKk7T/GD72daGOmGyodD8VgTXC6HC+lHQcSN/pDg0CBkE
KotFhPQDcst1ok2hzpIpVmel5bjgF5ggxNxAd7uHAU5j24MWV2w8s0QBU2m3c/Ok
UdZxqAeV0sI/uDPxs5yrtcbfPS6OB9TLv4GyuBhevVJQnp/bXfCZ05K5xfslixo+
M+Edd9syA2xxF4fv9NLwtdpgrnyCurH1SHrF6tGK/wpMDzEiNtDmcgqJ1GRlWo1U
MwTLZFAMoEVla0yBnKRY6fvxc2W/YnYOXeRDBE37mFdOmUUXiW3ctVuvPpxuyOBV
GcPePmLmW2ZD1DC8MwLKEEx3MVQS/u0eAAjXkmna0bJAB3DjTozee0iq9dSdtMKI
PJuNoqYL5k/I0Iu5WWAO5VCLFHEK/URjBpe9pb2FzTH2Di6k1ytt3p+mzkejLvvF
H7pyV06UBsU5vZ39BR8tWtw4A72PgFguzPvRvLApOARfA5Ff3OtZmX9mkSq2XNat
Q+f2I1jzMUS+mgrBv7o9SRzixsTnDLDLu3Ur/viSLAYySyAI+yzJxRlrTg2QtVuk
hinBBKcNa1dSuCntCe1w8LnH3v1g8ZYohrrlDk6eLOvzqpb6uBh07n/VfOznFt1+
GWcTB9fw/o410hjSgVHnAPRwQ4RH/YBnqKaQ7L7Qu0Qs5tp+gD0sCzTX/D9NwQPD
MGsESL5EF6nb753++ogzlKBm/tPmLfER2iqt/RPzhnUyFQ+Lw6xlEDujcgUZ6nkB
AQ18KQM21NXTsyHbjCguwnPTVB4hrU5RoEQu0SvpswT9nntMaLJOTkZZpWbLU9Y9
L1T8pUg6woZakt5BLV9TpHJvRRGf8a5Wbo4QfGtIFrKuIH64mgktRzwA7arZlnEc
Q52nn/ShPJV0FMGUeejzhKwJ6ad9NS2utBIQKKSYAqTf0eYm5iYhzyNc4RIRxB9E
vXDH4to9Gr19Q8BYuWBjv7A7H9foryz/V1OqtZ2GJdoMARixSeNDlenfZhSveFLd
Dqi8VQBOoNS+NFKFOo/4MsQkj28+rsLJN6vqtAKUfR1A2gRnKM7bFaJdE9soO1vo
sN2XmNv7kaw2tjDeS2XV8NBzbJCqjgAOK80BOTnWXaVJXrYv3Z2LKRXpxNE0n4nb
hWBJQqM6cYryBr1k7+7AvzDHXJdkcMZgQnCIVjZ0x0/0YYqsd3x9vsiYvBf11LpL
iCfDIpgpQlP2TEkct/H1bj+FSsjIH4EOeut+a+EwhHvXcHU2C/fxuFbAlGV5MkTV
pZzoQYWRBvm0rzESNxgmS5jIRUgHWlkqnUYvaboZiJig92C+rXJA+UoEpYbqw2bt
8eadd3SZ1K/ZvRD5r8ycnmEf5ve0FnM2Hclw987emuLIVLx1svULqcijsFixCPIs
aJNdJfqsVtRpyGx/+xafRipQs+Qq+J+Du5vP98CQXpg195DVMnONjiZmp1qE2z7y
jeX9u9PhcT7pUJ8j9/0zfVXaHgD4L/HJ8F58zqGCbnt3ZjoRKTKXNkld7SMUZXWg
rDPfUtrh2c+Vg4v/DFnUP3ZhNGpLTjyZTAEDuQu/Ekwp+Q5SvQ6E+1vvGPQJjwot
KdPKkt4QRTgK939k6GHEEsQyDGTyY7HLgqGHR0XXLvEVUGHenHJ7iYqrSQ2zfRQJ
KH2Y3Sf4mwL7pO6Lt59UqS+7zqPbd336t9C0O2V067Q/XIYAh42NUN5pu0vrss8v
OpeArrzlA0/okoV/+qQ7On9/QnWjUtyH5p5KB5HqnncdMrgWpxXcd+KeJb7wbNi8
EYaYyvvsNHBxgak0Zd1E298SZhh2qy+YjmgH3/LlrZT2dOO3gX8EQnA5KhvYRl4J
SNwrzKkONghQkFvuUkASYVifSlp1SZxUGEEgRI6Qpf0lplLYw7GPmI0T1NgMxlYT
+XZznzwyIC4eqw6giTZsWO5JJcEyM9SZ5YE9cmdFezyvQoj/k3rqHhBvjX/aUnOT
Xhe4h21IVL4kScUi5lE0kd6SlKKtF0kwQvHzlwSpk8SYcQs/y49tIC0iPg0db/z+
mZvxobKrj/XadyhcBaRAVyrbE9imXLbVyt6zVJBTwV+wqOI6yfxTXLXC49unPKt0
NuP5ObFWQ+pDkIRwPngSOqHrcD9NMKuTc1Ctfklm4XaKPKSMx4Jb24vAIFFdiRhK
j6foCh7KMsm4T3vHxQARrK/t6T8Amo0VZWp2z+AMfrDcZBXbETaDGoCq5fdZDivG
N2DIZG/ZodAd0wPoELMd50DsPVqOmFs4vziS3w8Kk/mfweGehxbehzngIRuDXv5h
8jeA9tgKk3SLmDkit6ZiVo7e7TuLnTSycp5sUbphWYFMrcR22GzooTZHwCiYQcbP
gLw1tO6OvOIHXX3E+zSM8+efOzaKjNBaJxYLySjjAWzSxwuN7g4dXJL+nBv/8mKN
W3YIVzPeMs8AVmTTMZQtPDd4mElh4Tnvx+5T7S4l1PVRAOc6KArydxKGKYHr08E/
vFuslXVkdtK1Xri3Vp3wkwKBOhOhqfAuu7y96k3iOgpYRn8VF6VWHLOuH+F1jEEp
RnXHxqmpYGw5foIhm+qcYWoSpGvDIoy0TeMD2c2yGIqFiUx6V5X8Fem9vNSHVyW4
QthG42VrhxKpkDlfGupNhjKp9J0l2sN8mPkvr2WxW5A1c0PaglJcEQaxvTnKwPIe
kHJm6HHhpmcvUIfTGBKqRYMMJrNrNhUlaSJ0QFEP+jYZuCAieNw3MwXyAq67gnEZ
7KM5Y8ZISaFrKyRDV0bVLjiEylWmAtrEMYNkmL99Q/i6SYdaZW1ScNuTeMdMfYPk
yVYHooPkpY7f+B1m5n5jJe6QsFmuJzGPUMjDr2i2z1bsCAkZdpCWpqwjS8EhaGQK
iM4eiLasqAkKlKdjX6oBeR15Eds7CVAXLCaBIaNfHFPJ7lOvY/ID/P+bfMepyMop
VsLxLLgLBkWP394DlRVLVYyde95i4KamsWhk46mIiTNf6A5cUueDueYz0IAb/8Od
dRVkNX/YYqVrr5/dM+bovBVRC2q7zf4biaMxcJbnSLqwi6GmGhouwK9Xpe4l/1Gz
qIXX3PkZiKE0dX+crxkGeS2i/MJu7O+jSuJLsEnfLofUqwwt2sQ9r3rtuqbSegwU
MoHqaVMXMvDhSM5GXhoqgWWSBYcb2c91qKaU5CZKYJVySHn4ohtZ12sJbFjmCyFW
mCwCEhT2ha6Bt2fSrPtwBUws4sQ4qSCB7F35baB9BnPUXhDesb4o+/BEqGitoyZT
19iNdEHYzFM9ayNG2FLaSfhgxsx4GE6ILCC6jUycWA4M8Pb1IOCRgwpPF8GWHNcu
tfMBkTG+FHuhXZJY1Gxy8upS0OjPZKwWN7lzR3VQHEKaN9Wuwp0dvlebfztgiVre
9WczQgpdOMQZeg6Ff7/26zdGg85bhpILkBAHvz5oslFowRiCl5efY/mNq+0Vg4mA
ICMgbSKzBg/ccXevkcCxCXWPKTpMROF/C8rm3LTKxJBKzR52RJForOsm1A0UJFHo
CVGs8u9XwWg7zuu5SZ34hg3psJU/wACAgDpGwqqPRj83cemYWhAq8HtMOAtx5/sC
SQ24Nf1CKqdh5509JTD/EItlmUnQbiXeSJXDgEMUOaEMhYBo85E8WSmBEb1ytty1
9srvmynzYK7naHCKyfl7TZzIzSIIuR5BeIJzcmN9/+lv3REaPy6bmUGaD74Xm7pF
14V4L4of7Wwizyd96+PTWIy/hFsSUg4acTPjJQLdDzY7PHTWZ3orCF8a/+7ezxY5
pY/kYQTrR9QS+6Q90LhLnXUF472wjldXLJ1fWtRzg+CCNqXcuTmA2V4Ooua7e+6a
g1pe717ilnmKLZHlzbK908nUK2F0FSYu0fKW9Cse/YbMl0OKSt07oUgaQKFZLh3F
JqO8r3BtRy342770Znh2XhxsQ64nExzDdUx8Ao6gDup4dtBuTsmGtQ7W47fMjoxR
LSY/0nT2SvtChkZ3uAVXyadMENzaTLYujKVlvuQU4DpEdigQGMMpE4p7LzacBPP0
GiGQP2SmfgSqJJe/xWf68sPDxRBb4/+2OAI5tHV20mhaPqN70y38VJwRJiHnU1oo
sNKGPxDPIPJeLo4mb+r1amTkXvh6rOIYfOKT5i5QxUCxtRH8toSaYR8sZEyP3Rd1
teQ/rKIFIpA87w0nPPG04pS9pSnad1zOmGp9wT9kRsl+I6lYTezkjCtOZj4hXIrl
aFBesCjkPsS7oOJ9NBS4e9a42NkapgnM9YLebv72TK1lxoB2L4v5wrXco7UgJ73T
z636RelCWqxiR0jH2cqW+pGU4tVuBncpZaVq4MF4dt3Ky+VcoecfUVLhGk0V79D4
Qe2bOHVicJrTtbqohqG5Y8YrFi740BVwr7KsIWzrRyCZXHGpZqWTxkXMiP3cPxHT
NxeE/4/2WLRu2/ruKJlW0QArFzJUrMkX+k0sER4XavyTIW97+zRnWXMTjbEW07Fb
FMIUkmFv71VzTXsbp2CICfb6+gOZ6GkBGaaPueCHMcctzoRNrNzkMj1/mmW5lIsb
Hf1CTuDjizzJuL1GDHqnssW8THtrrvhmvq18zg6JLpvnkGDVT6ZAsJ5cD5Rtfs8S
V6b42oNKpZsHF7CAe4m8Ot1OMRLzvMjjWUFaHA2MlN6cxn5OkA4kkplzOvAAfkOF
/f6u0d5BOdeyRBzcMToP47Q1FHWK0tnK0q/DYn3KtvFxyBgtyHbPgsvGLRLa/AZC
fYX9MO3zea31WgxxHzu3d/9ypRBY3vQVM+y4qiG6gvusWoujovGJrtAhy2aAvvVH
YqEZpa339XjaV6pNIcGL9XT2+xQ/WWIQK7jduj5NHg1Z75K8iR44m+jSSYcI/XdK
M7DFgeK692zgZ5K3ZIAp9uecd9Fj1r62sJO9rISWwc4K9nPYgATswZkXR4PQFxlu
lGwPkQFQRQD7n7CQmJB+ZBowlwOHY7yi446l7kuMHhRkb++HDRZtD0M5qO1R8m94
730obu0I3f6+4v965xUpq4rdkiXjbfvFzP5iJd/KPzVxwQ35dasewO3ErowKVAOA
7UiWtobH+JN4MVg2UiHcgARxyOipnxYtoCgqtDmmXoS9jDCiUjUTQoiW/ZqsEd7u
a+xUXQDj3Dy3N1MBqpj+7/Eml4JU1REaGaO8V2OSAyfJX21Wom0tI0vNC5YCvu7x
Oh8YtYGm8vAgbwR7jF362HE09DY1DR49lJFa+crxLNn724BnLCzrMWFksum0pqrr
ScrhyhFYQHqQanO4qzAPfTVXVYDh4QUXGLA2AGoy17rVeJfeGQPooBvAooqmShfV
APt5HCQUJbCtpVoGvn3WvrMaFwZ3O68J8f4X58HCV6Kx7U4g2GW+uEDwTgw7kRs6
VT6VCCnyuzqaweiWGzr0tFhg+UgndUJzG7eUGIXL+NwNYBADIlMIyETa1QChX6r2
HpYRPlzGiBhglmxBiyRepN2+lY+wqDY1qaoPa67fAQCZnVnQOetGEL/BPmYSD2ck
0IwxjVZCP+Mk/55ilbIlbBVoH+2ZQNsbIHOnEx9tk2Wnpv2DOlJhVkA4w2QaiPhF
jYT9CMVCrdGdf/Zu3CuvDhhlIBzJAnAdTzJ/zIKBkcf6Dlyq6TpHIM+fNmvHUC+5
FN2Iwc9CmLQTAIkZXcNt5EHfktAHlIcJ1C+t+c7HaguvrIvBglBZrR9OsW4ET9yH
wTgpXTObJgI+ixAATsnOMeYteph+GaQVor53qftCvMIQaImqIxwt1RNDQmKRzC29
OKyz9X34htfbQqKK/zAlJXQGW6VgfAyOwhTdlgFkyKmo0VHuBoezHDhlot1CXLUF
DhWY68i0f4XIdIYeRYIbMnBQItKUepCHxz2PgekgAlnf5p4xMCtAqF04E9iEFzko
ODDv1kowc7+q4BElfiQ7UcG5THFaouMNp7MypyscE9jPBnIcE2zEFjpcWRstXGTo
+RCaDvbMPRVhrCmivqEnAIGbFWr0B6VbU13OLXyoAp74S9a0Pemj7f9dCLeaqTsg
m80Ow6adiSwp72C2ZGYHY7zu2+NsXxr2qf5OZ+acUdbnyBiLXNqFcbl+iQAQZacP
+LaRZNKu8JCBc5Eov27WmgLUbbPp0J9BJ9VQk4zQX4tPylotfElhyf8GgAGZEaDj
0HeA/6X+3VrY0Qv4/RcoHsfFxx/Zsdmt+br4LXeBCdADZUEEDSUiH1DFCyuED31a
SFNX+v7kE6Dx+BUSlI8d2qM26eqJA713woDxKDwnE0xF0/ulGI55Cb3ZJWZQnGkW
B9SvzWvX2LZ7mjCo+5iLqcUwqRo05xGZdo4spRWJwtB2usjUJc+Zh1DN/IifhX43
aZpIJEMZL9R9redB1WHQyAs8/K4gEyCcOkaGDAQzKn8aMT/7TllwHMAfCmSMLgcj
+Dpku6xW9QD9q/KqsHlgDLcSQ+e6POo1Yk705hx5Z/zjau773ELuqOVzQA4tsqgF
+EBhgAiWgcaxEdq36w//sPWKamQlmSMwOS7XSe1D01kpJf7JBVaW8iRCQniGiCGn
xZJEbW7xbJr/foS+sqTphuuF0H+zVJDJPr/z4R87F7fHPoe046lj+ZMNVSV7Ojqx
qv/sNpyI9JOEoI9npHxRNTwMEI+XIFHSuh91grfkwH64tXZNNNlJkw9FNmER7bjp
omKChukjBTbc++7bpB6QnKisHKbNIXK/AD1xpwiw4WrYgMCXZg7C2U3JhviAxzbY
nuPFIfyFxWLvq7X2N+LfbmuTsHc+pqmzC5MfyZtC6DrMXVj12lbrLVlHuITaxEcq
Vsa4UzxdrtVL53uy70/WjZbptdHct++t+HnBjz38QkEITmgNrZbVXjkkBUCvuRmh
zoIzqYUrM0P2SGYINDZrkU2uCNSkQg8eUw/98Rp8NdZ2hNOpDMbzq0DmOGkmyaTa
jW2HT0JMxWX0iYeUnM+mp6utv+XRUZHFcAx0PHSayk8GMaT5YlopOW3xaZuKHyWi
JWDMsMt7CmQl19zRZl3DZta4OPpTfjFAmjn5aMG7Lgbwd0l4eCW2i9YtbKCCJLHl
Jcc8SMC8JjNXOiFlpR0rUC+EB8Ge34PfGVxfAfuOzhGCC/5msAon3+d6Oys4THRL
fLvMhm+LEeWo0UrgqOpWLdvShoTkCNijPXMZ1R1ER7fFo/Cnn+vSZwRSJxYhFyxE
G3d0qFg9TIa1B8/jEnrBF1XsbyDDDUzKHdELrfuqDUXyv0VVGKAvvIRgd/RXKbXK
IEfcQAa4CHqNtu4Xc8zq2kevGIwBSPQ3UvaEzvTSxRQk0kCLLSOx7U3a6Pjzso8l
1sIKmsLGDR7MwpLG8FGzp11wC+jnHGSIMCe5UNtbMKn0QIK7EMPXOQeJ3Y2aw6QS
27hKqF0lEQLjUdeRcm8+tEByuj12/CZhKowD+Ikmbg4dKlJWWSGc8sXEuIZ38Eqx
ox5QDB1f+AbE7UNMSy2w3RZYZkGvLlPNfqlmF2URKT+CamzOBI5xQd8gEAGXhNJR
WxofajcM9NlGzg0A9j5KqjpFR0X4yWH5gRD5YO+5Tq13hUg21Q4LZCa/u0LQYT7g
mawNJX1HN9AlEFUKAGEkxynOGorLS1PjArhBCV9QEOSL+oeLVKKBRzCe1H8cw14+
GlrmzPGqVCovqCbKLzUPmaWzd2fAG4Nx8nPhaS30Z7bzYL4xdZyZnloy1RJ6Cr2g
V3TcBXxm4t+OFiQZVvgOLYicuA36tCnW1TbAhcaZr7z2yHmUEjP2Coh+4I1/Hd/N
BssGFlj9SNPWcX1aca2sGpxVg07bqSsHtAqDp4S95FyhIuUsFb/iKaRNIjb3WNL1
OPe/oVu4a8VOPBezM2a020LTShmQFkQM4BwfhkzgpYCqQPKMpgjUxsMsIosScCeq
pfyJWpyNT7oT4QQxN06S8KEBT5+TuIX10R+flRG9lgFkjbuuKIGV6y8ObD+SY6bt
EtovFlYYXpWrsQp/sMDyTrYXoYCujzH4wInLhlYLUL9/uLicgw/psPnYePYCvXmD
PyxoAM+j8GwGAhPz3LAIFciVyymVf1LDxI9uMXUcVm13C8JKaTD5/n70ii/FqQEH
zEq9aPt+i2wJ1dGoCt4ZxaxbdfqbfQQhit9BhQ7usSJhXYTAvDqwQXRCgTQFSo08
SFLyLNY8fiTOfcHugnw4RTuSkZPgxV2+0xW43uWYygzZ1XAeWbgsB3Jg7yCntDmS
e54obPXgg442RHxQJajNG9PeBKw/E6ZikwqUtry7lI6C/ewmGaSRFkrCQ8MAVNId
79hotLyLPcsLOBaC9jklLn+6dg6q9jLBBE5JAbaBURz1LJXirItIAFkV0QP38/Mk
WgUOCK0tfPPzZX1emd9Ho3n6cSeqRtbiYVfazvLVEcX9I2s3AzV7DYzq231s84Hk
ssdblumwT16/VqLZhdPdSYMt4TgV+UiivnFlH+FssH4rh9xGWRKls9BGJ0vlucRE
gnU8fy/iiJn0iMueaUWWqbbhy0EIXv1kpoPWk+HgCg/qa4ZUuhMPibaK9b7+D8zf
CTCBG9dSfYqKarbHShDRLYfzGyOughDxl2PO5Tq3vxpohdlIqVNWsXowbDf3Yljl
fU3dY+Xv4RFm+M1nPHfugDYdKlNFd3rvqaEgq20U+dbqZ8tqfLoI/2IurdnCVGvf
9c8aW74+TL3ahvx3hZdOnl/Rhxn64347Ha8MeSH69GOPTEI65FB/UvBxc4JMX+Uz
ICQPm8ed2+XUoHCJMfGsPi1TIYPEYlMcMKDmtup46sq4vJUh62A7eX8a+APbIaje
5El7RPQ5ecAb1P8avxjOFyiyqy6eDYEEUiygL5tOpRhXizL7exLL35kdVQqBOFWa
2/n0wBv6vNWi5H8fzoyov2F8KC4kW9qazunfxOXpWamLWpTSb60oDzXcevozGewQ
NpFf0YVgnScl6z3vsUp/ZApgFYBwH/qg9dstM/Q72EeD/j3uv9+pqAEY4BzF6Zh/
H2M2toBAoIKkBsgzqv6jjUf72kQmw3jxo6rSkCLT/3K+Q92qYtnSplJsAhdfRrfO
vLkurP1cSQJX/bjFsFeMXKk05b65uyZ8an+PoOTyOkOs9K4f2/STm/5hm/m8hOKe
5nTQss4S1gc2MHhMJy99MKXk2a9bD9DfQgfIRKUXyogUd96SrnhHKv7eR5QK+QXh
WL2Bg2Ob7eRRm5i9PLLeLHPQ88+6b1/PM83zNSFDB6LMebXhZPOc3v8nEk8p3cjN
6R26zgLqGZMciBxvgCj0ZgVZxuismXO5uxrLmYZTuvAO3fWKQJejgIGparj9M2zi
F1GifZ/qN7AHoYpt5CDdFbVnrqSSMRxp4qAxeJYuXM5GUhikE5HovZNhNFC19wy5
tQP8teFQ9fnDay+MAefGsWSeWdhktYbLux7GhoACZwIDBDBW6ca8AG1N8MgWewpg
tHrFCHJFlVxi8TZtyjwez7WHk/FU5n/3jiRj+2joYLjgn7/GCgvrcdmDCYA0xzX3
dfd2dB6aTkfFRlNOaVtOQMbdfE1enkmqfqIrr6qppySP1exYkJ3i6PbjifB28Oz8
t9qjtHub0W/YbroFSjK30CEviXk7KK6Pg8mtEAwAR9ZQIYCRxHvyGZ51EVO3R6RD
eQJKJbqqkAP8Ik5W5QfcShc2x2ZB9UvE1IEINK3G42jgZFLRkGhkVezeKVxuOJW3
jB1Ij34eFmF4w09Kyqatl5E5oBCuevj7wZwUzABx/KeXmolivBFW7RJpDiSnIt2i
9u2IZe7bjWUnRbIoIf2/CFWD6BUhMb2Zwnzs4n4rvbVDhSg4aFMGJg+v8prJY/QY
hlgnqx/ywy8RMtxhmE6lcytnJihp88VtacGS8Q69pPRHUlyp+nHw6WVts6Mho0sp
c959v1ECNJtw3i1ZWZrdBvISfDOCZ8qv6r79Zfd7nPAx++M4oxZmjBxi8qqnd9IZ
+Npo7q1jerHfIdyMUBOpSVP+biuoa+RjHrUqUiTWCBRKWEixT6cMkiNKVlhhNK3H
d6vKd88p6gfGv5FOC8zrjxZSvA5JQwztuO4z4wnhCZ4Ha66ti3HipgA4fjuLEBQd
dn/kzmkvoXmRReDlAk0Lx81NzMVC2PTOpCK7Af/ep3QP59j6HxP6drA8US/IrtWQ
CCV7AMu1UFSZXNILr0Q+SInY2oqlzlm4r07aFha1a4U7NMFaVYvNyBUJpBhEwT2s
M5S3DqNBPnJfe7ByOZxZ+umhG2umttB3eXoS69vw2z133ccvzt6dRrxbwZUsfdHC
b2A1h0qgG9ojUanntnXMyyqNAk/Hk1gujE2C74OUqNQEuwp/v05N4c4B9cnHu0hp
kAh6jclya57SyuXDquVqWGroWl2CkhKJt/5dEe99ZUAUdqdvywDHv1YcQBfzQlzc
tY5POkT/z9AAeMuGVyMBcXm6qdHsD7tRAvg516OHaH+76reYF4YuspZkf7owWdOV
CeU83Gaczkg2Hy0R+8yvliASpt1erHU+V9hG7hyCQkwDtNl6o3U62yAs0LW0r8zs
JilTqquA9Ds39MtftYu+HwpfPvrFl+i6q9V8CONWCj7/lycm7SiMe2ORzQzYve2t
LZEoXViOJKWBUVD3Ny+ozU5M++z9eq/EAhkNKuo5g1pA4aAS5LngAksDCKBc2fiS
ldNbqEp27JmGwzyfMkNHBuHCtn43ddE+GxAbVkLy1IxwOD/K32Ra81xc1gJQO82p
9u6rVewx78Ofgfh6Ve3ocCNd/tLN3T6NiLKrO1fi5A3ccCHUnoAhQtrcqY4JFq5I
nhx3SGa/l0wX4YDKYgjFZz+/Q40YKDlfx7R6Bzcrnkw1p5INFsqBGcZ1j06oel5x
aL5FQzWrVpYZgQoQS9IjB6m4MNXtl7qbePDCFEMSd4GFlAjx34qnh/AtLRu2WgAH
qTG1oKwwQsO0P9x+6BJ0HJwJLTtOa01Z+ZY4MqmYnpYUaSz/NjyjxlLgPGcJMEnO
2IGkP5PvW4IzzqaVUyErihIpzgRIoGgSr/PpzAgPnmxIXh6N9JS/0mc/gJhvUp0j
Mic7+pitc1u1HgIsBbZQhlIjPRW+4qod7Vg609P5oixZf6GaLeR88GuS9gasOck/
1RLF+qdJx9xu04Y/4s4zpx0PbGAp4v30IYCegkfzZhpPdiMJFKt8/kK1apJ2pkqJ
DuHv9cRyUjbAp6jzgRbYRhAqlDX/8+uz+Z168swmdAuT1ky+PRKUldBIedQCBX3u
3e/D6++Hn4BUoLlxf3N73gVFHMq5/U7YWYw54E00wmyySPDJfbOSkHU5q9Zr/ocd
2z7drlHI9CNeP8cCogjusdlf2gh2g6N08fCRm9HYkpZspDbjJiq4Xz+fKxz30mHC
hGMVlzvu893WsPZM/tfdwbkBBb5rGhVV90XUhtF6QlE5oizCI3wPePbuAClpU1fW
+7K4kkXuZxlX058mt3jTXEeBpPHJVB0vosQRFWNnSCuP9cmSz+3OZfnYlJzlFdc8
oD1eHeVRTnnBN6WGNaKm9QWBY+IBhIyInX93xGVi9yU4WYZDJIPhNWiIy4LAgelH
bTB//IjsUGIx7YwxAWOifOogv34sf4tTjKU/JiFi6huc/SL7wumQ93mT7CH0EXyl
C4hw53sZNiKm/vwvXh0ZsoM3ULI7d/T0z7ocb5QZP8b+BI3diAipmkaFEelrgBr2
E1EP6SyTPc1A8r7Ggadyk3ZsFgZ/B+bZ1G8HW+HfrCG+2gdhAGk3NX9koEdGIMqj
zNFc2bVhWLSuchoP2ktisu9m/p0041zmxaiW23dD2bDbJeirkQqMhSOrfhdLSWJJ
ugpr0u1iD5bAQ/s6gCuCfZsUTmgxDBIQLUFsX/EYcG7zC4m7cEspxMX3PGqWF5hA
kqbsiKa+4k10t09fUf/ZOyI60Rq9EvahgLLliVeR3HdmzE/bgMNNxY0G0Kh2c+XE
5n3sswUqKvb3NF9wWNbvi4HA1cgtc3kGtyO0ScfWXeDptMetNOcF6QQ89njjl4gN
5N51ReZxX8l/9W7FmZCSXAxbvnodPlCDcBpes/Bt0kTyHskbSnYl2tpC9KxGZpmg
IezMow5MNP7v4mtsnCN1BbYXmdVALX36+ArQUqDJsoXzdYRdHZUVuDuHpZC6lFfj
cRMsOyZfCbM59RNHzC/j7vOL0Io6FtW6ZD2JQGIvDKqo3Atk6ij+s3dU5xjcg01E
pWxYpbKstVdoid/JamQkASJr703+8n0fA0rG3X7a99dVlvzzfYy+IMEo/l2t/Bkk
u+3+7FChyDmgNWuy2M0Cy3xz9bSI0Cmzc30Keqemj0n+X/sR7/VxYjyqruD7cF3l
JhzVqpV1kOz7Z+m2WVk2vM0RN8IXJ6jz9PZ163eYGs3ZZvWh1KcJoOWN7Q8dW7Y5
ypqDyvfDc33JLVSFkgDWyCgNyFqa+s24wRpsFaZ+gU7Hrs2dJ9bCp5KiSZxHgZNW
2+1QADGksfELPvkVbWZZRLsIKOr0CCHlQZHNpaq8rqFUYnBazI24ASNlvkhSEfuP
MpF9rBAUtgvucUlMglMgrzXo/ExT8qQcb7KhIWxag3nUQeTQ5Fl//oZYXugYMiTp
84sUEbXUWCCiryiGnJ0Fwwsu7Wo6/o9ggxdD/KVamrIP/Rx5gaTV5oVCZEnszaji
mEW+V306ZMpFUND0RhU6rSsdyU6/M2HUdv3o8jlNaWw/jeJ9NW2G7+qbIQxF52AX
H9RaRjuZF+I1klushrmihg910D/9ChVc3+fO1CT272Hh4j4FDaAkn1Bf+3wtEl+p
ohvQCG0JvVE3XYwirCd3dvnYbAhh5JSrce0HgUHadNJgg9assyWnoSUB8BFz3Mit
hkjWPB0M19gBQ9RuJi9gyLMmRfZJJKuX45u76k2ND4F+UnRr5uMYkPfTXKsv2CZi
DSlTWTlnOKGcQsVl1zfQ54Mfe3v9fy3uoNLVE2tsSZedIm2yviGgFxbakHvIHhZ6
tQTNQk5z5iPLcG2D1vqst9CKQyvuITqhppe72vSV5ApNlGXwb5HQtxYhsGB46mic
Y+sFBLylM44JFlS2o07NuBG35LuZUPELZOoqScCLqoknZA4WAUrsN1IbdVFxeOxe
Xl/gOeDnONyLFrho1TtpctXUyJE/5RYhG4s9i9bcPFlBs3iwW0RugsSgbIC9khTo
az48EGPxeTOv++FAOPHbq2VgQ+YBWZnmztqkyTpJFDZ+RF1RhSCls/DsMhLbC5BT
SUcd0UHxs3AyQJF0LS5zBbl/R4cmNZ8TDCwpWPSpCZvhHaZR/dTNb5ZUpC9Kg9BS
ilfsbAinIkWyrC3z1M+/LFmFknF6hMson+CXSRD0Ow0ki6wRAzg17BgWlXtgMXTk
7V8IpfIt8N373PtjvfFJHLNh9573ANFqUxblj1Bqwe6uVbgaJnH+bvPG6tSybWNG
Yh7X5D2v5BbvbTVmok0cpZGo00EzoFzb+DdZjiSz3V4UTLwnRGcSO435WVLaUXpx
f+Ss6Y+RJbQb02CfZLnZdn7da0MYqWSYNOXcqvB/7l834l0cbZ1FR51h5K3EbexU
INBhxysTdtC0j1+U/OmB3nkNsL7k7eLnWmXfDwejKOGWrUgMCAz60HC5jXUKni3Z
xMsTviMwf6VW++bJ+G07VYV6OpvPgUmiCmZBQGRrWscmXzlCWoeIAd/XrhunNGIH
D3Q7ecKtecPJDL+ykNj8mxcy6mo7IrNoiv15uRTDpllhTrPjOFFxSutS4KxEopde
tP0yBaU9cgnK/cATO/kWNU5+9slsUp3sVEDibF+QDqDOuOrhIEyDPsxG2CLfK5+7
4wOKeVymKKA2gGsF0sMdhnI9pO3aFISG71bUdU7bUDKYVZyC6eytJAVwdSn42dJQ
LloND0O1hQVSpVTRhyQzwYIPfIf6u0r3fjacPl5wJDFcTuML6ETKqA7vqSr0Zh8G
ARpY/TsEDrUD5tubdffY+AKO6psaik7LX0V95jJq3wAvgfE727Apg5jSeDRjSP1L
bLV9at9Rcf7EYDrngJoz3r1OohZsvaF8TmBFT/A2HnFHil4ePfOi4cd1zxJLxWNN
Nuy4AK6U+9mG0TBMlHhT8CLyBAYz7mRylHZardJvypiLowhVDGYGuXiY8mClY50G
Ysuu5tVipEN99LKAfyh7XTa0BjpJalVcApbufUr38YbXZhlhYCV+2OvChHG26N84
1RMnd1r0Rs0n1wvV6MwhVBPUNrOi5ps/59RA1djbHcDwa4F3LahcBjIMx361gOYj
k58MX6G+xSDhUETEObvixegFmI0WffNys73aMyCM2+KryQIv5l3lreIyTC72IoZ6
EkUnh0g7NJLnWz8k5Um1M4yksF6eQpe8EIdGA3gUxVC37mqkhFnni3/2zvX6NusX
BpUyPtUpwTBPbycdYb8LYqhPoZCNJ3vYyhil2yTQkQu5uYsB2wezIrJcJ4D/QPiM
63QtyZdnU9ggkIS9bkCGNzCpP/h7gBlRlmmQo/ByuZG/kQ4+IGAll0Ego5ieo3oh
YPo0cB03LXJr1JKU9VWDclE5mIQHWrIXgaBRijKBmA/VmFvi+pG+I6ElASOoNvt2
oa7Kgcolh5eGmx2/SEZXohCwIHYQkZpAl6T2kdNXlmwJNz4JDSVzqVzjf8557IVx
sVQVsu5I+twhOsj/w1P50+C3HC2NP/p6Nb88aIXiPo06lLovdvFRqhxtuupWGW/r
g+99o7VbFc9LuApL7Xo7yKMMa/cApJvYD8NFILozFXJbTfUkXuLmWDzZQ3FyufCn
A6aBthGBSuywh6VCIdEIhMKdPWJDlB2kcvBFqTYvXiZfimh7kxbJ0aG21tDOWx70
SjyP8ywNYaSgpbkFg5rC+sYMVcuPmCmFMCO2KcPBqu/xPzh21lj+3BxdKgzHYzFg
PlSHifNf6zUfPYIZpsba2RXBgz0/k/51nAB64sA1U1L4QzKfGSOSw38XR4SpkG/2
6ruWP8DuCVXPswTIWOdW3LmGve0Cfp1vs5X5ET7bGy5dsXoHE8hXQs8n4i+OkEYL
yulFjGljPQZCRnptw/g+9RwYo0FxJNP2FTpZfr34RZvpg+Rc2/oRPJ+QdMUxc5Pe
EOFvZ3/K/p+iQWNwI7vGvBrwg7pYkOgxt3i+nc3LChfoo3Zay2CTz6pKFZDecefN
Czuqz1jj2+295xvuOkDAI4AYDYVc1/mGkSwnt3lQERHG13iFujdiML6KsZzgxRyK
Cz/MzttKvN8bBq9dEbCObJMNB2pcv8yawDgJOL9mDLLHJkRCJBUcfsa99CwK4hLY
GXkVx7WtxYOcrKW+0EQkPQoua9ugCmJ3LXOd463pdDMEguIJfLcO2ERhLNLMX2Ae
5bDfqlNH0C4BUnE2naOHMS6vVVTABm6iChY+kS0ffsieyMCFyzkZhbmK/qaYKWdq
1UJlWywDsjfANGL4f68LiE9iR2gQvm8YsAngjoP0cuvNEEcnU6qI3tBMi8PYcJ9j
1dDFycUEjc45Zysqv/ByVLojsX6KERgs8DDuI9zb0CJL/uGeLcaAPOyOFBufFU+w
3zFXGE1yz270+ODpIApSxiXixKQOnGt1K7Nam6Xg2n6IJXxAafinTnqpextWoMHe
XoaPzgKpujfi+HzWKT4MOAi3dRNdLDpRR9Wu5kZsgPlPqndH4/hxhrU5TPKnVKEz
D1Yq+ZBjTfzTG05fdMY5hEVeEIbO0IZ4JXiJwEo63Vonqqv9IDwExVnVLAiOSoLT
rfDuZlPyWmAzrei2vntt4dyJ7s7ZKJ+33kF1ofGb2Qp+NozzuV6JLvrvg8wKEZ60
oCHdABDIkhOa5MfgfzaoqvvIkRcLy7reSDmhugIzzmt7X2cbZdn5+x8xrcAp8FkR
zyzaAmD9dUBMFDYLP7NrFT/ALcoASftWkx32jZJY4LYl5k0yzwgKMvUpq3K49cGn
9afTZl/8nxKA/v0Av/ccjE2MafQe0oBUG6b4JkgEdvjFrRkLiaiDla+k2f72C/aZ
TDKUm2elyAwT2/oWr4UOtU68l9FeNZuNldduAG+1ol+w5F0bCWI8656D0TCbQpOv
a32KFzJ4WD9ozyUgI8fMQCwBUrMVcKcChqr9pQuJLo5Vy5zf+xY3qyGzoch57EwB
5i0RsePSSdqwW1hUYjYjXhDx+ZdBHQQVibj5CogAfqyHboNqnB5OE2oYzYk7Mygq
54sSvX6tRaUFwhVE11/dOX7crhWAe4TR0g0bmf6dTDmBZkqyfNQghGiE0zz9pbfR
3vTuSFlMx9AGifm7U5JD4bJLBPTEkPmWWfwDuBflBzwzd10skSg3Dcirgi2l/ok5
1f8E13AfC70WCUMyD1fpX02/15x6LSNpHMJ9NvFEFed5CmF+eb/qFf7iZi7vvsJh
MYQBB/utgUo3E7SCoeb6RKaxYnu4MXXDnTvu3jVCDWSTwQRPVTlEJZK7IwIWu2kw
vV3cnC9IzBfBzkJWSTU7kyXEn1ImL6PtaQY+bWfvIto+jg9tjWy3wrdjtEOq6dkK
lBtC8LzgeeMtwtNBC4KgzTlXQGfch3hy9RpWcg3osoyF/Dzz7/HFuawNTORmgj0J
gX2zP8mjoCA6fZkbdV5Fb2ylQqesRfypT/sbregaCbaA6xlub1hWXRD6NRVrproZ
fB5VAqYJvexdkDycvvEUO0m5QLCSSdRYhzH6Gs/gdFf7HXyJ6NhG4zoOEkFFlr4M
M3NiJWze8EAga2PY0Bf5g0iJZSOryA5G5pubds0jRRrKEKsJUuexsqDwWOYDnGkr
wh8MN+oYNwvef4ZVC2gwMzkZ/tWY57Qzckh9z5kBbEFcgbursCLzADrSKdjKMzww
CzT7+cE+yLFq+/U26YEYnJbBexhdvKuHIIcqQJKazH6ykj74wwxsjzs7KxpLunSN
x6o31w9c4B5wZNFH2zinaRUMuXMtdA9J3n496T6AB036wzqgfzgd4zvD5EFajxRF
vWwrUPx92rj8AxMtb6NgUpnBEBDBYSoR+xjG2r0D2NMuyu3TiE50UKSFHBlffJte
UEJLrQ9Mzy1CFzFaBFp8eZrqX73c14iR6WnmREw7kTEzhkJQjDflygMSVjrEaKkQ
hm2+HK1MjSQxEAV+MfqQWvV3uzySMb5iUpRG6AivcGSVQlrbc2NLa8UDhQSoSWT/
zkYH+NeWeFzpMSpZO7vPpagWjzefVszz2hUmsCh5CW9mOY9ercv1zGD5OebNGHpi
E9HcLNWTs0AI27ZSmoVX7A0+NaN7lW8lRxBPV/NyzTIvYwo0M/IS0k5oy83+sSWy
N+bz6GZ9p7CyS0pJ3STrmhz528x7BD2CmpLVCdmvzfbJ9mTER9hTtseIoGRsqba2
AatsX8mnUce1SybwocecNhPcLXlSgLorFg+P5cZfA2A/6Li9XjSM/0FD0XdS4SPe
FDSGOzrntMxNsToP5SfPnh/EiFZyn6pWIPfF2gwFQamKctBPsV2jmihtl57Y9XPu
8gBJOIdqbkj3X5+Vb4YdHj8kw48YC/Vs1VOrwl+fdU/s/EWu0VQD4K5u6UwiOwSx
SdaoVfyAu2KVt0Pa98VK7WVXcHmUF1RciRslOmBsyqp9MJM8zJkhIUOgC4N31Qdp
aPAQb/MSTVGdqOXh71dZ48qEnOCFqzoQ/8EpMfNjFpAxh5BQ+xmHvnJXz/ht+3OK
DnR/bFBv5B85jm/Vx6wFWKy1ZOHHsMqx5MOcGQ4hFvs9rvA9GOAwdF6OdCLW50oW
hRsV/GXw6nX15OYrAdl5qWN9ZQR1i4woIRtcQwaZywBu3sMV3d2H3mDR0ML5Viqt
g8v6CIdTPetYMMLZWUoqmUttUl5/xtKzKIwYTUc7sRPoLKyG1G6aaJEic8v9IBaU
VF3I0M5OiHvRlIhCKQ5N0riHhS3E5zlqQ82OBk6OOb+8voswEb4AWsnWcq6DlMZa
urAuHb10tG5JjnzGOPTHd0iDYII/BuzKMoIaG8/pyfM4ppharfyisvqpRrnMMJdL
DW2VaHyk8Uq3/YOTa55xrAkKteTVlHJkUliX2zdtK/bvgX/mepcJ3PWJdI5lR4Th
iAegVxkkrGHEcaHftIg1krqPF6Vi9aoH+XMv0R7nSPTTi7+jVJ3SHRJW3vLsbJs6
BmYPCjAmBeNSKX4KwSGLeUG2X1cMnr5J5AZ8YE3WFU6JIZSP1PzYdkSGQX6FGYfe
8gVIKBMkwRs6L1YXnpXXv1YDxBzJjCgGsaoWsgmMNg0bRHb0QOt9OOH0jzLYymnA
3BguY6856D175qqmqdqgh8Z5vdWiX2GmeIo1o6coKCDl37Blflf1ka9/PaI4ltXG
5bn9ZI1wJFBgphB2CeYi0G99j2Jmqz9mNdsGoISRWMFC3hvbYqOUSgR1AojisxXp
HPEi2S5Tcofz2rOfk6MpXwJR4eYvNz3PZiiCu+R012tLDkhA1iVKCTrmioWK3lsF
UcHFxPdXyp6WufeBOOtPqSCcpB31Ny1osqkIUG6bkNDPfUHw1DLZ2H/2aGzllmpb
kPZ1d52IU7nnum1L+DFaWUIZ6DVGMKiqu/sNg+cWyBmzIBE0aOuGx4rFJx4Op3q1
X/OKJ2GlrknHMIsNlsyR4ev8mnc1wJQcajjIIkyxNK7wch0Pl6ims6DPvFa/q617
sc/cxRNLiZllIcBoTzKiesR1lhqgfJOBbyNXhm0SpIfeHswt4omSNLAoMFU1+N11
Rez/HVOplxhYOp9UUWN9xDG+O7LEJl5YTcEzzYz3rFRQt4lowa5Bjt6nMou9+o+D
FhK8bUxObtmzQdxms0Fl2a5pUCSUlNxDpv9Gai0wsJPRlWU+2N3INAqXfkV3eam9
yCIyV8k9dauiquvd5E61unWwB/ou2iDpb8/3ffDX6s5Pu1Vn1w7z1Op6ADD7mjp1
rr8Ici1r45efUlhsjaIZmwwgruIYxArEVhYjYcl4GtVAwGH7bjhSIBGhMtPTwl/8
D3ArMaCW0YPUGxQ0FVwtToSHBBF37YJRnjKgJ9xTtXrR3X+PQflnQGUjlHjgZrg8
TxlOQIq8AzXY1I27ZWkbC/NqZYyb79jmLa1wGXAITuO37JqA/7ibR+dfwaG2zT6B
HuKVYSf4H4s/fIr5GLU2PbK500fUsWf1PWFWZsD0diy03qjp+GPrsu89tBkj3aXx
ohzKzk7Rpu+SK6x9QcoQjF5L8nQn3CNqFoiPpMBXcuYcTLxDOlJQIRsujlqudL2M
1xUnMSL9bGYLxFgPx8CTLD1I285O56amT19zJiSxaFIfTCzwveKZBl5cxLBBIDPn
ztvDbBS3UABYPOqLYhaUN9mDNzd65HqA7z1Zzc/k4prdeP4/25KX6efvhOUsNnEL
i9I5+y7f4b9K0Vgf4E5gsloDW/59MH7cCd3EZyAEXuDalMzoLWHHZk+OdcVwq4sM
TkrDu0hbb6GW6y8/xk7lumqnz00x2uIC64FyVH8FkznMplD+lw7+12JuNgbvqwim
qRR7euk6KRMPcHgp03xwDfoIe6LZS0Amh9eWgX/G5za5lWxJ6kbW+a4leifcAsGd
Yjeai9V2CRJqi3LuJGAd39orORAL5ogU17OPwedc6WOo+O06/UG3nQn0NhQsTOAI
jyfStGLBCEdKgDmiiT4NiSfYhP+Kx0B9ruXzbfQnvxVLvB3xO7cBGStmMY0w5rDt
B8B6ISszA6OCYz2yoCYiz8m6sUhtYZ994sCufrNPGI8c3NHjq92U5bsAvTlv2k23
j79vChi+2TJ3QQi1O+l9CHJp/S00Axhmwnf3qGAJk/YO4puWGxZCUU7uZhprUU+H
2zq6Nb4AUeyKXzXp6kpWyPfIQGutGRSQmZy3HeyBQk2AzEcij5F9aAjTxlDKANfo
mKyBDau8Hea3ZrrFD0lR7f6+bls3ab0I4EFlu1sIWDtijrTDR9yLwragS67LVeH9
rYyDUDDaUzrsmI8ZyvSIRM1/OSHf+0Ln3DfuNF7+0LRX8yFQy+9lA/kQjCvEJpdr
0ekzpcGRao6aRk7TvolTaMIiHEDlue+vUYExFgOCXHH9gHOypIVHy7Op9DOtWdCw
XYrjXMBqn5Gb3Eo6ckfH6DjtA6YhDHqS1D5nfDPbo4HL5Od2p6Z9xqXRyr1LgxqP
r8nwwyh1p6c4Gy4FXWaqNxf1tL/+x1VhZC8DVtDutmPoAJSkozjFVHK4n1NO6btI
H7+vzb5/WC6g1gBhn4Ze+QbIWXDdY87a7iFAiVvkTBSG8njd5zOr5DEqxOB24l8t
zX+0pm5KPI+Drnde1Dz+ekbJ5VBdoR0mFpPdpmgTdgT3eAOyxS5IzC3KdOWNpUmN
4snrmkrcbkd1ggsiFb1PxykfKpltosJWvzuXuCRCvMI4Ttt/EpyLkJnswH9YjeJV
MPzaEmCwdh82fqcOCvdzHH6okfyOePW0d9sJISL4mQr+Lp/PwYuJ1F4MD5se/9gL
iY6TvIyl2EJZJ//hda0zlwTa3lGMeYZNfRSDHrSTLgwgKqw44QmA9PAxkWVDk9rs
7g/JFq4GG2kqzySzt6nvaLTNIiafGLXWWdmtCQ9otlmRnOLFdAHKhOGqHJj9+WdV
GtGddc8f9lAjubs3Tf6WJ+REmIsK5hav3UKe9283YK2+Tvxo6/S4OWr6ECjRKIdW
R9PgsgL1ILMQ8eMacA0hk4x6aw0hJi1N1Lr906/R9gu22hR4j6qyXZbHgjgIvsua
KOoNTn3tRSST4QLHGArwSrPE5+4bevt+Bv5ByGwpveAsdzcPpaRjpGzCSQE1bnZH
1QVmu43tfGCDrwvKQwipmZtLLCkieXzJY05zI9gk0OQDzJVZ0GylQUjU6daHAS2o
oAxhCCuZgLNhqI3gvvJIGZdw3DeoA71veUMCgUj38mFdinovbN05xZvGGzYGgJsC
M+QVpuuFtAGo+0WhWM/GeJCmVFZhnMaSXUGTTFwIZUAE0N7R3/ZYXFylMZLoAzZQ
DTEby92jeX4KrVfT8wwf1HicllwQnj6cTUx/kmEp6U+RFpLpW8EYTvuxiN/ZYK8i
Z06JcTMgNkP++bgtq07mjhahXcmWEBAiCKGm3CrXI6aYqPEJdf0gYYVapXWiW070
MDxB59M4QZ5cb6SXM59q1La1y4WMq7COgY1HKj08X7wRDsRBhyGg79dsQbO/OAV1
GKZMYNDAClJumdRtPD5d4TtUPtkw0soTKJ5ApLLY99924ZBoRA3tHUrGSNFeHeNZ
EEoEqxpSH6ZBWKMyasTHf3PtMAkpDSQMXmLtuTpFPcnyDiyYLZoeYT7kr9yj08G6
nJv89s1MsrUvTBaqhxxZ9mClL2viMT3LH93g0C/u8xgRYycDbYmMhfxbjmD6HzmA
0OW1sFRUJuLw5aWnUPBLTHoFUFJBE7KnJULw9oncNdBrZ3XhetJzs7FZU7Yfdklt
+3LM2y1bqMf86RC65yqO0MaJ1TLy3JH2hTk7gFJ7419gG7aIh3K2LQl4USyLQSve
CI7SGX9QzbxruKaEsVIRPEYRKpkhagOkLczWG85M6QaUUL12RanZhjd/DRVZYJma
TnuHGsnlVCbwNJPahhGNfFTB3LQXOU7zRvX9w8WL4wuRf4PfmUDUQBZWwtJwVB/U
dByFJB1NTnii8He8brLJ0tvUfNUYmFe2J8DQl8agKRHvtXA1qXDirpJ+vKrG+yOK
SQoLXNfEnhmYezugIJI5wy9UCTDItipaeerGKJaYbPrix8M6l7B3r9vlCs1StWxe
sVztH1pusMx+/WesebFfuazZXgo69VNKUXmkalFAwCtlrKsh8SYQYUTAmxXogqql
Xm8DcBhr0EJBRidSqasaoNVdtb4sbRmA2szqTHppTZPeMxpOj7PkObAfevjBROBl
MQGD3xqtRk63cybMCmQawxFWTQYtuF2eLqPGFYaFqvldLxAeSHzyxzXyB3iqNOVE
dq6W8GhBUxC09NQik6HOueNAcl/HPd0kvWJa8OiV9kQmZGdETO89/Deuz0EEdJwV
/CvCYN15z+z1mvKSt9Y1X/QRHS3tgfG/TOXQgaVQHyjEYL3NuJImAfbzcGoC0Cmw
37GeAd9GL3uCA2dvh7uRMe8/QxHttU3WQvNUMit/MWpCvNuqYWj37arQDzKaMemd
rvdFdOM5cblBcRgoE4rRnv5v2xilYwPjA2SjV6b+4W3k0Ig7J8EzE/8wYH4S21qz
AJfJJRQATSaM9LX9SeFQc0G1nuPkj4/05e6PE/pFxKcsO6pkk8MhRI4iB59ddtJr
oXSUfSO5FFqph8IHozKV1AeqhjkvJEXNSdKYp8rEtSOV5gxd0JKL3gTeqmK0HVHj
0t+kbVGwFI6cpK682x5psGd4uqKsunqjUwapCNltq80fniHc155OEL7IwqN+zG69
4InbyEyWAyi9zt2/M5mtdYLypNJwdZWtVj11KH9zo5P7Zynr31M7x/J9L2TL71LP
3Dv763jDwebVUth2KuI+MbLtiUwNRE7faXkWgH5IPRdpp4clyID1HatOSayxI6rK
5Ly8Byanij+kJElI9iL7k3h63s/j6nMAWT/iNaGCZvjw6HXSb3Z/iG4IlvTo0HiP
V1o7DNl09pD5VeSM1bLyAumju1mBaDA+ZP/mrUfMp05uJCt3G75f2RZPODJBT+qI
KJwCpPehUd9LrlRhbxeQLRjzjvpCacR/gvq2+zefN2YzO3Ojud3hy36LqCFA70Ds
/bmowbmwFpLCmMq1mDbU3BpaO7YR5/lFs4T70HzEvSAA1wtjloWwyQ1jbPfkA2EW
1Rjzms2obZn3Zg6Esgz6BX5tUNjlseQKi5ijjrqqPdNjSXKopQ950MF3+wvtNgna
0ENa0vBB2kY+879UCRhITL8wt5coERPPDE11Y6HHj9tJk4NIqJUuPLF0M46nNdOk
HhEUrihtaWWS+jONSfkcLC6mZHM2q+HyhPyBQxwzIbgaXnXmeJxtotS9Xk8VPCLO
SJOmdnDKH5ICJG/bHH26eGb+httOL3c2edQFb/cHtOZ3tTG3qwMtRKhznvLyuh4h
dqunjbDF3MS8P8AIRAPAsPyQX8hfnWuWiyapvPgp0ibhlXJcenn3yH1kZNVYSOEw
ExSOzniLydM1K4mnuGKHiqWkOgXuGTicemxHYUnh6h+bs+pEtBjX6tz4AAnLS0LZ
g6UxTwd7LjjWqXUcrMEV4ZYvJTvS8RJIOJSZXSuF+5rAmeYlNhzNkdd+1rKeUoan
dWYtKKPI0g3cpvux9fhSo/T2XXj+GiZnon13z7XKCSs8EJqCmxqoEHQzG6PZEQ5l
sHBxkjSXpE1KnC5h53UoVnpzzHPaC1kO62GO11lhfmIGoXDfY2OHIRegpJy9Ae76
1JWJSZcCw5S73jRW+nTfkqJl4lvyGG7oBr4CoxOBlwtlCAL5SITHXtaemzTtJn5E
yD2wyg+ykD0BYaq2SDR2ZsTZc8x6meO/Tg31coJb/6L5ljKdBIJ8p6PgzTVIWW9z
HSPvR+reYbwsHvlFiialr8mCTSjCBslt9rc/Tz6/ItkTn0QMthXvhuD6MXprhNNq
J6ubS+xwQTu8ZF5YkQQGgMq0ktuJW46D4xDY47ZWe+9BAl3lIzTBNtjNxPmZMdl+
VMuZoXfcSs8X7bUi35fu/D+p7iWp9SyuxTEyF3cGgTC1O7pupgJYwR85XRni4gYy
FJiZtdhuE+ajvlsgqDl4vvdcUp8uAU2bGxc/l4sRueCtv9BNBhqtPPreO6JUFox+
ubCmtuQJkpqlOL5+21WjbtQgqT/JH3OwGXa7ztoD6mt5y4JaGHuP3TmI/eTnvWwW
XeGnU+o/DkD4ttL5023WfWobBrmSvrMHZuIyPF9iF/2wgYVadEWx0GORIAIvGaY2
9GvOjsd5o3UrmuzRW4/rIt/IzEmj3/x8mIhqMAYDipvdrF3fpqh8XWJ9FhJkahTM
045WL3QqoR7xcb3qavSOQCGQKNmLgZIungjF1gL6bIGH5b8b/ya+l0/nLsJk+Tei
r+NfBPHtCKYleSnGtMONew5qBhT1+yB7TjMcXVYk9D7/RKHMDpW4Hp7czGapgSu5
0Sk4wHabFDaLpA0jaBYujuTrGADH3d0VpJ3SLEy1IXCBfUvNhfyUaXhWYuNeix78
3bD3W/d4NgfBNA35RWKyeJq2a9YxwL+9z7kF/ckm74OVXWEmOYsO+tiPp208xBwG
tkL9L8yBBAPozLfLsoafL11hADEd92UuWubJlqbVAvmWXZvsku09cGDjn6rdWJtD
J+aChOlNIsxvO8uVIDYvqBZHjCIzSj9krVjUrY5v/H0UXLUVHmtlqV5IMhj7oqjp
YmNVMp9ELQom54PLTxAr65ef20huOWnr2WuJ9jUdnTAmoQ22yHBW60sIxi04FkK/
YsUWT07HPRgdSTJ5WEOJ3VXG3iIViW4Dvf6j2S5i3vuyS+tBW1AU+wlw7EAN5MfO
4LI7M5QuYNeTNT7ABUdh0O4tZNrBL+j30tkqeMnKNeRHmtXqDDH+GPB4Ay/FjQmQ
C9WN9F04OGGBl6SOPgFicG0T8kSacHLzDEtcBbjgooqyRMbAFQLyc58iff4/MtHg
r+uRJqmhoY7lIqA8p7X1h+bA8ghqW98CB/TAj7bRP1plCXbBdAgHl3ykEnEJ9dNC
IzZ2bntd2rDF91lQvwyUAO/9tqLBDb186Yi26+sAbEsIpQcVPm8/QKEzF1crsU00
zDlK2vwed5JJ4++ol7eFRcYj7hCmwGXalmLmVYj6UV4dk1HQaht2wV1NSGGihUds
tZ+dQAHZ3NiB7YkJJ/xY14EZM86fiwXJ8GfSNzC+fV7+Ilwg5ExKAPIrpcuuRh6n
/gKLEo5m/V9AGS8PZnFAsNe5q8t64QE5DR9kJKiABubeij+9N/QHXxLBNLe5HvuC
R/P3KdnDFmHJXHalmhZR8AX1AmudcuBLg9aO/j3aSmNFmZ88smaDAdwsc5D5Blc/
Bk7HtNmaLE2w6pKOSdP0ORhFrkigaOY1NTy39ViSptKvJjdS/3W4walSaBTEZ2mJ
7tEwt3dEfazT33S3Yd2A9fsyVVop9FKLHgKOkjR9hDwbElp27WiC1TpaUXG/GgvX
5BkZ98VBHpO8fEEG5nhqcZJavJX342SZBvpR5MndoyNdWaPWj41y22FF6U+CDcOh
P3HTZtlOJufTbGF8GtvbGvnJ/FQZHpY5dX93IZqs8cDZ/Nma3zrO4gxv4kpa3JIs
jpEWniW/m7joOlx/Ro625o4U1bXAeSXjyNe2bqD35G2p6372a+CWzMajW0n/yL7g
a3+pi/pYMyGpnY3yBCZscZd+osFLsiVPrxYF63ubS2OtkOsNcVXRcaXsC74kntFn
8QDUkG17yX3YLvac65Su5On4lvI6SPWXbQtch74XRDb9NT/iJLwTKedckoVLmtpa
Rlx6kGhAzXYp7HhZqBugH6EY+2tqCSZwjJN9zeC+TCa+uyXm+cAMkR+2JYq2+l4W
bbhsrpPpzkDucIsr8uiKF+Y0hTgkpsv3nef33K+vEOB7YxUm2vgRggHGHM0A+TEx
M3Tf7SiEjgQiB8yCX8b2Xpryo7Lh/Urtoty90pTTkQo/WBVe8K9/ynCWtBo8xsHO
q2vZX7+qSh1/KzqSLZk8thS0/On1pz6UJ1fThESC2FkNIBuqtQERWpLzNODYl4BR
iOoikJTxi4g+Z0EoZHkdrp9weEsTe0IeMhZECRw5EUXHvieTYCsw3e3XNlhOWlVC
QQLVJ7XJ2K4VIx5uhwITPU5pqaPtQ1dPBvQ/R6f5++vmn/zdAXvA4fK3v9+IoW55
ggU37prlFZZpwD3Z01JOvhyhQmjZ29fI6Pz9/2lmAgLG4xEZyGeV74EJTs70maQO
WwNPKxSX//DXK6omNDr9aV9Ds3bJ1I+ZjkpkhoUq1YDwzv0yTuhcyasconAnfdJK
1zhPHyshpk8jPEmE96trux6qnD1PiDUHlGQkh4wOD15h/XH0PjjBLlLyT9jqnctu
cN2YcMFtnq8/mEd7VB+A6ub/6hxacK9rvyyMjxHQA3a791RtCfnuLzD5nWKs3w4Y
T3u7iz2DfZ5iiVw4lst06/6BbP6EXmTsJCbHeXqxPlfI9WUrhq08SDcmj1hIRD7n
FTWiY3/uW9bCREI7/eWVbfDKgk8pCdSa8aYDor8NYm1q7eC1NhpT5ikCF5LHytNX
nRhctWS/QHt7nEEUXIBjtOYgG17mKiF/tIcq5x9tuLmilTKLCgV82uyz6QiKaXuF
Pi9pSdRnTSWOgG+U3Owz2ELiW5cL+OvdnxVz1GFkAKIyLWjxjbjtbIsNNIQYnN9O
t5tUTazpXRw07gfYFBMiQGhpDuSSVCwFjAMrMLtTe9PP8XYXtLg73Z7vD0PX9bJC
TO7XZ7FCKtG1ok4FDjr5lKvmXebNya2HTzIN9/2k3cXEWgwb6re/rZAve6LZ8Nq1
2P2JsbzmNWpCcpHrWlEAhhCU0HWTxirSrq+A/Y7yfdaxXnlwDy3hoguVX1USRjI5
+ajad17F6iBlAvO/KydlmUGXU1JohV8V4934gafqTSGGh/3StMGKmf1f1sSLKgUr
tMJIi1JV4dfZd/OkqkstvGAxVEFksvrlK6c4SqCHJiCZ1rghp4wa5UYciBARb12r
I9z5OAv9BNPZpB2jCnuxtbcDVQDm44pTSWizftaQ9odZZ3cTYbt/qu88V48ewwuy
D2gYvvnrT5+z2pg+jb4cx7vWSHQyNmAB92H0lE5aRq5nrcXYrp8O01QbgP/u+TV8
/YXyAytGhDphhmCdagplQb0pma4ytFVgB7pOLsGPuM8aaevYVw6xDaRxxzVMe/MX
Mnwgd0kbVPLFMNsHmVPpAs72DeZ6G5ATYLi5KTHuNtWmm6behesMqdEJTzXEcbTt
GRtSlfYU8Oheuuiin1Wpo+I6SHlBRITPE8HnWh1MpgV2Ac0/6Hue5vDgj7Z0xr55
fEMhrVQGT4XAJg8222xBlsj30pS2Cll1QNNHFI6iHjGR/12dS9HZwbwb9GDa7IaV
BxqGsQPC25i3nHgTiYHLS49bV+VWI7NWf+vuvL9sHT7ugGFP76AJvZb6hdLKiwKc
dzoBHZ23aeGIF+DQUIdPwZSTwqiStYdwzpKSxFxdN8cHXvpTyYPXsFcOMp3sp6du
MrciJ0OqsPHdjxkp+S3DOkCybfAwxAG46CgdHJHbf2WFQOp+i1v4/ir3MFWx08KJ
3zIe3aIatiAx+xkj/Z3hdKFLD6bbbhGF2RWypOLjzMEGhpV5YIAiz30RI7EVXbGa
eB0fEclSkrvph/etTDZTaSZ32m+JpoxqWKOIywS5vAHNtq7Q9OF0mDkWAJ/rwZNc
35QRh3BPH+UhUe/oCrnrP++WhHE6XhEOV8M7djtIsLeEilbuAZgjwcAwwGvbtRJx
94w1+AM6v/1Gc7XKybtcsBBc0EfXzFoekHGuSbq2iyTKdk3y+PGT3kiNTOmrP8BP
28EZ9WF3T/LhOj4rsU2/XoWgBzM6sTqhfuzpcROD5UnFGF45FJMALASufaIlk8Qh
QAxS79cndnEcaDDoFiK3w1zg1gvuSH6xuPTooWwAEHCz2LL1jbv5WtrQGDrBPuye
2wBreK99PUmjni5pRn/dErb48qMz7wJ+v/5MBeapnscv5B3VNEHN95n6OE9jCL6L
KKSpDma2wdEscbJJmC+syAHijXWJOvjhRXgmFy4oXN4URMcr5CKTQer771LIfdca
YbPI8SCCvKeqqrjssCqOAqTWexUhMm9D99ACKu6innPUUVNKalVL6kP9FgtyNrUz
J4wyMMXiUc7gvJVpn/UGw0bxzBOrBRQkqpKBubxHHjHgF3lQMmICKNAP2Z+rHNU5
fD8WzAqUQSLzjrkJqv2JWDEqY8uzyoPLyauNEalDzP8D3IMBCEoQRXk3tcGHXW6a
6fjbmiuxwPOKZf4W+g5bgU5jUPQTkH3jnRFtUoom5+miwCcNY5bFGjHLBLI2i/jC
5LrtUUa0DymjwkuQbyn9uRbspownVK4LOSVdz5Us2GsSKzjADvJ9jh4XICkBFxdX
q8T1ms5yzTVAPmIAZ+xDGgIkN6txBwfko/1t5frCniBwjKrlG7uRch5GzfetXu8z
z3FW+goUr8a4TeGeyCgG/hTa55hRjcOEz8mYF0i6gHEzVLhJJVNQT0XbUBNBleJy
HiOZYhjRAetf+CUiWCwuYMzH9xcXMRJc5/ETh9aGtH1uK4KespoWa8MCQcjBDzPJ
+4ve5/rJ/nqFD0oLKWeU8XYa3cFF8ubJPEZPnpUOH3pTefStuwHmcU/Q5mBOmRK1
mqY8yJaZTqLp9FbKRRdWifovv13QIVCkgad7KOSj4u3g49Zx//RDYePJQMxj3JyW
2zP80EhFjSmnWfoy9LSaM0qwckaKvBKjffXx3Lpm4B2oa2hZWmHfzpOxJUCIRMoN
ErjDYkXfPOI97T4JVOf6QCk0CompfgcKWus1kU/ZPGmEOdPKVURM44zxTJyq4msH
mJZs8lXMPunLKYLmGN5PikP2of0KvlfIrWEQ96LV8NOeCsbE0UwVV9FJ3hWbKMXK
a/JEEe0QGlTBqeMWkhvVM69gEzZ+7k1+kPSGLAQf6TPlgC35H6V3+jlioXHwk3ih
Gn+V3i1yc7XE+yooEVKTk33aSU8hfDbzLCiMlxBfV2+L7RcufESHPOdSUWbb2ATI
55z0wlsaalOBLNLbUdFj6cEJPpkYz2LZWlHhmV1O5VwZrillXI6lsKcBK38fJfHW
zYS1GeBkg8QOtMzw3GnKE3KBw5US7uxGTZqQ/PBFGBjRSeYmMj3wpqhCDXNSyPB2
MhzcgvCif/k65LX+ZGq9WCppwHAzaYGt5tuflkW34kCEWdTUqcMFXVBbN7YoSVce
DbnDmJ5Kt1Y5njCndgawT3bBgQl0iyFJnoiT+EHXyqzreLSlBDERwaxJtVhc2jaq
PZG6f3ZNH4Pe+DxQwJl3g57U3bBSuQanuOmITKQglBlMmNSK8Dp968E4HGvn2O88
nWLDkzF0eAVRK4pJzENDHp45Qm2D6STg41yMUENLL/VVdYIuHXa4ZCHrFrqfOUDM
9zCYoTqVoULhp+v2j5Mt7Ibx2AfJcXExRHCUIb1ZwcMbBDT8b5PIpmt9QMRF1LXv
HaD8MKpmDndWaGZIJENC++erXsZMXOpnly/peVBsCQykJKcK9LLzZtYrAZiThgap
jPe7UwfjXCy3wONFwVzr/IJMBawQOJZeOK3Kw9EVtSnEWKXmJBECTy4Q61oTmSzn
rN8zJxCkHHkmI+dWf+oaqss8p/1ooWVEejX387tmD35WDu5TW5AhK3F2CcuYMxqH
Imny+lCEQG+gUnzuZQvx2auD7rIT7llxbtH5J5/AdGNBzpNLihPPYGoplfSf+wFf
5/FOR3zXCcHyN7a9F+MrSKG+123ZLR7kK5ubAbj1pxIrXYKotZ8cOCX6k6iQXs70
ma1pGkUeIIqeflyLcXh658vSaJIF5Ai3AJf8NH/5VjIY55y/ZdharrBtRMbNzjyl
emgpeIMkd/v3O3COwJUQ91lS8EsGLwShLrR0Tr2Xy3bE8FzF0sadWCT+szIrcBos
qlssPFjetUrggxSBRQPrakzk/ZDq6cmac3oCR7ifWADQJBL1I+ql3Z5bIIZMXCkO
FCSFT+rPAI7rOzdpmH0XU20VdQW4WZuA6GMZcr/lPPuAGyCFJ37R7F+8fVWZkTTf
ucAtYQSGTc/ixWgcxuzXFw15zmkZ6/SSLDIBkABv/2Bzm9kEMmmVqm3qiBdn+Mc3
uvV92ngbpkEELK7QV+42U4s6Vo1my5uOqlMCcNmCk1b4iz/pPMB61SLAloKzlOdT
5YE10o3ZRoweqiWyRvEH1NKj/yTgkcCGQ6D8ob3S1/KwRFk0tXG1/Zy1bTq9l4Hq
6hJRQviGAB/ouHRp+m5uiivYG9B9Fq5vYsBqOHR2Nq4j7CWijUFEWhDz3VogYM7F
O21Gra27YOBtxDFkmW9LN/uQHTio5uw213hI0o8MUlf7Iq1YRiF5gKTinimXMmHP
HRPQJLbULxDVRzI59k2+rpzJ8HhMrEGpXSbuMClDO9kbwH+UnC7G/ISc8gfWLzs8
x3AGxqZbji9i+L4MezLd2U2kC3zKkL8EoKPQNf8U7KuKYSR660sX1b5hmPUjrrfJ
8++OLDoS3RKWnrVjm40bmqllE50nSaWZ6m17BXvUCu2VxuUipJs6rf4/FKUtTvcg
Y1wd4TRLU7lQDOHMDyxobsfVbit69Kn52eijKqC/9OolUGUHB06ysi5SSIHJZbw3
Da1oUoPENZKbaDNtVh8vckqcUhKel+rpMT2uKlqVvK6cqSuM8GxmNDta5lD4jdEY
tHnAF5nG9PaCywkzeaaTHnlyWA4FsW7gaUXV5PPYL42QurB1O9VfY4FcOCOjEEa+
kfaf0l1KvWYfdTCoPqVWE5xGyQILpRg3HkoBdQKrkijYTWpa21RTZgNScyG1QqTx
Z0wkfXsBBPonBCUvd55ZUYcV9y8vYCD40SVHQrF2NhIDiBCAZFzzbvzFmZo/85GN
Z+GRuEv5iBr7aRrL46eObwAnk0uoih5g4xkLODwLaE1EOfmbILgXXAJLeBxby6av
KUDu3GFN6wZl5BlBBkfemMYix+KRHFTktTS1E9Tj+zGT2IgHQk1YgKIFsMgx1GWm
K5cpCSxhQgECLG/+98teJpXRMk/GsgrOfxiDGOsrZrgUsXY63IIEapMgMJuWT9lv
Rnd3F8j31vTFUCe9eFiQIIhMGyaBwYCJQPkbxi21zu5JidhhFVfN7R9xEUsm7s6d
j8u+XgylJloS//HyRQSEK/E9swqgfGeu4D+W6ZTDhpyfzEdq1IWMKrDypyHC89Z0
eXTAdP709mY43qqMbqgjCDCPKv97mOoC7TpKQ97TNbWPBIxzKig53k6ePfJb1aUG
2KgXZhrl8f4DtnYy5YKRS/JrVjEf42W3dpyiK4qdWuub4Szpnac+VySxePNeWFXE
1wK2jfiHw2pSEcaI8/sz5K1eJ53VJWkF8lVW8/MH0SxCQcclqn/iMQ1F1UsscUDR
/3YghyctNzfXXxoPX9bhK9Zibphb3IAGutO42hF/Hx6CG9fcfPSXVyVqxENPgbPq
Q/OKNwZjZYwlEhMjUzJWqvWEun94caNnK8im+edC1mHzXYt7wJwYvIelrqU0up3A
cNrxH9gXKgMwjn2f4Rj5YCyq+BunR47v+amBPjuTcLN8/fbIAD1fm4XJ7muZxVJA
dlQ0LNKw98obpHBUwZl7GsLXbXTBDiddsRcYZm1z2dovL0ros1876V3akcgETB6G
ZlWz2DLSTvO6MwYPH4uYtYM4Cvp2SNtqZNMuQAV7jhQwYPJpf/YocRZI3U3Yrd6g
6m92ppOFSzTXz75A3t79Ar+GU8jscCs/Mrfn7xFsrZRADxpaHtd2I26uyvXT/tIP
sFkNt9gUuVmEyWKyqm1qwsSA6HXi40kalA55s2+tvto01TGpjDO7K4jEyZcXCKBP
GFsgZtI37TFblodn/+EpvgKFJGNbDsTyQMFz1+VmbiF09YV/iNlu/os404p3lRHx
TgkVe5WzEKX+SESKReOf7Ghb/72CuWJv1V39wagzWAukfdTN/Is4J6AAaCV2e18Z
fiN5fXaBZUzenFEVMYaRSkRWTpa2nTeNwiy+RmT9AS6LDpNezZtYuiA8Zyb+pFc/
7CUoc84aCXg2XltYBPF36admkwNp9Lv9Z39KHpfwLh+dH0ThPATxVyqC/WYjlyxu
vTfa2zw29GPlvDEn4yV9cGF0x5AVkAMIR/U6sP+8NHQ/vrR1Ed0avlU+rxUbtZd4
Wk6yxPWQ4ZGoUt1BnMXrlOC32Zkwhg5sre2Kzu7jceIhcQMeiReTiLm/4HUoqNLz
c/ODketFYTqsr8UA8wFUKPDhxNrjOtWNZwmPdPRidZfEWCT9+Wkpt8nap2CvC92/
wtIDdyw3LbjbABnl6DgtteSwI7VpaUjDwdZP3gvtK3IaeNc4QjkZmbRyPtiWzfRa
Bei3+ieVZMaywSYEfaJjC0wBV/dOpdZe8vC44OyKRkZVW3ZcsF7FpMD2E/BF6S9U
lgmNJWP/pEPWc61CSHO4U4sS2UPG6mtBWpxvimK5M47kzi8awNO8ihf6qbEV5hYw
EW0vicQ+LzlSga0Ke3wqQmqwXuP3olVeqpzK75MieDfuPpI6UMgRaZoGuBt8rgk0
ENrFLAqH4r9gLJuP1qS2WDSuG2ToNVzzXKba8vKNJ5plPFk0Tn+mIksPInYgaMDj
91hAlP0Ri9MPETPw7G0VNXM/ZioAzHvTzKTjBPxy6FyfIhRcXgXpCDM+KZ4h3rlQ
GXgc7SilvNMJzgcNyouF8knmjqDe6bY2UrR5rP/v4f0NfRa5HAzdnRxgRD+LH0N6
KBwPW/dPLpbbAyzbkfvF92V1eIsDiavJxW1iJkQ4uBMwMEB2YuakFTWSa8GdaT/A
xNcNYke50J2U/DfFSbYchqWuT5f2CZuEy+iZcadaqh8+FJBfXsESNMLx0/ZSTA28
zy1rWw1F1NP21yw2iYCdrZO/CBD9psLLk8yXJpu8PpyfdSkYHxoM3/bEU9OByJTV
VmTTf18E1kvQDIbn75mFAz/XXfa8/0Eg0t06w3LyLSVJsGqgq0+DmZXXuueZErrx
MIWPcGizwmy8rnO7GBPoSzcA1qPJk28RvjsjCo3sHnHf9KLoS2TzJ9GzLMBA9Qtt
RGX6La1O/X38k4gq1rKjbI49FXNGQ/yaiqEiMKJZxqCcw4pVUVsoSXKGxSq6dwBw
Id4FGAV9ywQN8HDwryrYjgAQ5DhUB6b98xqmFs0trREI9czdTU0eQ9M2pTlIymYe
0db4Le6+XOECoBKzTQpbobUl14rV7zGzm9iMVkru2KbL09f9Iog9/tY+k46CBspq
b1izATAT9f0SfnEg9faz1ZvaUrwMGH0fNqfs0fnFjZC1t0wx67st81LvX65hkkT1
AbqXtQIaTuiWl3Z49qLbD8sPpMy9cwIczzOVwhtlohZpmQs/FFvGykhHs3fMBqA0
aDEX9x12mhXAzAycPB61dzRjhvQFP6Y1xfWHh9F71i/yywUDTzjTfEIbc9fOTDHZ
NMe5EXwYQLatuEqKtXsmLQ+rzWLr1U8Pj2Y+7Ui7ndMR4y7SOzKD0DGj7FJcNpa6
xNCJFD+zSrTSl72Oh+K5OZNts/QNUtpz6ePk2+B512R7wdUeu8GtpO2s+iW1aWf8
3tBY6+0fcqCQXlcrLcGgxZcr87h+RfQPEY2ATwcFuYEAj3+30KgSeh7ASjgbXzbA
RGXw3JZH5EdqUNMjOQnqXoY+eJC7/EXWPoBgnjDMuHOIxVRXmuVSLAm+oLmz8oxS
GnG++0F+pHoyxOsORHvw30K/Wb9TxcS30SnjyhT2OpmuLjyJ0d91OTatpONm1WMH
Ivh3rR/67w3m70nrLnB4UvC6NG3iGx1BSmQSuv1aJhy7b6DE2gN6xlMefEnnxsBr
QK6gvd4MRTciJe62hnMpA9DhjWFlb54D7PXGW7DtTYANUutTuV1gqXyFKreuQc3v
04IO7pSxJ0jsNR/z1Mk9pHkuq2nqlKdMRUqVCRCuAcwtKcQoC8wchBnC29Fn6w2L
gpdXhOjcrKe0KMlNl+21kjTjYAuzy7x7K0C8N/D1dFXCjFph0c9BppCVYc8at+dL
zoahJEqMDtTy0QDM5wjwFET0Rx81vBsC1EBjlTEgftSqRq68JdmEcVJy9QlfDeUT
NVgbxvs4pXYvC3KxoznrIwDMz81FuYWOnaKAjLf9GCOX+Sj3MoD4kFhZjxH87ULO
1ymK1gifX+3uvE5p5MqSMG4YQlDdsbEJ3Fc88VdNirHHnYi9JvxZtXTxu18fTHZz
6d/2y4Ja35p1ITvs8pYTRF8PYX5j2zLmIP6aQMlmAb0cXsB5uwZtjCtlQsKwpwUF
XSQ+tj1gk0kkw7SWmVtDekGBoXTerGZDhdOSkDoB7FUTaK80vqSgw1niggTG/NaS
5pb3tYLCtSl7CuIyPHrgrcHXNGWw7EkuAOm7QWN6WUVlHtF/efuEMTypXAj2znXb
/XW7jMJGlybZVNc3LHr7xPOO5sztORbcHqQEe0aPckzMlb9xdWcLqvWG1tiGEc17
XkUk1KX3S24RigvB0LB64F+tuYLTgqzNfvEXa+3b8rmxHJWTnZqQll4hSeDCBWVJ
NpsKhjY8dfvh4YB2NLciLOc86k0lJBZtlITpyFut8CxaBE4He6mZneZveB01l7r2
LFTGM2LbFhj4bSXphO0xBa+QjrUwMHMzZPOWbiTg9twqTW9rRqo5fE0CEHARB0E3
XNdwBc6jbh2nYRr6eJzEBWIDKrV8mbk0KJT7dlHGjptwn180gHbMZKhSasJdAnty
2BZ1UnO3OJNri5bHcGJJ8W4JQm/XkOqPq7QoCpeIcIykbP3PLCO0sMtRSCL8OsE5
eGTOq12LgPRYAY8S77vJDeeuvqLxv3j6tE/YegIvVCYpv9WKTNrjKQp1aY9dl+hr
pNJgdUsyAAWFgX88LYUo7sPMQ9WZQGtXcSL1dAVT75/P8ZGsnBKamivaIbtY+r4G
YBVNSRNF6VavvMeQcOMUTpdq3WLx06mVx4+scU5BKwZBEmVqVOjBoW01BjQdvzhF
Glxl4296oOoAYw+tk3w9rC2AZVdT9LHElPgMKfUPSB+a5nuOsoFchp3C5wPYws6C
HuFMSWBH1U6w5s2AyoRmgbnqYsEkMJGtt+7Mcgu1y6JUwVD6s1D1cWPUoPZpqqTs
6qKGWExeBSPez90HAFSWyvd08ABPkvmCcYHuxCP3/JiMoZo72UmVhQwo5bXc/so4
XV12OBBF/3CCJDg6qdXODTMAbdco75F/9oAVhZ+/uj+sB8BzoaSNVpeyn/VuAysF
mGnG+PVDC95Yrs+NrDnbC0i15HWkXV7sx6wZAMURdqvioBguJ/opyC0qTTerUY5P
Hk4xr07M0/9xkWnsg1eZ9fAPtn42qBWJTPH54lMYRjuVek79PGn9KWuBnKOdDYhu
NcdEHVyTDmRWBE9Yefsjc+jHEYHi8xRW1buwH6/KsFUiG+rHG+iCLvm4I7zBuUNX
BD3GOrwIoLjHAmyYd5vyfnDHou5VT4wO4yqV1KxfQ72yalsw73dFM2QO8TqqRe+g
hOJYcY3JVFg94DVI9MzEKKNc49lPekTeRIzlBN0mOLYGknZMHySSjfHUJZXxuOwW
vi88EI6FEmcQSyXdlLggcEABDMjkAg4adY1X24Kce8D+TiXaSBnwJWPGZaO2jKeW
6pAwiAi2aUmwY2u3OLIFwuUpuxzeKZuSx7wUWCt/qltvIDhNn3ajKON66mWhwnID
btvAU2z0YGIKRJCzvpG1sJ6NFGy2OFxrxXk+zAldsle1ZJOgnR2uufEsjl4dvFse
D8EjuJgTMKQRheQI458OChPor9ovePcqaK7DejTu/h1OQQJ2fJzJqvIqS8aq/qlF
ojhvkShHhsPN7aI5fEZykmMfFt3GIsUBjk6E7bCbTHZv3ELCC7Ii/PCwlnIWzFeg
TIfTCwMltbpxlEeW5n3RLgnUWJa0L8NbXFRD1ltVvJpQHAMWeIxHGrPa157gidJe
lBJIx2eiDk0M6zbWNkOH31B+DD0pGzCHumiOJiieFPyYCV8bHX6/M4iY18Hv48AF
IpUEk7V7D3tCqVibJH43yPsCbWqy82ySTpQhGvdp6srnAdHut31ADPQz67OwMhJM
8nXaM5MWLKpI5a29ThZ9/KasiNZb4yv11hxfPJsSWrjJK8nMy3DuF0lf2vwnoUnX
mK8ifuVUlb4F2wrXAhrbnt90OvkGqgbOOKSOTT18zFXWp95tPCxYPLTsjmVvm0QE
Z1vjBrK7CUmithgqVyykdWYfRijdh4eS8UCAasppNcRBrPVYEHXxX+nQEsPti9V7
qtFNvA1Ud+kz0lBdPFmhKwHNM8zqdQlCVM9Gif4SBmzNaJmD0vUDJlwwCnE58i1H
FtbviOeKnLTGdXamiel1hARhBtN7Gr/crCYRGg95+/bM13NoBNmfltrLmkJFY9d+
mBtbWPdh5jQ3BGZqlz7PwM9R0Dmpk1XFsuvXlLHdLC54UYEkdciB9Ue8yjNHa4Rl
nCkt696WhzcXyEheuUppBBObVT+YUbQ+5SoE3ddmkcMcrNOCmfBymhA38yWSK2ig
hnQTceS7nrMkNwJJFw6igA+Ou35ZWZw6w4US+KKOzhwQhxEEbHwY1IpcwFYRm8oT
qz/Uz84CPQZMQkNsWQ2WK3LnlnkrGn2IA5/49RAlw/53NZG21KQY7rUmOnvt8P89
+X9SzSxpF7a0/Cfujby6Pdh0tBes2TsuDgTGZBkEaoAknwqs4s1eKhoFDRtnkhkO
gdCX2PflHLpMPfGWtSnhGSqyKRlUv6SdiKdvWJgTMhRBHsto827JUsR/1AKiW0Wo
YlJYsKOppza0pJVrJJIUOg1Cu+1tt4gXmLQhuk8a/qDvuYDL2AIVLr6FUPL6dwgB
8v6Sadz8RbeJXCrcKn0xnDQB4ed4R6QJiatWxCjXQX4Flhi2Caos/nv96Ozs4YTb
7A9X8p3915vbDhmtbzCPJdzmW60LngUJm9/SjbBD79iTF0ZJH/xc5HTC5+rlaUu5
IAiyv6dB4lZjY51GcZfCzexJpC50you/7NXhVrJVg+DiKej+ls3odjQ9E66xhm1i
nHKX7J1FDRCYzpoivAacQgtKHHiqxVmW+fbO9iWH4Y3XnCVkfDeUGV9yHmLQe2Yj
OzU8LCSOJwm4iwni9uuJEan2B7Lzvnj/sHPELw82w6oQ/deompxScIFUGZ6aIgNf
8W3eq6tvkZb4IPcuuAiJ6ibN1Gk9VPU1vmkjwTN86tIjQ2b1ZQKP9V8Mgjh9TlDZ
G0YN8d/SIa6PcXLpXkxNpdpnxjieBycv48gbu0zEkz+f3jdijMWIUxNG/2HPNpg4
OvksywgSUJKtg72q/yJVsR2FQx4cI0LE8YaEzPfW83QuU4rIZaOQzTYNuEos21Mq
VSteFGrq0ctSLjGOutBWYGu0WFjR+HQpxRrjf9MMgFvXPsnAqlt8hMftghyqmc7+
tI2eN7liQ6PS8T/jSG4OjlCPGK+WAnqd+p/nwUy73VMGIbmWer15Vwhs6PCPX8T2
54/+5jfYbl693RA/d2v1M4k5/gJwSs+bIzi8ohbBTLH/V/znr5TOyBWVy071y8pu
tskpT8a4m8akjtZkEMM+QPBYksSnj7G6J1sOziBn7hShvxT+BK9/1JeA7aRYEU6o
u3uBLiwsVZO9QgIiqItPvochyEUlnwPEaFhf2q58KtWQ3iBnvJW8m+gqnW1f40qk
hOipqj5iETcP9nHRb1fPTYPzuMhq2l12kqiNuEF3JKvAlaGfQ/YPqQ5Hx1RAXs4p
3ywHN3nqQVZGqwnvOk75S5qfHo+9b8IlMHlHInPZGm8rhWWIA7xVSY0NUPkWbz/B
qyyHXjbnxwhaBKqB6TyCwpNLvG2aK90SLRVkqiNgLknWRFNgP5LLJSesliaKaNbt
oGUMPXvz1+cSAxJF/Ato4KXWNAMUaa9dlvn+LLfX0Ho7+AL1WzU1eMdvBFaMC2mb
yVZg/tko12DRfo/xKGeuLtz1pGMC7cEwT30NEwDHnVsvu9Lsd4GdCpGP/seNH/SS
wwkQ5vGsTGCDekACPEQTrCPzQqNu412XoF+1PnplPyRoj6GWVAT2dTILq+S3EKWN
+me+1Ynkyu20r0hmqcZqc03WEHn6PdnC5SPx2AxAFfIV4PtyEX41r6ZVNVrhk1wj
MTdeXV4a5B2V32e4SICgGFWOOPKMWN/sbRCh4H3nk0pVmbOoaXxaHb29X9mv86N9
xiYiAOjdDHnE2/igEznG/e9osGR0bHDOnyMoUz0sBNPqmM06ocHa47OXFTzLPdoT
dnnKbUglvrSvWYpZzdiBjeibUjJF2/GRG/kze2E/O0Oo9I+WoxpAe0lEFYE+JMMw
7NO27xHkEpti9QH62USlbg/7Gy59DBnD/pQwQukeUTNa0WNAvjBogzJyUx9er5dv
8Rsaj4gzp3A8GiInpA4Z+/V0Xg81I37JUv1KnlpoHAY78AU2GKHcZa11RIYcH1vr
RAgCDqeZBUMXJ68KiO2eHMOqBRQPSRzyinR+IoZU/sVDzHWE/br3yH3T/p8uzxlK
IWFr0wtNKzShCh8pUDK4H51MdLI9Y5n3159tWxMFRRc7BrIc69yJw5AVBBm4LcBF
zI56uDu7vHq1nMS3EQ3xyY9JoJkpmoQhsBpm73BA53PIWVs+gbWheE6+fyyMK/b1
4m7fsMrLJt8Yby7F4KvNz6YXlY6/7qC/aJL5K1BLNidslQH5mkBQmYyOOHHkqnnj
02BPXCDCNnxrAhqtiosQMEppuYY8Kdrui0jV4IeEwvrKjEFGGUDKgTQZi5OHPnpE
o6O2BHyc0ZxNCIaQbuuoauCVsWBgqLHEhjmWhAOvf0HxtQ2iGfDrCiIrdri4sL35
1u4wQliU21RClNVhC+iaLyKImoQhrsjefh7JTy1vB4Wz3yRb9n1KxFbpajTznNfi
y7U2uCeNO+GtRSTYv0scS+s6UN42xuLQMostCU3De3SkwxPar8q2Zlu0xHSG64f0
HTShn4ocOOi9vljzyy1zylYZM20Aqs87khM7npBAEEFQRazaoARQEdSWS5P1jqi+
ec+8/PxjGQE3n+YioMEF+hFurXWOHYUvMesWEwivdqk0y1uRykCjyxz/5kSFQnax
IeyDFWCXUNj5S0txR+608AOJDWxx44/0cr+uYPBRTPuzpq4EzqgWQ8AyYWeffSrV
VNCSpFp2CVTpqVazRFGLBjjvAzy/G/uzUFt0EiU/F1E02qOCS9POknfS6HLgiOQa
J4xeku5JJidmX7l5TOH9kFN+gqF89sFfGFAuR+oWQw7HnN09B5sCUsQzSeWov9Rw
cMIDXWQKDkTovqpp2SBujsDj7nhXBMG6UVZRmWKmYZCNd71sDWFuluCWH7tnaLOQ
AtviX+3FKjxDo7iagdJlZOrrevoPClUVI8R9rRz9OPf4+GZzZcigrAWCbG0RgWDz
e+TeLazc0Md2vqErs4gOUQjvRNUUAFDCzF9UM5Z30GZ0w+QNCD/FQUgLFPv3YsOL
uzdbvLZ5T/GKk4+Jl0pRKVQx2FrqoYDgn1ZdhOWkL+YtK4/cBm1bRoxopO5vJ5ho
3xD8ynu1/QIF2C23Pn7YCVPQ+Uoy1WcL4QgblT2zh9530hhU3eB+jfs716CnWI1f
7czOcMAFrCn/zCSNtH6uxBMVAJt/8Tnp44R5Y/kSfWIrXh/u5qmC0k7LjEdxiIY0
TGPNbVQOjyzarFb3DJ9TnrBv7rzdOda7RyUrHYoyJrM39s0v8tc/u6zdBT2iD2tn
ukmeEwZGtub/sgl/Mk57nwBtc12KX4hCHkt5g1KJ3yPTxIeo/FplP6w6EdA9N3ez
7vLJyKDM8yre66Aogq2S3Kus2X2QhivGDftbABWnJaztr1rxQmpyBw6tyujj1KXC
74DcppIML2zGJ9R/PtW0IkUWm223d9cF0rMuGHICzLpKcJqWijg+4kKbjiMc5DbU
Bgo5oy2VOs1S8hO/0VQJtwahfQtjFQVfiHF7jte6RzCQbef6Z09l02PQB5EbthHa
74HsPZRxctPCIGvM1IdfMRfUE78E5Cp4+5yfImK2e4GtbATFtbduzW97Vrpls6b8
J7C9h+KYVhriGpfzfQZB8Kczl+N6HngUF5liKht+jYTGSuPSDrh/QcUzxzNc6pOE
ocC8Ss/jBQ45JgQ3xdjqL8f9xKzycFZxuvYS89pxpt6VV5jiKFOS/w7FlZpSufzW
ZxKp/jEwC0pnrVQmWiwrDc6smcHDjYhTe7+Dt/G/iRNStw9jmyQnTDTwbPafM7Z8
I4Wr/mOwKSQ+Yv/W0jvtP8ih5FjLuaNr+seChK0Jbbo6//ITzOF5qGLt4qkcLaK5
y2j5Wmh5jhbPqvRAwntEuDsnfBte6tTRt4JwQuupdf+ONVmkP0DTJ6jdMjwIfbGs
5cjqXEYFxYN2o0q1KqkLH4p6gnBpihAGTM7xZ9REYhbRzYlZo7xmsdt2mLUZIn1l
JZQa1D8L6iZcTWUDJN7qkQQNrYJvv36UBA2HnL6706CMgOQ8JJ/8wvY/oJvlyADm
MNAbt/14ZiyStswDAv5sBQHSii2LIPiAv6WdfSrCVVjvOvuUlNirLqalU6JDNMiL
BZXHmOIUucx0p3Lw6CrHnRj0Q6P4p9fHc6beqEFsCfzXWWtHHnHwzY8S0DSj58RA
upxVfTIBXh79VpouYZmMKnzkvC448l2Zp3RQlu5ygETSFtildPEr7BqyLyW0++7D
9jToqwS8JudNquFh00H9cUSliKzzzF//jkwhGref18NJhpmCpE7++R5XdLVDYluA
kln0BtSztOE1y0L61n3M/2fYMy2rpJAdINWL5S0kmk68CE3+9bqTbn9C3rcH3fLl
kw3CS/Cku243IvQBc74lD1ZdJ61NjObDdxCEzLnEs0GRPBYLUJV7ghySXQyG/vNe
qa+4rDsojJT1fUMgMf5y9OEAhzyWPFqZEREg8hfAolGHLBXzpw4X8yUQQeEUUXaK
oUoIydJR44pF3CglIfvI0zU4c7TGLY441OmcJ0440MFT4MpPDk6s/y//NiDXZOpy
iW1+UQH3+oiQ8CTOTzYzfuABZHK+yHLamEnxt9hNQAUEJoyaxr+9uMgSqY8HgeL1
IuLUrRa3eq8euIfXx9RUHLkSnH7Iuy6d4J7/DoLcZghZRgrDzhoOIq10nT2ljqCO
6TIx81HlT5ftt1oSg58k3sMJMssIMD16OHvy1R2dVKmKu9hMG27uMQ4xTbkYEFOb
BFFARUmLCvlfMbAHJDkafKMZlJMoX4e+dx8VlrDkjKudmrkG6rQiSUqVxRlrGfNt
VGXMWru8wztFSlA063XQzuo0zCV9xXknx1Avz7xJs85kBPFmSsfQGoYazOe5Jj8K
TY8UD9azzIt8+B9ZRa9kP00F90A80cxEcRcn2COGbT58TV94YHykwjBWoBuoV/6Z
T5IvgE5k2LUKcugmaX6tJLKRmeAa/7r9/5fJ/wXXSoPZaudgKxsxuDxeirnr078r
rHGEmijHGyrInVLSYufjLvIcH7aZMhIUIrON3lt4do/zF/O9ac7u69KbudQv5U/L
XeiOAiN/6FzqzKuyIoNWhUC7FhZ3BH7Ycaa6Up6UvOz9pK0q5rAspsz/UE4h9gE+
MdsPQndJX78FvX6OoisvX0/BaHz7SzvKaRNuNxGTxPDFZNMG7Hv6MuBaX9GLG2RW
Tmf/RHTfcfQc0YMs9e1nQ/bZNFPUYaxHvchdKgXLYxwyJ63Ue8mBBs1tnWBb7bi4
9isNOZplYA8WjVIJtQHUlMFTNyWVSJ9gjLTUqscWwLwl5N1F6wLj+tQr8an9SFDm
vt//5EGZXI1RVHR1G0LLK8SaRCYGSK4zi56ndYFMMfr2KuSIX0tyfantYZSlxO+J
LxhelB99FNBpw35dpaN86Xpcr6PqS4Ym1yXEDiAQ692SMfWF+LKdq5est+a5qrEi
Dc3iTyUoz7DcQhNP9sqjIdJSVtSgqXennHSDLkWJl5uzh3G3ropZiEwUhG8GXmI4
s76dE4jXCv0EHPMSRCI3qKjTffyq09AWbrnOpmt8VySQ0e1C/Age0oWWWQ2xQvqC
Uqrl0YzIByCEXIpZeqR7qFoBB9R19OCc0M2plgZdvqjqFjZBHCXjDHLzJViRdvtm
+z/++msGm/YBSHzCtkveSaXvCaE6iFabvSnzlBE1++H5D/LYkSWTwdSkCpNsO9ub
i1aTLxqj1NXmxCMqqDsGj0+uaw8ebh0WTy8HOJEQgIOd198Ix7dUWPxYMfxv6+85
x1QD07MEdjOeef6v5Dvt+T0XKCglEnRMCanmZnSSS6f/yj0mxUyFuMQKtMj6zkHB
dFNKgLxtKIavYU5G2/t2JDYShxyz3brVerY9p/cAe9INWGDJkPwPVTeo419gHAdX
Llz1K7eQ5pE4+w/r0yPL0seFR800sf0cqQgEgLMKTzkx1Af4z2Bd2ipBrWEsF4FA
pS3N/+cx5gZ2g+Dr+Ow63bIhA23vhF6FOU1QCYXO8otCoULjBfetlmrd0RitPH9w
ZJTub/Mvl/rVSjdMNp5/F0zBxMTj2utllR6nJlwUt54Wx9MaYaQ0i/veMSzglVAt
ZqAOmVbO5nqGxFL/CheS26RuHalPYCLBCTD2b6/ou24crvody9zqPvbZQ16ZA7B8
LVY3PsNGZJrcE4tRGokP2XRcE50CL+XcO7LMMFSfOBLfYQbIEHhutMsn8hF6Wk/q
Bw9xqWrLyItLF/kididderbxt/E05+Pm0QBSOVl1kNP4OeifCQmwFyftUdnyc3/h
Es92gjcSTo+TOaiFZ02RTbE2aipGr0NN8OzOmANfxRZEW54IrifL3TqxU4txNwQ5
MqUIsYPIPn/woMeaFkrYRGfXyj8SzR6XGaz2z22OOGfhfHMbqfj9c7JmuNcUbW5R
SdhE3uU0NxPKAo/of18zhUIESUPK0/ycgdGwZRPPZXoIjjlQVL7xfWN8XB75Ojtn
AFdD+p60awbWkSZUMtCTk1PzTvSwxF1jj6Op3kakI1e16t9zu5lSpmS/FzCQYtUr
1tdFgSL41nzNBQepq47S4/11N8D34xzBRXMuNivvj6i/O15UcN35vWLh/Pl4/09M
lULXiNOnZz67NKGho7t1Z4Hj5BZgBUAR/BvEn46Yfj9xxfo4AbWGj2G97SDlmEvg
vVqVg9FpTOUlm0ct4QKgtoo+oCvIfxmLkL2Zj9Sd9VcflmPr1nl3Eherlw+ZrmLT
WQPUVdx+aV4ZNfk3FAMcTyJ4Vgx4N7tDC+WHQ5naiLf7s1Ifv04gX6ex89lkH1Vl
y0EM4ueVE79itqMMkidMNELiCTocm8QAr6FMndO9UObhhsiULdHK76j3hbsHwxFR
mA8wnzMVbIoRmv9JbJ+NsaUNjYd7h5glVz1W9S8Ma1LYpMAGq+44w2fpbQnUE/zt
dro88rEmnI1snJo9gEryMKcZ4GG9tG6NVAvglBGElEHNRLosbtyy3WeOlBAPX9TH
0oQr8lrk6vLbL94nEyFlSqFAIstDaIyohaGm8TKOUKwSypeAlB1IVDVkuvhBKfiy
yqtArelMLe70AwK9lliYdesH0hDY65BP2ie20xhhgozv0vDaq/1Agr9QYhJ1eI/z
9B65chfix1O6eYc77SHJY39PVWyMKLiA1h84ZVU5p1radK7QSALPEQsN+nt57zoI
LNn07oqxvo0NQcD85FBX2W5vUaTQk60SuCLE59Db75Yp+EZtw0ki7HeFohkpner1
FzMmCVrW3IR+8fbjvpVJw+7cBfAJfONd6HBub99oLLfSYHeSgHx1DZtEz2LCsI5I
zkKhjJ/tFJwI3xJrbUzYnivDLQUZEOOrG1BVkBALERlIwDTNXXchtoi4cOWgdfQW
73v+gJ2nkqTXLboHzcdlNG0hCK2I42+UQvBjW8X+yz30AtXhSKsSI8G8eql7C9Ra
1thLFYi4TYSt+2lIDhb4WWIZYVMRW6YaHK8aBUR/UqBqDAjE65AH+OO1VtO2R31R
e9zULFRkdF3gAOQfsvzmRMGwo0BKwn/fIX+z5D7UJleTpUsMJj01A65gnpjckvrI
wxaBJvmdfLAcGacM9j6uwNt7oz+F6SNGUHMS7xpjTqZ3ezzyxaV2tXIEXHqdgxjx
n0FGm0j2eO/lF/GOYAbOo5+nN6RRTJjhlTgSV03t4/gLE6IEsgoYYnw/6KYMqLTN
5m7SYEaNucLLBgxevGWU79yp/s594tfjPHcOE2BQtxMYMzWzB9f0+b4WBSEkk/tT
uV60Retytth2MDk5DKRIhkuawgAv1SgH24v5nxh7B2596Fs2a6PT372I9VDmFxI6
lzMAY6j5K1sYq2g2PGtYWKYiKZ2HAlzgJJZimcIcjo13fEr2uAUQz7yYQAk2piYe
RgOWzXjLKJFzIO/WQukp/ge4R+DCSgGbVZZmpJviBQYV2zJPRemCFcid8E1OFfhZ
Lzizg5Hj1ryRoM/VTylK7Ac5yI+6WPdXsVr2RSCIBl6/r/VuFuyyut+1urrCsVfv
w4gAtmaGM/Wy4NckxwyN4AKwLgTSykYj6120js6ZO6xmksHzlcbNmYzTA8OSpt1x
YYN5OdyvuvTVg7pPnue/TIfQcNaM/KfAfkN5s0/DR1eJjvzlIHuQ+duXRDv8ghFt
ziq7XQo7S8X39zbcHrEYzF3nFJiCntkMn+7596nHxnVvlSafu8fDs26eyj3jGXM4
/8lwMfBats/bdNGpoD04XprXJcMjwfG0DMvP2aBEx7OOq2NPVjYhec6S3fXLzwTw
r9bECjaEDpIsd6H19uOSJcTozKq5KzXy9HO5VH9BriOhyxuxrww6az/gg836hcF4
4m/a89rcgXbHWsPEcUcagBCamm6tqQ49ZMq7H6NIL3O1ClDXO1eoiKEB8+/wRJqW
4tRPBSXcq87RmBQm1oiIMLrYZOG+az7YqDSiwHY87q662+0AUFfVKB84t/g2wZ+k
6W/Od6+0+Qsv6eX5oqESG5jE60wxtxdBh43KPihXsBVO/MHxpsguPUZ+3moX2Q9T
r26Hrerg29Lwn6TLfWOaiadhfmAUvCYNrozh2yPC+eGyKIvp3L8c7aKn4tUR0L9o
xjzqafcCJTsswmQJxpIsUiC//hG1VJMxI0AsWwpPu+9AKTTSenpomu5e/agYd3d1
WT8T+NH05Scpah8mY4Shpmfnby/74Ypra530FK9oBtlCqGcF9l6rLdhuw6sNyEJE
Esug+w8AoQ7cLVEH0DL8DMn9vnMCrwCvN5a0oV1XByFCmuDtPlIpJH6o14kxe2Z0
bcKaUw/rFCo0eS2lV/bfuP7I+VxRyBW4t6/0WF16dtZV0WTCwqP+oaElDldzprJq
hDpkDM2jujBxVIqOONffNHXw1tjbH3pzJOp7VN5mhuAEvgxVkrOnXxbPCFUDqYjN
KhWrSgtASSrWqjLqzbWJyZSJ+WVFFGdtsvOlTtJawQKdH0b1pez9aZoyXBKI3YdM
EzDbUufdxXBoa+GonVuN/uM4tfLmvx6Y+vmYvy4YwAy9iX6kkkJ/S5Euo46wBAZU
nua99PIzGe80w5+SGq7WzS+ZOnUab57KKhI1jwKYLtQn9CZaZrE/ueB7MFUz0fLN
QEuannwChuN1MkPLxeU+OLdeJYi6Y+ECy5J8zhatedOZnx/A/mNsP3iaqqb9mNDX
nKB46wc0D5kSY1dYRdJ7WaE6uDG1aQ3F1BFNS03iv7fJxa2t+/Q6FMgvtrnuuV6C
sRtibR49HiWSwsyTNZo+aSTdGz6Kly/l0AY2Lys4pTPj9CGzkKSefAHURjnTLye8
n1tKT6ARaAkCwGjQqOQEUivqwGMqZao4mVd6v8hNZKiNiluNpkGxl5znO6NkiwaY
6PP74pv2hiR6gSZzObnPJ0QcmHA6r4oSF9zYSBLcJdDhFcqng0MFsVyzbkOlcUJF
UAR9mbRFYDcfcEorYDgLVfz0V+CGaOGlxavpokXgOSMBHBKSGfbnzNzl08iaYPib
xODyKg4Lf3nvs17zIrZJWnc2h8Fb2AX8azMOQyNDb7kgtqBFmaka3P+NsxVjKOSN
dZWbizPMOrDndbph0t5/QarK+KvjcXBb1Xf1U5HfKeIoknWW2V8hd1FAdy71Kp3O
PrL1yLNgl1sWjVxIctCA7wxRBamb72esigewfg+/kf3zMhAdSaC7pMfbKtdLS9OG
JlU9fKxo5tQ/UzoTvdc350UqfwhlqbTZZHNV9Nsvj7jmgnbb3qgyL73S/dQGvOFm
T/p0d9PkzdF1Q5uJAhjydSbVnt364pABJb8YDR5VZjME1A51vPvyHPrmkce5yjgO
P9nzR3oCSJWWuGc3uDuZW9e7xSgMkrHE0B9Fls9+HZm+SfbxBP8dzXSrIWNr5Fuk
a4Laa8KLvL+2xyd+tMVzVowmBmA3VY4QWIA6h2dveSbNsfGuQxe2WbJc3Xl6NUH9
dUqBBBh/IcUYSWUFDRL3/H4BksAIsnvLYb43eDLIV5HW+o/Ke8LVnxlU4Oyw9zR5
Oy19Gdk8vLrL9u1Xd7pwJReJK2X/4pmLchPlczyCy1XJov3IEIvd+oVx5Q1nv7n5
6PC1pO0GIPc/GXEfKEFCZF4kb5EpRmeiJ346+eCK0Ow9DRMrn6d1p4kOFekO9BTf
+t1jJ6Vr/1lSnXrssJxKa3YwmZ7a1dB3tlvmwEkj5bk8/GB/U+gFhMza/RyUYxUH
YI80HWCZn7n2oPO59fNFZCVlbw2s4ePy4GW00pR2/lOm4jWczAYW0kALnlET8+G1
1cyIP1zL7G4zn5mS/+p3+NVPqxMep4gzX1EBg6G3wW9PoJv0dwRcjbJYaobmaCHY
FcG3GLfhUV/dl0Sc202NtNnBub+bWDJ25vbEVKKz7LC0e4N3+yeSAYNxoHyiZ12C
2raNxdLTlf5BLlyJ9ojBvYiaHPfRgwrLh/xzYaXIgtLJKhyU0jY6wEOL4DWC0Yqt
pwpCllm/8qYB1SWsU32pqer++X+awvia7MgIkyZyjLQF6VYTMccqrIJwPuqlH73d
+TUFIX6DQd8gQrz7GyhuIaX4IObsshHnP6AvIa2Q1XONe6pUIPI2FHfnd6+zJRoV
Zreo1a6vC2fIM+70zXp/lGiU53/j+WF0Rky3x4AuRUF00sMVc2vfU2/2YcuXcKgg
+gc1/4tX3r0hQjOITJpBdvFh5JXeWSAO1B/sdlc73JiUrPvC/X1U1EB+WgYFtbis
K7w9bZXIZafj/XINjq6VtfxNlJGosDMLs57zLUj0sUZB3xgztteb4Sy/habSu1zA
UxYdq/YSEfitsy5nF1uajveQYw3sEk1hVKIbBwvYPALpwAqPVUHNxHNz1zRvtb4W
5owIKZapl1wgU8b9uexSMhGCcfj80cjEuiTaLiQCxl5KUdUbVe9sO3DhnFJotqon
eF1dY8/2Hpz4lSmenisZmOWbyOq2GavyiJhnyXXsSmemJAsN2rg5UHrg1aEyvRXN
ukm7BqxgzWaQham1bEH58u1sM3sh2QDOD5WY5LZnppFpxm9RcW1GGQrxu0vyUQgM
g5ozU06C14cxnaPU1SLb9aNT3Xdl6abHPa8NnVY5yY3AT2hK9vgrjs0K0LAHo6S9
t2unW9GpUuKhF9qhV1pqGYxLybTT4tr0CRmFXZEfXSltkOTbSKYU5RP1rzXbq4vB
ZivAzWSZNbMtqIoBS7CdLWgywqHbwGahFNNHjr0hU5TMquZNYOs5vJoK0rswfNFR
s5Qko5MYFAu8rIdnqqK25aeK7K3Ca/dyNI0ySyQRSvrvXQaLxzh19d+CYrPqGYPC
xXFEFs54zVc5VtKWougvC+6AlU69Ka5zaFFHhG1vWJWWTuoA7jsKspCrUfL3DJMD
Qw/swL86HKs0e1tAH0/knjE4Yt5MdZ9T3cmu6Ql57pfpeoaxUn6JulOqAdcW2VFO
a7a0mKHjCV0ZY4HyXO/C1WltbFsV345d9bW7YujyqAUKWLYOwiykON5MD+wGS7Ju
B66SR3oNMZ/anYFo3b4fnOuKObylA8324mmA4on+AESjt2Lp/5nkTqbbRfzlYvft
z0B8Fq+m7Tpb5jdfUUHxT/QaoPuBxO7p1WeogbD1KwjAcjy3cID6yZLArRuozFV+
AZurgZziR5vvEeEO53qYtF+mw2jlUY9txBgBVuur9chzsfOC0MSV6+EqpV9hOUwP
4qpAz9ITgqzScp6R8HCvoqtS62At8cE1R2IF8tVU2CCuc7IpWs9lIIas+CdLcDWb
RMXRIHGJMVksxlyW1aYRrsJHhWQKo4EAr1IqNP5LOI7zWUlsFWS4uZRuOAb29l0C
libt4gCWmra7/1+N/cuTpPBI77eRUnamclgkubMltoIX9ab/pHtncEmqJbjcmPRs
XamHMCHsVkfeQiV2jmLA3rFN9scseMMmTo7K3KB4kwTqqsvvP4IR7CkdQ2iuKBsn
ZVs0PmpiqjSp23YBFkIXRqDAhJfQZ9BYec2egk6NKd8NZR4r2IM8g4rCRWjX8WlJ
UhMvIs47cZ03B946qhf7mhYl+KWp4Z20cxDsCzwFaH5IdzhObkcYZY5ndoYf96u/
jwBRM3ekz5rmSahucKnehv9wKjYE6frmrZ8eJcTTh2PUoLseYGeUOl/pMCTReeRT
khSo9aFliprwXxIUS9P7aAsRf5X24PX0WZfGtzAQ9Ai3R5KYUcCL9r28n7ErQZzX
byAMlVtgt4gohh7g7Jp6NRGD0IsGi+Iw44qBQjfNVMzPTTQD+T3/lyJwBgLH3zBx
Y+kkqp86Fk9C+4OorNhn25aVpTo3fpG3urX5VsQi9OziTRunrIB0jgehlLq2IfzL
0d+7ZOo5ZDKvmE++iIjYU2SAITF8NT1hUwhC4JIgDVCeUyeBTnJZ7X89JzawmXl6
Qi6IQt0M2kbv0C4KPEvpVJDjwvgsj381z040+PhwuCelOoF53NRDk2PWAIG570Ri
baCAVk68WpkELLmSMV3n3tCAscYjy+6vgh9f+FyrsnKChUU1XC092PH+uejlb5J4
pBENcgaaO9xLsQRYKzbUYtf934cJuH053MgmLfudfPrzsjuWs/4Rk5RCh2IzLbWW
pMMq9yPF9ALjQ4BQiOizGIorD5iHwY9IOV8DkiIb9sCZ8+/UrwJHv5+l6J95yUzo
rIfVvu0U0gYKWdXTwdQFrOunscZCHK72A3KeuyfU40WEpLz2ZLPQFEJ2TphJg70U
G6q3bruGWRuhqTgEn16WMr+GveWmi8FArVDYRhXEzOo8697w5QyyQTvEEDCmM9TQ
rGGml9TkyZeunBN+KIbLBp2NA20Icg3QkwzrEf+uCI/TqtOMGuRMr3+ssp7xOdyi
Ntm5hK61eTRQ1KU/3CEJYGF4UnZ1m2COV3NPvfgJS6BRUihAkL8nQ4y2vCSMFk0I
AkK+xOx/ed1iT2jQguiKar0Axm5l5oHH9lNQ1VjP5c/WU62kvAUkgOCSEqVT6pBb
FKL72QEhdvt3bIZ6FD39ij9KTihsDGUalUCkyuxHGtVOXvqPCGwIL2z4rYYYkDo8
l0xEIY/hg7Hyl5G3MZw4hmlQ5mNnYeWyIj8CDhaHw7fsNQKsfaHrWv0sUWXWLGe7
GOlYh1XUrbbN/JHJb6RnuBn/4BNMygd2rIDka00VgOBrPLtQydYmqWwAAA13zV70
Y/hQT9fCRiIAzLtiib6HxQ7XQJ+vANqjvLZFlSU2/KDNtsDO2G95Vo0pgvDo+IeT
kzBRozcXaD9RanUQYfWteTREVjAQIt/zUImB9eb3EqWsSEdyXY6HLSEZ3zzyeiu2
p3kxSEu7skOau0SOl5ZWdyZHEnCE5P2a5Mfc+zdlPn+NXYXylbXx/v/OGdwqncgk
JsN5HQp7lyq1E79mgHcVVfCSd1tc5kkOLBKGeUaN1QRrRhCY1FUcJ3L2I7/x2wA9
QBZYcapGtzCD/k/aftnuSTmQNBud+vBk5xgk/MgU/H/Y6ChfrD3V7/YpAmQzu7FB
jGBSk9UCx8su6IUemwGBGfL5QVA/OYlezbSOEGWPQ5jvLdgrkTdbWNguswZwYsjO
g7/DIsVjgXNZgVFhzQZN+Zugf7u7l44W2ZibTfSouuWZOLqdhLInXpGd8mUXzzvI
KL5XXUvyvlqDIXR4TFLkszOEW9CZAIRAC3VxPpLek0650iBLUZ1mWdEPYSF6TwB7
6zOaVd3O2D446CZQ1K5/6Q==
`protect END_PROTECTED
