`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J9hlwipoPVWpSXXZz1KuEflAg3KMyQR1W9MZFI9kAWsgY3w9m4SelueZtlbY7CbI
fr79XNsYXiglGWQUFXth3QQmkyewJtl3QUdh2qAxwHq6urXULgk4HTGPVzR1T7Yb
WAqdgYanlCXSLpzaUl7YH5JgVToF03gDanGUhJ3a+08PNek6Lt4qsDJU/iapZsRI
4ny4nZg2Jz+x0Q1eXeo7ACRbkJ368YpCFmYwEy2IQ4HRkUbQblNuUPVslnonlJ76
yPRAVSJd2z5f2QnjlHincdT/0lfFnn//IEeTrQDjt512eP8nrCYm7i4gGco5TRkn
dSeOpNtIQ9wFjpnZ8Ldo5TaKQGLRWlC94HeCOn/fw0wSzqWb1vHOyV0BtfznwVfz
`protect END_PROTECTED
