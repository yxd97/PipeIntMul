`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XsmvF6Qf70yZmZJ265w1mPfz7PCbwKZZs9hHnervnpAh11IHlnMHt/IQxj9wfwHH
P5I/Q2BrDtfc7oTQTFFjSqEgM7+mM/O0KtQkrz9mvGCgPs3dLVNhDAA3+/evFf0N
b6jPzXDIwlvw25n2F0KQYYk+WJB7w1Nn8x9WT5zp01GxqQWuFUHBGFUTdEcChMX1
XAYGas3y9cLqFC8blDQwqbYm3DBWUXbyhaIo4MJ4u6X18d/hzcRkngU3OisDCIHz
8In9LPhsjU1vun5Ry0whTDC2rcqSYs8TEztvnXJbpm+S/NLQYGbDUjmfM50XFuxw
QBJfJfYoF+JFg7nTAhQJ3g3NLha0vuiKqlMhtcLtUemJj19mtjHOaXCIGAR8n4pS
2HEyZPSO9QjExmpql2+parl5G4j+73ES40h1UQkPFHQ4DoxYTbVnSqlP2uJb3X7w
a+Ax4/4YVFuNncvNoNaiMrhS+C9aSzNXdnz3pmw5A1YwS2MgBREIiYpQIB+Xk/C8
aPwCdAnkmuBbqJFRhKzj6Zo+ZVKZfv2Jfziqt/iGzH8V7Bd85z5hnH4OBtUFd1Sl
7Uhc8soszuyI8Xe0QxV1WTRYIpZ7ruRQLBi7wknp4oyaW65D8uH+02EycaXMzZWK
/lCLS4yTjM4aoBRYuX2y6TPlNZK3MvCTsEwWuRA3u4d5JnFWeV1ZXmdehzYTratv
SbXmqgRbXodEYIcWkmbRp/Czml17L+Uz561JUlFCKUPIDjnAITtEBcB8IPDJsJ9P
zBvBnDUa0EOEksY5GN+4e9i3p+qRgyX8ASVgz9wzEUdPHdMxOlndYxZkH4w4V7Cc
nuZIxjahDDQ6bWq38XhIZ74K6DH38JVYQz/IyRXvuWMuBKuj2nv2zG46fppfMO1E
R4ZWUclcHgQTvdfBZU+o/A==
`protect END_PROTECTED
