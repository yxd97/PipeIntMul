`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MYb2dSRTmcxeM1m8O1QVK+WcEu+MmlBiPxELDKmpbtaeOUO3bMkjxCgcdKgTP/OD
gl+rrgCnBpbG8ja1VHCAieNhPd93DLFUey6M8IEKyjV2Cx0Y28Ry8LKF7TpAZILs
2JWU0WNjOJA3IvMqdUGcy0riNUbzZOWu9IqDNFczWcx4NwucKPqeLWnlVGLSV8DT
Vh89nkjHjgYcuf+cDM+n7ZtKTfp0qTDYZpEGN9AzNVBhFBBKwuq7xwfD85aTyZPg
EoakVg98pNinTgscVpvIf3kyQD2p4Y5HEWUmrkltYBA7oznwsJrE1KbZ6DWeM3CW
ZJTwhO2ZwX5Xbir+vZS1WX3IJ6PfD4aC9XR29VLdGu5il/5I+3HsKNor3WTZqgKD
I2oQ8ELUrZFf74dKWBaP+g3irUXBLOGS/VZSDWRghaOVBXsL5Pp/9fZfMIL9RQTy
3DMmvbqplkMvjcK8L4xD8L4T5LcYTtGwN/d+U5jAAJ+i4GtPPDtxDPDBU8inEeqk
srt0al7aGAcv2OuTZV+T8T11jK1WE0f8Yf2UKrlvDoIk/nMsRpQYd8E86h+TwIG/
fQ8ulvRyPafrP9OGfPlHc/iwJfa8a5t8kDnKNNonS5sn5yC5xl/lOanVY0UjB0Al
qxkp4178dIS6yvyI31v6wGGGH7yHJoer38sVFsUG83PF+TDUvDW1wN9uZESXr0SI
X80FzhHHduqEZWjo2XaR7p1nSKfuyKCmnVIxMPipV8c2wCSwx+5FekswyfenvaHI
5Kiz1v2Zh3+tUP43y1TEn9/yycnaqvpXcbN3y621wAkt/eMiVK2VK0+SwnWqaotG
JCKSwFMA9g0vkxoY7OC83TmScC9yXa+xJXmqP9Uc88Dy6RTNA29KwsKqDQg5/fqs
cNV/IaHiCLQ1w3sZHqCKxQmNxJzw7fMTuOhE0+nh8WIv4gwQ+bGDSXhilF9xd5H5
iYuhUNBSSzmiT/j9YrhxsHblqVdXpQIqthIJCiuIbEogggaHQg/82abvHx8EiCPV
moCWSyawQxgRAtGe1/eA0TT1tqW2CH79YDhnZgaUsA9csCpo9LBW/UMpJqD1zTCn
w9qqxy2cge0U5idOZ0MNMLiXjD2tOml0x6D4lrmEAZrCxeAAn0Oqsa+x9Ll7Hi4U
AlhMP/LSxvO7sxw0avRhis/KoICheTfby7IuKhTdg0GX2VBapXLe11Yrc+CD/9KH
mfsGzh69DdWtgyCdiiSeGkRRT/Xsd8LMN33rQqxzqHcaZpNCKKfOC5TvKokah3Gb
zyEzIiG3m1d2eRuRUAxZKJBgclfAlmE91wPnPy5Dt2Bfjq7BPJ1THgVGVeW/28Gt
ms8ZdqYix8ul3pRLp1CU9YI4gcxAVwgaM1VOKKsS8UVdqj2dpzjCWOdV5aOhyx7Y
/OnOhiQnt3OcI/bdwW9oVS/hDCb7vx4uNAu/L5DUT44df0Mu0ZH3JMcYcFrCV3ff
gIXBWUCgxW9l7Jdf4fL6gWbOtSzypEeCzSEoekCsuBeyWSlgu+ENPEm37ber2feW
aH0S15+S0NoUyyvExtLOrTlJeGmSVcQr8/qV3S9FNB3aK6LCdajVuA2qFljnoodk
LVzTzU6AtauLj5nMbzNWRgNU00tg0ytcR+svaqlJCUPYks5PcRLJTgpMAyjcIdsE
eyJCpu31AxPmPASfg8ryvFNRjM9j4Ia/dGy1GZnjiHeBExAlMfaroX3pG+pcTZrs
kN54KhxaXn1FE1oF0TC80wbyyuJNgYL5Pk6Nera8FavgwZLpM5XgL6r5xlPoLOV+
6sQPqt0pHWVpxeYl/U3ccXa1+IYDDKZA/5IjvFAXI7/uYmiTCnJF3uVeIlbteuFM
S2TxeJN4VZARbd5KT4s/ydOUJu/l9DdRsShTD4hJy2qat5uTRv88Qp2w0uc0dS43
McJlKbpuH6ZsXY/NCbCR41NWIHLAQaM5Vc9ByOJh1t3wMlqO2cuQIn6cOkWArTQx
XnB1eqUuIQqTjQcPgP4lwIecL8UTb93MorjMBA8aWbDaNAo5CpdzkEvDNjfOtHwZ
ea0aSdBM2eHaAqlsHWBWR5IV+a2M7pd3bEY04toZh+w2RS2xAXGjY6/7pFW3w36F
p5wEe8Yjxb8FloIksCtzk+gPHfQWC0dwRkTB+PcnHPtKnnhY0m2hAVrPWnUv0Bzg
gL8UIUjag+eCoo3YSQb/DztUP9iqJCNRRX6pV+l55Y8iheNsz8boFGsNNMchhHxh
j+Q3y3FPvt7bPlMsCD+mRLqa1k8Y6vaFfcC0S1tiO4GWw5p1xmvtpZ/qtunFufVp
obox7ViatNpBfL5704NlvW2i6EXp2HS/E2ceSmSNhpmDGpryV4t++PZS7Lf4TuPk
vXOUFCUg51h4QIrVWCTfYG8pCcPidwwWy9JAaLjSlQVgyNug+F9GXVSzAK82TMNi
hFTAdz9CRnHFURAaaFakFg==
`protect END_PROTECTED
