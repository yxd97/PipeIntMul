`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OiskxxJwU5R3akMq5rXkzq67V7tueCHDLhfac0+LKNn/ElGhBBo0jOF0JeRa1qzE
pRyU8pOXbtrC2QAtlOW+B6CFwTs/09YN3ZUBVbfxZW0Y3rqZo+Q/BacjcaEdEz27
nnRPWMTMP7UGAop3ehCfu1dmIPLUBORdrIs3Zmv7H2ATOrlnDwqp+eqR9ulK8DMX
nggd2q39jyV5vexFvlvVjwqweMWhEvi9ESvqJ1uz1c1xuQRn32/DLlzS+a1axSz6
fDQo0SU9K2eg8JpPtXohhOcpbmMo+x+xdKD8UsPiKF/HAn7U8xn/on2juyb4Ae76
ZTFSSnmgbLXsQjjdPty2niN95dbyuMJCg0iPegb6E4NaHaSLhFcDGGXKjESZ7KqJ
oSdk8l9m3Ys8WYN0odO/y3K1Naf1PvrpOY2TU/xOcebkcphJNwTV2ebrm7ssotXu
Q4seDbMQG3hWWOMjoa8ODrn6kcilIzuM3LYNReVJJna5fGrsfKp7C5i42NmKERl7
TSUsD1YF/iV7y51wzybl6Xi0fddgPklXA/gwTjVdwI0yFE82glqZtLnM+KB55iud
FnrP3tud9czHyE+b7kgg97T3o/8aLOu38gLNu/05vOXujHDpqKjl4QuCPhr9+fJR
KYyaDm8RPPmfArlTlRX+Jj26jjvhr8s48s2BEeobzYxrjP2C9TMDULiYose2OOlk
DjIb41jxdABQVVS8skgn3LlUTNnxwYvfzOEkm69tzJbK0alpEE4rKoguVAJd6d+W
tF1E2+G1mQx8T7cm50E4p6j7NhhOcelIsRcDMhhAYedWf0fRTajIEFWZF+TKWiBy
KPv8sh4UX+2o5VgafaRgiXzPFRbGF1raUGD7X7yb3+g1TBrqyVrLK5lJdOMHk+PY
2L+MiC1ClbDYG1+wA++GbIYrSa9f7mZ5UGAfIWBLClg3PqfVrzr7+Mmc6UNf6/wM
scPCfWZeQi0kO8EjTcG1tQ632vPwY+gM0IQntv8kamMXtW9BX0rzc8KKKehihdBR
PuhyGEJTkGJy9FhtUMrcsFgu8YNUbDCGY86WFZlailRfIRrd//tHGBmpFU1arMHs
MW2h4dX0YaisfJeS78QLfYTIq5XR0a4dAhf99Nt17KJ4DLKaFAukBpsKnKuHN+a1
DYzfm2clFMUh7Vx3tLMs3uBfE9MYs69++p6rD7ALBbwSRTyZzfy9bqTgM6IG84rd
hx/c4MWZajXI8ZWuIb4fhmLOo8qguCrqsUz2mJtvabEznzYgooViDSXQnlPqLsdy
ikWgIcW6fnVKeD1z+dfKif5cqKvO76FlzvEb75w00C8K62AJ9oc5nT05cdYg6GxB
qrpoZuy21P+p1s43tmQ8O1QzUN9TZSGNDxs45fgOFjZtEvmQAzzC2rrMzX9XyngF
mM/C+zZTPAJGMd/6C72SWQBujrgoKlV7GKodKv+A13RDxXTjfQy1qRYL5IYJz3QY
ucmHlEBjSxrwsMuCRl6p/6SlQS2DCUBmyENurEjWZOZ86X/yCmjWhxOuLiE2biZE
AjXHho4K+89m2qDf25+R5TYPDEpysrEO/SaUhiRq9WwbDGXQNrDsKane2Klimtu3
mz39nRAdOrpwoRorUlV1+dbSSbItcqejdBTEtmik5fKb2Ov6D33ug2C4h9b9Dpl9
PyiDdus7vrtDnhG1JnHVU5urMfNxUJQDWVvOGIPR4IuTPASxxeX964Br8LwI1QVp
GLjaNPuXd4Zh9BRpVQ9fRbiHA6u/fuRYAZGhGZCEb5Y+y0/eFQN126SiSbpgsirM
tU/sL5ZCOESU4XtYAC8bgVcbBR+U0fw55OIpRKBUESmAiZ2rswKBkwlIZE2jUMDa
kAVSYgoQIZSzAr2sDnfGAG7QReMIKkk2yva8yWVwB+Xz8wvZ2yUJZnx9/EL6lAtb
6+PNkZCgvkyMdVSpbMhn9NL/U/gL6nZ13MBiwJbbYuBBtJTNI/hm1Z7qnFeaDqEq
/oXIonwPBEwg4KzXJYX8BQ7RL44G5YGQTenXBlkvdYrzEMMn4Zg13jwmSw2gjQtr
PelyKn9z/t6HhXuuOu5l4t6gRgcUJpCgUtf+W1zMNRtmZdUhTUcldj4OEcrQbQrk
MjDZwlV/YkX7tez5UVAepvCL1YR7RsXJB20PT2SO+0Id84oBVamBhiS8MO0y7SrQ
CA1uQLVTPOyw9hIyLhZWCLHBDk0yDonLFwNmZuHiZ1cQ6zWVehmh+KTIy9GpsWmI
p8MMM4UYbzvf0vpbQEOtJZFzBb6qYLH3e4VcX/TR1G1o5PmvKAXHh8gbqvpb9fuv
5v5N5tgWZ6TEyfJnaQUH+Cl+8JHGHXVnueHKfYpZ7Fqcal2dS653vTR9hReBgOhL
XRjLa4Z2oZIpGmOLuV8x93yhtuI9S5FekxTTAWHRvdJmmBv/ZlZudGYbIUZvVVon
h5J7aAq/lZq7BQdDmVW2YzQMqK5+wGyd9cc3lH79C1qkpoYskMA1xifkDFy8annh
kD6z3r7F2VtLUpNw7ohUjkD1PdqEawZs+JV6Ke7ycNG9tQEJ403qqSG3f07BVXIh
kcislPetsUPt2rIGvoDEWazg5NbAQqJxbzsH57DdzdRYBIxHeWpGAagK8/ZRpEvi
KFmT3aUf28qk2fWi3x4/3gmM2inDQkAmAZ+akeZyEGQQ4Mh8/0i2N7a/S8PTjtkF
rkQeZSlpsbFTVPHZjaYot5BcmQQPHpsRAreH3r7jCD2FlngTh51AF6GFw0CqdZeJ
w3tCZvtrkuD8+zVGJKt5J8AyVfFib4/l7nxpid0ZHOmezqYvwgPFjo0Wzvvmg6MP
RIzJNF3mrksTHz4qUmfqjfd6X5AXYUkijLbEbPUJTKc=
`protect END_PROTECTED
