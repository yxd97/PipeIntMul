`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ddZ46vPQHUmYwpZdhZfndHwbq4zaJurwmlHfmZ/YKyQSvrlrfdbFJr4n2Tnbs1vU
G0ybaJgW9q4XVz6+4JU4JfjQg7EWkF4nGF6DnOTGav/YeI13zV6IVTNmencz09wu
hhktY+qWjqLD5qRu2BqSWpSu5baCTpgLmoxWGDtSbcjnz+/38etcg5K+R53ZnGaS
gg+dAquKdQSW5pZ8Co8HS8wC237kE9iQ6+h50Hfyvd05nDw6Gt5DTQxNukdI0qdX
hFeq2WeqDhGw2ntNwGO+jvQJsVNvthO2+0wWQog8JiGaG8EslZJ4P6EVj3owMKSw
nmp7E3fc9Y0ipyGoqzllTA==
`protect END_PROTECTED
