`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CJT2G/U6NyhGZNB9pD2wxf0h03asj1kYKD9QfHS/dnVWB0VQ3NWRXtgmrv+mup4n
MvxOvkMvnVFkWhT85o1TRZaCwafW+XKFT69YpoUeFPXYA6i+d31xKnNnYOPubRwa
xicxZnsYeeOGdYJxt6vNrhbJ6VPNxQ4O5buf+rP7v0EDfeQNi2JPZSCLHb1Qtbqt
POkJixL83QlDGyjVLi4k/NAtFqYULNbJHTboh5qUZFhYw4VvhoIuDZNhsuTdreTR
FXyTwfOTGwPROqQadw3PBHaKa99cHxzXbj3e29gWl5a6T+amz+8ZUmlQw4cfcbfI
fN453Gi7SJhNDuGnXe5RjvgoqKHhMarhibUCNe5W1myxD05J1MSDQiXAcPrAbtFA
`protect END_PROTECTED
