`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ef5sabGFAZ75sdXmG/NiPTaO508G8rQpwhXlbvrX8YJxOT7I3cJB62raKji/Z+3i
e5MKQHPIsPCdgVYSYJQPeu1bWPyerxWmpB7G1oPVabEAgPGTcRYDTBKLOKysaGzM
WmiExGJEQntwl14ynLLOqGmoV6SFpFXW9KmtZxarcETtRQcUjN1E9oPo4X1MDhH3
4UlYd6ofYRcIBHAJPaAR1hXhnnlOV+XhQnb4H/eGIzV2eK+zkoM1sHiHmq9p3X7l
Tx34cqVU+tqCjx1+Q2w2L/LqdGx8jatmNUqgHF4sof8ymv/XsWmvdQydoXDSRWKI
ep48vgon2KCcRHtE164FXTsJK0m0LeClxuqFd30OITnyLgpCvwfx9Oqp5WJUR+VC
+Ov1CloGfQEjabuyVNLZFZq0eatgozF5R8MrJoVUD4oHZ93HOL9Ad0mRwByhKUEd
R7jaCOkiNGk3IVLqJtpsC2YPWRQqZ0sUjwZV6RUq29TCDhoWd/+n6XzDUItS3Dmm
LFmXJ3A+8mBVlgusLDZ9gOAMmwDkAl63m5TlUFgx3kspH99oNQpsqz+8FAWjQD7/
NgPT4fJ3xeGNWxh2foYc7kFVmiIw6AiDfnk6LUTHO4208jt27B4bXHlq8Y2iPGUR
i8etynWa7D7bY++z8rfX3g==
`protect END_PROTECTED
