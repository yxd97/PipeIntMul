`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s8P8EgMQTgpq6JXFmYUNb0eWkGUQEutOX3h8OtDsQz7tkeKjOM0kFsjbo5yDmAc9
+AyteNN7qXjoEZXqN2dt7F5HChPhCy1tmT49luH66tfj1aoyobTlcBn1196k8Ipu
zbwwqoUd71sOG/rqw5NnfXcCEnj3zHvOX0sYrO2cpewrrJJW/OZY1D76sC6PPr+v
tHYTPbTIfUtVLqmag+nOgGzVVyVNGsWrWdNLADW0jF4l1/SWl/vWrST2BFebdMcC
bx4kSV+NTVwd4eIbaPDWClXOrtIKd/GbmM6ioI2U/vDJ58ArGvfXzsZekEO9dPcC
oEkUjFYWoCFleFaoI7yE9dqpDQiPeUgubEwz10H4b09faHjhpOjYaQO8V6FDFHmU
kyu1nE17pQ41+EZEjVzM2HhcQWOmo5kkdd63wVdvl+xypXD1d73CFic//YKqLU7x
9IXOiyGGOA6W6puA3iy5h2cEtmf+OlAfP13qoiwTIcLtRqmJxTaJN2HkTfcIhZgH
20oOf930reO9VfiD+aawEoX8naeIoJVEeB07PR1SRk+4ZC2jL03iyALwMLm/yGz6
eH+gK/uWvmaRaYa3jL/brx48EX9fEvEbVK6I3GLPz5BdfLciz4wUlegx0w/M0Pil
MUC9defF1dK4ZnNlxqSE7VzXTdPau5g5UigTCnJ3DsszEzk0ZIaw+ykradnQglQi
kKFP49fxArn7CAZEBFbTNKgU9lxFPxJ3qCRM9J8UfQxMVNAGv43UeS4Nb3eLtODf
r4N8usYOYJfNiUk+6o2EMg==
`protect END_PROTECTED
