`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2F42mSAhoPcsL2hXdA3Mo3Wi3M+aCQsHCAqMIMlx8M3U8pjD9NHqqFc786uz+xXk
QhRdRN/xs48Xty1t41SHt/ardOc65J8cKLfXN8qJFra+Ej5dBoS1aX8ylMyyEB8+
aCxBAH5ZiLl+JCpZVxO6CEvTc11VMvQwQEx2Cd4wXozFRJAsNj62PwU5JkvEGeMr
f1QNq1yvIXFtKB/VRG71kekfzUzArZ4xcoIMq9ZC9jwoTK9GH2/3WW55Y0uRai8G
Iv5SfFLRWv4y2TVLUiGXGQpNe8WLzIV7tmP3BwJTJiw0V4bKghHKZoyek5B5x0n8
IGcmsijbLF5/OiEl9A+88OQ4GB84GMRTTlDKU6oVjg39gdbQjkfvmXr/VW7sS8X5
npF+AZRjJtQ3+tEs1iU6mQ3ckzACsCeUBq7Gl7+mNF7yzJGyvO0vw9U98LMYtvXz
rj120cZ4Rny6WJDFT5U4qFBjgXAXOn0aN4l6UmBwPemm7BF2T6/pH/RR9L94ZdIb
ti5rzXeFTykH82GGXUxGWZro9ONKPJs54uXg+VS2QSGFOfd6Ub9H6MkGZTjwddaO
efAV0k2/SytS3ekLKFe2RlDUCwIdm0d4UyYywtxjOySN8ZGjnapSWgw6TV76KTjl
EUTtB8RqBdzEOJGyD6fO53Un/lq1eimWSRTy92xRWklEKZ69z/Tmz3O7PeOuSqiw
3aC7iryZ5XJex4KdDpMq/UfFZMSKk3EEOY1Fd3SQE4+HTZDb9lytKj6Q5+EnyXRO
bSJvnesb/e6EcFtT1mkTuM9PkqRwlNnuNAAblYeQLLY2xWjhg1zp8LYNzQKsk1fK
WJHl0DlRoO/G0836KFJzmj7fYEQGW113fERKBxPjGe7BxZAxx9ZpFDWwB5IGT0jA
PwmVfdGJQ50dZvGXDWt5JfvaHtWqWr8hej36PvGO2tySZ/HAprKiqJu1/lDSEwKM
UF6QfX+bTXugJBHkHGfaaisrAozQogZVat86AHEkuMqotAL6S3TtcEwY3Z4dS4iA
y1BqPIK2P7aW34sDLx8wwnBvxZntQeIzkmXksPtheuw9+Dp9buqaSV88TWo5PfFa
Le1eKd/7ZgzibX4+GisZ9Ulip6pWkiIPj8l1R/niZMla8cdezk9asKDHC6vsLeAD
i9GDQZcQMkIUPvB/nJtG9n+IoVDovDKoNlhl4g8JWY/NLqcbjKxKltLcwke/T+eL
DQ15XUd30xrHTytXJ8zE4Lz9i4JsFrjMOeo8HJajX+aBOr3UOqbiatfpmHgfqRmg
Mba1jl8itIvq3BIuIVR1Rr0C4WWwab0D6/xewZQGi+da9iYfrazbA0NOEa0Gvjcc
DAgiuh0T0ZO68CeMFzmtDSmQLNsLbB68M4G1Ac/Kxh+Vbj6GuO7KjV4ItNUCBUMl
FP4pK3KLKXWT5+ITLn2zFr7SwSJ83vJ0pNLKtxRUuYHEvLoaMRJDcndOHnJqMzNf
TyeTPAkh1/bzy1bxE35xOx5A8joDWQSOZ8vXr4gGPezvfNQglLntz6aGSmir3VFR
K2Txc736WfzjvQ9RI1mbZyVsNOPp8mn3/M8sMsBS9ktYI98wjJs4Tw4fnQFnwklL
w75Cv399KZ5DrSnWKaxY1qlapnOi+uEsPlJR2XbhGcYmuQXjWpQqwFfg0zfFTBUP
69KvRFKIbNe6pErlGlDqSSHWEsQmJFTobmHeE6Ueo76zFQeIIQnEfjrgDlj+1tdr
rnbnSjjWijCcTEOjxZSsOoUmOkF6ZdCjaKdVHJ4pY/1lXsmRLrwysY4r5z5QnZIb
umaZx/oUZ9UFwJsCOKbLH/F88Q2jU7dfqWxTvyNZoqZZDN0lj0a9iuL0ZJVVQKcd
6MZph+ZLHhfpf9ie80HdLjbLtpflCTHQGgPNCv1LvTv97dHG0ZUPRKfhfHOako+s
9fmTCX+IjdJA1Wgo4Q5kfZ7eelNJtKWWAsrdmcL2Vk+mwc4aNvxBR8lWpKWaIFsx
Q4ok94Jj7YQELuM5B0r0DbA/rsM1tn1ROSF19EKQ56Wz/BwQGEChRMO6IXAqSLzs
jaD3UGOAmQFadFmX5Uh7XTtwIE9x9p8fAPaR85/ucKo=
`protect END_PROTECTED
