`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2rxvKtFeO4edtOn/puN2cNT/2xwrULRQqFxeJyZjM0Qj/3bZobDj4mvz8xPonA/C
/il1E3ZYkfTs2wOs2QilU4U69E6ATI3nGhT5/7XuGqASEvFzbeqJGUMRxBLuya8c
qaXsHDNlGC6wf7a7C/Cd9P0iliDQxN+baNgOL2kahfE2HwZK2Vfj2dkFvAhs+yTU
5IT8MtFMv7MskL1p/y2DAenM80Lame+rXczvnVYA+ok8tkRA+oh1xQHi9IFOIVNO
ucQwjv/PWiNN3X8SHl/Yhn2+PUsGEgPfcBp3ZaObkOnAgTddHZHxcArZhjhi1J7i
GnJnmb3F9NwsfltBPlH50a93mZVS53mwisu5Mdb5YkyY9YAR2ZhKhj9MssgOGeew
TmnsLoAgPrgR/yPzqrDv0HrgGMeTGaGh9i5JrXwzPtyu3tSAlJ/ffcx02/2Xsi82
IPXwWnvwpm6XtRK/max1vfFiW0DdmwO6K9e+UExgHAcurw5Evz8CpF+q22wlIcZ1
2bCFlqqVx1ZZ5OiZ21qekBeTlAJrPmlwPrL90L/j6IaaHyZ4rHRuI/yJPv4I88Lw
XMzysJziOeoxf0Moa/4OlVF9oM2Bo+zQa3gp67aFhFUjC7GHTOAA0nDikcyhr20m
FvhcAekNl0fsh4QiUqNtG6GKzMK2BKN+7D6CyGJQuGpDlY8cN3gH8VjMOxvEf4Cm
wX28JhIajeBVDz05xiZsHJ1Jb8dWyYEKAGDKcuWpN25Nn4hqX/4JlfYcpZTDCIaD
xzZzjH+YVmbeDEVI0MaCqN8R/x4aiIqwdhUPsWlhVDGwtTPOGphIYLoy1E8ebG9h
kLlyVY3UyPFUlj24pu148p2dDb7GIBJ8qB7FBJn1BGtkmiQ/TU/LYILq3CFJlsR9
+Vn3XlRWdIAG82L4F0U/+W0qyKnK6FC61F2m9Ojpc0G3PDllFbOgq5dXd3SHAFr4
TZYjEzEYNSW0sM3XcpLv5xh7Cir346FDuucauzLxmkzHYapry27HSIaFo4tU8YWf
GIYLLvBrbDeQoh/NYcCTptOx4Cu28bww7BKuPlExiVsgynxcy7vWYPfMjz4JeeAC
//jybGzsp5rgHs4hifGKhizBEgtenH9tA3X2VPh//DU/lS0exp+bSRw+4tqXKrH9
X89lxUH8wUD/OKHibWV6LTX6R1ofZ5/1knXsH42dk+F3N0TFPuCk7mIOtGLNVg0N
QksxT8U0sV8FPopcFcry3QcydHRfozQnI7lhfQwdNN51HWbqYZDXBoCfmYBNkDQc
LsL7YMbQgoN6HMgFyFo1grfwoLk9gtnubvDj3h9XRHtTX1yBI5nxX3y7T7FQR6N5
FlU59AwdBVAcePg/d0zqzTWoCyK0eQF1Hyc+QrVxI+NhQA4qXbk76yB9denwLR2Q
whNVxo0JxqcdOEfBhlH+o8WfGBY4Hao9qqTTbwViRtt4tunfhQCy/ETbJ9GuLbTr
S5L+kWnGSWhZsjtXqg9fN1eWhtiALlwTQmG48TkyQr2YclOn8DxSNBO3gGgbe69g
H8Mr4shPPcRXGB/8WdLvWUWjV1z+fiE6uL9psIULkp+HoxcpcUZtIyfcwPcHUcxy
P7vFtPw7gBdQgqDcPCoKfiEWL0muiK6bN03M8r6SRi5uDsAWuqTMKnF57V5EWWUY
6Clacw3JP0LEvoH19g2hzDBdeVO8DnRHwNYpO7gZ6wVljs2aHu+pfYQKKiiQAnN0
Xga7kfgW1FoBkRz6VyAJOFOs0/8t+iHeXJtlHc3PRMHHVdsRtzUAyvY7Fh/hY9LU
HorwtcArDpTxNS/rCFxW9WbCdW+VBAOixxhv8gvCGC/VSG5bAAAow7nYH4uZdQx9
iwhUYUEtb/vIWC5Y8qNsKfytfEH/KAVJ0h47dE+Prf6zNz4P02hSp6pzM2lYm2JQ
6naw4iSJQ4LmY9lof0/Spg3nb4ujRqU9Rl39qANPQd2fzzUjVBDwya6E0OKPyezT
y0B/MTceNQRcyhD75+qvci7V+yjfH11IuVUXePE637RjyDDFvICP4s0zMby+TE6L
rsVkISB2noXJ5DEsmHUOvlfANAGYaeIMTk2RPj/I6WuzuEDcbHIlXqf+xXZWW646
QJpsrJ8ghieZlSwid7ph1/iE+BPDWKq8oAB7SC6tLlA1BENm5l3anhJgWv1YQ96k
FvsLvesz8xy+4TDQ+UWoiRJU7HKi7X7SBDrcmJNZ6Xc3YoybQ7uUZoZ/oBkprnac
W8gPxnQT0eDeNxT0KgpYdJBCcSgjMriH1Mc9JllqvAospsUkHSjPttOOTVA69HeN
iq+QNMRx/yRvl/jbm4sD39p+wdBmSUe4j13B5R3elPZqIWIRIRVHHcw/wabjakA1
xRXhXfUZ25zWXkrIY0z5RiyhxEcqgt4OF3/AlR2ZUo+fHNokLwDy1Ct4atIaU47s
iuOllHpc0PdR4GQ/O5tdJsrtmTld/TfwBl9uEwV3q1v59qobTPXENDdq6O+sW209
upBXolLXM+1iP7LWa12InYrQPA6cI+yUypNwoBJKkbgfxneZSP03DignhK6RdL2D
qjhsr4wAGpfrIVy9oLJUAVutndLHDMd493Hdro8gg2CLt8rukF+lwqmlVJe/Js9u
mQyOYVFucTkc7OVV8UVrzmsN/ZayUZ1+BCRcXYP8gFjljuUSXd1SvZjsRj5VlBmm
qnmJlA8b9pTHD2YdFi/MpPSh+nMvUMfz7tXXNeB2bx3f1mi5Hm9WA24XCnJ+Kn7s
iHbRvawJxjbCWi34AO4q7CobAD2O/tomx3jPo68XOxznSDFOC4q+4Jtz4HcTeSYq
6B8jpAvF/AXdzi9rLN/ZRSySuB3Y1w2ld01CtMed0uJkNEXDuE3c+QBgqX7NNCq8
bp6BxOUnsrHxPYGF3DwLM1reusCnudwe3cwPdYeY6APLDMcmOrJPCu2LngNULGeb
xKzVTi6cUFMZoJ6UksZybwe/zSI665KK+nW6v/GnWc+nvXTyumXqYL5LKjXtAk9D
5Ve01iKbZ1Zp64RgxSei03bencoLDx4TvNQjesFWHosf5L2S+bq87R/jl3gFE1yP
d8M8Yq20sAxx0bvz86m5XluYjPHWGfRZJNv6qGAU9A9KfoLJgJFpmXb/YKYGZagQ
3qAMFhpcf9UEPAkWXZuQvBMI3uBBhmm8lPWhy9HVyHHmNRFKF8ul1Rsrdnd1bRT/
wwr9lGhVHiniXLevRW1K6pGwVRuSHpqbvuY3oq3lR0ZODVKahsBCvizUmd/4h0LR
dUuuEeWMYIGQGZlQasWBeeHrl+HXRdR4+3sGkiqG8p4hQm+o8/v8+vteh/3/+4BQ
d7LSXu24W+QsqP9PRs/n/ED9fa+LtraTXdAjW4PyI9lYeBZQWxdOk9QAAbbugdeS
shxxTlkeLeOiI06L4k6B2i4mTpa0sDlxQNAmR0rOjX8CDLhc0fG/BwxlugEXmVwu
rBnA3yTUwTvVRYZ73PsEy/VORBLy3Kyv4vgWgRYTAZFbej6jQ47aJUCxsANbimxN
nyGEo6feMzM4coXrUvBS3WUMjRXNZYK6tDeVJgrxvUVftDjcx8jMvjHc65M/ygdM
mNkh6WIEqRAPgkBBjqD8GnfbGhEi972BsMNgj+vCewQSnZuE4uWNZYUC8JZWSdft
A2srcpnSzamIAjjY5Px40PWS1fiU5/6BVKkqzj2B1v7dRvgFEqfFf/IQmWssYpsU
QwgI+tKgAL96OCEN54zUkBFBSAZzZ6KIsY2D4TxKp0yQN3fdD21HOSmrEA4EnuVy
VtEDd21Ia3jmHSviDNmWrdqncaCTNrqbklsgGFdCVv3F59VxOC3ILySSybKBni8s
Ys2E2w8LurmyQOjfjobwikYpyZIJ7Lf+6WxZ+KvfqDlY1vh+hM/RXgqjo+Ua1DEV
gkyU1dE1E4qE5rRMJzmsiFbD8noaynKOPvf2ylPWZGydEoouAaZ6iusgb9m14Gkn
j2EvwTbcLQ5t28q/a2npRNYrliEAoV2YF3CU9hWaISBVDD96AwcdbpU852kazKJI
xPpG/lZbwAJatnlZWU9ChgJO3qsA1VmMcBWlzRw+ucSFWWfwBZcHpbIkJiIACV/0
gNMhfmNuVYLizASCGzpSNbT2po0RkVCOn3+wLBh0pP5pDFCtN7Tc8rpqs/GYST59
1VxZkZMh5oEpuZ32il9xrHxJH034OaCVxbtA/Yin6jfMfCdnc5Ra3CWYZKminCdf
ac/+iuJnyy8vUrwtynLfSfszYkoM9AaqFsCHarSjwljbn02jmMTS6XR+Xz3RGHBo
+beNHlo+9tR11MYmrFP5uq+vqjQ5IWD4cuFqkaNm9PkunqdfHRQUX61frZeZ3ORs
ND7WF4qTeO3IP1HPRaPLt3NjR67SIbK+95Dc0ytKhSYQvcU3Bw+QVnItPo2Rs4qA
eTmo7Ln1/UkofH6OEk2Qyb7131uXUn30X2e6edeQ0RukQ9/fMD/FY7DTRas/X1Mr
rQMB2Z/XZL12m1AWIwpvfsTsUoY8wKKN/XPSNsfiJpEIE78o3AiOFOjrJ1pqoVMo
jIa3B2ZHkytVCksSL9i0xMFOwZE6PvuPxd+wuaCKEoiMNUh9QyNGG9O9kC/ox8p4
syG0b36MyInTFdEyLrWXD7vNlOYjdc2rfedX/S6tEK9vJPWHHi04XS+JrkW1uacp
pSubm+GjWaKkY/UN2D9YilfRA3auqd1fXq61lUWyHDoLmwsyYhVHcVYZ//vvejjO
Pgu2Yux1OFaYz9C1S3vDxUaLa9PDN7I+EwKdSV7yY10MnnXfWIdTLLozBsOZt7Fs
ZT6anLdlanTzIH/YwD/dq8wRIHcynRQ+68nCE+I9NPKtNtJZ6NXUUH5zlvEmfdj9
m9ZalKRxbQF0ZW347S/o5K/gv3DpQc0Ag95mFDlgu2Yo3bpdd/Czxj5t8cxqBGWG
KfHHnz4SeZOoIycdlQKDy62Ocvsn3mgtNuXSLFGAr5NALkG4kgGqq6XTVU+rdeYz
O88XDV8i5nRblKR1J+aImL68qTOQCSY/2mQgIGwuNptkblF8N64bXClgQkdely6a
bFugfd0U12FMab1Fg/QRP+yqtJ24ScZST8JsQ7a0AnL33aqxbXdoMkl/2ZEUfkUN
aL1TtO+XAbJ01oyFf9CH2AlFEr81n0WbTt73y3vzlzSpHmACmJeL1zoz0N9mjaqm
lIfIlNzALm3qlUjBBbbnYjyPm5Q5lVpuniXWlWD4ni08leyAyDTnRRftUCY6ObrD
4lYv75nKN3IWxUonq0YHSYjHuGBjDKO3Uqck1TOFddEKyWZSYFyOjJZ++2nAlo64
z5XBx2Hmp0y0dOIMvQnXbG2tf5yDb0fQnLG9/WnEa1/1ltvMLptm6EmBOw1TDy1l
M1m3Fvhp0RWf1bl6QkjZtXJlip7HKoFQuEbZD8gRnQXTNVCSQkztAXAxK8il3Cxm
XYoVf4vTBYu6MrwVLPccmBydJeBu0UTGDXXXQzv6wLBeGUBL+rt0RPATN23p1nxF
Lcnp7MNFvvQzUeldEy2T5CVnz8cApJ7F1KLZwI55IQ5E6ZO3ntVkXCYM3DDVlAjB
+V8ft55DdiRhH6hpsikMot9v/PVefz8dJuR5tjPQFCzBMk94qhNK2OqH9G65Ifqw
r0Prl8r2lK+8wJvmMMH5ygBoB7arc39bm7acB9Nc3MBeGCssqTE+q9pE70/cEIt6
O7/ULbgZVb8czZ2GpPWacvYuZJeDnQVoBXmqLVHWeea4KMm7i1+7VoLwmlgIg5Vy
AKkjLXTJQXb0VPilNbij9UU/h7Kc2HoLkFseDg5BapGpT5NYVvMjNm8d5tz44lcO
7TfrFAQ1/l54Wd3/jmtJtOB+5NuRomNGP+zIwAXgiEQEIArKVP98A6ds0setlgRb
CMjdHBkfoaax5tHxihTN6y3dtnzsffTQMvwpNxIxtSVlWPopMUdrSRELwWhZ5O5n
UD5FnIdMpgWEhFYP2Hy7pCZTkodCuRQ9mk4z45yU/fc5Xwnn+HP+tbTwZwz41lFO
nGc9te4ZXPWzoI1jbDuiJE+ewLGzsADwwVZHT4hTE7jcicFTdKDDiCUL4qNC2wku
hfmpFUWjvMZNeqZVGk8csevJvmqQOUgZgqFLAO1s59G8wJKbu6hlixzqSXbRnASt
fkVMHtrLvhoXH7fiqhtlPD43D8iVkDLiMjmcSPG3W+gx5uQelXdyd1zhVlhr51OL
EDR3oI9eKVsNbYgOR6mpF68Wxi2omNya1jzrtpTf7oTyw6vZ4wu7ifNlSyVaXxkJ
bMJI+PHSg+H8cw4aCLqv0pq76ZXkcvOxGiyZm0cexOxZ+Uc33QU+/kchFGbJy+7d
+TINnjU2w10+HnxrId1AlVG+GZEFE0O6PI6H0BhLIUZQHxyX+NS9pxJoVlWzSMvk
SDWraNmvW7Vv29RRcI+yVWKNZsBqJ5ld31NUAailj7RsxtbMZwejddRnNDSnjmlr
C/XVKbqTSiX6i4IZh8DFgRgUwmldfBVIFsrJQcvqteTNQzjCW/JkRrcH2XKKp3wk
CGbCwAuD/pP2pdM/xz18chLIdyGICwToIpcdTmBNISmHCWCgBCKJ2AwF159e03Xx
NqB53cFt/y+NStY+CCuwBQOcqmET5nkz5DUvBB0zWRrPbju35eILRh2y5BJ6eY1G
7hcSVBDeiNEGhQ98Yi1iEwdd+DVPcyTWaBbMInzvOuMujq39WWvGHjEHFRgiuzeJ
mf9eAbnNseRvsBAo5VfDgHxLikGz1kk8vpMrVyBbyCZ2VIoPZnTW/0LWC/2v0N/8
OoI4KBC3WYMU8+I3iuLWzquj0TGM68GoDhSwMPDWclwAP8Rzrtcsp3eRlQLXvqem
4b0wm3UbRkHU4Y8zalirMLGOZm9PJ2vPbNXj9yg1wo58+kyZxostSasvetEUnyaM
JCEEdSbzhxr23hkXkh1Mfm5TvPSKutpWS0yUuJQAJ2RVGi/kFHTacCj747lpByii
t6fq+lxT05zHPn3QY4c5mNp7CpfKMfjMwpN2Dhm5zcpglPLM2Qe5pWm4NvT8TJ9+
WD5BvOUL8M+v5dGOvTGwRJ2i2gathyu/GGKq5CEzaAJFNQwJDecLWvJ9z2tx5JD/
s2CfAh9XCtPom1pWLgYmRCP4OslD+5V1G7zVQUQgp8Mu7+IXkJBFi15ydMRC4Hmv
7OGHBJcHZ+VvM2dQtepxmapmP0zkMiz+OHCVp6cVfsa9/PGMJp2nxHLdtEIg+lyI
U7aNYiGYdZaKm+4Vj1g+xTAbVuLYd7i2Yeeu4h9YYI76jAY9hN7k71zS0PodYFY8
StWvU1s+V040yTVqiahDHhZOWqmSkJtDPLRWC6+5v3TWssk6I+GgPfYkV6cnP74q
Hvn4mBr3U6ORprTISWBpcj0RVLEtmCewPpNdY6Iv+HqphCSap+W5b4CK3G4qK+84
LAvDyehawAlVBbG5CnRGu4DsQ4ni/swNNWFJVlR8RTEecO3cYUzdroJ5tRfoXnsW
NttUGlnTFsBdClTNMABUwr3DVK0/b4WNfyxpy6abWgi/mPoQQZ4tTJSXimxZolcq
1ySkXXgO/Af2vwRFfNtomRhdCn0srB2lJbFvagceKzYQ3NrliihTQkWpyGHrkIAV
1kWA44Km3o9UgxHz6gcqBdYUrHcOd8GyZZPen0cIJZuLDlHx1wLqXYkzjG3JRb9Y
wcU21iQHIhKXxgatjWvLpFWXqgoT4p2YnM9oRBBeKOjqnb2G3sa4C6wd7GYO5Bw4
HkQZwEIREZj2bimxqZHSjzEWdLVnxUndqfGU8vUEEYA0wlzxjucUKa6OYTl3COxA
0m4utLx77ILwlC8qVs0zCTYA8x9QRujCDCppaI02q/eVD3IRaK+fncx4NF8Tbfqx
xtyb8muBof5kOBrqpQovb2qu3lWMUCXFLi38+EkN9ghKpJxNlpfTuVNYTG/gji9k
6p6S7RYUI4XdXZyujUWqhZIaIVdFG/Wlkl6eLTw3BTjOA//VMlWS26c2dRtiIaSw
U6pWC6+XZmT5aQKfsIWp6rh/1rzJFwW5gPs+eZ9ZswJyKhwiZunb5Fssfeezvsw4
tJiQ5XWn/9sP4iDixMA+TtVkDtRtayc8AvXAiMH0TwjQa6pVwQ2EV5pAa5bI2z5q
q1h/oq/aboXzgzwxYheSXaH6UrpTvW4gcXLPApjQOCSJ9DzxKIMmxsTUFxtc5Fa9
CT/3mXQtD85csa+Q6iYeXBpLzL1Iqoa9NGvUbma4w/RpL4484wXf2YBc8wTLjcbS
FN2aH1n0k78XHAIsjQO8pemwwujRID2PMO88M+Q601NBJJHHRjaxsW5PedcA9Hrj
7wM6gjfv94QxnBqAxt60nTfnYGyqx7Hv+oRmklSORpakpu0x5R72+uQrLn5Hu2LD
Qk76qrucHJFkZwkCHOAXk7tl6RY/4uz2xq+BfGilyTKweTqIE1YsRM2ZrZS9Jhve
CNpvg5HyHJSTwVPs66J5GP1xomO+c2mnG/0iviuMqorPHbgTEu5NUw9r1wFEIgDf
VjO0JOwjdmqUeJkcGPh4ZEVsQv4IK1C2iWD/1WUohT7fAPPuO2LRXPf+aOfBgEZf
2m65fPNAxde1gGLe6hUWq63XbfVb6MNy3FsM7HOl75d9ZG8xmx/2+DwUs1dmA/Q9
uGczl90mXyBdc52IQtTNgtIghNcCnuKfjBGJgUq6lT0I6FFW/8hmqG/1dpIn0tC/
9KsUSfX4T0dO9nH9UZ5Yq/6Z26W+nwI5yjyc6aVhUlbCFUs9C40U/RnPKUprcwbH
P2hF2yxCvhfCT4Lh6MpwgVQ6C7LIhEoYzzFKLLs87kQWEX03C0eVsZ0FZgGWYJBB
+vilBjg5kjuS6gWe5/5j+Jkgpd2ToDURpDI84NxivMD62zPUHTT35AXN8q8gAfjp
V+dg5yfPfzVBx9rT5IXRkA==
`protect END_PROTECTED
