`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vx+DRYKB/THUHWibiKoLRaJYp5EvnZL6k4dQRSPBl0AJG6mwNWYoiJJQCT4q/pDb
E3URuDjzRQX+ARvLFu52aJ1VVVI/tzfQCk+cvx2OvveOeUuGdxFJNlQjuZQopKtD
bjMVTqku65ow+WW3fUpEpyum9j2XPaq9GhBmTfiLFuMNDE+w67VcUu0+8J7iJAel
S6zTuakJF9hkAB273JD3wDSwRd//ITCHp+IAudLQ7ETGPhPgWXTwE/c6zoC8Mkne
d9BDD4IXDEh7B3Lu3tSy8nIP2DKGsX8jvLpd9gkBm+etPCXGdfPNfSSmhcik9OWV
jCTXJieSrK6Yjpa0RnkZ/8O7ILjsMPSLgOxB3agwzwwSe4nr2u1UWglCVC6WArkL
Dli4ePPWRIn/O7BM6vJ9QoB9oWMiA3y0o2+4vObEubXJWnGAdEpS0b5TrkXV2KI0
Ry0kyzuCyFMzUQb3OGd3yRdEMywDM0a2LsseqTAnqGb5+c2XyrLhxGyFYu1l+faS
OJhbgRJ98R7yduc+Di/vlCXNLrXtKPry2kMlByzmjgIqjCfwfu/4YnxjCT6K38J2
gndR52iCIi/efyU19KFcSS2iUTs9vWe7R57L8a/8waT1wV/s1UBQYO+HR6OsXbae
VGT/Ag+5IFPYkEqz9gtATipR6On6STbJxaLW1PsY5rVjvLiAMFWyU7dfxUN3Dh3q
tUy5M0Qn3V2D+YFy3GGjl5f6/kglvY8m+OHQ+5ETCUm5bGcDQF+88jL4q5BdbX1W
xdCdtpWAU7l0FKiG3nw28Q==
`protect END_PROTECTED
