`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s/7sSUMpJQ/V/0S9sUMEcatEujwZ8sZ1vB1n2Fs3p6kDghmH745cNHL7lfzAg7MQ
l4z4/jkvGELIwZDwO/bvE7khhAT91WC6DHS5Nc0gDVUAko6oWnA0DLzvNYyN/D8l
/3gZJllG3uC/NibpIUspiw5ymIYeDJK/om0I0RE0KKxyeel74C7J1UJ1IixCPbYD
w35Tky9mFHM4okZBkrZJ/eOXrCDvvlmG0Fl0mZt6Cm0eQv+S3A5EAExV5c6M5GHj
B5s/UlW4QhLv9y4Cb7bJrrlPyQLRWKq6XTJeEvVGuZ60PeGKPzcbbiS6aYkvyZyV
sa80gFrNEvmGsQSbnappv8ziZqWr0KLqsbEZRxZUTHPW3NakshnR+ru7me+5vt/d
I11Ml8ha/E52LTfQ4NQ/glA6MhfafVNSXdfPDCaWPOsoDfhrj8RlZXTLA1mFcmIY
4pAV/7FGyj47offbb+j3cQ==
`protect END_PROTECTED
