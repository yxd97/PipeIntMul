`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qRSZgALvKSEGhpc+RerZqAK4ZMINTQPnCQLSklB/rh7sGEp3lsdVPGY22sfdBcpk
Y62biYqRjPBW10lGSlOoY876uXmDvWoHjquKc6JqpkkOZVqCo/s6yBseoaUQLsHz
uAeh5l9jzQO1e0UR5t9rUFN1jPuz843kg//kQg8YqhqCT9Vk6RDetjadHIUMAddi
UI2WHvtShybzYEgVaT++hJVooxwzqUoe3u0k5t944zNMJS8vbQvZVbGhzCTDjh9x
dLKYVm4MiuL8JmgubRSMz1i0WHxmhDSqO/L9jUaMCErIyVyDFgk4378O0Ruy7hYH
KtpmpiX4Qwsa3/lTy84Ny/r5YeArhOmeBDvPgYyLTG4Dg3/gjHCfI0Q6otw4da4T
4CabVBncV6dvRkXcsijHPFML7+7rsiInjXa+XQhWHQTnm0Cfi/3a+hKIi7I/Q1pW
OkB4TkRl/8SQfHKmc5kXVhTzNqMit2/GbC+m070uYSCAKBhFG92X9qGWoxED4SVS
+tFkeMUhe/wWItRwPNHdzPekuWunIEo3EraMA5eqq8LAiWSOlw+wDMySOxEfRSNy
lp7z38tnZoUpJ7GIQx8zszWmaKsz3V/t34oV0x3McgHslmuU/p29EgLMMiFApqXd
++H4OczW8eGfsZ59YDTDsH81VrhwJ+PO3r3ygyU/zQrTHqqoTDpQBiUjBMiABxop
t94l16pDN685pAecqrScKB00V+KuMH7RL+T2es5e8OdeUmvTKIyEoHLiXYsz8TnV
V/0D0527038p8hcCmT/Skz7o3DfaTrWP4GG9AruAaOytpbhqygOxkuaEuUYJ8rlm
qgrNp/FwRgpn0+8kOP6Ef8QfVbixry5F5+6WHJWqgx788gONJ+S/NqmnMGhJrgrI
69xPRdSi6XvdEZ6OYMAuOK9qaP1SM9Qr52PVrGBDGHvtgXa4LVDjrR3laHKmhNLC
YiI3/ocYKuIfXeT5+oNBe7CbgftONvLKBhUW0DztpKI3FlX5GiyG/1q/KS3RacEA
L/fQIDkGH9w7Kazf+Ozv3YkpjSMijTJ5pSCNfGPaqNcCDg0fEmpKdhJIzt3sCjvo
l6TnIMtOvGv2SodPdsuPFHzERmTR/CGhtHn9QBtybDbJGwMzNEbXnhchGph80uzW
mCp76u2ar19mmeABtcdCrQ0ZXCDdT9t7g0E7ZSx7BypvbWo9UQ9B+MVTByj9AOxT
sHGPNMjCv4kLx7jTdgM8aZEXetbDAsglZAbgr/uZdhG8n6jkjQfZsq3fgyivskwk
PAN6QKuI7Qo8/UcZrhrdNoAhdr3tHeGwTd46eFna3F+2I/3aq/dXPhbC8bXuzgYk
fOU464kWahRwZNaOX1ZWBYKRhOSsMCoXXf7/9JTArfXRqg5Y+HkvG3Cy/Dr2DCj8
/YxDcA/kvQ+GlOm/ZEC1Lh1RjUUYjYu7c1FcqlqCz9b5tUWw+mak30CYSFMO1IrG
YhLjJBj9xX1WIzEt6XNuy0F+AE+PsGICqEs7AhKiVsex6kZgTQa5Fm1M42KlicmY
+1MXrM9/vZgMT9dzczUriyeDHGlwvSziaojFA7ZKWG1NRZkaxOJzDkTydS6gxnqq
+lPaBtXopPVTcuH0pl2Uxv/t7euJ1xxCWttjmVb4BoTdbz+reeM5kI01NSGwynoV
k+n+mwkmcUMTDjzwGTPbv6rM7+uQCmX8CjLk2zj4TRLk6tw0j8liEIiO0Am/uTch
idWyxyF2xYGNT1M/wqdDbCIVwGwPIPUSkc1iyieQgFlY2U6SB4/0Y3bWHN3j6DJB
LULW9s6h8NFvODdv6bnlvBc2d7pDKD0X9nkiurW4s4Rc7YZgB/zXvkORv7YNX2+J
Oa4HuGbVCq6YZdNnxNrfP/vENNlu+j45usN/LqRq/5DWqNoA6xYhaW6lSEfGrWdP
OzT9iG8GAe6+2tEByO+WxbcIm0kMbKb1Y2sHrpLHnrasRO2zA9Aw2gAVqpUoqHqI
jQBYhMv6RAvcziF7+C2pn4iu+6HihTWB7hLFd7MBllWKXt28NE1wKZv1R7jmWc63
KMnwAUievkRwoHayEhvsM5UzrNY4kKNuH1I7sbYpeLrwyT7lRlIDTZ1m60ok48B0
E07VTB4hlL6HvYOpLlNkEZQcLS6ABX4V7QP2tCTfuJ7V58VjfKiSuLYQ/PWmZKHe
LB0LMNRNQkgN5nrIjNgSH4WhVlIpNOnDhj2bPNLQzOeCYr2QlllxSEBLRiwpUdbu
soKittZctNAXzVhI2vh4Wp106v+7wvrThjlj6AzNqoYLmJC9fQBa2yDeK4IbnsYH
5S2lqHI5EvD81+F+TIp4bjZZfXBMywDcPB8Ik34/IfHXt++rBCxOJUQT2aXQPPG/
ZuPWounX18QqpkAETkQHMgqr1V8PsIVkKJ4Up/bhH9Qxll7tlCHgrfFRjC/cuU14
YbpztAYOoDALQHgLwqb2U5qJ/iNHpklotVAzC9i1xHNoZYtcSv4xzd6nqhhQBGpQ
o2PD2wMn1y3w+E9hg/ex7vtexwRYL31z0uPTJByhKS3+AVwUhouV1oX5mA5Ad48w
ICd9g9oglIhIvEh0ea2c4cADSfT4TOyYQ9RpdRcMOclj6oDrY3ZZx+UDqVI80Zao
xX7xrPf5D2dZ86qrL3eLGQ2XVyBvgVX+7UKL7hXIdTw4aYs5hPVyuA1cnhGaBOm4
W+WAp0lLGMm74L5P7MelzO980O3sD8NN5BsPQ3Qlwkju+7R/ny1bTyk8SIz/rMOZ
oEm+REY0Z0OqdFPYy6F0/TGEZpKhf3quwsPcuu3WORE4u/heNbeTSBUxVq7V0Dsu
8PBrEa0MIDmTLfbecS4suVHadsSWJUaYIr7YvQQRZ9AtxDAUL6LGnGzqbdYviVMp
YT9f2uqXu6XJjxKXnWeHfJCCesJyFsXYF9ID3gnXJGjxYf7KKl5oPt+xZv9N85eQ
I8EbJW3KiRfZ5P7wxh0vp/4NtI1Q3F8/OcclRXjlEuKYaw5KxzvMOe5TVsKDMWXd
JsEKkLmopCd3/ZRmbLK8gG9E3dy7iSzXpBAtWXeyQ9YBncDC/0xp4lySttf8rlsV
5/rZFlfjeZiiWqgj8BU91uRXpPfCk+w6t+t4ZZrNGI4JJzSP95GdjmNzKvgAHGPB
oWp+BVVlZLugV3X7qV345+SImx2bwMmLzLHzz+TOlu+r6WEPDmGizptggXOmm82h
8ZL1JGrOqXtHtymBXKjkw/GWN/F9E2+YhgyAbOF+uQuuYPVbXoHXR9GAjs+lVhL4
YXK1WpG7LP08AN0uCda/k7m5vLOH2BwM5NsaaFed4Whl1Cxna3MAGGmEXGUv5cID
4TUxLmxARVfPtDIJX7K8UwvkkfjwaX4FGkWImJQQvc3pOXk1+RFDcvj2pO0FANq2
HjHHJYBw7pgQAeuGbo6ULReRwG+Pf2r3MX0OEZ1AbiKNntLYKyVLBNq64gsYnriM
mpBZ7Q4Ondgh1DKvn5hPQV0trHgOOM5YKG2mOs080Kni4a95WtZ642lERk3JmdUR
MEgZim8McuwCTctMpIG9q98CJnnR8TfdShO7LbCR9hcFTeSswMbSsvDuMXuRe4a+
G3lBy513hmPK0Ub/G/FYH+p1NtTZNF/GXEdMj0h2FawpUtEWPFMnjvN0JcnNBsOR
VbZOq3sV+jIrZ9T5bmuBMVaYr7QPvxlL3H8TwRKy3WbkPXhinxEzcvYBhmEhbT6N
bRIDSb7PS6FHpZwxfDjj/34SU3aZWScWhILzo0ANC2ZgAfWWuMTXx1Uuy1xKEeLf
YiqYMTTEWX4HBH0Tnu8oCIgwK9b5e8v5aA94JbV+bcbSLXumNoykMnAX1gzCC2fY
7+yg+EmKZK+ZtFLOGRGG2VpHnEh9XeO1A2JowlmVL2YGVCI8g+khY8TSYDmgZi53
6lkEdQEGoXvooKNaPKGh1tmuIp3zXEWZci7wneGTQF0TxMNzzhYdRfzdBRSqhsVm
rpfSgq+LKKEru8ItGZQvAqGocxT41pNf1dYCYtbrlx6fgur8suvOZqQjPyLkFHZ9
mNC+k5r8laAabQnlrshSU0tiPxs+vjky3dxmHuYXL4jUKCsXql52bEcNn73pPvJi
JFTe/CGUxTY0QV5UI6xNXGgtZalJEq/QPv/ugg+wBuLkPe32npgeFBVk9prQXkpa
f6bSwTFfK22mk8sqFErVbaEUskceTNOxlxvX980JkaZ9Y/ZdqHim2B9+tO/a1jnO
okfCX86W1MHuLoZLqR8ue7o1fZvlSNpzSGsZRQ2V07pwy+iPq6Kj17cv/Hf1Adl9
WT9dw04KJScbZ/LMYzHNnTWURR3vNBuJib1nJxCMI5WD+r4xV55TS/GFaJ4YVmkv
ghoIIdKfnv13pR6MEiBqYm/oAOEL24JRsootqtAXMWqCmBGOlnmT/s3zisMrVVBg
Uuhzbzk0Ws8KyTtKxTkTius4yWe/Xsoz7Z6f5c95RMu+z2b9Dlj6+MRzofr8SpAD
oR9s9/QVJFA79g1KkPDcpmI0WF3bW1f2rh2kLAwPgqTLNYW8Mi8ZONnRt2CdM4P8
H5vMGH0mN+5ywX5so7narF+RoZNIMNyUN91whsryJLJTNlpxjBu5YzrcKAUVrVSq
/e9f2Og0siB0UHslwBaoX0ZCNgd9mTjVQBmaKmU+FVA6xFHtvRINn0JJOD4PtLvL
xH0wuoppKBgwH3VJeYiLuJwPRowc2yVVZUzt4/MtFAMSvBnKCvXCAQPgpPlRRAh8
f0vyx1Pt9eWUtyw41TNqPfBDmmRxtrdjr5dcZFo9egBVK0LX2J+t10+bl+Rt5fwB
ZY2SPpm7CWA4szPozvKV+Z/pSClTye8ARg8HXSQ6Td+kBXbK7ckamk/L9gY1gU87
EplHjhcA5ixN5hnoOJ131RJ14bapZsrN8CHNCrCbjnWn1voaX9X1oGmvNcuCALE/
BtJ7Cm8sTKaaSaNXHMGG+WfLrcnGDObPWLyWJvjsYIjB9B4YZe1bHrxtVZvtf4mC
k2XEiN90QyyA93fFbX6wxBKSRSQGXjyTDNl2qJTP/Fej4zpKTAzSrakLp0hlvmrm
M0fU39oIHmX0kM20UyhaY0qdxIqlbPmjhQvyyPDLqNfEiYHZrWLAMwXmO7X0tBYq
Qg1pNOCUhy+8u1VDyNJ0vRpNJXi+5Y6OOsdzNn5HbC0vtV3OPBb4V1Ua4oLNDyHc
pwlLyr1b4LG2B5nUokxVnJntlQCIengY1FjmvkwD4YGln0Jxq239WNwRcxCjp60P
8AM5wMVkZIr38+ypRHoRVHWtOQjPXoMXTwABC6/la/bGetvMPQIiKp4JvS/0G4jr
qLFGvI6mzcGLG5eeRU0SZbGhKfCBPP62PnCCwGuKJ2QZcYy62+s2X2xRoKFZiyC7
+QdYwQjy1mtknjX6gbUWkO8zNw/jmjckZVqhMHtCYtSyVsyqXP72iG9mN3ZuFGnE
b9WDIMWN7QEJQ2L/8glkGdpC66xaHBlVyo/wY8CefgjC0R2xzQK4T9d1P67yBaXR
z9XpJsSvaFAdJjOoMKrC1TiO9BXjQN6BnMstug4FltwTE+SVablLUaIk3m2p2SNw
GKcCZEeFiNAE2yjmb3gWpacLskNatteEMVeGXTPOtPFvgoXTC3KHNJ8c4xUvhJMm
M4t26mbIHGhuYkBQdDeD19WAfspFbq35m5swUVfgIOIsTsI/Fnc1wgADqAU2yZBL
F61AR1XC4MwiW0aGKGY4YTLTwaGlE/BSxLMf30G7jCJbWN2CxWeGAF970KCzQnKu
jJ9G3ryMiDhpJ8AocTwaqj7v2t8XrFd1jxKewutWjJ3H1drMgQQOQRNUsy3qXjt9
Ip5V6ZGq6+8T2B516wDh/Lr2scZYikrfWTtM5x3KuTV131vpKI9K904yAW7E0t2c
ctw6R/duOhPIc4ZV8O3JMDohg7WO8WDqCXm18GZlLx2NNb1ny64ejeR4kLeT8Rhk
x8KP7XHpr0SgUJK2FQpsw8knrQMi8fdZSt4rq5MQ+rkrVaI8zA9HHxYu0gOBS/RN
pmRFXL4PPcETe2Qk77sBkQPPsTfAw7I5tWGRW1OxAmN+np12mY1VyEiJUq7xf31K
jCG8K+Cd55sVqtb0wQTbC+sn7w17a1ebX4pa9QDrswn/04LpxyQ9OSOotd4LsD8G
qaE5DNY8M35tWEbSrf4frTLXr/o5YtPTjnlKFv8TuypUEYzaoY/MQSrosSIw/DDi
2Zz7N521L4ITg1kylShcXSNvIr/vS+7MXxUYooY4rGEvqolnooVDEuA6Fb976LS2
3qmA5WYHrS2SfIjM4NyDLO1xMMjqaUFJk70RL82c9rDlbEt22b6eyQKfKb/0dnhx
PismoROYkMqdA/29OScfwNgkz/8AbbAcEpXesyjbQMMze+WNdNnRNgKB2t0d7XFb
EodfXnnunV9/uCfYc5lSdGKjDDeB8vtBzmbwS+SoLeCQsGu6SpTbMGgQUYlskGuk
61uRoZQs6PAaSLkgM/Chh8+h75F82m5KJrXOMpaeb7FHyeVLaD7Y/MQ4OT/pRbac
Uvkf29tofJrdQDgxFfk9a5dPhgxKftVD/pqi8x+pYYH2DXgqulcl5QHZxml2lLyu
MshneGM/YMjaZgJ9Ia1y3i40IpG/Quzljr5tRRHlABdn0sASLfPmSPCvwdtKSY/N
keR9m1PyaC/nwpSrsYcfPYx1nBU05V8doVbqrTviS+fvMvEoffFQST18k5nS2H+8
zEyRWpelAoqI40+t6windzhKQuzqELqIRv6Rkx4JYitutetZwqsrsZ9alTC56CM3
UPy6tjAxl4Bj2yrAgPS2QnZoeSNPyo6gbZ6/btAgWOFk71RrWonFCZj4Gi7ZhG19
TXA2dDX5f99vFE3oBrsMmID+cmN0PXLRzBb5xx7O7pY/y05md3Qp4toiFV7JJTMZ
8HjP9tA3OmSlUtiYXeNqFLEtMfTys20ZpwqPBZPI//V+YOOoa/S3ShYFdR/hD9cB
acqZ7Mv+J5Dz0ksRjlTxeSkrr/Yn3wNTIKW1E9Nhq4LzCztMiu5WAwekH29MGrP6
9hlgDAEzNpKCrr0k3uewyI2jRNQI/6y71yCSaRMAvWE9IoS0ix9JBYEzXwb59B1E
FI5Q3G56r/LCtaQwGnefTElrrmiriaF67QJA2VRT8dm1zzB5BnK59apZ1u076Lpe
i6sgz+HbrnhG4XXpceYFcDZKxjkabIww85eFyIbJm1H0cbkEHcmWjhJgYFhlxOhC
InDKqAEDTo+M0MTC3YmaU/RAhTejuMkkIw6Nt/1m+7nFXz5oOi9okQaoy11LgoLd
LqwqKNdjcwcZ9XnKjupAFbzaGGcwJsEKo1HOfMxM04XQKg/YQotWNHFC14dMOzxc
1FAaAZzYLZaQN2VVIyCiojd9QeO/0MnFm+TrXZPjrOYMi9I9xWIQCyA05Sba5tdR
PZ4Tg5Wqur1mqMfxV9BirRz9I2kfw/L9w6HBzuYR8TXFMZR03ovPRyj6Pv0obAVk
t26pw/DLq4vPR1Wjofna2etyD+lQPSRlBlbTY37hZbBDsKjZGrR/7Zb8Zh89NEu1
qmwwt4K4pUsN/mdzk56XVsO2C+sGnpO4sO6LEfXyv0QztZ9KHOma2bkG90Qun7Eb
Z+aQ5N0UdDdrmvf79FwjPdj2um2P5KJRQPz3aFrX9TWIZSqNBDqu58eWn1r8a6Fm
5Ccm++9jIPD+M2O/1ZoHVNzN4XQOQ1zxBEfluUkxMME8pa7FHVGWYOE8jsYKuC+6
ygxJWdBuwU7P2c9pXYgg4jaeOZ52IgkH6SrCFLyCtL+txxSLb7M3SaT0zgDpUFO+
bjWOdeWAGeob3TLWljef/6qe/U33i/GTYR87JFCxTsL9Pz/1LpK2AD7GUFnRWmya
rpva9CZuf0oijx3TOtz3xfsigJi9ULRBQ3Y4rfRXo35nbPeCbc2g2u9WArYBmSHZ
sy2MtxHytvgVmL9fUpjcq3YvXz4wdby/U2dSssgyyPQwklvFOgOw3+yRVk71Hgl3
bqDFlqP+gtizebyeCTlN5nCbEGrXYvlgiDe1Y9g8xyqMhnOuXZjiBuDQgZAxRzBy
jOCeUspUi/9jUBXVXncc9TOXIQK54PiF/KZ/wBj56OisHuZ2JNjV7VM4vlEpNoha
jle3b0SATtYBEYd+jPiJiJzfWCoqzk2PsaZ4UUWapwSlqUWMOUCg0IIu6kWSPRvx
5uzGTKLyLFDH2dcjv/GHKHmUcnUDhnB3txplqNEWSTxDCJh/9s1uF/yCbeo2Myn6
bjJhGmLuuyotmRkHuwaKpLbkNmBLR4E29a8/Osb6xGz3shObwvZGzEKyuCO5grEW
vlOorrI0xxCVo4ij4Kr7IWF6qFySpX6eGtTpT17EYl5iRZJtp6XyT9kFvAnCQvrC
deFG0i1InHDT7OH7GTQQ+1fqFuvkxNTQdESKWZR2WUsIFlqEAQ41ajyWLnPwjP5E
OUmGXPInxKiNRufrk0XcVeztkXCX1cmTx1Uq07iJi5vDlXI92ncgi9TeOKKlRUwC
rQPOwfGSMyk6mBkvV3uLPl2Z5qAyzOSJnPAvLJkhfsWrGZjJJbfhk0eS7rT5olrl
3VXsxvddSJFghbL4Qu73YQaPjYWBHrt0ofDy/wDal42IPUub1gPuR+tVtaaKxxHZ
kWDRo77sTY58vEMOT4ptigrM8SdKswOwBFP2vra8KJ57SJIy7rF0qfOuv97o9Oyw
W2UGRsdTVn23HdArzr6E5rpPt8Th3oSHtATpNxiTfOHzCcdKxHwQP6FtiWE87MK/
gGiRDyKskWCgcd8Vh2/EcRFC0WFxGpKxvRfZqF4KyxdihXY3Lckrh1wudvYdyZqg
stNZeJ8SOOTrwPxy69/RTjhTRGH2KzJhtnIH47wFQv/ZBhkXSr6mNFvRxfCgzDjl
qteOUT4zyCAYOjZgSjcqQOMqcxthfV5vPh8c297gzoGMR6k2G/QUW2HEZddAcj3E
ifN7xnKh88ZAsS1ekDBFsCq7AcVrEqlCVFnZQVV8b+6Y3oltPZeQVHhHfoZcVOtv
svsEGh5AlVYuz99LbwWs9qxQcebjG1L9pJp/Kut9QzHRtZRyjQ7gGVjSsqsfxApX
Bxe9c722Ln+4TMoKUcxbu5o5o4JoCosLvYJ62F7j4ohuL4+EDerNWy2+66RX7wDU
ZENoj7DXsgnYxxOWv1pns+DwX8jZLaTaVytZ/xQ0U7CIPUpYto4HfnWqyaYVtAey
ThEWpdED/5JHauPV+bFf7KP/RdvOLfvU3mnthk98ol6kdI6kZ8pWopUl68XHN5V7
3OoGnzuFSuEMNDAAN8dfejo05pltpeycu24ZeET/c/uXGkEQ8SX8uGIGxiIgqSy7
e1ZzsWIXB8+Kcv1Yq9QzI+KWfKuPTUYYqP4uqPhNtERIOaEp8TKAJsd8R83yoQJS
YQZXkF6EXCUonDA24Zq3p22Gm+THDYZoGNT8d8tIxQTYuwswNoy5k83bq6vDJ3yE
efF4prpF5jDv2/fiV9+lFp9GE6s7s6Ye6bZgKFi4zC5goIBp6plp0BIi6LVeEIvX
IouPuvpueYg3vXWBC5cAnuaYP6AfNNIiFIq/QFk278AIDNNvuDIaKYIJ/pn6oEPD
7nJdDxv1O+SBclUNR4UDIWzmWF6W/5Bf6YTrbjFmDSTMy0ZF8ZA4DGQxL9rys9kt
bC22un9b1s5p4jgWa1OB/GA3mpbWIq/LeKA+LSqnnAP1ewpiS4B9wWKomci6h+E2
PjPAjeXfd708BYFtDKd/x8t8AS3YywKaEJ55OFuIxhdTG03dgrVTiwOfilg12Tuz
IJLi2xedW58ID0eyOBspPpdL37escPJI2AwNKslPYuzJ9L1Y8qTUo+OcQlFgwAim
cWQ6NvY0NaO5FPqBAiynt0JIjVL6djC3vQJIc0HeoZBtNpeBReb+a8G/tZ2O5luG
ansMnco+R9tpg5iTYtwjtTKN6jqZk4yLCSCYmZBuL5ot0IJN0F+Mg3e3m/rGctG3
RneCW5zPWNk7I7BK5u08BzjfrinVetNOet/B++E1ByBaAsDujxq2kx1j6lNVzZKO
Vhb1IBm0eoUZZtNuRPAV3in7FRsuqC/J/nhLrBMIJXJsjwi2RtPUvhAHMJerS8e2
nos3MlELILeC0gm7OsZju8b/HJJKuLWn+YEGj/MXc2xU41kYPxzKiQuQsBEmBnkB
UMz1LMCERjnCAxfyiA5BUNL6Fpg7fQRlO8z96KJvesS9lbkHQIYxXJBV8k/ZOscs
tjIXSsXCiQqaHnK5E45suWNfKfeENwsx4hMVNfOVR+fo3iwOglNdeIzsvft6g2qa
b98+msQFfwWeY3LZYD96OeVXIl+lDv6fOfUHLWB78NyYUA9YMkXEZYItQqmpmYMk
yKviV5XTftPANyzIzbLPxI2OOJZ/zaRw6k0yRG+B8fX3gJcgsNSDH9I792Lslj7G
fw2sFkRTuKEMKTWvi5o+c4BsS49/bdt8Dfd+ssr+lrHtrnHzWHP6uct7+yrdheL2
/n1M/rxX7MVBNqTVGvZzmW9RetHHTJ/E7+b6JNGuhz3NgQRiwn8vHimaW2JCYEd+
lryxdRnHKxIruhug1c8atOwqTjC3Ilwt2fXvHUaWkKKDmB05JojGcrIbCuEoHMe5
SIT09Zb8NDV9ADCy0bmS+1Ng268XLAEb2yYnoBcA201p/n4pkW3d6VlGe+hueXUY
CjuEceaQvv0lWNc0fwBa9o/Qbslqm9jUxhzFpvPKbvygeL+tEuZVtJc9u+iLnAtC
kPSqaFNZs/n7E2p2Lx7TWjR1Y+hWN3hAiVpa19I5aA33Qf5VdHuXiu70HPGfHM5e
yvewz1+ZJCR8d/utA/wNiUZu4/94rNqt/pOE0Fs0GiPIxjHZ4xjeILunpXNywt9v
gngWhcOcdgDjrcb9u1ukCFLXSqWnZ8IBQ4UHc1hq9nyzcqKHWZCzUU2B/QUqABqW
j/MVwxHb8bbuBLWBCcl7/TExn4tS+0m7FZNNNHDNWV4XcqxZEaJA9tGW03gxTwDo
BDgsf3GbmmY58xhvJspvoAXj0NvbUek5UfjGNDmlP7NEp/p9e1CBunoOPHKmnxZ6
xEqdn+WP89MmWO8aJlN9k9Veku8vhO2JqThNfa2NMl3JddfjVL3Gohl68DevD1T0
BSIXd9CzP+peh1LaHlZg44HMKlqXUdVWKeA4Vk505Nyp7h8BdhYRZde8v7JCn0QH
dbmqCOGqmK3gYgDy7F5VBomfFVnspCxBa3TWjFdhKH3FxmcCO8a5G5CWjxq449Za
rJC7GqshINfYNfykFNlafWPnPlqY5aPWbydHMGooKSIBtPO2AYMUwrkEr+n34cMn
OBODpl5fE0D4184ksEbv3C7l5ZDKcix5Shm5eKTOr1kyQ2bTNUlu71AdPC+7BHZi
NiR+kX0OLMLDK5CqV6vemaFOcddZbXSX8LFqVW/tPoCwtVUmLMmq4OxfPmI+3ROu
TabLduULOiLvmjnMtirA3TZkADw5GNzJzwsrYvqH8oTdBiUZY3hglLBQb3FcV96v
oFHKfesJWiUoX38MDUuAQEyhIh+2PIsXbbReUHs+KRQsgHwQWg+NO2h/aa/9fiCP
bfTN0tQs2llJ4nz07DHl5X3vR50I1XzlXb2QKCYgCKglB1IGePqy8VJyDBZu0ymR
ls165XUcyZU+nXepnjOnPalP+2BapHEuByWnwFp5xHOOeAjnTB/amUXtN2+7Vj3Z
TGl+PgRNYKTpvy4u5/P+OG9dzz7iDL+VDgVmyDs8er9LOErUubISLLsc2dgPc3hG
RAMo/io0+N0ui6TX3q7C/5T6/AHzuO8kZUzZPKJrNEnwNLZHc1k+JJuLn9stq1lJ
y6EVvnKVjsDX2CL8zLfOPtmN+L3dsoio8mgwvUt3R1Y7wt+CHK8KJuD7a79hqqCG
4I1fKmyGG9ejUtGqsCJ1lwNJGbX0hecXC7ZAgoTdnli0d+IN9dosjR0J5AqRxw7N
Ela/3D5T12xupCd18BHTWG6V3t1uZ0Lu1MDroYWhrolpn+/X7MiJ2ufk98iEBzRi
rm9otoRJuyBkZI/SlSf+Nz+0GPJAWW7cipmbdmdPvpRdC0N7JRMYYnPt5yeKmgv2
isahzabqSarjEVBuCLAvfeBs2dsWQ4EBMT5QkgFs9r26iQQeq7FilCDdhWSjkLKw
hHLGTNcC6Jtf32gD+v6PuuzJLx3xzIBzr4WuoQkuAJgTFtdbTWFMJkYyLUiQJjYy
MbkWsv6bcDT7N8WwTLZfJtC9S546wZz3iVQjszcmLyD6dZ3Mkc4IXpImddjmOtLi
RJHL8G2H0tbx7DmVgkUyIzF//76bWUpTdFIm0OMKOAqrWrHrEQGqh77fsPTK3PLW
ZA16Ooyw95MAa75Q14oCzF0neFMcyr3C1oGl5hl2c4p2sqiyr5XoE2t8+Gco3Woo
xBwvZoLpFvFbtKL51dnUK0gkKPzaRY+M8OvmOpnzIM/s3FFfYsCgYELb8UHkmXK5
1t4XZhFoHKJlgrhz2YOJ8DKKg4xQU1oFS/xeOFDx73FYUp1SzIms0A2ER6JVF1pL
j0rzLnlEuKWBHFovlj5w9ifmDfh/aEhGOP1m3iud/ARogf/Bok0nMeZOsObf+X6A
yve01wdstuvDZLfxFmKVpdPYmACID5mouQ1y0nkpYkxO1B7xYJevU7tchsM9WjCY
7sMWF2gpd7lOxLRYgNAeB0TdNNjqA8PI56iX5u2JT1PP26F54G5cNCgiBfKae0Pk
MYQ6988ex7zSJ9YBI5BxYwhyVR6N+I2gkqB3wWGppgwB+gQ6FxGTlQy9vtWGnRLW
/5hzSSg19YB1eQqYNp884wzY2KcbMve/r/O1NbF1j/Mb59jics/L07579OJ4AMio
ISPbUErDCGCieaLs2om7456pLTqciFTYU4M+nvBJF1SJFw5o9XpSa16aD/NJiv5c
+p1Ehh4qQfOv/9qQE+ki9y9mf5snPZEcR+OpGwMRxB8C8pRhTxL+a/i5VLfpwOT+
GE4s1BObI5HhIh+YExs/vE6J6G4BUe6RA6QRmRwzE8jsG642Hr1d1UBnceCO7N7R
UrGQTKiBCXAmN/kG8ig1zL3E7W5Yy/X7eTF9Y5xArfZ5rQiZlRvqCI1PMaofyprr
FMyMbGZz+o426lr8fq9kL1AMBLVU6tv7qj/1vDxQkbfQtkZIMjbE9Rq8hvpIldYg
jCULE6DJWEBEyb847D/IYo4jUJe+68SPUiqqQbWt9bP2ilXrHrHHzqA1cYlT72WX
Vqc4nS5NzFJs18dzaaloxGI2OxXnjlh1/57KMNQ3aVZNPZqYwgsSeT32wjPvbO+B
e5ivOIyrQZ+Mb+i+JVbcbuczGHoAjLxRgRW8XlgSldqa46aRoPQL77OudXv7dC7M
co+3kmhiFJ7rINecedZ1VlR8v877mEn0hPnLsAfRMfXcyAxwnFRaEZIyYtvNmCt2
V0eDFu43DetgiQBNGkr1eccjQ+KmdlRLdXqwP47XG7JFL3a7J8/Nfsps405M20py
GALBh54NBlJkLYn8vb1MmL9sxBRD7RLTEby1mS3HCcUS+zdXkvdlKaP9Ua4cMUNF
LCxspdq8tqsjVKd6KZAl5ckyeOOfjWBn7TSolQqHrv3KBglt3e1oF01ggzs4yu4C
NF3nrNPs2GOVyhvPQEORkZCTF5NCrn5lHh9fVjk+DkLrYiWX34AYrmAuNhew+pPh
kMRfN/O7QATGqqhmIjIg0oT5NaPMjHdrhRE/c1lowwMM+i+SSglQjlEkOeLr4EJx
Kq3KB7StLNd16C67hGI+unv7LRLZDG40MVyKSRfGG9zZLO+jPini4oSFUqtFXyF4
EhePjgf5oDVmaAbZ4B4rhe3cjePMK+KqAeKtVJNRej/Brl2Crn/SgFVOV4UuD5bG
+11+8MqgcixZU/uEFcocuRSHBjJ/lE1XRn2Vd12zrJiBbvFPteE9g7XJy6xpg9S4
XeExbvTwlG5jlz4sZviWGjALUvEhX64BvfaXuIrhKq+ZyPdq4r+VA702klsS7iKq
6RkVhujBFekyIzTpTKtVAFtW7KjJ6sUMB+VlBngQDuEa8LPuUUUHFbHvoow8Xaxt
7LaClZ3dkq3RR4/HNhZK1a/vgUIEFNHuSR+mSYWf335ZC7npI0CvEZJ/rgcwoAVQ
F0P3XvW5kXA2TbHwBps+3BkfqPZhSU1cIgfzt9WpeVewPWMF65fP2lt1jGe5AgV6
UaFpB0OPYecw+NoFkHYATIc5fwf2w62aQaOXC67BdeGIL0jJNeBTkh+l20zm05yR
iKkM5h1+WOsfXrPGRgQMaxgLvfcmUy3AOMTvGQ+av3lw0+YvISaTr3UK/AUoLQeH
hCH66J3fxt63ajilsIw793SI6K56hGF+x10KLcXfC4QMcMn0iIS0eXAJb0daC47i
MJS8x8SMnY31G55GGD+Z/HXU2yLs0B+v9ndIKYFx1AODcgO9tqSnIPv8rxWG4ftg
Fg/GzZ69nenc0NtkNgqTR2Kh7Ty6n6NFGKb/5DgtcwmZ+EaBYvbTM0q8xSoA1vA/
n4eO1aWK2hBizGsWkY3MpUYbXhLMu02RWdMUXsagUdwuUeHXNsFyTesZSLNld3t3
CAGhao4mJeJkcHQa2evGr4haPb0VkdD7yMMWGFh+Ll7tNfoCsJRpJ4VO8jCLN2HF
zbBdFJFD7RpbPizyj4vG9OY/5ljofZ43+52vV1JvPaL6jHlbzX1F7UeMhfH2Uy2O
+zMIB6ytgSrt1ppC3w2TYjL85J2sqscAeKvWAzhPnD5tt35qSOrM187qWi/GZ3aK
mAtijlsh+oMFM5b5OmAzmW9zJ2akG/SyNqSOwWXMTcRPk+LJ4pXt21jRDLrpVxtk
W5ODineLCNfl5huAqo7eIiUtdx4FDP+yHLGNo0MuSW0SH4LwVwSA0WHsPYvwOWg9
qHw9Kl2ggcY3OFN5VwHdZMwVxRPB9rwwysJ+W9v/Kf9AQbgnljjW0Lgkuk48mMEz
4q1xM0tIsRWRZwkWCMzd1qG9M9o1k3voZO5UnfrFNoasNDAI/1upwa4ZifGpNDwD
PTDpfYaB7L6khOFSIcUTB06/bixWQ9ew4qopWOL1Rrg6jxvTElBojBmJffRGunEA
6oaCpDjzs/NjiLrz/XQDq2ghc5XiJGOXLey50d7q1PQCO35OYGqJ3uXg8cxXOn8N
ubzTFcC5czPHAPPPxX2t0YW+Bv61aX2MmAqPqwrqWPvqYzGnlQ24K4NPIoU4oHcn
Ebz8MoP/hd2HNLu1JeYef+vuf1oPKxW1mp06BABEa0ARkrl3HRCjJvLGZhok1emO
jg7LGBwJGz3P+r5rayQnw+Rn4AldSh+q3uDVVSSkie3s/PirYfE4xd1Zk/ILEJhH
hFCERhG3U2ACZktNm0PqKFqmzxhx5Iz26Hj91y4m40NSbIaOppK0NvrVKAXEOOxB
BPdfWtg/eU6j4eDHyn2ySqiJNG33xuNCMHCgmjk378JcgM2T/4za/Wx37RzPacIP
upkLtweDUyTjvX3NYwwkTtTwUbzAaDmR4YV3Wd2l2Xhjqzv508UJ2WWX/iC0rLKX
ZsWF9383yu3q/0UiciZyxph0FFq1L7vceG1wHvjD4lnXQ1HXJfo9QiCgjJ6EZwRq
TJGIOJA+tEPudY1HcInQFaKsneEghdLLQMtaVdJ8wAmS1SM7vT09BAm3PBtmGG3r
7F1ijneK6vwl+YFcpyqCuHxpt+/IyRZPz3gIFYDedLVeaody6vWdQ4/TPLXfMs8I
I+zkTlr26GmYOVEVc5q9GPTcNo91u8779Kq19H3/uAeQ/QuhDZphSZ5kk7NBtJVE
4Dw1PzuZ1LrFHa/f3hgER/PTkUKISFO1Ube5gbDX0IrlpNaJCgwucwSjAV57qCIp
+Wa3gWIxuerXfSr/DHGPNir4duNRHP9sm1icdhbZ18JoxSJ8ziPQg4EZ+CjNYVYb
XGIrR2rKEyxHcFrkPekQrpxGe+wEu2AASoBtnPL/Q+uV2SzgX0uOz1cuqnDvRcru
Lp3KdKMYU/fBOq9XDjrT/+iFRkgWkPr6yHeV6loSS9Rk/yjdoiokq52mZkW59AR+
I0Quq1Jbu2hedohMWCZaKpXtrQ2Ovx9q9mNlk6aAO9J+ijJXbLBpp5GLf3L2D1rY
xUDi4JBSkMBGjLZJRjS1bugmo+ob5pLXnUZ1We+3BbKRmoX4p+0+W4Mau/K8HU+6
AMBsq3Ly7o930u0E1yZBd9jtU3NmvFc7+g0mXKNSeGslmNasAThQls0+lM5dgFW7
PbyHYVhb8VXBrXTOJviDYUZOCpUF78BfxEENDGLZh/Sp4BzX0LiEwjXMbjQ3dGM0
xbo8UgDEvk2d0YmYDYl7MfsawIbqqYETsWhKSr1HKPTxQ9+IqFDcj3vyqla2oq7h
+RQXopHVu8xmf6oz+yCssLOgjE92fKm05bSa+oQw9SHZIfDMtiWJU8J6RAclaPfV
XjshDlcKFrIdv7k6o5NbVwiCEbgyEdRkMstRpc0F9OkNubO1bJogL19PiQQYLjOR
G3yl4L4ROGgMSlzrE6PBtkDOkhb4lRxka1LkZQZ8lbuZNMpPo0PcT1uBJva+vPUg
pnW7L57jjS3hmq/te+FhceJYgUJADUPpldU9agr+HJtK6TyWCbT/Eb6ygOkK+apX
AZF3QLFErG1h0QYcLR0HJhTkUykCDXpxiJw5iNm0axnIyLcsSs628Tr3ARY6r79v
qp13pjtkunVpbsmX/gOx90agdqybBoKVzuHyFS/NgyviHBUY/mKHY1y8/vE0AU78
XPihucJxDrMOWZLBt8cM+oSr2RWhxQ4wDZmQp3GnFo+7/0xGu7x/cI+6rcZHqrK3
piEzkYs/MIocXTcL94xpgTlf6czVoKMLshsTGW9U/ygw5jbeQs4kEO2vjqNoXS7f
N/J/f/pHcBBJ3Ec62d+2F1by7UrOltM2/GVoP/88MrzSeSbap9fzRZuSrtS6S8Az
yQLFnrVbJb8NnqeY1G/vH/FRMWQ3/Q4VdMIgtLTUNh5Ux1cJNKb60QyYDruG1OGJ
zEcUyAzgbC47Og3xxk6r1iX1hF1GLUgh+IGmAkpSh0NU150BmlU3T6F/kABHqBtw
oggkKaRNYmim7XpVem4TNnBdDLE9xCORXMaAQSgzojCWPV59y8KJiNkFq0nD+sCr
pRUF6StFYq72KvqqpQk2vHYJs/FvJbsmUZAahk7T+jvEM63CLP6F9T9RMQB9YgEg
9DFIDuviua0aQM9XFfQ7PLunwG9Z8rJeZWoWZ/1qUa9rRh0qQ+3x8G3211yeKjo7
emJO0AwvPz6FA0meWJiUWAu17eab/+SsYVmSNstbSTfRBpeR6BxHbsfd/xEU0cPF
R1TCsFyk04wsmvSQSMWt2ZCj0WdgDODWo/tDqSZj4xL3IX+lVdQuAseqxyuCKV5N
7MBfQ7y1R2PLb7GTAIsZXO521M5sWKuhXSYyVs7VbzVXqQ+14krzUynSyn1TIOw2
5nT5g9oLPXSLwRsGmVDytNSzLYTc1XvPfsOu+rJH4sRDuT07vJ6fZjpyWJbjAF9e
jS6lsKGgrz7phS/JKq5w1ICRX/lyHLFWKHMO11Xwx88aa/c1lxKlDcakkHmGc0Jk
P88/GTiNJ4mAmF9YpgCjxpDBa4kXwcGpsaV/3yfJClm+BiwXH8GohEUYGqM/84dM
pAkR/MsPIv3H5ykOHHX5I1ulbON6Jq7ALlsC/Ig5y3oi3R7/7v+lbpE68sS5e3wa
7UFHg3XreThudo+oowM47umtXfiOAXBJEf1xawZq61fhHzw9vE2ktgxtbUCHdihe
FfaYIuIAU6QaI5tMMoh3/jT+/yWDlTLutPa/1gtOvowxQm/W6RncnP+RBbS1pNxj
AyyAIVR2slgdYaKHsO9n6qlGoukVSV6+UyDRJ8kanaQ/EkSeieeLS987vjNQWQsw
2vjYWJfumI1EVD6ZKjnJ5ekn2FGyjKMf7Gold1iMb5zvB1NmojuXuV3UhKYbbDOj
uQerimOqN8vpW2sCoHM3ZQ2LhK0s3RfMwnlSatF67c3DSilyULwKKjHeUDGuXmFJ
GzbOn+eESy3vJF5y9FUg8aAWMf+CFpo8EqZCEX5bhPmjn62sJOqeNSvuzrP19Rh7
E5Okup3TbDfhaa4sCmZpctp8HFw5N1gXqQ4bs9Zqjy7d7WA6oFWU/KPa3mC4amGX
VHjs7DvlXdL7UvQduMzVgphtefZq3MIiU3m7RX2vcvNrwNfu1pih2wTFaqRV0Nyk
biV8JxnnfH7a2F6raU1ErkFs3+kgB2Jrm0INRBjHpV4cjGTP+GNDnWXV+dBTx9li
ZwSC0oepSb6k4XnMOtZZjgAErROhOtL3woD7FmFq78KrfDpfa9it/pfXPvfsUUCQ
4chg1NCRk+haoQ+j/j3aG3ItBedFk+6CYQ9EwNzY8fD8txUNt1HiXMXFRy//MYie
F71eI1DCzDhjwTnZNEcfGT6gR5i5F1VqbLbrmxxTE0gU5bLCuddl7lOQaSIqDaEJ
YZPt5sMiuZMb11XBevUxYkUymGG8+tRTNBHrCjm4F74KTk0kyXKY1Lk3ZxS3FIwB
WCtCSUUTXKF0f8d27EGwkaYQjx51IS3xeUqsU2egI70sLnPNDJXwebhNi6ly/wuI
q4+jHPeTBzAdFY18ys1qwFU9acjycXrSXfoklPuPd2az4AexIlkkzRjIj0MwslRT
/1Ot4Drw+/Es+q3nzoHE6auhKSP7FIUKxQdAPEH+0e6Iqiynyts7AW6WDAp1+mW+
46tQIx7ezltWU+XjpyWuz0GgmUe/ypivKGj3osYBW9WZOeO4wDyIqFhhmko3mjAh
OeAApjCeEu8Qu04fQHMHP++iq4AAsjYdmej4mMUM3e/slPsRsfNi4Li3nHk0D/jN
IGWo47hj7J02/1SMSpJLClrqxK7J3QN0/6fMM3ECV4OrPJXljGZ3t6eBYs8w7BVY
03T0sJjz5uTzcmU1FTpqokxxsc1yN6wPcx4TOu0KR+XUJJ8OEFtoRrl1XK3K0WGV
295BCTVK/EjHaitwWlSG9471vRRLuPVPjyyaXYqnTK/QCJVltxXqEYZymIZr80GR
ukULwRRj37lUussnyloMVRqIanbgw1Xb+x3tE5vi0koEUudl91C6R00ETBzzH6ku
Um0HkEw24WVKQmBRXVLgq+6MKn/n+YTp9LPOzYToXundeYW+7+kD4dvkdzQ3/hNo
2/mvlehqRgRkwP6Ss1BnwQh45BjSpKrG79fBzU/2qiiiL2vG5RhnZo3xPFnjseic
D0F9biiUC26LEIdvQovM1GwK5p4dp6OQXSwBRppBrPtEOolj4XH9M2ptRk5/6SUL
EQMNL2pt3JY9ZYLQ9dOgv/iz6vHiE9ekMpnOmgnrZ8KsawAdmlaFUvvQIE/WCFLD
btHYIRLL+ck7Yl3ecXdO1zuLrB72U+gQgWEDIkwgDv0H0ULUv/V6NbdZ8rZjmk0g
Mw9ryYjuyMCJNSKfINO/BRHYM4Ixv1n+H59+8RYLBxQuOb40rFBtMg29sG5RpiQ8
2Gm3hhPKHaBMjChbAdi/njvHYF2x2EnW+y2BcwYf/g8pPOi98+RGu4zx2jeihSSY
a+LvvGInroJ48OdnGWaT7lwxSU2p1U6ShvOT5SmRX7RUX/+qqKeXSAKCcxR6sRLW
VGh3xKrn/2Oo1F78D/JzMWwpldwieL7ttd15UNUkqzfIl0IgCplD/6qAL2GWTAlN
CinSWSWjvm2Y6OeAwvvW6MWTC/KEXcoo97W4A3kckCZBvCN35sqUCMeNtzeKamhI
8GXvBvS2JCPt+8RWfw03fGqvpwJdbOoe472PmLVcyn32azoY8oMtMAqrQ5FG84st
YnA5QyGtJ8xIaPdCUKtrHFFOgDSz3g5EGzsX20LEEqZR8kB389PjwhoVrmfF37DN
Mut2gNrePCkXUINX3vf8aLI0hWB1lRJOzhRSNJr7MmwAD46a8nKXSgPuHCr/RlaG
6M5wSjnWtcFy5tkRVj+eqCgy1B6oj+TuU6FuLjQ0SBbgZL4byTkw4ZWlWL50mBAP
lTxhq3m4hK9vAkWDVe01uNl5lwlIbOAfLSrQ17j49MOEg41IiFL9RaduYTIr6iXC
68TioOCZwoOgv03ZvsoX/bdcEkekf6jPJ4o6nY4SG3O8OD60e6Fb39pFI783jt5A
2kMlbt4FMRlF8u3ST6+sIRLnSTKMK7HWmv/K7XaIu1+XJ349NObQV3P/46ECYXke
n4i9Fx0mtSr0hBNz0jHDgjcuhnhC+swFb+n93W+hqVBtJ9oEAfy0xMvO9VDHlSqA
a6U6aUBfcg1sFVYFSOtRXUmpb0+4CRB0HPl0NH88aN3eHL3MaSK1DTVW14Cxpzzw
28XaBmKaOx1KxD7ogjnvA4VgVxtornB1+ZfCHUA4iBmpN4u+Ukgh9II7MEODFPwQ
Golyqeiq2GZGvapzVrkaniOE1DWOAJNHOr9N4dp+6lgY8w9wpWQhGAAJusl6v6Wl
i562Hg9cZUhabUX0jZTiyOH+D4xvsI7bFgb+wCJQZH3KBtwYozvCJl1tHwAe9gKA
PfpF7CpaP5ZIRkW1ufCHou9zMbEZpYGt1svOw1nLHVe5e5fBGBFDxigM3QuaDU82
l4QDmfiJxmVF6dYX0xvDUb+oirzy36wKbGHB1SHDKjv/ySo8ckiYWMaXSMmO5lTU
3EpZiNpqf1NiRiu5flD+kqwi9mk3+3cnSJEbKDzlcmmSf+TmgsTJ60CRzqsia/4T
7gu4X3sOHViPQv5KNTLft7On+Dr8Ax8s4a0cXFUSkU4MYeJTXwAvZdSp+j5lhW05
corFJSPdTEnk7V1aGG+mcOhBJqwwfocH/ceMgdiRL2o0KvkS2X1EgTbN8n34g0jh
h9yWhliAjjwBtVMQ6+M7+gcjR6/FPXvQEyn+4Mi28aKbkr++QK67mgNpTycKrqDa
G0+D7V0pKplwADfDPHd0dpH8xl9TIfEXLHcHizfRp9SeaGZoRW3rInTa80Ii3cD2
+cKG0JGuVKI1UGJbZ8S+Qlj4hITkoahymh9O1KgKiZmzstvIaroFPBL8BsiZZRoZ
2+H8sAu+oC0Rgw+0uR4TjRC6C3n9R4Jv1n9GWY5bNSsuMAnqxT+BmFxOk0ir2xaS
InqbQ50grMD1EYX8+4v7jKiCrQyRmgtDkgmvlswiaiAlB5zseHROVJ/Jq5pRGSM9
xPM9cCNEVsvzpcwPiz2ekXIK9oEHNc0f2E3fnDonBHy/YgsGsroxiAvmTg16pjem
C7pyvB/AyBKUKgL1KzIWZEC7Vof8lH0HT4KWA3UndO7tCN+hXAtqJEz4SWR88i7U
gb2m3mFhMZYJoe2juxaNWk9o7aLJjsoTlfCM9cAykWYm9D6zcS+keYlb0bJY6U5H
paQuezF74n5r3cwOpWy9wPktP1fV1mhFSZtdjAeYT2dAHKTMQiqxbtnOOvOxzwhF
UErve+ZejEnGZ5LiDeHCnqL+ge4VG0wNHRYlBRLykOpTEpLfqik4U//sXR8Ckuvk
UKi6n954cAvpsMabjI9ViOCvWb8Ph05BZ7AVdEoH3ZQdPdTNTssIOhu4fWroyH9I
igOXwEtJTFBLfGT1eXatHsc+bwb1sEP45Y9MHgIimxNAiolGCtYhF5GVxZsPIDWM
AfwEyB0inBwHWz6vkR1H3axTpSEDjfeaWMd/3ZPHsb43/7lBgebit2fVDri+ymU4
sgETMVqjy78t1pPRmdzSTtHA4/EZjTfMgTBE3HlzOFD0DZJ8zT8TkrU4Qn9uNAO/
ABCrVho/1itgwDd6Hfwvke6XVFwbjIhexgb2i4Y4E5pPVMNWJREU79b6DaNSnyYQ
9SgJt9JOMWlCst8Wy851/tXrfrxMv+yIquDkDrI173TOY9S9OyU/sgMX8ytg2mfT
f1IM39soF0faRwQrfYzKMgBbC9ummtKjF6bk6IB3AfdFgjsoDafDZ6o7HtlQO8QI
3lmEe2WyZaKtyJK4rjJVEbQ17OOVnBkGEskApUK4LV7u6PdgFh5n/+bxnvOByx45
0y+HmAPoZlk0Hueymbk4fDm8bjkoA0mflyrGQeq2aW8YpuiKrB+3ujTxpQyAzgPQ
FVa2DKtMIIsoIV4EupkcI/1Y1thrmBnKd4bYFkAtSCZn53/Vt+cKhcttp8OA3nJI
+9lzKzRr8e5cwN6qrsYAf0AdfTOXsujceN1WJNwap6TIY/zQzj1mQHotwjpkfmPy
YOy6BD5oz7UKVmuIkswMPrz0o634R3CcFhacFu13itxmh6At+u8pAInYWyPwxuZX
h+yr4/IqPyo1FL2l3IYORz9L+dytizMdjodmyl88XxVfqkx/BB6C0bBnuYmExQY0
9MxadX1pgkyST1pe1NdR9ljlMHrmq1XzGeibANbtl6jwKnum/1xMYugdneou7ZAj
LsM63Ix19IEhuOCifiq8JcHU3sOIQ27jnS7oaq5ft+GzXZqsxjdK0PyxZ5EUNjW2
kp3pAWvDN1nrYqD089SSherPuSkuLRjtehjslMNO4OgB7o+O5aA5VsSdPB4pqfSR
HJAVg/xrkLFi8RNDA5UE/tiDpN0E9bhE99GAPa9zaP54GmvsNjz3P942lyLvNJjT
Wi4QkkwB91lEN47FqsdBuLmIbK+JunIKIh8JutexX6zn3+Vgw7LfFn0piApohWnp
WD4PWQF0Te2dqVfshtZcybLxxap5K31QD8FUKAhvCHAQdBO58adhkBHK/BRC1pCd
O7aw9UrcZ/cysIM64U/+yoYrnyueUXeNPKFxQny6RmnlymkLz6vpIq7WqEMFG3P9
5KGl7+QdZKQH05HhtM6zBkmEpreCREVfn81ItZhNVlASX84x6XswIVmMCm2Y378Y
beRFYsUksSM5Ddu1uRyXjOwywGglEkjQ6htgg+hzUub8vm6wUfCgca2AZ59u9WhO
QFyYvr1gk88Qu6sCp1pNlyuBSgzu2KUO3EA0iw1Oza3u7+dME7dqyuGJ1ioVujj1
ig6XeyfnAHYkTRqDxhBBGIg9ZQdFi1epzjcyraoMMn1LR4LhZRftQTD4N+XyXC/d
lto/SiaWmGhSYssixqVo+WquiZDHe64yu7P6Nch/VgsdUX1A47fUk4t5P0xcz5iJ
1KJqTSzWbrom1+H3r3EKUkmYOJ4l6ATn1eOaMVtu3pFHxaJEqiCH2jfyhOPE2RZ2
TIadjKITDWQKMMBbdfrtoTeknGRaQ6qcuHtHO358uvd3wdTgl8d/382Kyucn5w39
8SztrVgvignVf0SKTICOCsvC4oxrcjwk4H56sDIHgG8oCsXcGxJpiN9AU7O/hvxl
Zs/Ll7915qO3D8xj6WIrgsvDLkAkeN+j1kf961yRlgicXi23KaXUvpLg80Dt3ear
2mxE1uGFQ5sEivcyWzLyc3fYe0tgT8xtSALB41WNPKlV7m+duklCnaqSVtmAWK0g
S06G3qzWNJ6UR4BfEctXUz73cg37qi+xraxZNnFCGwXdQYZhPqMnfH+ouuaHzs1V
eJoKXS5Ypz+qITgLUdWmh77AdaJ6tDdjVSZHD1lc+fgBk6PHRoduBMnJdJDmF9yu
Tjh+3m1047N4Ip6JecfIa2h30PzlWqru/xSnGrapin8IkXkBlfUEXwi/s1wH67ca
SJm33/UIBXCRvRRRAEDZy26EdTxiE/aoTHunA/eVmHQeFayW9IrEXe1yPc0FoKpD
kw6KZwuTifN4LtxUVjtOPxVT+X3dvsV//N6GIeXMUmNaqoZHA9iCPvMjH/oRDn60
zLIIJAERFaqEDxdWNQb1hhSmQaqVMoxnQHrlnSmSc9PHcgocgJj5GkV1eixOEwGs
ouvfqddDzrCZ+wrBPErK9U4rDQgn48gb225YEtLOj5bRrKAFfG5YzS9IoHMnxAn3
jC0nL/gQmBvAnRXQJ6TwyWt8dD63QqCwhix0t8U+tmwWvaSlr2kkiWVNYnWjQSDp
dfWl/YvkMConRzVFgzUweo26A+/qyD5zme8UOj3/pIPJ6fFmw0VVvPsuhhPxOAub
IhnP8eRCBk1hGEvd2A9HdhRq7h6hR9MbYYAdbFg+WrqgR2cvov/0Q841KT5xkqL7
pgbODxHtbUera9VC0Blf+fSA1ZZCbyCgLA8apFn6Tgc4f1PWPcGvMIp4wbOIFKpF
pdBSHLegAPMWUoRrZQIqKe4Z+tqi8e2f+P3lkYrW0oepUyo1g7X0bJvuY6CCG5x6
ZvgZqyl5oo70BxDkRVik0T56xUL2dmpJkKXgW+TBpefu7h8I2LhO/5WgtNqhmW3o
LPz3ffOZ7r065PYB6XkwWVD32VswomMg49bnhpotpMbxkC/QFeFBnwVaX2cBdT0r
YVMcNqR7eSRGm32Y0hLvNfB+/h6rUhvIoAFsLE1sx+QTNvaaRc3P589QySTIdv3h
Y+ga1xRDG2VJ9vPfJfgvzZ2Hvvd6+3rC+cWgmPLHYBZYCbpPol5/2Iclzi9Nigv+
Yrr2tJtOqYlzLzriIJj9x9KBztbnNz39O4K2zCIwChXs7nQMKNgUS4cjCcGZoqZi
cLOLiWGNMH1OySvoeIMXPLAjmOmV+alHB/Zz1bDkjCqZ7zHsSyZMPwJ11Siowjvm
GUfPO1Fgeijr5mKHit9RMRSt0mvnZVK5SGX7au0oH8cpow542a5WM6wCyormlN7T
UhqAI51zQ1ye1dgkOp2OyPo+o5ZNKeYgnI/7pzBrtCE5LVpNjrpF+cAGlLePprJT
ydL/7tHswoOK9nzUDuhm1Q7QfTD8Zf/r6eTkR+vuApSOHPgKPtvDygr6lNUu9Pqt
XEl5AoRVYqWhizTnZmgYqEJImUReZxLRa/37DCRJQy0UnIrFl20/h/zAaA4EqJRT
6C8UJcW3EIFE/HuibJ/ymNNkvhn0/H0cXoZF8iOBifsdXLs345ENJyvmLpftCC21
8BTC+3yzAxEPoI8IFmRzmhLPuIYcKKRR1o4SQAPf9YR0xo9fnORRAAslvfULs6vr
gMS0vDFEyAllPoGlsSjT/OSn3C4HPc3sozxdzXzJbarf3VtrNi54nJeFB2eGeTNY
25+0ogUrwWwVaaA04bKzjuuwPClN7kfXVyH1Zw+kDnrdGdY3Q/Fxn2BOfv7k/eK9
vNQvsJhsDQHUxnDmC4AMiCyTeI+YGStMDr2FqCfwFnSMOIw9jc3t3YKaYoXiTvha
rmxWrhT2jOSUjnFxBd+J2hUgepUgOZSudI+a4eQtHQOXT3I8NTW0gVo32ENyAFYv
M+R5xaljsdKeSFB7zqpaDK7tOy8IiWPBuvRMxVXfv1Oz741Rt7atKY9I4JMjK3cN
NQHwOVlpJzWKJVNL5QlK0viENiQh6opVh0YPVwEk2IdOe0AyXNADBHZzJhhGkN4E
e2Fjyk4/qPrXsy5B0HT3Gfx/hhRzQ0xI+KEchn0iy9wGVVZqGBi2bGsOo2FLvaHs
pOgy/LxTa73xJjDOgnWpl6hNJ00kiesHBN2qzY1G/OjT0gyedTC9SYEHdQzL5C4O
G9xt0wsc01iR2igIBibjaB0ZMdX2N3L8K9ROu5HNsYQRAR9VlgRFd+rB+5ec7l5p
/Qy8ZbGOjCKQUyPeEMQ5r9Fkm3+deIcWX0ckPxJy/tB7BDaQO56WBxF2hJ9I0CZb
KqSw6sF9+/i7fSPJ5KZPwE4hv7YB6P5V5txZi622xhxk/Nq0I3/FrgzyOF6WS0oj
QUr8RVCgec/bOSV08bSYrAc87wl/oBMGx69BZQrTcle9jWMt5WsliYKmbcs+oBWv
SPie9+TWGGhnboriKyxPByUWglOwMAkOBUFLXOhVRcQrth4h9pIr/DsXhjtnnKsd
sraEgjaEfqNm50mjFNvDbCnvVNeVf5/y30pMKdQY0tdYVQFyhC2RM0FCqdNiCPrE
mwP7RGVkz/22zqxwLUx4+6EUREc83Y+2VpfVKnFkcOzXnktkEhWdFGewVjWhnuI9
W9lGptdXwchR/8O5k8Bgb1saVzJSWQwiHvg0+NTs3izzAwJ4g+U5/7HUMN7M4km+
VgAvMt1VYXLp/wcGA3wx39XPH0hLHaBekVsnX7VHS1KhDy4iRMpyiGEEh/7KY1ec
Y6h5a0UoWAcFLJZYjPka3X+nM4uFo1T+dx5NYY17U6fyeGJTZC0loM0lupiuP0CK
Mp5Wf+E/R0KdzE6+eL7TXJCNVunPRfenVgDTd93HYGcru1zQ+IUiuI/tmstcIApA
PQKI4p1Ik41gsDvP8Ui9uCaV0ov78F9Ir8eiQ49H8eSWgJePidMBGshTGyNUnF6V
uuDl51vXuLHuSxaK4FkrxpLYNk18++ag4XswH0NB7ydS3NQkaBFr4Qbjg8m+TWNl
UEe/R2+Chn9aTWcL6+j3hH8aRtACLvt/44hOQGO1pN8P0NTLtU7AfRUX+dvjbaTw
2PB+B8g8flJjsODN8H6Dd86Xdbfp6ks/xC1SstTEFfMlE1kNuYiVxTv0Ku3l1FrH
H0HdaHpnnWGriNttpLl9bKHpGO0bzgCs44lYKi1Bnf/Fc5NKnsbkvQqQvwo/Jumb
nJjnu/2jMcm0FAPc7/9LjYwbedxrNvU/w/Dh7BS8OjV66kMd5XCcTUMJ2NvXJxA4
3migTgzr1jnhCVVZboHkvQEblKAYXTzUWJrVOaR5iirieHWEbktedRRCUtzvP4tb
20O7RzRiNLFc81K2jtqDbA/7Bj6oQVxqjlhtCCpsV9mrh8Jg6oFkTcA8f71d3mjv
pXyZtdDsUsrAls0nKqdijF6U71H4kngVDLG5hvdIIOVEbxNW1k9/x4M4jker0fp/
dzmIHgCpJZ8bbgCCBGsixXR4vKlxpPr7aySNQhxW33V7/mzkoNWTqnSy/VXZYm6H
+YSyLMkex2LUslLJrihFu05VJA0OhlDhy8OSS1zNDVOuGcHJ5nFn+BumTocIuQg0
NFS5DW6JFmM+VGvK7aS+ktvB/IiVRGV/x8r6HvDGPftV4t32GeeebfxkJLoZ/1QA
HWafODOgfKR0eVOZ5pUtnEiM/GMyU8+8R5zNoe21+NLCvSy/CYQuugsuYFZFNpZf
PwcTaOBpGQQ5MVIXEnFNo7FTgKqs4EXF3alahDxYLLsrLisOBsXxv163ioMWrBn3
kHME+CvElpl18zWZifSxFD5BJIQs9v4c2cgh3qY5gDo7WyvwLAnoJjkjbwxL1+gS
qsN0BE8/CVRU4nii/xLwKWGcgiCDVjbVbgmL8Ni2PHfYrISZLEL+lrJXBkyTkl6m
opnZV5/abbAVo9WdjYvtZjTvRJQa2L+eh5mgYKFqlUGjhrVrLUJQMNFCBoCJKtEV
a1nOKe5NEOckmHdLjjQr3Zm34zaP/A05ITox3OU8DclilmsmnU9uASKvmOo79l4q
mb1Zji+TKTJaklRPzlQ5WDY2EaHJl8E+2oR90ZtSQol2KomVxRbJwWQgnrBYCfbE
EwEVnOpoyeWBil0MIc2PPt91e6c0y73h9ximZIc40Pm9ue/T4c8GNGXWg4eRhJZ+
aUUgxf+4IyvYaHAnUAvaWhZJNXBGUUl6MZXtroysRhOdf5ogp8cJvxkp6htsvz9X
8jfrtBvmG92JwqnN/vbgF04L75PRKkxCaMOKGka4tQGrvE6+Ez/6OQDIPR0WSijv
UmN3Ebempgr1+rFena2xeAeU/UYFkGwGfTSxLXP3vh7AOgkNfyu9S2kueJbHHYS/
hp/V6dZjJzLhHgOCQ8jsIRMhOAjHbEetN7Lo1+UM56h8uuMTTBeKDTn1GjdsLL62
D/u9U+4R5WXALNSebEoJDUDb9WwU6sFA3tZrncazLAQVOL3djB6DW1VAaR6fq++k
XHMNNuvlNmDNPcvZkGcYy6jh7A92KjGMbfRUFRyyFb56umbjq7/klSQI8lddwcdY
cCw07JfnNQxd9phH7/KuCOwN3w4ntSNbFEiQ/iwS0CHwZqEAYlb+EWsBtLCFuay+
yvM+F1XhWudnPH07xlK8boO9LuGrkNaALtFaJ4n63pa/MrPZ9NhlI9RRyxD8t8Hu
qByn0T4ulrHCwRCUOU7LAI5KaMcEVxh+4xz4L4eFn9xVRBVJGlpLCJ/icONBnmQ8
u6CxAwUk+JGmnbe1fqVIV/xwNyNfHHJRsa8P/8DNA8TK5V6+DtEefqVv3gM04/4R
nWZI1CTAkzLgUDs2xNpIf5AvsrspGSVlhNEJOLHgWz5Y6wELUwBQijuC3Tts7RH6
BCT//Vcol2JUI5Lp3WzXcj3d3l7txECk5SojQnnkqbIzkheFZUD+tQfcXTsx/yfT
`protect END_PROTECTED
