`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PnLo/bBeOHd138aFVXmYr8pu5Acy67vf3QaHjd3tZGKNiECrQt/RH5oNp5MOGsMK
4ZTKC4vXAO2Pw1iJYJk0pLo0Sy33AOgrmza69q7m2mScHsKGzqgEcMquq4mI2DrV
CMO69FqAUusc2xzKxy5gpQHlq4IugZG+XtPbhTpqCLpJ/BDvVa4sol924Sj+9Yoc
vtCymJhSB+yw+EGjH+1jur4zNP2Fb83i62Hyvk8bxOzkQHG+XXNkT21jG9x84Ryn
W4r07UVjDf9YNWUW71qTkQ==
`protect END_PROTECTED
