`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7U3ShrIaUyocg7/LahnXwGZlmvCDBiaz1MkKSCKp7viBmlbimui6OsjyI+0r7AC
QssdbncjEBlttFD28A6AMfPAZcfNcGkK2W3mJfHW8qHsxA6zdxJM4aAWkma//dAt
PoiC6BmdwhW1oMVLPAtwKYoyqHuzVpx6fdSYaVOXMF/dFK1IN+9jsDGTzD0JB8ig
sqanz75YYLbHPL3TFjCp/Px8uDmTcjD6IL7kXvE816A9hiuYGb269yFIXxUPJjVL
GoXInvWC3KvaZIPUinxK4JqCBWYMQ/NGYq6fU9E3kIqVHWzD+GQ73uXc+sML7XRR
O7uuT18IlD1kAdGexE+iygOED1mJQGDH9wmJKqFGz89ldHJkHIFURUklzVK0l5zk
+3wmo5ZLqp2DZxwkDf5CF9DZh+YG53ybl61X76/DcgZ95UKKABfK4Z6SC2si/6Ck
dD9sAjQ1HgaaJGuwSrPROLoErRFQ/IVkFHD8+4fRRvEQaxKSBcmY6i1j0FH6nlVm
o75hs/WzhHCUmP1lpqTMcZHH5k17OzSfrhpki/FBDFZuEoVocPGr4nZCfllZV05+
MbhWnM8/65DwqtnPnvPJJH5E10gKgbuCmu6hid0+FhFjQFCEdx2lXk/JT1fj+m10
I7qAGMq3eu3LHps/hDBcOgPw1v9nbqGn4QLOE1vLpokDXLr4kY7kYUgxn4rr451+
ljBUB3q4dxQsWqmuIMq8lhj26ncVt2V4ob+Lc0CqCQaxdOXM6D+QCDIbCvcUJ+fL
QJEpz+7cvdmDZwFu0rF5HmLUIn4c9p0aIbKT8PGxdU1fvpOVCWFhN9gYY3Pfwfvo
Xf7Z9CqxLmqtj3pE/8vA4PDz+Md+K2AvXcjGWSOSOnBVtSFtUZZgMlqtjIyjEINh
+dXUjDeiqT3yzA1gI8OEyCLw4w2PrRSA96WIZOtg1/EUwD81bNiCd5EfCDgI8K+l
QYqjU7+hGvVb5wnZp73ku6WAiPvZlRyl6MwAh2FnDTU=
`protect END_PROTECTED
