`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I/WZK6UB6H/SqzqtC0UnQTu1atFIc2WKotzKweyhQZK0VQwiAbw5QDT0+6v4od/t
vGo8IkWRa0fCwuU42BrF6QJzEAa99su6erhxiPpg4+muFRr3eakngIfX1jfYUlp/
lkL+JQuK4UP8TT0BZK/5uWEPCJA0dMP+08BwH9N/mw2Y9X/2AYiXjeNQFW1E2T4s
t7k+B61GfA54Hx887HkQedgp5pyWDVeeremtCHbyZtbTMONb6bSLfPbtfSUd5qmP
oowhk9wdAmbEEka/J/iic9H5AdPGPlmg4xrItnqhkPjtzMmdbZp/ky1zX9t5H2n4
LNHUwa0juTAFrHFJPYhH51g2pLYh+H0nVEiT74E3WHIlZP11dMsrU+8OenuPYwqT
DaO8HWGSc73IaCSvpcRej7k5byZHdf2TlCS6qYZQR5+2QrCkm1YriTYc/DK8NnQz
Y5HkTjPJFp++Ldw2Ki8L8JvKZiIn37RegJcKSIUvHBLsf+pcDhpWB1aB01lTF4Xl
ukTiwPqAr49DASRI9O4lq6duJsYgl4aWLWabm2qw2oc=
`protect END_PROTECTED
