`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SCyiIQnxtsF0rbZtlxBX0MlKa/hpk0HpUekTc36IA0l+xaTOkBV8g9eFfZQe5niZ
e5LvOODbsOcwDf7mtQC8Kjq4l9Pz4pCS3CT6a+cghhVVWmCB4Jv06Bo3jJz+46vQ
9GYqvNahWHPhfQr75C4W0gLBYWfFDyEQxuxVBi0tdc+VGptGlFY34UFNoZyBK06i
x4NEmwzxgJl1hztTqaW6TGGQkQU8pLQzIW+gCNRMBcTiZI2q4dAj83rY/VTaUGzx
IdLmfDthXhgUhl0AlknKty2k/bAS/KuaeiNyUSOGbuM70Chl8War4JDLYr6B6p/H
+nCd72Ocl7endyAsXBywl9dVwgxKDIzWyqb0xpZ0kK5ROVO9TfTCf8acjraXathY
rIuREOrzJUPRx1LZPlhAS4WY2rjZjtw6WK72q7T1sO0=
`protect END_PROTECTED
