`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a3qHwfeQ01zuZt4Mk5W5BPIcL3BYO3BPn6mnAOoxPB6E2GakEt3/qzHS4jnTWyA8
JtW2V4KSHUQ0uErhnOpNAdCA4KMo4IVRxOAuvpUr4cCLHuEAs83rPSJKSQ+sB9wk
UVw7ZWwGXWs4ujEmhJUeEuqpo4ZHfj5CAlEv4gGABieINFWJFW2zUd5BOO+6ZPih
9iva3+P/jHfRccaPG4OZBbrhEA4aDxelke0Qv163wmC6UzpdeGbNirinUcUeW7mG
BJUFYytHdU32hApwm8j+jhxqZt83IqgaTY1xdcID3Jngqhhu3yiYr6uR6U22xLmW
AwS2kbNW8IYinB2etkxOQE8S36fZHhBF+eqyvQEyBfz7wEDZ0t7EQFHnmVFyV6I4
vHosd9snldT+Y5zLJFRE3OHp0DGSEeArsw3NDUJkdTH33VjgeXtbJvEl8CUh5y/u
fQm5pyhpe8T5vmZGBY9x4/R4knd3qT1hEPEoXWTyFDHscP6D/2RySBsDfe5zIEwj
SU5dWMYoXqK53TSW4S4YN0+H28hCIgHvKgq4pei8AXTFzvQHtis8HKr86RRmGBkb
WNJIcm0qX4CJWJg9eUn7Bw==
`protect END_PROTECTED
