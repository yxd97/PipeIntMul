`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JGQKdrZ4JTufZdSJXviCikBCJWk0lnRtj8S7YgZTZ0JYkQDvaBU5BcNooK8W1/Y2
U+4Kh2nkDU8T8VfN6uJaNe59whNPLUIrowuiWfgz+k805V8wYVYO0+qKPs91tfGC
HT0xY3LSIQY6zZDfArf+9bepAENEgvCfkALIHGVhqyG10Fe94IUImADGlzKiwIAZ
ndJGHGcizcgZgOzG/DnOMFDsq6du2cTpT6oGcLjZgxuDux415Hq3C7DFSTwoLE5D
VrOgK6ezh8zhMDq3Jj4/udaW3eMzPfd9JENXAxEMHuBNFhM+YPrhRZkJiP5JbY6V
n6mSTB7PJAt0fHbDs4x9Dg/YRdCat5NbsuDML7ZbzEiJT9Lvjj5hi3mM0KJZ0Xu2
C14WnRL/PTapenBapoDl+t6OGS8Txp584ODf5RjtfJaS3x4GE76WPD+m07c5mJtz
Jc2nQ9Z8+tr6ld5IN1dLhi5VutQw3YSIxlXf3ucDkQi74TG1TeIjGSMIbx8ntSY2
`protect END_PROTECTED
