`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nM5jLMOkbdRGi0epiacgi2B8MB4PTIW/lrb/ORMo5nkSxFiIhV7oljO9lY0E2+RW
SgUsCAcsMmvP/l+TeOpQZx7svHlMTebjFnFCJgtZRUr9atvEnNIQpjLzg4w2GYGr
hNMGVgUbYahBRYJBETSdgiCScFkkOOaDrOmJxoLuKyYiE9hzRGgv0Zv81Rk1bPQp
dcVHL3+BmRg1ZnCJ1zvqcxg6+dZkwkIanY2/RS1uwBx81rspI3LjdTHhVDOqNcSe
gxAsKo9HXuG3pIuUzxxA0AL6ehMZcpaRyZwJCUY7DaYOqPS0Z6+zXXYQuq2Pu2vL
AsZqvUp6KXD7+qqENER9XnUM/3fXoJNZJQWe5BPTXQQctoaZ059pTqVgqLWgrVMi
jdnuilhH/LaKLB5pjPHI7Q==
`protect END_PROTECTED
