`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kzqAtzB+80OYuy+OKKgkyMkxs4RmXD0/5bTTK4loiCbFdjtPLFDJiLdkgHZt3vMn
unl5SCeZWL5axbUjm53jtK0HnBrhZuEgxFEtQ+xo1L43WbNEMDobJ8ahcf+3UN3Y
tUl8QYXKT8UCXxTUY0udV7S4pG05B8K/gbY/qCsbWUn9tJg6meNAStn42MSx7kPV
brALQqRJNYMrZXVtQg3UYrjTVavgMi0Zm2MvgZGETWUXssOL+ODPa8PxuPRkq0xb
e1PLx/QpKr6ckHrVgHcH0pnlmolG0Bi8LhOr30f1HiYYzqsfsvI1JIZRR5zbHjAC
IGNDSgEbXQ+U5WR1RLIlfURDb4CPlzHx6QLS78w52QE=
`protect END_PROTECTED
