`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aUrOePUOyKM37I/gT/ahJ0DaWA7cB6GZ91A/Yt9V7FLiEnzyDAfWt3NDDqJvU6VE
GnyJ6DnTJYaW8LFv0F2/843gU9CrEYsKzWupQRIaz8BZuaJ9SlncuL2bm+pzlcRD
GEOAoHPclP3Ut9g0PsXSdenQqeggjkPpg5+W8jNy19Iu5w6j2iSE5ZbY7kjg5iUH
dmc3wsCG3ygA5Jb2b9tfDAmeYsuNj5L2hzk1fGXWLTW5Ee8ylb9FzHGRU6kMSpdt
Otpi7+U2CyQYB4qtvnexJ0BeWrjJuxO8PgQDoMxCdrM=
`protect END_PROTECTED
