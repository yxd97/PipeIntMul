`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p8HQCPMNadMRWQozuR7kBl2mq8oDMIiVdAlEEL3barY85JhaOZWZ2TpksCsrGYuM
qG1sD29TQubj3HbXRoAIKrVirrlggRvLTOOBqsOUqWgZE9lAkqVXnlhAyZNSIIyf
rcAGOKax15Irvt1hV8GWMaK6CNMAnFsP4CfLi73AT84QSn7sbsG7CYMDannGGrtp
mxz1nGpemPlLpeIBcka7oplmKoidHmv8ZTrRb8r9WdyLcmwiCuKXRFEt0J9mF6za
G9gSLX/D3hiy9lChB/1izm9+Eq8ppx02Fn5iAAEnpAOB+zvLhGuBb0Ncqt6/7nDz
9Ol79UoMZxumNDUf5QPiLQxONoVK9/9jIKuP5CoPtSvBgLhlxV7+fVG7Of/5gw4g
`protect END_PROTECTED
