`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbzWDUjdiRZtTbJ3CsyGNXI4yIIIofR6+8xqlNLr7R3L020dd1f6biE6TrMsjjN7
rHb/Wwd873KjnelX4jIFud6J6g+6RtOEXFRLpNXmft1mnq5MnhfmwMTfC4VT/3jB
tV1ztyBYt0/sKbYoRf/Zb4PlGGRt4QeWBi//fo+LyxZCuWUdObQwpi4mLcktdcZt
/8N/e+dsqfudRBLDpH/35s6pIOY6RMF8XwpRfYKj8UBIX5qHYcVR9wgrFMV4d5zm
nYPFZienARL5qDwBdsxXkHM0DD26FnLBLpNDQn/5fUwqExmfEXDgUJqsz2wZPPwl
D0xM2gXK4r7hDHo9GHtECndfUkUSyVhs4sNXSRVS7atjfMCRsYZ1CZtz9J99gKYD
EaaHL54PSZhcE7oRKo29Qh3e9+F7oe3CMT7yzIOxNdUzwarj7v4yydUGHAHh1MmQ
Fx1dWLMSRyM18CBK34iTlTxtc33FaAMlnmOmBP9xTzamYLW5I8y1M7u/4JJuJlRB
OrqQeuwqPnfIjIWtAn/ryyOlnqFXmnnA0T22hnYiML9FnCrBI4fj5X/fOJumLpn4
ENgGW54H1bPRO+mg60xmBnX0kb4qXW0RMF+9ROhFMkd9He7ooQvGdQyb4XTtPXwB
8FfY9QBMDTzlPvK40XLP2EPbQdBuPko/QLWzv27Nl0o=
`protect END_PROTECTED
