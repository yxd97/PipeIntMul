`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D1csdZh1PwLtCtB/IvgIT0NfdzCX/J3atWplxyCsyYIEAx+N0GLeLZx730N3RYY3
GmXgdwSIsD0kw/wi6Neyr/mP0Ks2pX8wx9T2KR8vfPEA81WCGPE4J0IsWKbRACtG
QsE+/M1iOwPWjqKRq2BLrt+Zi91KJPTsaV1kWefyoDlgDrEr6Y7U5tYdDKsPA+SK
yuug0wFUEAiue3xOjfHU8S0AS9veXG+oddiKIbyOXddfCFq/MEV2L4s3tpmEAcki
PK77TsncqfTTowS+pfxKONbLyJHZw8a1dj/VYc/foZDRdlxT4sr6KXhh7pGg1MHJ
3a0wzUe3Ow/4UTdjiktCaExD1ytMB7HOGP12bhsbhruTAZtZzggEDPo8ha1snpGY
1R03cfqzwcWU+TbpR5ULkK7yN9KYse42tQXECD9LHeC5BAbnQQFdzScTq5m7t9+I
k5mHDxRi6ed0E/6LG1EyTRLSsulGuKQyVPO7OmeUj5xE4m9is39bWPFrPDdIHpR4
X2eiyTNdB0jzKP6RVNCrDlyX9mgzK5R+wVnzdayA+/wcFUjWPslOE9pkuwCTr3Am
kRXlp74PeVLv+UD+zVA4dXK1xZEFAXVxhguIfunWZIl5ULpZ4I25ohwY+ryTU02H
KLn0lhAtc1Qmfk/7IG3meEfpKysA1pJKbN5P/Lnd+uimxKjz/wsxot7SpeRFOWKl
+lnefwm89NuXWh/JAuXgQ4qlX/kzcM0PNNAHlNuheJQenrewAhdUW/zGFUaxj2d0
XXGN4Etbj4ojRxhj+Y7yM+SoyFqpG1atq4EX1o/qsXx66KX3FNQf0GX8sCJeR8TL
+vH8wUvD/q+aw6dY9NFJjS+Ra8gfv4GizXZJRfkp+LYJz9oME8yeJVetMiKn/No8
bMLA3z1TwFNCGc7x4mEHsx1+1BlKPbtUvH0ETP/F22Eo4aX+sjQUkWrI6IsDcyx3
g2uXVJeQO6o49dTbuaK3mE+PkpLoOT1FnoSPbzqnr1o+LDAb4wnfEZVTYLl8Mnb5
HB1DW4wC5GuIv0nGbhbl/J5q2hJKpHfA+4+r0WlgaxADxczavxtbRqOcioi5P2B/
hX/Jjk2J0VN9QfMpXKc2Y6XA/DCTDv0Q93wkaoMWLy5kMnLRoeoB82jZABwPYp3a
IkTCEzI9qWub1VX4wP8KV07ROgDXC/2fwjtOSLREWockO1tD5erbTXvQgWCoil6L
DSltvkeJFqweA5Cf+JFY6BK4VG9QZFyY6BFQJHB0JaQhQvGPpLXI15qChaXL1FMr
yfyVIff3wWlEsQMG7urJUNarR49eJEKfVKcI1jSALHQQIr7LLfzJEviP2Nb7I9E1
S3SA66HuS8Y7GBwPb3do1bAVJ7HpQ7MAdUGzbqbJgZrCZ/JAMYdIM0e/XxTFPN2h
/wV/shaT0XJNCxA0/M6XUrSjX9231hOKCq1O8rQk8nUtGWFbN906708AbZVqLREk
+0UjiZTbfKbUTR1V4wvh8N7XIfDhdHUEL3UjrUIPcj18gLt5kB+z5+hAyhiL1c2H
I/6mbc/PASynwiHY62ibjWbwEbibcpwo7qlpDjlRqrCXWK3LBdlu2kJPhwUdKau8
jd6ZfOO29PDnNu7HFH1bjl3J3hQTBvVBhrASWLS6Wc+OQNuvbQe8M9M3ZnN49Tme
hSW1rTxQEEPYCi9ZACnNQrvrL6WWQMX+RseWnnVdstu36LyXQnFBPLzmpBXebL1/
B6XkRWuLzeaR1lmz6sDJ50qA4zpV/KUmkYafh8hbOa5BJJahD8OcyZTzlPUtT7Zi
puHJbc0yIWXjvX9ZSF0ysvtT5IXJQKhjG3n89qU2yZ0yvJDP49TWNGAyuir+whp0
ZrVO1p9hbqCewNvY2SpuXXCEBAfSE4dbXYpmSFHC+pirSgoNw5q4RsmA+1rA+ysw
dHMnI9Cbr0yy4fXBEJpLC1hlwB0wvBHPhBNYN0+0ibZ0JwF+rdnd4Amxs48geMEc
B0JqhXaPH7PnR7eZY8/oG4xDqnaujBdMi5cjmlKrgHjt+kYbLVZWl8CVhZZmttsN
l7t9qnuFYDEfvXTF5Z3b8hr2NSxTBJLwF3x8ZGF3rKFDIi9C47wFEhWpycWpDDp6
yHfAwN796m7gNVN6RxnHF9eZbQIPYtEKnR120s0nuLink3sNUH1c4rWYVIK0ZAJT
eDuzhnZoVIrYXJW0/VsKAv1JXXbdGJibwjAGhB94yZN6SnSEMCRgh9UF26CNw1vh
HG0bq2Xfev1hTMNfJnmkOIRxf1sfxyCmre0sC/6qEjOcD+EBvTjy899ncfbLIT+b
OrxZ4sH9bH54NpfOINOhKfcDgSw5qB/eIFz03OChPwwT9HRIRiVcmtX/Bi6uW37n
7BlD/b2GYDAvTidKxVNkNGXzesIHCiij1bvU3IpfgQJZHvSUuSSASh4v0973Nv3R
i1KpDIH+LOCUG5r62+kkKQn0kgXVaxVEBDUUAKl5kHJGmGifIfrT4EAHp5DIEaQi
D1OYatBiNsYjjkWlcC3QrJsx3USWQtySqqKkk0MysCOPwo2o0QsZwM8TKOaegK2H
rw5G39nNSjQZARA+wBFdkSkZRm666QRwyee/DVDrjy2F98jJVE88mqZQqHtY9Dg0
OstZbxQt1RQre/oXOmpOSQZBYWCyUpIbNMEBHmDndsOWSTPe1J9bpenltOCS+LBc
CYdPu9HhpiEQKvG8jwbXQ+OC+KzeRbPQ8uk4BviKgkihKPMmosyu4tKFqt8GwxFu
KfKhfhcLu60guhj/yxsnx8eL+4aY1lyVhpkWihMKLq/1ukDQuSwx6kUU6LJTxfPb
Up4uE6o8lWsvvoecv8+5VJZ3OtBRJji/xPIW1fTHST8qRAg0dCfeuPKRz1UaQoE5
tvihDeaD8qCMjGdbho80iy4Id2PjSZLpIOrTbM33G1GOQIiTwgijcDO4L8XrGrey
q+E5/TRBUdO5mU6+RhfOpsEwJR0lU0Nq43DV3TPN5PyApMTinUmUpKyHd2cT+VK0
yGAaWlEcYLy8e4BwMZOceHuZs+zP2ix1haf8SLEsZU2SX8kldUTYG9EdF37kzit4
s/GaVKlxr2yU4bClyOaorLWiC0ZdWlFiId/pnsQyKuC6EqzeJkgtS5e9sWSkNb1l
LnHBJGBzSXWuS9/bcJWJzV413QXLxDNR47wxdKjZITGSgMPPdKbK7uIlygHevypX
/4e7RqUVY0I8hKy8lR4NS7LPVztoa/bKYwrtxUFU2rtDu3LU6/zKEUmZBz8d4dur
zKVEJuYhgTXGjZrWuiD/QSzoYAsu6AD4ixoZHhBSITcdJ0Jczm6WzCp6ZfNyTco2
+vBQPIyj2r/42iEX/HJOxBOzRfdGtshE5L2ivtBrjgDc9bsR+mVAgAQ9a214NVh0
xcpYkJbd85UmenqfWnOsHboMuihW3E1e0j2LnkI+BLegWJBFMBCqhlxniyV2Q7mE
/r2TElWbY67xqnDps5+L09K1NMxWYhfBVYDVnIQGyPuAmdu/1ZsVuSE3jgpNZ6Qz
Ppe4M90s2oWobAmdjcQS+m/MvGGXpxwTZvJtvCCuMbRivlJoANWGdZ18CJOZU70N
r5PEMQc98CtNuX5QBCo1ZANooPxfpsBec1SQ7nDTFijH5cE0lYuxUfq41L9o9mTk
mS5lVPMJGJj4TNIG25uEdOJ5a0QFtclOwyR6iDfx/rMQn50dQaejTlmPMBRHbNNs
m9PJzKPQNYkffj/uehz+Qi/bLGVIXUBE3HOKjm1BxRoVUenFkEu8MiCy5U/x1yB5
PKNDs11mqWsC+rjr1MkWUHDjOGsXiHP3qxLPPVCdOE8RN49UhkrLaPbTHIZduFXI
sXFWFM3TSZP/MBZpCeZv5C2pWG+Eq/y38flnU2v2lC64VItSnoyKe5MO0a6OFhEh
8DfYZ6sVV7tnBRylDvx94UVlqPsqRX/OcFypkmRBaCB2JkgjlZYD/jmcsaY8w/9R
wj+sw8yQJEjeYrkXsRDJ3YJ0uH7c2QZBj7XnaXBirvM2f3DvdNFQr1GyMCcDuQm/
iS2/1oJFGqK3tLYv12wk/qEwU5Ie3Wfj84qOP5u4yiCOllehVch3qdEHDU8eF04s
PQMOfcYiWAXdPB2qM/h4U+ESS6AzuT1k86YaL8mffHAGGjMFGBZmUEzfKRkQajQN
zn9mqNbxX2kUDA69ojPB3hD2zptD92ugWY7ZZzUmsgln0sz2Ik80qDtDiJJTVDlo
+aUZvt3LQ9E7jj+CCeUH4nFhG58JX9TCfgJEUdga04ksuAVvtcjfIT9NLpPjWMi+
In55zyYFPJ9+1B/QqAS42MIRYyMZLz8J4pSUnfA4lCouIxNfiQqROFOJvwgx2Kzh
ZZUFYRsqTxq8tjy3a1R+B95yHmPTfoir0aG1kSRKzdXd11het/ccnvsHeFBho+MF
sccbC+OYCsh//w+uicAnec2TlW/aDvuMsbhleeFIhYVSu2e09Lzne/9JwThasHL6
GC7C7FddACL0aHtylEnaNSu2rg0AWRI1sThkWT9LZwrwGBauo3EvLbVo8rfjp6HP
bDi/+aTxg5uJ5nvfvcQ6FnVzxdY91uQvU9dF8knIE6siIMvwd1MKp2rp1ImFJQ6s
RQ9oKG4QD5pU5j+xMtnMEsUjjP9tLJjBAXOjOzP+2ozOEFk1/6ywzMSypwpd36YJ
CGJce6Qt6Zx3WGqSMxny2i0bQfJVWiOnaCJm6gXnrri+cbIbtX8NWAD2hnG2xC5C
gGGZwbVDWSTYdI0eZ+YLLai/T4vgB3tGUUsyWd5sNO0i5Z5i6UH8Owufy1OhqAVe
kOdX+bfWNrfV+8L9LnAEMnKk2HGtQ2r5aLM/XZa6NdA8Y0ea7dOVB3az5OJMSNQA
MBzR0aqOYycchKcnInmKH1U4ptuqHITQQ2ObKfdfcYHvxrab8BSYT8/AVOYNqdhM
38YH3jqJ7R+RO5O6FbVAyUP4suVdGu9svJ0ClOQ9n6IPfcrxFCQW9+sOrEk8e6MT
gXOvtVI1MBUPm9hYx3cueoVAJvNHjKuvuXvEZUDuJTZpVbkdNL9a7gj6d0PF0JI5
Ral0ZpwxA8+iTzSCiPyMmx/awa36MwOUW4cDb/uvikW+Ytu/M1hKPLkDv/BecZEt
fEGRY8E+bWjQM+uReQ/hTeiY6STsP9Mxd9/zWCoGrMRRvy5T/dkjkcWkHtFqkwj1
gfxX029jXr1MOzXDM1Mbz1TezjQ1fr5EvZLA99eEmJ+h7pJpfDe4Hhn1Nt3KQawk
Z72uMcF+01EyZd9M+30AcIV+UvkMGlzXBNouzuNj6t85xNkeWL57vLt63dY5bh3l
FBea2h/lJDpHAoDqCryQjQpP68Y76ZMy9Gbfr4oBJDywqa3Vy6BuocNL8De7Zn/1
ph0qXdGWQ0X8FJWyQ+MCOD5cZrp80jmJyK8dIK8FMUnKD09oDyBWfa3boQXpv5g4
CSBDic6XWPx7cm91o+V+p6oQPYpDIQlHD7L3AAK+oDvOmWRIeg5yNOzmPhNpvGEp
utPrWcJ4nhY31cNHUuxEHJ4kvXByC1iw2ywsfmWRnEsjWfpZOiUGc1Ie8qwcFeym
SW858lEvvzlK1mE7uQRrYGuoEXn7PTd53vQtCnyEFOHJFRijAHiw8w9phy9LCm1E
59zEKenbmDtEApmUH88n6joCSaU4utpgjdmETI0WVd1WmI3NSyAwQM+fgdMmqLxj
ZGEZec7tuzdgfb5cp1DUGlyRr2LMEhvep1FM+v3O3hh3euvNylv7+MTALoKJfaTw
8Fc0by8x8RP7gkgzhPUu8s3SaXdzXH8kez4uxXbrCCIH+UrEtXnNO6XpwW05QDnU
sgUlDWEOs+kDWJcAk1MwV00buiFt698GBsHV3X56sjHAhCmrfOGT1IRbtbxAaqMS
xTBlVb+Ro2UH8mtyERSXn8O0PrmIw8ZMLl+0XU/NA+QW9YmQw6FZKZWBP1flX/Kf
fU6lHzMCoCgVmbalbD+kX2S9tBj3AO1NX+PozIjEhALL1DgHN7EX9x80Rwk9O3jw
RcQ0l3jd1jwxPxFxS4c7C67U/5uOBfbl5O+rgmiLoscztYXwh0Ec3uYqdWuhTdd7
ho+RBCqoaZfGRnWSeQW/BqRXitKjmKxbFh2tpWvHrdWwq+vHnImE5FKW6fbyvjcU
W7xOeb52TJA7LHc7LLyXu7bQ7DjG7oQKSEdQPMy9W8UxZplOx6O4uvIPXvQAXttw
zgo49oSn7FTeTT2dHYBM39UzNcr0hva1esLeN1Natb+AM2SaL5kfG96MYeVOpNph
x0vAFxEII72FDGKiranOCpkhoENgNxzdhJ/vf2kY3DoWCAg+/KzoxSdKFWWj80Vh
OzQwxUbusg51N80SOSrt6ohFWXg7j5lPer3hafwJ3EVJ4jMN+4XOucYCUN8+SCLO
5dZT3Jr/kQJazJm+51IcXZndQmRSMoDQVbR7mSDQuVRuL2AY91zDXdsd+51F5EbW
54GiIR27CeWamtFzMRGko4evVfblzIEBaVDDnATjN0K5yzdykKc5Qmo908VO/Gq9
qIrK2N4D4KEZ76TSSHKer7b7sdbOENGlMq1lenxnPhuc4UTzPn6N1fu3f/+z511P
drKRrp6c1Y4OIQaPdWFNuYaUncjsuGxh5Wp+Fe1QajLb7VpK4KOnDD6PfOexQEnI
2SzK+PHXa66sfOMZ4UoN0h4Ul1PXuI5NTHh2td1LXRERUR4gF8BM+3ctehS4aSgJ
eZD3AJE8HIsSwVQ9TWK78NT4ND/gXHWrP4bRy9bOBByOZwwlRGr7xizaFfryDmBd
ssmGBVO0/dDYKLfAFdT9Rm34mRSA5oF5FgbehNmXavT7JgxXk+EMBbWkBzMlrdma
FeRPISZnL7Yna6OMQtyRTnxJAp6VrxzqQnHaRIxEuLAWmRkaNbC+ByVUI1h65/gz
TDl9q95JdoTctDcrs6UU/uzmOmvWJNNVErHSs4Qst4liNSIt++zJTulfhNkJv6mU
09EyO6zduqJemHgdSTbzfjC0camajYeaM3tCm+xmqOGNNLNTShMCJuQ2vbQqWgAj
67jFr1sqUxh5ctbKpYe+wcQwCm/vx2slOk48XsMxWHeYwYhbxqvVzBvVwYb7uApP
BmF8AQBj5oJuebKN+xRw7alnMKxS2Ij7AoQRZ67UJ/iKAsAxac06qvvUWgliJHUa
7ZE2T+jOFqnkWYHM3uMKR8N2RyYJY6Wj8YCgLi31bV/wuzAX2k1tKHUEQ0+e1bKY
lQKBnTqmYywlZrLx/b8MQGWEq8NPH8QFSDZcgTITWRlq9fytFIauMxx/b0a+5P+5
EUB1F3bNApmfoaDpVlgfsJug5NFw7ya1xu8OxYyOTOaA/EoOJQCCUoSESr+meij3
y6/ZM1EZ1AcNfhL0sfhYHr2j+Aa7PVWONoL5wStNG44rxbDRgZ/a2cwj3gIu9Jod
uuWeVJWxUkIJ8xVWUKDIUEtentGU5N/29WRy2NuogXMh23cYKEE94h+AHrIlyNIA
MZa/wXaZcR8yQYL9FJB3V72mnAnAJ6E43ue7LlpyYy7jRDmM1LGf2yrAJ1qu9Pk+
zCQiAwCEmr+gubsG+uSKNmrjpHyrZHg4WU74oMBRSwAODnnS10dq1tth4IMf8WYz
7RP7tlJvEpcgxmHt8ODCNECY2YPXhDvjTO4te5kXsWq6a+V2SM5cOtF28XtSw75P
1k0aup813qfWePD49a18B9bcHhvsurFBuozoOLq6P7GwcTbWf/FLUuMOrhGHmC8e
KbA1htCduBc/vGWyWxi9I/DvbfKZ96+TOMflhrJWXbLltIHu9dms6oVp0/yWwaWc
Z/ErS63kzdL4LeBH4eQnKcDW1Waz9sDNeCpB4nV9WO1FCFBlc0t8bCKXQ4vV2iIo
V1TDYojIYVxMkM58A412dguxli0xjWLNHfSH56jYzZWq3KNUuZzS9Zp17kWRE94f
KYycpZIRXjlDmgjEce9dkYcpG/ChpZ89EBAaHPv2eOI/XturBfPJwCfeJ1L9iPjV
nOQ+q9uD4mdZhzFF05kZDl9zH3TjB1QeQ4K9M43rqGFHer43vt8kA1xaxBORMeJA
SFnrGboCZKvMv7gtouNM1yLrN+XPzaf6VJY8avB4NOpASb6WOyEJiMfg2EfvSA8a
yk/XO0SZFOJQBOeIPT4P7nO0u0vIM2L+FCLPS+VAGbnEfVGajPjUZ12QzwHRT9Px
i3x7oJJVOtcn5nB1EOhIrzBQNgw2mJVen5J2EFHggngW2c+QDq3zjmujQ/L+Vj/q
T+SdsaHnQjxJ3wO5Yxp76NNnI9az3IHG+0tKgspEOyQarohj5D5A8T3SlsUTH/0H
jV7a7J5skHs6zbYyxfEqdglVvcXEZUQTO3TCynwgZSE9k5Jq6v/CctjEcEda6hWx
vJ22KGAM5NDv4E1vyz4YmQbdz8sQHQZPH3qw7ZO1CfQK8R48UoLq0jAoqLoZ3ZGb
ibVGFtoIvMpojps808WP+IX+3XJjoO9RWJ4aGxDgUBQHQ+zaBT5grOafZdIi4Jwq
S2/1EhMh/oH4VAYvEJwqNkyenNF3x9psTehq76Hm4gSeIw27PnISwN2GxTQKSxjw
qESgNSr8ntf1JhsCYO0gJfuJ7xv/Gi1fWL/U/aPcDmQR2ztkQJJACR5Ay5sDuSZK
4J94lnqD/mVVeJEwqjA4WmdnozhSpOpIODgLhdVVRePWX2Xlzm6q/HS4ReysJNla
Oiv9gzDUku8M8t6BHBJ2lXNwR8vH4q/s8wMT/BgHpW4N8U0PBSiHKxCIv/dNHeIC
m5h0NzIKeDj1ccSgaM5RcC6vixqbwIWe3WRqG6ImnSsZISRzLi5XfI/5Hp9EwqVz
fyhMi9DzgOuDtL2X8xEXH4WCxH22hHpQnQ3g1jUnf0z9luFRXiE4uFPrMJl/CgxQ
lF730eEuOZ0k9Px+YgfjPzzc+rEeTtmkZrDVn7LrIH30Kg4Ic48Cq/g4XyEYbMPe
6WJWY+WVPQWcpJHnizihg6VOzsKIv2ba0O/iZeg2S/1lpK0HjIdVjubgByEo4FUD
9ucnz9InkJYMl+cI+kaQdNrDIeolI4XSp32xUS5mieOHZwG3hXLZla3JfIIkgDqx
fRjhQgYHbYj7xlfuM8Gce47KuGqbMES7JeyJNNlpXBIO2Wc63JNyyRVQ/syL26L9
sxyjYFbz82a+VytcC35r180YBpSPj/6eGiew1bHD79wHXUsgBHA3FiUkSpLfELDZ
qgQ/rioFtf5jP6NsGBu2ggp+Xf8VQm8eybMBf/t7CgEqOfci2UaxXAvl/c6yRnVj
CjRBYuXBb9+Pq4dBWiVQXTjtxtBa8oJsl8QKoJfbR2FQ+2cT+dIM6qs1phP6C33K
SvEtCn9APuUVjP0F4VZH80DQbF3B/tzMkWBbnFQ1wBJCSRQ3cjhnEXBuSsaDQYVZ
jR+ev1KfLBy0kcva5YU3LSfqEOgTEJ4jh2SbbwtwouRXQDmTfA8FtzOge+a17qM8
ALY5rhXS1J3YE4jm6ydHgK6sJ3Gv71qRAKJVzBcF47ISKZw/em2q7xTOCUyMDzrY
8pBV9SM8HAenr1j65ZGQufhTpMa7V/+bGe5u7LAW6GlU+T3VwT4RXh8mi4zOex0+
jTmu8XgA6+4nFVLwEMehgusgrjiJv7ko5q+3cuH4qGVarrf+Qy53xbSTre+kGDkP
SxRI5Wnho6wyc6gfO9Ws8LWVB+6K2OYozLgS4JjjFTt1lEnPxk35PPIEiiuGJptp
JKmmTyhud3PPZIz/+/pxR7MJ+15uSIdKtjI+/cX3oQVXlfR0Cp9nWG0uI4K3eiZ5
PRmTa6Rhe0w0pRiIhd5GSHvdNC/a2Z6LM2ZJJmfu+eeM4GQMmFxqK/JPxNTMmklA
45/4Q0YtPsSIBm2UVmKjiUyXYOV6wa8l6QMUzPhdrEbUb0MjOHE7QCmxNt7maPR/
roPjaOxRD0RYjbd+K7I+CvsYnHRcVuDcea4oPFDD8CPJSkoLfkfBwtgwbmdX8+vx
fkX/bLvR1iEw34YaF1MPlvOBK8eLWiBBd0hYOZ25B1DeyrgeKRg9lOSjEncciIro
NXPZs0BvxXcyEhHVG/Rw/OboH9Ri87IGv4yLqvNBlT7ElUxsVnz9bjqu6IN8vV6M
BfkG/XNBKTu/aRam0nhBElN2aVznBFdk0JC65TrJHQkwNt/y3RVl82km7OoUemb0
YsEbhxzh3lWYJr5b5QGST5vikIlXAIL65vGrlgSmzFy6v+CSjHe0JVG32G2/iG97
Hb76Qo+ThZYH04X1Qs5nLW/Y1KgbLjEh9hVxMzY6UTEodB99YhGvsnQl2pW7guMU
w4JR8jp40CzzVJC5oUQjENCoIE8p9e+zbt3d/xqRZypziry71OfLBdivEYPsQq57
l/YadvHDFfdqBZNpOrP3w/PPW5PBIKS/0LUjMDkzoFzGrR9lAfzUye//t+l+xIa3
2yWaHjt7nOqA/NgpIyi2ufczO7kdv5Pax4MjSY8AuzfU+TBkRi8306kkrFbry7P5
PswIGyQ7ptmH2pV4i9NCfCzHE0o5vuSfHxQwfcNE/1zezAZb1pe2YqHmZg7Nb8Dh
m7gfyk/EDR+MjCqjsylXtAewyXLzBA5VWvoWELs61sC06fugpsyBESF5ND4brTjs
Ikas2qecm1EN1KO5N/1U2Dy+GzM2FZxFCoeRzYoTKLDgFHJUi4qzUFUeNMsWiPMG
oZSqsS1OzYY+xeUeGEZr47ixUiqeuhDOD/SEtKFgyT7G/ZNjpR23YcGQcCRkzytd
42hhpzY6UcvGukoESkqy4G2Q6go75ZXWsbSUiOdkNTbT8dZBbOW2YZipqxrsfgIW
2mhUCkYlaK+EsZi6AZMD8SgnDN8vP6MqRIFH3vlkDZtIphtNzX1xmrZLqzIe2uw5
Bnbiat6C1eo03RqEB8UTY+CbjfKIr6XQhOCT4EHdN4f5MwcZLt8L/fEVcgqUbTx6
`protect END_PROTECTED
