`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCUAXjodC7v8lPolmgva+9eacsKE3BRy3IThZZOLl6P2QrhxHPrT6uN+5vOI9yzp
Bztnm+WoeqIC2T0YLTsKx7eYEbOAPpiOpY7dJx4jaIlyNCdjRHlFPmp//daQ+WBA
R1Bmmo7IbM8qMIte7YrDWpA840YEBFiRjRV4LvrcTNFQfnc4O40DyRW4cjt4wwwH
h2Ee3PmsYaCZkmnWRJArdeML54RLl7dNJjmeVN7i5u7RJ2PBHEej8QugYLlTgLvV
d7JvhA5qRE17QEIlteJ+2H7a9NPbvU/eZ40gyn34wauqJ7x8svSyLzZlERiAb+6f
y+cBwFc4jmocEBwlPlTER49hkv/hzhtMWBelL2ahESC1M/B9wZ/qlfvhECRYyixT
jmJIlzJcPllIKbfsbmUa/f7Hj5x0BR/nVK08DwElPIEwkHXGPYfpyWkqU/3mKbAE
qAR+PGCzcQGLOY+Fdv0RvV36REiIkQCUxEHGlhAYrCu5/AovbVTWsP99/RLe8Ule
l8Bd1++crerRarxudaif1ca59ngY2b1Pv9clxsHoUgxrtH8v9FVeIvBcJZy0jYTe
8SYDgz8193ZwUmccDF9AAoFtCqNhGccaVuccqnfUyQfPKIPku2zUASO5r29QRUFb
rcBYptgDzDxn+DV0nzS5JikdyYQkwuPWmh/jrfinXoeQ7BalBSwhVZG+WcAFQSfb
Gvtj1z/4it/o92EFwDR9ZMw5SKuiUeefxlQfW2MLqog1SKtHFmyNLUg5KHfTpf9N
rneeHniITxigECGQ4SOwtTuiGBOQerVTSaZf5w4gBowQ2f8icXUVhFdHuifjw6l1
v3s/1lMLG+j4itutSe75IFmLsY9DDicHe/raeKGOSIo48SeffYez24MlMvx1aSul
qpGYOgd2ipvr9vP58XDwTF+rgIm7j7DTZxwfJZ/ZasI93PeLRODmr+44IVpGBUu4
Q1YOPrk+2jDZ5GbdAuqodvvP0w7ZhsXO1MEVhvTJi859uZy468qZKAqu6foDZZGb
OJt18vVgQMApsWwCmFoq5hMkk6KP4yYLhX3ywsL3XMIsCWX0DiRwYI3a5YC+khFa
+TBx4m2TuPgk4pohKy/5gww2lKrPwWkdLYOUtY4+dyTjZxdtqtr//DiNJ0P5m081
8esdS6udnx3hSzXa21kj5j0p/jkz3fAOVoZXaCX8laN4ejl3CkJ+ULxM+bdCQacD
Wib4UKKNe7pAO72rIHsnO817WFhgxhZ/AfoLumI+xUWT99pdh1ogkd4H5tewOYof
w+3S9PY3bKBnNHZZesF33O2xijtHbL5uuZ19u02K2WxgU9iTlPSzWCG9JuhsFpLw
kadpLQErZui+RUH00ucPQ5OB0gWMfiBlnQyuoraC+jwfVp17HzRay9J+zRqfWFOT
qqOw1HU2MMXHHoQRloDMysMPonL/qwu9d+EfplWJIkuEXftMsjNIFDlJuVVXZPP6
bxgc+YTT0LOfMFO0aBovpO5Dim2RAS/E5Js0/hcBgWlhAFH0HLXz+EDE8gOsqXAh
WJZ0GQdFcRA4nUK3LjpnptWfZWdGdXY3+ogjNSYWvih/vfPuDJIk1gGMRp/CYeG0
qxVyJdS5jNfe+T/wm0g9qYcDpWrKEZfE5ubS+pvWt6mftbcMfllyn/Bv539oZNW7
eG+JJQGZaWx+QJXGQOaCwqjSy8kZh2e4l4wnZ8NF9FU4IOS3t2BuTxn82Ofj7XnW
IjX6kuujRSMsOL5DA2qdw3MF35+JThl2yL7FDoqyCoW6jBGutSHyURrkBSNvyOiV
lV99qwDAJJHvXKQTuscICngTzachWIN5f575QYWVVxbmbvYXZE5LlgYcQkSY6WVz
0nzYayBee5Cj37q7JOhNlaF3ic6PqSZKfSgpXhJrVlEBg3T8HKiH88GS8wqLBJgF
CvrSsFez61yPJiJI9IDbVH74+GeoZHt9aH1N03lUIAFJlK6KCgUNCwke1Du86tvT
rbbYB3HIF2yPfolDqdrh613hn7rPEAZhn1JviYEQqQnnuqpC802FDQyc35VP+2SA
Bmsb+2tsqGilLe3n1QjSUqHkOrHp8orX912REwd0untxMlHvTf6TKQtQSIbJqd9G
h8GyJ97hu03r1qTLCcQoAl0E1t8a91qXsygXYfHrFqjk4WGGjD5Yod1GTIYiqhZp
GAZkq8FB0cjh0MgKPoNLxJnoYEMrzgO1/x/wQiXlZLi35ExMf6Q0hPy8xvfEE4w0
9EgCHeT46r0CHzC/S7W6hglyqKAgGmsNxb9UMlxjF6IBBbegxc+PmhOT+G9oLs0q
KT6owpSsKg/qfE+JWYcrOcWBCl+iyFu6QL0sLtyOJ+Gb8+y2KFc7Bn4h1EMuf3S/
1WevlaVehvQ8WulWugrRK7UNNL5wjJ/qdIacCJps3DFY7oTs08CY9XT2U+9nVeic
J2G4PmSU1vv9h5oMPEvFollY9skjlqiEXE0Uzxb1I4pmq7UPgROx0OnuTRpvICc4
n+R2RcKqgAxuKyl1tFHuMvykRb8m4dO2vHqLnd0z8xIo5EqeNS1WYktOJz7w6+Fw
TXOpWKNHCMmi9USShayzOqXeo1Sg8aiULtVD1givHwSmn5NZFYz3axcwVjcdkGKS
NUYXBoq8JL2OWWg+WMi6+bKC6SPuolzGtDMzKTUV5/bAKf6AxKeIQqB34n38XfG2
DAuttZqjrAQS2urMb/cJEeaBU74P3u7SJ3JJCgYTkK+kk2QGc+bcNTPUYPfKfDYF
Xi+dOuUngCkiVb40CTIaWzDE+PeGmMmhR3TzwTeQxnSfzUdq5m0Jh6uf7dpVXRD3
2/7AmPbvCaif8GmTlTljgDwxYwSE1B2GzTLs+mSVmwJduH3N3Q2JYDBoBSg1nayJ
Vv8e0W5bW1Uedhbbfux3N0BhlL2umBUIGNesxilyScv+ynynRqUBFmX9nljbnaxX
48Q6cNfdNn0GpZwDvW+yJM8kLnv/CG7kqGuD/NAA1JcDxv1enJQG/F1rK4hcAufk
Xv103ad22Xw3xR5d0E3Kx0foB1EGnvktLmwu0tUUr6HYfX7IOsz9QRLz7wLzY2Cs
O6Pw7U8dIwFLw090EdicRs7x7u/Zj7QFEbhuL3qyrB+/Lre24KA6bGJ6XrJFnZAj
8YFBpEoB0MZEyaMrEfG54D1n0UDpGHXKTymB6/N47DAMK3j3HNDnivZ3kVY6Qgdz
mKsnz/Kpor25fajf5Ou8Q/WmKmsgf7R7yosWgCM8lNCnauGAFZPZGz9y3re1+yKT
Wl0gPQ1zUrDwaJR14HrQNRwcWnKp1SNIGLYqSBx2mGKlK3YfXkFLE2mjQ3WjE94M
TuxUESS0UVCmhbVmAzBF7Dzwt9I5jWHhCRp3+g71yyQGMv5kTEx8fcAJopK8YgVh
hcW/wvoILY8wVz+bokqCBEjqxFiQnMBN7nHpBLu5jX0YeMR8AyBdWGswCFno9riz
yNIXWBeWUuYWpiBHQG5cgOrdcIEibH42TSDwLLeraaUJgLBBniGSt2fajuqQ2udS
ufA8E6NAaQEF+1hosmzEPFHvKikMznLI7DfBEV0eQtYdvm8QHK098LRNbPSvwt2Y
lBUsvAp64WuswHT7ywVJCUavFj34NXMOnYmdVLwbxGD5MRQWKltcz5YYr8Uvbzxo
XH3RoyKus1Itetswk6NAkYo94GONQ3AaKK9YHEuuFUVH3tg1+iPKmapEo4QGTAqA
g4h8SCCzD+xXebFGOGl/DyoCZVviopg9KgLXDeWWJnl6e+uOi7yIdv8ceClayxOb
TohhqkXVzgWb6xhLDlJdm1c8Wjk/JHhTqdndrq/JmYGBhnVJPp1WD0q4U+6/gF3L
vPHYxeDLBXuBizOEuGlfzFfvJEPcuFY3fMwLVvhdlmrE5Vd1KkuCTY0WTh73tUiu
uvgh+/+bz4NJHFFCIg6kDcqdSNwmmrZ+ziOBRokmHlFcrFwrSjxtIQtJmbMutpl8
LU23k4exF2Dzwvmn1b0sF36AUVJAV0T40RUs+FMU1spJQDZuP0WrwhGop0RT0KIT
CqOfUJW4Cz15PQj08lv2cGmJs76wuKQBXUerhGatrw5g4oqYHld6H7VycDHgb/7H
cVOoze4r77AGlU1X59AbpvUixW4ykHxvztQpMBJ4SYKD/KnagrmyYmw5K+nnluop
gmENyQpEOpUjMohbRXJtvEwr9l01lqZPwihU4dZkj2OQDKssVW1r919TFL4pHC30
u+MZnuMHQLQjQt4iCOSSnCEtgcgsrMlFPI2S2i/mF7KyTGVH8x9y4FiI75fb1U/Z
X0cb/NPZvh2BfNliq/XTrFDvfQEmtxz7AqVF5lWOP3l0cNlmzAv+lTNw4+SRV7xU
RIWMZ5RVAqcLEh0Te1WmsL0CmKK6G55XMfg/0oVhtIkLymJbcF5kuIkm33XWmuLQ
oVPE4V3uI94cNY/wBzv9MkKPEQ60wqjISNlqssUu26TngFTWDfagIdYOLYqm9yDU
TLAvvRZ54dAPaZaZ6Un3Ea9K33/BmBBIT4ton68IEpLdqahQGgUoT5xI1EyZ/x5j
/cWwc5sKKEYs5LGHJAtnwPoGFM7sotFYrT0K0Pifazzvgc5EfZneDAG0iRGPo/79
xLd5XaS9egZu/ttFlckCLYhYQHL9X4aqedU9K8krTI+NVOk+dcu+6VtDgcN9T6bs
sjtAnX/7B0M7L3EZ8SH2ofhUEQS97jvHwRvAEkbk/dRIY9q7cXoXkfCeaJUqziE2
+NeLiQ/kUztejiL7S5TgRu1DOOIrCwKz6aNTIsMlPsAmWaXW2l464s98pE0g7N7u
P1UIdCvikO/qYaNYxM2NXtCGmOa6KUeZ8PPN37L6jCPJqE2MHXjB/73L6tifAly9
DWG0/ZSD9CqO8N7aHvELsk73KZuC6YGULFWcX70826yYaFSmIjtTaw06vjNnIaOf
`protect END_PROTECTED
