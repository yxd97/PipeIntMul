`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GkjN3jPRXLYdAIAuh5DegdZtKsXDObB7ih0VdYsHAh7WVCOnBWuDi9PLapOZUQiJ
xNwH2qLUc65269tol8SKWKKeZezUkjlOLlcRhOtUguCyvKABrWuHX0i79gBWo0Jg
xm59ELUsaILy/oKHgTl0TozT3X+Arj9Te6TjXxE+/MO0RAJ8+IyFCgWhaT0hVHy/
IcHHb976fzxCl60eQvW9M9660fCMi9X3a9W9Aa1dYigQJHwJjMH9Cwp60H0H8iXJ
6PYR31w4qHfTCyLiRkL19cjb9qegDyPcq7i+9ZV/bv1bLpsLdsY31dGmlbXf6A2S
hdvcGqauNXIZP8veQwFudyj7ru9Plqe7Yl5SA64RrOoPdneUNsCe1M8bwL/gckxx
TcOphn+Cj6Os6BM9IJcBVQ==
`protect END_PROTECTED
