`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCG9cmJLJxZO1ID1MV+BQYOxqSGd3/7Z68xMOSfveaKPMZRyrit0E1MhwuvmOo6l
b21mbjxWtgex69LwK97sYCGJlFslPT6fG1mz/uOCZt8p0dy/31mK57XjoR3Ynru1
bmEll4HKOUHkAJXQJ2y5V8bF6H0JwtayEnbiovM3jhMEDYECbFg4cCfUdUHVClrV
chHaROBwWLoSL6pDuqNvHPB5dOn40hckFEHNSntc5MGHAXplXdkYSjXsuhDs18vE
497St+Y6RNm6/aR1l1TTWsFB+A6HyPxpwx/vlCAVQx1qqZq8VT9Vt4dV16M5nI5i
UJgzEii0n1g38JuRPz4UzNlKS2lJ5FJrddFCVQVx1FfA3yQWKOTWaBLqbD1sdnGG
07H8pvR3M543vyL8nscp4fVbZR6teuZLICOFoQ2IQP2N5k7iMpGLdNNuOy9MNUr0
`protect END_PROTECTED
