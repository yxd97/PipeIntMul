`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/uU75yFV5rqwUXylIwr0G7BFl06wOP3uSJrnnBSMGoXVI6742k5R1YTRZIlzgoC1
CVSe9hmRuwa+TQTdVDjDaEiEhiENmV7a6GnYv+NFe/OgM1ZtK3AaDhP+u/SqdeWe
gntzvxGL+hC9HOqwAj3QlSw44H7cW71MgtH8qq3n9HaFVTxbeHWa1kp5QThkgeWO
gXBVvbMo2OaElwFpgyjt5xYI2tIzEYqpzpGAvgQKQP9lkzPK9FohEg+51Yorlqge
q0eMMUX+Yvahl5UKMX+eHKDM0Xa4AO4eH2JWSkCIVz16lh+KUCf9yh8jeGjDvfCV
oBnNpJ3vnOoojNlR+w3rlgg1nG1sHYl9KLkhxBLVhmtS0PAOksRDrXmeQ80eABYK
FdOobqjXj/tM1JdXaCrrje7iXioBJ/OvUEvxBrzCJ9QZy0+RdCdun4DwBwbYNnbz
P+IhqjC48kej8FIepkN8hvaCo6eH6WJUCPDikVeL/erMjLA11U7QTbAC1cPrXcit
PmEBgiz5Dq6nEKDWpTFGA8EAW+Xl4yClSKX/HGrYfyo=
`protect END_PROTECTED
