`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SiuijauESDVebfiIviqjI19gsGcnXjUFtzdJZHoA7BeQZkurow0gGsuRGbxH5ndD
GM+QA5s3YHU7ztRrRNwxBI/Kk/4zfHHqkqwJLSBMLZIH2Q4o13fikSXk0bhBG4v1
r+D3AE8DTxd/jyqns3QD9F4cMc3CT2NSCsUalA+RhQJqFqdSt1crZ7cTsFFW9FNB
QZQLXvmgjcZfITjLaoaYPZa1/Py/tIKRmQFPmbh0h79MgWJDEyAhA8m5RqUOFe8G
KT8ndT3T7DyqxXsG4IZxsql06xke88JnNtXxsqxXuwi97cIA3E+MmfiGwbzuWkv/
MNH+FPro5ItRbZgxuCwgXmPI3qqXl+MvtA6tljlds7trOIdMczzE5Snxdn/GHKG/
f5Jnk41rIo9dtoTCmtSsJ+ZogTUViym6W1ANnNl1N86sPOqpjQucATJ4eEroJV/K
STN59dC6jB0JXLove4fRhQviH0D/PXMnJrjLjqnZXAV/q1B5CRj63XQQHFbiAyRJ
BJ41IgcqnaeyhbsDEsXgfte8+m5ul9c8cLdVSeMUyoUR5o292b+RDxddA+4oaJbD
ZyISdhe/FL3ZEl6ADe021jQ8gkdPHyq2bhq/GwUfgjc3Ki0o3EvEjSZLkCIjqm4L
wQONgMfWEOuHWprAij00Omf0/j09akn986OasUnwfFTytdaGc1H8ZaNvxAGb3p5e
hmLIW7juZktPfLoPWydw+Hzb7sVZPcFuov8gRdxzRZTQYFgfRp41LrEJJbect0u5
qJZihYM11AAH+GspOi2b3vC+YiQF68SXN67ILdsfoUrmWgbyzj8Y+wubazmkOhkB
rWbQVhTp/loNMi2uu8j8amZQT2RI6xuOG+tNptqDokucFaxrCxPDKEj9GPZoeOU7
+KwF31P2YlYhAI+LvOVRd5XtVDAoinWE5H2XG3OUT2TyeZ7Z2MtLWaNtrI8XLpnP
kNongUwnOcxmrNY2p1/sMQWt7vF4/nIe1g6OjUuFSgEAUuo9RqOsAj78VGuSCv9K
TCwxygi6izuI83KUFYPM39/GxhEyQxzSXoyyS7xcJhTjEPZ4Jy/zihx8/92wk+8N
UKToMB6Qhb32kqJJPppOWZ1zKXMCXj1nZLMCFmN+Z5zkgi0rv+K5G8YQ0zLyUvUf
f4l8WdWNZVWOsJOqFLTL+H7lftXJ8AT33TyDyG8sCB7RgCb3ZyXfG0orSxoatxDb
T9E91xamP92jdRFYZUCQZsp9QoEpiwww+xi749GKXC3aWqzDEK3jfMMLZjhtyGro
Z6LSt3UB2LWd8MpPwAFPHYWlPeiDqiOETWBck2K2Hj2kplLjjIJRjBFQgOWE6o5P
a7BeoTKaNXzyFkUNJlfPxvzg2werj/swQvqKfOycyPLmD+5u2rUGlcrLz0d8YAqf
ncUUp+3Sx/vHdargZTbVy3dYLiaACzrmjFuT8aMQA9vKiGx1N5O361GSCtC6WooW
9FSkByZcCzY48BaC919B/RvCrCmmByKOAALtOHg3ULIsGAlJq6Ww8ZFB9SO1c7+j
uNk+O6jA7yFrMoWlFbfVt1NhHnulSddbL5QkJvBWi2J4b3jsdWqk3TYqHsc/m/vN
qT8V12yjzET355AfrQydAp05oSY9CnuwydXrE6klJMg9YGQmlmSL77sPyd/Jepvj
QFcGK1Dxb3fg6PTF8Kb33FoD4pHHo4/4RbrEo9UvC7M97AytHLN6L8uHmYxB9yLI
50dYgoaMtMfU6+1uoy+AH8KADFeYe3TQQcMgheiZP7LMbTJPqcG20iVWEetvwAFq
Q1Tl0eCV41RUgK/aRNlAoFxCrJTEhONGu2KXgMcDij5bFJ9sW6fNBpjW5rFcIUze
fENU6++yIh17LB/f0GP3htyNAYuANK79B7AQDL7xbKcE1YsiMeS5mu8CeD2zagqu
MOBi/HPbIdv7RN5I0If/+qNg5uyQz84Z/RVa2OqWVgTn1zoHgVZ7hlDKaLYXZRx9
ovJV+yUZHLn2K5R9p89KfK8/6wocmtiw/4MA2U/MW1uhQoeUjZeTbiC4xWYFjYA+
dW61cNZe42ggRY679PYT50PhmiVlVTBEyyNG82zAwBRJCr5TVI8fvaiwBIHwf5Fl
PBYfvKx53P6LRLlTMBRcwlLtgMiglsJUZZEDpabSaRWE7uyA9rRWx9bZnjurPMuz
KOxlqqwI9kg4HlspQ+jo+sLgl+QEtiN+H8jWzx8ddokfVAe2+dsofFvXuwXdb4yp
vbVzTr0anFMICkcvMB23aMGvaS5dGELjiHCxiqhkINwmawYv4ANQJqnKvOy7+sJ/
nhuBYKcpdERzv0Oc6uJ0H7COj8Ewvt30VrjGc+F2STqDSN7RTxfWiblb/DjrZLxA
+z8Qd9E25Kryf0l3dYfCxc5KRqb50KAGdLOUh6FHBY/MaYzlovZtCQZymsbJvsoA
EWz3xjHU3V6qiEo+Q4MiZMvFdjG/p7uEWn5/fuP4avpJCmqYbhLreWpsxHmzdYdx
aq60uAe5CRHPF1O3sSB1Fk3du8yEW0p+JtwOvQCJ1oXDGqi4IUJMu+mYSMLgD4wl
+OVVqDf0dBSdz8TuCv47mjp/LhIsHkjW6bosOyrNMc6lOMhPgQAz8X+H3EohlDsK
A+mS4oBMFF81f58cStDJluc7ba5cFPtxNeBmTT9OYjcl0+bBwOf6LbAoqiLXoP8g
Oe0udzfz8lnMfrc7bsDofNzAwUbA+7Ig+yzVtTD5hAMYpX4cXqWYhrvxM+3YY/r+
hAmr2lXcAm6yygDg3GcW1OBp9RdcvZFOgfyuunDD787BvYqJT9osFwGQaZonVipa
J7Mw+1u0ZGtm6y+yDfWd84BoRA4538xPI1pbHrfSQvy7T+2//u7utnFrJeCniWdD
nDdK3Zcpp006G4xARKO7qLtatZG2pseu/9aUhzMjABET9DiQX/zpAhwaWxQb35dY
3B7OsDvMXyUsil+Hi/kyBo6AcBG6gKO4V4FEOcVwixMzsMrm0kzjgs7by8nLyh3C
EdaorUeHHUzzgfCTLrdnjaDBjAfuRzOgs7825WoWOoJN5+9jvftEwqxJ1X79YWCw
GIV8dHJ8Oz9+DVr7G+zsPzL2J/L/elaZCCPd1GzuutbTXNU9Ga56C4VOwNw/va2D
OSLZfjte0Fm1rnUy0Sheea9kgf+5SxzK5x0TsoFAWMHFq+fyaxCeGXYlG7PZlVl7
qmmXCTmEunQq2i0w3rfJ7J+PSb2jyQ65i89KN5LeYG2bQjqX/zYOILKho1E9mnGX
4kL7saFdYYfSndBg0F0Sym66VdyRVoRxlfmH6k42mFD6HZ8N0J6gebVFLXnDDwg3
umdVPTLk1rrvMHgQG9CCRylGlce1FVqN0mLqApQveU5hhMOGM5EUkGtlgONVbDYs
x3685rVFkBShG8wz62TD89C/SwDT9KdVGT4O5VyG4El2eSy1GowM22GXGxGQGZM1
XTabcya3BdCmoQfP/iwh2beCd3A4HnuxcNkjeeBgDQ4lzXTqxSVkdX3K5nltLK+E
+oi/4UTDsugxvnvG50S87dOdiOSIzKlz4Rx6Dba3zEerdFbwCKhd5lf9GeZIMSVI
ssJ2mEexwoAIs9zG8vk0p7Rv9yCE6FRdhNNLi5A0s7WL6B+DQlcG7bnCYZg6QHdW
TvrFBkbJdAScm09jLB3w/1vsbWzmN4SkMyz4KlL6ZmDTKhVm3HzUP7o+Y8OM40Kt
31is4mHIYCJ4vIa8IodUwD2vtVV0SC0wSPCKgR2nuchgHAqmx+hTepihuVuc2FrI
YGdv9VQf9yIpEgMOQhN00bT7xdhmFXUBbmfnCTLyay4cIJCRvW+icKZyO7TcsvA/
iFR1ipAtAOHGwH/DzW9i1f0UhVcY4n+ufX7zLcgzJ6QyW1IRVINXdT8ao9CuOSye
lQT9hZMTsZRir4++2EK2bTtStzl9+ngmakGnRo3dUHHV4EkepvHo0uVhIKDZl0aV
IEISTbmFCJiOys9uy7yxv0ftEJND2cahZHQE4rcD+RAC8VV4O83dJPpciyyQ3wvG
0SBPlPumJovuRBzAWcG+McoVQyzB39Ehin96vi/En2NafOWYZK/FOdVdSqFSCAIU
Gyo0nMEwWvUrJlkDp0gJ0A==
`protect END_PROTECTED
