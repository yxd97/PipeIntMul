`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CQrq7EEHaRex2Fvaaalvl8ETe49ZmZG4Z7Qnzhs7Po3NJdl+B7jgCix/hajd6nOV
mIizeO4shmdemwB/kmDTrpdyTqJfqa+LAdyOIM744h7D2JjakYKlyfVGsF0zU0Rw
WwX7E4XPs3gWWcJlyJgCQZZbWtbow5jYbemgH3y4urPSARW1AkiMWy1k9xFUIId0
kV24sNNRfhAgG3Jvj05TxZaKDoTVoJx7nXlDk1DdLFzYLztk91j/SLvj5HCs5Zjm
t4RoTaX5jS9FTE3U622fpQa3F8fX/33JMxB5+OGzXws=
`protect END_PROTECTED
