`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AoR1PJL32FciMVr4jQBzhqGqIzUPIoa1nueCSgNC7Rk8mETAerYDJQ74KXwJyHyz
5KgSyf+a3c/CC8756D5TKFcuZ0cuLUa+o+so/voH6ZLZ1LPt0GFPqyIstaZ/uA+h
qEuOLQAOuZAh/wxML46BXYDqIIfcBgAD4u+h3fjAa7gDYdpVzZI4KM7ttpkXG7dd
N6EOchjlTX3+SlzcwtIargFItnZbOSbkHzofBrd1qHMwTLixZS0BvBnKBVs+e+2B
cyISwUTLju9dcGVdBA7USKgrBcGLslXEAEdKkcJehBodcC5xJRZuaPVixfIfB7s7
Dx2oeGx7mR3vFxcxwNf/dq8GNU5ZfLezExedwilPEawXp/4hGT48VrLji+8hSzsg
pqYQWNxtAyHBpxA0lGFLJlmwZzP6kK0sE/tLZfLWJM3sggxs0UHEX9NZLKfbDivU
DUIPKdsJRf06BjwY7hi4k14UWrtOGlwdbEOb6cBUqtXln2S0FsTNQRNR26YFQOuv
`protect END_PROTECTED
