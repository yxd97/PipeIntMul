`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wRYnL5k+Y+VNsBZ2yjQNmMHJlA1xsw159oVoye2x70/0Aa5hYLGiiyPnuY9HfwHt
5H0YivGBGANZ6w9rHvNCBr7Pp0NJKg9wUXiySW4hBVTdgBb/mcOM7GK3xadKDzzy
A4k45BH497U9X6qhz86MIVo5bLty8n6PZyx6ny+B6FyEmKqCjkd6izw4M7KG7+v4
MKfZYe1rkjWiQukUlWvVURQWV9mZJLNBeRIiG8mcRKSoTaiF2QZmea3rIpw10bRG
qE2BikKBM7J/ckambbSwkNqH9yqd5tJPQEZxDmzEkX1XAxal83+HyCP0NcJZOM8X
fRM6J4n+5m0JHO0+ZwMM3UorPezXZZ9Uh4jnHZr6JWLQbvVdXuXh1TvUaNDfSSjd
v8O+IuUIEhsdVNz29cwotWCqzsMP3GgIN8E/KtpdxS2I/odM28nQ8LvWc6ulL1ac
kbR5xzSRQEYXgPEOTA3tUpONt12qXAa+sNf8rGjTMdL7AHW+2fqeRh5hLdZGF/AO
`protect END_PROTECTED
