`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
252roOyipTZ2isKS4PKQdpXcGE+7UF2tCenJTOVEVGpOFCM1otMx6FmhLgS9nxIL
+B+I+q9lT3tR291PyfREAgcUt18Z1Y/DvnjJ9YIJUUQYFt9XMTp2Whipf2l6zTS6
8Dt6Hxp97LrI5uvrdyYLE3kYVcqVPvrc1qD9FQ6VKtKA22N9YQoUa/agRtZOtL5y
LJ4TKr26w+LZ2yR3gc72i9vJwAjuC3S832WBx4z+kd4cjcXDLjynXoCu7yMMnPao
cm47MzbbRLFIdVouP6A1F4+ViN05+YdU0Bt60/6W1MKSHo5Lyn25S3YCzlzX0GCg
L8CtcdS/s0c29ppWleqVXbzkDRRoyR5xibejNLonzlVnky0TfCaSC9S13WSe9Wpc
Hb88RanMqmvOGeyZH9/qEp1xgHXjuhf9VTAd3qiztPL/Bx1mKvazP7or+fSAATj+
czRV0prD4qviY/xqIY87ww==
`protect END_PROTECTED
