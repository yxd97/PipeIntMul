`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0NW2FSmstzLtCv3wVzLyTaZS1FLSXXdAOfuX8ugYdB0rUYvRfLQdrxJEgTzhFvpK
dtf2rUjpeBk89uEUey05hiH14GXE8WTdNpN7z0Vfd6C2kVesTBS+7nsx5K1tBPi/
khfoLGpKpE/pfqOVu/w0nG7V8PqhuB8WeMaWCsviTOrWz5AvvvneFW5byGCNLou0
j3LFAkfwlNGrV1e5TkiKCBCjnzE7LW1LcPqOnsOyLP9avRaEEShqfjR9q7ycgSvI
wnNWByh5YMaoRa58sOdHALn9Bng71YnMMfaT2QR/zUGjvjdE82KOl3BZZ/GjjI4Z
Ym5MHoMPoUm0QwwfKvqgntnXRrIPqtvil0h4RD7/j/o=
`protect END_PROTECTED
