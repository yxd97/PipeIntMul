`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6HZLDEIKo6VSoAyDeQjotXyGaan4ZOxqdmjrnQ2lWHWQTMSiPmMGGcvW84JW8zpQ
gzgI/40YhInrtBXbznL3TEusvITRSAOUaRBGvRB/mFsvSuyc4lMekWRNjByOgLUE
Laj2hzB9bKsuKumiYI+NAxcBflECy4iwUa2+n154xDdZb67hth65aKcGy8NHHXAx
IDJ3fm2Do7JBt0yVmx+/pOKw9DEoQ2jgmBAmS/jNbZhHGngfS4gg5nHZc+SWh4wi
oktCnt2P8v5BYWVQ7sPNCHT++bymn8725j9tZtF0JxNbdt6+X/ZqrULRjNHpyLVC
+irUhYusL1q7Ki2C3B3lFAw1Kfk/eBlAyD2Arezi88RJdpEGi9cekTXyCdkXk8ZY
94B/+qrvl9ldecwvChRzqurvkcg5+UKQphPtLRpvxAFJm1V9coRq+hMT0WHvEKMv
ACxAdo7Q2t4gsK1GHzeh+Tj6RnRZ4Ov+EZiaTdEN8q7QU7nMdX91YsT80hWhyy1k
5QKmNKXKawXUy83osMb+L+y2uS4q9296cJKnENFKxYSmlI7ZN4SqaVdT/uKVcR7Z
zxhYSyg0NxWjs0au39+6Vg==
`protect END_PROTECTED
