`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7shUrxmXpoSTWB0G2W1J1P5YlNCn47+8nUxji3Gu/NAe71sYkY3BQZTEUWyUp+v8
q15MzR816qku1JRpCTY3a/42x/sgYmRUAOzmhd2I/eV5x4UeV+EMR2IxU0ha5+3e
y4BNuleYiGRa6wSNXydIFA6M1ZTlSc9k0ay9jJ0Z3MV72z0pGFYLKAnpiN3N2fxZ
uyWDMCZyHwyLYD28UAG5c9zuROB3OIcYoZO6DRpEJP6e8v2tFZMMwWPLwbrl5om5
I3TGglUIY19xP1N4tcgVr90Xp3kG1salT2wYhi77LsU3gu4YXqg/1uFSsp0EholI
L4A4cmqSa9ZjZfHQelszolgx7N8JDn0JkUxVlwFafLQ6M40owX93GAytKcFfFZjw
bMTYJhN6qEWg251mJJuMQHk9jy+YVNneYmOYX/6O81+loTlQvDKJhmh8kW+B0l2j
OCkttjyAe76YhpUTeLn3MtcjF8vNJZ/BQbAgNKh2bqs0vcJCIaItM2DmE4GhiT0R
XZY1CIptqU3QeI566ax/vdQkr7JA+6DFiHtXuZNpIqJv4M7g7ACX45T5n0cxhe1y
WqXzrle21V8+XQ/VMvg8gz8HDy2XEFEMiDav50aKAcZ1QLF/R8dhLtgSEHU34R2s
Pe9TcJsLu/sszcfY8MBJHqdYXs63FmIA/4oD7eTWSCc0en97FCHZrj9sHop/s+lo
EvlVer6i78B8mbWFGZ+GbjDNG9DplNOFoaJ0QBarY+uhbX6y7L2AShz4citcngCa
iSWuXpKol+IuOO2ffe1fwfIFocDg7+tq6KOQHlAbjM5kxCDrMcWkcW5FDjmozLiG
zMBt3STouqCbnlh4Y+HM8DVV96BZeZa4f9DO+QlWYuuC3odR1m+N7PmAblxmIyKw
38pQSRhSszfdU1KoZBmujaMBpyNGLtSjIHa4nlWCdZg4qTkvU7dNJCffNHpItpmK
BxCtUPn5AiQxN1tZjvhUj8DZtrNOitYCpf7Ye1EBLgh331hjb9ZXY8AkYwpz4Yt9
`protect END_PROTECTED
