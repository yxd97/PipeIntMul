`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YMpPVgVQ6vWcYB22aI0m3bjcznDZNUkvLUDaZhOeJskUNl9yvPwEBi1KrRxSJNmT
t/8y8QRFR10orDQH2EpcvRiShx3a3CsORkTvWWtaiSFYxUl6mMjxI7yIhKGK0n/W
0+paX7+CYyQk+6Gx+jIrlaQIVdvRwMwNruuD6iiuNK/RkHVq8fR0AlaW10/1r7tP
sLPH9vm2J3b0GffKXpaZN4ZM3MfQ2/DAtedonwlbxIGqzPZap3rmeOPTm0UZXBGO
u4c21hdxnvzHb8iKgC9u51XrzwZcdupv4Pi1mnnAUlQGOfzJFbJtSqiBDqVhjuRR
MYlGS0r2j1kO+4A7WfS47Q==
`protect END_PROTECTED
