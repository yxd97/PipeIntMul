`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
alz9DqyX+nP6b5aWQuMp4arTwgfo6LN4f7OV2OueYjbMIQkYyp7nh7VmCoPqgMx/
5EkJxrMuNg0BjlggYHLUHlxUhq0iSqA4gtDki5dm4G1yTh1cs/kaDI6Zq46i9g3G
ffvqHYutf6eSnKbnj0msMP8LL0nQJx7Cb8fSrMVxuPZNBA68TgLKufSs1+hQJ+dR
l7W1gqwZQOrR4s140ln3jfx1DCnoCF5PM5uSMlhMZVbZitrr5474T+wDSrBEQ3Ue
LZV8hIl/+v5VoaVS0WLw37W0JR36gOAT5hqh3ccTuu4/q8a/ekL+sLmMlu1fGYce
SfgqI/wjHUqeVl680z7IahQmvEbg2nTylHN4AVjdmP6XF3hHlNwTg8qFcd6DUDke
C6GAmcR7E1xdnCorIhZlzYv+GiXar/ZQrzK4R1feP+dcUHi/atdPNLjXP5Np1qw2
knGTTLoKFIB1kSQQredQlvGbO+jEeY7rdAditEofwV8z9SJxIygU6gs+kfkrODvG
kINHFOo/RnR+HDLZ5S2VCPlmwcUPC0fZMBvpxm4AfLVhyk0ifYSXYaliPXM6zXwC
VM8KC1GhAfunaDnM1BnDR1Vaj1DDzDJbNunb4tQrtcgTVQCJlG1FTRmRJKb8gZ6h
8cL4h4wNdV2td9uPxCLMnnIDo1s8JMwQBpveKiNQ460KaGG09VmvAkOPoVuXMKgd
JMRrKbdXE+nbzJUOuUiLHpBcvSVYGeLhWIieEg2LSCaoJYc27zPAXJ0lsQdbyCbu
T0JyVaWyO1/LgMmNaVmp0svQN0ST4pUGpRyl2kypi9GU0I0/zgYbsSC0D4GVhwuA
iu3B1F1hShmryYiW5bWJAPwIbRU3Bi1V4/xXwm9pUNYZEc5r5GfAv9Fc0JUsxPb0
3xz+dGa59+lqr2EgB2f/LTjf+keciuKBrknPQeBzpvg0VroK9BjV0+gDBQnAPS8b
/Asko6NXY//ZpuzpVn2NBdWWsfcjMna0dZV3DA9kpei9SIv6f5wVkFDXALO4Nu6X
nSnTdK6g+ouGZ624s64qtyFgnpYBm7G3BCOvl+TVOYfTZhqU5CruUw2fsE6xD/Bu
A4NlSmgReVfnXpulBRVlhPa/vn2uqrcv+3mDu/YZ4TwYJSMjzAJ2joFXxWkkAwUW
WSeSUY29UszupwPyRgPFdGjBlOb0nDRZrdsUFnEMsU/l7BbTaD1qKMTNjwgjh2MC
fmhh4Ey3pX02JLFpDiY8HKyFryZzJTpR4uxbLCv2wswV4NiAcT6xfe2C9BamNzAY
POQ4AFWg/idjTp+1K51uwXFTr4viYhyIBeuTfEy7NQKY7M3vQnvT4AYxgOWc4fKt
JLtTQhWdH0Q6bMeRFBrdUcVSrRI9rRtVO0psPvmx/k9OYK7x0SDaZeZkLT901Dqz
vEbbd8y0a4/44Sk3EPhQd6zXRsSZMbIA5uN6coyDT8QNdouYgRN2Iv6Mu+xaWFob
pIK9ZPIN3RErUHUn/S7HxdRr2HQL4maStY8W/vptzrCMPcyB5pX/IBZumGvHrsE2
SCQ9rRgbMpHgcKpgzQGDaPKfMlyFYfbltCLxGvol+3BjF5I2pwpXlgNPKwKBmeXm
DWAuEZnJr8aoMVUrjE3xJmLXYT7VDsXboIsZ/8vM6xOu58EW/W3mGv1tTIavUdkb
+hO0p1RVXdlqyb2F9hpIL8FPV0l+xChXrPbJ6t4dRl+IWMJyKGMq1rDRRk39YLS0
l2ZeXOK4XixBcZLPQV8e4GpwcZtvCasf4mzpx8tsSXdcn47MdErxsbwlHgnwYCsu
pK8IeuiE2BTDFTi5JVHCU2jn2IZ42Boql9fB1GyqJK0WCjr7FG1COpZNMcmQ//sL
gOje8RKjU4QUXISHNrkg59UL0ML+DK+eudshUHStTgYEkRpmerJ+C26VEn4OV6mk
nqSUFVKhH3NhwuLYERrHmGA8W5SvNfq+uBNS5JsBqQnBOTAHU6tkr5IDHiXhGglJ
615D+fzPg49gDbqrTajchjdbVMVnDL58y0YDhwiGk0DpsepFVpeA/C8/N32+/Hjf
VmcJ6hqIU2vPRNz4VzgA8zUW4KVdeAQGM85S/SB11bMp6P+Sss+5XY5hSMHdY5/I
XOqK9RUlxPrzQEnnWMeo66xsl/Cn7IRUDpWJ/f09qHLN+PeMxfynAA4W1y54oI5Y
yqa6kMnBaryKO5hCJrRgNdLP96xc5DiamLGm8lpgRq/aM1TllAJwnBz3OaMOOX3B
vRdVDBvBaraCiVRoE2Eda9pUC+zc7AHtU6/ymJL5TDcbwl0ATyAYRrVB7eqz33up
3JVN5VbppbwO6E/bgsLhVx3IC537DWnZEtg3gPErHwC+YjFHnyW50+CNaBxsyQIy
j1UTZtVZZo18/TfUYTNGfEvQmR+1MckEBs6reH8daKia/yTeEWFviZrtwLRbtWJ+
S4rn9KriiC26eJLYbW1qVnq73RiHtqV8ug6FSRtf02q9mJqc3w9R6AoO7c88Hy10
YhGp/Dk349DFP1lylmg2Lw==
`protect END_PROTECTED
