`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IMavoFWFeGAjYxTdZ6yDg+Y3A5m04L4maiCOgfv+3vCGQyM+jlBRQF06UvJqx1JV
ca8uF/vOR8LbB6u7V2rgPsz9hwaWBUYnyCdCL4AvSzvOB9I+jf/1FszETzr31FW0
dvEt/uW6V+2kBbrDB+DjUxbtCbwKb1K1Ojv3Wy030p/Vu55Cl7md8Y531O0hT/vf
4N0LPnptPQCsPytXGd4aohaDGis5IuGZaLTVzLQF6qKMNg+ITKyv4+UMUDiaYViT
iCPo+fi9AkajF+3/wViZCKoZXHbNjjCZURD5HdKAAi9Nbamv4YDApxRLl400ry3o
AxQvUMTf4IZ27o97Hai5dBTLwb4uvg8Eo6TajZFQN87/cjMajsyTzfkxITroNqmL
1Uxqlie6TQKvvFqbnYDGHXszDlGhsXw3MFF/A/ww5Folafx/MZO+h9OXQACBjk7G
`protect END_PROTECTED
