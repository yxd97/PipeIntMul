`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YfMvyg2W3rAVyZ+2YIeVq/z+qr+qGXqw60jEp+PlEJIvBaQi64YsVkXw35ITsHUd
kDt1wVg6TU5WGh6K88V81f2X/y6/+9+CRRjTp0Qe7jv+zcasWbYYFO0WbYio2rU2
NpN0HqwLGImIC64OH946dGVjdAXBHs3raJCglR/+Y4NZeawy9pKNCeRBulGaP2kX
zT6gvHg9hGEuDZE6jFCURkFpRWnWYJBL4MJV6uAbs486zoUPFrcCRR9dTWbNa+m6
QJTq2rBJ+jGxRuEVauPIC3erK/+eM5zk4eW20g3vgpo=
`protect END_PROTECTED
