`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JlYdX0TjEfc3mBSS1snH8GAOrFFpYwy9sLJaTLW0tTEmLb9aEq9DklnBAE5aQSyM
ZAfn4/+2OsfBM88S0MmXwpHlP3aHQHsIK691LkdyikrUWo0c17QyIOXmtkCPcB+y
yIcnu4TMbLjeBvBeB+gym+5jV4xaTWNZhEOGZgrCPtWBYvw6GgyZZZjS3doFSrg/
l1axfGNeoih90AiHfruP6/hGTU9jwTeiFxX+8+2jLBvN2eBwPOXbhm2pKj+G6sob
HN0LDgWpgzuF84+bKXioq5Wkk7O+2+hbEru8Gzm7GWjKtGfOeUn+KfqrTkox4roh
EnCdyXZLXt6UkbfD2Smyeg==
`protect END_PROTECTED
