`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w1rFjFqWf6aw5e3cID5d2vwnzGYOpU2LF/ypUD+BgQD+gSN7vtECH/ZIzElq2z6t
84ZlbGxlD2v4EFlElmp9J1vR0sAk2j2bTRDBclU5Ru4BcGXnI9ydmhpxg2dHDvUq
zLjLIw6987xN/IiG5mobqBihMHvLbHyU3Xwmi4cCV1ueozwcPwTOPz/Zd7FR6ZgS
0842OCnFFgLaqQZpngI5ABtf97ua7fvRdOJStAzd5BTglqEEbOrlgJK1LUZhRv03
G8wLh4qysA9+E92taBgXtQ==
`protect END_PROTECTED
