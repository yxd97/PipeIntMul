`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WKQdVuvRwdgif+ADyMMO4G1LUG1Rgcd5MrxNSWCCDFAyZiDlyTZjZcGs+Ic+ejqs
DPm3qcMPxyIeuZq3xfM1iNnbP7tm6t0PLhcl1fTe2NFNvQ4EW600JVlLcJVcDlOu
yNLurx7iM8HU9YvjqNBIK5naTxzZwWGZtb972CznonuxVy/Lpo3zYOUnpuua4BWC
OtoM79M7FITW2KITkB9mJ6mCl9bxsiErQD6/RHgKcac6f9sxIkxhAyNhgdknqKU1
u3S4BFnOmcbWoZjYSmnpJ0uqFMDc3BCJ7kKhHH9xSLPzF4QPhE7lLrjD1oXxuacn
YzL9QphhQ8Xt6sknmmQBKBtIexP+gwKcko2oWtxTuXce4JAwjI3LUzhGR6hFyFf1
ArlzQuK3W6IRClngvXNo4AEiNs11bzTlSJxDrD0pVx3+uoL0aNqL9VMN91S/q/1G
2hQbQ1l/La0Zak1dTDZDF9YruL1rq2EksTgeAgP6jxAAErQ9uouTATTe/NK2VOpd
XvBw+nxD8zrQjcyi16r8eA/XxFAaJExl4qPbmcOqKIIdJNuB23UGtVuVcteIyi69
ICtSKbxjV+/JAkqZ7Oi3yD3Ddf70CiQA6wsXag1KVr5OSPPge2XcH22+5VePRmzB
khalwdQAXwrmpVDRBQCCzcBmZyG8z/te14j1bd7+kR5xUV1j1GVbrTfEnS1ct6Ga
6xoKElRUcYySY6o9ZAq0/4XY8Afg/cBFUZCgYAZdg6kvs42jU2k/b8PPo1CrrSRg
ngkjdAUgceRG21e8jKS3th6r4F4tbPF67sJgZt02YnX7pAvFxYtWhVL3bBoH4dVj
ajYftcYoqH2Cy/bWtPxZt3//fXQs8IAzN4JZbyrUdPbe9bHyoiwYBgGm9Nk/eNcn
VAjfuy/12NgImFqFkVpHvnSyNXqXdi5KRmVwWfvwQqkj8MXfv6B3/UTVXzx3oo1L
5/gaUl/vgeilbf7FBNEjBqohneOX5FPABGYOsGkSmhrY8G8LYzMUABWhPwOvxDWr
GQ6YCzgzZbg2eogIfcJ9+kGqh6jJtuHgkBlMyOeV6nKElP3BIH9NdtXeGwJHsnC3
PyGRmtNEPEwrSYbvZFTwYi22BOFkgnHTByE6WGlBJURbfV0G8QY5stvrOM69WfpI
J6bTdQ5OImN88AEJ0tB1dAXeOOFgUY2KDEi7HgFcHHE=
`protect END_PROTECTED
