`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q68/i0A+YdWmYjKe6PamzI+C88WJyT+7QPuNSICiSFoplGk2BjjSSgv30b1CI+XQ
5mayH5SNcBJ+BuDReZD6fRSsLW7FFlhAh1nord4yVM7pMnSzBryoRSYM3cjPx+mR
kPFgcTuC5MNw5IgfAYqrr/oLJQM8bZhqSK37fVoH8sDtHbnuAetbAXL6oERL5sfj
nSVoZRb7BZPXNxYaJgjKb8e2Gc4xA6h8owUL/PpkBYlpZ4OwNOH+rBGqk6jw7Prs
dvF2Y8JE3sevYUVHuIn2o/Orpt2cX0T1z3B39Z89APyfOBWnv1yqBIvvmulESCXJ
w4HduPkPzVviwrttV9av0g==
`protect END_PROTECTED
