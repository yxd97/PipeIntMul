`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qbk7Q2MXpvj4pDm1PJBLdLb8hEW26R3Ub7oFxrkkOdBgxUlaRK9T2em7+OACD79f
rKxhUoz6pxk3ls3PYEQGBHifmll44ii7UsTrR5ShQFMZ1bCOZDhJnTeHy4F9rLd4
T5yM93TU37yj8kQqeA/JX4awkEAwb+F2QPoyoaxfTRkkv1SOVeq2T7SQf863TWFu
Kr6La+KW/O/H5OKPhUc0+8sg3cDQZZ8P/IEZCMruLhBV1dOUlS/X3y3GD8v82M+H
J73fSO6g7tri/0f7Aa2IdQ7eUYpqgNZGRRqvVGO6b/iiJYzAs0hg97ZKazAberxV
IcUvDBJTHKl5pX5v54ckIelY6xavTLmFAyTKueu5jCZPeXn5NX8WrlmXM1GO7hNz
PjWHd/yJda+Mg9cYDz0qAKocL1UYZPJDBcnhhG7vgjkZ3ZT6QiCLbA0quN0G1HaC
h6loLbY5iSrsJqsMpDx/13/Ia4ExLa1FfNFYlIS72kjvgn3OS2wbq43dHSrixHDF
ZX7d38B7D0o+u59XYM7wpKbGjjmWVDqrPUHftiDFTl3shwieTUyY+zVa0REoFK+z
eYkM/1kT9pTWq2d5p5IFXRIpr8K1lJYOJLk0OM7MfCWiMC83iShxd80VXwxLDTpX
OaNw4WqbFUi+aIyoZgO4yLCHjVxyBhxPnBhs8t1g9k9ezSlffNmbN7dKtCSOTLNA
SMRDk/Am3nIU1vM4FNOydJX6iStiXGeFwj9myNfZiH+W7qITXdFx+qVn9U/oR4O8
YyIl424sq9r5M7aU0ahn84rTd9VSKEBNUjtPCqOnQ6UsoUFV8LdAT3kHskW83aB1
OjtPTICK9CPo38umj5cTYPSDspJh7fhsJUHk0u/VVBNFpz0fMeRKaJdl+6lwqtOM
7i7HDanVyaGFlmwdvRDPefkXEIHfKKIv/3SJoWZpIOzQBW8GYBYGrawlk7t2bCAS
RVwdQwJzbbgtrPZKO+PmaS0LJnqQUc+MHrXWIzY+FWT8V6oM8IAdh7zS6+YeLfb7
6fZiI5SBlMkamXTm12Cpji2I3gOwB1sXwjI95clYrtMKEa4LCHLLVXVBthpZA+YO
o/mv09Dw9dAtMYfLRNwtMWgrpX4B4S1iY7pSb6MYRWHikcfjO0njQgJvLevypMfo
eSUj+I/PzxFoV2TpAvOH6ptUj8rP12tKZqLmwxj7R9w/kuLa+oKgyU3i0RYbpmV8
eLqtpWyxLTQ7SEJnexlZ6pdUKsCHO8jAv5B/Icc2AS572nwHLRksMUDzIxrfSAam
gqjNAatOwojZWoeBtHF53LkKSYJuO4zgfAAI4yjOK6uTzMwLF0D+aXhNForHUa7I
Qov7KAwU2kDSEX4nztg2V/nVm8fH3mKEhC5MBJSDAopkW2zouNCHj9QdHluOY8Aa
oTMQyPMYfLfcgX4xJme30kv71SsfzBsIpn6Gu5iv86wRNocf72mz1i/r6Bldcu2G
DTomiYE9Un7k2cwgNa4WC5GL/Tg1RdYIxbeegB+TbE9tj2D12khOnq/sHvSnZQiT
0KPfMeHDjyOaX//JOkRgySyKJJuR0JXewlJdkcQTySo=
`protect END_PROTECTED
