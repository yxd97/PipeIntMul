`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QDlOQn8MNF8SF7vQv5JggzMmaXMkbxj/tPKV3uXWImjR5S1Lz7+TkkNQM/ZAy8Sd
M9DTmD+o8qbkbICy0Vp+90QE7pXFZ7hFAF4X24HmlpOdseUTT/AxPkuZRlkZ31Dd
ZPPKLn7VhHZvDGCu/lSm8Z+GnX1tQFxVMfQZ7c6UpPUufNF4SuGiQcmrEqNjybbc
7QRYubi6R4l/Z1hGI8vfEMtunBq5wOfoxdOhkAtIk/uxdI0F/82RxlACChp6fC05
28FnaPWeXEDCeFnmJvEYZeV/xZ8mqXfGiKKpWdJaPDhUbG9uN5CG1qGrxVZBgNi/
wFElDPH/MuFwcNvHAn9qHCTqtujok2M4/vTzR3010sdS6XYA9pJTiMrmSx7jHhvr
XRuLiJUykJcBDQFYMtUA2uaanP49sAI55aMWr6a/shgTeRifS7y8HhghgicnP+at
VAtB2pGgT6DsTGcvNbE9z6k/B759Y+VFwqpLAX9jJj8=
`protect END_PROTECTED
