`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zcSoiIsfOqKf7DeauGIaASw1YmSLnl4pPgm0AF5OcBuFL0FS4G2xCjgxY60BpGo7
KlZJ3U77Mx+sFeYj8K8dsikNDUWqZHdkplL5IZ1AY3QRM39OO6sHF9H8ixJiwiaJ
b291+uL6aQ/vTeJ4bWHM3Vk3iiH+38C5hERPM6ms8HKVKFlwxJ1Rvnaxs1jS2qkA
JELx0Zq6CCn9bLcxGFDaItnHo/6YmXhUAdVFFElFHzbuwhje52JgseEZjv2irmce
RDXURLdkTyumLadr5NQJW9usHNcqnn8EZFjhpiQvm4hwu+Ow7AaDw2QP674vPzsk
`protect END_PROTECTED
