`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7QiMU3UjCEY/Fw4WKM1otf1Z8gLaY65wnndhd9CxYbOAUhem9L9XB4uH5/kTx8IO
ES3foxF9o9q3iKPfsk99mm6DtopID80WH8ckP2CoHwllpST2mQeXTJbkLGz40Ko0
Szq15eAaGoRXppsPARAL/eg53Av+D37E8MG2D8mSc3AyINC6yOZR5u7BkIGk4vRJ
y5Gqo5sdjNCUgao4DooBPC9b8Txrvx7GvJM/UBUqvra9HIHPxw9J6bHdslv9kpf1
S8UILkfgpUIx4V6x3l0IGfH4Wlb2mh4yhCNMAeQ1NyTZeFWc9o8GjWePmz2ITIcC
`protect END_PROTECTED
