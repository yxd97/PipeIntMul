`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pbCM/F787b4DT8vAyJ5GNJB0blnr/kLpKe3VyEGHMw67aZESKX+nqytH9U/y/j7G
h60AsxA/77Pyk4eH2XRO4R14PY39idBh4/cwgTpA6kYf4lXGAEXJqLrQV8KfPwsE
/HNHlF9DoN6IihMLu6xcIzk4vmMXc45OOY5Joef8TfoQBAzHP01D5bcTq6LJ+Did
YDAKJWov5NWqdPpChAKiZv/KB9ItNjdsE9eXJX/YwqJbO27pMFMD9KX+1dNgJNKe
jAsz6eM+JE+QS76JEpFrBTnv91407BpMvM9DJXq8FPXzKqBs5qEI0Y7AOExgl4iT
jUKwHfy68Y+HNKpDbyQe0YHxzkxqW91TRBHBQwWFwOFcJP7LqKYf2M7N/JOVgWNZ
4L0Gb/NlX1+72FTxPge7A57T4XM+YfpeviaceRc53FOvDkST2baNsExWFNk8AbaU
jJP4O28VHmJOVJZKzRqi1frQ1agdLyxLkEI8voVaQKe5uomh/Jf6dfbZ2j1rFKnc
7l6GJOWbd7phWUGOvo3ggUUVajN/Oons0ahSjAVzFAEEzWc6H6J69a/ScaN0sybi
l41Ky8jKycUzFsldeX5VEYNQxH8gisUBOKRDoQIqqWs=
`protect END_PROTECTED
