`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tl4iSxNgiORJgh+QvbRgGq6reRk/CMI08SVgKvnG79AHQJxYpnuQ7LOaqAfyEba+
ls9aM8k4CW7JanT+TJNQOE7PgfGurE7y6OlDt2uO6PqtoMpZTUPJ//MzNQR/6eIu
b2mgWdgY+gPhsPmXIhwXNM2CZakcetx1SrpXHByTbkDlYsJBZheU6CBZODme2QCW
5YdqvQNScjRwyrxE6DuhrqYuw+2KDL6Qn9SvHY3KU/MGYOWHe9RDdy4REia0Mq4D
q20g5lyqJR/24fw41b+JjOaguJVHTxE4eDZzoaH2NzxAPa3CK1T+2L9qqlIMxgxM
cRQzP6/qdtUOZGu57K14hzVbHEVrqzJdyO2SFBBCY+R9yqjNQZHS5xh8RHaB23tU
gJ1lebzNkY77dO66TAxSwOoq8DgVqYcGJwsPp6vrzDtavWogprIV+vztl3s1+PVR
WldT6HrxHphIVk6405dki2HRoIyDrNBZpPsBPWIKGwI=
`protect END_PROTECTED
