`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CaE/DRfQEj92FwrKTOIXnA2i0VsXw/k3Eq9b3pjIQgPwope9e0h1HyIFsBMkMI35
oQoEVLyT9b6rd2qi0hT8Lpg4HIuHbX1d5cPhRq1I8KBxcF5bXQPUQSwWAWMPPE3a
G9L474DZhh4TObtABy/FB+px8cnvgivjWV3Seo+HYYywPs8bAKJ3cGKb9E9ZDNNt
2NEaQRV5+04zDnRGOkIBNFHgW9fgJ4YLqWRdTV9M9euPhbCv2C4CFcnhv9UiYPK/
e3xbo04t9f+y09RMn4lUgVIsPg7kQ7/gei0qiAt0+eUa8FUb8PcgU8Z5lcuQMisM
GfKL4Wj038kgKq/x9PnJFaXA5PIlqV1HU06WKnHd10hetT5QAOCrJ3hT9ERvsrhB
rJ76QnPO37DaH8ml8iMMUBihG3SqdhQgVxNKlwTsIY3/wgJjkqj+jSr+0imLKVXr
9B4+si7BinE1y2n/etCgt3S5VY4BI2RopEMyvTbBipXNwGGMKd0AZgCIb2Qo4B9Y
KXzGGfnadpEbK28bgV1xWXb1/WIqJ0WxdJWuUzijhGWsW78QrMfhoS0LM010BU7h
ISsmYPEg6S3GOrBoAEmGbdIO2u0Hl83Z/Y33pb0Hkhk6Rpj22wzCEF7JJ4Oxf0/t
xk2s8qXdJA+DmjP78Udjx42QL54M+15H2GbwHZX8vjPH3XcAYXyonyQ/EXh1/FRw
`protect END_PROTECTED
