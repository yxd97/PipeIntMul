`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h5wwLDXa7V7x3WUOVBNHhhiaWzMiQ67xlscZfdPAJn7wiMmzmj/h/F06MmkLAv9Z
nrbeWhdrPuXxilDu21eGYOUz/AJGYmHskwjt9bzdb0AwdCtDKqi94l0MO4N896Fi
ADzApybBPDF6yGbxzYGOWG52c8zcvGOSZjGjWWRNDyKYV5Hw+MqApItD2pRSSoxq
e7aMHFHMBh9yQSjXoths6nYpMSq6VxlZRe/z+DfRye9peJCFpRFIHu/K4lcymENp
X0fVH0Y1mURymkEcgrlEBmPmlDI9yVCLrHZphGbZrsMP/MLIgUNMnmC0fxZycz78
F0y+dzLIwWGdT/08A3FiwJwyEO6uWEb9M3104xL+dUXsA1RUUkvzVF3pTm7RSXUX
uidcDwN7MRcFBDeANS0TDqz8opx5n5DFXj4AaA4q/pSeso1n+jV6Ko+068sADcU2
0YVi/3lsF+77UsBMfefGRXn0lX7TTWuJaPsn50W9sIUSZfXAxe/79o5iKQlDePbz
oRfC0Z6MuJkFYzbhoHAKUsdfnZ5M9wdjXTwTAdSntoP77oX4k2QP5d4BokPcEoWX
TS0OsOna0nqdc7cIpi7AgyC0cdFKJdC9oNJXx94OqsD4dQ0iGAPe/3W1Yj2DmVtk
hjQwMNUDecYPF5uUWW6XD2Fhu8gy2ivyUduiAnr6CCOdUFSvUxb9Ipe15ScPWxbk
ybGn4mTRcezXrUrtRD1/F9UgeaiC48ja2GJ1zZk4ibcSVlnvcE4p1jvBMSDNpI1I
DDxIE8cVxzkPii/ocBRoZkgdqOXtGXjfYYngrAhE5NZGAtbuc37IJCD/RmYysnAP
IuvaH/otRP1+LTI1KAoM9g==
`protect END_PROTECTED
