`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1GBjAGX9dDhkucYUQ+E6+hVBtyO5ih0FBowPCH6Lk35TukQfn+oXK5rMEv4trCyE
ULiDjdDfHkIrdnG3zVGGKy+BN0o5oahU2JD0KDLjwyfCw18yDEpezhqresGa0fL0
0oowfOWN//nNOryFaSmX2Qu2A0BUKcA+3VCtxSeRihvhQq/qktwnOqD87w4j2otS
6Qp7WDFLFmVovqR46ilXC9dUdmGlUUsYqGgZwd0rgC0REYqMHGHcDOMsmQedje5W
`protect END_PROTECTED
