`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0PafM31DkI/sTievLlxhp46TTVYGNqMsk0Pen2+SUA950nPeueQRefHt/eMDDiR
Kxat1DI8+xGOyJlPTxfKAvp6jdThAX2RBRrzIXKkFnsczQD2HHiYtdF2wB396gFA
hvril1OC3VIDbv3HEF1hTTPvJ53EPwNVLvrvEAi4GAQnZYJRgnFWieC8zpsuwBBi
h9BbQ0ZIfVVrMrzGhapW907q10aFKPfdDDH12q1Rem74hsMWm9VxTHarjT34BFCu
IAlzq6HDJJem+YuOluFB8n5zHAdSriRwlMsXhtBlx3jLJE6ZQRcdROvclgq26gxt
X4AgxXH+c5kaxrkyWGcNgA==
`protect END_PROTECTED
