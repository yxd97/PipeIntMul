`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XBFOKjXbu6NtQ6dzrycZu8rl+GkH7Ck7XzPtHOGv657PdOZSv4/4azBl4f5uq2dA
otNslQ5A14bnjoRSeUojv0ZErO+Kn8Vy4yx2cZ+LyGGWkpacTThaNZXFttoIbid3
0GEqp7NpQ6dpYneSOj1+nf/gwHk8Za5Io+PvE93Udn69jFtQLRxgvZLAM+YlmO5s
VWTQXF7QLknJh8fvf5ZqN+Gm8T49BXlgdHEYVR7H71ieDQJxDbH6hUN49uyOlZwK
REtpfK6k9d4Zd65ne/pjMJ6Aaa4PI5V4FUA2+ZWUiF480k3fuBr/l9wD49re45ax
CCnXPfJufF6p/s3clPdwm30Dy6QRJewCJzFuzomS5o4d4yHJ7CFgxz2/ZW4ON5nW
Vorohv8hcX4EmpIhaA3uA3ZAdFuzfxJecsjE0Kf6Q1opGkY+l1PGkt7dh5Jf24bL
RIlOhFWn34fwN94G6oqKdr3B4TzLetuSF7+UMwoYBuCJ3mQQQhNTUJ3zPsMjP6AM
FsGeIM3A/bpDNuhmWPahy1gC2GGRbSMUtZfN406bSnB69RC+ea/IUQnsEsgt7qZg
lnNnjxxc4Mf1moWHsZBlHLFh5dldD3zj1tgax4Xv+V3J3dQDPilwQC/TUii+7fTN
/HR02yPvxmwfMs+faz5/fV2AV9JJTxA+eoPrWS93wewsrGHnzaMAmofYYxliw77b
`protect END_PROTECTED
