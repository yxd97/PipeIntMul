`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
29aFCXRul28VNlKX5IYOoRP6nDNSbtAOPBrHstwTp9P2V5feukw2DIcpt3hmkbPG
xen/5hYRNMg52TSlGcHLNc4neA5eaxoy9g035fg6wzgDCOMjx6ZhYKyWPCEqLUpj
zPeIf9rFHuxAPMMlpN9668V/UOEhJCgLNJT9cCAi9RujKfnYv0pIlCM5nZ7VEcAE
6mDiG6QVKUN+Xsa5FJBFhLUi/6/B5GZt+J8WxqT0AMQ5TOPG8YQcYGxJ5z0fexVF
GSyA/pyg7E5SxdDZ+Kn+nPsUf7/kzdRvuBlvGJzPsWWYYNzp10wp2JL7ZUOt6Hys
pLu59WQBVYsDoYngjxJ8LcCFuhha8lMRkNwpkffjUVSXjVeY8Ak+BC5dwAAQGuGg
2I6RykkhrEWUGgd4JXgoF7orDbBhRsyxJLbIsok6bp4w8oCxN9Vgie/kHrSr/bAo
QSJOrnwdM7rXSbr3vuz8ae/365+iH9id7CWU0U6uIYwniHF0xzzCZFkhDf0P1L6x
2xXmelfxIrrPzdYY0n+JXxndT0JlZ7mUGLHPosk+wSzYfXbzchitemNfUqRpVTxo
v3+2xg8SKa5C+eofeUu7pEzrI4JUISH3y9sLnSL3xVsWFzWXOvHe5d4I2atr9/I6
GQ7XdLcwVOOKg0CucY3JwWLW13g0mNQlzxPPNkjGWaoEdNfpiL+TOPvNcZT6DJIu
TuUTRtDxhLdnnP0JAtpYMq0IpwbuiE3ZkY44Z4wc2dUWaRnC8pHtW3GNkT5xpgqi
dSgiR1qpHDqP2oIApIblJDkIR1TmjtYi1YAQm/5RuEaTDFXqSFVZgGXAJOnWTNyQ
PtU2tWxtSgTOhiFh8SBm5E2oGkX2+cC3fIoLygyGzH/KW9W85dEpfR48AWAVWfPE
ArfULQ9b/1Al6CLdWvkBxIrFeY7T+PxRlv6q01I54VEjb8x/1oIXLMC8lifFDHkx
LYCC/TbHHstiD0ofSRQozcqzUQ+6OQYT84K7wALo8E/WCsCC0Y8Un0nRSkcsKyoG
`protect END_PROTECTED
