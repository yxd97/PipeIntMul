`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C/06qcH+QlQuhoOpmyp49/aeXMb9/hujvNlFnhyBjbd9tGarTsklU3p06rOy1Pjo
kvpeZGatKda61ZCWzs1bTnS+AgGAp5FKA5KphFjp7ubr7BlL4zXFo8cpWikuEqMg
7ZEWibBVSZEA82bEl9im54n1NEcMHBUpJYinyduSpZx+bnZXxMFhCKElrN0vkPKF
+uXy0otz4hg8l5ftDigI/7bfYAvlx04AGep5w2/0MYDUi8Mu7TcE9pPcxDIoZUwI
cKkQAwyxsHn3nrbrapl+AJIAe70HdUQi4QC4M1uQs0K4G8KJzJa8Uagk0q7xdtiY
6E7VM8EhJrWCDs+iq77t3A3UOHNz+FamVS/6KsBAH4B8RA4iqn0WJ1bWtAOsBHou
j+MbEyaTkCm9AEnNL+2hfAbhbcRv2KpQONWZ+NHGXCZKjUCh6ozkSvWV3Bu9tObP
ciyC+rrBSGhAJ4xhx/wna37rYIcJDQ2FcU/C2zU1/nqBXbeyPCsQbRYYTe9BahWv
wXhdv9Il8vhHZKk6M6sL/cXse4SMk40iGjekdznCfMItrcr74/fmSda9JF1LtZna
i5mtaYTh79vxswDbbM8lkOWH3Gd9EKf9UApTymz2PZpsbE9aW15yYCnfABcCe7dK
NkTlgnphn6tirikM6AlMgpx66d1mkgJCuJj3yMX/XEmvutcDld8xT5ffgIAgmnCF
t0UElWhQyWmoFRiFFokqVmf9PHFp6X8KpScPVQBxu53+U4JwmA1seJeNsGcm/hdK
EXUd3XlF8DnyWCFNvvK2bT6HX7dyj1ozcmhAM48v8N0gVvcEdjSCLihAyRXVz5DY
OgOdgI0JxMN3Fr2ffNM/aVhZKtGfa6iP5p4FD7ZRbTfISkOEXh3qXBwBKMLzUo7I
B1lHTD6660h/YJRfuyWfLjgcFZsa93W2y3ofF6JsVfenumyd7xCelSiRigTrYS3W
ADfQIqhzjuxMycTa0rQxzBTOKPEdmSaBgj1TW7uUry4vo/ED1TrLnNhIWH0iHRa/
49PGP3M7oCrnSCDwTQ45UPWqDy6BQf4bbaDwm6HVv0/8OXNCN7B2Cx4FDK9vuJhj
hIYQMZrVul8hMNuqTlxHlXPIywBgUDEX4o3l+vCJI2rAYChGaKjwtAHMmVQjqjtW
FqiQroBYoGE6kwHi/ecp+zZY2ymMV4ZyChkjLfm1CatwI07Fz2Toq5ZJ16VthL4y
JFBTqjeyTP1gP0so19q+0dwYkLN1VkA20Fl5SZ7bsFn7F5jrJHXtlgRBhdXjYWFy
tNd60Ucj4/8+sz7yY01tt+/qx46bEbJ5SD3iY3GUi3azpRKpcEvo0qZMYk/h6OCc
aYaSSPR04VKL1WJh2y3fGQa+Pv9i1OdwM3byF6qm/2X/VyaopPfU5Jj/H1FQGEOl
tKKn3Tnay5hi/UPmJj4bIYHjFiolVTDJNGE3vh87nGbb3L/ImguLPGXpTzv+R5x5
Y8BUmPiKgmjeybCllYgZrw+T2m0iOxne5r6Wtm69N9Gfu7ldWL8doPKH1PZaoyDR
`protect END_PROTECTED
