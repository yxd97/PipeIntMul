`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
15dzeDSGqKL0As/vJpTagQJ5m8nTg+4kZ5s0Jl3687KMu5x5dC2bFWiPMNHwSC8H
S1PnPVZU8/d8vHsoEgjBAl28xYghe3s8Vea9cnv7Ogx7NOTsISaDtjVvJq2hgNhj
mYzco/IZ8tRMo0p4N8xrCFw0yvunEWFWVsWyNcvyCqhKS7Zo2JyKQTwo2u+u+JjS
aA0jkivmGxxjQrio0nuMuxqFjbLQejWACkR0s/+iG0DbAdGV4Ys9SjJgo6K9T+vZ
iqVATWTyhI3Bud0KY8ca0u0ImvQ3cH2ZFfbIvonpuFfMAb3i0nrLE9KyGDS043f5
GzOZhciiMF5b2IhfymspMd0g/rbiwAOA9Mx8r8JbcTO15OL65skvnhuJ78Oxk02n
ftuV0qjlcWHJZcky0/47o5vUDcdMDbVmQtCwir0uOePc7A4IbqRyacHjdGG2MvQp
2fOTGABeKCBe3/R00Q7yp86tnuUS6F8qzhlAnxtqW30bOuoxFdmCDzoT+Huwy1az
`protect END_PROTECTED
