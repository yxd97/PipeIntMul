`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4EFZLRbyKf4xF8clPvlxgXwdmjHEqNVm0QilYmzVFaFlgiQfniE+bc0dcmfUQ23P
EcvptcQohCZFobKogZ+kKCBHMeCGm99whmi+zaoKPLWk7CI4gB28XQl7QhVX/hrB
eQdPy0igXDTdKgaztXf5spZvYZsFo8gdokAa27OC4dfWCLQIWXEVGe/ExnDkL4NR
xZQFX6ZJniUz1n2rT4Hp6BDzEjX0Genm+6frjPIoT0eQliVZ4AcdmtXQd8H2yCox
/pICeJnUj6Kj3O2Ry2XbUrYyM0zWpOtIOIpU1VZEixbmEqnGC+Zw9OCGl0kROw7N
y75xiTADeX4M6dRP6bGNNURaWZcbIP+qYzoeD6+n3MllBKi5S/V1Lg7HAXFrw1Wc
4rbZUHRyjB6AFLvxY7eWycm/pw3zaTCX3+zmGaps5VN+woFL9gm83+yi3hTnD9Th
+3ZRlIY70X+hLDPOij/WiEe9gwa1LnDgU6f39IsEaJE=
`protect END_PROTECTED
