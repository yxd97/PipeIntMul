`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iP2jKd6A+U8/ToFp9PPxfe/0wGLAh/NC/vHOquO0+I+fxyt3/inX9hWg4sr2jb99
ffHfSHNydcPkPGpqD9r3aRXBWGVxDRHWVFKzBwqbn0DzX5FvBDy4FFVP2TcI5ixu
MYBCiLFmPITxeHbrUdXzXjPk1LienchnsjdcUnVaciMg7P6WrOZt0sNmumfz3+ov
wgEhWNpnXP+m6S625jSOAE3MZGiOTMBlEaazT0BcsnZ7y8oamWuAG4gF00yE+0Zl
dTmO75ftl8lFGRy7YSr8Gg==
`protect END_PROTECTED
