`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ui/5bVs3R1XJND9mgKDhGMxDmvdftgyavHlpNO/n7NVjU9gKGcxhMd3dl7g+vs0t
ofnBYw/hx3DMWNBbmc49Ve1Y27PVRVtI1EitwELg1qt+03ygDMcz+qUfAxubaI3Q
JPsPPVSLwY7Rk4G0Pi0EfrAhhMt9lM9HEvBCX/i1nvjC9RSxML9cKp8vEyCvlDwR
R4ES4/15rtPH3jjV5nmsueMvdNs4Bj5hoRqshx8HpXr+EK8dILxSq3yOBFPjM7+v
7HEg/bdDCa1YyX4YVgq/TFxCC5Kf/AkprruW5OVkx4ZXqEpVEgo/0aMk5wlGiu0V
VDiDjFsadgFUHikeKY5zwx4PlbIrE0mdT0wCX1Z0/2NPbfXbY4eRBxZrEPpLv53h
ypwZ8Vr+QCF/f0Z4J6YIHLIrVDBRqdtEhiMaE8kmNb3tr5eZXKpEnyyRQCbMUd7P
Y2CPwwrycfgi7+cdh0VrDYjgfW71Pub2XJoYE4ij5Fo=
`protect END_PROTECTED
