`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t+B0HO3JMs6CKcgy/ZuHYfllVpuVgVWtYXPIal2mpyvjg98w/hXc5ofrk7vgPQhx
pje4XllbZklN4sib2rygpzolJdZfYrb9dApSY6KDo2bJp8LC4jCXQKgpCvjpDgDM
fC2WnEFBgn5b3jZZjFr7sXJzTcTqPmU4h2diBddD/WQl7GC/UMrDAsSBt85CcJgk
FkAubIPAcQWLbZkc4xbmA29nsKuxj0Zti7PDzg5XpDz1jclfnYJ5v7InkBxZHL/j
y8DS8ZBTZw17mbS5agAgv6f9RkKKUTDu/qn+sX9APuUVGhPVc3F/VTO/guHgKPEF
n81qYrWnTId3wvBbJQQ6X89AW/HzqkiVF99//NAvt8T8f6p6lpz1UMIjZGdW87Yo
5yshBC40IkSc4hjtq615JQ==
`protect END_PROTECTED
