`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lciYLa6QDxSLHa2YXNm9B0bGqIZIwGlxjWTlu0aCxFrvMwv37D/eQWrg1kT09z6k
34PUArDVn9C4zkXhHys6lsqR4nQCXgq95jZmDf41E37grHWkRD551GUTVTdT+FmA
vWEB1pnOze0yKhZrTuJGBYK5zdO5rIwVk1d5DSU9NpaRIU8irrsVh1r8tFBwwfr1
pkcO+y2FAK3ad2KUZJts+a8E0mYRNlHMSe/vGo0lT72eF4fApWFmItzGJJNj0otM
zMUaJkC2jMfdrClfT0JI2g==
`protect END_PROTECTED
