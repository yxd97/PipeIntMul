`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2kqCJ3jCgM3zmxXciBAIn3hiPSjyfItucwtqVWTs3moEMRqvaT6eTAY4ESQ+32+e
RDduAEnR/EGWt/D3xAyMr82MZjv5+VZOrFlrMw8DIYWW4apxvIXp4zkoN86d2nVb
LuhKG6JkMGh2/7tajseZsCP67mzZDeLA/t9FN1/D+kt6go5Su6pkPV5nLR8emqD+
431l6PDoyTX8moQuzTpgI9OAyeJYw/3hbV5A1ZeP3H0kqdZJmgmxayUyeZ2Fh1OW
/eCS0QRm6GoujKrU8oL1VFJh4YP8s2M0brAuTNkmapmEhOewdjEHUT2HaTw3RFBk
4QZ4XbRbSmU86vuA7yf4HQmyFW5hW/WsWPt9O8YQ7Rlsc4PgE1JlUaTJdkh7/1SH
`protect END_PROTECTED
