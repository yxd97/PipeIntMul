`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7TT3F/PJ4DqvqomQfS4a83c4nSjXRWjculQEwEt1+u2TpNiqAz3kbGtB2SpHNoS
dUTU5zU5layb1eUa3YX5AmRr/JFTflk+M1U2j3Yuzn8CRx832tgOxCxlhtyiUZI2
LYl0m0zceLnHpkWE9K/TsQ==
`protect END_PROTECTED
