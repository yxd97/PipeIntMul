`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KRofBtXU5hDEBNxw2Gsx76wUaRQ99+cgUrYRCfbxJnWs05EOjpkGkRYuckrWoULI
n0qSDDm+lp5HZqRHVF8XJe9Nj6tAda7q8FBD0kAIqB7X6WYyQA3mf0s+mocMXroY
ExRNYU4sxpHAsYWIMRAKl5HB1O19Sv4KNe4UOmes7ILEXS8IIGpMz5gMc2e9nlkN
rUL0nZx7wn29DLMRZdHqk5UNmBJJgBhSVQIPu1JqRUfZXeMc/vuBI01/k5QLQ0L2
awbG1ofK+3zheh1vFcj1wEYqEcnu0wGdZWT7IfCQTFF7P4nQ1x0m9HHwVTrCDT15
3usN87rF8XwKqXhFX8KGOX6UrY1+t8wcdj7Y0qMRdB2BW/u3r/s5EHHpoqnqIcn5
QHhU4lazTH9oznd6FmAVye7uDmdH33WF49W54MJwpjV/AT+LjiBlN5VepS8qo1rg
C/9s44C+HMTjmNJ0Nbg+m/l6b4G6dknW3RZNm7CCsH/J9/tsl5HvP8J84xmr5ven
rlpgMmZ6bUoXenhFcL1TcwTpRrn1JyY1+AtlDK3CbqWu1TmMXU2ZeFSeqWbbIGHI
OPbeEiDfszro4GuSOMbZqjKW1MzHcn0tmOq+nZd1f4O2l0O+Knv3qg1yguiMdWgx
J4Jz+6wjCIqjPlFzPypZVMYiIZHnaInZuX8iedj/nkQpvN6gLUAe+RTlYzlv+CuW
Nq/NSvq9DKO+BoLwVaNSf9bZaEYqwVWLna0mmRUKxkGyTvavIJI8Wm+YdlMw5uEP
B8Ra+zyrfV3CYJPDu6YRW67UVrv3XJa403Ao7N/A713XAMYqQYx7kTb3GSvuF0b/
WnVBbtZwc6Ub/fj3gL3oqduYt+vTGCZclgj9DtFIDpqlS8fLrd3Vk/3NosHwEX+h
WvWUkAxhSV/IS8JawXTF4CAehFHO2iM2f0IiGXq/vgUtShX4RnU47/LVUGtQZiB6
buExL+5dekSImCYJosVcmOSpP9tmchq5LE6MK08V/+xeCMXnH0CvqHe59RpXub/j
oQylpiR9KhceB5PLa5xfxlgcPZS/yQwue7xWqQxvrUbZRLrn2mpURnkNJm5WF1od
7Ho8B9mhQ84wApuILhfQjkaFrCU5tIBkjsMtRR7q0TK3BGV21SUINHoVSUKV55dq
Gs8c7L/eWJSF1LshVlarLp3m0zuKNvco5b0vo3EZrceQxSZc3OkN+0BF/qrkoUEa
FaY5UmxoBRWeAXmVEy4vdks8Ivzt9TvfTXazIjk7i+b9JHl3sDD/rBR3HqGzGldG
qq/iUoVGqV0wiLm/JhTh0wrv/HMqdwH9PK9P1jiLrsKY6Hyj3Cl/tXR/MvHKDuOq
oEKhgVCez3AsAZJtaaN0Q6g1QV+pBCBHj/ndrOUc2gG5OxY6bzH9iis9SLiPKnWk
w5SNM5KJHLFglcMPSKCq0s7LrBaRJNe3/soigZKwu8xlGYXvmbIChXLDobYBQu0u
WLqF+lP6CfvHSCaelvnBtXooAJdibTf9fNw5gL3uNiwdCndZrNfu8TE8KLibcUC3
vyPeGd75OcGgHJKk+vei98XgBmjxBwBOQuamdr73gPcVn2no0vyiLU9oYTCXfinE
fNNbCzBHyCflAUOxvBXG8Maq/XM+KMS63aBALlJQghngJfJUJlvbTqdnl4OeaCfP
slklMKgzyKIdIBjGQ1qFMNoDvQsgmuWW6Hu2LCHCj8WlbwcqBCPmIO/dMXn03kq5
AaxVOgtUF4B+80+VH1UVpLgWNi1QkmbQkl6BQxrrKwfP6mdzLD2cHzxU8lh1VMeJ
xuguQfMPgWWj/FEcg6CtKzfkZZpSnbRgo/MZGFyxeBMWWxpyoTHNwZKd9/fGiRFL
Xn5GeukSHvkWz3WggtPgubLNLdgWcfE53q7F0KVPDxIEm8+nem0mh+5aLlDZLUBv
PkNbO+E7Kfv+CTqgCgOcoEgQBH/QjBfChpuRRkVgA2/foBDV8IvGirrRS90EofmH
oA0r9Jp+UUe3c376/Vf3KHLERRYp86NbI0LSDViV/OWUJPXpbT2hD0ne7c9djHqL
ICM1GSfHu4DyMwGnJ0eJMip3fKl/J7y8w+zLJKHrdAU=
`protect END_PROTECTED
