`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tKefYje0wUObG7+8ntERT0CM+Xr6WhTmUqEibcJuND5IPOqoySHRu5lCnCsKNaVs
R5GZbVgXgG9M1FUnX8jfLPAjSArP+YKe9RDIJmsES4+SjV80Zt1W92ismrYB2Kal
Tibw+iqGsYLA58S89A2dwHYC7qmOpLU9tltPlCMeRQEHuzs0hnvAvkQ4wrMUc4zv
YbSzb8/Ikx5GsdPViuw47wKWikX1Vny0lwg1s1xzQTo2I/9Jk4nf2HGxZoqe2rOT
q5NcL3F95ytxXICbDXvoOAUl2Mpe4YcfMSA9mVX3cHF3u/o/P7B6a2vjrbNTfHoh
CiWbuM5EAJaSiw6KimsGTOEQOtRDF5uxsnzbvvTFpc5BVEp8cVlH9GwJp+JX7NJ3
MI1Qh1Enmh+zCFXmkbVR873bcHGRen4sAzp541FtpF5U4vgjmYupTAa9ZOQ0z/k1
mnGU4K22nEoC28tjZhOfgzfipHZOUT644McZBh730QTroaC8Tn9+wyjt7XDCk0Wq
0OjKMT0rxZG6CVqF+m827Hw6xicOcQes5pHMPPp2OcZJzufTM1wowv0eXiSnjgZz
2SqmAoBEL9zmPgzX0f+p2QwHRd5K/v9YWnPBRpLhxd8eiY2uxA/0za6oz0Ip37zp
tNv651Op9auSSrzro/ifIw==
`protect END_PROTECTED
