`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GlDwiulq/bXoiI7KLmRKN7Lz3ow3ctEBaH+vPtDllip42OrfVtdljUKr9QwKwuF8
p65bR9XnPddAFXUYwpmvzbvDIVrSXbpmvhhraeNpA2MHqfUE/PqpPyCDclqycXqN
icCCtdvA+OEOvwv1XC1fBBLa+3vJeUzyavVrfikiL7aA9WB7zqOBl0R7mDucI6/5
MIAhcBm1vncJT1e79psZn+MQ4itC+9BiBdXKnDfvASaprX5Qh+UI0pcw4VRblVxl
n2h2zMl58VtARQ+mqmkhONUGifFXKIUXBUma/PdW+htdB6dHxCeqtcDgnprVcvQa
jNHGxbBpIcmkIDZEcVMw24Np4wYbLdh7vkKpPCW37YqhR0retCEBfLnwOOXByEKD
BEctZWglEi0rzWzto1ctiMgaPmxJtD0ZSetN5HwpCUeUZm83Mvyi2ZgJs42IAW9R
q7Zm6eaZ4rdCnC6ZhFq6uF3fUahuL9qUUUscb98UvQzh39tyIPqOY0EoeeOBsEeT
O3Lg51Y2tvd5wItphXHPQK1xiRzhPC6zcod36tkLdjMaXZgrKIFj4IMWhtV12xhg
5xgT7Y9i0Er2wrA2jkXvqj5HkHz9tjduLc1dbO4gOWVpl3K7TMh0bgYJjH3rE0l4
LzlPazv9//W070+jDZ0L2VGcu+0USQYRuKqJ3jmUsWZt14hs3+aUHsca42kZCR6m
1FgkOnPOzBcmLlWClH7SA76fc6capfOsSht9G9KHzx4D/E9rZFsdE+FywF7RbJdS
jUFeqVNJNpcRMLZcHv+jesJdiXkRBqr3CvcTPVbWyjHG4NNQ+5qR2NtXGKnRl9yd
UoTiDF9dDlKoJOB5BXCJG3mfdVplPqHB0EBGvdz9CNhPfYPhak1mYjZXi8ABtThb
IHeUzH9eyone/y4c+BlecjB6PEnSWYr70HwKnc+Cfs75p1Fg5xl9S2VnvBD9L06m
64jh8/XsqzvK3MRMkS+stA==
`protect END_PROTECTED
