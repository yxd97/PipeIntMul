`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nd0q5Mib9zPIktaBRSAk3D3oWx/c3xJNZilgxrjAHpl5gtMdSoUbpcDKl2QTdjsG
QDcEpIlJwr+6ECfPYef+ov0D7/OcyugDjvj3GTgGnhjXbEoLNL5EbzDVO1Df+/nB
M76+GAsPgJa7/PthyCMrmSAwU80NgkAohGkJ8XVJWlj+3YvvhqZswf8lLpsoL0ws
Oz+yQqq6LNz88zQmvLBcabaUCGPQaKf24I9ahd/mXD6gHow7HifVnJSDXpNhhyO7
w0ox8FuTtLzaHGKLU1RK4aa7DhZqjngyrnVXHKGGpoHrULuQG+f4lQwnZFCWXy3D
j2ldiZgCITiEr6wjhjeAxLe521fKolEgGZ4Vh9wfx1iKgEX2WdqDy7KjxPQuzDIj
fCA/tYqdFZm4mziwXvYfccNsMvCqqmXK4TpeUQdjXNPLgcOomMH+c159/EKjWDz3
Xdvw2beYDC70tFlq2yVeNg==
`protect END_PROTECTED
