`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k0gAWMl9x+lgBghLR/uSA+E+wq+KwH7+6X85/MzKA/ZD/jeJCuFXrWWTXnXHjSzv
Gojf2HK1QKbXfQgiB9RNPl5qU/X2a0T94Ovjgqc6TUqqDn3eMpRpL6Iz3jkOE/FN
PlVbxsNiu3pKPlUG6ssZlYNEtJEwduddAoOC6UaeBGvdb9gvlPkgSKdRjWqDO0oN
uzwpEdCq0rxtFixpq0UqipMtPOusLS9ajsa0y8q6Q5OfF5WgP88q/Mbkp4xoSxuv
XCZTrGjXBuO7FC5WZIEki9jG/BbdDEk4nJupNcdrNE7AwolZa479LcVV0x5kuibg
s8zfQaLklkEBcQ36ywO/eSuOboCHOv4BMI2nJ8XjfoHCkUAeD2zlJojoOoWYuk6z
J642BDT3CU68XjGopPhloz2FWToZwAHqEYo1aWV6Uhok3z2Csxj5pvwEJB33YuRE
71no8ORs4PgIW/JlY5h0w2Dv5EXIeFkDyMaec2XXAujVUmvY72yCBjcJR4up/plu
lInLT7uzi77FMldMYLg5qLOfuK5tBQCwZbihiHjitDTlpbKop3nP0TCaPemAjjzf
GTXKpuGhLFDvKkR4scgeHZpgWj4mQ501/V5cxM6zt2aAGMtzAhohMOIg3Ug1uaBE
xbdRKafMCmQywhP7Hr5XS0Pn4gSXN1/Lm/BlYJShu8g+FmSzTP2iDM4xrsfS83nE
FPx1lo/e7Q9jivvmEmStMCYk4SZ1UUnNJHoJK/EeMKVymX/echBk7lDwl/2Cru+n
86YxyzlUlSE76x1FW0kxcF98P1XgDUcjMMw1lwkdpf7fRKnDfAwP/5I1KPBbJy/k
Y91mowdgAOfbICP90IaywCqARJBsroa6VSihGBEGO4aPsK1j+Qu726a8F89UWSVA
2M34DdVL+lK7FQ+WvRjJzL5U0ew1AQE3VU9zx/pDDhntBWmZQuUMCbtYw4xS+uvA
bwxG5vmA/Hx7rI+IdUxB5LulJgSh21j5xmSS/4k7vPHb1A5sNfDx5fbWfBtKI+GK
a3/CP192c8US9aPnhgVc2tqYVdXPuSeztUsk4khUkCEu0nCSXlxgoWM4xbO7vrck
XtEit1fGDPC8PzWwWjJ2n/xMQ5qBiVjN1AvsRRTxHSp48kDAKzJ6+2J1mf2c2Lo4
A7a7GWs9yRjEmOkZ34w0Ppd02nF0fxE4wZiygYY6J01JTYXPHZPFhVBihwt3i4ez
5fo8CYOo8vJcDEnjhgmIY3l6Mk7JN5QhJyYcQm+jSdzhmGqoDggtNVopDgyDxiI/
lAvtgl6Nr8YQwG+tQhGotL3KYcJYGt2bm7P/nMb6n0S0iKxox6JrQhPxC3e5cXZt
gp5pn0Z/k3OxPmH7F4Iyxp0dzP8VLgGdqS4UXulR+PGizhzIcQ6JYxRDqZy/X3tG
1A9rD5obuX4V6+xAsatXwov2oeHlah/RkDJIzEtoayYMv2bgIBx9SFHGsWfoBNQ0
52PKsV2EC6ta0i75iRXXHL20+4rtZidTLU0qcXJWN6DSfH6kbs29yu8icgGvNDKl
ajgYIhLTNqLTInwucuH9mZiB1d8Dhtqa85XbBSIG2IfWtA95sOLgzRumx9uZjDfa
WOfunTayXGscCEicjoHEEG2XEdnEQgZ/HJjwyGI68a7x6X5Hb2MmMpAH/NuCqU3j
di2Lrto9zjknRyQBB3SvluRlChHtLHu/b9GlGaDGhlg3QfeGK2LJx7O2HZiYJpZw
UDdXvQIjMmU9M39R43DbjI+PpbpysHhGOq/sWRpY9gz9D+JUHJ55AbvL5bOv/bF/
1WAByxkwZ5z4n6SPp7+9tPmGSNjGWS8ZyLiTY1hUIb1e7dl/2iyKvB+tIPDneNZY
tAbZsahFvywcKyz68muB9TrL5wL1J3mFhTsc0HRvnGoebCCs337oepkMDaWAoTJy
9jie9VeU50IJvTBMC1bzn5MNVmG+3RK+AOQliS9sWFZQLcCnHXewrQC3A/s0mLta
JBIdpOGsVGsodhTZneo0fJWKcjXk7VY+In3f7GlKp4c8NZkBWKmcVhNWN2WGeQnG
gCVjknjY2XdAdJVzDLR2juID97qrA4GgoSlj2MgvOpCk/AJ6jvXwO8XR9R/n25fZ
dYEwY4IAs7yy/6q7QZKkaHag0+nMLwmbbqeU2N0JvNkmd/XgMHtS28C0+KJt+3FK
arZMtkdLY09fpKGmcG1FYnzoGtdsONnF1vgYqzw2aX9bX1s3RN9/B6DJHdjR12Au
2KTTygw2T94H6UW4t0+2aNcvq0S9WMpg9iKDiXAYS7UjAEjm/cmXqStMh7LQVrNI
EL8rvgstrBglJcNETLDFlyiUXV0MspNxgWrlHx2nQr0fWed7O2qmiMrZMMUQgVQ2
iBhRpEilkHl+NGDuV/hyQW97eZNPx1VEHXu/zT97mLTXKQDGWpNd3uUu1CFQVUj3
/eJeV3G7wQX35pctY3nZyqfmwsUflHrx/fcW4dg4QfE/Y7SJ3zgYzLgOBB8B62Db
r4oh7X8KWqvS5xhmo5hrXi125VawZB8FHuMyCQ9SN040KYDJanbas1fkMQT66ivs
e3Op/0ocS3mI759+9Tq4VLzNrxZ8gBHiKy9qPWTsikiJ9f8F4aAqsYs/VX4k1vbd
Ld0x4wq8+aXpDJA0YEVPEotfs4Tq3ZyRmqfgr870XUYgs6cCgOmFjS3c+hcNJxJt
aKnWY1D9JDgMez5HIiOamDRZ4qxfFGWndA1Qf2YPnuiG2peViuAZ45BAwVOss+EZ
wJj6D+1rLpd2MBL6kAQv2mDwfCPYYki725sAPUUGoJ8SDatuUcWdRaOwUbZwGeIz
VxzHE0Cjty6BEyRWsee9UKcR6az61Rqk4ZkR8u3fl1UvJlj/E7GAy7zXGTPL0uua
It4lSs/ONNNbBmWi/jpKHovdDcPBSzt1WaOYvMPPZrfg8h4AmxWpfzTcEMEcVQcD
ThBLM4l9je2TMoycv0bm8JdCsitZKHLWB9DO7uFI7LDlLkukZQhCg70TNtnwGtpo
DZni2DfWU3R94RE5a4hNMdlsMnKibJcAUDmAlPTPfWNVmn3qb9QZp/RDowKlBQ2u
orVRCBk7HPgggnJe6nZkxIoqJ2u1wWYDSFIy6xlUuXf2vOZxrZSoXZv3VPg2NUM8
yO9kPA8bn9N/XP1TrmcDhovKAHvwF12kyaxyfvfeJPSSfWCcPt99kGRX/pc5pSjY
4k3EISqv3/GH8wI/OvmrlNi9QYwxRiOlO7LxLbnfOf4FAXvvMVlEf9pl3A8JYyek
5Prf9cCUNnMO4fIAebtPo0/qbai4ZtPcRef0RJLo0Ho07NQ+wfHWW20FcJ2/IVPM
tfUgbE1jMGLd+WBhYJs0Evn4in85HMoexRxNsASziN7kjo+fIFHM411ey26uMegE
4wnlGTrMF6ITMbYQA1VILs8IX3R/FBO6PkUVLXOeBoNlCesuXeFKiGChhOqI6fDq
SnQYJI9PGR9nU9Zx2zJBQMijR3iij694ZRGoJvHYJ1tbLNi65nzwL+Tj8pEqIutU
u+pmwabpz5wm54Vt54EOC4EEl2ozBKEc84ioegAKK0BHc8dO/OitbNVkOdspbHM1
vq8HmBYOLss/wWc89Ws1ELN4N7i1pHaGi6Kf8H1LH6J94iTG5tjmfn3GBhEDLdYr
3Vva2YwCu4zjqPghtM4BvSBplmUpfHG86S4mSKdp+jQMjn/zCjgubenz6gaVC1Wv
yBjC6yfeqQMPIj4zvrou/WG3OWxWAq7KnZm/yp40uJMjj3ah9bEkn3oWTCQ7UtoV
y5xI4RGYghybxjLDtyBmgmJzoD8C0YceB6EuFVfvL49NtnzLRb3udIzi5/ACf6z6
VB/RJBOuVdtJ5GMYTtu8zOgEP29OeBxTtq0BeSwlCtDi7FRngdUGeGb0mGY6/GAf
q6z1NJK24Ilcs+b0TGw3wSsxdSWHP1AVdU5NbfpQRzjpXzcOxybFB+5X6bpBJZup
IS6JrYJrrSoR05GZwlCINoQLgCWE+zcW/C0GhTcBh76r63e7lEO6uT/CDLQU39oh
S7EnzLVZ5yDr2Coyuhdrl4Yb/iMGlvLJ0hlTIVFCyW3u6gtn0GUwQSoy07Bw9tc2
awYCoZjX1KsoMxAj2gQfErayig4iXD+U/u+0pDEXACHjQcfa3DZqwO64nVklRfS+
AUSyABNcUkDKsZTWWEWPJpVj4hK06fIHiE9qqKfjTOwnTvAJBQr2I3wLn2R4SlbN
V/L4Wqxxy99V+DDNIrfc7NENkFsKXzVImefok+PcjBHVjfujU1m4v9Zksmoa/kme
JSCfV7qW68cA/5eK3C7TUWEDLAFhxlcgjO2BG7/2hWuaF2DjpmS747qOFDcNDj5Q
0L5X3SH5cHWjmgF0dvvYiNs6mUejbQJHqlNEL+0J4GK/LI80/x1GWb/uJ3W5yiXy
2BbnHei0oe/4Z+lytUCjPnPwJemRcfBC8lshT1bNFIZVOdh7439MuLIKymQ/OU8N
s8LoqrFovyWjG6DJg2FkgykVKE4fDH8/nCuAL4Rayx25fPyxPoG/g5fCqokO85m5
b5pQ6thX6rHYFcXqjZkeArLOo73s53RnKYbBiXEltri8RT6kdIBv7ZUVst3HtVWp
K08DEh+t8vseYkwJU0P6B9+h9UgbgH9JmZgC/BVAnV39bxSg0+2AP/gvH0Tfl6Xm
V32v4CcmlhdcL5Wf48ftsBPlifMN9mrcDVDigQ7B+1TXRW6VJfITwYR49sxCxduh
gSIFHJBUyxdMV5/TARp30O5nCLkMThsjBSzX+dPRRUWm25VWvwuia4MEJGGVwi2R
KQV7T7t49FBMkXyz7//PmMGw8t2qr59MtZmu1C8DHVDfPAC/KnZOgh7oIp5t1Pd4
c6K2NwRE47guYivLUKZElzPvZP8QXdHgvDvNCLErrysjgTbqawGfCLuNzh5JfdPU
9NeGhyvkarEWrEw/NcbkVv5TMZZjBYzZAoL0gGHlILtQ+gx+ntiXrDN/0BrgAsjp
1u1LRzGzOWpyo0Y3STET4EYCGW+q2c/qWnJ9N7El0z26gyPnIWz5DT04ZHyXmTc9
KC80+VyuD2qR+12bjCt6Re5Sdmmog6n3AMr2dekkSxIeVKIZQmnckIvROOar14Dg
Q2BmsJ6oJAZf/bd6dJYRTnHL0HuT5x9kg1LJKdGI8WbTpMGwQ0zcnETfpID5PmBv
YAHVSKGznHEHYLD7S9/ltaT/h2ZDg3YAwxunIkhoPPagLZ633KcAy5sY3h8aVBHG
A+V0lBIvj75i//Q/N5JtZ8VmZgJm/ZwxpMU1jvMAPkLPao+6/KiGVUV7tNCgr0NX
Yfdpf5BM6btZmDWjHxRfpm8aag/Lx22CeOAQGBhD8EcfS9HJAG4j/jpOKtPSkzvm
uQUe7M0Hs1grY09wVB8v+WirE/h5ncNh+ihbzMuq92r+imVWZfYc6qbEh4SYjDYx
`protect END_PROTECTED
