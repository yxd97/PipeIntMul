`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cdZR99Yc/0FNMvhj66lrWYAuHJ61isw0AiyJ3W63qVaBRxBgAnR3dMoOQTGJcnMr
PXGf7mbYOeM3o1x8SFAVsdYjBJvCMgTdVW7Xy29qY2wi0FTjQTNb8DZgicRPtEZe
V9KwGTaLYHsUP16yvU4hKGbbg/7yi7uo9/4ucViQs07FbT1DAOtahJ2Sc7d4uNnb
6lnrBjiTdhk+ognNHF/XAfbmICGCS8+PFyiD69+XrxEp3/f6wvOW7U5srpYiryXO
SliJf3Rvu2EgzJccm/HmipRYW/EF2K11kyE6IYViZrLRgD7GlR2gdI1ZsGylKId+
LJr74/s2o+OVf7o+XdQj4jjA2EqByrlKSW+zjR1CWfgN+r7/DAPaHG+d2wqC82NB
e0WyGSOaR3zA7ywYSpaUw125yudDuAt3rxNz1VmOWtvvv04txJRYWvNzbjFJSR3V
Iw4q36dcHB6SwE2zhgJ1AFLoIjO2y4oX5wI7BA4gT/aLPss/TZUlxWNZtEIso6aW
0lr3XWwWWOWO6ZQS8H1YcAJ8SPVFRyxcn5Iv21Uu27rnPOajCcS2Ehu4TEh9tCyO
nNgk6JGm8zv7OB3b3VJskYlJr7ZY7m6mFjieyLlAhEvObDBISDTdqr2EV0tu966H
0p+LwC2OYadXmpOb8Nf2RQ==
`protect END_PROTECTED
