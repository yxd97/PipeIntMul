`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RnNbNZ26pCsN4yMOlXpo9hOjVXIEztiakKmxueORLjDjNEzmGFVlBwB9TXu8A7rp
I9ln31nFyf+S9eJM/ATwHl7MIJxQVa9NySV7xnTpIuXXXlxDa8uZkxNF5UMePkNb
WifmwHg/5KJzMEteEh83XTQRWqG8FkHWpj1aEVxntL44BcMcCK/xjbADnxCW7B4s
Vi7dw0tas+WqSq2lJXuxiqz37UX51HL4Q27OzJ7fZsc8CJw7hORan+zX1Sz8SYY/
GxWusSfV/7hCwMC1F/5No2PelsWMYV+f68NXuk5AV56tc/5Ae1/fpfnlZAsTTXcv
YsXj+EZt16Caejaq3WCttL5rqYVxVZgZdOf4xSe+jlD/OryIuYdfcUlDA/AM4M5e
T+LVcATtdkbJfEpIXs3rTEjrYpYAnYAD+sFLqD8ahFBvf+fPFD1mmliQF7A4Tgmw
epVUj4KcXTTXX2pjoYYWO/HICWvO9djPvEepNzwgANwoEz9tDXoxRK7TM9LUJ8rp
`protect END_PROTECTED
