`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7kHmlW6o92mC3/wP8zF9bpC+Tt0g4B2a4i3xVF/7gH+y/wOrgD2w57GsImzApDg1
55zA2rQeByZbOth25v3li0zpidwyeWXZ/CwKMKlZfxExtmK2MN+BGq5hJsJj+HX+
UUfJhDKgk7UdJaA79XT/WUmGwCSc9pW+98IqfDg09lqD7SwWnfWcQw3qkNUKgweK
96NZfWWZcTVbefdE5pBqFs/uRONZHilrKiMHfI8qwxNbMXvXIy0wUQ+RJSFaSf2C
YGH0tw2/MHw6Kb0zJaBY0j5tfckAd9PjlDtjswo64sejqSzWJAQUWrlXLwwHYiUR
DnqPZd2Gk7g8M+gK2smnKx2RyZTQ2glO4Q6E0E0NQ5I9gZR8mvbRowBfgLqDNFJu
/IQMWyYM5RQSkRLfONAcYaUKHOWLYlC15MfVejpChKiFLISo9bkTijTPCVzdO2ez
29RGgJOb+s9G69uqlLTJnSPCaFKpOh4d9VcEGCrZQdlMyNAVHeBS3Vjh6A8yGkQB
fQQse4hYFukIMGCNm6g8bdj9/RggwtBiafC4G7ynyJevOXEyiEYGRChaH3wK54DZ
mCUaBiyVI8FQDWO/E/Ds4xottGr8TZVr0PEQi/i+n3hdQpS5QOyFbuQU8SZRPRdS
9YgLh3Z8NQVMcngCXMg9msOBRWQgC6V0wuj+C1B4BttVyAz2itfDL+W4TaApe3y/
+20D77rbvvOI7eg7P18KmsPcYXBb5DyLZgiy+Wkvj2LuRNk3JWKcXfnBMVymg4yJ
4yHSM1+HK80wQ8gC/AUNt2r+PHwWQ5o56b8si4qU5srmHucUTGfw9NUbmxD9TGFK
6dT2jYV5FuBStAC7SAJa3AjVFq32+Rx65w0clOATfrxMUMQnEYoWGYODZgkMBqsz
DYpzk++L+fSDUckrEJIB1DvDZhyOGa7/w42u7FPsY9pOaMZS3dwZzCatp0xxbhQx
p++XmpdJFdyWx0SysEs7IIMUaSRD1AyhQf2IR5gAM3uUuN67lvlOt9BE/6t2lyWR
ZWTSWeTziiPetyjQAVs7T8pWKzRmukJllfFfC9Z1nm/KHt784ZhZGPxEJA+QfoKb
Lj4ySwmPMuakGar7P61Zk2li45ljiUvW24F4jOHirAebdokW3PLs8gjQoMv/EEbc
83jpnmXByRRlFVwEglvGzsuA6Sg3IxIcFbmbBk7pAlzP4X7muXh7YsvLgPHq4Reu
TjTfp6PPtgWuvuoY0oz89/KvYUYAhHQNDBM0Y7v9vCLgmRDyN+cp69PPjGBRy/Kn
cKqZUfnKP/g5+A9H5apGYh0HuIO9lX4arvhA8okTpYW3yELphtVDMmj6op9yImth
yhCkqjFmTPwk2kGU4gQsZ6v3h75eITO6KBB6z7bZobOU7zLtMsjFG6juM/0UhTQV
`protect END_PROTECTED
