`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAWfxuICwVEdIXLHu5QwBBHKTBo3y0LivPYfp5v1ue1Ajy/v4HVWug0XZA2tBRER
fBtPPmcwmFQexoX6Anw28g+OSMhlB8nOujRU0EDfuRvwIhXVM5k2fy/defLD43r9
w5QsaSe2uIN3O28BNtZEXZhWZBXphI56x8jJfz69009Ok9Maw5UiS+VECFxIScsh
NKQh2617JaE46ZgNzc9a54FQE9OcfmkKCGmHC1YGW4I0CTEPo6gSKm+ejjKbXz6Y
LMxWu45qTifqgsSUTUVYo3emxkCy+AylzyyrA4jo6nN6Ok6FbJSVC8ygUNES4QJq
5kBnP8oSh3bqhHUOC7/2tA==
`protect END_PROTECTED
