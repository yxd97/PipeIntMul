`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VGSqa4b9OIu4baYPvXS+e60sq0YhlONolTQDFkzW0OdG7jc8/kcwfM1kXcNoMbFj
c8zx9HDDBjKBDalgP5ZPhQnF9oeHyRSfWRAdbl06MJf5mVH0iEVaavsx4vic1+yk
8mgr8c10bAUOQlQc6/hG4F/dpdQHwDl6/ASrEpr/7G7WlhIj+EtllvoXdPc15/DI
LpfvhrMlg1WtIJcwTwwM7w0/tyoignqDmcAoegqaU0zGy+HXKo/nAij0nwQ28bCd
VQFC7yEhTUJoYYsQOzkP5g==
`protect END_PROTECTED
