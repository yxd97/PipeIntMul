`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7peTLG87z1XbL1tQFH9jZJ/LZ/EzQZeQ9njFXuBdM3MIj+NQlKV7jFV97rJaX561
OmtQdq1BNw1ir8bmljV+DmqU8ieDkTHHWkfuseyN5ae6qWizy82WiBX1bChJmu+C
L0NAmNRolxFXhArcmKkuDT7dwAvyVHb4L7xUmPhNAJDvqXaYonWwPLuzbF6/7HRA
7cjc/0jR/CsRt/7zjUaORmx/8ouYlqDRO/2oXWzPRGCik5jNqVbDZQ2sB7npjbPs
7ahvNezra5b/TY44IHJEKkZLNER1W4sK4VtOPluNhjB8nP2yvXYe/ae0K1/BgOuG
ARUojsdX+iqC6Ni96/dEPNLUPKdG4VySdCi0X7XHqmEPj7TovNt+cYpYz6oYH8JU
WLmJDy/Fzol+7wiG1i8prns55vcLroiJ8xy0oa1jolfs+5TsTG/8/cWlWZ/0LwC3
EbcqR8rch7aqX62huVTrWNRBI/sa8WLVta0PLvADeBDQOHVzCgDM6VyY2EUKJkji
I3GkDVWAuYXfPIkB+irYnWmZeKSVF7hT/iVFXTUCn5j0PzrEQVEZ3gUgsNVdsHot
COGKWCidA5tY83tD6IO3bn9CHhWC6Is1iCbMbl1ufjYWgbuLZzX6fyjdCv68KsGC
gq5U37p1D5Mn0TIY8TK/hYqBh1l2Me61165FWwUEpqxRZRT2eyru8rjr2H4plfAU
`protect END_PROTECTED
