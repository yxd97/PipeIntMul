`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b/eUC2ytLf6n4//Zua4fsJT7PpUA1gKNQ2I0BQvF5Ks7TKkG7I4XdVt0zkEPJkDx
g4wynytjOAEXWhkO4h0PLl2BS4q4d2DHXeKfFkKPqVSSsjnxXk8jUaNcNpJ+OudZ
0jF9gw/7Tp88FkHqhbfTZPpwuzePs5wEm/XVxjVnPx3nhDMYxP3h8xlZiYKjfqdY
58sE/zRy7Xmb0UZF+iOptc/iSfC2UXNtxrdsQB76syncwofT5A2e5lZQ+nNRTxfX
mThq3nvxXHS2Zt5iFyQ+/uZUumdSMmhNBPEs+Aas2JNjuTfXKtJsVGtyu6jRCQRG
wRRnVk4IF/KPJMtRMnmwFaWVJ/CN5VHC5TWX1Mk2Z+qGaVWIjYylaq63XlP6FZpV
m1MHG/qG7sHMNbRv9KNwhdwy35k3m75glMmyqrWYhU7owDfELI34tVZNltyFdXz8
NAZRd+/7b6J0x9Bb9VleSw==
`protect END_PROTECTED
