`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aozIiTXDv6tyBGiFG6Dzbcg9ULDFPfZ6uNFfvm7WFZTbu3oDNibM4FHx2/OjXYND
HB9gfxgra0lBp9ak2e3RYMhgifVN3Gy/cqT2ImX8Nr8+pGmGzvPrXOd6GotvZymz
tNeOnOn89xCIvtExrKRF0URu+OXCF1EiEb7a/2qNlauKPR57eK/1GCBWl1duhwId
wLRHde7JZeGaESGywPZK/MsxGamLImKv7ueIrtIv5SEYV7WI9Wgem8A1MibSKjK6
FWti+X2o930ZWxT2Vv5ASWkOOFDGK0MvVGtOE1WxF3ChShAiOj+lXNMNeG+7K/us
5dpyt5Ds6A9xnTT5iPd7VH95Y68ltQ81SNHOn4q6p0s+r7kdKNlOrC0fM+1XCafI
pKtXvyLlrRiHa34zWxh8U6hjRMc23VdCu6dseTtomltq+GrH3zHGeOOA3bsB1vCs
aC28gCoqlZc8t1RZNJbE+UI5ne+JBVRvagfqfai+amYuoh8Q7R03Xa8kars+LYtq
Azy2uSjHt5p1RE2jDPGgTpz4Z5db4zU2DBiN1vziKak=
`protect END_PROTECTED
