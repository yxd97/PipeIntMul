`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iXQeX8f+oqsxBN5qfZQ0hl1/qyDPEyL/4TrCmiI6oDCq+hbrM3gvZ38cszog9DU6
TGhwSr5OM12feQyLWgZqe2L1QM/YAnFKk1JYkUG3yERvpwpG4Hb5JQPz447cLCR+
cblip/o7wWetp8hDthk876k7ddo+QgHBq1wVh56V1xNaFbW7nOrktB12eigA+yNx
BwgTo14SnCN9fsFzSj1jG3vLFW2Ywl1in35u4oyvUj4Q+/AkF5/6v88AaTBNOWjw
it32xOGxuNtLOaK3OPYzDHFpfqMvUxxXhpPHjiRLsOgiZhwcI3eyUKm/fuUBMX0o
54hLJEORDmJI7d/iRcX2HIvVSd5eORLB5k61xxdmlmcfB94CGpD4IGe4rGeiIgbU
1ycQyzUKbS1rgI90VUIwt/3VhyR5xoesZAL+Fm7n8s+ozZq0ot9ixjfjRjOoMnxd
WUvxHLC8qNPxW1tJTjJcQ3JReX7oJDQicRojqw5xcxE+/aWgEJ198G2HnUpSSdJx
BfCqMwhVHePuhhCNfd1XJ2xptKO8bSF6Ghyn6ghk4SDcV4BW9+d9sPh0aLaPcW0O
fn7XDk/3LZOLJb2XWhaKhEMHC2a9DcgItMxFqiycSiB521Y1IRDR0xCBdbQAD6v0
blpS60m1W/1wrG1MfLjA3HNAHsCZTCSgcLlJM96yqy+VVH2mNEy+r6SRVEBU14tw
qZtpju97Lh/ji+rxV+fRwdvpINJfsDqrGjMGPWwmuhUO9zgmVeuo5rc1H8pyuzBw
fJp7G4xeyRvaintuNdoCtg==
`protect END_PROTECTED
