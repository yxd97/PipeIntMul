`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1lggqzsTam+BAALTfKQb2e4vyXnSiWsNbcpOTJRd6l7V65L56kqVRuPSuzRR5rb
5gexn3FHbs0CZjCuXFysXMStdKdTQWGph9xu2qqBBLFWlEmyjkt+gyGa7ZULTQac
Slyd31NviDO9UKTrA3JqfrtT63d7E8yZHgg9nPte1Fsc6UIeWH2RhV+ZiMBQzayY
TqgCZflikvOA5XvE8v48ySIg2zTHhsMwCUiJnIilvCJFIZPca4KyQAws59UQazFe
UTnBMd+1nQ96DqXRv+GjL/CdPQeDiSvx+qtgYzsvNJA=
`protect END_PROTECTED
