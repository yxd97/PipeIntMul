`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sMEnLnPuZOVK8Cacyo7kOj586zDc5Pps5YBo8G3jOtRlWX0QsdB6tcysXljvN85C
CMYKdw1Smsje1NG7JvbMkNXaFW/d6oPq5MeuKx/VC6ZMAc0tpY9aSRyZRHi6+AiM
YebQNIArgwx6i5VWSb6f/L4SZjg51lakeZ++BYeIQLZfx7oNDlhrdMBltdxT9s2I
r8FvIPY7W5gUeg7u2mFNL/zFPXxRVTFdQitZ+F2sjClt+2ZIOQ6hUVDMmfiFmD2y
spOfX8w5BYONWBXaV1Iznw23K4ntujKBVusEUdzjyvao23XcmsOZ2QenNPs0B4xD
oDR88Ii/WDLK9q5JVYLmDrRvZ37jjztyJq9be80z/yLWqt7LAdP4fb2XwEWb38nx
rx16kOzNhgbgv2TDGsQ/p1+cj0oMFsilDjo8bxQ/j8PEETnXdbygnsNqIPwBtL1n
hWMFRDQ5Wf1Y51CCrnCtmiWKlVN7zfLbudUCBiOo6LU9R5VhiF27DYt9O2LFt9IJ
Zh9WihT8DmFVpmGJDCzpkGpA43lrUoUZeWUiS2p3E2iI3Z6/KQlKEfqyOuHIIWxE
vZsvK5UzewYpMQTVhuZHCEwJYsSj2UkVSDmXFRbCdIm5DUstHF/BVJW0r0Wic0pN
lYE7af5FsiPX4B2VZwH1GIUnVpqYfYDSjhEzpz3l6YiCufMoVeDZSqgRGY7xGKY5
sxq5z8xUsVnPNTLsB8Cn14ir/lVMmFEK5rEE5Q8CDLmMV3KuA5TNKbV07jxqTMDo
dtA+eG6xecyvaxeOxyfA/6O8bHQCaO6z5JtJwH761/wAJQqFRQmkb6SHfp6DWicx
fDfamb0rAU0C7/h7o6s2fd3Ekrc0u00qEb0Kpl636091nAGkta2GPech7gNEIf9L
8H2MCvmKgUNFW3a02nk5mJHihHouYNpADzR1r9l2GzBUiM8wdux35n3SdoPvFiQ0
PjMaSze//28/3HUCsGYlP4qNwX9ofb85x3n7A68QfQLKBR7OzBEdKWyIHthFnfX5
u1tjg13cslPt5qEgjQroU7ZR2/5AnBF/viJGjMnlaj5pvtJmPlHuEmUGAUuPPv17
rkA1Lw9QKH5ZW6PVTrQug032ri/xvxHBeEg8gs0u6t9v/9Yh7b8k33zG8fbR5dc9
GtihdOKlVTKhb6cIhe9kHv7tDm55mgT4tl70/JvtT3eVbabYQsapLMOWibDUpGTW
uIdDRwtknRHHPowqBUGtPI3pbqxGC7jD9+35VhuFn5ydXmm3p1pGUKIKOM/iLIwz
BjDTSBkynt+GkiyYBtgVKyAPFGP44Zv+Q7LeHiQNrvBwBAMzzy7CTBny2LFCbEOJ
/TkxXTvVkjR5FaW0LCOYaoJvfVgv7hR37gbCa0lKbhr1+TCSkfdeAU9EFI6moidd
leQiKgx66RfKDkdZF+06GkPBcCwpEknDtoOv2wQcolH7qHc1d1ltY9Ow0E6nYDlu
OBcNmKhvoylDBdjuexnzjvofGapZVyFwLcc5nCypLAvcCxgNqTEXyePoi5twGQj+
Cbj2FAWtNC4szK35VYgcRsEz6kglmqxbrEwsK3eqIeC5W+MrWUjDMYS+zXbfPPFU
uK/UecOx4moZAo7p9zmBNutocMsWSDsT+CFL3iAUVoK3AKxNKmsuUDbY9rho7cih
ByT6oRjrszF7D/QzSfdkyxnynOxpX7lATEeGv/wPVwnxyutif5LdLS9xvB7nE/5r
C3evEiR3C0ZHNFp2UWIhmMvnQfb/rOae5HVCR31Bp7Cl/wMXXd4c+BNrdinu432r
N+Oi21NlU/Xbs0ZVWq6sXAB62V4gXrxrCUxpoToPj/9mJS9xkHW5NQP++DEa7XEb
ilROyBf3W4YLU0cW5p1ZR4u1MKmNJLiELQzsz5qsrfCdA0IjplsP8VwR5Ff8hpWR
+jv5zoo8N0uPkpyqoCdmU7xm7HIaGascGnXen+h5/2W8NCBm2IujhhMvyQvgXYzk
xIQhfESzkjqAa/nF/tjudSsDuFqgaNmzjQLrIpU3stdOOTjPgpmw/1/PgS9gWxnf
KHrUykjrby68Ie3pPkuVTKdUHY50OSfN23dIltn6qBGkVsQVz9RbvA0q9UF+hIc5
+TACEZ4Q6Jlcn2Li2dGKAjAK55gLfN8g9GWeqx6xlB1Rqa25C37Mt+WM0oHuITNN
wpm7qbsZ6WBOmmjCUIDBfTKxpDeYC1mFS2bPpWYidQBVyNoKXVhsWghPX7A+Ls8j
G1lsnnEaNofsqh2boW2EBrz7q9JyMShKUXMdYugNSodC4iRh6HwhpUieZIKj+Wob
D6SODtyxbW26KLzUiypvziRkM5h5GpL+mLAtfQRy5+N0vTzskhqGslGHYfWQ/iNe
ZzDw5Gd4IhObq9aF2T+5AUmrILqb6L0I34/emcUI9DwG2Ad8m/FOm6ozaPMWWcL+
tNc/8ESWRaIO6KJ96d+95m5gejInRjM8CaHKK8o7XiraZ7vKechYa+95hDllXgPp
Eg3xPEx/5Y6JsjHXH892T7kC47C4+88paHXr43Mdy7TchKhCiKkTwI8NkOelqzY4
/JOt7G5Uiwlol81BVsN/STMozYSnVJpo5Wp7r1YyESXw5W3R6pjA7s3Z56fUR3Bk
zkyWhg9eu3UwPIUcsazArxdS+o+qBe4y07h4jwGyWM84QGY5AYHbA3WUehQQZx19
GXU5KKHHLtYqdezH+0nbHBXGN6fkCM9XCFD2I2yIK6if07VObUUKzOGnT4/cPc3/
ge6fZcwpi3HibZ3MN3m/4RAU5HtsiCD0YTVPyE0Mq597etBPM13ZBtauR4Rmmph+
F7fUZn5m+ys0y0hUwGRU9iBP05pIiLkc2LQ1VpEokoMSPxjTDOY2zvQubiLrtG8j
tXEBJokjbcAvFwjbfYdgD1pXqFwTLour7/qxITg+FMJbVrprT2Li5htiQpPZ8MLq
7LWFVgs7kr90Dv8YcRC2rP4VPRKEtt4DE6d0GodkWUcD2ierDhiAVFn5Wk/W3Mt8
ErfOjRfQ3WCnS5JFCiuGrZZ64TC3uXsUKhk8L1FmL5zE5ENcVbj0jcJGH0pCyQuT
YhJX+7pL8TqUBGhhh0w89uPlxlPY52v5HYK9s9Ae+B+Yle/D+7XZ39wfIk0qHfYA
178k4Ep9oa6fSdHjLt3f2tKbfxCjuWmQjK2VdhT/JXkvmoX2K47tl+AGUPjlQsJc
DKVkmLCLYMVK5At2caYFQY/nLucBLUVHGTEVrNa3keYP/umztEBkcSrbZ3SryjqE
mMXBYR9LWRVh3HUwB1CV5r0dpnDwCw917IrrhmZhd9WpsqpkOf62kjFZn7GNy66H
3PX1v0hJw8IfDyobg+DAi7vvBw80Ou8m9G3DOWSk2zVHJ1KuTg2yweq73s4TKKM1
2TtgqAWH//4fAFoGaVZnH09snEAJDFfEK5AbGriigVsTwFbO0v81AF1HO59Mwle9
pbf/i7xfq2yH40NofBnWfWLndr0WIDujHbOagJT4xwe4I4WwojE+G3j/atmPEH4d
93mTdCXvhXojJLrvIe/Y5DTWhJyndg1wtGBzMUkRG1mPL3HHbVKi5V3wR3syNdsV
4LADa0L9Xjj14KwDEEOAi6yn+Bo32SrRNe/kqHE+umkRDlY4X1at2Lk/kji/B2p8
WbR6TqvbruSvL0RxiOOVZAnmUE+7MSAfF1Z8owCHkDa1zRQ+fmNmrTEsJhID+hPp
Z6e+v/EDAbA1NkHxjxfPlK5iEO+w8mvS9z3dQb9HqiKKAV2tZrOy4vFod+5QP13r
La/uaU7Gn4IrNKzysGgndqvEDu0IvRY6rbJuHswvLz7xwW+42yoRtUsp7C2cALW1
VGpt1IaU0+Rjd4oEJiS6PAqagCN6DyZ1vIJIF/7x7Es+DyIPAWsQGdiCBoxc8FxO
Di342kbnwlLxhwhxvDu9b+eK4pjZbis8UONrhurB1tOrr8vgNxgN5rvb5Dv5xtFC
9k5l5MeX+sj8/ab44B9yV92A8FuZn9sII/bB5UEtf8jnDsEaeewXR8CBoeVFumAB
pih85XnS3zdHZWkDmr5wHPL0ro03Vo8kQZqSbWQLxAx92yGLYII54Ei0K2vtBkUB
b/NZ4i6tV+EXdhakt1C5KLNLPb692b3P0MkwshOefBV+1rCHG3tNmf7cxebAre3t
n1nkZSssQrcOjc7Ij4k5IhSAdxWPsTbxLudUJ2qBKzO0N6w+r5RWeBJJq6uefUnv
Rz6sTrSIz+8SQgdbIhqQkBsJpagTBys82vlCI5cnwl5Ie6fv6hpJW76L71zFk1a3
xhmXn9KCfZuNlxXUIL31LWghMjmTA+Vss9oaix5IXC1PzKVpM+Que9y+WHcA9Xj0
8AuPwvO/qRpOGOUc8BkkcUbFSMqzwfIDqgY1GiLzJG8XoJdCvvWACuLs7OtRgcJU
OkvCUZGOr/wkrWOEKA46jzeHfqrnh2bEWcNIsPU4UbON55UnwT57uivC76YhznyQ
DeQSsOvPGidP4ERAEVYTErleqIPdYZgeJOHJujFxLkZ3eo6L2CbXs9pme4ubLn1w
s0iIpUL6/oq+r8QyQvunYi9mUecjWFJhWDP7ae3txi7NaJKpL5SGYot0Dbq8WC3g
0XSg90W4HK7z8krI2CLocAUOPXVfv61uFqwHKuvkGR7GhrIuahYXBhvcVD0SvIAE
CrLfsvZX6zLICewnb8VwxrJfrglPpzIObQE9EZkr5lqjX9L6yYqcvQw9RMKxmvw3
dCkD+fhu0jAgJl7e7kntsgrPWbKU61s8EDhBSu4H/ODZZ3TCdMqP8BEa+w6q8ZjS
VNruKoC/h38nJREZyTBIpiZ1E1nvFM9oZg5mE5Po3MPxnUgpGYeJEqzjLQbG3LWD
o+CRFXqVTiMVAQG3oOKe0TTD+SsJ9UXBSoQjhr1c1rEzhjZVrIqtbn34u7oFmyY7
HP5zdP8TeWl0QG8/3xAquyVWAStKQAGlBXdyOwYNTfirS/cpZAN7nOJLut+mamxX
cM7cgIlOsEdN0zzHMlI6Y8TjPTi07e+bSlO/7P5dOCFzZqChlhzMy7g4nxieJIaF
NHiOk2BZBZFwmVZVh+JyMOu517dcHhJCkhViMlA5aXG6DmgHgIcM3g/j3la//iWF
B7MJZcuJ91apjc9q/UXaBOy0sYj1txkD/2KFuOZNAgkfYwiFm50KPzfPjLwrL0Ir
5/uFwPiyiNdDAZpzKa9UxymzGgQStx3DNFgtzYK89Bj9yk7Zw3xFYoaedv3ic7PI
bLzpDS1VDfZ/b3l2QEn011UJ8bS//F9SdMg581DjCbjpxo2LRRJyGAvOQQK/ADFD
ZcDXe+8DcEPl26JWV/2+F1eA7txVhtEfTsQrOqriUZRO/hli31wAvdowqUF03vw2
DVK5kA0kTxrQ0D6cmtR/R3VWI5+YsVqaRy+3Sz3xgLRE3iGS5xo5y7U4/zwGHEgO
jSKX84l9USXqVIBOY9QBUwE0cx2ANT945n+IZlLz+4zoVXLOKxzGpZV0HynAoOzS
T0uurzJWmUJNws55ga8p/co2gqnEoC9YT3UuEXxCuKB+0hRrpE31tkLcm8M5X6eC
f/NbE+2Ee0ssfY4TM6aVfFFbV0hMpi15F8kg5hj3BMViIJAGkMD9luiXvC5WARjg
BEUhgU+2+pNWLmG3tqjn1LnYaMLEpATOoDgQQk8aJtiJyFgVYQKtqx3jAStIk07W
CJzZehRpx5ScvOm3cv7rb0Phtd8NS5+xm/bCvcB8YlUZ5RqMFq5B+K2qibidVPtO
jBx74/3kePklhmkGgxE9fHXkndpfhj1BF573pThpguSGbp5ORAzOsGR9CgTAu941
jSpOzFGLMCzVbzL2H63fMOBa7ms8QxOT7WALItFe/aRFgKzwc6LqJBXbIv7rPtwp
uednx8I5aHodZre7dVf7pvIVckrznCEhZ1asEy5ikqbFFxg69LiWATyaBkfTBaLZ
YgziR8B6HM6OT/cx34VQJqqh1tYjxdtOvDJCqoWRx6EGgD/bRNthKGe3nya/hgIf
5PxpHrQAHxY1xwAtGdBG0KW1JJgXQ1MC0H0O8WQMEWWCV0CTDEH0XtyZLr48qEDJ
BRlmKVLthZ2eDKZ2lB7Z/nROKblTnDBBklYvItC7HMj/gpaV7T7vZqEIJPjnZpSl
kL9cwy6MFcmRHOnS5yZ8tDb1KQJ0mbLU/3hi4FH3ceR2IcBY9TxjBsA/EmSFcNfZ
7kuYUozoCHu7qoCDEnKT6Sbx5QA7mNmQH8BC9Itwgd07XOjQUjRDdysZfKEB5CzW
jO9lYToOP5Gp2OQ93nv5WPlSdCuzsAqUr2fr95FjTYR0MHe0kXAuIDoAzAgrX3wS
GGk+k5sT0N9yKOU54Jdta4QpTQjHn1RVaWzUEgSeMlCH0NK+5gCA6SIijlkLHwRX
x1tPOcYtZeszEsFWDHj2hJZ8zuJ7EzUyNvRRXTrjCyfBBg0Pf5Xykksq7gW/Qeao
YcowOc7TyBYrcMN1zwYjJvr4WCUErXfCPxUMJdAIR8VapTtjtn74cex5XtT5MVBt
CMKS1lNhZhCILZq3uGqttH3I2kOH++MCLCi4BbZb21A3bV7lihpRy5zIn+gMdCit
6+uKj6MWPW1+m2XPq7rAdTOa2ULSv4f2fJk1xVlzHh7Kkjbw2cv4GWbSFjA0AwIA
ZASEPffVUkGQngEzNEiRsVOeOwfSg+HwGNzLTfcjZ0BcQUZakJ+x6RZDeJd1MQym
GoO1otY9mu00s2LO7SZUAao5p2LKUDBQWbbP9L5sq1yt19zOjvGlbfuI7vXitj+S
wxtdBY9asAmukO9PBQD6LhkM0g+KsGOrSlmPrfhaWHUqpyGd3Q4mGQVB4Uv6QDGv
nOBDox2hCrK/wk0QYFqtJPg4eH2K6pXJGRiD06gYxw9AE7CHoWuMmvKaD3Tg1Qum
ydo0bqJ3ipgX66lyvTG0/27WkAo4CuLNo8Vv5dFoNS5C6PugyZKX4VHj084Dep4Z
3GvkJaG38DZZEmgGUffst8uIIXOMq9yjWJn/WuFJXSDS/qg0I3e8pw/8/GE6pLPU
OX433bgSnCoPVg1SOLsQ63MTMjGrc8RWMINKwy/UdH+uIs7Fh4DXXLiVwLuGKz8k
oexRbtKuuAUo3yAxfuZLLzNaZThwkPkfUQvmtPRTy/r6U7yuIIy30wqc/9fB7CoK
mym6xAh7OtEROnnKMe068exmAVo3eoWRdFqzVnxSJGUjhkwDD3ZXe288f/RV+7kd
R5pfm8mqF6lPKLpkGIdMDiparXDs8WgCkEmsnzdoLhOAhpW/zKku6wGC7opaffZg
McbFm71RJBEc6vFAOK2fZ0JyBd+rM+PvhlF7Do0NjxQ1HuMBTQAvuAQ/uoQA1+oj
Emu5B60UtGI7NlbmGQc3tb5pcdZ4e+wiZwTVp016Wac1esnHqCxJhLeSyjqeFkgh
kpZFXblqbuTEpXyWG5zO+xw597EjDJKhhpb6wmB1rwDc6T9Bx7yuMqyM8sQmPIQU
ayb3StLSSbbVryy48m53AkHtdVAwPrjof9e2V/hww+jQI//oFnkscxLSDqq/VgSY
8C/vs06I5unSrmf+fW8ImFaqLRt6p8FGa8JNNaEN0yarUWb5h+XOT+uR4qoT1yUO
7tDkXWmfgIRZe7IDUzsBMr6eRDLxqCAJix4pOv8nugRMYwUd1amIRaW1Dv31mzxY
qUHCsfqMIA50rQltxqkxYtED64oR/Az3AQNvQq22xFsq5lkUa4U0qjxwsYX9xnqX
Ie6ihLbI+4FZj5QPC5j6jBpo4dKz9AnVj6sIHnkbxsp6uNpcu5IFt4/CqpgwdNIA
sGaXoO1ellWkrckSnu2Xgpuj7jOzfwgRVf1yUNmk/yfxIXcvmwDtlOWva+CDb6Eo
G2X6KyucEjxAQFMVwRosOFmrjb3NYaLd/d5Ahfhqze2zbsEmIYlxNASRSzBHjb0F
g+ewgSNbJK9Sek92oDw+St9MP2b2z2sMXU7mq2n05iM4XyxZBEVQ6g1TgUtdn6B9
gfH7Eudg5RWCfjN05tyLGVDSv8+Xz0WfiShzHEjUzYfAqocMl1eQBNV1yMQhqm4X
QpQONr+J7YjihX9pffHsEIc6XHZtGv7TVGFMkjICkLtv8nYIoEvoq5RyfFJ+dKD9
QU1iu1Ynt3orRTZfXVzLvdKSap+c72TqpDMvjI6y21OTlMHYzIRMhLeFMTBzyZtt
dlj10jYcwezPyUehSUvuMf+RKfg2G/Q7gDkxLTvU9363uYMprRqYuTmnoN7NlC8b
G1Jg8A52r7WCu9y7OlJyjpzpcr+7kT7DxpRhNUr6b/Ki8g9q/iCN5Q36OLdtyeg+
A+pH/wh6qI+2/7NwdzDYqE9fAUbnQ/S1m+FlTjgJOPqDAlOZY5mmAwiJIIkbFHqp
atf2pQQTtLTGCgYzTIX7yat9atnRghRa+oJtrYiDGNw4DY+gPqPkON7KGStMBr2k
wQUUtAyFjgOV+ynchrR7KQbiQQg6XL7Vy2Z7RAxG6rUBarLhFhrOoDNW473xUvKQ
5loaF1FKCABozaMAiNBegYWz67+i5BNUimE6ODOufmnMVr07jiUzxOytm3YzTtj/
r+JotMtKSNaL6flhG3WV9QkC3YBwKeyz7WhXgGP/HaSISutQhLNpnhdn4f/6wont
k2Cv+MMSo8Iw7iJSzCI4YrvfuH7oym/vGkP8lwlDItuP1jhkn2lkdBRMQr86FQ6E
WaEACVv7ASHblPN3UmBJZaupcGt8HY3uWXYzvhZbotHokskGDBBG4JZOWNl1WaYz
VWiqZrl8cW9I9mTo7UaGmdfKuquT2I5Q//VVNnIDCMOkhky2VmDj6KdX5tFBJTV9
RxxZVNgnz4zqOKjIoL58xBKlz7OKVzJZebXTzHkpk5JfiZAxwsB3yuTkk+woxttB
VqG+dyDQJbhlvXgaR+4uU3+g/qyiv8Lt18kyxKeP+kD26vJHxk4q5RxYvirrQCqd
+I4Hea03VM9iTQ7bT2oEsn345PS6CRQeI6ME+mrxjrKKkmIGnMjgIl96usSIngy5
Q3dktF5h2iyMI15/FPByl0csp1roMkAPsxHm6GFdU/yBcu40UROjP6Xr4A6V91eF
6NvB0E+Ulw21sxQ+yUVVWW0INmIIhDXWi36eo3YJiLonwPCpWYLJibsXDZ5Z8LJ3
T+uhHv2e5STv2JnB1OEJTANyrf54IwPK6T5zbk4tUi4VLsN45jDQyqvxIwa/JoHt
RJ186L2Dah6Cia6AJYCFM0nMhHwXOe/5ee2PxHfytB52fc7TXfwoPnL2fF75JPMj
kdxO2dd/HuiATMNGNnA11/I1CaQWmwZu8PrC4QHkfHO4v+RsLPXyONdwH1uW/Xtz
QM1QBoCjjDaWfVlIEuamC0/tXA3F5P5JeXudDyf+3SzN3nawzj9oZRpBwKhMeV4T
8W77PhoRWHjTC7FTvkYIiXAgNK+Kl+QgGawqQu/raAvuJyE7f6M8uwRpX4/TfCsK
hLWKXZ9FzXZBFU1Tf+k5LPjS96LXvX0T5H3Ku36bkigDmHdZ1EeiOk4LMkPHr4qC
rtt+169SlvS2MBpixzRaMKgDwaxx8amC3kmLaAQCQeF3mGE/LYsNZ8uwA1O/k/4y
+DSCl7No32a9FE2+/zGXKqvR8kjoTSvf+j8Fpy43fPgXO70o38+y8neWKdn5XGc/
GedqkjKjqzSmyTRFoEJ6XKTiJRBEWcN2178jJwg1yKDg476RNiHi5ekAkeug0Zyo
0+xjzMb55lug1djvAHXd6+uFzzqmLRovr16/ZRBE4OResMkumLqruukdmAtuG+3A
L+ynaZbNsUcCx1T6TRSSeFndZeJLXJoI9NPWvGq495zJ6ipm8K447UuOwafJNcGT
gRj8IGt4pF+FjmfRLsNwFXZ0ZQ+1AkujnBdGBnsygSn/VEDv3AHSsfWAkpIkY7PE
5lXvROgEI0Vcir+TBtlQD91D1W9LJnhaX1Q7AfvWHe45b23+h+i2oCQrVAFWk8jz
nWmK2Yjp5G8Cjs8lWJLODOT8xEAgmYPoznrSXh980tBNXJn30/sQT3gEW9F0OYkj
047X0l9HhKXbFPwqoEdIm/mvg6mF82WbYW4ZEWd/Bv2kdM3VAjeXvJo+nDwatnBk
JIsuBX5JGgQsz1psQ0JO8gJz9BowsyGQV0XjMg0jDaRW8di5Jihw2ogamjM/QquI
372K2LPUufpdJ94cRNN1orNq6U6ygu6wZxQzX7EL4TG9Bj3hSgBe9j5LrRkgkZHc
vUJ7bXpB/fV79VOOye5Oq3y43U1PHNMAD+0RzGaOG4jQXa+16Gzxv6xvPgb28n65
lHDPK/JmHSLsZJcBivpBodWYkrvIvIH08BPxz0iZ8tOMlQss7jO1L8kLsZujpN9k
NaWwyeL5gfZeHb0gPeTaIb0UiXqpqoS9ADtRt+yVPOhWMjZRJaGN/Jsum6qzi9pp
88rtXkjA9fKED5+i8ueg50LrYYAP8vBRasPQuCTz7+Y+T0InCTk8SvnI434CzU5V
L7VPgb5MR+sYRtfPUE3WHwnNTsfkj+mkhNGE/bAsdHCbvoCjK4c3pDhQzHReWVfx
1PVITbSCBj6ykhZoNKaVpS3oZE/LkKYDwj+2h33m8EC6ODS0UzzV1SCTtiJUN8xQ
bRKcHZsTb2+2TvBbkK39d3KLF8WF8VG3dmqG5V6OtTgQrzANMHGjk7nb+lKpnilP
0akrlt8ueCGvPuhjzVqOO+RiodxGl+nknEa7BP+TXf/YTE3ewtnoEj/7gNvQVzj1
VZGzw6Th5bFSmdZ53pbpZNhuH3OQbQFIGCt7/hlKd11ozbnuT9i0QlWV8MTA3TTW
uszW6IcXln+GMXxuyOvGiUcGAseEVqnCjtQEny/IphPqCmb19r3f0Kt0Pnfgc8nQ
YPJnEzJ4hj5ria8uOGtuSYq/jb0pfxZeEhJKQBwscaLYUUJSFkuZeL3mVbdfg7wP
p++sd6i7GlC4KaMV3g/+6FsrIFwmPRpYMI4g0he23ljMeXfT1wUN4DG9HXPmsSiV
EhJ5RVCXENR7hY2DHPCmr+rCbxOdAzRTcqdB+ZAwWLLx8CkBzyM65EZopySKf5GU
ZOTd/HJ2hBSuPiheA1uJ5vp0UhKvtT+/ZmP+7586CxXJh1MH+LSGxOI3f65pgxBb
301CAJHoJpqpwZBVz5KKOAZyuTXJ/3Kr2goJyXS8326pXh6WgSi6Gd4b4DzxyKdL
qrZD+8JGLsJ8xvOFAzWjCp/0EBXAiug9rmuMoBz4SZAm3UOmVwtcehBcZsZu4y2i
2t+eqDX1m0C/12EfjBez6nVRVShqQIf+vqJdhDKa0Cq1niEbyl8XNqN8hJx0XlcY
SyhJQsnvwTsshDSpVIcEArD+RkKLstyP2SLQqkUjytOSCb3GMO0DVPbe2/sU6HLH
IL0FnIS4Ba+YxlhPtV3u7AJ1JTr1huQCKcsjJiuWlBs/lyp3YfqHvb06o+tDWAwI
hHGEmw68hsoeswCG4FAqM+MBSShRjnIDx6jKlVPbTX6c67osf6HQVcQEB56qk6w4
gfScWEWn1EO+1T/bjoo5ncWoVwxWAzBtbbOaHbQmmAsWfVQHYRpG0QfpfB85mxQ3
NHssD7R37XXKhCopaGk+xiatVichlicDCCFuXHw6K2Sjo76F4pCMxpxmxCpa0+/+
BGtZfUnuZSBZ8iODCROMzkS7SVtY2Dl/QqSIETngUweA8mH+jehXLNYTdTBukDgO
Pa/OAFVlnYoch3r9bNxSDTUCZmCb/wpRxOLXFuLPhjAmozvdnXfFp9ETCGuC8c41
bAOxMJAU8rMiJ0OzZRT5ETIB9SsnuvjQSnUeXqfLO9d3RVknEUzX6uRmyCRUDMYx
iTGxK6WoVVIiJEqSD89DJTfLUC+cXVnSU+d54qYaK7iHe/SOCmPfOoHtB6ZHFhOj
awwIuS7hI/D+2yzH2mL8wm+cHmx00bDIoBKiW0Tu++vVhv3kO8qIHnn1APvZyidj
+NX7BHkBP729CAwuCAIpX4hPJCAX8OGcsX5mp6QELpTi1GUPAuEQ2qRHQKeH9uNH
un0u0eNokbxXvdt0iAhqLoHREByNUO03ZY95B3mYsf6a2CBRhC5ABQgVLeU/xFPc
OMyqJbQWXNEOtdjP/hHDpcAMLtW9RstXqn5dHtUA6SyjOTkTNc3gCZ1FMDek6rOD
ghhUuMPwjZwFRu5Co0Z0BhGDWB1XgnMfuXTcSpjUpF303V83lXsCTlObRw/fNrBd
D3a89o7jA1We/4HVU6DQm6MhQGi9FBdNLKkalKJm09pSHkXsyyyTz7wNmH3XiqP9
OCU84kLpaXOtnci/VCSrmtLROGxWH+4uK7eErtMUBbpSkQ9OE2Rfgk5zt9LfJfUL
8uqauC7xp0KcExi0uNzgWcq0WuiZOLwsNZjuNwoE7xfOVU73rQPrW+URmJKV8d+c
/mfKZ+sf+IQuLwL8cVpyUo+zI/z4Sr0yvx/vEbnWfR1trSwz2t05UIt0s2iflPni
bRtpKOf7eFtsvDD4o3eIi5NaCdYS/6xDMLxh25FYC2kmAnZ+DOoR/OhuhEslUG7w
C+BWs0vdqs2d1asgtExr7osk4IE24ljB4qR6MUTVgdbLUKA+vJeG3pM2z+Dkc4OC
xzrt9QumTdAzMuhN+A72O3qyY+OAHaU7M4twLT+oLvG503Un2OtiBgDI8VocVf07
C6Gz0Oip1v4IyfR0b4/YjPJaUpR9IYkwnaQDswAmfYeVRcctDJK+xzEMW+SbFUbC
CO4zLkX9dZ3nnspIrrQdQ2SW3bpal5frZNguiSJjvJptEGWppTW3UlhPih5w24C5
cQ12Fh7qNHlXmfTtJR58UqLftg6zB3owWUt8sKuDIlnLvmi9YA84uh890KxrBiwx
sOw6wFvBuNv5xijHGfz6gBSLyG1AGfKFKypD6Y1br7pMHBxdZ2+PVlY+Rz4kEFb4
/SW/ibmoakdHbEkRKjh6UP/Urf1etwWeiEtoZ7lYr6VKtDUrx0SNuYDMhnKYN18w
+PPMRB2S0n9ELLSjjnnnzqKQGxsD8QdAGXm5HT4PcV/H37fwfJT7Qy5VNN08RP95
l4LyNNsSlFvahO6lfBPNkm51bxr8g4pywjED+05xcXNLUjcxNum5D+rJB6xJ2KbA
6OnOZzzVUJ7i69hd8ycJHmYQ+vCnzQRqLmTVb5uMoFMO9tfrcBr0bh3YhRQLHLNk
3aoWJsi55zvtjziQ0XLFSB1WkSuKJ4MhDCojwvIFNUasznaMyW4Z0eSZDN+MISt3
aWApDpAiVSw+z8tJgjMR0oqtMiHdQebg3aUVuSjN9lECJ0Yk6Mv1qw6DPLmCpUtk
66YDh4kC24KxFNw8XhDfVBgWRNM0lI8BrqxySnMkIPyN8vLhcuqwMj7n1FicF+j9
SPcSsR0PQMSVac65512dJ9ymXueyPbCp45nOA0AzPsb50jaAhx1WQsnTe9ayANBm
zcu7pIcNJv9RuLYX9z38XNB8rmM7IZjiUMCwr8BOMFZnsrPHScEzIlZhWADiOZo3
V7C47wFZ49taDIz41YBtnamH2PJKtOJHmdViYoqUJ8/yAJIVIEieTWbYjUpcPnFn
K2xCjf1xnUWAhRgp/MUOLyKSYGSfK6x0umbFU3fNXBMergCCT1InQ8XvVyLIornF
Z5T51TBQvviWCaXIMnkSBA==
`protect END_PROTECTED
