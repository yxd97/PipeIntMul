`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DW4vP6EPnlW3WdxgeGpNHuQKlYM4v3rYLsoLmt5u5w3KVZgUg67/KJRRv1L4whOe
70CUPCPFoiz3vjXSibdcpm6jMU2m75ikmKE4reZz8lafq2rmofiNeafIrcSHQxAD
2Khh1JRzEX0KrzNlsH3jQhkKZW9dUQJDHgDseYdg8g9mWVQxdGhY16so+kZgPc9Z
EAGLxnAnR1uswYvli2PB/sqhzwSOFMtKUflPDWt3bqUA/8o96c5nmmFDqbvIjGEn
OPXUK9QhHXw46366SjD1/DLXwMNLLIl50OJXvIrFa+p/UwZdr8GHUhgej1MlC4TB
iMHhof0X38CI2REKBXxHdT+OlnavYLOR2p+v1wPCNbM0yVOZIcITCALTdZuJC0EV
0qPvegbDbMHM5c1GsZcD7KYqe1zeTqDr9N2v51jy3rULB71EYC8dICOioUF9ukWW
yk8SUgBTYAxFtfjj0Vpn9mdmo9Bf6bkjGyH7QywGTyl2t7iMIGltTBSHLjVgng3k
RPTg+w2UFtrH66JIcIFahA1fMY4tY9mbDeAt7tdj8roSWivaGK5ski76oq7JT5fa
K/o1NmDZZyticyYhrxHK+J18JZckaXkaaHi0OoU0E1n8kA/aPDQAy85fPJbQ7Pt4
FQ4e8hx9wAa4NWg2fZ1iA53jlA2Cz4ElRlvqTV1+7p8=
`protect END_PROTECTED
