`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yuMz8Bn5YUrtHRykv8odlz6hanDLpSotY9Ss8KXdSu/gk6fStjxwoPTny4BWcSLm
VSQ0zYa3hMhI8Qk6VJDVCG+sNjPO1H3nSVr9EBbxOsY9czpudZGu+2ZYPs5g1lT7
QtQisuVUKKsBXjm6Ee8j/kRaCsjoTT3BuvqMs0XVjknUz7BUqdTsNQ5xWiw7w1DF
3MbB0EtT1Bk2J5hG2PQQHU1VmDR2/OqNc8Un15PGnS8T0abW65bzfV63uDLU4hZu
AewZW9PQyKR930hrdkgJYeuK5UKq8Gaw8cuTLCM6zJ4nEx9nO7SQ4m6wBeydALXm
RjKGiiR7HkWfJKjBFwY0TVNr/cSJQSQNcqurwxaroBVoNFuRFxEJS43K+2eRnFDs
7tBCuYI4QfzM3v1E7sqJQ+zUeoCYfQEIvkz2cNPs3eRvT6YEZ0MntW7f402YeXng
WfQhNiQURQUW+pRIx57xveqRRAR0KefxqnMdLttEzVxhwc84f5DCIXb2qrx0qEi3
A34eE+IbFug7VrteGxWDynsNIcEVNuG+6/rhGl7HZ+j9zBhrmp1QwPN90iZrS2MD
uzhnt19V4eqeg6UHopsSQWMXTxuNsNlCTibChtZJwaWiPrH14rmd3pS55WtpXmZO
qtpR1jcJFYCXNMjABW75JvvW9vkRWJCzQA3xcOqNVH0dzzKmEp/Ed9uKOqaXrgrS
LMOazKEhIU1uUm+IPycxpuDrK+hDKQAWhF546ppwhiqwbAOuE9GYsyKa9BM2PJHB
0f2/bPGRD/jWOXzFJtCQyPVPLwdEkKcccIowkmSvXX4JtWjoKMfiiZU7CHSCub6Q
Bv3aUDcgq0RftvsNlVhxbin13j/hGiK8twnbqcdlERkbY2uPMKlveHvrtcuUWV+J
FHFEAsNqURIcHCircG+ooQYCvkejgdaPtwQVkEf7cZ/gLnriT+Bkrt4wUDMf3gA8
jfbEBE3H2cGXoYacEByvCevTWjDVanA4yN+cI83nFOtypl1otW8hPUVBHMzJkq0o
ky0ChrfU2e4x0jtDhmF9ckNqZqN2aBZRAUVM3XHwCfhVTX/QX5oWf1++ANuYcdmv
+gERlU+3bQAohXZkIKsxxiH4Oi+ztCVFjDdBDCkb2wFN7Z1ytwWDBCi10HDqw5Xh
WurhORIgFyV3d9T7xgv5SglzklcWXfdHohHUxjYAR401Awelc9eoWEQBhiQoJN/r
fli+lyJj6Ei+i1SS6lQsUdqDASNhcypSxF+tYlCekPjPGsW64hed7JcTmEuFX3QI
NTmQzUv4siIS7HU1vyvkK0iGCJnmWVwjwqwRkjeP7K/OsBhi6AgqVmA/XYJfjd3T
k79ijCKmfTtX10jqjvfFI8O6QrBAgU7C/l4hIU2SOfr65vfLybN6a5HybDHeb6fC
4Rb02pPedsvcJDParrUCc1FqWIDOZ918EY/tB1ZzTaH43aNFwAWpUn3r8m6kjgzM
HOvuKn4rBUBUfBAcWBsUrVBQum6jDHnkNPHhI5ft9x4GGpNkgPglVQULXBBugEre
Q8+hbAeKmg8FAVDAW8pYAchSzl6BC6YttmsJC2yZdzJwVv8cuWGaR2VJkNUHkGG9
fL5YDAIgq9DrRggE3an3HWRDU490euCox7o5lsHZkEcd+99nWuMRWDxNgsX4Uk7+
bp7S2PrB+8d2KyzZms8QOGf6Vb3b7ThXsiVHzhsXQktVaH5pLS6LGf25XMappm4E
OyvgkC49ExmDrML2BkPsWOYA9kLTewLoPKjZqiM2ScnmtHeV7GfBUW/6Y0x/9v36
cXS1ImmDmVzfkx0MVXObewmTMxJ7eiXsDcGey6dO86LmsX8nFpGpkc6mirszC8nM
4gN9n9TZ26gHH3d2ACF4ug+RRLk7cBlY2UpjVpOO0UoRiQXOznqrYDJGk2+g3oUn
zNhLzA54syO2AgySjSGYScUkyrVg231+RVrOHN2WXVbf3/LuULU2ow1/VIhKr0Yc
f/hUFCngwNnppIc30YNFucD+O0O6ny0dfuzCaPHEvyfaLFqfizg0ASbBkg03jr0f
j3y3UtHiW7QzzqUmTJhsouyhoFmslpOmEsssmzg8Ot1HmMAIEaacW7JvuwApvJ59
jg/M3XcT1X4poVCC7FE0yvLk9h0MrPyNRnXJA+PkrfNrncY1whHGWIavMh0ntbd7
b3Y3yzqPYkcRLTgoxorUAlQP2ciolYW3HyhkS445OcFfw1dtD0KoYgyK4AxQMRN1
u0RW3ARlPwWS9d4cu/WZq/ptMf3oW7vjYcvIq/bqtGuQuMzZ3Xsf5Gz3Qzfjp+Ma
UGZuescd+oiYSjyTwIjdU9Yo15ImrAkjqbs+2l0BLoAuwDI/SUjVyJycjnteHL5t
JySJSFrKiAwUjQmN57B1yPL1MDt8XpasbpkgZ7FhysIMBqYHuYdrG3KMIFQc+Pix
SrO248HxM2jEG23O0s/8tfjCtEdjTJudHlYKsNhtaGbANRfn5SSbkImCBvuMnboQ
/+rekHI+JhPBkkxuI/Gs4+1xQHiAXLQwRYDRTGPZqxz4vc9Ws9TCpHEwn20uBr2n
pob+jx3g1sIqmFWc13obHbqQmau8sYlUgWetgdKdXKXufPkjQ+u6LpGDPJ3rD0TH
4+muQSjEd0vn+7Pqrh5hqdOx57LCQLC8JQ0B0B3XQdiGYpJ0dHiDtj7qBuJQGbS0
KhZw1do51QX3DE8bLEbd42H9KaOiz/8pAYMWRIyrboQYNI6T9pITimmXJjYzpuCs
p8cQwjlza8j2o+3fnXCnSm/ZXkqjZqUgBYkOgaEF+5fzYMsPDQhhdLD73UR/6GvJ
LQuDlspgqlRXWMrnvPuuObq4paNaSwIyYW+ihF3smTQDqGqDkCCxFKbDyLyBWH8k
oDebrNT6lhoEqf9fmV4oEUuzhh36GEBgZbqq4/uKHFQe491S6pA76DysPbZrTHVs
YsMfYlstw88pk5PVcR47NsU2b2b14WhqCU0rdfun7oUdr7EFV0hfr438F46ds6oo
Ue2aXVVPAcdoNfT7UGqKgy9ay+c17MKjcAiUX+oy+lVuPTZG+7xzIoSi5GNYygS9
LHmBZDwH9hYSo8ZLZ4jNoFkxj6j31Z3BZcrUB22a+jo4oVbs1tAq0MhX+0JOFwMe
Aa1LkuYqfN3hyeclTTNzfj9XbEtNRPlbS4dZqPdt/YC1GntSygIF15OyfHsRtkDp
HvsmL55dEQibUQiBKeOEuq1wVJMi6tTsxGgmqfdbaNxUp0RK1QMjzaq5KiwreLkX
9JH6JPgKuJ3rma0TRWfE+1xvE0TR2gj4MHY1sjo50cXLpvewXPVqZ+bFf8ac+DmH
LrIJXebcYsYOol0LPCtF+Mw4nFRkh/A/SSDBhEoSnprfW18iBVN17Sr3EBHMR7c2
hk1k5kQwS5aOinb9wYHJlqIQNOavGeY6faLS7qVuKbNyDrAykKKLiYpiqyTtpMkm
5JLo0HQOr8vsfe0rtskPdN7dZntbnrTHHEU1kYjiQFuZsa5o5vIYtGlIseg/5Te8
2aKZt5Tkl4d62FiEtL969IktlLQBLOLGdSMTUWnNtKX1C3pUSJDMQDs2yY3eGWJQ
fYt82pmuKEr4LGXHU0xLbFYsy8UGz7k/VF2hUFIv2vPTNV34NC493qLAnuI8TIlB
P6cuvlXz7kOPo0Te/oexNdtH1Z/mWRt2/aEQCD9mgKnNsxLxWMTaBU5kvJ2Q6Pto
HWBx5AyA9ndZ6v8sZ8lCG5fLySrtCJy+RFWzAMlOQcGO2Jou794tKKpSycAor3lf
MtAJlEs3CAsYGLDV6XHTc/NTuq60ec87nZM6FJjgZBzEM9xYzCt5cawv0qzqmPCT
RrzoaWW16LAziDLhK3A8iE5mVAxtXuKSZu/O9OOvhE4sw35YAgV2qDU4LZSHEEfw
WnYkqEejZ4nfYDjmxfTGBzkQjATIKSwgb7n+1nMcO6rmiafGWKaK6BElWex8+7Gs
xufd/mhb2N6++Ad+YCk3fC3JCEKA7ivec1ar06a53D7sWUgCLN3hNXtzSG72AXPr
Z5REVYwqJ/TVV6u2em2ByvGoj517mfRSXMeSRo4HuoqdwM9cuMNTxnBs1ctqRSrb
cuM1E8uVsTetfMpJYGx5PM2bmzKq80EDhd9LYDwfX7+WjLgHBCfTmjnX+ohVmNhX
kinxMCN6PHBkBevk7pYAhBgEp7NC6rNwCG2Yn7xnLSM1azGntumarGZmAq5muf47
QFFG5347cWIBKsNd9ywie1tIdTNYx/HhrdZ0AYcg6bo5+N3PqL2nD8jLPGzoBwZL
uUdB+wXi29XqnB1WpwdWPz5g/PXWicT01mm9s+MK+xZ2iV8KHIdQD1D9Ed7ST2jc
F89/z9OmVuuClnwIcaP6eRUWsEyF/nVO/d2rUgPzD255b8wKvRjuXsdnteO2mLVX
mV3odBb2ecnnI/7S8LXshQ+Hombmjd7G6AklX6KGj3z4XGWyQMcEUYQWRQo6q5jZ
lCdXYKZf3wkhLXEWrK2alMW0t6mwAi5QzBfL7tjgGtoQZIGbQVlUyo+udCA8moYZ
0dRgZHoyuzZ3zMJKVWD1vmWCwAsCxq8a4DvgIHDy664KN0pDSCkqHR8fEUi7n5D8
tQhnys6YTOT43+TJzJouLD87hpYWvjcViZzG4/j7W7p4tD8evGgCcl+aqe3yl11+
m7L2L87RBtvepkWKXG5AXycVMNbC0VhuwAGXzJ0n/X8Iv52oCkHyLBJF86m3wBYf
JjvyZy/EAuMizB98sb5QsHp0eO/noY8vYu83ep0obI3Gu7vZZ3BR0xVh/ulFtUwg
AlIyEaUGsG8FrggWaCEcNopYTiQ6ikIYtmpktlRlJVrIVrbnOIujJKbnIRH1ojDf
DcFAHBmBfrFu+WIzoq3iPGoQ7b0F7NFrBk+58v6gVi7Vz+WmFE0J9ag+F7Ki8pB1
BTdB+zCbUYV2G+glMDfDnArn+2N5lsByE8LWhNXMfyiKNXzHCHMPByHa9rULFogP
Hzhd81yQrnlNfj2i1Upma9rBhQog+v50EMs9PNRpXCMh0Ojm17BoaHBgdkReSYe+
o7D8fmDS2C9AEeXi1DAgSAICUq2s0vxa6JeLGgj4ZqzurSHb38xZpA3jXzRndWZz
LG9v7+MSv81j8AwVBPI6F6hhjUiGrcJ3mI/rt8wqmx+la3yXEhw8vjD2fkWTFR5+
5B7D1dBTfQQ1F/8mVZDsDDFOTBqNvHNKbQcj3FeGFx9UJeYmJY4Ge2FKZWCL7O4U
DoijJQuLp9BVdPzaMy07L01Rkx+fCXE12N0fjJplYKxZwIsNmjO+dBEHMoyPqfk6
qw7FLZoCJ7Zx8ZKVfeq4Iy7K54Av4q0y4YDWhU2aeAhRwWVhOoL3dMqlES5HnCao
tnzrtwNPp1Rk6fgMVltHTTFg52W+iVmCwWfcJb5ikEq49iIQphC89sMsCmOE16z6
5ANfRehZUMDX+jdPb4QmZSidQWHy7RfA/X5GkKb6aPSwjroNHxEzr1CXZ+8umlRC
95u/8KSvitBenzbEw+lAiruXFJlDoaoeJcD6dskPVs2AzV+O4L37Buzqbk365q/O
g1P4cu5OiQ3uqmGoxSHJmBUhFmf7OHYCd2d9GoKHnuComyJIQj3LOmUMYF+TfUti
KEo5gkgMB8mnK2PLGSCdKiTqiujFo/onlQVeuqovOiRzMdxMs86ojwfDHRjRfW/4
mfVhE2dvgtkFpavRCtB0oXuT1uUk7na7CFmcD9rbov+HHqw2PtkYUT4xdWNhc5yg
4mSs7WC8psh3ty3fM8c/rebEGnaSEefUf27rKGp52o1t7yTsWw3umqNB0WJESJN2
1Yn8uKwNsoXL6bSyQWn1XRKdbeopCoPmTJmh2b3Br6+LEC/RUkMdLgaKMxO3Uu3f
F5watJbpLF4pf9HGGlPzYUkuiHzQFb33gCe27ditG9RR0e+FRBQ0twS8Tv1GveoV
gSrsovrCeWyYqzIdHg6j2HCvuJ9pOFuCopyHSRvYixw6p/XeNC3l43doX5+beRmU
K9lKxs3wb0qhWeh9dFKRwUKU0pgEFDZJHCH1GYm9ky94spkF+bN7n/Ir3KdPs7ST
UmhZh69VUX7bpPBsSb5cvXNV4Vp0CrCs39pD2tERLdMN7gXXEDrquzqskoucfPyQ
RWmfL6hPRluQaCgyhVYABi+Zan8H7RrJMxCJDwflKA58L8guy4FLZ+wagxMwpGdY
UUieeoAXzU1vU7cHKhWFDVDrrlqIIGHz2fF8ZXDq58c91AJB86xzlUKAYFZnujpt
neEcNPUs6NUBWYZRVLH6Tm5ys0AgFFa/NOlAaab7+wGceVfTbgVHbZq5PQxeGPBb
Bk/iySikedDOyPrY9CqHaorr8dUNTCuFYC3lhCWvMBNtwlUuaNz9mHHwpz2EAuk+
4XAzI5E/LGprqdrbrxsbj1Ow7VwWIbSNIenbfKP8Flo9bFKOMPJddztCHJxugLNP
Dakk+eo6tltxHyyL8tYRkHDfefUdMQUYeCq1CsVHSQUn6FxmR3RZA6s/WcXmrTOz
v4hh8mr0FTP9L39UuhvLX8DV62bm/G1WlVIGifuukqNh1HUiqNsY5gGVWVzXUY2H
Ws9J2e5AnhtHkAJp6f754KU2XmoLC0OWXgmtn51yMWxCUDxASUjCBCPKzExFu2Y/
gLXkFgdvRZRlxC4yoo7eKM+FVZ9ErpEcVL5NVV63ArDdz9NwmAT7yO9LQKIwOd9u
mE58pVKwBvtXXRv1L6i9IcLnMks0er18AviSbVaTlGtXE7iG7ed4RZMnWkLMpsQV
IIkJbPC+urJ/nDAxDCFrczE5pxeEoQFElVY+fdBbA5xCZ5nCtfaJx097izmI5bAd
rf5zds936GTb9KjRbQ+p6GZjOViYOryxppI3OzxDcHjgR1hAg9rvTFQNMNnmdnYs
bAFVTWrsi5PrCmdNWyhepAZlfehOihGP9Ag3f0IoJ8D9TUrBtTYLIh0bUEYftMis
GEu3iy92EtJDo9UIfVZtkewp3Ec8wOZzcgUh/Mdr6I98niqbF/gdm1dxM1ClcoLy
LVA9PWSXPj1NYQmcGTzt8n62oA74GrgccEGM9AScVY8/4+dtMpC5lKHjWd07aFpe
KyITrHHcgQ6ArFf0m7y5fXFugPqCcQs6YSduhKY6tjdJYdrM9jIEeYT0hn+ccfsO
cFcTiSVJdIm5Sj9P8ML2/t1DKu58nFu1WExZ4Dtga504R6g28VTirjyS8cFfNBSU
eFC/2G39uAftfxjPOUK5ELKbKdTFCcqxxLu5Hy4hFm/DUeBNPcLbdAtFy62QrkzT
G4XdIhdMPvlz0JTrSXIKqwHjaPhdi0SuvqptJQks3f7PflTKeGw8psWk6eoY7nUf
Ku4rEljhetONqptAjK0YI7jQBhZ1geYioJ+8sam60mOMp7wOQrquURu9KvwicrLY
CSR8722bwoNLDYxkRRdlrtfH1YP8R49hYDfrFCkQOl58Zq70YTOjFD3QfmgTG+24
y5covC66KOsIhAzHnuvrFVjQ3XotmR+eUfAZs5VWZR3IsRmLL3xXEv66s/gIAYJA
KT4dDhKDee7pNAOoMoVakpv9UyrPADe8sZvq1y+eTyix0Qfp/XriCqnc5KsPI33t
1dniPvKjYjQymWJUbZpq13M5TmYZHzAcgys3Pe/bmujtpVzkXrXlKypxvs5gBQys
ZAf6iCRrtGWa6Hkc4IYbKwBaNBfQr/nGJSi6tsha0fUyF6bowB7K0/VlxXrHG+oF
7VDVoYecq7ynEnxs2BqXBsHZC+wL2kB4SSVx83ok3oOZIQuiq5D3q6kXHq5ic2oV
SCuBlIVIxiVKK6JFgqotICGbng9FQ5dLt6mHE3e7nQXmEyIM5or3S5ROiNGRKwOl
flWEgVIYYpcYnFNkZcd9ZBCIzq52JM2FNfYBCIjmXBlywS1uB7nGx7xDdXgJ/H/D
RmljwG2pfpGnDLG1E/DwAvLhA96hAh/EJY5Wr/nj9X1e7z386J0rBCexOSQjZsUT
lumpTC8sj0KIkt5RQ3BTSHdJu5LfLwkf2nVPgv4Wt0+/ZrSLjhGwILOiTB08j2TZ
NiOhgFMRRq5ClRkcfYlZ8cyQdruoCIhsBVdVICslu3vsbXSkxXpUIFN+YLbFs6ZP
UCVwo8iUmgga3fDEAX2fMAXdWddRqUwp5vej5B4IFD/xJYot02Of/fd0FIhKszE0
RPa7332CPdNf09MYOH70mNAKT+ctqdVw/npUbkCxbrSIpgHeTjGJ98Yq1PI6SRaU
CAOmKXI5R3+PvUwbAWVNrnF26/LMOHtVz1oZgdgbGC8FCEP77dqWc/SGM1MpIoYc
Ujc2EVGjjXPnfRHlFZxBXNSH7Srm5jYE7oyxJtiLr/8ZCjqdLOrJHquCCkaxzx0j
FcPyiFu+XxHcjyDpXa/8aoALQh9G7lek6RLfY3efkHAUP7FLEcpRfQHgK0NTPUci
iE32A0EP3A00IpHA5iS2EYy67JvuAOAOXD6o8/PdwwI+5wshBYnBE1UqSmi8lCgT
8ztml918YHovGJ79bb0wFAgV/9rIUmTBxKMBkMpfzEkOpOb9Dt7TiqtD3ajJ1Gph
ACWycGm4IDfyhyZneJgp4JwquJ7G4Mq0pCXe1KgbgCuERs+cA3No1nlJhqgIfUXp
UshVBUArAmBryiQYeq2CRC0oshrdK9+7+5spl0QJ+xLjnCAZQQJ4LtmB6fWQtgAG
M6RUKA2lpLvqVi2Lzk1qxK7xqw2ja6ePZnAiRDB8Uwkm5D6zR16aHvdHsMmB7UMJ
SVM4Ht5zuCX8Ai3cLEAWfNpTrv049T/xoWzVIPEosWPX1U0iZO4NpsKCJ5QcV27v
GfZpiqPAozbQ5XWPQ972hpsMdKlYUwv5orgugo1o57ezLaBJFJHJFRQLLNk34F+P
5j4uqcAfAzfa6vpvvyB9ZwtNtspiwxo1lQfoxaejf/4E6Bc8yvfoHbOy3ZMGjquC
5LdRmgNmeJCSYG/2M2gEFiWiHPcma41IYsrXuUzR7gKEp+RA4nAK/O5lo3YogRBc
b1WfbbrMzM3ySnADljZM8n9knL8CgUp+uiCSuX6QzVmFO+c+vWFTJk4SCO5Ptc97
IaZvXIiDZaUP3tJqRC01WgTyLmO/bDoDLoOFILyq2q0EEVhhtFGtv9LCxlXqyGla
xRfyqXcAOLNmxZ57h+6oz/jT5mrXoqMcAGf7R3NhnmOppWDaPnHxw4gulDeUbSpc
M2NzjR6+ZNv67juJXAmvR7z67FEK9Hmztsse2Rw3i/muPD+2NikOQGvwpvRJq2aw
8LiWduVZBRQTLhqPtLxqS8oeL0Me+9n6yUBj1f02cmPM7FGzoN3JF2UdkjK3eG5/
bCFNag6liWWC+JWAAYdLlRNQts1zZct2IYd/Fg1J7rhkXaUmtg5vxNzfP5jYIIfx
NJlxSt8P95AV9oArbF4fEA6uph+Xjid+/+exowv4YzFEDb3/zch7ANF7sEzKu1kU
8kvQwB9SLe5DP6hv/lqaC2cf/99S+U/tDlCzzmBJ4Pc9D1y2leOErmFVMZWHzjYe
yxgONfzfuhfB6K1EVexARzksIom5WeAEwLCgtBmJotzXeGpShEk1yG/L8kfgN4cY
hZSXFU1aLAmDP88n5GASoFXUfbZ1iy9LiPzkQwtnkkuvwI7SkkDVhb1AIanHxTpW
SirFXub5omm+lcFZ+TVzMt5QironxX/rHi+yblvzdVlSWSPBHPP+vtnDx1ZuzqUV
YbMKbI78A3aPQXFH73uK3X9aDXFMxK5PE47qYIN+/vBNXihVB4KqWLMPsTljYRh1
/IEiMCEITWbwqvtb4aXPcieX8DJEvtjxZ4Lbtp/oT7EYuKMx1QEhUU8FSSEsT6aZ
GFnqx1CvTU1EVSLJHhFq/kmVcU5yWlWkUpAfBaqU3xydvxydqOSttPUQeni8WKWw
GuMV3OoGsMjPhmHHG/UJP71aQGlWFbuismzf5Z7XRiVRAwu2IIRKOu7in8o5HTeY
V4fAdOVYb31gL9h74eKGx1+HM61Z1NubsWqZEqzm7/rErm7w1v/r78cEN3NHS44I
RT2hF5RHmiv1N5UncrT+6jKvTlDsJNkDfyyaaIsSO2RYIUuFbu76A0O1tzrIK4RC
aJ1xFEpnc152rh+G8HIOecXVFPsuGWBUmp5h8l9JcXrl4HCvG03MEMxe2sO9rpee
bYwxGiL+Fmou+pWBisoxONwTOazAA4prIqBkAFjR7/uYxxOubpBzhe/LvD66AYTe
lTC1mPTaNEJ/fqj/c+OVj0dRy/6hHIp9hkv/P0nImQm6/mN7Z/wel4dtqWSsI80V
vo7jaXXUzLlM/zu4bxwppY6vdipKn/Y8NMUQH2ZROno7iRBJWTp9gd13EtR5NNkK
xvw8l0gnfpqSt9av23hh5XgSf9Hku9ZtcXC+5sLslF7RSMVcFAWmrsPCF/+FLaFz
EH8ifiwf46MSIIZNu3+yTkQ8B1ZWJeYryASC/Uma7ARIwoQGJN+paFL0fpDIQI9k
BIIvsB0LQgStlL1IfV/9X1OarJ40PC7hoV2SPBdyHjZYKJLzbhHUc9sBnUHqRbSq
zvad9rapvtUEGkfbNZyVoYTxAWKpi3gHskiAqmL88cCMWU2fl8leJ5M5kSFIJq9C
rJ37Tr591UnrwiKEfegRun2MBxIg85oAJ79f4OIhjzXYiNdeyhmGIJ4sb645/aO0
jJ5dyPZ+5SscaoDKxEWqmmWnOEP1SdxKroNetjOATtpGK19BF3eSnf1isl8bd0kF
3W30mmBuRnO90X+xWlISYmSreRGX3IxncOkD6+UHDVpJxclMXgIbIG+1XhHpvQmZ
dsIHd8NVyyC+dCjN3yZv+rnlJdDxyYZ5HbTS9SC/mOlreNYnRsZxdpU4T5wWmTDW
mH2q52vUPAxuGXoGQkk+D8QFICdNYTIqreksfTiovT9ekwcTBkhcaGFWuLan8B9N
tBJv1B/o3SmbKsG7aQis/OT0gqgHTVo1fi0PY33pmawX0Rh+vV05BEZ7WdC2+b4j
Klsdt6JWJVS4p/ZrZiV0yLUciuga+4jTBL0eIUuR+WpMbivviqyPtMjlOS7NAljR
BJ0vCVgFC42rnJyehX0QrrR+Ayki4KvEHXADTzeKZ4pMBjR+jlTOVyWH9T9puPp5
imCIRAXlqOIhDxLHeUv4Jw32MAnm6tF9ps6Z8eSzn0JEBvsEByNc8SQpdAx8vGAB
2LVpoj1BQHtSycRydg01O7jXeECSqqanGOupiqjHYvS/jgGxopUv82yYKTogOZvo
ZUpGwFn5TJ3KmLBy7RkOrNoAz2pE7Ey7IJUI6W5syCFKYWd+eMGVeffD5AaGQLj+
SzwNUghqEQ3i9ybS9lOgrYNOcvoQb6L+sEsjnRZLkZmgFEJzJ0v1ELGj86VCtzEe
JNuqvRf2nQC3h8AzOU57DCepeIfzXqKAEHH+orINclACo/mbBudGDrKQ+ZjReM7E
Ch9RrDJ3LXFAkmsJvoWnfhWJIEDMwxp23b2+FrN7kKR4L9apdlQ22VdQOK+rjXh3
pf/LZk+VARnEfklKUgXkLTiIikSzV0PEvcOWgi4x3Eqj48UrpBcq48UN1I8LnSDl
ep2pklgwDcPzOIMahc4U+/mlT3YH2fB0TKfxcVdm5jXzSW+EBH9Ho/mNuCaQ/Xma
ab7i4656CbzkI4UNzUlROrct6EMnI2qwi588yi782PKNdhxJHzZvqj5cTE3x1o2+
Cz46bJ1IkzYX82wjKt+LvFubn5nzkSI85Er3DE3MzI4vsB9sfpc1BjWucDLOHtg9
StyzmqZA5WOgHiUI5HxXdUvfEWz6BnKXYepn58WV7o6x79pKV8yZLN/Mn5oBzDg+
pMR4ahL3Ik8T78L62Kezc3GW0H0YYqkWTHhIc/OvFqefLJbxyW6LNF+F24hsevU/
KhoGQ+ArGERpos7bf5EKbdCZSDo+ETuZR6c8HMLJbrxcfr0CNlEYk1/jAN6Uk70D
qevlh/jnHXWFIwT0GHUEm9cTbWjnyDSfyBXSGEuMQVo/WgNoWQOrQyQpROQ7TCU8
zO5qHtGk8OycpB6X3sWbu6Hjne6CiTFSvrTrL091xE0bqk51faHJJ6VCyTap+mxO
/vpz8YDtfK38+H3624Ksd390QULgyv0KMKSZS0XgrGvM4s7aMh2MpjUHvIYmHo02
Qhm6HlSacpECCQLoW5//FhZ/H/XQTQebvZh4HwjOhlQno+4qs/oepi3b/zoXMZNi
npOLU0WyM6WT4E2UZWk72lulp/BbIPP6ZrNrq3W/3kgE/Lqij88CThIxflcITuEi
JA3F4T5hTCrBPoLc79i0uSgyBQb2/+GFWdNzxjsVusxywuzwl0VQ/BvhgOUhKAmA
VrXvbUp5fAXRU+EgkJrX70sQoK4hoRxNj4zxayvhcvkIoT20uv1kqczZm1R0kI62
w2oVNuGFyRhlYMd6J2T797R8lo0YLCiPE5VHSScgOz2o5xggfjx06YFCeulOq/WX
Tr+rxCQhC0Kb/0e01HJxWtcGYP8OvN3QemZo3IXIs3tQFa8p6b7CcYPvydT6Zq/r
IBG9AHwF4mjelgH8bMeJtllWarcAScGdEObdm0tmuzOmx585rtIYwSpz+/64zp7v
NOCjcZViOxFiWhCpSBm6V19XBnh/sg5eAPFjGqEUrQ6LF72Zg/iH4UBFYBAaiPO1
rHD3EmqhRLWfLCQNeszWJAMund4uh4gXz4QplJGj4lNuODVbrCArCTqUnOhx+Mps
DiL14fKgBhrl5S0QritPv4cSYslVZHl0q/T0xSNQOzIw5uhm89RjVpZMfSSgzmMV
FEcR/A/nokZbsi4mQmAjawrMCwVqRAnFfTwIzptJ3K2+xSOYZ+f1UQn9OhUjPFOK
snkB+BqX6N69d67Qi94SUsl7K9rTotnHH6ahywORS9lQbbqyDzV7OjtYftncFFpX
6mJUId6hjdvSoQGWoaC0s57Nn0bKa8Jd27Dt0wrc+cd2fPOSvfLiAYVWZ8cjYAF8
8lni1hObOOBtsjtUQCnUFZvPlUCUrVBm/+p6qn7SKCllBWQ1CGHJ3/cqlD3Cg0XI
al9AFCKyDTCKz+al7rHfFo/YMtzWnVU0s+xeLMh0r6XQ11QDwSIHaDkDeriT9rQU
iTLmVdsZP2NmPJpxrEzCQBwu5cjvrb6+B8d9OGXvOnqYu1P6IrKf4lWNLIo4pJDf
AwQBAkwd02iBastttBjd8xjMXPzmHBX9xCMVBT1UljCbk65djs5gxeD7F+PCccyh
Vib5HvRTpuJq4V4EkHh7mQ3q5Dk01FRXw05oVi54dnCV14NALYkGI8KYEeye2c2I
YqhtjfwDsvVREOyLp1z1zNOI2Aal/B7jVFoK1jHjTdKdTL3otq8/aI5/1jq6sAU+
zxvDG80py21RmIw923HTR6HUiuJT7q432jUKe6gMm0MPnRCnvwOEhSy8DZrxjYU2
KG/l8gAdOsFdWT74GS6VtLlFcutgMk46cZ/PB93ZeKIMrqQYljhnIP2uxe9e7eTk
vGwaWrh5JMRN0O0OSsP4RWHiLrdSdZ4A9TMWn5BVmvGmbITXjsYQki8nDzcEIgsw
LXMuvBKWtmBTWQuneBVUL+20YDPk+KEJUkTBT7HoBZIEVVxE/dRI6+99iAUAuivF
DCp1ie1RO3M2tKrxfYH/49ul44v+ZRQ5No/x12ay2WQcXOWGqHP28LLmg6Mh4gUi
W++Ep1De2Gz2yku9LtuwI/c2fnYZ9IZejhhB2b0CGnrAiwN1aXEaOmdJPQJuUTi9
Hrp0KzzI7o2Db9HF/T/SIaVGvNYkyaimyIcqghH1n+aLP/tfAs878DPDUhg1jAps
7JmnIWgLISjH1GD4lPE+4zgejrdKwqfiatLLG9s8ND3G0W3Y+1JBeYmtNF20EOEz
NVUzlXZPDJXw89uj0A7eys7db/z7bmeKiTDsXkqTYtb6h4yoQOxgUAJNp06cKTvz
ZAdF6/c2SUKW//Bd04Ny0mQN/SjoPccrtrt4A49iR4fRNHBRgcrxy4NBYh8KJWbl
yE4cUvBbl6B+mxWNGBFTQZ3k1PZE1uNKCY0BsdTJR0jNKwewPXVOepRMx/YQH+PB
lReUiNhz3TVYwYz99PG6sBjxBtlqHYsZ3XOEkV1/8zjDyCZKxy406aDFSkRnyXbg
RMAZiCznMlBUPx2/cXDxvjhuI2yzsSzQmMldafcocak7BINbIIJHX8muXpI6fTg4
iBPSKOoyd5jlIxgwj77LFCrEoP6q2PceiRsmU8Q0djUwt+0fR7gmLA4e0fDoXkjR
WXTTsnFrm4f2sjwKoFGfPj2QtnwnSYJWi33TXpurDv/n5DzCz2KNkzX9UEDG+h/I
67/ldAaO43EjIkdKGrZPE1VWrzT++p6l3U8tXqVKvMBSjWfeClCNoXBiIqjmhyl+
gfd/a7rfZ5yUHajCtCf8PxpDGxqWO/tVj5yg2XsQ3zSqnS0iQ5wAloB7mMfCszp1
gStNf7Ol6femkrEhzvw1hdA+mSHIPUVwE48uFWVwJTvbnH89PohNsafACNcaD5+d
2hgUO8palGUNnpsEYjOkyK29RzztfnnYn49EXjKD/auO4LCwsCv89gvz7U0pxCxh
P0DWUjMJsHS3MzOWAwAAEgPL+hOhW2NnKRD6SpCpRehyEJ6NmArcJZ4LiADRZndr
6zG9fWTM6UZQAMg5Y6DZK4FjeMdBiXl/HAkV6TgI0bTotQ8DnmcABYgcN8K3CVL2
DRlGFCzYmOhZCsVaM7ipVoWohbXauUj2oPuQIsrxmZe2HeoD4Xr0dIm9NTmilhjb
OxsewDeVIItRa5M12qJji+6AOnRBSaO3MKWFzi6NiUc2hKk+zONxbCGK5SE/PRbS
vz5FK1vGNua1nSlpsiSAOVeR3xV7cgjnfBKITGM2AEEydxKoy9qV4t7s9AGSQEx/
q2pXfUHRR3KHfti1kmztZZ0yTKbrfOAiYWQ6Z+Due37L+JfveNpyajCXRF2twoUN
9dEH9Z6UvwabQ2kv5qAx9TPBqp+TVNvIZkS8McpsaUBw1TOWO562OFnKpMB4Io8O
CWb8GqkxHWWq78HemOd7H88sMQ2omoPxCexCWqC6XPvqxVzOWGlDgOlZiSiDSvH5
LuBZcsxbdS8om16AYRGaQXdi9/uBE/DjbuWOLBKqq29KS9HhfHpQJS4XuFBuCjIq
3SRRukVG7gLvOUZdvoly8ZgGwndsPWTpy/Hs8yj8gHPKKNqruI9PE7cX9ih8QCND
X44uzX/488k9Sy5vifpMJcMhdNwjB3t28leg+oBfpnx50ar/N1W7gtW8lXvbBfBI
zmSmgkYRfc3vor9JHBo7UdYgKm1yC4H1607qNR60UARmsG/FHw5i4wmZYntF+iq7
IgizdNBBMfbEWrGD6teSaRaa3wkFd3+v+in2WmG+Cjg7eQFo7ZHX3jKp/l0WEHC9
4yebdbQBmduPiqLYHJABkv0Yv5jBGGwpTXfo29KZtsNSE4woBzKHj1oZaST+phT7
adhAmk/nMQenT/seBsYUOtUWCJtUQ6HpI1sIA28oYycyF4ktjXyzbDNDm326xTPi
1VyTvI4hVjaTpsJINZYADcR66tKvplrPKyBXn47TIXxnmvE2O1QpScD7R+sZJ/nf
6+l6PvCysgjQaV2zPeVBAVLWV5rEdekM6lhD1BS2dBc5ojYcqIO3WCUkOnvfd+HC
aw38nyU0opbmTm1hlf9tIxcSJMcOoBS/Bxvk3fo+Q8U1yiP0QcnZlgKJNy+BiLqR
xO0vJA841xutahDljAVFNlcoCr9p4u788KEoMNZDOjHpIaelakHfuhhqUPAMVrLY
y64dZ2jqs1aAUwM23IqomSpp4wAKZT/F0m/1akpesrGZ/gXQ4rABxqb7+HRFf1V6
eRSBrkkAoZ2FDUN/NU54t6zcY0E3xeb2PjmA1k9mb8BatT1KP1XhzQy+tea/rviu
WnDfj/F0Apkgyd/1k6DOeGjChMhw/j3jU9Ma9JXd21+jo5IzqTi824SY/luBmxAs
oIsNxzUakiQTMLbSjYc3x2/EcY7nUct3qKpO4iYiAlBtt48twXwXSsljN2/TG0m4
VbpsbKuZs0VShuMx48d+7NTBlIwG5F+3+DKmqjmPMPuipfRgJ7M1nPp40W4PHOeY
lL3isA0ByEgsRthWWn169QXfMbxNV9AwlLWWzHvDeEHYFHrwxZiF+3/oPZK63zD3
V5lt4XyewEJxa74vdJ/TFnjruwNLEoGi1e9ZbXlmHDl+Fb14AsLRmOfBzGwVUQJ5
9wdaf4Y5r5/OzXmjYlkNbc8m8HtF5OUaU9Z4HtnwFCGrQ4GnqhPxW4V8SvpBBu8t
6c3Yqey/IDM29rZvbcZQfnAKZ+JgYVKdzi1WaLnCTDHnp30WjGfNwoFrNVilt/GE
MQNnRtVvs4PgLFitPqmjOgyrBnpnFT8tUsbgtJg6Jzg52WEedMgzBsfcQTyOpZ65
oPMnYuKXB2MX+MoYVCZQwvwyhmCg05Vk63sD9VnyNSIaXWG6XaD38JSBpIU+xmX0
qNBXxkRLLzVvzDjayQtELLoJM6f3XBGD+rRyy55opRMx19xsOU6uckodN9NxMMwB
WBnoIC4LjayLxZ0mK1YQpNh50jmxoGOVlyfEnrorPKOX1EbGQ/HYc7PLR9nKCyfc
wBhJDKzmKSneoVqh3k9/9TeehmNRiBOha4TakQyWPjVZjtctNOUfAkg2nnVU0JrA
qg8cO5/H6sT8fzF8qpSTeg9p10O8RQNqIgwN6t6EnAQQCEJopOEAFC6pqtINIc5y
mGEuNiHbdRb+w/0iBuLNcsHVdzxd8K30c51qp1JEf+QqeXtXUcHgohGFdaCUYwZG
exmtwNef+TxEIxRQI1MMBq15WbbQoLWjafb9b5qODN79qMfAmhlTicrxjBZLU+SB
eU1+sZrR8Iz9oiX5xahtsJzwY/gX/nNMWZSAAk7ms3q86yDpaHPjq9Xlv2e9YHpT
2wsTqpglxzPegxy7Vp4NtKuapqvuQspuLS+9LKLE/f5FFQKERD+6r6YxDg2ZMm2m
EximP/kfsUxIqwTScNmwWXJF/4cjSHl+2a8VAj1oh/KMM7gxFU5yQI1WQhE8+ZzI
daT3We10p0XDPANnrt8QZbyiu3a5SkOYm/RE4bTYSIQ0hWZeb5qWtkXlk+dHGKPv
laRueAGk4TyEFIrtBp1vZTjtj5YdVodPZ+Bf5eYqgHrIIwPDsN1FiAnfUvMlifv5
JYmbhxBdtQcZhvTr3XYsqt3wfaMHNMituSKXsnBfzxc0BUQuB82zJAvyFJBXPJZ9
Zz1kt89qdZ5TwtUAt1e28IrOdbBJpvSgRdbktjfhvq96nNEo60tVzFIfL55jGzxy
R4rK8kBvoFf9yzMSCBo9PG8+0YtPHO4Vtulmjtfr2DRsW4MyKL9VUeLwGyvEbgSD
1IO85spbiTdPAtYPeae2byd4/aEDouuOHH8JV3l9NCPsSAYm4/AgcOT64pjbWkTl
XT4TXqGaWknMNrLNV/TPa/OOB0ZcQJgO9HR7fcBErDQOk1OxXyia7dE0IZZbYkuB
kLdSDEeanfs/7GyO1ljTtCqIaap/5av730qjK8kvsMBQFUIGEVrO91Emjc6PTiLr
4LgJE5aZufr43EKoaXKPNu1Jqg4YhhGj1Cs+umX3+QmN2Xtsn8DCFL96Ojy9tpaj
eGMff+nvQgICTxpoUo8jJ2NUy5qsUyGmsb4EgDdf4mUqgajk9Sd6IP43MPdAxGa/
cmHEZTfwipK2vCv3znRCgEdKFdd1xkZSQsJcg3UxThKs1KMZDDtODgi4upeUmmvU
7kKHBOrAly5EwY8L82WlpploSOH/juTr+bhQPwEE1dtsCL3xFqtap3QyAy3ZfGqA
u+C6En21LZQb3T4WOSD31WkjKV7JfOH+n1BDDNhgl3u9DOHQVXFyWSpGFJtkNw3A
EHPJtDNd2Xjp59xsO3+L5VtoATR8ET6LcT0CZJe8k+dCbAOotggqmI8Dk0/frDWL
2xB3vZ4abkA4KatO624TXAW827BQU2p4fshYjFSIKeIKohTu9bevTdUJD8qkOv14
kS5tgev/YvBPrDIEcrdANMAV4wrPojR/Nzjuqc9sJCg3B7TwZqhSaGx7EXiYOBYF
yb8oYX2jgL7OjjjFan4cWk4h3KUEmuq0vv9OTIYACOdTjikEQT6ZDw2UadttZQR5
qA9Cz4EUY+vwQS6472QYH7/oi68u9GZXgjhmJzO5uD3fWAoGTBjBhp79v6W9XL6G
biAtWgZEVYSIDVo55r9/xyXb6lGAzISyzA9CB3Vkq69f4NVSnl/TJQfnzTdc5ZLJ
m87w89RupHwt5y+13hZx/w70xYV6h3kmBihh2ylM60dZD8FV9e6G6MZExuS6FM/Q
S86TLHQCu7sqomOf/jYwY9sCT2fNWzDZD4HIQQu1/dq8JmqqAJ961KLWVTFvIlW2
8AB3IV/y+eW70VJSwXljpsncvNFwUf8yJS+FtcD47j1kF7C5JINrufYNLhbVLXxg
Kp/geOysIJ/pwu1qghZLk1iEB35aOUpieSZWP8OAH23y1+P8En31g4XfkxIwNcrH
uOmcUkGSo5ROTTtXyqbx/TD/Q9spGbxauAph20girEJOUDbNvNTkqvijOym7uElJ
2XfhNZ0ElWmfOv33/EbUVmvwiwrg6oMGhU21+Vj+0kW9smoHbtZcj+LQpClm3mwL
+FpnWwINyjXvCpAA3FHmm2/GJiop+JYi+KKNd9JDt8bs7ohUH51MS44ZtpAosfYj
9I3p9SaTlLKupv3DY/W/seLsod7xgYs76f7r4s1710alikgVruYIkT8rZ0sIWVaT
DRoOf3Rp6lmawjg9lcfNM2PhhJ9Kedn8kKizYv9we5vCHZli+lXuFYKsk9fOPohV
dIKaRBxE+4t2exOjOe/emypSBG0sUQU4NF0W/uEoMFlpC54KJJshP4IXKAjJ32WR
E9Nv9OU/HLF6dEkW9Pr9CgELJ+oidWAPYAv07NDJXVYq9AfCfhe8SqvgfO7pWGGk
ljn5xW4BKV5W6qxPa9dq/FTFnEQ8FM7HctSWzv8Psyj16xqGf3gyMSrjwZQkPwU6
mQLJTFX2P7oiHjZ+b4bbY/fVh1qFoVhZRggecinoScENupJCVrcVy+OTWSfFNV7A
zJ+yPfuElYzfNzXy8qiTgPQrdIi5aAbdFmDkY08UPhM4TLC2Dg9QxUtr1qVHU4jB
0twBZB2TW4cJPQ4K4UDAB6jlWOgPhJSYW+GGhJD0eXnfdcx0N/pnro+SEz14qbH/
Ilu2Av4a0gGmgNsMFUl9k68DViAWUbSG6aofNRR1WIrfI8wWopApCBr8eoYJEayZ
reNxt3pfyvMPIOe2VClX0G5scsWYgDZmVm/foCvVvHiDdp381R/95d6LuBaV6DPJ
s5XqqnvLDD3Tu4oenkZfuzUL1clLYy4neUquPhYOdvPw+Bv3RQS2MBx8s70AfL7V
V0ieGNN8Kg/ZF8XnEq20v0KqV217SADxyMpAjrb8xtgza8Y1xv/CRBO19A1TNXxo
MGwcLU626aPCAxKppn0COzv6e0FDRjeeMprnE3wtOj9LbfJCMeup0y/Hr+mSOEUf
+QKL6VjSvq4qYV7MBWqAXtqYKxMxhlO9fLtxesllvMHnwTHyOHjIPvFRBqDowHlW
NvYMovGz+YTqfiilD1Ur9GzLPk9lkyhttleIUOi9IpXLCuE7DehSUJwiB8LstdX3
dot+7SkeJK3PGfeQBVMrIyt784DJts1+06mxE3tjiB0B0RuCKft0+KolHTinKSES
EEsXRTZW5E7krSdZMqC/Iki7Y32dJN6HBx6Lc7zwLCzl1/ZbyxVRuCsNbJeOles7
CKT6EzQlvrpBY6VOwNtZP3dvizEYY8YTUy63G55p6ZMHyzwU80W8HB5LnUr6vPZZ
4tDpSYeNywDzGoCRZsj0BEMMwAADV//TP4rzEx92k3rHkt16DmPGsYgHbRMoq8Ed
iSjgR9GEmkRjS+njFTAE/Fab4LtwM5sne+7AFRIommHR9wS0W54+G5QSzb5v7YFp
Z1bACWuDKfiKTG35xhe3W5yxQEKOBYeoPSG0piGSb5IMANA9/TGc4lRkycTtnuyr
GEn4yUPE9a/WLMZ7H5W587RxbnwnJ9tU6Tcb1xUshN56Yo68ocdokgf4H/1D1JF+
0aP+xId4uxxZAm7wUqitud8Lis7M2ji4aR3xRZ5hU+EAS9rOjUYRKCLRji9D3IFY
AdjsNI+RCJvhY1hU5M+6/zN5qAkilTV66UCzsXrZyRs5rJJudYJzRt3QohOkDClY
6LWU2ePx44Pn781Jph6PbzuU5LQUALrQMg8vtywlIgtIXQ/RepMzxwLdbzuFkUIU
6nq3bjMS2RF3Gf0FZqoXTH7wGxZr2C1/FG4YY+TD4fcq/0b9VEbWujN1eRNPZC7h
d0F/m/U7FDd0sP4W0GkZ14lI4nPjVMNGq9nNRV7YdlPhgBB8XCYc9slt+RYTvyyu
`protect END_PROTECTED
