`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
19CL5D+CdNWb0OUkQNYlW9pwwrTn9uVM942+3OFY081yccZcK2pLU4KxtMLY69q4
ExlwMSWlcT4DvCVrHzepVuTkzBY0jUe2tbrwaW6EM3MAt6XxyEp3aZx4WDP0QtaW
XS/ZU2surWhM4ahPyu3u/39E3vnH5hl8PF1x7sxhKiV26gvgbaqSrn2EPykwFoyP
0WQVxm9k90UTR2MvgNS8SmQa9DQmfLWOPJ2DeJuejVpzwAMtsP+xiq0IObmhPmSV
zLUEbWYyIfpGyGIyUN/xq9BKplTqjv/pHt4sRr/YU1qKYeGHVzO+bvEovu8WV4kA
caCAeUPX4D8veFbRQelHD6KZxCOCuRQPgzZ2qSZpfHojOODnEyr3H8pH8Jngf/GL
8WeG4pwyUgA0XBaYboQ6vlzvbC5Y/0BCliDvoCkIfAQDK9msiCCFiKTtc0K1NuEd
8egHHKLpk65crm6fBb1RZESHrIlGRfv6AwkDtt3faihhEeOfNnb4ckgvgILWhEUB
eqqB+rZX2a73eGZ8LywnnI0JZ2c+saS5EoXDz5M1BgaB+GXnQnPj7E33+hT3Jh4d
tb+0C5aZ5mqRrNJe2ErnTvK8UkCW/GilUP4ssrjg4xhyYpOnOQiCTaaGv6nTwggy
FVF1cYNTj9niuPwC0meLyT/rTMnA27KhFHHuQM2Wc8QHkkGci8EI7pvc9AaM3IVs
4/8Kr59llwMdGbFe15w07hrLwVmH3Lh04bc+z2PpBzrN4JGsAJwSbvDonr2GOQZA
8zsEOyOuuOzreCwc5EMsJ7fMCfU/Gyhz+D95RtFzrfI=
`protect END_PROTECTED
