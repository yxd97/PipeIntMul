`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vXUEMv1nWAJFntOIVYeGOTkyNJKlxmkW1VnuCGApZ7ddVfHkB4kRXQNGxqeuVi8j
sDkl2fI4YtYKQ8UozWDLi1HqOwUUB4m9g7bAg5y1eMgC1yFWw7kGH2Ng8xp5Hmv3
lIZT26kkery0J3ZtId7hXN1MNdw283oovbFlR2xAFoBxv5PDpxChYy4qaMP5Jt6E
T3WmU5XWOSF3/rI7Iw4TTJOU+CaoZPXLLSKwXf1Bs8lPMMLiMXTSPy6vVtgbvbp0
yR0D8JZFBIZ4q6yo8KjwdUPsFPHoD2l/1jFYOqgixpeVAn2KBZ9pNCc4Vb2MXKdG
mzWqSm16sEsw7pTlHMQlUrF7UuWse0UI0FqfWsDa91WucR7x7kS1nKgZ4b219SrY
j0pxRVByy64EPmQo9gNGUImCsuEMmyw3oipLeOyHdQMIcevUOY9ws4RZcNPNjfXd
u6Kv4YhlGg3KWr4VYaO5XmHR62+GqeOIfOIXkC+2waMnRg4eaKdlHTFmqThJjg6v
`protect END_PROTECTED
