`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJOMRf4tTifWazZ1vFUoJ0s4x0Cko2VeX9RwWDGoL5aogFfdyRieC1CN0omRG5MJ
BTi3IPVkhHhvnQBKvGESADek+ZNfrXe8HjBvX+CTR2BUQfo2JH4bhwfYQTZssAti
Bx8+b+gclc8CH7zPUSwRIqYjGFdvsndncsN5nbxPWmiVwsxazixE4RHGCuLV1TtV
6+5SobAgTJm9PWfVQLyC7TrR5MJeAIh4z+/23Xndj05UuihU2ids1CmuKF9DXejB
L3/t4WJarKtafM7EvsGYOJGqhmxojhq3VcnnfMnAgBHdwDa4l3XayEoCwJ2RkpH5
ZyQ+8hJS8cSMepznGV99fRP69r+eRrnxl89c5FyaUdK7CSXqyv/Vn3i27O72To14
r+UZ3/+fo1JZnFJ1tejRF0CSUmaDXIYkd0AmkFVV+xpm8AHakn0x/PsjIP2DsslZ
Fxkxy8lQr6Qattlmc3Gy4z4VaggvXRxhDN1n+O3Od9AqB21skOxekasCNFXMAgXN
vxqJ7YYMYA7igEBFRR1F2wA6qFsFWw1dU7AwU/WpJmTBi6YSc3/Kkid/zfigac+F
kxWGl98tabkYiFez8dyuAWV8zzDN+fPIaczeA8xmOtTEKPikaMhii3xRdMuqiAtR
TwRsRtZCr0RsOjO0h1/u+4rc7cA0hWZIWJw8JHaqc51s5dqiByZPe9WCNhTe0vV/
F+/7Va/7HcFKxfq61pFi5EuDWeUM/g5m57lnLP7++X8=
`protect END_PROTECTED
