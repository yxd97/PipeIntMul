`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vdo0feznmyT9KBZ02PHNwPpRQ6V0JN1lDoj4l+zDY7lyaIW2+FQ5faIK152VKzv8
ePBy3B9KA/8xfyYc11kXHrgfCpr1L0egias2+amJK+o+vCUCVbMNrxjYmtV3VDd0
fqCye1B7/utVfc7r9L3ETWdKC80CZePQfFzNowEpviHVq50AJTukILGQXAKcLS/E
QyD4lkPuas3bypOyS0Nq9e5AHf3QoWWLZ1+CMZvu1MD7C4GKPSlBY1kP5Fhb9ojz
cW/1dd10xic6nc6ElY/OEYWDcKWbNucEaXCSiLw/1555ud5fF0NhcBf6RZEdxNZu
mDTg77epte04dx3tn+sDB7ra7+JbIZscztHET8VRu53BJZ+qqL5iMaCHeyyw4h2c
IhpR7ZAkclQsRELdg9A/NkwWtpklv+lAREZw+qIzuR8z9ls7f2uOLzJPSoGFdQCd
gNDPN1HKEmnXWgNb+fKZDw==
`protect END_PROTECTED
