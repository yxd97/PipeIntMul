`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Mj9G185P3ntmDdZ1js1rzZXnD20EvSFtfw+gVM9mHgjuI5MWfwgEfuHH4Xh2pTo
cPBcM52iVjQRYJ7iOb8FyIVWLeiwf+CfPr+0sMHtbK0Px6KpFaeeeRDMPCLfKjXo
hqNet9JhskF/4aLeFTYNzOG6N3Rz2Mk2IMnOPIm1kulQco2Bz2+PRe/bBnOobnjR
BlfIzQJYFL26JQgKk0wsqmciZBBKPMYRrVguHWcsVOy0aP8LE3pXB29kwOIOxHh8
zEW/r0eTt3wgOCwOxrTndXpWuMFudVBuKmePXL80E1Tz12EPPYkG5cml+0lMjbic
WZJ+IhISG4x2rM7ZbZadk1bLWyVjKY/nsuXFQcmoyFLGU/dMzHbJQ89Oz1SJSDbL
kKaMTL6/p9R7MBc6Ft46XveQBzBBBP3tX2bpb1xaxMUQIpx8NR9fftbQ1XbAH6Tm
R+nDRYOXf5OM3eMebhHUK7OR9pZNbuhK1Z3qEx/nP4eMfIZpeFDLEZA6SA15u7Qx
b999R/Pgkwv97WI/FwjsZcex2EVEoh1CpGrl/F6HJa60dVhH+ZG0Hzb41aqpzPs7
tnbFTEb4pbNLeouisZquamqClCNjlxB//PN41PlKEYoPLfvlugoDQKoDa0uX5rnJ
N+7xN3iJhXVu+HjPnXMCdZaxYWkdRB59MLAcwBsUSx4Dc2m1/QE49L6/8nMlPFok
JXWUxXgis2dGTAjVmUBQLujBp+kiNq/EFpZUb2RfNd/xkpZ8nT+H2Y579aSQRwBF
mTbSgALNDMDHakKywyLELATIpBMmMW45xhH6WFndBinfnVLS0nirCgkCQTBoIYJz
Bylh3WmsmqVbx4gnCECZ0cHfiK+ypJE7SoAeS8Ap+dI11jwnAZJ0c+Ie8aOeNP7V
h82JMJoFoZ9lEi1vrZzDYQ==
`protect END_PROTECTED
