`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+YtIpla6D/53/A+tUwyVC0KRffltiJ7h/7PQc6bn78vSmcii8qxMBz3ohIGapPTX
QzgTSq/fP8fSsTKR1hIaLeQzlVcf166ccRYJhPM1SaPD4un3crSUkHWJFehZ8cmo
W8J1+edduOQzD0VIB+Rm33LWD+rlmzSlbRgHKj6cx1AxL0LPjL+Xc5eoemNBYqFX
qauXUHX1qsUwv0UGbRRXkIXMnWpaLmrR77EeYq85gIfxtitRh5HsEWd6+CZaVk5E
N2dx5oMr1a6ETxLbodnPxLEyBlNpLjwxBgKM1FTdFE+1y8+P11E2WK1gwCl9Su3o
yUD9ZOLl7AAnZaBdF2skMSQOPTf95X0TSm8BWw3+EaHuJeQA6zTfhneuyOupkwyx
3CHnEJHSbaA1475UuGlELrQmPdwo9IqMmSBPg2UjBUqARAAEV79NAk5SFuRFIZrd
p1n6E/wQtRGIiCN1of0b4eEuW3v7Zp2Vo2tknjvSXTZ7JPKYueuofvyXue4GDSlx
xjA/U+ScrJaL5d1ydWQxaR0SOl67e7f4KV/lkKjGdyTlr+CA6nu62OV83UyRaUy4
+6YZ1BvnRBuO2VRdlA7W+++836T9bBVudRkXWkRMhqK2GMLWTxPWB9YAa0RKZpwJ
kKvflGmTn9B2AAXIvHpywJ45nM7gBIBCxEJoE857kRlFdMAq8goQbPCc6s6W/PvF
A0/+wLqCxt9eNPjjHGJJP3CjlQAkvu12nzUxEPIChVjtYor6m6h60QPNq9GHQYfb
JezhFw2hNvTUiaj4QgufPylTt9KcZ4lJN3FWpvebF+mMoetSuEmOvKDoszn2LNsi
0vOrs0E8kj6errWqv6qTRr6mjATr9MDw6IIXt029dfJWvLLWFFApQBVUTTwj+Tzk
TzucTxsfIzzEGQS6eW4Og/K9E784POutcr6WBp5DKZedbr1EpFSFE5gVQfhkSOVr
8gqxm/GPDPtikqehctYcVCA0gXJcS8yvSSUOSrgDTQN3QMiV+bz31ljHAt6yFXTi
`protect END_PROTECTED
