`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TRPfNIywJdK+RrDfgLWnReLMwxQKAz+B0nwAwl+auOKbA9RnzepQcgEGPHT0Nzzf
E7UO+9LGFBIFVwFYza5fF7+i3PWSbaPPIgvL+Ie1n68GZjMLAqGKSCfQMVvBZONw
YMSiB7fdSvnkc3ha3A2A+4n4nkhFph6906Tu+SPaRXNy/hFze26DucfvCV19oCh4
3VP/uV0h23OhmR0dMFBXTt/5SlQ2TW492pnRla0BhgQttXOGU78gpRyzjRvGwnTV
c7qKhtClEtomF2MY4oA61dgK0BnKmZN6O7pEW4iaFi7/cOfddQwCne8oz5jYUS1L
0o2Ggsh+/Bh4eFOoENAf5l+cyrkTl+w4FKs4wiX14FafRVlMjmiAGz3wEvmHpnvH
c6Xmky2FNzWt5lopErsvwtUJLKTt5O9Y8dSUy2OAzRiTb77njEnnOIBLsU4++py0
rJvIUUCjgqu1/EY1nM4IP3/asH7Mklije30rUamVy2Afu/qEE1oiTKh+Vyebr0i4
lPpVVIM06nK6vXgYBBhZxwYE3y7UeGHOhAmYIYIXhJq2ykTAlWgpiRMxMa98ia/t
rQhP812iqH8DT42JFeO2fKVehuHiWkTJf0n7quOxCCQ=
`protect END_PROTECTED
