`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/mTucjL1oI7uQzKkN0DIknGgofPzoVEjvxo+rCrnvFkFvegsGbCFKRezSQtYEWYh
K5m1uPU9qVv4oWHfaLCl1U6UeAQOa8ljSKqoUHOw3PIMzFT52u5IpqZXGvqCKCKG
VeTzjzGWt07dRyusChVmjCQakX5wwhzdCEdLcdX9FmU71u0LHb5MS9NmIu1QC72O
v/1qr6XzbTzAgqp0YDwFfienCIJdJGwFbHNy40oX0uNrZ9ibty4p7Qhs9h9q1gTI
ca7+qSzZtinJF96iSXxtFZqLrKP5hrIMSWiL4phU0zEqfp2KsQnHmU7x1zCXGP86
nagbtI8Wp2ClpTWe8G/JYTqNDsuRtqASdClFpDO4TRMD+skcC8LT6JXU6GEKBfuZ
oGerfHVYUzIYa/GgPU6/fohAV3MjEGtFJLFDHpRS/SlBgFi9CRHnheQF6xjfIQi0
GPesOlDcQlUvhqvmdqe4jSIXEhb7EbpDiw0WIVjC3U7MHcxX8buvTJHkAYs58hB+
vBC1WzxH53WRW5+KBOK7uj5odjlQLOVHjmVGbrrrE/dxWlKGgtFoO/fKuO1xLZas
ENtrsUm/O23Qg7VoC9TrKa6oK4j2S39nqKnqrokBVgY=
`protect END_PROTECTED
