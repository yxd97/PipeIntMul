`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7aEy3/SJr250JuserA4rqjZ6WHPnRe55wAQq+YNJ25iEQQN7NTypHpf0k8eVosMA
KEOjlsg0waWiCEKJgUE2sijSVW2PCtB9mPTw0j36TkbXo+dWdyjcnW4ZCjekfIVw
RB2iRPBSakTINLEddGGLnWOUt77jGnTtimERjpFksR0PGsgow005r5Tdd0WBs/TJ
I98q9681yOgB6oyMClk91YBWHft6MxqwjA0gl74n3GAEpULjtkgtGnLqBbljEHFu
9g91vgMw7ktF2sPnwsNsuBJawmhK/7ZoU2cyicZYdlSXwfUuE6bFJuXE5PpwhVPC
MoszeYa5A0uXDLUsUZMiWouxTd4ASXUsOJ5SCQy2MTKfQjjlnGDkiD9mQoRqUvSv
ElxM9e+ml6UUjMDLeXwq9Vua5hEK07SMg72nN0noYsXgaEtvWoiliAJ9Qr0vB2LA
h6dt8nJARZ4Q3GoTLx4Ctek9CkJdlqczWygVW3lqlnfBhlRK74pUE9+m4iJuBRJe
jMxm/LNJyWC7HRgJAlJFL/MqnjfOfUQ4v44QnSqbx3ej5Dw42i8KPil7TXMybgju
aJx2PEJN2oE32ffQTsEEsg==
`protect END_PROTECTED
