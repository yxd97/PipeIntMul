`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8wMpr+/olLqbeUbhji4V9K6nkT/O55FZbjWCp+w7uCsihqAK70FpvMW2Aws6kuis
hjxbKgUBNBOs1Z+N2YBb+hRa0qlli8U8rf29JDgGwXKrJNbgITtc9g6WV5KFuvVy
y884LpecQ1W+Y+Tt2YIaeOF5OHY5DumafzjZDnw6Y+LxHPG7ojT7gX3I9WJu5S4B
N5/8YB7bQWq+MJJSSr+q2OEk4ZxlGtFKqG7WpklpfLY6HWApXLSRnXa30bYw5UMd
JWhK7l8uIyagMLdfRdlP/CE/gj8alnsIT3+I94ogF23aw7W7AAkZW5lOH4w1B79o
x9qF65cKzFhTNqccpUPakTxvCn6PT/j4CNJYt25Zaej58opMZi7FljbjvAh6G2vf
BOYQ0NtFHyZBSTFHrAAHoo5A/RFhYWtZCcDg/842twhoyZNsFuMmBbNR/rqA8O8b
rMQBjkMD8q5d4lFQoJSfIZnyQmw7h47IFAcUcRziCEMPOGrSk6pw/ek5AlPMuRAO
ohTBXhriY+Cl5qrZKujnqVjbByFoyS4mXpbeckMAuBc=
`protect END_PROTECTED
