`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4SQrer9qtNrgLosCep2r89qMjZgxUg5J4EBhCh2HtH0j00x7IsjhtF2uRIizIzT/
kQdIuXh7A6CpztODsj+lNAIFJOnj6oPkyIaN1Aior/73oQaRtAbeFne/FxmqNod+
cJSNaHmipM8kO0cCE3kvRUEjgxP+I61EzrLiHzc+t5kN0CzXIfGEIddlwWa5ry5U
dN19DNl3lL9gSrgomZ+ot71M5r/+iuVIg4nspQtZhDL/Vd/wNuZnjGdPnMiGqL0m
Wvm8zJpAKrJ5gmn75gHsXiblx/vT9Dgub1676cuFw8qXuclN8ENYmJSuWsnrG7u6
OC9fEs4zdXyOuQqkQsnRaygWPED9CrajjmEWnZVclWfn37krJ+szJ1/JLwPcOTWp
/ir/U37Z7yjbmAIH3ax8aYXABqAEmR6A+swVaVzcdyuoQ6JzDL6vjzvqGyiCu8Qu
CRf0IEtAMWSZ0MTlevW7pP8O40fUlRO4bxtKb+H9t3GKEqW56butxq9VzO7Anat1
f5DJChOgaersr972qDqPRW4WPzLczQ37p20ncS3El0NTG2fvcppAyL+sq1M21CU/
c+QW3Bddud4o2w5RiOjXyL+Y9bVwIlVXaiwQSGtlkM9FTUYPF2HNQymV9Ppq9lMv
anX4FFqA2AgW21F/5YSGLvBdEljMWnOhKV9GemWhaO2AgKgz4mhfEXaEat7b3V7P
WmarDHAt/zGmpvqUSFCiEJ2o6Rn7GECO1wEq8yujV1S//NO/WePvjBBkZz9BbySE
nf4I58iNVIvN5kKyYjLelA==
`protect END_PROTECTED
