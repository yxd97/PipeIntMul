`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MbCfnpSCdIH2AcUX/Ehg/8WuclcOhmY5z/qCzRYx0N3fDajeRIjoUcAskPFPb/p8
B/6Gn5nflUvsun7KqZGf+KSmht8DVmuJGGhDRIrV4zs9z15wUPUHB7Z/zEx2LD8c
JzQrlrxSYKS3YkEGs0YvteHSC5yW6SVAfHa1D8HMoCEw8YO3AYXwrY2lnFAvxtTw
yoA7KrXFcx4njWOrGGAWyzQZkZ8v5gyb/HHuD6Bccyvk5eyvwFs9dTwOrvMIcfqS
z3JxGPdI8w75SSRomEJVmBuH67ABRd8E/U1/yX1TUNMOxyFivITEEx1uvHjBgaLe
`protect END_PROTECTED
