`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8n1dMAeV2VxBzkn9hGI0GWzj9mzO+8/QliCFbV7+b8KqVf6oL1w9Tf4Y8wMX2AgA
KZ4R2DiUw8RRKPKVLK4KY6vX/lZybb3qVbXE6jMGRYUNeb39o3s/BoyJE/6AqEZv
ZLMMwtrOqLIauHmevRu93DtztddVDhdrznd6LxOEDu/XdQkNpj5VUOy87pDnvUPl
vLXIcYfDTRJtuiiLuuH2vENVFoNIDLGz7/gm73nu+JT2cpjA+VSV/cWlLWIG9ruE
O50LyxBOrW+Ha+VyJasI+OxPgmI3Jj0FZpLLBQJbKV0+OZ4gibO39uA9FDxnU0wW
6EO9/AARkB1AAog/yBTV3k/Fn2e5GP5TYy4P7uLzJ67EZsbjGiE/LXmyiJcdZQ0s
CUWQ/VRuw8Rm0mrqsitlp4Wt+gqE4+NkHCpJ2fUhqN7OLnZEW/zQnGN/7B7Yyi9X
jyYc8Ike+cG6n0749yNoWT7YpnRzABOt3U9He1n4BgRsZd84Hw5xprT0bScaaa18
NQXt0nzmz/DZ9pFESsT5etDN0TSOIQ7qUIK3JAigAbJNs8W3SBWMG1qwl34NnAWX
gSJdF2CRKUfN1Og6/FJDw8/xq/GFceiBtJt5ZXVlhjoc0AbXegx09XmzbXone4yu
q4n7vX4U+UeiR9zktQThww==
`protect END_PROTECTED
