`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HWoRaqkSskFhfF4zqd5Lizy9U/oZSO9m5MxfGs47wjZX+dYe+pdYIWHDGENcKNsy
C9I8fXH/tdcCXAJBjCZikRf3KCBCfsil6NdZTYwWXulU69YnZkR8RxNfJOEdtrt8
HhIy/7Cr1729gIXnr8mv/GvGFaIn/FXrPzOVWPDn1kxOgKfk4JZFVG/za37YfJAT
UpiqJVIa6H4XftvBKzBFLDjXRd4UWby81rmFQe7LVY91GirvPD32MDIgyssSQoPt
44DOQauPMhnO0sKjhE0Jnw==
`protect END_PROTECTED
