`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OITlWVAwaY2vO6GEJamj+T35vg417uqPFL6C6ElHpr9MmFP0Rf7onhmuT+OgXlmc
BxoIreIicF0EoLsmEEmBzLTRMoWqFwRSr4QimFq9ymzOhPkVerZspU2QfXzQG0uJ
KGtUOLADby1JsgvShuw1ioLhwANFqSC2mvbCMm765uTimbToxoZlxIlrNDSCaE/y
ciNd6M6a1QgV16+D+hvwVnL6RwS3b3Nd47EgTgcrlI4NpVZoZ2NX5zTNtfLcWJp8
n/LYeLNOe7eshShX2w1BxvZ/nsj4SAy0DEncxCOrA8e8pXabySD7Mh32ZiVl0jYf
58gmGFZqhq2YqebQxjXCxvWlBLoYUeQ3W1vQvNWomgGeKp1+p/MBxmrE6K2p89GQ
sCks0InhUw+XjvxrQLdvFwmvdJsy7DZvcvO4bX97MXZrNraSH3d9DO917RQoUiB3
Fpn1K346/8o9ywtxcT2QmMJKR/VNQAC7ogWcK30ZfTqs2Kge9s7uMrMH5U5KQZ/E
`protect END_PROTECTED
