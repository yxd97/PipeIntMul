`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4aBe0X+8NkoKa97qwUtmScdO4KgrqF4leH2kDkPzZqpZ1E451gQARqtwKT+NZVxf
h+fVQfowj+P70NCMxc0LPcHPWASaZxGDofG/c7rssfztRc8tVulNDuI7fmzepa6h
wj8foWc2WlDV0Kw3qan9U6GqtIyHqB6UwH+ml1zVij8NxcTTAQVX1GzJ4RVHMLKG
mbJq5DTk4ABn/O0nYNdZHuJU5ZTjwCaj7W0IAuBius0neFMxOFeUU5xtErAXwEPH
dqTwMrmeNur1tj2IqPWOYmMX0jh+64FN9/ezhiXmoRyFZW3/UmipKT93kjRvidVZ
A1f7jBPZSmn0PJXboJe9rhUzKOwEJXIXJQibFurxY1brYe0a1RdJ+22nFfh1S2is
xorVvnZHnjs8FBOr51YLa92qqYzJNF7f9Xn1nrwAsz+sZncrVBg4v6hDNfAEZNWt
S0h0S+dZmS5kzPLxzWkhgksJOTRLclzM7ZcTogqWNywjk9j9gI/8IrDA/J9/clVz
lxkvQyMh1wu86pgr8KRAUndZXYT1BmXCl0sEX4D/0+hn848s2OxDCH0B/BSgPtOp
DQIPc9US6fw9XNthC4cDoc+HmEyUHaunotUP+7XzBARvrMJm9BSxG/g+/4rNLxfg
uG9B1kQoYFcdPZrH7WWZmKL25VZJ645ftZQ+Rs/dDOaHogEUdDMXWjpjod5PDcIJ
u/F3MxJrPZA9+RpXFqCLGr8Mzs14BzTk/GfhhJW8QWWOrIu9kk+nJ4rvZYAu69l0
N8fe5rJ7Wm03pfGKs7nwfSai+LUo3dfnmtTpZFLyRrMQqn7oLseuxdAiRF5db2Oi
nVnJLU5gGSAryU3E6PaigZePeCxbOx44efqx8BZMcxZOCPS21uWwQFxwEoZdQk23
OT1MB/cyVEpSkf1NVoVO1ClFjuhzpL64vYiiFKGqUoyb9VP7Nbdw+NFkocyz1FTy
K3ml2cFJtNSjQ7sVFMo0io6i8IP5nBEWIVYKv/N13+q4C7cafINfaFcUBwFEmhj6
z4zuxms8WA8otUMjYdlt8mKO5q7WBxAob3NSpDvBkieHR59NNl926ZnzcYzzrqaC
pwP8J5XtJysHzPfpQwcfysOxvqiFdndo2+iG7pjnlbfzORNE04HrOdWwP6alMy+7
K1AdZmn/G0nSG//WjmAQdwcb9cIFPZaqnfstlrKex2oaEtx2ZBxWVZ9ip5R1ea40
QRtrNSpSMZTlhELTBDmDFxTQHNsX2CkOFxQzEqAD4nkwrcifHF266o04jn59y8yR
aq5469uLfwLAYdFvWrmr8ykv0cfOFvjlIzS3yIm7QN7VR6hqa5q+Wir/kWmZQCVT
1IHsmo5rtTOPGqCVDkSmkPbrYSGDSPHtWSO0mu74PfOqmc1ofEKeEOfJNMEumSNe
XkLEPjPnJdcOPC2depySOTQAUeCblNJiOayggu4+yAdMpZXmqhEIxdjoFDxmyVWy
cCoZ+kLbC1g02R8szw+jvRcjfRPMHkhoS9la2gx0r264KEgqy8P97ffcaJTcGICh
Ee89QaWvIimkClxVuhuRf/GOjR9yJ8511z6iphVa/8w=
`protect END_PROTECTED
