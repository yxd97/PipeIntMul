`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n2G9Yz/DYw7HUEs5iMxmFDM+3NjH4CIHr2Qc/qeDL2detq1Lpu9Dry5THt2Kr50h
AkMW4roLns8bF1YzVoaTqcCag0q5U8/Nu8ON+QyWS2E5MlyrdXGYzRHPoE3WJDkW
VZ8atd1PHtBdEGIve6CV6HPBSWxoupi5v+EDVTPGw5hKZVZaLrrGw/zxk/fg2zB+
esMtINN5jj18y+2CrXXwaqGpuEti7s70VTCgqq+weINWbWAL0+vtO2FY94oyP74E
zsQrYtr5ZNMs5rRIKeVCM+KyoGi4rHc/TlB34FgMNdhbtnBfnnHNf5nlSvuAvfQn
PA/29iV8gESqwSCtd/KExr6xP8i1E3UdwQG4XB7kZ4ey8QFDjk1jooC9CsnDIhQ0
4GCro1oCtt5QeGfIj19WQHK32vqoELgx0fUuq8HxY3l5tLOmfWFTMLP7XBaWFfgg
ZbY6NbQyNLTDYK7nl9Jp4BPlpTSRfcf8OD04pNkcgGWU+PTM8AHaueeqUwojDlLc
0g8qJ8if78K9596e3JAbSMebZ1qy7AZuAvI+87VHBD+ZZZwZiN89AFUdv2smxTBY
0sXmkZbs3eBLAcRNAQ5SSsL97q4ti6Og5YH+LwSe5XrunZtxy4lZz/ICnLXGH7mJ
kKPjiFoFUE1zeC6VfqC4xZPs7w3HGdEFWBNLOsyzeOGVmaRV7zvLvzufqZuCZKi6
Zo/oVoEB3sOk5qBIg221VanWWI4C0IIf0ostnlrHVO9RzOU7zGXVFekqNdPBcoO8
U6IeFb2hMQwoiSI3SwDoaNg1lqPGE3Ngj3xdDDfNC5jPZXuiXB091kFvXifHWPZS
Gzt5p6Qharyzx0hbjQf2Bm6X2l97cQdlmJwaxX+J1cCaFGfVuuauP5VMroE4DLAI
gZXJDMCzLp03iqaR+lfCLikBhqsrFWdCKs5nbQ41FvQzGqg92yLCP0wY3+bztLDz
g8oRQtzil53BftvgXnIOZ+bOr5egPbJBi48Mra0Vdx+QLXd0uFzFuO4UhEw7yi7n
zjNCuavNiWGfMN2Uybor4HQvzlbqDbQb88RlLEUx9lgp86DnaxpHSulGXSpUKIXf
bfF8vxbzHa104o4XKKPvERhMAPjjwUomxDOydu9nT1EAb/V78uc16Ka+S2o5DNJ6
qNDTjASdKsIHdPi4I5EJprLldEeaz/ZIV116xYgckqZBZsmRDmjZaYVu7pe8Kovj
OZFNYTvv/fN2171r73RkiO7b9IcJHE2Zi2tWv9dGLjh0K54K6q60qAU6r0fxymra
QtdVTKMIRoc9nLracK+hCFYK66t3xW8Uyl2AW3TGbdFL0V2FPcIkVFadEdx9puPk
7rPvzuSL92mC+r7Z+Nqr+05HrRPtnxcWuq0Zhog/zEQoep4LeTe0NXXR2emMCYcl
AgDZFiFwD/L9ZF1NvK+NzkNOxRQvrFpeRosaQqOFJbWpsDpg2c/QFLBY8NObvfY/
lnwmz/yRv8uxzZ6hBcdZwmy5qaSPAeStd/uwWtHvL99SNN/zZL96tidEKQE/FmFt
pB3xa3plY4KQUQNP9P+iP+6Dq5DbH30G8Pn6EvbO/H3f3PZEOn7zYTSEGvo7w6tK
4x1BHI34fZpybJP9WZQ5pJMfSxZH90Fj3t7lcfzwNLNdmtkfNq2+Jkyndms9LGs9
WgkgJHXwsLgtUZVRlgnHOg==
`protect END_PROTECTED
