`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
69a7ScFoAomL8rHRouxhn9if6Y6QzapAT0DlC+75X9nChmISQ8mH+Jz/Pfm0KD/3
GOVx2s5TkSSOTNq8SLRN+6Yeklfn99xXnEhX3cfdcc7VzzR4Omzj/mSEKSyG2zcb
FX5vaUpnoJpZduk5M0EjjwWB/lK81r0LjzRAwz4gfTmK6OodUqy5tpjYGR5kvnpS
LWNUKcl82Y73jHAc5j3gt+WJRLX6DLio/FxCzVOtVRXnjkiP0wRNt4QIH8jXHXjy
yWK+zr52mriVJIk5fu54CrAEeXFPY61IVCVseQwjkjBFNFGgwV97BC3UEIJdz5Q2
VH9SuDhzViLCdtZ9ohVQTdhvX7tPI7KC1MEtfILQJ1SQ4wmLD3hVKtbG8c6vqOut
`protect END_PROTECTED
