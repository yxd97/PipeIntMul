`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qvnFkc8uBgOM89EBdKbOHgOXAV2+0gySPXWQOWw6OTpR1ilXq45BIePxsXsUAG8+
dPwMpLf6DGIVywDBTr8FAnU/PskUPhgJiikRZsEfYoUivkS3C8okuApNxDv12DPa
ib8vME/v5LOI/kmbSkjoHq2ztlwPWww7k5x+YecxLCJ+CirdcROMrM3a3gm+EqF4
S6Orq578HyKnwbc5UbEg3iyMeaJ7KP9kyedQ0uDZ08op5zIzvbpD38L4ElIsFoue
+HuKBefBI9p0jxBWOBoOvLMr34nImTJmXcUEG3yP9TKVt64iimQlRtHr7cRKsrVe
FAZAO24lJbkuAfmH7bFjI3wV39hex27XM3YGHn3nbOB6mIdlX4pASmLw1INDMYmZ
e+P1fnB0SkDRm3BUV4KhH78HlovDvf8/dKCAjpezExuvPiCA4OWmmajwf/a4rMnH
ivB8omJxduGMN6o6uXhEaO+09AQjIMCRD+AyAJ5VhXBv/uiV1UfkZuE78Qp53Xoh
oo51op0LLjW5/U0n9m2VlWKJMs/8EtWoy+IzUBoP07hRDDZdz42NIYP0v19N+OBb
5dA2MoPAhaxo0rClQscfl0rKM9PtRJL1zInmpoyYYQbp599romQJoPwa/LCSKr3G
TTu8SLRctVEJ66VrAiY+w8uQfgXeokB0MkWYiIx++rmF60mPWyTEJVofGP7v/v5Q
yNm4QY09dsDUc4wGrdYMxFOIQAVrKQwITZYhWkCI8VF1zH22cQ8tMare349bwcZE
PaqAhwtyi0g6iPwBZVCYWgRQy7SLkInn8TkGOOxWjhSzgp8tzM3gDBI0KmAm0tkK
crwkxUjHZ7WWRh9WWNj7c5OVuZYTCqUr+it+KNHIkMd689AZHoSYNlHA3G587DsC
iT/n2yih53I1vQpmj0alYz8OppSoWwrpwPM8S6bDmeuqP0pri6+NP1VgJwHtLbyL
DQgDICm2mPn6k/IGiyUuosmV0reQT6YaalD5CQVuxz8nHe+sfGTQnl0E1OopigxG
SFORm+iPIkdUTn/r49qx9vn/w77yt8unzjBcBYUSklybuVfMGZEeGa9RGhoF/QI3
xylwbgyE6jqI3eaW4dIW38qI6VGVsGOUphLqTSqeUr6OruPsm+gIqQyhgkQDlOIR
`protect END_PROTECTED
