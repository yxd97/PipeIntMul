`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E/gwIu9p2aco8eFAwkThQ+Uznh42/L7KRECNIkq9437tyGdSwfyFdf4KLRvvLhhG
xk4Omh0by7pTIn1VfAIiSbEp+6Vs6ZWqO+jzQPx6kTabE7Mqk/piiLR80SZKl1h9
571fRo7HuiaHdbP2KOJfzhIoMhw9h9UzJsoy4bghsot4EMa9JGdhN4P6i1nimAMT
FQ/xNUJRkL0EWVwQcWelQeVP6L+lOOfb9lruIz3+LqRQpgSIy33bSZRXnXHQNhLT
mBZ56L2qVYrFsS2LF6hcT7XoappIE/YiARQcD6OMX24MXSxLIB9QA8BsvfbtETxM
POj+PUQBQCu3vCZ+F7zYHI2Q+lpaVVJFmeQnXoSVtt780nKkncsO15B+tKKlFZ6A
1DP4kVmuU5Qa+K9ebcwVPA==
`protect END_PROTECTED
