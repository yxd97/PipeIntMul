`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pk7k85ce4gXPTicIvX77wNz5DObkQM1UB9LhppR55z+ddnvBZIc0VV09oocyWPpZ
CItDz20oumlt2js6o+BmXEDRf/yv4QFJ3F2y+Tb0xPWlhuw1FEpc3F1oXmmHlrU+
mJScjX0MVwnOGRfPvEAjH3BFTtmfJRYUljWB/ZsefYJuQWwOdj306aDtEfELxndT
3Cc0cOe6Ol+bmnDeAsDWqd6J92XOoJtPemWvFw/+oPVkB+dwL0/+aNeK2ET735WA
zXs2TV1uYkAPhjYkG2dnMP4HHhKIOZNXq1WQTRpE//TBTRAwNrzgeq9MezHL5mAF
gBNoU+Kh4qCRxWIu2yIqaYdQA0voAHu7firtP/nqOWEjv2GhEYdXEJeuE0nJMOoC
OrHEvd0LaKWpUx5f4LaZRe7eN+gQw+Uc6p5zh6v4eJQF95CFsJKLRcszJXr9ctyz
ZxUa3otdcP0/dhvOwNip3TGDPpUWUnmDBbf+fwjjSLQ=
`protect END_PROTECTED
