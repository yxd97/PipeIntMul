`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
INgSOnyflqJgTBoND7xA9tptzQQu7TPMyUHstezPh7PK0FglQOK2+0WmNw7KVVit
x2Ogh7EzJRVa37jejru0lof84tz+FuD7VgD9QcRtEW4oRkA+y8RYxZ0k5gUoVXyK
krAJo4v8wZxgU1ldRG0Zcu1BjVVuJPRoK0og9TNiPfqLX5hEmNpDAn1u6t0xVXEm
/YRs/BkMGoTMejZdpd48wv7obzjbcJTzXdPpbt79IP2b9OkLHfmKYYIjhm4hRQJ3
xJNvSaOPOV7R6XF1y8UKOF4kEdwQym7Jl/yxZn3d7ZSGTHbCa7+jIURHhNBoEv8c
`protect END_PROTECTED
