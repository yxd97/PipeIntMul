`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TiNKp0iHRuEoyiDyC0J1ggPA1LaqjqhPiV/o+aN8S4WlcB5BmPyxVKZxMV5jvtUk
fdpYmSRDN1OZLJU1TSn6roXAXBA2PB4E6ioBbQLj9tI5vJdPnQ9YVUUTvHlYkQNL
+NFrBxeRZR7bZqJr1yPeBSwrRhckJwNTjJOo4xuaHW8u8eRypx+a/pCagMzbLj4/
lYZJX3CB2akMyOyuPW+O+fd0YqPm34AOrOkZXB6+/OhBOxhjhqgEB+j972Jt8EmE
d6ZrY9xfb+AV8vFMYmfjOAI9LXqw0m20T+WVIbDnR+kYYsqlBeORlYnX/nQcwt9s
XBE7YSv3vCOx/3Nt3XIzEzHncpvC3ZfFR2wVYzCQHoKb0ZBbzlLlcFpx/O8HYZ/w
GixO4MJowXw2chVgGxdS4o/D71xSeG3F3vlFooiz+RgBug7DCLEfULF8ZXF/0yIU
flqWfwPmsPUDJpLdQwngYX/hjfMAfSAp9KU5rRZdo7wpJs6OiGR/GD2YsG5v7As5
+DAX8uEPKuOTMv/Zf52Wb4AlB6x7tWawY9RsP/8BRBiQT9eqDNKZSaiQo+2NeJdO
`protect END_PROTECTED
