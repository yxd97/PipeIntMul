`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O5AnQmW7rL77kvXb2EKQEoZViIHOopgBFcuQwKHNfYhsw+Um/4Z6CwoIZfihm/Mu
7n3wqQIKeqLNhbpn3hDb0pZGecvil/aW4ug689S4Uipynb+bQNQpqcitwk7IENns
gnJLnW0bIaVyQxKuinrQXQ==
`protect END_PROTECTED
