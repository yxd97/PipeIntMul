`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ig73XpyjL9+6Q+sjyiUk26/peEULf0zXdO1Fu7IWhz04aL6cNVXz0Y4rI1tJfORj
7a0UpCGGFvhDp/dlzh+mrd6EgAwmDXnyEDk00ihbhzmaiUWeLm9xs5zsnKkRn6Uv
fAPu34R+wcQBaumW00kpum/eAWH6/SkBILXXBiHMzQUezqkYoLno8CXCw1C1kas4
xAQtcfkvH4E2y+UE97EnxSA21+jCeRUdaTt4PfsSmwAXyWawcMt1+cLu9ft98xQH
/qnB01K2zmQFRjgWiocOCTVI3t2Nh75OLBwWXKIncTydhkWHrS6DE4a2KFfE6jPE
MKe1Qy55hYOTp+lYz9TW/uyYdlzkKXI2nxErB3587h5aEo/Ikb4znrWpNn6s7nGn
yMFLUyiQBFo36A4yiXorQUb+ay/6gsTtTwQDb1cBgF3uQ21+XX3NqdStE0pt+ZAD
mXeZgPN6yAfjRx4fZQL+vmBnlSQMX8e7CCtZ42wBh+l680qYngad8Ozby1XduIbE
3KeVK5FqTfLM6y/eDx+9P3JMTjPUcd+nltbdMhFTS3PENesvBj2PLNCeuii3V8V4
vY/Y0U8tf9Fn7VJqmlFxcEEJYO0wRAWuDkRNKtUgkFd8XeZBfjsJ9LOut6DIaSgj
8jT08ro4h+HhNlWAEOK6G/DgOvJmz547aXfdljZndJKk4cVY174o0HjGNligH5kJ
qyztqLEnK2Fh/4KHDEQy/HAqG4iK4qZ0SqDeucmK8ix3jETa77YOXPTU2LLEBqNR
JwO/CfK0Dcai/cnitlcKsPn62QSs7Wz3QnffnlqTcEZYPtgG7bhJW0cV5mBVbFaB
irXrgvYQCxJ/xtcxy0wULAKqNXY5HuqS0ek9NWu1u9tIeFhGuZFewFe8RjJtJHHi
Ap9Xp3koJmxaUtgLIR6ozwwKZTxZsWIF06vTOk4Ok7TeWPu8wBKJain6kQ6/Gd9b
3sR2qSU3VU++Rhn6vSxU+7F+sVZj1fXoiNUz9J60rNkBFrXyLNCX5YuELCLV/RNx
zSGtwO/nEwARkSpaApjusXDv7YjGzMkooom9DYHmHjrciX22cn26ThV51SmAmZQD
WvKRBppQh3xjlx1RX+Azqn/PPh6kVb7p6r1/atOaPBYbpZRf4Jxb/8EGTx55bHgI
xGk4hE4lfn52g6KskCBJ/zMNPCGb/mTK6GuI6d1M0/Slfr3TxpnzjcFECocXPxvm
BpvJ/P6eWW3lnfzDfWUUGz68V7zHnWJ6fIUl6iBpV7KbDSls56r39i/umxAA4H6z
immm8urfVfJohVsvkaWqs9nw6STClu241mxCAOxAEwezDxwrVFGIIJDG5HMtP0G4
x3fX/sBVsKxUpMoHqsy4xjLvSWhPplgUw3FFBpae9Nm2J2ZysQvoB827MXKFSMVO
m9Z9wKBmXcKGdIfZS7n9OA9WnVf084TEne6FHBawsmFyhrjF86SIBO3Sm04gYtl1
eM4Hm8ZbmPqsEoJMmwofQkMghfYucGSUF37CxcnXsH4whC4sXkdx8jcJH1h6hZUW
5Ozf2nT4vL6mq3YLVvqeCRx83eTuQr4MkxZwXjGDM01SNVZ/PChsiP1yB8rcH3eq
PWz60oAb0yPnxm7KqgkL7SBP4sOMOqU9sKcehbYwM+jmjJRhLPIpXWV4ce9qXXFv
57hzFxI7KJgZUrCrxaE1lT1F+miTe1SHZY4E3U493IT6vARgwUxQKB+i2i+vEWMo
ryog98T6NzuT9iknXnQjJihvUhFu4C3cl/JmJOsH2X8IIZpRAlANcLKnD6lAPHKo
zW29J4z7Nu28TugPu3MIZq/2FEHp6ZtoHL6ROGRzHVnI4Db5QtbX9V/p1cMFkFLe
`protect END_PROTECTED
