`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hIGUuJkzUr9kiQfGWSSx4Hz3TH/J+0XeGX9SoVbkUkAw43aPRbR5nDdNLdFrqNcE
I49jz41cdLcKoU/KwfcSevSwvLICUlHIUeb7aydj11GHO+J70sqI59gQhHr1WvOq
FLyI0/+T6tvyF7z8lX6mqWt8eSli2i9M9/zG21P90kaqwX6vDU8Z1+UfM0h6LtM3
nPtDSlwa7co89ExBbweus3/FMCrE06ntn6RcTP+WX3MVDDwzjQlmqVk8k+73Ipfa
PcrvJpWkVy7CcAdTCK6rs4cH/XRNeDPtXFSyFjk8mrFBchtKQcwwsWgoeEL6z8YK
SYNxcVFZzGEujo0TuNgCn32YAmoGBhwKKWwpdxgDdVuaRKXXn7J8IS/qwVQ23fzK
RbzRT69PUkJtJ9s13pjg8Ujkv8WZCMvOO3AtZ1PoVh0zTXjpCyR7jDyb389pRtG1
JCJfVWmrEx40Qe3G2eFcGFDK+rQlkLGCHrFFiLpydunm0PXcQ7Tb6U103f2qmNDx
2/nJyQc22H6EjRjyTjFaea9xaBrSMToi1zL74WV3PZnv0pWoy7lcrQhM08McEDCp
`protect END_PROTECTED
