`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kA03FY+RCdRszflQsRsVWVzN3gAkKQPdSiEyX+GnyO3BjNz8CmptMWChSztWp2Cl
uBffbG0nbwfyprYiThmtfjr4F+x81mY/5pVU5oXqa8WCjCjbrF06/jYSBECPTFhf
cB4mbHI9HrO0obt3N5J32GQ5Izt4bSHulmG8ReNFqTxWoGjoYYM4uAiHRiXoijHB
DF6swDrTxt+vpjhRcaC4tGyIBKlTh/9pcy79SFsZPnOD/wHFy0rmzzpTGieI8VRn
5jqIu6MlJA2qfz0LniSi/G8fd/iCFNub5Xho/tq41YCXgIuXID3XSyIjB6stWP6A
MgFGTFabDGiJ+JMTciwHkVPYf+3A6VPHlFC2dy460O0K+SeiMMU70lBdqhEiwy7v
IgTAQhC2q9Ha+wuT03LnwTPh1nkQvOWXuPnO57+6rbu+Stz5hatVk1hNJggwIQ3G
iFgVy+71IL+AWQEAkSgMioFKyqJDI+a9ecP60lhp7IUbkhdvuIYk+4mBHxj7wr/J
iWRJ44NCr0ntXatBZ6OMG343r02Tt+xXx917xy0mnTPj4YGjaWwPZNx36g6Ix3C4
/l+hoy6r9BzT4XEwrh7fmPMeQzOd0FtVSEfgE03+kz6PLgBlQO6wwjy+VzLYmhMo
+vdYH47/EPrI1JHvF5htM8y1ef4E2bKQA2XsWmTpT3br4Qn/TJAFugkixnKDGHRX
lGj97pCbcFz2m8TKECmORfeAJRNMeely1wtvy79H/m3mZ4AaHpPkTGwOu69ZUDuC
WXQlbjbmVWElMf6xvCN2bxDvUzl/Cdg7nSVHjPFBJE3WxDHrWPV+F5ms145Ts0PZ
/OliaFdE9/T1VPi/87S/1IVrwKbxO0a0yjdfBM9EModyn9w0+t0P/p4CqZzPkvbr
HczVqfLQbUegWsQkK1Xs4udxGiI9UQGlCFDFqrm3dVP+d7tKUYOA/xyCsoLrcUS2
`protect END_PROTECTED
