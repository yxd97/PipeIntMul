`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+2o/AZNqUg2/qK83LxQstvUVfawibiNbUTaHWSizKt8eWGZ9Nu14x3MyqRfYgM7Z
EXQl8+r05esfDBj0DbjS+1qycG6RQShTTT2U3domESCM/qrx/F7vclDSUn+1ImVW
J+QW+GxMWgf8nK3T3PUs43dVUmf5Ba67J9wYJ6Lfd944CEkpTLpOoPA2HaJt4rgg
4Ihw5QXRvkrt0xkhulzB9/U0sMvr9rQlZCLbrwD06VTrtMsxJ0iPgrbXUl0wMF7m
28a2ckXEtQkLp4oklAnIFjqLqG7D0t48hTomiqWIMPoXFeBUz1wqjPsKEcOeDYls
by/gCuYeoiwmso7yNAyzVb1rRVaUuFzq7pZrGszGbv5viFx9PK/IaaX+v+zQT1Qi
`protect END_PROTECTED
