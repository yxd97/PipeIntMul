`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lHD5ud2fWk1yI+a4/o773oSH/c3oZd5tpgC2E9+VVj3zybErWif2eUarD9FKmS6Z
s0J2u5JSciAC1DyFnICktjxTcAu83R19MAyDq1+s7Xz3YNkcRvNsRzA31OIeShnk
T/vXSIJJxnecHooZnTFVzCJ+ie/wllPxLv4kE2r+GycgEpShbkpyQY96Q70LUZZo
0+A0Sn2FHFa2tNQJ3A8fxxTRO3/U2XeMPyw2bXyTKPZSN0ViS98+ew08Vj9ClvAz
5sdSMHhtte9MNYgyO17qX5LXQ3vNIS2nb1sQthCnyEaE1DvD+1q53klzgOHKbTza
NZlXTIzDxJinmWVgcUud8gwksrOS9HU8nKBo2XR1IdW7SIDGbMaUDX2WXko1nqq8
MeLnFBkQP3eMbN1pXq8W5G+l2icj2zzkrsln35emxJFFiJZxI83G9j+fuuezDj/D
40oVuWmQsbG5ugk4M4uAE2+VrcHA/12c4NwUGGDjNafjlXxeDGBw2GvihcyP8twk
MMhRS8MmttxOajU7AISL/MgnkpdpM9KBi+qrpoe+FfwYhuUJsRMOwKYzs72mtFNX
9Q6by34mHn/yPN0UZuOH4/BvJ6xcKPNZOGTilR7ZLfFl0xegMso67xRh6/2EBf/a
DRtIr5L52nstKzpKaGCZVUWT98u01rqUG9cXYdg72sI=
`protect END_PROTECTED
