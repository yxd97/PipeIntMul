`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3SLbIZy0Jmvzt79Z1IjoEPeSyHlIdA0S7NgcFit2RkAaId93hUGjMk9r1lTMg/0o
kPPcXZNgELB3A8c3UCnNxaIC/jbfIPsBz+2WIrt6bPgoTxeduIPf9/kSIYq3h6FL
zjOE+++6UOyI70QBiAZ9jEq+iHYxnDh8Xej6yUtq0ApoIiBaqhMKvVTqbuI3DzFk
IxZa7RxClPIEY2o9AZqQFYp9yva3kUIe8pC8ki8bxHXHq8cXIoZxCrDtoPWg4Gtj
ImergRI08pB/dSkUbWRaODLc9u8I+YsQ+XrenLfOI7/M49geLnMDMtkH4ksc5+OX
3EVWO6KrG1JJCgbKjWU9w5ssxm6nBJk4ODQq+Y3CLJn6TnE3QWzTHDtvU/7lV7OZ
`protect END_PROTECTED
