`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YkfntaUYDrU4COHhp2LVT8nPDH4DrymNSMvA0gFH1wL/SyGX/YNl6/jDuOlEeUYM
b5G7XyA+FskJ7rVboCFOC16B/aK1zMW9oCCcUrTf+UETQXKzJ9nOILdxppmPbkuo
H0SQdZDAVwINJr6JNVDT2ZdQ+Uq07dLs9buwk8ux7OBjcVbgeHta7Hm9ELs217Fh
bFMmpeypuLMSo/F5VP6vzFU90yuT5hQyHQJWlDZ/6YH2lpxO15iwVAP5PdhE5U7x
LuqKRbvhk9hRQOSjd2doa4g6V6Is/WQi6sw+x3zbyEFr6x1hMPWfBMtWObNXYRvh
WwaLLsKo1ARpD7apdmhTZcXde3i6348xqu3PApzPlQbOojqK1a/iFS8FInLmWhMb
lb0yZV3xo0To5dGvMt9F6VmYgiA0aqZwLJH8dCWkxdpF+3G/JodEvloh2u5GtKRG
YRZj0aSldZGIQzXHacPu2liJ4K7b4vDExBPZJbaDuiUNM2pdH2HlJXnlV2/glg0o
V4364RbXJLJDxBj4Wv+8ysC6aENDNne0maQ1aoaP5OM5gnEIVf164T6SkJnvryFN
HVFBHuBC3avQeyQ1qOgIw2BkKu5dOokrwHjGzfGO8rplnKahBWGOWZMZuliZ8zQv
R6eo0zzt1Ck8+i3/lZkEVw==
`protect END_PROTECTED
