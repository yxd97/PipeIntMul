`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFVeM0qwNfPWwGIuvW0Asya2s+hlkGbrYaKg4T0EbGlR4Xuu+dCYWIixCyDZwazb
h/4is2vxPXPtjxtZB9xRgbj+EkxSAgckiwk9GTBTaPvK5yq6Hz/97i2mZruOYr7g
jd5glZUVIbWmcMBrkO2xHj3p4HQuZSK1j63g6Jwi7m12CWKFNoIZgrbhn4EgKhx/
QNLjjU727mjOviU4wO/sYla52Q1RX63szDp/FfIC8nRRLm8tnzT2emc2+5LZlGu2
U3WhPeNihCSiVWHooWT8hHOV01qBaTAbRY+MM/eB5QddeBC3h5u0Q2ews1inAAKJ
jVjgSPmfTbyAHgZ+966w/Bd1ApGtUR0+CqwxpfT7A5hA0+V4S0bia04G+aeu1iEt
G4fVXmffpfEDT5lBZdti5iL/sqSt2xDOwdUaKYnLk9AXUQb2uQF9MkkIGuEiYVdH
OdZ9IJRoXira/Dq/lnwQkoVAP/ld8z7wwlNx/FZq72rgNMdHRwiiDlM5hPn16bvY
`protect END_PROTECTED
