`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NP0xd6+ibiTFS9MhBuTHEmUG9o+L3p8bDu9HBSYDolrOYqKnChQFk3Vk7beSvrlA
AZMA9Ntwt9ZdJ3uLNxKRv7t3xGRp2COYytUXDvDsUbeaKupQPF97iWdsLt9Phe92
aCN1DlXtnRsl4oub89s6qL2+I1J+OHwHOSP3Y3sykxmUsDXZpYc/cFvU9yu/ixWA
mM9elCYDacdl/8UkuSGpQ0sXWtv7nZER/5Q74tmFrjb3t5i6MFaeJA4lCEetf7ag
pMkLUVb5xdlim6SD7ew68F30s3yMs4ORL9cnL1bIffjg4s9Fk4f3L55dbIyeLeVK
aYLYGi8J19/U9XZ1cxsdg/bpmxCtd06aisgZXcxup53zxVBU8SQlvVtOmONCxp1P
MyvB+3K9EoUR2G7pyl1SYqK/DEorPHJL0lUECRSxtZsXOpl8fGhbR3E/p7Jl7Oji
qFfJGPpn6phos9vZECWPDobzvUXvGVLWv688M35sS9jNIWXVLB63gQTXH3cJe0dJ
IYeMHJt85yJ7ZatsGlQD9viDsRLmkTFzjhjGy9EyCHpfgYQ6hEppSVsr3e8hh0Dg
BdXd1+ZynCXouBzjgd5XHIfrtGZVs1Ib0Uuncl/T+lKbZfYFcOntAR8jGDMKMJcy
`protect END_PROTECTED
