`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M456f/T4VE1mb2ctGsxCs9t29FWOfzM8jJOhLn8mJjbouRri3TQsjMYD93YXTu6A
zQYOQIXcjn2Rdc0nag+bAH+yu4TlmPWs/dEHg8FvLlMtKvt8y6NbNaWjfC+En+uD
fOjgz3VCLJQeOD+vDTgp/hyg2vw2K4u7azuzm2DQhKTu44A3Sg9mq28XPnBYD1xp
Qlh1+DPWqs/KyaBu9P180M9E/quGTsNOCF0FcGdDCoQ9OkNicMPNGzaSMq5vs7j+
Q0yE/OYFz7srdygIZB2KNLpZoP+eljxhvF3hv197Hy+AGI/HefiYnKOYhDjVqIww
g66iqpN5n1fUMF21K5Rp0O66TPKVTJtoMuZfQaNMSv00mRRdx7ggMAWZ8gpmm5mu
YpGn+PfQcdcwoqDGtv3kFAvu/jibYz2PFclK0ne0aKevmMNjrVhQ+wnEmk7Zc8HD
ACQm27/yygG/+6kiwuuuw5F3zh+DISXqAinH6EWu5eu/LM3lnX4lPK+O0iCPXowa
AbdEgDxWxT3VO8O/RosgqFGJKtpKnwFa6PMZ5ToL1mxAFMYwHZbVugJ6bodF3nt4
X4zuNt9Y1YY6lVrFiqqFFj+EpIWl5asnDjiU/lLLUo+SafoinsvB98ftFe0gRQCz
d+KtBLMTxtlIi+aYBMjHiT9WlStLAH/cP1JC3oICAMvVWX3GKeXU+qaekXGuuiTE
5i6NkkKBlcqR0SsuNvb9IDJ0rKN8IjfE9RzWcYiDXoRtw7qN2m6dYq0M17yryN7u
m6UxL2nQNXw6VBWrNKBE6vULIvxkq/5lmBAq2GwWXpKVnLA4yhRUBGaDnlzhJ6DB
aIYtKV6o/U9aq07Ll/cmiEygd212yTdzNf9+noyZXqvhMQxbXyALxxXCnaJmo++B
FCdb/D99AyCCzmK5FaQQXokdDaMAsWcBmKHA45wiDT71hbxVpleldzbZP8ZnP+3R
hmNZ3W6+9xq+Fie3zLtlj5vvGfueav5NLKYo0NILj8Y++9psZkLry4xLgskrLoXO
3olQ7Bc8IkjTSaEY+CTrThwu0wXqHYBxWwxnB24Gq+pQeVbsjp3Wo9c+vkdaEams
dMyzmVd5ybdFvpxZxkfJRbCrN/v2Nbu+r+asmkN+FCh036U1TyPG9oEVbBx6OKPN
N+xL+IRZSwGWMpR5D0qtyQcmwEACA/QbIk1KGCfRujw9hNPCIdSHowx81GhCoE7X
Zy4DBhyiLCK0RPTSTAHK95pZlBl40dqgtNOyWVv9++CDHEZnjxB42PMsxWlNjRgL
2lcclGdJxxMgP540yT/xrV9OwfE63MmcaQsLJxMSNZNVnvWcBeA1b2VFKmSAp9Dm
NDQv0glJRIWFQvBKobx020NM6SdsSAe2PHCli5Sh1djpj4qHKlj6s3nByfB9YHuc
jiSCYO5E01pLxWHGSbuPMtpWp0cSQRa6NJvFGl5cj1vOh+UoaWCeXipQXttwygnJ
9thVPN8W8wjcvXX+mMslsCX1irOTE89IymUkz3pd7egTHpCw11eDzNxz82EH2PsY
Ygr4frI6WcB0Ti7qzunr6fFq8CG5pQP4yqkAdojrN4lRSuOjU/v5vYNvGNFyFnEb
eg3PZaU8Hjg2BlQoXYY71dCLwDQqlDWgF7b9sfcuOwrHcISgqmyKdKVp9MYNDUKE
gKTG0spFW4IZlcnxZ/o0WhuKk3bKX4hBInxyTo4X09/KvR+lWcyiUVlsQ6KoEcMA
pIUka7WG/HU747iwFKkZXdalsmQi1Y3O5p1jjt8eCZvLGo+F/+br2shoASymsShQ
tHyLeWSbHEw7QC43aIWT73Ky5ZOSa7Dt/OZWzzleHYGPi7dKlF9V/WioLvUUs6qR
QDF+UYSlXU2dcgTiUxalaKQ2IWrsB/Um3nRemZVZf2q4uHsBa2EUt/RBph/+LIhJ
f493rkETYyu5TdRFMBC7htpkD7SpwkS1lGC7HhXHCjfWBI80Y0Z1TWtFEPm4w8yu
GwkPTwYvlgco3+ta1UU8Uj78RzY0ELBSgslxMDzmzoA2OpbD9DIIkXuwwZphQ1IE
famFXJ3u7hOcQKe0KttoLkWY7e6Xe4FlhrlP4QgxioUlrgE0z6ye+fTbFhYF6I3W
1KgEGcEISNnp1dgbW+lIY2KvG1jhPDh1mRlXqXAy8muGaickGCCsh8X4PlbqlbDr
Oj4cRD0N80URoiLj2QSd/mAinvKUr4bX9HYI+gD+MUDalKlg6DYB97qCw/kxwE45
BAeCj0IacutpbzBc3e41bFwJ4kF7oVgcBp/smKl4qY0dVxBtd9BQf5tZ1pvyOYiC
kL3+GGNN2/mHKZAIi+xQ4An3UkxcMBRYh+4+4VNuNKsKFSkiJsQqPBirZpmIdz0Z
lwBm8wHZr5WHmdEGetYVlCDT/rNTCKvttBgaeYb8fHofTsjoy2pI7bLPTSt5vpEZ
kWM/obf+7+bypf11KFsbYPd8ajMXDyqXAaQOYQvbM7H6nMqfGg47zRb/GhxfQ66h
Fp4TZfGpf82eXXkHIq0KAhhuAKvdeUkZerMcIy+o8OFwdz69Fke5TuEVVESwYvIc
IxZpgwNZWh3iSrzlSDVJW6WQTsoFfcuJdAUBFKkKtUfqfVjzCM96kAP2NLjWTIkh
yyirtQwHBQ0gSj8KCzZSjWr+0tI7mXToMjSAYeTpdnueJtElaD2C2weNFYIv0PqD
ko5XGzdPZsRNtK6rSStnDZkKKfEk3fXqW0jWls8wkLJYBGTcyP1O/YyUp/fKSnoe
aXD7f3gZ958RzQvSERaYOmtHK7L0lXv6lM0g22VB+8nL9bNKQLWKyiaW1opxMXZk
ETzHegkxTH4kyhSkPeA/oGxZw1Ixjf9rXmGa8QmYQ6pOcDCyzmL4j1JYcTzWdQC3
dB6u5Z6cyDn8l10DJfHddy6VP6nNI5pvHxMB35PsTedMmlIOVmOkvOKGBgJzHz0L
JewBkFeZQZH1HQ50067frGMfyFupcSom6+fmx+bkm+nL1vjb4njQIzMM5ck1MUtG
+ITJu12MbmfPDZy/BjB8CTo9qVBTPx+RgavjPACXK6PwdzwyP5eL0Lgo5/7tMzPH
YOUBoN8FaPWGpxKURAn/BbDguwaAOs3Z60SSIdYV6z+y9gnhRkl+Y8Nu8i2ZS8Kf
JklQgVhF9CNXhLXtZl5uA6ITLhFDmyWtk9/Szo5U/BFRJtPs+pGpuQatpjtx06qr
5DQ3E7EfVB5fcpK4wchmCJMmh4PQWFaSp+3LgwuZGN3haS56R4s3O+epdeM46o5N
PS8fwUjLErR5HZI3/abZgcKRUnUJpn0GMQ/z52UOECrof9qeGwgL9O37/KOsU1ux
kxGq822rS6Sh7bsPuyrWTgdHmFp1qA8KYbTeXvohuZJdbp6MVC+Ljh8icag0sH7o
hWxx5YDgJ8b3cJxhyrdyrfA411NEfIuQjeUhGCTTnRA85xxSTnmb67eA/LU/2eLq
Mc+PJqSlvGkV/93Z1l8mkz35wPp1Voui0mtJ6TfdisIqlbbUE6Z/iyg4YO0GiGWH
zBvcoPxbE2Cey8UyPv9FjLUzp6+Qlx94zGOQEgeS6McPoGKww4DBVkRLeZqTtzIb
HFnnsxboW9VOppnEluNOuhwE/HlFBg+bR7y+D6BCuixwDCGIhaTv3Vtgfr1X3Ls4
LyZo3V+c1OWnZlvoHmJiFdGtbUQggZIN3i+m5ADj2Dudk2Yu9q6/L67e0S1P9Z0N
zgYSNTmPQpZ2jRRrfM65sy8K+ww+AcI4dwpyu5N3Z/Vb/9Cqsgy+JJhcjkglxJR6
4zaSJWvgLndmbEIrjTZvtH1q5YXa/UZbBlzMW2yggtAwdi+1UJ9zOvxMtvcingmR
eSXOx1rbnvaurCHESaziNln6IgGVmxksxr8zgOSmvTTVKEQ2qNuHfD8g2fy1fkIq
RzEYCD2T8XE4/AMsh7pTWSMzF6xtT9g+fd2kMhV1eGXvTbjge+ZZ0PxiMx8cat/F
p3o1Y3DMkUvo3R+NxXNIjdH7E5LlA0QFLZztoudXOPfeIQsUeLEe3RCzTWnppdRq
5wejRqOt5kKRcVybZzbnYEtuo/nmYMD+txzIBzek4zKJ1U40wpOx6aFS/FuTJIZg
fLmNdg/bG36LlF7tx6eHp8b9/CLiSe7Rg2IHMMSXg4eTiyZCZiulSqThmZ3Co/Qh
mVISMJVpzp5EMfxyv+FDDAriOoDU0HA8+3Z0eSB0QqufuU7Vo2NTsn9UHCxZV7cV
eFRqSAlcMRl2BikhbWryUQ6HXo0Mn6CR/dO/9TdUTTUWCDlpLzhwv+8bEODUMHi1
M1z0FmmWxkQsZo9aQNZ/qP4UaytVyZUNdq1dpMKPm63JC5vs7TpyoPxIUsF6xhyV
Tx0qmNH2RoOF9+YQRlQOmISobi0RouKSdxUWi3xK+kh3ljWhqjav6XJ7R057a4AN
UALAtdFsSNeTs5aRbsdC1+Ek2EsPuJ+bIPK6olo2fwrIzxk86wMsWigHD4j/+iuq
lqzvRPHGe9smGortA9oM0MTNzXGt/IzhOLVTLilHJjw2jMWDoQOMZTHkmxMkQjGQ
sLlNmBc2oCO2GdLwpWJEzKji+T8q2Pd4XvWEKvln24QrpL+e5byrqpzZE57n8dQK
Y2eJ9jDyqdy35ftRcUZfelx2R5Bzl69Ukye64U9k+fXgqgb1Ey7qUmNqdE86lnrR
vssps31XC6nS6cm9oCz+qK4/WXtt1Nl0NGfIf/9stl1ebwL8ZBFgjza+OYLERf+G
Qey5M8R3CJyTvVWnp6zMJ8QIQYC0CshAc8ayTmrboZv8RZJCjrCXV+a/NafA7+dm
MDJcOq2Fu8c0Uww0e0Ij2oUIMGPyXwhizmLLnKAZn5SQ0c68L87F4HYPCByjJdfA
PShwlQ17Wx8doVwGJ3ogsplFh3XiddIpq8+PZu4C0d5tsrAhYCiuXyvqLn/2GuCb
xmdDNu4moPOGPP7tWwqFcKpnMx6AkLuUAf7ANzEkHZWrbmhzFe+O7oNmHQPZtYJh
5c+ziADnShSW+4DTmzzfaWiqF8T8irPYpsGlDbEOthByKpjlhoSiRJJ6ZeytXPB1
PZ+yhJETvIiukaJDTKIY390NSXsLR5Nwp/+L58qUzuhSDtZ71hKrc7UtTNhHqpog
JDmRPpX4SsQUDQaU7iED1TEzMmi+JKNqIALqJULU87zAXRlIS9F771RVPdX5Ugib
tF7+/JqHw6icGqVIiXIKKnvRQcsWtB8dmq8EpRjxutLb/8nX5CyNKO+NTSCMQcl/
KVyFvdc0K+ut4qMkG+QMgXuueB+rZBXuplU3mL31vNQnuBmCzXBNFuGJ/3EEn+qB
VdB2Lb+z73fYPTb/0hrJPmlErq2wh6hL3ZrfEg2zdyw46pO2GN2lX13vTdfaqYhG
PyHfXQSJ3XYMyA30nPnwBotm0DEc1+lDrIudshO7i/Qlo0GgHCZ2nG1H23hwz7Sn
YlO5Z7eH7Cm/uCGYYnGbduax+ptJrKXxNTff8SbLgDXpPNx3U0zSSbFPPcqI0p4W
HbGOKVSAq3P/b8jlFWcZmf+mDaQUuyPDbnOo+2QFrPLsUFnGX9AFWZ4UXexPidIx
7qZxG8KxkDW0o4ThLvoRuxqC37hyOAEVm/JY89mo8Fzf6eDc8z+uI3FmOA6Fh20K
NjghqUryD1zQCh6ObnTnvP/Zdv19i4Y7SLj7Xah9xLEgynpegtjkOXBCAabmA3kp
bGWmhhRCrz+mpg4FEDnddQ2kxc4nbhA3ermoQC+FtMJ2fmX3AfL6/9lpvY74LFvg
APBfRw764hg6pwmGGaZJziQDzjfxlmm+4QB45VNk4GLrsWTCXPyFRkZNfz6HKTXC
GjVjdaF6xQ1vylbc7wATcIX2Bo9VL9eawPYVchxwnSXJWDU0H06Hh3/4TTmQ+DRe
iuLB/1oSg5dbywqTxXVLBza2jFjTvRj4Pf84575eKXXt2vtKCr0DjwJLozTHowRT
l1Kkw3IJPFC6fcYAz+rQQu79HA62B3UZ3CkiDZVXhaw+yglwkN1mctTVZji7TugN
EUrrysi+3IVm7hke2UnuT0EojVfc4Xlcfh5e+xzYKDjJKUN2/IVc887I+axstkMh
ptkC1vBKctjPzgEZoSyfRXgFkMASTH8X5Bw7pjx5grN9dWKi98D8lTZibEnTFGTP
t54SgaoJjhODa1svm57r0mGaPTTE7O+PBdvARviOdixCcZS04O8ZUFxLrZnIA3Vu
jA9gdCnb4cZX3oab971mky81K3AWd7vIcen40KhJPzimQY/SnEk8E22KrHz3GvTL
YnR7DegF0s7rRtxq6OSLNr2EWFi7UpCTIYsnXQ1NN0Za3k5UOFOuCBcGeXVPinzP
qAojuw+zr6i/5+V0cipn+BgHuI5NSx8q5sqQR837Yz5zZQte05UNqkPRpXzZ1+f7
H/CaDpC5ZTq3iT0i8IlEmtkat8hme8/jwzRh6uZQSeVBKfWiI40/cUopihTGIATV
J2fPOSac/tJLBIGADLGEi8wke2McobidhxqdWnkHRBJFZZY1+29DGx92/eXQa8S6
dP+qSVc37vULU5wB6gswWI68PB1AMeQr8zjs+LyjccdkKW0Bi0C5OWBGfxuAWtOW
VZekBJ5Sr8n2lYpZy5mk4/89POf6FgQPEukr21v7Mo51XS/l+Ssj7LOzfwYJJLAE
Z7HlVUb4d0WGdPKH3bCt5dhvsz/Xmiu0xZU7DWQlgTytag3isodZyLEk79X1tp/s
NCT50laeKH1hFvLWvonlk3OJ/RY+EBgHEMMl8An0Qbl9/J9CMCpKd7EOz1NRgLwk
iIxBNxDF4aJAZx2ExP05F33Mez6B3eyOepsgCBHDcDcTNwgg7+Bk4tB5AATVLyJi
Inb91UL9RhQR3zZr682mAQz92CnWzOqCUZ9lvxu0Yyo=
`protect END_PROTECTED
