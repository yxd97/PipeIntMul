`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KFbRmqhh2W99I2KHYzNiX4q9kK+4QtbgCI8wczEbSAOld7D61wzoLou2UC8fKJdQ
x8528CFbWYGjtGNNhifefr6KEzB8Fk50liLHZwKJw0eTfdEyo67JeYH75iopCE6t
p0Rwr+iZS3hIsJ4hacgNLhyPXL9yzmYBkjq6Bp93yFGiVEuTC18qp1ubxM506/zi
f0O8sBXljJwZbTSSU+WZIDOU53IHZvXed3lC4053u1DWxObGQebiU7gni6QhhqRi
g46SIXMEe8z+3EIxdiiOFtxPjNovgqcpADeiWwiirBNiSIPNNFxy/8qQ6Pzx2Ruo
DWulzdz6A4OKmVB2mZ2WAWUiyrUYZhtg4nBsVal4WXzIaBNAJnAh1to4KaR1k4a6
aa/3MVISDBrPxqot4KW34z5qVYZr+S3cj29CrR0sk2cHKKMuZXYXyfF3/OysyKJY
FyGUJ+VPvUL1o+rnWtmDBBgigGfqpyeWFC6ohxB3ypMFuIkg8sl52U75epz2cIXn
vi+uwg5nnOSRumeoFe5Jdd7/i9Pwrd30ykBpqu3pzxqbCRwrXDSg0dtNAPbchgih
`protect END_PROTECTED
