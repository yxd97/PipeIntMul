`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DahIxq6SAQ/u0SsYeMiE8db30wnPNp9/vMoeCUUqFcxfHPHvFcUUeIeYnypSfcqm
xbUxh5tGzGh+4REC8n5E3X/6Ij8P2dFpcN0Hjys7WC7h4qDLf9ezMjDoFhGmSs+d
eRdRHBv7/dkj1B+FFymWZUuAZlKMolzmyord0tKsy/3doPh0oUdyeEAPm5b6mwlL
NfmmIypvptMOlXyZlNdVEcecRPJilsp36J0rVBXH4415NHxI83Az0Z/tKEiEFsVj
e4ve6gPOxKTgg2ppGLtq56nQuNcyQF6pfCQV4UGyVbQRd5c+D8cGyUQJYpJ7yN9H
`protect END_PROTECTED
