`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P7tbvCcuxhl+lJnDc3sf8jmRoXhLUdKTiyRosCWSEddrbaBmPj8ZJWeAjJkJP79N
482A5TjtzgTrYKJ2Lzs+FdThClgY0fQff3DkYhfpbRtkeZfpxCgl76pjkO/1WukQ
cLSRiw89cOWQGB82RZWrpvgGrvf8elszLpM5Sh5yuzs3l5Q6HfvVwZN/dZEj/2zK
fnL/rtLRoh+Fa6Vcxz94ag5fRqH8F6brbVTpp29kkiA1ZO9zoD65KpITXvBrclL3
ozbuyKJpBwNLN9mYhcYyYmCa/M1zApR/abMXSAOBZH18Cash3ynX+BdaF7J+3lH9
IPpc5HEzGtZ04DqFqfWJjKVAdZDvFQe44Pbmr9PQg+YVL5Fs8QolU3dSiMmMP6Wy
`protect END_PROTECTED
