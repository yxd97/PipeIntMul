`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l2cfWXpyXXKDtaZ63QXwZCOZIk1fJEg0GSuZ33qKSGIDr4i9STlV811s8njFKlw3
DVBay6CieeetmmS7p74hZMu8OL673XnzOWcacsXY4Fm9cSq5C/rPGfPlg7IOvWdU
VQMmscuZLNImduexpRoRAK+ItarBDfOp+EgBaGD3B0vxtXmjHz6XvaUhz5b4oTFi
+QzrlE9Dsth0vHjDCzGWDBz18W+5goCsCl1F7aSNZhhC5SXG2fuGWuCU01/dF74O
`protect END_PROTECTED
