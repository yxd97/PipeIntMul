`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BZwVpfRrRWZn7GoiaSlYwt0Tu6s6J2xiG1kfbEqAPYV3RHATvLrthB6rqUIA3+WT
fs/OOtFkISq4A0kXBZdNNC5UJaE6LOmo0xTzG/OT3xSbUmxMqNYXx/1ZCqQWTSEc
bMrT+S5iNZOaDOQBgzYOKSm7ctGnVviZ5GYXD+FATzG4BmuMkb7inHa2Ov94UIbc
J/PM/CMoWCc0JSaalDbfvnpWZD7A52GiOLmbPqcC6T7rBSmWwsNJdRpsUwgjE+E5
9KoKknYG64Y2FvXDDZ9AB2QETJyprVZhTuNNPgDLqg09U/S/mciMHX+BISB4/cvk
XRUcqEweiYw6FSSj/G+XRNvJBPB7MbJdsudW7MyHVhKqD51rd+JUTSzG6zxRz05O
Owm9Vq+2C4lqEvvfHTCbwxE0K+KZUfTx7KY0Ccq7WIDA1j5QYgMHPHWG4z61JFgp
6itZ3NgK0vzeVKHn7KGzvzULXP+MZJN10eSzguIwgyGirNGUBVStmgi/9YyJHZE+
x/2JxqXXWynY8u6/w581fsg/ztfxrjGT5mhj1qsVmP3stfDGwaXnqYDyBKejTeHI
NUPM/G/PRWtqUNb3/8iM6KLzYMpUA8pm/7QiitpeuhnpRxkSE3HeqngMt5ETWcvN
T9Rm7SXf5fKqK/oKMrk30C+qFLmnJILOywuKcjZvFplMHJxhgtY6Vid3UDI7Rv3R
2TfGJOa2aMSauHCgWgmDilyA8UoHvdWHtHZxV+lM7M5iKbHO6LJlWx0vzHhqq8uj
3ir1zodkVdkqHinXO6afXq6cu1gN5hRwuTyjsS8/SvM8p/02Re5Ca3bWtRZGI6KW
PZyWvXy4p2PI8oKNbS/R/pM6EIGSewXnihMWHDOq7DBXtCkAWJEx3LX3hPA+/k/L
Q6uVVs/Ca0YnCjsbxHguxQYX1MTUCTlUHN8shNFFBK4qkzLFf1qTKk215oA8BDoD
IbA1DWZlqgX8GqArMxtpeab2KzYazvkcK1k3lW808PMJF2mlh7GXfiMo3PxJrYr2
kTxN1BIZBXbXto7FenGMUL88fdUHoL/esKx/sVQdUbly6DMSPY+Iwk6Es1QvYOnp
JQcgNyV4SixPwxkz2xvubhFlHhG5BRQeqSgoiNp0z7yrO6J84cSIhCEFd1nR9bp0
AB5ITP+a4LiGF0KEApCzHdNjI+c3UmfIgmQTJ2Dy5XWUIgT21nG0Qkx2buNh2D57
Kwmj2p48vio/xrm7T/KN0f2uVW/Mqr9shGTvWbyAunm/Z+IIv0ud0oGtEpLKpfyX
y1eI4f8/zoSNinspYr7q6PykrO2VwseTEZH+PyF8kX+BApgy7Pj6vzM/C1biVTHp
RS9ahbBON0izmSEn26k/Ui1fVtzhoAb8vLgsgZO+F8GDKCCaQV1c6lD5hZzULk1D
wWkvEszDirJvGVjDZwTAyIujoRoB/HzQXTkBGjdDTWbuFkMdM9IXvie9clTEEGG7
uzBx9uQvA9pw6bp+q9RV/iLUvICRfbc/Gf2aozHKIq+OduJN01ToXGqDl7IRTRxE
xzOsL6E/TQA6JYJdgUD3wrTMxz1DGp089uX3XAXNkUw276hxNeLXtIG4R25GIHqR
RjstNrEVBbjh6pyXFoN8iJxS2oqJVndMitgkuajkk6hVHbYxVQhSi3StQPDZQkYq
kR3JKiXTomPdpWT78Vy4qi4Xfr87T/RNsd3EoqoSmAevY5eQUSNHYsOjiYJr3qGV
KKK5usv7lFbd5ybQdR+5fUjOueCELQp0DDBzxkCpGWOlqEk9z+MDiYuW8XFzmmyb
q2jDEFdPdv71Tn3yUPep8LFQOVVfBS8T8FzJGXdJWqa7VArvRy2T2TAqXpcE0Q9Y
JeU/MqdU5j17ncy96G05GcIsjzEafiZ4ZRbDJEJquyirL3PRC51peaKYo+dnGw3B
GoTX3eZwx+lmhGour0XUL885qNU0WGhcCAOU6tSZYS0vZxDndbleKd9HZ44IMSc8
4zF28WQuB3sPIVgTJmC12ilbtIJ+HC5mXvwSMClJgihWI7wrJIjAa83lqX0lUJlJ
Rp+lWdLohK61c4B4lmAVTaLWKrR94XKHsWP4eR4urPDs0aTqWeI5oAIk4ZNP02DW
PXU4n5E06Ldl+qtG+8bHI+kQZP/tPJbZWFqbYNFJtoI/R4hh0esGrPezZ9TOLpsp
BWS7vwCnmP9NYHqnKE4ESnJhuXdFpYyojyxMfXC/srDur8t4DEt2dU7AtYgnL9jt
kbf5z7v5SQsf7qKBaXZNTGyrWLO2esXu7RNKZFysgxh977UJDtgqJoOP3tu77ZdO
0LeBP10x5pq5kC+bvE3Qa7shQzTUO+SrsUNNPHWsz9PashAGjgmcXUimlJaGiY5a
UZxRqlfI0dHVyt1FYDBgSoODkFI6wjYYJFodqsYd8q6qQivQN2jejkwNOK236CLK
fzuhbLbpEL0FpeJ4cGkjRaZzEW+CQAJcRZMUeyRgFxGOIJxlrc5qCjcLlPLroF4Y
4JM+78APfNc9eOLUQ17TaC8d5nlrf6GhuOz/xRex6GTC0J5VEjV/swkTEhOCyAKg
wbU68jKQecMTvKr05c3Joj139JYhQsmKnJ6FWSIcsnYH0DSTOkcCZJZde8/lkVA6
ywt8p4zIkxx24BKHDju1uxcGDS2wAhFFVfyfifztSOG1PMvgEWwmeg1J5m7XMFVG
6EGpL/gI4qvVucywjg28mr77SJIPPjBSspkIyc4M9QUq1+V6FOPApnXilFo0B/sB
Hxq6VlcUE3maihq9/Y8qvFdlsy9P2mYf2fqnM4zpJ1KRsA2fOspGgnz+cKB2o/AM
z3rtAxspnhzGs3l5yZf0HB8Hfr9zfBGanpPqxpRD0VBzaXl8kwfgQn7TLmXOeMX5
LKzmNN/org3//GtBla/AMs5Uv0OcXxPfgUgjCbceQsyJKBGtj29SqUY3NRKTKVKs
e5ptR6H6lrjjF3da9K9A19Q23VYcW3A+P3/iGYsodUpjf+AzDLq6Gjn8+v97UVVc
rw5m1ZcletXJr8Hpy0oQ3UI+9+9SDNeohJjZTqpfNab54Pvt6IERlkjlf2mOCpKl
aM2LhG7NaznzeIIA0DNle4FWHf9h10Z5z/dY17yflIlTmoPvFVocJdxLSofoPrzq
uOyFBVHmVeJAAdtfT3qLTz0z3qQoYpoMwDL/DGGBqaPlrnqc9MlWZuw9T9aECVgD
B+9V4/ZIgxk+VIYddB3eLpJUgxECBksAxWWUjco8ehW1pcJrlV052zBXTW4HU2bp
iz9dK/6XLOcRNqe9RHe0cmYDqNDKnZ/IAc7Gpv5V15p1PvqU7RoX/xRyFM0A1hPr
3ZwnYOIm0aWLnnTL6TA1nThpu6ME0V0wDH5lWZFV+D1gT1v8yR+uWrBD/VhEXh8d
QXHw2Q2d5I4fDwuzIcI/jhQrA93fz3fvsnmCw32fE2sLwdLiI4ywac0mPO5FeWMY
CcWbpnTeMyobTeG1mdfTk6n2ZQNQTwKZeQsG8ESsEt00sLFrSi4JYq/mH97y+NVl
jFshyr5rcXmPmTAl1UGy6pHz/D7n80SZMbwBBAqyQQYXLpdOSbUUHxAnQH9FcKdG
1WNKuCKMZOXo/J+wqxC14tA145muXpcOTw20PJ5rpvi/WhPs8WJrRiT1k+QRGV7d
1ckTzo8PDt1SSFjJg7YdHwBoFxqN+Un1v3djiMAN8HM3bEl6NXk4v9a01F2eAjOz
dKnnjqKwcsI4rbqB+Qq8O/DmtqRthxrMQyU68GxRggfn2+MoRVUmdeILonixr4d0
gNJA1OEv2gddhSwQB517CtDMlBgrTu4ABo5UsfVsUviK7eIgZJOzYJjAXGZ53fQ0
b37UMoHtjDhWbnBpvdO0pAqzt1Pf7DvBSCLoBJIJ99mlKmDr/prM1zlNtSs6OmnC
Y2XlcUZQ813IAkgDRFIRUJIVEToMoXSdmY2lNOeN5rVFLMTqv9Evdg3d7AkPBrwH
F9+w37TkXzRjLGF0S+Xpo9KaR1fU3pvTmdsjX8Z5MKRpnZSv13hXpPf4JoA1kCry
mRzyD5+X4RJjcwiS1SLm84wUafAN8SsudORVDIl6U1Blh6vRGGoHPIIMa8/nqZNl
0xjVbQMyxwYy5tiAM27LFwFfwzYPkJX1nZOUw3M/95QTAMQrzpQkd+8WvgNuf05n
XyKm18e1s/ZjtUBUfNW7ZHslT1z3Wzw7n4lvQODnnmud0gzWQBsJr13T9zzp2ePk
YNNK1jiQcweAfU96YIay65tHiwZ+dLy67hbt/y061yHac2XHzPZLzqJqrrhguH9G
8+UNvS5uGscopkdJqjpHckJbI+eBcBjqHiPL6GRWRuWw0two+Npxw24XChOpQlzE
N/VBQNaf5xjyKJtPtIldCJ6o0m5Jo5zS+CP0qYPDVRJbYtZsCc34MBLmb9U3lJak
56R4Zptwp8h5Xq0Jmc3ko53IVCOFa2dFiu7gLnfHbXJQVb8eGLVM2nspqAt3x9mf
hMX6dUjlZu1tyqqGzQE41eSOkDcMKQGAQyU/Q0bzp1eCimNrJkERiR9LAeq/1Ho5
VMI5gUwolJO54D8zbWrwtMdbLFh9g5o+y7VUCTpxorGSZy8p2tRusRKxOEWQjrkz
+5YwOd2CKtjy0kzCha73elAfl4bhdodRfIk0ii514IX4yGvYUkCH4D0Bj8axiGAd
UNK9ZmaBxJCWkrkf02E/wWbh0tj9lHd056UIh1OehAjqfnyJPYHOz67pCqS/0IOb
dMqBPQh/btfxea/qhYH8W+9XxK3VqBYZ3jAFE/IF1ccKCJpYtWRg30q0Hu/JnJrh
r43bGfQ46czri5FUe6UPlF7XopqovlXUu6v34eF+FvylHoP37LpItcoliMR+tXeN
cAytaapctlGtFtPXGkmko7sKFmKk/ilsmzenChbrvSxRB/1U8RDmSudYtyl6KeUI
JkGCD9EvnuV5aU/Rq9Tj/YkZrbAA8EKdRqJWZhatKOJLN/rdEHbxOwGUX923b7wz
DSoziJBdMF96Ln7OAJycGmb8bR69B9S/x6E+Z6TKi8Zi+od2nrYajCmTcY+zfxGX
lXCOv6YTsjx7Pob0IskBYTCOufsbFpKoF9+8mr2YZ7KeZY2GG9QGPXBqmxQB0pOk
RKDUHhf91Yf1yuC0AlQOvFCF8bmueQVXEBHEwjndckh/ZQmGwdMCMMLMDrVSdd6B
TnE/Id2MLX4l0SPV+qMhXLIggqyILei410K+lAMLePs7K+TJqGnpqhEBlhqIIMVS
1ro3D22rvxUSq28gQnCWWvzv/bJ0By2v8KIGbuPFPBgcx17p86ucQ16cyPbHP7Z1
yhSwSmRlp51lyvQIwlYM+TW/pE+VbB29It1fkvx1mEo7Flwaz7IXmKfLCcpepM5j
tKNSkJ1N6VUOowN5gkKWDZtUshT3u2eqWXBRu1Xg9F4dFMh689IeQ+LKxfMVZSd5
Npy2gfvt4NKQpj4OjW3Lbb/XvQbKRyrdmXCiBbfkNChZM020HUt+ZCII9I2vCiyb
iXuO+AZSowpuxHNz3FqpNOnMyJr73yk67v5/EwFN2QfdcJYq7j2BIedFCcgRiYi0
YssDiHTAhwwYlBZJruM78LAk2SyfgfpAvWQLJTN0GwFd3lstvtZZTG5fsgcvxkYm
wz8vAntN8F+T4S8ehuoxMgleLmgMsJYxYJqSUYNFlRUbp7WOZGLL/KVWOVD2WpZZ
JvfSa5XJwJUibP3Mu7VoKWD2olyoPmZjuAOllkJZM/Udz1ZheVbt5jGMzRgNrwGW
QJUwS68vaofuWoCLal95Hkt/jB3T9jN+AuDAnoPEOUijnb7IK0nYcu9ku9FZvPmY
mrBURAlTvRqQRZ9lcUArqtPLVSVF3dcw2SRxGNf/eJ1YP/jv2VW+xpdIWJlzQlIT
ktJHj1YC/ei3LiPtrNXHZHYnNYbPkh8hqVhd8sFLPCuGQ0ZYW2hNw/Mg06KjWDie
xU+2AptONT960JWPl4Rnc8F29IdSHDuTkTk8kROmmvabgjXrl9KIgoUyVYfLiPxl
BkLX5fr9eoFinqbUrgtbi0PhexyyTnPCY5C09oc9oIsWLbBdQVyTfnDf2+BkszXY
fYxuAwRwnmpJ7lb4NZl/pYueu2pPLQgHSBfROGFD8IjA4rK4pfl7+Qq5oq1TRtUH
DdxWgDNIx+mwCwDCAJy92yXG6paVtMutVTGh3itqk1d6eM8h0zWPh7c3RMFy2Cmv
1ZPatFg2hEv6RvVb+Xx8f2ruVSKXvqET8WIqlw3nzPeMGMrZM4qgIXyhc49qwJQh
Dt08Ww9YvhCK7UoA3JflGVhJRUae3Z0ftt5mJRSmAQRXjksaWHQNvc6H660iIMey
3mgbAR5YeChH2MspbQLS3I7mmrDaSaMwId9EFwRvO+AaCbNhWCRH7Du+nwZg1W8O
AuYfz7e+0Fy2s+xmav/9HG2Rp7BTEUUnCDcfCAV/qf0e4FEbo90eZozjhvzWIJbD
5sqbVLX6a7SOZ9Z2i6gbbmHuOCVSeSdhxmMhgKgfoJtf2gIr6LlJv6VB7+XjhMEL
ldI6bX/gV4w/kLAkIwS3b3EtVb/OR2MgfxHuWm6W99wOjq7X9sLTp55WuCSCMTJ1
JUCcrPKfK5c2Pd0nGuEh13iDHM9fBpqQTdvb0Fc2FfgPttq+m341E89zhH5Yajq8
lkN3ugglbwciwVh9twKcA5ZXOXFJfpnIRnIacBCanCMZwK1fncfsCD37+Beth9Nl
uMYnAm5DzHjkQWxpEaf2fHTxoFoa3sqvHlbwQoNB3c+/50/AIhBrLCRNCf49ye0m
g+VDgQD2o6I8wvc85KiOQj46qEo5GdLZWFQaNm3zSDeMiw3lm4BG260a5YpH6x8t
/eoUgFO6krbjsXH989E/5eQaQsoYb3IDQTuSQpd8LST6j4NH79iSi/QSiKW1ps+I
2qOVgF1TzC3AZZXG3I+QYDQLZiUZXPv+YkyfVomPbEfwvOMf9XxxTjfXgEodk7G6
PvURMLwUdPVXS6y6pLXhvZa896ApGHfAzZwVm2l4NAFe7wn2fSnlxT6KWvmvijAH
h/C/diLoFxp8BZytHc3OV5t5O6uwsws4AJBHx2CjrbVI42nO6i4iPVe27uN0rmyZ
LZC3JwnwJ+FmU1SbBwAZcHl+9QGxNow3Cg+1AFlC3+LyIiOF9y/jE9mSXRAIVW+p
7gFaNaMqhM+e8MAdkRk9iWZ4zE44wLMpd8x0tT294JfgBxv7sopioJ+3sz4K4rbd
xx7TNKTZicr3tTbNtG+Z4I2xhGTsS11Ek9ySYGH1MCwOywwcOufiDfV2xTkRgHap
fbgDeUVIYIljyqLRAeOA86KhZSUYE+fiynWg0GXZ1MQ5xWV1PFOfy7aKnJQc1o2o
0RYeVLULt/THJSQKhAjcBJPmz3gNZ7aZAOUvZ8hgBc7/NtDoBNNd+1pLeC3lhMtm
1lf3jIVE5X3zMyZweS8S7bW1WpYeg2FiyGWqnLb3oiF/sVbmHHtYwI832ZWd0eNz
/9+jY4fePoZOVLe2QDqjfES0ii0cnmwaAWbgjAQobsIgsaPm2rfRZ6ECVThpiIZ+
V1zZA3ZwLntvgUTDtDOXhR6OX1ZfHsaJufDL1uY1PUxvUApfJk2LjZcU4yh9cvlF
tNBAPQ0L2M/ph/NfY0Y62x48niy9FG3mkfT/29CdxROz6nEG1pETZYznB3JFcEjR
mkWKDH9n74spKwh2YX8bUnyzgKxutIICANGWXaKC3dtDSivL4zNSzjT9+bE2LtA8
JVA6+yDgxpgQ+6taFK/cGEO2HOI2V3z+vpUEC/f3O5iQRrzGzF/wc4EMEe32rj13
BxXkavUuNWJDWdZIjOayKaXkRpQfwxw+v6KbhBdXfuEJK/dHS/AE5ebVo6jySx7w
F99sLXaagRkJMDSeYWlIH90n0dtRnOJi4zjhPhDBGA0YHmeK1Cf67siinwlg9ya8
AidpA+y0TBF4712toPqMGHvnneNDWsmT33Izto/EoMiKZv68ENxDTr13rDxsyddB
10fYDQQgemxPq5Mhdc30EgLnle3KxL5vhZ8kjgXKvcPJYHmwFxODRiU2N6/SW+dW
qJDS46y1n0lLD3jenF/NDEZQdQJ8iJtmYC2TB58wu72LrCv8G9iUiTKqFw7EijCv
tShUdMOqQJZ+hgq/n5QliB0MiUPqg/eZ7838lu6Sl3Y3nSu+ylhBgg5diO6KalKi
ApqoNoXmHxVfkxEhHd3x79lqvulCcAYc7kfTYgt06c1DbqDL/zGStrpD2ToDCF7M
35Jlo4GRgWTbpABcd7BBV6O8sag7RIaD0rC2SUaRwWiSJpLsfvoJ8Lys39nhOgkL
d0BXCaFAMANFapA0Cp8lbymqw5kfz8iIF7NcnT4KFfyVKuac3sBODSAq1wK8P+mU
1C6+kQZMJSDtLlKZnajApLSFUEzL/NP8LTw7BWPa7L5gNeDqZaGDDjwAL29vQcbr
T0c8Rwndh6zs9rByMlSB/S5ASyJi6TFaRUxryWtlM3VuAH3nSHTjUhD5Pg/S7V0l
8lY4oHOKiC44LV/cVkKZxR7hrbZJmTvMsQ5f5eLW6D6BFZB726PSW00zXIMQYTHt
9uUH21OPmLCK8N1PjLgyaO/djuR7T6Fte+riNWgnKT7fohvYy+SoePv7YI0czAj4
KWoKNYzvDW0B3lOHbjVlEXbJHtGaY/Czfvu16kN6EitbCpNQATMM6V2DO0y4g69e
seG1F2itapb3fzzgNhPO/L+eHEpFknvyhLRobw2c76LtjECu8mhHtzR8Yr98XFLa
FZmBit8IREZxxfHOCZA9nhe18eSHdAfkNC+g+wyJMqt2RZkHpYlhCXVzrlyc83SM
Rn9EqanTqtB+eqtnSszcDZtta4XyIhGPLAInkVp3voLHDbEpEn420ataaYnFNlQn
ZTsyRPQo6F81q52DJBKfZCtQ6mTcW5FY+9ksxVJPxM5lu++2/Uv5ATlfxQVm9G5L
RTWqBsSww/gF2WdjmSduqBlJwoouHPFH8ivPHncNTLxtpOHTFwR3ki6VQgALrs21
m+3LySPD3o9rYVqiwdP/ub+qhtjtdVvCT/8Dyuh51020umgzwJwtamtGMjm7ODyc
M6bnuiHgULQUzkAxQAw1jW9xYlgfkfDFGkJgFv1p4+bAq/GrNCYius04aFMLjqcH
NielsIAP04O1BaM5gXa6ftcUw0AvFvCNibrt6KICrjVCkOBXGoQo0YVl/k8Ef+xk
Hp0s/InllGs2W8/ZggfZyzcO3PmHEh11Rq+FUS/pA3OitGtaaIoJZmdXqr+/EpbK
TDY3Dwj39PaMumHWrZJoZbwlXG4AHUh4A3lN2vtC1Mf8b+TSrf2t6IKPPxidF6dn
yFV6w4uTMK/drvakSWUooRViN3RU/oHtreoI2IFkgQYb58AMh129qTEidGHUvtig
Nrk5JHUg5W5ewv9W9049mVVz+zvIBwOwV8ehFIfD3anuGfMSBRdHHxIg9t4Qf+5G
vvPxt5lG7Zyk+zsGJp/jssQxZf2nkOBrAFN6uxN5KcKqQdDdshfDJxw24pWlJrJA
8iQD90+85rDtZPWzuoJEQhMNkS4T1SF9jv6CQT61CcYreaF8ykRYJw9fCVNN1izT
FsXItHaQBl+HfaxEseRHw9GEHSY/EajWHBheHnKFZdYHj/bbWntSXsS15U6nRd58
oRE1Pl3u/A74+XgvpDoYegiAbv2EvXaionNO0Vmw+l1RbWwQw+awCJheM5A/XU83
dnS8zNiPR1QsA42vBEi+wNNUAMgNVLt6jWwuVqHwfo4byFXjYvs5AJ4FxsOZ+Myp
dxJVnRb/IawmTWA3WtemqPfFibvHDvQcLx9ZXh39pVwql5WW+BmqQ2a+S36X3Dei
8ai51KHffsVf0pztCooj8KG3/EGwsBTBGbO/MTirE3dPFBzf2RSVexyuhMLfhw2y
d4qRVd1Yw19vAlOVhBBPevSLQTLhugQ7N3sCLglvuhL+CzMBiDcsKkNu5nYjYjPz
VwMnR42DuTK4dOQbByutj1ijlzFuFslOttmZJZezgwnsjljGODKHUOrQ0SUkOB+r
lSEoKqCCItpcsN+7uUFYmgT7+bAVlgiEop72d5fimhSWAggnG9Ykan/WUkivgB0w
m27WBg6EtLKp5tFKGTyFlX38CU9ADj/H/4cBQPyuhtBxM4sisvO7zLzO+WbNCjs0
KUxA/9o3POwydO5YAs7K6AE5h1Pkmhlc0l6hPanz7zmlxGRoXEiBnrK8T2Qqn0Fw
nK8GKUxTbUTGNLLXwon3X6C3cVCEGl6veMpX9jQs4ZwkgVWIOMNDLzuJxOUe0Z73
8dEbuQ/XdtVmNeqvw9yzGyWWG2tjvGr8bjOnyiOKef0L5PDrK7pY1A74z8cbNNqn
rJQ9HtZBa63455Q68VlK0m3/FyBBnsihPL7lskZxDLbDuaS6lQLmQefjvhSXpaPU
WHtekf15ngOiR2mW5Z9pHH/ka4ih+LPwNVOaxzBEQfgjkQrVIxxwGWiGB22MvGl6
iQPlPpsWMbcMWghPdkw06Q8D5ZFe6i2Qm1z8TFbm5kOiR24Q6TEgIqe9VHq0TYSs
2hbF4s7m7HDY06cowWtRZ5Xe+zQi5D8hyAxuAuxHm32TAeGGSlb5VE6UcB5OFP4X
k4/1PqCN6D71xABUQW+tExoqUAOYHjKecKjThmgs0lbTI6h6vp/qIvJyyJkS1SPM
KiiRcEknIu0osHAcfWi8Qt2cUisZ+GVoRCG30FJYoV9RIETvY673dgcI201qsE7b
mPm7nBdYJT6xZHGX1GMNTg0U6bkVI4j478vPUbhkovq7aH4B9tT1RmAzwqHXEU9m
qreUp/3ZPg6LX2EwaCWZSbhnqFNa8vTrEF/HwcZn7spQee75va3UIC4LfWhiqNyH
gAl33w2y+5zxlADlCFyUosUhVbszzI0C/WLDv31zHdcFZ32lOMswMbpXnAfnw7oa
AM40Y0W7mVGkzPFPTk/lDBzGNe7QYkdnEBi5QguV10Hau2Z4Qvta7pE70yray0SJ
9Bg3FBPpTkiv6lmOKIbML9h4eErsnWbQPhSm7cc2ln47UiX0iuOsxal94sa6z5rl
PYSL7x894b9Ug/V5Ix8rm0fqdNfs1Vz02s16cO1TLcTttlkEtyGzrb5SoF/QkOUw
4J618Rw4EFrCgpeSfMxiy+2+C5/ePwhxuWGayC9Xp63W54AcdHyrmvTgb23Rn2lb
UGkwmFCYmmAZyUEzqpfLgSYwJcsu8mkMObLP31VQ6jraPHAJGqXjUvysxjjuKK6B
N60P4/t6W/P6y3jsUaS+Hn+Vt8E/KNIOo4sxLqNzFRdSyUR+Dawg2o3zsf3+k9Sc
6BralCU+czDzSsaXDZrKiJdpVqYPFmc+rUSruIS0N5G/oTlZorKefaEyBlHJCJJo
GlLGDjundH3Yx3NbTIVhEJQ30rMO5JNAE2GUipVRjhs0KP5tpqSyJ7jBHtBt7UyB
5f0oBThmhlXN7VC1w42Z2l5FCwwaUTrj0dA2X6/umMJmw7WYbOQvfFc9wk9gq8L4
lNdNitlLqC9FHrsxfffVRvaQ8Lsrs2cCNH0jHPZ3L/1in52resVrdMf3F5DdF6Eu
RHvCi7szVS7/jBPHMZK7ZEr6nzspkSrcGTzCbNocQthpS8+UvhDrz51VyOy3a+4/
D6M58ap7JeAuyqsT027JTO0c/ZR+/LdSDhHyzRu8xbiimo7KX/yBpiP9YntkNnWs
80NqsS/sMM4BM+rXH5OZ2W0Ap/q2UJx/OCkrQGnU3ZMx5S4+dUH2C7HdXvZ5qhYC
eLqBxCERjxCEchPXIKXqFaTJnwHwKcOS1xaJk/6kodYB4oF2+lDuiQiB773SSjNY
vGtTYU8vo15IxIAhvNSGz0Btp3BczaiMVNJz4whePSpn+LXvNESfXkHMBf6E20qW
blkVerjNGE6yXQEYHni5ciS/l6Oj/CnQD3FoeFSUjHuyeOdEV22i8LRvwOQ3iRd/
E8kEJ2XXM3bPDUs63/NFvS19tj+Kit4fvzSfemi3ktdVc8DVQQRllQiB6EjLqRy2
52O5Z0428Y1FI1XKQk6ADY+Ya8JHlXhTd8mjLDRtf+Re6DP/7g7CHds5n2mm6jXd
s+a3+zzhgUGZSCXts/IqU36kBbuapO08YoRnmTBXi/eD9iqrsQmL/U2aUMNxSz1z
fj1tUgQFcwS2DeVk8FwFDr74R1q2Uz+3lvM+06mklkpXky1gw8cshr6T33TYEKzm
ZiuottPBTooSVj1L0Yp4X2VwxH9ELGDfuy11Uj2A3qDBuvlOI48ZP40ACBv2DMx6
eGiUshGYydfgNzpVBgaWOBYQVLRsMwrtKDH6bF5KQAVshfv5k4RC4TwqzGZEsO+3
6TqlSvuk3NOfuna1bw6QDjAzBTb9kBgAfeHr+W1y1A81EbU3EVYTRZbjy9eAWIaH
Pw5NikO17cBEf1V5e1Pb53T9lasK8nBcil7Jj6imbJTR0HUpuwFWENhN4AaTXCC7
I81RGYskj26fqgkohqPrtzTgp66cEw0GmCkotQsyzq4W+uw9PTND3OAq0Es3kSgn
UCSdegF1do52+CKkZ1MYVKLK0H03VuKYUPt6HdHxmNRVK8ZXSCNbhMwOeWeJsCV4
qkXE0B1ZSmsVww2YFDkN60CqvDN3qgVQvlrm8XlEr0ldHR+GPiVXIOIFG1ceu6oj
M59MmSflZMmFaWat2Uy/BFgwQiviK08JOS41AKT6SKo120+MWWM5eZl08F7mOnVz
gieGzVsxN4LSi1n/ZeiZDx/Ee59tBJcg+fhZnPvGmOeAXEgtAaYoxO+lp+oBDjIU
KoDY0M2B3Vuziv1BZ9P9/hC2INIqcF06F9nKSpRlQDFDIQsbLSy2nUY6WgNNLCUf
izbu1paTvgT8w+j9CAj5eu1gb4L4N/MZN5pZHyKsIEsoXdZWfFvbuhC6WRzaL0dK
QMCOKprcA0mwkGU5cnYrIptaQ6oN1a83mlvDS6HP1sAt51AQUday9cFuR8xWFEHS
AsRJEq/OIBy4Bm4HI9gOumqWlatTjFwP/lDY40m/tifRM5RUjxJOmrJULabOjCsO
wesjAZ/mCOIUc2pvw80KE4OAVe85d/1PuJ4Kr6A0Aw+WlGMkl12exQUhd4KWoPwJ
BlK6SKQPGeQFcv1+Xfxd+3PIRa9yCSv0PgUuMkl4iygg4h6pR0se8UKy5vAZvp2C
iamvSgJuH7Z3vdtMojAHCvrtJcEeTG1gxR8S8SHC3SmU+RRmZ0xvoMVPGnSEB0e3
zdjg1jGj5Ky/fCZBvv0VIjoSxxZ+0gu/RMm3CAbYXTZKF3+fu2TyglF/g+YzlTbc
9sS5yedo72DnlMkESLx2DF/odG6F+P3RHrUj7QFZP0eEqEpWPz7D/6YLFzeXT7fg
7jR15DOzyAjl2U/hslYalfrfyIXLpIz4ejJcgd0X0nXv6XTdBzoDxrTTPwwG+FeD
qg+BNO9g8oqMK3jHGwIiZGtz2DNMNeuUOZPl9WwcquSaN7scqUUIQqwPE58CWwkw
xhLm5JzTmvghnls1HPx6a4F3UhVtXeBkx1PKAsZfK99Bo59IVlytVNhOjL3LoG3t
VniXJfVPngCq2QHzh6a20xvY5Rx6mIWz7jlxGoDZvLZGGzBoiAfRxi2sOCMLlPbU
jh7QHkc9+2TJJT8JmtnY+PycMETLvEztzIpjVwmRup2C+DNrZb3sKDP7wMTzdepe
XghiaTDH/0VD3CIkwesy/BGw3dpBsIcXFvNmJ2IJI0ud0dGxRQbtnkcusoq+xFBj
ag9ccYs04WPBZzK7a6cO9TNz4zEa9gfNHLOxqNcITTtU8g1RhOtOErhJ0ZHdQ+xz
0EPmSs5CurGmYUq/d51KF3BoERsQW13rDPOq6RXFZqt10WxvT1Q4iJAV/MS8b/cz
oAhCp/eO/6eO9qRT8hI+8+IftFkMKp2o13zgv7gQ3clR9htvmyK5jHjLBIe6bo3/
C+qDJEhpcRjKpgjBA17QjPShUFRxfvCq5epCOFJyCXE4zhs6llLR6qinwBrvE75X
v33ejdrNaXCM3r1JWyxRnpla9tOS6N5PrgRM2UdsbMa2ERLUL+eh8g8u8/sbBiIb
LIev8Zl7C+hlQND4kMsuH8n/naEP70o4Mb+37ik0VT7udAfLGttuUeWvt/C3W0/a
8h11wEn3FJKFDXjujQedYH7KZ7PBwj+GX5Fn5KQea5xaLYzeYoGRt08GmXjFHHv4
xuctKla44btshKTx1itUhnYcg6lqvpT56cDFtqO2ZbSjLKD+RaIOOMfoUXX+rby8
GWegDaxGr7OYOmwD+Y5z1fypG4NOMNsgdPxL7+FnFB8UWJEKb/rO5WihHwmAJMTa
vSuo1GO1J54MSuO12RPPkplPnSIu+MQAIGctAPgVibvoNNJh6PwnYWs0dln1GMm1
wfxj5GNw9Au9BLI3/NQoHBCIQmE/JWA26vcnn40/qL0n/vaqgUsoFR6FEBD0ffc+
VBTtqa7NI82Abm0afyRG64Y+8FghYS9Bmd4arOoBMr5fbunDUm+rit+0ajW81LU9
15biMuufz8btfEG6i9FIYdZwIxGV8lXDxYI8UM3PI1NpU24ePyh20Zg9lzWjPki+
KfWOwStL3gkBVI6F7AZUWIPvE+Gxg9tRn872OxZW9/MAhn6yaSTVWnT4N54mA64l
`protect END_PROTECTED
