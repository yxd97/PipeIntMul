`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
acfOn7q+vJ9bVh/L20ZT71gBh6nDF37rM1wwMcNcuAxH58oDYGW7B1kNE0yU0TmM
Eqx5QmVO+trCVCruHZHDp4sfgs57eB6vcI/4tX53CIJDP+4axb0g6lL8RtS0fDDV
H5MM+pt8+GaXF9UUVsTAOTxXhZdSSKmvOl4SqJD8GxPyyz3/29Hbk40cYBdr+2+Z
/fGZ/rsEwBsEw3PhP8lx8milOnmZoP6tByz/t4d3TzkcuTI7a6qAtpI/dfi1rRjO
TuOewY6JwUtkrcbe3Qk1Kj0btrC7H3SwdcQp2Wazr1Br4aPgdIAimR2kj35yqTRX
MRMPSz2lWgGpnUXWa0TrXjsEWzQCeSPjH/Rb6vMKIl4KKP11YpIRSHcCBcwa/OJ1
5b+GD1ecJRj9b22YjjspNw2zG0c1jn4S0dCks4YC+/fZ2Bm6rX6KipxR6nCLx3yy
q+nbVju3griccXCxxn2YClWiFdrnFfjZAuOpLgQ/pEzEc+g2zaCXGJ6ayq1XmV5b
PZqz5U5BxE+nY3wbT50c9Tf+ushdkA3MLuETyfiUKr9vuKPaUCFDZ4z2pytZbD9t
r3WOEpzOdsBbDol8Hbu8VYn9Fg0fL00KMQFivc275Z90RnvjDIdIGSk77rd8M9EI
tOA03nEB/lvoXw8N0XqspnWt+JFnypxS4JCTIuu/Pjwxp6QvrXu6FDkPT+vcxacy
OMSfEiskZlBACpThFqvT1G3BmDJ3IN8ACZemX58wWF/Icuk2cAXRgU+2m5OcFXbn
W1PZkJqkrLhLL1YPGAVG1w==
`protect END_PROTECTED
