`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lTdUaklTfCeJdIzvfSejTkd69J3W0hCSp97YgPmgw3JkqLQG4c/VLGw2d7xX8Oj9
Nt+QxSI6OrSeFybUCQL4X9SCxgjVHx1GQk/BFazIiGaRK5738H0E5onQTyWpA3K1
9RXTF9FdcnTgmhjgHc5RaBW1atAQPWFjouUMMK7mVsMccsodnr2TbS1DqmeM9HEi
W3gFjZeUK94Fn7p0BODJY+QEW5DUrMwn9lGNWvq90F7K8A12+M2uKB0VumNB7t/o
9S7T1qyFiETzptCwqJdgdnF3IdFLWSuD8OswhtKLoErljfVaYqT0K9KnSOsRSgPq
gzUHW6Dm4v39bjV0LLlh1PAdZwZQGDBVYm7IWM21fH8FUt1YtzShG0nJE7YrmO2R
yE4OojVM5/ZP0ZFsb1h1B1p8sU3LGj5uHv209VKJlVljrjrHjv9hj4VMPHspoMdQ
uBz5TfNWgrd4zOF/dXY7rEi26NAJ4porKMafOV9lIMeDAEMiQ9VMhOQ1GVDt5HhO
q5KYh4oCvffueUS9Kbk6hE4TJkSgqAnZ9Sjnd7UeGR3QF9MUYy05xyAQkBXVnqUl
3cB3UPyinYwRyBPBWeFNPL/ubJKV9uC+kvOeG5SBjKN7+uguNaSzDWGaCskw2gpg
djG8jaT7Xceh33AtFYJfz7THw5+NAZR/SrwazdlOUB2okEMPGiDC0maeBfzf/Rqa
zGVfLrlSxv6+q07xnzEp+rrEn7UCYkTdlilzyyA2eIEeBjBxWGW8OZCfp8MHgDN8
xUbCSnjzd3l8okf52PFDc0NyKkxwaHJj7tCRSeu9YNTeNELUWuFnuUuy2VUMal1K
vYULCp6dTYi3zQqTPn61vJJJX/ma2BBylXBuXup0NolYHWmG/j/53ANEhnqhNZ6E
mmAoZWuFEmZnmYsJVhmiVZskNPPbFc21twEBub1Y8sJlAGKWPQ5UNyWS1NP0rxNy
nT+L7AX+Glg/+ZX3m7wA4bcBAESCK8aeWR6nKt9U3skRtaxmXZ+bdGeOp69wY3iW
kzCKcMM0aUC8dYt0LDum1iKLi424t26dEE7m7YWCEIMFFa7tE+Me6f2DxKeXxAyZ
V0eaTcHV9Mq82vMfBPYpBPphaxnY4CtRTD85dpNMKawz9W7I8sU6QXtES/tu6GFg
0QfOv4TyA9pzUQ6A249snD5RyrQBWZ/1iquXvbqrE/Tj8kDefKfDlMOzOi+20hYY
oLdnLw8uJ+kRuii2Z/CxWzlQuCMhSd6jqwLC4M0adARtraTKKxB58AKwUDg6xheM
61YQJVGGRvS2SGu4oCG77EI/Eje1ZCHkPEbQR6PbOj4ZwLVk3Oo2/fSDrSPU6ZAC
2U/dfyEwv0QLjGzRI0JKIjvVquviLNCMAC1LUtw5fwMWPxVHMrbJA4GYd7gjQgiR
5yKaxU14QQW3zdf6sIadjLe7KT+tXeYW13IQ7IwfIq64XpS2HC7zG7kTEs5OqfV1
iHQT8UR0nmo4dSFKVckmxogJI9G0gZFvvdXSNNAFejct9WgGecouC7TuAqPtE5ci
wpUF4z7Zf1lElFchCdlHfiwptzXmpSAdieDWfu99WCDKkZdEuiUc4rwWFsN7c/Z0
w87XWD+DULx3pgDL5GLn/eptLI6uR2NNKTgOU3z78ppmcd++cANz30P2gu2hnwyo
ZekCOmnERHN/csBVyJ3i/VnOcG7dZWuXT5ykEExL+NMQkFPfcOjeWoxotknAaSbH
SFVDsxFAavnSrP4zoYAkkCjlxcJiaaHVQiBCiRx1DmTbQWajlMCsU1FtMLoLgv2A
lvNmX4llrfTw3PwqKy5EGc8k7RcyfASWmzMOJCcHqhh26HiK35zI57lrPntp0ejV
hwPzkZODIzNehWsfrTpWl1FzD3LW7bVmgtGUcZOz+PSCm2BWRfSl9JIKOhOhN5Rt
ck0rL0QPvSCAXvPJ6F+tyXjUTYNXx9ffsmnJkuNzuiIrr0ZaAWkZvdmZufgpBXq8
cuMiZ9Rk2tx29tyaJw7fik+CGOytCzxXTs0oAoXPELM3A00P2+Vd+FOdOK33sAux
fbmRJopuybSc/p07ZRTOrbkS8w4336Ero4hXcBQOie7orGoZsyydXgJ0/MeybLp8
9rmfheW2afJT0OAwO6oE1ysWO7yMef8T5wLzlVdQ4qxx1+KONZGPrQs05mB6pIoZ
vTgZEBfP4d7na2lIJF3XPS5L81gs9FwGfJWtaSTe1AL82W71Yx00mTXXIEZhM6yG
YBGgr1xudAwnD9RYhrjTTC0IqQUm3qVto9lUfigyVqIeXtcWSn8tETFaSEUtiAP7
kdXGxFKzE6IhHHoXS8/UiTWsqFA0dFwKjfbJnTdsgiF5i87wsZ2bePs30OKaj4hU
cYHJWAJI7VWYoJtcv22YHlFZNNszB+C6wSEf5sm9V4tW9szI30EGHEcvnJJvWyxi
Hq5xZEmcg653m/RkGQMz0kVsdV3LHN+lLArKM77pdnb/Es/z+08AHm8mV4/W0Kyp
4alQYHqzDAkrB73e2SpSyvBLAPXc9YumKXhDOCDYyOWqEYEGK9mw0U63BVKjPM6d
J73O9S0mkOgPHjjZhrpuQCk0kBsRTwg0pf2rOMZ4cM+dr3vZLUd6AXAQ8cjllNTl
tGKEFHiUsf8ug8t5I0AtztlOPLQdX6Cpl4Ywm1/kfOLJVLuQHtmZ4BH3BwBu3lcH
9EJynNBf++wDqiswF9dT2TDBy/K9ai7FxNMfq3zN4rPqQC2DWTvM3+MkP11DPdbo
lM6+wIr8325llsuMP3vH+LsdGtMoU6I05R6om6ARKvN/hOZxL8dnEWfNYDE1vFQr
egzwOnMA7lryS6HB0eE9bJnF6EmigRyRP/L2vJXHToqADqyas38fIIN+XzMnxyPe
ovHKnyKwQ9cd0jLRh4effHcZ7PDmARMjKxwSHzX/bT83CzvB97g1ENWwgpo+Zpd6
dIBfsLD/njSdiB5AYz2hibrhzvwiBbtRwXuApXMt4WMD0LYXUOLS8rPgUDjklu34
mxzHZzXkTMUiRm0Kp+jFuXaGGyHiv2Hfz/2YAHMmnQ0UEIqrPZcw9h1zjppDrG5M
/kGANobtZxiq3vYkVhyjpjhV+5kN2S+ExpKPXoAVLYwJOa4fyF/4ZMa+cJLDwtES
jTcEf+CbbQlVS5Isx5kZpx9oYBdZakvQbIYmCW4S+u2QATgQ/uPoZJbLFDPls8/e
SQFKYX1SamCzkkl/8Sw9oDn6dhs94dk6Q1G/3syPl/VnQTMQFlzeyW76ehqeSkps
yqTckkSoqLWd3YJVnu/DswZP1IqXk4nS+Gh16w1cE5FrQFeEBqn87M9Iw6uLHNfh
fIbD9eEmGB5fY9+ico+4SvqBuhpE+QSrK9qvqHCQB9pAgS/qWRpy4BDJP9GwYzy2
u2pHHPyYQJyPpnctChpwV9HUryIoON90v9U2o5JamHpaIBs1rrXcoG95557OkUmL
m9HwdBG392EAgYm7NJgZgl4KJVkVz83+Ua2CoQmDGWRZxRkrU0kDvf2mYXgpyOUF
oCyMz2Vq4D9Gm0ovuzED2gxA64YGsTzdnbleIF8WQv0wThgnpbSesjqY/UvuC3p6
X8uVVzkemzXGKrW0rfXFRAMgRWVhmtL5VibCfk5hou4kXtFn4j0sNqN7KuLlTwMt
Zm9Eh2sF+tkCfp7YwqBJgHY22lK+pa3e9qQi5GdyPfzLCk8HgihLYq6XsuDuOTsp
2nV04p+KBg1IZeegnXwck7YKYQOF5EPARD2xONCc4QZNrsqVWX0kf8OPPYbsfGbs
kj92Pr7gvS7fby0XaXtvDAabYWGD07LzrL3NKpDcrZ4ILpe/rX7KdHjPPVUUj1Qc
qLSGhY882ipJKy7BQDOhNkG+fZ5+hC2eijgfStrWTiAt/vO0ysrdPKuVZ2RmCtR5
+Pvg/4ayrZpatP1yKFYBfWow1fuDJ/8k1KBxxKmOo809ODwpZPFRsYpt1O+HOBcT
dWtLDL67pV/3HF43RLPLbIc9TynXHHCVG+ALKd4f4+U/m0hYpBVgbvjsgpweDUBj
xisiXSj9V1Z7k5wTbSjxmlplJMbh11EUap8iWrbIqpEkOkwgLBjW5bRXPfY7IfNh
Lk3TqJ8Mm2nDO88r8lxydKPNp3OaI3rM/EkDQuADk2Qe9raFTVys5m8s9BSuAfOQ
1zOwIl28HjijLhmjXdWfMgB5aPo4wrAgTW55IexeJuelRdYiQ0Li+ba+GAAiIyLl
dweFbFjgGgpPiaqCpS4eyQ==
`protect END_PROTECTED
