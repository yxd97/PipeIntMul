`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4Zc0Oqt0wogwgr9B9akd/bSvIYkAle94Q3MJowq1FMl91UcDdqAT67BTQou2SHTq
5ghcIIuJtR05ZYwBmodCuSDbih5xeJUdLmDtR51Tm49l8DEw7iDv70WaNUBz5ZoS
cSSN20omxMatwvBS/+tHA8q3Ooive6YBaPUY9CO0j2mlaoa6QeaJr1Y80zaLc5NQ
Gz7FI003X0uNBLBamCWWpMzwI+J331QXbWeL4/2j1yxz9R/jLzKmuPcjv7q7UZvF
bs1b7MK/LV3/oxBMkthkduxb10Llp9OfkYlsz7ZDsYZREOH8B3od5Wk/dPizFdVX
n5ucUyR1+DJzk/16gPsQloJeVJrv5lmO9Ixl784KifAnr7Cld2iT8YKi1lH/1DS9
gCsJzsW9q3eAA4K2m6C/nKTP0w6tJzbtUL9kKuoPjV/BdGD8vn0IBgzWXHTP3DmH
006PG3R4QLngRhYgRWIV7BZkA1ZbhHzb1n1fcr8xHBHmehikZOfGXIENhzCyEk6d
`protect END_PROTECTED
