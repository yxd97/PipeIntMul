`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PLrNNbNRHMVo4Fjj3aj8mk+WkeMzOSY/FAtvoE+oupgDYzvGdvuWTrsW+8HoNNtz
UqfQ42zcTQyvkTMizTpO1CwZwZOuGgxL+F8A3HjFxsYmkSTCHY1X367zraoWQNR0
S9iOLuCI67BOmztABSFZj1um5T1Gm10JxjEcGQOgYZ6fFbBoPabf871b+95NvZe7
SN+qcW0l5jlcne3bFjMYjVKwu3sURnqLOslqbjYm6Yrs9G+a+GflJeBAqeOs9bt9
zoLOTT/2NklxVFuQ9pkTDyra7fkSvDpbd6IG7cNBcftBrnsIS6tDLJRGXj5e6gol
KRsblwkiuddxia9X9z2OghInInywhHPAyUuye3bN5uZQIkGq7zS2Ro1plS3N56sa
H003H1+tSH0mwijBvy+APFZEUrvoRmiXI6QkXhlvdcrkOch3vOM99JmmtE0H1IUO
kuAV1AgWC8AK8FQzL2xThDib6aaWAqOhjRRR/SHmI/gbj2W3o4/p67c0ae3V3Y4z
b0sKB7qEF2iqBz8Nc5AbWe8xu9BspghGJjodUIY9CbUjX8mvNvOtalWXdcL0mFJd
6ubsKZrPOdt+KNuwUNOVoDfyL8TZltcVmpbAWhmXU/bBqrM5xzUGIbnfk6I1rCKN
Y4dYSKFdTSebYyS9f4YDayynnt7LT08JjoKdDmHz0n3BZI1eSR6+zymoKseYsJ2X
jBlTOOfr2LZvOTIHi74PnffguyvV+J9Jnw3V3jKk59itmauRLQAomoeUXtvjAiZ6
9K/MTYKYFdfIiO1e1cSWd+Gnyn0A9Vb5+gBohAio7aVxVjMKa0DD/l35X2SnE8QL
HxSIfc8A4GvQz+1H+2T219+ZGbQzkfcBO3cGgdotF4K8n2j5cGwquqtKNaCb2MCp
dPmBMnr/nXscNOVH47KiQzUAsVVaH6HDQK3BhYMdPUTDwQj6hYYFT49i9pXNsoCR
UIXQEn/p4LRlLLZ+iHjBB9Ba9nm8NN/PaGyjYdmBs6JC8RZduXa6tO9tzRFiiuzp
4NEj01h/zQLDX4N76KWRewqG4v+H2AvquRPexPCPuQs49G6XL0HORjqPIykNsYBD
2QA4RrvTFS4CXcmt/xzRLttdkUzcZDZz3DVxWG/kFp/ZK/8YGy7DsiTV3Z/iPVAw
GftvpSbfy52aK8ShWjeEzhr+iRqWFS7iDS74CIO8S96+N/KJRT7Y7kwH1Bm1wiV3
23rbg9shotwlLrQGr4A1XynfTUHQqnIgHQrT8tCeOIYOHhR9vZiv/1XpPYjKprKT
6FXZZzBIrA4R8o/QYsQaARime3YoMBy08NRrPB+jvLU8NrarOEuYYeX/dJqvQsvw
ts8JuNIlVS3X1+b7xm/GzrX1148SAOYEXu1E0ilnNijorJNf8R1zb7s4EuY0R8JF
/x0/lsbJcWh6mUyJpKSMhNMenki6CK9rPSQ4AxmUK8T0uEzMETqM79xfG2H+lFcH
qD9I4LQhwPMb/d5hn6J3t0WuEEeRLS9BzX1tvmewdHIWCP6KwC60BKCTdDWg7y24
oZl0+OD+1Yfr3vXEcOIKkFLV+t2S6Dy4wNBIo0bzw6hek3uYWIQLF6TxOVqlk8uN
aQ1qkkSV5wdgsCfUDnIabHoVaDjDTWgka4s0hSmXXneTuhSacQgP7517NhvvUGZ+
4m5YQ0lw7SrHjb1PbijJpgFiUqARNzghH2ZvIw22QSrkGiQFREmfrJeJ2j0+MsoA
JCxLYepXN1TAd5gRuTXKEuFjlYanT+qCNCmOnwOhQw6phH5JGABKNEBI25exCbJD
k7YENuSyG7ANiVS270efu336ZufOE+GCLYiI6S7Dw4h0POKzfbHuXaqy2o9pAFGe
LFfww4dWKZb2SSCDbcYDn7/E+TzzZPKR6BaSohYpdPSUg2Ep2GgvFCSRMbAwwfx2
V5FxUmffA8J4gFC8VWcX5zaRS1hqyA9Nyg0dD+iULL3zx21eLnA0tQOOf5cYgArv
OOCCL21w4KI4WM8OVgLReuDBx7AdxFJMvbq3BWz24AsVxGhTrV6Zj0cJB8vYK33c
QreGgM44Wte3VJPnL/jZ99lh5Lpaz7TPpPMITlwhEp0zvmVDzCC9pXxvZlAwomhV
KUAYDVxU2kQ44fiqTW3IyNrBxwt5eHqyNQ6F0lueKlpC4ZY4ilLqQTtJrfZNNjf+
76RRQd1nSXmJOrcscprgN5MEi4WoP8hVwWKwpHBgykFRljyhHOZrK6d07H1m4dgm
rjBdVzONbmgOsuQ3jZhCCIrUWGUDqnbPBfcDiQRDwbkDsAStWswsFNnXYLxOojHN
KX8Upqo1tPl78kkBDEgaK51MsDpZQpj4dGHYrH0WnS5NlyXilOx/y5fc5ysX7lZo
6no+5kb5Y96PJdC/n4t9E30I+7uY1xpkFwCHoX8uQE2dRbHc3s659DmZLAgM09ez
hLQY/AEIpEoNzFLZXTP1wRk/uS9B2cFOPTo/tCK7nZEkise4R/0FeNDSqry3uNhV
Hf/9Rd+WFHTFeuRmF8w6Jo37+HTtBC0LeliCp4xcaNPcWzUnNoMS1YU11bjEboeP
9alYloLCogX849Flo0sT422p9xqAPijdPm9zuQxVziZuMEVrWacXQelEq+xaAuI2
jz1VxIxCCiCJmgnwl/AB2SXwdIebbHyYMET+UF7b5B00qLsmo81B+Dl0/Q+TtWX6
RjxYkBDvQexjzBUPOkaI3dcTqba+CHSsvLWwV28hi6vpa1eQZ0UpPWthdXmEzvLo
UFYARkQDF7X6jhAzVcXr2kCz4NRZVna67wXtYM5K16iA2AHnrILXcbBuy6nv6NNu
vG6/K75Fi30drmWvUEXszaXK5Z/P3RQmtiKCw0cIUCsxKtt0IydpBHV1bKBbGSke
tw5IHoahUNFZAUba6ntZnISjmma70dWH8nk3TLhhfFaLsGp1i+igg5bU0FdqgBmm
25rrXo3e1/g9mCwrf/RJChZtiX3Cb2ow25a5LcpulcDOD5d/rQYdM18+9q4A2N+i
hK8U4TXREsKjbheSN+sig8Ary3qL9mdliKzzkw0uK275a6NpaqrWvSLhwOMgzicq
H7n2RJAOk1kwafJEedQ8stnC1OU2QmPdiGyLO34HhpRUrLT2I+onfne1OgQMiX1n
9HldWc3M47bAsFIE8C8TkKmLsppZICFSw3H4VPSA9HuoAL2ZAT4wfA+N77ANFOXb
Q84q+82oJrcDp4ydWiSVj4tFopzliDdjjMHPxcK5AxHu8IBO2Si2aN7d2FLSbYK8
HIR9MQdwO19KeiP3Jk6801UbqGDNZjIx/5zDVU4NB95FC/Fq2+aJ+7YJ7D4iktd0
5d1DBgJudYeDYWFiaIAn8J+WvIlvOrgqenjdeMa0o+tjqHP8LedPE1fIykrmteNZ
gHlWSmQQ00X5ghBXKMZUMVsyshlT65Q9hoCHiVnlN/4phz3FxHkOiD3BZAx44o70
HQ3Ep4JpVijHyuq36Gj+XF0d6Y2C+EnPIHFx2w05xAoZQ0qzshxi/jQdIDRz4zk+
putkpX3bx/EJaJiFPhzH+PXOq2FpcDt27rcH5OorMu+6nTN4l+cYmBW4SxnwTU5X
vLxoGlGCSHHQz/z+7NLTPnNtYMjQkVT8np9Yg+7CMsJbGaO0ZWaL5mbPzVSyqRKQ
vUJVHm2ef6J7vhheEyMQToo5hIB1i6cspVdKqlgg+7Rrw7i5obN5+FHDc7r+O8eF
MGXtfkVmmtXMt+CQYNHcq5WpIhd7jXCI1DZWeWFxyzCsvFuPa38kXRJWjTqj4HKg
cRe/n8UtM+OjS676hXvHwGIb2u8tV1lqF7W6ZRZ3ZQwWaYbIvnLmFBOzgAzXmagE
uvQjKMtEj+tnSHjnwPqL2ZHOpsEjV3oT/OrxVdgYsDFBHByv/0wgBuKuR3Fd4ZrC
xX9hICjUENL3T+Rr+ma0WcPmI/jtoXonIY4oTEWolJRJZ/ty4Oh/MBpOL+B07QDY
Fg9rPAiB8RzHgvCT+7fbAKUBXqL5O3Sb2EJt1Yf3qe7XSTkKbbHX3ESeeSCx6l1C
pAl2+t1YWWmFJllF2hvWFVEuAC0rVcIjUYWJJoYGgqogSHoM5/qdlTx7HC+6+EdX
CT3oWWlCNhc04ZYUJkbTfNCJ8CH1XJRltc3uAVANXpKhzlfDcSusCmv/WTdt86gv
F6+5pU1J149fWsZe6O2vl2e+GwSF77p++OtXYXJso6IuzgbMoLkAnpRFS5fQdEm3
tUwOLCTXXyBMnQefo4zI1g9uKtHG17t9eigxeRHS8wf5GpeVt+GuNtvlgXZ+fZxj
rNn4i+bnXRs/h7mqlFVuxzeH4qjGZnjsv1Rs4XMn0Yfasset8DrZBmEVn+21Uxua
3UxGSclyk+B1cN0GAluOsmPBtbRiKoWlyQcDIBNS9K0DtV4TDSd7nBmXfVX0TSIl
`protect END_PROTECTED
