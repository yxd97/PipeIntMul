`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+PG87JT44iheNFT3q4y3ztNpnv3fZ3OAekRylgyHvbaNKbHEw81m+nEPkAKiDjoW
RXgG7/o+zQqDk0H2aXmFQ1u1Gvai/PKbv056rwyycYdr3roUaeTIyWW0WUyPobzT
2/JqBjqNRlWiERkTLlOihkSSCW2tusUyFkd4P5q9qkipLdW6HjemxyYyyc8mg4a/
6P01QDrNSZtQFsD1zQAy4BoCZmdXNDOQ7S0vYPD9ix+IzjeDrM6Xy7y/2tBJfEDD
DfqftSwj7C/7VQVFrSljIqE2hP8ojk8LEYUPZKmVCQ84daj+39YsJ+lOyxD8jlfk
AjWOS3mrj5Uod9dLaCM6tAUeKawrtn10FX2+yhE/HbBzeTjuwnHx8zxHVz/qICoU
Rr9ORIVOzyzM/riAVNXH3v2FdA70dAbMZhSoHF4aDmDNxlonVxw64elvSCRb9dWL
wmk4Ny8lEpZj+N0AXxJ58HBrQE1xVOxLbRtNtojuTW5IX9OI+whX6qbT2rP3C3au
+33OokOT/Tz3i1C8KQ/RvjtZSm0wvbWtuA4pgu47kB4AN05YuxGN5EDOGigH9heo
lpkOPtcH/Oyj2TnfuOTg9khrdfNOnUiAhnid7xl1+HrDWTfKxTqrHEqNt2n7AkEH
L4TKpMPlIEbNFkmH5be4E7bgxYZfwTwnSFlwvnJ4d+h/avZK4kRXrpMfG7XmIVc1
T2kGq+moPUeYXwpQd5HONQERM6Cb6SjNJSneLGhlhTXIz2zslmcp+A+VZ+qNEvHj
jv4gxb27ogFZxsSYbgW3l9OTqFfAayGa98uv57d4vlaAmCrPlzNNj1vkiGvBinJC
8hAvTBXXnNRBDO1AbRLYMsz4B1llc1NOMXdwLFbg+5yhn5iI7Nx4vkwfhXnPgE5H
jluQ+WE5DGg4AR4jpV7I4v/W3y/mju6QdnO5KSfWll8Vf8NvzaudCQHYUPYPMiAh
pJGfr3rIuNAsgvKsB9SahnwswVUr0quj9hyVAOzuAlkQ7ozbELDbRMem6c5t6YOg
GaF9X6QE6ZtGx5t306uwemjJw+uwEWpq98revSsABHYjBS04mkoqUEzup9X1gAnh
ftIpmcum7Qff+a1q8C3uixBJdBr2wcuscJh1rwthG25uIXSC5JKE3tGitZmVsm1H
Up2HX8ZxyefCegqIzSyIJ1237Wp82OzaKmCVV6c1A4kgOR+d8fvTXz5h9g1o0wR9
nSaFAs5Iad1bjOr68NhL4CojNoTf6fkLkGzHPehFUDuS8yuS3QU6UNvfb064SfPj
wdTJ1owtmEWiE3qUa7TS+ZW2JH/saa4RnMlwUEfRw81ZhtVAIs8J4qxulDIda2ym
W2pWeYiJxsUUP8cVZHqyTW+vcJSz9wDWZeOe8tXCpB/7IlzR08B7rlnzuMYL97lI
rdZ6llLBzQ1rbLfoVH3yiKj2Mn259PXQSISv2O4ES0wxPLRSvegs+dqrC5nxWt38
B+xF+NBLgeGRoQj1gX4uFigaswoie9klsSpz2Ak7UnJlesknR3fvOQC5+WnsJGkk
AseMvrQyMGHGVyjYQfxltFRE1Cd64E0rUtxqS9TKMZiKmp+eBmr98EX/f7ZLwvd4
/MDr4umg+XfLku3JDja1QfR81pUgoQYJumi3bfZLDyeTEFpfQthz+7O5kcMuvy8Y
VeqX7nv9/eNE/09Kp7RFt3BKtFHTDJutXfvpxq3yiZgcEm/YKICulRGcAiUTDS2E
k/OuE3vI6KsgewcOPfh4bJSAFXr29+pg+LrQXvnsA7naS7eNsmKkLmNB6S46v5qi
mT70FmoS3scxVh915AgEXt7Qo3GsCdLJnBUC1zPEurY1PPgxfsey4//aWcRkWZs5
8Ecn066XSirdHuRWbWRp1K1jhs97lgpqAaInxrWVm7/+xmE6C9f8QpxKWURThYc2
qpN3//5SWwQMNdHBFiAAqtgzdOHIbhObl1dRes/7zEA49Zocy++rUI5uPs3VdGg0
DLuFnHkjMLjZbdEcu6L3YofEbZBxDggDA1/CPkiZLkKSmtgL0+pL+QqV39LOtdPk
o9cklJYMw2BJXtzsQPgX5HgchPrkf+3D02pG0lvbrPBRH9QPS3b9lQJRRZfQtc0v
H6Wpco/aMxnHENHjXHzKHo2/nOCs2/mJBQRX+S19u1239nZPDlrWvJLK/6Wvw1N/
Sr7/K7pQAbZM5k28y0FbQJ32Mnda0lTlT7w7TN9/t5thRsl8eEIMyzRGFL0cnr6p
ufOcrig2hJAI9VfSIPhgVOkHWsClmhFsjHX5K6yQwvXWFaC8HdVBondXx4Geb+Vu
chSKJ5k1kRTodmhOzKo/+24FW9HQZqKF4o0zDXcJJhZuPHW/qTqdtkON+LJCI1Nt
ZRb1hYgX1r1lyF7ImtKfILsVwxB+7hzk8lsavEJ81IbTSNcWgatxtc1Q51/7G5WT
Kzeu1oiV0Kk/PLEtO8XaiQjd+L9ee5K1elURqH1qou8AbzjIZ5ToPt/0amGVdRnI
WZC3Ba1SHDWU4dpm74/9+JLfT3Kc0kokXf+el1sFSu2GDR6al5rZMO+6e3tg0UUN
DlZDX2lzAyGm+R1Oit8zqod7JkBfR8opt5/dZ+ROhCC8OnKuoRBqLwfhLKVTKe+C
rMVjsjj2nA3j6Y49C7rc9vtolfVz/7zrgOHZpeVsqeD0cap4v218OCou38i/bMKx
T1XYiTJkJ+V07PB3nGLBMpjQ4P6SVXQq3vBqLmx8ZJeW07rv9JxM12sILv1jTA9B
r7HJEYMNEUFyy68iyrpvSaUoOnerswww1zSeTeW/pOSkROTlUBBihJklf0DtgzRa
fr6P2MNxWqonp9k+SDUhuxtHZZbaq+rp05VcW6wtikiDnnmx0zAS5aWX5mMqAcdY
gFnpDaVeEJdR9WAxyzQyVvW4iJSdPhP8gFzwc7q0QSTLXuo5sFIsnJSg3GDpZzTi
O5dC23ccFuxm7HSpsN7txU+AthJPJkPLGeLDHKrfUsV2j1D2rZC1RotJwzXDb3KV
XzuNbW/hHgswcKtVs1Bc//jFEXpJVOT4O6yiTMDl1f7p6BDyhIuw3b5vHBOl+Sur
SQ3kUprfsX3lLErYdTAkQu0GB64gB7YH8gR8UHGxD4LNVUPyXBiV80X0839MInPR
V7mmnCmbnkgbVjVE/1JQrE4JVy+z4+dx8mURLEBIDT529R5b37sdWQsrtgSng+pO
sP/zjpPKFyPEluWzjfM4ga4gEzFLo9VIuHVyZZd3E+jMTMBmAI1xolFGM0JvsUf0
dRwojiib+1mqyfgIPotrRTDAsN1oclSkYubYedk2G7PXmc+Z50e+ZdWovNSEkUQ+
bXee0VTNFcqyx/j/33S09TZBAjvKqwQDuCnKokpLrDHQ7vUJzHb+rfXzXrYNQQVb
KCcdrgLIDgca559UUyUnahj/an6Udoak6GfblkBRZQRWB2b8VgZJZXJfLEsOoqGS
ou4zmQcBEbCRCMs13TmMaOoyp2y1V0TOQyKqrQnl8OHVyoZop3JkCZ2qTrOz3t97
d9v5IADH6+f+hE/d08u6Xdlvf+5Rr4/wX391gRd2v9pGncU7Q3rSb/Dah8E0ifCg
HtW/DQJ82vrIgOyQP2AcEsT97IO9NOLh6NKyF6FhwgVHBS4ryG0q0SofzuzLDVfi
FkGrCxhQRzC+e7ekwRomaRMTef8shXqQJuSNhuHThgV6caIAfDHnX0k/jOB1rNL7
e7ZNbW8V0b0HmDv6XY10Es/XfAXt5zlLaaLA+QL2RmtDGCRujZmcccEoL/P/7AYX
BIPmd8rAQ1I2lRZClFnw5P5y3cKE5ybstDW3KordEDVfY5fl5/7SiWKKHT9SZyaX
eHY0U6yRXmgAPyEFDs0CEauQQSLWEiuB0qexoFa3i+OeHwAIjvdyTWIOk7EbZK0C
KtT8rzAlXWbrx/ZFlgm/ElRlqhu8/o5Gi3KWikUf77q+0yAPQhfqajcn7JGXmSed
f/fP+hT+YL+dxk4BQ4M8OxCSqFQy+O7FKWOPFGtjyW3wUlO6RFUEDPFMnMPNoRa8
PukRdgk1TYyfB5QJyj0pbGr6eSttYe1QANVf6svfSjDxWNYjTkAZEOEFPJxsw1Fz
hC7VMA5Owp1Gn9ND0eI3Pz2W5HV9yTQgcTkRAj4A3+UA/Et6WoNJ0PRznrRMjlG1
rshCZPz6A47vAGklkbjZ1YjEhvTc8sJVCfF2rFRHcZqgTIDqS0bu0N7xOWUkV1B1
wkpOH2X8pXBPpDmH7Q4evMt3xer8Iw9x9k0XqR0QgVLZfZ/xz5qzxX/3/e4dHPzy
VFliucGrR0Yv3BnlsZ0Uiqr8Un3tgE5u6ToazeG85FXJ0dBRoHmtDnfFvLAMjkgj
dX7+8SqNklnqus7W9vIq12fn38lVUPrq30doXdtT31znoO4aZ/Eo4a/uUeRuVOn5
D2iPNFhvqTM+pGcw693bfwZ2mHuZHD3YD9kWndBgp+mq5To65jdY6wWxsHQDl0jf
GTRTUfybqchoF8BIZ9elqMURaH83gjHd+5OB5rYLS+/SsE5DxR4MpQRGQt4vzl+e
0hoEmk3T7+cHwRMwwDkjMWM6s4rxev7AE5Qyygl1BhNMW26saXFnm78s+76HI8br
7IK1FElffHztHtHqqw8P8a0RM4BMbd3b4QHTibeoAwE/+Qyb+rpbT7NBXkJS+wQ9
51099bwC1oeeLYeJj/Ucanob+H0ceSYsDK2iZIga50la+Lg4d6zMwRsvjXXAeoC8
UaCBef/tz1vURem5scZr0/FPhcDaiFs9NTsWo3zGQa7rBlcHfpXLT22FzGMv0uEm
hOTRQapQTHuGy18nEjiIbDDaOJS1GLjYAXB/KK6/zt680MbL+o7snFdgcgbUr1g9
aSMnGNItz9a3cVopjDHwHG3B3CP4c3+zSyG5X1MeYBip7rlmupkUTwz5gJ1ut0+v
c4nytBBpmLvoBPki2RYAPqDe0GQgcHozKcheZ/wlmapYZbkWiKpENuZaiNWSyxuw
SIqkGvppK/kJb6ebLIcilyREAiVTpAff0cdj1o1g3Z/UB6FH509xCN0WD3WNpiI6
UtiZ6HifSseCvW7QWlRTK8odHOI1293dN0fch1XCN6DZyKCCU1mftBgY+g6IKclq
yX4rLNNarlnMeXnXvSlT0tntfxUoT7L/GPnjDJkJcbAtG+Lybg1TcH+UecCGWBuh
QTVrUoNsz58QJNxpsPrfcFStv7AOJFIOuhFOSsw/6GzFjxlibbX1oFPLABpQRHo8
hOrZ0306St160nF9A4qIlh/qYzEjs/ROh4FTprOuYmx9eNBh40LJ7LEZdR0j7EzB
k+a4qedcxlpWjPluL5LC2GzF6EYJ7AoAPoM0owAJiE4MyZ8j65ZV/NiVv/Hr3XI4
8qCCmPbnKgv7Kn+5jZfxhRhjs1VP7rhzLl+kX4pKXPJtjpoZIo36XIyD7awlpv3m
iPJC66F4K7YfdMMrciguEu+dKG89VThOqeymOopadRQcIVKB63x7+DFFYQZ9LsLX
zFt+Dh6sgrFAidAoNI01N5mPVReuH3sF/YCDpdHSMUWRwQIt4Q8uFsJtY4nQXK/k
1Fm7EX/ZUmrKC4ZHFZ2kGqW/SvB+kubBiEd9bGDNPGLxsEUgYbt1ZdUFSogwIHPe
Htu85IWIbM1uGN7eMimrh40IeK4IKDWS4gINHfcOZbvu+b6MWz6CVGBMwFKFc3if
9dX38gT3RB6gJRf9P9t1IFqQhsuo9K7Cj5c/qZHfH6r3UwmH7iKtnKx3vSaQGYd/
PqhR9mR/Vd7uRVEFSK3v8ScoMrMbd/+34Rd9KHXz4bCxXUxAcRBE6m9Y8KRWuOof
0ajqw8iD6NskSFggLVw/V2z9YcxNuswpQDxFjdCDSvlAycXsAspIiB0KFZsFBsnc
7IG6jphkzD5Zsz0u22sD16PxEt66UDL2DAmDE96z5aWNL3o2SbMzWLmYf/8J//Uc
mPGtMOqKWisdskrIkJxdrgi9tjqtjhPUKPKckG6H+ZNONl7XGo/Hs3/Btt65LDF4
6N1osfvP0zFMb28DpEAQ9g5FPxD4YHdN88kRVkAVqcHvoTkbTQGkIw7VrGRKSwEZ
J3OgyN2aPWaB1nzanSLfzP+0tWLsjiKDGh7bFOHNehN3E9g18+WW9F7UcI5CHZhM
Kn2hU1gX9860EZ9DZjXM9350fr+3V+t9yDFypjy7JkEhhBMGbiJFE9TW1+/oUsjs
Xlqra0OIDYld0spMZpslEy5GX3mg/WVv3ykBZ0Uk3KEOQInxSIysYSFGRhdrM+rB
sbi2nkYlXS3OG95zzQFockpOm9G50jfU1ctFo+HfQ7f6I9fPT+YUctxeMOrQKFzg
XHDZtzIAu4EvWQHU+jTXcnkyjLaJAl6YqvduK+dFDCt2lfW/afgqsDQMhSMNjPhY
RN3HJ2esHTvq4j8EyT7/sVmaPQLutDNPN9q/BvGCa0K1XVXJApZQ45WhtuZRz+aN
e6RzUKXXB/aoKzh0KK2Eu6pakfzFTEPGhIteVFJiCUkna6KCwalTjxYOS2fh5vad
8WNpGCcbvgaN9R/z/XjzQPWuV1rpJiUlUITp3NuGv9K6ByynLayFr8InD91nC0QB
TugNWH5iR40f9SBMacT/XlB39BWkB/vTZABdsUCvmhLEr1+KqJnUJ640haNdL/aZ
6Hgz8mw9HvU6+saYM7cPF4vRb8l3PtzcOBz8SPudUyrsUwxUQX4RYyttKLkeBBEP
O90wxZPU+vMTy2aGHLdRJVd/QpCwQisSWH8uhPo0wU7L8pOu9hrCc46sobpSkidM
4FdfLacjnpIkLBHcpJ3rR+hdk3bEeY8QfOXhn90Wmm1rqiHUgYJnJJTLfy4FrZWJ
8zaqcGHHolJ+pBY28TurUY+ibJcZiTOXkXkr2ViOqtMVYlWL95PNR0aX3IgSiynz
G2UHt/sgUKu+Lgd1rhZ/jeSik/qhNFUQfoVDh5Ei42YDym87hwlf8AtTkFjlNDHN
RHADzUFLU5/97KaXoctd/Qpgzvkq2QigxSEjBvaeDlAWSOOpUH9r0xUDhDwB7mzk
+usILStkqG0AWfYMF8djwi8aY4FrnjSMMDEurslMxJfpgwcyoTnEy1ZU1wi++/5R
1D4v4GleHdVWQ+rwgy8GoU+Pby/NzujUQq0To5YVrNZS0R2MC9dRIWksV8chWO94
ytmjUVqSXC+b/KMU6hHuudRSZzTQtPZ2pJQJJqZAX5Y9ahvk96Q9dxF+O41vy0OX
ADvySN2T/3pdtbZBeDBX5Ybyy5c3tssuNTlWR2krvYfSlJA2Zz6XpXsbedXViwE8
ys5R0cSoNkL6AJYduBKzkpmBS9mVlJE7k7dOXzWDaG1yGtNozO33yfOXqwPTF0CG
1nuve4OElrBkwXMqA+Wxi+KwScVqA34hY7cZ6HwBdO6b2uLQlAOqn9wwNEAGXeJD
ijHnyEUkMMhzJ2QdmCXLob7cXrWKQcSYliNYOC2BnZgf2W1MsNDv6iAtXjhckRb1
rZkVtDOhpUlovhK8UvyOxJ/KSxeZ7i0csutl483/1dpe1SGi4uO7svVD+pEY6tiQ
PcM1EQTQ5QJXiqikG7hgyGb1rFQMuukAf6NW6AtoZDv9xqG5ei/zVqtGCoaRGfWp
VB85sx5PPNNIkxuJu+dE8nZ3OYE6wetiXKG9oS4SWTVFqjqhHH+L3N8JzHgeM2eB
JR1Ko47e5Vd9A+MbuoXr3aprlW6HJga4tFAWN2cnvRGNgoECrqufG6s/jEHGOdQg
V4Njcdo7de5FLY6+8xhbAisGlEi6U7LFDTfIsISmuWRwCg0aIUp3sT18KmZXL4VS
DsP8MIrs1YjYhznlDnGTzyke1ZYUKuWeuzy/i5VOUMm6SiM53iKqvpgjI1EliEtv
OVv+uvC2qH6MYoGYNjdcXiWxggob/+AKxWt6ffsJU8U0MU2XlE50PS97ctDJDC8s
7o72o0RF+EtaKVdLA54mNFM39mxIpHS0LFG/0UEeq9l32HRGqLTcGcs38/rD9QWl
WVPpm7VTWM1fiaia65ADtrvbNzdkEOinjLqIXXz2NrsKUFqTh6l1uv9KBJMvrh6A
Oh3V+sd8lfQbTTmpyE3GA6NUXpY2kHWgC3LU0h2oU/ULpSJIallLK8vWOKgjlzBU
/qzG/Z/R9iyuTw29LD0EtO4n8Ya/Qk3QOxiRnTXQnZ5n6yn0Px0M1/LUcZuZoUtZ
9T2jyOkC/BjCCBDxCV1uNRXnpArPKuumpL/NSgv2DMKsRpVCst5RxGJVvLx7dbrC
T8QA8wDKHYxPUF109xdRkKTRnMNNDdIk+j/Q/hZz0NGG/uyLnPlcG/fKZYpUwnFM
V5kS0IPNAeNBS4QR2UTK/w58G7pUYwydTtMmn88yPNCt8XqMm55Q5rdivGxNFeQr
KCUMw3qBEgnzqiWQ6D6gMZnZ7OBs0NzRFs6pIiIKVmmtz4MmenRMKZUVO1vuXzq+
CF5ZYX6msmAR7ZPMO7KwFNKTNnU2yUDLtzk6aeH8BeHbNeMIfyppT5447Bui21J3
KgOC+XNrPvGKcX4ejQGFAdUoFYVYocrUGLDj6KZiOkrBRYNl75/AMs84u/XEw0/d
iANrkErpufadKBUA6OnEpJBRJVSMsCzDbqYriu8FQa0rIPi0D0WcZhf3eSvRnvV8
XS+q/Veb7/7OFO4j0NeN+RY1Ep5fy1HxAo2gyOlpH1qVlaRbEQoqYVK90srXb5DF
o3FIL20u0QBbufzvZ1nblqJQMENCmCSR6Un0ie3me2uxodJfM4OV3kVVzDl4BADI
lfEa/azd+E53WfWQWJgCfG5/ifYz35btTd6eQcWmGhua9rr5O8L9EHLMvuZUFwdy
6/rTtB7Qk5AiSvEr9w2xuDyCGV80B8OA2Qw++l/TPn/yJwJz8PIWiC1I1bgY51DH
8+QgoIFoPCktOspCLrj7aK5jprKsi2rPBTpydpGolavFcy8lVP3cweuvlfEceX7s
BvJbe4pTZ77FSdSfxPpyrGUZIGZZCz5+KdQSsQ9bdzkEjCq3qtt52BVZERVmUddF
n3Re3UIvHTCc/dKe7YoWvoxh6OwnkH4S++xQUTptBi3NUnjVMZ7vA1Vc+gNjeTpF
ZQJlZ/aXqLQF7gFeD7O6YEaliMQD3aj4MvgDJHVtN1FGfPhqOEhpRuS3g9fwKCW/
yiXc65UxOcR0ukvzdou1BRBa7DXR7EjF0IA0vRH5mCzeQ5FqRpl3LGpInhHftiY/
VY/5ErKhI9ggY5XSAslPA0tU0kd8WrACWJJfWAffMN/Tz6eC6KkDy/doR45fH5pN
WVjCbKuyRPyUX3fnjMWUbqpQmb2dctCVnbcf7VlMVPQA6XqFjdO14GtNpYyMnkCv
zGmYShAFA8El0Uu/ejMpArdQiuVP79nz9MUCwAAFEO3qojotzPYBtoZA1/1KDN6s
+3opsqeBZ70LuBlvB/fj5y4eTVbQm5QQrnHHWCoMCNeXDFdu2idupM7IkTzoXLtO
+Vhc6ZAiTTl6LqoY21BGmvpSvxdMf0ejRYG9BCElVHfLLF4JYdu8hudUjiB+0VTI
6834OwX3lEOEiMzCNYt4UvH0hOqw24Wu/WOz+z4vxDLSOmxhdf+sNrafkl1ibxGN
oHwX4YMUcyaQi9girm7NZQ9a4N643Q6JGD8Uugw2X+DQVT7R8zy/3aQOQAGrT4X7
GcP6LnFwgc+qbvQoHXxLVqblrUB4gs80fz/MUw+626wBiWV2dJ8IuDj3HJUDnqxl
XRuttGnrImYvZU8hajxB1s1h8OntJwwXbE7uFJE4VEW2x6M3mY3IPPohjIWG2N+1
JvsOXXwp7g/raIshAbJjKzDa9wPotVx78qMz+B1TgRg4Ycw87FDyRFyIunienF33
wnCUW7bwqrZvXOviiU26gyXQKW4A8AP8GQo5ioTaApSv+7i2PUjj7Azhlv5xMBuV
fayijI2VyjMkGiE9Yui/XMIWY/WnYI6HwyMIscYduvuLeUnpzD9n9zp+Jmi+Txjg
HYNP2Cpbt32vBgukc/tueGnacAPVplHqEY9XpJ1PSh4eWKZlLZ612LDNTHZ8vSmR
I1H+hu12/35e8YFLkbkHvp9swlK8OWrphrG1tBTvJY5eCwxFki99fvHoPap9zVYt
ThuBdeZ2/Fq01wsXgIXCe3X9bwaBrJuj/EcT7k396szpocf3SKCtWy9I1vh3h9qb
8MnUYzDV4IUkCWTty+zghsCZ2yDEba/EP6MsevM/t0eEigqDDdHmxxWzpcOUBHys
gHYflbhA7q9Vm0b3P2nsJznOykQdvFTZsm+bIkLYJfNhtv3tTTftgDk4vS43yDRx
9AkB8BbOY3L12cr4k2zO/Z4hbTEd0ow3ajez5T65QzBK2K3WyfoKlQIjjtIkvBlO
Kzavh9xo/hLqmiUVoT51qslV6Z4K7l3PzG0wHNZ7g8aEZyEl4W2K2ExiiHJAWvnH
RU6e5i4KWuSOuGgvmyXj0zeBFoaWCmjBO2xPcp+zifOXI6B5t5Mnx++z8lajCFjp
YL/lcbBItBP2+bv6lD6HTvBujRtxguV+kqM68AqAQJBkKFmUnR1E3lyFp1Ph2k3g
xlCHUC9e3D8OT4OpCkHwnZskivGNCLOY2ZE4B1dloCza3+Xu77yZo0BTos4LglxD
Q+mjIlfNUAIX0YUdsAAeiO0b07wPwCWlNsTDBtApvKHioL13Y1L6Kg6FwdZMjuce
aJD5CHhqfUCrgjmfMOAqkOuZEFvi6vTu1M91fmd96gYzJChqYUwu7SOO/AhFZkWe
H6a1HFu4G/RTc3NHsYziPdgtzdgqyi59qZHLqYPYi99mEhuD5fupSWkVirKdadnH
uqJRqbdtxwHD8M43yZb0XDug9gQW+XAHjNIYPlRtihmhNtQUznEsOCEs0tIWOAfq
FaLBj7kM5YGNWiFGqghAPZIhyr8ahmMezYOdbXsMqmc3y4ehUh11AkpVGIQ0jOeK
ikoJBWCYw096GPZIvxsPILcgiJQHZDTsyVfaU9d9+ffKr5p6a0IuqX9hwqRWzZR1
3aXtU+TkmkS/9cLFsecAeA9dBkEO58gpmvS77WrMLufkt9t/V/7Nfa0cCyPGZiSJ
9oxej25VHc8iqSU/ig2dMTMRZxos/ytT2i5xy5tiw0pRRerguWo09rdeRshrj03n
1QwJPoF9PNHBi7lb+qRJAqcGBgqyVQQe8rMNI93nGsvMSxaaQcohs4non3RQDxn2
ShHRYgruzeWDlJ0Oj8fh6vnnUGyR0uzhNHaC4kDRGNLygBt0NRWEz2BAExx5iPFv
SnhiZ8avGfv7B3lUsFKAmh0OCpj8Nm5IqiG6kPxaXCl0YgAUwIHTn85RtHGE/2L3
Pn8Qn9ACJRP/HMQcrmbG71BrL+QNURDQUPceRdeB6ZHw/QpwKCDuBP3fXhVtQPke
waOOOab8O3Qpua2bfAVvVvzheAt5jeBvgVIItawBBKuHQjW12xp6yyatAjFTBaXP
EAWqP7zOXCRVQ2FiT4B+FxIyGQyYavZvVpaMkJBW2soAxTiju8VUdqvP3zd0ouVp
5NQhy4e4a6AIrd3eAV646Z4vcEDUy9LCL901lV1ane9bCvR07quewi1geKg9IuaV
jFDuFUGtxv7PaZV7AquWF/ZD5gWnY/XjJisBQFaOzXz0q5gUFGAFZYFUWTu6WKdQ
Ayv3TptMVw+25r66IXclLAIwgB7nXNB0nPHKAEMefSYBZnwwaApEu+U5utn5DUr9
oqIFyq2CoYvvB3JNeUpcKE7TaUatPMuN3Pz9tm4eb5kOseexQoF/zhScFFfNIDge
aQprKsI5pu/ysW9hJ2HNJgb3Gddtoc0ae0EW8AHThAshYgibKOPncG2OmU3rIr4S
VIJffZdGXgCRDTREwTbD9TfkNFQw17/2OI5lnukRB5YjvGPEq/D9cfQhLsBDMSE4
Uub9HakCremHQHolkG6wkuK2QEvhUs51KF5BwHgq+H2Suce0c6tsNwEaMk7BpRzm
zQZ0QRIPM7fUiy6cuIDNkEw5pKO0FGYNg220Rg4PZZO1FBF/22Lc+d5L01dPYdO6
x1NTUnI7qSUs2XFBi5Jtnn010gMi7KiRXRRD11JryVTihgDQPI0JS+ei0tLQzPdn
36d1aQD880xqtscPt69T63UfVnTvuMjnyU8ohNNcatT0u5lIYchBBgyEzLe5M5eG
TAsAp6utxnyaF+sCPQUYCiEAmL/U7iq4hmqdZQQjQdA+H5v/NJkxis+eYlgDYrpU
2Bf3XMNPvy19BySuqYUsT9hm1ODYHDnhlm2eX3u3j7//7gETzMtxKLWwm9/vmMH3
JHRFFk0QxNmqmbjkYWj/3MzU0oob7w35uNU8cxH5UelYBcouA+moMbWOfgGP65TC
XvY0R8+Ai7guOtlMEYcKwMxJfKNFhmIkSreNT1LYZUaRj28xWrbJzCu93lCMGWqS
6v5ePyK8gMmZCKoJNS2bpXlDeoyuThiEr3EMyb0yh7Zrxb/cNYBaW9Obv6i5H3S9
hdi+tu1dii/X16N9ffL3peT0fEWBfvE18VDAXET5VqB/+vBAzXGQt6P+rboK7skt
rveZZhzZFHjxZIpbbSc4qMGn+6PRSr+UhTF2WDdck1U=
`protect END_PROTECTED
