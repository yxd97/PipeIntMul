`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9Tnhwo5u28JWNKDCDMZo9SgtBmEwpC0MjDK2ehlAhIxR9DLW0rPCIc55Q2O6r3TV
du1OaMYzf00mZolovcgAo2KlocRvoXzLVDCs6FcO+r2NAd9997dd+ZtrFHAMIa30
TjzEQzJLeePrT7WuMukYjibSLys6sIXzK8M/PEv/ytwWJDoaKL79qcYQFKQepnx7
Fr3I7tDeq4F2RQOD/dc2qFuJq4zZ70HCJ3OO+/pTSE/7gvxws6Np5j+PpqI4DuCC
s1puZj4no9gFmqMywKClawI7/bA/J8lCA4+WJast5LSFYTJkVMpGKdED6DFsm28z
SrL9mbeIJzMkYBsC7sxZwRG3572e38ELb3puMs/+1RbKZ/jG6kK47OtTCTBSqN92
g+MJqidr3BIMFr4CcDXrpjGHsSMo9JsMfkydTzAsklmY2zhu+Yh463oj1CjdlfX+
iJYjZbbrOOo6Eft77D+NL0NKo9oxQaVlwEqtzxfbY2FH7Zfz4R4EPGSmdQUA7XKr
Vi6NSvJZknQ5Yu0OMcxDmDUoZqeRjPkhXlv1nKU/6IIHAZ/8GA9KHsv0lH7b3Ugd
26dApFWNPTHbuGtX3kf27cc4+UzRPkbmxkn2HL2Jpuc=
`protect END_PROTECTED
