`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3tBo5ZVIU/dgNDJC0pObkNF6e821W4StEAFpAUBJy8XqdGFUQLsUysQs20KXF6v2
qz/r1qouGjLO04kmKVlcvgPoNrl7HQ/Cd3B/w7hIxNeI9zS+hWRTVqBi1TyPooVz
QakM4pay2Rfp6HD95sSGa+B7hLpzX8ye/lObCNLLh6fGkvXZJyWCh4z5mZ41A5pC
yNykB3SzaaEnBTxX9I6ml+ywNwlQ3JdImbJnM1W3yysnoPjNLNv4fSOXAa8ahQUI
Lm7Ya54C6kpz/181d+51+erMshxNLIu2EIWJ8GzwupY9gBFzrSgzV6ZAm7pPku3c
btQF8NyOaqvjDKJ55Mgw7DyGfFYUwbbaQJlE8SAUR+Ty2HgMeE8NmPJb5Mvup2js
VUVUFKMFJaizs8TQFLOl0gKh0b4HPzZ7f0ZezR6XB9He4WXE/jD+duQJM67QMPK/
vTMxy35maEyCXZ1zFESBUO6gNrShuPyHDLfmOse+EVQeWsXIKBkddz6Sqa9midGb
FwNOJw3CsIpXX13GRI7wnODckslzULWCCHtSko9hZDzaV545Cj9OllfRpucdOD/Z
6TSSRkYt2QaXFbk2T0Oep1byM3NangKJec7nfh2ke1wdDl4/W1zexmI6N/xLFCNQ
YgKpQDGgRLmmYfCSTmfiSLxW/MAv6APBzqRe/FuXI3uiwho7/ng+ScloJrlmDgS1
cnNdEWtmCyxuYrfE78pT4rwe8MUawTkwW2KGjkfaMhoJkybKabPSUgzFrbY2Pnh7
UaloiHtZ5E8k4VWL17jlo6MWByP4hQVq4N0Y29Bo9ESxm6sjfg4SJ/dMMltPZj9H
DFbhHasqKx638Tw8bkjadn/wU3N4Eb0Z9ehk5W3lEQCoGNRKx7EgQCfJvddRzzYH
BotZDRDz9BUkPOfEwjppg0TCf5EgcMls7mHldIjF5U5XmHY0Hb2zQ5ct+AkFb6Ui
S2WH3Kjq3SsDWqHTWYR47iVnVN59H631rUQhoAGQFCLEPd5RsDG2POwSdeFCSZ+x
2rweiQlGBdgV9z41TU2N+DYGjTY/Hh8VryRy2yPyA8krbhI+IFRmAtZr/dv0DWXR
piRwQ0yZtxWqWHXoXR5YI2X9Fu/kuVilGNajLI+WrRzL5ZqJUWAdT6ITCYWInJ08
Qu8ktK+de36MSVUnE5TxQrx90U1WRLKAf+R67vLDtOzTmHiFrTWJL4f4bukIUQk2
lhrfBeCcF4Lto4UdPnrvMWuI3M5a7pmXmOHmwB3yGQwYPG3WtMFAWrDYRc6QzMH0
lpA259lWM1eW8XtAZyikDi+LlkFRFTsmxEWoY8TIOSXUlJmp2rok84Dc8ESi7DhZ
bh6XZ3B6LaWjYVE+20sD8Anp62xe4xBbuOP4yht9taA=
`protect END_PROTECTED
