`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mvPrm6bPD3eYqtdzuuhP02Tb47Jq6LQb1DyB95EP2xOG9JbDCyHFPpa8ZpcnkW+t
hAz9J/hb/Fu/fZqqTpkTVq0fHKiXCEy5CgA++c4brUiJbfM1WczUrRAzG3UpF/nR
czMVoX1J8bgaSYNcsb9Z9m5vzwvYAdNNG/q1a7MHyZnRVNWU4BxDKEy1NUYe8krQ
Gg0Ycq/xIw5aMMsriK8ZhxrU2SPIrXOB/HxfGJ/5XkvOqFKuSkPz0Vcn68EIZOql
8Q7PjTRCewuyH+YcI3JupY0tYim4yl9fExfyu6tUGyQaVc+/vyuMk+fsIzvGoJQo
9HgZQv3yCxuNmCWvv3sD4Jtr6JFcnc99oKB+4tCzkz0S60oV11E94jqaS8gYQ/+B
g/tWg+u0HOFp5kG7iTDiWU2dubbYlAMbcbPyzG3N0inS5c4UIaK7RC1PqqFiboup
xWo7CO3EBx8pYfDy9BmYvxyqNO24H3X6ATdBh1bqAUJzaMFarasOIwl2g7qnt5qR
uLubsaVFn1aycdK/IKvaxy+iur01xCdbCLxH0qblqB3C4Z6O5+CkA+dNElRlw83V
3zZQHeiF0lu3qJOoWJ57+G9sp44TcC75RKChQ2MaRzskasarFvF6XOF2RWsWAoJ7
`protect END_PROTECTED
