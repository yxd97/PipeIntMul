`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t1SgQ1iFKCFb/Z0p/nU5LctoV6X6eYk9XD9OzUno+XuvL4OlaLjI9TiNJD6FJSmi
UgQCRuwX1AoVyjpD8jnHV9ktJvgFkzdFAUVg0UtnGoiZEF3exB0t42FYW0y0GXNx
wghhXFqj1DH8D1EjjZd4MeEBnbk5hbOU4zJtWAF7izGV/+rYBVycPqbA+i3Bj/FI
oC/xXqCzlmX8Ytqd/Ok8VT9oUphSHybfwU2QFBKVc6/hTLJH3TJ1YbRisnvB+7l6
A20n0qh+mfaJfzIMyYEVMQDeD6zELL7JftqS/Ru0GrdxA1vOeAS0ZFRtsk6h5Epe
33g3SxMGlufEiJhmWGOLNKlY+N6PCbl9HPLwdzoPmrSKObJCxSPiP02Ux0cC9S6O
7iHST9zHkL/T9ZbRPEjSyqV3SBtrYZZEqmolyrZSc4Q=
`protect END_PROTECTED
