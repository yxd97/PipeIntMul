`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ZZgdocQAY+Q7qPvA+y7lI2WlJ/vl2VB1ZfMx06e8ZktV0tC/OqGBIkJVJaUv+BY
A3+CVIdVA8iTHUnTAlixHBYJYqLufJI3SpilFn0E8mz22FTsP3sBv0QZB8PuEkUg
K2chwbzNvdlmgGaD374I8gHBCxIj8kPRnP7hv5ZuUFC1Pk4AsNA+YThVY+SLPAhy
uwkEzWu3jnqbmeNpyl8M9VOImsZ+3iLsSDyKpdjr3nqNKagI0Ecnm+ccyl3Ig/HM
ImnhUK5hBI1a/0ZdFfIMV6mPRQLsDYg9OEc/HUE0Ds6/mXO6TtZEldAi6fT6pgy2
fKAOBEQXtOabl0kbfyR7Nw==
`protect END_PROTECTED
