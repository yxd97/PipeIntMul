`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4gkESkGWzJaLo15Hqak84VxpIjYTzuH3avJ5Hb8R8NPovU76sFU43oQG5lHOTDfS
cKSHOpTvYbkLARD+m8gnd3M+k9/J8pWAyUT/MzMChGwgjh+OVegkrIr3S1QE/04f
Tqx6zoiGBKmQ99Ktj1XeIuwAqDG5bLyL0L2kFz/vBNkmWBfH7sorQ2lW1wy5iBYP
/VPLA4Us+La9KVl6qYnr8XWE0RY6g6XXs6lXWlC9GuLwddqaJ7kMbr+4OozUy6Vq
mx48u1xxyDqzm38v5VhFqwQcB3AtdvFItQ2u2EofutmtLZjgneUY/jHZA7fuSyBl
vDaeLMsYFklQeD981oyouQLiSMmWhoRmYvejTWZHARY+GKkoWAAgmxfplf+g86in
69CH9e1knDtII4w68+8bJXtaxc2BLgMY4VI+/mmjxuMo1LLIN0sIWGpQfrRo6OnK
4YHX+k4Ba2NXPAwjfqYZlNTx5iVdLf9lchBh1Ha5AWB0lGmB27+8zCbukoC2K9As
pLG0Fe+eZQlPfcf1f6h3mjcUvGAGcxME3T25SuhCSCKZzDXOGRIPhUyw6hKKamWP
bQ/Rtvba3egaGlFsrDV4+1sEei1HyNM1RGutv9Q12Kz12h4M3j0HbBrTjKAuuUwG
`protect END_PROTECTED
