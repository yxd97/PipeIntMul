`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EU4KyEAJubCpC5hlcmm7nRZ86iPonMXK9m7Q7OsNL0yEF2dEfkeybqct6JPij/FV
S+CLcH7w81/xBBHd0kY9FUEnbR9PaPL2dJUSlaeVnXQulj3JWKlx1XSWBiGFgR9X
lX9TSHZSjv1Gn04TgIzGf/fKORnKyg+aaVBsO+MCKKi8PKPJwCDRnZj5nJcs/JWJ
gdUaw9pN4B1p6SQnZ0KBmcPUPE3IrtHNORsoSXhOzfTfM05qYbnbFDmHUC1UGJL2
lE3t5h9wVfQyp3ZhFIvWOe3fH2Cy0phHQje72aSHo9f6GLC2UF+yxkyS4KwxtqVf
emVCYsr0BrwtHOGAzRoBstbfHPUxoQDZ5PRYrmKC1zQSWNz9CuK0Gxh7/jrUD53V
QNXVZrtVOn/+d4BLYFoEd5XjeQkebVU6HCuJBRHzh0p1NzZ4JuojtxMzoaeBucS9
H6B3RxHAzFSyO3TIhy5eSSAFfzvj6K3szfqB+ISzwu56iShoT6qnilduOOK6q/+W
/SN7QPuu/ZIJ/qA7ATANKg==
`protect END_PROTECTED
