`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6LjRTvAK7KwjC1cZ+0z3HvcF0rtQc6GkT+4BjaIZjzInWIohtJY5/Sv+wokjQGVw
29gZA2PBy/SS8yQtT84YN1/OdOuSVwskNnghuXBEUnyFCh8EDWFyPlbyJAok3qaq
Ak6FR5282PQK+kaM/sjg5hyVMGB3e1eoOexR1UXd+3YjrvnZTFsL+9ez0UF4E32J
CH/cOuWImkGsx+07bbWIo6rMzMIZbNyKyJMFco5GekyCtSyyw/iS1p8b1D0dhA/N
/Xd4XcSg9CqaUPYattl/fv1BpnLthTtTGL7dKx4GlXj5prmVL4v0Y16HnL0yi90T
dwxpgYiKCwtXAzHLpeoMZzKWeWuu6ralKqOfLvVUDyLGojhIH3f90N0q9Zgmk66h
E7P7ekOc7n4avtmhMcV/o1hdtH9TT6bEqR3YOS8vMVT57liO7J8BfURT+mXjsNI5
QMQFtZamfYRzslpDvGdZfCoCydgNtiS1xKEibEMaG3BH5/62yh5PC9tPmFY+8P/D
lYRVgpRwsflY5fVskFDI98pcaJCGvpDpiaOOUCAV99noNq0/3vf90o7o7I1d6cZR
eKO4bpR6JhrGmli4lXANiyxGf1ORce51hQvC8I1PoRn5dUxiY1OSdZYf8Gk3yC+f
KpY7sJCSHLaYu4CwMZKKoSUg3lcNSv2kQFOWINb34wzsgbAa88yoCWl8eEfucrcl
ce5NDH8flhAT3lAiQ3ysKYaPHLBADOX1qrpInIkUSF1rOwRM47EYQf8P7a/OmHZa
9HdTtgQo3P+5KLHggiaNTWFaoLDPrgvleMvq1yNpXnViGmmP2QNAr82iQ5GDKjuS
/eQAOtmxGy7MogxMwOWk7DCcoB3w5H6F/hFASZaK9wvOwNIu/VuuYQ32iACHDMUW
cLffcqUpcohIMdQ9uWV09g7j8QOAk2uafKSjt/64rFqi0ov4iJLiVUNA9LxEtSC9
kIUYqdO8IQAIR1tecFlOFqPhdsey0kCyvN939JH2o03vUrldBiaion86x+jSLUZG
x5bnd97OLqtGq9aarIdCrK3L0zU3jh1QnbvzS50dXGvszTiXKKyeCcMCU9NAyJsv
W9IXZOjaaeoHxpFWqjJ2vVoyw3/wpyHZHXF1slgyPEQ9nKUrH3sAUB3mKMJgkw2k
eVnbUJ214nQA37oiwYOMpEAJyytkoADUCq//zDqza258Hjk1Qf99MSKURGZrSArA
y/lNz4W+OIVRlBGDuO2EqXsm4+Pv7hxL03AegMoKbiEMuqlckjggvtLlvAhe+Jc4
XV+huD2bxmqU1rPrByZIcuYaEBQFppHsqAgn6UrszlyrO1AXQ1CwH0ybzfOdfJdP
/tqiv7ZxVGHxsjMjwADcbSdaETajSwgAri8/2aSvcz5Sz1YWxnjkFNLo7IlZRiw4
TwiefwT3TJ3y3mm36BxNQRShgnljYMTlOWv8s/QfAOM=
`protect END_PROTECTED
