`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Dw9h28yktF6SWasz0tMTiNXA9urFzU70IaN28Oj0qVVdqknrnkyeWj4roRYEXFX
0qNQD1yCBBnooqPUCfcA+Er/6OWfM46Kdhc+rRFgfO4IPsvFcNKYBfBkyyj5aB8X
UYDkJ1qnDwcylZmAtOfVePB8v+ht5fqC3XrNmgxtXF5DtuK7cCburpTnNwBcBZkO
X09c1DAzzhjctbJrufR0vOaltMtKKk2UwNF5Qb4z0L0iIvNrIhBvAFWr26NsY0RM
dJVwqnzZorlNC1h4YRTiG7+xLsslTJ2YGxlImkVSuRybFX0mzGC+NQUM7cZx+tai
zTk/8dqJ0SXA5/JjdR4l7g==
`protect END_PROTECTED
