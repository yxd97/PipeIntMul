`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
POeHO28ypDC0w8uZnxx0he1MlRNtsZoVApsDYqmSd5sZTrpZC64uhTF6/NPwYSDk
ggzMihTViibx/TYa5aezfhkQAdPTS2LXlJGCqEBD60Qkd/zdVUEx+2S0dSVmnKkN
ClzRV/pZrKFslaRfRvHrYov98C7StaHBD4G263V6PO8haOv/UsFtSn1mQfjdcazO
SHSrmFLNhZMhDvUEmHiaqVmg80jH0vhOphbZlkYdIJRtDsUhcBTo0Bh2MLPTDBvY
muZz545mT4K2wGebr5NngJw9tQMLY2QRAtVQhL2LilcGqmyJIdMIvcDWSnkA3PN4
URI4cRZA5duTJ1ncgspAevgSjqTscoChE/XXlP6MfDbL2wDRZtxvWzO9lif01CYr
lnt6dNAc4SDFRD5ZsgXv8w==
`protect END_PROTECTED
