`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t3UPh30GPHnBIUw0NvDXMOzPV4gcWYCm7V9QZm0YT57u7HcVfz93J6/VH62tT7B9
SnQzqN2JZ4BVByJzxohykfYjd/RjYS0rsftZX4PNRD4izz+mA7oLTU6DNFWkBwSX
i3CaPSNX4UcZot2ftZQuAresTMLrfxFZP2bsZnvHCoBtZ+coH55jB41Wmb7GZ1an
djvinzSyhjIlppVY6wlXBQNGmB54hz9TOgpQCJF0fNeVGNOkSZkpWjA7sAIUTp/L
wiJxBzYrsrIrYQJe3gr42PC3HOl4pFXZ4I5O/fikonJmYV0IwTf3npPiIYwRxJiO
DZRI3SUbV+QrFKpdhSGw6qYwBO4tPTmEMlbV8WogC9KetQKyIGe7fTre9L8hT+Km
GQPVF5H4A3hZHBqG9dJvdln6vOmacG0CPH8c9bsJatIX8odbR2SfL5NQQr+ujvwH
gE5ptHESIzhzW1ETaD6UbYQQQwevogCUff0H3FtOEN2/Rw/LyBTMYlEOdJ5knVVf
AOvulWkcrtSRFNvJuith13o24jxeIFcCfb37bXYtkEHitguiI0uer9Oe4N2UgWxH
BdDtgkBccCqv9cvZb1BQ0t37RxgXscoZ9buoKPVEyeY3yHdF69yzTGVOZjT3uKJm
nMm4KC2aUnSRjDBoiVlhlJG4/Q8vAowUUkklJOEuaCUsnybiTdt4ALmd1bbCDQ5V
pappT7HfHCud9R4VbDSDIu4aDGVmwotMH63CFRKOhDTzWQLwVwNHVlaj/XbJ3ZPt
jksxVsNwYgtPlUrKy4ieAJjTJ1yCrfjJEBbcQtYePyFqtJ1b/XSrBc6NFOrDQurH
sTIKBpl/enPUGLFjYpTAuJiLuYf6KhMUU9lDQmuM4ObRSxUpUAwvVhJTmCS9mY6Q
5QaMTcB9UqPM+qL5/see/E3G4f3dQNyXORcmcp3PnZmGRA8gZ+1b0ioWAjp0rwUZ
aASbuDP12z4oJ4FeZ1rh8OihkoHi1OFRhHiliSvjA7Sk3WO3CpS86o2smWmrBz/2
`protect END_PROTECTED
