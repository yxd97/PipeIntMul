`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WlFdhdh5p5h6ZLmG9laqJYqiXUfqMkr6SRXiiHuFPLCv9w7l0qF2iuHlR625Wunb
z94adxRpWKS9xrP6rCeFkXA7AoVVMmP1+XfzZ0DMxreomq4hM7MMEYiJ+IuLbDQ1
jMR/cpcWjwqmycw8jmVeNhD9Fv1zH6IL+kaT0rJSLlGuXH5v5yR8lSFKISSTP2Bv
43gyKatg7kEuTtIQQLs5EYLmCtTO5Y0qPTqSRpYhnYCADR9DfbdK67wbDcG8uoJU
5N/eCRsKF5VD6XjdGbSZoCe3OP+HMmxLJoHfSLdLOTSgLGDkbW7poE9R7wY3+8aG
1dDoQO2Say7rJTZ7tPeaoPTF7d9Lis1eDwmJ5Fm0ADhLmRLq2w/rPCLOtS1qZaCB
Ht4cSRSGPoe092kj2jmijGxqWGsveovzDU1iigCOGYGtnCnznDt1O0t/YxOvhKb4
KmiErnZSkfeW+gwy0O1k8ZuQWshK1kvkQn5lwE//x9U2qXtGHxrc3Urqi93LO/Fy
NfGY+4C+cWezKaGzow5zFf3PddLhVuXrFA++V0NwVMudBGtp8FKMRx3g+b4GzJ4z
eIlnHwFams5T9f8zROw9JBJFEBG93GCy03m7O2aUvHQepv2Hc8w/Bi74BV2c2T3j
vW+amMCzdt5Xm3IJk32XieeMo59D7e6FRZM6LdhqfgIqLErP6hIJdNVjyxAYMWof
xhBiFpnovVQnKwj5xdYsU1szY08P0KvgX+8MLIT0nIbbjdxd+6KDebQ3mrTxqn+J
VrSwuFg2Bb0Aw91XsdnrEIoCKa2e0hf8uUFv2LWeymrxzltaUetD59o8OMW2+dZ6
uNhYzRVyEsj0wVNzA0RGLwQ4W+Y1T30aBcI3cTB/5+01FP4UgCmjXQZrkb9ARNmD
2owYtH3SCxnnCry1tQoRly4wP9xSpmGXFTB0xZFp5WL+AuQ6hWoQOOnrY/Q+QNkj
13snDEwumq57wyYYeqISxXRhrmcuwLA7satUvUoV4J5d4omuwXmbunxXY9EInwnV
e5Z1WF54VorH7fdUaMJ5DXRliaeRV/OkPa9wt32YYNaYt+TADC3Zcd+9POA3tDxb
TxiG6kGII7xNJKii5RviP6PDcp0bDWuo0XRQBYPWlc9p6qg2eqAwjU++80PmkSnL
OEjvBlWbJswOHNB2i8SGPEbNPD9M/8DDh/iH7/CQZ/u8iuFNb6d7oIErUn8AlrJd
k3Yq1wmRqX3+KTfKjN5OHeQFMC5rHPG3bhXRAI42zUV/iLfh7Q/Q02D8LFz50e2T
hA//esLIfKk84DKHbEAidf0V36TWylGsUscOaP5ZwVBevMHgDPEu0PQK76leGNK7
bXlCOJNmBu+g6avypn0O6IZHalxUqvcBcoKWxJOZ4GRQE2wfliSyaiwMVTGTlGBS
94VCFGRp/bn+JRlVsXJ60A45w/WzGI2760SXUKnR28xWsMlcx1fswK5ftI40oEwx
F7tpRxG7uY+MMFvWQxwlJ1B3s0xem9tzKjWgt7l9SpThzyIfto8/G7pdtpEh+5Ve
zqYMeoFwR76TyQDWaqj+rfB57yT7ArSDYmQYv8tJWsheR0XfauQfptRyDrWF2s9f
UkRSMzcJeiV22LN4D53Bcw/cJMEJqdoewzh+xf9s3qrB+iQ59GwBteiQAeObpOUd
zYVHPyVQmxOXhVUgLbyPChEJfTLiW12d/VSYqqyBr4uWTr2nDjmTCMjvOvPUDaXC
Y7ZrUuisjhVI8Z1rI3TlKPkHHSelNB0gYfM9xKPxoTGQsG6rPXCACN8imyUh/en3
9zcRDN9ULR5MFAdeXbaKKXHO/0eX6/S5443Alh9oH+bFMPtCiRiciXkmY70smREb
S3wfNKXpXPYL3uwFU9nkBVVkHZsEVvt3dHqSce/sYOdD2RsxV+M6QuqfMkdq9azV
NuXWDMPcxSWoGzUGyJe9QAQ4y8G4VYNHwmumKExJJdDeUzioes+L5jYLf74Hz+Bs
OhjDKdrUd1KZz/q5WMzCzEi711YGANABUNANtrFhiE3nyNAyy94gyftijBeSGGnF
5utw0fhn2+TruXz7lVLYmgx0MNJ4qeqio9ca4vPK+qwxRRrs3Xg/C8nJ+4L+bUtw
xZz+1yZVMvKBsHyhxXLyug6W60Obnu+/QG4s0JAuKAg+Sat668Xfx8hoHCqo55ts
aAWvnfZIJFoup7E9Wvo9J8hzH+gfUKa4UxgQd5nDHUhLKjz9OFe+G86YkzHbtVaX
CvksqURw12ydsHVNTuGQLrZFPjVXdS9YlA4g2cvTs2C2nWHCXhr1hh6GAB4yYJvf
yiAaL2C9YSQUCBI+0LxSi4wcRFy01Tc6YdARhl+nvDj49sPUW3jkVBLUaGOq/ExR
Bh0jdZmArhcnIf5ots8RvdK/iD+eIPofkTeGXDAW8pxDqj4J1+tzbByqVsM4PcWO
sHbeSmLGVPTZpGyyBOuTWcwzCT1ccKrhkd+aZG4Py8CmukjXu2lI6vZSrzOuY494
k8bh5n8NUrn8zIN7QjsKbBpOgEOuE9r9PHli4b16djD/PHxFa6ywW8KVINdTqQFL
1hbXZjrz0tVKSw8b8AeR8MvfIyiCcd2Y+Qza71NCprK4UMzX4ALW2tBJpwdiCgam
RJqBSizZtWWUP9QrHis3QhhfxfrfYJKryqFk356gCfRMT9jWlXISdFHMTamnkngP
KnwWo4DCdK1RM1B0rMN5apbzBmnbHHcrsVxpoGBz5D3VJglRTD7bJl9XWGLWSQH/
FUpGPDecXoQBPJAlQTuxn7n1ANmBE8OzYSBu1xb/S8i53P5+PiuIcO1SQpcmoerK
fVxeC+yA2cMdm3jE1tzfmZrA8zjGjc12LNk/MEHdZ+aetQVXBCyNs7I6tjR0hPvL
DuE3QTgRmk0p2uIOsg2SrygmmFpcM8L/1Xb5xolnME0nNRdpBWF92G0YeB0l4Ran
5YiFm6UdpZ7fhgrDOURmHd5djPWHPB+72BggMzfYkGAzgcQ8w+nKqIEWKozvhn0r
9zaCrnzmAeEq6zWtkG6LcMIBrlFY99ditC82C57HBbQ7VxHPgHm/5gWOIkgv2r5r
NU5O9e6EvsVL2EUZRkJ8W2fWt8XzPcLEClRIf+zgiXG+ZfefEv/UycK9yXvLUGYw
udh7bNN6iuMMPE076bp4MUzF5/hRMx61g9S0klrutCeOWZHct+oCKXJRh3Xe+8VE
Y0g0vInwI4CozHH9TxVP1AThRuagLO6lrVR0lfgtOkui8p0wzYcPTd2o/V8TeqE9
ArHiU3S6ksUZt6CWdkQLObsQ+LA3CG/qax6CLTv+LxnaJGB+WiFEJsUCtehBrgdR
aoc5i26CtAHonKqKP1UcIWSAlOQJKXJMDeO+sr61fW4IiyBf/akLC458Lh1vparj
3HOX6aG4uEEquJXAMVWEm099E6g7JBmd4dRH34yQ2/4J6sRKlu2yxFpNg834n2CH
8HiJ1TQdhY46si8W3kZVMQ4y3C9Y9Lbq4aKJtlzt86l9oaPqoiQKpXpM8n+gx5gQ
lGZlPDuKdgon++vz/wNIhsL4cUxMbB6ehcO/ohljbklMllafno3pjyorNMf0G2lp
qT+fT2JKtmTbQTEACrcM02sFTCPg2vkKxRKdqJWmsAVBGL8CwtAIPor+3h715/DM
5nMxBOv5HS138WPTSJ6uD4rhAaHsg/4PsPlslDaHUTZQ4fAgf6SLgumya6Zx7LS6
u6YpOaoeVSgonrqd7ncWJP8reUC3TQvbuFF88xjmmgfJO0e33ej45fWbaSM6ttE9
71wQmjPauEQ2qIBPr9QDwRCGYX/F3KzkXdGz5utqQYGbo1O/vjcmNbPw/7yf5OPK
qodpAxJJ0eP8fHh4/HzBDq0tkRxh1lXxO1H/djti87avls2QYOqXmBc7dBN3KlPB
79WYWnaPD18FsB3VgOV/p0HiSUkRFF0nsrkU9BJ8PALLGklLaEWIcD1tgxk123iO
s7hOh8ONcsf75Ej6Ioke6mXAACdvAa+ayNJ9TIPWaKh3lkrSzCJS2mc4HkUlWR0T
SLm9ZCZBwAvcJmu6sqOGtx1Qr2BoI2imrGKLYg5fCAbNHQ8qQ7xyyJLP80+nVKMc
mVmZ9iQ5sVfFeHRFe0Uvn30H7cZWU3GG87L2QFOx+tG37gTS7Thxf58nOLMNys0J
Gd5RxZp9RumjtvJG64iDWMsVj/w4vSFd5yAQdLoEMQOC0TXgpS/GKyKiM2ZhSXEa
AwAhwy26ohB0iDPbatmPWBw4RJ8OLhhATRwRWT6eEnzNKc2t0/wE1rreh24xSwK6
k+pbwEM9KxqhUIcly3b8HyTeOrE2L0BP++o5jxU8k+gs3EETykwvQdF43n3jBLNL
D0sJ6Fqi0sp1LuQNhZkrAgASq0GHAflKmw+o/JJ12oGsimq3XdN7mhRdchRlmLOX
BQwv+dkKYDLCopQs/RTBxsANAkit02GG43HosZb0uXhTMfFHg8QGrRiDkFTUfQkQ
zSKPa4CovzzMbrg9ZzGMee8/emiysjw1shcAhGc3YlZiYmNeRoRbmnURmVC4rJFW
tjjlGJP3zd6xzvf94RjQB9ul2fT7hytXFYjbPK1KwtJk7862alUJ1R2pRxX/4J2K
7Zea7+JSFdCkK5dkDvKLyc0FYga8xU7DDI/3KjCEIfPW9/MT/rk9KysQGJzxRmRy
8UESmHWqK0D9m6z/U5BFaeED7RI2CcIkFbOX7kuUXVMDa593Wo7WvmI10fbuKw5m
24uJ4A9wW32ftXG/zdjHupth+mKHI9h6PSKf8Kawffy0fGIDauQvOUI6VeD5g3ob
taK8AJ80N0fl8xaMyY9fJV9v4l0w0MtHoH7sT6pZ75fMqKA79Z+uRSmiG/IX8d1P
C81mHi2zqb2RktxT1ldWZQYxChof4LbN/aHrZugfn1deBXuuryHx8Xc7hgRmsuA7
BwaDM9o/JnOsoytdDB4urUCfjyDmpgR7ryQy1iDW1iH8VJO3u93xJUdlujktf14Z
HMOk9amiLk/HnPAkr2zYENSQ8gz190QaUxRuU6dSL5nDcjusR9fob4ooKb/r81Eo
9f0u4Ve7WHRkcIad88YBdZCvF8tDezNYqSsIVRDaBp4up6UjDFyduRmNrDdUTQGQ
aSzFC6HrraqxA+L0qjOQr1ZTIhCj2IhmFJkeNJEiadMPmKv96W8EvD15eIiGsrNR
RlFVDAA68PmnJiLat1/UCBE0ta7/XhOk5hNbZRs8z3h0c+nmhRJtya6N3Jleg4xt
d/1zlKOcuFeVC0uG2oZwkNhvqXNUbK5kOb2NbH7nfVMWymetWcQMshuT8jrrbxf5
jDSUKF6ngi9IsVLR7E+1yAhmJ7tsvX+XE8CzqcxBlFr80Q1hb7KdZ/8aW6hRCJNp
HifDa9cDTLTFHWmcSUzANrPd3bqVk4ULmH6JdjQv227QCayUkZFdcTswOaGveS1T
WnPw90hra76uzgMT/cm5a405eFOGQGgnONUvJ0/eqYZu08Staq/ts3dtXO/3RR3g
LLqLtGIL4xhdFEc0zfTqelJe6tp9Gx6yPt3+A5v8QW0uFWUiPurucD4ZdsZVxuHh
VE0WcLD7TecXpXLFFZ/qmsx9gdcs3/Cf/NYUfoxt0EnDXio3efGukZOkpT+GZ/xK
UsIIwAFeNvLthTJX8vBy5LuQD4hnYp6wDjYT7MLGE90pDr0FwgpkwZbbDa99yRnP
lrxJGCoX3abbcnoXXyL1x1mGZj75XuxTKITTdkaeOo0fTcqwzyZPwm7kOQzcMpUD
7UYVTvqKra7hdGwhNK9VXllqm9kAPNq7b8oKGwcXKF4AG8e5B8y70Qnr7v1Bh/Gu
R5LoZXkOW28ms+aB29phvHBM8JY1srkhTk8w9uFVYTFJMjb6rUaKcYr4YriI7EWc
WAQTpqYDNZsLp8FaNc9KwfNI1W16zi6t0W+RKYhoX5GU378ijafbt1DKCbyT5w3A
Mdm6uenTw0E/h8Yf4ejteIQUEi+ZhChs0wuSOTBFqHRhJu2hc3qavBwDKXWAIPB6
lo76sTAByyXgceXAkLi5pqYJsPDy1TWO2fNy3MgHeZdhEMvVcz1GsUhQjp3RB7L4
/1Y11BsBXGjiWwY7ibIEhzIwZpHH+cs609K2elAVL8el9iqW3KtRL3FNt1VnU+cG
qseJ/PyErRTgkeBW2TeC8tqQN6qjwm/t6533AwGYXNvUT4g9XrOTz1F+Hr3iADqn
Zhfaj4TG+Io/aszCwSJcGmzfFhX1x1eISRGWSMxygnPtXMX5P57bc6tlLzKPey3X
IecauofxAXfToAEdJAK3niPzqrJ/vyM6ZwP6fw3lkwieliAP7i4mFA11SQETYzC+
6Gp1q0Gyn8RspuLgeu+TPdtRjgXxmt8LGwcgjOcdmZQnFxNp0G8akl8xfMbrVqwB
WV3NmOmwhjo+z7rJoLkVS+IEzQZzALfAjKPjIafAl85VLYXk6aBqNMILbb0YcrW8
FaM/H/1IZVT+pKOyrQBOyz7zOBxE6sJ0oiqOAwsqaXhGHplLJEKbuRVG8H1Ma9oq
7uNRFGIP3eYmqcQf09H1+yioLQ85OiQSoVK6LSt5D8//x/CGHRfbfR6XNqP5cXOM
auaOGU9iGltZkJ4GJgW0usnXuWk2TRFBkLcMgtxwJWHsAOBvM47KAwX/hQaZW1qA
WX8CISMUo4EobG8mzqIyKKFRFg94eBwIFADqmlK578jUtRVYiEjdHhSHel0ZOQ9W
s3iIJqPMe0fV7rApRLxZ06UFGikVqR0HU3jMo0xjzeHPyhy5glEgEKx/trP6MZ1H
PTymzBwrJJa3WbBD/nKERPIT0ucGwhtbV750lCH3cag=
`protect END_PROTECTED
