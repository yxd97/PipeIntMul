`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mef/l96cpKKCTrA2ipWaNu5hSDb9MrZsiAt8nCEB684RDGZrzQYwtiz4+VSWRhpq
0XN9Lma0oFfMNKex+EMbkGvFBEQqcb8LPZ+FwY0zLtXyg1sF1/EZ1KlJzTdGg27h
WHTOPMQ9A/kNeonAd4vwmWWmwIvVnYnD1tAEUBNNoolmgW7vgm2tn5WKh3A5SGc9
zLd/oWHhG36L/cQwqf8IJnSheXz1P3jYSvRvTeVeC8+CjRQm5G3zAHW37k/4YQtT
IkK7SZCpqu1ZVpAfoubBLFhqxk1cWsR/2D9p+EAcR8FQfNpxFFE6Q7KPgUgLddVB
jclt3PVH62w00NF6wo0u8Lx1T4JK4mbaPmCmLvvf7FPaX7RdulZPC18/m+l9krk7
HiU4pkSzbQ+DB+fchtbwpxzK15HyTNJEdSrJEhlJwhEewexcXNWv2sFtz2elRAW0
`protect END_PROTECTED
