`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wQK4Dy2MUugMDDA0+z9i+q/JI1h1blC5z3yrPRxfEjteUI5Sr8CQxNHZ+2/h8Xkc
NZ0GSSpTDKYy3zV5senJ83l7Zafw8vNl2GT+YlYbixR7xx/9kbgsoircKgUnEL0Q
5LLE7M86GzTw24wg226IAuvMvFcaj4Otwy6GSTdGIbjFffjrRAOsQ+vXYJ3LcZPX
egL7QOUIi7707I1vW7tOeq3SlG3zpR34DWKrHuwwTiLXSaPHbY1hNtreXzuZ/pKp
`protect END_PROTECTED
