`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s6zy221/8MoDY5aKlj4qmh/AR39ZNpqbO40VHGkx97jNUaSnRMfuTANPypKWExz/
uv8Nc86ujQZkj9z1BEyhjCJcKkDGxu97Zro5Bw+N4ZMUSWZQEB2VGdL3e3b7cdlp
qQQqM5AUFzTOvgHmBZqzfnKNQbCIiUMDa+NLPimk9TJE9MwlPyQ7MTbKvsi0YXBL
Oetclj4YFu+aoYUqpNriUg0UJxVbue7vuFoDB+8SMaUW+d3v0iXLK+rMqjR+1CXl
ga1XiYWU3+2aCwSKJOPOvjqsYs9k5/Tv+Vb/jYb5X+SsAAktK4P826JrUdqoy2wO
VMueKNcdFs0Bu8s20mzP0sMT+rrFXhmJ9IXIV1FxOgB/CPGCXsCBU6rzAD2wTaJl
2VgtgwPP0bWfcuh64I4E3noUIxLzpAA0BtYZ+MRyjoud2xVASXD6iiVZNeUk8QSC
N17V3M4+S66MWo6vQ7heEndVUOjpl0RoQz7hxmg5xI97w4LG6cvXrvGdt1aps/Nr
s00hO+K2YY0Q8RK9hiNzFqfSokP8aidFFOtMxfaGdynKItBnEOIoTonJleGMXqlG
r9f3hPoSqzPkMZQFXS45N97vb8RMXpoQCwMc2nwg/xK5AZnXDWYtJ0gro9vHBATb
hhb8ycnPWrUA1EcVzHXh64EBfcdiVEkNeIrgosPggJLF3Rlu+Fy8QTF6ZTO6ny1v
hj5JVH01Kvvs5iYKtdony5mdcuhwKp3qkfxcU3XekvTdOOV2Com41bdyV2a78cac
wxZwWiZg3u5Rz3vVNhbyXQsM9tYi8IMcJEj48Ug4Mqgzt7rVHOWtjxcQUFzDEx6o
+fcyHaajrwRd7SILUYtix3Pubng8y9nNJqFIOX7mPKs=
`protect END_PROTECTED
