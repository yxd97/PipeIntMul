`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E5dMmL8h2KzwZFeAZ/mCZezRTHbjER7M6CTQmaqo7t8Ef5Z6rusKNatncamkY4HL
f5Xdwnk5gx8zEpbPwOQPTM4xttkNmxf29mJS9tzjcOilpCJFcx/mACgwTtvMF7Me
itL2adwI7khps1YZBTWlewvmyVQEZ0PWW9/lZYZvgbt9D+STHamhDwq14Ew/E1dJ
G8NaybL4dg5uR7NywWOT65ma+ewWfoh+g5LlyyP4dRCcA0Q55+y/ow6jJyHVeSrR
YVRSpOmC8yg6UGovX22O+DalJsKswot2W6Cvz5sJxPZ7KAza3cWRmL80YvZEFZB9
TJ2WPgtcNigNJjGkHZqtfKWMfuIBHee9yqrZUsNkmC6UcgSY4wFBvp7olGKRfEn/
VkhevBPRzU5pZebMKoME23YVy5PjFqMy4dkMx7Kus2obi+q/JeTj8vBaY7NAede8
XnPinl25cs9CIJc0tVTvNZj3eluI3Yz9IWkgsu+6VHLBCzGT/Pno4k+eP5ElJdaS
zudzKb0Y7U8S4GIcjpndMH7VUUgUppgcW3ym9puIJ9q5FURKzq6yi7qrGTxc/hpW
/CPlZG30WZWj9SY5ngpv/CLgguhrzAlQ/CG3XBQjI/xI85+qs6fOYXSmxexiI5Ea
LOXTZOi0Vk+lQ7Cz4/VbawjKrJ75cG2tGxbZTy0gGkBifZpa6FUJBTHi2px4DLTI
KK+5/vGImi3SGPs3jdhuig==
`protect END_PROTECTED
