`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4rgepqSdDR9/kGR4jHMKMI+KqPtgZn+mWH5NZqacuXGnh+RmDXVejvBPUF6nVbkx
sN3UpPq2fWaJESE2F7gXd/iCbfm8M0vC+MC/a+mzbsDFrBfV599l2wjjdLaYfOfn
N8vaK7159PNzDyvjDHxx9C/lPZ7BJ//WgYU75mSc46JTu477MFUQCQzHqC0FZMsF
fluZbbD7MH00IGheOqhnODzUlsldIzcsZTxmxDRHLWBHwAxAbgPPSb/Z0Y3DmpId
X9m8bU9sYJJrhLnZAKA2ls/Xzq6nchtNkhxii7M1/wPj496BeFyoJ+2guszarARj
/9dnR1rkKwL7TBCN/FNUvxlMb9CBfK6Z+mepjsGQQn+i8mkrTwG65S1k1Aq67Tdn
M7AGA8JBmy04LlWVqyiVkoKVWkGz5639CUkH9/0HKWY=
`protect END_PROTECTED
