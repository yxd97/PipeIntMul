`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F6dUTItTAy8E3TqPngyUwt7OUkzDgGuAqnMQ5V0OBk7gmTjXRgm9c/+O99anxXTk
0ENVAvhQG99J/i5Aa7lGBlocGuehcMKcrWf6uB7PrapgQOurCwfI7mFbss1OpNr6
xavXWRDeAZelqGXHYDxsAsS7pbJnXpDddZ0Ano33gOhBdWJxJW0GgZKAPtmBYxq3
aaypFFNGz3jJk0thhzUM4HrgH/xtctwSlBddEHRh9pYhQXh+V4lEalTVL30TJVVS
yRypnnK3ePx/eDSFbfsdvJloIagUylZGKt8AXiEDPXY0vzYXJM/Rb1iMXqpjWEYQ
klPFu005O7c4XxQeF3DruWdh1N38RKppjvRNOza8R9y0UYA5AXWZCEJcrEwKF9oR
sbgJksito/3lsrVRJic9JbVPocoOdCXf10bSw4yqCFJrGic5v1tRik394y9KlVq7
tLWdGM8fPf9raGDWIyxzLIclXI8ZvCzDNmTH+eYd00PqZkdnrl/oG7k2AhoXukUg
qHVCg5kaj4Ba6aB+hivOuXgjRHJ6eHuur02eeIdSZyceeT6jH3FW6CROdGwAf5Fe
Wjgtm9HGuOjMuOcc43WV10ILC7bs4n9XgJI2uZNSBPi9QxZOzy8p2/TF1Py/wmj+
BuE+tZZbOfwtTkb8Yp/Ubunpg/qBEiMXb/qesd2Qy4kVbEisNQsuTVAf14FIYrUy
z5maSultx8mvStuUd+twDy0zK1KDl1eMIbn9j6WIsD8sKnE0FKkaH6oULWAd5K+B
d6gU1teR64o3DMgVaVZJN5lHRqme/UmIIZV0oiwmFvEkBC8IZgLl3eFzvldYjuoe
dyk/JHxNadMpbPh6v3tAE27tI0+ACIcl+LRFk+UJxvPf5fDkdSRF4QEj5WwcLZjF
tHAkXGfv95fVQkmY/IWEOxp7g6bZTeUiW2uHBzpblPn0beKPHp9fLK+b6zmKOq9S
jFn+/lBfEaZT8Cgzx1cZxAiH62FaztYfkNrDJbOK1E8y64ajYV+B8wC4GjJFdxs9
1LpUvPtOltEgg7D0ZNUL5cifpG49BzkYtByv+zXJ9upBlrS/yzhJwACf1ysLak4q
lP+9LxmFhpcPjDDxcvN4FGnp4qOnmkXcpMsSS8nVYaqa8QH7nF6tFLWW5iEGdET7
`protect END_PROTECTED
