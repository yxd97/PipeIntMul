`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
riK7195lboJQdWGskA4ZB/a7V3dHnzrwKs3/2ry6pbXdP9cAl07dMBdR4T9FKC3e
fXgtVIRFHGfuTDTprch2gL/DqKCSi/gC8gzSKmBeQ8ccEJLyq3eEf51LnsmEQpzb
Q8ur8GP1lnT4DBi5FPaeIK+ZWOtIPr+vNVz6tt/7R86xuwAoY7vO/q8S+/ESG+4J
0OKZvTd7KPSF0mJCGZ0AWLe1gH2oqIXzTYv2Ax3j62AmxAHM2CCJNSEJSgoatYuC
Pw3YNnMfINLvovXrL70NMWigyWnn8QPeaEfHignwSLyTCHPTKkrEp6xOCqDOKJk9
PKapQlB5b/v4an99PIeljxLgadWHPXKkeruTkT1KK4nDFuTVMmtyfznd7QzCrZ9M
dl5KvlZz2qG4MS3C6ZIX9UsQxQsLkB/1r0T9IUaUweg=
`protect END_PROTECTED
