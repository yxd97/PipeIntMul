`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+y+7pRKk+Sm1qokMUwkVk2XHUOvlHI0cqmj8eeJxJipAxU4SgBZbtfIFEZs191hc
spdKuN4ER/bXaSZwRqIudweOFkMGggUoFJ4WLIlOHyjLoazCfZDJQJwJTT/89ZT+
N0dg6FQiIfSsANM1Xr7ARegAsyObd6TrUETYmYlUZdIk8Hxrt35ldp4j9EB4Y7AD
eFp031WneOiTbWouf3yAcZ0ZAz5oGL8bBcF+6Xd3Fslkujx5gGpT6PiOni0tYamJ
Yq9GPVYZixVWng6se/Lne1oW6ahuuTB7YmvQFBFJDljP2DHQMuxftNX6jcl3POw7
F3OPtp4nJs6b8MLqBWssQ+uqm1emDV4Pycrs5hUDUPxE6itJGhEh3vW67qR5bNlB
C6nlMUbidd9uxysJx8k6UQE0h9nipr73Wl13ZMAnpuarKu/5Ipy/S6qbhEYgozfP
9EREZRfA07+FPpf8KnU6sxoncq2nvAxyCxGoHAMvCv2+nkDUfnjn2wsogkRndSnE
kVQpdpJtpU/9A5BFLYuSraiLI0ET/9pxwHxN1tOqwH7JpqYp/n0T4e3ZjjCqOOEZ
nao1SL4ipRJnruJ8W80Hz7z4NdKiHyIZ2uzQ0e2Ok6Rjop5fvkmmPTuWYT+kXCm5
R/O9jf79qYFGws4T5uBJSw==
`protect END_PROTECTED
