`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rdgJMMrV0ns5ZNdzMBlHovSntaYnSTZ1FjxIhu8a/VQVsoQczpHLTJvS0CDK7Ukr
8qapQmTFlls1jVR7QYb1JxeZiO8RCeHAzRTohQ/gfwgWLiC+nGV8ls1929Ii2kwy
H5sST1gmM3Mpvcs1YQHamp3E+8EC/2+mmXOVPTuZbSJcmWmGO9H0dFc9+QhCB2Ts
XOFDoDoQqt4X+A0ncU/uRjuN/1efuVENyC0BMO5hIx5wxB/TFr6jV+d6jyRBnLZr
CwzzS1TjoLufrDBNg61lEfLCE8EZtiFjZIJ6ewnRXZqmz3SzTIelQ3JWul3Z2Ixq
433ZGhxSPH9ibLMwokktDSxgJUdkCSUSIO65WUhmPBmusVgko+mDxCSSYGWNBHLj
LYcnmPM5V2DVZDh627F/yShF+aXM9oyi/seA17+t6SXCWZcMqE6W8FDEiAG66NrM
zzvHQgIAxr0IMbrcAb5EJqwlU/xHq1hL3oPxWHmFQmT8n0Q1+Rf1rC+Cyjs0sPg6
J0iLa7b3RQSCzz1CFN6zJJ0DM7PfJ+A3L+R/dQ6UgNCVUf4NxZbpuaShUYdgNLsZ
`protect END_PROTECTED
