`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fwwYSUBGezZANuZcHwS8u+iCmIBHht1OnjQTz/AXxbC2waZALbNtQR/imANxgX8I
c+C/6VaMzY1vg7Cb10+hcrcTfeMhfszBYlmQInAUTqT9qNsfyOnJgawMG2cCklau
+Zhh2n30fcU7qcKnaFPael97GqPunbf+2+IvBDfMKK8BjSMkyiDKRH35tQe7/JQE
N88aqkxLUfKlw0Tmf6OwOen6mkeGOvpqHSGNHMvjqHRzXrWhO8ej+Uy5uNPRhwIw
XPVOnM3b6udP6TqiB5a2arW6d20Or/lYRr3kBRhXjIo=
`protect END_PROTECTED
