`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Ik8hdOu6J7DfgrNokOD936iwGiBvE2LckdLH/rpwsmoPyrbT0UZZbATp+sVpppV
E60lGGWly09Dt5FgcjqndjzI5cRlujMAOLp86tU+0tdN5DyJUjFE+80mGOu5A3sw
8yPfATft9Xf8cCugZR4cwU4Z3T+IQjzgCQ/BAYC6THe4HSJar+qHoM1YKB0B2U5q
mONKRdibCYhczNfkT6zj7RnvUrtg6Zd2D8qGC6DK3Re+SfPex6P3ErQ5Kk2Pupdg
005Z3o5JWnOL3CPv6BdjEqCTmO1tXJDdR/5VfDJYXLGVR5hlQyPO3gl72R5vBCZz
t1PVyv0HwgI+RUeP6EM5H4xLGWV7mhiKj44vST0GSma/YenvRjK4J61dazai5xky
PJnf8szISwsW0ROTr2vbSeMt/umIFhRLYrndnuRQ3Jc5jT8xMlYtRazswU/yjTjS
`protect END_PROTECTED
