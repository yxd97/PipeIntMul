`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6oQwn/cMASbz2TEP1eoOJ+LY2nHwdIuH+szziDSzC2iME+OIodpifxxCzKlNG1As
3tEr9AkC+6gjcjVRe4EwBfdkFFVYMGmxd8P8ZdqH/W+qVhQpnzwFV78+I8JwvQ7R
7g1gOG30Q2mjXQGuF/A3f/VuXKxpOX4gPhvx4l3M6bozLhbUoDOB4ABDTUY0tliP
aYaj69P7Xeb31Z/4einmmcBF4i3z1ohysRj9uBw0tk+i4xf0AQB5nS1ow87kahgq
1uFAi4KIbJwqLJzI7e1Y3kOwTlHNdkVumQGXj36FWtnmiN35uSgrj2CVyNxDzLPn
8S14ufAWA0nqmUauUT9C/WDJXXW9za9tX6aZI4pPpRM+r18aEUAiU6IyXoa+l/i/
hefUAivm3ifJkk9CHm6D5BZYAUZPzOPCfc3plwK2pyM/9fhUwZzbT2rnaLp986If
sTDzxHXD+uh+tAeCkyrfmr8z5ajLI6cwogma2JDnqAiENYefdJo48uUR40ISEcni
sVe297Ue8Sv7+Ea8HvEK9GO9YQruh5iNwtmGUtc3aNooL3SBsgr7WV7lk7wldFR1
HlkAaxBvkGd1YAb3r57bYjPtcLNtgfsU6n6oJ14E7REDCzs6B4NXZZ7lte3oqNBn
yuNxFHN+wGqPsj8OZ8f11gYapeAg4pBQovjTn6eI3i7AumkdB/8a/JLB9I3rR0M4
P6jLSdjgV//r0QgfOaJ18rpN3XHmjbP7vTnPkIOvYQDI1KDPBLZX8jShI6uhwuFD
htMpC8KcPr13LZfQe0L58G9yo5fe/1htIApUL0ovfPuXnu10j4joz6dfLO9zUDsI
OryGxS8HQEbswzrEGHGUqX2fpFn8E3giPQSizHh+OgfYaeIydix5VMPI2h7O10Yn
4xl4D+X6LqkYpXP5fAKGOWhHYhUm/UTN5QsFjc4rr09mpZMH+gVdz1YTl1IYMY75
wftAYsQWmOps2Z8Bb7PKuFXiJlJXXkVSB/KRcw2gaJLWWbR8zSbR9F6q2h9YX+kN
gFCkXo7jA4oxqmyVYWhHR36tj5ZXSK+r57Ul8HFEhQ1/WsiGX2dIxMCYELkXTToZ
lDerROu+Q6zojMqA3171vvsR2RTaC1m15sWe349fIQCg167WXcud3BN7GIpnO/zS
UIWAHu6PtJS058F+tU2OT7luBew0rEt/XcWr5q1F2Zkf+g8xHxLSuJxDt1Q8W9+Z
dEmTEWaRTNBvuB273v8m4Pz7gYcs+mOQ/PQX2Klc4AaFqkHp0/54TQzUuyhlYpyx
n7OdesJjBKhVtlWEOCW0i0q8oS9dLqlbV9m1jxpoDT5so0uZBcT49XicyhNjYAAB
sxkx5hAOjE2NAZYvOnxD2r+/EkV4uL1Qak0trbCavX19hZCB8hm7ahlTgwlq60QF
SqBkTTjRNUlWONBihmwYjxVlQd6hqkukP1qluK8+ddrcM1v+OEjtLWdlYiA+T9bX
3BcUabX1R+54aOb8sIUuNNpXF8YqCAQaP9sCrqPhLAt420Ujv2+hv1mYrEExvgJi
ukh9tzzq1tionSaKpOytcIRXndBkEcaMJUGsKpW0hiFlplyfxVMl9s12BkSYxdyR
7jGUxZFwhpMpiskH9pfuXdAYpTN1rj40L5qf1vm+0Zs6z9ajX6JxrmQeXE+wQ1gI
uL6/ZXWOlm48U9RhUaVq1e024JwFT++uOJey/mT4vslUpCz1KaR4GKRCoQlxINx6
Rox9EhOTkXivL6sdyRQKUNiLFBQG6lNB5+DbHQpx2U7BHy61fq+HjMKVXWAEWtdo
L844+vvVjXaFsFhmknuiBQL1l0ApdNKeDMQ3lSnsfvV7LCRhIXlAIWoZpaEj6HLO
lGGp6AnAsLHNTDtrxf2QU0cDXWXjn3Ana1Fgg7foq9RHAHdOPWMVkH2P0kRUrrL/
AaNr0wqChZG8+Ih5m882t5gIV5kHxmrLs3Mp4BBISQNIKYthP5mvaoKWkW9qS2hs
JjCWlGBASsi77XfuBZxfl0qJxMXAHWgCKVLcGaAmu2DIlIcS5QNQ/XT+2+BoczX7
`protect END_PROTECTED
