`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fXw/4XZ9p0VJEJ270NwyV0kuyYVi7jp/loTip0a/G+CfVV4UVoUPA2086j4q5ZHQ
60sofxt5PskRMfD04ncglaKVkDLjyxwQqasxmOp4GTTqzIXOQVcKK1X8iQUFiXpY
mi8tAKQ4B8IPV2pVksXme0StQfSeIlafi5Y9CKugMLD5rEUN78vjZCSKd0RgW6N4
tZdWzqlFbtasuY+f5Y7Iqqetl3i4RlItnJ7wLY7bqCSzbqdP0pKaQrYyiAsOt+EG
lQuy4T7p3rWKUPK1KutYThzrKM85zIofWI8F+TpS/NLls24ndke0VWFsXZDQjHSu
A/NG0dAmSGz1Xs3mNTKhto+AqjgZpzrcn14l7TvSeq99au2YWWTKpJjzitd1akXe
Rwk9i4UecDK9aoJd6BbH/v0PWWo7d4v+4/oQa5G/tomSa2jUxgpx+ApgOsoeupat
fo/A55arzo4if2nzSbTjcLTZ1irqxEn8J/6gVxPl/mfVofVKbJGGJEBc3R+2cE1G
j/f0uWiGXLmo3Y7y2rRD1Fkevva1d6UbV+Rxua7qtb6gWExh7U6sUNVUw1ll/G+u
+CAw+vmv7JtJ/6JR/asL5++57u2O9+BYDISQyyplYSiNJOYxHtpfqYSc3rRlVPcd
XRYp0znSPYTdrRT2uVR4WeijQTMBG37vZ9NbXIQHNqrEu2zhoU7HnaGlWEPZDZUO
BhyURlfmA68uEy013EZUYNRN5J8xWdjIlQUDVlYnF8jmpXmfLPDYON8lnI/8lBwr
8r1L7q9h6nuUxlfhUZmFr2+G5LKEYdeE9c1H3DcrPylNOUtq9hlYvSaR8/tZrYLD
ZYyTiR982XH2qTwBch0dUi1VvI+B2UrpZJIFUEP0FzPH7vsu/7b+QHdnp1+9y76s
vroxetTVa7Ol7ftnOqE30bXgSKdFtk+vHd8XCtCqNjm5NE8U+yefC/MiKmhTXpq+
xwm5gT24IAiQ/NGJ39zR97Rf/cdUwmX1bNAreumTWdq9a0nKTlF6HvDGPyJ4ihB3
KVS43enOcJk06+/zZnflyogjaz4S2mk/Ev1dzhFdL1WggxTZ3YVIXMUTkGwnndgV
g2FsTiH+bkCcVDojhBzk1KHq34oMWow2vOtes7m/VlR37Fr63okrm/BGsunize9I
BrTYHKqY6sjF68dibbR+wGvF1isgcEBtX2NJxGuS3F7PGaHqgCkGKtrhO+h5ZlTm
nK3qBwZlIsbWbZ6YiFIrvM4PRSszNTyLWLPRpAGG5I5x0PaYIJBisAFE8Mz9MHOq
l6V6xF75fToK1QOG808WDQ==
`protect END_PROTECTED
