`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V5dNvmBCWgBivtrL2iF3FjvcuFdMqdcNCwX9CzvdveK3p1TthGk5/xslnsUkc5Ue
qGYuEuDMd4ZgnCNQeXmR0/W7I3pnlQ4ERWlgbQm0QEk6ZgZK8Yh7uYCkStp5rOnc
+vX54pBa9ljZfDtqNkTQJdRmDTzRG2R5W8EpqV/B4jlWL6n5v6ecw2FcmldSeKMW
OvlJQkPII4FkSZt1NGHf2AsSP4kGpHZoGazMBYZSOTzvsKCDcvyeGQ0WqO6RXHV9
FOc2UEi2tz31zH2LI+KDWA==
`protect END_PROTECTED
