`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RP/EOaeRJ0Il6UjckGauTfGqlUSbRpsfI0upuUUHloNT+Q9zqoQ5L12aO1qvyveQ
xNSIRjgVvFkDKCap2dWJ01fdxO5AsKUT91+4jaXShI4LM2FQWxN35PMQSPGOMK1I
yWnMiGR8ka0uu9GKyqkpJqED3hE2HbmS/l43GHeWyVNYQCKzZJUys6Nh7heBbasm
0dTffcRG2eASjafOBoGoKzUPDfRwcNiWnjsCWcxPParuFhsRVfQnIdEkttkRqh4x
UMfAv8Hwi+SYzBYhKNV9edpARx8s8ie6vpDvuzRWMpHFhJSeakdVEnfD6ztYKrWg
`protect END_PROTECTED
