`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CE4pAQkmcHCemU8rolWA1MxZX+1Q5nwWtFVulAh0tsxIufTrxZNv94JaTKmUq4+R
jVq7UyHV/ImGT3uuxcDbG7/cuS6f4+KVkCK5dHCFctW+Qtoy6QWDnVE4orqiGdmi
eMwGP6R8v+zKPdx9bQqS/jYwmvJnQyvNScsc+BUZmuduOZMgDxvhf9fahZxE6gnK
koM2fLj6/IwgmDvEfagoV6EPkKWDTVRFgaptudEfOqJ8MWDmBH3o5rBhTRZHFs+e
Jdw4g2D6wDJ6lsYkvJox996qQ0TvaDTQ6iHzG646AKKppympn3r3eeJQdVjSwfJT
6buO5oaUjDZrmvVnoIB+OT3aZeN8n7mb7E1kuqT1mClDwF2EZyaCN42xujkX6lyH
`protect END_PROTECTED
