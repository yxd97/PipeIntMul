`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9COR0MAVGVmDmbjrpTq2O+LlvNdaLpnOcfUWxWdmGPKgYdSe1fqgi42W9QXw46Qn
ZfEPwGt5SN8qm3ayrhNUBpObSGZSm/GTissV5Zs8Q+470z9v6l8AfJyy3MpxTZj6
EVUnjntUAq2aHNGpOgPhtBVrEpkZgqDdR0CIjL8aKA7pQOmtx04uGZKZgWv5KTyk
4eBPgFagNQU5tetfJ5OuanDo0aMJkl/xqfE7qO0S0qdI84zVxHWTn5Wu/cy6bj61
drsTEp2Av4oHDPj5tJzsApmmtgEmu8s9+E7GjIo8eQMIJsCPf1c6YiVqfKKfzbsk
GcVJd73BNY8XmqfOESO+UFLUCg6Sgff6sJ5WiS7SSt4EhiTh5f616t90co8etnx0
kv/7+mDFReW3lt7HiuBlMu+Q75xvJOmsuhEF1iXHkJHCXtG/OVQ+yMcfK99LdLc5
P8cmU4wSqbgzSU26zDsrx3EXXG6h57/bfP4ee3C+ZVNEpozQWYhPAnkqB9DRAws9
mYLrX/xt4iW0pN4nEFLNyugalxZ8eCH9XUtEmY249Nox7QNQrcuQUfxFEn/x5sPu
`protect END_PROTECTED
