`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k68qYIM3se+9hIi7qq41KDAPXJtpJMcEKs6k+nC7rBnLSrR8QK9R9GWqF+yNl00N
HGWKWFeYFQAgtoB7abjFH4sbP2LmbM21BpcXbTnI6abLmHEIvfU9SrWQq/P6L3XQ
erutg6Nl3/jiHB4uWlxskBE1JjbMk95vzVyy0oGSTKo7KbdM8J6kVD9gg9bPwvTr
2blarxXthVItRu2Y2afswuS4sBmM8FXdF/EzQRPUwSw+UjWRV/RimEn3kSAMmYOX
7ceQLr2zGTqpGFRTRhcc9LB2n7g0oTK/LcKcbeRPwV6EXNU7djlu+fXEzOYpsnbN
`protect END_PROTECTED
