`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vbfHiCGa1fv46+1z1rVhDxPhG/cLDEvKRfuRfSeCIPEaz5TS9aGNh5n5V+8UZJg8
Fh9hHoXYVNlnD1jEPqcdq26kD0Q8WVqXi387CmUKWC1afCFARfGjRs4cL09UzbF+
I3+k2ivxVU/VG6Djxg17MklXVwll1YYyFOY4lAYNaOE8B7M0QiVWwy4MGudcdRTE
xXIMXPF06lMRyHNZlQgBn3jHfVWxyMTlJ+YEdB7ncCQXfwOB2dQnHq67/TYxIcBj
yo+LD2viyEOB+DC+xnaAAQpZkKaPO5mBPqCYW0N5fLkPp615nrObU5MbBlMIfciK
MSCm8Llb6UL8TdJO3a3HpQ==
`protect END_PROTECTED
