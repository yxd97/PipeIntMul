`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LwoBLaumWLaxIa3EsIUJUcMGnmVxNLtXZxR/MAIPEnSoJgh0xHYnnKcylCJQwsEO
gfnN3TufYy+gEYCXdLzNckR6sfxTqR7XyVrfDwquPyURwGpvR0kf4xVcECiqRbeO
cbwsnBP9RX1LcJUIgvy1GdagieaMTVISdMsaULfzRHdMD76U40/X/bQp4Wd2agBb
hNT8/1r5BH84GziBhrhQtMUlE5LFm7AUElMvvtFqUPL2Pc7obM04fVeIjA5pNgqd
5Bbg86Pk+AQd4vqqmptSQax0T8Ou8LYIgjgd8tQxzWE=
`protect END_PROTECTED
