`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
szMaFG6QfzsVHKcyChY+mTZgDj0kkkQMTiSznq6plDhsBCePo7l9Blo3ieneDYeV
b2qniKzW2z8DSJeWj8P0PR1vSWFgM3ygZANIl+VShgxzGE+8kf25fePybYSEwCQE
C2Kzli1J19X39NcFd+uv8K2aRLwZAkvgwuVMw4UegaIKpsAhdfUr0yAwy4N5Zb9W
1/cl+rhhpwcK2gjmhLV7WgXtVZ/Hu1QSY29h1GXwdw8ry/+BOiOxKph39jBFsKxJ
UzHIy9DDvE6jXLunL/PmBNTwnEU1Anh0sX2jZcGJzmQxd22Z8HbKlgcwhcIfd/Nl
VqHvF9EPKfDbHpNXCAdcFoNXx9wEor71xj+s0ij9nboHNLXx7P0awdqolIJPHCRt
mZ09bgcr1r1b6V3LQGSyhc9CKQO8UJqWmI9WTCFAneA=
`protect END_PROTECTED
