`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MuTVRH9bBQHaRzulc56AS0Tbsf6f6T9xsUjuy6K2rHKW6KVUb574dCIOwsjtipaZ
lpKP+nrgkucc5RBUMp1fjl7St90G9hvw20ffXlrOwOKT+7XkkgEV7E9egBUOF+s+
2gIXN5MtaSoBmwe6nTtExjm9mbyyrHWrpjFNyfwXrp21wc6fH4IKM70oO8CdSxtV
L4O1KyIrfWYSU/fZ1wJP27r444wTe/jUC3p2jkce/tKmSGecnmNRNVIPpykhRv86
idN34ZtpYyKX6VOkAbhpfgJfR/0DFON1RKcODvHfs+SiB5JcUS7I3L4ccInnSJhE
XjLwJUj+dX3p66X4Bu2mdH6BbuDX/laY8Jg3M9uRCt2gwyrofde97FQbnW5FhCo5
tZlNWoEUn6vbJFOHxAHGdiRPG4erF/3slXNwwNilAM2qI+LXuuUnRXUzvtAPmdMx
a+szR2iMNvHQJnYjPbFcZIuF2yb2zmYdCzS4CcmwXj5f+4SK1VtFsHiCEPovS2tT
4CMpcdkGjeIJCnNQUgNipk74msxVMq9b8/UYQgUWePMu0hSSaZY5XdYIl8S2JY/O
Heu3Ccawr5k2YepldjL0dbY2SuuJdvP0J+CHNroFIoZuRoOZsC7R66JSSPa3Cxvg
WAwRx2DvOGnkJdnT1drRFkXRjVFBgmFPwgoO+vkZVG/YfjJnrRAAkbZBerH4EJit
wj91c3pTiu1XMjdkweGnakKWiVXi6pPn5dY0ZujwU0orp8aTrmxicDZfX3lxrOg8
CKF+jWcwd1hWn+FqEjtJnJfT9r8ufEwD0f2Llo57ThKa76w2YldLRkUyqlLOEUmj
U04fnZz6x69s6DCEtJQTA4MWAHeE/6wE9D+Uq1J2EBGeIGX0P0Zd3UwweGkTh9CA
Uw1/5zqz+ukYjZK2TI7zEH4BHZwlrhj9wHiuF7DrIrKIQCMC5GpGbPApeikPrOGY
LgT8XP4dRtswhVE6sl2JLzr6gSgzBm+xc3MHbJsr8mnuVs5papoUsQVT2vRkTBOt
IUSjywzk9iOrzDi0oumZi1dOoVNFo3mMLDAJJ7z9W5dwtKJZmwpp3Gtk6R+RPMjX
iOKcoC/e9aiNfi4nImFEvwJULjdZ0219bxZQamS7ah8=
`protect END_PROTECTED
