`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V+vt9d6U3P/PXeMJfoTpcU5/dkY2GbXXeU1N/VxiVr6AG8jTNJ+WeWaqOegE2fCd
tk+cEKefsNgTcRkznGCmtR15TFiibEkLw/KCHTjEd0d06UWt884jCjuhyPeWACw6
mYOOu51I/EjdqTUECP9OE8mNLif3tolP1TgEmeowmicrjacT0C76vAgmPK5nxyw6
6x1LZEuGNxLhMJIccM0p/448vjvJxmhHt1oWP8EQo4D/Ssk22qUKjOf/eASWiRW9
eOenz7FF0JdybRg1B1ccny6asth3acQFHXTeT5S0yojg+ZXZGmnVyskMe5fd6TfB
pGplbigKcAl0Q1wonvOrxIkrUB2FCTxHM6AlILjgrCTiRHZINnO1f4qTJLo9WbSb
4c7ys62jgcTR4Nv6y3cZjHSqHM4uoblxyl9K2n7mKQk=
`protect END_PROTECTED
