`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KI/CEwMTjJqqrms5VNXIPyoBGyBCzrGkmofdPnqa8izVIl5DaYFoL9jJy7Q21wFM
wnv/14eUClitiajYGu+6885aGDvuH4CNSPPmaVRdMbs/WEs3lUlG7hPsMgKfodjg
voOeb8D0kwOtqrTewbCWd77bmGB19XhLJN/8aKzGKSHlZHDO88DXWenlm3+HCyP9
vDrryCY/Xaemnd40XvN5qaSE3TakAIgw9WWd1FUYj5tQ9LVB502gQsCI3T5b/ux4
W5mSgvUbt6FazYnJ2Czxow4HqG6tYbSHpYEBMEIQ/tXHLfWqlIQNvsWBt0dZeAav
kva5SNjVPkWFo7pFZS2RfhXcK96itJUvigLhzGBNzygcjjON0+KWjBe/BTKsNvhf
Sk1TPkj0aZO/xgVfxIQ3KRmBvCg2B3AKbmvEV/dLJ50638Qr7lH2O1iSI6nzggKW
j+qnV5PxkAwBCtU0oNMlqlNPz4K6HxEs1moNEdxenEEeseSsOipRZUtQOk6HrYe9
rms2UacrhAsbwX3ZaXF/7jhub2zvy7xqV+LVNKy2LobWHqfRPjpJiBzdU7cIA/2u
o9TeRS+mHO1xV/tMkNo+GocSdJWZ0JRtCe4NY3Zdb6dOYsTHqt47YdipN9JCuweD
/RCVUjaNYkgmSiJ/r76enA==
`protect END_PROTECTED
