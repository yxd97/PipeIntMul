`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QhLPhxyVO687orlwMKDR8O22iEEEdSlgGQeQFZlZ2x83N20SdjhsbgEfS2WHQGnz
766VOutYkto7peEBWrbq2R+9emAEGKkuV6E19WLGANjHOPF70xEnqnVQUUI+t1ld
vt8QhloNiakmgxvn5EzNeHjAaXMgj6iIIgz0MXo0YCQcLDRczlY+9/9mfZLTzcZz
pg5oogHnRzwObmr9X+gftDwMj49a5fkMK78mWRcLASJszOF+i49U3bgyiye2fZoI
fmB1MmmUdyHY7EPl/SX5QrADqSM9FG/QeO+ND0xGd9pXsHjwInYrs+JpNEb7d5QN
YQWnzZpQ9OYFyIt14+EyJD5sxQrVrIiZ3q9qzlJQ3V+5A9Zwu/GmVjFLOVJfFRAE
LS7d8YPiqc5eH+dMXTnBJG0vqkmbIyeZcF/8B+fAP1n81qEj19As3lRiQZ0hZWBr
4KBCT/lE7HFmI2bnqCL4walAGWdyijD377VHWPi7WphhyitvWHL3eqn8O+S7szwp
cNpAzw1GhpJCYkIUJqqzSJPHptjvqEvDQ0cL1i7BaIuFryKe1HwFHtilFPMddpNG
6ABlk/xu0Mnfl6tkhcwFWoTgEYf/dqMUXmlb1GU1iJh1YNjsdZBF9/eQI+BOaiWF
S7HJy9FeWmERur/nw96H0inZpPM5Lf13bh1VbAoWRh+hlioQRbu5pObwQB8Mm1Gp
GCmunhys70dtvt3WHH9o6SEvk+CYAaCnMw8JswDPDkyJWIGnW8ux/9N2SLtq8su3
63jbHbQUxnk7r3dOb80w95mVZK3i+rEjgLlXUGSGvA09vQAnRVwG0IptRysqm9zJ
Xjz2f7ZhHhcKPiAlsZzU2hNroG/yS76nFeDAM83ims4rwrySuyTxbM6aIuaIeehZ
O6W68IKg1FnrFj7hcoQgCt7ESP/NEvXmagUaUyGRW8A6XMI39I309kMFSSne7Lxn
`protect END_PROTECTED
