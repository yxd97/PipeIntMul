`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DamikvATL11YtX/uwjRrM3h1WxOsxPbxWrkza/rJEQTywQI1zExNoaTAsaPL+p2a
KZxcZH/fCYjT6xkaS3NbfnH99G9iJFI55lSlQmBwu1Sv2+5Gajh4dMl0ZRw3UMPo
JRE1b9it5EOMNMaI4eXttUwCz23gk1SvXYWtnI+hP5vCY8GNQDZ4Gcxs8n8K1J8s
sQ4tE3/KUVt9Jh16nyHiEKHBBaG0+80cgVZSc+dmKOdCnYQg8LzOPPc/WX1KIP9T
5PW71U54sBc/p5HAqsC4K5b8aCyf/VCTPB2CpcrIjB8fL/+NCy1Ty04wT6Z7YMco
ch+76MBjRtqDH6fddqk64pUDXCJByjbl78fS1LiUd7lpxf1MWBSPUlbZ1gSZJ3vN
Bag8uEOugTxAEiy7FGbtaryH/ceSSfKcSGqxtFJ8l0cxoB/12B1dYyAwAFQwuyF3
1myy7CHtF8VRMS6869K2g3te2iu5NDnPYBgvHmq/Yy9186EZoL1I8Lth8MbGuY3U
9TrR+bg3CvCe3bBGVh6huKU4xw2GNSScB98C9UOZMzBr5+WxawKGKzWnu//hZato
PKfV7lF2vpL7RNRSMPkOMlZkElSUqj5zZ6rT5yC7yT4sKq1G7Fde1EXIfO7NFaqt
dv4KUh1i8xehMglII8YcQ/OoFcgZR/wM6znL7NiB6IkqdNiiH9wPXKwES9eIc1uQ
ec5PaXx9F+1I2fBk02Ph1Z0nr1SoDWlIUZFBJqRLakOTLZcCvNaOIaa3GGngq013
AOPv1ywHiofV+RWhwhe2FamtjPcl7V2JsXm4ulAfM0mwnqXSRsNJQy8TrSwl8pP+
KNYAq05F/MMd+hdhuabnCoKUgT4eJZ0ZM5YPeVWkWuSVGNp+wSF/ZhggQqgv6yNd
dAT8VaBKcMEb5aPpsZC8eRi47ao0o6g7c8ug8LKrXWpGTEkxojJUKFM0DFWIg3sH
syGO6k/2SRzQfYDU5BK8rzBCn5ipE2FQuUHpoIayicUTlf5POabVls8PEGQTgDkT
fxydbjszLMXv5SdK07jGVcxLIRLXQQ+7ie+avbvwO8kgEmbqN071AYUWnctR5ojY
IkUBb+MorhJCbfOigNC94sYf/prL24cmV8dvFHSpar8v4TM9wWFhKw16EYJ8L58u
1CHHWj694xfSxdAa4M+jL2EcP80TX2r/ykDks1J6IWG/HwYNTb0dVkjCP9+Fgzov
j+UEQTcPeKDI5SOLIIPtn4o1ap4xgWegFZQE2jT9MTUfrdwZrtAjAL/ahtl0ytOz
ZryygSJqQ69rlKSUl5zBB8Vwt29nLLp+5A9TUtIDg1WNoWdl/iqznQrB1Uwrf/J2
vjsZuYn06kAE1tjEIwR7xU84tbCphTanh9Afwx0R9nrq1yPg83usoYiyxjcpPeZI
/0Uc9ol7hedG5I5y2zO9UVDdN3cMsvzmB9u7Bl8dXE+iiC/zW69xgi6cvDc2gPkN
lgXZtnURS7Pm1zYmqMM6RerOrJMfIOu5OswusArX+TdR2intgXJ+6zVHJmaONZVE
qer4zZeH9M43xO1w6mmUCQYR2LYzs1Dlix8B9CGWp7jy+1MUsDE3UdlgxaTQ7CT8
JMol7P0GIBVmZ/TtexfcYXHrJCACd7Xq3lRz6Yy4DRxIM2aegwsxaXnO0bwHrW/9
yifEMpSf+cGSvhMpqo8m/+zFoMRNBUVh9BcymgxdxAsO85qaUeLJpXcPPKxqzDrt
EmCJc9m1I5Mf4K3CD4N+J2Dlhelm+RZT2BpvBcKcx3g4jALCJ2kbSR0t87fcgeHA
rT7tdbF6xzZNR/8YQiepjrD3/ME6gu2gjEf7lkOzAEjRg5E5LOz6XawgwBUIUSJQ
iQdBSE5q2/qxlqeT556TUXtDqHOQiY9MNTaHuLeZF94Q4WNxDV/ej2goy5WqsER8
9mlmahpq9Yaxs0DIJrkRLzyqDLR7hsfHQn9sUSu69FNBXSJpZlDJNvDZH/NFRka9
KYyqIB8OZjBBO2Xu8ppRP8FceFpjUykFhgAQt07Tk1eFGbe9MjMiayj0EtfBlecB
USKHDxip5Q1FjSwTUyMRZKXEt/SGp5duZ7XzawxXkfpc8VAD9u1kx6w+Bu+3nfBL
SVp5uv5iYcplAmAiwEfuU1w8qF/iqmU0zq5aOWM0DmzgGxE2TAKTnHpGag7aXRu8
qIUBGFYmfzID/O/53TwJVSM0cPjg6vlscFIrOs1mus0jhsY7bG3VMh10e8lDtb0y
Oj/8QdBm5j8LReAcZJsNqpI1wrZ8U315v9Gn0V0JHr4wUw8aGBtW10LoIO0t738+
Z7r1MdAQQtf+w0jECxK7lBiCof1zM9zQD/mJZVLpQi2D2ynNCjtVNfH4vDFJIG3v
KUBO33jvGlXVOM7ghBwoWpMuSvC0C+OFgXQEgqQ11nfQAeVvmGn0UxHe8iPJWFyy
0aDujZMmzqwRhNL9deJcwmQ8NFeel+JwdOb4YzgBUF1doWGl+wp59RFp+ekZCYTY
RHJ/fsLh1e2xuLfCk4o1p6oL5CniuV2L18bLgzCp9Q0qBxEFe66Nq5MRKV5kCLEp
2MjkqKy5biKug9hyuVTHiDhSplZlGt02yvBqpfiyfbfZ/Gy+dy47SVq7briBixZX
wP4Q0Si9db0zX00RC9ANa5pCH9gdCpdARFAOAeRAyenTp3yaVpFw8GrjUw2k3Evi
pnJ9G0UWxI+Fxf3TfHMQ45fCZz0mGk5WHZBjhRFZwLiqF+JubrTSYV9rj/f0RM6r
JM8qKorqecdTB1JRoU/9TMGcRQiI/RgsXlpdzwo6C8Cgf9uw0ssr4dmLsp2yshFo
SCwRXpBp3LxoBIh1EQ3K1aS1CLNT+Z1fVpD+f6oAvQ0lp7avov6jZBsYpQaL8ENQ
NP5mPP4gBXZjhgUvd9LiZ7C0BczB5krEQxkeAeZaIeyx3X8pZd/1jrTsG03J9YXS
KIeaDD5AJMgtTp6H5m94KSbV6fh4DInu3q50aJdrMmN5SYZo0bVKF1EGPnUsCQiW
5Zv2Or4OxjPx5v9pyH+dqipFYPPZCRF3BcTdHivm/XKjxRKNo6K44zy9bXqjorIn
ZWvyxEHiacp8qhnptTuUWJCE8ARgL1WSG1WsopGyPL//RowzZ459azekDGqCwavJ
ASyigU9rNkBkMEmWdOBZy9XWxm8U30brQ+692+WO5DwK+pVCnYuDPMY6SAOdSpif
O/hEcolPubC3ns7/gtS2+G8xlw67/pT5MsoTCcEmvut5GQ+TX52jcRbt9NqGkh/m
Uu4HdYfl4Ty3l17wkQjwQnnJIZgKEwTWIyBSlVf5Z1vdc8lmgMX1A79SZmxT09t/
PLGXZS4zU7FooPUDt55c+FKgemEACT3MLpvQsj1jX9zew/VpBKp3SCiGRWtGvUub
8+8mkUceXCym15OWrbyolQHmxERwFBLNaq9ZPBPDLrpHyrKu3rLqDy90zkFpI2kC
mf+SrjJwcDQ4Ko5IqhC1B7M2eUZUPIvZYbgLonBjL0SDnJyJdX3vJ4waKQ1VZdPQ
YJeht3h+WUuuL/WL8vNvy9ToIalXKxxinazbZAXQC3JtAbWGKOTeG9UbXwZDabl+
WWpUdf5eFgdblCFVT7/DfbUj4I8befAmbeDXY9HYrvMKBHxUy1lE7YrYLmE4yiFf
DKkKo6yG/pvHp3L4Ei+es6U9AdXF5o7d/je/QOL10OGpV2Lfb1FqNkqK57NTBOLL
GkoQLGujcm1poA3DXao08hgehmci/fTbZTpuWZ86Hg+VCdDBd5meOal0ZCXagzUh
T3pvYNDkHacTafTR693NDYf/xw1LAD8MI6ZnfXUe/V0CAAinCCshcdkM8D52z+OR
C0C4MTiUA5Ux01PHrBGIAhLeWvc4F9YhFjuwfHxLg7bRFvK5GcDBR/E7hqc3ZVyJ
ND5nNdoe7ffmYUwbdSZ0aU3OeNyQk1taDCVooSHUBufcRc2iPEgASuq5SoIo8u4o
R6W2FFYM1ArbmYNwToukzQ0olLpljURJH6foTwu4v16K+TzWvqQg3btSRPgPNGBc
PN1OjvUB8Mnv8HM3dYDP7L5P/w5ueUiJPWF7pZLh5w/Jr/e8mjwupEE+evxT2pNc
VBx5DZXfIrZlG7WO5OO4a+D5FB6CPIE/5ZZ3u6PjSe3T30YY75BwPAK3jFer9j+3
boiIvAf990HpgE/9KIOHI3sNUIBNlVNafuzAqqNbFspcUeZh7H5TpksOIFduHtwg
ct8CPHnCmGQYZrchOBvl3OT74qeobfqQ+Q1e1kDohbuGjhJEX76XE1GaZ8UICRYo
CRc+P9RR6LR6FgmctyqwwOfLDqMBtvETCHulMS+nscVbFbAKFcdMdEuT3SOEaCIW
BgIpUPRW7eBAPBDae55037fQRTmGXFWD5RVe7oUSesdYeJWipfiGFd3hbj5i3+lA
D6hZSQyGxagXAraV9zXNldXBF0gDFTfC6VZJicbE3dMc2SmqCEAjhfXqMk6GCFPK
pQEgFfnHzUt2/ajPjEYhiOPpdR5yCCSjn+KMDTIzArP2A0Ng+5qsn0S9UZ6dHAtM
vcd6Pvsp7y5p37HdQhS7VLaZh0ur+y/89vwglfFM2OtFnG5kYz/tIHcwsGIW6/GW
WymeF3hPggwuB1KJ5SH+rU0/ow4Eu4qBwjcw7lDAcIv3md6Mie8PAEAclBXLGkVA
GNqKB46ZcVdnyLqQmgDtZY9qIts/pQWdQh9CqaMAdY2Zlr0LKGG0fZvQaJqdKyRw
wAJI808MDovHZ3jYYzI4ryys/XGDzZ0bWdagBao+ry06yWXOR4gzsisENKWCoWKs
4jdKIyKTNCYEgwNS3tWNw+Z4Mxl8+/02xp2exUGwyNJAasjNnaPXGs6s9DSgQTQa
94PQL1SyI4vEkInKFKgH9dc4SulG1oW5Fp0+zWvStreTgVfNHYSNgkohnFfPG4pC
FHARHx2X1vYLA46r8OBlNeJMjVKuyA47V+596Uvt1B54HbwAdKshpLYwTMbPDHhD
NQ0y/Ikyh8WMgYXagkKIRLzGPEaYJdGOUzkt50BWWWzkLSj6eyvRmIcDpqnaDU/r
XD+pO9VRrwO41m8a0xZQ3g==
`protect END_PROTECTED
