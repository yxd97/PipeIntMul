`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lXTEuPROuHMBsIGCHygRhnKUn54fAqmU4Ly9wp3+T52lbNXiXVOJMxJ6pA+dQoLA
FxKEIT9l6+x+oN45dSptNl2CKTfGWDgfp558p6y/hagHJElv66zCgInk3Sk0RSFP
nm+Y5psUKQqHPLSyV1Mc0qm454GMpqgr1ROrau/LuD64Zifk0a4c4eQ5VqKea1va
AeZRXgXaMnwSPpQJjd58MLeUQXKQ70gmhOvJZnjWSlXxdP/R4R2motNYKG/OHrwi
dlJg57bUvewU5AMldtoCFS/4NFsz3Hb23tewpxlHDpGsNdfqgmoTtmwvL5Njboe3
0yM2z5zg0wOTT+LaCSXHsQ==
`protect END_PROTECTED
