`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iCdIi8PqtBxrbwvMCq8uldTCSLFoyjMYD+k36dTeuDN3msYKOGYx9bDM56b3Ch2w
um+imTA3YUZap+0N46ky9Pbj9Y9v+kUpwlJJ5lgUbsl50rhbOGez780xJVLmf1CM
Wys0USsR1Lt+VvuQ8PUlOyMv4KRqP7aI61W7jiAkOk5+0WKz+CFpTkspqUTjokfD
grj7p14P9Hz27JNePuzpZHg0DLrYR4NR551VRRfQNJHaWbS14gbplulhih4A8sJs
bauyv0Ji6XYl+4UW4GJ9VQEBWVl2J+hvnFHq9aWFmvf1cVB/ufYT6Is5c5Ry6ubh
F6t5xyw0g7o5KIIKoHNWDrKYVdZPAJR9jupp5g7zl3717vqhzgB6xkELNpUMi/NZ
R1gyz6/1PmMHaHH8b78fvTgmYBR5TCSdBYxy+mMrdCg=
`protect END_PROTECTED
