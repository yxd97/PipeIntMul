`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiguybPFvi+JH1EIXnklB0UyqNpo3n//aSadGAQHkzXATcJKfZ8sbd5Xbxa0hiy6
Ol1LaBw+pgeWLUkOAVH02k0G8+6MsbJH5bhmW30v1rS4EOKX3+oJ+G0bWgj2F/gS
GNK2s7ox9jcCE+NL5JydGwyE0axWXvM8kOz12rm9xKy6K5W6MjSgaodr3/6ZfIEv
App6hxn1qF9zYP1IjRA6Zf/d8nbcF5ABezE/D/1x4+8lpPiddnAb353KRM7m8GYp
kexr5wkcdI7Uu8Tr0v3aG34e0a9+RU8lXGF77l8chkC/VDT5WtNN+YM+xOFhKBvo
X5Ziy2IeAtiNQUAKx+2PHk2qWD/rVWTxWW/72ZmTwfGNg+b5kh80gA3i/OCh8ZQl
yvyiyzac6AkIBwhiu2GGxj2CVCKEc9uJ+o5TYdSkrwL19TPsUljjdAiHo2j50kJq
bpXIqS1KLULuEugMkV/6rNz/6vhVEYnOqjV4xWLUOh0ao11k0spVGlVRywkzBsRh
CdrtR0YCT9A0nqHNr6PhNfMdrQEM322lqPPfueqRj6WjdETjcnu5o1YihLeFyn5Z
YgPYnB3oT4Abb/+C0Iu3AV2v9RJuvKUExQ2cr12uxCPRPNWPx3Gyn/U9VvN/0cHG
zGMgizdMlT6aPqEUPdBJ64YK4yWRuS50Gbd7UAvM4sLHnJpSw49I0OjGTdRZTT7B
AIrubaspVpv67/JXW6Q/e+3aIz6ieHnbqE/ZrTNLTwwSe6ZM+SBPyZPbihBTZBPS
kKyWzbyd4nMiVp5Htxh4QW/gquUQIVWMwxhH4FKPVOErUbnoWuXKwWWMKY8zmHuI
EaPhM44HhmKnwZDDCGFA22QPLNZGQFCoY16sia09Ski1UDasxklvGcEgCx6/heig
keioKlO/2Y+yknbRhI5mDisMaaX0hAYlT8aOFxxYC1HEED9nRTWUGeTIWEZGnxXd
PZMl0S5Ts1csr3ssoULXhaD0uetCvQVMz0Yq1a/bqwBq2Ib0S+ORwxMmlkpMPpex
Lm3s6SC0VSzEPj97kWdK5mk+N14tuhZ5FtaqXXbV5ASor8gyrV8lytkkYcB0cRuy
Lpid+FG7JOQF5FoE47fn5FMcQcGwdMn7MGYmIaoPB4u2m9z2zlJ4GWhWyg1LBDSG
KLHw2qnVQagNf9uqp91pXmeBugGmRUE2GcDnRVvIXz65GLWIVWHi8KfTJ6V1lC0r
caYlNORRlxRglAxHf4/loFu+1j2VO9RFpkxrtoFvRERURRlWVKbRHU0Ji34zOwZo
VoYPoV9jI1d/CVIawJrgJdYRjfGNG2IsEy9jRhSxxj7vjmvX9GeDb+Llr2WXOjc1
Bywk1zI3ZrqerBk+VBdGrzVmRuZ8emN9SmKbUHuGQojAgUWIF3JiPYyCXNCNJA14
nv2xr5Yf/WrLR0sxyD5UEjSYLHcOFAGz17aHDTPrdfa2QV5F8e6XKHtEOQHMOL9A
O1B+SZqtqOMm+GeA9U2EXu5YFLCWv/mguupsBQWqWiz3O9jwue2S33xduFd0gDUR
LsUXnFYRMsIEN1A7nof1gO2+GLKiYwFlOhzoLjo47zlRkfCW+/5eQZAzbKsSqnS1
yQfs+TQ+mXmV+fpAv7mCl3CUYZilE7K7jCpR8o1zLNJ1BMDi+jyVw/aKgl67vw86
DK7CY4KmGbxcaQSuQOqrLF0POEyhagdANS4wUvg0OzN9CeQBGioSzLGqSqGRLpNM
ir14ZfDmltZKB8M4pV4I06LKx/cv58TXPcg7IrS9LHE9BwUiVuPqHVmmxO1huDyH
f+NLOH/oGXJleYJEEnszpB0TZ004wYVJ/eiCECPfGIoTTLDLiI9ibkr70Wa19aY5
wZ+RfgefLV8bfRwEvwMswotR1J+JXxU0CF/GqbFI+t82WD5NpiL200bf8SLGceno
`protect END_PROTECTED
