`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
do1a0Q6KKh77KiTD9Ve7oN5w+wfOseHxadlQTlP5NfNbBZkUkQ6eoeEHIAPbG+Nl
05VlZp8QMGktMuI4MgijxKO6z9Ui9/U7tlx1K5JWAo9O3kPO0iTBn80SBGL9NOtM
/uqF0UU27Uyumq5Nsm/NCicYyM6aHjjpB5oMpJ9QsbmoW5RbqOwnZK1QH0/Rwrbf
ADctunI4hYc/+BtzwNqejMucMbcJBN1e7/qP5kUgUYo12tl0usXL6tY/d1F6kSGo
bqLfe3gz8qS6x/HYXtYJROSlAsT3tb4Xuw+UihV0KVkkBvY3i+8bTu/bWL6mkK9b
IFFzw7QBO0utUiJ9ZSa3ty9SzLaXiJqGrUztHZr8WEbp9uT8164U134YSFpUlsfB
09w0cuarpo2k37RiEh3SpBQnVoeIFxdVIrr+ez4meYY50rkjL0hu1valj3wQUbj5
+iuoPkqFWmmpp0eL9BipOcM/o0xKHZQmqGGGgp+JboY=
`protect END_PROTECTED
