`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iHYM4PKl00UoM0nZYrWT2jReCt31zi91mvRtS+/AG9XAhKi4qaXt3GoDwgZwBa54
f1fkvleuX5OX3/yoNAJ+Q94BVuKWAcYtXFNRYWOq5BQAHE6yAz9VLagfae1Euc10
dcmUsa26SJpawKVf1+v7WMVLkvLBuE/7DXLNeKCJxmhaLaOa1eJjzllYJsxY6jo4
K1ZvL8r63ov+obiQ0pn7a9YYCP9Niur899ksLLp2NTpvhTLna5cUY8BIh13dQIkb
IvdTtmSv4V8mEGyA7yQu0L1lIAjvW88TJdeCItX6KvA=
`protect END_PROTECTED
