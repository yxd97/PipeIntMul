`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jISX6cqY48MFDIxoOq2Ccm5Vst2dB6Xoo9EnFNlB2tvJGATNwOXogBd6AovXudYE
p0d7FHGK/H6p5+XCQkDSKlZ2AC9xwQirfzrOe2qZx/K2/FhxBx27S0YGsWBiIkNj
4EsfGemqWshyVIQ5PEnVJxyAXocjRMo0J71H1f/HoyMvpfEGbWysbMd+eLSuk0v3
58c5X16smw5nvQPReIm8Kq/1gspwpXWSQYmL3dSm7KfgmYeJ6D3nmqAxkf6AIRAW
`protect END_PROTECTED
