`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TPDFQE+GtXCFQ+rpOCzMeZPll7Apop4qm9x3P8FxZr5zryvb+PxEiougMQsmJCnB
Lgq1G9pd1cAMShUXSh4R6mnxakgNIyZLDU9h8+azGNqKUcadBo8HOie8x89QQM2y
ytGPDNehcmy3HrvaxMT86sNCnpLFWeSnxiKAzyn1FGRYu8hvzxCBBPhO8AuiYqRC
k0WniU1wOGtfJvwwmVNp6sf2CeZMPrKJDMVKcgMsYbUTFlm8FZ2bH3N/szL7d6xn
fKrJXpiRUeO4iYLQKan8yrWr4GYSxWk70hlHHEj0XEFTQtOwsL9BLokuWxJpAQno
3fn6y/Me4K4MuyAmvzt8RIhUtwN4gcmT1gNNqDEdARvFLqLsSIJkYejv1t2bbNrP
I8Z701INev1QFMk9EXob4st6m2frY5Vhl9p6GALfYDE/C3qXc+1hUuq2OXkGrub0
cLA1bAV/Re6Yfe8OS21KPWCJ0GVOObf7TIHzm2wOOWle2jB5yfXv3N2zAmw3/ymC
4n8ZU/gBZvRVzOtdooHT2N7p3d7jR6LuEHF49XzxP/gC7cq4zVpj4XQRcP9Ns3t0
ONRtLAIHyEvl2nAxJgj8NoZcnGJgbRLwkIkIAiyaTUXWPczcHVHQ2rW0fV+sutro
5Y+hLeTEqAwsvUWDW+cuWGkyUfJiBFk6fbvQ2iOopNjKOwzT89CDn8K6w/9D138c
/R79ADAX83yUTbAGKlf8Gdt6VHJ01WG1d1Xr0OEy6gGDs8NY7cyFd97OobiFHgdM
RP/xHK/AzvE5Axl/MWxrH3xFccsmoXRgNQs75EhBQ0UO5FLfmYa3If0ROgoToAIa
6aPxUVaERyRCaa42kl3jrg==
`protect END_PROTECTED
