`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cbHAVZD8MCrG6uyd2DIG7KSKqdJsk3Z2ow00W4QEqEp4VMYn5EkSBK2MMaTwKOr9
wc1NTNGyFHyO03IaNwPW1FBS6rGdMznb0ufC4nomfe4YFe/2fL7tt2ak2MLsqSoh
9At838BPkXmPlb8r1xelNzNjLNIYp0cGpE1cSoMWEI2HcAYz7uCLp+rxtLuGpJCl
ekrpH1LqBYqx0Lqb9KgflquiNo0sgW3n1E9bulDwU8tLrVl+BWn+pClqmBmtsfQD
iOeYKJ3bM0n+NilFTUYP6BFwIZYR6418wB6d9Hegnt8=
`protect END_PROTECTED
