`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gnUjqRWVKeioNVoAYgz1G03G3gCjqIGFLMZ77mZSUAENCL/DLurjeBv/qV2hy1aZ
zRTxLBxTNQE5xhAM0FPjC29OgsfHD+MMzbj/Wy8/FapW1uEDwCUwx9R25yXnaz+h
b8UPBlVJfS3/weoorXaEg8BKUJMklEGtRWu7Nvu9IGm527U1zArGXvX0eKzJgQoB
WIL/E7KVXFfZFfM1Du1oFAazG7u2WxFL7ETpLIWCQYi15fzPBYKhcDVYr1B+TT0u
MDzE8Gn6nwr90+7HQjvpyw==
`protect END_PROTECTED
