`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9RDghc/H8iAYJrkM7LIcT6EIVOZOELXuYLdb4f/E3jn2kN8vlRxgkGuR/M0jratt
IBiE9DJMoMPrtUpQLRvzml7EMA2YO8kreoc1EbU0sLCgCp+TxYfGVSVH6wl6JNfG
mTEfcvhLnN0JSwY7IxV3QcjR9SOZbbxw/aFcMZdveLNRPD8iJd59jdCU9Rq6cvTT
WM112dlGLZw444uCptIO12F8/hxvI1w1Ft7TRC5vkOLzTxArjyBssJyXlp4SRuzI
y711IPMdrAHXMqo2j5r6zFe1Rqf1wBAaaveHd2ZYpaQsFCgs3hPAHA9jez33b8a7
4MN3fyhx6x4rw1lH2SvDit4Rt8f7JR9oKibv6GDV6u4VsWdLX0IrbgOx2ZGjZFXP
0J1PeCJ20uIZSya/ouQ05ry56DmQLRvsRAbdbeJ2JUo0JrnozWibOi6vlP/tORd8
Jgm2NtWXq5xn3+QHR12UOe/CZRFtCQs9UYyaPJSFpxzBwzb559irGkoh/pETv2zX
WPJSZNMkQI7euKgHXKBC0lV3D84nrBWiKxcUA9xCMDznKtz2IAvrjIGu45W/gN4S
0kY99vGvyU61IVo/PNfMq/g5gs322Mya5IVS/Vn18LQPoslyZwi2hWzFBocR/z3N
JYQLtOK0MSG7KLrSJRPqi4WDWAKzYkYPDQA2SqfBfOgk69KZnZYLQOzRIm94VcOZ
b3RoTeSVbGL4gUhcZH6hlHDxgEuTEHExgED1WFqbj8T3O9PXPsVZ5fH5of7h1VZQ
qbcxkLinpj2+htn4YPigy2yaochWu44UBRyhSv+h2py+qmBL23PFAVA78lAuASMO
tJnl+q+6ED5H2GB6aDgoyGkQPqVOODd37GMCxMzmIid/RgnRf//ZRF4q3agK4U3B
ZFYKK7c66n4Lp6bIucLejFH5QVxh5cCbUWAXENfBVlfqkUu9Ql2vQMKBdWORNEIH
qx9MHvRxHeDNJFxbssH0QTmmEO1gImkD2AFVvumNt151uImUYxH93z0lWm7CwrpL
N0jFqaODiMVVQ7FHU2wuv5lBe7CNp6E8+imSTd3sNxdPwqYj/SHwS5gTuaxlT5y4
hM/Inu4M7gSNallB/Q6wA0fWA7xLzDDQfzPZgUNmIBMNPBI1no0EPt7BVihAObmi
QUXujQSnZc/HxKkeAql600lRqRO6mWG+wqXsRaww7YpBg1vUIc9GNtiH2TkjBc0p
Mecf3mws+q0ivPU7UUOQyj6afOd7frPsg02GcWQUXi+lC8y7GRwwr8m92EwcCqzS
f4QLlWjRkSvO6thNviDLCe2pTaGEUtDXeiHib89aToKhGFd/aofLxPUUvNaxgC0y
HE5qxLSJITEpEUvDYOCiuspYb6ZuLmu6ZXGgjbILIEVxZ+H+cMh5oc6tMjFjdz0R
rQLP3XJSafrZNQaTbTTBx0RRDteBElgPT4DeQOUSNb2PUPkwQkoT6rrrChCF8auV
lBLTj/NmxnyauWW0UA5C0/RxkuKDNU2NOT0AvWEbhUXpbKslzTBrtfkxmeWrj7Sa
WGwXmbLaukJyniV1O2ag9BVIno6YbuBL9ZQDFzSVIdnb53GD2kxR/C+L1OS42t6O
`protect END_PROTECTED
