`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tAk2UeaMdCQZ0WvWCJKKoBYn2tOqhzNiOyUaidgmYZLS+i6fBvmT9ufIj9zrV9E3
ie691vsmeWTj/OMJQ68y4dbm5Rh/4yyw7DfIdsW6evpNPveH1IlZDp/T/y6UrzAu
JC8P97TmRUwuztuPlJUh0TfrzunXrbua1WWDh6jV4k/EpLdUuiDMNSJMxAM6Rf+N
X1pcifuAGW5iYFEiXXQc3+7Rv+qhLCNISGGEuDd3glWPQisBjentxMmjod/Ku5Ck
5x4riAi0J1XjkkXzLXYUx39QuMHkCxqHVw9gPYP9EACezYcneVWtVjfjo0kkPz1r
cE1T1OP4D6yEa21q8N4CKeBPO6viZo1nUiHEDbZF0O8EmATab/3LkQsrITWJdxJ2
SBaeeBneovbvfs4z9NwhNdLmVmmu+jik5YIQSIwmxZzYmNFd4nNs9Yym3ebSjbfN
bTztxymf/l3noxPyfN8mi8yYzAFKJGSBn2++3bL0xdqRLnQO5hImdCW6VGfUWovV
N7hReECOQHyCTM4U9icdjtE6s5cNSKthtyS8rkDExZlsjynz64PprpyqNoGROdDe
HS9yymJNw5svYyXNE9DeFMQhnwY1KQrfmP/fb4ZIazbnsPhl5CQ6VYQynvEMzmPI
FnmVPNaIrS4J9l1dX4Kq5w==
`protect END_PROTECTED
