`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ar6x+6PG62S/pR+tuvIEqOeRdRDrmhdZU0IYKRcM7SirCDYDXGDk+iIoAbcUVJwo
vgA8K995lDPA9QMju8d1vqBkIvs2zxliFx+l9hw2TRtDMO7NT3pu/BONz0/beP7U
qwyZzePIRvbiaPoZrLiu6WXzeTbOQi0CwPqlfNf8D6Zxs6jfv7W+J6bYb0WbhFfg
f/08D9LZJ7xNlYS8Kh34SHP1NKY1AKclupphhBVFzIdIowZnks5zHP7H9QxPRe6n
bq3aYD24VsBOlmmVSC2tSPwHNX8X2NZcsuQos3FY7fSRQUp/PMRVIEb3tZ8+50C4
kbFJTBvXcSn/k2T5UIfQd1Xj60Qs8MExJYeG0SIgi8pVj33ISWQdVLMtUYUVBmkX
VKT957eUYSUQOUThOx+tG9dsfn5I9dPYy9jq4+PIhrc7nT/KxfD2GYaPqJLtzuRU
o6BTtvVhvW8JF32fHEOZ4A==
`protect END_PROTECTED
