`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZssAElDP+Rj1w7KbZ8rN/8G53oezTuxBXM/LEr1qIqdo1dAPKAVLbyoeu8qlsxcm
Z41AoAUBJ2l0LPPvuG3Gmj/LqhhD8OBuvx1JQNMKehztwSrMmdMtnyXx3/xidpxB
0PX4XZbB7E74RaAWAPc/Lf6n9u8xLou1Ok2KzDpOjYDpjqc5jURPNBgfDyWiPogX
ASjDvehk6dLL43c4HlTvBWdH5a8tw1fYiolu1vA/Gxzw5T0LHX6wv/3Bv46iWX6e
pgFvO9BTiSFFWlayjadwG7/LRDlzA3NvokOJ/yGWc+UITCGHpqp5Y2VnV+yLVHef
DA1VMjyUpSSs9a4llkIbxeN1MHprofm93G0dYJsMg1bsY28TcrVLTdYQxuO1rSvR
Dvh+qpm16kRTbETqdA0Q2guaSkd4IXeIGBatXk0pmT6rPK2wqK9HL6usO6aOVke9
VoX3TMuVucrXKHUWTV4UH6L8OU6Q3Ig5lMQvxfZG6rs=
`protect END_PROTECTED
