`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q1cNBriSMxfOI1I8ws+PwZ73uplJ9aYAGNuqQLtyh1gREH4DttCTNoqHvnm6aiY8
/BdC1v56IcNODgSP7rR86j8xqaHO5cMBIuTUij9S3oO8LZpRIF6PYNiTbu9lSYwE
+ezmx8CYzieJ7HFzxlJd/w4Qcp/QU4jJety1iKb07pD44LgeoFqBAHmpe7UEbm1m
cfGxFl1/M6sFNzlvY29IORwHoc0MM5xbNVzWp+L2itkfkdIITIx1/hUEaSl8V0FJ
JDUmd8y1FUYwQ9i77E7ylkiK3s9IST86O3aCszCmIa4mFx1MMvSetcK9HqY33fhz
kMsI5YCya43L7v7Aux0nWAQT1ievwf8jBVbidKfPeogJJms/VjkBKoAYBIALDL3F
lYDTsfv4an9g4yL+SrcSyGpVX3EbayO6Lyk+mOBo3fM2LOQMYmb/k2AqvxIQFKfj
`protect END_PROTECTED
