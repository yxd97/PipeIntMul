`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
l9SCYWG2LHx/Bi37pvfeU6rpCn6/zCpDIFMarQrj6B7FrzvLqyaYpZqBBTPQnCuE
0F+sE5C/t+HsJizabAVMkK5VmYCZE/u3qEgPz/KFTOh5TAaWq6MYQrR/Qt+1XJbK
8/NCD2WiocXbjN4YO7cjhFV+jamxGOsBVqkiJ/XRKE33Vj77KuERrl+SYit8h+TO
dNJYhCZ4uqbFKjWTFfvi4fDJrmrmskcQCz5koygBBRC7hiOLcK+DhExKuy+OKkW/
zHKUsLiMmT05w/ggXXmZDcpY9TlKUV72qF8zi9EFnDpjYJKT47ek3pNW/Zf3Tw2d
UwYf9WcgnpTVAk+HHMw79sJ5BoKvqjWGoSoG/a5rpnY0M/xwUojO/QhAbMfGCsGd
two5ljW4aXNlGayWu8QwE9BdAy5acCwnCGz1/KUyz/Zegp7B6uKrV2oktHwq33mU
nr7e2JBRAAiQ/xg/Cbj0y3YriX24Rwxaxiq1GgoqBvunBb5yhkvzU2Km0wBt/zYe
suEN/h0Gre3vYMT/bDN4p1ccioTufmMoAT8G/eSHU5/lw8SGrGSIaaupCTxWlTqX
j6xEF4MXwbktnaGySzv2oT/ogPr/f5LhSyIDrbAqVdnqreK8uosr6lEgx8LOfuru
fh8PpmOs77/i46Ny/uapsKk+AQR5XvchLZiRRT+oMXZgD0SuXLF683z6ySy2T5Fa
5PLbXLD26jVPGOCWVKZdb68E1sXplpE2OSh67x2lQIYifybiShlM7zwS9V+boOZo
+8cRWY82HO5kAlkhUyxq9sQzE9PDHas8hHRZGU0JvrHXhwBfPKW0kgwgrGjoyYgu
EHtRDNh8MUWse53vmK/8WQpqJXfLuCDiqJ+l2exdD4MfTOib+RjZqlyDwUC/tH8M
o5XuExPHjrdIPtfvZtvrYPBinI13rg36I2M98ciM6rdz1W8BNhrEqBBn8YoagD0M
`protect END_PROTECTED
