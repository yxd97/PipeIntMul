`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vjp/DxcLXHTcW6Y7UpS2jVbm3/nA5xlfXpD+3wxUYUOh2YhnS2QOtx+qRhy/IiL4
4PfW80P1UG1Uea9EFCvZzOyxQJNXlz6L9PUs8eMCT5zguAK0yxRNWuor6JLIHWn9
0X9ZePMsddNbD+sLOakSDNAuk8fhL43Zk7M27zecHS3keglGhbJ5jcw9+FbLK6ZS
BRCXJmSnwXo1UBBuc/jZ3ydcLxj2DAB990A/2M0IG7t644L262uWIgsZBaXWjz2e
m9N1BhRKnm6kIxP8EjyXifYkSoLJsyRyWbtMTP1f5vuUkv6qxufXet7yQ5LR3EZY
KvXMzVBsjpqjVeKka0oOKIwc+c2Fk3Xs4XLY2YpBjQw487cLgSd1ByvIUf698HEp
NhA82yx8iWW7xlM8BrFWIxhuEb87g63nIVg1gPQfeUGXnm322nlsq5H4YktlR246
tjfsY1r9eoXulz8q5E9ZikoNoYXnib435Oo3zSmAdxyPuBl7sKR8kKJcXcZtL5/K
`protect END_PROTECTED
