`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJM3owbcRvQZ1Zii4sqKGDfULAb7OOf0QHu4nUilpyseUPv6HcaFg9YJw3QjCwMK
80HUEQBX1026l6MgUv+cSZlYRlRx8gtPB+VF5upH0T7sW7rjDYXUGIqB4zARt1a5
YlZich4EarX1nCB+ug57eAP7FVkR4D/iwXfJrorIAlxvuIMj91qFungE9SR/IpHY
mbjURzUQ3kee0mfMDZgZXeXl+mh3lGjUaCNgmJURxgq0KkhdF4kVIuYU91kpT3j7
x1+IUbfdRSFMXwUsqutTf7BA7h8VCAqGArCZm9P52ZaRiDNEsLxtRGJQLmDVRnJi
ht5YJWSeDqc64Z02QnvQ/QTohfakdGSmMeMOUEdjEf6WpSJ39GN2yEf+yOqbPdxp
XwlRhquOcmD2i0kxy0xkPtj/VYncKPSP5Pkq7T5kPTd/jyPb0tqnyKHtoq8Q/sW3
hRnAAGONUsyaHxbU4t8EZy1Jg5Hbm5485BBg6q5t9CmgZMVP/IC0BRehf94LoT3D
eX5CKmluEFzf9Kjf4FvIiAPeRx/hPSOyv7o4HPjE6Q0L/w1rzq/rK+Lbk9xKurlI
QehRPwXAwneZGviXKJdXRspz6SKH8nEUHb03Okj1ZINcZvvl2pMJruR4ZUHCcGIF
EiBjXn/rI1veqtSoCUO4YG+vBPUttv1amabrr/TQdvHVNhLCcxDNdDOeuIgeu9JN
C2UPoQ5cgPYbP7UZCeTvK8Uo7m1B2gH/RkMYljsXOEWi65LHiRuR807sYN1lKUJ4
MejqaD6EVT5yGCk9iQLX8HtcaLaHKL+iEuVdIk9qPAAViOoBtd5GB+zzvlX2Ua77
s8aev0DFkgyzsVEv90vVtUG2eVyRs3ga1bemNz7iRG4dJi8BSD7IHfrCLxI4ffST
2MuKYLZ7u4xHMEE6lLsi9FIVHVStVLSorAM/sqE/a43kHYqJDLDbtNaIH/TzwQI/
XQHdQze+3kPWYDMrutG7VwEmTsQD4XWdCvgZ1lhDdBSJhWKsZc1PH17+Z/iIPENX
g2CQWHZjFH9Df82BpT0vJwzWVeRAp1oNfp/uob1MWVf1eprBD1TBFowMWehIXon6
SbBjcRCdewM88zQN9gU5eL2bMq3ZxZG5DkwRWaKhYsc2Cojo/Ppq2SPZxOWYVAGg
Hpc7vfx5O+P4IB1zZlw5ffojzZmOSqRRVtuUH3KefWYAEyES537hm2oIkKdy7juo
3HzWBb6R0eZorFtc8084+HBq38luSUWbJkT1kNKdS0sX1BRYpZwSspL2unGJPGhi
AQmMIJIqZ/+Ocb8Z7GkERFqQdm9YR48TaY6R33pCcqLILrOC5+wqd52Yjv9ddYBf
MAjSBQtjoMDFwbyg+P2whLrXdpK8WbRJN0OIbzeQH5J06g7hDcC3dg0R9uW8D4Re
8pOIBbrSkf030xwTrWYAs8Yof4+bajJhqKnFp5K70Lnzz9w/XoRUCVW9k0h/GdPB
z9Szm3ikDD2z7eP25i5vva+u2ZT6D4L0nqkX4dGpDmlMMzw+k/pM1V+Ujw3Py1Ov
QsDQIiefdt8eG3AlSGtP3mrdnVvcLu1OTvziKi4ThKGV6VtwZXFay1Uv5Ai0MYFy
UwxMrBENb+W3+MSxs0nvF24HA4jjK1/gezyLkirZKOoc1yTW5dTRCatBaGVA1mER
yPtnAFB1uZslq+hhgxKI8kalStGWyEQojBPZruW8hFCcy/pYqfcz15fD5Jk/wV2M
7XJBKLW5cyniOlfD1VjYqORkHUI2B70kEssey9EanOypIld+pAJRrRoS6zkE9gxO
oUlmwvl9cmZqGfEVjBVYl7iQD17JgfI7I9nlCWSKLZrgAAAMpu2ImfI/ROF11PcV
Zq5PU7fesqc14IzfHaD58ix3mwL5lvcCkDquIoRCFwClyULHedaghwMhckvhRiWk
2454JnleEKNdT4kYpH/zrpR9CM8SUMOUvEFAqC7gKK0KGMQ1GSVYhLcZWj0nvWHj
+3TKksleKdR5NT7N7fpIuf44qs5ZtW/1MrBvYA1exw8PwaLb+88QjsL4IrOnrjbc
RnOA3ODe37jpJ3zieRKp0X3hUrEGkAahotgsxm6a1w+pTnx2Zid4rRrFaD6gxZhK
QgsoYJQBsLkpJiS/tY6U2kylkkh6LvtNcDQOM67+plQhqNgHbEmxsS28cj5kV1Z7
k6TPkKWr/Tkg13Q/KvQp+XZdSX+OyrqsbXE/9yXc2hoQlWV8FxwYyjJHniKksaBa
KnuNjAtYtr/Qq2N7sWOIeJLGF2nMtCbgicmlTbBdxNDVeE2TW+1amRBaORWUMwrK
10iX6JMxW1SfbTVGElITvkP3kdtrcyDnqEdAmhxZnxtR/jipN1bPkSAuoVTh/IOt
DSIzbJY/LTCdmtGBw2tnmlIpmZwx/ylM1vA+Outd3oAF7EOZ5Mu44RvVtqDYRXuR
zpPAvHjfGtn0QKfIYUdZoN3O5eefrJWpWqmXIMlRo9ZySlgxclcXISJB8CQiESEC
Rutc9m7OvD/kV9TPr2lal9Rd4jqG1fgoKiO8E+USK4gXncCK6HGcrCRalO0HYi7l
pog2ie8/VnhCigIPTXubRqkg3Ds3ynrD90uHsv2wX/NcXtbIMmllLQ39+Uzd5yrL
aa2ZiLg+7FuWsgn0yjQDRfZ2thI03+34MmIwlaz957CGtaJ/3TU4YJ6iVTccREI3
4pluzHREI2CGzUmdOcQqE914hgBCCogW0tkJr1QyMVtUzhgKGSH7l0EfI6ruMUDX
/ZwB12vPowrYPycAJezxnWn2Ljgany9aOGBMtKSJZreXrs0/2vHPey0nKVyO9kt+
7Vt6wQZ4fz3tZbiAw2WK1k/Pm2JxBVkW18mgFICgJDHiNKsuJnZJr7FbFCM2Rpug
APM/rfIN6aqIA/My302hsodnb6cuDTz4ys+l95A3RjgA6Mcsuu5niUaxsGXCRbT6
rchAFhEB6T/Js+s/UYlq/N4WFcNKKs2zhWAqrGxXaeS3X9waabQ57eXink1a1MCj
xTwCKbnDxbwTWpzGJ0m1+SBhwZhDvJDCSt51rBViUqVMpGdss3M/uqEebojQI369
X+zyC34S3c8+YrarXmPfGlonQ5YI69EicRVknmz6qrnoG6BS5Jfx5LpxOyl1VppD
EcXgh2HGIFGCaisbNZUjE5rIaDK2muuaCiCpUqTKE3i4BJmSps5pqlZxWbV+Rz21
v1N3XU2u7nOXvpQ13W7KQkWyYmJAG1Sni2ora7rPSSSKTMLlmociphklNDjtmL2G
nYVFwrdBGadw/ANX8cs1NUN2DQkQ3K8nHLjZCLBPX7HZmIXH0G6DSuJuupTQcI0r
sY1lqLj6jqNcEr4odvBTja6K6ZTk0AW0UJTsM2QwotxWhE5lwPHxxlyA5dmKI223
or0xcVXpyCnUns75PgH4O6TGBUUOmo+xlKcdDhskG06CbMdITZXyJuR1X2siL/Yj
PoPSIknxkqkS+sWc4Vb4sCiLCt8AptPi8xNBilpWJeyplg/wFnhYexed4kj7ky29
VEpOKJoSYBUHJU/ZSqja2FXoAsfjEenpZQ9yTM24yQGyAhd53gPJEigB3DXm8EKX
WrhJhG5tpkVWsxt4HPLR+pzTpTG/TvfvGvOUQ45+tHCBpjwiZE0TgytdxrhLZlTW
EbzHrrlibIPpGk06663+B+LbLx2eXhLOKPggletX26ZgNyBSVJcp5Qggxahzybhk
IYMmrlUOLzalailzSKq/2GQI+A5eF5ok6o4boRivJbiuKEaZ0au7Lff5pNEP3A4Y
kbxXC30jdkAYgTBpch4GnoXTNSZZV9ZPOcAOzlHtWg9KW/Q/yP6wcRfHI0B2AEbI
hFEXZReiarHc1cLLAdJuiHTy1lA5fraJK6kLyHHhmAbAkYB7+2vNUL/0/oNq3vas
jUgStjXG66aQTLFtgXAsrxickHbAxnVrr6X369RZMT+56rdG/YyCywALLWZa1pZN
RwYcSnLrwm1L9ffUdzli1JBr6snITU5zjCawqJ0NsrKtoE+i+4ZACdGjSO1Yw57l
L8bjDYML6oHKGNks7vwcA1mFfNngpb+T8Km/ur4seM2qLS62npA73QOK4mM3ACMR
wj3R2SO/Zx5nsD7ebciDDelfCCEGpVU6iDYQEXX9x92N4LYj2CqRcFOJERvmiVcY
MAE0UCZoBCobQVm50YICV8xxzk9XwgrZiJtNwb0gpSBXJGg76mIT9XqKNBI9LPQK
5dnixmNzVE7eIfSWujnsQ4NVC30fyG2vIETbrP7YNI8XrXHdp2HSTVl7gh9PH2zV
jDQGtVcuoT2PfE46ckcBhb/Q4xiyJXTC/ayxj7y0sYP6nFhx9kyFHDy5fGMaQPip
CiKFgHRaIh7DjuFom1xfc/+GU3SUdIJLcaS2Gme9fdQf89XSJmSg877k7tiV1lWk
ck+cLhRCP9MnbctFcz67EiNBrpQ3tGu1Wa9XmfEZtniI8AB06h+lqnsPekUtnpRP
C01WVGG4bKrS374RxFLLZ1AFLKRqnw+ZxAr8YrtH5uytwWskUzGBTJlCVyb4NPmZ
RCthN6UT7yPP6tLf1z9WPzZWR120YQHdh3dccC44NHoZEWqQ7cs7LTySzyhf705e
nicU/b3qNWvvbjRbuHwL8XDONXn45ITvA0AjcKQy+7K6vHuEOdrTlmFsEsfdrL4+
9uaJ20rK8IdndwvcE+sriMgtnai8JdVxX7fadFwKXp8kisFeIvAQhcA8gk8mIW6N
HxGh0WHCzkftI0IK07nJPG6DraowuiW6mu2WVCWouqPx1Rab/dynZ3GShy55DmQv
RlPsy/a+TLwQqCQGv0E0H5R/SKADMlPQNmE7/alP5zas2zy1VLZVbbSRAOBeMqHo
FbZCTu93ezhcX/RrtQ2EOPxqtvQU6ZfxVYwI6sM0C4J/derfdZk8E6LBbqj/dcar
NTdSk3bWX2Knbieh8Co0twOGfURilKVZURxsD0LFUft1PcoLiAJZki7a6sz5Mj50
e+7GerCIZzbtlQmCfgCv3P4QZ3ljJh2yfig7RcZftxvp0TMl4FRRv/fuQBhA7qwn
x2RM3EXGA3cYbFH6pxKgBi3Wi2XG385+DC39YciSBn81bgJ2c865QJetfzYBSFCa
VaCxRPURCA89NH+HgpAEYlVTbG2pD09/MTryn/on8V3lVuDVsq/i+05dFt3B2nQC
wQpTSwR4uwmVddeHznb3T0Vl3eepyx+WwKYSrt6eGbbeJqUvBtfW4gsg+TGIu+fZ
SE+7aF0StrhINyDPAl22CWB265gACnTlxsDIjUR9OfsmTSxdfZKmPCLSfGtzWWfm
sE8gcI/1ylnchqkMLGYMCMVNpiopyvth0tvoLKJCB1gg3iYkjMCGsowhl1+P2Mtm
b1vRXG4du71P3bRYcbqftR+ehKLIBld16lNg0Q4UCiwnvJW7F6sTvEIX8Fge9Zo5
mSaeAlvMwoP96RHxt43E/il0bh7U333BkyeqDDHrkTgVgXQPNr5x/+vYQlsZjy6p
REaZDy0aaI8/U8AjG4VEavWY6W6yNq4QZJoUj+c+P8oCx6bkabwPiSZgOq8JxKWd
wJUE9NI6MDFgHdjX0byPWryXbD9kMbIjkUMic8Xs+aTX21DTE4Jr8Uaailf7oAdi
zhG6UCZdOcxYYCTD4dX3Bop0VPdUChptafu553apjDDGQZO+c0T/nNfcDHmVRxnz
pzHdNhOrqxAILDAQUHhUv6ShGzle44BjAomRz9a6NfLla5QBsIOOkZmStjaOibzh
nhdREBZRrpOexKT/3m3E5WWPt6WTIM0EQKy62doKS/Wrn24eHEyrPRWPAd+PXIlm
EalL0RDzFo1juQ0+x7veRfXkMMAKC/AM++czn5jwD2xQjQY5S0o4hwXKtC1lrZ5b
n0chGS7wHhUZGdjDVa5P+IFFx9xWnGCF8HcXtnqZsyMuCcn3oj2riyDSQZDlkrp7
`protect END_PROTECTED
