`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Dbeao7/Pwje14h2kh6WEh0zoIxoIMobZon6s6F+zAMFOQ4Q+xFeVQmAVdzdCyf4s
MR9wXuheqgKJ0yqeJrXWkoDC8gu4t3Ap+toAxxiL3QGKv3kNC3GJ1UtQhZkxDIaL
2WlZQNoBkejIL+7UF0wMJgoM/nc+ZQMR3fBweoMKOUrtio0W5GmPWpBzTKQzBnAu
tbwlevS2fahFsZCkbitjZgBm+13mVPHvVVF4q6GGd1Oe6Pem4vDuBiJ7k0TjCudF
U7IpUuMiJp/Uzw9qNM3OEd+tUgX7VuVxEY+XYCcERHWJSgQr+XB2vY/eCtHWGphW
SWWkzX7kcSMN17ZERJ1GNgiKmjTyUjwEa9EJsMYDzyf9bePbhd6gDh0wVEphpbhw
BnY7Drqm+WaqlyHLfq7cN0UivxW4NPfO8xa4DK4k/jFZQin8xoxCB0hK0hWqfUK9
`protect END_PROTECTED
