`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1ISoLep4Oh/gria978/56xD1/fzScnvvBKA+tPasYh69e4zeS9DFxgVoijp80Hcv
qe1WjNQXugRuOzaP8LYymzAkv31j0QRBNnUNASRYB9XBBAxNlepzfI6hPWR1UejA
0ckQZFuurAs6QwDb0MdmihfMWtvksnJAPXPquZ+PIkPoGhrjVOLhWdBI5XfdJ922
j2E55aLId4yIrAeK6XQhd2P0Z0HQN/CfW4Ii9JEXJ2AnSgk14hxGpCjyK+G/ltun
4HNPXtjMFLma5l0haOrQuSln+nAsVD9HE/UmrthLHRvUzeTuQWnhqTbRyvm2I1U0
Gqz9wERZdYN35vjl5drEvEC0SjohiiNMcKMsaJiZiIgZv7hUl+BpR0q/jHKTmzGE
NH1FISiKiAE0mw5554oMrp3/IoYuookPaWEqRzdayuTLS76jK/6mZ+YSB9AAlWdJ
7m8eXvGhH+rtIjXPhOVfaiCgOYDnUK6JszIB7kbzVt5dTY7aqsMdUW9C+crrBeVO
Y2FnOgk44ELeWCF1rhRLS69Yq+rfQjbx6w5YAADgDKkMwQkeP9g6cRR43tcj2ihO
JbMRxIBiBmcdc5wOfHK8ogfZ3RJAS5idBS82c6mZ2i0ZKVj+muaZnJFKKEPqdjqM
l8GqizghvN7Tuo4rVJ10bAKvvIo/tsVMF1HUuU7Y6WekI0zD9/iXC3OYBusNtnR4
AvZSVKbcJFKH/8J2kwxH7DcdqTodAAv/7QFi5QorrTmVdxRd2mEEtkU4nu42amMI
P8bsnTCKS4itQibL/cMocLSCoqft1e/knLl9KXkznwBOOTEAQ7E4ju6mmgN6QGLx
ld8OJyAUoCeLRecICuwmaDIloix/nIOaIjdAWtKaRf9WwvQLKRCN3iQitK6Hr2ej
CJCVjbXpwlGzaPDu1cAeFBI2Dxb0/bvfZmgxrgsiK2D8RyGLT6/eR87pjKlFpTnf
1gh4oJeMe0YSWGJzjS2Xdg4zcw1N1DMH8Sk5GfKwNSvx8NK6rNpDOPoGAS5pR732
qr/HeX8H4JjI0B6qOyI5GOf9KQpc2WaGOlKV8iUCVdAmW7OZ5QTbgezJ1MMGEusW
g2Im8TOvQx+dOCcy4Pqd0R46tkhwEA/3YdKkaH7T3rhw4jIKBLiV4G4ooJiTejDF
rnhrC8w+D/moybqo0zLWHwkNuLlYrkvixZ6+/74IyYs9ct46AQ4ePsZJNGD1E5rB
mQjU2GVR3QQEVvSI/QiussX/MyEmW9NMG9qVzfTvcrJ6OhVp6jbLbA1vwGd6EyL1
FsHfe6KCYMMSz3BQ2Gb1UMjDT1pBvZc5i6FG9gTTuq5HbSlCBMYpcQIPxVvRmnPD
EpPiCAlCMsv/lVvZFxKMQ0aBZmoYDIH1LZqGlhmvrxlDzLSgMYJWJGRgapMufjIL
nOt1KPHzUzTRbpNW5/PEcJoR3Ao6fAdgyzHJTUOJWNCI7JnRKVSeetEKI8cHu2z2
grmkOZXVLZO3pcFKk8ifrhKYNoeXWldQp3oSj9Lp+9VdYerdW5CnudU/FTCNbwXd
1v37hRZsHJ0f0rRGFyZMhtHOQFN8AvXmck1MmDB0+K+Sa+kyzXjkg41kL5Q7oX5X
LbxXJjs9LcosCODzPu1zLCSmeF3BYw4ToETHmV1dywPGTLpqgNTEnfWn943AqoLY
hGaCDN6wl/udscSriK4vgiR01x/Exw9kfCOCozsWmjnu7Dj77ANN3cLW2arYKbSo
Aw3vJfIn8qk3M1v8a1jNRDftWWNOBtcFCFVylYWHMRFTnQ5keWYsbltGMTUPV/OX
sYBZ3A7XDj0C4xP3LicOt7XPM9rbJ0UjuGEue1uAlE8/JkGnml929yiRXEgzZjoX
07TBSVu2AM2HMNFaVCMt1ner4iVodC203jWI5RrGb3BhETm0DR1xBHo43COxVj0S
0RDrDUD20BezW2JDaKtJTQ8g2BXs4gx1sopqo7rBDr6v2N61AtcdGou4yDD6wVlF
OAP93IZLxJpTtPmu48R9+CzfjZx2L3pmXq0dEyKH9P2PucFWcdfZGrrwMGwTq0s5
zqrZaOJTY2uJ4Cm3P5/EpF039WCoMSt9zeN4ocn67m5m0vehCxRgxHn6rEgZ5UUM
3dELZWmBFkuqo5hCUG3rzoHUBavOh4ZPRZPkHkRePnp/pB5Gt23IRTPvXxd2hZaH
tfjMTNIgSKSET2XkUboHO3aCiCxWNIf1tJV2T4Qh2Tz6NxK8epJ2YNTAOxT3bu4V
yMsoWB9pB3uPhTEqgP7b3AvnQb9JGRrqXHMMG53YvsKzuO46GztZIEFrh4i3RDbi
csBvbDz+06PcQxIWKwoW4p2wkHARPKn0Vq1hWlBx4KXra86VOnxN3prnHwcGJ8uc
2dfBo+8cKxIICiQgYCjKGoZl3wXsaDvKngWWTz3Ms9dDjDq76WSnzGDTH+cH5z7g
s+IPmk37zdDeZ/qQsfuZNxuby0A35FYk/bOvzht6Sy9lJDyU3jAAAlzlM3qNR7jF
ylswj76AQ6z4Mgl6um0QPOEWadOxWy1pNPcy88RptcbksU/YEA1qdbdh+IHKpGZZ
yFQd9tb3jFwF9X4iLrGSWpkgISYBkCEVI4wyEvqXkJi/1nfTFXUrBv8BthyuDlb3
U7o1XcJO3jIpBmMswCrKRjgtwmqQ4fdVi13OIu8ijer3IJoyIIa1p/AJqCjb+TJ6
qS+m9qguCJgPqIwAWuMpoxl74gj3QpYLoJWn+0GbINGzBSQPCSJqLFwOjIyvRjyS
gah63O4ZVJjnme2SGq4zt5lFUCZGHWljaoNNk4tMkxpLtlZfyyOp/jgWo26e6kkN
20C/dvwPJTpdyKNgDUtUbJImJqve9LJyfDfrNtdYUiQxtVcm/aYvhvi03pRJ9wFc
wXfBkFt3ZZUrLwBEt1S4cwIVchO7XqVL9FlYzFPJRScnFHq2zitSp4AThc/rJOAs
QIicGGTpQTzLhck69ljk5QT7HIfuwZRM83fikDIirbVyMMR/Ha2590+fu067gaCy
03BLduk+i2wF0uemxYaGz5f2gtBomlJjvUjbG6XQWISfeUCZBDYLMRvRmTRJJ4ZA
SeP6CQIsju33ml6wXoAGEbMuQ598MzIFn/PL6OkTx9MrQfZ1YgAQU9B8Tw3UPjLl
i6agQTC52ZF6q6fN0b7Z+Z/IT8lmGUY4+1a0bQwPJrNwUKlEoYBuJqhrGKysZNSp
X5XYeaIHh/e8DBJDeXRQ6E7I0ogN6BZyLPy8U9AyJCxnU7eFBceXhBT0BW2krwN+
EdtcCkvtjED+8NTHg24J3iS7qGFCgoS80Z4Tl2G2bwSmdEAWbZI9T2e20M0BKYsC
kgkRl10/OnrTey51Dz62+PKzvLZnUyaDUZ8L6D8v9cjPi/Qe4IK21IbjKO1B420A
Ubw6iQM6PxzML0TovHsunu4Y7E0ByF9wNcOW/1BsWp7H/6sVJZhSO0Ga3lPQ55cf
yIA2e+VLmwVzz3r34s8TCTlCzyGspCRKO2EBMerj++HBEYtvqfjeJObnilw41m/5
l0pSsCbflht8S7K+t1JET87f9qZSyUfemLre6CNFIcswwMDQV8w2kMPRu+lIdgRP
Sbo2ZIf4bhU4KhwldW8/EccTMTWE3sPvOAMGrDOETqLafcVfJ5nS4QKvPeemGcn4
hYjd+NwpWB2svhr+BsFMBKzJKMAJTMwfyPaqgvZIpAL6nKFVjIa8C7HzW6RIghmw
+apW0Giq/8oJdWsROIxL1hrxHXbbakM7lrkuNmJ44SX0QBXqtT1pj88jfV/spKBq
dXB402mjKnjQAuGrFvwSPVaiXb10foR5OnXnQKOIWzqtNM9/xNkLbaZ90mtZtNvk
HUWHE8crUWGIs6wc/84gtObNgkbiTj/lqlZ9Vbc+yskefDPkZbFDBE24FwY+1xC0
ROZKcAoFgmzd3XNe2A6e9mK01qFXhA9PVutDNaYdHRO7LOxcuPyYnM3b4CRKapOz
GSqsIXkdKZSev8KfP11m9f0J+RDWtrwJjPy1hdHs8rF1scK5uoE/Txr30IZYRp4+
eeTnpTGDFm13xZ6e3brja8unsZeo2C8habCKIlrIIHToUQu0bEaHYiUrBRsV1rz0
unH5J5bKUP38/2YqWwxhpCKHcitHtkKtfoLQWAhHV73zcCn+B463akyWHDFGQCXS
uo5yuazcRW5Pcmobl3S/eiYMncUEs5OH0VHM9ENxh2YicWQfPOyANzLHCi/czdef
qov96+/x0xNk63V5KNOjBfXhl3jo8ZX7PbK4YBsMPt+Rupj7h2a/uUMn62EiImjp
QKXRIjhOgejfEcr2Iv99L8l+8C4LfKvp3DXbOXfvAqVYoxZC5ffDqk/kfijSWAK0
4KnRUNg7jX8/1fXVmrEEN8EoDdqAlsYQka/5rw0e8cPZIS1o44HbX6oxtGykCdYb
vO3udKfKb8KXzo61KdmqMPvD3WMXeGeDXMA6pFpN8rSoSGM2zvX9ApR0X3PEKeXS
dzWWD5y+ctzVAgsgWRcdWQZfCbSTxbq6wdLm67s1oZQIQ8HINUx++G5YZHnIcj9x
DxgA7JQqaU/JJp98Eue3Ms/ue8hSNDB0UHDFZPs6uuehpVnO1LY0UKVxyE9HC5vI
5pGepR0/HB4R4RzOPM6+qMEVi68Y0O26Y3dX66iu310xerLtvr8MVuxFe+WNArMN
whsoU8x2ROAFPuSXoCHk1W7jM1LkvTDj1IyXgd+xvRUzWWTRglDLI4h0K3MqYhxe
6HfhZa5icW2ok/VdBX5FA/4hao/yRgO9S4skYYpBzzPIuYy5h+xjQn7xQoOY1np6
EZrxG/XnE4QnXIXJWPSMm2OwEpZWO7o06Vje4vbrYrr4CUtWUpfz2bMqDg629H4a
8mA/1iv8dNZ0ygWNELUa7uREvi90+vDGvXhRF94TSEFw/yTHhksbaySienEtD376
IFQr/qc6HyeB2QLkyZ+YI1FiayTLajSezwkin4FS1qnVKHoBYHxuOLtjbBD3h3z5
R2aA6Nd4CXgNSKCUug0cUqxL9bie7wz/ET4cPE0llS/SPjHupbgjVxqFWWlvHFSp
M+h79Hjmt0ZOo70VWMifjDVvlm2Vn4qbGGX+CedDq12Mk9UuVMFhNRIAn/fto/XA
XAyi1NVI16PXeSAmtr386lLHAxs64kO367wKIyo6zPP5ICSakLsQ+fPFil/dDwZc
xxVC3B/7MSq8ZbDszxPUEn1C9x49w8XpmoT/au/OAUIjwzt5Q2zxD3wE/8ykkHGQ
jePs4UkblYwU5Dw8lGzp0qci53F3Lkg14Lsjc/uLpFrSHJOuJEo4S5i6QHZo3lOi
YZ5vaocliGUCscmPKyq/IuYvj154Wj2F+yLI6TFZVKJbVp/cYeJ/+fecC/WQvi/g
yQ0kjzAdf11hdr66QxLm5IEs49yKYnHotSdfcugAiofS4KiBlXoasrRhUXLRQkuV
+lw4v27omnENvPbbpfUoKWkFmV5SLasHr0fNTvT1HKOBf/fZZ/x7fgK6yxnTpbfY
goNvgBPHqkQklV78GZ488AtY1b/rX98jrKiUCBasWX82A9FUsrsVb5Rkg3MCBZSM
rHIbJhud142Cl0ur6nZZZgSMKaHUbQUXChnaPZ/itcuFER+cHmmu4hDht5FYxmud
Sfd8kn7Xok637zygZQNcb1S3M5w7YRXkHr9/HSHxEXTu2YfOvLrJCIG+Xenz5BoC
xtaOhZPdCQBJT8SogtqRJvazQbsegeD0dWlQmnIIXKnFgT4ceVhDJ/zLblp3SCY6
mJA55bmE8TlZ3Jdb3A0LEacLD1tKvIkuf/i4jT7xeFYFMPMZFKJBVRpdG9B18FwK
XODVortGEJka1Xg4P8o/Zzc5uwg8GBdajXPQmmynjdodRLe4n8pa1O4TD2XjLgO8
eIWg1LdMkjfgfzPYhvlNCQITov7/EmhH6SGfni/XgKcC8+IAt1opAl3HD3AMDjbj
gFTke8hGBaqLZSNrSfKIRMpggLHFA/BuUDZ463uXo9hMMQpgT15KlZlEb67A1v9n
P80b+3RhT67Mj9kqOQRaWBd1u06z0XILvSbD5omFJ0FUYoGTLD3WD/zBtQVDdS2H
UqWGc9Dd9wd2e7duIybVBXkpG+Lz5tp4x8/fx5wMUu19SSCxWX2ELdTY3GGuBQ8k
nICm7kClpHfNy8iJaZqpRJlKpAWQOlIPsf7HnbqrA41U2qun+LVHI1eEAPzCz63R
a01mmYGgY55IvqzM5ZYMl+T7zki9xgSGTIU8XDMKU3AD+nvWGOFSEIGBks4/4ec0
FGH+l+mz1q3oYJvzAwdhbpTNXp7Yed3zDtpbdTLRCwYa6Pk3dPdaZ2s6FKZVI0iE
nZM1QoAETH1V4PpkQqvPU6wIT7BY9WUSNcUanGKDCtItmQNULqvQUoIpp2mNwjmf
QjTqwa32LYlxPj4WiV+r8IoQqKDh3L6ywMBHrH7+JYGjwf3AOaboGCry8PTuznMb
8UWc5mqQvgvBVq+zLflAYYHY2icSbMBaRocxngYp2e6KsK0SXeeE1tds5wf00xAz
fBejQz0KwNV6oCivweTH6bSFYlpkbq7/Yo8looLy6laqYRCWduhxB6QPMkPtpoNz
28t+1lGlv8dNpOPXgsu6LIuBIv0eAQW0OMSTiipGkOrMLkfk+tlhPNtN+o0ZTk7p
pVXnifFg/MOBG9aVyHrnaQypSnyg9aPJQ2w7+pJp52MqWCzlRz1HryWOqNs/8Pos
kq4l4mFKD4+4CVPQNX4OHRxgp2+kc/XDmn9dJToXmySuw0RZjRzJPsJ37SxXHtjR
31ZdR8/NMx/+30JjBborxT1TlABiQKMZG253vm8FB0+P7IDTgkkTwQgam+p79Inx
au6kiMYddk8yBTt3kHhRWvahOqq9KY1hlPPhVxT1+EBBsTehVLoibz3qK/GaVOUn
lGYRO2HQqtQe2NWEqNode8nf7nJgsQrxTWmFdRPdexQmM2pcEnQGHEzxq7vGIFLO
orOG6kHFM+KVZF54DgWN9b77sNsW+up6UG81h+uunadSCueLLyMNhM5C+XfRBnI8
XY6PJtIsereyzuLQwcbp83mXOHqRMW/AhIb5xi9r4K39+V4xAuwJRk6JDxJCIzOU
tFyHcfJ8QSFTnzKPHuKZ13/Acw9z5msEKwVm7G6fsxH5KX23Awzk77/FBPi7uX6J
UZF1u7+7FgfstKtJlRdx2eYYsMYraHVeYhsGF7SMZVXaiRydUmGbRmNqfrVHd5NX
7leGGbJgVxXCALxY8GpccP1M2fMTjr/utXMabKEGHJJAos8wsgWYxnj0gyOYHUS8
4E7dgjexp2PHLdyPxqsMZSLls5Bs/N/E5SmoNZOao37qikwY8mljISfTBHt1/wvK
wA73KqqKpWkxeG5jx2E0eTB4fMEgRdymCtQLNhAug6vTOT/jXXlWWd7kYoBAbIMR
TvErWdipo1UAThAIlb0J67dwinsKFG5saQTc06vLyRWOgbHHcvL1A4poa1dLfD+Y
xUs39vNU9Dd3s8+rxTp0OAvuDgM3c46Q6KaYOQL578cTG0ZSx3WQAL3hHjsgPB4z
ofz+3vcycNFWyIM324FAMdzFNRhSjSu3XoWBSgmLzu4joUWyNlwkMfdvp/HUv0tZ
5/4qrCpphWjofkG9hnRAvIQ6NXUtTy0hQ0kVQx7D0kpOUuiuZYcfilG1fVLfeopn
ZFUOpdy4ZLdV7xePLsbDVl7RNafmYNfpOsgJWuy98M2v9+LMLmcqfKQSDZ6capeF
A9HF/CZnzmhEEg3AoFuc4rOUzF/8NYOlkjXoVv+yGVKGUgiYzJt0SHO78Kfc1MBt
PvNKWi5xZMB/ksgDbwrim4m/bA9VSUhih8XDBMatWfWoTQKqxTkMPk7v4pfoEzVy
P+skV199L39IGS9Cx5U4PciO0yR4LsS2XVCbobLeyo4cKOJ3RkGIvMWCYMo1n/XC
owuRkE+yuY9Z0zwc2apRN1nXNKmdClImTJXKtqR0xMswhTLCCgvLNsRXDLYRL6Xl
Cz7Ge3TvUlmFAt+zzG3ojMLmZKeVQ2sKo8WwugZvTuegz1kOYSsn/fNdNkD3VW8o
bjJpsRhQsEzYwO2b2Z6Dy9VznqjFSIgHXuLW4R4YgiXj3IF2ujIf48ODjEqvNkrd
kB2KMcUTvvxLyTt0dbhxJ3QR7SvKCmRUmkpKbOM65g0A5CehaknC8vlHHy9P0JNs
QszW8a6t66PIeQ5dh0pY9BWYVJcmm3n4auXCHyTSRt9f43gNPEVX3rHe7OABpJCO
w7sS4exlPyF4hL96ugAbiNo8KaARpPXOtksr7OJKFfk+yu9apfUYebwudb/WFQxR
rTwCAGSZHA9Gh9Z35sLtF4ModV3gyRGuGmuLJUxgVRPeoXeq3wl/i8KGWcwGwNnQ
fLv1JqUz7aSExeYgdY98z31ucOb35aFZqQ2RNc/h9HoovL7hLNogs5x6Tqz9eoLq
wmP7MJYCycgaqA+L3iojvrZcOLLSuXw1o3K4UOBYkWnVwzzvZA7P4xQW9wk4cDwI
cYpbdkgn6zirG6kyySe37YM/QoZ4kyqu1QOwmLacimchGhUtLsET/hEvyTMpYmm4
8HcNuvoysTYxLfTo7y2NGNTNFUrXNHkKmOe4LSdsTOb9xhmW3unBTcL7j00g8n9O
B6Bw7olcKKscmo3PPUa8d/KxInmSLfWd9rWsHTgzAlpa2DyLMMloGIVmIsMkzR9H
s9v7yrs3+3VPuF4A1+lOdiKGxOAX6Z0/OA7LqXnpANJ/tzjXlJKDThaMG4mkb6vq
EqNlPTh8DeefxTSxvsNKtLTHmDhyANVgBf21sokU4R3TVcoGJ3QzVG4imSpyxPfG
6AJJ5MoGz9qIlM7cYrfCgDo9Euk3UcpI1j8pkiKuvB5XS4cPgP6xqeZNoB20BGtu
LoIAph7k8zZcCdy9Y76puiqSc9TDdKwQUWFB3DgTSJhqGhFdp1XPftAh0o1Iq5TA
WxamLrFwgblXpV9VXTLsHMO+kS+8j8dn6vGlUPr7WbYcvD74P0MNO7Citl12TQEW
+jp7NKXjqyBSxYb28/+38HdLGB6YMi6rT6RneLyuhew2Irx2Ggupml5e3I6VNQ+z
oJFhq/RvuetzG84U7euCQuv1k5JicASjaa8kywkga1EtIlygKSkZSmJjc6CY/+pE
omvXjK/+INXpb9HWUO4tL3dt/yY5SwBhCzsHkOBugLOLfSlOxp3JhIDalbxd6VkC
A3LoDUM3n6gvP4Dy7CAp3juudx9xZz9urEi4JaiUovhdHrBm9+o6D6nCsUe+Khll
S+0LVC58gFrleLYUNzig6v2lQI/RKwsseDEBGVi099DsD1w/bb6ljRmNT12IQSBv
sJr27T7TC76lLbs5XyuDbRUKcI055kLU85ORHBmn74EHOnkX7cVWccRgVuoviMCg
gPU7Fp1YvpkiBpCTHGLxbZgGjanhzOMVEDNjF116V27MlIDx3BXd22oUYgcu5LwD
OTyGjQGO7SnfdoBd31pqLSE9/WxDZr8VACCtngdDzqpZ4jJPRCO6N/Q09AtSXbyY
npqsMCmQeSQOOlnpxjr/w6RarMRKuuWUpAB0iKizMAL88+oE/BT+OxjZiBy+Qf8a
WyHk3AKGTQPDCgE3HJ//qdccpZa8rZXVE1H5EwmtjshO1DZX34M8EEy6wcDUwjeY
+bPeZ1TEdZVj4YjlfnD6hDD9Ce8zGCHbeIHDzfZ7WVSW2C8GgrBtqco90P7hlUOD
LZ0WtdRTi9kwmI2LSUJTPS0+fBhyFn64KbOBg1JEkeoJJu6bC8BLq25WOBNIGvFN
Bz0Kz3yR5+8r+vmub5cw7TcMd2KlaS5nzoKOhojDTq0vOUEjp1a5ncMbzIL5V4C3
KcRPPQsJco3zOgqr9eOLkOO7T3k0vNST6WaHIi8Xi8F+GdtR9L8eNR2XB7ZG9IRJ
+vYyMxRpg9ZoK2iIrVksZPFuOol4ZvDlQSPqpyKfZg3Htu5Rt8C3QD02p/WwyNJH
dgyVf7rk8pwqkeKInCHGnH2HfxO831RnOeo3nb6OPIt8i7l/YnERCNUnIRZgwsX0
2vDAKmvAc0qYs4YZlCLfBmJBGY53cDmTRbo03gSnuVk/JIE0q/2NmaPgWJw1fM+i
gRzdV3FLQJ+ZVZaOn/qBOcY5ALK47aLOkZFElhk+puQ=
`protect END_PROTECTED
