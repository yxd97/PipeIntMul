`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uGxQVof4j+EiDLM5HucOD1CYNXxb4zxu0W2HMxm2O/DJ4kyLu2vBSIOSvSO3n8bJ
bsg3CwY2cf4MOeHBtYycG5m2qctWC16zcCXEnMG3KCHbji6Q2qgxxrt90CweFbnS
Lx7xCVYS7hgHrRLm7maHlQN2/Sm8EKoxgGLBYwD15tU3r9vfLecn6SN0FyGZOF9H
IIM6QATistM9aG0ovrPzIbv7JzXpd1YbrCQ0TA6U235X4i/D0ycaCK/Q1dhwciDh
JXZBsCYv3HLsu/W3esTbQXLFM+wWVEBbg8k9XPlv83j2dPzuNuAEOk9/wq0Uy2SG
nzE+EjGa63dFgSsj+rivtGl44WMORvYkRLA4gppdoT2SD12tbm+HGiJRvby8UFgp
MiHZSSrnXv8hjli5K4UeTQ3IgKwpi9g8PNUOeP4WAY8sae7avFN3kZSMuLqdvCEx
AWblQGkkXr9P3JSquU8oOlviCHexGc6klLpmmdODmVouRoybmSJHq2pdMmDVSnYq
8XKFOv8qalv6H8CzoMLUV9hEraQLrDUj7/RHtmJwYHjF99UU1Rm7rLKkuIEgtwxH
rrhvIgti2oqvs3fpnjAJDdFA1P4raGS/tWXs6diHxM/kvvbvwA6KyfoRRHoGfhqp
ByA0Sbnpdtbh8ZbbaqN4uQSsBUM54MzkMAVPCv2LNL2y0MTmL/VoMMXWsxsDw66z
/CctI6AaSi1M7OIRt5BOYk6vq/vmJJq2V8aNjlu41N6OQYTPXC/ZctMWWOs7ds+1
jCf5Du/pUk6gTFpeOC95fXI+/F/rItAF58PuaWhJXcgED7wbbutL8hqB6UiN17lJ
0j8fR8aY90zvHptXyv+ELVzQ7RYuMKGxW/49Ldv6BswwpsPuMLUrqLPas39XNOgp
zVbPFHhlmy0CMuMty+P2cqMPqyLzT9oQaM5LzGs2IOhIZFvqAVcIckcU8bI8w5fi
+maBwntTev8iFw2ecVnZi6jfZtSbONNJSWAIpzcCfWFqAHDsxwcb8mCROrOfLWJG
Hzvs3Bud7WHfwjnCFl1TdwyZTZR2L5RIywKuAy+0KdZ5fk8rEWIbU1uGGR+6fk3s
/2pN29x3lknR99o0zqLNfSE8QF8MXyzEMkA4evPmql4OOzpw90JF0R4gpZstL+TA
A90ESU0buTQHIGPV6FlpvxzAo8bfSQF25gRJGVyUaEit4dwbZsXheyyiqWYHe/eu
L0VEIPXZAkMmofFdZPHouWEOOT8tLblZIr1H5nrBym76hnCkkA8dv6LAyB1YGq6v
1KLHG1j+QavxkGlfPXHBT1C1WLBD0upFbkghvxCMGqvrgQStcuDHQyshedo+BkAk
c9UIHDGYQuPC2ARGlPANKYxcQpaNmu7dpHFkQDVlHZ1Cr+GmIRTo4Ob34jt7Eyuq
TlMc2N3+h5fvyVw/ekEZ1e4UIkLuQFr3ZQrDaN21xa5nrFRjhyHYPtgPKMy03CPO
bGIMsaEjAYRM8mrey7mfU5/vdVrr9BAXbKNkO6wyCXnUCupz/vxwHB8uRUncfI8p
ZFV2gg7gaUYKfRK3UtbcWDG356ATP0+qjDaC5BnsR91Pk1TqxJcQcYJwbE1fafnJ
tQJ9+aCaq86+OUf3CdW4y2esn+HTo+6SppqUhudaO6nGqQ0YRU2Esq4n6q5f236B
mx5Fn1wwyzhTqU8PTLEYLsc/GjQxwbpIhJOJ6t6GSq6vaaepsUckSKJIbic9W7Np
6g3Zs61COmmAx1ML6+bGF8AC+y8QqcBqysUknhsNFDCjASSN7KUU6AbbF4c6JMy2
T+mmhJf6wQeYJ3oDFdKmwqQ8jS2JIs+1wZOh9X9e/dIfyQZ4YbqTSJDXhECBRUJB
+rhIyOUXNUWpjolKGBDKGcZ60AzCa6CgtX8xacTHG1pFoCdob6BWmUIWWzf4TqPu
YQKFnLzBnJ1m9exzMpF4gJpOZ6i2yNMq7tRc5H+oS/ApstxO14Ylh9GwzGExY7vf
d5ZtQQ178N/RmmHCjRUbptfZZ9rlxnTLJKWvQ4JsjpU2rhIVORx7f1I6PDR9cwDm
aBol8jNF1uPGQKoEHX4totkMqIjkOOek1z5yTRyOPe63dE1RDHzuDd67SepYAL7W
AsY3dwmnMMpyN0LgYNLLvN3di66x9EW6ovbA7cfKbrK1XXRw8IktRfwARGmiFB1p
qUInxs4NKTx/0DtGkw1CuKkR99PCNhQ2QG5fQDg6dplwcu56N+o3G4zIHVSmKpc3
H1pc1DoQQkYb9hvORDoPtmqyNnHS6j194biHlse+uQwrAh6XgEO5efBJnAnpgoIL
S6GkKZk7Z3EU3v5D1NPOkD++bh7t6NcwJOzYvak8sVknuLx2JMqHyQh9vtSKv3oA
E6TOX5l09rohfHgqJWWAg6zCYyhMjsH727KCGJGiQySxYdwwGl2B30Xe4+pZHRyV
gNQSxpz344BK5QBWSSPcnHBDZlOmlslyUlY37YjqIgds0o1g6vcxsLV+1pcrStS5
4pJYJY138Z2nbwnWZBuKYWcssYgndy3yezOQnrvqT1b8oXidkDYv7OlTkn9VADzC
6VluaUy7E/L6jZlzjL+BfmdI/K/flW39E30oFBUXzIlhRVDAlSXkrs9mg9NIgtji
2FLbtdNABiqr6Kk5TOjgSfojjL2ATLKla/Rmv3mLuUNKpYvL+4Kx8S9W4DfQzOSK
tnN0OtJHMdg1dm7cG1OJHUppWr1iXbgxYcbh/0KIa+0/NfEqPigOw/3wA8o5yami
0D6oH+lSf7aVsm4K5ilhEK5jr+OlI6PDJ4e9JsLvJoOAIN0KF2tbXpoQfk/jThbp
BYlnn/UOJIkstnAQ3cITm7Ap4dazNHdXvnR4ABhIsZcI3doZ9PNd/KHW+n/9lSm7
FmSngqldnh7QeUTqmBsdaAgZVfC477HEVHW5JcH7f8pyYN17veRRnJskqja/85S0
A0wl/AgStttfXdLKbY/fj3+6ou3h9coHYYiynDbzhXg=
`protect END_PROTECTED
