`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7BgWbMe2zoiE5qx8VtH90bYQ4ecv38cBQE30MXSgZlvUbFcZX2OdN4KN8lpqm2KR
UAZrBCwxRz24JOCmr2w1yv59HXuDzmpNLMJq8z5qtjCB97s27wpxS3qSbvmrrmCB
aUR9rCQGfZpkhIXV4rZzL6LmGQtMc6T6xwjdpXdGHdTLeARDcY688qeBuXPIUnc2
R3tqVfxnzrqYeeKe4VyVL/til82ISGdeVr69zdIWBa2VRxTJpVJsUCsLBEJ2V3bh
OiG/CQDyRaehyF8ibjdVVJoi2w4HBwtGsAjT6QzsRyts3NKE98QSHBvLCrHZ0wR0
LmxeQf9LqSYXsrtBvUWMujG/cuKKnxCSEitfUaZf68LoaHkwuVGh9FPLEo62uKTw
MXSNvnz6EdugU/TF7aaXS/a33SSRUDedjGXOpXxOUfwdx8cCo7yj6gnNm1GGzZwe
R3rI+dVyvXyMpFxfWiVAuVijO1AOCpXi8fkZyu6RoWLjFvRuBTznL51t8K6zaQWQ
zZPdOwvcAp7BlwnhWJiKrxLThaKXxxa+EK+5juu4S/7AqyT1pNiq4TPlVpgGzusf
AW8AYgY/TB2e+fbmnSae6P468Ww6hKMiDB4SMwaQDjOnXBEh5u40NtABfLffBITv
lyUDtKXwOt6wv9500oBhyw==
`protect END_PROTECTED
