`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZqVeI4UeEyUQSZ86J0YZGmV1Qc0mFxomw3MC3zuSGrlrxPwe3fddh8qaWiGkUsHt
EPFWU/XH1AZ8B4B1Bdm/tesJLue2l0wQ87RsbwPeVHns1pycehGJY4fEyrn/YDVX
9MekUxvw5hNzE6X7VycyeY7SjJd+LAZj9DdsseJV+tZ4KlU6Ztfw0+Orw3n4BBX2
nPT036/yvPf4GC9xKRjjUUtvzv6e7owD3SmeIYEyybBKWma9n2iG7Qp8vluKWVO6
PKRQTlf0QOi0F1L5dvSzJS7t1BLxDelFQMT4R9i4Do7L4wj2n4I6T+uKUxYgFIzn
x2RBF8njL8SRezmISiKs0YEIJ/mvrCK263gpuJu5i8tcNhJFe36Mv9RdIwbBjxV3
u6a9nbbigkQK+QTsL7hXlbQtaNbGDUwEwv80m8H+Nyaxqb5ht1ckATyg16G9YaGu
QdYHJ+VSCIiydPZh4wgKruv9voZ4y+4G3cvDgYQgzHlFrUCxkFJM4PZeJn9birhf
w2zkQOEjJTRw1eyqH00+gFaaU6NLs3qjcfuEYn5WMTT3fvKBdQtC9qw0d12QXKin
qvn4/chS5rVpc9+FoukHvXrA1EuSXewdqTneVoK5LJC/RbZTy0NcxyUNw9sqOuJe
L4eNzpf6wUQHsXHXJRx+16oM8Ya+OkE4Y9qB3ZshBLWs7mMshg8QKO8asFlh69Ko
C2YXFdZuJqkAT9oP9iWKfpmHhjgPWHizt/AGEJWJEsnxRlLvBo9bAzudZW4HdoNz
0eMX4WZEX7UKS7CY+cnBQW5J3pe5nIlFpYwI/CBje/67V8ZRBMgY67kbczP8JLM8
EvuqahxYFXBOcIgOghuf0uOQ1HGSshJyiUyldigAWgik18z3ri9Yo02GOF+5Fxah
8Hr9tpKISHexwvZ9RmAguLXnMU87Q4I3RFBzprVUjuXmdAhxS5fh+tcumoTwXiGh
c8WU0RQOAi7k+vV9JwzK7w7FK3TlzPMkiFN7kRL4TBWjv0bmmiZLyS73IZgm71Iv
qaGW8DiXSn6UxoD84YLzGVAeUxIuwLZAzGgBnDdkfcJc6pLfCgEblz+W9Doqojbc
+USNvJ4NjyOJuezvuwr6NJzEXxF30vj3gyevDO3PU82XAgXGf1y9xlMVXZzFx5mn
pbHMTj5woT38LANhfV5TFtiUlihoYZKuL9+F84CcBc6MruAacDYE/piqJO4SPLR/
5anG5YWgU+FTV2JAbQZ8Rnse06HgkAMJlUMBtt3BqTUbF7rhUk2s3yzsgngWZNjO
oqFv3Amj9R0SYQsykKsYreOQeVMg6KjSUNtpM/0f46xDkK2Eq9tayZSZnmut3NXe
J7W+jkVoZocwT9ByB4zAquR6jGcNOZTdXrD10lsRxW5Xbr/kC7XpdmSGaX8RUr8n
uhCws8XqehCgQPjEL9B0BjUCrIOrOAT34Fi9Pg7QrEUOom5g7V0IAXD9pAlpeJPo
R4kTbNMK0IDxjuSZQmRsWO56sUdWcAIzt2XJ55kmjBlICLcuE9p2h8+qZuW50y4s
dc/hhjGpU+LPiXm+9zF00GXclI06jk6sY15E22xVqF4Rsc6od2lqw7Vx4W4wsXwG
6U3hLLg9D1bgUZt3QP2VDTjC7uL4U1k+Aeq/1rWU0bn87bzAoJpQ7FQzDYSkm6sx
mX/Ixs4vm9U8JL7Z0KgzlOfZfeO+LrOoMePVN/4v0p7palWgHpseg7Vz9V1Mg5IA
IqX9PzguJ0wJk80HBCcApqu6QirmbornSq/G+rlZec1gVFZWDOOaBRrc6bV6zkI2
RhZ4ifEWxUwGXiG7XSix+M1gfXoTWkSc8kzcoNaEnMLqlZ3GJiF85tsKhbqtdwF2
JjMCHDFx9Z9tNTavrOyvJZXS0/Y0XN1ARq1bghf6jYjq43NO0ZGxXVQBGLss1t+p
p0tjMaaC0pUL4oNYvp7bNsj4v5XqaIDn0Nc0mDi5WFPNM2KUkSV7JYRY0nL07dhw
po6jbimB/ln6VaLeb1WcDxc4WkBRWsmN8/JYcdQ7oAlkhb6y55JSDgeFUwSu/n9S
YrMdGrvxN2PH5ZHoS0zPIcAzVHbqdjwDN4WZNlTblK7sK4+Cf7aZogjUiS/OUAm0
iLnIziZ5On1+OQc5++iobhhwQv6StWt1El4rg+XS+v7yyMH7+f62PtyCvtxs89N3
iXuSt0uflxLpSDYzHNVR3YpZUci/YOi6aLXpc1b4f2gyHU9QfsVmVzUT2jT4+h5q
hRiPbp6d/2ROTiq0Fu4OxOx5Yk0WofPEWcvtzqIKn1AocDDw2tNHI59zmeobD6k1
tLJ44q661g2p5Hsh5RdPl5TpWajoPdKJPL7qH1Qj5J6iNCRCHIolpvGi2hxCtEwZ
yAYhUy6uWjEgwO5L9DlM0XizckfviXN2bR+hZnuZ7Unm4CHjA7zGA8SoAzNx7mHy
fMyvZOMKxfTdUX8PpYQrtHh29O6Z1tdhM0ELt9sPggZnN4KygpRyj6E0WiTDMKv2
UwhoQiaUqUjk48gkT3O8t1ECXNCsLUfbsB/M9aDS2fmQ+oD69tdRQhdhg3Xhj8rg
+EhXkqhKaJcfA7Aqx0brsjxxIzCjdJQ6+CZWI44kQHbvR50J8jlmB2BQQcuE7Vjz
IyqB5SnwKF8ipUPzNy0A0/w1YnIFS58gI/yZhbdKU3R5ZcMuE81IBrrYU4dBz2Ki
BsZcH7FGFHlViC0dnfWlthRD1iFu0juPEizq9OzQrAUYsrtWcPNsV4uvil0KzX7G
KqRAWhOXj2nuU4Va0YfCm+RPbd046eo4pqczzQXZlUH8Q9uxq3sSa5XWQQAMScm7
BCNyBo7Jo2ln36jJl5mv5mvNK98QBY+L0BdjBkcIO5sJBqsgbzHZj3scn/mbgkVM
kO9k4LqUoDsJNY8dt94QR5VLxsya2cZr/bC0kydh4kiH36Nr5lCFAUhEYS3sfI9m
Yu743O6QlURNlpnfC/EWVSwoO+TWhlVrHyQ7cVFi+3uiGFz/p5N+AfKs+gJBE0DT
J5/6+ssFAEIm8aT/pgyFDFwXyuZardUF9WrE5TmKdIlxfZHvCbxDc9LzYrIG8rkO
AmT1u486yrxJrhbxhDWSskROIeLoiX7p22sbAzQCI4CGimRMnKY0H9nqnN09H6TT
9NkH2ftJk2VuAeHh3bsPvXcvt0mLI+558jn76wSJbF9eiQrgjSlkm+KU/MUub1ya
Ef+erj4vijnQCZO2WbHyS4InkXc78Hy8IYR+OHtdFfK15RelXNax2hmh+o8FRnkG
RM7iFRLuPZctsW/QEYhKHz1N6oujfXEyKv9rZP+daRQjJptzzJSeTFOVaTOk+Xji
2o9B9FnPkdwjoKTNiIKCe2jcgHU+6hWBsUbhtad9bdXKY1+Qcmbv5Tg0lpZfL2m/
5aaGdGh4fZRw6IvwhuxUW9WDYZRQyci6TFz0Wga5v/Pjorv9/eeTkFl5K+GY7SkL
E1KbC+RT3nQAi3QpizQwdRZSrD3iEr/zE/wEkqGPFz+yppAzJR67/Q9gLTa4kT8F
gFWyKK9542lywqDj+nIJGXkMWkOwMUSJjsOujelwgfKYAdGyB6xrtadJnPrwB+B9
M7xcttUuEaXW+davodzKEhfZvRvcijkrVT3NNhJEFkHiv62ZCySqvbZyvDE/SBNe
z/ViO4HUdqVryUPutYqSZ188N/7y+9mGi8QUIr8ENXFdodMUkboV7n8Yf+CAsLXn
7oJAMHhg0Onxgl9AMr2v9A030gM8fiHWZPs1oUYt3tPJtuKmlEWaemtNd3cxRnOc
jPd5ttWzhfZcKRfmg89QnTj/iWPSmsBfMwko2qicykK2KqVSHadWxpVadIJ4IUJe
LFAe6MuODAL0VM/6Ir2tN86pQ8/NhkfFpysOiWrabzXw3eUDTPO0aewedqDtCFoX
MT59WiaolTLrvciTx5ZWEYhh+B9FGOEXXWMHmRplMMwpba/THo8+5TrYTdXnFpua
BOD78f8gcgLvJkrXlld/nEMPkdqN/AsBTw7IZnhtQeluhFK8ByPVtnqiAVMVP9zG
ETDPTVAB5j6I1IyH0NZIBYOGNB4vOoHgG6gkkLTbTinbwWuabG15R1jFVAwN5r16
sqUXhD9kThD6bNvJYOtOyR2NqJnlHQeiY9agODfW1ma/nEGqE5ClFnOvPjbdACk9
DLUogwfKOxmT71MwDZlcD9iGD9n2MfNnk2maZDjbgq65vKJ1tq3eBp0WCyFBi8J1
+hOf1ZizWeO1W9R+4HZRSqE9Cf7vmosCWXLfrAZZ2zhIGQfes6gwfsadenhjoj4B
Sg92Z9i111B0nKZszyBexZAikoPiJaZa/1/FYkpFTxwYQLJlT58ewnhFqK3aKQ4Z
Rzq+DLzX2wFBiNXPfz5ZsRcSB9u9fdASDY/GMa+g3jCCc1xIwit3DfWcF553GUaD
CzgD7HGqrWUqv+WmOzlA0LVXkU2/P7v4AS/9pIoINud2pXgWHqQfK2ZOpUAF1PlH
+BKoFc/n0nRU/9+SYDBXhnOhLmZlui7BC2/TVrPxXqkdqR4i0UHiQjBGqeslnNo5
TR+gebZEvV/zIulxYXVTnKPexwzySBHJD9nLUr7ejZFN438+BHp5flzxoq8PFDBQ
5zZOBGoGy2kZmZ+WJjuheA1X8qiyQXpf07y/B1TVHH+TE8CNHLulQHZ8/heG7T0Z
gKgG+LD5A9vlwh0pbo9AgsfAE3NSE3DgItUqVX0Rqj5/+QvA/37AKwE4SLzk9owS
JsZz31SQikk8Hq/fbfjbJWBtLK6VCIUN7ig7mvXLd/e8vZKPsHWoiGhhX4v47jhD
bpnrnw8acqvgqrTz98X/NRDocZZ6D3YVAj/RLlzZDfQdWligi7ObccrRGdSme0JG
tgtct8SHLAck/riiAors8DAJmVQS8Wm39YJ/AKlpstE7Z8O86F3JLqkceqHnnI9E
x1JMAnQgLmuzZg2qyojrzZ8KamMiaavXPiVVqQ1QE7URqk3r/e6QttkxqDsoxfUU
pBO4RR2wzrHecq501pDDZ/QgJw7Ve6IvEk9XzbvJOMc4IMgl3WfsXlBv/JBM5dcW
bIVDkUuFTa7loCBzl1NWriKkP0ay88ZSPNOXaf+Qrvb5PkHejoWaLGQ1OUgUkuXJ
BojIjwhYHk0cplHlr5XksZUR6H9rPAfNmzlkIaHvfJ10Ln8Pz3gM5cG8cKcnTLIp
umgOMsKZ065d5BkCrc7aGfyoPgzDVXWJN6nk2Ssbai3FHm1VNaEcLiWrX/R8YTc+
hshNqCsnDtikb5KkCkyQOJvBDIiVBUyIREp0/4djFx6jsSBKML0WASaRKqxBT5g/
Qo2b8F5MdzxrnzyLFHBARAUZIPx5zi6gXvm7lvzaxcQ5ik+cC9nQR7prmvBvi5Fm
Tu9NEzZVZLn4VsxVpEFbrKSAM5DB7Vw/JoPVl36zmPe5mp0SFqyFevT54vX1M3so
JBCIAdCfBGZvCvJK9zLmW447MhLJm6jbrpZos23SB8SWBtabDNn/xuJe3Lrfo5w2
7YYmaEmqcE6XxJvQdFAowuQByzd3FYzMzGFqs+hdQ4FbQcEx/WhwIq5eC9BuFT8r
ccL+aUh0hI/baKYz1dnb1ywy+WLG10f7kbL1y1xJ6F8PVIhdpYRDMv62pYW2beQi
rV3LLgpWvhctxFFdg05BCPPA6kNlJoc2z5ZdQ60GIHX/Rg5DdcSZN9TDBBo6OUNq
4rnKvAzPikwbXGRkgVwMfIruOZ8nPGIl7SVaImQHlvSW8cJPuTqBFOi/386lmuqf
Atp7AgNgwfYxo+riQjE7q3HoSuSzMCtVEtfJXoKEmQImruGdMQXJ6j3SfkXzmb1+
1j93e4JhkbYipg9hvyAOyJs564UGFaXSFPEoq0+t09BZ1PkclrQdtwbDMwOB9Xw/
qMkyELoKk3uaDAajY0ZeOWNB9JPdYX6RUwREfVT/kkJvs+dvDIPclJXxCZCmU7mv
Bfwe3nm9r5+2cmErTrClVkQ7kkQB7b9QrLbjawN5sWUQpbC6b+QVsxvi974cAA9b
Va9bVWV596k2SEj+cuh4sQksv+iOcbhIUduB9Pw/DlOuP6dJpemo+uhSOTiEXvzt
x49LN63157VEXWetBdTwTniXoPCp5bvoryvPyliH8sICJna3E5ldQvvRYiPtws5W
SGB6EZeBjaYw6WZuEdgnkWRbME13AGyn9r1tw4gkUMju3r08G3xdS49/rztOyS35
PYBT44oP2WxOWXEUVFP7gdSX8jLWWe3y4jMRvvBRosfguJxVnavIXWCyG2OAyddk
qbnZBDQdZ/pb5pTyt//gmPC4ZvkmuqiRQOvW8T/lCGCrOmHpQzX8tmzoHbVa9FWm
2Yy+SgWK7BfGGXydC0OFxeR63pn63E32k7hn7KvKYPyBrPpfw8HUC6hIuEQnvtek
G/+7Cd8TBjuVTm2ChePB8H5zy5WvaM602KB06L62+gbPucCSsbJUX93SefmC1zX9
hDTAB9MbDqm3vpS72Zv1klnZQEoyjrJ9ZbgJo8yIZa+droFtEnUZ5TMynF7DPVeU
n77qfKjtdfE4oK4GQ2l4tjHT8Yr22hlPMsdWFTU64qRxtz7dVG2j0VG9fthj3FCV
21Iosdk7PRcbL+jOxRPs45tKCp3olFjkEpt/mXXkhc51w3PS1dBmCwyENvqaMdz7
X2MpjgBX6skCoUXeZhezJ7Y10o6kthbu0FlGaihCIGTbp3yf60t995yXpVMxPIok
p+yZ4ky2pOhfWYbN+nHLOZp9NOjXEXXkfQ18IfR1nD9dibnZR6HW9gxxnDWPjNal
MOxO0ruNjddXN12n6hfHn9TJyul2Q7TY50tj21//a5MFuejS3MnSJyk58R/c4JpK
7f4Czu9hUaNv1VoTnYp23hHt3aalAnd6IcbpZKifDFOoIXaZybx783mttSsapqBb
imzr6RNb/7+bTO4cgBFs3TI9zrCWh2VICfuO/eDL76xvk7aTUyB7aXlu1DoeaHtb
ctqswmgt4yX+i7tDgg/bL1p4Q6AusKrMmH1dccD0mEHfqtOsPtKZjT4n7ND6CAT7
8nix2Xi2PRiw848v/RZPwjI04QdepEsPFWqnQklkvZW7oDz6momXGMvUTOBqXjku
VsB7RBfbblX9/Z/+9Sbr/5zu+7A8RfBIJanpKZOKazADMZfPDv5ROX0XalBG9Jcx
ahQpVlnSZOucxwvlxSRKyF9onW2r0B5owDHmciOTcCSaqOCi5o5H54Ve/npMgpyt
t/O0ymLO/PmW93MEXUMlr3d9sy1YpAKLlNCAs1nDGG/Mxsrk/1xQo3z9aN34ghVV
JEAJN7zvz5rkxbvNXgK40DKVsfmryK9oz6hI13eVhrXn7N9jJn7+gmhkozFFesMQ
5t4FSWsfEkQapB4aYC5eNtLz9Ryjfk4A5O00NI/TbF2vca5MASXjEBBNCaHWIml9
tmFZrEsUd2709XZkeDW+417J6AwYnIJTw+bD4sTY/rM8ewtR0WxfZrKgtIJOi8p5
y5wl1yNFhhGuT/MQ7A1TgR/ikgfmXuAlrxsIAvlXCU7jRSClAEcu4lyFJtljEVoq
3jvUkBIAO9a+esfAQtYoysltIePkFHxccPd3z6Gpkv1KTaI1SZAirnfuMPiFRM8N
3icNyFcevWuPjx+bPCMNHc5IoDcqkyB3wGSPmQ4k8nBIxxF+QfVmWNKWDzRUxoFb
SP3XYGcQmJ9q6sRE3uX84UGY+O+drAHLH6MrxEhkCXNN5TAQLo2MZowjOKbgD69S
/PLmI4BD4dTjxAAjJBBuEh2MtTb1T4nbDrU+BUyfde1l28Z1B6R3IyJEi+EDMbre
xMv5vwLuIOyHTkC2zOrp26hwOSOUR7lnFF3N/avl86cijM2eIrgQSVe5ea5B7Uxo
asmtL6xhaeZCsURKEIt/+aNdqaIMoOt4nMO03CYTYxYh2mVi+I19JUWx/fiH+2OA
LpZeALAlGljAJXqinA0hTut6PDCGdMvh4rOj7Jy5jQhICXRXucQDqEZp2cE1ePO0
rA7TR+VW5kMdAtuV0CeJ2WH+cqN6VF06cmV/xzXZg1MN7J37cfhTNVCV1VfGqkPv
bmIsLbEjHQsJVmdBIJHKQIICZ0E3/CqA6xjPcgtiEn8mox+IgAi0fqabEn+IwFtD
yf7pW3x7CyuMq7pnllRJFaXRqixn3oeIbsMOfqA9gwtEPW1Sa18XfBBbrwl77YOv
OB+ALCLmwzaSAN5+oO8PiWLhepYn+gb/BmuC32DJkJV6R9AhwvKARvs+L5uQ988W
BCIFHin+CLfeHZOder+phl5AXMhq5rJrRDtq+6q96iDPXxZyM7SRrYW7Zy68XNdt
Y1tkAzrQngs1tu9ACXKgdzuKAu3Pcdm/n0BlA8ToHLO9BJTtBAaFx939pDxxM+YA
CsWJAcz3oXL3QydbHVFG7DvMW6vRCBH1snOSFlqJdu9CeOU2/kcDcOmZRIqvDuWg
L2N5eSB2MQ/9bQkuMRN6KWjghH9uOAUet78vjDhHOe+56qOfVucHXWJMjSjLmVav
CqmDhYPtTzX/Ju9m71RQYKkI6dvuKQEPHEdXpNLMv5g40HPySkKSsDyIBFVg1gWP
1LG2BYvyFG5GQuWHQTCeCxCINWDepswIew7xdpxNbAk5m/J0gd/CMDw1Znp1X6HU
+QtrhjjA3oBGvtmTwlmVkj4uhWKA0jjnzOjZajGIbx9vnHRTVgUALpwzeR7ifD8E
k9/YdF/fvkACMuWTkUtBfamNgHbhIq4mbyj60x+y1XP8FA4778idF2w8OuoESNms
7aYkMdDCkVeW4DDCUS2qKsmKlFCZmR/rvr9kiKTCN73512ojUFEXOvi1x/64g6qu
5FGS05+EEqTEywb48mHb9Fx05vbtP+1ZB6EZCfka0zd0CSekLvQxxeI+cSuc3d43
AEPsn+iUjUGasISAEW6DOqJ7no37UrwKbumDtA4CghzZa8i/cvY2ioPfN4lu5Qa2
Kr+Ihnf24I6XhniUOyEyVKiV+a+iUmIk5rkT3gMHBy0Pq3O8LhlmF0jQoMn5d8OM
oDuaG1xOpkrHSYfCUmdMPF7ADG2AdNBEjwMYIIISjYpGQ3QEiwo1h00FNOSxy31l
JzkoAZMVak1jY7dO3mjtbT8S08IP5KB2nyK2qxmFco/PgMDoceBKWwk4j9YGH8Zn
MpRKGJHIdZGBDyC4DmPtKZbcV7pXEio0V/uu+yksp8IV1pqSjAnGFe++jxY4WfnA
udqSgSe94bDh8orjjOzmOLdIj5cgl1Mq6E5EC3J9S4ylas6tDZhYkpFYW0HXZy3Q
bV8V0ylI4z5bt7kmNfxZqAICtgHDn51iLTkk6HW8e/w=
`protect END_PROTECTED
