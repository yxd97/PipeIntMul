`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iWDsdT6N7v9sWPcT5vV3xSPZS1GRTAF/BRH9GbMYtMzwYVuST1GkKrWloDdOqOzF
fHXGhAoyIzOBTXzsY2virdYudmjyo0ZqxNFlMsin/himcz303SeYu5Txy/1oZ+cV
1yxVBmv5MxYSAaPC7lfNarDzMFDeWccGE5ORuRRTMRsBxaRcm3aFzWgfHerR70I4
M/FyZHpFLuO8ga9hxD4VrEaGiXF19gBlLH7+NzS683+KjdQbM3zV+fbAYchqUryx
Ty+H8di0G9WWsEUN/2uxt/qx7Araas8KcbtrQ+UFbcFDaGpZfpaJnS3V822XZdn0
i8k8kloMcX1TObtOR6ZRmL8w7lKoUMYEa+gftCvMfRJka364zv8to4+nfLMmPg9T
8LguZxvahsGdJ6YpqUb27Kckq8jhrDhOi09YJ/PBhHrGd1dJ3ii04NgBV+kNHqbv
hxWDlYxegTRY3wLnazOrR//I52BNX03E889NWr0JkNmAooFyQpdx9SrqC80mEgTG
vUjX9+HX4C7BSbR9hDbd0qU6jLuOftYrJWJyoaQpMlQVJGo4vMGPGNyMsxk5oZxs
zLncOLq/9O9nPEdQDkRRHmLXpSnw+mXFZ2wZF+N+WlgJ5cY5MxDmn32T28yx4hxM
SPwLUSC0t4ZTbCU+k6F6EIqEcCxb1dA19T8LYboHWxicyLiGPc7aDALq0i/LDi86
bLaGzirvPGaLBPlAw4MVeRW0emrmPZ4kYGjLZaB+kbZRG/PmfPZviRxrjjDTji13
hOyJRjMYYzkDGjU1APU3nHg8OIxlYrlcbGjiprb+iqjzmFQPCTv6sgq393ZbQDXS
9CWouz058uAg3N8gVllooRcbP2PtBuxt1rf14pr1oEU8bryMDvvjnC1vymoPXBah
1EMmEQyWxJthqkUamfZGLE9kEl0cc73tmOyOUrXdhojOnT/8E2ZWF/ocRXqdrWar
dcJhwz8kBS0TSe7/TUUYkkXf1RGjw7sq0LX5GSvYoq+QOMBFu1nf7VsP59G1t734
`protect END_PROTECTED
