`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ys3VIoP3H/UZ/Hvh4uUAcf8l6wGTMYul33hEwR/XbWvPZHmGqRhbCGSlFFTEEwCI
uBaVJf0zseFrmiCrvlviSDDU9csUiYvJ6S0t6gNZcR+gHPCGJwiWvYFqU4rwsCJz
8oDL0CLb1JGBSk5cq2dDjiMyrm/o6+hPT+9mcVfPWt3Uz7+xdSzYbb1G4k9lgiho
ur5ol3XcvLhmz3pwUB5vGnJMup0pzR/WqpiQZQ5As6XORyGLsRjPELGH9NE1Pa8C
Lh2p8Vn8wh2IFvXOEHpXIoN72QvTShv09pYb9JQ5f1mi5c2mXrTqoi+/7NKOJi5/
KQoZ6RG5utRwROO9ayaQGQL7zVbjqlSch9ELFGBmdnfDRqsuRkP8xEyNAAfxmlsL
XD34S52UiciSw8mZvswUfQ==
`protect END_PROTECTED
