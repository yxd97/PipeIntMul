`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ytG2NdmXJTElioVi/9wA69h40PJ8boHQn6XshvpMLh0RT9tKGnAeJd1Zya+1eEvI
ftKJkN+QlPG2KIqgj1eRja6qk4nYkLJ2a0jZi2pCI0dVJze0iZOxfaaeRCPceewk
9RX+Jw9OFiFALrjv1HVbb7PdTIxuvA7dGLXW4OulMUnO1lp1MkPI3uSTWzeK8txi
+ZRBCY7WpbJ4Mig1q+7GB3iF9e9mbWtYMjxArfhurHYS2gFJ6rYFlBNgQ08JaMZr
rw+iGSzCh/dg+yuyiAt8EdMx0XC6FY98w55hvZ/zguLEnDPtMOwHK2/7sXdoycYj
k2Baizzo4q+TAz5So5qJeB6XEWAjdjHSR7qGUb5eEtjsotakGeBj7hYrnM+ujvdN
noEi+9P8k2fTQ3XCRj9kJx2ZOZWWv1SvnyJSl9Ea3AOqQ6QJeSLTgiH0jm9ic7BH
8jtigtRQGEIbWcjpHr0ouXw1WiXqKLSN54JLOk03v9Ah0GKwTL8W7opn179XV60S
81jmeiHn1Q2iOCqiwThq5Q==
`protect END_PROTECTED
