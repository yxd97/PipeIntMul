`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OobTZUqFwGTNG+NtyVs4360SZWm8GmEsAMVo+csGmwTaNDz7k8kAAFn6e2XlAG7/
4y7pTHxzPZ5i/9AZa4f+WWf3fdFOd5SVVb7QD2G2AaqoSBV7YNytN+SduKdm33Oa
eSMliif16XW2j6RDI1jrM3s0DJuL8LrMpnI2Rv7GfG6R3oTuqGcdjqBPqPKZn0cu
hIVSPE1Es8g8CKmGrQ3RkZQLTa2Fw5Jz8ghXY70ZLb92P512wd5sHnvbyADLIfWC
oW/TAYkSrNZw/g1fSgqLLeYgg0uACLLjInHbfW2kjdYbcFt0nECvVUved4H00Gns
3tCU78UKp6LUyd7trEakAAR/4kzESoPySiWtWcu3r6lc8Lbb9vtWv86Q5kEt8TQb
bAis3YI/MxCe0zIzJmN1r2wMyq/ykOJn7JSP4PrpQKTfvFYh/o7Vm8wY919a2fzk
MqajXfLhxxMXr0YMBZZ2ywJhBNeDd0iNhY0XpQo3hm+4Lslc7ox/mwxss/+b26aK
KwJWRLTIXTXhyd5Zg2viPA==
`protect END_PROTECTED
