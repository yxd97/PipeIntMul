`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EUJAaf6HGok+AqjVlrJJCRF+nGhxKeq+B3RPqinx6ajwj5OecjyiwMJc5A1VBlA+
jK2ZAT5noaBI3yiX2kasZCojFn59xzSeNyBEUazZwKaAkMd7B9nEILgE7kcSh7w+
2lWqh5FN/CR3GlpjWWyQXUQ5LNpu1x84eox9OTqtte/eMMpq/6bE2UDS74k+Tmzn
cuVpfqZNjDZkreHYehhwN0TAW5pUI5X9Ta5BPKnd8g531AdSLU22YjW43Z6bL4zY
MDXQ/pDdyhS9Jw5lrAxlbxO6k3q8RkVYkrH7mg3PyMzwiqwPHEwDwbD9FB5/g+03
aBgi1vq0F2+yrsJ6VZSKcDeNJDSH1SlJFWWnIOvwT7Aw96EvW3VwjeHKiPV5eYHz
LBARJzaP4f6nIDlSo+3glNrj1bqOrgCfCK1qxFYbg2qS3E3inw0vl04UcWXKHG6/
Z+fFRmqKLtecNZi1jI9A5A==
`protect END_PROTECTED
