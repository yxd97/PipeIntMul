`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TvKNdp+PhDPEjAE740vrSo4Fu/uyMRtBSLzZZ7koepDoAxO5few/4bZ5oLSnpxaJ
F3p+In8l97/7j+++GKelcwb5c7ox0htoKwaRqSrvHE5Ilk6tB0hXmm9o9612Wn1f
iYaVAn9StCxvQzuty/XHXk2ymVNznqI8mrlbDrx5lkyvUsO/JYKZkmJy0DUQy/XE
x5M9Z/iw+xJfoM2SfTpkZ3Ry55t+YosomYt50TVr/ei1SvysBuFbIcrd8Rdsxj/T
ABc0nXihqgtjwsfhdwg3ip6A+Ijn4cqZNlRButoKBtADTLceaqlWVVL41M+GEorl
/IrSmXrFbj+f145DNpaazSOeVxowfi6Rhpxt7BRERdq1gFXHXcDnk+xIZT1KKC5c
pUoGvXlGbnWOq+jSLq284jZFglKFxGsANwzmZivxRvtnQYrmjPEtX+QBmIauKrSJ
r7+7RjZSBblTMLyCPgOaJlcxDrfOQd47RuSe8Mtyp7olVFRa1BCH8oC9xjG6ANqA
79uwDt6nTnP14xMb6l15bNSpsRjqNdClQy3gjtMq9F0Xna8Q9GI2GUFD/IMTWz3X
hYfo45nydh8XTFSWzIJmJyyNbGIXnvb9kpEE8EQP9QeN5oWn++ODU7SqIMrTtNif
16Na8CyuWYXV0YIScbG1wjOIYvgwivf+UqoHFXvMRUuSbK6dmqYI9ZYGi5scaxqi
3hQoH74GJ6m2ZANs7PFss4bKfIxsTsxZvKpGvBvONMVGzwLV8GyXaLZVdpDU2pXe
H5yLETqQ6uNy2p3Gadrwu1XdcGfcISiq5Wi2ShnDfQ54UAB+8yl0IsccbxdtGb+2
T9gU2z03SIS66mTjoyoUFbIaleZAPDdxl6Ik0U+T9tlegT4MkO/+9jVqxQEGpfnS
SLpofIgC3DIcNSCljdimmvxvmMrWYQ6239zUM0/as0fmbMQzrCozxxOahtd0d7ND
gkpGhzx8xi1ArBUSi/9HBh0zesBt9824S8fQvcmx+LB7abCnwSaMth2klLbOTUpS
VGCxBxbuQ3NmFTtfcjcGZwMEQPU9xpyQ8dNzZo00bFe29hCcsGLyNI+zqk4Ggls3
T1evhWlvHGpOJsR7qQxQ/lt5sS54jrWoXA0HnRXd6gym847v3+2PivfrZZFcI24F
6DNKPGDtDqQx4z/WhFj2XIdZMFxa3wpw09DkjaTyldLEpE2e56WCjq3PKIhjoPIc
alq+TJY0CAbhRObANuEq+9nQxmntGKOLMBLnniCvZB5XMck+r5aPPHWS69Ow1n4O
TFwphaJOIPuzooHNMMXGZJ5smfxxMQMy/ChMB+muxWJgqgPt1CKfLaznyUqvUwas
Yb+kCSaHO0RisRy47aF7bKkW0FyFcLEJtbogMKoHTE+rZU7iz0XhwbNHLt9h1Qsc
ft+UEkhdtsPHmiWOzhnmPJXTkzxcBDA4E1nOfGG4ufdszUNsYdhwvPJ+aRaRjaDb
YoC/u8TgUh+3gluQuUzapA==
`protect END_PROTECTED
