`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
30bSvAcRuzCaG1hXKs43rfUo7xsSw6wDx8olLpAv9+ExwyE/um/CeCzcS2PdhM0m
QaJ3UqbmzY6mfQPxUxeBC1w+7G+MirJMS01YNNrXQ4aUbnFqj1ytrN8qBfFfJc+H
qZc6wsMpvmCiHMgwIyOVZpEu0zPYRdHWpzgOcf9SA1EpepPtKYh1ePnOyFYXdo8P
Ua93ZXBcXqa9wmwUbDcbnVyBn5ULXHY74qFeBHESrYv2XA+IwEkeNOtiCZI014JM
IjikLI44/6ReE/RmGptkUabVoVNgEmHpjcD89JW60ydcmZvrUKaHEgw4jfGenPUU
mStuCTRCxfe0EM65F9RCFr2fEs/x2u2IqKNRd4RZfDUGNys0A7kOrVFAPI+08B9z
6x0OZFlJbirbLKLRS9Vk6dGRcc46rbo0l6BeAx2EQDDpy8tF1EhKAb0qUpprd/Sd
xZAP49kWJc2Rs6tGXSaiVYv3UTwDRG3QJ06rgSrI0CMViFijaS0geWRlF2h43zTa
XECvSKlEtrgVsU80Ti6CBXa9tHUx0Gd1Q0mD+X16leBH1Oxt+6C2yrHm2C5t8l6a
hJYNTEWAJJu3sIhg6RaTCn+STWCrfzeJiCUdKs5rQI9h9nEiFhU6LemDFLgmGKwq
CMWpH77DT/nJm/IoEiBe2B22OED7GRPpmnocYJtCnlaVMguX2X1DxuiZeGXfntN/
g1upvrlsrPyS0QH8+ovtWUgQnrn6qgPB5R+MFbX393JozKxuhk85CT2eo9+WkSDx
eVOXLerpvipu8gEA0p+c3w==
`protect END_PROTECTED
