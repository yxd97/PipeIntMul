`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n8sFsS/xEhfOpGTqzecLNBB7aSTIEubJOngIzlGzpeRhRNnlprCKYznh6MPxrFZ7
bE8YiTYnaw6L1esocAXIaoZlo4wpWVSxLZIncv/t7wE+uu5+hBiOIrT358z6TyF0
+//vod03BgCHu2W+CFSlgAxDt6YT61bZSxUyPfNUuquyBuLGMJqWNULHxR6olI2J
7WxpS+r0FC6YvDcuOqBsCIofx63OUwDIJlTgNv3fniin10JjbCxo+xYg2MSSOA84
Lk7OtgcUkyOqugLxeiUO/C6jrXTIxCkhNFeMjOli3aHiYz9EKU0ANKKmwWGQ3r+8
`protect END_PROTECTED
