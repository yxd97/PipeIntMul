`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WofG7FIlwfaIKy8bwNGkMRtS30GG1w2xNZxqo91ljbPZIcXatB+W8fFvfLek0ekf
hAVk5WvNiynoWO0P+sgRWYafob+dIi0M7ASc6qiVyNdW3TWAFTny2uESLcs7QIDs
54luXh3bEdrCHfkvKTVylnrsFeffa6Ycn4Y32kshusEofrZa4DjImg7vV8OHtI27
MAmwzH79z3c5j6q1uFSbHjYJ9usXsqt/evKpYeuqIs6W1VR/xfpJj3g6AHRw/JqM
HONel72tg7nRSGL2XLn89nTX/D9Gu1uZwA4q3H4YVmu7MfGf4EUqq9SHReX/AL9d
dfkuIV7//ayDim8eUjELEC+oIL3ux22ylCxZqfJqBawcYrVaqHHL0jV3jPocTWHV
umfXacq05I1FqHP2WSszrjMZHWK4A2nk73Gq0HZ1ak8KY/TRZ3mPLvcL94ZwEQ6r
9vAxc9p2ZA0h4qgIBmvkjJxBRwXfFk/8XxzbWiw3MDMx20KPnHrmxCF1K9kkhqU8
8RMX9nzzlvcMuu1yehXCvN++6gWYOS+HCAsKbWLD3Yc6K45yMu35OQLfnF2UbKeh
eSjbK/KEhD8rSQFMqptV8O8TSsNoP0YX2qhbKeli1De57VjrMsxkCTdxqO6tUB9G
oj/ogOWuwaN8QQ3jC99e6+fnbI3JM8wmThgldpjEJ2emMSIU0M45KolFXd36diHv
`protect END_PROTECTED
