`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8cDhusAgrTLPDzZYAJ2QfelM7zTuiMf+bHmcmjE41Iu49q3dRaniWIOcu+hwFdYM
huMEMwGuq0D9+ETTw/U2yKNINAO6xFhuqcPu8quVzTVU+v7vba+MoEdB52N/a1Nl
cbFe6b+DIYuXU8CKorzi8/7wVm69Pc8iNFa956xIZeipU2nVeHVgHqSG6ihD5R4d
Zz+EVBqcHm60pbr3nQ1o8RvQpWWlKqkvGEqnerwSrGgrs1M2waj2S9zHl57LUybH
Mc0jMeRzHu0y1caeR86TmS4cqhPaJImi0xd8ojTevEoBwkFfM7CA0Bu1nckhjDrI
HURPOLZ89drdtqJYEoabCC+E6k7W+gRD0H6La2ie6Bos+Bc9pIyjPkewiwrxFG0j
wRFrVg1HA66KqUElOXbGhg==
`protect END_PROTECTED
