library verilog;
use verilog.vl_types.all;
entity AND2B1L is
    port(
        O               : out    vl_logic;
        DI              : in     vl_logic;
        SRI             : in     vl_logic
    );
end AND2B1L;
