`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RUwFWUch1awFxzxYUIIJtA5VFMq35r3gkWPm9mQ6OEHOyqEu4TqzZRspfGZHUTTA
8kZK9VqB3jH/ZOae0PAcfO6IRcqQZa7QyfD+mwNf+6ItSzkEi6U0QHMaU7dWz+eh
Mk0E2u3pAOVt1VjADUcRkel+873Sbb+nofoKy5gR4RjBh5cmLKxn7/VY94FtTuOj
/VB6uZpjjnua93v2vOsJA0cLGVFPhfbxYgG73c/aUKL6shTq9xwGP4mob1Aas/tU
Xu0EL5n/epc3NvWepDjkagrKOxN+13m93sMIWahw0aL4xiHySBl1l8UrS4d08Pi9
gOrc1KNBKz2weahOzGP/NN3jQ26lPcfKxb2xld5MKEHMZbXZdOScXKdc787UwhXG
MF6uQHiveRCdAcRu/ksKqCdf2rClTLwzM1iibM0tHzAkUIVOU2jTK9ZuF7gREMMa
1u0QWW/7tjL2FEo5dx2TV6DVsVOzN/CeCyWvpl+w1fC8k60yL9PgAXs7dgPg7dln
z4ZtHlJaz0VFr0a6Ww91ryzoSNDwdyBZ59b+398JYxziwp5FdF/POLxyBHiJzjGW
QAE+ax2CLc0fN+KiUk1akE8L8wuEdOEV/i2vawJiMAY=
`protect END_PROTECTED
