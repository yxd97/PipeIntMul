`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VLvmhkyLa9ycz3uoURgjdf04PAOtqp3obY++oPPswsRZb6ks/vSQxx0sxNIcf0kW
LLmnCQsN1TiS0sqysBJyg/2PElZP4gr0v7IOgw03I5W1RS5o5s+H0N4GYMyiiCIh
Pl2i05Zr5OgYbdVJnEbCzWOez/gurP+ixURbyICO9HXxyKcO0kEIQFAO6QbgKrYU
ypCIeK/K09JiQHJ/wULVB/SQJY2uOpih4XeOfYezA6lKKnyWAfFEyWiuNuf2RPKZ
f2UoA8OuOD0f5ZGpVeVYQQSUYDbiQDqXTvXB1ohWYhoAS/jdPUazgm0ByaPaFqpG
wd6bMSebE2PNg3cx7/cxw10Fw1S3PIILzv4+mytRm0qi/giFWc0P7WuC5wn8oIwg
JaM39Wt5TkrWne2tCeJSjrS6p36EWGJwCIfu96XiUck=
`protect END_PROTECTED
