`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
O7o5P/RplBRocisM7zHAe6FV3MZP4qJx0jTcqs2Fw9hcQi/xe4IUeR5lHOP5qziT
wyFYlKM0PaZ+5IzEwTv7FNFXraHfe6qwVO++gQgEzLVP+YU9FAUoQtZuOdCacZat
rbf7GTcmjtZkmS41fmP8Pci6y6cv1y9lsbW3JGJaO9ZggaWL5x9fDDtjxS2oUoW1
BEqKu6hN2p3za3KnJMWWcbDaNqLCiMAwb1owDxBJAT6kWhmM93bImhnss0VtYsTr
ez4r6rvY2GycUBxkEBzbG2NZVSu6MICSOb8dMg2XdQ9wnTy/4yEayQMzC0T6kphH
hb6rjEqgXqclDthH75fTWayi7NDeaXSwj8lD9te1XOMehMlkaqzB9ExgP8en/ZNr
f6T+kBhLwNCZL2rHoYIhs/dOsQ9uPvVvX1wwPzgV/WMScVazXwy8ispBp0KFksp9
bTXfCF74hKca3xQy/7qUsZhsa5OFqUE90B05gr+ghXAckRVZRO6Y6UiJBcbviWAK
Hi/Kh7BTJdQ8p2rFjWWATB+Of7VjI/3nFN6MqkMfCHfkqZGgcUCAhzJz/RNCWwrH
aKbhHQ2TXKAgrEo3DhfEVtbWbgnrvYGEcrbaVC1nvzz0/2d6SzS/NhpNUJuUPkgD
2LaZOEolPv1UwxTo63AJ03fnuK2yW0PLo2uiIhxhBWUeL7J/DKgArOo09hsQ2hqr
MZXnVjmqnuMqhhOD3ZccUu2DWowVlUQd8GXtb5XLkPfda0o1RCrG4EI0+CXGkMn3
Jteif+PkCGtpU/CON9Si7P887rNe5a5zU++Dz0FENpAOtxxynzY6aUsMJurcOvuV
CEygdnGVto/2BNDMqanYWGAQH39L15goFp1kyThhZSSnTxcZlprMTLgavBMWW2aL
AxX/k2w0H4cwNUTn9jTcEJlcKHdbDSOAlxVKD08LHN34Epm+8eGEX+tJdTumQxjn
rYVCp4vYp4d51t+7g4CtyBArgx5tFY+de1st/4QaMVA=
`protect END_PROTECTED
