`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vTdKkp2epxM1GtFkRdYAyCP9k8VVpR/0GazBrlZeSjYtZeC811NCkp71nxLgkdiI
ncyHNT/CjrQXmP0Ngl6u1Pc7M1bFkSLHlOtZU6QZBxSymFZ8lxoGXx9YN+Z0brqJ
lwbDd1Adl9FIYR8NTT5wmA1mKvaq4f3jsr7+uuLw+b5/SpUv9TJuidygIWXbzURn
iVv62ANtP7o8henhLkK/J13DsWMP1Nb1nRlhZVvs1dKc0OR8EQmISMijSaiMMxN2
FuAaZ/g61iXKRfnC78DhFyfGvR2aHnYbh77BKGTsBEHnhDaWzOWQAiXemjkTLuPf
GrqthsyI5bbZbxatQwl3FbwSm223z3qp8Lnmflu3Gp5BTLuvTnRg4IYdAV48Ot0/
XvYyiA++CYE5w+Ee4M02tQ==
`protect END_PROTECTED
