`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U2B9QGf7+zS2kzEWQbswco2iGSyLWY87FRTIGsuSxqPKD94ASUrFp49gXPPjaWa3
zz34HLY0TMw4CyPJQXIjVOMnwTI43qqYZly+5awZNAK/o/GjLoHbFXO0DGG/tsic
+ypyfCpRTQcG/5jWftPIN7tPX+ADHcHlyuhypnMtKlQ7RLo+OgUTI3+SwEmHgrfO
1tC/teeBQvFIicyhHdmwLHWGGrnKcxZzL3iRea9jzsG02/UudBGzc587jXZDXTS7
pYNpuXhfuQEOEGAEBJUWNxqwRdXc8HTp1W4P2E6/4UcHU/1xWeyjJW7tt/VlLeg3
`protect END_PROTECTED
