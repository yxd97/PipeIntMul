`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gK6xzYF/Ukvfs8OFqDv1Cbd5UOtNha/kA1MLGDuF6mQy/wU9i488LeIBYfiigJHX
9CsVn7casR0vWGUIKU7KkqAY3FbyAuhB7J0C4Az+uFuYHuw1R6caCIF9w6jSh7eJ
XEUEc8d+1ZkQps7Sk70OHM1VmFN2EokE/momyjsb6Yx1tIR0SnAPUR2qQQ34dtwI
+iGjkL14fdENPxlsOvhpYlw8pzer1he71cHPgYifSsnJFEhmrJIT1dpuFPiNZayW
IEhdWohsBP686SwurTCR0o2ypIYii8QwUbf7dPSpDT8=
`protect END_PROTECTED
