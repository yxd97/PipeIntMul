`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgzdvWWeiGZn/q7+aZGXDnOs4DUKuL0iFXXf0OU9O7MIHHRvsDMyZUfHRzqJl3os
dU4veQzA3r9UAVd9HCu2UbRENklsx7Vy+ZD12ED6VUkl4uIill8vJh0K47c6nuGX
KNJaVD4YZQjqk2v+EXuRAmka/HBitSZlg+D85J7dUhfYzKv/uYHssMEnPhT9oZls
/vD4MteSkoodc5hZFNNl10jBoNEZZQTyJTii0ssMemmZ7xBjZpM8Jd4Zv3CFqK79
kOsTzo/fDhh6cvY594wnYhlKaCzErbYJfbiLgkm5JZjvgBiO8AaSZXqqwDKCi14Y
U8yv5Shru/mBp5oQJNNumrgrePuGpyo0L6QnWaLNa0mFAuzWlXmhfxgLyGrKuP6L
hstEEmGW5gNhg6FiKAMaxIe3SXJMJS2AKB30F7sZ/iErVC+owgioCCqxKofbUN9E
ll0Srdbio5KJ4x7s4LqLT6m5uvoRsNyPnpl4minTILzdFQ9Ilyy7y69g3hHX8uX9
hPkpCTeeJURzsXXnSb71J1tSO4Zz4cBjdyRiLbVOyuepWb49hJU9di7UWHrCDAJq
lB2WqWOE/NV5+xDZ0vhAsGveCuzJ4UfR+zY9b8olk2AdHalSUeuIWZlx6ocRXVUp
TKSZO405BS/9LdtFhPa0Hw==
`protect END_PROTECTED
