`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cZc9zf5aryaLz7qDHhkom0isVcOUKuI1IgZDtbnYDl/oDmglGLYB8MACUkXGPADj
BV39Vv/KMalNK8idC7g52cOZogT+7uczjrCFLmTsgvwyTvnsBsOBELBjN4o3JMe3
9Em9lCDHKd3dRq8RnVwhXM0BSk3J/9KsPxoDyQY9I65PSOyeOT0mWpBDfmm9axXs
VPcqwnj8QVZBZwJ+PmxkgUHZdEexSkW4uVS3szoa/yhWk+3iWg1F38HUBLcc37DV
lG0gu68R4cvfE36YhR7XeJgFSaiuHq2y+4ok4pJk+quZlx8YFzgy3hLZ2ONIfhG5
BeFRrurGQ6ghVk7QrN4iwpNLKUiS1HtNv2wWZR2ITeoThpMsSe9SMOJkxW8K3Ufq
uazLpIhbpstGlQuYR6PUjQn1DfK5lVVmkX5Y51mznVhe3VLjbuLaslFd0mCVpzdv
LvAvjANuHmKAhKU7/vjf8AzGfA6ZIPiVFj3UB1FcVvLql/aPnOTkfwgchQvsq4KD
Aar/39dXFTd76MLOyKIJlv2OmG41Z/vYf/cPQAShkW0dhBY3QxQwxNx7imqJo33y
o6IgRJcH96VSn88JpJ2FT6r4a8JIcV55D/zFs7qLlM7zEVPZHWahGO8WY6AlqyyV
LWjrNRFrzKDLNncvZrXjOwjL3puZsaAFzgsoLQNZO5B4kB02uYJ40TGcsAs8oWDM
4bnmP9Xtu+Cxd6rsYuAbStm+ug3Tlp+yNLUOqLOcwb3yVsrwG9736zcrkW/0dESb
ul1S+J0MPHif0HUCbFjJFM3ijKFkBzsxF4TSJwBQIis2kWTK0Tk2LVJdcsQCNh93
k47PRedniABEGOS7rJVoAzPSIX0c0uGZDb76VQ09zMU19GFtvr740Zj8t2mmlZkL
p4jwiNHT4kuCCaCXug+xmuAyvLzEphq2AK099r9eS5zPzMGz7Afz7GR9jKQlP86e
XQmJ6J5d9oxQYXfAwaSp5r3cBfjawi1QdmR0NGoFQyRHMJoMdfVEoR0KBJa0o3VF
TrKyAmNvIQQaTffbg5bgW6isznt4JkVdD8albQL6NRo+V9RdkroIAXkuv2csBoeu
pm2vtPiwPDYF8tlr2Za09lPd3cTZ8b684nkBQqq8mfAzyEMnv8au6+EOvDnFvbYC
SXuYzgfqveAuIn+4Io5fvZGIqmzlbzkoeOFYL9h9Y5RziZvEJNcgtbqAV8f6+Y+A
H4M89wyLIEgl04LTXCQUDnwTuTmNaO91SZhaD9ldw5YD1CIBgwtaLt0Dxy9boPz3
EVdR22cZbkovO9xIkW6BJbdfQfZzVgBFKiqLwq3CwU0PoSTo00MZYPju/56wwRpk
VlrD2uMBKmz10mu8HtSUZ4zu44pY9rP40s0GX1VIklGMMcahP28U0lF/OqUPNecu
4LwzJQw7LcgL1BN6PxgQegfx1ReqqG/oQGo+82EVgj1uA/vqwj8dJPFE0KqoIis6
ezUix3MTcdVjqJJJIIWercPnIsDSyAG7AOnVVytXnvou7dsGVupPKI+d9xjNVj+X
tBKscciVtBKr++Ud+lv3jnLeSc6ze9ULDd27PhT8Mzj/IDGOuw3EjiYVwCSycEBK
tZwHf5P5tUmkOAi9vaHD0oFwsjHp2Rl50wlvPZ+/KzCYQFJC+xvnBeDptGZqD7g2
ZfCRVv7NVQHJ7pew21tdywrepnozAXN75JPS7v/8NTMmMIwyxxj8+TtqqsZ5f9GK
9pkf87Q1NKx8a3pIPldIE9CqcP8mJXGC8HGsLSQshki7TQNEKoK0oYVO6FyDdcS6
5zCUewCeu8WheoGuKIcZwoc7fACHOnzzgE10mN1GghzMYfzt9FJ7HV9tHlMG6S4K
YvAwGUXddc8myVVzunOFe2gnpSKN8VeJ3hmGqvGhINMoM8XkDx5bQ0cTnpG2fMYb
sMCvCrdrgG4zxR68xBX7cbG3pht+nCdMilVJVFXALx8RSQ99Qp2GIy3ceo247mh/
NbiybBNJuEjiCtJStC/Q5pvTKWLJHEw/0Tl2ufieFrdznwCtmTcn5QpvuVeNdPQ8
0BVHD/+a99SXomqWcbpuPndMlVHue5mTJS4x4nZ8gjFWpwg4Yzm2Emm7t0bJkjYP
IAVlbtv6BXR6vR+TAFFtQekdPTpIU4xXf7SRgsq27LvcVJWsjiWIEgbsYfnsdXi8
mUyR8kW7ZnU2Raf1TNc8A/TTgS4AISy+EPfP5YwBDSLIFf8KZwm4GzZ+nHyZR+GF
N/yR8mXo2AyxldTV9Mu/fEb5C3+Mu6bhl53Xars1DpD+K3JjrFHo5sCZ28NFVhc6
A6wKus3OAyZIBO7rzoIzg+tDHv9+s4a+1mYee2+cCo9/31qkgIW76TUFkF618SDv
RsurDtKWValG9I7ZzUvnd4syjGO8rEDuSnYWXgHZulUiwUdEhc4cYlgi5AG1JhtN
Xk21ETjmzjrnuh2RztsTloey9xNPuK9G1ys2ULmuKa9cAulO3swSr6Ti/JN8pz3c
8J6ykNBujQlATTSfTWC+LaZtv0ATeyK311lZ9WrTE6rbwv1l6rcWiWjeC2+VbH6d
tqKV8LtVFX+cFc62Jy8Bv8KPnPNGMYhWqgBcstemDImkMo6QK6Vuq9sxKvheCjHY
CZr0K16QTPnxLEFvP6puuZp6HeQrNuaY6uTUVGOeawcTUSSkAgn2ic2pAMiEKiK/
onC88av9NwYzd0Fd2o7DPdPvyFNH8jWOA3nBcacM3ZMaIg9i0M7IgBySWCdo2RAN
7TJVac6tf6pz4ekm+vRK3352t+2aMyYAj8ji1/eBoeFpMN9xfUPAJAFVvxWhNTyt
cGlWfu+INFTRfFP/fP30pP6FSGutFND3znytKZujybcMhpo6xGFpLkW9k7HhFbix
3hOPnHbtaMslF6z+YHyx4JBrExC8O880NgLxFZmIeZKnO9YEgKXcESy9e8gwBFeJ
+FLMM3EYJGkdM8AMuK3dCO6Y8Wfj0lfwSNf25Hno/oWBqze5DEzmsiqX+ff2ywmT
3YWh8P4Pk+B2cFvmZWrAVv5VKVT9i9k4R1lmly1tFGuhOeMSXe6atoPcgT+lwbbu
TIha8sKBPgXH/3lcSBuXmFpS6gfjx9v3YMN2Vu/7tddY1j6s66n1Q9k2zCn4j+/Y
61V9naq6rLKHH4TzgpaXg75jmu9t7iNNCxk1YY5d1cGQc1pwOZgWveMKpnq3tn5u
V0wqSmq6mivVTt+kjxYQ7KRNt0pla5bB/Q6yC5XHI+DNWwTfmu82krFImNA+Q0+9
4jHvi28UzFbZ6CLtBoG2U7Az01k+iuENX1+bP/+W6avgwjaLYOOzSpWqdgTxsQS9
TrcRrE4bLENO1qZz6CviTok86qf9Pw2EiUsWZnwfpp6hNoyIE+Yn6NWh7N1YTwCe
t0/8c+Jtqz+VBxXEgcpUA34L77lOLUOE0LL0nfE8QqBy27EIBbb8rm/sN1H1u7+J
+IQqFLHXb34ch+qhLsW6YItbI0f1Rfq1FaHD/PmjPNJ+lVaWSBdwZQWxuy0pFcgs
D1dBsMEuGIeddSuXRjPnF8avnDOeiSpOjqwFp3kOQEVrLzddS8jBrplpYYkGlTXE
ksg1QsrAKf0r/aDdfggyE8bvUNR+F32ruMjJcbcFOyDZORPOc4wQ7BP4OZ74py4d
3IXVN48XUC2N26hCvkbi+PJ8c58PlTHhGKvBtY2KomiNuCJ7Ku7m4r63X9U8gaSP
lgXa8xAPV8XzQqWUaLPxWZ8FN7oWiIrbfoGwZTB1u2xBa6zB52qujtpmlpUC9DE2
Ee823Yu5q8qAd7jemfTrQQtadLOnKvjNK3Btt6f9IlrFu5PL6Nn3i854VYyVxxeQ
RxszPebFe1RSVExTkhassJd2I0aDz4XIhgStnbb2dX+2EVUn6IaMfz4kDK725Biv
oby2mLrdnesKvBKg3+6XRzAjAUjIAbqwOUYlgIetcdK8ZZt9klZKMNsFNZHAcjc+
qOhR0U47uJyBg6fQSORW9TqSEqLwb6UBhx0AG2Rml7mWCk/79ekKwC4jvJfUFglK
FDovQt0Q07kKXW3r4cRl7nq/3ejzmZK9nXLxxF59mxntl+II54N2VmrAdgthPKSL
E59wika4jl1ANryMP7aa8sNjIKQrtbOIp8JPWlWKr/Gx6iLYonmp8MFlixzi8ZJt
pyd8rd3IKjI/PKytX/DJVyeSgSUtFnTERIb6x8SFGU4EW/oNEcUIGDa8IQ53iwCD
V1ZRCSeMln7QnX6j85gSH0UP4TP3dd+a1NwDqN5pVh4+YcFpc74nv+K9ik/LEF8k
VlGk47HkRPGa34G8zBOEIH5mEP4jR+rxYHgOJSKmMB+MLdTIJvuG8tfNLcKy4J/W
+RGtEVTAKyGx5yoZhTAxLXOaYDyfccDIyVK/m+PqboKyexP5DHEE2SA/7Iu6ExCx
nZq/sghcAW6dfz6WmSFnif/q08KxLk/sYEhSTqLJiqJzOASG6xsMTKx2d51Sxprf
tBbc/batCyrdX/QjNHGknVA1o+1rtORqvtHOqD2qOfVdPO4uoFLyxPw6hh/MLV1V
yWnzCxVMSxjeoRP4vpIzb+pR5pkbmXQQRACSD4VO9JgFG8ot0neTPq9mzQIJqtQK
oZV8oiCtd4MQDq1xjd73WxwmnQOz58UdCkQS8+IUo33puSgHn7zd1PT8vCJH+9at
ycNkJtVmeAelqCAvVTU0dGJusNCe7J10Z755hVWqOv1ALEjLT9907sXV4uepMOzi
MOFlhb4cnInI5hc0FfePfK0xkMl8CX3JTXDIeJs/1IbGMfYtTeos8Itybi1/m4do
Iux5tZKi/A+DrGXafdMoU7d2oRNGCruBHaP4ulfo2ancszca4BXVLegE4ZfMubA5
Uixx75FY4X3fPXNxGX5sjhwkmF6RaPewiV8jkCsMz7r+laA6liMuPhXXutAF0/Vj
QmXDIKG7VANNl/A7goiBesU1rExsTlOF7ed8afYNxea0SMmtJ1mxzjAVLND2uQ/w
tf0P9cNpa/P/xtGyWuUckoYOhR2eUTl+XPcBVdK/Lv5hBPknlvZ5gx43avZ8dzFz
IMkRTWR5rPBtwgCV99TVfT9TD4c1xUmg7ugh/va62EvOXlu7MI6pf65YhatIKGFX
Gl6Tc9GHZTSVilwudmDKD8X6qsaSCvJb5Jg8Xs2LSWk1yMIdYqwWQisJO3dbse71
k8oXZPhKVUG118zXDehbk4rIurXP3JOqa7kLSJOxVNOuDpp1XMkRCbJM9kkb5ttX
sMdvGFtvbKOCIl11ORv/+Cvc2TMaDNuiQvSQhZf2zqyV1DvWFIK5FbcvLm85ga+W
4/4jMxjvPYBKLqYaQUhFRyH7Va/U6FhrQsB5mT5NQVqGQAxAIypehPax9JWGPlUx
2Gd7/p9WflObzvBzftI5iNU4rD+1/4i6+AuTHzobnciHexTdeYdD8UGkynLYZyDA
vVdIo2euRJCx4trz2ZJ0dYxDBy56YGRPdCaX+PUzD+HERSvaP1tzjozs7cwIdoPy
s0/N9TQFVwetcMoRuOt78sNDmY7wrqf8dyEbMxoi4GhVmTlvyrvhe8aDM2/Ubuqk
IfSc0S2gu4dfw60MaCAjq73DI/p9TkAbKvillOIAiq7ISfFL16Fm20Bz4hKBlrHy
t0x4awzUf7KWzYr/WxHEOx3zMHtTa7YWnHevJpKIDWd55ATO2fKSKcrscCzhfbQN
96gEy0sXt6uROH+J+qh4OoQm9Qi6foUB+pxuhOD7TcsS3dQUb5mCi8LobxwS9MaW
W8oZ48D3cMA2HTg98IXgEs+2r6Is3xtf/7XtLFQyINHYghre1VSh4B8dp16h7D7m
76YAFeHkx3cCM+H24Nyi57RnXuzWXLJqgWxZKsfFmEWEgXSBBQtbPoMk9WXk9mXZ
5kZ9cSZOspqtc5IyJuqiMwn6qbGM+d5d6cYNweo3Rpmi/2imLpp+Ge+NlJL3a9o7
u5a3YbkwjVyI75E6YsaJ67rOX8ii0EYn7MlEC4zV1N/P2X25eCYTrTzPZ+x/L00Y
z4CB/xC6FSb8n6wsP5d1iafjElZlbfdk1n3eQfFHSHLWOvOg16Yf0XXHSBzkxCOf
Ca2Fq+vctHSGT6UYZOuEVlQoqpS79jKPf4oMhL/Jl7u9fVun+bJ2Sy/OwsKATvkh
1o/lpO0Gmk2ab0pNPFToZL5u+gwA+ZEOT0WVnoZ+Z4FqiATK+ObJzWalbZQRp8hF
sSQPuWK5tEHUBDUj4U+QurU3EYiHD+bYTSKGUasy0D7zvg/hLG4DvhRARKcUH6mv
4B+QkSzBaqWw2hpPZGpU1BhyzoRnuMH2dEl/mL/s7ax1c5Y9XZqOKfkWTJjXBMRU
HkWXyBQlQxjjjunfizpwwgbAGsCb2qONJf2nyOaJ8UYOb6d7ZPqmOkNaD4xyThGq
T6WRJ5LPXoGq/Stl0U6a1Sgh1t0I7lxGYGQAQkAlAxoYBskwiD2ilxn0jHWU0Oka
hfUQHXd1b0N6X1/JvR9VDAZZ8Dm1gZzxOXIl8lT8d2/HukVDjDS5OumeGbg4ZmQC
uhWQSXM8xX1Cz255jP6szoq/hkRjFTm1Rr0eKTdMlWS1u5QhFF5+7EM4tIO/wCoN
J5KUuE+bFLbeD57BBk7sWDQ4Eo9b1G6asXuUFJ6mtt69w8ILTv4+zeNIl6thArwC
Od9+BBOUOtbZPTAinIOf1bFvRJZTBbetiQu8sbbPyGkavzrBJCjCSy5sLC9D9A0e
hUSk705J6Qx84/hkShlVsJHUnyWSF2cGQXs0h0hF6cSI69mr7Kz7cYnUSTyhX3tD
ehb9VmGrNyuXZBliQaEi+FoPzfYH4Kfo1Y+69SLqNzdZP1QpuayXVdXMYKPTdlFo
6oQBq/WKY1SEnjWjATxW2zAQxKjmSuSuj3vThD63nG4z3c7Z2UBdI9jnMXsKZ6mq
5quep5jhLrDfTyB9RZ9jAjMi9Yd/tYpPhnj3Vixg+Y1TkVKDB1L7b+cLxEgdG2wE
NkZX3cy2Ua2rztvaJgm5VNBrOw/QICqSoQ4xkV1Ofg19QA0Qo4u7NEGLxk4QkI4y
bL+B5ZW/UYRtF+AnBZcxh4SbAE3leb9uV9nihlKzvvJ79PWaZ+I+qJ7fwPVPAsQj
6C/611EUi0yzg2Nh6CHxfevhZqqWeVvw+gATfFm1aPxX1WZdSAkOTA6RpqwNyIMC
skjv0Q+S7SSuFeaK04odQwohhvL4MTRlxrvLXPx4sGDADqbjlMYVHHaTBVIhD84G
RqhH6yKJdm4iBq6RDY3F99UZtD9OXZmLT4PkT8Cx5rog9jylbeNeTeabGK/WC7Kw
KeFg60YaR05xMdc0CARmSjghjMvgdst3n/dbOCWg/QedqWOgzbtZE8wLy5Lv1d29
NOI0bDzO+iB1QQouGUYPHmqETsa79i4hwOhmdkKHyWp3mJw19ZA+Ut1lsMib9Q0C
jcH/x7nNYtx6bbGGJQTMJUk1/8kd3fND3zIv2PiNDnywPpX2jhdzSfPzcgf3LEdy
GMAT2bMD4QOIsGolQzU9wMq4Uapgi5rBAmGH9JMpQDyfNx3ZjYijSb/X6UFeoIoY
Z8OpKTIMKHAiXfEX/RACx2fkx/qq2F3of1DChhbsqDbfc0rP2nMjjdOmU23MEaeP
j4a6LcjL3G2XtjFCboOqLcSn7lBTX7i31Ool1bPG45QZmqeyf+wxBK+wRtxwfZBl
TmYkH8FMz16Oo2ltY5MOZx1iueko1YL6PpKYBHbhYR9TNvCB87rDknWOgEem4Fu+
BjrPZg7Oq9xxJPyXHyZRumHj3BajeUfO/TxGcoy8crd0YUxufEQJiWLxDQBFu4vH
2hXNJLoqmv/9UL7vpxJfoXQmncOcML2wCJ/Zh5FakP6wKaPzSVowQTmHK4irckTv
clC+jr45/LhKG1Vehmk0ClugGh8KwRA3K9+uvPZNsZGxJc/Sor7/TmbebMxZMopu
Nx+weDvOwBlET0x0Vaam9k8q8+C30JdzVorbNqCEx1mqUAQHox577bcfbv+jqRJr
A50yRjr0Y5VaA1JN/t2g0NwL718o0+GeWhBjSxj+tW4POkqbBsgv8ErZe/Xzj7g6
zdvqhqrZy7I4FX2AdQpSx1woDRqo3Z+IOR83yp3qE14GZKiPTAnl7387PWAxsyna
0vLcLC4oJ4cxaXOvVmQAA4Hz3Ad0911CMRTEBOh1+BnS9thkfrh0oAeVuHcLDzmD
g5h5LJdVByjIyX9uWaV1uCG+UWEoFl8DvTiT3DOePFRI62O5md24yBL9sSZEmh6C
JZK1SwhsxwD5wjDJ97PwUKCQOy1mviNnd3tDeV3m3GKHRy8QLnbDSAl0QDdDUeql
Lw+IseKp+vXSmIE5fL69yySzsqYMK8IUEgswO/URPvLdMBFEzb6JONdJDuJttdSR
8MM9OjB/GMSbuq2HFN8IQuFLDq9DX4ieWvpjAtiaC0viQOqOAaJw5sLEWODbHGn4
xgHVO8iK18YN4iH1LeQ3TPmnzu6rQLdZ/l/jZGpmNETCN/y8UGEyCh759B+7eFW6
4c6y1iA7x9wXtP9iUwAijdsbPpl7dsMnyCE6n/zLDW19RralbgoJaBCz1UYN8MVq
gUcysuyZQRxmjEkzYd+pH+pruh7MUXbjasJ/7RCn9xTFW4mqBUNglqyGwQWv4Rwr
NMl/jFHO00S/9hn/lajTQJKzdv4/U9/fWA47OYGdMP00Z19ZbTJgGRHOT6oOEdAh
xiBoeLvfde5Pk36RY8kSJxG464jQ7Lqp5ns/mW2BRwOlQcmbg2JdHxUPwb4wajAu
eoj5UiMb6dtjHwhfrXjKni+2Zym74dxxgkVH2qWDFjIUi/hmSitfK7JPy4iVNVWs
yD0ZSsbLtY7s2BZlrpuqXdHfr4bY+JshOWVtNpkSLwqmW6S3cIjPOZM+Gq20d47Z
AuQkGfqYCUnmlY5Ibpp5757v0DjT/W+9mTyFwo9s9iAAmCeWOK5Z/KmsN5+1uyCH
RK3i7Rsg/6639hw12K+0JogZ9Twz1mfQL4gs6kkDiJkAjFWpb4Vp8phmcrJU9Igv
oHacvaQCK6furzLtdzXqW8yLDr4XTukL/R0Lit0b5m5OAtH3vcXUbLb/LVT8dTy/
ywiFHoEJsVFjkCfoq6UTjKh7gDJHhv8ppPozmLdhC5KXQ1w58PjOYtMKZCXrRKiL
TOrnKl6r9bcLeFBAvaQ/WqYFE6FO20GwDc6zw10C1NQI3UZm55APYeqQiQw2Z87D
GLynybiYSlOTBImoY1LFedrtq310WdFXTG0a4bn2vzgHQoAXqJOy6u0zEvNK/O+4
hP4AfS0XlxCBM2eRHIUQInh8IhWUS7sr69Lj74aHuMisZaRBWoRCpsmTyoYHRB+A
Yzo8gUqosaEnvKo/0bkzddT+1OWC7XHiirN3WPXlmVLOWZQymawMg8SSzgJ0SQPa
sNGDRnUWcfupkdHyI81a2C+RDscWFNOgQ+eaVPboB6m0InM0nV3g4yS3VBJ4ehIQ
/+3vG00IQJXzaiq/8iCQcF2AC6IUhnmCP9/GeEPZE/LaBzGRs519LJEk8BcAgjAj
/0On3I2oMvA9nAl+En3VGM6aawi6w7UpmNGrCBR0URH3zkuG1ys5Ssi057RoyUlq
+GAIasYk64MIr3C+eQ5qDylmoKP+OQyjxXHhaCJETs3SXS8oskOMDmoWywbiuvXi
dv4T9v7uTtW22I9MFVnwloFSuC5p7dMVpAAY/bFh2ijsG6FtG3nouXVuHq2tl4h0
zpqJxki2YY7lOTEHo+uIM8weCi+0VpAkGzLkpKJVYlq5LQtx4iXtFy/dthG64U//
scag16IvGol47XDUCeVWNPeJSnz+GMV18vGHU4u981TUfPX4NiGp+cqpFJSfPPHj
+zYH+iaSkxXEPY+xeU/qARaTE3rK6XoqcHxRj/fBDWr8EKCLmLYWyvUPmHHehF/5
RRErnkJZjemg8n56fY8jcPoKBjilF3GJqykIH9nQaK+CbKj98JM17T4dlI5wQDQ8
FQZLlTGSaZmKhKfYeKaCAPvTlkK/DVZZEJwc2JMF1IrYMIeCeU5frad3lPBRLOQi
MuqGgJMZZGaLQS1jKofDIJOK4XMamnwxk0MnQfGjqL+I/7RXCO9d7AV895ezT54Y
Lu1ziIohqnoWy+KdSPYTeLC6ce0Lsa2aME1tlqu9ykdRuIUtuf6bY78DvZZkJ/8u
MgS9HnxRyVdIFGo6vwCQG6W3yaw3gVjrcyIMPhDf35It+FGAjs5+fUfRvsQZT7VE
yt+gX+X37SWhS9pnbi9dNFQ6cDMKavgh5LV5YKG6uaplGME9y9OTyUW8QxL7vm11
fy8vxXKmwYcYjT03K688PHKObYYbU5L30F4buFdeZwiKrZJuiPYDlqxOlBzMpAZ6
bUUiM8SqNlU+ntagfz3bYfejbgGLK0pxoBXDhOmfz+01+Z7hWqCHkIfvUvCiACoN
CgIoWsuD3Bd+zd6wTY+0d1066EtS2vIKH/1dVYSv6969DboLnfSZPKKVPUHQd1jB
utI/feummSL2mQJ1Ce4+1xXstowQ4JLibohngtMsy4UFLJdKZJjhVgu4pqN9EcrW
CrOido5HXA74QkMLkblB9lBMtWkrN2CocDFRuo/OY3sg7zwhCPFFjXPRLXKrwNWu
v+4II3wmUfu+97ANGCUW7x3NYzFZuVwBq/ZTwGVdrsi48A9atZPC9+OV087BdaWE
OecJpK0XJi9gATN9Izj5Cv9DWLkPYPU3yhdR5IagwLpurbTDdYMIiirTrCoCsNWz
E2fw8b0HbN/awNytiYIES3by4JnXaMb7NJzftlPLCD+olGDjRsBzC0HW9L4zomQ3
lhZUCT4lDKWj2oWcjcE6v6WSRwC39jeKrt1gi5SasfRFU8v2ZPcWFq7FyXrGbYY5
aY+N4/nlm/2COQHvQugPnVlv+6BdLOEyopUD1pd4UW8KP69PsI+QFAFDvBv1kEFu
NPBje2YIye/bOaMlpU0XbNyDkBAkNgkEf17DKT5cyZFfJFL7gSJEmZmRYGP/PTHk
JFx+XtCpaH/ANPtLztMUt+vtnGYUZRiTIMO3CifywyWKE/2Cc7pBDYZPMKEyNvZ4
ZIZ8mfp5YUBKmgotZoFV8CBfIWKrEK9DWjWblHL0B+fMIHwO7J+ZOA90gNmvnoc1
kiSYO4YPJ0Q8GZ0ShRR9DndBoTkzsB2cMSrIL11kn1+9JKcTbibnh/ojJfU1btev
SnRnpqCGmgOZ/2vkkSp/8QSVB6Ka83hHD9su3/ANGl7t9ksTznHfoC+fTBNSvhA1
JOLcxiiIh3NvCJ4lWe1RQuHrFDszw7TndbXvsW8oIHbOotPrsBDZOOukLnvQAHCj
lMtEldhgP9v0/bwjWBRUJ+SxrX20SLO60Dg76boA7M5ofCMRC2gmMwPXiKkDHrdx
pjqa6ILBPHG88n5hNBNLxhdN+PCHHjRJxvpepVypezY921o5cxbVn9Mxx9ltgK2h
sVIoSQTwyjPUrSkEQmMEOKpLstkDR/br5kpMYdTBLxOzwi0ogara0T4MppzByEWL
H52Qs2eeT+tWawv1P4tnOwm++Uj2TwwJcb+1npqRqVAICsckZ3tk7ADH2zZLJ5XF
iqIASv/EWpZ/TW0fQLedHHwtsfV3AGn0F3IJEy4fiP01kp6MQgrw1VcZTEYG0rrT
o+tYo3/av9FlDCeYtBfSxYDK+PS5/HffyUV/3zGifGRuJU/qhKMZ9tX+bBARDwnX
T/G00ubnnM84Kl5zYZCu1OI9QQb3SrZJVGlhRr8I6F76B56/VRy40ER2LrVSn/84
3fKdRuQSgqKLfOgnHLwZODRl3AJ5XAflwZ+Y5lRjquU71S0qzyT4yhmbR+gjxhsu
vUN5mGXrXemWfOFxm0pfbHhycDboSR0tvt5GIemhezORnL8nfRfPKtDEWH44Jf/7
nuHMbhp8noNNKcHaMxtD8mI22o3xnD40r28iCg+O9WDxNoPJR9mP33y96w8BOM2r
fKR/p7H9mW3nZ00YpMEvhkDK4YkqREEYauELwBsnVhqCcI0Rd2qAZVCWKOFUkVCi
/uisoGkqcLrYZV86P3grlgQH4Rd7WJ1WXMBTcj6WdAsmhjeBb7fJCyGimTLGhLoh
UGA6ajqtQc6OERkbvqXQUoRaQAEKHKbb7MapzwcdOVVEpUz0Rhe0J9DfbtT+FtR7
CeoF0EAGD4zoDhPLJtwOLwKX2qtcVNcjEZGgTXgCuc4GSPOdS2pgpai8BWkG+5eR
s5P80eaS0EV2w8d4TmfeTY1yMD7zCtYycpDZURdtkgMu/7MkqbVHjYQZKvuTTDoZ
yttnb3YgDx4+UDpfwuVjsgx5NqZSouw/vCB/EWAtE5V1awHBgBT9IxDHWbRQ9+r/
eWK/alKut6ZJTWbr/Hbpsm4oFz7L/Vy3Twyc+8ZjUKpDOD1eNOKpqlw5+59WawCL
F+GzcqEMf9InxyhIeR2K+QelBfhtifo69snPqvkiJm1q5fy9ubcj+TpD8y6vfnm9
9mKRzMY86qqXyHy6vl8UR6wXoXQVxMkmsEi37Ci8780Ew4YDxgmnemhZEquyJjtG
VV41E8yXLo6wv4i5dCjdJzw6BFNP6QSfwm7Ey/uYPBMTNTjZMteTbklJhnNQE0B5
cEWAM5wxzIsBcpbm1Ui9Oeunw6ktDK1rt8go0VrTflKZn+mdSvf95cM7EksBYNt5
Trsrft/g0lR19ef4eSlpXoP7S//5G6QWd0MPDDahsYEk+CwgUT4Ronuw8L5iZXud
IKtiaMKuy/lrfbkfvcoe9sKFx814K1mi5qBaLcHTDU+R77qcAWYTP8ksfUPsVtg/
rvzNv8G6NnFTjnZNmDdoFKVT4VaARBT0BzqvchwYfOstFfhSAYqeeTDJ7HSbghoA
iIZbbd6fl6TGbhC7Ei0e0wDs2DZRUmx2rgYJMGGAGO5oVw7OKytx3jaBTIUjpmgT
8xwHnJMEgB2qEelKhZi+uqWZWILAgApZkJ2X5/WezLsdm30JAfztrOCqj8KT0+Dc
tYCpQMoLYog0sX8ZI3uiTDxPD24y7Qpch1C8GFtvjVNhoGE/X6+ESa08Qxi7+P6r
iJFiUYhfUjM3/WxzLHTSjP+O1Z1UnhibicFTRUacJdW3GW6N02iw+S4Qf7iit7k2
gpqDJ7ja/rUMmJez7SYVfTaguJP1YX1JRYHjSbTZQrm/bLp8VVtnfdHO0RVQ2hMF
3YbVluXYxNzI0ScNdfw8GQFigbYmEInurrlVlZK4sDMrtZqwHueea38gTEC85T0Z
6S1Xow7m+6oUgNAJb1elkEu4Mrw/1t4lA0UA9pc2tBBx95dW8kzI79wuPJfsO0PE
d8enc4qjawOM2qne7+HYthGMpCTSrin5xK2oeU/6lGhqEzAt5HTR755j4i5Xs4cc
0Z0ZKPzxKTNCmltEVTHQp8Wr84oVGQOEwr3+9oNmPA4kj5Um7l8J2I22JSPdo7zI
NNTunXxrzRuEhb1xCIsI9kIJFLK21QiAdtqIOSSq8ptTlvWqSG1kWCc5rQcU+7cM
hGPZ35CmZgIJke1VspjD9bSUIZf+rXS6InNXgp+btdfAROdQoEZkOz3fnnQdWwoA
umU0hZzEKeSjkX3bIgv9Pi+gJ6yzvN+/zviHOHb1gNxoNtH5P9dN8dMfR35r9VKx
j9gIEqJZgRejmPUW6DSAWt14i9jyhUClx1JJRGJf+sqAEQfyJfATwvrVGVud5JjG
Up9YGWGppEjJeOSb9hvVbQvs1o6g11NRIUgH7OvZ4meeM18942YIV/45tUjYv9g9
CzcXp1pHZh8Cu0+tnQBb0cJKI/Ykj4Niu2bUHIZjE3g/PZEILds2lhMjH0Gb958v
eaSZQeU/QPXHufIefp8estVYFmQWFfI4urdb3dIQFgNa4/yiSUS5nDfw5eQGKDou
mwcbAPzP8UOEh20P44cCaEcCTR9klx99MHeOO0EPxNoOR+UvExKOUi2WpIL8yK2w
BDHWfaFV4YjLd2NOvstdi8Zeho6r8tWbjOa2u5GUEPYP+OTO5UwkqJnD4OwGaMj0
V+EyqFXq8eZskctuMKMBIj/t7i1Z8juv+s0MA70k9Ad4RvoTS/KzntjpXljkCpGs
uTWpZIbNxxlMFPtAFrBjXSUGC9oBFs6COO6Ijpjwi+Ji1XUQSykZHboGN5pA42QN
rsXroNNovKFk7i+4RHPMm6aIRjd+BFgnRgy+u0e4jmsVl8Ir0vFAZ/ux8KCmrUf/
+S5k52/KyXCf9E2k/l3zFrSeQ4lekAVx9ceJ60DwJLp81H+mEBAH+Yh7R0vUxdcd
aFRn3bs7PgzJoRaV5IREN3sJ99QT2yf9alggTLYNoyMm2ypTvHe7BU1/dBK0cIMd
Q5s1ZNJbKP1LdhDm+rFgfi2+z7ZHy15BQ9g+dSKJg/gpUtl/K49rVWJum5yxJf3N
66X9sEJpf9G/+efiq+AOeGLysOu+xb6GgeqDgmFvNV5u/RU6abil6dcI6UE3N7XG
v/Roafgn/gLQVlX55mBTj/AVIPhZVYroUSmnPagoQ0+tCRUW9vkHrshBhdJZwYaJ
XfiIwj6zwmezicDMFKwVPDq5i6XRLDf0O49A5w3OKo9JDbgogHtQ5Jir2XE6hivY
5X0a3upfyFGoH9ecr60x7sm/+4EEhyvUcUWhjrJoAprAx13rLY4LwLREydcbRvZB
LCM80RphHAwUsyMGi26R2eIi7TERkwy64Kv5crlEw3hk15KoOgBusywKlvp3BzZU
8Sjhyb9ijAatQXeJkA3WOKZ3oE2mo4fA5aHUbJ/EkDdJ/J2X7X7bZyQVuhdG+tYX
G/yUPVzy/Ly5Q6Kf4QStX/AGe5/dJyX5ElE6hzeD3UhV6LCLXDrg3Ae7UDM4kFXK
LWrxlExhEmxtJaTD6tMLX8qKHTKI6o0SqY5raE9qhWY3xnUGJMgJnVmolRPUTiH9
yDZSHwrjuBW0mkQbi6bC4JFhrr+0yaPwmuE1xgxGz+5GRlCbD/lOfFXTnyK9bvum
SpcDtXx2A0xf1cQ2JSgnE1N6cADbSn0mBnzc20g8md3R5m4bdM21vmyuOsc7ueOE
h0JfuwDwh3YSTgIVo3TBqi2krnv4R6SzeAqgZwcH+SRCGptlZO8YN1Y/XmqznWzP
xSwmf7lgjPVJKURbUJxFWNaNNYl3QSUCQ20hVdrJlLw85cB0XWFlJiUD0z/3rIpQ
o9xB/4151iccf8/J2P12AnWw0wjQPyZDtL7+Bd3U+EEWmNV2+MJrr0dR54c9epTP
t1lTYZKMhLO5omGrVlXr+SJ3ISiht8n7VI39RJxagCtxSStRN1QkKMjY8fHVrQe0
ssTbHBu2Q1JD/h3ha4B97W1mbOEyF+FuHrf1k/yy7L5f7TUJh9nuBMuopQJCFJBn
Px10HrwInELjPKZbmwnyD0hKWVF9wOgo5IFYBedpvsEZGJu4L21xExROLMtHqbJc
UbwVKzpt0WDgxL7SO1dMdpXh45bwF87LL3aDfEdzCn19YKdOo7lc8L0z6Hbfggzn
RjzRYV88sGnP0o2uJSiBIqWyVdEzvOSIt1ycKEASPZu+Se7emy/Idr4LrFGz8Khr
xOLtN5HBl1b8T4jtnuQMgMwvL9Txqa7D39a1vk0w/vEUXju3GN+jDTw1sf5eut0a
UmAwjD5qPhbZSPXLVYL5x+MEACSRfZX0nFbBGoEArXa2EciWyrnGxQNJ7LelRk21
vnMHcamRsO6ePi5DuBapHcKN0sMU3XQTJBaV5QisgpILysFyrHXhIhxGe9zkSvfk
lUa25Fod8rwEDSQFTvUDqiNQZ4qq7DHOgAL/rlHol3b214pW/Xp6ksMc/GwyMCjg
/OEmqZbyvtzOPh0BLTp39WixS2Sa2iBccByV4cq2DjpbPFCiDI9w6pgv/VDjE9Rz
elEQ6Xkl/+ZMKui/KDAOi2eJSMCf27cfBmB9m20QInuw26gpYMHgMUa3/W0LAIEo
zA5tLzmjDh7vX4A5Q1xY2BMokXbYvCc+3mg2a27dSAkO66ylE21clIK3lhoJho+h
VtIDmeH3eP3dMUMKBmv7N+LqkFeVmMT6alUglRiF3vkPunwxGYUTtohv7o5O4SSv
hptzxY6VuwNVmT+aI8MWXdzR+bls2x3ewTm73YAedgNxUJMC50lA5TqKoV+PK1qv
mWqRSJ5kfZ4JOmg2pcu4W/1vcac4PLImIR/+dhoOBhXRnrAncUZ40ZhMVXxKZDz/
caYi0eSXNAfoUsFL/BTtzMvQRaGQp1igwsDjAhAhZTk0hUVty6E8Cm0E/U1/xO0a
1Z6XAe/LDoa2y3AZ6r/lF4Ge2EaTN1M6ZFupBXBzjpy8ymBl000psmUcja7Ds25x
p6RdjJ3pas4Fb7nUskEPR6IiU0QTUOIbYpiQKzuNEJVqV8pYJ2K1dZWt4HgKooX3
78i2FovTEsO05ld3xYyKJeDLle4KDMYDpVayBCgoz0jw1Zg1Q5uGcpvuZ+xd2xQm
At3LatkDNJOeSKbrBnpPBNZarWywGkmzG7uuFFhGrMEpo3vUc5gvamTbsx8d/ZZu
n5eOu84bSGE5qjNCebXh4T+jRebqhRLq/IQk7PDF0uuzER5dF5gpJi10HZlORZDC
t6e4Lp3vJ4hFJXAi7Nejx+wGWDl/oo9dG736O2oCZFAITG6PpJf+QVoycr7VzsKx
J6Ny9WK7/UvzKnI7liWW7RgfFyz88flxs7hiyPIwd6hcPfFJFZ9W4v4yVtWeyn+/
x612WHb1m41qlLj+TlEfNod0sTuKUx65Dz8W6UY3GrK/J4RuO7IIjrrF6LJF7ift
EgS5mORhkjPAqyRGnlEEp5xsnLelgfkW+0x9dpcWlB/jJLwKh5NCXqkOJU4ZUVKl
kmFW7CUgJYhZbkY5Gfs8P5Cf3tRX+TtIqYObxUCLdRhEa5GeQQrTcdEzIMTtKMOA
JyfQMWrQ1is1dMyfP6rbYdJOxUf+ygGYLAPNozIVJypSAqn0D7D1VZLBg4hOA85X
A+3q+LN2k87T7r8p/tjs86C01TyUPazVSfHsD0Tfwz0IXHX6PF64wePUKR4iB4NQ
tOPj/GGHmRlzof2rCoOfIF4VYij7CvX3n6tKSOfvY99kXwAs/mlw+oWjm824esiR
3Kl/jp0uLSJ6Wxs53AY6wGQmemVp2OIPvwdYSc/vSRK22mJe+cYGTOAsD+yfFJ6H
mhc4kHFxMzlvgFrJwOWHXpVcpXVKT66/t1yv5ui/q8XJ5jQcV17Rttu9L9qJGbVe
BgWFhADp8Vwgrbet+Z53QxU7wvnYNdX+NC6jmjrE0swcHSbQT5sUtb/BbBOmD4DY
cqdTbidW0tce/3livJwMf5cueG0E528u/iGuSjaDV/f8+/zVFOAW3R4ihsimZP3u
6q8xUVyilLHoSNfZp6Eq8S83Y3N+PH81kLz7GiNaUXNVkkYhsjhYPgmH5BiStxDK
dTVuJwMdhfQwz1BVR9FY3dT9P5Anc0rZH7tLHPiRUzADodRKIbM1DwXZ9oI7rh27
XH5V8QnSEYvWIzif88GCbXPZcVO+xruHpIe8SoTcrQ96TmVm3Fj0Z/6VTNdwmF1k
NmSJA4mIzXBuwNkDVfdzsR6IVTx6/1NjfJs9r/DQSfc5uacGJEBGriFELLJWi0A0
VMWSkatGR9uXYpgzep8RnGztepOxfNpOdudBl4XrqGb3ZoeGQ+JY3MBtP4e9SsKm
BTcyGPZgIpZBSvkjJCxqsk+MICxQe5JHViDJiijA9cpkRnbj4ZYEjZLoPzScw+Bd
p0sP0HYAfjghioAPBZTwqoB8SPnbowuX5SrikFcLM+kkVE1c092aIKRj1j69DTNU
4YDLF9mvUxHg1eGfFYopo1tQyWfSOKCGF/V/C9y9qfUysHJ+H28pf0C8Qe/XqBOQ
lS7Edv7yri7mrS9cST7qaJgYrr4nZpNXEm9X42ptfqWBysk6nuRtMCMr3SbDFWtr
70udpJD4kWcDq8JQVjrYKTN6JIe5UxEQDCPBvQ4UAIel7xcnhyhk0b4W6640rezU
PkCOMV509tg7I1fNPxho3Ih420XyzjUJRxLqD8AU+B6ROQxQJmcLi6puqOm7ESgQ
3eeQq5e5B9F4a05nZaPO/DfDIk7G9NQTPvNqJcu9kNK58WE1pUfl7ZA6OZctIcfs
3co7Dd4EzsuQsHvb7X6PHND0cAcaSQJ1/D1M5NLXAjfvE4aHBv15355B6TmsKZYT
Abxs+wB10Tg8UnfQmU1cPKKeLxsPtNb5R0fh9FKKFcWopRGQFwUg2qj5YCFocM0K
+7e9BjAKzwG9XNNf/0c+4rFHZTGbYXzvj9LmxKBLlGKenI7PMb70L5iQ576IFQZX
l8S1qwZaXI7tDxCquWEME3HmPMBRwy7I2og1/YZyHnrCJc8vz7X6lpbQkejFXFtE
+8WGvJHJFSzxGzfyo+IWumCEEPC1LmAlv8lZNCTu/8nXQhZD45XAJg5yAusuXk2d
BACevGNz7SX906vRDfJ/txooaSKJ8MpQdTxqmxfmQFdzH5GJA9M8v8Z/SBBiMv0M
/ICs+1nw9MqJcDUlZIwtnn3d1cE6AOxC8CUYQJ6KTqhzykvd25u7J6EwAQXaGXla
yB6N8YZ1kIfZBFIVWQ/zn6+k2SvN0CRf9ukuvPVuv609wWpGYfGgUpJeVq1Cc+ea
SvAKQG/1MdzGahQJmc9q3Vvh1m05h1J8/0w2nycHx6ZCQWy9VMsR6hiUwFumoZWq
fgYz9aE83PcFJtlImtMgzEAvnreEQYr1cO+OYIG5pO7DbzrqwI3X5DDJn/Ik2kmk
oOGbG6lG7l0ibUEIiHcRz8Zi+73oHzslsCiQzfUUGB7yqOzz4VRNKHEVTmVE/Iua
2/tVMTFM0Lyqtf4HzWTfqkRiaGxLnUv4idaWaYOBYtXpipzxtVSAtMjODetkpxKe
A4fXY9dVkXpaCrorA8IdJogR+eytLU2020PM/+7ml0KQ/e7ZAHMM6EHf9yPDRA2M
Ay5l28SQ4vAC4Um7vD26rkN5An9t+O+ygGbo+T2PU47+doNtnJeZXrf4PL/J7fo4
ST4CcvdgFjiqgjyz0WDzXuGigryoDA3v5Hm14ZUMHDQY2RQ3Ok/jopf5iF7nKLsF
W7Sub5WFggXteDaQ+NpbM6W2562CPKKIiQUUcNionseA5dtCLMh8cpo42wZwMDwR
HBLQu5RTwwAJmVCLp4JbKpXX964f8OreTdnbqWZt9BvJAjsGaMMYcSE8VvzEPbKj
YnlzZ6ESBZcZKcOXfP0ps4jIEVnG7923D1M7rlB5KCWntDJAfG3hYeHRjeD6cxGz
Xtiu8zKcgxHMYuh3Y3NdJWR6M4SAE1aCOBIYDef7lhbyMNGTtCN9Ldj2LTxCAN+E
4ZXmkZ5SVFPeCdg5GY5hFjQX+YqT1RU9QiLIBZZIisa+xyVvYZVC02Nr583IB5GE
kNxp1uH7L4E54PW++Pcs4qWsRO4NDt4sr8+oTVzbbtbJWgJBFQ6Kwqja4DA+yYN0
ucNvA2I+PLHjnL0eH4l1zMkL+DYanlJqXJX4iuVxVMgXuEVMQI1ByfotLX5IKWfk
7KUo8QftcLabnoWq2PyTUdeTuQmuTBiVGRmtgxjE/JyG67KxVa0yMuE3oElaLumV
BGE3gVGVxbIXjTz/cPN0UWj2c2pUb+mEaWIffAEcrjiUu5imjfIi8lTpuppPZfcm
Sa+5AclImxoAwqVvV29ZdAxh6u8QmNHOXeOQrCH2jUTxLVh5X3c7Zwx4FC0QG/hX
kkqptaZEMJwdc3xrEOH1t51qfr/xbep4QOJEjTjw0ql3GCCljZDzL9e5snsYjuq2
9zc3WbXTv0yQQYDWAqlhw0HJsCmd9hrO0wvWAziuhrNkmPA3XmmREfRwzKOHpMK7
08Y8iuZz6ZaypWNM50Kp6yeWPlr+hZCr/n6GxW/KLL8HsJ6lTd/4fGhO5tH+nnmH
QSIgnmXzDkz1k2/KIU11mQ==
`protect END_PROTECTED
