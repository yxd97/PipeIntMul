`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
shjNUYVuSMT8NtBMCoPOOgi6Hw4VealAXPO5a/Zwe1AyIlNZi7Rur5UxOthNlUi/
3oRof3gQn5ZXKqVWazQQCPF8pU1nkMCNNbJZj6lrjntGY8JyjRkXa5bMTuROHnk0
za5ndyt6aVKVxdpY9vMyvfBgaUkGox9nqf0S1T7Q76sjydeygsR7/9O7DX8TU99T
Mf3sVZIxRgGOh19CnnYmc56cluV+K9cgkAYnBdMgqxH4Rgi0W4KoEoVvmlPy2/+F
/xt4ock9k6LBihRaxM87D7fkYVQmer20pHSvI8uxFqzmYsB86owtu1L6jkAcSynz
v33p8/uGZvPzRm9akYhothQ46ZI6YoNrGJ0v+meCJ29iOooERUI1UVujMJ/VxH0T
fa2jR9almpJbYRXRnTqEIJX/JYtsV9eyQ7tJzQmasUYv7Ayt8FmQStPnSuMNvJnr
S7MmVx2HZ19KT5nbEBWZsm6KwQ+vsxNanKwYDegOI707mlzGy1BZxZ7p572Ps08i
BuvFii17qwHfXr8SDOZ9gAt+2x/KLR9N7P40IZDwb/7zEdLyAtGXZoRz70a43mQ9
RnS3mrf7+xhxWlvJeQe7t768874EXAgPhZjx5knpWOQtesuZz+hwQyyd5YbSjrjP
Sr9yTk9TGRlABS/e2vQurKyheS7phhDl7BDJScXZ9OCl93BMJ3HtQqhwXV3ppbhf
Hp3OuUPq6Dszz7y7z9yIlQDWox0fMOY6MDGcCCWHK67PHalO6nOR4GXM2eJxX8s5
Znz1lYKekMEkGJj38qY3dS3d9A5OAGuHz1Tl5VkyUcFRskAH6QneDMDHRWNeX1V9
sn2VtXvkYv7A7bWNQvbgFyRzZPssJNpjPRqx9ib/STs3TiD+PES/uFj9vSbTAJTf
iGaJwW9ORh4glPx0diOSkjdcP30zZjBVafUAiU/wF18ADBJUXwCJzV5IwuiHTLo6
0ae55Pz6fnxlnx/eusA/w4uYVmqeIXvgDFZzKu+3837lbVr6RXibhLaS/zXWnMRC
RlOIo/lDwARjCIVfQkdF71z4Rc9tQ1dpJ6W38F3E8pIRWa85g4jlLAu5TV+gmSD0
TDxM4GRiCTsQmu1yYQQiAw==
`protect END_PROTECTED
