`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qgpSsD956q5AFJ0F48ADR1DVyxzVIY3M55yZ7Ixi8t5nk4UQsw2eyfNNlfpakRmq
KNCsSBIQAx4NVugBnjDbPIctaabru5v3Vx5wrYOCZ8g0EmnBNoxPfxgRXc5BM0qm
hBvCUf84bq5m5q/Im4xPspbh35Z2QPFxrCknijryrBedOXA47qn2d0+vKEMDwbfG
hdxiTCr2LBvluwyPmCBDjekEla+/iqpGdBEaCkdL8Fqsk8HlUQDgK72TXUKknWFE
fMQ5d7FL4EauFIWeCWwtZu9DiPjuI7pcjaeowyZLAo0PvUXTPYpABDttESFFlWjQ
yTt+ntuIKIUcDE5uhr/K3bLOVd1fyls4ROPc8eKqfA1ixcFQF6utONc30PrlILkO
eLH9SRMaP97h11jVdftXDeyE7zXHS+LPtMv6U1Nunp/PTHoFGxe5mkRiJZJ8Wwl5
tijbqCO69Hv53njM64qtbQ5iNgJNCqO14ynwGEx6WNFh09bSLHSWd4V0lmdo6vU4
/JFuxfLl+VfD5p/UnXa+2b7cqaKyC3lhN0my0ldSorFHrk+4OYkLFwrBTSWZUYrq
`protect END_PROTECTED
