`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dW5hq7UufgSGfi1T4tP97d0I1XBGAQwwsDjcne6rNhrY3B95AQW0/twAM9KsG8aA
ANJbf3gs1CTV8EmddPU9IX83r141Z+/9e+aom8grt1d9tuOwUN93W6KBCyUdt3zc
rUxMs7UqvAWi88N6yUeLUG1yBAlWeDF2dewS9ZOm4wlxHQdJqwF9s5UOEXExjZ+V
pOzI6bvIFCpLliPuWJQqAhxPtH6Y9oJnC1CZFDOJxS+tEEZPybVonPOa98HFbTqY
lfTeCILTLsk7j0JJiWS1bYkzBfWCLqjfxRnWfGoJ18oFEHA+Oz9e9vLR+xxQ41La
yuvB3Gfj5oiC7jV7RaAFMg16GvxVlhF2VYruP0eDAY9qrq6smyg9h69F4PQxgtu+
lSAwmMq43eoXBu++/ZD+490reN+jaNdjsHY7pUb94i69wHiJSfVAqpPNNTPRJa0V
KH2OuPKeARdvTY4s41IW83T3Fxcz3HUHKP8Kug7Hgj6Y+T8d+QCpW7kuxNrAJR0j
Rqwyt/mXpuD9XFxsCHy7G1QNdGRAAUpMERsWYMlqLXK6Y2W/EMcScPmNrGWw29nh
T8mdpvXhlBhnYEfOlS6t1ihivPi+Cyllzm/gXwWlP9yc8V0R4NAP6vJJryC//Iwq
aeNZ1a9hZZynpwxYZwEP/U8mEhUSthPEqWSERBk9w4+gYJfMuFTkD+CktlAq7sgv
N0KxG7dKXE9jGqfrQui3/jwSSLwiSLwx6MJrD7rXAq0qcFn11n6fvfqlVw6zLv5w
zXa7kGGPDH65y9WmNO1koenFnNz1IPxVa8XJ63/cRnsB2LZjqOjbjuP+DRMtDqnO
ax/UfUt08tGMjgNMu3fE075/BYGxw3if1UJRRO4H2RjWkDVYuAVtjyJlEGxy2xN9
6J2zfTbIKmFOo8AP7QXwY1LCUv3Bt0T/xPIXzMt07v9K1K5GHIVn2GrVWfKB7NQU
ICdNJn/49k3/pUHH/Wnqui0CJB0qY3i6Zrmy1pomJT0=
`protect END_PROTECTED
