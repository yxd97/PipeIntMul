`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w/E3FMpmk3ggWrzPCpjKfQeFWnZSh94ixg3MX+6hr8yCjVRzAGctTjjDQX7C6R8V
d+hJjmsn/pyMcjmYZnHPD/I9Y6h94g6V3k0OO8TcjDaI6GR2Qti98FwS1T0Ez581
sv8OYX6cu5ND9COLqmZKVl1Z3QOS+WTMVMS0XPRcrhloPFS4Q9A7YuNru8zjCryF
vNOFfeHpgBbC7eH4CasWREBa8PYE+Fzf+Dwn41Gbt73M5MBA+epMfza9W1UrjUBn
bTXVspmWenrUxMoYpJsaxrz9oVi9S9Q/zAnC8jI625PFuuEsxGv3DgPSBPIwSD/a
DdLvZM36MVQmEbVO803cCNGea9x6B1JDn4TbD4+2p3xjCfxvlOhtcfZPPmrLAakW
`protect END_PROTECTED
