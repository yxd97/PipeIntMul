`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UGTvB4C17x8beGgdDxmJYSPw/L77xPAD2XniDWTF/oSDurls8DghV03buszrUN71
4QeebbYedUfygnRqtvF6s4IWtn/UFR3Mwto7yCzxt5vJ07LbW4s+xiiJVzMTAg68
LWbwz2IQxNEHPpHKsAkpkx5deR5coCfoQxDsf0y9krfBCuYgXK+RBlzgpqgaBzuo
2KzRtqg8YWch1Fn511Jf+YYTISwUJBdgS4uZiI1eqSNL/KiOzB0e4Z/eRTNjZ4Ti
J+eDnp04dDXkFKfhvauHrA88pX0Zt9TTViHz88JmTOW9KZI2/ZSjW76fOMPVz5jM
rHeQ5i0LCPuCFO9vlpLZWaNbkAtK3v/RZGUl1xfabsGHdvmvIJwF9qHJhvf6ZggR
RbrmbO71Ra+HCxAhmwjz9tMNYzrFXiibFymB23JwWq1RR8JfXMbzRarZRvm7Q/1L
mxz7B8YSKcfld1ZGNAsdGw==
`protect END_PROTECTED
