`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
djqK8kQ4OV2G2KpLWgDTD4icbN+WGmBCKQ6yFhQZcAgAKEbFxRQNcFuMVKfA7PWP
YA4SEckH20Uaz/F4OF/4l29jWNmxd0ClYRQSgehc3oQ9qQXEO7fMZfcmPKNBuBUj
am6zfcRDgxBlj0y15tjxfosgM5Ez9dxvK170BD/DFikJnrvE96uswkP2VGu9tiod
thPa+Hns6IEDHbLOpKKPLZuKUYQFkdbco6pOWVxXbN8SUkgsh8rWGe32n/tlni8a
y+j66mR/4+BwMSTSQF78n8hoEVTFvaOYa8rQYBq4wwZx/1BCL27bf+avyMX3hYtw
96yrKvFWzpeesMBSH/eurbMsEZf2+N/Wlh+1Cp0k6kPCWrHJbqggDdE4YQTbm8Bl
jTIuWv/He0Y/CkjhWLiYHKR9V31/CdEtRZYuxGJz/7KSU5jAfWuYxIOAx7ngv9LM
yr3d/5Xk2Dmezqu3qPOK9eOWIA47X7QBJx0NvduRGwNKk79gPmnFeQOi6+s2Cv70
42LErdWxNyBMaErMCkvEvzU3vSfZX93kj4hVnpYks/bkmcZB0kfuofGmNAb8+WU3
tbnNidq83304Wuiu0gN9x0HdCJ8eNRe808eh6cPjKYfNICdLvFzhskIhhJOLTo/2
wz5sBy4pOSOywlPEUuQecSPnNiTE/NSi8wQb1gJVzObyRxAyfdXba3WMXBdPf0b6
9G+5z+u4y7/WHFmA3DDuYjjbOf83+tx/zsAys6bNuhw/V1wbpuhZC1BoSVpo3erm
0QcmodjfxwGrb0YdANauQ8vTWaC71zPnFtrTst1q+pzgVjNl8SvlKZ4euUyuD3lC
IfLE8alc2+o0rZUNXiNYrgvPIHmjpbKGw0lUfO7FkjyPF6uFJwS4pFN0mhsSMiI9
d1PywR8uf4ITzej8C6SVe9aUJFisP2hEBUpSZV3so0mclLfj3reOnm0ul1HHFQK1
AUXnE3SzJo3njmZlPijWz0CoFuO7q0SsPzjil+eBqJzIzP4zRdkfiS6RjRm2XGyD
0Wz140BqAeph05eNnxOe3g/AyomQOZ10tAweYIzpSKDTEnEFwl1+VXdRU7O2p5xK
bho4ahTieQF3bgnTqOE/9GqysgplgE+kf15jLZ8VOdaGV89wr+coNOO34rlhbE0c
mrfUI7Q4xk/byVszXujYlP2wZJm8rR4Almh6ny5EVxPAyaN/sW1P17+Nd1PSnBMB
r52FRmThjt21f+ac/xViRWlr/d7RPLpNmaV9VXIy170Z2FWGG/TNEsvpCFWxVHYE
+5jpbPM/gRHr7Ol+lqJn8IiBLhglF3IbieSXZE0cjyziyuWGMu8Xt+DbUFjsX2Ty
8okLCfvfQG/KJWqgZGKdpsCprVaivKVJy+vdb+cyjc8RkqrZd8fdhT34hLgFdfWz
elv3yeXA31ERpLFtXddFUe6UBHJgpDXCwdFDxRZ+QpKB/6MyM9mrmnvt91F6stJA
D/oWQlBjrSXR7OpChCN53ZnxdgiSnPMuriS0I9WbHkRNpY4mBMIqYYhQQ7mOhz9Q
SESrWaLc4+ru/75llCR7hhFh6nA4XulfI0vPScLg/stKKoqvU2ptzwuhGZgFYF7h
d2R1XJ/JlSB0fCo70I6pPex+pLG1K9xBkLUYwf94hzM7l3nwJfGdGKjscptasHRE
lw23Czx7RHMGNlhAHP75ThT+aOMcqjq0JvGJuZVgu72aVJhoXpapbKdg5wrjUDXi
XYJ+ZMaiRRPutrkwHkc0Ab8dDm3p5Eoi7vaw8p3N5GbWe10NgTj36fuZ4hbLlzLF
i0VmlBcChGxsnZUkuK04fmtGcMlP8ftU7L0l76nluHYpiNM16BHtSuJm3vJdiG63
HNemghoZFMO6YlJsjVBPlIdmwHPwlUYspTchD1tpbRHo8685NpKBYQwrJyIVVYLm
9WAGU4cMc0QBgY51vc8gmV96m+rsjS9ms4dUuSCK982v/kuDiEy6mHNHmL/dyCYH
7nPjluELMe+bNdHGkDrZSDL8D+U9ZN+Kw+Tp2/5m2YE5WZJt3H0Oju26XpQq2yL6
fRFtZwXf4qQIXcCBwLszFcL3ZZ6yQOGGwmC4otXPPEqYH9lbjrDh8XuVZYUCIqvT
Gyj8eiaee3I0q2NlHUZhINYqEClkjeW5IKpkV7jJKpVaTTFwHq5twhIIKwcNEKUw
mUQIMHglPTGj9ycsM3BAW4SifeWOgZLpF+oUQuBulslo592QyKEOVTftCltfalmg
3XQk56bDxmYVPAfxOfwkVLK9rMbEQni4SvSZiJZ8PBmJ/KU+aY6O0AcIno2wwt+0
4JKISGmzaiMXaQ3BFokGPWyIU39Xn82Ors/RqHM060slJmH7ahbtL36NZ+a6AIC/
j8FUQkU3qod3AHWYuyCmDUiw6A7pcCWS2Gj8K64GzyHp9LS7BY39m1t1VTOqoxOU
/P9n2nirThcWjpGsjpJ/pQ==
`protect END_PROTECTED
