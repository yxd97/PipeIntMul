`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZbNNnx2H0fqx8IHMBs309ouDt11p2/IjHERgWQFl+sPfQpwEvcyWA0ayJSRhUq1r
kjAmC74sP5Wg3/eCkDaYIyCF3aL+u4GIfxiSD789AEmYIal4O+hLOGQmBKq7pRwc
0mr/0KMyLBmSyRpMkW2XkqE+QaFMA9wF/CYxcvFRv5rr4Y2N4fSVPUH6wsJXvSs2
q3TB95oFKDVOCxb63qKkxWeJmfPuJoJuRWiCAFO2w3ZjTovTIJnbyOtIzBEibEGj
0GR/AHhPtoAL27la7/zIbyXQTWeqtMi+LiN0kBS4JD/sncovuZXrKT4+m9d2l5vZ
aqmhk4BiHdXqYYjZvNIGEI811lI2IUh3mhM08KbBmOPHCi1S8oqp11+t+l8fNkvW
o91rbYUyn30COI95FvMIWw==
`protect END_PROTECTED
