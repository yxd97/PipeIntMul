`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
admf+QHOeXRqOf3vGRdeFvpbrMIhzZ5J0gLpNNs/r4UnP63/D+e1z6X8LDtvH8ys
snL0Lz3CvxdaplGUerN9oAp9ZUEz5ks+euJkVgMRMAXIvJyQ6/1uhRUkzWvt3tmG
GLE7AqD4AUQb+/ToIdQ1TD3KZVKExj6o/egehRjj79rtIwemH/+0kuV6sy09jNvz
Xnvb4B9ZA6D5kNb+BA7PB4XhTo0IJ+YTrahCjQLg94GqElCuZEJp917KRaA3nLFs
NNwFLiL9U8xaPpk7QwmVwIS0n4DT9o+1wuKsV0qBcNR6bHuKRHQJXTvIA6epVRRk
BrhW0RXWcxV25fLxWc9xoSI1Oz/hkYlcxbHiBq92LNcXDB5aoyzb7yJ6WBhTJEFT
Rn+FwIUcbU1XxmJKyzxIt1W38EwIjMOQ62dCbX4s5nHJoyOme1YUTVNc/KBv9Z+r
ezhFCEq05SQLBw1HkBOP1k2Z9+0dB/VjiRr6Bh2XXbr48qxsayJXhL/1fMo7zEc/
wbFwR/CwA7QM+tBMgVuaftP2s/vNNs44DFE6f2+77DvigiqCQaS7GHUfAyXHhMK+
Hwq5Bl1/ftkbqFBFj4dXOD/PaYQt07zYVyNMPcG8oYHl0ZFOojf7U25wF8ZnSisW
LLWozm2Pm+g+eNPh1fvODT1qHbOUoDfvHSUn6FmDD4FCQRaqprJEy0xRht+TeoWZ
q8TJL/ZMiD0UcI7pYvYLEIyf0lpO6dalseeJP88JdOYLSo9eaiAxAO22TpJay/Pm
dBJpjwTii0APFzDHQkI9jiSsWzt9bxr6Ld2PQDkY5icarxvLADYMOjRaGc2oy6Nt
9+Qqfb/kKvfCAKheeUEUiCqCtZ5q36PYJiTuy52iI2/GGwKVmaheGqwmqz7+gvfl
VW3mrYgJvZ+A47o4pyI7K2dzt6hXxSY4de9eizfOAGIhX0JrYVBlAOBUhvKwP5bu
f7bcHSXqIhDFk1hI4m9oisymeaNgyJ1AwlAgqzQueV+E60lWmg15CAHJ3aO3Scsu
T+USkKnOVhXWGWu9HFWbwLU/E3Q8P9mVGhK6F/Jn0DBCavXgMJLaMAbCuIBz801y
j5EM1NBS55cXIzJD8Fr9rFdjaRN1rz1M8Zs29r3Db84aDvzLTuG8HDwYvl4E3gvW
dGrvpJT8GGzXM2dwmUQT3OqsD/DoeGzYa9pF5H8Xu9fCdLXn31F+9eaDxfObG+ht
flCbv+kZLfPmp5v2KUAFAKNjA8vkp8sBjLlGYLSErqnS3UruvRdFaMVLunCvloR/
GcadNUoTcStVK1H+jAfRrFYIMkfOKgKoKqoRTnxCeG5oscRew5Q4Su/OcwCvrjMF
OSM5r38lTdYrf4m6xpLdyDzbTb1rojdp1gCUWUZoWzrpsnsEPi3XKZiDhX07c8zi
xCWLo1IfVuqd2/EQBXt5oS4saw/NiW/IJ7uVHSOCsC78hfoaZ326toLHOs/yQcPQ
YcxUqZrP07qg0Ygq+B83PFfhMEkQHBqaT+I3BaSYYd4z6TNJ5bLXjNbmZxcekRjr
lV/0kAEm6VfxWTcgcNqQdKZNAWA1li6p+fofJct+L6y8HOT9o6c+wykkGZVJ5Ai/
`protect END_PROTECTED
