`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wr0xvY9uDG8YeRdSL4LaSkirHzaTbTG0/cA4Yo1nh02u0hGIA5PCwdbD4NPkM0wa
cWWCDn13681MPF8C6y0KDNMZQ+jlzlIdq6dpAXOrEwudqBIzj6vtYAW+wA8a6XiP
SeBYGTzQXb8E1jAIOpRjxAQsGbFk4cddLb4i501huezCYD+T96ocxzWhaJH0eJzr
gxCjTnKIzsDANJW3Jvva8fggpzfmVnZusgZ4VE3fel8n/oadvmYyv5LC6uUz9tHp
d8HB3C08Uqtrx5GeAe19xsxsxEy1UwA60TfIU50A/6cbZ4aX8SNMaGFr7pIJCddP
dGLyEjtxpKYmQUtnIN6c717KuQlbk4Pax3MI6vzD1KQbJQS20KQOrb+EJ25ebigx
QlnEZHvOfiASM3R3IvnB8DBCwbl8eulzzHBEiUr+SnyaI1GOuGZP3wCW0U0Ekx2x
UYuZTPIVmsq+prCsMsjUaLv1dIIiMJq+F2AnAS2dIFMGa9SirgJPXp21ureKD3c5
fB+MdzDOg24V5OeIJISRbaciv+hLhtKrmyTmBk0haECko5GkM0Sr6d+TrePd/+68
bkEYbAs0v2MclPz3q2Dd0042EyZQx+5PQX+pSLJkYfDO4ihyjYIJFGU/Xq0SBhiQ
VVFpPkf0Oq1unfb/P0Rzzhg0iW3DR0yBvlHO/pQo7uzKx6bp8ZI6TVXuohDk6jsD
kvXMWexDPD8huYaWaboCBipFgrjQwcvpFwfkre9+NiLKjokVYoRUP9tCoTa+/+Ra
`protect END_PROTECTED
