`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p770E3sbeq768aCQoOK2wTq7sIUddhrvB9WHaLNcy/FZ0n4ifdYOMx3axcnWMGBe
nIn3j5e6GtwLjIHy/cEvlP6EEF0KVE4o3SLcISp2IUA0U2vnkvibBnBGPjvBbVZ9
Py8Xsv3tejnWFbfHpUcV76BNk4zGjzdYcmYTRP/udiYVjImSZqtu/EbRawhx7G/Y
oE3vA02uAVLIzmwU4H19ujldXCDdk4zZ1vIm2PMNWlsIaXaPsrS3Izk2YRU7Xnvx
ANjDbzc6IHpgcPlDbO+B+FWUMpFC1L/a6eBVdjXGTthHmHYGf7y3arSVUBGDT03+
454+6dBpSVcZBHrOYlf9N6D+5A+4asToBfFxqM4E7B30Hfp+NP/sKHVx06gOA3fY
qQwBh6ubjgsU/XJNp5OoOXQKxGksj0Sy8dWVrkFO4+b2eO6for3CyVbN9h9NdCII
wHy6aw24Dp9jS7sZFZnX57GWYeuQz8HvPR2o76QCYXipKW2w5dHDfBUTpol0ZqaI
MA+GC2r5uIldcW9qAx6lgVI27fSvcO0enz4RFT6ZOWeEJnlcD1/sV/dXZ8Ub3LCS
OFqCyVgRymbU7yAWAe0sK6KhnifbffLJh0X6W0cDVBQ=
`protect END_PROTECTED
