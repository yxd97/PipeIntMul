`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rAq7jyFKASKQlBJ0ptedTuYhrBLot4DGznSf703al/xV+cZVtCsTsz868QX7BrS+
D68ecCQPcyL7/2/aSn6Ak7+U4gQP89MnJrn3Y/FSAIkfeWdC3Yq0dYVmYIGBleTZ
nbi+irrLCIjR3z+8amJQSNdz0lof32Tr0m3CyTRIVmUzvHm1v5mklcX/O1yqu4bL
lD3SOaqdWljjq01K6X4Em9l7aOH9Y6cq7VQAGR2/Rlcy1nB9QEYOd5jXLm5OjM9I
xFcF1VFhu81fbFDtB8q549oMGojVnzdECnPG76X0vF9idQ6j6eaLOUqXdWeBNhjX
lo7LIXBQee1PmEaegxtFTF5GEOqVIRNRf1y4cmXHnjr6DF185Q1494FoWbSxvud7
Fn1mtVSLnDIB5f4ypBuEIn80KbsD81hlnTkTuawvTEcZ/RFqNF0DhE/YrMvaGFlN
`protect END_PROTECTED
