`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZDTbgrE6zfRJgb1dZmshsHSlGV9LGtEte3aQs2RjBj3gvp/hcIlju8Ep3TUzpyBC
Ruq6xPpoJxKSfE/Li11ZYr7Hhoi5xg07eq8PKX+9NdJvw3ZkeDjqzfQSyKI+F4Ny
lRoWkbx0V3LJfZIFNrAwRpTXF2zJHz7BTgl9oFsBLVJO359lxDpgY1a0nFl1717v
GJwrXEE7JiVLktT0LHmaYhBiz7wL57BwXQeSkY39vtqXGQ3nmwzDbHmVVXS2Gn6C
tzeL7ozEoPVGZIzA0tCWGWNQ8aJ5cICSUG3dGk0DUyNwJogUa1vMKd5K3c075vpt
sunvjK3YY8ZvdSEOxbSAeuySYYN/LT0wPySxSTUPmgxaYB+pgOi2XLYsJ5rllgXn
cAlUAQ+0+Cae1VYu/ZSkxySxo+GEQjhcTuxseJp/nI1D9Yoaag7QuzORl2+7gU/t
06p5GV29A9GHuBDkT9E9pPcpY4M8Grre9RyErowgV1YsYdwSc0OeztvjOgUKduUz
awf7BRj/IDx41Xq3rLzzIhnkQwTEJAdLRzy1z9Xs/rvBtKO8oOq3760tiYBVRA90
mOYplOsxRxV31SLdSOknuqYmwSxLQysnKQzeCijkjV4cTiYtOOBYxy+SaesXMD/J
tXuvmLcQn7DxB+5mOLvNxcj3fnSOT9eNe/J/vzgcq+585whc6TRTd4es37v/nQCL
SoY+De0uMl/IJp6fh7EzUJ31YmyfeeRLKdPj/D1JdFNlsW3VY/U4gZNJ64aYF4D/
SARzhD+eNAJTPiaQipLRVN6vCvyPHhoHQI+Zm9QxC+z1LVr5t/PxrIKdxffrBnYy
7zFRnrlAGOLENP1T6vXRo9Eh5sw3FWExzTYaSL254sA0XjFFO6atq+8lMdNk5Ife
Q9csao35oxrTN0B2uo6T52ezV4q1mpyBhIImC+w7jfnSRgsDAWK2WARKaLGj3XZ4
D4+BGVJ+Z145IS1MVf1sIYfs5VLiEXHF27Nk0gcJtdM=
`protect END_PROTECTED
