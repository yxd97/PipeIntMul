`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jpvN63vamu4bx9lJ10NwgQrZppIs72FK0EHZV0ewsnCCN1PyQVdx/D7761WyMy9M
dGFN7wvj7FNMXbkZIaTaTm70IoI8mn9341jGDfZbXDrPDeCwdcz3REIPI6DCy/DK
hUMBg+Aox30mYJc5Z0ZsudixBrAGqd+CreJM+gOdMe5lO7jxuENhz7Rs8MaieE14
lDE3iMvcHO/qkhtJ5D+IbJDAp90M2clffcocWcDNtQtpL9PvjCPdbrJc9xzefDpM
CLDsPA3/GwjaI8jJtuRGp8gm8EKrfiC4fJK/FaK4vRttyGOOL5m3EKQq2TvVpmpu
wgazbP4S7OicuEei8GYh6amLyUgXTkEkWV5MEajlPGHjkfb1zhJ+ZDxYmVasC6LX
6h/ddEheyA+5JZZMdxEl3F1nvEvWPn9550xdwiy3uwuHbVfTK2bpdtg3K4Rk+PmD
xWCNW/8zOvOpH1N5IaAbGOZH+ZnuiAelP6pjFRtEER9XSa+4TXmOIox+BlTvDPUX
r75axxcLI57miY1vvfavzg7S/vrmo8X9evM8xigWi4oYUFezK/T3FREvkSS1Q2L4
+LlaaZv7QzuBWQyvaB+SpyaPJM/tNvQMu0dGyYPnptt9GG4R5rWEvk/fjX8sNiV9
EOqtYL3rW85mbCCQuq9CtglJ7wj85hVE26vRzGVAzu+vgIScnZ+1NGKDLWkx2tBP
I1eQUpZoC+74qiqYxPU+fh05DYDUsDkfKETb1WSfvcKdAR8tzr295AArCXNnlS4S
jFW+qovEf6AiNHIEQwYaV8yFVYjvW0oqBKnguA0Uok6mTn6v/8N9gHC7Lj4p/D4r
eziu9M2NNxwmjxMMuqy0UMW+TOS9RW+TflWHhNCoUZJ9y5L8OA++PY8P9+Tu60Cc
pEaQcNWwfQuG23mEQeLr8oMO60RQz2PzxqgEPRfqrpKZQA4m9D+ZLIQ9RBW25KFc
N0iSlKFuSYYx9JXV3zmun/1fTih90ycRan24ejSS4C3+erNop1ErwBtaY0a0zb/U
gVlNj+Qk/MFWKj9f/JLN0gk6ScrxBGJlEy3gLERucfEx9/8rK02SVJtdQPRc/Bor
Oc0TdrVOiXwJKZ6im7IBAw3ppu/L6o0rJqVtyxBfxnIfokH9+goaAW4aL4Y0dN0o
5fqCUbYnBLQV/r9pAkFTJHbpsC/MeTNty9dKVhxX1CTLTyk132+TbCHYHOmum3rV
mb5v64KnYusqDSQUyGJAjOPLuaEN3A9S/7639uaRIG9xyPyYRylukKPFbYSN70iy
4XXGRn2T8JbpAJMfD0oWBEM9qtM0WtkzuWOhiZbZHQ/DC2JImVm17SrEiscq0GBf
RTMe4JBUKKkGkTR5SMAOXWsLz54LjL2PhxYf6YMpSDdmA4FFdJWKVsRej7z0z7VP
Juu2DLZKckyIh1JRxcWgs/8/t9i1PT1DTOzSqaVKmUvs27URdIHQbE2231tPoxf6
eUBfNvGk1OsOBY27olyhcQr1jUiMQryUNPfIoRU39oTq5GcyicoYs7BFZu1xLtK1
usPVlMYVgL6yddJ+r5EwCVgruG8nzBIZd6ru6XwH59HxaW3BFXqITVqp5HpAYj5R
eTo3AeRE6v7QI+HQEIwp9LPEQ0TYvPiAbdhBuw/UBS6AB9x/3qi/oEw4U3FULRc2
aWiQ8x5zahTTB4pId65sJMHoDOJDvOFvCy5F5cy5iI4UgK1FFASEzT1eNZAEE+Tf
gEsrNjVRZDy5mMI3M29OghGpD6GGMao9NnVQYJkq8NmYggG7pG7qqP1kFEoVDCYJ
QnNKUf7FZiCmY1HFKuqB7id5Ja2e519lgQcWZz4TxpnDEGVoQbMumd0P+TUR+ejE
YogsLo9g9qx9gM3rQm6Qj5ykysNkcAwtF59ghj4QbxGITCn4hG6L7V23468K/VqC
phH5ApBBhTr41X1LQX5BkvFi0Vew5m8zWb8cfrFqvwJr9OFO9lGLW8gzstl5Kv7x
tczfKpCKA2dXaQxGUi70POkhcP7bkKCnfEKJOtpSnXZ5yUeplGEOVLopZbf/F8MR
d56goo7RMLpQbwpibG5fLH1GITA2UeM83oBF8Vhw9NI/qAtmL7gsLMvLK8ZMGlfR
9Te7tOe9JGQdZ65zfYRVEwb8AsigdpDMEt/vl71I87xO4rriDc0Xn0N9xsiEHHc5
NOkLxRATVcBM/7u8T4sX4QGwkh7iXUrsTkRRiUBESMrQi93qoPcINnTHdgacgf+k
5sLMIPzGmnCnrCejyPzzIDe8S10TZPh4G49BMIJ7tmGwa2yQwl6L7ODVl25c+dk4
3xkne27wX7evUmFbYt+AOLGJ8f1lfgdt8V9NjBQ+gbKUKL4UCJwOtM/636YgPx0t
eLD3uVz6ZRuyst20UFaCcr/A5kd/eMHhgG+SszYBluzRSHl/VTdFnGPyjHhMs+eQ
O1BM7WtGPIyaIssglbwES1EuQKsoWCuoDjNAR2rhKkArV2DcmvQBHCZLQheDqTDx
GUb1EhbglM5jPyeUdWvK58pm1S+UvqIGgqPqpZIdyYu4gl9XCZSFEUuC+6m+4lMu
OwvifilpAqBApthBmBHLw4z7wh6SVCI4djn+kDG++PAmp2aMfOln99IC+k1IhbXi
PSVWLmHDCtD4ZlH9wIy/Gsh4uWdt4iknOOwbxfZR+OdBQhSx/lvvv3FzVhvh14J5
/Cd7zuNLcaZS/OvQwRRuueCN5wSM1vhMjulxUxV0eCnLPfbcUd/0aACzKCihnW0R
0QXAJUQRgU7jjdTusLni6gqsGHIJcO2Kcurb3+BsnUKNPERr38KR+DjeZP3KF9vS
2Ab9xhGsFikd36VW4lGQvEX0Uk/Q163i8ywHX4lFpBkK/Z3RoiYzBrZUQhn3BbvN
/3ghMmxJ+xHlXplslaNY/7xAbhyk6oeRLC1nILVxKWB6mo5KOUaSfBR8phV7H/L7
0dTxtEpkgz86UDKQXQg/oBPlxXO+ie0DF71MDCslw785gAWKxdejeEQOYbfEHeyk
xZQfkiz3m1S6CyVioIfB1fi29QouffaOc2Uq7JC23v38f0mD32H82Pry52yryfqN
VQRpGdxMkrtDnDQsQz66mBHLQ1E6k0tJFZv+5GR/5A1SVqJs815DlCtuh5drOz/S
SQfDtqgL6vrsM2h6PN6EQafuA4WMeyvn0pt6yRFye4wZoULuodk18J0qVU9xWsdx
FC8JO03kC4BEnTMxrCt/bhAsV1h/84sZ1zanOxNL7mDH5bNM9sFM2L3bxPKwXHQl
1D4Jex/2Hwy75choELYwMQ4xSiausY6befCwmiOcMPcQeuFtOIwOfecZNmXEt60c
eNGRbwbcdL3n/kjRAzZ5zD1hMF0C+4pNFatcz3EqWMPiJV9rjCNzDubQWD1+C+WF
WDHbCgb+00ECgcTnD48gf+1sjPCZrddoUC+DK0fjMirEeBH1rieQZ+MNCMZSoMZ8
uTK1R8Dn0alk4tawi/kZV7pXh6UzkSvcJIIMwRn2UR9RiHgzgtI6RZuxmWr81h4m
sg+rODYTAgK73LtodjzfaCMMhN2e5jsHLYkZMr28Zo8V2Xh2CaEYPwb+5vJCduyV
xAWCsL4kOEjCd8hEJEfp7u+xaqmiirW7/8cHT5V1agVC8r/0V8pzQZ1TyL+un4EJ
DLGO9TuAy2HxB5n+ATKVgNsXgidKGyL2mWUNCB43/unlOgR1Ummtlft9O2BD2eAO
/yJc146wq4UR+LJi2jvyEq3xvvfG2gPkuOujWJ1kCZl15fYSCP0xitgsXxeP7Qbk
vcOfGWri1ta8Y/XnsWpGcT4N0totNEppJYkpLU8VcqLENKrJWsq19J41ZSDIJKig
l9vhaD8XhR1IzFJOm+HrQjtom30VwtOwOjli07I0NPPS6WCGVZLkW0G25p6xAv28
ngjvnJ3k+5sGZjtdmm4CoIKS8aUhwrU5UEVamMVnFas++2vBHZzjdFZMCVsbqFXr
n2yqab18Z8s924VJ8ogIxambt5VitHLm60NKTuoEf6M4pXvOkyIFSpqOVuOO/wy+
ALQ0nmY1heKTuf9o6O8NtxhmzG1BxUnpECL87WHAkmL5Y1R/TOPrrdwHxjOss1ip
ktUfmVRJMjBQXnaxxV3TQEbkFZ1a7Qd3uYAAtKMhGxTz3GtTkSZM5Oe6+GZX6l6v
`protect END_PROTECTED
