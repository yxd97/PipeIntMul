`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iFGKLQ134k/B9xcoXCC8mx1LoKoxUrhXXyD2GwiXohnw0R92AYiT4w2nbkF5zj1m
rXp9d47CNTvQqh5x0MoNY6jAqkKIJqaR/2uFiI6fZ7u2+/aXZD8UDOcBdYvX3L/i
oapOAmvO4EMiafsgFKvzW5i3oW/f+XxmRzGfQsQPk/lLwPzXhQIxcOeiwW8fPYaS
Qc5jRL2pY/D23tosZ7JL7xa4P1XgDZpt1N4vk2vaN/mmrk+o90HnvPyvsduMhM0L
lVtQdYmp1v66sC3h0+76SNDdaecKF4mQAHsu5dHEMLH4UHZKSl6GMLdsl2mnZABS
KypM8sgjHkLBM8F2JERhD8cjQLQ9nnLmVptD3RxZWXrbevKTSGUCL+EXPHlbqvG1
YAXHTDXhqc0AKZhS6UD22YeFm2g8ePhaQYhFQmWCNGwioBaExW0pjrO3dswY6LNb
lRnt6gp6kfJdZmXoXIQsyjVtEyuTHZUldHmgLF9LNT5hz9tky6sV2/DfHEBvinkz
0LL+CdDtkZjtUiCIXPsDjb+auiUta1ornF3MDfjFCMmqi+lblDJJivTL7OZ3GGzG
O4jO4NiGbSIxAL/jnA3oJWEKeeHAUq2vJlyxkSTBfFZp/nkOzc2luBs2g2xauYWQ
tuRe2yCWfO7veMGrumxtRZWaAUCFmHrksGWthqJefk0mCSqlN9CMYxoB/8UFVd/0
sm+1gYs5eNGY5MH5sJ15B1Z9ZfIFI2uumpAab7SlfAZKhshV591Ebt9oguH8pm5c
GH+ZKYSPrCaf7a6Phu6oLlz8U10uBBFHwfi2Wje2iBid/dnCoKd84/WXt9VFA7OU
e3hbea6GNE4WZMk+8iI+hA==
`protect END_PROTECTED
