`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kf0Lzh6XLGvvqTkPxBCPnsz89vNEerMM3nrQ0JGJePeMXq5Dh0b391P+j0Y68yXA
ah6lm/EaNaJsWG62U9mOLjahj0hCLhWJUXT9g5FZTcntUa/Xm7jWaaymjW7N91kQ
WQ/ez1sqPyr2VbUo/1YAmhlwD2wLxWNB55BM+I7tbe2aN6Q0/8y2GfxbhwRhjg5Z
6z4CuSjlQpKHMC5lfBmDuSozNb3hNSto5hD/vTo4DBLVGMwcVxoBMcs3ME2JjLAq
kT+Gx/388MJbWG50xyCFH5nUYYg0ndTWn3lytewj1qG0EE93xajSV3MPPTeq/XlZ
veC3FaWyCyfFgjPk0N0rlxfsLwEJ2DzC3c8ScNk8twRe6Bz3+/Jmdel5bovda/Zi
jfFkX4XdD2iU+U+EP/Vingmt2b42bpVWvxAnAZP1UNu2EnH/4jtwEILWVNch/Euv
OPUJA7CY/mSL8oGyJ9zENig8ztOv/Xd49y824UC/ShWcFRO0m9JJWm04AQlU8x0D
lzriqCJGPxSEYpqnV/VOI40wxbhDwJioDD7qfEdx+rkeesgNDh2ez7rlWWlSArXN
1UStdAuwotAskXUrVf1mrCbR40EbW87ahFoFnXrxfSs=
`protect END_PROTECTED
