`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
akR/5/n45sSVdfHF3J5CPhuGCNKYfFZAy4hauXICaLL1SEKAg84RkLcACyV2pAmQ
pWfMkATcn5vl9zxD8sj202pBPW1Q6vHhq0DDKyaa+24imuUy7iLlOOV2CF4b6tt3
l8ajUxTGjGsAO2/Vkj8hxiqYYfoP/wKZ+X64nuZUzDZYqghilf1flW0ovJ+HUO33
ZZwNLWjSx+BlKlrfu686CmMEq838qa0xQQrGjAAp5IVmUNb4iaY5oXQf128VQMET
a2xtcQlRQ4ogoIbuj/3f32VGMcJL3BWWt6/LnJ/yvEx1P31M/C/nB1QdV4mjBPJ/
d8CXsa8HnoJhUpuV6qMOgFpS+9vahPf21EvpIzmq7+xhbwWpg/U35OL1Qtk+9f2M
QL/gplKFlvigOpcTAj9HAQD43BjOg+H7B9Iw8qfLSSq0EDeqMrHdvk+OXlKyx3YO
BljtYRwkSC/nIehqivl4xwEN1I3DCiJqpWHuzj4Vxq75mPqqkg99eDi7w0wa/e+y
0oKH0t9IA0DvAeE0EarKArGMP6V+JmobxQ/lHEVJ0vhufU+eHhPPZSPxjudNF6EZ
e/st0pyDRiK/GesS5X5oChbJNR4vv1r4/MpesTpwqQqRzynmAM+D7j3rKm6b8DVE
CpKPrHzoG8pHahuOVksTyZ4tko5cZPGy0t7wyHZR/fQT4f8OQ1C5cswB85HpqTRG
PHJ/nQQOn8qFMHIdSslxMJTHhjzL+qt8igt4LVz0GvsjQPm3xmeBJ3l+IC7/dRGS
lPUI7s7mYKgkJXkElRgUBrnjL6ISkLyW1m6uZ4+3pryvpWA/SE0pupVdjVZHPO6P
flU+9jmFaZ0PVs7IEJTcT/BmTlbxTDislZdamjPLrqTc+btbZ76ZM/du4z+llK0m
OfwAP9BBprVmp0IKwIcyFt8oUAGUuW7AEQYUf5TFJqVAXso9swz1lRq2atAjOlqh
LJxPKAkoUYgFt+PxOg3L5bdA2GJDk+EsUXnfsdM4WKuFR8aMPJdE0zMiIuM4gtSG
uQsrpi2cCuLjnecQWbOPT7c1OJAoxU9Rrq0qLf93i785jPbjfCmI1/1S2Sgr1922
Bfs1dkpM3V74uqGJiZ973UCl+F4ZcbXtmpY+cfms0TjoGaf1660sjaYpT/hJS5z3
oPStM74YUpz0N6nFLPFf55Kb05YsJ7bLSPGv8hBfWW9EkhSzjyk2KWpeKJWpr/x7
soeNrwnZC/zqoB8UhKs3Lp4VsMv0f0Rze3plda4NPa9BttzN20MS+jk2hFuRj7Qe
5AhRqTp+IBi99Drwo5+yDF/d/wZvCUg6DqlG5P0duvWAoyvqOXISUnP95M3KXyIz
IV9UDLbdr65ReN6jtjNylpVLC1xqYjQkiEqQJZKg9cwm3iqAh/U3OMIR23Cvfdwh
hnIyGbXi1wmTi99QBJJIY81LnnpIVh7aCGooiI6rEI9EsU0Fkzg7HN7pULpTwzdM
t6pNTsFMGfme5ozGOnBiBY+SrEAE405GtsF1lDR9WcBc8SRRSfIOu/4p9/jQ/VNb
1Cq/BBwj5tOg10ftcqUiZ63geUSKh9c4hY2fNfZVKI+uQpKiGpS7XLquQZ+K0RAW
1+PJnrcfJn6XJWD8xCffGuPxteub3m49OHWAEnCN708/1Kar1F4vZVGT0dU5/YD9
f2CW3LtwUfYgozAEN1U5e9N4CuKOi8tHnGStt5opdyDDLKV1RZrclV7Nw+bdQAf/
5TOOooI6+JjBwPj5yD3mc8L9sejRJi3OIzfzgCEq4+jaMcymAuE9WPs5sAioGahu
rPy0hk+hd3UXiaTrJCw8r5uaFjS5b7H0blEFgxDMJeAv7ES/xCuMNcBC+BxDc9Uk
JaT1RVM1BavQwZbAi8Q9fBBlZXWsItaCQUCg6bJ49aJxYV1pkMo8SQyJbOXBky/D
3gKjoaDotsWgffI8I1hZW254VxMMGE+CxvIOoYA895KsszbJLDfyquHQgJUuMPvG
nSwFEMyz5T8bW8lnrlpf7iTjvjqXi5jMqcd9v02kVd5WUvnt7xN5b6TCkdKFyFPK
luX91QCGC90IDYUg6/Jcn4lsaKHyiRlehgGgqFBsHjjTddIzqbbCCNDnNqB/Bkz3
AoEcdXAJZ2mYpnVZsqx5w1KhyOUBnral9D13/QXZDhhhEqb0acp/Hfie0psuZX9d
lSWOXD5r1BCcCNmXjt5xlG4q63ui1pRu3bV8tKSLq37v23OIlr0HFdVEaay25q3O
351HY3RmYrIU4U4xVwg3+fC6WmSj+YrB6fx8VffqLAXMY51wLVBovYpexn3rWToP
6cNmT5b5RLwva1eHebSgl0C2e3Ht0UdRBEIvEDCRjs6QOlZslUqt1ZYaExDMf4gl
0g+51ab2LvCCDltoxyqhnBuCXVGBelTYR0Smr8+qOKl2Ug8CcKsSWFl2HTgWV8OE
lKoyMGWlhVAskolFn/sTwXN7Ehd332oi/2dNnOsnvw6CGOIf+eBZcnFHEUYkhQKw
qyRZ3ZwTQcTIY3TCLQUkyWcq1oUJe5807Piv9K5DNy+aYFeKbO/lIw9Jrx3GUQBW
b2fyroFMjlWxMy8vK+BTEIadrcUEhlCnzkh6ctJhXYHb4weIvAyPRUziagwdatXU
+bIdLJLYy7ygamkDQsPfjCG/arC8V/eD+7ZZNzsvr+QOqcy6siMg/JlJuinQ9kQM
N/ZsfvT2K/SxzdHOnSR/UhvrZuZ83KVE3JnFPQd/jRrmoQvvmjKk3MiiD9Dh0UQ4
DgAXtQprpr0JHs7A43l8X77xkhqXYBjppjgwbqkNXzR6bCUAESeOPBHpCEGdZX1t
8vQq/aYGvQ0mfCySLpmyXKKQg6Zfo8gTeLCnRf5ykFrj4rxs+EC0/B+VvlYMbgXB
cWzIMNU9p1nSW75laSAgMn/b9isXzsBap/VALv1KAzo9HFdOBYziOV2El+Smt0MM
ceRqEcq1bG6JJteI6DL6T9aV7Zm9o4AFxa+oLO2W0UgIIfjSLkl5U/0K5fA9GKL/
19a3l86Wz8ACNdI7LW/5a8P9Mm7cz8YECnRDU6ML4LKopM6O5zyiAdfVEoGAMZRc
FWizgpMZPudWytUrvmAzk/IKtvVXRTPyIaxMBfdYD90l6rcGEx8qydEX52vdCGoK
QySHLyBsunIhubBtE6gLKA9ondx50wuTLw7embkdYLFa8vc5sue74A8MBn4MtEp1
ra46EZsY/FhtwcKszdABjbuupKrs/yfhVT0ZiZjBbc4EbaeDhMW2suCkoPOeaNUQ
59OJBuw9MIwO++nM2A1+GpEWkIx9YY+0fNWlxU+tm1szeFZkaR5a0TVCoQ1gC1Ad
RfmUGBudMc/C5XCp9bzKWEzJ6414rayWmdsK3d4J330=
`protect END_PROTECTED
