`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Bb8/HzkjvlboDxXh+T+wTwYl+2W3xbZBSGStozzKKAxnR2mz4q3Z3A0HEDR0uBIP
UiDqAC/2WGKPHiljB1zAkLMx4JyR3Uo0oQ/heyqLKVgH/5I6QR2BheUcCPB2W7mz
wQoILfKXAJDwS4tetm+kk/IEb+DjHp897vewJd2IKgiclYTbzKibu4HlIxQ8wT95
TuyrEajqYUHyiECFiDH5O+Fg8zPbOCD82WhDieA7yf40opBm0zKhJdbUthehh9W6
`protect END_PROTECTED
