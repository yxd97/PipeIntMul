`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
aFm41EK9cyVQGYaSbujoVjmYlUZJTa6p7NASnqDzNPwnCZDdNAFT31Gyloqw4/DK
PHjNfNDlcEcSCpoKEp7ZIobY/E3+I3bwuL5b8OHfYtEJfWGO5UEBrfW1YaX0c5Ts
cgdLy0FQBrHEW5OKWrQ0BJ8X8WYpa4yeWJqdKunt6545w9AM17SP0X22jqEmZt+o
/MtZ3kkhIgrWBXLGdKILMf+Bq0nJgzMyj0hjpeDYIpS07fe/Y5ea8467aALJeD5s
QMBb0KlWmGDIPf7Y9Yd8nF2w9dEXnpTmwNI06RGM4slnkGGIAu/OKHVye2fcVeTs
JaJmOsH4FR9ztlm2ZnPp05ycVzuh/n2i8idJ4IDhb4Bn8faGFKYHs0M4zEmT2gEj
b6ydwTXc5Mss5uGIa/76ktiMLOuP69L1FI10T0BqVkbXAWc+44JPgD6dKA6tYG4l
1zwXf8gR/QGAx93tmljp53T5V4bZ3fP4XYkXiB3OmqNxyqiATkvbw0HVKiMZey7j
um1KlrrGj2f8Aq/Pe+dwAWbNYuDFbcsT6bW5ulYDlJkR/2aqxvfWMywUa0JfyVM/
68BhXIx0pPQja6aji4VXgsLCI+LGdAO0BcLU/guf9k1IxTCF2ebczjEv/sOc6LhI
W0/3k4ocW9NPqQTqsvHjxF3OLKUfTmTpwVkcjry250Vf2rPQMAEsc9Nf1bxEcVWz
YiydoGP0kY1HhE6HsiDqDBg7S4dLjBF+LdXlS3GMqe69fAuKkHt/sJ+kWfUPPQlE
W8aP0G+vQvBEaIob6AmY8g==
`protect END_PROTECTED
