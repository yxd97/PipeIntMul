`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f8iqfWYwPyRCsO7p2i3wsS8gwxc+4EGoIHrvYqQRDWg/mCu/1xeeNFGdQ1OopiVk
OvMHxu3CB/Cvhzj4SeFwRlgoFsOkXbTf3MlwYujsVjvYyDixtZ93wD/yyquDwo78
Kz9MS7qaC3FrOF5O0MMBVkcTiJXcIK4xz/3UeMfQAoCidcqdHry1IaZe2k450kft
VCCt9iIYsnCjaBAL4pL7Y8Rq0cUQ6mn8ytm4y9K/+OxZ42Ix3MJZnWgDk929YwOl
mthjv4q97F75J3kPjZRmGumCf7gX4FjTNhfHVRRdmqkIvWrrs1sk/8p5cScTrd5t
C2Xff7iX6ZrXRdIu++9vKjXV83B7vDqDc2zI9fAhd90M/L+mDiCrx4KjYKt+r3P5
t501rlsD1Kp70gvhwW25BG8UbIDR9jub44nt0LeqfcOYE9fAcq0QQEJQ/p/6ujz7
Fww8wbNHC3Z2i6ccuLapaNBPCX9m3+aUHaAZ5wXy03xCaFTIazzVfr9dT/8uj6vq
AsQ2ev7p2X9AvrgegLXKfZMSryis8bHpKklhsXS7MnW2l0hZyqbRUrVTp3uw/FXy
pDFB1EFKJ0eH/uJB/c51jhuz1k/2pa4NYDIEp8C6SfyPm3fXNjqMu5nllrdXYANV
/uhyDHGPyODwZoO8YuvpOJBMflNfWb8Bor//DF3/0PxrUX+uR5fcC2LSoUK9gplM
YzTMTyfoZRarmAuANhUt0fGW1YK+6iv/eiRhOhbzEtSjxgGKc3gfjFRGvIe2UbLD
OriJ0Hpkzucn9BE8R1i0qhT9xkb0HNr+5GLN0YJfPw2Zq/0qbhiJz1GbZfcmOb/w
rgrtWxCnc2n9Z+JprsNHVM2S7rdEC81RQvbjuA+SnJU9YU8I/M/4g7ZCTMMPamoR
bXikiBcMSGofbftYPqr72ykYQ5GK5hkc+Ok6/8J9aX2jRhY0cZ74q47cwkRFdQjj
n9R+/Ps2YWBNmvifpgB0GbfB/4ivyTh/t2ecOs96RLLSg1rZptOfhz7MhHDqD827
lGUmU28WWWspjcN6McgaN2p81XLD3BC0PQMDStk5qH1lBfhYhABH1nXF6MeMxlj5
WshafqYHGhj5LHDb6qz7vomqplD+8iY7QkTZmuSotA8UazMzC/fR3iNQqRcWF3UW
+9jQBEq5ooD9gqQyNr/6IO4yan5tSBUPSqdrqv1DYdzMySoNQbGcqYfZ7mE61uJ7
OWxcYgzalsZpmZxtoPrfLo/RCQpgf/LpCVnu5hjibUlYGD3/sDu+b6wCDjRp15KP
LsFs6MAornZtAoPjbtTAflkbP3bx8p5nHMZ2MIsBs0qF/+r9h5+By6Neb4N29hlP
tVtqTyoW9Zz8lZBnOBwY9Z9KIpnccWLJF/NmT157wn27q1xE37njcVI+AD0yr0XL
18gjer8wZxt3aukg4DnUgPyZc5/Uy4vFwF44ew1/xV3WDmzddzWYPjcHqL9WwUWz
hbbebSmZP2KGmypPhbdx18G5X4USj+5qnlYU9LdttnlGEWEJNryQU8o3AaxQla7d
DRcigNNwLAypNTcvncVpEYkxZQ7ZCBKO/f16rtLl8DLZw34kyz2UP3p6hjQ6K4q2
atd0kGrm4ktNlPUxVH5gFmOsUUsIUe7RZfgetZz1sxib1KhLiAIZ9vTE47q5KZXG
i9rebn8QfANublOL+hWLoUU/1Q6wVI+4ovh0N0iRzs2ObVmngaA43xHV1zZBVJgB
AjDdI40QzOA7+KTGZu21OEBTkXjXur+18TLV4850omvnxsAqKaxmIFdj9WLUUPtB
h14iTEjltFJQAe7qJnUk6z+IFujiF5RizPbBndh4683k3jee9ConMaMDeAqJTCJo
OIhiPCNodrsROtA6D0qDiAsQV6xq7s96WJJJw6KUt4rrSpicbXMf89HkD8c9FjgW
02hx60kT/3cXa5u4WAgIerQzDI39CsxisniVFpANwTomciKEZ3efpYX6jBciNmIH
hEUxtV7MWB11f6000swMROiVW4C2KHguBiCQxKBV2TYgqrD/Lks02ppOZ7wLkYHT
QJR8vm7NhrAVdT9zNQQpbpt2h4f5E3Yt7sR4ZlcEZM5LLvGlArj1QXk2vmXjcYqw
woCw+4ptVRpYHVHfAw7pewjlaWfT8+1uIHOfKZg/LMiJv9WgX8w6n+Waefb4gSD/
zlooFuo60rNqI6FMivDzXxz1kBa6r3jYsHv/N3b+3cjUQF12NZFNb9/dCq6mg/OU
Shc0ZjtuFD4H684yyrdJ+Xjg2Y4RsCykHwksTydW3J5j615jyeAhpZ1tB82iKjia
V5Sbsy6NPzKYCmvKoLeKvdBfv9rH2f1a0x/9+zfRVo0WCxitlml1yXre2lBeRicu
ikJpcyhFqkYvgQfaiyAQX8za+77U7gzKiTKDoX2eYXkz3d72nrilMc6NnO0zWmRv
yzjIm9NCnpQ1V13vHzHQa/5lN6llQi7ixekBl2W7580VBf/3GARj5OcghHpz0Xj+
8a22w7pq5fOIUDVD0Z9Iexxjog44X5vCyRyz0fVl6u/soxkdFS8DfeHa9vRh+HZW
2LRJezZE5wdqDB7W5PGwa4Do5AMeB0+JD9RLh4zX+oQZkntwG+CdMIeKV++cK7FX
keCx4ZF1BMplYecIHghaxfEbzSc/B37o27H2uIBc+FAu6Vs418iEWeaZSsHeksJa
eT+j8/+Dyl0J24X0uUw8A1BJdteYAkMbyBH0VB4Mu7yNyUOOY37wy8QdkwhsydBB
BYkJjny7yttSChwFSohELiePjYX3+cZ2VJasXpvlJDeXSTJqM/CRt4ZjBxv1XdMT
zFQzaDMFPW5UNjy9JFZxQkrWMJD43mi55SJrNZYzJLE=
`protect END_PROTECTED
