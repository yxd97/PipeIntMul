`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n/J7/GAFlRBa3m0uMCMjVriUhnpTHDJEJtG1UYc6edL5+T8aeQNadjDB+AeOoK/I
Ya8+dxKvJu99iYeSpX/sRxhq0D7t1WafOaV7Dl/ygZNUkSg2lYppl8DKeJ2Fyws3
zJQo8lpRopBdH2Smt0JQ5XQnCmwttE/ByKdDS3CopIW1+TLihKK6p/PRUdOjCiCP
4cNuh4H/VAyIq2JfTLtEKPASBLJvMZJuQDYTHsa4dtLbnoRA/GLNCDHEFaIpUFKa
kd2lH9/scUfsL/0u9JVz6XlX06sAAL3JtH3BdNsZ/OnRyF1jKpoH6+eVz+bne663
2nXtaW6eVcJDgNFyrh+KuqZMGx0PFTRzBvz9QCMio038K3mCRqrHi86AqBf73moI
Fg2p8sSPC1yw0OXgKUsRHHnV8N42fIM0E9t5sdKytlJ561HxycqwqlHgQXylW1eP
141f3DhVys0AdwueLyX7dQAgG0vM29dHkwBETId9o9Q=
`protect END_PROTECTED
