`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfEpggO+UZgSp5Q4jHiKBKH85kvLl/FHoGkshUeyswOm/JuRBYcGJ0H7KZ77ZA7p
McJV2pJkbIPAHg3Oi+TZ8/qQL1Se59rKNabEFZf47A4VJRVFcqs+u6fEK/bxguwm
iqWTEvv1LjfQNko5l6WUnRMEBRphb/Cd+VGlnT9BaJ6qhxBeNwt+MlkLueXY9qkM
W+/Xxx87wRU2KXRlM5x1PofXPh6FL3xTIb5mp6ZAiJKk+4qp88fkJwT7K/FXBA2U
zmntPVaY9ST6LVB4p8nyfbG0wlNnujt0UGGMNmKRdrZgWmlfJN6UPu/PlaVTAPRT
SDU8vcEOztF3YSSGrQjrU4lQH/u/yi7tLifMGwcN4Mks5iC6hWmxG3YEbLZWHviM
hzz7yf+iYLxkfMII31lJxbk3zwF/frOJ+FN7N24z8A6+uSLA5dY9sTiZ7YiYe9js
4ybccqJlgYT+gfsjCkDczRxQg90wfJXgKWl6BCBp4o4kiW6R4B/2Ceth98Nb3mm7
TpK3ppfUG1LTwe3V8eEVXLJPnX8hlhqWtmnCz6sZXUGKC8Y/mlhZ24OagjBNpdPo
itbz3823hr7g//MYet55vciK+NjalIVNwPd2Md08Op7fUc9LEmCiEYkfwrRqNU4h
/w+kMM5k3dSFLkJrLrafj/MN7bm8BJT5g0Bw8g768E/u+ye7GJMx83uRf/Ds0dn/
ap4DK4k86+e8mDi7RoW+VBCUVbXgdQCOx6QalU/JO/gVDSenmEPMDC/tGAfM7yto
V56afoSUOiw0ndBzVD5OHqZ+o2G4B+LL5UwqXTu7aJIdlwe4yAJUCG5w+vAqnrcK
gX24j5Gje0Q2ZsGZVweaB5+UwGM/OW0V5kpbGl8HyG7bG08NsTVe7IRIxjrmo+xA
mGyvO23d9jrD444eYFjP5Nbw4nDiCUbb+POF9YD5Yd2YgtKJLXlPdSYsUqzWLK0C
zzs3ZT0phvW7tK1Zy22kof4+CCpa/lnG9iusvsWyCPlMuymyt9vFKHcv2pHUkTEU
Cf+7aV4HmbIOcLlqI4P7fzVsWU+9HgwK4+cgkVbs5eSoC/k80JHiB6TBvykt+CCq
4eBH+9u0va9cCxacpvNKDJ1FOJfGyicG+6qJDZKSndsTazXq73RI+dfadkkqG3fG
qcmKWtaFQ6l4Th4Op3bdywdFaDSVwTs8A4llf7ZyxWN5nQ98spQ5/iyeVOIgr4VA
n+nwvW7pemzA/I3Xg+ji1cjBNdGwFBIwewX4h/iI6o/flJBl99NPsEAiFXdfvVhY
S3roAj1fNgwb5RyN3Q2dGIzzPM9GdC1KfTbWvEJzLxp5dpBgA9LrOJfZPzCSKoGb
ynXmf3P1lEpYj3gMHElNRYSWC0xPKwupkdmlUp4dL4yxuIG45UNQBvtHSXAlwboH
n+kEWcJZgOtHSBkYmzMKPAiFlu208KtwM3ZpEIox1R+6D9kPb9C2VJhL9HuEDTxb
pCkK3bOk6XgH9fsv7HaIsRX+SHxOtNIh+1SAFAXD613Lyi92k8FQpSg+YVjZVKGT
q6PZ53fshF9X9+rM3qhl0x99/whe2ol0s9Cug0TG7NzL2p9gc2bjQUrh9oMxLU/a
xaoFkyapCidNwXVY/OGaE0gB21esbrezDZ0/5eLloVQad4/waP1CRu6d7a6SWYoS
a4cGU3KA6z4wdIdXEyMLiFZ7zXnB5/xFHHp4rROaBEFA1jQrsbKULGP3McKRQRoA
PDlo2/x9xBKmhu1IU5leTyy1erbRFk9UPdovdt3ifo5rr12ZG9sG0cKLz5K+VzrR
u9xnQspQd5Py01pyFWAdlaGxCRA8Dks6cNl5YX3+U/joYNBqGqdwmHkSWed/lEfg
npYk7dl9CjMMyz+6pwRP2o03lxdOlX0yitRyj+z2SHB2LMXLH88LsXXWne0bKM6t
WL1od+OV7wDxU7FMCxK9EA==
`protect END_PROTECTED
