`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5S6vAwY5QgcYw/AKCaQne6hho9wC7j3BcFUmHge0CATxnuPuv7dq4a9Std6gt3+o
2BqK+2XZ2/s4mWrGY+esnByVDDDvwln64kSFrEteqp3HA5qBLdydTU1repVE2322
vzPXbDp/9Pai28SG+ZAhnNDIj+DWonAh0lm9P+HTTmpkpGFFLPM+L4fHMKhvQvBV
U8JiwrcT4z45Mo+1s9VqBIgWJA/PpYHQPnSzNEPojr1AnJP+Eua8vhZbOK/ROdyn
eJ9RWG5ncegdQSXhxxWiAZKO56anLuvQ3pGreRORupQ=
`protect END_PROTECTED
