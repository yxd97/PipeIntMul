`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1jbtyGPJwL7r0AIkypDUoKOumoYuiCmtxLdHDsvl5hk+olqpppBmL49A05Xc3eDr
3uJj+OEkB502PaHYWzj10X58iNJ2cVRx5JSqQGfEqurPKCRqu5sDbLAH4JQDbJoa
YleWhbCMixJRV4Q7Eom0AO/tuWEbB7tF6XxklFwogMrJrq7NC1JH6NtcONMmhr3H
ka3x7CkGthkm3ctV6KQw0CtfJmulzLw2ZciLzTkbD+ltoR/2SieK70Ri6U6sOyn8
BI/OTvwHCHMY09WpCAeZ6Pi1sKn4lClTmf/Fbfg9AC6hjye008er/nqJ1Huu6Tge
GqitPEcT+2lpVr201XSo5ZGWQXbq73xaMH0scgaxbnKyfCkblO9px8T55wJo1lc8
voThBNbtRyKT/Rtc76wDIkgrsR8AFz/ZxZ4s3qCVWEdFiGeiDq8HvkZpnbt7Dn1O
3kSLHRJkiPjiya0ZD4BdUBKn3C2pO0TzCIfFuN73Oq1Qp2t1lqC+EszFvNTOUdGk
IeZ1EXVsGzi+MMrEUAk3YXWWupoqOGMe1IaYEqh7Ot4=
`protect END_PROTECTED
