`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JI7Llm0kELCeklnXiU0vdZ0jwBFoP2rvYXLa3f8l5P+N1PLtm+cqXGeuSlDBKUoI
8LvKMv4j9/1O7THpLily271UR7Fxg0LWN9cR6jeFhGwuFGguoV0+N78pS1T28Co9
jyU17x1ZyFgzk6WSVrB3SGtU90o6sLfqB+7hs1rKiH7OPU789Mscrz1cnYlly8gk
zlCpGtXXEeakgTd+AqQeeZGXP6lRm85QbQBittaCXAYCorJrqjMQwkqqDvkK/Pok
uGfaXldAF+w0vqq3ZSUQOglOgJj99qLlpqBGRLwbDu9Iu0GmPwCSy4ps6ruIAiDm
CnhqjTcniaI2efcWPOQ3d0+OYTSHgKOvSGEiTpodYMNaIM/przsVWFQMaPK5qAa8
UbhZF3MVX28JVp4wpqRbZobx2F7Y2K+SEOkiKjHBmFfTnNEffQzXjEdA+qXqs17W
Y9KU6TAbIQhEsMCRDQa/9ehlEJN2Hh+AWyPFu7YAtbwFaV9afS+zRwjAvWP4PIes
jq3MyTswSK5yIg5r0+bGxkCUv98glYMn4pI1NtKVvDqvx9EUHeIUdwiJpN4oF47y
1BcIW5IA7ZqvYi3DMsWiAmsaStTcQ4ehHzCCOWt7BXsgoAwsp9vMkFf+CIHJuT7u
XU93lTetdnF3Ry2O+r93MHdh6rKcR8xcK6FUyzzglLOw48jSXvgFbFEnvgR6so8F
SOori8Xfj9+kAYhnsOIWBjmbgIwVveu4Phu30r78EKVl07ki3v5K8atnyyDfOiTk
frPLwmDDGG9feZfwsbHRCc5rK5AYeJIDu7Jnr8YqVmitKDTPYjNI7sdLPQNjlxDP
aEsJzYgJypU6BzeP2NTn4CT5rq6PNdeP+oVzaQRIlvkGARa+Vg8MbKpfOg/u3SvN
Pls/QEwUE+MFOt2qeUy1GRZsi7tNjpE4YhHsmRS76XHqlYf4ZmsumQNGZNGTA5YS
Btvm/cy7X0WlV7SS2VE6tpbOOAretNaQ4MYgbLwHE5UFc4bFlCy2Ma/0ygKH28rV
Unde3CjkLSio2KnncbkfmM/SSQkuASDZ+tBqkeqs51P88JN6m6r1AmVs0ruT5Wzt
ev9ilvh8967XONhToHq8Rw==
`protect END_PROTECTED
