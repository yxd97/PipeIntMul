`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z+i5qD7R6Mz1pac8pc4NDMGLyssxsqfCWDovifqauPMw7UewJWJ0o6TWyQ6iyoWP
BtXmO07smZg8Ky20vFf0RyZZlcZ7refiCMydJ+O0ww7ydOEoqwZ/g4aJJRsVUtTe
T45R+R6X3V705EZZorWkOQw2dB/qmwkELxI9M7mPnOE/nkbjUrAtpTHLhID0CnF9
jOZG2Kue1HtcXkdG/W55gsQNUvBI50ASwiyAyhD7QVTb3q9we0bMrD9sDrt4nMq5
WT9nziQMVfA+q8iwILPTcwtv1B+NS3ttzSmFtN3a6hNNR3kCqwCGqKj2lVaqBFjS
ASoFb47WknpHGUCS+TLJqL5XFxJEDf6vZTKf/0nf1FXYcngpfuVjlSCn8Sjf+ar9
XThMm6ecMsanhQa/TKThRcTyxWjBb/fPCJYK5txrope1wlaoVSAs/zopYMT/HYo/
`protect END_PROTECTED
