`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTqoSiSuSvz3BlPs+p9J4X0NE/muQTwogVukhXdkXIFmHlJQ3nk3T9TKkGU7dkvo
J1b8Gs0faIV+k+vmlXOOUQgTrIY/56gGoaEITzQYuO7avc0q5esSa1wKIc4zzt1I
BCwCZa1RLevZD/8G6f5/7uWVLRxWi8JQt49IQROIt7yQAugHmmu6PgywEWREPesL
6HzS4OZltHEoPSBPkVMw8hd3uiQirvn5hpmMR3L5hXlju6YJzgXas+a6HgIuhtZw
Hwp9+MWlB9z46Wj/FDO+rQd/MqkXA1kYl4Bcdsk7JrbGM+PVHywf6Dan/HbX9XpI
fWuZLy6kvIM81lK1lHiZUODuosj8c2c/nSHywwgbr3A+symn3t7QlNoZB/ClZxBZ
FpNxhPaRPXt+4rE2RmLMgCTNF3suzB9ecTCEpwGYnMlWvFRnvx0oht/3Y6xrD33m
kNE9phKFjndbnIviZg3DDBw2z1/ulbcH3fbGDCcDw/s=
`protect END_PROTECTED
