`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
59l8wv5Ru2jcoUG0L6I5P1nymSGFOQlopT8KDko1Mdx8C2gVunfgp7b4PfMWXd03
5YGk6+V3kN77w+MXCx139vN08OUMX+gQ7TYiKNzSMAF1jSa7NbjMM5YJeEKgFe7E
uhj9Tt13MqZ1o99PzCuQ92JkFwsgams/TEqL4/M+9/Re2Jeho4Jkn2q7fTOWM3k0
6MzU9dubwyqicKkocYkr/PW1aR+XReqZUaRbe0G46IbMe6wy3aQHvvPJFYrRIWQ+
y0tkKWpKTPLpKBurAiwHGfWIhIH4cVmt/k1x4SdMh2MqcpW06WHlNn/x1PZLLcMT
3gMRwUpK4LHoj806Yn0NjiYYSO2vqGitTwwr+kcHCf31QUFigp5xVtAJT0lybHcV
wpVBrW94gy0Be0ZFAa/1esI/NpC77EH1V4wqzXgl26E=
`protect END_PROTECTED
