`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PgpIi9BVIXm8zPA/UTmR0DURi6rtK5e3RFB3ZRaUtBx/ILADJHTyzp9BQeiRKs0p
L3rst9ZNZdBAU+5m5OUplb6jyHso/8GO1TEEoGEPMJXnTz0CzsL6pWPpEacNUp1q
Soa3t3U7TpZiE+9Cu6WJLwAL1hzJ7BW9rvKei6mg5pPdQ1jQ1jw2iqWxc93ueVKP
Y+OjJEcX16DnjJR2dy0ZxTAbdXTwAn8adsix4NnaxDBH+DQkyRfrh0OGGeguITS1
/0lFF/0wudqHYRUOPjM6Wcf7BkqrM6LTyph/U7H2h/ZNU+7cBqXtWfWM0bXsRcis
PVrIKnJcdNyd5eWk+aPeqinG+vMwHReQ2DeRE8NXP6okoJv6AVP06vrX1rOt9SKW
qRTNHTqjc510sldBpTteTVIx60qBF6HpYXjhx+q4Xe/H0AZMuY8LqfTVEMm3ttTZ
bQGWV+ASjKhxK6jzkpljH90GwKbNwnRJhawcGzz768ldrqcAjD68LNNtoel8FmE0
EHRWT2Zxd4DF3arWcjrc8JgujyN/EOthT+NrG+TweIBCIE5p77oA+thSQ7lQtOhm
FzrBtbkOpSby6x9eVPq8v7RUJKNB/PiFifpBOmCMfA+U7R0cskMMqt87EF1wpv41
WXx2AWYz9X6ECgmIKC+9CV9Zf0Aa1fKKBRbPVN4k+3CLl5LS57AR0rUnpA2TmZ0y
Y2pRioz/C4vKRZnzlqVlI5BX8mY1WNSLUItzooKtQhnVfy09QykdQ1ghXNCZs+Ap
QZOwCz9kR4nroOapmZZBKWtHgwAAwYp97ocYpmRp+Nlq8Ka2IRqcOwd+AZuVIcsV
QbfEcYwr/Z4qCTOg7BDQ84uEgO/K2oa1KU57gEHBijm41sb6PAO6L9DI/nqzwUm/
gOXMnpDUt0odXG4oekF3PZo/5pOCuX1RdatI2oetLpFzyfkbt+BohaZywpp8BLIh
DH8c9fXz+gPMxrbcFdKRh7T+X/sXTpcyFRaYu7ABcQtvBk0TjmyP9i020MpugYV4
SOCbe9GPAMT/rWgAGaRJD+eFAI3bVv+uJdTpa8rizHYeEFO7wMZaT6lGioHz7WIx
+MCo/mjLtFW6wmXS/qY31IDiShmx3PQpY4a1qGebKt2KAXueFCjfZC9wKpK7/dDC
4jQ3ez8t787whi8uMGG6GhUUsrL9ojhapk+AHnQoKdsu6LIQaj49INdPjLOqM2+V
pRygDKTrp82LvHxM0YLPG2pwSvSkrPqWWDf1dBF7mFDEZfVjSwfDrQoEvDf/jozA
9Nd3mUbG1HZiHjPmpJIRhw7hLZorbZywQL7KzqSAVORZBxWkayccsQtpV2ZGP/91
w4m2uHsFL4K9w5F0KDVupe8J/Ymz0Qc7JIkQTzYwrSuTu33Eft+SM3XHDMI6Vuc9
mBAoqWxUd5czi+zNF/kVYpMh0Ay3AZfdK4JsMb5yIgEgLPCljRJ8j8eh/jOMmfKT
7cTzm2T3y5g9BkBT+sJMffVruuqWs0PBtjv7Rd7MWc3bBVcBER7j30ZrJec7vm8v
N3nLhrhORExhKSOGeF6xq38s/HzFwlAzABdbtT7jqTJ2s4vhZ3Cd5djfPpBbco6O
7E8eZn4SNjBiyOmueLOVluLapSYKN7/0Yulci87j15wO6wWHJRI2pNJRBPVOYTjl
ewDqwk97Vj8oVo1ka2fjQm4apF7+JeJlfr2tHTa9ZRP4DK6rLI9Zh24pcfUlMfQ+
l5meIYyonj1HGyIW0WGeXoZ3x+6K7JFzjFrnv+Knzq/6ZeMtFX7ZRvnUNAoDvcFW
9/+SbQqJTrpNJLpISCr7j5J5rS5vevJcHTmMffQ3L8ttCVSL4XRpPZ8X5al1vbo8
wpijACck2gIl31kVtdndUEYm3G6rcra+ffvYyRdIqmdNyuNHrKCFRXegMohbVUMh
tZZpRCzE3KwCy/XB44I1AtB2gRI7jKkrzmRgHm03sIaanGHNx8nii5B8RGFGb99D
4VIliZxeI6WV262Bmu3tnNGAwmoae3EgtcUnIAcCYcF81WKKj7ghjRFSWKg75n9Y
u0lqsrlPJD2u1BJJpFAsdw/SOD0TfwEWNr2MYycspt2zbkuACaq5sGd9pa0FWffR
/bY3M5S/PHYIMKAof5Wy2B8JWfGp89JV7YCNCX8w8v4R6v3UJJvW2e/C+ELNFTiV
`protect END_PROTECTED
