`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpJBSJ+c6wZW/cgTyU9OpiGLQDNhIPo0qeq772wQzk/K6Lm1dOmQeCNGS55Alg25
KvV+bJvMs8DjXPTrnjn3/4AHL3OWjHjSeTQW4taJslPtgXtPn3Z3/ne/XUdae22J
s9Ml/55keRz3VDYgAamQRk6ywsk8C/qAwlFoXKRQVWVM8c0ODMZkUPKSTdxQAT14
NS3Hc7WRgo8YJ8OMep6zVnRWTAyBEE/0ja5+xpRwwE0ldwHrCTYKmODgcJLPWoE0
KrFeQlhZjVWqF8WSa4TYYrnDYbQNCeDiXPBR++sgnJgpa7N0BpWJZUQsZq++SZP8
ju4qNVL4lTSDtmg4tnbxu0QwNGGochw8MbPfEEKPmA9riAR3moOlCt+MhBYcTxXz
Zbd18TllAvzgTUW1UfzrHddWJXRH7IVcu9mD9iEJ7Jovne8JH8ujarB+8Or4xe+C
zQ5jnnuOPgqbDnM66+nFVljBQZ1HjZLVZJLLwNKnWA1mYAIEdtcpjh6KSKmkqqQD
P4+LEXHhsImPAlUdJoYQaD5RwiZuzEAxkobE2aSM6h965utFxwlLxeHUN3HiYhSy
J5UHy5QXPSNe7tiFgZLG87LjJ0DFTQvPVYjIY07MQsSTYrcYWXBCZMUrUmwMbVaW
I6sd6DC8XmaOmXF6Lmx73ST751ClPMkNpxD7zcc+Gs2T4A5lq1zembY5ifIEhjpT
rY0vQmSyR6jGTzA0CJUxGZxg0M7ZeKv2pVb88AxUt4HRdsaeqXjkSMiLw/coUP0m
JVCp8E0mfAIERrHedI2y93VQZKXy/G7mWf+qcIQclUv9tDu7CfSaRtRZfs3yTjq6
0544aqyBzdWS2wHh3qpD39Gn/5/1WbKO4KqOtqYPIRr3ILyV6VX+att2AiC1ATCE
2w2rqkI8mAPjF+5y4auQYs+gWdF05QgGut51lEHBra9Yn6RUPVUVt0qCuz1ksl9z
vVJTVMP9TiN5FflydiapqhKKh2DGGp0Q5N1p4Rgto5bNf9h6mAxGAexI5GLXPKbM
E8mTaKdofW2NGc4g6nGT/Q==
`protect END_PROTECTED
