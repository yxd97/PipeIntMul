`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tsVGCsegTDjor+7rWpxlPB2yO/iZtBYIiDaKDNlAteDh49quCBPFyCLstPmzO3n6
lnXa+H47nBEQPu274/RmTMhEM1Us2AfEpmNi39LdAbK6t2EI51gs4jgu1KBMRuAN
Sp9dAFLvHhei58quysFD2ajmdh5PfIaDIVj/+4aDiGdlYih5crsI/7c/OafJJubn
kKAhYUZ5lATbk/SxdJ+MvPSePpUVzs3Bd9aVD7vAYcNSOTY2hzOUrFZfIGx2b0fG
P37yCqiqr2dl8jUyDbzzUsPfX+VdM3Ngq8PTDPQN4Gwk5CaQ7qD3oX3HYDgKBjrH
jSp32TqJYIoSLkHHhe0gk695zzQPmS/Uj1EfrWKw7qsuYk7JRK2ERSHLgQb64CEB
KrSmHx2jOq1XG4Y/qSZzjGqSYOaLuOX96HTtlEGqxw4=
`protect END_PROTECTED
