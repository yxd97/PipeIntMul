`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XeWmYWGZXi+P42gxMPaItO7tsvmbcVM+LY7yw5hzXSgOeRIomQeqzLZs90rXdI1i
87TwP3HSNDxrUOWTgMeTo6vJpleZF56NAW4CJk7LLCTfxIa9G5BHVJ9jeZ5wQHn2
Rn0J/H0uyWx5j65GN7Qj6hArL4sh4EK+4/ZiabrHO8FXieMtyF7znfzCPf7KbrD2
XLkN+CmG9N/6iEZS/M7JrFuBiz8M+rAl3j1TzQ/i/YIPhx3WQO2RbrcNpNATJ9G+
2ddxx06nTJJ6bNPDg3TcOMzkHGMiNsyh6IogYcCd+Lvp5J8pzLfYf3CDEda59xFF
wYQWtNwh09N/qZgYMoIBLSPbtODCft9ShAA3KcXldUH8oEWH00jCssMxJhkvdJNy
MyLiCGuQRVP3hwcyJqQq02EXdSjVwrnvz+N7W4zqFuw=
`protect END_PROTECTED
