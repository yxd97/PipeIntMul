`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPpTRvWR2PEEE5+Ueknku8f55a/9tEykG8s8DSKAV2kT2Ox9naTrGmPpVxPoiVcf
PjpPxY2NCQN82KGBWPHdmj14MntwEt6M29IG3rmF7VMdqxWKUB7vSvKBiSLF4qbE
heo4stjzrn5EpM/KuDQ0gJrWYYjyZbzjIH+/19gZB29xb6T0WYjnT7jOWuI8mq1U
XAO8DsOg6sNjke4dmpKFRxJ1VZ4Ga2+pt1U+cPLlUVHKYj2yUvDVYXgPLzQlEDxe
4cNdyrZs/hjw2R0i2wGGvPVgNNGMXR+KnStJNN7MZ99JHaw6WkZsBy+f84QntO5o
51b0I3mX4K2rv8ZzzYbIGW1DbSAvyKCY4IBUH8TXUMXxib9LFzkfxYkGzw1GH4m1
s9ny+A19IcRb15uI0E/uLg==
`protect END_PROTECTED
