`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d8z18yWEFXEtiaPVnbELAzGg+y6XR7FmEphG4OrtTjhuLCOHOkMPuRqcke/K8CkQ
8/jLN+GLJ9ywJVhcBzofo2mSyAtU5o8z5dEpCPNLSDde5rBAo/06z5p2yPzqvAVG
lv/q/0R7/8Cc+Br5gIrM6A5T/iJ1jb+k73KkXyW2RvRWPiSwT33SoyZ8H0iBkSO0
/PJ9Vgz64ZurQG7W6w6lc7Q8xgq0PRM4vEjZTo2hyYvOWZyp4ljVoCQp4gBBWXEG
EJ7YiO6XnJtIIUol7ErSQqsJV9CAnrH10mVCBesBW2gSUAjT2bQGtQqPCC2OeM7S
kKIAW6F2TY4G6597LdFEFlQUgCOnQ3MZeYuSD/rHtN8Ix0YeDEGGIPrEKETLQJw/
hZqVpGJkrVMzIRp/FMVTZ82ykcZobyfuJssSWpmvdUSMipDBgLZBXfOOQhQLqatp
51kCFh33FZwcWb6fNU271H1bAxzvBGKeoMW872V75LunVvNPrhTfGxGwsd5jjgM+
sKqOVq7Et8sd1OqZB9uM0h+I6tjotvijeWItmCGzTvSiP6m7OPpKTxN2Kc0gjmQd
0BSMdl02Bi2P7Z16sWgxNXjNPtdmrW58QfelmmrdfSjQz8/H4JNU12xFvDd6+QIh
hwQ6pKv0FVkUUMp/8lGOmjNkxLE/CPSqvQGbnfjWbKiDVYFk2w4r4qzlhX180VhJ
OtgBybKizv0A5yaqIesV7yeFh0lBUu6Rt0IA/rusdFCLOf1Kw9q/wLmgGZveMoxD
lCw6MHuGBePSPIhRm2JEZscOn1iH7I/72c/G4gC4JHKskKYavFsuvC6HlCbOgyy+
2GBChFLuBjKDlbgFxkRWRFkqO4efE9oKtLZa+iZ9IKyr5nZXii47lpqnNgqIZGTg
way0DucZTZpPwaUstsLBeg==
`protect END_PROTECTED
