`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nA8Tp0dbJOTt07xUOKKVi+/G9+ZMLwWiLlaxlu5COZnlkpT/1zCv1SmVQHm0xnza
DruP2KSOpJv3WEih124LT6h9pVE4opnDkoNzQp9xWYaAj0uQAZdAXo85gZyUGTpg
zegw/ZIkFsBymx1V2bfIZnMwxqfKzJMMSTOC9GJvq2Ov1yxYdF12H2vaNDnyVPCQ
rBNwm6OrAhQg+h97Y+L3Rgf63F5+DEbdZzNq5h+C9dI9S/gfwXikvTIX1ioCe712
NQoaR3LuXDdHUqdKfSI9FekmOqwT/TTS+KSP3CCcsw+Es4FYmxk7bUlEG2F8Cf0C
tf1YlLSFVZylP92wY5nBvKa4crBWpxhgDQ7xTz6YLn4HUjKWXX/k/1fgGqhyJOc/
XZ5BRhQyVfXRh8lEclxdwS213R+QuBJNDQkissjbRpmqP2NvuArKNKmYzkXhQefH
oegEPXNC8l8rAklgoBtNGXxkVmUfQLmOxxwA/xgw/2fcXf3d96qArjmCxFAsQvsR
3etwYmkG0eGYrBAbQnsDCe+xtF+K8Q4V+nj2ykcrgwfJHzxGgfr/GlV2LFc3pgZd
0f9VnI6AKXDo/XE/500cN+BQzpKuZ8mFb3kDkRMH6kvQVoD08+Q6pbdY4F/uZBnJ
rO7JHAHoVHNfziLi+MTYCAgRRZ6kWsiPJR9PbyG3oyhqCjY3A/pkNJuJcpPcdYEL
KERAbp/ZOE0/kuNOaHpkig==
`protect END_PROTECTED
