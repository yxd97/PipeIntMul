`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sYkOzO/lPSmkyaszqgWTMPZbQrlvQfNrAmCISK8pAjnTPOSg+5GuCE6DBPGLRUGn
bJFmfM8pdZk7DxHzlAOqecIhrOuZTRZC3K2+co8xaZcC1AOuGOcg1RE/tMqZmPRN
FoXSyxKx4xm8Kz/mR+dTp5x5GzbWZuDeS+DsYMX9KF39GQen7/lAA36+YZ2EDLSC
2MbBc2WTacdKk1HxbR1EjDRfocvylbsOgDZoO6vX5wGksmCycmaOm6aKm8FWjlrT
fE5+U9kLCVILpZ+yPMokbTT5IOU0MsXXOPFxDJDcbedN7JdxQRP7PFBPTZvCga7R
ofPfCIM/65xv+utyfKW583S5kxDygoTUF0l25M5LoE31na3YiwulyPKdbH5RC49l
7hl8RO2UnPapS/6nKFmk73+LWMcD920XztuBVNUy3G66RVafGcnO8LeLOhfaSJBi
B9U5rjdyLFiQ5jsm591Wz8FpWbOgQ4lLpvAdzKIA7HbXhOdMXSPRN+HbNLile97c
NQ3QarI8oZO9mZhLsvHlLDBft2kExbRBtygbwe1fIDfsNLtCzSbidNEl+EzjHzIS
btMwmxHMsg2+UhT0Y51wC3ejQDmtGn9+FpjZqUVpTA5nWWXywmE7+vgw7ltXr1pE
yhrf5JkmZa7nJOHV+4dmMu83kB/hZwUMd1zoSTaECa71QkR5Zybo0KwEugF6IcKF
60CKfCXwcZq/CK7nBEk4yfwLxcfAZeXUZ7Nzrzuq+nDaKClP10/nhXnQzzE2octn
11D72Hn2fasSLMyt0Y5e3AWY8Xz3++PeRggbpGd/0uLlqCoFqD/pqBbJJwFa7kRg
ZKtk4Y+44MqJHKwjFMb5jE+WePbCbHHLAJ7QMnX/p0oaGrGgvN/o21hbwUtcTdYR
PkgSalYsbY6GSK8lV6Kwnzc0YV5/h7govaZFhICQAG2FhuugQ6wcW+Dq6fect5+m
JnjIt6aKr68GP5NBvt/b4Jpv2Re0p5X1xStU9I+lTXmU8t2wcBs9LE9lACBsmPlY
Kv8BCfigRy5cH4bOz3kTZgsfCT/r2QRjVCpIIv2AxYx8OZtAeTkpR9ev9EOzfoDp
C6ADlr75w6L8So3QnynPIHkYSavaEuEzDqPa9Cl4qOVRhZQS0h15eVFFMBbj0gly
`protect END_PROTECTED
