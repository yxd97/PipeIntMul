`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2lAhKmXHbWRMkB4vkzLC/MQewKcAqUyC+Mv++6e13+Hi5LVXzfo2vQPmPvgFe2U1
ynbsX5GtwndafbCTwXTj/yfi0wx63DdLZcuuLF81lHxuEKB72RyYnpDJEETc8RW1
BXJK+GqxkOT1eUIMHyy507fN70aHXD80eJC6AF7j61GJV/6PtML82UiDYyz1TIHs
LOi1SRBW5aA3uP2dODq65vdt5GcnD36/aIKIA/LbDMI7aiSQrUbM52BLzp1KvJT2
c2uwTcEN1LoOytBkF3kSidQPGXSk6r5d+9FR+gUiW2o4hDfKeWtInCUDH7D4JREn
RIMJ53Yc/h0XAttkXDDOwvLriHzZdHZiYVhmlone5XUR1u72wsbEPtNmdiaWpoVD
sn6Iz4Q5K7sojGFbER1rPAmyRU1ofToRTh40QClE0w07w3OV7LwbsKfOHQMuZrxh
u6GT0NzIkYNo1E5ASmRDD6BQ4bw6TzP8ayPUlbrg5/WHdk3Wg2Ob6buKOEy/mShO
pil4AajyFqDO7ikf6YZvp7cgrKaRbAwaSqsmzMSQnJwNb+X5cUHqIX433SaWZ2cp
wkTPX4uoT8Ztdn4Nea46o9nmDxmLQ3dpiKeBSNoqdZFcEeBQUDzcvOwz3fpD2MOj
J06wGvllx9J1Smo7irpyQA==
`protect END_PROTECTED
