`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p3anwpciB551DxipyCGjRr7PzQJBjjfM3V6BEQFIQk48sjPSJioy9e8XRw1Z2Lu9
B5deOQ+L1euG45ucCuynLXQ13nUZj9A6w1xuhhiGX32Ej8QG5At9C5XSkRwKJ2cI
K7ahJ/W2r6JMA/phO8fdHSHfjPs+QH2GDvoLCbqnC/xrvfk3pxLX/S5OQHppTTDg
cZB/O7V/JoDUABpSOjlFZ82uezCUA0tmtVXnuJRxcPR3Nmq+Vh85KHRdTMQdcvE5
axQwyQvu3bvA7C5LzeDFPzaNQnprzSO/Jo+H2dNPaqyGjDwZiwSka2Pg7ksokJqb
LXCyxT8mtk0FP4Ikp6ijK5SxY2a1oKX0Cn8iWFO8V2Q2tLx+P+VLEXbdpSNmCvoK
sBhnQwAFblxMxnKnAwezVS/tnlo5CGXaC9dTr2kB3hcqR72ITzPM1HWOvXzfZTsd
Bedqer0ber9+C+dpqFdq5vm7jl0v6hUoXIAI6B0TRDPIKnlKUpcbEByHQlbf75or
16Fu9BIiGQi5MozgfJqoG4E/UkhAM8cmXgI9xfiCKhQusiUs1qUCV2Rcke1+ydLd
8BeUZy4k0GQFdjHzZT/9gmQiEACNfUt1y9BQm5bKTyYGnRGQ3t+nXR4hdJSrSWTM
MswYGABAghOG8kgahgjBVWS18NHxpvMJAo5niDhOUyRX1tMdQO2kYDmB3W2adACd
UmCt3zjvWJFGC9owS7yh5Kit5ZRYF8FtF5u4935ptYVwovl+antXvOV9GKbdQl0E
Jx5oLTMUS2rLnltlO4a7pHnTK33BKddpgVqOUaQUr1wLOJQkoYsgm1pyXK5a/NxZ
ffE0Zta7HB7aZB4RRMBV4DsxieTq12mmYUx8rF1qikXq/ty+CL8xMsgrUmNdlCeQ
I3ZGlt1uR1FDp/LplvHlN7ahgQrWvy3OSsZFsWBc9YpzuSX7sB7Gk1LDYUWtDKiP
+AQ6WmaBIUAgwYddDyeWqUhFp+2Za5yNjlwoQIvuQB9W1YUMKQzsyN/ZzIyGH7MF
YxsKvZr4sE/Bvef/p3NLKdJreyrCtsIU4uWzMLpIAgBykTvXIlYntBsb9RCDg3cS
WfDMLzmDefqTqpXE0QENp3D6IyAphqjQoZejSWhvATlgBJL40t1FLRP28CRHZllt
vlTbhqP72GsRpOt2B376vR2v9TzcltnqshXdBR33wrkgl1OsTYw3FiUaWBL/7zDV
vXrXvkfWQDkiJQGRNFoTGlAy+Hem2qpk99fYK1qJqcyB09Q+pQB0I5zlIgXvTpDf
7Xoxm6iMlcaBXefwB2mwDkD/La/TJKKIENTu0WKoYiPGoK2VYkZ+UpqhojBHLTtX
9QzgPQNfr4HgY1ui28THb0ooIDIEraaUBwfN39u2+QFS6EJZNIENccelWuMd9im1
zvu7oygxj4P6c9auuqOydWTnXhv87RwByX87LufyGhD1Wjvz9FSAQtTdPqJJIgC6
8SGcKyvwAMlFXs+eZsVr9wc//ZT/dThXP+8zyjSEgOJbFzsm2pKdTn6eK90fCYDt
WlFukn0joxNeaW5PbbxeLtqjROHGUTXqndjG6SUGYcruya5swxwUY9gv7vmJlWLH
hDvh9xKQWSxSUI8LfbDGviTK5HTiXEj1sGDL/OV2RX9gfPLAzPae4/VHsWMJ4ray
7LLEU0tFVeJE4olqlqyA70t1F7x5A88RlCszYeV53HqfSQ/I8eEE0A0q3PPf9m76
BUL3AWXcJUDETlXY61bE7kQ0b4k1TeHPukkl7ADLwgQinEL3RbXBSbCLmMU366Jt
jGQKR/sZCOs3Qzx06Ik32xRjeO79MVIIhoDSuDXeUz+hP43A1QxpbfLPyiXvby5x
G4x/A/VUTwa7SDn7tr2SXAl8Z74deS69pZyFwPsfwddkkK43pOFu3xDV8P0INxvB
LwgtoBch1L68wmnjxJFZ0jCdh21mhbRCAapkOmeFFfewzUp9kg8JAEVDe6LwWhW/
QFtvbei0PERwPUHCtIPNo/yCM+JPjWrA8aFdphQ9ZKetftSt5eSSaypJAb4MBAhV
W+Ii5dUIj7hJvsZP5WnDVvjlkg9bymfeV/mtMLIGxp3tjk/J32EAud9Fk0wEG62L
AoHF7kYcf5QFOsEDbu/dQz2LGpLxf/rTVrcwKbUn8s8FBEfbDEIpXR3yD6Gv5oGD
CgouzxdfbuAL481pBpB6/xlSWx4qB+TyptH+o23EdrycOVarfNd9L3rEytQ0brVG
WTAKUuLoEHzWKH4eO1EiDtBY4+ETRkAkIHcqTzm59i/c69aCRq35DjXSKLw8OjIM
cPpBqMFmvD/CMR79K0YJf7KT4kOWi5K7SEhtsRb5n6fc695LdJ7zA2+UBRxMwUrZ
H3uL+fPCpVo2sciCiCmJqFwaWw5EZDLVMM08tz1OlQWuqzvK7ibrKvMGwow7t5TQ
iSpvyOr2ZSFf4l4KMWsZNbDeXILH0NFENerZA9Bxkvi8hdh3hKSGrNEUJRsQ2ZgY
aYA4FjtErvShinjsZosuFtEzLb9R6knidZ6sfYkktJZndzMTWXeX1WY7AfoeWLGC
JKDa/K9MwCXkOxwPxcCiGhOVvXMaWAWoEtpEz+QuOm6kjoLiS8woLTj+B/tv1rBR
cDsNBLzgxdzOt/wNFytLXwG30GZLRT42l8htPYqzu7VScjPlvdO/jk8n0MageaWx
GdLuFkaj9K+IPgPxp8MyPDTLemKQZtmbKFs7IwLLRTF77v/5+tlLDXRV4N0iDFk4
XZwusAJVGmEHoMVNIfp9ZA0grMruRLbf7YGhTZgusWpYmd4MgWys4JPD1GrTxUhB
rJFtJ5Pwig5/oR4GTUtuosTftR3wK4Orz3M5RpiVwJApYtOu7yEoW+uygJZLVNc9
2d529fXhCmCGFOCEhIAQKz/5/ydeLHKANbh+hFGXvAIf1TKq44lEY312CubN8Uvd
IpzwV5Gqei1C0c83+3rYVRsyAUWyGMhNdCiQZQas5bNtmvLJL0wSdnP5BiVgnJaC
s0f7R4K0Bjx+APpO32/ZPx1Q4ErIHoK4tOCqilb9yBKH7LXVNVRVV+rOkWrnrWZV
LmZCjn82DCRL0s17RrVBywRSlSE+IfP+1l62d1vLXiMIAhkyWgMXLoeSvt2RI4v9
RDh+F2gPMWg9hFETT20+dchqpWzYDGC/JwSt1MCkf6ZHPMR42UwCnhXRZVoPWbe9
p9Na28DRSZmaZYvKYl5APd3DXlGro/AaTQGLV8PVf8QE8t7iQHUSO8FrtVCJTdQk
ZblkRB2olAC8BX/QhKWnvRyJiuoBRaIcnLhOagIHkl9jBTbRvVezYRNhn8wF4+70
Raf6gH2xYMbRQ8iMFoZa/BS9dBCBAMsXIUvNflWvsxBpDmIEzVvubACXwSx4F6yZ
BzMWIygOjXxa2XiPJSzxyGOJXUAoWetQbyOxMpn+HagxQQJQwMXrZsBV3Uf5tadV
Rguh5Y269pPJyub41I2p9sbXzt67CykEqRc4H4lnsjci5t0yaF+BfUQ3qORjtBMI
aKdGi6I5Rc0oURFGdYqwH6cZwMRmnqZDBmuO0RD8XqjanZsyQDqdEdtytCpXKyEd
`protect END_PROTECTED
