`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KZxU068yjxPvOzdIbhKzugJbREWHuLWVc1+fwygxvm8qqXZroDthZfRJrbc70Z/c
XfmpgC167dqv4sLR6takMiHBViYBzf2UQ4aaxQiF00whzIbI9GUOrxHWdb7hA6nh
B7nmQ+1EfnP/TZQfxh/6OtHzrJ/MXfy/KgdWq8XPRXfpxc+iwwaQN1XtzhO3EsCy
ah6ypi3q2nM6jY2D21hfuthN7HAziCeaiNzpObhaKHlrzgsakMAfCV3hhPDFTt5O
xSX4vpQ3ZuCNin9xFm8AIiPqOriLPPNIEobBIVA+DvNMHg3vKUlIW2X4R/B3T9EN
DQena+3rN0RI4fKzHJCzHi1Wt4TDRnG0fSxnGjylHHrNQ7D6yHemCmE0XATgVUKI
TEs6aQjwkQsFhYXXjpUlkSdaex+AnL7DSM1u8+zDuCTnB6HvOqwlJiSXBJ+PXD/Z
bW3NpwpLhYURi8CxBuBuDOUV+XiLHfVaunW0wuJFKNJsFkE/l4isa20YCrDihUQR
m+2VMGeyAeJywTT5URjUQR8tFp823NdS2qNq8E028AftU10MMGR6uhfS8M4oJdNC
I99ldlfy6elpejPdsVSDYoc3S8wQgM3KNBCa8y6UC180k2SI9Uv58anGsfaHO47E
4O+XbvD18IcKny77wHMKqB+E3hPHDJaiyEXIylU0qLCv/R+4kEqbl51wwY4UQ2vU
648U4+vk8vDZfF3X3ZV6HK+rnxHckrEXVYUfF7CasAfCQvnrWT96kUVy2U3kk6FR
SO/yTp+5skFAS8PadLSDwlEvKt1OBV5mJR9UYP5VdMLmKuh+XBXeYPizrIJrd1eh
0yjGmIl/Ydpt1oczJEewfwoxflCA38spK51ph02GX84W9Iul27k8vJKOzRj4ceY0
/+LMIfglJAqHu99b2ItM/9NBOo1i/IsPu6zfw3uHrSHT+myzdGkvWT98w8nZ1ery
2k6Vt5TBhGyMl7iF+wB8YqU3aDQspkxgKVzTNHGB1j0teIk5LUdDU1f7YDzOxkqU
Zf53ZGsnIxd0L88kUlrr6QLBx/o7tomkm5odeXW8d8G5SGxm1FqbcQ38VYTn8Yh7
gisyzVSrxqmI+kZQNv56+yqHwx6AOyVMMjeoEMcL8I5qJctypHZPv12VAbsf1IcS
Y6mtou9ZTWq+q1KHRxAScaE5yBdY641rYXuQU9bz7BHucf1TmYrgj96OgOcNTaEk
sgR8Xo+CKvLNsCnH3zGX0s03on4s1Krnf9uIRXLVLDtx2RUMUM3rpuloWsAGalZ4
EbVDAcV8w9XjWsTHxnJOXdxm7gGXsuSacQD4fMjFSLzBbifx/2D4Q8PLuUQAvT39
Hik8/Biv1Wz5M6nKkMN57p55T/QXdnvGxIfBloulB2wYSYLgZEL1HWljOMvuh0PM
MPYtHVXKY1S9EUeIV6YSnwPCj8yFECt/laaAJfdWHOC3KWu6wBX8iovl1Gb9HCvV
OaMXlMWXtMsOC8uOatPhx0UDfqLrUCz4GXLGjNPA1cOhUhpSIrUzBL9jOCMvyuyF
KtXXD7L0VOjwy/UXh1ZHNzuD7Fn2TuzRmGV4o2h+koS505wqf3Nm0onr5bovcaUa
SKZhXL8uZGdd+Mvs+XduippgiTs9QxsrGv5Sdo+/G0DPpOOnzei/aLVmeCt2Fp6O
bxjjD7+08eqF2GQNjd7fVGwnVnkj3LgWA+sP5FrchEvJDNWsZWrcLLPIkmQlFh2s
Is4q/bN4FVXS0NSMz6nI+duBBu5Qxo2tRsaP0qiutVbDXDe8XIaj/yu0jJdNP/x7
`protect END_PROTECTED
