`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NvEJKYj1dQEL7/0n9nt8G1jZPbDhXnyOiStxIwGs9JiXGu/Vg/YxJjq5k3VZloEM
8wz73NC4TmjUpp3bpXO+/fB7R0hoiPSRkKES+O4sEmq2m3Y80+tn3m8dAQSAmiav
ZqKsQl+PJkG8Wg+G+QbS+3nmhHNdKTDAAyIkeQBiVdZ9nDA5YMaHv4G1/3HC3VCf
jMGELz8wZFTXMSJWRDXeQiXZ6enc+jhIJVfM+9XduFcg1hTYgzbPhZrASacI/4xw
+N9JG041pvg443IRxI+yWM+pw8XNc5+0OG7viyHlGqC3lUFFKyrbhkb41ahzL6mF
IoMo6pIkaedJSryjGLwh0LScGRrxBKSX25ivF+mupbEW2xFrBW3SGIBimIw4FE5w
nCaH+KewzAyNkYHb6f14SEIJe0GaALDo1CTSr7cvx30+u7IvxePMVPfVdnOObzhH
q6UuIdwDCk02lgKLIXHiBVvXxUXmjd4cEfmW6VRXlrZy54Kg0ttWFzrd4cx42U6X
YC/vJ/gkh52U3jmVFybKIjEZoGqGU4xARSaixmTn70Fq3h5LMJGeG+S50ZeARK0h
dVYnIkx5kg/yLoHyuuySF73tBa/P60wOymSDPxFGb7r0pU1PK9kIvrpZwVnKM67D
tBgaxKbbjpkKf/ZsrUUi0gAziQWnXuciY1kRVqE6ubHMwqh7bgeSlC6AP3Mjk3jb
330XlAdMIOndcMNULlguvXSGli/ex5dZComHNuMiEUL3+6tbQdWKJBIoU5vJd0mY
XOS4+iTumGQsdhwPSRcDtX8A/cxjziQHPsa+P/tcbJajUbtdFPMx2ObQ6ecZTuLQ
gdXXMxWABz/wXOpOwektTJE19uKhz/h3dy5tp5bxq7+ugu1hZGJDOuhDaPkQjCu3
9aBz36372Op9Sb9zaB6/TCr0Bwcm136tua9Jhi8LoXIIWavUxgjM2MDyul+WQ1Kz
Uulle00QE/FrNKPyfH4lkBwLYSf2NncIXoYgX6nVs+Khv8l2MwiDp6sys1rDT7hW
ImV5Ppg47i/GTg/j/rNKhv8CkETunvRKLbCK/kYlObuVdL4C1r8tmLlRHfrosNOt
4f1dCPTut+ku0BXCKDNIKRIMHA9rq/y1scxY5zjXuGBDHaBKzEaA9IBltqf7LIPP
c8tYMALG//MwkYUN3ZrA+LxfbibuZDNNFGO4ELT8JbUDORfdg5+MYFc0XCHD3bbF
Mxy9ONEJlYiLs6daq/JvvoBPbt9Yc70vd+UlLvA6uGvZqsuVmTLsYuIgRoUusZoQ
bJthro9hZ4ey4K67hu6TKtdyl8c0KUhk2Y35YcCV0UI07rTmaE7IbwhY64EptSiN
cT2L5qPjQn6WlCM5JD1BhmXaVv4PMm97mjHV2qdGahhowh52/x8ucV3nmluzOaha
ohwXdNyBujFrE1Mlhb7DqUSDnIzE5LGjSs4PFRnWhi+EH7QMum7nm87f47QZhX/R
uBO64oYGOLgvfMv/LVPCflt36DHgTz5rQ42TxMhtA554dwXQk7U6a0sHpipdVON6
wRALfNIjtOooHpYlXVZmltLrYUGmGeNH4b6VMmmbZeAc3YfH0+VDO/fArBDLv+Of
Q0qQGuzCiNWY2UjvgWp8MhTN1GmXJPoHf0Qf7ivJI13D1wuLdoRWBQ9nrkLAq787
bJ9bfs+RO/ssfr9dta9U295wz0ElK9eVP+I5F0SLTuVAZW2i9PICa+Rr8a+UgiGe
ELbql8drQvjTX1KAr6k7wvFwnkaFwFtMfGJAMFFT3tiYpbEnLX9bkYAE7Hmo5leC
XwppfM5rUFc+qjlipLWnSYxwCl88DX58894Bx+ZtEWhAvKtXaF+j/yrGmpxGpjvu
6VaeBXPIIh3Yyrce/QlxyutA6Cm50Q9PVNh/T6Ga4n64Fp3WI4FIwHB6YhUFh8Pt
JgvSKnMitTfAMKhf8Cd/n5D+Lf5rizd/mKAFiSlPeU0=
`protect END_PROTECTED
