`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cfbggtJaiCOm+/HXPCH6MxLqHwUdqBfUIlEY2yYkFfTsZj9Kfivu4gZt0pfA5muL
dpdmKBDyxasFL1qSK0e0+WQaHtmb6eByfndV2sTDNoWQCiADnP/7iqFKlObIV27w
1jQm4Bgfo5gRGvfTAudDsBgLSNuD6wiV4m1LuHfqwVff52w6rf1iEhH2L/iZs07y
LqmI4fIbDN7+Ho3sLNLpl1rIanxxGjdlbIT8yeMMetpCYJtdfMI38dqrXsIPWpcI
rL0Um569TozajNJD5z4YMXTfkh9qehifdFYNmuSsuak2JNjAHk+VgPuoqw5zvNCC
QC/tIt0d5oOfmROjq3J2r4bPaLBZfVBTy6mzeM3HOEuWNwNAC/RVzs3hIV7aWzkc
v8Z8L9W4l7iSIREtUszEB7GXAqG7Ja3uIW5jEL0AeQskbBdKOywWLYf7N+qw6v45
faoZnBpGbd2i6UB8TALRyseBeC6TXadk0/EyZNz4Qfl9EMVa4f1m7QuSx1W3i8D2
kJuDjBHNmYy4EOPDA7s0HqTLe7Q+4/Kx4u32rqe9doBLszW8sAWlI59J7q5ud8lL
MZ/VIoH1Kedip0U0h+eugDY2yCklyIB7gtg7GLjh+DjJpA0+YgnJCEYRILWhWO0e
Y0obbeQfBr8EQh1dU4b16Jl7ILOyFY3KI5gNw1+lF+6EVAwh2ncfKH2hsZTBVxuw
pOjtgNr0jCCqn4Gh7mqrHWfirT5cVP4GHtZ+gN3mTbFSV+ko7cVYwfJuRfHDxump
07Y7DERF3PbeB7BtWRCiS4PojagVcjqxKVs3rTcfJeuxPepu0m/JrCd0YhfKy8nU
0obP2GFM0fBlcJw0Udvw0tak/5JbKKVS84Gq+409QEfClvwpyy1aS9BAg4p4XOjf
5K34r5oBJzlUAGNRHxjqdDL2HJm0rOmMhNEZBdzmtl7nHLxSdbqPWGT2WVHa3Fmw
J67newhtp2VkaKQQQw9fJiRkf3R6LeowcoC/h37shxy2uM76HAH+ftDGLZxGbrIj
0ltX97U4JbPDaVVqqs76ajdL3z99vaHacJB7n3y1kWMQBUTg9UFY48VZsTGY6mLT
JhuYDLE7zuiJZls69EoIEydgnU5Mgu4W+S+7QDThORGhR5HRcWhZpVTIMlQ14d2B
kRlu8mroksrF162rFxL04CsEPrtAN4iYbUsyJVD6ae+6XPP6y1Qiwb+fW/elwtNa
EjO1czSSKRqyjpowxKC5zvIAmcW1yVFWH/amW7W6qWcNSVWoWJr1zkfdQy/7R80U
8hAvfUclzw+A4ZhtVT61kniqslvwplancOaaJRm7lObnauJpLVIXR3fFsq+7Y8Vf
V7vJXil2CovxXnfGTytJwxoF5N0ntXZstZS0XOkQ5iYX1lbU2i9xIHxHvuWawb+U
qnoyexjbPBZuN7N1me3uy8u+wIEEyoTiHh2XGSoOvDJEpuD4kxLi+YLAPgK3VJiE
e0bmSc1Abov6bD8ywWaNuASafM2YBGZrkaTRj00X1oK8BCpLLuXqHD4oE8TB8EP7
8KxyH94wDyY13gnzsPmKceREhtjVAF+n4LSeJmcs6n6P2myxdLcLt4QfxiNFHjnJ
K30NEjattcnAnBq/fTLY/EGYHc0OL1/ciITUb38Okadj9mOR6FGgTK4R/egcqnLq
YcdQO2rk4eV+thHPghE5aFIcs0w3/Hae7Ctay0X7W80GqMNmECe8zSPtfKAGiMqM
UcEuDSMyc2g7A5rcDzrT+VP/lze5o3kCi/jQv1e8FVAVStXbZRVOlIKcrlZpmI0E
NhhSAyO7a8sGX/tZwmeJLYPhyGbyizPMFj+tlQeT0DV1P6tFOnlHEAf/ofwG6/Hi
IO0egW2knvpvz5XopNv8Nm1BfUnEBZT5ZI5DKV7k0kSukRcFu6/kaUd1Z1Q5jFaB
TWI4tXH50aaBl1OC9ojIIw5XcTabrGZh4szl0/eQtEVE44GnUWZhnLI2Tgcfrp71
H1jImWmITjK+V1rALRJBQIyUBGYIi3UNwH9/TQklU/E4L0XiEaOlNyXzpJjvjTSf
B4FtiWUCu4iZaukNPurhotDrimq/FPhP/pn2HDQoHIvTl4Rlsy8ywjFyggLpsQQG
/YXx1fPBq7YrlNl6MnJt9/LPGugF+BO3KBR5hIqAn7sofT9WiQGZn6SQcRkaPtQD
DVZujzpBULNWzJgrrmPSHft7gQv6DCshSJa2tiqybixWTalYTdc2A/hSpqjn2JFW
pMJ7VKG6IxDTyqgSfZcRqfU00UQQtsstvP4+rEVUWz7TNg01m7K/Muo8VgqFHaPZ
CCN/eFy5nM5wFOXn7iJU9UaJVT/xVDVZp1Aars8t949ZOe/Y607KZqrepJvcAFIm
a5ScxALa7fTGWXmlJoORx+BtvScCdWQmOqsyWmayd1rtHdS1DsLhjfT5sMnnZ0ps
l/7SbO+SQyrLucJac0Mxv27zKoFrMybQfaZK4cRs3/B3I65c3OIhr1IQcMKtGjGH
dlcMK/E7e1SnzwConyxZcrlCW7g3yvL3jYkfDRvOxZemi2gTaQwWxUsc6/emz4BE
7nH7pHqGU6Xi0Uk8APyUHEJ4by4o35s64r2L7MO8JHYZzUdtb7Fen8vAiKYqTI2n
hQlt9LX5PhBnKc3z4A0//ZhkTPkeNBo7JlhF99hHdg9gvxfC3cgVyZ/4FVeE4OJb
P6zZRHgeHGF/DOW0gOmnM3Ni7eE05KOehjHuk3XzU6nCUC5lRshbDYejQuHDo9RH
WqioTye6gAu8MkDnHi/X0Oaj5gSAn7dHoW2g7PVNS9LRi0cOpU2ZTD0aAkn8g2fS
UwK0G3vbYTg2G3m7wASmepZxINEIJ7Sf6y+QlMMScamxiv5cmwwch81OCyqKppid
U453OFUvb+gJepDjoYa3h7yjsP3Jz4RSvaHC9G0lUbWZHrDlgypFSHDHkddL60ug
pdp8sgp9DXzzhkjb0ADxfJjYG8SBWunJfHd8lOBg0JE=
`protect END_PROTECTED
