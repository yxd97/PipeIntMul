`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pMOXcHW+H/310sDGd+gDeFvo2YjYn29MyuIDPRvAZK69Nxxvg0Rp5ebQ4o040IFE
dyireLvjRu5vGhjT6lPGfqKZs84o34fy97x/+HU+fuiWzC1Z+/M8a3iEZlnvU/4G
eD8khAFiMeTGhbT78299a+m5dVmiVEV9dEyt37/xtPZHh0xw0hu5BqTHr6bh7JP7
SqfbKc/YyP3+UegMcvp1GjXap0hG8yuK4PAwwoHW4Yser5kvDqgj86TVpgrTXVWk
I/MLEjO6qChqqgky1oq/8yNadk5YBLRdK942hDJH+OMkIkzjXWlfT8dOJuG5mCjk
8oUgs+pVclP/mr4rk+w9FzVTjF9UVmwD5cy9sNltGqhdWRpgvxt55qLXGeU/QIA9
1CWQ0lq8yoVXttKzWdgd8LWKGM3TJhyDKSy9IN9wAQQTxO64/DFUA1y9b2LuyY0b
E3Zfjz9Y+AIeeh8BNz6gVsuxZ2sLi41Zp3v/KM57gOitNb0znGW08fwFrnrhQaug
1goPyE2i55oZTvYoU3bbrZ3SsvqCCZZnc6V5FnzwrBxEw6dtb/WuFWJHI4bLyciE
5HtLTMDNrFtDthC0Taqm2aKMCDnRl90egE6ln2CEoXowUWjbjlMMI1lCpyfdy8ZX
IK4WY/ZjG25PZb+DkwPChsFbFSIfe+j1x0VgTMqzGdS1IXTEVGNsBZUuJqZuxg7T
AuBJblBtd+GbT0w17/h9rYzGe9b+dLqxsh7olg1hXM8rQGXTAhzds5HPi26GPgoz
5/c1QEq9ol0LqSTjuFHE8nQQrXHUB0LTZ019tKDba+UZdu3SwmU3SC8JkkDQiesM
MwZXF+KjP1xubge0Dd8/PsNJrdlakLUOfETzGtwTFhzIt6BC2Qa0Fn2A7v1/g+eu
Jz+a8vYREFpEUAB4gMlmSkNKcuvXo0jl5nMdtgtfQ+uIWQ4lmrMUBp5IRVraIBEz
x855xlp/AEuTX+CZORyQjjWTW70qHLrknRnJ4Wn4TCNlb+kKNVu5JMiAYdWxH9xf
N1sGPJi8luMLsMqx5wi+g+aYPk7KpDp8yAdzlurYkB0X/2iYiJmFNmYjiQ5PGtvr
S1KlyvTE3WvUTy4Aca9BTwsSM7gyyONtwaB3vyEtDCkJ5MqOifkftKABsCFqdhSu
nLPuvqItrVBgCInJWkoaWCz/6SHQgWhd4Sj4ptTsPSgtUdaGz3YbBgZY8ojRXCzo
7fqw1kDxAjxZFKfjgO1teu3sXx0SIFj7o59VTIkmQV5O/N9XVGj6ByGotZUa+dpt
TM6ev9AQSbOMpqSTguRlGwRY4cOfsoEhjtq7ZVt/EQKnQr8rMsW2I+Wie3bSSF3B
IKX3MbrMk2fY0sp8KVIFILYAIw2KGZWC9TA8CuIi2lIdALlu1lzTf5Hpa4oyYRkj
2KDnK5dnDHFq9VLiDzhI3cOcGzVspRx54Ls6EZhEofvSzSNarBZ9DSd6vjRSdKNw
L0KjVwiDHIfpDsYIbFBvwt33Q7NRwPND6R3Mj2Gi6i/CrYDArhqAQ36o72x8ysTe
NP5q+d/iPJarXfjBtezT7RvTD2nq8Q9XHJ90+vkVJHcdCMcxL+zhZAteMw9si7pU
ZF/qL8odWDLKcOTI4/hFCsz3FkKxr1igWdLqFjEhQgZ1zW1spaxJeDMaC3IJCf6E
41kppBrQVkVej+vVh9ZXdkVRUELQRw9/17LCUhGw499moDcBhx0zHxiYHTTwvG69
7Z3Fo152w1aD3cyQW/inYDGEyOsgAzMR9iOhXvc3GIOPX9jGQjHv8wa1UL8uWb4l
DWdA/XK0n89TS4iKuCDmRLLAL5AymCGrfr33piEoRq8JQQGipNkwCnJrE0zzNzIL
i7AvSqBD6SPjFaHjHTamDagNJbIISz+bQpfgwIj/VbWDdXa5XZEkgwUREEjfehw3
EU2qbStvCc1C8i6I4fy20srppiJKBA9FFE3nNV/Ix4bvUg43NjJH/+7mHqKhcceu
hoVOIOd93L3m2xsvSKTsZCl+5sPyOIAtTLucEA4Ryj29u0qtoB/RjbyYPdmgsit4
JdSaZ9c7M1y0+tB5d3w2zRDAHDW9+wUb5ChRxezk7VBL0N1rGyXyIRzo3/MwtRyN
iwm0cmUJ/PaVR3iOs+xngp8XhGMUgGdDsjKDFZVO1MzNsA0kO4D4NaQZF40bPziB
cRuVDuH3JHK++vnopVbO+exT7xQO3NOw9JvAR7ktHz7okTE0d2UYrceejqnS+wcL
m9vbTM3aUG0Hec5C6oyVp6jVGy9hfN5UUGA9z1zn9jKuUMzrQa213Z5Q92edpkjR
JifT+FKOkbSQ8k2xzNMvZsCReuCGhC9JYdFqPjR/imfHmLGB6ejOhWMVeyS4g5f6
Mk6UIrPINoWGU02B5Qmzuh1WFNHxbG7a99bHHD4ZmpJLf1MAo7UlQ4BWEhUg5V7c
uSDn3d4/OH0w/36zDvjoECQ1zkQRm4Iw348WZEkfTLtDkwxKU9MypV8v+5ENl4OI
CN5f1n3shWclI0eTGkF+QMzh55SDBLdPyRUYWiU5perc6zZqmDLJNpIZY/CAMeYJ
zVA7ozAIGGHDLrOSNetEUKBrxoUu5xK2UKVd3mhp53vF8NEsnKpvOE5ysf7nGpNG
vr9sc5/S/DijNGZ5cz5s1ql13uql205OluPq9IHc9p6BBA5Fr8y1oSXyhQdxA7+g
ZUGty6061re0BoaMnES82Lb8cSm7Qpyl1aihhau+761dTOX3796p0OHAVsd0r0Cq
DydYd52khKsXAZ/9I1YHiPox/UWKv5SGpwAbBT8i+HrZcTslLGXT62vbFr9XhM9i
DBhIYKn2OezNtG2Ds//jTJPbP4agqxziIVqoyLLy+aAxWJATgr+vPT8Zsd1zDppG
eDBCXDdgFv5IEQ8q40BeNKgmpaGdFIm7P/O4+u/LzMDn1WZj4TcuoLl1d0Wit/Wt
6yKi31ZI8X/l+88tjTrJS3Yx8etZJw3dXqWp7V7Jyz9QO3sKagUGAwGXUy3IVjhu
CEBbzgKIR1sqeSZR29coGQG/CG0bxYsJqho0lYCN+NZlpc1RYZzOZKmm9ZRbxY6G
Wnh05ulz5ngXoJ4YpP5pvS9nKga8vyhSmLfHTQR6xJMttwsn/wHJAyTmxQRKf4AC
ZajVinyOK8hh/Y+YIJznIWmhmwoqCijRx7VJacw9mJDyfrHv/L+nfnoTH0JWQFfT
yVYl7pmbvTmlsCnbt/+sVuL7t2lyOihx2c0hmlkUyiDJzKm90SGftDhCKhSnssdt
omRoCZVnAwDs3vM86wvQFM5AGaHZh5EP6ZGZXWhtqF4Lg5rYsY3DYADRKuH4ZQlU
fUDBhZfZYKxxL//lEzXjKZg6mIsiQNgtBxWgUPn7LybxK+xnIPCLlLe6YcrzPqN2
hYNV+WXFpyX8NnD9/sTLeQ==
`protect END_PROTECTED
