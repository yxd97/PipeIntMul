`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pLX/+ZpXJ55FKriuuSpGnJ1sx26aYpj8BZhnokIY7a3Jw6iY9DgFqqDd1GqMjn3x
ynslWiFcPvn5pitco4t8e/NE1kbOiatWC8pKXIPHmzmBr9EFRGmYVNqqRLC8jTWo
zO0G+PsVQi+7ohfw8aUWOf0mMQ3LWRMO6h1wArojHbZzxYn/6qNrl+mRkcqlLADI
2g6FVzMN/Ppmpy3HpsPHNIYw1fAiLZcOVSbFrwqYxzfClMkuJc67K2e7Sp9JuUAC
ERhtYvYTn2I7YNvOoUVtBjf5P1XsEQN1T2939RZWvyTsoFceyoArZNZzQiw64niG
lTKFa7ilmITN34vIFz5ZlXsdXKVpf1AoBvKq0cCZh1CAOj4eB3y/nUoJ2j66WMb0
0oko3Oan2Gri62bbc2nK3zsEVcPQd3vj46dswVt7wtdpfiruxbgABgJzF4jiI/V1
3pd3kfXsep9quU8YvtniFHnyAui7IX9rvPJTjKrxNYb2ZXGXfINgshnv7o8JX2Rz
dCoIeWxuJtIIYZNTMAH4GasxIDB3YRNjiTxg7Zy953EuXiOLzgbbG5HSBDbwduXl
fbyBx8QwkTmgWlFHO9AsilSx185uk5cLqyJGSnof+N8tD+ypkmwE//Zqu40LaMBf
h+lZLFcUY/CqMpKMWXLXHuWhEZFu+Ha3/6KeP0uS4rLVPayCTmhrZPCocFimwT6C
PZ8esz40lelNrxy63Mc92YNIX/BmJGsWZfO8duvDpYbzroNm/IlzKLANlTRNmIwI
a3GKRIyO5GR6UI3zBsGSGy38P72An+xbc7IKkQxQOuJ/apniQNshvITplztSskp0
z2bQLDYkhdS4OvJU+P5JKQc1fdzLriuDtXRoBQne5ATu767Cy1tx1+eKVIMMYRpZ
39xQOP1FpZn9wbsI21IVT44PF9t9pBPSUSp9YHv7LmHj9BM2Q2isAgtxzHKcCCBH
RXYXhcHBNFOv+n5FoiE7qEFZ3MSVAegrtbbfemmb3XbkTHIqgI5Iqga21o1ASOiJ
GfnOt3oZAPehbzmGQnGJrrzUGOaI+loFtd0dPXLh1GE76LSpOWgF+Oh8vr2BS5gu
/MoUFac3t6sTl/Zv/a3LUkZWfC/8Yag9mArqlj9FOAKzpjbbZPLVBrBfyBcxqjvc
OFTMM8j2TjthiqUOPcr/+3//WbkaYOPDpC02wBr9AJGPX6twvPBJ97Rf/V0DAqwZ
eW8F8nOI7Azva4vPDhYL1JfPmkmNIZDY7jcCedWniGfYhsoqTf0i9zx+oAkgsDRK
yG+dX8Xxve+962Z8BpxeWbHnKA51sE9vkPvo16M7WJEeDOy3tZJ4RasHxJ9zoudi
ipPLEm5+IptIaigrL/azBchI68XvMtGIgaPUtUaKlppVbTDJNhTyJmvRhg5Xp133
ZkW71rPEZiH5s2MJCDb5jOTkRStq7nTYtOYO85IlDa3e4wQtkzscr9B4fMK40/Vj
2gV4GwkoQ6L7j/GNTUGtu93k1Xqs+I7xZqdUR7kmygLU+ETcCtYiJvotedFOiJxf
t5kwQP7N6mnRr7c+t5s75tL0rew1DKfpvN3kxwP3W+Yk5axJy4NkmTipcophY8LZ
cv5ofoJhQAoHpuQM9rXli79l1DykJdhmziTD5riOkzkkX0DOr7CX5CuyX/hwxKGa
vcvEoEawU+mp8lpY7+7JkozxTY7eep34PE1vMv+BTDHUx9XEvyJFspxb4GeHC/S2
j1sCNf0U12VLns5NYiIlw89rtSZ4pUToTMr7DWv13isjJzn59EiEBHdL2Ebi5+Qd
oVyu70LnaSfAAGHofaVNpf38KHeXFZS9PppnMrzZGyiHBqN8SD8YNNHgPE3W4rhK
8zAcAzycWWVNxBU/jKanOC4zGyeq0v2nmLycRP+lwMIZuZw60OdA7ndOHHv1gZ3f
hk+daxLKOdkYUkvlryFGvvNMk+dY74Qp+3/ULJTZ99aXkmR+dbWlwD8k6E/HBGLv
ilWX/yVovvYShzyzyS9nYw/xDtMmE7uB2E3ayxuCce/gHJiPAXi06rH1g8RFiwCK
IIFYW39+sBTRC4iP2iYNoCxcmrnXjHpXRqWJmdX0C1S9FVlLUiR482TfhRXv8HQ1
Qj34Z9wZwb2x8ayvMOF7Z/agOrjy3MJTx30NlVvbxJVRpfbBa+Fj3kevDlcYOss+
/q+lbEwic2yDF48Tg6Max5lJMRYAV2Iyvk2FwMURGrhVSmtwfeeCX0x8T5QPazAy
BUHzr215fiNaB7oP+E/HsEW2lLwm93asUzQP7ex9v4IpeqOSrKnNCyV64f+7idnC
5NQmSA5AaWjBxvE5G1IpaWiRMu+8hgPww9XbkTL/vr8uRptjpabSiXksDmAYR9WQ
JuXUpCGPEtbYdlAQf4L1n4+H83OfV4tHvZSFCpKHkagm46f36FnLOfSnBbkeRsAT
GmE96uWYniYWaY5MwlqWKWeKlM4F9BuBUR92W1onhezVyum/mQeS8l69p9e2LASm
4Cv+Yg4bls23b7w7km6lif/S627MEtMGdWpEZZTv4pUnRIY8CCBnj70tOtV97hk5
dI4CTTLM2fqpFjhPmzFixmZao3bGqFaDTMfRF0RdYOroIyKkmdrZ5l5NqPoA1+9l
dEJX+S0mf+FUA4vI3aEGC1ClXALDBnuvyYOSMmhfLZ1bETzj1FucGNRvwCh3utvf
PkFZyTtcnZZHvyh1lhZT8O626kZvoFwZnfhB4esqIfDvfP+Rye9MzxN3dpTm1aGG
YUWRgpFxxfMq9z1RxLpRtVah0syQRm3avDlUF1tuTcTPdWNLupZtynOFULZNJKOD
LTGBY1n3RdhbX7qgiFH1KHWTWFS1auJC8uitwVklDpuxfNOO+51lZ0L7l7VU0/yU
co3cbXo3tFFxnaFHbaTM00doTvnWOCd1IsKBVfJfQK1b6Yn+RyZIkcO+BO5EE0j5
f27H1UoukKro2Zk6IiXgyQBFMV7UMxHwBXiUxceqsLehFcRCyEHSOPp/dnXmd4Mk
YRwl/zd8B1paLfQOKPqHpODefo8bDXXqPNM7lxV+WaIDaRv2v5rRpoi79uRGTLFP
DgTb1kigsDoID6dSW/kLqAKfMCyqHHhWIXA5ooaPiokBg5c6mm1iCoQdw7RNQ3dJ
vPxkoQzqOtlE6Dq0ykS2evbMeNzFDjRzTKegF+MSXpA1vTuhXNpYYlsrZ+nTir6s
tuz3OABHOuyLJ6rq7cnwvURl/pGA23IieO3vk2YmvMLernp+r6e2NNKH/4R53FFW
81g3048XfQD7Cfe0QORJ/1Dp5PE8bnXjdSDT5Yh6wE/PNtZvKqDHzoRgHI8sIFQA
bfMh+j+HL5oOSfK+MoYbQ/b1on+UyZPDNXZFXN6tLYd2scwg4CV8l1znBYGZ1/uC
CjrHfItnpuAgvAUwoLj3sZig8qieYgmRyGaNWqnp/68Y+Y4yeumDCQoS0agPImnh
DcDHXVSrx0JXu6vYJ8yQ5+a1IAeB4rN4F752Q9rf0RtrOV6UxfbZCEoy/PZ64xcD
ENJJXc889hWVZ3T1t69eL+8g0eyFkaYcZcUOb/Wirk++ERO1SO/ooniRH79IO61o
s5IcOucbV4QrmTREgToZJBgbW13A0XPSmKsFA+/9kNyGY8PfElno9vLbdGD/MQJm
FXUAVz57hg+NRhh/T6BVlEWoKSFJ3bcxDU2FaaJWP0FNxBU1cA305nHasKUBnp8t
O0kJLvDE9Ko2+UVX19XXtg++ncmb5J0FywQ+kxWGAhINhuFm5cEWTY5f8LGaNG4W
KTdCjCHolo2MQh0W/sDBpPRijTpwlPBS6oGyLfPHYYnvyRkzBZ8LezNwGKgoc32c
aNMaqSDqJM4U9KJH1LisP6ORToNhb1nKVTPNQlxSb4LAhFv/cY/9ctvSG4fPUTIH
5cdRIdqEqHURccqnS3wMAzSk/xIrMTBhejauoKTcLNZJUCilSYvSHG7kMg54FSsK
pZkiRQIJg9xfyB15uqfda/LOuPEl/VRmAtjiIMkAkYf7F0cn0YClLKAzuZE6Yi6H
TzNzm53PbRshrTIaD3X51hj8MNrrbg800S0z3282462LaTRxbK+0Py1vN6++HymO
T6CzG0F04udpI3DOIpKUxrDDHc1aodzd7EbJIxVDRER9BzW5pvNA4do4OF4VTbsq
UWcaneUMr1vD4u/nn8Jtex04wnrNhdlBgsJ9vUDbH9/HgvDYuHNqm4+ZAanEtJGA
ro7zIp3mhS3ZkzOuyr3eYI2piC9Vc1xRliDEojTH6T1aDyswNWbWVYA0atmxgq//
Fq0JMcCD3jNkrkht/wLVqwNiHSVLsajHZ/zufnGwbE0SqJYjIlp3F0b9NVnXEbf1
pJ5A407EQLVLGTVyTEVdgMJWsCXlnq0ynevWZiIuzfBeHD+jX8vdMEPYCcoFKVLa
FHtjCWKqD/efMhvmRb/euEmNWn8WTlENoNq+XhPV2KT7YbtyiGHtCRVGXo7p995U
bnsScV/oWxN4/H+X7TU9AfgqJCERQ9+N0EBBeVHhlYVQx4+KIlyA+UHecnUQ/vUD
Nk+7ksu9IRvp8Qt+pn/9ZZmCrH03wsab8iGpdmoavuXSnwFaIs+njgcKcvwT0b/1
QuX4MI0jGjdpb0SK3U2CLNlxlXPtj8UKJ4UzNl4a92ZULvx/829wDqlm+yeu0waI
HBCKRWPJL73BdZK0vBBoR2bRgouilAwsDYYbdoMD6prstpVo2bz7HKLqiVBumh1W
lZPv9rS2RNUqKHg0uWZT2jOR7ZSG3mIlY0V5alzyrF8HlgZ5L4ZHcUabrDdGpUde
i1nTzEYwYtR1UPUmbQJyFPA0tJLCG1hLMDTmSNxWO8cCos0SPPzoE2fLdcTGXoiP
c69FlYgWvnGvRc61p2eQkL9Kt60FY5XKGqBiKE2/7cSLAajh4cnkJhO07vrx+KP+
ldScBBR9d56qQEkNumahRncW0GCr4HzX0aQ0UVLVF2lzjqK1sLOIqPyRtKg38GT7
IRKso1DmShe1ynlcUdymqVNRY/lLNBI04aald2FQfCjLrctX+5fLCtNIQlLiwF5R
D+Qel/V1Nu+BAECxHig9CzjmqX5c2ZdecSS/tMZ9GC9WArHX5A/JM8WR2aKXkTcg
uutAMR/Su1UFBOf7ztjJa4wUz0XgMvDYUNVptbEVv5YAtjFXPqj1lXY/ecumAVgH
87kGtSUGB4TU5zsD6QacPw7h9cbzyDRbPBNpA5b2+Z9i6HyhxGd2GBlbeB5NcpN0
24JNJd43MS/JHySsC+vU7ABvKvqOXe+q6sGGpo5HUplZE5PtjOsn3stg92iCrMrx
l7dPSocQKiff7DW4q+6AfnE0cQ5RmrRA5mEmT54xKH2tTajWKRRAeAt6Mo8EK6BD
i/jWxcZPw2lF3GOeluFlLHag9BMTa/EPiWbsrRWGIGtD9uJuvdPBEFieNgWUDuOn
mORtF7EhXNrA+vBvknUa4UwPTIas/ejsDzF+3dZXY5MNY4BadccMHC1ETIEzniRm
Dn4KtK/gpunzbfIUvjYT51KJGpHsYSwByw1hyp0uneeZT5HOSlS08DRPNp/DU+pS
17E3HK5IaNqdT5GyTYa+c1Jfn7hHAIc5CfQMKKWxtN0t3UDbE0rELFk9Eg5khjf6
zccnl2B0atmGEiuUpfW84k13tNdoq9xINRmiUz1hAWv/t6w98kaEWG1X85yvVQ+n
17Pb3+M93QAy+wMtPTgv0EZvkvM9Mc42NBdy0BACh/l6qVzx2rMlRefaRnV/txlB
vaHzKj22SWfGlbFVALQ1U7ccDuGhsriVYRnttDGlrFvohJbwbUxiK0KlAJ5SCO9B
hlYP+TyzPEXfyqnUNTlSqJI5qp+MWvbRTsGc+PBplt2syzVEix9B33PsKHCe7R64
ScyWZDQ4UHd9ZWvHqRVsF1VgzjHXcXQdyHjJagIS3bcNA6IWAoX6iO64S1ThGve6
L8kIdXNtHg87I3WXbb+gHUBC469nE/Xb00OiqEKPM972BLmmsj96TzdC/hIfy9Jz
PUBMrMZlYlfKVonpGax6bRfedp5qudNooPgGWSTKvlaKMaGbV/PENhqxa1NkVIGp
OJz3uet/zR0rmt3Sv7260q6JroFMNl7GnnZy97C0c5WygdPd2y3OY+vkrg0tQAm+
LnTkw25KYxsBN87sdae8UNjZ+qbdhk0ZQmnabxV3ur4ljZsEpj0C9ERlAfYfep9q
0iFqFZXnbGB8gMCoovuGVxnN30eNi18sl+rAbluWwaKRf/8XKq8Mffi07WMbl0U0
apRnW8382rgtDUtYfARGJrsUWSNJBg7twv7v9985hgUTA3OOkCSKmfRoyvNhw2ib
3d0TpMV4Pfj3ygPiJ/JFU2FLr4yn8U1fCe565JYBUtOkkUbp7uPhtvBxhel3V1lI
CVHFmorN1TKWVQlEIMx3SAwJL1Ra4CDoTk3oLVGbZFKodnJ2DvxanqIgYrCbkvgq
Gh+8Rc/F0KHtQ49OzrX9aTtMG00wo2HraY8Pj1SpVCu6ceb/oM336QJrFOMQWjDw
MGBpE3YER4JODboksZIkd6dv4BElyh1Goe6fB1+26y0P/729qgb4Wtci+XcNEnqz
5KR1TuA3d1IkJ65RsUoFoy+KOQYhXFtJX6CvdxFU0jQ5ySX4W4mAb0WGsg1PX9ax
4SBHF5h/JbPERpFo0IHtcGyQMGEuVUuoMzexPvLbeWWiYhXdMZK9nSw8AcgeVzxP
/LRllUpOj7P/pEEEJTqnt0fgyYWe1NwcJ9Vp30XkjbkloUav/IP3MvvfICqGadOj
z21DXvSUx6IPQlHNvtFdi5Rvf/y6ZjtaCjG0oH6eGVlCwyaPvW/PZlHJ6Vfdy0Dk
3dCsUjrRQND6N5odkznwuw+7CE8Fr8nkYLiIYOX7H4+A70N/9GRsGjaScHIoMtph
y5aVsPX0On/aklKFtC2EVt5TrHzaJWP8cDNFSLHEDEV1DEJ/Wvzi0j4KRhf05zBA
zun9TpvMFXZXSPEv19kCbzVuzK02ZnK4ZdY9rYlgXn1qLaVNykKZGYxtBjC4zEsf
+Krf5EY1m/+YazFneEX7ILRLJfVAq3xkuUlrfIwOogUKZVS4SIoFXnvIzEsUEefQ
ZFwYQMYatw1YzJ8oo2A0PxmkrXaX+kpgv8F2GocoBaex5emva5xJVaoxEMEMBfG+
ieSLUs2pq/odFy9A3RtQ4kuXX9K57NtwPMWq5iYYcJkzohsKIXCi6I4s21fln1Lo
cHbjQBy67aMEHdEI9mTI2s7BmFBo2JtUxPMz6DKOl7exFZ68cSgYIRLDaEDPF4pB
mICYNcT1YEo8pk84Ww6bbf1t7DZ6I+j5ItFMemWc9i+gdtYytKTGauGpezw2fqA8
klKIw1NRUoKjzrnkOHc46Tm+UlvDzGirz9QYNNzkLzbIUNjZ3rIAoiyfZIwc5587
IX97q5iDKxkJoPwV0uy9e/r6bk/tLDZGoE8oLv4y2xZk/r2Jcf10AK7Yph8gsPTj
xG9OPqgfqznVIoc3epx4R1Q3Jn6tmdwRGlkH6e51/417yF5iyPlzyZfcEZ92iDVj
VbW1taqB+pxMosz377WN1lc/tqVKHReICwBg5Keco5/u8EDr5c1+VaD40wT3wjfH
FSnkulM4zdyxBvLbagff4Qiqi0IFtVsy+iJeD1PmzPAhP4hZkG9dOVtbNplfs+BT
imTawk2QVuQ7LEfLsT1tX724uf+Q5we4up08HO0lv+qgvFvWI1rTwXGEhLkPXAJV
FH7R26MsD73CMu1pZWPlK9g3Iq6lUUlEeBoCcjk3cX69kZFQEX1tJJNWyMOf06yL
fCf/C+zCIh7rcn3ELu/fTzDCPUANE+k/t08eeJkTgdy4JgVGXAhsNqiGF99kKvfA
TsthLVEy4oszx63SRqqWw0YNPtstu7c9jnJlHPMTzTnOGwYnRfqcAoC2glzNuo1T
hrOv402SB87vf9jQTvh3/wR5Mm3T+PVzPfwaQm9tIZfAWOO6Ql5lxYresRCG8x1c
Lg1I/N/3t/QOgdPY6H1xTT2lYUoPAPavQi0QwMBpIETX8Me8s6GCP6Etde4WLsM6
NNIA621jh2JLgTZGqPDr6KVZh5q5TCKPIuSXGumf5NtJTl78i3L7ErvGjIgJKzei
DmUKeEfOgoW5MRQLPIGwRvBTJ8Z+IPeX314G4yA476LYQvJGJNrUExsJcYlDY9nz
Rq2NxhTzYE7wtCt7LI090uDaCpp244MiVKyJXImuRyCLNvm/NRFPc15JLN+qdK7b
+dIrwvwjQu46qBtvH+Eko/1Ue8bJmNf3KGF+740QPwD1OpOMA8qCUFg59DyV05XT
aRsWxv5iBY9LQkkXOMuusSsiExOkFGxdkp2Dey2tRfZTfduVfWZ65mYijjUFUh4E
qUOA57htYPYZUFEH23a0WKhQNdrzN1hTbALNbhu7ELZPb65KwH8nRuWPQQcfcb4/
qhVLxvGPnnTF5ge+AHO04RuxZyRS4Xs1DRascSh67NPODVsCh/Z6OVZycqQ3R4oe
OsJKUMB6Ig39tnL1oUlpk/sQfjbquEFnYpO8EUQOQAvfegPm9uqd2rPbBAgZdc24
xRuCRyhSV3OSznZEqxAkhCwARN7GYsXjJhiBKV2juZhHkR1tNxCKFmGYuBJBY2BI
xIQINHiKz1PBqL/78wqFco08dV7BeHEDsZxj2rDi/KNtFz/9TczeIwBLzDY52ck8
wqz/SEtlqjQWH9/Nb4Wk75MO/TocxyTyuDjEiw2nnrhstpgVWYFQ0Cw3gYQSkdoJ
hPqBzzNRRIdRcAerjNGyFiT/zX+DZG7ekEBTekuije0iBeGMVEOOA9bsF0v11sWu
8WTNl8tDw3dKoxCc9tdiSPx7PkrmkoCMGamgSlvH48VKvwV1cur0Ec/XgJv/ntof
OJ+z2aDo7xQjWZVs+z8zHvjALoDt+hQBrayR9TZhx5JPR2RvHyxlxoOu3vEcPlcy
hNLfVti0vMC6T8dgD2Ctr0giuLNFkIePgdB5IyIZGmC6LlM2ICb1pr/mzbBvW0uy
EDaBUWVzb4X9/AgYmsQqaN95qXkJlh3OidIhgizNUpdjk42/prKlvrqrXLJGM8qA
/bmM8yd5vFxKbUE5mN7DHFdWppzq1HErWmjtGMF8XNHm5b3ct75rjh4GwZEqHEkb
rlydK8rDFggvQCIQs87EeZdUUEGEqh3w/L+y+hrTYNMjhU4K7ms1f5bdnACIrzpR
eCCHY1j2GGsw8MXgPeZgRVmKjCtGhQf6D0clzMrDwsmC7alHL8riABrYhspBJjnh
caXD7Z7JKEVxAl6Tsu4W+pGjmmi37RQaqkXHOR2bpj+5EK7zGd6iL3FWK+U1B4rF
tbqMQT9tePHuNvmjJfmX4fMdDo9T3AeEEWz8wY/Vvwq7SPxNxq2dbHxveGlXDhj3
6JerGKpt3Nbrk1UrQTTOm23nD+BusqebzvNWKqvzPigTUY5jVmXmp07eOVwuk2+q
/meVzSEJsr9rpVt+qMWvypNmssnsZcFqkCF9DSdCY9CiDhRx6eVI4fk6kIDDJtN7
pjKWFD4zmSsNOmCGdknRPPWbzmR1wvTLGUZ5BYryu57o2IYIJkGx1IrHpajBlgEB
CTgRIVFkQlQ1XVwdkKAXHwMisnhn/1vfcLxcm4O8Pz0IFfucHy28Pltrm4pc5oSu
bJagH/WDv0oEz8PKId1ot6zkGIv8xLcaCkVsPcwcQrBtJYSj2AIJlVzWZLhTk86v
t+bX2bDbn0rxrZbz1Nq3PzaGwtqR9dExNNioCFpH/T66uO7zWkhMm/7wJD2ZjruD
a7Eb0Rf1G+6EIl+g90CnozWJk+7JtSFogMvhS+KrSYlV+CMXIdUT44Q7ryvFrwJu
nKca4zBIw7f97C1T7UAqIGcSZJqdQRRHsVQD3jmhWj0nzl+3puWf1Zp01egaXw82
7TKAgE1VnsZkBjvB4lZC/26K6W7yvm1uwxQDXFjXgJxPL5Vd9JFFHgSzxOrA3+QB
JZtIjk+yxpgWPnPxwDxEGR2Y6HBxAAyj0FcOJetmKSM/SXVtwoHSbCZ8Qm4I4oND
/JZciuUvr5k0QwcQaiVoEMT9YGujUim7LZd9qgDcYCtRHrRPTG7nDPO9eYOKbKf4
No+gVAx1si45ChC8jgaGuw==
`protect END_PROTECTED
