`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BWboeUgF7v3juGeFUIJ25EmVavryzhK2/HYQXMLb4jR8CiHW9f0DbuqDL/ImdG8z
9gg/EtpE6ZGvJfYxB4V+K3j386dWUI2FBnl7YHugtTuP90i/LZiyBWwLgkkjoyEz
fIwocBrXQrjcNPTKJfJgsnMawvCJ9TwFd4TrfeXmVqOtf5ZeL5X0lxygtgOTzTB0
zAeIRhnD+WW4tIWIRcPDfK+O0hr3C47lkLcAYDFElN8YiwHAnyEMVbeByQFMcJiT
liH70MlpxRtd+f2nh0Kcakyy9By9fTvHUd+DiZIF8rS3ECFMGRb9GWw8sbKWyOpH
rzHiOISdQS6yvTKdjk8ybL+15dO6Mhdz9fEvv/N+ZSfNgjHpNP1FACFLrb8mOj1L
d5qSca06O4Ol5EYVStEIcCE7vgYprkrztSzzlN6uZ0VPEoQ3uxdjjGFicDfY6FlS
LWmmiIejEvb7LHz2KBbp3LuGdl+mUsaxk191iFNdj5qRdE/dCmnaGqVC/iJdKpcV
4HQ+00lIcFnVFI0PJm7oe1Stp5KhFOit+UYTlk5WzIxtlAGIB5qONsMtem2YKWAz
Dhsbfud+ClBXXdEPMyBp7eSrLxsEW1UzDp8NfPH3sN0+zlvrjZ3Pgpgttoftd2gT
DR+fpuXNIdkgZklC8yL/1H1Q/6Guo+rCIhzdYK/H1/5cXR9LaQYtPy92aOEbFjYI
W1e26OoT5ByYytjoA72PxlwUAaAP5HRLFRP62QdIP4W95g/975/pRck5d3T+ncIU
`protect END_PROTECTED
