`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BwJDhOfd8uDb7vbW9g6f7Q4f8jBltjBkYGN3LR/i3cxgUvL/A6O9+33tKzRI9eES
28RhdTZt7qksSuGzTwuJTPYUXLn1MDUB8EFJg85oQURFMhXi/UMys9t7LNA6t0s2
m+UPpxi/kKQITs6eAKWhFAmoJpER1X5qTEr/BUb8JwBMs/CegPw+jC7iNS40op5S
8YsLFw0aFI6aLF6MTeq9789N6fZC1IIuiZLB5Rqgj6o+gmipji5akAfclxGUUDmw
XDJSET3VKjgvUTtU/mRHJbkFWZr2k2Wq8rSsxgovfyg=
`protect END_PROTECTED
