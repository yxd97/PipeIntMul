`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vqfsy5pFA1d+MhS89YDrHS3vjGPi1WPj5NGWl70wCQdbdCdRP9cHdx4wRSr5IjTW
BxLqxEq/Zrlo+fRgL2DwSSfEejY1AXttKDTUKMyeh6z3CItwDIG/+a91wUTUA3c1
fr1+MONde8sfwKAJzndOeaWuwRinjmOSFCZ6RQLTYfA3KA159fnBiFzrRw6vdjLZ
T6XqcH7VmUKI+wAtPPYCsE4l/ZYwKrydUEXyrXZYaa8LUgkw1tlZCV8vjP8Bvv5Y
svjo+3JonP6YPVtsdejmqRMN8FIuNa1FnVN1b/4xGgdc/9KwAfsYSHN+L9/qCrEI
XbAzwjdV2bgrctOL7EfAw46iBL9gHZ3/VVJF2983rX5wF5UkUFTzxiX6uH6QMjL/
2XvEZQV6LDzhjy00OM5h/+pOaIpw4fuSLz8pZ6bKBouMyGsxC8XeTPYrhQWvp/G+
6j+4z7mjMj60dP/zIu4hQDdzy5ztY2RCO9jbsYiOhzsMZg6d5p5ujbOGjdDVXSPP
59E2QAsVAU0SwSgfl+22QDaybf0DwdFkCko+G+wDx7TONqm/VhI6dhdBhkA+7TPI
XIyNPhxDrqc77GBTbX4fAvya67FfIbEqUZzm6Eu+teibEzpHdb9mxB1dhqltaxY7
ot2mF/lh23MxS+OVbbmWpBao0Bx8kselN1gpyvDxiTmB5JlEy+Q0h9g9Nrok3xFp
2HH144qid3PCgXgwuETCwKjhXeDkQUA1PUey9T3T+8Mrj0A6te4zaV5MRS4XeOhl
JYCN497dPZVJJ33Qejj1tMb76vWcN4ZMRrJ9Nyn4IjnHCzVspjE6ETndhZmR0cqa
FVBeev+IqEsLt/Ijr4POaNDaSWsS/B7+YmqTIlUvj6CmR2GLZiiiJYR8AsPqmFtR
MINioYXMyF+N2xfxmQplWm39Y0HgPjgTCYt0ajXlvbBS1bxiIoNNL52ZK3yKO/QL
5Qs90q8MIQ9Od6xkGnpJwQ==
`protect END_PROTECTED
