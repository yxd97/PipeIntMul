`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Fjhfa/I+LZ7uA7yNoYjQK/dtlQFWhRefJvkyFbYAoDB7wHk6lqnKBE6Ya2dSFbKx
OzTod2GjhKlvBk7juIORso+GNCTGtgg048CVRCO7Z+yvOvTyzypukqXggCem31xK
h2hvmAYuHacxza92S1rkfMpSVvhYHn2PuOfk8uh2dDQ5QikpbGxcupYSPz6pkgGJ
kXjhaYDsUfiPNICc1gBVufsjZmZP8pHydOTjzOEllcxiYkZmaCjEfvDMbp7bP5Ma
PiQQDmPjyGxm8mJnyXFZpHNDVV+S1CfC8sLzgTmHuDBg1IDe4VqEWmd5SYd/J+Z1
t0orneK44UILuJ5U6GEc4ViuT/fj7NBDXfxMdJE9RzmO/0eI/74r3HYqyzdiRtrx
8XdwcqOGlrM4xo+4LxrKWg==
`protect END_PROTECTED
