`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rzUSBChD28eDPeYDLYVqhiEe2mk0G9Mvrd6zdPybBTyzUQBcYXVgRkJFGItINM+7
YS1NWePcHpTr8WUBU9l4IJXJt/Zsr2/SPoa1bXv4LqqFGmvaKR9xJMaz9t9D75E1
b+iA3nCk4kGmexLJvEma9YbkLohdlk1OHhwiCZrUZB/P0dBxHF3+i64fc8Nm2evN
fX3fgFObjgmI3qcmNLkp03m31I4phi8bgsb6WxHs5PbLejhsPWEmMUFBMUp7MrUx
tq8v5Wt7sIAtyUA2XJHKQodNsF4a0f9qHIHSC5xAgjCY4ILWiPPIFHzxuU1YSylp
WyZqcTfMcvMso/cnca9QjT1mMn3rBa4ivc8KaVIuL45AKjDLEVAeKdXICN6swKLs
zpT95qLhKZfj1oOsPabRajQKT5tmpS+qGLK3ytTPutwNWescs5xdk6Wo8xjZpsfd
kpICAHh2fxr6UfhJD2ocz+Ki48ziN4037AtGEAlY3RH1vKOQs+Wzi12NUFt0V3Gr
R1PI0y8EVVyEK7YHMib3YJmsTqVMIChZ13aFXzluJ/5OHVBvXNuBWdkf0+d/YA1Y
Nas4ukreIESv+cm6X0W6HIsaaZuVnErZARkCfA+bH2j7883J9eoXJSellwPrSIRt
ZK2IATW+EBWowFTfxsg4o7l4e0MU+qEqrLjdOFaOLOL2wDkIk3TET5yJhD8zfTMf
Pp0L+kv4b/iehh/h2QUSLqWywhfiN4D5mv59/0jgn0qzoKWOA91HiF3oGzQa+EqJ
vRTC5LJhsS8UNwcLiq6K7bgsIqlZtVxwbJqjgQ13i9S6od7f6M2auHi4Zm9l2DVM
RalMsclO0Pv7ZO1VxTe9kv8hHEhTarGVdHDAXawbEkk+kPxA3kGAvMhCiKv/pK04
0DF9DwYszCl2qP5r+7PTCaStFH6XmznZdz+sPrRw6wpRJpDeSRWCHfelQGBZvLUJ
1jAOjfAun7Nu5TrkJuVbuWGSUSg/ubCClZyQ9bJ11Km9zxFGMNC/frCSQX35cI+9
pbj+SbOWWdUhhxKPfQ2/gZ992NLGOXUf7A2wr7+6Wrz/KXkMASalF5HgkDFBmo5b
vtplX17IJKfTK+oPULnQbHy7Jick6Y1vc8gRTYQ2zTyg3PQn5keT/G/Ut3sQyAh5
m89b0F/sjov8/k99BPFjkF1DhqQh3s1WPOGG9EnXD9mRQRyQS0+GJHt11SkS+bKR
fjMux1mN41aRTUtUnZ0RdFK77G4NXBg5BDB2Hlq16gcYN3Tb2tj3TAZPbDrHR3Pm
INdGGCVtx7x2PPwma5yRfdLM9fYY7ReirmclisNwyFdczyKxIFdzesRc652byi2W
RWPUWKG56p+ZFENCl8GDm1261CWdDBiaPuozqvptR3VEje9NrDx7VJDDockNx04i
Co5D9JNdxrpthH/NpYqoV8CgCjbL/bl5FPprYngUrDLpDDLWLz5tlQBZZWGvvCJI
gCOIpfRyuugckULZCUxZEx2v8kBtcf/tR5NRnHRAFxnNjqTWNzffZGopwf5n/wfJ
d42X0htL9grvkj70sZxtRJ7LGJ0+YbSIZJwAl3H1wt3bW76TRAcPhuRxx9HOULBG
vvIz7wjKq4In8AG1Wlp3d5oY7zaIYu2XVPGGd+aLM4+KTgXQpvUm1dRZe4xByz6O
ldh8hOUUiUG1pmFZ8WPNnGt3vzEHdnvVA0gxo8GbcIbKBrJWkycGq0sTVr54Vjl4
taUoM/zFSc1CZNnUruaCUDdfjiAQrEjRcUZbFDSKGQ2J+NoDLHVWGh0OPlZqd/RN
tSU7enl5yJ1fawoSGynHbjfB7CiMrEDjjBVsB9Ce0jYT2K0aTiqgr2DZLYVg44Uz
XeWQIyLSpNCByXv+7vpeAw0exkSU7lt403Zi0ziCj0O9rgj9uw7e3uPH32YPWM52
xJIGMIw+z2egnkOKe4LU8muOv4OzHblfTtIwBCNFwDhKD4YpoaY4qHo3g+EgjTaW
IvH9sefoS8pQyFyCcwwQWHOF4C7IdIACtNBSVyEwMLSQcKv7rc46ch4LLaHRKGYC
XD5Y+D4E8FGbBK8uSjBepuzkyigpdta1f2/koMUQ2jXY0H+t9hGV4CVs1LOGGBwE
o5xt9z8WB6uH1bEQRXNX89VKEhQOdUxvenX4Wr8YSdWyAsEeVt40N7VM+vp1fClZ
hlaUMHXxWGIPzYhVXwAMm/wzpHcALZYJk3QaOUmhS3AHcTTNK7Uxsc6+Ufxc+UNf
n9GkFf8/TUyDNPFzxFlnb6xBVuiQiwqucCbZ0MeAbuZCtsi87sb9QLpPRBD97hBj
FMk7Bkxpx6rrVyf4EHoAqZR1x7ZCTfD/sjBqxk2yiGAF+4gkh65HSuhEw151MpQ8
qBLTfp28LhZbXtHyQMl19ZPfhcQIidSLT7X3J32Lmic=
`protect END_PROTECTED
