`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6+8JqQUwz8gTq5vtgiGd15MVLampUWRntOmxGaeaIVVyOcCYdrX5rtrapqSVLKi
KDIq8EzZ42uQRLtPOGCietfWLbF13ysQPO6jzDL4gJE7BLiOD7EuaKDtMJcpofYl
uQDqhFFNSf3VJgmULLCo1CVaG5MZIA0hxq7j/V3kwezIZZjf1dIYMRWtdHTDyK/G
9eYCFaewVjFrmdm+FDwjeFkxqWpAkOCWIUxwe3Pq13NHfZqc3MkY4PnyKEuFI1UH
PmofCVgQzCePhBv0dR8LZvyIIboP79TVFbTcUz0Dss7DUrJ4U9JOZP9kOXz+Ua0S
E1cTkVMuT76rE1yLfCzX3ADqdPT95vuI41GaG6j2BAKRESc/Ltuws0I/9cqPhvZI
1Od7/Af+sNAxexFT6EInIVxCXwLCeUY54haQr1hsbpb70Fn2VByioZHn77jsXZ9r
S2hsTaJ0F9jr3JCPKHlcU/ZqW8TQgOyDr1e4LSlumNMS2Pdy8RrHuoWevKbGtvRg
tE0MlVy17CpWdSgSOae694weF5RAOOljr4CzdM8CmSXLnLH/UsXAJZNCqVDUsWvZ
AdYyN10geNKVS1dwq8l5m0RXaYKOFx0/3AJQvn9bO/ZxiN62Xk89kSGahzG1gZgr
zF6qrjAvP2j+VlBTHxSEY0UnJA1b7JWGSsfAhV3daX1ufWcl7KNBHCjLXE1kKzKV
cmI75Yvp/vcXcgNwFDc1VsjyjLCDpcXp6sg4AWSPig5QTHRJB9XwSKUXBwhzqNNQ
zBRzex5rxVmCkh9YKFVW8AZp/G1kL9bv5lQv34JiE+24wZhQ25NuqcqL6esHLuYq
NIxSU4R0TtYhQUmv3+khYGOY4H7Y1Z5i/Li6mNCACpOaxi4UR6v6MRQR3ERDZDXe
YioCA1X6EOBKY2TjipHb4C6v6CF0y2B/uIlFgvoYbJIMeu/rTwjj2ol0KH+6Lcj/
VUCgC292BePb1vOUKx9x06+tKpMrkUetviEjG36ZhK/6PXvrm40lFB0q2iJ7kA2Q
mm7Lnsa0fVzUFYTMfdy6LWAjLfEXbcXEu3Hxofq9FvNONWJ5rCENK31e6OWCEIp3
/USYTixsjPb0Ly0qgS+4GdNFf+IKoTImKYxfG31vrD5wJHUgRJtKDGGjTAHhzTlB
1j9dml0KYnJtlXJ0FkefG8tEH7HY5KwOOSO7GKkz/Qw/ots50widmyZqHRBPu1KW
D0lrWrgkIggF5LPlclI2+udJ8SjixwTjoZtDN2MAA1V7v5TneMZBtXFuxOiy+MF/
qzB90KxOqe/iOYOKlLDoKaHauYdP51kIGKTWi4HBsz6rowr8gZTp2vL+hYpLtsd4
I44zpwosklGYdhtJhWqatISnDAakgHs+WIlUIiN1xjx2J1Fo7n+aUuXywqz8jkfj
B4bTiV56oL8EVhhyFkMz6OwlPqC+xvTOCMoyQGLbxXvxA2YeSTbe4QwOCWoaXxVV
LgfanqTtqRoKFnwBqo6iZAb4AKpNwJ4qAgljilXuQ1Oif7iAniQfl64VBdwCk1zf
ltRU4KpP9xQQ7rQ154O66oajUNQtDP9MMY6gnyxxpsPZiM2cMrpH4S1T7PYt7j0t
aDNXZ2DIrOIGdOExXSONTRkNFWIXM61FeygyAv0kIS9SWe7wZ1Hj6MWM+DCuItLA
ARjmCY3lEUS+pg6ZP5NeA6cOO9A0xe12yZ+MFXTIEBitMlkOpjZ47nAHPQTWuL0M
MEvz5aKP1UvZE+B2uYq62X1SR02VhtJcXVsyM5EEBeLbLKtCCLUanRm/b/mYij/Q
r9ml572mj1rFNWyggP/4m4pzMqZkKnYLGbB+KG4lT/V6YZFMwUX7JbZZ9ejHkKb6
CuMmRt+JHQ1eeUV029RSWWqRvHkR+jpM48Tm9h7b6KT3W4n8MbPl/pnTzqyFBb5m
7Q1OI7D+MDDdsKZemyGkD2R8W+5xxL4xveO3WoHmbWVY9wnDQPE293F60XZXZxmn
Qu7J/L4O+5OSxbYC+jT6zdlBaX2nAAlRyLEhWwgZgKx3iX0N0Jm6kOy11LN/TKlC
4O13cXIQB0fJHV33i6nRV+e/m/FJGezgHRZsrmpcADD/12wG0yPHsfuIuiyT42yo
FqlrrAp5L/O12AVzxNrczi+JpFR1L2xstEoRYjSg7jLQ3kIN3FiazdcpWqyZNP7K
er7c5juouzo9i/QMirQX8g==
`protect END_PROTECTED
