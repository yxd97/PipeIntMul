`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6qW+CnoZ7GzIXmwPdHDFCKEDfHIaVnzIvLVdrEOzEgdRmbX+JVlOmBkXYrR77BW
6VxyTaKW/Un9r21y4CUH8LX0KqEOZyNMLS9P7/QMeccKSEbEWHy8iEHayJAhmFa3
kHoCpEBjqx+RpKRG15CeTaejWIRHK81ZYHjnbBhBq56gLPPxNwjdSaz6NF9LIy7E
aP34cqy0B0nIL5U8jmfBS5JZ0ba8MEv7eMk4F6L+HXAnPBgKczMDodaJJs7A0uoa
lulVKagTGgeKgRl3yb21Ptg/EMDjUG/ruTgl6BQBFyNDtAWGac21Ky2m+yxD6Rap
5daL3rYB1F8HupEPrT9Baxuv7L5qKQkKcJ0bOLeUhTMQR1YWy3Nz8jbV4hSec/F5
aG49SZSIaA58VREabWO/TeCHtgtOLoLWV1NSKNCdLJauR1Bj5Mj1y7UvqrgyfULB
egOICsMF8AF+MQz+4+txzuj/Ije7VMS9MZgBSVXeLCDoODi09HZJxBXngkecQJl9
XJz0yx7H55KbivwyS9Wj7Bt9aXJC7i30S3oBW4J3aCCuJTtjPCeAWqLnurvJGiDr
mHfzJMs6DEri6CMyntd7KMP/xduzmuqStZAzpJU3s0XpisJFAm01FML7dZL4mUrT
voLXQ3Gmkv7J7KrZmxDS/B/HcOr9Grk+HvtPYqmw4ujJ66XME/XC49xuMneCPg+F
AyGD0npVtouDnujaeRfpyk9bdrLCxrwyc+Q1Q5WtkpaGXPw/3J7JJYTlGhT9Ofmk
uMLYMvuNMS1qxd5p3yTyp4NGXNtM2uZkfYcpioULVgPGyB++OnzxY+65yLD+OpPA
dIFtXGj41GPxV2sxG97dd3K2YLWuxcMpFKlJQWkDm8UWFYUGVXasRBWHA3FXG/LB
FZc8L/yFc3X+GpcwN1ggSWsLcGJRD5osPkR+z3/OWvwNAdq4QtA9olQ35BnCb238
B/Zuo1fqQR1SS0BzEDa4PFIEUYDIvgx+ml4Mb79WJLfHcU/N1Qs+cruqUeB1TsNm
W9UltzOIGrQNOipoaay6pSV4bEgXOjgr7VX5VOEyr4jyA7i/wotjunKTDhUhIBPn
Y6NXNYiadPJ0Dz9sJrmBsciZWA0yoptIeCu1Iu8fqrGCoBVR60cvRj1tf/UTAtxN
Mla1xlDayy1Jl1QKN/YT1RZr2KX5pS5WCYzMH2ly4Rl6QznwC0zKYknUtxHqxvHf
HvpaZzBzPN1u15ZkzLI4V3MBkQaeqpeauzALyg7HgKa0CHWM6Rgj0g9WWAbRrWOC
bfoR1ivB3YrkzV4ws6bSmDMv0LBl/0FH96KJ4YoINRDMOZ4dR9O1p6LwDLb+Jl7T
q3hLLxIuJ6o1odbxwYJA1xqc61iM2d8xdEoom0CzWldUjk8jnfLWq2lcahXyvido
ojkN1zO9uBq7gUs9qE0A/Qzunu4xuji02SDOtRYv/dt0iigkI570lwSapgr8SQa6
D9NBqiSk+NiOi7F7qpw7MkZZHku97fBl/+sVjn40icKvX5NRoF9DzRC5pIo16XcK
1ha0Ny+f00Ui3Mt3rRCztngccX+G5atnEJAw3sSYW2GV9bEE+BY5R9QiIztpcHnt
AFqippNLu1l21Zr+QTHb+XGYreZuDjBEQqseVn6+chGdWlb8RVMofmTiNbelvoci
6PEQxw5SDPqCEbvJmi6wN10+jZcn7/4TND4MbUho6O7A9DQ5ua7g6zvxDopqulnz
oAHyeZ/lYXWUyxpctt7CyeEyLXLKXgpJZiJMvl2o6lVUcocvWLlea/TzERpOSBjg
8BhlMxnJE1RTwo4aIP0vS+sXmUODSulbxWqMt+WJMfKxzsXrv/aFeId+Qbgq4XyU
fYPUWJY17eNplxJJfk26YHGxztkhCyxvzC5kZaqiID3cwOQqz63nWD6BtbrNuHBC
izjBbcQJySVsLk0A56+Uifu7L8q+VBr9zikCo0GG2QKy9Fv88NcpG5Gnzls2SmrT
H2Wh6BTC+t84wfF90WoWTC26bSvCWH8mDPpo14Jy0ct0j36GFF1AOr+zk2lT/Uf3
yGRMo89IZ8CvPoolLUZUsy+v7ncZEVSkzyjADaYP88BvTEFogJC0N0qi2M5mLQC/
SKLJdap+JXeVb0ozCkHrPsAjhzN57wvcAbWUsVt2jRWoyQwdr3Y0UbClhWDMH0cs
quXhqxDaSeQxvBageg0HIyPgM9XVSLTpV3XQpuWOVWxRY5Ox2nasB3XzGZVYgFog
zxChujnh0jFnKnT8VRPXaZIMmzRy3WH49qLkA/GjuguHdmc5Fik6przBLzjWZEbG
oQ5TZOlxEX5FMUSM1mvMsLed9SREPgI/hw0bDoan7M9UN2VtSKEta8QmadXvP0F2
kNgJSAxxELZI/CkitJfIhSp9F+adsJg2HKFbBkb6rIN/vKuWzGQYstrWHSRe3NUK
38pfEsW/QTdnW4b/zyx0pu6K+WxNbWj4aTYZqU6KNiqSBQ/GK2+6yxx4nWAiEoPe
G9UJRNAKMXg2x2MzRm5dUwM2CPgDwyUkvSSWl1Zj23buZGAAkV2BEbCZC3jecryq
1v9bnT7ropT3KMvBYJYMGVDIIg0809rNqEsQQBEzZJ3qF9XW5tCB744ZlDUSJ8Sm
0evNHy3NmAuN4rILwcQgne678voYWddcT87qOqCb3P2dSa3ZaIVdUOz1FSh8vTrE
/bgScrIhoPnjYwN7nB5rFA==
`protect END_PROTECTED
