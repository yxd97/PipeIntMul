`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1g6z3S+vuTg0XsLuRzHnhM2ocxrjzLNgJvh/DF66JYADE64LOxu2XLFOQXvZhF3c
CIRimyQneIo636wMB+grK8A39Qd4Sui/kr6vch57MvTLngZQ+t0QHFeC7DJ7ecKE
xyQpa2OHghTbnYlEN9etgIOqSItiFE5m/cS0UDN7bpDeqttHMgsDj2N3KHAQ3Z9F
5/U+JoKzQRgQ2yLYfEZ8XCT4uoAdyBqGNjvwDwGYl5nf0rpLB7gs50Owda2T//Jw
5IwivfLPxNE/jiwrtJWcZZSZtwp+rUe6DRQy5vSwaggQWl1jt50eZ74MIDDJoHT2
KsrJZRYGGCtLiPYr+K5YE0PNxgVosM2+ovzr1lPryxn7rrL0zXEUZyHGiXn9Yda+
ig7ybP/hyRHKvolge+qVmEQ9iMz0rEUiJScI5Fpx4W8tjxpP5rTO5/aoSBUdsuOH
FC8siaXPktqFEnzeq5Z6BS1wIien4+OXfU4KHRWUQNye0R8Xnr+I5YwxVWWEBotI
Bif4cB1jt7g/btYvg30rONEN7buWD5HRx5aXbwTMpUAMIln//WcA3+4DjizF9TLI
CH7+6QMU8s+YViC5dy/YngqTf31K58i3EhXiSf4ZEvcuNyyHBjluXkFeEDA16++E
6QWIBTtcWFI+dPZtq/1aKdLkS3nqDS8X0O7csXIy2Do0MVDkXBlEQFsqH0RxnmKe
3rS+L1dFb4F7DMy03o/zRrF+2C34HlRMgt0WVqffEeTKkWlgcCb4Urcml7cl7P0b
ajaYUyRNq5FLCkn+ZMw2RQ==
`protect END_PROTECTED
