`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DcF+GJ3vCUn4XFbeDaVt0lLoSwS4GE26ORGFq1iiT9DvHiEHMTTxV6wSblI/KRbD
G7/C7vYZiIJAOAxvJDOMA8IM06O2neLadppRi9wOSMgSZLUcpT5qkCmp2S36Z2Np
7WVEhMRQsWtJ4PX9w7YKM/cKsPudj4qqBi3BzHQB06LYtAO3KkVAmL6JFw4dFuuz
lxaBjThq8ycShoanM1U3WG8Q7gbLXuHGTzfMOthjQCAcsD9GShN8XCFCdXAUTM3X
5F17QlKa1PhuewdHJ6dpETxu6lNE9IHxQHybkAzCKGvGtNEGMMpI9SSGklHMcDJN
/R7fWAT/vNJMGSEQzCEDlpX82A2g4iX7ywSEl9GkxWkd/N6z4v0Jlc4sm/7f1Wu6
iBLLl0cn4NjIruGUQCj20HaIPQYjCMCdf5EIsoB6f3fZwXaDRNfmlEH/6e91pgYs
vMGuflhpcpQt40bqoKhtCBq+8MToakQtc2omwxu66nQcLnlCAlyDC8q41V/Qz7Pe
`protect END_PROTECTED
