`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZrLvlgqk1/G+WE+iaZKGRy6WWqQ5hbco3ap8L0xwiLVC3AmI0MUBCl1t+KnzBwBj
0G+6lKCSaTukVPIfORj7I4oX9ovMwOL8EEVGEGgkp0TKoM03YUP5PGqeT+vHHFne
cW4SRyJ4CK+YvzDOO1kpADz8ZRiuZOQq/JsG4VDvArlq+myIh84CwFJAg+7oGHV8
vGXcBiyCKW17/irrgpYDgUAPumpnB8crUbuKpop9FfULllC/B1escUHwFY047Ewv
6Ege14O3smLSowTGIr63HA==
`protect END_PROTECTED
