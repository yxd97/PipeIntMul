`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b1MvJL62CR99S3Tsnjbs7x1NdLKFmCOOUhPhH6dOIyjbqZCxdfN5s4G3silpSmUv
ic3OI6OHTpd+zx5iUhyH05otQ4pKnW7ZOKBZOmcFaLwWhzpYWfnabBfI/TwpMPkt
JzliZ+n+09UyWHbGbUeC2wKNJd0WTpr5Iz9QLo5pZBIHXagzJ1IVEsKS7St1d0RO
6VDQqq6aRdHYjuq9RoxWG5rvrNwEg8L0Rr6hYTHSngQIPM4jWRU5Gs7yH4NITYHY
rZckqa2Xk4YrRqEQKO54ujHjuegJrjXdTGy1ibg/VYxgv2GKbtYcUMF7To465gkX
YP7V6LkkteJULM5iS81BXyjagQ+gDeaaIudLBM1Ie1IdgX13PBZ+ejJYw8U9OWpt
mjJ32zu38GdtA0DtOnKkKSbVWj/ADhIBIbZIEhCsNc1npn8t7zO9uCFB9+ObvlU4
DItwq4xJe63MlLVyhHvA4CezlT8DNEGZ5tgucOv9JNIKeY/yhDDCoBMQUEUd7VeL
+WD+bAK7g4NJ7JtTBWZcqgkglMMMxgyHtNZBYtQys6MMyWQpdfvcsFwC5OIay6nc
Vnbqyx1AIe7IvAiGzi7dT4mSh4WVf+eKX04PJ93pVwxhegPcjvjd1KgZAKmWBkfG
YYcVNW5urpTq2yHEm3Tu4GmAPv/DFpglpCbQNfPtqT6RbYtE8vpfH7K0JJ+TADtS
X8Nh0lVX+RDNxyvkmT3SOUQ2JfEMGbTnYCWRa9MqDIIhKM2J3yWTSoV+FE0szy9Y
o8wZNnEEIwdHBy+tCfjWgYC00z/P9fv6DqIVoBUkqIs4N3dHvs1DY5r32VDyzte4
4MmVSwheZDeps6CVoZ1BqVpqieb4/UenKXDuRtLz9T2AulSKKlxLTLYl9JQyuR5v
TxDpZR4ZYPlAl0GKFPUY7b49FokC7stQvZLjBV+Yb7QH0m4wqEh2jpNX6bQXuGXU
8sHUtHb+MdvEttQ+IgNWnwyH4GSV2QCmYu+0A1JpE+py3Kta7et3EiYnCK4iytVf
2jGOECVoE6iwIV9K3LI77tlT7aiTBdUJe5RJP/DcLwuYYHjfjj8zzJkZ4/qVbPDK
yPi50iUGkxNLiEKkb8GRcL8Wjqe7KxJU1aJ26Jsl+TTeJIuFGG9WdzeuQgS3/yy1
/WtdArpYvgtBio2nlRpzGrFkKJObZ7MJQsta2wDjnf97SI0jhOyB0EX+yG6TwbzV
UlP4dGHfLnswy+QkJhf8Jg==
`protect END_PROTECTED
