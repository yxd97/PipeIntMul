`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eRU7tgPkDO+pkThQbiLmod8vy1Af+1JZN/lP2OEfFhwQxMC27v0a1nnjYaAqtEVf
iGsd7Jc3BM6hLRQnOjbt5aU3g1iDFMX5say57Zipo80IP4+pHWRtPSsKy/lQDxgM
MAX7JWrfLmdCj1zqOTGUyu/u+IZXYpS9+ENKfO/hVIFQ5vNtnBg1Ir1nVohxqo8S
bf0m4xwqhrJbeXPhaihmlez85oIILAaxJQM7ebMRGfc1BkoJqk1PjxlSEOidGL/T
CSYAxJf3640qRtiKz+DX0y3+UVGT6a/odWyuG2eolBwVx5S+61ZGT9m+smDhkJ/6
sbfwEOvRND0Hw/u4F6fj24SGOAeS42+r0Bjj15KiVK+UNTn/Gclc9iPvijC0Xa84
xDq++fuWbT4qveLQGTt2txA0h/EjKbyc93JyN4LuPOAKbTU4mJZbsvQwFqSOs4VA
0hcW8E6mvP2IWsIBjk2kGXrt0N3bcA2Yctsrjciv6F1ZCcGpwO6KYpkJBtQ5lo/q
`protect END_PROTECTED
