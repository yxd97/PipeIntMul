`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q5VZL1+nBg4Yo3SE3CFBcbYMQ5yqyMMWymSCN2rS5qBh+R27o7Klb7OvFWMLnQGI
lcyhEqDLgGVkPsb3ZW9KaWZIXUhS70nLuZF20kmAXUOX/l4VNu3OpJx+GXHkLfsG
QzXXLh1rs5V3MlzwiEUZJjkfRWskNrezOGSzpFyWFSLdmTMEKLV1fkJmFSRlutwb
DPI1jThRjGA5eNSY3PxT0NDLEA3reYNRDrcf3jHnBx/fpAo5rh+YRccGa/fEE7U4
vjtzOOpNfrpDUlmKLs6yjKwlIzziV+pz5T76gBPqfaolSdq2VVGIx29OmpcfJLsb
MYPClxQ530v8Z+yEmh3KPQQC0BYcKF87vfMh3AAOl6zWx7i5Q+pEZLoN04jQ67LZ
g8vBU7m5mmfeDNwJHSzPPA==
`protect END_PROTECTED
