`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibyoIAgz3eurKNy0LIed4DSU2uZjd9f2RdumZGvm1Fag/y0aogNwnPeDdcOREgev
ogJbFTU2NHNxRMynuL8ehDntX2YnO4NYsOC147qQl8sEd9JGTB5ZDLYrUobgHfZA
kVOwa834Heq87XjCn38Ehi+gORG4DC5L9v5uDeO4qNdrzPHTGdNT0iZV/gSwUZa3
IjNXfhgKMiV68po5N1rOfoXmGusVSLAX4j/0dYXOnf+3r3ndMLiU3Sl0/mekZj+S
fijCh2uGXLmTiEsU/Escd/RFnJGviqUCnCdk5m5huQv6HcpfIpPUAIXU6HP7rGjh
1q8jPaxKesBJ0VRxPV9KD94+PXlS6e3uUibdbFDN8uNRMcyAQUCUNt5X7+0qDWz5
HWyztkrr9pGZNAgYW+LeUT3AlcoEHKCR6myKO4JSqVQ=
`protect END_PROTECTED
