`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFYCLvKQb/rYHYZjZ5YWsu0k24x0w5SCNWrcN+u5fVTGWMDQDvjHDgznrioMNzRH
wkDYe/q+7pnfX2KQcOpYOln57+Tp/Q23z6c2tmK6+GJM97Xt4SScIOqIzI2pgcfE
uOZC0Nx94XXgNjFpizJl2DxSvVelPMll9+OHSswwLsmn319IpXCAw5wwzw4XWTwh
ZbZlBZk+ss7QNy+bkNEV3IxG7gWwPW8K+YKfWGSXNtZEB8ONfh5YgEPkLhBl0Hle
vH4bFLXk/2JUv3TMfzhnByOay4YbvlQ4sPDgUjKaQqYe0D8sNjbEXO01MEw2mtfX
rNosJqd1Q+G+fs1rAhx395tvZIln9VhZeZMdzgk79aaOVhegcP2drvzIY87DXVY/
RavLb7CXTVpEUJcRjgXLxKfHZ4nVL4kpgeaiseEXPxk=
`protect END_PROTECTED
