`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h8VFUDFINHecw8gtkcFQGIAbRqxIz6rjYy2qIQOIEy/FcO9F4rfv0ssy0hmatouo
wrdYXjScNhVTLmPcuRXMouWoXWTejJbFPAZ7WjJUW4CGmSUgzge7wYCepb/1AFbP
+uthbjXuF11QmA+or9R0dGWys6MskIOY+ss7tTEJFvbp7BJrLvFQjKV641rvGgDJ
/5mOpHmhSfuEqmW+STUKyFvRHvB5A9E2IE3uruUSyet+UMTguVuGCaKCbx9v/ceW
lZW96XIai++sT9BWaiTzR3pzjh5McWPqXkOaF9g4WvI7NmYujf+tPuBakYhUsMdu
HyTtyrnVM16L5mzu3t27aIHkkLHKLy2cNRdmJlAc99CFEYvh5IbdwtTYjiI9PYrm
kV5TrvwpD1Dw0Xks0nnQjk8jU0YR8RcCaSZyrTgJqo0aYOYugA/5IjJ8NeqieRBp
fDu13tIe7VBNMdoIPeg+L18PepYlse0ZGdqLnTcPbSx1TGrVK1+31Qx0RlCWtePc
nbbWoNKbJUYku3QYS+pY2M8aJpBL4FOnFy2xiaXjGFtO6IQMB4JMFkgUGCnc9l13
MPjucXMw0bAutiW6dFOyPA==
`protect END_PROTECTED
