`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5sSCtN0+tZfHG2QiJ4WMv+Xq+CgES+s3MoS30WTyiGUBDRh+w7E7r3QpQgwhMmys
yNg29ri2AKj3jZduDkQ1POSDGIjETGohHR/1ml46C19qMFZGeuIEJzxQseL3uwRy
mZbMyNWbt15U+gpI9VYdC6BgLmdMMNZM/cD+ikatwmFf2AwRmaPkYwZEkWUqz95J
+x7Sqd/k9KpyCszI/JrqhmaIBVzJgwmfNoEH6d8kncfdAsbrPiXEznzHWrKv9mW1
MEo9sbycFHvJ3SrwH5KFMibHgSHGesJZASPycXAgIqmb1h7TyywmzoNJyXadg1ph
u9n7ukBLh3nookYIWUVj4mem+ARkH3jJyZpw1DRGHQbgTTR5vkzq9FxSTTSi/VEY
Bx9h3w34Tro14Sny/e9ZTC3BySfQuorIF2XfXROL9KyFAb7qHCbnd+JdyBl3NUi1
cIR7c82VFvlAD06xX0AXNBY6h0P2vildMfuEVmyhPlFpFTu6mSpn/LkB0J0PquS2
S3Zc4lH2Pi03MbU2sumWc/QalVuN7yIuSRlA5gnW/0dY9/wIgVNpnFyBko2r6gLZ
q+q07U3RfYDC1ET/sYmeouMm6RW2n/BHVZwRHiAevr8tQ7uI7gxAvNm4upFTJL+5
fknQxzZDqKrBTYirih9AxCZFCY5FVvBFCULnaeQZv2lv89yvh1goJpe7X4itTsCd
MPldx4pl6VX8/2UjcEUyhgTDBgKNhrq9vnL82NNfFIcuAdnYuVBl79xrxP5Grnn6
apCo54C/4l4cZ8GopI/oYPrQNl7JsfvX/EUio/83t6TViE87rXpMHeNtBTKgKr6u
F2GebIa4IcIOH671YMUfbHF1BEKW7e7Qv9sXjfugll1+jq9Snd/s5pHxwsTAvI+q
BBw53bfzQqyDZEQVVIqfUxxrmaRUgZZ25BZP2oRz7+T5ZyOVERYGvTPH3dA70cRH
S31fUQZMsqbyu8H19g435/OPKm6ht/t9ZT7/9sm/4l/Mtq7S1LdqLSzYPCayoMwY
mQiz9xDBaEFkFIDJ2/l5uNH46bG5m4VzP657oAqoZ9VmPNVgTfrzDdQz2zW3RxMa
IXyhFRNvfPgHG5vVCDIjS3CWcvlUnClJfUt/eflFNV4aLRZXguc6mIQx9zhlkVlm
aWZxOWqodumLMxgU6MdkiWfGFSIx8DrBWyDVjbxDiyJosRpBTlkuUum9axr+RWsq
ubkNh831MBPWJQaH1ZBEcLRmy8kuYF75RrO84iZ5gwTUHTd4vvewpyZJ8SCwrv8H
7bF0iYja/144XVThvuYqb6OFJbrsNBgwG76/uTndlUOHNIhhzf00t3YuRdzP/edi
gNZs0lhlFvUssZU6tUIpE7L1L85jqrsimWDuLWuCNwWCTvzfOBD4QZWooEOmfZs8
wnMTtImCnYELe2fXYts9OsNIT7v46ByJOhp0LJ9EgjaxH3WK1MYnfo8OSXzj5Q6X
hRFM/WE4bFOgYIuXpyz6VDfAicKm4DKVNmX+VzLldG0wALR9mE0X2bpCiyvGUW4p
W40x+jhug9JyAv0oqOOcdWy+bHzGSi/9NLAC8e2g185h9wBHJUb5iaX0rLo0b09h
GKeT4sI/obqQdihIlgIqK56nErHuaLlVS7Mlr8pS+2idCTMCM3b1uLK4w2u+ToJf
/qf8Qh3fRM7BYX7Z7pct6CfJoLzteKiATpTSv2DQvtHgeLd7SgiK2029JRF0V5g0
Qhb6W1NCNJD576V2RTfXWo3iR6D8mrw4ky96MypqnKc7krktcJo4xtAUI7ebE4r9
/bYW+5GGGJ/rtaRSYIx5MR8hP6sJIzgRtHoRv+l/xYJ3er0QvFZB+NjOha+5dlW7
lJqYdu/3+3U2oMssZyLF+bU1wOcNz+5yNSbF7JGWFRA7uQFYbcQEtnJI0QZ/xf5t
f1mr3ZHpTHlp2AhKDbNMDqwWX6HqozOGDbz+KZXUTzPcYaI0XXBGIlZ2NMuJarV8
gPYzODcznRluOV74cIcnpTJIiG19gpmbfMqGI0SPWeUsCaukz+Do1AC5G3NKW95Q
`protect END_PROTECTED
