`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1an2JE3sPmFjHXcmOsv8I909S5yo8AUDMzb7t+X2IUll0rSqM1dT+Oy2ef7ktdmw
ek4yCgPsKSAZB2l69JKtIwQzo/3QkKqGcbOxHcwFL6QrMfGSsuEFve3Gks4iYsDC
Ae7QrPGlthG8yzB76SFXcF90T1MHw7m59J9AxATsHmYqtzqeyb41SFesW6irq3cV
PB+pkweZjJBeGfpU+93+BPkRG0SXo4992Hpjf86/0lHE5oTdpxSPXgv8tAufB2k8
tVkUub/tNxA9dqrKyS1RoVxz3PlZDSWsdwmrdO9iCBd3U7TUP8OtzPnKRVlVkyD2
MUx8K9gmjTew9K5EQ8ikh7lbxG5elg0A7iqDUN9pShb6QSm+tyg5HrlMn3H6N8ka
0OppN0uHyaYha8GhObVLWMT5hQwRKffOGZo+oqIUwtvwZlld8LqcMJtC9dL0Ez5M
2rOkr7Xa3k5z4pBit0GTbIAYxqawLpg7C8F7rWQaCD6uUIfmYxGyGOyECemWpz61
N68xSAROzz2d4TfqfY9SyMTLoP6HqTIryfrCh+BmWoCfKRmasPyQJ9e4QU5GsetG
7k30NVmYShQdAqJxPfMIK12oUD71ehR08xhV8p3JHhmqJWbFpUnf6HxvUU64Jg1P
O9+iOmTIeeoXW6Cfc2h6kAScK6AcQFDTUh+0rcPOQTDdVw4+OJ9ivkjZFs/Cb6Bg
btn55fkfSiC0PlclWX0FG+00C/FR1Z38LI71QquSEZoBt4ONBIcP6nJkGy65EEPF
YqtKC+M+MOvFDte2Fz3oYrv5XQXA5gRlNJintJuNdLFEaKfD6aKwoHHu2Obk14st
+Rh4AWDniTFaTZDKCOdc5OuxcnUjtsryTXW6BjteAFYrt2PA8Y3NE8pQeq1bfUQZ
`protect END_PROTECTED
