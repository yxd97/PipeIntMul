`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ek/kXZHwUSvAurQUjs3unoDlcdUiVeZpRPi7m174jaV9OnwuDLFga3dc82vY3sRC
/ceu5En49w9PrLFLAGZA353TvOr7yt7es0FeJDrySuWIJtJ+SK3UBxV/jquOLYs/
N4yC3fxHKHQ207ZLqrajFMBz7jjd1NKLnatx/WLo9I3f4o7W4b7Ch0HJbi9DoBuV
GifGDDiRGnDDrpQQYxdCJYpMCwmdEmqIDC33kSO6H8cARnfEb77J02Tpv9qVtsGt
qZ9HyAR4DYfzOHJ/RaJck/olEOOK3WDuiQv/4JnR3Iplk3IDFcAqobtAdFA5x7G5
riwrO8ZnfgOx9PbngNgyoJS0HNfQVh42EKw6r8iLBHA=
`protect END_PROTECTED
