`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Vt1kz4vmiQFOtf6zqw6yaT9Zoc2m7DEDRSayqb7M6dC2pH6eesiDOEgoxXiXqjXY
c3wO+wAdbJQj9M81igccmerLD7NVW9wiIUMyJmxPy93Q90ZWBdGokQzFc/cO11Co
bodG1N5ou/4ySxLLdAa5hjQYQ3yVFNibKzHu1X7Pb2lciFqSPw1wE4F2xnYy7jy4
U55rxPflStBPWdsqoPxbaQ==
`protect END_PROTECTED
