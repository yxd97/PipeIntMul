`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kiGcOlYJ3TE8lQvLRgN5SLzPpwYisCH82p5FCMeWhZ+BZ5hx0rBjaTGZvM+xG+i1
zACr9LB7HY6Z1VTvcZM1S/DUmWrG06yiH208KYOHc3OlM20OnUwMVX98uoKGnELl
6ABnvN8R1CRYkOHtGoZLD74S3wK+Pc9zIIzaSd0l1qIsJorlyXw0XBc0tNckYqoo
z+8GD4Tb63bfNNBloNZS1ZDnzBjZL3WsVJj5F7YosyZn0rljEkGOjhGUcmaHZGZ4
xdX44yxCH896X4crqb7hirrQxIZcX5SDyU2j7kfkU5TPwo7t06BxKDC9ZGRgn8E6
ZoV2ZEQzLJkGfkIG9FZXgCWhp6N5rf8D3Q7fyl0fy7/bKk2CqmHkZgPkb7CWIs+V
7mXSfwZqgsyq5eumnGyNKI4KUIYg1OFNpz9u3126eCUlAANpyc6pIAWnsFyUCK05
/Zv2AkmSntc8o19YENmJrcZeslyzy6PJLUv8FrI7ocrDT7Oev0RWT04GP/OkTG+y
5tnpSq7yNvBt3/mPX1AW9eCf9tYHhtcJtR44yvW2OTKzQp9ksE1U6OWHnnvR+5bX
re9HmXEOQCEWWHdIo/QFlfgaY/lW//96084WTNvqTIwNgbVA+aGFf6mOkItrrLNS
CbysEMPGvA/bJHDscS1hdg==
`protect END_PROTECTED
