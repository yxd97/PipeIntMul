`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c5YvwmsJ4OFyrf88yvaJl+qoMjChw8faD2AqKOgihhmol9H1MVcI6h81sfZl1QR2
TxYISesmgjMhR2uAIoYieu1iWw0ZQ6pAUgSUr59q/WIIcYpeNBPdDkoQk7y5AyHb
pQ7WOWPtwoKMJR6fdgBD/JTb6DaW1u2qdOBueF3a3ns8xJtG17SHJZnmZ+wA7QdI
CC0luXWZns3o1zZT0R1tjNJ8pS7x7LnsPBBYZg3Vwbs4pVgMA3UbJrF8KlbsU/Ob
6ncW1rG2+lXyxHQTDc7t2sfxTbHMEs4k4i7uGoKApHxMQRbkwGQkz1a6dE9Lvhl/
BHlZ2lKaEwBi4uoDYaOHNfeszVlxwImokAOPJSIlV7K4lkniyYi98Mmhd2fF1TX8
9Yoa2JOsAQXWtuQlJgZaNDLh7B96GvxoLt/YZhSMkVUgrPtlkgTpKtYd/woA5O9l
EZ31tLk1v/i8XdHqkMf9wU6UUmbIglyD1g2Cu4Yc48/Iz61OCItCRJ0aPr84q/+l
uzaUkNR3sG01DfcJ3KzNWsMfG3mkUiC15Dg9KS4FvBphepGu3Yjxgmb+AJz+iDpu
ebYpCwqDOcn9mpnHnUZ0fwv1MM/uuDaJ1G6YFmu1NcHerzACWzUzi7CaJbTyTtiM
kMxhohMtT/VhsH/1SUq4clzrNWKPnpsuVDCggQXWtMEDRhtwYo5XDKIG2bo33/zc
o5M1LCtFLp9tGmkaWA0leyLkaYcITEyUIfFBGPZy7StvCC9gOD79DjSh3G1TbJa6
gEFK7DKABXf6mt8t3e1+9xIAabDCgX7VAErKqjJW8TAY2bPqt3PbjVaZBQRezc8a
o5eVHj8ydbfPOdy9YZdYyHbsZGcbs7yHPWE0+1ihviaViHrMCeCqdPM1+j6oSscx
kbWwa/jDDhBPqW662tNi5hUKEUvk7SULIpAXVU3d3jzJLeiSlMlZTLCiH2OAItHF
m+++05aeU4QYSIuZCf+wmyvlbVnfnKZQRlo3nL5tIuM0vd6sZ6ff04ENf37OszEN
zpCLexB1Vv6/QtlefFUNChVh8f25poyRqUxc6OkuQ/8z0+uxz5sEZRsnTI8EGZ0v
859dNQTWYnvYBINd4Cue96cKgb5ZmyBPLR5cQswr253RbW7cBDaMS7F9pss+6DaM
cciYPBC8xr2u0Aj9/580hABkWLly9s8Y0BU/bPEAA9FxCSPheO2BRo6/lTm4Uyd7
8oWpQZONoqYJK+i0MRPhafsd2I35zzseBInl/xQEudIHax5Q9BhvPjbIcSk87hos
Mw0UVRgqgmAf31GAMCrmIOTpdYmHbj4EvVJX8OzTPHp1N0LzPmUcP3Vn1PwrJy37
Xs0M938mToHpYQon5L8HoMLy0bNqfOg0BqjxXeykob79E+326/qRzq8FzytJMDHX
NhrG3pdAosHNy1AL0762ppR1bXdj4VmB0UbJQ/Gha3LltsMqFqHTHEy4kjj+J2Zr
lyYEZ1180uLi5nPPaZsOuMEuv20db8u0UZMnVK175akCBSoTjc4/WM9/TIpeW035
pE/5tt2ILIGSeAOuxjVpsyImmwR5UqScmxFI5yClo2qxM95KumezOEsy6WNU1fu1
NJl1i4euCml+ZRHd0gfkpcCUrl53FLvopn3thRjR/L/POXyka7+jN5a9ABH3g9Vd
NhFT5a+UbABXBQfv2qVTaPmd1ioI1w9YAZOrSWskmRJY48KKcyoAV/oqxcTPzzaR
GdYa8daq/jVKQQK5cYQhcDcTX1rkGowmwy30xouhz9vOF0WEfFIqic8faXwJPd/M
Ozm1YfVZ4usbi+zkXIkgYytUpW4IKPPhST3/kjpPvcRvsRE4hWCbluds2Nq3KJc8
7ame357eee8Wk6WSZVVgWfeEJFjMBBerJ2vrutiihVUt7jsHrqnELPwgGtOaFqXa
q+OsyCKJtB0yjXrXh5T66bdghNBPdMPruYv829eJYjUognfFjYlYzIEKMNwTTvWe
TxHCw0fv07tvanlXQCzVj2bczcYSIVMkvP+cXpGASDYEPbOymqxHT9S9EY90bfrD
6MzlJac4IEw4VQQtIuZZq1v4WiJ5FyIsLvYd2pxcVnssWBf4/a/A9grcYdRF8wnu
00nB8iOOp8PAwo3LDnUh1D5FwP53e3eVqDbjmlkTQwXRwQDqiotrvoJ+4FuEqoyE
udaWIDAe+dxV2uNTNVjss9Wj0PUhlMR7jhqDNQYz3q9lZ/QmMpgFRAjKBKQnvL64
rqfDs6KduJi5O0/ehFzKo8bCWHRbBAj4/58QSJCxHBc8Cg6mM6FGNMeki1Jk8d74
UwKgvqpaq4UsnRULRmBWJVynPTdCnBMUdWaCJS9sydvwjfj5m+/V6NsbOSCLIni/
VivGpJHoTJThiZl6cBMjzsE7S7Oz4OziBgOpo3rYMzfi9nfxkSPSsHYhusZ+fKJ8
z6rfgSxx3DegxANgPWEPk3nV6QF1x6dw/3YQc/pnpyxz2Wj83YJD2IgGTkJA7uu4
I7wbDRRF5qQxszeNmx/P43jIS8+Dcd1Mv+plVMCFAd8V2sm4C2hltNe4r+9dwe80
qJbYSSvIWb58Qd73bFaqg43izwN67qoNTwKdRLoqreeL+yvQhNmNMP3mEpYHT1PE
zb+vTKHXc3xpfAwKmIkPWQBcNCvviwMABSx03kEmMjk4yxaRtMOf6WwuqxNElOf6
JR353WDoKEH0XyKbR4XhV1b+haZDAC8XY6DlXyXI51k/VkNtyGufby1RBJJ8EPh0
/fC3EhnLOvyqaAA4PqZogWIk618Wm0bIir9CeHKRvKIZzHAEqjrbKt8qOlSAKxSh
mQ3Nfto7rnJWuxD4+Wu48IPE3k7bSqVW9A/fqoAveB62SwZSYLSpINq5IfS2dowQ
KXCp5UVkvQKNDqLuyhG4NvsnSSb8v/NDRtfUoqm4Gsoj4gJM50VO/KH5sBfoo2KG
UIdAmM/yKlz88pBE/rF4+sAKJy3IAxytT2YEOjC1H67GE7k+rbZ6zKEs0/l5CrRW
2sv1MrFq/8dNmGKtOEPC24FzGeKri5lL1st/7QDUpt3jr034J8IehjML8HVJGRkn
QjYPXeaJXhmax0GeloQfZgsXOFgzGTBUFuut86sa7S+numluFJFmy6qZrbl1a5Fx
vvqlRqEpXifc9h6qlSiHV+zTvHA59eL5nDsosea4kVWOrr2StRxhs+ayOF24TL0Y
RH3lRzNCyI4UNFFM5Pc6KG0z4PbJHOpwWSDgcXr+9ZY/1jtb6lcJOgoAIz4a/HDA
113439g4HeWyUiPpHhrbS0FVxuLsab2SYGrkCDYSFLri6yzz6/xw3HI8zLniFd1F
MWIxFIxzs3TvBQ5QfGpFDCWbj56iScO5NOL7wQujsRnirJ9Z/SJwU8+vNvccxeh4
2uh0mevGz3IlE6+maYp8d+f0XBjqkPmRhrpaSfwy89XMUVh875KoMCezt+vx5duP
uP3khF+jFNASDvYU1Xv0VPAxtQkdjovqITDE43KVKQBszL7qZ2Wu3FSUYUvEF/sf
QQPM4fIVfYfAjXAdvEiNVmYhyN5uiYtrkbbFHSAToQG2eltU4Sll0ohEc1jTx0OZ
TAiVxK5OFpnOC/CtHoL1yDmozDpuDBJgPZ5jK16/Z3oMFluLCNGrlUdTXVk88y5T
RoDYkzM/kXxbDmEA9LvW6ePBCftOdOCeuUiwbhJkDBVutIe0uLmPSBWEmJl+h8gq
H80Bj6OfOThRH9nNDM46oIu6HnWtePSuBNh1H6uDU1G86GYv9+X23j/MggQ47j0v
p+sGZO+7eeQ1X9wkSIvjyA0D6pcOXhm78rLl7p1imbXYlG3d2+NqG7vlOpkVfXbO
94ko4qnP9ka72n/nxBAdL/aPZMBxTVOiD5+oPwghOVxQvzUL2ElxOWzk8LSl5k4N
6MAMgql+QvzpGDQDvsR1NT7Awba91xg/s1nwWSlYl12PFHfRuGeUXm3EPD4AENai
cPtSehljXyQu/sH8PuXeMybe3egxLuLuucxO0z3S52Zdz2k0ompPza5U/PYPpL3v
IocHfy+UPrLKdmI+IPEH2D0JstzhP2BknBBS1QC6QfUS2o5k8wVYk1CUyaHVXW9M
fVKh1xFLhp/rMYTd6n+mXO0PgWosBEqaIR9Q1W9J4nEkU4Eq3bc83SI3wssRUVw8
l+I7FRPaSknwiAVtSs7ci6f+VEeTXUmXBEAql+LuTm5XWtwo82LL5MO4yWbaZd0C
XWkbOVqwX39umBt4oOdGviUQe3TLctjtTtia/+t1qt8ZfGYFIUAZDMEsdlA0qbIt
58Md8t17POmt3ijlTJXvNHN1i/Ia0M6iM6VI7jItrROaS7Er1QtzBHwGvE6ZRuAh
KqtHT9tIFGzp9s3kkmtQgdA0tnAOzTQtz3icFcGWU3iSMHpM8YQagQZ/Eh2yLrWM
gdBm534G8NBgIZ7hEMYr5rnbJ+kUro6grEJE6edvvfWZ/cK+bBpmZgAGkBnraA6Z
i4PRhEBx8rBltEE6j6qJG4kTL5EidgTunWhx9NTJDRNAKXG7ork+Na0jqLIhlBmG
CjlzKgajIL1GaV80OLJtcDSMmWHexn5njrwtkKLFaX1j5moi68v3N/tXH4Ort86V
vhCSGIyxxU1DOevtIRhkFOVttlRV2pHTeI8lxkWGKYcOiUkuxcqjmkQDSKMjp/Hg
tChWNJ/qVSodD/4eVuSybphb5/xNw+B3rmKfRBo2X7837l8UVmw/rD479bdPeN+D
R6Bq+MU1r5GyifYLCy1I+6yxBrcE14Xqb5/h58GGmY7rTCR1U0ZxnTVOyF/u3mF6
HaP7HKj6Ibz3i1GtYG8Y3OtcSbZOZdJNgWIOZBcNgDqyE1kH1dP3cUu4oai+pWcs
8C/FF0sjzUkS6OtFNXpLfVDzxgaabEZXNW0bvWwyPlf0eu3WeJ7vuU3pNA880DvO
iNy+mGjmWvSlXXHtW8nQmXMfUfTyO+F/nvhIA3S48hYtDXXGGCKKBRrynQxkMOXB
CxauTMP0ZccR9Eox7SrKyNtQLwClBOt0YuA0qZT/VoA1G5zhNl0CVTgA3Ctm6V9H
2glmq2ocnVrAx1VAHcWsaJkgO0ENwU1vCVEyzdKZDTHPfu52U06d422BYPfqyvNU
DWt+y9Y84/IcAWF9W5G4y7fR1hFC3qgxTu5eI2LGrUx6v7bIoLhFqBiZdkY6v77B
SskYWzWPXJH12jRrfh4252XuoaSc50/mVQI+dAjaYZgjT7BXLOD4/07osHgIjUBu
UD4XuTYIzyR/Nw+O525C5X6fYPZ4Qv2jSJ+AFGiLwIDQ3Oh93CsTlpm61jR0rtmi
8kOHXjYMfhny3RlpDPD6XbSWl23ip5wlICNdgpzKA5YFAnbdCFEKRGnt2YOTgfT/
7ccuBd75J66m/xNgsl0uDcLqNTDBeCIqH+YU1yWRJ07gigEPEf6uA2R/zNMfF9iU
0mvT+Nv0V1C8xQ1dTJJA7I/2+SyKe6wZ+aOF8ycRfxMh/9ecr2FR7Y7SIuwhsB7a
/AOykptgOay4fkzzdzYVXPPYKeN/I6E2srNvyKgmqIfmtFKAlxfn7KF2C9E4bPig
joix2tz8U0dkDME9hTnM06WNWeyeuJ5cAwTlb/1iYA0LyUcnldD1HaGl7lMraxCf
Umjj9rErKwRQ1+jMnx6gESbR9rIF0UneGnEeWzvweF9Dr8R44L1UhQJtKxB81VZ+
8VYQeqCEqbaQGfdq35FueghDeJK+Ycmfpy5JB15r0HugsXLapbNYjp9pJ/XPmtBN
cDp9B1tL0jOTDfdx59NnG+gPCNXOyyHYYW/5e0mK+ukY1n2MYSeiXX3PGShZdJ9M
qocRa3uD4TjECdfIafTKzKOnQ6JK3DWfmUszEMXBgMZGB80MUmZ0shSRGBTAkkQq
AtP4vwPCPAECCeSVafr94hf4GfsvBT+/6OLKKaBojnT3/GRIt17KuaEw6lB9+G0H
j8f0eTYyp6RjnfdnHikuNVBK1w48o26kIYgv4a58q3RzvZljHxzfrNK0jTGoyQih
gDdYM9myAefuQXiceTGNlRkiQUxtBHqTJtV3YuJk+U2rBPY5DllkX7ZIX++DSPfc
u294QpzwcYPiPwb1pUgc/4ifzbM5B+XKwXQLY8vLZqxX35U692tgOTDqjMLBKFri
FXfk+nkQBl2a5Zt4mnW+KZ+uwE8MphbNeaTKOSaTp3YbKR7Q9u4nQk+AH/FClbCf
/j9OCiQEQj3YoX+B1dx4CVcPga3/Yc3Pys1bHV3yiybuWqT4uuJu2bPNANtJ9AcE
d+f0weI1/WV+JCPsHH5y8Ugq+6d9U2/XC5ti90jYAXnr9bM+MeINuriWUC9jA4iJ
Spd4hKyH0TyHEP2Sm8L0tKedas7HS726falDDkRA7TqCgoyXq0ptJZuRwrCeQb0/
b97CgAU46c0tqwIJxOyQtm202DWPdUG9HC5eYlF4gLRJHZ2U7fdSZOSveOFj5GWX
04JXP9dBRr6NJ12jZJWIyYXSIbbvexMfcdwmxJ8eNnwLp4mwpoYlRrnP8Mtv+VvY
rK4YAAzRlndbBIo6Z7xyQzX0E6AbQxw5tJJof5wLCLs8OCs6ZRvUJBvQwmxgbALM
UrUhfaanN2W5i1YbnOIDQB4uMzSKK1qkB+lJgZra8/vI4o3jE4050R1tQzenZiaM
sE1GRb7dSRd6ZtoGg/KqUT27tGDkc+asS576XcCb/EVMO/d1WJ8PWVjd4XSB+xT8
dotRsGLnK839eZnPXc1t8A4WBvyQjCU3wsP27KUCY8mNXBUbYXAZJI+Li13/sFLS
m25D2gsB4H/enoVQy4dRedAl8RGl8Gj86Ka0X6ZE1JkGZzKKpjGBjiON1l4QaGHC
4NnMoWS8F7U+KYRaW7FNR+VUiibdNY6hVryhPffaaYOm1S6Zg4LYfwqS9v61MaQU
u39dLdXXQlOLZ0G3912SIZX4rQIJlItsBTH9ELc+Io1r5Y9dRwiaxzW1oqtrmXYi
JuwQ1s5oJUlYWWkUk+p/2ID/E183q0JCiY6/F3IVilCC+tpVEbrpVioC6tXB+byn
ceRn8siWDmpikWEtFXe6hCLaa42zMPdSr/Qe2cgQT4QX2ooQaQ73PeBt9R1nDSTr
L89fRj9yQp00U9Q3dKONdc2QbNiSGGZ+f4DnGV3k44i5lplRddYSavEHKTLszB3J
udNcaESDZJVV7uqdlNh5q8c/48Slia8xFAtLvhqnp7FUWzyP00tFxJ8lOCGrwqMu
hyQo6ffp+FMdWkscec1L2FMKRW8T67ZHLhNh6MDT5vokC1GCwK3vEEHOKnXnI96a
VOc+SEbo+OAC1/kIZFmbS32doN3AeTane1Pt21zYnYDAIB1FbC+p3gCE+Zv8tCHA
AWOAtLAiiBsC5RjIgVn4c6HwmztHz1o+R7yqv/IpUulae4DaoHIMfUn0diAm0UFe
C4hnIVUgqT56fl6X86pcYAUpikBNWXSx3o67kcRkmJz1a/FE7DSyjunQ+hW55c1X
ubApc3THC1B77bwiscVGskGE5RNGPmzANpAXR6QUtP9ngEZPHcFIjXnvXQj5nKsv
6iKQ9eESn2f5Pw07vw8w9Bdrc1Bl6wopixnuK7asv3tnXrcZssVrX7LQVUv039+n
eHrnKaSmX4BL4+AXLFHZlYjeStpynswunxueuL6w0CLRAWPwBldf2ixOwRAaZ9NG
zKAbw2Eg+Hah+WDU314aLFHdc9MFalKAmh8iIk0c3hv7CTsBFQYkm4qmxtTI4RxQ
2OutCTlZ5uLB0dqf3ZLgn1kbm2UPVA94YNF92Ll39sg9Mf6MglX5QPkoB5Y42Kmw
BeZ3bQ/bFInu2MUS+71F2KtPDwnBKyqneD/PGCu4zs1HaL9F3YqJgus4knFcPYmD
aZEr45EjNOIkof2h0wF2XhYrh/vh1Xd+nXJUVUhMgcN5yvyAjmGRGnhaxLAyqJcb
FiwPrjz6hXiWFxHaCNRUxU8rpwcdqYvq6EPGxnjZcoDbTR5z5esYIXTpaouH09BZ
h4e+RUoSyzoFwjG6UbWfapijAWdctRuvVeD3RteZhUJ5n1qia+jdAWfUo4xLmL0/
7zwyDEkG8BQLjM+16rLbXoO4w4S1phN3PU1iXiyqb3CuI96dxQkbvS6pytCLG/Su
u+mghFeWOk3uaRwNwmYhYagS4ZF6wv0IyyuXvn41ZtBay7PsqcAhS8OvkuGFFTie
zADpJHXf7PF8QOk3iVJA/WpZYHaBUK/EOVaq7GWlcB0tTYlbeuRqhMq6Tc0+cKEZ
z6i+r+RI9YV8Kp/Yo42YMHHbS+Ov9qa9zJLZIFVL6DePl5yVh/Hip0S35KgvONnn
lMlomLY0Us4LDxdv4hIP0TsF9cdHKFItgYRoYxQHnqiTXbTUJxiNCJ5h+YAl+199
ECtJatKgeGuoOu5hWXLtbUtpqbjBStdqcFhOTJdIdrUBNemBr3V2D7xZ2CEYn+Lj
dOUgvpxCLoU/Rri4iLfKuhYkYDIpwlJ1hFeuvXHPqL3n/FcMS5zxYA97454jzHAP
zrwu4SCoQRoZUfSLXzmZ2dR5Nbwt2H7opUX/8dlllPOCqhNIlg3H6CVv0kI7JnNl
M3vR731T3ExRqFYhc3jBr5XQZkYlXDamtFxnvTqVP8ajaPg2mOr7kN05kCbxhwOb
urHDwJZvxHX/Y0A5toQ7Y2mVQiZO7dPakQ7vdTW+x/Vuwpugo5wrwb69QmmlqYtN
ryPK/pfCkHdwQOXK+cKnJqnx0KwPN/EvzUmCSCFD3ckA0x3Pk/WT8R81vZCwoilo
9nyRc6EuubBUyO707SBP69959UpQplpPSf8CYDKGHWfUUY+xptvo/ctkxgFh+aJN
PBadn5qBtuEkxZf3GA1SQ9e/jk3DxQ6JYupK9G29Rx7gVYmCnSM5Hcqj3uGI64P3
bwPlsRYgUa7uCy2/yuLWM9BsbbWoKSOIglCjOPD5XoLMSJ7za7dlUCRjS4LDVBDa
510+3RRN255KLfSMNwKIqAyGL1tPjLP0h64bYqnGdhafWJn+PWw8Eg/XHuH3FMao
fKB7R+Qmv5wDID7188a8Rvi269Oa6utOsX4zS0xR2pwaGQd08Sobl8WZMCiQyELZ
1r8w1C/Pw7/7c/PQz9AjFyg6xijicoe43MH+ywM0lxcIi8WEuH+XUrAqPUFH5GFe
Af9C5fwHlNz8/CHd5Hy9ZHxRZfIBwBFAogrkZv0AdraS9o6+hP04F5IxMZgesN7D
w2GyB2vKY7yUs9G5Ct3aO3N7wS1D6iMNxG8JH8zIDOycdQFXFPBm5wZzoMzjMrcC
zIQLITxgNd4yj57SF3z7a1cFfpRy+DgGwf6InD0oqXt3CYuFGMOZFQixgjB5jUew
kDjY3chW4r1NfWE5l6DLD2EzLnIjrVCESNq09Pl20P57hwu1vxQmmfbcKVR9zrJ6
ojaeQXe5E5LonlpCVUhSEVn2hcow1BvOVAcnRW/nCs+y4gE0K2jsjc7Tn8De4NQe
wrJNCCviA+kUW6PSOYdABAzIDDc5ciGSLqDzkOb34bZMg+ejRQzh+so9kEgC3Fhz
GblJhKJPRB3nAH+0ZGWcAsYRM06xiyCzP1q6ambIyEyu2meobteGQnJuDEpjTaca
5bvRgbFbixe2wCOgxpDBzcmVcMTLIH0giFJGAA9FqlpzK8LglhJxh7T+0713Vrz1
8bu0cDXQiQA7ne6MhMXwtx0UwPKBTUP9v7T9rXWmkJSnaeI4Bbb+2/K5QJk8YseY
RV3MTDi0RwFU400pUpioJmcn0i4iQtJapX/og/Oyx/KIwqpaBLFScEVdLGsH29eW
Ecky8C6XuCHgK5cJ60Rf7zj3C+gkPLIN5jVoF2KZ8KlJw2HMYBaE5hqIBv+A/zCH
V0+pG2L87ErdIEnXkSYq++K+VLBdZUmg1gb+leNwkzfjSCugLftahfEw2R00iY1j
dZzbTbRvyhNhSstA+VmObJUGphykUwulZ0A3LAw/0Yi8cAPny5l+mrOuGOprMx7L
xQ/0hSauS6ya8L5Pv9DDdPl5/X1vs8vC4GqCDKpzAhODMpC0qRBbHyJ+3QoUho2n
jvrmPoiP/nj59LgV5EqCdm1mMv3DmI9o8rlLf1EsKkyb95QhF/5S0TkrmJG+Lex8
t2dTaT+giOJL5Cc54bQlWyoGrC9A75cvtYV6wQ6gckYA0OxY0Ijv3oKEXAS4dxNp
R5V0jG0tJz2lLl7i605edX5UhyS1C+m8cDKdc/+G8nBGybn7MO7It9ej66EUk5cC
yc4YnDfoWqEnO2VnJ1BOeRm1QVHVaBNFk8nRVPvyNKc4yd4wBfKaM6x38DyCY6TU
7xk/h8J5eSEyvo7in2XElSwP+mAQJpFPGSRarIS6hHiOt1RPwTZcUP4tnL0ODr71
+oPDFrX3uuItLonqDCWr8XeRJFuGwbdchx7sJHc4OUWn2aLnONKZ5SR/WOYRCgHk
7S+kGjtSJUcbkLqmkY6PDhQi30dZ9kPTPoFiifPYTnshCRV2JxwpKY7OUi4mNjbF
vMQyqQsAHb6oZSu4rKX5R/IJ8jdNZL1Se043Dyf1NQ14nSRWTsm8+IQfLM80uh1P
fUqkz+DS8+PxSenoJhqAHYygAByTEV3Sng/tyumgQMsiBOTTGZYRcm0g+bYJ5DWs
EkEVLdFB+TnFTC4lEQr65aaazHU5r/iGtkpKgWnpSfz3iAY8g8MBJBfd9YKai6QF
zu6k4DkKwE5hEFUDN8Kq/bkkMzWZADov5t9+GnYHoicVk5dno7BN2hLGa6jUeVho
2rDpEaIwJZ0Lox5gNtPaLG9yyYRnWG8XrWDwelN+45CYIW/nGsjjg5F/+4oJJ4PY
XVDWwsaRD44GmzqSweCj+sQt5PQ5AuJdTlXGmTQmp9UhpkY2d7PMG4sgolZOokYx
4+mNwVPkRfrxpHUXNoZRn+iweTNRTEUFhv8Nqtiq6is0HVDXdmC+fWXMQwPA8lvx
Tf6E9NEaDoFGkn/XpGmKQQDk2aOGYjn50nNbmgdouCfJf7GYgBWIgg7CbwiqdwOx
Brnawfz4oxO7eUG3FsraLvr+BTd3/sEzJqUm3EJGvPzn17MemZtmKGsSmWmIzH4e
jFdZoeY5BlUJdBR2eOhOltmAXE/M71Uwvlb3MJQ6ic6tfdIfo2Z2BqrxcKFzx8wl
80r2Hm2nnH/TX9HM9HV6cvTardqGKv1N+nXR1Zwrt7RVsQGpVMfG7K9o76tbtfW5
TJCFrXgs2Hp4d45i5i7U77RBeBhaqWBGtScHU9Yayd4NhEOxI6PrKbBjcq2YHGYo
VbG+lIBArhfILRsjTAxFMIKWPNbmCMqL/Gl/p/Y9wrEFs7M0+Fpo0uws+exLS7cT
dhtAQ03Z1Po5zVoVm1FkpAbCZmV1OAv3XQvHWk2BdCc54/eE77DSiwa/z3nOF3QC
lU2yLI2DINpyv61EcyzgGilzmGEVC9e/Mm9mdRS9NOPyqmix4WfcXGMnmPDkX6RU
fWeOXnwVc/QG2iyurSnUPNuwrRqQdzBXfuD0GvEqYRlU9BSJBOvVpHTzJCPZE/Fe
kDLfe/X+i7NAmNxdLvbKkX1sqRQYfBwEpB43kO/CrE6yJTjvWnJfdKrvR+P15xbA
kKzrcUKujmwWktVsCFrGvDVORwMfwcsAirXpVhePFTeH3mVEztiVAQM6QJ9Lzphq
XjcISDprnjWoH+/KF+ubNp5JBgmaNnnfUxNrX1LAQoSdy6KMekOd7wMboKlnKjBW
5V7L3cUA7FFQnHkkS+gzAiegYUNZCaj0h7NWEO262Fd35K/QfQObffRvsD2ykFWy
65iKhY/2VvZS/njQWtGaFMRWAxH2afLHggEZVvQICu9NezlVbePGmevkiCaOsaFU
73Xx69BQvDnilouuqVEm8VtlhOsKRWL2Tncw1Okn/iH6VLn7FpsFdUkMQEJIqzMj
lGMiP/Pm13fhLV21d6SYueB8BjeW+8PT+0SMCtJR7Txeg9F1uc+dnb2JoxrVV3n4
EDa9sM0fEgTjrHlfN0Vro4nPQfKkgN/LHV0QLv5Sc+2eGhP9jOsstP3ty/DNaC4y
ylYoFNqOhG0Xm+wa1X+godvGf1IGUm1w+zPJz6a8q9Vpr0I0GrC0xga4iIS2BPyB
jUtaROPYXD9bmj3qzIgDICSm7hQD6shP8xiXV0X6B1wLQ7GZedV3LsgHD854Sf8j
SSePoikP5yyDXd69WZMNMzb4vHua/UVmiq1MH1UitAZtikjGdIl+fqodnHG+h2gF
yye9cbb1O2FCP7x//+n/V+UMfxJ3DtQwDxUD0oeK/Prwn6lVqjTWUHSL5ta9f4us
Tq63KcjwKDfb2HWVJmVsY8atsecE82NgBlj6h7jniRAFHTMNdRFb7paUZO5Geke0
xZ4ea9BCJDQbH/iILJhFAKzfTOvLWUTX7zmuN9LRIpke73XHd9pD1/v3hu6EYvlS
fV0RjMuRKY584BoxvedwCM2iJu4jd2fKWOeS5EsHTp6PyYxUZc04mN55GBrZOBq0
ClL1H9qiHlQG02mm9nO/neBqqaRKhNszot8UyP7PrvGRdggk3ARJWWpx71xsjtz8
eAnI2es0yFIh/kqNSB2LAIRnk0DXKXchSiVOwc24r0ab5tYpoTimtfyoLX2CAeYl
t31Hfaw+WEPnQhBH2vPwsHMAsjDlAUMh0B2NUcz8jCc4zGn0hnrx6keBA0R/BxM+
4o60lLyJpDXazPh/K33oyDJpTEMrxulLMy/48HbF0SO5zlGTgOFfyZmSCcSVVsK/
DvGtCfejQnX6uB/Sdu6sqtw+r6/j6QhJu8gGEQkp2mRq+CF9keXWd963xJ2xRGaT
Gcj1Pd+PoBWlj5VQ/91dz3fcrNvD5gQHzWsQjbwj4bx7y+yHN5tFA0Vrz3lCcHRN
SK2vifglQnr3maASwadvNb+Kne8m8qurXcK5GD/u2wqVQq5dunCedP53rTmD7jko
8oDS1bKt7qsQ4ALB9IhuyOcl4Tv9wMbfYTgSISkHKZJ3/y2kxCo6xOlq+HOFI+zY
j/rK53j9cA8KkQxgXuGRw7cYl38i3BZSTVwyCF+uT3R1GIOMZeT9HG+E1pc29yL3
Wi0rgJGea3pMQEQlgGrJPXSYzTS3i4SVFvBxF1yr+EhXx88b5mWFRvcMBIOmeV0h
Ef7IGXCCGTsedltR5Rtg+v9ZlTqpbW1axoFl/INpU8GnP+/FATpJyVN2tj5LPoLC
N1vqwVRW0Y7U01djhed1tMGLIIkZwFD4rvuprkjtHsWb5C92slnRg6v6enPoWQR4
T1E48oT7CQQROqB8OSpl1XbmGq5Aw4JFbHE5YasshifinnqDfXg6o3jhGAVFxqg4
408uJ1jhWvF23qMLFSX4j8uIwdN55l2J2MsnK9kYtCtoBVqZWZLmlsoEbDh0/JEV
g6NHCOEMNN53aLTyDJ4lANsfGLaLOWEj00v5qhcRlFfYuHY61LJLCniqFTozan9+
HQLxyHmn8Duct6b4mJ+Qm10V9FvgsvOS/prlYvuNJvDUqNn95Y0dAOTgfwa4kSgj
c3jibHBu+KMfvj3AZVbOEnLRFgAFzqnFxaIDMTYuCkLGqMAjb04gXIHVAGYSPplH
DKobmmSXsIjw+vU4vv8iccCHdBYsocjIubRQuFHkj/Tiz096v8iI5f3dt2cZuWFU
8/Ra4c1m5jtv1+1kcEjerUxNOROOw/p3jG17iTXdvEVc3I7eRRb56MqiQKrrRvJZ
Nhf+XazokKpePc93cj58Gskm47JYZ+gfBjjueDzgXeFntEiQxsswF3VxxD9z7t1k
Md/QDP28/xTGpa05nJCDVmcTsPN97opwpB8+dDBq5WGxNA2E3nDeCBCNS1y/VQQR
GGtKmt+/V7WFDqL7WebiYiwOPnrZJJsiOwpJruXqk10XOuvr5m5muV/r79twjtC4
iycNkeHgavdacNe/1H4JEPCZOAHClH40dSaNCUQ/hUR0WXF8Bmf4nrcni/zIpbQF
vVbD1lLlNuroSUDzQhLggZsT1hImGiZypHdSpWAOrbIo5EAMnX4JtbN7X6PGwbQI
x9v4uQDAZN9nfoCZo0NF87O9c0Sn2/2ZgjeeveArLxpxNrmBNMEHrPJ7WukCTJYy
pk/2Afc5Z99GxRXtT99CJUapMvmqxwwmjLBJfgJjpt+OYKgFHJDRcw9jN3TRIpo7
IhARbr1nF6zh6hnO5Iw3QOs5tr/67NAx92Q6x97HcKFn19Qy7O1uW1sNPHFH+ZRo
uvavXU+YnP5tcF1faKZomHzZTSbUdpeR3J6LCfJ2vJS+oKKx2ZUxG3EhbJ9PzSsV
b3rtZu3NZQSHVDzVIgM50sUSa14Z4Ykx/z23Ido6LDVHMNCSaRB4LGDFrgchs/yN
ZQJNjNWiaqqqJoFlgsh9wOyvA5nDPTc/z2q9EDyqDCUU00BJvl/IN4YR6YB5ujIf
B1uwR6PF6h95FY95IhhM7IrVDv28kUF2dk9ByprLeRXD062yZM/hmrZVgyafMvx6
CQlWE8pNFseLpxcPh2EOb+x1xn20PWNI7TS8+Z27TDvt9dtZsHe5qITyV1q4lGDS
zmVp0+5LQdJJrYYioQHS9BmTRRkLX1+KNgpNO8eXb/etV0waicssZ3hEpM/UbEjc
ENBPuLbdu9o7scTmL25LqPcIxtxQ4C8BTqk/ju86KTS1ATkLRmjPGJ4en7tfs8+k
WfiErfeim0XjQatokeYKsqCu/9JTlXXMrcRCdOlZbZyLQxL8ymNUAfYJfOp2+QKr
dKLqQ9jfIbKqp5oYY2bW62j1kEh1ZBR+Egpne0wvRvsMciiFLgChsB2jGIjE60jx
xYw7C8yfgyid8mDTIOeM9PEKVKkk997rES4BOvgrvhlF6QWuVqa/4PZwIGwL41Rs
sBG730GneoAouJEdCEtmWi8P/RKWtFivLg0Vr/wjZH43OEGb5yRYAvIyVqjsYP1P
gqNv/DMBN02KJTRXrHHQRhRWREdbMosOjEP7fV2GypnGj9lbA7bsSeuBmDCK6L9C
j+8r8oljT3tAf5tkwkGwSY4zRliY7autCSj6/bEEa6AmKq4m4RoWBcN2w/zR4D+e
XXq3oboliQOD4E3wqRSomzeQNGSuo1h1e8CZwXtr7ORdoWWB9STzbNAT165RXwxD
AXGduUMv6Qqas9oNvzmAanZc2hHcW5hX62KJVWv+gwxnioZbtrUalg6dyO0aF7fP
e/vJg0N10kiPJUFSQXqw+h/N0700ks7CDU3mGbBpC6o3ilSS0Ppm+fiFWkOe3Qv0
RYSgec6P6iuKUDpHE0frpz8FiafRNkusFzLec7z7FZFpYutZ2cgB3YDM9PD2R4Sf
ngVnlMteLXVelVILm5d9ywDKQTe/nRT1NxbL/ezUsHM4ws+dms6JI7dtVcaH+1JR
w6jWOlkbY57TshthCwRd695Oom2jYg5TdqSI6/T7cnEphbD4Y1MRJzs+2SDXI+Kg
rJz/9LsSESsz8UEl3DoNotQQf0GNuIks8/xvzGrsQrDKfLRkMx82DOqyv36WTkFS
LXfp6rxaOdydL3e/vmB4bVwPByvRNX9xWzmgyCYV+HI4w+J/ftesttfGwSfJ47io
bB6/nuY6ZXO9ZEE0o4hiEZMJjsraKZiXRavTL5pZiu8I5ZWkdWbdl+iu0GS8irZi
Ehgc3fncAxnWhf41lTjJ9COU6jZQwzcSxeXWPvnwgBnBLh50wCOywCTLP58jLqdU
Navi1fHmM48txBa0a9tFGVvIG+n60e1cUVIGK5fvo/M0vS5QjbBOkSCrl5CWSC92
VPUQLrZ863IlmGUP8CVHfvTiHC5vgUDM0utnbVn6/sJqKcyQsZRsEbwqp+ksVVfZ
PsQmcjvD1MD9sdoUN5tQuAGle5YHXPmb18/GNTg2WABMMhhslXLOJmCVTFMqbz8v
QjAJEH/Sndeegm3T0BO/I7vBxg+ONhp/x9WsYGIP+eWAEdUmQ4geAtzLobeYr8ho
z4WdIC9UhsZ4JJyk3aYRTGlcotyhpTbLM0MnR6PwdlWLNUee4BOTuNO8eAUr0FJ0
iquQ7r6Qee97QZ5O9xMVlJkEfZWj32kfN3Qo8gbuWArTjWbKqavPIcPJ3HFTuncP
1IxFnKOAsw/7Z6tX9f5vUMKQvU26Z5+qkTgiOQ9+Gs7LS69NGT+vNP2SqfT1higw
ABlxEmWux6Z3qXKmDSxdUQwNSbZE7ugovd1mX+M7BvoQ7QW8p7w1aH46iE8dEMjH
ug+mTOtEgfOZ0hr9rr46hBcEOY0jrAzdCI80P7UJXWqSHdyLWSvs0HK2gOTEtFom
ankQ8JkUhsQyjPiAqYRVLmslMXekno4D7dXe0bRbTeHIcLbw/jDN5XCPwAwLGuoN
vVvL0jBcdg9GZSL5qkaOIwCBPi5yq3hV6Y1ONDOK2vh5wRLb81WTLZRD6XRp11vW
uz7umBh2+u9aWWNOKYc9QRiVCK3AOkrAHFGXZmoKItmAicU0NjDc+rqIVOr5Ghhr
3A3f5UDTL/GVYBuisKh09mXC3blzAvUK08IPpywzXZHdCbYbb4tsFU/h8NviO12j
wggvwz4ebjsysREIO2lLkYD65ua0LBo3FvpqMPw1jG6ezYy0UkJauN3P3mT1pSPI
gFqLNhDz+359yQxiUtAJkGLYL2KOAAB1dUC+D9BBIo8JFlacAOK2/M3gO3hIqZlp
Fk2E0KjEdr+lZBJn0eFKJLuDdB0kr4j/0HmtM3+gM2v/ehiyng+kDAnkmDnp0FNc
tDKcTpA4HVhIUlcgayo4lB6HJBAo4lJxYy+/OW/5ouH1X3ojO+jFlrXR03dytVPj
fyhQ3IwbTB5AxhwF+fmJ8lQHtcAoqfeWqjtWLJMgLvBM0nX0d3VoQFjFLWPl1dnf
kdXckcFYQscraZpZ4Hf1t24fMUhwsW4PhIEByLiO0y46s2GUwtUGL1lzMHNuoa+u
fb/Ug4kJlNgsp34Zx4dC6CpyUted8y/Jz+0pByJM5VoNKTw30mLQvQsn+a9gp3ev
I1Mrz12NyWmO1ivlxwSXOMEtXSvMfoRufpG//ZtytPaXRvtfgDdkY+Xao6HTQNyR
XTsuhHvp6Ycq9ru28noNsG9r8HsIbSohZv1AbS80fHtoUXfO7hHAlmbemoWKutgE
dMzFXQo5xFgchTLSW4NV5nBcf+mV0130vqeiWBF1G+VAheFEh64AB4FoIR3UQshW
GWtVBQxCL6k+bq46lesSgC1LS6QBngtfhPK52NVVgqYZwacoiYl6QFQBUhbmiGPL
1VqboQm1zf1GubwwLAsOuPnST8LgVVqrXShYzqvcHEKgJ2dMFR7EgFuobBdNFO1E
bk6nziz85ibGUST2ZUG4S63VDWhdUde+xsljgsKOWb70OTRU34BnCz9pGsPpAjCK
9mgcM4X+0ClTZ7QHA5n8Hb1tDdnzvEGwE7iINMUjVOPEtBz6Ky9McLYvTznJLGoq
bOAwwrExgV/4QQWMt+xMZObSRcMNiK62ZKam/Z1BouQDCQDf+NMHYDkJQVJ5Ag7x
S95pn7zdHa4mZoY2aRUJDe7ju++2GcMTZVU3x4pVKfRgN+OCAGtmpOPup3G7uUsJ
Pa2+HVUQ22AgoRqAPz2shXNfkPMwyVKIPxmoR4ErHLZASgIOw+Jfnc73MV263bMG
hULWTgCcz8lPGuuHGrX1c990wpZk7+B8CiAqMRfpSmQQyncPKtWYLJWfeXa8rO8O
QfTZU8Z33s6ZG82DTYcUEf89SK7PFY8eLWppkFWKEslsL8N/UcU5kHS5yRWCG25+
4dbm4402YVMNSxAGo1OoqN6asnReCBNAw0q1G4t11x13A/DwLMDsK7t9UEbwvZ+d
fBD1sAHQNnuv+QK3D7liVw48gqNIR2afXXj6ramxkr4/aeKu2+O7rXNV9ISNV1ch
3Rbkhg2Uvv2iJXL8TOgNn9FYkWGAy1Sc56NvUNm2kVRzKSucbqKjjEjmNH6MBkRb
oRojFbHnza5XoLkhx2PJSMm2a8EHFqkBGsrNp8xJUy+RlYEH2olN4KvPUclUGaH/
0jLqR94ZaxkUIoKGs0S7esfRgsxw8mxwhy2/UiE+m8SXqpzazlTI30A7Z3t0WPGp
IfWuC5sa8yGT4Q3ILf6sA/mgCEZpTamLCilAlUTxeURUsXmWCUo/kyfrQmUHeI9b
tdL/3W5iJt59WzX2SHg19UrNGXiwLBI8qVt1tMaZT6FixcwAV7442orh9oM4EA0S
3yN7oDOQ/kzmaMyoZfeDf5g8ARtnAYsQ132cBI8i04vYqGEq3Cmn4r7AU8YM48Lm
GVuQu067VYx1RBjmrJHmF6eUmqQ0yClI8Fhq1WCnjThokClUKoF7GydsXKa7MGBc
FlgMEWXwvUl5ogw8o39D0C8aRpUeYMpz9iSUCfIXYvFV2YEfNxjhBnLIXlPbGupF
pPxpGcXYZ2U4zNoZ/KAdD69Mau2xoqI+dmzGH+WpQ+/h1JdQ3XbsiIlUqxyIuYEL
QdTR38tqQ5M0C+9i9K6Ur+J7nK2J6Xo6RRuAZHk4SrMcMxspURN7/SeJB6hb1jrf
FjfJ9Q/hynxWF1gn3pi53sBhwsD5qdBz8yZoPSGRLBabl5oU2I/iZN7EIJt0i6ui
JQtBEbsuK3a2gVNa7qVW9w9eevL2iEMgy4ORYL3md9wAei9/NfBikct3zHNB2lAM
CGmwK7mckI2CZ+tcZZafYLEEl7KCfnQD0izv49GMK0yTZvQ/6Kgz16jBqisT7xLe
w5bpQV2gk6SRBBAo5AkyE5kJ2gyF4VlHErG8T9FIyRuBmu+mMsj7DY+SgpFgC9mE
T6x8sl/mkdujMdBl2tBQaCoBIiCO+iOyqIZvt9z6/TpdVuQyaEhUXXNyfcE06AIU
bZbvW/hxwUxotqvCAsAclyx18f0qw2or8k3L3mMcvxvQ0B/175vOphnBSyTwBpZA
5WepbWru96keKqr4EC7vPcnl0Ko28Ghmf6gKqNr2g7gyxpCEpSwG11kyBHhlsIOG
YzpOSLu4yC5oXxfTknThOtx5FKD7kuZiHvs51FOkJdCNTYSrEzAIexBiuO7FZdxX
/0sVx/PBhlR4v3SOMNZp34LzwLioxdkZk+gFOf1eNZt/KQsUsju7cdRGaJ2q+Vgw
/+FZ3XnF8DtNJsPSKCtIk3PwrfpM1eEchRl254wnU4m+ckSmtY3vd2eyWNXgMJ0s
K+BTKmaDBIzhTCtrOl1vhBr7N4eLAwbLj8e/U8IoHYrHDwC+Pu3Q0+A5bkeCueb1
RYDq0PqGb6g90WqyRhXIEjRJf2gqKpN6raIt6svxT8vwjnuM0o5UO9JpekK7lVW8
J8RNjwO0gqxwNdoiQlYx1M5VEApwj7DcIlwYS7SuZoSuBZiptedoGp1CDUoiPEJY
hIIzSyb4wjASuQkcYoyYXbfuD3DTKQIk+YRB5F/Z2YZM2nrqnNrZGQeLVZDA+m9r
Ruq3QXSb9h/nl7+aAL0R5igU45wgwQ3llLTpx76ZgI7dr0FGSFUrHzVYoKolTz29
BTvrjBpPMF5mZaQ60NlFdejSp68YrDTV+dZWxR6y0P9Xt1I2klEGqQvVLCOe8UEC
7f2qEhZVzsUm+RsDAc7w1wSK0jdA8HwCIpzHDkHSXbBabhAnksSwFanvWrZJU8yj
YHpVcb7RcJr49T7IoqdO8QoTAEd8aUdCGk/FP0+df1mX0I0EzPzmv7xWK8kCoBtP
REEgQAzIGtNtBBQB1+cKDCzk2360SCMwaGxXfyKKnO8qaLG6P7hmn0/0vUamfa99
8Yh3FNmJZQTKmAWFlbA6RIEP6DCTtJ7wM2Xh/RveZZPnlxQND4rVPQowh1Nk5njs
/RQLm1yB0QKl1gfGMiuWyNQ2erCTQDNLA6xDYsiIbRLVyg8dF81LI/VrdNxUWcY+
KNGGFexttCmZJbzC9jhtAT0svvSB7zclwxWva633u6rzEgRjmpT9vcPhoYBAmlcP
weYuldmo6I6rMN12rtMeDsIiO/EYNegAOCsuzbMoA8dFtRRA8c15oxsCtDRYEWBX
7FmWKG5AltL2K9f6gECj1xTBjZX4VavLMx7VdqKc3Vxaob0HS/tYXiv8vpM/9MY5
O8NLfpdzxxNs+ZS9aDizhGxEXwbTPskgNXYAZlVNcPvmRtaQ9BzqgjV8BOPsMQcQ
S6muXPxPlNTEmTVa0G8qiqLc3EVl/7RQKMs8v4n7/p2WzEor4pz8snRsqQliVW/j
/JRvyAwokJIs3RR0FSJ8eCETG3GgzTyHX/6q4KC+VyTYuGnFoT2VBD3W2Ucd6gya
/merSD+1m7a3R81sTp/q5R2f1o9a0thnCGO0eQPYzzeAK1IQyXX1lIzRj3a1VuzW
DKM4Vw0zribp2aYUSjYpukJS0SKTV4FDRWqbv5QTcNDirVMJZJvLX2vL54/jxgOU
kbVVZ2QDuM+3MpjVMe+SS19LIC1NrHIym80Rekbm2O3tAM6VON544xTRzPawGiTC
ZFk44is0M4/RwTWbk5cYyptk27V9bdMORUuoSpW9MInWqXuISFoOx+hu16msB0XV
L+InxXJPwmUm93gGeDNmYZ7DqSJK8EmtG4EEUtez12g+KEVZHjjo/caW+OW5Z5CP
iyL1cPVTc577rOEt2LfU2yDjQbM3wgU/rkIHMTjqojF1BteE7DZgdYKDMRELLZnr
OhfhSw8+C7s333KnzR6bm3A5Z0+60xW/+eJ7aJy1NaFCmwidlpyW0/uJK/sbenwF
exLEaNn+H/HrHyokWPipnrbPQnSd8hoPJIAGz4BQHrIJ86NLzrYJ1xcgryy7Jgj0
nwqqEeNBQ69igicGswvVAA2gvQrJVpAa98W3nyH6oTWpHhLkumDdEMYK7svA8dRX
bHFzYkSJERp+WKDjEHsMgj3nfm3xE5C3usJwt6XgRtXWFMvrXWL8Y3iRjSR0yTpE
UOWZzAAU8dYysVIMCeL70aW8VkwZZTOjlwf44APco51x0MK+MRMN2pPGqDkQlO+o
29za2girtpa8+ZpbnH/vro6Rcao/XLr+inUMWu0Evsf97ICE844n0kuREzH6ceUO
RcNWQhCTFwOgtPLEhd8LbKaUpyb6lLHBylCWqmGK/DMb/HUSbeuy0BPJ2EFiDtZE
DTnBKdAB7av2hF6yRrYjh854EpyeIMhwZ28cBFqtRAeDEEBNQDBYEFhrflUm3OJ8
ocWsSBKn5iPPxXULmhdG0abtfpPRbkQE2cngZLOEPIytRnqwlcWujVaDh+rFnK1t
UseSa70z9qRJ5aowsX4p/P9uEuBq8cMRj5n22r/YralvfepEAPXLKx+BVIs5I5nE
IhJ4WEhHYWv0qDWsBcqAN5DK02/Tu1DUFMKt0JDhaLeEqRDwmKO4qmx1V//+N4av
6rJKRt1XVXUiD0igKhWdCX46ZqlZxvExCaykUjKy4T2CICvQHQKVKMUQ5m3uS5/u
e69CtkPvPUuOGUtfl1V83+Pcb/X4Epfqa+6qEg68VgfNsQSSas5dGR0PuHCgtbGt
w0/VNQmFuvBBIJ5iz/dn9ZAqp0tFWjEwjiP583lIs+vSPdAbvBFM/FnfE0l4PPWg
49T+SFEl4ytsb+P+DOnwktxavr6e2kd1Z3GmpilN+0O+yNTRw+9On4tnQ1mhHYFN
AbGq3fjLZrVGQqNjRtXN5cclbmxJPXSm1hmruYpWMDJvtqbA0XxDgGKoPOZXtxss
UrmBZx4haPEU3cFqOLlT4cMCXh/ugQ+LlpLplYlRja/gCPGFx1bx0td5uHOS91tn
gzvtxV1NWwcfdThpwi6v58gf3e/dbtGeYpapt9lfm2/pufKospAXVW5qYpJzegZE
2EpOAZlfWdqay4irPDZ8cViACfVyCsfbsNb/dLE6T6VWBEhPaocjM/SxsBxdjmaF
sO7AUpWWztJgDcEgIyH4XfwQlIP/+2f2kH/CSz1/A+/Zgp2CXLp91mYScMLcQgiN
9whrFR8XhvRKVWfSi1G87QpPgyCXbn1+bdlmtfiVn6yw/UaelhOtUCxM5NikZVkM
v00lK87hRpN/7JHc7doSIHJLiQ3K5yZS3ouHK661+6rrXshWA1tqt2km6RgDXP5v
6mTO4fQDHHiGPxwnZhkx89VbRQ9FuxRPdrSTm+jujqosQif6uHY6Pqw+UyF593n7
VV06ahF+HlFxg9OvqmWpCGP9f9teE6z0R4zLY7UikvwNUswHGJRdpzgemfW5AmO3
ShysRlszr//dMkkph00JhielhJG6nkiTKwIY53DHVeDCXTXTLTGQK5VJvjNdBKVS
vzaTP42rIdCN03tKldnNas7gDDjYPUyLxHbEcOY2owT1yUymTMFQrQl3IDO3K+/3
3qyuHToAaPPbF9MxVN+VqGKm94Ghw4fAnp1MY1U1AA5hPivNYIjsRDnB0o7XSMss
O63T79/dPzzt4Pkt6mWxOKBGJ4vTGYVW1F7tvOYk6CSOAA1FbpTu0NN7padAZCV4
3typBRDRI6OTwTzcI91cUYeGFYVAiAvcKv/MbGGws/coFyAm/BTzcMgOciA6pMRp
Jq+uwiNuJ6L0AkNY9R0nHKMX80bL0debJvA9qeRseosiuOyC6p1ZD0tJy5PotJWG
DUpKohuRB6CCq/tJ8ppKTidjFPG21Fqnsd2G+k4hW7ZCF2hf2lQ+Aouo1iD501Cl
l2/KqfhXIQ+3BDk07g/pwMkYxks0G6fJQD7XMLmlHSiy4oovC/2A42oNKDY8jYRn
Ce4eqXH1cNW+/fQh2J/cBmepj0UBDE44Ad7K4BTevZEiYKh+X4bZEdLvtc43pqrh
QrVeuRdYYUeOi/R+GNAvmh/JKsEHSVnlHwIpaUaSpzZW43TtQfVQ3LGkuaOTCPhH
EYnetxmG8Bb4ilJrcWEKfK+sgbpwQ4Yf0QTKSReZSXl9mMoQLgiSM2CPpLHDgMI/
KYkyg0QBY/t2tBlQLGevhVE4AbDKgTOGyR8hOwlAy606pA0kjuGz9Z9PKSDa4Xak
B88YN+6lxoz2E9JeEp26K2tBwMP4kIATWrTQBo1eWBqxkl1zmd8SvZ4yYmeRSQz5
1z7B9fjxmUX+Ni4BrWWehUEduj+8I2YUiSCUogM4WYvQALigpNg6G8XsoRd743gk
1uVLG/8ZMy4nEHVyvk3yu7GLhZKqBA4HVw5iVivuUbJfd8p2sXTiJi6FcrMfUUZk
tU5h/FWWe3VLs9mQA8bAygRe815n1QOV6MksxGuZ8OwB6wjXEoBtcdILkPUUTiVe
uUgvc4AKjHY3NrHdmXTfpZh+h7Nw8vizhC8Dw8kovZ9az6k3/+kvJ+iuTLgUd00W
llO49Ck56a54dlNNkI22xiH+4ZdkS7KuSSI4fsEYZSDJ8VHWANNHNYY2CczT0M1A
kfaU2YJRuyagzNsjWbk0t4YwB02aOr99zpKxEF5WQa6gjWFdaz+MsS8ofwhYQezl
3W4YE6/5HhlOfBIgowoZdYKgcdB3lpprQdizEoGPWS26GWxem6h1PN50JW8JkPq7
v+Msyog/logEGwJw9gjctOXl75QT786QJn3jL74wCD8Y4jTJd8DixTf60x/XTXZi
RJjyl2PT5BvWJGfRuArJzD99gNTPvULiOW0qof3UMhU2di8BqgTleW4MI48bEesn
kXKc6zwoz+FYRMpKxKBreEifsrMMbFCtOFQDOtKac62pMcOUanuZ7Ok6zkciXCp8
uBp9wPufQqcODw2nInl0cGsPEmwKxojcejdr7IA9T4ycSn6ic0tm7DbnMBW+jDFe
Tnopew5PXdjFr0XLu7peS5IboNkfzuCu6+dRDMyd5jKUNAvC3XQel+1JHFIBzTDz
FqSC9xN7ZQB2QSy/jAENi1w2azpdSFDRgu5AT/qzWe6MPb1h0vZwqfQb/E5hBoXb
RGf7pcN/fiaFVeRw3fBV7qHykSnqmSPnUWFEdfMu68l/Td0ZAUcqEyx9XgnlX3eF
DLc/kaRDgGzriQW54Y9VsG2JtMG19F+f7qPWypuC/plPevs9kCqVa/pFpOCTOkIX
HbzJRkbqtU9JaViHpB+2znO1Lu2oSwoJ1eph511ojTrU262+WhBLpzMusfU5/SqQ
1WSbx2BuOyg5o/Xg8O++4GBzDyWBvYUVPhvuM7mmNVdnKTmumW61jOpAtypZ05Z7
5Nf1VPn8ytHKTNrOZnvac1+zm5sX1tMvmTzYl5RLxQtYGUOh/pVYlpj8u/e+96/U
w0XQZzo1y4Xe1oZ/a3BDO/caUF/O5c7XRcKvOIhXmX+OoBHFa4JnW95RrEbUu9Zt
C6cdmnsvLsWcW5GsYlcGBR908GornBCOfBI5cCzHD/eNZWOtQdC65lFo0gMNmc5+
QYBw32cLb3YU+PDCuAYDtsdBA3TmxuXc+u5ATtpLms9VD+AEL/wpJu3cVXXyZDko
yNo5v16XmBpdXZmELK3jNuUpAcCjPfhb1DxFppVXKiZOT2NVnrJTvI1c+mETRwV+
7wxcm9kM7rKXZJEUUdL5tS6KSWKOvj0EulrLtJGiDORhgcxZc+8wGy04jR7Lp86B
e8J6PnqDFQ2pIzwUCiRgSz3K7ap5LzcqRhmVQkSZwzBOPAKxCq2rAR+dzO3NDVE4
VsWipRizubnBQWjvi1XdmgpqEudPed6ARsJsU5u/rv3nyU8qd+PcrEDVxoIkiult
byPIWh3idi8P16LipkMF+8VRV8X9CgfgLmHB4spRG22cedIgPfDCS+faOAvR4/nW
g6O7+Ng2ZQHHDu1r7/iWBryvDscJ5DZAs0p+ZY6hJy06k0YZ9a34AFZt4vuqggeB
yfGe7UOnptLqHvS2XlVEU+te/dZJpfT+pu0FSHD2Zz6fXhuB6LTHaCsNwn4yJFN9
zeNcQVFswJ7wokSQw/tFBbCPU6Uw5i9OZs6dzBvTwCPRbRsw58ztmV7n3NMn/AC7
gYJsviHeHZGOsELBsY4mKsd0Yb+S7fLPJ40H5OS4dB94X+0z245gduv67/39WLbU
nuBKaIYb56ZDJQ6xAY3laLCi66TX18Jj48k9Ep4+kqDLMmnJHMPQGKnAE6H8H0QM
KGZHQd91el4/ek6dZowvRXDE+7Ihly5V02jMTv38Pwzv/yIAbIXa1KyRGADZhe9Z
Jle9tO9MDu4ssG20jogFNnlpVomMfD0fPoF9wX5S3AKqFs3DOTCYwIy99NyoQfrX
4rOdSpSDCdEC1LOMJG4PIrH2ID8rEx3tFACrW/ePQ5yDHvcIgvQVtBWW5ViR8MsE
+fIDohkQu39A/F3frPtxIveanoNjDj4otdcktL3hok+owL1MGtGqW/3UebUC3Vb6
xQPIKh1y+KakBNXBGB/QKTOoD4dkDyUc3xGBPZF1DCyGTbB6j70nmw3iWwB3U538
yAUo+2sPbG6de+lKXevDvfXJuJLh5/AtOZ63a6xB57VwIu268UYc/RRMo51TqFA/
Clw29dEGghOeavX9hTHVtWMLGgUk3AZ/QAqok1pzPLIvDevfdNN4DJTdW5cRqgtp
hnt0baRvixSKHRJ9sVj/urQN2OiJX8+6r216JWe09pBYgjHqi7egmCQbpNalyl0o
5gD6qmIMG+0kZKA1Mcs3uOz1Z6PClIpyIsUnMxblVY8XIrb/7YYnT6oI61Q2zDCb
XD2nsqdzMpQLiDzpqXWNRkKfBuMf7yDp1764gPYIkMwG2/4Dp4hTuCAF4+ExDrVs
WY9NqojpZxeVydXAjrhussL/zgSq4Kf0uTndqXO/ZRPwdvEOlPM7LR9nEnMC3dAc
+zunBbIkJ1L62Ll5cGAFDFgsopbXXRmnOBjoErnOnNIYF+3ZeOMFM1aqDfIm0Paa
bCYDRDHCP1Y0pn18xXmneyDRTERzI5jM6p3RgU8LAaLRdeYWcPJ4HS4ivnppZGzg
tq1fCAQT6/sH69meyL0XyTUM7x8IRKOMOqQutPhZWnjvtxo3Cly7fYSvUY7L5phK
WA3bP9VXHvjpZyidwhm2uruMUqjryDKgCCukDbd2eLJR5uEAtgZ00+8OKLy7AOg4
OqsCxG6xmKM5dl/geaqgNPPc4o+61CQUykw89uFGTW+eBTyRhxMM4Q8F8KqWtBt6
lVs1BxKn2J1FE/N+JsQld8m7300mocoNBOJVqDaTlat+Ev4beIdZslsjWm/vS/2n
bPW4WaJ6V0uWKMfy+4P7Ggy2km4ateJd70fJt31uYylzl6dShY+/M1aBJSqbxzcn
/jpZuQJxvl48++cXrkBTYddMrwUYoHqK8QzcnH8ZvlbI5Yrd2Y9vtg3Sw33YAFLh
ZRSouoRFsnBknqXs6wJlc+8Vdem0lyOiT/sUqvksFGswlgBU/kGrCI5CWPqsgMC5
eJdzoaFd8xbj1yh9zS9II3dnOl0E5J/jphWZeOZYRMmzl66FbaB3wv+zSJUKWAlu
EFOOMQhxs/IYEjKSNk1pCq04HGFuT1ebkzigmQnsw+KH//EbQI2nyGxbywBm9HVh
28t2lWDG4vGQpBMVY98otimOPgVujYM3lUSntFB2GBZu7+bGhYq+MOdfsVrKH9tA
uydMesmPXLQ4vi9SZRFGJUp8AcpDx8fz1PWa1WC1QFGEz16wLvR8x6PdMCwAgp6F
lkwJnaGpT97LMf6/2Dl4prkc3c24dR6v/5bnD47m3zAbvLr7UfqCB9kcE739rfgQ
zwO6K9RMRFnKGoyfytn9yG2eRHQ047Qv3ar+n45pQUvqRJKH9J0+9vkT+OPRhagv
gCxjJqJWqYpi8XrKUQxzjglMOXmVx8TaBmrpOtwhFCJqEGKKGFM3Gy9w9qUpSp1Y
UpIjOHXNrfRYhNrT6x9zevOKl0q59esQaKSiV9avBwT6qTNnW+dBmuHIxNNdj9ZY
3XG6Why4d0JQQ6KB9ECliIw2iWwOaDaX8ToXPPCFV9casdYhimGOInIgSdqnqm+N
xySWEhZjIXZyfDcN4nmzWqKI6asqq+GBHBGYy3ruyGtk51H3qLInSl6Ygix/SBBu
Qnr5453xk/nVDz87PG6EeY+/BI1PrrQSgbRSHlw54vbAqszEr38zZlMI+zvQT2YK
6Rop3bT88zfP+EOAchrsFeFvbsbOrlbUgSs/xJiXRucp2d331CRcc5wR6eHq7NOQ
FbU9R+s93yoSffX8GhmNcJeBHdRGleeuyQxLBwFYjsz7twpbjWfPEgIS/1xzMAok
P1P03wC9b2sTY/zMLYGwrU5Qeh/dItWIZ0Jc47+BUJz2Jm0ifPKr6gWyHuQZiaci
JaSM3K4Eh0tF9W8ip5wQupU2zFBbrRDzquf/3GpFjaDEL9w2Kjx2KpxnthTR46Ft
6VJy+eGaHTXmR5NjC43iJnubTtB3zde1TQKUNw2kuqkTvydUkICo8Ool6i1cAkK0
XTnCzzNwxI8UmxqSLlJc0H7QISpsjEDr1li/KWeZ6IF7as4B3h4zGVc2JHp+Qkfw
uThvTos8x6yxpU5yg4QySx3aiuIcNvVvjhKM6aVeQpmhnUKNAuGfRehdrb40ESlq
7fnlJefUCRixIR9M35xoXZAPZo/XoxvjvxFpYUiBmug7FG1E9Tou9gxx/bwujl5a
5yyy8B2aL561eClIOOIyFaCiSugIpfzQLTervGYgBeT9CwTqEXTu19NpupQeIdji
45nHp2QX5DwTs+l47bQg6y/DnDmfg/ymOp26/OjZHTEyK5cLgSlVILZu1WQEPQLH
LLGzy3cquOY3cofN+2DI5kgNLreukNQDQk/5aLgusiIPZEQhSSaOrcBIlTfE4QQg
kEI6i5QFr16NrN9s16txi6wVxdugSzb5+Jx8uQgsWZysMSD0RAEB8szhmipoAE1p
PdJf0R1AdJKyMDTwLuLMoFJXrFychF3xZPeuSG01KnhySvzlGUKJUPQg0y85kXPa
Eu/fKwaKOAA8ia9+8Fh1lEozqaM34EwItkkH3w5K/AwFzEP6YZ0tIG7n7JLTSt8J
czr4cJz5BA2JkNSVcztAA11qKpfkZvxo5Zt5hXs8SufF/TmlJnfi0luLaum7Z55/
WRupWn4ABqpOHOqRQkiVfhS60Y7KiRHUq3ktLH3huu9UIHE1kulW4a3ym/N8MEZ8
RcbhXCUp1q8ShtqJ69o90i7Q1+XwjG3dbEWdeVpYn+BSD/g1j4ZJkDay4essOAzQ
lCh8E8+QzE7hom0Srh//WJ2vZnKq59AOmvEnTMSyR75vj+ejsACPmxNVZr+qNrI/
plDP27/TZRKL0UNuiJZjryGlIL2ynrLN4au3/jEh83gTmsz0O3ulfBiZDFU+yITN
RFNx8jo7EUX8M+txKzrxlRtIdHpVAg9tRbVHLcHtEMYxRdAd1J6NQJpAuVGPHNe5
MSDOF36NoJbM2cLeGnHVYfOh57L1yUmaJSJ/6ckK+rEx/E5yb9H2+Ma+ZgQ8jYqU
iaZ5NcOcu00+nXePeucZZIbGF1JuuAAFYa5PPEOuGR4HeLU5MJKTQ71OiMr1Eg3k
aWCCNwOEkdpQxSgJ0RdFhbYMpM/WevWTWPoBoyq1RW9xCx1XvB4a1XG/9nZbucFj
irjAhqeDMRDPp7F93AGvH0m6ERJqD0JWhleRwUTJLAj9K7dxJfPdTpk8RsMrnIm7
JuTtkt/8NOXSzxgF8/cPZaCREIKMqhMx4jThX07Xvsky15zoohiA1qgbq4l+YE+h
Y1TkyIeMsriQ8RQy+QPngN5Yy3+x7XYsxwHcxYtNTT6Vdhv9XATzUc0XQ+zb8PmY
ZTZxdRyyc7o0xvCg3aipVMsnQ6+UWhSFZb1EqCfNRpwAk4eZRmBujQYMy6g7SxxM
Rr9amMAsXzFiF5bTWJD98mqGdCujTw2lhTWAki7XFid2C6EA425FuO1KqPztg9xy
9y+BHcS3tmHJa2BQ6uwTe3CU5VbZV2ud0BIwRSPUMPv3AUT4PwkFA5pFo6tQ6U9t
+M3aafmXW/kH0qJAgGRMhi1UjhUl7brbyiuP6Z2QOF5JiEWtn4tVsU0Jw54B7B34
2rUo3McTkrAcv9mSVNFr5l5e6QHSp07nkXF58CbeQRDwgL/IfQMiv2m02gmkZO+Z
SEU9erCN2IproogSB0nXpQY4+OcyE25XcQZd5pfF8u2BqDRwNzIoViYZ2zyOi4i8
/pfnd23rzu+V/5Us+zBzzB+zx83UQsqpOOGc2doy1OxINOAejZrWnuIHEb0q6cE/
hLkdnq31/dLpBicEZyfcstUgZMfZoCo6FA6ZLSw65Mh0QxTNXQmNtToWEFoTp4dY
z4ewqm2FDdsarcm70CSFRadixvR3JrBY8qcGK9cMrax5MRSKKEu6z/Ke+K1P/qTS
KbvbbcFRKRAfbBzP5ldO+Ktp5q0E+ewIAW9iXrq6+AuBfSil+swsicAUUZWXy2U0
8XgnQ9irY66GaaF6i3ea3YIfypktjOQPoPpVyMKn0vWrDH0pLs+UwzRq9g7KkZsX
Fo1DiX7QRQcmcuUxIs4/ds9QuDuuG0EQEOUzCa2ixgMXnKHoaBV5eFQbY2NL7W4i
yxbCWC3icAgMBW7fJ0jMsMB14KccTPvjjguM+IMUsgGhSljsSHuWGpsI5WszLxko
Pr0f2u/cmvX8gXf5hGh5ttEMgdoFTTnelH1J9uBWD8sjrcYaIQVOZfqSSYdDSTr5
k2VmiKX3MQ8aE+rZGnp8PRZYd0NUANipKBsjlNaxB/BuXTKBnzRRF4AwCHarK+BT
YrDxmBqCMIsG37EnmWDztGA0w6qc6pic4VZ79X2OgxNLYVysInSBq7PUyvSfrCTr
aVpkZPQvEIl2FCMd0Pt8MUiS4uRf8AMlGXFQI0lsjcebL2neJ2UUFCs8rbI/8S8H
y0xEk5csufr3FL6/m5pJZuggREiT4SF0CD1gV3OvjW7KRcZd5dvCwI8kJRWKaoRD
s8L37j4lMIKfpsElXBo/yDa5HF8u0myzPyG97gI9ULrMJzN/TfC7E+PP+pyzeZcu
qPY6kXEyb5j0zXEBNeWKiSYjFjw2BbRytBFDeMjjGnYk8iEpmZZfmeU/kgzWthL9
P2nLdjhQ9fARDI05ObF3xWxgfWfCSNG77o0nkzeHAZsuBJSpchn1FejNesNHBSh7
4ceHBgoanahm6Iotuaqa8Xf3zUVYkWuGb/grIm7MWOt8V7FxHbMaKkhaMt35JVnX
lkIwD/Zzkg3fCcG+G2Pm3R/sqjU9L9Rwks0t7zwREtKjU3WbZ6RhvDZ4ozhy77Cg
0IBiJYd6sOr4GgV5HH4NxC8HdgirpI7St9KkDmnyIFqSz1Dj0auAMAvCiNg9aBd6
facLshEBoW+Vx9wfr4og41b8/9XxP76S+JQ5lvh1YP/GWy+JXol9ZIyBICmMZiNe
YxSx9Ku5SZIfLj7pGgx+Lr7/6ZttZmRbYTnsZ4MFlGA1rBNWleaZu2bkf+Utd847
Kb0PNQ0xCPuaNDf04EEGED+749BBWslXTGDQUdsIeFCLy8hAINk2S+TcGAGHOdjL
hrJE7tjwmndJghhIv9Mz57lsbpkKxSLy1ZHkABpw1zsKmsS4XRMrZ77zIhdQxOl2
WLnOOfICZH1fvYYrHoSiBFeanFoCL0ER4Bwqfn4HBk/xy3mFz8UKAgn4DtiT8Meo
hzf7osRXs8QAJN242meLpYFFbFevzHje9MGR+WtbeUGjlvrutz2fGawS9nY1/SqY
QIaPKaRNUj+NSqsNAKOVu0qd1jXrci/ALULukL9YM83QG2e7lDwwy/TWgMU+xG2z
KpacSjNE0OUwPkiOPgnz+sFDuY5mPl5A2FHRg14U34Y08KpIoDUDBuLDv9SOI0n2
h4+6lPSzLtdOoTND7J+MvJ2Yw1vXDcMaJSDRA+YfamZMdpP+8UuEhMihwXVfBX50
kE/b81dip7y2efsPC6ChZBKe6Rw4T1hnbAIK57HAs2mx1Hr74NG7bxixrwyYlqfK
On6FFFxcBbs5nzBdm2emyyMdohuUUA/g9iB16FCfpyp3QHbvYjoMfLrb7NG7wVco
nVwGBX4K9kb+DSeRrRMjKljEL9KL4atjmjRilbvKfTMhOHiMV39+72yCIbISBUxK
A2y29X4zozVJFgCbFfr3j+/kBNWBN8DLUtmzdBBGaOlUq11r7n1zbNE842L9unmd
2WSsxNbtL94N2B6vS1wL2BE8QyxQroh8VghdQdE9JJFV6NfKJ8U2aZxDYhIsuSTK
bLLoZh070/nNHyEUC4Al6AHC2tt5JDPsSsR9cgNHp+Ef0IeihW/TNBPYetruz2aN
JBgfcEwk0mstwu2u7bominKXiI/fJKWEXNEmiRYLtny7ArkkQFZt8zIYlFx0g4Dr
xkfBw5GHr9hw/9/nmobEStaOySrpmz+PZp0GtKJ/fqpmBmNWP/PlvCimdoksAYDN
gPFMKDbqahfTjE2DdUdTH+MSuUD0OdrCmrD6PUeqhJ1E05lKGgMdG7qOn+wz8lCg
ltdGcoKjDlxDc4R7qKg3Lxzh3yr7eYS/rZAn7rp9CcweNZtqjlAuENZLdTHkTjbu
W5kY+zlug11g82M8Te8I4kJVHBzCafLKja3aweoeeR/38gsjieDNqSyeKyZ1X8Z1
IO8/W+KZJcc4/qD+F+II3LjpRYj66eLHlik4ULoxuugvuy0nwX1wwhAxUJ+SKh0m
aO01KgiqoO9G1519BeoKE4FMq2GspuSW2MQaJM01N4G7Fl4F7ee2j8mDaqZDmEhG
xMdA8ETgVKjrVLbGPjpTec0+WhFD8Bg7Y4AK99RbVIXhMknZ1uig9+yq37ViQhS8
QwP1Mo62GScQ5opNI93SCq7mWYgNhc+vZvj9KQdPyplXWO1vtbI2RgmbwIxd3qzO
AT3iHok7lYnQ0Cv8u+yleqxnpgSmZygfI412/gldbgXftIme0RWbdbtfKkx0Pg08
XSRSnWwBJNiqD5WFovojEYT41WC76/P1/h7FwURi0FR9ift6qwjm2fZg+L72DOgA
1D2damxEXHZ6h/eOodD7IRLZViQ4Dob06BdKPtc8tYAZbwMtuQHbd8Tj6T3nHDVu
gFPv4KYfsBaz9H8pcy2/vfp7LcLVoVEswoTYW4wevRFGrJZqO0ZygIRNAIu4JG3N
6ghaPbxlG4bW89pOhvo+bWIc6QiFtL2olKZSSvruTJCcNNfB+cuLzT65F+BNBJpN
o+eLWnwgBAm4w7BZkfXKwFtgNQtcQc0zr7MZj//ue63qhcPVg7Zoj/tOEHMLIKAx
AjPDMA6+3Q6r1CTOyZOO/WOg6HUi7FU1PWCNq/buD6PpMmGQgmdaflFERsiKEDph
FAeyC/faLcMBn9FJQY7qgwfsJxFyICjyUACAHjEYvOvssuJ2xJG1TcT2xOGu1tR0
G4J6erY8uN27KhmnQ/lYFOJ/oW35KbWy821eSAIi66j9wVAKE/FGw72STzHBzDCn
/YoKMUcDg69VqiIg1IhOpEaZJZjFmrKUkr2ZLK6UYyhncSnVN+PRwVesYsRZCMtl
Ec33V/cK1iFcDDlzaYwJ64MnnJG4T4RlKHFc5KgQft1M9zcdFYZ4xl/oNlpsdpHD
rGJwkiFwOTZj4Wp+XWjB6o3Kow/LMfCQGvLGQgkasRjnFY1Rckhuq9A5HdW5UuFs
ES1MwO9Q5sOZP1/qHQ6y1aZcNamq+LMDFfun6FhijlxxZspyXAm6cRR/IpNTWwpq
vKBVyjb0AZfUQyi9mCilrYY7tOPY6ItxPFRXUGVoXIRDyMw0KoeRkjqX+0kfLxqm
FDKJK/bXshYTQHvyQ4pKX9tHEuKyshg0v/PljpGSjyYJzmCkuz3F9CqyqhCAZ6DV
4EwsUoPhNlhTyh1dGkdiIctIrsCujqghIRF9LGFwYtSQCGp7lIjU4ceyvWdWd5xR
I0ypFF0kE0CineovdG0S3aOPSfGXyJAGxZmsKKKDV/14JNTeO14hG0FMoN0AxeQ3
C3SI2ZjW2VQDdOPRMzYahdhdZIQA9mYkNYwCQZzXmDYjzWnNJss74y6CKhgTGEPy
O+nQh/o/jZjq1HjHrbW9I4XSe0LEnPPwMcCyc4kTOUpSdA04jeV+5jMLkUf/BWZx
bftxl6N14e+l0taUp4ZYgLuNNEk2NWYs+sOgNzAvfI96q7DZbZQhZaq7qzaCPssJ
IXGHgWKFWz4VTCGfKA7c6pVVfVMEPh6B7fTD22bEvir3Z46ZELzBHfaCEhK6rkHq
X3I3Ol6QLppF1dQGp9Ama+Ldw3KYS8aDNjRaKIP/3UBzCtBSQoQMJzDM/guLEdZp
lgPb6UrKy8Ly2mlzSUMi6tECc5fAX4VD8qOyQmhsr0WWCBri03Ng9NdFrkO9PONs
UYfs7vzQv/Oo9EqSCNquXidxnqyWHhRwYJ/nyv0TUu2hqYM+lu5E0G23X3BqaowL
7dQojOYxVSTqzVn3CemERD8DrVqpfNZLn+kKBUdktJWXn4ehyV80QS3iE9Iv2cda
RCSPONRSF8IDK/GYRLzF+rbEr1r6NCbdMb2xq33Ju6hgfp87T1KO/8zzbESpzuel
kyeqe65mnir58+Dx3x19Xag+I6HXo91J5gdJvm7MBY5aOP0Svth2X5571M2ltKwh
vtPc/5RVPGQWm7KeEnuv9xCdPPIutLq7LL1hkA8/l8g/cMmYHxHc7cuyNP7cV2um
9BNF3Ms8ht4iol5knyaSP8L+Q0eeI5cx5rO8p2tpaTGIxTEewgQyg0oI+tgNTRZi
k/Qlq1V1BopjvVYbC9h/Es0bdZGReGiB1s2xS3vnw8yLs+cmir3MALNvzJnfEz3C
9tedKNsB+58Vp8CXUMCy/X1PESAMctpTwMUP9yxwoBh0v+4Jl0jL6s5PxJPh/B9/
xsohhcdSZoIsYeN5zTZ8sKj2c+X25sPrX9JQA0NBxLQjA3ybCbN2XtSbXehU6lA0
E0JCe5q2U2SjrdY1MWLmSvgQTVwM7nLemc7KBROSqvsF9usPPlLl8q1FlQN535xC
r+bbiLQOOS8AMyQcIZoa64yTGO0RKrMunWU/mYpFkTL5jlM/bpvJkFOF62+KaJwZ
FL+anjyYRbsIXw0DNm35SDQ5+tFy3cVWoJmqAqnhFIT8C9SCExPlqKo1HgBjJREa
z1C6AplYBLjpj5F9H5nRDp3CdbGRB9RiAtDfekV2wi6cRV91bJFgoPtugcDcwBWR
Zh0MZFi58vlPpVehk9SJUQ/CzI/x+3c0ZdpfIba225dZCk/tBSydusfuw5HU/gAg
LapncftI5DsTv9kD3QH3Tx/J2QctWBr+nxGJpiKkfjVsmXtBXOTR7BeNaRM1ikmQ
vi8U7iBOOnDi+5BmRETtSWPEvd1u37wQs1VK7fqk7hR/nwp9hiDQLSB58yXPD/Z8
gmKCu/Db0l9ahOUCH9glY0AlzorJa75oW49e1RzoUZKHM3rGqaW7UQjruHIg60L3
+7vPObBJCZG9ZAK24lsAGMJtN4ebPzOEDRv9eootD8dTEyLwL4bM3/QBSx5wuAE+
azqkWqcgYNFE8cC+fW/SL9NkrawKd7CqKNuyWG57bN10invdJ6LObBE4HAoB1qsx
RPDtEbUsEEBHFP08CjUZJsWhZwj6nZUmUiHFJeprkLOeGsMqrqYHnvevQ9S0IRCK
9DTnL7sB08wl502O/gzaiMEr+rSUB11jL4fjwquDMSMDTVWkA2+sah8qlrrNWbpD
h9VMf3Utk/JtAwunup9+sUZaDCLBvFY81JDxf3Ui2brXILF3xNiDvi/kkCSdtPc4
WA0z3wgvaFOX/gmbJTmJjATlKY+/eVM96NoYiFoJhXIUyIOi6plwKADGvh+A4Um/
9gwBJhVMQ9NyTfpkA9H5qvSj5ARFNI1awyLMx7FJ+SDf+VT3vQzQHBbCHCuGhYoq
S7Kfdcxd35Zur2nbisR8m9TccFzSWRvhfpU3Wtg+DhqugFHUBJJVU60HFrCmsw1W
kq95hTl3riRBU2LBY678DMzNG9xW5ZC1krw88K/MOziIuED8pTjo91qYXzM0reD6
0PnU7zrqljeujow0kDbPeJggPVDRmNZmhdH/qh56pBO3b4AA+M0PwUMb/28PhbbI
2QKkZrUbfJSqcnJrq7+vSC6r5KTO2NZFbs7SX87r1aRyeU1nm6e7U8y0ygZ8sX+p
O4dTTy7jtBlJ2TWBoKq0ETxjUZTcjSoEPujygZiU+LuHer9hUX+RxRSO9nEZOgnT
XT3ySvMCslQFVqni8INH7GCv++XkWMA5bcRejwemzLk5vzIeLgAubg+NrQRjS7ZC
2ftivkIZN/3vn8b2is9wHvZbAmdwFZwjj7mBCmSO9g/Okk48H4+7tBGE5nlAYp6w
dVDhfaalnHwuhWQ+TBwStGHfRXHmMhI3jODgSjnrojdQGwdGjzyvYLuI661TgYGy
YpqkXK9g+ZWhHmZR0I2uF+bZXtNGjTDQMpcPT/7UAYWvlJLA+Gqy4mn9tSv3afUK
ab7aTcop2rMwsDTZmEh29PsZHaywCSTKuUjkLph19BLmcJE6L8HUXzEtYLUCxOey
aBh/t3gx5Wh7wSe+ZRmaEoqvpMwdV+zZTSeP7Kx0wHImjKr5axgI6OGRJhVgnRYl
5HqAIKl0ZpDcxa54gkuejPb7JKLPVanhAK2laKr2f0eSl9cBkEtHvwVXBFjnT/I+
czQj2wsjk0PcfC35FkOGEHy9KLe8RHv0xm9XP82p68qk8uHVIKy/RGXyrzX0I4IM
GTbUo+OXzlIfkkRz/xFFS1fZHZcoxg9abUC8t3p0uK5CGUg+bCJfWrQDzNL2vPZY
jVdQ2xKgY/R+eBHn1SODls6m2irS43LUm5kwZS7yuu4tABiEAKdNDpJPSXIEk+3V
bjC7FWLddIDWtblvh91pimtRYSSz3gzu7HYVBCPSMdK7SrqxZFYDpCVsjNTcYvD+
CHVFfVKWLfNqBr26v9Ww0caJtc6s12MddCeJ5PCEmqktxyYhMF+E/qyg0OFEGpEp
hs6FaTu03b/i5TpoJT3/g39gY+Qo/2HM1A5LmWVmfTqQXuoLZyUB/YzBtmKnn2Ro
zRHIHLMeL5HsN3gktkdrGHlB6YURv4V2MI4oU+zk2wkck9q7wh4YxJxSkJDO0Ajy
iRbZvrX+LTFpbQdv1qjSvmqDJyqz0zXFFril8LN32ftL9rYjmX0KZk7YU4w9P2DB
ztbuqk6BlweHKykIkvP7WiDucBrYmQx/siuiUqFW4sCLlMU7lPgCyDs7gwVUHmpu
y1qm4WkoSXt08f8ZF+eONyjhhHGDub5UbvAl+YXWmlLxdZe+WwtlwKxkdUCw6OuF
3DR4DR9fkztrOhwGgo0O5tRhM15xDEE38tyqoSbm315MEC7aXFd4CoK7scAAUD+N
l4YN3/i27ByCT62vPRGXslMglkxfHysms5yFtNLMTUX5e0AeVmiI9BHLcAIiZxD/
zrsqPnThEdXN8iXwxwzjbQpDeS6vhyZEOYPhToxkRkNre5tV2J3trCQD4urz1aAo
u4xg+3X7jS6aHwgE8sJx1RZoHsMApc8UHRkdyOyKlA8cMtXMXE5/ZBDAT5dKv+K1
1i5ioN7n0jgmVlc3WRxNt6afi1QrGeqaL7ykCPEX+u5sSIove3H+hg4tEHcJD9Lm
wWedgUusSnCxiI6sOTMxw995gnHeR1aSsa+sZE2mgq86rolCk7CqofE7uHegonNG
5RJGtEPObSWmHREEbzdmIDxuAcbW++niKSZqw5J5QGo66MkCCtTQEaSyCNAkJu9I
3wFNTH+0yn9jVhW5X6dyxWri/ab/TL/HNNa9ORb/gd66cUDfG1+Nqk7yaSAX++H0
kdkFIRJTUspVR9V1RGU9ykP+BcQwZulnqbaEBd43M7CW3ErFN9Pht3Pf8NRIb7nk
bc8Tt6jTApyt/mEcvWvpYno67ixIjYOS/hErRPlySDUtAnQseQLL4iNkQ259GRY4
/FH5y07wJyaZMnS6nAybik8bdPgxngyOq86/smBcbXg9Sn2iCdXfSOhdHKR53GXQ
B0gENzT3Zs5yfP6ilBncDc5yyFCwSjUVONfHEtBxdJohE3PxXL54EanN1L//EjMU
yhZ4GaiqOAzawEXRhX0+dohblo3d6b/xiBitFm638sCCMo7Ra7gDJABYNs5bkKzf
s+b2GxNG26qYM0L0/GmAaEzCZ/8uWpy/tyAvHj9bC/FVgQI9m3evy9wlH0hFSko1
NR3+e6pHBBZaSZ1+nyqFopVH1NK2qREdaIaaWKT03ew1RBIpYtHmINHPpgktuFMu
nXV5GbWR3P9k/j9L6xflApfkEntIjDdQ1XdV+IPerfxTgDa/s31f1Qww3IISw2+n
9JmzCjL9PUM7Yfi/QSlSMUAVckOJXWDYyGf2L/lIqeVviVvghxWcnMAdNQpFGAzC
wm5Y+TX9/7HjqRLScVYOXbHW3FTU4ZS49nCoQNUwYryf2sKsikRVIQjn70vbKQ6R
aFDfmon3ilW0ZbqzZWbAjUL/myMszjn30b6ZZGO2nk3dn0ztHzf14B0ywRP7XMrV
Ce/IKb2vPanbHk5Tk0qW0xKoVQyzThxh51Mk9FZ0ldTCoG4SAYMDEYOkG2/xb6jh
HI+xlUk8GRq4XB4Q+/lCZLl1Gct0fC+xgZVS9PP1TIf+cNTasSeylcM001IpBkUa
M453rAk2iaEG8T91eNgZDxBOyUErd5ZCdJbc3u46Wa4kOdFJEckvBj3eP5Rf2aI+
OTRJ1yOQXvAY+KewE6rsVBC4eO8bTd7HuxHUrw7jNZwTYyOMsva7tz0v/5g3puZY
PVUef0tnsjXfWfjVhBOicjNd28lsRKuA2MPlzSGItwSn54TCDhYnLXjxOiFUJ4Dq
w6IR3Y62ESnAtNpznwZrTY6ShTbOrZjvwKIf+thCu9Js8nzdoCpLHTyKs7oMUmDf
gzIb3eyArxMO7AuB3dt6CoVOXJCZWO5+fp4iD0UvsT2+Se6oKrsFAs2NPMCpAK55
EAwd8xXdaVb8glUN3xAXhpNY8RAU9JbD6g9FQweIUBx937hKUAGu56y7EtAEyRgt
USiYJol5EzEqikI9wBBvM9T9Uoa2ROAOoLoQ9svV/rgmm/nsfeX/w5KCW8sdzJux
H3HZrDBMMbDQyAPO9UF1Gnmlym51mZywwZ3CZj1MQf1VWxL9EyJ5u/nUZ5eo4WXm
ieob3/8Ggq9aZuQ40a2cv3Oms2vF+y/Cjb5Uy1L06gW0bIayX0AXrOoUI08b9Egn
MaE0GseXM/Xwjm8SFSBiaVY4N7qRBXdmchdDg1dlnEt+3TIf0MLSOqLstfBWAn5A
jma8OwlkJw/4Gvyhmg+fAaoC36En1ydtQo9lRDYsIYdoYHXqCM0pcTB6ioLUWLil
cIig04iuNZRWnY4HG2sTXIs4l6fTgBzcGyDRg6RwhhQFPb9bI9Ef7PS0rhVa2U6K
wUbtukJ5OPUiRD08P/zSKCZj/XkZXAT48auswyviHGcCe9uPRpVMHvSQyN/mPTMO
mKRDx6nz+3DdLVKoxqvbiVQ0xWRfBlfO1V3Fl51hd/6j00kwuCYZ4wscqo7tkVS3
mh1wAevCARBKJJxCShi85z/qxNHpJ0SACVdkI/jilqoEr0gvv+gONShaBi33zZnv
tnVW3kplf8UfnG59DQLVMP/YF+j/yMlEpBotk72hhHYjcXBTay7XFvg0YYhiCQFt
HQko0GJR4Siqk0npHckvGDmiU8ZV+3pwY1gEpNEbDWrkW3UQHjrJ4e9idEmbpEsX
tu2WPeLuFrigY6V1kfMNGn+7K4KREN13rvkDBrJX8V5WV3UV7P3B9mUHgFYmwQQ6
94P9WBvLn7OsT00QfNdeOP6hPJs9LXPw1LqJG1wa9TI/reQIB3tQwQOdO5A3Y8TU
w0ZOgYYw4Cf7RgbtXtXlHtRXFVmG82C/5fFmoD1bYZX8kqE1KWy9PDmQtCpkKRSD
VH1+/m3PrCkjBgPSvMAPOcweLkG8o7U9K854Zl//Lp/iG2PpY5a4mlxPC5MM99F+
WxPYz+qYUlu/Aq4ooC9jnVDgoIS6NmI7ZgMwXyWVgmY+gTGTEoJplX2xrsShA+Sq
ehSDYYxjaMhuxxRVBspeOhmLDojxswvUCwFjsc8be6j9gjdKjvcfTnTNlckmckuj
3dUy0e2/lnwDFk1MSr+hAnL7wa5vffwhf8QB4knVE9wJONsA+9+QRM0lGNAZHejI
qRLacC/X7uoFjZ09GGa3u4P1gcG8WbDc15Vp+jzBjAqOY1nWd6o4RXteeU7+6Kzn
biqzRt5hSPG+mBxmo/ftfS/JlAOYJcS6QbJyEQQOEJ5hPSZnyWYnTwTY4R/96PTd
`protect END_PROTECTED
