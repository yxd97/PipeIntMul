`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XDozkt1lSYwr84vxuyhbx1lZzjv7uzQlGwgWXw2/+JfDcILdKM9yI9OojfZEHR0T
CzfDookDiKwE7mZ3w8xJocLf/KcCr6fiDV1/nAfEfklJfwm18wuactEKaXZycjlA
hWBIQSHCl8orc4YVzk7dvuz8bLbKXrFBrVJW9Szbfhwe/v8yhajEIJuF2ZLgVzNd
7fjqAZzqhOudbrwv76ZrYisNPHe+Q/dEGeJCFS/l2D8otKwDMjjj7wkK9hkVbtGu
0/pEQqJQg8b3+woogTX/8l2lzyW0zty5/Jte4IgSDHha3tagb1Zof8J7x0QmZH7z
Fn6LPVosFbCRMFaWXny2h80/qt4SmiTXHHsyDLXSjFyufJr2Jl6VuSkHaoMnm4QY
hM70TwBm3RR3YLBVPzcZ8QcEsbyYveKuTBoL67SwFN/KOWr+a2YPaTGJ6kMBy1bH
zswjxFE1B8VCewMAkmg9zvUShDvqwzfvL9P1pW8D/rFunWNCkkn7Mdc+JgV2tlXf
msfiqg2563Jj3wrOef2r+92USRIWMeKHjy48D89+IZm2DpdIbvfIQJAJbZT1aiCx
OS+RvLOKAhHQ1iI4EFkpXu1aHraqlRojbZ3EkgVcczgTmcZCyFlQGT56ax4w2uFz
pXy9QPz1IFwLYqBCzLZMVQ/VolWQ6mfm9K4D7PGQS1/OoPLudqAT+HcuE2OAInSv
5znLM0yWb/VY8ifef+vXqBrcUXyudqj2R7QJpe9JBejKaUnwcx8XnuEFAiVZFhFq
7/W+3KRE8wBW0/6kAsj88KpgqSquWy480lzQwgN+Jm54fcOXo12z9adLqZ8qvEGS
uZje95+ROovOLuQrtswcF5DTdyBF9ZvEPmVhy5xe4BeNkGxyV/0/euTRusEWGKaV
PmCZ1Rn98yV8NXqbQ2GGspCFQRX0Db0aQeyi1GI0r8TELTg0i5emFK12KKWhRAup
3eQyi9gf9LQFEERoFf28llklna5nfib7hl641j0iRoLDvK1h+Xfe7aaSUe8ZtcSj
59fkkh3/BHZlXHx09pYq4k4tkx4/G+/W2yN30wDEar/A11Ykjk0q4GIjFSvGZsSM
tVfsiMjti857tvsdcxTTyGunou1wGHefH+E+q92JhvjyY6J6zJ7cbxP/gHWLhxSY
gkFGSLF5o6OSwM4BLk43hI/Oww+HHvb33/0eFbPVxKiY7Bx1C2vgjUwzqM9xQwmB
+lu7lxZXZHgNjuGSxBYEJG+GLxYBhy33UcGtLshcojO9AXsaeRhIip87RtPyYOGo
1Y7Smv9Ew4mCTbSlt+2NWxE+Yn2k+gemyAlvXBcY7ZJb3lzjW6mHsktmMuYqaG5h
3rCZdCnVFmp/08BwQ04s+xkWie30sjXcA/4MR/VGBVJmldSY715P9vtVyR4jdYwy
K0fHThVtz9VaxEkYh7FMJlpWYEzt+k6/2fZH2qW3s3K2wtr7S3qKr85UQbQBqFF+
IZUnFvTie5mVTIo7e5492CtzIu5mJIaG+ojhpV4dV4ldnakbcu2U730dZOtgIqcm
CHuQ+8CAlpbdx4W6WAJVrOMSdYuBtJkfzxFy+z9bmOisL6JTnZ3EqmbY6+yzc061
qS2qODc511b+NEiGO8ULOGzL8or45QX1ltXAwNzAhvJkaPd8l1YI95SOerm7zPkE
r3d/3q6eLbmpfbAaB8Sdz026s4cmoQdYmdVZXLmDnmuUF2VPrtSJwtY3ha5LvMXG
eonTDv3O5YFcdrjfGwpyPLDTnK/yGPHERZEAC6L2mi0vBzzjfrJRn2y4porm3f/+
ECJVfP5NrPzOyqZ7nKeJCpG0Jk+8feiGB0JcyDnDhJs+whqMfdODGXRzL38uNNlQ
/ctm0/fIqeQIImqfpx3Unn7wtrf383sWI+slYAzwBLIRgnsvp/2q2oGqkyESF+AA
1AZLA1DTIGsdZCa7q+nUpO+xOUBMxfHjRQSrfgazftwuIbrqEfVdCODDgNNaAbMe
b7VuknGC3mc6QLOdL2+4Kf8N/xIZFggj/pt1JcrtEXa3roSGMOSOBXTtsPQdlnPK
Gx0AElGVX+8FvqfjdUXrSKwHcbP68Pis8vfBqqUjVY4HIQPPpcjP8XUI7XuAa1WE
NMbQd/iUqkw5h31+QWS4I45raUGFQ6iFbN6q6MGcKr9OEoT4J8Wtst23/6JzwXa2
x6IpMWm8basYPaJ0Vgxs+4pAN+jbuawwCn+vPD5hfGLStZjQGyw3tvzRlTPqJyDR
WRMx8MFMjzBQ3WgNirBV8OUaBsAzFWVhn+zpBKruZh7bqAQvMQKU+M8p6nIaxc7Q
MQnhHQZ7d5jbSAuuimGFBx8RTb7uTVK8b4xS0lULCSrWWGLOWY1J6FrpAvYxdJFL
V9xvPOKhTjASsCHFqOjvkEGHVN6CPQTnD3tpbl7VbPu3j05TUP8D5dkijyL3ce2S
2WzAu1Uznotb0k4RmtPMblG6tRXLCyP1DuczKkE4U/0dqvw1BNL5Ut710/7f6zYl
kw/D3xqGAs6ay5TZzGAKc2Ylow952kfRNwi+QjVVdG4=
`protect END_PROTECTED
