`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D6zkx09q2/urshixjt1k88R2k1aKQMd9hJ5RS+M2BOAu3oAtToZxM/rjNKabL+tq
KfBceVQSOQkNB0OtXueiMCG9JdqlbOo5gQ/M1YlHj2LSO8/qU432Qu2RJd6SOFZx
B8T5NRWeW0YuIkvlErCVFu49VtDq5k36Xa/eGXP8vr3oxqRfDzjmPvdaVrVrG6qt
uN8rs1ds7CVPfF4jaO4IZLzo3QIDzz10VCNpsrW+LZ9SS39G7CqdvlQt8wAXHwLN
/btogiUPBhKO3Ld23WhqkZ9Lz0/WrjQjScLDjJJ4a11mQ6u+VtjT0Ik2CG8xpzYa
3WFXoh8MO4uIzrDDE9aAMn3DYODRviYw+9VnkIKMpE52KgNkrndZLMFPDE8++fzW
Y5uuELr8EaW4b4vbcUBZd89Fx/QnTNgAo4f3RbiVz5FX3/C7Ei4O5SgH8KlHCjX7
YGYbHPmwNCYPQti8UI2dy6I6J22cH8Yb5eXf1npV/9E1ayamIlkpgLZNf3UOyc3z
XxSi6SqIIq6ahPuWk8649A==
`protect END_PROTECTED
