`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mAai/E0/kBohI6h7iNc3oeYJ4dMRKaO1mH+u9EPZ8+Ezs7J8u1yg+3Zh1RePNiG0
SrAjmlYHM02DSXgD/y0VwlI4r2x71ir6YXk7XqSIoFipOJWbO35S+clH7v09wVDQ
qpSPZDoKQWY9vcv0GmmwoubCIxzK23C596Oz3eAiOX4nj/otVRtHfacWPDZQBdw8
UFNeuM5amMfxFJEqJqy3aQUViHOAJXAmyhwVJf0xtx2YhUjuN8MsPAA/vZLAEedI
rBlVzGALaQmOeHeVopj7PFTFdMVbkb0LilZzk5VCbATW3WNrb9UsZ/FDk5uQbo40
jtKLbpq/KJYeyh0OyNjfSG8Aq7dw/bwVs5tOiElSNDWgB+YjzGASgMKOATFuqiZ0
YMfhtLUFRPr2G8ZsL6RGbbZTFZJ9xdJ493WjkGo/dYOGveJe3SamLP+88r9pRUZj
XM7p1Sy9ciomYiV+WmO+8IRJmkVlKoih5+Pyd8KVdpjtm1J933BN5wsDGZqsknR9
6WKvsuM8l4gvYEYxyN+n6Lhohkeop/oBXSkBS1xnEISIRkb3McZd14fWJjPs3RuD
mgmbuZaMHkxYIAUi/y7kmE9gXXhYqj1YvZ9KhJmMZLYjUccXY7Sxw88c05tZOpBl
nfbkwSdole6bf42FMkNkdRgfuSPYkfFX/tYoDW+J8sjz5vGz8XYZFijMFlBvD46+
bg5rplS2MFsb1jkdoZxWjtGzVRi3HIRQu62vXGF+pfuykaFFLXJKHAKROU0dDJNL
KuVC5+NC3br4dpG6uTA7qQAtq4ouC1U5wsfA7sK7OH0az8D4YFRYYoKJ/qbBptGm
OC9iljNh0irWkwtpgVQMb8Sfz1IC4W4SF/F3m/z1uLSz+VV93PxCpFtYAVG8rG1E
lVLR5SZncrVycH/YT4tRiVxpbTL4+bhsKqczlT6wYd5aoO9JulONuyPN1tW2Nna0
6EA0Z2aqJmIn4tPosMaI+gVYslem9IF2fKx8zVqJw24KytnWNw/iHcx9HE4LXygO
I42cswJ0ZfXjkzCSJiwxrRAe0Mosy+iqs/BNmYj/b17oNtSWMd4/CBuw4fJ4sePf
4Wlx8heFfjPug2X8vYfOE7YfMNsTJYlapwN/dFfvDpRKVNTFpXum4l7emqeTECmF
xOBdmrWpSJdVCOGa2mnIyL10DrI1hCJUqovVjK3bfRu5HyUdlBASPg2aB5wwCuTK
PaZuZWpoAAK4NHsurjxOSqthcoGkTEjM/HdbXI/aiLMWKZSvoagk7u+TUbrZElQM
nQcAIYNrXCZGOYT7aJu5AZ0zxp9Zgf/La7xk5zRBNJuo0+YJM3yyBmzMGZgSOrPR
Y1tRtB4kEK5xHIrV3qIes+/BIBowvSrv6K/46CiANKewNkmQnzBsWxnKJ1ue/JuI
iewBn2pyTzgn14cYhxdZRXbQsT3P9At4yhe5QmofqRHNMEpSKDRK/5pB3RAARsji
+3/kK9Nfz1kdLg4palwacIyhkLFNqcsPcXKjNqMDxzT/V3nTQEQ8j3f5RdFGFmBq
b1hpgCvIwsqniaZvvs6ZLqQ3TQPUKi0niox6sfLjT8E+Iz/SnR6SsA78yxff131Q
K0CZK4Tc9xacEFC5hwASzCT0Yc2gH/oAJ1YWKWr9s+9DoWa7T3iMlS3mvwZeVmSX
`protect END_PROTECTED
