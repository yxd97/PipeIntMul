`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xxyd2jkXtJ1043OOwOGEta3HxO84D8dL+tYPFaJqmLceQ2fuJH5LFZbLdGTcL1Oe
QImvTkadXsv2NCV6+8UdNt7ZGm0nUPAFnYAtQ2tRtak6g4VHV6KCUZ8298W6ik3s
RiVkCVjkoevbvIYEsrcslSkqR+c3brE19rhUbVPe5+/biwyzgwGS4WoBnhJdfFaa
xnGXnH1v7b/dhOnJDTtflKcvFLgmlcvm/y/Ly/7n/n+v9/PuFlTfQ5y8nr6/gJBq
gQpL1+S5o25IUFT2QsQJAQ/PFeQwQoyBZrBJARCs80uMZApqSZ7xVGBxdEkDfxfa
DbpnhPQni3kovGbXmo3Lrwt9wOmgTjIU8JGYs01HRQds0WQw5PR68aVRDRe6SPDa
pHcf70oRE27MlzUu1hN1HqYZGHtzUmEh4mVOJsDpjSzmDQRn4wKtTToyW+/+Ucsc
bGUsj0kztQUwXQ1DkpilyCVSOSZwISgIOA+FluPbXS3b4gMDtg3XuFajq8tlPHhD
JBZ9s0frQBGvRRHtZgzqI/yKckq4xuYxOV42FivX4iQc/4Ymg/Q8JkuizSpD4mzd
qz8Tadhs+Bv+ix3nxZMUqxykmEd9mv6178poh9qw9DBXFqIkVjeGmJwfthYYSiNg
Ia1LUgZg/WYkuARH4JzpQK3hKo9Kayp4YMqJbhyrJKTNNBly0Dqu6whir1U2qdol
jLbFll5hy1J/K3xn3bk7JYrkWR9gTUQ7o/VZHovEFb8=
`protect END_PROTECTED
