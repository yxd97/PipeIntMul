`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0obTNq/fcDDaSHF5v8Ddw54iU7LMn/rzDAWclWmNWUbq/Mci/cp3g7TMkFZZqxZ/
WrUD5YP+QFLTLLKZ/QlkExkB5Y4jwwceeGyS7USmTd6tu7hEfcGB4BTeRGF+FIGc
4kEOrXlEJyP2pvXfQkru2uVsEaAgzLf3LjhSTIeBz7/qf0gfLORmp7CWBAZMnTBV
bZ60mDQg6YAx1D4e0zfXIvu94KqRqwynR6S2Qs95P99feQGjDbiizLWKhiDGHiIX
C066bDFus7VPTskbSbXWX+fBamQAfvSvBa4b4MjIaDcbp8Rx8946QBHGdeMDpNTm
d2JwrAe1eCzlh9xb0ipAKYFTTRN4i7Gkh2kegZUqeddW44ge5CXRFNulFZgD7QnY
Gjj3TDpLNLG6lkn5eEq7yE0OZVXin5XHaEp0qcsgL5cfTUu2rAuk1zndPscUaM32
myugEz6wY+iFFr7rx/RqY+ZPjVhITzwcQfWL3wgs+YVxzsfMv+uOlQVSiEfpEBQA
HLz0itMIlhTsF8OPvSC681+bbnP5pVKOe0OLYcvEKVbc0Npz/L2hwRZnHcpeHibo
Y4N4poVRYmbeZUfb8R1ePndCwfk7LhZWiZyMCph9EcortW/2dO3XZWt//wgaXvhF
sfVY6AnMstZlDc42d+NXuhNvNbBtKGJn25MUvIlSdsscIl0m0u3mtOHNJ/txBIWG
c6Wm8CHGkFu3PwLTnqfxCIR+6RjI9uIm8zXldU6NHpe8X61TSgZJceQjUmfkvzrB
5/M8Aqj5kink6hp92HINunsEZNvQE9e2cdx4A9anp67AAI6GlVXl6moWV7UyDJ7C
VSYZOYex3uqDjNPX1o+b3tJIEPvLqZP9991o6FRfN01Q1QBHIj4EnIJwNcLJbS7M
cExXGOlRT/hW78+3VHS6URWlzZ/C4OkDln/aokHJX1GA0qnQRjQwGKIrmF7lKYmt
CZRENgvOxbIDrGztiETq1KTiJ/71PHesWzZQOtwCsveLV8qHaLU5jtZhMxg748la
O+gbmwkkDggGTMEx94n2unlKz2h9NkmSGV3OHJSNe7ZpwcaYdVufYETY2BEt70kC
`protect END_PROTECTED
