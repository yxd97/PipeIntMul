`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sFSd6bjMofLTgkhNDQDud4cSiKRbk5JnuV9abNlnH2nEAvdP82sPERch82z77F9e
nHbPoX8cokJu5XuoZm/cl+ik2hUHRr+n++pER4XZmkbXpmWoodFM9+nqBsPycg+G
c08mcj9dd37REEyTLb9QTuWkK1sDz37usYz5CPsPXY/VF8VFo240Pss8FE1KKMbS
2owTVARHRqrt+WYct2+Y1RUk39nhQPUzuYqGdMyKj9j65ohRyC7mCRiapIfnNroU
ZohGsHEAD5hg+P8Q+51/SCUh257JsBDPoR+YRB/ooHmImIIhjSPoUg8sJIqth/Nl
R4GQ9KJPf8JrfIBCgdbGxLLrU3lxY87ypUrzfEUs4Wq7jTmC6sGFwLL/AbSWX3x9
b2gaSJlaCjKzbgrXS21j176QOMonI/R0tQcTM+Yted4=
`protect END_PROTECTED
