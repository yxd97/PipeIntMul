`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wfh2zATnX8TwC8813hiJUmB50jx4VDCHuswrgss4VazizSpA3oFcL1ccm1/jIKZY
iumi1ylgGpk35sUt15rbmBirMX4EdNRUUGulfm+Mi3PK+LJiFu881gokQ2EN2X1Q
+hnnyIwBPfiTvO7bFCQiFH//pZnQl+VWiADcsNsVFDl5cAkmg2BYt7i9b79GO2Ce
p7PuiO6sSUEMjEZnQs1wxSZBGMRmayuUBjy8ZyNb9adf0791fXAQS8CGHh44+91i
Cq/ApoWyv+5sStJTvEqXXnAHNbmj8mdubZ6GQGMcQRyjqnIr0bOMoHF1cpsID1JT
aO6ZoFjHh1JgsY/CbYCuzPGJIrDe5Zq9GVeLQbkgc6kGbQ9Mr8H5DyL1oapaloEH
lezh0Kb74ARePSY9NUiVsFH+e+3MRRAGwOmoGSiDtTB2DxfKVgmMGGLHa45ushDP
`protect END_PROTECTED
