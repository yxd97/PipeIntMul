`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tdV+qZwvHbfI4oTRvdIGbOCRGGOva/uICf2CxZMolyX7Ks19ksYsbYNjgW1s+KQw
EIfli+Mz5MgbydPeiyhYLezDBTfw3XxnUS/rdDrHh38gYKY4JzCVUDpqz2hChw77
+xWlbwC9plImCTOZdHc0RvqYycC9p3HSRrwDJyGV4NrUJOR4UvFlDrUZg1nUnTJ5
H02U5rxt2cU/4PoyvYpDrwfvSumvHVq5yO1mpwJ7AXYH+YeIFPyuIaOBLag7dcsu
9izRJcNnLXdkdB5sGjrK14zBQH9egjZbylzWranOGPsVCfNWCcJ72p5rKeWa3SZR
55wqSczE0f3iuJmhMeKalw==
`protect END_PROTECTED
