`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ufp505BaggHrgRGvKWIiCL4+XUKnOf2dvb5anQ2P0sKPrPQKW/OI6rGXecMBlwC7
FEhWFc6N+oZbs4G5DcPCuORHu41wkK8WaHfywWJ168KbHOmZFjeVR8qfMOuhkxw4
mP2EJ5dtohC4P6NXDeS4d5ouLJ8HJGWUqQg8hjMkzPr6D0JvyuFa84Cl6qYI4HWF
BNbYVAQ/GJjyaMvJ75BLkmK50Z1NCIhmY7YH84gjilBeuxKv/k7xkXXsCRRK/fTb
NMLHcvx+4D7nIJP9Vcv6UaP1KNSRQT7DVMm6W+mNckh8a4C7Xz8pg3vUjgj5ShXm
BSjHrykQIvILOU55/lGRZGGzUcrRUIJbv8JgZryoCvzBgMIj7jHwTnjjeDdbIhxW
TmSVFuXH7ZXvO0zwAsSHCKoyTtYfR9tySFWHYA92ITYcwP/P1aMpQu+fmLPuTBxS
uYzRiV9lMi5Sw0SDn0eLfcfsFBXu4y3NCtLh4vVE2HPgqq2/+UXd7SGWSnvyB+a6
C4zLRYCURCo5GqdMX/Iu35vJr9XPCLGzQK0+bDlyE6Fe0uQBH9Ye0knXr+4oxh5K
ueXTxLtfvVh54c+Ad2TQvbOqKrBkM/JWm1ZXhnNNZRwLrOlmvYr3KlvBEtsqsfYN
ay4306Ak9+3JpwzXgspZ4CD9ObuG1KyciFcX1VCWhhMV8Y7JbmXj0Ag7fdjtH3yt
yAUDCvk6yG3BmQdWURE0aj/pY8blo6NqgP3VHQDOPzmEH1vsvWMd+OJfqPZ8/v6t
ZS5WBclj5pnn2wjWfX9r8gT03RR7AW12FA/+IODFz/hqxftypneNkg47Zfs6kM7H
MV7z0FX1YwLXBqV1fkUaQ4IxzItfrnb/WRxAEslye7eJ7oi1zFjMKT8WAAlWX9+1
+NsJD3BuxSJGMRURrpcYL8AuBZxIPcotQSwCKgwrdgPFbfum2y6Yghyq4KVdy2c+
jnlcALc3KvQzYkIqvGM+apIYxVxBXNOzic/5U1MLY7kbN78twTZVj859EHG7Jwj1
KObMjsr1OqH4kTDq7J6yv6cYcwAqzQOQ8L7bd67YcVR3KhD/1Bxl9vZ44CYsJX2u
7SIyaP95uZUXyz9PNM0M7rk7IVCsvlizWLZl/Goh+enrCJxyGbPvqiNOeLB2RN/+
Crx0sV51AF7eNn9X8RvKf6aNkz5OUpuczwwGDuRZyK509VtIirUbwNEXPNgRLXRO
iQoc6dNI29XTt6xqc8uZsJYhzrlsnw3NmalMlJMsm7VOnpzMCyrdXQfoqns2Q16H
ADMxb9qKQ0cOUwHaS6sMydYdeHIenolveJj/3ZvQH9YYcYmg8ZAIyD0xrpxOGVsU
dQc0hNqz0MZLezsavI/frh+8AI0s+72xkNbZynnezsQjZABYup/ZptZOTA2Z3ssg
2rm1n0NJBIS/2Dk9jAAEC63EkRnplCldo5jSiEunY98LY2iVzk4aCGFNH1xg7jeC
FLP3BA048kE4KRPJO7RbAtBFpPAp2GS+dQ1E3tzGbCTIzSz3zOcv+XQk0EIHiG8l
OxAME3YJBih7/bHxY6qpJa/MODc2wl1FW1PuGaZtyLOpk8LZ+px2UBN+xYdlo1Yd
rGp0chSAFRqVZyHiTxqPcWW7MKCbj5p/b1SSbZuNM1pqKKXFeNTNWOSgcaV68+zM
ldYeaqbWrgtWcvgkobFvAeSrxImqIVqaOEOKVv320UvNXKhAGq2evNAH8yCc4zZI
DLV85PnOcBn78hR9IZ6y9SCuxx1X9NHBAgiwSTdwZu+CgfU/ZeqLgQUcAPWH/opq
mNnSAumK1PSSlLYdx15uSduRDBzi44Qa698+GccRpuHu4JtnUSGwKMlc6nqxqlCb
x873dkrHLTZIRHsB42NzMSvZ9unwYwyEG950xVkl/tcfyCHviQNb7k6HdAIzuQAQ
AN4n1hkVU9zFyVjnWqXTfw8qIrhVjOqXp1YpHNSY1VIlTziluUYROMKD/DJ91RBr
vNY5WBnmr/bniy4adXG08VG5rKYYxlg2isbKgJHmJ5c=
`protect END_PROTECTED
