`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZiGr6Mx9+c0KePN+bWGvKG9iVDQY1EC08ThYRgnpWKGi59uW2tpiXKD7Q9xsBkS6
ak83hh02kMJAatkVJW6FKqKhXooP/g8bCW3EUld0TQnvrUJK5BYnWHnib3EMMkvm
P3yjALV7B3V3pe5TYgUCxdeed8pMSq3Da8wZd6vKMnwip/cCAYJk5GhIo/+ZLe+A
m/DVKGeUIbuF0opKOJ2ylbQ40IeSWoVJF4tpniU2/AK85rJZYYc+evT9jN67sEsM
9739Dk3DtJiTFyzEI2GoWW07d1bNimnRmiiUDH8limPeSOExduYjQOPJITFx4it/
jzqAbaY32IG2LUccS94ueh7I1VLMxQnmWOBS15eZx9AcRYXCrQyEgu3UFiI/LrGh
v7Ot525+SnpHG1dCdN5fTOtaHvl5WSPRZh8mKyAvimLbG171bNcMtciBWCAtnhFx
2FaLQqEBkWsuAoKl6P9Fmm5eBEPdzk24QJBoyYAVgTFeh2Ay/3mYsylU8KCiJfJV
3NApQPzF21Ay8MNVt1+FMk9ovc1eaqmNI0PIuXOEDHRjS0/8QOMWqGXEkOqjyR31
u9fy+NFM5KYMlgNQS1WmQodQIlMSKYVknlltOBbm4Pe7Bir0Sye5ftfIb+7HYPAh
6zEXh+PPOpwtLHBeBWP5K0SofKEPjWR9bgmsQmGaEmKTVhLiXZTYV76cpbyDWA8z
`protect END_PROTECTED
