`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dkqb6bHDKNwANBO7IJ8MH51TSDxO9Cqky41lLaz5NcJwyziq4WZieR94lVRudSNu
fpzOgdFvz4RqUzu3UqI/W6sRE0Tmc9Wb8fEClsUcyZ3IKvF/tqJD7NBd4IQOQZqR
seT+mwyjdXOiLV5UbBThkK6f95rV+DCjM15AZSRhLso50385HZtb2fz0GsjKcJ58
a4L4PBDO+ryRYq6wz0dloJbd6UJHh6wruSGu1NILbMnA9MXiCp8QC/rNEm9GRks5
/g3EFubck9m+BfNFpEDh2M3lGANmAHAjQurOeGD9TJKU7KzbVBCcI08N0+htT3/m
d4BuC0YZD05dWkQmQwpjktiiwwxJ1x2ZAL+Ce3M/QiXf9dlz6GbN1gVTxGYbROuY
ZuXE6c409JM9Wq6Vw47XfXoTnyCPxhroWEF+fmkFZgHXvaWcm1PoYFRVDkytTCvn
jVV5VyjyHndVPn2AyXoAUBW+N3IvNsSMpu1pAvFp2FLbMjXcKPNde5Aytf1fnY/E
ritVb5z62aQX4GIXRqZGHutTXGZBbGd4gCBOiVUrWS6I4cjyeAv5XAFfgFEdY+8W
/tlbqLrfeF0dWzBriZ6zJbdUg7PaheOAg++D/XRUoB0kmqgFiNL1ePuqiRMbWUFW
fdlfCN1/MeoqtVPjhU3qLZcg78vy8ey4WeXxjJ24/BOa1Jo8Th+UxA6WAkXlfdxD
lj/UriYTgbOY4Erp4vnZmqhs8MBIKojAAXXzztyvIjJGRkfPdsEVGbFqXbHy9rXk
n2tqbSDRWYx6Zvnxnx5IpdMad/lMkpcMlZ9lMOCnEoQZO5bcvECe2yIOchdNJI4h
AuJkrOMy/N7Ktaxa0F5S6D/2VGyO7lpPUa5lSoPBhwxg0DuFmkBMob/MepZIfmMV
GMwPKIVP0X7NYjZSkGr9hy+NMsE+Q12ODRnsFqB6Jigb4ssCJ9bUk+9JMlcWnjQ3
ifEnxwpoSc3on7vzsm2KkhTAKDTuQQqr9SUpmrUiJdVm4sMWRrCBgdbmuty4VSb1
d1jkH7QZNprbY6xhJpa9l7L+6zcCEQpb8ExQedcTJYSZrXphQ6BsvcbycllaohAJ
wtdLrLaMJ6HzuL5ME2SFOn+iz8PdZZNDUADuUC6Bsa/3Z9/5uauydWo4VHT5V4Pb
PTBzXcWdKfg7b39L5XZba3mkDlK4pFDYDt47ZriozDj8f2EwSRttAIjTGLSCyGpK
EBXvrzU+ks9UbCaZUwdwCMCyR4IpJEQ/lvyN6INyeAyNCm5GcXur9F/XGhrrhXqo
Iu7Eeu4QHhyWQAAc5dCuk7yWG/lAOx7RI7YeU02pPgwPAj8dI3QJJo8N2Dl4zMT7
jEOoGxSXgnFaVmE7N00QUz1XjDK34Jj0+vt0zSnRPJM13HhfSIFHZ+ZAZtAZWSpJ
eujGcAVCy2WiE5aAWT+vnnVsPgwhrugb+LxRAau5hlaDdlNrxOq88HaX7BG2dYzA
U6vS2cit4RdbXJckRz9Gfh+cZry+E1toj7CC2qynQym7sra+gcRQl3FzhFrpobf4
4AUIKTbV9xGp/khaG7k5MLd1V/xsfApo6IzldZu29AashNwgY0F5yQRwhI4b+kpL
RyTvdWWXQXlYFbToPU5/72yl0vuVEWM2uyuo28zgM3sfmQOQdnvy7gSeHQsL+5mh
X3w00CqtPpZhpJpT16/sAAIEwRqOuGgVGi1pv2u7/PIl1KP5GqbN4GN2vcsjVULN
lkIcVfevoSEMh5Y3w7mG3ipPA3LRWpmxn1YjpRMGqhDmQCP+UMg5g9Jk4lbT3I88
Gw5OrJaRAfhJDzW05ExZy63Q0dVEin39P5DTeOBsef6s2vyBjHZA8EWsc5SAQWfc
OZMPOfUZ93YYjFQcQntQOCXmxyzmAQeu45B9LsGtc9fDxuwZxGYbs59HzZW9lVJF
9/UIPJKJeVU3ag1OXJ1czTHh2uM4tKWmwXscFF6xCu22cGF4aF0IUxv8ePpm3Rdv
C0zwkYTvimPItH4LRSNyntN0oZ3xNrgD951XRM859zHcgH8K0CVbdyf9q1ljWYfq
Loj/jiIKpONJR8eoAvSxU7TYICN7nm+Mx1JUABesOm5PRW8OHNdq81rT9UNMyKaU
5tmUdHMkwwJV4/doquEHPsOIXJSIsGw8oWWSeZA/neYzpa+wYpzOcIQ0jTI+o5VO
mOQhy+0kGFdKsLOwGfTB+k/Rro7qsUALbqlD5DUogxLJWzDLkqfZw2ReSY81kqTx
QxrxOQfofKh9BHtEsxR4otzvr0mRiPTnP9qPoJKAG6YUafU0woyausuvgT+zIvX1
NKpNhp6BzvKcEFE549NNwMek3mxC5o+BDoymt+ak6PceishUNtZtfi4zxNA0I5Jz
Dd4kWjVFm0sOtw2bsFmZdNx+3crqi72/WJOW05gp/Ahc1xX/F4xUdjNSsYtYX6EW
ujXRbklZHXqc6gQRhiL+w2veimgE8ErLslbrGDKyfHBof+4h91FNMfKsNxVBY7W1
2vdIS31uMxvtUVYPF4F8lSvIXfH9cR6dxUHdkIsFCUMejIiy/JgxY5O/fz2cGwJJ
cNl/lxTO6YuzV+ZVCvTgyoq+0cf/XEy1cwczeCCiHdkbgpV9iUMvhcwqPnpZzLnh
xT2NgNzWm4Zz+c1MVaRO5Yl7nRHuqBmJC8Rym5/9B+kcAsMIqhmPGJufeqQ9ZvDf
WLJuA9+HCQDrkxfcPlPJML7C8O+ZkmdSOtTG10lgK3R0k3kxOd0gwgXK5ffdd0Ey
/yESpFzzkfJYy6I/nrqrzQ6wmv4GYSwp5Gy3NOqqTOQ2dKEy1rDu8MiTzvmg1rL+
xXnwauphEZMQw7etLhtKOkK/U3VmdwH/aiG/CghvssMZEwv+x4owjaX77CwBMujx
zJ1hUuKUnu7HKfYkxaGqPUhesJ1Np/GGflqgAuMg8WGZUOoiYXljET5YWUglldF5
WoHnUD3VUFhiKapvI6p+HGU4YYXaSOtKY3gAZjNGkHDHVxwVfxotiMFdJr2PEk25
rmiVonw95EG3/ELEWOtcW8tLMqaKXrBHkZyIn7YML/1rm3ANR+26EWv7cCKmlfIK
73CVfAcH0hr6e4M2K9Ahle9OZG6RJLnl+ZuSJou/8vFBSvycOp7i0XSOQkwc0IC0
Ao1Sx8ho/JThHzmlRfazRYMkO9lcwDc9iTBNNFf2pqA3T0oob3m48bnZLNl243fs
VfUG+hfuGEPrJqxoyWLYwlL6GEjnyZ0WU8hOpKU9M0XrpTBAO7zr1ucwjvTXDx7a
aEM3KIsIkCh/+xRtwI9Qnydwta91/aJs19DdNZU2cJoMtWAaHw539JDDKfbnyztH
LPqDuHiQTEWg+f6eKDjSp5srccDzIO5yY3xxWq7QVs1s/ly318Ifx7bcboGPj9P6
nPdPIX6N7ZULVk9u5drH9ZFcN9jk742xMdiPRdrtt/+zrO9Vg7PVnvL+iZVH1brd
L7roNI0X0VYvThT2DMHipVNxKRiDpVfKvoULB1j/3q9YmDPBAyYRkip5x+8R+xEb
CnxF8xa5VDs18a8xnQule2t/bMHHp/uzwpDCZEs8mjKacKRdRCaA8urDPJazektb
Bqyz2DnE96HKMDscyBPrIulWbUX43vTpiw47jD/hmICmN1bHwr3CQXUm53UuqVAE
OT6FBQmvc+e/9iRCIcE7JH5CtzE0EjF9bnRNptSk8sL/4sDl7z5z2pFVYl711YRy
kovAPxHzNCuuZOWuX6TMB98kC2/MywIGh8f6B1vqxd0ZHOuoYsF3utfVOtBo3FW6
IiNyH7BKY7aVz5AV6LqlqQ==
`protect END_PROTECTED
