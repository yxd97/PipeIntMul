`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U9zGvo5kJ02v/B9jJdApH9JbNA/vbbX3uN9HxNIJaqQFYgpAPnQ2TuIKBzlXCxPd
mQfpA8AeRgRzbB4l7EQBAq8FwJ/I0KgUH9ZE+LbP+b8wSh7kyPrUzu2/OP4VaIAI
GHXkFK305lmC5tNAHX9jZflX6Ghq/uvejotYvNYnMKyjLGSgxgHFj9TRDeFMrQWO
oYU32XA/Kz8iCgI0RyH8dtoA95qwK8S8fNxG1fecCWYHZp4flrAXH8UgQf1OpzA/
pizYvYsclceCDrGXIJcCrTn3/KimN4v1iI5jykHyZLAX0aBmTm0RI2avLNXstEX2
LUk3vAZfXqhtMb7qw9GiA1ZLjYlN14J7lmgHuBJe/ATJzP+dLINYywPxm3L9EAkT
mSmTFcLReBAe9ljj1p+h+JdSIgeSlMvDwk4vcY4YDqHtH/CK3nVvObBTUcndDyCa
xyexwARDhuWIeSqKKAHrlK0YENRCQSVN7Pke2U7lnAGqVIIWpf5ihipfOIa0+mIg
VHRRtxhY2itctJPd16tT+TvqGBA/2XYkpZXtphVmtsZQI/QIpgRTZZ3iB9Y3KmUL
5CmFlsFSW4B8ikV/61j9Sv92ji+fiUADenWt2m+S74ZJbqlxBJnOEv04ktOj/xPa
9+0xjRc71bv9XDXuQwDyBog7TLOkMRnoLZbUgrQOUoY+/8J9YSWMv2pnCEY/Bzxt
OFF4lo9ua1uykxFGD5+Qs/0ra81/IGDnO6TxY3lglPI=
`protect END_PROTECTED
