`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ONk5J24Jb6TVbgS/EPJbC37+sD8WL8xwd8S6SfWxorZYvuLFV5v9xo9Oooql14El
Y3QoqSFcmBNafNOpyhqAraF3K+H8CSK9Ag1sKuLB5imEijONX87tUndxEk9DXVtL
Z9PtDU7kvz4VxGxOQFktPLyfgGislzZGijhUzm4jT2ZZn0JSghaICxDjUUFORXTB
tdcDjEDkbFVFIKsqW/PeNy55twNFdvURqJAjD+1EjLli6KKZVwPc1HMsa5S5PBqr
6soUuiA6EtEFR336WtbZn+HkLFRuijL2wybKMg4JUj9YgIOfn5GZ3I5rsH5fQmSh
GbMSYk2UblbqjpdVKsw1QqydO5589vSO4aIPWhkjno7xG+BkA4e1rQqwEDaMJvwL
fVSmGXJHdEVY2KyP67HU6/EDMyN2w1CPU3pZxab/Qc11YJfE5afjdwCzam+w7LBr
zV0wrfclI8z7/Jz3ha84UD8/oyEzY6fmAjJ8Q64/Qkb8Xmg5WTMTMLF0HxhxmVaa
/y0eX67NmzKSnK1/haUEvXWHJ/Qs11P/JD3AM9CPBJ2xGEstsXENiQVEfcf/T7aY
lR2EyusKWt5K0iNb0BXdUjBUmpOrtawT6L7nRbmKmc75uLtyF3ITiDwnaIQPwhbf
qAsRHfhnFi29pTQfMJdxRgaYM4U1OJeBxJn0Oo+ljl5FgP+we1NZBNrFsIBK+54p
G9qV6kQKbgEkATZsrOwSqUaF3P/9G5HDs/swuUsPNfDMKt3oQU2tcXU/r+wKtAs7
eBhGNtf9tvZUEefV5Ic8B48A8YHDOoSQK8Wvpe2u7Ye+HjQvtAqbE2jHgLcqLhKr
xcbWFnHpMA3nkZh/vRckgoHvkHTJ8Ac7tfHVivLaRoXd3GbedYsIdQExp1aytPnQ
EDN8wtvWZXmJCM33F3YOXqhbXhzYqmceg8YI4Jb2BJL47r7kDLZoiJu9njt87PfA
RVGfISOrCg1If8ClcCJISzx8vYPdVe2cCPYUxumkbgSm9b5VkkuPrdhypvijMCR9
T9FZcbtRZ6X5liun9UYXAUiFh43QPW1NaMK9KnBPtH+x36AW8GUmhYOksZoTlWyU
FSUA+0BQGk/FxOVsKv4yG1SzNYDxd2Q7bpkjgO8TkIJxSy/LpvNJExsRXSm5fa1s
Q9a72LB+9OkrqnmhqbRKmnvM9zh6MCdkW7YcmdEFd8ZBLCR+csX7bl2E2tvAWEnv
5qpOEC9HpNvmLiyQ4oWeHZJlUwnGW1VzNmDXeTaDcofMsitGanzvH2LBZdLUQNIO
aKR7JtuED4YAaAu3q/YrqQ4D0OSk84A51Mn954y6Fl4yTSSLheERQGDpImiKBhMq
JAzjaXSPkTACYEIbjhLjYpHA6UKBZWloLUiVeyCY/4+UJxo+taqf5VprxjNnqGtU
Y/jCWzTZEH7NlK5541Ss88W8dqsJ39d+cZp9x+r5Beo/zaNMudlpSJ1mI7P5ugCg
oGbJ6e7P5ZmGFeaLHJIywSiznMuIvTyp5MibjUfhLLrKUe8Ygv1pOYER8yWcgQBV
2NW/37MUy3PdkiCImB1Bahdj5d+v7IU8Bx2qm4Q6dn/aUUI1NFYpji8wj4ygW0f5
m5PSenEsIiVvIHj2ur9b2V6hYOwDTDjyg+ujDl66S4W2B+xw2M+O4W3qRChwhVFO
Lzjj3BtJBzcF7dc3u4PTCC+VBQe4NUmhjiNOfh22FwtTkC89tui7WPZU/SQZgiY8
+Qfl9PdeE+I1c5kF7au+Y30ITdL/Iqcnkr0ntnktdt+aesAh/1mR1eBpz+y64oHW
t1H176nu2ePwXQRcxgFSjF4xQQ4lkRVZ+1DxwUs9wlLG//6ZOgUCuxeo1pzk5lZZ
Tjp+/QoUnQNxE6tud3EyhcygjaxvpU9IRavZAI5rediYFvOGX62Ad+E691yCvPjz
VPbGtN1y3QwtLJcJvHjZaZBj+H2NwZH77OpgINxkmmcHOrT1aNX29OFrPlKiE4Di
S1EISpmpWAvZDkx+8zazdSEv7TKbhgfeERwmIZavnFtLf/PsvIrDnn9f2G+eKSRk
zQ/xG/vawM1Ei0Cl59ObUet+Lqm12orLApGnlYGZeN/Qm7G+5hnefq/XcHb7120B
Aw6P7QNb+c8HOqoRXGYNwjt11EoudD/2MpvhLJtAyNmVqun63qLhoi40jBbk1vmi
TtOqN9rjUd1J+TNwT6ZEkF4VKGNp0a1jxZ4Se48R+P0kc4D68auwl2WIc+I4yJ2P
9J8sKpd4fs5vZ79cNMUfkNvmoLA5KtyrdruIhUHFTrv4RFV3YpLRBnv/nLoMCQZn
3Ddo4nbzOIAzZIs3KMnK7vEVptWS741tPyhnlWLa8mi5V7oYnE9/bJe7+uBnuASd
ASOKWFqn77n/yGOsBH/VoWmWKvaGrwRLCQMDdEEDGt/GyB4h3XbstZds9y2idGsw
OqurFt5TIl9msAzFH+b4hViYLJ96DRcqiVH9ucxQhSf7Dtx8QHxNnb25FY9TKJ6X
18E6Qphoi8CQRe4I9JPGJVPPcI6OQ1Kv8Vw38SU0Z2ZCnIL5GQrC7kB500L+Kv86
knKJlY1GHIwMP8xfGlADO2DXbK1vcczNYZ6ds2DY0PdXesdLth1d4EQlrb07rxlo
4x54eLEEEzujNeFVV4zl+GG1ae9NP+4tv3sPeElUk1XxQm8UcYtUElDJawIWWLWB
A02VAf6I88NlTbg2XVJv0zyAjsErCqFHwwZf+QyAww3wlpTRsmZ2ubeid7RQDpwc
pXQF7vviq3wac1NAQU5yYCudTD8w092bvZwyAH70a4zNaq1WQnYCOXzHtTuQww9C
uOivGls21iBkl12uyEILGu+G7KhLnjptDSG8XVGIYUUooM+aft7utTVCbLCSvxW2
ESuhvO4yE/VcFJbEwEqfnkyQI3agRMLGBhn1RzBGM2m9ea8LbFLO+AKdc5c3TmMA
CCbA0yTo1BgDz1Wlt2LgYiUJK/O6TFM4gRewTAKPQjo/lsFkPvAZzZ6wb9c+0aqr
grTecXGybr8j5RnU/mgl+Rruel7u4a3aWy2LE1u9KV4T0vHnvdpVpKOsEfQFkdXJ
Vt31pUSpaQEUd2hGw6tHre0IKFBeN6C8BIBfQ8+4KscLrlYDdo1qdtVbzQX5Zzm8
RXSgLRD+VuI8Jw5wjyzkjCI4/MD+tFt/j6ZoJvpwYHlntzZKniYXhyhZ+EmOElmb
+mAOivf8JmM+sj0ifAgzGrd6MI02OVdNi41jWALby8WYq7qGAWE59QbtcMBRlTzs
mFhWsUOGGfdlfy0n6nNu05EN7/SWk+/LBmmyPNm+VAsIHbpTAP2nT2kUxew35jD+
fDU+LTRtcl3FEddhTa6drcxEWR6WWgFy++BbXgdQyxAVg/y9xpGN9+5XEAejaw7+
0mnrAq1XeP3mmMjbLIrMkbXudqqHZbByYyXkStLvjbJcVfzZ+BRl+5HIwg+IhtpB
2/xWcPt+LkVNDmTuSd2L7TleHHWbuEty3FrJl6wqsE0xc831IIfayLYpULEhsvFH
tzzJe23+nlqyBXteeTASOUvsm3jbXO+YKezGPklzVppRhsWohnQXO/1k+oQDSn5V
2IpTCZgpTswRRm2nlJzjW962/OtK0Gr8cJ49liaoyIhT7hZpvC8UZ2KRbYQS4Wji
NoH0cIYPE+n0tJ9FhKw1clpumuB6YswRQg8GgfXJ4XaQVq3GNxQUbbCjbKo9aNA+
/BjyJlgVCY9AR1CZ5FwVEaMX1lL3Wnm3tEBJlirsG69ZnhQwBgZ2PV30S8wV6PUw
LEhW0jqayLnYbqrW6lY0PuPChIpEBTD5oj9Ibv3aZQ2NX7RXhZf65WGOgFztLsvR
oGkwwXskMcEa6R+hoscQKHye5MdFbXl1pJe5GzQcNBBoQ3WPP6csnaHYKuxHtIuy
cv4LYKpjLCqlCzWIyEPs0pb9CHTy9wW0qzHqpPPCxwjb6kBClPzIHxJk26Edo5pl
KjTjG8eWEHiXLlIjrsLzbajwkN8zWE+GCFg3j/xvk1Gd6DApHzvmeS/ChbLn8hrY
sVGJalNtuZjzs+8sHBgZTiL9e27tnxs+yHun0TgYORPLbTtPagezpMRALpK+P2XG
WbaAzP61oPRv76dUCEmtdRfX+u9IcKw3kuFQNHagUpSVea1t8qxN6E3CgfXQes/l
UEr96gLk0hS8q9dfiJBHsRVQlzMiBBCaxA38KUTkuDC1MhF1C7RoZ16AsTf198/J
qduqrYZhwRvAdj7DfpND0DzErSrQCSmJm7YtCIi9E3oDS+71jJUOgbVMP/yN6j1r
3edrVF0zlBzsqTneE8rKyEFPxrIzsjN99sTlBJTetxxDH0xS/6FTsgjNgxHm6BHx
BLx4gFRhGAq5rafYLLOoDW8xjCGIeOtBYrTL2nq8B9KdHVCo0wWhBH71rOaKCl3L
jc/7SfrgkrPgcyYASTjtAbo4rw26O77xkCFXcD/l1e6BupRTvYOTirkFdGqVxIrw
YvXLzRaJbuu3ZYdhHQrTG3R5Yg0ASA4RFTTgi6hnhCVPvROB5p47FBdok6nYMmXB
tJTsuxwLYX9Q/KLz8lT653jlmIdYOudbRg2NvW/EUM4GXiRHWJaJQZetqStWxAHc
3f08L1697tKKqwwNSG/O56j5m/DGWga11uUx7jdelAHBELoKFI/u8cxgbek9Ctwm
1+HMa8CHuPgHB10A1DBYjGv3TpdRmbVfVBdjwvN8ltNEard6I6TWVZHU5JAfQChs
QqXzQvHDtZrH3WBd3+tMckuSX7aaujXb1+IefX5xf1LYrC4j/RLh7I8rl/sNSLsC
Km5bvFdI9t7TncNyczr+arQhpEfa7XuttuorZOA8ulQ+ftGJx6vIHTSw6Z0RBh/D
K0Is8pRxzqr7JtB1fVzHsOCrYfI/jEqBIR3KXYcvNnZTKEa8mgNhwi9Ov0bra5v+
DlYwZw8HRjTumXmM8kfk4CxttylH2uMR0Zdl5u7QYOLS0KooBWX5GVC5SxNJJui8
7ZdZMUCVlg4qF7Gn+Ea9SaaQL4rVWDKZafk/WEcWHlLgIoEdGlGmmYw6WwjuPXQL
HA1L1pxz7FMa/bSiERjmRHeSgA6YH6noBNTPCfyF7mrXUA0oEvlgLv2i8VpSuezU
E5MhkxH3+pSTDhPlEHEj2FFzFC2AH0B+PMo7cWD5LnidzWvM/DnYOPxRK71vs6kw
1oKDgQ9kBeDALjIKTiBME8t9W7kpQnbUyUFbnebQKrU28pHlrhXDXT9mvpdv3oDA
VnmmnaZQC4TC8BWt+D39UFrMBKM5qiPAj3kCBuYrASiV712tXbjr09mWqxPIAvS5
E5gpaBxRuV0nb85W4dO+vvnrC0yFq+aoS5TD7ww+RKPFD5XdxrsX3ouloKGUDkJV
NBFj7PLi1vxgfTM/OIJuZFxO5M4wFrgfI2idIe31n8yHDIqQFiJXTfiJcYKInlbB
FapfwnkNoATbutYqCazR2WLX6E6ZbwCcX5oyG/3PyIsE/y65VKRT1ATpQ4ImDkAr
GhNklMYfY1hl4k9CJmaQVTyis6c3kXGkhZQxU1O7ZQwmTQ7o1orQBhBxsXbuRekn
mb6jvS3phEr8v9Pxrmvdj2fLaZSWO5hUd4aUDGsyMcxDO9jC9VfS/hZJ3MJ2uZ4/
2SPMJOwgDzgoxS29ZRX3WhiImAEFS9IpJjsDxqgdhtYuFgQTxTgItxtmAGtTn4yb
DQdUmviPT1q1wbr4LJuZVP3nSTNqhUwpRDNYfv2vAAS4eS3CHGJewbkxlEVRibG1
Ylpvf1ZmVNEqu6b0Tjebx1F3vQfcaAyE1FySYFvIgRvAhRbb9lTP9TaIWsWhtZjw
Imm9wxxmvaYxrW0pb0ouTasVvy/q6JiUgR2rfpHNjrpSZ/+EH8F10Zi7xkbwPb33
xfaO0f7rUn4/OBZsv94EPE86fzRrQWeW/o1WZsLC9rv+xbmOMZb0de0/cVn6LFH2
KCz0mvTOGXUC8DcQrjXoDxY8PH0dxdLIIIcLiyPNBqWOsDyMfOz+cTA9RGIDw5oL
`protect END_PROTECTED
