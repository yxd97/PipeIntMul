`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T4U9aARPW57nVfl1KYGqiARjkvXyrwv/sbscLAFM7GfrofKe5SJ1Kq3tDjr+sEJG
rXTM+uU6Y9x75o6axREXdiMO6aHPiDT1PAKzIn+CcJdSlrHQ/iNPZk2yhfdfudCp
RpHHrXm/mwv11LfmE+Z8DDI2q/IHSr1vd7gYxp3uZU7leI4fGhrWb0qXC0RZU++i
c972vPP8V50HceITWmeU3NJgPx2K0VMPxbDwfsm7UIExH2/h4PI73selzgyd2wWH
6iR8R9N0v8r0PfvGliFBYtjDUK2LkJ4ysbORTZhcUMo60Eh+I0//mBhs0pR7yDcc
AOSCO33K06/TarTf+4w3nNgUEUwe0GD5b7GrmzzS8UtlsKq72IHmPdwu6X4AA0D6
UHuYKRx4rsbL2VjoMse6tpC1pz+Rgk1IKpUVOVaREZZYHeaQC7BUgdliNSIfUAjE
bmxfKmzvDL5zeeG9LdJfRBPk6RfF0EBxLKZNdTyHPLXDmI5Bh4H7LQwTRVYTNiqT
LJsUv4zDqCc4lETGC0M4/BLKdk8NLPEv8r7MfXEpLUKe28WGowRrYlGvxt53RLj1
5WV2Wx14DQ3s0qo83BRkqW4yKvHIXpBsKNnQ8ZB8HfX283Qj+J99p9T3VSiucNfs
hqiuDFqn4wFYpXz1pHACBFxwVaNiISy+AJdiDNsh+emuaxXoymwj9Z5uEU8l6nb6
oj86IK0EvK4oixY0KxMJwxn7s2nKc0ab7e739GI4ovg7CcIl1r9tcEI8UTn02m4T
RkQ29oJJuNZTG7bEST6Gqg==
`protect END_PROTECTED
