`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HpJKFVcbL0JOuy2JjqgqtE+uFBJOhF1p58B+kEDnL0IzIJQDIb2S20FEYGmzZwuY
0DGoihqLeL37enBIwBpY79T/7DtDU64nphz+qee/WQVSgvdSZUCCg3m9xC9iduNi
l1+5gx9My2RJ5KpOuQm7Tp7zTqOxGBeZIDdtrB6bYeaJ5dGvulP+D5jRM44al6nG
O60XO1Fe1JkD2v2ig08aah+IagzT8W+9yOxrYa6FsyU5pnz4gHTPdf3LaBp5GiLR
N5RfVnY5wUkwrD2YMOI7XRi51xKLfBBQRN/aCd1+2v8Rmjp4ere5sP2ItnDhK5Z9
5V5AbaVI7AvuFabKhq2YMQAXkDD/8hI7TAsPk1XJImYOdRhWsbB8AtJdfI/wrl/h
MfXypcLuX+ahsJmqPYi3tRKtR6NtfQgFVdS6fpQEWlTxPFj8MrqksGglUP6ZwSYm
`protect END_PROTECTED
