`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9yrgsQH8IYKckxuRc1NL4vIz4qgXoZDposdMa8vaQghmfbPjMksI8I1BFZYbutcq
fIFIyGussccpGTedRw3vn2OBl39rQInFsoI0dJHjNCiqki6m/Tw5fKivNkMIkqRy
iUpoXJkqCYfzymQ0kaJiNrdCfpenTQvId9gHeNAUMsRGEjnhQ9sGrezx9uHj4rck
wWVq7fSEnK3reHwpAwCl26Fzq+dSKsXbSfz8SLc+hXPrpblGzBYBLxXhYLF13il/
kTCfj30g6ncBgvFRErDQ4HTiRINZ4Xl/DLGJb5GlDhB2iqa2EaT4tDs72nwOyvsO
HGGQGayyoCUS5HJVKNJj6DpBtPJ437Mj8DITnUGqyvOcH2TqMAyVjB95h5MJdf8u
Y8qUvcWywQtrIlxM1PqQ7vz9SsNLYVuvlqROXYdO3WNYz9cn+THnLZ9VLX+pm6t5
ib7D7yAw04XZml/OsuE3o7276knna6rOznQ8v/bQ7UTRfD51tp30No6rqNgHVWJo
d5Hji1PMlPKiWWi5I9hSfWHG8wJLosxNaKddZipCutEeVQ1JeT9cEDHQViLC9dnM
LyKEvih8axiVn3CBo6Jrx7AkblWzefIDxhX/yCcb+fer0xg/4OQgUgW117EDbaJA
tqGlIsVHSCm2+htaZe6GT2fCKCS8x29OeMioocU+P9Az5mH0c0VybHhG/aYY1FkM
XQrP2nW0cOHOmKSTiNUUswz/hKQYRavVul9I9pSDhVbEfNHvMdME2DJzJntGTkre
90u+lwslzUFp14uihQxxTUJe955QEJ0Z5oZAaSUXGSaZVE1yZmlHKgm39qCApGTr
uQxmo1q+KTmvGCOgamFAMWlnByGjVphym2JhD1AtPp2gOU4tJCvgPENo3PAZgkZq
IqGRXGmY0nC3VmHK4mKx2Q==
`protect END_PROTECTED
