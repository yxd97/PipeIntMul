`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b0lwZIoCBw2Sq0os5v6a4Gs+8UQYuUj07g+bTQsEOAvN5gR3AbfubcXgUrNJx5Q5
pbJWuy28tLyIL8Jf5Mb/rDvEtZebAj1MXCw/ZR5s2AD4aCeqBNHmqr0gdAGG0bvB
PbIcd0epmrRkBUikHjHcjC7MvgEcpVxW5Fp7It6z9F9A/OM9tkJ0Few+Fc+/C50T
Vu815D+Zukx5/tVY9vtLPRXl9Oeo5p6IiLcT+orGpxQKFRGUoV7ESIpFfVFJ/CYA
yWOKmUSJZSKslDu70v0mStXIDJBmVECSyLCENZsP4nSUiVn44krV9OyFbDNC13hK
3YaoVLoFZS4a/RaSR+w3ib0wHtLiaWLtF+AW2nQafEkSxNeQtVuA6s1QJ1dwkX3l
51sbR6MpyjYhWr440x8l1OIOUuEDzLdTGo7mO5BgmdZ6JPf7kFtsw8aKv3dcXy6p
g9e/I3zXLju3pjVGpGv55dJFdQ4CoVkpakTwW8TnGkXdk/u8kP9Ht+RicRyCESzA
vpXCLy9rNvDGyjSU502HAHer6+u1tXOYzUIqGJLmg+xbuhsqRZFw7xfdUmdRbQ5a
bwR5cNyigLta7IhdYTtp7fN16nXzRDtabGMbVipB0Yt2gl8KfTSc3i8+u6srS+3S
lEfptQCXGXyrbLFB3o+blw==
`protect END_PROTECTED
