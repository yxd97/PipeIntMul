`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V3S7VHipd3/aEV7U80xUuK4VYXpLOxDYtt31+zSzNn6qfOTuc4Iw+8sWjcvA+j2v
vObeMV5gDWaxloH2juO1syycDRthqJARMjv0wxoa86N5ku6r9TPO+6jDZI6AF3Ib
qnbwXqmAwC+OGi8FLS+64hVJIh7yMdWTrDoDnbfBKEJHSOhLXG0SE5HgIKjvgQER
8eL2SJjZl5tKOgBWFwCejg1tESK0sQeyIBHuFxpZ1x3LLqJfrw2YSeL21rVKbR67
kaE4/9QKGY7RwOx5dm4eGVEK+9l//ccLiF22sNb4M6vNMm2WvrsUgXyXgtJK9qgx
ggzbyselh90NfTp1s0dv+3AIY0DuTLg69xnCwX1CL9o3NWM3kI0xKVIbKdV9/hFX
5wVcVqFshIo1qUUWMyZBWkQQa7mtCVm/o6H4dVc9nyPveNNbjFGx5Wt46Emuu4p6
YGh9glxGR/a4pORhD8UZVUKAtUwWoSC68jIEQUzLW94v0H4w8fzn5JOJIdg96O3q
KS4ipb3/1MIv3T6/KR0XGe1qx3rIBK4c7s3B5/PIKTKlii+0IOc1kZ/QrMWE7A0u
WY7DoJDv6I8lnkgliYi9pR4HR6xmVfno5vR4HL1HGI6IN0YJsM9ZmWq/idrVR8St
GZmwsJdQqymwoy2NhxqkpwU663wTC4uSWUO0gj4K8DO74Tqbmv2PDoQEvGgOC8OE
7uVTBdpMYdj9NJJKK/FeCjlXIIY5l2J/40hZIsyb8o5f/aLa2YvPkly77duaP9Ri
TdIg0hZZU9FM2KSyRtgIuQ==
`protect END_PROTECTED
