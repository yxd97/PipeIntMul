`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lY3ENWJaEVksUyj7EYg3Wia+IAuIUwolPOIOR35GNlq3gDYJu/w/UVwzEvzKz9qO
qwYHwhBTkAteGugXwTM8kF3weWy9XCTnSiPpu7XU2KNsaBBSopKa8QyEpzyFoFug
5g9nCej369eAqh/xCCZXLQdRJGyrEObGfq59fVBvLj5HivfvcnbhqzcA2fE/zQc7
sZNZV1QycUGF3Mpodjx9vRSocbkbn490+PIQhnlJDhba09HTPE+d2NvmaFh9x2Iu
8cu3EbLxEbattApsMT6Cm9/4c6AtP6iYkDadxOge4Tv/sNPh9zydU1h7qIEfw2PJ
QXxISi3zetOedkiwBfsXQHSEXpEn+rBQpSXvdWAUzfcTjp7zj68KkrLcePkg9NKz
`protect END_PROTECTED
