`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gk0/ZGQ93jq959WWei2hUGYm37nnNzBCLWMQwf+lWDmeCTq2taylfy3PyQXiByA/
Lnc/1WvB9eKrnjeQEUyZi8Cm1bYQi/H7WWU+LKRBPPBiNNMPUBu02smB8pXFDwuW
JJnMIJJ3+lrIyYQahFt3LHPb7dYEXi62bn0Ax5KFZcm1qwyRRnFq/5igjGO83jbr
Qos5/2pA1srpUihIx/X6mM22V3zlhVnpsZUZU97sVO225hrmA33SIXes8uTZMSH/
E2Fzp5kJCFsizgiPf9RakyVthJ2OUb1xYGBoWQ22S0Udk+44rZjwAp9Brx1sa3i4
IvAWMD/1XzAF4S/AJAWdQKKGA+nNdJQqcS9Y3SM7EpJA+4hZIrPK+jpZNLzTCB2D
Dvn+XMQIb/g4QhNbXVPN37IUjQWTXZoD7T7TWMGAP/BS0R3yMB/uMv7uqG33MAhB
d57x7NoO9Q6eSvc5Kny7O16BSX8Wck4Sb45NdS59yNB43gVtGSGRmH018+6qxmRq
5MuWSIWa+lDNklM8BHD0pwuiUNWx9cvk2mzE0VJvqZ0NX57AfIIDuRT/WE56EcCt
guiAmc15AqDK3Mv6bemtahkE5Cl9R3qhMoBJKi0zGT/mj9ZWjob9Xux/JFaotjIF
/x+HvT4Z+0YknuPYFpuX45FciaSkH/xy7lehO5pExUja1YfPbwdEh09iZTuEARWV
Jh6sOyJZsTVlH0vnwU75XQbV4HgeaaqLh9mD6F4TlFEgDB0uyUuxaUfgnOPh1C7N
ls2VxP2fuSDmyEcVwa8LrcmiX+m++dQTzRDtG7fRK0nZ7+Oerdl7lE0bEaQfD3LS
GlgJAvQddOugP+O1NzoSGUQb/Deb0fokWewfmW+ktfnRULJyocRu2qIchZYxIUEp
Jse4hLe2Vq7aGE0CYv+ElxqCDcqelMgftigHoBjTLaLBlNvqgP2K2fI1fZHoKYRf
8PZDeOz/RcZ0cdkPlpDE840C/y4XGrRjrULiqYWKsfQVkmuWTV4W9ldaTJeMUKI7
Z6Y5+i9l/BhUB52tFD6AsiTIqwN68DMscTC8AgJICtRgXLZntzLf+E2oI8spWM4P
twgeGsIGzrNsPNACB/98oKFaVbFIjB9VHXMSHonuimPG+bD35XdgXjzRVjCV5uSB
vYCTwXPSBvud8G0wTp6RkYLBSweFWeX3pGZ7fBAyiMfZTHg/YoClV0c+J/JhsUmX
scrLU2JE7GwhkvAc++vTgQ==
`protect END_PROTECTED
