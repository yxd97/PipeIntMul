`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BiKvw1WT6RLuMHWLMryi1T0qSpXc9HgA8KIss6sJzC2U9qM17EK9SevMId76zqGk
vFjz3535wB6dCU5JZ2C4VXX5aLvFm1dv0iK0pknj4xpOaipyI3eaLsN+ttPPJjDA
nM/Zg9IAulBFliUFXmCfC7jGILR5ciR55XmIvb4uZ3fhh99C5jVpUoLdgM5BGV3W
DdKf+TuaavDhvz/Jw3gbLTniZpkqoBpFl2JUbF+Onqt2qNxIXap2HYfMEKdp1ew/
6snBuXsom4+BMda/eQArhQ==
`protect END_PROTECTED
