`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MKa1rlZSaHxNLf2vjUl56NfDQPizCH2N1e/8OxS6ydSegdDudAKCqEPYz1S8KT6L
ARNsfS4gTEFwO2K3uRb3v4D0q1tBL+0t1U9LjnBoCdI/fXkGLU6PpEbSLcu61JRo
7i4ow+fZ4nfHJyGDa20jN6pOoUzNd8hxxllUk4U8MHvj7gGxUaWtevK06xbDV/Na
EcRX4puUwgv+GYkSg5lA2rDvYF7GMLvbh2qoM5VXp5oCDrTR8ilVte1Yix0O+ixs
qOfZBFKxATCaTJOKLVoBCJgFuryNLFfSdigZUkBQQLBKSn43GIo2deKkdYaCNuIa
Wh5dTHZcDjbQlR8WpuQ9kyMOb9Q1C7csGFQ3EY5ORNMRaB/S5z92NBXtIT0/l/8K
/6pAv4V1k+rmSD0gD+TKBHx8kPHr6OPhGT+frYFf/MV/ZwKMmFd784cj8mnbk/Ks
8dEPYPwfWflYYT5fwQcIQbAiESKsS/TLSeR17/yUbZtC6whD6ASKjk5OoodrRbBm
V6U/leLdJh5EgQMgPySEJxOIJ5ZNUVq5MX6uykAVIOLmfklchZWMs2AAe96IXne9
8LN+xDMUlfyCSgvLwavsiQTD1wu7umOO0P4EUrLDjA4=
`protect END_PROTECTED
