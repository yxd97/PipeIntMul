`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z9K0eMygfueYE5/Z7mDXc9wwcIGrl3abW0c1eD68CO5ZFN3RaOFoGXmFEQVtua0b
vlycQEr0TPdKN8mOkPGCXS8vHkJzw0s31Lk6GrQ8p5pkieykjYhwHB0dj9rrMjJV
8SdcJjonjUvvTyGLz8kUDnBKZB/8qoIhWpVh5+waXmMqdCgxfngPX2ZmHmtHM4rh
63GdeRTHA82j2r5G2AGBZLP2ASY2I5Pg9umqEx0e39McVA7fD5k8SQRSM7vPk/s9
biXosuMeIF5sRqqV0eE7piE7t3VlWqzAO6uA0ZY9g7J16Wr1Nu1WhSLaRkEwODYP
IdmTn7/mE2i1tzLBQMD4V98/SrxyWnCXic/hBXHniPCftnWCXccfBj2ovlkdfUcX
dTR829ndOMTWEC1tnD3eXKX0MrwmWM6h4wmjn5Rsxuplgz8H/EnhEOdGYlOsfSyv
NurA65bh5yNt1VUBdMpMRVJ5dBVWQ1bU+DEmGZ70hpLfP1qIcTiGqMElG23QhHPD
M2yOW30J2iVL12zsZOd/C5YybnvHfIAdrs3HDZNdT6G4ovBAEwxnqdKVy0gGSjIu
VvlXNkXiiA/SyCJCYuU+bkEgwqDbfyOBP9Slg3q1QIpX9ToMnfQ/MPkJnL7O/AnI
C0/+/SK56EuIWdOhnakDr8H5taijVvgCYF0Lc2maixhHWwk4eZRxlw+7vhAu7SHH
sA8BmfHnh8gFs60Qf1xIFyAlIE820ZsmQ2yPE/eGwBWR1r+0W+hQmuRUCC/XOmZL
ALKoruTOCUHkNuv/Mfv6pThr7d63iw19D9ssp58PC+JziXOxVOUMne2soxHBQlY5
c2wX+jVADHqk1Ghaeru6OUZsR8m6EK+ljwCDgDJ7ruekAcompadYfIhHyjT62tWe
2Barg08dR/crfCfOelus3yBFGO++0NJfunwUMPo8g3B+uiwCE5soGuMlcpd8SMx4
AkzqlT4gzFWe4i2nksxe9PV2HeKbS3Fkl91JuCkqWXjP6JEqxpaFL1O1HULS6Bmy
TlW2U+6Gf3r+MpWCwBnCJpB5tJQgqCnNOiQ6cTRmXI3jHhKcEeMISRZeU9Dw6m9q
IJd8kmpQs9ZrifBD28UER/oba18vjAo9uhxaHTF0NiUNBzlXHCcQUTZ/bI+dJi+K
Dj2rIXu//eIL3cn8OKj8+Vj2Kjoj954yzO4jhERvH/HI5V+emNuGzStKYq+7sp2n
Hyqgy3+2hmeCIM+TyJVzh3v40Iv41x6B9Fhid36jm31ZExEhvYLKhIicqlnpf2vU
ef3l9NRKTMPazh7Z5ZrMvz/DqiuRa9x5k4RUC1RwMQUjeWpOFboK00IfuClGSUcC
pds9vX1LcRBcvYPjk2U+ioQJ1nzIHPw9dJ9Q1GdIUI+ajuQSRwuh6Wl4A7ZLwdba
WZq68QRQx27oCUkcVJlxx9eMSiRF1QPCvmp7IxJVHU5k3rTFNweYeh1tll+fVYwe
RRPGQ82dw3zlgaRiQjuUzRWE8oFV4n1RWy9oNq9giLxYg2h7piqbBo+Amd3RyBCb
VtbEj4aUbH0PnJrpNPwh03xGmVG+a167jAizImWZBL7YJSYLeKEX4hZNvxRZMM8q
r/Pca15W5PKIbJ86s0PbL7xZtJj9R+g31s6A3v0RlXnCDz54Gx5br3amuiL7SQpE
kaIHXjtHlWDFgskdZ9txK1IeVr4hcn9/8XMq1B4FcSgoBEnw36hCiOIhuXxcmYB4
UJsUoPFdazZBEBZmSX6mkkBavEzVf0m3FO58cIKJhsh+3Hy5yVy8bGZqV35ZE0Nt
j8IAE6b4vaoYE+Gz0zTkSxOC7iannBpSt4HeAx0jaY8wanJR8WTddUk4SgrC0MAR
t1NMQMAGFwk058osnBqZVhsAIhXHJ56JRqOhNO5UINmBKkBICnMBM1Gn8M2fq7K4
s9egeYXH9LbXegqrhMdWPhBD8nqVeT45AFk7k8Bu0Fc2Az+1dYTwotY30ldhSnaK
z2xLqaE8V0ur3jMUnT66Pp0X/CxcoRdc6F9wNoCNm0NViscTtMVsc0NN+furToOR
FswuKjMVDZV6D+aLOJf1Yg3WVpb6vLuyL+YUsq0lFcQMGgN4W6X8LwV1Q4Vjlp4D
wHavxdWBjBhMezoulz1fMQ+sFL0vi7OEQWQ/W7FQlopTuOQOes6o0IkC31/hGI7f
P/YRcWwZ9uZ3jM2dzjwNahf6A8SZGW74ye74Ym8qwTrokCk8JMbjM7kkKQ0z/P1Z
NG2bFEtW/XPqCbcenz3C6sVco6nIFmVn7vzA98JqGR1+UKaIdXk3OIoxpG9Oflpi
eQ6nJ1NOpa+pKIlMmDdd5/SKNTwdx4viTUvK82TCgfVuAiKj7457lsA7xnzMg51l
HHWKp2Fy6behcrpLrJsSa/Q803rfZ8fmZcBucg3nh9WNdXUGZThlsJ87isk9zFcJ
+1IzgXm8+ZYqMUaM07tn467IWFx9SPBvMcrfcMBt6WyqJQ3ISgkE1wa6baABter+
/c9XgwieQQflOEmEOXC0vFSX1DEuG18pqxS4d7OfszVkvJxK3TaLpGwdrJ1n6B9u
fMDeN0i7Ku9mFTSDqO2VKdEW3twArC4ub2fy+3+aUh65TKOgpWGPrIhjD+RyCZwi
CuHF8qZE5sTXfJPGah/Ey0BFiJ9xXza+Sq4F4e/ANdmmn+vHiVQsnO7vOTWVvTsk
sd3cGpL/49Mh1vDlUZ9+DlGBUXTE4wr13UI55QLINaxQHMHK7DaxK5XDOkF3JuVF
`protect END_PROTECTED
