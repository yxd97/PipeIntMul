`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Phd0UykH9N/9F4axshJCk2Ar3M02vyBqIjk5ojSJSb0jPh720DJThXV/+XvwZc1/
KDQbhh6x71vOnxQhvsvQuZhAXkvyOoe7R3CjJNDLMj3S1a/figdI9JR2Su3yPQEr
aUgPw9haGBfTMAt2KOzL4XuEOFfXKzJEpZUFgkAvXE2ES5iFyxj1ao+P4uHRAU77
BmmN1RcIuZdP1xXeQFTdUNERozLfWZGeMAs9rb8tc5ZxFFVm2TezPPGRdkaawP1D
KtACokDZW65owt7QfhPpn/MPNUujMA7o0MdKCtEcF8tnpp1ZSvnOe2hFwFcHsWhQ
d0yyx3RIxHBx6/HkpshWvgwZUEDR0hSNoe0kKz7bLRBj+VagRKbcGFojKWYMppD3
nL9tPwf9MSSlZF4zV7kF6hQnlgMkGZ6Ms4BnXzKJVDgMYQwyJV5DY3BuU0cCKA6P
DCsJvnU5nKxmMwTeyjQsgAxWdiWUQyUR43utGwxh05uT0N61qKj0ZymQ2p+yfPY0
GUf1vMDs8QjT9SHiudlNviSFWqODuXoZ8+UYXO+5RdL9/O5A0tRTlt7t9eg08ecH
XoLzUjAtXKB8JspmqO/6rVrWU0ig3OfFL1HtxZJQf+ZnTbcShZZlqk1TA9o7gHos
HhS1g3xGhHb2CxPkTAHK/8Liuh0SwP5My22dA2pdZpFvIt30VgU0NON2xDzK6Mvb
w1qm0NyK8n93Dcy5Tnew8ZsV/fzhc3JhCa/JMCtl8Yo9e1F42CddOC3hQ2f9vYp8
TCreuErkrCK6dD9EOWDof9OpN8WgEkksBErk32mrOuqWGQ/bZ+iBVMOMPMjmwn5s
OIultsQX84Akngnl9c1xAfeWrqJMNc9hqLcdTsFK7NnNVVMbOdDIHnZwgI5pro+L
t2SoAH+RX0nOiWgSwNr7NPgbLf7IkW5ycN7dfJsvEsNamt4aFOwtIv5ia6rMT+c+
`protect END_PROTECTED
