`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/Wh3cFebBfFcqrOfLYSr7QYABrr8jwygnA/h+V6SRTVGPUjmpxWPn92GEBfLZBGw
M8gcH34keo5G3A8/CATmUd6G4tSYUekwXRPb9RskFL1Ey+QtoXokP/H42WL2M+Od
EtYDjJRcXRErV6bXWjcIuSFddZwUteYzxaP1891KE0wJC7uWC3y5fhNkp6iSNqhW
1mXcnsfeL1iaIOF09NsVEmyOLBSrOeNwbt6Yqx2iTgv1SCXs2cJ4Ad5u4mkbhp+D
YVzaDO3YtdrtIJ8E36iUFcHWP8UOCSh0qIrNHw0LMbDcdaYspf8DIxbAuFI5OUjX
8mSfPMi3e2mgDHQHrChfoxzQrGQhDcp8C9mWC9TDVYzxBZqaxFzzwMZmw6gv1s3g
Qn47xJgECwvfkzCU8aFW8k7Uzg2MZWDNM9Ix9TPE/RxiK4dgWs/STBNIQ2ZKQDWk
pcKTlsL1JDsHlvYiQOp001bhszwjLTfnmfDdoeRanKurmc4aew8tmrKdQavlVpd8
2ehju7EGGWR4xXAKbgo+1eNUvowjtA2gd3ngiw8uYNb8pyjJt3+xJVKCXG5fk7DQ
/A9U21s91lJf5SrG54d974zi4wtNGMPTKOUbASYZOyQxoczlUnIYjxCB6dLm9XWC
wP1ADdGlyEbm4spfvVo/tPB1Bt88BEMjuUnULBwqYGCK6kHtiswrGgVX99OaD8wJ
pfwm9R+sopYLw2jEmAAhHRqRCkuvlD7Rt9RxL/bafT4=
`protect END_PROTECTED
