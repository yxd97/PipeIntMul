`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
I12LVv9g8QmCkrXT+PGhWi+ZMyyyZabjY2tJJ6nslJ0jqtTT/2WDf+tOEpUBTdgu
jo61zdwxPPpitWDctrwVJ75v4/jZDYWY2z8IjccALOWswc7A80rg2BxTdj0zXiA5
FSuAKFqi18FMtopcQKcLmva4GaZWz4Skzoelo8vfK/T4AMcymFqMwegjzxe1q7og
UpZTlcfirvLxQhAYgTJTrvvBL7M0LXGZ6Wm6sTvZd23gpk9eU3qiLFSMFSGl0N3Z
y2oVZP+hX+cPJlEwlf3VOA==
`protect END_PROTECTED
