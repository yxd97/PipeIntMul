`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/N3Y+3IzxqoQVbViw4h7Pog0V8ui6z/TRsaweIM6FEngk1BAmjXstxg+KzxfX8NA
QDCZyrXPJ+Z7a0+Yng3Pj5zo/Gf+ZcYttDgMBT4dT8EN8TLPgmwEZkqZEkg4lwhZ
lt5oSpLoiv4uR5aJ/uTRoI5iJi6p6SwESt4M7jbCr75Db7O3/sbL3DKFudQKVF0s
aCYI7f2Ymci6juWDg0vt2ALAFq9iBwpIvYDVMiUBonnnxmh2SY/KNw/wFWt2cM7E
glnaRpnryTp7hNbIvkX6c6xMY7+qxozjwSXStQ3Wl8DGgBUQeyRrFrDl+0V3loHE
7qhW3lg6IGvnnVu2U1CG5hJK1PnlhnmQyFBgOFjNqnYx1++JH5J1hdWXV5Z9iPpC
DUSvHdlm9LgA1dQ5crVDVGIhi51i2S3sImrH70sA6XpqGhVV6JbdTVmbhtuJFsi/
sufeQGZin5cZx0IMAsodhJdX8DrxFI29gMOprle93+mzMWaOAU8Tcx/qgIemQoxP
SVZC1pjZxZ2UX64UHHXsYXLiBkqI9Y8Wc6BTxvbQUMGajnvBK5rwjrL6TzUmIgND
l0Zu2eKEW+vROhzawFIyszRAa09rKWVAa9IyLq+hKwgK02pdDTdk4tnNYM1aMXb5
1Vew48wCbL0qAX+318MSOB1nvPUXlHarjjjUYs+OSUfFE3hYOwDjDV7GcmmZfq17
SGOke7aiEXYWyd/xNyFrYCS4AkQOoz5AWT4bad5FcQqGY2oTzZPU96+Gm6kBZ2af
285bETz1OiZMr75Ya8r/Et9V9hj0elXW0yriExvnuyNRHXwdV9ds5bdfQ9ZDvztA
wV7iPLHHBCDrtQBg4ShfjdsNeIaeNLdErSQObSbEeLTnxoNlq8H8bVW98sU2WdnX
Uy++LNHXP0SHKPLLIfWvUxiQkUDF3PSQ9vnR1zDEP4NzvmEFlLVQX+QGiqH6i8OP
EBpE41C5pt5qohyILifs8ej9pNLPJRUFVCQ+pdeFdjuZEH8XsEjZ0eZ5U2xHv4a2
w9tqNPy9+0IJjo2G5HjJgBg/j7Y0lR4Iw4oelT8XPBqPz+mSSGr38uk7oa++c4jb
CG+9PC6i1D7/5fjcZKmrgYdzztR473ml4QUJP+hDhmRDjlHAAey7fTYhpOk/LhzE
VkCPn5Sh+Ms5MNGFbMmx5bcrSMedolaovzWN8Yyni5fe7A3CShNNnwzCKf/YUXa+
Q4lWoMLf3zKnCiWR85RzjPijX1QFr4VPbNqVOm3501yUytiQP/lUG2dfof+tuNGj
Mh+L78fWopdcA90k1NPUrMkvoByY3N6vAWvthBWdCMpgvm3huH0mhKnLR7/f+vDD
9TkweUwsVO9vK1RYtDIM9qI9RysRdtOsIY86LwS2qVApaLMQS+yQgE9Qx48X9Vpv
kMvKa586ePdekGEgbfb93jnQob3MddKmGo/w2LT5q8J60GKmIhiWXviW6c4TadTw
7JAUJVsZZjwcdYBGqn/MIxNsBmq8eDSvaJjjmVye8Pyw2MGuZ5jnYUgfBP9htuux
hNviHy7lWS7EZJX0ttiXY5ekBTK9Ckt+wtrAJl7Qrgd1OqzHkG2CyWTApLteaWtP
HVjVaqP2R82fK6Jm3euzh5aFwB3eqwMdH/oHMCzLcvp/fIEBZF0m8VpIFd79Kxp9
ynR3V2CcZHo7HCEnItk1uirIbuRZY8t3M4tzh0om2SRXedVYOSFPGVNnHiRmYuh4
2j5jnfKqlcur6l/RsxszFK0pW/sWlqICJxqee65SWqW5TwJBAORmIISnQtHRo4kq
7+6QoPaQx00s0RpjrpP5SAW8JggXa/bUVzF7BPLXpwhrrRn4VHe3a7XqpnXuwf2G
RCLDGHqVAuunG0GN6mRurrTR/1Ebz1gF+qOPD166yalP2eGpigE5r9gllYfCqPgE
7dsyukaj2pL0N+JhWBl4XeyfjXY80ncJdcSuKFleFSdTwU675T/Lt9C2ZkyLTOYn
T20OSce1FsxGXvHSCMNu7otBi3EDIFha974D0lrzXvxbgihAcXd4A+S3fopRPiSd
ZJNv5f4Zs6EAPMPUSZw715KEMW3IPiPMzJQ60+oQF18mALtCV4wq9xPsbda+i5pg
l//kEfvxhTnJWUGd9eUl7gXZ2cEszVCXeeYodgqaimh92q/wY3eypOOv3fLNdpEa
9Ig4gWFLOoKmcyOpGjydFiXqf97/fMSeHr/RsvMVDwCicHazXQZYqc7Cdyw7Se+8
pJQtREkqkP6WWONsDgGInMnzKlgxgjmF5NOZQHm5OaMwJwxktabuenr/4A50uxpF
w1Me2zwQbac+nfv0cetZqURL9fkin01HL57orclgHazp4mcxw2HjcxyuEnjIfQwS
TtwEbA/nsXJEWNXjOuR6YbV2V8zrsOmkpLtvltGNilTfwCfcJaXFtjzX1duGMRrh
NBmybbNQv0fUxyjbKOxKOmbVrIH5qyGKh6dOwFj24Mdi+6vxLSuqD9BSgADK3NNY
mRFC//I0hHrEYeWZW+Ai/HKT85d8nBxM5gumRFKOiNGr9IgVTicEdHsF11L2xEmh
iF+9brvDjvUtar4N3vwVnND4ELzUTPPmetoyglmy1pTNe1j+hycA3mxbQrLxKCLE
eLjMiLoshQkAoQh0kieDgfq0aONiCgJiWLZJRxlLxlmNvzvxXDkQACN4L/gdoJ3+
aDELW6SuvdCXWDq0xP8LjdTibCxaD9k63JOlSWSwTRH/Gl0cc8YzvkS8/L2R6W9o
ON24rzq1xQeTMpqLGm8gAOo6NNEvQS/eZVksO2huXmcLKRgy/oDqQYhaAQlnbAWk
eW2JsDJvI+S+UP01o3Ciw4grSThiWsbz2tM82V/KfjfJ0RRSBPwhXYgcxfrk3Xlw
6TQYKUn37b0i0By9NeAB13U3P6sSmO7u/m1A0+IzRfc4PMATk4YmqMR1k4v9cGrW
k1TH9vxxnSOGObUSmH8l1wc5mTdj80uSV0HKT32m2FrwCzFnRcFdnZB7TMsVN6aq
CMQfZnTMGlX+Kw94GFG+xrDnZ+g6jbS0Yg8r2CwsJO1kYa+8mA28S3Pht0ilCcS2
sPcQYD34+oAtYLDu4kEWtxPGwIg4byLEYmIRg8zqqS0EHCs+o3deU2EYfPGDjuAr
H79rbTOCHs35IfQDpupG6tYcGiVzcd5nH//+8D8NuoOKmz1fDFBRcUgaueRTCLnf
0I3qo8nDbwOBdf2wGvTBCJds7s46bwTwOrImE2NyLfZHKO5NF5lNE2AWHAfd9t51
o0/wOkScodE6aVXC9MXH4WcrMyEUXDmvOyFGoXuj3qhxoIYOiNgv9hAfNwmBt4wf
ttUt34nIEvKPlyOnaRNgqKkMXaTZig+oGydw8fso+d+fMuhZk1TlZlSMxw5NCLeq
84VJyxfx1KasUy200TpYAvi0jvYZww5hYEtSqlgyce8JaxrKiy8ceQOvKjdABSqb
815OeWaVXRvBPucEbIW03yS3V2fUKcKygeV5mDc1HhRXNxbHjmX2N8+GbPZNEqF9
ny1+LF6n49c65TRxUcnXIK1ECNJMr/gzmzQq4gHIQOKPUSym5Z1++i0xj+lRCUFx
oHNvKo0s85aliWQaH7yU7oO0zJxscnikveM9O8tAWfmRssV5ruroEEd+/GEL0H7t
qJ+WXA73QduEgzcSYdy3rynGUGtdYrDhn+4Unp3LltON/kPpgQODC/yCCJOtVmnx
1qZ9hb0EhbLMpL7FbiQol84UmMAH+0jVFhOYEsOTpAGShc+iKg9oD/Si4RGyJ/9x
BInTaAoSzTllzrNVW8te0jM/YZAlpR50l99h7EeuqcKIsIUAxEO56d30PpQxLBoU
zRQkLPvuHL+gX1BLKBxGmYAI0oEtmH10JHOGHs0rDTzsp9D66I7F4kp2BizyP5xM
5dohG8rTgoJ7pU2hzzEZa/e4zKZ6tr0SS/rpEuhfh160s3vUjEYYc/WbOs1VlkEV
h2JBy0LQ7/HYuhRft31IbIiXcXRmF0gCYa2cST7UBzDxh2TAkd6C3X5MljeUSF78
pJEMn9tEa2Lyy1gVpn6IePNKvCrNj5EorcDgHsNydoeh7zz0pqiWW3DQsi89UBUj
WdqM321lfdTnmsg/ckIIQt/H3tSU0L/feexD/zLZnedfid6Adqrf4t1hUUG7cRx1
Q0sV+hPbdrk9TmXZ0XUKfo79tsK6JEjRf6DfhXE73CyaSmNCYGO1uGFNDKaT1gJs
BU3Izq0Ixv5DBKsULxbJakBO0GXnrg9kzyREp4tMbFcAUwy4yxpxtV1BhXNbxo8b
IOeRNVZDMcd4LV6JTcZ7EWhiGGtuM+XBm8b7EIiEK4JoTbpnIa3oFReVv8DZBJ8p
hKgyWJi8ExsXMqc+fRglshALULmXBY6ZAyLEB7VQnmTnKCXSpXgoWhdpN/vOvKX9
JDNEfO+16ehwv94+T4FTP0kIqrH/Ppxy0q7SV8AqOMC5dz0ZQqO6zdhD5gvxjIuj
88j5tZ7+c+mO9bhqdN4YMqW0IXmTI20sIhHyhCWAbLw4Z/lYwEzJpSReux+pGf9x
foJzDMCAUFpeRlc/aKOfH0s+1saz+DR141tFAJlnySFRphDj86vQPbufdZbEeQ3N
qEYHc5h6WQLlZFcTuzGYnchDyA9ZJKbgguszIilFougznpm6aye3dz6OrW9KX+Ho
EtiQZOpWoEIyzbZL2H1LSzogoEq66M5ry/qpd2eWHmPQ0X6hd+Q8Dk7zFUd3y15z
UuHozmB7sdCJInrmlgJnYnGcqvvcg5x08Tc2gKz9opuYv/rnSZ7lZ/LUzLoGwR1a
VkXtXvAGOGvkSq4PKu0iogg3LxHy/Gh3mQsl9HNbQYFHI+MqUrMz9LSmnhg94kTY
wXI4iOOpiopBn5lDPiIWghkaFpjpjYHy5KQ9IHqMeZnocVMhSZp/0Lnv0gnfsGMk
uhcUGo9PZLDfrw3YvpfmHmu50vYGRilInKPqfpH3N6Si3NQEvMXv9Ta9rDgJ4v0m
p6DDhaCZ2RwHLQZDfYEq4pFVDL9jQ+m+elyVuA9g5Ay2LcdPmzzME9d/AEL5GKF5
WhzVVwZOSzrhQ2yATjE7k+qZJ9rwfzfoII2sA5+H5+qbZj9alqh1UCFUVy+BDPE3
rp3Wo4XORD2ddtLTVK8SiT5sFDauHuCJ1pR6i5podiA/btXNj9BgfXdS2y7JRMdY
YMxkMfqJI7vjJFsxWppU/Urv4reG0X3Nkac5X8+7aHXkH9mmiiNLloonSVfDZhpr
FAdJ86m7OhVD0yQnz/k8xqXW8b7KNEx/3oSufsM9KDKJEsSQoRotLaMU/Jbks5TF
NQTjJUdlaFKudAw0yOSy5WKbiKmgHArnYo8HCKMd3XyU7egEusqnQr3LnLLD30p2
pbJuyjM/Clz0X+XXeQCBNn71Jc/TwsSzV2BtBgYZZ3PtKzpHKZYCsFHsuEzre7Xa
B+GwN4MOs7Fv8L9PKCrvp8p5ZjWDj+AXjj7VI9+aDq6YQs5gsaxO0mAeeK80BKoN
nGGqSPxDYnqeGrQn+CbT6EVU2Hs1Za5bY2MGbPNrV7hAWzhs3fhWHXwfKEMxk82O
UHT5P1aO8EpBEbR2uXpymSZSlalm04h3oMTMEhEKDaO5zOOhGgmqnhiftGJ2LhnH
+8Gj+ymHx1qAX3mUuh9xvE0ymD5RYeoSM70m/HZBEaUXdEpshfSrRSEM/Gr5hoel
kFBsX1cJ5IVJOyOsyWWSiYZ04irwqZIjEj6kHgO7DNuBc3B2uTUmogCUbxEd7nVu
F42riUTfKYl9ONwTlzE+lXUKcXmZwBzgxkvVzXS61cuQg/vWewB21JdY8fE3cHkR
Yv+X0DO0zNT1V5JQsXxwgz3dsS0Q4ZlLhsVeqyB7UniMvakqs1EGnZgENwJfPFsU
PdUhqGIQTQrx3EXO1+/zjXX2qW/NBtaTuRNYvKi/4bohyIWNMG9p+VKOZDGaK9Z3
uHAQ5XLKrZmey28BDBIJf6h1SD3zL1Mb/mFBsTy4gWK1p5eDDVOuSczofb63UbN4
g5rQPOB0n0PQX2h0aquWimdjv2I6F9XeLZFp58c/iYfr14W0x51BCqWGfIZNZeJz
FZbdEvp4EdHn9jHSoE/fVe+GYWQBKgpOe0+NMppEp5ha+6gpoZMiG189g7WkqfN5
7F6n0DspiZ4G9zpPcX+lMaWNTMm8sbGfZeh74vDy87xNRvFRqlCLo/FEb4ZQoMyr
Q/1FCpzmXF2oT+qGLkevRBvaKMu/WrkQ5zeYc055xmgYooRL8SRFVlxN7VR2mMxQ
ej/z3Qi3PRyn1DlmXqo1A5boPSoX85tb9e6tsxzwUBYP8rI9bscagv2bWphZiWgD
ubnNlFC25N1mX0kQomUKZrQFdmKXe2y77hoDiXcuBMapBdPk5CyiJGdMfwB0l6nW
y33fWcdJjO8D+OhciFJTW1HgjKSAnSPHWiuNYotA6n+gxynOUB+HvOMJucJc54RC
OrR/1UJ5H/pN2Jta9dY6G0biurhUAnUABDDk+40csDdcai1jRjOAjNsfLYz0BHr+
QFn1jmQti9itrVNw34EW7g9+xfXu7AsXzkJpnbyLyuuLinEC48c8mDbKIhFLZfM5
xwSph0l4ThzhJfvGiiOs7pwB7wKou9szv3GCiZUcgHOhYdtERb+UJFkYVTuOiFau
wKg227dDxW8q2gH4al01Eb8+ABKQUVuzpXNtirKudZkP9IHQpvDW7kzAuIG2zspI
YYbHdIey1lgTmeQ64sRLpq0JNMwzuPYjT89ASt+j/QW8lWeLnm6rwc2pB4Br1kLR
mz9gw7Ly+TRl6/zxGnVAok6p+rUKdG3vREqRQHHQMCC+nfP1Zsd9/bJe9ZG1Ub3c
dYKSQpSnsQOiN8/SSIE+HrTLkayfZhlPfrYe5kJEByU+6FuYSZ7hsLmgAA+atVve
N9PlpYrw/6UrBYm/PHKU/c1mvzifIIR/uZJjBxmVipErpg5DExLIcFQrZMiwyAQB
hww1v2xNlhd4bl+EEfSyW7qAHYOJE68ohgKyEbfvrK1Jk38+dXPHNDZnaPPJsfgL
fvUh+iMbZLf9x5odCQ0cbD3WqlKLmuuWujRs0P3V1DNwIbqOMmvh3uORJxmAQATn
5V3ShR0GZqrput+C+zQpXDRYhkk9Bs2k2r91NSRoHs01JnNmCQgnEye9JVSJdVtg
uHE9PlKm0KpXLlLgNMGKTyEUiiS2tisXoHRM/kQeHQ7sCkd/Ua3ogxxBQ5CHp0D5
uZjNLyM0N0yhp3fHF8Tl8BiRKIMAP3QSUNaaakBbXNM1KaTE5qWiwPXnphJeNzZh
Moxi6R5qV0N0uIzWisxMnkTBDfXTz1hdvLT4V9+eIXhTJc8e5dZprFQ16cvPydy+
9awfc3aqrfrF2cQbgL/ogao/1M9SiYx/NdZYUTS521adDtQsrCCCojGCXC4zyJST
1AzlJQRvnCiHbpN5T8cFlJaqO1pMhp5w7ShxRIDumcIg/HlcPOdYMTwqowvBTrg7
TIhYsH9BWgw0Q9v3GacgxE+AK4tauxh75MSX70kAwkKZZVUAz7zW2APknNNy11GC
4xLE1y+7DWGAPy9kzcl7BvU/KQWcrsSrQ37L/Ukp5lHjQAniEl+1VwYNnegtc7zf
sUHakPPY8iEu+RGdwFVLOkpfT9vAgn1H4uovcLl5EpOi+L49OK91TmM70Z0RM9Q8
PqXNi2redNQ6ao9TxDWx5z+9rekmqEcJJ0YaOm0zzwnHx4rIzA+83vMlr287+SNn
O3MuBtaP0naoMVtHJZhhKiU8Mu3Yriz8HQMSsmRObCQtg4AGu7W8KBKAZQvv8PiB
bqsG8I46q5/FQBqOAGDZdn0qEIMN7d7ka0Wfj19mIVkADm5zCLSdS1foCkrbasPv
PIfjpro6nBrVvlHvSktGxiBK9aIpsFMvTA9HBpi44omN2fCVosONp6Iax1htMsIr
aDuOM5Jwgp+mhSCU26zku+8pOO3BjucM8e2QXAkbzVg1YWGdJjyxVjEXrXYNl6l1
Hgm0/NKhLybdzdjefuG5318LSZdwdtjEcUplqw79HDo2F1Yi5Aw44t2KNqrGV+Uz
PrtLb5zPzom9ve90/Da8GbcmO0iCo7aD7ub2KnQNCiIlDd3uT1wiMG4CwbblIkNt
785rK4UGsqukqMUHStsnbZn4x0CyM5glEwkg35Qda23WLmC7jD2fzyTSITpX6zwP
JlGPD45MmrjFIum/hcQxqpEyOxs8YE7AI0O+zyUYZB1KT89Kq7gpm/+a0iFlfLSu
WEIGglxik2gll0Fkc0kbcRcWHE4evxh8SSq+y4Ga8TTXjJWEunN80TxvVvf9Zk5h
7uwC4oMuBZbE/xkq8mWa4BeX6H4WVm8NU3F52VXxvqMK64qzYZFu2fHOOzpJbq9E
mBELLykAOThtx0CVecGBq6227Oh0bE2H1mKEuksiAreOjPWcnUrQvxbQrwdHqMq8
CwGQdpCg6411ns1uQN2M78QqPMPS4TNW3zS0jWdzehTB30ik63HMfzY5sHSYHzjG
aFU0WUxqZHRgUij83/DRSQqJDYvWeYZCJ/PM8okY3CevkMfjFFCYjD75vEq8CNGE
nlDrMEUPpTWoubJftR/nEa3Q7wW0s9N8ja+nZZ7e72CbollUDDecyvCs9YkDZnga
E/o/UMq4wra5gC2mGZUAVh55s/KzkpLnMjJL21B/zmutlCzVH5V2yRGkn7CGtl8h
EP+IsUl3AOlFUVdIXWfacTXimjUV8D6Kc3S0P3g4ps7zyc9PaLBRWXke2XsqOO9W
rJ27MXt4J6b03a+Y11QJW5u/BOE5ebziIbXDn91L7z9BlfRzOn0ddUwiVKIOyz6z
bvs422Ci0GAgwx3tO1mY2p/G8E8ng1YdcCAuU7OiRipbl/bqu6mzLWCzWZNCCCEo
bE9mCiICgWHR+AwbLIuCX+ovezKebmbvcfFKAzG5kHKYE+AW8teuSEpJe8y4grrn
6S4huYfwXN3KtxIOHeOz+DC8D5PzjSuGQuIbsC/ngCbHkbPZ9DI5o6bmgm8W2f3J
esk1LFdtWaMWR4LZC/aIIn1D9Px3HjFL+Ni/JvC/AUrYIDgjIihzJyWi6C9+4cd7
Xqb+Gu2hR7e2drvoXJerlRifpKdJqGaLIapaEWuZAzu8rEb3nTJc2B5Cg1q5xai+
exUD0h42jZ4nCV7nShIEet7KwtURU7CezRCXSd3WVPB9ECtpsnHIcp8IOZU0Kmxz
fzTjfp9qThJnAhmFGAwQ2x+5+yOkZCpdvYS6qVqtnjhWS3xdt+2tKTAnnOLsjQqW
qeTyllQIE0YyiEOlsD9ENf900UZRQioVjG2VW10ldR6irajzYdz9gZkrXPT8iHAe
fqmA/ooQYxs/SS4LK2RTW98zpIsL21WrV0AHruOo4sZumq7P8qbQlVghXA84iEVD
ZC1cuMLphY7YN385581OlIv87LzeBCG2oD4OikuhmF05Bd+3Q2Y83GS4mSm4TLTZ
k7yLKcKzK5AO4e/zI9ssy6dSZ/IXp4A8llCE7A3Vnml4teKLO5Kk2XqFOX5FEFV4
RnPsxgvvGbctXxVc1D8Ee7XKHQ3Dn8xihWFX8qi/T0mI3PLzBZfqDy18PU0E3WFF
p/VkbkXx5UWZqBNICBeaUrT7iqEWzlF4g5vpvbpo+uRi5ralTDF2p5HsLB41BdKt
3BCe89O9PlcLLGHMkJTzluSMlL4NxfxlyJ8Tkx+I/nlwEmetuSKDDFanfWQH+/rX
gBzDvpHFR+9f59kW/tE0ZsyPIMsHQqyfgserDEz2VJYgkPTq5B+MiMyBgcx6mueI
8mclxU8/qyNGds3GJQZEkmNvOiXO9xBOuDqKsgNnbd8hhvNubT7qs2ok4G7mW1NK
AQq9XuG0eN31WT3P9ny4jwVIqe/vlqQoRo0Gw2un8Doh0aRDWjbS47pKR98y3aLY
/600KoB2XwU9aUVv/VaipDfYdCxkCG+/DMAselG1z+I1YrDeTM+26C+LwH4QmlcU
C5vx6R4X/1xEe8uk3IMMYvR2jH5L1d6qZa2MxKjQL65dvC2U1+W/YdQLswOVpiqw
iM3O/l7e9JO6BHEzdm/DoZ98LvCqbFN1a1pHohIrcG1hiGojPZFYRqq2m0MoUzx8
hKW6THldLCOgSoNtTi89E5HrtetvHtzFTQcSE+a7lYPHdL1g2AyaBvW7EiN3g6w2
K1o6Us405leIk2b8fjNa0W09nBR7a54UyIsnAu5S0q19VrVL90AScM1bDh0OBlW9
DMRKHWLJvQOiiWm5mKl/obmgm4aCc4pxueTQb8ZRVMVVjyN9TMHTIKrAQfFVpGye
X2PMAANYQwkRyTm3exMv6HRWZYiYOYOwljVHr8//0LCgl/78bt6dGBlBgQnjKcwv
dJ1b7w9zogJJf1TIQpBGZ0l7m+nlAu79Sc3hRZuwFm4i6wBUof+3Hhfbwonb0QbR
4ycfMfhaVs95j+CgSuLAEFl2Be7ERIC/9kfj6Q0KP11LeNUUWdrPSaiQKCvwxxLR
GTQ1eplwPJGdvXMHA7AiaDST7MdEpAcLtoYuZt4hun1ypb6QFJo6iIpiSmzrz2Wb
UnjdqALBSOvUAD9WcLB2QCXrL5vQMB9OIm6fdNeA1JgVcAQfOUe1snAerfrtiLSQ
KscqULnoZPzJpbxJ6AAj70Zs4kdCztj2aF3LCDiH7Q/KQrQEQxpSYeWJwfJ9aH7r
W/sr+6k+n+ADuY/qSjVz+0s9D742ENiQbWj+uON3uNVZ4m2fgDP0DJS4I++nWZmH
woL4K0QGZeyp6r8SEHrpPYUVfn+FHMu63Hhvw0YtZKSuP5zRCzcizt7lGeiT7IJp
IdXBwi+dwCYe8HpO6Tss/SEC3UNhS9MhZB3dNWl5MYrAVTj1Z+4NfTH5u1caeFh4
ZhcP8J0QTPHwAVOraff16z7OJe28Q52k7kOXu2FiOgIeW23nWQgAMDA5MB0gsjdw
pnVnLqmCuv6UBuetEZ6g060wAbiFV03rfccBoifubSUwauBtp0tXb5lUfGu8GXzN
edppxdvKyEYZP/RVPOyp2X4ncSxZ/ozpMAiQV5gdaq7PJzlpVXtyblvd0M5dc1KS
SXkONiVZJfgvtIlxO7duanGWxcgSetJreQirvk1lCPy8j93xaxQvajeIlAUz2HCC
YO42GyWdN9SwyS5hhrMnWB35TUTAmsiZVwPrguJcKH1fMCvJUsdlGLVuWEbk46Ur
tHwUAKW15IvHayUEHwkYwQrkpTAdPwG++tAUBBhwvp2fdmw5mvy4KpFaq0TNvaX8
9jC4693XCjlmw+fO8S4tCsmrYKpepjZsXtxxFgm3E1UBilKw+KuJJYQijODphkdE
oOPAjwvpY68Y8z21xcIrUoT3gxcRFP6SxVXLvbv6mnUhTVsJHteusccjxNblqxRg
zpc9tHCOQKLfGXsSq3axcSvOWT1Edb6hKCCaXBLiNsamiTNfDfxP3b7pYYDkC7H/
1n9C2md5p/JFqCeyKcEoaPrvvIowXeKGHaGkg73G9q9cAJYtagMFOpAgz1o/kTGr
6OOXPggqhTcCM4PkTIrkSVOuiy1n8s71JFbjeXorjmZJEZaMk4oZ6oP5kSHizSqV
wwgx/KCpzSbkV+2t+6LtOt8tLHW8mbiqhLN5KoaD2Swocc+xRzH8LTcPRau1qtUG
eOQAt9y7kZxyC+uX89ReRXv5sKCLiQjXU90NOpKDyBjJUQGBcO1FhnoRQnK2Ouz0
uQJ2pbXjqFeAQvLIY8nLc0acvX7OrQCyFF2w/gI/p+gFCd+tjUy+RBms7k+e2zPa
/tM2LsJM1IdI6BWZJEBoMWCZi3RsEmw8gKSCGUOs+ZDn11y9w02eTqLcBJAomO9v
cYgtBCIv7nVCHyPZ+hV7gKNYSqv2sB3ucsF06FUFxwVAmugQxIc2FGbKYB12Gmce
8SedycRkpgUGaZhdQr/p709p1s0zMp09Nn9SW4Vxd8gm5u5HNu9Wmvy7iDSDGOjO
5r4zuKQUfTX7lbX2ei6kbpFC1OD5vtEkoMtWh7zCVnTIpL8Zjke5dXDFeLwVVAi9
Odz599TRvEU6p24dJC/NIyhh2it8jdiq/JvVc/VSHD+OtPLvBYgqmOeswjj89ty7
9HUIdra5XDw1pcyxThh4/nyTZmX9r9N9xQZVipKurNK54Fftq0zl/inEmwyHQyW3
ixhRj2CKPYUcG2/sXuFarRVjpNdg/hSdIJdzE/M9eWqD72IiDfzf9BnOv5YnPaIE
Gr0lSGHwiOY1FiG5joxhKYVN3L0AhtnPIEpBEl45S67LjMqUuwqbuwKk82PQCir2
a6sJBhH5k/EWhwnEtZyhnLkEZ4o6JXNTzZM1omWweGeTYpfWtYcuf0SRH5NcjYV2
nmKPOgzPSNzar0FLn/k+kKkK9EjUTkyVLNFQII4N5C8IPib+n2IHnGTFdXtKBUKc
6nEzLW72hEw+gflzB+WSXjy8h7GUx/xM8FM/6wM0xhr//UJuaZ9kcmlr5ZAWLTTg
44jtc3ZwHc9b0i+9d+Cxm9mx5O74QnHftTzqJD+/bNxNzgg0G2ffrTgRPqycz9nJ
rrVA7V0xtP6ex1Nqb4kfgJdDs+RrL49d3NJDo7WyLcRfJ6MbB4dGURHem7+JgBUD
6tGdVOh3xmwHiOMp3lJbpbt49IHVg+YZJ050FTXqHYScDna9z/YDXgwyVAcFvNvZ
iNvm/44IFJX8BbPM+HIXscUCUVESef6MH/T8FIc+n4gib/9O7f7nRCbrEI2enYlm
p2TvZbaQXAeNscUQ2D9t+3NctGvbQY44/BXv8J3NEPvfr3eveXp0uG8vE/5fT4pz
1Lf3n9bfQJHq9dZM5WLzWsqzkAiE72OjlceEENyQ4cX4y+lVPvao2/74/6giE043
Zi1BfZaIhnBwhg8z5E52rBZGH8ktQcghjzTlXxoj56Cwj9UlUPnEqi9NJTPR7t1C
r0IIk8UOet5eKvAsoZRIBtC8R8SSr9hZCfnn8sQCRnFWOQuQwfEJYMVl+cNtHkSe
wBVm8QU5uQDhv3+TecqQ1So+APHlH6EWsKG0PauWQH53SIIDkCUSBT2TcNnJ0v0e
Tf4FbwmWJm+L+Zon/BLUDbzZJDp6QtVnhp6oAvUeEcavv89xScQ2USwdYHvIxwfc
b9uceRilzFwjdJLpBQz6SU0jmkpJQDzmArTpf+1Hmg5Ydkwp0nUAF9UUR07V7Tfi
jv82g8cA0BsxkZllwHuxlAYy9rtbzK2swv02So/9ejtBJrl8xNIu/+0ciN4aAwbU
xDewP7szor3WvIL/wRq+uHDjyXUpn02+iAjN9ZZwuKq3MZT9xNew87+9Z84sng01
2uSgFIZrJeNvJ2InIjiLYK6ibxnGRoG7/mrzKpKE2ELa+GTE936fybb1pEYKMSS+
NEYMvF5c3acqlLCkjYFDwxVmuQklRCQ8z7u5Mr/wb9dJsb+a1ewDmABN0xMFnkav
EVyqnygL8ontZe8raG1qcLid2nZ2gavlysvLDIWMTjW3W9c22Htb7Vc74P53k3g+
lVDw5TAqsTHKkdk23snswPDK05w7a7tBXRz9V43ro/uU7oU2eQgB+5YdAkoM4gnf
nMi+pT5bCwsttsfJMCzruWgUg23VxxCToriC2BSTJ0BsucPClNwgPMHAJkeOa14l
vNj4DH5/4LDO6L4JVaeAbIoMsvUtpz5IFHYsibcrBlLFLalPBnQeHbn9IJzBzGsx
0Y+k/7MSFn8ADUDJfcm4CRVmUH1Zf0E2njlE7cUSsAvo1DMMn98C1tbC4ngfHa9D
PPfJs1r8TW/SF1HIMWHoqqWBqMfmUlNAW4TKDsZplB7A7EkfIuyg1Szcmsi+FEST
QJ8xzo4ZmkMCsInJIq4N6eQ3Bu/ZHJdBYL2MJOcHMGM8aNcDo0n7uALoWN19wR4Z
M005lw8kXbBPfMEOuyGueiL8DjE7HjNcPXxx1xGGlva+ilcnx7ys/kWZJklk3a7q
K7w9lUZrCkJwVXd9jb22jFJ4PKvvufePN41igZLQxk8JpWl411Xp2cIJvzg2fqIT
c+jQjaTBelt8Pfkk2UO0MCiMHSn8BMsqFJBYJL03Z+qPBca4ads6g8o7F4utxn2S
e0Wi9aQppI43cMV5Eb1pBwU/ZUg0owF2QP9gUYZb0EWLWKPPjw2J1tioxkti8ES4
LWLxFzzPA3r0aui9NF3NSjfB1Cm8rTumQ3ThU761UaPU0HYc6qWyEO9e/Rokq2Kv
ycarcx5JkH2d8FX6wO2Tr+j3TQ7yGOp7Nwl6mmYNY4MpZa9zZalOJahw08DnLr45
PE+XTla4lVIemvFoQqvpGOHrurRVY50mhlqVc7zUibndRi+Q1GBWKWZX8gKMq2Bs
FLXY0ygehY0v8Asn2jZXmppztg09mpjNA4tdbXshZkv/+9BbbMCIjST/F+bzAclh
uu8HTMlOD3zSLpbe89lHYF7Jrv96tRLNC4+e4o0f8MzqxrL5rxnFSxu1QSt06NrW
vA6v0/fVoUb5wLTGtmWmY2NIPNOZiDkxaXlbdyRPVxgkz4Yor2vhpwm0NfJXoF/6
EWiOwTLjxpL9UqRhsBt6+90twj0aaL619UmLZPPpoVAzv/CzKCLm/5CBhkq6fI3E
1h8R32v5WvNrPjLCAuw/CLI9lpfUi2XHUHcjst27qg73zckuin87Fdgc4O8nJrph
tyKtynN69H97FSLRjgQsdiTrMl3/apkCqmOo5lpZKLICcGRK7WGKRv0qGqrAz+FI
QQFG1AVyTrl1BPzlDWSZPrjtUPRs86XIU9GMto/zTMdsJq2Wi8mYeL7VazKoKLRU
+E9aZF15peUYO3LdEHe8/RtS3c5BaUQe9OWJNN4HRqjOXkyewHJMJeVIJlZLmgn8
RhIIbr7SqDnFRQQlVu4o6TDoExgVlcRMjyMIhubkoY1eMeZIvFkH3XM0kyweqpaQ
Nu36EU47GaGzTvyM9Nr2LDVJVGNMLXjFxAg9dIP3fOHP3U9n0C4krAgL8eyl4eTp
TMi/dlzYvHKf0xGDNtF4jTuSyxeIabbj/REMpwntSGWeHbo9ua2XLQ5amT2kNkHc
nQ0F+2Vh5waJY+4uYoO5pgtwcAdXtS9uLz7AE8xiTzaH4OYtOUYTjmhf11CKjVk0
3lEfLsudgjDkgxykM1j/hZf2gZZZEZZZwIXiIPZBAD+Ie/Ze9zHgI+ZLRTbLwUGm
0CTWsDXTnOykGrd7BbUbPwjO/9GUNamsGVdtBNmtZEgNNlErm8VcBDpBbpMhAXGh
9TGXg0oFIUyPVekL2TJ7sY7qgmeuoCJ+XBwB4O4NIkz3ghEQZuUSEHsEs+2r6uWu
eBdu75t5lQVgrB/YFIzu1ws6ggHFKdzoZgDr6RAMJgM917RMI2Ujx64ZhHsn4jqK
JmfBKpkvMtXD5RcZ2vH2gu4MnbAnITuCXwemMk7iBdmBnmCK2VIVBt9fd2aHHagq
wsLKE4kCbgrgpLxApCjOVUJVDBxm6SIcIWKf2ryy8cloYeHHVXjZtqsYwS5RGqVq
ksSn+yZ/5OhqFlIX4oVwADTncVUrL1XFeIka1AwnSki2b+acvwPaAgJUBtwSNnBr
wFfmHciaa58vUv85H0kULIOv2CTtOUuX5yo86JF6XKeZXVfrTTRpVQJXjv1Cvnxg
lOw2n/Znj10hPhZ9PZJAkIku2lKUN/5cZ571G5q2EWrBIWShe0sRGHiXkQImPsd4
r/JLOKLKwyLLmykg4qtEy7ifWcoplmwJhMuuX5OOwD3UXjWr7Aa6/AUANZTq1OyW
2v6ZFyfSsouaGQpFd5gzUwmmuCT/SPOIpQlsr4NIUq+lEkw55w827uIny8O6mlFn
v1SwhZ4A6LY4aoWvbQ+dSsFKWn/a+gb5lp3LBJz+YMuA+BcA3VGQEUku1b0cmZZ5
EL06qzKq8GDU2BoDs9TSxxDCT6RBDiZdWKExuB9mths5LyA/9hWd/wN5XHbMbwVL
l6cCrAsUgC3qTAoduvGy9OA6YA0PnnKWvDtOYfMcP6esn+bsC+1425CXPzk4oDwk
MMfC8NyFWCUOvdfXo94l2ihyUPmf0yjj0sGSZLHUKsFyyKbA3JTkWJfQ6wgxsRcW
IKmSccmFBExz5wBmbXYt+NAXWEB+17LOfF6DGkSZLGIPl4fgYBLMH39oz/PNvZmc
U4g2ksPAxIShpsqtjIgU7maHzzVcigmCj6Yw+BvwL5NF1Y1G3DwPH7hzYFgaLpXj
k7h7KLeEvaoXMY8l18SXuV5e0WkddPxTOnCiYirQZL2lcD6naeLY4xMZm8CrC1mR
4/dpy6BnJZysvdVNbmjHGTRUAN42AReM9G8tD6sjMqVr/XaBMhfxGH43zbDTOV5d
Md5Oycnroejylw6kJScD324zSO+XotE73c5JulvjPwCJKEQIshBqxh5qQuKzOETC
AWDFpm6icBVmUWN5TcXNVk53uHYpGy/Vlm74VH0i/xj1Nd3C0DsK9g1nGRwyHGkd
n7MU8PTygjc9B8tFMdBNFEy3UNxDDB/bbzye8ufX7TdMcpq63XofWXgcZyJDafCx
aXmKXhYHZm6pIbtdR68xibGyP178Vz/MawmNCPKbkqcC4jRM8SNxU+KchKzmB31r
uIgzT7qlURC6P8tM1pYMXFpQlBG+z1HSnu5yG981glCLGAtxuGcjPgGfeQfzUnXD
sXif6JbS4eyInZgC/wUAhrwASVNbnfeiuyMQakC47nJ/VO7gn1KkLgLxDqroHdWF
BO62Pz+XGdZBSgxWGWvNoLZc+Y6GXWb3kJpDuAomrfS/OrcNWtXooG48/+S+r1i+
YvNuiMuvdJRA0D7c4UxGoOIOcpE8O0gxmo7HtY1CUqneNVNFFJSwNBleZEj+q64y
WrZRvVZ7VFLaR+0P36BXWFVeVLN1OuUymtBoCnq08uMq7EqLEwc5R5BI6StG8tY2
Elb8pnYboW4euoYbdPrNxOSl5R1UMMCgC7uEEfyyALWekUhA1klcppki5fQGE08K
UJEXsVS85dHJLXapJH+UegewA5lVWgCuZdjJ2gG8Mb2ARCspl/VUNJYy4DyZPYvs
/JOO1uEwQmEHRJHPGF4co26sPeE0dcKNfrmBXd97dW7tvdFQtcdtXs5Ri3bGEzyf
Aq0X7keBOE7ENDIVwpn3rn8xXuP/jBFK9lOKyrfUHAhnMyum6FeLLaICqCtbi3jB
YiSim+3FVRZabsJdxTyUfNgL8YHi1PZmH+DBOUsyOLDXpVDvC7f56R6Q9ITbMuNL
8vmKdI4oYWNVDvA19CEwAxsgtI/ZEPHKFbpEOIG+LKRUS/ByRE2m0zbmH4sIdAae
ViViJ+GPYIhiuTTpZFYquA0NAii2mvBSmYsRquvFzDMjo+KjaS82XkRrczGLRU66
/F8wBS/y/GFU3aNq3Ljxjezo8gPgq/ZVNI9HbGXVqQj5/aYrgj8VPQ5w8xujiNl3
+seqaOK8fMSg/dfSI4EgamBbIXvBcF4BnuteFMnJBZ2GDcFaz0mVJkyMwmHaeQ1J
nLxJwiELalVCjl2H0TPxFHyMVQUNGMvYUcH61tcp24euJkM2nLM3CazeZ/ncV/Qz
hMfNo/bth5TaXQKMh3kguVue7+W2NvKnZGDngZuJC6qMk8IRKyE2oTLi1LZP3EC4
JZN88eEIQ30yfZBKoCVv/sSatNYhD9IVqujzun7+5exGZt2z2YI/iZ7aIEpU40/v
NTt3bpxizNOC9JMrSk6y2Rb1BUV3By84pTIXTbQ8bLpznQohMCsCjvPauyNWEEld
bHRbWWdhtkAL+PqiPEepsgM4OqQZPZpbME5K/BT/tJjP6UNcYS4eQKxdT15Byy++
Na9HJ6XqR4gHZ0jF/1Pma2xVDYR1OATHhfJ/ncLEmB93zjcjnN7lIBqLzE732HzN
iu+Q1zcJ1adjtAjeq6YVmUvgM51c8CPBqq3+AczmpSltmKBOkrFF4O5JXdq+5d8Q
IzLl+QZiNIQeN711nnR1Ij9cq6Z1+Axbcy3SHEzR9GHChJ+3PYuugSAHDVH4Hj4+
jgKoHilKf/xQpyjyMHlTfZuBi3PR1pXQFgkgBXVjZkfWR0RUse0cj89V9T6CLz3v
M64ZaIZFPW6tn06Q1OGghGYf51b8nnesFK90DrEYDMnbGFaOR2MiSb4DeAGBzUz5
qRWt8YOX7X2OaibuvSq38JtW5wLnFlv9zmKK3LbNu8QTFCfkXfmUA1wEkfpdMrlj
B/B5ESDK1Dsr6Yb0ucy44EEoGtJ2ktclVp9SxDJcbpbwciOyKgyWeY89wgFrx24d
iNDL8T6FsbwdtirqktNCzaHxoiPLRGL3Q5fJZraU19n1iO7hYwUqIrX0uCoAipIg
Q5MPgQItsnE7kZ7C6IERA7C2za+M38+TLhBe5CZ3JV/RQA5EHezq59t23srINqcH
SEQrf5UV9O27XDFVl/ufyiQOvuMqsRyrvHc6QxYaOqYNH8hbDoazFnvuL6gO0xjj
8EvJ5rTZKYNNQPLE/ie4JCKEe+bWHeclnvrKytVJMmCDNgByH940UwDCqJijUk4A
tbiFklKxMMiW9DCKcYWiaxFklHV+DURhktvuoMpf374uMGvme87KWqDw0RWAGCCf
xXsdesT8pnPe+l+rQ3Ygx+33VwVxxiOPvEiegXtpZs/xICdeb28Bpwj8wNtCWEzW
LYB+fIFFetBvVnMOj0z0IBhy3DE1sunMT+4LXXqwIq6tE9aSG2fPG8rlrPIY1iCb
GwO1GPfmjRQQTC7ytR4W9Svbt5AaNMvoQ39n6ThBeQ+XjvArV9COK/ELSl5ALwhJ
K/SgD+uMxuB1jMMuWxIkC2+/H/mrd0QiRqxV5IGdZNRPGJZop6J97Xdi448xaYgQ
C5g0beNqZ6NpNgaRkm40LBYVPXsFFaT2YKvb6DMtystoKXyziOBNtn+l1gGkvocI
BtMYOqe2tpcOtmy8QwFt+LzRjHYqKwsQRRdrGf7jaIPvtcdYqYgzODvdqwWHK4/K
4Rrkr0OMxAj51kXR9Q7NwhDXDOUqdzkVP5evnhoC2YyOLsTgfaNE2U3hxsOZwlZI
/GBubJFIB1F/Zue6oyOOKkyLArrRJS7s0So6n/idIh80VztrxAgndmBk3+8zNhqI
3RJc+fcraAC9nPaHvr1GeTj/vTd4DjDUkolnskokpMj9onIU+W9AXPZJnTssm/He
V0szgfY5a20DvhxlQMR/IVJrZesN0reYMnB5pgOriwmL9M8iepbwNXO+YIsODCvY
yFTzQQ7aQd8WZvBjAWRfXVragKTiIccwc2Ts5cwXTh2rkoSERAhCWjcq5ooPWwBd
A7tfgc9SMSBoUJ9E9033J4dq6S5SEJgLcKr0JPNaEoUJ7vbXoCvYgXTKVeyaj+kV
SPUDT2fCuw4rRp3nRFyM4A==
`protect END_PROTECTED
