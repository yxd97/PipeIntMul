`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M94Rz15Gh4yyEgXvk1kKFDPIc54RkLYFAjyjMleirrIcB9S72VuMzf44uBOVbzgy
6NN+SKVHP7SrR7xgRoI7Iiu77OCtIGQh999T8JrAZbvBn8xj+fqhMNugMjSJFzUN
azQdO/BzwUnlcyga5l5aInmiNIH2Br4tqhabKO93xUjwcaNmP7b7soRrNu1gmQaO
J3bTBME+CStCSb5d02d+YwvyJzHIt6CeTIB06EOIEXLhJyIwkAEs8yz40xGR512J
Jqbj+l0Lax3vx7SBeZUzTTFgprZDrb8k4x9q8/Czkr4UflFe9Tence8/JdIvfxaK
JsYwVJrhK+xY02zHkLx5Z3JeiOkxs+oEBsxRDrWgg0ZmdvhTaLajZJCI6TPj1Ic6
Ptd9w2Ech3JEt/fzog1WMxaVO+lqLK/g3V3KfVijcPcPN19cvSVpKFr58IrRr+gx
NSOnpMaqfP/29ynP/V3gUhLJpt1NQ3zuWtRYG3ONUFd+M8Y5f3iFU+nQNWa85BjZ
JWDw94AZaOSR3jdmx5Yb4DJK/OHjhIsMiObUWCVDc3qcDL7r6oIJcjNHFex/4DKk
RT/KSwakLZ7wfpLUgAriyN1e5gJtrKUqSPdyD8WuKu0qH/XH4opIA0g6Cwt0C5LP
LdUoftgS+/FCt4ZNulTJyi2d4klvKf8ND8ILgUFVZKLX40u74aJhOwKcBgPXgXL+
`protect END_PROTECTED
