`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HMY5QILuErrnJz9EBddWu+EXYQG6Ik1gn0v0uK6c5MmprOzsTyG4i3BAGdzDlbhM
DGIQUHxz/VoTZ7iAS3O2mGhLjCPSFJmW7igccnZR2oS+H3gRRQTYwG//++G7RsZe
sWxifyTUnJ7QuxuRmnNd4N5ncG+X27vgdcYpZazIi7RQTyt+L1pAojVC3urslrWw
izndFQhCjBvqmIOcyXjFXk9xbS8dQvrMbx09a2bQ83iO9HJcleUF+7wp/CMuU0O/
K+AGynvH/nu0irfROZw6ewi1qRFwDorpQVw7QcE/nAOfrbUxeSxlCOv8Uq4INKKj
FUvKeMsLkQ6MCHZl+s8GSBEBCeUixFxx+poYMJ1xTnF2aj/hTlUREZboMDkZd9GU
/OCwYiPbGTPVeX+U3N6WQywsDGAil9sCTu6j4Hm1nHjIrdmftivaRDn2iKI1wHB2
E+tRmwb+DDy70TqwWeZrSYSzTBQWES76+Mp/+Vm2QPxlOcD808bjb/DlxOmhjlf9
/wgrZ5cRcFA8f0XtpdYs2s5Swizpdg1BMNEUDmOdPGSpV2g/Cjvp6Ef+7Tp8SB5P
yNPYhlnJGvWptrobJfcQra13y/UUPy8sEx8vIgDwGrf1sJHJ+9jR9/7RMnJI7MN8
jqQ7/RHIsFZCqVMNk9oOzZPiLHyImKNJwxivaxrlxUQsqHt25LfEDMBY3Aw0pCIb
BLGQxYj2SkQ4evOmjNUWS4fRpFYo16CrhVGDiawfdAGne7XHxxMbbnvPhKqecrTF
1MjMMiaN6LOOJDxF2SUWYvVLfTdgyBCVKKIt2DwHqP6AfsfYdTLN5xiCIF9/ZMa6
KB/nKDDNjmkcq4E7QzOKyahequm+MMEdbWiAxXYTvH6R7CMFU1NOm4Zk+3wcjf+p
D+s9IyVuzLkcgvrQYLaZlPiHShDGFp45T+yOxHvD6BzPydSC8116F3YyVCcyC7Gh
guOREV7vMhfkilP3t/k3b3Qbtq107ViVGtau92X6QbgxF21NV6fTh0P3we66I6Po
No5ntHqfJ2aZkfH6T8kxkG5XlGBt2QcuR5TsBcKet8U1f2Jr3P1ivx+s7e7DTdHb
vVusY7iykihRqDNvte9Dn3Dv+KWiHH4QtOgZktVXamvNEOi66sI0eFg6kfpxYjEB
gZ+mYs6gOpfUlryvnbxMZOp1j/5OSz5ATTg59pq70sC2NXv1cmNhNIKMAdYftiZx
KAIC5hHSpWmthKqaLSo3kT67t5HDWxxmKAa7jr70FfOVa8oDdODPh5oPsWlBLC7o
oCDYg0yxGH/tEFyIwEnJU0JdcM6lBEGInMMQFcfDNTqU5ZZxfrfQtJzKQg/8xf7e
julR31DVC/SlCX73N/bYxTYmq7UkvfpUbS7R8kJJ943DPd/K211vstrNc49vWhlq
uAShuHSbqR7rqddNm7jZZ8UCSv/rGLCJjtf2TzrOfTrUsAIN+YB7fIdwUVETMKlC
o/O9ilQiYoHYXBYoYhxGkYkua9Uv40tuS0kwIcjYHoms752o8XtI13R2z3j5jSWI
Nk7VZddoeJrHLTH0yz0Xg4m8+dwhyED9LI26KvYRcFioHkF1jJWGyZ1TBMPlzSvH
qJLvzUFLvSCYFR2TpsLr4ixW8FzguqgTAh6s/3fNCwDQmEDHe206ym5xpweqT5/D
fyTWiO9ttIulHW4SIDcztrl7VfulBojEFUjXCWvFvFwmPSkCv/0NFo2UD2blExgZ
ENBJuVmSMCxxJlsEnGtmMfhWK4jhZ8YAobjuj/KXi7rbiwxzGj3ArPoxM/oNvqir
TWtc+wq1qndZ8M+JCXH+bIeLMpbOU4u7FQ3SB8frQXQspgBeQKFf4O1DvREaC9+W
wO1NkkJhcn40iORAAbP9RK5hf6pM3BT/R7zBLglADbp4mc7TUZLXtWXVelnmdGev
IDVsMtJoiy4VJLVUgzoctjJKOT5mf7G2/oVVcXGxj7Dq7yKD6IX7GNEVVSHyR4XB
aIqe2Rqk/KQBt3wYFfi/QiFBOubaXkziS7rjp3AJpbl2q0hQeocxcTc+Ab3kLqMK
P7u4SUy+d6CfooRVzmosMtNywVugXZgnVapXGPtiIwANPld8jxirfVxHcJlwlsWu
cXgIHHtVxRggRuNvCBAY3cvtgBh45kvhPv/m03JMn0klqElVu+bTS5xHXTsmlU7s
nKetnxQYjb225w8uHtiWBHtYIvueahBOSVqvkuxyZwq6A1ny9fay2Jf7MrXkw538
uT3w1F5rRdTXtnZ1OkduyXMqSN7PW7WnzzIu3Jjs/gFVh0Md8q22hGiWpY6ddoT0
iQQjTpUXFert/uyO5I/iT+s4MJLSdLEaFEDWPRTyZ2vn74iNezw9+g37Lg0QLD87
EzVUANGDl1oQmShdSKMiFFAeiAuoQy0ixo40PJgVWR2qw5Swpr7n+D4BmeQVwViK
BZe8K0dWComXc+Wua0K3Hl7sb1+wlWivDaUpxd92BBfM+t9JCE8Ao361i/kAV+/+
kX8lMvPWjG1f/E7a7ib5oEbb95WQsaeAQKYoKLyX5XKjir8MQholrMLcKV6r9DOd
79md88qkSjUezm2FhBK7joy6LZVzSd94fx0KQ8wcJwqypqgLgA3shqmmhqdfeaeb
Iq9wX0lVjFrSB2dg2kvF3nUbNApG01EmkFCVTUe0qiSL/DH+/F9YQ2WxKgUEz3g5
HNa20iPZ63kWQXZbZpIJJ7QiNGxy97r9iRSqzVdMP0jt1rY+xN3M9ZPax0pxgfyK
COyuIaBKA4r3ccGNpDW4ZbFneblZK6gw9h9K5xnmW89BaCnEFohoSpDzUQR+629g
kxUyHQvLNwjwLmMdxPBzXuVtQM1vpBTY+1BIk39e6kROr07OinnBfU4VdrBxh2Sn
XzCMxvR4C/6yXGKZRMikEfxL2moc+O9dT2mH1xbhTH9NCqEgIhyvztwUGW0MpHgv
jyH7vAvZcgLr77Phv3+6xhjabHCXawVu7Z8WXIi7eAIZc+diKPAoDIXO3oEFkfs6
mtZ1QJgaQ9kj1jo2mDpYvxTZiLh5ErzMJES40n5rbVpqo4CWDk7DJTCR/Bwh1DSS
glbOFw7hqk71EbH0RGRsxgS0TgJhvj3ezr4lh1N0L86rAbZduBRZj6D5sYOF95qV
zwYPPDnJkf8Fn2xJbXOAf9FGHOFpv9qFl/kf2VryfddJZjBCeffponJ+3NbOgfVR
wcY/gfSMWAhh/2QCDtrIuBfjoX3EhPw+ug36vnQhcvpwc1mTE6SuqgYLuw8c08gz
UomgwgAVIpXppUL81rj9Kr/5lFU0aEEy/0s804BpAbXYThXeWIhC8p6l34A60KW3
ynUY2fKGX3rOi/xn26/gtSXXSBWRO9+FnWNeqLJ+ZmoEN9o+7rtOlPkydSS2ZGLs
HbTzwH8xsjNb7Ce1YRndKWQg8sZtT8BFOo1wQgbqKsqjXLOeDTh6QLbdXYxyHzLk
WzKI5+hA+d2yaqww5Qgh46gs8NvTtLNDPJe8vv4beOZi3EaxQTIfPWafO9DhhWWf
8aVSIH6qN2Fc1Gk9YzDyUHHysORRRcMneU3iBMjOtzO76NNM+gb5N9N5xiOjDJun
uRH4Jecpek+jUKIXfPOpbjA2InrQAQC0ZPjB8IDirApYiOi1aCa4Fy7JIMxDJElZ
CAGR+MkXb9cTxHK/R6i87giW88bPZ/nVid+bwjVm/Y/xoym7zLOL0KId0cCTJDJP
AbcyAKDi9xoGTNpspXNBIfbVyNuJ/nR+H8c2qgTm/ooBEFun2+wtgczBVdBYWIRr
7NXD+OcX/WBvZjSsEH58tcbyTsMkayR6oUQoFpDrS/c3T8wq3V0la8HDf5Xg2acr
mCyndtqL7L0530NpVHCD82TBoYown4/2gjQJUTIMuJPuxmfMxNeLLbnTNFZTvxY/
RH7KGDljAS7yUfvSnxhxjju8XYJ50Fa9RvqbwEAH/W78/doqp5xZRV5hgLFURqBg
UAr456sPQYUciGA2kAfDe12WhlI2nuLkEM43o2fhU5apVRsxIXTU5LGYNmitbqPK
+4V9vWnKNcF7GkKxkpuZDdGDYgrS04brFZb2aJrpETwrtCBafuCH792bSf8LHCv6
BbEDlOjHgDJl9y8m1dLS7q8VoxDmR0g/f8glApS1+uedk18qKE7sNs9SoSI/pTIN
kh0GMEWbM7jPBDFN6rHKEm41AFYh2sSdF3w4LuCHbG3QnrqAw15OXFEr6QgIYO3+
jdvb8vcTGb+xM2sLTy5j2M7KQgKL8WVPtY/81uezVfOTb65J12L4qRdU6Ktim4x0
apCLRWTk9+9vy3FHORflUoDBD7l7mCuq20NpNKYI10KC0FErRJoMnoO3/UIBhHP9
KMH9YPCJElDPz+DpkbL9r0kf/0nTbQzAeRzSi9euvn/b6sqmQhPwRmx95WREomcf
EKqz6FI7Ubsuy5zwsqtRUbkthRbV/+heiJa0FS+55XgU1KN6MMkVEeVyy82xRHle
A+uEAPwdwpubUJpcfLQctQVnmoHXZI8dDJM9i6LK21hlGwQvk+hLWUBsGQbDNLxT
vvhzZrExQ4eNsr4Sdu39rJlOxck6sHSiVCZGIFWLr5HlulKb4DI2JCKMN1Zq56OJ
Urw1xYEv1JLptCLEuZr5VgaRSuwEBOSDhNj1m7Juceu9dw/R7jBm6YKNHN182iCv
TmzAHYHAaNqhTh/rWJxdsmwhA8/ROH9QzwK8oFjptE1l/sSqowXmW64EDBLs1iJA
bPKeFsJTI5U16tyavu+UOWKfKb17QHOCkd5WZl2bQVjYp/5ithCmQgyrc1S6bSan
ON9vKcfH4nWG32hipo9qhcGiYjWLxwS9LStatPXVxU2CduTq8OXuV9DG4ien9bPw
sm6Vh3kGQYFPDmOwLpUYNBY3DewHRieLcaNw1PLko+4CXsiR44NXOgy7e0s/pN4q
5AEbxBTy7pt6EAZ+Cug1G18PjUx4r80oka3KQgKc77oprr+7kvKYjN8W3ChLLvGt
B0byKwuJQKZF+UiOkvWy8EOAhJ8kosJm8cNkmL32pB4MvD64eIMI+bg/+WIywlqC
BuE4KUP+c4sto8Nh4/Ux3KhB3YAGbi1clPxLOVT3TtLSpTJr+jphPu3/Q7DvWRx4
AdujVUWjIf709namim6BYZwLd+OyzzspJMwU63qSUFXzxL8aiH36QDTzEGS79221
bcrigGFnzwg02xDa8p1MqYI/dRewooXoxcqsu5v3JyP5WXRTXZANqSSVM2yXeJc7
0ZhnMfMM6dwcPLGwsKnwXsis+kxpV9XO5fYGAyBoBKFds1aBVQ0GbKTFS5Azd5qH
mSE2O0euOk87NB99CTBD6O6SxatS9vZt8LOz2yTY/JHsODRgja99dyT3MV145OF4
JAStEyukqglrcZ/wpMbZ+BpVQukzFW5Ms4avyXygktM8UiSPEivCffTqpv5cIXKc
Xr3VViEHLm8QrgixreyzHwcYb3Dyur+bnfJqoOYqBadFCR7GHtBvRwUBwZ7tSJ1U
EeW19kd0QrmVAGViP+ymdxoMu0qCbpIGLWOjNGSstmJOvx+xSTyMNA7V7/pZ7aJN
zPLpYAhb3cqtRdKv6y6xDyf68Lue37z8QOUF5DVJDufLOzcackNGfoB7+dFZ09sK
Qkmcin8nE5Ij93xpU2v+BKUvsfJBJT0/o+DiPtj72W+fnlXOxaQHn2qhU96nabvE
F9JFtvGs8dO3Mp2X7au8+w/Jq6oSnmwvPLwD16kXZgJ7CSnnytynw1JFl+csOZsw
3UuDtNH/ZCoCq/LBw9RkZSNHXzbrOGKp0Mw5bmdoWANgY/8E7e+XI/LfkHvsmyvj
dgd0UzEruwYeavsLFMzKKwYTVTVYeEsJsC5Pv6tGCOwmo5kUdAPlew8qTG0lC8Ko
4oH2P0ttq/N1OvLW2TEnZ+gG9yIdk9lWurIseZgN3rk+C9AM8JHY/0cV//S0GuNj
6bPHT/pfuUoE8oTgdDiqro2EuUiCTEHLhzHDE23fyUPw1Cv6nOLaC8eMF+tu3TAB
3XbwqnPyg+FU3OR9iNldcOMDtQ4cjIbgw8QsrxRr2ii/O6yKCJiV4DQKL0ccp9Ho
NcmMRYw63wam8NYkwCQb5+XQslbOfxx2g8+GE8ugkudZlUeQagp3seimRBMsywoN
vBG5VooXhq5NhJ8Al9HBr8AqYmD/bQj3zIPtu1Wu9DEUyYKKVjUJ0p0xwTlWDEjD
wUg7ozp3BZicDP+N6pZjrMkoovwRoD0Xwy/pn30hhkHpXOO+5Nsfunxc+guO291U
ZvAs43TMwRYXaxiFy99/y+cKRRVhZ+sle4g4VfhALmjH1lO65o+GhWJwKbVA25NG
pKTl9w26aFGLeB04/HBM/I/twRLLZVEGyAaY0CB4sEl5mwCZPwtU5WR+7E37UJFX
wnEQBixtpe1kIE/xIVX3hf0ZhlKUjXOpyzIS0l7PL0gp43PysU1X9yahrmMhmuA2
z+nRR9TyNX26S+pXkwguhbeyyEmWiig/DF0KUeI1geiYXY2kwu09cqZM7vH8CiIc
ckybiYuLkTCnSUt4doSYzXlvOpvd+7FxnnAOne5aDidhGrr8P9VKnl1gNPZRDc42
KNBDSAai2Y6Xn4a1DcGwzdDAWm9jqxAk8hAJBBhG8MahLmz7zcEY4vq2iuoq9LDJ
/CUiioIhNZ+aNqrxGGSrLRzdapMXsR1YlSKPXRtPfJmBgU4ocTizkMU+PWq18EsO
1dfOxiys3i6B5ofFdYhSPNpQG4jn3619H8rY/AhvMsjelpgBOD7qWGNM6edcyhHT
eh3tyk91nqZLIdkjrsS+epyPlSL23ADsP2H/9b4SjxjufnqlRWz9INTCdCjSNgLY
GT4lKjAoYTeqX54iWa9PbjZF8XedjTt/Px0UQ9Q7MEapgIN1V7b9Dz6SpVJTtWBT
dLM+LjkSPSomgUiC6RWH58kZLAEU33gBWkAE9yxNZVXA8np19O9t+ipqbZZEZrSH
K39y7IasvcnLzTh3n0c5X9GovLFuzDOdwRfSZHL1FchXlAfS9McV6ULic1deiM4a
G0mWNkPI7dR2xS3vUsiiUvOPr0TKS4eI+YIh3abXKak8majPOhbvy6QagQ9rdan9
+uqJoGmi73x9oDyU2KYi7bJnFuztZ5mVGgkJ29M6B0vXfVm0ai/am1Um8m5G2H4D
ojEjO2s9rXKz58+lYp5o0Cs7IXsFE7Zbl3Fh6gV+VbVlWTVK1hbuYNLw96RarPJ5
00TtrpqsyO96uhglmJL6E/zmCXOetb2GHOYljgl6QlGDSiJApeQVGvX0jJYLLIL8
Un/MJTpHsE8k4hZgN+VeUmMlQDM2zwu84D0V2rHzqRaWciilO3JzhoqYFg7Zc/9r
lpFDBirvWdbRnD+T1n9OJq2F+L+6gcrHkJ3YpNC4qNHRsOai2Swyytx0FGfHh3aM
WZPi14RR1vQo3P70EX0me1ndwgUy4jhGjQ8uRnXkuIaU3/AWGpSmjGzI4QFlDOHF
kXcywSPQppraqPpU/PJ0fUqRQ3gf3XRMFfp1qKnPugciI2pnpfhoyOTYOOYu9e9p
17eWflRne07x+7pLviU6NBne3yDR+BF4dzA2ss6bXG4=
`protect END_PROTECTED
