`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SvO3rXFlekPnYL3qeoCFcLMGLrv7dN5OR0u5dU5mHOqsWpyZiiZDo8QtO0s83X52
PPXWCbfojNoR7axp6CC9xa3yasSiS0USlL58WKGtK3GFmhob0LTrPpjOlK9OBUpd
vUFE3kIDZY/q62TPu69Lj1Z6+xq6PYCUwti5ej98sF21YYLuzHOBYn3KDTRNIE3p
BQ7YsZs7xMEHI/j7wxzx+8IHdfy9oU6/jQww2X+302OJYnyb/qRk9tV2/Sc+h+QC
Hs4gZizxK723NUO1mkES9dONaYW5s+t47imLncM1hVMt4A/iWkFqU4FNM4hlnXtR
vIGN9XPX7R2SsYYP0CHtnp6baUXJwJvW3jsV/ETqi48=
`protect END_PROTECTED
