`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1YpPMPQld5r/zOmTJI7sZzsorDxJcIOYQ0Eq5ZOuNvDQta7g0Gb6d7CUTgWxJQ1Z
vX0vyo33MFSE5QRBrkpy3I8WMa49iIwWgwLh0m6BNZmnK5BtuI73VUqsfCXkTnDy
p6ui0QQLRbnNJtrygY9I1s0NuQcuvk60n3wuPf+jKcj3MXAkAc0ZPzHtfGYFmyf6
yeB/wp3yQ1gGCf1ItbflPsw5vKFV5vh59ivP7orwilvxKujX4GMqkiBgATHndWPf
ai0ZhcxvNDYWLI/AnDK94A==
`protect END_PROTECTED
