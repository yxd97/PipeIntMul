`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Mts+/EXozRD2gpPJHQPUQ6eul+HZw0ndSqgS91rKIsJvpk1QhzgVMYpxbA7voxhJ
yxImVJDyqbMro2zbuhyz3pxtncIfRMZDLu6d+P+6ZE3diRl4k9uEpU+Ec9kYOguX
0dzMQNLQ9enFDvN+OJoSuxJzaEhQNBmhointPiwBO4A7qAmBkh91slNTXivZLqKS
Gsac6FlxjBE4w1b1oMTwHqzt8XxVOI/+8QtPUzQ+4hsQtEpYO9yPbP50AIVc97dN
49yIowZqBDlv/+Ff1hVehv8vnJxGhkZpIPCkv1+W0lVzX1zht9ZfHRDLR9nObca0
iTxmTqR3s1aMTLgxvGlVEakMaDTl8Zjwdvdzu8o+MTO3aQ5QhYrViUWTad9lXEc5
OJDGW+yItydLKjROozawFKgG9W9khEJ3p3LmPSx6xVkyK7UBOv/iV4zpt/bdbhXu
qukI+80cmkf/iGAK2GGPZ9oAVn4M5HSHt1GWVnHVQDQ=
`protect END_PROTECTED
