`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+0DNabLiricWXLavOOUQ8eVoIumtZnjIS1KJ2EUK88fzFMnpafPf3rtsKy2bCu9J
h99s58ZHnWtf+6ctzFWWfZSHFRQizX+dQNV+FTfPnBaco/B3x+w4hgGf1+xtVy97
cumjs6S4zG8KWP47sOTE2g1KrBvnC8LAInTYF0Ulbz5gCp3R883aykqEovZmjDNi
2OYGgEL9vxh5RwZRAeYA8tc/CHw0bN7s68kYuskv0U76cU3bTaxlbcGNEbMqozmc
OLhgMPhRKO+zrimYUL6M8atBX2MP9AJCJfxyINGQVsHq7vP2/+Ur04BI/vk/4FC4
hrtGLWVrAwbXqchY8v6ABgi4tGarUE3g58mv2AyseZz2ntEvySpLFQ9FSoLrur+e
UOfq81kpkOA0KW/ckU7ZscgFAT/N1jmytXI0aq3ORhqNGCyedcigL2UGoOCdFlRk
aJ7dvIBWPwV7bHL27LpRCGyscySvSA8yndWFDpfbbd2pQKuMldsw1GnE1sx/DPzj
HGiMrK70FXBbgt3+90kMNfqJgkH46TaHi1OAIFSBKZfHpp9y8sVda2Qben3c1U86
B07SZW3T/WaiU6fXMsghyhpXnJej1gdTHC0ouc2WV6I8vNfRHlrXBpwGai29rLd+
ruYzDiquEgddVQ76baRyCWHmzlvcxQJjupwcV2Qkee4QzFTXVfvUFF6Vi38lgBAt
pgwu/AxNe3fHwLRD8nItKPmEuTYpYdwYkjxwstMeaK8bGK4slSLEz7pHzUYNSL6b
+Ip6OJ9S7LJjlWVNtEHc2nro8iJrUuggwFWAdVRJWOJT4t80d9hEJ0UjSiv5qslO
QTa7E92kSLWOn0e08nLqRUT0cfXrji8Fyvy3oi50t8QGAvHEhoOETuAO6C5i3AnF
o6rBzv9vIJwFmT2fTKxPym5kD9m1c1BVLTH74QZsGcLZ2xzv1gd7LsV5n4tJShT4
umdK6f6I8VOFabXkPrav11m7+mENSdxrD3j4ruovfeb1ZUhTkgWEYuMQjSBJVgM3
IoAGWB9uiiq5wmpGxYTf3aNQCJiwieBgwlVx4X/v7knX+yFuchDLL2RRVfQL1ggZ
gf/SH5T5RD5xABi3zIhsnioLwQNX/mFGNXruCxu1QPMpuKILFMzMEKB6Ei5YDabN
CycaYFaXyYh1cV9eZbDsFrs6h6NkUyDevHzZAZwvIQVdwpXJF+WC12uVxTL/wURx
0bfL+T09D/xXzXRpZ2Xc+HwOmAqNHgaiw44yDvDzFInFE+mRtWLpGRcVmpc8bpw/
iGZG+RrfUVD3cZS5abR2yT6RKu9R9jsLBQ6tdGrfH13zWLDuSmP1do7c2/BCaxfF
xBiE5c5u50dlWapRT7Xdlyi46o/bAOCtf2N9Nf+K3Jili9K17eqYHUFNLqAwbhKm
EoqI9AFu0ZXv3/GgjJC19UwTzV5xBJ0XlXmtXlexXYoQW1gznlGro1TlnvamjNAz
8sIDTRviVu7G7/1TSj7fYVmdZ65oyWjOAe5iKzIyOKMCq2vqWF2rMN2HrfvUFjrf
rR6BC2ZTEYZY+e2Iuh6bjs5IA9b3uvvVX9iGJl22j66dY5H+v2b+ZsPi7y0yuqMX
heVbelxYYFCIj/u0NPcfWntaD3DIRf1RvSTW6uhWnlH1rnbMMA69dkaU3TUoyzwB
3EVIz23ozEAinXZz+8AiYxTG3APGcCwBIiNVdFeu9d/9NooKb2nUmjgGc3YKhuCx
XEUVhjLgm3WT6mSrsTxuLFP/UPu6lROBMWhUgE4xg2bQamj9JlTo5BswmTlyNG9C
Vm+WazI2Ss8XSp6eCLFohTcxCeKpJ5hVL2WUImySRRTnwkQdASsuEwza+R7hwDHA
bBVCTHjf7GzfKhLI4vGf00l8igGmK2oEVNEiEJ6GohoHh2GqV+P8VO6sRKroNB1X
9qE8D3PXfIsirEoSjSkrRX+USRz+2PUBVNs36cQYe1QritqimctKFc8V3aT/sNtu
96lDfyX16vSlzYbq5iTROgPMIip4oePDAP6IaP9qEL10OehiqAFSWbw4YqaUDAGo
xa72ALqyJO6e7k+9vlEJ3LOg1+Z7ApHhMhNAfgz7/9UFqdKqI7MkCbVMGVuPvKFO
yS3H9NGh3D1p9oGV+Fc9TF9+8gPeRHfLtHG7Tmtx02cIfZCzhUb1gc4UrF5+CH7G
0waQKVRCT0bhFwJULHS5J6xgjQQv0dOKpVWBbBA/YZJgcs5rmdrVxUKYkDayfjF2
B8r1vlmFnZzD2sjv+KLc6q8PDLvxI3q+p9f3X9LLMKt6EVGY8RSCZvMz9ouaXN58
OGS+ujbuvDz+qfPF1pHzdRYtGsrpZO2yWPaht7W5qcNJ+LGsJlaB/vZ1hJ8EB/sS
VXax8RhbiJhKRCX9bcW959uww8AU2gylF0zjhgIf2E9hxgPI+CRFeQN95AlRzww7
8zANpYD9pJBCWQsjr5oY1Yc6aVvEe+Xnha4AIa7gTzmomEoq29KRJ8OL768B5yRu
JiwzfWPpbWAfn4GVls8rrPXPeU3cGA7d/qqq+GDeRRkvVHs+9IB/ISlQhbS/hyfd
inZFovvVc8SpNW3jE2LcAlW69WioBKt7ajPo83uXO1igLN4Ap5YUVApzeyEp5iQB
bqkybDlVk0n2dlr/2JMgvjDjlBMm3ETUGvoOOKgvcgIM2mr1D8ZE+WIvsvE9XXqP
sUebZcrGYLPx9XI+NOo6dqg3RU15Kh/6Mud5vKJ2DPYXXUBqmBwibBrwIO2H4nvG
hQYYJl9X7NGBP2LvTlTFC/UVCRoWcFVFLwyXcr4gxvekCFh5EK0C8S8MSKPeCIJt
2/6yJpvXAGuHN3t/d2ddT9eLDDms7iNUmBkXXJ0UgWtJbM/BwNX2Y5t3Xckov2nv
oGj8CKwxgUA5VdoKmkjXf12NuJ8BJdbfB19rAvPWUSYiHBzQyzhr1hcVLUsZ2IKY
Un7HuPSnjTwP13DTUpCO96r/gq/aZWzJg0pIQA2C8uIdY6awLEZXXfurULXclAHr
UpWVnYAo+IOqT5rQyzz2LoAEvPamEnDrILAoaumgqPMTpOkOGEsuPN+3eHlwjftt
yDNzylxejixFJ89RKBpRsDzjIPelCfdniVHfzvwzOphmMWNr1HbA7mOFhvTqrYDo
xjM6Q1jNpz1kISxJqB1yrsEqtvnnfO/On4aBcM98LTIzYH3Aq8k3Se2kXHvSv65e
uzRmjgplZcQ78C/WkPtnog75YGocCyjytfWD+5BGFMQcPUGWB63tURJhlhGrHjSD
ZwlSmn7gpM92d0Vbk/2RiN8oV5OBPOwQLuPwpdckCKUfFfjR5HVPCCZyOXywZzkd
rQP/4o32n14ZYLyPnx3iroRMbwd0qXWg7Oxc3KhWnsTLN5wSlUThULj2E1br8w7f
x+rZ3VgDETdAuxtayES5ik1tFOkS1kwW5qF5pj5KbnQ1Lt+sEnFE2Zw1MoY7jmCj
BXliMG6fytqurm/CrLTQuVkyXXKoPXTC/fp1ycUmhNShtoKabVkwxKwtUXayUpRe
siQVvyws+X5jP78NFgSW1AAwQH6GXlWWEw3iqoex5MhecLAxqr/t/uebmOvdZ9Vt
w5/tVreX/DAYw/FIjNDeLPIGDE0iUP0xUp1bl6zsjd+3CDtTAGdSHY103ozktdH1
zh2vZZHJSu1KwG7AOfMFRyK21Dph8QhoVilkPIjsvlBzMQ97yTshBGw2JGz3tlRo
l94ZrmRj7hu2pTu2G91kWaEvb7yw7Jc5eYYv96mnumL5nQAIamF0Gv0t46oa8Tgg
JkzI3kaISTmGO2ssIfchi9vMaKZADaM3lOZqfcoIZqBSpA/LReaHs46s3udwAd90
XQoGa9bLAqMOc7wShq4CpNft0f/foLm6wCVh4CX9NMu5dMg0mLLI4Os35pkEjLU3
UrokdUk1E6u4LndIdm+P8rv1NNZPIkNV1qb1Ha7sJlcsqEtq7AM/VLKQOApI/nrB
FtLgfZ8FaoiJnmD8z3dm7ss2m07A8gatwBaFkXwDV9hZnDS2iMxUbvQK0FqjG/M9
7OrA2mF7hFPn6iTU8dwO3KOrzE2VZS/kgAqlHVtEIu8n0zYqifbWaIbYFzUP/Ka5
YP5n+WLjMRMu9PVGhXS8qWhAtpeZigAZbvFxz6Ktn0hGKFOJCF2l6dcrpwyVtoHj
24/qpE1E7WvNGdvQbUgSbd3Nv2qiuu1pwUrFxXGcQVXGtYUPXjwR9t6oi4i72+5e
ElH/Amx+bQjB+PhMqNhFtd2bstRgnTfuxL2z9s475kCS2lAqoHBod4X27jWYhsER
pkmkv/enEFAKcwG12fN44c/HEtZXXHV+vEOTOfIMyUp8c803y5p73KrH65FvsRhN
IQkEoRqPeD0ASqZwzQt5UbiXb0YXXsD4cbn+HCLkss2tuJtGRhkFZmRmpBO4kDDn
FmG4yQWQ9E3FsY6AbL4ee2M2kHfDO0DstyuTYme+wj1RUs11jJHKLsipJrPokgAm
D0pJlMBCKC6An9kMlkVqx6EMFqMnAGytdMWv40CiAspGCpc1uVdhXEVcuYKG6CYA
InFklUkiMpULoJPxpsjLe3QWJsRIh4jMKDkuERKOyJuGME7KLzcRfarOIYSyN21y
nTkybW5DfHluQvBuYS7q5J+ZdThz0aT55JcSrJ+NoHfSio4uayK2Vg733omeYxOC
rXmxjR60fnYikP7uS4Boafb9uc/i2VxwKw4NdYL3xxQ=
`protect END_PROTECTED
