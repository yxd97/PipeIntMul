`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7ZetbLOP5Uzzxs2MTrCP7EgKKX7KPeIgAPRj83SY4ixpnh9ocbzgsMnLVo0BEzrP
9gnPc2FxAIcu/yPXJto1NIYF96JzCOv7RMC4ptuuVH6j9ZWptERK6agwAb3kl/cJ
PwFrnpH44W883PyiTKwdYJAgjg5vzco1LnsSTu9RF05yrqi/ty2/MFG/u+wHSR8h
kSS91HvkCDHAs+7mArF3V+LKRnwDlTbnhP1ExBrIfJ2QXHSwhvZMCn2I+dSg7TTc
rb+EErvBUuqiRAZa57gWy4NTrOuLblJfn9P/B63S0X3VT52Na3kX/dZ2Ski8dxO+
DPj9oZDAaO2PkhMiM02zzN/0Htjnbl7cpY7NSzps5nyeMyVcM+PujKLuo8nfTnfG
MC5yfsXkxWWcUOYE2SoVNsdonoX0Mt1yfCwmLqnvLNiB8Du8GpUyCRNGmvhRc0Fm
rgprq2HBzAomkx2ry3WTHlLyZfUbWOaLAG+4QKCdyABOfoi515whRvAGpZkd5y8Q
bjxpUCfCtfgbGQVBEPBQLlRTzW7bJQr0O5Sg4LiDcFl7q3IH6JmNGUrA3GL7VH/z
QioDMGNMtMUYuHHwepbtDt4TdsMFUr6ifpc2g2EKAjlImCm0FARXG2H7E8NAn+BX
Gjzd2EHxZ3JAS5G6Rc1lZtL6/YNy+Lo+mtc7wO+NH2B3p03LquxebNGhdTnVDBD6
ljyI8WolexrRp0klTxzTNeHpagIA1h4FU2HrwaRHr1WtSX7PaCUYdKfjpGoM7NFE
9MjrduLjvj+xexhTsBzMC2J8gcpetwM+A/qHdTpOmXoPI+Q09LoiZ8G4niH27ktT
FKQZSDuvpoLIwHsl/UTV3AmsmaaIV805GMIixdkjKZgx+kHqARcjTS9MmsVVBiKN
t+EUJXkjATvyA6zufuVnXWCiUFac4joCGNNdcpz6BDVtQgXQJJJn7BD9J+krFlhp
OUrbEBEAH08BlDAy15aOasfL52YcNOAEXpc9tC6OxqjUHEMEcLEMa6YOQYweL0RJ
JeTjvWoAwcqv3Qa3uw7S4qWKugjUgPUBqeHZYqzaAtJtphVoKdYxao2d/QDumjdG
oAKIIQG32oQyCA6K2gAmjuNBGOuPDCjLVhjaBvqUeL31NsRVoYBH27e7yYx9n9Ap
ENSC1irT6Mq0ooUCdpcOCzvYoaWiIjpNKnTaizSHqodLCuAqBaLuclj0OzLPgMHb
nJGD+g3IhL/iDvDdgt7GQfUun9kLg126SpCehDfk+e2Xm6C78xvCE2UICxglONt1
ftcUf5TBpHgVhjO5riChjJxyRIUvizkFJmsMknZDhDF7AyLyRbgpgDrLI64oxUPj
gji2lO3fdMPfo5qO0hZgtA==
`protect END_PROTECTED
