`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kd3C3iVD/G6bd/ocboebM95xrOOosQyCw5TKBuLl5X/woO/PMNs04IMEdysz+8J8
mTR/BRiLX1d6PYbgsTsW+f61utty7X7hnoNfKSMQ8ey6XFAHBVBBnJudftOarwaX
FK9xTUwIvJpJnI9eUSxvZLuRVqv5b2URMQJpWPTykQHSF1+pmsv01e4nE5xEx7IS
pWSpLufhwKeVQEAB379e2pbE06TKu622FAbejosxlmEWCs+QqkAyCW1u1iEySlu5
qBZERN3kLeDo5D2u84r7IY3ZO6pLuAKO704b5Ka5KIk=
`protect END_PROTECTED
