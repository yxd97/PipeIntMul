`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccnZ5nZKN1ERIdWv19QtYoJzdtmfwg8Lzg5xel3QWCVpYNZz0EzH4EUU/AOFcEOf
dk3XxUiCdKzXAfv4vLXUGPWlDLJ+CEG/SG/PjQ+AesPAy81PxtvlIbW3CQCGl9NH
rb/igkdcMxxS0eLtM7YVcWpG8V/clqG5GDCCMU1QzLgZR/mF9ZX0KFTXQiVEfbJF
K7oZ7YQ5ho8/QxdlJhSDqt2LAo0wOvBuevfyhIhx7+44WaelNboWM2AheoL7+VMO
jRpMPuLh1YbAOhVaYt11eJfdXYjplZOIVXqqUBSORWyyZ2zw8V/dol/TrRqLlu3U
NAKvsTstcpcNrJJqLFX7rg==
`protect END_PROTECTED
