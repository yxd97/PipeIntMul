`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d0B0G/vH4i9IN2jnK0/VRJ1RsUDdC2KXDNrea0djvvGc+XFVwcEENuVf7Msbwga9
AaY/S5RzntaHTTCCok1DbfnptTWyRqGtODymay1u6BbzM5ffbRS0XXgqr9uBgrUx
uEwjHPStXu+YgN51QeE+RvQmNHRWo7WCDnZVP8YEUGRKIffPRuvSIBuREf9hi6Vi
UiSwkmp3FXC6ImWEuDnlYZ6j+cn5SOfzG3GEPTPTvkozxdToaSmo/u1Y4blc+1Yv
LoHVwjbpJEJkZdWBsCiJPtGpVEF/x/nqWjEdYDzwML1skfy5Z13KQcJxD7O4spGL
nFfvJRPeHRuu6LJgkjlnbKPadur+pt+GW0QqsNF4g75pGVSmnIOuUCrOw6r+3J7Y
FHH/sTQa6VS9tZJSCCN2Ag==
`protect END_PROTECTED
