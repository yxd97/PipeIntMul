`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UJdnr0OmtHAjUtlGhsp7vmzJHhZfAEqMKTmrd4fJGVsLW+gSoaMBnCJ4KVxOJ9Cj
kuXblksa/onfT4gGlheRTaiKKsymmiJ/XFJPtN+HcNNEkpro9Zps9bIBKX6TWEHw
9zUQn2q0vKa7zfxj4xR8bo6qHS+BDprb2FDVQ4wMSUNTQH359FnTF7Pzs23KAwE0
DipTSHuIk7Fqkfqs9bhsXUleN6RjOeINqcpVmkXkd+PPEMypLdzq6CRcecgdyp8P
94tUQbelKUHfCoFwx8Z2EVCFxhOppP7PBMyFWj9Nd+u0AOawj+p+EHqQvssqnx1N
4XL+uw73Pg+fiN9mHr5yPZTkDYfjeDAuXEk3LjSgS2yZWPQ2uboSuYv+rCDlBke3
8fJoS/Nhsd6k68W2AQmujTxOZDUF4YMQ/W9Mdrj8oWZl9fp3SvjlF0S6oHFM3hA4
T9qmt6sUq948CGHiEi1nItEnO8ulMirtM2S36aRGzWfij6Blo6DJpKrp/rGLG2pq
gFOK3WiTvojlvwIWSOFsn4RHCmgiEr8XJNPTbTTZubqlBDEhEYvTL3AZa8lGbY2b
uWcJQceIjnUjRlM10TkXSkjR+mGgDY6/W1HbDn9vTKder5AqmGTLAAHHFn3N6cmq
7IQUspmD0DjUeb3z9DVgZ4vzuW+3l0/sBNCdK3pLiSPDqgNepKi1zZEO3Ey2hgKa
i90GRcEPEjE5QjqumBi70aI3qdZ0Dio5UkSrIvmeJfjJID3GbYQ0JTmTZWBf4QSr
mMtItWGfotLOhYZnBEjdXx1yedqjL+93qhyh8MwMSN3huBkuwRkDaCeFRoxrC7jQ
xXRgs5y35TajhRtmXsJH8wrpxMkPXbCHeyAinrWIIsYrpTc3mmiNgdVz0cKhwYC0
HIt3htQ81IAfqr1Yn/+EdlW+xsNaL5O6sotsnGAXy554Z9U8l6J01wpa9ezwqgSt
c7EbmnX2QSC/vRcEhl7FtvjkNhZUF4832UthcuahyJrNNrDR8fn2cjkXAbV8bWYE
xijpB0V9ihu1pcJjqgwQvNlH8j7MqEduEJmYablOIPEK/8LaeCHPuOLog8HIMpoD
9oQ0HXs6+Zz/pwuZTkI1wfs09oI0d8SJZzHutkqHs2TGyCArC6Rk0g7nuOsGvI+T
Zc3OHmkUiiCZK9UcuQn8wydQzqjCoU6PPAfrSVqb3P4GR2omIITkF2jNEpn7IqIi
B8CrmD49vqJuAI3hUVjX+aMXuJKUS9QoloIHkLKmzA4qYV8MKSAVJuqZcoS9/3Hu
hXEHeE2D8lgEFoEnVFUUnwwkpoYlLNemi1TpOhjIONomZU3Odkpi4oCv31YhaNVd
BrczRVYzSX6Zs5Z2vgHBvNRpqD9gOOwxD4f7KsseXH9IZ3iyXtxhAXPT+cBYCEKw
VhFBsdpvNizAap7WNLHisLkPyawnUGRbITy+HTw+vmK+XFKrkjabs9tiugABoq/D
FFNDO+WcDiPzKVn6t0Pv74ZFwMNuapJFBRIR8QlFT6xpBX5flp7kg+Mm9sRyL2DL
PR4mc1SMszlO1+YsV2vCJ4TjPsfTQ4DjxB6kKtjL5ob8/6JcVsVoLzKq83PfdlOb
7Sw+nKDdUlt3KQLQ3EG9lj3kn8otwIeqrt5Xc+cl4xYMMWk8WQDoIxo5+YcbQiIw
uB8L/RjDlfzNJ37Gwxa32amxdtoyCIpV/b9wMIJQ0pjftlTwhfuI7j6rGoWyjKmU
+YpMk/8KJKAl8bumP1hwmjIK7q1bZNeiZcqD7vxmFFp9jyNL139yfyqdnPL1gBQH
7rrp4LlQr7T+fqMFlg13RsiVO+KEAIedElfrYLzJjbF6W9Mcu29jip3rThWzvw8v
UFS7BtfK3EY+prmqJ4wQF22U1w9huzXX5WTUC7jMaEEIL1wb25vTeuejzyNtuWQf
DBfVvPAVXahVc8pCk3ZFjfQfFY1I1PMSMIeaQldMFyCz3WTgeTKh/JwutU/rLigp
xAmtWePPdT07N08zEU37chp8yJWoQOwKBGZgDJ5wA5OAsThA37FXCxcRxUAsfkbf
A3hBbgu2cUHcCybV1/7uq9UREcBAMz2py4U17e/gNoyg6EG0tlZ6rBQejhZndhOk
MDTBnIRO0rExw94Mn6nwHgtK7y8sdyi/nANrtc89uWCARt9E2CW+el4Uz56yKjjL
GrhfiOvVFIiAHF9Bc55+ZffP3pkEMf6NF2SFeS4x66GevY6RSHSOewnu0wyLs87c
Phq0ZMZkXUvDUdYDBEJ0vHdU7Sfo0nXmOYhzFwyAfuGBFKojTUkTZ1mUeliEYqLe
BeKIEgTi1LL406XqDKA+AkbENR2c7MZRbgDpXFc34X5kL8VCp9KAVLoBlPLlD7Bd
c0M+sk7bIDMFJiaMLekBFcERPY6O0nMmlE77hdLsRq5VqCisMajHYOCgGIYcLyEt
EuQPgijHgGzazeQ2DHAUbxxZE1UR4jM24EJ8/15gVJe0iyAMTKpTTiM06dNdoRoo
4pzmo0g7F482oA6hJfYq1OcOGcDpc159Q14oueMKLXwgBdeMAP5sME5zHiKTpxP4
6WAw4Hxmg8YsGFIfggpgOet9or8W6Wx/9MsBNmv5G0XNQSgxFiaKX3zOBttCbsbz
szG/TcAc+wYd8HpWHLU/vwl6ntHdAM9w6tIvdfucLrP47m6OkY4U9EbtLEeSEfDo
eTk4+0h+2KmOu61/kR/2wHGZ1BUqIytBL4scyXpHhDtkdQPw+lOHOjIKVJ71/fnu
R9hxEoEb5/ZjnjUjPPTkc0mhKjEyW41WArLy8pZUd44Ask8ar/aG4yNlPnm2mxfW
laevBUdDhYqD2xewEpF0jWZJlGE53AQCDmURM/ODZZr/VWXrPiDcaoxC1beBrxLs
wEp/IXnI/zB96sRzXh9GbAY5JK/Je2vDkp6QFORfo+j6rhIpDwoHtXUr7Y3oRq+x
qyLzYdZu2nrzlKbxInSv26vZmphDR/+Amfm9TcPpBAB1OrEg8wikEmEfbPcznO3o
XG9AeYySvvpex5UEIkjBghqk7RBB1aOdnGpj/72Yt26dF3DjgGsZW0+Lb2yqVYOy
plHD1gYL6UhBqYtc3tAiC9y3L2wTynl0b6+aqpjeqzqgFP4bbj4AytM1WZCOslj3
F84irNVMgfibp4q+XQTeKTniqFUqVS+1mqXFovAHNLhEpVaeWnnqj407veHzAMEv
boGVqc6cKDpVKjbEYAwhXTOo9ok9h6L1TjSw3Y0uJFmu8xHq1PPWMRid53QfsuGT
I1hmX81bbB4aiTNJ2kfzBc6X+Syk6iUHOWut6AT/0Oxtt6N5oaP1Crk1FrlNanFJ
uQ7IZS2MHMGut59XNC+01gf9awgekUZQuchFMhOARRlkGZccj+SSeS22TT73NPct
aGWCXJ5VDQmSw0omVUzmbEd+bhjSrQSypybCQ1MVej6PDvLpHfDELOBrKjtx3wH0
jecxlMTw2aQwNnYuoV4jQPuVVVZJbIb1mjP4lT67yHO3egSvM6GTjYg6BXwDYaJC
0fuurEzLiKROno2YQfZU7dH8xyAnwEQtFJkLk3OfQBXpj+YuJdWz7+c353LncU76
fix18fsMhAQAv18eevy4qZTWnK9ADScxVaPV0cobr3Awhiw+12c8WaIIqi0SQ8aO
rAyAm6hIXVVz/8IGPRJWp3Sn0ylP6ufU4MEnf1pdMH3GjbY9o6IU9zLYATusJdGf
50RTPill4MLHisWFoCvmkhK6puITNwvoQ4XI4ZyVCrgrX829dFkkxJKE9moHwA/7
tURduhIhiql8Cmd0UHJB82HcRZyViucxbS6JI/EHMIVaCIop1PrEIM1EskadPCYT
FVQHgXl4sy/URdD9akGW5seTrENpS6h52gpb368mBov1rP8PNJtf7QvwwPvC4IUZ
Oh+JOwn6GJ8ZL45sSuzNXre67j7M5sWG/WvedYC9nawM/aF6yDr/NFnWOsEVSwM7
6cB6p0QIyaEGEeL04sfUBBuxoLZouBa4nHfLy8Soqxzf7UAUSgDro/uUsS8y6uR3
JZTXQPFlPWi15HJiGWFaVcxVKCnr52nrlCo6b9g6WHOwor6rwo9GHHqSn9xcMva8
PSJKia6wceqib8g/LK+RMcNsEFk4UBXN1g10a5141JWyakenU7VMVU4LGAj86S6Z
TnPZvNd03BMA7LySpW5dlj+KBoxoGjeDOQdndSSXIvXsNh1DlQdfznqgXvYR3eFv
9uP4oF0PH5keWTOns52gNktXj6dVkfrIYaxqVXPQkuSSJYgMVro6C5tW1X9e8JWy
cHxx9SP67aHzPDW1kRC8f7mKnUtURdF5MB9gqc0PbbVrd64nUiArpXWpPUlIhVwe
OSqEqdUb/xXjTxM9Qf9hk2l5uJz0js/HKgtC+zcNc+BSvBhIV2KmWhLD65y2jsf2
ttxp4rYaMeE1RB92KgtDGmjsJhhgj33aYUOK9nZZD+1303VEaBpZGy9Go8fgdLq8
oPs2dnhSCdCT3kaDa//0LlGa5qxqNn3Y6WQ7gEk/bvkUHBDte5zgX+wtfHZqlVeu
E0oS1z4cRVHD8WYfANXTm75IXzjsDVngaEVig6igdWDLr0iKuMiqmjYzTvsTh121
bZYRCK+x9/VEz6yOCEhOjxemu6FlYhrDwgeHg1G44MlcjARK8Mf4g/coIf4b+jrB
ta/cBqlPbwNzyl2Pry4WYnti+aJDXmpcN5UKXpeFZvbF9UpOPLDoU2i9J7lO4Wlx
cguDA9piAzMwqJPTU2z18HzDvzTfVR88uOgmrX+L54rSzmhjHOEHKaUVG50hiS0R
Tz4ONTQlVp16QIfe35X4eyp8Vwa7GiySlpTV6Gb3OBI6prVes6d7wmhxfr8R6yYi
/WQGx9rCBdD6O+tGPTu+7chQxh+8864vwdMZBAc95d+Q4tuASQsDwl+6DiTJ86HP
AlWj/DjSbebbOQcUB1ZsKwEo7HwnYW05Slj1jXTSJVah1jvxJnV4Tdepvb4PFsZo
TU/RL5smj7FRZGb1wCrKfFc83HxYbt4OXAaSqjBNGsFbPXH2dov7MPMFinF+/kKs
lds5rtGtlJs+W2TdyDtvy/rn+YCfEYgw3Rt8dPB6wQX+JpMc70FN/VfmBfes31YJ
UQzLiGXm3+V4GjTtdKEzv4E7Nc7vwd/e4BdkdUN7WHFgleuCcZ248/hI8asnZ2uA
WJQNiIq0xKWtwvAofngi+lI3/VyYjPN43BmJK+2n9o55sbZi/mFINdMLvXvR01Dj
pfRTWK0d1Yu5PbNAmgynSvGbQXBUXUTZE5G7r8dqCZPDp6IRJA62u7J8UklJ4MgG
KOh+P47V8GYGeABryBF6WZZg3UeArlmYHl1oivrbT+HOpQ3Tv41V9yoMMbCw77ql
gxGdIcj63OyQRYfr6CCJHBjMbI9hAwoi+CJeiWRuuf/6p2eupmpV/VRaEPewBIfo
N41OuU+mLcaXVnavfzjjB+39v5h7oNLFKR1lC1uuduSceQZSlCs2F1vBaVoAfXg9
PHvd9RQpUuW0/ThMRDzGE4BtwVdeZlRII0ehlp5gruC57g7ysEyALyrC9Yz011qJ
6tA6xrzHQoR0K65XjmxlJf05HE2CyOFxHnjMETRW9l3KbsvHbgBBFbO1R3ypi1p6
hbk8eN8QaVCBwfi33sL8oZ+I3u2ThsFOA7lSEauOx/K4Oa11Ze5wUrU7ir2m4Qx2
lwZtVn8Zw7uBKBpzTvEDjLAjG8wmPoCm0ZT5Kpaz1p0EYX3g61RK9jHzT+4xjTei
E/sXjS4rc+PKwrTzYN3bTyN7GpRBYR3EmLh+ebCntolMutY82YKmwG9ZxHrbV+0R
EQQ7RorjT4Nanijb3ZMMyJ8xOm3nOfsZWL3qAXs4HDmjVsZGcmvrNFn8i2Wx1JSI
k05pd+f0O7VudrRN7QU5O9bvVN/JCpTKVldunUrjVpGfhQNCdv9DyZATKWcaisYS
gIH0fKnBYmLmPHKzzDmRw+SMmiUCAJO2TAOBaQ5mOqlZTNldw8seSGRwdevFIxs7
pjWKgOU5L6PxIHlKEYMgTzgDh3hqMICUiUgQYGQc/RHhGHNV6DaOw+hcQh8g/kaj
tguLpcdJ+ejctaadhg39rSmZ0uk8N+1P/o4bC7Q862vBZVt9SE+8cErtHnbDgHrR
8fSh33QESPsSNEoinQZHxpw1VT4wLvz06rcA72d7Y1u010q82sHkaHPuwO9uaOns
f3HdHudcTsFj6SrKYs9u7GVL/wIGeKVC82OXgfEMt+sQXsUp8qZLYULjP+lbBIjQ
PFEb6WDz0qBiA9f7YNpI08xhKIlFhT2oAs3QHysv+svdpjLc5LcXWLYFZqPoN+Qw
05UPlUYAIgDN8L+ZjpJ+Op2d/lRTSlI0NPH84/34oukeWDj6kQ5Jdn2munZRbT/x
kudxfkNrkYRIWR5wg1b6Lu/wjDPiHJ7I8T+r24kD0yZ97gV0WnWzSjlpkrsomCec
vIDe2TkT/CTHmELYxSBn6EM665C2C+xk/8p1EELNtl7BcRBEZ92VsNvjfWl8Px60
/AYtwXu0OsNSLhApoRwREkXMA2MHuDs6WJ1FmsH21bN/eyqNxR7Gjpi90/xlIgGF
brKCbjo0ZSEJsea2e+RMddSmAr3AKR5bkMjydjxiLH5xRE8ZzaNoMrQwdOLYGc7d
h8vKcimCCrAFPTccGxRwuPoMFt3bpqQk5QexmcSxXfpdHtTRDBN0Dstm1BwXW9J2
9IRfXc9tMeTOtSjMqD5f8IlRB/PHkVciTMzrCpPTQWn/nECkuz/XbZ7YCfnoJMu8
6z45ZLQf+9K0ak+xBVu82vBX2JOrskLAdS73V85oAqJsuqNzirOcvyd1+x42W5U+
u8Vq3ZsaY6S4Sn272M4tRWJBw8aDxnwaC4EHxq2aUkIQjZhTZExlZmgxkywF966e
roHR37Wyfm8H5x7DsMGm9W3fdTZUPIRPa4Bm/GjlWDN2VhsitLPqhYesmtsh5zQ4
8IPTgO1hWUYoh+HJT5vbXUv87Qg8QxQWtix1FhQuBFdNNcJPKF3lwXTIQlbi9PFK
7fr82E2+PeH+iM24/evxARp0kzYxg0slMQcySaoJfIh4nZJh8R39PGcL26WUIlp3
DXmTEw/6GZ82yY4r3ERcFg9an3KQi6O0k1Ost8pxGiiHKCUyJQLu8vWbhXN+9kF8
IM//ej8L+ZcCXJZnH15u2u1qcjgNHktWHF6Ype4kBnT4jnPPNumQRzsjBiwqF9jC
Xm7cMzHfibjeLgNHnS+12dZpr/aWql45BS70S1E9yF67/b0+YGJdJ+qVEReAN6h8
k3iUcm9FIN+6eW6xm3PIQBCy1VBb0S8I+w6JlXBIDJLYOFmOMzzcGdP+VYgOzl7G
28sC230EJZ4mGC/m0CWVaNVrX3nDPonqP7hEoPOJ2t4VThIQixT5QrfDHWQBA4aR
l3HaJlO5SOHq3WwYidHDJKzNVMFb4K60eOp3pj5RKdxOLNgLHcU4ggXz08+1OKOh
337fiSVw1HY/GF+HroHeyM4Xh7y7RiYhKkfb/TKlOYetAHFMd9HKpSTcBvZVGew0
SQS+AshI/ANaUyallC2xKWKMbez8IVEAAQEy9tI5ZjGZUfSyejatQrTnsPDUEg2A
QEPFj9Rkq12+4pmOu3AVk3ndgjs1mnaHwl94JgOVp8x/Gr+AQJMnrAkGQb1k9Hwv
3cQSmZUHXFihKLqAjxZ8BQPqpeI+2LCJ+8gNjuxMUsixDqMR2euUSyuela5+UivY
ltz7Eety0OChB3A4i2blEcQYq8JMqbxLti7dKqRJnmhEJCydj25XX+9X/vv9Y6Um
UQ6HeEDlVi5uZIYBEkB1k4XMh6K/XDQqzCNXWW5Hp7opiyEWjA9BUQoxMdq7Mh3i
K36vLyty0rwJAoYeqprfSOZJN7N9e5tLF4bTK56KQRXf1n9nrSMe9ZbyFT8QvuRn
pcqUBLZcYJgNH4PD6AS5tV8rJvqeZvhH/cTnDxbURojnhjyoNjC2AVA1JsEO2edc
XLFgR8bXcvYfIXhzz0b4XEPdQUIfMH+D3ARtDxgDKK6VtjLmCLR6ooaL+BcpQKlk
eOfftbgNU6Jia4GxADlMgpTAC2dsbGIBo8nS+n3MRZ7RqXgz7LNF7xDNu9htrl4Z
5yfuZrUAMh6rdDfzgyfIQuUQDl0SRU7OvYQsM02BK1d5OiqRCS/rthlD4TB5zz8k
Qi1E5LuXj+G5Mz4T++yWwviIj9P2OESJuJ7H9nsFWtHOejLlie5+GUmt0l+bCZ8o
w41Drcx8AFS6o+Ky7kRiojfW64UinhGh84+jC50aS3ZVjq0DA3adzPT+H94vjUim
k2LmLqX+mtOrif3H0GAlQPsQzy/6XjorBL47yhkeF/Q5y97LTFy/+azCF7NGlbYa
/WccJN3VysXohV7ji6EzT/8MfnPqr+W2lUAzq8S5D/zy+vlCbygS12GJyZdq9jbo
8rvRNNH5VmG11FyRla5s6wqmRfElmfV05cXvphKDBHFKD3ACHHT/kWE/dR7G/C+T
xNeisD7JtkIBVxIXCifNWz7c1MAFp7C4iCnusJsmKqVtZ12nubTVSZ7O7/1rfo0w
heQ00jm7AmtX0iUWbmG82rJaQwluOULKJ2NpiWe1oFwksPysW+KTl2xW35CJqz0U
HZ0sGghizCYbmaGRqhNR93dvQrMhWkXhYWGUo5vlN3TLFWIcdyBHOIZxXgQUsywE
JBturvbTSsfTqkdYF4KwQjLJ7XILx1HjLzgr6f8NwV7tDKadn7AZiKHTQBTig3Us
OQau06RZEF4kfpUjuiv4U+KTQ/7Dr4T1jSy1OyjPZ2gKUGFFzHiJ2icD4O5TQTFq
NDbXr5a9BGuYj55ZrpypHewv3Lu67eKJepbIGM9X0bOgc95LnqkHhyQ1bgktGrQS
7wyJOSjqZfEqeCIo0e1yy2azQ8TpC7oc4DcriYGWLnEOjsCRPpzArRJgYG/KJX3V
2MCQ82U3fyta6lJTTxjuOfp/fIkXSIEP3KibiLi8mG1klNzev2w46FLiR0+QK5oK
uOm6hSMLUEPO3ZjsxLezyjPg3MYZgeANmffuwjTijXYLPYN+bEGTIgh6HBfu6UpM
TW027Go7TP0rwz+E3scbzd6T6c9CjMiKoF7PlJD3FlQO0nF/y6GpXUjFbd3AZBql
6kBfMKQfANuE8ZrfVTzW6wvAgMQjYhV2a83qpnc3syR5O9Wq6DKYeQU1dzz5QtwP
t6xR9Bs0VHeDIIoOVOtMnqvB9boNbRB5doa1lwzKMudCUFW2PmeSLWm9Rn8Upmni
IfWazvBuX7kd7UXZuHICgnJKqtOkKup2tbf1E7ZdDtfSCh8izW2N5QDN08UoXs5D
I+tZ3EyO88Ca3iiQabfGb1pMmZgsBqhWr3fQfZeVODK41Cko/qQJBqhDbaoYa86L
onQ5MQ8117IXJsj8Zk2t3AYaV0zIlWQvdyUvGfWToD973S8Dovdi+8VnwvDnV7Gp
o73b8n6EQQbKCaNMdAxqJr6FOdAtghABt9J/yc0FMeRYdhrk9APt+IfrTXxhJn2o
PBt8iHnFhBCSY/3PwB6mCZIxdVKuO5UK3XJa70c9xAnSi9PNX5VQSyb/AgL2wsjD
wmkv/D6/PQlASMMozFoTpp4YDuFhyDs+Xxb6ZRjueOkCe1nsVEib9HkFIifszQrY
ppDUFPzfF6MgrVSI2x+1Sir4bvupRRv51OMGJyuxbjWV1ZEGvYZVnT5RUbyRj4Jp
ZSt66h0lxFVe71OgbMjV99Gq7jvZZshIF9JPx+JRoGsgY0tKqVeRqPZfrl2votKc
9LaIYSjcCp2UTZ8U6FHP4kgG+RCwlCKrO7u33ZR3AugxU9tqSEce0tV8tlLcVBxg
423n3UabbqqCIdBQuvDQdn9xVpDWBm88hUhjqmWNdtrZPqo97kBZAS8JrpoOR2rF
JxC8ThQZMnJMxV5LQa5HM2WArGZxzlfHk6hdGRHrzhiYeMwGjbRGsCUzbP0hCq/L
Id2bCqXzOWWZ1qykC9MR4HoIRbgqDzf/4/RuSljz7JOqUYCsllb0BhGV3eO3VbCq
XtPKlyuuNBGDorrcIgfIs7Z54w1Z3VnyKFgYL7UGqkK2NT5dZ41bf9nsUFc4kpHV
sXi86B5Xy7osQYFpJIHaB1mOxBEwV8f+F4RcDlFUqMRxsXs08ZT9HDRPIr/pLQOX
EUMRP0YOz0BbBo2ReSvkO7aep7lPm+3LojGHystfzZ5pBsmlSbHaBzmoGwtMlbIw
SqcR9nKw6ROttvbyPIbrlJhrp83bZAtgobbk2xH1wdj8LOwsm6J/Ov52FGmmQvOW
cyb8mzgbCY5a710z2HUCVa6cqzuo6YMWxgwdj22xI0h7LNtkvwpk7307W2u1fBQ/
/qSg12Dizas9JnzZ/f3apCvBAI2tnkYIVqi2PglgCnDQ83xYgPePpTscBuJhSVcV
RHQKWuYXQ46z1CzcavdHBx0rwEyLvIBxnEjJwCp/y0+/fFFlZaNhcJjZUMmWQSvd
XfH8BpYOqvzq44p6qcrMJRyxwMo1t19UZV7XMHUm7/UeKm4W9oRQJ52CbxOFM2t5
s/vrKUTwkxq3+iQ6LTRcpGFW10X8CvJzyT6vQBZmbc018qFZ6HbFpzhbJU9opeT2
YeaE9OnezkcRB/omD1U9B/asN5a/vck1NZSzdAxJBT8BZzUREyg5bJaJH8BTxd6y
M5xpdni/5Fz31Jo+nrpsHalJaLyzHH1btkV1Ger5+hdeyunAJb7104kpFjh4jQuN
N6Gmcfja8W27K8R8RcGek/VEY8y21E2ccXHEXGlF68Fgd12l6xsdq2rjzniIhypd
f08scMr6Of39+cSSHaTHdKxw5yKHBHFnJCjeqQpECMKKa7xSWxTWDPdbN1iHnQmH
WAgeducJqebZ/drpjQtcXdpI+S9i6LygqCBgkubAsIHIYC1rAOXVSsvb8HaD67q8
ydwKD5N/GslUCgXZDjWZefNu/RZ5CHTcCbIUFu/znkll9oEiX5p9Rnb9CKVDONJ/
Vkx+wYNRXa1DVYhLPCZN346khqQVJOtWGAkGNqGBSEHXa7/4He/jasrxxRIOjgR7
SHXB/MpjdoMi/nOG9PF/ttN6UkYA6inZ+j4MY1QZeUjmpvsrXynXWNEYIqmDVOty
kip5RDy0ZhFn09ORMSM+lC+1xzDZQO0jgM+jpsnyDCrl0xgsrlOVM0ULlDNQ2YiO
vACjM6PfmqenOzLvYTc/Kl147Te4IPiNauQmuZ7jNxNlMaq+dhRvfQDkPCjxizen
U++JN89wZbpGdY+5mFnuMAyoofd8Meko7NCOHa2Mkjn6dc5KM2WgzFozUwhnGa+C
uJGl5Thgt/59mVZnjzx2Eqb8SMcAsYlCuViOYeC4xaL33gCw04pw6x83yE9lzLUZ
m82Q1MCPhVsddFDroD0wARMbTY9mP2SZG2sezMiXPXOeG1D6uuxwIa3X1wRaYm/x
iFUbRyvQebk2KVvmL7Y8AAbRSO8vxAy9qVo63SApxY9Ma6OttVG2dXR5Y4fb9ExB
fusgU9PT9WggSmqoxlZHxPDD/qLveNy2s/c9ijGiIn/BF1v73ELPINPq3rLk2nLN
nDDp+EC8HELhtW7Cth2XpcQdhr5luXxti4TxVKz4HvwW46oM9qfrvKW2hHD/grgI
hMZHyPdkDK/lLkfLYSmdIzlue1whRfjlnxYSk6vMidDfEK9tQuk6UHYZIIx0colc
THoGrcfMbeQ4RF8YDO7izVbf+cIoDlznAIeJULoHis7XXJ7tqeB+5KqEttDropmJ
pDcndCBFbampsAy6chWVDMxl2B8crmqeug5+eXy7GzzGcWB2lDOqa2DLX876hKrl
7nqk7bllhRfJcg7iiKkpWOpJ7eZzCB6wHVnGGTYu37ZaiTaMtI8eEu7goRDlnzqX
Zked3ZVJVAAb+OYGaRd5EuxC2YvToDQBSqB9Hvh1zGzbegVimrLn+hCtOCo8M0dw
RW+7vvojuNK4EJ11yf3JV1sRPLz+ocTgnA0MTV2XXxcKcq9uMzSHeMI1qgGkXJ1U
3cmRagqfH6ac4kxND3/lkdgn3h1vr6+c0jh7GJGmdBU4txE7KifjkYEiT2IFYL4b
VmLvnA4klT9mcaE5FDGrLDasDlf8pxExrHCToOyPJxdOYsKzifaln7FPPVrCL/Jn
ns6XYWOmK3vbbp2ZC0sNgia7AHgFEbCVOahaz+0lS4Krx2oGXFnxTQ/goCxwhMJm
/Ot/JY/weYltUjhmqCJgQ/xb/4F+aCCTWBgaBPs/gvpgE+HRNWFBFkuIb7ljdYbk
I22m41XRr5snJ31aBwo0DWT/mlh/BxHffpHYfQedOx1E4FzwgnYMIhCjnvIBg7Kv
rQ6paIIWm1fUzIK0P5T0tZQMlI/bHUxFZu4IZW04xoFIvBSDGF+aLviAo5dPeT6w
4el4pQ47qQsrY9ColwJoD/GhM7ZIdhu6fVL5LTK9n5RMIYcA2hHIkzhkEBS5zfCd
EPTAGXG/1hFveTIQj9wM4O9Be/7Meaj5ev6My2quBtyKdlQL5+5oaGf2rhNnELIl
nE7H4sISkoj1Uxwc/ElfKaCUMP1AHCGFexilRceNJSafqWDKl5oJet2kre1mupIQ
fcKpjDr+qlIlTkobg7NVUT8Ya22VhZH+EsQFQ/9DJd4wUmOEOfhk39+RdtagmQOS
QyRGfznFlhmuOODbBTRBiunJq4WWhv9S5BoCemnXlMFIBW3yc3XLLLWF6GSbAffr
U46ZdqpHmlwZPvF0mZrCdUrmHUy2TWQ6QAMqq7/VKkv1sVt26m9xt3YCSC4l2fgt
FqmQ2UOGlRKHjQN1qe6CLmAvRI/0yMTjE0BDpnvhDhUvShE91Kp5wiCOzRBsWbJM
P/3me1cNuYtL5uoIIIqv/3w79C9XEpU0CSNlbw1UQXg01Nm1dx5fcmcrDvSf9PKl
u53a9WQexMDPSQIOJ1TQjxZalc/cSXJysA6W5KFcd39MyYT0PKd6SmChLmcertqr
Ju7HcVqxhKPLvd/Fe8TT1tN682JYQMN81hy29yoYujGqEkOCgJ639LBCxaJcpMjP
vrI2Ty+p7Vvd0L4EwQCb9VnnPyk+QwkCFi5zGYdKb3nF4mVap5SWpZYuFhl6xRgN
sUgWhC9Xhibxh6S6cp2OP92GzSSfEnQL0oIChkFNlQvKMcPOKBaoETAEVRpPd+Vv
VdZ6G8mPVHbjfuGve40JZ6VPnxQeVwE7vVS3eRx/OO6O/fcmjkRIsbBYOALVxVTt
tBQRKC+pWi0cK4lTPnCW6R8LitHD9Xgp8RapPP6ds0GcMtHpz3662latfdf7xETw
RssZSqNTg5dZdEyrefpXkpYqiADQu9KV28wkOwi5eHs6ueq8xqpJYYfzgone4B8P
4m64T/Rf5iccZAS8aVf9N77rLJsnxB9ZutijbuHrG9f772EdN+GH7BB30Ew+G+Bm
DSmLOlIt4zTWx7XID/TGVwRDuwWnOMcYaEAijcHNg91wDy8CH0Tb8yzC2RqwOUse
ucKMAuuM6VjZ3dkV/pP8Ri70+bCOXQ+IkE+wlfLiZHM1ChLATyVI73eFiOol/vVE
WSvo1QMTK4LyHS0nHpndtLQWFvO1l+LzBNP7AxQgzg76b+b9kO5x/Ia/hYu39TCz
JzQstR9ufpgNarTfCTHIf53fzz9CGTIAmebxzyVfriHU8dLHPab7dwPF4wc1DMFu
M58oVQTKuEOvax4O4hpA66MD7ZBTH1wO0m+6r4wM92SfiAa1Lv0fOoSfVDEOKZyW
zHgIxsz5lg+JsnLe3V4DeUoIIolYGswwu6rQ4TVnZU2E2cpwiMrdfaHJgzSJ4SYp
tWhBbmbuWCO475rWCELqoJ/iy+d0o+fVfg8ggae1f/umfGb1lgseNtfktT+t0vCY
jsrajVkomBZ2xEf2WBwCPLWoB6PqFWcm0NY2jtTDtDcqwZJK/oFuSMVAQZs85gXz
T/VfxcFGpkdPV1plRCDna/5oVK2eZup4SUvxO2yOnobauhP46+FY54QMlBfoLG8d
IU2W3BOTzf0cP0ZqULZkjnFcNRmgidRa2+bKGD0MBMw0fFAEqJlZzLTcdZ1sGyeM
AgcGWcc/tRFXZASXHWsXdq1VVcNoLPGmSmRc47OcrpNdtxWJ85wFNbV+1EfUUeAB
LtABxYiQrpw2OumEGTXNmgll/cs5QsqpR6xGoDZcl8agPPzlJQ/ZjbJJv74Qpowg
TVqOn7GDP//+V+aUXGsa7OEQ1WiqVWPCxBN/MTeMNtVcbDcXU8c0aXNHVi6iVshG
`protect END_PROTECTED
