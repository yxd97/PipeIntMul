`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50n85s+mRC9krvj8aXwDXI5PaPG99GWaFhrjnK0bblkH3SsHGRUMhWCsPA5abY1G
IsVYeTXPWubtOagFUthC+kqicHBpc2HO8xfe2LklKVOg0lOdJv9Cc6zzYYfEkbV4
IknNvZtasa6N6U4hq62wHsy0JSJYuZQrwSEI3uIiwV+XfohuD//vW6RolyFFDBlM
K/YfAj64KqO7ZReDccbJn4HvR49oSwj57x3nAqKR7zfawQ67azewq6ZexWWKPO+c
I+ADoYGbrjP1m9Q5o8/tzNq/koom6naWzPTWRhs9GEmosxiVKq9YTtuGdOz4H/e5
kHoSW7Zi7pYiV7eULwECfc/4+PM4Q/RXt5f15KLCOepJncL7RDZEntEtViUdTjHK
TGv5Co/ve5Gv+FnQiJMPkn1nFhXWzrk/auoLHmJLSTNlryUCSSh79+8OQmA3/HSg
cxOB5Em6tvvUtjvi1pKHuQAidsHyj0D+iw1LD85Y0Cw=
`protect END_PROTECTED
