`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rvuqcs+Eed85OuDwRQ4XhlUmlNHXHfv0B9GwO42xj3HJYPHzijJ5TckNXvpR284
XBkT8eRKdtC0NT57sLE+bzySZ+dSW9RuVh5hgZujFr3PnM+EFPX/kCicppbA9yUC
tZ4b+TMlEmoaMH87yuuqEvijAT0y406gjIeS8zYFdU1UGBgtbD/FzpMYGZwgKEkz
rxx96hwf/X5zxKHDbH9FNozZNXNhdRXNVcUQVYzsRAg81n68bR9o/9kKh8U7UFfr
zfHQW0k2FsYXDXrNt42IuSBSqXoD6KR0NAfsOu4r9Q9uI95qFSbhoNFVlCh4xYgz
cQF3Rg5zQAlZUqe2cGMK5w==
`protect END_PROTECTED
