`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGFJZcQZ8BMgU6zl8GkcR8daZ4Kfsfsk3OKUm5FlJ1PbRg7vrXG8V8Mgaow2y78e
Helnic7UC9NXlFJZcig2UPHINihluwoIe9XNk3CYO1o106FtiZqyqiFhoexxr+ON
uDxGN9wCvypMma3slYFaE7Cay8pjuaor5xL4KJD3fEUDv84fgDWonGA5amr8Ehyo
HKzjavx7uSgeVy+mGj8KBUFlsSxGr0oKFXvjyny0TZXDU3Akk0oFI5IDDYO8HxKP
FEPR1oS8kJr7PEyZFvsCkzmJjT6iDIS7ZXMi+mqtnzz56OmeYNKHJOOLoRkOR3L3
R2i39siee1FsyADz/HZywZbyWCVST5x9KZMfaX7SR6Ymq78N3oncDBu4YlaB4mSA
WWFHRgM1sl2AZQgPs2wsGc+tHWZCiaGmPzqql0JnI5w5K4z2r1RO1ao/zNkg76CA
vRmNic3imwCieuWdw+Oun/ECiFOeNtOHk/R0l9iJh0OEYIdubmjQqGDQQIzkNp21
820/yYM1Q/VFxyvPayK43ENHRm/R7izWT/HJ02jX/m4=
`protect END_PROTECTED
