`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V1GFPC4czPpDbjgQRGurcqgFt5XUk6FWenIcwIoINgt5ad9nNCwaQSb/X6qll3Fc
Tt6KlFSe3Mw3cB6RC1z7edNSwv97TupG/mgUdRRyZ0PmLj6e7krBf4NbSxP40wak
pCQSX7G17Wwc09Bvrsvql5oTIClaK/mye1UFXt9tGfESSAKgR0ri/v0GIjKBf/wH
VcZ6sIhrEfgwrv0PqI/mJx3S3cl4/yW/f6ude+OnnEE/vbggs9Omclv7dJEt3MH4
lpkXipkdev+ICZ7FVRQzpzIWgcw0Oe00/GrPKi8HMAoJkvFH3q+tMzEGTDkOUWEe
2ufYybttVnxIwxwnTmVs9J2wml5SqZii+YpllGOSeprBhn0H6kefoeXoOE0tFerc
vjbADC8MSjP+MHoYv2TVtpX1omBdbQblkzppbCcSkhtEsTiH53bzujRN96zHfak0
`protect END_PROTECTED
