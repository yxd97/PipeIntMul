`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Ta5tITdljoL6KFbfrznxB+7zm1e/cIlTmzRq8Fbd9JDYHwbZO5QB8YUjdZC7hDx
SuWUaarXmW4BD5PSP63NC2tFMJPpwf2rJmnpeIj+SWmDGSIXdMmR2q7r4E8p2nz3
MG0Wn2A4AYf11lljqYndgF5Lu0ayxCuxhxHF8GW7fjJ4pMNirKoO62yR/VBt0Ydm
WfSSkGWJMgswK87uxoDi7eP3Y6WpeN/h3WpISpxDpSJiS2JIyVQkYo6hjd8D3M+/
jyRB5HsF4mCthQV/M2pck/8fbRoquBkBWUfsYqfZE/EPb+Rgrhn15eNGSOxmsbNh
th7TicAGqhlBTMcTuvQ++bhWB5Ahhxe1Y9UkCfunQKbqU8zogpl7XhTUAtZnAB9+
vuvSGHAzoCN+97o+PcPFSw==
`protect END_PROTECTED
