`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZES0W9pUfCl/ouLdKRrjTirLqsRIZbX0CotBVAfW2y/kJA/yDFAI/6n3nozYuLdt
KgqunE2WD9AD0srmrDZ6kP+Vh9sx9O/TmUiq+dSAlkKu15rIziO/gSttssNSiPX1
Ov471eWI4sMvwWPEYTMovoH0WsrlfUzdWYHA4A+xUQEcCxSutq/t0rDgWdf6R+jl
e+7ZnwzP586nV3s75EHtGplFPZ5yoLHVLxeUhKQtEPXxaeKFXaifsrrMo0Go38s1
+rvm0a4H86jWvHsl8wFgl/ytszxeaL7uOHgJJfdG31P4V/qIymprZsTdbQR2aeRi
stF04ji+5D9yM8bJszj2eSP89OeOpbbYVX+nNkAyXw7e88vKbdIlkCebOd0yaUyC
fv1qHErO4Rd9HPy14FMbfCyFtbkMCilzFss8qAwbfu8RNHu1iVBTrN+llGcJ6y25
7nw2mnPgX66qvPZrZhdV+xIG5Q32d94zEX9/jNKHEX4de52Af1ma90QO9V+smfD2
6sbRTtbxJewtes5RsFoXm8o5j56Ox4fVwAbudSVtN/sskMbApYCKhiKvAVaVubxr
5DsqHBOKbeGhF03TBbN/oTTRGWCBnFS18UerEtoNZaPl9N83QOfPtMnkLchgxZJz
7eu6kMHUzP+UvJqPKsir6FS4yRgC7jfVdrIyBDfhP7l8wrAIBvApoq9cfcPGsEjF
1XvnEeYav6tZDmVCEDiJubqp9Bsogv6DO5c3/bNKkBDKjsNxCyXi+E9uEFEULdsg
OQCLQhtksDOIP8bXblQAamIhnudt+R+tNx701YpXOvv6mYur+i7uNygI3gXWt5jM
zv2V058CHn4Cn2QHbO9gs/kcOjzk9yPIEXW0JKn8wxUVa25gil3gAIxtDxQyV2i6
sOnCsNdRkehK+JrOk2zFRo+R/48Fow1msVFmwc4v3K88BFIcA+Dxa+42evGKrDn3
5npdPRuZ83wMcT78//c+tBWuKpAExns+OmScUpKc3AL3Nc8TIAvOpNhkx6BPD37R
auY/wKidmm5ARvg8NMVWPxFKiH8ZqGnplUKY31siIywIuLf4TFwTQzjbSe/ZMnIQ
Kk165yykimlzVOpK/cxHfowxp+NQ6rgQtcFbeKOi7FDjj9ogjxvDTYH4nbDeZ3/3
`protect END_PROTECTED
