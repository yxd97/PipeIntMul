`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JbYkkY9j3/FvJFEFOJmGXE9tfqQz2qkpVmGr8KZ8CZ9Sun64/jaNYTObqMYnXFIy
eNjVfhUW9KhOPZhhdEaVYlGFsDqQ03SY6eoJ86bPz0qj1rb/nqVK05NGGlWXEIye
YIRj/2BtjdvlgD5cav5QNVH1t8ycZO/rgIEM2ldBSk6LBmaz8C64JetAVjsQqREO
KmtR/nN43NkoyQMtb2GiZDzcBx705o6W4i4O1PE2reFQQu6EQRF/EVWqsSFtR/1M
Cc47gH0spI5GgYw0DNTys/j4QOz8thiLm9tu88oKGcdxn4EvghEJcveePU3MjYZz
CyxpYak4gzdkCLNNyZUxX3fAdvN5+JU95BoVTDQy9gZ7qwQkgVUSTBHSkY8REhU6
IG7VMolKNascMlimWh3HfN3+5NwwgFFdJvvr+7KFibqUg+k3NNLjAWvMzaHk/e+m
XXo8QFT63aEbQb2+9JhdTOksWSRNBTfPb76tUm9Pdd/lpmPYWJZ5W8HSHt4T4QKW
hrNN5sIHnMTOvINrOBJ8PVdo0/nqVGZQIK6fDZXxicQrytCwLrgFxUEjVxpqKQdB
Lpb6PnakPWbyW2GIvcTyOzWVFv6lbHf18ERQ3LUUqiiImtpl9jPMa5wDQCXKISmJ
J9OhOIQl5KwqmqiX658Ku1JP0VmzT7Cb3Q4NSEH8MokX+pQiv1q5WafzCQMHLeIt
Oo2oZcJTIQ/kDc9iM4icTsRsIaqqlurecmutm4QsWLrWBqq1Vod2eAaUruWGuoTS
kPAajVpysT3XVul4FpzQsQQ4q0UnKTcf3oHx+ngtTdMH10THb4JxqPa97ENZC+83
Y6c0PgARXZWy+gXd5xxkNkPogYItXs07QpFOxnSdCknXugWOi0ljiLCSvpLtGnkI
`protect END_PROTECTED
