`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y3sGc3FzgZVyRjuTjGM7hb5T8AB/AiUjIinYNYBveTs+C+Dpyiktiltk++Y+zYFy
ZfsnFEMqJyg6m0aMui+0pUcn6hgIQrO/WTzgl3UfddPTcRt6OFmxDT2OmH/MYkHL
dSe34ZuVCAy30XPGJVyr9nP1ytY6dX34Q2gZHWGq6VqxJz3JfDSeL9ly793QDzEJ
eDvnHoatzdMK2St26f0NioJL0mc7BHn72qqsbNPYh/6qr3ehhi8yj1PFCvgqbxCj
Tp+HDA1TyW5hoOCJ0FW8eM90RS6NiJr+rZB0axKND91kJLbkeUPPw4RmhXVA0C2x
4AJJFx7miKulEMm2KDXTn9GOnT0r8qV+cZQE3PY6Dz8PXv70MXQqG+x3BTB6zq2Q
sQ21ZAczgyoF1/aCi5pKD52Rp62fJs8JpxnlyHgMU/qWDQwfsnHI3UEKqXvIbEy1
1tv9uaeBEf1hXkW455o8zmlAG2EQgOz/y1amqa3GRDjIiD8xm7Awt7W9otoXDaI8
0ednWpW9V6xA5NatrLTiTmQWOR6/4BTqkVzUEuUG63iNM7mHx6Vja9XGTkvU1SAq
dQW2JUkTqJIDRlKgJTmuObmAaMcqeX2fhvi9L7wN2eY4xtnTRo3zP+9P0/ZsW72S
GhR+oS2rGnoRbW1GICq8Rq8VQl7FnEwC2uzbvCJUHMBs1VhdcfyD30VvPO4g1WQX
2grTB3mAa/NXeot2B3zAaHfiSzmOQfE2od1ETURTS0l0vTG9C81pE7KnSRa8Dbxg
Af7DjzQMDjIV5uBFgPxXoEsl5CPgzKgvw0MJk5igJB/KsserMxtka/IEVBBHiOtB
oftgIbJksHgAjH1t2WH3wSrcZgly0R1mZKO5jxCfWFB9g0zfSBf1E4kCGmq9Vpi1
28qq+ohQyU8Yu0i33jq+vnMNTlEeyWv0Ryy/TIU88onTDNoVM0aB/Rxvlk3OvPZM
7K886c6DiGpxwGzBitSkORQiM+0lZRCQJ9guSr0hjO80/E5sHP8WbiD+QpVoBZaY
YrBNNDwk8sJw/bivZH7E1GmJK6Hzk/FX46vHpqnz3zVc9mEDW5cSkpgTBoqhtsPe
YfavRjCqUkNlEZMFFQ3p1Q==
`protect END_PROTECTED
