`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4fJ4ZX7W6c85u9+Q+mTrLqVPImpxOUiabO/GfTvRm8PY4b3e9KwHdJ1F4Lh6FyM
hF0j3sh7sy8oJa8ht3YRVBk5cu8nX8N404t1TEmvotEfyAunxWKvyQ7gKq81m+z+
1wasitR5FDx0Z/tFfrJVV0DrLdEEEUjjLL/fFzXyCGy5soy3dz4i/M2YZOhJQGt6
fEVgn91l4zxcJl7930jpShAZ+ZIyWS/o/fG7rqmdJzPyezrlh8U+riFJPVHW/5/C
Rct/OOgiJYbkBFSLIj9l7w7teNhMf78TfffKw1mRNGde5uvEmZ4iQdTQrYWixtad
iMH2BxyVef4ttYqZWTOpvWh7MD6GC/taJIwVtZi7EaYPe/LvlS7Go/CX0ydbv7tV
pxXxjqzlfg+88nqv90y3qxTbVbsuFDUAdS4hGfnb5Jd3ozSz07spJPn6Hu81vs+9
Tt/dtkv5utAQI0oZxwH1K7Z27PJDSPSs5hEnlJ8VWtGQ1PkXyFvwu3pXttD8EzTq
Rys7pyNvFJs/wfY+S/avsNSngmKjftzlAfqBcQrb1Cg4vZAKgJ9rj6gHbz2uVsh6
fqZ9ZJ/VQ4xmzpNkXHn0SrH75TGu0tvzFEW8cNCNwW4ypcd1FlyNkjWnt6Mk0zxD
YiNmuNpWJUF6QLtfq9/KdcKkf/R+iuGKNAvRK9+h8DEndTNcx89LMx4sELoggelA
Xom/HaJbOoctUftChJebzxvPf47m4Gu+CAFLZbR6EBHVbshSOcNF0AdKx4FBIIMK
UVwWV1eszOl5W9K3MoeZyFRUJVHPg8J62TuqYL/EFSKLgzKNMs+n90oTO+vQS6Pk
20CsXQLabZuoafGUlO31LteSibzRMImjKcMatxK4ZVX/68uamx06hvuuRJbGVEBC
ezmXUZVx2n9Npdysdu1CUdc4ZKcQx1k6W2tEglxNwMpNmd2BAs2wfE0sl9AuK36z
/5BwPb8TiTumqhJkhB+wLbsPhhHNbat/OJHlwyY1oQLVt3B9JfvNayAVHjmJOWoA
UyeMhSrv87IKP+Td9KWOceuviwaAVE/E2pyDgR2I2D0TlOVm0BngbO1EW2CD7m0U
Q1Jjm7YcBb8uSgcFk1AJtQBEeKZ/2ppYn89/egesnTNnkGn6zoGjieq8izLQqrKW
gVExPXB41azXu2G9qgwgVL/iEyhluDxtR1AuUp9eddk0nEt8YfmZR7F7IMcgHT5a
xiCYzOoqEz9XLnnjiA6wKGckYmBTuTtpaeczPXotJkTSEcHpfHWubrLkKR1itYVR
DNU9+oJFmN/qq7Y/8qKZ7uLjRXJjTxfj9AzSQwn6qM3oA+rLfPkfj6TNMvLQj89N
UugafqCLvjwkRpIjfjRsBJ2+zihVAgZHeS+UhCeVQb+Q0xnrG9jnCjhloTcIOSJX
NtCk13mmwzyAXzAAesCLG0eNlEmcL7oACjNh0QFQTFhwoILv/M0j66UVZvUF6OiJ
c5s840uvbJNaTzqsFQ+jvQ==
`protect END_PROTECTED
