`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HNrkS1sUZiSLazZSc6t82ubq+61DNg6Ht9UhSkiSnFBSye654wbNE5l3gJmbD8D/
XS/+HpreAlbwAMdy984KKzoOHbpxU2NneQc+lE26PQc7BVCJ0+p5mGtu28WYM+kY
KNHVzOegK/6anIpptyPWZLWFQlFmHVZYKsE2/0GLGzzrGn0WiP6x2hcMtcyzXNa0
IBM45hY1vj+GPAygEtA3iPMDe+Xx2YspcoMtqWThla5K9yxFsmXou3lDOGfBtPHJ
tdCiIATwrJA32KLG6DdhQRS4jKqu1cOxJkT9ILZfHEWNx1kSFbzui7jy82IvAbtV
UTCMl5u+nsJI4/ZbKChDP8OaTaaNaOSi81nFujrcHCA5uJgJ1IVV8lnWXXfIh7We
Fq04qR3UakgUYF0+AkkDraTvhZog6uTPv34GHmk1i78dHlAYKOHtIjw/JjNybmrR
jZtxmFEzcjfYTfmz/MpSWB/SbKCM22+NNJGwC5NFy7iEEHgFIVTl5HF6fvE4Il9V
xDrgYrxTBnOMtY4FRuL4Tyd4U0I7M/jFZO3bqIHnc++zOnp98yjDgX/ySsno/pdP
K6XGuA4Sh1f5hfBEYAKf+sx6m2faMwd/zfbxNZHoc2B9xMouzAd6BMiWg4phGngQ
viYH1olpOG6HTr0cHvtMzwBTmlW6wpd3e4rekCT3BPcTWzmcc0s2Z3ApATKNhAhG
8aUb2jsxGCTszYbcBgHbo89L56nM9eb+d/B9bw+YwIp1vqnK+NBdQ/RBwvgS41uA
atIbltWFqVv9j63bUlcimQk+8lQZ6l7qKMl5oS9CbLrH0N6OTtO1quzYokDvB0FN
NYQ3qI5wYrwMBmQNreuQ1J8B92IPm0EQRh4dNBF8CL3zfnRztWNBV07cRDS8gpgK
bHy0j+TSoGlCeFxrdtdeyoexv098Z1GYPteiGIPG2Q1Swe5BC53oQL/oQ7mghLT+
IrirSYVXuRSwP+Drc2RUbg==
`protect END_PROTECTED
