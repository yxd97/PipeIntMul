`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N31XAtwJc0JTq5JVaIk4ve2EJT90K/kSdUleLpQVEaLHCpDjSeSpPFyNxIqenqmU
zjbhRRLjK8xUXZtSVwNC/eC9YLZqdk02PNcXNYC308/nR7eiZ521n0b6gpt/T4Jl
dgbJRxOdePuhg7eGxfTSvuvVX2BREnHKIhFuIsdfcMCSldY3lLaFc8oMW+2Zcgv5
AjLfgkqVNeoL+9EMwWmzdo5qBReegS8ci6TswDi4HBksacyhxIH5wcSby3n85+9C
5ffrigWctAOqs0oKW9aRSSEHo23EhXh1O+Ov2wc8+KEU6I+7qvqvdJWcfm6pz+BL
`protect END_PROTECTED
