`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6UxXgucssXo6l/sUadoOEqn1Q3ItOZo0NQQwnmLtbF8J3NBFNq1eYtirHBxk3aKG
95V9hPgeeJxTU6e43EjgDI2yOVQD3htHZjPA2zTjYn67KhFrASBNVMCh5hri7XO0
r9aRvtNPTnrpGXSvLPnQhpnNoSPDm9Z60tTSirwH9IjVuIW5QOgSYpmHHEVuQBwn
PUh7Lza9b3oc2+xsO92zR5cZAtRBOpIMTIGHCJXBREVyUZxyv9SVWD+6Vm1ibzql
8vaIEykFSK3Ki2s09TSV7qdpdeEYxoUvwecKNtQc9CFx6gMYi1j69Oy1o5/2z/IP
n/HavSrjfb6KXGHLdCWlIZDZBTBhnkRp6nD8STX4vveESKGYumCTh7sJKoRKJRCS
issPav4IV7D/EAn0IzVddjdav6Q46zcoyoXDcYsx3gQMRg/IgSAmcZ+AOA1MTFxu
ch4jqynjopNtuatW1pEFxjBLukphUXrs2NgUb4ofePx6lJfRHh4hqwaXtktTm+Jb
3WOWxMzk/oWXKHJIkEwklGW0n8qpDlHmrwlqpIapAAtCifwWXfLSBX20uVkzQ5c7
Z+lC5ywERMDNXf1I/5W5s/vOs36pAXSnKjRkkQEra+wreIk36FYwUVCv8GoKt5Jz
qOPPQlgIWdBYm/9GWj58YjbgAb2S91eL00i2MYZbsGsON/UbEu19UGL03Gyjr1y6
kd/folwx82B6OW3wQd9nu4gWYYMxFKIsCCYxZe9CFOWBpzNAtVtOYOn7X5P+sX1L
uS++yLhwUf05i7f/nSCBr9RNlfhW8J0bF78gzvs3MXsBF02lywzUDiOMUimWs3TB
P0a05Z3bejnDYHEaR4ci0CSVc3x6ikv1TBwYN1vbQkftDJ/8lQeMdIy+LbeUjm7W
uxMZAaykmofOz1yW05ZWvsuhM1BKTF/afkuch9FHHxjrA80cS3pGwvb9AYJ/mkbZ
EUwIXkgTuGXTjZW18558/wIxmzlR4+Rb2uoG6E8A8V0FIYMbVoMi1I+N6HdafPuX
8jNtpeYDYBSEonZmR0FHmi7e9iJ713sE+AQHZaW5FH08ivp8V6LZA7SpZ0S6L7cL
MtG63EMuA6yd6F7t6rki/F6BrDQt6uHkXlmlzhsj0RZsbZeVTtr8rQG3Z3Rqmolm
BbzEOZb+u5xSTpDjJtvrs3GUuy/5cjogEJZ2D07wtI/C/hQEgtBuDAE1tRxzBCXM
uu1R2T3bhKgklaB7BbN2/pCBOLuyqhTTCU2LD+igetnRvds7Z85nc9CuRcqDNo9K
`protect END_PROTECTED
