`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i+HOU7Z3vBhGrGw3lOBtZKQhK5TxC8zNERZ59rykxteKYAaKAYMTRp/4f7hDQhya
G+y4hVw6lzqqSbWvwr0MCqj4btL0QWf9moRWdyQXkBJnqanwoeemyeWvpAgLsWe1
00rm5NliYpnJQFOMPeiZd5Ym1fsXQD9w3imT40RRRkIvoQbeU1rmZBQBiaueWrZV
CFC18OuoUaMBN5dFWOuP1E0Z3CydZjd8VuC2rpOlbmxmJGuHjhVgg4Ny/cnsDmpx
gXYkQTnhXnOFoHkrCfeLIQ==
`protect END_PROTECTED
