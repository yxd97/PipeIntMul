`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8CcW+Oi5Sbja1nYVpKrt9d4X7pFCRfETMcc/bu+beVZSm1EM/M39G1Y8otFzTPRF
psRKSlM6fcTKmh3xRzblujkev8MUU09sPQ1jCQLHLtxD0gpVw3+kvXhJbb1YDWW/
/5mLmk77soEXDEOMreusyWCd4xD2CwWy/B8YUB4Et3NruiIMxKXiQ4BKe3Se8UGf
H4vur1a7y44nmz8UCG0VuUNZG99r45bRXaKmojEbVppYgUt3/0ht6YNiDv3eCuLT
5LDkcHKLPhzIjyIuA35vUgJL9cXmO2lqT1fBbtew/EI=
`protect END_PROTECTED
