`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tbnbnCwGXhEs2owZTmiqMUk0goDR8R2NCzC+ediNif2iekPwx4Ji2v7InKVQpHx+
ECpEY1qfpjVEnnBAmNZD/NwIFmBQJqzDgurK5Ss1bT+xXJ2aha+vyBFEU0Amk5DI
avFyYUZL8LpaX3aGfxcdJjG9NxHcgTVAEibK5+SFSEoyRDY2Ha80GRWC9FHAhViZ
SneMTlhUk5QiIcieUv2mOvTkOMD1vXdnoJJKRQ5f6lMcM6kcHvEMAcPOcIF6FkzD
1S2J9EBY6tlaXN5oK9FkgA==
`protect END_PROTECTED
