`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+4B4hDKd4jMAweK2vPfNEOPbshBiDH+hBcmB1zwWk4j8VywAA4Ok3449uLKS0UHr
mtyXQfjCSX6VnuIH4aSPWjm8PmuBv9+uYzihgUJKvFi4VX+m7D3yOzfl9tqU6Dtc
jnXRUMMeHnypkA8B4CZPibvhVWqsxycRYa0wc5DtqHjw485SxhU0xuCtbnKP6cpn
FzjJOFQYZkkwgMXUevtfm9nMnj7Io7r8f58XPV7HxHBrstkoxtiOIAfBqXi0rzZs
wpPcTXoOLhHx2nKVjvtnClRvbqDoV5GhTEq6u+nCbphsLQcm8WFqtFV7Sg/xea+3
6o8yDTeMedOjP/Jzu9H/zDNfB2o75JIZ8wvRtTwXFD/w1vmWsa8F1s8r5QRsKNlz
WaNXr+RyACJE/bxkT+O3mevfFbcmiHzCiumsvmGZtj42x3CyzHvQA1mt1M+uRoza
z94lkPlKaK91e1rqT3Y1o1p0O09y2uf24rvLbIy+8/mchuIf0/3uf//olJS24oHB
R4TCo9BOkonf5ycYqpvwDZ2CxIusmlYpbP8LnBvy0ChphgKhiQy6U5YnNRZCRAgV
ZYnmBs7WzN+cDjNLfX7f8Wbnwcw4ulv70HcKokA4Hk2gl9IHVeugnYo9p7yu25VB
+U53knoMcWOARB8FntGpnBGePZiLtJi3/ycccYtpvUXwMM3ke1YA6b0gyl+XKFHW
eDmqOy/7JXxk/WWZIpIu6zXiXdF/w35+xuqz9RBI9L+t/mBXgV/SfLDaLCxRZ1d2
f4EOPh77gq/CARBMKI8uw8bymYurvvBBK6J3xI16OV2gyG5bPOcmY38lyUr8WYIL
R1+t6WSGrfaxPaGpaurDrYb9UJnbeTuLm/pkmxCqrwZvLYRTL/T+SX4ZgP/FJPF8
3vPqI2qpPLKBpqhDryH+K0mRnzE6IHOvGwY6cB/nSdhSGhmGqkZcEASU0eypwvoP
EtQSsO4xXQPolU1YiXpm1kjSfgU6inBCaeBkoFAtpHb9EPo3QeriXsVxppfRGhNz
EVUiTcU3Y9uSKIvWWaLTRR/dBkbpPMrgaa+XI8Gg0N/PdyOMGh3840l5Bn8N+7Me
WBUMRxnRlP5m57/eSNaghERODEsMTkyiZ5odMDJC+5pstF4Ky6xp3CyrqwgZDPDY
OJ6uq7iXw2bdlIXoAsHItVKj9QkmSluc1WokdChhJ0EEHIyjj9yhSWjXrMF2ydc2
XdgebqBOv1g/OHmVneBO2WhOR9tK+MEJm1c1DtfaTrls3Dd2woKB2zMK2iofIUho
AGkaHC9JyoiFL9Nze6qRpEN4IzYPyIvPDICYsgyizEgBrR4TqsF3NZ1I0CYW/tx4
7T7qzQuN22u3jaBjAbikci5MBSYybg8nnT5hyrad9Q7cN4E/+k0HjgbakGfSs1RO
q8P5eMp8mAWVR9wS7cRjgVWJEIagMcBADyU3JTdOzxyitmAfvgt+2M9F/j/C1Djj
4CWPbiWg+aResEm2Dd3cPTGSjktUciBkcHqbZuqf06Nle644DgU+q91yDUT/ycUX
Z5Efe8bwTFgo+coL+WAb7QpzEwEFw7+l5+gmSGdmZ9mSOvzFP0s0Fgw19PxUc11a
V0VaQJcnOSyubva2C+4hAwdTPXLfqLX4FeepxzRzeWnyBZTFxehgUjDX8hbLbJqv
HTGdzmxgWpDZbzpXV3CuPsT52wIXbapb3LBFrRi+2nOzXEz2eTGkjWqfvWQHWpgl
ik2g1+oSDVyjm2/MR7Uf7Lf2ymBajp8KcVR8p3/uBjL2OULFPlFnyMviEkHMlU6D
gU4rx39i8OxdNy3qOJVCT0eOZptBK5o1vrv/khZ/ANrsu1wI0+yVDHs7jF334hYo
u9lSA6L21CBdcmChih+LOzERKrOAv2RenEn8pYLzCNHTxUD6c5WA8EJG4KaHIXam
0VtOJyZ+kFFGNl+6KGK9nc04dZJJ3IAwn9A/5gma1ltVudqpIKyjdY5uh7oxZOsj
z0eLa9svpPqQtk/AhExy/9HMLlSztvdH+1kdp/T2Duar4XIaPBxlbbS4VROMX8I0
pdLptNoa4Lmn+s1/x3ukt+qMdVT5v7Oy0KiYl1cq1JHvp9R+9einmaBEiVrtfSig
XrwH+v62FBPQdpY6nMndXN2310qY//1d2FiinvVf97utj5GqBQU2GYS0ebqX9VUS
j4T/ATzAdWWrKMOnMTMAJwAke7xjDGjWB2WCuF76QEaEWj6fFgI7K2vSADxptfMz
h0x3BWu/67KkcQ/qN6o8eXC8SWXbTrBOcYVLEuMLmcyo8+xgqinjc1iYiaa72iN7
`protect END_PROTECTED
