`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ahRMFPr3PMAgLsF67uoICioXne8PFuTewP0lGukxJ2nNtlZOp3p0KO34Bs6TPhjx
Z69CsufgoXurYDcDDMNvG/5wiQMq8/t0dkpMF7v2ei7RoZe+VtRt4eBdpRdpWWi6
GMTLvELsHyvlIlDGOLKZmV0E7C4oWg4HgAYTSrEemy0JPHj5wh/uIC2yU1Ee+DBg
et7PkCLc136Ogs7HnIEficAeUZ+JB0O5BPIvylq408JuzJGeuGUDP6tNgCZV2Lkv
Q4AlUnGikPPs3wUqNTeIjj9hhv28gAUHB5nU2KN1nZzYGGqV6ZEcnnLDOhl2cdXb
QOE1h+dS5HfvEw/6NRZZ0Q6AqOyvZdkHY9IbW20zcWdIPsXwmKSH9Xf4T+yG23jO
mCmNhIiihhWdKTNzAGQ1YMckfkgtpnxYHA93xliGt6l/0tjY17GuT2X2eE/EX/Su
XIG2zM6ZkHavbI4smwNSsNNZJPICdmramAFTHPIPOYjI26d2veht1h2WzxKWUJ8m
0w2Xp3Y9JGEse4eYWwnF6PIyEzRdY5MS5O8DKUIK26kJf5xKq4JiC/ruA5joe6yk
ZiiHdyxz9DUK68wE4b7PykkloOTnJibUtS/HCx8/paQv+vjK5RqAubSSpTLMlD/A
LwR4rboCMgtxx1oJTauw/mlneb/C3Wr+akDDWWOF98o=
`protect END_PROTECTED
