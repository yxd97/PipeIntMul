`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qpkkLsaGkj7Tb4Tqz70bC6tMvRVfZ90era9BTllqmtTjqVbiFP6rQhyKMmOv/7qj
mpjVSxcZr7vBtOXiWlgz6ONjygI6h0lBbrnowBMKsz+AFOh9tz38NMlr9oEYvp2w
8aXlGfBhdNBQM9XsEmqUl0b+PuiJFIrm1DPqRsLffYNgRxy9IY2NSNZMZfpN5De3
8fobaB6Nl3UiJpAgFhYrEMcRgSfm83mwRX0U7mCf54eSYW/a8CkQqQIFOi2J+ZhD
M55X0gz5G7kXV/rhNPJfN308tFpldhPDGV3n2b4OsUTWwOJABZPwUDaGxhkHXHLf
OBbIg+yfXKq05IiIVdzQKgNTFGZ12zkTVbEk0tPTlQ8oQo6QX8zCtOv3yzYnCXzB
GLYR5KjYTRMyBi6U8UI4u65DcfgZgpea0qv9PmC0vQaduQs1xhy201ZrpN3T3Wwn
gfH7qNgzNwp7Ix2SL8BUE1TE3zqeJMLUZwQCNX/3hOI1sbY+DMRkEm9eVGPMsS1h
lB1M1I75a62Cul7Hk7Ameq1ETBpDE4BH+Up4KCffGUaMp0ZHQd4ZbaCdRL1B5ABR
tsFyProGf83CzDiG9mMCAuaSNZYWm7xAeqWbaPMv42EunYgsX9L3zc/4ZKa29MdS
IS2Q+m+FbJ1std4Vi6hoE0YLVsBMVt0gzaVcF0JEsJPSOYa+e91U7Msg3NyFzN2D
Js5W0ZL/rRn5d56HQjHFYngYdecc81P0OA1tRuCThIcC0u7FcfUcWipNf3Dz5nfD
Zo8zwfzcew8YZY8qH0P7IlIdAu62elBjAsKUqigGvXg3VwOF3j1jYawZDWyHeGeZ
QUCUgv0PVzg7yWRIbWdhhtD8OoTvvdUPxnlhgfDFPYk=
`protect END_PROTECTED
