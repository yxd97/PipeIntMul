`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+3eLOeM8nMTA7sfPJyR+Pfgh6nYZxYRWApnqKe7zhUKYt/zpnh9ydnWd29oe9T8o
oxsCK9pLGGWjsT24Tt8t28B3ZzvocU9d/etp88GdUDqh2CMMmpMf9BJEAo60fFhi
pe6IrXbFcAExgGzJxkKwhgWqcZheiUkNJxKgQhWYiprB4K3bCO6Oj8+G9duy035E
dPFJE3pVOKLKKY4PnixSPAC8H37s8kJaooJ1mg23zXuQfsCk6WswqPv6nsczNHU5
MuGCgIo2XVbsVT2Z2shnVIuO3vRrGX96mmRLyGC9x31z08gvxtq/Nyqxw4foCTob
HkUrhN3bkyq9QJHDqbOYIg==
`protect END_PROTECTED
