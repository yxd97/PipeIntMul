`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jQtS8neLHCUmaJwjuDKc6e73I7Z6kodU+TBDUyCbQ5tggrj1V+EZHSFfxelN7O0J
XjLvdPgQ2tECDPa43ua34cogktHd1Qlsg/47wxm5DcH4ft3RH2obfmXbh2J0oM8v
zbzg0+caX3mMnO9JkEwRVn8E5tyG0xfhqkoq/G2PDklhU0ug7/Ya/3Bhs4IlNhwm
KAq1dijpG4hye+Pl+FwDph6rqC1/9ZwzFKT+DwnMEXEqjPcAj2Ib7EKev3JUP0Cp
XiHgMtuWT8yoaG7HbFake5QeV+DSTbm74k0buz0DQBX5A7RhBueKErnheekxw3n4
as4T3QPXO0lXsM/76Wx+wnG3ljmjqf/bxMIWaHmfrN6wHIqQ/GS0NnGSLnuwpPjH
ctvCOz32zO5yQ2NBlaAFBna2pYVEddTgXFnvAcdjTD/cq+m3ekgwUa4iWD42IUeN
ul4jEX0l0n20Pibo/ZQlZvTT+cxRQc2fM7jVnM21vvHWiOyfHX6t8br85myqCWGM
hHBelDsQMxdNx+gheOeZ9mBfYAaYGRRKGzUwZ6jDYx9YjUxm8k4NpZgF7gIVfHOE
/gEJzpYR96cYz0b9w2QEJhjc187qvsY/uXXKaDe8NA1ZyY2YBeOiZ1qEVmK6ucfI
OZWkpT/XrjumKcYTUHhBI8cuaIdxMb/od/cveOFOXuKgcShH2cq1BHPQLx+jZTFR
/zxE4ZFjJ3MA2SCzrJToBf2pI2EQ88GCYf8PsSsJsrj57x6yuRhYyWQ8NFCAv5UW
uAnwhgAzbrOhBwOTnNUIzl4R8hDNvUlNIaVA9mSUQ0w+wzuq9iI19AEOSOvlOBRr
/N7IIAhyAgli5XLoHbKNGW64MhKuRk74K+iAOeO15aiRtQkVW5Wz2K2hCrEvkoqO
Sj6ukqA00ZklviRIsRUsV70bYu4xrm5LWMhKe9rnmro/i+oyKYXeXGsbvhcEyvHZ
21JmxFhikhAwU+HjNn2hJRDDB/JawoqDLCFAU5U0pNKddsCrICy46MF+XXDqEftv
51/V3vT4Fgt8HykcHyC4rjynqfIXO1Orq/FBOFHoQchvMJlRmOdLLBRbnXB8/rGH
iHATaAQ+RQOA5BaOhZUG4ITTsp0SZxTpx1kge0MNxcAeiVfMNM/03eHYwIvfuXi7
N7yBpOWHvWRZw4yvM9Jg14o7Q9nd0qiokfSCUK8/HBSfQ3Qo7e6Cb80Bh1frrXeB
WT9hTvtfHZ4TiPf+mTDo5MVN5+qGyHFZYHujtywXtMYUJi0rJ4OThaUGmwzjgfHa
Ue2buOpl6vlv/L+aa1u/vMPg3i00eFF1GDgF2VYdh2BLqHtQnaBWxMMB/GD2mbRC
VdNd3IGdK9s8Hr8b0D6DN4PyYrE+wammKsiiJas2d9UKkBykcgGf0zpKf9MNJPv6
iLPjYQRsRyRX3Uzec8DBEr+kOz4jjtLeS76oEqHHUpOgaNHEvK4LHvF50uiDw18Z
89RkJTWw0oBVs5GiXMNiNVBkG9jrevumbCeQ+Q4EyCBUK4v1xVILcQbbedWtwehy
WfVsR1JGJod9CyDFppalLHoAdFIdsMUayUsn62MzOo/Ndd9tUVQK5j/T+jkIQHJt
Wh/tUNUsPXNxseSMN/MStZ3wTWptodAFjWfnPWzyGVyFpZbpDEkPMYp4sue+1ec3
PTdwJShSarfsvGDlUw+gyvNzeo1hl3rSP3RXN+f2J4Mchxsmpqv4SkmEeyavsu6I
ow2SmnrGhybYXb3aXbJVBbvBmeSf07owUPLidYt4Xx+HKJEHT7A8k7UAAZd8fdr6
AvP4YEYekH42fqgmqtnRL4VxgkXfb4i+f+khwsVlH9ul7OE2JkouCLQJ+uKNFwie
H8zmmytWDXfFgG53MrRTugm/MSwC0KCZc9jEhuhwShHKbuWySfQ2uev7DTOuF+ui
5h+GH+jfGDFGgmiq1lCMux9Vp4h02DBEDDvsgyfKej7PoShUNu6P42g7fvHGo1Qm
RFgUKFUiFUPhpJuB/JN59101gpY+fD6Vy/SKC8OP+OwEPoTVD4bELaVigJFbEbth
rG8viuBtieLJz5asee4fbioEGdwULqifF8xP/rSwWF2hs2nIHy4H1UVFuZNllMmQ
pW26x413hDox5lAJ5xzd57GTQlIuVkv0oi5rwMUpXqbggcnlETDe/PHGpoDuoLmQ
V6ThuKlekuHR7L3LixdguX5/d/ndsLySLGKwcoBsgvinyNZKs35rLF6jkhsuoUNy
PgiiAOqHk30ZGZDKa0BhoWwz1TIzOtfZW99QtLMxJZDzwo77SQQ/1Ad4RpZfiok3
sfsYgdCSSR23PU8V/kqf0dtA60Gf2+fECqVd+1mb6WzHntnh0/niW3NQ1ioIzLl8
CdYDkAokSbXBNrNbJO1TySC7vQ7tHKSYkOhf81eob/3e3SGJ08m51KQOJtONXKiK
NhsYczB5PS7GJUK7YXQVNn1NcJMmJP2Q7uJRNSOOrnpoNQYVCbswNgJqYxm0t2nd
yInz2+B5ygH5whOtqnL6IsF3UdGc0NtS7WlfIG77erpg0XUNAPpT/H72VhtfZfwE
H/m/8AgWjykgc4cbBatxSJr0JhZIaPTeL+F1Xz7TJqGS4ssq4ldI0Vp7boDrb4jb
rtqXwIqSP4SLGWFh6pPwV76gE/FEY9B5ob9geuDBVG2UltTjoGXDxANh+3dlp4zD
xePg+dGhQBJp3NWKuI/gwO3+vjPbHRkFz5Wg4tnVRq5vRF1Mu5T+kGEJSqvRJ5ft
uPf1K8dYcG+aGrI1ny8LDIn9Va0q9S9cDMQI5ybFsxcr0VzxLAfdjYxMdR4K5qT5
D2maPYYhOIwMp8SEUeOFATf/F+8bjVVb81Q/rRtGQVtoid/0/hXevtjr51chsCo5
gmL03dfomcKEpqj0TpQymXoYnvmA/Eld1rbxM0E4INybMNbqDMPgsDDIfIVqeOUO
I4wB3aSm7Lf35G27j4AJIHE5E1qErIsRSsB94MOzARjXkW75M8+TA+0FOHc5zwQe
bPNBkK13b3UcbftA4ios9zhW5DNF0Ygw2ZDjzN4vfhtrQi3gmxcwk0qWkbu5OZlP
w6Au3KIf8h8+X6nUJRwfHhzm7bI/yz5LcRUjg7OjTV0EvvcH07LLFHdyLtNbJo91
w8pV0iKIVrcB5uv/w02u9YYIc4Si2S3YIw5xRALAbnOwURke2sJsFpHIZPeab3ac
deWR154hR3VBlF75i4QVvxhF0ZUrt1v3YGzzDA0EOWdJuu7Xqp7jhuRxeLrzNUAC
4Ak/fazLCOaLJDdn7qgZb8NtpQ2K1J+o1s90QqXJMF/12JfDUguo50n+nIdyNJzs
FXD3US/gp6P+ttKry8KWFjp3CRY/cxSx618zc4ERRzZehRQTiACRM9kzzDI+x3/U
5+xmEAatuSrnwXRop8GqlvJpm7CJZuuDIvUOX4SvsirDrvgxzqmebWUmBeWnBtCe
zwKiK6FqiHHpTKtQim2MFfZX4s6QCHoI4nikXC3nAbxJ5FZF6Ku69urO6NDLjqPg
5ND+JGiyfDqCEbi31zb0Q8bx8a3lI1sYrFdGvQvscFolyxSwILs9SJo7T4lhZXfk
2QCtBNURQXSmZI8h7dnSeg8kY+oSTHMJ1bDfTmygbdORGYnrQNEDMdyRWIL4FM5l
RCaJQFR1wXeEEAW8iOzAbrsgm5alElgTy4OVe5C7KZSY6/b94tUJmH+1CiBweu29
sgWayIiLvmLjksNIqR0YFoQJR9NfPe1xgyraYFLT+46F/1iwV+vckrJny9HtKusB
Orp2jMObSt7dL8pzVB4uersftljXN1qg87rNMMJY+rmmtPrvAgNgCcEpbrEURCWO
kB/vCD6lfUtfKPZQkNC227ox3SK843j4vIz/yQjYBXKMgTLCfDN6PpoqmNMh8wD+
/w4MYfaaQCMSYVGLNSzJQxFK9OSKmr+Bjdohv8AyI+XLU+8ZtLJ0Tgx5WqIaJ1lW
/HoOyi+eW2l920dyDZG0Wg==
`protect END_PROTECTED
