`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o7OVy7Esb6OZMmWxkLwUxap3p2fwQggLwnYelnyQDp++oIXSp3Hvp6RltvVGWgDA
I/VyzBWoYxLWaQtvMatxhsHR4dhaQlLeIO9CXVrU1ujawxcae0W7YBYkVyNbuLge
mzEHXap8PB8ZtA55ZHi7AdKexsy9EYGC0c+qicTlCkT36XUHd6pFzQs8MHJDoZ1J
AlcTFmh2InnlCkWiA+qMZBIvRKAzNINKqR3U5J9j6LyPfaoDHZFWRbU7evndWnNF
PGml6hIGeX1Aq08oImVDrPAxJ/My+zK1rdVNvyzVgyRnSa8fEoFWQZKF1Tm6UDgf
FXVX9fWUPpW0fHtArku+Jhud+fCWE87FvXcCgeYcF3aERvk0LlU6ODm7vQ5Bnp66
8AanHH6qiernQM8HVhIZpw==
`protect END_PROTECTED
