`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mCQa+rjHHg6zBJWVGiRarw17JO+/gWFjAwpcuXUV1lgbfkDL2zXutDPn4uOw5TbS
rmiYwmo7yDYcdFFAMt7jL+OnP+VaQ+qiJtPBR9dSYzIt95c39eOudCCGdxFeKgyH
hpeMtNyEGYpAzyWCdAZsGmj37aXXP1hjhSu30i0VJnOyZCbo0ylrzHyUEukinZ88
OPQbHt1+fU+cy5Qb+a27WcRl78GBZ9gFPxBL71ieTnAvoEaN7/kAgCMxlTVyP/2c
CRsdIgjLtQUXk62MX16nmX0fEiE96WpSEg6PLf7yLBQMcxYg+FNsjBgJZ6Mplt92
BkJ1LkqzSIp4GZb+MYOi1KKaE6xC1dm2a01xIxKEjmB3bAlLvfHiqc2g0M1aYdUm
WDXAC40OnW6alffko0FEm27IR3dGDcXrD+9rOX0VPD4=
`protect END_PROTECTED
