`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1+bRxbvGq2rZ0A+3GamR4NvDvpTWYxiVVTUVVO7O2UcmXmAX6atYLIUQ3yyYSk93
nH1NsOZjY3jCcFNc0BrynYebOPXfY6It/gmr2pxYAmaAFnWRCRFbuwTEzjYSj1F3
xgZpyDC2Htwf5016vGT4Ffw6EPPeMApWV9JtjepYimWySIM2QK672xAjYWwzCqWC
E3oyJBTeFB7TNQhPGJlDUOpmGW8uKdPuVuKXwHBuoFu19/rj4uVpF7KFCFpW57j4
AoBRKzUgdG59AMUM+ZikMpLQM7dHFigvPdl9Y4Q5MOJGqiEVgCRHitvBvKZO3Qos
m9NmZgeaFd5aHImroAWW/6W+mOEblAShCLtAKR3qOURuxA9ACraASY+p+hhaUrUg
1aILXaUr4Szti5RusCtvwQ==
`protect END_PROTECTED
