`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8rCD9tmUb5FkfRRneEO8o42DY67Gv0IIzMoshyznHMJ0+LwC9iBnl3CKrUJt83Fl
FRal45lOZ/rmsR/DwYDTjD9iVQtx++Cibo4WtZHZnWHPTCn/ZeZ1yaUyJU5fIU0B
x7o70p3EXXBocej1wuwrVLCSoLsW1YvvwTdGbcXAQBgmoxtFBx0UmuFPLGOEg1G2
5XuvgyfD0YZGAeIYIvadNDIVYwkxW4Ipfeax7J7lMQqTjO6CRGykvIWSiT3/fOYG
ahP9XcugPCr3v1BE6Dpsx6mK0ebTba2QwMBJMICFk0KRiZl/Ke0b5jTsbe3IBywZ
/p8XM+i2uZ8CyfPbWn573KBG16rhafAyLpE0RIqzzcrMm+yxxxh+ZaY9gbMQlkaR
eNl07SmMsVN4O+/i1qfBVkvXqkoSoH+6xJqB+4N+rxtCvY0XUwEjvIfhZXrsz/VQ
XQy1uiyDP34hw/lPvfk7jdB8MjsDHm7fcJD5oHX5fT9ra3o4zM5PwmYwRO5p2TpQ
hcYaI6eBNDJaB9UgAPltmIKf7MDOASCfuCKPMRNFf27SV/VQ/HTJFt+b6gxpZDtV
2fDJs21l5bHLmwi0/LVowkjqdKJiAe3CYiTHBHezl3s2SEDjJ5DKhZy+pl4bHhx9
zl0XXS8XkMnxnLyQcyE4rUDzCs0Rb2OQalDr9V57bslhOgqHf4EnphvA8rR9U0uQ
vZ44zVKJUy72qNkVw8Q8fUutK6yQQqKbJ5e99XoBEybTjd9UOXmGDPUKoSesY8fY
v15lbJd1vnvhAR8pqYdxjaW+DKlXu3hTW+1gMRTXaYHGfV0wZspwxtPSzi0TiiYG
FkPnIshwTT32hf1AL91yhEfS2MMJ8T3Rre+8+19x8RbM04tYzs46xypF9wOV3hUF
cziS7+oBi6Fb5IHIO4PSi4y9oIes18qVlT0Ro7hH1LoKFK1ssav9U4IHH5uAQiDK
2miI3HicI6C5FO/EjGlm8JvbtWpWSRt/SN4UFhykjSZmUC9ZLiceswhqT0N2copK
80t9PwPo87wIbmQqG+lCE9QIiBGbaVXbeNz/1UJjxWsg0cdBnUgnI/wcuUtuVTAe
lH57mVRTgw0/kbWadmD5uti27Iz6iC2UnmM5aT6Wv0KAiv9/s/WA2vx7pzjzo1Ev
dpGs3wqR38RDp42h74ziXzW9ixsmKAUGg+UzJE8IQbJKBQMpSDrwBhdwugQMrIJA
SGWCFxcznW4mjCcYpj1qMUt+mTgU3zKLEWCncpOFXmpYUk1FT/EvmFO0cRIPMDcG
eoA8f1KpG3q2tPDbqlJ2FpyVZR/hBPh0gJ6TpS0RwPELUkzn39tbvEMz9Mn7gUC0
pY55RioM9MRuX/hjIdA2TznZTQTs4e/Fl8/cAPQCGQGqBxL+YbtF/ujMySk1LcLI
uZHtBd9l+qFLuru8xxo/cAPKK3s7xqrlnxLyF7t3cjghkdnCciZAy9MCVyJPDl88
gusBOFjS8AB58/LX/XKuKDf9U8hF1vXxa3JmwocK2yQy+17vzFltiuR01UFEDn34
2/+Chezvf97Z9txf1RQix4i0wKRnTstySzZJGcu5VO9C6ZiJkaR+6UrZvOVHtFW7
7uFm/8OJO0KAEX+2R5AfcqEzB8q+7Ll73nWi7YK+4Mx/GsE9bvdHR7DDaeCor9tc
FeHI0wgWmgNnsbXlTaSYsELKOyUl1QN9ck08i3DcUTVECEEKFuEM1z36PeMnOwUa
d7fprHLyLoTvxryxAb+VdmTiJVJHaZA8V4gp6nM2P+8fcFScGE1cJZ8x3o9Tx/7m
vCkgL4cc7PA9KCDJjkKMkZOHaCjd6ZnNznymXHDmA+Yls+VrId5n890RuuM8P3L5
4PyM+UTc467jNtaT2W4F9kzEHrPDDgoMuE3+qxX16UYtCynba6WTrU1r69rEhFxm
jI5NvRc3ObT1AbxXjGTdDVF2sWaWsDga8z3yngFqERopUkG32tR9F0J7MZInqA8z
umyhJL+QaI1Yc/Kv85rD/2xw9SGlq7UxSJG95SYkxdTOEcFFa+1xp8QACRG++Ntw
ImgCAdSVbveHogP0b5sPTWUNGuKuJ5wOQjP76jDiabSqukJx9gBZ49wEbQvJ8vdn
W56/QQ05GuqavQ3vkTwYY0oasIdAigdNQU/I9p0Cia3+QaZIAu0tPB23mDAnA+LT
XvEiwAYsgCQyHnIneq7BGBwmYV1zsdQBDLYDmSQX0PrKqhwZyb49X/A5NRIyiHfe
NtTcy8S0qRs7c3PmpWWn1js0Q43n7aEhLaFPEObodTK8ZJKiTgqHgJaaabkzCz+o
jJr5wQQ5mguH9zfXnk9ffQBsSnLoyrJ/RwHmGihc+xd2XoYr3G9ggxGk/RWYf1Y+
psHzrtX5X77gZIeYD5/03qbXX2Oln0N/iATfuPg5FIkO/WxIJDpEXj3SxCbNSWOL
uM1JeXOEchR41HCbm1jYsnoeKs2sM105bx41Br/fD6O/PTKT0qdXJ2wfKXPibauO
cXIJlsnz5kprOnqIYx9UpUjlvQXECeJW8XY200mtD42Er1yRevkUUtoBDDjrpO+2
FT2GT8YGbkFgCtuOfo439gJJOGieFQ6sR4u8WV6ZUs7yh1doa4z7UGd/u1V5WXKz
gr0e24zPlUQ4otOhg3rcy3zPJ9ZxVR9Y8a/k/dgeOJ2Bg7Tw4GHk5UVeVSjiAWSb
aQ0mYfH/jh6rg+iuLHvCY7XqXgoI/E5wdz876VHBX+aG646K7wBqhlTErw2GCCDM
TRaAw6tKNRrdFOoALp/lQnQANnCyAQzjEHHfbDwGzOdPIgu3HFSAavASAvkq+vMt
Is++mbrsRMS+TBn36R7ewKQbqpJkyVftGlBqow8AFlGX13sEqSsYtkwQr3AGkZJ6
ysk5n9KHfXh2b+CibyB2Uz8RdN18qHdC06g1ICp1+iyMY/kl/y6DRvC5TvBNmwy4
XS5oE/1iyM5IsFWSpQaSvV9YazbD+9WAOde+N8ey8yeLo5YVY4Lc3ETHZt1kSHCy
x8aDYORu6wjyVL4741F8LCadRfNj3WaQIwlloNHrgOYa8rPBqL1zQcbj8ERjWFCt
hgrgweYfmazmjjtgBC7pEE3glusclemsaJVONDKXF0dJs/udsh+D8CqH2x+W9gv1
QplJgvfQvzLGjdOdaiHcYF7LqhG8P4S50NsAe3bB+6gk1dB/XohsJkRzSeUJKSZ2
fD0IxeoVEnilSnc/re4OPTjpMr0bOVr8kF2AnTj/8UivEVC9xUWkvtd46n55mFMY
Ltb3+pS30AURXycheLgkcuSDy9gv3rkQaialtMC1vWXRt9xuyPQKq55awXAnxJKJ
C2GTVfARiyunpttu5hikQMFspdrYvLr4K3tX1QvkgsOD9Xv8kNb6rOlkH8r8ta3H
QL6mI4MFi3H64mYexKQWDmrwXfXR2KjMBsQ6vcuHR6MXwc82/bLskBsXwLiYOArr
lcg42X+BVqVLRzXBZ45EPpRnCzDiPFoa4gH0bRUwIjR1wMiKyL9vjRGRqFesIMQ7
cKIreVkcphEt2hIrwiryLky2Q1R4ON/492tvUH+NzgZfbM52DkDwwUCqGFgImlAG
9vAYpam0hlUD39nFa7/khiiwoyVqdp/yXnjD64SxI+t98Z2LAgYti3KdiqZAmJ7q
IL5SIta5n+9zE5C3lzKVZxYszWhO9uThg+6BAo41K75dMnkaxn1srhMmRbXm9zYQ
0q24FDjFejwSYVuSzL+Dba/1vor+Q2dsCG3T3OUgPaua6OSFv6fIEmHyDEEH+39f
q5QPutB6GLOQfGyhVXHoITrcKlLuSXUt12TamTgs2QKSoeiJW6J+QRyQpdV/qUu9
MGP8gYMv5oC2rTSqRyu1UBYFso3BbJSdk4hKzRG85dibLiIVXARB+s839P5zbmMR
PmoikRHVgBr8OiXZwjBA+017wLwqfo70ldeVigk2w29XIfUt8oDAfnOjsu/Ugime
3KYxMXMwM2JUXYKbv1k62JXXswdm96PJMK3OjGOp49Q4e25JSxHnN3ejO250pwDi
me5DlXtEiyiW3YWR+YxK18+3Td0m/ao8rE1VwUcNCbo2rjkgF1Cy8UI8oz9Q/rO7
KGwGFPMZ+zqcRQ5LgRQapCjELQbr9K3bYOVDeV2+JvxL9HcV6Yel7TrSdUPGSX7Z
/NIXv7dZLZI6x6jb7NVCISCjDEI0IrB0DTe+kiKqhR887N4NjZ+3Q7u/GEFKtVZW
ikKB6XGOr5wUF0tYl3QLR1TsSrR9Q5uUJcFS3ZIhD4yRYt8p4sEOvLEH9lFJIgSH
XGRooUwIL1rrflgpUXyy3LvPvXmoK8sXfd1VE89LgNwwQ9GJHs/U44DxpKGf9EqC
FsC7deehxpnUJV6vPk7V38fTR5FMJO+u0QMdVQiqojB6TmDF9WOZLrsZeDvfoT39
OHcTHvkYSpMaU/WAwVuGbit9wl12bOgTf7BliQN63c2K7oYRrB054SMHK5hc3TfQ
BxrVkON9JBeGIkI2l2AlHhEcy3pRNXR3MzFQt+qnnGL6oTpYpoYQjx2EaEmaj+uP
L4xZAs5fbcQYbn7RT1zX9vF5ETE4BjsvB3aGfWXWotFW1zjxce71FdIYJnwvJpKC
HpZrItuwoppE9+ZfI14HAB/j5UCJADO0XmMczeRMOfpBXF13slxDnw/M5VXb9Zjs
mllvVVtxcEyMZNS1L7yCflgLUWLCOiATCUJCJSOFMPz+BrjH72HHdecdI1re5YHy
AKrQ63JwMYGdzcH21ZYuW0dQWv3GkfJmEJOgE+TnM0IcggBoxfnT5nz2dMGbKFtn
I/AQfrvmRRsSCQBglnHTR5ZhKAREYjjO8c/KzDWqK62HKoYYSuAHJgRbE1G+6hYa
K1nLS/6iBIGRhWUfUgWIJWvtSZtMoQq/QcphjCci9k9XIQ0jHCM3OxuzjrlRCQxD
oAWFd0w8c7YDr6Ul9Ti+Njx1sJBI6knuMKPquMENpbLB8QrK/jPEIEzQa9buj7bJ
81VP1oQCK3iVKfN8bFBuMRAMK671m8F7m6j8+ODFZKpVw1hK1vRYlN2vQyvZVrF1
8B0eCuRRm7OgQCM0//Vysaxwo7y9Yyk4q6MPcOudvJQ0xPNPW4ffjbx11RTHWqnT
TbwcO345bDXThVrfPqVUzKkIUVIwjxxw9ZD4X667oWE12Cv0yTzv2+Oig8AnQMTo
uwFXbm5qrAC3u4eG3QR/eVmNcCSmQyYUSzIwZsK3PlhwUw8TRIRRBjPjwr2+vagE
IzTuH3WkKqCt95s/lRZuhVFDB/RzesjPiv2Hkew6zGBpdl5HCcLU6MtIavEivwyW
APPrc8QzEpNiIlwNJSl4MP0AYjsTnjV/Nv1qpVH9j2y+HEhOwepAz2uDayskyMDW
42Vr3ncIWKx6a1llylKEofUpVhuRPYWpSAen2qz1bMBvWqwuqLXgstOK7aUQ4bzc
tERVKhZVGSFKAG5FDqi/3j9tCcvvMrlzbFibUqibgohQpkSEhblYmCnFA56prTRe
zUP1a8OodkFszVIvXqFOd2XyzW+5CymUSjdOHJ6y2P3OppCt7zOt1JLoHrhOpJXU
HtZoyErIfaxeQ6nI3CpwWP274yml6Fb3UIYrG492dtvGqpbab3jrd8PjniicJwZ8
gKQP8yRd043DavNT1XYEkYEdpe8xikxhDZr14iBseCod5lNE64F/t4yZRQFqSKmO
fnipg79LBdqAXY9fELotO4MWJ9nFuv27Zq8C1IHei8A57rUDzFyMIJDaWtHuPXZ4
HhOXNH58mAIUQJ245wgmAA6wCCM6TDYETWzWqIWVHhJ7rtZYMbqb1UQ3LL/bDqKZ
eIlw6pG0wSM662+DPfXdc0aoPXiO9yvKbwZEIubXsL9uCR6kCK+Rn/S/nNKrm3R5
/au5D+SEfwcpuXoTpxvshkGTaM4yBjYxkq+7m8TzEeDiRVak4pt+g51MtR/T7d/m
uQQP9F2GIBjWCLvhQC1UKpexeY1s3bVhgb/uphUI65ZznpGz7dUhovJWMtJeKzZK
EfaPz3uxTFAuk+OChtUxa1QKnBH8Hgbpb5IKW6mUQYnrRzrT3PBlHvjb6pdf/s9N
tKsXKPZn1Pu+Cl+gO4S9LlUYhnFHFGTGyfrpedSgHVoTDlzDvDXWQgbG+POUHlMw
8/1p4pBICZnRKVKHMkoC7uwoN8/LnmYJgEozGogLe3OLM68GeH6bPFUhHGXvWSOb
g2PDwEsAMZGK91tD7fFsBOxb3CIxMamKOEujggDUv638kQdDFy9pBcHIz6A60qy2
35B0TdTUwakdqvuCcWM3rNbSFhJlTUn/iwZrLTrgSOBopqJmiaQu1PE5HJYECpgU
4uw8kSYNhkvAp0J5mrpXAOIhWy4P16F/ItdWjH1tkkDEXSPq2Dy1W01+M3DSbJFt
DkA5kX0CU3NMu+/yOg1PV9AP+Cn5FNn3L1jlQKGMGiBS4RZopVGrfQpVc9nc9xzq
6zQvp1tKnqYo7V1QxtsDIu6NlxkUZ4SIKiBYNfX4Yt8HoxHSk/a9XPm/x/40HjdO
ad9EGw3IfotSCZJK0gbA7Tlpj1GJ5s8a62bGGXOkNbQMkfXk1O0w9h6XkIIp3rSU
xs0QJGMsXZ9enYmR5nq3pOrL71eRQwtFAxtL/iXmuE6q+i2TLZMjcWGmQL66LSjA
P20RaYwVv4NpUkz5HlqAben6smwr9sbL4X6Ks7emkJO4u59LK3Yh0UcfDHPucTd4
LsHbRBavVDpiNxz7l8AXSf+YyY2RhBQsiq+P1ZMdDhZqsKvAgudkrrcxDjpQCbBL
3FoP2pyBRVuLO0x8/f38dtCtn0ipq4z5587eE1oY/YDvGBwNLWbattO/GoOKFaCX
uHWEi2ErumTZysQK87lgKWWvWLRveAXZmIvPQICbVuVZXqOAfhIR/V8TIDj5BCk0
wfAvSKF9E+MtbwY2pBLtWAR0dLGud8nu3PsXYDBmtHEeqFB8P/TbZ/wLn3ZUrEcj
zwL9+rSAy6j7Ox4NyR1y7NmkkoZ/yxkq802DBDPZHHVzRu6Rl8Wiz63oEQMmpCoe
EHP75PH+5nwAo0kdNgg8ARNDKoUs6cSDRRLCLtAgypo3MNgySqxJsidY0g6Y48ZP
Uj+WEnI+zRfatpY7xITK0rvyNDpfh6NU+WMOGML5QOQbylLQZDP7qmIBv3NF5Fdx
gOLrL99RziWEnEt8Khekv6IDcMKcD7/HF3Vv241O7lv4nnk0lKusVMMkM25uknCw
qgCex+NpUPY5lYn08uKzsx4WFG1JcjweBVml2qaARSm+IYA11vLTFf4ar6Z8jVwJ
3lhBj2XhyPhNC2aEGQnsvOlDYSyVh1ODPaGA6zf6q2+3D3tS7iTlBMBMy/cGTurM
fL7ma5uLWIxhaoSbhQdYxYu6FQ5Oh8qrkv8oerL3EpL4xEy2ZWGXhZDTyfCYkIdI
gedFlc1jBgJ8fI4sg3iWnc4xlqv7Jd71R7H+9nVYmH4xoSZxTuBId5+5nK1r4eya
Nv0oq3AXoW69XV+CCeAmLiBNnqueOQ8LqK3iPDzcBFr2PxENl7lF7lDUrSERUdwd
ooK6R3wRLld5bmbW6f55uLSTRui2I/fMB0aRSOwAM+p210GUxf560AUdLe+qL3YZ
nZQdkHsmf+l6BVxvsVZr8nT3VGQri2haVFVcSOz/1meo+rKP0OKx840IST0SYScL
8tLj2Ou5QEkifim940AAEu7k1M+PQyBvyggmBHWBMsaZW06UwJ3DPCbHoX8Q5sY+
BVCYxDZxCywUOAvzMaJTHDbFtQ4x/xAnZSpI0/sukIWmX/Tb9RyKSVbAM6kiAXEF
lslCyOV/W/OjVwGgwrvrNO1LTCL9cQ2y2fQu/f9/kQwy9250CR7H0DF007H0CD6h
fIeFJz6acYiPkUznV217lHpHf3w/8xRAqHT6Nxz0CgcksmjcadG+hOg49/7lW5FM
+i4Q9ZuqQBnmi1SzHhYPyVPrB49Txo4nKDU+mdBqsKrmsm2k1aa7heYIpfgKz2Lp
JTwINFi49ZZU3M+v5gjEmrCfj8LO4IZD1Cx1B54brrov93kyRvMNjRSE+/qSbLwI
td/YIk/1Zauk3UaLm2QsWamXmh6cYIEvMv+6SHXgWFACoJUyQH+GJJXahhIpfUtq
lq5HoqGXwm/fCI8EkAQY6DQLC1rtROIRqCiMDR7yuP8ACjrFGrlOaHr/edPySM6Y
jUpQLAGyZMNJongIaBY5ziqmVMwqgtYHsGT2zKQE+Y/LhuodY14vu9JBBcMdw20M
wp3jwNpvuvx5LS2PU+cNJxAvztS0M3E7sTLZfJwPZ6Mf9BiB7ljFkq2OJPo0YfFM
cAM+jPisOP1guIsS97uNO8CBNVezjKkLYL/NG4Dxq539xx1Cs83AiHluRwguSo4k
EqMVqPhGYi1vhPw5xVx1lMxt71Y23+/lcmpcKWkDNw4w4UYHQo21LHYBE7MAE2Ij
x3X/MLBgvSMEhcmOj+kgjg+JvRYXJ+hPmt0d/mszyEON3gL+MyCS58tCzTfllfQr
/nJNLV/6F7I3Uxp3eHSJqY9OYFvKFdl0LT/4zSrs/PKACSRhXsdptNrf3YFzohDE
CWM9EjdWitLivqRGC/Tt7sSimbnYKigJxGOxKMg4mGVPYfSamO/kXjgu98be4wi2
repPUFBcHYg9LdjZF7UxQgfpyDP80nw5VkLeBts6BeHbEqlkwUaSNEIYlEOg1Kbh
cKMu+gjaSDAMGTZ+bd398EcmEdvwrzwIXfxmZFsN7cmwdMV9/r1FhxKfn5NjVt3G
Cvy5CjecHkPnbjPeCWc19UzzV4gQ/z6vKVx7nZfzkyL/ZsJl1kt/tG3HCCRV9iX3
hFcxxcxy7lhG1vYo7B49bbwQMQN0bI2CzhAaqyNK0J4M9O8mskS6KXfACaxK9PHv
5emJUf8Q/ls5e1SFjrCHToOS8srFjojSns6o1yttz3u+XaWz0ycOqlXyWsV9xnHr
OW+EQNIQ/xuPMOc3a2+MSkvskQXZJgQIP4F+3tFIIXOwEc3GKhp2aqcris9TZuvx
LNniRdTaZqPqcouVFjnqs9mt6WtQxsgGdFUGr7SEtrB8pP90JmwRwe0u2JQHWwL1
pPXRYk44AlqX16B2e6mpUrA1pah9TAD/7RpAFweCyYUBL8Mnlckmhi3MaNBqLJLM
PJvRgUY9GAotKvEgZVY6xwAyIrE5d7GL9y9ZnTTzccMVswh+GUGXJfMKI5TM0P8h
/r1ORsjbKdIxYwVHWkGKaYtej1eI75I00tpTFtzlWlaoFh4D90Mxsxhttp6ev/Sm
VGgwvFL6qoaYpYGtoC5ZtOEnzFa3d0QzMlDH1kwIE43TNaS1CugLHuwW3Hoxn9iM
Xs1F5aVk1uEcBDCG8XIDYyVlzr0ekjhYBUIxnLbpOKl2klcJa31UUnTyZFAOrnQH
jPED9jcABbWtaFaaY6azmz+evRUnc/8RAlHQL8ECKJprtPicFeabQaZDMjPAGTP2
PK9mxzoMy7IfA/wUnwhXG3q0OTb56JxtjhfX6aJ+BH01q1wpmECpBnBTCPeQvAhp
UoEP83cT5QDXtSu2HeLB41cY+nVQLHej+ij4USJmFqcrQC+m3eXR3YyyTjITP87a
pD1xkrNuVCmySaWtSMr17WXGljuqyTzUkpLKdG9LxLsi/ByBNfZxRbFHrXFCbP2a
7Up9AsW6pSl9kTiX6b4y3pvnU4qaVZnfOqt0JK1UCOff10+/NMUgsdrhqw0b+Fw0
bym22efBkbUrPxNKz/ZCP6pEx405TmJ/l8FbTwb13BTqbyve0GZ3xn42jdlYM75X
KUJhIG29aHAtPU7oHBXYO/2X1FUQzrkCmqa0G51Qpz6SKHa9l2VXgAo8SrdrJkhw
bKx48vch6yWmHy/226OVcSzCT7BPK/a3B9LElEmixemiEn6RCiCOvA6QtiBb9PwJ
uR42UeQHM5VAyzX1XCSgxCxLx5yp1KLwKIw11Ud8l6+DaNZSi7LJftFSKc/GlK2b
op+TppICkFM9v9BX/HBg3LrHz27aCofzTivDazmoIBEO+HMc/egR9BZ62XntHmxB
bGlHIvcw2wGbfCwK1QzLAk7CWtHybYwTewtPvuT9zzlx9sEtFWHXPPlJeU6O5T96
OEjQ3r5IxttneGU5K5tg6FNLGquOOnlO8wYK4njz2gvHgG5nOFRccavgq79l3e8I
vqYKl511MCMOtRQ/FwJplZ9occFJMkOsnvf0Up8UIILxDqr93kocvQtUB1SU58SF
ayHBeXLXrtWon88bMlKNYnvbMSqsjBujpBEyIPKSxDCVbwHoixKJpxgoAR24KDtV
hb/PKU65X8R0fwMyyBwGapDS6Pu40HWmT/2pmdl+xx5oDytSpRjMpNvLvMbfVOxt
jo4kQ8K3yOEQvkmWg0A8Xoj72LASHAidKERIygNE+bl+ROtkKcz6hVHFXCuCIWAJ
KDkeR3KS4d2eQbD0MpKxkyp2q53JyOLjHH5wMv7Ar06PkH1O71FxkKj9suCdrrK+
dDckRp1uy3B7go4zFrdUoNF+uhRvDAL1Cyg9esktCCvX+dtiR7G5TAbNBB9tNbao
/C+Q27uhGg07YmXxtOdvRxi07F/HYrymjTy8yac9cCAiIkmyi+jKoPPbe2Rcj5Rf
ZRaZ7rc2WZCNX5bgnyLf+Fb/iEArh9Pvlc0mrrwSvUKK8TFg6oNnxIkLlgZE3uBA
Tr384JwI1hbpSVs5BvJ1UJZN/c965smHkPR7+yq4wD7mQmzbXyTw3hANpTjFg9uk
cag00W61fwOFQ00SmB935mXPKyZcOTXQi3MNqba9RxUCJp/ikrKFv06MTueSnZ33
TefLW3NDMzm5mE8kiLFrqX7JHpxD0AFc403WY8zUx/+9g+74aRoFCM33tV6YXB+w
SDyo1w7VAKtzN5+Hh3hKNr9TanyjSlerX9m6JTvJ1HUZ4fOK3NV57Cs6xmqX9Nfu
gJIVUI72mKxel6c0Vo32ERLeJv4fRIf8bKWNuyfz1WKxtTRehyuniyVq8rWZ4uOn
k0LCeb1vDIKTW+GQ98Yy8+4j/mjMvJVzAJhljO6C+KQ5IIcNKTGVQBrH16L5CoGs
aGCOc52fkrK7FFcVpEDJHyqZdt876JZl1ppm86sJZCWcYaSeLAOuKy+qy9+n7IAX
eXjhonSylwi0Bvu9o+PULZsEHUBgZJwV3wzPfvAqTomf13BLXntHmhXmj0AWznMK
6w/qj1cPTuqGI4AOmpzFONphXp5383CgjDEkg/swR/LgCG0DOPJybilxCFXiavF6
i2gWwbdBH6hwL/Nl0o+FdO+PDIZX/ow5NEweSv7B3kA5vN+jfd13VKri7sks5KES
toxhuofXbkghUJxY8sMTzM4MWaW5/9Vyyyzy+lLEcZWi2SzI9SLb39lOaDU8M+V5
BCmpS86O2wHJ7+RUOGu+Vrm/7In/+ja1FqLzs1cuNSCUZgN3gi7Q0eayZoeX4QSt
YY2r2PtA7QgWmKPTgEMPw9jQkL2fHwrUGHnx8SuLgUaTPOHyBFACFfq3UzdRcprr
4lFFmNqS8pRSmKT0bJsHEQwQkER0tF1SSleO0KtEn1TmII9QQ/r0n3M4gs5QHGZF
93Ld9agtiMLqIefI2WlEycf9ds1CUxVcHC26wzZTDbC7jm1OZ1cgdW+y7ax2xSJC
CQ5xL7wavi69Z49giSZckhLAaXdqiV1ny1X231wOS6VUtPnEI1kcvJ77y94j1ayz
wd1jQUcoG1uEi+bBp43rOg9ezvzn2sQDKNenTp5sTwAZTEkOMmNtWDXKIogRGENR
igHNeOdy+rJwGbJXTguG7z5xWGJJxCymNw7G8hNLP4/IwQLg2RwU+WOto4Rcpc89
4KnynFqS5iOyVK+rGB5iKJKbKw0TvvHOM/5SjRMPj27xGGdvdIG4B1WT/ZGlwtPz
BniWXXCjs+V5KhpnpryBE5BWccwtAG12EXNyTwPwOobsltk2hcsGGcX4xfK/XI+N
JHLCSxYf/YmHpJGDxODtDiJhTVPSArLBvqurY8rVNJfzz3uCu2opbVFv/VhGH6JN
bLDxXubMuqXyjKfilY8vmJwh9YasIGofO5KNjlVXRVc/UjEx4xtpdA1xDkbCbExM
QcTfrYEJ+jc67vMGpq730fulhyOzCkmPM8MpecpHrI4s2A4/DdhwvcJONsugVVpM
k1R07bijhzbBhOwWjplUhpdhHIW1DTE7h9hTzFtk9X/H/UmvGYn6Yi3r9MHO9GkD
Jc+DaXCGY4IknKhkErBBai9P36IjYAOzzOvnF6FXIv1xlsGi1El6ptPCAaFRsV8z
i+OGO8UKAJxZw6cxo9mwFpjf1clKh9122gFC3zNrKnyZMi8DoloNbj8sFpxxdh7/
DvlYSv8YIDlRiOZdldp21ALB49utF14HXLNApTLSufoarpbBfSdgnQ8Xmy4VhnFG
c7L9K/FfxgkBwUNb83YCOu7q48oIdCIDHgivGNHgWskcY5+yLhfSj5cRa8Xs9WPF
nXcuw6rAjnVkEr+Wzg7zNnpKaL4i7wAC6zIbQ8LV+Eo4KIKEg1e5ZwqdwNPy4xOR
YEiEe8A39KhQgm6v59x/BGm7sq3cD/sMdIXLXm+PNXKJ7pUMRG+QKqLdRoI5Imr0
M7/NHigEYtGNFwlRcylDgGxOR+DqpC71KvRxwdBSoUIIkMRvzwE7jRAInDn/KgnJ
fesEkF2QSXq7wzedz9/TXWqwPPYsuM2ds2/wy/LXAlvgq7hhBUG+DP+HUbpGMbNa
B2f1LjxitV+8l8fqXD6H5t4KOJlocLOcLLprYpojqdTZD9HUOl4FapdtG14DutEm
KyeNR+mcuGLx1AII3sSyf+mrfPfWkCCVOhbbSRcZOoREIXoxGFgy9CqvD9lu7qob
4MAh+aRrnCX4ZK5skdtOVLI3wV+i7W2ZF2wo4GTjn7YlcudFJjDGc0RyKPc5ld1V
zQANQqN9M5slLAYdZu5sUj8ZIIlxULyF82o0aI74hVaO95kzvIVDLPDq0z7p0x/O
2ZkV+y4Wlc+urtQX91FG6lUxfwPc4IE0tL3H85phLkysROHsfWSxA52xX+AxsHLh
IdEw8isWkkNyA3jRHWs7+jM2H4Za1IptSh9JxH8lBXyZ1Yu4id+pg1HeUeMLhP2k
14APiggNGe6k6oLDAgtnrYqq4qi80mWSqqAsnVlEBO3k0padvjxPnYIU/hqhk4QH
S2/09Bt4GrWnfBpB8uhXJ1JCcpoeyyKz3+Ryhog9uHTOnzFXl5qy3WmYfno6zyKq
GM5z5emQhFwQ19m4SplVCYUpzoYDxU2GKx8Wi40n6BkSC+DoOOwueBw2VREwlHOO
EUnaBFsC07HZzUmSOwnzqVOrQJEZblLc2u5+249rmDTV39TWu2zdG3JEZLKwi3wo
1hN+pe0RL/qIwOHU3yTnneLGpDgUz57msuBo4ej6rc9aWSrmVmzOldObxkSw4fsw
4C1nkEs6xRvPtwvSQWUHPUxJ52guk+kqA90tQS3Zmv/3YTwAYMkepX1HmOHq66kj
rZrfhjXIz+fzLKgxOHUdNvBAQmrAbdZsj7qntWtn1LUZbUQUnqKlfeq2aC7oT2+s
Jqb/IBHdYrIJzWwC3MaLXq8q6lWaW02AXkip2iOmFI2zrbbfdirea4U9EzuQqCJq
G+vNqKKxy8U+nDMuSKSEMg==
`protect END_PROTECTED
