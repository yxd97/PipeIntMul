`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
APTztzCazNnQO4Tq9kvfKSOKtD2LPqNMn48I1VzNvYtjnCzsGbUzU87zotc0ciAD
nbh0ziBjTTWjzNVAvxJFrb/V5B5QqlSufYmfUoAKH0A5DfbnYvnybRYBtT3A50Jk
01GbPVxxSHyIklp/7whVeARqSEqyhy7HaHvRBRfeq/w5bhN4cvcy98pwbUaSMCtz
jbWi1XzwqP9PA8fb9m6avZnHiFfZjV8ccE1PHUIhCDvzB/DJOWY4QDdr8+8IBEHd
dy4DxlM11H3OQW95rawPE/o9Br9dExR6opL4GCMZ6Wtgn+Id6IK1+aqcDa+Snwzb
+BApudjINXehQvBXE10RIvUQJigokAC7eUC/sJ80/sX04kmys+DQ9tJNwvXAQDum
YiqNKhUL67VLvy7Ndm9p59V2SS4QBKnZoTDTs1rqK2DQwS886p+V2KKXQ6nzr22v
lJ3KuKMOQlG9bO1JYOFw589lm+7tJZQOwIELVsnvJvBmoR9vBTYvWKtjlcm4DirN
Id4AOt/xas3z934Jgg0S70tr4htwY3Apv79c87WbOqUhmmgqQYmiJzGsTWUybbCU
mZ+PTAZOC4Xp4GtL8jv5SHYCfxmPC5ireIc/vPCS4Y1pFICgedr8xzE0D1/mQkkp
xqmKqlPkUsakak4psGNiYM2G7vsOHFlpMPq9n4+CSqwoMurI2fd6IZ4DoJloG0q3
HP1DtIM9m4hz3mBv7rLe5nXSsMFr1likFZkert7hA/SU9T5gJnSt06O0r2C/UfeM
gsfCIZfz8Ecnnynve6LEFV9fc+5zbpQEgLju2KUU+UX+dwMtc8R3/OGBD2x28i26
yZGHC2NWXdXPJdwPpfXYcAo0udCU+pY0huBKglQAf/944mpDeorIcwR7HMUi/3dS
2ZgsELvW2Ke6uXestPGDo+XAoX59HZybAqf0j1EQhem5Uk4PcMZ6mdFHpByR/SbC
evyY8IaBVyuIVRjb2kyMtJHIlElDWor1jlcoxjUd9MABKCdLgKMb/FWCrdMBxE7K
BO1fVaLjHbUVx1qbGNHchfxePVRe/K9/exiyVf6uJqd1v7cTcJk6hT9Sf/aDQtl4
PcjbLRXp3Fp+UiYkRmEndnmB1DCnTQPNVix3DM2AkvA=
`protect END_PROTECTED
