`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OoEqEYXYYoeZ88dIkuWdN5KzSAVpcWzTYKvKwIecxU0eMOFAQ9YOHw1HvPtGw4kX
IG9Wzr3q2okNgbH3wTwRTpiXDgCTlzuKtk7qfkKkz0y+r63x42tS0noANB2h/HvV
4Rkypc/H6B04JrT9V/wARsXmX8JqVVZTwYgtoMG7tdh/jPj7T9pWPNwJ8hBb1qjO
/ugbzfqCnunNsbQEaydhNfdlC7TpooiawohiwIL1sPKeX0eOTNgtIYgNUL29nPou
Q17vTyNeLjgv2t23ERPmXRfPStkwLq/KmTdkwXoGOqcdJ+zdvzqSwpEnMGZYvgeY
2En4xLvMHrqWG5ifSRceEDfn7+41c5F5Wp3kjuN/O6SDJ9+R+jNr+FUDY8e/xgjI
QPxHGWEaS0S43k9Won6EsvAazOhc6qMObHfua9zTJwqIWBEvv4fmP5O5i5IFMCXc
ZTIwh+SELcjOgAaVAcd6vbuNM+vse7o77rGvxwpBvLnVSMa/FTPIFaSst4+n1aDC
6TEWOd5nGE+LVHg4s3Cgzgk0qcd7ZyccIJlT7LJD1Rux/08M0ilUbUkIwSkzFNaC
S0SYjswKWqZrCEHB4RVx7vUuIGB0qvqT3ANoTJOF0QubDJQcrygLODB86O+PbOfp
YkNJChhmApZVNkRp9lEe0zZ/F1glPSoMAVgRgdfXhiXPvWRZ3PL84zVtnNb9XtCP
kYIEA42qMHWmZr1u3dtjQvXjIUjXApcNGzWbt4w5z6NjbgbPBVk1IFoXLR7g0MTg
yXW7mOheAygaUFpAV/xWGi4uVhvu6k95QBrjPso5tAlXjIaBU62FX1x8kK3X/zuS
OI9XeOTLJYWeS17FsDJKC+/84rgkf1EYKC46CzxFgKoRqGEzr1yXn/2dEyjg81rl
j3EIiJ4E2HQrWJtyaRshomPbf9dCKDhE7i+R/vsEJQXy0mGwSz3SmPdFmRv7Pzai
H4q5ExYcytswfsNG4PZfYP4o688x7mgJHUychVppROi8CWbXLJ8ZZmQxdxzCVXqr
h9DY8hAYsATLwjPlunQ31WYA6K/G8Va/cWvQF5uFNhq6UvV6WIdTRPlCDs56khFa
NGOwYW4Ffs5qHZ4xsyDN5azDpGAGpCCzyHk16jn41zmvRDlP1zNiXNU30G+20i/e
Cy18EcI5BqTDZ48IOchMJXBGAyxN4jbNn1/txeKt6oqrNMf+zOyolJQTglI/N+Y9
jmLOV7yUIM2s6FL+B79jwFX4ShoJtsaGIW2uy6xegmMB4oQNxeP/tJ3isv2dUMfP
EakpHo+7xAyrShhTkLPpGr9ME/xD+8rLhdWob8Kr7mBEAIG7WR/6j2bf1cA02Da7
NmAhaNAgyPpniGE9G/UY/4x7aahn78fz2FCxWbX1gqN86Aq1FuMbn4cPsxO2Fkta
vLIXQzmc+JCv/BL5dAQzbFpgLArr5V6tXedkt6HrIcmTPIITYxYBEEdaNCQdbq0C
3QNxjC3FvkNRMFxVUUzSxQ20qUTcHmHYHA4L9TO/fhdLSyjPDYo7NfKgFrfA4ZsJ
FvbC+wEbmmNEL3oEv5WOl+K71r+xtY5gqL00Rto7AyOUbRdrRyQtM3xo5C8tjxmj
1G1L3VXkEeFKS2xIv/2vtqeecEAMcvLc3N2DuwHe9peXPWh2J51bnbeKPzwbtWHT
s9/0iaOQ5QYc/pgaewNwT4qbZLFffeSWGygpDqgm/Dzs/joH9XDVdPafdmK0RzkK
aY6X9/VBxh891MR49fIDbSMGpDGKfFzEhFy8DK+n5ax10BdhAD/qSaajA1UfI8dr
zyw6562CsQJljKKm2/ejml9r2xUXtMDFEj5+yARDhsldQByhOat0bXSpKQmW8HE9
7pHyJj00FHsQcZLj2SO3QwXTvP/oZvIVoVDT0eyS5p06tHDe/HK0t7fMWZuEDLjG
5flDvqUJK1QgMfKodQsX1XulKnykMpGnorC20wxjTvrdwpOShENiQ1Wn274w5HoB
KcyIvT9/fxVzySg3/zlsk7cYmFKS1GWYbUFk6zo63U9lGHxJp5pVCeTcM3dMJq5u
h2haw8yMT371OQnq9YsAs825bikDeCMSZEa2dCP1TWrJtLz9MFXSxR9CADCzo6aA
vE2c2medR0DpEXT6XQcB9VjLJxw6qxCpuoF4WNB9p1Or5+fXBHO2Q7f5oJgH6HrI
mghlJFrGpCaHpZMllhOwRmfxSsLS0lPkVMlDPuHmxe83+MNxHbDKtiIrY+igoS5C
owBUmeODYZJYoG1N2qUoILn2Hx9djrhzj6oSye9ZEpRJO4FEjRH1b/Frsu7nfGSh
UwOOYgafYAI2H6Pqy+iAASzUAs+fi8vgeGRALv8ECQy5ipr4j2DluAm6Z/W2s60Z
0OhPggtM6Od5aXUWKT5YEojJA0JLP54wy93FGzz7Jv8SiVFhrDu5HhoorhWs+zWN
ZHZ8nL5JNAYa/brW5ptZW4bo6KepKzHx0jlyTUma22U6HaUauEAuWD18VT2O/+ED
vIQAlKdNtIHbFnFwd0i8O1XO75leqboRPqpkZpdFEy1LBVUNOnAUQxe50Mmfftk+
wbLTEqCZUB7HG+ytdKMvpmjQ4mkqmAq3euSrdU1Oi8tyUxJXO5c4jnfZVB4vpiy8
lROsYFw/ukISeaFdK087ZxubL4fgojU8LheFw5dMJP3e/IsX2LwQdqxIW8dzGFDm
ondpnajCRmDpBhK0ZmFvK/cgzx2tOmkzFt57E2gbUmeQapuv0f9HpyXJPfLcvI5F
zlrx5Yq3RMw88L0WVIUiun92VyCVwtKQ7nAhD7Cv4kB/LPu5TH5B/XGlL5/k8yO0
APdZZEyWS+IrU9GOMPsJ3565ow5bcLI7YG0eHiPad6cNplHzmKdWE88ayjfww7Dd
GmO5AM7JTo5pp8ehYdSMXbsu1MrMeEdat7kYa3JdPkwO+sZFxB8WdKBbwW1uLOJS
gIesi7/yBY4IY/3yQyOrCngh1v3Y5sh69IK8XRZ7tapWf8RiboiUIHhIG2GQak1k
fvkooIv4hAb65xvvr6PpH+wnmAzJHX+2xuXkC49niuuoMF97quckI2K1gRO9E+yc
QO3lxRUFygN1oMTH0jPaG7U26KNY+3T7egvIglz7hNg0s9BSlERKvXk5Tdn+EaA6
b/HS+dmpYv2u5JHwVeuJxc5CGaJBCr5GE/aEYabEdOjIXQGFRZLWHIo+CGnBh0VW
75NcjRj7cmvegP1KdqILCqSKf/iVAzp4QjXfFl3TcKzsxyJAoCVErhOw/FdUizVv
rURW2DA0Bg4EWFP7p4/uS7j5CdiJIH22HlFqrZBtKAO7Z+jdExR/9l/iysXr97Di
6LIwaVw1ox72Hv67u8PVl7qLDfg+sFiDIpva3gbzKFeuMoGwcpMTI3qmaP/8sStu
1SiAvyHJsv1hJJMuIo7jQvZ7DuYxTDcr9eemY+BOawyjyANT381ETWW7IFUL3lDN
wbrNBX7ArQk6vQZEV6M/lIFcU8pDCvMyMzbAEpcjOUuqNs+EQeg8kQ5O5DeCoyOi
Y0uPIWFGRCtZSSjnVYPURtTQ9UMdKqImIFdVBVAPE4zU/TD3NLmQw9Ik5hMiakvP
RYvGVM5fWRPilTLQfE3s/t5z0NJwYitK8rXXpcJ0m2CIUnny9MZBF/9q1RPEB/yn
jfFVLyozvbK76rB/jgdmZDx4Wi/maDqX5BwINUUakazmh/v1xcK3KmoQVX8on5L/
tHFD5GqoLSYjfcx9IR47+4eFfw1PGu2n6ckx7ERrzO891vaE37gc775sCbFbWXsp
qQmqv50P/LarP8hXzIcd5N1nrj5WJ2K9XFNVGzyO4feDFG6XQwbaN+wC65C93n2v
3i7AxSbPqnJ9SW5a4eT7onh7OdFPNyfYzQvULcFk4Qw82M1l42egwUlJOGTQL8rB
AsdnvkzpDsEVVVkMSPSBM7/iTusLrb720UAzmVdiJoVsz7B0G8A02sD1T8KP+tx2
AdaXqahCf9PZQqaVG0f/BVCJYnbMHb8O//zxetuxkBodJ1EkGsjVrESPtFXZPbTs
ZQMUiAZos4E3wMhrHq2JV6HTaLImhEAZQohZ6fwi/z7TAvBR5C3BodkB1SvWA4OY
lw91IRkL3Qu5ZZ2ScMVdYH3ylJWXf8BIRuJ/vCObhNYLIe8BI9rUR/tfsTGIslp9
tKOH7OnQD3PenvDbo/oed9ekJkeVu9CktNqYl2UasKojIpumP314ERVWN65GdtMf
l75l7aiqYw802usDxvo3ylJctFV9XkhVnDCvFrEjNOUu+48KAjCuCTJsC6taqFjN
06p80Wdafu0dispYWqOjzXx93Xprp8I08rWqCU85gB3LzpGlK+Lj1VvsKRxoeeMY
wWP+U/yFdT4fWYoA9Mi3wIGmoZXCDyAD/j189Mlu4cmuVQxEZ3lzte3BfW8Rek6R
BDTPkeo59f+HL4Yp5quAydXTUdzTJN6paV0lBA9vqWtVfdKBgXVcdGuNSyzR+OvR
/9ZlSM8IkNZPiKaYhQmK6capzYBKlMkQ9NRcYU9hilCJR3VugoWgBV+KQEknRYUs
Yvu9WS4fksQ/zRbAaPk8ld+COX5YzznbYkCbI7V6cyk/xQBc5VjysFLdRXk8K6B4
G1IMSZvMAOi0drrpeMNyvXdmGm8s/NE+abSKqAjR0b6cXKo288KLtzf3yyw9+6Zk
xSmQNKVKTNDRR0QqjdR2KZs77G8J72KmUDwAMxSCy1eOZcc5NOWCZMAbxV4fnkj9
/oFCISSfzAH7kHq42CaMcqjuAXC75bNdht2FM3gpF9h5IXZLFr/KgAcaJ+XjmL6P
xdUDAAC7lPScwKkSeJfTRZ6VdgpjpJlK4iYnf+zyDdYV/8gSevHI7C4WV149zcdY
NFlVb4MkD6i0RI5dF+uB0H3tMhJPzF9NhgBJdmZpNH67jmL3bL43kuIUHOvXCpiV
MzyhtOHG+wstrCkq5Cjqzw==
`protect END_PROTECTED
