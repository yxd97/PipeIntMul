`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wDoEEaCglTIxBds77gXO/zDb0SuLcbIIjY2D3moCmQxm7eIyQllqosbnNkjDVyek
iwfOBP0OXb2hve5gIyubrTzLZoBhaNvM38UUwE1UZXj1/fIK29sfh+ojZWd/WT1q
3/fUx26gX/laONBVq3Pi0SKKUcdVBk9DKweziQ/whirUU1pCDpfnQVEdTwVdf6hU
o39dWcTkOgkes+m80VtrqFHcnRYIQ5qIOASqV8iowXwaR5+L0n/5pptAz34r0dPr
FD6AGDZd+ibAmce7DZDPr/U+sueST40i7yuYRKFSLyynTCiPeVdX2W6zpau8IFgJ
EjcGOs/8HDFsD6Ta9FEM2W8ibvVlpj9neGTXYMe/Jqi+/431LXDybEi0gmyARZLf
ptZwEyibVt5lfy+PBeVcYGUmb2BzBwiFENkZPcToNP3mpv3Vvt1L4ZFeJ4d9LVSz
ZGFxHKEyBSsWUEtsvNFdUgnI3W/PM9OxWBVaCk+n9c/nrXR//QIaLlUVpwQKgiwp
ZVzWBbWjn51/zOTZxeFpk4wmIN5WuqSjElGS7krgya8d9T5NUSx2T0Y+A6zErnFj
fan3LbF2Qhr3yrlaRs8g2n1i9aXaa8vJarQ2JnaE91xAgUoTMMdM2K2fDEW7Jz1N
faDsTYG+3FrWNij58BeXht3MKiftgrL9hSGZT+r+kqmi3tYyzvAk65nyeQ/5Rdcc
sYQ/egQ+po2EIAJbtLTSlJC9r8YXlemR95DUQwdnxEAdZ6tUe5VpNC51mfH2qtsN
8MryAwYjxJEbd/Fb+SzyqlWnx3bk+kyBOCLi99nXTRs4KZBwyeabTxmHHPfRTB/i
/MtNDK9iHN9TaxzMTBGpH6Ei9MlLmuVLoBXY1KAaPMoHlN1+Uq7gDZfC88vsVPhx
tSx/qkR4WMJ+qjPP3USvxRDZtqad3W4mStOZCfASxiw3WjqnhYxiLS2/aBQRjNSV
2IsQk6/YKOpk3WXpoJ0U6LcZ4FWmi+WprBsnKHvQjh5lgEpiQeA9vB9nT9eTvim1
`protect END_PROTECTED
