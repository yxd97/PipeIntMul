`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0cC857A/ZOA6ObfY/sAZQy8nvfFRBhU4zeFhAJ687K6+YOHNGjd3mwfW1cSmZP4j
AXVSxJOn7yBH0+1HdyOwuO4hvLQJUjO25uZPxnO8lf3giqcW1yoLTeQY9dcAaz0y
1ZCTT9ZXmIS4hDsKJprha08sfxvAtRE2TPfo3Goij90LpUNh7QbuH3MNEaNhA+82
/7pmdco4YClzWNb5olYIpLpQ7yWxyjl5/I9J4o9aqN66jsE86IErLDQOM6EOKHKL
mY1uNVHdrZ5/NFTnjNgWZoQskCk/7fuRLaNtRx6+XcQr1ZMvk2pZlfHpu11CAyHB
inQI9mVIGAYam48MGCx+aeh5Bri4JO4Igr2MmSTRHSPpoY53Z/O/BSJFfiZuhFM6
XeUjXCe15a/DfaBYj16p45tCvKtdau5shJuyWZN2gy4=
`protect END_PROTECTED
