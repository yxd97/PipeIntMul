`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N935M38QM3kjIhSO1SgOXygNCSy3iJW3JdhYtfO+tmnzkepwZmfvWa7vi9I2Qop/
/CtX4yTWuuPNm7FhlCWW+vQNstExJP0hr8QltfybtLhoZfEKSXAAbctaZx32RZ17
Lejh4h6/mMKaoFb59NxRQqrz1UaIYHIbCun4BJcEbuPVfxKOejUJLY2quOfKxl/K
s7R7H8yaFg+zU8QFx6S1EEEiBHf9Ie29nf9h8zldpjI+TLc4t00wB5/bIPpJXI9K
zmMBCprI83MeOcHEaRGEurSxm6iSJzpRQoZoM57kFAyw/2AcxDEL0UB8ViPFpMBg
2LSnIIJqa6jQYv0rKmvFwTzxMZ5tZYwHur/tXND7Qgw26etS0rPPB8Rgp7/DVy4K
VMgKZHA0wJ7GbpB8XaX9372Ewt+Nkix4Z7IXoinVSAv9OqZLSzLyeSA5D/2isqBA
xWTVXYVeleb0v+4jPYzvczZfk0Lllde9PDsGgom/WS+JLbGUeLd214OsRbR7wW2u
A6plJA6t/O5YWAA+i/R8WSrA+1GYEvNOYOxYEwu/1jrs5D0dq3cKaqNmIi/d+CdH
EVFhkagjFCqLBaLW/tBpTAoonQGEkhkx8MdW1zpjeStPeZSBdGI/HgLzBujmeFf1
7oOk6ZIfK5ZOQe8oGjyjJS2Bv1YInb4194E/L2mBamylemINS2W1xULiULRw0OZ+
hCFV+URKcYiBcil8tfF91AqUg/OLzoIOwH0GgSm/jn5wjfXqFu43b45Qs3O62Pjq
xeU1s9MER6ASdJJfvsSUjzx5YMusYA/kec4rchCfhAqKLOe47dEQuiA5QfGnxrEL
DPIS48DkjjaDhmQPkTp2gzF/lIsLQ+qsGirbwvgvjOTnRvrw9hMb6guUg+CXx+fO
jpbkOdLXKCNkSI/BkGydPtPXFTcrFp9mbt8Li8dlB8ZcMJZy9OZWvo+k2qD0zgWq
+FRlkpIn3Rtsr1TRPGA5Coi99LBUec4vscYFcj5VxrK8CCrXV6gZq9Fic6OwChlU
iZEoo82FKd5v6sUXHczb/vK/Ba9nk4N61c1gQHsMMzuruh//P6Rx8ipTKNwMILQd
7LAW0docnrTd98RXMuoSq9ZH/OIhYnpXUBplad6rGV4fEgeRQCbesexp/nvfGRES
ixCUfsl+yJ54WZg/1EL2I172SOq+PEgCjFbJxWPZg4q8136KUl09BdGmHG0lp13b
gR6gdKvF/1tbIo/ATtbDzApYo433m7PryvEvn511SENbatD3OKwDi7Y60LAtPce5
TAhdnT9r7Q3P9M5wDwI7dw==
`protect END_PROTECTED
