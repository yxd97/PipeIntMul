`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UU3UJdjDthIR8j2KSZ/jphAMQlTJ6OCzARxqrtJmccRoSq5zS4JEN8HEB5GWSa3I
ffDn+LdO5WgtUYP4n/bfee0MhXg4TUluo8zLQjQV4zBt7LPu2w3P+ZN1sdQ88elL
FBYn8NQzL7CJ2RABvcUBY9IzP6ZwHJvDS5MA3fwbbuat61v3wFIKaA91ukHS+oz8
OQe6+lA09E3Jns+AdP/aV6+PjGk9aGLlyOs5Ji+xH+29MTo8e/W50oe9HEAJxNvt
sRONlGp8YZuEynqM8hMOWPv9eloJY9eVsZsflzxSyTn7KnNFTo6CLhsDHklmHW1Q
4jOLnIFVkoGnQZ9Y61nKrpxRXpIcMobeNMeLp7a2j5E=
`protect END_PROTECTED
