`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZFJhkTQk0JBjVsw0vsfJcCVecNIOxYHuMC/TU9M2/x2cx1Owv40VNqt0J2nDz2pJ
rEINM0vvWhHPsGUh8NCdtOC2UepIUnZ/K3CTcDmPrIkFRZLjRjdnvxEhB7Hd4cdp
eM/OF7WR0fu7Eq+YVJIep9rSGIsVANbzTyMmFjN1esUTWPATKtrNTUwstewaaa+I
U+sbkNmQZyNJRcZcW5uwQzXCKBcba+6s9vwAjqNCcHXbmnlNmDasQLNxArJDL4Hb
gpz111+q/526eX2dPxOfa2Q+ffbNjDauYQMldWFUUkjvgTebQ+bTNyqyEwi+IFeo
4pcFmBtRd+8jzsClva/tEghRe34GkmPPl+uvm5fwOvoS87rjGN+5pxDp0rSjaopV
rEWHZrEe1FgSZXJYW9SsliDL9K6lkwA4NlyX+kIQ3bUXNSvxRVhAn9UvMrGTs27L
BYKSlaU7PH81bVXRBUDIlSAstkLD0WylWAsNpsCi0dSbOSr6YTlaW5qRDKm/6Rh0
`protect END_PROTECTED
