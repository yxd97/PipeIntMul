`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nuo0Od6WsloEQO57iuO3ms099zK5KqMBmr0RTr+fPup7BMPonnKMKMB0Qfqo11AM
URw3ZEYV8aZ/m8+M+38wXEMqbaMSaXqkTIF90mmiw58uL/6qsglY59on08Wa9k48
mFShQGcIBm2ZAiDZwX62ob17K/lXPfqZpqjMiTlO5hI8fO3QyRPSTInZqwaS9nFQ
ljzZotR1lET6W9WCjl1zRtid2hSojfyDThWpC7X7GvNUX0ReijpHNFS+rUw4nXiG
Zmnd9smPqu3TIGDawJb0BkVFpFNjn2EvcTn39gUnbVNU+ImueYGAE+spPXHuzXV1
qiiU/FRF6tiQO9TZomkh3tsLdB1Skq+Hs15WXT/a3Iyn4vERrDWAXJppRN4xHpXU
bUa0tDcapVBXu/IbUteHavQylVIfl7aXHPKNryRXwpAkaptKS4JDYdxW1wIaCE+w
g4UsJUpDBHbagvyIys3GksUB42niauAXqCBRIoWHRlg=
`protect END_PROTECTED
