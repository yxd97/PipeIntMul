`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QcTJuDH5e9UXKdBZYmEtLFLFmj04CSEgC5v2m2gnJguzQyvbS+IU3QPsNHCiA0JZ
B29lKbejm+LdSJkK/fdgNmA16cdlDuSLcqlhUNj8iiztARBtrfUHzDRDQboFK5Ze
FTn79gPjaLRo4qMGHfl+fd+bOqP8XS40CGrmFDpcBnuJDLF4S2zLXMyUyL4Kd8uQ
64dD1d/5cxegjcdG8RfgW4KwimOaJB//E4XVS0z5J7oxVrS0EjRet37hrASg40c9
dTjt+KYPbzEykjFVFmqrPVTTCuqD/QBaEQwpWPab0y5yXE6wtpCqHqXxCdCr28AO
X3L7ShMDoR0hlMQ9Bn7sLYfweAUWSSSaAVGcDuQu7J6OQKA9Lvcjuoq9mSaETrAI
nCoUf81G+HDbQTOXGvwS9px6pVGD7GHerjNiJHKvqILj8Wj30hF2yM0bQ1UNsC/n
5oxQ4uS/W3HaPOOe3lyuFU8PJ5mPupieRqT4UrvOwz2BmXG/Lu4ujJhfqgPYNLEe
IWXxhyihjObE0jB1VE66mIWy2n5WRuzrfAvejLD8fIN0SdBehvdP5T/t/lVhSMWy
rzGT0VslWoyA8aEvHpt+dz+rqztT3bklIbid7UvRN093ZpJ0ffZ6+S2TvlCI+IYN
m494xKj9SWfJmb5wnOzEL5U+ypRItD4WEW4NbEOBV3zisQff+vcQrotzCB3IAfx2
RjAcJbcKS+uhZYWkn4C1iM8Sr8E5guGVP5622Q3CwsYr381l4sdywRqKP7T2vczM
90o9Qzsk+dZgvDc578akqvP6rlF/LALPpdnSshO7MmZ5e+6uihKyvX6rAKNFee5r
h6NdkHqKH3R2zQxiJdCupSp4ehrHQsjO26ir95tzZjbBu9RzsQO/RZSDw/w1gC5s
mYf8UrcetuGQDwbTCdoJpQ==
`protect END_PROTECTED
