`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LIEDfqV/3x5jwA6cC7OhP+LVsRyvNmTwr50Bm3a0BNC9hjzQ+5C7Hh9QuUQiccjx
D1rKJKGASCcZFfQOKWauc6pDg1v/7dz8waKZg9WRGVSVczKwPeXVrsNVRees4e2X
OhAyfO20NYxfIbRHaWx9S++wkzEOo47fdnxcT4YSUVmufhERYDQMDs8ZN9PEmYfH
JxtyLYs0yGLibY1PB30tami687QL4YA5mgXkj3ECK4TgK22NKQ8s6oW4smgSdHTZ
lz94Ex4a50ndwEfHoT6fdyyU7e9ewEiUUvov3ZLxzBivVCudkVL7oErH4H7QJX7H
+vXxJsKby+DcJDnwv+3PaC24OKNMpIp9piFexyV0wSYaBD61Wbd9+QHoDKlYp2K9
8bO65OaNKUqKuWzSE9UZKacRLQS2g25tuKfXFgK7OCff59rInUvhpcyTALs2Lvsg
pGjt2kCgfhjKWA4DLO2UwJFmI7x0g8kgEHEkoC0ew7YKd01/KmAp/wIodhexwt3E
5Np5jXPj9prfCrmY6nKV4lSu92xj6Yul9EJbLcMTs2WFL3AknwUr+52YCe6dC21E
`protect END_PROTECTED
