`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+hZYv5HhjLxX4Ud7ptCXtb6Y+sqNlWP0+dxH4ICXfFsIIeSAqpcu10xKZmIrG06X
pItKDvUjyB6qYr+8r4MTE2UDBCYytah8fdPsGlF9ysTNgSNZYDIqorBz4s+eSEIF
sZw64+cRCakQN2W1RGcThV+/LFNeHbwNBxzoEvJPjktD8CactdGVlxSAi7uK/UOC
kWrQa1DsMxwY4zmufETn0RlDedKH6OxVMIPDuFq5DQn3EU8nhJi6gK87/VaFLoBt
zrPY5k89N5FwcZQIpoF06C5s6743sqbYE1dMZ5xGnuiUHBjz/UxZNKCxJ3U59NKZ
VR1wGyBcaGLToliPpwsDq7Q1QXE0vKf3ksJwrPPKZVRELZrWk5b/fztxIdglYiok
9ILu7JcnHxhwh6I4zosPklSDPby+TR7mODOicrofq+xhIj2WGJ1Lkj65a6JhIuQj
vCgp67U6f0pc1mjbZi3bso2EPssAaVc+DHMkJC25Dnhlq64+GMxqDr2wcUaD7tgi
IXPHqB+mofg9c2BB5zYfPoC8pS8BTPJpI4x+9QCTtE5yy+cCfEl4JKGTad/kstfv
x1pp8yLfoWDgOcjCP6hf33xaUX6IDrQVCuzmozfjJ9G/egf6ByKLOQ8XbGOk0I/E
WkL+rO6vkkvAekAAUhC0MoAq6xRPn6FXALogh6bS5/LXLcJSl4f3AZuOo5PyQtKv
o780dQJUDLn30oltVtSbVHdCbIowYBKJLPNevObSNuZqFMsn4HQhh0H9DksjuJsO
mmb6O3882w3SKLEZwssZK4I607XxWIFI8ruSNea5z8Lk4sVQkQNlG8D2R8QCKLYu
zdQq4f8lZ8iFGULgOjH/HZitptSEZnnKzc8z6aHp5PIKozCO4PyXPWGMelQ9WWgi
0t2tPY9BW6DzOTQBBo/Y7SIekYXQVOr6iVHYfktlDzimKhIkXP+kV8kCT6smK6xb
go9pX7VRdOTeMq6XyiOKQ57RiXPdzAyHkIBv126HFkUn/VjE2j+fvD4ZgyrBJMN3
lb3dHZRpFx32fQubEkjlUSQr+m9zgnL+6DeuSL2ROysK+ZYPpdF96Msx/rJTyDli
EG3dcZ+wcpqzrMfYuxhMvgIo8uOj/fCYsArnrW2uhzhVN88mR0lJOeJl/wv1pDR9
nO7goTa2lU5yp4NUbMvtS1T8c1to6ebYzs/afr6gNEYfUmygki+WwTShSzwmjzqw
i6uSlnrrO8iXGFqJDxF18jUE3Jvu7Kkk12kvzFLyol6kFQ5WS49Xf5R60fk5uwgk
EeDYoc3A3nKTdYUo2J3fmw==
`protect END_PROTECTED
