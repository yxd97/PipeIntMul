`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dB9VactJH6tpBuBVld6Cj4eNDms2dnDyQf+FEIe6Iaos2n4PFxLUmTI8qXBQ2dWj
CxJPS8AS4HVjOzgtevUFgiwnrn38f3+g9lh8lBJ9wQuB1mTpebptEnRjKssJrEzt
c/hTTSyxB1uqU+eRDEZXlmdJDLTPz7Dv6B/hStFWp89MRGVYR53vSaHXamNDZr0c
bB7VffTxvojFYt9y41GCrvZhhFW14V67JF5VCoRR6CwZHa+OOhJMKavKEQyRGOcw
rh5TV+dlVjo/qMLVdcTG1GICy8XGugk/1SwEzC+qfSqLVbnrAVUsRNXXDg/nbrAf
f9bsksr2tkRKPwkG2aVucb9cRL75J/6VwPXOZUqFuKXrLSSoMTLCUiDs381YTv7Y
C+WT+OcG8mhk4vZOtigceENyxTBJ7RKanYqAAbPEIgYiONVro1DE6QMwU6LnE33s
SpmtiAScFfumWM9Jqr227xapEgKTGqhg84/wRUIuNo0=
`protect END_PROTECTED
