`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QwVElQv82kKnrhZKkYQ2PHJkcWgmL1ZzRYizztf/sMcXjBUosiK/K8zrkM+0io2W
2zG9wwSt6D25/dtQNEe3+uWABtFgJ1ryzv2iSOFfB2S94neckS2UKJLcS8STQCYI
MHbsVbnMsW+svz0uzvwSSciCs0HR7M/+rc8K9zHaJ4ygjMunJ62eiI5kuI93PsKX
FyAiXytpLEDQUbfEaXRg7jPWmYeF5uNRKk/IO7uc65V6vWDQKyRY/+IV6GzZt2TQ
2xcSzfXg7UDgrqJZqBniKfKTz5pkQaeKCbeXRK+FGb1XkSOjvcwTK37wURsq8syu
VgVxe1JrDldEjJ8m0Z4CagHfqtSHjH2sCrxECsM4tLCBgqbhuD8utLXVpwTFbkdX
`protect END_PROTECTED
