`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tGZbDDcwj5mjsGaBntYTQr+gQBXnlGfNrzWdBjkO0fh7TyszY3C3f1DAzrZLAVu0
AWkFCHviGP19WlPZRW++0+SNyhcrDKSi1dJLUm1j3U/yolzTWoGrrBc+JiXqiqus
9xM4ZvXTF9ieeAR6fW0MiQtFp5xekJr+l1Vs5yEO3WvOPH9VI9MQ5jiCeahcokLL
q1zEAoepEYuxPpUqbWEJ44zNkRo+16y0V1CZalyT6HZqR97/l9OIhYlCaM+b/WsG
KLpK7ljqJkrrfJ01b6/afw7vxMENccOXI4reFgLpOZPeCOuyqol0eBQ0TgZ1O1Eu
n3RP9AhYLhr3jrLVk6u2U3aIr+yx4nJwU91ZIx7caV23wY8ZUT9QTVVg6ug7hnON
VdE/za1kgBzJErivQ0An5jtQnWeAjRxhKvj6c9FvBZm1zzgZEZtMOvOWpuk1rt9b
WRIGt0h556JnahldhpIuzvd+sWv31Wc+0YGbShnxRStG5+yYjyKqjhAVnkUyihje
h3kYhSKijcPWXWPMtGteR3ZYYSqC/D6SZluyVlLPXbuiip33PxtRH28RUWqftb7J
Zba1lSSMS6UgiEVmrB4NqZvp08RsAXqFA8NVQENkMqtOmf+r2GQ2329NJQMJue9i
mLLyDLNIJVSZajxhuBNGL8e7VOg4EaDKtQOHhy+6z73g9/UlxQcE7KbXD1D+58+S
d3KZnD93VW/bGfnvfJk/nqjxmHeXGnzPlKEWxLRDZxx6Lb9YruSA5pooST3MesvC
Bt/yJspFXbteHvNKwYu/dsc9jR6FPDdbBtx0QBUtENzSgN0QfIu9/4QixLT4wWTv
loRiVz1AlD/IAyUb6ufEgqFR9P8h/HOBSs4/wsmtg7ZgsOSdCZ00BNlofy9pzhVQ
KRP159GaMHnbcsDNuwWFfCANre4FUNnafiKRhCOD5yLZsE8ozggb7h4aVrFJbMlf
ro0ZoSFK8OGFoyPDHGtEKFrQjj6tRLjhcPhcsD9F3Q6NUShNCygVA9w1NhbInaqe
MWrb08ZONYJGkjD4D2h5MK24QmPxZiPxtMQ4W9IVdUQ=
`protect END_PROTECTED
