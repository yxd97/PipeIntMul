`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8AapkV2mgIQLmrSBAIueRQ2/SVh2lHyBdLcJA6++8k77Lbbohuo1XJxoNgjtugdi
K5ZErtAsN8AvEAVNz1ROyAgH5cy09NwporF92lFuKViYNkJftGrZnn70/VQBCJ7j
/hXIxtsviC6umPxWHv/G5N3TKnJSxoV4GCvZHyrElQZdpmZJakKdek1k7G93GHMy
po9vGfUaVRdPL0l6Jc0sIaw/4Vvv3fBg3wn757I+MjluJ+xIltTQLigvw9RYZZI6
0UqIJ8OELi/1U+4Xgy60S3tCFkuRpCe89mCxWi/iCJeYXaByX3tJZdOXvMbv8Yte
zv88SnNcTw24EcmOi5aCi9syi7upD1VZWOEk02BrlmEw5WeQnRelh4733ganQ/CQ
oA7woskOxfpt2x5GMokcdanbUzxpCtjCEvTDvE1RjAHOCDzzvKGgOFr9H1Evf3ch
`protect END_PROTECTED
