`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YQ1nwPFh9e3BkYDp6eJZ5xQJ7D5cv9dPtYZN5uFdve8iyLj5SN0b2ahoRbkJaFMI
BcxXVyVax4tmN9gmOOtgQGCbpJAlyCZIx0Qdhx0+x+fd4Mwnxxo999LHxkU+/xg+
NCQjIW02skfYA3qp7ScqNTwAccPh10FZBwTCiSQ+YSj62d40fTnvzZDAe5gjlTHN
hK3b7seOEDKbSzvbnBW9vN2X9esXr8FENjevnAd2XDbFWUYPjed4GsQhhyusfpth
2xW7aOHbVczkDfthUoCGpQu4aO51xkt7I8tQd1KEr6g5kxom8w8Vdxc9VafHLP41
dTWfTGDtU1bvkT/OnMCyqpzZeFAZh5EZsLryufDWfqs18lU9C9lD14GGYPDG5un5
58TXFyDHpjvTkQ+fJqjzSLx+3M8fzwfSwATortyav37aa1Kq8TqxWCJ6BxyL5Tcg
OR1vu2Et0H9j/TKQ+Ev1Atl0tbe7SPVAQqInQ0tGk7laTFojHsyUq6Ts6BN78s5L
f6H6ug1a2FAtS8YTTQnGZAFN+b124N0D3D8MMD07A6IZLcVxyZnDwyfrcreT2Xwx
GBBTexY25KmOL1ZVcKDDvtJyclGgjLL8rNPn/ADzmBfPjvHcU2oOBv0DlNPjmsY8
`protect END_PROTECTED
