`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
J7tb1/vv4pfRH0nU2qwdNM6sfkghLXDla+IkfS8Gai7GvZ477JUR9kUfaCm4zIHg
5gqhFir81PKiFSnYDVjLyCowamiYajBZeqZ8cGlSfNkrKUy3XKVK31YWDoH6tiJ3
h4lEhZ4ydAAliZMIWvBXErtJ7FUhB1jbgXMDkSGkTaznVkVifbG+VOJDPUmDA0mh
IDuSrnDkEaBOEPPoT766JBDvRpfaMgyoAaA1DQxdLfNrbIj0dUiQ8JqIckIa/mXy
3CgUpk4f79Uu/y7ly7tV6ykZGxTmd7avbC9rCC+lFv4HmBfc2AFB53QI4VZ9J/Fm
ZYgd2ZmDSb2MuC2W0EGR4lR63Ysx02zfcDLk9Qg1VixZ2VpV2HDUfjk0pM3Amsao
RR1J/Rp9jCNiOB8eubylloExBXA4la5nja/tPMR5fE0=
`protect END_PROTECTED
