`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8Jl5L6LS3hywPFF4G1D/Y4d4h7E4A3tuTSUOVxCluHvc1iKwXyuxVSTDbMVF03nk
GVfUHUTmnn2G22c5DzmXfCQ0Tk8CynneDXfVM9uJTSWqlje+CcWzGA6BHbizNpeQ
mruHqWRLXc0RDE9Fs/iem+K5v7sWF9u1rGrpJgNELWTKgj8eM/RdCwFVf9MdZp3f
A55jKn4CYmF41S08YAoMS1WrEDGudQcnqHAnWqt1IGQ1ltJmXmrSG1a/y3Muwl9k
FJtJptbTxDYIeMMh5Il9fQMyv8IS3OB2U/83xV1LOGOHp4qtpCrapIoyKZvbzG72
aAVUPw6kLjMAIoqvR/iaDafxKDFDv7i6jZHap2R3NXxGyMXlXbExe3uAygf4oQjJ
tz3SUUI6CnSqE/LHW+75iYpVCH6eqRPdcsb7JTDRL+lRoNJRTcuucmKOd+Zw2uZP
RkhSUv5JF/lc67P32m88xGX+zSyr44rU4aZnCz7xnTfHqEY6G/3ZOATxT8XqoLkr
nJYaLIknIax3RwDoiRpV+gdcySs4Jo6IfLeYKFwqqKyJ7UhwCsyF6tWBZO7xCtTQ
U309VKOsvJ/ocL/Svu02vyPYDuJiZY7ALX4bc10UBkA=
`protect END_PROTECTED
