`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRjCuZV0W2vJmwL/9ZQ/nTDWuCCXkoeZubeSNz2YZOo6/6LL8n/EinMgWmIEZRRw
wP/pceYwr/cNWQFlGD1/vDUzb/xzXcpX0dZBqaZU9T2NdUAE7+rxXX7vYdD7sW/G
20y7G9xmI3DsMcQQYmeapdSLSzyfqe1l+8KKpjXi0NXDrriGlR7umw0uiT6y8WhC
Upm9vBPZaIppsmrNv09LQjvyNOQMGe/s4T1J9eRPejhshtRS1rjggHoA9ZjUJv61
XOKdSHcOLbJ1WZ6mvDRi+8ylwiqNLkLhAVHTkCKED351Pq2+oWz4nNO6ASZwc4it
ySev/wc5tKEcHFhx1jo40vrKVlbTsrQBSVC900DnVS0HL57SqKIMzKwQga245y5r
xUOmGRtmdA49Y/isQtIGRoISxMQow5+2F1n/sQXSvx0l1leOmcU/of09sbpvevY2
QmLYurwY6OvqTShDXD8RY2paDibqkPhvMR2Qo1bPlco8J/1lNlt1UanInOTpcFRX
4sClEuQY9V4gV9lLiSaI7llqm2+USolk+e2SLRmuC4kSUfdiUAlm3gOwH2mgP9mQ
2vWQDlX2ecRyiWIU99jLndO4/gTFzlgfiRhK8En7L1GpHf2XYwdB72HSi+1VNjTZ
56OrTUqcg7U4LVFoe56jaXNURATktNf15+d7oxTtWjoJHbjjt5tdbOFysnnqfcyK
rDWvk3bl9DuHcokSIVYMjrAeWwz9Rnd1WwG8M0tRMwa5Y+8y9WdUZ+dzVPLazfMe
tBspO4kRB2AEb+BYHTJit35pztFSR19SfTcfx7nlkSrXuaE2VzLkbMwQAHGJcSXm
g4a8iMdwVNmt8NaFjh4HzQ==
`protect END_PROTECTED
