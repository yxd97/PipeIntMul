`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
63PddKX1EyYq1xrODQblMR3Ypq5MiDDpvw+lvIj0k0nyYqwa+hgcdD8lHFRg9RuB
8hO1nDlSkGh5jYVglT1X23suBPdb8nhbnouA4Lk2QQCEz1r70ea8Y0Gczzx+K5/u
7aA+0ur+CuD876FZnchmN/LHWAzaiPCbQpCWd2BS0VqcmdeHximpmPnFe5NPmMuD
ZVGOWZoF/E5SiKybua0MzJdve74vqMfP7upPaNyGfFcd7kcuNuw8jKgoDe06raQe
4qoqYE1cOCJ09XQggvCmLA2aP6YoKiRg9pfFVAbZca4mtfK1LCD7uqiRYtYiTBTr
l94UOhR9w3fTVGQxuS6Q3EW54SaiQby6u/2rPM/m2OEJ0ejEt4L/eEgCJBNaRkzI
blajPx1qBmv6DGHzYTC4yuJtdI/jd4k5bt8RomPwJB3ev63+jtjtJCjSSj8eP41E
`protect END_PROTECTED
