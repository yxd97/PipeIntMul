`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0fFsTRNiYj67mIDkJfa/2CI9q6PhAUVbiDVmMCezq2o7jrCP11uKgfm3YCJZGbLb
3TCdESneId95mUVKs8dlsrnqTu/oKyBKwHJkSkHUW+AjQ6dlEkbGoUxvNuRvQq7h
zPSQIs9ocv562aRwcYtVTR3PrTaUQNiDjrqbX4B8ITzDNGUoo4FilSMW/GgxzQp3
B+zV7+T2M6taQe5ZsNfbQaFxVcZXJyhIF2ExkEFFTCbqG6Zukr1Ec5iKTHxILgDS
Cq6TmRqMpn00Oe9t7LIID3gae1W6q8XAWsZJDnrRPHxLxTE4eBdMJZaqGQrDwisF
Qz/zmi6aDxp6xRAxzAo7Z546W2TKSEdFstcI/bXkHm8z2JRiHGm4vcCZYIjzr8d2
ZW1SN4y50xU86WhJN5KyMjuBiMB7OCBRZ3Q3pirkV0/hrjkweexpr03YSf+xaPtJ
8txwELKhr4SKqkb/AhfBDV1zdDicGQLzwOjNiBwCSH5XnCGJ92fla47sd3SfmpUX
Eq2hMH8Rt0mXSrv3EaLfdWq2K1/GuzZd/f1k0Z61/WrA/zXuzVfDoFGRPRUyBf48
i5DdKcy6LwM99RA6HmMjcI+JCqQmpFM6BkcsU1Qp8PGpC3HSAAII/HcziaT+IRIO
Se0dAnx0LzorYeLFaKR8J9dHcNoDdFeDpylhzbpvB9aFuqfRnJ1MiigfcXs2CtD2
q4Q2RujpcvzBFtVPe6lF8ysgt6itF+fV0y5QToL+V+t2fb+cT4EywwuaEQyYD/xw
4kfV4nkhcCNEZ7ISZ4h7PO0BxLux54AQCBVcUt/Ev0feROqY5MkaG3xAGYHlv6Bj
QPcTx55TlmrVfnMKysdNRx/goTaghTNSaDMBwwHpb6NsIXNqG+zKOlCzXhfOECbc
GlbcyJnb+gil8vy+qxcWUnuIEEIvHtt0qHEXm9H9EHNoIcE9mcbw28pTWiJEo9XU
65ifEDNMf/rCG6dc2NFjLKbsQ0nX5zKWj3RuZa7TiT+7ErBbQWaccmqjd7uYl+9G
UMS27ax4Uu9YpJHKTpoLcqVPUXYdaFkykUkToLTn+Jd1Rd6Br9wQFLxOKCsp4YGh
n2svYl/mCtY8wYXwSfF9VMtdZkrkuPYe9oIIE8mvEeOvg8NQUP3G8Tshej/KnaAg
vt1tGwPQMf7l7aAQCSdE1N79mWleVs6xW8rJurdAhlaIo46HFepbCeYzAM0wMKKG
2JSBMFabXJoh8kEHsIlUclOWC+HgZAvh+K0WGiKqEg22cFcxK2ET0Wg/EWyV+zBD
Gq2p8Ewz0RJlIyoSUURgchsfhwCclHgBu+fAa8RsdTLjhO1Y96nXv/4TG8liyYn7
o6jF6Dui0UKbFSdHx2nHb2/ROnijik9KeWyoTa+ivWar140ZmU1OV8KHZSoViZjK
Vc5zNhhg+azA46iuKHYKkQ==
`protect END_PROTECTED
