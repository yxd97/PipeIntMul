`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SNgs6zHb7odmu+ZLb3YVERi4i3QyfSDqGGZiqsyeTxM2S11uw9kgs6CHfx1G/fWo
97IGJaOJM4o7A2RzSYc7hgydZILLLF1EC7WnLPeCXBsIqPFQpLNtPOKYGx67RuZh
iwZ9YFoYRl+NADcVJuqBnjCOY9Y7Z9OvRuHzzhPHtz+HJ3cfuEPyPdoP4GoD9zOW
wmHAjU6LAfBifbhsyvuWn6fk7ljxX2vXvGA12e/mmatzyHaaNzAgTIQowAswV5Gs
Z4+TSIkIWiyI+saJUOx+0Y+xJE53nCuKSvXipIGBtTqp67AFremb+vNEU8VHZXT4
k31YJAwD3OH76T3BrAqAT3dcR4YWZHv72zq7o6Rca1nGxH2okxUrpTXJKGAYUpzX
6elMkxzUJv868y44rG9u/wMH/x0NONQfrilmYlREamSMP2RhQTNY9+gPQATF2Y/E
`protect END_PROTECTED
