`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UyBYaVIBy2uLBDmSmbDx6zqx8Vn0n6qD00beqmk8ZNdmjpJ4N+bAYcKLktjtWElg
TfARLgjq9+n3Ybc7xi1L9p8PXwvq/O0DEv1r75J5pU8QCu7f6xJAbg+Vw2nZBpq0
NeNDjfCIqh+Xks1SA31JYTurKOCKmTS0NkoG4oXRh6mNYxuaHzhnQLiT8td1Xvpu
37cNQZQNzmya04OilVZ+aUIYfL1nw84drobFkUb8kSip94qYXwhdQb2ev1qYNY0D
0Y7C5ccCVjd5204qjlxWQydSFrRt1MguqezxTp5R08L4taNSX1GiVvMCKc6c74X2
hICLcV1ZFEDVhuhYqZHSXgqD1NSyuwy1k2RAK2ghIsNWIwFjMXVFxI9aztsWu04d
iDsW7BXP7DRg1Xiq3V1wS/3Jw6w0R6fuMFTQu8rWOswyOB+kuQnAFv1BzniJrwsY
v2kNPTOvX4cfHh234mxt8gXNbwgKYM0XJdfI2MxyEW7HezMT6EI3INwrdB94YowZ
bHsrugl/B8dxY7Nn6VJLpP3vdoKXPX2NrjFBTSrtjcVNqIaV3aGcRiGXkM7dfjhd
Vj/sRw66nuQxcHpODqozHOR/c1tj2YfJIGnJ9bbTBQ4=
`protect END_PROTECTED
