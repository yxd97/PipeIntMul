`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKvjLklvnvuzHciqhCIuNP2yTAMBXO37/p4YZ75T/OnXv/w+4Tzb0hFaQO3VMCT5
tk2eYNY43gmohNWgUT35mq0rNRlK/HB0l6tha3ERhQnQLvg93D5YovvhmGYxlqJ6
BkxfpuLousVu+pQi4SL4vRjb3ltIbjKdRl+WGOnrk8RdC+LQoPa29d3VRN/FiKSH
6tg9rFR/0hpUJ8KIb1CBgPWJYblO43ypzs3g9zzuzaJVbpFydH/nl9f30G6zYggx
SRTrlWzKhK4PtPoKXYn32g==
`protect END_PROTECTED
