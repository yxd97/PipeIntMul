`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tic/N32sxYeNxo8iP1LfSS5bT0kEmqR4/iC2VZEaVsxoYtW84b0sw79sCE+bu7KN
e0Dl3nMtvDO9vBoJx98VRv2Nm7fc+5y0vI72pGu7GpLKqWOBr1gWj16MUUhv7i0V
/LZw2t51ZLqp20mJugnrp+f7YTBqIvGqyb7ls61dH3dEkAp/aHVxDuKk0w+7pFUW
NRvj/R+3U0PPXjcsDx/kk1m3h2lDJH1iIBM7YSexPBdHcx3oqky2ZGGMwgAWrQP1
u4sFeXPCfhmx4JFX5f5gZQ==
`protect END_PROTECTED
