`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ydiJwWclTw25cAJ/mitmRtdy1e57f1UPl5vALUXgSxrR+4RTf5aYGhINZ2hNypsa
YgpxIodpj4+McP8okc6isLciXL/0wsCOHKp2PiDQca8rKzCsu0z+T6q3iZ8z1/Kp
n1m65oDBJnHoC3CK6xLFHdfipEJ/aP/dDtkXdRZgLKcHDCa2BGLWPRug4R/3GaUi
MEgxwVSlJ4Rt2Kr1DFF/5FQsCQcgEeIJH/ROo3vXAyO7ujvsAh64Mzu9D4v0f+V7
awoDHfbVxlEDa3BmmUpxUFBy99JN9hM48frchOMOPryHvrfrq+Uki009UrFyMFE1
p5TAlLir6pO+QiOjzBpUDn8RwEga9jDHmbbOeayHNCyfRxQagwkRwMeZonMubf0o
oZxHCkppK9LnvNla7wAnLapAsFM0HDp4w96jdGxE1C+qoKYJnJpbzd72dFJYw91c
8W3Z4WhFzb3gnzFX10HBCcQqwRTB9HyArtODRFIxLTuRd1g3lC88FsfC+M5xdZlH
q/27/WhTxmSrkUjzJJfWrlHDRQQT/nHZj3y27eYEp1QKEG4vKMIm1VMJod9r1Xl/
9to8bAuqQm5X4WmAYj/03n5QEW/EjDyI7BqTVa4o01SbK9Ss9noh/bTAQyk/P0VQ
OjtPmQ65z37uTZPHA54Cf+fBMi27CrevFUz55hU9dp1WAZXXls5FeSpe1dzDmfeA
niIzH0nxxJNulE34fYuBNwvh/zJYaCDpajcpjVLII8nutTdNWMU9/pHrbDnzL0Si
8KSIkcrtJBvjnJFn1KEaE+plDrqvQXPWL5oAhBbzfCnfGfCQ+sxNEae+VD0u4FdN
T4ZgpM1tQ/y4Oni/Zm/WhzFbKoATF5Y5DuDk+Uow2DxHm1Ib7DDzixZVZ3whyChA
vSGL4vUKcuMQVMJHwrBmv7cDSKfp91uluiXM3IoFq1uhvDg0c3Xc1MGGteP2cn9H
xc6ve7VxC5BpAGVoKff8o/XC8K/i+g/VisJS5r6Yc/k=
`protect END_PROTECTED
