`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oumWISdGNxgA6PDc9/q0xXxPqX84/3gyopAomj7eW8RvzrdcLviSvRc/OCo1j+H+
s+fROqdx6SoQ5UjIpJKyL334Z2PK0ZHr1/FqIyhbHGGxi6dVDz4OfHuZuVumTC1Q
x7T3m97GcvkBp3z6KAnHpjVMi5nESvP2vl1mlKgy0S7Xqkxpvx3C53Y/b2wBz/I8
+qCa6e2QgSDLJ5xahlNSaffR7OM9rHVyuZ5XvFKcYx2+sdqbFCRjvJX06laOHLc2
xaMQBes6IodlHlo1i4nxv/QdvH/xvrR/mUxtAoKIm/ChrUDT+JnGlXaeOsF+crHV
l85nualETPfXgazhzg+EF0PHIv+XvcIYdnXak0q2n5kUG02/5rKrvGrgqaJ0IjFZ
dBWqZWXn0dKqL8XBe8aGCyJsre5pdkkX5avClCPo6/unjsDSVupCvNDdoLkSzEtd
HYaucXXWJLDmJTHXzVOVEvKdC+6vpmfobo49SDIo2MAZ2dDRqfeSCfi2BEM0S/1b
Xs5KDYGNV19HJcmikDVgAdj2FDWZVyzd7CD7uZdNKBE6uhZSxQfwuiLnTVaIJCsP
8pjHnF2wiaBGMqQFU5akDqdo8l24o9JyyFOI9MQOwGrteC9aOsKwuYJ6no+/MBT1
DbJgM2ADHSomvXeERhPGtaZG9Xr5YBfrr/j5w8+sqGPxCwEduoa66HeNrwwlQixC
bIHV07b8XhAqAeTIpu3HSUtU6gUw0LT/iGjPWOmHA6pHMZX7iZ4IjaVmH+2Giw/D
N+4JKPIDInmCKegMnWoqpQE+Myzi4nE9HG3DPJ3kFJSUxIGofJBJS/V0j/KIoo+a
NwJLN+Ea6frvPX8Y/FKnmZOgu6keiNftOLYNFwLcXuiekrvonv8/yLvffjgbLPr7
DiXoUhz83UA9s93W9F+P1xPABhGETwDtwO9O3yNqF2H8JwXbm+OdQ2ZiANX17ste
zIreB+kwMJv1vIpJQ0celzMZh0jQ1rpCAiuf+1cnV26urm136cYPAXFaVt3f4y6H
fFKmJnyw0z1OdRt3Iwm1CjjxilSQO8lBPpSotNkjjemNM2EZBHruGZ/ztPR8DrRw
coWNDmbfJzbPhPc9FdTw6FO0wIy5seZUGx57UOdCiNoDxot1nlLo0JJcr23IEIey
2U9lphkLXVFDwQ6TpQUCW/K8CReOfDFz2Rx0RDOVK1mOq7aES+KwVpiIBiPRFqPm
SO9IRku67yMl1fYphrj6s0HLhAO6NMX/F+aoIatQkYwM7QSmFPopjCQ5AR28lX79
mBb9dd0+iX94FBnvtpWgMm/XOqroBGW5eGUJA1l7PStTMNfIXnqHX3xO+++C0ZDM
NtayWKf+JzxI8Qfl3rXjEzaIpPcKcd3348pwEgsYexxbfBC1lp0xUk/1gl4Xoh2g
ml4EKrL7BvW/R6sZU+TOgvzRwZo5acdD0Ok8HC8hy0aj9J679HdM/qv9yxfBboU/
6V0vHnLl3gW7SZ+KP6d0BFKp+TdxRj911JBJEaJTCJo+TDXC7JZC2iP+dvHAvTyA
ebNEO1Sa5D9bT8XIJk4qZqPyWw770//v2MfxWWQXmDgPa+MXzakrsqVfSg4OlUZv
UhWu9AZLhna3efK3E6DTH4YxlEChIDu9GjyiZRuRqSzIV06hw+QNG1P6XRySLXZp
8QSSEgngAH8Fn4XA0czu2AFJ9McjXKBiXsI4d2Kbyo4IlJzmejSJV6WPAgzaVTyu
M0QksUHtZRIUrzIhjMF9RJj5g5Gy58SHGsqRl2kFCIKgUpRArP8bQqu3nt3xQLEf
GMSAOFpINdgAd8YZM8+aLGUfIlQph2LVerUfO+QbIzb1miCznx2Gh2mY3AwFUZBT
Gkk/6FF3KVRaoc8dogVN/zxqghEW8pcYwX1WIAUYdc5/Q0df5wfkwug2ZfXslPO3
UHpaH5Z+9pEttBNhaNG3WjFVFuIK8WIQds8O/qFEjiLcMZBs4jkLBR6Jf7b1NDmO
umB2izMPW0X5QZOsDU3n37ZeWKAnuDpU0qN9YlAxOxcVwvz0L/PwVmNinQFZ4Dxa
nO2GObQBcy8ZKUJ61kKNOTPb/RpYne9owcjLhWTP4rrl4AlHIFjC4yTtfYvLgEur
3eMUVTwYG4abGc8IGcJpk1Q1dyhin3aiodMBB2vu0wtHWlE8a1PCwV/Dgtw5xRMI
Ks5Iexj+wq/TqG0qKCEy3OLbCC4w8KHIp14LswhcYT5xAslE90+KgfbnVRX7YCKj
uTSvU6TBdOwciYNWjik2dFB3QB3BE6N9wcqB6wR4n8mONNm7uDLEUplS6KThw3gU
aNzyT/afCZbv5oeuT0lLe4qoIV2fWbLSYWM/yIEpwGg0CNRaKaS3RtjNbP6sAanY
8imGCByG99Bbg3vL2C2eMsA60ZCTEvRWQQXFtlQGmffWhYBYg/8Be0O9fA9Yt1vS
YERqm337IMatfKoMv0nuFlAGrRVN0J/sbd8TLDfnTIlhurJU+sx1vjiHC4S3f3vQ
VHY87PPgIkSd/njvSloVTNwB/S/3xd65DuQEZq1fSsa8dm+VrxtvMhSMd8/SgUvz
thWLCUDa75Q2Jlw5jGMvV/yts95su0ixuB7UEowKuAbaf9LzhlJFnJGwuojeQk0R
+dW1pCha4BNSXLhd3IMDt3jCDr+jl9q9Jwi4mPn5gDyf4nXuuwt9klUUiEJ1tAuO
+X2AjQtQFKHj+MXciF5z6AJPmBgemwnyDeaod8Ra4jo9aP74QYdjlFzuVDukaf1Z
G0uwny1BXOB60IaOLzvg4tZEgwc1ej2rlDgOTja/79xeWIlQcn7pjgmKyY6PKd35
EjbajUsRvE2dE+syp79MzJSFxCZ/q4576b4IOO3m7m7iGImIXFd4VDy8ldxuGYsR
FP7QSgG+ApBEidF0ojJHJ8TAYv7n83CuR96H/aOainqpcI3ETxS3aB0p7uoXjJqS
maFw1QR2uvd+ieoWSNKS4huAwmw/xaS945L768VA4DEDjPM/e/wXoUaZd9xBdnr+
Tc+QZFIxilPC85unJ/+c9FVYzvHvoRdM5rgpfKEsdyNnc9psngg5mPpzl7//yELj
/vpwTT9dIDqFOa+FFb1R5YrKIIIA0FY19pd0zdYUmGx20duQoSnU3MYYdDkyKul0
ogjNgUrkdQzNmOWbI0go7WdVlbdG7FbUYrHgCes4QEEo/17RxX7rnuiGoAOc8mvP
aIGKe5q3T/cG+9QayOZktLsi6WFUkwIoEw/5/k2H5rNTrIU32/RWY8rS8l0o7KfW
qcDsk7qUr47q5K+wy1OODbpgfpaGs+9cjY8jbCX1dXrvc21rXbEgi+n0UPaxfIUr
emoUT8DvbrJmujADqU5BvE1/uDBkfoS7NPUxSUNk9rZS2VnYzUh4N3qhq2T45QGt
xy4xy9t95kdJVXf+AfVKlDW70QptbGOdcxl/WcTHtLsduu9JibC/vd/q+mrWO0i+
jlNsv4egatWa8eBoVC5VrjgCFYOx2jA0rw/ZcTXj2JxDpJ8fSPnPd20mcJUJ6Nis
SYFXiZI1BH4khRLVQCHtvzP+RMFJuD69iDm0d8gatFaCswoVLppXxXOf6LHBdyY2
xOlcxUSgKPHDQofV+tbDFlkd4yQXdklHv5VI6AhUiAQ=
`protect END_PROTECTED
