library verilog;
use verilog.vl_types.all;
entity TIMESPEC is
end TIMESPEC;
