`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Og6DeyEqeikejCfF92EU3zUirXOQctZqQpIQRU3QCfinAICE3AZdGyzFy/8C1KZ3
PP3ZUfBgZWQggVTqmyW0Y79cF/1JmNZzO4Ww5WZRkqZ9Nig3UnFB6MOJLxyiRgeu
/OUz06oosuJNpnQr3AJiT7vJTd2qMGb7Ce71zEJth+Btwf9hvhfoGEM36xCypN1u
imXRD60rcVkDdlKryrO/9HJIAygjTW/Zjdm1ptm+vBFusuRI6JvtXQs4y0RIG8XY
Rc7L8CSH6jLdEZD98WHN2QS070f2Le72JUfVB5GstHzbfMtRZYiny7nvdmOHnrwv
6lwONFpP2buv1g8UEDmHL58sb+rpdgBLZsDG8ppovpmgtdfeJVQ6Xr3U8edn5hin
51sg1/k4/wwjD3DyYDJrTv0LwVWAeQkXJiCZdvUD7XrRcXges3WDcPqPL3dp2JRH
`protect END_PROTECTED
