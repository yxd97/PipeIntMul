`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CVsP/Q9kTbXiDHT6onPMExDPDqe6flT2A29CdPdL+DSw8Z66n4I9thDuvRL0JnqW
xcH6h+kXUFVfe9oRhvpQhifx7qjyjwttMz3uTVX7K9Q7crx3H60xAxORELeYkLJg
OxfQO5ljfMV+ksELmU6gWhW5nmoSj8dlq3Xsnyuu89NeLJxOJejXel5MbqOuROB8
EJHFoHTgYc+7rl0kBMrDWhXRBKUUz8Wq0CVg3cx7PN1M+JttX7Z+FOxZblhLhIgE
swwrXg0OCaGtQ2W2w2F+pBdngA6fTm/0hQ5Y5MbYbEWYshE0v3w+nQCP4pfduMsL
G39zM/JFORjOuWcNZYGLbfiPO+j8JtiEv9FiySsnHJFj+9nDjxfYgdMlVjikef53
yCz5jKp4SWCWH21t8W7i1xGXj7nvz1GVudjTpm30FRQr+j1mQaC0t6jN8iiyap8F
S80iBEVQUB+RM/EzQSesQRm6UZldT/FZfO4MKa4Yz9k6frZ1y3xH5sYKXzAOTVH/
pb7/lmllUfg01Dz+oCfQwE5phbk0Q49+rWtwqLsVNxbRpxYIMY3pVXicMr8iGva9
pW0EKilT2/CURqES7oW7J11tTSCNUCV8AR0UlIYqqM8=
`protect END_PROTECTED
