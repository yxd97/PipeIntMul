`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HeWGqj5jn5+t5gQBnaEMEd7zCSv13Ns2T4dyd8eUN7O4FGX9CAfQ8k8geeOzvKFb
XkzVs1CQ3a3q97kyPfZhPXX7/jVUBDYAq6nkq+h+3kFYWMssy5Qo/zqEySjUcX21
en0AgAc7tDPVTFRdFStHrjEEHlSoJ2XZC0S2uJDBx8lRqgIJkkbtmEfyX7Nkc7mi
jwO2HTq44OG2wUGj1MCPA2W3tMhZXz/NfEkpdH2PoyDPVWzavv82H6IlQrPrq4E5
vGqO6FiS/J62ZFRh3dfB9dNu5G3uf9S8tKuWJzFgDqK8atC8HYzIi1Ja4R2I329T
889zFZirSJ2Im0ij+05hcVTYuz3wyUvzt5YCKfti2vBuVw1+YemscwwGUgsBKpCr
KqaTOLcI7oRQF8TnrFAanZ0Dy878YRVEolaCnrdFS1PyeTi1mgsBdXf005FV3Ykv
9B8/QfROJ4M5NJW6vlCv8rNOuB6T+t5v9QCCsUyF5UH4c1DeS07WRO6nWF88HKh8
A4G62pKwQlbi8OBCyzZPjlULLUY5pWwxDRxbndNh3hJHwDLFydJAJe+LeYqfbYg/
zh/xEnFTCxqBw/+QoVN0khyDMqlzHiXL9Ig06CSugn0yi79ZlB5GAkPiwqdNNRz/
JBGHXgLECwC6yIIOY88f8+j0fFpPTXoQEButJc2fjbD4dy/Hc6+NgtMfNykzW6wm
uLwyjwGQ2pPWoN0uLUNCaFRyEFmIchl69wSSi02GHCb2NQ9dtxCthYj1PTuYoLw5
0WnjPveCNaOGIkDVuFnVha1SGxrt+qNb1AedsryuMd7FYqhhgFUKohkbtnDqoHmu
FEuy2E/5K9oP9CHbtp9xVDMoaWY6YtPvOpig5XsT6v3iNJVAZlNpjxFlXkdKUTKJ
D4+YDefwWoAyyNmAp3dTTWK1XNU84i+BNsJxkFJFXKT5EFGiyPWoF82NT8EIuRce
E1g+P1cPI9Dl8e0X9KgSU8+9vVI6EdkIqbPs4O2sut9AMiNVDAwEFH6lhPwtCVtY
5+9WVPjNCOpWUG3aEqPJ7jyqROU1+DY0NhDetHLKZYtUIra/+N5zNgvVvgxuEsVl
FYOVob22w2HCfvFJC+ZA0amEQVHu4JxJkRP7TYZyPnKFT+W83BsRgf2wt/Al34mG
n5tB9GoNqiGqKwPQ+tEP5oxbm9fFLON/e0glruw1wb0EviCpEOjbW/2OwchDeJrT
X2Ju/jjDcHgVCE4BHLjrCCXPB8Qki2hVZcZs19VPdQXI7wKjEn6liIipgyyjQUYD
RXzm22f/fvAxwtYosqXf21DSvT44sqILIVDf/+2zhsVeZI+l38KZZRNT3bF42rlt
N98YAOghvOaWn8ebUUSdgn8PVS6AGn8mDqVVwAtUt06NiLo9GGIDJKayPvBNEZ6g
MRgWday7gJ6axoFg6PIqkpT6M7p8F/GptX25I6DD4HFQMsLYRRTzfD/ibpuc6NlF
GA1fDPQSrDgDFNRB0SaPL3BpsJrC69bjzL+DNACNgGzBYLLshW4elAe61U6FaCK0
UC5wDGSxwyKln7+NpHMm89jia4uaoeaUp79WzPx4gw4BaGPFQJUmCKnwPbjq9xTA
M4tI58AMlUuFpuf8SSEiDatl0iV3SwVnBPdiD8LhmA+FRYXrlht4L/foeb+FBZ25
cTRWu/fbQTG6PIBKc/HfGkCiNgnBE+aiKGTpJoU8XKjKft2DKKa9wes7Qc04Qyui
zUmzhmLHQzI8sU8gP1ozr3KXLPBOT/02R8MxfmJ3E8L7TGJh5NYHcz2kmayRMGUd
LypTpBZz6kejZbIG6Rt47I/3W6+5CM76MjI6BeVzqGo0rKCag61QXkRiH5jY9DpK
0YncX1/apStGdCJPaJCV/tfcEwXgTsBNMtBzKc6PHfYsgLV7XeILnUXxL188ncWC
SaVWISJJBeNNqrIRFPC43cILaK/hqKMY/ALk7llMZMr8q2bfti9d1TXJPZM5ilwA
jsJKPTGLa/SRHIYQo47AkXbWGiJ73dMz0Aya8CGwIhrKPDlFKzUb3edVx8IBZIgM
lQDEr1kdjSsh9j4uyS0xYG6He7DVih7d9K4O+RlTSmY32e3dkX3LhPRJ8nmnyzDF
IQXxjaupstV/TZN5bhYPH6sn/37/XwPqWw1DaQ2M1y20lIWw5teotBYxafR6Ugh0
k7BqbjEQE2QtU8QXqJcBMsHDe19gW9gDxeEG8cmrSGKRFPxyY3eonxpeGN/eSg22
ADacrYA1uqaYNvIEXXNTQCH803qQSyRfC8VCMINnXZreQUGJxrjnEw4Ncq42b2XQ
QBiekicdlLZF5g4s/JHU4ixZezqEKe2V1FO7wPthXk/MVVFDGEClURz4NZVQPPE7
wsM27hYiGc2g8J76G/uziF6IOLErclusOeZf5K444qlgh2gj/LDu/v7/uliHOEf7
nBaqrbj6BBqVDcLTjTh4aH7A56HLyOG4+vBEAqxi1p6aqjm/PqLlB+WNaEP0vrb5
ZFCop9ReBFxn9jV/qVBmsUlNPS3qyxnDgEsd059cpObJg8gRwJvZU9wxa3ipiSFA
pc9iF05/cLuQzZeI6/Dl2DCygP00qoZOGParMUkYZwsBefQ1RiefOCWqQJr8DThg
AVf5rlNbkyCBDP1Gh0uI9BfKjlbj6igpn7SpeNCziXy0qrcCCjw6HiL2tjAl02/h
6bd9W21SaVlXvo/t6dAlrpcKMwWSl45fSclfYv4FRDg/yDDC65USo2zSH8wfdiuu
V29QlTMAmDJkLRArUO+dMc+M5YAulnzqsbTXX7J2ZEf8nmAuy7OZO+FCllC0la3r
U4oNqSeUX40RkI1ULOAWGz0qPIOvuwYGD9qpaqw6hIfEV/ddb3uag3ThsmIGsAdq
YUPh3zC7fBEs/9JVGGsH/S3Uy22XStIkr+Nw3v5HacM8NTctVfJSbKyGj9pl4YZP
qig3ytwNEk8ICk/Vi3tczBXfYN8nXwPnzl7w2PO3BlGU1J1L5iFtVBXMBYZVpoWI
K/arBKoe/gDSdj3MroDx4f4FMRlnfUdPK2Z9AVeTJeeKy4zRqwGU+fMxtWM5xsiG
Kdo25A5dOsVp9PX4xtMhgID+67/UOk4kakMdhue3uS6FvwSB6fRnyWFy3ClYnMA1
8z4eS9Pncz4TtbxkUjkD6jZ2yOknp29l4m+iI6ne8pG9SwIev1C3BVclFHyrxvbz
D1gnz1zxBCVwCpP9YlEAFoJRSPknZCSBk142pW5K0mjtdXEkYDFhdaysstxjexfj
7vU33BbyFZDXWiu9v4oVwcx6KAoRoRH2VtmTSitbQRki+e7yQMxYDcPJZfM359dT
zOtXiqr8tRcPBjK/XwI2abjFBgHPTBjT8l2t1kOvsJl4XBQO1vcB+8+YEgPZ7QvM
aBGIpI1KMCm7KiL2rfN+VYGN1ue4lO0/F3I2jsuyso7y01GxCWnb47YvovcvlgUj
NU5g0dww6JSkgy6JrQQVWrGGDc0bJYg4zZIYAJeEg6zkcSQmWzi82sa+llWiglsa
PIGVqXTcmDZNvzLxEcNie5Tn3+rry/L1q55calhpB604i35wbY0YWKnJHG9e9dDJ
RotxGj5EZJfEQsfEkAE6Jzec/JI6/N6ZjSYycXZa54uvgxCKE6Gl7iv/N8FXObRz
D06BUp79Ykm5PeKSC8b2YAnO3IrLKQC/6RWkhotdsmtYTCOWPSgaOtG7VEHIsZfk
FgY9Jhx4CHHqBtD8D6Iw7d/vx6LgCWM5jEbV/tjdiTzPXd+uMxjq3icZQDEWtJPz
YQcQM76W4EMLT72im4ofiCfS5mtK78NX6of5ejIfM/jcW9+6Fuy8tG6Lf9otDw2Q
Uxvc8orMYCS2DRhUB1SyRZNAITGTamUjbjXIp+bcihwAkestJEVhiEBudUbjO7i/
DJZi8mdgxWipLmwcSpJs4nAFLLLi3Vrzi//7PybKCVcwhZf+4uQLAichpQSXA0hA
HPSIAxJ3zqZfbxBTt+bYhZkNfGRS1/PHCObAdBYpCoQC+mmDsUCxx/Dpg9o3QiLX
OcbBD9bSlFJ4yguYJs/9w8wFhF3JHBBFNWwR9GiKPklKdG/Teb0LNA7OOXI1nZWA
wUVjBhWICYofgbr2d/MZ9EOFgL+xRpQZQDM8iL36nyKbtY+896Jn5byOpa7M58gw
tEBBuX5qIOD4OYazoPJ7STZLEnzeoVHEYka/ZRPesFh6L9PmE6oXxtuP7IMj+j4E
remV+0u5xeCg9DKC21Nb8Yw3tbEtbC5FHrY/FI45XJbGitvjnzI0nzSX+rqynytG
QSoqnR/pnpRiYAW4y5FJu/TnqGGqYv3xJZKXKchYQGUnB5dTe2zsfwjQlB/GceIU
z3wu//iPxSB8q1/FXovKHhTaThuFYwDIOdhMFrOIR9Fzj9DR96MOCvcfkvdKxnFr
aAY2Mtwz8cPE01dsT5o3lB9BpLDIH5mqPXrvDlK0iGy086pSzrRjR1fwM576BXMN
F8Di9oePrrugeFuEopegvU0mrIe74FXxaDFek6G++TBC+aZQ4pBlmZ86ol1DkSRf
cP3RgaYIrU91DGcmFnzDeN40utXlzbI2K03eHuclbJIGCbM4aVH+vLZjdDWCTALU
lO6bdn40NyS9dISuXs4fnJy0hRyl3ZNhAR8d446Uo9LpjkpmcNYkbz4BF/4SBR1q
qmMQJ5j9VkAp/otqlUL3WxNpJsNzNYeK9Iu/e4I8SfoT7RWw2dVbroSx6QTKAfvU
CF2If8Dk0hhq5rR+fH8Ubg2NmiBPIRPdXc/qK8xbdyCRL1TdvUeCZ/k+jGuAd22/
9KHs5DWKKdXaoGxue5o/G0UBmJ+SDCYTzyghM8zm+c7Kqi4OQxBpC8ARVjdrFnk/
PJR2HBBhp2qYYM3+DvDTJzHnF7+dNjYBCoHQp47JSeYHk7x0J8Xbeqgr0pxhxJd5
yc7Y1ytFDgy0pMOHstnp+8DUaKW8csP4NpBKwI3W7JNEihwQqTQGsfCcjjZsv+Rp
2mcL3kPzHkVGZlnvxw1MX6hXoSlxXnw2YW7tC2N9iO5pELkuMESj/3BXx7K7WAG+
srT9QboArU8HLMAJ6vOaG/oNb46zLF5zK2Orpnb6EX5UMl5u0oZ7vRKnfbO5ODf+
x5RWw3omNndERl6AJ0rOEjfTPfe41HzoiYPz7DKWSf+aCNeRKFPcjTzCimPP1c7+
NpqajS5khUn9O+/DbqhQiWcfKq82+75wVgm646nRFAMKrRq7ETZwX8V0mM92jjKt
Xjz60MHTjh9prPcWjxsFwOKt+LCkSJBNrZZACDAyHC2rcPftXa91/xWCRnkvdz7+
1Og/G5u8lS/eZzqQ1y22MmL/qQaDO28uZO9LSpk9/e7WNlIt98USZ5MYh0sg2jKF
c694lNGHmF2mXKebIqrikz+yKliBtO7PcCzD1Hc41Mg1z01VQw1iGV4iNGjxPPuF
sTF1Wjoi1oMv2HuiC9RLZlpcskw+ovqwg8IUcGCYBz8yAnO4KgmoWOo/cWNmWlXM
UcTZD1PKBSl8LgMFXWsy+yVu08Lhpu/e7m7a/buxsHI0vyaIuali9ajH/H+E30Rx
A+oC5DOUlg+4H1q1Ch3M/OlMmWjzpkb3NtJKfjk9ozEmPrRl/TGG/6z1SBK0AebZ
VH06ULmSd5QPiTBey+NDk2A1rf7T5EBWSZoS1XbUi2KNbb/8HIl76nsB501KYcwW
ISCELk6GSG9VyUCsVbdMM+rQU+6YJme/KISRjqbIQFUz+eC6k1eDLFJKnpB/a2w1
dfm3XzXtLT8ibK9guLmypyiNMdGhTqDYI5sCUegPlD1btOl2Quyt/r3kzp/ML1wc
GYXNdpJJR0WzRXDcv6qqPepe+hyHifKAgiww1gxBx0TVoqgR5yGmqxvW2HrJJFLh
tixS7nSkVgTeBZZCZg3+mCS9hZUcrks2/+bp/UyPZifsqkkFXOLEhkY7VvZ4eoSn
jMXNp94pLpiOvftPkfA+E6LUuUW6M4bvGYMCntnYSy8Dp9HX2k2VSQFVJ7R//jqI
vp7O33tqrRscN746v0syseKv90V9lE0oSCkXUYUcMU9w6+FG9mx1xRC/hF4ScgNK
YEb0tpp7kOMZ4SyZBJKVtLxxKPD9cDzL0WJHzLJHxlKzMfAttdPt8KO49wACzjX/
xhgz9ByVBVVH6r8ShSoCdK8ImkMF83spQYde4kpOjKTLaO2ZrvXezxpaHxml+wt2
qqj1bX1dlSl6Q7Wl2lJp9ygG0EUTxe/FInph112Q7+SssBGOaAMUFA6cuqZFAnq6
kAHBvKpzlLtFJykX7vP9dGhoKLyxt0CJ+hSRJ7NFPmCJzP9qHW1WccmQKfmI9Zgi
YWh3BX2k+jcdFknaCfCy2WiFPzZDdZQFFOKE61SIqUSIUtaBprIxTF+aCCTnkcMb
esTK6TWSTA/2Xo2PdduAa3UPc+aPUSyddYM673qKrkwfiUf6ufNb5DtaOxd36130
V/Ih5XvkY8g6dHrCrvKHD6ZzeaRV5IE7wuSla7NzboaRTvTzC+0XE1KeFb/Jk/62
PuUm5mKvSDAfXMccbe/VTvR0yP18E6MKfcQ4Hr5dW9RR9A3EpPYTPHqBLfYZphbC
JD4AH7pa6o+IdKw3R3MA5Ci5Sfw3MNPtYImKqrM6x9SRQJg9DmlxI3g9m8se8jI8
/bmfZ3+FtTrkCQ1ZBPBwUE1SBgz6tcMX9rzLleyJ7bainF98vSWLDXWGg67Lu+C5
GxhPCgun8qDQldTyxmz/8aQhiT0o6pLS6F6FY1INgMTO5eS+a8gR4RTVjiX9llhr
7lAR9SKW5k+kIOcEAwYnJz32KTun32nQfVYcktzpwSpYYC+2HRDPHm+Ss1rBZGMa
2DqJlyxNYVmiKmyY7aJt3GJNmsoEeaYP0QUu/WeJgmj0rAHQgvpKwFYk8TT139Wp
HTV7Qz+Tg3OoyoPEv022hzBel85lEwcu3r+l40h+tpOHdZYhZlF2E/zvqSr+DcCi
`protect END_PROTECTED
