`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rMRTmvoG3sYKj4q7AA31ylfe5qURF2KoVMeqYtBzM2cm3QMZyyaQrNwWMfUsB5iC
UYGjHR2oUflVpwj9e+teuWQQA4Xn6g6L74gNoO7JkXiene3EBiY3LZ/VOlkqfAyt
902sMcRYUaHyugivnmmNTF0PSjOwoptbq2RIKiDY3C6gbt3gTAoRwHJpLWQD6TIQ
xGA/jsaD46u6yINCbD6nUvBH+Cx6qxKOpxP6WgjRPF2pxlq8L2JaLUqQz0MC0TRu
XTymFWFc2DICdBG0hzsCNHXJeYQmAw06nUob4Z72dHX7818ggnve0sLkqNDO6UjX
Jgh/4tT3uUtKqjBeZjHAaAU7sgAt+zigbZaBGoV3C1TznbeFuTmXX0ShHi7TBRA/
4g5cndix/ccRmMYSQZ4Go9Io6vnP1Rr8s+X7jz6/kc5gX1DwoyRTUjzZB6auEAHa
0E0KT4SISG2+BqwzIIDkehlqmxQcK+77yDaMB2HGsf+VLZYS/jmKBfja9E+zal6o
q03YGU8vCpR9KP1Uf6JTFiPHIh57YTjuiMhhL1ZePXo=
`protect END_PROTECTED
