`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RjW2SC768ZmUegqWowpDolXtsdy3lH1oUPwBhJLfEMfuy798Z9ro7gOGn/k2DQxn
Oz8XE8CmXNlYgNyikpDhD4obGRiqn70o8kkYZul5QcZMFyvvU8qhmKJaxYdmFbwB
Kqc79jF5JucejTxYBGjU8IcSQRRlCQ4y/bHDNsbxMEJfnVWdH77sJ7zPKVQl4JqT
t+SlK5wNyKs6g8TZ+Q7tXIPq/pILF829AzEIYfcRf3Qhkk5YYUWZoWPwdyCk5AG9
1TDKKeSp2OhnWgl0OGxasOf3av4I1hfl5nYp0BTtI5QrlNnoTwTz5SXW45hKGKKE
tgai4Scx2Ez33TTdw4+2BDJGmAlUFw6XRR/Zb0z1Foc84+XBc/HIvhHqcFQHr6NG
ykUR71UQTVEShuPVUjFdgl+amhyUQZycMYxvoJ80wqCcVl7LmxvPLLILwLV8NXoT
`protect END_PROTECTED
