`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dJgBRAtZuk4vn5o+itj73iGkV9deh5OU7NnchkfJ4FLYhOrFOylbRPNBoEteroiX
TnU80BEIvfIT8GzgAYdj8oG/hBbUcF1a/bqlaKcfa4mMUCcspeI7cvqSEZv31F7x
XiNBfU1xWG5YN/f4rTOvUB3go4MwbG1+Jy30xqoSlfCwRfpdOnZC2htVqflbQ6JU
LuSbNRJV5mOdD7h2XYfbTJ2JtfgtAKEuZyoKzF2Odssh5SbXoaEPWYqeRUUaaCTV
6Qq0qgX61DClxU3+2zeAnOYYbHhm7BHm9mR14KPVZCdvBbKFmtZsix0himf/2NAo
1BOku2gCCcwYZM8M1IUvwmNMIGV1tdEFb5DvMGLeM9m/dvq6/X+AyKGeGPL1IWqy
`protect END_PROTECTED
