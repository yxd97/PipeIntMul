`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hcjucN583lRutODna17HhxvvaYFil/Th1y0RqW4124N4Iglzb6nXQBlk+Yr61I77
1zgwjJBSUjOlwiVfViUAqSFb+fuq8VLcIPRt7484oxuUcc5ey7bUmA7dQnZ0m8Zc
4Wkle9Frv2D/OVbAmh8bePDNdWla1813y/nM24qyfgUYeSbRTeYuM/e5w5SgqemB
bfzmRjsZ5jmgvJJmn2kBS/YVCVrQskdkHtyvhh7pSp+Nsh/8TqP6ggneLqLXKbHN
/1LZb7spdwblUIPLx2UB2C5ZBT/c6pilh55FUsVk4zCtzSZZqe9DMVEsXnF23uns
bunAST6jHholzHfIZP2njgo6ATEajBDBa35oVqH/XPebDegVolQKSO/hg3Hprl07
3vpFp3FM6oJNe5KdPhJvUN95l561K3os15KYxv04pRR7EnjMyAd6qXc9jCnDEfVX
OatNoc4bPETGuun7QdZbLSbjqv2094XQC3rkm4Lx8yw=
`protect END_PROTECTED
