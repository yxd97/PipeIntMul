`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FHTGUPC7Y4O7CBZiQZPusQcb+I2Rgm/aspcGPSrrcS+yrP5qhZlNOQSAdq95RQWD
liBC1xMVEJykglCTUZCTuvYxWO2WadLcze64PAwfNGVVDu1riDuK6bROAK6zhE5j
7SkzuYqN18xvUw8a9PSzwck0Fko15NcBO7qeK6yNTellmPX1u5/s24yWr1+Mhe/L
wSlysvfsmly+d7NzDrOsnte+09TELLpqQ7kZ7X9aDCYnu5C0Jk4NUFmVPnCxFyxC
4LHRH3YplLVQQKHGZnwx+fjP+or81fsIDPsdqzCiV6PEEkZy4rFa8NauoDHc2viC
kA2m7ni0QFeee7Sv9SDTO51F+e4eam4Hqk9W+5KnNFYeLu/+e8ltA0ShsgKSIcMV
3UUb0HPpD22y7EguMrWNZVdzTrGZIjxbX+KddP8YZFJlvNJBm+4aorJ1jllcqoO4
`protect END_PROTECTED
