`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
X+lIeJyfsXT4SPW53muTs/A1RpH0Ccr64OdSpJhXR1MELJsv4suVKcfPRzMOinxE
/sdwRMZ9h8gse/a0mKxRt0k8qm8Qfpf3L3NFL5xKcQEu0eo3026PvDP7+EXQS/yn
Ne2pG6ZCit7yGAGND+s0Rx5hLSjRkeLFexHgkgwdXfWZu0BUfBA6Z85B5q5ZwZT0
Y85w2WaYigR7n4uR/3apAhtC6MGccbxYHhfWxN+P2/75UY327pxfmmC7NJiU2Hdn
gKQXnHLqYB/5oQGwJLfAFFdysnwqKGViJ7cYPJ7PbebNku8bT+i3ib1z5ATmCxqK
D6KxHcz5aFf04gYG6Ol5fYLNbWhHFs2O0cLTryCvNEcFgcB/wRWvsvrcp9uiblnd
GeonCgpCw+tNava16/3qakT6tvpdl9Z59tj3nEPs1/BFWLaASf5BVstle/0ZBC5A
`protect END_PROTECTED
