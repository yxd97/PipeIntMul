`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mHQzx/5CimBSRJ4SVaxKQ8n/Q+ojiWE1leIo/VPMTL8i+K1CKC/5IFDUc8YO4w78
lIZ4ifDGzT20DVV1VTtBJfzHpWfhcf/WmIah0laaIuJcMeW107cR7d5JnxG4s+zp
nhhWiRJkSxE8nlqYHZVl0f7dJ9Fse20IiFk8vT4yfCG2Xi9aVN5Uo2CWliNSgV9C
t0YTl5qnDY0bwsrlw8FB5LAaed/aQ6esikXKY7M2K93ee08dkb4RbyHBqPQHOxTo
xAPCdVACKrxfcC26V+PuvJh/YgSdoU/ta4RmSMJKpCDNHK2fMreTQYbmY9sBRk84
2sBVOMg5B0Hn5XEHmNv5ZPnBxMXYKkKLYU7YeXA9FD5MpKA7n6n8KR9ekj/Kh42b
w1nANfCD8cadLzarGyRoZPi1GkOOYGOtRZ+hxa5hXTv1cWWBQ+zvUopfdNpK9ego
otp5qGUjwaPAYqBhbRZXy6cUcCfAWfa/055lLcDujUYZNZL65Xja8QhLHcH26RxN
MPSSG97UAzwNnBWVg6gsPcpe15lPhJ6OI2Dvr8p40LotCTQWfOLgeh6r2R9zL7jl
b/nKUJ7ClJGgaUzKMlwmaQ==
`protect END_PROTECTED
