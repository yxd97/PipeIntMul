`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RrWqP5DAT34N8iIPkf58ROB4E22LUsAGlYvcysAqmfjL7c+2jP2kyEhniN6AiOa7
t2JxWlUfn9xyroRZHUS+rGsmEXOGVJT3pDrp0qhfJb8PL0i3dpwr/cKeswLn00mY
f0mldXJExvJZi8EH1uoRpRUxJdXbWreDrAowsmQL24B7hXKfmcfuBBEP34qDlU9K
GvkyodunwPVm01foc6THGFsfIZ8g0e5y2yXTkyJAGrOwEy4e6/B7uPvD/5PXj12f
Lfimgm3RAiAGiece4WRruJDfLoO0kR0Rvn+ikCbVr42Gz2gS867BHI643EiTj5tg
lnDsPEu8MUyQVBsqxnqCmWbjHMj8dlRaOtHd/6tDO3wxgLxvBzEPzW/xjBkFcyHA
`protect END_PROTECTED
