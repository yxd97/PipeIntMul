`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y9Ux5p169II/wKg1ufpXkCLY9U8ctvajhhv3AtevOba6Pi8BYEjXTz2DBrl59zbS
rpTysYs0HmKLKWMudD4lK9cHJE3Bnm9B1cepnkirdHo2s284qP/LdjjNMyctjrU6
pYrj4u2V1ucgbbp2mdTW9djdlaBxkT85Mt7BBDB4g+rsdHfiq04Hi5nKFlK700za
ix41F5QFHzqzBc8/25Jg6U5IcWoUPh67MRMHikFjv3+cCixky56zxE9UwoCH6TE3
VYXxfaaSocS/I5kttmiZS2uYJD39mADhnN1hR7GvrvDYli3GZGP9mwF1F1e2MmED
tpyKA551/ogOVLBDfz5J+unJTyJszcXOOatPoTecPbek+UePf3ZHJifH25e43FZr
kpHLSb2qQyMTGWQj0Vkbp8AGKU1PkaJyXWzodthKXPk=
`protect END_PROTECTED
