`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F2yPEhnY1838sFu1QX1fROTdw8DQ4v0bycjre3PwMoEznL9PRJQrFeNvE35UTV6L
aXxeSBEbVAsSMJJtLxRukcgeeQUtAU8WCATKTybud9ED700lfbMP0G3BBUK45DAt
Qhe5i7sBUoLG301ZwQL7dYosJ6P1oXbKoXVi11n1TbJSf69N6ro+0A96IC8HBvZ8
FO2H5FCNRaCjlTBIJOTnuNL2PLmamVLY3Cy9C8MtO5yrVjtXkGPqrcDDEIGxR592
KadHYA5t8YtEuXTZSJDeqnJVOWZvezUF77c8c4M/DARix/h22pX3O5Sb+i5wiUKn
TJWBBFRPToMg1mYmIOZeso0EZOyoMMZHHR25UaE2G4A5g6tj539seE6+YwCOYcPg
xWIbZPNiwADlNoSNnuwAVDsXk9VZdJPCSNKCS60xnun760ARzJ0ag/eM6QjI0U/0
afvTNhxXJapSnQwYVVpG3mN1PWvifnNCpTVY587KwqJVyXkaAp9PKBPXm+vCdwWh
`protect END_PROTECTED
