`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xN9mzHwOY1eLUx7BNjE5DM3rcl3QcvHY/ARBrpv5sKdTdAAWfzkeBh2WvkkoLzsx
f3yMhxyvpD35vd+AfQS6nq2zp4LmG4MP/Xm58aVI/bRbKMlSk0quFkNDCQruLJ/9
v0DkxdcRyZSZsWvnaTDnRJiYwXPZgzYTByGHO/8ueP8GU5WODr8S8CuUl72TUYVy
PpeifyhXRNXdKm0hIjSN9M5P/93xwqOwwxsNmC4kt4A68u2R+m5tXeg6MwMkP2Px
nPHcCtWZASKevW8Q7s1REG/PysZkoKQvpDKGoIeFoXnOzQc6wskqLD3oQIwjfWgE
Y8QFfM3NXeGP/jMqnwBX2ncP2R8rcCbDDmHjsCozXSH7ld2MUfIv9dQ2Alvwo2sq
+psdm+7CYEDgBiGBQpQt9wA9JqK1FYSjX7jm1KLGIcWzWFG9K+8XGlLdhOf6Szj0
7wRz3oAqa+fQ6tQGxHXe8gXTSKxRkD+yGk/sOE516wnmyZLsw3VSJts0nCEffOZC
DeDdCsg/4VAjed/PbRwBdNHbtxIq2Qg2JvdKW0qqawRBBEM2ixoBovG+AkgI3vxQ
qlJP0BLjKp5IhIyhKWTUb98swFoB6WQJeKWmPIbsdRbhxGJWb+uLpSLPc5sk7fDm
biEwRAWXnQnhpoi5Z38zUodK7T6q+QXZMrFDXJyzjF4L0NDxDu/HpOJxiszrBn1T
10SUH183FqutviLam0hKuzZzapLgDw3+s5o/5P1zuCp5hl2BIellib4maCsc5I1m
3LcxAFU4H0CP/AQ2gTR/zRSHG5T+A2YD9JUF/KFxirzcGGSaNjMghVzLQRumpZZS
GMBsMNd+lDHO3TC49l3WaoryXSU8TnJpvW/JlLYzfwfXtfFQIRFJcRW9yeCi52oe
wrr4W1NfXFxBVtkycCS+wpxW1u65TfMgp67FmjlJo5iagWj+fs1AUgGUOUjBeLNt
`protect END_PROTECTED
