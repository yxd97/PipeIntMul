`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K5w0PFmBOd4Ms+ZWT0pKzV9GLXFm33yrH/IZdYTZIG/OkWJIXuOPrCt2ybhDn8Kj
OsRIQUS9qEIw0epoRs3I8Lni7kFZCDi3eIvcmFUXiqRN8A2dJOnCUDllYQHaK/4X
cpMsjAW4tStWUPQB/o591kWeb7Cp/tWwRkSpekPLwL+TwqjZ7hFOPNoLqvfJXMe0
jp1co2VxNzC4qv2OyyQMs6Vi5axYb9b7KIe6hmVg6JS2tbyJ9y+PkO4cOgtGuGOP
+TBVJkfDhc8plbw/tvNS+hzj6E4gGIUNnX9j6ctM1NrbfG3CZ6haBvHwubsGKiEK
wjzcSm4EAyNnJ12IDAAsbXAQq/U79aiKOWZ2V2nl84P/F6EnxpyNOoYCe2+fnf7+
+Id+PxcLrzEqwV9gI180hGeVxQUN9HNx7oMnUjTQfnYakzMgV7bM9ZObtRcU8xj0
RwxOJSi1vdDHtiMZ8D6t1TUkT7wUQbQ5yOKbh5m6c9rtoEfiRblR8e2GMUe7qJxh
ud/6gAFjOuG9j6TBuVzRhG+gPI6MUp8zFxK/n8qi+T1VJJ4EkKR6SyOby+At+3o/
HUsMq+xAaUZ3CB1gI/ZXIJlCFmuxDB1XqHDZjK5sZPURhxaGbgnOe0QbCirCS1aX
zoAZX57EpRQv36C8UI+dAQ==
`protect END_PROTECTED
