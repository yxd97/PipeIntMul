`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ttc5xmOtnkGbBKVQ8uDDgpfh+1xlxWfYHSej4UW0tkvs6ouDUDk/JJHtedLDNyFP
8GU2A2Pn1ywBZ0+K44adJpY7qMYM8p6xMyFNeQEctKK5NX7QKGg7oWWXxPx15LSE
Wbze+zpCBDxxFmYRyFHq2N2vpl4gLssK3vVLE/H/C9YxKNXpJhbKKE47AlYn2iue
q9YgOzQC/APv/ZtLxtfv5/UgqkKhG7vUtRMbeWhSnvRH+QZB2MoFyU2fi3SbK47P
3RlVas6Jp0LljwS3nBhDgT3M/Sf/ShkTbIdqsLFRJz2kWwj5IwyC/StVAo56slK0
lHId9+Ky+MvUAN6IEKsmPtpQlL91sC4iNfRQD7nUr9W9rGeH7Ob8s3N7aF2sIpA+
OSOijYXrWFX+eJ5fG89QrKD2Ji60hU9N6PswdF5fTHU=
`protect END_PROTECTED
