`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oUvodOr0PcrpiXvmYzKjzHY1LiJvJGGteWV/JM383go4EkI84iOyFDgwQcJWTUUj
Z11qWrzs03vrCM2y+rgUJvxRy5Q1UIFtt7iK72bTIIWM3n5t01WPWJCUrKtbCxqR
aywPy4UFIfZU+K6RKHLxJEV+1vJJ2yTIejPwJWqEDf8VzDYGNK0Es6tiolbmPvSQ
W7arpLkP4ZZG+NIC5ouO7FMJRskAPpvCBLn4SBACM84E+OyDmZW0rJIN+eiRGvUd
C3fVmkMyVNMTTVETUidWUUX/hOzZ26BieTNllMll0hGuBlTXJCsy/vaCKAegypf+
asa0I9J09q9rO9DTMwEgGOxh2h5cDRJrLXtLBr5/rkY=
`protect END_PROTECTED
