`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QpKmRECPRxAi8r3xy87uaFEWg7gWV6OxHSZABziZFBeaoer7uGru5+P7IfuS8hJ6
KaMfaQDXV3uDFol9xv9b3T8GZYylU+/PpvruzIWCAASQ4F5CV9tOmdKdFldxKyH9
3WIOjHXzX75I1tEdNFy+J1ydORZ3DKcY4G0b2RCI0h6gGxOcQBEjU2PovNXkjBY4
Sn1/mfHO/saXS/hcImtkbq229hHGOf4aCshEXr1pGQF4qCaGhgos1hNdGtg2JL++
+7Kw2Wr/yO+Cb8sVMIru84cZ71g/7svCyFpYKIseERp4bV0PkMu4mCB+VzMe52UA
F/GCacfiP5CpluEvLDC0NRAiT/M9QAoa2R91C05/iEm5/KakplVqydy0y60mc7RP
LBA1a2MIcJvB1zqj9b+tDx6EvfWCEADWYrPmck1mu7HX5wEQq26zUrMadAPoPM6l
TpNqgxTJ8u12AN3qU7LPyQBe47OFY/jMOe0ZGULaerudJVgjdbU2JHPbYfkr71PO
CTqCUaF9o7WbzcNgG+sCLgOTQ6kCVnaDH0xE7xmw3TbcliN/QXeUIoypmcZtdUrI
`protect END_PROTECTED
