`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZHkOl4j/p4NX2JNllSYm7baevQbz21LWfWI0grP72ukem93je33YmmwgDh9Xik1g
+L9RLbYlTRS9l5ktiUdwRLVm4jZ1VxxTkNlooN6CvduI+RBaYXoSkgX1WmMfDSSZ
HWDqoWfY5+LTRVIr4LwL3xxVUwFpzQHCRVXwohdcl4LlKk2g5Zl7QXHtt4zh1lYH
GJmQbfNUxWi5PGmSbmP3avlOwOX3e4I/Kj/UvpsQp4TmL/X03HY+DNCJB9b68Bx3
JCbZx+k/ptaDiWxRhA/Xcl4Py+1OICgWuiLNZx1E7wuVwZdmekfWVXyG6WOFY3/6
p0rNi4EXp43AfHtFBX9vX40ozMRIcPQqyiCNpdKoHGbz6a3ET8Z7Iy+Mr494fJOp
9wk0uGm7Mv/rBk94cZgzUXXCfngohW+0vPRMX9hHOM9ObkuZwApjAQgyWc/PiXvS
IlyE3qM73B0xqyW5aURQ7DAA8OEe1ik5fIsgFcYhDJQi3u4SRo2VH0WLRdATTaj6
WWe/+vz6dFIfHgDSEAAisXu4Z9cYCwdxIrGwzVUV7rJU6IIhb8IqBr+DGUgbIDFT
bmN4Ks2aUTUWEizWZyztXtTVreRfxcDAtKq4WZJ1Xfv9BDXycjB7pcxdspYKFr3E
/YS7d+/aVoRO9wryqwdwYA5R3IOZb/6U/7tZroinLplX+LKasG686T6db4NxRXhJ
Kpb7MZp9CWp0cNPtyQbEcxNoSxzkrSMkCqhqWAaKIUNlarPBykFvd8pVO931FKLV
lpr+RbAxaXcsgeTACgQ5wgcOr/g7L/2a6VPVVc/V0x2pMtSAXYqTQTBWEGtsclx0
QCmpvzB5N3n0HpbTucfFHXq1tJnQaQIXncowiDUfyUnq84ptQ988NdG5Dd9268bd
AvokR3s5jnBgPpwygZqWJhLTdBBfVQyq6qvO1xmHwb9ROSVbv2+5Ckt5zi4TUh4h
hl5VleJZKzj1/cSBKhr2fm/1YGncf9qpHGKZl0ip9eF4rE9c68PyZcq5tVZW/M1B
KccFzZfyvR/4D/svfSMjkSWn8EMndVaCdbdVaJR/YF8v3COaLGAtRBHCodWTi3gY
Re/F1a90Pe4FgYk6T2ToeHCLH3Xl6M0AzpPvjX7i8p2rf73kLcjbYU/+PJBEUJ9q
q41s/0LzoRLBdkBUG9p1y53ojORxXDypUh+l48ghAuZBdFHYS9LfFRddT8pWBDR3
NjVYkaqqsBH81UggcRHxF4IAAqG/809to2iOBz7UUGfGxGQ4MobQGU+xW6OiApMH
vWV8lZHTcnBdmpfLD00RafzE2vxj/8/mIwPKTdHYbEtgPHVKS67rWK3vkLH2U1gU
/w6ZttSptZi97u4/3077GFHJM5EofbvuFq21WRdSlBZTC+djLKw+hpHU0xYQxeZL
0QiTOwgMO0DPdNGG2KV0UivWYqhxTSOs2wr4xTDVq3pGOA/Z0MjuN7JZHBAWVWGW
ckmaEsLRy6aT5IouXraBebY9EaUtZjJ/0NKaT1Y8OxI7OxMzszv0CJ6/k0BWBlte
T1laKzPyrmX0dpeWtjRDDiCzvFdMMFoB68onYv96NZCmyoJIzEirG208loxn8x/5
YQ0nhGwPaRphykYxDipYpNn5jLARF+jGXs5xpqQ3uKMwXMcYH7sWi2HEOWYxuDk+
FVS+Jot6vsAj0g3YHvR4Ymifoxwi3HbCkHcN675l0zciJKDgQ+SvjpA82s8J77rC
+Zw6bSMmqUsuxVvcsK3RAm0td7NvzsD1SPggh6SU4uJdKDAJK5/t4U0Jrx63V9uS
K4BtOfvPoT5E6Y0CtiSJ82/3nbCzXl5DbcgwqQR3UboJS4SboAHaEc06QHOZQKMp
kcUXFd9n5bjvoc19K/8jkEG0tj7xgvLX4+QLHbDJ252nNtHufGFKkX4WoB3x9xzC
le2hd8bxmcBYjJ0HgyjtL3u8EVPH65Pp4GtDK1XUTDkWF5E03TUwvI9t6mCX+yUc
As6PW8xmkujyhzgPudRu8UtqXjoUwKsx6jCI7/+9UY3ZpJaHEO6njsFj9czttkN6
5QYBFJqlYQmM3VnsfBBvVqHcoCVrW+Hs2ZPMoQoM+9R8XpFbkaD3XCqRClnUJxG4
0ZZX81iQJnii4hB+CIraZwJYs3WKafyN96Fa8pgl7arPXfJRK0CzQT4vTSioOGoa
eJNx+TeEgwXnNGjioeti98laxVhAPA2FG3244UHpsamvjerQpZ3x0A5RKmcQCsd+
+MRMXiiISjT3MIcmNQixsnEmORz9tWngYd5k7cm8RvUuBceqa9y9q56WNAl5cR6S
YRfIHOgtrctrDmX9Toye/uZ8Ee2QJ6N57IUGckX5Lrw9b6aDhakKNodWoHFP0UX0
ppT+N45YV5QAKpNofQMxtqqdJmfB9tnuIbhlA3rXHAFnFLKi1n98VBn5TAJQXC8S
1LM3kTq/fHR9notFSwRuG/URBrI4TwsrecVHRJnT5oUfSgOYTAbxYdGch1bPMb6U
yZAmNR5bjNOgzmX0RTsml0P+AK726Q5XTi7S+LDPRypudeKpIIR92PKLiJl/QPuN
RqXb5mLIMx0UpIXrb+Gv3dbR1VbiaTxU1C9cC9RJuUsZzCknVLg6uKyHZj8pcfJK
aZEmwKipI5xscVmmw4Dgh3z0FeDsH8+7e0SnCiPE+SJD6eWbz90Ik96t3/pgtcqS
K3dnC99DB16FNd10WhlyLJzvWx1nFshl1VwTHDbtsGLhNx9NTvivZYKupTYzSdv1
3QEggwWspAYvJHbLhT4GPaFoPLUzo/mOC20mBL781OnK/Nu4SFYsKtjjrpOJMSsG
lkCcstbChBOveq1SOVFJkUqa7t6Nl0YL1Vy8V1P0MIDiHPHdL5qq7dOOwFpEH8YR
1cyoWHy9CVICYR4syf8wEuNjlZ4FtVu+fwVpoho1EgBbVCpAXcoqsxy/cVdByNuy
020Ge82Eyo/IiLqvJ3CD1g21RSBVzTV4H8l07Ih2E53XzhfZ6/x9Ogv9VqgzR79F
ICYT6zp50sn2s7UwQcEG+kZ38URNpemqGoIRS5LUjo50Dcdl8zOFbQreedFEacYs
xDEryVcYg2KZ8lofFFx4YJLMVAOU0NyUvuzboCZL07c=
`protect END_PROTECTED
