`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hENcDyELQfhNtLnHa5uMCeCs4RtOmqpSFKqCAlQb4c7UbDH7kgmpjrtmeuZuy/WX
cKPeV4BixymmJCscyAxy22lS5IxoFMigHxRefXOJDr8n1HMrG9PNXWpNis3AUoUk
WDM+GzilPKnPSFG+Sz/zZVzlzSKzdXZv2fPkiL6z+9D3hkqihWxOXXizJEvkPgp6
jCKHi7sXn9iggGLZPyRXJD9FcXbIMAIbPlcRjq1Bx9oHHL38pa36bwweWvxwgQSO
V8QlfHHwhXopcRu3eQLpzJwUhxAsdUKposIbQz1jW57z4/TZPEr2Q7aBFdyFdaMI
m81B7HYpDoniD5Pc4KqBCCTu0m35IIAfPAYcrq4OcjE=
`protect END_PROTECTED
