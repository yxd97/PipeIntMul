`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
arvoOFhMoHqI9A1xKMT4EekC3ZsE4doF//8+Gi/cCwSrkfTxS4DvwW+Gx4Ge+Yrn
RF30as5AqY+U4cZ3t4DWNcXIweXKZMs4/WmEmIHp1p8OEvyHCXFI80GhRY2WZRNI
OfD6fEQrNUJkEixyRUSPbJCuc1Cq9FSK5DQVKb2CuudW0VfBPLvjxOTnKlfZMMbf
xluQ9aT2Qz/jw6sEYnQSKfhzNihnyb/I5fAUVLnTTaIjoozD7kJJPwvagZOmAnGe
oYrtL5lV/d3MLf7b4C/OtFr/NQrQoXRHmSug9yqfKy/ib+1Xy+PwOwa5IUOnOpsa
`protect END_PROTECTED
