`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q6WkBWXBQvWSb1+T6CLBjXVaWSE3T0JMTwZz0rBkFuIJvT3VSWqxr3vjAG1OsHGY
RNTJI1a7GeouidML8wxGx4wZR8E1MYBxz3XiK9iqIW0HsgwGew0BasUh3k9b5o1b
7vQjcefa0xg+Pnh1mG90K1xUn8z8+IJHQO9p+NAZBfm+/ALsO1tGtgzGzPEiPZIN
OKV5wiv578Qv8Z0Xmw9DoRVVfe2N8eCT3ABCl2dQ53AAYTzpBF9wwVs5QMV+e8r6
eRLSHRUsrsQLWafGj4ShiF36NDqP7SRzrUwfOp3SItV2V7PyxBEyVUKi49xdbT40
7pUoXZ8+oifvpzCaUV0HIcRlbSXQMuu0MkWyGazu8HcFERrZ5DKoxLaDO67ftooI
yTWx3q9/fSG+Z8CyTZh/BMC89bAH2g3bo03w5DA7gs4=
`protect END_PROTECTED
