`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
huRedmKnKvLZD/i9o3Mbx+JCSRvumC1YyLZyp1hEMl98lYHefXHLRXwVQHw6fLfJ
ppN5B2z1oM0d9ax91R8G/Kb1fbDWlefC9MuGKVTfDi+X/JHKqRIA5/6ERQ9rvIkY
BSdmIhrWYhTHvyymqA/FTqEcJI5Dw3A2IsNKg8wBrmZfYF53fljrM9LBVqN6TxlY
ate66skMxMLicI/CInla+ROvUs60yW9rRtqJNynlnWPYbdqUZNvG2lnBrESSi7Tb
bURNRqacFtTNaIxtoTgQjmDPkbNw3Ei78UjEwcLWeGo0OAYeJfv2zYZCKKT8ydqh
TNiPZ7RMD5eoRWZ3JlA6GZC8NwKUrMWM9kfbkNTwtW5J6Uv6L3Z+D8iHqVdkRKST
R7/TTTaFb2+wjUYCTmDgC/rCegRSghiuXtWQwfK3d6KaGcp7ETC+JlrjwrCQnXVF
dK5qTCdI5E5mZm5nq00fr1qYDSpEtTLXHq9/Q6hXbuCEn2Brs+2XvZeui50cr6oh
VY0gMBUg9VUsfVHO4yA6pEMM4jOXFqJiGVWGoS9bUk3PADsfhstImKbQVGLwESgC
ByJU5Vbda8liexNxpT+q+wPeYYb3JrzECqQxUaQRtRE=
`protect END_PROTECTED
