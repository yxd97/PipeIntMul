`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
r9nYlxAkP82klXWzQ9LGS2RJ5gPvbZXRx2Z5z2ryshh4gj2yTFDKcza1j6/ND9gB
544XwfpnXdc5heYPmIJ71LdlM0UUSozlHsxeY9ecFJCslx6I5KHToq3YCD+/g0/J
TGc88J30xJPbdLaaOHLB+i+eTL2bsCpYIkhXP+sctkfttDfH0COfbbbKSwACsopB
s4xTrKYrGWMwqPpDu4gIFtXUPCLSb1QQKkpFVx1jkfgXE7qL/QkqwtqrBh7UnfSz
BP8mcOF+Xp/lW1zEKImXXA==
`protect END_PROTECTED
