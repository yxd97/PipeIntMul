`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FV0odlQ9rMoAkseruaNN4flkJTve85izNheXil/sXiN30kJlxIuGut9OJe6uc0RE
KyDwOBXGDu+MA+aIS4RWSb2NzpCVzNi31PEy1I/uBrVi8dZ756wco2XsVLSV9LSI
LnbSOsAbUYeyaVLEG1MF8IsG5Vk65C5Vh/7NcVHFfw6nPokhoit0/9D+hmbtDX5f
pApOU/l7x6OX17KxLjNP3MysRy6CHXRVrOyfPUsQD3hKruSyIisyWo1xN8a4TslX
sqXFdOJQzFycGx9iDkhiynDNJNGe0RCJmqh+xITj7Jg+HBL1AW1wRIh/FaKiOC1K
F6GSOjTbFw566UA4PBz/ezZ5LMVz1oyrHxc828S0jFiAScRsYjR65U6ayWsCHE+s
Iw5BLWm5Xf50Xv6ot3N2JppB0jZcbWs5sFZGaSV/Gbo=
`protect END_PROTECTED
