`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
V56/6HyIIlXVtnly3oI99qU8ui2jnP2E7QSRPxst4VE6+RtduV/IYOILQyM8cjif
gkbCxiI68k3ZvXpVrvxy730STOGe6hs5tstPl+RQhSy2x8TYFSNTwptQDfmnDlpV
bzIQ0sUwfhGknmpSpnBcunQCpPl8wLjeit+8cxwCge0nNYnYoxMGhNrB0MUgvoMx
mwfIA9uBl4XTMv99lU0ShmmzKu8JoQdTP3vUfIfwTQ9v5DsD15mBF7a2wfgpRpnz
ch1aEE3SP7FwiPtfOsZwr+EDqi3mUV+IknTFpv8dNBQvFsliCAtHFVid+B2vEz1+
epxrcJHNU+1Sm703sm5gJg==
`protect END_PROTECTED
