`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
coxaRu5qCsngL6E75uchMPOUkpmWo0EJN3yBARXJGdL5eQ5DCb6Chk/6w2CYy8/I
cUd4etNCOTLZ/UfyYjN77ZHL/K/LQst5eYEBIIVn2EKIuCDfV9kERM2Z4i+x64QE
2D/MxTpX7UF+uWK5hVZNJNFbuJAusZqQiGEdA0zc0m3oiyAgisSo+dbTogbRoB2M
COlEuD9S7DCuwn/wUsUrv51f/pE1ltw7IFpcuROosCslTwga1hJjIIX1EB6nHNki
jrakn6vn/bEzcM8q2laxd20GYypwBLLbqoxqO3BbAxHSKy3jBceIqorCAlzuJcQN
DsvptB7bKfKd+wnLkreRPdsWvcsookaLIG2ErXf46Qbln2gZaKZLnv4Yeusp5iyu
t++cmt4/GJQax4kllanJEFepJfT4S5a5MzxfafrxkoQ=
`protect END_PROTECTED
