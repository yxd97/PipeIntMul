`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ie+Ytrckjr0qW1sIYuP5RBwTGvQWbfCstKL3rMpyRm7TiEJKjTxvz7NyWkM8mHbU
e1TuBs/r4aDhQ6KoPH0Erv7Uiy0THzKkpYImk/LUlFU/UU7bLIDJMxUVZUdzEbki
nRsk6pz0naloyfBztryZahFmM1BiSIyuYPK1CkqyPQq4rAJbP7AK0bHIy1AnnJWq
v36g1me19CY58QIzXM/Iat9bKHBT1EmQSH6UEZKT7kFhnIt6bN0DlMYdot1ENvA1
3X9wb+rlt8wVDuiE4mD+NeATT9jx4qrLV5R42WrCfaDjyKKvlG7Mz5a6nZ12RWRz
3zVL0/t0QkWT+pzT1FTtI5dtHXkj3h3Bmydm63hS30V/hLdQMSzHgrp4zLKUXcLC
+qCqoYfNe3xFfuSV4UfDf2FFKlsQyX42h+jAHe5ixOyFnDCvADihEseAQluVK4v0
2U6SPBIIMsP0ocwgCbpYbD+zwPUzi0WnEfgrWtlU50NzD6X6Dzj/e+LlGIBOmjK4
eN9EYsbP4/Y+Ccm/1OmkDESQse4OCKPmPXemBRVYwiplaINbfAZjeXD9LOXxa/7q
cz8hDyOXiOlUvCGVFiASpgJcyepOvfXE9uX5130vbmqL86O/8HPTq0Xd24jeZGp1
1f1ZTEyaQbqGw4Ewehf1u3QKjYtWsEQvuZMflD+aUHf/fX0y/Fxq17BMEjoKFSjJ
8TeNrfaE8e18od1VP3iZKnO/vZFhuEAaCV2fbSl14wPMM9guwgtm2a7LZewJ/5oT
o2nTOSDDj/okIYxzN6Q87/BkgJC0mgWLUY9PjJdGxqEDdfG1TTllR5aEYBv8XIFc
pOpx8kp6piaZ4Yts+32GAGE2H+ljcDDvcM1hPUb28x57YXZAY+bImtq723585tIx
5iBIXUmExV4xVGA2vbjcRzJiOlImbrixuAYoNUusCwC8NSA41fE9c0sjgUAsKFMC
5eQmZNZtt5178KzU3qSm7WoDq70MWpkO28qeDsUNEqgue0K6YDmMOPR1JL3nD9Go
Uxv+eh2GLUsZC3wHphk6J2ZiswK1PJcm7osV3BMfbaKivTNHgr+ZyxOGvUNU93Mp
4T/HltEBfJtF/72ebPrlV8mRkhUXBqt/PVwqjk7cAjiKrf2GlJ+5H3Th16QyT0a0
B3LT8Mf5U101tYoRK/OG8Ez5mGjLiGRJqJL+5f/5TYL/PhpZRDKU58Xj51BY5g9X
Uw8RhyS0ig8MHGbBeOjyNtMK/6pfvwmOJowER+7YAwz+4OmVAwFgcm4rn++i69ct
o/wZMKFmykaUiZ0y/8hztZUEp+tAHp8wPtRy3cTR1FjZIgmkiF5Grehsl2W7r16j
Rbo6Cgt9UcjXavx37HakLeFfh+wKTfGGz5yBYMecJuDu6i53ofhI0qfZAOeHEm+k
Ha1GzZiM+M5Q03MzOtMWOX2Q9l6jnE+4APXVWeZ47rMQHb7obgzD8l3wWfD9GIbJ
GZDbJH7BjOw4Z8j2VobLvAVSi7DOwVqXvcuomx9W48y+jWt1e41qvwfyriFyZE4F
H5McCXXmmYKKs2YSqiO/WNzrAV+mXMiWd75fAyefOiY20nA+PP2pcU0VbvX/le2l
4FvWULAMwbsMGvPqmlCcsRU+jDDbrIxWae0KBaRNuLlfxaA4++CoOcPlEjIxrVnC
5AXeE/dHJ0+omAUX3l9CUdBTVXWJseGCyXgPsOJpP5MSzBGraSvtJ4X46VZXHURH
kFYFmC5i1G36y4Nmt/yaD6h6jSEQnklO8Gavr9QeRz87xdiispYToQ8W2J0wTBWG
lH5ksTjz0F5ZcKDouhP/F11/lqo9X68Mxo/wPKnRwh2oGdgLCHFb9oiZdaHOpWhS
q0RkOAxEGlUnh6zvBSIa0Lug7iAUsv0sAwkM+OS1/Aq72zehVEAmJbYZlKlth9Fi
gLhKDvje5HDHyeb8YA03wDQRu6fY/f0c8DYR0+90NgWzCJqNMm97qKo095Zb6rDA
VZCkYH72GJk66X+5bN0WDNCFVYfdSTq/BIquaAGrEcTaARTXTE5ukbR+FhOrJuUv
4DDSVr13zKhchgp1lgCARqEpujw13EpX9uFsi0weZDmxIDQ4K6ymSTOC0vvBNmRq
MkBdMrhWMBmvP+Dxk3CbWZi5Xw6JdqbkbDsv2YwWAQ98i8Ifb2cxnXpHkDbunRvt
LgFeAR53UPnz9hbPBEBNnfDuARE4+0+Lt/pkPZFrfEfRYyO+r7+jWQLXH/e0W16C
HfXWp/XmokhfvfeZc3gD/syjKSrDgbTYAkBo/8jH4e/SW5UwiK7A0QRH1MoD9anT
kVSvFSYgVPAuNlrubgtvXW6pPklVg6k0g1vQ9UA2jEwi4XzGCfi8wOyq3bTKHJxO
ju9Q818MCDhFb1Q2myVbuSfrqM0mqopubRittXDfoDVjvcA2k+3nWyjyq92ZgpOA
2dVTKBGhsr24dXAD9tZ7J17iUl1it5+w5o6Cg9YyTJdylVK/RLDN44aH0eLsMANZ
I+zY5RbgUdcdG20WDVVORwTNkEis4fdBSLyG7P1Si1e8hat5T271LfC3EOaCGOJo
MOUIgBh96OqKx+HeSg3tklJLPKYGR+zWJNmRyvk+is/E9CDhad4N2LbCsPKy2mEN
mFhK/V01cA2NUlzG4SVe5Hc8g0TzeevfIdqGTXhTpsTD3xC0c/x6wVz8zmq+Pg41
cmY9Vl7SJ/QoUfs8uPiOzk5TQzg3Mgpve9/tvRSwJ2ryDIYxnPQhxvDib3iO+uJM
W6gWtbMB2/hbOwAnS8YQ/OPFg/bgWAi/Ku6RLVH6QZhuiuj5kukZtkkb2Bm7IXA6
BWqC6dZhkbL2bkvWgPDOn9Mo8T4OERAJ8bvTLSWJLN/Hpr5nA3DY7dgsOmpSqdey
dbPeuyILJwhO7zrWltZe7ApY0ylXcK7wOatSZFfSHWlaLp1C/IlJl15S/147gmoD
T+fxoYqz6j7G3h4HdJ+WnPmKUmfmOZ78VJWItlS9UMT7MJT+IeIXb7YZQM9x+Rl3
kq3/+30wzS36wa1pjd5pIG+K4OHYh6X/APjiRD4RhhM=
`protect END_PROTECTED
