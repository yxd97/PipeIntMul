`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nHqvFCwz/pXX2rqmYSzDM6fl4F68hpXaO2OyXWNyrqpW59lo2zxsKuS9DlZ6ufic
J5CeLwqKUrtdWuPGuoYovziUnqOv9fQLGfecJQD3Ca8iaIJjDWkX6OIZ3UJcMoTd
mTli3Amvz2j88bM1cGPT0Toap3i/9czKmaGeppzaOhaiE1zaK6nG8/SiS3WsmKaV
anQXHqgWPyHswT0kX+RF6RkfyzzzSpQ+eHpLC5gTSk6t8SOBbUginyCzX05L3jn6
XhLI8UJumDJOaDCpB3X5uS5sVslgf8T7QfHhLLzon1woQxhkcyT3WtIu6wmtOZHe
QSPf0AA0cxGEXDLeSoyqXSdvqAEQqpLWEMRcCP4HiT6IHTALGlmTqLW3lSRIe7hW
JSqrokOCO44JqeXYCQUDJEF635++9Lf9W8OjPpJThWl4qFlt09IB01dL9FCSBgr3
/cKYTH/N2Mb771nG2DSOSDICrY2xKTedpZ/65kzaJnDZUHeRY/+urRNks1VTVKIp
6zTxIAsrMzVOFnT9w8bWVCju+4emmhEI+R63ZtYnvDNHKrxpqDKb7cFviL8kTowM
cg31M8q+Cq/UcUzydNtwA/YxRFSQ++9BVqlp9pWKpghhDB3CVes3S7/0LUswZvBw
+Jqb5H1WaE/qsV4BRCfX+o8QYAf6t/04rhevSHuzr+SOQd5Qnjc01yWUfAe/YPNq
AjXQJ1tPxXHhsSe5QxhEaGngHeU7+5j3Mwlzhp8yKRCIQcqXoOdqsC5q4EGU8Yvn
cLe57Sra8vlXgXp97ymcKj8vdFXJuj7RpZZOQF5EvjSXm2yjuGVxg975EADZkHus
WFzrxjyqU4e553z1PLf41JBD0lXLFZAfhTpwbBTTRmFamm1J37AKdVgkITasCBBn
Le83ycAfyb9yf2+iQBui6ZrXNK2lcn99fZGrH/pPtQvjitG1dYQbol92rBD+DoRt
`protect END_PROTECTED
