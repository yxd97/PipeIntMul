`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c9B5dLK21vBdxKeVQKMI/y737QKB9LIFwOI2yqYrcFG4OzQnscCObTZzbBLABf9U
O4EsKHCSbUeQ+bUJ8hBXpXCx3136ufFiiK8SULrp9iM75SDRmYzJQCPrfKhm/R9E
5MOyTRkA+Hjx++lYK9XqfPJbksIP3MjhDznJYRv0cgoK8Gg+xmHNkbue/vZWzfMD
DWRHJtx0Z3MGTUixJ1gtnp7Zpvx3VHm4gucddVQ5zAvCkfFM62nvigtAljUvQw2D
zzZw4TgeUFA1e2jRMRSBcupvhPDHJ49ul6ITpXRZ7fDR6I9hKwXaYy6WOf0y187W
3kxy+E8CXNdJRef10bU2TfZM1l8auu5MBRY/d3T66BjLWnyyi7JDV2lvSjBpBOq7
/8Jqkel8TT8vFKwrCv32Osu8oLcvUGPOYQC9nnWSa2opYGBwYsq7wqg5fVnOBPtt
`protect END_PROTECTED
