`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s30KaFgtFPrEaCog4jg59bSQWs5zSOnKnn4vWp9ctxKdBr98IL3zGL0QU4fJAaGD
pFb1xVCU/0XxY4ItNNnyh7US5k4O2TiSllOrJjJyH0ER0kV0N9IP2Pwh5fvfz9zD
Hg+64mrSux2fYtxYrh/qJR4gABB3+c0gh70BfRm3XMfIx+Jbjm2ioPf+srK3fZPA
/zBiKchpD7My+OxxM3H8i2XbtG5PdYqnMWsvKBseP14gzMEPDva8IoGtH4aJWk/8
3dCBy71HaaQBtBxwgudSh02XnmdbREdQyZ8b2SOqtR21N22so9ur6LOowSvKP6D6
Eh8hgERlqEHMeiaRBaWepUSMBYaC6ErdPzbQIv7THMsD4Fd9+bsE9NQpSvVyA7pj
9cp+fjTPm79OqktrfxLoJUnJ+wdDWglSa8iHhmS6pxpYeCJzf21KZ3yjyz73mpWh
`protect END_PROTECTED
