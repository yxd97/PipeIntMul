`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qf8i1KRJDi2hKEZbQFJlw9RU6iQZ5iMlAuRBNggPGGAB3GhJRphPVl4TnYwosqZR
K5uEX45UGCAQLjpKsviaUIX2+Up0wIew1Nm6guNGzqzhW42Ab36E1t8Rg2UzZwSI
XG9TAskJ+o8YelHHhkz+O3S1+R+3ZL7Fp7m9pB3bFNzES59R9cuuF7sbyv3uEv69
CWitwQ4p/PLbRBRlYMoOvmxCuVhScEQIzoGA85/uh5hIxj0v/TiM2fhtdKL8RBgU
il27xJaO116rLB0cRdFnivWGL0t1q2PkLHD7GOLkYwZBVxOKWhw6/3/wXGaP4cw9
uXUVK6yLSqCo8qTGhPsCRmsGdiiD64/c4g1BpGnk53jnEDr4i5W79YziywW8TUKl
59gorRRLDvCHRbcIVfvByZP7gU3yMoOvhfAI2PHFlykOQkm0QkvNqOA1mtm6+E5h
we1H+hn+dPdXC4OEGbl+7yNaz1WnS+Ah93gXIxE7s0g/zQaINAHsZoKhEbuw2BAQ
SeQhxij6/chKgDju0N9WWmSNx6P1YEPVDAKFvR6mgeKGzvJM72VYROnCr0VsUD6z
jnoSquJE58S0/pHSRXn6rZ13BjkOeNx1515ke2KdfM4/gEQrtesXoldQisDLNGuv
YxuyvJztayLrF+iMiuG1KLMoBMP9/QE52kTq/BHJFLHUxtFY2VbCM2x3DqHjSQdQ
rftkwhhOieGI/lKHBEIEv+CmKg+lIXk6miYyXPxgfD6seBIFATjSZWWXL2dtmSpf
RE06md6xQXgzPZaKdgecFTe6tMmmFtqAmUI51DOYsO+CHQFm63jjcsEkaViKcFbF
3SLFVqTuqtS6/gDb5+Itql4EuKpUrqNzenbnF1a6FxCNqhruh8HrlJUzLsrJFLGp
ihfjpB+GgxkktKCuJbPAHxGajOG9XaA3lHzZVgfPOjZlRsVl2RWYbebeOPwZ9spl
zkZnDHyDsRtCT/nJQ6dS9J51zKW4GMMzBm68lzer8CohdMwKR77QNoTKKu8qNTzT
iR9ACKXndtVPmcLChqt6GxQ7MHVckcjf14Hj7j62dWlyGIrcZfhxGOgjhczFogwX
vaS3YXJqvmDhhZSG8BzBS51dEgc6onhaZojaca46u0F4VOyKcIsVsAGkNI8PJgs2
Zs4AjPsfeO5CvBToXVgiazxAZnCnZsXawY2O+opwSlkhsNtLZUg1RSHquoMxusci
ltn08D0NRQw9kXGqtzt9L4M09bGKfi8GwzKfpwYNprO/5VMWRBh/AH5POsXNbSTn
aYnsCHNCsleukasXGqL12jKavfQnqrEMQoFShz7SpceTl8GJ22frDW7sgEb+327R
9SxxzPGwOYlcd3ZBAiEny6aiWgkPHioyyl4BHBLbYpsLDfMRn0uLGyAJmKgme2Kw
1Gh9xrzuqkQ6E7vgc9gXxmsnFjQeDECnBC5ahtq9vWFE/aUq6LeaJvOBJWcVaOGW
gR9Z+zwqR5bxQHHwbQWWS0kyUtG8aX/9zt0mnmynIENA5m5sqpe2Ux8wG6FTJgc6
SwY6YhFcUGbYVF3HtsuZYvOl50MKwIA5+eevoM5ceT73BRmY5G8hM+IlGHAZvoVc
oNIIDRT/43B1oAFsbqg1AQgpXz4T8juQrAFn8zZD+4jYYK4paOeJXqiefa/e/hg+
K9tjpEa5MUpyvSXJi/w1B1Vjl3bXSU4wdIy44EXc0JiG+YX2e6qIs9rIXM021R3d
JlYw2nYKloLOowZyQ2GX2+edzxRvcLH75peQzc3he2JGLREhKGqpKxxl6dXYr2rt
vsxRq4tyVX8e5b/QfG4SvhSGFA+AZv6/tOiA3XqPeDfHeYz495huIggGmmh0dhxq
p34bMCSj4VW/vyJuiyhsWEUn/K6bHl5YIQBiWQm+DZHLwNO9b2A4yujHTbgr4Grq
acfxuevNVhbRDlSLEhPYjCtuG2787xILePFNbfe4rzqW0onS8p6p/L6ficUe+paq
lxgxMy3vQD/hFxVQkJLQLfrEUW+JFZXK9owHfDNKuABg9+Cf3a9jX5s18UadIeT4
cOwSn6jFbuRSHv3WvpWuKqb8UCBg5LtGJv8v6oVkRC5vHBBkq71FHFZh16jXWKln
0hIdpQJKTUkv+Xm+VpcqFaFI0tNRWvc+trD6lZGGHotFnfqjHF1EOfEwtGlYF1Ev
q+V/upqM5TjpeKBPaGJpA0xxTxSAZzRjIvr35lXLO5mmQPaW8R7mnrFY6ZpHzSGe
6HIyV4Cd10RFy9rymJYPc4p3cKMKodHmDeB0ZGidizlvtKituGhuIVxYAffWGTUC
1vLLhbDyj3d9RLlw7elXPh0aR7o5Qs2ohdqKcxOKUMug9V8wa0T21sK9+wzaYyy8
3F4YICZLhCTn8M7bcJQ5oObrlAzCndXErVCtJYsGSKbebyYb9TK26FufNFyKmk7P
BHYZ38O+d9KwgHa9mjTFjCzL2PMtBxlTRfcz6BGOs/z+AgEsZUZFESO+YCBHElex
FtPJGCaeF48Lpqbe11LZnQaTiP67M8EnLotDhVe6NAE/hp5Fd0fsJUWit1GFv6tw
SnkSN5/pNXNMARdfy9bjBUsDA5jAc/AYg7SGRR2wzAGI5UpTzz45FjWl83O6v0uX
sSO2yxRNEJPeIDcJa7qt6cIkaviHj2VeVPizFvXL9de1mZIwU859cH+zwbMoa3Vr
/e+XvUWhCGTEoLs46RaGvMCJCwyzGwJ7h+MJYpv8/hEAlKP1QkAdJvrfP54bdfzw
rwnxRiCLwlf3V2ajN+hLuRTM+4aY3CpHaS+l94PYoE+62wJ0pZaiOwPNX+nknmMc
aDoGQ6E4sWtK8WY3Tex5b0zbFRqL5zY5cSLd5nzeJgsl9Q89IMfVe/d0npwTfqbe
jBUhp/v69w0SuhOOTUrCJwRhvz5MGkdUKrcDP9g2BAQNOlV4AYiX7W2LQnB59tVB
puWdJhw4N/I7pnpumJIefYpe0ajYryEMpFkcAT/9DldQHsbfjBANlIuby1I5+qJL
/C5nRLGbWrarjhaze2gZ5m6a53/kcys/KbTr9D2nYFGdlTSDXqXSCft4439hfNU3
C93bArJAA4wXpEKwdOy+Xi3IFFKQfsELjqVo4v74XbHVexD5j5fJyKX9bpDQjAYe
wHuglwg8sxkxgwoBz/vv/o5cP779mK/asenUvFm2rhIcLgpRQGfsN6fzOesRB+nW
XWmjcb0Lzl07iSG7DVEHq1Mnb20TWoPXcbpmdtX29HoqlUEETbn67g6q3H/V5XcI
c0NbqwH5jPMYLXVWKyGl1rtCdqzc3Skfe5vc90Avf6YCP0kN8hxstch9aSyyFhx3
RV3t6X43EuSf/c3xxjTgwe+agZe4QfiXlIoLbWdtw36dkz8GSeBor9BALR39pP2L
eoU2ghsmHpMhM7JIVDy0XuQ2is1Mr4Omgj5dHEPqN7/HJldNT80adQLYyVHTOMHL
W1ARS4dfIxoVVIHqLYq1wK7I5hPwBKCWSnK8DMaY2OKljtlHamAHRemUsE+kKpvO
CD52Bgd5aJTmNzCK5yxtFh8qSBsZNVbjZErcxpLGuXMrP5c/+HRbvieyR6DDtHnV
LsrA2sAPiH6AQAArBitA4E0byDl6GPBDdXwgopL6u4zE+BKgpxvPuqGuaqASUjNb
5A4pfIARJljQWCGOA8s6eYHDVlz0vEMrndrZhfKL8slfol044GD33+v8PRMzTj8X
TpgOZTj8uLH7Ce909Gx04DlWylECZwDxG0SESTEDQfwQKFhAmkjh2lqJnzJwAeSx
mOh3EAycPHsNBpFTUVUNtu/dMDXX3QRlIvqqE60VSTM40YjA7tLEgU7owSNWnGn8
WtdjF9s9hAZm66fRLZVgEYTMDMC3VCXxhObG5cwS+O34dCX3ZRZYzvNV9E/agUPt
Lq1jYb6T7fG4QLmjyXijH8mM7F4YRgyemiqPwRH1usQEPwp3cnBg9S6f+DgMuRCA
d20Fz3qWSbxfrrPvC7vgWeWg3n62VUOLJc13NK9yiWUfrvxgkOBSr5xldf4rGL5k
9vNrRgVtvPm8qWkEaIjUeJQk8QmUgaGYyUr9xYtz09UG8DmDnS9pVLefz2QvkL7h
jfCLai/YWxdHz1bYpNAmMFAIIopeFXVJBVNi1O4w6bmHw4kte38sKDRaU2Of1y4F
T84Sdcf4PZzOgEmy6M7rIZ0e+Wjz9eaIJ28zjqk1v8ht+7GNSIzLet9+yKeybJsW
jeYtdAOaz+GNuxeHb8UGJO13rZWEaTmRuJMkwSlyVNzi51h07cdvV1Z9exfuDm/X
Q5XlX3GkTUARFO3IjLX26IhWbsYzoTYzAFTL0F3OS4bAJuUUCqJ9bXbetNOSxY1L
Y5I+K7FrAUrAd0Uffqq7ovjRCN/H0UchtQ0GmtqTuUMv50MvpU0PyRrUUWWuQ+3u
ri9lOcZ9OqcuZmEnlT8tL57qaxRm5a9gfby5tLzj+Gp9sTp8R3VzhlCKb++M0RpQ
rTjsLwbbBryBO7sWHwT8/7TD7FoIr/1i5PyWaio/yQ7dlZELufeQOtuUQNv8FJEr
5dd6X2yXsG50yLF6oZ6WtMyY7NLtxGt8XxScUvkLUi5Qaov8FUs18RnzzXsOS47Z
mYgPKXNAN+oCvSR/JgALe0ANz1DutxWuTsPNh8iX2oj5vk+bYz05By//0di83LDo
+UlhZNtQXAaL+ytngn7hqkxTMmB2TCtP3QgaA62zyE0IHAjYjxOE12sBfGxOaxaf
PcMIwuxBp/a6Np68nqxQuwWrv5K9+09l/jJWbGabCeLQkwke/Eb3UHCy7nTn7TcF
IFO3vKQZtWoIY3THFmgM0mqD2wb50ek//MtQbjcYkcvqjuVEvFJbYsewN9RqVZLr
cNYnrlmHDBdZTfkbp+bVWghZ3ghzl99gaZI/2yVTW5EoAS+T9wrbBJmyRE0AeRq1
mDix1tZbw/nrPxWeu8P9tJYLQFZtEcAqU5GFIdFkqU8WQsOOlkLt17Tq8zdoRhrP
MPizlfLh7emPHCuqBWpC8isHcEathe8AyKb1B5ogyDVSXXBFpaKlzoGluhTBNEq9
aXe77tW2XSxOORyOdhODgEk7nkCvaa3EhZ7rQAOW5Z9IdY7vD0/gpOHst6lVX8Wh
+Dnms56gPFxUBJFwm4qGiCsc6pRMYijCzCg/OUvb6bU0wEeki3b8H1s5qdFnVtRp
HUoNLcKYYsNi3TKpBusLJS97IVmGQV3ttwEaJ6MZ0+q9v3aItnUPas/9bQWafIjl
2N/4vh2I023Nh7htB3XkvR2poyKBI6N6bBF7UV7K1j5ew5bUcKZK0oXGaoz2NeMf
nHLciUaEGQGmdwbZ3qMP+34K7l4r9H1XwXvhslm3f18jGAvM/54eoo2dVedSUUo8
H4CNtG3cPWm0e3EsFXGmdeg+5HfnSDreVSy9t9aWIKN7W5NhPoVHK0v4iB8lxztN
jCL/IJXFukVdz803IH+eJyGz/3wHnShuwPxeothOYNFtuYXsRsCFgXFz7u4xgADr
zlzvMs4OFzY8CHQkp1uVbR3ImhjkC8P9ZyWhbEUmiBcxbiUYI2fV1vfmT7nJIoGQ
Ro31U+2TLsdzMvF+AMLmGdrZ++BW/BKJBm25yx33GlnpiVzOM38HqAlwPQJwwMK4
FldGBMDYIXo7G1zIGH6xasM6CTWcbcSSnqwOyvcZWf6TO+Rp1vY7IQhBKAmbuUBI
zkaTrLfQnKISE5E0Mw9VlelILDoDbIO7xOvT1DsI05UK08diZ8r21CH/1gAIphoM
XsEEos2h+NfmVJTVvuxySXicLJt1XUwVTEeLE8oPWYUAWXoxg6XVzCO2QOqkZ7C/
ZgjjGeyPfj16qPuMfoiu7X2qCKl/0DTsAqNbA8yRPZ49UzKa/1XiZTZPq/5wz09v
E+XWZBTp6cOdZzjvlosoKKchqkXHXfAC33CHCk0R+44P5I4uX3pHGi9m1gDpR0X5
Z4t/DHMg0BavJCMBWpyRk8wd7NRYpFndwQpNQ36vyDCK5b4GRdHYaIN3uGTN4fjH
/Bua4WJPxH6iysyv8K2b24hhZDwA121QkuXDvFSF5mhmtDWmGtWDWdWB0a5+GNyV
vWscBW2STfhg7P+obEIWW0Adb/zZazXNG/zHSpMpNFMxM7DrKEyNqkI5LB8PJmZQ
iaWS7j1gyokhvLF9kGeXs9cbl2lk5AZm5OwoLQsptPp2S8X72wuJqd0Xv5+qUtrN
oFf1ZxJtWphs38iafzUJanYEtCJb88HNEzpY+9fA1Ygcja3DvUnAEi7TWXBDcToE
7JY2zw4HWS/H2kMrhRjFEsCFcyUrFKacnlJ2QCkvT8O77X3bRhSaG5X2Cp0AHVCq
Ir/1ZPfiWwNNVVvXWqnTki21Nuiyb60AXv3kujT98iO//bFU2yQc+FflvtsOCVGM
rpoIGBr22LP5EJaGK0g4wKZXPbNSbqjNvygpIwPZcBbSV9PFe1a6NzNtxgLwMJJE
/MDmPvDsJy8y6FJYoQ+kwC4ouUWm3QmZCKQmi0DqYFq6d0++OjnuzoFiEtIzY39s
fr2yPdNSJCflQocE7d22vafiGuWDOAGh3sjVSYg1BXA+SjlJ4BmZd2g3PXZqrfja
tuMrNtLCdle+gkizsYJnSRUmTUOmv5QcvVJCaFw/4pe5OlhAFlsdiN/uYTf5kvht
l3hszFoAWaK/R9WlD6oVL6aBpQcsZpTUlvvBDr1bb8HA7IpRm9fTLWZLbospPiG8
9oIN3mvk+9892REbfHNMxE8gGE37NVs7XNB9oJrPrQPBFww81a5R1v5+R4Khpo4A
BRGZUZGRoelMTOVE0JZFPrKBDTjYStowLRnli5xz2GqS93jjcf44pWfVEmGBJwS1
h+gQy7iqnugF7hwHnOLZ7eT6WohknhVczbG8GyjXQfX3aSgsYsWvdtGuVfA3lSO2
Ful9npxkt9fcvagh4hWlDPgOtCSvTCf7ESmARlFKdWwS0/bpvkDXXLE9cce7pOIM
WJ2NEHJzL3VsV9Q9BLz9x6q7MZJztG12g1TcpTPKnd9ivG4M+ehqFmXevU4dqDsU
R5K/LEXOcKAZsL2Vo75nAlkEg66k8BJQE9ohy7v7x/XTbZOIA1J0toId+hu16qZA
W/mqq9TzLaiOLlVrEPGITmpmI3QnEUZHN44/NjdSEqBT3CO4ynt/+wNFXzj/fN3U
Ys/Afj84QuR3Iw6XCjJ3wBCeobh0o8rKPmSCzTHVQXEWBZ/+vhqNE68/Fu+79ycW
KhZLfGLixJVSG235Vbmz3M9NyfS2BZqPXPoQ+w3ktk9UvPGIWSNkp+0pxVH9vGD7
JhCXC9mJu90lJ8Q8p46w5F+mklhk/5YZsFzA/oqdlwtYCdVzYlJLI7JxPspzlOYu
0jcT1xuDZ/2diO0ck3oHAvYqgLd62oMUgRbmm6Dxpmy3c2gshgGn1jesL6Q95Vay
pzikB3SJnK8CxH1N8t3e9ACNvaiDx6i3hWmqyfWJo99b/3zTadWeEApWfehrMKt/
93NhQzEPMz983cZ7A8btDf3LXIqs1SUCjBnaRFSuXt0N4xdCi5lqZIcBJAW+pYHj
WDpj48MYdq/J5sAYPK+RH1zyxkflf4STT90kVWIBWv0RcjNad5jATYTCyFxB3k+K
wzU7R2WwmfnhNKGCeBVY7+/yGMoRBfKxah+WJnECBQnTpAqKKFNrUVAQDB4aQTV2
WDY4cdMR0lEgRqYQpmyH2XkZgzT/liqefAUPwAFBAmMcYq1ZMjvqoayMhXEkhdtm
9BJJ6xUHc2NHbeQakGQg4OzDnp9kC+CeGdlD3vaPI/vp/WJXmLsqE9qElSbqrKyB
2HlE1AaDhLnr5t4/lCuRjpcKkELl1QxVYXQ5Hn7wnonJRpmmD7DEwHSK/7aj3x7/
FMmw9GYBH7+Xd5IUry4G7laMcOBwGXTTJ+BBvlgNvGn+attENqPlWBK4Ez8ii/IP
E6Cyj7uGUsHzWxBH+VpW5d2WTQW3r+M7A3dSpfi8HJQf6JSZ9+de8xm4WB1SaiUd
7uiLTj4Hll2ayribB3FhjRBNMIxJ1YThdz1Y/Qszm5q9EvD7XZDPQO/PaQk2rgZ0
X2Z0+Atfx9pofBYG7bH4KKLoQXDfqtR8PiNBhfalKHX05ooc5tWD4TrGMSxcOrxp
ekMSdRD9yfvRvIX1ZHZxhY7LJiPtf/Ql09ZqfcaiRjBdMrCZg+WLNOVTwDMTOPO/
bSavotYH/aGqEuf0yz2zDm/U6EPU6ueTze5BHm46hlJctRNmpvRGU6t+hHi6E2gm
0LyyO2F5Zs+sQ7EY31Q1RCa4lkKLjfJD+foywZ9UwN3LJ4zbBnp1oIijViTsxppY
cNzHfMorVAfLuzQV6Z/8FWVLkaPSsBqFVN9V0AZmGd6WU2VjBkrtyOBZEmoieqxn
afJMYhr1Y6cshv1o8UXIW+Xzs0GDF5kAynGceS+v81Di2u4uUme5wJd7gG/KwunD
P5CjAKTNuwZRfCuXoooSMePAg37ZWWKIEhU2mcEwo25e+Js9npWdyQhtKXI/gcCr
7nygJdZy/y0v4lq+aexg6LcWJ+bIB3aQfwHB874QXxdyEGpdOWEFsg/cJb6zaoxA
bgE5ieYmslrG0YyuzJoKTPwLuFL0hTTL3DqAqXNCNTtyVZaMZZe7TyNPLysOMdEU
aCN0elqJC37y+z4MUhaTk/uLw8ZrcDzdf1HZlTUcovgpnOc4qtBT0jPjjVHCZ1wj
PE0QL3BHoRUpHf9EX2Xf+RlvTSHuOWcO7HP6qYRYZlhkqgJTJ61sN+sqf0GMDOX7
YXmG8zS42hrDrlshC870RfA4Ji/f+mS3hEIb7byMy4cTEfRnhIF8B2hRC0mrhinl
Y3tcv2m2BybRyMGh6+LpclQHlcKOoi1VZ6TIVp/iBIYYnS57DlOsKPPDV6LP5o1b
EbpbNycVNONlJ7mbAUMUDIIIGbw4Jvj536bfTfx8I/aQ7Nybw/iM9brtiTPUYjJH
O0a09oDrnb44xjgfTjbJmiZM/fQn/yxDevWqEl+FH3DRpJsJAorr1z73Io3lSRKD
pMTbuQN5nAVBDWZVMkp5BX+Y82zlFuOvjcCvCm/E+pDyAHr0TQN1xPa22PHcdvti
nHm2gDAvG2qQluWZ56PBQ96hr2vAxrXVE0lH7PiywS+HtkwPje5Q0Jh9WtVmh7/+
lSwYRZEYbgjHwIZb8tzqpJGADdLchRqXu3YMBwiyMm5BqQci+nmNgExB8joMFFAv
oXcoXVIX+U8cOWIghveG3BMN9qn1hW2fe4N9QVkunTPoaUWAyLwQh5FcQlEZ7hgH
k9L6W4z6CDKn+/hFNBsJy647lQQAFg4qXohgONdCEXamBr47qiSudTXcjJaDnKNi
8/ie9K1J8AwHKsyH9SU8U2Q5+zdT3CAYTFQTbBFm0Jn70qAQa9muHVg5VO8DvWgO
cn1ABxjlLYyI/L62iWxdISqaTafQI4GJi1BGPU7ME/IlIH6Ni14BqV/A9ta8EfOS
b+Ha63o2RpTpItIV52Wi4AVHta79CX1UOhseg+WSSNKntEx5w2KZgL9AXON3F7Aq
jpYmCYbj9xl56+WiS5m4yDXRWDrbdNq8LaRb6nFSu34KQO6wA8lcqCjlFm3nVqZE
knV09d6LKorjdEBYg/+2XYgzM7SM43DKTZLlDwPmcSpU2De5F9tgh73EUAYwQjfs
f5XvrEpKk1Bl78YmdP2U5eyFroiT6N2o7dvUFztKfDh1KJHE7X4G4ig+0+TZcHcX
Wske28cHyOR7RENrNd8BkXYOQKpF0zcRQ/kPsWDfjeW1WMBFZv3In/32lxuPa763
P6bmNDhY6qc8na6xQx0gjg==
`protect END_PROTECTED
