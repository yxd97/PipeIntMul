`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DDs60Ks6r+rTcYMr2YyncRAG1ZQixGnxGsvU2pHNkKKjtXO2O8j3w1h7rjjOg8pH
Fk6jNYeFANI7yofd/qfvOgD+hligcJpasPXkDkPIC/OOeeHhjgsnPxnrD5aUTLZf
/bt9gKSTjBtp4TC1GzAagufC+VDbV5HkNa03NExdKmCpWv77N2wTnF5DVxJXYtMB
KU8nMbzterGDqSRpoQefGyg4Oyqxg8SUmxFmZ6OENPy3iTALa2wiFZBfJBeJbsjq
VpwEFObxrtrhUz1YvrUT1QJ8CYGK0FkTb+KK9uJiI8gyyDVQ0jSMxwizA7S9uRHs
eSq6oKq8wkk1/DSk3xEfZVryOvena8Cg2vvPm0opxv9eP5GSrk6c82EyQbRZrm76
dJgHNKWBfVUhjs61Xpzv9l5ibSWFFySVhcejPeuZ8W8toAhUlkloDT+DP6JxTrvS
hWdhLQoDucBNgbHjGs/kp6jURQe1HTcdurQ7woGkLSai9Qx7BDD3R2jegrUos8Pj
E3sk4LoLeUWOi2CZkgxUlDM/oCuWF2qkpXtwh5Q40LVTwSIpT/JVH8U5yJaDEy0Q
s3+4hay+kTpMul1q4YuXbGYZPrDErNTWyJmaHJRyNauMAYA72pJMw3jzNXlpNDi3
BIC+nAcao6i+8boTciKvU3KjL0jTIAxXHXYkZPtcz7MisUiHvzoTPVwtf6eGdQkZ
AAOo4rK3mxDg46C9fqGvo2PZ1zW5ZI2AEYWKwNPEtIZ1wJHG3l63oXqSdKULPi0l
VkzC2PRjAbL5Ew4mtx2DIvsdsiGS+2N1ESYzmxRkLq3tmczIXn1kWw6WrYLIhJvq
zXttTRIF3fASTYtop6khqYjLqlPMLC6Xn4kKIej/SXmy593o16vf1E59HyJhhbpU
jNcgsKhbIUyh8HZ3LVzglg==
`protect END_PROTECTED
