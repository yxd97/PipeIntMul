`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uV+HFK5x5qqJgSXvWt7ZYp4kzhMNgC2bFuNlEqNibMtAFqWKlbqlpC/fA4lC0KaT
UL9xVKCYZV8TNpd2p1mV8lRQB8l+Tg0l/Iis/VbS2rrija2nnRFpf+g4iK2QJ0Gx
H7S8ZAjYNtPBLe/dliAyzWHwrYPjyp05JJyGUkpe3mHLIDz5Aow9HE0FYOsmdx5/
HBjuou2ktmL7SqTeKEKo3sjSE6QZVPir/D0Qun7CCsuKk1FRzQ+zmbbXcjdhbKdH
k+nmDesOPg1jVftWVcZrKfpTj+tIjyabEiJW/XcS0PmZXYYEf2giR8XRfYMyd/u+
D7WuvSW0e4AfrfWdM37ExaWPc6Lm/ozkBkOzmlITG8DuMsXw5/IjkPErRMQtOea1
dcebkLHvWdp8Fgp+b+TlcqAS/7HItYaLSeK/3kfYqwXyQIQX4IusINipckSokN6t
`protect END_PROTECTED
