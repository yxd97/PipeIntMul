`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u5fXfI4t3fA0Wk1guHYqgZr2hzjabaTBcKdKctO0VqAozhEKItmO+rXOubxya4w2
UxVHopOR6+PtrNJHmZZrtjZ/jg7OKlLRziyRaviQJna9GqT2l08tUCZtIBc93bWD
qJkHm5YGdZOFg+4UUrb3mnhj3NZ8TSl9ssy0P793JAQ5qZoeQUgWUNC7gR/mdNAs
+0dF0HZr5jzoQ59sC3PS8WfZy0DALjd/eMourBcaNNMSjYrONGxzR+AbhNnlgxdf
T3i1q8IDqT773NAvkJXieAAlEx1Lmgg5HG4ELYaysH8xBbzv/jLE+KMMwbRhPaNS
G6PjA5TqmJTsmImVM35x5rvwkC+9ud32G5s41F8qPJTDgX4TRF6jpERclM7S7EhR
FqS0ThumX7zpSaSIbD0oBIQ7KhoYH4kqb9jWUzDxjBwAU6k5fiJGgC521WfG6UY5
UAdnu+f5ssSHSKtzoXoMojj/w61tpLU3D0o5H544YhGyOq2JjRxQMs3JjtpIg0a6
4pCc3lmOOCbORI77bJBDuHCg0HeCvql4FOv2PQ4zQwlqnvt+sEGg/VvV7uEjHsVR
BFs+KJutBmaJ3ONotBLqNGJQhVgRHTGm6z7N/Kg5qSxyf1buSsIMoPoUuFLXhDej
Fh6oWrXS2ODJIikzh+0izb7HAnrmyxV+j7PO11Of9wDGxGY3MhPHhIBEpMR7JBv6
c3Uq6i8Scb4dSCb6R8FrLnKQPlLlouYknP5AfkxK0x2Ci7lFvTRSUEhM3Hhy1d2n
H4IzH5LHZnFEfKL7GymsAG4m1VqnFl6VVhnUR6ZLdrSmXZ6jy0fxvEYnDC7iR0Fk
4g039owPFcc+Y8SKPfCAcYSBmOzIMQ+n/j/J4JHQCLXE+HeI8ZzPpktkQnp06ypG
ZU8HkbybcB4ojjUicCzrmGBg3veuGDD4zgK4rJTefFkSysLYbOBvtI18tBOcRY4M
j9WIgZc2+afchxwKJhCQ798OQncafCRExFNJ52Y0ngtZbZyYiqFNLGthimyQ5ARh
omkhVIieLpZy2FTtpIYs1TL2bGTK9Ln+s1uI/5mbVfm4he/HcTj4SVsAOZHMxQBs
KxeLxQaNitE5tZrKQDmALA==
`protect END_PROTECTED
