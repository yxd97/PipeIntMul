`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2I7lLpD3FjaYX5clYZMIzFMFh+AellyOJnouE4ISmbbs3NCxESv5IJxnBrr7ID9F
hu6BOJSxsoRk7IcRSTzZ62MsPxRud/nBQkyRvA56kkSAOzsiOgax9doZ6kJYuGmi
mF2c2C1FtblTOcw2qOmWhqR7Ga3RXS+BTwn29tRTeb2LEM3xwypj5JRkr8rrI1GA
VOXvFPpRC094CxQ5qstUaIewpg19+YILe0lo60IlVhuN0KU68dTfw+UQqbfUdn2D
yZ74alKh+QUEaQYVDATxp9UlhZa7/sLoWOBD8FGbJSrjtKm+HNC2w1mOUkbOb7v0
MqBxmJtlepkOs760af8Jl4/UKhbMHbw0f/kqmNcBDUNMe+icxJAUlLVnf+X3CcQ/
ACXwWM2NHwuxMCdghNfe5MgXVU27J5cwfCkxYQbsu5FpokxZgrC4vB+AA/Ey3iq5
kSjP3g0ens2KvkzY/SG6f0Litr83vdJq9sy7ZHtaUYseaUhpvBNkXZZcQ+VFt7Iu
6LcNNVBYHZvqVcTtuAek4T3rQIRZVnvjhnmGvCVMnl0L3Rx56u8krfm6LiLe4KlT
9rcmhdSnmsV5/2kPUW09DeHAUGadzXeBnyGjlF2MHVxRu7Z+0fNhU3ycJrUfKR2P
yWL0ZML3fojht6Ito29Z7hSQ/6AeHs2lPGfzNN9Z7KVHNjD0hOnUjucqbOcT99oW
jjw6/rN22DppTJXDHq2h8mWuK13nrjmfmSfPHHtDeptlXX3jHXlFjQM4pjClEsIH
a30+MddGAP9i36DxTSi4cdvaB9C1fgcP1+MbTKKQkZI8CYFowFCnH7PxgUl6SR1j
`protect END_PROTECTED
