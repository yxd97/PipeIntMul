`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
N4qpzK1Mt6P8rpV44T2ktAIluYLCEMXiuB95XFlR7sW8Jkjfg8EF8Wxlnkq+39DF
5Yh0IejGNb+Vmjk3uAmy/F+rH53zA5xMFpPcb/THDeGsO4nR/VWBPVXkBNzzqg77
jr/epCXeW43/Ge+E3MYvb+jiAwKRljdWv5PsSR6+owiLstAFJiBA50CdlqE6NVyj
dj2EzwEattd3j5BCpVPs/pK747Bom2HaxyK4bsuies9A/6sFha9dF4iW/MwlFwFt
ATXwO5aHtYF9PZ08Sr4XMWQEKJeaiL4S53u/aZTTWxLjEhEyOtewltcHSEEtxp8Y
zGR7I70baka8omCLAkAaNoJUii+0m6YVuZazBwT1ha72Hk7P7qWOxD/AuxQGLTyu
/OyVvedBkOOJ1ZOGBOxl0ZeRT45Y4WqAZOMCdWaMksM0X2C3Nd9F311vpV/HJ2B8
8t65emUUUmlOR7LPsiMocustlyhUHPOgKneT6GcEPGM4LBROcbdYwlJj/ozXehje
PjyZcUAkziDVnwz41HWUQ6PLiKCf9zCUHhcIhlNoWKmCos2aSNwFo6MWOjEOQ7MW
dF6oretfwZNH9NE/pw8iJX/k63i/tMk6tWYXGzKQjj4=
`protect END_PROTECTED
