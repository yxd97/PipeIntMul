`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
616gNFwpyP/6Ofg2/x5uxelWnbaHcsgUnUgx0vjRVmzI2F0X717p4xNJHgLuiomI
z4DCrICORclW8ZFcUWdGUym2K/vhn2BrSvMrgQWkFD+4uBoxbzbRaGSpgy/EKOkB
WaKtdy3ydfNBdpFMoIJ+DBC+Istajts25liaGzbSteQ5GMbelEpELTf8pSMcVLZl
KiZWBV7cYGgU/2Zm377shcTwgt/ivm/7rwiIYlndz+EEf49jdAv/qk7qwrO3oixo
okqSIeIw0asdbH3g+kpHqHHm4ryv23yyJNhKiyS82CoPAgDxgIwKJP8AifK4nvEQ
GEwnjkbPaduZZdS93MFL23ycy8pKgNB89QNT/BVUKIyiY5yWLGQEqBd/Hf3EtNhJ
unIZ9Z3LQ+ujJT+Mh3F7wA37icankzD4FRcJJMOYXmQiekydlMkU+cu2B4xPgOzW
NcH5eDtDkyfMuopN0w6aI5MBxKEcsDYdUmlKylA35oGHpjX7HrABhZPfiDXZSwRx
Qx5N91gEhjMBPdgYrKwEXgZ3AFDG3lJaMiAOvYcm9cH6zDK9lur7sTGNs0Q6jNNu
5ukaA1o91CKsLeJARdCAqxYYmkk5ReWd6poIxGILBgFVJaXTV5AEQelOKHdsYZw2
MdHxyEtjxCYCUd8h08ql5y1UDK343sgJWn2lg4BjnXmJAJhgw5lCHE/hQ7FCLMlX
jdCCrmn/zRQYAAiJqqsq1SaFKUTFxoij8cRI9wcIXtB4i6+8Mi1L9zeRJaVtJdso
bSxVzH4KfoFq3sSZkaRqIBhWYZxqdtqGpsl+scat5z5kX9MYV7Vk1BvAQEBxv2pX
bUXZH4L2liE8SA2v2xE48si79gRt71HMR3ZmvJ1auKvhf0XQHEzMxkVDdzZPt0QL
24UIFWQqDGSMC91N78t4XpUmGb9eLSEPk1Ga/r9/pnlij3lGbRn7RLIDnV+0xrAd
oygyNQ0T9TZlly9oWLnqozqC0opghTq1CgmUHSPxWPAtzkCldt4Iu9WTevS9TaZC
TvFEZq3zfAAUyJzrFy0xPQ7jLwq+81Vxx7SGP1nkxhevggNOZyjD4/2Hdxyh1CFn
qlzoxDKGEJrSYFPfLuBIomWNGcZWFpkT/Dwss7lLbtmU+lWJ2fzW2mf+L9dFG2e8
yRuMqpABuoogrXMVBava2/E4ARK7s6R6F0HZLAT1laA6cR43stzkOgLiVsMeMq6H
Q6VeRJ01UDvzPmFe+d8pw9aTa33WMRDX3NvbDTnn2QSxxSaf/hB8ktF0g9rgbRwj
5jSp7jIa4E64Pw0Gs+M7/xu1LhQ1oLKYDLm31+n3Cz3UGxaYc6kpQoGeLRCg7CgC
9N2ycWpNcFvyVI3WCqSXMkQU7U6joTm6n5zL1X513ry4FfUARJzwsmoD9paESKGE
VrNmUKkXQjGZMyvihHSOfzRNP6Qr0/tABM4HuZTsGfxkFRes5Xy2jrg49ehJNdNo
gbcn2SooUo4Ub3NvMezl6Z59f5cQx6u/kn6p0n/AmqhXSfaj4xSDnlpeTb1Wip9R
gW/E5vpNDyaKi+1nql08Z3BlOhyscP1/JWJHLocVy5JhjT5cZYDGLgPinU6Mjues
V0YFNS7c6HE4FyMP4f4DqPY60w5573xVGSILtvb9EpX0AzAkOn6A4xgR9BhlPzEO
rHAtGcf4iV6zFoz4ckaWBZ69bLtRIKG6ImV5AizQxj+/XegiHzOdfsT2akTP9ItH
QI4qsMu6tDFkF1QuNT7KKxX4r2+tLIWzEdheawLybuwCds4overncMCcN39LKIMF
uzHbI5ndJIxN6DV1ewVfi3mEZmXKRzXXwoRwMP2xL0cncQrnFsDwTGLQ4bhBBNdl
pmsUhIZKzEzIs75BuFoV+3WndoymWUFy+zreQg4XSaGk6NHL2PTp7v3xp5mwuQSc
gsHqg+vzCnewoIPOMpQ4yCRM4XL6o+YkHsSuOKys3K2XP/Yxw2VDRJonMPzxTVGj
OTTzBzfb7R13T7ebu7gEcdxqxyPnoVpzUJJL4sp8WmnOznlVB6S+iNKYIsRdvk2e
5rjBWo0WoYsM6iMk/nsO1cRXFyXsydhdbNfMJsUlASoHLi41vCsyPjmAIz5otBsl
3fn6KfvOLjvBapiMKUGg17gMaXRBBdBeiOm5GV0USdeBrsLOUMLQzLjK5x4hFM++
e5lv6dzA6Dw7x6fv1UYlmnMzoH4Sc7sXOT5UnOGlaWcyGWhm+9VOHnr5KzBGjXI8
lFMJl/9r1fNNzWDxTc1yaxNwvgcJmWRwkkZGXnkWaIsZ0d5LtBfnmbWtUQ5aW42g
/DXH261J3N+gF0iDZk4TVjbEpLCj71QlzQh/CYPaQuh43fNRiSezooyR5yVbM2T3
6wzJylUM8+/oqGtkAD2XKY1MZg2ulom2TT/829/LAO6cOSxezSgWw7OKuUZnChy4
3L31q4/3xo3KmZXT337aUdEuZ10Y1nwmr+7Kjd8peg4KRXlZL1KQ54rBJ5DG+/ks
cWsgKwOIU6RhoIIPzKuMMYyG7Gxp2VhISrQc/a3+NUHNnIZpdZ8WQGY//XO7XIXL
kVJOnpAKT8PbtJupiz9GTc00baNqOnV1m3dhk+D7CMiSn/jwYjfmt5Y8UnYwKqRg
u/j/vuCfFc2tetJyQfJDmQar0E3z6JHRDXRoj5ozdLodZk3IPx/XZKLpOHfNd4O1
5SlpFQG6rfw02dIrg8WgF2KuUFwDo1FjmkBvhQ4sdWwoo2nIxmkKpBmupldLBCJr
F9DTEg941w0FzSiNiUEPKIVIfIANS/Osc8mQzqN6Afoba5oX4M4W36/xBfxX83l3
c0LlIK64mvczxTsAT6OZtb+lneQZlW1MVSyMkGeZ2NKPJVdCZqOp2Af8zlN7Ciah
FNFZ5tHp5DxTPDB1GvKK5eSEhcpSCu60PqV1C17ROs/WyrzT3m5neu+Ez6QSNZzE
D7SW6yfNgBL4i1aiUJUTHa8xjY7wqdhr5ORxhQoeZ9TKAFOpei4QpiKseBDcv5XR
utJlzRPK1qb2nnUL/346fW52tyQJpAqehJvBvYPCasdSio464JPGkpuNkxNBv3Kx
mXENotwmxjHThjEHamGm8ydyLBSbB7OfiB/h0PD6bMOC8nn5dZkVx3rudlV2HnPf
GKhhRPSKhOYNQ4xp/M2W325DOc2pFEjPH3Lln7mYWA+EyVIjTdbpiltVKZ/qinM+
+JIMwzxxD5exC7wuBbdWeW09zl6DCvHPzoNVPqYgHTJNyIdDdS3yPEGfhR7kLD1v
wHEHuhaZLPyW4JusFxHF393PXHm/8gixOj3zqnEU3rBPLnxhm/+f0vfMWeQO4HG5
GyON5/TI/xLXIDeFaZSZXGuYQyOjheto8C2gm++cgsl0nbd1mhHH1Jw1iUoWmJCa
RvkhVuB89+3QkgP5upbVOBZNdhMaFw8f2pf8l8dQ28dwl8vj/l2JaSs8SEHH8LPy
jAI7pS2U1MWpUPqxz1MFVmMCYvBaD2ZTQjqs5QgaC8hdoA5SHzv7MBa+6GAVBBeP
2ETm8okEIIouZ48Yfffa7G0ipN/tlOmhY8oVGXtgINvD5LVAkksPItL3u4cIbBtH
8xTh5WdtogX0PFcvr7spJQ5imVNmGg9d3bu4TlfMqwA841zTcM2BF5zV5wXI93RX
ShbmCtC2CIMScggRELFgvGrvpQ/Oz2r52MUDKaOgr+m86YVu81hQU0gFC8sXEC86
vW7JLCCTJDtAW71gEVzlRkcUKweIN+ev7h/eCM+sMvR496fJW3DgJo+kFHjWYggD
/4hMMCmV8xBaIInI35crlUUhw98dcMCA3jkmTEDuz32FZvgnZ+5g3dPxdb1sFBUw
m5r81gpJqgtX8cdy7Qr7VYZlw9MIWc06lJSV9LZxWxErW787m6RGgJC2OR4E23Qv
9bUM4aH6qyqPwkrD1VwS6EvSctXsSpiGHdheQ/j+YhEUSvaB+V749uA5Wj4zlBu4
WIyhxQEpbHBGLnu5RBgWP7iU+QjVUR+3YbHDKTs1QiYJyu7+QyMoIwHh/7MdIf9D
WcL8bGzRKL7pWugSKvgy3ziWhzoE5DJMMA3hKnk2hmyN3PD5mB4xB7c0d/IciDM4
VRD56ROBAf41KXdSBWCmdZW3YPnrstXsWMeo0qO4++bo8yHDHWcMAROBmKH8O6Q0
P9fer8Jfx2kFjqdKVeqmWq48dUFJ8VcGJy3qGRIe18kwS7rZld+9EszK0vXOplbU
VwGT2GKdvv4NVOFY+fdTniPOSB6xU3KCAAW3bKVlWU1GwMd1MBK3yr075O4UkUUP
EIC6JwuzrNQAtCNd8RJQcttJXH2pua4Exsj/HeMPNsBkdLz+OLvlRh9WCFlz8Wvz
MmwvK06f4rnLV6Zbg3yP5ajW6pfKx0iBxX5LG5iv7lGBtl+HcRrs8Ank8LnOgBpd
NithulZX0HY3uOh9dqVgHOlrMQElgWcl8Zdf7Wwy/T92CqvY6ZeZZOTQ6ZW9ezBU
R8Qztb+HMsXvvEPsjdZW+c/v30dot1FocmrQMZxfvtaXLoUCyjlYYPGknVZSO9UK
nZ04eHJ+Bxe9np+d76OmEmXN9uTs5wMlsTNTpML5r5Dd2x4M6vDu1XFQutHBjtzg
gLLBzZmp4RNWX7ds5HETA+6drsDRIUY3TpiCpD5jBhQBCfZ7pl35E09+fz/PN7u1
cK+Ckx5fBW/c8yXwz1LV/n4mmBkRoyplMbfn4ujYnw9yJq/oRohcdY1NHocd80ky
twFWbE0X+SE4YIal6WMxOva4YMNwBQS+Afb8aMAFDwX9ffFvCtOi16BkbexrNyEq
nt3HPtd7V+Nf3o/P2FniGcz2gIfpUxu5M5Iveox7ZgvI4p7nZwVhDkI5wlxKsHvj
dKGY+Q7WKxxTI0ntQSpo7r+FtCzZyJIYpBbr0RpUx227yxbq0npQP91U57EiWasj
EjQewJwFdf9uhHvRR4tZKNJv+uF7s+xlPZCnww2oVwhpKZ/IOOqbX+8jtqrj61an
h0pjueIhpSBmsKeHrQ3HWimK9W8UE/Z4IbfYPQwABdZbWm3nR2f1wdOmFXnpfaQS
jHMmY1iNR5Xc+Ap4CQCsMldswt8r2uKfDrRWSnB2QxE=
`protect END_PROTECTED
