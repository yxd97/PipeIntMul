`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sfyuiaLDaj5gu1PJ60rCzEd/dDVzeN9zhyeQDrOnRYyYdh5q4M9YFoFSg02SaEEq
2xIBqwznVzYbp4nk4lyLQckhtpHZuZeW6B37LBzcCOllTyOBtuQ4XZkLxM2poIAT
CR9r+qkR7ZVFfNB2DT5MabAiW4hKZqBBoW59owD+wZ8u/JSqZl7WRvwTI0O2IBB3
KqHCtSgP06CVnCNTm9PkLw7oX7VsjvyfpzUxYhzPplGQNGSohTEYRfqQU7j134+T
2CgpBsQNwjCJCMl95TmRmt7zcwS/Jp2N5Rg6AjweOA516u8RnB722GaKGzlJmTCx
OZmRgZUQsIkPFIGyioe1FVF6GmssYulq+PRMmGr28yHPBZPkIxQGuKOi/UojqOq7
tm94rGJvEfZCiuzJjNHvv5He8RZ4108FiBvfYLpZ32rzszpCFHQl6bvZrejuYO83
xyx7hyCWceT2AUkpRkIpW0bDm6E1dBTIHfUXjHpCRJ5dmfUv9a5DoQfgU2XHciEo
2gKkCQp5GnZ7gt26+OBMZ56uVQulddg4O7qMqnR040fGgMErwWKbSkQK7jBJ43HH
zz6j/9nSH1oeUyF1Qg9QlmTUP7HMayVTDi1ssHFLh8sI0iKhWhgv0/KEwCS9cIf3
PulGR21iKUr0GDzUCZcI2TgSdH5ikWmkmwlCQBiOqw2o9oi8BRKOenFOKJbXIsFj
VF/CaIrHkll5MFRMOyEuFtg7adcEF6lTEtA/tqIfCa8bHspzhuTNn88B+1UfMXVd
/KXjFbhcotOrgHoOhPueB8Fqm16W8mVjaSmfwyS4vX9VuTX20nAjwDBu+K8GMnKf
cqmLOAm2r1H2wffOy0wSqLIwfQY4qawVKBV11X6yuSY=
`protect END_PROTECTED
