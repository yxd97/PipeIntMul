`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSrIzQahknv4q2tGRhSxAwiMIDF26IvagTSUhGegl5wF8b9uV+FU6kh/RgfVW7Sn
nBLVbPNQN9dzin1OdgafxBwEfUULZDE/rT/5aFnS7aComs3Zo3OTrzstdXoJKpog
iEBHORNLIFkuUe1FyM/RExDS2pTTJN9I2YMZUOhuTAGVwvAu/9I2Mx0uANIvHEui
qMvxGhVaCa/hLN5NX1gW6P1iKfMw5Ibt5ubYC7P4abu0stqd71Rf8mtZmvOSGZOt
KGtLfNIa8mjHCrkyAJhKvHV7zX+/Zpj3jGMKkXfMrh81yabCH5E/cNV2yBzCZ5LM
3Og3Wh7vJAGlGs2acDsWLj/zoKB/+d9IFkJ/RCfHDppfWylj8jSLzUqf103UY3eS
8HSQqiLLt4wa+U1cYDFDh+Y5woH4AB7izuNc0ERCM3nsXY+W8Rvy5JKRqubcFSHK
D/xH5zXRfH67OIIKovC4pV0DYbg9L6atuBkTr/CdDf8OGpSlsDNB15OmPADXXM+Y
M0o2svyhvCjox/AbZDSjwn8SVh7I91yY2VMEuwEg+kN3CWaIjuV4oAozZ3nLIdEE
hk56zx/YvXy4WiZkaYJW/5TogRmhZJe8tkuxjJzKyOGJui4Ex1pCDpJCDCdzNtbX
Ti3M3IX1gCDAJvgTsNrLh1O4jWgr7LqsvnR4L+SuDU9kLAZ67V/EG2Kl81xuS2HC
eBNJRQvg46KKnm8Tqp3J5R1AMYqjjStF5q3/65u+L03ND8NcduSQ3Px/IX6al2xj
El7RayleCSnTitIS+5r3Mg9BxDnMtpiWiKeR9jBpeVG8PEAdKKNdnJnt+0WZ75hX
PDECdyxIJ2hI0L6es14UuSO52WdD0HZJzepEbXnNCRlbPJFOvezoz4hffoSfMmY/
bXkpIDxTstWLtFecyal1c1wkiHfjyZXnvr3vqB0hlT4n0xLg9uRgGWneCEX6E13L
PW/e/7Tlmf5Gl7E9tnrWeVl9caiX1KAhFOZoIZquepUEWoD4lD16e1k+licmxZAf
OoIJBARXeuhy9j+ZWD3B50H0okVeihQAoDRb0O2JI5K8APFfjdzeBuEmPw5M+Xgb
Hs2rccjtD5o7jOy/Dm3gJw==
`protect END_PROTECTED
