`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xziOXm0yZWHhjRn5rIc+pAgWBYrotdnzIKyKvtPRs+8wUMRNs3Bdyucd7EDuRWVU
tNW6uGbEU0LI+CmuNHt6/OYQQIXgYkVhANjigWmix1PWw8VIeoMxCAnrjRarue4x
qD4DSEm1MK1/iRcPt5Ou5ZRheVki/EvkgSF7AXM3o3ZXr4nOvBFat/BiOJdXZFZz
PbveYxhB0O3mYU7w46AnT3sWKU2nuVd+5L9a+e4+Gk3u2qtyCzTNKJr7DZ49UVuC
TKEfKRg9UkA9uyTWopb5Xe4ZFjvWSTFiDzST2iJVpZ4nx1LPLe27mBu+bRC0fn6A
nQJY6ZGRFT+cWX/TPjZSpw==
`protect END_PROTECTED
