`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rn/+iJ7fdq+o0WvjfoBG/PtUFzNEllrXHDu4LqBoiZE+3r7o8UYIMiLewILds7kE
O7nxSsqUwBUlr9OplE8hf40NKINEAVpaX97FehkXSOnTenGcYdhG7+EiFH5Y34ci
TwPlPTZ969hCA1lbmS2p+HYFte8jSKohtvVwrDhlGO9rG/eIeAAjI5Uhtu9CAfvF
94oW1he9ocWqx1XZr5OWyyRNVtwl1707ZPdGiv3MzMVzujgX3+b4j8axY/5ptUuV
/ImNBiRCgHNJLQpmaql5a3VH+d5M9C4PDmARfNIHNou0CspxgYITEKH7da1Jk539
2WUBrVgeaEj5r90CHmm+QC7hpSoga0P+yw3s0dpFeQusoxaGZQWPvxnqBjOtalHQ
cZtmWEEdr7MG0qWEl53G0wm+pLljzU9GfV4YBFK1MU/V8NWqb/ezrHIYVfw93rvS
m0WpqeZVSpbtC5IyxhCbZXkbfX78Z5jZoOLl+eorSQjdd1LhDD4JH7MwhvR596o6
YmMR7OZ7mdiIAGtVjXvoLx9TBbYVOtiPNeJpH2lsrBn6SvrA/Ws061gr0zcjiqFP
xg9fPZix/wI4uxfybbmoFWEQI9Dan0/qfcbj51spg+h9mK6n/yUpD61kt867wn9O
6GRbQCqBjuv/42GFucbn8lHW/tKLoyVSI1iLBRDZXzCUTlhP4jROz+SEVX99k4T3
7xZ7iSVwP+2+RhNhKrdaPFH1RoJ7w3qy+bhp23kV+RQuRDzjFeJebW3u96FMkrpQ
G0fy+VIywBmBBXgL1beHJo1MXafDaaPuUJ9IgZN+OZW0RR4fVMKDjcWqVsjBd+lA
a4i7ETS1NRmY8rX1elELWaIGoVFuw1bHHNuL9RQqlPtwyYddBllV7AtZvW4bYFr4
MF6n2qryIvgVNfsSorZmbbyM4OXaw0lTT+i1k0hZvdxbXHNgWmlNy3G5RAHF/NDq
/gf8+6YkvofkdRsgnl+Wdm02UTUaxvTBitOH6ige9fMIJIw4w25wbFxQTmT/LI24
M/1CW4SjEkGdvMFxqD0RAoZC5ESLBXegATXzwEOl4G1yzuUa5P5+xwYbX56o6TnB
zEbKIceB8ySet7+3/+WT47GfNfKcqrYtPxmjPOrKrVTWaFrd9IK28sXmRVYOL7IU
5CxYfCPVSAs1r5vO5bgH8qe/g9ze4EHWsKNUPJ8qc6svnGvAcjZmjG/mOQRCxGS4
d/wfn2r93UoZ6LOPxhsn5iBBX54Rczgg+hObW10g3DcRqoXCaaGCitqTsJGZYumF
CmgqQxO9nfnlEmZYSfFVdxNYmgEid7jZtQYn2AShKK/8aweReuiGzV7xUYWBx++X
hXSf5MQU2QOnYiyVxnPfP84QXqMKaYg6LMv6DFAbZI4qXczq3wyWPUwF+CaS4bSK
TiS5HDxOXYVxRCAvG9vrObqsqQP2eO8i589jGB9EWiZ0BeQ2Lappbjvz+Q+IFYsh
/HGAfMnEuuI9zoPieqGix2Xbrx7VSyN/cc6mluLBOW72ZRW722yqgY3mLDQhBrYf
gGMwCrisPt34NPGj1JwLF7+Zhdj5IJPiCOYHEKXocAFtgsCsmdTeU7HnzsIq0Jb/
I4WvhlrDwTDlbQ1CS7WFjFFcApY3cwA4vR+ol7m7SFaUhJeTXQP46YzemmtYiLQm
YfyL95T2Alzh9xf/phHMOe3SvS+wDvRhiwSLxqRR98YTk2ffoca5aeQFyx+CBbDY
z/rhRqZ9FGgB86lSDZOWRpImpxVHQLHNjWuTOiNxGU/aFIijXuWkNzxVdO0RA2bh
rkmrXduQzr+rmDUr5XyddMWEIzVvTfqeRVwzpN+F5xiZvzaYHokccoHVy6OQiJv9
2I763V9MYLdQ7qMjUYDhS0erLCqcRS7SuQV/xlaY1LgJRRqcBQZW81LUvjQm92Kb
GawFJlSd8CsDiI8ZTCuo6j+FIlho/k3UK6EM7H7DsDqelQpCAxY53dU/jjOn+x+j
Izfvt380wpD/dMUlMXwxgS+Dc5By4DRsg7frntXdEKj7KoiQcY8mMrT7q3UrkVmf
HWe/yQvFs52VDxd1VBEj5J8fhXMja9BVGPnXmf4WD7AhpZLKS8qkvyc4tFB8+dc0
vEEr+NN6fUoDkBMHnC6QI5KKo7OcqRwLYsdrH3NoU9UwCcyDssw38GgzylMoRTgg
Mx9SL7IJZUjrzEm04a9TMyg/pCP61NHOOrHlqodgGzTsfSm8ZeHG22fGGg5kjF6Z
aplo9PRuKfiPqMf1YfIktmGeAuUhno2Lam/6d2HzZe5H/7eCWMjM9yyzSDBVy9TN
C3vuJbzBD27dYpH/ZhE73MtY64iGY7fEgryqX9AvQ/V8ASWaJ24lUpv4tfGAmUle
a74cExamFmq+ywbZS996Cfiu7+re99WrTeI5r3WpLu/p+C8/CXXEPLpED7L6lMU3
dBEzaQWkaMiBjIQh5NRLVy2gEHmthxSxyqEXENDHeLm+XQp+DGEFe9jwSEPw6Y6V
5u0aGErmdubFI/3OO9L6KPJ3tXMYJ6cojVioWna8LTb8o9PREBxywRLiHzkRWXsI
gnp/oyJjoDeFN1OOGi8i/3mTo9UGkSh1ABJrVDfE+d10MrfX85Cmb5hpnGrk8aHz
VI8cG2B64Um/MjbOSuWwyKX4pbnCiMYVaOhqJFBTCKQ7EtURf83sopDv8RItjDYe
Ai2fjAkRDmxD6i9pjUC9I7oISgGK2RHoaIA3RoinqIQOPhKRI3AEPrLmwMZpVeZQ
YsDgfau+3E55hFPtc+ZajusyVKWqej8Wwl84ehD1LM0PdMq60qqyHHFyBoeQxZrC
EJyMneGw6i32m7Qt7eq8Gg==
`protect END_PROTECTED
