`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7NERxMJqpXTO3xTF1E13Bv7RPopGsnHlySP6ccdXg6Z7JkNFhDiP4fnyNy9XnVAh
H6v3pNBEHwHS2qabq7teuUgbvj8Sm/xaLxJV52L8Bc9wmxojEUEffsqYlyDqAYKx
sX73d3W6Iod7JUz49tO4uK2lacNk+cn6yvl7ywH6fDOFA4W6OOkQxmk/k01h1M2c
2oQiSp8ZzD9Oxpt5lpMRQEMLL4y+jZwgn0oX5PtWQD6OCRJjruMXFm6MMXv5I+IC
`protect END_PROTECTED
