`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
d1xYQNdVxxsqbp3L8+4j5bFrzfVP7DQk4J9pjzu7TM76/3V2+rLoM9+VP6Q2KR7n
BJKDdd+c6d/VcT03bEx2yzxXTKOMf1Wbwt8hmU9hGJ8ovRSZGkxV2XbLTVPsk+Ut
sCzFABIc+bY+Nm+NV/eG3GtOkFnvL2W6KP2vHl1ed7OKt9ZR1LMLZmGV6+AQ1uWX
PuO96aEaUOd9lpuxYj8ToKVZjD5V/SFLMuxSctNjbbESFuzPdtC9Jl8HBVIuNxqf
JmJjwpnQ+l0dXYP0aZ9+Tl+NAPdO+PR77rljiKzTIbv6IAA4FvR/WsBegG+I0SLs
d3U8Zq8+giXefbPP8ALAbegtukX00SLirNBLMx90TMNZyXYOWMcun6BkFUM8h15d
Y0+wzTPlTw6Wr1qPSOAu1ruzfxB8wJbcLvtNSPxp4q6cbMD4zrLJQjkUse8UdH/3
dt8Xnqq51Bsx9s4f2xA8aRbUlMdJUDQ74OInn9IWxHwX/Esi1vQ1lWg7sWoXsWoM
pQ3nKbOSPPg6IyhSt9URNolIg3Gf63EaD1ZZZuvouxXHseQKgkzPfzpTZ7uN3xaf
ufYFcnB6cwmqnwYP59uZJl07VSA5gbga/b6AHSBlXaXXljZ51vPa+f47llP9BjYo
755WaCrz1Y7iHXilyFE+DFEA+4+sFnwh9piIlwAmYzBmQwrO/gvaHV9oPYZozMYL
o86XEWFKfQcJdIM8/OIH9L/XJs1283mKVM+NdIt+ARDc1tuPsMIrfbobhXsqkauK
5+b9LGLtZ8851eFVPrlnm9/VjEnGYlJ4zMQbjnhE7UNp6yN9Q6FyvsHLW4Vm1HQ9
Xy8pM43ju1/XpWdbOtMhZ5gw4m+OIBFOm+dekqI8EN5Qfl6ppUsvvohywsC+JROa
jOF84jydXwupA4dtacdHLw==
`protect END_PROTECTED
