`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PjwxiAHr5JEsENZ8d/TbAaGFFpPKncoABGeNLy0fxyIq0TCmCWGpOyddOsZM/9s/
bWgmkPPUlpkvboVNWDSh3J7Bh/Ai6s2JuCGa++60mie7yoit6Vdd7phRfFIKOrX6
duG3hSaiimdkCDKo7Ka/ZL4jBIGwFhSsa4AoQra4morQJb46vo2bYhkJjdU8cF1I
PtUqwgMkGiBQmyCs8VtBFUC9+pi+WqrpLFlWQWanx66ERluBCTlWBGqo9Q8/XSaF
BtJf1oozT+wLqWhntm17taiOTPqVY/nl44MEXYE3LPoLYqR9kzzQhqCtvQpneJma
SHiAQv4AlrAmxZMx3A5xkHsIylxGW531hreu3yy6zNugdlcOYTeliiXuzXmflLaJ
gsh53gkG3sYTz2BfM8D5ugv+2dLuJ5o3mDgmcuFWGqY=
`protect END_PROTECTED
