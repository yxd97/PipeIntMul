`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5Auf4S1cLvzR4DAIDgZy/5NZ6rPrbLPahp7J/1mITqX1ntW0j2NjBBYKR+I2ChM7
S2Gk5l/TIbrmuVgvv/trosfmcS1c+ArcPBCKXvjeiUgH3pFcqjRFJfAPHfKHFbcS
Zoa/RcF6bMogWMaoutqI21ZbiJG+sCnR9Q8C0+E3jImGMtfVrjWWoj/tp3vQbwLe
QFGkqDIPAIi/+e9ipL+L6V9hRUPI+VRcDbk4v/kagFNrBPC6TfLzzaICy5ZfScTi
n8uGnA2fxZpxFSmtjv0dsA==
`protect END_PROTECTED
