`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4l3PJPnjcTqZqIandBJ9ShOqb3HZaw57LYEeii3jsnlU4PJzkOrYVpxB9Dxx387c
72GsWyhNekAAs3bQ05DKwjBvethU7vpL48TBkd70mgXnC13bb/cXt3qWiepJEUFC
lAWqjCkAsfQY3+OOMM4bdHlSGCtXtH4V6sdDukB8LNuaDuW91HW7v1lUd5W/SRma
riQLZOKRi5Krhn8DQlHd0mwN2UOKCISQbggevnW2roQqBjBobXmTHJhtCo27FP8x
a6RLodpbw8jhUh3RW5zlo3Xv2PohavErgV9zrIEonlkzD5/aNlhY7752NGXJSQxe
lg9eBKTjggJIwMbsuVOJqGx67kPvCJnE1y4ml2YNl/zWGHhBl3z5TKeUOEndWmGq
MPuNIzjjkBqz/Jc6w3wr3kRY7A70dUf1MeNcM3V7F1t3MfESvu7Kh/bUquHzkBlx
hl6XEsHYTmL+PoH6EjIUhcJaZdwwUx8vP8fQvwv6TIylTi6YCDhEySt5L16fmOQq
`protect END_PROTECTED
