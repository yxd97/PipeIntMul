`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zfkCzTXbYRsengSrjcv6f2HbaMLwOOO6b6dSTshCaN1ay2HktT8R3GRciSxEjNjp
6WeCGm05Q/YfjJsGAeVQjaaPmeA4BHJ0i7Kfw6dum005Buh2pQbonZbYa3CoA8gk
uG1fm//faW8xGss3Kd0gAB+X2RVu5yKYuEGR3p8gBXXZHDUqVpF5h4IgNjgkGMej
YwIl8SB9f+x4Lsthzj5Bs7pDHhXpOg8+wk/Xhv4ai+JFMDCTLRBIZW28nz/LCT8h
yRSChTyNC3Jk7YG29SSgOrX0fKhR6mMAdPFnK/jRYLObJhvD8djVVhLXiuMjGU1E
3vt+3X2dtms4nc3ZuvirqkpvZtk2CGGEgn/moW3NkEV7gYNDAcdqjWea7BuGSJj5
`protect END_PROTECTED
