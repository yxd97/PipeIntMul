`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0N3D8vZe/vJJuXEK5UqHQAEsfTkKNyAlHaW5CR8tzgkArpOB2xmS9sb8Mqly6qZm
Bzm8vKKr9JDee+VcNeiRlJBC5WP2vIJgkBdkWyJpFwc9JDxnO/2KZjoyrCLrryd0
eBnD/REcMfh8ee+o+kcRTasuEYFd17NZD3ocdb3911yZdcUtkzgdebQyuh3AvbkW
OFPt1gtztnKw7CAdMCL59/r92c8/GzFVKAstZL+ftUgcvvqX5AbQ7zrNjdWMcloZ
vaCxVJgZ3XHYSLtRcxiODmBsQjNF2L5PekYyX5pO9ei9mCmiyLpRYyudeMyHlVxT
tDQt191Dmr1twTUf92H1He4VuK0uEo1m/aAxKg8CngeV9Lp2Bj2s/Qy8RCfcG8od
gjHKLFk3ccgb6EZM0UHz97z3ymCXF8gQl/BqRykYpbR/n/W76SYDko9qzmxsUbCJ
A2HgpAXo70wFjfQZiG8Su1pXq/QQh3JamYwqpxeqw8ivs0zkt4Oh5Mz+spRSvDQu
bfxBkUs3oM+hV9oA9h54jVbqHAP7S4nWGgt85wT2OxnZ8EHoe1k7ZqnK3jHVa+FG
hPr8IZ+Y3rj7hnqKytrt14amlwQoXybcUD2ZjUdEz1QoS2o8bVVMTEY980sFobw7
DkKTkq/RC3xQrScDphPlMorhNPRx8VXDhOPBQ6+5FyO+WARqS3uidkYlACUwhmp8
OYWRmcF6iEDjeQQ0/GHwSyGUCJVl688d5g9ZImZ18MwIALKfxMFm7KxcVovAXg0K
MmHZj5GLg0WKW4r3tPzebZcLu/BAf1A/1cZL9hx6Os+Y1FZuTqs3+vtcXo+0v7Vh
CiiTfu1aYAoKYcGnDPLNQA==
`protect END_PROTECTED
