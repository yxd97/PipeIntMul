`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtyKl/TzM5AEXNYwqOc3g8wdJoyAWbpE1MuUcIG8c24qXaap7HKTxGsPVxinEJIT
xf4pgcJxNLTG3rNN4XBRTdXeOgcDTtYL98uQMXxtupV0xjd4AOdxryWkTL7xoc5I
kWvxQ5iRdwRdlH0UuqIqkF9nSADbBDnto0ib/iGBDyJ633QLYJbfB3X44cLyeoes
RdzXGk0v4cp+mc99gcKzwr8Zq9gngtz2jfV08tWooN2Zplr8iJ7lpQxRG/NdSiq0
ijIF9Ne7tKosuyOEXy2vlGrjXiFlVElyTksFILnPMRplROrSsgMYwjXf3az9F7tw
/X6pGs6R2kXWI9RSPblUPv47cnqMgSlw15AU5XCbmzQ=
`protect END_PROTECTED
