`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2yH9cTUYcly9eObM+uR0e/IaWP560KfPCb6wqjOHa6232zDPjWrom2HRogtTqYRQ
EfplrR6XVYr3x8ERxQZakLL/dcm+VqeieNmntpiKXQXGtdm+dAigcPyDV/Yzy5TI
DOF3UfJDXZdXA8gfSVgmLTgWkGKbAYY3JSOh1mzFinDOqatAt1cOX6y4msMPyBhP
oa3GXeqVB2KY7A2eBCc20Zgp07s/F4OOvC9wt40La5cyXs1sFbg7K/n4aT92ldZP
TPrXItXOWGHXMDtHprRrenAu3gCcE/klCAZ2XsJScXMxr+BmQ8Bc3E28Dg0rGkml
F0sMx+dlPi0BZgJyk3ges+8IVPM/gZLgsoNgofoHmkcqz+74XZUuFVx9z7zAVajv
sCY7EX+k8kEXnmftCI6Q/pUenLP9tPh3mfI2XTdGxbvU58S82hwLvpjin2RCF/bQ
hgCLiuPzv9YGlfGdbLyKWI4OYnLtjJZR/I2yM0YRHu+aeKL5y7UEMsGz6LA7n95G
Bcp6V3cScrUQe6BhasohEQDtqUmDZNFR/Btci1NFzDLHfU+lPNbTKkvRtWNN7TJq
tUxgQ3JAWYHIoXpBPScM6xQzf8uqo5CQa7iFLnaqOucYMRPiZYL8U8h0MHKoBOcc
cZ5thY+3uwZuBM4Ab4fPf2ti0Y22omVCqg8nPTBVABUyAUyEpPWZwoHO0sg0UIZO
MPP/AQU1RkM4YvBXvQBowO6EDMoIh39rmGKQkRk3w6ppReW/+q7O1T85htTjPpvj
3LLTRfLbbQtWp4bU2JyIRNbl6A3cBU0pcHWO87VS3HEOdSjIOsR0zxoQcb07xYy5
TPCSoFYYvGdeTTT+3RCIF+Iask5IRf/tz4M/yU3pG7I9KHQNOGNNAWVgslSnPTQL
YW6N5ihPfhNgLFs7yLAt90Exjt4Iv6iI34h6yEY2O3+MqBkODhGqqB3KGiHSZyY7
xSWopSbJaez6gbglis/7MMNnk8TE8ZMQQAO/t22itOKdugu8ZgGT5RC8+uTgObaS
jnZCgIxcMqDi8bLvHyWXlhME4ehTlAubDumTclvgTgJgqp7K8LpyDkHEsvwwUEIW
lnaJGhac+s34L7JjHnicYhEQScy9Zuol8DsdvlOG5w335RizPQ6Wwcy0n3g9dE1k
85blg9ixeT6xwzsjJp63CJTfGkTeS3kY3zps1aUm76udWPX3ntJ/Pn2OhhAO9Y9G
6W51C/vKFP77tpqXjH82fuKlpdX3moG+OI94ww5A2r8L7Y7fZaRQKOJL8WElOOOR
CWHOEHFKs1LRYGrul1JQAHzyh6i08m9oTHsbu+H70jtx7rE4JObHFfo+Jkq2txUc
hJT6EuqtyatF2aNUSiC4PsljV0VRiWbg5vojELWzdZ1urcy/0T7kvszOTCQhabTS
coi+UItXB4C3AXkLTH843KhfFJEGlwXAztmtDNJEblmPgFOcLzVDd5kT6OOU0e8T
GR9pWFSdaW7pe5K+ChGfYFn47T7kyjLcC0yMoaX99CABeMM1/scqP8DzDireUvkB
Lg3P+pZ5qOAIW0ZlGEY6F7eo2YDFPiA8i/rCMyLsRr9W21VSWCm2lrKWMPG5jKo6
rEGeyusLfhw8X85h4rYYNW+aNUE8PMGeWk2qM2RAQC9Fn1iLqefB+GljApKrwa8B
vg7wsQCB836uE1S6+w3rjTB5xZFGjtNP+7B5WZ4TwSMo7LLR8pvMeoAQgIHEyhrh
1V6EdXgBCUlbNS4xkTs2beNCQr+fDfAM5B3t2nZLFDcyYYoU9xayTCxK164hAz/4
Hr+a1ney/ui1BjwNmqXTV0XXgmUkyDXSMPQczwlTTL6K9sl+gI0wPx0Mnz0iczUZ
CNwjXzRkgRZgFIbdvN0x/o3E1yP6cfvYfzGZt8rHqhchk9gU3EDubobIU6uHptVm
EsIBx7GY0Ettu0sTE6tU6wXJGlWRpkVzm1Arxq2ojOVbEEO3MLtDc31NFywivheT
MXae7fYgmpbDg9sLw3zsH/+OV8nh+gcUJjHCHTSH7zoVEK3NnDTqZjOG2eOGgqPZ
807wsLljWMXlbhpth9CZZIccnTg60SUQga+krCM4htKUGk9oRf3O5TQS/uN2vlRI
YvLNNfvtd3LfjJTj9H4ELsWL/9WzwlUarO+dFUQt0Sr0TSgozbg/fqMAd9mFTI7L
db2hzi9Yzz6fBYFLdrwlgO0s9jTRj+b+ZKzrvZT+RsmMaLslTU3Bb2ZqzntbkDum
PN6A2WvIH3L+i4XWiuOvTS/l5Uw5K1+63c1qQg73JuT6Xv8/MBuAeeY/7UDhr/3J
Yz5wfdURZ9T0pgR7531zJWCpQSMQKf/GJaDBN1gpZgbRhSQw6m+XGIL5rupg7U55
CzqhZaBUZFdA9VW20oGqglfhFhBgRB6zT4KLStWhJ9zu5a1qsybUaKjP1SDI+l70
eVAUDi48sY0n0hLcTTLAlK5fwAqMHfeJ31Qu0fRvYI5XL3p8j56STRXOWOtckVeD
AyQGsECIuj64cKfiVSZxl/Q3ih6sQGL3IiXBPNy2pvLFVEp3ck7wViJgryh61Ssi
MqH8XxPAaRTAn1FJHMM4lA5xwhcOZTgUrUhoqZuuP5gnPFeqMHbT5+NoPHRpHwgh
yOlj+WOb33QWVifIQsPPq9MIjlB76HE5lGn/8GUwLuv/9Hubzx41JfGl5KxlD5i/
2OKpLTJ4d82ZcVZi3ZwSqwoHWuKb8itY2+A9UZcMc1wtl8STZm7vFGIU4qFecBVk
zFAnsw82NjJQTIoeErdxRsq9hZcaYBsR38Flze9/2cutcJqLJXJkOuydUhgPljAY
ER3TQjhxE2P+2kJF1tQ1pomZrDfxzeQJ+vb7qAG7c3qYdf+KY7FKjNdBuh5B1ek3
VY9neQa9Pug58lVoogPAb8ttq7yZkryvDOtPZreyBgOt7Preuw4Nrsa7DN+v9G9H
B+ksY2BWy4zem9nYIl7mRdUpmdkTKbA+HSqJftVb4yUTlnfVXlXDF3KiStiVCQC/
c5lMubg2iSFljbhUJiSAdAokoKQhfKLTyiau0u2zGgGKirJCh1OjmBzDrIibp1LR
oxmWV13Rs4Boynv7u4jUPiirD0LCTkDX8l3HZDLwgcaOKq20YUdk5N/LuUrPqj8l
21FLzBWRO9gCT4Pw2GKzvQ4+4z2/4YWjCbpdzj7ij4d18WvlONHsO/NGpSo8fVVJ
Kz0rItGIgnPxLeOWLdLAbNAqFvWaXq4LQfx4UuamqnIyhWibtq1F1xysjHpn32KQ
/J1DA9dDOn2oRT+PfNzTrAILiLLz5/Shb6uvtaaVujd/C2oMnglrzDhvpLyZmZS4
o4NaRVJWKjVpCaX5FafW1Ngh6uttV5+nJskn/vZqC4ziC2IZx26YUTX3p+kvonhc
YX3fi5SQVkrV3shRFBpZdhyrKS5UVM7GaHNr2rWkGHy64Rljw34bCHuSrND7lUJU
GpKhlLou3pzeINER96YdS9GRcuxy3QWCA0pFADbRzoaMwhTti8UfgEZCR5QXFG8y
49qyDr3nEWaGASFar5fzgWooA4U+w1kpkxKqZzY5WiN4r7leZvEAs/BgnUHCfM0G
NCYxoA4XbHIkyWeg5hrtXFUtmwFo2uOF7zI9/qB1u3fFJQlWre8e37X+hBgUAE5U
yMwMtFvraXTMNKTi/bBx8XWkluz0hvGD/UTx4jl0T4/CIGKpok/syN0w/Rm81Vbm
iPc9ZpMhgSmEtYh+B0haLo4KZlkGbPaDOU+GyXjYNlcCZOoBsH+51HsqnnBp3LjS
2fuRd+v0U6aFiBnvRY2754uotsF5NkfjcbMuM/Wk6bvvv8iSD9Ho7kWbVzWyaO/d
/HjaScCk49bKco/nr59ossmckCA4wUD3pfk+xHAb33PWu9QTCwPCtTQQFtrTcMN2
RIzJvZ4m1y+kq0zaxv64ToeVqr2V8hjjjJqlld1VDUtpilJGELiVTW+PXEQxjTBt
RKvyVs8Pzzc5o50koNpZkL4du7J+L/7R2t9wVAHJyBWPEqgUMzVLbVeozgnX0gss
aRLSQ1Q4q3Hy2feHKpxnQJTYQTQiKoMQCs+ivIu9ZuHpco/+/wI+/XeAneytovOK
XbGD8nBLy906S8af2EiqGdh/42iTl2EG2JdGVis/E3/bCKm8y1P7XrxKgyIVLkUY
1Cnn7Siclm161rZRm8zfcYz2vppZM7t59xvkKZhq9YLWTTzrwVvHejKd9/IoFXl1
bbPSV0Psi2ACWyeOxDhorAKZ4PqNDuWu3Xr3TV7p2em4r2dUcPFW94a6wCBPy3g5
zfhlaYsTwpiwe2ssuVpjs5y9Z8e75UmgHt5GJc/1/pyzplF4dDay/EKpPCSkVZpM
heBpyo7ee2qsmIrbrd4lTRnSH8RzgV25nkg5UsQiLAy0DGyEWvbXJIwIwIxAQPo7
DdCa+98aV4KxszJBbWQywWXGK62Pxq2nzoAa3n7qGeJ+eVfX50r9DUNVH1wK9Ua3
inOVs83AcweDUOYsRizI5KH5M1iAtlHGQtErMw5O3qcL8p3X5MPSmrgMFz2tr3XZ
TNhzmXP4hEPQC/m/6Qo491N+7UDocguWueVqbAZ/omd/fN6W4e+UzxPiXVxzPet6
d7S2YRrNGUNcKwhTPa/k7CbrxOz7HunbrgEUTSBO6MR13b9diAtUuvjPfvbmWGD+
JL3XspidV6+zWI5wjHdnLlsLtOMl3okuu0GJE0crDVIAAPGUN5/oDRUegI3CGp5Z
UHnMcZbs9yHXZb0vYrECNct11ui6C8tE3RnDimvUsJzCvl1Zgil3rCs6hoer9KY9
T2gBRm5lzWFklPXx9+jZEhv9mwDFa54TcksPSyKn1DBQDED2tHdHlAD0XrgnREHX
G0dn28zcRaoUrvJGBe0/qGj3oL/qWIXRqNnHuMhbuFd0RXnl69Vs2tlwPBucz5aa
OItsHRDR3iRPA/YWzK5g3ZRCttUA5uJ1wulOEgqryvx5B5X6jg+DlDtGND2URvtF
cpQl+TlHngAP31iAsx55kCln1PjMDSkBmG6iLhQkvQBbHtZ6ZAp34x+ZPdUdIp8Y
zgZNuGjwBprC7/Hs589+RsqHww0fFl7fdfFzhX4U0kg8Vnr837umxrs8vIRe+6m/
9dInV19u1g8KYjl3m0u2/3QY156nRqn1r+f9WgYMxziHvo4aQUNpK/3jxhJQEqXM
NI0KzX2QHM6sxrvgYksvchfRhnSnPM7TTr9OiYz9flnZp96zzpnXG830VfOHpwqo
WbM7noO0Y5eSTbtFlOJhxUnJklYY83hNLh8picVwcXN+1T1k8Y4GOGsQT04be8eJ
bKKb6Dexv+jEp29l7MzImgPGFJb3EZqhmEMlZeZJH1MhWO84cuuuGmSKEbQLVvsQ
KUl5xDjLzBoi7ycadUYx3LuwvzhGOVjZZ2fYgVe1eFLEl7B6QieK/4PPMi/uXIZm
0EnMft9rFU/vuyvDYYelgaFyukOUmPK0iIQ9O/SbfMVdj6EM0ExT24h93bfBC0Rb
kgrJnQfnT1j1HI+Ri47JWX19+RNGfogZoWst6HY/WO6wrB1G1xNjMj6KJKdyEGaS
Vzdhv1t30EKv2p217SBiq0bxvOephqOgD49BSOGb5nIcHmyRb2aYlB8wVvUZNvau
GhOu6nNs0STFVc+Xsx80mhaJVx4teM20/hptxnQt/KjwYW4ab622u1tvUizRpl4w
QMbONXKZoD2m28xiWQEiqB5qYwGOLmvx1fkh5VHlAd92WGmIPb8JYPhvwkBhIC4j
Z6/MMw+AbKqKA6acY+BO+yQSrYXJAJmPgSE5NmCP30Bw4J5h6adp/m7JpXX+DLMV
svFreqe5vqhS6zGpKHBh4OWMyCtUQnHIIYjLTI2yWqCuNXgyKnYL09oooo2ANw2k
pS205BtsT/PNY+u+5myqJLnjUgmCndmPsHsuy3/7NIyO1uEqqqh9ixRi+dBCK/6g
UJI12mGg1C410RY1aCreY+pqy5G6QZrXol+qxtBDSUpFb/RY05PgWPXdtOWYTRpz
JpaGs78FVyT2CPJtl3rXYoNgLd1RcPuPjJnodfzVUEGxPZs0KYqU9EhBgpc5fB4z
yrDWAWWFya2yvJa0MfEHs2FaAKhHMUKpXunEPH+Fdj6WyYhEz/gewPdtJF76nW0w
mVAaS3isVjS40TP5OH97ywwQkxipTVJpvwaBCeyWTxXSQAZMI3UzRo5Figgete5q
XZOpFSw9AaUYopU74PwNwSAZTv2M/LUtW08DQgXwdDz2jiLrlXxVshco97W3z1u2
1YI08kuvIsnfM5JRPJpfjwg80AoZI8v3A6UApLM74Zy7QW9dYMnVx9R676bk/wB5
G1BQd6FDHn2m9LigpmqBnTvwh8SWhgNiORC1P+M3jJHH57d0jK/VFKOrevLPCECN
Gh3hG9RWwVcZWlSwfZJMvZ7Ad9qdQXAD0bWQ+/NjT8SelsRzcLhvOLGWHFKlo3k7
svCcsujc4edQ3a64xx6JYqPob2CcoJ4VWyBbWPWJ/UHInmpyP4CimcOceD67sUHA
U69rX1w6zxI/Ld/6G2T4WXAMWRUprlaW0C8YVUFB1qQLV/9SUbcu1jkaZFlL8ky2
8XOzJUnafHUE6SJFIQNsUZ8kUORH2yDHX1DhcUAPopGp0Fh2QXp/aZzyh6/pz0D7
CI1YL4WoWhCKf3dIlmC34qN5xSv56wYXVR4a5/99jbjkbkMHRaHS/9/6VtxDlW3x
u3QSjyIvoaAejX3f9P7BKS1lHduW4MvNV7QWpzYtwV+OsnhyYOgNEvtEAwrVsiUX
nxnBVHzZzDWD1wmW5S1HxRW+VU10mWPxDY7tdH4zDIV8CC7kph7doPGirgioqBMi
XRTtb0hqVjfyOPT+JmOK59a6J+5wmGzEeMVE4sUyM01BMXIlwtteEkPK+VqEC0qR
sVcteI85dxCiIp02WDoUVUE04WQd6JeBQTCbgSTPXN3bNZ5GPhrc95WTsmC4AC6P
fK9qnRPpL05jVIsnAJknxuShLlGrJz1MIquMc4DauLM5tePZ+K/IRJH+iOwJBBhA
BKxfkiayRf+zGNP8dPLn6TuiFBhjElmWa7p6ER488yXx0X9spyCh1MMPV7lWzJI1
9M3mTzqgqvcJvTzTkyvovkH30TyGcud//DB4QHzWUfb+r02qechigdbXRHMGPoGC
wmGkKzZgY8lcasfGFjKFv2o5O3oeH/yLZSh+FvcIIT37N2+bZ4lh6LyzloKnkavJ
2hvpgxwHPZ8nVlpBhYwcokRQtO8oed/DHR52K7hK976wvGwkBuadaXkP6BmTLzJq
fJLauxClG6AnYWD8MfXzHODaKAr7+udlGD+x5ALZgTPJ1fAypTiQmXFv5eAL523c
pQPEDHAu93QqHJRG19ND5+5GklqOe6BGX9IrwNoKlD1tHtCi8Cn4KP+PY5zIT8sX
1qbrImLkKwCtvzIJsJoWBG0N4NR2t56iz8wc+kLJ5LA5cCKxsZc4Ah8e2185R6g+
qqNxq8ttN4SFNl8U6ROQ/xNgGRd24r6AScDB+wuI1oMjnVp4ZJFruUjxqgOF5JtO
QYGKZcviTJE4N7H8rFhc1V12OB2+uoHqhpac3UrsDJz8ArCCBgj7QTHhUULcQFqX
XzMhbktMXrl6+10KaEObQheE69jfD/w8ZIdGQxNTC7edSMXSjw8ARs/blffy19et
FOcbVcU9gtjHMsEnCAOCqn269yRYndUxtWA4mvdttb/gdCWNUjS5k+T7ZtYAqtoK
adeqQoyxxb9QUVqht9aAvIAcDbzydTFgTGaycrmMnjPvuFXMHs838kVqF6dpoS2Q
hQTeu8GydzTPbOGUvqRDtcIdGwksKOdVKm7wOAYKVze8jmeWEAKb95Sqh3SSB7Fc
6USgei07qKT/t8cmQU+gQrdmesh/yt8fl1il8WrDTNeayFxMSIC00CibiKH1PFJu
VEmbemMT4wpZ80GMYZEAkV3+yqQSFdz1i4rlUF6bCIgO9oUY5MfjPtfwnA9Cv2En
J2SCSkq6kmDmjMj2j4dtNq/neURET/cRhupTdlvvBmQ+PymuuRMPR1AnEVsH/Myu
epoC2bH0iUFHNSFbJ9f0TRqSiiIb3bWnauhtDfK41p7MA5gv2ePJZbnvSy5ghlVv
HzhEgccdPxtUiyIXA7b58PL1RLNjanLRKPG8J2fK0mSZIWVgQx9n8U2N3hiBeANu
xf2fubWpSjbFy5MMqePC2Me8dwKAfvyLFDyuBveioKBwmO8OlEEjovt5g1nSL/nU
KDJiAlrtceiztChHkmWY8v4XobqRO5Qbh4bq54xDVA59bDZO6NL9OXuu7/5QzIUS
ygbL53aS17BQwf4pZ7aqRcCtjY9a7h644RnamPRO8xlAkBcef5TBKbypjHBLvf0M
mmQphs9UV2w3rABHEk8tk2cWfTAOvy1RpOXRNhtAiyrblP7LVfNrA9dyf7HKItrh
g4KE5aCaKT2oYK/z4l6BBj0HkJx9zBl5uabZS5Uahy46DJ+3TEU901WvyoP+NbTt
o3DD6Ur9GkUaDzRsgIOj86rTl0snhQLlz5ADzCUzo0s0MfHn4DoJapgP4ZC0zgvP
vp0gaflB/7ysVAmylMLBakIf3QlxTGDX+sx7rFd+q/Xc4o9/GUHDXMwxAuJfXJoc
cpVYOQiqQcl3UXoCRPoIVhgjj7CyO8Vk/W0Jep9PIJZa/lIuOmiIk4mCu0UyoZ0Y
g3wR+idHY0PAGG3x+Ni1NCVbAFLukdvVk0xXWEQgStWt6xT9GE/4oPSnJ8f456B8
GiYI545Vos2R3d3j0pf65vtYxsRUA0j4eIJh+g3ccUDLsBAcVYYk1+WbfhcOstdP
4+BtCDwrrHQzq29eKyjutRH95yB8Ffzc6Gz/qAXMlaJJhhS50DqPtU3QYW+fzqKN
PMgpbcVTAX4My4i1fg7uGl/QG8pGpRno/I8+Ju8sfimBOiLui13yyQK85rBlmL6I
7fOUOX06hDdyIAkFQP336Ln5PQrRCpllnT2ef32RfLoM59AJFwXpm2bpsQCK9yH4
3cm6A3B8vCiVg6u0/gk93XFbeoyonKQytVfL2Ej9Jt23d8v6AxOlM5eWR2arAY1E
rWXnwc0g7cfl52k+wQqh4I1vW0F9BXXEM4wvDEXia0VdVR+5YB3dXYGNNutV4mhG
Nobgpj3yT+KoKTxb//ALAnr47iZglkQXGrVq3gpx1168aulTG2NFvJBwZt4f58rl
i2+6Kl3HUrK9j1e7Cs+7fDs1AUSN7gtVi/FxY/vIK0yCiePPYhOrYrQM7/hLrL3l
CfRdtSH4v6J/OgZWeiolBxCP14/n5TGQiAVEjGdGERhy1QHrutt/5NMN8w9d8HaU
E0vR4Oz1gmgtHNK3glhzafMVkDbX64pmbJTaMvsKRvtfjKTxHQJdjjK2CBpNLVxe
e0w/edaRaknNZJf30keAOcd2MFPq2WXndhVCSL86fFlOuB7Us8kUL1UXQqrv52+r
hbBcBdyZS8ZXiktD8+DQET033bx1W0YjMbc7AJmesoXV1XcfVX0V1Lsp1s9UFdLK
NTXeIaUKZyRz2GA8dbcjX0LOqW0DN/wuWdO9i+k2fvxEqSD07HDKH5EqDPKjQLEk
/xfV+9vgS49Fe/KGBIc2+644ajBU2meNCauJ82d5XJAKhean+/D5O2IRaeRJNTkR
aLqcqdrhmxSxwwgSi81OkXCWaYq3/MpkBDqbDDC7s4XUKHTP2Wkeb3En6hUAvCed
PLBoGNVjFbTB0OGFGDaFsIKJC7vfG4FbDF3Feb8ixnbBWk578csqp8nPpj4nUqiD
w3NVNLXnM31gu8vIQbJwXOzUSG9XHxRFi2+v4ja+ojPQcJtz/CHVVLWhKiZEY1Z0
gnWU0Jwsi+2B0pmC0UT6xZJJRcuWNcaq7JaAayFQ8bZ2gBTI9ICfTCjnU9FaCMAV
TZsadfaKGXqAuxRQx3BX3OZ/GU+EeSIi0q/YnQyqWKJdnLLB8FTjzudLYxNB0z5a
GViYzLNZ6Q3dZUNQw3E34PwtiVxaW+LxVcfLB7RvlWgwD6+MwiY1XcWDF9JruCwg
XP8MVHQBEoD30CnksrywxgmzbkAOYC2gEqkIcZo4d9r1Lo7Is56WXpqLFGqwSNCq
/e1eYloxBhyhBfK+W50IVFrm8BHmuMKE5g30NsU4YBzvsrUFwrUtNFeamrgA+eLE
P2OJvXTTOleL60yYtLG1fUZkhN2wzQnA/iWsXbDGbW5pmRuTRofRzANyrzGQu/lO
AjMudFXkN1B/PuHLT7qruCX3c0nigOQY3pRmHtTqsjczQRFUg7HktkbUTntcWnFn
5cKW2GN2G9UwtIUlp7FGAHPfuAd2FJ43tfFd3OhKPRoReB6Wwp2Mxsviel5mopbM
vPbDtbYv30Q/UQhgJsuBhW5l3YkfcY9Mcaw+eNUTL5qEICrqQShU5ZKMiB1hq7EE
fj1epqzhkxZa0CjJz0t0HAmIa/5yvp8WVZE9r4iLm8/JMwJqFuMX2pU0AoitOv0c
IlOpgiBxIMDA9WEPcb8i0n9zsrfpwAwdyvEwnp9dXS5YRHxOlF+Q5FHk6lmfKlRA
O1ZtogrdTXiFovl/g2FLitNlR4CjaN0GUNeedUS8+8T+p+s6H4/Ln7JXkYIcrrbj
up0nEKvr4LRwJV000rauTJbUMxF3KL8wvA1WGDtC7UaplOOUZ0/tuBKHM6xMj+io
zM5RMdq0qpGNHJdnXnmThBozSrbRIQA94O+ylfN5V9HnTriWFekDAr6JDUzQNGGF
+EReQ0G87JD9daljWzDiJPZcXDkhPB6CpY1c+PE/vQwHhWXhoQSOxb1cP6khkIsV
Ofle9OVmtAKy18yWCs8BVfC3wYo1P6eeGGVTRwMJvc71Qi6ge556CrGGb04wV6JI
2fqN/ylQBpulYp15pTmJVnk19w0jodQzXK+TxDbwe1yiEDLLoE0pDAPG34SSsQV/
Uq7+Q8qISmWekdqVpajcUH6+m7jqqvZo5fnMWUXIpsDEgmt+erSnPvnXbVvw0rwI
kw8XY+/SyY9YBxBtis0DCQFCbSLIqj5KG5Qf1SM34HQ+4AI6RTt5ADd3U+b7i8wS
MJG2VqxxWULbnsaro9e3vSToVodhxxlbmSpLasnrToOHPQLxz39+n0chD1u+04Ev
iGzYGqAJV4KTBEtFee94mOwL11VOGzW8/gYkAbpqDVW7qv4HqfK5+f8vcYmFQN6j
TKdS5q7AQF7Tp32nas6zVyLg6FkA9soBMROB31aidCDqqOeQ/9Rxv+ksyBBGueFI
ETr4c95JKjg2iGrUToRlOQV91w9VJSXkP0fPwDyyeEpFbPuxS9wokQX+ndT05YKk
YZkYqbmZUz/QT2Ozclzp3qn5gTm1+lonK53MypeOi2wHLTpyeqLX7KSlIN5dqcXH
LzGNn9R2jgHZhtMY/R9FR8FXjZBcV2o/j3UVqlLw2vI4z28dFsvV0dl+Qqna/0yi
LkS8jgQIM/vQdLQA1wbkQLhgh79XN6HlrYmwwI+8maSXmQAt0t9cotW8Dxjnjc49
eKJ9vLypVEVZmxWjrWm601AOW8zhWFi5zsrsiEWVR+bJff64FAeYJZuKvcI5Kfvv
2A80r4WG+cm2BOBSNKcH922AVa+r3Tkswwp6ZpzJ+285Lhd4Z74KFAvhXIdI4bw5
1OBmsAGbKlxiFSkIw1//K9/6mpQaIVjAZVc+/9EP4A5ZxCyp7XSVVlx7MAxnroY8
5lI6cgQ2PTlzIKu7PNdP/VBF9xdyRX9ogrlElfk5tqtLr8WhQtMhHofGANw0+GBG
whNJiclBRFmXHBRKXkp6XVH9YUrKor3ndkwK5l/UQ4JQ89S87RwWNy5eTOE+6ZZG
XsPp8FkBvjEDdPh/NeNrf6VPZeZGsHWID2Jt6MYAJC7ra8LDQyg83Ohl+3wuhdHr
nxK45EEQHdSTECTcmzchhvIV8A0Wp+MIN7zxQCa/Krko+xs4+9vHn1J73vLQ1hiq
8VT8Wqdc8Krs0M/5bZFC42rhE9TEAnoJXXVo3TFThleqZZb3vfFJ1nkl0cod6iR/
dDywR2g/9/vbhLywZe8CdKlXmY+kJV/h+zZf5AFBcGQgAy5rgdJkADBm57km+rsB
SUfyG28YszHu0HF5IYcKUVCbUJgjt+rTOsqOCUXJyQ4OcJ4OjB6qLp9rvxaC+U9E
R/aeE5eFpcL0glglpxvIxMHkoy8RxoYXMJJW26tBopyuQFgGds2YWoPPgz8y7Laz
gIAuJrRq5ThvjgTSgxOaSQf7PNHhFamTSX4NxK7SOds/+mwZtn3iIMBageQkEoAB
lgzh2vHnNKHHOn2JwmnJZedvBIsMoy/FG0UIk1pJFmEArX8qBi3AfkqT7a8qHoyx
Dd4f0/UCR1WfJhl9WRPKiOOZFEZcs/4qP4rToJjU2vZgJ4orCvdsSe/vQgD38tbS
xUYx4zx8ixk/vxRtsGh/OIw/g9bUPoKm2KiY3qzfXWuZW+OrMYQL1gQf5ge4tOFv
xHiludQX1hKD6np3VDzc9M0XwGqiZRW8pRD0nwHXUARjRoOQlL5dKGgUOyunTQ1F
mYuzZPwJO3MgCMGpbOq/ACtaXnN77xvrSMnAZBkLy4k9RhpLWpzdFVD6mIg89jRU
9gJJ/pJgBoYswQc16bsvF8PafDRGCIjYU6x9CCpetCmenj506ibhDjnLmSEm3hR2
iY25PmFnxrwoeHNbjSVNIWO9YYqjnxgtTatTuLyZjFY6KH5951CWSgiw2/rCMNs5
PLUux8d79JUdyRSlUvQIiROfk5Q04xpJgy+Kxz8h5pGBNuV3Ble3R+Tf3W1mauNZ
qPwRj5XuxuALFZ9PucJ6Y3yf8Uyrhf4tdhqQYJxyyjaFMFjwsF41NhNYw5448/qR
Ub95ThwzxLutBAV3XCtvPFb94LBxJtfIb+Urg2+fcyvPNDzxPZekHHa4e1coakVm
x0yUCuNCTDPktYW7lL3IX+jb22TeDG5Wyq68eDl0zy/MJAw+QvVVSAo45+9Pt7UW
EmSvMkVugh3Zs6+8Ac/1vPmnGnkLcw0p+Z405+0qaaqPv6CnsVLnG5AkMKnJXoox
as/6LWgQEsZDiWf0ajHB3u/3LhFm45cqphiSlZ4SU3gk7crsOUkX7NRXJkHmBU0r
CX6iaIC+d2c9znf5taUDxMbMy/ExF1e+FwvUB9D+Eg72ZU46pCSiwwlm5MNXBuUh
eFyzTKdiKhea+XhCUqJgtwWPMeZNWFdOewzRSabruKb5UjTmyitq5X+mMviVn6sC
rZ/jZbeSkEYac8pzLZ6CRtspP8KndneKlDRj+BX5zJTAX0Ui5iFVOk2G9u9tdQLB
NVzp2GosXMUFroZIB3eQt559DfKOEnh0lHpyxuDd/HayPG0WH044tO5z472f8p+M
Wet64Ot1eopuKhqLLPnXw5JD23NNiBoUM/mSKLaf6he0nYeooFYpEL6p0q/W0ave
90y1WpNHUpfl1TL0fb0EG4DT0znaAf3EA4YV+JM21Zmn0GxySzWvAjd3RcI9wcJV
2IPVzTkqkCWEMJziTZ3cbWjLYZYBnTKpc/SgVyWLxuCAbQhYfip7i63hhCcp9JCU
Z1eMhm08HQkrB24+SwFmuhJXQJYM979D4Cek0Z7tslhiap26uD7LooYM6YBFCE9u
e4c2qP8es+f+UTvg9rH5nsqfg6MGJXn05XDkBbj2zu9XF/D8PaLrlsI4Ec6KT6pJ
jHOkPbCs0haDt67742peoh5Xlo0kt9FV8A6wv9IxXchB3m+rUmzn8Av2gK855imP
TA0D6/lMIlBhN+ElL3bMO1AFAccuOV5u7e/lOdfN1wYkavtsh4oIgN6kBRGtYsZM
zdqtedv9JfbcvSBdEPyRdz6sDAZolm41H0mYIb4xVn2E39CbpWQW3h6PTc+kC4/f
UdR3jW9i9i4FQwvSjGYjxBiJDdd55eMwKjmfsZAKNQfVsV8QSKQuWwQfQLV4r/61
NN17JJFo3kAcbilxEDt3QauKHNxMr/H78IWph5h8ZwMOW89a5jMNdBGgGJPzqNro
dPLJbiVVCYtNkUA8wUmlX19Eqh3GnlDacQGXVi8AdHogdYS/1aRQulKvG+Rq5w8c
Cjau5KT412VIUknmzJrizsKenlRJhq0i15dvXlMPRDsY5mseb8158w0Vc1RgXYRz
JNVhvzqBoGzeSLhmlh9Qz1iTTaduzxHYXmO4DoVLnuw6pUuNTls4D6rTd+GMPqMW
nb2uNiGMaBTYzGf2KpV4H68/9Gibav472UxvkAdnudfw4m6O5aLG8X232vB310Vj
AoLPl6WTGdJHzhsowKJwJ+r0OQkUUqiuPUks24D3y2o0L9ACIchm6UqVboDXu2GH
BIgkLAQeDyjudo+vt/u8wnJI7ws/UjCA/ac6GkoHNPVOV1JxzLwJbl88bHkPt++u
5+/I0dvyZkECRqVHe+uA8eEDHU1mqbfnc38pfgwEAeqorAGmWAJ3RxbQ6LMljNKA
3VtXVM/GoshO3Gg2NYXxGz29x7cTuKkk4wwfYQZSgRpVixt4xN9hYYCBWuYoDnyH
XvvG7QY2g4KPZA6kNuEwzVQWlQ7LTUaJ9iR5Pz+hx1AVyju4/chFZSH39OZs1Sfq
cD/GKGWdBk+TRghQ+AROv80KeWFkoZVcswW17/Cst6FyKXqFScFuWq8Ssh10DF3D
grsjcLOtW/QUkendnX992aPq3IG1pRhQVwk2ioAUqdQiLCsJT50RGyeSg7OF1iXA
W9nkudQXvXcxjefMStJDaAHjSZogINk9yAwecT/uM/SAgrJlCp2J1ltVxdVlQuA2
gBix6bW9ZTV+EwrNHgMxug2c/kQCAISjkFzCRKSHwImQo/MXAo94BCvDq6VqqX23
bNjT/V820d/HvDS+TlNUaUSpKRESKhHgvcgfYI24CkYcLx8ABtcs+FJh2xk3qhHR
Oqucc8tESYtfNEHXZmpEEoV1Ulg2fPuWBSjLiX2tgcgqspADMmCOwk8lVKfpq1XF
+mv5rZ2bnHnZ61fOzoDvR1JSKx9EJfP7fN8TRarF+8CBoz/QqgrNrxhHZseL6qW/
z9NU41nkm+hIFwvFyAnzq0SqKayKDVw/4sBz3HyEXCWJ7YT0fiNjbpZZMME0cwU3
OytrEMdqZLKXQEIO6SlIMf5MiH0VV3gb8j4IGV9lJgLldKe4XISdkbXeLmlsFPtf
w7cdbx7vMiioGxfKvW6CNUSPm4tCgzfrG3IqCjLr8GaKAq22Nr4v6effyx4EVJKI
DVyYWRsYXog+ckl0qrApWqVvZYJxg6XIQ72E8G50S/jBdNrTZYBldOT9n/ZLMPnD
o1oYG/x6H2bORxGTnmd7KZTqigvQVUQJP+TlMLcGtKOL69GrqQBatSSJLAg0Ero4
1bXx8tskJBEYej/zLyZiCcT8rNtboInauUbsUzeBcx1BLWKnqwYamZSxf5ZskzcM
rzGFGprN+nKbJu2AdBaj0A23wlVbyMKX291nogAKcHqV9tGU+84VSXbpALJKgAxL
WGFdym4mkoy1djfDgfO9ygqajEsf9gFqh0o7fTWkI28GDMT81Ca7BcjyJh7Z2Tn7
bi8UYl0RfmwhW/icVP7qDcoZy8NHPjtu/uda9bNH7hb6Pd0P23qpRiSRYKsh24Ir
qpZ54xmeUNcloMdoqdxQK8TRza/VR8I0aYA6jkQLD6u7PFy7LP9rkoNU19AqrKdA
w2qhYxIEwpKdYw8cdJWD3ZpBxXrJTQqLcESv7EDTA+120xwMjP8q0RnJr3neoHqw
w2Z/H0DBTdbg2TW7CZU3Qx3k8UD6bnum3KH9JZ47RZn3mpsgDDzOKpsw2BjrWYVX
fVbWpr2GguRZ8w9mZCAuj/7tlsSt7m7xQMwYaCK0GeJWnwZlg73nFSeOpxRteUMU
BMZV4uZR3oGrfwKnk4mrQVtk+5aiu+Vxf6fEMT5P9nw6srKBnhcKEW6X6REFGa9l
zxheRNRxnNTicbxKrrZLL3yZCWSAh5sikeqhoBXcZM81H1FT5Ww+IjGOPkDyio8K
nDfqPEgngkcxkw5/UUiDHXckAg9hDdY8xv5OV3pwVfC1in/PuBI87PF2nsJsJH/2
yGLRyOt4zdAn0XZRy2valhrBwACDjUJDZGCydFjUXNhrUm+fMgk2gKEw9k6S9THY
6oMLrlC6+fs/LcjOynyh1eAQq5GELImUrLVJigGFZT1Bq4XNDoSku9omG6raAVGD
eVO3AcSiq5P1iHYCcpdVv99NK3NXSSnXBTq9nhPem6Ro1/WcPIivQ8igZjP/TChd
8rXaGQnwikDQONTY3zrYu2PbDm9Y1BjWiXq2gbtnKV7ayX5pvGCKT+IdAALzAUlP
kUt1GsMb/MLP4OfyirCyJPlQEes791RDOB+cE9pJry9E1k+5pScO9Jdti0Zw6QPY
14Q4k514IMTFPxLiuWZE03hWIlgd4C7wGBZ/qTcO7/x+ptEo2SiD+k8a1RG9QHs7
EpAWiHRf1xkACvyUm22UrhKfOsaZwJwteb8M116CvYdK0sAa38wmEhey5co+9nRL
ITHBXWVh1j1dud4Mgz2UHNGJ8iWav4jCDP8QFMfog+bsAhp6LuOxSotxFt0sUlnK
JWUTv1BhXM89ynKu5L1uu1/+LBNAaB0UxEHaR4JJ7ndi3aiLOg5YlOdJ3wf2K9Gj
73ISpTG/I2P/s3DfC5m4POS8CFrMSOxoiFn2SqS/eVezOscyu7A5rSHfEgEFYelS
weBt+iu86niWxYzWNAeh3e0JQUPH33ZjkGEPCXXE+lFARcurW67uBS6uC4aQJvqD
u7tm3IhGMb5fb7Toq4u5N72k+2jiqM3KwsQ1yhK29ybc93NNgjyZDaxRCKNBjmRS
d+uvUpMd/pM3ba4yRVQ/HEIrSGgrx5PBaAS7bgxBI7SWSGYNwJprJi6y/QMapwGW
1umgI1pomcTSrJ0FDNgGHVZZayYKAcKaJlJGgeX/qu6CFYc+bSRrzDsgKKjKpyeB
IwSgF7k+dWPDGAQ5ApyfZE7S7wm8MgvRD4KsUVucKXiP8zQogAH9GKAnXgryLnLh
07XS5qOc7dJ9bkPP+l87QEVfPVUgLi3Ip0VBOevqyAQwsjBYNtL1FilSqBV5GVbE
l47zh1+Eho/cqjZpm4XSnUJGH4EtNgfL/EPLqmGpcSf7rlRrXMRSUKs3OTHGHHwh
EDGclbkvLUG76y5yQh0jYX1+LSyjQBGaACK1PEnrB3qUx1EzyN8Lho/PGnOqRpUw
LCUKb+3//63sH4XhZMlxCl1XgiP3h4vk6G61w+GBNp+GW1Trtxn6yxq/HYa2jfGY
tl0UsYGswBZQDAnXgMNN8b0GFDRfcddd3aO9H8oaO3l7BCfTvwYSeY0w67A05xKe
VZjbv2eNTsI9SmMFdB2utB7PVG4Gg42uExBk6vZCyHMmKSbucbNplf8oMgDwllEA
QmIys6Dao2o/ALNABzkLxNgQVxsJmHAs08BJ3s0lBKF7Tj61JqOQ3ppVIXglniMc
OgidLUNSBMui+8E7cQD4rzmgy941T8v2k0nG0S44oqLI2fmD0q6PwtD94PzxzfmQ
RWp8xhUe5csmpnolby14rha2JlAle8MKCIDggKaTZmzyeWdveRaWz+N3PzpzVr3I
PSa4MNpGb+6jIO3aDRATw5i2Af2I+Fk2TXHIcqe1d4OxRRGGEalZkZnOS3Ql5n35
N7l9dBCnLDYAtKJ5g62We1iHnlBPJnb1JlBz/bNY/pRDZL4ihJ6LNxkhw5kzUgCP
CP+rd6SQUlncU1rYaMUN2ftte1DDFS3SESXSWt589RTuYbrTTvLkldG2M0zPo2kI
/cKYsT4ap0dg1KpytHLoOi+CRp9uXLHY26kU4oJxbJ33JqSX39PHaSuJNUOBPqGy
H1Be5DZbV+VNVuAmmxVaQov0GJkUj5l9cxR+lOcakLnbd3AIAB7I/cQMdVi0H+ry
4R+zI8hHAi77FqbjKbgUi03Y9jg5jFLS2BJdSzjv0ACsad9/kKAOroyPjiIiGYX3
zGBTueDRnUO2j6nrDQlTPQRDlWJ7MFagcRbI//O7NDIfxdSmJdf0LrgPHfhiyEL+
OWILiCRKnZ/A47ohm1a4o4yV+vz6SBdmI9RKt/gFDWyNHtCflHEu+c3aT0ENaNbO
Vpl+4dsdielFNjVCaD2Skdhps3mDpsAuf8IAmS7lYWrZT8g1illPLEQuUpjc9tvo
4vt6hNnfaWfWVF+VI1oTRjn0e3ClWppQSsLz0NJM0e8C0vGRRmFIi3GCZpKWo/56
kMrWrc5AYUwO6UJaF3UCDhTtdqxvWuEE9APOJgXkqsbzQLV9uyH5nk0rQS9FG1oB
eJCLNbkmqFUmIAztB/C99uGoCXlnr8pofVYubFil0Eubo+kC3LVspzQpzt97kTJl
QmAUtsjuRZ1TrfNj4F7/aHh36JhaJSboLhRoRhU0an/MzOd3bSl235jideADdE61
q2lGnB9ga55YQhclxLRq06yf2/Wjgy7Z6/PIZyNT9ZwKQnh+ValFF0MlDceQFHt4
Bt2831DgD7FtqvMzHYn1+8d3SL4qys8PnlVEerw9fhDnsa277EztJ0HOd9ZDffEz
poPaPMhHI3A1d+gWyMi1+cscIBhGqOwEuY0wvU4+yZ54UdGQPnpZ5wV36mIISEg2
VBsFlbvrkLPA23vvCxW9gIbZS1rn5pDGkjZZb2um4BCbvSbMtDgjYz4f1tHdB/g4
Y8R8FXOPNgOLCb+bTfFwjZ3OuKlkXLsQXD5lmLBN7JmhqMnXq3RWuAk0b+aBC+oe
TysPhehQ4Bw5R76Mq0iBQvfn91FqAuiC0X2UNR6NcGEH5XwdYhJdxn3Fdoxx9RFn
7Nt14214NTZZ1wl4fWecLI3otFnSkMCRp5ganQs+9rctUk/ZPlPjZHX3sM4LqbFj
4BDccEQQc2IluxIr3r6rrNfgs+Z5yQx/43WXrBvJoHfZXVS4EOV15dhxg9Ar3B3Q
80lztEjzn85TEK914TWm5dCX84FzC8wZ1cOPUm3pdBngNBwCCemxOJGScwZxwakN
gjjBJWlCThkqgQ9KBd64YNb1ayysELnoSiwlfofWCXBHKdXdUKxJQ53Wc6aEdCn6
5OVKgGkqkdzmZhpXEW9eRKjUXVUlLNMcVhIedAoFNEf7QtBg7reshGHmWWZIKAAx
qyTD3KQWex7tHvOTn6prmCv8bPf6pSKUL1zRVCw2FUTbMOpcGyjJY+Uj/pssVC3N
vtuRfHIc5EWn8cmQq/+yCh/ML/1IFDf8FYY1KXb5JJZuLUQkD1RirT2ztO+zeuil
1YN1pGhspTFO/EJehXV234U7gkreKjrUz1Q6b8PXySYeE07JQIQtUQpMTFz5Ujnv
NAk8FPMXsQPkaKxDfS5CjTuyE2zIjbKGPG7pSqTQUmix5ShKsB+3sb+50/IiumIy
o/uYqoan1nApiPv4Ohn5OBwPd9n3ewflMH9vEf6Uz8XInPm7dZ5L8REXin9Ypb/Z
fnmDAZzw5x1++pasgku+/y+Xz0uQp4IymDavq0SZWbJJ72TQDPbEl6sXKFTeEEiP
zt/GqQJbJ78/WXReX4IhYhYGna2EYlRRIoWcOCwNuGnON4hrDAn6FeEJ1SuNJZNF
+mYyzJo+PV0jtccRlEEAX2xXlCOZVjP4zRjOt1FHowZ6AsKysjwKSURgl2n0gzGK
GiVhPjUZJu7u8eOL0LmGNxoW8zip5NzTMYSHtrkE/dfsh1W/+ro7Wz9+NnsznCCu
p3/pSi0u9T+8qPIVgXiKRFyk+wl9LkYnPdhOJoVIyQR72nR/Hhq4CThRFaA6d0uu
ZxhvCYkDxzeJgUu+05NxopcSk245xfM7ch0IQ5VlAhtBXTbuXTrh0t8cl0Jpk+XI
qOkMzh56y1Y5UdbAJewVsglEHN4EhAPY+H2bEcX52/NQRMmAJwol+IaFLz1NzNW2
M3JpxvCTzZyR/Yrhdxv2eVQJ9JrhbA52AUZIrTZ4Ewvl88Q1Oyq8ddZBH95vl1o7
WyjN8UUth7IzbnDe75gsD8aIB8J8XtlRRrKmYlA49+MKgQypePyPeFoxFRA8F0Ep
8E9k4C4gFqliUIFtyHCCbtgPZ+LE8PjE+WHGQLGMvx3hfKOf7QkTLrG1QDNwi/wd
Z7FZzG6o0ZsHYG2QVdK7SQLcS4/OgnZuG57hfn6g67/w6+pqpuUIbVMOVtU7qL0E
xJwI6SbGiFEoUVPZ1yuUIFVBLEwcPrhEQa24HJtHG34u4Jbcw1p+hU//ShFBRaMr
12LuzuuB66siMQdmIFbc+ugF6uljHHtv1xCrkXEC1hrVwpJzNvVW9dmoNg9cv0SI
7nu5NUqDm+WnvI4nJ0g0mMg1NVqq+tvMTZR6dE7fZn3V4K0FSB5Gk6XdqZCYCCBF
9oqYZkZCHK1/ngZTjqJCqE86w/MMgt+Vy7OsBxVneBs92XMCufspmzM8pICEJK1r
12R/KxQ4gfDng/RX26nCB9bhsVunEQTNJMqTz/CwFNeQ3T2dTfqx7REBn7zp0+QL
fneg/Dnth7MShs5WWxyvYXsENZicTO7bvqvjXg1sD3UO5T12Sxc/RcV5Bk8BPxoC
x7/guTteJK9VcfjaKFoIRyXJcL8HZmzHwiaSaCIkGYthHTLJBTox6oW1Tv/wt0hn
H58QMvW1G/ezHbf1/2h2Xn5EwScevuJ8C7FyDiQgZNunouteki4TX3512E+5rorw
fORHC3ieO3l3GVOmWQ/rWzb2ROy02Dor2WhISfMtcjX/8NqeZ5TQC7u/IIB8khEB
wqlHeTwFsJDMZJw8fOW3Uce8rLh170WTJWoH3/Lma0Okd3lU8lvUlvUkdQjZG9KP
gQ2S9L+wASOrxi4lOCDyJ6nSf/uomCYOiH9LAvLBAt+7cjHHEsGb5BsQN9L/GGTH
1HDXx5mptdMzZX7y5TcVLOSMyxCAKY9GhqJu2Juv9geti525JPWkuJ4eVsyPX7K1
J7o0XJzyD14KIIzCIDwiT3O3Cnjw7wET5w11QLxrY9pWrMAW/JE6CBmW2mc4OgMg
9pz0cmHCMUoqahqUqmkhvgOMYFjkcdG3s6EKu5fdmAyrNWhcw3DhxM7At5CtjTLo
4F7WhW4zM8qHuI2ZcseFfpQcF92djYqcH0cndLpdTgjrVvri9Jn6dwtRP8V3vdZS
7jbUHM3fyjKSTrleiaFvVc/VLwYlWYMKr7x+vV9wOIhSnhCB9on8INPbT+ZBevYP
/F19vuTBbI6EGZxux0fGlR4i5rUpvTnAZ0zBRaW3X5w0eVr9VjGBjAsjGTlPNEkJ
FUiaJ6tVBDPwxAQHYyOMGGve59PaUlcK95Yb2nQAs6Z6KmnjgtcTHtZZdQk3EYnp
RuyVCp5LBvQlVmvA2d1fOWqG7kL0JQi56hrc3EdQjXmCtVKTgW0Q36u+h/dLLxcq
Ex2PzXoYSWrA814pNclFW6dK4TU+1xrlw1rrkqpXQ7Yj1dUqgHx3qLYB319kLRWB
Q2MZEN78490UDFsvQFPNVHd7ZLrXWdxxXGdu3Rb3mRwTXAfRGFTId/D191iTgwG2
nAdgT1xYxMU8uLt4Liv5g9SxX+AueGbPIlkaARlLmVXZcstQMPJBI0eTM4vSTfCN
DslG9/U8aHmOMwmxEiV6N614sS1d9Bya/I89bZh5WBsTszj0HrcRWHMjs9mwIE3L
KK76Z4vijJHQ83P9TSejzfBPsgPKOfg+DdxKPg/BqOMRPG24DG7yQKsmnoZPhnUN
NG6hhtwRa6klMz5vubLDJKoRXyA/YYXVCsGQ2ycLgcTndm0cHdY8jo9ZGCUkAxZZ
866AqrdpxumllzhnI11A/mXhrCdBOJ7BytmR9ohqF45AjjtBKWRiEThDJ2O+/ruW
B4cX8bAmnUPZbqK24G+YeOkxnWMEl+Qj5U7g5o8i03dEWuxyhOlTwuT1pGMjKI9y
7rFdhplTyfSPebkqQmGgJes+ZjWxkpDIQwWjz8Ftl+NVVCkZla0P9oj+m04UWHnm
M6XtwPpU1Wf4GfNGIBCHh/zRMgzg6Xnkl3om+Sb+zEVzPMT8qpjPV/TTdV51YEyz
nuOoFZUpDnh0LvCKh+ljFxDurPGvdZ2OH32gdKkDIvnwYPaymamNIF9SegsLL7ee
5hl5/AcaGZWJmnCpDD0jtBc2S1+F3slZzzZsHwp8kXlWhDY6JHpRVHTdY8mR75fE
739j8qaDYBDDsADa7F0ZWXtI0r0gEm9HEFFJmCXvqZKXS862dKSniqS93d9cSEwr
AUIydEHFOZ82VRDtv3HuTUdr8fKrlot12MY1dVcbqhgtE7evGUqNGkAtx4tdv7hq
/RNanjQXaezX/l6l02HjAjaYX7se5mHwBTPBmPvFZ6kSlwOpcmUVpdBnDYs1q8wv
HLIIt8udd3HriXBSGll2S20xkjWEi/4S3hnLGKhul/64fhjQh1HPlqEemPN2z+Zl
0UgrpTMvm4WgAT9JVjnwNHRztqyExrgwNzf+MriVxlFpnNRrM/DhFeSO/q1EoR7p
gxTJU90sqbDL9WRyRQXRCHaMiXmzniUxeOdbcs5rezl3o7wO3HrzVw7tTv8hhWeR
Khwj9fRKubW3NsxZp37ueW9P1thwH8FiPB+OzVGuaFaKLVQ1Cg+lL9beuK+NNwYQ
lJmUjbyGybc9VZ1sDXQvI5PU/p0L+lGhaTUnDHGhsxaEohIYIX5Za4yX153Ejhsi
2pEz9635nAfhULOMGDdQLNgSlOsBCHAtnxlvgJVtKuv9eDKFGD52FPkruWq4IT0q
IWuiuOAvgFmI97huVAwtsDvEKnm/9GrBHT3YJs+4PbWZP2EEg5z4aNeMDREfgqQK
Et3dd5sPGD4C2ZqB3qkQXTfDSn/CLfHciOuNt4D+Knn17QgnvqO7qwG7Gq5BPjJC
qyUa8agf6rw9yTrfodmaIuIWuUgWuTPBHkSjQQGILKbIjdbnxb3FdHg7zMkpcLLZ
6UPFkvxm6vZvefNz5Kd+M6HYIXkljixZxOTNx43Km3bFEhrZsq9NArxefck0noMX
8ZmPApJeddGbauDnOi+U+CaPzOn6cra35Bq/FKpB9aQTtgXEw2RP4DWb1YviH1Z7
jP30mbqquynHCV9+Fz7pGoZuMuwKPQhxcpihqtdYif+NIgKKAjuKHbfHdXnr7Jwf
dKUjlQjgnSVl0gr87M/1tR4SdXfdQOdIqX0L16/d6h5oyHCbraSpjTgNZ5LBL+2n
4S5gpHB4teq68M+xbERsa4p31WpnR6muUKHfLWNVaTDtV3aeXKC489+rvqWlwHYs
lA3BKHALI9gzAcfzzMPhpH/Z8MdNdHfdFR8FDa+jFRJ+RKA/L/acxIYl6XyFp+ns
IaXXJnPY/udnErVsBHs+8foaMaUnT89WOBjRShT+uKBbGU1f53aJ3b1LV/dXc30f
v0rmqDNnzM9gS/Jwpd4f8WNsRBcQgQ8PFUB1gFaH/ZzGrvsWIWMdLIxxr5yADrV5
rAo0ktWnUvabSCqXL/FpS5G+K1kuoEcBbxl/iXlsA/mOXkUVPg/TFpYKdf4FtrX5
uyP1Ctges+d/hk/02zBa04zjmIZ9iwCi+qEP84W8XpaAM7YFWDmEaO76Ga7gCuS8
+XMcRWiW6f/j8J/EhgeH2N3C52r8c2SkOljtTG2874tuflwP7hpDgfJxkWLSyCRm
Whslz9cIw1Vk996PAwdmjJuXN1yZKk80UjiSVRdTxq5N/9H3NkXHnDcTSCcgh4/9
rblmHZPpt+gHhc1XK1NoEC1TwAUylVBRysW03500Zh77plZt4gOKXziLSSl8y/A8
+8Us3Www03po2qx+wmr0v7kk2dNck/Xgfod4Mq8qC4uk+aZ0ae/5KsVJborthpKM
peqmB91HiCR59bbd2lSUE6Kd1Yyu6dtXGeC9DDebI2nAyrGNP2juuV5T+NXaUTkp
C2Jkf5+CXZAXenu6vuc7+0d6aHh+h/sPgVxHL0aaLtAb4yFBGmD+ACW8DSMq++J+
lqf/5nXn2oxKBRdFG+GGXeNAh1Jq786S775psJ7ClHekhslhoJeA/BA3bF6vsWQv
/lz4BVNQp37xnqVfj6pxyKg+VwCMdia6DpNzfp92kLNNe4iHmdmNpjzkGxOXZAgM
FwXSRukgxbNiT3JHjSxd1aXIsn3ajzpL8m+Ju4h+UyFWa31+Bm3henfwE0VZ9HR3
MScaFqGXzLft1Xmq9kLNj3wyexrV1TXb95XKU4fSeBqioVT8oy5ndGPbawflLyIN
gP8HaKkWl59NEC4G78QzhUwHkqZpeAfziipFKu+Lb+9853w7R0t5cKv6ilnCoGBQ
q2l5rkKVqJ/zeo9qeSQvGtYrH7PWGdOTTNqjjKuuwpR6aAdkPMi3lS7qk8Bip5Rv
nqnJubDhaZFmlvXIpw5eOfDVrRhvXExQcGtuLZx3tiA0jFEwXp/IuMhtZ8zjJQQg
LbKo00eeqQuhRx4W+OkKYQ4erWckFWTRVGx0i0xK7tssyFMbM/nKXhrsIYK+GOs+
tgD3wtn8/T6UodtePSTmBgD/WSBHf7UKuuR9aOYWySuqcjlhuR2kmypbQ0eKaBQ2
46Ub9UXr2lFeRuZ07FrH4o5Bw+tQUrw4XJIAlcOmp59UiAu7ei7hKAQOyrAnkX+x
G+FlEewrM3xwy180Vi8/giCjbYn1W3in5c/Iwr90+4Pq1a4zJeuVoixXO4R9APwW
vSFHeZKdVCJA+b9pqGomToyL1Rz35tgdV4Okl6HpYQ99fcg6haollDoDhXgfZGNo
V65IwXzjtVyXbAyMb1mnGhNTBCo2qz5khWAntpD4B5Sl/gf9cxf+h9Z3ayuL0rLF
66uZA6ygmjj8z/RL0MIre8zabGigHOWoVNd94P/alm+rp093RWbNLfmimvuQo85t
0xpD/bLcBuS+di0WvVObc3VyWxeRZ2eajqa+Eqop/cSiqjfCzJY1Hfm1D946M/GS
zw/SbDfuVWRbK+mt5byoO43W1un19g2ZHYYkZVsiuIKm5WZBMIMRwsyUYysp561B
bUS13HRX8YXiTWud02g6DSFJt73f3uFFWlVP0xhP4O0qobeJpT7l567iyDyeOrd5
LuZsDPcfBofZYOIiccfFDdxHYBOBzSHursxK2v/2JUVNRGd7451R53cLQ/fAE854
KilrcycGexjorBdAu7/67GXcyuli/Bd/zrjoDOcD8OYd8LH5GSOPImet5VSsoZ5V
t7jpLUcq0UysYWyxX89qGWdoVeELD160sMaGw40R+KGQNQCXf+2HlPnQV6+v8Qy8
ltn4ptcoigZAyF5mOdVHZpfENxXtLSt0NZfdlc0Y/rqvMc0SAq+eSIt+1dJakoPV
8a7aVasPqUXWhRfGRIO84Cbxgg6mKdxQ3K1q2OHnHR7gvAzlUwFWkpaDiDs48JyH
4atgmYctJ/3cBi4jDwwapcH4BhRjnyF1M0FSmgHEqsHwdAwN3ih1VuyvU4/hPI4y
m/vJJvk0XZxDV/eUdzgAwVOsN2TgEXQAn0ZC70y2Z+GXXpE7+g8AQo9gg42uDQU7
V+jcd96VPm4AaRjZk6trjU+SK6OqlvPIXW51yIfwX4QipsOKOl1PyoC6QrinTRXV
2wQ3n97Y3v7ZWG7iL58WAmGe0uJjP0bEMeP1xZLP1615Emtg9lDCyfAn6/jnuHal
oSA0wH4PiG8yyzskbuYVg/zWoaWvJcaZqgM9GpqZr0OQ2lCPGQZzKyIrVylCinuu
Q8/aIYnI4MpX3NKmAhNdKa+X+5WnYqZv22lcF9r/oAONmSZFtM/61592O/cdL/t2
PFWELp4aMjB2JWZg3r9CkPB/Ng64V2lDTGe4VPJ+VcAxRlpkHRAs+CA/sxpD9ppn
n5XVBFVaMD5nW5lRMqgu5YCrEEZSZr7eM4z5K6cpPpHww2trnqmoSjzIFjG2M7Xl
cwa1s/LmFWsTOb3xcsaAZytQlUfaQIPg+t4VUr4f+WGoQvqxDRxVmLhXJRQVb8MC
HFq1vYVYeA68wyFPoS8t0Fe0thc691ozOHOlAEmE/7qG38sDQ5jk9V97b8lg2XZ4
Fsne27vAexswZ603WZa9LWNPT+vWmWmmMXhLhL+FXQZCEyGHjf66ykkZN5PeGMKF
AUVVcm53lFOGA6h3+nyji/o5QwGgBpO75DR13phX4zSi9Mu/0bLJpm6/nWAdc9TN
9d0SqO5O2njHiRczC3FVjdfIU6rJxc1ylbNqNIlz8B4qKQs+6EcoBTLQ5vT1knwR
7Yn8HTfcYEPYzpmxXf1O5TwvM6hAM5dfEWCE1hKc7/c+GCNbsQfI6oeLm3EeSMeS
stBojje6eFh6OFQ40RwVzbFJpT99WXB9AbIBzzdKcFQq1LYxlc2n7ZPtANsoYNAS
HOVhsyw3sxf/oosdMCuwECtfOqtvA7fqPq6vwJZTxSc949eYqfRcZkwIlSnkrOGS
etjpE6NEb7rTwrtf7T9IfqFfjW/kHSz73vMXuOZgVVW+qQdNkiFhKBZJ236p6Kw3
uOHUklIT/KxgIdfLWwGWkZ/s5RRsC9h8hPcOh9REHY/ztf8w/UCeyXfOJq2Cb691
WATO7XUxqimE5iTZuKE8f1ZVx7s8oURLIxWbL1G3NBguk5KWuWU22zAR32o5jYoD
AEa/ZeavIlUuganBmUDWxkPglR7QBDlhFXD9diQ5RLEo78E4OlJ37OA8/IgnB96O
EoXu1KWaBSM1bvRkI1GZ17abbv1tquV2EwdBodSVZJwt93EMQydJC+EpzrtsiM9B
QBiYYZdNnxTU0xoXMBLjJMYbysMw3SAo2egP0+Xk4GCtAvDNhYllDVnC3cUblhft
epYDZFx+wAUzpG6Gws0qP0grbLOwJyZqUttaq9tnG/u+A3VhmUMDGJCC1jFIA8K5
gvdGzR31soSVAWybhhpjmzFNvKJlULsKYLrJM/mj6Xr/8dtCmh9mMa7gET7FZT/k
IvnN6ffNwG8lUSUsH6zqK7Kdahyu0ZwZCa2mCkfa9OmBXMXbRzCodw4E1A90i/WB
YDTpwm+aDWRhLkasXy/C2p+iOc79KZ0keRNFcW4kKPugT33Fnfz0xgdT3gAIvhpH
UjIuoJk4ih3uQFFAGgnwMSSs6Y8xf95Qael+drDAxMT1AGb/KtBfDBhKYoRrTWYK
axN5+YNgcU+dqTRTUdS1LQhrOzOTQNOcxOryinN5Ob6whkpGFkxksWiWgL2Wh/8/
ZJivc7ejEugifdx5l8Cql1/aSEmraazwz6A5nZzWkGxxZYYWgt6/igR5A9JeDXmF
Wz63xaFUJdohmzOmZoomg/nshLDDpDMAEYAta1YN1yV31gh5leb71gpDsWV9AvsU
+ZysIegjwQM1oOVVH27AdeTF/TM2niB0eWnhPHxidX5Laq2vawREueXLt6OPVd3a
dSj0bglnubTd7OUoNoqFH/efpFqLbsHd5uubjr3Sfy/DWPOq+hIyvaa8c9+ZuGmT
3SZuH8CY6zm/uGZxYeKOltwCEtldZLt99SY9idL5tpSv81Wc5oJUkHF4TsUt5ZDM
fA95jlfQMcJmUi9+7+xGa/LT5oEQKPOsbfROTh0GEGGSlIngsGwU/C8EeKimwTOz
PhN566JF6kRmqmaaRM3zFhjblAyOO40+AQqtf+NBFgH0220zptvAt6nt5XFr1HV1
yUjK+3dKrrJpOXT6w1spAzvXRHfOBiC+Ncceg+UMmUg9k2Ge1K3uWMiB7xuM13mr
5c0FsHr/6xoCD7AQVi8fQ9U6MvFNruS9VgTOEhga344m+QwB8GJ9Bw14M16phz2L
XOezNvMDWfTG8B8teY49/oqjeZSAEH3YlBAqJetEeiV3osviskI0oc5/utULpFiD
DhD/zM+ROmoVj9UwsIUbQjSAjzLWhVJDsAuYPPg/jpRi/bm3Kll+a5DtVrrs1xjN
eP7FrisqcoZNxgQeXaQEHljN8TPPhX/pbCZza3ewS8jLbOqbfR40iKAsrBBV5I2s
AixjarRjWFxReWzVn6mf3hgIQh+ADHqlppDfD/n/Zju/yEg/rTBZCKsRZEU+Q1NF
+u9U1gt/+bRUuyoPaREvxdA65KXZULYwIQyrebwj8Vs6zyma0ZtEzAFlQy+Nc/9W
pe4zdoQOjPiN/KMQIWthxGq4shamvp/UDd1RrcXVTn2OK+wwlmSgW5jGQj7mfyI9
fvxUWDa7NMk2RWDjOjK49Lw8wETLbjImIhNsitDo1Ch6ZNpEuXkC2515hA/G38cF
ZeAD9tROSeRQpVsc3cVG6A6+BMqR3roJHoI6pIEdOUZySvEnJYLdlZBmCBmCFcRV
G1/XCBonVHFhVpG9W+IP+n0K50a7YX/c0wEddBknzpbn1eC7K8204QyNivz6VhGG
XgLq4iMeQ/i8VlYjsqxolc2i7W+ICbbJNUKOwbJySDfDYWCPXgwphX0HLeWCJefh
sLYW9q9Ht+7Dk9oAhKUeUmYNDmsvJt6K7rOjwdyp52Pj6xTkzHIaE26K9hPZk5pF
HZsZ6QLbW5mOCq0VfahfLce06wix1cNsoCVvCQmDWrq8IjlDLQlNeq/mJDxI1iJm
dU9d/YZhuakb0+rlG8GOlfJlZNZodMUoaxJpMLsKMT6fnWnODhB0yJuF4HICSLl6
YkqDr99GZ4n5i5wv01oWwVdBbAE80VGdBK7eRIWb9+Q+qboYtlBxwj957V2nI6nC
GbL5TBrLM+fSRKMJ7mWiHkdQIkwZ8i2fWL6mHBy3grsgonz6j7nGyWQJbWWy+z/x
TVs7+1Af9ccVf4rToFxq5kmfKcPwdxlwUjcqlt3lCRrLzsZG5H68JbE5RV+OliwO
0bl4gC56d4F/qx5SNaM2pmwhy/qCY9ZqrMMLEW7m2dtPZ3F7uJijTUuAsuuvV/IQ
etFUoqsq4nEMjT0lnMrkyLxeiFrAOv9A/GQwWRSI+ihqj+dH5PKnCc4NTOHhQLsh
lasP6431ahQF6e6WSZkmbPWvOueRdBIRa85JrESuYtTGPmIrNKmSKBTDYfVYWgaQ
f11X4Dr38dFwgV1asnQuaZuPWmjlPTQxIyBSCf0yazgjjGPNZEN5y2ZtA5eEREhR
1h1QwTrFpnvZIj0FequZqj2AALNG/UDZ6bhhi+/vaPMQK4RxPRd4rvG5/KZ74DGO
MXGuea/ZNOLGScmxP+9HQGMwhca+8aBdDV5Nm5YppUZHjlalt64VIUBmxIRIgJ+b
GmG9tigEVBouuzV0cvqyIm0PH2Q9axY4LlXQhWHTBPx8lkDBB6Fz4EXLYCz5uf/x
K7p+QWfHsAEPXDPJGyzCInRUZ/yuQIqI7QHudEYIxG/lPTu3bFmfbejOOPSluTmZ
IF90IogHghMjq+oD591yW3TZzSO0i8aU7Ftef3Au2eE/Uqf1CpBYoaa2f32o5mRi
G9Te72JOYJD01OKgSoGBFEQzYoDVu7fFkGveMmtM6dJ6V5lDAMsn6UZ07bkpvONT
l0fCn55SgASitVUbi2DaiQpJn+Mnrh6+Ykl2Cz/90io7xarzht84TI/LmMOGWqbh
qQQDCq1/rCRSnpRoFOGwJqqNiqZUdLB7UoPQWJ4586IA8usIL7E5OJi1hE0REmil
Ma/DjHduf07EulZMjdfPlB2uI1ATwz3hYnZH1p2q9SYSGWXheXLquwggBjnb97A7
iFYFGGr6RGLHRMU/a4vf1C4bwxn7Z/GrRQoLCW4QDXSLGsGckfw0WLxQUx/Qu7V9
x/Sd4/Nb2WkjHhwf0cedtMaSuy4IXLhoHu8I7LNQBLXcQXPs1H50kJKtUIYuT8OR
xu38EtAHWA6xWchbQxa+gca3Jp5Zw/HiTFw5uUcDkgkB3qSdFpTWfIkbnJ5Bq3x/
Quy8dZbib2vVKeBYtG/jH3+KcxQHTIfmlpJet981eblLrykAY2EeQxwKZYHu1NxE
5TJP/fbfTcsjtq3YzUz3Iamp3j4EWPqyGqHjZrIDU/YP452WfHbmJ4Rk0tnHbp/w
DOvIsdvvnjmeQNcsh9PNdytRkj/9IyE5jTscyYI5GEDP5/EjYxwV0ZWKE7JxxkML
YploMQq/tdN/ytkiY6JHfCDDM/Ig1BclxYTuz3guErxgqsdCsDA5iW8+Hv/PmGMa
y4GSGqbRWdOMfkUIyv5q+1pJqusiLWbVmE3IhrEPjj7FLbWRpdSikFUHXIxqIHQ3
ptkGxsc7uPmagaXm0oLTB7rFe4YcAYVJT5xeSEWy0+gElV6YdMIO89/iphg2px4G
WIgPfk321IhAWnKmRWPgdIYlUk7lUPD76fuoHJUco8dq+3RKayu6Aqq2umWYP1/v
r3TX2q8plfR1tUGkbWAfIFFx0irng/m0vxNLUYd5x5EYNbMwfl9cQAKO4XHmcjpf
8hqHLZvMnAbno0MOjvo5mxNev5NFbCUPHyiF/9AXmaXIrrPnyg44vH6ApfH1zIGF
sKrF279UR/AJuZVe/81kLCWhJ9PPF6mDWwKBpXLR079Rbc5t76Z8eLI6oS4GGb6+
Zp+rBEGNfAkczD5SwTH78r5asdNg6F7+U4sSNMX3ySTOPH+rsLD93EuO4F4YjusU
bdg+t6/Q/Je0h4McJfgymZNXL/Hzrg1k+VPuKWh4ZVdX45iOKWeeNQZ8T24dQx7f
ZDFUVccogHEAsFPm8PQk5OCgUj01oBX9Mm66vpJEG58jPj+VfMgzz6YPioERmtoD
oB/GMr0T0+FHLi1St2YYBMlrZCrDTsbuucAEa7I7u0BmcoYUuAjwBQojKzpe4sp3
C1s/+MHAoXHJuh0O4XQsqfLLk05NvPzypN/mhjEZWTyc/yoEtbgf/IMvjKCMLNld
/czuQ6PRyQtO8x/bvsjTrlpZYJcPGewaIu7j0LAbl3KUq7fbhLoQRH720gVyZOmD
wI0UP5nT1bfMlpNJDx6oYePyHmh8/FXbUeBCJv9kwIsyrXKMmzP7d5ChJ903Nwdc
XYiSbqzXuOnG+lreTbzdC16pAC+FgVrUhqzPKLHYcnwLnyX3l8DNM+6hf+VSBW2g
9dStMHjvuF3BGjF6ZSm6SIv6ycbkZ3dliJLdJvyhdREh/UkBuyCUulKu/1cmy+Iy
hICd55/xH1IE+UyHz95AFbWyl1/Tf9sT2PdyRzhQ/NYsQkHacAgBG59TqUh/GwSL
autR0EL3ahCoH0XbbpBFTAT3cpDbOaKPmf8GZ9LKbJjZxbbwunUzO5U8Ntu8a9Yt
BAGSpRJwCcrOz2AnahAEObBL1NxQYrUN/KHf9xhHhdTJoewImNx/3W3tsiHAmsOf
Xu76bgDbWn0l57BoA/yU5x3+XETYv+s6tXSq87swdqyNlr4Gb3ba8XfrpAIfa7Ll
CUMi2CEAAwGZ5L2DcqnFkDpO3X3Fy+8f53fRDoEpd5BZGD1oPqwsoBuCQg62zjFJ
hz7ASp4UK4C14TaAnPP6o01Jj8JWi+rSVgwQEMHI2gi2XpWVNjcnS0hJ7K22CDxR
N7/lHbgFUCEAHM13vySn49DGIEwj3AIN7oJ0I4pYPjN3OIUeA7nIREjvqfuZ7Z+N
tctQE5m2B5HJpDiCpGCzhVHcFiXtlrMyi5J30FmAjrEbyPAf91ITgrFJpXadsK8A
hkoyKYAcqOiMILxegNXJlGCCQA2ENowFLegNkqQew+0I2hFrJyMdK5Vx3Vc4fEVX
zKOtQjTLMV2POW/m+70y/waS555+g31Hb2CPpTciMs2bPLu308i1O+nvXREMRgMF
ouoopx9V3XkbIi6RiZ3ikZvBFCrWeP96isGRezrjzhoeMo3lDADmC6skvQaGThG+
gU5ZVFNJCb/a0NlSZAhzC+V3v2KMHSn6awVC5AvDEt2Cu7un8iLMExNYg6nCHl1J
lNqraHSLUfNecS5uvIjMzFdqjE4S3K+u8ylCSFv7mSOxtU2Sx0LEM53POSE6H7eI
wFgI0E3L8XwIEhIAyWCE0HV7AHplrZzm80QI9uRjQ1rdpTo928aRARqoqMItDTbW
UU+/mCPmGs2i4whdFYgt4AUbxosY792HHjC2kRr5YRjAYFhsp5j5dpD/rCgDqcTN
v4ihCznGKwCpx/tJO3tr0uwXieRIDlyJyoYPBxpEfGnzBzOKqJLASeN5+++SM0Da
Rzk3VRX89msbS8c2+BVEhFUFg4vOECBvXVA+ilE3UupBTZ5dftxb/zJwEmfUBQZQ
mEIktplhKZBTj6TGO/LqzoPU/iC+pSnydSg6Q3UolW4mXWJBhY/jhsCeLMxiNKS3
rho/wKvLMn9YDjXtz0Ne01NHXtGtYOMEkRY1WmRIJaqFYS+BEE2pK9SNknUv9h/R
+NCjsQYvTjJSa/+uvRPNrcGFEhHUUPCnthgfBOvSL1C/8XNEJnE3sOAo620sTQdW
TSjI42brrptK8reYl1DebLfDImlTMPP3z9JU9VPWQ6qX6xdzWWYjIph9MrNkS0qP
TFs3tH9Eq7edr/18kNZgghTVf3dSzOUBUOsm/wsM6oE/N5xd+9cNro3Qvr9zDXLm
VFmOiEEBF4wTRXYlRpSp6465NHqrpEC/1FgByFs/YQLmOSudZtxzT+cte3nkCo3q
2dONlcGVSQH6DyQGyvsjP+BEENEiVauNTT/8LRjBXNs+Lt5ik38AfjHwYZ402jCs
yiQ8u4LStqVjf4l1fym4VZT/93g/teiJZVQsaiUEnGmiKfVJBv5n2ZNevKePaooo
imLn9I25FcQhzNXXvbfcgn9PmEQKLFqAxcsJJHKVjKqQyYbYLmoDfUdiI88CRr0a
alShyR9acvR5SWVeiLL79uSBaXtkjXnj+/xoW66QmADQXPy9AvbFx7WTFEBoesKc
wO+Hz7l1f5pQhVjsvscnwst9tZQ1tm3yFuEWPnCNQKoT3uzMNBviVeV41reejPiu
OEJadaSUH9II0IEpT3Gv4i/SeriHe/JxV7XeoAlX9RnI5ihl+nSuiO1BRnwBnkdy
F7lt0Mep3nCufLVh4fhYm1geg/h4FUzpHej8qKUIlTGBdH+WEMs+R8HAKdtO2BfU
XXQn99b3CtTMDlKsw7MYsx8sdi+C2rahj1RmlRvtfNQhRJOci8xBL4u6BpH6+RGf
bGOuQnIPoN7NvRJsJourELYts1UzFkeZyX5C/ON5DCau9jNsySVP6W1E5RYyRRFc
WKJ9ABh9VtPiZAY9olrJGHfR7ms/Uvm6JsCJANu7aoIOy5fBLMh6ZApDoVgydYIe
HrBJKHwbosB/0W1/+BLX8obKVfH6+hTbU/s8mkyvyKYF3nu49fAsZs2iLJEjOzsv
4oggLQRfZ9rzBlWDVOzIPTPFouJPCWSoUziufwcI1Bwaab7tSjYhBEcx8TSGAf2S
8KmGJc8KyI8H2HE/zQicRKTPQzLr3DwFko1AU3absmaij20NK8r9waIhlaQsmmay
Juie1YvriJTBvoJA2FbTXy7qagaLHL3ibxU/gDyT8zM+N01/eHVnyBrcLwMKHe4U
YP5d2H6gVhVcX8NMNP5FITB+tfiM1palT46sev/rk0yqxw480YqIF9pNFmGcM2Gz
PXD5Ttlf6tpSfG4XwjJX1dHSDzwkZ4t7ha2jlbXTFO/one6OrB2+Hd8DJUsWm1sN
ptdPGYc4Ul6qFmmQCG9pDVoNwLMkqijxLWoV23j4QHSVMBlU/T5qRJzG3oxdkUJB
nit9Z1RcruoCkCXT5rOs00IQ2voHZunAXLP4GRmoDyupMz1pDco7+wrc2jyovkSP
WlcSZWbaV5DG4gJ3Ghs0cI0eYP2PS2VMD/xqhkXy98QnT9rYON17GfQSbcWqLpZP
Z0m5rvYcyDWBVNEuw1mUmE5UxnBj/V+6CvC9pCez6e0zSIj3Yyy3tetKBV7+c29O
ZNdq74Z6HTh6BnhtMoV9oEUZCmDw3alWiqgO39RcdbK7ZvoOZNK/tnWzlaWzfoNG
lcscYW3I5o4VV6mkRisaw2c11TjJiuKTiDk5h6D6qJUA1I03IXb6TTC2OHR8LMxr
ciMC4BVU+8ymbRkeoQH+geX91sd6m8PP42nrSOYNoLzi6WMe9Yh0JaMluujbRDRN
7jHTJjdt68Se+1LTaAF9bv3TramAOE2NzNa535vQBdRp9g+6vn8l0iSyqE6aNurW
Y7086DtfToDhnCHYgZ/7YCXCywJo9GiCH2CyBHrOeM7CTycXc/9RwQtYAGobpVq9
pHoTqFx1v2jR3Qsc5jj8RLE8PSdNpPe1oyo77xEHFY4+KhfPPW8xP/WJM+Irdooq
SjdBboNarHvW/ilftnb85JpsrKIpYs0oBMtuOG6yxGVByfSBZ6/8vH3SSfckmTxJ
fMrg52ifJsA9mxS+HcpWYs5rkKQ8vSIMeoyQD/kBxu9Ys0QaNk5xHdOSBUQwiiac
nWEvN9/Uv2vvhtirV1Q74Dj8TFwnV2lktMdpnnN2AN6fuFlY9l1X1zqb9nhhtEhd
Tf0us0hr3rVtmlDe5nsZZuECkJoXsUTV6Nfc2vQ1y9xbcoqLVXolQ1HmhNgz3jVS
qdAGohnN1rArmsZBHf6K4isZDWyw2QJ0OaAHAqNA9Z2W6ArlFgNFQaviPR7zovBY
drmVV1L/9TmN+SyXezyxCfOgf+pp6D670cD+6HmXb2yzL7j3zPXkjGb9MLeiD9JN
zVxMRVUXmjnVCu3dpapYCjNm79C36MBEcRMJDBlxhQpaAZdq97Rgiic4Yn0Fxg++
n3lleM7hvq3qWVo7xiecxwv6BIZ4uQZDDgXpeeAzlbPKhCIjNIIH/qakgauosFo4
0EYsC3TxGD+zIMT43K8Oj5i+7/wPNJhYu2ZfYLccXwg9fNNA8liUtjNcF4U4pvZb
4ku2daXmX2QunezD5HRKqVOD3CfAZ280W8LOZR8ryGc9WidUbRM5Bgneo4v1fmaD
uv+t0Y2MFPLaiCBP17RPgnQQrrMuZ7iLsb31dDdZtc7UXO0xDy4BtYRjQ1ByO9BI
FL8hPySCizHgX75sDrVLdggqg0F1V/J87HTPlmSY0aVuE4x4+6U+06PA4SLRT0Jl
U2AzcBD4HrtGFp97SO+uHw3ubTVUAQT7XfmpHKSG/qPtXChy2iIwtaJNefNgEjb+
dmd/Zsy4iD7ZF94B8bJMCwX9lCfbhK373uztF7V9MPQqvnyv95Ik27aejUWv5ide
nC/2hCMmd81LuHmNl086s/kH53Hf40NZZ6khKFvU/7kYGraN+ehZRvrWmRo8d4yM
cYQGUdDZnsYbA1N95tGdMIGry63GbU8KlzACVndPeeVpiJJ91Mw3yLEa57CCYbat
b6nB60Fw0TUuLgfhFuksrAXZIDybvALjwa7qJPZXS81l4IIChq+4SYJYLhEzZnxc
WwemHRxMiMonuhUZYf7GUG+CFc/7FJjTD0tkEqWur7lhNU3iERKaAn6XowzWYhMC
nwZQ3JH7h8VesJl6yC5RTOO3msOtp/HI0RYW70Jc8qdxWWaVNu9uBh7IoayK/82x
giG5+8ul69w+Kx7Lafjdv464uPEXTwqP1iT2PMMFwz0liDM4mMXRatXevs3d3RuY
zEFXY4PckjPa+wIuNTq+pKiR3y8YBFtpRVtrMkc3/yJc9T7XK1sifwbqCkhXvKd7
oy1nxiiMmvfMy0IdvnPVxSkDSuKy5ZjgWpIwWcaMbUuaxiFF3X0lRi/HEkSYjPCf
azu17UYAzs6STVDsWvahMz39Q2kzF9mG6fArhhYlXNmj4CSubPYyCwxOipe1KumF
+ZG+K9tcBFPEPRjOZfWB89WIGqPaLZNA0nuIc7nE2Kfg1xY71+hRZ1rozWOYErhE
pBR8QxwyvwmQtt2Qr2H+A62mLdq2xZTgSKAg5mfLAKo9QxReQAUniwycNBwg8WVg
DTx1zVYIu3Re5K5yVPW0LPMTZGwOW7VLkAE0a82OyNpfdHG1Khu/95P6FlboH+sP
CgS5a6BVfjj82R0T9oKmbDpl2C9irLsBe9qss5zizecvHljuTlpsjoIG9iMJmMbR
raTD09n9Q6lN8KMNiQ1T8Ac54ZUDArGGAHw6gFARuFCmAaABc/I+7dd5Lmn6PpoQ
rap9p/LKObTQTW1o6S8eOWifkwu9nMIhq62JiFe67aAsiHLfmphj6thHJDrOPmfS
ptrXkysPy6PIOzscmf/lMXlQ0nd0ML47RkZBRVhQzRSC6xxdpVqIM16wglJRTRt2
4qmkADmCw2phiFNFYxnDjTswqaqdcGGtBnSXklYkziYe968/ujwIuO8m5dS8qcHG
hyS/lSyZIxDdpEV+Ko3vuDmM69NwgFQarGbnuffW0eLUI61YBHYVSRUCw6ndA89F
9FWzG+1rvwrJPQNLFV19qcuVqT1bKoUf0Ew8g1YFmbz65nvTto1Ms4kIeOSmTy9R
E+wrAZQK6RX2v85Y9u2QnltXTFUdqAgk1MDNNTorVmSa2QaodSJqDli5VFNbiDkA
S8pPtcCuY/eI8wtghQCYIIP72cl7xLbvN1oonwGewcDXfeJ8SnXlHxJABlUqt+Pp
K69riBRXKUACznSagxCZxhjTid9Ss0R08MezV5Nf+sSaVfgmovyQ+vI2gUv7Y5Vc
/FlgU5lBDZ6D9InMAYS8KbeJpk1HKEySUmtIR3EzVG8KboDCVsfg5NCauh1j1Tt3
Cda5nQQMCU5z7unwMH0tGnvmKVoBujAlOvMyIDMpz0NfqDDxWs8XGOs8ozUsyy1S
wx4OH+D8DMvHWKqmV+5PsIzX4atQc8OU5DBjup46G7s3k3Y2XhMF3LZszT2TqKWn
VaDRgNxbbximjFjrYh8U/XDUra+zOkxRMtMUPp3dE+KrynlscfaG4r8qIrv/hj+g
qADFPMOo4B+xgDxFNZ+9NTzJsCqYnTLQzRWFqMUGd9X/WOcN23VWYivlNYZ4bMqS
w81P3ur8UlemcE9H0aUL4bMRQm6I/2PhWzflE7AP9oCtzOvX46qbUBSjHEMc6fLm
C0v7++Ll41BpOvbDqYH71IReQOx6xgIPFDgaDoepSnORZ3Rlz9gFhJ1eZ/dPG1Pp
blJJ8mxPUjipjH1LmoBXp1futfWoD4AC+zCbR/KGjujkwm+sxSN6dttAqMX1nIxl
MBOn+YTQrzyTc5Jtn7WtRKEbEaCfmT//1Ce6GzK5Klp26LxfwTK9P6QFfTvivU+6
x8ercGN7EbofDQnfZsJC/30IzzSNhATEu2LHnp6vYXiz9axP6g+t9Ko5lq69HsvC
X5WOF5ilv53r+ItdZu6MFMs7On9iP+Nqazk/oyvwvtvDZiaJuf5AuqrOsd7cKyeO
Jh9h1O1GdkrHmKHp1z9F+Jnuc5cRTyOIhzY742wuDWSUmXiy8FFb9KryvW1v8Sb5
FUoVnsSy8MLByYyQCU27vkCoIqCxDfI5odfsPeyzSpOJ2Mu8E/SkHV4JZEPUPRvW
AB3dsn5ugzJoOzp3B277SHg53PIn5bRJSdkQ/OheBpko8POMMhqIq4IH1H8Yqrdo
zI26LCYyovtxKcmjN+TbCarW3SpdKgPTd3q+GROVK2iv4EzJaPhhAWdVEXj4ex2s
irFPASE2k22ObTh2mcJ3BY7QAqQ+wnXLezjVzlnZAc6DuLKCsW0V6Fg+ciMd6Gmn
jYsbnTs4gtNe2WFbKXhPZ2+naRCHaTLazTLclEva3ctXXSMxDOcteyYKb89Mb4tp
i2wfpxTZEtlXtSbe1XxuaLfcWIbD2ZtqYeLVsILRmNqbBol1/86vU1ZnP122nXPE
j7QlfEE6CLcXXoSs6FqDzNu4jkjraGgINoinFrakgGvQRe4K6nw0d4ve4Q2ZBOR8
hqGhzyqkaS++3iaQ67hihwR8XoInlLZLebPD+OcTHF7jLBFFCZPWjQ1baX4AMCos
x+goJXhrZVwKpD+11NrH6n4JKQodE8bzS+CmMQBM9oxuuetOJ1zrhacl5oU6aUar
3aQq0VNtFcJlPFi2v2Acukbbo1+gqg/vGvNyPwga47eyncUGLCpZRY5Q2kpR93Ua
EzSstT8RVy1L64aOdyT1hkopfKKa6dwWN8pSMSzAPX8NBq3R1avpc7D6GZn58q/5
nSxmVDQsGKZdoaN/j11jI87BW0tUZgt67q1m+4W/k6afGeJKBJDuCidrr0HGB37u
00ymNXEICgcxSn0BjekaRRgHnSKFd13mWgPvohpgGDhUWh83TKOKRsWXmUP/QkYC
KCe9SqaffmnO65s2mHgxLEMta9MBGPiwZWeU1rgja+UNVYhFXL6f/BIbYLQpg6iv
F5mufseN3HGt8SMkgPdGjSyfOuYZwOvTaymTG/fHbr2FTentP7ytJaST71keDU+g
GrJzzp8ZdBfGTDAanQgKojiiQb9VXz1fdpQhM3CVAdcaIcR6SRv6szKJdhfnQCmD
SBbIJVxRJ6IW+/HPtELsY+rOpPLiMUmA5HkibOlFzdcYSUpcN/ILE6uXSxa64/jO
jQReaYYjGGqc0nCvtnB7X1rXZwpihNkA9uCLQeXvTl/1bItzoSGDEMD4vpBRr/Mp
J0Dbg/W66pIQDmSRkxUMXnS9hkIEqAFocVsGeO2FnRZz/H5MolvDAD3lMPk6DIp0
kuOkwOe7ThirACIsNmt/IyQlbHS6ZHdczgiHA84k8eP/XjJhwXStXsImrJig1elm
JMQ9F5hqmC4ll7Xf+1LpbORZSfRRi8456cz1iM8e7hTi7EeLOCbRtsDuaTuxlmm6
6Ro8gPHDABVESxXIgR0lkWNJiqeMl1iU/jkYfjo2xvhCSzxkMPHWqyEdMwYHUy5i
caTbjQJj0V3x49khHTYNqVLlUKJL38ncEr9HqAIFq6b4XYoegVpo74IGE5J4P+xj
+neiz+xcILhrFZPJ1/Ul6htv20ISl6wB86DR1sH/CwgeP9UeCBiiIwq8hEiAkgoD
K2xyLBpchYVTODg9NMKx1+0DxOA18S1jH4OgcQZJPXRPDhLHC7qrz/vauXbKZK0Q
VjhdiMZQVEl9/IFVA8jVOHMpyzCFRV4EgmaNfQN2ckFiuB40ij+h6ObpWgY+D2Nu
iRxNQubK0UyD7sM+haqRmFyP49jtX/JC7UeXNzT8QmxHMGfWRUSRxO3bfeqK5/e+
V94O4K01vhVVq7ooyDVFKLmDB8WrPoyl6Gxb8QhB+n/msDWxMK6yfAUrjcrrEW8R
l9kBEiFuKxDBO9IxtQKVgv/MkRxRUF0aspGT0tTcQQ7fUBgxjmTvnxFZrhF4If5N
gFfr8YJB0p1GKVw9gY0lQ57ndBNoRruQQYN/e9wPMoEuvX3qe7iouXXeA4a3BAoG
w7B+Ia8be/+8fIS6aTcPxzDdXXBGeO2+ywlCZ52b8aTk3MGoqEALSAMvDs2bzc++
rvmnK+/cgmKOLkgndXgwNnqi2ri9JJhV0BQp0fbnWBDJTkpMU4c2Xxh97aVrBSIA
wnaLdcz+SGZ6FEMnbovMb/bw9tf5hd/CX5rBXHt42sUBiTMlH9bSH1P2Cn2vK++8
QSU8gFBOjHLe5EMLv2+xql+ZqvmfCJ1nErELxxlC/GqDmzlVTHLdIr3bgpa+I1iw
MfLM3Rktoznyd0wN9KI2keXao5BpLU4FqG8rgMMrvlxIh20QZQDls+qr8BH0YoC4
+V8ArbiTGpGWPthDZddWqrX74dAvmLh3moCAkRBNTx43gvIKfuS+1ekJZbgX0qjL
UZJc09EpsTOdQnomtbjOLi9fpVvrs5hhQsnqXB13jFk8lamkdFQBkBaQBk1lybaT
T8QIgxCuQDKJ+f8AVbpEYsmn5KFVG28qLzJq362Nq6qytErxzbQ6uwkvMmSzA0vs
N8bnJaTB6CHo1WZbbdyAHxZNb6rtuhv3pGtQefWematsg/GNGRHlQ+jEB3pvac5F
4AGcDJLUXY4WagZwLgBQA6ghBS7IPFfnDph4nrdJ1IL1vnFk+D+K3Sw1u0pQGsL0
TywQBgYu+/qvn2ChBT0tQtMGOyjIOVAD+h9cVTHEyl1n+idsNFE5JebNJzpFhOjJ
JZLgNfj5QGdKdaY4lSES47WKTdrtkJvxZE78bnV614YXW+drGs3CSTmF6MKf27Yy
FsNDzGc2dyUyk/SElqVi4LwEad0Xv8bV5LHHPpRukZd/gTyYUwY6IaQ0o+fxbJol
ExZH9rWTvDNdaZ17+7XlzdknwhVmWgp/1/xQxrXaGw+kYnzDtuGtj/lMF6Nm/uym
0esO8emQRDNnA+Ztd/YPeHDsEBMNkprwgyEQu15TeplB/F/xpEyze4D6lxsutyqw
yoU9l1UOf2vXMQTvTQ2lzaZz2vDY3/zj2zRGeajYDYZfKcTLOWGa6gpMa2m7Xjy2
9HsB2A+9vXlGdscl0AxC5tSpnlYDPMg3eAJz/iOaJewt6kLtxHdn9QPv/85KsN33
ODV1SgUYX7d7VrUkyKG3h+Tz/dKsBdxEjcngkmIIJtbVpCj8rJvPMp3cL/oLh1CJ
jNbR3DD+7IPvahBNWlUh75bFRNez641I8RNtyI+qdpn0VVcQnLgca2wRKSG47+Zo
hyVmy/1uMFl+RcWSQG36/7YxLe7AzOVhDD12YhpQmynU39zFM5bga2N8AaWd8d2R
Wy1+zrHxMIuyFgo1K/1zyD3EmAIgQoXlG8CanvP+dxFWxXe1n3AxMRgmIuL1sq8N
zs8p8cEHQ/7/J2R9iBoHf7i4DFFYDfaZORkUHt4CIi135omtHI0PZ/Xk+MDB9UE2
MDntELifQbOLC0MpQSiHK1AtbQyUwIJUq3W83X1XvL1aKUbB7nUJcQk3su0DDZjC
PxV4p10ahky88QMVHvkbzyKrvMqNzZ3iKqtiHhXMS5HR+MKUCXaP9bjRwMbWRLXO
iw32oOqKmGckOCbLyYN+t74DejvkIFRoJT6Je/7yE87jh3LdxFtaDb121CEc7o96
gSHXfRHX4DHR87Ej4OmP/h72FNDQYTl0asZAKjmNlJyX54LtNEwUKBHVuyhL2cX1
pMWlYrnTlKT4B5sB35OzPqBmdEFOR36QtH7q5BUFX+saI5+J9ivhxbIFYqZTTIJc
jjvDomOKO5xHhZ3e4pZW6laL+SQus8FA7bCEo6Wlc0LDIWrR+zRydR/4kyGC7FRQ
CWQe8aPM8N4UO4vm/BeBECFVR0HHZns9rErwDRm0tWPzYaJ16FSZFpJHlmzRPv9l
o/ZlffepS9syQY0BDRGo/K+xpFLHZX0grhaI+cYdMRLGsVSQoVIYIN7WmPuGeQ0p
FLfBRXOoI3LLL/RxpriN0FVK/ONti4UjS+tT0NscTFE2mfyNvSDUfFLQASHpszx2
pV7DSQ4ho1164LUOM0cKfbu3rnFbSqmzv6IkS4gHpuqFVJ1M6Acp9CaM/smYxUMs
bA+MUsAp2hfule01mdgy0Snz8ebSV1LXgVF2s0C541QofWomczomOhGeqLxPZilA
z2v2RKMWlq3+muTdO6Pn/blykmYS//TXIHg+LFBXDeriM/t60ZprX6+YxCfA5LwJ
a+1a9na9zj4CAtofmiyxgIUNuVrS8aOR4xZCzTuETCK755zJpgdbnQZoI4tT8q/u
UkkqHFz+1oViyDO5Oyb9zYDu6j0H6WDelEUm6HUhlGIFOW1F7z2Mlj6qqeFFvR4q
IT0uZ/RxKsjpDFDcIgwwGY39DZ0bEMb0GGWAXoaplApQv4JHInkebOV+lpnFhZdc
F8YmilRW1zhIK0BKA2GogjbTVCvqOzvhz/jOVKqVB/LfG7ZU1dSJ2g+/Juk9/mDl
xSI801QfXGXgIZKDwVkCfh5irWfg5hwvDoofHPjf8YTSWJz3qUTMaqUmWuL80XXL
2w/StBQRMMeFBVW1cqnYPIE3x+Y/S1KbguWyxxZUKdSHSORBtihYYwikYlVsnVTV
dLhAUodIcE/ORykLMEUsB27G4v8BXVZWADCkin/7gCfQ8ISX77zXohSJ4L9fC178
jgr7ZCxbco0FHfsS70YLGug2NNtnNo3pmtbs+SIMGnBvFxBRv68rC6pLU9rs/OEe
z0eiRC4j3+xnpixTFMGJmCwGDC3mWONeuhF5/oNuhmSVAv4Ai3ny/XJA06rotfhi
zARbjJ01J9L0XOmAnk4Ry6JR1NaJuTN8UE77qdNsS9WjdLo3qVPxgiKr8ZbCrbp4
Vl4TdD5/AILX4cPalSF4wOB+mZxCGFGYV4ZySOonuq+oMJIc7F0eMaWYX0m7/GIK
QqOpg7rrPHt+kWQDuj4aHnCo69NpEcWYISOsuOquFbW5lO99684W1VURAcgwCTuy
GAa5lc13NqqZeVpZks+kEro1ZlFbpSYG2V1lZhjwf/fbEBUJ/boroVO0eZLWoy4I
DXEOVvJupz2qeor/0JmEwHO5bNpa8UwRwmvQ6SUE5S4kgB4yk3J3CuF04uhozn19
1Nt6XpFF2R88npf6A7M0AmrNGVAn+g+lX15lhXI6/pQhalX3i3pV4YSoMSJMQe16
ZwDT3DQw3X5htik9ZapsqJikUoiE0qdv0Nq13tg4Q+/rYpv/WleSlUxruzfHqw2A
ITneWd09pWAnjMxDdI0rueL+VxECZpvaVejjIWIcoDBd46CTE8J4bhrzNnhv/oW8
8wCxHhStpb8gS7APjUbwMrGgx2cGg1vM6AJh1xZhFSmSdAHRv0ib8pVkaqgQrXD4
m1gRG3e1z6EGwMIuFoLs9MCCHScelO/5j3QLdsyxH4u41pxD1+xlA4KgcUH4ppRT
tnxS7ZeMLC2rJxtgTeilBB4bTxXL4/7PPSlU4xSn3EMw6bG9RfId9p1eI9x8S5GP
x9ZdRMFaqvQUhorOCb19XZwmjTPt/Qr4sfGorB5DvK7y1cjq+H46S9C3+IGZZxSY
MpT/lg9Li/j+zqyXAec5hrxFkvmvSmYyzioPGWAd7f3sKaEqL7jknCpqz3xPERFc
WmdGmUjCUjFLiThp6cwqvGoExQKPrAWmRcTYwPRWH8Y0Ce9mEQ2msoBqXSFGeL7z
2A2LKuMW2u+SgObYNEfx6eMK0iVBpZ1WwllaWSwuP5VB/W8x6AliuMfgwYkuInAV
8wPu7YcLM1QiFT09CmDoPvLCikvWk6Cv2sQC3smNLk7KhwanmeFj3JC+KE6b28VH
R0otlCft0it7UKA/yGI71Tpa61iDSOi/6dOkodVyycMxwaqK2XB25UlazCexTYlk
iVW9e5Ys5zxMR/hwJSYRiNchqtYsYRuXFN9iC8jKqby0oWxaDsqxAbsBChg/ZAnl
IDXz0cRyoW+LlNOq3YlX0jFbSsL0ugszaqxiLF28ojDVG3/1/RpgDQAetOmxTg4J
GjD55wHZnX8fQAupFTIJ1CirKnMUYJoh/9dBKcrUA7JCTaraNGiI5EV2Snh6F7nl
pINmDaDGrgCjMQ0fwENSwg==
`protect END_PROTECTED
