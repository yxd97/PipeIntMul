`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+pxhnYxB2yovbpHKvs6izhI5SK2/5S87UiS6+qSJlebC8E70cDO9bBTI9fwvPTDr
/F0PEWd0H1GJKQaj/riRi9pdsmcWyssx5krylWJPX2x6+RYnNLGfU36BO9zZlKsa
x2pnt8DUbW7srHF7CGlD9q/+9r5EnAR34K11iCOIjwjSRSPWoL2mfAOD9U5pQp+X
xdJirtD5MkPee77CsMnDNi6PhhYuW+CG6WzB9+Q6aEIrXsC+NrxuHhRcRY5xZijg
XX/ZliQ2K1YtC7Egyim1P3Rw/MhgMN6o7KXFME7chAHVefjKqRYaMLGqFTApiPjk
WO4hA65TZNMUV6h+gXv6vklM/m0pkFfToqbxGhITDQUDnO+Gm/bAm/e6n/Kpftgy
jNS7YPDfpVFfEXXUokRxS6VYaNLjd5xkW1yVB/UmrXKSNo8jA4b3DhLetmynEGXw
izp92QD+Mjuyox4jJ3lVbtzhTXbEegayylVoxeVp3+4lt+mnhk9pl0fEvr2DJy2E
t6nGJ/QtQe9SixgaIr7YN9u//psPud+KXZ1+xKFDfA6XTLsJHiM9wSyu0MKHPPrJ
f+rDvObtamPbkpD8JaXBd+eE751Cy6zQ7pv5ufWsweajZsqo9sw/8ggXYvQioVPd
PpXdc75DktSoTAEZDokm4WkoGDXB+EHzUcD1tgysNFTlEO1hThwBVFeUmG0zsV9N
ILZa15uFBTnRXStOXSvHpcIow6ilQH2zaMfjeimNKGXCGKC6vvf/XPHvcDJfeFKi
th5PZyCqSzJEx4vexiDchceGyF8CJEP2/wA47OJZUwm+04x9/LDlQPUoZR3uT8Yf
ybzZo0gn/ZU0pi7/NqPpLPfH3Jgy5EfdvwMwqT0J0aMuMoyJGaeiOjqKEqwWRtLW
3mf11n92es5ljQ5Iu2d+ZFYKjkix4KBlg0ODLlCWs0LwoUWl4pw5LITmuo7JOBVz
LJ/jPs1NPS1v/OTg2lVbtJheXnRqtzQCXdRYGiSFZtgKnJLt43C9H936wxulQTXW
ZP7kuGcAP/hIBrLCTniofBJ/xSpitaHdk+Vld+pPiWzXjpZaBCPkKsPLmEpN48DC
BJgIILMvantZ4D2hxKv8T82nNyjJEX5L/uTAk6XvUZzX++qyZAh/8jFDs6jDww4p
Nq8iJJFbktV4A+maJZGh60JSuRykMOnPUckKxY8Bc3ye7pHRIBnetcvMTD90teE2
nAXdVvvlIT3GzU4xCn5emTV/8TlhLQAicMYpx8yzHtpSSEE8iicJYzPRBDHBbPn9
`protect END_PROTECTED
