`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wXspgUopyvkGYq/SbxQvubb8UUtdGGQxMWq9mM6yUGEjLsqUbPUSzATjU++hB6QS
/N3TpmevYZc4A6xI2O9w1+kb6DmcQI0IFOVetleBZHqzTsUr3Cs9/s0XJreM4lQ5
1f5JKICIXMA8CkksVvYxfrkMBRql56TymCULH9NkNmblbJGDdpoBxWR3iAo5T4ir
Bew/kl2rrTb04JmmnOYHg5hlmkTUr8zqH6pcVYAhKz6kfKRYaGe7oHQhr+DqM9yE
lD/ED+gHSdbxCWM1Cfr7pwXDIxH4uTYB+uu5N3wxGouPb8VleEMWz2bZhZZdcMQ0
FNIOXFJQs72zn3VCwo6cUm9MiFyOZyqfZqmTFyhdXtMJlYSKvfRt43AydEwe7Y+e
Ggd9ne/xlijUDpklEXWB7yTG1ZKfTy+vPHhH5XkWkDGuVXwQ44cSMMVUY2QrvVMb
kP8aarAHbDSMpUMaaQLEsEqempRK+g1qVdThDHT9ZMiU9Zb+ZRKa6SRJfN0SIkOE
`protect END_PROTECTED
