`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kEC/E554hRDbAeooHpX9AxUcDxX4umxyGZdugLGi8TDE6GTiZYIu2bXKFiwe8hmu
TkvX4qFT0Q/90RGvxL0Bm1aixNq9M7sgY7m70b5NUpjACgoHrFpiRplCI59R+xdx
iKx8yQM44kczCmcsT/gNmYSWw2eVvS0IabGaS21pn32JzxKXC7OMGHz0/UD8Eavy
QLMJXc6n22BKO9/oDi2RwdlXhnAEv5jG5dtZsyEKkJRGrEZ3f3CxwfBMw8kMMDDF
1jRTI2hfeUQFilnIowYwg3nDSjQs6VDQPwe48C6u0mLOZX3nI1ilFOPKqzKMuInT
CI4ArkakvCUmgk8keAxRn1OTt42b8VsfbnsyUEZkOaTIqjA6bkHDUJtanzaYjgvv
`protect END_PROTECTED
