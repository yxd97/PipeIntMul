`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GBgrgVp5cAPK1Jpwbl9AlIyvVKi+8ocNKWu+1Zrm9/DeNWLon3K8uNjApOEqi0L0
f/gijt3r8fbqX3FXb05O8Ay6RdFi5vFopc3hGKDHOPl8K+YJ+HC604qxH8yTEdsV
0GnvyZehFvhqHr+NfDw4/fmv0yxiALRWJESXJaluFxr1Nc2GMPPF20Y6iw9KqtsR
U2lM3uTsjBFiyFg7fKNTDwZxRvzaAhrPLiZM9UGuglGUEG/kQtcRy9jgQrW7/V8h
DhjrKD+JW6XT/UQuxJz8oB0Ph832MDRP/rTq6rhU065Mmus/GqclWzgF5AP06F5W
tLiBtIV7Ycj8L6V2Aip29NTHaobBxudJUcz8BRq7+waoHfsylgA252BNBtEJsXRX
igyzaGvBBROBrNyb+xb0G/NkUXmA5x+bYPsuWgTHN9NhoOrcP9TZlPwfCAeEzf/8
t0n8YqEMvQioFP8LrlabddUJ2RurlD/wMQJvIRQNApzZfF+Jk0Hzh4wwUKTwumlx
rjrZic9FXS7kI9sLyHfZ+NKCt0k53h0USEoreuNlXc3vvaiDRPAOKgvPvtFbgcyu
eERJx2LC3pr8vzUKN7jZxfCl5JiHzuoxCBpCPsQweElok7h939EWTWTRRThWUEQ3
z6jZ3uGF+UwXANYzXJWg+Nj30bNyjlrZr3WoecekPXZRKT4UAGdSwjTl8yIyt5an
OVbgrSs+SMG1TEHJQNouJbMoc68LU1utXq8ycU6hRfpjO+g7sBjbUXoTFoVLLfXh
jpEtBkUvRvd1kFSZ/+st6nPwyCSSzUAUXUbbwtufbva02SwP+jmAZRRlir5el5rH
pEQkibjJ1u+B3bg2OKlT4lIHx/CopGOvCw0XZKPa6gsssdMYWzsVzllSZBS/WCI0
7njKRgN+KdZ7Sgd2ZnEwfFp5Rw+vKAu6IqwvCckugbqbbjyDcGR1OUVLdFVowvJk
H6E1PyDrJCPZTReYn5Qc3bWklGO/LdVtLYNkxZhAxPcPsSorJ6aW9TdK8agi/O+G
2nUuWHIWtl6Hs7xxzLcQBIPTcd6Uc5P9Nw6F9ITf0emPPVEhJHHeVa9OdKAA8Gqw
b+xJUkZA0DBX6buEAS2VNFS71Qefq8W28mF7t7qlB2Y8O1z2c/BpYJu/xd3HjFe8
CWm9uZLXbbgmJKHEDr94nAeiaUl9O8yWQd+KFkYIQfNRVDXn9Aid0FgKoBTs6OhA
Iju5cNCj3P83ZvyIjLv8g7KQT8WrOGEAdGfrB1FjpyP+fDin87RGBxQch6Rc0jS4
7D0NEyXutoRyV0bMdQNz6bmnEZ97QOvTZkGQLECVQPiREDX6u/q4GRYsaiprW1xR
3iqVG7WgEAGOBDpY0W4xFM2zHzT2YwwCNKPE/z+tnO/9DP38hTzgrqG7ivu2mqFy
/luAAL/LtpyyCVqrIOWSNzaQTiNkFSozTzCyV+BQSbCm2l83zWNoFeAv+cDJOu0a
QrfylezM49oEZ0f3ciWBjwQrciq3XVZ5Cx2LKsnhH6BDDkwZBNxoa6jhGfyr2imr
drw8CyzU8/KFGDfH6z4D0MNP67TIP22dluPC/qQbwR3EScr1qdvqMXz8rG6L7eb5
lEdcwO7O9k+FyzULMQeOpKckM9V25/vjksfqvSbpqebD3uc7gfc2+4aTFKCHID0p
zfRIJlKPWTF+uNfaKNDHjwBCcWVtoDUCKu3i+/BesG91j35G5YMo9A2TdGFb+soH
`protect END_PROTECTED
