`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QuR26S4BwB2jnSS3yuA0eqYqi7odZPvwO2Igs+E4bg5729gwu0IwJHISDAOt+qjZ
0iOnCTsuCOwAmxlDFKPA8S74AxK/kFu3sdBAJ4oYB5TrddftAsKiOux2i0qXN7H6
wOYVt44KLXHDlBeZ1868EQFqfIfOkQwATILC0zsssW7yUEOob+kkY9sotHbnR2O8
JgbkKQX4M5W4bXKcCYeeqEt2LDloR9g015GLt5B7hqkVB+Sc5Sh8BITXlsO+86V1
2XQnFx1czcylwi9c6tDKqgrr12X8EEMLPT/5btGTsoAFZ2zFPar2i1wyPemKtxJP
8JQKpbxkeXwRrZkMt5KaTjWbKb85SbF5R4R2i2opGl3w5A3roAwEgydhl6IJc9VR
VMiLuZcuk84WIYPd5XzaPvLiWT+pUIyUYpumY1+uqcACx1bbTaL1yZGtibfpZjSZ
E16d87rK7yR9dP7x4j+4w4QosLDMAdNO6mInOX+TS5Q=
`protect END_PROTECTED
