`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jy9NCxfqGbNGXA7Wfh3JeDV1Z6yketqrurvZE4tE0YZO5i9khv0AZlfXOeexIxXq
D0I0eysxNtNzk83IsQUrn0o3raC5um6XsmHreYNcZ6ky/SLiRDLvvQN4/iJ53hNv
fQi7AKxFW6QSf3jcpNE2Ev4xAUVf6HvoDPW1c5/MhwA+5q1qyUA+34c0ygiljadL
YkXI4Ifveyogbfx8VrC7tkM2VW9EFdMcCZqBbkG9W8lgwPy6wGFT43r37F3wFlfq
hwaotLBARq8ISPBQEWXTjqfOf1oAmJn0l4sxoQK75cIkgJ29WjO3Kjxg7ZMN6BNg
GGUVTfraSjHvvFIVT2M5xbFWVdidLZaueIcaN1cGhyTxHezGDlO9lJyO9KBA0k3f
/xVQ7zKevE7ClRpxh46hJW/tyC9w7AdsUl9vpMn7gdhWikFVje7diRqXyetEiQBC
`protect END_PROTECTED
