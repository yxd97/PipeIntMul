`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CsZarG8176Wu/FdhodMN4a+XpEVUytdQQV36UApcjIEEIjZqPusGZMdQmtnZy6JD
6fxtROR5QNmNe0qOGWdVs77ej/v14HduOJI+ClAXoFvsHKecOLFt+dsUNHYDl83D
apTMKVHeniA0hXb+Ai2iWVZiLdqtzUi+LeLawcssIJKNqosHm4v0+sxODz/+fb5S
JWsU3f/ZpAHqH0REhxqXAqmTexZ4WededozyHbHKpzUhiKE46tRhky6WAJNZMmfs
CiJwEEIu/YTZ2YH66HBWPa6wapoX5tWNb1ZJl6W4Tnu8SO8C1+1MBCkxqTwLt6mQ
k4VgUIGlAWx4lK4/H8L+OaDivJSG+eg4XfdvM/fepDXru1ujxCCrHUUuU0929tKY
wBS0d+GY066738Vck2FOi/Dpo1fXbtYrqsWWBrignl5LB0nWHz7oUK/Qw5rl5tri
0DMouMEKQO4X2I4yukwrsO54gLgRMWeHYTsIRIbkqPup/qU6fyyE8jk+WfCrgEb6
2bfwOMfKo4MomG2EK9onK7X6/EZv81wYQtORMJ7FcFfxG6hF8Jm33718y/iMUSHQ
gP+Wrdu8mkkfzn6mAoDuAQ0KNC+y762tPJhSEMGHFI3mj9a3+2vMSPy6bgOhKDeN
D2C1IQBGaxq+M49WlMEXC3C7iXfS74gW8P+jHyyIbMZMQfloixceYVT26pRzCRbL
ZSSkH7WwHJZRu2hD06BCVu5mnE8KyhcXWMIek4IRPM9zLLSx16BSuIbkbzccC8ph
6qGDcRkcwok7RcgD8VoLl0zAjxGM84qAsnsbiHWDlBeJTdfl1wpC/9C45AtnmFFF
AAc2EDxJMyrugrFSQKRmI1FinwYe6lSP/qZ8e+VbEEdOIVSd1thOY2YXZOPXSkh5
x3MYRaptOi8BIHAP9v6Tr444GDCuycBOuvUjfeFkZCrWQi5E1a+CEtpm4PSi9zh4
EY3MFXO4G1nYmEy9KDGIGpMZJx9oL8KOuY5NlXD2RpCLHY0B4FQedj/wew41YhBC
l5kH3zekroOsh1l8NM7G/Z43TCywnexdu0KRhX/X2kLhKQ3H49T1QMvK2q5OSVHY
3cZgshGw3qvpwSqNiPHH6dcQtYgeaM+aa9umkK1PHlTu0PwAztiklVmymOhaZtvb
SNJZpCO+QJmGu5OoSwCrEhZtDkmxY5MTmcdsTX4qUcdFEWrQRWFDVAlxNQhdObw/
osUZRl+PZxXGq+ggeBcHiS+4Jyec9SnJ2z2yL/e+30mnXBi9DLd57f60RpX/34Ep
UVTDw1AfDYa3pLJRmdBW3k7sZelHJ9JR/Htk/Tin4M3I+sT4TKktgIvhzfMG/nr9
AXHdjm8vAFCDBCn/MrCtGgfVarmYFxDVfJtQoPPyWathdBZQ7fYIjoFYu+vrMfZw
IuZLCk5mwRW4hKkvLBWL+3wZtViy1G1PS8DuVs+6jDi8YARTO+cUmY2Wt5WrwsRs
W5wVkuBuuoGME9EoFPTPjL+Yi+2GlujesJ8MHWekGwUq+OfRzLvADBXhXM760QLA
dXBOcSZPIiU1WAmHX2QumWPh1mFYZ9qbnLg/BiEflOh67oMYfMmgxow6oN+yP3XO
Q6yaW8HEv+MY5q552AvcEUlYF6mLNNUmbcESCXWgsp6uMlfQgigs7DJM8gs6GQun
xUothMTL2CUJJ+WfpCJz3Z+D0eEuUCG6+PAcHWhen8QHq6Lz8sFsIUSzt8sNvHrO
31Zz7rKnz7yP1QamlbbruquLvgJKEmwOWmw7PMHtx386LyICr8PRYWd2eRCX3yIA
e6V78h8SwuVQcHZ4BNNzN/979pF2KHnTiLS9s4ehNxHVEY69qi+HubSDYlCBvTAw
rb8TgUhGG6Ac27KIgjMdMUKftTi5opeoClpuvxgBm8TC/RXsQqSbOHWLlSULBVo9
u+FovpSjU0hgVq4F2ovJCc6ilVvadBt6OLUxGuc0R9hyeuuWHMw5viNuLosse0eM
KErCeZQDRb4LfEfVeciME9p8j4nkSwqGUDn/9nWNIKbiEzRj4NPa7DbpwKrEyjqQ
Oc+K0ytlL2WyJGDvljSF0c55DNbp6YI0/Z10w1ta3Id46bB/bRgJg1kditPFJYzn
jRU3Pkl8MGNSjJdB6RMDeAIHkur7iuyO8YlS6wwZIIZqF/AztDm07zxGnJK8SaXj
mIrYa2tMAO89z/gL0HjvNPlGYxYT5JsvQkiRf4pnCc4dg/B8ftdmty4GCgkJT5+8
eoyrOSYKuPLPVR3qYkARTStjL2nwK5gr34fap0lBiy5FzeBBG7ihT23sJZaxRGfk
i0LgvUCe0jHmPQn9T3RH6cQtjwO4WQ7ITj7JlsYTLGxW9yIK7haKxl6hhabWqqdr
HTm5SkHs+Us4UTnl5ExGP0U5FU43IGffYwHtqhSW3ExsMrPt7uUzjmufGrCpG/e2
OFYKubzhZ1z6G7r/3x4AclY7OYVIqchdXfrNZ6qA40tpRc/TSYaTK7GIFr7FadFK
zKv8BzJ+JY0h7+bsY26REw5slMSxbMUwbcAVDr0dSjVxns+z3G8gzt3Do5RtLzKw
BvWF4Nt3o/jxkCJcWwY8stEiQ1K01uP7HYxJnhfESGIM0U58xdI25FsbfbLGzgY4
AjtFz+x4uVSdyv+G9BB3zLrcfQECz3fMxHGQUrjFc7co4eJXe7BsjwoyXInKXrKd
Edc/4gimTG2EpSo1Dt8o4GKDBAQlrFkf8dkk+N+PYowyG4uZnJK6zeza3mRbADGa
3y9u7zZGq1S5coenROk/8+TksjWu2Lesy/zUemfBD2ZL6L/DokEMBBPBq0svWIIm
zCN+yFvlTNdqkxsTnU8Bd2YNQGT9q/ijYkNlfb0JTEo=
`protect END_PROTECTED
