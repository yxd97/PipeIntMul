`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C7kxs+8uS0NJbjL3Mo6nqgYsvetUfa8OcecOuUJ0PlA+I6UyoCuI/swp7YRxGuD3
SoDHNx2U1yWDrNe1WqvzK4WAXz731bxwOir6k9aoL64SbmoWZeOhmN1XR2d+Dcbo
5iaU762x+N1ZXUOvclkhTJh4WkJRzhRSMB3I+U/POl5++r5k8fdeg9yCBcCusbdb
uLY2X89QJomLJI4+MjonU9BpFa6+UNmGVI1cZKhUIxA5jtUlkYb3JuZVfkNYUs/W
eI3EiAvvhVFgWYU0yCzXDSssE/xN2RWBuGO1L+jUj0t+pMuRMLs0ryl1wzL14FYl
mFMkI9NJdSOY6zu0JAhRJfJAR2tg/1Kw+uW3LZPChEYVk2GlaZTBFDgX3UzRTD3D
0DuDlG0jFrYMS3GOU4ZqNm6dY1Ek2xwcvDThau+yztymNeeceEB0CexR//7YQIdR
8b8pzRTpl7mnmz/NLQQT8a21arQg8kPxso1c4r8yy7uH0+N670Sh0oMYyMJ1NH3d
63CuYwV3Us6wEczYMHSlnlNQ41JX0m+1xHIravGoswt5Zpwpi97YR3Lb9EygHw2N
s0+ppUqJHIJvK8FSjYGvw/6gYMxu010U59QzFPJ1qvOGrvEIz5SO0++FfXCnVqLI
3kGCe61n3AYABtm/hHR2ons5qn1qFNXbsdB/h07leiQTnfrO8cW4RJT5lcNEOp2Y
hfbTULVEgpC+Q0t23tGtKzVGCVA2UsmWTyIn19o4TUaXYW2lSVUJo+ZA/dnh6Dd1
9Nb2zxEzAaQZtAVZ08jLQ2z8sOibrgmRuw+bv6EOiAvuetSdakHU809o4cj5K/E3
PwE9nKqhSu/8T6iujcfMBpAn1a+b8d4ldqJktSv491Y+tKiKP7s6x9LOi/CoCfEe
13sx6CIcFSBeMau3EzE+1Bo5/WKW+FOVhPnyo3n0EQ2l3O9Yl67hSFETCFFp4pVv
teXrgWdrftYp9LMIj8UR7O2SF06HXfVM0QSRuz/YoTbpNiTsJrE3lKr9OHce6A4l
zIDGhrx16LgJTyFc/kahYSb+JX/b0OaQ/buDFjq36pk9rMtsIXfhonp1syxudfzv
pcfe59UBc4GyHlojMDpJkKKLPVpGlRGCPKoJqxWC1coVMFqSSsq+VjNlm8KXTlB+
TCEvw0Vx5kh+0+MrQinunhumbaZT20O16uWnQOR9ia7V+A69yKp05r8N4TdClSAf
FeX4+4ZzKxq/ER23u4b2hbTXO1frHGk2n68rH2VL5ZvEMtkqlm28p8uErSs0Prmn
+abFdP4DVb1bkIBnX48oDwyQD4G5T/fc3jrVD/F00aU2DNHT8GGChUfYQHz6TzGf
59/woksiq2NVZdbp29RmAu+qT9oQRkaCQEOnZAOY9njzVaATgSA9FOUpFX/UpGs2
PCc+TMkNNhkC+wg6wtamqw==
`protect END_PROTECTED
