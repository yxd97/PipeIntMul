`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h0qaGVU7xmk1MwV7tD/L4s1WFhonCUOVefUqYcfeZCxTjCE2mGk7fM5BrLOF4Xan
ATHWPkc6mZWkyG+Zwb6OjKOZnLtvOQgrN7pC2ZaZdyn9mz8+ExTOxNF8svMQB0YR
ET3//qsPUnADUoh1MndVCUYeOz6DmxrUibqTzE/GZgFuZOTzZlpZ1CbjKQo+h//b
ShQ8It/uBdqYBsu5szD6eZGTa96ZKgldAIUlrhkDoIlRR9qXOeXvaZaHbqN4SHV6
E7f8A2hmjY7/ZHxop1UUzgzA0bEe9wxAcLJSUD9JF8kAnl2NpADUq6epQ1s9lmwj
x/fTSb0bcpPwvlpYQtUPTaUUFQ26iCPAmmfyBR2wOKmTMWZ3d0XeqwYUzIBFNwuo
0NfOdmyAEDmMzhINWYK1jnK2iAD9+Q8aOrL+RKmeuOY/yEj0p5XvBqXn7ZziJRqB
DKqR7iIN3xiFmbpMJsPNruqDj2c/r+eba4FIQw/DVjXyoPCRACUTYwGi5nzPTsMB
6L04k5pJoO9XFNfXGFfN5XvZh0GHq+UVuyHImGlCle1lKlCdGtdACwDyPdIlTK63
BmRTk6oev5HCkA0MRPbORhiPK8lYN5dITBwOMp6eEq2FlNIx0ebPy6V3raxwTUyb
j8gOF4zukJMro+E/oCIjz9l9s7Moms/c+zp2d3fqc22v6wF1hwj0syOMyh/G+FFX
yxaGgkJjJRzAUUJbG2uiK6WsBz0p2gA2h8fVRKlWnc8YmkaRcLW8mXekM9oN8sbU
xktG5/2UTpM7Rml2Dh1A2/U03upCI2PrPKyzThe1zDV5d5qiYgrsGC2sdEaLPdOl
`protect END_PROTECTED
