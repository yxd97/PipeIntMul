`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1pRJJ+ghlEa9y5OgAogM0cIwAPsgJRMVcKemA+sx7pJAxmiFmuVLUq7XvNtqHwMr
HSdp/N9qGqwABmygLvw7qIepSFm/GrMXKzop3bbH0TBRKmqLdHVrocwk+NrElBRl
LtCAHoWWAqB4n67943qlti2XPFUDrl5dyJ04K0chEoDUAvGg8KBo9YhpsO4EOHXg
WpA/5Ry/LDtBalb1+fcuKF2g+kMcyTqHMoE3fetQDnxv6KLRDuKy1h+x3LKqg3Vw
mI6DO5GPjVIUXQXVTQXcs7FM4fu558KyEaTuywergctqCpcIVJEnx0bHmGjGTjse
/oq9fEr2+ympjU+7TNjlhuTQkxo1btrtQ0gzbvQzcGuMEQTlo9+rJ3Tp26CfAWbd
1QBlqR7+M8IJbsdwHV+VGw2Qt3I0Se6XoE+U7mAL2JvHfa+wiZL09/UFHQVLGl88
r6XkmbubgzlxA8bXC7IP9qejwIcijdoZEIdEwZsgydL3UxNva8WcUpDPcZimdUr3
1VTwKsYSVvZeiy+eAWY0Aql2ek5IAVp/91r07r2AnufOYWrKY2BEuaWMB1Mt0BCE
6nyYynfMx8CAOW4y8T8SiZKCVhZiwCTn1I71ndVZKsEKM5STYkMb6JtkNBueW3rh
pBpv1J6qgOB67kaRkKwIi2cHPJ1T1P88E7WQ7C7Ipajk1TW7M0gG3wjkKORCoTKq
dg+aGdgFyBvs5KbpgfAseVhKiYusYxWDGEqWPpc1e+s8gYX/CysKNjU676aNYdjJ
42DKINUPco2RiCtJYoZN09ZAJRCX/i5E6Kw+WYAR2UiHuywNA29wzpsnjJtT1kIy
sRgWRTddUGNCC5Mwp8JBZMDO2OVs/d5FwcnIA84EMT0u6QB5+I7CaT9r9Z62pu8+
yXphS/rvKVuNfSyDhdA1gXDGzAptD4e8lmDQmiiVngdPHuVy5sLRyfaT9I5E/Fj+
PHFPQLenFBqkZgJIhl6yyXtck+FIFFzf9kqPhFqwIckfjq34iyQ7hVcbr9gpfsp/
5Fvh5XbbN5vUq1wfxbL+swbagoDV7gcR0ADvso4LIWBy2K7PhZeitVDIc1ixgoyz
oAHfomnlzZnWxWFKziue+Jsk4d/scgKHdX9gk/38ERlW5Igbtpm+NsSVBb2xBX3X
+83IO1USpGirzlRWoTwSQNBumEfhTjbvkPNcYa8y2SbakiJtaJ0DVhhCQfWU8PTL
niLwg9CdA843f8Q+PWOUoehFBmHrvwX02FnSNFr7tHGr1fa88Dh9Q1NS9ofyqcX7
vXGAzwvu8Qps3dp4bh/i7JMt6vQ6gsWfnN0O6vMpBL4V8VuTUcopmQg7/bixJgKL
`protect END_PROTECTED
