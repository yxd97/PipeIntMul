`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n68MAI47fPhOb/4Yr7UJmsDZLG+Z3V7dojfLOpH2X4h+9LS56gwdGLpuB6jEO6Zk
4B0vXfERvGwDrWo1UFVjXN97O5OG4Q0yStrUBiLsiKRM5hTWwHNhGhgyabyc6QFH
fvtypQjFacxXeb1yB2jLf8W+T6XVUbbdtzqyDgKIJWlg5+sgpMExXlk0+of2tce4
KEZ7pDQbwsrVQa1q0P6MU1IeMyh8OFniJ4Xzu8+N5Q66c9msR2KAbVRhlVHsyGFg
Y3KCTOBqUG8drRZeSNzuYLOvECr127K0JQwq3tGRxbikjR51EM7RaGjKglZwSnoE
+IGEe+snNUYsaGEFS3lfsQ==
`protect END_PROTECTED
