`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qFC+ZOQUVaNQvZckPetEcp0kqj7x7XtL2HHo3nZ5cu6aIAJGk+vbjNCk557lRtL0
AsFaSVgtE1Sj7kYrgOH5wS/Hc11t7kovh8zdFmAWv51GbZR6JmptpqdzpkZRY/I/
jM+lmOgTtK13igVU7FkXNVpWCLwwYq3Az7uMNEmpe3Yech6Vqfd2nsYxb+G37XDm
FDd2x3PlDljJUMN25VnjDqJTPt4I2DQd7CX2bZFd6KpP/aRoq4unBV9myCyz44U+
BW710wwZIve7SOH92lWYTHOBfUq0KqYANV9DDJBBXRA1mYvM8LNw6QvYMA9XeG7f
vs0vcfetNvAVOKcEiSmILBamZyIYICMnI0i1Tv7fWA5Y4TtqBDi/MKDwb2ZmWy6v
LJ4Y9O9fU8JJ9WNjjtf89wPGsgNImZInLTNbU+kp5cCrGwjhKinjW2v4ILj6WExV
jgY1BWqwvWkt8mVTSzjzoMRh9IatgIYs7WtLZLdf6zVg/h7EzVT8ulKDxJAGugtB
07i0aWlzXKLMrSl3G0VZ7FVtqgQBDNZODsqzAFXukfsO8rpdXdEzZI5wwdzYAN+m
MJpsOCMeJghBeGc5a4pCSbjm/mctMs8xnyioJivSoDwMFj4RxlBNkn5KlqtbNln+
ajZC19E+lfKBGWgKqmiEiX2Y0R6TNth7HGaDS8vKxLo1OoS7VBpckDLlgME/t9MG
LtMlA1OnwpupKt30Z0hi1XV1f/+2Qnk9Fc4q0v9KwaPr2mcC8PMwBAk7K6t1ve2K
2PZ/QzlzXLLRw0oxA4BSQaWUvLFYbmcM0gIlhybbGfvkKfPiRs7JHM93qjXC7aQ9
66TyZWOrrlt5Ic9+6wkEJ6Ni/KH5UqbERc/xmX0K73UUe9KMlv4Gmo+QX2wtA6QA
orVJuszXOnZKKJESHbI8BcZ3SRj8FQ81j+tz9atVYCSgIUoxSJ3CjMZ9u9jYErxW
WmubHFvOaotEglP2ZwU3nayuCj7G9UU78wop7cMnLN2cm0tMfqS5UBGKv7+QqP5y
JZa9UmB/fHcYotc3QA6VSY5SAOZChId2ReM5746bmxNKxFqwQdHCbTo+swzY89CD
zREDQjTaNv2RODk4uTPWusQJiANnuSqt3xmGv644VwpzctKKdxE8T6QjHb+l+qkn
THoUSkZYRUaW5MqXz8jN7+C2Ph0ri1HkUJfczWBhJBPtaw4Fm+JwHAXowc/kT7B5
/tLxHVPL4XWbdqaSZE1Go0pH362hkNTnZNF1miO12KxQo81YlWjtBSZU1Ys1qlis
Wg9UeLds4W6j5rj3ONwEcZwVWicVbURYTManoADv5bGAhe35SSnIEMs0vkWSO/3r
qMhQ4pQ7KttcHIqkOCAkbfdrnCxy1I0KpRolLqzoz2TItvz7c6lHPWcbZIHBkK3m
fzFKD/Jr7RNgHu0dvzFSNoKo5Cfa40qDsxwMeZL5CF69Zx/To8e5kbkBLJRsIjTV
fsYxeh+k43sJGcMB2vah3PAwcXiQPFLBicfhVONxWEWjO+Ip1/Fq9AAjwx7FDMgk
tLBb93JIxitdcxdl5LsPnSUxEAeIqPTu8pS4PVWZQRwCJ5CBDvNJenR7FWNFnYXy
p4bzUhro2p/2EMs+gpoSk9Fz8K4E9Gda2Msidc/03Ns7WdEmZKLDRkZthEt1J6Mi
lEURv6JYB44zCuO6rCGlcHOi2hVe3O00UdkARQ6aKfeI6fGWLAIxqwQ5y9yJ5QuG
Efw6xfNohtsJZ128tRd2htOC1x0/6wWOH1RyInzXx5xxzaxfPwg8HaSLaCFxijhP
arHx8yvS0bJo11oorzVTwNzB9Q+VRE89FBo6h1rQ6elcbFWmsD95X+283Mi7sBHQ
LqI4hiXeQX12KjDeRS2elFMmERzurXpkjBU7GmiYiJzGvyHT4Ex5tp1sqKnOcHXM
eaPalpPpftErpSAdULfB6867VThjJSV/WzxFD+n6Jp5HWCCQobWKDMJwuaon1DuE
x91XCMJI9hPUbTXBpOmpbfKtmAKrfL6xYs0VB4FC6dJlGV1MDDCbQxeUKQWa8GjR
HtBfXyDW74oySr7Deb6uuJZ1LX6lkaOvzweK1M1zkgzdIpKzeUVGlSqda3uvzw4y
GEr2ZvSCsNDXGGYe4G9YhOj3Ym8o/QHASGRx7sOFfewumI1VGZbRywRZzas+gae1
mPp+WNxrDVUYrNGGW9ginr6EAcgYrXsYbfu+RrTG8kKKfJuCqe2/olwGxbRw0gZ8
IbcaDxcLSoM0Sx7t4An749KqZkAapz5EyBtQq0xC6jAYsa7dpO7+Cj8LTNOanzkM
L1JJ0mchqoDwILxngyAaqVQD1R8wKABe/bPLr74rbanyl8PgISKJPqlwm99RvDJS
0Hjfqo4tAtBllscYpl0xhQCmTXwNy/2CbEqBddLKBDzlipf9CTleMiEKkXFvDQK/
S4jIUSPrn/VdPUTCcUYjbXjM1lr7Gml7qM8qMDt90y34zXCZykPjibhXOFXnuV4D
orhgqs6DQbu7O0QEkfx0S4x6nLtBqEiQL86QncDlAr8ZQaM9JM5iqq4KUzuw4MQG
14nulr/9iMoY8zLV0DEbnUeslk9mE5M/x+Ko7RdAso3IwyZXj5dbjIhaJq7VPqSY
VypdttUG5jMUlKu2eY2H981wxWz9SiwLr27oiPeo/5nOlOacrx8QK97WiK0aBhMq
kz4EJgkFLZnbSJm0L2M5MB6EdMb3rJIF14/J9z7Ggjzjgki0nHN0muObEEHS2VXR
ZINXNFJpe1wCdaUyvrk3B1D3sy3AXBvUnCKwHUIHrv593l87egi/wdr8ZCtCNuot
shmLTOlupctVOdg6/v2Jvz9Uxcog/R/0FLFKxbN8Uhyy8XJCvMo+8RP+6X85NGiM
/KXJkKldIfJsSiUzoLDYAuLYuhv/hIlKws3KBjlZiSvxcnD6HxnTPGBUgxjr6vR5
V2PUHp04PqFwL19lI/5OnC19HSH4orL0cLim4faHWMzbl9uKRG2kqEi8GSNvjQPS
+pV+//lu8mXOFVXZ/fVZ2FaxFagOPtVnoPaeFO1z2PeuNolKZb8CVLM4MHMGZbBp
tduRsmASzVoJdeRD5POW0/6wuMAQLj4Ht61P3XcCSd85R6Ek8AcyeaWBrH202JjX
s27CNjGs088/+CFCvl4C/VJ6jxpPZtvyk/vR1hoXHqaXAn+FoHDomT3WUGtp6YVc
Gl85trbtRyYtcCq5DhjBgXepNIo2tm8bMCAIyTG5DJcShG0YNkL3CfwEGE/3ZUqJ
S2owZo5NurGCRDvsR0oE3hksbVAia3bHicsjDrMiU7p/3zkOzw3In4SldbSa7p3G
6WSbd2QWDqvxIRHrhpI/zxi/5DrC49y42ggGeOxF2PBGQudCLbCkrZJpS/+j4FAd
o6pQJz9BGCH7gWPXxWlUuWt4CXL2vToOgVJU1JkJSbHBkfl+Rn1ieR/ZzPZshGB9
Hd+H459UkjDVDRcdwNymtzs0fqXOd7vL7UqPadf2p2/WE1Sal1/80xQQbx6DW6yM
S85ju/RM3L32rmlsnoUz5Rf7L9K1+ZuHP29EgUSck4AI49lhpRO7wUpDBXP2rM9N
Zg6nepX6cTEirBFCovJALsRhiULt0cNp4sLmVriudxvh1Co+cKU5BQL3x6ZygXBr
L/WrI+TTZkIqEwkLGQ2JlgpOeJ2SL5rGo40k2rcSwhTj+7IPKNEmIXI0ofV+caNO
`protect END_PROTECTED
