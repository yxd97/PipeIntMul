`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o1HEU3srSzYV+Ol3U7+JsPFGG/YIDbbnOD7QBFaangPSPBuxBjzNg95+Kxwmc0Np
makXst67pCbu3hxbqoWIp6pH7VRDsVm+Iozpx4vouMBXooe/GPl1j26/YBVTiuou
4fdji4AxTeMPk2nwaDFfQ0hgAWhVcjp8r4zCOrYdA6jbK2qSE1UT0iecSc8ujAE9
vbbkidx3sMXlsRjuhVLCVgvTrO20XsWn5NfvCfxRoJr6CnlIcAtOUBGe/Og2XNSe
fLvE26bnzSAHYPu4asrSRNm3iLGHIjw+T32CryMDj9IG2UKtVqISuGY91NrzIX1G
1WeFe7KeoTKoMEkbZH1NvSotsFVBfdNaifVl8ewDFic/At5DlCRtjTVHk9iY5ecf
A3m88+IxMtxVAaabHSovsHwLTYlE/AT4JRK0jG/2cXbZCg1/fxGqoC/BaNA9OmZo
MkGvxmD67S7RjcgGco0f3pU/SPbKNMuWezADyMtExp72xkgG45EtgZ7y7my/b4oM
fxZC3kUcMG+/G8J0JA4PxibyPQeudxPKn/dEBp01Mi+0adyKEVyT2iJ4pnHaSS3g
`protect END_PROTECTED
