`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hZJLe+M8OXF2YgSat7ijgWlgecI0Eko0hU4yjsUVJm//rgWaog/kcitvOp+5bzqm
YRJvOHgzRuTIl7HocbQntbXPxgSko+ZEHC4Ze7dpqlFjx9yxEhfWVKDsHRBJxDtW
moJhdsFRHmMhn77vzsHy1XYJVQkHQibGqMAHPPCu7KgPSqqjlhyHvWwBxyjrH5EL
TgsxM3h1UGBV6+DPzzmvvbCF2nKIJuz/CCgGie8+mx7Cr8KtMDeFKVLIHTxlhmNl
VR5TTh+zKaFwguCYd3tDstYltqoZS1ENR0LMojEbiX6ZanueDb0o+W22hopI3F07
P4KcuiS4fDjGo+Mm5nJFYGYWrXLUkk0EV8FXJdKqoGEBS0UGqRQRCUGbDTfTaaf4
AFxbCgf+T2q63XzKZP7VvKGH0mjUwTFHSKNVlUy5+t6xHBiqXUZV17A2mgYAvqLP
kIi6ePg5lZqIg2UGs1nRHHt83Tmu7r2o8SnXek/pa/37Tt8+55ob/NR+5nmPp2CF
H41kw/bakdDxOjoNnSH3XFNotZRU2bPGOkJD3ZeGtNlhhAIL6Txw8lbrkfD8n83Y
6H6VvHpVsoEo7njZpXCqzXOttQsK2+J55W/N2zSAupKF8/d5nCeCuvzI4iCuxvPy
D53SnWJcf2aqbDDMyDl4Vy64XXyNuLaCNWXgJj60p2GF7bMUpedlTiw89bqDJhMb
1iavyDDyCfWOWHPnE1Wgbg1PtJXbZCV4O8+tXchjeyNsXiTu1lKzdxGaF/yhQwsr
oX6F4ZlnLHr8hg4SnU8G4g==
`protect END_PROTECTED
