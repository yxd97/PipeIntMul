`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xp/nisrb3HlPHAzTPP7WN8cvf5r0qPmRYiXij9lJJ8galCiwatgy7ip48TnXtrFN
8dRAvw8myWS2AcXtcBdQdzLXhz14uD4v0n0GJQKPXBXCCSABePIhg3Ths768foEx
03S2BeaIPzKjmNN8bHMMsdXMPKT/5CYAejDdZzau8K1YLScFrvY9Nu9n95EKVANl
xF5bJn6dQbjLu9FxRj0v3hK5dKgjYJ5SE6/lFd51LxeJsuEnahdqp9VKwFN7HiRJ
rfMhnJSNx591Y+GyaLaD9HCGyj3r7v9QJiPAoM25ql4ZN3YjxKnA03d6Rixh2UhE
I0TlYfnoYiaEVD9k3ptV7UNdjaoZ/QTNjMhF1ew9RMosQBiW9yxOFaqwmHisvZVX
K5gc4MbmDfWK9GvhmbOvhsf3hxzlZzP7tSXgAJ412lcGUfD4Ha5Aq2CDAzZ3LMyn
bEaXKpiswgPVp126u3YC9o6ba1YQxgQ3POA9K8IS6cmDDrV3FI8zX9OBrPqz06q8
`protect END_PROTECTED
