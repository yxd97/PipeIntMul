`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xyzSNYjS5M1ZmggNPWAoIGwRa5pUhLJ4ZRKleTymPZ/26tVyAcFIgenwUZfpoO/T
CDjrZmH3x8LlJYViFr/bpeXUPkIeCsvaL98eWuZzqLK2FeFsmyJF3t5oNZekTRDW
oC96awOtxtRJnbspm2RGMT14v0/YGTEAh+gZpie1lB8K9EBCZ/E5lK3nH4GOT0SG
GT1gQ7ic1idKoIJmhFLQx3G3v6eYChyfgzX7wAEEc/QcwhT9pF8K0cqyuUesl/n3
0UYsjcerzQvyi11QLL7XG//2TPj6dulyKm9WrfLboF77H76RJ6sImX8pZivoOs4z
FbW9SBcrqhKXdFJdSZTzzaj9oLrbk/p8q7vhbm7okZ9J53w6NVvzHdxnkxhjBnBM
d5xVdaK1jNYD0j/+nWbJCeFi7JvuworCUAKmBLCBI96hB4Uqgh6cEv5lbLXeTSq6
WrHBGMWqz2LUtfgdS0MRa2/ZqZmN+RHIndO2NabyeSZR+zB7DEzhsIueAgPaaJeE
iRrLeIGXlbChlM2KnI9ydNLM+Jq+RhZ0LuCDyxOMqFoVwrFV3Oi44FOjzlJzm7SN
u5U6A+FpAVX09Qsi7rY2qMh6O7l35jQLNB6y5cz56NVjJZNsx0N2Cs4NREZiIHQA
O/pjsEjIowjbOjRgZEFMFNahd+EHCz1+Hh48dgGUtTFcQrim4bw09wOENKwR7CB8
6ND2eVW3bCtGeiuhZfK65WwICPhvm/nazgI20Sz18Ij81Iv29dL1A2YHZXwl3sw4
dgz8oOLlUXv6c1POT7PoksafUFGkjXEKTtXY8dJp7R4F9lSfthFRG2zu4id9hI7W
mOv4me+HQlko4nM2VWuOWSxOsK4LfvMEWA8zhoWR3B1LglbLaao3MqadzCLwLhp+
9tsdtOPcGG5vqbEF6Fd4b9EjPFfv7wAdRHHTN/yloBn5R0iN/FaSicDZ9GdcBsZ+
`protect END_PROTECTED
