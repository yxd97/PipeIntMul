`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s7tR/MqS6Bnj92tE7AfZOA1m2Q1L+qYpbhS8SEVPI0kGFhgLOdY6WbAkv/fIL/r4
vobreMX0/RoIAW4tc26zewtAMLAo42Cx0uIqeaT+llpjO62LMkuhvSHOkp1DBACJ
Ixbog0l2NCBETAhmThxwkIKab9N6Wvzcv4ZxKYr8QPvloqzO9rNYdD9woag7QshS
/AVVhBUw0J6L8J3BqeX2aag4lfKicZ5nrUJ6sDLROQcMOm5i+tF4P2gP0oaJepLq
843h9cnD6hyyBO790zwIPgGNJDn2kLny9kNKLrYvrWNZn93on+HDZrILgHgFbqhF
nD2wY32rxQIZGF4Gyd4U2ZEYiIqVyTAyUy7OOjOWcIapfbH7oI3mvQtdm8aVYWfR
NqhMAwqhdp0PV0Vg17h/TQ42d7azq14IdR4nWY9bgmFctl3IRuoeattsi0+ia5qL
o44JEUrwb/vyzswKVQKHi9+SXFjzzstJy3apqFowxr7yqbDU1Z1JJACavZwjY5Ar
40Al+HUcYbU8OniP41VMUA==
`protect END_PROTECTED
