`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/cDfTTfbgSXZpVjI2kRUTFtazMPqI99aj8kSCDIujGZ4mw03y/7Au3Lvi2e2I6Df
n/VK1hD1bxry++9o13R7dp9H4jrIm77KMoojlc0+sPE7wpPOT8idmR58Q2QHxRaJ
MU2AGPVrqN6zvwqvkg7FO8UwHCPYtIeoA+2pKbkSeZ1KO7ZmNp3HXDbHsqOEzHp8
KJJ0eJNlsDq4ldX96DR4YxJklSL429WLtYHaYUFTqpRbUrx8SeweXzpUOWUYSRzS
jKp0yMJR7ZuDEansCSi+R+YeN5LVMzfs0Uwyw7TG1jSc/Mbv1CPNExqhlqnu71RJ
Anm+a8tpkklAknMZ0s14WZ88xdRTE8W24P3yKpkOERLAML7CbukriFu4PGjsMsPB
3+CfjS37UKW6f2XSzNPsgD7kKmP6n0sqTYl0Ut3geV+QT8F7DUMWoVM38H0fwdIf
7izvjPPHPjp5ojSb+frgMK4osyfw4zYu/GHvJhTjQQhtH5AWwPmwn++8eHqu3Qmq
jKd4pMuZh8Tw+WRO1dMJTjBu75JfmVCaQkBbLYXBWPFMAZOAOO4Th6fQhskDJfNo
tz/HpANYka/qa0YZZu/eKQ6x/R7bpSJHLk0D1WfVKkBAUYv09p7yG1Za7JIHNGk0
sWMFZ4SVHjx3TJRzvwnjWHwr/Y6PPQod/gz1HTRxJ38tHvu2n5IxjJrJw5bwtYNb
yghH0yZlW8hfzfPoNs5eiNHuJHz0UaiaKRsn3yMs6VjPc0YgRQOGcshLPDdC7XiP
3xK538OSMsxVWYzIcRM5Wkqo4X07b6VXxgNmRWcDuduVibPdjKXaTNKx93H5Ru/y
U9xrqvwRHiwVdHdqh4ZETFMoO1WVvCP5ze+yVLmU7uJ9Rpl089lyK/FynUsAPU/A
7t3hHI9QcbQnNfPd4XIdRvq43RV2xJxL4gXFMKBAkWg/tK971Y50QzjZsNx0l4Hm
k+ZA0kFxCx2Io+e26IYestXiXcopRmcCae/d8/JPDmh4+g5RB8Udk7d1UgcxO6yb
7/q750pPv8fdWNr1dFS9YplbfV41a1Z12hQeT9A8nm8yFu6MyAbL3cxMOoPySJE8
Fk6IgM1xUjY0qwec4r0aXvWXzLc2UE9lwt7It/wDAnk=
`protect END_PROTECTED
