`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WkxpWKNh1EJzgL2J3XIv2YYIs3X71OyW4vdBwuhurEmaNffgJkEUwAmuv9P7iBAy
3JYpNrZfiQa3CnbvM52Sfdo179ajNuu0DWZrq8D8Vr/z2zO62fRbjt0GORwz1f7U
XbTmt1hNIQ+lHPi7s0OKc4bH2unlItQJtQovt/RGqFf7ACEDCVlkd2gyRwqpJfxD
LLqD9/U/4z0iE54u9Uvb/iFm9uSK8gNDTHLo2kLsTtkC1xNIqtyfIym/YrPPGITU
T0JULo60V0AXiHfa4F5OoGmW+7uVRPe4pPHGqf68HwtFsipkCG2htW3ab1kIObVj
tvoTxWEr2ezPTtnPt6u7PR4yhcfb79fx772JYtXGPivNixNdDvrGO9jtJPWRwcDC
`protect END_PROTECTED
