`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kVb5EEOhEX+eiE1NiCB3iwsGK2yEt6BEth81H8t8xK5FDD7KkuXNcMJUre4Bcn5y
gt7q5Zkyq14qQiQl6/ORTpQGMwgpJm15zLehCWQct3ovO76qxdE/HvWQBPc4hT4y
N0TA+q+yTPSuSD1+Uufrlx4v3wYROXVzIjF/PjAEcWNMXK0yUEgLBX3ROl/vXr0V
yy8hV6yyR6jjD/s35R1alM8Io/++BxPpRz76YJmSDAW1y/TtBMwby+OMtpkmBKMP
w6kHslpGgs/Sn1CD2UsP4hW28ITuhVmNVwNAN55bNFN+pZfJpMuTEOaM5HTe9D/v
DQdOB2RwU/IKfvX7wX2IRYOKfx7cSNKGbCC/AGRa64o0cuDNO+yd0QzWRcvc6D6q
krNUAi0dTr/1oy2KXN8L0c6v+FWUqUF+YWNmaTRB4GhGmTniUQxbXGCDwTiasFHK
xZAx8d5gKg/ojPE/dhj4NBe6qS7uMBH5svCp7W2Jp32p0y494Jaas8IHi6okmfuE
8imNLCyMR4RVipTgAqejoqcOKoXdZeVGvonoQ0M6ekDEyYIT+Ib4sE7wGZUW2DJk
tJCsQ44rG/m5IpPxf5xIrAp8TJB3T5cfjOdqNTi3sxxEX1Sm9hu6iHuh7ggZfVcS
eZr3xZS1ClROYQxeeWjItzo1SMBS3E0oXqXFpQ9lFJLg9yGKgKfwx8XTPf3+JR1I
/QxSID2gktk0E0chw07pThv4avDsMJtPR+x0e7bNUZAamAs1FM7lh/yd3iZkdysl
Ul6kt/YEJlYTqoipmWGSBJS1Lfbixb6GxMaJxxt1Vo8e9QPMmomXk4iIDOR0FnNO
ws2glSzcuUMEUJqkxdXopJizqzi93yiJrvDUTjxaTANWrXQBnQD+YWU+DAeNGjX6
3fsYzyn48H1vVmbWrQspcH2Ez3PQNu8kXLpK5iWU1D51Wg6hxXL/pvgECfBsX5xp
chBRxTqgZKSiGM3axbf7iOcaHewHgauKVNNmyLdI8kpgnYAvENDmQ63FosEWHYa+
hwD+83wIJ4zavZq4vzQkjyh59I9Yhy9bNkGzHwPan3Nd8QdZZzRgKbcOqsVLJVEi
u309ejL39i4BuS0HnnB00EmuZ9LqYdrznHttOs82gm4rpcJFBmZKt7tL9cPjDT7A
EeeNkvvWbUeqYR25Rq8uVlc96oBFHyUtLHwvE7Ahkw1PxZoTdqzrhVBGkDlZCw/x
uByZ0P+fremtauCo+5FIiTnatH4tFz3BY6/QHsmlSUS+7ha9+kHgto4it80aBoNv
9HmSOjFsZzvIVtTImih/2lvWiETv3dIzKnKiCoeMc8HJzyT0Xh5QEHK82fPBMSib
fiVCLydPDYZU2d9QmL+ze/8La8hW4dNUy0SkJgiTlWo8e9HiBxMUmtV8fo1bphqn
0alV8igXb9vhYB4+UwZOUNcKV+5CUSsXxbRCISuM7JY/pA3ZoOCzbGjAgpLduG1l
0wnfuMQqDlpLobvf4vGsIEl3HE3DErKSLwN7ghUwq6iDkrTWAYtFWGJ/7yq+cC/e
uZPQpbRHDCkuna601IUsxHPWjSoKJxDTM5S5VkStTpub3c+1L3X+WQzu8qvml2KH
ZMVudZxp501y/ULt4cus9WTNDCsE74JYdU5ApQ5HwSY2jtlcgBA6k2MPvtOmuNdP
dtMO4d1j81w6lTNHkLO2DGk4vtmGzBPDMReYJthP34TKvH1tXLj8z/j3tqoNeSc+
Y9gdpX3DfiDLBtJ//mmjiPosT+gvko1Ki4vxjnvJWzeA3zmXK3cqWfq7rPS4UFRM
szdEp6G3PgoHLDdlM3ukMI54PLEOtoGJzN1IQ10kMTMecMolmfLmUznLeKgBwxF0
eYJrDQ8Eiv4XGhAVLmXDQ83ZKZqwPxa5QONJ9B3gYsS9Qp7PpksGWi3Zze9LgtON
sT5U9lQaYUEbKGeRvDpMFD2dMm3XJ0PXDslDRVUL8Qg9NDCYQ1G9dm1zWN47k0mn
ruK8J4EX+5yhzUWuhwVIiGEupZj/Mti4ug4JKxw/+LNWdv8UStVHIcflLd7WDqPD
JCZZZsnu1CuWsS1yttY+JGKWiL+RmGxzZqGiQ/iY0lMYv3GTflIz/KjuzW+6McZ/
qrAKRzCUTGJjVLt3vix7F74G3F+5PNsQyx3YUMPXP7YDQRVK+abqTyNJsUyo1eLo
Q4BH6n8Acox7CL5IaXLzL7M7NJMXRUDZeBM8Db4eWHAIxkIV0IT0BUWvS28/J6lw
aZOnHuEJXQN1xo6rFTJBDd3TszcoF8Ox+3cWIgFj8HYEd1rlQDCSn4JPYLLC/ZHb
0BQbvXoboklyzRA0kIz7Xq07cfGgMs6nxP0+Qb9oiDTW9PrZ01Y+DkyDuGlnHIzH
vCjMisN3Z702AgCADwGi+rGE5YOFQhVELhlusPqWoMo=
`protect END_PROTECTED
