`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4YgkWhCobg06F587XmnjeZj6obh+1l1/aX7kY8OQnASFsofF7fOe59+4+ofrS9rb
qBb0XR6qQqJAwAV3TTquCtgjJsXQMj67Tx7PnuHb2+ID211xXJe6X/nTkg6+ogM/
XhpUogRCyNz2x8ctMlb3tOOsmvDCIYAMZARieuIUgO4r3mqIoX1p9kZ97txrmwiB
MwzU1sWrWyjMoAcuWaADn3Iv94XR63Nuv8m12k8sWQ5WWBCSITm3Lj6ZO7yNE2mR
pTsM8GY5NLS+V7yTtS4JokJ74eDPPEGCKMlZHCZ73S59gBJS5s6tAje9kbNrv+KH
cKyi8f5KrgTC9WCCUcKDUUiWQDdvFqYze/73HzamtEC6W0mb/qUw6PqjzY44kGa/
VK+WuRpoVVA+s9TzWpcbOhI/obC0dAnWgt4KD4r2v33kWDkZ2o6ZSg4x/JFD/I1k
bRC8AQcgpMLC9SC4jvEw3mg/9+wIo8yegqNCm8btcRdO9dIlTTrjI9bIv/ZkulSk
B2QtA/IZ6QLR6Ay1GEZmKPrk7jzqbE0XIDbmbPyfb5u66qVpqTKLwB5wSy7MO7IT
+VV51FnsRPayRql5+/RC8sbzewEHljZ39KI0gRgYQzA=
`protect END_PROTECTED
