`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DoyyyMmUJVB7oA5gs3fB1NXdWF3T5uvhwmIHIchEO98ukoe5OZjLIPGdimZ/BJw5
gukYVwjKPbcadV6W/9+f0xMIMT7zhNMxl0JnHa0dsbKt48zWD4dkt5iJIDZoYNMt
MLcEhU+PGtzye/pyHBl1UIPYJWmtFzpObcTpVN8iSXStrh6W/NPit5xGsAq10ZBO
p2LbKqPsdvb7xuEstR6lBbxxIa59roF3EadBwaJc3GwIoNP2IhtSTot5Tdo9zytg
QNSmkd+UqjMmeKIfQIKAhZ49qpC20G3i1A31oTKWWRgIQjwpu6BLnWzd6688JMka
Fp5opCrEbSzjZB8QHoNXU6fXPOK9nwHnwDIGAH+uQ1eh2Dy3uM17V9KCIGt3qugA
IxURi5HnUvnuW2A/c9p7PG7eE+RyB9jJujgrl+Q0nA5lJZSkRY6rnezBjPym2P4j
b6Vv9o+KPj1I9YBQnX4p5kta5ujOJJ6FZUctv9H53Eh7YVe0P5kBc8krZ8lzh76A
`protect END_PROTECTED
