`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JQQdRJKAUqpVnIvfxB4EAjCm9OmdBMGnzhZNPuP+/iSEaa0kRRJQQDmae5gpUcv
bcuRCugEfRdRHDW0eCTGDt6HNnEGnHAp31+NNd3noI0gWtKom/gYMicg/R+1xltp
s7lOP0HSt56pmslCn/4QjZan7KnH1o2wa73ZxhFwPhTjXQVa+lOvXgryGEXV5FmV
IRfbSOjvMbIC4wMNqppNXDHh+dphKkaHbe6mj3n7FRuQrW68BNUbdDWcFypz3lsj
w7fZql5xuiWqsYKFTzfsrQjzqfyJqjYgtJqq9CmaxiYUZPFotl31NO53ZugQnsbf
iR2RW5Bc/fyw52T/3TWNw38ndEHGgpelwvWZnqv/GYfdUx+78VcgTBT8znJZjkeP
7masfrjEutl0btGwRCnjNNAuqYlJzfNAPAKcT5G9W7LpJ4P2jEiIHm/IJN/b52Zu
17USxy524xsXKmWOD6LityTIxPXLYd6D5Nqr9+LZEhGGTn45FgLbM0o1+OfH7zWU
YvoNLv/2qtcnFaRaGv8jX5/U+ZLfNPfB0tVrw5cwaJwVKzhwxZ8urFTT7i01kUU6
Em1C7/qLFbfkxgpZEPZqk3dItbCBOeZz2/ewNq0zbXUxlgeAD3P5aeUWIGDZNGho
b5EO7jT5eaHWcAF7znbbeQ==
`protect END_PROTECTED
