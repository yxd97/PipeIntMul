`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y175AaMcoenMEAlDZhzmAgtM3RB2mNW9Skz2yx72i6rKYGEDbwaXOQYP87YALNwN
KZSFLoq91DVWlMKaZaXNmjomkQTkCWiKrIMYRF4wTJZlrMAJcUjwk7r/nY8CzwU/
stYaq/dDPOa3k0j4cKiJ7XAHpeqjrHER/awRrjmg5g7hlHkVnh4nqnh+r/+AjD0F
3xhmHode1uHNRw1+E86TmzovLg3+hNiONlUU4RCDOv7wbJ1zBcllPsz+TvUXJo3H
0HYufDc5BpVySfrl9HGT9bdEABd47rZRjfU1iBrL7KWkxEDcF6pELrQJ1Y1dhiqT
OkQDIPRsAdA0D57I/s3xBqCGmHEDFy1wUGYLln0O5H3VtRvzwn19IHMAaKWpY+9F
tIqNbWaRkPcc3EppT/HXnsmLW/uZmG+lyir08OdMgCJecKIw1RPZqQRiVwCPiNKQ
`protect END_PROTECTED
