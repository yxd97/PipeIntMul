`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xOIB4Jqah9uYsMxJHRPw1CNZitDxZzR/y71k6rBtKwMZ3oNWGdmyn7b0xjalTWkz
I8t/8Q43XNCqYyVmdF5ebB4UatHZmiIkHlQDuXZR36zO+6wXfltR+V97/yKiDKIH
sRltu1F52Vmgl9APENw5wk20gg4Kpi8gFy+L6D79bfbvvrmNYCc42RxySRdOPMJx
jy1qNexh217bknvb9sggIHqzZyb+s43HljZ6riJdm8PCVJFeapPloW+DqRFgaqSF
`protect END_PROTECTED
