`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/RCJDrrZHwIlU+VFIbAYFq1u/JtSjnAMLlBqR9SOp7vsSKRfC760scxNQO+FgOox
1w0VfRQjw4nKDwVxVqN8zXfKDfTxqgsWReFiZy6z/2dFXSwYnL/iLACYq784w4wV
v6hY8GFF/RqVs2iZmCl7nhah2TdHJS4d9eHr0Qk9PljmwRpvn9ATIDIV86WToNeU
AFa0ej3b5F9UWml+IuxaoaBclAsTumARMrIt2sQXf/A9sG5/4ODEtvwGoLpSYqCM
BZuzw/91zO7LHF0rGkeuBgCbFwMc2uFw8eYPiXxDZHFPKrr9DLtLSic6PfimmB5U
696iG7btNepzr3nfo8poSiw6FIngACU9EACAZMVHH6h3NdhL2dPHyLJIKCAeBsvQ
Ua6G9HfevxS2k2WU6M+3+4qPnNt3dC6N7FRpJOUcTA8IhCpnJfiaVD4XSkF04XmO
WAdz3g6v/FFJNKEGMIECB/7rnl5AebLAyLa3ga99M26h35+qsoqciopI/rlo9/xz
1Oycng0ZLt8nv8LtRwMbFQ==
`protect END_PROTECTED
