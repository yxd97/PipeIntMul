`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bZSF1kqBcV1QGlGmWVS+TA4E4HZY2LSprAqFTMtAn6lz6Cm78ieg6PPskAwNhvCd
8ELjnIblHFO+kUIv2yYRK3s2czOcAaLaP2koE0vmmGb2T2biBGc9bfhnqHjeg+Th
q9h9LgK6/EKFqEzk/LxiUjrIp7cFvqwgJn143P2hR0gLB6t6kYa3eZv9YH7oUlI7
+BnnkWJ5+PwHgI/WGlwZ06nnwGmhE3bjy0XSwa8JIVHfjThnQ+W4zVYkOihSFOeW
5OyMOyrxjsCesuz3+mO6rjPAujxxQci2p3thsPUJ3FCwGCuUmhMdFajyzJim5ls5
WJ7teNnuN4Bmy2/uACm9ib/SNvR5d8IREpU2SZCPtM6Coocl+JPTbq3FTHvN69j1
TsqWruendCwdNgzXMgwVxINGlBGNjk7waS/U+gCbgNtsCvfsu4g5XCal+3CWGdHU
DP9evXqJPP/t7+gYEjaRxVq9asFufhjURs8JyfcFweci+dCc0//BzzhXCA2bpQBL
Vsx50EFNrGB1CahSzs95dYKrZQKSkvk1m5frAeMTTta5mZGyXpazxZFSVpSwBnJA
2TooD70HjxLMGEH8hPprELljVwKfHh5HJ6vy03mgAgsTo+US9BShuDb21UhJGBEm
R9ZRb0K2JosopuW3LNyO4rN9p6WPbTZx2lmLu7q/Qv6JQpop8IyPvqf1rANOKnE/
qNXwEqzZeXfRna/nimUCEJi6uOyxiqy2tI05QcTFTZbmoBDjg9JzRXERKQWy5ZAT
kPz2mhH8m46hrdYMoLXmdz4at5MLvDPC+nkoxH3jCc5xSLQ3/x7GJe2S65t9rdZL
TbtsEjiIjvbJFkHRkW2ThqXPOTbGQDosVuz7eWSH6LtWxMuooeyg/5wNv5lLPVMb
+KtTVsyiWOXFaQ9Pw8pK2oWWP5s+cdJrQuZzl2Ma27k1VUfS+fnCHLlfcL4Y4Jq6
mHVnffL9qSVt6nxYnFFupLueQtXfHru3xvgQvNtc3TmM/DhGYHyQEVzCNQuzPtZ3
ClzM8sdgJiVskY+C0h4ZIjDqVKvtiP62mJEIMWjPri+I0puM+o1OLyt4UAmI5eJ4
3JrZjV26G7AXVoXL+1Eg0CA6oXV0kDMr03gOLfILd0W6xftX2PUZGe1K65q99t02
J9vX8BROxo+M3GF7nzBx91DOPi/8vo6Szem7DmYanzEpXD3RLttQRG51o0YEwmLR
vhejbR7POV2OidD8V3LEgWxGOmYIAw1vEemH+iNWRD8st+cbJ0fvqHuzl3g/vJdX
1ykQpPkKU8NK9vfQAadnopWUTqkpjQs6Pqbm4KZzunW6xLfnpl6juyTW9MnlIhBd
L9zwwDiqnWypBA6ZKC2y/T7FdsgNhAyKn2qwTePn3TB9QTu2cK1b4UAMliSdon5V
gJZ3AgHNyZOSjekadjqBKeedOsCgw3TATtUlDCScPNDqAXSxvE7MMz111eRdygfz
1X0HCXBSW6S5Y5oIXGLyERfa+KIYw5QbvC3k1Nsys636uOeMMbkWXQGDGgT3LOGj
nNYlUNrSXrVLacTLWsAGvlFZO4l1PGThD9suyjhCpP+7B4SkKfMNPdunAKTAS9fi
IMLipZx9xvcFeJOR0nDJqgenBV6iYvWSMWe7d1drL5b2+WJUVqrJBUdXGYeo+sIl
jEzld/DeuF37XUaz6bdERYtwRIq/JjwI5wBwAwbY+TLBeLnn2V1OJz7iHfczxOqD
M8bPZ69oJDt30emviPz+6V51SKOxFSnn7LxP9/dgdxf4Ha+wuc5RaGadLjkfyzuA
tU0kS48tTgG+RsUpLRrFS508mnLU4YDjsD/djoOyW1L/2Vd1J6FVzMxdwJBTWUi8
w1nvjv49+IpwbEh6wVuyeZLrKpEBuqO0LriAXVSpgnPzoCzt2kH14gGBWuDlvOiS
jSiBW02BX5Hh1flQDoTTtU8EPgngxRBXocnxT3ZnnosXqJNNA0ZvdoQL+NhcTt22
PY26KUMJeJfqGonQIU8kUy8ARj0GJo9mfhvremCRgYX74glRyOpErfQKFkt0+uQ/
A8dS/kDzqOomuIXx/E8Aew==
`protect END_PROTECTED
