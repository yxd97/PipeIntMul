`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nUNIMWC7FPHdo5uIfxl3X+CPY5CHejTTE5Tt0k3D94qgVX5123+6Qym3ErPzKKVp
a2j77ktFejbRzo/IpkT1glHm676IsHpdXAs99oJ54GA5TgYI3lITW/cQpIk5oA8Q
bfxhJ2aob8i39PvcGhf6R+BZI0nmV+pZL61HdL63oAltrc/iuqpFoM3k0eupihwP
nPr0EN/9PavX5SfHP3JvGBbyvKyzZiQyWSO4vg2gTtcn0QFO6DEcIcCiE7J05OH7
fq6z3arlKeB5U/xiUW11oxHOe1IJBzsQUgT+SURohzkqbigBPIIz8YlrGKrqdZXH
92ZT2cnmjEwzkX98IlCKMsxDUv/Pbq0X+Et6Ee9EPWajhOgT8lTo8HcWjgIUbliM
Jbeqz+yQAfi4p88y+bcx9v5Qmx/dqMxEJL7P/5a5D6wQ+6NJgpJN3gw7qxgZHg+q
DfTGP7xKjOhkPPM8qod7+uolCF2xbzeCIrDSaNOeWRs8g8v8x/dMAzvE4bFFFeOY
JwJIEgHU04xQ3EoqWOsbun1jRnF7TF6Ku8dWXjprTpyYu09DJYyvtY+XMfaG+Mo5
7KEeHKLfvgDY0HxYsOU87skUU4pspXVhYZjBzF8WyQjtCsjDIui9Pg2qsp9Fox++
qmEoPA4ycLfFGN8q9ngkSPJ2YDJbh5iv6yZb8HxbvClVncmmv7lvR573XLdC9Z1y
R5OBsTdToLOOsG3QfgRbUvbwPRe8G6hxbDz6KsHEiVqeuAaDkitpvlyOasw/fOn3
+RU8gDlOheIR+sICAMR/leKlIAoSeLqKzo+D2ZFLMRbqAVo75B7/rs2KIV0APy84
6JVdLmIZN1Qtk7WrEi+JBGR3LSbc7GdfsCxwzKe+KL+00F149AXjMwhV/j8u2gW+
jZ08xs2mO6THWV2csg6Fr1CXFse+MoSQuBcJU7iqKsh5oq8AodoVhy/aCA+Tg3u4
SKZLy1e2Li25E9oVwVGIA7DFDNTTzZNWL6OZ8NDoXVks/S3EDg9CpRSm7mJHsjGP
4Tkox3A0CiIaohXZ0J9tTe/8nn0yUzSuqcrQl5hXw4rbWE0AhIpGNC6qgvydVJTw
hgUKSPiu1dZKWnUEJS1J7zkt6BRUKZa2owenIm/IfvhikwS1DL0ybRQwt6Xf9P6T
1korOY3F5v4JYd7vz0xgMBzKqprx+2RP+OUte5K8UwJkugFuDBr9wY/kBZskgFlJ
pgsi3PEfa+jjPNmWgOZykKBb8Wr7ksfLlTxI1yYQB8yZJiS6tnbVaL7HkqnfcHTX
pKGaSCTaC/MqLkadN3xA/U4Be/XmLTmK2pRGBDAn6SNCE4dWk4zgBVThmjLKDSVz
RDc5wcyuE8WDR/O3iwj6JRTtSxCOIIIBy3WWhV70G5MqdAm8yzD2HG72iXldyKda
DLpcU6B74yw/2tRVGuWcI0M++VXYXUZZYIvMWUivRAcdG9NV6eIpFim/7pKn+bY6
r0+ZZhSWgrfueVwxF/pTKy1wM4lizBvWc4rGcl0nZ4w6kCC2sNZ+1MyJhFDwBpzw
e6Gj5ybNRGeiS5ACJujFNp6CopOUbgAND4U7M1oNZkcRDsdeqYolAau8HMTeDsUz
Hd6y6PNYEazd8yQkIziYRUX65WUHVK3xI8BxJnLWDPZu8a1i0Agjfb6MlRz4zHfO
TJfJ6QZwnt8xWL++/qDoi4BKndLgKlcaVgMbgzsh4Ct9h6tqxv+CGAaVymIUjzaL
Kd0GtEDTnXUyDro0MefBCFYv2GbMWzxqDIsa0D5l2ow37rh1AUBNDqslD64e69UZ
jeSduTQPjSndHDH7HY8QgyfaZUM2FJJxUYrjv43AGh2AZX3TAJDu6QJrDgMT7qtl
Wk934ttJk6ChzFaHTIrAEmweoXFV/7onkhbGJnyy4RbHJw2h3H5KrNNIHqQ1+6GE
SCqHWDUl9/pSM7ZlZZEP/eou/h5qH8oYZp7F9S3i1SoL6vWN9MnCpQK6gjfcmPqM
MmA41NMJL2Zp3xbpLyMerMpA2WNgsMbOVO25U6U6gtRLbwRxKTf9VtrCwLNiLo63
2gadEa5ScAj4g/dFNio4jMHQDlGPmnWxtlxor1qdIHvWFVA+Qn6qnV0dLR5BWEZc
7Qe6bAmADGZUfNJkK1SFWQfly2b57iGeKH/2mChJzygCSgb24E8ZTMO0My5KcZKB
6O9Y5eQjT354HlOLJ1c1+MmDLhkkAicOLtKBZfE7VD/hkO3LmuBRG5upeKl7g9Vp
pDwq1Q2P4LbuUCetENL4/AtRktgd45pNtJ8QZB6hnabtm3+6VZ/szQaf6D57qesn
znIzsa9AKn2Bosh3lbr0BHpiM38pagNojPllejpTIfA2ZLFs5KTTwaecD1Pp/ILO
k+hSRzuKIg/Mad0B7zJqpt3qgPPe4MaZRReVWTKWUgjNxgTx9p9TNrpw4AJTfllh
Jkg1QRkfS3WIRLjtiURSJ0c9+hkKo/PWFVpVc5k4Gj0qG0SPcw1DmfdD+Re02kp9
wXxqX2PTQURHHlZzsS9PzOuXK8fxAHUU6rMaiqISDtK1QaNa+zI51Yk5oXBE76S0
GHpTD0/jXsYgs8ynpbd4xIFusxjVzKFK8othlkZbx007iONbfD67tz3CMxCucXZb
GvYNTdj4uUv7E8rZLUSWLJeqJl+7ZoNHWDtzQHBbAEvK24cu+AXaSW7U2VfGDG+1
jJgpiOaIpcPDdJgTiUyuWc4CDm+v7f/SUKHxmqpSBW3pPy+4n/Ogc+mWSG3E+Ktj
h+N6rdjbNk19DhMp2RysTpoDRmh7elNsHyF2zEjIsdxqjGHii0eWTc8nO8v/NMxP
OXYwrxszT21B66zgv8S71McutRBfC77/+xFfsrXMs/VOTKcDqQQDDuFJPhVmNYYu
Lxll9UzcuymaUwru76S83gmXb/S6GFRz/VihKRBXXMMEHhQ88Q3yJRyvv3fSe3NI
bd7oKMIHHgvHWb8OgFwoyiuEsWcMTp3r9prgJ0B5X8M=
`protect END_PROTECTED
