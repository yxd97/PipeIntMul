`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jsue5v1DpK+tt5x+xPa5lYiLisuXdRXYELFGW1CONDd6d9KRigvzPQfrt826srkg
QbKjYOQmYNXHllRUYJRX5DhhM1HgFc7HV8ICuyXYuU/AEuFjdVsrLzN/gSb8XIOX
6lARIzbkrSAAUAAbd+/V6wFupkyYi7buYa4J03WNAbUAnQ0nLtmo7rrukT+tbJXS
Q0YhkG3f9KP3/0dpi0OPz8fFIj6iD2LN0boIQ6gcD5dsmC+Zi9cP7ESOeLCiKjdh
u5NcfBEvrHiYIRySzYxixeueW3xkGjp0vqHfLeK3kE2ke8uyH6x27VQ6/RssjSjb
ZsS91HZl0zgpFn84hUs4TwIaBoDPfoXYSsOl4FcfmLi0veQoFoGgTlznbTYq8UPc
h6+OJwwyrUp39tGUMreOm1yHdaMqzNn7bb/UO5JtD66WE3swVkj2iWcc62hXQYm3
zrrJqumQtJB1jyF69m0MAA5N2sSovJJmHuTWO65R+XAsgEXIGI4yr6sTPJd3S2u2
XrqZ53WpzN2yaeD4QuUUbZXJSiwQzwvi6pubjNaf6f3MU0F8wYAjZuiQUCo3Opdx
K8dgsTKk9WaQysMayHW5JaTWENZjHPcR5TGCEMpqq44=
`protect END_PROTECTED
