`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
euoXrScJ7fMIDcKgb7uMDVGRnGMBAtyMHWwWyc1bTffE1QV+mo3ImkfCTABIVxGb
Tp1A/B37gKvnr31aDW8fqlo9vPzmEC1+4eXjY/e8yBmKdpeULNE1Hor4zlecAs/7
2m7coBsd/XW0L+6DHCe8m6wDOTo/YOz9pHX8DWmAd+4oEUE1UsxWc0y9QpxdeSGI
xrwhcS8xljJvZT0TZd3RlPijddhNGzAmhPnZNa3Ddzie/mmuT8hXz7VrYdBjDjVN
bcQUn3QX2934pAYYzpK01W5tDGbVazR9vmU6h/ywiuDOTqVHX5lA1gFnU2YlPdl4
8QgPBB9zjW+yYQGcOOzjuAN/O9hRFVZsIdYxG67kwzwRCM+FRlxO6TwfoNbufcMc
eAwY/vvzkHkQnxRtAc9/Y4ddNKjLVJJ7WiBuW47Bm24gB/qeYTCW6LVriGOL0dz/
5FqpCGLLa+QEE+uAZ3H6QMlUNngPEXYSp/PCVjQWwCG29D/lE5wkX2GyU+YHYG/j
6512Y/FMhmZqd0IjmodSSySNk2ChIGaTWZG1d5nUcw8NTB9cUvZTuwHn0ncgyzp3
tL1Mp+/3HfwSgvZ/JpLeAMeReMflIQUGjfQM3wvO87q+Azwpshj+dWgURKaOuRlB
pTxry90tzsgwBaXQkCAp8GBY7l/EQXPqm0ULPXyHeR+dTNrzDrOO4eoP1OzK+Vu2
N8hz1rXWEaj8VN8VB6DZR7VLWps48DMw99vvgC2xrfu6arkKmBzPBk16l18bF3uo
y1S74vzsRgPwIP6orYa79N8zMMYCD1YsBg5uhmABv/tZaiDsbR4eLSm1pep7jCFH
BBad1rusI/8QVL73Q8pI7Q==
`protect END_PROTECTED
