`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zTbiFWSuwXzIHdp5bkTuFu7/FKuRf7W29fwv1/lvN7gcckwCqq5BZrCnUiLC3dPc
lpysYyNTVLuCcDRqXBx1z5vWFsPZ3aC85ko4xwDP46cQQCKQbA6dFSiizw9ba3TK
rFa6RnG7B89XIN31Icna//enkAA5eduJBIW8vJW7iRQMHOLeRQmwTwEjEiGeAp3X
1XALTjIrg0Ah6sOJAEVU75hqUjMAPlpa2etVxJiP1daVDkJtCro5k+GotIXPnmpa
OyYyE3vGJKP4p7erD8cObGczJdqIdfMAb3Dqb8Ou42A=
`protect END_PROTECTED
