`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uMtmUz2PaJ5JgyimIZxmFI6hM52KSHz3R4tBSBiys6rxzOKjpEuuj/MlzHIZCXct
HJkuI5cLEzJ2MinbbxnzDLeHkJuv/fGzdevlgH+FvwnAn8KQ15BTiJ/RHuAQ+23F
SE/zwf+oWnB4T5OtIDzKk6a4C86p8kXSAzV3txqvu2o5QlQIsKrpbrRsYpZ2+tvn
vrhe/2bqtzQCcKio2sp5yUNqJNhkzzS1cMxcd/XdBNISKVYEO0aZBm+cYlyf+P6j
0TI7XieTsciVPZbXR/8fFMiLMPE/LfPBOgSWb6WZ+PmEL9zS5BEax4X+JsT8nsov
YJ2AsrWgNWHDtUnp7pbJV46fGidy+LSUfmWQVho7VNZOj7Aji6wqA7hwDmJnAf8N
e2mfXaZaLuAQlvgMxWn3+TDgcRNe4aNt54lNRPxrqTTyhSJzG5k3jhXoKWWeogzq
v9zE3qPlEUpr4bFewvpWrws3XJyWpKaWmq/Y0xybVq58pravVDbWlBWvLsbk1skv
p7tE/VIBJyA7+SNU15234wlNUBxyWLYQmhB3O+4mWrra5UAqpSrVt9YMqfjr7BW6
5vfJAnwhHvDPYXsZy+eBVoTQdgl3S8vc+W4MWWc5nasGeS0d8BZsNR8ybUcmpWCk
0Bls/NjmJU69Rw+AoLULHFUyCe3pznBSINrj8vK9U59GyXfv+kLWZeJoxq7BWAbB
3XRAwyYvujGvS58IkiBIDlIZEyD16TZDuotgHsae389eACV6EvrujImyJUi9DZn0
3VvHiZBMWGCnkCSMxT5KrgsaM2GrhxypuksNz6LByB0vT2DqCH6p8kNAA91/jbx5
2x1BwZ8A9HZKGa/c6YUjLOS8tREj96mj6oeghd8Sy5shP9XyJP67a+mmaPRP+zK/
jAImacYk7bGy0NtQrkFAF0vS7yCBHUh1+Zzpsp2KjsT9t0V6VXOb8+TtZSmzOHk3
AZV9fSpntv3ZHhV+cQ+hZiQhp6oVqzWnBwBAnINXJe5VO81uEK7allAvtPj+7s0l
wCooN+o+OigDBS1hC9fBECRQXpj2nwApcVkBtDOkHoBAJdG5SfGl6CICu241/bub
HMlque8ESYQvJGq3hGflHBNftkPVJM3sxIvYiiBWgdJ22Jf8LeUgtJOy/yW2KUFE
nSFBnctE3Zr1Kk9yXU/K57NYbmnbF5PFu0AtbABQ9LeZV+Bb9drZD7jtZVrAYJVA
wR6WpQja7iEbN5LUjw5aqnoOeFCyxhg5FlgMV6CC9pj0sXYMi1li+kADKy2jtmmu
sQH132/r1RnzebpQ+eOVWfhyJBg2Micc8jZJYBIE0E5A1GqbSqXgJSZcad/mF5Fk
VJHHo4Xj3OgHTo0kufIEAqzgqoDD6x1pRtYqrqkyHNC3Siz7j1X848n+hrQ+mh5K
dakvawQL7m0FkuiNVKoBtjvL0maKEn/d09JID1aiBb0SmMBShZIrp0aUUXAvs6VB
0T+h4VJYzq3Js2xKu/9qs/P/mZVPWgD4NFs1OCKcPlKa7yeVvW/KIKriNHZ6t8NV
j4mn3mx+XXImA8qctQk0ptAwNfR1CW9xyWvgV5l2uoYKnKtTZOBD8O3bsUGvTejV
AktjZ25QYHuWD7YBOZAZCu26TzocxQFV5C09dQTTWOHHb23Rg/Tdtqm8qC1o0unp
T9nqtVcpYhBbNyhDF0SiMCut1om4WAdr4LvjXnC55BknAf++dvZd2HcjuT5NBkRY
tlsC9Y/88qzHjCnt9BxIYQQwXcDK4h6dP3kRtdCEfoSsyQJbLc/csdpVMSXb9iVS
cyeAllE6pIjkKxmE+HWZdEZzSqOIb5xisg3YlPxo1Lzdjix6tav/A+8RETIu0fZD
IYM4jJEK30l5OcduIKhKHaIAt1h9JyAIdzirnOJzKvVpjL7W3ak7s2oz3oMEMV7c
7N1LSCb0jLbyDNxN4iAKHykuchJf/gxvbQI8mPCEOY/v9v+msNmlB359pamhrSkU
SdJFbd4uE2mqDrVNGPIDrl/uyfEVXOUQ6itlZ7nVovv0WCiHqgmFFAU8p93unJWz
eIUCLQAKUQLo/iqu0VBOdtXnwISUEUqVo/O7SaFyulGoLuP0moUcT1aKHF6Vn6gV
EMUiCm8McaQSTvbdBvIZycXxr+OjRIUjSRi4rGEpvuxWQ/EveKLxR/7DGOFuyBEE
WIUz/i841cEx1qH78DGaRIvMXIACT2rCZj/a8ReGXAEvYE8g5j9p0/EU0Gi9eJMX
i6uaWysWYVmmzvCya/ubpIcncIwXShVctA3/vjfW13LKIb0rA9GEpdpM5ey/HDox
LRHTCQdIF5RbiY9WCZnkqpTtYO75qCZsToG+wSPDfkzRezSfaCU7CWsM+hdqEXMe
rDUr+6apN9m/eD93IHVRF4+PMh0T2zVF5SHun5GSKt7PNwvaMlcB2WOuoIL5BBfJ
0+xqNEjYBxb87Nxo+3tZaAzncIRKswDwVumlml8F8IUvJAHJ/idS09EcL0+uPhbB
o74FyG5d/vtW9za4si9Tz7NSlynG82LXnb8u8jIMHYJ8OZ/eR+NtlVEa9saXnmLa
4dqIcyNV/sv9HnR2PpknXD3yx1IYw/6ocwx+Bvf52qCCsTW/hF+gOl1XKQhJJjsd
iqdpUZhioKqlwrddqGf6qUGdB8w1nSKC493b/lifKgYfapUHAuHIiTV1nf91WzsZ
ZnaVcdd7+yfDTSKepJ+3DHcBm0wreYIFGICs12cmJT2vwY0G/JBRMBrFNVX77fUD
nTgbqILAX+P8ZXqMsMAQqiqiXAGb5BnjpSo/sLo2RZV2p8QuNYhnW5CL8M9EjaJj
9GH3fNO3kLBYZPqvYIVMOT2ICPEhXoP7HA2NTXHtWe79AkSWA6f7k0xcTuhLImCd
tq07v2VauDDsNW8ckOlQ6gWu4cuKOMK2PBRPDK9C3xuUvGzSSuHYUHObvtIfL3RN
Khemy0TeBAXBtB5EHmQ2utn0bkwBQomtPvKgGhScdZHxT6GAQkxO4BustfVjIKtT
jdg+QzNDCeQSXUQXylFXNZ0AC3uzrTQ9mDM9sqESZAQqcBm6TfGAN+d3ZP3Rjd3e
Ta9So65uTDApaOfY5tV3eQHDJfjHhZRK0ssyUtlyMwW52yNYlEnfwrzPuLFGEmug
ta+micifCaQynZpOIh5ZPAiXNHaGlN2KxdZ/kCNskRohV6OlHOrsYOgj5R6Thb5h
xdMH2cuThyRPF7zL0mQj+o3Rfn/JQWMBFaJJwzvM2b/hWmosN8I7Nt8tGyzKqDhD
GC8yt6n85UUpjc9i8vaRlZaHfY2sDNQ9sYneDGcwIVRRJ41Z0/szPKYWDV7EZc9O
LIjYO4uwJCnlvu5tylNyy/A3IZ89TSoJdrSsgjAknakAB+Vr1OjdNTMbgu0EO3hA
wMGVQNvKtoTugTx1LExlkIVuiz38PS9N/o+k071AtiSPm2WnEAOLyzlTG2NGVN+B
EPO4LPeoQCEfDEdAYccXKan1bpzP0n7IWiqoTj2lmMU=
`protect END_PROTECTED
