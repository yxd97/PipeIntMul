`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nA4wr1GJ9me2nSNDUr8Ukix0P/LNMAwKWWFH7pB/rOxKyNvreyrwJY6inmfxPcJo
s6ojewppnymaqzgHkAHe19UwbgA4rubWqlu/rt1x7smp357RhFYxyPaBKkeO+gMz
QeG7m2GrRZKtvLqEABmz2ZdKJdiEcxkuI8Xs3TIZ3ej10UOTf+f4xtMes9xYqOt4
wJuCAXhoUcO0NgufzzejGAIY5PeUJJcK0JrfVZdpznPoInedof/rgs6/pRj969W0
bDY1N3dJv6raCdG8BGd7FI/s5wyoDn20QvOm1kji7dDE5W6bVFGVliU15tnNqptg
tdyun8dLbdp/wLpkgh7VKCSom3jRNbs91eQ++MMs2HegeR3SP33i7ciu4aq1ekij
GZX08fynt4fQTPmgiTCPQVr/YbDwMc9IJVdofLST1WE=
`protect END_PROTECTED
