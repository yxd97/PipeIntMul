`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TJaK2WZv6jSP0CfdwLGcWbHlju4bssfTYn2e21DbnPk8LSsgtldXb2ETog+cCwX1
fuHiy7MKt71RGjH4G0WLlXgo06kY96UAcqz5nBItYRrV1Svxbwzfr85T7vn4p80B
bbeBHHOTYrtx9g6XzY3UJaLSoK180MeKGCIcXRqbdqBXDw5K/5WMSCTx4O6bNqLo
Gi8DDMpSqDn8ZWewWfuYIKI/jKviS5ae4AR/d5JC/T6FkXLky+mVkKMQuzRc3qJn
MkxaF/IPcarbaex9D0Ca+cEeFtWQKRAYO6oDyvx746MC5n7I0fIUatHMrgs9VBrf
rJjHLaK+inW9KhpiMS7LKdV8QZhKCoc6Rf2j3E5lQtYJe5GLff+anXI94Ioc+9Mp
2F5fXzl0+IFCmj3qC20UW5hMVwRstOp2TVRfderkKNeOXNknbk7MiHZqNWKAAAYo
NdEtWSWek8rQmNEb28yEKmvaDEyVkXDXKlW8yyKM2YQsKVgKXK8Ty2DPf7iF0+BU
0kP8UL8BQpaWBkxxaGhyUr5iRY0Q9d9KIY2MeBFNjH1X0L0ZUMBKlKR8uAg4uV2r
rAoERjN1zbpKKzQTevmDYWs+NWjDvqN/8FBEhzItAyHkGLaTvOlt6U3pWZvDpnlO
UhViUuJOX/BKM3t6Nng2rr3yjGjSms8mzxcI6bM48d+ewiy3l8p6Ax5bzGzwRx8v
AgzZxcmXzu/JxhGLOXDhxXQDOntnuDak2FzyKsdjttrcAZ12ILNW6HHeT1vBnlXH
GRnCUjMwvEOm+Vmv6BIV/lME8FeF9Mia4zKkBPR0CUZW+J5aN2ztcNnZrn5vrfFL
luGLWkPjnVmv4juhVrCbGx7AM2t5euzU36NvgiO15FTiLljUjBmFf46hC3RWzi/1
FS/ZUJiIj/nAMn8AfXmKuY3ANSnsbf1dQE2ryDwZkfZdLlLBIm5TB/SxQD0kHos3
jqOB5jE9J+nEGX7BWd5+Xe2EIV+EF4An2yBOR9B0rwtJHNyG8GpefV4hO2ylXcNb
w3rOX7uHzky2K/pxSnLuqo50MPV9zn0L7JTZF/ZM02IPiYahKTCNtpzmkOr9cOje
dyJdDrbNFA51/N11G0uOAVpHTBp4cO4u90ok/p+cSSgnTcbFxW9GJ6RfoZ1Dirco
Mb6IIFDwyD8gZyaUXOQ82aN+UjT9t9CoCWS1sNKOgN/Ge/ZF/eYlhbyTFeRrOY8S
iicHgFDeKZCxDt25WtHNKZAkCV3iWMU0ej8wghJDnPsAU0v8AvNkRI+j/8J290TW
9sLx7gNBuWAhQrSt+lcSVMVo8ftOOM/hZJUCSZ7JYGvCcEZxR8T+OrYMwDX/OpSH
vWcH+hIGU0082PyQXs0FJWhov5J+VWjzxbhf3XUlwcf/s370I5y5XdsFIqU8wsBu
lSQt1vfNaN0nplkXzgxohoirK++GWBnKkV3CjLeqB9nzHfI82DCITbf7gtVABUVG
cCnbDOUT0EIELoq7XZZ6pd+ql2Vn9jYqV7auJ7XAWJjiju5lTIuHGmc6nGGEnuq6
xjW/akFOntxtOGpM4nKF1WYSBh90UX8WBNdDFDVjbmulov9pN4666LETd50ASqJx
9JOvEwBqqAXT9ojjgydGJ1Wi9IUvkvxQNMFmf6tZA8yMDRzX/Hvgrid9Ab9Oq2tB
Id900Fr6emfpzty3wJCZDHX5okgBmaD9mOEQygGnoiNwWTm87LYEXAr/cAUrmAF+
maqjb9plVZDasCIS0LZZojSFKpIWeADDBxyQYJ9siT18kLDzAC4TSgO00JNrjfrx
6fg/izrnONTWSpInmkaxTkPveMUYZ+84+reyxOerWZWd7OgaAVh76DoIPeofXm2m
Gn+IuJxa2il6cvz6QRiHq44e4S9zACTjhT2wGA4r7ga3HxADg/BEyfiU2hWB9XZa
hQ6uv62/xu2yDai0fbgJqC9cmOyCZ4EzpO9DBvGfXI8ml0IABO6piuIQ1bNyCU7y
0u4W4Mw4Cq81nt071RIM7jCXC+VvMOqP4Q85sf8Mav8e2gokzWflrSEfoSV+fijU
qvKW7epevmIQVyRor8nKTofbL+4FtyKaGROYcw3nzYq2ZKAsIgb3ALaQGKammoBQ
7wD3H9xyEy8F0HDdbu299IhyicBV9ITcdPtt9ueh1EuHApt7f/oOui76fbonKkiw
wiH8GQJKAeQi5RV2AzYnVRjg0dL/Iy69bBclqg3TJyTGENS4xUe6xunVIrsPMCF7
vquYYku9sZXtToAjPmv+YeEWKKjb1/DKgGt44Xwx8tiidAAxQ5HizNJQqc7RP58/
Jm+9oEmyMjDh0mMi3zVWMeXUIDU8MRgdjDVgIu56t2ZInOJQ6+DHvX2WRwlsgw+Z
vcS40bssBqHZSfW6eh5wugoVoQrIgAIh6aGqdWYNaRNAwJnUs6UIjo9s1fW+Ol1P
qM3lGoRRrS4aNJcSD/MEgCJC002eSIWAi74krA6uwUuN8oV20Rsz2NjLZSawsr89
04fr5II/pthm+8xDgvfWlHlv46iCPEflaDCJka1Hl/r17PYEKGwJ6SOJ7g7XQPHp
jDkP2USV6MG5bo0i6c2XBoMN/FUE+o4wjEsybuUka9X0EhmicLDDzdL+AdGrgxA+
48MUGRQafpqUskgYnkvCszsIMV1VmpVkAKTBK27kO8yWNjarF4Usm6sqiYIlpgaB
BC6O/sfo7LPgiC0GEAVb7oHgkhvHp3QMSfE7tl8OvxISM8K6Yu536wivZf4Tzx3C
IiqQEfsvDknCoYTdBuKhL9FMrt5ZULKAL7CbKLfB6Uag75IHpKrfVpWWNKcCinHS
xa7VvT+R444pL6zb1WTjHNNtR/a6BeTJZH/PmQEgAwXzoT8dMFdFMC60pamWOa3L
/msuEw1RpD5cOlrajhwlUJLf9ZXesIjW47AD+CpGkUtUlQ1DsVgDY5wPf6WtV8lk
+Et4jAyvrXKNB1S6a9iMnXOmJXA97MuPBaNrDJomVG5qTMc+WaHsdqahhUgkXTO7
BWndr9FJ5kDJYehWpEnIpZMINRa0inRnHr3z1e3vCPwa4joppHrg8f+Gry2PZY0+
+Tlg2kJxhBnk6xB9nsDLyy1XrijhDElnhj8qS46kLhkElBfh/ZL/ibeNKS7HhFqE
e1dS6hmJBmWqzq57Q2v66QgLNG1p/3+69am+x6MAcmIpKXJhk0RLDrttskDP/kNN
5I2Ibwo1vsO8p377BrapjRIYKlyyXYkeA+iZjQCDpSyYDhMc1hPpZwo2QC8nHn+m
eSGH+6t8IL5PE94O4UzyZkE7gZOvI/XSMMd6AuyusrJ7v0TIik4l3xRbA3ccCI0s
7DMcl9ai5fVZCeKCrG07qjg0vVUrY/d1Nc/LmaySk9AKcF3tYX8FBosjGYFX46N/
KRG5hUDqC7dCMI80cBshJckuyF0Ou1XUO00yt3sV5Q0iv2vFaCe8yj7nLX2di9JO
mcjldtXxXUeg/MHtWuieaA5lzDw6tl36np3hQKH5M550d+swHB6GMcMKaDmTrT5/
iO83Vv7U7THIwyhrM0dxhGADMwrKU6jn8tAYH5Hn+Aje+Bk57AXKCFTok4MTB/+n
yRZyqowlNOKUWlEJClJXcDRLy3uWHG1pyxItwGLMxg5f1kzZqNsdbEXDXGN/WPOx
xMas432RjblP6vFt1RblBtQXaljBrQL7z3T7dFjcBNDwuaAK4gb/vY6ZVB0baXEr
DsDPUnY6X4TzB12QznqwuCnB/m8earOhTGAdT844bCX98ubwStpTX2fws/NaH3jF
pknVYEAJDRuLw/+LT5neEF86bU3s0SQFYRzglHKUMLPTc/MH0FdbDyTM1sdTtWup
Xzzf3rsYo2l7yn1CIFWnzY2BD9Depf/V4qmtUGBgYEjpUx9oMTPuyNZQSOIdMIsL
/CYXbigOOwIlx1YmrmfLn9LGTtkZ2uFWTEVUPTFXk2MymlekSzsvIsSbJCnAtI/E
OTj4mStnL1dUOJveUPM2av5nooQu0cFgGtcYgKt0mWRmwP2iikefQcCLY6Oi8UWw
+ZVhC/Rllo6WjaxlfdMhAefalG28B1dnZwhn6fTsuo9cv6ZmT54kIXoLa1oJj8mq
ONoZ3CFlwsUvVNFwUhjyGDXXViixAIFrcU57C1tuW0kx/WC0x3u5eZ4EG4XY9hfn
Jd67ya2htoXl0/NMnLD8N6KAQ7tAifDy3vKtq9/h6rCQs16wdmDPd18jZxZRiuPE
Y1uf4zqpHlyLKxC3PHpc61MEeipCxSRbQNXW2QP1vy6XWnfGYtXPGjv87IrWa/oO
O1lV8irj7pKYNQlWcSmS9Oe7C2NVWoCth9m+7H7ilhSBLseJ2TuyVQ6diuFgmsCY
Z87dKx01ciHxyLBEq+eH5nzV5ey9RhM/DWNqNZ4hmcvDzI+KuHxoObCzj90qxusG
RKcsYL7gdSRXOyZ7MnY2hSSXPBnsT5D0BrMKDMBhgEK9sddmCr27/Pi11FywW50W
w5P6VuTUsgUhuYH0yov4iO1HVV6M0SeIq/yS9gGuJ1pwPxwKkCXiRjDbqNNJ6es+
fhE/PXuIDSP3NPSdsNG3OQC6wS/PzsSzyh3rp7fZaDCEmObRUBFP5lLKeQCqMEQI
kQ5P2PsZpm/mTySDtFfteNAPabBiAqe0SDCxF9qn+7o8YxIgtlSvtzEd3sDwS/40
VQ8J8ublXHEebZh62hfdmqIzftQO5lt8Spv/cvEqqssFWSIh2xRSTymBaBMzrVQI
7BtQ65osSn+mghHVyQZpv+IIMTrlIWeunyNecSb/9VzPMipXazjUjUvFzQ7BEA2o
RAPvU8BGGL3/7rR16/ESS5jvZY6sMrLp/QSYPj1dRO/uA1KtWQNJhBmOejYn0cMl
Kx/p6CjSjtb2dwVBkJwZ2AhUWOeangDf5eL3VPzOV+YHKAedv63WiLIgKnZYBTWl
A3pkGK8t2qlLvm5qFKek0ckzT/AZjLjNvawS+lB9Tkefci6xN7/tkP+0osAbNTyI
u9cttJjLCIS1//YnI+OI1SDdORfGAAdpflW+5PmAa9G84QQydId4KoCwBKK8tUGY
4XS4VOkdEX0smVOR4pnfPdQY6NkF4G24NSx+u4BPuP0jeJnDX3EXgTj1+q5LWxq4
wYt2sG9ATrYxo2SuuPUoVIPIBFFwDcEB4NNN98A1RFN1IIUzU8xs2C+3rzenXC3H
UEz32UMIYghJNCk5ez+HGLolOlnz9JdiSdE2cKY/v2Lb+o/XrjRfJUmhJUsmrByB
IbMGAc/Lt2QRMs3zIod6qqNVsVbqH4I0SZSGxVzaLnHoftc/NuiT57m+yZnPE1a6
SaUfTR8E0zYnd0UepRSZKfaroy/5+uCqf6rtvqC1XMUdgPbVS9zP1rCn1ddoHZi0
RPDDCNkJsfWLwziqzSQOuHplleydQkjyToX9Zb0U/KEpeJ8MpsoBdaNyVPtKo6UR
D9XUpqpG5CVdeGJ6Im+dip4xw71GSQWqaIAGUZ5e+uPFtI7ILlsMwzSH5KfJBVMN
3Z/wS86Enoj1+l616TbtI6Wl7Vdm2XN2y2tn8eDfgZQqAu2qhJWxnFVT7RxyEbe2
Ea+2tFf9b4UykWwMOyj2/Ho/heG5mFWGiG/5vhdbwVltPvXMkfVFwZjgYWviBwqe
FPFtZta7UhfqaxIjtRflB2afvn4XhfRDY1xiEOy0LkhYk3A8UVqwvhMtYKU3Doo7
hs+oES3Q3MUkYU7EEwkDw9Z6/y604yiiKIeGsiya8B31jVozYJ8zNeM0PsLaNQ31
c/2sYxRkwNQZG011qVLb34bwpbSINP2jTTFrEgJEIQI0uJ6dRk8t/W8/g/S1ZoQI
ECVfVmjsDGD2WcrOUVydP9TsyPL2Zju+jbvm6+qdlrrXqbvP88ElmHftACYYVMz/
sO/XipA/kaBEUJt7dvX4pzDbnZcwQoo3691UwN0vqfC/gJ4rp0avDezIhltRyMWM
RxLKiMLzjVrBQ9I92k3tNDUT+9b6E+wqVQUEviX6I/E=
`protect END_PROTECTED
