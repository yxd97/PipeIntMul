`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M/7nFACL57+gfyP8SQ6MDWoRs36VphV5HC26bD3fx1MRGikLiQnOiQ4Y09QB1Lek
pBL0A6pS4oh/vEX3WZpzGrFzy59bXTPM8n8+Yz4G64IArJRHC7tXCSk9ZHUNRBRf
h4Osj0aKuQNy7E7Jcb7l3OgaD4D5yM0u9dWL2BGJ9+40WPntoTKFzqEf4y+QmuOy
THJL8CYLzHqadM6Bi1iMlnY99t61Nq5aiycGuUpU52pWti7bD3A0AHvCpPI+i5jN
YwoV20KGpo7VGOJTdISomqHL6pwWrMhxnJb+I796oDQCek+sMLZFOrloVLHxQf79
hoqJml1tMQcM5SLoMGIl2z8tXcHBvZSEbu/jC8SnW9M=
`protect END_PROTECTED
