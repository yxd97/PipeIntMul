`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KV0EFWzUj+i37A+MCyJQWlxcMD7di3I1Q4HdU2IK7i/0Ql6WGiQu9vs7NMGA7U3z
X9+WTxaGzOm4Z8P4El4C+E1KZKK6NN7P/ASTpuUc/6Zo5e9cyc8PYjfcXrt79h6w
cCb+h3F/CoqXd+WbejnQRQsRrCaHzIOempzA4/jUv3MhhS8/gTbMcv02W6JW6Y7Z
og7QWxx/WxCjSG6IVzVT5E6BpCw6CDijTdKgum+D5gXMagdUe6EWwCRxnIlGlLfs
DSKZBB2cFvB7KGOft4GwpQJmokmN8MrwcBkt+D2HtFijbM8H5EwnqkO8pinq2sju
W2ZGRLLgwqCS/m7JQkFR86CYpywmGZKPSj5jxfHOiQ+GaAhcdG5ow6QIvfh5CgqG
yiT4BnCJ+yRzX06uCIb7i4KybV7dU81YzoPuWwBmcBg5k+E5f2462fMAquEkmRXI
Dz4nYKiHtOyYNOXixJjmGW7jp6NmBI9HCGVamldMhqVZhG0KA04qYeBLOfCw1/TP
JRJIM1mkIj3PtiervsSQx1GMapykUCTWiMFd+wqnkUAaKTatQSv7xcTTcXT/nq6w
rf3cAk//mFC5kQJCIyzot6STg+GQVopA2gy4yv8QGjqfqKI/ko6SK/1i3Dr9i1e0
QT2jzd/eo0ZWg8nZ0etq4w==
`protect END_PROTECTED
