`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zigiqddwTT8cU098GmD4zuy7lL8PxEh+3jxpWpgaadIjFUsJcTzvXbJ+w83o6wq/
5EYsd+4XJBQItF4vnBCZNLhDRh+ruQs3hIR6fZpuwjLiK6188MikKnLbON4Yx+Nb
9QUvcTKaE7rfthX4Xjr0b1aQCVHxUa8snPy+Xu46HwlyXYVeMCAWP/fWuvI3CMiJ
kMoxcQl4apBBfAjdO2H8GTgWPqKzYdi0nnFT1o+PRuGTLkJPQ35/c/6LjYGTusnQ
dYEhpVn0el3OLY6yXsgQ5QaXPAye8YKhhC/SiPJj7GNNn9PwxVVuwA6WaLaoxBy2
GNCpt+HoLg3YubiMUE2NVhvG911nJgOEDQLaA4+E1Gk8MeJweOXI0xCjBVQcxVjN
3ihsiCRMBFbcuybSKusby78jTb+rLAYrGxGumc2dLhD6lDisZOUJKiVLonxdOwBe
DOuTKBLMvmv51gGVluWg03VuGn3qTOUbc215V4wftM7LaDx6onOMQp6J6mVzWH0B
5f4WXNRCxVpCxHCGk0QtOgZkxlZPfRPSt74nnXiUl7oIwOTYmLKwI+tapn4bar99
`protect END_PROTECTED
