`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FF6jE8ZKYrogwc3qBxNLhmB8zVT3kkMjgcvjU3M8P97/COr5F8UL+b3bQnvfCkvt
UBcDjKlTSJQ/hI4OpYdpWupFVO1OtSSk9dxtzEz+5j3aXV10yNOqv0wZTr5LvXWn
n0ydFmN8m56ChTRhEl4aWEOx/snRkOjeWmaxXbrvJusYO+hVHREJXGdCsROCLg7v
6lxnQqZ8ZlMmzbyLyqr845DKX/PXYLsd53Xvcoq+r22VdjFMlkVEi5enK737pVjE
qOsrAr6exSmm3CwRVTj5WmoEwZ0W518huobgzIgAWdGxWvKdXrqmPOcB70iB/4pP
PjWv7MZ7/+TSOZixmbtDpIbxxTF8AZj3iptj+TWyMjripS5Bb2fgBwQ8kgTlJdVN
MPPX28KXgH/41Fde4WuT9aQ66J9fa9F//uSMlCa5qFB41/FWxYwm+f/vU6YcNJE6
GKNOT0jLdtpAH+041Ub1NZPCBs1qUXUDJId0a/yXvinTpF0mWij+kG1RW/b/ynI7
3cVfM925lgird4Bq7mLz7YFNXWTBjv7T8QdMRbsRmg59rwR4NjD0f86wC72w9lS9
WQDJUMNZk9VTsyf7svwE6JSrP5xs93agz54SVw1wg7tt4tQJBASI1Y0XmKYH+l7m
MCRR+g3IX6ITQ2CikQBmSg==
`protect END_PROTECTED
