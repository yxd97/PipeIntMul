`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lV+zEpBwCgOh16+3fqFhv64K9edeyQbbQ835gLZjyrYV9ShC0KYc5bbPAcrCSRj1
cUW2Vw3+UFB4fxtBWQu2MT+OhHlnoso+YJQUKQMPS5CoQj2hUqK1LEA1Q9rtylQ+
N4NPfzabub4yHgBUwGa7JDHJF1+BXb2/TMV3jwH2Jqbl9gmpbvFoFFiFLRWzuB9N
mO5+GKMUt000Y7cgk4XWwmZwAKzbt23mmv+xuTkuLWkEicR2OXlUyWtvQi8ep2R1
hGfF74NEbtBPtne5Z1aARl2D2CMCMKLSHXLIcPvstw0WygowuDcT9XwAtT/tWTv2
l+wxSBWwQfyF7n99miqY7f8/YKdjbXbj/phrl+xrrTMhKvz74HIHEIV5bapWrD/6
N1A1OSK6cUCXBx1UF6tcJR4uOwKORoElwSvrZfRT348=
`protect END_PROTECTED
