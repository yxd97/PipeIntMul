`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8e8uK0uJmdjxpSGvbbOrKWX9e1i+7hBRXhZfjJ08Ew1w5olZnZZa+piZ1QTWlDcP
F10RRgKrHntbBq8/LuTnMNPb/OsEoytEXEyNmRHHEqCRUdG/gpdS9lWq1j57nquw
PPr17Ate7kZOE/OVpbNZliuWVIomAbEtcXWI6oBrN4qXVEBISHK1H3QVv2DkdPHX
pASjKARIFqaux5vJdC9v3iYWg0NqZkFic3Zov2yk33vs2BhiBDCqPWg9a8Tr/bm/
M19BLw8j9wca6ztr53s6ReVIaNHL5O7F3P3Z8XsY1m/Vv7bPHlsgfSHd/TpCgtNh
1RzEagqKfCoj9dNbDNqg05xug3zgGN4jgwf8A54/Nx3pIWZb4lTELXQJBEqin8+N
+F2D1Dub4us+ixjFTJ8/oomoSUzyqHw37hwczezzeiw5M/UL0NpFSUq58MeYbHu/
EqJE3i2E4Pio18bCF8ybKKAYpnP/4avsscmzq5WlDGXfgzFFLPpkY0JFu2fhKFqK
0FE2z++EHLHq9XwmQQqgB7A36IWu2GykFpPcGYMae0ymHButrd8SolUkCffln5ET
MNBUyaGxJKTCn1GsWO8tYOtBFm6QjKBccF4S3Mg5Kggl1utB8MTPm8HFWuqN0798
LzjJYXprmM0zkPGr71ApvE6sdvuqLghqYso4euwgdYQreIo82/xFrnR6YsYqguOy
VHVp94Y4lA+Qvrda2u0WBbOM7gUFIogPNB0G2ZSDuuNVDBWCvH/F0KhSV9Hjcm5j
kxPZ6oysO+Oae+SDhdxjmCONMoZrkp4+10Lzwl3ScIGFNSJv57Mu92H/2ouiuJVw
kgFOuKQefXFqwHtfWvYHrAU72DJYWNij4mDBXGEbhgU/ROl1WXnhKY/gzTHnRehQ
/g7VPeCPQQhyn6myEqEaS1KtDfE81vp7ByxdbNv/ay8TxfD5oYNrDAjvjrUHM4X6
`protect END_PROTECTED
