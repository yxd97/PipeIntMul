`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hdh90gmZT1V9t8z5+FHoOZ+jrvAt/TENu3qvxDHiR9JOcAQjPMAZjXV0i9Afgz81
UCMHB9GMqj5iFYhp8lLTe/zAXJLxeImPssjHTqgKidl3ZOkpLu2r86WNv+7mTsWD
4D/lEu7S91UgxvV4yYcb7II2l4U8U8OStdbI6JnTr4w0zZuEkPzARMOf2NXWM4kw
BegDSZQX+bGz2NrdocJJY/PQaUpRWqNlRu5+uatre5VkBXI19KHBI5L9dP9Zk+cH
0yLWkeuZkbTCPcR+n3t8rBmYcdk+3x961TgVXKQvf8MY4pUqEfLNm9+ADsZPa/qe
E7I4iv064fbjYFmTsEMqp3yLk6Z/cxSHd+a7ImJibWrwumiUuuXtWr20DLPpMskt
CmIKISdSKZIEZLB/lcLWOA6Wql4IgVj3aSsBARAAELvAHbmK1n/sKOai8Xv/iCXt
jtr0TuTbBoYpRnTHh368hKolSC/Qxf1yddeKf9GWa4hyNttSxYFO8wuKA+GHIe4W
sXTU32zDys8it8ma4g/RNgAtmBJ92WvseIAErcnOkYcR+McoNcfrhLmUTqQGcqIJ
ZZu0bAB20GK/ADeAGFOR8B7Fxpb1cfyBJKAGbJd9pMd6Nu0AWJe4HJ2SDBt6J4lN
9QaLLWqpuO70pGwKVVmMNDBllAUoBwETgA8eqDYm9MFLH2HAgw3bfY0a5LhlPELT
4WZRBVvpm+xmpHxSAa7c1nQWU8MNChFzuV+VB3kawlw=
`protect END_PROTECTED
