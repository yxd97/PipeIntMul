`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3XanAnvAoFT0dVu6SoMCIEh4XD/eKB7Cv43uf2LQWdcp357QoyUKSy7M7X1kHePZ
yootTGNJN5GGzi5lWA+aewPcw8PL3p/mScdX9Gd2C1QW/MtS+VP6IG4fyFQcrwyS
/5uW1COzGXrkkIw+ReSeDpUNU5wl6IFtorckeacVf1vFYQjbabMEXS7V/Q7ds6ag
/UklUzk2/kTCq7Wdz4zH6sXeFIuSsxs74imHKIF93KvaSlgdpDsSFvQj2uMuKcp1
CkO+LI6EyRL+NWqhojpm4NW2K8H+mB23XTWTxyrhs2kXE0qsOMwoekCzPAVCwyfH
DpYGimLlrkQ7oFccbPbv9MNXBOAvAvmv7HUZ1exw4wMwSNWvpXx0RQrkniUoBCn5
LjJCDl385SaebDqyxdO7BxqUVBjao96VKji5t6voSPnP78B3xUTunaYe+B3BitEF
SkJH2uo13G98ycWLznMhm2tU4HrF7TtzAMilF7mySjrMht4U3BtblekFj81MvKng
bepUgaLRJL+hzELl6WWGJeiDVgsCOsKiJql4lxpmh2QwUxD62cIBHGv2G1tMf9MU
yMMMd1PHybkp4BYhMy75TWfvwoUWyQtzF3kpHgFGjc4=
`protect END_PROTECTED
