`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPunchkLbpD+7jLB3ihtypCgSu+RR45RYL8o0q2vWC1Cpy/12E5EKKug7pFJ38cr
eXTIr2uC6T+GjHVZQ8zdEWbAebXxT2BK4hFQ4Xih+BsgLsz12xT34T7EqOs+4y6m
r7B3ek1/zCRQ5gDTG55u2o2TveHEbZVRASUpum6jaxIZjBMqYSZQNekF7FN/OHAn
lU0o3RM37kGNEYAywrDHMkA1ko02iZ8IiaagPDX8KgPoJ4Gtpuvmb8J2GtouauQO
h+RENANHYYQs6OagXSNiIjqYvVrwXO1GqsDIbtoXptv/b9psTICPKjtWivRInEe2
hDwQQmyOUv1KZe7XQBpGT4nRSLjf6p1JNYXlcWSd6XiolcRhMtoAVz+f8YF7YSVr
i38YzF7jIevNJG/sGAwKqz6yDLHimmEZI8BbfPTDVGcpYGEb46STD94w0I8Vyxq/
0KEP5GbJPx3m6QRFUBv/7tG6A8TCwKkHnvdGXf4t/OcJXbfUaq8rAZzh9mFRhv6R
PkP28/z2Klqf0FQ+oYei97u+BNqSC78Y88jTBFbSrGt0LbKgnhwNAXZLuSvuN08S
nsMDRWniYgnEl0Q5qvOB/3pMccTos+uyOxtdO3waDY+Axlr0/PDwOYNyd2Hh59BA
kHDhSVTWEC82Xtk0lgEFHWdBFv6Am5hWIRI/6y65FAIm0dcbGyQ1F8OB4FOtHLOU
KjgI9pHKdP93cd9b8MaZkiKWEG6svuorQ590KA/aob009zSd4iEi9DWvBCYP83ai
tFa5OnvVOobdta53EsdNTVM/sjWZ2huAbEixFTwxWc8XzRRbj+WFWuhJqiKbdhZ4
J7N8XGkIwoVmvZGcs5T7kI6lVGt1cIC4sJWEd0wZXvUxA/0e/+mhDHVZ7eGvnw9t
YmU6Hz8BtrqBydubNiQNC+zdckptTSoYClTSXloa3S+a40TWL/BqZ1nUXhDXj569
V6i7P+sIiAfyJ6EWxJiqG6jghQm4bSmGQ2PTG/SiHdehkXNehaZpiNBrPyToqfr9
+dku/uu6Pfxr+7kloXaRIkjymwAv+JOZUFEMAUPoMD23IvbaL8LzAKibEi0AeOab
U1RUB4L7TQUiJkRzskZXY75sT+iFjtOT+WSZVKoeg1CJXQoEo153SSwhoqPjCZkg
msSYdDBchRlxkWo+BLubpIRHXRdCsud478ONnCLoe4CFdwJFbvOgXfw49yU+sbgQ
8gAbh9+T9dFp0mkji6HBYtmE8nsaon0S5mueuWsCPyDsaUW7TSVHNUbyQG28PkTe
LoeEVaDTNpwehBdlvkp81i27TtO/ayJwawWylf51sbq+0tUtIwix17Hr/QiMhxOh
tEN9Wx2cGQKp3YYLQseznxpnkp4qlBM7qox7czPRV8n9b9HAn1MwFqXAMhQbFjjb
0xIWhNSujgS9dfhkQJm9KFSH9u7pjacWob4g/4lxHfyeV0HT4h2dpEW19dCXN74Y
LXVVjIxHcxInCQh84/IG55iHt0HiYysSeEP7Ht8HmCzckfRQ4oOXbz4dZupvqrDI
zweVTGmkAx4gHH8ewEU74cK7l3vICe4BKBu40cVOU54911tvwnz462/PAt8Mxbmq
uHAeeHNaKc6yZKC2VZgooU/UlStsQwLKy/HbQTSQfKdnDsQeOZ37mc6BwsgR3d7p
BBh+O/2i0IPYLo9g7O5fhFx7DkxRxcbLbhOcVarYMbifVZ/TQodNrosyo21YETzn
2AnwGrbLba+hPcli/PLXl+TKTEA+Fz3trLPu1iGQu4tIlUk16dtMT//33CLcecbP
JKBfsjzUkdjiVwxl2XfuBeuXjCtKkCpod7nhRACc8VpNu7oNWhSHrAAN+uyFOSmU
tNkpIZe4mgGz7d74YjLf1yynwjHoak3RX50qDIfd3fSy7wyezNsJShAcWvkXR6Mb
fvIOF1kJjAQYlAwtIw+Cub5kV3qPCLtmG8yhzBrl48IyxaYaLq4pQBvM8Vg8s3Vn
FlLQoWOOYS1UfUEyeOtHreWd2JnVsdV1QMuHB18AJHZfFIVM8hZZ/N0NRL87IPe4
2wk3xhUOxIE5omskKASLdzLhybMmmu6k84yzJ2Usd2ErYjopRvFAlY88Fjz4rWtW
ah40dde+WeE76JxKIzZwAhyny09H5+9kB8wvW8Pb2QVUJeO46da2mAfEzHTS4zTf
r2c/esISlr4FV5+AbkVcljuISY1/klGuWXd1FqYxVh9S4Ii2ETlnfG94npPps/dp
7pQ6GhYJdBEwdrhWtyjdlPjHXqTMAt4W6JKGKqeaAts1b+QONPmNchhYhHwPA9FG
7hWq3B0O0CEuETmTdUuA3g==
`protect END_PROTECTED
