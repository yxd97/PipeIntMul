`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
j9PjDsk7FRS9wxaOQgETHPffGB+oz8W/Mq3LdkpT9SNolkGyB/J7ZTh0O1B5LUnl
XyfOlSWmJrrlN1Sr/iJ4khu42MGeE0fm3s1FfwX/rVZQ4gWZr3TuUVZ/e5pmWWh8
XWjBKrDrnCHy+XhCKMVGXsnhC+lxsLWAEtUOd8lIPh3CMCbvSo+XghRTmC4F/cQc
HWheGiFr56zI470bnYgUFyrebgysh8LRXNnAaDOsgvZdNsWYwt2JkF6J5Zm1R2Ff
MgnvXza1ZHtedlVA/sboBYVVcnQlRtEETzSt2PtOCsll0VXw+ekfo5K9vkUfs0Cn
B4T8c9mUwpBwe6VMjyOOeE0vrekZEv+1bW04FaOAPxLVj88VZV5KSW18K/DMw5le
ZOWjs91/HvqckoO0NY/9Qg==
`protect END_PROTECTED
