`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rKcNNB94lXPCtAqy5eEVFlOovmABQs0Sc4AGCJytK792U5i9wS3iiGoHO6ZIIpOj
xVz73V6ccws+hMklsPnGbuXzCGNsIjnYKAvx8UUtsKKKr4PecPMWzvcB1TLysyuu
MriJ8p8frIbgwKF4fFe6EhJuqEXyfcoWVCVa8xMA2QLI8R9zzOP5pX/hnzjrWDmr
2owaRHZfKFlH/sLoFZLAjjr4kHCRkvtUAy26seCOhTUmlioKMtSRhFtotashupIh
iigID6NRzQsMbqlWnJTHihihuO8luJtRDAO9MguD41PMGCI2Gfx4ns0wMRllrfHQ
qMuVPWgVhQRb2roKK6vkNm5RENItqv5YFjL16/oIM/ROJ3y7zy4McEm5ylxZLew3
vR4d2M38TdwnN/WhwF6P4KtQB0IS8ghsGsy+mNpbXuGPo9bDH0SKCNYsgvnuDodp
u0UDtxEnjCI8Ual0nz8fKe9fXhY2LpAYPT22Sa6wNW7NKUklwWsX+SVkSML7NHw2
q30Wngiy3pBcQlamYJX4xXh3YxKDFg2H5MxFUB1MnTPIgzCbE2YyJKUMqsT25RGN
z/NdU/Zvz6lrlRIMROhEBzBt3mR1vweulx8TgMaYICy7OQOu6xLyrtg1fWS+fy6P
hYuyR4NomyomMIAbnfVc4PkS2bfW5xBAgGL7FvLec5Ht+/voc2iKgx7omZzJ68qJ
Qp+sno6rfhoInFMg4+eyy3IP6mnAxitzJpQ/dveYxDYH9jWkRRTU+Ck6Tmq1ISGZ
vj9e2NvdASJCzPq/YPydrvDytSX4i9LkDKg/FD9WSt6Fehdw3mY6hTconh+L4xQs
xiFOg0bBBy/kMSOJt3alKPSFXZiRxEvnBrShH+DuxVensUyVh1N5eMf3hkriCtPd
j+fgwgB73G+2Ii8/YG471NhdPL49Q7fuvumY4SIhjlTU1vEDsGGuyOzuBXHWYTEC
LgcYHYmg13uvWTzuxZJlapA8TjWMDnVcvv/usT0+Aj/RniwcLigaBSRZSBZaMItm
tBOcMTKJP1ELovfl8l6CykfIB5hy8DLeF+AD+EjZ4pt9HjDEB2esccAm+Nm+YTuE
gN9ISMkKrLxuTxKTdNzLCeP3g1O35ozG9YY8ossJg/wJS01LoyPuOOl0eHBfS3Ka
M3kzgyXgwb2jPR3Z+jDngg+kFY7LUku3u7zSScA8ZwNFE8kgxBiCApFKpv/wl9A8
gduzuG7dR1zX7YuGHd70GwoburwjM5VMRvxPtwTXoAMnBE8xceJkgys3FBCsWZzt
XiKJG0jvrYVazagCqFP8mGM0/Rnbe2P4naLkIUQQiyHO93F559D1ebHtlEQTAmLw
raYGLDkMx6HQtXL6R8EtlpcJg+/kwo3zeOYpaNTEUzrAO9Vkn5O98+whkelRrKMT
0LTxmFNAlE04DorAdoQ3Nmbt71kdhZ1qbvksHVu1cCwnVtOIHIWem7pHwGfvYcwy
Kii9kaARKziSP4l5YSeHBpjm9SnsqVIvuWeDKETFOKVeh4TIPElzCSEQ3x3m9Kxc
wgw1XPgM/JelyHQzokv5WCTVtpePj6/pTK/JuMpsHRgOVkcKrY/iFbct02RtRnOa
UZTmZJofzgg3JUj28Okp7CeFiEpUpzRVnEG1kknTyjy80Mv/J8ApZFNYKROH4pLm
Hu3zh9LLlJb8rliUOQw6CSoTXMnEpPkfnqA+EowwG8x706eEC+v7wTR9J+XdUrlu
eOlYH4Fn9cDyFaYgEs/YBQfOKIj7w+X85XbgZAs0L6dfXPKA5r2M4fLYM8u0F4Id
v2tAVLoUK0mIHKQt1tTebG5R1TxD9FjPirqZjV9GJ99SvB5Ht+vXjY3683AhSm0b
I1224AxNSpMKPflc0M1DWSEmdekbo711uV9wVgDXIf2jy2EE4apSHj0WK+qAJAxr
bozkPVKKtKV1E0c1PrIn3poIR2SIoUWjUmWbaHSpC4idLGj7uCPxj+YfFr2sSe0/
yBhTvQ8+hs4IQ+hXx0dPbr0FSnj47NfWCUwL4Yb9Q5dvRXD1HuGts+jQKwyPxjBl
HjppNICNvf9WfdIuM6IlZRBy4r79asqGRShGjdg6EqUc6Nh/Ba7ZiVSgONB52HwC
kGgDAQbkOk+EOXkyiF3g7OEMmEoJTwgjWeJ2+q01lbrrurqjApqlXa5bKLS0rSsn
1HjkYw/oAwNj3XnA/1DCgS1haSBcHWmacbR+knGZTrsA2s3pU0DWzLpbRhN2HLYh
b3SN1+b55cDmE81/6KI2Js+jxSmUBgI3p+X+6CTP3t8hrok9XQSeCXUP/0DMPHsp
pZALuYofSdSPRNtfyzwKQsg9IGbe/GIJdOd6BDgdN8umtK6lJXk3/Zu92SURduS3
J9UuMi4hRFazrjKmn/fkEcWUDpTDIhxT2pMHN5dT6+KBU1ne4WxEaEVhG3jo5YCK
rcBAaleMhVrGPrIdo/QIBhWrO2Vb+yBOIepmj1eCuxq7o8LiOq0J2NFbN1achDnv
NH2t2+eBRLKqQS1bDANCV+4ukKAeu0G+ZVSge8knozblI/DyCjcx7Ldy4Av77ZjQ
6IMVkO5PemvrgcTyjCHYky0k48y42EW2PBQL2QZ+iSi9bzDW9Rnqtqx9nfTE7RLB
/7aoXIImRo2CbkXzngiVyv6dtu+irPecBgSwsKFTWMIEixRHB+E9gRpYAz5gBF+w
ZUEPypdiaBmwpXQi5s5qyEEPw2UXRn9rKaW+VarE1+2buqP9Kx/i3f1Eti4SN7HH
6wtbiSUVuqbF35BLTZA3Xlu863ZLNLD1I7rjrVQGl3zkNw24v7s9Dk8NDP41msZP
DK/wjK0zkaH8wa17PiO4mseUl3QeGOCedRwvFd3rp+wd/wRsU1edQyOlM+0NdOQ4
SAxQSOsBg6uOAi6Pfa7GTg==
`protect END_PROTECTED
