`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HGIiRqZedS4opLOpEQFz8cXY0KD+N9B5Vy/joZH2MwVcFEXwHkGjw5eYIeynrqlr
jL+yvF68H8Rz7n4uBNdwe9F5IpNYGuhfA6+LgILIMTo3mysdZXcDCrsO98YTAvYu
X4NxkyJZg6Nt+ZmSBhQuRtHSNleiOFnT/O4BuhaAEm5FCIVkL/r3CUlNZjxuI96x
BZYjkQByfcX10BbS55qRD8lJi0e7HGZ8d5+U3+O81g6chsTcuyOT6WXZ64mU9kdW
jGjwmfkf47LMnvZxpJmRR70YDZKqFfPoqH3izqDbfYFETfXGC2JnUGj0ImkZrv/9
x4fDX5wjxfqRvHnvSVIzC4oUW5z3ppNoQpXYrvhjtu2BRPhblMnMlgZQtTe6WXGw
GBm/LblHR/xWxRlaAhn/WVKFlhnXpklHDsMPj5H7dbKOEzi9/RHdlX/s3bdgZOvm
z1MqUJholhe23z77iJmkz/oSwYJU2Pjfhb/d8A4Q6eEJ7WJj4Gk2PqVO6oUk0vl2
ag1WaS+aOdLQl5fYwyY6U4FhawgpA/egVzk5B7OakXxFBbInQyUXen2KCLZPko2L
DUJVwkyHlpwFRmzVzR5Ne/XlkxSw5ffQUnGzeqx7sknR4lX5WZkr9jObzYU2OCHl
S4/y+7z1tWI1R/jJggl3bh/n0RKvINB5FUkfQcwktB7pCR6ynbzPbpNPe7V3oKM5
KFVVEXD4AUYFQdzb0cE0KEg8axb4s5M6ndQMS7O7+MEZx2vM8+B21Hah1qLcom40
Yn0uF+i3l8wjGoIDALEyB/QGAKb9cYb/7K++fNeeIUFZ39MqxxqwswqS2iol+xMi
z6fRdkwJZTVXLiGPIKzPI9aNZT5ApB9DDHMXu/jzfjVsOFavKyrZpVbKCTYPu7U9
Uk1+eV3YyDJYOOnxfd/HmabkIhkQwidf5M4lH697OyQ7D1Oi59+MOIA0jd4wzWF0
QT0niRMAqDmfvjjubN5k8KvLuU7oJKBmadmOiv7J4JXigL3DAl9WQEZAnz3/LZdN
`protect END_PROTECTED
