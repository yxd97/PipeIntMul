`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pURQzIgHDDkNZpqbS+ZdQZAcFG8MaNNkkrUmZQ+Ngc804yGu/ATkZTy/A3b1NGkG
KSCb8llQlmzBpplrc7FwgSQM6EsW6Yh0dCrCqn+U8OJKtULYdm2t4kEG0K+3wYxb
p3MTSBPON8bsgQTDbKSeaOCtKMfWDlZh4WdsdDNx8F6nRHPtUBDT2EGKjinpyAH9
XmhLq+Np50V8AMNkhJ2GaD5jJyJTvHeQ+FVnBs9hF2TvBdA3WZyW15P07ZPXjo6b
owxumKMO6Rk1E8izI1i2P2zAsH5j9gKbvnS3R6bHSvrxL5anBSivGdjRkjzA/945
XhorK1NBgUC22Sl3QDfw8GnBP+HvqhQUoK2+aGNPlWRTmlDHS6k03MACwqVVAyg4
aEC8Uj3aUSnmZVu5yShbDWOYXUFbxqpEUYFfIXh+2NgDMvcYkBVNFo5NiBKnnhcu
hWW7GekxIzNUTXvq7o7e/ySdbBbmODvA+IgJJ5m7PY1DDI1UAzaAhj1cZ+6Y1wrT
Kzb1U8gxa8c26DQ1UrkkdgkOj4kPDan9YzQuLI9qhVdGtbCCngW9inLyosExTjb5
+JWUFdUcjSOfH/ZdyyHxNkMkJTt+YCjsVOi7d0z2Kg4KHYS4ClcI5AR1GSxurKBR
kKQD94wFMdE44mkxvwyjGg==
`protect END_PROTECTED
