`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Qyi3mJlt6P4Qb5vNnL3pfyH3q6OjndM8lhOS/1uhYVhqCpoT/bSTiEjCClY/tMxO
Zs+0tQB2gfTbEv5ixCqKIF5YgJVqHntSaITXJaqNIP8wSnLn2R1xh+UNhx55DWZ1
K6Ik4OsUVyXRrjMZZA1FeWZWTaVAKGuA38BMPA//B5rUXJcAuPiWZVn2KseZtUW8
zwnw9mIHT63erHkNafs1hJCFpYHZIjzGXdry4AOYrotHEqHvYDviZe/EkHUlQBgR
iPZdIS8pWMugjU/WzwZY1p0xI+DtVwrzTziKNCWTNrXn0R3ezPtLhyAIEGLCsM/w
7MpLETXp7JOr1xy++tQ9xcx5628Wze6q1rBhCb21z76wxxDng6iOJWqkxvcowv7V
`protect END_PROTECTED
