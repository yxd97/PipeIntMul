`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
056Dvzxg+LPzv0HEbUFknNbf9mUHzL9P8qOsKTtWpYi7uHLxPndpmr7pl+3ngszx
SzibaT+WgrKQHIb7bt3X7erZcAXqAkU90xp5Npbpi4JyEXitDZZsAlMuP3PPWmKf
ZQwRx+cmgcpBWu+0UCo6ZQyWnRx2BKKK05TTYtVzdpQYSIVUcfwa9GMMFfoGWrcM
/j8TX+QxjGCnHxgRte6bjvA+o84enTUDE83DF+P0Mb8e4WKxwIhMU4fCJPJlXdXu
PFRXuhVkz8ZIkx7D6Q48xlKq3S92CBPbn9dkAD42/myvFgPSWFCtsJMgyjU3A7pA
vhe1tKOd0UQ5Mdbfqfdlv94KXdLtNbzng4FQtnFNxhvA16UiUZF7yaRfA2of5sGb
qK2gOkma16430BQt5Ywt3QepObDzCgSeeGLq67/xIJZkJwMpd3nrJL9YmsACAAGc
mu9SDcl6Px2EmpPEJaWqMo8ig5CI3h4k7l3Fs06HiGQCnHDA3/FHgZCiWTcrlko/
VsJNHqwLZSvOlfJcWhc7CBdBFu7WokM5A4exURroAuAXXHnY0CJJrzeAankMh3yO
nKQgsgaBLhOBvoX8E2yjUMv/B5As+HHg7e7CKP8aeueemlz1Vu89v/FnwDtUl5tz
Y6z89FfwgzWD26Va0H5SCKkxImZY0oj85rXTJpwmIjUZNJFCWsE6oDyRgms1a6US
GyLoyI/4s6T1aRvc3+6WBUUxuyedrzjSlKJtb3tjoYtw/fgfJ8VEGM2CLNiwkaaA
b6VIwrqrqFckceuFzNzzBg==
`protect END_PROTECTED
