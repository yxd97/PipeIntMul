`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SJUvapTx3KknL3wQ/5rI5OvuLZHQ/d+Z3SeQ13k9+e7l58gRE5utzo0sCOJS+RXY
sw8g67g6BSPghafpm2Ru0N+fvS0+oi/QVMqnHsaUENDQ35yablu/L1MNJTldIVpw
TH27h7DgfQMZdYxARGUpJa4HWAHm7gLFgftQBsboLsWlVmn1sjzCVGQq4hIEmkf0
NtxUEf1O/GgEsnzFx3/4Bg==
`protect END_PROTECTED
