`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WT2pkNomhRgRzXyVUeFKbzJPwV0zH9z1HnUf1L/38yfwODmVcHxDWQSLx6HJIGZG
jHCKA+oqVYuVdkFJTsW4I3SykEnBpQT7lqSDsSMsindXfydWpeZZH6lBRI+uM6jj
QGovHR1KeH/4PYFs/DorbA/jtVV2qRXJwux5olbrtLn1eg+c0l/QgXgaH8e6hyT9
wO9lJLuTUW3/BPYBBcTeUplSxB5yyVokiHJU03I7RqF+gqw1icRVXLvNOw4KPD80
+BnNuc4C6a5MIRzGlsjxTUmbCtPmO4c9/ioKhNu2Pmv8jPwA09qlpGPVmG7jSpDX
illEcwRFQj0CDajfr6Ee1fKB5/gc7qiHo+kFhkivsPI=
`protect END_PROTECTED
