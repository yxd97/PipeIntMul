`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8MRLZjZWF+Tj5ocemds7h/cRvRqEPTT+A6/MRWzF/3frR4b01cFWDs5MfD5benS4
ex30YX7i6b+2XKfNwMwScfXaWNMeNYRuQlSza8bUpls55duohVtsiblC2AZ3fNBi
0XvEaBR91wxDh8jzmm4wkbODNhdRmOCK63R5Yce0YJ9edaidqGPlbFN70v/5EPTu
RUx2DqrWTBeau4DPw3RRYE9FPB4/NAex7LCX/8B5VXpBvLyHpr6V9ZTw6EJH3WVq
xiZNF8SioHp8L+6pl3YQ+x23JTVEePhXlABZWVUxe/D0Jkr/+lDcFPxDLijkTVw2
aVZFb5Drq733cHBQw1x8u/zp+iHCS+UzSQOi/wUGWLdBD7JJFDXxTwsDU1CPMf4j
Uwb5JFSB0lxDC207p5tECmpX/WPlqCIKpMVgeJziiDQV50cyZUHehaY0N9v+TI0K
BMQrgRf+H8k2fYq+B+mr1f03a1v139Xr1B8PcG/79MuE7CUcP7SaMkWfV13Fa/th
5uSf0H3mMzb/TQrS7x/B6ek8YHlhLm0l4y6uF8+9iSJE806iLjDiFe2zE1jjlsjc
/4ElDTDzxpFYYc6OB569oPIRQ1XpifddNbNacIsDVP4dBujg7k2ofTbPQcP1MUPD
VsNniMkZMX2bjYmBylQi99lVVMqBu6udvHj/V8xMYrMwplrBX7DVJmw5ILwY9MER
72WjD71atCDiXgUS8J2z8kmIa/ieYeiKl7+h/Ky5uyNL/YJzhpZdG9I89g9pUF7e
7mjJfeFxO92LcQmRgWjl2q18P2VbRqRLKECdDdhX2kV3MAJaIoAcBD3u26YQRyrm
Njfnkh08SHEpU0QqW0mtx8Rm+R/jaUKAiYpACloP1/MZ4K1J02zQUUeueaqasRAj
FNnCY7qMcb7KlNT2P/mfTPce9gUoTAEGl36wm2QrYGOQQ7veCBucAKwoHRnxRUyG
bCTh62aDtsFb9XpdSNc9WeX6Zo6aViLhOW5wnMsbXUunwS/LCwDwtQ6ieg+vc/ql
IdGVy9p+Duftp6HHFZz78Q==
`protect END_PROTECTED
