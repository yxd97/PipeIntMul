`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BRpVPONuYW2BEdSsxqbbSy87+xAACpKnO5WbZtv7ebg7boqqZoygG0Xylzoo+SLc
6Esi9o3vOarY2yFVbn6j+GKOq+8Hl7YygmfLEkl5GKVNV05IEwTVAz8sUnZCl1an
5Xql744acOCi0YlCRm8sLPxon3/Mr/k3D9XojCvcTWg/KrfcVQhRYlxoh0jQNt/y
LyAavhcZ1qaKHgYzDWSmWiDZpti6MCWcPneoVRvAcswa8PjcO8yl7Br/Sfp3znoD
zI5JsIN/LvR8OYAmXzpEeYOoT/kFCx+hoRYonq8zbHewkNXoiZG846/805puRCd2
52jXA34FxpEC5bW/TLtdo3ahjLHlp9PiMBYBWGrIIfeV8gsaaj06ggG9MtjJXiRl
6h8sfVETv/50zh5ajwFfgGEcNZlOynxL/trdsE6Pi85ebpxfNqWQoLxLLyEejDET
`protect END_PROTECTED
