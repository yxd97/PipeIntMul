`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Jj2PwN3SOpprpkiS1I38zqPRHrTxKP/SX3IJS56R9VzSdG3u13W8kJ0SYx0U6ZCy
RaFEccFGjWR+ZNEnqnmKSbbDoOgZi/oihWmg9ELRHOlXXo/dTI2Jk2IM+nPwiJ4i
JUoRbJrag9WU6NGvAB3Jj2n5avQRU3UexuLd854oCytgq6nvT4JqsyApFhXwAac6
sJVbo4bP8bTPg2jV1MkceQ6b89483mDJOXjmv3Wz+amdTUxugyI2thk5c6/8mrRg
4MQLuxhODGgwYJwLAEHAUyYhiLBFvZv5rgDo3SK3SDsRHCZljIb8Dwn8mr8FT4lm
rf0pSKXnbDW1Y4nrPlpqx79Q40FZKY4aPu2zzpGKe+dv/siNyicr7/rgfvAzCBJJ
u/WSoSPJA4uQgChFq2ptkVqdq1R8/kyqqOtiOf4FvISHLkbESagpXVG/n2WeGmJt
jnvTT77tgauKI7kPNagFV7bqDFie60nURk5WOssB5JE+pqjLHEeo9BlPc4CHoeKy
2NmmmonvRHxFbfqOSp/mfWbvdbjRdfsuqfdUFOxQshHl6ojxMHgh5MHaBTZOtHfx
9T5bxxGtpH3A1m7HXdyTXx4LC8oWgLBf9QoTK6m/OcDykXLZW4LmdDqkqJgICxBz
SVaVVrLrcm3QEhiVdE0sahg+mGOmpx1OjLmmk6oJdNnZCtyWhY1FUutLNYEJ1wIY
Pm6dbxTWwT5VY12VZPJD/n1CY1PzvMGvPDuwZMDZxf8p1lGKzZ/j9dR/ONDAugql
6iloNhQMysK0jyPRcFS01A==
`protect END_PROTECTED
