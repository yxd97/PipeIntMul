`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bHsxtl4DAkkilnrHCYrZVRAj+VnHB6C1fwsRkgkv+xy+5ceVZyTCQB2qh4bmRRbU
gbIqHfl1YrAfF01xon5TPgbPYPPxK8UjWygPySpBl3Tm1ChJugi5cmd5Ri6HAU3A
nf9mXaQnDOy1x1Q0zLIJ+hE1/4DhflMQqnuklja9TaG6V/nlQBStRUASksf3LB8t
HaqypheF1aFwX3NltLHX1B3LrgbUHBmDmWQ9mvmW0zJjne6DGpwIGd9LGqHVjRiY
c/CwugO0C66iZfvIYTjK1qt2stcW63DNibvr+O3z7lS2PkldHxDnx+PnQTQKt8A9
t3O0N9p8BZdgu2gELqiA4xzBXhotUr8rURIIqcFbK9zHy8XyMoB3/Qr+TZH+fiid
22nM/7rJw3PqDM0x9VwjatB+QsB3spd/j/XyOmambss=
`protect END_PROTECTED
