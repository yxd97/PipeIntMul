`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/B0wFuxdvixkOvigWMHvDbiuGzzoqsHP2pQn1I+gLzW0vcqCuP1zWHJCEPD5CSrH
rNR7LfaN179rXdxy2lPdXTbZFEmbV/VaJ6746Uam+DxDEVjOawAcqHFZv4upzc0A
tzNwMpoajR1ShV/HjB32sY+DiGafnLTL0VtUCj7HyTfrg/MJydXEHGi7z+mHAjoF
iGalLKgqEDro45Bl/vA4q7v3CvuMO7k/70tH/ZYR/iE0+TZgWcp1WPkrE1yJtznZ
DTjlrCBMhPdH356zQ933+bIKQbSSrRmFL3ldPMbIOLC9w17fS6WyH2wKn23drvi+
CnTTAnCUhhiFME3+Xu5rMHDZNYXMBF1w+IlmMV73vh6c8oXT/qoDsyuImK+D5u2/
RNNokAHpBKCbJnR0ZGQ3paGYwRO39/TbA/QWKGCNItiK0V9kwHEjhDeCDFNud28n
dwgVyH9tot7M+BhAWq2LleqFuQYifwFo1qLFnVQ3pDwoRcp+BwR7XKLS2r5MEnDb
KS0OzJdt0QDuhys4YTlGIi3Br/qgA3w4pIqzZq9LmzLa9uV7jV/qDOvtQyuN8LCn
9DmbFqEBL0iPDY/cB+/Xeg3j9z9CVDkGyz2gutF+p0rH1sozXS3bthMYNZGfejYn
mZ2OQ39maF8LJaZWdoeZryNR0wMlMy6nOQ/bNUu/cbCSXt28gEClxe4zEl6g2+93
Eko4WP8w6fcY5OCSbbA3p45ZfuocfLLdUAN7J/oPJGszOC+EHyJ9ZtRABgzXqolW
D51EHEoPhK3JM0mY4RA/T9yazDPba4uHE2MTfIsqNKOgFQHxNg7rqnIfN0WDOwvd
OiyUoxyJ774dDIuv5Fq/o54quwzWJWitWdab5CMQc8XEdlUgncXWUGgCesWq5ltk
zQac0SDCDwFhWlQm4dXH0jcgncf6rr1k6Q0RnXD1k6v86mQzvj1IoR74dPa1/ZSZ
Jx3UlapzePiHJeEwS/VyVShXp/J0OSyDOrrt03AWxwQBwdelN5wVkr0lP6jhlCMe
ll0aTBz+9BX2F7BsBUg1F0Xe0XFIjsNB+kXNNKdhpqkB1ZBasOhKeNmRwyouK/YY
eGnEe3ecp4Eu2+fOYg29cwfbrJVvqMFdvffyF7/BfBVzMpZYibRWXmXwkrKG2TqO
35hAAC+oCIJtB1pP4J+ac1A28tXzzzqw9cHDCGFKqLUHHTHONPdLwIB/3T7a66+g
vB5cPYy12oCCaKvvMUCun9DkhWb7oBVGqkI6vSst6+38RX7bKFU7VdtceFr6IZJU
OjlsFz2eyAk8qw/7JEi+Zp4C5e0+WgJifN7KvsWUIQcoXJF3JlIlImbpI+HHoHr1
ecFrnyAabNmtcuNp44E9wvEkqZyW9Na7Wpe4oFxjcXtNs5mfbNHylXOQMnXPgiKE
cp+yXCC6XiMHYmKU4dvTF1lOKZhM9fyn9jUT7IC8W2U=
`protect END_PROTECTED
