`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JvG6LItVHg3LE2R7vOJmAcuU7vKsi98Bu4vzJZ+lzA4puEYs4u+yv/tolwwgPhNR
fWgSXbnzxNbr4ebAoc7dQ9ouZEO17gtLxLw2EW5VM37Qic77zcKuI/p1dAqI55Mt
LsRDqUmosOeL+c9Ey7f3PlCo+Ay2+yvNlMGLdjC0Fz35sdpQXlbVnF4uEqDW04nq
/4+zAF0Juc/iDXVsFvm04Rc6+H+6nWx1dkkQBqG+pzMF+ciYMtHK3ZTMzrmzQPcZ
PeyBQol3oO46z8UteulL0KHoovgz0dgYn2mxD5Fr7Eb5NH7J1M/yaqR5p+TLyki3
V1l0XrSv5jfUZ2tzHNBYeekg7UJdKzzPLLqzMAnA3YwpkEXngm2rL5/0pYJM/om3
N1dtVtsXIGO/DQrfdOL9wcPvYwSyZ6og8vapTiDbxOjmsACM8wnkjRcL6Ngujrfj
MUzdVoruAak2aD/THQkkJKfoGOmD+EhhrC1tAQmYFsGlU0fKhFRdXkbdiPYzyS2n
6Hd3icDiptBmDBti4aFJYXNgcly2lsDZEif1+6+3LIrwvyLcueVPD3Kh6oiYQsEr
YcMTOreGlk3OP7+DWQqG1yU7VT8dGV7RFxu1oWkl1v3CGx7Sy5PAVqkhL+IhEJEz
t8Ug/EN/3kbXtG+Tj5YYxcxZxdPkfDaLWy2tQx8vuU8R+iOiMaGf/uk6yDxRzKP7
snCWtlyKQOUAqhpZq31fxNGRoekNgyhV4hK1aHGKrmkvjpWJ9OdLKd7H5BIALnrI
`protect END_PROTECTED
