`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
i9Q97cKdinn15WfDY9n7XNgrczJvpzkxzmmFVLzts/pfPdNX7DYYXB7saE33Fxeo
ZUwZp52tuFYVACVwKDmJlw3y1nl9LXQY06gyBYtwrFRYrsOlangfSDSgIaZZ4u2p
Z50QgiNcCZt3jo9/QvjBcxRSK+iXMoIHrygLkd/59VFZn51t4SLIXhkJwJFnU4FR
5kxKyjM5rs+1uDZGS00y/7xs9hBiA7AVDfQVgMfiw0lB1WnshmZfzLf4H0S4T9Tk
T6bNEpizuiv4r4Sm6vmfRl6kLFL7XfwzfVAmEMAZBeKV4JR6WaqiDmhqwlVHBS/O
l5lWoO8mT2nDXrDi1xN2qXuyYYfkf3q9LXVcsk8ct/YgfP5jZSNI13PUjii4Rs68
IY2CMZBggr72E4QwPPHKC3z2XyBBOuVoBpa29JplYGl2csnBOyeVT2KXn/RQ5eTi
KevDeRjrKRd5VDHKHj4HOIBLGjINBj+oHAYfgE/IO5+Ec6m5tcykls2XVit5TyFH
LgjWv+wsIhzTkPy1KSbYOPMrbe+EDcxEtMV/GTf9bkoMn8eOYtRWd7DOT3fcOiq0
GjlwwRbPjl+S/k/ImtovZx12lHjdgqs8NE6mRyLkPOjd3OAjUj4NI7qoGnGZsMWd
`protect END_PROTECTED
