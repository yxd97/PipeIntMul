`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FEcA6cswpS7eBFJfcsWQQmT2unxHlvVQUpaUSi74CayBBmgRQkSI5iNSDR1EVKpg
qeZlm5B7DDRi2mhmb/2lJgP+B0w3AK4AOdjhvaDOAV324abVS1tyCMHJtEttKJto
18CgqVBO0X2Cxg7cchSUJx1IcZF/xRFApogZ5BHcP6IXmovbFGxd0CYcZJkTtzm3
Laf5Qo1NpGDpW1mgsf8y3au0yYElp+sfqALdWGZ/MmI9CvVgsXzXOlKxJAUzwU51
3Rb7xKS7JZ6woin2rJA0ppJIhYc9xNkoEYUFeocF++R8jFBQSs1N7UxZ0dxQU2Uq
+dKCn5jfty1uV/jd7KSRyVkC0hL65HPjwkN4MUkUMHo1Ln7+77T3WcB/ohv0ddXZ
X6lUHAx/DbEXB20g+vtclx5/jpeINkiqUHMsYodNCELvKsm3e5gJDYWq90iK/gBB
I3ydmynBFFxtSPplguNmjCY6i0VzrYYp2ah8S1r55QHLxNfLYvLiXKUn5wM62IO2
3OYT/nJDrvo8YOQq2EJ18uow7XKwHaUeLGNIkNrJgcosjyFucKyILyFtrZe9FmwO
ebuvHe3C/cKB419YHejE9LNFJuJroPDny9blXs7U73HL++SwSsqch8/+IeqgUGIF
qc6oHc2nYJ5xruapcJMb1AG7645UPCYKqe2VHGvDl7tOEAK3N9jsCnC0sS75RNp9
GXsdLMF4KkIT1zfHIaTVUb/Jhj87MzUwzBYwNQ9u6cmby1Z+m2mDlgJbrZDW2ZCN
gahZx5OLj9xhziBdj/ppu68w0hv1VkmsGHVO4qTsBnMaUAUlz5l8t2tRl6g87vSm
I7PXm7LtiTF0//4nXYadkORyEPqUNf7aVcANw+XTUzBU1tly4c6GIo6LgCyQNlhm
aJrPaD7blLJCiMVcyefn6TCSl0K8OZ6lJAkddLKnqBVr1qfZS7u/3cX6IgHhiJgz
4oVjGJrOsIbKFWuOzwtaRhC/mT3GIdmWf54qzm2dHfH3tDi5Rhx2gOR4szXDlnV3
ReIboqPCaBlRUFUo4IoiuHWr7cGKLMmTA2l97lhfLhsJcV1D/1M3bZ+zaBnaSjy1
aE6XcfPjMCG5RESMxkWrtCrz5cajRmg7te6iyyw/ywf0m1Gqoimn54IPsXjuyG2T
8I1bz1AJXDw8FjDFo/uYcL1TxBxPEgrzxU/8nucaFZEJ+WO2EkkI7KEZYI/iDmuj
a4spYUOEA9TnAT2rsU44zm1lyW2n1UkRfYHCaMvtQAYYB7vXQCNMwDBXDLtk515N
paBfJ4MNrfUJlI6ccMKRZ1fslex9O0fCems1LApdvRZCOPIED3CgABagzI2+6DJM
d41ZXmWHa8WecjmgPr78BvhohQsTIK25tXeq0VGYEEllzUmIgUySucFNUs55Oglt
sOD+eRw09Bzv2IwIyXsoz/LUOI8AuBUfLflrGxkv2Vh+iLm9HIX5oln0r4+e4Ez3
gDRMVMALoT20WLCdySfNhjZW8M1/0ZyckE/9+uZsYFKmCQlORGdQrQ9n5relA5s/
jXq+DEnYg8LqiXKSw1YaMvH4uNJobt6pzc/1LBC7T22MX7MaLNaHzfIWNCFXlkBR
CElRn/vai7flJ6fxy9oysd6hpo7kEUzAKZ5wIxG3DFll87ZAIHJapaMa8PCr0iyA
kO0UOc28lL1MzNBoboYy39AVhgnun/+GoM5N57VyBC8UXouIBvkj3lkpJ7PvofR0
cIErnVZTxSckh3pq0DF+NzjTY7gb/5gvCqewTHnzX9JRFVaeK/kk0oYadwBZvnkH
z5J734DtcOnLwm8YsOuFy74lv8Dswi4UEbZ8Vi6sLcAXIKTOiJGVvHa7n14GmiKo
p/hMgOYHxdFRuxPVbHOe2VQoJdRU97L/CHc1iiA9qnKzYRZ0AoCp+NSc6VIryKmq
vVcgeOrGeyZ4mzjznV2XYr8W7AGIioEX2GB2K11Vy950cyyfn5yCk/d027XH/Yqs
MnZA/731YDVNDDvDaLHQIyhBrLt6ZWUHLcBvRECdnSPCjvOxrRCEPtgte9oL2C4i
jV1Vhwzgm25VJV6RFwybU9wcXDi3362QYOvvtmnrM/9XQ/TkNdorfSldVa04MAUV
sRgslyE8vIXs9v/6eNSl7iYKVK2+EJHrEBCXdhQZeUFtDUIO0WfbDYD+Xlmn3Zzx
+VP8ItbasRgQ8l7RiIPHXG68yWK7VsO1q7b4jMw2pCTYypXcO1Arp6Av6Osh5g+5
HNUjERMpnfYYvmyi7+lXOTMhYe9Pbz+JFZKNstl5Nesgtl76BoHlz78Ru7iV9U7B
K4kBhC06M9ohWNNNvHDjPjCfpHVEXXVNGnmXBpVaQgRjQroZIoJKFX8CMYuMQfCW
HbUni0w/1RkACebzR3O/LunWCQr035jMWWb+FUv4djQRfNftY8uHCVJFBqu66M/S
l8YLttBdAmnSpLS1v40hQyNkDOWwEpzLXt9h69oMewxCqxDN0nFaqz0HZJnU4q7Y
R3b2m7aWyOZMGmLjaRA8hmcj5GGyyMiQkxds5LYgTNZNgsx2faVovYnJPGPuTX3R
76LkMS8PnhRL7jR4ARqzth3ZLDM6GCj3tUcu9DaDuJYfu5uP/07u92Y/WnvDj/G8
H4rEDc83hPr4tN986XHIKt2Xf0FSbNH89FMufTmd+/lh4gZ290Cza9NsS7IZFjuM
88A8iXBbOdC5blJYG2zyHd/Mx1ltNwNCBm/er5hxRq0KoOi0qHR+SVXiyAMa+WSc
Ub87Texdxett8bNyRrIO9mX0qZsNAuAm3q/G7Un1/n+mJwZeAak5kkenfqIaA+vK
mfQVxbGsHISVsZ83X/qQCUq7aoMUraKlA0THUFV2TsalHP1g5//cauPJv4AFcXnO
GEWWuS0DDUGc1S7GbUGUI25X0Lpkv1NiX1nYqvHws4mJ87Fyisoj8UNWB51Ty2jt
Xpig5Xi1MsvrH6Ck5ZC+Nmz/I2ZHmfUVXom56Zm+7H4BW5Mohzu6bVP5K+wVCVww
/8RAQbAmtAbhk4ptMMGw6TgeEQSeIdkCLZwP+z64u6hPgHr1qnpa8vqfVy+SbNsR
afb64mqcbPy6TJoJLgnAjWr6UaNXtzCo6eHh0Sx4shW/Yrd0wL5jwuf98fzT4mvs
lMxlnfsbCZqhDyUhcbkUIyWDx11zZFxveBhhnpMVtmdKdZHY+TzrE/Sw7RUDRjgo
kisfw/dLSCEruqhDjOi9PN2eu9Oh8c/l9peAkbapUUZIBfkzIM4kBmMkQKVvN5zQ
XpshzRztHMKC6oKgqzWfZkYyU9hstI4kRnnJke7iRjTKVUGALLHNPtIQhoWLRMru
ENl1t/aA9FX0jowUc0qbSmn5U3M/GDCxAN1DdPkYAr9l8ux+rcbFK4mQDpW5xp73
b3zzjlujrSxYDlAnwogs72manrkAH5q86xIOHzL04GbJu1cGO7NRLu8fMDXxM4RZ
f6hYIU951IcgNjw2sPVakbrgtHWcwN35J+OQaAqMB11cR4kvjMZZ0R3O3FGxDI50
NBmAQHwgV20D2jZguOtUBVY64Z+hqew2P8gVnxKX0SWAjJoAwPghL/v8vkANjfbz
xc9n0v+ofRf0403Gfitfqqy82ZAjgTHT/pEyBoFb6kpYzFwV67nniakxfR6I5Xhu
J2O/zPVYYpuLo0yJuMTHrkj+wWTewF3YDYw5GUc0WKNQ10SEdAHOcNVlU/6Tetwo
doyrqHXHXTwvyd/aBxNjpKJM1pbbSKuB+nN/z44pL9Y+vBlQiM0ScJ6DgncQ2kI5
uqOEla1rVUNkv2JERP3ULCVvdWboGuNrz6PrsXBwWdYTVNN07bI1JvHEke1g8034
sHYujvbYxI6E3nxL7vCGoFC+HNWGVFVtz9vXuMZwyr+rYy6PLmUcneWE9HVdSlrW
8Ot/MJLEmR+CcI4XaKUgFXZJLkOlr+f8L54VpaNJ+MOibFcZmxR6ikAzTWS4FOeB
x8hhpW/ORFpZCvZ6/Yob5EyxQVrpbr8cE/2X0bhcpgZNGzco+1KkPTwkLMzh3r1r
0uAy96yv/DMNXGF/seqesIMBZz47CH6F7joFndX5jkJy6+pLl5dRqdrPGKXqONn/
73kCK7Y0Pc0K7Boiq5804Dv6203UENZfCYbIh2LHquUxBC7Ap/WL+9ASp/t5fXR7
jxnRn/bDSmUAEKxKF4g2iwKxHJCY1+2ODHNzm0NqMQjw1pdKVPuDhvNYuBZXCvjr
AZedlhUGiPXAS0444FXGhu3AOLrzCmhOe4cRCDIy7ZR1esdr1fudhDJtJhm3aYIn
2GrAxoIfCLuCtlYkl5L5NSc3G1VPY8Xxiyz3HtQM0fRaS9hlWGo2owjUAlLirPXN
m/LqIi3ntGPWa0O84aMcLt6RnxVKVQ89x4y/GsHRPhPloJEPv6VnyWpCFre8Rhh9
6qNdSH4IKkCZOxv/MFC2iyjAxFwXlgBkAz6t0RKnjjbVHIBVUT1ZO+QMpdhAdkKl
6zmt0ERcZhz5P+QNihTsS5iYkxQ1BTWCsVTSuLxQGWgGRQm59kMWkw07U8Ab3U33
1UBaGa+bWtKf4rTi82ot/aQbwg+UXG21hQjnlZeJNRbEz+KNd7aFTgQyUTZDOa3n
HhkT6DP0Hdbyo610ZF1vNgQxAMdumvXhZAmjum9GSsw7JtR4AW98u9KEPnbobJwd
mJqMN7O9f+t2EeQaWAR3gjrcZSPUH3eeZk1x7jBx8jKteRsqNs6ST1LOcc3V9Six
91nz5QE9k5YNG3DTyI5eduR8Tj6T0HuJlUU1JIPVezIwEKtvOPHPUp62RmjB2W+p
O3MsAF0RF3cS2zs2LaaNV3CCMCtcUTxtAr7UCRBVRcCAaOGpPCwXvj8+cqyX5Y0v
9JlV0eBxYOKAjZNK31uPfwKeQD6vcTeHk9JEhEuEaLlMSN5pMIcKmVP5q77ypBbL
dt0bvRKkQj8ZesfntnVxoabYsLGOoXMmV+YkHe1fDFIe+GevxDmCXCfPIHow3UVZ
Ou886c0AyAzSFBcuIbYspNVQYivsk+y+NM/mpVrAYBeNGsFpKl0b0FMTv8MWg8ar
lsgqBksxqtFQoOkFjd+nN1/jOWxTmWmn5otHRvgbzZeqjWsvOxle8CUXsxHAZ3Rk
PHkf0HejE7+OHlSO/OprBwqpymgHyPhpNyICqa0ZjO8oHjtv1wrVOgfQ36hHvTAQ
MNm+zMG+gFATFM5JhcodAVqAaYp8tyGAMn6rm/9Apz6JkCA9jlRdPpnPK19vJQkz
97k4Nk2HiVlhxVsu4cIhwCnqbm5duHn+YH9+hxpYry8IdAgP8Uvf87GuJn+kTfZt
LttGyNRNj9I9ns1IScFR4a4zKrEf/2251I+9DKnpk9ktA3HrQYPx6sG82iCj/AI1
pZGTLbY/Rx6eIxov3ELZ2bK6DMe5zPBAa+cNgewk0QaMhJVjDbn9PsFYy00eYYMd
RbC/3mq9H3ek8uFbwcIJ2bVJ5t5GMFrlbBmqvtEhqFWvD8Rq8pDf1N00LAwKpsR3
kg0rknvFqeKyyRoVpdx6LUFdZGRD1xpDJSW6wBrTDeKA8J0EyXK4FowoDKTE+4zj
tN8ZV74e/lDRcz2tWDspfW0E8Gq19ZaJLJX3S+6kaRbrnLLtKFM8c8PsUbOultag
01IElDcjsZ8cdc+3bGyabbUDD2EQRoHOFpN++1uyoB8UFHXxLAm6defrKZh1j8Xt
xq5AwGlLrCLQnC8LwfSkJEsiydAuCdkc1Xjd9IMAPiAj9VXbOZMHlcXTkuygO8oE
IDJQ7zII43d3HfI2DuKdMbA1RtmDgL1EXzaxFIQpvBgJWrLRfqw76rhlBIFE9mvT
gXmZgevWFGgvcPuYlqKTwTmso2KfSPLz6kn9ng2gfBc/MxxUc93xkohnj+OAjBPj
XwBvHSOWOYfmI/Co7iJySHZjv6sBpplFZO+/Zq8hPspOXMPIhm40MKXNRkUW21Fn
couBS7kd6/BPmQiszdhx7gx5Qe2JGTbI8LB5H3MczvXVbcX2Ei+w2+9k3/4ers+r
38Q3n5LRv5c3YzR6klTzkYETSTojHQEPHOTZimkP7BDftZUu/9V4BDNI7iSnBvsn
xNZfQUxVoRkLXmyhKkyMJ1TB4KyMTRhHAnQfsm3lK4FOqNTZXiRqEUCkTCW+Q9hu
ixHF5TdOwIf0ZPqiIjoIUswwXGbuZI8VffdG3A4kRygidk5wVv1X0tusDl53JTjZ
MDxVdIv3rd+mrFcuGWE43LwyFDMdqcha56DqnHIWAv0uahXhV6dWpmc8wwuFnffr
OSYalDVHO3fcJ9jkIAkRvYq9O+mvEPcAF3PA7jiFZZfY/rxIChhhq69MeEziBnop
vbW6KcWdSZYHwMVztao+PI+2y8u09keGHYjvmWI2Ltm1S5QdUSlkdPKL2FARIVuo
UJGhTbRCR0lNA5hmUXGYUKJ7TwDg6oWFlj4YOPAcWs0LqqhegrtVc3D5BI6avPeK
0lNYkRjUFBKKvvGIv1XvtvbBv7ijFFmYgQIhlYmU0ubHEZRzd63WoGdubyu5sKWp
wmBCZ2diKJQz2+R/3T5A2c0lWUm1vdaXwrdCaqMY7k2Zuzyg8/NrmDgdSK+ylraX
KZ3UaMloBytiK0zLVaTV2kZnOJG+UqZugOf/uAzbB/zRN3O6lSJmk80JoeWfqwH/
keGESAWRNIS9k2SX3x+C8bAuHTy+zMB+DfMvje6e9QyfZKkZi0UDJPGmLqOd4L0l
Gv45n+24IQVsxHAFXq896gl9l+SBxsP1Q+K39ZQ6xOcEUcg1AEBEAiZf8NJkzeOM
Bk8jE2/yZpnhyaFszvgproyBAE0RTbqFD36H61nNmwiOrcOOVfV+FqZs/coy33o5
l0O0Xev6sG8xas3zm+ndaBCRPNveO8KXNAy3UOEf3oeAw0w1FBYWD4Ksj6gg3R9x
NVRYQetbQ8JgQGd4YEAkBluY9tZdhp7jnM4czbwWP9kb2jZ5hb5+N6rHKZLZNJGR
G/MJDOuUBeVCshEuI3lGU0tJ4qhrcR3p2Bx5Ftb7h2lvAjB4+ju+5fW/nvHzVlsi
KLAXFuYf14oYBE4oHVx22xBnIRNX8bBOoqPBUih0qLZnsrbiitsP7sBHNFCvyLJE
Y/LeBoU26SszMrXQ53zrut0UlVUtht3T/DNK152vrQlgiLVxoLUoIMo60fkvE19w
WaO72AXyQyEeLUaUTTcei1v2gxJc8c9cNRDq8vSG9tyE/Ar7eEXkPktcuqLYRXwh
BhgTOiqXTXEISXG6adumV+jdKimC96X3Q1Dwb+nwvKs1r7IZ3I4PFxCzNMTqU8pe
dbX03WiRFwz7uRL5lmSe1t/nGeaCJAGQSEi4xdFi4jYuL8uwrHgtkgQCbmkluHSx
B/7f0z0mufqgg50U1lvloW+bt1W99vm5MLN4KIttdsB20qaSCND04MEk+/2UXdg4
XzhriDW9J5aII0PY4cTpiyTtpHIayis+vcKPLdrtdY40n5mlhGL9ciES5izSjMfC
Rl735Lz2dnHtfPkGKBBIzqZWzNfawaEa34m2MKN8tdOcqAZZWv2HJ6cYCyYzsgtG
YVs+9CSdxuOwEob+U9vzprCY9Onb/2nLolc5I6ccDyfu3uewUggC/HIK/VS/foY/
YYhh66y+hjSp3BuW6Fu7ooK2oZQK64avqSDFnZLC41y9yB8tPWK1/hw1EOz0QzkR
cxxhOXK68Q3K8wThBP5ywxQx7wmnUNOfGbYvgmISnlLabUZbqolHWVLzs+vn60hS
ao1bl3jzqBosMY+AN2Tdwtzg04YnLwNL+WuC0jgOWhxGO5IAsWjxKVZUFyL28kvP
JHzsN8prs6S/DGgb9Oi45avXM5GWl6Bx/ftMaZu0BP+q41XotVn6D8/NyWkTr11Z
+h/lsPccWACWvuDrtV/F7XtR3Mhap0QfLGuxTFd0nfVkSEn40WmgIrbctVtmJazL
mCun1G4XAwnTP9a2Ju6dcDjSXSsBi5iGvfCSiS0eneIELKqNqLgqzvwpeh0ccJf9
5+/P4U6EEk9OtdVnLOxhehE7wV7DY7NyT202xFSSAUfptYLKS888NAwO4aP244HP
GOUAeqzj91l4+pXSxQVt072mjQ5vsxJF24C//pIeQqTReesKWrOAU6m/6vNeKYnl
2Cab6OVeSXkIdWdkU8+jaZhFXPqeadhsPymRp9waRmt1g37Qv9qGIHvCDsJNUIN2
a2YI2gwFrhBni69lhLHrmwbyfjso9YUK8gDg2XYVAY7fcndtYP/RbgFsYr/xvxa7
hamZqZS6/AIWbavvQ9+TcXHYlBH7YjSaV/2cxBROPJlDW3K45HRk3W465py9yZQX
hGiCdxu+hjnIST9QeQ056kgzwwNzVI8uID/rRV/fo+lvf5iz0rcu3FdUtlZxAHDV
8euT2otFUgUrPPint4UqR9VMYBZNYj7+3ncbrMjDtzwalJX/cX/GmhWQaKHc1ZHo
TCol+FTDZbzroMeAKqgUU4L78yTBarFEn6cmi/p0JPwtwW3BZELrDqiukYWwFqXZ
CbVr8DgiJBGKk/NPt3gAJGlOjdEl+RSnnKzVQHDJzzxws5c3VUq/XRL0t0Oivj81
Oux+wS96p7C9JpjFaBYeFrvxJVnw2Lq0JetHw+XcFXqDJTEUDt7uw59wNabSfaeP
rD+R10Qcsr7uihDe3ADixZtDeb0dM5oVX4Wo5h05pH5thxdBQriuS9pl26kVHYUs
YytOA5EswGXAETcYLzv7HpRW1k+cKo6swT1vw7LMjw+EijBUOIh6sLMWGC/o2mk5
VHnjghSO4MwhQPCuypRW+8J7PGGqQAi0+9fNhtLXGV3qGdNTQTsrSnqZSGuTsZFN
nqYdj/Zp2EVMx+khKmp2o+XDk0ZjJrepPrUL6apvxF+KB2munI6ZOozQeafaVLjb
HZ+BUCoGA3m/znHiMPCT233Lu/jTJ/sZ1VN7Y7AJrimc6FCfLRK8FVjH7XXJ5PV0
kSPxwpuejqN9zo5EXg4cIMTxSybu6Pjv7+0mL0mCXUNbIm1oLGt5+gBJGzt6C5Sa
iWdJ8JLiN8RhNpBBaF6f9HkVyh/fbYYIzUC6FD+IcisOX5K4D1njTT6G/gYJtvSh
oG4Bx/hDjF168Dt7B6uYlzbJCDh3ScotIx+qDf93ANFGQlE6CWEnl8kyTbxAqMDp
cV0ikJALZuAL+JWTPn6RVUz6mh3Dt9dzPjoRSEUfE0wTmEElcHE2PaW2h96Ysm7O
PfOoCc/FC88wo9GUGIY/rrm4qPTdhgjaWIYFRInfVzlOj51VHPpnmUU80uYoSRos
ojPORmtKhbxXAj9f156OLbQ3nwhLSx6uS3P5xQrbI9Ji3W96nHx/rKS3KR2A5Ius
W1xQLOl25595M8qvGIF22BIuW40/wdk9/LHE/gCmGhmo7EVTm7hhTzDoFrSyS3uX
6Gjoc+wg4CGQjF8XqhDaeaA0pzyDuHBMIztvt2kytK/ZVd0VuncnZ1LSlwqLeVLt
368aSBzJP8wYiKz3FOkGv5wNyZbBgcaGYau7KYlGzBxK9URdvblb03eTAsR60N/w
Uxef+nVy1fZ9aYGDMDGivsRz10yaVs/qpGJXuZwGdTgfkBokt2LgsL2MOTvdKx2/
zpRq7itKhgnKYHj2c0B2rAgHg0JUUmt3faa8o/zonpIckax8+LPswoMpn0CQ63tu
7vQKGZsRF/PUZKLiGC7KgPmq41/OKxImpJFO6gka+7BEcENuSYNONkpFuI676VrF
kDPUC1vXnvnxhmzWIcoUf4VFx2O7/aTzYQY9PqoxKyaKeqFGDBLhwak17XuEJK8H
Y4lsiM0W2KoDSZ8iLJUwpOIU5d5W6GR/5QSAZvdn+ZyYxDwgHDJ9WqQqde0+LbDB
cG+wM9iYN4u4sXw02sIJu3rodR1KqYB9ANlwdRm7Mr1szKJvopj0Zo7XiVDHE1S7
2UY0agypJerj4ozGNizlP5XrgdVm8+liuWL4t2dxUJmQmkwD4fVUScYVrqKMb0X6
wBUka2GormXr4L3Ol8iPc+5+wBxvCyRYjop0Fo9NsRl4+fVA4NcA1FitPiVDvDTp
/OZN0cqKfyiC3DNEX6crcVDfa8gnHDZvUvlYv+7J6xfyLLVA8NrXhRYKvL/2/gvK
f8Iqw0eCG86cgoWACo8yK3j+Mw0tY+Ic1xPYSP/vKNxjz9COtS8zHuEXPp7zb2uv
zzNsV9RjnIde/aFj/BvuaHAw1TCvdj4JmBHSHsoGwfyIw3+fcEXTc4UA/QT689Vj
DcLZjaGJO8k+21Kycqlht4tbvQ+lowHg/LCkSxqHbX3UlV0Bj0tEipy9pdXzgrB3
uKMfEt6BV6ERGxG5sj+hFCf3IhN2VXscedd6LZkW0+ZthZFJmBp775BI6YisVaef
5CVQnO2uhOK09sfIQOqo+8K5iShhSEvMJJ/MEPZMR+sx1dkXsOuBFfoqpGmXzBCW
gtJ/xtAqEw3GvDnM4ep53tQihCnXQ1XttFFnPBlqdN6qgreAyCkB2JibyL0ysRAS
N93LMj+c1tNmXR4CAO6X8yqcl3s60Pg19PYj7w79zy+sY314wlKyebaQEXCcQV/0
cTb5Ts1COziwD5WzDpd4C/6a8sMGL3mSJa+Luldf3o1nOK2eiqkbMsugFRSFrvIn
W4swY0CQCwzk2nVY8BCT94z9S5NMXZ/U1H4QHimgpW0zfermVvo5JItq1ZHXEV3I
U+EsAZzH9BVWfZVe74Jub0xY7SsEqlYDVYk7y0MMevmL5c5guWcL5h/69Yeq00f8
OLXnSPVf/eNcznPXhWDE11wT1weEWA3I8xoAipgLHgXoSZFpufllX4n+HYo55/Y3
R+i9OA9QMBzPEcIqCFTrAzh+Lr4smFwS3qR2Z7YTu5c0NKxIUqiqnIFQEqEoxuge
sPtXgdA6yrsy8xa7cjyJ/c+pGfhuH0osr0rBcY6Yv40FkJSF0V4cSdj8tQHTE3B6
pfHOnVps7KWVZhTN7S0rCyjecvak6sd8i8QJnjT3p8rsJz8eZBCnuUQqMYzTzFKt
mL5tvFabvhMvBnVQGQ++zYb5YuyH68CfYzN/KQ405AExml6q87nwg7eFUSQQCj22
RlTvrzZfQ3zBZERDnV6OCMaPuyDESR7zeLlzYrWm3O4EupxVGaIbLO6SgPQSNpvR
zkbPu/uJpyuzSMPderWnGJt8pM8NsVunt4fcbD7E6XM+TFQzgUIefOL7DSg3Henv
EK97xgWaXZJSeADQ5jwFtfOsigWMOvm27l0zgX22mhLFE42oapNiNEtikDSq1EJJ
cT/38/bVfPxDZxNIs//FNK5nofKewlceUEH2G5VPFg1jBiUUQ1jWNne7MEvdB4wJ
jwwoAuMlLoYjwhj/GaWGnep93GD7PIwCyJpzPL7bHHejs0pwPrffTDDLdv5ij6B7
Zr19pmrLBcfLrbTjiGa+Adz58rH37xYRKB5B//p3WTqsyo/IP5bnhYO5nZI+wE/D
m4oqvU0/BkB55Q5iYbVoEofcRgYMrcKD0ln4VmTS7S9kaBXLKq77gkEY7XWyRH/N
LvTyd28M8bw7ytjVZ+W61YEVxf1sTVvGKDv4aICuxnt3yb1BUT6K6KHTQuMg8FGs
uDagV9AXsfzOf9Rr3ZksmZ+o4lJcGkYI5QOPOHnm9AAqcq+d8ioNvpvCpTmN9HDq
chDTpPQ9q1p6T/mmGSvwSgSp/HTkB/NIZivJ7US4RKlSii/i4jUTl/PqwcPwCW3g
p3AAwYwpDWK+HhaQtmk8Da92w16kW+sDfBX1MpQqm9QaJpyg4b9uJ7FAtC6k0e20
MDqy2Wq+L8zWVe6feLOoHho2cAOeEhpjxBJTnTCry/OpIkI7nhT9T6kKPsPoifXd
gHgGsooI12dKMYTYdQR6mzg+qJ/NSGhSPW93ETKN6ZqEu3jmNB803mmaBvljtCuh
X6PLeCGDpwqB5aJ2IRqw1/4EayvtFajeQ09VKYPDGDS6axqPTSxcmUr8cKo0v13h
Qpyxs8ljKEOLJ5hf2fnEX4LDDSXRI3+AMCcDSwI0JNf4J64qEkvJuE0NcmRFZc6f
fm7HT6JHLFmcfXtscaOwET15cLTKaSbYe2dxQVX1JCjYsnaAqPeb7YwMCOaziPtH
STp8PbWoRua63TlAkon8FptpkOkObJEiYRog9tGSsJqnkF0esW/sUrLLCIydPCJi
TMXgVHviFIlCGkwrXcoO2/eDdmPcmmuiQBEzFmgVFs/pNLbDLeYiGAXr/y1Pfunv
5PEzpxTLWVFx1Qsg64MfVuXyFhZXCK9JbR2XvbqSn9/W87RalNzx2I3BC5rDOlTn
F8Ks9mUyF8/WdbqRxHqHKIIKWrNuVdl0h5fHq4W28pRDmv0ESRkezfU7CxfSjnKr
DiH5uDgcyH58cekmN194RYLJWEn9KTnHJFlwkl/kRD4AqLgzozaG7b1Ltnb24cVY
uIB0KTOdPgEeND4CfiLNmo//dTCidCaVo2RqM0mDJHTC8LJO2FIqzsj+ioFKmGO1
wvjzYNZ3YRCHlsx9ZIRoo4h76F9WOU5zMYUhvmMArOZ9s5jYQXFZYwLsyx3wjbFi
GhaENmR9vZQqgRNYjEW2vdb0U86Xa/7zdXF/6BlIWBw05QsZtpKCmJYsunh9BQ4i
CnILFo40ng+Y9q/3bWWwvNgQ0cfR0NBawlYUal2KnriCMvOyEW/yjHP0FEA7WMy7
8mbvSPpiFjtwZS+nMqiu3iSHGwfblZUGDbdRU2+Olnc3Yr91Hz3H4xHqbOezV2qL
gDtr+V5tW+i3lBsQzoUt6MpIX2Nl5lPjLdQHQMY9jKRtdQgvAP+G7nYFzCZtY6f4
wc97hCwyRJuxFSLt9CwOVITWpBVQZtM9vt2kMJwm61dsbhZBwPRRACVJj4DTK/Y9
Fff0Etl3P7iWeRxEwJs/KGKMBOFgEgVEIwtumZulLpPphFLEBUn79lQ8RmnhghJ0
6j0j8YlmE1IIbXb9tEFYK8BDQRuM1Og/CLVWSys0reqRPE4FNONuoyDIbnZhC5oG
G0MuXeit+Hs0d11TX+OwuDznjEjl8n4bQ+v/OBLcMY0OfB8Uo+ZSTBvhRKb1fIXu
gHFuv1uYwenGL/in2BQKCCVx2oObPsEpXfAxHUrfD/9+6/MxGL2dcZjFwlla9tXz
U9LUiQKKBGJb74RWnc0LvH4I3PGtGftV2aZBCGcnCXwasBcJLjcMec9dWiRt/+Fc
iOEPQLMpGynwe86UAChvKE9ceyfVYq4MY4AvBnVKKD1wQwUq2IG2h2f5zPpzSIdb
OTz9fpYXai5aXUqjLoYvqYxLvIL/NmBdpPHwqFVYWBnVEXBiSsBPlXNelyav7D6N
wtCJX12V0mQ1XVCGgY2yWMfSKXFiLr3kUCaLZyCzB8LV4osF2nJZKPjw4lNZ+23V
Ry9UTflc3xLZNglFt0umJAAwUwwLQOF1ITqOHa3kZ+D/MEpeb4EuBF/KwOhzvA2k
cgYnvL7aEzD7TSHEjFNvaP9Rw/Gm6zawu+qX2XuWF/N5D99+vdN4EwnSjXqVZVrt
JqTcrHTsh82CbDTltk5j/PQU6vsuvcasp8TveGi/dJoOSJT85JKyaFzBEUveA2cs
iSqFl0HpXl7hbNBcjzrULc/KpGXHLXm1+vFxfzkZACaqNmNQU3ULdoB/7DUSCGBY
wTJ07ZUGzEJyX+80xPVI4O49XEhZdl7WEPiGjnu3d4IPBDGrWxMaIEfYsGkLWfGW
XnF2RJjP+v+QDa3MUj1bXqzhEvSwvCW/SDhg2Sxdkp8h6KYmaQLGJswGE1BG92iB
nmSYscHrVHauuWXvgoLW+BXxUnDzjk6sauCQKZzcek7rDTewaPLyfor2cvTQbmco
/8qRy5U3+3ESTvMcTEZtbY4Fa191esTq1qtbRXGz0FMSY9hAthtimnH4Lk9SYWj/
FmCVN/yro85PiWXaxTxodii4zlcLI1YbtQR2B0JLGF/OrOx8nhySOj/najvXtQ8H
1gKzScNWoSQ/YtZA9BhCD05i1RsTaR9HTwCuvwjrXw/vHvWak3NvsG+LJ+MtDHfO
VhBFPX4VCL246+CmsDSYUhiBAFfP3q2ElLPJRYgRdor7febn19ZCcn+ghuzb4e1F
XO3Bgthpd4+wsd7mAuT+gjJYC8kTijbVj3FvlUurTJZyQgxZQN7SfBx8biC1pE04
RV/6F+nFK5GWDjQiJZ2HaSgL7vAbHgSLj+mo5DO+43gK0F+2RfLjhWi/HRhvGje9
Bzkz9DI2MS8fTMOXxXvfVB6EZJGFP9WCycxaMi4s3BXGAUjwWHULvo8rBAFcS6Li
+2ATz0XZhsYShXl6vxLleHC/RhSf9TN+CqC1PwF5du4lVtbz4Rzs2TscBsQ+++/X
VGGN2ICnjGFip7HIkdoXTFB+WJ1gOz3ivG+rShCb6vuzJOHL4oLEDdSXIbyQDQo9
PmRHdoE0A5pkI++qgZiG+XNfb9PKVtdGMwhHgRcqtjMPu4Ecik9LoQ6pLKdeiWq9
BDarax49ArPwzWU4xYNz6jiIuvpnmNvU2eE529jUYA65LsPa3BiTu5jGe04JAPgQ
WmhPHGxrfLaoNGIyLrih/KM2Dl2wcRH3up/4zkwJKdus5jAolBklSW3wjXRlGTqn
Uz5D6jH7egRff4DO/BiF3lm2bmOSlK/InKVLF1Vq7i0TOGxoopACb1BvjOANNcBh
yOcXM3D5iQo/ZH/3Pin4saCuEtZUCfEtUcSpnQ+mhpdHeGwYVMbYUsXmDPoGyoaZ
vmGlth1jRfElhaO7fJEjexxOMUUo0DsiHz7kBK9jDpwJ6fS4Z5LDfhoEamwnSSZg
1GTamjfEVl96MbjjHZl19Xq4/wc7/X0LIMg4x9aavuDHw/LQZeUyp4rsaA4d4Vmn
CBOA2q8R5+mczP5AaXroc/x5adwR75g6LMhQiylqWGLi8BTeYKrJaqYzHNluEO8S
Lce0tPsSuZVFgUJb2qWPyv97MA3ID9SaEozk6LRyh0zCcr7oF9hMBa0arxDcpAtB
7mFE+p2A8MK/avSw8qIJkBAyTcruY1B4PX9QXJKl9+kYUpZrmgzQeubgI6vMS7lM
LUXFJ1iOGKiTqsFDAc/7i50DlCEDJ7yByIyv16HcI2+V0DSHP5NoWxia39OODqyh
wvaNf/o15/85FxJH7L+Rs+aWbT2W2cmLnccOZz9ghsgyN/L+UdYd/Hx4yWAqB6nW
RhBhouNgjf2g8pi5jYYRteXjKhNWjPJL31RCcPZPq51fsiADxZwT+uXj1p8lRHr9
+/jfQRFnQ/lAXM3BRy9UVAW9At+DwVVfrUIO2czQSyXV/vmDQReKQ2Y+MI+7SUNY
9u5DC63JX+MKHs6c25SGRwFl9KS4fw4lM9KblbqJ2FeCuHBfdgGkjR6qhiw3dBDH
s8Xnk6mun/CPSVOI8Jqu6RRnfl4DwZcY0fxX2pNvgjvqp0DZNo//KmdjfO9N8Uit
YJpNM3Dw3whm0EBYT/+BKL5Esxb6BygEbrWUqLuy/z3eeWB3rw8wtlJk/V+qfHY1
Nz7M/SkcNgxb/hn0dTAi7rV05bZLUdReQSsJCgJpTiUC+vIHNs+Xhcg7oKb+wV18
MMvrbmMZbHxCzUuVjmIeC0IJI235aGyaPPlepcAGRmT4tWk1CgmV6EZKDhcuBR7B
CI1BYMtF9M3870JsiU95JPn38EWIfJin6N8hp8VhpPfKdt1rdZ/CrHdV+KIiERiv
A2DDp1nyjAasPo+I1vW3uBhe517c90aX3+fkWGQgBQcflSjNwUSC54QOSEAGtj8D
QmjiYhsJ6X19mfRLDIAxpnmPJ4w3oHLkDIclwnMUUolTlBIeMQ5iCh3DDBpfcOzG
LCAHsfpbcxWOW3H0YvJ8CLQCfc8w0mpPDJEfiny46DNByVN8CYd7inYOWKva+fjL
TPORtp+eKcKtj2AfQlnRDpjfYqoZ9mw5bM1qEjxlwSZ40212Wa3HFzbWSwsklVkT
4/kijbMib7LBZTO0w6CDV7P2qxgGYTPnBMRJwRE68x4j/l23Yg6vGL2glV5U8koH
V1aSARFk5dUOWtKGj7Pz8jusyY4l+BnNbXsj1xHMVOXGXBLSl3Ut55rc/TqJX+Av
1VcPQ6ezjSzpbBCp13hdnWGzzOotvjAriDm/fI/BsFCY6JbOBZA+zvs4nzIPZiT8
O7KS/exX1V0oa5rZhf0jeLVIoa8INs0sw6Fc0PS+MabGhs/CBaCiYGkPm/dGFhLm
qgk0Aadp0tdgjJdXmYV8fgi4E6EcIBTRpHiAPezHoJYRsjKuFwpco8HjTo8uLBGJ
I7JCiOZtQaBBvjq2RUF+2OVh6IqeTnZcsQE3rWjM7KnGr2du5sbv5EK4woIaQNDW
0E1Nbg3bsBq0n+nTLyUhk2Dnb/fnbw7aeSa3VjABGeZUe6RzEPmfMwkfheWX+pR1
HaHggtij3ezp6sWJrV3zGTde4hQvFrJA/PDpc/575vxEcGQ64/Ku7dJZAFY4hS01
g5TJiDvEO6U1evOx+vINKmWsfHECub4nDfWLXHZs5FH75pmF4av/gdCQvpVg2l1v
M6wr0BWpr8Tx4obgWElFGR34xXnY0d6EJOfaqvj132mS3lXn03i7MDIxyOR/xBRC
NtzD0o9CFAQA+TLDGXsEUgEY+Qz89NBhO0ycdfLEYVwpzsETT8UhcKAMrMrmlQrF
tv/qR2rq4u00EBOUDAP0GPuqFF5n6dbpoBFyl51fZvxWGOIUMyBxbn+n8gTpTjwo
DNbgXZRkDEY5RMBY/+HYUsVYdNOSMG+uY8WDrxWoBYkppUuCNvw2InHAOjwj5BIH
/jjDpNMHu+itWd+fK6FNqVT588s6QXmRFH/isOOA4sf69GPZHTGDv6xLr86S4+Y3
NSR+6wv8KKhsF96aVo+CnYUJkqrnyWn53ejz2rtTV27AE1Y/Yj6ahWRSEG0ZQfir
gkCIwVlduH5U7/vifpyN+602cQdcZvvIb/uGSAiwpzSm+YBKxxs+PRtvbLCyyRlz
auqwd0xFOBFz6bJK0AOTImfvZMrEqbY4h1a7rd3Ie1hryRr37FCF2DIi99tGbDvw
J9Cgc55SXotm4oIoABv1BQL6UPlYXg47Yt2C28CZM6d9t1qdQsdY4tSiZFQ85PxK
RVRc2R9ZYTiygRug2Sr1EvBdgIXLFV/IFxs26RAOphijYD1XqJbNA/fWMhn6diby
EyrtshF7JcKZPajEeScWrHY9iocT5iDqxSgTr4ffw4wXbJn2X5QSugLh8+8jWma7
IOstkl7SmdVP+XfLFdVPjb3PjOXQMC8sgQ66F8Nlq/ay6QReIuHHu+ZNbkWVI+iX
/McSfZ4JRGFvKoAt53/uuGSj4fkK56TKPNIKHXzEkIiDkfRLnBsNvEjvnwltDiLX
WuvdJKyCUFMmxKTizuLLT9VwElZKH0R4uvpJ+U4J9gzWGdLAhsar+XCTJjYscKSP
seQrF0RfVlmmaU5zRxyq51ZSZ3ZuyBx9QRJ1xmZzoalOCh6/iDFSfhVVg4x3alTb
/1j30ouie6xIrJ985z8cu22LDQrodsG4fiZHbY6BpvhDtLI0w35iiuRSROFsJv9c
oyLn42RAgt43RvjnA6dbhfFnaWhOXL5SkDgC3ycSpjbW669k1neWldTB4roqH/Wz
KnkkQFZ+QscLPwlA8ya+wuCe21FWoh8LLj45n5UD9i+D8Wv7wql+XndNpDvJalU2
yjaiAC5QR39oNz4CD1WBA8T2aPm+miCulR4QUvJJ8QbSfIjOiwfWOcIGAmyrlFW6
/mu1bWKJJ9+vJU+xmrXcJL8g0dcWp2AzFhGkX0h9ID0iV3TyyLdx2rnWNyxLZFSA
lR/MzmKNmXbNDIQiEGVlmcpenz/cYfnXi5GVjvtrNMrpN/jS+M3cm1hnQUholwB4
JMNidjCFJcshIyeBrZnb3BbTJbiEq4jMdEZsw3FkJy82tAYz73fxYx9eOycMCiDC
I+HOd8Lc+jMnxFGBFfVIRmfolSbkuC63yKz3ckRIwynyJisjrbpNzQ4fqc6u/+yj
J3FTMXEuSH/3UuY5BkjuWO5e2uKWFpnEpnme4cB4KN8Q3LUcTQC0wrh23aW8IW9P
ptx+G/bmMxGnAkBCiXY9U7GVyjeey4k1wLKG3ptgOlTlOsw/q0K2VJUV2maZhglg
FAH9PG3ZW2fzJA5JadbhWobDjxu/a/gXJ/85ItfsQ6LneFbRv4nOA9JdDrLenJ8N
otFE4RHxEq10B5nR1WB1jWXjp34axvQN0AI5Uh1a0FHogPfK+z12jlUK0HIF72pf
RboHY114yhfb3WvS1s7Ri0ndS6xT2IpauBzaZK7sLyVZ+adJS4RNkCgdbq+GVAyi
tOCV1AP52j5C9Rub503m/jtr8ZpQfi95pPbZEdvpVdyvp0VHjUlC2UoJrDMau/TU
/ZWHab4FyW8iB3cVVdLoJBPsbePLwWnqr/0/xYeV62pG/Rot3gfuqJkLgpKcIfDo
CzVP+u5PeDvYAx8Tgc56T8DGc8NHPbIpblNxRSj4Od2CRcJxtq7FpyMY6wDmNg+d
KOaY5VbNo70GCZXjaO2IvURN0W1nHP9uCK58JeNte9Jc91iZBuY5RpHxNvrJDxub
B60eTanuW/fSadq1RdhFUGJbA3ubQaZrC91SWgtEqW6BojYqAmLN9UA/d6WUkF5T
9AaR1d09EAmDFyzpkAwERrq2RT8OIcIjn6u6/DG65xqvYBlLXC8OXZbBIWJ+arzR
Jpqij14+WM3zfryeYxlJWgyhVSGsQeFhZ1rVhPHV8ShnF1xMqUo3Q0TGLLmSzyAL
jOXgjwksZeCWPw9xgNlsFDobhm7DzL3lUE+dO2WpfE1u51IV3dYavibVtImzIgOc
jgI2H+fo/lreDQq7vHDCq94uRcsgA4eVI3KfEQPgFYPyiQYVdxt3dXXRD04VBt75
CpoTsmD/WHhxu6GwClWkmtcdEJNES0MpMPlHggvsG9ZUauMHoXyxXDgJ586jr0KE
1Xrd8IdYOfZyLfIoOucVSEReWALeytKwY/puzIdIAU6gbVEnT+x6D+brzDrO5sDl
OS31f0Xi/2gHEWZWPBCFcFJgezilpCjtBPN9N0RZnHJZbFL9LPb8RRUxNu0CeHBg
UxrI+OxZTpOKnewwDkU3/Y09KNvnS0nAG1TaMZr2XxCoP0qz1Snpd07yOvbRApzc
11nyFQKj55i2+osUuAlYgIxZSB7e+Jq8BIjIY4UQ5jNHe1n+FCNa+7p+MI0+r9/S
OEFP4+0QHOb/SEuTqJG+OEpNZVB2sQ0GnoBrNa03Ad8xSRNW07FgDu8ebnAwNDCC
r8CnrFYS0VccLMqnKp3KUC9fLAevvQWx+EuvsOUluMf6J4BaH90ZoTSgsLWKf4CT
bvm/xuy5FXzd0ynrFNMPWmTcytwbZEbesFRkheFai0jvpwHcSXQck4r8lVf8qBRG
np3JlEGTpWHQqQm37+apNV2FjBcVnE6t4fTpvnzmOKxYY8r74v4HiiedAmLIrDFB
SFz5lXuZA55iZIqbI3ZN9IojmdOlfcfi8vA3gGKEb6CDcir6IqEnO4X6MdIqBuH+
nM2HYwdOU5O58/Ce/S0ik5UfoOBMrcSZoJpB1ceAdRmvFfB3OrWoHZr1Jc/be8sI
6s5ODMpwog3KYkpxyZ9MrHKVLZhGs/0GfC4ZKG5azBSTrhI9YBqSGOWXF537zr58
xSfirueMJGfxcTipLrAJmNLePTpQTq1M3cA/8OY+BYhLxmMsj+NYQ2eIVMdHubYs
kZekJejYFY3JX8bK8zDVcltCDunzBG1BK0XrnfwscfO58LJ92TP0kJVIP3xW6LMu
d0btZVzGnxHxk8RtpcCNocvVAZkJheYGMtaEirIFwcwWDcpEMzYC76q4TgIAZYB8
MzTTgu7aO4JDB/MdVxtqJxUzWmRjNsgStkdpiAguvAOFH1wr9Zhz4nv2gNCpikEE
1rx8pKHe2k6y+jz/evbt2jx+LgGMFrVZ0uMjsN1/oOcUC3lAeZq2AHg9jjhqiV7j
EjWDclF+psbpqlcfhaeayXhrXoSbV03HWTPxBeZq2gCJd75E7JZVJXWqgAdPHOsl
rr4kk3LNJZzc9ZVINIjHeBqPv3bRsnXbNsKb8zbEgFsaob6jhBttPY+7GgdToEg4
5eIBxPpyNpVqc1Cc+86q7GQcwixh4TDLsZbr2OxXc0YaBn/XCNiCS5bnfbL0qKF9
430edoDKs2kd/qrXAye7Y5MBNUSZDVaepqIY3KOTS3DRb5G4VaT4RCdmvNKctPZo
5QIC5eGCrfvsTalQHQM6oGAx6RUe0OWOowhQcu4KE04aLm6ZMzfNqyNUC9Bv9SE1
GbffVtFLXA/pV/3aEoCAXcfykDlojm8x1KzOq7Ii/TO0LtkhL89nz04LhcgjcmH1
Cyvg683Y/da5oA/HH4wv6cd3CNU9SW9a7ep17x/EmFfyFc4i6qKLzbgNDFj0esqN
lyxGxyBb3RUOcHNG6/pwYSjwfme/OGluZz6jAakVJyd3GVez0iT3Lo5PIS23QlJ6
Uz3NrkmMDRZAW0N4SDkaWqC155ed8UjTlAxzyUo+ccU0irpwgh7Y+EdkFwf5dcvd
S/hp6CHhNVoDvG0Tiu3HVXan58sOYRv+zMMHJd+OZd+PXFkA9oFwtRp10fA8L55q
Oidk4x0bOV5zMNOmxF3Eaj9w9gEkTnksK4MPCsxp01fLDpfNArMp3VBnzXKq+PfA
HqUVT0w9fPwAfddVVjY5xY5gLacir15L3vG5goaOYLny88aeiWe/5MdFE09hQfqw
g7J7YQi5ot539xPg7m47JPJzeMihS5sIfqP6Cn8iO0yYE+TdMnv0e2HC8L8Aoqm0
V7ha67B1EBuXPi+ACLaR0D0lzojT3fn2rui5oFNl5z/QYR9eQlLnsRrZBm1jr7/9
ZPFfloMuGM8fA50OKoy9M8/phVLJ+AgDyuoL0ptFKQDwu+cZZtwxRU43SzydkYbu
tZWgdeJG5oypRpvrCyvkBcbHXczN4v3vJIgKZ+RxprijrpJbodTJDpN9PLN3julm
zFmkXRpm/rFpj0u0nhpfX9nm8zE/PUT1H0YA2Mt6mK8QPDcyG4t20baXW5oVZUZV
dVDNdizFd36q4M9JiR86+BVIy1R1k9A7SL02S7V5cdxz/cZ/I+8DY/GeOokEscYQ
VvrBIcsaQjUFY1dL3LlNtWhdvQk1nDcl4QHKLD+McQPp8O1j0hHNE488iEPTJTJo
1V8i3i/N6DP1ufGPcMCsZ8i5JG7j3EWhHvIxcaM5zMjstuzFWM4J9umgiXWhFQVb
aCquAT5U7i/zeG52zfLIXqpjoZvdB2oTdzqwCHWfKQD/Dbx+8V3ZQWhgCPAIUUt6
ans5JGdNWTwtgW2ytGC2gdVYfK/YLhhW5rZYBD3iTSK+w2XbwmsnF7ippyD8yuES
5ZFnxGcbZrWOL9iY7VpsTlOnnn3j8PIG66SyI4uQzkB7le9f+fyRBbBY7rYYxJA9
afR5NBYzXsZstKJaNN5QfcnREDjIxMOz5nzLeV3ZFnWUIaAZvzL3+g/zLIO3LOg2
fBg8u5gcCC6fYMN++c2Ha8MMqkA7gv52zrSt5ZA4V2V1EnSDgJHhWqWPFpmhYXA/
KTzQ5vCOama7djF5BYop0UbWXZoHWk8ZA6gxTF5om3vB33lnQaIKF9AsBYNMg/H8
WzEofHFovn/toZLMzFbEpVgo/QS2ZFg027gN4DbsZTslMiGTCa0Xwiw2ObldLg4v
mZNplSnQAj6XrRz0mu7h3df0WP77kNYtmDZ7ENXUnq5s3/J9b8Eb9TIeqg83KBGY
EO4120HWTG4II1xmHZxhZ5z/BsnPNg0ghQcbfm0wLSTkoO3hPfdsVaYIGXaB10qf
3SYEVUlhiut3evaPMdDhHTADVsmxCxX/6WB462oW2KVVDWYipydzMNwh55Fw61QH
PjGdaUmtO60LaFdMa1q4KfCoqyFwWDHubY2+QCRJPBdUSjyaMW+UwNFOK64+KZVj
1xiKEza3gkIRkzcQt5pO3yhAv+m3Ma2yMMx85HzV2sFZ/X4DoN1pQGQ8Q/OmnEXI
eorHjTO1am9unUN8v2o37VcD4wFqGYRxf72Ejwc3XAxc9WSiZkCjRAkblk6ExE4+
NhqGTobXLJsrqGR3s51/FlO+6bVOmvBHM8YkNoAeCxwq4z9VmB3fzU895/NriSXN
MQ23BfDLnyy0g4n4IBW1psGilVJ3CZEtQ+a4ZhZX5s52HT5k7EfH53vCl9RpdhJX
yrUbH+n0BeIVdViaeLW8NQSnTRm41uJM9HtGp8FV2QvXnyO34yHHwXKwbCpKjc+r
`protect END_PROTECTED
