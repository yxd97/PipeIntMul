`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wmp7I2y8p1499CLuSZn4sGVcpuLB60Vhtx0mW6HXb1I4MECALAZ8Y9CR68K4DrYL
OjGUNvcIHjtX79sJUtn4j1crrC+Su/MeKHmkY22eBIXSSsjOslLS+wr0GO+hfQm1
UK7Sce97l+7XqX/mZ2hyNBxoaOuk+AZ1b3wFaYLWBLl/oKaqgjc6BuVWelGGnZQi
3aYd/RySPLVCsrmcRn1p0jPKg8B36jwHqja1l6IBpAicZDiXbLSlOVo+1vsI9Hq1
4h7ynnE3JYZ9DSYcrZCE7zAyj+qF8xnNff+VHI2XeKVg0nuFeqYFjXonj9W4Hc4e
bVybLzIigFhVKKcfCAb7IrvCdtXhdAFuQCVz1Rlb+Cg8jeCUfw4Pf5bSkCcgB2CA
ednpGcdmYk1GD1G+E8Y7jkzdYDBSRy+ZT2QGF/gdvJMUVQDto8R/7sz4BJ7BWSCL
Y2T7VlFphudJZl0oEdG+ZEso70IjLiCEoM6Rfrbx7eaVKi2OpMqKnp6AoyurMyYS
PBqEY2+uQGC+nKtlxYCugi00DlbPY5hMn+kdMWVezvHuscSlOiYPkgV19NvioaWG
1J4b4/MknWCRgTxzstoHu+IJbJiEvR6rhgztCr5bHTF2q3mAQNCIcQxbWP3CS+/t
PXlALEkXXyMjyaTqSGNzVQ==
`protect END_PROTECTED
