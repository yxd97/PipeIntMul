`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T1VsFXsax+M49+gn/cv2SWNI6JheLj70nIvfGOHj+2gllOlCPEUEYmOIfkRvw1f2
crUiNXyNz/eLrlNVsRjy6xtjWMrA1vKEKTkSqbVtYVuQAEpMGSYt+0ryRy2yLrRt
JwotHx8ywr+qy81ISq0TwnWJt18sl1GHrxP85v6zteokN4AW8+xzrMsn1X78bvvX
yDfL8Q4ovqIZYGIcM/Y5GefHgy8fSaKfk/NkeNI/y58lrQwE6uj+XV26fhI+MZxD
sHzH7rk0P30S3hBGMlx40T8wLjlqSsw6ac/xc5mBs7Q6VsZ1B4M3aslkeClmUzcz
`protect END_PROTECTED
