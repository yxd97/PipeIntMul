`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Pa+iH4Ygax00+FJ8E8pIF/sfHNh3H65aUt7Y5AUfzGm7pkt1oG1wUOovbN4V7DAS
9vRvqJBKgot35NqxdE+kQ3+1AaVEwKNmOopDv+ctx6+PB2WZTCbNO+NaaVYC1i0l
/VpRL2t+LhJhELO/OdWi/GE2zJQscy97dTrl4jXxHW/NNT31m5VF0aG/ON8de4gq
kJ7G7AY/zfJ7MDndkm+WmWzGZrRojQyCkAo5adpt2ghsVCaFJ3e/C8uybyP3K+d1
F92VDnq4ZmpmBbHn14jD88wcidtajy3HVVSNa1R8F5hJFbhwQKHTMgV0ub88qz8m
8WFUQ4KtiQR/2t8IfEK9hIobujDip0VlH34ZHEp66mwhMm6TMfVkHk00sZSzJlGH
Q1apI4QCfsyrA1qrmZhStWS9Jmm+/+W3EKVlSM88izdsDyilwYB7w68jnBht9Maq
bayBeOJda5lAhKxN0HaGgowNgoGr/7SHCUKrGWZf2fjwcq0JPugUiAVWYlnVzNWR
bvo1569LkezVvAAaO6/t9ZOTXE9uSimDofxczDZvhDJ7oUH3oKbku9iRuFbm9NTx
JBRmqWdDfXMHu+cFjFcbJoHaCU9kvnQ2mBE4K1YOIihlqI2G/huwHfZmH4YGM+S5
Uzpys3uL4wgFci8MMegcoMuQo8GIwSCJfUNJKuPBJm0=
`protect END_PROTECTED
