`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iggjq2Oqn5wh6E6KVLmaNujYYHDZRn0hFVWZgRzmHW9qvR3MC3oOFQerUdeh84NA
mqUNhUNY7An9mJDE4tsGsIdYvIvZDhHnzyY4aopvvkhPLslA5s65p1GHhh2Lbw8b
Xq2wwRpBjzovEzP1Nn0nwqEwyzo8VM1AG2w/rSczfo1NlrSAx75TvH+Lu40+kOdJ
s0wvl8Jwf5+1SNDpuTkmv6d2QdY2iew9+p0lNlnwDWVs0dthdgvq9jGuXZIriWlY
aidypea0mFYtgy3cLw74b2vB3jvHoR1x/ixKCRhXtGm0HTAfbc7rUbMBUAGV8xWZ
IHd17VG1Sqq/V4y3DPmufUhSZcRzF8ZnMAQrrES4FWf7wBH1sC55utFzKgWLEC+P
hAFx3ghiP2JIkltXUn9YhGMzi7u4T/dNmQyb5qcIEMGoXvToXE87bEO7oVwgg14B
7bRLl25Mae0KBoTS9ANRybPfhw3WTG4a9n9c1Xw/zNRnHBITniIRZ6tSSFXy05DF
4Y6S9VfeRCwpwVQb35Dx3OUw+CBo11b8ouQbJwCEqGuDl54pMoaHrOeQ8CzPW7KV
aEtpxXApy2+iPHhVyrDsTWRBRdepN+bUxietsa0rlm93xvxSerwrccHOFKncBhPT
Jy3/7mOs3jizFjlcVzalQppatFHzgWUIK0KlnOGkWh1OmDnleXevztK6A7BPfvhO
UlMs5OIuqIA2o1ialxeB5duQTmsDavdaU6a1/qvz7OCwMH+Ge1kIH3mIt7CURdc4
c8jtsusjARjb4j+wHc9IX8rV2Tt6cCWqNNJcnTo8yg54QLvMcch1/H4in7TPwGSl
2Je5hHQZIBeZf5sbxaRof2kf7gn2Gnfn8ehtd/rPbTEXjXp4B5mPqmS5F7c6oAdo
K3elXC8JxgFvJI5eXV7u0MMSTJ9+9V5iroZt9zKn80NOGIVetAZXCScmAha1P0T1
L4Kqj+9GXdBo9MhpmRzP4B4VIbwxIiNRtjLt158ZBdMYPf/SpsKmxUNKzosodJok
l1llcHCQhFQCWLMf76qbblKYaY9Iu5eyTwCssHxGTi+J+4sU45JXmOSaOB+twgcS
nPzDeaX3KvM9n3C+sB9N7EhPVHgcVY4YrV7yzYEOGaIVX14y9jGbbvDd7FdOgChK
RI5oPhH1vDut/jNZ5egi+mf3wA3vWkpKN3U7v5b738WzIE+h7mcypoGo0g09WeJg
dqqy0S8iPYAwlKpbJZDfqKl9hdOZXZe0VCeuToG7RS1ldOxQ6dp5elUwr51CukwV
`protect END_PROTECTED
