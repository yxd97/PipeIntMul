`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e6LGqlJOr1fJ48rRKqffg3bbSOkO1Sket0I/hSR2l6+M+PazzgJRpHk4JojMSO2y
Wh6GHypB/j3tjI2XM4/d/DNajDeZUmo7WAltahLoP52dM8FQTwC3QonHuZ0njpcW
oWzoOPHRDShlZDdsF7wAGr4X7c1ByPARTTRpnmuoKY5AURnmpjUt5Bq3CzFvFYC7
AQBHf86o5tVXAUJne5dEmKQ2MMKHUFNcAgCWRzos2ILZTSABH+ngVgsI5XLpEAEL
lVoP3vm/vjJltCrGBaqQA9p+h/ZnDaAP9jBN4+CNr5ITkGpG11u4t7onM/2QQHIX
sQMvfsXq0fVQqQyaal0WDm0cP0G9yIqbEvtwaPdZuFzNKFWEkBAFmAapMRNWOoM4
lYsDFRE/ExoqKAexJYT8NQ==
`protect END_PROTECTED
