`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EavW0xzLRgpk1CwZnxBQSC3SGiXwHOyR4IJcJKrIDc2RAekNa2NssaoX/omGBHo+
tH8hElE8RW8y7mx3gaykECGHdRmFq62zMzLONhNvYiw6+/9HVURju+3JktRCeaQ+
DgWjX6Hu6d53JGaSDsVaaaUd8fiut+llmFXH9bHqH+X83REqQ3ngacexA0kXb/h9
dWNnu565/MLmHVaXkcotcLqVAzLkxSgOJl5IxeTSRAS384OqUlVVWdTiwMoEjqPi
0Pri0YI8r15QIPDqteXIoE+hF4q+1NebKyBKFryQKQU4AfYc5bPtiZSdoEVliahj
o6QswPGJf2QF3fmOG0txi/uHu1Ocswbeo09AHtmdAHC7xxNR/IJj8XONQmfYkiTO
nAt6zIaWbkUJYvYYUiPgubN6a9CWQT15PcLuny+qO5CxbIVX/Ebr6pKYcqITIyK+
cL1oUmIx9sN8ii4vIZ2/z6NW7AC3Q5E9d8VHr/ctU6b5ebiYt9RmefU9433aSNL+
`protect END_PROTECTED
