`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PCrQ293NWw2c7nKY6aNzqaYU/62bu78eBt5e56GYWaEAX6irjPL0rT1+LtyJyyt4
lKF0uZsw7b/f3681IVEOD+em6HFxGXT+917vT/ApXW0Q1D3oas9/n3NrTU858tiE
lwJgc6wM2CF6q+5I9Cc23DsRC4YQ8XM1pS4ULqzSNte46FnjRq+sp1WSheaH7r8F
22Ndt9OTmQg5Nqc2T6E0QkAUkAWVFMbdOMZ9Yw4fWM5SK1mF3Q9WPFEICW8xpQ6W
b0c0YW8/HoaAVvqVEUjYOGIpfhpAQ1ROBy++7nIURuFCT4QcOrkKrYeaZZSROApr
Jcoc1MLgSb+S5BUumQyAuPgcDOGppgBqPGTz8O8cDlicpUL0RQH4mq7I3TvseMs8
ksFtYnkz47HpkWIjyb0AL1Mw6Z/YFLA2obgGFkhSvIuywes9HTBzcIhYtVMS34e9
`protect END_PROTECTED
