`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AojPOhnOy6KIe45CCxibfZtH+XSi+Rn/vprHyFjfRuANh94TZP6NEbKlNOq/oaGd
9ropQRi6OoSC2t+kDAkfTa7ZYaNC1uGyWioYwYmICFXqZZ9SrNBKC0E1OtvCcBMI
Jtc2Ctqt2851kIxPNOHdJ8Zn9iakx7YYTq7ttunQbPLLBxcFkwmbrzOFro8rpRFC
h17KkvRKBiQ/wvriFPEkoVbAyfUfif7P5GE1uX7QsztX7w0SNusk4AP/QUjTZkNj
+ShfafTUEub8i4qkIf/uL30gu5UEhiwFdZSlfgDw2eA=
`protect END_PROTECTED
