`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjihPY3tG/WRjwzsohpQ1cEi2xLaGF9Pf03hX7RAznkCNKRzx0EuSZ5j9DRtUnJn
ni4gZ1aUyQZE2buQGhLTzx9N3TsEcwg/Saiyegk46qSJoRbxU9js4CM1rcbfOJNJ
M4i2y9ZZ9+5nVlDagpEBIPW5IkI+j3UzJ1C6wQgcvrMmLgIPYjlxiEny7ZvsilJJ
kVMRDqqgg5rPOvQylZUPisXoDqBFSskozuIB+1/jsNbCGc+i5FvcqpI0OK6kguDT
bdvQL58PNn3NnD4nhs0RvWWvX9Z1gFQm1w0t8eDgxEDPY33T+eX3ns7UvQoGmFX/
JC3cCPxKN+8klyCUWfcv7z3aFgVfL1prgQACH4rKQITrBhKJm5+SL9rH3QhO5uuE
2FOGfixMi8WsAa+hmWS2rhIbUKLAjtypzSSPpfOpNa4=
`protect END_PROTECTED
