`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EaXp7d0XmqwtSqwKmuuQ6q4wtN0UOVFaTa6jaNlWqgbRo/iq2Yk+rMU9gzJ8K9NW
mrBzwRqAjcgLTUeh2GqUcZVq+3Lpmk8sdcb2s1fv3OKX8Xx+Ot0sVbbOlDd4pzK+
p9Y+9jAeQ+61KaTQJ0R8GOLXVeBdKe+lVRN3MUI1uk4IAu+FoZxHZu2jmoAc4If9
M3zwQnM1Ml2KqktadHTOhoyBuIu22bAurRiQnhW1w9tKbSfYG+BqmwRYFMGZ0Ohw
DcSh3E9PaStoAuKiEsf098lhx6xFNWgy38bDxmHh2B8soxfBQPwpi/DTODaAWbJV
`protect END_PROTECTED
