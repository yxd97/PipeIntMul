`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCA0JjZ9AThdVCHWI0YeDrmmQuuI43/0QZRIAFu5M6heJvzXAnxtg1q8uMI2iBpd
lHK8Kpn9kTv+VHgroUuoAvidBXJWIFHPKef4M1/g+CIas3Y/KktmNs5AcMkEfaCd
4PMW2nu3MQFjmaOXVvxW1/uexHw1Aq+4+Ol3fXGB2/pYWrLGfr0xMGZE4VLhzybf
djHQgkOKbTH3bfbSkWk6Anil0IIojHcH/aOQDlX7HrnB1cZsNgFnkYSf7j3TOkAd
DH5Jy25nS3WPAE7iqin2asbMVHkcDh4XZrx1LPNK/IdHKrg/6cmUXyq4cY81MpKg
FEm29Ks2Agt6oRmZt8RJ24a1MtlCThzMXYgSyc2Oc58kee5LxOvmAcYRKmbaQs0X
MS1L781d0nRB1dRSdqACLcS9+oQA40Zjxk4EjbaPN67kQ88cBDAMLyoNeTGtKh89
e6LWsKDUMe6Td/kR/GlqTuoqk1KKs9gkYNnSl5YmAE643OITixvPK5w2aNQzTykx
dpS77am4abZ0EntctbOYtWwNaFeKzKqilUXNR5/wlv4RQFimOc67DuQmZOGeRt8W
RkZKc6yF2XLGBVmvK+JOnNwMzsDDuUFKGam8VdJaftv8mLi6ohyX/9WtvVsbNajt
XvljLIlE4SYMcHkKZn0W+3RLYTlV6OREOKnFNECqEylHYOWRPkWxk6kpwEWXBe1+
nRQcP5AhyeVlKHwJMO+P0bGbyziFkpj1vD3iHfcMd6hYF0rLyARbwWwqEF7+OXe9
DBcCf69urukzX2hYOYFstt6SatrK0I0lKJ4lXeTY+dQpNxqHC8uG8v0ZtaqPlNfS
u7F+e8GbhneEzfi9xKIA711dzLINPnPI4nJPwipUoe4dcAHGsA17QjSQsFu5nz4c
Tf4ml24Kawo3gz8RRAidJkljgu9Smyu2kWnhCAEUG5Ich1J0zi+ZXbSOAxqr5/91
ng5xEOInyiz2RdObkpCCroXZpgsZSgcRToW8YH7UI3AKbUIZD7VUIS/X3DCpH5QL
DLkDofuwlnfdHdbA7xExF9T2Fgd6DVmVs7cSbZYj7GDHYSE9ClZzqCfdp3lBcko0
tyntar6GfkXniN8vfXhyBLzEBV10i2iMDaLHjPbdOtUjkLXOwdyBmGKdO1UBGsEl
QqB/NoZveC4tyQyf1FBtSKJq/IryHLVh4zv47x2nBI4bYM1wACwabLX5fEstZUnw
v0rQShVrNrQB0oecZ0aYchVym9c8rBxFv8nYFOE56cC02rc93fewpeAi4Xhp4O5+
nBe89HRv28Qx1IffmEr+IeZgQRA8fF+0fTqkUsVDmmkLBEjo2Mjkh34PLQIlc3kz
C+J3atUmXHxBQ6Zp4r4f9FVsOF433s8L1KvQ+mXVzbC+x9eQcLkuk+5KyBJs6dXa
kTieS7aA/i6ET1Sf8IicVMQFwEJLWmjnav2xbAbdHlqhlQgY5QhOWvEQZwhutAQJ
`protect END_PROTECTED
