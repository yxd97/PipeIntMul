`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RLQtaZqe2a8GiUhcI/uyTPmjXIrYwkYQ07ArzHBz4tqQkBRY0N+10V6rw0Ltno+d
elFtC2OYkMVt6sKzs5QlNKlsMJK1kJI1vRieuM9d2JxZ/cuJtoNx3d7cMIUT7Zom
Zf/qFRlEi82oPn77qs2szXgeIxMu/kdzDaha5yNdws6HBTnpxByJeMuhyLW/XDpe
ibKBIVEKweFAAknf53nB5IJ8gWhSDoDKCXALJnB6OJy6/ZhKg8QU4UqNEPueDTy7
lVh1qCZQPC8bHJWFuEUNQ7tIVf7NsS9lx/JKw/6d4s0=
`protect END_PROTECTED
