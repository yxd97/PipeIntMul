`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
H39G26CaRhQWKTCWYRdQiIOkDa0a10C8jBfvnPZqmwLPqI9QxfVZD5jwAYrp7qMe
wdsQTYwZbY77jejDZF0N+gJNJ2EOjZwtgjIvEZhICCkYG8nAeRJNXrhxZnqXJiKJ
9bMr3Ep5XhFgcW+lDUeLwgkr/PJPo0JBz7nBIwyMdOKHtwAv/TJoqQeH4BYX9EGz
LXTSdmkpJjTbV4yRS5slj9AY+EGxzKuim5RI5atFlwql0zvUIpt8iMH9huuAWi+N
2mQOVnu6kqC5xObelyUyF5G8mghJ5FtLK4ABYkYRxVA30kHz6CcSgTJq2LucY8id
arvJ5viRsu9ujRamO0VJIOddLw07vu0BEQHK160Vi2wkKosGkQjXhiifHRe97cqk
`protect END_PROTECTED
