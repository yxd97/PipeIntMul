`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XY7o+0O7Cr5WxM0ijwmbW/+8h/DvbEBEjutqQvmdmxEvkt2KrE9WsxbXGW2jhn72
IoUMapG8ckfiumZ1gVrZNiGV5pt6r3cK/wyM5+FxyeCombzlN2JKrprzB/6AxDbI
sSmJ7u0o3uFB+7vGAxiZXMHuF4Ba8VcVDmYlAhkcfV7vgD3nu4CJfObUOWmt7AYq
hg1/rtBS6Q5jrlaXN9z2rHAR5qMIrKdBV0NsRCPkaRNPNizBggve17nH/LQ7U2k6
rADqHA+duCZNIe0EfFIv4dzEqZ6OjmzQj6O/Php/ZRdJU1z/jK1gQcpqPssezgPJ
s24gRdc1/2bfIadsxeyhJFV1ZE5Ff41JNmevtfJfWHaTFN0fZoz972PhGUwU79lf
tCKDaIJnX6UW++hiEL9zojfma4U1WwmDw1agdw0BcUibUGS1k9Jl0hton5lBB7VR
FxColc9HwXSpz1mMP7p0aIDCsYhU1fUNL1ZdQMWpXrwuLSrfPvcGwhTGClXSc/1U
mbvoslVt0Te4sku9TpMYXazpoGTqvWuDSKvwdPs4sW2GcN2JxPvyaPjv6iX4Tzcj
`protect END_PROTECTED
