`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xa9oSL0FOWykuBcMOkK5OGdrdht48FnRX/VLaXpIkdOg50vRZTG3jA+wZjX2PIqT
4HyIXnf7Ne/d/HaxIitQkXpVDAdQbGXI0CGpO+TBwT8Cuje0Vm8XswkL6mFETmud
ijlfa1Dn0B/7ulP/C5aRaqf3Jp92WkriSZ2eVGUuSLuyhHdVfF8PuJzGNcq0FqmH
Z0AkTuiyrkzLg7BRSNV9w6G0p0yMso3a157HTW+Ug1A1nnj03DRgNqhZQcfPB7Hj
sDte4pZMywZygWiN5y3FuFm33Kc1T7+yDJgN0qX383z5OZU3eC0W7TCnaRfMwEsw
Xn602PALToRcG7zOPmxJMZF1Ug2/pfwm4KyhXfGqilM7IReuRC43naPE4tFaEIS7
3tWulySxNP+XFhLq62PDcXVJ/HdfEh2XRw0MHStpmD5kXRSs2iegg0CHp6I8VuqP
iswlxyHazCsmdPaUZX75zghq98haaz/Nhz7J2bUu5nuAW9bAD2oXHpqcxMm14lnq
GetrZ/n0sSaf6doOeu8BjA==
`protect END_PROTECTED
