`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oY4cmuvyfmpluoh+HoO5oOjNtJvwYZCxHiG+QpDkF9UPVi0ldOIwaI4J2uHeccMD
p1PFgrELcCPs+qgD96wl6HwS7n/lQHHdoBRYWwA93UZLMLs3rq66Y6tLHGKPfbI/
RoqmDkEX+akKLWDAja+O2szIGK6bx5LGoQmUYfmIqTh1MhGkReJEm/DLlx7Qh6V7
DDb3G8S9yhz2IizXa16Ts0TWHjuYeA7aB+bDP6ZnBk3rLv0SkRGh2KkScxRhJU/R
VhYyZK/eTRQHOGOpRm5gHOq6yEA0Sd2uvRfD/NDUG+vPuV3LPBuhVo5eT7sMy2ZR
fXZlM0cdk13ciLa2IGXgxTezPYWhit1wp0NwTRF6hR7gP2wArrDasxPFVhORX+cL
V0DSm4V4Q8ih+FPSBeOdrEveHDaiWlj+1nf4urUsvGA=
`protect END_PROTECTED
