`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OLTmoH+mccofJwaz9mDg1JSZ49/8b4dUVrBeGkM0N4z4h0S+EZAH/B4Q8m12NTso
xINlORvUwBBBiv/6fr8qOf8lJXwrRbZAxqprrAsx8sHm7o3EqrXZhdeBtu3hallt
RqgFwPcZNC8o51H4C0t3+XPq+Wm/n8v9JEi/kWM1mieUlT6qtzSOEiNY1higWh64
NLaD+0xqBRVW7kGXtMn/PN6l7nC/63CTXtYpzw/VnT1CT8BCMA23FmYs1MCmxAhZ
t3SMVkyl9FeiOfrNc2T0S+2bt2B2urXMr3ul8v3N8DCNia+FBPo5yYtbTcAhXlXT
x9NT+z/LjqaOSpScPnO3y+OybWhvu1C1JmjRJOQMhRXvKONXEE/k13sglq9xS7F1
7NQaL6bnOiNJdgkqbvBYL/A2EQe6/ChopO7ipE5tqVxcjgu4aNWlx4LwF7rqM8Od
`protect END_PROTECTED
