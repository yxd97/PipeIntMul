`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
czTBj9SX6TFRwHoBAj+L+tP/HWZko8vNIrV5Gxr8U8IMNtsD4WosWwq2uVLtPxJr
RVKe9OxHw+Fy0OJWBCcnwJueF+xs2s5HOyXJCHAQsk0c3HY0YI5/joT5ocgMaSec
iok/cjuHPYo3yojKUlrozQaf2xVQywtOv73aJhvA3toQxhClS5OZfU54GWPfHc4h
v8TYLyaHne85OsyXZRza1GQwvhIjvKXGu6XDxm2przcZ2jEo5q1eUa7vXi4ZNyZb
GwF3jZ1YO8BXRkc+ZoKOzzJItDxoipBaV771U54HxJWMQq5XEiOsLupPDQRRabHm
VRJBbqwKdIbNwi3NfDvCji0aRhyf7l0D8/aX+4lk3SKbgvNrqpKod2Gj36/EVzKM
DIE3ArvZv71JvO5qwQjnRc7m9tuiauuszWTg4OYRFqT5Tg/HaeGkN5X+iIEugZRq
3Kyr3E4Ho+HQWifmnKyc2v+zCZoZUYHr+UgigJyjCDiNFq+iF8llAaS2T48/aTnm
KXmIhOYrFFV3IYPE4jzaCFs2HROqVX4iRs9b9LGOPUZT1BTp3Wkk9ANWPRmmjmoN
N9sehFPy1/dRTBkGPJny34W6QXpLZLtbrv5a1blyOON9ohVjkJbTQWZbc0KBdzXN
bFGiNfdfgkhN4+rPXig0iktLHQTOtJils8h88KVGRWytEBXxpxjnL198lLigqxLQ
4YEJrPhsorQ/obsDhKxiStSDZPWVrL/mKsY3md4fZKteq846a2IerYGfgNNeISEq
XmWg2GUyPx4ytmH+1AgHxdLnaHADsTjlHMHER0n0D+iSXngH1kgd+hq28M1vHPoN
iTyRdPhFO5Vg+gWY5fwv76ew1MZ4wcz4xONDGHPApEFgzlSMwOlR7U7p7nkC+VZt
r1+CnMdBGOevK2tkUS4NTBsDnMm6ya2uc8NdmwerkPxBbgjzKe5VQRHnPc8Lhxiz
8udeQQJ7AMM47sFNiRsyv/8B91eDWfucVvZUYSVzcIqez2HwotY81+/QAj1F0nKr
/J6a4At3QyvqY6wFJWmm39WKHluH5ERFcAqw5hRBlKvFwKpgi1w8308QRhR9MdiU
y/Bu0gq3z+x1+wM/mCN2DlwGGDGqvRhfD2kwP6FOghReiBUlMGAYSDbQ6fF/jRfC
m+QqtUvnGagBjSPcFqSXQLINx4dsm7IRTTvPevuS8WHmno9KzyRMEX7wv+phLmnT
T4Aeb49XaGmJIM3IBE3f4JJ6wRTZ1z/fXuag5FP3ItmkboA+PXhDr72+N/plAvwP
ygUqXAUzyGbKSKAV8A11fPZZlAg0avNjhXyi9Xug3qtoCtdhi5rI8Ke2kPhUOYYE
azWfZH3rnNeKkS9gioxA64/z4l+r8ZZB8LzEXlYpYgr0l+S+Xg0KMTfLY81M+XQ5
MOBdBoTAFgTjv+M4XajD9Hxm0zvKF7zpKDR6Rdo0z2FFC20KZIDlgSzwpAlWSCWc
QUUQBXjNgb3iTJsSQ7A3OgRfTeFUg9hDV1fxvDp0/oFYqLG31PNayGzHIBx5WWbp
TafQWXUto3KO/szuzHGFieXfJq5x+RoVpJE7fyq9iWFiMsOctZkvn+fT/GelIkfX
AnlaLCOETKQH2ITN5JWgJGbgovquPfcPvZvvdCx94KGtQTW2Ek53IpJyt/+mOpGI
579ZjtG1rEVnMphtMSq2KL22Bec6GrHIvPRMu6Vkw/iQGCZsPBveDkzw02/t4naS
9JemaYHrmlirv1BDfPx6qGScAuhz108rjR9jmk75Mfo/Acp4svla761QcsPYrjUt
wegCMOWYgIAVBz6KtB4H10/ULxGWb+Jfg9RtxwSj+oC1qagXR9DCviJM8nq7fp8I
wPqUVqp4HX0aFJzdQFuZamhKsQf0MlSk1UDNFLjVdywozHQeagZN/tMaqJc/leKQ
mcuO+txN+UY1dShC+ROGAfaGM+qRlYBwEKrn6SfwWLVD+c1cnhH6f/X/7/RmG0F5
lHp80oFGNDcDmjgo1MTtWad59FReQhd+rGAaHBBHtOV0g5qCnFMZzE9gf69TTgvy
tIva9btf2tgX4TKJRglLxHYPY0M6yLX31zfr1koky1dbON3IbhUJHWFQrPqbSAxJ
yAL5pPQvdFaq+yKNROA2l68BvsmuQKFA4ftxPO1eRHdCfHWeNaa4II9/LmyBHfj9
BH6yGmqCwn0UifQCwiMtOYaF/uH3Ab3OfMU/ryTsDd8Vd/GfN3JK4tJi7VUfXf3I
xOUE6J5W2PZUNuHlzeac+206u8OymhKhDNLH7qTkCVgd/vnGhBIAk7X/XR7Jfm0a
PT9XLxvkC1+vGOX4+qo2wex8lzKGb3UgznJVYv+6JZhg/unHBR8vYwyjxyHbzNUv
Zi6XJJeDIU7caN4nFSV8CCna+d1MXZZpEvDheCN/XgMyoRJNpN14dqYi6FvM66Qd
beykWHqw3Q+gr21zbPYRt7GSbm5PEex+zDjb4Z2NjqEBsieOLNSohqrrCt3PthUN
5rn30awr484yYVMhBS+frT6nBvoxhI2M6eppbBDMzTRYXQuPoYHH//9qsX7Ytc3l
`protect END_PROTECTED
