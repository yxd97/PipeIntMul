`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EhxIGGUXks1+lpw82NzLOgiOhls5xdBb5pM80+jQjQzMQ++vSmIvn4P7a3ukmIlk
TBkGL0dKQ8k43CyOCYseQ/MMB7fO9XkJR7FQQKjqJW7p5ya6opZaItqP3TJ7eKk3
85XuBv+1PHHWWgEHUtJodDRmIAB56xKq+xeCFcthmvMmf4vbYaqhkj+TMTILyIFr
GjC0Fxk0FjfcrGtWvLe/ZCB5nw5szZLQ3JjdbLIK+U9uVoWKLDpcyah7Mj84wKmq
ZNDXLlqBOS0XWsWkiFbiuRKNSqTXIBQvOA7w2C52UcTH7OrUg8SmN5maQbqe9PiQ
a9uorsyUb946RNpKZXAgPu2YTbB5FOYmdmakj8rL3oM=
`protect END_PROTECTED
