`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k76B3e+10Q39fsLNXJEZbeOvqlyWS/Y9Du9cTeL+LmBaTvh4Rqn1DyetgAdegBX5
sFnltrx8xu6c6nGt3SpCFieZVnbZuyJkbg9ZM9RGrtN9bwpRbXk7asojr7Ulh0tT
IiDaLd2UbNr6vnCaeDgS3PSukCGv6pbIq5kDptWNEysGL7psbJi1TpZlryRZltQf
nojqteGWOnB6gzJ6GL/lGWE4scSVNndq76CbqtO898DeHfGLC7xdf329GazVXHX+
ssi9Z6SngWbRIV+y1av9tyFvKyXP1vjiy1VLPnUsTRVF2DHuBHD8JDvreEkjPU2C
325N1yH+LpOEjlAimb5tbLVVDXuqKRM/iqatBsyQAoRg0nSHsOZB+AxqiMwimx+R
x9eF8VvJ97YHKDOsXDC1vrHM/I1loumg5C7BUuq76CImBu0wv1TTVvILdBqOUVE1
rdQNVtue8OibVvzicvUoR89RS8R5cMPp7MTEkIj0tdQ2Tib4Wls4QSdeC+33oviw
IK9zt2zdzv4glKs9+PrAanrJlgpAhMWG1Q0u6SDpMacjWj5q5Ot3tTwMykckfUKc
yQ75v3yBS2rMxZl1HFrS2NS2KuvQp2JoYjtYZuKPlzV6l7yOknMRLq+OgNyyQ7Hu
OxicTwrTMDFKPMiNGa1Grr9oqvV4cX8PaGPUnwpd6YuLoera+T+dpPrE5sfWyS+f
oO+2rqrbqjf0pAbxJI0oI/VCagyi6N9ousguQGSoF6VwBYL1L1VAOsHj6/jHybph
faBzQ1ZmvFhPkxBiZd/9LnsSoEk44TRbzbe6snXT8x726CtJq3zaiIs3WPf3jhHU
Lmy7vlLchUTgt1tqg0WfKAG70vNaQz4qmtR+Mt1CnQhvkfMeI1AS69tjY9Wwlvtc
ZMEeS0IaN4DHVIQTnTwV1L1AvFA1a3SSsYjZEAvByyq1ooPKCApjfAXC4VY+V2+K
VJC55u/3nTaOKT/urcbRiFeFDlyI1RCuXL7rZ8OwZced+hub1I5RWItORX3egH7d
INrHkwezVJpgcKtkD4PMQ4xDeX5SNtuK5pgkgCDQ7fU1lAy0G8x3TGWeSxfICTz1
`protect END_PROTECTED
