`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
R6Dod+cQny55uoENO9yS2gc83bZnqS87vN2TauldJbj4sVZMmMX7GWJSytBfXCAa
M0ecIU0SnNMSt71El8d7rHh7SN4Fkh7vkdBeqllfUPEQSMD5tVhSYGoJq425KeId
lEXl9M+svDd22aObEsouVKcdUonKwahZXHK0+qC3J1DtsaSwcuy4MYkeaPvLfJbW
xI6xcwe1r3xXwdp5EqSFLl+yT1OA57KSQ5MiJeDalNVp9Qo4lBAE/4Se6XC61ytO
wxMOcp0S5UOLvljp8Dggl7Czs5mnPUWTTwo9lCKdj0RkPGKgk9A1oetBNLbDeIqc
czL2jrEQU1v3kQaZtUh/owAEuGJreuDbfln6KJpdSsUoG1bH4KRVgEtzlSW2hQyX
XO1IOMfh2TYaxi4wRicp/w==
`protect END_PROTECTED
