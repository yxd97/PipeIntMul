`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OqnMdXGSO+BN8WClc3xw8tYSd0zISlRPynrQn2bjDlFv//jk/SsTDGWUxVG973ch
19sG4Nwa/J97bBgyUhLufW70aBEiJ5HNSdoetDaZSzpba0KbIj3IanmHrjiRpAsj
2k2czADKgm6wJqmTO2I0l0H7urnlZleGxtF4rcU3nVoVQiI8JGhZUleYMG9M7/tB
25HmSTqicoYtmTEwu+HVufCCQXt1FFnM3wA4te2pIkwkycd9yk10fgflMjt/Mbiq
I0LjlalDbTEMNXuS8PtGYAPb627hGhpwoWTekKfxkNNNHWKo7Wpt41nhvVKNzz93
mB1p8EA9x3GrqmmVAA+XQIXzq0GWkUX8jqH3hpdMGkG3DEms45AGE5iByvEQL+jX
aVSbfhRociiepKqwBNN6gn4UoS531WVxACe8F/vwVqYJeqUsZ8FI/hXLPEmMqgaN
pPJo9VVsQRkx6jr57SdqvPHBa/FpPwJAJ62f1HU9/Nhkp2ax7ovq1263iBVYYqhX
XJ7BDAfKqnYdBYbgX48PRxhZh6WLlqVqHWaPHfaKKLP60vO9ApLlgNeWBhxBXW93
C4j2nZza9/gIdcKPFMi5MdhOi06cH1u9Nkfif/1PdmHkTxFOTXZkQT7MxE2yabGo
nckS6mvQOQ2ZBnpQfpiJaYX0Y3INp2txPNAYa5evSg39ET5oTEwpYakrfBgWZrE9
G1Cmr0AowMQOwtbjrzcjTud4/y/3RFsJdWdx6sgxLRLPrPryyl8/fJDvtzd/3afR
JxnPPyXREN6iO8IHxXs5Zp77K0U2EVX8ryWJjXJr02U7G72nDeEzQi0ItcQGT+7s
r17QKlXaXrqZjGs0WcduZ9391V7DYcezwTA9JKm9fkC66l503hp+Mb3wYLPOe1Uc
0u2LaLP2lUUcmU/sQkrWhG0U931jHqsWewXsywGUKlDQBxN/P0L7olDNuctPY02G
1B3Mq8g2kb14GANkbU7etK22D6fHaerlctXSDV2hDW0jlX6x68aEG5vBcAhiR+vX
UBm+LkPDZSDCKvVqiZydWvkjwC3ks8xY2HHWWtbu3Cz08toiPkJXpMjU8kIhPGt2
`protect END_PROTECTED
