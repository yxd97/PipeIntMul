`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zRGOxwXddNSDcUz+EYsN/6dBbfpIC4r9cpAUvAa5YR8MGBXh0obw9N+OzJdgMAVm
xa72VAAW2TZM1vv8CndDuc81YYBWDqI0m2MEjRPf6iCIwELXNJA1lIejcgA6HTKv
nz1nBalvgLzBO34NgcdTyAfJ5bX8nob26VYdrwHxWgbOH4uVDGHOQdX/oC3ZFuf5
JUP9sXLVEBYQcbwMP9gSV6VVYPSC4J7ggpA4QXj7LTqGC/1e+byuvElnRVWj8L2F
fIRuMcCBVoK0S5TZWupg0buBdL6/Zw4cNx4VN8yp+aWyYcfLo5qcYxsoNvPJrKnC
zy9hhVhCBCRygWazdF7fOhq7dpihHZOoP7mrY0MPn4ISH5jdcUicrITiE0fdgJ6w
dKYEjre7hfuPLzSAJN2goH9kZnHx6zaarBH9SJmxbf8uXn5g6r7P8m2sOgzaU3dO
44xEYhiQZD8MSL9EaofTWKAvtwzcfFpZW8k0r+qyfNjoewqR3E16PWSXmiKaJeKQ
mGYF+8ygl+fC4SOw72j2M8BburttRdfwvw/vlWSJ+UEPAULNijllhGq5ZL9mxWWs
jp6IM4zSFb7oGPnxT4N5iw==
`protect END_PROTECTED
