`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OIsdfor9HN0f7Adu3z4vqS3rMKIhe9+W9WbHUqdYeVYOc2SJ9zJcJZ7gx065yfYz
yU0Cj8nOUAXgCIyUM5lDR5dY1TsqeCjxJZDEhRNm5IQG2axxi016N4ezbE5KbZK8
GgCRPNqB9FyZUUjSyC/+8/9YC94ISFLhxmcv+RDppitfAb9dnj1IU4dopk5PlYgO
3gHMwrp2tjf2eqocbkKRA6gjWmo1CFmG+1HdI+aeCtJSV4ANBhTEV81Zw0DPLQfC
wR9tBMz5tnu9LIuzXX9/tXn/A8voauaKLs23z+f+UgY=
`protect END_PROTECTED
