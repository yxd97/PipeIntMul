`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6EQtmeGFJEhgUxTwfIOPMZsJkBZ5Hd+S2kt2vPchtgNkupcL56XlB/CdnGc3s06z
sJdQCK4ZprRaBX2pOZVBzISuOtRUT9eprqsfzTlKNqiXr39UPKiW4r1Eu04iQV6w
KycV3i1Qx2uZ25cIgaDU/KkcNN4dHqNzK+v5RSTNU/txYx5bGKxHhC8gpgTlIBP0
ejYrUaLdKrIbcMeVw+Bwbf6y33AYgITkSa/teXnXVSWTr9ZCB2bCa2v+HI9/d9gj
xIFXsuuJyoQm1A/CZELZxDUv1fBR4sNkl+kXlGQFR2h1grz1Ws5cHOJUBgOWzrXQ
dbop5TLQQ9MWRx0ankMJ9fkRio1vYwrPvo1vj+V90lrOrR930GtSMBiXmIqm6FW/
JsBd1FPINCQX4BaVm3vKzj/+rZPX8nBzu8RpyktyOTi2kUsAAdPT+EbbOM5nBYvW
1lqz78IJXr2t7MLFXLogKXvzM9yeP+Tw8zJTVv6ML94KhlDLj9PFvGL2zuSu+fvS
YtXOUhlzUc+nyJWlrjuTNA==
`protect END_PROTECTED
