`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rojR0Zrrr2Yv1CG2nXBI5Z350bkNkQ5TAX8sezrwHfQFHmgD6CgXCjAe5fPlrdrc
s8VvGXOiagAVf2fV9lFXuew2gmr8tnvd34pdB1JHqbPQyoMyErIn0fFSZ4+M++HD
AB63F56zqfAkCXA2i5WSRILWLRXEWhjwj0CUXakX7rLTXkh5wNB26llqir8E1bqu
sHigWrFNv1l7qcDqnegJ0ghdMc2AHxqaOWt+YXljXOdi4qiaU4oIR6HwOPMFux5R
VmSQP8J/wOu+rF51M2VcaZSLS672B18UE0EYEib9iMAgfZJzSpkq8lcZX2Noruo0
2b4cdAUOG/BKfwFhcNVrgI2J+s1+dw5eC49g5F6dPFGrJbaQ+MRL1t7KO2DeiLtl
fe/cs4qMTnmf6dwkCOx+uG5m+AilYP2URHYzOFH/X6ZmqMK0HnDtCqNu5RBJk/F3
BFC5c41hQPl9U4C4WB3FexRuAKPR35IRfwqtJP/ygxD+l5JLGCa67AzKwSsyvoPB
kz4yMi+lfSdDsOuBOnufv5q2IgLLIm98V/OLAYybLjc67sNSIv/220uNTBIgy14w
g0OAEpo5/0Uhsi8QR5nsUGV2+dpG1hn6DaRjLbNtPX9OhhRgKu+67rFGK+qpVWUB
rsBF3XC4lzU20ak8oJPatd+i97I7sTgOpOBUENq4STmmwwE1y9HsytQX4XGqY7rh
f3uxcUR4M6T8TpYTAdY8r0BebzVH4Ysfhg/zteVq1DRalKhvLRp6HoG/cH6Xr6sy
Si+hOa33/a52tFmpZ0Kir4iMTntJHFvTu8YcHgYuyzvRUYQkDOFW9oK34dMIjbBL
sUSInCzBdPC18kA4NGmv+XY1NOTkUnwsGkj8I8+g4ELyOy2VgGchkWd5q9VuMVZw
H8CY8qQhhW/2Oe3aL206sbX39KNTVELVvotPwrlAX0uVCnlokh3Cqst2TW+cnxFr
zaQCpFSATa3kihAvf161GxJoW3ApW8jaktSooXPvQh2nqh6WwU5NGfKkIH4BHg2U
cLhNMe98mrnjz/K5kXQ3KkjBcyF8MILmSCRXFrowNTGn0mEmxbcenu2durAzsEei
SlNLlWp7YIe2I4kgzmRupGwyvNGN+KMkyxKlgeIySdhuqiBYtNhMyLkITNUib+yF
wExJBK6Q9u3fitWnjQj7Vk5xW5QiDThAEQWrUz7IiKh4Pl9JgYfH6yFWhNVMtgpG
FWaAQizg46xaHNujNKEKRt4ASa49Pq+CLTLwKXb53CVwUmnvakbWpuZUdwQw8Gz0
ITmYeHa56sEYMP5IzCfdH4hkvWsOSuN9EBHIm0a3bR4ZI74LLXIV6ylmhVkjnurS
C1SDO8gFkECyNiQ2VCVfu4MOBQlb6NUDJqXSvm/F//rr0grS8MG9kD1vk9BHbFRK
7ChBUxORJObA2/JLL61ShcJ0R7RZGafRoioxFUBBr0txlWsPpAXf9MQ2Yut7sGHw
Wm1anYGgcvi+BkW4zrqI0n3wqGsmP1ZX9zScFnVhQv6FQxxmhY/4QSG6TGx/rHAc
uqjGB+bqD2M/0CspjNr3RVUfvZZHRrNEV+dyvSxBXJbQy5JJDzA1SDU8MHdqONxh
HGKwHtp2EjGcDZZgOZj4apIYcNiKtCS3vCfrosbvevWAtR6wr6EpyWz8UBJia9R3
atwh7H44F2bKY6VEpWxy1aSi58tXtjx9o1YNIROLj2Oess1uzXnA95fxS+128cI8
pMoBdLjBIq8oP2n4Yh59JcO0i31iKymw5ayYcQz4u2Q3owMq/8/56fviUrjezIC6
KnC9ct5i7UtOwLehZ5pjLIwTYgi1L4XikEsWbnPo4FaAC8RuqY+aihTkYdmpzWJO
jOxminnE6NJDpfVE7FPw8DVMlxYBPpE2eHMjrulo03rxceK6XDMTCeKhOGvagg0e
AxRqGGmFCNXkovP9lvTC/Pru/SFzmmTd4QfjmPPLFOmx74zgiiqhacVMrne8az3D
erL6wmbBp0eZuCHW4cIyqEczEPcRy8usA7C4PXYbMB40hCsCiEyNGSKF38rnPE4e
+WOCJeKb/5rIa4Cypzw8I8Q07i54Kq8gVPvoy5Egicc4FDkXauE2NAaouwA1+tkS
H1imkEPcEQ+ZR2pN+3hxsfS3LRiJUQjL71qYHXSlYy1UA7fRjbDHE2m6IeQCbIqj
KpMvfEywcWU7m5X+l6pjYJJESZpzHfMfUsC7iS9Blc8vQbT6weRVFvZ2kBjSYypw
LW7uA/452TvN+rP9Ti0Gm1mFWNbPVZ9pdlqrP/00DyVmkCZgE/Gethtzq1Hq463/
VPZiMibAKkoB52RQxC6Ph4TeHN4cZ14ujTRWpbeCmvSHW4ptE6ILvJkgnBpBa6w7
TGlhzr0Se8tN56a2EhQS0SwADZSPiFQYVeJu+iG8uP0Pgr2AmtzT2ZHFymJhfC9F
DTr6HzPuPJxDAzvwdX1SOH8nZajf8lLLrvoe/wUm8uWp/SlJJLowV5ZzW60GbeP+
GPO/xTulmUACsr9+CD2ciyc9/Xu5UDwLF3cktNutvN8iAHq2oVyjk6S364mNXHgn
r9G+TwBFlG2ERfDv5lxNUOm8EGB0m8Ss+HOZQc2Gg4y3mUGctgeh/unicOOv7zK4
YI0fT0d51mPs2V3pxlWZQOZ9//EKOHRlcKPtoN8M5juNRK4h/l0LruKR/9JUcIoV
eEWvG0R0mEMz8cULGylsfR1n7kvLxO2ukYMP8pM23Ppk3g7yQo6WjGx4LSo37mKc
97+xACz6+j29GI/qVIIGYd1Sv5kuOxmFSfRXInfNC9cNmpJx/HUXnMaZoWqEruOF
Npk38V3ZZRIstRQBOfW2dA6m/uFORD3HDLVoL25LSzoY+/HApeoklgNfHH1V08aI
DMoG5ujSgShSH9hxdg8wu3JDM+ovd9SUHyXbytYVzee7mJIanEglQoeXmMIpEy7h
s9hSyaa//HOQpZjISu+Ekd0fD3zoVEHbHTnwUebPZSSP0PKyzx2oc42WSkM11RC8
1KSGYfnlGctFcRk82mAMqIIrO1Cmw0WVsP1mq72LVdKy2EYF5YefBfszouxMbglh
FGjb6Su/1q9VeyLyE/QsX5iRpgsQ8ckz/aFZRp082DEKVEARpiiw5/I9aQGhZaK9
qeND/HZugLEMX78kE5jdMUqHceGYo+BJrndmS9bcWDGD8xYHpTTkm5VGiRMqC0YO
q1eSDnJ2rERO62ZqDbCKZR1s5AgjYUcPvJTGGr3uUJLAt7XcWAEBGXbyh7YywtPh
JNoVqKKdVfPu01NTT5KWNmFi+3f/X+L12Vj5XA3zP8xWUUn9Mq+7dzEXinL6vmgS
Kg9TD/Ad6+QgwtKl82rpOSkEFliUWY0lJW/rC5olxT95ihdmdcmKRTt9+SY9XmD7
dQU82gdO7fZERNGXcceQwUFF4bSa8cEaOM9e5HK/gxLuA3kYHhEiaLddPbAyZEGo
DUTGdZ2JPgdJML/9UZ+9L4ypV9y95z2zvddQEQS2d0VRpNE5mGED7Iqjiq50/wL5
wGX5Re3KyPAyQrIBOf/b9+rZCm+suik+DftJeivgmAcW+FTVHMzFksuUF5ga0cEA
g6L2pzT0BqwEgubMEImNvVD24MpoVZU8viFY4ZIu/ydX+N8PajkvNF2Yn2jGlndo
EiiPRWRe+fWcjtpFhbCRNOps/4QkftKCNdtjJtgLiyossHFgNrsKflxdBvR6IMtl
tAYMaVHBDUI/MM+/ImGM9wbuC06VqlAJMf1moRbyeY24yt1r7z/6YdXfXg6I9UN0
bxtMwop7M0dORfZNwhuRbtF06Nd9oS1fiKejNIZxnoJyw4Sl/sYinO6jpxs6NjId
T2YM/EdANCyMwBJZLV5Qkp1crzQrubo7wYuPzxvTBkZ8WzpwkwEEVrocTPb4vXTl
nokFEz9nX/0AcpLVlnhfOdi+P47wqYMXGN0AgJHFOUk8FGkXSwPkNOx0DWHgzBSb
TeCe8zKmIaDCWzAhHwX53VnxTFfYJHY6HmhUMObVnGuquoHQa6GvftMkgssYs+y/
j313KaZdofeZMlHmRYDo7wabbz7E8uPjAwrrhFHvOuxLnXodXCLIMKu14G5u2rr7
9TFfgdWrsFf2wyR7PxfKwS/Yg/pyey/Hw6r/bfqrEBZM+Mwuc0pcW5gQ+Yq3P2TY
u2SH0SWTHCVHPrPIs+3COKaG08nvWxYWxnRGvScpTfwDL2zB+DSwJzk899oogUhN
BQMUTAYiwZUVTQISWJB6UWKwm7Ow0C/ZwMayKkvaWQX5mndaOpcPECpnyH7u6bkp
E5tyAtmwwfHTGBUbcuW0DcrLl+pR2gkFBH7HraZCmWqLhrFG+T1rA8olVrgXRYMX
riVHZ7woJCmloKBSWc3OAOy4NTCgrjaKb9rJHB/KCWluxC7tH6JxQRJLFyFujuDr
5PHxuCZxszooC+S62lqI9/0kI2klrTZkPSUcP93flGtkB3XE848sSDwYs7F5mF/B
7M4kVOWDUzbUlyBw4oeTmPrOSnTY/Hfzp7JAIe/4RhgoWi64p28sjehvvqKJ7fOb
ABk/yo2BOfNwbl+69rnmXudqzsqznC7d2Q9BA9B8tf1u4BtAVwYbPt01PmbG/ouL
zF3qX/t/NxSt3m+NaRdaScj7h2dKNB3ObsRTELEaGWzLHEkTmvyWJgR4AgpmgeF7
7QJOujVMx4H1Z7oQceewWaOLXhOayT6S9qSlydtFal1KUwMky5hXf1OxVrPr+wKC
fUzRIQb4kUO//D+LP+TOsot7/OrfYC4A0ma1ERwdb7P3nffX5JyLylXEwBwWmaNm
AqpROIpOPFClQOLSAJI0Nbbv27JTiYh6q1OlN/jGpAg2P/pvdWl1iZQDDvUEYdFS
K6ht7yg7pt7BffwlN4nluzA18OFsGhb5CtUQDsE7N4Sf6MnxRe+U68v3TDRrjDdN
qXAOIuHZZbOm0D42bvnh+hvFBjpOmcs95sRryDege+z2B4L8HBpH8IVyjP+zlIMS
Rzsd1Ryxo1isBkI4pxjqDuC8+/xHRl8VuGH/7FgteHahB/DR9tchBazvicBih6wm
u+b2ssDDxEIUX9NboY3n0NO3/5gqCq5nPTmgPnoV6Py6MiHDzjxelPi+Q5P9s8Z2
fTtlj7jAIODLvYzFGQqrFvFrOZdqPZVnNymxAi8UfnCrhfGRmhSDW22sP0kwZRtA
0CXHfdwEQPyhg1tOMC1qJcZ3OmbNsCqHPz/KhyDUc0WVGIDCTpP9kYtQc/2s/XOn
BWnEPfEFVeSnt1tC4gFwjFZTemD+MIFuQjBg+Fj69oYH65sNj7jXVc1uXW59Ds4a
3NDU9uXP0OHO1LH67i5D6DFBB3oCeUhpnT2PfRn1BmkjqbjJzm/c6nXFXSxR1JS5
z4o2W4NPRT96FqeDlnAMWuzhZn4R6RYRXZT/d3sk3sZPtNgHAHemMBAueTqTCvju
Ruswm27qzUxBLxPvT9zcF4Q8SVcHa3hf4AHlDNxJ2TEitS4Ny+pZR4BOj2KYk2xq
YODc9VpGfOLr4q+BsF88O5wpwGQYScQ8Js3XOeV6CMu+shSdAC3jcTxVjNAfPrjn
CdMMB62u07ESeyAMT/6rSBxDekSQVDjwbKzhtpzCXtnfSlLctqIriMpe5DBHBvMt
dV1XM/OaN0JSORm+9EbBz0JIbLlq92Te9WrYXMS+Z80gOJ3Gkir8JFqVf+0AcjCn
A1DI0ylS0dtH8JunQiJrX829pjJ0lD78FMLyLp+ZiBXzhWoSHVZdFierMLXdOjNv
Pascjfyc9Av4as22U0yU2aRnFLWSR4n6oT8rV5Kvr8ULcVV+cKCI+k29gLgoMkWb
YuXgkqRGKuQm+QKiQQrR2WOTTQogmTHmex+xjGUarU9BW1+io2sstAIgUk7ElXhi
opt/BbeHFYTUl2b+dpWGKMPteWHs0rkJrChtk5Cq0S1ZFL3ReHb9tjPSg+FK+RW+
o7pU94qy4m+jpVrWIdhPRyvhfSGFYOrFSq5/tz5si6TM4aR6e5tZLFkRMtiikhyK
uMVeclt/emiCa3RJ+f7LeI5HeoHvXTPY9oWGY+MnionEav1xSJd4S6iBCsMoVg8N
XVmi0iWp5qFeFyBDOoBlYGVkEU4UwzsWQq0CZcJhS5hxwpGW+J+2IAdgk7CiYD9U
1nTbQleHGWpwvE9mbn8Y4FpnW8CmtKvv2+8QbuyWuBd/15nEPWWT7JvJ73+Su0dv
UrVCNlLnpwl6RHGtcYnJFdOfyMppX7+R8XvGAWgzmxxP3q6OLyJ5xq9Vj9oQTTjk
YqSd/HqWAEVnynr1ouhyEFDOVRhzG/FxTilLI7U9d5DokdedCkHuEWm2t7EVHY8a
rr2FyEuiwdvWZplHhI3pz/EOz1637NBmieKYNpxA3lGW9d75wum6rIpGrKQQoC0v
ROqcGMjj1ecKqHQV3FG/2gj7P9Cn/vsyaxcGt4xRdphFyJFDx3Ju16Ww+KoreEJb
W5T+zzcl4VEGc+67qeQ0cJ8iW7AiPwSZ0aIhRHAPsuLgXyAoncsOOTfS/OUe2bgG
Um3S7VHvRszelb/HAhyEGAdGKcm7azbsfnqVP2ih8+uoHf/APh5pScjxCrnFfMNF
1Ar8rJayzi7cfdES4LAaz7N66/QyHvF0imnFXZmktaUf80safdU3ZOz24TK7CUKI
kZaI0rk15yMuVEt2AVv6akuqFhyXbtXEXMqXO/59ROakcm+vNfy5tqe41gxXS0oW
9p5O2T6AWzVUvrztpeyidREFxNAOZCH5F7au+biIAilZFCqPm2L2rCiWDZT9JxEV
qE6FPkfAaXFD+6Oz6o6yW6nhH5At3PxzrOmFmkGa5kbIENvMvlNZlnVfLtQYj08w
/wLqZxOeWbuuKMLFwwClFsbz3Ey0TGVZR7CTv9OzBA4/5i1aJhDNVUegRH7kGViw
5ezUfMgnhwKzn2NDJiSlR6YYnIkBvksOQE0H5S64vcUEuw4dC8hoI7C+Ksg/nKCp
XjEBGMzVRVpD9yEKF2Ka5z3zUeyhenFsYZlOgAPgBLxmKIlBy8Ye8nsd4Xt3U5jZ
qL5Uf2HzpDmWc/YFnixnwKnrv6SzJU5/3UPVGYWLF/gAkSucUdsgr6cHfq1HghcD
n102DvsUiD4qfYiQMdJ2saw/kSjTa6stp/lemllwXsWcPyr2FGUI4S9Mz3ofmXYV
MkNmKI/LcIm/TvmI1INhwEVNagHwLNwlEQI/CWFW4bSOtflyJHNs7rEmizkRfnPF
zNPaOHLHZ8/3a9L7CZIDyD0zdBb4UsauWK7BFsLOGoDa19we+XWE+6Jx/hVodMh3
nmVez3hjsTcOjJdRlnU9mkazmeTrZVfbDdzmnS6Sh5ishsrMkk5HfOd2wWD5QiVA
Hb1ZK/F2SB/Xjj0s7Y6ipPHOgif43cJXRxQ0sVmtp9r5TXgslIpRpS/wW756bAFn
5123CJSjg5Uh/Nxu5bcjj3GFi5ygkmNZnnuRaXnmnjoIe99mkozaGcz/GqB6g/wZ
1DGPgAsOLLtsLlWfRlIA91XkVqiWYVE1A6E35rO2hm4mmRgKySFM3YDsTYD9qhS0
ZFJEXk4Q1k3+ASUp4DB+DVasGLBTqAFyomKCRs2AKjIjKEmddH3dq4KNF0wtvwkz
AeO2j31p5L3nXmp7SY+8sYpDalzrCM4i96uhIex/Rm4xpW12uv+6CyHZAXFq6jAR
jeqhfTyugx6H6Caa7CyNIRZmYwGBvRfh8gHlv32P3zPws84w2qfk8PKZDNy2/Xcp
iqp/D0VcPmPX1eY+7ruCLnizjdT0rY2z4GQtrRajgL4vDuqAspWgo6A6VodBG45r
ImpAL+TqBWhzBcjy4FFmmWofR2ZIcXl+2xiNxuKjwYPjxRLH+fJ0KdS2Vh3PObrW
OGHAuDhqxHBAEEqQXf/m4FuDdCWCb66GhADogv1uF1Bsyl/GQY4000O00p00OU19
jIe4mx0j+HessdmWFq1vSToBLBBZB1Ki16f1ua7LTsVrXmREZvzZbd9Vb2CVL/Fi
hJb4ySl88oAiLHXrlP+53FoitplQ6kVQzbX5r1tVaGMK89/M7LqeObUCrF7G8S2b
8S0lPe41i4KaJlKFyPAqk5ICfZirAcDxMaCzSJvzcYmR4In0EsRRiiFEA/7CUJGn
75SukllhTJap/aL9ZcGsiM/BvEE2jO68vdESQYr+w8a2tSujBnEIMNCjWb8FRP4B
mwBQcP8ef5GVnms/FfVmx52duc8JWT3cQu1U3RAKhZBx2FG3kjYXivYlFmqoKdeZ
kFiR+i73Rfy0sekmf9DF1N3dK418oXM/xN8Y+Y9/Ldbd6195uzVM3Hg4XTDPK6et
kiyBHt+RPnpCo+hYyZKgr1BYd+jg7qgfgzRXp1QR2OLIoXa6bas37Cx4GS0mVqqZ
6HKBvc5cI9WysQiEWwy6MGJZ0NZww2hIoHoR3vnbPrPgSdKdtm4+1y7ovv5HfSKI
/IkShIBFerkjRv4pPp4ZkvW+ufeIupMXwCLK34/YY1F1iQsT7BC3Vm4vRBnIbRt6
bUy35yT8y2KT8WtZp0H79zxVyzwOf+/UzdU6WFlEDOVkg3HkrF6okpnvJxF/5fc0
Hfhg1cYflDfy2zjFwkF3NyCHcFnaE64t+Tx50GWzULadEEtrgR203Gaz8KkS3z/T
LCjER2+Z9wHxnIqe24G8TX09pA87KZE2NYijWDcL9uXkeWwYaLk80sKnqTs7kVS4
aI1izSf2VNGxfzr++2WMTIOwX4pOmoBbgbpLJBjEu7RQSyTpjd+zq9oyIGTFDv0c
wbfjecpPsPCgahyMu4sjLoMXq/IwVURbaKiK15uQYoeOXszWQk5QEYrinxAuChlO
vKehVNradIbqkRzUSz99MFrTrUVeL/976vt+FNa5H6lNHZKznub2XBlh9TI8G2FK
7YeCvQbJzXAJxp4SgSQ3ErUxreY4A3lyK5PqrL4yLHSLqquxVYMUlbHAZTIl9qb/
Q841kdbvpoAi0Y3e4WbqCvg9hJWr5pQyAB4oa6LNO282ew3hPT5pt/BnJbDOSh3+
4PEIEmEduma8l+TaH3Gzl4ieuo3k8R5bUI5FjBWxEBAbivF8//l2E25ZPFPBX3zn
nxbDW0H3mGhF3LUL9DbXXFym3Dfn4G1WYrfKd7OH6f/ASN4NnHdBVq8FocfG/g8Y
PgykotVA1tWO3tOx+0h18Qc4VyRQhaHJJJI7sa5MB89AE3kgRHL2SxXqOUkl36Mk
U3gzjJljv9Dym4aOBvnVVGMrUBMzh/T5EsPDYsFh3EE2BQip//xnEiyL5f3ttzPf
OIpAUP8EE5134jUJRuGKyzWr3aBFn9eLBoRA16MwDmN39CuNWawIglgKI9xYD7lj
Re1J1tNHCnWDRDl3vdOWuxjwyyO2EL9yXvq6BPJgVyG9yMfNlaz2ueNO8OPHvHbh
7zSTmdd6rtvRQjpmoHtfVx0rb9l6c2KqSyhdkVajyT2clhRx0Fy6esJm0DocfKSW
+A7AASveH0/fw2xRIkiokh5SpoCe5x3YBIu3gdA/4cfpFCLUyLM9V+RB0pUqtCBH
GvBWSjUNjy/G5gI1pfiGk4i/UDUyOqVBclYTU6DDOGNuVUySJinCvgmkr/YHYEWO
cYPoun989pKlRitFhRTfiX7OgYhZQCUD6wyzHBLonKDtIy0gmyY7BOXHHvYPTAZh
0O1LHjR0aVss5e1MhI+AYRw/Uoj0WyotGnvma1X9rdi0igt0CNBkUsXs+E3NYEBo
IiqvznItv3en1Q32jtC6DZ37C1gZTJGlEBxRZ4qepexfmC0aIdUUdXErlrS9As3R
4OIqEc5lhs7p4BATCVjWAYJiMAWj7lSmmXjH7pbrUtZM29d2mSrtE6vz0Mo0Qrc0
XduH/WS9FGwI289CZ4opG4j2feD4rwxtr1gLdrZmPSrC0L+GnH2q0fPfoPvd8vDR
x+XzEzuaaq4W6mJCvPp/r9nCPq2Nv8X7HAcNhrhJxMiVn96jYVEZwZo+vz5YnETU
YrKyh5vGO70I/Ot8TDH7O2LDNoixVGjIwmlAmd4aZV73X6XBSI1j3LadqF1VHysA
oapngkqsldqnaTwBZO7LjHYdqP+hgNNBVsg14hbkY5Gj4B4iQFlr8qY6pvfY65XB
ccIv3Y5ydGLE+ZoZv8OsZNBLX/oGq0aNxdLms9ax74fCvitYZ1CnleK/wSGeAwJS
vEeMzrtKUErFB+q7dUFXoXvKcHvLjPyN9QO0oUQUJT/oLK18sr3AZnoOMqj0bGvN
bW/hS4euNkGiHSQxhHqV9w==
`protect END_PROTECTED
