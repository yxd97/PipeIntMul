`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SDgsFg8oZc/VuGKBhFGNn6t7LNX2ZNijvYSL37isHSfymB0Y6O+jCUl3tz+1cETs
4SNJxiTEO10KOoYdlkS8y/ItAtpOrfBhwyzvTQLLq5nU1AKnv9dbaKDrAfdO4hsa
TNJR10EUZ/k9ZySElnaeBwwHkb44hJ1V8NQXXwCRIy9FvmK7DWAsAI6btCjMpCqW
2v6rGP17QtuXlLYBt4PCfBPW2K396WNf95wGoFnbIC4+oIAXyhJb5u5ZEa10yxUB
6lqazyGyiUtnNzBNlorTKhbqf/mpHCl335UknI3yH0AaDo4rihQSdgvAIYJPgN4H
OEubIQiLFm2D2uZSCjLcL9SM8KqtI1IUuKcj3KdjfXJOjlJ/Zi0QJIrs0XiVbdRQ
TYFsVjUNyw3z2ccFwWaJX/BAt4i6oVj2uSqx2VAHDd8=
`protect END_PROTECTED
