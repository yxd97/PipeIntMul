`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
23EFkvG8hKgMMbSYlPC3kMSKMOfAnr4RDc6FRdjt6UtooO0MEr4jy4thJitgyZ1z
SvcaUgumprOYvSDr0+UOBIlRIK03BclbV2b1KQ9x5LX6H8NJkQCjz+HvPCFqiAqT
y8GDamHgCNjsYPibTJplUHgkBYxIGhgbvI4eb9jfcB7V9BvT0aDS53dYixERglGH
nVMIpSvRv96nDawnSGI0jN3OSEBLdulthG+xnXJCSuubheV2WIV7F+vS75jUwBEr
7oVE9dzkdP81rEEiXCZDpo/0uazVdFQLQifyhd6os+y1cI3/Gq+I2A1Ksw4UhPAA
X+bUwuz5svicP1e+WEQi0a3AUT8zDR/iCbIWLiWjats/+WSUloBC5UFRcUyv9CjM
m4W//gieX83MbHqnwmzTpRbB8p07e5zYFrn4uEY/CYI13ZLBYJ7aCh9kDDt9NyQN
lE/m9TrgbrfUdqZ/MyLVZYRaCaqoLvPBV4q4QNay+Fot7+AZe1V+LlzNJ9LNVYYl
`protect END_PROTECTED
