`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zw7TWzBue+xTOj6P888RZwbmp4V7r6lHbmu8XxX4Bb4fqTwYVp57fD+qAHcTsHYN
kXIkdjQHUbSPh/tnecHgxVvGB0z9NcSBpmcp8No7UG5jLRLvwI3yKzh5PwpLBHGz
e+QZnLyR3N/pm9IO5zvxUZdQ0+ogVr+6xhNBoXcxEuAwOiKKPFrwzpp9QcnNgF4j
Q2IH/Nzcnwa9J9qSJIdVPPWb1h6alws3MsUrmnVpaqRdPt0tSktnDZbmQqZ6ww4F
va5pHgFwUsUl6syB9mJ0ch1Q/zgUgDk8cnY/igibt+sOfJOC2NNrRRgx/c6r0gZe
TLUAvkHnxjK08H2f9RZVsgrcaRVcEoJ1ZpDlNtZV7iXaw6O0g+lUSz9pienzYRgO
8hYjkZ3S23nkbAZHejPJmAA8l9gJmt1j+5Qv/9WITGfhcryBWGAreIn6WpD/U8kb
LVv+ACXl2SN3I9by5yb/RIl0DiIp3xXiMnzoDe57ijPEvLlzraMs74fudu9nBbMJ
QpiccR0zRgRCA4ejI3J189P9jRay1W4Bb9b1EudAkpQVBDbglv7WbkjbGy5puo32
AbbTrPYC0SKYgcV0U76OZu1Lfg+XUKG6YRLxr+skR8p2Jv4W/a7atCafC+mbsO8+
mD0srGvcmcq4zCBWiVr3Lq3WD21iXj7Fnlv0u7WNyQDI770ie+OkJErj7pGAbK4z
xZd96LSz2M2ujhANn1uPHy7V0GWMTxdZsYwjqFphnpkNjOE1xmdS9fuLcH7WBVJe
V0dQ6EFA5jOLSpSOIZUX5gbS4EBNxxo0i4geXWMCBKJMcYnF6cYGnoKZuuXSIHC1
kzjPx9RdwyEcxyNbVu5zhZYjfjIcEQ7Th3zl+2fkFfjR6McD4jsVpsor0RTiuqjq
d/jUwAb9m0fQpY6Xsqyr++gfPFv8q+YR6EYEYwWF8ArzqsEJPXuC6sN1Wh+dyc/Y
SF/TLzkCNsmV565hYhC9FhuB53wZJUPTbr9TWFreiD1SpTSB3sN7EbypNfiKynCX
NavAuLr39pbXr+VC4lgqfosja0YBwX7TSJCGjIS9oOJCmLB/Jbl53S1eoC6BSktB
LimEBO/CsG5xRG8EqYDzMElrDaTEuGKTItMB+qTuAdWEpQmepInJ0+QWwLu/n7KK
PwVF/t6D/g9kl3SvkVyQ2ntLVLEnkRGM24HUgA1N0drpbQkKydyvh/eQ3DR44JhS
mFnNwu4xPNoOuaqMw/NXZKtrjEZ1j+YXdmNYcUv37D9QCvFNhVbScoiLkBPMRBLm
qDVdgcyDgmFhBj01lBjXwy2eq8rProrEjGiRc5DuS9LZ2W3MBCPSu8cQy45bhak4
X6jr4oBiNy1iPUGfG5c1SvGqvXY6o7/6pvm7YSSoYJgvmOJHj144jeICZJyHBKt/
YtHyN+DXVw71YYx5SvSB39tBk1fs+7N61iLvmcWvfsOXVQfBbSBpiKAdLN1cuA4s
kY/r6TzhY6CSvz4sSjGShS0BhpMkpP+KRTADEqTaevN4IZrh7ISm8HaorGlwP5tq
e9JMO/lebJKEGwOFZKlQKb6ECYpXjvGMB3njBu8XPzXDE0eabJmsbIC4UieR39W4
u9hZNH4YevQPBkRC3eEvtnWUxI+mFkTn/bk55b6IrTN9xoPtgdfSD87iPqAQeQe5
ctJ3EBylBsbKiQctqr9tbLwKMXYNHcl7jpDKnZnnNvZlK0xPR2GhWWwwDKcDC0gI
/abKwBd69X43RIt4PHuZDdTEl7EsmWWROtuVkGmnv+/tKbkjRr1tVMexWOOK3AQ0
DLzN7x09DDgzrbRwnNWAWRr7t4An2/g3TYAopvR4P9dqOXxhjPpZobYApKvIfcDf
BMEt99JhBUFKqgBlevVVqSSr4d44GSrG7Nmt99ybhPF5AsDLPgoT2/XyKvHwMq8I
HCJAIC1QzMuMa287dDCLdFq5kR2ebJGwRoRN2THRl9ujCnwv1B3yWgxzSxxplIFN
HzM3K4YVNS8C2SXqB584oClfFay3fNGjHd4pMLebWuaWn2r5eoKdp1AGUxJu6OyT
zVxU+o2mcXixSF0C5BvQNaSMdWQkT11X+5A1mpt+n6bV31+nzOnijp80oLA6njIN
3YNhyTumMZI4w1btRAt926uf53vOZrPO5BQeAUCpE4xA8InmwiOwCLk6D9GJmZQK
oIzlkL4OHupZVC7ubvoaN83MOBdc746IBMzCWV2ojZhvmTzoi3yMsIq4Afspu0Lw
1jL7gnIcCIjQhJAtQMp/6009+3SGuMfH45adwNkoHCLWhn1FzE7hYB7s71o98Eqw
Oed732cQom58d6YsRNE35fBHSRInpv5em8VKgYMFnyGiqHbxXWWChWTqhCUY5bvr
yaH5AoveOlkG8rknNkC6gTXOGkvvh/WbKk998AvFs7nDObzG1uofLoZ9gWwRKl/Z
MUYVS2Fs8KgrQAREItfsvXUsex7NerDrjh6oddHPqbCEpeLS8ZLIjtxAflrkghsG
677of1Moj+IIbqe8R05rJT1NpCKHnstw8o5bzirWNzcTfovjgJvYMcsSm5HNft7u
DOMhKHNJDSmf3eE/0L/PYfH9j1s/Wof323HYkT5cHgWQWOV0JFkA/feSBWZkbGB3
NzP4rqaaTruUH/6QBsDCs21F/598HbobhN8FdRygiNG6w6rxQsx1kfvIPbYOjhSP
R0DgsMB9BhcQUFex6lF1p2/atbreaZe9bFyZVpfllWwmN9YDaMsumRz9/wbanZNJ
aMzC0bKa6oFwS3z8QJebamgihdey8zHCl92SDmbQwAJwlEGGgMx8Jf7OwD62An4N
y3OOHnTxAkGrjgGKtzVhat4ywnzq/vGPQgL7Go5mx+P4WuDPHjCi9XRlVcItR+50
y/Q883w5IwnPP9eNZhqbbB1IoHr92LvNkq7TGLI4baVbjuyF6FzitBB6w7VG+34k
P7pLFRnBvP5SzoeUqtmuMJcDPgdjROtKvboev6ePGjJnHOFircG39erMLkKv5pOr
40DFiZ+JlVyFtPUdgJgXudp7oBDfhlChoKIrZpI/ENeGH5jlA7lt2CB7SwLDl56n
PRPxdHn672BrYeZEWnwtTSbNbV+j1WOkLXpjSKU3Q5rwb4IVyX43/m2AWeuRNu+K
S4cZTyt+x2TShZrP9ysFesHXXZ/LK9RmPoi6UC2R+rdLgIlxj+Gr4OHJQGo+0W0e
J6gxkqw/hXbNxUnpmSqaveziTvloSMQTFf9y/QQ4XhB96XYhmLzEQkJ2Ij7cNXbN
wAiKVGoVKmr+b36JUNwTK/WohAR4BlhAmqHxo8whsKze+B5aTQ94ZXxxdQSqqYhU
2bz47K8bdj5OF+Rv9Ly323BHgQ1hgH9iD036P46L9XIRrM2J7lq4DKsdoS6V1wc6
OFl405Mdp/qo7R6kh2+5g6MIEX/gGTFbDsJt8XkY+U6ZCp0wswICI0tvLB6kA0A5
Bg5hII+KFseiVbGkNgcEAEkLsY5SNTzg6we0FIzjP9cSdmYTiWS1GWGQ1Dzs43rW
1Odp4tp8ZTkDZhUSJ1VAtOVunY+jPs6oxnikj8JxpDtAZoyjhyCH2Je/hRBk10LJ
xfrUpYXyUzEo4a7vUwOuJhOXxAC48yHozjq/mlAkXYK6UlGFs7+NaHuqQ0dE6jcy
`protect END_PROTECTED
