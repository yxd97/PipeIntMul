`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8DVwZYPi/x0Z2TOIAElS6GXLsgHkvnlfFudrHfMSoYty3je4QfEsAGIwFrMp4SG
4aDf18oU+jRLbegOo4+rzPU3PsXnMLESBEwUAXO+DmidcqnSM4g54bxz/1fvq1r6
nLUr2tVd6NnAAmx8Z6fvOO0T1BT1lVPmLuNqj066bzUp8x0rjPkFQwnc+y0gs2ds
DTm6jKksyiZIQpULW0eyaq6JLjWHbz4hmrtlSk0tGTD2JLVdPm/tXCiGp6KbKMkC
Pk9UhmP09D3YIw8Wpj1c/Lpl32vKkt5E811lrjwo0HeEtCFemuAryYncVVvFOxkC
cJqxfLQ3V5en0e+W0Z25ssKXZMsAMgpo6dfn/zIampuypaWxdJgX55x20TrXx+oi
82G8r4Mmt0sPnFLhfVEF/tVYIKC5Mah2G7rFLiZw/GW9ezSUn4Zon/iQQpK96U+G
VX6vVSchwoisZhQrN+/bkwLJuKMXjCtxoyB28qghafYgkjAc0uRZ7q+0wgP9VhGt
FMAtq1IrPb+79emBbM4ms56WElGafAaPMbZDb4C9PvGC0qAZ1USgHOpqOhiRY/K+
XSZojVjXdBQKS7b/XjZ/OMdL8V6MSaepC3p8iPr8HPa0OGq1CNodL9OgyBArK7wJ
e26pXwOwDK5HX+MPZjNFgHCMlHw9yUFmZym1d0Z09Q6PhtmqcHC0PMyHyBXtyj9t
sfuFqC0tX01SwIrkxzkg76ZqDL2iAP+FKdXB8nxu3VXSvIiZVy1WwMz/lPz0tk4G
`protect END_PROTECTED
