`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4nTnWrDzLbJ3tmc1NNpNUhutqGAR4KugzkLORFAjENh4vNTXaEiaZUO5XP6rywSo
GXoHKeJFX6RfWSjr+qwjwQdavguEkleS2/hU41ToEbhI2PoTBIoYDwweJktPP0pa
kLGLDF0vm25aC7vtLrOCtQZjMqcFMcAG1WGxT6LOcUSueTtjz0N2h0gOF5Jb9yPv
S8y25iPb/FmsfmvY9ac9u716mlsxaLbhEVtEJXJgxdC5/zkLCJiP+NaaIo0AHbaB
9Ulcf5/7/sF4pKRRwiozWQ==
`protect END_PROTECTED
