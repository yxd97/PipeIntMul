`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rH2J03gwGhj6KwxS21oe2Z6G5oQo9igBYPNVQskfPpMB7xh5fl9KhspOUc0DPBia
F5L1DPbTLn1E60HBeWHhQJUIknGpsnJIWmqy1ZaRC8jj9VBe0d5K253gfyVr/D3J
hEIBHkFS551Cpi33J3RSe1MJos6TPh2LGEwueNhSE/Bd9AhE+R0HdNX8vkuwAqNs
lgjEwBYb/qZsaxBW4TesyKBeg4Vk9UPJGDgsnwAGF6AHBZuC7VwV1QQD2RTdohn5
2dNIwd6QVlZMJSVlQCMA7S6RlrtjyuamkvPhTkbLuk7XpKgFqebQHLlhorI+JYAt
on9FDAT0slMNHTUfWdrt6dgKk7N8VGnr8+HQkSqHaZTugq7zo3z9E3nU3HIsB7p+
xhQVy21Wm4WTFXVC9wJr+9b6p8rfdxLsapV0mlEZK5NmuZr2bUKR78SRIJ7XyxHD
LvOu+9VfU8jVq6LgAawQJmVvLe5q4zzn1z8LhIMRbXs+eEgCWQcMQUETxkkfKc+C
zzBn+3MuiBbDB7hwEKQ+KM1nndso3Yjht5ryCnSATbj2rBg911FtMjphaZ9J1h7R
hg3f1Ub22Qtwl2Jo1MhzKWp9w1rLHCQmT8HUsbRuloT6oAPzllEtILJDXYdwosgp
lBEv+0W+hxsnah6AGGI1fITHiNvhtj4Flj5j/xHB3W7TLTlgeJA+THBvBSXAaTmC
AvtsqolS6zHOsc+uEYYwWuCOZvNpJujaKtpvfsNDGRRAdNh9UaC9Ko+9AtBxSwzP
zsq4kelAHfVV4xu0a+DN5qje6OgDIGuQb143Cq9nyNJvBrbK5DXlaQbwjipfaljR
OOLKzvQw+Kvu4qERlZeJKtKcs/fsWu/0V6CoBQgM0D54072ZvB/4Ac9YKd4dJ5q+
BuK11B0t7x0P/lqZULQ1yoX2hWRXZvpDcB+2A8lDClwOq5TdS29icCmx2EcjI7Xy
XBW2CybQu0Cb03BJD2UvUNORtSM24v1yZ3Qmi/qCHXPovnZJWDsxiHIa0IMkJnVm
tn/wlEojgWowvtA0E9WUR1OYgN6QGxLFKWlLQrDdwqZ17dsTuesB5hDo5zHuobSj
+wxkHXt4XkRU+evAVn5ztAZdeJABmfeeyIQI0rwec9wQgOgT4b7pNx042rbi3nXZ
NDWd+A9YXb+ec5awtKrLGsYlsI6TexB5TnFUCbpRTMRVl2ZxeHIkMY+2b5VaZd+6
MenQMu/csYXUfZxM5toAuGRT7nWtzp4m7X02iCzMBI3ivxWGkOTnkUD8IlYhJKoD
s2BpFjmJaZHSftl1zuUnSt1SDILIrDsAdC/99FpGcgh0g0rB3oUhbVyhqjVANW0f
G/ypj3YNX/y7nFsnzQKqw6NeEqTAzgCp+JFUd57CiaHpdGaCVK9Yhxlge0ixW9R7
8LTMxE+fjFKRa9a4Yv+vSYS0utDeb7skEoCCR20aDfVc6o2YkJa3FzHi+13WZK9p
pq35yJXhOEs00mSl5gaXyk4U9KQqPtvIcx8pJTPVYs6AZnS/G7TqNbZUOGzBPjYo
33jnNXZ3/gR5GxXo21E62FMrVkkWiBqpzaOypmJMxtvYH4p8wMnMa5JgilcEx876
sc1V/NgIKPZ/bp2eAetlTtdo3hXpmFI6uJzaAp9bdDkufvUS/XZDjnXnk44CMGTH
6fMg552WXIBFGAzk9RbHfUXKSK1rLzf72nD6+J6guXwWM+Rv5A9yTbNrZ/F7yYxm
9iSDYtFiL4cYLgVeRkFS9rGbcSKpYViIAcJo/6X7dAKALmkR8vlvsSNF9e5bT52t
6KTKrRJhYinBbpVGG3FfYsx5613D1q4uq5yTUABaVV/4sfsNL2x6DxpH2OtAcFb3
U93ZpApZYhkqZPFagn/vZ7wME1l4qjndd/r9WvAZpZwdvBmtB9CkNY1nK6OJctru
SNGY217roqvUd3LFh5xgYF+/v6s4UN26XryxL/fLxyJSk9fNKCDDmjs6ccToAeM9
erdSBo0585f3iwr4gBUq7fhAHlk787xxErpBxoAqKJToUuEwimjY8aOjIm4OYgPJ
RxA9RMltLGajTDpHrKzYmvtKhTASb+c/dwORYn/XA3cH/yWEFX5o1vCXiwpjC3qk
5+Bts0+XSTaQv84N7jov4WmALlJN7u4OAJi2Y/0YaoL2Cew/atquHpa6oiWP9Zb+
BXZVb0OhsHhXfj5YGDlsIaYj2qeByhJy9GvcQNUdbC3qyVxU5JwJoIJhbBy8eRV1
C+oEAdiwe9p00hNgqgH84NUYXwg4vFCdu7asla13T6+zJPwhVsHc1pg4GS/fEXL2
N60Ddu3oEXoKnmMhMnOq/WqZmdjck3olMf75W994A1cFQfb9imlb1SMWK7sOp4Kz
0wMQuCXrZAnv/FPce6aRdP+tX8zw5scVvIJi6OF+w3VaNwvXFTc5vJ/DbXLRSJ8/
2CBKIGALJy8sU577zah/lG+LLeW9gzY6u3qWQTcZobmNN+WoBkvm0vPq+be8+oTm
VN0prHDsauxuRlKWroFMafJlQXgXmDrsTwaYB5mK/H7eF3ChKBzE83BI3nt0LcM3
lXAjsJRFQ6atPzgsZQOMyR7trjZwCTvo3A1o/CvM4bdsHCylgDdofxgy/5dkjddX
+xlg7Gnlfrt16ye0MMuUkxUnrQ3poU6WvKezxKzy9/xxMMz9aT5AETuDsE6FEKfb
ddlD0M2mtO9Er9nxHttt77USum4OSP7mRvTVgUc6CTS6lugG897nEHAWnGUfFgEQ
Mfw+jAdimMkdSf8FDGdM9hXIURg7hN1QVzdDtHYwzMuH6ZIL3kpZjBmFzrPq6vOV
K1B5HrzI+xzltBEH9Q9pCJEGDrI1Y+6cYeTGLOTcV9pGBLMUfkEfuAr5vMOFVlrv
tDHsaWBBTdQafY+92A0mVOsA+pDUpa9g6YntAjo+h7mTGaU2sbRdlfdrk/x+c5tU
JZfdBLAIkUusSkFF4TIkCOEYfBjnPNM7Qe5TrE5yJKJrk/nFjUyDlkcSDo8xmaBE
W6ZlX1jx9VS2AhCyjEkvGHmxES03u2OpKpQ5+Ck8d/uYUikDjF5kOJcojRF+Fdg0
I013eXzUQ7vsyWTVQ54/u/WFFGdGBZ/rAJgeHK8O/uI/QKSzE3nh3lvpSRMHsJ5+
6iMBsL8+3+DrStJ7Gal3j56JWE1xuiZqGm0L3XvZp6TNrTIuYNpAtqgOiQqCvhsk
u552wMUfEScUrgCqbUrXsQpTB0U0y6OpoWAWBllmSTsJdEt0nqVY2NrhvIF0bi2r
iYj2ivJzvhqVmnr75EOq94XqH2Fqype+ugL13LGftShAa0YFKpiFZMSn/xO+BaAx
uff4QPqXI5h7S3BHFml+nn4SogTapyqZA7moJvZgaCalfNQ3Zgiwt7cLvLLIFqN4
20U1Rx5YKZO0h+8OGvG6Falee55c8Fyem/crNz52PEiFQToMEW9OTpQF7jrh9wv6
5INhRuHxDkjs1LBuCkSTvGMpD0pWnjb4NHtD+2XMkY8Eg090ixp2vzmmZy5gVuSY
5/OrnChso//LVwChWPH3xldMpNEd8JxG1nju3Z/HKooZou/GzZ0sFnfi2TOOr1Ce
G8h/v/I8HVlgKYO8K2J3dbKeEv2vi8qAQgcD3yECcQGSGzJZOrXNNN/ixR2g8zy2
7nKit+dFph0qtr+CZVnHmULnAvUtYSBn3sBlmqQRnzLTpgDb33l9qy6WzC+plaCX
cIcCYQtjAQzTFUCKv+wmSZAD3AY17/rfMpN1gh3DJQGi0NH8GIpbUZpasO8lMJYA
CZxESOnI+nnW7SrzIqHh75lAciN/1QND0JZqDsF5EbQHpeG4PFIqaEB8dXXZpe7C
5T/oyK5i6HE+4ClxJULUdWBKQQDWSmUi2RdDMzw/0MwcT0+xDMBzdIg8jNCnkp13
FSzZyDSILgOtvlyAvDRv4Tx8b8mXV4OopOndMF+O9jvtyNM3+AVJAvtSVY0BKdh7
lPhpyzpi6E1mMxvGQfU6q9wASxFA9WqmbsRYMU3VhEmWHQspdL7iPpENGsMXW6RL
3TU7FBjhgFC035kgr4CSSZusYCTo/MpvdoidJk+14p9IKA8sfiBjAEv7mAAvy/Lf
KzhFW0vH5+hhrpVzoXM2f4Lbd5GuPIDwwrSKv1xXJUYpUWaTHeK2KEFifOsRrZDE
Jwa0EskJnImiVRbvm6t8I/0DmTqD51HNbfxUCtECfYFpE5ST9noYBFf9lTfcMpKf
x5Y3EJQgSvCHSBDpJrS3QpwgWs96yvYMFdePek96qkq0ma+fiOOC8BSxkJz+EVSo
l8CNXJ55gdVu7gE2ALn3v3n3Cd5utFdtasz6P/gC6j1lzJQDsV61ZCQS12NLIP38
KuIGkBFUpmo7Fxm6K+tzIq2N1inAb7p+ZVf+Y/qdEXCUmHuN14wRgHNMCD5oHXCd
eInL6MVMDPAxIGSOgdXAfLUGdkUmDBCjZK6kjFNNnGqJbJ8dFfAq7nCXSololwXo
4yjtzw4z1UlzSYxwRHDta8a8M0mPpwje3WsFUEy2zrUmODfdWDzxSe+TbSGorSE+
XtzsqRP+WEQxAig/2d7dGUQzoQFVvW1SCUSUz5xwiM16rPkriHPG8cwmhwwr+NQo
/bvXx2aionaocO02NsChd+0RmMa6MW7tqGbaCyrMUpCJyCou5zU6iQ14jUKduBaf
M+OoWlEabpz6nxl/b7d5xFu6+/WvHZCmagJsNJng12DXA+97qA48lWGZjjMaFNr/
wfHzogbTkZMwFiR9f32EUJeRVCSprSQxTMNaird5f2sLvVEQ9Fz0YX8ofTKTEeWb
+1VUHXVTNR46K4v1sIyJ7GW6FWrLGOHQnmaoalfkrHn3ttDeqL+cBpExJw9D++hQ
C+xte9YxmJ5xn8K88dbSmu16yOE/tPiYRjS5VAApjOLmT85wnWl2OUfJ/DQAVlzS
Wf643fsnJptRqCQQw7Yyh3OZW8gKBC8CQOouLAqQCWDaJg02UXZh3lYRi1WOhpXS
O5pDGMAR08U5wGH+b9SrYMY11/JcLvq0KkL0hDzK8DpwjAK76Z/3gAFjwqloNBBQ
A3BzKoEZrJOJavu698fLIEqq434zpPxi+SDJPA5HJdAQuAJx8lNbKdW1n4PGbyE/
QgakIO34w2n6rVWkj4dFrQ==
`protect END_PROTECTED
