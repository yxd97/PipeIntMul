`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KoLdaT33x8mCGgY/fVmE4B17fPAsslZPbVyc0uIhuwgAUVtxj58c/xClUgkwJ6Cc
v9MfUI5q0jH4vvtyJ7JtzXz9Hc3X2fDVeGAZTfRIHuX/yD7edPJIwnWxIDlFbz5q
J882uDdL7jTyDC5ohy+yQwxUK48uJegWj/Oco0TeaHfk/wOuAIvNgU3XQ+dpIywn
1SUw/Vqk6opA9hwBSpgH4dXFdoCGzcOuS4VzvmIR/tlCXyt/cSJ0JJOCzjQQ+z4k
KX6gAIY6d/+gPJpAj4KCP3kkJdLQPfORGSF/YCEkzor7ghm6RAWlWOLIGhFgqDvp
eaKW8+kv331Y4z3m76pMrnqZfSwhS8RGBL1Gv1XOvEUlo8/pJskYKhMWd2EKmE5O
zpaWDqnM2PYYbQ5kOLwOCeCqnuZeGCjVSY27h0vzeObvOksPfUwHguyALsaJDGep
Ch623z9RQknqXs7amOS3s5l1iGW/5dtIgk52ok8u/bEwUfiaq884Al/YSBRaxA+a
iv526iXEe1+0AyXnx4FQon4dbo/R43Gm+t6f/4nO6B8HdZPXwx87YIpyNYZgvLuh
NUNz7CJGNUbe1vmZ5OeRgb4xGwBQg7hPMbgmANqiu0k34Th9gmtPejYl1XK+3MrE
QCCC/nKf/A5Tv4aRiOkF7Wi7jR76/jyInOdiVEs/phHzeDyvTRwGRTwqasWiuUaN
m3K87WeK4On7RVy/hieXfCpFyX/O7gbdt+cYZXUuoy6f8DyUX+Blp2DS/zLNDoNB
mCjvFIoTi1iOWxj/W7sd8Jqnns0u7Wf7I6qVrWYjrCRexDK/DkRPCWNlQgwp5VpW
sXZjp9/54D44GucAI+ZYZjZNTX+kwVHNQXZ0XRvXKfQF8EMSnEUPm9Iib+Tgljyz
oS8qLg9xLFOGQZHXlbrwppK1M2HlS05jfrF75BBCbDdfykDZHhF5/cdpuqmzusdc
O97b8QvFYi9W49DSRJ+NttsP/zo1R3jlg0McFeP6NQa7v8K1uyBbEzHjh1F8ntvT
x+1iQ9wIwKCHxp0GjYwEuAP+aVOs6bIht9S0VGa3IC6fn5btVJmyq4U3s753BXsv
BKzQxBqKL8jeEvgFIH7Q10HwY6WcDgYTtQxrRlgBn7BWtFmS9ZgOcouuYLjdL2F+
xv6MMSdGM//yz97WUs4w5bbnjZjyPlMBIF83s0kkaBxn6EtYy5MV+CYeqoPV00FX
FxrZGzN/aZN1Pftl9iavMAv1ylTrwLZ6xFmabWsOLBS5hYFthwjiqmW6ZS1aIi9V
Tl1fR9bHrLO0Dtr3VrpOWTZLeNEHml7xc/lk1s9Fok3wie0hG1gAf/CBC8x7LsGy
fMFCGyZefnNdYT5pbSG2byMajBzSlTLmjc9n1s+aOMYy40zYhuHRLOrJpMo6iITl
D0FhD9A3jntTed7f+uBm9yDdsWsVOlewDOz7CFwrB6d3lGtLefEDcql3xdLWP9EF
DLQYPdvDJl8szBYmiNRSuzY9AlCySsSb7egI/OVjD05aoyB9bMpv2/orjovQGJLv
QUe3efWc+0JSoSJ8F8MvTxGqQ3vYsN2qt+na2syOOftSQQ9JLECRvavNmp9nx920
Ld4oXZ6y6527h5uMbYak56JECmox71FfeC31KuMdpggejMJudFBouvPhtnqpaTyi
PvNZLwZTJsaolXEw0Ua689le60+wKWJ3fI27GvEgMwaRKkMtam0/lN5TrT3f35yp
/Uza4dWhAEebfuIY4GEkia/jpMMl5mZCjFmFTX/Qskj+NxNxuFPjgGHf7r06tW1x
i4SI9YdN6JFchpatpOwQSRls9i3+/L8amAb3QwaGVepJFr8ob9IvPQ7QX62FmFuo
RHVlwSV/bbFMdm23Iw+4447/rMCoxNT1nVG1Ab+uW5tvxw4dP8jyi90JWmVAcyg9
M1W4NgXA2VtC7RVLdmvhvKn8nraf4qPk9+z/90R4zumqD6BIBlvRwEDA1HR0lTjH
a3pKS5uzNyxBIObbH8rS74YSSkArZlLH14LGdorPqzi1D/XEzrntoG78bvgFb2B2
CS+5vZoifsW0NVp11S75gObCIswHwKiRIzBfLIsHnsXK7XaRFXuZLcwjahMFv6VO
kToPJFbIaPk7nD60AHsftAN8O9c5gQGuOqtml7RDmomJK8PkLELORgTLhnONLuV3
DD2sVdWKw7YdDLnc/1qllZmmT/T2Y+llsHOVOBoAyWnbKXf9yUUMxnLLTKEh8xUr
dITBKzOej4/tvvgQuYRJWlQIivEZ23ohZgXEZFDW659RkluZ+B1AAHL0Xe3FwJ+0
29kdxiGJGaGo2LA5cVULPmUWnEVMtsf0PYnTWkpj59la2qAMLF3TX7zOMFGQkWC7
ymqvm4PRcsV1OKU2Fx/apY0ywQAP0m3rHn+OfC2VZI9VRxBqE5E5DENHFjZv9lSS
sWN9Qk9wfb+nxyGa6Ef7qx84wfOYXf1nMVg70NVLT8j8+6/9YHbHpNcZDLf8vm9t
U2byBdGQIl6LLIhKRNt3YQsayz5MMs5gTsyA3HArFv4vuDX7MoJPoVw/fj7CMeM0
eUZM9j5YtPCkKNsbIRTB+i+OWfmNbB72Fz0g7NZhLXrNzzYt/AtWr0UQ257OSKa/
JFYTKRpAvyBt+ZiiwX+5fj0fcKLvB3225YZMRvWSyLSr+WWL5nh1TCd76EsYb7qY
suIWp0UuiURRa+qNdjgTDtptPcVjj+MiKcq7kHsEGzoogTvQ7top15Da6zosZIYd
GIkN5IFRpNeAHEXCfpc0jETgn6AMqOyRBuII9AU4gf1uH6k5WT3+d7TQ1XjnBj0U
3lSF9RSCwXcR6czLpyDG0UN932NJhlf7uJ77sKfcduknVizbdHXDf4ROMKaxqMMp
x1Ir+jFwIyobzSxymoXSIfdfOL2UD2/kL/JLhr6g4LG8hWJLmhSln6cUQdAGsetH
TIlOm5MbpYT+hAbWsa/U0ep4zB0BRB7r04J1mIiGr/r0VjUkD/kqv/OMT5tr69mW
hN/2NdpcQgKg1KAA89ZAOmAwVEVBPzPjkL/Pih7GxTu7Ppi5IvBp1oX+RVfzANm0
6KymsPTyHo1Ul7cnwyBOAPXXbMidKvaaDhFBVWrVsqL4Gocro0oaCAhmLSHJrIgn
KYxCiB9whY8H7hoRVHf3ddQ8zA3/FjHy+p8gGPVDtJxM1cTYIFoPIaS0BRT0khFN
nUlmSGvrZXq+s2DzCSw+7rq7BHe1ojjovEBnVq1Xq/XYMtaIjUoNud1CSiAlMoUs
PrMhaINezIAh9nsPtp8ZZi+PAIv79NsfWwQ5GffknPw6J+0S8Dp0U4cNHPmPvGR3
3jMSFr8WcUW+iQOidGHyU0e11JcVoFqo5aVx85Cs0tgCjcf0AfS3KIgRLm+/lbG9
1gokjMdBL6At324hBmLMOxsBU5qAFQQB7mSnsz/InQNHfvhQBvSRApInVJe4+ARD
7Q5m0Z0Gn545lwSIUELghZd5LQ4grBIzXt/lrNQehSseTPHeg/rczNa1m24JIhFL
b+vUtjRhjSoCPLYfAeLvTNyMo5tcjv+87Au/aqRBK4f2JP9i/Pj8YI2v6WSIVQm/
uXg6GAre0z4s4zdb6ynlUq8Y17JYvTthq0nnG8a3mYN9VNeAmhv1hRjJQU9kCZpW
uaWUnsxVZR4JU6BYD8HBY9Dx/wTX0TDnFGC85p4u/7tfdXMEFntxNU6NkFySneC3
C8+VYDDTNn+NftCZLuLgYu+ZxYCfM8M02laSLVYE88SKkdJrRvHWUKzi3clprlRN
fwV8cBnWqzk7absteCNJyXfpOujsop1ol/ObygjjWl2eo+9gxaVO+i4Fwt3sXBE4
RVcx0bbZuyhv58tKhY973sabfPxqmLLNDokPOq9/pQtieOHx4kwUDrUQ7QwC+5DM
joodhLAaLdosvrQLcUCQ3pqK+LofR4fjprY3tV2TSNVtDu8n4A/O/WxIi1529TDM
r20g2ZZYfFkSaJeGZNswzs5Ts4y4PsUlE1QR0FKO4YlAHMYtQRTPzYUMJhtTi/r7
adnNcg+9MNsqh9TLPcgXbBILCFad0d4MIWRoWeJajzhMdTqzLFBt4JVlg8G6oJ8A
5L8LCCA8IbH2SUXqvmpNDQNQGiNVBXiRT6hQHb1kFmeWQGaCuOpiLbFfUIaNzdts
sDp3/jE8p+XWuLoaEMDKEnFyHfklclnLjwk+vN1O73SdLIZHL//B3LwFRuQSy6N9
EFL1aOV4+7YvvgoaCUV/vsuoNx2wllmLj3yuI57J8Bg/hfkCOAD9k/CParNpmCGQ
A7tmOq7XQfDynHWAxCFbMmRDjjnHaqiwDTWHNYPEDa5v6ODP09+I19WsyRC9qyf4
cHP7KnuRPjUf9qCPifK6TVeO0eHWAGNRg1PaU4UNrfhWDAn+ECw8wCfbK0otZt2U
BQMUir2ljjpbtvJ9pB6jtbns6BFFDfAJ+r81ZW6eWZmMAgUeE7oSJUk/2NYaKhcU
+llPP71QHt8mzZlO92vgrOnezIjSoUKwkhlX9Q6p45GxRa0ZBKuzq0Gg5fSA5tfG
BuA4MQnNZNCRsGrNSoiX6QY8LwBylML3l1x4HtT2WutbEzOzFsJ2y1hWOptlx1yw
utEnQhEcPt/2FwfwMP/VZLcs1aTxRd9XXB0+zUT7+USKX1SKxFbZZyWHmzlqVyM5
jPZLN80rFMDWG3XeRb2KjbcrVlHAR0zEBu1gOMhsytaKjFAIn5psyfTkF53DM2sq
pUzfo4C82qKd0EPrHgqN+Ap1dLM6f6AQ1r9FmJP+suW4xW5aP7ryng3i1VpJ8US7
e4O1NjFFkhjx9X+69TJUp3MSos7X3bc9PObugyly1vwGo764sgBr1E89MWHxmoOl
ipyHpE6BJstwoZ2gfczqlGq58Hug1kohiODxQgyLTzLfHjFxHjQmG52snLtyb/KQ
gnFHIp2o7tdJmDlcV1S8eq/3vjQFr8SqDTkDGxAexzPwox/8PvPfZ4qVtwldlKEj
/OmlG1DpuepnS4MVPEqbNDrag8BoZhO90IY5M4oP8P3i151Lg+wsT7/08KC7DxQe
0E1RfnbaF0MZe1lisut01oA5xwSFxOLvHK3j5zS1Y1O5b1qr+u+bdGW7LC5YcRRl
CXhuTaNgFf4OWENqygMWlvTptmmT6OsXfwI8PU3gPWDdQ0Z0mtcCsoGjd5UaX1iC
i8hmhcaNPBDkM63iTB15jV9RC1+5BukauTP4MHV/TAVvhwBcTz2NErZOCdfPfHkb
9azpn7k8Iexu2KxM8XU3qEC9k/MCCvd6Cl7uqAByG5SDzebQd5b7UmaJTlfWZJbZ
fU1d2Xanu1hU13hsSYAVRXZfPw1njYV3QfOGc5SL5VNHQd55hG6tOs7mI5gixSmR
tD7ijzPtXRLqmGVk3V1rRGciHd5g384xyTsTR/Bu1/ClkldIWJmsPHZSxq/BEtTX
M6t08cg76FET7q35LRu3jMpqSAfc3ookWZ+9G5Sd41X4u+Yx6pZ3D3/Sl/TE2pL+
R3OqyD9XfbUr5v2xPT4UrkiI04K4X7Jo9vz2zmSGs2662OE8baXCu3N8ZErYBz4E
jTxcI6xKJujuyO1RsC2ibUn+D0ympQeefXfLCJzrgJ+lQD+TmXpV6ytosY9lKgVC
BT6ntQDmWEIj0J4rkNHgh4N4/ejYvcyBansnRgrxxniVCD+kyl+hZuTKMz/dSfhP
DNvy6wwsyAJ1C+nj6N3+2P8cAiZV8NYZR2snjJ2jFM5abrXL5Z3fHu3/yxQuWgYY
MIvaf4mrHnLlJL/DAwpyQUup5gCeRTMvm8FKjEWP9j16632J5roeEd0d70vQiV9d
YqPGv901D8olO4204P/SOuGL8f289qW0bYZP9d2GU593z1bDG//YkN0tu4eB6sr6
xfIUvanBrlvspycZogisDzG9hJ361x6t0VIv5569q7ADmYLlY1AyTCIaAIsMhJYD
+4OMY+vRF/KwE9iIIeSYWnyGIfoa+mGl3ypV4kVagvyWc3YVdz8d3L59bxheS1Bg
yOxYp+1fhis7KM5MbAQdqgXwlTFiUuhj+OyLS6RPdM2qQN8/H2jaeW9kEGmrP5L1
bd2DcbNG/n/qJgpiVNiu3tWjR69OqvOexCxa3u4M4BT7uMzeeHuoVuU3sGZteVCU
xeFQliw73xNe599NOOyI1zeA4lWksoTt2ZCFxmlm9jCWxOtMe4nf1lqMCKFdAFVf
AX0gf9W6Kh+yoLTImKWrddNCrBY2ck+ijWg+Byw8zWWGQHF/o0Fz23mGSGUYowZf
fR0fLD4qbW7z3H+R3FFzzCwr5ecHJvKRUzCZT/VH4w6PJ0gvRHwPgxxlNIngVbzU
XtRJ08LNLFmT02OxH0DTi1gD599Nk3YJ8oulYbpYz4sQAAqHRyM9/rWlHhXExP7J
vn7Gv5ZgGfXl3DXbOlBTk9kGJ0wg5DVSsD5llw+J4eT/xrquFPZQ8bXp9DGYwIla
UK/noTjX60TXBDx7VBTBI6xq45tXkfZHpolCpPW9OS7NjM7YOQGvxW+TDpXE6MEV
wAY8OuYZbYNLEZXQoHxA27UXRu+NbOrD1Rc5C3SISd0BVeHc3FQ4DivzR1Tr34hj
N0K3NOeIqLGUx/a04RmBJhjDofcpT4fj7xmiHdQwPNtacJS4wL+ssMJC0leACpE2
1iVl9naTwsXIQ0z7H6OKoBd8+vygR1S34IxN/epO/FtfiAkv3VMJHc+k9BE5Lm21
WQ8t0ZLUAMRx28gsCUF+eCPUFavxMHUlJyth0x7O+GQJWSKb6ZR0EfBD+vEziyqm
10nRxRaKB7MjgX6mRihj5xJj7aplAR16VTqRtMN5bBGeO4SbXlCldWBg/EMx2Fhw
EyaqojDPU/gb3AU1tI/IRO4V0sZsY8DB99pgxLXsUHn9S/pa0CIzQlC0NKibJIDp
pgq7xPR+Eqa2Ix0SMYN8OJ6/QLiOfaCCv9dwRq0DR1ut0B9nHR/Ar+nLT7lfQpHS
J/BsaBK+Z8J7Gs0RdvbCOqtaRliYOemmbfgU78De6BN4aLya2Xx8jv8esnnwDJN7
/KNhClVTAgz2wi8+HlEo8vlv05mG5rQhu3dEQXsipKoZyk7PvXe7H+YooNG5bVBL
VhFbRQvSVQqfYe/4/zpXBAD6BEd5g0BEO5PFya5mCRG3iWLZg+LGiwOerdPtwPRd
lP6iIcA/bsI3qCKi0yGHTrEAIqDVhOpy9PIkbGtxvcA7yHQGgZQBscpyg4qkuQHf
wQoPOE90TudPHV8nlUA4ibipVxy845yMgcrNGQFSRy7bEFJfUXcO0iLfI30b6d6Z
SMW1PYni92N1mm6GQWuXQQ2ZTuhLiyUXsxUjhUi1MJdaoRRwo3E5RSxF7d27jTYS
J92MZxsYi5IljhdU1RdJxWCZr7Rc1KQv6L9IImiIYoo3WhjHHFrasnnkzKckoaQz
lXizNPLK2eCeCxJ29DzasyEs8lNMZVrMaeExK0/HfADSjglm5kvZTpfGL2sY+iBW
W+paFaKs4HrEcnENd9WvpBh4SnQNLWlOvciXNFpf0jKTHMnx9H+IG5sVrloYYe0M
nlocGt8SFP2bfUzftvvYIjW6r60Djsk8/eSe9wmX09/hvUYbPjTB3sgEE2cp+7KE
6YOlAL7wPqWkWdsbZ3cgTLyYdALl5GX2eaExi0RCd+rxW8P5rGKl1MGyXZAcE2Bn
e0nWT8pBiBvv+LKdx8Z2VYi8vt3+pZptZb0ZwOkj4sl8PlWepblVVgO+dyna4owm
++jMIhvyjdo/6saGhTXqH6kBPQkyQOxEwsE+OlHkrl7rZl1omkF7Kwmr22hyycsG
HxRE2Vc+ysw0sgRslaTqe8M9RuPxKKhLKTBtyB88YtasGUx/BMRNwwAiuMoJC0hu
da77kB2By1yzATLDoDgE13CoO0FA8c0YfIdz/XE3Bfh/pVpMSFVnjVou75a2mPlV
Wh2ulEsY0GCmd3IxCZBhNe2Gi05etc9VYeU1CY24NX0FpJdx4BhrO15FGwRoLXz4
pEXGagle4FS3DoJp5osWp2VTmxLdLneapTPx/xGplN6YEXtwBVbZy5++39dTjUrE
zsJcsHDKfpdFBrUMuFK+5Sk8sQ0hzDwJjJ6eGnKIDSHhmedaH1424QaxTjwfVKz5
R33RRjXMF6pa4KBp7tkproO8z6mKvJASS0rJK7hJaX1ntxR0QlRX6XpsYz7EwC7s
wp5d16517s8x12Vc8Ld1eQfkkDqO01s3Lb5E4epUzDa8Fl32Mo2smu818Ym3S6FP
XF6z1GpuzMs/kvQVVcVnqUgpysNGiqpcdbUtb03jJ/xJzfg/iO7rGxhqNESatK6j
wJWlRqytHMuRtgIxwHuAoBM7CYNI77Jr7WwTLyxTV5H/Qk52aGIoZ4VbgJsp93yu
z5rlxytTSpmd5xA1/3AjD92ioVIIrG3wnmCasSMS4UtjccT8OH7VaWcqjLHF0RrI
MuatjMT7PbT2IXR3rlVjYfje9FYQhnv8sNlwjoM65mJUlCwX5cnhQDdjTZT37cE5
8NQgX1KUmqByjOcSczXCmgqqqsTq5ANMKUSVnTkY/XmlDkxgk0PM41EP0QRdcfLl
rxx4TTFpLVgbaEVest7xItR2GgDIbWnODDXesomMv91Jr0J2jLb2qhWIroVr3VNV
6tZ6JZ4f916Nft9oGQ4GMuo+/keJiyvNEXjxJYXzsZ1984Tp+7p8Al1y1CdgdXgP
1v+ncwllzCa2B/CYQcXmsRrQve7g9qLMqq1LNQRFcccEtuGEB7FWiAZPlvAysUu2
tpBGBPongknWuZTonodEFPmHBYoJfAuyOVEyXwr0OvaAIQVY8Mm2TEZrOpf10b4i
dE0qVo35jo7Xlr+HDaEqWcNJiQ4G4raQcd4s9Lv8RV23XCFSajzhnAOPsb0dNjU/
ZmRR/0aABEuikSBX0ODk1v9vR/FVU+VOC0hXapeKKIQ9NUcr0iS0jSNagjQyZVYJ
qpEIzGP1SItLxOacWy8TmHRLxkJldd8r4CnaHTWxbzSUJeVjs/jkHvHn62qlrAU8
7OchZ5yH16ePWjFLfW4NWvMgn2q9AOcF3ZaZxct8U94w+Wtyzu1cvOInD1ZezGdK
QOuhWlAlJdRioBkc/P2WJ8h2c1gh/NcuLTh4sn6V9jQK/75QK7AThm1jG+YKFUmJ
wqH3LrOJa4f1pWK35fm302cyb/uPW//NhxAVQQrdmxZx6o3sxZP35Jznfen3Ce1W
njFuLMY0X1UpdKP+I2j+MT4Wdz535uo4cxhSjeDWnu/qK0DUI5Th7aPL2wMVdlY+
OC8mwDQbH7wCz8wDzmbanagD8PYMaCne9PnjFgSy34nwLNaeFiy9PjIUz4cGHjeI
QXjwWsxSmkdAnICSq7tN2ptDqgflBKAvzkPXfoxF/Qwlirpst7G1mvs9jfcWO6y8
LnxvSA1kABZtmouyjdJfp//cyfOFzq+jqfRu4gpf0wu9fGmXxkSMwyJuO1vfzn6m
adP1osfYHuawpJnYEZwU8h2i2Vq3BA9d/H0juhGgpg6iGZkL/FkrdIg5iB8ifgYa
X/y+CZlkc40Fp1D7fdquf+QEXb/ClJGYbGl7trqanjKrniFuIwbHb8kO0yCmED2k
m/VSbgRibF5A7V9jcSsDCNJpU9HzIj9KYEvgfoCRCtM18nIkq2jjJwLF0TVvszIn
Bm+rFnqj8HzOTpcojkmxrEevvHvQFele5m/puBJ2+IDKztDSNoNZWCqtDAO7N/8F
PZGaCABtoNJIIWFC+sOSMCpkuddZ7n1hX6P2c7osRIb7+2hh3iurbh7lO9sGh+c/
kGDoo5e3Yjs3+TmlAbOHoP8+5RDnGzDAUdQC9ksEZwPeDTCB7VoGi2QMHQ93+Q4+
xZdPC7t4bCZJMHEPt2+6YrfIhH8gYiNJDKFYBvSGbTa3RFGVG1RPHs0/4lPvgDIH
HdhtfYDpsPw3DJd1OOdKbOYP9F1qq+PSKLCLZwlfMwPyVfjnT4vkteavQZKkaea/
c/2ksV/zWUpcTDKc1UgSfnhtJsUrs87TJIiL8vzVg0xXyrlyi5yKwZtoo+y8iO2E
lJmeDJgo10jyP/JMF+K2ZVhKECtWI3jY5VjvBvYXv1+5RpuMFTqWKdLdZOZ/rCoy
ljw010xmalnNBUXH+dZjTOZP/SIvieX/rZLgSKS+8gpvMHg4XdF6OnnRd8ucsDq2
gF5Aa2ciBxMiaxJJoyK9cj0t+oFB9CukKJBK/8PPfSHdh6oH7c8h9YVed7A5YBw+
CRB4ROEVXsQ/iwbio6ex6egjxK5yrqMGRPQQXshmA1a0nEi6pl/EdMCTwfru0ePc
8KUfBqPVoxeZ4iXGiqRBrXA0BIRMUz1gqcGTKsKgZOIKedYLkAf4CR7LCi9SJm3j
NnAnwGZLmPn+T8lwV4urkHAixjvrrYH8n1u4+ZA2sJEZ/OqlkssO4+gCC34BRJ0I
PxC5e+mHSnTnJFTE1Xgm9l8h76MAor17Kn0uPKQo8DLYnuk2aPbwoitSVviTwX7Y
Lk7wEFzabijff+x7up49phJpz4jhbIZQ9U47eCMqlX3xcMj63EFlbAnYSRbq6T0X
NAtpyYv7aEo1Yzz6Ufw0AFd2D6bfIC+VsNnHYQyRzZ0BYo6DERDExxDVB0vavgEG
iO3MlAjTXUH0hI2FKSfYbUryITC3ypO64y218f5st0ALwgt9lWEnDZWNRyUaXw5o
dpRHYLANurzLyzJRWJa8ygSuzegSLtM0GTY3T/cuA4Vj86pC01LIW721F8G58fWA
7WZP6brKegiwZhj/sCeTVTofquoxGDoTGMTh/Mtd/yodiuQ1bMjCEmyJkPf3xaar
/1EIpzyA1A82idbrZ2cXw8YgGltr9RwTHZAoTqbtnpCRAj8Vcyg/6IqRPNbPLTRj
Pda9gdE3JPtOoFhZM8PTpFeHEHxghWyAIfwOEigxnPx8idLx+hI+jNCbaE7TbUT9
BmpttW8XWljU/FdhS3ooRex5LzSL34YlWw5KEnYlt9MB8UlrQfwHip7BiE2m7w9O
5oghkjo7nSTUke2YFm/GZWjSwrW+BJYBh15G/F0h9D3nknzdl78qB/v1vWVoWAUw
UKdRxxDyjC8W8ynL1xDMPZtcM5e6WqrYyyLsnQGSnHDnFJkb1SyY54vpkbNZpm56
bXxVhmO7xdkahI/32uyaIuf6mTDD661MCX5U1CKpIu/G8Y8c7UugbH8IG8ZFlb2K
eS4qDw7UWwUateyNqltAKmUJmDBu6orN620mQzwr1xsi/YmWky38LCX73OSeh4jV
ah0df8rXc0/lM7EpsXOhDGQys9b3ZMhCN94v9KjjZ7XHJlTqE0aQQPp7+CALbRJW
4YEQ+KqTHeCm73cS4pN+VoeTJhNIeaOgAScTEDeQRkJoMLB97s7guMFHFHh60N7x
QuXgjvf4AxbanWYvGIlJ67SYZaMCQq6+442CR1pXtbNKK7hrttoB1iS7Fq8i66YM
CEYDGs+DPGeY03cLnu9I8SQ3otYF6FdYev3aoLSdbyqfPM/Lq05yt4VVGCuSEXsl
UXN7oToM9h3BQITm+ZQW5d5NlJqFLvwF54rvc+ZZKp2bbvKdEtNH8L64lAX+V9jW
fdQ1UCBoqujX+NIWkb/wjtOEzuICOFPSfDxLCebhXPUT7FTPx/4me/BtrOErMVyr
zhJot8FioCzchLhfPmRik13pzxejMUrNP8iB0h9yZSOK+Nghju3H5Hzf7exG3VCa
+ErJ9TB8AWI3LLa+PU0QrGDor8KIL8OrrSyo/13l6BWM99DZEkOyEJu2IjzQTZjZ
nEU9DdAgV0Be0z5ckwH/4YogUjEusZmUveVBFrzULK63lB9i8f1KnHDaLzh2l5bw
ucSgMlacKRPmPhAfuELpvigSkDkQHGAb7vYK1rzzhMJQEqDn/6baY8hEFPD+7mVx
1g9dji8HmD0nQ6k3RL/xwnwh5w1bPYrBU49N0heqiIFBpa+lBvYsbA1A7spCHe84
NAruCzPoiBo2FR7Wd7h208lTIdkSYqlZxTWzwlJ9/hIzS+oWsNNqkGMW6x7iuWM9
7kT+DMDrEp6rR3pEbxhNkfRE3ylZJMT7JH7XhrRWmlpl4XdGs2re7DJKPKqI16LJ
CZrSbcUyUbvacivDq5iOZXmo56LSirFAUVn/4YNpFlvGQT/G+QulzstLV8RxHUKY
RJX8/r+GrGEHsbDcpijzFCC30tTOT9qDn5IWe5psdN+2/lkj5tnXDmtmzC786Y9w
gM0EcYtdms2fp+jP9hJ87EhkgbSfyZdEhH6Jhluv2pdHM1P1rDHKdZVxq6mKRBdN
dglszydrPz5DrL4Niu2P4h2mV8UFFuUCL2sw3BWyXuB7XgmPDis0mAJP9kOflUDF
wWLHjk3zVbb0r+8m3u7BaJxR379XISH7UvGMrC4UlEALYPM02nChPugrGE/sJX/R
jOR38Qx9bY0C2Gkq1F7hqjXwXOsoyIUycA22vdzsOtdFoBpRANAwXzwCeWN1xTVc
10a6ilEr5sgpqeXbKg8MpnQug3S8Zniso2qa3c3y/XCgZc7AF5JHXSJRmaPO8K4A
+aXZS1L0+GLQXSitYuJlSCMKzVzHzgWuXCQtBQF8rv+d7YM9LJNrTFQ33mYvChKB
QP89Yl8U/TYMhFDi3aIl4QHNNo+tLviWSSyjB1tI2j8SY+2sgei54gKwGFRPZzZY
vgxJ4eaYpKHkiO+5cO595vnC5BVx0vdPtGBosleQu7YSQX32kCVRGL4dtF0nejfM
WGwNDWnV+3gVJbcwGk8bVYuK3rtLGr9UQbJJugB0mD5Zdk3i2BW3zAXaWUYGwYvD
WOyK4cwlysUqyt5oCWYp+28Dcm5dKKqnf/kNVgIDdCqAOh9OoaX85+q/e9zRsqwx
yGdf1tbQrWkC3F5BcdNy+BSzizkdoz/boi7mrueQKWYMt1r5CRvfkgbTGNDO/VkC
CtKjRawJJEooai6ox/9XhKB/61WYPY20kVWw/PgJlXeROy3T5gbs1urZDgAE8QPO
7Nq3S6qF5W8KLtbv3t6nZKRQDo5S39m/XWIc2lKsdz+XqvQdsVplkfrk6W61H+vh
kwHEVEgvWtfSms2Yp0dLPq4cmDe/GXCYfKtYUAGpo4KYzpw415PTZitHM9c0yc/1
yne/pOaiFio2VSb4dmGWh6sqUBofZ7Rr1kKFbzqQlQw89xiLjG7+yMgc5OTd0UH0
5cc7YLbeEI5jJcemuFAyr5zg0LOyFJKPqkZmR0VOsAPrYg11LpFeP81Iw+jzDhN/
en46kNk+pZblbH+eeIb2OHco07KWB7KT7rCcnP576o4RNIcSeySZ5sSzjBVrRHzJ
XFHMLexeXiqQ2dZe8cNIgJyIYKgf0cuV67gk8fCOqoY69jfQinTucgNcb/KnjMb8
wnuJX8PEYPtTj5VSa0cvM3nRyjOBtNBkNxBu4kDaYbLDM/ZyUeiEUXXVPe2WIUrG
C3BN496IvzI/W2AifsGqX1kY0MPwi0mJZZT0m20yRGimiUtIy5fuappwghiNRM3Y
kFFhid88NZfTQRwCgcpK3SLX/MDGT14rHu5ZSIOWy6lsHE1fv0eK37wFwSwB7cCa
HLwDeMJBeR6erPTrJLDM+WdGDkJJS+kUFYbid0SDISD3v5PoAari5i0V0hfGOPIf
ewAx1mJGcjv8vHiNm0JD8EIFWWC/9IsnD/HahtfunqLY1qUWXsiuxGJTVChOHP7v
lIjVYspNuLrYFjk+RtLS02mKI8P/dsMvgs70ZtXi/2v5iE4vc2Q7YDZALNr6uS6s
MbbceN69M4soj6g0yTgGQ7d19zvTZ9DLo5l5+7QBVABsR6tZS+LFCGy0+MSyU654
BUPR+b43KEUqgZx9RAK3ofVJT1rQd07n5CfmizFcowcA8lgArSKC6LOf5lNO2NaN
gYT2TyTb5gG6lWEvD0qCUtxleryx2JVNrsFJmoSxKhmAYn4ZH+G1aF8Lot4gIVSR
4oSMZlsX0NZkuXjKGROG62TiCNoOuzzmWqKaa8LypDlQI4YhNE8yiaLghRm70Uk2
M91el+B4+cdz8OtyhqSjPqAA/9H6pEOT0YqF9rbRnpnwGhss0oLfhltqJmJR0mTp
F7tJWP4MRrEJPEqtfjcbb7CLIk1GQ5jgDKhPgx0EQtZB8lZPLYeFBNTKk+7mL2zY
8CVHoSrpBpxEOY+K8aoDzf7jJ1MhLqvFJdtSRWmAHlQ+8aexY1QC5agpEc8fYpSi
kah3JgUhmtL/vtr8CC0FRukGDg1hTDyNcLtyE4mXLby5KYg+1twSNFFszQT3Zbn/
X4Q6CkCg3SFlgHy5sg7p4b4kAwPuMwJc+Qgl5HRlaocgc/9jetvqpFijfc2VMx31
O3Qak3PIZEl1RGZr+8jymLSxSxaqyhKdByTVMpGE3ITVVi5/pmNOl7h3ZGhmGl6m
l07qMBtloXHcSJKszadGGid4Lvzi7EztfmG4hJnfj9HVHiyCtL8tjRCnIFS4uzNv
HTfELwODIghyBKaCnlED7NqsmP+1QDINZj8srsJZnp2jsUsKo2JZoLkhZ3eio78Q
x6EUw3Q47PzF8bHBTqsRy1SFntFwwdUP0f9vv9ivSE5U0ht7jMy6YRx0PDJPR2f/
2trhpTkylNVSQtobi65QnB2vlujA/qGyuWjfxhyKxiGgxaDHn9kU8lBLY70WeWQq
8gZmMSs5gCChEMgkSNF1sJmHM0aAs8Fuf6qlRCL9DAJmBjKXL72XFP0b/4VbTCdQ
wW9l+IBE48BWTixbOvetnqVs+UMjAgznRMZ4Kc83s2qZlUvt1TeM/m4E58RlhaqP
mMVEuX8z+3FJZPZx4TlzUGURgzsgFOAGdF+hLk6+XNGH1lsKeSdolWsZkoOFjbwl
2rV2nReCOF3GwM2ORlaPtqZwnvecJXcZ+aqQ/0IS49ABkbwJToEPiApwJGr1Y4Uv
PCBQ8tATEDsRAezoWoVDDrCHgNd2nsTRxXqxabRLjV5pfGxnaoRxv12G0cVjjv7s
9BI78nXGH/JRPCKU1IiFzHFyUZLLtD2c/D2JmTXg5MjAWDeYsXLdJ5+woIXNPoUu
X2ecFh6JtVvgSFzBTugIHJsHJc5KWctqPDh00F1Qbn5GOyrjuIJho6SuV1Hurs8n
BAm32cRl3FORPVeRLJfgtT4EiOAXq/MpFcbzIxFLm4JPnQ8yumLkdxYcXCWx6sV+
hFNcYeCWR+2Q2TblYQ+iiSqFnU26lXN8HjWsEiRQ5hk4zLA+4kX8LF9LibYjKt0F
qjOx/PgHXwwFxBZYB9zeuTZW98WeiwFaRlYIcHuR/ldL64F08hlC5Fo0whkzSI+N
L9VwrUFqpMbGaUc1E60jNUcrmoDhih0BAnf/k0RbNu5cdK+tHA0b4HrHCQoslFF6
f9/F8BBYwzll+xrryYrR1TarfwP7SbyPyTRVRoYunBBdwJQAQBGUo9QzlQy6lJGh
VMAskVHOzxQYnya5Q5cqSIvPWmUBsuLxbAhhb4Ai+9NO+31H2SPbu5uQ2y+WuWie
iR9eTfbAVj1/bHDiWLu4/RBKt1GTk7kUzmsIhQBFxCDxUm294A5vfH+LQk5h7peb
nB8jurQq5kTEj6nOL44YSkwq/7GeZXY6UDebUiD1+M/xqR7obSb3e8SqKbV8RGH9
owp/vy6nNYuC2RZZdeSiXnL3TenuxdgRxrtUExDOYQePyympbJDfXxOIZ7Rkdgtj
5kfswZvfTv1mRN+1V2Ydy8QaTJgiISSJjtWQH1JOLIIUztPBfzBgSi71lDH0ojJR
9Ar8jXdR8lvK6CJGFBgLQouDJ3B4B6+jDgA+ITEp05DnXqpjL71XP5cBZlLOC30k
XJLeZHHeTU2Rt3j58t4HjE5ErXufxEAF8XxYPpvDOxxjBSqKS6hkgpTLSuJZ3HkM
AUVMRj/kqEYNZrxmZseVdEeRvwmDXcN9WyLbOc3s42N6jruCh/R3N6y/VwV8q59y
wG40YCPZY1VMsb+AW08cEH5xao15DrvgPGNxt0jbYjNJVPsngAfQUQai2r2ZxvED
P15yzRq3TfwEPA6Asxv9vfSaIZWC4Jzt78ZzhuDFC44p6i60sRqwOYdJRk/ZhjVO
4XgEtu+wq6yaRkPiYOpL6IHzs1gekjrUhev8TdlrywCessgSJm5pzXfoInJwc0/I
qbY80WK2n3HiEA/Zl3+91/hIW1J7JonLhprvwfVyNFxnijJy55+thPtLGhAV5zG+
REVBC101EqVPh6yz1w3hproh2Vg39Zkbfw/MwfBKioJONQJBczy5zF0WNIsY7Jk0
ANg66MlpPHfSASm3zCCl4LA/kq9S7jGC2CIHdBuLjKcpwGRA4Edle7k7Ty0BUrOh
KdhQ+Qb9thUCV+KDvuEVNspHJV1IdidAWeo2Wvw69bIsrl6+AiYh1+PqjksM6MgM
tyVlOfrjUecryhjaSMvuaOG7GEjJF5DBgZlLDByzEyjb4qqpHm60E9pRKlhsHkPB
eWr/beBvYCicR7igadE6izRzr7TQbiHiLixYhbfMjqfuJynSqRzb2OGqrUF0gEUy
F4/nDJR6qDUS83WCEkbTiqs4TtzJpFLMwj5/wy+e3PdE7JXpFymn0fMVOMljb2xV
vDkEUzYPwD4my6TFVsZ5pHLhVh89TEdxQHptAw4WST4ntaQEZypEujWzPr3+T7bo
SSc6qUHQMqnRYDMCSoAilbThbRtgRKrD9U3j9ebMUpgl9BTIKtyBWKWaPS6+wevS
jRLwLxiy9Rj5M6fpSFa8QYUDQ/PxFxN1NvHRy5MlwnDDwftnLs1liYUjOrg3wDJ4
1b/qNoLNT/EtrMaNpgLbBcCZEa29E+gYhGIJEHBQMpmPJWcyXdZn+wwNYOEKhtHu
TBgK0Q7QTfQjAImxUt2jO2yM1m0wv2pmYAgqzZDmCfdMUubUukdamzpaUoZl5+RN
6ETivXVaKSmU7hvuFeB0xL33CHJjgZeZyAxPiTdrHR0PxNCnh3UWWe0QR2kWdGjm
4j5MDSMjILLQ8v+6vTLwdo9jgUTWf3Ivk+g0RqBm0ipfrl9opLmorklhNGN618iQ
f2AkjyH1oVBcquJM5gsyT+v2mGeALSc2ca+gvissH+TwwhCeWVvw29ouuj6KU/QT
kQigeW6C/aXRz6fUKm3NoPMT7BbEIpkUoOji6ZIWCwJIlyO6ks2Rz919ltPCwQlS
k8Q+0KoxN0r1D5JWUy43pGvn3cnrNfGRUBniHsyTPSInXysPyHpUmib2yfLJtE9q
1zxXYgxU4JNDUTDa4APLUEqy9wLG/4tgXZKaKJWIYAPMqVWFx5wl/C2qjvYq+DFh
BinjO740xStB7XGwahQd+Y1zztbNfiDCd6ZeMPjvJq7LEFWqw0jxKBOR0u4DvXCJ
b9HIWMfVODUv6Kbtlf5pFxmXJmbGOb5s52kW63vCBZQAG0y6QBq7eToMqjcn16Bu
H1TCT42H6mY93SDSYXnYsls2/uSKaj8F76l4Ka7wrWOqFDlffHe96sW3hLDr0mRz
4Mn1/ryaNAmpyJita1G4HlqzqWg68xt25abK+ZGsGhu8sPkDxGJvaqqwe8SXYcZG
hmSO8mMM6/fwPC0Zl8fL+wtNYFuwMG0w7UlCbaq/cETr/qv96xVg5cCTAKVohxG1
fEhYjEhLvYQeEql4PPmnOmkjY+2p1PY+G37R+tWm9Kd8gwn/CXGH6MAi53zKtDJV
pl60iPw3SOFvndn26DI6yQxZ+1eLHOOojdE76tMYRMRIY/iiH9uYinXS7J4e/vFY
BdDG/2dOzO0PX7+9LdT6jpjiB5jmoHLD6Hy6T7HB1dDvO/YecPoRs2ZNy/DoRI28
gKlQq2D54XkIKCP9OIauxn0WfYdpokdzceOTs+4MaJaEEUk3f6moDbw+Gey37pr/
iWkz47/sYcM5SJt9WXhS74EgXK/f0y6AMnNm0XDbW43K22AxaGyb5qW8D85FubDX
u/IW+y9xXDap/ZHyTfD4oXkQeuWDKiaeTB+6vx88ceiRLe44JrBMNqTI82SLlAAA
T6+P+Rwk5UqQWDkYNH5zkguQBo1H81LtJWoqTh5pYiTX2BdLdneStiujNGUrF5cy
Urd+58tgF94bgOg4lmKA7JDF9P0M0mJ12UsiO1T1FbPsAVGEPUXdu8N5ODb3unic
7/jdIX6q/paImE7c/jqgN0xwx5mDqz7w6jyCfT+6mYGFhMKZbLZiTHXKFQRQE4fA
iBKCmEKCH0md4rQsmztm+6I7EdjhvsQBMSJ/hPDdzY0qt9Z3IN5xBPtk8q1Zc0XS
UnQxCN/68xzuO1Fvo6ifevjNfu/dkvrdSIjzGffHFpJ3RTsb/gHXe4i39Sbdssxl
IFrryq7dx4EbrdiO8CE1ayHtBdiBAyXV7JndGfeIAPyt1QW5bXBllEkapPBgWTug
6qMQInsUvEiXqRLeOkWHJHUmDrr6c0jwGisgr1JmUYGYPL2eOuribTUa27PP8fKn
W0OYI3SwfqRCYVaIthbcMa06stHWjvcQ/DV1oe8qzEWIeexn64Wvs98M+r4XE5cz
DBbEWgtfqHtjv2SWeWRNY9BIdMQjXr03cKHC1+Oore7YR1PxgOgYhoGS2AlK60Tc
8eOfPuO49h6fhouTBK9qF3RUuHazer0ogeA+ILWlrOsIlRBnZp2FMB1i9KQcfZGa
hAnTGoR5HdISI21DQLnoZBtxeWak8KssaiL1kUftVxpqdO/6x8DPWY0wD/gB4fE0
BvUZ6Hpb/WYy0l1X+MH8dif/cLDCTaW8N2TDbQqgA5JtGOfKszme5tph+s0Mqor0
v7rdQAZOWueZ60p3783/EJ4lTMw0J5UruNQeH5GWSVhQfz3q8W2EKpjGQLiwZlNy
Y2dQgxaLaaVJmR7xV01KBFbB5A9Q7ukUcXi+iVO5znE86Wy9nE+rfVZav3BTKwbF
6dg3mCZ+jvyS5Een4u2lEhLIiRaTzqoaF9mURdea+j2aTDkWpb1M2F1hXZj+Kl0h
ByPme3LKSGIah2kNkZdHe5I5zQNrbxGg2yLJJMEFJl4xWTIah4LiLx5WGAZuQVUA
uMOk8Mya//mnDZcI49W8GmTGE8hNppIYgn/O5VUcqexFfdDEK7ktNqGnpHnotqbv
6uPRmZ2Ai9wtTeuVnXa9Oy/9Od4Jmg8oFa+9eK3DlDLp90mXLrGbtm3Mr+CD4Eb4
Xf/rcFLBxBUSPu8b6MvnH1vla9gz9KcPVf+sOQ0ZPdoAYF3rrQ+rz9A0szJFgzqv
G1uJsk0Lg9gAPRn7bICBseFnVMJJFxdaOcATh3CKCjLWR1PIkHf6aaZbM9IPidFC
+v3GYb4VTPgVzk4rRO0AyGA7UDl7DODayaBAcz0hrZ1JNCHLNkzwXJj+XCncS6HA
j0FaJl129tqpnivhHiwsA1ZS2+Vz5NsNaSx816mrOmI0DtOKInAsOYzVkJ11SOcl
EcC8und+8SaDCcqDhdn4H+90KmKr0989a2lM9dLfMABmy193efdlvPIKq2Q/QLKA
z9bDu89vf33fkER4L7z2aogH3wjfCT9Ne1iDUbF04Aa9QP8ys3rMX+21K9W9kjgY
uA/p0niX0kYfvfegRCTIXT+IZ3D9362ewGVMTQ++P/9Shg4dodUrfx4Eq4IPG3Fy
uQhzTdBESANtqvhplpLvYebxgF4vEgQ7/CccdgdTMlok2B9YUdkoQRUYZlASR4vB
IrBaYeAdYIXMPr/IQmyH6aJEP4OWVjkKOvUpsBXwu4sFyQSjrOmyKX6YwYFNyX9c
HJk9rkn1JuW3QT8mVLLPe+3az+jgqBLal/wNTFsvtqMAn0LvWP8F/ca1LzCRx5Ck
XzNq25sJSe+2/P3bsoiittALuZjb8+ULxMXBtQfQMehimoeu98J0UHSAPy8us6oE
PFs/IahMencvJIpqPJ86L6gCua1x7CjHjjnOUvM4Td0IUCU/UnKOqwN6EZ7SZUbF
joAEEPbyfLMKzqZZCMnpLTkl1xRJQNPHKQttcCx9UaqyyTtAa7abuf67tekjw2rL
y0s6d9wEP9+XfDSfPetNcJmRNHoIgx7onhRGH7BMeYdbgbQzgDA0t+v4+I8IV3fm
yqE8YmNYzCm1GUvLTQsDMzt9YyKyupnR1Yj6KkyaD4F5NG2lzkPTiqPIEQh7i1i6
QtZk5fn4GEgI6+bPcN93tKeqY5fV3BAn/h/qr/2ROhbGiCYL1hiXphojrk+yRkJm
gaPaFL766BqTuJOvMqKVDxFOXc8VHuaxe+zJ38zyqvbxhGxLi/UL0iBXMtfdrsiC
SIRezImYTrQDyBU0rS3Qs07Hjye3+YjbLHE3pIOYSyu2QJBsV9m4cIqRSmdqV7iW
5PDcbSr+rfGIWtN39/oBq8bcXw96GaX/wGWs9pZVEL5XKsjgeIniEScfNNC0+ngD
fLe12x78CSJm0o6F2UnhmJ+2VdWJ7jfFGx238GLQooRHPKQgi2lwkRZYHVOtqrlC
w35Uw8ynISORQuXVYndMmZgEuvQxqoD+fN5GGh6QQa9y8H1fBkh3GfVHTccV2Cuc
YP+80GdO5O+eieDcjtk9A95XY5zjt7hDQa0/DqWZDh603LsGnpYxW9faFvfnMP8K
hdmyXDiPaGqVru4L9ct5JqYvMK6dGGZUTRC0JNF0NJozAo9PKtTn+e5Vn0FE0GQT
9vDKkbKEiIH1e2j2/VO/wEyxQJtlhjbDdc2IsAWBjiaA2FHNghkhvxsVX7F6nbn+
pI0UnoOVgPBj/51RWc5AE4AsJj4jDoNjMDb8Fkd968uWLUajjK5JW1SH3Ls0FqsD
3WjzjuvpKY4sPF9t4jzGWA8+ifM1sKZ67oF9syHcmahK/E7hJl20wc10n6dTSe6j
jKMLS+vJWJjhPvKsTiZPFg/abs1Ir/MBv/MvTYsM6M8RO0gUUyEXhHOKwUCaLWhT
+TSgUG4/J4pFi7hTjN7OHZt1VuBsIf58+oLRbCguCDanSnsdRcvhyPVx6sbx9H4E
g1T53TvS0lo2RKz84r0wwIrDrGMEd6iwB16cDTmW/nyS/4aKQ6GpnkX917VM3SyN
xkZ8AtIXth68wXBzrkBZdEoQ5bCBJYbm9SCHnh7a4NsEfKKDCCrP8zQSbx8yPpDd
2R+WzWJxZAxZlbk/TQI5HaI+OTsrAoJVZEC9xQZ7fgz80RqTdNWozl2xJI9Sqw5Z
AopxLJJ1yOBO2CV8YtrUWuHFAsP4FJi1lfKR3GlhLtBcIXOI3SX8UhbxCeZsdA6+
pp/G+JoUfEijiKMfowT0cvtA3pqdJSBcV/2gzLc73g4f/nLQaQPaFY9JDKYDL7cW
2ch3uB+5oAX5swKMnZraq/gCrdERogwoH4F2SgaQLkqr7FGO235QmrsGVFA1gC7M
C1Yg4wcv3VbqQLEV1+4itrx2SwicnQR0W+ZpF/uO0YgL9hFa9kNH0XolGgCIjIAv
npYiI9EcfZDUFicjIoH8R67ILKnIKd5hx814LreDfnic8EbpiYn5xv6DGM7mddtE
PGoL3gvIYzsJfgooSAHl0il3R9ztQZ8qpKP4GVmDHhKJy2bpklW6fGCdBxpj+00Q
n8hbNkmZ4LCIjiqOsI6EOjMIgIFK4kmEikqXl+wpbdlmJligz4qGxiE+Mw3ZyLtg
16jTzCF5bKBIDkbEd2GL7f49a35F6lAWtp+RGbgU3P6vbEssvMcNn0pBZElMPuzO
5cJBgbZWsrQFsMz4UJ6AA8T1Kg+ojJ59YwEo6b4bnX+xRCO72vI0rDkHBqtM1vEa
f4VzEP/ULyexZY0+YTGnAyNGVRm4UPM6a754bbtyHomlPQF6O6T/8jme369biZ4f
ive/CGo1W2abdQWRFWd5LbLBibRJQrsSoJwQeXg6eBAankSx12oe1QFx2Br6S4jT
rP98tGk1gHGeTR89K/OiLD2qo+9tR39qM0HeOecBllHWldc676ItUdqx5cWyLDYP
sxyqzuAgBCdmkU0ZQDIOOTPAU/ZYo9kdnY0ZvPq72uRPMW0v6nivs+YXpgWb58nE
+Q1/YtGJwvDUF9bYdZsQMafbBrSTRaIKVQdRIrcP5rhRQV/wOtfZ/ZZ3Vy/lTQMJ
CXQS1oD8XrBa841RMcTrF/zhtsmbCcKN+HL64RRrUlnpbnbVbf3+8z9lnkftCKq6
1o67AIw7yjiL/Ho3qkJ2n+hVd94Bgn83Gqxz0IbiK5cITSfMJVu6ZTLncQfG1Zs9
3OIPpFNgicICLJUKidHU/LMOPIWQgFTGIPACxHq9WLXzXgxfbPBv04VJBxPkksdT
WsrMNBkF2iGqOXTFN3dS7gxfgNWCm/R+TL/zgQNrqWeX0wxECe8cjKLczpArFXaI
v2UbEfXONyUPFAfoPJF77VA8bBHbXTlJw6CjHRaEVd20siNRxZhlWbQohXIc6qzv
ZP+jIb83iwbTixhhlUad2PaMbKixVQCF7AYhhOMQLE5UttK6dr9lfTC1Xjx7tEhg
ONr4oGZ0rxqj3P5jJLyFWfghi3Ik3FfCrrBHxJ5W4amBU73bZIZBp8it2KDS5Ojy
zRncura7eEvCzce4+00RHC2A1eQwYemgUQhLL7+R1B5siEl7s1nUSefurFiTZ7c7
W5zHuFtSd2FTnzuMxZNpngyQkpWAP77wh4RkGuwUJp5ix6+N8Sudh8ar9C4i9TzZ
pYxHrImroX56jrVzz9mLg08ZuXw+QSvdH3BOjnDyA9BOw7tz8bQvdU9PeWMjfzpF
exQGe8nXuCnGZsH/NQGRv0YBAYkdlczs6VYcscgPOdqgnxAET1JWKlwqXyW89MDH
sRaSe8BRtdHHunpknXuqpWAB1YAmpBsx96NVcTXCJzR5rcWBBkDMTf14UsiSj+WF
MqoLf8hIPrTjqsqrZs5z4//86gSpLT70DR1Rfe7dL+pHstyt8K3iEAUSp4HuEgLz
AIXAC1IYs3bvW8hfEo5BNgzseC2Sm4XVSlnXWdgZU/JxZajT0q539LHTmIJuC/P/
2I1VQww6PMuBkWIPUH2v5Auy3p+VYApQOssph0bDJoG0HaMNR1CKh5sJeqQRjubu
1R34cEWo7N2nTOXg9UssZu9kijAPN2K6Dqwf6HvBjZqclNeMG4C8BA+Bpvha/Yon
gJ7w4GeF+eXCyw+teI6nPRoBptnnBdMVqRubrGhhGIL36+eBxVDaYLSpP8VRHTUT
oX0bnVFHOz2GgNS0ifNEIzNo1DCJJfJ72WbHr3wtsJfSHPRvLXu6w4gRaUl/rzjY
BdudFbsq1wwNdirAFeaO8zzLWlD92vGyxjQXq1L2kZtXNIAdwYr+i/ytzAwFxUJM
S/5WvLX9R096g7ujmLUtA55CsRAz9RodmHYKAwz6qQzLCuT7csEDojrHOpD+2QU/
bzop71YYtdSjSYdZXn/LzphQYS1iDRe1XyYGF+MP2glo/6yOt4sES6lfZ0fLRptt
vdj0kX1H5mLRA6rmZdGgMGaQBhJyojrSNGK8mKbdrPFH86QQMN0VaXdaYricjfYa
2Rq1C47LUcToUzxtbyvqvHqlFXouA9DD1Snp8YydsmR8/qD/FwJ3ntruY3WqduEj
GZ37ZDPb6hU91GUwYerHJFvyVF8xEashAaEh3guAlKqJq71ovNPDG85kLrra9wrx
d2PID2+x1GsRruStHW4g2uYqDm4GzaS9foIuPTRYnrnXz+OQBKAwv4FKim+fVEOX
GBgUboJOvsSeMGoyiOCPWMghidW3dj40BfG6kZ3tWhPHEwmAzX/59A+RWG5YILec
BdZwFhHL3ML9jl/yUy6DRNEdNZr4tNuYTyUjbG1QOeWfMGGQu6G0ABJo5dnYL4w8
RpdpWxKvYKQc4vHlx9aKIDjd4Op7ryO7nAHp7G4cUj08WHzopPKYMzZ9TUbug+to
mPQvlhfYltzwBo3v5v0FX8w4mP4gub4GCo8Xm460eUUYDbEo8ldZ7r51HIZN8rYg
Yhg23K/QZYH2pVCdzZ4FcgrPy4O5Yy1eNlvqQqK6IUl0oLDDt1QCJjZmhR/0OTS1
ucH8Hna6IvZCl9Lmgbe7IVI8cjilXXlzaiJo9nrCwjAF9/3a/a0u3nj5UOu1U0gu
6IQpcfZy5lys+6dyA4f/p//px/liIPpgpxg7nUmWuE/eyRg8D3ZD+gKiIwyc/jLU
NryF/vIwdEGRBb/NET6fUPcFj9IwxX5UfdzgX3kFGqfmajS4TcAmRdmE8g+OdTDh
C217ZIKk9ORkNgC8/BRwNrpbIJcEaMg1gIo9mq9j7oF2c8qRS0gYyHUb5TkE1bvP
KSRiXTjpsX+UcfmytQdlQKBz+lEpEL4WHhQEo1Xi7FkP3KCn5yccLDjOS38jCoUH
2auu7bSWu44+qLWp6j3kyvTZwUXA0Ha3umNiWqwvW2fM/flF+YOqk5laO92S0FNs
46iiJgVAg3ZzTTQmDaR3ZmaMs5YhMZRchzwh5cFJRBZd/t/x/4rskgPDnWhhWVcA
r3ZoE27YsjE3wXCFaXoXkT+i7EbXJwdLfaGtHsODr17o6uuCBzqh2773N3Z4N9Qs
5JnpFBCGoBfaEyYlNeRQjc9Xmna5k5VjmQ0qn90s5g+avv4ezBWDyXqGEjvo8Kxd
Gs9IfUnpoAo42acMSS4EcdZ+a2n/ZOubfoM94dGGJ+bQw5ys/F0GH+K9ES4cNSYO
vQG7eynspgx79ipZpOJwGmpFwcE4RJlrvQXZMSufcos4cMEF3b3MFcjcFl8P7Oq2
fARNC+HbPt5hkDux5jqXOXkgUJDBFgZEBZ7M/d3kkxOcq3UrQkZTH04uk9KNlucW
u/YaFxV+LhrFkZcAvHjz86ePQn2vMStrFqzxIvc4OUafVuSArjV/2V0K2H9S5KBg
C4YXPblTFpiC3PldXamlCi7TetiXIFYq4RgMCylMOz/q8WKMFy/OeyGI+KTUqqsz
cn5TUDZjinYih5eV4DUx2SBKfRiaCDMqOSk+A3r08YNpxm63DtOYkqXuVv9tsHBh
4Gvs709TLYfF1yFkYo58ewP6d+EjrfPCQtgCtFLOxQKGPOOX8+eRoV7hfchZ+tMU
mtKE+rLAhWgPJ71hiKYMubs5izTkIV8VWvMOWNmrzRqoE37wO2HDrtwZGlaQnYH4
XXz0TPcP1yx82Mnm87PzNp1hbky4tigtzyHY7KRXiRnlbW/Gv0b9fd/1fLKk4mLt
hof+OlR7vcywz6U+lDCsC8T/yuYwNWmAYgsfxccuQ9CsyOuxVWWhn+v5P6reMNPP
CCZ/jAXPP52T/FOc8jGgucbJwV9vwJMdWYB+xfL/1mgN5eEBQWspA0EAzVFbwWBO
49Va1m5qmAEk5jdwwZ1YdX8DFKJIVSpyQDfTmmFL+QfgO6v1uQgGQFsjRcHdb9Ow
sWKWCECdADF7+sWTxR3KBQ7JNCWLE4KAt0VDhD+fpCu+xnKX/X0nHCD8ddvXp47T
ZaDKtV/P5b8r4uQZRp0jrLyZR/LYlIe3SnhRmmuYNhN3a3MughaZqChTDfjhsU6l
Nnmn5/X3dTc9YVFYs3kocSpHoBIXBaqySJs+whetArCbvlMAev19HANUwNB2JlPI
0tkr+8VceaRmVUCnYqllkpLgWCisRF+RSbRwAkx9lIRlw8zulhOhajPlu1GP1UyU
+CYBfxEwpM1iYHDe4YAptlZHRa8jS5Qp9ow+tXfuxLISd0SvXsyVfPG6WreU7EGZ
KQDIXHwlGVXds+mpzsy5zLjhGtaUIw1kUvJ9SXGOWLstIQYdbERPLBgtPi71usni
GAVXX9j0DKWz4q++7g2aZBt3YnNRHW+bnZqlmrCaDogwQSX5QOtO+fQaJ5ely7fu
l+gJ6E+IOcvPeXJbLCw36rbfB3JziloVSe7fnLJNIhifd7lb6m3TvBt+dn8/Kdnl
d02YSIWm+GYM7SiBk6Dw67gfVEIa7D/rejIfGEkrSTxm3fT1VINNbsCatatVwH8d
CJZLLTPsaJZi7/C1EkFJl0bF1J2nurDfuUbjg8kHmvG2KMZZGRn8afc+xUKwIqbT
QC/mxe6n3HmN1BRJVfoJ1S14nJ+ALbumH33E5CI1MLJF5TTSmbsnWJj9eGkmxMdZ
uqh55jqhoMfu5IXVAcTB5R5Smg+Ho8S15o4jEdmNkkpDU/b9iNJWvyy6xkPqlXmV
FKswxP1TqNs/9J0EgZl2R0RKbKWKsIPhpAczQhG1IAhO3QQTHlkR0W8+m1u+hZfT
6eYOGNI/zjGI02FYEjkGn9FQEGa8E7oBospHPMLr4wEK3K8nkRnx9b7D7FQ48tI+
sCN4GAMCnfkPMWFEUm+MJCZvWlEaDmhm5JMbTyBhuY8vY6wB4Y2UkPx03B1PXMav
MmTZo6ZiU+4TW+gSJ9ggpkmS3WT4NeeapS1CeWVGReCA5dTK4FPBRSc7HzQ+coib
kbDZqFR5ClGDnBEV30Z9/F4NNI33IpcWk94Qbqyn1nnPnKFX+xIVZLUL0qqiZ2nP
0zCT+J0/YEAdArtm5MOzLAco0XUsMChKbherO4vL612ridF86dwVFuAVtG9VzFVo
3Cf68tssQI63nMUBbGzvacv8py2Tp27RhhbVRO/GKjK4SEHNc6A4z6M05Q9udzmR
DjSI1rkWskQWX7W82gO2wYiLxCH0vqe4m6U277QuUEInQTGGNqe7pKuKuGFeKxl4
x4N3DE4J+Sj4vExUiImbhCgO312xn8TILCEGegxJA8/pZ2szEu4m2MB4yrFFKJE5
rgiVGcpg7cGF5IHq0u5euG1gDLzB/3yOslyKlk9vzTOgiRMMuN3Wh9X+fIbRCcGu
pAAxAb3U7GcHcgal7IIyU8NFAjDHByD6cEykTKiAuDxbPe2pfHPH4Q3PX+zVjcIJ
Bc7jqC0LJMIxG/mGeAj8tUJeyzL9QQYyhg+9twXfZGQR9sRhPo6CKvZMtDpf4a/l
okdGPKG6A8Jzvg1/AVH72NeDb5VQoiNmbAhP8wSjpHKi2/ONNNZIhV/W7qUNPust
ugQBmj4YuoGvXsoEhNqBt4/EFphLmGPg1aM26ckW/8nLgV+jaK6sIte4UmduRfHH
hu8UZpsgqGOoPk4lA/J7bak2d6J2inwiwJ3RORHmwetCNFugiLc56LjGzDAUU0OP
b5CO0liNrR43bT5YUAbehTK0oNC549Qt6kegCu1mxAZi8OXTrBsJIAfRscqkD+J4
tl2rLkLJI330gu5I1t6tK8IrCWZBZpZn8KyZCICB9kHZevSHvZBzqiGycj7AWQWY
/3l4yim+usvrGOqy3ecU2MXhPIP1VoCC8iZOp0hPgzxwVM970AXl3TB/7xbnybht
PeOuGFdHeVtCCzbbGtgKQlWTXUpxlVpMzKM3QcsdMMBwF8S8jNy+IuyXelDVkyly
ItRA5FwB+TBPzhoB8hVlZ34TeTkl/4OLH5M2+Ndj7esIXVIRdVP8pefM7Ph4PJFw
SIeYsxymIHDGtRPRwI9v6jv01lmb2gp5ZlUYRGWUOCnMvBOxocbOXSQjYCV/SdLW
bbkRjqeGlTSHgEQ4TNKrs0RrUWEGwov8wAkfFNDrf36d2yY0QlG2IesIPX1MNgoM
ACyLigUxYdAkyOCdzHJiivMYYx0m5Rf91eavGM8hXLyIMYD6rHGNsAl+mwoM4+Dc
GOzsmFSTA7aByIEVI/L7ML2TrOqIbfxe8IwWpHio5w1UgK2U3qkOH+Q8edEDgvbQ
i7ggTyiZCJohyiiAMOETLOPocIs0XqV6VIy68Xua4Rv7rhg/XzVCeqcyZE6Sjk0t
KqGCmzOU0fFDb4J3hlZbqIJ6Tdo2t5AX3h9BrPqiM9Z5rQ5skqrV/hlhD9A1gNEO
n1/rxh138NCQzTBXrQS4iKthYQQ0LeryEW5pZM6YmdB9s3RaMfd24+78Tinx+bKU
bNFe9WT3XyPkMruBvNMt56SOrZA9UQX5M9TDqVqngEFSlJqqsc81AHYViZPBEeXl
4hLSrPGc9hsKsW5yFK9marhQtC1Ld4vEOEfi/8hcqQ1eXcqcDRuyNbqiww1evuUw
hlukSSXyLdyPYcy32mfWyUVpTbpvTiG1HyUzYnw2QDgYeZ/CHeMx+7S1rtKJZKpd
yzdF2TSLRke12zR0NlmkhHM6ZN5J1ki6dHpPSagfW3aL1YGcuzL5jtSjg9LWciEA
q6Wks1/UTuza6uAUEl/Penu4Cr/pWH8BPSlrHcIYJCL953mTzLa0HrkJxuHeCaxD
RnT2R8tKDLm9kqMszAuOCbZw1l0783g8DbBhs28A2SNKQG04cQVnF+s8pMJ0OxcS
vPHrGaFfFAar0LzkZreNj7ZJpohPli4sSHA740rkKFQqEA+4dVRD2Fz+oLiSoqli
6KNB/JyvwbxIjX4POKWF/IiQk4MlKvSfINs6EUX5B7rGH5nkFGkzcF3uWuJjwP+i
jzhovubwoKRt1+DPYkvzm2HrF8uXHPsjPSj91eXeyFpKBP1Us2MGayteuHSF89sv
d/LptwAa0SZ9hJ21YDbRX42+R36ctBDxI3TRnyyrTtzGHdSU/BzsFrxank02WVro
Q+OeolJK1FEa1fCgJkF5C557BsX33vXw/hAd5nz6o2+jpJNAnoghVxg4hwYSfKem
QB7wWGGDhsaEBI+rcEvwWa4ydsYHUz2c6jv5C7MHrkhmQ+vNK2uxHcMoBEA9UakQ
XUuSjGt+Vmc3ACZQBRacdVP8d8+Opz1ksfi0+5hIWLWDxA/EzpbhhCKwuukGlnow
uXEmm8O40AoOu4KYto+NB0PBnS2fAP9ljzAvucgDy2QJq/hn/gMWrsc87NSQGoma
ysBIYA+D8yUfhFuoiT159bD9QLNyf29Y+DH7RXI8iX13DL4wbICzzyofTaqT1Ax8
gnbiuXoKIKIE+UZcpS/zAIl3nQUHCf5/XqH2kp/aCbtVYrUTB3Ys3/plhi1NBoW0
vZ4fz2du4ZvPepMZczQzkFApDDX/P17iD+NGfDfVmNtXHidJm3P2dtyxBYYZNd/+
LILZ7sCvLIhl/4tSaFiVkGvltEqAYrnqzB1jQfPx0qess10C8RBGvLJDIpfiZTrE
AtEINgGvhWjcCinzsM0Q7Sk9i5PwUOkIWmyok+15HR+YYIe3IyZcARWKeZ26NmKk
3tSiT3idh7sZT4uUWoMy0wIFPcM0BM5tvOQXaj3zPDjdaduwrC1yVnH+xFw93jgz
DN9J8agIQ3/U32t0Irp8nb2yW4rrsHTCw+4llC2VwY0heG6xC+b5143/4n/2hVqr
rjMdIbaQPa2x9GT0Je5Nks2FmpbVu00MVU7g/aA073ew2ydpQhgJon9bTfo6KAHK
WaxCLgJr1GnxjISuPW9cgZwyHtzvg73aLnfpVxalOV//WkYBfc1iIRdc5Nnnv+Ja
dJz02sMSbp6ENwUUAlfEQMiRHT0HjgsOhuTrh1bmhMSfnv5859rfMGCsRVVG1ejm
zS9IES7TkVppPqh3YwZsnyk1+xUhkjjUdXvBkBeUM4cHKmO3M5CWi5dzJ+R3FqiK
WuGS1evVUete+Rfgz331Fb+n9CMbRyb66xFmSm0bCwnHt+Sk/NodvVTSeiarOs+a
cFO367Gq3EEOw9bgAackB1fdnG6pwb9J7ooL9l/JwWvdo0ehhFePm3b14Fwxlxju
r0WX6Xyd1FrBrqvfYH7Ifp4RuIqciIKfIErzaIpyZWNaoj3aDWiV7S5YIuEIU0AP
cnvxhDL3l04FDeFBIARo8FRKB1M+1lA3wnmsUnKBM7IwU50o09AfpY4TmXECNGdG
+WVbqD+QcgHY8sbPEjSC+8D0RYbzR8h4I31ZC2rMYQb2JK5KHoVFckhtjScQylY9
hCWbZfYYjjfP3ULTX0RIEP6F0tU7DjBUO75VJdKjjGiYuLVD9aW5ILD2UeU4mJvB
KNuIqF87BDgSILdf+jalH7BTsFN3DFbMizPlsC8oTUkH55UOLPdn6qFZF53Rixcw
eMhfbDOQXZjQ05ktNm5ilIzVMOJL6i1GSHfjUUM6Uwd+1BCysx5UfFT4C2d7qglT
xyUIUOKj1kF4l4A74lFCrerGNOJXl4zxxorp9ISB219dVhAZzLx9QPOkXBWaTKmp
PYVsc6NtI7Wnbggn4xZUWIe8TQ4tAXIeXs9jSUKl7/IodXme5EEPevls2yNuOsU/
nAhSrPHxXuPLPinJfp3lEsELVi/2sPzTo2t7oSPOEpwE1wg7wiotHIacShiXlEZL
jZjdb8XrW03Z3t6VfJ4hLZWEHrgaM2pgPqF2fCi0JTcUrF2MVHL8jWWznnLxF0y8
nDB058cEXl7NMVou/2BsSWZgUwZ6hO3WP7AHqYKCWbrCI7pU6Jozjca+QLXWH6oY
JXSfVBy3V4hy8QAosum8vqWwqenoNsCnWQ/3QEGSm1TT+9DStH18Q2okql/oycNP
ABmFTn6zbAdUpTdm+lCXhTuq1HlQdNU+gamPQKzGNASsITzJ1l4jVg26xU0rytGN
dBZ952ZZiGEczIV9RgImPvv8RJOU+Mgggb8dFNFy0BfZLqdJitptoawMZUEYSEn4
4Qc3m1hI+ls50DL9CwkjbzCNZ/POvNENPVCipM7ryLuSpaXZacZp7hvSSfqnrH0R
Ue0iInkka6pDcjh1dzo6oLm8QxstN+PNs5s8cGKe8i5Ap7S0zFPBismx95ri3YOs
VKTbC8QVdfUMMEOquDWjPWUGDBcl3qdJkqMx3opTQ/t//jQSUeqeajkUJ3rjhbUf
1yCoylRwFKv2pS7lgO2wDUXdDPpkzdEyn9OG38n9bzNaOyyY+Ez+OcUCALHy/lYA
7Bi4utgGlC6mHQ/ryNcoo+G2XMsbBoMBQ2GP+S+RdejMD1NCVsvVJh2FfpZ3u3xR
pHHBTZ0qmlCROQOR5Kcj0X7cK8Bfa+3ighnF83e0Q+1gxAec6k6jMRth2e85NABG
guXKeNJ2DKWF4GAf38Rm2L2Gh8zkVoV9iaG6FiT2K9jgkqyOMGVs5pn7oyf8/K0C
3CcMlYIOIePYy3p/O98KsfzWh7V8wWWKWGMXbPE7vlmmjKJz3/T1Hrl/nx9hgkR+
LW8C+1eHSXqTjmetwDmPE033QhjP0aJj0Yw0Oxw5O7xkisvTY6dDQLxN74dLaNZc
qzzAU7mRGQCo4CeUUZNMAUxk7gLuANsOIrPJPfIbdBZYdcV8L7nDDEGUV9vPG4EB
cpFT44GONQetEfzDpcOwaYxbBXC/ocqtZzyTmPfoKo+XgA9bL5HLChADhUtnFg9l
2WZ/c+ynPyfZ5/tnCuhXY29FjxAvzOP+tflaVsLgSVPuE6G4M8PsexjSiD0ySDgK
Ge18+LT1hbcEY7K69bUE1d+5gx6+ohUZUsONqGA9JUZHI/oVWDGCDTR/PK2tFamc
LSZRdrPzgSOzL7lH4ygqxYBh27dBS/aff9QSVlF84KhTpdAgWUrRyLu5Qi4j6lZe
4ctvYLY9+3zrI+2SreaAoXJtBtp6Ss72Kkim1xUMILFFi6QQKIIX4aMJ9hvaI3CI
g2fxASSyEZ66CCWiwPAkndf2XLZgl/1eENAmdbmXkkV0vGQIscRnT8Rihoa3/1OX
J1iCGSCb3VGm/1tVVaZXZ9APy8rwVtLwA85MWlnCmxqkcIxXLfrvdAEx0RAuDF2s
S74EtY2VpSFROonTuAzKe3E4G2XvrSOPytFgWGNEFGiRd0L8sVeeM/aeCDMxskxc
dBM3L0+R6ASyiLQPRx4QBARqVR7xuvIWQGZmqLnHKP2BnpDUxuYEy4+ce19c8tNL
+PI3YtTEM6nK4Rf4VGLs47mSew5cuC+F9qypx1w7xlP5/Sbd/GSPENlE1hiMHGUJ
VZLsUsL34qd9PtxBNiph7vwUU6SuALiX+YvlG/piaV1g1NTdkfM7Eh4rvAWl2bV5
rgCsZg0OXzyicPIRepfT9qoUlg6jzwMQQAZx6+31EMyc4dYejTZ2rzcnbrMaFkg0
nSy7jABq6EyyZEgQJuivJD0qfQtl3o0NEsarwb5gfQT6IxPnaRdiKcSYAfB0xRaR
DnPwBoWiv0o66vCwdwxAl2BvrobdRVHKor1n0XqJyZpUBtZUe8i0tT7dojilNf10
5k55eGRysyVmEYNuz0OwNKsesHaXs98RaoRkzVUf83MxjFuI3cIo+rX846YSBJAi
Anw01xRWJIqfqFgCGAQrqxWxowi0c4nPwkYTqmZYI6sEQvVK0Fvw09Kv2hkHFT+c
ZgmvFPd8b6HdVtPS0hu7Mt+65b8da/3BCoONL5DRT4lOPZrNTyhJfPwuBk8CQCe2
Olr7EuBwij4NwT634H16PT5j+KMtmU65/OdovyXFCgvS+t1pgxADvMi/EF4/C3gZ
18q5vg/uZ9Z5d1V+27tSLJ6NIt4rrGKfn9f9oXUJDX2ewIlR1Vo3OUiRqad7raXq
dvjUBhy6pCNaZYxdVnwgestSdo2Rs1HULd9UGmwexBFjidofOvYvyurp0FXiTQgt
TtHghDcXoII9mX59u7vm55/hWRUOliwBOaFaio+5qLF6Fql/0JOMieIQXaJNX5cP
xeeiTFbVLpafFAVAfdtowqgnV6wS6q6ccndmZr2/DTGz6eA5jZc6bF4psrEK2Xjy
ESCFfpntsQqqVM9FRC0pycaCWCQ7jDAfW94CQhoTWUrp4iAnj1rSkp8QynAgyim9
GG8O9iqJJ2m8z0Py67FFSGG9i7mlBRHLkzi4R9DDkMkzR4r9fSG+LP2dCjgZ8HzN
rVI1fen4UCBYUwtVuVNOAj3TpXpLtv2vHwS8SVSWmUN+Pk2R6OKxTnuDZ71L0i8s
F3WbiXexQG67+1oQKGtF24YSgb+HDw99uVTNigBYN/0yzXauxJDaAzO7q01oo23s
NEURPmxqR87/h3TIDp8NR5XZqJkiXplgphOIJsf/zkicOTownQahbDgz0dN/NzG3
TL9AOpwlHoqvFtT0rUFXT596tMfLgUEgkLYWeFzPqcl2p9rjqrzAQPoXiEQjQf3O
4dtAuTfkfq0IUSti6FidRcLxKyiIAWeP82jSwqFKjuwbbmOGcC0x6BtXl8vtQ25C
Fzsm5zpIjrb1FX//jBIGRqjP7kjM47PjpdekTEgmmjgQxcdNBh2FRhSgKG4a0iLg
uUc3KdhnFflM53cmShawoNRZZOj10IRfuNc+W7Uyp5ZJ1TY/fzcqhtul9SVpd3CC
IToKSprZ5yoOEfw+4xNNqXzIM4xwoJIBF0Qu1g4getMZt99yV74dN0DlfL3/rjxr
yDkMXYJFxS3zbqwjp2b7e3SKWTdq84aQDWgXwJ/aYhCTQvZbkkziyRp3q7FrXVNR
+9B9Gm4bHad+ulUHfwGykCvHe2ddsIk4UleIwQ9Pj18kSqm+Qw/K5PGrG0arNZ4l
lYuvOfOUQlhRylcvRkqUESMEZ9cegh9vkjNWgCi3pgqdof7dkn++8HZCQGcjb3uO
Kp/U/GwqUd4Mhzrv+AqyjAdEShLIc4Frr1CQL7H/0jBsL3GZ8of5OyH0s4z8Zb6h
zYxDOSoARmqNagB569aZHqSDGphbQMwzmnxHhnNANOqauT2yNJ6uSFP+OQ6GvgL4
ozuygsYxWTr3sFqf6887VuJJY5ppYg1oSRXfe1PSQ+Wl5uHVRzz0Y/OuYXsUXeyu
solGvCPatvrDHn9TNmu4e1vBs7QcH/lta/S7XPZQTGzdz0/s+nDNK4ypM/xNmQ0C
rB/wv+jLRdbWUn3LkLcxxrDm6i16E9Y/PoAGsQJDBnTM/3cGQTgI7SXT94j3efCp
93K5dH5n9jKok+KR5tffakf+k+erED37yqYcKQskGmZP0kZDNbO5xtZqhLeuIHcl
E57mLngGCoMGPy3WCiy6lk88N66fEve0dslAyQ+6aBYbJGyHQTSnW6B02Ve8jt07
dl4FHJ40MQIsPsvtNWc2eJDJri4gKMQd8iW/7wQR+FsmkuHdDJAiwgeBVbHa8jcN
r08Y1t0DE+RGlo25oAGSVMlgtw+dRPYvaUSPTD7Vs/nsEHt5xFA4bSqieSEENtEm
tpZ/w+0UXcT8SGSp/kSTzPz/tWvlwancX5XVlFDDbJtJVmJ6SESj53UvEKLHhNYe
dIQ4WqJXssVynpidOgd0GlVB0rskI9BRmnoJPGdrOimu0U6f2TdJKnQkWSDp7yLj
fDVvBq6iD/mM64IraH9bbdpoYvnSPtX/7vZIJfyixAo+S9mEPjkjGLZHGzqv9z9F
hsM55aEWSPnL/FHegJlPdEg5zdyFLfzqWLaJOA8RJbz0Ir9jfx2LIJa89jvk+C37
QFRv+RApV+WjatP3LOmQUT4bQMi4N+dq7pIUdBH2w50uQJCA+JFdno0bb1b/krX2
Kfqqd94vKcD1VSoWM0uQCwZGJSzjsI5tRiFfWNN/Ng3JBxrLm3fUIe4sIOVrvTB8
XItW3SHooEk4RGRRp2fCXHqjJOgQKB6NxZlNiWKZxqCJLPlmKShYJ57OvjRt6Fiz
kix/X6tqIDUWS3PS4uKqK3kTnQRYWDMQ9fVBH8lp+s/e5WNUEu+NXeqHveNjeYWv
J8OmMm5rGvvPa/1VTlyGkWIizLl4nk7dw2rYAGK7RbK40v6VDWF9uyk0cs7XS8m/
nMuqZiaL9Ceo2RdEPvUukmpo9UU6SfkaO6FoZDLpxsg52Q+hzAdfCB6MGGy7J+V0
z12+KX5p/qfuN2/Ne70cvmQPRRRrUl6Lc26vJ5C69raGah7eaW+Ru4BG/g7dCqa+
qkjQNVQ4VJ/kjBLrteK4K0CM+99G+UofShOaeLuqD3/sXZAH5MI6xeSSYC6Fc0tr
daFM90GMlu2EIC79bCcm/4sjI5d9vz/T3NAazeVnYeo755QSpA+G16CSeEwWy+Rk
xc0byLgqxU0Y5CSGQQ835LVHrfnu48W65OHC9SxPtzJfxpchek0t7go1S+AyEN2X
2RDGRZSnFQVA08yjt2gRfbUDknKYiqiM31zo0NvnnfM3fjKpZpcllGjk3qguttBI
9kNO6Pv+jDwXvMQTBAUdmDQLnAdeVMPC77dVproM5jWlvtfnnSn6+eS6ZTTD+5Ie
lP2hGo5uF0t8yjQOe4cBKny0SuRKvdN0T9IgSzDqoCny9O2GBh3UC3TOED7d05oD
4ngoVMhJRpeJnFfXv26z0ZXoAsyjH3RLTzSjOkJnS/66i0T9pdbMgMjR3JwLmCdM
Q6aFgCTx5Ae7fVs3iX3uygvL6jV5XMk+iw/N6PvMgTqXEqD0Ab2rykssIrz+bCG2
QKKMAmvj1Ec1PIyIkNoPAA2bDhTRzf92xtcCpzHoBna536bXp59ZUa0TeE4f3wFF
7ScBRrD4qb/NJzTsUg7C5Z7u6eefQvifiMBC3v9tJ6Xrz2YkmJgCLsPELrOvfuA4
H4H6ZACm5XxiqJI49vi0d5tmLxij8RtjYV44uv/uN5cgKCriVx4YS0DlU7+2ILyk
KYbzKRI7RpMZglNMfAVth0bSRZNoUGXgZzuK92p9fnK1J/HSFbJK41WZDs7TLSK4
l/fZYR+qw1BuGjLgfHV2SX/TWCtAOBuVWC4MYBzDxip0QhjxZFn2tWCUKA9xXrDl
IzOC9hbc5mKaB1CtTQXWwLPN/ZzeX1WzVAFVJRUvQj35FX+QhGBf4qdhrq2DbpcM
2BqmilUehG8vGBbn2t3Kk5XGoIcOMHWzJ4bpd4gg1cs3tywhZcd9VrYitWiGmrKL
WVLodh9fg7Mcuf7l8qCgijpblaMBQhGBwIdX3+PL1DQ2Cpn/hMPoCs8qdyNoFa6r
QoNILWTiYF8eiJaJw2bu7OtzQfuLPBD8i8brfG5ERxCwKDTaua882JJPdCuJe4ZG
AbiA2JlyGrG0CDDwU3utbcV+r8Fb7olTvJ1h0xeEQ5zMxzesQjflVVkVZDyBlYo3
2wN+UOjRQEDh4BqNYfWMomjGU+hvc2EHHjWo87O4inGH8OTZj0TL54BSrSFx/iVC
nWcB1cIiQEPWEnvhLr5+fuVg2qglzmpEoCUtMmzvxSaOljVyDw8HQF8A2tzZn+9J
VIN3nBEDE3f8eMrLv1Md1rHT87lqRxF7PaEvdhyjp4Ww8ORwYgE0FsK4GtnEAZ1n
cz/yGabvd9i5zjlZe15rajsOdLxsICNUbdIKjfNEYa6mn4YbSPpq0bYUE8f0LD6y
Eoj6dl4hLft18lL4YgucPe1b2pKG9sN/q7A1+z/X6/jvxxjnIcZVhV22sDhUnxim
QNMRZbT60r7od0kVH94tdPupZhFSyqgjlWDNWVlo+HzUB4utR29znsGvvIQlc3AR
NhbUAW/Rj69pPZkQWz8Nr7ZieGlfG9Nm2sBsx/fVCxX21ZCFfRKaiafvPQ1tfS+r
go7n+av4X3HPzU0pluH+uP8u3rAWANICnJbRnnyuB1PauSo94kSqGfDehKU/zuYr
EzkIQt2BMglCmYA99DqPnjx7RcRoy4GTiwzjiCiGF0v6LL4bW/pL64+jSrOEgwtI
Sbg9cA9afSkq+CqF/2EuNBZedCPyPCnvDznXPOvJ8r1eNocVAWoe9P+vpM+5TgXZ
1MYJt7PPngCsBsBqUJ73XA2L7+Ea3k+7gWHCwRxGLumrdV/4QfrzrulhsJ+9iDlL
/L6W0NGszGf9IIavgAHZY5u6wvcQgISTHqiLdhrKCt9hRcUG+3kP18qenHDbBhRJ
BynlTx0YfH5CQGk9napPHuvGX5ofmJ2D7pn6LYnlK3YJ4e1ziVsP1DAJoQzQGDPE
EqjSlYSsWIi80llmGoEXnfdOMigAj1f1sdI/938a4wY4jTDR+qM6LB0Wgvhf4alP
i3josdgX4f3q3Wzb8dd40y+zULoBJxHrt/mhjz99FYE8S5Br/8Q506XB2yGoUgWp
cHi1Am2ztuniHbTDChKZdJwumXbONzH9ku6+VlJJUIAlojp2fVUN+3zOOz7be9k4
NhY6T5+FM7LrZ1o/hOeqBrpk2hIJparpRUC83ChdRsJo8+Q3oDjP2IpSME64DumU
aGo1DAD+VlPxIYjRIJGlj5Dohz1+Y52RRw/arIQ1o5JGja1QRJ7Bpt9zShTM11T5
yKSt+mPnt5f5FUTv3iYuWVn8U1mE8y5X2Imo5rfcp3oXySiHT7FEMOS2S8Vawm3i
i/oLzWXAFKhHLpBThJIk2YLsuiIgG0YDXlARoCpQVC58SEf9u5KtrXvXVKY/xn8B
90U4gilcQlQHn6V4QtqDpLoOELWpF606RF8UCf0Da8Gck9kjVud9yDwPbU0czx4f
ZJAlK0+9enQIX5XIxJn+QiXXi/KkNRuVYrO4ZvVB3Iz6XfpN8h1yBtASK/aA5oqK
I4h11N+3z4SWQZqnV8LSr1uRLAQJtuqRbE1S4sCzOT1KiPXyxwTB2t04tPmXD51L
TJBaVCi8FMnXvpcnTx3DjvhbkCLYTLeJHwxhsgrvx2bK/h2rGgih3+tEJ22loV30
PuggxJpAOl519EcOZx/vbjYk5W55H0DoBELl9s5CLOUqt3J8O6h4AIcTD6KzatRo
liTrESuzPHxYtSocDvxrK1Cp8D/XWUPRdpM2UT9oGtCQ17asRMIw06vrorKnGBLs
xICYmHGqclliQvLEEEMJC/ighd2cDt9wClKjdW3SKfIcpRV4me1tKnQKthJxvWD/
rkV4Ugqd7O+/H8iaMdz+U/SD9mH4oZv8Yg9v8EKyI7wJ1/DTeI6x5SjwY5ZD5Aa8
aXy06B7cMm0c3v96ZVOzeKy8idvqdwufArPTDmEa8l4I9EjowTXeS6nEEpzyNzzC
s6y3n2K3Tjcm7kuD+xF6bT+wMAaDYXhXhBJLHdYkEBPDhhVRgCkClSrzXfxCxuJ7
u/1dpE0F27d90NVzNpHXwhh9BQl3r3byGh3WmA/MlJpFB5SA6EBfOkTPZdtxVzix
OaR51cOm3fnYLVyRavCGq/rLGaMZnP5iq8OWDkMoOnEIuBqY8RVvQQmovW3JbOXA
aiRlxE/msW+l6RNmCUjXEtHWw7nPRNl/uBalJ0KohNl40Oe0wLkx2FMynXndQ5aG
nUrbINXXpVYwmlBvHKbGWqEVY5HkzeCOYtEvxxmfgmSdf4WcZ1KyRAPQG78oPwzA
O3kgBU+2RNA5Lhf4g6Ds5pdZeBulwQbrVXYXJqazmvNzZGoxn3kmtmWB4rQfYw8o
HGn0/GcwkWyoRl+0oXX+QhzOBtJdwPsH4KFKXthpUorOiZ7D3EaggCbZbJj4cCIh
mIfIvI+M5JM9Tt87ELZ31Fi58/DKMySRWd/d0JLezRjKdX5xh6kYwBplzrqVKJ80
ZHbUkLT148T1SGAEhlNvzd+q/9lTmRK6jST5G2zBelxLMTIyo0jodf5PMdLIwT/2
4hlcoCs8+Drj05cu7soqZzbVNxIAv8Sg0bwZL2nS9hoVH6GjRrYa1kLCeOQPZugn
RcbuyAY3S0rAuFcrLSqzXH0u9tZ2dfMRks0chfpA2sxohepMYid2Tq2u2YwHODVs
e/ckdHJRRkLP9vy2HpX9rcQqAm/ESrAwOmR1FTEW66QlVp7cf3jfoQN8xs7/lYfq
3WGgIyoBxMqErBRFE1U8UMgv37bQwO6son0n9dZ9oqzHaNtiTzcsUQi1nUwEzFGw
qEMIPI4cPifkinE2PfeUWy0uUW/08pp8l9VSEvYXw8Ii81Z29bhOaYckrzU23+ka
6P4Q2bz+CljCEjOjYD0AIN0+XKZZ3sExyqhxCUSRJvui3aMMz9ZCfWkAQ7VqpXB3
ZDOHXPQUoAcrR/91DPZsIQh3qdp4rKEzuuzzDhPc2/1jIBsOrupKAHDcrwnIxwwG
sJ2yYb+J80/QEqnZlAdF2n6PQ/dOSV+DS9skClt5VgUWlnL/jAGWfnNaIHdmYcZD
ygm0Y2MtzRk8UWEBa2T2pXhHOg1WbL0C7fIuFdXWNHXgbD8svQ6pBwiQRGIVH0xF
T7lNKIh2IYhhemZOInx508Ine4LJyBT3BrpzDq9VKJy4h0UEEf0L8xSG5B1KftU2
+7j8yxwkotf2HKH0KYpdMr14nRGEfQiSRkcR1nagTRF/W8tYH4b8tLoHfgAcPoQB
Z4rkqmrkvA+rf9ymPi+5WeEUgc4OYnFATW+CYUBG3K1vcznZYRR0Wvdf5nk2tJrq
cxpbLkUmmV6/qu5FQmng6niLsogzeIZ2yrev6QYKP1PbUvTnqxX3f+GEICBm7zro
q/l01GlkzwWnhKslPzmVyBiz5Sedp2yMx+TF04VkzLDtr3SRqldC7XGHFV9j1rSZ
Feikwb24Nj1qXvMkBqhObT4C0M7Uh/wIWvKxTq7duAyZdGRob6tneXl11x0bwawe
8I8s3vcqP8WIeFTzxDsvqW9aRYxfRRBREwnBHwVURI7DPLLOrDG4gxYes0qpgKH1
8a9eBCGAjSHOOh8YU/nSx5ndW4fOWZM+YJokHoWaav9pOhefOv78/vbMfIjRVWlO
qZiJ1B4fa3ZhLr2T+uSXMBzoDuxJwDDaHfxnTOt0AgAHELSFmiS7+F3Y3IDzumwb
gatRKfMg9L4hTbbSrebGPl5b30Bi8g13yTHb/G+MY1LZy3mWhyNt9KFSBpJs1r3K
61IrdlVgKGCmfDdFqj4b4YvVF+ENKmB53+tOxcZy/tMucFv4VaHeKq7uzCjIUUHE
gvHqhlPEMSFd6Z40RsmQJeujb1SkOwzax4dbC798rOd9RBmxpHnV436FcaYF5dJq
rXovGC1jLUXxxaZXgb8NYXyJOxmMJsWeF27o6BnTUFOhnqK0zBoxYJnAKXzGPskl
6OspA9+p0PhS6NVjkwHRRbR+aHMOlLalBvAy8YGLd7Hc/unBIp2q0sppTSYl0fMc
mhoihwrVkImft7h8PoVZpSTuMKSpHtSuJM3Ax4298WpR05a+fC1M6EdJTVv1UBNC
PeMI0Aq7n+vwAjWYBHOsZC/1E0dbAaoX63itaQ3++N4TJwl5viPFKT3LOk4iv1qk
V6NhcHN8Sr7VUTf8WTwfLpDyuxo3FKq/IEtNcnK5HWxX4xO0HmLUs2BKvadsRp8R
ln2IaFeHUKPD/NsHVqSe5WMk+tuOgy/0ZKxz2biYvQPeIh5f8V1VIpqR6oLIHFhh
63nH7qrGU5Xk6vZeTndtNMxfUBwUo2NZQhbErs3UAlwe+NXQnJ5RNLAwHR5G4R6M
+xwqYFOea4Gl9QOW5PqubY9pkLZbmTDs77NcQ8NFppMpxF43IFSS3U0QoQs+aLFs
hC4sa9jCu6BaByH2ckcjXsFzwxgmDCivUJpyC0+l39V7LT/wfnmv2T4Gdb+BIznP
xBYkDlLozZH31cbDf7SVQ0PNuqWL+4r8Pk+ovW+lrD/AUSfmxWgvT5ml4NjmnVob
WU3dSr7DBGi4inFfl9c0BuWFaPJ7OYIHR71oGRaJuzE1eEm1v7C9dtN+mNnNxqFL
lvVITpdl4r07iIsByFoExdQbpcH35wf7/PN8Q59SWqS6MKP6YcD52p5DXBIC6FeT
vHx/Wk3iPEK6jVYZvVIbvGEZ1M10BSI9kLo+F55583VAhwSWXkMLKorWyhSESZ9z
Hh+m2zvdDgIHj+UzUyoftizMCryXJ1dTWPtVAwMgsijYKs+8iinD4ncXEk5/NDlh
x8NithVkALjsCDOzikO48BvQQTS4YqDFYeCOJNGCExVQGUGztaVY6m3NkV6xa+tp
bYJ+uRh074KFGBAlSfXXGCCvCf1SHwQ4Xs8NHNNTBpyc+MmgDiSXTklJ0E2/TXWS
Oq1K0siUv+7RpFIpWKF0NYDUu6yUQiy+2U1cIfHKefXxZmf8Xlp+CbUNgV/dO/iZ
htBWkTDdhqmV0+KZSC2EFfpnWuVjaTMsEOXKP9u2an05UXDCeZufSwlqf7lNaAJR
kqr/f+utlcbrjabMVO4IiAoizM08CnZfLmKfVfkW7ML8bSK8knpidILSXOfQz5Tr
R1LgjwgPIid9RtWfbvBGufmwPc0sCCNrA/VGEAJ8UnQpZqt4NHJYmeNpqiBA8rCn
juJeDYBiq5RF+oDvUEDaQ/b+LPOgh6xlUIMqtnEEcJTEGRei6G/TEOe1VnE9Oj1j
eWKY6t1ReEO/Oj9eMkGGPE8CCoI8vBN7LYxAreH3qnrVsTQp2E9tjOUaEbcRB1Ma
KWDO/O+rnQeHywKP+5JtZLQpQk7Uhdq0v3VH1KxDjdOnWUQPjGcKxDZz/DPxpjdG
JrU7yhq/QD0AVUcUD2TmLM1eDsKLFrx+ExmCmdmb2zwW1ULJvnUl+oBFgwunGi2O
mx80imtUgwi1olwfueCvpmVymcv+JfhNPZ7yhidG5ecYETzwzLjZzoa8AbEipXT6
ixP/9LVLEUhZpVurTSJrwFoQ/dNqBvsdCt4+KiLd9qeFNlnESA3XbMQ+l9FP+e21
XOvq+XLa9K5dO06Mlx0lI+M05boo7nqtyw1YHoUbh9sTODBgn3361S1BcW76rJpf
6b/DU/BI6ChGC6RcWVIPNeYaNjHRbz2GPWiho16Ev11J49UBGNUQeWqDC7jGa/33
JOdhOfcVGZ7rTVANPToEkazA/UYfUcMRkSkGk+bK0tnpaQ/M6IGP4MNk31GgY8TG
V1Fwe1QESlV0xNyUzbICqC40T6jodZRh3lhQ9nxMJPeC6JfU1M+9k662Wb1TeAcG
TZzaUqDnP8rDi8ZH16SBH3bO0fraJUy6ZLVKXby9T7XMyypBFicPwmjj1eCQuZCZ
ABrdauzNq2+hSmh33GmppJt3w1Jwu/LesUL0ZgbXhBO9kw5RgIkI1Yvbuq94nzFc
UiRX8gxbewNjvt1YYcuW/R0ddV2ANhktfMUziURHVe07MHKdsrJCPruTcI7MRadg
wMB/EVopd6g4RzVlklpjOD8/3bebjVaaB6RJfTE9xAy8UvsItCtj6OK92V7wSme6
FKRWsJ0O1HH25leHeAVJlpEbd++cNMIDhaj9M3dBIE1oZsVS85mJd0W+flini7sQ
nLCqJq6lm7lL6fVTWJhJ7Khu2+U5RhaTa9yNV0LqsguryUcflqq1GOmxMbzZgCza
7zyvGuBVchLxRlxsY/mevtPu2ySZp8mV8PM7ZnikQXDTGukRaoIdX1u1VwVlNaiX
t8xn8Z612Uq0G74p8axHimWHy4cTCj0McYrCvk50v1iX5eziZ4gl87G3pg8HUovS
t0eFmzAGSSv2cWfDDBoBFgey1ckWqIKSJT6857R+fZ/A40ih4Uq5Ikp8r2O6mp1H
lImaeIoE9DjiIh/Se560HxO20UkpP4RtQI0jBHBtDKo/53HyNdBX68Dv4lnlq0zB
PoGgdbnfpAtSwMtgA6FA0dVK99LEdFu3NtDEL4LM5DdvZ4CmupDc8ziVesfOYcEg
K4TfhEcBHHvZOkCFxW3Ij2XNUss746bhlRiwRTUDKTIdiSDBiRIbl2DahR4FFp5d
HoIRWdJlfAFC11cEYYpJyyL5wHUxytsPD1XFg5iojnPKC1S6ai/6TK/hr4SXh5TR
MFXKN1XulFDNWMOk1/BatBbcTEx+ek+XHh9MlGZum4PLwqV8uuv0q9RRQfo16Dmt
YQPfgevWalMGhtDd9cv7HYOSgmIjVxlYebNfGfSRQtOdkKVCOImoJxUruXOrv8ME
A6B4Iivb45Dg8UIXMl2Fl7mrWaq220qXXoZdJvcwPEAfRBzur1vvhc9XuXTaCPuo
WsJN/kCb09AGZNiLS5jNFKOfJeUEVxmhHUDnGM++LeqbO0QLN3qIMgIGVLyzwM2D
W6YPpW039FBrR58uXOkHVuj+vPDe900R0csFXY9tURC0FPkoZm+KaIujYKyjyxCK
NhGBFuoLiq28LC4ub7pG1WwNVaqmbmC6YZUIAbilovZMszNHInz5u5NIt2qeHJgW
N/DBsqspYw4vA160kWlV+b309IHtK2RKFdjuiuTM+LWnTTNWtZ3TEkwY3Y896SeN
qqgfepJu8I3s4qj/1bbccgDG44AmW/tQAT1JqgbThuW14qbr9yBDPk5rTmpb1nC4
l1eCpGkWhRie6Fdw+gHuZW6z2/kNkmNiq9e9zu/mZz8y29X0mIl7Onezuo5svGj0
oHPy/ymHo0RhPzTFJgyFVBan1Ooz9LVYpcilT2FP7bM1B/FbdERZWBZxk1rsg6WN
6g2z8ef4NIDLldeZx5oJBmvKtPgOWlcNy/fEHWy046NDYOca/D0nl9gA/KsUcizX
SFiIebbxrJyCXe2EweJ0pDCb7/bGu5dxzMKAgLiYm9wYlJRhbeTkNdGu5yPFPY7A
gm8JcE6YdrBPcL58HjTXMQk9r2I153zB2syLbpDyiiRm1gZ4p9VZQjuL8oXCogDA
mp5OxqpCmmmJq988kkD/hXkJ4yTBjyNSs5G2AHJvQ0vScZ7crFUFtpaA13tcYh1k
GlN3OjaowY5mNGVlV/2YEM1x7+eTuDofOwm6cNieaFUak8O+B1zRcdHhVTJAfOfr
X6gy3AMzvdpw/BI4zEO+jOdfDpIgF9Az5Yt1heVbx3Bmh4zZWF+B1wdJjLBJQl5r
/X58LZTOBGCgJonGpu+Qe4b4fO9zLF6WLp+5mygGuOd/97m6hk+rXtgMzb9XNkLL
CEivTcOF2ZrYHVYNhx7l1TLIqVv3/GdCj/CSs02QgLKoP9QOK2QemX5nZf9mv21s
cKHm9DOdC/ySkwJlR3ZSCU7RuyMKwSaN5nFdn9DG+Gu19cLrzoQprxEPunMC4PQr
EpL/0bOX+yO5Vqaw3U8UY1jVS1CyWXHmL8XqpjtMEuurUj7LWoQHgruRLSxyf2AQ
AD4+cJ8mstEbm7dp1bhurAU3yLGEjqVVip6oaX5Q4LNM0ZWq4MdtNvUSemyxCGHm
UDalPECoubO3mya0AxqJqlh/MejJFh65G8ZKgQum5z8G2VsVAOV/9Zghdf2YOgCf
BqolY3qUu4CG5l2HP0obae9/GX5Ps5PBY5GeOGt2X+Xezs72valULU7++jF/4lxn
yWLQr4SIczHYgUVzUnPEqSGYIpPOgxXY1O1e/iFlPZNb/DoInEcyUsr4nPY6Ce6q
PGYPQvTuVvmALdXeTMXxxkgUVDiIn8H9Sf8fnkcA/xAtYvr7SPcxmagXJ3nqlQN3
HIPH6+AaXYii85APFUUrrt/YPuSo7a4RUXcmiz1EH6O9v5INsEUYpPC4FMIhoQJZ
tg5IXh93NCMFZOpcgRfieBEJaMCZ5IWSeF4AyViCJwVM2Nv5krEb08OLDGiREeON
cr3tIhQQNYm5qVXC8Y5ta/pxKqgy5rlxLOEGE6xzTkTw66+pxetOF7l39RLBTqoA
T93Z2BxN9aPxIOBtmOPyMO/77Svnu6p5w6l7PrkW/XkmcnKhTr6ycf2BdIHwHvYc
U06dP2tVdpMGhaSLwsRsm/whYqqlHDvTpnslHPwIOFL1W2zb7HWhS8jbzPOqSaKF
6aA1MvLWrLrS3QGB6wH6KIOM5ai8iJwdhO9DNZTCFGwN4sprpv6FBtIa/HSw38fn
AUsUWbJnW+xSClwSo1yzqP/GpBIgSMlMhl3TRzvKqCROsJfVRB8ODIYyfxjYwpyw
6Mt1Xq3Wd6UYX0d+Af26+mnjDRqObHZjNRQudUTxYUeisWQMJCvMz7pFD40wQD17
mx9Rcct2yITGaGN/P+fiAkpeOoNgQf7O27WAXq764pBKKtLnFVA3C+8cTOlRa53U
K5yASFzG6oKjm/qcAdg3nXegxe6w+fl7qNgD2donqCCrqzXtEXBujaD8d4eg9maR
OFBsXll2jmyTu2+VJXrtwP72G7ED0nAdkzufQFNKcUeFYIY8wPX6wPm58l6T6YDl
HHRYc9wRbU+2Sq0Nq8BhBxmo3fSOMjmlgQBSbTEDh5pVEpDBMRSS/ZUoaTbIBaOF
vnk+k5voWXMVk6G+WjiMm4T4smK40m/to0kkaLKsu2GGSzSt799r2JQbCDqp5kJV
aEs6oR4QgHgaoQ5TKnEq05oFbaaD+rlOjPpj2dVRuYnabXDozr9kcQHJ/lRPy5po
fzJGVUoEoGmJYnG6Z6F9EOuFTQvmdgUEZnOqlx+hcKnoIR9RMEHChESzyQE0dpHZ
87+q5TtDJYnOkC6fkg19sGBTraTJxmqI0F/aLf/aADXHjA/Qkii+vbnuvGRmiOSb
Ci/GClmkQXz/iiPh19X1G5s3zdexjgA3nEwvx6kSllwGFeqM8ZRI3N4H4XZqnWIR
uEgMNXkJSQc4xBjTUoRzkdwtP0yTZM+/+3IYR5e6MhfBPUt7QEMODQvAR6bX98dv
a+buRl9Ofa2V07jem2X9CxCmfayERXvz6uWQsw7dGQRNXtGM1UeXxz0z8e1peu2v
eaGvFSmYNUDNoJQ3P2nw3eOyza4xXhs7hZJCmggcXNX4xJQ/0rnDzjMx2CY9vn2o
omy6q3nRabC5xbpYp540Jg2UU5zzbM5EkS1Z5Cj4sL7x3uH/WUwO6gL3kH7Qq6xm
QGyOz4JGSZStHIEFZM5qb32JUR7xATof5p00FswTHTpvBCGV7LCjCxw2vhtQeXXU
EmYnRBP++BRy6PJXzaOqeC817ovJKXAYWKvB82MMW/zaId543/U9kH54WL74C1g/
YK7CONHFEJK6p810uYgP8qEFCNapPH2agHhLv1+GqgkpPlFXbOeh44SsHvoL2t7C
HOzlAPFETEcnWw6AYsmIom3BtRWzMOiMxS6MRPs1gxoaMqmYc121npqQ8dzvLrtG
T0kdAKKWB03dEa27pz+YKaYieLzN/F6Gu5xKYxOJdEKZ5/hRSuoDsTm8q2Vvfc2k
KAjLrkWQYd0kuY4+7zuPKlFnctDBiEKIzxqUA9kLEAeYFqDrt5kaIWYHZHtQnfPH
gvHwLEcH8DnVsGSi+ZTjUXSR8PsAbnDAgN/DlLtuXDCXvfwjseRoekZCMyfR8VzW
SfIkgIMtb9n9bDUYzEeGE1ylKdObsCH+7kTYxzBfYPbrbj45/46At5dRGYLe4qkp
VknSays8bv2HQIS/VeHEsORnAw3NWyuEPtsnTPtURXaCAaO5BSAwlBcOI2lwCUDK
qXXiYYDw5Bxvm1H1v3zfIKg38jLfSXUDFiu9H7aW0/fNeRGF12ijmZB7ZRL7LFJu
ppWUyDshodp1sQOfpUgxHL3ctgEgEXmz8ewk59L8BrxwbWKsIDuUc37O9lo6Y+pV
QKsVjJXoEs3QqBWG1i/PJ3etWjIoOT7f1PK2uKa3XRgAj3QDuP7ajVUUAbwpCu99
QM3YGyA2g97/xxIt4HJo1gJmQdGAy+WbnP4VC6W3SUDGyFMbne6jHhFtDzwlOvK1
ESHsrkO2omwvtpdxHPVuKjf1i5rhJUjLOruiaV1CRg3JK0DD/L/HyyN0hxVeQfAF
ey7FIdCn+LHT65V+kG5S8kE7Aau8FWq8a+5AKC/0JCBm+WWUZZjOxuUF1wOlZmVh
isNl7HREKm0QNjdztPslDFEfw6Nu3hWcgYeL13k5vxz4GxEX4C17GZ/z0wc+Uvit
m+a3FBMxFu2klTZoW8ZkoScPhCoc7jVN042y/MTaLbCxH8vEXOpgM4pQ7ZF5pLL7
TAPzHDOjXfKqVLSnmUBM4IjDOtNaqpqD6FwemIhMOLzNi5udfMP5w+qZ+Dc6xnGf
HAvslEPXsTGuIM4S014tIJbs1gmYR6z4fPc63F9FZonWYZh0KZM0NOa5a4GAw862
F+/9j4DWxxgH+surehtu1FABkiIt1917sIwwTjvs7y6tuTC/Yg8YI5Ek4MVaWPUu
JO6tb6OLg/zrFIDoM8AP+N/PrhoUJgB28MYQ+ngND7qRiWHHQFG6aJh2w+owNQTy
K6iSiya7KKR1k3FuuycmYoWiRrM55YhaLK3L6PkZdzJYsuGT7YQuI8L6r9yMrBVJ
ZBgf/HzedgjO/okkT2WRGsGnoLPKCFnkVgjmbLcCBb2+Hqift6GGdwAI2fC0T96E
AejFSIlzhDH2GYPG5neJoNHsTbkK4KNP1bjTCV5vskPcxE5VdzqNFssmDIMSiWxW
bQbQ/nwOGQEu1hB8D2/fF5iDLB406I3EWxkunN0UBo2b1I8lav7gxOscN8IbEsVM
e6y8MmuF1AER1ZXWEshLG91E/Li6Z/WuBv4j6gDb379acDiEt/wI68KXUraekady
OZE8lD7E5eukq7swwe06qJvTdphxe05ru/U5LObtrOmW6v6ctZCdpi6Z2yhyYOvk
1XpXu5ch40GBfcNZjhxzbfWh7pKiGnqWa+yw3d6x1kO4UdVg9aOb5C5uh02gADdi
knZ628iM0DU1VIXP1CBeeAk93s3ihp2KaRTkcqlIggXO/EosfVfZ6tk6tAseyf3D
sr7neujNQP0zVbQF+arEIy7m+N0ke0+6XaVk/1at+jgzcqOKYKUmgAfZCy0GxLZ2
HRqU636SrjxsFx6MDIjoikIUq1zF1mQe8xBFrTDvH5c2vBvqgp4z/watfkWObPGg
NauTlu6ASBR/GJZzzCIt8/KuepgQqztqVzHj8ggWlCc2RwN6jENSEJtq/fO0vJba
USXJpqF7X4yVW5RD44hihJ5Sm926cWc/5IFQkeZrZxT7JMB+QLjJ0E/TrCkOeSK4
/FdYGBdl9Hr1+3Tcf7tlKniUwSdtlKMxuboBB5B+wt9VIAk0szMG77wdaZ/HTCtR
7ZtDFBNeiODfZAWQ0arrExFCo/UMcy/fFsNVXSJVM0zl9yZRanYTcrSf6bxQY9V4
qxRrlxbfpRqs4iLsTuXg3KBrwB9P1T8GP3XOpzcb484LKSY1eCC2JwMYDREFsZk/
rXPTE/MS9tEk52xgh/aPMhYnOt5k+xJKPu72u1uwngwvhzK8cSGNrkZtneY6fV5x
hIMuQmCM4vmGl494hR56dUP+grIvb3CparNMnZ2c3wvZOKOEvjkb+WYVLWLoIAVf
GeS2Mb//D/fGfshP5q67bMFQ1/iytazps5FPzj4FyYK6m20SPV89qQTQaVUsLsop
sQRgf4/iklb29AqsLNY3osD2br5hESKdFaZ22g3z0lNPtdj0O/dTRIBET6sAkeoz
bw+Y+hbMcNCDtSBXZrHaX+Kdpo4tJhmdE1u+yCQSzgsIhpZXipx/pR4JDlEIOSv2
laT4Vrlu+GVlg+iY7obyCpoJydI4aYfxedPDS6E9AR3GsjGRoEeHGJbUT14CMkCC
KPlAFUqcJre+4zWJwfbhqyjMORyBJLMRnqY5ElvkEhhltHAu/mPrWp4vOPjSlDgN
wYYen4LYKVmCg+HHG3AYmpzY4+S2OTAEDGC6ZqJ/hMi0HTilSvIkoA4SMNMZwFqe
p373huDrfObXEo6seeoVXPD7p3U5P7amDWZMLkTBx3CiimFCzPJQAIW9z7jbsT9+
Blj+z43fxMfgQoUAyzIc5KJ/1q4m8FytgG3Wr5CjB2l8Z38XlMiN7MALFdO6se7Q
p97WVooRZSfiK/KX8C/c2OB41i0x3PdBWG7gBM32gpp76bCDmhLbzcQEJiiIHR1N
e/Sm5waeZA4Fw+xfz6fc8VMLLSgYOtZ85wjJQw8vphuoBj2owLDFdgvmf7lksaLI
n52Cld5al4tuAYzdUs0NE+jyrPraTOyMdtbj0KvuSBMrmAeCjPkKJ69f4VXNc6mq
GplqPjgG/zaBpiQ0rfiYfPfZYSMzp7WU51NDe1/ebSkdTF0IVPTxFwTtf+cHohFd
bLEU6pxUivn9rZGZ/7DJQjdz8sXQ++EilriC7jDYLgZiWkgsqFFOO0na57/A+UdF
F4RYg6WKkP2Q3EBqM57Wysgc0pS2BaLt696P2RUQ76WrCix/HMg6Gv4xM3POKLMR
gPkephuI0m3RpLA0TSSw9ySqGZApAPmKdsRH/KbPsOSV2N01wFbCJrdqlCuHqPFS
xPyRZQ6e9X3eC39cWgtUDrApNJnD9adDzh4NiIfJEiJayrlwg48onBMddhAXB++k
SKpHvtkQ9NtIHGVmDMeERI7NTXLDyB/kIXvfqXzcB7is2BrRkbDaTyR/EXaOLes1
qYGEHG7UxV1gnBqaRDe3mPzvewG72KSAr8L0IQI6q0y5m5pJVHwD/esQbLp7le4p
jtwKpevP+7OcPubcZd1/uPkkqPiCsU+EXhDm0qBp0guAQLshpYH9UsPnN3jc7Ws5
nhbUGAB4WXQQDk+5pjiyq3oAuZLawkN4ovPYD1sBZtMdDF7RaEQRGoNZFERaaZq1
fyrsSLhBeETzajbEY/YlBpH7jakcRGL9cbJMZu9HWmzJ4awTgCbvMiVebbGW7Aqj
Hh7PvqMMbki3Ph7wNJrJq2lhA+dSaCPyYJ4vHE4/oUt4xiaznaN4CoXXJuw8ErP2
iIe2Y3C0hgP30KQ98oiupwdbXqKiIJ5Za+Wu+0+O+xtmTvh8Ig96cxFmRixFtjXq
QC6MHvZOc7B6dCFCVqTuGzmJVPzO2YYY/zm+m4mQ65e25/jURP9qgq4osJj8Izbv
FOn4I45RixtWluTm538rIXENTQvojX8maqlu9v7Nrei4Gzf1HkxvTEwk1dvHBrmU
T77KqAH2G2RKdiTEnJadivNGe8Li3Vyz8Eh4OtafHQskLt190/h214iTiUXS3cn2
EkBZtnCDIPkTLluHlg1qL3Ar/hEHn9kg2+n2ZxvD6+X3BekjWOBEYGdsxgPKKPIM
oA9N+yUy3dzAsp5fSFe9Lr8meCY/VEOTafhEjCwq+edXCHHDaZj79NsXWuhqAjmH
212mhRxBlkH5spo/jcQu0ZSRtLcQyeoNYcVySVMMH/v0J/ytq6sw7viKgjE+yB7v
F5iATlXFDEATZ9JxIaB1FadUtIVnq7K7FOwNG1Ubsy6qfXoOAzGp6J2sypWStJRQ
6uLqqFKKAvLOhQtQRJ5+jpejlgNiehB8TXVMgHp1HB0fuTx0q1X5XFAfFll5h/Bk
XZD0J6XDTOLVJv17WgXI4sswdUlK/nTGUX1xHvwI0ThEcv/VKJK+Kc587/+alYQR
f5clsyvSjZDoC1m1wWdwnASdcmDCxVRva7vNdfNyqQ9M3Xfrf9ANMQiC/JHLvYS0
hP/VtmI5kk0zhFuTodhTsvpkgi6sLAHbpZlot3qZQxpvRLwc5EgcOO1xaB3xgtOc
QPOP0T/XvPovSUfgW9Xerih6ZZ/cA0ArA3VqKXfEKke8AkuHXa2J4FzEMrFWAyQg
CWCOBe8RahOopV0VH2aS+83cAEi64gPadm4FzDNi9mzxLoZqOJmER9+0ZnpUQKIN
SILEPP4QsszLziJLoyKwdqCJRxCjoexGaFmiotOVw5iCq2dFVDZm4DTyl7B/pNTV
tunetKrzBkXr5wVHLQ/L8DaABASl8TsofGxPs3WaHTa3mpfQ3Bgg3+y4AlHTLMQR
cboH5G/uROfM/FOxASSwIXdi+vd0gJHA/vd30MjDnZybDeCrEV50N5u2DejMGBJH
NBlJ01wr0tOxapaRhrQBm2oy1Ff6kRmmJ/z7hGt43/K4ADtGHrEy047/jQBmYN9r
uWYd0DcZeL7DRbz15P8aQtNhPYWswngxVYmAoX6fzuBkDdSYk8QVb92Nw6NwbIV3
t8wRynEfIZw3/BqrMCLtbrS4Oi/1/qR9pndknqmSnIryRH1/g0KAfIQdOrFdL9s6
59FtFyxBKQhzevl8sq0XwMjruo0B7U/4NjOiWdu39nQDLl8RsR8DEZMpS71O7Tlo
I96mX9c/XuqEJBgMgZ0MkAXk8QquccLboyABBLd8hGidGlil+fgphDy4Iz8Wn6n2
vQ/VD59uoVJZ8+jVNUHgj8ydKcPm5Px1sPeUVPe1eRjvn3tcKFtxiAu+T6ggVriK
6CK4rQp4PHo/NukFrCNIzJkYT1QT4BeDRYXvW3P1e7U51qOUll/b3uhT08TjxA7t
K0DpCPBROjlBOY2roZdbzCRS243OUt+vkcOezBAndbvFFpgwGgPt6n89colqHx5Y
FX586KcfSvXdr+Q0yidA8FaZIrB1mNA/FElP/m97/+Kc184/NkK0X5898Ra/aVKY
D8cqEBAmqZXF2oQr+aOP8JcXT83sao7P8qyGnrfFQvAikIxVlkHAOyGG86xq1Ldq
f8becqk4crK3dcCdqXR+gj8wMTon9PIzZhjeiLM3/yzon+OEdjAZv6WTyv+Q7geO
asbNarMuD7jo8iPy5Wnt+vtTAKVltCke8qikSQkDPnDV/YlDhCH1WjIsBwRWkcPU
rVtDuZF/JepzcSIIjYv4GiNXCUYCiatYSK8OibTljT1sFX1EqRr0F92Y7XHQKfRU
1CGQPanJ689PFI1U9vGkso1Vvo70yZnsWgT0uTM6aa3bezNa2PYeMA4lxHLS2i0d
AYDCK89Ws8lzGI3FSfSxkza4cRt8a0uVTvSWEwX3xZDzUP9pSoOeQ4p7Ca6eCIhT
oGcw0j9YrpCbjtTWD+cWNJT5tq/saaKxCDdGD6QioUlfBxd/mNl92gl6/IK2QLaE
+7XEDDihIFfAcMZ1Jbr/bWoMWdgMBzIXI2TCfQUBIgcBltPKY7e0iF9vs48NlGCc
bcbPUiDpfFPZR1XSMhJPnDg9nYBA9/fFDfTYiJ+sQMnhFj4bcQUlUn2Sw1S1eeIJ
5W6m7nySEchq3+9dzJyir8Pxr8QkH2LZRXTBUZRNqcOwKr37eL7PSXchu7RRoh69
wArxFdfxrjjS9wjOIAtqIUGDpKy9lzsoBFmiU1TCCGOszbjj+OapDMSkj2td8VWU
qMFZd/MdcVK/UBPIrYzIzIPPG3Fy5yl5j86ag3sVGicP9iiUpMzd3dvXFey3N+tR
MbQU31PM6b54/9jjAKLXvjH/vX0Nj2BdK7sl4NLvMkj+c7rbw3JwAJ/V6Q+WMu9D
x5Eu1+Hix+9UhBXjQH0pNCwVSeOn953QLo3Udy8acZstR31wBdAZjMy1YQvM/gb/
B96yICXsQH2TPpdnTcQSHCdlmCQD9c2kuL9ovwyb9WqVfrAMm1aQNZIzUhsXQO3M
c864Q0fs5Isn4fLt7eRd3eUyYp7WwrdEkdmonAOGa8zYzoIVL2tH6zZ5ODScZJxq
++L/Vm91ew69why5wCy+YgqAx0iolxAyHMeOIXqscbE0fZL6vZXL5dYWERJ7rLdy
GhBSLnjILy5nVyN+biJJHfSs8EkaiQWHk/QOKWNz4C7QB4j3OjbMT3dmaCmnM48K
hvYvG21nvLrbCajBLsObR3yQ8KlMLMsg8Dp/Srjvr8sbB4RfIzGUHYl4XApbJl7n
L2PKkmd8+FJCkItw29iwySH6kzZoeCghLT17lkg0ToUs37DKNIkWHBsgw7/mA5J/
uTmtcy6peCIQ2ZZk8+YCsxS4X/diww8v9RUWO0vLtXOV11HHu4rxPhHU0xq2iSX1
6b0OQ0fcp6bEu0MN0b532etScmLhp7txM8VeeV717NIZMTqpKNloWX9abjkpczZd
qwW7DPYyrA7cDTcs9OQjVfR0cC/iWgY1QP6J1hko2Lucn5gFnx1kHwJAKrxc+bhC
z1wTMElNfq6gI/FedP8YyCX9O3+oT4YrD06sgauxntY2T/WVcP1C+TWAZ0B0bi9q
H48jal4v6+GxAAgm5v1KlB/40ZsOqlYjAv2nuc2R+uJ1aGSdlMXRAxyKf5/uwmjF
BOk7WU1YN8eB2yAyTdtPoHoF2KLjqpmF/y5pCyKDlbpemYJeLfbv3uAHsO3+apgj
fIJ4ZmXdxWV0nJxl4urlhSKn2h5+FEA7bMBy4iCqySxxnfGOPlSQhDLrUgt35Lzw
blEl9V5XwE3nmuPbAZeyNKkhGKyekSQ7CzNnaZpTRzu/+44+dqo/pQwj9tKRIRQw
FzpdwQlj7bO77DvFTUuwg8FEvKLmBumc/rnFrrMPbSO2MK9vJLjg7PP1XQw/GPEr
0XxEVGwI+BlcgL/tJHpKDbl0fjNUT7O0pmcx7WuEtOs3+jfdxCfbZY0JsXcHshu5
J1d+h0k/YYlQOUAkHkcbsv7Lpom67XOZ/3JOG0ZgMFOFpgdjkRxvoqxdTqCHxFQA
7EzvQus1g0KVJBdH1UbtdmCBFQ6zz+0dgAiGvLansGNXN+MyOwoolsePksRA73f8
bDGDEhdFWy5POLBSf1qCycAPg5bMwoPMbWU+3x9jsrKwzPemgnPLBzdIz3CzF9S2
XrZQvEFg3sKC8wJEaE0m4ydyxAortZ2gJgBX1aOLID6YHiwFTHkfcbri0FUqdgh/
9efj3KKbNyGdE4GIB0rOwis7I1QsApEd0yx5M70U+zil1F8wP2SRkQVbt0/dIHBx
6z+OSspEfY7IO4Xp1LuZXwyIJgFcq5POLXgvaOOH5JFEUcq+z/EKdereGhRemHQH
0QybPfnnAozVxTLozgREY/95swFA37uDHFV0oPwe0YRVCEfiOYvoVShPpMYQ/LOm
djGwdtKxJLb3lTzeP74Ry/VU/HiGwaupaR02mTEDRzgGESDD4hIXDCjs1uADWt4V
L8CSKaPHC4eDc8jzmz3lnzJ1z6u0hEY9wN1jnIUyyk1KrhbQ1EV0o2ozYMuejydE
B88eAIwHmQgmhSxKa0/Vy0swfRs0mz9WcRvcixzGbUYqmm68Gvrx+soYij9useCx
36Qs7p822KiHUw9dxWr7Cujee+o5UH/Tu6WZnDZ2eUhAzr9h+vDAX2pxInm6fd27
+Vm1c7Flx9g+X8NYgBJ739pT0b9qXmSIes+MzsiXWiiETVaX60WQrX4XNlbAGVo6
y9kvHvkW04/ma7W7YIITz/x6XPC3nJLoMH6aF5OD5XKhn4Hh2jXzWDAiNrxlF2KZ
rl75msiyGD642H5UEQhVCcx+HGhCASm3SKM3RswcIeFZAhHsQl9Nz/wOwsNP0Vzq
bDnjUj6XelQfXNd+AwEDEQq4UMlECOZLdPn4JvxnWh1Gs0GzRiEF6LT+tIDkwcjp
jRbZ2eoUqIschH15JA/KwGrRmnC7PnDakl0448ydr3Bsl74Wp5MGADku0uEdZiL9
QNo26lvlBJIQXsBGMxlOPWKQ8aym0E4uCaFvxp1cxhUZOW118pXpX+f+7e+m3vjJ
4dBJl1Ffg15t8X/Uiqn3/ylg7EaUwtlsJtgPGa4R/iMiAvwYLm0DcBs9wNtZrlUn
vnfzFf4yDRtmcKn4PwDUm+nExHpNV6P1NSxVVhYr1ByPGOBmBTgM4WYhlRTn2u46
YG6hUYQEpFwZom3JFq5ynGPx3VG2EC6z7nlJEhSoB7ePJb4cLXLef/N0iFY+HioQ
PI0RZeL35xzPIrHLOc0VuIkql55QPa2K2XPKEiIQnvi7utk7Ob7khTPuk7ewapjO
ukp0pwfYOsYbYX6Cv5tHqPgPhbJjK6xoVsORGxz983YX6T9VcaV5mswP06/PHGE+
NO1Admap5G4kQKrnr+a/zj8xCMBQZbhKIf9Na0+6cmCUzOaj3y7pRyTT2Ks2nYC3
lZi0Z5hmt+BCMGR0s5dYhsaS7sjvYZc0Spqdn2g12XXK71m1bdmY2XoGLS57xUFo
72xxcbMAiahE3/RBMvFUaww9SLqdYJU90CDmdzZBtwtmVqHXwMdOCeAzLUo57Bp+
KhdSSjDIyPZlewDUgOvawSPd/tTPepDl9l4T+JnIvqP5c3QjP3GB+K0EZZqNK/CC
LzVt2s7hKAln5x424/zYq0eqM666xklGBoLFXY7im3lQWpwfRRwkBJa7v0k4zzBX
f5Ioqgr3Sbuu+e1g7JYdJ/c4tGv5YU1GRxUqh65Pne1UMVcdh0ZklgeZsSq/A6qW
h8BtjV+uiTQaYiJTpFLqVwnJ9xYU/joni6HPQlbzwRW3W6pkzGrtOslGFRarJ0SI
NExqnebZ7bpeXmkPCO88iT0B9abquIq5G8UVb8mE4YyIX43yqqnqnMcqOO7CAFtD
cfzi1XTGPCzdjTQS4xzetd0lemEc2/h+zwPeqNeVrj02NmOnaxshX3NbB8r9wo5+
t2UI5p5+gkuTPK8iz9A4J5w3A8gfsmoRCdZ6KF1eV9YQ1s8sc6R5w1f/J0RnBaxs
S9hpA8F5Jj/1X3YkOswttZPx9TBwLRMB0gD93jyKbbSo07mRgy0G0X4qjmutSsni
6NNETvxrfpjpWd8i9/IXyUMieDw6N5jeFLyux/n6PHPvIvY3zumtwvI4sUWBqDW+
PgWN8RXtCvRPJUviEObTqKAF2vdzsuM+neQB1FMq/bSAzAH6VjcsEHfNVrdU6CgC
0WsY9/R1vZhkz3F/KY85Omga+xs/9gLY9Dj2wcRROYmbI1Gnj/9/UPCOKTj6WSu6
HMZuidOlQugu6FJtXdUq5mb7DNImnllCKPID4CxUl7C+zGxw5HwGa2o28MFleZx+
uBNiyJzf9wkotY0mjOA4NYQnbTpCayL+hI7l1izCDJHDw+pV0D6tTGOPRt/bBgEm
KW6hrnlKk36Tk45Q+lot5l6Gr3NjJyKcgQzHSue2pxDZFZjHDAW6J1Aerv1uJ5Ao
/GM2hM2nkVTt632lqBJIdOKcR1zECQYqC68DRYxuKGPutVPdMU31617kqQtmXgY2
srM3A1NxKhbk0vUDA6iPwiZBH22x+mrcwCpJyB8VjfjS/OJzfd1kGRaGNNbafZXE
m24DYV8dr9fGowNjSgEtHrAwWr2E8UAL1gGIvp48Aat0VADwccDkl7dkZxWSj70i
IIPUGe1Cg5ugAoHZp3+CDkuLlZjQdTinM9nVJ5WlqD0UbXYT84QCDAdgnRSz26nd
K5NefahTr7Zf5OJ+g0IYbT04cCo6/uFfmZfFotz7u4OK2suPPF4C8M7XVUJgD9s8
CuFaGDgdvjDGQKkyLas4LZ2eNyNSzHHWhV3gRLs7nd4H49An5AdYQcWyQHJ2oSW0
iusJtbXmrkP++BWdgwkzxtshQZlWyyP5eWAwjbaDt9idQJzmPggP75+x5dtibyZR
RFhYZgX8WvbmD7JtN0C1+pY3lyTMN+5aCzWwM5tIYmAOTWwCnAm6qOrl9EBjuXpn
Vm1mJD/R+xg7aAE3jgEb0NA52FRHfQ/FajxNG/AYHdFBw5oHL348haNCeSEyFU7b
8uDs+0wPL5oaoen+y0XLh2JnjIHcuFWvvi4mW47cpaLwtJNUBQSIADCfNGbSi1/w
Jpo+D/v2i121Iy1FCRHGItuEcljtTbqjLJWYO5B0YylqYfyan9174X522Mg3HWUx
So/pgY64k40Bqw4amaobsXvdS5QyzotJsAHEAO4c9/+Ahk4TprtuiOb9lA9X90/a
S3j0YX4Cy+LfDTjpsH4Kyy1E20KEc120Uho6Y1vweNFl1rbNvlsmi5HVost/9qCL
AQFxeeBhCStUqwgKKHd1Ca/xXPNMWR9tSFZ5VzBxgbb1lyB2VS4Wi7+naIIMmLsp
YQ6IXpJFV/Dap80Z0FfQf7CEHpWqKDXH6CvKeckUAsJ3DhKEk7GTK00FSniycY4O
kxK0dzvkyG53H67frC0zUuCeOx6PUfKYlJ1wZ7hljgTsNdjilNFJwXRn27xg5h+4
+8h5da3l6kqkuNc14swsYpxJFTPF53NPaBHuLgZbSftBpXp0dZWgz7QY2pYmZABz
6+c5s+wsykkiKoOiu+9Ij14BdsTT8I99QuAOqhWeCzFoVQ8VwTJWR8EeUB7DaOtE
b9CWIzSxV8IVSPJDTJgsa7yH4XRLnd+GdCtI/CcDk9HLJLKBlwBWj0OFG55rxXFP
g05ymXpl6dblAyGiCooBbqRNwFtQjy2byTD0rTvghSJHT5y4mENuLDQKAA6Vuzp0
LEXo7vMHvvqfml4qgJv4o6ROh4a3ldwYPebPwqajYNVsx5TYcR7aaSEzf9X0sTnB
r8/PiTkzTk/c0UwHmAFstD+rzULGWfYuRDW+vMdkg8m2dHuDqaOcUtOmNWgnFfe4
UM5FUwuU+ubq9bQ69EixnIxy1A/0D75LJ0JjzjuOodGFx3JZTwUyopBjXYJRQWIW
nuMtzvRaOZGKZrMdBSJ7LOR6wYzoYlWaVDFZ1R5j6VBBLoysLyLHUAyJR1g/DVbn
1wppa78RHsZX/VM2XKaxjYwzjjYohV63lS1bt3DfJzp6RJU85kVG+NANxsjhXIFV
R7bw+jU5eWdvF/NfiqrWv1hiWIFgb1ehvOuQ43EANtHw7USF0DzI6YK/+88n0BNA
qB968ByWF0essbKIZO1epumbQgnXL4KaqXmgNAHAc9QCbLEltAQZRMfzAKF1Uahv
KtRAbDJLN5bo0iMAOcaIdvhz5x2b5r8dN+GIMlETzho3yVwXOXe6BMEbs0/zxaYM
jNaTGlP3FGiaUzV1FoqWOlbWSnbULWoQM09/1Zrw4xKcOrJ3P+64QRXJ4z0DpW3p
gtDBEKe9pFq/si/3853nTU+HmWhpwK/tjIxKtEkk7+uFc28o9Kz3EdT/YmXNQ/TH
8nPW4YFLhm35qSE7XQsp6Qbai+Z2WEZlWouVM73dHmbDIgEy/v29xAQki8O9GdT4
hcxn9M4211eJO1c+s0tKxAhOPS5K41Qd31C6Cv2zivRvQztJ+xzOhE/jL6vF1w1j
8alXCasPWll+1GnmGZgg7i6DzA6dDBrAMuTNpy/XmerltkYZmet1MbV4aBAZLrC5
Mn009j4wvtoOF008qDP03Vux6qNTyWN6K1hViEya/Gj/Q3vZhJXXPU700c8kiQHb
WlhQ0dxLsIv8hvfM97+4dH+JoClSUiF6XHfm8ie8V6ts9gdRscmcVqcktcbQNm9s
abbLMYBqvFy5salMOTzBiKmJZ4xeS1eol9ronz/gpSO8lqD4cOn2aCcZsGnksjeG
6NeWjVdAIisx4EjCjp4TjXScmG0s402I8bwKAD9Bwi1u87w9IrUPUkXqQgqIzTr6
doRZOKJDelEo7TBOwsjWT2yzd//WnjAU3I3WIm+lwRMWtPEESj3Xn55IxsJ/7hxh
5kpoZ0yzdcbNtMrZIjs3ezDXPK+tp2OigDDeRkTUsaQfzNQR2hazgZAx7Uh00z0R
U4ITt2vIXpNnGhVFc7pLbC/Qj91aLLSf7RIeUkZNTS0Iss8a14ikvt5siyO6MP+2
IpuzltxlxFccOZ8eaqboJnEhtLtI6e1dhD4MfA+4Ma58ZEMS0hRh7AWWSbV9gz8M
oLJCVL69MPPcM18KXnxUx+KqkZgYlJ7baTHjcIKPG5SqF6f/5mgjGn0GTMC44B3Z
qJC2t9SAIyDMHK98+j8KulgY/jBR3AsGiV9R6K+I58NU2xXis7Egck/4lLVlXcpK
e1ugEzQ189yqxaFcl4gIdjkY3fR8pqpDDSSDMGZ7WalsV+dy7u1F4wboK2Dzt2x2
/NfeZKW+Ql5h3elSh9HyAiQOcgU9FZU5lSnEwuIW4Gi/CqRUWUwXi8JK1GWGQnWJ
YdFh0JBfgGnhNPwJVbs7qdOOe0KEK6UDWBl0MtK2FpoGfM1WetPAUnFyfEJgFXKC
SvMya780psAdI4ONVBqZml5CtC09Fxgibe4saVTOmbfTe43YfX/PHtfdJQDXbEpJ
GzxwcbLHkJ+1cceX+wb0gdEspnWzBkzwA67WScgB3F4ajXqU70EJDlEskynQB1h2
7IM8aQdL2Z60BzWt3F1yrb9eZiK50LIh1A87OemPCkeiUOqlnP8zFZbUOz7V6Vdv
/SOnBuOx5OyA8BkoqLrrZVvJh/C9gOCkn1D7ly6J22LJqHYIJSi+VG1UDYEWsGy/
K0yoCx2/Dl7rM+C1KulMyyU5qv4/t0zqR2YwpQnxd19UaRGZrw9N/b94ZVHcKBt4
uDfWa9yHlV+hMXUEgOvZwlXhMFnIYdTu33Ftrg+7Qro6fL3Aag9HdbJwERZZuYCq
UxiyePPmCi1eiObRjyTC5PcIPjT13pD30/ZJbL01hUyIb9cm/YnTGz5OEp8OJsKu
no9ZNBsCOM82jTnjmlXgZaAdvgWP7XlcoLAl15/PleeL/cQkyU4yeXQtceUTSKXd
N/geobUZj2nlCe+5xLnWbe/3KrthNDid2czZ1iV1IIh1UE2Pbkd9isDqdYXTTsTt
dv0d7z4qZkgbgVuBDYC8dzbWjBqbV1PcMR3JW3YDLua2xpzbN9WL4tKfpxma1pvI
88p6z2O2hCsxDZYu4owwE4yeefvS9PckwTPAb2woKxjvJ8hyQMC150x3rqwXcuxS
Eb97Q5LNUixCpdmEz7oyPXoFK9Cqnf+2mgxEukX4fNuguHwmbrqZcRIfdyTIqwuC
A4X19zJpDrHpbB7Q4Xyr+x7fr3iE0OLDc28NJl26vdfJjED6TlGKQyNDIcRIAZmA
L/R+ACQtDGUh4YKLAgSrZXOuuKhZCQaPfeD/1d9fL/T258h3TARyb2VIlhay0Li1
z+fF+pY7ugbJIgy2fQJh6+buMtnl9F0sbKjhC5i+mGu5P7Y9z+DRXoe1X8ULb/uP
7lnTBsGH/eYzP6q+Np9s0BcygG//vwZyu3lwhZw+e7+DUllxQYSU++OEaxMTpcfn
4PLDkdjygjwdjhH3moTb64V2OuMsRs//pW/evKZBjKk5IxvO/G8bsKAXdHmP302X
rhVVKztN3AiPwzI36+TmFOnRbOqYpPwNwhJU1xIr5M5xDZ2IedB2cTyq08uN6mk/
RsRG8sXgRqagH49Co62G/j7YEpD0rw4Qbh6rP9ZSoJTd2OIfKDgBTmdHunr+N2yS
6Gm+5f8+0yiqxHOj/ZefAR5iSXkflfUqguwo8glPhbRfvx2M7G2QC4GYN0UOFs/q
XMrr0Tcye3Fvi8Jv4kM/bOVV0Cl7buyNt5I7scxrJYahyi9krjg3WvDPVar9zUNV
DwFgU853OZHY5f70cyIWfjA2M7SzzgDJ8k87q0NyV3BFdZZw5coePl8DCcZ0eKKT
G96wmex0XgVM16I88mhbURPkU/I+PEDNO3ObhsqkZZ0e+7LKlAvUfdJOHIM3D1sP
kw/WhX+oPzpTr0jjnJh1b7U2Jkbk89AtptfWse+hIFfUWov3fAVqNjerHjD7tFDI
zMHr0oy5eDhmx3lg7rsoOgS/7VenkCUmjnK3nh9y+sHbZU3y8oK/XCtulHksSpp3
X3JJsoZYJnX+1qwwnvkj5O28aEnravgOhH3kVfK9yPbm/zf5tpVy6wktkPrNDjLE
Ti7KmVyEW7E22qF+IEPwZvg1U1GeVOrJRbtCwqjDXCjTbsdvur3xaJ1I61fvnyVE
E3Sacaa5RBW2im4scfgskty/RUtuLOy6XFACTeSQyxTm/9kN8HPwgkNSI8+T+SxE
nOR2p8AeiSXVgodabQfyBdTN5WtdVOTs4wZoEewVLxfEpBopGfGdnLW7QcxC7bWB
2jieD9aWFclwrOgfJ+viCw/PXQ9HHAAHN5dXA4bIM0ETABsFKNW3w50HnIEqZaAo
DYLx5diqwou71tmUAsHkowVux5yfkvs5oMxrvgTnRtfYHxU9cBOu9eDFSiTTi+6L
rvu6irAu7mOkLfpvWBzyQr0LpScOPQdrhCWXSJ3ZqTRLK+/pZctn9m3PuHVGEAib
J31YlhbXyc8Xe69QbrYDPAANx6RXbTb8vRD3+YoC2YHpL/9jmU+qmTrI8GXNVDA2
kYOraPyuOmBX2gQZVZ9HEjGhTn7xtKaTVxCZXPVDMmUQb3tVCgZvAP4WqJrvwvvo
UNo1nQfPmsZr2o1zHHogV5ZFXOUbe7/6fCGtxRAhiSjaUn8WNEzQcsIxBwBBKvn8
e5j/NA2fp/+TX5zgmgk0weXr57OZKPh1HY44jr9nmKeD830ZSRk/WlelmzD8FaS9
fQUCpFxMNMp4jgUAMMVPd0L3XC4L7DSCO7F/WmpgI51mJnOFWMhPTXRR7CIeabla
yePGSPRDF8LW6TSJuCOpL7Ic7qwnERpWI2TtRdZ1miL0AMpkEHtERjjeCtHCDJDc
QiUiEel/PQh7b/1crsCOL8GbV8QpfpuDptxzHE7sqB8pcaCHgoZWab8mTQmOEvI1
u368kVnsJz34HCbs56FKaMa0VBnWJTLJxaFtV/UVWK6KQAEoVWVOWdZ0IH/U5Any
WM/U1ZXXoX5RNYGi+CaQMIeANCbRmOqreLXr4JU7oBm9inLQRtxI6xQoaO8TEwtF
KTed6caK11X6oSKkDfYcY1fmXF2/LxWyjrMKm8sllhV+VTu+lfsLN2XG5XQKo8PS
Ai7pxlWN6Gho9tG0AJ5eYZFyL1onerRiJvieVc+VpANTU9wAvpM5M78CWOUgGnu/
9nIDnLwL8CEYKz//daFhPsljq4/wS5oT4xkROYDeGsc2hz6qc+lw9iL1XprsK99e
4p7mgt/BB/g6urdQPtnUBKR/ip/Z4GgSxRjbX88AyahrKbpCdRomse7KhBnaRJh5
JbQfFFv+9Qzqsd3zjJ9i/i/f34zzyOtTOnqGkFe2V7Q1ageh464GOO1yDG73lQn9
DR51fuNg16OFCNFH1MySlSq8t5kF6qFe2a/+1MofzQlJD2rmnJ34mW3ky64dp/fF
h90EeTKz8pbchU3i+kQhMol5JO0gmo41+54ErmgxJBcankj3MXdKkAtfUk94/2cd
NPxVMFNQ4PuxbMjaqAw9BgMeI9gW+FdwChSvadarSzclwcoveMM/mwcNZFgVgsKa
ueT4h5hcoiHqnjJQ/f5DED6jwaxwvP8l4CYViDOcSPhEsS5zZ9Hohu0vtLltTYy9
WlM1GIuuxRe6a0jMjO4bYGUzgpq/4XBFB4a20tulxlJifStuICYr8jN/NWp6WPKo
lDORl3O5eXuGkuL885+kB4evII7iBKp23AG/n4Lz3r2WROXhVV+Ag9f72tz8+hDC
AreooT35HJ/y/TXTNl1KQGMDFQhF+ecI5vLARC9TyIOKaSGNt7kSvwkao+kQHdD8
fHpl49ffBVoYjEazInmSUHbR/uzClDLDht1ug5wv2HMPkLsMfspwJAlHqsfR21PE
oA6FSSUF+LDdFUAJF7zsbjPtTb0i3Yn5QuZ97B/qdBABkao2TJYIURfS/qXC7EmA
944fSutXhUsWRMBood9NcuqBm60snoElCya3yibmt9QF/XaLt2eoTTbmbjsncXmX
mEMOqftjM/tmSpFa23QckbE2p6G0TK/IDJRIYlkXxUHaZVbcEJ9H4eGpSKcS/1Pa
36GGVnfAY5A/JpNN5qLvRSVm7mbSX+n8f7CPL3lbzouUxIbbU2cY0p5jQd7ZOzgg
0KjQRHbEC8IEDJAbp+6NfyWE9C07LQ3BLsIYgr6lWO3/l5hLkX61OKJjBhHUH8zT
MqsCYm8kB/+NqKnPqgZCbbM/w/ls6uLx46VCA9bWYwKtm4UIf3xo/L1QTkjoO1M6
J9jHtEtQkVa5lCSJAQP0R8a8TQ/nJHNISkUuvs3U8FSZCEFUT28AE7PVi3+ihVdi
/2dmQIao/fk0AkF+YSXH4xQ39FIVA8gefQpKkM2vm3yyjwnW1H4uQBHTQUHcrk8O
SmCozG0oO9demMpR/wBsX7a5npnJy/TRzYiPUuLb6QB1GofIcQH/22PYrO/2WecX
sXqap0EkJFG51AiZq9pIUXK4Zb8j6wSAb83GfYgRabiMrakJ6+Q3RcBM+IrAMR9N
1L4nf24L/4ZdG3/PnwY9CO7oF6LW6t9tO1z+kkTxC+yF0QTlag2pQCYBbvblmQHW
kd5YPRWMJ1AZ2Y2sNHqrRxxA3rG9xB8T3loKwKdWSR6wdz4cwlrOsbznf/IMQUuA
biCoW3I8R0orXgXaTj+f+PjDbvJgNC6zztOalgQqiQnPBgs63jb5yxSOekQbbqRS
YCSvlBSTflyuFanAjS/iehznsC9cnCYn+I1xIYmZxTl1O3aEONqkCRc0JYMh7Mhr
6O5B0otqXv5JEAQiIiC6mKqy726mM0oHhpkURIHF8/n07jqgQVCkLHWX+f6nMRNs
jH3DGx5NryPuHvpWB/kJFdorxW98HpoDQVf2hmPFFn3+mP6qC8shF9bplIAu+EBT
iiqCe8Ba0BggDDOAkcXSYecKppw5R96qzBp6+qPWShQimx8KZXON1opmY0Fwd+O/
vFDTCjphkWP6fcMxj9JBgf6Z2eyChUO0jsrcCI1sDCJN5DDoBVITBYuI486HW8e6
zRUlotEZLqsYhrEY+NbS75UvMEFA0QLjTotgnp54neklJfO1bm399tKQ56rEsX2+
yFG00SuvUpkkj7qRjxtx3NWka4VCx0Tlb1m1/xXx9Mdka8x2cCN/v9tSEw2WrJkT
C8QdG6S+08DdU1EajPrz0DPporJqVWrayPj71RpLYmY2ifoqkBrN03UtJmnC8U6L
OVoDbWkSPHThsbTmeeIMOcY3w/5Pt+BaRDSGJp4lvvGRcYkUe7ECRnKtFhEzVeYP
KYmsYUIxmNaNUQU/3QOeSXysUKM2v1g1AgIDkiVb5KRb/cgzw3Lj8SCzEBPgQHiV
xiTQl5oAOCVQqDw82QU9aTOeNttxLqAvd8tkRdr5yjHGVhPhZTx2aqxPd1LCBrn6
fAcyu7qwjVg0I8JRXYxx1DZWuQ2ZXkiuK+bImfrxyNyel9i6vfQwpIy9n9ZDvfYh
i7d0FRsE/2i8OL3KWiW7LStRbzE0rdhHgJKyC5KFak2NfgKdrinNoD3SZ3ZanRmY
sMUSMbLFpcpMtR+foEX5I1wkHzOMQwHBJTevk1mgXAGhgZ9c+xPsGC+cxnH/QGXF
0CqlkT+62X8YB59BZOwtka7kKxt1utb4D3DlsGoTskKXEmHdvxrmBCJmBQsw+4mO
637xjeEMUOeE0WicoA50TlDyAlJnYwFI+lddxdy9R56kDOGWbD2GA4Et1rvyv9V6
s2POtNOTWtfAD1WBOrEGq+1UE6HbKn14V6kyMi5oMhj+s4Zqj7r51RUP7Cu/e1p1
bSwrVqOdtK3v6p/jkubATmCCxuAUyAnV9TrJ13x41aBmo1WI0n7lcUNsQpgXGoEN
DkAvzFIhLgyVnET+RsxODpfQOjPcEtiEGhWeWxjtHhAURwuvT9yfFomt/crDBMDU
alYG8mjW68bUjVPRNJlxrcXDuyISaSVz3yORMB5MYbT5uz4EdGUuo5RKwYyb+6Od
fE1SXoBkrqVDr2feoHLwGDi1rAYeLofXjzQw+NAuTCxAASA8FGzcgtQcFseT2EMf
XMr+R74kVESc26QusnL4kP60DfrUVhMBxnwrznLk4bTfB1TRWdW502WQXN5q/ixP
H5DPHlbPHBTuzFlp7ELBlkPOF+9jn81TnSRfhnM6rsQDQY342fZ/eeuMaiuxvdpI
iwIrJegEkVWZ7WYAu4nJsE6i2FIptoO7ZMgvBCMC5faNukl+qUA9L3AiWsmGmx4Y
SX3bSgEbXISJcEqbmkuQL7CZz3YhS7l2Y9CRWVdeuJq+FSr99Z9CeeRhWF+pqqJt
P834R/o3wPSKprtJQ8uXMqzRHbS3hXjZybb9jIEqk/o9p//qCnIJVVnGV065zLr0
pi2oOp4LKBhkA82rWsjBnnPmgKtZkCcs44y/WQ4t6mw4AmnCmNsGlbUgCLIOm18N
rPjFVGbNoxvGV67/3uUhV3fq14Mh1bv0jdHzf4PMASYpWFkfSjlZE3+weWGMrjma
AfmqJFM7wPmRxudN1WOuH0K0qmjj8uW5LxaWitnufwGWlAvzndqpeRCulQf4z6fk
7fvWHZ9+Pkniqp+/3bPixjFbXQEnjNHUAGgOYZU8d7Q9xFWZfGQAhEPwsaiGMHA+
BajZjcYOoKlzuXH+Q/RPVlP7vda3Wq04vm599akKRHGpOpiAp0djxaIdTLVOfPou
sxldOQ8E1c46uZ0bqKl6Nc785SI0QJIpJkLyAjIsOrkqxpMlPekkTnTgCGZkMPzs
2zXtpGcabFp+Jt2+65EG9HdwRWVH9MYeGnNObinrtaf8Wms3PoZaFIBtZNuO9Yy0
mBrwH3m/ya3idox5QXzS9zDBa5V+X2ChI2dKHmVurH6aYX2ZZWcQisNZI7cVcw3r
dPztp56lWRKkvEex2ZTVv50WYN4uso2cK1ORUW8f4WUtzkIQycVcW0WqK9DiGfF6
58XVA7or5HmUTG9u6bBMwWZ2nxgSBo4gIukon/Hw5Ek/b51WbcxXgSyFaZUTO8Q0
7DweE2HNSUHmaUvzRsq0b9BSrWRB7TxtyhpoWbw79KIzwk3gBVOo01rb+xGgRWPu
OadqrcW/wooPL3cd+48LkgF9m/M1S9Fbq4GT932T+FdnWzxssoCzvJQHCvC1Nx5n
h/7cMzzZZ9ah9xuVdrHJs70B58+zs0Q8RMqYWFtUG0d7jUH4cjEIYtJvWadV9osf
fPRkpx+ohr17QXSuixJMbpLfcUsmFu0y/XDg4jAGAq/8OgBrc2nDO+ockk4Pfi9Q
9MIFUj0PJO0h0zymC0b8VoZjxAY9Q3Fqqr8NMxHPliorMenx1nDol9t42nAqKvXL
izTWEfFYzT0y/kJnXz6fFHeURPTnBuVdAeItGsCmRywd3r1D/Au6OKmi6lLpjLb4
09lvnOyr4OeLPUltk6KyRVtB1VPv2XD9CyWotZFrETRLY8FGIZgVrPUyuTZ+sebX
8RfrGkqzL22Wn35icZH6t90YK54n23HP+pKYbk1S0xtvncOGBsfyvvfnGi9MX0Km
ps9yxtTzQMJNrrlEtA7TR0Qc4benTIowvYwWT88zhApzoM3HYiRUzK5yrcIjGwjl
mlhFI914Xf1mDPAUf0ceEliQqOASgu2YyVk3CQ1iAxfDR7NAdrb/tIpVIYIdKGp6
4U1sLJLWZs9U5znDowvXr6Mrtz7ps+cssmK21tk3oAi9ucxlUWnT0xJTemTfdM5r
j3uWWUcPQ7aPE9vGvNx/8xBMyor7RerSNigrYMRfe0P3fkN4yVGXung9tUD7NKxX
AcQhRbqv6Gg+lUdbTB9cULLsc5mYoQfhhkfL+u7DPg/wRzph/2fEthc17t1O4Qyp
dJvJ9zOSX4kqcaZDWwx4RpLnKukP4qdkTrsCvxce+frgHSwCqQx/dGuAhjJSmXh8
LLvgaFdGNJ2SDSfZtte6/U+JCh+zuf1D+pEo6R5hH4ZFxkz8PYxM8Xei5FWCAdrT
tazwMAMc3EJjIUQCm2TARolEsVt40VBKulVx2EOtWlTiEnXuvYJZvtztKNQ9x/Up
IHpC2AZzM3i0LELmXbd16ZkPrG1F9vQi56zRa7hWXT2/aEWIXN2S+jsZjBuk/TNK
0BmXlU4FwAbsGtA+jzVPAkrvIT5Mx9rVy+55XdQgypsMG0FrtVZdT1SVOFexUQhY
pS4zuZ2mfPdgjeDUufqVNLghz+SodmENwECecF7B61tnYU7+uWo9NZRloj1zd1fQ
+ovkWzH1kP/qdaQMq3frbIVhURqWyoanpU55gaSQpxDey1zBsFbd8SLg3Z2RIorO
yMd6XSMNw9uIlimG1DuEDTgGoRV21E2MW5o2cTWfgn8cp1/SEcSeavsH5fZmVibD
5U8qCuhGgwiNhJMtICzubQtYYHCHkacTIMRsBkUIyys5CC1WCz3sfGPyGGRkaWQN
VFMnCdsnfM1/4AhlpEkGeEqbmCigCd2JKVY11bBfFVWvj96C0H0VQaVq7rx1kGip
IHBbtHeQfvnPJRYrW1SWlGxRXm44eGSVVMZ6hyHNcG400yj7yMuzt7oLMWsbYoUO
BPawmFPLU9VupAeqqKq4/7Fzp1HnNPtKEk/bmKpvjDOzT+Gpyh1pnYbdRnKIJk+5
oeW+wFiMQDA0uZTFK159wTLPhxKY7pEBOpvM+LxJHZcJWTcRuFIq9US90yzxYNqp
QpEG3L7I1X6iKrqg48lifYWzR4xySu09QV8ZX/D+o5DldiHIyr4P7/AXzDNTiv6t
zjncrSFTVPpCRbic9DjP6BtXTgA/w5rb1fVDDxhgV8raYucSjyr9cNmcEAhBTqBv
Odr9mWuQvHz1RGANnv0go4mBnjWts3oPwmvkhk0yVQ/9+AakjE4mFTtv2cyNCUSB
e1aDJi6yn4+GSeM1/KkGbFX4wsVKdPiq+OCb/LdH6qPXnpExTkXm6M0GM42lIwPQ
SP50bP6mCEt8lkfVBEZIqygraD+jOtQAsb92STPOB0B4JXUXxnOZy3RlRFFxNxrx
YJ1zN1xZIiftjOBb+VKD+t9ZtRyR7tiYyPNixsW4/hBIQG0gDpjZWNCSnmltougU
Wfp1Shs+TRGv8f1w58GvwVbQLDwsT09cJsZ4LJYpksbD5z/1CrEwfjgovFITyurO
EV3eh95hr3q6aTnGG6XGXlljbSx7obvSz9lZaGISpYVt+BtEsITrjka50IwGMIsM
k5GyjVTIezgcDi/NDEY2qcbiBvla2Dx7C6r1RXunPTFotAqWi1SCZopKqlofEM/C
eYnzVg0GH/gkSINNslTExj46YR3LBKbYmpTcFDCCVT+j0Z4mBE3kc3H8xicEW9MS
RE51MkA1COtSK+HxIXpkrikN+dcFDvauhHw4xiAgvG8oZ3soGyPx/cKiNoDXIm4O
5F9KHXqAb64eImPoeopgyB4MejNjrda6TmVh3Leju/lZMUK2bKzeV3V4Vvs+GrVy
ihrO1+LOR0vmjnkKMRdUk2VmDIWGpqu2EfLOiQtov94KVFZ5YbfCfgXDIkefXOdf
fO/A3AGHNSd5QHZP4swtwHaXCq9Dyjks/2buERkvKaBpCvddNniYgRUja+9GUUSO
8GwHVSmRE26DMgrMoqIRDFLiTBocd8K7d1od1MKkkV/ItZsGvitsce9gONRVn6B0
lmDiReVV4ZTqll0d+/1H24atYmfuz3BQaxwg61BBJlR6AQ2oMh9IJv0J1abrmvzE
ipxQrY93tUWzDyUJEyYwCbQ5f8HEb67Rm4FtAU20+77T8yQg8TXTWrPYwOOp3Xii
t3TQBK3Svb0Pt9dAaw2Kjj6bK17KPp9oz2DGHoJyLOqqy8tah4ZxhwHRkXocG9mU
WgZm3co8N6pl5rI+hFc8NO8FHCXpvJfg8y0WwMqGRGLPgx+ZtiuwZ5hxSMjXZzaP
2aLMbYe7CW330n5REJA2QG/kaKOcQMEgPpiISedKTM0/LRmWdyWkItt6Zk2KlVDo
3srXUEC5h+Eq8zk7CW6Ne5A4buC6H9/FWSZ+mJGyX5HY7vgZV2tGacl6HKJNIMcc
wdQ+mdXjuQtRXbU8/3OCy64WFB2ecXtmEefAeUIZRYL5X4u7HwEUNQNLKGzDmKLG
GCT7Hj48jCTdvX9u+BQKAS7DM8GDsVn+TKk8rSebMnmbnSp+p2tjbby0OfwAgGhV
uK//L6MgM1vcnA5xlsP2rT2l/89/dqtDz1UQrKK+vSehWZk6NCCh8RkKOMOFNIiX
1c1yzPNxOrtItJ2C259Ima7/QUo1boUrTON8uDUX7s5vdZVqLe/MKl2M/Wxz0r86
jhNJZ3fRoAETUvg5GUSC/W1yIZi1QoOniC48PVeF8U/Lmefah8bSQUvXhMXwTpb0
FzNXdQzgwFhb47oOCiswV9n6hkW3F3NzDJV33t1QI5Tiv4rt2BFD/NOUlL/nA26M
vqpCY2l39pZkdCHeqwokXiaCbRDKU6VVfU3ySJGGn+eME+6wuzbqyTCOzmOgDzRa
6Rbnoe+zJxbAtHYTJRWxvmxKha5ZsQeV9PLL7AsubiH3YZ+1f9vnQvRmR4JyVpgN
Bmytc2ita3EKz8D2ogHWr8XVT+jeT29NWKgOfyARneDNwMfq4AIEl/cM5GDrnyOp
ukav6tfk0mnArQ59z8TqjLnlPCBT6Q15bQR0UQqAEKaFFVu2KGUjOv+TkI8qGcWO
3XrhriVzhDti4hp/iqxD9RG/APkNlnmND9miLbYgV9zSRhhgVF+qGzQUh4x9gAQz
Jjvsl/NA6bQw5oplKY1K04WfHddoEwJ1Kn9KegSNQ5uAoCpVggeQW50TA+6yqcTr
0NVqmWwQmHyYw+vgOWlGiPSKTQysQ/gBAzBa8ics+T5entn+1Sln77RTZSGLSeaz
PwqnpbInwtedXDD8nPA4a+4IymGHS5I05jbOVl044yxLwvVC7K2HEvOkKLQqfVoM
+zttQhqOEgrXphYA4sm7qQZHRHHqCu+tD7VBUSmwDgNuQTJdNv94ixesRHerirlu
97hGiW7lnK7wtQoHAY0SYspIm7MxdSHwrlUQaFkAgGZNtBMALzx5iObzRzzj5Z8k
3SIkv7Nq9fL9RPfvG8M4FZgyHG/mpJGLy5BZz1eRcKOb/5IeuxVq/gMlNv1Am9bP
ktNR3/gTHpDF7w7pLnMlxX/uyZXFrVhor9lELBzp0J10L7gxetCF95XzmHnbDChT
9Q+NVqXyrOZ/6g3HWRCUBZRlKu+G9vn2Z4jBKPL8coARHDpnxTBqlRQIv0eajj0o
DhCXdJD8NylaXyafLnmvmdmjvkx2nlXbbG8TNHbJl3VeuwA8FP29hTSD8pGh4RSN
vXbib/spsIfeKuW3AbY2eUpSBOrEyJC5Nq+dQ6XkpqH0NkZ15PAmiR1QoquRgRyM
JXLN+wNBM4aKsGq/5DHjYYqGRIYUCIqsWDm3qgPJi3Ylyy9hIqniV98AbwWLj0Os
gpcPLuN2HagKWdQipdE+ZTfxlw0703h+o+pEXBCaYvoTSS/Rr8Y+05q/Pme+3mQx
Qr6bLrRekHD+H2PRekYMU2Ub6MWyz7gWNpUdhucigdZDKUWOJLqWwq4000XZ3//0
jt+GMKTKprdEtPJG23qT/fPpZd6YCutoxksDWbGyyS79/qYFykuCJoMc5mir5bVn
ZLx/icV09iLI+VVyAx2NISaMYc5Ot2Rks78kw+f88Q4KmB3agAna4BAyVJHJSoz+
UqVka2ihmPAXj/JazEj/Unj5wZ0mG2HY94MOooiRqbhBnI+UeRl+8LwU7zv/EZXP
8gzPd7LyamE2JoSGqLyZCWntYCjPx3fnSn3sR5fCDLPOQcxxrFXUaI59fcaJD88n
s7FFp9S8eBl+pCwKcjr2N5NsqNpWzplBamT067zgDICDYk/+bf0B+2VvbqAJgq91
atp209YT7BVZarrvp2U97hd8qe54lNanul0O1rPnnyuwJ+3YptLIpIrggVasKN4p
tKORtTGbVpiZv6xJxw7xlBzDBKLaR5zAOe9GkDfkUwbEprPSAW08/T8Y1qiwWsaU
p7ercdtOvC3gc9PcFia2s1sck+DsAYBSHj0SIIuEHqwCq1yfgXWCKDVFn0vLObUv
0mvEmULayvYCGD/cbx4+BgwWsg3gLhwWjs8AsT9HJ6xllkrCh0JHZI0T8D7j9WRB
xosH+TmrFc2gpSS05XRwNWVQdks091pzi3TcrHu6HEhIvLbPlW5Agg8WMyNZONxr
Mfwn5x7RAFjMpZT6Zx7LnD3klQKqwRfyy4LOUkonk2SCbX3Cu5dDKkxztvJwpzN+
1hQjccTOZ/rllMD8j1Vbrjs0iCx/4U3URKt//XrQ0w4Va4O0ihk/rCeyp5hDPLcK
LiMy6URw6su43wD3HKj628fW+LfF/KIlZEC5VD9WivzBuYLoKyp8PHqboUDTYuXL
T/8OlOwXPSoML/klR5j9U7wxoN0cDoxb/p3etnyAPYdhD1pwCpfDL/3SgJHgH0RW
ms6+cZ13hYLIomtyI90dfkma2H+wNdF2hbZIXUo/fBLqfNm2kBB/ysGJCTtk8DdE
hpUYind9h6SJn4IqqPA9PxlEScMc5Qhh21Y8tymmdZ76UUFPDsTgS6pebnAG5g+B
EyGd1u89ikTWfhbhzi3OliiMpgxs60Qs9CFCQixyLH0T0LpN/y2+JvB/lGImluSK
/GXco6TlZJuDnp9nB/zSURVp5M2Ykl29ill73nSKkkOWWSZ2HMNSo4LrLPWqdwYt
Aznp6XZ3+TgYcVzTGhRuk1Lu0fJNUkd6RGLW/DkvzilTO2JFJM4KZuLEXKyh0Z1F
ChtW49I8UMovwhcnJn0ilG13dual3/oWO9ZcvqHExYM8YqsUt3wJ8LQAtaRQIfYU
CR8EuxL++CcKOAUInK4cAGAQn/fH5nMDXQ98gO29uVxTxeMmLW9OTy5PIkQk5y6X
olADZ9MYEMSpbxp3DAF7TgtyRtKh6Jk2Yi4rMlxTNBEBzIp6nuxDiocsgSi1/zat
HAt9QnCdpEAzUZkllN7He0vQzFAtk6ghsXzLD03ehx+bbxgFs5bYhvVbjpyVDNF/
adD7NRecGMQ9bMq1x+s5DAzW515OqwS9lNZ3gIPhev4KBHoqU++LL3wS5O8wLHr7
ehdNOg7JxTNcL7Uf5noo2RvqV4wI1RUmRHsPGyhkJZj4i8OvJaIh1nP6wuf0AYtI
B+pSXXRB/oeaCHs+Mz0fXqJ22K3WP8xaHN0VVJ9v9k+VYy+/xqwyko3YjY7KTt43
pZglWue8lO78Nv9ZVe8PczIVf7S7aTvQGW22MYKU9y22M05Vu8bC7QN22cZH3xHv
dCxH9lI60n4o6kD3kCHozZQUtaCwn0KAoKvC/FEiv3S8hIHGC9Zp7cQSPiC+hOwi
g7rfBDehZvQuvo5iEpbpgmf+bGBPe0v2QLSSmiC6UKochtTFKOckn27KSQCoaoG9
xWmiLIYzLbFvG2PGrOzjjYGnL0GpDGc/okEfPSn3WS1jDDWwDrqeBi15StsAXv8f
8DgMo5f80M7fp6SOcjUzPjByUZSrQVTJprhqtzEazlAw6ezI+NxPPxJNE0GutjWs
xbXmNJY74VJWyFARYQcSGEro/CyIhuZlJndjA18ZTOckvldU7Jpx2AZqyiq2J6rz
D81xoNWL3h7Ai4JnJ8YO/4F2/f5xscAKrT3WZooJ54oTu61ng8TBQrrGbkcMcuWR
BHQc9XKIDND1fsRP+aZxzS5rgLoH/I/cKYTfVCNrnahQly1nhv/crhZskNp6xJnP
OiCSUD1yNqOPGG7kJAbULvE5Ar37FVSueas/YlpAvS9du5PwrO9MTwMZQW72lB9X
dipKhCJXsiXYp7gBbpBJAeg1bXAvnO8hNGx+5k3GTyzbihoWFk8rZDd4Li6794S9
zf7LyREOlA69bdGBTDKHB5m1/9aXMYcyHpOtY+es6lLpEExCKtp1NQ9XQME40Hka
uapep5pIr6eEqBx7dpWsNMBoKESpk/SY3KBSU82ZWfV6ktKAEK8zSweg7xaA4+iX
qLEJDBxV7sCLA3UnIPCZuu97qLuf5khWHShtzt4ew2/XyR+i7+BZ4Mlh9M4aMOeZ
1c3PVBwJprOW9SswrXT1zJx/jpc28rNEoq9Ke9HwwuMmUbuVhU9zffVo3LS74BmZ
kXUOTGuttA/R8YKAEZ4ikKlHMImL5z/85lbG5zqmBA+CerTvFf0X+ICGkvwrCpmr
c5kYfJ8JaR+ld+jI94JMio2ddfX2BDjX1uMuVM4Y4Q1hEG3p7c0Wjvdm13rJiCJs
5BGpqNsN+KmXG5qp8h203KhUmlQ73B5HYtooGOHPcvs/WA3NzdtPgTQ3lwyO4xpM
hDUC8q6F9hZOzNI9bP7cUQM9zF2ehA0uM1WNcx5uM08jBNfHg90174tnVFOtLozg
5GdnXhq83QTGwH29505p8P+IncbzMWXiJrdgW/9llSM8EuHt8m7hm8ezpBhP8JIb
BcKeUkDazVfnD00w5/jAMkE3AfTQV1MgcZtE/XpTxLHoyQfZ3rHy/lpauOzUNiMy
TAoMobUhuO0NpOU3IZT13ng48KrHIRGdRwUvZimGN2sl+ru3L5SwMASbvhkVp0YH
EpYWTZXqbN5F7vKpLWRjCsLUHYCxCodnGb1tV0a9bn9Mrf1LSIHQjXjeuJ9oEGw1
cvaViLBpHEU1pevtPwMu2WQGb+feLtmXPqyWk4gfk2x/Epu6cqarEez9yYKFcwfL
VdvkeD8dhQGIQdSmGpLNbSQcbK7KRbYpxyGL1hCo3xt9F8ERpLkBbd1sWcKISWh3
IdC+7ruaIstkBmTfddczzogcRkYGWV4/AwQCIVxx2L95mt6oxt3Pi+lM8O6owuax
m5YrL4mMG4wjgZ9022xqojnlCuhllPVATeAwzRgNyQ2BpRoFmdJjeONIP3D3Z9Pd
6TntLWov1+SK8+CLN8ih9WlVkT3IDm5Wb3Nh7bkRrNFuHFycueRFYkJhH8Md/qH/
SpClvx3nC//+9rnG+GuOgeWW2Zt7DsQ9Z7Onzm9NJXcrKPsI0CTVsfm+i/n1zRSc
VNd+0x/Eo6kDLEniVbx2QAUFgFmpQgPVGxGW767TRsvZKilh+dwfNd9axEKvE/W6
URxbIlGA4HioHJnKUTARAoq5BpV2eiMYQ9nzqYgIR3QC9/nkJM4mEUO+p6Gmilo1
MwBC3pl4pgwS1jEN16/5FUk37qHXJ0DNCvfHeWHrlyFDE0rUHcZFp9UP0lxBuf8t
qXcbw1g3CT3JBFrcLvbI79W3dbrrzpEHsFqzgUYgeWhcYDN1uoXu0Hw6c7GpScZh
2mbvz6nMka9KxyunWM/Qt4OYBGLHb7xmJM2/Ci0X6SwjL92D4G4BT6HfgE4QnbYr
enJo7ryPeLqyoNtzRaIxfiN3GngI/R5LGFEo4wWo0Jf0tTT3GcM6e5vm+fv+nWXq
qDWaIxmiJ2gxDs+gMPFm1mra6nwovLrYy/eVoW6CDqgbcTt4Fyfr9qR99rmrcZ4F
2LJJIcGPv7Myu/Z0NvU3J2SVJf38rgZe+9J8Nt66RUj1ubqNqo2cIOExXsFmHTFa
zrnRIrYtS6MkUA8VY7Svc3qMmDHcXMlizb+sDQUcL2T7R7WK+Rdc6KGUrdT32DpV
2NF4NtlYJsuUyS4Y+5wWP0gm2UymVc/Qwdnd2tBlhOyKOqbQUzb1VJtrug67Q5Hh
SOx5cLYe52J88wlcPnUbjyJmJcaEe/FX8P1VNNZtEPURVER+wDX7ZExK3npqh8el
XbJeGS5J747YOynDDxOCO/QrwipSwv71POfj4vEpE01f3xlGYwvm7kyc2IPirCC+
GJfew83CAGYdgWcEzeOPx4gxTuVKmAvYuYg/lHPajMyyPH1wZ8YQp9toXq985UYS
tu7t0tdGvcLXQVKVpmO1QyWyvqLmGStZfZyt+Q+7nMmZ+fHQof5VHE0wIySYqgxS
5Br1SFVjKS4eWanzxEVatF97Cnh+f3BMcSEmeyLX06HsbDC7JxPuBgyyTykGuaCA
DCvSU/sNpG4TBALHjKnSrXPHxFy6B4shMBAnp262uEiokE5J132ox/CzL7OZ/H7/
jgla6wUaQtZTlkw4hn1+Hl2vdo616tMG7z6KRogPhBrv5OX6X4Iexd0EakV58T1+
anFNvhY+GafBn4+oBOHtVTTulE4E4t7aM8jSce9z4UQBN1X1pW92AGoT4dcntNRX
kK7k6aZnagR+ST2LkgJN30q7sKE2tweWVdqyWwVbu2FW7oatS92dK3mcZtq9enIf
pdXhXro5EIgj4BrupySFzyxuFm7r6GR5j8VKM/g43BIh8hi8KbFzG+dHvQNwuJfp
FU5zS1+qNb35Baz/QvRt1T02udJTW1JHehkgfFYi7H2Lpj1MVKlGLvqKKnD6L1Dr
gc5dtc8Yduz3lu0eYxY9t3aRlS8UU19+hpxYq1DV3GPONiFYJt4D3ZSe6wjGuv6p
lWftf8QW5G43dRSdy3P5QbcNmlpTltyVmAQ2hk/tDLI9euxY9jdLC4Knx3cDcZp7
rKINtkXtwZyacXrRU0Ppa3Xryr/X+gfUSaJceOtcxOW1s2e2ipBS7LNa4dggXWBr
WWIKuBC6MB8er0GA2thPLOn+Lm9TFs6BqTuwytWPaLbWsp35D8BZnesNFr8KDM8N
Kxq1LAT4Syh6GnuRtHngK1SaNmL1oALnaF/4Kv6nGcMbuqGDaLNNw0xi10RQ2/KV
JdLVHTcBdn7YogU9ilNHHui9PhVbxp2ygfNWEmV0WcHhSkm2gVAWWB1A9lQLfHVZ
oMJTm5Uwwoogs8KrixZtm7lxCnKTRBnZkKm/3h0XVjvjySI5BwbXCft8w3wGf3rk
JXlEec83Y8ammpw6KZJzoq6mkrYpUcK/aGSSyRPI3QyoXwShf9fHzDIx+HmRYoge
akMSHQWVqT6433LuVy8QLaMiiKu1vt9+6jYNjyF6AhGLC5Rj/CpV55W6mfupWY35
Cj8KjRYvURPvdlnqKiHvr7T0ZVcim6R9/1+nFuN61mBPpU+KNPz//9NAicCEnCzm
Jfa+C1X8Cqg71zVqgcZU7JPXy5J+4LONDSoqD/aByX2VRn56c+yYD7bZQ8iM3jRL
glG0xsYGxgecwx0FsV+qQMUYcgVUDu00WE2C8tyYEhOPKaIQ8e1uOPx2QDBCmdgA
d5cMoWMMJ790QZPXFtTG9s6TmnDAFi4lz/BKzspdzXIVT11BAuZt+SBoFVinYBdw
VQHh4p5FP0fUvYsU1Ub07sPlEpXM64Ms9gCmu+8FyENk/OgduN8/8XfYb6Y5Aqqd
JliFDFR7CuBE0nhmu5GMhVGo3LhQL48cFfT0cvOu0NHmjhpa43kor9AvlINWhBV+
RTQ+x9oVpUAv7/n/1832c/kaEEfGV8oPvzBlf3cPv5s3SQwtyAFRiw2p4221IWfn
40GaBgS0kUjXm5qUEHEjivhv9LUy+P9vDZncC1x4qGtRrH8kiP1K4zF7mNUUpCKd
eumutCfnI4q2oTQknEYkriiHo4jPO3z3Y6/irigKuYU+RmAlZhRM2a0w2EQ1unn6
nvbkWqYGRHjlNGixnZftXTYHDHh9wdFUsfmLCHaZfAEwbMun8b/d3kmsGJiuHFl/
UXxCDfO/oDfQjy4ziahF6sj2c8Tlt2Dtn0pR/uoYqMOfJLZ8JXq3ldoP/23nTnGm
1Ro4DccByJJcpruGIova2cxwb+J+pJGxR2lBfj/tgC3AsIAUYe4aAdLdWXVPSxk7
GSq7OxAJNXWReBVDJWNgV21O9Ml12stTumOxMUveRd/gpJOF0oOdL6RxdZgqaF3n
54j7ezBQqbpvYUZMOSEurIcRPwpqNePw3RvrsBRMHsDYz7NJUVLJpNDk/8L6uRVj
L/2y0KVXjkJcGf2qDSL5OTbTy6CgFUG+KFYSBMT4dxMOgae+oY7MH5z6rx1ZLdfv
uuHhzx35287qlUmBq0zdNZGM4xZkGTeNY9RzKi81mCdSV2F6wW0pM6BqM+uaLqt5
qFb+D1E7I+tmra0PzRjEK30fWQ935eb3yo5zop4KE6e1IMhyjIScfCApen2I07ZP
opXf7pXV9Cc2QCXjdV5K9Tmgj/yhol1miivqTa8IfiJj21jjbihu9s0O+UtQgyo8
RlHgr7bXypu39FB3vLeArLB8uB743YNEU41EBcyltl0d6cxZ+7DZHTZRafJwOa6S
nFHt9FhbimTTTiPKc4p1sEZkdAW0W+T7daHQw1507DFxgzsRwUigNKZL622KvoJa
qtAhrRx4iH+gV/7jvEODVzRX8LN1//iR/wjYXkUkmwrmMK5q++3xLFiunNTG6ruo
nA8A4jvwmQYDyIRlgd32Ki7yzt75t6QAkiwnvl+bEGnaUa+JSweGECEjBcAHM7AP
d+yYEAEDCIWYZWKxcxSuamAG6JJxKjZ2oMBVukE6RsQtmJpAvNX0ByeX3CsbovY+
GEb9dGj+uIA4m9THeuxlpSO+0ehZx+X15zY/NIiTesRHLSn2InbX4cmajbBTX02J
Qzqbxxrt+l+a1N8SC7PDFoMnkNHyXCJWdaKvKEshLflmPdzwkWOzKLwpW5mpuNir
U6762ELcjOoZtYdZzKSS7ZQYf/A8tSN1UD5pYfG4KaGHsxbGTNSspA7HSa0E9Ybt
a6gWLf9Ol/gVmMDKq6bYHN5DHFw6gQyvvcipDKm1g3WVl0IJWFJRv1xaxb1IU8ta
ln4yhoUdERcVFpu02Tor8wMlG9YWmKVjwbMZ7GY8S9yyEoWuhm2Cb9/QuFtVCREW
F/I20F0DZ90rPCQO22t2fcaUnEOK9jWCDXmaIYi95MHGMmMuRj6pu+KNKgqqCOF/
9/usB6IfRhU7xEzWjtm8aDZ2tRb/Fn53yDeJE/ODkWImB1CR+KR2I3X9NLY2x/fx
QNBB8qg7ZJCGcGk1xLEJl5PcU+UxRv+NI8ln2WL9lOThOVwW8hmt0ZG0i2NZUZlE
CZlfJ/i4o6a43BDnghcoMhSzE2jvNRx3bM2LPVyXVxdR0E2C9Xe/cot7JTum5XvO
Esgx+6+u2RReMuyCaWkET0fHJvxsmLFANwwGs0dw6k6HBgnF0/+GTXOfDIY6Lt0K
Bk0+GpBK9ahRVn9k64UZ4F1qbvSiIUVkeVW4Cek3OyKfASTKMNTHyN2fbr4xLl87
y9MWVjI7IGr+M/1ENnH4wSGscsNWG6GITgvy1N8rp+OSboM4NXfD9QxN+G48vJaM
9iPQkjUnrUQD/vfs6sRiWhRHh/EPQe8M9qbrXhUS3BeTCfX/ki8zeTrcQNfcJJRv
ttcDGT1oP59mHvW10LvL64bAwR2H+uvoS/I8m7Qr76nVy6juBg49cQL3GWVE+FF0
Zv+S/RUFsv/U3ybAn+KDa13ulEr04xnOMJ6iDkSCMh0dWDkurNP4e/GQo4t3Xu8l
Oc8kz1rgtSSn/oJS5KUY1Pdp4qcBo3LimOMJvC7rCgCYVvlrKwsFoP/CrR9Rsr12
9v1D5VLdYoOWqQ+tMbCBdJL9vmcR9XNd1B2qMEAqOQyTRhvHkmtfRXkUZJ8fKKip
g1EABUE6nIXhvAd/HEcYSQA+mrWHZLa2I7gGsWvfMCu2JW4HHl2jTNrHS253EL+g
xX+/bG2z4fZKZjfQjEFSLI68Rz7loSXLaEVCY9YhlzVcUrZULgNOxD+tY1IZtdSM
xrwFe7xVGD5NTCkO/kZ+wrMwIGtXU9XwrGb7qrBVrNga3SsEbm/YIDJ44DyTz6w8
Ejlg9vSTDmBLH221roN3BDE1dA3aMO9FwvVl94cECXb/8eA4Qy3fIX0fplJv3Y3O
Dh9uYGsn6TLWesw8lpLbiS3ni+pPaTr04y2POZ2tDfOIxrEtl8lNuosCQ1oAReip
/gnptIJLeXj5v4K2KLrRFGanWlKh63ejaDCkbJvYRv8n51BgQloSu9hP4/zdfebS
lfrG6FhHaAtJjstT8QTGxqM+UdXJU4MkaIc/df7ydGyx6yXocv61bvse9UIeWmSI
9tDi60K5/VosyCYDxuaAlYwz5bp8UHNJLJEIYccg9CdgnWm+zEiq4QMBTNP6zIgA
Ycy5BKdoCfLOk2eZZkPM7a2vV6GmrXXdcqD7+ekRwaxkPeCz2k5e3zjLFB46RYLa
bNLKopsC2V3dFG83ntqTlFQnFgkLBEj8gXhzZw8T+WNjK2bCxHQGe9oVVZAjgQml
tzOfKL1/8cNSLXtxHP/ruE2Z/Z+juxoaJ6zkxe2s6lxGqQZeNgxCF9Cv1A/ivcZm
JGWRO1PjUR/3OcmM5p/lswDGbI2Am//2eCDnSSqKdAxJF5zwppHWq8u6wGyqforE
JWfijA7jgBMltP5d39FBeI+EA6YrMhrT8rbgGA+UVl62p7i242kR5ErOcmmc1twm
IoiKVxyP7BkHooPTS/Svhr3P2cTrFfwlmbl2sw+z7GmEnvrTo8kyUdoLZjaMhNbK
LBIrFPIQdf/TEZpE2XZPiVm2mcgQtdfKall/VmXW6lsNoCu/CVKMwblZqgR1du2x
ZaS3l3fOZFyqJyzP/p+qrOUw1YyT4ziAjlQCCRLAzU97YoeJHt2mA4QXBir4qmv+
hFEeyjEE6EAEFzXuBLyHzhYxWi75Ybam6jgeRxfIVigjTjbJ4lhuVKD5c/WCyHxV
3uM1sWiWJIFPkiSs4jwpXvzy9vGIlrMvt0RTGlKiGU6rb5btPb+O368y/lnoeRe/
H1h27vEMklPmScw0dW9JzLJf5D2/2M0LPITWD/9NxOdQObPp768dhfoT1RO0v8QQ
sXjClK2/qYnoxT+XG+Szitv2O8q3jxRVElZsIuNVY0CDrlObnj7qbVlQGixo63GP
LII3mcb4wPwp2mV7MFI6a/36mCh8H+fYv6iLYYDRyckhIffW361sV7m6qBd24v+E
eBGhZN9K6AyxeNK5iQXMi7foUxOq8KGLg4mWEyfUBta3fwZbs0OWcZfVm8la2jCD
VpGkPBn+dTrChlyJC2XMBoedML+V7qS2ZmsYxmSIlItI61vQMLS+MPRrUop5tYa6
lNGXOI4xGYs4xQeyjTIS9PD3bghe/LzJuUhKpUV120OvN8InCZZOdYwEscP4xWGv
Te6aF/5ucThFVlGCv+SQAs0dFe+BK8VzLpryVRYkUtO36rjlZ9v2vGNofsBLxxpk
j+rfvEI6TzotZJjSJ39rSwtpSydv0BkDGMj5IZTm3qUIUrFoPHkOfzo90SgH4pp+
ojwKEAfk4OCxYbN6URBTjggyeEAWXn5xCG73PQbgwJHpMWTL7LQhqJu/Tla5zMoW
DTdxXGxm5I62A4Y06WJGb0SbB74mCJ9QdO6Aa7EEKd+R8aEuYPKH24cerGKSJkHn
VmpJtTv3h8iEMQqAutYXGgPZFSbf8FeVvQIlxKHKXjmdM+tg5RLOuTla1S59R9vO
mfmIkhAXour1Ki76GOx/l2nPXkSHY173+ZAbKmVmoXcwPp0qwbXq6g/DdpaI3A9e
NIcQs8yLM1pZl1S9MRK2IcQObgOwsFqYHzPDQPQUwJzKxpbCOtZnomUiVe/Gmwuo
5MRhSsbTk0VrSPn4X98M1YhATWx94TEjAA0J5Fkf/4FxJaaoBaxewPGSvyHW2E2p
5rKRg27i1RTJ7G7zmk3R45ihvMt53moyWNi9lsxsSih65QFlQBx16hxeEvlhffDA
HFA6IFzvrK8TpQZOz64FpPbGbXgzpmh2pOILF+K+TzJmJHuRotfq6DHssWzkxez6
0JhzWn16m3Ixj+Zt9MkMYA5QDCvnJ2/g3Cj4C4haCkZNHgNNImcxMEAydpFj6IGD
vu/c0tEFokQxiZ4vrzFKD1HzvQcjyPLrXFAoBWkmK3o42+++OeXPP9zsDrz1ftQe
fg9lM0EuFKk7GYUMANL5nw9Hhn9CVpLN25dEhBZCEFRZPShiBvgk9u15T1+yANGP
90OcpkgMSobrA24Vv/K9np0j5sY0DCZTkqdrWGac6lquCKkqJQW1MGMDHVRo62lZ
CTj7KNMednoReKLL4zm+pGQdrhWcxGOyxXrdsAjUJyuY8ESbF/yYegV4E95bHVqi
d3J90x6JbKFSP5B9QMnVT2ws6lHusc2fIrbtPA6xwZs/zC5Nzka1vy2ijRqwphvU
VC42uaTX4dhq5xeuVCNCvw5Sk3sqzVA7oEezvsFvJX9os9+by29CEuVecXBXeCgl
nBQXFnWX8oc4syWbCcHXy3N7iRbE+b1b475OeyN5yAMtN6FmO0y1dHXcrUQ9V9Po
o7rvqEHxomFN1uyv414muDst1byTnZ2zDZnXjhtQPnn9tPG3p3j06dQjsTX8TuyQ
RfuThH6eX1WB/fv2JEYcPryDMXRri/4Woo2tItPblK/dXiAV2PsJkruH9eRIkaEY
mNzOUNB76UxIfTKJ6p2bN7TDpEluNJDNTIoufYdm5mrcQ8GrhAGF8kc/JxPS68S/
x5arDAR8J+AeD/4JDqG/84oRGoe0rE91VJBUXq4vQE/j1AUp6uxUYQu35dbsXORJ
8tFJivrsFt0hVclF3Li3dIKRC5QP6Un8VB5X1LMh+XPxPN03uEk6mw4W5a4dzAX/
JDJ2cvwDPLmmdWruNEFugROrEpCALXvEpYz3+vznQJFvFcE40GHUpSnJ4yfcpWOa
pRr59YaAEHrzLOcF4sB5EWQ00AiSbGbIkGc9jIcKRAo7CoN6OfrPt/RbOMFvWCoQ
EarwpHrE32DcaCwFGefwi3WCV8z2ukna+Wq1TarO9JpsUv1p+47cV/QMw5tL2/dR
JNs3c0H7RQwSrjteWInqfd9/As5W5va7eMxETZ5oX6GLqcFqk2a3sTuswcFVTns1
UZUoVtY4JJaNUwokO/xleeJ/TWNF5LFvbi+OcUVNsNYkjop34OEWR+Y0H1ceZKuc
iL4wS5/OeM12+vatDwfpUjdFiKdK+nQJHnybYVogDUK3xmHAjCmQwqb6W8Wswchn
ZeL7NzvnpzG/0+k2+EE8iNcOWTDqdbjlTydY360a+w5sZdvZ7G8OwnulnTO9tlvl
/ImhhgsdK327xHGYTn3YxTJJJp1SMWjrgMv97Hr4rTfpopYpu3MqN9ARkrvnCLRn
3sfKiCLmf2SkuagMxYOXiUJklBa+nZ/0+uEjyAvhfiOAZYkl4Y3IiL0+KMJBgNiq
Xew8COLHU8YSeEVhXjgQ3jfBrSfYuePEADw58xSjdg47HOrUi2Y4/Te6iFE9TLAp
A5Cv9zYJbdoPegFykm4LsRm9C888uo63BHX970ZxufFUUeKiaq6zjL+HZE+hk2YD
EdsWOayMGux47Y2ns5moX/5VxkDO7LBCIrVjlqCfL5SNyqWmCNb8FLveYIVIk9/s
RuFkZBTmJylwknuffBzUlA0qD19R6POVMKdSR5Ltolsk4edV0UTIRUZUNvIcigoC
uPXpMkATc42wUuv3jlIXiVrexp/yQkRtBLLZy6AWBIVi3yrQxG90J/NHbkOplG+w
iSg8qxc355vg7BEYxBZImlWiM9FirNhYfjO/cl+oVnCcj0dyptzpu3O7pcanpHD0
66dB78BcuzZOT1vIWW3LUhuT7NiLQeGm7wPHTUKMUFZX1mjQQcM4Q8IFghMf/ATN
RwNOIZU7crPWKbZjik1NRI+r0ZmGoV5DfCDeyeyEGKZmYbkEBRj+fmuzCjJTUear
gNrdNuew3XlA52Ke61M7hVatk09uk/UHTuAB8nRFM2OBDQ76EQ1Jc7mwQQhmYqCI
lZAnQXywhyb056DNt4F8W5MchqeUzYNhiM1Lvgo3X//Mtd/Hl6mev2TdVKiyIhAD
l9TEi7KLEtVk8dECQH5aIA2q0KMb0DV0ROBUVZ9dSHRmyyYWSFlOIteRBXurjUOA
bQWBU5RhUenKFXrKraIwmeqQPGwR+Q0CN1xOFF+jnUrksKApJMKj6cMWsHBd9+lh
VJcR1auGLyb7sZiDdU/21C05l7bvpwRZN3RXrkxvpUfcB5N5lLCtPXaxHrK6WxuC
lcuR6dC7BIDwxMjNWtpc5VDFyirLSotkU+ty7GQ8gO+rx4D3zig5YOgZH4931p2K
kHJYd3ehUanuWummgZJgqt3tyoaGopxceC2qSuOQ/VnQ96v3t2HKoCc/Hk394rFB
DIwL+bwgy64CIny5bNCtSFaUtty2j8Ej/z3gBlQjtVUTxrkQeBTnGSF9m/mFkrUZ
l2vuCwBPkY8gK2IN9yjhxogqeJ3J+J5+kkqxCmgQqiWR/cT4+t0XIrEFtpNDwgkc
4nJEpZc3IHDzf0b5hVmfbfNo3eEeiSDOTbTOmSk0Uy3A2TB2eN+jRaKJ0GZFnXar
5kQg4Dj0anOtF0pvODQlq+qBUX8ub84PEH6Z7cDIQOe75gxWDatbcy153Uq+OP36
ArBPh5SJHuJWhBngSdwZugxhs9csWs0ZQCYVDCxDeiWDQub1ClI+4mwdFM49nnP3
AnYZ8bNgtHOSZZZN11RZ3RSoEmvAl1N6anOQHv5R0DpPaE1MbLxJQlBcL7OYAvcr
2+Jcyuu/+BUFI1MvjyS0/tKmWETVJRXKEzmDQDxZ7BDLAr6MSoKrBbfZa4lMTK9f
wKINXgWYcyf0IuX9x9LaubkV8CZlXx57Bq64hD7tcbSP0NkidFOAEhbtxhNbRpfF
kz7+gavWzALV0rG3P5dIPLVE4pRPgal0T7XueyLdLKdTrU5YClD7YTLsqMheausZ
D5qpbzB5BF+ZqS3Wz7Qs2MW6OFdvhecqXVBs4a3gN96gynqooDPSK9Z0p7KIksRN
pSDWrIE89wULVqrNtl9UXgwn5p979Cd98tSHfGn7Yv1MiXI/C7iA6U//iVhMnoKv
2sSbGN8auOFNejJDTDo6xayB0iuj4A8lPgfIa0pQrwXnHvPV8v1GyMqG14LfQkV7
aIlw1C5clrcdgIuZtzipJX2EzBWCTUFv2drp57ZECVs7t6Ve8q0KmFqJ1tE/HZFJ
nQA+nmJ2KYeLZQunq+Zt++3YtAFmWM/rHHpUJ6LIdVGL2FQtk2bwmdr23LB/3gKe
d33UKqIV8xeiQiePKD/gTA9yz/jbITi6mvuKcmJhbxn8+n/yqLlS5hZlQqljc1pI
gtQWPXIaWxmjoD7FzIuDliMTeneN4+PPf3hEMRqqOKbNgfrXVaxSaTsmfrTrmijp
3O1p/wgtXvH2XZw8yIiHSc1dl5Zs936alHUM+jOWXRJlhVknomsFy2Am6Z0/s6FB
EXQFDzQS2hSgGcdX1n0mDZcA1Yy3jikaB3FsIchiWqdCizcLQxVEqFlT7nhvgbjD
/tBIr5RYpLY+jpkokoIOCRmlxi1cBsuEjoAPapzCQFToVaHug+lKoTHsRotEf18g
l7lGQ3WOdJgQ5bl0H9bGkWRyZapIe82LpbJ0WvJf6PaUVncWk9hfG7h8fN+ILmiR
ojQQBfEHTColKKZvhIx00Mt8oAjKjlYQvznLEwOJuBaOdfNoHZCEleFHZos5LDIl
U1qNXPaprv0sJ7Chs1B5T3cyW7BxrDBJ5cysf5MP9Egq87taGozmHboQlLj2s4A+
cFAfuIoo657SKmCxLR/D+zazQQCJqA9kUs+e1FUZZhTRrNKleLX3JG1oRPJnK77o
xGZQt8tsnNSx2DZjXqrqf0chWgdryFcWVVSGCLUKMX0MdE0YakrIgu54ncBpI9Ue
oqj8sAKHfaCZY+kMqtjd2wtfSSYimjBmBL5aI1/8XZII6NyimlU4g0ijxa84+yUN
+Dduq/Q8xq6Ow8FOorapIOItz62LIuxXEcryFuGv331n9su5IIb+MjZ/O6i29Kyq
fHlgp20ccfsy1XnQws+cBU0i+6mokQJ5A+L1AB6azYihAfdV5SrqI566FlBChbiO
5b5R2QUser/w2PwyrjeQstud2uVYT/3lFasQqCVb0lT2crqkGKw4ESflGlFdRGxu
3aAkTFAROQk6+ar6VFO5bOck97Qbyh/LL4gKTZgjdinz01+DjZsz+lucCX/qGcl9
r6ANNN9rgB11Pg1q+wT6qOQ0Xe1q9UTKejNlV+MGuN5nSZrgVWY/dgzkQimP8yxr
wvdPlJs0R8V3d5PMX/YBuMe9E+59nUlHsvR54FCN9CNjw2U1hBN2b+Tm1RiL4IKl
UWfi6oCX/0Cp3vsEU+tfXk8Cq4aSH534dCbgmrAk8V9EpzyzUshOi/SdXMO1I/8N
X0Veg5nn3JoQ1XtKa+pQJIfFPj1cQcWs6zKjoFJ66O88X8vFHxvjSngCKDapZdW8
EOf6OWGq5lC+VAXUrRiOIzDZPavPdiZ3QnxpxFkE7alGNVdTf+/8wUlg4/HNeS4H
g/aExpvlQ7Rmf/bzIBYHd3eek7MCSmnRh+gM7JNaSQpmzloPMW8QOUm+OcgMfLLH
aga7RzEl9yzlqSBAT7T0hA7AGnd3mGBj+dlg67szXicrEpDQenp/8G/tX1kveccT
LTC/6Skrdke9iV61F7SvRwXF0lZvMcB701JP1JJxaOboAN5hU8A4DD4RRH9EwejP
fAGUTS/9HLaCvwdqdEkq0199GpgZj7Z3uasyZPKpxfCliqa0dIpnTLx1cr6UrC6g
ixGWpfTxWFbswZSnUh3KjTnm3LLNMHo1ujUZREwIu7nKL0vpCoZ+SgfFKT8xtl67
wj1HGxFN7ysThpdhmEhVDJpi2aoM7M3KXc5BcjVBBphg0Hc3fbieBoNKImigfMXC
pLLQGu7F//Ve/JcXqhYEEscSTMiKdnJ3yUpkvj94DzuAoFWebFTBVZrrDHKKva2E
2eCOkXURECpDK36T3iQ39qgroSLLXakRgZcw3/oxV2BiEdOiCY0U7srlCkIOHO8j
FDxMKT+5Lrl1Bsw84HjN5LFuuwFRUORzW1TFOcnglyu3K5nn3ah1Ddweij1kt7ot
HBRCS3zfVcAizrk+zlKzqaEcEb7hIAVd2OO6b8IUZ1+QZY/jwovXe5g1WNcRZYgT
L5V8ecwPHwlr2hhMdlXYtx78Uqslz9HUZW81gqx5XVbWa4F8WZ3jwgSXqiH5WKZG
1SywZuvkUSPI86dc/PtW4dGbAUtOEeuvGQjCPJTnF3xpFWMyz/w2tqO77KFl/JGO
I7u7pQHNEeUUWsKfGjG6wlNLDNdP0PZg9cMy4XJj35msV/qoEWX05bKNBsDeEaMO
7mvGTjzxfbJCwPLIB347Ah9zCQ1gDux1Tk3WwYVH+8Es9LawohHccWWK1teIB4Q2
bI/qBjzENf3YN6eZe9Rd0QdYALFRw1Kd+y37cOaItBf+5NxmwzYGiWOEJ1PVpEIa
P8WcztaLDcfo1V/L8Ex3miqdU1Dn/YHFbqKi1epVHZ2G9F3PRUwBprTKkk0nyA7R
uF6vWgDL/mPZKWAdjQaYZsnzuQoOfNHKBkMQgJraYZ5bq9rph1+a5bffjxMpXfNl
BOqTXaajFrvMiVKXMGXT8viMMQAJuksTmwqOV6OXkUdIvKiIaVNhbghdEk/vtOpG
LGM4Lj3ShxztVwuiAWjTBhkQQwN94n0sDYxOurQjx9ddEnqldUrtNUcMOlI7ROpN
hnJ2ieIDZiPWH6Nzd97jDG2dMxh52PJSCEmyWco3EXuY0l82L5hEVX5QOid9U9+0
jOncMPay+7W3EXXS15z/Ogeiur3+lhklKFNLo8/p51GzXw09X8YC81uB3tsINyZw
n5LBXp/LJOPxA16OjqzQj1BFg3SLEtLmU3ddykT4KeRMsgvp+wiYbMJKwyGrhfJh
ki2bQV4SBv6+FZiRVbhxRmF6n/P3OdPPKREfFJkDhtm2/xQt9IpqWCp+JOJs6Opo
PX1l7cRSSmT8JbN13HDG+elgAdg5548mVSeUZUqGLSHEtoArCMb0xcQ7Juf6FbK0
pHzYJD69ZJC00Ixu3oTBgcqX4wAIdFtNl4ejBipjMNdc8tDPpOcCZDyQ24VeyJO4
R/AvNPlU21qN3D0SsIpJ2UalPIVz51a51480kjBlS32hcerAjmUmqG86B8B+4uh9
/H4mQgZhaDFa0V++Du/xomz1HoHTVvIH1CFGjLoMNZgh2OCOpoLmybfozVWCfdQ5
4YktyL651apZE34LrswQT9vXyUd9htAgncBpMrT0e46/GgkdBaRt/z0pPHQYnhwS
/UXuh9rV+i1cq+ckzjc+JGc5amqSvrwOdIM3N6bDfCcOPfQlWb9FDMJsYc2k/lz1
+RXekvXKBQM7zQbTclXpc20tdYw1wk7GGTgyBmUH0RwzfO1d+AAkf/d/jbUStRZa
k+cqq81sG4WPSrMmVxwfjuTfdb/WIVyl9SmqbPSEWDVL/8Ugj9lglbmGQRR4bCe8
TxxH7U3PR9XXMSiIv59k8pvXS61ufD2ajDgfqXGRqIOISpKZrKh3awlmpRq3jEsd
gJL6E3yGH8OGuW3CFXapa3+S1ViDPgKXfEYvMOBxZkxoFucOuQuWvG9gMdiq3LmI
iAG3JyD5ncMF4YgTvBfvxNfWtW79fGMXrJ+Cr4NzlrwwuL9oJzQTc+e5LQqtno+Q
T3tGfxkg7PAN+Jk4k7wYeFq+aQIFt6QfPazCabZU9dlMJ9kJ4jTiTHFgnJcsobed
Nt2GpGDKK5S6LtmjMY39OHQRlHZdyHaDgPih3ecJyscSd4LZ4IfC8Ysq51UHfc5x
Q1k3n2739viDg5RWuKDJQWIXbatvK7c0c0Pfa5jD/txtU03QLrG6sbIrL9lwHvZW
SpD7tkJ6pDxJwSMfDi7BhbGIoo0b7NrBduU9ue41IGZhULc7WWnr48XO7PjOhDPe
RGd86/P3Bd9JQjsyxdHan2ijLmEziPNAaGjKtX1ef/K4Y0Q36cq09+4t9UUt524z
9K/TXNWhLRbQZKkLXv9bP5KU9+EWYFdlxhbPS8VzhbwvmL17mmg0WUCYpZKr6blj
+YvrvXCgbXWzfPzH8lUF5lEHid9F2SOtHl/C2Q6JNjBTKk6yfBrOgwnAd7F3O9Ih
APryPMS7GHvtoJuccIjs6HgqOphLmLXXqUkmjqvbovz6VFOIf6gTVg62dlEhoujf
j0no9/rsghZ1E+Q5fwTz9dtXgX5Jzk6sHpXQcKK+64m36R0ypXn8DDYgkjEgw035
jp7Lj9ajkOjkoUA1806wSQl0OX/VkaSQkYCUCSNCBfAthvqKaCGkQxdpH/VHjcx+
BZLZFY+Nyjp/LnandFJbnG9IQPLa5zHAylQeCjVaPtBMzenKKzMj4wuPOzh24jEG
bSCpl46UyGmG2T+uClcHzyEjgiL3fE3Rw/XijAKwZkulVfKo7uRDoJwOPTW1RUui
7zXzBI6skBpiwYPVIjJ2OYprb6D15fsT2vPNGI7hnhgIGiNEvcPV4CAyuPE4PJHg
r1x85APSt8quYo0o+5PSpXGvQQ9+ZWZLoNeMT5iqXeG2udxkCyqpjl1GD+2lIapd
RNIdUYCXvKZrgaakLVwdQNNzDmXVWAE6zP8lKbRZwy578PJmpkTOnVzSd2CNFDIr
DU9ZMxSS0loUj8buJWSadwYx0/Yl3oaW88FfXoOmfN531LWTj0hQjk5fg8EppJD9
AYZg5dFpbq8sti+uKPLCJN2eic4EirJjbCalXupVI9KWK5tL/AtgJPE2MCsjjjrJ
PFo1545Y/E5JvgGNqECZOVWJpBXtrz0wJdhlBb71s4LtACljHzDXWAsZ4ToDPvmH
HgnxXu63Z5ORbLORnYq4Hz97Nfq/V6DLbBIaLl8fgzH1+U9Kncz59jgnxyms3rKV
KEMjDIrY3B6O/gwUd5PEHVBPiwyILiM/4G2a4j0E9Pj2y9pY2zQ7t7yw3FGC+eDy
9187D6s4Pel3JjIVJWoxANSIgBJK5tJZdszTJEx7/He56LnOuZFSHAeE4Wtej5oj
+8Pn/IpkkslgwA5WyhI+4Be8aLJ77IBDAV6H7ZoMBza3VfU0hRxD9fslXz/SinPn
Te9xyFSWkaoJ4BQ+/QGsB7u/kPXkN39+npHn7inxYVuA5a1tYBskLrrNmfC15lSN
B+Vl8eUWwRXrNtaMc6V2WaqqE96RX3wU8COvf3z4AW0kCdOr+aEk6eAfCPMO/1UX
1NqQAqJN6I9s7gj5IFh3boG1LhturldAB4vePIKUHQGuo7QvxpBt0nF0dhfHqJr7
FVWIQDc+Lb4nXoKrWiNfiROR7HMBCqSZdYZohgn4bhUlW/2Yh+erTblHmL8eovW6
VHV/JOQh5JBb14en+Ge2YcYzIVEExM6q3Nq0dzZQ1tRn2OzZ6A182GRqP/9zjPh2
pdymQBglA9y6JLLPjtGQ7UIHJ3EXHPZRpamYvIKMTlHjEB7qjqKNGdDiFxFJrMcT
jQSRjzjpkwKL/i7RGpt7748P9wyaqObOOHRwwNJNVpad4Ca1zblmkjJ6XemEUum0
wXC/RpktJnS/D7Q8s5NOY92prVfQD4RY/pag0n8JS8f8WksCe/tXpc+OsjYImqfz
4fyTEV4aottrOWh4B2p1iutExzG5GV5asYRK2ZhB6oJQ68dmry3FsXttW8CA9VLo
akYP1LncUCQqIYWQNcml+rZVgvlutyg9GIqDq90ZNRMkSSoqdOIJzfENnZ2xo7zn
kX2dXyKK5Emxd6QuGyvX5bPlgAu2gN72HoieNDYbD9rspSfsgFHBaQZa6vkRR5yZ
NbV9GMz7WoNCBWXHyLWRsLQABl3krG+rFNa3CFUrj+13BEma4QembMU4wz4+tQ6T
JtP7/mKqgpeYonFa0Pfrxmu+BY61K8/yssqQlv3zsUyKGwZiDH6GNnKz/KuSLuni
PVkycGhnCBhaktFOuHTwWl2s5ybx9oMkjuZi7g0jaebtderdQu8tGDfrwVRtxqk8
sKqmOtFvhjPoCLJW5gkzx3h43xmCTd6gUeFh+bMAk3sx8keOn/jJoQQeeMbMkkLM
nscsZT+aSbIW6y1yLNoK/gZ2nVGF0z+jbxZKPL++P3PluP6XtAKBVeXZuiyRwVFw
zJWZy508ysg2FXoAbRQPRdukx6bBP3mWXUc0iCnnGz/NJdgLQPzkAXkrfJR5s1Ue
cTq6S6BGYUlh/CorZIfcWYyJpnWuHQ1JNW21ClfPYUOATyAHHxCw2bwwQNX9WOuX
GMDnWJlw/RZbZtlR3Kngz5z+F0r456Yz08UVzUxWEgbD3kFjdjUY0iErITQjVxlj
bz8rezpv7J/GfzOaK4htd/JxQt6AFQAett6d/CFpLfUpIfldY2QJkUy5LTUXZAuE
HhOB2E6qfCB+ZtHoMQgg1H3KgsJIoMzGGWpjmJ3qSPiB9FmlYD5mvFx6ZcT/z43i
ffxvksf1ysko/6OlyHVUPcufhu0C8/Vprb8pq5Pt5PIb4+7FJOOrBlz75zKwin4W
HsPbUNLC8vGVwI9hRviQI/7m+luQnA+lyr8h167azEQmnJISfWQmBk3xxL/L23F1
7vIsz3Wowy/c2sPclfWiC27Vq7VW9NRq5Sdd/QxZbs/Qam9t9WFhoZYzXQWAgHh0
ayiNl+3gCUrrbqwlpc+KFIga7pgEJAUNRLXrkFg2S6sDRy/OHp1olJF963P8wCfB
SiD8OGO2I4Bp9qAtB//s5BjZFUp9Sv05lm4EHDpx9N83BOEs+XCt9ihn8bVCKszV
vsFhbkMc2fVQ5G8z+G1UBUlhiYZxVngwbXakNc5wq6zc12xDDX4ZiH2FnYbk96Pm
UAEgr66GpT/IL/LmRTIOdVbOfc4hpOnucwo9dIP6BVF5t7wvPLeSxi2/Sa92N3TK
+P0eDECi6BiYk9a/M1VWYhpvy/yJmcV+VInER8aKX0rEDMu97Uf9fSnuYu9jKuvy
7SNQ98vaYXpshs5iBc3BK0KsphRYpm1fUW1j+X0P5PfY7mzd3jqKVSZQENLyzv4n
cbTLmXqzRN8Z4WYBbyw2qwkMHeEhcT0ldp4pqwVW+tOIsmuhXJfw+By1fCCCIAng
0l2Hv/AiFlhuOg8rBZsBW/RSmPPVVmriKvgha/Aq+hQRT8p1dRW3YdjbRy8RT8b6
Ld9mUMNDNjbYQlRbBwWfBra/hiSAuFKjpUdExeSEIFvylFLzPN606lIi2OSU0nfm
IBPAkf5YcMv+j2V4KOtvn+caOdagZsJ7ZbpyWHmA6SXdNqYX2iOlf4hFndOZchVA
rLVOo0bPJElLMHuskFEerkeS05sPjyyFIU0MYIaGXbkjO6UrKANJ55BQaopWicQb
19MCjSTqeUpO3kSFaLO0Vy35UAghm9fC+t9hvtK0xtNlLTBXydO2hOo01zanq/rf
N8jKwv6Js0v5l3/Q+/7RWfNhl/GqMSn1St9CAdIx+Nd7cS9sFzqD2erKKcbcWvh8
eO2ASsSOQW//Mu9DwLqFSPrmCf7cM85njpBOwYHWqY040ZikxbYBRGIfSMnPXd2q
42UQr28aU43suOJ9HBRMWDbNyMZJeVJMpbiObELN21KUsulAeTOeaOEcuJeyJ3al
sKM0pqE8CpaLhuVd19zzN6ijqKy3atxi5FFybK7HkdAlA6giuW5FGqVCNnGdvylC
2UtQhMMpdYn/9W2s66fm21UXpX5EJruf4pUGWdk+SqNhZglQLNOrYkGANvm/zIe9
oTi7r0SIwpJYEttWpETepJXRyPNrYloIhVxB+K1eDaXQg7TdWGIDeZout5FZarP0
6matgH8mYefA8iIVe9g996GKqnO7jcMVSfWXZoDyx5TfdIlz9oq0hOf/1X3F1DpL
+FWPwGx8Vqr24O1hhaRGpek5qKKHJYTS7jUPz83EtSx6I3VDtFpYTxfCnlbp4Djh
Y/2v3mdFZmmCexNARMaf8eKn92LhTtaw9WQvjUPRU+5PaK0AtbT0hpe6+O1eOdu3
GcbRw89rjUbyIn6wRQdbuDGL5KA6qM0xMn3iIYwnIbSK2w49rYY3EDrCssVXjjyf
oaMtXmqjmWlsr6LG/yomF1VuKku2wc7k5fSwr6kWXUGXcS+cl3a3z5zBppRvLJHj
8Q+uyP8bCRXjBdcQ7d7AMxFs9TcPHdO4sC/PWMKbyeQR8KFH2xXkqr/vrTrNhTc+
9y0cO6PD/UIIacKvw3q5zDF46Ca/c9TZUHzZJGSVhMjWGyp2woopZImvhkno+KWo
nN2JEHx4O6LXpWBgMC7wglMNfcA8aLMbaAq7yBXsk4tWVvkwPLew0yECv5ssfivk
HJspPBThFVtQk8dnIUEe/rxKQ7xPUZ0taZSAljq4AHj16F6LFf8YzVD57HeBfXMY
U5CDolLzomXDyFcK/czRM3Phv45DPqfFhzCyIT2FQdcTZ2oe25YqeeQEKtLq4Vsz
bq3+r2P0MdeJCWeJue/49IyrpGSrcI4E1tMApz6fRMYlOI3Wb81NlaOvmHviIsv+
jqsY8hvTEN93ABr8P7BFPeL9d2qqCbwuXE0LrYFS5GXvsdDqkxiCE/nGtJizCJuV
tAY0ceAkkLpto089p5WeObLKSZoPhHXj3A9+p0lR9kXP0Kt+ka3VaxXqZ307lx5q
YERcWlSIa8HWx5YuHBem2dIR/GLH8c7+TeMtPN5v7gYtr/f/2XItmGN7Dk29kJPZ
b5Flzg1FqBcZXM3hIbSir2E5440qk8Gn1WXPQ6m0FvH6Qf68mfsrG0UcAGO8EtJb
11kTd/Fu4KJ2p6i1SjwuJ2Rs5SMI+SNBHGksIOTpzwzsslmPz0+EM8dz0cx3Hrh7
XMjRb3A5lbC4sxkm+IOEa5QBsevyB/l/7iJ2DjOoL3mtoubP+J9Pk91OgmrpoPz4
VQILkO7u9cNY9LlVgsDF0rtIaQrY3twCwJupGE3P4ke8d+zM/aUw3s2+9bZwq5bX
tNADyt5IYvvyu/zMXxFVnG/5BJ8f7R15ZV0VTKftYPXezrUfR3PIGWhZgX2zMM81
txs+IFJ/TIz8Q3V4yQoQVL7DFuINwi9VNMBE5nYUMKIM5PMY9SSaouSnQ9n0LAQO
Udua2U5zmvUwa1Aihmeytta87837ehJ/E1uJQq8t2HYOTBgkN9PEgmPPAN7MOC9O
7UbrKnmLkuBul9QjsqrUKoDnCJwAby477r4rQlJtPyfAsA7iZx8jrA8o0F+2xSJb
vJjaZhK9O20CW7Xs59u5ZUaMRs9mUTa/wo1pdl+OZ6E3JO5aQJBPA/gqNzsW1drH
RI2ROyovsqkjfRlAdtVpsOcqAG2CxhcZ7Ty+KM7ay6IFlZ6davHI/I+7NIxJ2rS6
yW2hVXd/T2J/DXZTn2GkmIxyf2CfVjKU26y8sLAjcz9YL9kUHr+cvf4occikePPM
VX6lcSyJ0jPBykoRNCTmn19Ik71UVrOjn3Vz8nZvp5tg1fltXOFfgqvXYXusRLTj
NZB3vcwdb9kQLlNTgfgYyfAoKSx1Tl1wz9RxUxgjBCN+v4ynL877HePhWsaznl/e
U8MR5gVUK2yUDibLdCHNDTl44I3+Z+vdjurm7hA91lG82YONVE82ZptLxIUtW2Nx
EQQxqjnr0MeP/zWLZVRuP2lRe65MFpxXMxwNPL2RXNffKO04vfKaHVz/0MH5i6/k
Gjjdn4ua1m7ZTIuA++UhFk09fdZ655wCFHhy3ndhiL1AVHmlFBqSuV4SI5qH2IL0
MLvAEOG5BALk7ShCBjlDeQgmKuj7WeW46qILlXDFP1gpP1uDo6xnhUXx/mCIVfEL
hj4/Tn1wzt4J05ZIjn3LqTNxclR+zxm6PiheGNYEmOFSGmilM/73voAIt33LVtED
uty0O1U2cyYFbrUM32n8oLUnXwT7ULaUx6fhD7JIn1ywM30CU5Epy+19KVIuwk+M
vG2Nob30uN1lHO8mt9abueGv+qawt5tq/tOodC2kMLlk+AAXAmOyZpZPeiYQujAr
r3wR3YOYYKOUiwj0SzwQQ/S5SLrFwNvFwzp6RFft7dcVB2tcWm0PEtJ0gJYFyMPN
rgPQfj2ixd+H38YERM2YaZohWhBbfxEcTHRdmuPBEgfMfd7XJCteooonh0q2Z1Iy
xV1FTMKR9epMVaGy/mtswlyl8SVcLCN06p4G2PLlXQo2+6qoJbrg6i20gT3AOIb3
SWLZ20gK8NiY9Lsn3sKraIGoLlw+wqfB9stKAvTxkpA73pvMHwu9WbMtg4ZjSDab
QsGRsVmZQ76xo+cwy5QkEXLYQIWC89UzRI8/RkD+IbH6tGiklToQiwkvDdS4ZwD7
HI8eHU0wpyceKUOLgZx46eY0B4gqHgI+82GiZgRobc02Hhc+BmVObsMmDZs+hxm9
hFMXvLAUkqHyS7UKRAMBfAz+339NmrZD4U4qEHxZn4rxP3hDjKnzsNKI12oRHj4e
PcS/K2aFQ1V51JGpdJhMYbyLl1ku9YBzadgZBwvUstsh6ObbbgHc6PHU0saYkhsu
ljAMnTJQ5NgketqhpwmdAQ7hOgkMoytkEoKyhzbYKdrU+U+uqEuUneeM3qoGw4oK
qxf+5sfwRq91gqIcFVEFN+FSLn9mkQO8eacx9YnR9i1WaKrr4WE8AgopQhaFT7qg
jzTyE8IkpC5uLtoPxcsAcFaimr/QSow/SXlxORWBdqd9HMROO2eh16yi3V3TcUpR
nT4KKFmdqFqX0SVuSmuBbM+S3h9q5cT9Luxq2eUrfubLnlcAvuQlqrhkbxB/nhbE
BYeuK60W5aOhDFV/6Irmb8LaEIyNJDwlvbPyx0e+ljSxuZ1ZQOMHhbUZ/bf13Ikr
6r66lBRfpoJsYLYh8o7YelqqfPI3RFdSTycTM2NPB8xiZ9I4imWq0gWi5TjNVelp
ZNm08mggi3/W5UkKnvXO4oUudzZVharPshqWt+9iqHYfxkg9uoPOC7BByy8mTXWK
ckz0yOzswAJ0n960OjCgAalUOEQ+FKnrZE5ytfIsts93o1wN13i2xHBwRCiq0od9
82+M7l0Qt0wnYXiszGnHSvA+fiP2EBwzKHIiMyhSLz/dPXMRceswAJm3q1C9FNnB
+r5drOowdWybGjUGyKfGMmpP9u41uCA6IIFyz8K9SOFuuB/lVVOMIziI3hEuqDTv
teYn++wQSD2qW1HYugK8nUpGfinsA1hs6gFBlDpAsTjoL3TRo27uH2efVhlE71Qz
357mDYD+JKmcfJAJFeiQRBcwitrH4SkmyqXjyr946zvYXSmikj70sYwYfv8SW50T
e3Z43H/QftUGNW7x2uivipWjQdgBLQTEET+uTv4UI5MsyHjdYif/X5vDkMpaLB9B
sf8xiikBB98Tt65DuyL9u7oAlmRxO1g9qR6jxV5wdlTQo3Mjw3OQ3+hWdQWOoEIx
JRat3Rp0cWeVQCqgbFrkm1zS9B/ude0HjiibnpFOtitYqFzNefIzwCli1Q9R8M0p
L5ZJG58NSJauDr9ydQLYZNq+FusvSGZbdxrZ6awrjLE8C0y6b/C2Wf9NzXpmRyyu
LsoTKkqGQJ7zIasUVZ176FAnsCBHysVcydk/BlfTBc3xOG4FPPDu5BDvIyP4j3Bt
661ow4ABkJR3GOr9gkWxVYlHOCtressiU8o2PiiQixBzMjIRbP5RP7T9r/9qJdvH
TMSgQvFOqGrK3OmzJAiEMFNak17osovau1FKQ3wQfWA/LQ8/RcnSNOTBwk0wO+Zy
qdWGZ1S5gTwbkCqEvvEHCANwnFiSUVF89/eNkOhm3RYOf7snJWVvie7dIgLXluhf
wieas24O0GD306idm3rgzUewjSzINO88esUJzilDbvdWgM+lQp2Q2XkCqX78kqZj
VSY7H4qoqBCrgve5jYxEAvFX2MSMuIsGx3+6EuTPsMr89oW5TzrD4VCTQAtiv7Sl
RzaBL3slxddytLKdc2tV+aApQoAhgTuhrM6Spy47TAN9i4buMCvEd+FDSzofSGy9
Ue/yHNAX9eGsBfg1Ip9MoYkO4lMzgb92UOPekg39CHwFN5IWAz57gTCAAjJewfHW
NTf7oDbdrTQ4JjFGyNOHc3vBXNp0neYp3H/w/XmRVS9a4U5P3/UtyjfJDZ3hDKzd
QVZClPCoWQhkQ3wuj4w8VYGC3CSLT66LpJZb+6RJZqyImtk3CoxcVqCFLREsft4n
C0MpuM74JsfDupo6eGcm5rgM++CTjFU8wQ4xkAeODh4sBIexFPqnirITxP8KPopN
GiG8AlmAl2AUmfvaFh5ST1xVMpc87+/GGuTw8fb5A1Rl2ZDPYYC+5OKGyOKUDCKV
vbHWMeAyqrCRrKE/Sl1XQ/cnyZSDpOyQsOdHv7BU5dm7DH1SruD/TjpFIQ4UpIuj
4L+5iFrchtMqkRFviyuEPSHOKwSyxU2brz6nQm7+aL/MQWSj7e+Uad3W1++RvRnw
WIIX7JbB/U9Q3lzLF8nXsU/UFkosxgwfyg+0bkSe1T/E/Ttj2rCQeZWMJnt/3AUE
jFOE1YlbEllPLE99D7hGUVibQgzP/MUcJrgz4QKneRREe9w/lDGyoqhvxl+2cmsv
aZycjNc4di8rk092HxH1prA/053K3lIQtD8KYuOh0kwyhWbGe/0Zuukk52sdx4kh
w2kVmvSHHtyHZ8xfEnqRDlyhXBMggD8gy5UEN/OJjLttnTDSyvPySSx0hrrI72os
6EIuxtLGfXE9a2zpnhECNhTEmdNxh0XapdP4wP4DsBpX1mdJrpevLnTQ5udx0Cxq
BAmQD1vAKe2DsLMmALB6DMdgY9v5QWmjrxgvrZnpLSqIjykgCshc/Sj9jyI0z6yk
818bRxYwuRaKJku4yA/bGMRcVdieu3edW+GcysiCruMkDjRxuXgfGd5dLjItUC4T
ODsabwvNslp55qy66Fnx3hxTDKAF9XKJmPk4vYkeDQpR2i7T223+SBByj/4IFzAC
RnJbQn8nfhyxyObsTpKESeuPoUsGN8gAFLBah3DGAWSb+8CmFNsl6m6Trtg4EtuR
q1TkO2OqmQPfFhuB759R8kxRUlvV8kdZkmmw3B7qk63cDhNVO1FWecDv9NCt0CML
X5qp+sH16HNLILPU2ljPhFbZ+6zoFx7y2EOtYJvev2M1KC2/ncLHGZsMcoltnDH4
FHrwDH5BROewvDhaOUnrKxz5y2klwaAUzKxtFPfBKbSw4ECNJTFAI8DmVWZ2GjIq
2u56WNkT4cMAaqrNxUcom9iHdttfNMHqafRZm/bjq2tyF93jN6M/wjwXLOyQSN+C
ixZHz3zPLjZlPCfOnnXqLdkKU8/sZ6TN+wwFdaaKflG+9dyoRysc1K1GoLYlQkXn
N+5NFJsohF+khPE60vbYJKyS6fmUmMXe95Dg+uu4vzOQStmD1GdHr3EjhKJLskzF
qtjp1TUPvm4d+C8uTsFdJLnBvEGOPpUN2FCOfmb62P8YUL8MWomaUQBDI/DX+hJk
FcGEMM5KxG9GwJ5QbPMHnpjprvHl4o1mFHkgQ10KsMqBkepB3uw+rccJJlOxkJTv
rkX5MPnuWRMLM9sadFfvmURXYd+IBFG7egdJ8HxFb2MdebpeXUP4HDgOewi4caRE
Gh6nqr+DJHtxNlT4l4iFgwE+CxvHGReGSm2ibvzpo19ebyCRK0ua65StaE9mtJ5a
iWr8DYwU3gMAZxBl+C6R+uZeqeUMer89RY10b8ClOp9goieVP/VUfpjBHFk35whW
cv9aJ/Nt6RZLohMrBCOa5zVKS0ChhfKVEoYIuuWeQYTom4hsf0k4n8HBebZlyyF+
rCKjXDManm1IgGq2XvN783FIeIQfbuPg0xND7XeZpZn2uwcDJx2LRHBQqoY60OZp
tt5xPTJGulimV1s1YQLut9lW92B5NZMGUFiRIRyK+1bqYQztRsLB/nxdJ7j7CH26
UM04CpJcwF5oohxz0Uj/kn2W/Zsjn0egGofRYRw3fT+nSBNeiueVnjY2X4Uiw2kK
aGgE+3SOZZ4uubsCNABiV2WCkYxiVhCS4z30gKSRoRyeLNxQRAwn3UzF2FYcc9CI
2XouDxwQpEuMowdH8Gf/y5pS81vmUu+ijhy9g5AahUwUocWu4yoSPMv3Yb6WfmKP
WXZrnU7Cx2gl7APYNLjNgvNrqLBxMz8iM5CGXoCynL4Gdlqx6QQvaXUXBuehv1Fo
/38vY/7a8yKO9DcttX5CO3xchjiYaueMWedya1G4bkk4GjyNn4MmhaeAuy5wzdKS
06b1r1ypLHRgAyIRaAUXdcq3XGJa9UW7AbosjezfFEO/35fdMR+t2xaw4SyJioR2
V9GHI1SOUU4hCOV3A8ZtbZ0sgbtX/MwHsDvpoCBYArkUsTXr1yUJXcTeR8v4dqtk
5JTUuvyohjfupUlv0WH+fCY9wF2Yi1SYFiNqfx8BCLltHWH6bS2ES9u+YPkPb1/b
A7DzLc5QkHOU6pKKhljzEhd0HjSldZZVUOEJQic5g61v7oOx6mJelzuaZRuI1HT0
hcuEkbR3hL6X9YeDR//KGjFF+GlJPUpGVZxf8m9OohvdVUj1oImheeLJjju6QqhN
p6ifQxtRN/UBOSXE6tDpilk6uxLBedaNEQEJcH0VMWW3+JF52++3lewuX0Ptd6WX
aNMVr9oBMwhDBg7m9+3TnyscENWaR53rJttaVQX/whw03CC0YMapWZqD6Oy7dSjh
VZD0iCTVZ7QzM62MiUHhwGTtU1+f2uj/SqF0NRikP79lPVlH++6371rU7/74/kSm
JzyAEKdqB0Ho/BfiMDbUXWxSGjzpUHU/obLUl+Wg9hYYZyHuqrN7h0carjd4Rb1b
vk+cSHfFGN3U7vVzlBugTdXhcnnAdERnB60TrCgGjjycyH6lO/5QpCGxWL/asiTq
eAFZ720XMJcDJLT8VAFR/wCAvo4D4l5eE/0lowhwm50D61pD0yt4aTyWa4wdl/MU
IRPtkruIv0/VLap0FmMMa059V/1AKYbfQi2PModPa06ru4Youdv948pj83YHbwxK
Sm0I8gKp1eY6vLxnKfhHf8FYI/qd5NzkGh3pXH8HmH6oVFHLBmF2g0VdKqeGtZkU
I8wvoGysQufHfyeAIXGx9f/vN8AaI30VtK3akaVl+gE+IEqs8Lyl3C4WIDpYLSiZ
XRHrYNg8OtNhOcIXtY2PoJLaBcMnjUPAf+izd+Yu/1LdphAGOArEO+9Bkg/ZiCu3
sR56X/doyNgpNuQ11TML1OQ7I53OjjP05jUw2J10esUuFK6RA33k8XhaH/mzy0Cs
LTY8oGP9/bn/I2U6V8kumXl+70W/nivwEElL2GzMi4kPzlDUAFPfRgioSUp2qGqc
uqEKVmm/w0619tYuO+T+iM45udAf9/Df0bCFT0EPAPHIbQGYXfwu27k3igred2Rc
gAEj1Z21MNPirte4mJ1GDQr2pM6ZabyDnucI2dEbK2trojeTmrhSSp3rU/Rcyszt
z6yB6dVTfTTY9JVlnkPHDt4wHGz4h5xFL+0hhhSwpKmdyHL9+Kkw6o3aXlAsC5+J
83fNDHSrxMXHs13PGuM5Bg9nS44zPnzflusyu7opgpxCSw3yKyAJvtcYvDfYw2AM
HMXEv7ThJ39bcQ6zB+rO3rCW7cqTkx6VZzQ6kdQr+EXFRgeL3NvzXYsFeDOP0Iry
0Xwq+OSlZctfcNxmX3oQMdpUrrTDjvGuzO3g2I9ZI2tiPSC6X8JJC8rwUbJB99Uc
qnKDEVfdwuF9jVpxTwJswarsQnaX2Ar5/9I4LvASiQebF5LZAquuK07m/KPU+kb2
p8N0oyJZwa+A4Zg3TG8vDEFYJmjW/LXkav0KVOOIV9Oze/VoktnXaxtzWbf3g1UT
CxyRyQCsxV9vBYv0kI3DlcWvJNz2chfp0c5HYPgsTsRsEJtrUCI/OkfxuRcPs+Wi
hH8sgmYUZceho5GNs7Dm/2NT9L052QJkqfIwz8g4YQ0vvXLD4FoW9C3+bYionT7c
Vq+jbCTtIxkWuhBiuFG1XkjSVWvj8JojzBAdRDMZcpBP+cnA+vtZN1xO/Mv3gQTC
ucj0tNR9U56LskzK53hA1gAI22KXLpH6uD0x9RjHFbOWRhtMAw0c/W1JT/XiZXTZ
hotxmM0oBc/VDdN+dkl+GBWtVz43Kp9V6gY5VFENzckcmsBGa6iLdLJ28U1aT/bi
X/75+kfyi4jAN1jQUhk8WUAp7OhaRvKVe+Okx40IcDXWAsPVVVhJfzOGGdRSTu2L
4t2lMWK5JHNdEMcl0sWXqxrK8p/YvYZ6eRP+/LAF8eUWAcdwh7kwhvfJZz56XE5W
i7i6YS+5b/IZ4tH+Rw7JIhvMLdTrYB+PFU1AuOlMV85vBZqxAQkxWKqTTBaIi30F
kH5jBWK1WSORFltrbNJkIAUllvIlsioWNcOM60L9mSV2/7jAZgQaG/PuDwmA8jYS
oXRg6QFPgyUKOMttQvtPzbA7xgSXzF1uQJTk11bsZgyWc9jVEm2MZ0cDKPDICd3y
AMumMyAjQjPFAaT1PnTVxcAF3b1nSg5c5XL9Bdh8ZTdItnff+TSdiaS6bpHU7mPk
7XQhDieajtuSVLV8CXuvmgypN+7TQ6qyix6Nqwqs4VutqZyGIWsAqO1rOz6zEIQw
zCuLMQoA0G6Lk8aB0et6ii1Y1J6OvenPkUNK/Sr9pag+bzJmnWGsHgY/5yzwRn5g
w8puFgVGfeslZAek3/PrWaIEZV+uZt54ejNW+bFvDvUzun/KrJw/KWB1iQPWO74k
LacTExyZD6F1k9kFz8qT6PFXxCjdD9lKPy2+0TZTtwkmIZFpFK3vk4NOoTT+DfcH
vjg15hr1u4/QcO51/NNRImlqucNYqkjoUSrOeibrynj4Lvouu6F3zrlz0FSzOiFT
OEWPmkLzxitFexrIG+xRq98LZ1OJ1qldPpyxR2bFFXqHZ4rXRievrBajEcn61T1T
/OFsVhjRVl3flONdil39j+P8s+oT5vYSOj9e2R/1zFggInen0vymFm04yhGlzTVf
gdwruutC8UDKZjPyVpDGDkwwP7VGfUGzmKbrytVCI176YWUxU1JxyPjGaLMQ/aVT
/nVIY5BImL79g4tAc+nrGIJUvZzmaigbJCN3IkiTb+OSSRvHRoC0/iCisVlbORRw
vEqY+7tfBpMIQQoqQkRXSG6nBE3sJanliVRwWXyq+OgHIfeGd12JrbNaIcB1q+Fl
X2JndSbmrCr0ZAf6ogsGRv6QOp2XdGiZo11sy+80Krk76mKrOc8vPMb9EK6fuhk0
6mKnUUiPABARuMVh+RMs2ZDI/WhzHcDvVshZsdaOOHnfNCwz0aO7vDoizElvGPfL
7nfoLtlZGXggfttCPLX9UFjptIgXUf5bQv2JBJmYSRE1xECjfc5o1NR0wlAtKnu7
sTyAx4vYjMgiopifrdidn2zD6ePYPqjyCPnlLnccarp5jXOAuIogTM2EzoTHDyA0
OOPUPWENWBmyiOgo4iXGCLUnt0+ao0uoNjBuSq/jLTRYcqVvtM8GFcM/3tQB9Kc0
JFPHfiHoTrXICwbkuaN6B+VKZ0AXfzJ3wKYsW79P6wSV2D5O5GtVnd8sP3yW6fnC
t9X1W/ONc2Rxovic7YInG+ZK/wXnMogUP46JeeTMPICVWG9/LOdWuCS+kKMoF4a1
1nQH6F/2vsdXgYSsD9eU+yFBNpyoQc4qeE28lYlgsF68X1jO+9CGaXO8jwNUk3I/
sWivKVOHmWoRI3fwINS3nXSQsqYx4xhGjdJQ5xobliN4XzJBm/IgWk2NlBgjpUNO
mgl58dN2DWq/FFdtr8Cc7pglHM8bIThAvUh4I5e35gurwDlMAKp6wn+b49ungJb4
FeFESbfAwVXo66ZuWZb7O7seKKv04CNiJTGHF2GdBqH1YloSAAIxV6RCBcNdUhNV
xHr2YY7zpyjTa7k5j6cJw8sdVHaf7HGqwRZ6UBtHwcqkocbN2l0e2Z5cCiE7csw/
sRLgFIYdlrDl9fi5zIRtSr62IxsVEphYwyUhZefT1U54dBHT9pVoczJnaoZS0gJ0
ODaOASx4nfmvEBHCrdfcLEjoWea6DqxumBS9azmYPiwW4t0SeCTU3Zal0k/DCXMC
UcutObJ1ejE6nYTOzD8A5tb/ux8gxzRW9LJHVwHmfT68SFkvOIRYD4lXpq3yRf1r
7IgW46V4+pZWW9/zYTkpCujy+r0o67uhZK24KnfNq3oM5+8ZABELuiIL1Op4Wv75
6SjJxcb+qdjYQ19mQb2z3CrRYiRJYTihJ4R99GPMJnd6eQ3FTd8V6w6PoEtibgdS
NxDBbjx93R0J+ZRZtf9W1XhgnK8Tksbc+GRYzEnHqw7bFlRrNK4I6TXA2u/23N3/
2RqHgGeQaow0itq/7f4ZnZczmxugGZQXukpPIXXeJX7ZEHOWV+/9NEfyy1kN83yr
volXrLQ1ZyUpKvY5mqvr1xE4SJriv/zpPSPWKzquBNbCQi48ujMVu158QOvbRJRE
Zio3yKAgHWbZKeiQbOkRDgt02FY/TBU03f/qhKvoXwlu16cB6aZfLMPOMmchZFQu
eugvUOOHG7E5teV6j2JnLFaHF3RkIAJPLkV4R599Fa3uHzuG9C613qT169zvg4Xi
oWBLlFyj31iDb6oiN6NrrygVfjTN47RvxegKzJPumR9OGS9mM7YEnHKFt46fyUQw
dPNp6kO0SpGwXaI1k9WuUk1skHsvI/T7H5Vc4vL1sjd61HUQScUTfIc+T22ym6jV
AhljyneR1FNYmLigxMkn+9p8PS0NKPUkzP1QyZBk6abPb8heBA4iCj7BvD7sK4gu
RGM0d4UVBCJFG7sE4pjlqrXtknxW5h3RdqqmzC3FL4Rfbq3PHZIMUomDxJQ62mEi
N4DEzd3E3CBP1akV/uhoqb9N0ESoukswHTxjuMLzvMrOb5VeaeKuSRdu7ZtB77F+
mbvYtiQ8AGAO8hCGziLEP9Q40+/AtKODwpsIDTaLnDLuQuLU5ASviptxsnCBdvKN
mBtH2DZXlc5iz+CrXRPrSqaJrD2lG3N3U5enPUruNzlfydjkNyl7TKOwFm6Ojrub
dPL7xl4ts8AcM8Syoit9W0UTfhfW9wILfGjwKT+U/qhfYP7FeSw5gTllpY0Zyd4S
0wI2pdjAlg3VDBVSYjh60cZYNRUJSEpo5/J7xytwCqpPojpvZZVmAQi7sJL0xAQ3
WMTIg24iG7isDNu4P8adgc9Oyiw1+hD9ig1Ss9Nonma0i+8HYSShKrMYG36pC9s/
GXfJaVXyBnUeIw+6eQ/VUjE/+JDu/Dk0st3pNhskPndyZWO4vxMfzv5M0wdrQcQg
IP7lPyXn5d9G890Nn07PeIdePudk38VmWElupbwBKFnDOz1PM2wZfhaeK7b2ZjQa
08ePvCXHDmuoDmuVmS6grYOr0l6iRyEeVgofscNotle6mEX0NX5Jsc331pStw7do
HiNBRLY9B1L3lhuguYC67k7eyIfiXijHgE4Zu52Sr/6ZP0ho4CeaLLoHODLwZRn6
dq3JuMohqK14enjzH6m8VYfwHBGHbBugCAVfdFixIpHsZbw3kqcvp5OLZsJKXBR7
1YkfodAuk5RBCivQbguXKktnR5YnK1n/2VoRghneVNQnRsoOYC3oat1chp0tQoT5
GJx5seqfSdKl4fF1HUkcOWXZfKZyBVil7kLD9iU50hCTGKpJ0HAll1SLXa9zkMFd
2bvyiJQfpXac5CmbloFOtSnxLSbxGfHbc6/L145yITmnbxjvcduUOygampAn7e/k
5QZjVk+DqEkc76i6IvhNdFDshc7wXxB4mjxC0M4dKfELgqMO5red+EMO3cR459cE
CcIG+VSnjXwbRdGHQJVZG4e8wUbrObr/TnU0Y9n/WQ4EMHlIdBGOJwL56CoTJNEM
u4dmwIE2RAE5Et7D1h3yjnqMJ6GWfWv/7RKtjJZFbxwdUNXdgwD+67m5NTSY7/vY
5BmZgidig0UhsJbMVj3Nlybdf2iGcfZI/2XgK8vJ2WYKdsziqYsyEe/X/f8lyPHs
yhNvS54FrEKVnBk4+Tao9Uv0Sjs8Uvt0PZYDu5Za2QiIQh2uzM6eb8iUXRbyRPUU
YrzW6ohn+U8IDCRuJU5OLUvkzMdI5igce6HtLVPzg2bXHlHcUnnhVBYEMSQSFj1r
a+dYkG/SvdyegcFOZutz1o50+y8brQFfaMP7DByUH+Pg7Ea3B2XS64ICm6y7yiDh
nPTrXU38Uz+8E6LjfLwUQSPd2HjUuVXQjNjk5pprrh/+RpEvc+kxDPSjEVu9FQ+i
peTIegwS3zrLS34IhzovtjvhgmqtQnnVY9kWgpkCMAmOjtJOW75C9fpg1eNKi83I
AVIge+cEwfkaEadVRUMZEQzF5cTbSSS/DP0ZitAKHF6MdlBLkmDxNEKZNLQJ4LLn
pIfqSEdje6ZxbYHSANYgDMPpaPRLkqXMUmXyR8uxfRiuc0RxZpWIO1LTP7d30b1x
2x0N98r7rwk5C7wWRuBUqpPcml94LeSqOUfe1CRHO/3gU5MekKS2vvfLTIECJ797
v4irQvFv4UMLV6jXbg1bj53OvDVVhj2ACnEAfMk/Zj4AMZ6GKkYHWI61s5YOUTxb
9ct4XLyfsS/k+yE6tgcn+dsNMEcRUMphuv7g7jYn+HjX8lS4930fkI0wl2ZHm4D+
r6IXdxWrTGpoz+p+gQ4NUKha+YT/IwaJ2wVM4Wn9w9KuHER+s+n5bn93CYdHE/QN
qBmoB6LQFPYxszlqYkx0wvM3xIhsEH27KBjszYzYS7+99ClASWC3CrGcdkxtpvJy
w79l/83XWEVxf73FXeZyzirvzczf/FzukffCem86Iq948qMnanIGv0kgJXPli1eq
xDrxMlqaO3nxWc1QDJhqxxSWK4meztrT2hX2eYCuKX2WBRD6GYhrayZG3VkP5hPi
MJqKaZCmaiSkkDeYBc05s/AlBWZ7Ldu7zYByR+tbIoaeWTdbXA1weBrKB6ZTkuVF
zb9gsKQD3xXGXehdalt15zsRZnh6OdTFMJRhQAq0/GpB6v183Nuy2sBEQHvfgsfo
mlJf+EIJkN1jnskxy4+JsrVwIJmwu6WaCc6h1u3ypY6Uj7BvYVuPn7NWsWk9KaEy
r+iYKdlThBbtVgMNi5pyVZ8NDI5a70/wxHRvNjYdPdOUuGT3g7QDZsFYmsD8qlyY
5MwfjTQBbLmJ4HubM5vN10HwYBnZcBycghmkHkknf82jG3a7jP3aZ8Mfb28GqFIn
JHXNyr/wPuD/1BWBGTTjIvOWsrEYBDzCiy3tzIdl4a/Tn3nAaWxRv+DlWCaBXnyr
x3C+/IyeWubcfK8lLgvnGHiUqmSSBEcC5P0rtltzOQTEEwhIHW369GM/SKlV49Qr
BbItOzSBeO4mMxVNPSqJeBIuKYD95t8i4ArWUQON5/j6FheA0NZP5PdysMk6iiDI
5LLesmpx2fgNk69+KltqgThCncKUAxKihqYj73hKldt8fE1ISiBMVDFzZ09N86R5
GP1Cukijas5bCJ9zx7gJnf+razOBopBiV6R7W63hLhnkUtDwi9xiq0UM5eAPKRpB
zZAPuzD6sFwVSVLL6IYbmI2WJIHSwgQTyyCI2z52KRdJziJ4lnHWE1cYnCJ6955M
tgQHcCry3vWP4dasGnVkjvKPnnP8K7zT+rWnV21xVhqV36fLJc246R3vYr9BoGkn
a68QZz6XcQHWd0bCeTd2PbETDUI6Md8TRcN1yLXd0U+lPapROIYkuxJWTxnGQc8J
QDxODTUxT0LfYBr5zw0e85Cb/k117p0zVdwpJTRqMjfBPEc2nK4swa/ulKRfgXSi
3Da9aU/26bz8OIrSJlr+U+eRiM+1EFdggpmPLFem177L3B/6Dn91j6ugaaw8p4Nl
09fDInYTgZxBVVphXMstMJEy5y0VuJs4O9tWoDbFeX9C82bPlfmdB2TOwcpet1VI
MQ+eiz2gO1gPZrtRZLGLHphM+zGLpYKuUCY6wsxgQPVo7ET9JoL8SXhVbLK7eEC1
uZaxKGZE9u8cA1JR7vdZnCADHjwSNZgJJi8HVGfV20srVlY1k/IpMbMzm4rfjoLb
FW0yP9HAO/PXxh2L0LzX2Z4zu1rkb++i8Rtkc0oCR+JKZWRD050EvO8v1i28VAUs
0/g1volFLMRE1B9u/JclkYbOqAlH72b/VNz/GYJA0Bib87sVT6FduF1uVfVBL3w+
e8MHB0vkoZ109Ajr3ywGyMMhJSa096NC1epIyzI4yCspCo48kb0WXLNQ2ys7K4cb
geobviIDNioMAnn2RyokWQykawWl5FQPorQCenPCkjQckglDy68kTLQL1JqbYEzI
4kWuQ4DHkMTpOOQZbFlRre3gUBoUQtQqsCX9++F8b7ruN8gnWjZhKcAggXiMJR2e
Ygy+OBQKPDNLC+SZeMfNCrw30h3r42+iGLWgsKu5/+ExJWRIfkJggApH61KdVB2p
bEMCxIyvJwh1f1bJbwGkd/p9vhXM/cRieBv8wxDAQyblye4MyUBoiWJa9sbWeoqi
L1hTMaQ0pFAAwt1oyK5+rvnv638jpl8FBVzfuYwI1pIpyxaOWVBTVoZafnjy+9AF
iju2qXRpJqT6sRDG6Re9mmtLognl3DuZWASdewoS6o6SrmG4QaedBGQhq4lnI4MC
8Paf5ku38paF5OQ4c3+jpDtw7tQZZorFVmxvsN42IvUNGs0W86gmU1IbRbsFJuvc
nQNKhMuoXpoSRGxCVV/jwF7f76pgMrDcwb+33vsu+SZuQEcxqNthyWc2ASArJORh
sRKVjIWy5Q7gncPqGTByZzPTgBAS9eZ67RwQ9NNi3Z4T89E+Q1ONyHFltnP88pyi
C9RyjKSWL/7r7VMz9SUf6qUmQ6cCw8dAZafUjplz7sSIqEJStCSDlp3bV/dXE+py
mEUaNc16OKI3TDm3aDdzK3jnwRpjsISijqXzW3p7ArFzSe6U6ozkwm09eybR+BpI
i1P57tX0Ok5iq/JxBCoJ3V9sSig3VbV0BjNB1KpGM3Q028LYJjeJiHvQbu3YMQAZ
dPyLj0okcRWE56WnHLK5+AmjwdeMspssq+7YTia9htCCaq13kiUCieP7GRA/cBMD
KSZowAS6f2kRUufrNJImj01g3ex0aG5jenyb9qMAC2MBEyFUZveGzFVbtXTQ4vIx
6IO4JJ84IoXE8fbolYl8QEyV76RzdVOuN22Ix3WXkWkjq4miiuq09+ZjM8Arrjxw
pORn8ssssH4K6j5NP3103KvfVF2glnc4pkiHPFzu9pDBzkt78iZwOux3qBT2Yynu
UZuIMFOtkQk6G7oWjGO5xli8ariqTw9JqzpgPsxioAht9qKmpVRqAFZrI8WbaC9l
WefsRKeNwzaeIy/VNjdt1TJBH4XgtH+ezF587pTEHTM4P3Bs6oqolc2qWJfqu/Vp
q4brE50bOU2E4hjeNufTrb3TmRYHowk/vM4ebpWD0v6dRf6o/bK3O9t7GB03NQjs
kc01xnS9B2y7GKwADVzp7DO9KeiNcpZoTHB4013s3jl6mGmtlUqm1htQP0tTC2Te
Ac7pT+aGbHwv9eBpdLvIQ2cFXu2mEsJMEdBHGpHpCPIIsIAHFkwJOeg4UqM0ampO
ZdSXkvzBBx4OdoQhjCQkh5JLTuZdU81RSZIsAZlbnEN7tcx1aI5wmEGOpUq+BmR9
N/gGOUzRh+UF8eay3BJBJD0d2nbgWrjyhwNJvx5rJFGY0Cy2c/6tAUD2foQmEe/i
WOt+b+dQ6vhiXPqytoX8k0+/UJdpnawyRfCCf2avv/iILYFAGvgIwCgxXHidjkUP
HMZQenFu40/VKXl3Re+v2v/P8hZZxRAUZrKGWOqcMGvAHsURsXFAhMUElReOH+L9
tN0lsqZaEvgkqyS1DRQxNj9NzS2QC2hjM/QL2gGsG2Gfm95QaxFzEH7gjgvr52Im
6FeJR5Pn9Swm5W/ZbyM/DKGmpVqYhIwu91YFZ4MEYhSYgyhbPoO5JIv6CKmyrQdq
Vf2jTIWq6lsSPKW5S8fV4wEHa/h/5Ldcv+gKmcaUGCHrlEXTlSOwK4v9XRoNycDX
zXFXwbpsvCmPi6s8epwpeT+Qh5qnyYJtHilJiX5Mhb0EcnXiA/vSFBtbnd3sHS6l
7uRNPgwbZciftJ/NCHllrspUkW8zautcG+iJt0Pex/gWsOoO99/pYLb37B/7r+JL
v3Lw5hXRVDcD30+ei+JPTwLrouoWHxI5kvtpvfgypODqc75DHgXJkvnEcgFzE9/q
yNRU1zPiacn1XeyjT2WF0Zd3pCyw41FsC9TOrayaTcolNmSrc7e5rObUo0jrCV+q
ttq6uVsgueABZqzs2TptKLxU+giWlWlacz/rwhdO9e9psL4v5bYZzkjj/nD20/gI
ZHrzzY+k3KN6Dn4Nzc7ydAQQk42RKa9s26G8Iq2DvaxKqCk7oK85Yfw/eLQnskVq
8L4Q1R1boaijMQzVMK0P9/1sp0Tca8xSfOc0vhz1uK2VPzLCGQcT1SBUTHmKyKlf
HUilsdjH0jkWOXcfRWbCdQExb0NQioVHwB6IbHUwXjOGnxmAygAZ7pUvxobodUbI
6Au4XS9d9K0LOn7pvm4gaYGK6yH4fCQlz0S07Vw52OcwlcWKnL066SM7VezC/Tmh
U+5xIxwqC9K0NPRyfGNGiAvrn+BtOEKs8GImbcnk9SMyloXPfoG6HiMqQo3uyFg2
sBUnb0MSP1w69ig/s+pyYpQCv1MQAsnQORp12J8wdTaa5d+iSZNEhttynQWQMKC8
ySxeqAZlivbZNnGVqqR0jPO6f23cK1/cCuM+Bq3WHuZeyUhKlprlDO9rsiEuSJbZ
xjMeH1jT54GOGcaDT6A3LMTCW0xMIC7eBLMrgJvCqIFNQOD5yHvyLz3GKA6FB6BJ
NacFP95S5VP+kPTrNguRodATJtD8278AIX9gCMJDaQrR8wQ1X65Nnku409PsiCam
wSE1+wMlU9SwHn7YO/I1FemF1yijbIM4HbC35ltznp4Y//JgtSroID3qCCgcJGbf
uJsya7SJSRoFkxKrESGB65W81GFWGU+Jo93l8/wXBS8x/yg++owNlh10X8EpgGvn
QCw5C5OwXbdB5reURMfG3K6331mdo32Cy8eecxCyIf/XYxqFuRVrVOtBpb1WTlGQ
FNUjE4fpQMEIAUe27b/Gq4k6b+vLePFiU6WHsK4WFZ0kAIMP0mxmr3nEU/2z4Ojj
4pl0dLtcmqlB+8lTF/gsrddQF44GHCU5zk80CYsYHgnq9OJ69fpjkNCm1pxi22C5
3LvGIsbxg2sDuiTEOxTEy+JlbUv3Wzh8IaMMbTWSIaJ/2Pf3+QSHqasbqKbpb/Ne
saVD95OC8z2kIUe4nVBPCAB9fkHp9ZcZUrTwyXppfJ3Hi4Q5GPYgJ+z0D3Rgrf2t
Ggksgg18R05JskzPxThZyAmCDWNS0N8D+zPrjjZ0qP4Towi1aVNfX5YgiuzlIMq4
FtCkrK8YOG7NgdF52/wnqsvNMwki9KmC1p5VkPz7LaCBbbXXYUv91jQBDcPylhmm
y5eJj4X/BCHVeXGkgPot+CAjWYrEnr3jJxPT9jtbJbgeEXRyzoybkwE2BnDwACFO
+99F4bdDOKmnhE3+VD4D73lzOge3U/S0PnAzCP2UyrxLO6aYepl5XlpCKkcXoY0T
VqrNk+YPAlHRivHTM7MgWEPuzP1LZS2+dnVzuMdCYtPDiS5fn5lH/cNe/mDTnCuP
bXTzgUa2pPGns41rwOb/Kf7z+6lRvq/+36YBphrdcY3hIAEWtENqH0EEVOpr5QN7
OY8TWrs3g79uLHZl2PyV7KvI2PgnCZElA517by8GpKyFwQ5Apj9DndJIE0Ls5WMz
c5qyDKW5y3ZYN4pMnjbrMnMs0HxJugt8KKnqY6vc1nj0XOdCGPD5gJCDcFX6p1eg
4Ais/VbalY7Js+Z9SU6zr0eYx1cMOc0qjVYvFtAN6kRpN/BA45WQdV7E//tFbJ2e
3tzHfBGcL3/YJxDx764fYnPrxSA7rBNy48U+1XLJmQozz4CxNEpQuFAPcCwa5Z3j
Se9oySMsKvrzpzPRccE20zdKvtl7ThxU9sMMzU7IgWZY8wzKt1oOGZLGg9qpF/ff
87oX+F7+p3RUXNvyWuBkBEsfxNApsbMoA4AoAQbDQ5JB5fCK4s0D6BxvxyMQLZ+k
9S4AVJxbsKa5hpuj4wH7y/Kew+uVxhcMYwz7axCtp/TFD4H4oyLYI7ayEXxGKPPH
bv0PuaMq7X5L40NPiIycM4zMK5sxIn5uroxs08lgYibv5pU1cnfczNs5zsDKTLDm
c/HQW12ax/30pVTB64baX19XCw6oNHhxhpDDzeJyrTk9Zw3kXyNTh1W7zLc6mbz0
z4+uV8XCkjfKO1Jn+AbNuLh2ahax0wxdYLlgJgYUPypvTof3pVe4y3FI6+uqvyZL
CsbBfZp0cZR5eoQf6F3PpD5u3uNQA+eSLtxZAVXpKWmb9KWGnwPZVMZFZBLBusCi
ovZBHboXjRXAHbXButIrZUBmdei9Dw9wdOAQEatnd6pWsIsk2C6VxqtvOvr1e5hp
wHZttoQfGjsG3rvu/op0YG6lrwqoFJ2cis6fLHln+ov97zppcM5LrQyCrxfs8CB7
eOy+rEuBxW2TekVlN2SX3gKZMxhX69QLTC2+VwKVd4fSsv9k+sJYtajmieXNElRi
Cn1Zzz+/YGiG99dQzAtJHHRAd1LJMux9H7rQBgpFfU7bKLgWHAxcrHM+K3xoncJP
dH4fv/Kb3QZ6wb7nPc5CFiHMDieeC8CV08cVa7sA2MR5Yq4Dvgk94e+iY/hC7EPa
RIUE4kVFVuWw1wF9hU9Br6qzYAaYttVBEJW/IihNYI2aH+k0Q1pZcFtFsOeOSzfN
7Cj7F6bYjNTsLaEqoWLbevcLFjk1r6gyBnuqHzJfybH+yZ6sDDvtoSq/X80IBKue
dSS35Wlltwa3gwYxcwi4HzFG4SS9Xuf9kqTWPdn5kRFUZm3C9gZGjRvhZFop2QfK
mVviZjt3S19EiqAkgnFPYRonHarCQkgU6kaaiUv38Yf1WZH2QUMt3B4fH4lUt0eo
ydihO0K+MFsgtAfaZm0C90ZMdS6g6G9XXZrJmoRUx7f13G6SWS0rA9S/P0Gs2ez4
GXVGOYisxzI1U8WZxLK5oNKzDLtuVIC0P8cACgeuqLOA008ZYFCNuERmFqGcxwGq
h/1zbZywjtoTnvW6XGBVy0sq4bDFtH9p1BjIsuelNjIAiiYr0NMC3+5g1rDoiMGD
+MbLpu+kd7N9cyXsVbG5pjxBci1sq24jFClL+kH9rNCmPB6fUP5o502UId9/IPpe
fyO8E5x4LdeLzu5xdcvCnhVXTwv7e+CobniGeAnNZU7Y3TYNFc+AIPKzmD8PR8+f
+nk6mpl3uk+mjZgS4y1wiHrhCCZq4+7c4cqCWxBWVcWgohn4K+B/fnwgaECcql3i
oJZAglqC8G8OuGJVpuvICkOQF2/unj8dhMO3rgNZeKQP6mwU42BORuZFDhJSlgaq
dhDYElkEanwIFkNecfgEPNoE6Nugl7ZCuvwsSDCiNgS32OjZ+Y+M6ngWolAKUR63
Je7GGTxJU0JO5PUnYaJiw5Cf1/WHQLofafpGtYuv2oW8sjnz5Le5zuff+hHTtIa9
ofls1XL28oJWtNnYvBhlUj6h6R0B9mahF5jxcb3ofG4rvmZl1iVJHL43MkAIhOA6
dMzObjpWB0DCxd8ehFCLtIq4ayqIlfIQAYufiX0Nm3SwlLfVomMSD9Byyf9EjhjJ
7Oe0DJJAOVCjOPWHjC2JntG3zUWdJzpyVTDlYDHRGg1GK8+rEso8IDCR0zWeCO6L
C+/oKy3ac3EZN+HoaCAXVTXcrhoWPqjk5Hez6SemJ4fvnKnf8mGFOokQ5NId0z6b
32rEYdQD/vv8Tou6UDnE9jOUg9iwzKKYLultGo1G3lA1q5YDg8QEhI6sGQb9Q2+0
sFOxNA42c5lSkdICQMbiTcliihvFDkT/ta1CVZ18NEQIAGP3FmP5qbABwetQyra7
h3lT1/iCZZuhPSwzSyeBIv90l0aERhnFM/pWUUJMqFOj5d6sRCIE30YGGaLc7uCh
dsgIPhpSss3I+sXGMjNw0nlRK/XfOSQ/slETPcf2kaOC6VCplWZwJTpwpmB8fxmV
Iocr2hN0Xk6ChrFtRp/1rrx155ik/P52DKo5tXhX/XvLSSmfHvIYgAjBKszx1kwo
JNKbVAWR5br7s+NV8kAWHQN8ZFje8vel+kBwIpbR0wx24xJUjNb2ToHkzmNqM++U
mfwEdgThuFMWSyNhYyVGbgOyYD/TM5TmpIfIJSdfdgT4xtRQFlbMuCOw6uiuisQI
M+6PAKiLZdkttjXCSq+axWV2d3pCLeuHUnvpJbHbkGsW7xzFG3flCqJZWT3KFaoH
4IQF9detbTyoHSHmqVmXebYRC2oZGGfKSDGeprUUN7292KuxmtMeRT7usvHTdSza
aYSqkwZD2blLyYRUkk/Cq+bh/GINx3fiJmgYAIHBJMqGTYqL0A7TAkbt8b+WWDyw
PUvWgxWuBgwvD97k6jZ/MBccVlyKA8btn9ZFQ78rW1j7ybVdL2J0d5a2byPeD5U/
KzKn4f/cOtk+5JLRhaTzzHo+YHMEIrj8gxtbvCvJ6zP+CgTm+eGieXB8z44gTTKw
sI41zXi+9S+FwwfD7ahgFSpsqeIj6xzsplTuB+n2HngHC6btWmGpDr0wgv+mY1/e
ff3J5bYvXr8vlgOOYunvECtv0pqZFFfFUgXBy4PLlNUVgIpQCAYB6Yflh1cmezAx
Hfudtutq+r8wqrl0FYzujFQ6ziOTfkkWhYbAyHrrwQmPRX4JIXO+T9rEiVUTJST6
a7M5mu7OG798rGtpaKMoYFhEI4KalbLzbhABFJHfUPK9mectnO4FjarIORdttfqZ
65cXkBmTIzRlcO/Da7KHYr+UT4OEvr1S1Q61zjqOO+p2L+Zvjf/5Rs3W5nzYrLzA
li+WIpIBs07TwReiGLATeLu+CBg+5u8aWqCCczNDgiOBzq83C3G3nzc4n7cN064/
BWtrWk981ZSWMoi4VPJlSUK1chvfgTZWT4jtSGRfg2qdIayCIwlDv2OGuwCUlhr1
I1nnApspHSOrxMNOMgDY6JIK5LwEDzGeCSVDTKUf6/usVA8DHLOIChVydap7Sfcj
VFAOcTEF71LSVIHpD6TglGCeWayJLZs0HA2gLY3Nx3lz9kmp+hgMsJmTVDQEI0Wu
7VnotBy30HAIADE+aBpeyYw1L8R7blyCn/AdKJ/qNIQ6Ns0h+fTeKGrdXxQ/B14M
HwSWZhfRIUTtahRUrdaBitSW750xOEYj2eBEdyV2ufgZk3A9IHOPsAgVJfRIQpQz
MaVLmY8k6eWIZ5viNQ5fNBSBJSHXQKyUMm3xLWdixX8xczgHyMqFgUDH+Bs8KpZI
kKlADmH9WOvR3DxnVWtYutnZCk760XU7Maan9d2T83raLfkFry6eOce6sefF91RB
ttnNGLB/OjNgYysFY5OmPtqnALoVVR3V/FeCxYqahKrC0Hi9kkI6HxYSQoxXV5DP
IOlHibxycSeoqJsZzZWVF65bHerXdgjO2pXuFTnZ4qfxg3VOpgpW1c7u03fU7XF3
Ltz2r0XQDjcjKxTNxaic8v9gzgJr3mZi9soSoNojRHzmWyY41qB79LSC2yqcpXfE
e1uLrT4FlfnaE4KePonPWMnxPqSOgEnqSKdI0OcqxUkxsC1Q0gCUoW8R6hhLgCQW
QufxfbIeZ/VSX8Jz7d327Fj+Y5QeEWCo7T3UJVEqExpewSwd46Yw3cmBoDGXIvNP
uVye+EFg5JKaWpLqENT577bhG9YWbl5s9IwwLPMUXrVP45r3lTMnCsj3SrfjseZF
DpPZxo/6PTfr4ZYIJ5LdyutRLws5U0c0USZTlNwE3mVtZBK4dJJgxp88HwFS1En6
KYDG4fpTStIxwQme8HwCPXiZ9F4qXuVq3Y6ip4OOe77nTH5pBCSbGMKRJAzDpysn
Bvvt9kaHHPg5JATbt2zO7A+0c5n+BhZ0lbUahbhRNcNCiGEJ3pb4w466DnVrauKh
9ALxzX9idMiKmeIgongBFCH3YkF2CETCB3dzVoR5p7xHWde8/ObTSiWMwnygaXGZ
xElrGKpEyPpdaEBKVJIVu2cpVjDtAjTC/dDfeYdCfxYV15cvB+3S9LW7kp1yDJew
b19E2MKTKUyLMnLQQZqyW4o4ih7msG61k/tYo+wlU3wYqEYKYAY+uhLPqK8dSSFk
NmmLfXQ7inFqgnkV0CCOVlXJs62XADI9GQz9ARlQK3n0hcwaBY2nNt49YgDrmTot
WqXhNDPNCA+JanLJHnwvR+mb1s4I68ay3+Hd5ZqXc5c4vtPALeFcBoROcmlYCur6
7HyoIuY4yfXWnsrAjCzyHjzq1SNWU2cWTAwaqnVZux8aIpQP5zMViKQ9ySUdYC8V
P2YHctqNnuWgRNK9BI2LNiELnUCqUwrXCbUB/SLBAnn+HS0r/XP4h257hNE3LGtX
wwRFiIH0jeCwy5mydbFG+S7qvY4XDJDqhGxwkBYkuymn7HwFOJ7bsry7P4EjQIXN
w8GW8PAX8GR1lWjnRbkSG+lYIdXWDcdQnCDmKUMr8SM+CCgoDVGbzy59d3MWb23x
W6bp7wstltI7e/foTllRr5FgiaZqx8NzG92K/FS1QZL5UbGM6elHk581AnMcQjFd
tdsE4YHZXY/E8Mr2cddezsYYV1fL2TD6NMjODUOtN0IJfFBdlVvKph4qq+D/5ghK
dwhYSyhUO14ktEnr5QIvAoOFNRkYNFyZGSV8wmCqefLjcYb7prqTw33R+7FFgmGM
jozeFFPNAYPOSLa5yX6E5jx1p1GUzHrU+/po/GNmPjMraRpo21g1Be/YyCLxykOT
GLppYSuWA8ZctZv23SQm9MXxHdq+9+R88U6HedjD09K2iQbkt9bzhqW/daMAmp66
rxZod0Bwt6THB4BOqjzURVz/pTerGiqqJyyA88QiECG8kC/FujOWgwcZhmYzzS+W
alr7R4vtwT1IRYiBhHUIQvy+xx/FZjMbtsnuPgE1EMhhD1t8FHGtoOljEODQrEI3
1L36/PqjOpBs38/xbmTUt2DAz2MlnlFhR5HYfOfSp5ONzl2hS1Anc3keXHekjmZY
0crFDxprCwQKBKxdYPQeM2OFX7oqgLHjJfl9M76H5QfMuAviTvH694qTtb0QvT3b
h9MtfTVCH5jI8PifFDa5uoXpRsoQxY/2W54w33ytua+xRRyiFLekCcFZG7nAOq0L
WQlrEri+WBRZgYhZ0xzj39wK04TmK672ip2TIhvX/kRcIjmITn/x0PasyFwqFVqL
Ila48JjK69J5WXCn4a4DmHMHA68cScG3lbyGhlTPbIoVs7Dlt33leRtJ4GdY7Gam
C5IIEOjSsy+cZAGscaIpvDB6XxCTU8ui39W98WxVqkWQkSy/6Vx89AfP2WR3Q08y
sJGfi/tV7VO5TNoHYv01Ww4D6K7HFAXC0GIYgrJdiFz+ZKqV7AmlEzUvgp0JkLzB
qDrJ+yQ4hfPHjesOq5wIzIP4Xhka/jbzgrO/rx7cvxPpwok9eq5iQg17kfusT8/+
VuzzuDnqyNCN4+yrf055YhpD7kFTBxw0Y7C85HIk6pNCD+3gLAyCWOkKlDm36q6K
W7u8zi9+6IigorIC8NtejpyVuWr7d3pu/JtqVw1i6qXUZkse0Mr+lMMja+9lTZRk
QwlAHARgBzOudOC1V45FY01Ve+xem6LtZmWPQRB7fQhZSIH1th1JaTtgn8enISu9
fy9TBqXm3OWC7GUR59Y3FPEkfDu9+zuj28XqE/5NXAvGyxtdhBWc5E1dY9Q5l63h
4bYALfViNgG08ViwCm4H+0unc0bkyjAsd41YrUJhZ4tEnj7HjdfbZA21xkzai0kr
2S+gOiUCgkMeohKoiUEgTVswaIlU0yaAQ42cho3rBlKQg24hclQlB0HZW3VmNxwD
rbqnmrgWmBVDqUqTKY7kF0ZPQFwLhJLp2ytQY88DVnXYUbMui02m6tqkiW1Swfz9
L7s9UxwRHX+/bxVbEXCqXomMEm+8xnv1C5TYBG+EvnfaSaHIBXfCnuSaOCwJBbk/
5q9D2GL0XdLs1i/HZ4UW/OrqX0CV19nces/9GfEHni4PWjcL6JljBkFf4SAxZyEZ
/iD6PZLFgRbEYdvKjXD1fYHEObixZL2wI9yMgvWyxU3DcbEZbggNNI0YnjbIL+Bj
eG4s5XWWrN7grSfBiIR1XrmKHpRurNfMPTmozqAuCi2LuvQ/n7O3Fi+gTT/w2KnD
DltvAvo9ox4ZqQYBznA26P0tPxJFup+Jwkv/RGPF9YYhyETHtlwCJIPNmk0rt6CD
5vsK2R4Qn8TF1MU64pPakMmT3Pr4LbyuC3r5MdwSUhHe37HVSseVZLB0c6gaZ7Hz
lWfdpG2ZL8jfdqSf8O7DQP78I1t5HX0DqUlxYFuRZ0a0lIh9vTy+elu0LqvXSuLt
/Q/xMHPWHvQYJ8IphYKhXnJmopm+piZYq9vpZhkblFa/C3iCs2uB4COPzk0B/uwz
Y5C744nOqLvVB1aarrKf78m5PiEUOBm+DYiyuKtbVjg8Qtzl3RSLCcco6qtKiedz
ywfRsHc+SJrwPgjqUMddqxQ5Nbo/Zk69++8jhx7smXU6pt3VzyKNU1C00TabsI/n
36LQyxIWEkm5l2ubCmrDCwVNPeW+DBQPGdWsgLydozCbzi9n38JTxPnnlbjibcCg
Ayv4Zji1E683/XMv41k7VqhuI27D4XMqZG9HtmblMHXqnDz5a8io8hBuyH9jT55B
+8Sj8NO+/D1d1hm9GmFkquWmNEI9jcw4asp6QRER7t/8tInDULEutw+U0vpP2LpY
mW3hEJ52zQuKLjglOcrBqHoW7jDi8CL9TVDZN6olrFdghalMwlSevxSAD03Cx9+6
ee1FFRP9h2g7wQ6IqvsPBMAU2LIGPrUNsTiwD73FYJN/7t8/DKgABS0IXVF+b3uW
4YM2/CvfOdhIBFubSTlbyEWCrUlAafLqebxQKIxAu3wcOIrLTDMfP4BW42Bd8/uj
r7I/uxC3L5JIujmA7JCFGSGt+EvW0KFGvG9QUtKEFbEGGAeQX7gOI7GZsTxml0IU
it537UxBKcV0cUHL4qGfHEIEej03EZoWhgYYVpKJl4aTMRKCIAGWEDvein/vENlG
7V3YQVDTSU0Up2Bpkf4MWi+xpbIlGF9uidhWY91ltsrg8LNL/DW+O7xOMq/t6rXt
q/R6GE7rA1Prb1hXfCSRf+FDaNCPHaUskbMxZxQXMI1olsNyxOvEN1NcaugcUcIS
DcrZUw3nVR2fxYBi5Pq4V7tNHU7vSXvbbaz6ED6ojf1bs3BckJJEJUxB7lIcoRw4
1jExkEiBxP5szc0CCM/awp0Nxo26Uf8qrPq1X8kA0c/S4OsbU6DKyirbC7diPsex
kPzJwX9SiwhhbIS6kth4mMXPCqeJYxwIcOyEzFRfVV4N3MNW9WkwpXY6ep/wVvgx
M8PJQO7taJFALR8b2lbcc8bRwh4tMFTq+39hYXZZRbLVYCFc//mlHgkyPZNKbplw
P/Q3ym6WBjFHybtLYDLvEYr8pImiVJClmTxeqiD9i/LK4xd3LkrbI85Q4w1opnFU
ZBThETGMm1PnHmjm0IA0wlAoxJxRGUvl65T1GL6r9Nu1nEXjLCGpukGuOT3GfV18
olveyeS5v3eBH1mmkj9mEkZdijYgt0NawQ85nhX7/XBG+D+Md5JN5wxkFTB8B5rt
6pUdPNHT0pRPp4U9nxJuY5dy0aa6rQGDJMjsOeFK2sRsMJd6htNQY7B0ic9zys0P
aZxfU4vsewkSrzn/NkN90Szr4rzSZjFgx+PyKxuPrePl81FSTbWdTRcz3VCtJsBQ
mpGmoHorf4BY9QU1fKgy8RW/0OyzcXqWm0ltsOOvsEw9sx2urtHGO4/k71QNqUjV
p/wqGA707WF2H10Q0D3IPiZbPv4znmeCrbeUppKEzLFy0489YWNzgM37Y9X98ix0
cQjBFQ+i3rEua6hj3xtVfzBVYANKrOaJ6Z62EpxU+M0OnW6KaQgBgSdWf+JzVGta
d4mbtF0SYsoC0TydAaX5WGZCqVMHGKi25KeRQj3SYYplsjrLeiZsDq6AfoAd5Wi4
pYlfK0iIxnilA4Gs3BSLaAzK9ncJbEyHPZ/lZ9gp/mgmhUjC4zF0lqa/7MfOEWEC
34mmPEggyDMFwu3C1/0YkD5NYSP8/KrjfTg0HNn4pPDFCYHD7Ype21tvczEQOiU0
9voBMCi1E8bLtaepAswWx8sNGat1P8ETeiM9r81olfVHxrgyZTMN9OjXQDwk27v3
jhKt83xzexfFSeLUys6aqlaCLXvAd5sbJDpeutkLJw5TTpBF0xSrY5FpDLUr3srU
YQN2725sAex/wZgw6XfeVhEnCpA8QgTniX4+JD1ywCAXc1hpAuevT22cVPy1LwKg
X5gp8j2+ptjebUPrldCLULIejjgI9/7+JfrcVXdNep6cIdme2PWp9oaPeXs4uU3w
WtbymFxLbJMhcss9VOBvlS3JDI+rJqhfggcaqgQped+2ZlvqORhECGotk+7kPdE4
9oe8LTf0+9nZlPkoSV8eZT62aswW3c9ZuraAtrBoYasdfhcUMJIghVJXEeqAcBUN
PRIv7ZWB6UXQaQZ18lMV/0Crg2cKS7thqJHQ4E8pPb0slr6D4OUyiYrICIqHouCD
e4Ic1SIXvtz/IGg7PXhiYZ4cz9dcaS+zM07WSH9fjDLGd4U85o56QR9xO28a8QKU
W19H/r2IyyTke7xp36N4tJthmFRzeaj2ZWRR+JYyO6NHxlFKE3zVCu/5ZTI6MOjg
Gj7SndmknhL/oSzLMQ+b4QgFjGESXhVWkdtUdwSxEJPLU4xJggCfW5XvnVqbV0N5
ObGHhGrlHbH06Y3BJSfLPbpQjRLeCQtAvFgcrnd/RWilQFIkj6rj3ITPZwDI461T
d99MY1nkxRMW5b5uSjptvg1GTtwoFblinalhzd7RdmHDaE1LY9pJdP3+vQOTrvKZ
agvoWTh59PmzDkb5xUjcPpu3g3GncJaffchtU4c12vFggR+dfceP+HjfKHvnhii8
FO2QgvEH1ERaC5/xXQsrwdt9iTx0v7kU6Wvz3OlphSAUVNeSEYj9xOKuzoiznx+s
xfODJomb8gbquB1fUCx07d/ONR2P4Ltsx46Pnxh7xK1PGGtfv74d46F7TkoBbkOh
BWDa+mGi6nEm0lo8tYjRub21hKWzBdRjY+PUvjrn58Z1RtDAOU/aa5h2UuNdhd5x
04Cz2stgOTkcAzgo+YPvv8SvxOiUoQE3IUKdgOsG5U3bZM6pqu80KdarDY0mF6aW
YI+hu766IO5X6E83XgETQS1HrEXCeNF0Bzkib4gZqkRmoHSKtUHFHxJcpnz/9s3n
frzPe31wiwdqtgfzE2XTSczbQ+4aEA0CCiy6VVjn3jUt/IWdvXrMIRVFsOI/Xs8Y
9WVwR2WmmmBBzyEFcDJU3ziyKkXCNxzrIx4JUlFAW0umVUMhVUVIQ9ThSCcp0llN
g6xC57+hCYqHAYRpKy8P+UMK14b+R2RxI0k/gK0DBVfqfhwcpoN95r+J9oMfEat9
RNbzuN3eDDudplG3yuF7BlwXSGccXX2qrg1pE6hAW5zQEsIa+I8Z47sMOPb4F+t1
O+2idriJXteUIHRKbWQlhU7lklrjae6F3KZzt6ufu7p8Luwk+eeJsOqBtd/CKU1b
Kzr6+Dnb9avcs6swwXRL0iCKfIjCOhrGnK+bwkRH6J33o9Jaqhj1+3g22xg3ejYw
vC/aJoV2rB72jM8W+altE3/AOhak3pKHsZy4vyuv4+nYpKmZPtsAtvNQ3+XETrQc
Ihx0T/7Z2I2vAJ9bqNHuXlYeSCDhzlWgZQiEyJnzg9B3dak1prC0pAH+cid5A9w1
4g4ydPs14S/9RErPKiUsE7RMbF6E/HKrgi+lR9y8kZCzSdEyfzufmudklgTxGebz
LGZIRJwn0ev3wpDLHrom6PscVEXshHvtO7CG/0pa5AObF92qFYXO4NEEDwccm4oh
DggSLsmrWrHLNiKLIpKwqGYqmHXZkAq/wAFwR+Fq78Dk+HH0mGjEcUl98ogx8l3N
NJClOojb/U0/+OCCyJ5zoN35lxNNqMAjUVnrYDy8Qq7tZ2sykOCEliSTHMC5UJIh
jzchBqAT9fs5/+qFhBzIyRyICcgiq0zr9W/rjWIBklt0Dl5KvKp5cuvZT6sbwV7h
qECqt06HHLtjm91G0/XeM5fkXZdANbpX6ItaBvAyF8pcG5RzIZif4T8jDOEYQ+Eu
RYDMYz5C/9fsPJmPEYs/G0oJCxatbh6cMULLYZ6dx3jV1FJYIFh1DfAAKoUVoUUD
vK1ngtbwKp+EKtJ+c2kcErjGcL2gRGfawOJyWP0Dl3s12z9aMwevJo9UIwkZz9YW
3qY1aZn7oYLKiuycOYVd5vNRsuLeSMqcsW5cMUPTdcpJmxgaa/gt1VT1rwFs3ONb
7zKnzYFWKtK1mDYKdT3fSGi51JISESxd7UOL8+JGU+Zq+r1ADxm0a18aqrWooRhS
oHZpYa5+VZ5WqI0gRLBOY5u1ZS4d8ezTFFYYoYSaG6rf8uwBH2HNHz156RpV+wYw
qnQJLX4M6Q2CiI14spxIzF2bJFMN+jPHjOEtFDvoNAwPkuBoSlFtq1w0qMa8BQ+/
/WstcjgKqeCHFe1VwbFPASgKTSx3zq5JdRfu4V3p57rfwyq+j+8XjSH8VvO3fs+A
2h1ukZDLH98+fPEXg50+tI7RkbQ/iHXWF3HcU6hnIqml+bApmnIddte69OlWDjm4
IGqC8qU9UB9jrSl7TLFlybj3oNlKuC23ZUY79S/Cqd2B5REE8V4RtCJjR143V6KU
VreHH5H+Q/cZq8b7Fc9wfRwO9QbB5f0tTQM4xzSwtIYne8aYqFR6SZup6pQnMUn1
ilSY/CukLqaSVQ7r5w1hcO0Spy7emUDYhDSbvOIh7/WU+p0VCg8gxoTcjIi9zKoS
YLEzhZsVNyocJriPuGvfmFYCRmlWpvwYz1rbu8Cd54xJnIukeY7rvLiK33Fhm6rC
3n26YL29X87ytIymSzM8980ptybaAapI2zALzhkT1manatfuafrWHP9rAH6b+HxG
KqQSQd6wb2kJqseta0hYnwOwJAsVh5i0iO9EIVByJtaVv4qV4Eb+sIf2ErawvUVL
x0BCbJSaoVq8crfWhZpVtC74WgK+88H5AvJeefAl5cqxl+HFDOMhig/41BlD4QG0
g6j6rvocxl4W6RzbUNl7taAWBuVayKofvFwERFshRZhmpVFqJQO3PIQxjagjoMNT
T82198gQCaoDsqVu6a96Xe+8fEEvap9LzgvIQrKppA880ZgtzWLEWwICkUh4hBtS
yTKfvyuZAmP/8DeCal4WjS1s3xi3bGLXOdrpI/UBkGbvDz7w+YcwSvQ2TV6z9Sew
TdnkKLHgyuIioiT7TgoerShXhdOZc9VONzwykzEdAs/cZSesN5gzBtizREUV5r18
sJ5upAeDD4KbGGtugDhfXbQ6gE2/bH0gL7YxTdhnOZeFFVBDo6t/0+EZrpv9VnyM
5fe2u7OIqkCOYYNXWytB9uyu+9hfcNbEyTgSaCXJrUNerO6172N9BeNaLEPQCPIr
hkDyohOK5K65UDQd5yRY/ykQiRJKo76ZY/MthTBSQGdQgQY43KPeo35GX2OPMokU
FJHm9xMTdRsy0chxVIiZxDMr3qz/bOUATj4P+jYB1StdWh70lUIKpyu0Wv10Twh1
Qut7oUZKAEgg8yv8gKuiEjUSadNWmmEjg9v8pi5pWMRy3GwR14NGZhBPxxDtO5o4
7KwFaqniGHOTU5+asVuPpjlsX6PFRS5YhMBr9kjlbLvuFO0stfhLMXsP4+zNF8SS
Fjqqfw7+AtDyQ1wp3NutHhY/nmW3EHKkBOlQK77eh5HMOhkxcwVes6hbf7EOqH3r
/0WXdVAr5k++wKrjXBFzADDuo595mzrLL07XoSwpS9Wc8/jObgcf7enijZV+k2eo
+5hduTco24jM4kh/UaSjEizcBzz1VnbDPh7mKHLeWLFgW0f6u0rwmon5qi512URr
WWctHo6Lbewh39NzMuA7NDaBW2NHwvUbOhKddTVERE1Mcg5/CZQtiTzWmRfpk/EG
Qq63uhB7NZF4RDHaKHCBrZMgYi0dTnUyqXJtXDNzWE7m+43P3HgiFfpy/o4Sv0vN
40cXKUedR9C+MvRVvWkziZaTmYJnmJIYNPGDDyLxkNYZ4hL2j6G/nckl4yCHNANA
w5FxQ1tR/gl/tv/IAh9DnAlrevNu4Z7j9i/iezFjOIy00bYVLe+9ioAFOXC/wxwE
FscHOd3n3HK7O10D1vMfqOCBOgZ2JynFJREJOYvJB6KD3qsU6jp+naLJW4Wd3/mn
ZfcCtTAyQeAXQA33glcjse54BfQmLXOHngsTmjkxlBdnBBFYkpkBBaGPbW29NXc2
B9GUQcESpOBoiT4IVtRfPWbrnPQnANBHtFUpfbftewEEluooa3kB9DF8zuHxrZ0c
Zvz+e6OZNB/UgeHHHluM9BlbxYPAUJvcKwFbMe3Sh12yftjKwqT7Uqgm+FCMixsR
4OFLQQ5RHQYRd+3gc+B0K0jeZznN/+V8TcesKuDPB6SBJhs7hf/HI4c5LlX7gxub
gldkDuz/XqbJL6TH+Dh6SdrWTnzwwK5607p6gpis+5fuNymW4C5Q0A1fVjiVPl8J
qnvlpaxxzA+RbaYgl0af+FFlpDxpo+hZZNaXzFwwC2VWXe28e7TWLtUVq0qVgE+6
yQIx8RAnEjY5nmcrfHSNsJ84TORyO2WCealq7oQ16mpBqnuq88BkSnrIp7PS2kyk
VTonL9qG05kTK7WCynfYNIsKvn1jTGyIS0N8SEL3ZtwAwHPjDgh0eWCsWtkolHFg
m/nkrUscsbA88i626axJy/UU0/cFWaV78FFwwHmYLrd0f/7iGTQ60g2mccbawf2E
IPBlCSCBSqoCt6h3KQX98pDqdRP5zHxUD9EMIyrg2mPG9qwn/uAkK4xieV5LCchE
lQzTYzYRk9TF1Gsa2dUs1WXRZNiETW0ay5Frlr1VU/pad9x+zG8Tc9kZGuIVh+Dk
dbz02VCTdqWsantRIRKCZqdQGji/LafQmk4NJQMkAUuxA+FlA3KOir78X7KnxDfI
x7K6jhGEpbw7Tvg9MNGS29Bd7AR4nPZFyoHcjlDHjGqPBKo8rb1BwbW0xuOe4kqf
TZHz+fSB4l0C65IbGsPjffVfu9PxN+QjAXBC1H4zA8S8P5hTocoRu2gqiFYV0/9T
BnVaCktTR7ofiAj49MSdy84okyvqZ/sp7PXUBnrwQim3D987nkk2O1GCRtaB2zC1
EtW6JfUyxTQeZi7PHBw/oMv7hzTWjHT9mCDYc9+IW8PPi9QZ2pdv/vqY/vOjdTYW
c1e0lWjkGiMUl55B2RdKawpIAJTHc7wGU/MTmVDaz113bx46p6ecNhdkTI1YR+9M
mj0W+L2xRXrCkfK4hz7ULrOnOfLGAAlcvoKxcUq4cU/Too4pwZ1UElsWhw+Ey45h
2b0pICgtsI3/NH8XHPTSB4f1Xfs9wIepEiJEofQUQg2/iNGdKVM5viHn85D7rWIU
8bL2TV7cFA+NC1hJOXB9xGZfapwGdBeORmEczRO8LEHIrk2tFkb4rsYw+6qWYIYA
zavR3Xhjcu9f8n3s1CkyVRPPlb4L2m4xROU9ZJ9yE+bPVSLrD2qZ8L9+aCCMXz6t
nN9bjSF5gtoG28lVbQqi9HymtQxA4aRJp44c6bOzNcxTUPYR9y7h2j+LD3AMe85h
qaV6BMTgtkRCTLBjeJftQ8q+78TROef7XqpDTnAVoUeyt4GtfDl0vFrIb9h4jnlj
OZy7aj1tR8j8YkSxAcZ2a3TEjvgn0XMyOiR8Ar30faYy6qgg2v48Nnh/hQ7Ijnrb
5vwrZ4ApAA1Z3A4JcLWZTQyWtxLaHQAK6CcyZE+1AqqJxxsOdssyCfb9mtd17UEm
eEqHBrgLSWe461wL6XVglcHhrdHXuopNLMcW1wou8+mBjVCF5u5yZwfUz/u5LwZo
7eEBM1/cHDBkYYVLGzMtLshpbezQba06oeoqoGsN2VAtURaEj2YNKWMec1yD1ClW
UALiyA3qYyh+MbcQ+zW9VG/Fup5eBQoCnurngRaQpwquRupNLe7ij0vBBm0xl9C+
+f+Q/sCDw6z3S/+m2sBjcR6k5ji+Igx82uw+7G2bjMZ4D294WlTCmr6jKe04Atse
utxQkllQ7ct+/zV0qSrpvaouvEoD4UWVqlRV5PHb3Ide3BclyGJEJak4haQfXSE7
zSLskMk8HlT7gl8RTM25DyWDt8AjpgkMwYbPJ+tBk9ljp1OpKgWrXtniFab3oB7R
9s71aNzRdUrWfS8v/9PO1lpHZfBOk18Rpnr7OPQcDdqR1oUq+TfVV1Cce+KiSVGy
949MXRXm/8GLGkaoV06Adbn1LtPDZSYP78fFsfa4x/CIs3/EcAsKeVF+ruKZiSzU
oaGwuNf0Ai27OZXFQG2xTSaJCUqqbAf6C+S154PVwavp5lVR3yQghH4gsGPikgqQ
ROad9gE8ufJJpGHZ2FzuY+z1+TKJSYiCfnA5qe4NxfUa1+DfyGx5NdQb+hnecCIp
qx65RM/LSGkOKp9JdBIBEhXWyWJfFficC08TUqtTGBpex2FYt52uejkU26uLEzIh
5L1r8r3eV79R6zyIFnoKhghi33B3R1K8LnGt5ZCaEbg7Wfml9KnvwxItprS//rTh
SRhg0xIbS4nlEqKrK4v9wu/n5j2FK0AQzKyMWbMHg1JXL7Ukwme+0dr/k1xK6mex
1dDlh+mF/iw459LbZ/yf6KJ3SwKUx8BTbty99OAvuhKIbR2X0WbooSm82J/oQR0I
ee5asbB3BodMwoMsPUnP8e1iVGbrYn/ExVB7RM3Wcrvg1fWJaHEkmQ9SjeK+8o20
0/ltCDHpaODizQlXpaEQs06AQHZC6019SRNd4iw2kIf6i8jlo0VcgPJ2Ed+CTa63
Mls7T1fq8l+1eQbcuwqI9Y3vz3s6aB+Hd0etkEP+HkDekA6IE8VyEnPScOV93O36
mDGzb1WlTS0QMnWOLWFtdGNLujYJj+5uDgonnnRIFJ7D3FqtaYf1zwFxMeKe28U5
labZzwkgWP7swTsX/N7Euaiv1DH/sAXBB1Zr6falaJFh/T5UPsKfRdt1eBLTS2al
bvmUPeZCi2YEw3H/9UlSiTUDrxwSbvk+uGWLN+0wGBVeUUOduSnQwVboEjEPPWUj
dx9gXwNiC5K5S43aWdAN4VsUi+hHXz6NSS12QJpNw7CXyYjEbIiwUiZsKSlt9fkB
BkbWsZ3j2VSv6tseLMfxFA+ylEpypNCzDLHxXjqPu1jN5/DiEzUy5E9Dsz6YhsNq
KnwBgvMBLoE8iwtOHGeRQ6uao318TkMozgJ70Z5FMlz33VYKP4seA4MmQCTKoZ2t
hHLzFhdt08nG7lWgah87y7vp/efSXTWNeD/J+xGEdtVAcKrUrjxPeqj9pPtjYrst
OMwzUHqxlMZh34F2Bb++nC5NUE4Psv+asBE3d/B5Q2+E2rS2lWLtyS7DREFBQfgQ
Kjrl+on3PCmkbAs3ve6tsJsAyg3IVkmFKwn18rivpxWEu+nJp1VY/uK+1up+AuNm
iwTiBvRokxoRrE4VReN0AO49SFcRONad5L22oPb3SQYA4BD58gq8eFqYmIVHR17l
f6efb+tkFbp0eWqKpvbH/QXn2vSz3QuMISOYo9TC3HAnHN+JVjuPHnTz284XaRQB
+bBQaY8FLv2QUrZhT661ZSpQHmHCoNzJzAq5jrAJEdb6m9G6oyKcezmJfUYuTB31
ZbXO2H4xF64zWqSR8ot7gjPHKFcEdIHRFy5F0oZ7eR/D9LkhETuCySEL6IJwjRIG
4UH8cc62VqngbUOFFlUbLj4HkCJv0YxCJ1ESH0ROJ3FNG1wK+toytZ3pguIru0v3
JZUoI108omYXSkDSNBBtrqs5s4VJFekeKCSzaCbYoUZaOzuS4hJOyKrJZHQrmJkl
awxXAFrsEqUqn4jvU8skkkCxd8zoSyQaRz8wR7xkzLodjJ4sgIzWAjm+V7za/8X9
CT5479js9gcVevam92p16r4jS61tjA7iiV/30coFkmXCUKMu0QZT9cZq86RMOcXQ
sIeJW1wnNuMkoX5XscGanwUHdFom6oxyfJOmfoBY3LxybMMGnkLRaDe24VwD68sI
7AHmiFINbNpSxjgetvv5IgMWw3MVWDtpvudf5ypmcBTQQlGgPKrm3bLB9gGN52oC
zoYL2w9qHmh6k3IFMofTomlCzUSICneCqHm5IR0mAXYeQ8o+k/UMd4OEib8I1lI0
agerAAE4oL0GQgT2OR70B/V6NWm3kCzp2MBpSo0xmPWBRBNiuejQO+vZThXRpCRq
8xdJfHyx1c0bmAmL+C0Nhk1ExHZqsXO1SAlVlsiLdULr2k6zxpKOTaDveHDvWDC8
PWJK9b6NTgiR9ZFi8JhFAgONVtDYxC6KThs6Ck0s+a1kOkhPRlJXsu9CVssWUnf+
iXA0F6c0T2EDPkJnjE1oPoXcZke/wi35OGBfEasxdy+py9ZmTEgUgYT5iC7A/qSB
/aGd+pFDVEtBFYVY0j7J43qDQEdlUs3SBr6hSuAd7dQ0+aaOY/qhfx1Fq7z58wGx
bDCsNah9KXsC8hNIR0yEK+kSLAxNcE7JdJe7UPMFo9qkfIUv0TsJ0pszpgyKUv6f
t8/oG9MP6GR51yjl07FsE2a7xKo2YbyQBYlQm1yjQg7BP2dUPiwVe0ANbLK19O2P
3H3A1aFmKuvJes7MR1RCdRhJvRMEqtjI1aUkgTDqPmBRx10yQB0YjM252tnCpSNq
5i3PTDB19NILhEV82x6wdPaUFgLpV1zUbuJ6Ue6bcPZ+OE+D6p8RF32dXYzvpq6A
NPq0H5Ph4s+Xd2MCfWjwz1/ZWZyisW4I5KbLeZod6Wc3/lzNcUQ7DmN10qbaQmT5
gg/Cpn+21bfXTTasMUEUVmA1MZHVA2+6D4GJCrp6O40SqWyX57gTSedyfhsNdrmz
w6qsKFIXUILeywnF9DqP1uXewCvm1PTfJFz8bFAskuT/myetB0V4RwjQBEyVHF8U
J/UhYUCgG/gfjynodciZvY2kBdIGg72r8ZYiowXfxVG/GsxE91G0FTUtTzQih7Rr
L4Taq4SBjCZDUVbam/mZGwXu943Ael0GjSKBQhXBtWsXYMPby+qS0sI+xAfFBYSo
juwTRHQhVvLcVF+slQhtKNn2BmqtKiI7eoMR9nZNsZvshZW2M0qViHXZCPyz2aLe
h0+LXQSNtYHaDa5I4gOzIrNu2gjxYTfhSzZGROMMVbt9gtsGgSuZj4a9OjtpZX7o
x34Q5A5MvQiz9YjpSRuLmZw021Vq4Q50MTn7TksfEZXyF654rmLyaWVDk6FryEG/
XVIAsRb0Q306/9rdj69MHzoeNqfBvzxVvynd9xSUrhI2Fr7joS+vLXlqj67lLp39
mwUH1MAPY9U/uJYcY8sfCkEsEpkRBlkx5pMW1fOnD7WhMNNId/SHPBibfM+5lYsE
DgRlzh0kuVlyrGbdMwMX8wy638UezVHgBZblgwQROKkVojynu6/YY4WzFdJo/mDh
wEjrcfr1ZQyoD9G/Dsu88/GN/OUvMslVCADiWKO0Gmo3D9kL+LdaW8rkhfC+t4PA
qvsW2cxXYkSilShHESW/W62JLLpVHobNmwDZoOOADC1LaupafJwb0JATQYxjaXy8
QSKK+Jdb6GcYqJXfqFe8jZZ5cLIGoEKL0QN3UVbzf65EwitBF00jFFEclTzyqD42
kWd+y+d67fTRykVbPdhXbJSfabAynfyxvdDzJFHsGStIQu2CDt5SBc/A3+kQN2Ny
vP4wITVk6bFZv2Mv0beoACQXK5LX0PgHJkPCth1TfHgL05VhzwyDGYqz9d9XdZpu
MdEJrQJwFlQN+PP+XNIkJ5v/hqMeDlId8Egv5ZWsQTdfmiBUnqMZh90lFScVmeEY
3ICZI+4Jj5enQ+bnNJQvqNr8OgH8H3bf7yw3pNza41xB51OyCecbA0pdUFExF5Sp
qDQEJksMMZL/2TxmBLXztUG0ubXaVxjUlpbxNNw7KQHZ9MbMRt/7kUETrP8Sd3j9
3nCSiul1ltBXPt/fvEWBkG/+mrbagBPctnuba597PYp2FGYuP9sIPqO8u8Lun+9Q
9c2ynCvLSXwLZukP0ECrz+pPbpJIY1IIirr2woQS9nkXEikzHVuZw0bM/O1ZfgSe
k4bX6axO5v8AS8jNw9zI/yFWsPwULgq6VA8Uh2THNJxZSZzChlMK2E9gsijvnfkv
EktDdRyaq8vUL8OQ3ZxEdC18MeVtaCgRXYg1b1a8Krs8REpD44pKg8jA4wm7J6K7
Oq/1SBCpwr7JUhXDyOFcy5OEh1XK+sTGl58cYyxG7TeBml///QKqMXRL9l49+UBI
+rJquF8CrrguBf2yON+Od/lmYz3jatabvYJeaE4r42T8PGfO5D0+AEgtAVW2m+q7
R1sxmtW4fG9LENfntrjFB/xYlX5dWQoLBCePGdzo1nnwkyDZeB6NqU+o9BQVF5Ti
0MR73IhvoLIFOzd0fKZl7t9ExZYfoy0GLHBgB0U5gegI7OBSHnRmhJNDkK0rZOPk
KKHAzHUodMQNZyV3tIw3yILGhHD/e8yBfZNkr6Ba0PZfuBGKHbyvlDMmZ5dETpWf
O0z+tzrLuXBUIoEtv3rRpe0KngWbTxNsB5tmkaasivSY0p9uxFyLeuqFc5rt8pa2
sFe2Sxq/sE5VdmQGnQ1pKK98b7m++S8+jUJ4Py/2j/uQppRkJUgbFJSdwemyzxnw
Tqj4rZX7acbgBgVI+6aLrHxEUdkK5WocJx6Tf4Go05yLfwJtB6HkarzWZ1FWemlu
b5kyFY93FHINvrF0wsbihFVwIbXhx/WDr6jlk9CygMJOXO5eKNJ6WoSMSLBFl63d
7LRJ4bmhJhi4IpudFje4AaMF71184amQnG6bx0NtkXbYxAQlci8G/S7hUd5Jg87E
NVc+oNc0P1nn7Pm9JGFsJI3Wr8SxK+BVirOn2EgaOYzF0C/r2qDDWU7r+MKaDLHV
uf3hqfIgwMI2QaKvPUXwJckomcfYOG7429uFR9ZRuQHyPxuxw+6BiSA3VSTwboqC
z/rp6xdCt5oGwkF//aE3pGPmmCku1DZ6Uy9nipkI/EolL1NLW6Aj3DhMGr3gIg5L
chNI6jeC8jk+6witKwvHRufPO/ktXIoum2IIaA4MJvmYjO/w6DW/OQ9/baBy8T+/
u0duRFjj1jGAqev/2dCiV9BFGV4kEKZjOvLWzKryQeiKL8NcK3WimEiVkTMpnwQV
RuXjKsu4sMQ9zb1Q01JIjGV6s7SOH/+h+cOa+1zyfO3lmQ77ezRZ3KPsuoZ1nrWe
eJDc1kLVD3vDsv0l4l9r1ODgduBlMxFDVb6KbxW/pfJ2icLeu8Whrj3bPzHssZW8
6R0LIYJobO4PCKFKo0xPkBmvGki8Aj/5dmKwqyGxXAFzC0QcA2GF/X1pbCWXufzy
gWgxRMa4U6I8DRkui2v7+LYFjywADPZfdKaNDqE9Vw3IiAqluIo0wxZ5TabbHbik
x6u5Xik5IGBG5dBIGHh1/aCX5c8vvrv6k7XYUv3BA9qo1jxtDJUDaH/mYecGjpVg
Df9O0uJBAS4wtO5U8j3e52j8USbIaI7jiVLmPA/HMswfgZENp+FAPWMXvqEXk/mP
cOPgwmxeh0l5/rnmdWVsWnYjGJa1Zn5pYVc8twOjYl5kiKFeswQJAzE3R1HWDA1y
G7Ehy4XMWAAxQ1VqzMNscRFft6ACD+FH9IRZcBTlwHAw428/e2qNzD1wfrkX5sWz
OhoQ+us0w5FszWG5YNOjfyJgKdM6ivtAYl/kH0qIyXQ8A9ubbXX20L0XqYB9iXT8
4y2r5Ez8zA9+Rle5CDkI3R9hAcv0FYdU/pNtp21utenAlMHyaMpxwN4kW1oKSqF6
wewYWNiw2HxefVV1f/1MrtSwxAkcsN6gog2JBWV9ZwNY/Ce4P0DMYXTrAykRcb8a
3janqvoUYNfMIKpelWrkQeupq+Ro6sbqAvYU0R9JGBCmysmG88IUbqCpCSIX3pRk
AbKoTNBR0lbfIpZXWF6/MwPolzN960GhNY+jz5LrqKbnPMUTjm1q00JjkguA/7Ef
wuflTcbluOR+pyoeTakdunKC+ycg6H0LZhJ5Y8dfugZ8akYCQcb9UtBgGMhTLQc1
GrTszzyv7HO5UaCGVJDaduc9fOm8Mj0PQ9xJ0hmQv/6IovkHVS5FyLZt+NInuRHh
UdY8MvgayLw0cAMaFR7h4j+nWvDym/977IbLOACFqaf2c6xykqKbPwWlfs/ezOnc
QygUfKK8UnwuiGm7WPRsL9igYqLKDntZiM877gC7TkTCizz4UtxsJUWnGZzxWsjw
4S3y6HM00B27HT8Q5jjBnzWIbR/y1UGrfMssUlaZXSOoZ1Hm8T+fnnbsN+PLPnxn
QA6QLYZjfNryOhPjP1Djl6QGWjwERRJB+ArKvdn5JpYLUC3ENJFcYQxTSBdE8Bom
yVtKBHLBIZaTnLI0NWREMRYLpHQi52xu9sYgF0qBzj3YGbXOB5+G1L3Dd+zFNB/V
NLk8oxbzoIzZ0cGilmYeL5cwFHi6BYOQQ8i8pILht8tKw3EsPCKHvi+Uosg+G3JJ
PHV3gH8hofaRI6thi5gwq5g+6nvOTiBfrDmU+/+7dEDsU4vakz6ucvKmkp4n4duS
Ib4hgxzrgQID6poD3TYdnObrOMlPo0Hw1o5ncVsSQiW3d0fI/dma7SQy6kx3m3gL
tibHJNRgD4Ow0fKahZUDESayLncFls2pFt9pf3pqQ3NPI7N7X6eLfHcbkDKiHM/0
oCmUuIZeIwRS2md6kiURwe0phE/MsfACD/xisNuXNmzWiCKasR8X+w4g/aSFTaFo
htAOLZZGB/YLq0R80rcvW516myF0FdRsk40NMqmUiLNaa95voQWDIf/QZjcCPD5t
c9vCFK529P16uRluY7uze5Ro0CFfMBQwDbi7ZjdR8nodVfTF00mXhttWuhLBrCsf
lLOR5dnSWZnhZ2bxFDffDl+Qjq97bXxxZ+NQxm+ZeVS+0qpAtcXvRGkdzQBHF3VM
sgz/PxS9L78fDm0zDJD6FP6OvOITHj9kInka/3nHhI0yUbc6pwFUGGZElSBb86Ub
leGsFvx3nyo2ZI4vK8hZH/8UeeCGriQsTSrCOa1h51sr+qEpmlWH5jy6ZgvI6k64
xcZsw6mvcJcI/51s+//AZ7f6s+fnYoErrNusobUMLonjwLZaEmLqgJo89a+ELbPt
+mrK2WjuLoJMbd8qKkcyKoOiLs7/jduLaYKrZ+GX5/+tC3hkGv2c+5Vm8bBajZN7
BRKe22hKbqZR1gGqzuhPM4gwW7OWdt3aJAiZcXCfdcANtCqaFHQ6zkuKWeevQwdv
//zNnIY7p0XjbTgMpvNjSIWZ8HDv51OULO2sg0n3eRKkiPL0unElKLpQszLEuQzl
J9yeDIZOc7jq1Kj+OX5h1huBgzuo7MSxp2bk6mX1ssfUSKLG8O7x4AzJFvwkXfD4
6hUaKUitgYWcMMN1fVLC3y651SMu39EEgfsT7AdZRzMxbKhh9NbJMUUOdpcFfWoH
ou2T+QuWyOv+CT6uqbjWLHYrMqmrWSL5sSulliPpFdqQmQT5n4VJePZcP/cikaUx
S264DtPyHa8kdm2Kl9aLzJVd+CsSMGYJgnggVlEoTda4+fBgEAIFc3pUo8JcD0ps
ClRt1u0B6dcscrvyyoFAg+QkgMU3Pg8NWBQ6KzqlgHr5wacUCjUsjadF+b5+Wb0V
9ZQe75Yc20iYMlwZRWeRCck4owpT551G+x/GVIjr466BmW/NI2ptvYwaP6pLNhKz
5jV8HsmVZANSOvMAgdxdRTMDonM3V7OkDsUmCa3pEEhlIerqR6ToMSSvBI6bfqHq
A6BdJrQeqxQZXBumS+kKIFMrLwn6zxWyUVHtcEGjRpwyDVk1Ah11JTzRpT4a6X2j
WADSLLGTyjs1K4RTqW+XCRYE1yJn9dQ39+Tw8flalz/BFxK5YFTe0ud34TIDPgkR
9xGOCk1YB7NcWtMG7SYdbXa6jGpwZ3oyZz09C7HjYLtgrsvx1OhdAr/6X5YpmUuC
ViNOLUuulLJ20sfVWxcX+Rh9VYkRWoOKZiClSOdVYnWhhoxCBKhHJDdXrlXenwtC
BJPeudRKkcmeeK4E/4nPRk7awdZW9zilYATK9TTLDHgoIAo8zOdYQrk0xf5v0ipf
9bS8YBpNpBB+6PHKZYG/Jj2aqmV5uRz43fbOyxaumMucW7BqRnigrw3Tphe7cLjT
Bg3YUluV3fh79iNOPsNT1CIOzzBnc1EyM5HfT0m8FdY4V/wWb1x4hL26M5n1X8RF
Ar9O7yTPryKojR03uuerX3ubYlYIPbioc4oxOVcehgc3YVWzXAD/Ako5Z0u/5Xcw
IFDpRJuUemXl6Tww0vYUAIx+r+jA3xoHlGLBg9yA9AZT+lGGevwvXJOOm4KFYavh
9uGpgUVYEFsmfZ6+dLN0e9itT1W4QIStNuwXnKF3K4u8jBh6rYCrUEYfGK4CoDhl
8D+u/oaj7Krgfjeyd54k/WHpvlrOKbnYRz87O2mRCzmBbUBoyBdapbWCFTBeAX2P
HDx0LETXEqTyer1ujwwnlQumgKKRCI9++Q4+bAW1BVtEhTNUSxp3b17rWjKokhVu
GwrOmbQY2fbp8HcQOpPO7x8E7Y+vcWg3LcCjc8EmHComNI3ro7YVFiyNRB6j05CV
ono9/8P+6Z1Y/xIMgAlm2aqkCN5NnAcbRamnyS6IugmIfzuzwRHh0GlANwo7UVh5
LBkVKJILbcBRaljsClXmbDdmER9QbBKPHgGfvs5IyJY/laHk8v2iEYMnhAzFVNyV
8dZKipt8g+SqeFYsw2EA53oWlkphXcBCQisPjjQHH4N6y9/S7SODrvPhGqfdORHU
HFDq6DK8mLGwhoxn/ohcpWFfpSJkjpCOF/uaGMdVSqtoX8ZeIIFTI08OJJ9ceWs3
HN8iJAf3GhcNn2o3i8x+l4mpWxyO0VkoEGxj2gIsOz/JQPVm06xMa7FEzwa7HW56
Z+MNRAf5QRkQxuOucz4UsMlJoBVwPamlM9NbvYb53t7xMSiXy18k/UNASituQEj0
zqPzY+vED0oQNXMJEEM37oiMZ2eKOzQCHBWn965rEFei30/oRk+3gkMZt174RXdv
zwRyHd2c8Lb6Lxy9Jz0eTApIK7wOO/m1E+3PNBrWUYP04//+Yr+eLea3pylp6RSg
XtFyqXIDLQkTVxVTfqSYq5miugM2sy60soA9U+lALHaCBlmnWKCeM0qDrofvz5oC
A551AboUz0satxqEra1X5QyPBxGnqIa0JAKAD3HGfxUMrRDNk4YJUr+uimX+3gD9
5L3tVWHQ3fi5pv3zXhBJeAKV7+T55WIht7JtGLliSJjeOscTrZaMvbIyNnj2JEjL
zrf6/2aoruiDtn1SSXYzzw6kxVlnDwVTteeKXRJsUOLB3EcNjfrwNygTpvK/7EOg
BC6exxFs7/xUQY31AzTPi6Thmda2YoeSm9GFyOI8BlFdzR6uZe8dQEWysG8xTeiI
mLQO9vkciup9oBUWVu3GdHZR7yrsdXbpLLNAhXbldPfU30KKqw087ZZ3izNTgQpG
nCCiiYgr8GmSeYs37mdLulMRyjTdptb9mV+AnJdj4Ln+62306TeBLNbBHVzcslIq
BcpCnt8xG/qdzhc/ny3By5s2v/pfUiPOhXD8qqfcIf+UMh84RzVuYXn/cWXxrJnQ
S3AMUu2JD5PbN0BluEtmAkhAmczamp1Q2u4bnIKWjjtDiPy7mEl/z11REq/E3LdI
PDIL5H2yMej3MCxHxOH+w+WBLzdcpI7Z/MgwwQlICTVntCKBj87QCMyrJYAualJq
7DfU6CkN+i6Bks9g1awTZvi/8L6QT944WwSwN/+JxVQyVOKHC2j+IHRnQETqtgeG
ieOgJnpdJAqvItgDedD11cSNOU4dnoVzEyDfqIbux8dYEscTsZrNSxkewR5IFFAS
GAohGsY19sq17HPM9rmv8IytIdWZUSYSwbUkxcnyALdmihJxaHelkvx4BlFuzV19
FItamYLzx2dXBN0cwyfaqkzKriinKJx5VNH3D7CLKVkoOP8iCtIhpvk9ZXt90i2K
/fjuXCv6NMpFzIQXnH+39ZfrolmYaVZzP8RtGX8cLsQbHedOM8OcizadK70UI/nu
UMcwLF6SlYDZ6rs1/tcduDR/Ai//helMRng3LSnaOzFd+gt9l1aZ/24nPsenRdWL
9ZSmueO9yaCkjP7h6+qySNZ5s5yRQt7rzoHI3iY5sFx/AlKdQf3CLR8WpjiG2kGx
opiFrI/lRfe7ZGcuQG/NlTkeWQEmCMlHTmidZrjqlXvAynuIZRPwj5Q1sYTZYcgU
Ine0tE+Xm/Oi7EfYnU1TEl9Q4jKK5lcVsAl3NSkTg+IvpYWyN4TZLYwIzCsO+B1c
WegY4TRLLhW8Dgl6C5x7PVpU5OSouK3U3LZ56a9rA7eD74C98Wy4glunsAnxCzz+
FnKIPPfVJxP1EdqwywNWqbobaa/H3cSKmSZy1WAtMQMqWYG+WE1V2FqxDXZKfHmb
V01JYjhyRqpGg2JIOohkPdMXJiSQUCBXEnzSk1LnMj5eMgHAnllLl9Hx+EWkj0SC
/13ysklj1v/5fzq3MzK/w/LdIoe6apFr8gejOFDHJic2q1kXoZmyS0Bu/OjUjAN5
SZimGDQHKipNtIbt19yeOS7MmTVcUyY7F9YtCoN8wswpWcunf5lplzP+awqFY7WK
tjBFTvJpa6BaNT7XvO3miZ6hJmrLDge/BKlWRdfrxI36RODElbc9Wi8zQsTC5eFi
rUVZD9ay7+pd57Ut2e5SKWj/HXVxF++e5nlRIlC4IRJhE2t23zoEB+WJWLhjUv/B
NMsLsZS2OGNPtgr7uU6ngt+AXLYWpSAJqJ6vSV0sEGwpmoh7vtZ0sLmJiu+8BgQM
SBR3wChtXzhp2ldQHfMZuW17Eyf/6clKEZALv59xtZKbRfOAol1rdLzEo7LMFZiO
nai15jgpwQmgFPbFgpRwpcxPbNDNy3KcozsUUSdaGFhlydWoHKy7EtCMoxc78g7u
JzSGfheeG16SvuMa0XdmhX7bZqEeAhedMO745I4D2cdQAuNyTiXPxnYBAclodeK9
0sGQiODGK83f2UYGi8qBZYusH7VM411eHDPLr/Cml6PHifzlOAswyMP2knX2+P37
XOUn4L3pC3h/6VaZhXggRi7gndEHTE97nfPjTr8buPctjs3VxEFDvT/1wJwhtQ6G
QWHk240BxwV7cYlfqOXmJpF3IXB8QICFSGSC0ue3NPF/GMq3LTJbC06Ou7wAY3pB
sJmnWXUoVPJuGonVL10dHKNyesCMJ0Q4VegfewRkQj/MEHSsPVFjakNU05pGB+F9
C0/j3uVYjDPp0MpAKHrdBkz2lJRbSVcDsUIEI1o2ILl/qvmpfmcYH4JUs+Yhvnk2
SCu+z1S8YPJlLf+t/WDIfnwtyYAXDH4YeytufV+Uy/w76oLp+UWSa0wMnn9kfUY2
5aMMJih7Ayl3TXXtF9VcHGFqrw4xoZ56MmBRPl9h3POSbVh88RBdPPdpIF2xr3P5
078cTSG8ZybRwqqRBK7zbI5GunMERluh5BczWUq9Gtw8JGTWTGmQ/4h58G9sAaP9
RlzC+3cwb0nmAxpVtq7OFnPvGMYXl6DcPY+L7RMje10586er+CCAUCzukTglxXQp
iBy3vt/cwBxQ87gR6dVqHMRFhTxpERhGdQTDl/zvptYrhdoinwgHg0NaEgaq9bnz
9x6H/v+Vcvu3djeZIw283590qvy8eFg836Eq5H3s0p/A1Jaw2PA3wzKai3fRqQ5n
z6TfmtwGPAoVoR3LqCmDMvQDmaesGXv+KmbcBwnniOlLSkfJ2Z0Is3Amw1MFRiQE
dJEIFEoJXSwFPVmjgPmggogSpgxKU9SLr4pi3Eif1DyvjpWSBMSkxWegD92u6bkA
f0zgyf5BYEbs1aM2TuPMF4brW9auFKiuKqk8r6WAb6//SmtVh2KDDLiXT/pr2/r8
xU1ULaTpKZRh1FBo5T+gytJQ6BhBWouo12UvnGipCfXunDdlSDW3AFs8i3Z03j0x
W7LJQ3c0niNxTNpGoyuC0UrGB35I4803uY81mSKxS9hNdKQTfYh+QDhOf6CjHCjq
SlDT8nNYCakrX8VYqY1PJuKub23AT0Aq6l/+EvMQ5pHmS28xdphR/RHl9xgMrcU8
xzLojzi0tU0X3NRdwp4LKjv4J2iLAQJ9jC3K5oUWtgiJQkh66QoKZ+QnqkXWTnM2
ZTXhITrDbWwQq2+xN6ouQu1p8lTauGoNJJrJeKU5++z59tkV7YKO/c6/ZzCVA6p7
j9f9U8/CNXieKhc7GT3t3qaNPqbNGm6hKc2VsnWA3iD0vRcudc+CG94RfW0avJl6
xSSOe1ypWiD1XO6C1tc27qdtWvt36XXVtYFmjXkBqANQM8FsOTQrSmayfg5N5eYf
GHzw/T5XHCD7DEWjF1RMCqQhIs3rqfXK5oxPBP6tFemMMRTPszIZXfvNIcsZP7WX
hNiHrUZ/BOaUbc3XCsOXomzpxX3aYQzPXgnMh6I7czsvT/j4fuBkIiCU5oFAGPNr
ighW5En6BBfU39/pLuqsLobH1Q6cxgbKyNgZPaq36nzvV8DksZZ2gxKAyLpdgMRf
3F2V38U7HnRQ6T/C1wIlMh5xOkzM97gA6ZNyk7ZICBeofBybOLHENrxDX+nh9qsM
x8JJYq1Lhs9J6AITjdUcnd69arhjPcHs4CJm/U6IMDXMzEnLcrh8MgSBK4KW7qb/
UAFE94/ISGD852a2UGs4YbvO32i8LymOdcjhgRo/i1hEyvyGi+R9R/2SkcIPUKoB
UMs7kGvd3+SEpPBGpt+Ooq4+K4rUbEqhrbxP2JabWdaIsGNby8ExFDc1C0vtcmvM
CGW0XTABFZFYeBpEtdbNv4mVrr8kkm4ExLPI2Gnua4newfdGHDDkTM3gRY6YHboa
OGMX4pI4orEqdTMWfDk5rmP8XOe1HyDLaRY5CdAgWrc+6VZsHFyCAHgItMWBcB3b
dwDYSTGJzW2uIYWLQPQ5lnvP+ZDNwmtH6SSgEXHh0ohp08uLEzfVT0I9OOs5xlE9
DMkyFx27OXnZ27YU2cW5NarxhdKJnEOiLUWpOW3lfmwWXUfWFuSRlqgOQYsfLciG
ejQEA0GThfLzgE/gZUtZ3ZHt3tq1MDh24OT3KsqYa7MIihVfWzz32PU0cFQ+heD+
lTE13CLG/UOmYaJX+/UCoE+jVODmwpKQLFJmrVac8amCLsDE5nU8YT73/U2poIeC
sw008KiiyjR3Hi/lkggDp49PvSi2AvguDRywnQ5QQq3wggbMStZgrJYwGhPKauDb
6Viba47q/SnNPlhlbmRXKDacID8zWPseC+KgLteFaL26eT1tasYVJWvx8PsVGwig
9uwEIDVOp8OuOQuyBegRvvJM5F7jcXmskeKFExZGhiCFDGuxg+utZd9WMetXmfw1
qw7+AnWIdhcDM38Cm1eWSPkLsUIzhPIZfV6nB3EIIILvdZvONaRi9pV/Xs2S9abQ
IP9GW/EfpHLY3aodNfZ2DIbqPNwqGaoB3nUdNppL3wAuMof2QbFFyXQgYQDfIi2l
ovswLR1yZGRVgCKwKCxQnXf0Xj0m4PLdWl4OPeDT/pZp16TVAuPAIzHQ+iQnETGQ
P7Uyeai842221yxiuz325dymO0DsBVEibfDYoqMyfj1OnFJdLtPgJFz6vB4uR3QN
a/zbgBv2DHFbyMhHlaAgl9l1jYapcrFFRFaBQe8ZsP3F+X6J+yz+6FKavZLxOMkO
mkZxYudTLg+LqkCU/5EaxV6OqL7HkkZ7BKjqP+ZBBfwwGOcLT4oBahiiPkxJoFu5
pQazmohrnSMyXW+3F5COssExL5dpr/siW7VmteD37BFiQWjMH9ZW1f4yEwieEWl1
AzT6qR2912Xw1Biw21mgJ9EQWGNEqMChLWfJxm9Qi7/R+sySAKqCDstI0W1sk9T4
zHmXQ9ZyrrQxDfGtBCrppx86G1ef4lwjP+A/giM70erKIkxejTMJRITJ5V6YT8wG
pQkz6jKedpp4QPrdX3uF+n8Ap4tGXd2bgSgWMGfFNUTP3V7Al9+m2Wt7a+8cVYZJ
E1KnPGPs+i9DcZdAuR6/61voQRvAap8QVqVV64/ErVdvASbAGAK2EOnLYmH0qZb4
3KthCv7gcpsSoBDFYLa3P49LrCQs1u5X2+GCFDi3ONDHKRJ6GNArW+pQANDZ+NlX
/EhgnwMxUkGgCA85LDFqN3h1xjjar8eNu901LByizseH+l1vURarVfMeAx3Bsvq8
/1SNbL7iwWGaxc2r3L/kOE2QrBG3bfdVvZdevvFsw+dqNDGaKDoHOlYDGAjL8P54
A83UQ/RUqAs2gH868XJpHDfmCWlTxVja8E3XrLx2StUwRQyP73YcoDFjs93P6SRd
FUzVBnGB/2pT5peAZ4DtnGkx655ERBdLLEN6wLoKrrqzv0df/mt8yKDKRMSDuK1Q
OJXeQfycKAhv3wrFO+P6oER9jYe9YedA/fiCNwf6vByZMytX9z96O5ignltdj8k/
L7dDWFkZHU/xfG6wiYlHs7gWYmzPUHzydMXjep9GbtA3aHqzYwUe6ZNHNS6cDRCw
wfsw+RwbGOh8zZAtFO2hKr2c9TGl57EZnPjrsES6myiMREiyiEoT2GGUv+XUAyHc
VfCDuR3FCAuPd24AmLyr/SOC91W4TJnnNd2Nku6t5nGnkGZACx/Y8hN7kh7nzhGM
huCe9/l2Qxt696fNPlBG6zUnMng+Lzayyy+wValPASiI/0uDJdGKFBeU4xsnEr1q
AHHjNK3gxUfaiUo/U1B06HKqAMBZHWmoz4Y125zTf6qVr8FlTTwIFz6X7gf8plb2
NP2XAj/ufjALXzDhRr6D1lnJbux5X6zRJnoELu9HYjKgTkC0w1t7i+KDbRO76DGC
OsJ4C3qmmv+y9Mv1SiZrFW8Sl5gpY6S8u8834JSXXJ6XHey1pGB8HD485my+5cXv
BIWS5G4uz8bfDBIosRni/N52CDL1B+6747vQKMPPQj488kZ8NaKSuMnzul71RO/6
k1hFTboZiRj/TKN0Q0AkU+qCYUsIUWOrHvu7SG5Ze0T+qndebUUbrasxfJ4moPA6
UzgQkWX+iZVydR+rwsHT/VFGUapnhPYI8C+Neo9rGVhK8gNAIQeyl0c0exzX8CDm
k6E+2KsZ1PBGX6LAyESiq1Srp5QAGwpNuNVJzB5sJwMMdFyf4j++r/sUkVN5cMLF
uc7kCv1PHRGTZ9mPi3wL/fLDlYC4WIqEv+LzQ93xRivPeo9++TSp92c4relkXnzA
dl5U4HLwueg2iC2fGFqFPv3mwsP3AHPD6XRS/bN8hQSX63RXiOtpoZAowLnF0FmR
vhLvRpSG67RJtX45PApNFoll+MfStf+OpcRa1k1cI8Z7lpQnJClNwuWP/ezXVUN5
RjXG4RzaQ7VacL1zFeQS2C+u9RbiFUGIFbo+MpvPUp+i3J4DwPDfxnq5FsMLa4h3
wim8/cxwiV2nHpRkR24DQi78lz4C+tuTYknhJ2WPfUTUE99uAPAGYNEamMBvBN5u
paSf8qarIVMBSZWkvlOMTDh0DfdL+7Hb4MRcmvbFyL2+ayO+CjuxdvQ1dlh1G5Q0
/HlhB6gl7tMFrUtkxwZZzLZ1jmBfAKNsM9oMrO+onGG8W2avrEqyENZs0VM5f0X7
7EiQ2i0ou5W3HiK+RN3UEKv4xPiNVRqSQwJNMSbkUvBItCAgWiWFtmX6FUnHqWzT
2SwGxJ0FIMx3h4nCicBaHYjnc3bsJlqQjzo8zEt0r7s8nwIz6Mh4ABtWCmt1zgau
nXFZ84k6LRGxb3aUxmSe19F2Fri8qYfM7XRGTWGQidA7i3PubMMom1LRqozANELZ
cnh5s8ZSE25ck5FiQRstqM+/yVCSIHmk4DduRjC7XoYchkhubgIn0l8RKE67PjM5
BjNqLxeB97E+8eO++4DLVZnZlKmcyD2kdC9sAtA1RPrqg1IDN25krqfHOgr/0upp
iPPQ1nBPQptit4gtcmPARX8/LwR+apass4JTA2c4DVW9oFxbbXXzt3+sFYcNtXBZ
Sfgq8s+W+wY1+pwplk7lRrYNuB0lflglu3GhJtvWeydr+lgMkWzJpFCuSRb/zDeo
AFL+P7psGFpvxMLvxQLdXFdYjBVb0yjg2W60SHAFU2UDEJInh4rWgIP5kBvaRrBw
//AK38fQ3KR/x4IxmMEteNKpqpfpFrsIBBCCNczru9ApBKcGtDmPpXcMLzDLPg9A
HF2C6t526/KpTqBKslfswvDJR/6Qpmlr48A55kW70vtrXoSU27HALwkkZMDwTyyr
XwAcaykBPkJyRITowCdMZ/0vdcc4ZVNJCbQ5dfi9c46DQD4fruMYmoob8sSNYa79
TUsG3o/MjBtW4fuPS/xxS2GGFORN63W5Zdwmit2OVGdg9mTBlzQm7R6vvCf1yFyU
4WK7ovbhhZlmh0Oe9U5tN+++vf0K8uXrX6AORNmzJI8tDeBzoPSrSgGHlZj5Dep5
OFH+YFkHuvf4ZfHa0WjjOuSdlJh1BpKnzOMRRCQWOBfVlSn5Auk3LWc+APmb+9jK
/pNEDe2bl7cr/idVJwMRR3kjUZd2EFwwNpqwsb3BbmqMHaIVnKUoWV9YSDJBqzql
F/WRLIMtQ3oyq3GktNozNgxgrLz/499rsc/LLnr5fOHo69FQxnelJGuBdeZoQw+t
IQWM4ZeXT4iMEzNIcKUuU6Wtu2B28TZXSe+PvPTeFkcFZqrZBI7qedZho8VjsPLT
cJPyDp+zRJa4zphh0rnxZQc0E9I0NY8Rcw77k7zAoqfh40agbP0CAODW/K1U3BLk
LrhboaAUTtd8VzN8F2NIhz+uyHmwYJLPnzSjfOtfFtVyhDZrziubkUEst4Wkcx9P
Bxo+fJPjFO0ANuYvpotkIg32NWpkfUIqVOLoDNpfMkZOyIYyfA8oodKuXj3HDn+y
4E1lzL5kWsKWWBCCnNfs2OhmgTXYhAXs9A436F1zDQGS/Pfm5dnBwCChTY/B3sfn
1nYs6zMOUZ5bi86sn+5NyYPM3muzn6iLIYTKxaqOULRYcROJlRMcK36oEMRZRk8L
xzxc4RTDq6o1oJHMjg7pe5TUUboQtnVkFpY6OB/nUjHY3c7rOL+O5Wn9IViObtYQ
FMzbHmHELF+YI8B1hsef6jyeW3rc/DgKjDfziYWdtoXOcNFbQkwuc0LGW7yGgb8F
CBSbJmTH9DJzcE2H7BhR+IsiB5NVZdFAX+q8T86m2lzdSi/u+mt7JAr2wrfhbtlb
GIrJ4Fyp1kTY0CxvOpo2q7LFJgg3S1OmmO8NneMJJXGKYNsSXkvwriEn4+gEZkYo
z7mP+3OgDdPOuzYm7OTC7Rnuhkp8jaeSO9sRRUrgLf1KevEmh+IkdMXP0BzXYgXO
PB3ZIunhoCU1XUYBViqN7jmj+p6EzqfTwJiGjOzX4SmKa700NlSdSS7vVXUqNjN/
G/f4OoLhDQXBVrZCTm1do+xO4bBRPhi/A0W/B4aAvHmpIO2Vf7UJUyDSlDI7D+w+
9XMZY3MYC/7NlX1KSZZ4oUqoMqtADnTlJYEJFVhjF2Xg0B4DiXOS1k3sC/8Vq/wW
viIzmeEr2D6viEEg2RBe5I9mLd7O/6erPNf6pSB41sPa6h6wNmiRnf8/JrMjZTSp
dyUeQhZzAPDEr2Knq1akQPvmA6SQ8BLr4vCaVM/tw1aZ2ZmcZJxIJstuuiBO5tGD
XG73tYN0XwuuwuyY8jZ8gJz2Tx39wQ8EvBlSBZylmTd5j+OG5kDEwQJld27Q9TWx
kNNWEYde820gEUxo0EkxfOFsEtitkus4fskqmzD890ETSDMtFYPvRLcKI+FQIC9y
h6LrvjowKklCGOc7bTp3Z93eKcyiX6Hnir/OtBnzp+XiiD9ILChLNrI3HLJYhgVE
dMkw2dok7z7r9COdMsLk9ApUwPKUddj7MWGDWSg0nmnFhlD1fmgpH3PrLsEqwmOY
8Jh5gZlgOglTMEEnDW4PQNOgCc/rVKUg15RnWwiAPe3c4aO9ao2GaTYNf6OkDGBs
buknVUvAH0OImETekTObqdgCfqtxrekTCB++uAn9564LNRoIGcwZH4WPVL480XR9
8QP/N+X8TWAxZvzsDgez9sK6KHl+DLQLKicbU9LKo4HhRPyirJN17a35byM6qqQ3
dkHL8FdAZWguGveIo/ftXp9uKpfhRZ559kJUkfjjQc9HwD+aZrc7haiW9JL41sv5
ra7tSZqwKOWj5hl39MBtJie0Mk0av5xKV265b6jiLqAi8N9+HK4A2hDqeAhJ0szC
BWsXv491uSm4IYAnP8HxEXLeytVdt+gCduePx45RsMIn4hDjhngNnQoQl+EJhG42
GOCz8UUeUtzO6w6r4XuwJVNXznai15kQc7n0azNTzXaYEzj37so7441MFsNSSk19
9wywEN/9nYlA+kgqM6dhDrJTSGnZxj8Z6eULti1NHGpicOt+aT4Xuzg74hfvpYOX
HM9Ebi78qMaic4mUWGidN6Fc+MB8UtKB5wIEvH3akCrgR2gaIr9Gj9WjbPBvKTeT
meufwjpqR5BzAiHHuKEIL0KlHiT3R8+/VQkAepzaBEOvHrU2SMO4006mlJ2eMVpg
Ip4slOkgpjtp4TmyztbsSXi1GRqQtIeTHYuLdrmd1stP34PHP6pNf9uiWISQnayw
ohicLEiNoapK3AEgUBSy6jcPwryHMwiMvsmzdglHMveUZcR8McL7KlE1Wb8BvScB
jt0V8JVML4HA4lG7c/Qd2m/l4pe32XhxTHM8UrTJ85sf47DqmYRfVzAIJnKAIXzc
lwt7RKEQBfjYrYZ8RXg+t5i9wyHf2o2jMwtyWNkcBrmIKSSYdAkDO4tiPO3+au6/
/SA7kLJb0QiYlL+1SmdcNMWbt6xgOmsLHaf561dElbjR34y+GBHtvrzj/hXrxvYo
rt+A5vZuj3JqtTkLgr9KOKTKa/dRJZmjh58tQ7MpIRd5GsE2++MwrUzvW6Bff1TN
iq8npwbYtA5grz2jSLhCxw3NbNGp1yZt6ssJHS2APfq7U/MVCrxSzlKopZqA4hyC
qaj1aBQiMm34RhhsgJf8Cgx47GgDQJTjnTuEuzzrhJzlBUJivO9MttvQy1JV7rQd
ZFfWtwvEJRplmFnMcMmNsH1/nNiphFDBMrck2p32VpuV7aBk55maKZwC/L19zCUJ
Z49fnVizz8NpxE17VrrdxVZfPPrIAg+NF1HqaLgMU9K/152a8cNUgeByCbEuDfpX
/M64+OTmLAZzxKgScHwGrN1I27h7LK4/x5ymmNeUw8jy+Umk6ZuqamOYp5b6aynD
uIwTN83O/xD/MUvA+5qu2vG4AaYhl6TZs8cu4ZH5Rr0idL4LhdcYLlVfBS2hOSR6
uySeYN6B9/0xm2pUed+LgLiSTmZAZonV8buXtVECiBwxg6Gsh3CV+NnuaM2Byrfk
S4OXZLWlxhAOfMQCr1yhWtNmw2K5J/thoHbEsQkmTdnZ9/GJbDRL10F+IKVB2NVf
GG5usSumjd4B0W8thDVH5FyWOdepG+80QMQCMbelBptw92VsLYkHmXIleidpoRBG
H8mBfum/B75+O+pmQkFZBcD6Tggf25UVbiJ7D9WSHmeGUvl3YdmSRCPWWrrhlhLY
tBE0nwqExi9m+UpEIu2Nmyk6j96hlu5vBP5c3gk0wzaSJpLNVGqbkoiQB7IUZM5e
LnvUtn9DKNG4uQoWgRrNtiVbz1OSb78Qxk1ogZJDMPnaA8A+uvk3F8lCZnqFLeJs
0AA9xQMGB2Qqiq5G//x/gpYUH8mw2C6y2TqDN+NMOD/0OLfOZEL4sMR+GhoSTie4
0FAqEp6/u56oNlleTmRrkC8A97Rp6V6cRanDVYjA/4RRBTb1sJksLHbxq2pLnHNP
RWYGQ1UXVYHQQhbWS4+MB7l9ULecx5RoHtv8GaOsVw3KS1rthdCI6tovN23RBXEN
IFWI+KkSY+CWektong6atJc/TX2A9VKzu6G6jS4XIsfh1VVP+zmwL8AOLUAxj914
WmgjhtrTKpiAsZ34mio1jnGOGhfrHn/+7XOGV+gy4D887XV8JUhvv0JNZlaDB8Yh
wE0VQ1Z4GrmIKfHjEDKvONDjAImMCIyaLz2wi7gmijSlgoRvz3i5i85CSKqboLml
yLNZTFceYgzLnarMj/wKs3OJs4tHXkSpYoWwi+cE8ZtZnYHz4x8veeaUni23q9/p
DCCCxE0Cu21/ErpCEOAiskbTggsOicnmsQGDX27xEpi/ReM+Bf+lBo9z1J6nZHq2
NwlAZa1JOHv4RqEOwZFK3aEuglTsFMoGyDubgM87EK3hj8iF07tyPWjiR+Eedkn6
z/TMFXukPgqZTvOAMMSlkCbhW5StqLkw0ZvZ786QG4UMDIp8ofUhzMOqgpA/bg9E
yXNVNddy4pJPTe80n8QllQ965VjHLCcEQWzV4/wXsFSsUGQr3DGXFM8jNcYUg54G
v8mjadD2yihg/9CBo+oxsNYLake++ASRqicI833jX/5Hqbm7gee+r4mJacWREJ5p
bK8MmfUguBqzjKDrltl7uiLip5YKauX1MgIE1z1dPCvxLwHrSEZWNtau9yNd1c6d
6wlpsxZJUnJuFrSTxoGOrbtdfdfxyEGDnnprL3kSRrkbSjwdZtJB9TQqxqLWv0KG
4e8KuD2Duw5PX/mpLdvW1tss+AyWO4lM5l/Itz04wggoT85tG4Vvn4ToWii6wtz6
ctT+lFwW8uz7DHaNgRdbDBB7Qy6TRuSK+Du0NKrNJJIzMF1MEEkZykPu8X5Lt+Ye
VmAp9MugGq18J0Wmq4lQzRFNYKSYtw+wb9yB3sA+mxcxpIPPwORagWZcRAMbh3IX
6HATRgCM8p8vF1QU7OHDqMtmRQC34lwyLPyPBeyI7uBBAZAqVaQalvyXwA+tNLns
6ZSW3aQGQdyo4/O3wLGc2NVkXPZ6ouNXE069E6w6DKAHktxW/nJIn5mfvjdvNSZv
KRFm1lmWXQEOzUhOZz8dGAzwdnNjJbS5ccnn4BP5QI3OPGTL6U/vU+R3uR9Q7yI9
vjLrZ96Jg3eJW5Yrnj6Iw2WFeZ0IOsL3sVS3WXKLQlkLyXfJ6+FOsqYW6DH0gL5/
f0hdBPwVj4F2qUAHjKQKvbi/QimTPkqbNklrRJjgx/k5hRrVBNioJNvgBfmR0zle
8ibmDpwTNAq2TELFge30EmxTSuSJLFrj1dDADNZzuQ6MK43ykUGGIThHkPzXj/Ha
LfPfJsK6HXsiYJxHpJimsGoyZ/KBsNazGEwOBUfpwQLkAkC1BmYtFnp1eGjcB3tN
MopMYqruV9RZAEAfoHfFixiSzPOhZwRHlMXVINoOuAtqXLgGrlGejfQ8D/ikRbQe
PkNXcHORqUv5dn1LTdtF+N+P7K/Di5yrHer610Talr3jPW1XrBPz0vhM8K8p4qMV
JLVw5B6S8c8yF+cv+SXQ1JEd52ctPCEGcX4rKyUuvNlXL0h8x8eK+CaNpc0WWUaT
GpIzc8kMoN0FJRAwimlXJRadcnUme1L/bQLOe2j9qt+91eSkVlcCvuEes3tkw83x
cdVoXK9GLSQeMl/qevqyIylEp4XmxKDi+PFtJgqIFNsnQxjufNnZapt3YQuX79ok
oEplCafK508a6LAX1iT4kGtxu8Ct504DJNiCiXPJpmRBgPy0H5164EXUzfI6uPnG
CX/NCsG9klpEngO6aaUpKg3aCAh8qD73vmeuCYMHxoGdTVtf5J06ozGj7LsddXM+
YRnFQ2aOfsUWzehlpZFocwa26UOuYGkuuqhWL2uKsMApGgLqB93U/nneeXahM20F
JVQtElGnmbVIw3sIVg1QTkkeFoh/IIMQW1880NQnO4c/5VTrrVJ/v1v41GXgME9Q
MrIb52MVu4JYUZtuP6FAzKHJIDY5UEU7xpYArPnxXWje3QZ50FNXx68o83dwMhKi
iNhAr0uLZNBJCZ1h7fHJD2qx5+Nlw42smihdn31NHLIkqKKhxiLKXdPnv8QoaBq0
F9gd7mVWuRjqoeChWVLRYmfCPTh+vVRmHSA5MumNUi0xHYUIulL4YP4F9jIFuh6v
bu+WhtypH3K18rDqsS0QYBL79bk2yN+c6VdoWieMUkdwcsPAI5v+GkRD4b7UpShy
iwrVl6UwcNEaQRrYVCKg/lS1xKLkYSYtS1ghKrMG13UV0V6Z8HhIS8PrmAuCA5ux
CoD4PBrRsGxayqxAxdDSw2W7k04bMOS25aipLz/3tisolYQ8VYSfuvHGFIa/GCYC
NgSevqlmnYnNUpWSC6gaMlFC0oqLM0uNO8ZW0nqvcEULiAFFzyzdSwhXV1PhAncu
E4BeVCvi5t2Wih0nwNKQf6q40wX7I+2IK0ashpyLzrU2kmDS2aMzjp38PjzYk+fX
1d4v1Q+AWi4CE9Ify1m3JsZkf2elCePSfioxsmVBE/2ACfsEgFmkdrKPbo57zHvi
RcMGOPRclVqeIBrgy4QnFz5M2eaXa7hvEv+Kq8buBVFnmCbZ6OCBGp5tEwfAux8u
kpTMxmF7gk8bIAOTCAfGxzr4xVC5dIvsWCnD5/aSbbONrTr1V5nV0idBOGwZALLR
eG/FMAtw1JscyT9TNdC31GYt3qjF4nMJYBYDBWfv7kD1CRYaqEAZlix+ETxDcNcV
HdEWuW7jrAKJZ5qnIJ3ub26NS2jKIRMN2/RjHCvqYJ6wGVAui+jgy+P4foXl0lLp
iqgNXHO9HwsnFeiq1/sJMSGCnIMTAEWk3prQ91KT9UxeWV9WuahhcEkgmZwkbOle
2NHMP11YP/ZIecZDzxN7Vy2c3+Qso9jFfk94rxMaP/Q2J3M3zS3qziIbI7uzzJCh
/H3BFJF3hWqSn/Hvd1cMytNBp1X8Fxesh3VhTsfJhKLB85o0gI5SDiE4ppdlFcjZ
6o+GeWEBgG0MlfbFckK4tDdUNRWhof4GWQe0msKFbtHTTbHkcpzI4t8j08NZxmAC
jyYg8yc2AmyiIEisKbEzzUKXwR+/Ai3zNNhqj6P3vjsyd1lnRMSOsn/L1nnV9OEH
PKtyLWP5YmeNc3hJsMmSmxU3UK7VQJ/SVCpmANOcu37IXiQfAjp0hna9d6cUoNZv
mdWWMTsRhIN8v08ll6ACWTZfK10oBLa9eAM8lXcKAbJT5kiKrgDskJbQ0AZ+pJgn
4QwWR5dj9xwMkpvYYBhO8VTv7tiXkp79yqZOTSH8HhviObY6Z//RNx4avQNITrPg
7gMo87x9e7ujxWZn8Ru9OqDwr1pVeZktFGhRG9nprGfQaIE5L2WhbLXvmvIgFFa/
5EBukAOewmTWQ/H98XiuyU+cA1B4Vn/qipq63VHtDwDcM3yl7pmIEbMXuu/wUySU
Cid7XPJRHZOYSv+o2UTAlhR7XwzPb8qS/GqM9mnpuV3BB/nkF3d49hNIVvLZEnKB
wkRovR8kHJSAqQbTq0dBvJYRPMEivq2jTGC8rVlrveUUkFlpkPn5ZM56gmEawXtU
38irnxEGjdyxwnYDtYRiu7nPramAebmISEZNOC2ew9av6ONi0bISJ28SeYei2gFP
3WetO73bnN6TApXA++TEcCjAi5kdn3/4xDsIQBeAtb+1uuQNlexbUCJNd5wCauGA
RV2u5fpzJ2tvk49QL3Oy47eQ7+uRfI10B1wpnLhE9WWA66/h2yeRf35ADbhdmOg7
WifsFMSGndzvV2Sr6yhgLAC6GjBxbRDWwFp4Sxtx12KTqciWAhduD+vtQWzfpJuW
xsINg19ebKZ90bF8TmnXOCsI4vC7zsNWDIBFtp35LRTVyiC/7c5utobz9qIVOAqb
DBIiKNXfwfy2lvLL0dDefw8hbTDkZZ4qWN9ymj57bvTnnI628S1enIdUj7aZQK6S
3ckTGRqS0YMmDI6MD7GvsbcEfcWxp2YWCbAQ9xJU31AuyNhHBdCibGhxkT/1bCsd
6zg0FIq8eW1bEi5bMuKIHltG57Yu064Uo/gtLQ3E/Layzh3CgZg4ghDXrbzVD042
2tfdEX+X4HiSUxc1bb9L9NMi7wtxfOYsHvXyFI6vNjocpHad/YGgAkbYOdRHgtQM
j8aqX6RCj4ii3rrIWIDEUGSOTweOzKWA5leObCf1R47RqF2c5NE55rPou8GpqaXl
W8Hc1F/10Q7zPqkq2a8sZCoI1UBxLC4sjkbuoaRWGBaZstYPvTUqxO48gtQVWrYp
f8YF9wDnS3tlNi09oxwwqVGRmkvkrHSk7ZdvMD6V4PT3VH33osSBoU8YW0ThzP9N
D3nypaSUQIogPRyVfpN05Hp4zW8+7bCGWnbZGci4tTfqcw2X1gHRMs+n8Od16Kez
hlEdS+cy3Y4UT+1pFc3Th1yweJM36QV0Bxesvg/lo4F/BQJMtPuPCiUKk0XmGYPh
VUG9B+3uatpwiMND6qIEoFxvZW9f7sNVQDiedO4fUENAhbBkzCSjxUt4x8QQELGL
FIuziBzuJeh2uEVP5BSOUBeyq+ZovbxLVqyOtq+xZBYdIA/U2YaFI5l4GOANyvdI
q/iTqBIlGthxSpRp5MaN5RcS3C9vfVMzKJLAp+X7O8/PQ13tjCjhvUddnHiemZlC
BbuyslMRRw9J45bMt6T8P5nuoOF3lCE4jB5xQIOohaPxopwTja/98KCsNDD+WuRO
3r+h8UoFgPgUJCI5wl/P8mDC3H07h7zWX5b36orBJTWRzOHxWaCtUJd8jXTDqgnB
uAgmAQagITppkMeqIcWwZD2ROLAOaCzU6PEm097Fe6YDSWW9U7AaQdfbpYGT+HpI
Tl7MvYfMrnaZ0BanYFcCpvVQ/wTESE98yg45JS3o7pjCAj3KhjKUWrPDslbBTIXK
l0KRz3uFnZ/YbJz7/j39rjyHguFWRFMVdtLF5eEKrVvpG2kahZKg0dPPGd4QhYXr
cOrBI4KMjcVBbJemxOC5rx+TqegLp0a28BAM4QIkFi7GYa67GUMR3+LJCghzSlfX
S+wZfVXMmRF/wA1kV+I1uMJyoE8bUp9JtqYlWgQRaDKDwx1Vbk99oHBfX+oy2LC+
mTWK46QdxVawJVmbxMwakfYKEy5+rDcsBFKjiA6ud4Tp/xTyQ6G9FKLBIsb3Bgr+
54YBIrxS+OGh8FiNWXoji/3nR+zcv7G8Syb2KBXZpWchjD0qGW1Us+pEBOPM3pIb
dFNIkZRXbGl6DcgZkobBScZTT9Sg2pTAAqULpKHLRMpvXzzUHs2JicEVsA2Cq372
lSB3TrrdEc3Ri8tHaYuJJdCCcuWVcKB/B0GDMxc3IhbMPtU/lWsrlX80WT94QURr
rsyrMMIg/ju22zhZJuKRQoAIAEo5LV8IbEOE2hXgiUz8IOA0ZKl159+RxG9Y5mov
f8aHtBSxs2rZJb10xoShS0l+TB6hvi3nf3b/95nZXRZVF16zw5vvmQSFdVSJMrSs
BE3WOwuEOWwsxpzuY4M2KMgpROze4CjlrnQp0PR3Pa3d1GaVX0CYnQJryt1MVV4S
caOR3ambZYG1OXKYKHa1HwbGyzbcLtn0cgpvUL5uqyYuPw1DQ/8sjmi6g48IOkNG
XIsDNHCjde7hc2M7OS+xYmFYnXKr3cfh2RKc8atiNzKcge2anZQWE27Y9NfJe1/f
0FFzGcpgwusJiauMaq/V/0fhhFmfLc9epoWx2AxzoekR0fFqjfwRIaLLIPqAU6bk
+GEhGaJ2LYbA6rf8cF7/t+Ayz/AADAK43qCs6UyJrFu4KS7nw7ADcJWGKFDqetOh
9qV9f9w2sNvdqoCDcCQe2ll3c1WjFw2gygq45y011nqZ7ZhEZ5jKvTBtUMeHDPv5
18xcqEzgHnIeXI+39IcYVwf6S6sL/PeBkPBeoUoGC6EoWgvx3+lL5T0yYlvVLgV0
zoCGbWja7ZzagvnxwMIdbAEB349cI+GstyUyRLNlN0GtYgjM7jikgZB+EB9tC0b6
sW2thvQw0Feh69duFtXBISqBfZSfy+TqTZ+s47Gv9nO8C87asFAGw9384PRNfy+H
PsangQmeFLTOTRTcOpWC71VXqfo2WNscEu8hVnZWWKlfzBWwNm6JROy3p4J8U+cP
Hv4gcMOZOP6IPECJVtP2cG44HQ7K7U0KayqBx/XBCTAjgypxcxYoHnWUnKS/kS4K
r55Unf56MRGIGqhs3tJZICBqHLM7Nl3QE5CPXkW0RA6E/SseUGEwutIGe9wnLYAY
Pj02xKQ5NJjIo96JKLvHCQSw56cWN59aByGicV4G5U99AIv7r3b5SL0cVogW/hS9
to7hwBS3FbvMgUIqFAIzXYtaY+5FQPIjrC4ZDDjZj2EJ/JcY9cq1WRpcyYAC6crr
ZHFvz8Ecumofnt76uR8+MQ5ZUeFF1oOV2LpBHnVACcmIMuP0VHYg1p3s1QnbNXna
alu/7eDFKoIdktlrMTn0ZY0MMvOtYxaNAIgmw78rO91Qx4rDQzzN5FYjn7+gpIPD
blR9xfyBoxzw0h8bKpNONiaYQG7X4VdbWRMdULfErNXE900TnCzW27kJ8bJg9K6a
gi4ha+xrRl+7M2hnRmero7BUI9OW1ih0EHwrdF9Cv/pLDuSgGFyEk/UZDFHeORe9
ORj9bll7pV8nAA1RZ36oGWe4wtsjQmcDzGaKR3nD3z3WMOSuO1xZtFA0VODbz5Xw
dftqcT1IC34aKKV8I3rNSTx+IitwROLFnOMCZtIm459XC1wS4ePkTzcuqCVTpT6B
DlLRq52YEebRGayZKvjWGfUoZiM0paWIyRBkuku4xoEXKw8GY6YN01TzB4/FZzdn
T8UyvZsAnVTN4Im5YYfX8vNtKYQEp5akFiLVquosK7MuwtZ/H57mxINlgdnufjAA
5tn58E/fuIPm5PpEdG+o/bGlt3g2HRiXZsFgW5lbTdNKzJ89ZNa7GhtEHtt6Mv6p
e2G2AurxepWcg8EPjvjgcYuUuCYFiaXjPG3cVqWNu+ro8ZVZJ7c+u7FeN6ooEqLC
Krrz9JlDg8q/tXRNxf1fSiD4kpNnpVUtZsWiu3K8/mE6bAgQoJwJSle8WUp3T9Ld
al/3lsKx4FDpgEu8Eh79Qlx3y7npkcoG/9k9Fkvhkt5EMGsRjn3gfF0/LrvKGH0e
7aVqxd0IXapAbVNbrB6Pnb97Q7wHe2jozcY6Bp1FPxkaKuoEHLnMWoBy1mtzziXT
Kw+HVktuXPU57yfzLA3wOkhjsdJGNxvT3mgTu7XUXnWedISMqcbOUYlbHROr1XiT
s3XMKUW0CqIkfI7NzguoYM77E4DMiq1VQvgcayeN1so1MyyuMhuZgZVmR18CbjPl
YarphYIHnmHCxTUgE03hPTYIVfRmeQ+c/oPi4zVblzRH9zQVgbbIdK17owBIpD1G
DrLvcEo9d1/BIt8klrfe9f0j6+6gBg6ej/wb36oBVMbFWD7PfTPc3t+vHQkKGH48
Qbq8PXuS7AEdcCsbhEWTvNG5raGTzPdkI9xSsvc869pUkoF2nfccHEB9eojXy7ke
0xL6LZ0V7jdRgR4ZZWd3bcpLALOKF0G3wmHALao/g0f5YnFXfJ5D4b3PwR7QsFe8
cPYFEq9p7WDOUKGoEOk6L0c2jg1Z677ZKWula/1/p13xOA/0n70mNQSyVbpsc9h1
oCO4TgPG2BZBPHiiiImdyUV3ufDJDQZpBh5L5UOQ5o2NB/XoN4q1PJ2HfIY/D4vP
YOQ6KLy85XdwH9W/ICDSZRp5Z6763JovkwQj6IO8nKZV7JTGyPrm8mligW+te17h
h79UBdYF49U8dT3v6CRDAfQ2kSsREKPxhXX6lecZgKyxls9FmKzyqzhiJ5oeRNzw
Dcr7sqMAgKUlI/FN/ol9jyf6KjpFz8BF4+2LRJLYxwmOUI36EPQSwSoDQtLa92YE
KcP80KKeDQFNbxeSy+9mYk5l+CT1KmIqZXogAri8x+cdXcWHQoIsHm/ooMV7Qto3
4mSoNwEf72xuDMZN3j9JNWZYHCVkFhGigExgYSXQSxQtDfAp9MnuNM8WI7L34kXj
iCjikSOy/PzmlZXK69+pvMCfM0oe0ZsbcsgLMAki2qMDPAMgtosIohckbXgZucnU
X1UrcIA1Qw2y/TlGPAqptrl3lRdCqvC6nIE3sXq1wHo42VpCKRDakYu3SlejyUZg
E66dSXXslLzXjK47h99xEiuGzpsJ1VP44SFpxV8C6Fdx3KEEM+wIVTr4ZKkXMgC7
GHgtWlzkyVvMF7nt5W/SdUyhcv/5WrNqT15mDA/ngkXJm6PrGMNsw0cWjB07ZNAy
wQwElls/no9V9gpjrBMGzxQFuQ7Beo4uUdwyHmuUB+YhtdWRxMbGNY8uHrqbxOco
ltLsFN5NWzfn7aHWKJ9hLI+U/fAdqDLsH1EpTJOivP4Ev09VglE7hwCcaEpFcRU0
Om0VLZG38fkaEZDXrSE0j/mCjqvFC77CG2Pue+GEFi2uyZKwxkRLTotHxmF+dAbC
HPsUPWLtRfn0wkarwtVtIu2IupDO8a7hokN4QrF5Q4JBKpLTkPPfysjbD7o5zNst
Zr9cJ6c+oorSvuKnvFWsQx8VhdkqxreZPsRkB2ckdEWkGGpyl+c5vqdJt0JPTrpM
acPLbbTGAR05YOpgtmR9WJ2VAKKYjlDIgafGhRbnKW3V+Brb4Oo1NpUtgE9pdlTT
rc66En4baIpArsu6Fy42nQN6kkS0PNiU4rkCCbhTjaUJWPy4zUF/4n0yr00GouEY
HVsg+OZehASMzFrzc/AkaHBcs2aacjPuarFIHQ14mg21wNPxugpcH05wK7jLv10d
6nBhMUlRoJjMuo/qeuoOo65sGzP0fhSfapGcPPrGaa/xS+FgbZ9P7waNEuWDsDxU
WkaS5YpEUj3qwfIBIvd59Fs9Gyic0KMLtbA/BgvUoi4U2RNwNwie5Of3RSjLn/8q
UwnlXxf9BJqOY/OWBahgf53xeanOwqF1Iw8dgnfGKMLuzwlWrcGrRmi4w2n4SXEK
HK34y4stzfrv+F6CxA5NRRKg+mS22LNSRXEy412oVSUW1FjiizXHcKAOjcTmDozY
LRROP9pgLR1T0DN61k76Vm3e55plchNFODyLbu5HDz112AMmZbNp75zEDdIEQhpH
d8qxKc/w4g/D9ehKy4jHoXHeRShN44tC4JxGxirUGnbA7sh/XQOzTJPBdXxINFnp
31PKK3FC2RnW8LaeOo2hZ8NIPthorXQR/LEtLEsx4y9KemAlj2u3Cx6P7D03nSgg
BX19ZLdgjkYNIHsNvcsgYPwCCWCRWMIFUr+EQrlbd5YUoq/h0/y6mfE+35GRGuEz
OhK5gkQbhPTxZTUm1icE/P/dcsBtcLfyExRaXkWe0PP6SAM3WSH5x2rgr0B+pWrg
flgojVhvMBnD7oiHzqt7byL1HKasLlyD82JCUScEXDAKKdTi9Av3F7PakDWTjXiF
n9tJh3mmA/hl9TPaIGRr/Aw+jkeHUAPQ6A8FuGT1gGWkbewEl0MJ08CoBMXHTmOb
uHekYkNk7BKTxjblHSyVUiF4MZvDbLHEeKZH1PfnnFxy5oIdZr/70MsMH7vXziGV
XZYO44d+KikvqUtfZot1HCsU9gikAZ5DH3FbMCL0HQKIoY7fH5zotZKDXPKOu86s
YmSUG2G4AW3zsbBmtBGOZFplocqg/2TIzmyWW9xVsTEad/DHj+zfrWrXyYpIdCie
GowuWpPDgTqORZs0+Ogqklya0zsUUL/NQbfb+LJK5b0QOVy8daeeFhl1BxO3RhyO
3Q3527RxKfCSMlElHbBJCghtRx9K4XxpQ/V/FnDg1w3jaE2XcMMkOFTfwdeZ6Lkz
56HHfuZpu6q98gZ3cswfdxBJTvsN2hIiKJPTBPCY+8nVAvOg+7DCRRUHDzWGUw9L
0/kYgJL2PlElbb/u3sIFUMRbCVFkKPWuCX0nRMvg0AGS9FTKd3L/cr/HUgCc6gWZ
t60x66O+MKfHHi015/D7EZHETSJMl+CfKTSPzsLcWu86L0rgQzyQyGllCWLu6/d1
aWa/OdjBaARXDeX+z2NvwjCIC316DMmAF0gH+FbkOxffFfHk49dbozzFo9EZX9tr
5pySNhO7Yp4yFThk9zHyBMgzR5jl2SKxj0Nsn4iqC4z1f9VOtjigNrNIznR8U4Qi
Mmrtckyd1QwBB6LhUT4A20l4r/40LKanlCKKPl1V/j0xG81XWQHSt48b0w81QWvn
Ekhh5+crMNimjoSkkryyBv75Lht7x0THgGGi0AvwHv4UNgHBDkGBXX/8hWRaghzO
9AC+Znzj2S0Mp+ry5oMP81HKJQ2nzLODg9aUNxAPxdSPVgZoHwJITk4Lg9R+3Afg
GDtkl9R2ycPBMmLdJv6+BphjaPJpvhu+I4wlrHV2/iZGoZIBVkgHiTfASwsGObt/
7WsTqi2iAy7Do3lSR0zYggk/3P5xw0XCM7Oj9M8Lko1ejaprs5BMp1ZXfnGrHkk1
UYWOp9KPqyW7wvDKXGreJtp/NHWyCurQufAptmBCUplY9sqy/BHA/usabneqOLwe
KIFLHQLzb2mze4XjvDTD4XlmXXNayRIlfjSzOV+o8dS+M4svfXdX9tzRDWqzMOzC
xkRe8Y0L+la9euQ/+wrAYu9a/U1NeI57VC1I84TiTIIskF6hUkD5NUozGFV3zpL1
bze6p/cruD58eBsn3AQJsHQ8BVIgwIyn9dBEXz7oM9GIXClygctNuLBLKrtF+SVS
+70te3qnAfG5EjcCWp2M9iHe+a1iTpX2LoyQ0rSgNr0EAeYDEZeMYABcqcavxZvp
RatPN/cRI6sawNfJmXrjSsIBudAFzuFgb+2OHITLPs+Gnm4vFFLKVe9KvpgaRI4D
t2JXAa4mp3KwzgiLhCdjGMEEP/uMDptuJ8thewrAzVfOOnxfeYUQPyffDewzgygZ
OnQLKKqgOQKbyI103RLY93EqTdusVGj8OI66UmtRrKKM/VWd8yRW3dsn+gJ4Q5K8
Bob8PImBTsYlHYYsyh4PxXuW3yvdISSfWuel+b+R5GDx/jTW6zFN1+35lxlrov+4
J/nboT+CWtusPxIZnPQ7jZjZwHEOyN0EhVfvA6H4C1hNIdLf9UK7qsSSUSOTOKgB
/5t2ugWAVSAC1SzynMFdhEgIGXKEYk+HtMQLWNa7TIQG4bKxOXgpvx1BkGMxNZMF
jbyR3LK0sxXwoPXA6mZF1Lva5UerIXJO95ZFnyTI4gV6fb19awYDzrPv3KwlsJ1x
W7f6lkHkooD1mIffIVvMsnS6Ef/CkiKzRIUOkkdTUaAG6YU9iuGYCgeNXdYoyANj
pXwtoBSc8ZWIrMLJwZKJt0eXCisl0W+RY1zxXdHa1EA5qgNQfOxynXaQXkNbwhXU
N9DtzAK+78pdF6xigDDJYivNx6kGlUROxBS3wygYpqc47tIphx7+WaGQUmTNSzfB
G/0qSLI9tKLDgWbMPhkLT+gToR4xFlNlScvwnexOvrrJu3+f26SEg/l0jKlNfjMx
jPUYYFzpDI/Pqw7k8eU8zO+hlr7IJ+4qu3OyHX5ssTpEHq4U4Ot25E3VcuXT/gk7
fqZsWR04gdIpVFThLQ8I3kqgk1G8csfkoHNB4gH4EAsVKQKAQw+OqGJHtCipVxtT
TPJXulQIa5Qi3p/8hJZzTHJ+ym+nhhpC5KzzuUKtzyol42uwqhX3RjZJq3YVu4Gr
7S7L672+LLSH+rbRojt0LsbY/+WpHphRykIcxJJwhnxiuvLq3cwlH10ZLZbLmDT3
uREidKzDL3jYZjQ2eFFKM6S4PHDrQlw26MtYLUhkQcL9B1OELx6zHuVvc3WwlnhH
TMMAyoZk8z+8GbqQ1/DX9x4RTqtA95Tgxen0rIjtGSjYLtV20zG8TrYBXkr2YK+I
9jVCPKia5sq7Ut3uBMTug0O9gU3XGGBK2n90xxbHXdKDOyb/DVivb/kunfrvU452
M+M0De6qsO5N7YIB08bzMQZpc6WBWrWL4qd66v+4ozL2d3UOV+UxiX3Z26yujzQh
g/rcn5OdIDqYAhgnonHDHf8MhZsTid2Nhw3c076YGbC4aOOGXszNuM9bPRr2sY9P
i2VKTTkJUVuH7uEpDTjrC6RBGHlgQGY3YXJdo4aSIMuVN3Sq9MBWhACXFKxjh1bR
9nwuTNtjN9d2K1uKytyXHbtM/Gb1VCV5cSgYm27ZfVx9NfsHYYAeve7FTb47AOuP
EpTJdEMlq16vzar6yomfskiDzGQvgiOCwR+XybLfAJIJ+HE0CgXjHKuOMvqw4L30
GvPZnc1lXy8zmJy+Sjmzo8F9GCTenGLqNKAdVc/JY8zBWz7FZEXJqGclAwi76WNn
+6QlEZROvebJ0NA09W6oQDGaRv3AwuP6JugL4lMG/7Vf8lP7mMNDDwxrTBq8mlmH
zYbZi6KqeaZ3SXOoHQn9VJ5mTNOeE65cVUOYKSUOwFcVPI0WddeS62zwrNPQTZB1
4oMwi4BHO+CIlL+6z2exVIrubnM4apshbD/pXFJ2GJEqtI4h+J3vRQ7OEdrExdR+
o6+Ux1PRgf674vcypWwPWeWlx3xzLIlQNnBnpZKHQn+RpqnJIIOYKdzqcYUdyfus
L3YUfnhJcI2k7xoRIXm9cjDH7odrc0B91EIu/f8gKbCyXFgcZPelotCJS1Mt4rpa
AldQx1s+K5Yb6qBOGaOPGSWyt2YvM/ibA7Ma/dDWiXlJOpQpDbaZM+atRJRNpOQd
7SYWNCj2b5gXC7S2KJnDN6uWES2kpmhJh2jxJuse14ZBMYTWedv9i33BpCbnnR0y
pPri56IQo8CF0g02DBX39CjpYvsKorexSfJKhXOfx4KxK33TltiFw/9fcgY/Q4HH
/zeRN2L9xO77mLzZLwjON/3IidTuftzHasg26DnbsBxZazvgRZvH89loHA9SUrBv
2ZQ3uJg6NAL/KOJzJVjcwO+7bJThLuN8OXrXj0+OvvAOmIVzeY5am1o15HAiGwyb
v81qRGmEyYFviy36jrLmXeovrxWRB01HKvmIaSFXPvU12l/SS59n3DzPud2TRioV
q6cAjfgRJXQFLyUWDbv7I9DRzfjnD3LzvOVIPDja7NdMxkrSALgyzHAG3uLAql0B
rlGS+ZC7dkkeybda04GjhCkLemhUSbVXK/wsM8wkrzeAglgOHkO0Nt4q8ZqjZ8fp
ouObQ2sIOxiv1VaDeITmuyWsLRyiPlOzASNp94GpVKLwdKLTbY0Ue1qewx5IPKHP
vPHnGV4uBSLjwNqu0wooEM0Ghy6CbNs/IplDUKFt3tgveQFRT3+cR/d+TMetcPqE
bO5TRBlzlMVgSq7BijRH8qjcb5n/BkvlT4ZfeEhHHZ1pYcPMqsut2G64uD9Lw4SR
JHSi6pd+Xas8cdgSsojgg/R/XRqBLend8QCVNSkzGG9LrP+H1gR4uxOf7bo/e9/H
fYK/4ORVglrGMxnOwaDK22sJwr689Kk3TJGYxys0Te91xJASAvR6nI122+lpbsSA
qjZVz+P9xIVHWU3KPbVmLp5RDeBvQEe3idOJ7c4j70OK2QkPyGG2+Z/JhFsxBDLw
a/Rp+44pKcadmBANUq+pmC6wsZh2r9K7pyQRfYgHvAGzTGN+klLI3IN/ZAki3jSF
TLGnHXFP83fd/b1xq49GSxINSC0dxIAEcyP47W+HNkkLqZSUviMfHph1ap+wS1w9
udbiAgeJS4RARDteDqb/arOQN3VvxtMlJOMuhP+xVYhUlLApnWMAT/up35M6RNUy
QuW7qVI4VZNAKEsjp9ojPsqfDsRGBf8ilRTKO3mGCRc9VvAydYC/8heTR5XcRkH+
5BdSqkks7yeOh+5kVjJk0/tclgu4qGa724S+L5pkwLcxx2WokYJ1eRKq1zqmE62x
PmFQPC4n4su8f9PWTqMQ11iUkw13BVXTn+CHVZTm0hZHE//Mbn5mJc62ne7c5U1P
j0WY/RffL2hjx/01/UD8YGR1Sm1Ue9BA4pnpLQvoC397DvO1K76bihLdSMNRofzB
dA+HeTDkiMkeU9Mrrixqna5o1UBW5HUx3hfQEFlJLzNitgq65zKILmC28bbxCv9r
t3KnmqD8jbUu/SeqSgZszAfExHI0tj7wLwn/7x7BtQ5Lh5KonHHzOZDQ6Q/WeoBz
2DV4vPXihED98VvgN4vTlvIgEAF8rcl0rGX/ZKUcqi92tIif8m4xYrvV23VyIUxd
tU9azYRVCTQRgOjF34azxBnl39addrdzJTSyRDfN6UNPLWEdAkOIjbApD/KwlxIE
mPs3GIZLqtNJUsbaHEDMpxhWqCvQCoBDwKxKgyahcBdUvH+FTaUnU2jM+Gx8+uxv
0Gb1hf4ejOhddAtk8XE3J2GfvGL7cbbtkbcWzweTto5nNJUe4KCZZGiSzNFnUEAp
H6tIdRSK0UoqDuDHnI8ljiBwII0lGa+ER1Zp5cXT4tfpCYZ3dtrUlhDTvBs0uGp5
FfJYwmGpDkrrTZJbHq6sybqPH/Oz5z8a/XNJY16Qn3+k2a7AgpEuLt3psEuh8qz1
SI0ewPAZoLW3MPlPtwQTiJN8fUKIBM6eddo65P/MH5vhLjIOpdd5YNept3lhO7ef
XmPZN7UrV3RL6HwVqGd6vabpoep81epzeIACEvATQqdVGxqweRc+FJLlRZAfXjTa
OfvEUD/LONTT9E2qMH9jmSecbcX4IYUsfnF1euzjtou30cXiltw6J8/SnDH3GKjx
/elwEbqGUrQe9SHBJdnlhzHWHZHclqkKaSkAhGtgkKAk4jtWPGmabyaL1fxHbFGU
ejkeaPDRafYU5VHvpY/vpixza0pHf2Uu10iP4SkWI5CeQ6j2m7kf4iYThhmXhmFg
3T7vbU07MjTxhax0Kdzx/qBb93kS074Pbw+S+OYrHe8waZiCtVI6aMWr0JtPvQyh
Dz2SexsxAlD7pPjtM3czLT+Jmys6zKLkxO68wOwdaS7k/LsjcxuZP6PNA5EMgxZV
79QQXs8MSIFbYb4Pcf3mfpWfwS7XRlBvxycCjUCIQu3wGVlp2t5j7WlieDA0A390
Hwbd+NdON8niDC8N9C2FvxybmhvAWZKWexjF/KMuzAbpU+lSLefO76t8VQsW+xhT
vpQ17yGpwR3U+TCr+ahpV3+qcBBDoJmVG2UmPD/Fp5Z2zGlfF2S1SlQKrdu4/U1I
dyccYX4LN2jcZnygD525SgjSyt/5UXm1BT6fzgtvTFDJ9Jdbr38wFSepuDoQni0W
XBxtd2qZE0dyHvWMXq67z9tb4CJ02YwwI/Eqh2XBIvtIag9z3jrWKK/IqaEUbI80
upY5nhLcoV073JHWVNc0K5qLw/6st+HsM77rH6RZCVgdNrz6Q44T9Xcs00EUmjxL
G+8qhA8eOlG0FLLOsRC31X8PY9xGVIgKD6nep+oHk2YbstTlxSoHhizfURNhd55k
z203+Gc6tzh6eka/8avEgSF64sJAkB0XK0W4fFM+5+pQnCBibBvMs/OHsjptB47b
V2Ns2nsT2aSokEYBBDM1EYUyJiyGwqERjYYBk4aO8PXGJ6kVW/0e1CfILz+gTpV2
T10UqPkLKfJIF/ZbyGbnEWUGgTqrsGbBKABInrngwNyhvnhefOnMR3U0ImnBfEHX
q8D1NnHIiHXHueO3nC0UjFEHowsvZ+qSL17sVdmJQZ2MOG1ZpgahT8Rmm9AFu7VM
rfjO6+vEX9Ko3cUw8u4r+iwanxcbMuyAC4j5OmmOVn5gmGpI/q/DtWGhLm9x6Olu
w/RDEXSVr7qa4Eh6tKHvyhHEg5eG7cpzjCuCzpkdD3G4fHimhzSes3IfR5MiLByW
DW5vKlRJ3hLnYS7WivTKQnmvRk6zgRee9wzEHKNGEEzlAHKgBDwrU2XXR1TUm55J
8fwMsV8R/Yhg8IoZqa+Iy8YzcrjbkWSBkvF8lr5dOIAxBxpDjC5+V8F3rt2TBNjZ
NlIaunNE9MQRIVtMTX5FhcDARer3xZkUaZL9jCEKzGTGDFZYlGxcn1fAWMJdIvy5
lXCgSYCL3sSL5HuA2uW+USbaM9M2fi0MCl6s25sjBxNvTUIPzgnafnaMiUJIal63
zgp7XFNJIyhUgZfXx51zF1SfOIsyo34lRUq2K8125mdnWDs+aPaLUKiH8OLoyIGj
ugsEqEDPwGISeE+qyQ4Il5yFUswXMO6F/4jYgfzAqSkRJMnPsGZQTVv1KA8g5mjg
1DjWP7Hq5HmesvhWr4Mtfyl8pxf297lDPx9krPPTBaDHPDTzx3yCVHb48/Asc2S3
rLndZe6Vk7FGv1smLbjlrvkJYO2t26Hs6t7YLWTSTeKrPt/MaqwFyE+PGoR/ArWx
+3U0swduWqrLoAGFg2ZA3tjAfzN9110f/nAOuzlczUT4rhBqF/XqjTu0mTm0DBXJ
7ubavEqVnrq36bKS5aR9uNPxT2Ewzwt6hUAFY874QZoZdWZ8dYbyzqgsJbVrISzr
tKuNhfH+zHSwSfmVo7l6HTSyv5VHso0hxYTKEIFtrGZx6Rh1hRPZfL6sDqLH7Xr5
ME+CeThjQuy1vobefv5/8zyMuZ14rIkNSm6R7T1SS1Lb9NRx2/RXO5HjSoxviwBI
BsFOh3EFjYQdi8/55iERhR+KUi3AaNmgm4U4cv64mnrG/avSfkL3iKu8sKzzfuTO
GwzAxYqcxtXuSvEIXplL/dJjVY3pOgtJMBA4G/ktdKaVeweUKEaGdSm3cjVkpZ9j
IlsUxfyeITy57x/MLB4PXu+BRDjZfufAHaeCE7wMT7+KflyVHTIhl2xYvXqwhRR/
TAQYOAIAFuOLk8XQcTGb4IvL6n3wfqEEohc3wxlR43FxweqQN/ybopo1FJwj3LJT
U9qNHrHbSfb6XVPZgMbfRh7hvBvzR0bpRHxVbyttTSfVlynCK4VD2Yr3gMUt+V1h
okDLb6MclK1xxiGWbxttPJj1dCa+E6dR7CaNeB1TA3BHs5R7C/BTWzZ3MMkGUTUc
zhXExkftzKi7ESSTx2FR8+5b9tUMWCYcQvGODlOdX3S6D2MFNL9q/oCDISUbYtaN
V3mtWSfpgsQAQXMrkTgrUYCFPYm/M+0WRN5S8qm5J8RYgMAbLwQXTYZccdWL6/0F
BdvbTib+p/OyHN8ZGsLEtrurmwrQRlVfqZX2b07LEGzUpteqN5jlm3Jz5/I+YfxX
4MWezgloLKMIjIfJfxi24eAwUhV0XxTZgu2sMOneo44I0mUjP4fY0biYB2vF9lRZ
mSuI02kGmTWzkFJX9zSXmHsFNRd+lF8KbfRq4pv4iwbks+0imQR81N1b8IEb2PTN
qpkH94VbvPIOADfl7/7MtEOmCqkOA79W9wrXjLz1xWWMQY+xgIF8M7FIr5JjkQN6
2I4/979lD9Obur6P6p5Ybif3zw+ufC/kXoSkF0umoUg4faOSc4ltW3zQl8rrfnXV
NjlNpHnF2aqVmgaZK55oujmycsmdDcPxig15ajfA2nPvkvN7mByIBrCJrtxMPKbt
lOkL+4BdsesZWoHGkBmRGMQ5KuqnZnaPwkzgHvVwu6BJmdvNuyjhTzl++3RY/FB/
JpG6YVJjP/fY1g5xSwqcIYWW4r2XyakQUZJRoCbFaOlocXBSE0K+l5I5D3OwMdpK
VopG/J1Z/pVR2Uz9iSWr9TwTg47raOCHMo1dYGm7ZDphzAhi2W2g/EVjfc8PZLJ9
ScSUtYRI2l4wHo/gra3Rs0hGPNiGXJtqOQ+GifPv0r/WmWipoazkPhuaIkAmbCNk
bowhOURy7xXhlKEmmtXfNtKzu21nJW8O19cjVuvCEFswlQSZhaKQ/vkL+BcZNNba
+hdyU89gOxpQMqFYL4MkngLU13Y1x6W+ipAlDGlpl2EjB3IiTtqZy30/FmT6gZgu
xEPnRBfH+zHS1ATEnUpuREPet17OigOZcsCb4xg9yVEGxsqigRZfoSWozl7HRURV
wIvc5SEn428SjUdO/V+S/MJ/pIvFrFauOFKGjrlYt7dZz/IEgBXBe9Assd7G9yCb
qtBNToW0vOYyjNskf1HpFJDJleE1Q23JwAffnREwhtuP7x+EMt46p19CjTE6SYLK
GnGYXsaWXFHqag8gkdWRC+UYNQXNrKDLyavsPApbqWxTpzki2k6YXi2zSJTwh4E6
fNMstBGA8mE78yjBn3nw5luaQyuRKyQJVriqNY/siDgefxUD9At46zKslp9qwbze
jdeyVDrOjTeAo4IElXjxmZbJW81HH0m4n1WLOn1FT5z1GThMUTOtDBpocX+XZ4Ba
5vE4SQtFK1bsHI8wwfcKF3Mpm/ALpjRGTOvIirInoh6pfTmE1SdWOQlsG4rzH+FN
DoFjUgQznn3Bx33JfDOimpDSBZ9yzIx+1rIBb7asExByGqm3P2Ony1SdZ7WPNauK
uke2d9TAWJhjc9S8Psq1oWR0f5mchnpyZLZ9vuw9rB93QpuyzpD5tVy9VdRomarf
WlzeTwlvuDckoD3J8yJFJebifq2tkqJ7JPtIOmO4+aRzXk7iiPGlBQW02S6VA18E
W/hI9tRyb5sNrHAFnEoecOrAEKrz4HVMmnfAHqNMYyaiCfynsi+SEAeSj/dHRuwg
wEzXSxSOwhLbBQJJWe8TcMjspfEahnC71S/7jeO8kzTFDW/R71u55Xcr03qp4sOj
R8G6+0I2yx4j47g5YncraC3mcy4uQo4KxL2jiRyQBF+901nuEJ5Hp4Iub94L56kr
sij0rSCBkc/0eYl/wg/fwSN549KHTyU1NDcUjYP21ZziGt8xweFB73AERJpK91cm
GOP+bWl0tCGhhj1YkVXnxamFjzXOkEeXDBqEqMq1qT6VluRq6kAPWgHdCzX4Zo0K
bwL2TnZxQrNEBiTe9gEW9aLI9888Ru+8Kbx4H2CXTktCbVZ2JsrBaHj+rVVn5sWD
BJQslX+Vv5m+WVlXyJUFZIzBv5k4p/LHCua37f9eLCPrQC2CWjCUUUrySudoQKZw
5RqVJmoiYGzeCecnOBlZUc4cO3myUyKgajE9WKS6ZEqKyZuhQcbZ8u1wR770Fii4
9jULqoPbkvYx61/Wd2hgQA6rw3tRFdVov8odSNJxtLipPpV9UOd9QLMnS606F5/9
SRfOD0VijZFauTomA+6gczef5TumSzv2iS2Haym5x7uYcicBtXdAFl5q3Y8GIMUC
28d7I5ZqWUWWZtvgPOOb1GPqgpE3qZYB2zBJFD/sNgqpZu4gjkNHyJPRRshaIci+
CC+ojM8GXbM5mAQMx831Z33flXabOS/aL1V3wmbv+GpiEJye+64uLPbnmQzhD6D9
hVAM+BAUioi0D6eRWCzNIt7XIgRepgMOhduYwWv15LzSzjYjJAP0qRAFA+qoec3o
rp+jc7liSoW3tDCF4vCKG1tp6N9aeChxCVPRUh/3ocJrObPQa/cTDDXcN9yIKTHH
7fTtAejbAxU/JG8xASeZIAJ7BVQ4mYUBGPmbuuUb9NlIcJ59afXGB9U6qM/yPxw+
dhX6bhd0Tv7m+DakbRM9PRGok9wXGXT4g/S0QovR6FQBgx8ZDNrAjYEz1/8s1Eku
R0EBJ6IxpKsL3KsN5ehQa+2FPpnirpbqBH4jwwZozK6i/qhj+GNhz0wg7MTp+xWD
WPYavs9v8+iSEqWH03XsQs8jZ6wENWnai1lhtEoWyLRsiMIWGqsbP/FYG2V0kL82
VF+BWyjjFz1fKcp8v/PkzSxF5IF2//h0A95IpeqOvG08BGVBAt9BEJspCQce2SJ8
xtGBRRL69Hwz6pYWIkH1naS20aJncwRVnhQ1ilHnf9WKfbt5/oCOJA09M9Vz2ET+
N/IDUxvzC4RId6gmToc1upBzYK2YN8gQFcVr5S8GWbi5YEsIixsCHg8Lj0ltSnyL
qF5AVpzKR/A+Ecrnk81T5g6J9rosZuL++NlWo3tIMne1as7L/li0lXWFLK939Uy1
zxUo9fl1+gJJ00SweX0XKaA/kE4r5UsQPn3uW7Ei/XDWqc/4k/LgZ8CmroxeR9lj
B3cVKcuSJ/nTreBiry85zeVcqf8gJJgJgLSrTzSRbUYTVCBEwOYIYjIIAqTHTGEX
vjPRAVVN0dkZkH9dqEUyq+RymN1AfAgb1gSbtRfAnrtqsqsklRnfENfsGmqawaZz
aa1ceyJsB84XmF4atItbxrKMhWN1Hzc7ykHLwC3tC5mXI29TV0WCfgkezCvBjbIx
V0c4LOKh41EhhdSs0/TVweD4IZ7bsvqn2qvUNaUmAtijczrSvGVc5mcejbwSwP4o
phVQTdbXBpjCRqz0S0wxoVjZytl5+b+3Az3AgwojkvqjCvZ4VE+h+6sD/Xjf/KAF
y9pDqCEeiiGCBYQctIVr5AVJARPkzNadEDreK3z0um+12TukzUNlgCoRHRlOZEO7
xJENXbBQAs7YklvoaUmjFMxerAlz534fKAxIdEs9kuEfjCABq6HfNmiUfUi3OvN3
+RzZoCRKJ3gZetbxrQXQ4SsjnA7ueHNShsZBI8a1Vj/ceHko2FMb95s8RLWTXqP4
viVLe6US65aDBFTXyo3NXaqlEei2YdoomfRnCs33ARHwUNK8mM1YipRrU+HR4COr
hb25NaSmihYZyQ2D8yws9lk0HYXw/NFJLHEAUOKd9wQ2I+EH/Lo6NsO9c/EfPEq4
OadXQ8qo6+dFv9BJb+CVyYvmEaXC43CXJJj3U+6beAQnxoGJlfFKCo8WjUQ1av+1
YnqYAusrRoOwDE0aJOommetIvCnRJfxH3Oja80G4T+gFXUK9xq90Ef+UcO0+AJt8
w0hENmERKQXnN9PE12DqRsqVcn90zn2/rHhom6k6KFH9r9t06zKfI66QEArSZn2E
YSDn4esNidbkGS6SQuOJJw675hjWYRoElwDaVXeLcQwbpLUfXssHszwKX2JYttVG
GXTz+d2UUjxP09s6tsr6SF4THKK+Ys6/RD2PuHXSWBi9kpiqfeCV7ffkdd/8FPQV
x2nPZ85vKpuXvEB9c5lJ6uPFvHwI683utX9Y9sNo3kklwf5AflidNegsXn0S5EVF
WfHmK5HmSfYBqYsDHooLbVwxjubSI6TONIjEEp+chJKP2ct4E9bw+H2X0TRCHeUb
LLuYKWCoJl4t34xhkyuUiuj1BZ/sWAw5Mj5XT6klOodcbxjpspW8a8ZZjAicN1Mv
PiHz/v9ed5RFvEfqKfC37yqqwotvkC40goYbxiP+ZgTlT3yKUrJdVc7EYBxpiEJx
97ld8mDKPfV779bLPX7tc/b7cTb7XbZmAtUPTeiToSwDWaRG7wGZWrFJWzbkVqwU
zV4BKxwGZqDtH/NsVfsvU8Q2eUHbimg1WjVk111rrF5UpVEC/2hLFFsw1BmjNNNf
VNksAg3qG7a4Am+9MN17eenh7WfWxokAXyVrvFIx+qhhLKY3vZPo93kbuLI2kVSb
wM1gMDCRV7+rk3yqcyp1E3cVdYRD22UwXETiH7D3aKu0SsiNVdSwwBROtFGw3uwi
T50+GmjGVaSBGhI70BAZJvleNJRWlgRbJPHvZf0lVGYfu1otJ2m3xaGaqHfsoppN
YJYCnhh+0F0HjBl+jF/J1miih4FjaTO8cug15Vnja61MN8Cgb/KU1ev9yzAQW/dN
HHm6Up1yq8fjU553wbDGn27DDKMX2/kMLA2DQDpHxyZmEDb2XKgU8U9fVB9OVCGx
xUj+stD+sWG4xyolFtqerPsFkaRwxHKvzmGYbgl+q61Wu5nr70gsRE7AYtmOQjus
J8XYfgo1qSbH8+E5n8nggnY5UQPVRJYAZEyljWGI9riw70RsDwJkc8XZa4fMDRg6
c2zmEHKAcNmIR3qWSQiNBuWGjcIj85UWPBTEbs+e2BSItovODFSnlx3JpZ6TPQUm
3Bw+goldBJBIWc/CRmgerruzAcVDVnIX+8/UAAn5iTHQgttsdoWbflTYGvzX9Vld
zfcWE9awra+L9M6SuZHqh4oBgj/2LZfbBi1xWbkDK6HtHN0tRJMGSViEl44oc2mg
LoLYmcQLqs+CyhN9/PApk3mYuE+5KioUZDrpGH1+bpGy/P84H+jvi0QUrsPe3i/F
IZ+mgUnBYgWsY31zbLQ8jFGx5DgbG7K8U8RQYhfgg6QdKcaTZdqoucA7yogrhho6
bLjbBaYFT2oGsItQAGiWjfAqY0QXU5rpSBUg+JoD4KFGWYSpXCMwLr2YrlWFsLsZ
omaMuYbf5w4Bn/Oa2DhqfNWoJlHjiku07vrBhr6X3bLt9sBy80fcOJWS1mFuozcq
c60tm+HX2sfooigqEQHggQzb5m0i4xqsxpxqm/jxLjEDnExa3XXZ7fJMjSI35Bp5
vFQGbeaHp8U4V1Mn+CSUgA02FaRDs36hcZ2gNOtLE50vbCE+oyGVI/MPlem/llXz
YJLJkyY5wf2VFSQ9DgOCm9kZJ07GKmyJhPHRzOfnkbYKsBIKj12U32jQv4R3jXLa
EOsjo356R7TR5+kk9WFSlYTMkCOwkYa0FNHJGjNCMUF50RcB/9sxMvARzoWAPEP7
7QhrtcQmhKH6s8/uuZQWVYB1kyJSybRG0AsRvN3hJhD+FLnOhz+s6PTiQLeqv1qC
FWNaGYFIrBdvgTlxWJgEaXsx7KXxRmJIbS7rhoYnd2B8dwZ256C3ueVDCkpVOZje
kDv9VgyhIStLgKHWmnSqrS5oJ5bPC6x3TOIf5R2YDiE/0UQOnl/xRqmEV4LuncH2
y/C6a8weI1cfR4Qrr7P4kLWZwXjIJbKGaBs42tcuILz4UKsjzOhl8uslWWceMKqS
3r/F7zdGaWKWyqorFSEhIIv5x/nZ5+E6wNCyo9LiM1OP6Bk6rpo7KQPhRfGKpiw2
n6u1MhG6iZzjUElY5SsTBVfn78CM3KOSpCJ9mrzhTJzEyfR/3jZuDqmV74YlCgnx
r4NCPrRUr4rfvwfIWglAYpxOZ7I3ncgz7h+xVVnB0s6GfIfN1lerXjKugW28UcVS
cjkCNSWeIAJPvKJwFT1xEPhig9SbtT4o13wlz7eJaHVarAhGM2Q+KPAbUyMayzAc
NeC44mzD9A0VOTer5ohcU3RSyqq3bkT0YBv2ed2W+Y26ptsDsmp/TTMUAz3DIiVq
qUIqAbwVk9yZR2gIQa8v+sAWMPQSpEQ1peasXr7Rit2G1IV++2ZRoPGk7aTKxmkv
mLp6AdAo16s2cQO5DT5u6WTf3Rb9vzQTyqj+ap3UreoQQjmnCOQBE9Eyc2DWJ0g8
VnFxx98dtNGqjq6LBB9jQYqSc23e2nzgD05dkrYiTpIGwSFWqRNwY7s2yd46BTww
ROWmbogg+TFVEz25VK5r9oMsIsydAwJm5KGi006wud6Hs7iMb1lVKmR+vrWYWuSb
nvipNU4HJTm63QuzMOiqaw8JP0Cw/iiqG+F2AvV22hHNXUTh+oPY9GSfwimNVzrB
r0hVeSzyrFVKD3s9Gi7LY2H9+p8G+YukcVt4CU6n+rx88rvVzHnrBQHxjNYOC0+o
Yv6S7dtl/fyTOvzI05nBd0dclIYXHXy2hww43+qHKhtN+xKOhXZIhDiQ+1eIjGIC
r/V2P3sclSIVy6KqiHl8ZYAWbQdRKHsBPDYAQuhBi/Tbuf5U8M9dkBMjJs28ZPL9
NLKS+BKPrzl6mJKn+BGiglZDjpO0oEoB2tdv/ggT8FdJv7PwkmZsUOzwYe5bfKDK
7mbeUxktBAczCNvPmF4kUs7bltVT9C1/CmyemVyEPq6KAy1FGbNPYim4cZoCoqD3
zKUQF2dZpkOVnVtMQO27gJ1Ll6AreLAo0kMHmXsymmZlqvWzV/VT5M4FKZLRRO0e
umxnqMD7oHWfcou2tH9p1cyRCFcQl+G2tD791MEig23zR9sVMostKQuJp1BUwIaS
ZVVi2W+xj094DeHHd+vT/4EAD1xxQqT566DQnR++msIz3S9+lK5k6//JL1EW1s5J
VVjozS0u7MtV/8SGAVPvixxHr7tfCx8dezKPBR4gh/NOxbdrPsJs9LmGjrAMWkzN
kJBvclc6LbfzJ+L8+aSh1BOvOz0LJsqa/ayvuj1T5woj+yQ/sXF07EhShNlPSKm0
e5D31aVU299xV2gNgMRK9NFVZmZJM5sKBRH316f6tVsgm1YeNCU7sfOnFkWiKGsj
tAgifYMexhbK5a49hr1dInN+s5xAp1b5N0lV6ypKUvT4/stK/gA7Sp3vFQx9VTCt
4nfvafntNT6qiWDzTD87Eb7upi1hPe/xSgAOjfKzIT6tRa0UCHmjoGegC2Jtf5bS
hkiR8VzVz+XM0th0fFnxZKTzBObPH+1wEerHKaP+q0F0OuooA4oDcQgRIgYo7RKf
Mm+JghQz8yhKySwSLAUBJ3c8Hg+RQA0oUUy3bt0Zpk0WSPGlGkffKxQWzeZHrqZO
N3Vc4iBMO2aNth2s0Aw0KKjU4Dy/HfmTyzY+abSwkvZxUAVdcwh+4prhLf89I6bt
5iXcNZVa211SP3IWDrsjiQOvulQ93fg8Id5VsWtw0QCIqL48iHOhYtKpds06ejfE
UJhfE3hMSyaCoAaaBRadTXY6KiVyS7S2rNbBTJmZd7ezYBgQg7kKqZtuHPGw03ll
H6LvUgVNfcUb3rFf3FpeY8tAnF4gxSzxX0M55jt/GUen0AtRRFrhMWwnJw9+FBX8
KrQUMmTt1qvpk1EQJYk5JxgcVdTfx0mydhJVhBcBdSxRU+AGJLjaB63NYmQopbf0
V6XHfSERJMtuGqMZd+3uC792znkaaoBFbpR5JcBluQuosYRLgmZ+qsE+wRX7SIqn
C7UlqkoAeOzzyLkZfTBg6HTgH7Eo58USdqgzMPfy4kRMVK0OaOjNFbDr6uEPEWZS
eeSsSCMoiJjqkJxMu9cVyad6WDZ1LfURzDI2JRrnu58U8W3qXKSHGYsdwuQNodsY
18yVdAa6qMwTOV/Rtrr78Us3x/ecwaoLqrJVdNdRO/5CQV8bt1mAv0wLXbXIR9y0
bRCs9JLKnf1GRfonhVAX2zI+GwQWKPF5OWeA6OhRYfVZ/qh8YQg1lfduLbgtJL5S
v2oCtzjmWT5gSvZ0MvqM5iVMaE0P+AiPZdylDQqeZGc0VDmtZHdKzQOcn3w0YROa
NF26fXQvhkLOKb4E9vrWEMnk6sPceJXjD3N0GJE1+QTmJ8N8vUg1RYfYhGB/HcME
DiIAE97oul1xHw39bX6rMNBzAv3/WHX0PsX0tYD1EyCf/w2y7+vAcV7MOcDT072b
EfBF6Nnqxv0lIn5aVtflcUGS3OUM0ybjCXCojALCP57KaI39//UtxJfAh6wKNCxc
H4kHu1EqV0QN1Rpg1m/tgWTIDKBikONKLXoIfC/JT38Y1qeltJG/5geu1IfBudGO
VE7uZoz0C999fkdbCP0k8SgCdaB/OOwrLqJl7TwD1w92NsNRbPAHw18hGQxC9jPU
qXXfGB+eE0jnUy3O/d7CszDqg3q/kk3kG0L2AT2j4EiEi9XYRZcSBg13ZymHICac
JRsq5uUcdhaSNhM73dWnI0M5uYH/+xJtGTctm0957KR+EgdKAHOSI0Um7OZJo8sK
w5i818r/Pci2uDARz+Zp/zWbrbJa4Nbuu1cnIBbHt8MWoNDNb3gcjCm1xEmnNYfs
sAk3vqs3UbPjwRE0Kr9BJ32XSNNV4QosLwPg+rvLID4A8g7KTkeBTz1Z5k5TZV7J
5RcA32jACcMWQSVWLHmZ0Ua8Z1ENWSShCsnbwnU5bMt839V3/9rebofeOplNexSx
EOBn4qCX1frmL12ggVVe1zL9r0ax8KqYb+WA9ST2JnARxDrE1Y6UKCcgU4Rdwdzd
bV9vJ9x+9mC2ypWjpzeTGw8S6CAMKPTVXDvZkLWomM7jLtFYSAE3EnHrozwUoKeC
siHblza3vHFdomQYXGLfLCzPeFEHIEhA58WjM0mZzBXhqXMsqtGoYubtw7DHr2lN
EDmn8M0X+8vnFTDlfTtJYr2IwBayVsVVCm3jxQwlMX0Wbz/BKbXUyVvJRhx/Lgsi
MCX2H4o6Tq1LHJydk5AbHJYSl12XUMnuaA4SJ4/wTtO/CdksTHyLF4aQ4cSUp0rl
Xb6TlM912iYYmBwp0AXfgjEndmGxyJ3xk3wVO0bgNXauIY9cho2G8k+BCxQzHAfw
Im6C6ippfbujwUtjj5QlwG6R1n62F6c4OIb3uFYUNC1dqFuSyjcXpSYZ0J8rQibs
g+rGw6maOoXTU/FQHiWfHMuy7CTTFCAiJOTHf23U/9WmQJQX/bCPO994OospLP//
DsOftcuC1bS9Uzg3fe4iHqyB85fyV+TxmF1ni3ZenixKtKt8q1uti+vvzUZDEHEF
3VFpuL0EWYPDB53qTfD+1Oxd7+gO71+qXgduJBzSPuhAfCCh5rCmmQYrgGuVbNk/
htqpeziTDnw89jm/OY/MeL6yW8q+Uhr1fv4d7RRlA/3fAFH94FfMgalcZdcXsKL7
uSkxQrREfbLBW8Q8CXy+7FXj9iVUHE8O1lsQlL7TGdPFoP8gd4aTEZS+90W/t2Rr
QUiYtmnwUyIIvHhZ+5cDInmcZ9wHE04viQtu8WaKkvdZLOFYBfkpodeS/yPjFeyo
JDKC9nPHzbghIPV65Cjt7CVN8Uh9+1NhPqJF4Gns0qMmRoObhVTC5mlL2wCIU/fR
GUXeayXz0LHHhf33uf+Pi7v46MYGwux7zykdct2yyvFl8JsVX8ENCOGbqSmGljqK
g7H/NSl9YmRGq2YLuE1hagEfUP8d4Q0u4CSmkK3zIvNRi8mgQwdeAUrXlA4NabXb
zfkiAQ3ZpukafOb2+/W+gKyQ8Zv8+64LyfBlvmMiHRNtu9Ym0VUHfHLC8aQA+pdO
KATw+p9PEtLB5a+mImVGkc1YVoEUqCITEjErY2B1jjuzesWX8kXk9SriKER5/OwH
6o3wgOE0o/9/8etm5AgMpjgqO/ifaJILiosOC50UnfFB1zftA8QmWNaF0tBUFuyw
qww817whrxNdns8M902WEb78v8G+lm+Ir52SURol20zGo93ApYaPlaNCexe7mRwq
DHsMcruuRsERBwsA8lPWjtc5n/etUtJO9y4CRO8yDpqFYxhjqZUoZMen2ySni/Vt
cbHDfz3ZauYTN0Vx3TnIu9cCZU+ZLh1yKHZ3MGiRw1Ho5ckrirX73PMnG3yorlnW
rAeus06llQGAteGPJjF5oxlQCD/aEGzD64Sp7KFlYB5ELLN8LC7HhCLNytZkWCZ0
byr81qS6onMPHKey+ihjnYZZ1qQ+iJLwK1AkX1UGf7TtZw+fW0mgXOvyjsjAWXlw
mO8m8YrKoR9H8iNoF8d8RH/1jblFBU12fMOKX6g80RwdVbvvjgODwl+nPItlxTm9
RcqS7Mn5m7agGT3CTarcG7opQJqvsPtVoWlkXdoH6m80F0jCukdY9F4IBLoJoWBQ
D3KegIBJEguSahfmzgB3f1+oYpFofCCfe3G60ykyDU1AISPBLd8wcm4Venui4wNG
5hpRpVyicFvyxnbFkMgde9E/KqfYlblF0bTtlb1uGyxgxMapuPDO55Y/j3zEEEaH
fQW6mAVmcbPd9qK9W0sKxZGpwc384FPF9BT90E/6sb9/n4zSwscOPrItArvpAy9Y
zOsrS5E2ZyjJHAki+k6BEBvtg5YhK0L19mMa4UXzatIO7GS4nAakV+D4jX1hXIAJ
8WlsmMZ2xBmdxB0f5BMhZm+0AbbN/7kauS9U+PRxXC7fzW+eVnxZJynLk/1gcxV5
V7Gy7kenOkWZ5noclTba/VrZl70sKrkdEXkS1zmpS0VLFqP82qLa9GqNJXFTJ+jF
trbBzGAb59+YiAGf7vsthluIk2foA0IikjTG2vfBQwc+3PXJd97785PWuNkJd+4E
nMx4F8N22EljDyGsQyiahZ4ZWkdjiv/mtpRlAE3y0j3Eae80an3KEqGqq5loxvry
XrV2AC/IxiYkk60R+Hudo6UdU9ivhCml7OUwSyL86cOeBcnrMA4B2POl8OtEEVGG
EzEgzAfzXcBI93thxD7qAU3lV1JEsxmf9o4OAkUaEuyDgM30F79lHBKgvYu+gTk+
WVlqLqxRU+JD7Dv7nCB5sKwvVnODjMZB38B2m/o27jCq/B03fN/+/9/Ycx5AgY+b
+H29SwnW+Ib/t8Ww5pLrbBxdXgqGDW34acohAtT7RpwwFpareVntCwRBY/BDp21Z
v7+NuadvOqrbe82n7+ebdQ6TmPEcoz5vp1c7ddRb8rdN1Q76/qhVQHspyE1Q7gZJ
rCmMDcT4ixCOlaYSk3o8fxYOohwqt9QHF/rn/cA1Pf71IhjkjZ87DDbSsJNIPB6+
JpqOVmPPuOzbPT2sVCf4iw2KfPXqJBwK5Ka9UyqU9e+Nglc526ee0MMzQBl50e90
MK3972Mmz40CkHPU14ZGRWzcRCkt7ln8ZqbhHInOdOBdRDNTPle2aO60DsjNISF9
PS18tn7VX+kjPOUZXVglsBOfxp2bhuRQ+HY9pLvRW5Mpf0gp/7Qund6n0w8nYm1a
gUTouOgid1teaCxY7K1w/HNxMB7/izI7Uq/fFB7VVvIGpwlsZc4g9NRMDXcu23KH
KK3RpER7z3cUlvsLxsw1V9T0kzFzuN0wmstibtW5QOy34zb7Ub/bKo844WaW4W82
hc3Wh0PcUn7MewHOOcdWqnUXbc8Q9v6m3N3EN+vDfmlQJ2U7mlSnXD/4M7L57UVf
LMEUbdT6khl2l8KplWA4hYsIrrjDT5D3socgJS9Af0b6OI8G907FMu9EcP2b4ABr
RExdZFwQb2n84NWktZaL+tJgfSWjLnb8650w2aNzeiny5/WKCqQloJL7CpUzjqbe
tPQARuyV/s/PHL4zyXpCnodKjPHP5eDVzhgpBP9EF7PCWm0cHfXTsdXTx0x7jq2r
ozHkWC0zLRx+B6B6duqa7DIdJFKUIRC8iylOSeKT50t9ZHa46cJU/cZ4QJ81t3oi
P7IpM5reJeKiWr0m6D9+Z5ECyAUyoq75KAtvAib4RT5LcVZwym4lv80gsTIP8GsY
CsC9lWRFLMbGCuJQMv6PCJTBlC5M7Cq2HmEPqGmzbF5ElFC/JrizEEZd1DodL8ao
7NJDk+WF1XsRrfZAfaoJIv/lNkIx5ToyXNLQ6AEBDhY3zjWgsY/Za1yEZ1oNuPcp
VOot4i4JD/mNgcKiwRvOt0DlsQrHYsy2I/Oywdc3IEBoe9mqF3IznfbrV933jIUF
ZoGATl0iSoNPaC+55Gx5Y6F6ZKw4gkBvHW16GVGj8IkSEpf87SP8udgo6rmiR+MY
mCKpTq/sXQFSDrqXBn856AA9MsrV+3Xlz5X1l6JELAgv7VmMab2qT2Tqo/y+lnFE
YQncNfk9gH7bx6cqfjPFqYsAM56wucR9096th7EBA9rQL6PrVoOI2cHM9vlp7qZY
zINIjqOV39GLTuAcS+B6DrneXyIZBrt3ZrWM7BqpYiq4NRktZzRh/bHaaot8b3Vz
Je8eNzguI6E+2CvMwGKPzGDySOpd2ju+kUg+cpRjlm9GVgU+o2QDAcTNFaicw/Ob
zFHUM+4NWCABA5DJX2L0Svu/Dorq61/gp5LH+PNES0PDUpFhM24mkjKQx+Voj+xI
oxHCxuTabnADVNod9vKp7E9p73fg6jLQEw+QrAhSaaiqdbvf8ouwtNlS2KtNU2AE
CzaLUqQvt9ekLJ9VGCC1iEMszMqb9uBI074+g4uy2orjgzBYAE8P4yx1ouihvwS7
AM8ikg3vQuVBmbLGPQM6FNg+2QIU1vKJr0bnQHfOYd2sGmiB1hgJgOTwIdodejLO
P1zorCp8kEsGrbiPD0CafjGgUa/F7lM6HDRrsTiCurwhPmAc9kFRmnW6vIDD6Rlg
gym1wdrBpWSXo53jY5q05Kd4PCcuej31THd3IWqEcKVohM2FExlNE1oMwDg/eGzt
e7N7QdfmFXIeVJ+uWIrRdFghIBKI0XjOBbJHOZ/qeLzjva8123J97Y0+eUXJzcXX
GteITpzA7xIKz6e1DtG2qssJVowWixfYuPnsiy+/PzXUe6kYti1otrDCuI/BL6KY
hLxfGEhN79pZK8BwdXtd3ixLShw6XZZ+J5lohdI8AUPRugvuLzynfz+zA1gcvlS6
JZryJPRANBTMDosicNOAyqj5MT7aTtQZkgHc2n0cVqfDDdGpR8ZvuhrpvNTWkhU6
of+3hX+0Ikug4g+Rjtne2Deb1OrACWh1ekx1Q8u1szf+ax674ASG3RvjnhUOzbMT
OIJDB5hbtjeeGSLjy0NUYcYf+xXyQsB3Hf3X4Bbi4/RQMnEp6Ipe8okqPIiU2iGN
P6DxAXMHuuNQZDzO3Pf+pctOflHsCIRo9Xahtu8E/HFPEFjyNjNcRR3kTD7EiOVS
Ihd+J0SMFmIwZpX/j9KGwxISNNv0soaiKVaNZbhLrNG5b+x7ynBA7/mw5tDqYSro
hXoi8PVyuWyRLfW5ZMXR7LnU/OO/oG6XQFwvgyctXGfDxiDBmmWVZBO4p19o1jHl
HCAdCXZAUI23J3u6SvMoYmI6PVYD7YgtmJy1prH1kTTq0CQH6IHLX9cq/6wUwtdi
YyOr6zcs7on7fx66QkFQ5DC/F6RYDcg0qPADEG7YfmiCfas2MjUmLVlMGOwU5f9q
HxoXNaJpXod9/aQTIBNEFBaWe9AVdFyMhyYd67TC9fG9cweKAyI55x6jMf1U1bdK
S7QSWYgtsrw1IaDIdoI95930CZzMWtVik3OuTlOn6MZohHSiUs6uB6a2wjR8DIuw
/+8HTJnqiKjpsKdvvkVGQXtov+0OsjDZhjWA+N3JOgaEXBbO0FUW/3qelPBhJNuj
JbSY2tL9pD0k889UYG7az+VcU9L/EHztuEGdV77AOih+8BsAMhOjybbAZW4626e2
sd9zCFDwR6l3BK5GXNZHkfa3QBPna8LDeWKeKl2gBkPz3ypxzmfI8Pa9OUcZ8V0T
88SLBPHgG2doJ1jKxccudKT9sHMtT6rV0oKii0uy6G/2qo78ZtamvcAX7TZfS/i3
ORiJZhiRcwnJQwZqLpuLVgWdZL8AuE407uAvMk94GyaDkCZ53cfhjbFId/kOcinS
qURvNzfQHqG3NRAtbgSqVZeL6fChSrkXeY7rD/sAQgF4aQfKC+Nsyv/y7mlRiRwK
Odw9gn4ksCJCfipSsdYtZ8K2GcxumBApC5Ctxk4i44eahpEpQGFXdZa6hVOPlDRO
u1w/A/Rs78T17zBcnp//boHQovA32sjm7n/7NMbX1W2jsqCIKn134EF4+whFEqin
G3wBa/JI/T9gd9qC+8t/+h9ddT84DGRbe4XijSUrzYBMk1RsSwHCIFHf+6si7Sqa
HvxJ5evz/bCpASSakEglgCwSzFBTaqozpvIQDgcTEhPF0Q3WtsvnN35SgpK5RSFB
Z+JBntie90Y6LPX4yw8x9t7RRwaAKAhD+qme+Blh+eMpJrH+Glm9DH71/wIQ+Tka
ot9nkbKa9sO03BYLpRWBN18nMbpimF+ijcvA7giu3fUsY5q+ZE81nPEQrxP2ubwZ
qHgzVyjIQGXDd7LB8x9f+uiXIUWcGNqHugueS2+gQZuw+BAQfwiRODfD9ClFKlhv
Jg1W+RVKB31WNXRbXJPwOv9zWpwQB7jaeAmVuiJfwOqEAAF4xhBPr+2OOL0MGliJ
o8v1sGP8KxAs2OHfj9FjgFfalPnn1Zmzc80FNeCsz8CJJ/8WyaBs9b4zjEQ9jTID
pAQCzbysojxoWJg69rj8aQwrNVshdKTKNKcwEBf9B1+r6vyH9n5LzGHEj7xB0LQI
S4Gh7/jA1c+oXzoeQeisdeDSZwWbu6m5ps01wecejmaGFsPusw/SMnYu6UbIJR74
jU0aYvycnSgy0UzTIHCxOEU8NPj70i1BaT4VLRXxpWSZeAYfeZb6Q/KkrUNnMQ1D
1mzVdpEikCfqoKBqtbeR58sXkNj1G6tjuAsop6BNy1lhrqHOfI4nyLQZYUSOT8Wi
d2YeqlnRCkZ8l5YnUs5RDM/003IOS8KjJou6uqev/dyE3HPstE/wNqV0ACVbkXIa
nIz3Y7ayICKiitQAXaevJfOUUG/goVDeu0bCY2d0zvr2z5FEUoYDpzEKFmW9Ga0r
hlNl6J9vYNPtFBLHzoy+6a5Xwswda5/u1fz+ABeecWzrcYiHVlaMUt+qMcjh3gX/
sn5Xk3re5hBlQ5a7ye3WOzY4q9yy7ETr0BmsaJLBHXbQvDF8nXLTJCzOsQTz50c9
+W4OmM0lVdyn1IEzLLu5RPDfT6gQURuSwtBPP8kwskiw3mXcSazp6EYWgbikKu5a
dwKxJV+se8P3Cz5ffd/Xv2n2P8iWtLAKNNN0YDiHYG1kZoHYy8inE6SlpQx0NM6X
fbroRbtTiz0IAUWolEI/BWbJkeN7QiZnaH9rRC0eYjWgbNKh+hMde5qDIyrQopb/
Cu6Fgre/VOhxeQZypL2CYc3i25jWCLJ1Y874QuEkypNvqwTbxLB5xQzBq0b2W37i
pSMXFoFmpdoFvd25yDES6Ww8Yu+sNXZA/1elOIoRbhfJ9Ki5RoJYLTluEJb9H1Y5
Aybm/38RSuLs4vx/ZphEfOv8LLJtU9MNyxgB8yXz3lhe6M11Bq07BdkC414AZyjJ
EDZaqLn9G/TvBK29CBJUpen3U/bIHrdZIds5fuftG/B1rs7juO/ZbuAdrwqQxAVY
SVEmxZUx6uXMOPJQ6J5egScFjN+IshnKbQZeJyAIsOtFGHfkiiVvARp80VcppdnQ
hA+VpU7JLfdMMsGFMWBPP3I1eub/4vRpAtRuMZxo+BzbA0NpCHD46RYNWAvGxxDl
nvf8dDi0es77OdQlW/RYHpTOgwv1Psvfs+uJ/CXCi1sJrmz3TEFnRFGu0KUl4czp
93Qqyp0941jAj4oMK0Yf/KrqcWPl+cJR9rJiUjjEpeoFDTsTcMAvWXjHn3xL62pj
Ugfp2D6KgsyuPUmEUcJOXeyKtz2MUtFZsq/CgRNwYueCze+xH8WZvToZ//uKPnps
vq1CLr+0s/8E6/ypm28T0xpBUJiMFAS46m1Pu4bGj6xZa5isTzUCNxBxyahcQWNu
N8hywHEKCiPVIQ7FxJFkbqRjk/EWaNIsDl1RBGocl1Ba0XMOhQ7sZaztfqe67OJ2
d+aqoeICsUmdVgHPEajaWd4oduy8CLopJJMk+RtMUaKSu96TbDc9eFi/mmt9C0jO
YMLySzE93wKuG3zPkzqgmoVEFYI3dV9s5DqOYVM9KC1ev79iyKiBSEVYJfXckuSQ
rZ8T30b7xel9bcUZsYQmUoX3RRkl4fEBBLO4xrRhhTx0Ys5FSsMETUfkrPZrDB32
jw/hbUMN5kzkZTGljtuqD62OyYA/hoKPIYoAkF7gcuqb8aUp2oDujh3uGFQ1oONF
+pUzjJCudtVCEZ8qmTok5XrXWAjZCFDbC5LaFRsbkaBOJ5zynD6bMuSHCOuWW5k1
2dtDyhHSV9eQCz8Rr30UHI37wYY8J9CI1exKFa+fdPlBtzunfg0FEUNIyX4TT7Nv
eCdOpVZGdZYVd78owf2IIRhKSGyRGIa261qXCprfV8LKkCLrUgB27/b3D+8qR//0
LowlxosPB5KTBuDVyM12bJw/QbjjpjG8D80RvtOGSX9Eq5J9YeIUibPH3DXAJ1e3
m4/2bNLy3IUtf8oNF0CcheFhoXW9KRIY8iGKbE35ztL3Z+0NQ7lNuPureYyd1IB8
eFRxzwjsAULFRf1B5RAylGUUjMxrcUU15jZN0T8jsrZ1Y0QzvqEsSlXhJrwSDEYv
DH4AZUeuA/cc3NOtN5LiNwwrGePCQPwbG7vhYDbPZVGhsED0iqIUYy65tsmdciT9
urJRbSmd59VBgqvLVx1/70dOPgCM8YtGksH2DkzooV4yaRYQOumpgTGlZ4RtUL0N
lQMeUYT3n06dDN/5as0it6IagJ47hV5H39UkzERUx6tT4WwxiTga4SFxx+Fv4E3w
sgBnW1lHdLFzlnRjcCJpdKsO4uZ1SGrG58QIzn1NkoiAzDPUGHGgec3XBjFE80GQ
EQqC2GMs0QbIYGb87NepZ/oi2LL9pGcuXxxdHWuBmA6KQOJnzzbhde2saB5xg77e
CT2+CEazEyZw/dj2fC9DB7VYOWn7S5R2EBitZmMQlujgRvMIw0Y9oRcKbv2VzuZc
sY+2BiZubfUBJPDV2gPV94EmoJn8j1CZQjnqt28SGAphzfrlGRngKLLpuvdJoRDN
RPT7kyk1ttT1jCg9rEYmCvrXMrXQdMPvh+tzWoBksCMikYSgsAKgcjVrbp+j7fFg
BFSR1RnCZuFZ9IhAZxqz63ca5HOYUwS1gZgcEuj5bhtwX38VOyfc1XddyVF288pw
6NLEyES2rSytQYq209m/XqCRs7C5vXkDgfTbf2cXSXWm3qBpspGntWd2EpS2+0jI
yMpqYakTTprWnvIW4gJq6fQWwoGL3Lw4MagckP4eKI4r3DlRzt9AXkoAPJcZDClo
GCqU9weE+Uubx7d9BV+Yvj6ndJ6LQyq95bn9TyFwc5/U+CliHSjLSOOHCzyQgXaB
2mVPREwLC6PDhWpeOWATfyfW588frvoH3G5Tk8bJotSENt6Y6SKiT2PWryHTAXCq
gVnfp8bftXmxKo9NUWgQKHHod/L74CfxxpDOWYwVBTvBrPc1i6zNtfKrtaxoqCIL
m0M2CnsSA7fwjsdGQqQK82kQmLSBV7NB7HcWEr4xYHvP0aLt68AXHdSdeYu6iv0u
I4T1xUYMpkJ7b7APKFnM4fKSebPvJQtsA25cw4TNEkd+prOFR3KC6VRlFVUFaQrf
n/YBbbxKOYA3BeV/fdMoL/7BLNVmPlW48Ea9sD9D5aUdI+1wyAY3c+wClOfUofEf
LERcw7fBi1FckoYkKuPyRReWfvU1nPlkSfQVuqmC0ZUxnEjrzl+bPfn/f/9RDQ3t
POXkSHXC/sl6umWK1dzuaHyWM5vmfeyLL6W+7GcCIfmcHZYf9hvm9BiTTJH7FAi6
RkX0shIy6Pd+hKVbO4foObxahOgktZr8oYO7CsuUYHZxqMvnVrOArS3/uY6YTuMd
bo2hqpatCpUzqukh4VkGv/Vt3bc1szrNQ9CAvOX1wL/O1BXYTY1mzDJeJSOEI79c
B849hgcCcfR2XUaMSd+A947hl87ANJf8mPhwqAbxIBkqA/x4IY9Fj8z8Y2Oz+RgC
FTSjVCk3OVbnkrn+777po+fPY7df3XcGURBd7poQPDMQ7tCslGBIlSn96tMfedIN
8PMNiGoSAJ0Kbi71r9eGbE1OWZpsisYQ3JR1KDtG1HcPws1F5mfTIMcG6g4Aoyqg
Q6Tv3D2drTPRh+zqOumL679AlRoWY/C1CtfChOi12YBQL2ijvb7aRa8Lwzbx/e9/
47xd6wfG/WTEZS8bnhPZ4gbJhbkmjUHJ+N/QPHpqDdILx00vQjveFSsMpCOxCG2+
IS/qJR3J8GHulLCOhe693esZX7EMzRyfuW1QO3YUPti5YetPK7Z4JLCwawuhNdVH
mM+q1eEg9LE5zPsOCtc5uorThMTNi45AVLnxjKyJApoNkH4235egvIg83czeQVeA
FnT0oR2T6pv6oNKaIJ91KNpPxw/FE6jDGCqDs7Xya2ZoRdYaBinDSMQuppdMZlsg
ewKA4iDfGSAbvKo6FxCtTjsYy8bqE5oI2ewZ4n3tjUcwQJNUKZVSQtWAUG917bKu
A2mbc/o/CK9RE36i5tpJt8FwDnk7QBTM4ZVnj1v7ljgzpoxZ5AYKgGcycyNkkUas
ozlamGYnNi8kqaAob7dhfZ1nJ/aND8vgcxbxzKcPChSBgyxjIHCwFs7grAOY4dwp
EGG7bYOeZhZjm+aY0ute4gN0F9wsqxzvn2IYmo9KaWWR0ybl20hIBJKhlVM3qGkj
Ym+mqkHoe2BL6KwzuEIIECFqnpBdWEwOgHWyetJoo22RsQw2kqoXawZI5f1lz3yS
t4aRQmHlTXAXDj/T/Ojof3RCYw4AzVKQe5/O8oSICzFiUhjK8vw93ByNqPpQZQVT
KtUm0xBbUID1cheC/uHblFJQWAe9WLui4EYQ40yhlOqFG3Ck+gcxMteThCOaG2Gu
aryVk2f8PpbasT7hStNVeMDjOO/dIAzglu1euH52y1Y73uJuA0eEpjdXSHCH3l1F
R78I4wDPNkL8O3rFJ6Ru6coKGP4YpLgWd5V1V6n2SavxgSDxdmooz5KCWQvRZ9vv
pTVT32hp/J8Ug0vnGpsBjkszItwPfCLWCdw4vElqz9upMthzrHdSp4IkbBH2pTmE
qWZPKsXFN+t86ChXjma/14vtb6TiPVNk21BGKEiaBMQdPYsMm+uT3fnHbFZlSJ9s
JKdJVHol3DjKGbAV+/jEnbu+p6OXqaaSHX+x01aeDe0A35D9zZCNQALL1fNAeds0
tKt8CWNx2GQyqOJ04P0H4/NNjwkZGkz2exRqFzrU+XE2zCgow7BF0Ag4gWxngmUU
Z1MDcxriHQwLxn+gIW0k2u1oiO1t2og9y4wHA7j5IGdJ23k8wIvnaPtmz6l/vGz9
NHLZHnCaqrQd701gCNUfvRq/6HJTexqYMNX9PFkZfnq8qMwZVHtHRZnpxgRFoUFz
k7MZFqjiKwdCVTGZHGsRdCW0qs7+doLzEggnke96FjdopwbS+nBSu8vHfMpUh8Pe
11Fppb1HK6xz/mqfr4x1YeZzzhl1Q9ic6ZU8NEjQCjn+viydY4NzKDz6Ga4BDiUN
UEZfUqODakhVWpMpAzpvSukGhfTtFkVaAtDXLmNxPcPwnWwRBe3MgyZC3lHhWYWT
PddTQfk7/ab51TTB9hme1KIzY+p1b9G7o9Sd8UR3ADJeQ+5rWzacvfuZQfoFBASD
uNnIUH9KkKEj9oJdo7affMDmJ0CFKwGM9B0Cc3JuDfKGQaRBusy++Uj1JbZCh/1r
FbDJk5z+k+9n8pDmhg7mZ2C8dt8glBbzBJ2kOOK5tNmfoPaDd1pJcB8BAzcqKYBl
xsWGJdMQd+h82uAIZs7Wwjws4//l6fiVc1J/jvPezBT3ozj6PlR67usWBsZKxmCM
pbFOUgws4ce7/qFuTFHXXYJLh/WVVxvOeuor+Z0HgOeAa3OHhiUBOV2gFNm/QD17
5kLQ9loQdbVNxjGD23c37c0uRXQtUJWYfa/4cUqvJZIjTbm1PtGcVElPlvFGTxU9
zvqVotrf38EurRn0bpC6u4nWANiR3r2rYous0sk00TiRDyO1rGsiSnYybuVOJzP8
2Bs6604OVZ5ixPcVIm0F0c74V2ugkl199hI1N2IlHuzTOzykeGM1izAWZ5jO9WFf
PJNgLTP9eiIrmoeSu/RDBGPDztXMIY4/WuMlpGeuOhkPK3YQYMj9U37qon+VHv5f
i7QzC2muIIE+E1SyeTvVqMYzQHzgAyAgCfZNUgRt7LGP3arqHxjtwRpMtXL43/ox
DPLvr4T2sNJSI9QbH08G7hU8SLjLkx4LOl+G2SKTr8b8gQKeB1L8MAWke5Yl1CuC
aE5GNy8MQe9sbVcao3nuqx0NVtpWfLiKt3TvBISuCOCpuLlbeFLmd25XMzL357vv
pQPCv7ZttV0sozJcKAR2ukRjF3N9uMDm2YFfciYYe/FAHCr1QK1GHiPq3j4SewOM
mgWMvmXcq1zQR12Ku0d1g31hv7XLT1NBujRvteUqW41L/yN7y1lxCbtW08CV3bNS
0nOgP8A7CP2P7/355dcZIVriMM/LLVmAvERFBoO0whh/AFhJe5mcWOcRd/aF3t0E
nnBermHSVNOTcZP7raTGoGoFFtW9oOzPcxDgY47fzSjMNGm0aDYiITHrxQd8NJX/
tORjSgT5vR7WMF7nHW/8uut95YFMv1wA1A+OB8uCnrpDiGLGelbZkvtHGBtsjryF
ZHFaCAnz9Z2r467WdBz4zlpZRD48VRc6rOgTQMymEC+Zr6UOZ1wHXdQDxy88nX5m
zy8OCi0SqzuBo6hyxOeJIEEPpV0R4Af1RpmUvBNoYYd9Q/bEhT0KbtEmA+jXhqwg
LfU/EemmJBZebnTPoP9J8+86HE0EVqd7V1rHwNGWu0qD1d2exJPsAtAZQGoKFBta
FCyetrwE1n3OAI4N06YgAeyP4eEXj/iIzYzzqZ+g3juo6KaH47kZMh3DHZrK7YXa
c3oiHrybclMnKZTuUzLOpVxPJl4w8ZueNLDedpff4y2QRwUaWu09QnVihHFw6PzZ
6L4SjUsLgBKlIyw6heM1/7sR/WGEVvdlEA96NecqCGHKEUtuFDDz3bFEI5FG3/33
AqbU7NDsituja7vpbLmRUgqwOZL0MhgfTqgqblBb60tBbShBT9DHQkMrlRv4ox5i
FcWJMgc2ih+VshNYXM7urRJOk2VOrknZq+x69/SRSomEstAgegY1G1YA6xqjKtfQ
XK26GxjFy5drdfBLMX1zJttMYO4aSC5YWi78Lvk5Qzvgc+g26rpjFigDedFHZdD9
FUVJSkKU5Icq8uj/wM0CisVAMyPXyFrUofWedIKq59k5ttdKLPzzGQpecZNlBCnU
IsjlrXxFQkqJRmegWNQ77Cdra0cK6I+19jXkWB5YZuJZXyAexpMvfoXns4aLs4ls
QBHOctjK+Fx80AwHmRB2tr5PjMHa/RpMbAFN51mH7iKb6Lxa506bBweVw7Fo7uuz
4D1JjtMsAgv4mU9rOpl3Dz6747CSBG16tT/kbRokdUgSOIzF4BxouDwyUSYTBI5T
0LTzQTPz3RcD7VEz0jDLfIQFbSuDbpev0qsOBo5c8HHEyHXbEBvGv+CVcumuaG7/
cE9oRWctIZELkwhehCTplqFhm95Wx2uIpEUhM0wpEmUkhW1T4ozh1UyuYWFCWnT1
OguZhMIVFSEyBXjCcl+GVAnYCP1UjSiYPNVV64XTJYTpaLgXxroUmOFwmSTyUOMh
YYcMOIwrPjTbZuY4U4FnEMoyq3CRYY629NnaDUlLwRlNXnFXDzn/Ic1ofQ4oz4bm
vve8JTCzEaySYM4GqES2tGFShbMm60UKJxzUnw1n4rdVmyqNhHDS51FrPINPaGUM
J8/Nk1km2u/z9Ih9x8IVNGdt5AqNnZyKf52F+LOFhI577pvKgB5ep+TQwJTduDtB
CdaDH1ygdwweY5RQsHUBl/akAMakfU87Fc2PIKlNCRvsir9HmLrn1NmHNAAO7ncs
98zILat/XGJkApKBKLcVMIcfAtwk1BbRfBY9H8hETE2lTOaYXl3kd/Fky0ROXJCA
wP75Cw+hgBePQTqJkPgmlrElxHAqNEMlzE1aVItJAFOkkEVnwn1Hz+7VRq1x5n81
bk0sAJ+Hk1ovgoBKIZfIYdyt/LLrLFkXgJEkYLARpXjXvtffO9CC5te0fe2RRiUm
Zc/E5a+ELHa+YCwpiz8YPb2PdLTCeOTciQOMw9Ynp4pG0Fd8etKe7Peuj22G1Xto
S4AhAUfJdDgVlZ3+40c5dfD1mtxlf7xERXkxchqn98vKtGJVWfIG8a6uOImhB6pU
26u/5NTbUQs7MFSWkUbqDcXtQToNGn8TAfaDjEhIDZypcZLABmfGO1Ld36ZlPASM
KCB1RChpUR5Xgt4XnZVuA5mSXzL86Pp+PRmgAAl4ZBcSUZu7EE7dCmcHPT4EVDiX
tKF51k5FkMV5q90S7lIrGcMjb42lzW7FLTSZ/o377neRkyTzgwADml+6CnRJ+yTx
psFKLVcuhpNrRu6K1nPy2V6FJvl1eONxzRKPFVjfodHcJZhMCBbtciEUAsLtdsyh
UazPnX8u2JHukV0MDtHH1W1m5UcuCqwS7PADR5px7k/+ERu3P3wfsKFj9t5Wc3Sj
BXQ+WlzbJIQWVmCXGeVmAARMwSGNEN0thY4lpZn5IfHrS4rrmX3TMAENAoI26uee
W6DcG14glhNnFwaxx7K88hJSvPdjIj8x+3YTRUbqlapg9YCVJd1tbNw255o2FHpW
hY6Qc0Q3aeeoO290vdtM5WCtorey5esdf3/XupGCgVJ6WA8vXak41XxkRjqjwtcT
R84UrG7EptEKkz9mw+kF8dv0VyaSIDv/kEQPs7zv8vrRQAgV76ak0FETIgbYfU5s
StmVaMfpPCfFzGNs/x3EqeQ8b1Z6rXicTiP6Pwzdhl7GTolsyAWpNP43ffU+emjg
0C0iLBAPgxfq2j1e26egOq4F+NOWZ+pLGrUaabonIrPcAZDbNtFm2gsQZHcoUG+M
nI+19EYgrhg2ZFSW4t/N/03BCWl/caB2tHbkN1l0NAXlK9p98PJCInIYSblsaso0
ztZGr4rSHV4Jdnu2qwrGfHvnlEDvBGowitFiT5VjCt9Zr1zm3qUv0w0HSpPrYgVz
3yafkyP7u4waxRjYBEeOB10x9emCkQ8cmdhx6zb2k00VIr5VbQ8OPeETyVjw6HKy
rPl7dZpKZidPHmMTGhSgd6wOBH18PRM1gNZUxdjNo+GA+JFHmnNDqpenchwzy9cQ
Huq/4HCgf89T/TER2//zmjjFy1/CCCGOesm5YKdsTBFwL1SpxctRJK5bK+9qMXyP
wzFp8GHDoLpjbTmtu6u7RlZGZVRaG3ts6dEeYKZF8YlpbqmX/DB42Trl/kIlW+tA
s1jByh2MFHQDqqrMNOy8nkXeVhn8b9C7DXwFGE3nakK2qd5WISK5U8yUtBEKIpvd
b1PlbAsYTf6+PDA71du9Wnb+TM3BCN/am9BphGtWNYld4XKtg9fCnKupV7oqayIP
8se+pguF0ahD7NX/zbX3S5RaRNKM5QmJpOrrpiN/UP7OrlxHqFjqaCF4zt7ceMtL
1z20eOCkJ2wf7k5TDKM6WVmKi12Sc1VO23vFWBiphBuDqTpf3QLIVAwc3+qorwaM
3JK5v8dUQwVeise9c9IOhCOi16bX4dC/KwYHzp+M5X7M+9JFcP1OQVp+/Z4DprOU
7HHoy5vw42QeyiE/D2aN1fNROata7NrR/afv6M3dyZ16+90QoxhimXQNu90QDleu
iYva+iz9DHmP1Twiqg2zaLD2QfOFMTQjzMMqVx4Gi80+W+8zzjnbJXbDc1r49Osp
MdWdJzBirxT9Ec+xouynYGEWHrf8DGrgw3ejm94TtK4H/gmP5NN5X55/w+rT/8ij
KIpJamDqFbljszMYVPNU1gQHPovb2UFWtrsiHd9QGwzNfLJJGQkyk1ldbbYtJJhF
u1plElYU7XpwHuAfUwWETcEwDAkozadMv3a/viFOs8+PnlqGqrlrLQs25Bl1XigG
vfvBeap9xCuO1Rw0O6mCqOC/fOHNWlwWdu7ncrR0nRPyKD1nxNREf5+Hm8z9ZmNu
D5Gkps77rrFnw8p9hNttsoixH7qifPjaqY2gHpj2vx5L6KORpbptag3Xt64Y+RNL
4L34zuwBagoAsEedfQhU0at2Gp/OG5+9sVjoShnfNvTYZMgszBWlhjRS0Toz6lzp
/w3ORXZJ46mOSz3Zyza8eUs9x84Gvf3+RLMaFkTZd4gJBNrEdM7FcqRkDEc1wV3T
RG3/86oEtjXzDJCJWWFyZ3n0ihoRWtcNmZ/AD2aHA0XvboB6xt1aRh6Z5nlvDslF
EV40w7zqNZ4JyNKMNxjxZ/PjD5Rh1rP4nV3K+ay+h+eTUMDzeTCCyT1RncxHfba2
B2Yh6Pc+NcSDMVX3Mzy2Rh9RNtyyl+FpjRpcj8XOhysbypM/QOr+KRnaxiayX6Ni
Yzd2WBjWYHMXE+cUQhR3Gdvd/cHBhAK54yVd+IzgIPcHndIffj75zFiKEeyfVqft
47RU90jDimtjAdcSQt9HMchP4H1IDIYmYrFI+iiGNFUsVUL10D3vQ6He0I3/GmaO
4Lr8hfyKZcbGWj0+dP2eY5sj/pBRFSeYixJXTRMoEozAjZta3ozddNvNvL6Twj4g
LrJa255B5C2+EYyHVP/i6+ltXdjYsuCppGPNTpc/sarTKvJw03X17M7bMlV30oI3
SI7Byl7TZ3Zuzgj8NJKP+X3wQh51ZBjvpSRwDWoGLCKCWCFxuzS/Yz3hjlpwu4tP
S2ZjSROMgZeO4lHukpbJRCXMfTCotxOHaeUKLLSOVR6tf96XIuLJyOOvPsnadpO7
qtU6wbE2qt9qDjq7ERIeLf875H8zjyrCxrZ7+ic+y8UPp0QI9gz7ps8leibWG8RP
a0bzO07yJokKXm8r5P1SSWWAF8D9Fv8czqj/TEztL4250ZORadYgyj9jZr4AeVIT
JJFiFTwJh432rJmub0r3hemVFCf5v+ednEqBvqlBHHBRHMxirVJJp9pSMHGdAPGG
NTmMleYXtxuZlbuIFI7etrlHROLQa/q4jj+zCl2gtYgnprJPVtO7hb/DhCrK6T5D
So2X7CtSWaxG+wiSUWueTptvh0UjK/VYsuVykD6TpH1WtogPOrQF3xC8xPE+ofqq
q1RMbig+xxK65T0wtogH9iVnhJM4H5QBUEdzhH271PymijaZrAIuTC7bgIk8eQwG
71zznscfSnBSDV3+BfeMZatRaRR/PONJGPcISH0BiTh7J7H98tHdkb1KMjwtoxFx
r5WoApo3xSX2pSe/j0DDxpMWXVt2kWbfz2vkWw9JTv8YClfDsi7MzWbCLqmLl0Y5
mL0VuWSgYZmLgGS/P6ma1cvQnm9+FeCq8gVzE4n1xM06YDZanlRkR9igE8d2nB8Z
RtoskZSgIGy9W64XmVyCgLvuzqEES2tTFULSSBXYedmbE+NqvWTxDeNdWX4oxPOA
1j3iWxdS3TwcZDi5cpDSw/enY4Q6juCyQn2xfIaWWqGVT2Ozx/k4WZ1OT12XkMw7
/d15gRc4HcXfEV8bGeMnLlJLs0CoSXjYMvVf2JRxUmK09ntqf719clZnTs91Yxya
TcnRIz+zNt5ut4PZuOHWySVbl3IT/3QyFEd9oolfXOf/fY9vF9xvtbKhQO3kogAA
FR89ZAGDE7BP0Dyi5yKw9NDgbB+luVQHl8rNBiLXYhY/0MqHdwGFqy6K8YZiXS7D
qXfanEXDDpCc5UWawWk69gEAHQ1oWRfO7+Jy3X4+vqg8Jv1E1rOCiuzEwn0oyhkC
sOZTfRwE7+JXQ+qocHK1Qb+vwUq+INM2X0uU0cCVOAyQz4CxExn75zriQNxyhG/z
9k2PGc4sbGGnUHVXxOgLyf07+NP7ETSQm5m2lkFcaBbyO7gVR9B5+NkSh3MupItc
5ysOZy5GZm14Xm6vm73CIo+PHV65xVFhTc/bhYqzdkOjb5HxkUNpDPmVbB9LVdgE
UmIX8pLKeI6G2sRZABxLlPPezTCDuEi730cSpy6L7TuUb6o7D/XeAZ9KcEm43RBJ
RDdbud6yTKPaeR7ug17aqaUGggUCdKADqtuLS52i+s2ZrqYX/3Td6jiKHUgNQsk3
9UIIXiBxyzgj1NI8vkKk3Kgdb8t7J9jyU9RRI2wEtbd+VGaH2UAFxRQxHOq0sQu7
cXjxOtuMJxGZLbffenq5Yxtk4/juVEOXPNgMwrcd5beDKW78PW6CjD0WDDg5sQ00
5vtj/o8h2oHzKQSOr6H+oI67dny3weOp1+6K1wxVGY+IHybFr5xJ16u8CDsjhvc2
LK3Y+s2Bhozaj6soUDw73xyMkRENsEZQPf9HMkGOAYDPXziiRcPwJJ7pPbfGpiqK
ge4v0d4iXVG/hhaK+xIF2GShDWbUFQTbXmhsAer7i6Beol7kJqQk29Qx+4Un0ekS
iScKXpFl+WiVl8493pPB/kiipbbu9gWnxK2TO4UJyvvnEUSKEAI+JXyQvOoeqMhB
WBHv6vpAZcGh8LgNoxUoFwA7XHEDGxXNw3HwwXUBob6QOl2ZS9DjUTlhLMTUAeHb
Tho4GEkkq6OeDwgefUHCnpDlj11UnBCNFl9Bf6j5HRUdTZ0D3Y0W3Woz5BSNq/IF
XetIbWP0oeEejQLLtVXfAHCb3d/gQ71A5FQVrW6E5+R4TBwurr6fwUb4Gqx9I8LF
ccU/MLBeZMeyhg88VBgLv22JVVXSkhGtFRwpdiDERK5u9XTHDxJf4P5ENHMlFs86
G3eDnIGdFVIA0UGhwQvUq8J84KxcIJ6AllLNymIUlAegl5BCMZxMoPQpIfKpeC+q
TjQgT01mm4HzT7q/qfYpTtwpbAfP3V4EA4H7/6kdIRZROdlh7wOX9DhgXfHS1Uy2
e4QNFNDzZ6vpGN3d28nioNI8fCnt7bzhAeqFMqYrs6ynsxc2/oPmmSZpKqf6/arM
4VeLsa5CIuR1cbnda/ZIdMir0XV+toN+TgQgzijGKOiijwWlgTc3CsIdxBxDSdKk
3EEaGXwd3w+rwsQiU8Pbiq1eIK9VnFzyY/iz0GVWWA+USWxSOlvofdNrOtEnlA77
LWuFEI4PwX4fnA+c0xoU60NSH3VN7L85EYRuYqsZQZ1oO+Gh576nSLz513ZtugRM
MLEl4Ehmr45s2HRa6k+0dO8dW/o+52n90v2TNlbNTIK3T4DEKaAAcYzoNkRQjx/8
I0xjOPPqIRCcag6345uU9vh+Semr99V36+gu6rkHkbiULX8m9qXjIYS97P0rJxTW
U+Fk/BLVfg7YMf0LkSfc+DRcLkdoT4D6kwMS/cp8k3CQ0OhNZIAFSJoxMLZQ9g6F
FktwgGNRFM14xADTqBLV+voMK4Kfn0RDJMQfCCXe8RZ2vcvMxY8oCy7wSSmcTSNW
sOdvEsKziM2OyxIVIEahsGUWsk+KaVT3pcT8OEgeEWCkn5kAg9hEUghag7r1cmX0
dfjd6LRRMXhTGfg1/FdWvtd0NXNbps0trl5JSNG9UG2l/5zTPpbAiuS0VexuSjje
slq5W5ba+yfWefbVvzHg18wT2DZ4/9i5rwsMIm8U1oPnFfZ1ZlmUYLX8k+HAkGJv
9ecanrQBjgcHcxvDAJZh0OgHNAgo2GEnx8DfuJZcBazfXcpug9xYT/n2WCLcc51I
pqqKlvDS5GCGD44NUdvzUP6uDys3HRYobMLRhsfhhm/hxTSEqrUydqk1ot26MUZ7
ArShfWtD1yEm/l8xinHCKwXEGkQxDcomsrDeMPjYgE6IezeVWIN6/1hgMczL12t8
5Y6f1lhEr341gV9UAZogH1fcRmIQYiql4WKhTcILPGhDCjAZF29zxZQ0rZvtyoh3
rxcxz5lf+oupUxO4A1gkhAgw42KgpC/2LLDRZZSfMuuNQ97lIayd9oOjesHygEc8
Lg3U52n5o9QwZqb1H+Hveb++ZoKgAET0rVXk2Z8pdXNWkEVym+h6Ard4A/38UYLt
xe/VKZkH0lUFcj2zRBc+QpRcCZhy47kqTgxU/0uFTsQHvxGjdlCDbYg4MqyL2Zuo
UiIABlwGK6MdjHJpkf89lxr+t4obgPe/4P5lPlY5J7dL9nAqokbVD8NAqcZOc2np
xzGi0G2g2MyBDPnv6+ssW2FoTM06kQustfe18/i4+2ibwQZSS28cSN8qZtKhfIx6
Cj1BP/0hgu6O8I+cqFWyYdeYOTch7EO0Wnx1bT9tUHJTeN1cYFEfRh2DpLtMGKU+
d7o/qeKjd8hFgx9w73BVKKGC9+GkKoV3pp3IshTooNYgZ96i9libFqNirWTJ8vc/
RaOId7Bwoq+pWr8DmSfGG0Dw4YlgnTprEgJX0VdQ1K7kOgYU4rlvbFxFRTUcNpCN
WDNsaEDGosqI9n0RR4JE9umXm/u4E5ul19lKphb8Zoh3ONrexETiO5xn1JBB2srm
P3dYL2gt0vUWeZ1Uikq4StRYIF8d1CbDAzIt3LD/LrhBoixvlsLDCCpVFs63u8sx
5+J/pzFDOr2/ZZVVyhgKDMuz1ut2hYKzmHlgE5xeKIkLNX8AtjqA75PjR0KI4FWP
VNVPBVVQF6VBYsLWI7uwlWjYMgFxzTGEbtYfKIURARiLfpYvzluEz44CO7z3gab7
3YvsW/4R+WQOOkIc6PE1FeZ3MWvB1QnlNk0uTfTbf1b5XSEMVGktcFLcRRw6mRQE
w1/LYxul752OdB4GPC5dbQhYZluue2voA3+FK4x/QUBP3zKWRv+2+1go7o82fOiU
gevjC8yLFx2oproRRf+9cIAi5uEZoz14Yrq1Yfeq6Zhiag8WFMi6F5OkZX7TMXu1
p62E06uVSTv4kYLtq43JC1OpoYl8yyt5ZvG1Q7uGQ++LjSMMpttgMFlDbM18jfsM
xeFYfaAeZ+Qpa5qHcC1tIsw74uQXGMPYKzaDW5E5QshIFb1bKIaC+As/tbDBfaxX
8VVaN1hzu2BVDMQPwzuRegnnPN1fnCNlfV+hKWNXH+KQ7fxqfkmdPRkf21w8X1/6
vjK7lBGjCLKxQIKGZiIwU6PmH3DggIdWlzYYjsPSCTaJktJxplEXW8FNMALsJ0nc
hZKDWdJsJc273hExhy25PY5mqoJbaYqzhCdoxyuWyLvdROxwkpNi8QuwNyc3TgKF
2j7HK1nn3sFdUajicEL3CXSgYIGnTiJXrQX4pFhhBF7NxcjwA3exvwIgcamtpN8c
R8EzWWv5wKsfifeluoCAwgVDXPRVleZBdFdDgFuHyKeSgjAPPGnqZN+zvPirAHjn
5KZSmhR6eBcAdjD8LETGJbCtbswrBQYji04XB6KaedSyk7w3laB8S2p/UvOi+/a4
cA1NCLwDFChuFHYgVdAt+npw0q5e5imYNXJ3Uw23S/XUr9kbaPi/ODPPXkgST3U/
k5RpehZafQHLXzIBDE/ZWFEd0PznyHpsasOD4AHHTisx08DWr0fdxmx6iRIeoPe8
lQsUWH1lEiJMqT5W7wBV809VQQjkTDwzny0pzM6CuW2WNl+eD0jtElwvj2gUmjX6
udGQwy2XpCrQsvYoCCW9IXRF7HKfECdP73Bbh8DAvMELa+ocBaOhq8O96g3k2iaa
eT3pvm9VVf1XYsw+mc+wgnaTu9G2vWSD8KmVVlZaVgQZmaeRnCrT+0LNBFnX14tv
gJUPuo5OmlbiJnLXgIeL2EVB/O3yZwRK8eR6VAdG6kEE2NdbMK8xca1mrEPJiX+p
SArZrK11bc3Jj8LBwYqODIRsFNixHpn2BwV62C7nk7cBGfNZnWAlrAJgf8VDzkCv
RjcXeJkMHZXkn1kdjOtsVjAuH/dmk+joUMaWca0M+ty2kDA5sArsYS7cBMicCNi9
8qRz4Mo+PK0vasHGan/ApTED2kJQoh2S64KZgrzsb1XJ7mcMwgc7lmUg3xX1/0S2
chvraQLBJV9pQ/GGU54xr/RqvLkN7SyzJKgN/KNhXKeAJN+KcXjJg8hSZG7peS80
dq+YOfyiH1G+pTcs8aFdHUEMIpaVOG3DtD3gC9IijK/s72rl0y/4ZBZqpuvzA45+
pgXqcYUVCBSIH+8kexkfBVqMevN42acnJvMqyRjxaxqq+NW+iWnlFjRsRk8VoTF9
/C7SqB9YU7ChWEFk6nTmiobrI60isY7arHxrzOTVxbZD/aCcI5v2fd8w9JfU1SX0
DgkSo6bbQAOZ9u98UJm9WXk0b6LKQ9vEG/h4QW045bvVChQw5zosecKT9Z5t+bjw
WDyF5eKCfVuU6ogVKmQD9D8IlYPYu3mahvWzoYywmWSGdpZGrZgkff5pB5NT6EJL
b68CkmYBVzi1goj0FTCq7n8RX5oUj4VGq5W0QcwQ37XTIuIMR6pRAEViUcAynCWi
Gf9m1kCd32jxaW+4aux+T6NxhlNHEJ9rswuoRqPwmwGvQojQU3HCBrKMd8QyMqiG
DzoLdU/yW4sIdFgaHNyr11YMrgpzsHlYSz7/Uas5X2aBxlrGy6Y54Kd2rDoAZ1s6
4eayGcpMp7j9fWY/gx0GQ9Q33WO49jwO95ITRSYWwVHpP+kG9kVQVHE83Rd1hQl1
3nLis+USfiPS7gHRrVOXunCCyNxwJjCdmhdTqZtThLNU8JO9A/USdGUXrMzOlVsD
twVbSRKGhfWj1ozHpfrN1VhSbgtwl2542oibQKxmyE/BdTjBleZOS9YQTrtt5Gy1
ulxVcgWwsCk5Nr9pHyD8TgzAcDeocK7+yBfHAmjTYW67oy91O8ykNyv1Fy/bt2tO
m449IeAO4i7CTXc3nBNv7WXSSGLFmWxmu09SeLPWOK7W6U9ec7TQVb2xWJ4/37UP
BOQer2zgDDeJsMJ5Qk828/F4hrm+g24h9bFgwR2quzsG2Xd1mrhrIW9t8Y9Pp+93
m0VJfSKADPxKOKlAKuHU5sV7nMtVIDznhwVhk1+JZ0cHwtBMO0ayzK+rtTBRtVDW
v5QkX+wqYHkUYPJkFhw3WmPGlr9T5lT0Rr4VYj0WqOhvCt+TZom8qWEr3zXSVEE7
xITknhShK+3EmmPS776Uz9DGLLwxfBGvwuoOg/sGramoY8XJIpoEjbbaYxuk9Y4U
1NkGfZpiHgfzlQQf/VA7qDGRWV9UK1VUi/WLw/w/3IP14Km9Hj6AgtnKc+GniiKD
03tL+uQ671g8JTZBXInfuosuhwF13TK/1XNRNqmu9Vh2AXwhRpkIA8xFHSO0pGuI
6OeAd44ASd0gCxiNSByxyKGQV1oQdUvizarj/Nw9+VLZWqPhvkeT/yeDQy+hI6g/
iTTvbg4uWFOxIMnfmk4rrbExTc/52TuSqo0w86UO+9IPWQMKjwTLGKJGNYqoY4yX
KI7mCT0CsrRDR9XDCAHZs26uxMdkC0SJ36FVSQrhYrLotLle7xO0bdT1oG8t5KtW
p++BC4l1Dhcpg6XjUxG1AC+kxCgxirzLKSnfxdOL5b6g4shd31O0XrkbPaPLOZkR
piJi2u/uSS54Z5E/TdtXvwHNNjvDbNl6hrPZcqd4fZyXxzephcjZsF73q7KAwef2
jWiTtlKhP6Fs5WsRpFv251c6Jt+cyvzFQ9WJtsgiI7OijkSLaxMXRxo/uAw4sRVi
5XQ5Rb7dmGQlduPhW/hy+A5Duh1u7CN6+SBm0iqxJRAE+6sTe6Gyu1QaqDbZsqBM
uAWRa6HRrXTdhUfBG3TMIl726/v6Z771yZD5mHlb14UPPY3YdWvKBcKCjZCbYjgw
oWnbcy0vdfstQOo5d5lmT1/Yp9CQUk1C6nTbNN1Pmkjsy8TjnYnZleB8ujYreXe0
shut6GEk6r2M+4dndnY4xFxsAmxL89CjCITTdi7lqTt7cxJDZYkEzstCNP6zzSxj
rU8Kw0wxvJjRjOx3altg2aJ1A1faw01BFdC128eATfGiLbGzKXNcRv/pYm8LUS3U
9r1UtjpAsEQfZVaHryE14CEvRwIPsup2QN9xCTQib/SEOuWkVC3L6msECFXhYeku
jdZVyJo6Mw0EQsd7HZJyuztU7ULjluJIYwTNwNAicxUl6WTGjd217x5CXsoAnAm/
hcLZvqVDYp7IRLvWGgLMVNCz40KkS362fgdVw+1POvEcr7bIqQw3eLR0gxSiPgqy
+M9tXNhDujE2aDbiWg8G+4IO+qt4mDxeRAEXxVwmW7ISBDgaidWD4RNY+1b5/Z+a
nIkJUjJK2p6SZWNu6GedH+HLGlZSLQtctFDmm8nH0LzMZa1tcUgihJSXiViy06Jw
cML08uBH99hfDkIpwLWqYHAdhmatTDpQHW/6cxMhLzxoAuzQLJ5sEC7b4vbWT8a0
mA5778njisIE/Vn7IMd6g2KwK46oEmYzUBQynRIRkpabHnZDDYGT7FAQzacpaU8O
vaeRR5CQwOk80a9mce90HO9LZM8Mr/+qHagnRoVjbQrtR9jObeWz2dht4PX4kbp9
0tmoGA66dyh9oICpxcGqxS54ctq4OoAtXyuZDC/gMDCuo9TpfDAfKX+gRiG4aAeR
9bf23Rb9l7UWlLkwctx293g58JLdypYj8dwfumbVyPHJOmS4LDatttc4OzqYhUzx
wnb4PQS1hG1Ez3n8HraiUHxn6JfSgn0/1RS5yPsMAS4o6gR6mFMIdU4UvZC+UXq1
XKG4c2sPLIeigKZpdD6PoK/fyRieMZaDvQeE69CvE+6S2tfKVfNRPLj743cs6p0A
wf/7odJ1KCWBp/3mBZvhQ7tzuK94MczZygTROjnodu4bjp8RUvyiFJtZt4tbyI+7
e/ILwz9vJqywrcwZngfC+Y2EAeBKrSLwPEr6fKstFMreks4a+JxxrQuJtwQGIsKG
aUv95rA7ZG1r4p+MQ4HVP0a5ZLmnpVNZcmoHQ1yvS08OTkfVS2OwgOpJlK+hSwb0
n9RAM039LVBmKNCySAwfdFSpgVDgNoiWLQR5v1plMa12nAjN6Z54SnXyecDW3aeA
Am4JxM18Qb8Tl/JGgtBVDQsYE3fUh7fGrvoU85hZO06cpFbaLjeRv+1byKpRR9Ve
eVuneG4sRTETvxhuKQa4leraHEkAi+PiSYTDeGn/q/OCqP2TxPhwOI6pRjkJrpkw
GK+IKNKwWkxm6aVPeJ1MLZD2Kyjgimhc7PYr7ZhjQHcllfsjpBQZthDV0Y9SPlEQ
zQV/O8qoLBzklT2td4fIkbvrcRBD6TEY8zS9yOFmnrcwQbiRHW4l833FOptpgKc+
F+Lm+f7DZ1Pgdzo2WuqCcD3hkCpESkAa3f6fz2iG/09VMf1L1okgiCdIhI0Yf7XF
N/FfUGKstG3sR11KDf/AyU6y7vVHeihZxVTTwyEL8Yk5nz85f+eCS8UEkdmrnITi
Wz2mNBTABgQIh7r3E2ehzp0S4wRf6S6M73P1DCkCZj6mCVjaK2qOVbQ+tkTrNoev
YKL8ZxQKoAbitc3lBOzfndU0Lfh9NkbhBNLSF72DdklyYCls2ht6FGtWAmIDBaWB
3kdeIfgAFX/grJxqKtc1cCGII4KzS/QeRcKxhdIZpx37ylQBC0mjQvr350fGNpCZ
kAQmFkp5XdADg0iq/pbl5Q5g5Q2Z71YPejfIYJoUUVdtRM5UmDcjP3eJiEPoVwK9
KTxTFsx1UwyL4oVKdgfOVI/84Gs8ryvibUycLF64+ZbvEA8QS3YBeXN8QQdKvSCc
p7afYQBr3w0ZIMSzgPchx3Jx/6+Ie7PuGMemHYSPD5mCQG83LDtqvrZuSgIFDfq6
7ORfGm1gsihlWbvzUPdzt/2JOzbSaVmE5YzTPSxXotOPK21/GyZQqGSflmDmagxr
GbORK6zBk8E7CwC3d1xQYa+PU9ndOGUc4RArAWXGy9crC/M/AG+5WtfC0qMe8XKz
oyjTEBATLsXGsmmmvXwpoVuJhychWKuutvBKG1G9fXgSv3Ae+xSE/WY7nWnv6VY2
pSU+5wwxP19s+RWReDmXLu8fTe0eYSqpV1qrMNDKefnr9sJoqRmDHhKVOG8RS6RV
kvp2eHSIdLEG0JVTaokYpPPW5Z2hbuaJTnv+CKqY86eONzP+RQN8FudFb3CO8QyG
QuYg4MFStjBtXK2yPsq7WOdTbwU8FxVysojn05DeasGx3b91LJNq1q0fHN21bk9v
L0vYvedL/tcDcp9OWZaU4R8ftapfchH0T1rmCAgEmyrv2nUwWUux24DY6ODLuv1a
qDX//I0QNHdD9+jTEkViVbldN/tOXrcTnMx31kP5PyZHvaEjJJr/HC1wlhAgOQdq
Jbd/GCqMw9esRlBmSv0GlVrKaKgR8nMKmQ1PLYKkeYXJ1daRZD3H8tcMHazC43yY
3JGgBqxrSW7/692vabxwOrsMpTQRw+Lw6ROrkOzKYFydE1ZWtEMLHoI94IcIPUtt
gQX0Dvdvibij+qNCSfZCXWADajkIQl7Aid1LMnapyHsLarDjAuNyCSuI5GH8LOmi
wXycgbx4hLSwZdCzJ6DqlR+r5y0ewj5jcd44iUlAPM7abd6L6V1G7Mcsw/dBxHWM
j3BRZHQCeusET8ugD79gR8dhfz3YTxt3ub/h8y3YGMrmMU5SXJgTB0/Htr1gay1L
rPYngI7b0BBmpOVo51QkheL0LvZC6Yjbj+x5z6enCM8F3T2GZAeb8WYX9IRvr2z5
LgrA9yh+6bv4IMGmyc54z25bXIChgxJQShOsN27RPwrJ/hrphA5w6RDAwLkV/KOP
0h9Qn7oOI+UaF9pI7cpdiBAoihm5KEovSQzU7fW3bprXjbTiYt+jYdrM6/HUIKJ/
LHGpCEKb0g1swSsMqDD2mlAVjq9/LkAvDc5dF72NCH+YqJhuKCwsp+N+/kk5oVNa
879wRNtc/RXOZLZZK7X+WS7jXIzicseNlmrxNKIrOgKRE2YylfweN2FlmlUsS19n
Ou1YRMuOr8l7xZAooM12qBjFhCk1/7eNofh67gAboCD3Q+8RHFrBRIA2A8L6t7WV
c2evlxLUAjBfzavhRK+rzvE/Q3Zau3abRmQ2fG2++sWRxfj7aA/5DrS07OYUG/mz
TSsTcmtotW1FyXymIqM1JhvhVBIhFfpfR/P7Na2sDnSjn6gHEHVAR/s+mAMz0+2t
d2MmYW4pp2IVdNPi0UTFTn5mC6ADFQVBpEyhyz/2y3OGYeOOuXPWsQW7aWNM7qxj
BLAv0a0qX24IjnjUDxZHhFtbOAMHkAivEEtjABxFzD4GpmeXrGWCI0MDhE49OtNi
iGgYN92XprwVx8EgtyjyFnn7BhduRvywswKly4XK24qJy/eC3Va+zpNJ2JJ5M31Z
9Zz8EM/vdglQvuYsqxq2sS6drY6qhvI5JI69UH6sLedtQv3RqKkeZ0xNNvvtUe9H
WviKHAGslBc8/vRastRwvihMUn5FqkUx4WfqdXfqm0JhIxtqh4QYU2eqyzzVx27+
CJJQr3OpRZXb41zcQXyhlegqLCxK9PLVPTbUfJBni/VBvtR5H08IPSyYYgUrZNKD
O+d/+Z8GZccJCkgo7qZTceF4sMKPmaABZAOqmC8P6sesb5LN7vBBaMysGCHZ6Qsz
u1HSVKoSbjRTo9/nb80KXF8KXnPNMYujTOCZshfcNLslCfY1pidY0QcLVmoy90nb
EsFq2eBcxt+yf2tiJQ38C7fZ4FtTnE0bpJ9UwKPHRkh8+4v6+TnfnLS8CMsWz9Z3
w2B/+YMv+85sEPURS/Q2Zg2cpMGIi/C8EKFeodHIobYW8pPcJ84cUAHyU9lngkmh
7COR4d2k+jbubfgM2JSr6wXzB7UAazLbsP4N8fI7sRHo/zGOP2gHLVt+cJeYuVvF
gBJ/BpC8nuasRUzdIwE+yy64/Kp4eVAeiUjzaufDv2Xi2Ru0VDgv+GYw5gxXBqsy
5v/rK9jmwk908bvxAcv1+GCGUNJ5z48gFNCC3c6mKrzpbm6MSa120iUs0RvjJ8QY
778B24+MAzYAwUglthdqCwkS1ssQw0wCm0vQmz50BXO+Vd1kIDpRFLsmlDMlo6vg
RcamapW9UBbHJHdnbKu/aJDL9ktlQMh5eyXLzFCH4oG/sYYiYH+8sQLXE7XfUtwN
eev5Nnj4+GKFOfqTywQFqi63pjwb6ylpmI3mPQNmNVokkZgMr1lQ/I2oNBDmQNGc
QQxb7FkNFb+OzTv1es77dAvH/8tFf2v5Ad9QqTMjfD81DDgkXWYa0vpl3dsSbV04
2g3W8KKANaQ/TGLVqByuZhPtRpk4OCvNSkn5fVu4J3MEfslJ707Sky9G34g+qwoA
Fr2s834Pkpe3r8/iZYT48NUKcdVXEgoV5y1z+kfsYMZ5hKVtX5oIiGaut+4gwIo7
zTrQQhJlFKd7lYRJJbKGwZuaNPQFqYsNtAUBz5Mw0wX692KLi65364mJX7lblXx7
KoGI3vanRmay6y3EZX0rrbTYFSmYN864vSvcVmsWyyeUxK+Oa9ACZKETDcCyPh1E
Ki+MkzmloIcIOrGXjq2PrUZvKn2O7oTYXqARG/mo7zwGD2lnz1UCBW5Gq65Y9hsq
hQFOoNCOZcsBBVGoo98Jdcf87Jio3+C/jwsW+DcWr2hP6YrGikZjFSCUSc/7Vaks
v6PBV2ug+0T+2OHVg4/F6egHGz0rPUFgULjM1d6BbKQY//1qx3xbR3PbEIlDNWFs
1JMYuoGWpDwQpjMobghDsgQ2U6/v5TMtIl3HPHftNUnfqrasjvtWJr3On5n+9/9l
hveCrjW2L3ho15nQ5HZ7GlvF2WB3OxOk94bB0+XtyQ7XIn3/T5ZURPm79PV6xpm+
pfGi9lWEKNZnxaCAHSehO40ZVXVj4xchEolMw4k0HeKvSgNzizQCDop2V8UtBG67
MBre96nZRgKquq2rNgRtQC5QIzeqWB0FjXqi//bB7qdHFGsqkJSEUASpNEoRoFlz
3HuvPNX6/Ma8ZA/x3MrRkaikFeDWgL1MU/5RhefI/TR8FPBDPTIbdJdbmzn8T7m8
wGA83ceFph6HKsVqoaRuU23mkP3dBBR5PN9vtymP28faGKHbLMXNC/sDDs/QOsJK
KOHXsz5m4i4fmaPNUXch71Wms/TZIk9F/GYb3uIo43fSqhcgaud3NJQFJHbsqPJW
cTeoDfVP3xTvqGxWL6elx9p5mpX9b4h1XnzMjqRLUiOWTr7CljA+5t9MbG/XbMaZ
VWcsXiy2f7RxInHNdJRNIxI8czGl3iEQaWHM+eYuK4UYSUQM3aQ+/vgCUneSdWsA
rJ3RUyFSUQUqIeba/qoYIXLPcPawylOKMyoZPBdiRtFZhJk/cxQ4K1KE9t8OtYVw
MUskra8fQliB+2PKMnfwhz9+UBTn4YgOOUxNfO4z96FHX3rBk5j1k/wCABolt6Cp
g4xzvxg+aKYjYlzIGPdnV5QJphN3tFIVsGzOXDFq/yv3i3RbmfHQQGJz35lzvezI
fwGueKh1BEdjQ/Iz4Ir1or3j2Nm77lP4xg0fwwmHw1TMc79IjNZ6cZBFi0HfRKZ9
iV1temwOchB8WcwHvugh4Gr9C9s6M0t+shoCfdMBrrS5AAkolWIpFw3jKPffTFSz
/04XlOAke7V++wGBZT2HGJ3p8xSEmrhKIpgypo4zkvoWu1Mw3CxTn02ohGFJT7Ep
OqaBVvEVoDw1eBrcEWZqyiXHdm+1zxjtIKKWLZGqcLu2k5lQPpijeAPNfKagEbMZ
pELkpFcs2KLq4PjjUVC0TqKWst9h3DeE/CfqAhaggkZ67ZlmphtgC66UDaBzXzTy
vgL59H+nuB1k2OO943bgl/Fk8ttlZbjlfakLa9BHmfEgiwvBoEm0EI5T8ozTj5pR
Xe5QCmDOBJAAUxOBy+zcZksxlfRuD5phcrNkZy0sPBVM8GJbOiPqEQBom5A+2fEc
woRp6ALUDV2IemGKHBWiPsrd37YpAuPzIpyMnS9P31XXIhkhjqL5LbKOrglGC2QL
kxZ6PuqHgW0NmkukYvMlYQjrH1oxElE4b7pnSkxO3DspFGVJ49KMMAkl7FqWUj2C
JD0OtVq4qkLuSwgjSc7keJKhtjPFw5tJPmZIjZIow0T3qnE72HW5vrK5e6xddjqH
jWqC5ZFkLQYLnp5veCUAY9XD53AHh61CJzj73X5aSC07jvmTQIjjS7LPjoeTMD5g
jn52iQexzPP75EuPYaxzTryoE9DmXwlFyr/93GuHczYRq+cw+kgZBref1CsdqCcw
BjxsFAp4HxxfaRF6YHTAlrZLPhTq23/0Ig4TKhDvzRSGiYXZC/gaQaSGi4jJ+s8V
XjC3/CvRo+mbfs/NG7L4W7L3NvOfs9cQv08HIAsCikh+j4D0362hN5fNaRZ2302S
XQ0S7ThmseIQczkAYNpogdrZgX4e2/7116F812SEM7Gia2zJLr1Rv21CrVxtXF1H
SzdZod+LjFiunwzVcniZCTclm7JrLBkBAZ+mALxGXQQ1/pCyP+5xIn1HuHsjw9l8
IXYPyZn77kRFLyImcMoyS7tHXiDN/MI6CC/0ZuQPgfatNyiEdubDmi2leiD1q6GO
qHh2PsS+MnIIRM1UmwHCqxA7OxVesN9iHepLUpmoc28gbhh6QD+0ahCxdFK8aEh+
rW7YleOPSllibQr9rt8GQYp8xXZW7xPW6tcvyZRKead26GOiNxBd03gGDOm+7XbX
UuGfKY29ZJ4uUDpRVvDMXF+eJFqvKV2YygSVsYmNeU1PQt+qN8rSUHzmMjoFNUTr
Ga9Hw4GsKTUlinEmMH62q7XgLBQnW033zqFcuK2eN9VVrGfep54XyLzfCSk0awXm
MiwU19zwZIkI7jW0auz/de+LagRqvlezPwFJxOEiDIr5pTAKP4LFyyCKSVz+iLPS
lDiDzhOlKMcrLKFcYlpe37A2PfYshFA98IrCLNwdQ90b69iH1U8UjcyHPlH4LvqM
o56DxKNez14TeSwDiL6OvsMFPgxL5Zc3SQCOm12aSxRe27BqlZs3rhg2pmb2R/N2
OukBfs0YVR+X0eMLOxwA+9ifOUN12nYNPjlBm1G5DybrRPIbiq49jyDqteiNWETJ
zHwBBh75nWpgdnYVagS0+n6kjHbdoGP9MDN+q5jCGGfXCx56Ija1B0pd5dzz94Lo
bxhNAJEfdgMkUMjHcTIoa40yvzapNnQdTbesbJwdJGXLmGnP94g4kcy+1pfpvEJT
WGrRVmQh2KboI+7yX8O9pN8/EVqac2xW/rqiy8J6Pw3sdjb5mEVijHlig5IkkWpT
wmMh8Pu7qgRkaEdqtOhp4KqksohhGUB8pFaLllCeV5n3tCRgP+VAgxSDFtJWUR3S
Yiz9L8Y3/OAIE425tHGE6OROlxWdNU5XgnB+17q6+GWIQCqlnALN50+ihv1DG7C+
NIpNh+X8R5/JijmiPxZO4j66d/gRIXq4CRJy0P9Nlg0y2ltmLiitkYTFZBGmVVpl
xceizoeu98YiOAi+EVgWlQ7W7m66g6mc1YpPIK7BM8sZE21imNJrnEDL38fsYoEo
ln+FvZ+zn3HQUkE6Qxw6rlhe/jvZQHXus2rzvypzrHRkfODAS5EdRKDTlbNEG3gD
WrexYKyGHoPvYtjsioZ9WgBOgt0w1JdGpLSKwgC9bPpGd3flPPorx1A24kPJV4hw
5KAnO0jsrjP56hDgHlqpJlwPSCzYpRZAndI4ek8EJ9ixUljYgW4LlSNU55jcklbX
c77/ftSqRhpc7FDIeX5desFOKIWn8dPsdpEU9b96/6Hri2cJ2UWynOoQnxT71cZM
XWa+8Ac+TrLmecAwJcv4tsGH3SjGwsueiDDvDWuwB+VGsfYyhxuCbQzln32tsjbK
SWKPuSZ7qiLrPywzKhQ8P3Su+ISYIzo1kZUMITyWvYMfvUEMsWDo/0Ljw2Gf37AB
uPZXEyc6wHMWEdcaiBDidnSOrWtgoRzkQxhcSNpt36dt6IfxcnBic9D0pucTtBoe
qy1OVN4MxcuQLn5rMlivTKIGVj4YBrv/okrgV+kQzlvI8D8SgR0duaOiIIX9b4Jt
Sw9B9yrYm+mRwsnYeP5vOWnkxpePE16xtPzyzs0fu3VgbKZgVxlhPmDUEOZe64Vw
UK7kU5iHPnV80uD9n4dOx17gSqaX1QDx6zrnESj45vPWx0Z6GF9lAT0xCFq7j60T
9JIUyLrksDVyWelXm8T/eVa8cj9Gdz1E0whfmzsZ9A3ye76U20GiYM1YInZsa0nL
LR70fcjpy0L4JGwlCzx0qAS9xsnCdnG8zPxOHD9scplIgZxm6zoQhyTUPwQqBGnP
FrFaVNPV4w4Wpmp0QHbnuB3/HoAAY2brCjSsixeC/9zTmhRouXz4BjkciTw4l1aq
FNDp+dlI98gY7cyXE3EJxwOeiKzDl4lboP4n6n35g0wucVxlgSyRyr95x9AA8vpI
Su+xsbD0VKMkvG7QsVeIYg+pUqHgeRP2c01ugs9vqR3rQhtOylZDY2V2lKZKk8Vm
SnGBaeTAZC6PjOmwkaUqyoqTioPrTlMxknmigLB8QcnSouZTfrgBfVGyuPFUHtLH
QE32/OJotHTxcF/xjUGSNTL56d/v0Iwq0R55Tz8dsKXJXbEcKU3h97ScdtAoCQ7R
KIfYNZmXan3X1BRf3yfIvtDL3RxbCkdytipDkkFhb5rVGrrUv+3FJNkJUjknDDNb
ZMhuG1ANwTB77VhQ+BWG1mrAO/EILuZjKMe3Tgn5JtoM//rK7yihJ88ZNRDub5K8
AthwyAQUSC+z9IZAYJqV8cL11lscDNW/Kuv/duW2nNFcgeE5u4jR1oSDxVhQf1TG
As96N98sUlKNJuJD7ec4Qtl2BM4uCkQTQORZb8xG/COnTtAfSfCs/62QWRvT/RqL
BFMHo5x9TjsiK/KnXOy/giPcULMDEggjsmuNUUHqBrtif/AR/zoCm1WL8WCoxhqb
jvh6G24RPq/nkqB2qaeNOKoi0RQjdP4of60wFusESmHR0LcqgePPykt8/8JuIkyh
2aRW5paNg4MGVRDQoWYjgY5w0tSP/5rPV+mJuG58khCr7KKSlCU+1RiZcnmNmZ6R
Yv3Gzp53NEqnKP3/vnyNJ6zSzxyeZCGb28IiyGaqz/+WkgI0eLfZBInwMrzCfLmC
eRbyfHzELveWMFweeA0Bp4GhbZPqRWyMlb85JqB4J5G6Bl1ebHDInMrXCS+NuGbf
97w5inSxIuoICovWTrFTE2ZaHM8kbFrBJnKV7D2tljWo8HRlmIdwc6wgmDYiAZbI
rmkCDpTuWUT9NJ5AJfb6KJRyuzRSDn02/6WaSgf70eMixR674uJRWq7NZ/LmdNjI
HqKyR7jzwIEqso0loOZ4ZSQOImC0qVHbavXWr0fVEh5ZqxJHtieFfhPw6j1nImbf
i3fOpLY5JlndNMxp43IPukE2xODe1YX8su2p7zkdCANIqQ7YQ61Scoqwt1hBLery
/i5tHReFZpDOmQ42wfefH3H/UlUMRT4QamXdkt1qChxGSQxjOQqesYf9j+VdpJMe
vLFdqEZckcfSzAVe2AHBHlztRqd0xV0KLd162OL1JibaeIsRAyRVlLzVVFm3xLtH
4TDzaX6eiCtame/GpDncrSA7MngHfAmPwxDheWXGr/hkeOcUnLFbLALI8IclsAVv
95de0p/udTYFclkhQLhtDonWTf0nNiiA8+n7VDrtLBsrGP4CEYGLDie+NF0AspGn
VAKSEFcQ2+u46Eaz1zcd9DtRU4UeyYcuYUbYlTv4MegDpIlbNYHsIkVv6rrGjy2v
cfNtcFRZ0ZNQb/cwW1ThsZsQ406x4KL8Je4xyUQkZi0Y8hixTzGCvVX/WShKcNjn
WwjAZ5EnhqMcv0z/J5PfK4euCPdSMM3j6b7LpyrUfTi/7UP8QoycwfJA8/l4CMdk
70Ki/LjOeTVOOE3ajlvfhNKv42S+9QyHZwo2zrUcVWmrUvpsBRYlei7Pm1VUnf58
HqdLL2kZL0nFjsYsdPu8Qfeaqpad/F7XkCW9+Sf5oafBAv3DJ8BoQ9uKcCMuh9hR
tDW5+yLvgmhioGTHMDI+PRV8r3GmXXZzBcs1Drjc4BXGfrwzZWDpmUVo4fOu60nE
M2EOLhvygrijR0GOoPei6Z14q9y7a0LnD/6Vh5kyMIB3PLUJfuQcPk+TAUW1wvyZ
WtxR6CaOxOFq1C2kyr6/tPQHbRwV9Q8wJTofqYqwYDXovSpsXxrN5hCxKaRsacjI
Z8eheoDnlmQkClJS9qtG1ic7OaH66XbYrIZiH0zUZiF/O/SM83ee4NN5oy8dq0Py
Vi2VbpUloPuQkGOyhseZS+fjnFj1kY20AkTuo7wBWhH/RH4cRUL0D7X4K3zMOdH0
JhMp+ukzho4sWEy2RloTuj9KsjbeN/bhLNG9fZP94r5n2Yivw39mdtX6rkdFA17E
jPRtJQ0Yx0emaFMCmeCOtELoMJm693t5U24gLcipBqJjC76hCEBsApduzAH21ohz
Nt/ReXVWwVS5LALkrTYTZEupTX0EvICtrkVRn8i9pBeKkeSm9RbwVXerQ8LaD180
AL7FYz80cHlbqQO6Q1oEn+7tNRVuK9o9J3qkNKuMDPaNlpm5nnkbwNJ32VBFDy3V
TMaZDBGhWjQ+y2JuVqwdS+ZP4xCqnFTBakewoo20NVYr0AT7Vreh03oO+rwysY4j
M8bhFCnRRddWKwytrHx680vSXnq6mqRHmXdKnOKqjNLw7zTH6FFeZe+JWrNHtHl/
sWeysubOCz1tPUPk8X3PS1gcjbEyrhPtuQM+z1UiNnNM23uJkhtOXss2dkT73/AF
Nr9TEYjD/B/Ch3biimRoMX0712/jDK1h72oRs5agw8ETXoeYUVZJNbuVSCbG+EPC
dl1k5wjdqAwB6AlctTA/XpnuRoXhJW5yw8H6RoW7Iy/d8g/vafqbEfYcddJTXp84
zL08xIl5GmjnDx7XO1HglrOevh6PQWXLKmdq0STYPEFDth+lPMNRI0WfAlmvguTi
k9hVUp08qEIDxZlBUuT+OoN1GYgH6dxqJ5uiuwyYj8lz30Bq4435rWgwnxRJtXtF
+paOeMrzmjDjnikEwM4OjWNPcEemAulveSBCckEc1Jga3nQmRDg5m43Wiauqb/M9
65gzGGitKmCbCUhz3AgXUr1U9fl/t+8zI0c88jFGu0rTe0RK+wSSXZs62JJv7dP2
GLrAVV4TXnqR5NH2GaiS5m4fpk3UcMBUFUN8ktyqY9ncd3esZj/Fxp8KQ65aaez/
8Fe/LlG7B9iquVxXUnzW0uQiTRGbHj7Kihjq61Mfgi8MSjP81/rd5VdSN2El54Nv
Atyh2ZvQDNBqnTKCuguiM7YRWBvS9k6S8KfgGrQaHPbgDbWsJRdC9jQqCxe6v9Hv
sG22g4lbSpG2DWpUp2SUKK5ebbIBKsCLk7mDRGRAAcbkWExiTh9Y6FnFUBTylrUR
i7Lf1QRhUfzpmmLzkxojWh5Pigy1TbRPoAuCdrZEqQnjWog3ZcD2sHZXqCVwfp6u
Bta5Fule6OG6QuY7UhzpORHPxcHl+B+rKYHeNznrUT+LaoEqYHSeVBWgfVd1pYHD
lrvZaoW1W888Ix6ElIXvPb/4O48tgcwtTnXrX/oXl9oGBC+x64CEE0d3at/tQODp
csDL4d4bSxfXa3/flH5Fib9Z7VqCpL2NDp3rNLlGbIcawzGNTg5cndfca9G85+8x
Z1wdePn4KcGfKAmqKrEmve0FXkXdn8ZgcNfdgb3c/Rsg82YDTE7Cb+x8M7f+vNFH
lpFqk/JrwamfWvcd4pz7gx/6YJ39l0J66YFhcxPigr2gqhMkCuNf2kdhyf/6N90r
sSHFAa6+vczW4SsAuRn8RDHXv4DLBCE4jJsrsZOXgUwcf8wkoyWvXV+P+UTxexC1
uaSbo9j8qCx9HotPWQG/JEqJ2MnNdLv5FgXSWEcsKYP2divXU1++sk+nv+9BWFCO
2SpuYEIUx/6qHFzg8K1yt0vNvig/uV7PPCLlVKxoBDIaxYaVScAbboD77DmTnV3f
RVH5B3TFhyO6CR3ZgqyFjTGBODTMYKW8+B9WR1MztqfGaM254AsyHIXDgQF/3EkM
VIQuUIkCvX9rQR9BoZn17X40iLCz73hs1vIdFJ+JPMzb6qa4MZxFMKuiaHDtXgK/
eqQEJKURfFZNOa/Z0uyyYwqZ3nL9rQjalWd+XM6+cd9GB+w0vGgHmcP580JyVNPB
RnOPWimbwbr/BulXO+MrY0qUClD1Oh/q8hbUZj5JW8jpF29O7Rk8NAWKZkzSGOvi
SQfNM7nRTEMKpUTygbSdV3IGESZ4g/pXUDOfatYATDWt0okcM6e9JeUMl37BoDTA
B1sUO/TUbz738ib7hXmS+vK1cCiysPsaYs4+bQ2djNVTsTtsX4lDOmUG0TKXVNM6
Ek8sqzhvl820n2Ol5YxEPivm8Y379ObYh1EMOY25+QTqP9Vk9SyqAQP3vjJyhifk
N7tCBGxblTPsub1poR4d2/D2WxeF+VboLSC95ydMd5luNyJ7rqvOu3AUiM8bh5UX
fMsVz/CNHrfEeQerLEMlv59BYd0be3a1xIaJ6Pl+866NrTi51C5Ukgg+EK4AP3Lk
0BeKLi8k6qruiNhsE1QrSM1FX7lBf1XqcPK/tDPfJ7fSlXkF3SQ8fIs9+rwvbUQM
6qBU0yAsa2fPPLZV3VAgZFT7+iHsqNFj9yoLsdmVF4qZTfnGBbFSvnDCxgt+hFVX
BHSH2/iWph9j6CXtMF23sbRjk/23OjkyIw/jLmcsLDryva0srSLYwDg/L+ZEvuHz
JKWrBJUj6AlIZ88IhEMQZY1BMG/P91KzYmb8VUslnVuLmYExreGF+cuPidwxc0TM
HCvL6w50NM5Tw8kt3JhuJ2i3dbS6eKutX4DmaPRhE4VE+7sbP/z0dU045ik57gh8
dcajgGxFs1c9kPxBj6biC9Tz251qwQnPBw4N6qv9dXUe/aaS6Q0tMRsDj1FoHtgb
qeOWb/EbAcZvGu8XYvEF//Lmno155vEjgp6CZTqaFeQ8arLE5SrVA4dPxmEJu5wT
ti0KXZcrVw57egvakyRENg6JE2g5cX7JhMFdEfZIBMamMKZUPO3uHEk5/KaoXiMI
gb4jOKuxX6l70iOySbX5HTFED/b2/z/IWbVUoIlWEPZqqnFuLaUTT6y0qge0C2Z1
bsMPv+fTAPc247m0xIVdEkv0sGB/eh5akFN3Y3fJ3lTbfwzFzVH3JfHakTb2BMk4
BQf9u8Vzu1KYPfS89yNYsfQ6v0NabVjmY+Z768P6Tn1K7NzYsJ5eoVz7tyogHpzM
DcneRMvjLavYhz4Mf0viaCo9i7wJvcGEbK3vv06HBuj3dDWCsgX7mmb3OFMRMQAt
mUTlKLoIQRy8oGq8c3F7RXZ3DxBnzKvi3lm+joQ6jBJjOlDOxbwmELUaLW4jj5ra
Mj7k7AKOxueEwm44C2iFDz1KS67k9r4UQWu49qYJ/9bLsa8dblwREwYAZSTxs6nZ
/Dbqq0lp6+A0Cj46tGWGAjFzzDvoUpxPXu0UCzWg1mVt7MwJvU92n9j4YYNioYBw
oyhdKUSXF6wsee40Ccwn4E/KOUNgBu/FRCM+T/RRGsYCUoK0rFDZJo/VMVNwaB6N
4MffyliawHY/aScktEf4jyWp+vyfBBImsphJIvM6YtopwhziBhFFFWSFw0iwTT5s
7oJ5VUBJ8JKlo+u9GtAc1A3v/qP636W/XE5zuObiYTAYVsKi+dDQHHbwYUOM8P6+
XvOQ9Wlx6+6sMDIvogvxWh5YwuO3KOCGpRODvPMJrcyroBGSbESIJGSMpWN2vmNE
7RAA3FJymd3GfSNpYKrP8Sn+zDqwK4Dbx+YKCH+3mXvYYdFZ1UJfqoCctxcUm+92
oh/f2FU3xXhlzBRgsLESFTYUT16eGG5W2x8Xi/evmZczime0gBQliYzES6Bpriao
IVTIzkqPep/j1NgLDjM8HqBtGCWpNUdnvvJGvI4rQQfRKrt98uHf9EcaHfzzEXvS
J+6DsaF9H1OhrPWgx9100SkLvsO1NmLaGHEUSijhiL91vEaQAq/PqWprcEUzMX2N
k1CH1P+NkzzczW0Uod3ULBbDPc+NudeqfoVz33ymrvm8MNQx88KNtcs7dEmaB1yn
fsCW0jXSyV3i1Ty1anPNTpIoq2Y8M+qnqxy3wGx/+w+03BE+9nRWcBloJ7w24hnI
rJLkFNuSEWBQou1nCKxkdyrTNl+Ghz4f2gjb0i9t88RqDUuVbjq1UKgAvEFqvV2L
6Fm1H+qhhCaYyUAZmbCOmarz8U67uhHveOiRbH9lgy4MdkbjkM+yWUmgl4i2aSbr
X8+3HTE4fhMZZ658Gn3hYeODLVeq5rCWZCLf3lhx1fNkh5kVgXviujh8QjFS/tSr
qlMOPYixed1V9jCFzXofSbWj+oukXWVd8oKrWOoUXZR2jlQZa02+nEK+v/Y3JFFs
JdsTvywOeP2ALKe+4daWgPvmBAdHfgzCugnQKWUgwR4IdsIcxLWqP/mHwe6jDfF1
wvng5TyTj82jLYnpfjak7aGBKr0df0WxXkg2AM9QunUKmXXmcn9gl3fiMlrvLAV/
krB9gQOXSPO+CjiZDRmrpDKtG64AS8MMu3P5scrLhJseCvGBbqy5NrjU4ur4vIee
X2rw/AjZ9IvrEQo8LuHOO0X17EZKe+zqe5nPYsf1shLDyUo+xg8GGulu2Dw8WHMm
J/2cklYoUOE3i2AKZPm4tadNcm5Cu1VQCwUiQ6aF64Zvyqb+xgdsf/PqeKOA23pc
KKm0VA5291esvN5M4BfxKB/6vZ3GXYAC+m3zgec5a9rNQqaNhi7L9gI5jeSosrqT
gbdvJvvqk7EAToCWPv4opFBbLUKLs+hIZS1VPKNDse/hSv6gVTQutNr91LuJSi8K
2oPbajTYbztObd3CEx7EirJxywt/NifBjNvcWtbUKyKJjphmNu5eAXoJ25RxSVsu
t7MGMeoJZDakMnoDudx8TFxCsxwDJFmAWSmEQxCtAz5h+ijOzK/RV/qx1Yuq7paA
bBjsEVzxXUgK3OKhy14lt2+VeMioGptyeR1Dcvu4iZKw3TEWPyeb2M5HUhRBPo8g
1wxPthGVy9oMelOXG1FlCg/8O/8F+MwqqP/HrvaUMzv5D8Fc4gINl6E3N2KtTv8y
PCZzidPD+Q/6XnF28EnyR0m6Fy+mRNP6rqTle4F7pc72V/NKH0/2fK3iWumSTRRJ
PR+h6yMGyButMoOa/2RbMuYEGemtQBklwr/ySZIGORFWHp3A+dWIF8m9ZtcSqVz2
L8VG226Nhj9zeWvKpR2e7Ybr6fzEwVAOmJQGDI0TLPDCFWHO1OB8iM4meyLwT9ta
/UHLOk8soshKRcDajT0KsQrxpIci+MmVk1rGLvQtTEdvO/KKhGKziJ5TeRNiXJkO
a5vF0DIKl9Rrhwy/RFk+Fd/k18WBos0pzdw2+nMuTBpsyz691FIdpdUQqj2vvN0+
BN99C93Jdn9mJYiuJvuPCd3XYecw0gJMNE0J01tpXBRNuIWM1qj/sC1chnLrvGCR
yHfUyysoxZU7Ynhx5Im4WIMKGwklgvb0/Y/C0n1Qd4RZXD60d+QcbskUQQD0sNrm
CgEcRVXz9OdQdG+wAAwaeJGCMuy6+VDcz3L7Q15ND0td7WoPyFN9tq1/YtWMyPXd
zGZ5xi7JAe9T2TtYpXP4up8nsboHvBI3ghJAGKfaeJOfS9LS6TgACcDOQCiszOor
aaVO4l+lu6G11wwIdGz592LrBWY2QhNLESk7l9pygQk+tdJgn1GO3CqklBbzymyI
C/rb1wtpQ9TDOG5GdkAPGZomS3mdCmmPyVXvAsq/6QnoxJ6vAAziaEN+cNNafKUb
VmZXCRCcPkzPCeDhF3L12T0Wd/FvpERnOJolAegjQWgJ/lvhnqSAZOdsTfDzz3KB
bkOoa7fXw8DIoRpXVHEadCr835p2AqAHeeKOvtr7dpZ3Xz7bpFQ7bIWtDgROYyW2
CMS97zLlTil/thAFWLd1WoTC1tHmMypgBzCNvrEB/Lip60Z+uRpZ46qNbg3rVpmS
MVmphHKq0qcRiWJ19avU+t+zmi33AVl0D35VfVz2k7Li+4Xx2jAjOs1fajfhq52M
12W69c72MwOwx01L0miqGIGnCWzXs28gT+dLOo7xfxLMvnvPp1DdMW7xwgIWEYJj
mbUK13LbHj+IcuJ1qR+YFXjrxdMF6+FKx99vvsW6vKUlMdp9QvPoFdL/Tg+070+c
DGeUwPM/NIl9Nrj9MCw7IVebBj5rMkrw6C7dft43wRDDWK2bn2o5MQDHRvG4Nmr5
m15FsCaPB4tzjlXjjiKCmEv9V6QX3uF+5r5MUHV/cmO8NDsmZVewXX6Ot0Xr/HBd
tk49tdD577f1txbqfG6J9G2zcuAaOopTyrTr8bjaH9pldFjNEEIXcrvxnD0m1If3
Mc0vtu6wfzEsj6CSGmVNAPa9ioxLpMgHppRDPzsl7GrVtapNcJv65ZgP21wS/o8l
EWyIg3IDNQv+vuJyHm03jpdSDF6nm39aH+0TQkYVOT7JM3lAPPgpNgcTMMqsX0O4
U5OWy0qmft610zITti3uuYL4kssMMBWtVbfvM1XvSC+J6pb4DTj8TMzi7CTvub+A
7C+Qkel8dGkj4FdtpMRBdYWahEJ5hF6oJg03HmnBqVkoapIb/lFZBpsYXi6SSjfv
pGVYpirEK4FEQpZDAsjR16q0xmwZymGLonqjhYjPuUbm5Qt+/Vpb9h4Pl8lLXjHu
A01XG3gN1U5FFqqoXkc7TyjJSgCJ56KowlijF+1JXk9/6GG14wAoF7Kj4dhkSkaw
m/FRiT1KG2ZzRHew+gA3VCu1QzV+kogtWwGmSMzie8dYATPEkthpliX6dFOJ1RJU
nuB2shHfQkSebHH5mwcyJYxZgWIwTPvLNnnmALQmG00udECIbMHFFjyeDQQLjIre
pREGsRVpg2LQ0Ph5wm3t+OZ9RuVhv8pimIbkARyJp5y+A11/O1rkb0Lu0vGmgh4M
NfqFAZxebfDqUxXPSDnTnf7b19yoVnyVrSHEsamm9Mx86cd8eDXztrjLpQ1SMYUJ
10W+AvfKVT75UB/kM8sYabbV1CSnrxRtAlAg2nrE01ITtquGDSdchAUJMtO7LzpI
E2RteyWkCiW4efuEx9Cdu3AwtHbsxXdditiRtsvvejFoLMg6n47eUBW7DN30tRoJ
z0AV+Pv1V0zcWpMOaTEAjZrM19rIY35jRwNqWkV6+xdR9Kf416bJYmp1XfIUvofX
QUFN8m/Va5OLOKZiUnPXbThgb2Niv7apNftKNU17YFqDdN36EqdUmvdB+9mz/pJD
nz0rNWW7hOvZjtj0xhgMb4kjTTjHE+Qu10qeODZn3VVl5tvbzaqeuG12zlJq6Aj/
2upQYzNx8DOlCrb6370uGFLSsq5QMNGahEpDoOkyiKdhLz6TMBqsV+NDSqzGmizi
ZmHvp0GgftwxfzOIgMEAeJ5Dcojhji4chpMlKBwxi3PRhzVLtYBpG5Ia6Zz42UEs
9RJC5Ncy5ohyVy4UhR6y2p2MPzvremFAo4BLqu5mQKfH+7HhbFd5KyP/9zoaDqMR
F8ErFXQQfCXH44V2fIzh9K4drpexrhAJN7Y9QLZjVAjOatk4rB536TmoKd+Sj2hR
4nBi2flSFXXa7BEVq+lcfft/8Ay2lcQZSGieav5DMRTAv2Xm+HzRxTp9OfKUDWWf
DOvAndFCbzNgaFDGC6JUof/Es7Ed0yADvEabwG+hRAzyo9CW7aKa2DpJzwgyov/v
UKVo2nTyX6b3ShOC/5YLv/A91en5zA/1DwBE6EbSdkdRSMQdugp2Ak1lI77et0aa
BAMHj07++DBymwHhWH8JbaNUTCNPvGb3RyqOf22Gy0kF+pXFuL+O4RK1PDtukAKI
aHuWFEeDW32Af3wYY3ujjbY0YTk084jvQwm+7itn3xoq9BjzAbSM9wYcaVNVAjwH
2KAgMcXG8zoSGJx34hSaeDywvcgwDPkmmwh9Pm8TPWE7RqwmESahWoZC4e970AfF
2dJCNBHAq/GfYU2wDHmCweuCN3AVrfl1ZCYrXEQ9WwKdcOhxKUGQQ4+6gJMNcuEr
dzm9VHSnDOM507pnhhrCLc/LomVLnondNKXuhiWmWwlWb4qvt3JjQPYAAyhTmPyX
QuwX4451rDkKXJFBjGjpUCC0tSk5ndCB4Es8cFgF9YiXrMJO/C2VGqEitMs90NsH
lPOxugORaU2pFUpHChgvIpKz1R7y4VFpG9uxs0bI8rODkCBdknB/UAWWkHYH6sAE
PjxrwvOa+PijB69jA0bAIavhvDtqGxTtVVBpedHSCoVBOJC9eFHXT/VkFKEsgdV1
2/8w6N+P2+B9OWmrvgwn9J2TzGjdzWbDHazMywBMf/NmQaOtTqm8pCqqkHF600iz
HbDPZMS6YKfqpOtMaK/Qw1yZv+bX4eOtnxi6SxZH8UQL7ZILIn8WEs9TANmyfQ+w
+9/E5Zt5PRpzIkaVng5MS2yQSee4Vqd20pQf58V/E4nDsRtoJImnsMZsn71y5yEN
dtr8E/ZEHQED+U5IP1hKmcKXKt/7IFXQHOetqP4SwgaG4jvTET2LFaZ0zQb9QNT0
Wctvilzg0jvz2LU/hdZTfCgv4Udp3lAnUvCR/6o8sPFujG8oU8mCR8Ib6+m7yBDF
ibN7hheION+qynGfKMqjxd0jI/jzeUJ4XYmO0TQIzQ6WaM+udUEMbOeRy2P8pAP5
IyFDaSaR4MByEcPcUEsZsBtCt5L33LLvX6DB8jPBQvBcLHv3uBImfldHsVveGOLc
3QhyT9p50VUeob3l4Qx4ldjZl5j2u6+BXqdHU/GCjuChNkQ1nZTO1Fy+2l0VwsqS
53zjSRUGCmWmqFz0iCvEvmJe8JpYxDYG7hkn7j4YvRwf4cEOlBleXCxdzatR3GQx
yfuxNx62vKZ5yDzidBllQwFFp5cbObXdpzEDMzahShPePTHk0ykN898LpLr2YljG
ubw+bsv88rCNGMi4KghEZbm508NmqkmpVN8P5mN2OStBb+7k35Z2WzYj1997n6WZ
S5IuZGMYpMGY7PH/NdM7cjAPTaZ6uPklMZglIiuaHGiwfa6FtJKeewEXjCInERIu
MVtyOnm5+8ZaFGKqEBnrLK6MvO8K2Od1bW0BB9yPrJCioZyeLPjEs+UzdrztUznG
trfssQg/DPZkE+olg9Q+LzaoK1CfTQaR2UHW7cEgsi9YMbshAKeeVkiNHc4rScX+
yVPPPtKDchtgMaa4LK0SDLz3cuIwB787jhOymYgU/CdNWXdyJMxtHMnPQ9Gbntjn
nVe+z2JDELtG2nVDlO7T8UcrBltQKEEYVJS5wlzOO3sdZFQCLDkCZINmTn8poeUq
Vw37qLFscxucH0oHgcqy0hlDnShB+FGgxMZYnFRUGR/WRYWHG4W0j0wklv1g8Ki9
hANnUeGUR18tb8OyHE0PxMPKRTfZ9xb3kcFjO8xEDAPzQB94b/UCO2aV5OSiqbBg
bpExw+B8104AlvoB1L5uA/eiwTeElg1Ww5giig1auJzlef/mjiBKnHTY5YxlJ1Rh
J3TZzef96UcbHA3bxHw7QJvhDzC1HG/RrjSPs1TjAOb9TG5t5iPK2JICD3/gX6xK
NUrirWgRdExWCwB0kDOU8nnMeePpdJ9g7bYzmWvo9trw7J59EC0OFVUYlMda6R9S
i5S1DW0D0tcDAlFU0EIBe6zobwpCrMDOMZtBW80WkL3aAKXPeb9Z4xWbszK7SqFt
4UCJuhGyDGX3jR2Pz+s7V25RiQt7C5jAeqAvlZ1KUKAqo+roJF0ffsdslHup1pkH
SofWbgNN+sp4cAtCd6kE5+WcGNU+5e+XRPpW/oVYRJ/ZDE2RHk3H9I9F+CbBY5vy
8uAQzraUdYt87DhwV7rjz6oJ2qXCLVEJ7Q8sQMl2b7E0YYs2+/HzxDJk374VdUPt
+q1kRFK+PGH51W0Biv0Uht9wd6wIeQ1n9gGzzFNzWgBMVD4Oe53+mgZTurMHJ6jf
F4OjV/Dmu/1yzWBVngZS2pSpovCrwzrfvc9n6Zy7iNDFlPTYAbz/JI2N9kaFyscP
Zd4tN0FOWd+lDL7b3hrZtbQ9dgw/1LXSwvTMSNTfoqwAgg6bqGrKxpurn/NGBEf6
Pn2lYZDg5PW5AwPaK/M6QzYHFVYHmMHpEJYvAN/va7zGiIvgzpC3VPJiAkqVnlnH
jNXs6l0S2FrUWe5OBdutTC4tF9VgAPeabPjMG6Om0gNWR6eM6QAerMAgeuFYunQT
wRxmt/a5S1PCGHLRTxfAYN3t9rhoJsxa0vtwqlal+n6yMY2RTYopS0VUxXQcvO2C
28+zI8egtz9XZXuN+1KorQO0knqRxBgEyra7STv1Iz4ninOPguC+b7lWBlLwXOMX
/r6MMyv7iCtUVlYZloQoX8F20RR76rjtcbgdP5XzWqourAAnAKUOVyo548Zubgdv
1heXmzVzrAUEAbIoXCcqpH8esm1kscSLN8DwqFdBIohizLhBth+wcEReWbNGFSH6
30l9Affcd8VMB3xJbKd/++gromDoge5RqGFZvhfKtD9bInNU1a+T6f36HtJy04Rw
Bta/iWIPqBSZoSzJ5pyy7lDWZq0Ik7S0Uvmqx1URkWyIl535rdAvjJzEtAvT8YdD
NouQD8U/1r/zlMTSYC59lvrOzzmLChfIftm+I7LUtpF3oHkUI5hmajmTSEY8TTcb
XHyvazZchjTp0FomeZ1uAMUwp32sLuw9k5lguFOjsxTcK0r9Ojcz/oZl2CdpVMPU
Yj6qUMrAAFoKd92vYCFzRsYutSi9MkuuT1q4AjE+sC3td9AechiijptTCaRJXd63
JIVzAGYcGQzpVFzgMq/0LGpyJO19Sg0ViozQWfc1cJ5/ZFxMdrgFvT5wPs0VULDA
zBVqcCzj3TXC/lGDDL2Ksi51pk9ONN3wVdZJ/Tg8vz4dstMHRBhRiG/xbV25gako
DxF36s/A2laylPPZxTjGv0OmCEUVdHHCINiqIHnwoaJbGfbj9Cclq9AChFi9Ts9E
xbpjyOrppx56m9n07V52lAr+GwLgFQV0dVhMqbOcLLdVTs542FQ6XaVhmLtQC1z2
VgVRNDRAj8M0r8b+X+5cMccsaWu4377rhFSoQb8DRVGjOD6rO2WLmD96uwhuDOtp
BwG914Yxz0KgEnTo8MkZQ0gEEPXOR9mVzjwwQL5v/f+JdYqLfH1eXmqCB3a4wOXE
zvqRkdPDERAsxT0ZzKC3J98Ppu/X4/Er+BwIoUo5MGAp3yhNkNXjNQ4RFld6lq0j
s0enp0rP0l2lu0O7SsLoeBJ0XVJi7Z6uxjdoUQxy+BV5OilK7CCXUT712mHU2OK3
EfXnMy9SjfS87AakbJBs7UrftnXwh2ZaOj+QFmzWUHh3UbhGQ7u2ebjDAgPQwmh+
kYI6rGwlTww4c1PSOL0loHbL9ykoYjh1lV8pii8tZfg2YK+Ms1CoyhpSsSh9OS3c
YkubWWRspm/auhiSgZCqb44JlJZYRn6LFgxHTZXADnYWC3/+TaU6mFUazrwqgvqp
8cCVmzONkRql0GHEn3P+DNJJWYFfH/DYwu5WIFsNdhnaxCKDxk0ub5eXAF5fIrei
Q3IiqkGRpgQaqhgfqY+3pYSqVe7Nuv4t9803wOWrDFd9tu+Udl8vRfPqpKkwjkiu
sJ3hczIAbf4dP3uBOSPBL4THfq+Lpq2Qwt1MZeackr2hUMGSkiUJDbs0iBejUXQK
DBkWD/BAnfwB4rskzKS5vWmnSGnDrTMJfiBqAOLLbGg9j/NCDfwhmNprwRbh4O/n
is4OtVPRZvWf0MXFwhtYu46NEJJK363e2yVzRN4Ze0jQ9+Tp79YH0S32DyyjhsAl
VPQkd2serUiTo0C3v2GN31gJN3XRktmVuiHDjBX1f0FkX0GYUNkY167eYoCJlFYe
lExfFwbqLbb9TeA9nYs2TbxftBFf9b9NTFzjgaFvzBy9/ILcGCB0YGHPlScSEdvn
UqcKrAQviKrr6gcA1I/WtSltTRRa1lavO67jEudzLhBkAlV/aHv/G6A/1Kym7Jgb
zbMKAo83sZqEh1iyV+tVK7jOYg72bX8n8bYTR2d5c2TB7j1NbYaw9iKa5ZZK2h+j
VW6a9v8ftIoiA2jSBP+cXhGZ9Gck4XZq17/2Ddv4V7c2Itk9hjdZgLd6hQKnHYyf
/8DfD/26jG1+GwRKQ01nI1HA9KDB3r5VXdkJXkDNU6W5K3FgGFKnlO9Y2n2+cwhS
HxYumfGYiAZUSE4qLz0wxGC47FOq6LIC8HZmFSly8009EJm5AAslstlEXY3xkBzo
k9sXy810Qb9MvM/ElHLcjOK4+claCGygkUYlyAAlSoo7WpSoqy04PdEWTXZJ3NrM
n3f4nzWa0k8dL9zlGzCnKjZg448vBfWZB0nr+BTEQ3MpXmJAJEbvrQk/jL3vBMgV
4tq8+RyA82cmBzW00Csju9k58wMRdNNY5eKeDEnxPgN+aVvERwYOTqnWszCnjTEG
pZla14VWlbXdSLi+v7n5N2mF7tq2sjXgRjDlBVmsWR7BsKoRNh6wwIVchAL7UEtE
NsdF46QLhaeWIYfbrd21tIKDdOPzjHzi6IrpNEyjoXl56JgaAW/V5FsTA+/DbaqX
V62GXBEu9dyj2h10mRM2P+BN9NGT7TQ3i7bqBejjwcP1udSSJp+Wrofwe9u7R3QD
ozCUbGdu2eNo7if6MKYnwsTvHYH1ATmBmdjynYFSb3O7jcDNJQlmtVO/XFM6Flpr
6pk4PCil/68jD0eRmeMNjQcPy2RNrh+/HhLGXzN4fyNKFB7Ramq7M1KkE3TbTy9o
RrhjJJr/4hXJuracv3NsIr56wFEFB4sNKOz2aDlL9lWtRvg5x41T5GXZ/GTPInVI
JrwIjGCXWPrwam7i46cJCdsP6mfDtVE49LeVAIzHQro+nS9gEY5gsRNcLmcUpZdr
+JggMP84U/tFJVBcgcSxZB7GqPngy8Y8sWH5zOZoOrRi5uy3Hq0bdJy9yMBwY1ok
PhGC4n9QNYC5H6OWrut3VoI2xzu4dxilbL6ENLcazfOmqSROI8OdSsQA9+Wn3nBX
BcniKWtLYfB/8sNEQP7ab8QaNBLvgHzpGN5t5PYcgiHm2bx1njkTJFIHM8uzdrC5
9iDI6ZHiqdPxR/knmduIHT/ThDw2oLizObtV8xFaAMuUCVmtPbr6R5eVdSFQRgTb
X30oXYtpaP67AnyPNuJgYLfcDM4VQB3JfHCdyZuTd07pX4fw3LMrLOS6SMVJpaOk
KyGcvymTxK+VVj7NAyXTvmjBLpZ7qxFnSsDxJpO4WiREkOHSnDpTWJc9p2T22nTq
WFiDLlZ/tCBkFxrATuk2oQONv+6lEKYI+owzSGeRSsDjUrwCcUAHExOBwwiJRv3r
TLAeNM788QlBuv5EboH4u4zFg/ehp0zgF11dEkXzX59ZO6Rgh24cIcgaavulmhNW
41Ks/aLguad2VCHvmLVNSWj7YXnlkg2BnHrUKNTxLmo6meWHBCDiEoR1n3lRvwLo
cH3DV0ppLXITkHZhHEnpLc8DjlLjZjOSi7MT8dQfWqA79XsjxmXJB+2DARaCkpSq
FjQDuOQJ8I1t6JfuyEXcf3bWv0TsSUxZjGF9p6GzSY+9y2iTzCeAw1TVBp9f7I14
jS7lI41PjPmPA11b10hNaBtI3sTItAuEWgfQmtuoJBzz3Xs9HVjlICtSOykY8DKq
q4fTNrnvfw+dbOpK+DDKq0SVc24WPsXnZoHv9GSEfIQ/wLWVRmzio6Hb3b14Wi18
5CKwKBT5+9GSLxxhe/+0DKN0PKsFEgwfuCBdizwPuHghne0jwB5lQcLbntiBCyhW
B2Kz5G5d+gGePDGNVFUfReZ48WwLLW1l7I5sCRU+BqvvBY8f6F1y6WodGENQkJ+p
vym68Jn703YdRWlOCWG9rqkCSUpUxmgO34678uwi+E5ga80N2/NZkiqj2zkCJXaj
07Kdi90Amg7HkI8qDeibVeg5x4ZzT8oLRWypzRGfUg0TJJAG3k4vdo4v1jFBB9t1
wkHc2FdEyZOr6UYP2t5WhWYQ6AKUiUgZHjC85bUs1U51w0uIIkBuk8Tv639AW4Cm
jX7nBvGU7D7Rv3+AOHFNPp/wLvCIgM7E2XnQVt7s5g2XxwRY2v+NOrqbdibW9d8p
osWiCWCL1gZaZ648fPElTSlKCFsU6Athpg9ow9W+8W94FK8vzcMTtJC+7Ba+nqV2
ioVfKwIJJQNLQ1NXVjgxYMOFh0HzRPz/A82x0AHLZ2+TSP28TUh+NsK6RtaOcY+q
AZJDBWblmToYM+GzdTooja+6USFIbN5hGg0hUmm0XNhOEd4RLH1bxVWEZDDIcTyn
iXTlHp4X2QZ1+EXS199R2W6Wu/7Axa/bUyNhFd5G5bNHZVelqdyGmUr6YBA4IiJ6
F7+9BBdGjsDRYzmO46Ky603NY9j0mmxm4cpCJS09Xw9MjwGMIBC+XChbE3WZRtxW
k9TlwQqhrlmZizo36W5RwcAF/U1jniQxhMDMhQ6qYs+JIokaTldVnrGDpNlPMcEj
uimrQzi7rdRBN9iFqLyfjX8VB1nxkjdEYqqjbgCnis7yKUGxCt2WWy/OoZo49Rkd
6tD3pWgCvI7dP1zwo/Oc/dZ/U7Svn9uxA3FDiS2HZRHSAQtH7S3GzQLIWOIKBBn4
ZPjqqGct8Ke+55Z4VjWuvpw1iDodT5AEADZx9IVclkCn79KrA22YgyS76hMoEnxE
tgsdLgk28xqdgTTvX4BJumYmM85LhBdJ/P0ahgjN9ptCX+ooHlWClWQiK+EzNE6l
nOH6DSu8iJruAXAPyTX6QXouc2kwJ9O0bYHrQGdQ6J69yapNEtSKNqxQuMUiH5sz
QImsn62wkKgGmN1JNO7kMzR7AWwEFblKbQ09orV60EDFalZZu8v2vLfYQTqJJNgF
dE+H3RhxKDiZbZX2HWSkvyIGYHBgW7YC955kuL6/oLW+xGOn7p6PeTArJjf3qs8x
/DjjzImk3XgkNRYzyIAfNs58YoxaRtlkO/G8qBIQGU75BuASxJIy9w5wGk6OCNj7
Ff34C5S+6cJ52bhUoawgmvYEgccv0E4kyJR1+Bnsadzm3IymTOzpZPtG7ilWw8Ta
+4Zuk0Gfxsm93El4Y/fJo8QaN42nkLx1f8fCqlfHyjR/PksZCw7jW3rlyEbZy+my
iQw332a167Pz6kOsCrkiefTOOdf6FcAxpGjQ5mHSZfeZkna1CK6kRefnhTl4YcM5
IkR+Ra9spJay+bzHocN9LsC0ZpvAtpkdOrFVWINKiy5zSCD+BcI66R2WN3cmNNQ1
3qNq27PU1EDN7JkDqDCkcOQNtiHbpV1U9J6cplH16W8lMOIzRhGyO2SYfyyohBg+
2poZDz9nxfEVr2UOBnthrrX/Hi7WUs4cNw25Rfur0PKyNkSZ/tnzR80XN3sjoAFA
HeCAqEoKjY6b6wRPzCJnjhtR2G42l/71OGNZ2qfpfsk9Edr97oWGVDJALQylG2Ns
Wl89PBLqnPBVHdc9HFuNxrLCgL2fJN7FPountEJxNbK0vjEldQbD4WG5pWjuyYd2
r1CgIJdqR3q9whd8VC3Cnkudu95EwuYdbAxOjhSBzUJ/iqWoauZfpNRMl/nOBsWU
3+Q/8yIeLta3eQKim4uemAKrVImExD6mRssnXVCHsBrxEo685A33oE0nQ93OskTd
n89BGqaMCJEmyIX/y1dbnX2cifJbi5XhoFimeEnQB+uGCPMcZv3+RxbKYe0Vd0XS
51tRfRxBIJ9dsr2KdNkBPgJgue0apD+avSqf6IOdhagolhvZ6ZhKiiLJZJQR1VQR
IKrGJ0tHjoJ2unMQ6KSodUZVQNLpf5NpWTfzYTEv165BJSVyP2M2JCUCS8jEtAsE
JMbqAsPQqjiNXUgeYxFPSGvDg+bt2RmjygTscIodhp6E+BXXsKNH5lfLNiyt0eao
J79Jjl98p0YvTPqZoJ7tdxmhqj3LR46BKYxgVg7dOUCVDrtS4E5smMH+oVSgFTB1
lYlxnSb3X+ETO8wNwrcxE4Y2mxFzDR//QvyFtVKY38ZSlc+9T9mTsn/SUlmdQgku
E+wddj7Jly37hN5RQQfBuH7JzLwE0yG7QTE1eUvC500hf+mFR0Zv5QX7wgr+0Cqx
zsLGYeu1ADuNFqq2XIMmA8jfkPGHjsxKE4noWIg3Gp0HSCdi7aazje5dyV9Pkecq
v5lWM+BWwYCd7AdJZCLuW4j/7dUbq1C232FwQI7LmEHv+UoCvwcKI+0mV+ia6njU
7YwzU4Xq8uRLKzp7JKfqFXkW9gVXYS9PQie/ymTM0fr7Frs8tXLe3EkZpDYBG7hb
kkDFmGh89StCywdOo/WoSwPIShL571465NkdYS9qJedpGDKCzcq2XJE2Wd/h2+/A
0nKIFdkUFkEbHdx/E4vVHoLRtr/WVRtmRafoi/FcLdwoPJWbJbmymERLiQ1En5gg
qllVk3OneigjdmZlySdOIkdTJU5i4yR7ltAtdA1o+1rwsoXO3a++/I0stqnZajXp
evrDjhcVM1DtgeOzRtF9be8yvBsicnql9hBNw42w+jFanSedwXaW51MTax2hgByP
n9To/dDaCNKvRIx2rICcJ6lQX3C6lpURr3iSfeAGf7rR5rNGgqU5Xuvoz5RAvd0S
6r6fbgAdc36eab2/CzXzJJkUszl5t/K2gu501D77voEzZTC70ubM7Gds6RUsg7+o
MQmK042sFT7m4ppePLTnvOH/PqrD8s+UU50GWwvV8/mibkt310DF4+IHftal7+dK
G42++l7Mh0sy8BpSArW+Ta4aS92NwE2DaDcG82d1uXPo6aQpPiWIWMOBiuWlxzEX
aQ/IhqaLYgPHOTbCjjEJdCTOjb0VsW2cILThjA4xHKCKQm/+S6cxfJDM+jBRTYw/
SRGi4AL+URqsdKvzbFeKgi1ofzGG6V0GUgk45xPPCeA2Dw1remYummfJ7Lwk4SNl
HEeQfsfSVjhhN+B07uEI3J8tCJaaLrzPnoiXRdqtnE5h6EqCpfrDAOloyXRqycK5
gDTPfCQbDCkUrb+BjH7eS841QQqZ8HyB398mLojxlWt+LRpMtRHUNohN12AYDTD0
8RH5YWn+NXeq2sARZ84Lag5LHe40S9X3ARkI1EnK3jlRDFzYd7MQJavqvlMQ0eRt
IBGhOa4do+hOY0K9lKSM6z8eRIotFXXHega61fqZ4tKU2jwMf3fuwx9VleiKxmoJ
FhXeYqqYbIJ2NW+iQbYmeh4mh2jXOt6KVT4D45Q2COGqOkau864D7BwMaK55IqmV
vtkvUPZ2WD3FGjD9SovIh4/KT6zoA9XWpLl1E77C9oTpO1uT2DUKwRSdossbOAut
6P1w5MyXh5CaKwfginTCrolAU2ZhvNKZOnz1Q+DcDVYgEBgy1hRG8+G5jImMvA5m
pqubOADTKXcLMoXrZUfF0TcOZLYQdnpEtXw3so/jkYWLt9uqm3w/jdtfMDFlT8BP
8g9AJHVHO3yqc2qGU+1HjYHsfMp57WzbuSoQwDNm3gQm4/Ml90lY+chZV01Sguy+
V/29evJA7HCwHELdTxLP85VAcefdC401OzGAPn+dbUjKDBVgSf8RaHg5tBu5doJw
3XwyiOEBv1q6Uts/9xZdga9cJmj33Q9sDFAKEoWoP14/V7aX1KRGZSNZ5SFE5iWC
Loz1mnvgzmF9v1K0F0P9mx78fW+GrSimJWIUdOWDz5s0WzsCGqrYNxYOjhgYufrz
vzZ7qHORAfh5F/1HJUdO8BJzNDdPby9IYw9mEaG16qK71ha+jTMnswx648LjpmGw
xwTzKpOPQoNbwGRwL66q5dALgKKMLoMnRwaHBG9jPVmbPztISrJ0VLKrVn6yTgOu
IEkAcWE1WNrlYCPOevE+F+TuJKE8PLrT1jg7hkg3GR6iFJ0yymNPUgwaq/nFSONy
cdU7jZrhoWNmHmULDVumOdim/O0fRQGyrRHJqzDsThM4os30nueRhWQp6O8DCeru
W0UtSi25HRsmh7Ra7d9RTnaswXwqDIQn+yKVeFts+Ni5m3jrqjsodLg+oejLC3Km
ees27F/hCVWf4WSy6CAgqleVMwITbZfwamN9/l8HVbgDGo/tq63DFZaEHYkVtTkB
w4iH3QvbcQDx3W13QKBaUza8lFBTSQZE/5ctDIDwiDaJLzAO3whCqiBqNs68qIhX
sZuvoFMnz3uYC+rIovlw2GAFA1tjf+Do5OAYtbnAUQytmd69Q/n2BuXcH2jZvkwa
TuB0BCjxg/X1x7NHUJZz7y1GLmYWB1cyyXbEL5yw6GxU1ANAaaJDY5G39hQnNa0z
cNOYEVRbsKvPCk55O/Y4q2R9wlWuRuqCsLA/g1i7FpV/kT7M3+GN/i6lKfkHLc2p
2JvV4D8TvbpsoyoQMIhHc25KR5JzqtT/r5cDPouPLJQ1Bh+UIXEruu69gwhoDChJ
+BKXnQW28ypJqPJ+FfKDT0bOeuGam6KQEiAzN/GyaH0v8GAzBldPtGcgv5Q7kMx0
470vBPbJ4V+ZZBgnwvByWjf6uYkKr6D/ibLtEmL3ANPWiWpJPUKW5q7cciF/aPwC
St7rF/aiSWqxvDtAE2C7tWOtNv8n4D1pisCqF9iPTkuLkoZ85ZgFOdoKBIm6vbvK
vO/5mbDBhk/XfsXcyF7yR/0AJqlDX4ADnUSid197OpS9oWJzBNnBTLL8zKa37zz+
UCFgqVNNZ90vf0eWlcOB4IZqHW+Jwy9/z4oXYqOR7ifnJpw2x9V48leURvLxocwq
SQBozqBPkC9Vl8s9vyqJ18amB2Y8+7//Ypk6mzufg7bPJ4St3GimL9F1clMwxW32
D/FLYC2zBx0bBYpVLiJzSRVAh5n1DhrUY0i61cOLxEjTLZlVc2FfXbgyio2IY0i1
o+xnlZ/hceWjLLuToeb8MtOZOg0m7vP1Xp9qfm5fuAVqA2277HGiCEbcN9My3KtY
eIVgomUR8Tr0fKGXJHph/BNOswNjkyf/pKp4FQOouWvEGyn8XEC65J41OAnNhZZC
kVBf0V5bE/2TvZrGvWqwe7cBQEZ5Vm9SMUtuiv6IXAPJkSEOS7+CUPMZStGW0ZJ9
WgVcSjKoy/x0xeSn4dHsveNMvFZZVa9Im+w7P/qOEZHXHpr7YBmOKav/knA9+Ifv
TSjNOGd362FT3iZjcvKLAf6kU+FpELsGRzHYeLQYvIT5vGxvCtrkHO5qZ6lcLq1m
ONnwDtinOV4IDdFm+WirT5fEm3lm3LCanOIlsSv0CtoMbqMrfFLuOEETZqMHwhAm
Lj4LqcnQLCbgI8mNBlrswqi0vO9KzkOtJzIpKThfLOsisFmNtQNTYJOtzBGzn3A6
Uamrv457VqYp+4snNcGrDy4GKgHj8I2JSjRnNhSwYKuPihR2P8S+hjyxVpbQXCpe
y82lMlZ4VgG2WcWpdxDJALg0v/zzcV84Pq6Z4K98WGFbB8lYkcX0Rim9es4Rj1aS
szdf9d8g3FcfzgdZRSKewz3Uul3klH+MFPGhj+YfNxCbtJiVPLeyFeiPpbD9/zcW
dgIBxoGuWlcd0ELM53+BLu/7O/3ByYKYXyBqvfDGu2q/jP6S6SVt6gKAiSYsi1lR
/0KO0hEdAqmVGFjmgaB3KnvD2yhn3lmXddqw59mQfYz/+a3kh4MRirjjF+jF5rn/
HHuXzb92/ZfOpOuQecmD35eDBHX3KCGzXr+wNOv7cMelU83THI4FpfuZxC3KBSHt
rNRHrhIz7oKAMql70n3liYYmWeZfN1YX+MUWxya7QrJ6PRou9aI7sJAICqL5sRp8
zumI8aTzOnOPO12ltK11cEHM1x37AMuGhkIodOXzAo21ALmVfAeVicA+RUc3OvQ+
TXul3XA07miWdHGcXlrW3qhUXYhZSckb0+GXdB+tJwUjOLq4RoPTjB9MmXieCYqB
q/wPw7CDXA0Pur9Zhcw1NhYW3pdEfaSMnvyslJsOdM4wf/DadXaXDG6nguYSq6e2
D9WUwNxXsDkADOLmotam09d+2mzO0P7dfwvFdWUkpu4sPo5uTP5DuPh2RV5mOmXo
1VFENWpIvoXzMJ2qG+PIPzRNxtvUOeG70ZHG+UbmYpoRkeDwHHz907WYQsuwQjlY
ti0Y9EbsxJEZptVT8ws40My6T8+WIXaryfmTA4p1Q7KU5npAGDLokUGEF2rRhlsi
wEByVL/tLeCOIkTT/5yVCAop+u2goExA4ezuTp9mY++1thbOtbHG7oSHbNQ2+TQq
rYafE54bFRbdwTf6aci8PIbu65BtTl+b0JSmHC1n5VtCzYiuK3dqgerzGfyMFsh5
l+y0qjbOuzTsmZWv05Fd5FbZv5rGuX4d8KQZZyvLppv36mzzB6yNtGKwBplXCGTk
G3VXWwxvOHBggAjYKWbKv67P60AoVsI28TdwpvSFtTaTI3NuSzzGgBWR4vHa3N/e
nqTG62LDbvUWvVAmiz3ZXHRV/0wJZ+G7CcwVTmQfe0jUu/+nqDRJg2wjfhkxmywL
noBmnyQqraCpGETCXXBLpoOU30LYHhMaPHA+/rtXIimTxgp0WJFYB4yPXd7LjKrJ
97ndVJVDGeAfwvfHqN7ybFyQpoQlOdosni2N5R68WZb7KvpgAjCk69kyqaVkwCM9
5LAuUWRt1ko/ni6wPLqBEnuq9HEoPfNcWAQfQb/dtu6y1XYL+sI1KcldVQud3+lP
gPbFUisLShudvBJL/OhfYTNc3S5HZr4cQhXs6x1o80FI+zXk458I4k5XxthWOY24
8I8dNL4FzVIpqSur1Q+lNWGMMdYyaKy/RdL/0RnbaBEHT8Lj3Ga81zCTsEMrNq8f
4C/njgGJeJzuifu4z22CyUFOsq/yoBt26TTzOOhnYZFlSPVMj4hwTgC3frCfyTCD
lTkUbOqSY5ulgarffQfk+qku4W/9YqwU1fjgS2+caeXKQ/+DaImtfRKm6JEOGwsw
er0F44PTP8NnZJ0CQvvaRH858sOXUJozLR28Y4NqtkM3t08EwO8XlOh/He0ME9RU
3Vnpe3X8tEAebh4c2dBmYPkRoeZODzVmwQFHNdtrWjbskroWTQFRosgZWCfh3ipS
GOwwWJbgoy5ApCf7E7+B2wfVeJxCpyhV21wrT+IsypaYG72VbiuGQDAagiNRDOS6
MfcVqPxaT0u+iOh1TEgOby/MbmppEhBzJkzYZ2r5rP9C1xn+o9nH3WMTzfay7O0S
hXiWxC6TV4BeSszQACEKf+Ktn08j4UQ5GQMkopX47da1ZUJoAH+kDLWz10FGfx5F
oYK6G5X28AKTLQ7aGQ3xnePbmOsQ8evEepCIgEWs/9DkfvrssrQeAhp7HqUKRDMR
uQOHCgEWlxt6ePqzLyv01WH7Iej4QgWlu8grOwR9+AUXxfgj/HSdnACL4K8jInTv
4o9xoip765s4IQw5ciYzM8ClZPgG9dcveefjlozjJAbvRDCKfa7URsmrLgzMKTZK
lfAVFrhyEtUWvTU72ZDLyAbkJCGFlDySmCjIMAJqXpr82RP+RWpRKsr6TJcAWkbE
or1N/M9SHwAhVB3GY3QmFgB2Hz0DUKs2ACsR5kgn7wu6Gwk4/+AzSvF7hstgBHsX
ECvuri5RtKMKYU1JWufAOrUb4c6Lz4giUuk+Lz0qqtvkdCjF9WO2WwxptetA9aAo
HEtwtpRO/JWrH3IJPKGNHmwRuGr8WxgQjCohpP/SFja2ixG+NxRCrfsBWDFLoLZj
QD1auee79zsaZ4UJVkaFV91NUh/DMJjbquKboWMyXvz/mVZ1TocfHhf2TQMUx/jj
CpGjEPOjrTg6Yk95NZ7ZW+c/4cRl8eUYK+C6ckZFevCMyuZlW4/sqpw2/+Fzq7K7
+3Dq0iy9aAwwvIxTglcNftMt4DK4IQN4OWq88UJ/6iKV9+rcFUdi1ltxCHKWMwzk
03ZNRyr7fsXO91ZbS7dTqYsQGBKZARTFnZ/6YhkV+gbj0kFJurMy4r0kUgv5GiuB
p0cqSAwe5+W8Gd1uHjM2/uboj7afk7eM79hgIGADfLhobQiOoCyF/skujP650Cwa
OeSt0r37CSIeqCuGvG8lWdiNmzcyBukst/tIyC3cSkaVdNIrciwP6b8qZeS3Zsp5
DxfCIfce4BNmhKRdiBGfaKgMh9zsDzumwXcd8wo5/cd/OblDzDAdyGSWTAHKOXzE
u1TWSq3xldIiYYdDu+88yziB7J1HPakvGIHQCtBB6HfkMi59uOFFzGfIhr6ZxLAk
fbe6AyFLh6xxr1nAwG7cJL8mHyXdKtlgklgTZahCjoKAwCfi0hnUkpJdHogxXar8
MjfPX2kAKdyiAabypGa5UEfg9F7dthqXtRTKpgbWvbx4WulF1XdFOA3fRNu6B6y4
UElkKezIWWkQc6L0vhug66cm8RcOf1jDDOTULlic6iferDV5y9SG0ZMJW0OyUG4S
VnxfvV+gGCXqEjqVlbFdZb7yUeMxqvscK7KFYGutysA2BRXrYPWkoF3myCkB90kt
Ohygyw2X5zDkfpL0GaRKBLVydqcIxJlDHfHnTVlWlUMzfnfo2I61jFml0dFGZmwn
WFwqBiy0DEiGGMVEh5yAJpQgxmmiw+Xub0i4nGJ0FzeYCqiOO7QeUodNkv0Q1prj
E9vXP1kDXWZncctqIz3TUcw/QSA/YlGTVLfIsn+hw/VvH1mKEyhptHbWMNxrXuYD
il/l/3KPuKW12UlDDzMDql4WNPuTCSM3OpvXPFtKKpyzgJxwKJUYGzr4BD/1BrHl
cg1NnTF16gcngpI8IOi5v4nLMpCneSkTVJW4ntu4Q5EGFmU9OqQOJweM2RydBfFr
IzG+BcSW0FA/y7KIWsePUyGmmkzlZOcvIHL+jxu67wvf5i40s+k6iHMzEEyETcET
PYGtE5UYg128DATonJ/GEPm6y6Mjj1YiQ9I3Qsb7zB68FD8xaJO1kO2YYNnJZLcW
9HSL4lCZ8qI/xb6vAuDypTHMtpOcuD31bg0dfD1zEj3xAEuYY9a1Wx6YM19aYfi8
T+xbrFuaCKx4CnZOL2U+jpu/gnut8wAH8sTCPbX/kU0XmMbQvnrufFFT1JyUiYlS
jWLc0vnE6J2BwiE2FyQdkAluyIT5e5pcP+1tA3Ke6BrtTIIt4EY+2vJ60ygdBCwn
jLXruG3CRUMq+BST4tWQznwrMvLcTSBTdrnciRUQXBNfHx3G4QiHNAGKmqo366JM
isMc2uPwzQPddk/kNOWurVRVsAfnvVt7PUiwqV6zbBJwnj7efVHFnQ1fogoPF8Bb
Eo6RmsROwWxU071292KIYLJ6nmPCDtED9VwvXdN+Bf3jtJ5jhARjAtfu+0EDTO1K
RyOs8hLeg1CxLB1VZWeeVH4jsv79v2T86kQH+8GV2N6mtpsNxhfX8hJdVnHqs825
5QES66tf7YzNs+9fcysHE14B87Bh4ZsfqyarPrL2ZWwMI2Pp7U7BdpI9wILwpeNe
vNcEmSd6OKr8Dg6RJiavBw9Z+RTUxtmhlsCU6nzTgSRCydY1FdtlofJzxdJP/BeO
6P6zgz/X0s+zDEbsRlRvzhi3MUFUEfoTCnUDRZ8or3ak+9ZJpl3+xsci85+k0wXm
QviaBlQau0icmqX/W5Euk4yqTrWPc0EI8vWLcKSwWzWKYZUJxhLwuz2x1w/4I3d0
kv88VeoSlrj2Z6yBaC0Uxt9nNIw1i7k2wq3qEQurrDu0WPuGlAgFrKP1+vTCwQx4
dLmOwuBbG+VUGYJFXZXqOn2lbBi85FB0PLLHnXLrh7lfTtZbbArdGrCtXEGLuYSC
sSoyWE43Y02QAeNImCrKGF+1YjB3w1FGcgsDdJPaKPYDc1EV0RNZNxCRiQYMdtH/
8LElWVrhYDYJ9WHPGJF1ve/MmVewEmRShRiH7oC6K9QM3UaQJeC9cFLamqNA1zZf
eDsp2XgNTsUsK58HuYiZh/ye/dEt0zvRSaBJS071CkvrLo3iGVOgYXdejt4kjnWV
OEvpWbSGoU+IhQwayyWKT9wk3nUI4Wk81jEFwHgKReIcnja5n5EaYWiXoF2LXSpp
jgv/vL3MNOnunRse2NucyplJCwp3LA/PCnzRiWYvQr6bU48yJwkeuH7VDpnt5skw
A1PmBKnvIAzRFGPvJCcDlVkCrNxpegi7d9QmcBXd4yqc0LH/nqXsn20Pi1Gmt/rm
WG8Oxk31cp7YjF2egCwm0mPbcNAQZYl2DPtH7bnA3RWPv5VRWhKDZiX1NgR39LfM
UvDiN8L6XnqbJApWsoru9opuxerjJb4rFxM62k5BW1z0+d0R7Jj87E6auGfpTHha
PS+oZNgf2JQi5lHYDyCQ3ineovA42NADrM8C7i1ADnwag0+/Twu0yiSXhc9YzTt8
ZF8ku/J63OLNYSgrPQo+PL1ZUYmtUybmZhveiBbl8O6NPfM5n31h1kVnuiJ/QULA
X+ePSkVNSOjVY3WaTtULMEQ4xJsGseuB+wobx10eL+TvfxbO9TrSQLZQiXB2IO2U
GDOYPk6xMFGi5aPa3hnPNNSiYLqdCOq/Ye08xVSDJC+JKhQ2NxVZrV4oZUrw7aWs
dV/fiCzvsYGCrRU9o3K9Ayq76Slvel86WyUclBvE18H1EfI5NUWp6SmJdb+n+yML
6MQadsvr7fWCeCiIHUfNIFUzo6N9FpO1Pt7I6dRVHF4gwhVU8WYGK31iQHg4vfLM
r34Bi0aet/Pgy6QWng3L2SMYSoUiMTzE5X1/n1KwSdFuD/AMyNRhN1lyqc8jSwLp
6jDP4UlqH9Tkmbilz8Mw65SluyxVYhbg+suOy3JO+40vGFd3FOzzC6sgW18v12jZ
3ZvpqRsglIYgXWgoMgaIwmC68f8izkEZiQSuFwr+Xpa4Hf9Tp1RwJRO6Ui9t4LSq
thJ2Ar3skphlSlb51iksjQRMYfitP3bHQ6VKHnsNXBeVullicmZrE3CZ31hJjhNZ
yLrrLie0vNBBGaoC7Br8/0m8+NFt4kh68ZXWM9ehKLD/dtD3efraAfl5OCDMRdFJ
klWDMkJIuEfM71SwSEzG3A3Lfnf1HVo7SiYl8Vwt1ZFg9G+qYnbQPhAGf7RDNeq9
gS6BEA+vZQje3T7JDKvsUCXnTbKb7PMsNacaD6jMN5R4sMY+2bo18cEBDSeMnHCE
7Hu617zSH0dLOogDn/xksM/WamZYxmzT/7GPteDtEjSkDE75SHwjI7njTJPurwPn
g82piAOeGvjIO6pZDYnmDRpMSZRyvBTbp0b1Ze6stzLOF4AstXR42hlkHGSHAr+r
IjxpVwYkWS+TY2B41dnWb2Cua+kTKu8SvbRJbj/Bx5Ht8Y5NRDoC+OTlE50Pphtd
dQoqfEiwZ0trReKayESme+FSYYyBw0kBJmEoPepxSuj2qjlUwT2DDChEidMR75JQ
jojLfCK02EIyi3lWnfc3zp3Banq7gj1dISPZh19qHOzDca1eYDKzEVPRMRylFozw
1KuLgQaWYFXZt9Ti1SRuEkvZ5ktnhLJQafN4CvFLxuVWw2Rf+rcirWfzRnSydZEd
PkhkwCPxh31k3SwYrg6GIAiRDE91nYmy7uuw+2AjM/raJxP488Yd5B0hvi3i73tR
E9+u9eKWrfowPnVRhC23SP0xWrayv9CkXEWgSvzZeGM1GaLhIY49kcud84Gxw0th
EoFB+LRFTS2Ag0/bI4w2VIjp5ovFx+J0cIHbogOHqcpnibP+uoH6u/h0bxZC0IKQ
vuIyHX3xZ/3awIBPr0SWbfASS44NHQ7QV9p2VJyDYBFRetfLAPReuULirKqe7WY5
O5EZeOEVwlNKb5FMSCQcVj4lrFPXVP6wo07YMz7hHZakxtRqJZM07gZg6ujbpbu/
62K3BP7B4QB/ThP8OVqeaiZyn0hNamlX6kLSfsC6DQO3+qHy1JrcVhUvdwylYc4C
GFEBYPzKdnNvD039ENJ3SfcWQf47FwQ0UJ/sT9ZIVw7QctdMOlU/VPoFuTQVQSwX
Ilk0qEb6kchoDwCoiIHLKv76Iz0JzIZ4A0rzf5mZtRAnzaxa+XY7tB23W9iY+Oe6
A4f34eCenNr1KGwCn82njsuXidxBJOiiIxC0Oei4OdQlD1rnbch5YpaBz5puyUeF
ly+l+4vNVzhqBpviZ+ffc+EBSptMMR6M/XfnpogC+DQNj8ASOqMZbye5G6Eonzvz
Ce3q+lQF7KDC2p0FQVFAFxJi5C80bsfS8TyRPK4ZLOnGgI+JVFEJ0yvKXketISRo
hnq+AtYxiavZFZXfG5N0z+LgnXT8Nwllg8xTAYwvh5Rq9L5qy6vf8AQfMLzKAI5u
UQmT+XpW7W3s27JcariIh4+i7qM9ZiP09Y1q1IusbK8teEgF5UEGBoQKuj9wE3DE
m2mUa82zgw9GNYvis4LqqCa3u8KkUKwhs4iDdeB8/b2asjIs+wuIWupg12YvxKXE
iZ8FLWC9EifiiAGgrR3URhAyltaJRYdk55hWBy5fW7QtNBnT/AHdBqDlZep4tgs6
pDb8NKed54mGm3sVNIVBdgzYW6LMHNjRplz0xzkG9zx4Agh7+sOJmDU/i9hXEduY
JoCgUtrFiVksPf7wl91E7a9ppMr+lN2FjpLbDM9sEMEQppxbL2iac2fqymofD+84
eG39tUOHlGiplFr7rMBSzg7dG2LLVHlwXgj7oF8WhpmoiV4WOW2nDxeNHoA6343q
CH2EeX4B3wT98US/neZYGlpyXhBzA86V9Hj7XsFlM5GlFQKS82PAujsaEnYPOtXo
5Enz2PeUVmF+SGax1Ms5qkczZ+9SnhqyHeddO9HVcb30ICcOxbHO8Vn/PMLA01Vr
bSqLU7RWfs2igbWQPQ9yAcz/IAzaG1hifUWqlB8QVwVmIAScp3KbrUQRv7ZdhPfe
GYcNgroOtjRNhFskP3JVZdY2IJxwT8tPt8dcOIktvmSP+DNDhdTGZRo/V0YslNzc
UNQgSKZkbm7TibcxPZZrFqm2FUT6tKW1sMDASCsSox2ufAHudWuIpOQGPRu97wNV
/rpJunka4WRcgiz7ubQnVRkuhnqRS/NAXNAUghUG71I/LII8+c6W63CJXQeCJDFm
+6kCbzWBxFijCEvUMwSFzTCmICK4vHR6THXDZ8iEvmbwXnfxAOrs//yUFcX0Vcfo
1NFfZWVcfSFroYF/LGsUmxJpNI+VuSQP0p3V5+DVyTZcUPq2d4aAlZMDGzW9UBDM
z5qkZB/DUmiJg1hycemwt+ajJYx1xq82oK/f6AyPPkTAnNUE+XZmU9LqTA+QNqG9
5637SVrNf7OyvXWk+MYp2+/9jAh+6wgfio+AvFdF6bVX34JxItPmZY+3Npu0qQsn
hMcE5gMTcm1uavf9JtYXoDhqy3mQSin35BtjltV62n4BjN0dbFUxqJdgJbKC6u8s
SD5Sm7vyeyx+CFP2jWtVJ1jAwzQY88C8ZlN0G7wHyY7qUgntY1eSSjQzFqgciUjD
jcukyhRyUOg67BHcf8IBBIsur70KFres/SbX5ohA6tg7gZ/jiwXbRJ7kWeI3YGmN
Cfk4zzEnRVFWyWxJAsyeDPMuSg8UK+0/1bNozrMP7WHA+HPyvssgfY88llg0gOUp
doTxjLDZXy5BeqHbrF9jQOEgqasAj121r3GvLaKXdb8R4TSTPbRlNDccQRS8zQ4V
C1ok3gM9HN35G6iDZIKI+AYDdSOTJeXKgrYELjai3HBkbOYmDS+7j6rNW47/9UT7
m86pq2IsJj4P5dP9c60Mt2txNfClHZUFxXxSwmg+YhdhRWguqoxclDHpWi105Ne/
g/6SmMaayqEbhrc98Nx/1AvuZmWjSVG/YgZSkxj/dVydTeKK4PWvRr3k1dJ7FAK2
JJSdzJWhP/15NDlNIQOK5u75lo8VZEjWy+fMPmB8kEVTvgA+pbxI7Y6VvdhT+yiW
8CnLNtsuHVU7xVU2bHtuan2c1xLIhyLDL+1HYBKVAoG8YRXES8M55Qg8c6scXuPB
8uRDIiFCeN9RurBTvXzP0eMMpX8pVVJYLjNmenSnKKBvT4D2CVdAneEXBY2vlc0j
ldi6eHR5oLg2lgsv1bwfBBWTVTFWSIpniIluhZ8W7NfGlJ5GHKHk0/aF8iuJVjeD
owpm6whAkumEbPUS9kqXoVSBeXI/QyzvZXadrOsHebfV2BgQAoreG8GzUSbLRz3U
+8eEiOMLJu825qtQBsczVxuoKnLOH9GkGWVLvdbkmoSzejIQodxX1GqU21zfOyhT
mYqhJI6zhOzyoUfoWt+M4Q9wAUZVbCR2yYi7n9XKhASZ+hHOkv4tdGYUan/hVwxF
uS8xLj2+AYZVUFUXzlLzI+pHSSp6n56moohJwlJLeKCes4WULgrBXTw28TmsDT6R
ZDKHHRK0KoUONXAy3h6EaNTtDLninPMihz3NCCXzDqGhbS//hUbShxCZsSzAZqIH
Kb4ROdxHfM55nFIG1/2M0Y9VDqbCOrkj6I5rhC255v0w0qt/+5/A9dOfr3EqaCZi
qNnq/YCORJ3iRM8AollNp4RSNLdvAeU0APGXplhGpXk/eayw5oLA+4KfI62gqlfC
TwODxS92h7JuJevepOisruddkxbJ2nr4KEib+kCPVHBJkIu56RFGBSzJ6/B87KIT
jVA3MS8ML9L/EIktND23lYhLrNAY8jC6iRmHI232J5jgkZU8kps3Ll0ZKJFYITTj
Kf+tdXfdZ7bVNMbjjOBTu12wZFzpSof2fsq1LLpl6gZ+riFp1rYmWORijc+ibXLW
GinrTVBvsCRvYzO/DoUbViUbj1BslYUL+EV80T44cY0gh8hZKcetU+XUoIazpJ2K
TRgFMMRwTbFUix8WAwxlraL6aCJ0E8KE1dCTCJpPJRWrkmG42AAd9QY/eQGPugrW
SDjvKZ0rtChTEBIYfnA/IdK480j8INU90TuBqpuOVPnIbxOxPub4CdzOcZbeo1hE
AYJstfBJLpGou61W3a+vK3sCFKQ3aZsDSqAhT4p18y9Fu/ljEYXpUmWZ6bia4Ii0
DzMiQcDO39ljvq9nBZzA9XMlG29t8uL4rYYWXy2/ux5BUna5L6aoJcLlUKEJ5bte
86ZGN0ippDYlSJsNTwq+PbDYJupLX/wIp+0MDxnfsyIJgwby7uoiWdU/DZLHoehZ
oV+SiymENmcSYBVF8Bi+aXCF5ehB6jrMs6Z70ZPYIdoAeyq4UrTidxmINy2QW9Tc
pMPv+4Z9iwrs6QwPED+6/UnhxhW5EsZT22wfq0uIwhhhBMT0qFR/n7q/43ITiklo
sw7DlzBHAwHnMt6A3EoAU/Kv7cJuYSbc80eoKIad7Y9bA/VwzYSTNeOPrx+z3P9g
uRa718RwH1x8qjVRTO0i3UhG7mBV+ckK3iAuPeNgT4l9WILrbJf6YKKQT8oPdRbv
Vn8JjO++mPpU6t4GtqIhT6McYQmORjCu3tbn81gJei64PM8O8fhqQWkBNtPw2Jf7
iI8FFyjA3c9wOI2TQCprBR3GMMfPsp4vOliqFGqxqBX/kX50+bZp877iIw4aaGRk
on/DhzKq30svVBuH8Pk1Cpc27yyuEbm8YZhvWjXh9jrUJELff9cXsoizUIGLXgQW
SQD7xQfm5Eujo9uZT3OWmAPpFaiWDYxuKtb5PhYI96DxPOWIsjAKiP1AeHm0h4M1
wLzKSNJ0bGw/Rj6IdO1q6qThrZRhkns/MU2YUTBmS8HGP2egsOKlhoEJi9S1Lvs/
0t9A9103boV8S93qHyiHJYcCHqiBcHu9UMHRJlNWBNSfddYWlFGrfFixI/CaWENI
0N+9OXt33IVe+YoYmhlnCE/scEiTAiqVlS9sNTL+/ZUabTvW5727BM8Kr8nqqkz5
N0IDiibo/W9GE+R+o9PdEkBrrjcYnqkXj0m94Exe6jVaR1g4VgZd8yFoTrKzvJcZ
29IVq2At3Lpe1Z6h/dXTDz/FnNgzUZaQLOFXYUAuNTm6cH4mK103AQ0C+2HkbRah
XIjuI1DS1VoIjk/QH+E4tx6S8PkQC2l5W6BvVqQgXkJexxtpm78hCQFsEoaYOLRH
LjEWRC30j/V5sMIcyMrpYxWSjoQ4Y072OgE3WjEa8bCD2DdypUG4SildLuzItXlr
T3Svt2JdBXQISL0Ya0qmjkb7oj8k3O6ZMi+Y/rS6B5jhUu40q5/T7LlT/2jV9CPK
/tCduSeuOqsm1PP4adf5l9+zPVyJYke/BKxpnpSpJhFcshK1cwcI1++b8tMwV6YO
J8Ll8KDto7tBGUFsdaEYWz9efXV5hV1LuX6COUCLwGK+f6EgY2tLsMzMCHzws5sT
6A8dm0NDCw2cL7JLj04y/GkQRKaW1caUyp8i8ao8gBZK4BqaheevLqMJu/yIx1yE
/Btn2A4vbQMGynWbhtdaOCMzhb51L0lLnrzM0JCvTSLGLuBPQ3V53yyx8hD1Q8WF
KrW52p/wwtE52TFTbNfYopMlejHX2MK4mnGPoMZ1v+B5mxx58Sgbqfltr7Lk6W2e
omcRPWyMFod/JiW1d9JCcwir62+b9fhtx6qaRe19aWvHMbGe+E6jcMO17a+Vyn57
w8yGJ512plS65+yBECllofg3DYXS7u0ZbFbajLFludzlEn/sMec/o33S6aTjkf3x
JRLlnHTisIkZgLZJ06sjuv3Q0bC08XGuid+xYeV3Uq3nPCiTPqSVFBTwAkCi1kgr
vuwAV4zBifTHqfkllGHvP2qPJlnB9RhGS2f5JPABOXeRBhkO0o+JSwfV8OxkOBcV
10/tzNbs4qtD4ni9nwOtdAQLucP7L0AZc6PPdp0I3Tg8F4TVZb337Ny/YZqr2X+7
nNtDA2weLRT2C2e9NJ1vrb0gntu8PXSks8Ak9kM3ynDgwrm3+YlY+7IZMqi1P5px
4x6mMeWMDqRJPfM2YMkIq0GtQ/KFEorqg73J6zPBeESCxEePth8XeEf9mC/O4OCm
6dVTNQtvfo6gzpX4PPwzcSRAk/Ofl6tWsquqf2VYvqrcErfgdrr7OmMHIYc2NFpP
4lK3jKoRKBIix6lIWUrCExoaeLQa22Qu0e07cYPGlBHQpyGFpTdfcfaYWBET7nDL
3NSHZGbKflDCTDPvKWgWvYTO5wW/E4yaPAVvYNjwyr6HsS0MfnC/RDufIw4AY7CA
o9lwQneR0GupuqatanmaC2x1sZDqPgIC6eVl6GiidlA1couuMVs7LcMjiU7rIbbW
BkOzszMwF6tTt5WVsblE0w7s8Oz9fl3ZZSu9LzxVTDNivZhdBRHM8N9WyRuayRUs
GUijMSYhWrc2/p2TIQgXGKC23XGZKn1Glw/on1YXBgu3L8ZRj/9Twx8Up18yH8bA
VzA2yYDehCYsIiZl0e0VoToWZL65LYXw7vt/Ed3dqoT1QqSt0q2UqeFEXPpurmg7
GoKB2KkE1Er6LZebXwp37i6NQLhFRpfEftbR/UmDZj9SF2W4lAu64dCZSX5IIpN0
+NBgxFUr7hnrHha+k1zu1JH0XDoKK92D1L+K3K2ruf49U3FyUvgABUnMItuP3Y1m
Cna7bqqoDcAIPLT3dELqRk8OhNJWhqhM1kfiDgOM2GjO0jSFXmtzLr7Dqz9RNGmK
a5ggsmYd1aDgs4Zmzq6iPS6/DF0nUxHNlp0uoq0IEy1H7ZDBGt09ag9kjMYADEn5
xIoIXR8+rhSFAcYmzZGBUrzt5Sv7mrmLN+BDCqXnIXG2Db9fNwj6uFO30vwdIuqc
pwpeI92wtbbG1bChlFXFOXGajcXPzzyyYLKInm7la4oOGEBmANDWvzTYNSrurCgo
3i2mLeNbAO+QhgUQlJPxkWrKpE9yXMw4FXGC4oaIqBsefMHKevSYa4mgDsWVSVR9
2eKVBDH6ST4TXk+1m1bfWfOpCPfXEqEnIq6JDOECcGnLUORBZlFqVrtjKkpQ9poV
Q31GF551UgpqQeWQRqcbEr4Jwl97Ber1bHMraRGbwNyQK+5Jb/wkVysCAR4HJTYD
H4+eeEqQjETJFewSOGuWmnvevNJTrUI8B59IRu7y8w/WNOyId0syeQQkso5pcXts
tZScRHh1wkXXpEjLD1tTqn248CAikvaIzHACBpTPBbjTGQZJqc0fvFAgexUjhWKR
m74uw9VvavnZRIHsFlr2aH2wocbJNeMSZ33bUuJpz4VMXiLkBDI0DVJvfgVWmTH+
HNHM6ueeIkbofevq+Lr/lm3Te8BTRMuv2QICT50Wmfms02JGREFRzsVk/BHb6fBc
Ip1GBq7WUjclcJVqX7A0nP7vXBQR1py3HyN61GpyhijjT2luki3mMz8HNbcarz7X
CphjYcwQgQ6R3LKWWTZD0IUmBu9PH7DzbFh6tfgavORIYljFZmwReZ1J8k5n1jKr
c+vk6Z1xL+3uIhBoAWjL+IR2L+rqj6Lmv0BhsmB5ZPll4V9kANOuBdLtsq7eMTeL
FamHRKkw4ptK533Cg1XqfVaUwpH1qaCmDfHZyEwRKImFS52sY7EbKyALBJZn3WtU
QJP58s3bahP5069S+PmF0/RlfK+df6PfLBC0Shj2Vnzb43xHlHuHaCpi2AOWhz6b
TtYfwoW26lmy5nKSmfSTuqu/eXZ5TsxY38AXtpa7pkrtt6/yUw04FXdWqVcnJAKh
IoejfXkZuqPUS2UwwxO7XryMfiV805lvm4sKty1ldQPxxSpFMfdRQnVvW/RTc2MQ
QhQam1WGrOk71Vg2rQT4I1S9I/N/dKlT2cXGotWLophiL9aM5mPehSXWdl1M4xZL
2ml2iaJlaJb8zIQsbsPsMGgI8iZ7OsVotQaS4DQvUnKyEgPh/aRzINB3RN9+jBR2
GzBAkxscXjxt1ktVx0fowvWP49Xo4Z7WjSyGz0f4OvwH5YBRhCjheL9HC+qq0ZIb
Ycr/YsTWz5vlboiVPyURU6Qap/UiPIrmX8kJExk/dwMpt3vmg3WG+6i6S6cgKsG9
fbNkNFc1qVd0sCzwuJaTRRLPG2FODOfNrTud9nyFWIXEJtzQwFrA+FeHV48AfZU8
9RJxb3JUPwjMmubeIkr9KM7lFFKQ+SYV6RglfTo4AKc0IBN90xV7cnlPyuoBNhOU
YAhhj9dTgjasrdtqJ9baO7/Ga6EFlAVIfXJaYd1VXrTxhUbQio4JqdjaHoPh1VQe
kHxznvwB33ZV7buCLylR28OOuyyCO+JuTs7y3Bzhq4mZupezivDJNtdRo674Z1Fa
JomHnNTT0Al+Y7Q8jL3ugN0Qn/joN1pi75hL3ErsIlHB6PqTPv7Hureoy1GOQCyw
kVYSpgtdRayhl/Ys+pYJ6UEnjR9zQ5Wcjq0RiEyimNMp8oghKZvZRYkTENhSbwyo
d7n9r75kw1sVd3i/qOcddtwkGXUymjcGdMihNCZ5ivj2QzN7X1d62p2WVwsT0+MO
I45Z/uGcw9iZMzRQHmw1uA5e9uZlEX3bKJeFGdbOvgML6i/KW3Z19WSOjEUy+4Tf
7Iwwz9APEa4x1ZX5J5/yWD3q0nd+KeUY6xzyKg3i3pUiItAkGtk7LxFyOEE6zDVT
VSrO27vDVhfg6pGAoxllCxOVoT6RICyg8r8ZSwecF1gna0NFMDgEo6CSvk01xkdi
nvC7b0JvYksCgyYLaXdKslhQ0XJ4ltBt6HuroHY0k/4m123C/rfar/xaz7mYxNvH
JRuhL2YpMyDWzZZp7nd0sJoQjyP8lDRskMuuccth6XVePjpBMca9Nf4kOBC5cb8r
NnAARnhQmi3W/A5VYPTKR0Dlim0NLMyh+6eSD9IYU6C8IdSNPwzt0AiYKLO2Si6J
kyoQVlsItp3dQwBEHWabpdOcIpuKqBVQS13h2wkayXz0M9Tv6Toag58L+m9k/XJA
rMTu2G9TF1aiYmWz7J0s5psFfHBiPT66rkZosig8LbHN8jawg+aZtU+RwqBivta/
xvQoxjlkaLe92Ztlp+4sxR1tCjZ1crnSShCJU2hkptxVFN1j+ogceTGSp5Df9wJu
JhavVpMrvXHHTiEOtlgNY6PW47N2hHUUEv9WlzAT7RRfvN8TH3p7e5w6X8YyNiol
tT1vUiXaEgaKshgq+4kAdQRHXyUdEfcLU7pJwuhTemk1/XQvhGKqumzlByK7GoQm
yEdQ4IJOTeC76UWtM7qmy0trf7FWNcLZlIryrrB6DJPY7za/xiLFfnDTdJ5sTuvb
rhTtiqN+fUhtZCrI52M+uLm/ZlVRleZRyDMnItqjek/uMvmwbroe/H8CyvGFiNBr
QzjMt7FB6hLSveAWQ7S8KnFwtrtKtcMThky76HzxX7VA5SFvgH++XlPRgx3cgWLm
TqiwjsNZv6nzCkzLq/WujvtetoLS8CDYf1ODm5QPdqouuWJKw2eQVOjPwi/Ee9OV
xGxyp6em870ROmexWx6bvBpkf2GZ6p8lKQfa4ZwZL6KRKBV6n/uQfYUNe2LXNBRT
ZIIMjc5wM6zNYHKVMyzWmHlcR53H8jN612UzCFXd3h+QjFXCiO8P5GSrYPeC8HOF
ZcQtZqwydR72ia5f6EFn7PAcJ8KASHGqVfkGsCr2KOi/+SiBty6dZkmS7llMOgc+
NBQDCZ1Pl6FZ6IYxjLMI56xErj2GFnoehRVIC9MpvTJqzMt75hXoiVSdZa7GqlCt
59ojsL32CLbLTMwYKEp9ZBkRUWWFJs27zufdQPGHgAQuE9H4j3/lwFqhdKV5sBfW
OcdUlmM4WJRmDbq/NSBqwc4J7TSyM/Kmi4ttBV37mrUkl42TdzsZLo2lWJZysbjU
xFZZp2KL8N5pAUIwktxc5avm2rT0JE2wxWWnN7WVqZ/OOS0j7Jcqzmn9lyT7jOVB
37LF0LibOMxCwfJzZXDjIwEPaH6kirQTdW78owIT0zB0fYS1PcLxnY3yBTC9aVnW
6UsaxE/Ar7RdRQwBKne5eKn8qfCdm997zTk7TNH5N+9nc5Y6IMPc37R94Hj6vYSd
lwIAN3drf8qO+1SSYz3UK14a1wqh78HY56WwaUnam+dMgGnVZ9lsK7qrGCd7IpEr
WZ2Zl6cQd0biWoytjjyCtzKnoRtd2pe9obeaEY2a8T45NaG4cS0t9qylUvm1lj96
MdfyTj82fpT1W+V7F0P6TsmO38mNUDl5X2soZlWcoIrzGt17v/Y3URzLqUaBgren
tOH660rgilpfsW/HBqXnjHxq8xvmkboYxul6HBf7zxmO7BZJ0/6ewVGFHnwItR4U
Qv5LEd9i1vCUc5Ash7jtDHUi0lYlSyVw8oI8UpGkhrzqNez5K6Xdc3BEpmcZfVnq
6LJh1EiweTaIgDrGnkk9JPQuP0UI6gcgQAb0WHI+WJd183xqOG1ZVT0hYAHILaut
5tvmJ2bIWiiljtGaUdKy5koiIALycj4WENTW2/uXL+YYdE8GWIypYo9iZoKrmBfu
0t//tQFuz6jYetWPYOtpBXg6iNCG0NOu3KutMKYf1TqFl/WHRpzr/EHR6qxodqhC
qMCG5fPInzdV3/vYp3MIC4w5c+UTKct3li11nxWX6yW2YPQf/R8qvjqUBEiKIira
LdH0TMb2ER1NpobNkGL+8ps/hrcZoT5+2B40n/IdEYwMZ3zKEX0VBk5wBUdytjOy
PUFO+1JmBRrDVUdESnUdUsxbQ2sDBl7CbQZHsyxyVjy/y37Vf7WLEUw+oekrjuOE
fDu8I2MMqj8C0zfcAFX+DrYZir1z7YchpNsy3GILMNj3CnfbkK+v29y3Zf7Ed0RD
XZPb2/Dd75X9/Si5JKoLIhyPX4bjENGeEIqBDU5gtgGpY9TMYdIa5mr8f7On973Y
tWYl2u0OuWx/7peKctRNWpSDQbJ/MYkU7MNQOxPA7moB2Qj4/CXqhQRTR14Cffh/
zuxMnBI88QHm/DGvPEyZzNPheKJs8Zc7HU2sm3cHAvm+vZiseT8mzs5Aoz9i623K
3okOAiXqd+Lxn4bhEM/Flv9rMD1zyWOga7yD2GMjM1EWLmL5P3uNGoC8vloj1m67
VDO7x5vyX0L2qW/Q+kTw7+dVuMnnGBUPFlnYFP9SfQ8WenRoItpGZnQ6xplqgW9l
f/6n+Y3CwxT+MnRBHsbg5mWrEA6VkucKtVoyTPtNDbctffbi5XvmdgugW2ZZlD2D
5TLnQgVYrikHSa8XjsZUPHYcg0Mz+Rp/W+s8W5CVJ7+ARdOlCTIILvGFDX1lVlKv
sPr74a7QCdf3HstOt+4Q43HJQGbM6gSSbBo8O7NS56GnTk+LzxXlF/WyTDqinXFc
QnCqbMxqc4mMeKE/xsyVply6t3mC117RygIJWvPYdzWDDnzbxBo+lYnutW+re8fT
xl51Ly5LHsU0HkWpCaFql7W+M3/2N3hHXgWD5REThcm121Fzmfq2wElY2t7kyJVZ
eyIoRPxBE7oxWWcpr9QbbLEtwL9lkJX2x7ijIDbUS9z77nZQTd/VhFEUcSZAdda6
MmHavZ0eC3KIBvMaEm0KI7isb6yOixqI5HEgcgLvd9cMIon+Vibbp7U2SoruuZzj
KSlquYqcp4cgWMz2jr7w+Bt34XpxToy7wqYd2/54m++MPomWoLHGPMgA982cdlQ/
47wMiKuwCdDSaMMLTp/lOgYuJns2cc9x/ZKCOCpStiL3FqnV3g7MaaqMImlX2HTn
lHTN2fTpLw6E5yehdSAX8m1H2A/Z7cDxIwT1RsMUnDLDGy6+trK/vxhXjv3OR766
AbHvGQ64uzfE1XhB6AtguYsSpZJV0Cx49n6mayYRA+7SY/7uqZ7jgDgd242rPGm9
2NraS7u0p9+0Oc80/6E9Hp20NUAaZaRfdPXohoZ/FrSdErBPaW30MEK3d5uNtpci
ZJiCHcKPMFd1XzFw3GEKcKGcEYegegGUyO0g1V3H5TAWRv0QAueC078OTSnbJnmv
YGyWWpg8usEm7dL7sGWfeI9sc9jgLJOwprqVQjdpNgn2HySLSj+6SDv5KfifcCtW
XMKl3fHbpwXJvITBtf7xIsO705RymE3pCGzK9lsZ+G4yAai6CFfZUtnvoE/32D4K
5bGGwxvh2AJ80hGv0by+bOxEHHicUJIGnob40HwG1jxwLuBkaA6PeL7QtD/N0RwK
0Zm8Vbhbpz7hH+zdfo/qAA7N9dnBO9UJJhgBEzubPMlpOH8VBaeavD0CkzIynMjW
R6TO2jNiK0sAEP29sziq5XVS/PK03saioBQ/unXZJC/FeQktKe5lSw3kXLrlTXN/
dR1dUpuOSxrH5F7aufjJ3ktukFrj9EApymuo37z4cdWj3S+eknh6+wTAd79A9tlB
GBSzVAiKmAcvseb+nPR8nVX7du2HP8Qqxg2ATr4MDIA0DGTY88AjTF2KzgipGBOs
JgeyKEWZVBgMTZdHZ/feHspFW138fHdVBjnR6sIejuxynZQ6JP+YsYUkKeMXUOJX
alNy6o4FatjJwPBOTXIgxaD2KFtwDeC6er5h7X/SpcmX47tN6pQLD8eyanxTSk53
6zNmz0WW0FA9+IZCyfoecAHjqD+aF6f5C2bBEvW+4cUr7NfMYjAbYfumtrxble7Y
BLAQCOOJj0cEuUxmN2gyT3vfr6sWVih50FxxzARId0CRLywTQjHr7QMDRXtiYQqT
URDUhZ650qp1L5t7HM28io27OjSRTfta7fkE8FDojFSrTEdQq6ioLnM2TbEZLn5c
A1IlDE5Spc9153GUWnI6vZucEV9n+NQMps9FVqzoQ8dhQd/i/ERodjcstbXLNbaE
iLI1USKwshjF6FTTqo3+STRIoL0Aaaob9mOeFGnHP5vIBHrzkAJv0v6Hte3U3n0V
EO/cr7dTaAS2L+VhRYAXA7eVuRKN6fAZT40IIPKQDTk3B+NDcmKgWVhaHcxQW5z1
Mmpc3Kj6JzJWKwLcwhesQVXT6gcpYUquCgCwc4XA4/KT6SXVXWqjPTjft81bB7Bu
vQpPZi638mKDzLiDwL/ZDmsnNTyJDZ2UVSVvKEp9QRB/FRC6eCNJkXejG7IAOSSa
Z42ipbAmeUaABfwfzxp/lUTrV6nnMaS858TnYUwwPW62Y+uAInivzBkXQ1OQYow7
+byqgqQB9HRw6WRjSU/3tccsIevJAUGXfqX+OCwgbczjerjuxJdxeelVJGnpDJl2
pOZRMCxOMa5++2qZqACOt+Duk7efpZNHmMsF+uJpvDKySjzO6pzcFebGGnydGbAi
cRDpyG6i23rdoCDknP8VNXqNud3BDyUKmR+GQIBpY6FCbqOkqpTmSxPDaePaZsOs
C7veldu68nbMQW2YF4fpK+GzBytTXI9XQHllchKKMw8IXdTyPdriExu1JV0hSWst
3d/r1BgCRbWutfdHw9sFE+7mnkXAykm+kIFNVtc6EQ8Wn7B/2t82eM1/SVTjapCi
uK1ATiY6kfcpq/2kWUSJa/uL5yTBM0ppG8KiBCEhDAhjljElPfgYqtwoXhWVdIVB
BIUTA+moB52wCZ1fHLUhODY9az1loj0r0DYsff1zRIoNiIJZ7ceamA+V6YzKmL6C
IshBow0jQ7PuK6rPNJTAi/q3to8QTChjJ/Cr/LP8o9MW1LgK4q2qeL5F06Pkxhlq
049QtLJyrFNN/gHSW1O0RTRHmqvRNONpkDO8IcWwOogwBGeEDFW12vw8ofzOQ7JT
7QwOsUIHvDZr45rnQ/MZMNLzw1szHp6YXhDyjwyCDFRjh6RgTN8wMicuFBVy8ADA
zc3+W4d0Tk7xz5njmg05SF63AWhgqH7ZOj9U2fRuATuJgC5Aqj9yy0+JWCcM91wg
wvrO8NAYj2/koxnazQd5arMduL9O4DfY81VXHnvwRDnVJcZqbW8sx5GSb8mKpKhn
WxCy0b3KFo4bn0Ebwu/bLq5jXhDAyn28HGmX/GXxE17n2BhfWDOQMs7lA1bEYhFO
+FrQ2K7h7CWjJeSySymKhFoTKbUQ96g1rV3OO1HUlvu7045dZnRVsX5bgWLdh1nK
WG9Pyaw5JXyEI6n/V/3miT964HEEHwParPJJv7z+ouqecr2VAbU7jSq728NkHJQ0
1pZyZSzrTbQT2IK4qRI/YBN4T7lPGee8H2uDeEwWsy81U7GCjRSp2ZSEXBAwnvi0
CovDvXn92fcV/+zGEbo64zga9LzUiQ/gr+8Z7xk0B+yyrvTnIgBSc304VcQU/Pr3
2ZtaV/V6oL9hzD3eutFfayXUU2wyGO+gq8Hw7yL139Wel7NR+/O3EG4OMZl7OlgR
o06h4b+Oii94gjrBrXRkRfKxVNRU6SBdjiknD8GactTzTLaDb1/785V7jbYizDsh
g/zT60OwLZ9bEML9eSQZPRoLcQzZ02vsk/+lx2CI1eHTai21hxGeVsfHS4nKjh6A
swtYc2MxEEXZ582FfB6+MRq9Qlx3DGHN6YWPXgoEIxlFemo4Y5jGVkdqkxUk1rHy
/IYBzCHawiFnQ2HhjUbqZfCYOZplwfvyeJ0V9xGdkrC31hOwpmiRgPdFe7lQbq5i
jT/NMIfQEFEdm2K9B0/PVfjEcJZ44H45BoF7IheUfovRNYUHRtd/qq8c+fxfmm7E
G+swrPY+fOdeUwryZ3s5YEMhCEj9mjFoqJLlFAVMy62vcDuhWDLAFI9KlrUbK61v
LxDXAn3A8+ZJEPXxOqfHJyl5yepqJYAfVhb7Yl82lAXs/kMkf6yFnH/BWdSL8rFS
lOaf0OxlAXvSh3O9PbteX1p7GrZg+cnU6prVfAqPIL2qV0UQ6fdimHpQ9915K57G
2/u6//1PAp+7Tc4H6/S6PFrUW17Nrdm9i6migPqzERYsAWpSTliHaZ/mOODxzKuk
BuK21nR5nBL3rKkw2sF+8y+VLS/SjAdhlzlbdItQDoxwhCix0Fr/9UdScQPV6bUW
e6Ne2TbDrb4FGZ04rnHPc1/oeFhjBZqSt4YV2nsaEgfZAaCQ/xZa2b1Pi3/XR3na
N9TKfPTZRojFa+Ql2+R0Yo9SUr4sQVWcjj00mXuSacOTE1R2w0tHDozZVfTflnou
ysDrUjDCCkgDOn9UU0zrB0iUANiSmI4bcMDudVV9YRTnjl/QR4tVk+CvKOl/8pbL
4ZPG/xApykC6VNo2yhFQhkt3Tj/VNuDFcSwfNv27LnsXH014bwQj3j0gXc/B4Dri
zq36AkIslTrYndYjr/Rx1/vKHc8iksz43tzn7xdGiYwe2sdKRuNHtFPH45CxPWhB
xMW6tk4ht6aOzFzjr41EkaCwt+Y6y4g1bIdH486EX3oJu19APdFHuscJ6BrgJs1i
AhY5pk8G+OZdtxdYNP1j3bFKaMlzpW3PA9EoMxjOe686iBQapSNGNddF3fk4ND2e
VrWbxfstg9b8/X46dvJ0yEfKj72e3GmZ/GS9yTO6anw5VjtgMcSiSjOczr5HNzCU
LLvKuRxu5viwnzlpNzzOAosMSZW9/sAoLex2P7Sa33n0tLEW8lTbRYY3F7Tj3PMJ
8F7pA3vm52YKlFe1vQDxL0zsTRE7mWMZ4dlLssDdjxjiYafwWlnJ+yHF7lG7UHjU
Bbb2TYyxATFSPf28WL90UwWfL/uU4TPP8pKUMurCsZx4l53A7y9qaczm97g4N6wj
kVEgDMCUsfabN0O7TRNgkia+Jje6DrSOO5jHybo/NkIVFS1/D57FF9sBv4yFqBwt
nHauGo47Sv4ekH8nQf8+KwPxcdcZZ/hWXP1HwsPzALdNwtA1KMFFRPmJOovmIePa
mNCnGPdY8wDlTz9374gDjQ/RlQ3n8UNwG2WujVGzr0Hz2LvhuPV05uKvxRetFDyA
cAx4z/B55EeK/0sfRsA/v373+9oKUBi43x4lvTm2fkJJQI7qp/N4BaYReT1+m1TW
FwvwCqy7/nhyx46lf1dnNdcPoXmw/Hh25yceTdnhDn4hmV0U/yOTT9NP/oz+sC6F
YQMFVZdW5lv3Bw619XKzcLdRKfT0aLgVk4/gqVuc76xWlM1ROsTqSvEEWolOv82x
1fQ9YfAjOV0lPi9DIX0asiCV2wX6ZwlEoecr5Pg+Joyue+od60zckxJRMRtvhUhp
12gxvBU4aM5dPhY2wOMlltyQeXINPb2nhrhbIL5L1sj26B23SgcApomHNmw51lup
p4lrJBMP3zb0aq0iEoIvKBdRai40WhA8hR4gufyvOaG/A8tVC/JDi3j3YR3ra0Jc
f2rBHVOAhI6g/QyokuQHpzaroSvfueQuFywsmpIi7IqZ+/SIl37mb8i0X5PYSwUx
x78fADtgtsIq0azNFLAB/dyDU9MwNQELLjCIrl6Yjo6msgDGlg5KMw34AoTO3xUM
R0h9S3xOGoMhhektrzv4Z3bbs+w1l8pIF4nULS7FewFbtlU9t74Y1rLQnaUgXpRX
tfaT0V5Vldutc9hHX8SPVva5slbxkEcYaoGBkofwWTtWnBMOn1d4ow4rSlXMgETX
FLaH4IqAdUaVn904yukmJ/ZVohKkOFSStylzOeJohbyOQJ66eGmPQK+ekA0jQQu2
U8bWioh1z0DbGGTd9Oq0Ss4qqYCiHB1tDAmM35WecHg6NrZsOxBR1jIvWCmSunBt
h1siZ1jBdcdBefHYIaz+osUmYwwQvQ7S4aHU5ZkD3y6mAZ0H/I/GPNjc78sFhE/b
0MRTEb0sy3KE/X+nr8uNDkcWtizUTP1bHXLp1dMJZCVBWpa2musj/nwlms3O92uU
rUfXHBq+WGekxUaqYeDa6yt3dr+6OL0lGKVxS7b1U6GAziNEDnMPseeMYjcO2ITK
FOOb1lsQg6pJATC5fQedOafwzNP5enUiITrcGjbFwR/SmikZyiKZntbkfmVSj5gt
Zu+A/016v/AFJXjX53sQOYwNju5+4d26sweN2yDeP59sFhNrP7Tp4VtvzOHdlMBr
KzQne0gQJikJIklLsgHU2T/IuTdNQM2mLlU6I7KEJsQ3Q5VIqs7mCfqTAu++2dMR
sns2CGbCQPrFIlLoBMRqOa7C1zH4144ZGAcVhxmVVskcBUtmjCTjcM+rgggIKMcG
63jR/ni/fDi1WtDcVF+80Rs0Zkf2O4+MlDORY8rxF1ZqHoxzNEPcnoBedt1Pzl1V
8SJwrb7k4B4SRjel7Pig+Zehg6MYgiM9nCKS3WAfA6RJChWi5Cj5dETmVhfSt2TC
9Ov7UOh/P8g4424Gn3cv6rCt3u0t4aJNp1NZHqNCus1vWdBGusnxrreaCFlxI/YN
OMDxxzV9pMZ5jHJnv8w3Hnz6Ac0nPz53ye0abe3U4DWlE05kJJGnJie2Dk3y8UXW
vjefReL/gFGmtDhFVoB6//N1CcchmdpxKXI3ggrYDPpEfdJK5zgSk8f3sdek7Ee0
xO8mRPJFEDpVXQ8wdUBsXg2JyYG0OwrV017seHeXoM8uuoDe8OA24rSyq9r09qsP
aswestnGkYC5EntHMnWXa5LPjBe1KzZqBqwwZryA34PcqJDZDmTuP7OCIjzDWpXj
hHvc9EOwZ/uxvMl3bD/CV1fNQP/0KYisohAVBG2sMsjtBm02cosJrHEL/hIzAH4x
KEFvUY/yhXmS3JWuqQz8DNe5T/bo8MYVoXPcz340uVZJhIkV4+8tWvF9hGRRx7Rl
eK2Px34s7iRbsezIDwrq3pMsjpP9VoeRK9ThQlmSCSuNkw3Kgi3u94Yg9hcF1VSl
+ZskL2doMGNzEjJ8w/shjcCparuBpk46a6Nh/LudIAd5dGW/kZ6xwPAjKSpcULIz
gxgX92/2kjf2Zg+ju8EbfnKe5WdP9SrkN4ZG3Kkx8XbJmkMTqK55980sZpZye3/l
/tvXKBDWWYZobCX+N4HCUAChZ241X7+CVXsfqjjKcsOfRr7WWfdkvdrkMz0112ap
QBoPcsKmk6Carkq3Jcowikj8N62vlSB6jALe9qxJrCLpcAy05Tgbyor9MjQ12p+r
5B+skmZqJ98YxUoQQP0YrlreoXI+yK5PvLCYhdtpUcqIPZtgcuJKnRmROkPv+9Tg
ekhwiBSWVhVV+jxvP/JcOEskFHsJkS3RZ+VNeQqFOkGUAY43njxH1KlM2cNPEGO6
0r6lhQ+n1ST7XGMduhfQ1/e2J/qAddZkNHVSHM8SeKp0KPokHzShG2HEDYcsSgjy
g5U8oATE4O4fNHEwJ6pxyL03eUimnaP/BjgV67OG+MK///zWzLc9QdSy6VyZvaX5
uIe4T1EGnAKbofghY1B2ZAEqVzd+X3jGerZ8Ugs1e8JKW7zqUiz6A2ci9a6uxjiO
PoM7+UjZVlxOoiGsx9N05/2KVFdIqtiSZFXEEOZDKIS3ltLPFd5LamdcRZxLDK+A
b8UEFyJSKPFomqaEkRAxUlYCoUIZT3MdSAZ+jCtOXBuvDD9gmre8QdGimeuktOKa
nch5ORC/cpgtmeASUgHkh2/q/XzZNik68eVZBwzK6wKYPFVKocOLxeg4QkGkhwCR
vxi40u3rLbCugpgifuIG82g9QmxnaKXGwdHHt1TGjmm+I2W7oTkXqI4CrqUNILyi
U0oVuqdp0/63+JABKtXtlD5qJQFzzlMHQaShc6Kj61lwKnachTt9oWnEsj8vWQyy
L5+B7CcpNEb2vEBzKXecIrHIbfkzsFm7RXPqDuMDyv9zhxtj+qEIzEhO4GojgcwQ
1sZfMzsKxiliNaKtck7CSIwgSRhwI25vVadS7xHmSbkbrzsqm9w2M1Mk2T40rNbK
oFKrVyAZt5C7MbSxHEERaxQlFfNv/oQfEKccSV1RWP1WID5kSHph6cGkk1PCt/4G
ccVROSYGZoztliZBTiO8WPb+eLMofF4hahl9MigV5taLEnBl+PEzYTnnyPFzVAOr
7boYseSYvaxfytAEMtOLq550DhYRyuPR9d1E+lusbhBcUWVs1mj8Km2IlENyf4d/
bM6f8Zs03xfk/HcgN5rOIHevAlaqqqK3wJ2kMEwbLaO67ndthXJkU6CNUb/ZATah
sv9ga+Ku1uYbr/UJgsvtPsGnCyZwz5f0f5755B+EvyfGeTvPyVwYzulwTm9XzD7P
xfT8DffC0i+4ROVv9QNPo3BEpT1gyxxDgJ6fF35AoDnv0h/KCeTjBPoTtILca3E7
OusnONuMj849ZcPyOGPOhvwpagG9GSFzujGVARWjVcfO/+nmJEYIexhxbgKqviis
SLsLfgxfdPOTGSMPNkZ7twxcGsUo638ZlM+Muf+hwKOeEyf/Lc+tndsYdrw1WdK5
bm9l/3+SFserIdsFnbc6kkmmasSGhQfLVEMde6o9gfyseF0yIEh9iH12WO0PD3m5
QV6DYxFHcoMOmBAMDza4FxvnLWpOX3jxtk6hC1LLOBcX/WdWYOaOp1UQqe5mUaW9
/v0w+wd+WaQMnaC13SGZJ53nCDZP+fNge+e4yzSjVLV7aLQ6vVlm/fJeyZNur5yJ
I4RTEkrwj5NCvHLeC+Nh3JeMf36mAxOdSd3+DGpc3SLv8EOlcGyWI1Hr2mtl68bc
ksv4RNqPFUDuMU8nfp7jNyx0eK+ej+nfk2nlAvgjhEo4gowSZp8jtxnt1Inc00wy
+MmngCyqoBD4TW4Mz1Y0RXrf6u/grQqirPf7bdYbg6NviV6Dz0zMY528xCCzk1mx
+Ot+MOB0pXqRr/nbk43Loj+M66d3ThzZ0MQ94G7SFJh/bpLaCp+rw++DZ3hLtRh+
4ORDOiDTFHYr1fV/N7tr5VEtN72mUubgOvTfnVPR3RiNoX7P9HarqiC4U7Ma+hlE
zpBzP4TEZ7nEhxAb9Lg2AL6KU3tR+sd73H+yTErHx5cM78fvVts2IimqWkf8Iml8
+P8htu0B8jAyoYtyePA4xMhMgtuILJ+h1P56hG3SzWbymBfiL6H7RTe0U6pUBUCT
NGTFR7T3CxJIAU+fMJZsGmHr/fkk/dgZ3oyx3qG2oVzz9VI2AbhAWQsWatD4zjrc
s1wTBU1qFmT+hcHfln2G4bHRhKZQKwJXZGkxkp9Aelh4ubQodLLdkuQ+zjdMJ24f
hKIFMEShkucdxpW6W39DAWJeb3lzOPmCxqsD1Gk9Cy4itTY96s40UBNE/ClXgmbM
itFS5qbEzCDaqPxKnWwc+Z0gFtrUG8v20AQLjamUQzUydOxNYMcIPM7jjjCEjIMJ
ssETlxTVcWe3L4J8wc4tnSG4R9ujdsjaFz+0Qu5H/LIvW8zIh6hfPN3RpcKfldK7
6FphzcRZvOsLEleJ9r2WJ2VOZqyW884YTUNrhHM4hen3DWx1X0QRrtekmtKTwAgp
yKrC3W94csGPDyGKj/+6H3RCeuwjmwrO6zAtQfzO4JJJi2lc+md/WK51wWXgBVc6
JyBrU3htdtcxEse+GrkAQVYvVfXJkdE5rfPEYS8wsTGA9p+zyClG31ofInOOv/VH
F3sHzvMWevXes/+uq8zYZDdB45mh1ImlJe6ZdIHcdY41l/adN6f0rsgg+jgor+ja
9UpaGVBLGbzN6AU1xWa3ZxU8u2l2w+HXA/oobp+s9Qv0PKRvKxVwJCSR2s+ABW7N
1hqFZygA1SKD1/Y284zvbLD2lkFTruVpijW+UZ9XX6aunec8ojqps038wbJNgVse
HYkxx4Io+qgEWeu/pr49Az1NuxHZ2IKIvazMma+B8uhC8lprPTOZlkgS2g8K/Rws
9++YW3JFvgJ4+WJ9/L6oyEpDCSIdJ6zq3swzHvYrC82sLUlEX9mYvuo3pXvx4l5i
stkMuxwuprXk5OfO90MCetN/Ek6OR/V+3loSEWBCQc3cq249Lky4G1wj7sOPNPj6
ayIbnl6izRp2AmXl1yxtmy0oQk+21sL2np8XbhXL14cTWcMZc6edpaL297dtdfd/
7sXW/jLTBgQxXXs2DdDAtYgikG0XNlQ9mcHjNT/tPsutPYxhzDR6MS7XYLsWk6U/
mq2i4oP/rL/ah9mgez1ZHzyClAwAAlgYdujAV5wyR6Jp5/T/dAuClbQtMy+E7pE4
LeeIWAYuHMfiOJx5Wd2BCjO3HsEmdRo0moSvGS4rX+/LpzENhOY1WMTqtGCs5xNc
MisOpbnrTwQ0VlO1IheVOfgP2xfKaqoeAw3JTrdj4EYcLcrJID50ZGg3EuiJ5mbK
9OOKLuFPa15dkaJiDuzpT6NulvS0+y4hRkjG4vqlyFMx5dAzedjCkIMcp5d7sV6v
AU2USSHpi3QHc0AI+l0iloh90/8CC4uUJ2t5DT8ghut2uoLxgMUn0ICaHmifQvSp
SVY8vJ0o7bLyhAyKLBXkgTYSyxSbBgOXTUmdWuD00d6PrlCGIvX3weyEBBg431xn
ufl/NAJG8xV9LqNAN2SHMjjiUxKZrn505kgM6joK0hkODkuJVQ3rfO+PpeyfJVRJ
hvb2pRBEmzOCuTsHg3qczeXOR3AdVzZryeM1hhkwj3lvWuTmRCycWMhCiE++Qeir
Khi194eQBy8M0km+USc4KmfPsmfzq1HmfvOWiZ8xnhRHJmVHK5jwaDYIqEKLd33G
y7uYlc0aDqQ5sZ4ktHd1IHIgqPq+AIEhPb6oxnGKxesCFfIzIlqdOe2EmyLrGApP
TeYWBQA3Z4VqNu/6wM/Vh27ETZ9UPrCKl1YJXAw+8DpJnEN1o6pNcnlqMUy39IGM
sn7zwY0GU/+4He7SbFcZQERBL+fieaiF3eCY+uE0cRN0tezSZGUg4ATS9mWIJz8C
qwwusXGnb7EYRe0Itt1fnf5+j3Jkqizl8dOPNnCGZ4PAIQOeyhSY2XHqgfxxWriY
UPODe+3svUCyRKYRMpA9EfDQrQ2dUOe8lKiv/JtIz1lVgJ0DmjWarFmNpoZpiCvH
Wf+oqfAl+aKb3gMAB7dx/cmjttN6l2Qt54w03L6FreBIZkHTVjWG3IQoCldwe3GU
JJJOUCABc49itjJ2AlCoPWXQGxYZtrsmWw+zXGkSOpSLLFkzA0W7aOu59buCp7ib
YJ/pVcoyMWEqd0q7NdJWvJSKGzMk7Nv/hgAx0lW34hT8mRlRM5WjUzeW5c0OWteX
ZOBTa9nolcN3iXJK50s55uzF2yARpNLf2cthi8Ueg8eJziB8kJosOKnwFt9uEDoJ
JDhLVO02E5q3bmFcxtVFtKo+dodGD69dOBy/TrdIr1FOWEYsqEA06SEIfo7QfzWk
FQeSHCwgCOjcELH+1VHc2hw6W/Jc5hENgfNm8hLR6uIGF+xi392n2RVOUfhkbjez
uZ101ch4Y3oZ0Qc8pUDXabvzpGYTL7kNiKhrCXmL2qpU4KLp6qccpXPg6KXYOeoA
4tbUrD+zBb09IXGJTYYnB5dny1QTZatVguAAOKgcvgrL8suZKWcKIJG3z+UEPdi5
T1CUmwumF5PZucmUKIN1UMFtMncWBBFbM5ZOWSul2qM8hKVNRKsCmluTQ7M72Ncu
dyB6lSSknJ501f58KaIwnKooYcrCWp8rdZJDhc9CEmMDRUz1D80dLNB9YtB5e6BK
i5xdzpvSu/snQ05SW8WIa7JpelrlnDf2GqQgt9PRPFLmQyW28b8Y+wnJaYOMokip
2CQdNyiddh1amfPZX1dU+5qqpFr/nJdAKNi6MuIRc99K2lk29/wP54yoVMjkN5bA
2CeQTG3Jj9up+20RhTw0fT1Tut0KptEjzoHhbHYNRRiLn9KaOb7y/E7KdzRKESAW
5ddTrNU5/gs6LRiRPziPHiD925CXFmzOZnIaJrIhqezpSblTOwJeRPKtBwrGX4Ir
pkGNisoRo0lZjyvydySWOQtUH+GlTbIx2lGufxsaSPn8Un5uaMMrS4AiGchycA2G
WwJ3dtFFLeBlzUUgOFGl61hMrBczRkkrB63yE0UheDdkLXKYXVE7JRhkMPJjw6qP
GdiQ2S7ne9GCeW/U3/UlpOcrcDxsiiVFnXVZE/NOYzf18TaB1wxc8unk93UQ1x9h
0KrHlmdu2eMwxTYQsgqkcDQ7XkDrDCFzlaWCqDO1TMITuKFDMJn5u6kql1b0c/Ww
BJCk7+UqhJx4AlLQfx+kfn9C5NnwkkkO0vtkGfnn7Z+/hYylNAOt/w9XpenN8eb+
T61JO/li3s1nY/hc5jvExKt62mT8om+NRVhG2+4SP5KhlyTgimMgP/3RyjGgKfXG
V08hxiTuZu+D4JK2tLYRL0coQQr67yYh94T/eYm2OZWWjj4bYOkbvoctGpPY/BW5
svsc1Ds8AIArDK6OS9uGF/LShVJTkwIEJcS4duGgCYFRcJeNf6OHWkkEpclrRZe9
R1a1jZshKALzqGPGOh9pwHpgqMrH+p3UqdVsD7x8oBqls8KpAEKt4eEO8ZTyTa64
j/K/7qV7ZaK283xshXlq+7iFD8GG0+VL0Fe52OFYe0mXDtNCZcGWJzZqnG/dHdvK
oOfJcXmArxSlpFHXEEYnobPvssayPDfpAN2lvO3pL3iLozbgeTdlvPRpK3ElPkGm
+uhkLAvocVLphxjzLKjvAcucsQ1kFyIfLRwvYwxF7te/cMxwB+Bn9eiJoPmPviGb
DN8CTmkNQi8hMRO28W8XbMvmi/9hh4XSTf89qMCVNDaaWjVkpSbIA4w7g3shI40r
jlLg459w6ACq78v99Sax6dd3JRnOJl1GnyHAnzr1K2az6zRKV4tvokkkpXBXJL/C
Spzgc7uch1ufWV43Eyj/Yj0oXmdoKWheG6naxdm1W29DdsTXNUhnBJ8D2Pt47cGR
eUDSTXAxjZ9QGO5V7M6o98sbwGK/IerfYrNCL32SeAhbSDQk8S6D9jzYIm4YQUrQ
cNo8YBFjYIDdoK1tk0PH/OvSKtgk8TwoIqRRODMoEhvPlge1Jr/UpaK00Jjy7aWa
PYwmA3JlRyjPt4LDLE1DtqySDS9MbsNAEl6IVuxujmZeJiKt1CgK0SAnrvgXjaQQ
kmZN/et3sRP/W/nZtj4xP1t4YJoPfHl9eiU0YYQ6PUgmCsSV4lVlDLdlS++UCToX
wsioCBiP5hy4w+HqxXyLoRfo87FxU7uIii6EQiyzVbqNu8MHeGU2G4WUuEPg76tl
A4asq7G5eW4Uy9v0GUYjrmVhvt4Eo1XR84lRrMyhTo7lapwJ1PPIUjTLBo7w4HQH
odG2vmuAFiGTvMiHZcANpHA32eFJzpSadeTkh2ByphCXPhXkJKJPETjO5qvnQEZW
4Xt2a5PBjmF81GZvW5JXiMSLZd7LrHc3RxucrKikyaB+ekTA+0u2BIqJBAgoJvk2
mh5gzOBnk0FKBUmWjRi/+x2GwgX5P6XiocsAjtGSu/G/2AsfjoG/PQUqucUxUH8q
z0mrsXb/IdWP266COpBjKhT2BVwwS4x2LRffOKkr8uhhRefazVbpzhz84i896fMf
GaEmpGd09zL94bneET0zcCUa9fEUSHD53FtF5ArAaDmVGCkUZdLhGU4IPWRn5Ohv
NoITLUvulHG4FL96jaeP95CpzDt/oNV5y39KNxga5S5lqApDA0xXRIBGG93a2hLJ
Uxuv8pmuMggkpeiwtdLZ0Ziw/lTL59v7SF4+J5pv7MiivjEYyueh4DIvDH3SR2Np
Tj4erSS6s0pRKe8lfpREdYp4hNTzFw4BkWb7QPEf72njBqUHQlnDfG/ZmTyyZMkg
NaLD7lVjuilIeBrIxvZlBiHy/8MDy/Eo1yqMN85cfMEebz0Rt4kmrup3zm9GgdxR
YhUQldcoCnPmfNIIkqhMtudtwFrZHJOSHo4Eoxzdf+zDDotfxipoLfI36cw5DEQQ
RDIsbOHMQjS7wpWer7VXS+5LXQynOLZCdN/TlguqIcnRQWJOOGRajgGhvB+Vpl8w
jhuL9jlRdnB7SWUxYuk6QRT0CP9/NEHMIUJX/uG+vTsBGMnu5iLCfBvFknSO7qWl
sRkUZakIAZ1bSMCUJbKaTee+mdpj2gjudtgwy3sj0k9yQHk1VgL3lWnoJOzXIWF3
GG4FsZQOfJ8Js/Xx1TzhWNUjimOvG1/oRBJ2SWAtc7jisLuAAvqdTkvFBQ6/Rs5r
bs6E/cvU/0Y5NDB+dB1V+bQbcqx1Wm5romrg7r/y/R8KNd+88YivsyFeXxQDswfN
VLN1eD+Yb0NIF6g+Gg9tIH3gqyyKl+aT7p2DQMVXuU9ICn65lA9U37CqZRYCC00y
JEalK/taThV7QS2WCvJ4eqRVa7sMVWmXlqQWRqIjdtBqs/TkADalFMzTFvEEs03i
egNKZBA5TYFnPk4mYfC+z8FZESIM68RmUDSz5Nl5H7QPbm2c9EE9iN5pSrtDNsKv
ZwEswAINtXQWcU1hXOR6sToznVhHuGgt+mLYIKPQAYrJIrBZe+mvEJXuLsUji7Cl
qNpz3RRRYPpGrIKRV3rZadkleD2sQVbRlZ6EaWU1VkxG4ICHulfQhdrO2tlXek/p
n4NYcndF82Wd12YgPYZDnCO2CX2wVGn4BFNqeoK4GbtW+Aah61duN+npLMqeAhE9
MdrCUpyuYfLwU0q4X12IS+yLK4eKi+/VlRs05+LleGBw6oVg6l3i1cL3cuepiLmq
btBryU/wRwl8qrWbqnCqm8dhigpszEucUeHponwbNm9BGGP9j60gA5tbv6sRz1aZ
TVJW0hBjzlBVWM+R7X/FGL+QjXRlQOevasqU3ePbMMc4EQ3L3ARHp8VJETAyO+pU
NcZuSwSDZ81sFk8tLBlHL/JOJ1AiqQBxwzz5aSbCkOpWb2NE4jwigy0CEgx1J2+u
X1RzRc5vceLJja7wofMnWFNAVvPTg1IWwbgseLzeUWOkKWbaYPh8Y0YmBzF9dhvn
wXle+/CYMbik8y2FDG2mdCT4ocGL4tJiWSdt4/+FsbgP7DY/8xm3EKiMyqsmqZhO
9ebJGDeuhhn4hJooIMem4Acte2cs6mBdwL8w8CIEui7FTrUNQnjknUxQHpzdMh1v
LXo5bf0vbCBT9H+zEG7Nw15vmIFPDOUfDdV2z/V9q8cTzMp1nJunD2ZAFQUtwV6v
J+dUBURMm8oKmUMwak+Fp+1cB4mIHT+P+CLSyPFP0ISRwVd5uzM0whpHDnAnrLUw
D2PRNVW7b0o/6XjXD1T1QpH/35bT+EqU/hELPMY9UJnXY6XsmAxw5BfTECIBG6iX
hZxndLzkXG1FebhaC64FQM+hINCAcc1N4cj8KSq1BisYaoxKMqkqiEWRKztnIM4L
YjqT7LWzY7hAJ2FE2syRm5JbcubH/XrRHaZiyT49Jcf5Vj9MOpNh6OaR3JIYv7Qf
Tn5eZ6J5XDoDMa92ihOuJnbt6uhYBbzt2+T0SqV1fse3MIUwrFWv7oUZTvwKHWlf
X12dxMU3ZIHL8O8EYtXmoWvJaGL2YqraJJnmGhC4b+eJJnsvdZJBTDUgEw+SuavT
8794mtCxPHyM5gQUGoqRmbD7XaUMRnDffFSUmIPPaW7wymh9lzsu6Mt5/93DPhFa
OnGS9JsSXE69ah4Yjy4vmvIR3T1yPxm0Kqb7AVKEDWjyU0J03Qdfn2fBh1xOZYuQ
hH4Ba3p2mA8RbQBkbymBz85n03z81mcvO30cbt9VeZKx1/E5Lntfy9bH4M32B7/4
PCtf10FbqCTRThCL0Csmo3ikb8eNuamSF0d6MAmIPmuCREFQgxIU5mH522D6T6pS
a9r+gEn9X8C2ajT3JZZK9RThHfLcjiSAdv7C7woBLCXxEXGe6MgRgnoXfcwYPrV3
ShoLhHbz6+5HfqsjC80dLuf5pVmyy+ojDCTp631vtrDGvOBpacZ3CCogtlaXG5zC
5N5yGZIYJtKEJXpfFZ2vn1p6tZs2PxCvCS7P1dcgimAmpdHxRCQj1FdFS9MhHHLU
oB5nD1bSgmwR7P08yzzBVlIocJXHHXGMhjY9MpnGdqicoVFuwiaSOtlLSwY4ec2P
yLCim6c/Nn5WB5IlDByQDUF5tW25wEK5VrK9qS1YALb3PC7N2jsCG75De1KoWuls
3nGf9GRlbOqu9r/OlWQmRu+yHq17dNQXX6Oz6WqziNlyAAIPualmpG8r4vxtXK9v
C50N5OAZ7PE6Je1H3irwdai6zRIOXIZIomBxsF7bu/pS2doiMLXJOyIhtGen6Xln
y7Pg4zMn1j8t6l4wQM7aTTjhnrSZjPepAyG5VgYAhHiDiR6Av6PJq/w4E53SXyWx
XZJ0pBNNPDF3atfpRGoRGv8TT07PkaE5qf+I9vqM1vPA+yoMYZvZdU/RcOBgx8uX
N8muxnMokcxCGLg9q1zq+URUIxb5NifcaUHxTWmQz23spHa/LCcHS3KGdXVA/mpU
t7lxWlt0X/mtZSKtsG0QViQLlRl05f5tvyX7Q89ZtZAEtV4zmrAUB7kjqnKAGDeW
hYQ5a+O3iojbOWsAuY5YNkK2dQGjHBH8kTywpl6tjjSwIY0KpD8a0cRfpbE+sLJ7
/yC+FlrIsJK4cU9mgWMPn0RnNm4+Ixzrn6nVHVTfZdgAufMnNpOiIsGpzcDngOxG
QKig6pI4OsJ67NcEiUNBAhsA9tZSzAw0vbIpCGlrSd8pgtHyss1DLTRZBNIRTdl+
6ds7PnxJpDVgRjFHUMsX3ZnSnt2Py92C7Gu7z1XMy5vaxihuTOl2AHXqIQ4qlzlo
JSY0U/52KHYZ8KHgl+/FZWNPIIFm0LU6oEldJ9wySNA1jpYSVFW0rPDQ8bQdqnXX
GrJeHbS9o4fIGc1m1zkWC5565apBw0RBu+WameppDEBtKkt72K/HJ3Iv9Sz3xjVf
zcY2KBhVtleKsGqiKuXwM8iuI5++NOSfR71ZR4wcdlJLiVcRmkPKT/pQ5G1DCZTY
j5F0rMMDuVHhxcHg90TR95VAvtF503/pY1xgk/T6gFhQ+C7hMoqeUHLLQGuQNxn1
CSzHGdjsuMKZgU7bCRL6wjtbZe7oyQLrXNK4BlvNhKSxcxNHQE1LULj8GiTS7lT8
Xo6aTw1CEpFQAfVrIoHPbOMo25akc/m3xcZy5XvHI2WU082IQiWZfzW1UMLF9y7B
f25OhzFX0uCJborprLoh14tNCw8tTSjHkQfBc701Lb+poNuWjAoIBfk39uzAWVdW
G5GldDu/S6IUK0xXeuFplVlaxDLanmut0MCa4HAxsJuwPtmbt7sZ17lEwLl5Bwpj
h8Z/11CC6wVy5GPD/hYIkjXdczMUIpoAKT8I7hqcV+b2zmgBJMq/jmJBh3rR4qCg
xgR0VyFPULiTve/3zh7GyBCUzFLQMmzCnk9ix35IujlrsAjvO2rcV25/fkRJ96Qa
gU6EgVwZ8oZU16uhQTi0b36QAEHCtcY8PDeOkoAcIXb3G1PBh8ACYsq1Y0KkOjaW
BFO5CoRmjXC9hFec0wLOsYkrFn0xm1He3fHK1JCFr6XPbe82OvswejgKb9bq914W
p269KgvELf4SH/9ndj3Gm618J9jBab4f1iQTzixH+F0hWmTthAoKObVDuuqt35EL
gZUjqzGTEkjLnBlTRcKxQByUC/NfRDUwpLMsKtxu5Ld/0FjYdBxvHOx4GVgmG9Kn
CB0fc/LKf19alSkiE/b7jQcYHdAxufSPEyLkNvTL32g3SiP29VnIvlZqAniAzTEH
C/YpZ2f2BKWAMkpnMPB6V+35FuCK/vxJ4bDXkqclyUc/mR4p1pYfNXvBRmFMYgxL
n+JZDH7zEksgEQAJqXlnmBjerjz9tt5I5IJEPJ8LbU34pdeT6mTKuNNs+TL/Wwux
mLRenFN6+qH6FQ4kTQefP1DEfd9cRkjoxmn0XFL5G8iHYu8ELIZfCMCjK3TtnLyo
k+qAQIeaOxKa/apD27ow7CecYXz2bAJVVIx4ffajdr5XbP9TiTAYaGc0EiULMG/v
qp5CWz3UINPIPkF8nzFqbk3PgQedxuRIqJJMY68ez4H+FgZPg0spbRM82OSiNlnf
jhJ557SofdZybRsscILSU6PyDtHx0AKws9FSZSRutzCdl5i52P4mTkq7aJPi0pXt
akFTjFlRULcXi3Zgy+T6N4uQNYmvxMhCJHiuOwVroEkOAiw57xRhEPqGSdn6TU75
g6XIAzGMyUDpNXCvWff6b2V6yn1DzuCXa+r1hXGupk+JiMDIkhhYDZK3aUbtQqb6
pAljPis/ALAQBQl1r8ketSNDTKyAIBXvsJ2FQGVONbdyzz3gaReFmRi2jAAIoJ99
V07rAeQPg7T/atscxDyFi6PGN504lOi+z6ERO38niEo6kYTvJ5tM4SEDju/++DfO
e2xo/3m1Srpb0PDF66H9+CoUX/13XywpJFG61cACnMj6y6KAwEtEtdmLnVOVb8KV
dV3yNl+hagiEQ24hilL8rmKccvZdkuuyG72tGgSqdzRp4HU2XKCLokslF/9eeN3S
85+ryfqCtXV9BJLlERWuLai0SbUn3UO1Xnkcfpoi5nInEqXVmV3tt3MsMKA1t5MA
QScCXIy1qQDJsp7mnVV/I8YKt7Tqf7vYQxFz5WLfdSGxE1djPFPm5QoWZ7wZMC82
zZSETFfwAmr2/ce/NdLs2oIfq7P35us0KiIyxLGXeAbHS21GaE0F9qxXSFfs3HP0
Kkf6ACvXgWsQFtJccWhZmPSL+gFITTTbNmTW4GxXp/vjZN5QA5DmsKWFaAfPZ47W
2MYpld+wbK3lezAzpH/zwM3ptz7mNdrLCdmR2Er+TXkX24CdrGjCsU+8Fkwvf/mY
50kGzWpUn83SnxCQCMm5tmIvjsp/WsOig+/FgUbarwdGiF97HIJKnWw0Fz6E1zUe
uvbbOmo83gP6aXpxiTfY/NwOoONtMwaMJNFjrNvTcbLaeKPiQDSbRZljw3eFLRNw
/QVTrBpjsphx29HJX/31p45Y0MEqdnmqdUlMBJJVgJ/Yb6z1WNT/dCrEnT9nrG4c
w2g5ayJ5/w4mnypl/yFR76+TKRF47Oi9j0nKiqW3Fu89Ki6xLhhQ6GIOFjaV6GAg
5hRwt7IHfsZbU8b3igcJhhjRsI/wl6lsizn/xa1u6Ntgr3cd2gqkCeAkUi+Sql0I
yIxVamg+FuVLyy19WUA4mFS9vuuawlNxx9ZYaN13AdeVt+UmK8ofJ34+3VMSBUq3
Is6pJPbQSRaPjMXMVMx92heaAaixmh1zfEJ1efUHVe8Ru1VURqRdS8VZi8c0u+ao
aGSyyMuO34e2+5P6cEx64GvQ0FEyV1k6efoM328D2fiGuQcoSA+IwK9ts3/2N8h9
Cd/ezTclbx90TUVx8DOSO6svhgH85yiIulZCJUFEvmM+8PCvLseqiqnjMtk+EE7B
YZFy5CwAe8domIj5lzOt4oKy44KXQdLaAWKulnFQeOmvXcSI1Duk1gisirGqB5in
qHl6N41vgTJTQYTBw1w52TnnyOGK7VWROEGD7sGMz2nhMySLnYJl9Jo8Yc3QOjP4
8ou1uhe+bYPL7vpGa/eLj+COwyQLBg76+HTrIoZ5IBLv3OAr3kqREd9FZenUeH1N
nqhOPlmIij0utR6F5AYsh5dhflncbZsCD70W1qEKz9uI4cD9illkOvV/0IFsA/Og
wthnAs0D39p2dZ1Abv/4G5z4GdJWhpxToMgfY0tjJyatxDeVIAtPE1ZhkOsQNU6i
p/3riSkExioIqQEf9+s4XQJwpE/vc8k/kZYHunBOEwy8Miu4Ik9ya+YjU4wYCZDA
t0/KMZbtIo8hjuTTeavHV4kL/lZ8MTjT2LJPNtCdaDKMQtsdMPygernzcem+SLpK
SQMxoc9Gc8Wr6za/ojCXdSDQzj3jMsG067vKlmSMrg9swUKwM/F0NzYQg1EGjgyj
KUypjssnszrtnFgDcF+Tb6m7NS7eS7pNXdLXtMS573+IQ0LvrdmugwkliUSRLBaL
aC0xv5qR9M2bt3GAhidBeVQ2OcFFN9e504B8DVAB+IFJ2F1jk0Sc2+IHj79GMuWO
Nho0nseBzRCESYgpcn038+uxVjvNObLIK6fw2X2at8rEbezIWYxxuhL04tTg0aRD
5pNxpJkeG7Doxd6+btt26ZCjMt6V4rkXfEu+nuboO52oFUspKBB6pSqQPnIFLYUc
UfQz2rVruhMROV5oCeea5SmuSKRiVlOVosxeRQ+VbqJKFJKvRrxvFaVOog0eMuiw
4kuIrO0UXY9PR062DFVZkBcA0PtWB5t+oTHNn9QxNchQ05r42rpmtosk0XMZYk9Y
5twc/YqhGHeXWCosnCdUXyZcOmMhzGoQHJBEJUz8qFrcPhz+LuSSqjkju00sT5sS
sCl4tKjLGj309JDTiBN2bjZlExt5kJ2nwRYMXRR/TTPG5eVdnadp2zTAABv/QH2A
ALPeSpYK/Sv317desecFEaZ60B0QsWeLbAVo44FcdTFl+Wjc8jW6PQH+LVi08GCA
139e9JUaBb9kNjGNccdAGFIu0k6f5272xteCTU5PaXRBrNbDuOUL29q1nxqa3pz3
nHF/xS2/rH2fB1qWtMLumt000IweXCm1pVwfd5TFs7XhRbMa+CXPkVfxYdY08dFF
oP5SGjz4foKkTZWuZUk1bmW+FyBKs55CCl7lqjPFqXzxWKx3prkKBuLOFWWLJ8mA
awRLYjJ0p+nMH8TWBdUsgEjJScjSBYc/gRsE/+TCEyU80dZatpBF59TV0mSkoudj
LhzR/9IqV1arcEhLY07wkH9YIxHF/+Riu4WH+NxEbwa5IcEydZSGyIves4s+TtiV
XHnvaISgcJvzqPoOArNmVx4CfevEKswVfXq0XnGK2SodkhodGGDsuhMZSaOuZ6xE
TTobXl6JmrcThYO1dbg4cQ6g3T1BueNUJ1mzRMCuhvGWDrbw90NjQHbbsgeulbxf
RmhzTuuvbgttjN+BHeER2hUBOwsbMq8cenPzW1qHUTfjQKsEhEnqaiWsIvEoYJBN
U2W50Oi7FoQRh8MTU6CFceTk7KR5D4jsS5NAyZLM/294jHeNPhAt07H+76fSFLQx
oomrGDuhPl7+uZdokXUQV9c5vRQLhhZg0cF8+vrs1BIfRPGjcKSMgpt1mEU9zD5f
tSGWRPLTgte9VAtH0wc7Yc+JtUEr2/a4BRzryBERsq1gl1b6gBDu3bq5n+4lB7B1
BOJEEQ/TuHBzVqNkun49jhcoaeqHY4uFIYNlnq0CsjNe64nJMYFChp2bQyk4aXQg
HXFtpTL4uHJIytHZK1xTk9SvSIHY6VmWu1sFNrurtOercXmyBhY/is8ad6qBrEF2
dg/WfzPaSyk4aUp9s3BvwyzRDijgQAsKze/YwhUAeGWbDN3dR7ebqaJp571prcIq
ERP0T2k6H5UzK4DgBzv1zZ2azcIQvjQj1CWOwOyaqR4UnslhXr/LECHUKzMlK5QB
4V6RnjtbxFF1WDJoqptNrrpXIS6aQxyFOwQAqz3Ux754UViy5wOk2PPBFx9kjHtf
iOt2iXDyfvepz02VSx/lMfwhjJ1GO79SUjPzpBr20d+alZ0ulALjSKU1rgfaD1mj
JHEb7PLny//Z7B2g8bO8OIYi+I8iEi2iZsLTnAMV6W38HT9FZm9gaw+xt+UGnTdM
z5ruue48JljydgzzdD3v/WCe4IQ8quvilubW6R9PTomrO2f4tuClJMT3/d8WJMOZ
NGAcBwbwYizJjK2RdP+UlN+rbbYsTUQRNu2BFXwRC8h+lvsEDIUXsbvvuMKOcv5+
z9Cv8VNfuk+4CZuJe/byapAwy55fJC0VFh8yDyo6LwnXOHjasfYc4tibE1t1IXuM
3+m1689AzBOL5jdsQ7LePQO6Sr0lx0O2voY+kt0uDyewzlDvT5XWF4wHVZ9Kynet
YqNUdUmpmZT8IXylIx4Ba5a/Sv6PkUa3JLcMyxg7Kt/Ojyl3exTg28LbhMgKAf9U
RRh84p8iBwE+0Fom2SFzsn14ZW4OXNPEo1Zh7E/Xh6jsmTFlbn9cSArTzGaSbZHa
+BkNPT3HjF/WmC60Y1tlm2clSd1vNahs8VsD8XROdI87m3KsEOVijgUxVVanl9M0
Z8vvKkrDvKasxfojwQHCEmLrxEVmASp6uiGPC273gyRYAhLqQR5878CYJ2Ap7Yfr
5yvl6khZQFa5llC00DXZMg/xID99l+dNTQamVm75x/wq7dWE2VmAZbsJk5XBKJY4
QTaZeg7u4/ZWrFjWhpzZA2qNOg5FYfPqMa2oHn5G7bdgiLCBjGPc2Wzp43NoKwXq
G+EtkWj4Zzj4xRbImJg1LtyulG7GJT5UEGbVJ/FG9FfbhC0w8wkKQ/1f9egE4l+o
0/A2Q3JZtpUrcuANJ7eVu6mb1ZZYK8QgVI4hkUAl632XeTTS41y5e5AooL+qDtWd
i5xzSK0Ek5H8y5XEJ2V1Porg3lKbGJCetpd8yHSBiL5iijZrWoqWlTFb9ESUtlPY
DmcYIRZ35QO6PlEwH+gms6RcprUQ4OgzGFDw7HYsnAS7hu/CiA1kyj90TpnGj1jm
QakJYtNtjU5Bz/FA0m/j4laQCnUnmpwEuQ6uLd4AaPIPGvjvN8ERZVGyJwm+zRjd
uYdz7TeHRSVIe1520RneYqiFutCzSHZla0+Q4aVU5xMgfj76ZpUEYTxhd+DCHkFA
7oJg5RFC0sqfXMdospkJq+uBc5DMqxz1kw8Pfs7ppjnwbWMw0ThskOP4AIfNefZd
IDnFQQXpR62IrJM1fDft4s4qF29NrMGYeStv/o3yo2uwbnVo6cLGBwkEwjp+F+FI
MD9A2WgBHzY19SO6su+/npBKpgejcnM+FyeL8vHGTmRYT7IWvNeZLBeev+bDwCF8
yK9T1rbRmQ/cOiEKTANwkazIOYOlFPfcJ8/RpT74RgH/PzwS50/xZexFXGFzxwYk
hYnYSPqOiP31aNvgcaBy634ZhVzMeg/qrCvhBseaGgv6h+ndLeR8swAQXuDg52TK
SH/rCuzcyNB6nmzSN4i9n/+2FrFrlNLR3zETscFRl3lkbGJxRPnT+AZeCdeU8av3
qyEFTr6Wc4KgAzdHjjPC0q01rMcyaDj4mW0o64aWI27k4AIr59BBJtvrtqmkXCln
W6DQslvxVQAxGASvVv92n5+W/MhLyTb3LhM4AOi4XXQ3tPn6ruXI/cYOsQqEHprW
CcJeFdT5UoIQcqahgtaKE1fiOh/EOmUA6HwLzBptBulM3lueL45NNe2F0K7jF0p0
V5A8vsULMlTYb8Ht1uOhvm47SDXLE85uwPqbAtVeiz3UP1RuBivwQan3YSlhW1vz
paBalBVvkAtr3dt5sWNZ8wfwTlh6Y4VGeWSvSfqoWo+T3DGLRF5EKk4dRaE+WyZQ
VNuXPLhBjIFZQbR3y/VOyULLrvC5u+zcY2gEXDChGfrCsoyZjAQfpUsQorVIZjBo
rqPgqrfqkNBfEQ1HD8Vz0AKWzgdllwcS2E6K+UPZD3SzC/whLxKU+TvJSqo+QSqa
AFH4EgLVgjPONvjDt0tKC30faN72A3Y8ovsLMWF77qIVq1qzf+pVToU6b+mhi22w
WAZcIXU66uu2BTNVO0TDW8k8CFiAbDG4tZ8cZ/dhjZWLnbWNSQOkW3H0099v1/1T
UUiu4CDaT+XQDQ6Qo0ygm9dw9MNA1iQNbc4gMus7vT3c0FPwCrt2JjSpfo/F//IB
lTSHbk8PoWWKnOHa/ek2z6BXdQPoIcNH28Rl93lLACDiP8z0WldrFhiqLiKN4y7/
FV/f7Qgr+OvK1cQzsecBIyAGc1nIlFAdUdRBADjAZ0UTwTMsdockyJ6WJG/CHk8e
wZbSyW5VOir55wnNKIP90KvFXQJlhgmAg3tvRHkiYE+ZfYVll90ZDWui2Eb+AVAZ
0Oczx0JXRDVc16dEoZButoIjtdCZZJ7KCK6MEKgerQ1xOc5DwJ5X2U4FXcp1jcWH
TSZjcmzYo4GtVSQ2GpNkIZq3JQDziwnnRd8I60PPKw4Lz21kFHsyqySggc0mFN4m
xSqYfT5nNF2/32rcP25QA8FmX8TI1CHLA/FHwsIxbBk0zF4L12tjcfeFj8zYVmWo
gRUQAhlXcdk6A0wLpthF4O+K6+y9F9o3VOGLBMseWG2W2vZi7qHzwaVXs3AlDhGB
w8qVYIRacsS8aSPZzkUYWNXA50e+XV8uBnzvhcpRdSGQLZ5zQnOjYZgddb61FC8l
xkrEkMzzjnbpcY9xgKwWdeRncdTnBhOZ9pToQmsw/RcU2jeqh30AIPsQGGWIdYOT
kmwD/UnHD80AQMw/4I3RfSpwZ9LLDX+REGcE/Tj9xTtLnYJ25fyJq2kG9S7sdh4d
O/YgYYQrPHTCyS7OlZ/1xbK5rjbl78H7kXjIxrLYjMEcaOJ0TgiVW9dor0jctePe
xC72GH47bZCLfBRqPL8OUA1CULjEygzqX3Yfl0Wy6YcRjFHEKfryw8CZsjK450/3
n5GPHiRH7ofkBsC+MwhY8CczRODQj2t8+HJr9cO/xV3kuMMFVkgQJyVfMdmnB2/g
rO/o+79Ft1EkLT+FNsWfpYnK94wAl9sT0SarblWkhN5L+oql7eCWrmgJ5ZICPZGO
oNCw3OqK0n+CeA1lm7QJUXNERGOSjwcrMnKAHqqCAkQMyi4EvC0ubHgb1ae0tWNR
1hBJDhJLiPFErj3E2oj0Vwum1aJiVe6Vyek9u3jM7lbta4gKHr3b09ylBaoH4N8W
0C1T7vRNfBz/j3onHTIGWoirJT/hgEYUE8QME5G11ax2djBtcHmcY4F2COjfmH0o
2Ek4X6/YbCIiKWde+jrcm1aAdTRSuf1rmNNsOfZf7VNs8CLrY83/w+AyV9FOrloI
WTu3sU3Z8MfgnJhD2aFcFOhTvATEd4ewJwwrRXikvtuo8iglCf4MFHHulRF57nHl
ZwEzDXaqk82bAgpjjql+3+PCZyVjsAJXXjxOVm+BQdbRZ41lfs1XqPRIqqQndcSP
3aoM139TWi4PZRUzMsUTQDnLydmFtdLo53GMkbehyzvZOuqtkY8mjHXAv1ni5zkg
gz+58sPLKzcUP8MQJFyCx0A6TrhKzc+ZIJ2eWZPhKGbEKRjRzFJevNGyvdrA3toc
gGhUTj/n6Ls0gQux0gJgaQm2Ob6ut5xbuYJJMfzR7INImldwRRLzwFcVN61x/hc3
f3Gb2JfPBBAijigTY3DtWM671yzLY1XhA5ubx/8qBWjw0oy1/aUqTAOPUZlax/0d
rxgMOqCIgkzKZPED294Ji295d/vG2pgv3hPZngazsjJPR4udmv7tQX/T3COV8yUZ
k+xgREjN07TwMxRx4RhfArCFDTRhj2PsljYR1T79t1yoon1Um3wsFmmpylbAsxu5
7lZ3MCARUPJsZ3XpIXOq2FLXS3VDPAe6AMhnKyClmjcGlj9cSTZcD6jRUX3Pb3h5
vqF6Yiw8a/82UOMeVMHt7TDLFilWeFsJnLFAy7jsmBaQYEw0Y1fNQHHpZ7W6+Sh/
aEdGUNMI9/yCG76k/GO9WI58Qt3TVI/xzGrhTy4J06vzMvSwK78yfLRrVcI3Ezgw
WLIm01GLO1QznEYodjN2Qw5hJ/S0P8xgGf6v5tA2b713qStLPRmxBp5tNNGGNEew
qb1LUuVddWpt3cUoFbH9L57pR1PnvyS+yQSpQBaDvS0mv1RmehnmrXlHGHL52x9d
7WXPFK9CXgWaQ0DH5m2fMZOHxAIwAxenztTNabgld0XO8tGiq+89i7Tns9RFwrZx
eFIVjAdAVNnoYhOE7f9TOsVCi1CrPYVg4Xu5ohabTfFZUW0eH3+N7574j1LpWgUE
p3h6CV7e/x5WeR9uZwzAu5dqTWD4cmxkKiE/i7f3qHqd06uvvjAXlSzPMQFz2/Ic
Dj9bX1bM7/oT6A3bVZF5O3KJ2G3fXY95qL+GFUjPMVI5344qbnFVbfqnSgEYbUvC
wHiYi0YQa7W0EoX2lHhLLP4U1PJlPS+2fwm4geEGw5efq7lFWTr0vWVob+okzMQM
basFuYKAdWdz7GO7cNcFoxjX1LT61Mz0iA/hsDYsphpPSQCTHMprt6HaTTqdyggY
HCvugycQssZONQm41PKV8NfAOOD6MHArHw3tZhz/La7R/JHXquIHRURypyrn8Rif
BIvt8Wea+Sm1tB7Up3uC3yp9n/2OnAAgywMnzbZbzAACtxsYz6sqKt15j2+sut8b
bFtqtLURNMgovuXMcZBTJZ5fl7J1zRXLkdrpqmAMn3wf+HkxqAxxPyO4UAKwFzmX
U4vcDz+LkQP8wk6vSzPjz7MsS6w59CUQSNHjdunj05Iqpqnw/nLPJH5vyMwfq4Xt
cS+tUgWaNpU+og4k5fvz1BPiX/TzLT4ahj4TwXRP9fzpcdZISnW8IAD/ZVwsBDK5
TA2sa7MxhJ9g3V6hQn2s6ZBBTuFOL5hF3dtMb8MmK36iVqf+RVS/i3eKReA1CPJW
CF2KLi47BahaBy8AqgAouAu+/qo747xsZnzd9aIfnJQ6X6rJYBr9XALcexUhIujF
5K91/3DfZJRSLujJbh55qNpoL9FpUL8E4Enb9tN0HEWV8MmcMVamtFafMOnE57JX
SspPtsslhJPZlObuo4kGnnRCAk2tnK4DYrQ3nePQB0h3TgxgE05AI2hG4qsNQfO5
ziXRoygB80iydRCcTvip++YfzXxVV8ix71dhClJX3gvQhRrU0aTvHqyXgMgSqGxX
Zwv2CJ47KZ2Kp+RtDVx7a0WzaWEujHLv6DY29eson6Ax7ehi2Y++Tlu4zz8uDCRB
AUEqeRu840lEyiBhCHuBSwrxsLBqF6PiuN4PeA8en/rMrdLm7kRmo2hsPnofNkbQ
MYFVRbzIhOFFAxkb7Vsw98MzdSaB8n5p+Bi1C2Mcm6WEXn0qLbcQMiDDYruyIM5H
f41shJ67d05kJh5dZI+YVWzu/07czsMKcNVUqdCLWaOR5OHVxGSVZiIkit38yhNJ
KDEvGL7lBx+CGwT2N0KFoQvs95XBwDNssCwW+1x/Je1JBfEsGn/O6zvZwnycaeU5
5KgwNeDpr55P1cNO6XSAcFjCnZH79skeuekmkUaH3SC/2iTNnkwHJbx9vu+efz4C
ctmm8c1DtVxdHuku7s3oXrsJhPTQyrtZXAH0CDEw86J6xTsLNccsblZb6K3gkDvW
yKq0Qx8TNCA3oNZ7zxvQtDlla1Q9sUmYG0zCU5Jgcz3i0ZVmWmM6ozUEZ/GPaz9Y
T6vhW1FdtDaCceEMut0pvKMW2NVpgDaqEkBwdsrc5NAaZJIg3owIvVcTe9nuh8Xc
DjwMFfaJp5uZXcbDmEvtMZJikz/gp7T4+LXYf8396xxFbpo/XnnyBmqDeF7HzEQ+
E9svbjnCZcStvLQOjFLtDdfVMPd/DSFfp5/OtgZJx2IW2xQTE0g6iZhbQpfh90z5
3WefBf/uh+aJr9k39dyJqSQte9sfOKJsVqeATQZUFRpVA38uhHTOx5DFzt6AqwbA
tqiqAzXSUU3mOuYue181WUh9RLPYqXmaRg7qB+Ve3FeeLyknjj/OOgRMlMZOP212
r1K5ZAwN4iPT1f4+9fiH+9rYvX0zKevPLpE6lMJlGm14suL2+ob+PF3BNyT9wv8W
MMUAvTuO6ffw3GpuCaIPQ8TDYcX9wZ7Jb5Rsr6oz0xZdmKm3aRcGStXiaUOTrDjF
i6IGsAPnHkH9cCozdlHhJrmekQ/+xylrWsU5rEh5oJQGBHCTMbwAfXIaqHsHIHnI
FPUQ7Pxjt4vwNAGT7O6jo9av8AMkwDRgVabjQ6lFSpnzv6PsV/bPPfsPwelD1J1e
sHdjudWfioyEOs5sDI57XPnk68tqqfwQm9j/E6Wp8BaC5lc5NLDB2SiDhQ/6QXQL
omlqVr/YXgWs1X+5Z8fSr2O4C7S1l9NuTEPVcKs9p/bqJn4H/4sLWbcIUTbexBQX
weRBSgvuMGKnYPdvsOT363baT5H4OyA4cDyGCtR3lPkV4IidUlCa6FQ3VQiW+Q3a
bf6h2ADOWVtmW3JX4gKpY7WE7xT3l4qd0B+Izy54CfhJaqqfrwoaK3nn322yt5LS
j2hZHz4ZxzDaioBGBNKCgtl79Usb1GmpsPVkJpvhv/BwyS+/HgnaiOnngLfft7qN
pihVe+ElK2QenuVVkPqWFyyu9gwF3ZcjxzzB4GfJFF2+ZVJQ6urUm+Awu1h/nqQ9
Hke6x4Nhx4Y7+e1Rxq+SIAkvDrPK1pghSFibsv+G3wKcPueQuxOQcmZ44QZzKva1
I6MoIo9AaeLO1kmPQA60/IsfDummLjyc7Q8R5QpmAGYe09dKSYSqK/0rUr3aHwDH
Ingv86Z6S75aVnPhOM+x6ABUOJCxYmWLjkArev7rl6su/Lgetzf545/mkIQK734W
E57OfB+/q+cuU+FayIyn9VrsgsuQXulRQKNyLsNT6CkTvoGeCfWFfGwHnEYmY5XC
qIh2wkl/SO7peCagTxxLib/NzCEnRrAn/pEY5+CLG//h5Y2GSUG86FWG1JhhsX71
+wC6JydbgOynDtovpVoo9HE3hUA/CUgwZIuebwqyFe/hOXO38zFo24jos5A4Bee8
LnBIoqxfZpMUtKWn6TMUgXYxLAiLkd8ooH3ToihS4E0mL5Mhz5hxwRBpDpKvZUGn
e7S66FVs2vHUIkbjrYjc2QUTc/Mc8+Y5jqYpaYJYANdQTfRUM6eczKbX6R4wsDxm
xNhgdVodjQHViPoVqlYr37+qajRWngcu+RqBYKpUUlQDKLBTKjP6Om3IJW67RAFv
gnu2ea8xUolRWMgVqjnMtI3IPIpimrh3GgbYt2PC+h3a3WoMNtf0ABugqi9gS5Fb
eV8s6maD4JCvn8Xpp6FUALHpeUQKAsEJtwxRlEYLQ3zS3nBrgsT2lm4MNH+JtG8x
c63sb2A2c1sw6gMPTyF66yFdRCvuHL0lbbq7KZw8TDthKrGKe8bng4r0qxoyyaUU
fzFGsbCYBas6QmebNusUsoXec9KCMN3j5C7b30oFwNlxSWkQINAd4ggJEvJJAN1j
LWNBK7/oxh4MjGCPP/HuaG4rprjpN/Cl88tWBVfx+mAIZOERFRashhaEviYshpxt
5lplzeVS0Vk8XnDAbrih1hKgSu1227quDJ8jbCZt2WcQYTvXDnHPRb5JCSvA3t31
jVlSfBc5lzWa8QqhaXft6SGwG85gZ1q04lhin/DO1vJa/wbSMi+IzuTzgBTGlqfT
r7XzLBZ9tlw0VUNRAyHRcu6m8GV6xynkl4UFy1Ipq83ZdzeJrVY0ym5H7m+S1XJk
N5yJPGS9slkV4ANILfyvmbwgaOg8Z/Aeh6aWRueaOJ8x6svkx2l5JI5shD0GKOeF
3RkhVkssQ8ruYXzsvGmakv08bj/oo46EaKv/GGyRvggDTmHfjaeOZEr4JpLGP6ud
GPCu+87DdgbGCkiAQ+STzkxpbfJBvwNWl0TVyY2Wx4UykuIr5cUtPDNuIhN3XWbg
ocXWJGsV8cYxF0M+uYM5Dp7pJQ5iCigAfOKUXb9JBv2oNoENedk92R+YNCNBCjb7
YYYuZ+kQAOVVt2uM47odVndIJKoJJY4SIWjdpnhTbmC/lkVgClye7/spqFNQs/5u
58uv9IZd+pVBp3d7QYE0Fz1CEHnCXegMq7nCXHWC0mI1TWRmPz9xmoVxafUWEpF+
ojqzACh9Slzt4Ese867SqhPR8EZ5d3LZdaKlE/W7uwmhQvO8CCnrl9fhg/NrY/iW
8MuDbqphi/TKxaV6U+1ue0rVM/Ed/WGv7wPVhJF1RJgEHH6eDo641YaHBiiG3YeH
rM0oxgsy4MqUmqfrSP0a0OsZonjT0lzURLQLfBsWQsabw66RBx70F8B9IbKnkni4
O2oLIQA6TNth2bIcSKDPFXLh93RgBNscpoPuccGteV+e9qydu3YrfjzK1a5qX6I6
4HwUXpUVKbheV3WLpuf3uaBrJUhbsmgnSVaTZ8HCzvzqIgfL0WDkRxQKUcsCR4pN
wkLsiX3vOWy1/g/XD+rL0VrGkTg6vBIiluAIZaZTuRWFapNVvZ7/gZaS+ZqhXWuX
DqU9oq696GjbJ/MulkuFL0Iavu8u5vui6Qp62WNHjiJR7rtCrzvaueEiH6W+BBYu
X4kM8H7/azu5/Y5zYJmgNSwSaJIm/vV2pzynttHhDdg4cmt3TshGrEmkLOwUGu+Q
fkzDH1ridZT2TZsevJyLFGMPX8xsZshYHGmUIEvYACnrUp/EiieKWpR2GM77u+VC
JBzCddRdinDtUlK6Znp4qHM3BD8tXca5g/TL4hcTwOTeGWXMoWgGBK0A6BDnh+6Z
R8aoKcfDiYQQd3diPtG2e69Rke9KRt4Hy/rr1sbwAeCWOUtqQ/AQQ+J8Kn1TZ+vT
HfsUMExaA6h329E5kUcTqYbPpKSEiiSMfURCViXFxvjBr7e9QoYs45TU9IMy1og4
DJVR+HlRfk1ow/pPkP4si8wBzKQZEQb4HIosUl26l+KeiiGeFRMTMiatfG6aSCUg
If+KesXqsfeTy/klRshRLueacXKC+pGKKIQUQSegufqAvBJ+PPo2Ex0oSsiCSkBO
2I0nSumGFkaFoekXaIJgCSvZ/Tb+veLVM+kt+hBoisna10Da+O7aMaACMWksusGf
wSME67lLqy2VxjA7D/t2qCQEFvGym4lj+HZRgOPPjQrwJGvkv9qybee05135kVCx
kAvGkvuLu1RmVQRWksX7V2DTuJiZyXNgAloE4l1eoq2Ak+Uc5wP0mUgl6sGf7rA0
4vibyLlwGo4DF5D3gzDgSyKL3ejJv1Omug1OimjFi1YqjmJyKxwBSvrtpx2qfwie
g90qkMXvnvsalhjssBXlA9rzN7hktDG+x41nHKLQ/WrBAhM7WEsWIJCQdPDfisqJ
7zbkg4qsmKIntQJAONDAqGRzfucbceeEGzBpCuVZ+pzZToTv6/6WBHZhcwG6Bszp
Am+p5XJSnsHNDPOXQEeb8dfAj8oua9Q9x7tIiIaVKKUWTLeHcuiY/inhgY5tTPEK
yM/HTxujOH+Ix5FpyI6mAF28kbOxCUcvg711c240WI6DbTZxRBMj3SvjqdUOB6sr
R8gFJWZfyGMwPzxeu1GrdG4u2Cvi70CuzhKH5MeNSg0VCK5O4eaLT51ba/3kvbUN
kNBhNsLaOlJfF7Yn1j3EJYBKqsyc+daa4cRSL/lJNrGSIv7663DV1l2VtgW1BnsE
Qr+zqp1vligX2v5fi1ZvUVzg9h7UMH1M1KHnPApAZPZMqf7HzfPNxI9ByI0TWnAr
gC6hzlFraNIsWtFcly6aSSj+gQ5Ub1a+i2zWnOwKqbhizq5A73X/CNkGniRNKXGT
usPBEbX5EXN0EdSwn4KxWSsI9RRzWjS7nrOAzTHF8qgARHqluymzgEWizRXkUa23
iMXsoRhRo53mdUipqcy6YUyN/zJmFObHT/cZHGx6uaMCE/HOVJ1xs/i8oHoGXMBN
VHicNWnpiW9adzdlm5QHDJDl/07GhWVGdZZapceM3uv4fQw7Sv6MddBmF74bwpr7
M/OeG14MhJULI/O0cyK44HBMNtz9XUsiIbFJaZRBqTPn40asF8J21h5EtsSjusaC
aVxzGD/qscAPCvC1SsRENpFQxxBNdkTlIArPx2T+Qo/quQ/HwnMcTHD+962wNOWK
EJIMBc9NEIyzo0j6At/WSomifjw3C06WcwOnYSL+EpUnYt7SCGgGnqNMaOA3BhVi
Estv69bXJ8qHr3XRAmmilBDXcDzEawWxIYQ/5Io26d1Ir5A+jywY542QZdSjE7sV
EXW0kX+SFC519dJwFGbFUlfKLYMky9+mS7L7ftvAx6z41pvC1wYyiAve/VbfDV7D
duis3bHEb5PfUrhHeC8exv/MzVLkJHgQAuZNNspjp+O9W4gA1yqa5GAC4wpS88Qz
FCXvgMlbeDONATNHJkZsHYLFKOuVXew9ItO7Wjq2JDcxSH5F1Bf3YalJOkO5XxIk
47tyGjQgF/zX0KzETwHTIJichGj9dx4vVFpDuxGLarhay8vfQvgySXukLpW6W2aD
/vbmO2ghXHDpr7InfVa+MLRdPFBEAjwzq2wUqxsxx/KTLyViTwi5n6TvwmJgpRnI
j8dWRMtUG3EvoOsd1AOuisvlGuwFn7au83sTD63KUqlg+WsJFKdErym6++O7teC6
RBevQjMCmFXETB5VbLzkitt8QjuIoFT4u1sjrt8GPTvbcLifb9qU28IEcuPvUWoR
F5ZpWU2gv3+NOv7F8BoAQh+hOBn8xO8e4vzYco/vSEjz1YV3xEvq/f89ezBfTdLk
pDdUr5noCFg9wzD4cpSd2bIXx9880K/E/ixcX1InzdwbJ9gZi0B6JgVMn5Wy/sQT
/5jZVNbMmsL3ATn/Diuj3JeTWbkQxcb069nJTwS45qGMdCaB6rlKE0XnxU3Wvc+g
Mx9tdUsi+UDtU8Lsx2fdV9IvYSOOawtnEiucnIsq7g6NIDWrBkGOhddTHgcYyg2K
a8Yt2SQ7nZzDKKhazSSfkCgxbX9DHbSsmpaONH1BYgTvJagPH9f7KCeLzM/i4SNn
D+Lox5kBEhaCHeBl8JvMMJFwPfMXRFDLbJrAaTA/1u/YUYEjK30Kdq9GYdyl/PEW
4JjXJ0Pzl6OMJUJTZ7FVXgN5ZM7uZXqTVCWcgek8AjoiwgtBXg9Ymiq//zg5Nv8J
E5lXKH7WkfvP3x5yypEDJI1ueDincUTz6K5t54sJ/fJjL1khpCV2nXcKmz+bpc3B
5wMjm57UmWhtdj8T7rubthDGNHAdNtlylHa7PiGZ1C4MNxijAMjBQ8ejK13d9SqR
G9vHOzGVerZ3gcSHT+xfUvetYfdAWQWzbw1EalfC6Y9YfhyLdy3x6/lPo1rLU1xk
xzObHSdYhPj/zkVyZG4aoJ4RtSU+epcuxKZME/SbwHrnVVgMtVN62fKwBxItlv3/
LuYsS5XsVP7LblODZOZ/vA37rGc/l2I7CqXhIH+ny099kTUsql5NmGkYV7/2lyRE
qLURa4dWdQQKTfeC97FUzMLklGP1sjHqp3Tv9J01X8bfrLliUpf+W4aSs1xOJjH/
mvLohOXC/su0yc1N5/K6Ng7iKoeCymxRexldUqZ5CAul0KJfT6Wr78+Agj1emTL7
P/j6/ryM0L9zHcT/Iy6011pV0FN80c8yBcOdKwTnjFqMR3L5bnbmUVirO9s3a2N/
wekWY19OQFvT/8rMz/cJs0GGZZ8yIeVh7QM2QeMi9OnafPqDXTCM5jDZO5An7biw
ca9d1kknN1UXT4yzwa7rfDqTen2jO23E0hfA9WD2U/DjY9T7Gkam/x9xgM5gwksc
1IrJwTRvt32zZaQtnmdzniyrHC7M0u2Oyt1K5bDbOQAWDOGFrVV2AJqMHy1PyizB
nV7yd/2cZurx7+mQnMbmD7aAYYDnIHJOGKEfxdMn9AqzRQC7VFgIcdz3yd3dTYRS
9DYG0chUw16XM8N47HdEcjzcmDwiAHPUvyB/YIsvrSTxpcj6R//hIMBOdKqkN0qu
LuSb3dUYg+PdXX+2KipRi/pRhr+mLyK0fqb4QlpsS1HvRL3yZ1D3GuD24/55zNXx
7WDQdx5CimudNFDay01Xyl4L6L8r7vqkOb6SUVE7pdcfesPWLmNAx3uzQkjen5hX
6zlLl336qmje4Ja9xl8DhyGQ0EYr6pkxbWf5m7Hs6X8KY5ylXpYuszRuuVMU1jkT
BgcViyoVECIO4fm/NVM/JyoF08U5YC+VTIKv+KdIQrDtppn+DVIvOjXP/qxqnDcJ
g7L8uzwoV3+QzGlDgwO//DTGooMDz5FpliwK7EyrjeFj1e9FZwns/iM/Psq7xo3G
D2/OhxFmHcK+Cv5U9/p7YTc5vg76aZTUVZz1j7TRK9bybngibb+gSAGMX2gIvWU4
+ZD+Ul4K1jYwPhX9Ox7P60BbJwC88RzGWeMg5CCgf0XvSev847s62aiJe7kbex0P
BF7sTbUXgKnFRtdlyRvLl2HLwkvyD9fTzXQMy5yPsNwmAXgvoRMzArUu2+gafZoP
QxuLtdrBKv2276vBMaXNBOtasEh306PVF1AGmUwkycPf3T1mMfqwtJU19X2MAtsX
+koNdfQ7fiozz4lXMhanfZ0Gyo/HQsTW0WTToBk0BLVSEW/ebY1mRnHv/cJDAIEc
JWds9Ua2B8qlkQcJ7edXIU7jAI8dBdEAytTnjtfzi30p0OZHN8c0wAOiQzdcbEXS
Eac1trhG6RhudAH3ytYNGV+DLeATIzZeki0MtJiJCN7kRfchDl84WEr2/b7/NbI1
9XrPcTdaGdS0W5fOSXN2MGI3YVPp8MMLrf0h/4HrDZ1gw7mPonXqHkgTULQYhQvb
T41xUcJYCpqrFyxrWsNEjT/pZOaBUrIGveYiqQKwL0fJvex/P/ZUjJY5rd/CoKcl
2iil4vKo0L+G77wAncwkiPfF6dahZUpTCZYTbyQMFlGsXCjukY5xDfx+2eXFrkzR
cSgQhh9jaoSiYV1LkzU7QqLVc/tQRiVApKjQKENS8ocDUOavbxhAbNYkA6QZR0sf
/rbZtDudha0+qMuFX86jRJqNcH4iZ7fKLHUQaOxL3RECeA4WZNWhRwWAT931YMnI
37R7N2KKHoNqjpKk/1NoGVnK6XrJeHJpO/TNybpjxAbrM44KNhsZeXQDmHVcZX8Z
xVzi3st7tEitaMTqCxXWy3q1zFV2JaXzFe1aVbCtOlYd1vT6YZo+9mhUuspCARSP
2Z8kYj3+u+X7HgwUiNL8fh7cMneABPTd42RoYJAy4MjDKSZ/gPKpZm5Kyizjn9w1
war+20XC7GbcET1oZ/0/6PkM2bcDQBr0g1mYrcUb1qQHuIF6Ri6R9d4FVq+P16Kq
4yN0E4BOtfcdQWcndQrgn+r75g9qLVEexlfh7v7JFh4orUrsYZyZKwMLK6c6vW64
lizYwi1NRsD9CaGNc89A91J1DHb6YXVTbZ2d+//B4xlOFaoYqRdU9roVAsi1qzP+
6vEgD4/tlpNQyjv7+cP8vYMlkMHtuNxACzDtm74kQ24eXQZupcPSyaFao/DbvTnZ
3IJqYB3X6gI7wHA8Zf4Fm37KhdV+NEtuBHLLxlybz+FmUhCfn+MnmVj08wFqf5jF
XWWLVvlv2dDLz+lKkWoS5Yjaddko4grQc74NW/0TA+LD9w5dz2t6q8EdHtiyAb0I
TsIIRC9nrK1KH4XyTAblBgDRWNXXSDe1xGS2yRAKv2qEsoHhK0aEtnS0bzbMKzvK
eKJc3u0cIuDoO4c6QPqpMRb1L1J/UTywTmkUgC8FdXn0b9+5ex6n9mTjuR6rUOn5
Ul4aO4/XttpHiVGFG470jsHiQHCeAeDftyoV9G7scga1nql2UDcOUKryYUfT7wz8
4zzt5vM1Rtetotuq2rktXXCI6t4uYHKq7WUvksq1WA1zbt2Stx6V7/u+pjx3rECN
u6/SPCCWDQrG7eDSFa1tzt6tNuOfI3AkNuRrzTgA1NsoZYTc5Io6USbUoCccjGV1
ZtDBoghej5vVfUk2XaT58bh4WJANtcvlN7vH0diWtPHm8flKrNw6lgrAQCiuP2Sc
5NDw/xWMLlh37jUlh2Tp0ysdllh3lB0hJGDY+ItZjFozmtWwmmsvW/jUW3xgFsKW
Ym1JwkmDWZKlqHLdR9wtfFd2/2sn4ma240VDdH2oK8ZCFWkvBbpSp1PcwpqV0afQ
z+yNSvounXfmqTd0ekNo0JpuxtrH0KyYhGlPaFokciRovzJosM9FbLgU6VXUCT5n
e4rUOmKvRTNX6j6zsgNNbgHhRz4Wnuz3N5EZwSAlilfcRa284p9YmkWEcQ8aylIU
e4RCvvuJWijlSqiFwflbNg8g1c+XWMGrR9Y6Yacnql2R5VawJIHopG3PquJ+i9++
Hv2BtcRKAYytxrtqGE9Rvh9oXSHRmoWDCjbthZx20F7dffe3zXDwKODm6SLtqBev
1fwRe2xV+ra+otd+1xCWLwRQOvv1PHo21OxRPSQww2S3Tyd0y2AGafofhjofn0Ft
1coAIUq92s9KgkML61JY5zGmystlmltCwo2Hqip2ThMqB1OmYdiEf3qLoljBN21i
zH3nFtRxGz76UywqWAm6nDRB+XKjclOZhFa6CYfFg/B1gJHAO6xnEjrmTAgsRmFj
aL2Hw4ZYhinI9XJhbQGd1wjFrBGJQ9kNNotd8HivUtKPZfO0yyuos25N6Hh1gnuk
iYW/nYDD8kMJlx4NFMOvnoCVWeHiMgFQdXICPrS2KXYF/WS97xI++7pEmQAtVsVq
rpo4dpDjZk/A5q5sP76zhqGYdTGpPNCdY2PxbBZgqSW24HU3zFCfdTUrgdmr2u+y
/e11Owt4/hmbjU/FDPkFKrusg3wnbzcMA9PvzZh5gUfa84fmkFTNeDmfXDeKpx0k
tcDM23atELwxsVT5s48NKAqM7BtIiGrj9F22vkoxLcyrLSh2C+TTXQb0pciqZqOu
cm+CMinEkIZFL1v/gxMssO/F/EjRUDvM5hTurpEKGX6ZiDQAnQ7/4+PVrsRviJOu
mWNf93iYtg1PFMBF5oschQ+bxKdnJ4DgUFGxNFUhcL55YK5aJn8ouD0yJwNo5xID
5YCgczlTT0tyLm8DOwYoMYeztZWM0m7+2dpsBAuUu5X5BUOuvJ1qCGMvQDIcjJYT
PLZsltuutL6vOZDzzccXlbJOcwjTGcocmbDdW/TV4OqyMGRhrvz6FoVH8k0Z/Qjn
nglMp26EcxGDIqMrRecL2lji7R42y0gn3KjcJhltYXYVFHF7DzDmgPPt9Fy3FfpH
a1MIhEvRDPpGGzIM1fpnXjqUWDtybJDDG7RBup+iGkvA3FKszG9kkwc9yjCRIwiT
uHYjibRus/mGBjfrfAoQpl06cypYqbIFqTsrRXu1BlryydrDw9ftIz3cZJ/VC6t+
b5Wfw7HWw8/ob52VuxajFexdiX96x6sAV7JWzmgTH++wC9gsJ2yh7cvU2RwtoSdf
JPFt0sweUQy577RzW+Wa+hkwRUGzDVvn6iJ+O8wWfzm5EXU/4HV6naxLIS1JRHDH
D2aB0/tknjiepMYcQMjqK1vDbrLGuY+M5UbW3iuqiLh2FDGBmdvV67LdCBhiCyeG
f7fT3rXxMXgHokolAmtN9Xz5eFk9wlXaFiZ+DXZg13kE/YCbsT2MXlhimcqJid05
AhqQGOrn/XO0x5iny0XtpkQFDRL2quLs+UZYFldjflzVJZA6O90ht6MEC+OoLTJ3
oloFtXBtw3f9SzsvFFeLJABaWfFow3ZVqLkVNw0fmOrJf0K65P/o10gOj2l53x92
6zz6CqKcWVis86ugjqh6eF7tKVbycqy+FAMVnU109Io24++3OHOkC9Fg5hW0L3ny
w2fHtkAW1Pb28jR+QQfaaLNbap9GEMtZ0VFvxR/joipNoZJ7iQ1oWOtfGnO+6b+X
tWK13f2fUDQLojteeKji7DRtJG2sfnWLfXi4a+i6R02ej0F/+6g68Xnpow5hB7jP
Njic9i5+CIPQ+1+fELkXLJ/EVM/liwdE1MQgcdZouzy1MSDhZkZMpkbqEfZl9j6G
7ULBCRLYw/uLYQM/FEaaR9YUg0vvZssejpEPUGu+eYGLqpELE3UsOWSwsOppCO3J
W85LGHY8bshApALCjd32Yu7fL66afAUpSfyFOORimVl9viTD+bEh0gu4dhleENyB
bFgNBsut/RP/gxf1WWitRzCIQhJFo3skR+nl6ph7CsNHko+tS9+vQWyeEXKr9pbs
FPXcIkLIGRjx79NMRqF6Reai3KZx44gTW3ZH1F0rKR7wY0jvTIeEKbBY59wCrv/0
ezkyk1oP49pRTvIhEr2mdH6XViExq9K1Z39Tg53E3R+43rFunvtZx6zwdpsrLu52
vXBWneFgwag1+YKJkSXS07WTmyHFnvIs95WFG89+SPgv11HpR6wVNWz8IXUkP7MI
VS/qgSCIwz8Z3ixAkns3i7giyAGN6NnRYSTlgrHxTB5cIN6wNMjFGLit3c2oT+14
3nSW5afrT9yFirJKSHJTMRn+Jj9lkDNcDURk790Mq28UaHvgWiuNTqop87DGlEMp
P8a638I+2LL95NYWxq5ObsK6zrW5b01Dg/1aS74LfzulKEizyrWJmYCLSlke1fCi
cHhxARJ6sLrAebEpGXZhhSohHUTAVmp9lBmNBpolLGBNX7dLQmhpWCBzazJ9RsdA
JRNkpHT3i2zh0S6Tc3fUZ3+ezat3WRO6ijeSY6tn6OKwV1hHjzUDC4ItqQY/zJ1P
Z+xHERu2B+BKNZ41bU1dFUFO5mJNQh8ISEjWrISzm0o5wmMern76AVq8F72/Aitm
K1j1iw9dRTz+O9D6Ttkz5Be5WaN76xQlfb4zKHfsYHmep/bb7dZR3c716sYEFn4P
tQcgyoEqNeYJhmuzHZcj37cq1mze/Y270g60Qo4mG1qg5VgmGTAleMwamtPRdVZe
fSFqz+qN/7rUfSf5Xmoy3XO7p+bUppz55vOBB0C+eZ1DQ3d7duj03n5hkUKwXHYo
ZixN3V/ITbdqsG5sNttXN49cKsmfTy8TwIv/0fXkPtvx5+mQgbQGqW0eMg57GQ2P
pkDRPKbXLUYAKAnXe4p9KbJKneGP5G9EXjoUa6W7odv2RA94p74mRRao/Z61phf+
WBVDlnUQEqDJCm7coAlkDYEcRwmXREtGuNvkb6mgsGgQX+t9iIUw/UhaNq0C1dLo
Xd85arJf6n7GSxi3VZJZn6J67Xy5lRM6Bm8caX8Hz3KGXztLNOoqTh1DThJ6V14Z
4Fi8nAuWWVurxruMhbYEcn6v+I31dTXkhLCNetd6KNKLphTRh3Yjf6V2wr0kXPBt
re9yHdUlbbms45XImyVKsepeK8NIWdiH04S7YqlPx2m/hQswYQ22PHcpzGt8gRCo
nndttMenzR9K2VVUgayqb+btswjOp3ITdZW8HW1IXUHayDgqtLU+vClatv6VZusv
iKDtQcZQQnXC5noswifhe2btAlWZlNAAJvzszPlDU5RbnKUw2Wh6raD0IRzgcM4X
Crm2F3loLtrPAHjOwDhjZS4SnRtqVpRef5aXmmlLWSRkcz4MLlng2EyBX1w7cwZV
MOnDiaCcQA/F4uwa86OpO4MQANz34Dc+6yDIx34VJOaBN5BEB1VVo2Q/yAUKwCcW
JcoiqrkLzvME8pgR2nt2HsnBzLdSYgYNBoFEeqc8vo5wIz4hneB4bgLp8/8P5pko
BAe53UYuPQ+a97fB/0WRvquFvVMxT9jzeYIvEbIx4Iz5+ZI+0aX3q0wwEu5zFeNG
D7f2rvgg8o+orHfUbm0QrJq4iPeDL5OIb4NOzJjy5/CmhT6gRhxuWxA6W817DPNL
Q5ufsZxjb08SamHUx/jDQbRV1rB3qhW3B6YFcYJPer9eeGvOawLH/Lt8ZJuA6PaD
fNf2YJ2sWVi3WlTy4HONsapacVIg6Cr9W4KcPpZiUKEiNwT2pFKuRyxP3yZJUJeB
0fEB487ZYRA6zdxUem7k23fz3A7RszeCuZRJ6SlofOZXsYviqbuR5SwJ2m5usUGb
FnkrX4brdOT2DN4Rirphw5bNMUxlVha2j5TMy2BaF2y7fGNIwGptBUXtrM6On/7D
S8KDzNdAJvWEhWZ7iS59+x/jCusVTcDy6lKqrHrCKmaiVpVK191LZ/6sOoXGEAPZ
fq4ahJiiKxycquxEyK1qreDU4AfUPhCkcoGmIK/Gmtmb75BzmyhvL0Tvxj6AvecY
nll7GEOnvaehtHZICHrEnpTGxCPN35Sr9zD0XNMb1iCuXfLwub0islTHnrrz50kb
HjuoU6oyQhIr6iHT4wI6RAXIr1lIPvr9mgYIqhfQxpJgixuhYx43W5DLLZJJn29Z
04q37odrmZ+BjPC9zDb1/IWPDnWe+5biH2TjYTdFIrF3ZotIel+qj/6spOEhFH6n
fU1FKRoGmwcJPLgzd57hWogVP1ALf+GogkDWcHDtiNz7J8OuuSQZPx6XT1wGN5Wx
Z/knyInYaAT4NKwFwHl2go9TT62lO3KEdXWMrxkOUFgKN6WE+KhR1HiIS6rVvRSv
uZ4MGzS/JxNj4wcymzzdlWOaU0lKR2rNvdX3aED4in8M1PPM9zync6pGGlCMbIKx
xojgcV5xVsUe2eh/f90Pm48oanhnw9efQXEMCbPcixoZrJvilx1bzdPo/PqUEIh2
p925h81PKOnRu1tIKQ3ry2/l76scsuCTu5wz2XRuf/lrJpwO8me0cVQKvg+VM/B7
JmiJ7nLt8o7BYfNOPSM8e/YKK46Gs8WG5q4o+B8Yg91EnMMUPEkngVdiEAcO4Slk
W1ao+rMOGpiRRPQLTr53/l9Q65g4ekpoDUaY3bwHl0VLMtXjk/q7njP4Ag3rAmZk
t6PO/HpfSgr+N5eIsLe0YM38IfwoZJnAKo/2zvwuYiC7dI3QXaT92piXdFJkSPvB
1GuMTGoHDMD6gYG7OMf3+9LS4/+q+iwhAcLB+bBgCPZ2gY1cvO4w2vwC28IK3KqE
Sheg+pNCL0JiluSPk6aIH/yvPZ3GX8k3UKegMfGUSkXMdF7Wm2k41GguFjZxROmf
jJ/Q5E7QuIIPl6ltIyNP9sKI4q6+LwyOo4TYFF87bFRCmvSLdEPN8FLABG0feQZG
BpepB6sbts/Dnm5M43YwsO1igOM89O9VLl2pUAQjmkdYnUnIFWtwQRRvK28l16uE
kBJi8rvAcgA9HzzbF8qMxnzIe3QgppSnaxANHNCz96ejZCtn0zTl3EIgGzI8kMt6
tk9ngebX14KZgAo+seFYBJ2jV8a3oAAr0lNpVwRvR5mbsLhRyHUR1KWB0x4xSMbW
/iZ13l9poS7WuITFjUT+BHrM6YhdDTStWvrZyBHNSojPDODWe5nzcKuHZYnyZzBM
Ef5YYz/2LZ1mtkHqJU2YITFcyDxe9VEXDAXtJLHS0GkmhHaGzswgZqT5kC6FWxwo
MBnT7h53oPOXskYrNtw5WgdtnsNWYVniSe5sqaVLmwQ4cMHD0AJn5gWGGS0dwlhJ
6l72g1PtX4rqUdPTAXKLl/DAQq7Y/RB2zL7wwToSfPflxfMMSFtPqcOHzf8j63oV
WxF8t3zMYxMXdV60AZ6G2uSRiuMZPRxb9yFUvFsjWLy1s9N5PkXniDflnHS/FtKo
9ya366wBwvY09IUE67ezO0gftEdc/z/QHbeEwR1D4sABQ6bIZhsQndyPJiV+MioO
Kbbu+511Z1/bgHDDfBXaCCIyhbPp0cJUi5gqb1HNaigsO3h/oo+6QE2sj/n4Sz/H
RLCG9YSzubw3c1emktJskQ3h4dwkuE09Q3kNMwr2SkAmKw/Q72Xjfoj0BDPy4/d/
wKmF3mi9VRCIJqein7QGbuO5++/HAhYI8jDHDApiOuXl1OAHXTYcRJfUJ1sv9UIx
GWVR+mqOL/wmxNu2p/wv/3a/u/GnvHm+Izb9ttK9DtIrd2+yYgQftPUtR0Mq7UET
cHmxRJsZU4YmLdchecsUjQNqscCyucS4NrGrvBcC/FnL49IKdR6Nmehs4zQy/mUt
/ucxdsanEKaG1vlPAS5sxv3zMDJyOPkIkhQPsLja+AaGPwkHIHs0RSbStWZIvMse
7edgdNDFCaUT7mJyYNwJfuGZAcaozCnyB13m84cUmUFAI1uqGd374S0hLopn6ukP
nPLUbRmdUwupMFboQWCb9B/7PDOFdwn6FTrnPjRJBGIhJWY1Mp1OuB6HUXjvfwKz
KBe71q4UL1xuVwPDKEVx/dLffWnC7AOeSfdY7/GeGita9qJdg02Y24sJqIyS6Y0b
IHOQkqLoaIE7isF40UH6vQoQAXDsUP1zwOt6/BhSoazX1MYhqiCqlsHgIv5b57kk
nEjnEp4ecHNtBKgWsqs2SXblI/4orPcADwtRQ+oJskgc9ifcGCbCJLijELHYtexi
KQhOA1suQNI8cgco8+j4vDI1oZTh77xRaW3mkkBu8MpiAG6qNSO6FR68b1KdEVZr
rviWtswuoIGicdITBUzoyWkmDnp8nb4gO2lFBoOgfscthjTNzlR90tJ8ORuIIqFJ
N9K6zoujGZ/kW+amxyuAadBcjasp/IQ1eLMptoJgFdimw7lYmdJHRRTePphVV5TT
bRG6rY9MHxL6f1sE1x4boIS1uEiXShO8FKEayNJhfaEKYLAqpX/R/NzZXODQ2Qna
pfaOdloNyYTewsPWp067SHF0R5Ss4nqU9vWX/24qSTvIQvDG4BKg7nKmTRKVvGCE
Ord/b44lp3fHdIPJH4Zp/uQ2kHP4ZJjB9oXExRL2MucrccbsyozTP2h5TUeVInKf
H/+n6CyTa3QqcbDc7rXrx9lk1fBCJpnEqKUTLmoZ8sylPLxvdKx7kmG3AVFi9zeA
WJuv6TACUAhdpkTUDG3WMKYMMihH7xj3R53cV+yChkMwC8Kdj6jOEPfzhPdEf+cg
fd2GbXtbGbg9Ba6t1ZJ0dGxuW4AOOY+aU6zDHSalIHlGXdvizCUxC3eIVMS45MYj
jl/U87kYmgimqM37EsbbTXXQCuzqKGLyOX6ULIouMxBmIpZM8Cdz//R3uiBOVlDC
A9oROmKNUR9s/XU3qDqDHL/qyElphZ4zIdjO0vpLylNeEwHLDOYo84f1t38tHEuY
LFwv+2SlpNUcuHB2HYRYFwf2sJLsnJVLlvkco3YdYTLhMz/1+h3/jYeZ7f7p2f9d
zOjBSHFuHBE6EkWnF8eK19ZiyPtnCf3pn2DWh4mlgxBpiw7Jk7YVTRoJxswTamYv
jtgZ3BMqMhDL/9yY/ZR+E+AhOftZ3u2WGPU5RiV0pnglZihEXtWXq/FtWOADyhAN
0m6MOOg7mZbrn7FcXZbqmAx/q7tnNsdGrshA2sDVubNri4UD3cbubP4h/p3aS26e
MOU/rTk5sSxq0ckgXi6xdvlF5LUpkmjMnvy/vgVrVDQ3BsLvVushpJ9LjCLDp17D
/WcTSunci7fbBmuLbkah7hnM2rZ9DTW52pjFi56DZjGPPVYlxNCttJfrdTAzgImH
MCQ0WUn6mL+9vqeCf61apcOV01+hn5OIGtJ5FkwGsSYRjnZVE+W9oHc2Rp9G85sW
0F2G0glFfRD8kVu91C3NeVA4Vc89J4DvbTEO6RXWuq5eWFQH+JYDHpRR72bsPy7w
Mlht3GnnSIXYWT96q42aQpA0gUaGxVksbvn/Or13z+v8r+3KnLQZpe2SLHUKSjlL
tE4BTJBpEgXUyNiyhmSFfdVBgLYVMLx0nR5WjuTPodofBLFssZhy7oQEH0icBG5k
0XcXZEIVPcAfeuFYlkTT6B7fd1l3AOiHuWiRHpXQbfPB9iRAqVjf6iGluxpmRXvE
s/lZ1+KTC137Gd1Ue/bPpCJwlU1aQSRS24/ou0Mpz6i4T4oc8+FxjgXSzFTB4KlI
M2O4l3njZvKx9g9Te3LXtbf/QF1cajV0QizhJpPx1Pqetlq7hSJ0j8cK0y9ZYMTQ
Woj5DOEV3AHad3lKwSrHJC3ZongMir18rfIUW7vbStzYB/WRcbtjkTqeioRnMZ0u
O66cFVVfpeLCs1BIbRMvXu4M/3L4k/PbTweojPjFjOYM6qsKymGDeOyQ8byn7ZBy
8nrHUZCnGzHcm0iOBm7GE65CoC1kF6nst70k4tnnJ/+zNg+tN4Ohs4EETigo6Z/j
3gjS77JzJd5vIlHYEbwPj09riBvyd/HoTJdL1SZal4pgJOb4qsQwPQQTsNk0Mujr
sogRzl06/QEzW3MnxuttKeWheugFo1hfrgrKhWRSUv7Py0qbECJNa7Fin1ZgdmfC
eu8yl4MNYSgd1d8a+nNQFaIvjhRIcU5lWqqplBRYwQbj69BSxwzd0UsTqOmax6LD
7kXTY+xOLJt/SJ+KOl46XDDJRW2eeEPP/893dIpwJoUZt6wCLb1maSzpMV+OOzIp
aDkD5XJJCJog4/S3qWBF6BaiRd2cGtBl01Fr/I8EYANAXDG3ML3xIGHqH8aE5les
jGrd778UfPAfZQuumfuSp9+Yz5tyKrwYggC4DNfcp33gnxe6LmHJSZx2CpwH6qJC
3aKaOZMNsaCkKdVBkCfv3o0h0uuBLDGCHuw4d1YTcxQQHsfqlpFvRJGx0XWVWdyM
bK9JYqgmcx2ynzUYegafZbD0S7MAayx53L8z6nhEsPuehHHYdMvt7FrIoZ4RVVjg
d6QqQXsPmzSHlG4A+wlHYlJYv+ZX3MQL7tQ5pzToqcXYvkRnLsv4UY31qurxawcF
jxJzrSpf9sJad/Tvu1T7TUzok36vLgstLKMiQrfuhv8b/tbrb/QakcwHizPlAHwH
MHVtmm3Ev4Ge7mprxkwxEJV2JW5PW3doaoFdtZsNHpuQZyfawZ6XXnOK9dgE5F/D
4Ffzv1D8TDR6IpFEsii+EXBwqVnCvyooERxPIsA/jDncSsjDOBMB0s1vZU20FQc2
AQlI37Fi6hSUoRvoRrm3cmSG1GB8gjwgRtKlRdTB/HHHpxHP+2T7DTOWcYBlabuv
LB0Ihw0URkmOEsFehh5LKH0OLBCwhe86zHiWYwNdiIcn59bpJzVTHc0f5SYaqCc9
FIXt9Pi/5NKz9xuaRCkU/SvB9CVAOAJCEelJCn0jzK/rJixAlqPau1Qt1qQTqjvy
xnAHSkyu1uUqPWPXlXEYGOrljjYZeRdithjaC57rqyUfhRI0TR/hvTBCn+Uyo45P
5sGOHG9oU6R1U4O62hsosZzevXRK9YaSuHwjgJJbuUijAh2WVDWrP/as6BmauyM/
LE4zDMgzDuBjif3IYVuHukCgxKhRwC6Ad3ByXNVabGHklvHznwh8UsnXvjI1N28K
DakXbmm2iZlwnZoIN96vlK8LHJRCWThOA52/NQwKVfoOIjhSMoYnLMAQBSlyyHWL
d0zL65VmFR1pJQAKlf06Hm3xHecwk4SQSI5M5s8dzCxVdWtMd5rMB1NIRQs+4qYF
O0qSJjJs/NqkOo53bYsUCcWIncBA8jDl0UHQGHaqySHgLuVXTAd2rYLcZW66T0v2
4uW/MoufM73sZrtDM71ZtnNUn4oNxufXfuK5SqVVGgA5Yvnzt2J1TO7McjU2II7i
tJgQvUOcmBLQ3tgL2A5QH+lxrVjgIEsce0GXi+SAPzauXrkynPT2+P5fA0p0VKGv
Xa1purP8xXhU1CIyM1Z/dnC9eCtAN66P8RopqIha2rEEJyTd2asiLLluFVB6dmfk
4npVL9gYfpfbb6ucKWEOAhdU3hdnO0MmAVjszqcxqNS2+sk3lFsybQtTcOsJOww6
wR9Gnu7Fh1gW7uMubt3/6I8v3uWJv4aSruDtZzaVI8XPq2/sdZ7CCE+jLSzxbiOD
3646mRNbuntzOoGNlQMkBGfOPRvgp+/XxDHqDlhSR6piRMg7+ZmYf6o6x1inOUWC
ovdJF7G0umCRXC1OR/5WtU98ArqYnfspNuMsJuYpsAlQVc34GHRZUV5VuVCGOO2M
m9mpxJBeVT1GXJ4TvK5KoK84XM1OAnnohEWe1XYvpqQhk8EtEGTk7evPzVViIk+M
uNBnGQ5kwKsjRJ4uYBbtUS528O5bvY+L5lv/FP8Qq6k0fspj2JzJxBRJbTFNORQ8
hM3hcjJ8aq016vEkKC5DnTlShgZ64+K3fvY5Zfxm5CLqwLZRZsmka/75g012E0fu
zlc8RJyuXGduhn93zrfOBUEQ37qcihYcawCabB2Uqjc5xJUuQk34133RLgJ8DVsh
Hdqzus6HVgrEQrISPQsseSA+yx50NHWmvR795yFH/cO5rTAyqB4miYDrJYcxC5f3
bjkRx6wX381LfMm73DQBeO34Njt0AmFJymQSx/3NGqWGzBuxvM0pd6Kw1gPHhJ9t
PEYZmCypDAoK//4TmOl5o9BlTlRhV+FuhckhZvTf01kuOp66kXEGnMuD1GJpv2Gl
DWZUvoRf82DsQSSRyrfjOBG+k4ywxcPa2C9R4WNnH7U+tFD+XUOVPe7pWQiLmQGe
AkS0jBlT6d7d9iI8i9uFd2MvvfnAKsv8MIBdla6m8dSKoNp6YHtyMKrj1toiZDSq
UHR9aZA+0pkg/lm4BSpbsjbMB/BgaJh43i0mY3iarxm7xyhINktq0s3JAGdLsfg3
FVzSr+Hx6fSN4vWntilAez/NK1pKeTeRE00lEROymtc9QHt+8icXAhA3kPCBzsy2
+FCjdk8sCuAlKsgd1BnsQhIzrRYIE9AViTG7lLyfSwRgTZLMFIFprgclqvPQXwtS
YTVT2mHfl0x+HLRIO0I2ePygc0WsqZe6BR/yRqQun43eHSwAUQs2AAnT/3X2ix0P
Pgt6mKy66Tsa/KmrN3nOBOY9uzHYaHNk6QPIdv7rnn5d0GeajYHK+CE/BSJ55pN2
yM9RbvP+9j+rnFWk4/s5RxrTSVKaz8TvosjvDsxX6iyRl0H3kgnEwti4aKOapZwr
rTS3RGt2Eo4K+5/7FM5rXYUS4z83GCFQd8VoEZyt702PvZ4Skj7QuOZYTsgVIZjn
ipmu/zjM5CA2fGJW4IoWm5s+nCamt0DiMOaliqxCrVHfML5arvNQTpEuKHJQbgxv
f0c6vQ0P5MPYLiNFRP6njcbtw03LwsW3UiTLGVtXdC23K2hzkhvBVYzrjgZ6FG5e
lQ98bQ/atZWH7ubYVvIn0ZG3SOXtZn4TlOsoT91QFOH1ku6PPSGtRgkM7Gxp7J9a
u0Zo5IjR5jjktWFYNoImQ3mhJqHpicgwCbsN+HSf+yWAielzuQLRsgT7X3CKAhiQ
jfQnGllXv7WD/loxlDSX++CDqxgyUZYuDzkvz2T30TvjCtw/1SBSBH6S+nJGSEvu
C8ENayjqWx93w8loVr5ZCx+7Gko7JIRbVUL4U0TXlro4oH2LgxryhMYgPkUfRyvz
MepDtMJZTGfqWMA6GWeocsHCKoOF+bJjNxKpgshr7Wz5+cdGObbJHoRXmY6MKIO6
QJ/5K1FopbgN4SfZSawLxB5BoInAxpSr/oDezM5NcOTFzyJ2SzHqwJrw9bms+yfB
e6zKeKZp/u9/RTDEeWglz9sHO+v7i9Lu8IbA1DktXAd7OPypxV4gfPI8ce2PyKUP
R2cM1a9K/xGpIZ4Tt6QOkivKC+A+1Ob8ATZKqGJ5KRLoJYQbWT1A6A2Vn2a2XHBk
IeodzM9QtbNpaKKzQh/cvniM3f3kzb3Vv5DdIaXYKcWMm0jsgJTa3uVbaQJsnA+R
oVYQiKEGcT38UO75mMJil8RKUSiRhXYLEGx/5Jj5nMBnpJiJX90xnR4fcP8dJOez
LhQbVWpXRWwKz/tWWDojijUdWi6RhnFZ/wMF6SzSMrF3cbZxKpBpO+FbZ7QjdsfE
lRAERv4VxDrPYOcJ02uUiWE49yBMW9JmKYXC6LfVcoCTiWwWW+tiOMz2+7nvIgJG
aJb696qlYcfw6fPbMQHwkQjBukFXjHcKMR+NYvApSdVsj20TSBDl9l2yqvK78K5q
yLk7V9B8Y+P+I6xrZvOLY0FeORuKAffRSo+hwIshEBgcF27Tad23mOoP4KRdIIg9
fyViBzQWg4NcAHDiMAIp01SBNzdKuahbauaJ4vqY5ySvIkBgxaeFgjufEGXXBACK
5FYUnyyYY5lhGnEoRKfwY2ojfqtf/Jd5kDpeW3lQ56UdSvXC2fXJfln64tk5Z+cc
OJeeq4aV+TI9RcYrXCPXS7zcnf6RspbdBQjcOYIY8FtFKo2fpJfdS1fq4aix6jeh
qShlc93UcMzJTl5hSAlJ4fodO6UHQbygPp3onaLHx5XBQjj3dKEDf5aYKGYiyAKs
25+r2xlYF123PCuZ4WOxJTwxXhrIJAGiL9kokv3gL9KMNnEuKscniLiXiN11POf8
zRKjMoshg5nxgSChzPUmnazTTj0x2YPQI6PK/1zQluPSHM987lLw0Fx5/lbuRwKJ
3RafpCPn3G8STIpLezYUyE4PEuAvQaDkCovboVVun36OG6L75WgzKggZjrhZu3dj
ReJt74GeLrvei0oAu3Sfz+DYp7aOIIuXgGPTJV6juQn3H29oR6bG16Q9ugEX00u0
s0Oj/wPBC7Hq5K0GlcC9aFajP9sLbA18b2PNqL6Uh1miIQsEEoEvpc8yR1EkUBdV
vmcDWfz4jvMj0NWfUYOftEgvZMZBzUxFOpwVW0M+Vaf5nnc3ZcUZOFoOV1HM9MVo
+931WRiolEFRsa23shYjW0woPMYlETXEfHtPITz4tC8XrvkKB9K4AS+kXXriow4P
aoxkkyxwoDDfCGsuzsFOF4cEl3zrAq1vwq6ruKZvakl7dDTlF2HzNqrVrOrBQ3RO
+xyklpTEduVpq4Ebl/XvrWTNxFZnAR5GdxFpoa5xmT9UZ/CDRkFhAB1eqq0BIeQs
Li1+6o+iNLJUmnlL9WRcM0LqtO7ctsrog6+0Tw0cOxor2oBbrd3I5QxhVU4ccQrH
8BeCyNEaMCtlliTgJLEDQmUik2J5R71pzCTijuU6wwx9tt4ESb0KKqPusZyvDMwo
7pa1z5rN4bdazA0IFfc2qqKccHAzOe4me/daTggmc/XVRL2NE8eORGoQQlbWbDPv
DX7FWJv0TQQnhE1yzp0nO7WVNHwwoiwKhJXYTS9ZhU254zg16wjKcrh+hfjWUYFQ
4KXdstJWgIO74ZgeMOENcgo6KDViDlEEs+eISDNDNrsE4lHY95akiNQzcDJuuME6
K60jzELlmn4sIBW0cH4QwVJc1KzLq1Uq0RruEVaODtbJnoeuykEfDP66pO+Q5xMB
zUZmycbJVr0/tkmWTtJjQeVGenyhJd4x3x0YsnYJjvkOMVERDo3p1KTM6eVJkd/2
ooUQpv8GLE9BmNILnzOErhR9BWBtsxAIr1vS5Nu1Pk+Xa7amFjEd2xKxTbPBngFt
GSt/XQ/ysaze/TQ/XQPodcWICqqTs1nuSIx88VZRsiN/RSifTeqAMja3H1jTswwf
gcLpiqO9N1NQcqiWi/JY4/ovXi2RQ4y5SkHvICq1qtPhdLR0vdd9bVpdO/aphuas
FjPp6BdlFrKt6LligPueOJTmWMMjvnps9icXbnnJOduaT05wwsroT2sWdwvLJhvn
h0wk6QnagIZBZDdPdc60gdC+78Io8VQ9RBr4c7XUvoEy9chgSkJC6Fray84v+C6+
QlDyQTkJetqtdfOez8xlZ0WcFh+VGBt8Jyv05kzz340B43kS5Jjb10+AIUHUOptU
ZVFoDe215sraMErLnRua2LKsfFrPnKhAVNQksJLslyqOk/pKmx5jxd/Q0zwcKKQI
vnXyGHCgC3dJM6RNzFsC5sJWOsKJFs7ff/Q1TWETEK1k7v3F4MN3E7woDdH4LcV0
1EVS50Y6vOA1WwZ6jZaAxMPcI+c7eCyGHn67T8Sgml6Ad6QtQFcCPjfg3mgK8HyE
pZQoSEf4pBW1WacVGRr+ntkuXvAiLzqvTmeZnsZMP4RvEeN+ABxMU3/srhOAI/Br
CoYRwZACmxaXwHwiAOxkywwoPKw580jQfBv7a74m2+v7uxoxOqtI7xUVfFed8AQO
LbNwgNbD9Kbu7PKeWGhEyXYRp1VjX7d+i7+eF3f+GeAuZwC+xD5fCwhJPElGsTAs
GzwwxMC47qRkUEIWodc8QQMeE31+OcFHCPyHwB+T4yeYNdMnfA2L5nZ/WS6Kv7Qc
EiAYPeBiDsPWptGsktwgGh38vKlOS44glS8D8u1B0V0GU6is5vz4nW1XJxdJ0OqM
G8CDVu96klCZCgiA4mt1Y2kmLO0K9/Hb7PoJeUVtOa7xtRr5eEkojWbkFPsLHE9C
oqHNH8tb1TWn53pHH9P6rTY3Cb77UMWolyZ9veu6asxKj4f8PSKmPixr2VLC12lT
CZ/dMxQzGYyjmJCHWaMZu3ICvbFF4HV+mZWQ8OLk7LJ7zWR+vi/LFLySNHjcM1ke
IgDrkU7FCn4/Jzo3XG8qmI2yhqxmj1asyzcr+BuZJTE2fEFpQFaMmECFprTnJL8D
uXWzGCjPIOSzNJrZcBPqsH4XKiUHfBL6MPIYCa96FPwqBpaEW1GREHPlCrsVQDlZ
foVPsBnBsW7BXUrm4avfUEClzVM4n7TM1QRW03uVPAbe1INkchj0ZDgFg7XH48Wx
ijjJBqgGip070grhE10GQzlj3J1ARbQ6TpZGNWOLLvXgQc6Yz9ed9opE8VgE+ubp
fbbBXI78E/jTlf6UsKNd1IOpVPhdzaOE+Ue6RJc3nhqswYbdvv4FyXZAbPKjyoy8
yTJCQUpDjchqgk5CDNJnjJwVF9JKTeAjyhSWVB4KCFzVHHcTxlYnVUbKyb/t9BHq
qO3NsnVeQIYPyTNhC5PB+a0L0T2D1XyW2SgFI6527qS+djHExGO+c8YvLTsxUNFd
nYhuqVKm3gHBPj0z5HuFUbkDbLjmpRHUV3X9tqik6rovP0S2O78+alAfAfts4QwC
UME4mC93DUwVhNSt0Iv0FiDcW53oECcmIZjuPZ/R4LeH4mEvI3r/vjuX5JXTs6/u
COenQjPk7v4z04JPnc7HBMLtMugqxT48+PMAMWt1Gt6efd1WFgqaITlmpcMZJng5
m1xg/WqJNHhF/GZq8Mq/HAgNu4H7N6vtnPRZNKU30D36msG9D36gMzxXokTGDg8D
PwzfnXSLvYlSADBihmbQZB2qlpm5tw7hW+Cujt8L+fuVCOE6lA8XGYfIQ92hCY//
NX2hbPZ/ARP95UJZyMCetCojOUY9gdrzYuRGvWp27t3Q33qEKFsCUcu6myUhBE8Q
PP/kAj5KCFzUC2MdQEf4cxkFvC/nYCp9MgwqOv+k924TZH4DASVHoUUv/k1kpzmB
t6y/DJ0r5IuyG3NJt7Wumq7h0Nn0f4HCmC5gpgrOQk7D84o+3gnW2O8G2RCGJsmO
4pUDzIKmugJdRyI60HkAFxg8tFb5bXkr6y3GwX7V8pkZ3kaFlyQIiOApiOKaruWU
KuhVWxX7DMiHtwgPI5olPKT+qAWdWn+W5VU8F5qngu/umuagwU7Jo12T7IRl0Wj0
KaQsPck9tmZxriE7F1dN6PjON86tw6EToUwIeAn+i8sRJKFwOKzU1I3BiZnDKx8/
ZlgnN/pqANK1jhMnJDgo5T4rjG7VWtt+9EvxHO2wLrCa3X1B26X6HPrwmbnzEQWT
JB7RSR2UaC6AfccFjRM7r7P5eI9HyHTzT4hz4OmOKzaA7wS63T7Axdg1tVowsAfp
yhzbC/aaxyQNM6ZGC3w4fAurzGOqIvh/XFXMGJwR8AgwacqZrMA65i7L0JSrJY++
Pcz7yOoehlJiDPdmMQ5I/q47sb8RrPyBYXovtqCxles0X4ED69UEg6TNvBA1TxZJ
QOfD57PNfRTL6OZuXpWWXu0QNcO/jHVXLoL37NhbTe7TlsIugbsE9Zd2Nr4VMOH8
0AW/0Fz1yOhpsI8n6W2RZ3SnD35yhwX8NGQDkXKx9W1FDrqyjZAuzxF5igO9KVVw
B3zTXWTx8SwpeNg2mCuocdTYslqnScV2C8j2JUNL1hBx9IGaLKhQs50Ki8J2x8Mv
3UqBRKMqoE7sbVe/03c5aT/YBgKoimDpYg4yToEyxH7Ab6lBaNxjXJ1QWBsEjkha
ii2ieuiWvonycaRYA9mmLYz5qR7djS2pO3/m5yYpSsLh6IXh0iHTuN4qP63B4H8l
AilMf94iFQdOkhyHUui7FWdq6+epc+nM0Mqi036vhP80ge+tiLdpTGFTyUnyI6sZ
kQlqpon/JL+jJwI0qrW7YqzPAQHy6i0FaPcTOp5UwKf5LsZR6gjTxcq+0JguvBqZ
cQ64baJXhrY7t5kBn5LObV/n9nCHVWHZdtI3hQoVrvWYcZnwjdGtLGnfDlLpyx7s
RDemylu8s65F37PWiAwpzB87wZ0ZztfmoMNX5s/WKf9y4x/0hJ5jInH6cJpONFuw
I4VOamxOW6jGiq0JhaZvpvuCASK1niVxhbLGZgWEYKwvwuSWWDqeOubWRDe6+2f7
Wg6MInXXWONVdN4JC6fe1vK7L1JhI0oJgkxv4JDSKv6UnIk9d4yfYdeTciMIDo7T
Wu27IH8ktHKqKTdD87vnG7RxxMyd50AeLvZvNHvtmW0G/vxm4aC1YxJPqtkHZUCb
iteHkesg1/m4jipEb2uHEQDo92ujeFtplNCnQJxukYnluNGambaXdjU8my2hM8Ct
h+6NfPy/jtlJH+jgOYX9q9Ib5kr7OQh063lN9LRk4Y1JHPwuLa85Xtvt3qRvdRVx
IKVqTEBtEuihqlSR5NU+i8Xz2xAKi3VcNLpzcuN6bWWLretKdey06uxJcdq6hZ0o
XZCvpAn7hhUeLYtCxESnkubf4afA64FGCKf128wevalU9Uw1Dkw82Qh5FCFJLJGY
+N3HrA/Pg9mjTLLSgzI5V8s0P8UXEIbT2nngCSqBckcUQ9IuMcK8QD07ohH1QAIT
hGs3jSKIZ4VxSZhRh3y8/tV31z93Hla7gjFGOOSuImJu3G5eDlfg4kWdVmIpCpzk
tLkmSotU8OPBd7w6V9t/Qj2Hz000cFqda2UhJGzLI2JZx9Q2krVeG++IKad2ajIL
eIbkRhoQwbL/pjtPlmg7SHlLOnOFk+igvv1TbSt5Gc5oU57O1MYCUjcLa/b3eqya
FZLR6LjS2jwFaaFfCQkURS+E/qW4ekxrvZMzn9Mzuo7CoKMejMpa4moisMVyitww
fdi1LIRGDl+MZZSqqeaXUNtt6FsX+DdqwqgZdytOw+o5gdXRjU6SQp52ql6/I3Xz
tJTHF4xKeqfo1LMtzoese1pQ2NElD0/plZW6FTlNfLpnhLRhNWRX8KkQBoADKErV
5se0uyAvELEeENB4ze4XRl6OU9Bu2jFtSFQwbCkOAUI5tE5jnKwiW6s0qlm4GPQy
QY/CmhboHb56xdv0pMtx7yNZ546jj5zIgFDG2ZhhZd4zfeJeBFkpQdT3QlIjoYrd
XEka1XJU0J56hhirNdxBIGXIWPujTvSpWQl0+xeAE+vULxlzl2aB3fm9PwdSqerk
4hyzN8LYIlmfOHLEMmSrJ0oe93rfje7v/+jphqMqx4jN9O0jY4akRKdMTUbjq0Ed
h3My356RhSBRTQmB6y+Ngio0rTB5+lf8BHKuJe2jCZrczx2HDAoYl35Z10w9d1/4
xTswIxCGiJsqrEE0R3xcviVx5RAo1KFP3pkK/ugrG35U412XgwVG1FjaUBHlBRe0
qefh1HJVY+wHq9BcdB3YYLp5bWrkXMEwpE3x9/hx66/KQUyuyZHTVBkhIixZu1gj
XcJ53fKnxW0yNCkdVilB6dPoEL+/LBIHezSfEHbrdOE7jUNsMfa2UGRxUD8J+KYu
yy4E4uZEuJ5+Wy4S8uJk5iKHDn4vKURlxV01OlIo/kj4se3mqiIGVx6eugnbPXY7
LYRvMrqW/qmuQutwDeFMwufEKpYkKXrH4Ir69cEGU2KhU2ej7Sw5DKhaRAIqtQrv
wqJpDgOH/NjN6XasB1NHxcUfQ2Wi+qfgxCcyVnzTa3Bm4lbNfMa1f//Lyyge1pdG
kdS2rKPFcuvbnfxwDjtoMSgrjLZp1lVM6xJVt3ZEyvjCXnD2W4LOFCRtyZDJpg3A
IGA0jp0xCMS89wTrZA+Nw1AE4/2JjIj0oe2EFlZeQF6j5a1VDv1QGEsKpkK9AhiJ
esmkMSbhw+BZH2nj5JcEbevMY/3LUCmiP2ogAK3h7aZXtRj4bdRdnSR6nmBJ4bdc
sC9SGBxGIVHsdBePATeDf8k8t7u+xllNWujbqDdoAYixvmpvf0DJqZwDG0AZW8jW
UA34GWnvfrHrX44UFwXoSYLrHEtoMb3/mPnosV9mG4BsNADWf3K0Puu+rTgS4DwR
WWU/pByUmHhnylFSLsxR+hFGdFAniHF5HVuaO3BbdGep75+jgDQn/j9keq/cp3N3
yzCWmyL2S3ghu8wOg28+8XU2FTQkhXmezkICcTZ7iPipOsr9V6OApzYvC+gsyRNK
pjZP5u+uFlOABE//wJmHiy52HnTpdAYypLZv44xtasAedJpBV2buqmP3MD+nygGR
swSG6FclfwP3hxtp7TlAPJBdNyLH5DfQy2fuhu9ymfX9zp50RDAvxgJoY0lbSNAh
mFWNjX1950d/tBWwAmkuO6bWR698fTQmTTXSbBWprXvuf1oWvax1Rz2m65N0TsqJ
e+FatNe3z61Gt5bPKq8wmZ70SMyXrJ2QikuQ1SR2vQIFt2Icqf/ia/orBWujcosg
fVWz8Ge256TI4xlRHcT4X6d7CP5p6SMIKqpd83PpbW7+qMFWDKvok72m0ESej/2q
gkZ/yy+S4M76Cm/2QdJMl8cb2lJ5LAUC/KTf+VPHsiiwrW6008NOHN+iUNc4BIo8
3HGHcE/YRG3CNTMRQ19tApTpsSOt/sa2azvwIuDef4qjmrdmGrCq3HKUWbT9Urg5
mw3IW/4i67LH9jRfdUBm1PQ+mNbZgZ8/ovbVNAbZI9dVW+TWNrQP7j3YHi2jKdN5
EKZSkzCyvtfHYkj6Jmtm/iGPmuQ+kcp/gMm2mH3l6qC9InZz/PreUQeYtQenomqr
aeGgIrkcZCRU/vJP/4+OviDTor4ryNfAd/tKEv9z+fqQt71TAwMTwS2dbc1lCuc7
rOtTCJ0OwcWAWRdn9KrubMvxSsjSAfP11jwzGydPyTWOfzZqBNipBBXD9njLrbAt
e6GRNu4sKMA95kIVgY205NkYx3XxWwbMOyzhQcl0b3O3seV8ms5IEkHS8t/MrsE1
pGIy8WZeMZzzM373e6Y+S2NvsrGtZ1L5z/EqvFGBJylje8zK4WObNBS5libfJB/z
X5IvkwivLV0y0nLX99epJ+2OqDgU6UihpmXqHpHPlfB7OJf6syC9juUIi4REs+70
tc5WaYzdXmPuGLKRi6fuZT9I0cvxB1UMpU2VVjevJntWYFg2CJJDKn42q1zWDpG3
8kSoLT2bwTdO9/k/IKW6QaksuXsdSZUp0ig7rF9/AtMqZXSSP37zd1Yft65rMCqT
z7ZyTUIwLUVX6AVy3Pom39/XF5u5cQhxIM1qnIGC4KCpiaN9fZP4/LNOiZFU5bLY
PtA90vS93CVxPHeuWyavZjX8qM1ffv3UyDizWRzTlNU74NG9T085J6h8GGLHRz5a
b7JI2SUhO2hrIQedhhfJ1Qu5q7SVj+KrsoAMO8vj7UCT4yVv/3l8gjqMPFX5zcPL
WHQMAlTUYwWRbtJdufWX9t2Ppvzh/cwfQydOGcSd/bDQNJPKbzRL859migK/6UF0
/c/pfDTesniwCDk6TLh5PYR3GR9oqMs5lGbh8IqenaX5RYlGsnu1R+El2FXw/3dK
21CXV5OumCQ2fvN/TJyOxWhpHWJzj14KtR2Eg0nTKZuY2ELxID0oH6xxos6Xudzq
MPuTxcAJsHeGHMMGhpYwCSaM7aZTeugvh7DUbbTMO/8WM0foXC+pHOuCTQ6VU7eA
7r8MB0hJtOHtT7l8PdefWYQOTrH/ZBN2AeNmFd2nFf6gAaUdmZqnwyCaZK4NO+BE
iL42VcIcgQsebvfdtyra24CNZLHhcYCgcrpRa5QMh/UPr4Pbl0BvFxM8U9d9MqLR
jm2jh8qVzDnrL0TfPS2PBZ6P/60sr5ZaTZnvvC6pe6+zgOVlQ4a3cnC0Wt4URchA
fjnnE2soauIIYOZtog2076rY9+hJ4CiJQFl/VmJIsGjU/dSniisfrNmfaxtjVxTj
tpF0a/I3RJZmv5Xj01ixQfyrufucnOOG9mHaQ07f8QgX5gdJaAkcVR/1xnEDIB4w
Gi1HMpuV5lS35t12SCrWTxNN+HfznWwNBl3KqCL+SA55kJ1x/T0/MW8QrPTePz6p
JIfrhW7t8NVQlMvWP56BurvWNWBEkmGDa3CDv6hNsE1+DIUyNgtkmzUc85ARhzQq
59xrHMayTXycvRMreEW1P9/7mrTtlWxjMAZOD4q93GuHoDWK2yi3tLgTHu1i4miN
FKtnu6dd+EbCKQzj6gPHtLVsaUSnD47LF04ZX+jlkyRKGo4qb9C4Yepeglwz6wXU
7OLViz9n1sGIafOp/Hcf+2+J56BOa2KJXIIWRCFg7m8JO5nIVXYrpvKN0zrQB+WL
hXM3ITLiDVRQTaHbQ8lMSj0voLImoiont20EfDba8qH8Okl5SuveFL4wYOQxJfQN
NeXdUP3KZwMnHL6EgduqJzPV+4BzuMnLZPLCaKAMA08gXN8YKomvnSQv2JEy8alr
IciRrcbZztyUlO8C3oU60nrVbNyXYZqzNm5x0RjUsUBXHgB+0+xAeuOPVyt5ljY9
mFQEHSj8TBvIZwuL3Osw3uTS99dsXzWVH3yZV0SXRUr/Vluw8dtuKKtFsEwrYgsu
CMLnNHekXgPLf8FpiOkGdd9lv7cmb8IwhtBHokFBkuijfwWJQQyA+XHw3/c5nCW/
0B49PJw7sdqZG260pL5lRPfkn5wz5uoGicS4Rw0Mq+ThlRBCQ8nx81sRnQ0Cb6xb
xshodz/idAFtjhsxhizykB/bzMrB8YLnl4/eBk4qL4ECRDDU3F54Zvsmk9fZs+La
mS9dOpjXtQFuqtPfglRz6EE7+h6K0eFxw74TsFhOr1JF4hHcD3gNEDoTeIt2kkEo
6s9rPzeTaB3gNCeVOhajYuRHi/XvQdjLjb/SbcEyQAdXlRfkf4piJK7FS0ASLKNf
WRH0oQv0kwMAkBUiJeUAkBdag+h9uQW0/zmy38eNSYb9I37uTX/Dz/CRB9LAlMrE
a3W9TVb8AdYHpU9nUnTFyajFUok9VHeVMh0uuLciyRmXU5JG0YdMytRVGlANIT76
LuNulqrk7VHoVNnTWH/hbxgJ77Ftyly1DKPvpsmdoWiGy94ddoGLoFLR1/QnF65w
NPJX62df6XHJeUaAUO4XVbN5OypPZ5XBKe8IAqtHpxH1B7jmZCw41zasqPqd2KrY
B0ulD0ZfnFAT6b/TqeYD5NVWpkOL5In72HR5HY23F7jEOOirtGkiMQqVhibLv9QI
/AsXsrytVKjLsPjw6OWafd6Ki13sxo2v1B+v+SuL/rUyq1oapETjRrgAP210OA1G
gFM+z9ELVo/Oh5burzvwnGS2dZ493+2OZt10TRnOl9Uao61jKemLLdUE6U+5LhSg
2zB1hxT+qDOyCmBJkC/kNuBXK9/IOSob18Y2S6vWxz/xHH/WCcS1cn80vJISVSKx
K1zw80zl9xF7XEz2KeeyvUaEx/oxmL0/lxb8tHxZBu+6UnXSBIV5Btk/skGIygOz
hUhOjnK03/V31x8wVCOKamyWZfY4G5+GlvlO9fWfOB3+z2kN0WAxgePdW1UYwJgq
l8BCabX1tCFlDoZ2t3bN+Ms7OezdxFvuwPtR9KyH8hM4j9uliC2N37zbG3+n7LlB
O4glbAHcj/3D019FdiBNNEWUuSjKmi22X5f3xy31umqWtcIr0xQqxZJ0Z0bmaJq7
KF2xTOjUivT0sEQz0GeJwQricKhstta7HgZuPYdt+nQaxaCIsfEKdCM6b5ViPJ78
xtjr/2MPQ57zKbm4qCT8MbZOtlk8lOuz0WeDOKf2n5SaXvD+4WG8a6twkJygKb5F
cgLoKQG5Yk8AnSEqk1y0Of2Bb3Jkv8iGLBDa9Fj5FIn6sOSKMnkPBRE8FGXFZHnY
9fO80IKtFxyGVLBKHG25wY6TZYXQdktm9ViDTHndRtPn7IBwRr1LIDSmueyNFiEu
k5WihqiEuSGV1771ww7hFX3tPqxQFOxOxjey2JEIhUU94Cp6Gp+RrMzwOMfD7Sk0
xUSer4Jq0TUYjUv/vpfd8duhf0Whhtx75pvq1IJunkR6vQ2USEGwKd95nGy2aJBZ
vvDetYE8UVWk/aRyVB3ObI92nRfTyYetz/V68NlYriQwo5ngtc4VF8ch7Q8tOZxI
uZNAp/aDNNibj8bLw2e2faOCaW3WVKmuRV6apYRmvcDS9V+D4VIvrwHtJs7dgRoZ
kiE3JZRlZmhFDHOqlrkoW/2+Vf69uexrCao6ZF+SDbtUUWJkoxuU0hj4irYwndpa
dWGdYuZyUxMmx3OWGc5YnHA14Xa9Mvih3mtU6ZUZV02y0m0NgtO735wyBZy9X5rx
ocbbFogeVzX5g1vn3ryEy9OYwjdlG8GiQsE2i/1duqmlcAWZMqEL3QbrqbxwRYw/
/JiKVOS5FLcARSj4eLHes6/8xwmJ+oBopuCySq8pCTNSeUqeWeoDWTtYqfYcryz6
2dLN3+oU4wHjhbujhVOeKkmEvjTpdJP/XJLna8hiFOGFkcXYXOYax5XWVOEmd5iZ
LVLsEYni0lxHiYxFFB1a5DgVPLdQsr8l506LVdlPByS71CK5o+Cr9tC3w43PzQUN
yYGeegxum8Lw8ONMjR4Bsm1k9tFfhjPYyhmViop+7bCEFfjtQEbbYH7w6sQQu447
mVogbZNqUmxu3bdtw/SPzskese6YGcPbmrdDxMq1XN+TL7cw0clUrWilsIuIEMWC
2T7f6Ov0pUW2/roJ1kwGpG/K0OsqNJcC3YIOCFxZKS7i9KneXeKfTk1i2ALHeFBt
JowFOi6NmJrzk3Dk2u2rnAIoZMdMoKPVr1swZUZbqU+HuOjPQA7mxu6vsqcCH+bg
dLVYEALtefmN5fJyOVyiQk4sGHFH696m71zzijusURC6TlwZd2d+Gs1VLlq/yGAs
GfYB9jgAhyeO7DPZkOURfKTcvqfyhp99awXNa05qh5YOZybakxRnLfva6gi5vRuC
RJP1skoaq+5LjwkowoHS//UJjOZ4xDqWb5pyWVkh70hS6PCfxvqKeKRhVwAMVfyh
MwFeDDQm3n2p1weGrsznRmoLVYUwLD0BJqRgtIPQsthNehuNRPBb/B87KUjsyLFA
QC4clhM85+S6XcIAdHPtNUnc3TphFu9EbRr8M7Brz0CvZK4mgkcz+Wddg8X80kFZ
mEJTzWXkQZvKo4yPVbBrhnsmoAKxJ505UL52WW97lWd5t5IAi7CXlI9sJnbEMvEB
sw0VCGb9rTNUUVclmgVKxf7J6DooztmYGfY6WiUat6MdNUg6cuI1iRrYsjSZXUgY
voOk6Nb2Quye4rmnTnnFcGJD+B3xAkqYrivn6HUgMu1c/Pt4T2usuTH72/ywEjl9
T+Gh/xoSvYoHDIXV0Rn+Po9Annw+R9bLEJV7SCdQ6xz+8AwAZyhdoJWoxlkR2mWF
1jyeLFKudcmY1Dou3/cc+ET2Bq0FXRySBSW6COzf1lDQN++X76eEOJODb+xXXGBm
kW5nXkcumz2Ym8eNMBEz5TRZbaoRGUQ5hvabK2gmu2gRkkELq/u68l3nMUx0+yVX
qLI43uE29fuVlsIu21L6dDZwWXksSUGKwV1vuAfZGg55LGyeDLKTq+SojS6e3pS9
y3P4hqpQiueItc9dK+GB/JOx3qtbP/TnlK7BWoR45uNALzSPHt+17nMLsx8eBlQE
mGpBKDjfFSTQTwZvJvnt5Va2AShzbhri1iiCe/IASqDW6VGWFbUqiXvuLDn5L0i4
5kLXTkgiRsv9K5fshEFG05V4GTERnZ3nkV3l7x07602KG5pMZ/n/2dHJHxXTPfTW
t90cv2ATbuNuFtIrJmyYc+bPTHN0g1Jc+LZLpvslJ1AMUflRo2z2XZuhpzL/KxCA
jwxskBbLLbU0KsvPfGtiVJZzc1s6rVPQA2/pKlAf/MiXIu/hPDqEjb6Y/WDyj4f4
XELCYLq1PgZo0wsCjfCI+RQ33S1hwFtXWPWXwpQJGFCmlkmg40ykTEgUCt43c0Ln
HsRNvlRR2w5FGahUa9eRFiqkEwuonW1UIkpn49xj7BESqZdoRb91GqCmk/CVSXHp
bfAv5rfGgpq2ux/yn4d1Zz9g58vJ6y/xenAl+nZoyKjeS4OT8RbE44W2YHjSdRKE
WK/E79rAOfzNxE0to6SZYNKggjzy+2vxJyRi5rV5jieLQCKhbdoCMplqzHtBqmo9
dNeMm5wl4PaI96rngGTZe/NF2yokoZhF4dfpvp97IduBlirExy0sbNOLdjCTuSVx
yNgacNqQm8lQmd080v+Yr5Ian+08tz+4JGL5Nbl41eClWSMurnQRd+6+5qLMl30z
eJDT8r48OyM8PI1rMmQJWNvqKWzKvxuWBJZj74Yz4OdX5erHtR6rgITuOzoEviOA
gSti4e6S/yhiESElgtaREd/tEvprsP7oKhEXcbfqzpKF0/n7qIPSCulz3DqQqJeI
eWxgDA43n4slZ8lK2qKweK7l/vc4R+SxUsi657PAG/je3mMW7IAPsuGnaSWtuBsJ
2o340rr3ONgUr3TxyGVcath+aoSTjhMOtpo77HWwMs/8rZvk14xim8W1kQWxQJKO
5I3mNwEvukB1LAjfNGHQAL4jyuAZZTZFcUjWyyWdOr0W+DPb4yEltqPzsUX5bmg3
1oe7msQbd1+w2SkPaIf0nFK9ZQRe62Zs8TpKs0klu9yyr4PcEgtKyXVGTCYkImeV
5QrywDIoFRfNj7LRbmMjEL9LlMnYfSBGHI2UY388hiSmtNGHTru0ioizwERvS7DC
1B0Gc33GyMZJsIaJWiK2G5FBTo6PxreavBglIqLk/EoAX9nbe7i6FFN+IRKI8GG8
f1CwHxzb1szO4nFrunlWy3i74dQNecPZXRSqGgU4NJ4U2o5QSKwD+t+qK16oSSEs
P1zUJwXFl17pY8YhOj5E3SyMtT5FZrtrNfwaRkxqICyzGkjTJRlxjHxqEEvQTQ+w
1T4xOS3URGbyj0a7SBDse9no2E9FZu5IZDSrnJFD/3jC2xkXm8VimeeYyjivL5kH
hzyPmZLVbyxs4dRt9eQNAWiRy6dy7TlBrK3cCuwicai6KJyZiuV3bMm2nNkp5BEV
U7XBDWLILlW4r/5MAGfgDbx2GcnfZ5IrJx0e4A+KPaYLezdt9F5yQoou6pFq9LiX
ULFqRxBg+5yDL3jw5XGE9uspPU49kBeCxkMmZPfT3hz5KIFhhcDeWFQ3feGkIJVD
1FqVCA9uUWadWBuljgwfFjFiPLCSsQbRAIyr7KqQcklv3nkLRkSunwwcZGvnf54R
rV1WXm+Fy7uyVCmsJnbbZmChKafDRBolOJlF4y6OxgOztlR82gHuSuF2hkbohD8Y
OhFSt7ZkGMvYtjl83uKAfsXzCRD+UNmVN/wQaPHVokkzhVYkSmvg9czY/tHyVZli
52OMXj6OKozZ2ALdiuU7K48MSchOSaBjCRBEKaFLowKVhWsGeTNv1F/F7YWgeKYC
VLP70Mjm1MQB3toaNn1vJ2buU4hkEw+W9wPVUYfbh/TLm8AwxOwhvYqqucH5kYpH
ifuSE+2fI6dCDibeuopq1t+zDX5KDh7p3YxB0dGW9IqfqJWy+0o36Q4C/Oo5SulV
Z/9wYMCJ8zYQSHTes4NUE1AyfBC5z8+S7ZOc6UgVEfi1ZKHgsG5nHJPEJ2q3ecI9
lAcLNc2EwdX4+ENdRNYLzCDRW5KO3LKzvfuMOQRaDnk8NYyJ2nDY5RSaqdQrgra2
tPFkdXNJlBhpRhJN1Z41hePWeSAkFxTCGx+/XTBLnhV13VO2nApNj4iF6hHmowp5
d/HllepC8Kyoo+KT2DEixSzPksGMVmlhp2nDOnKL8wYiD0tsXOUGGTDb1JQM4msY
MhdUdu7ElqVeYmgsDZLRZC9J/Zeq2wV6phSE77UikZ8Z96vfaiP5xBZJVaE5MHdu
zg6SXBJc/ZkRxc/zR/OZMpOIIjth6EYYD5NXVUBlD7FLzOUPqxebhzdkFRAtwLyc
CrPzYiam3tO7f2knyrQbrevmMzk2cDEz1ZPlrM9FE6CFvS2MtEfSByEVNROF2RPr
REqksogHKHr0FLJ8cyWl2TtMR179ge3VYF3RrA1ZrjrnVYYKN3fm+LJwb4JufpIs
bjyg2Cx1Fd1BeqJpTnr+umepufwvsejHd0yOcMnJ0YRxHx53RATHp/3IlSjJXeqd
//GuWSVmqeB56uDMvJuOPLphTYMvXM3CfIGN8UDre/batys7QFMXS+c7XT4Fo/pD
CFptfFIvei87bBhjNi1zAgclTPL7Q+5zraKMsbPxYtU2p32Id6Xq8hcq+sAOtVXX
YIvdwLtRwIc0zYqJatnh7/T/hczRdrnHqEzw8jG7aEtfMA+bInOQBDyZOL+L9nY2
P5STEh2wNhPSotx1FTPyVfKAQqUCb1VvFqwgmd984YQKwyERp1VviC3aDFMNCUyB
FKbLxm9HjXcuAMMd81dDYjwkKL7v1OGMzRNk/37cvfU5nCvpWXps1YQbhX3YeK4M
TizToUB8OZk2Wwn/pozOCeVJlRphXFpU9A0kTqqus+NEQGcKkB/yiCmI0oziedY7
kxc0ZlhtGP/ybC8oCFU7d0IiLpElhOxfNJYJSLwGv3aRBbNC8EQEZd8oMwM3kLOR
bktmCmcNnFxJjJ8tw5FTu6uZ8TZt109GjXf8wqC/cWqH9RSfzs+jjsRkz8Zh2sLt
jd7p0DxkmnuV7yxddwjBz6L7oht776ZABWNf5rQBbjnKIqVTZPqerEtOAuKg+66a
jf84vilKSxxXQJ6GfMD0VY+9QSM04c3Y1buCXNHw3D2GetMl0trEdaYlh6J/WpN4
CGb6PzxYNtZjP5jpRHgSXv+VnTYhMEFBeUofD1fct3Yk9uscgFZixDb0VDkPvRWn
8eMQTcozZf7v5HtOBuy9L+iYNDn9J7FWayBlaUxYuRvb8eU9nvf5bICK7cm9fK97
AeQe0IxnxEyUIeT6raC4nzWTbGx8r00IEdIwJ1l+xg9Myhy/vJLGkU+gkIYQkYI3
fWOq6gdfOlLRV/icnz+acw4cLCHXKrJsuVAiJcSAuO3Bnlo9Njc1m0gA3w49Gh7M
GJQBw+hwOP5nXE0puZjfCvTFaiXWmflH9/v/sK7De2lGsyQa10W6pq6/d+1wot5A
zcAhwwXQKzKf+KpCxsEi+AUP1D/8actzuupGTl3a1UpNbnxVYvviYJax3p9bqh6c
ZjrSonw3xtKF/s89XxUZXYsAMlRZA8d9DoPfLQMGKDd3UHM6EaRIadc/D/GsVACD
gfq4zAYiWSv3D0dc8D/dDO+ERbdrw/u0xY9DnqIhi8S+aDwjCtdn6f9sWnaMF7pc
4W+8+MhrT+ZoQbAXNrpBjG+4zHT/gh2q8STUzi/V05ZOxM95XGuuZvbX+UFveGln
pQZtqMU4OzGYApLFwI1XPHzp8bmQ4U29trbO04JFOVK2ysd81lI7bvh0kqbNH+/T
7/SHLiTwqPXE6SvUi6w6m+LPAdUdIA18s/G+7x4o+9EiYR6S4Ue4m16m3cfMe0Yr
FL120EoS7+b5hIGfr3W5UJT0L1uotE2g5rCE3mxpHYbGdDdFNhZZ+Bl2dHI25CZk
Bu2l9xylfkk4i84ODUI6kimaxgphjAzyJJniB3SxToVzZoFXkMvYLhKUeF846gGj
NGtNsBKIbXx228XsuRdknn6AhNppqeMMl4q6jmV7SOI8hvdy3chgsI2J6exSvVEw
k9qBAeGV+hTWoCcQS8a484RyFwEvK64003wSsnfo42jTRcAi7i46GrqF78IcUGen
1AVLBv1XOZGnvpi753hV7bpaDlFXIpK4lSrv4TA1fQLMhbED5vsWKo+BR+52roaK
g1tcRsAgf4vjFaCbU+39I1+jNPWlN3whbkJKRXb1kTC8mFARAnqf7sgycoisptm1
Jidk6qx5hDBSPut/4GvDFOYXqS40Hyf7p69BONKu9lH/N3xmPsegRh5ppMJgKQOC
tLxCC1f/jKWiv+8pE3Eeg3rvbjML/rjCXFlqG1qJsbOOWbRss6tda9nTxEP9g3Vr
WRx8oCQd8V1rGXCNu7STHm13llQLrnQUkD4EDH0OkDQ4aq3yJoyM2hARoZubJNhe
tBxGKdXjQKRd6RKbTQz/rOM607Xf83kIN7Y57xMOgcSqU/YFUbdVcKEPhUuEz6wy
8iRpL5rj2wi4pU1Bb76e+5e3aAMQddit+78MMnchsjeO9nkYf/3SIvVrM76hddR9
sPVoMwKi8p+mkOHumBGCDJ5J3UM4dgVnz9m/pKLs8+MOm9ZW3jQ3+XCpRE5EJ9nN
hH63JexbSoREIu0RSor48PbILu/Xaxoqe8U28QGeyj1BqXSQNAok5583DBb+duCb
85OZGyID5hg4ctbJPf3lyhEQiakVL0cWUILOmG3DTO053viZXv0uJWtgy4M89mST
czR1RQW3tC7uSeY9BXhPGMHEORenoioOgwi4kv24vWNZGyS7hf/wytozyVK0watw
dzVme683rHnag36auEd6fJPR95mZumoPpBO0GzbynOSBmS4pAYPBCUekkuBBlDT5
ExfvwjAHIYdtI5RjWtB3giIRiBKyMd+5Wq55C5F8TUq/qeyJF/q8nlf4cUAmD6uO
ZVegg0xL5bnS1g3Vgh2zumOPnjE9CS5z64aqXqPwwkWlXRn5crPZUTW0HiHnkUjq
JN/hruXEsoo+yRiHjJFVMs4LwlgtVLkXQARkMj9mvcfAfZf3/653gTyPF8uYgFrL
XlHe2s0g5/94YyHwwyF7JQ6CFmm0f9DW/ms3lVGQzMtbPLvfUIqlS+2+jlTYA6ko
TgVKlpD1HXgFsnWEeIWdpQXxkt8sqpybBJxsH5nS19Nyv+qNfM0binZPuTJHoJpq
cELYBPGHDkmzhI8Pr2OD9+6t+7puw8MseDpmx5AQaR60CW3FnYvtHolk1/Vkx53S
xWdDBfjMnyGP6wam2X43wns0RiX6v+FpmIonUgz7Dp5ImI9xM9foDtMIG+ppH93t
tLw5YtO8deoPDED+O767JzwhDdEqxzoZHk6ZDAzjwHitCSmlyda8h90AChygOnrs
H/NX4h8MCudNsCecMal6Z2KgY9hnvoHhRRT8kf9PzgN6017Za6GpYcid2zxMWscU
aWa0Eyo1oNYUYLt4KLfQIjzSWLGp57669LSQGd1pfcv+L/QccJTRno24cOo9BMWL
XG0Trn5qQfNQ6gWm7CpNqwnJ+TLJgAEeCDtNbPwTELlLMfY7T9XyquNhKkmplE1u
gaDv9f8n20O8ph+FZB3+QCZlBM/gTIOWSgKk0DQoHGeOq/VNhwpT5o6hqerYMA1s
KVxkmov8IW1bqMFnqG0EaUG053W3iK8JA7E808LjrhL6rYwZGsJthplrY/1hYBV+
9cqGJmTceRC7HChRbbMRL+df7XhCK7Gn+oQbD5/jO8ylR5CYnzAB/jWOonaeGfDX
V+tH32BR10i8/du1G/25UBwVXViFo7yBlKxaAJvejJfzep1IeRMPUMqsXPKwe+NT
R6JEGzqqEyJxGwXLqNTKs4wTw54er7jkBu5+St3YYbyxGRGOeDh7LljF479phiqV
c0wnI9qKDDmR6jNV41mJRH/VUxB4r6+p8hvDqMU9rjgiIPh64bttMUaIH60c2r9g
GFbp3qS+E6rxIj8Sg3Dnf8cFo8p4uwNAmxt4+sqaelA5P9fNYnGJx/jYQZyB/CR1
/nhpA9GSNe8N7IkdxPHGIfdv28TXRLw2/vvnItAyTu3QSI1ePgFkSP4DZbssElbv
SYfuj5d502kcTMsunFjp0uBkTwB6i2C35syc+RzSybDjr+BDo64IeyBFzaYwPcoV
5FH8NUualNDcRrH+5Yu9hbxh/B+4Tp9F6WogMOKZFVnT+4j0tRmahxAot3gp4yAH
Sw5kmZ1+GjvzHWOQzQn8EHLCqSJrEFOCX8OjmvicdKtBqcJFaQPnw3yeSuBymBDm
VvJ9hNvoQvz3g0+2BpJbluL245mzZRTi4XnY11EmbN3bywg/mGJ5JOEsg3o+y7ZT
lK2n8v/1l3dz6zKtJa5RTBewmhXnL5XxPU4FKIRzNO0ODTSq6cbMVvvOPlq6RN9h
f5KF2m7nVKyDPEcRpzsKV+Za1YOLM8hbbrxG4BTtXp0fzojWO6h0yEMMmijIoaPZ
qKZpzbwbdSiEPo6D2DGPwaczOWTY5tQtreW7i8LECHNMlxxJuUHNJeGgCTZPYjyF
CuHg+ZLXWoVIW4iTzWWXkHl0HgZhfCArFgeGRvxkgNA0QZj58QQVIvhvBCMsKFWk
UDmCx1RvGH0gHqTcZ09hMPBb+p3/AjNNc2tWst+JCqWWRpHIXDEsD2gJdYpgvAP8
TwbeUeBIlZb/bdeCLfYo3gjLuVrjYf+bUUWE2/F+jt6ZdwdIWFrbvJfpgWm8osjo
kwVvMRoz8da89J806j/cVDJ05Rn0vWbQp/vYu4d4NXlwBQ8xNkYKx7kSSVMJnvbO
uWzGw6R7LRZE7/AdCGrO2AQhtbbZyUWucqM6hDcdJjlDgOL/9vE6G/VM8oKbkPl9
zUVqU16A0LD06h0rJQY3+63GCLcrmSb6/HL1B21daAG5hchvQis4VM6hgCuTSE15
Fz87a3B1iJzRXz7PSOlXcr8ZgGWILJtaSkUEzxovVRe0ttvsgI08cLKJHZMM3kIs
YY6NZJDMv1rv3PiR5tW7eG5rATN5Teys6ZsGXS+AbMWNCqVvXM/It3iAQttoF0Br
j1/m5q5iwcvp2RtzLQTzt9G42JjZ9ZRDK5/he+fAWOtJs5MnDPU+ZA2DNNxL1oUS
M7knot+iH1TLrPoEA/KCVGVchTQNeEtY+XRLHO/jzbUIpt2yg6QRD8FjggwyXf5w
a8WnAkMp0IatLQFic9JT/ZRxrE9oGt/CeQ3M7LVgSMgX1lB27KpjIuRfdY5Yonn3
asegFeV6b2howXdiETBkoHGhOAB9XsLDRW2bsBQCdmuktGUJAWJfqghQA0+QbLhK
L8cfhKDKgYpwwcP/B7I4BYVpfcrQ3akLjLZNJC98U46mLw41EmoO3Tz6BflPhSUv
w1phmZmg/jMnNagFAqVk0T4f75al39niKUgua6ffo9CgH1Ab7Mm9CWUCxgXw0OuH
juHLaSin5AdphGEoEeqnP/QsomNot6bKBN5H3Zb0u42LeOjeWbF8Xe+MiiayA3zv
Y5yD04Amg7ZE9JHYawfGi4TKqv7EPAo+Gxo4ax5Be3tC1oEDpBZa5rxM+Tgv+aQ2
g4EW6i4TDo7LufQ53UDK+k7z3P0wSbYyLucil4uBA0vzsyygjUPQRANfe30aeq0H
rrtdvsyUh8NaGoRimGkTO1A11SiTwDGzpVxgRkjsa38XOJTUImTmITtHlLhV9G4m
ZPfuG3Qj5OqYLbEFui0jfRIpbskO7QxMSB4KoASZOMt29sfuhT1CX6hVTo+L1Wk5
17DQYKg1Z+58z30ysSHzFaV+56jl51iTHX8E5aOmYP3K2SYppSfHwZhWFhFP04dM
KFd57YQJ0aRpB0tf+KBVqsG/bis9YL2mRb/VQrnwFvEPS8xQwuUg5BqBDAJxBYel
vHCQA7ZPyO4NAwnM8FaVm4EgwpQnIgTXOGyZOlxzWmU5xa699gn4BTTqS13116Xz
KvuFNkhTOEev8m0YwjtfTjPMTjIbwm7f4+PNIPbzRQht/FUVy/CgG/sJcOKXsT+H
ScodKVqKuhVZZdHVY7HGfb8YkCyv9LMt6cjMS/qr0d44WtR1ZTb0ptBzz0JSKDnv
Wh20FAuqWMvcOYW7sjsKkpGlXhfDahRgQdl4eoB7XO52YLXVOqK7xMmKizkWmhKj
+139lInnlbhXda2vQNRs6YlzQuoGmXeT+3i7LVQ4PJQcEQyv4BF7hY44b/1GZKeY
fjxHlrZyuo69DtuxloDBDnMnXA2m7jp9MvIUfqHgUey8TPQLxfwzAcamvtAAC/UJ
akqQE8rNvdE1WOxpVHy/9Az8xu2Tbzrb++T+tk0ryM7W5BC59vx3TRXW5sNymfkT
BbP/NC3NPhdMiimcB2O77oVtK38Xg5SVw0K7koSTowO9qi2aReDfugU+mW6ZjFrL
P5RU6OrvpwCw0QrL52JXmQKgUfh391KhfQn4Jpb+L0jFk9k6qW7kQ3oLXIaXX4B7
2ttJ8I1FFywsnXr74WH5belk72qc6rmN8EW9ADd0NY+ULqcVGQzXechgNzqDGQll
Ztk0MVXuYh6c9oaC5VOUfhPyYNWw07cp5TJsr0jJSJ1rXVUTCLunLNuYelCk8wmv
O4I+3MbUliyTDBl6bBvgasiAtKK43iPOH7zHSqc1+NFveaPrZp8n7Aq6QmSQm32k
W2kWA4ZbRouUjfNM0ullmczfmYAPk8lB/Yr0TwJ20J24hNShpegcvQZi0FB6P7mP
85a+ZBGS8CMoG3KCwPlPx1kGek9qlE6Gg1cd9/PTT0Tj5NdlOer9X/lGKdpYi06y
h+CGTOVexP8kFZ5iuaiXfWystWWneSg/Z172RAB4APG5H7dftWhFrSeB6ni6jOZT
zTNafPJ+v8vx+bz1FpvL2b9mvnpjL99cNyr43u+TdbL/6v7jCgYstGFiK8TcgVdF
x4Xehttbejk1Hb8tWZ7gbPNycR8bmWEHLkxNB3LNRvzvwP2uNZYP+GUcP3kp09k5
5YoNfyP6MfzRkBQPJCNkc25zq4Gxrck0xhz4H+WQpXN+F48BCPqi8kJDTJ9XhgBx
C3CqS8J8sKdp2JKvt5BLNBMSZ1QQoY50og34gCersftLfSRikJqgChDAD8tNlfOQ
h77EOXXhFoRMzNsBO1ZQsL69280OpxJpJ4my1nRtvbPJVzZQkVkhiyA7yE5RD8xW
4Pl/Gzx8Ss6UUKNPZJ1cbw7sS/99C5uHVMw8ILi4rhdHEugiyxfH6BKdqR3mCkJ8
xglsSYyCOc69sctzn88tmGuZ/4VfaIxZeCcj7IGupuOc1G3gdpQgpO6TnZFJLUhZ
GuizHsRISJaPiTPC9ffqSMak4yJdOXhjgZ/qTTPT84fce2S/SKyu4lulLnDPW9lZ
d0q9o817BhQzIlAmrzaIUx5VtM0E8foFsS8Qkp0XXjM1jL/2VYhhrJw7DKHbWcg4
uaK+FYgbX6a5SvKqkcyHriPBU3wxYiHXsnVeEAg4O2kvyKtjX1nKr+2hTv3pFEg/
HritdaJ0gB3nNrzYD+ybOhFcJ0NtHpRjxIdpaNK+2+H6IFdThVmnFCcPiBJq+1hG
9J5FVZG3iFB0GtgEfB65twH9OT4gOkUSgFczdtXV0liMsBuEt7EcWO92KS5iExuK
44AvCkY/8kgjryW6VfF3VreX+vILI2NNLFp1VlzpMYWvAedO+Xnm6cTOVUHNrKRn
ryn2PhF5joU2j+PiLQifxj0TV1CZ9qIlGgPqon+Doi7PxyenNGH217L1+vZjjIPi
do/KPPjpfP7f6ta2Ccf0/R7S07Eks66Tw8kPZuzusbmbJ1eHUWkD83u8JVphjCS9
qcP2oXC+HIO6upq7axI5D9akXikhg1EUO/yk6tdg0hKdAspYQ5VJAEwl7lZxTW3i
X3L56tRLvthdC+Uranz/A+/hSdvB+Rx+psBHHJKotDbUCa6xf+hRr3qj9l1zzria
KpIMKzseVve5yPbpDltbBlNAz6BZLkBaaeDYYPom5iWieJ42IOVCwsCWpTMPMuVq
+PsE5lDQiGEY26pMZuvwTA232kqX4Kbt+WyjObzuRcjnHGgG/6rJTakFXcrEBawt
2Fiv6j6SqqhopBVUs7b85IkGOmnSfekr7mTje0E1uncHFgZZPpA+UJrlcQVYFSt0
xXJjHj4UqafcVh4qiK3M9W43JPq/LNzaXSc8GfyX2E3PcUHNwptVqeXYo9fx/8Se
Ip1YmIQvQWDnCvjHa7Ug8V5XeJ/dXLKkP9q1+djbJ8O1s4ku16e3RGLAy9boCRVZ
LFWcNJOp/g2SECPPIX8uc3WJf7Ee8mvS4KC2Ct6zYY2tLVviiXbuFHtg8B9DmcBM
kb1qZnT+/46ALHS2Uc8ezWrV3jY53lXJR/fMDNJt5psAx3kgLlfPTNqAAAgj0GmV
PVQSGNYN/V7x9eLNNwk1H68eioIMhAAXbj6RagZdhH8wANtq+FxlPFZ+Y4iOFxkg
LUqXn3uakeUUwtVCOnbiF9OnswogwveaS1o9lVn6zWx0m2avtUHg9kVBMB0N0Xby
U/aJcfn6YwfCv3iootkJ4sz4lk8bfe4bNR+xiL3hGMegvv8CfutHnTH2TUrMC3rh
59gGpSZ4AY9F3fdEJeM/lOAPp0dabnb/fMuDdfc/2UlhpeoY50rdcFExBZgYAac7
u1JQqt/zfmICvzWZUUHpI/i1rsQVyzsT4x/0EIApl9NgBeEWrH4TKeQTqqzv0OC7
CcJzm29f41mvHisdU/jdWKJgPEWTlLsnSBIy2aZyTqPui0sjExFGntig0hWPzOR6
+F6FZL48ZvB2i3SGv3nsWC19UpskdtYIJv9VvwsKLCBwk7V+0Lmo4N6dQnHgEr4o
xNKqjqjzEXWMnYREgWRNhi8JZiDcBgc5uctv8Mi+bDKzQEQa29WPTWbuibSrJuVj
YfP+EnqQfZIohd5/aqHc/Clx9/8R/l9qMp3GLchQ/HSD6XZ0tevr25PAVhTiggR0
JlMaNqyfaymlXQeyTbxCGNTipyPRDEEisi6XQP9aAGxy311oGn47xFOULF8/3ciG
3ZJd1l54HDraAHCaQiPqfLvrDB5aEwEXB+9ERy57Yw6kpDCPOBGoD8jTgccjsFo3
OnVwhznz9ZKw2+pRF2VJPZqduCooHctbKG32kABRcjgpsmhPT0uC7QcAvuQBKdcs
qZVkstVG/ooJdywmvlu4c8bVkdAvo4GFUL4BSck/AmjZ6PlBbpmMKRBrLxz2wAcg
jj0mfr0L8FG/I+d96/xgU7T6HZBJRAu/lC9GwaJ3akIWYtKgYyU9507lMFKi1/id
yrSqleyFrQwlQfDlVggqvbi/QLWdePa7pP/pfGJt5OwfMxNd1/c75qKGII0U6RX1
wal9uyTIb+FK1ugyjnRO+8/GCfH+PNY1EyeiPtsSH0pHAWV6mgFoCTcr/mAG/eq2
BaHJU7oZCvSzqDCfUN1DfcfpHEs4/08D/BVQf/zvxA83izOtaq/+cudU9OmEli01
VDauRPe7qHIBw9HAL5iSYCRvQTxEjI+j9OjfJ+6aypq9sSGK/2t2R5pYyVO1QWpd
Dic/MdgXokKTMQIpiR1ftz9HpGs+MMRhnfruLcHuKvpjNXmc+VUX+BlV1mXADJ5f
aJLwHHdOAUz5P1s9Muc2L/in9Fy8hfasLZmxCHOjRfrqaI4sxodlkHQnlBjdjOsl
4yEMeNMhJKwFaAfMAGdDNYoZwXsvlInHpmS+YpfjH/6K/JzPli9L5CiStfAm7LX7
+yBCoDh3Zee0v/Ittd8EywF9Utxt0jVEQUhkVryWebkKuw2WzblFTRv8iqz2SU+p
C2+NoNsqT5WIRU/5qx8bHyhUN/Xwf6Eh6YkZbEK5mgvYYz1x9+Izfw3yjOc/zlw8
8pg6wSR+ONfzG5oyI/k4s8G9q0n4q6J7HPXwaahH9jySHD7u2/xXAFlZV1+S3vnr
BcKAHVeNLlK5XR/b688x9zgug0DB8ibIIF3zxC5V235y1+J90QLrNO0obXNHI4NI
T2ypE5la+qFtCMVJzJDYhMiWDHnC2WgsqY0RmhjYeaNWMQpP/TJOqLyUDaDywIWM
AEm1o4CcTkWK+KRef3mKHtpEUgr3gx5y5NJG3i9DWK/WO3nYZD80ZBhIYhAxv4YZ
yUHU28f3jj1q/nstvEWJZomqbuAYdCxvbgT9ckb8WVEYHN1/ke8F1ijVWdsiRVDP
Hd0rQa36bZuJTrIwHyiGRXrKRuYXSDgwvmRh1K49poZQD72FkDPsagegbQvnesjM
QF8nYXVVQO1tvzmftGh61nVoPegqPdaCIb237mzFD6ef7Un3HKpTlXnYHl0Zxg3e
RB0PEcntGwt+eoxIB1047x4KN1P0OmbFKUHFEN3nB57kiTyANPvapbwhk7gTPtI2
XJuEFj2QDU1jNVOsf2U4HWbB0wYiilNyJK1QavK/CgfPrSe10XlhecF2jc9sqtMV
juCouDB48RcHUj+jGZax3SpOp0iebTZ8PMC+WI+vi55Asy+Kc/DS3eAQkWJUBOSw
Yw+YFR+vQctu+dIEwPpI0WFkgR5Q7wIXNnRX7UZPfUB/RHPrkYb/iDLp44vYEJgs
t+YIy+TxOZFJzS98KGxXpJz7/97xclMkWzbIs217bIGH/5I/t0ZIwaDJkWw4Ro6+
w7sp7TyJDcY0dpJLfh0AtvL7iPmAv2OkUkO6w/sn6fmfkHApTmCcHHovuybB93kB
BZiaX7ExWyjQGW5CECaFe1NNOvRVX/eI0LJDHuWXngMqSbhfOCdPp3dbqCLP+8vU
F6Rd4AjzP5c3t8zuavDj0ALJ9Hiqpu4FbvOaYZfw6FKrj0+wb2LmlCQlYMWQF2ib
3ouAorvh/NeH2h/J8T1efLWIOrzfpl/cBad7KHL5uh4Cs19iJ655uDRtFsCP4A+J
UqUNjiAuQ95GaCxp46gZEQknmKcCLg+aQoTg05p7EDhXtxDTpg0PAtKBPzgGk9BJ
Z03IDf3wCs8YpRFDZyO7BD1Olqvwg5wNXnj2HPWbERQGKfvnI2X4rlf0Lrdk7BFS
f6GAg0l7UdQHDKxd4f+KZlOHBI9GP25DBii1EsDTRlL0zqRfXFAiYDw6c50tpDDO
KDxX1TTqmF3sg+Zko+IhoPhB0mfUwBPs47IvKrrLYHxQCYmLVuWPID5EsL1XFMAP
Kzts/PPOfD0Nrl4+wxoBLYiIYMeT7ercl+sTgYL7PI+4Bwea12rOxAmoVtcmaKkr
zTNy7q8+6thE7Ibi1JGqlO5SrqWhPH/Qen2AcdJizp0vlE4YeRiLX/9FN8bcAKgW
ZslJ7ZyRc46ShnJ91vWvtU02mNxdYDyI2KSwFYFSYA1JkxiFSKdL37xYW+1cPCu5
/IZxWot822FRhyQ1uYA9grH+Ui8/JUmRIQbxznLEBI0NjjQ1Nm5+UJOFbbcoi3uv
mb+iH3CrwMdsfkRGH196kEINErK6f+/Nw+VmgdERVTST+hRUpOfxA2vT2dkSBqQ4
plcOOtNGbmPK5nJH9bzDMllNY6eSgxY13aY3A/LEKjy9Fc+ivGPYMbMLWU5oKfZh
xj/hA3k+URgihdpiprnXIhzsNAOH/Kl0yIbiNpCsjIy2iOW5w6qNV8E3YMJR2auj
jNFwFdQBoP7el6kbvGWYK8EBSi7XmWw3QYM+nShdINx6Lx47GcRbo8hQfWR4t9vq
kd6QR3y3GWtHo7J2VFR0bSTV5VvF1KKU9k57Hvl7lXqDP3EICbgAnJom4io0PHXu
XWH1gNOLvq+HLvq39UDGPmq8KWZ6M98O2WES3E/aqeZcHRoy5BXNBJxSOitfNNmE
t+9KyT5pCf8O5qtGKrZCc3VLSuetKLFeouZF6BuqPOyw1sJnq5CjQWLT28v12D4N
jv/fqvwgdHdElOu2bJXXhGg/EAORvMKDxDKWd5JEMtK+G7y6c6Mi/ZrXt18da6TD
i6a55pVfmLac1CrjZ+QxmG4dk1SfsIwiLxM++4F02U0DNmF6geI8TjE4IV/cmysF
1J7ZSRUebMFMcWUrRtq+woBnHH9rvPhkvDbiPeA3/KIdG+SQeldACDvZA66UV7rj
AKf+V1KdMcwkkxZeCRzv/8aXfac3p1IteJ+NcEl1ElUl8Ds7aYyAI6ti154llgFi
lXw9GoGXBlS+D0D9g+9/wJ83eedVxeuI4isV1q5IFVPJ2gYMJNTg9hadVP4SLqID
evLgS0V/IpA16KF+Uln8iac8GiN5fPV0mof7enav84AA1L0hYwCe0Vozz7mEq7Fv
BETJ0vdDNsSW5VY/vO7IB2PosbFiT3HW4xzoS5AXgtdhAmHotYNK6TqxOVoVPvAS
AmhJtW/yQvR/TC1xQiWtG6Tjcy53AlmGAMB62ZYPdML0wvVJXSaRcthTHwRKZm2j
aoB/xYremPOXRhF3dlfp2SBNYs/s8osxtNKUXchO69Bo7jcXMx62z94LT+4VWHmA
tMvaHeCTlUB0csISaTgnx/PDJ+YK2WHhg4aDIJzLarnkhb85RkCQgL/8KssFrSBe
uIl/FuUQbBYydLOaZFeBhcOYMn0peS2dSMmaX1fBggt1JZxPt9GHVpr10MVGnA8g
CBiQ0Yv7btqxKLUqijMzKKcxOtUnLW93GOnRb6quEwucaDup7mLcNRuqaqSAZ0OK
3xcJkTFyuYeBiP0B+M/jr0AnmMPdh6D3FMd+QQ5Ec0aGr+PK8gktsJYgoHz5eudH
Lwo8JtxZdpAB9V+HuQVNH9mGB3+k0anALFQtaZ3MGzlMzUljgwnbG9za660Mpuzu
90eOtsOoPfVkYNjItfk5OmlgD+uu0jAcup8SrMpzA0L+g7XfKNHTbVZwRiM0vwyv
YJ5/oGQ2BKRPTJ8m8m5wbjzhSN8mrxq5BkQeZ6IcE/YfYoz87eVgoiliVcHLEkkK
xxYTCg/9HHdctS5klaDsg+3oQXVG//xm9AMv7juKAW8tqk2qynAM2NKI8GbDdsB7
alQ68x5QzEqm1K0UShFn1MQI840fUHf69/YzuCI51wa9zzpOmxE/DlrMBzy2sAiJ
NLvAWqoq+F0vo8J4WWtYn3KYlO+LIqMEUKKB43F+U1dKMx49TFZ4mF/1ZyBxwLgw
JtAfqMAy8po3KPORrPud5OPwxYmmS7+MCGChzkTtfH4U33X1y/zL1mgyHA8tuX5X
n76m5hUZOYfucrqhcOX/P5g6KdWyitzR4zIH/uhTgb+izzVpxYtV0QGRDYPY1nRm
OU6UreXl909kjberKtS3rakAhIJ79E/Tg6xrqoLKlrs3A5NMGsWUXfuqAqgmmbK4
TfsQNp5QxL/BkKDGk2eEWYKVDR55AzwvQY2xILs8AwEHZDEE3SgwaN7JrDoXoy5n
sOrWJN6lQlrJ0vUt1hfSKbDz+OB6S7HUUe4h/WFyu42tnaahVKvPqXe2Whm0JMb6
/xHwMFGW3WqZRYaoVMJ4sgx0vROcRLD8EEqGWptFRcMVEGwOab7M4rNT1/ZTqBD9
OyVo4TAwETCPX482/ustGWFU2SxP/k1DUAedOIVBP/9Yb35Grwy1UN11fiKCJf6+
/HZ8vP5R+luEl8BprSJhawzFbIK48M5OM2P2QzvSJyXcY3RMITn2Az5Wwj113nuY
o3NjmIO9R32e0IDG4/lCkhOD3SZ265n+8JtNyEPekNIEoSr2khD2MeEjRIGdFvhu
ox7b+8XVKcd4eTbKvdAtm3GHklWLB4tvSntunku7uJ1fxh4DSnSiwnTzlYBFsUNn
r1m2sSTM/yj+IcyYsVVRMpd5b7eAE9a5wvis3wz8V73OFlIguWJLZuDD3eklsOAH
kPDxDxzHk0UQdcgvtbbnZMYaJk/hoSR0G3X5O2JH4OAYN6s9QZnaHbE3h0K8aHCK
C0yz9mhS3xX9/eKFlYFrT7UFeWB4TXFOCgb+WaCZr4UYPWVAGXNjc4zKoTndP3a6
xdCamw6IYNJYy/Hvs2pnnUMEOUdv2ZPv74DzrR0qOjMC8KBoEzmw2vwTnmLwFX3Q
ML+OXyvvL7FsKmaRf70b1cTaKhOF8w0HQAsWnQfIgzFGDE9gZPA+4YnZLJOeIuX7
SUQjoOHDkxLjEtERtM+RxtopftD33dY+njBtfku5+RmWoOD6cDofboBzc2BnLr0d
nVYk6xrnB5YrLmpWzN6rUfyIaAUibDZ7q9GVZRTHSEqkDsfWg1jjF8UU9FlF2AZz
UqJ5KeaJs8xg1u3ztNvxYRwfxv5N3Z1ElsQEZ6HkxcFoUJVdA+CiZeBZm2OoXRNG
AOgBqd8z0uKnlm6SrlLX0rXnnXNrnRAgw7LarMaUZCVQh0pMv2V1LiZT4Vuz33DW
lPALFSU01LeFSxmZZNA4OuPClBo2h++wyZzcykKfgB1qFmQ68/Qa0zohRMIsC6tK
EkRuaC5ivcXlv8YfBADXh1bLnwL2uh88PPxXlkUPOF1en+CWKzwAGCSVpfHtDGYS
c5wJ95a3GMf6ZlNqaevaN4hhH5zAYlL1uiyv1lFPHx4F96tBcS6dXnIAYLWAwkZY
Vrhllxmar1HJjtxFHtSzjoiiSCYb3NcWxRLlOpT+8wZaKs40rLasAC9BfpKWw2vk
Mv+X2LcvZYqsteR20CbCMUjcrps9Oat9X2pEVKaVnFIX+pB+T8Sl8XERwVJAUD09
MYIIE/Gv2glf6moUIx7cLV4z9/rWM6wOHndVnMLzjSho/C+Pwy7kDSYRr9mRYREp
QX/a4RJHfZ3O9gXgQ7AmsxV8+hdS1axw+dxVKMRgo65M/kmEQH3XiashLx6ejhne
DVjF8kVSFa40IcCGLbT8RRy66JhZENidZfMPhQILy7xv/uHzGPrN+5DRdlj8t39d
KvGOBNasmSsQkmQEnFHKGPqFuh1YJXWsS+mHq72KBZNPxB7F0pGFsXdOklTXmpN3
wzXWZ7cmbOe9YhnqUO1/PkUdrtjtN1k3OwbjnGPS46QF+8UOObh/3B3MrJW0QzEx
vPVYrr1anqzmaFFTu1Nk1YNTurYRMlhkEKqEZq3uOVSxU5ces1VSoSB6AUS43L6E
Id8qfYaFY1kzbHFvQ6vZqTiOB/6nD1TdBb08NsJPbJgwdwRbVhukcZXOQ42kFnJh
/Sl8/WAzwVqZ0o3FIvc154l2uZGizwBnWYFxWQyHJTCbc5AYPt6TXzJjwF8ad2yW
3FAvsekwP5+hVuWrbvXd8rh2r8xgnXOF2kPYx74lRNH/MOGOq1nhWBEXRWazrOu7
WtNEABHnp7B4C4vyfF/CHJNXbLc1ed5rvMmEKFfeGHUv/vsXCvUtEDLxkgxgNpAi
PprqGbotyw2rTyONkxXpMt0npwVWWBZrWUA9iTMt8Ge3bqtrInJXPdEMIeTCHbnz
VvoP/jLMfUxSVCS18nPg2nxA9frWXDT8fj9kWJVT3F3E+okoXZrwxTaL/YyeKs56
sC7607WsJkKYlUNMQ85d3MGBfa6unwDWzEkj9pl9eJrQY3KGViWYnXxvpIBOYRdi
5hJafxyndxdQOLlGL3Fi6Gh6/pP2VIePw8KpWLbmDYf5YiK9Yd41W4qDNFyGXFip
5Jfys3nBzM9DeXzaCe/LfMnxqOgXfceh06z4bobG84e897DOHAGceG25x69YZA9y
6EnBsJA/SnINk+0sNQI+VZlJIrHVHlQochARrS5wI3VgizaC1Z2zp86uVHuLszlM
RKwLStXquRBJ7k8KnUmrSmx7u75BL/Px77M2ZnCQBiqQU8nVggHZSZbcTMvHnjNw
uc+tMeaM/u26nA01fZVu+w7bUyDVgpKvhYjAK66M1fyVuGN8luR1O1lEpCSyL9ES
P8U8WdhBbpcxR2DVB3haWTrwGQXWL6AUsN/2WPzpzfH0drxU+D83Orc8iMJ01w4Z
/VqY1tvI9QTtjsoUCHLLaEzHG594GONu6OdLC1Nt2L3hqIcOGInR+05uI25TH3KA
67GQj+UEUlVST1xCYzdns8U7tNOnNgBdQ4UUqhjkd7ugJYdUB50sW8k8IWkyaLpg
gtLX4YRExTce/oCo8f3xld9GPL9fcgdZ3Zyji4kJ6Y5se93ug+w8JQJ6jwXewwEV
xaGBFMf0rZQg+QlfHMw2FRkzMckVJKR5yc+7eG5ZYFcgXrHlLNLX88Oqoy1RnIP9
nwEsN6LSbNtWPrO+kj1WEt76wJ0a8EakbFXzX2Zh9LD1TEh2lTHpZvHaflZ4MvDz
dDhQHgAKQQH91Y743fxfRhRhOEfoXBUm7L3XyJwCsTfWlT7H28QNavwDSxg1ETeg
Pk6vcKPK02vbkBhYLt/kKU2myQslyr80wdhwERmsNiyn8X3TLYZqcu8hhFZCwzdg
lOeeu4xlvM+cyCkaDKjEFrubcTFq7Ke7qL7ny3pdfTltJMLrelSJGZifEn8H0AqH
qXjiyHxxiNc4YkDSt/GIpCbWeeyUvkIWkd+vs9wDrGen5m6ojHvhkEDidS9v8sMM
KbpRLkc3OL010sf9vQK8B9VXBHUbNE0oQO3T9E/jIyHFBF7LRLx1Owp5YirVjsUa
CUhN+DrZ1en0mcXYnATLwF4rq9HEFBf/pkcJOhT+EWegAXuvxbeclGY/cGKi+Vef
gPuPUFZOu8AA3f5rSCuzFrzd4JgcRxvweh/62/AmQ0kLOymcmBJ35xo8ckatfhFB
1BnQGzBKnV/8ILN4glWkxijzq/vBf+GpeVmyQnCwTwXtAayqeFZb+WN5bdEenrE/
YCfP7n89xF5ieqvXK3HSpGvPZ548BxeK4+7h+oObDxXkJsM9bcODVAWgyoeKz3+4
qSvmY/sh2b0ZeqiC4ZFuqAkkcMBxr83RqVm27rpAdxNdOqQfsl/nAc03uiKVs77i
tQt5vI3mkn29attIhOdE0cxmd0tOgwe+yU59PCZZuGoueYgN6ubHnc5VSxKtENa4
UzA/nTI2succ9rH3sJt/RXMLrNU7xudv15GAjxfyrNSsosZ8DKkMTLcvSTwtLfss
VZn15EKz8A0FBhpn3bboVaNagokEZQVuX+0WD9yzQDrj8jPAF3+OdJPCt99Z3kKb
yD2TjQsZ0xrQv6pIXQIndLgCqiQP+rFxeyigBO0rEz1MN3mvXCVsGpdyf7K/c1Vf
h9qo2kATHuwG278CafOZlJVjY44l9yn84aywQ0jpxdnIHtI3C62ueGSqaYWXVgJ6
RXKmgCcBm5LNnXN1TmZTDvolFAhzqZa9n8n70bIwjU658zrwKsC+zIm2MqwBJ/R7
wAobUGvAkra9Sl7LvAqjtkXUZ9HZgqL7mY7Iw2rj037880VRZza/ufKzbXykhAGT
UPPN4DKyiLib3tQW6LL5D1sPThenBiLDnnALqfJZIr6TTSQalW75b/aYysepuzPA
yFYIcr/g6VGb/dkplpn9HvXZ7M5Mt8HoIEAThr9FWgH/+lQZ8PQXvFDolCLx5Z40
be/h20LiFgklTTuA2dGORINwqeCoD9Sxg7E9fdBlRhEjslMmFhkDZna87v94NF3d
bgbClQpie7Ui2TtBt69W/ClabnTEIp9cGMnzg0jLYMHJdyWaePSerEtT+Ofs5Dnc
Srwge7ZGIqgBB/PdsUkbqld3u7+kgUWVMI3UKtOSfHKA96zr729Bgxgp1jZRDQnA
kD484QLcsKRVzsv7/ve+RiacWYRJZ0Asp75ZLo/8S378P6K0KR5v+RbiTR1pwoe/
tULltPcLWbpyP2QuqrHpchZi/jxtBQb88gTVutDCEJHiOcNGP4o+9EDE+HvRHDBe
WC4d4kdlxaJRzSN6NhJ+rcIvfFzuguRdiAzS+vTd7L4AlvafFOEv9C9qV6RqUzUo
DAI45vBhdh/WbcN0V2blCOMwN6ehhsiFg2uEvTW+vZaPDhRoH3uB28Zoz18darq0
w0uaowpoBxii7S1gXI/PDrwopJojB17AUWTAfsPp/RR1IammyPlMhCo8USjOQFvz
Co7PpFMLwAIkGUQRhaJL+5RU4l0s+kcoPBKPbIEmpnHEEZD/amuCcwYK2kixzRk6
KzLSsM8oakkpiiQKclyhzN5Sf4/fWRp5v6lZ/O3uJ/NH4KbraAA+zFMbClt+K/FO
xeyC6zarspwdNK7+0mpVwUEYZNAv2nFkWSp4wWV6wL6nEBw/Xvgr71ITh+xNW1V1
0inDdCfp5YU1N2Z787YH+WbxxiiWwO2+BmqqxdGHSFszGPzfBbNgXD78qdOdZY4j
z/aoF1zBuY3jCTEfl35/8S0xKEDwaW3v5q6dk/JzvOWVP8NeskwM7vzX3WgVDIEV
YdyvE8PIWAy/LxQlW/lXuU2eNr4XefJJyo/OlzCR7QW7E84c/ToWrtFGxJft/75P
OcnVL8iVZ5OvNgT7rSLBWq7aAUuP9iaf2ZENrJEQn5SlrHa0OFLRcGAWQDc0QLLF
yNygsu3aOwxfwRoZKB6XbYBkRlIvJwhQTnJXMwLctP9/X4ajBhQJUscKULSwlEb5
OKQ/o31klpqNwblVFWsMeqjgbCiroPvswQLd4sJVxCfxYVtftcSI/PO/fVVwH3b6
8Tn5uLO5ejSkiJEOfyp/UCglAh8sC85CwoQui3QPv9jUqaxCo93xPKQvbqGSQd4m
25Tr+QqusLAwUJpjwQhMuR0K4aXyxcD4CbTHh6Jp99tObv1+TXopG38eindeBGgi
KK9n4agXYaI7UASPd/KUSIHTUEnMCgcexDZYTOG07lRgxgbczAaCsDLZMqSQgaeG
eLMobNsRcMheK4QYwSbrO6G0HfWyYeNGIaaSXTIros0ysWMi4+kXo0gKU97+smER
f2zLzrazooPOzApmYIZY93yTGDeFwN9JDz1HMfkad+xEuy1V1oPi6/J/YYxeMHS4
tCIQN7hPFJ9QGYQ4xFZGl4a5n3wgJ97dIAAx25h4hHsXqAsJ0jzigyzI23xcI37O
qkRvgHWwKpmQcNul4waIWay+DcR0H6/5xZLSNN6q1luS9x5M+zZ4zNgXMwn8Ospk
0tgM2P6Dyb00cQaqJZsaVLz3v7fo3Hjd8B7l0/7qL08lVXVvtBJP9dSpgJFgwenm
VYpEos9C9Yhy6WRpHkXYRGEBw7CDgumizMq8zyN+h4DXSc/gkw0lBuyXPFB/irAD
C0YRlauxxazTbiHNTUidtxWwPObZY0lUsZyE9wvSz6qcnT0aSms+KeW1EpvMPQ0b
H233Wf/Qdw0xkBvIA+foIIbKf2GzVERLTgrRG8slsTHYrkUBPYdD6JTLs+guYZLL
OKi6boc4oEcZRDTPVJAADE8JPK+79xDUMkeEWd3RcV156dX4Zo9Irtc8T4I/xUmJ
V3ANdnecvkB5YntgGBqvD579gLKH159dgTKNLMtkFtg8D+JdcPDrX1LNYsuenRyF
5MPGSIAPjzw3AHe4128Cv4BKL3NpvGbVlVVjn9BTAPYMkv9wNEdegZEC63cRD48J
/T93qnhs2Eh/a4vg/WNjrWn8mP/CspEJf97P6o9npYtZnwT/R1FB8LRdcImbpMzU
ZePHH+QSEdAKsPbRk3PChLt1tmZrOlm8PPASjn31vz7VfeUYfDhWiOFOudZQ3Iqj
WooGVjAFLdgPUjZToyXmfXCK7Xe4mB175dctVCnc7sdp1s7N4GdPkLdEHiJig56w
KRaspo9Jwbns/uqS8kHu0XsrBmP+K3YHeDTgJ/uPeg2j+fixFPTSYtViUJjdceWP
rwVRrJfhSOe05f4IF+tVNNkVObfUwgkawyDPAXr1SXFB6pKD1SD909w8RDZ6fx3J
f2mAIwX90ft99A9XGwgHXSOsxigkQR6lpX4f9TEWmm0kZfxUMggP3tR9DFSnUwpY
jcukWlz6Frzl/O+KCzF3TZPiBh1Djus0iMs/n9y+IpQmQ+CwVoEXFQkF+qT73Ye9
HS4Nkl3/s4OK9BJc+15cvZeiHQ7KMoMZOJNFkKZ71vNhn8TuL5YfPbA6A2uXYDwl
+TYWZ9wsr3yh8lPrt7iCcjM+RsZF+Gw+I2ae0X5pupmxpHcDEQhEo8qobPYWb+Gk
SyL7p7ORd8qFhkcNyeez3Nw4D/tBnvaJBOipPJre10wMOdv9opPxsepYF8x8msKf
kgOb8W2yTo8kaGbEHuHEbSVeOLXJM5HB3LpG2iCSshJ8QAIehAV8qlAPyNE4WT7i
+OYXyyoTooSRDNoO7i668FCaPbjDQq8xglJ/wQE2JnCafPhOEJkO4nb7JadnEOXd
+oPnzl7QaiKqQ3IjjzLOWtSSXBI9GN8rdL8e1Z605gliaGQ77ULqZXM7cK5vrSR9
QrsVmoISMtsQ5ZrzA1nICcxBSFNKox7KZAgkQyjMLdNODX9LN46d1Kw48mVXo0tM
n6My371PoSncoURT+8vTaHzFCSevDnmk/11tGTvxkbfhz/K5NTd1mVz86QIqDS4V
81WhP18FZx2Df0tDl4/5LKm1gV7jKxrBCVmRYUG4BLY5AXDPfNajoK117QfMOSr9
d9AMatYePLpgLqvXYqk6h75sugz1fCMyMOOqO8nOUlDWclGuqmnwoYg/L/5VC1E2
mFWXfuUYPpHOnfRaDY5/24zOhMqkTrDgpC7+/NELYgxETsefaFyX+gLVx8zUibsb
3ur/A3TfVCqHsO9VCuIGB+jyCriqF05lVgBKoBBRVIYp35UcC26MY4w51TDPGykg
48qUv3JsvULWWuIDalID/eBeyxy3bRaPj2FggYMgVuCyDst30wpus1UUzsN6jljG
NieoPoOrHi2Sgd61I6HXGlZeWj8CPHjUbFG6yzV+qID85jqVZ2AqRrFbUrhVxVf6
qPJLaKaSSYLEp9aPpYsNkqaHUDdA1fjq9pjcI6ELp9xWnZM8gbJAxwmNpwq7Z6YO
pJOpMPzlq1Nsh0rZn7uugRTeb4MkIMYg9zKohYKcN2OWw+pK0eHehVnhPIR1XavK
uQ9b/Yp3dtZXtIQOGOjNVIRYxfxVgDerFQ8yxju2TsIVbXg/nR0M7YAO7nbu1/78
EhPhnvvqxe5xTQ4rjrW7VHbx54kSn09JIRPb4C3TrWrIWXdxUiVDqk72Ja3OFxjR
i7KjY56lQonDH+N1kuuNlxORlh1JbrNXa+j7CtmhWdRZw5xuPMZACG75vdkm/qEB
ZmMokvMZVk2Pn1OB20/qXwXtIWDOHXZvJOIOCnnrEJw6O7nEBMHx8HEKPLnnVDsW
lEYA+fpSPzwxDLxKiKF9iUhySI+TAQaBiU/Nj1BjCl/R455Wj81wSZhPdNQmGCkk
i+2w2BI8nDRCt6mExXkT7P5dVrt0eHwdYf84gxi1mMDcNytBkgjidYOh+fbesfHu
PmiOSORW0zbpCs9M1u+5Kkl1tyCf1VVL1HuVnn+Hrx5nfFDM6eXQu5BAgxIdFSqV
j9so2nqXx+KdZ2lE+yHeR/pRQfVVec2B78zdtfV+L0dzGkvJavlhiFCgvvAOppBD
GWZL1hqZOoETqIIe9RWWQ7NKb/XRg/CrMvjkMS/WrZA4BrcC+ihX4AVsN7cdbVpg
48C6pUZet0q/6ryKur9oNaQTiB7DHE4FWh8Vk+2FMAoKHm40T02sHP61mf//KZYW
gEDt6xduNhmfVnlWpJvC82N0YnRaZWX9jYA3VIq9Tti/EqLHJWKeSszDwxU6K57V
YXVRDmPoFi1i+CtF6C7HWvND1hf8DXVj0n3lcCX3XkOeqhjvPFbcFYRsLfk0dsBj
H+J9tv/URs506oClwrdlKHZsMkkwp+Y+jYmS+n8EwdJr9doORNg1+QV0Yv34wjVt
tsUJQRdtNtP2ZArJbn6CGKxuNvmVMtEHjhDUpCl/NoXeqYGkIlG4poJJqr/ajo7I
tinkAYHeNt2zGNN7L0eFkn/b4MOJbzTdjOktJghe6ko2PkXUnqI7lFqD7DpQsVTd
EH6ZLKVoIryMZv4W6+GaWnJhdRvB+1doKvMhBf127/AMk927ZCBn0vkC3Wq6+Y2M
w/5f2R9C99JNgmbxiFYrzMRud3SRFM2gkMsu+D5YBm4vekLrrLvCM6dyj7rLe/UW
BWwxni/eE1bzFIpNahikbTgyetu1Vhys+lpfXGFSrjPXz6LPrQDPYSlTVYifw9EF
q2EKvhPstSk8Bh6NFWQ3xYIj14Ue0oi2u9Pi7y/DhdLpnBd44r0baEz1axilAGOV
QZPRBrVIXnNeNTXx06nMXG/D4v/N4gmvcUCzg/QrUWfko0349o80H1Fvbk092cUN
WTVmuALy1f0vhS/ZhlGtZ0t0hmLi6EDoL+TCEhMNdibdOhi5/QFWPW98wn8XfC2C
lib9zKFqme3x4X3TV2O+vS9NxHevSGElySbSEjdhBcwalg54tAuy9lrbdkiYWy+i
LATYtF+wbOD6vmAS+TcaMR/SA6QAeV4dC252eUotb1aiYZUHBS6YTk0ug7p1GpFQ
EfymEjOGWCqP7gZ+d4C3Qo64hc1fwNwtranAecXVoaUf/7vCVTA/zEZyeANFnN1v
Kdf8xnAsOdbOg7vzvY0MoBIOYZmKPlBEg2pGSdYI6xihnoEwIYxatvV440NtA2IO
4Z9XIiMKiPZOD/tlXTG9uFs5XbDhGCIc7DvJcx/lnC5rVzWxUGf+oV6dFBZf7Vc4
LFIRBdRA0uglCUpaAzPCLDoRktzhDW6PCztcoA9Xv8YmknBIhjxYyV7zy+9Zc8NL
uHK5vm2NA62wpv5HEDGsTGheIRPNRgOi1b1yeaxLqaBC/AXy9sWeZed3DS5hN2pN
uBEQbjMDHqzTUYtMTDCxKMTyyXQdK1qinUA5hq+juwenDq5ULaYJY6aW+LJRrxCY
VSHhTmLoZsYkJiy3J85jQN5ywa/S1PP+Q2ziP6lnP/aYf3rkms2wqXekyjU/vN+H
g+sRiNzx8dKf7I3WS9j2iWX5vHOIP1Vitd0XedhFKurMsELv22hDbXr+zOZpbfOD
zZW/mbe/j403+mtkC0c3E1uLGz3Upu3hGiXkuFx3dXhO+6Cy+Tg98KPipumu5nwS
7rFemap2U5cojiA8G+YlNgsYUCtuvMkpANngH6lisc8vqkWapclNW6kKVs+XG4Jj
bSpehS9ZRPyWP/t7fV6Re0k8Uw/xRccBgvu0Hf/W5YJRFVmG+kSog4Yx4FDrFbJI
iHArVxE+TErleSkDTUacHwt6NkE4AGFvHD61/bAQB+bmBhE3O4r12sPlTYeZZbNm
ibHxcMZyCnyZQvbgu6by7JUq7otFtElp9SZwAp6T7hpjNLeixcB3wN5HAaCOvaz7
Tv2a2JvAd/MskLqQF7gRNhtSPcMFOhE4hEO6uKJVlIdP7pl1l3nZfVprJpXL7e9W
ZWSAj8qfVueQjUtnSiX5QsJix2P/hMuDOEoVwFOlxp3rPFSqSIAiFjHHW9/a0nvf
GrfGrFlJbCFHv/POxOa8Yf7O/1ntjked0bfkkXEXdWnv7+0gf8UuVOd1PR2xA2P0
V+RsQ0mp0uG4PcMrmbwxrjwZNFB5uy/NcBCi9GbIwZK2ZVUypnZ1kny0Y9OwRcxP
5PknXf23Xds7R+Pz4YyAa5FQqIgeZh4w4W/XrISiBWYYQcUFe4HJ3ongxsvvzsFe
lj16AxO+u+6qCcwz6EUFF3UUOCqayZmojrUaTCDsQq56/GLf9IF1JSrQVAjw6E//
d0X/c3xSY7/1fjt1LZwTkAR713Job/2O9/I604rFW9Eir5YdcC81hhrREVk+1ylN
GFmxuaNUT6frNt4PpDRhW7Yg8dOZ64TvbUvQp/B/rQmMGXvRvzF9eDA2psmdz9Y1
8EItcVs6JYA9ApQdrvVihU3dXel3TURGAiKZZBTYq9RbIbAfgi25xtna/Wa9+W2V
SsncpCaxeSclHEBGIj2gyWzAO1yxjTRzsyEhnDPuMPrNkU0nJ1bQwbaOStzZVyzO
ij2TXy7J7w+XYGTuLwKcluDBcoDg7J+8RKukeHNJ4cVOQ6jc2wSMqJXVXlui1Atw
iyH/QArv67F5v1XE67xbInWLbYubJdayl32RJLrlJ3ToUYdnO7ZoUrfov3SDjBew
NZMYYAGFCiLqAzC5A0KaUYsTeOSiXKUgUaNKo8UCeCz0bhT5LY6GIq5MKtTgimAf
mEaDQztpv+Zqx38mpWx3Z1rUeGC0iZbdqZtRerSsG8X5nxI8fLWcPu2I5L3LtN0+
EVnB/yY485JV1nR7fVQ/b2ZMprU+0hqaHOrVrT2Wc5NCzxeq4EL2iMqteNhEc/jD
AcAW+pOlWKezEvGO2wlGA+QpWR4cnU+rh6VCEXYmPKtV+bCRqgcQrc2OsZm+x7Cl
JUGaV3GEzhGMvoIKz0nYyIrau7TueQMAJiMhNvMSgy+Jj8KA+eyRgxIQpy31kqV6
96r2kZ5ysB2fPAGvv48RFlFu2M5rEG9P6nU0hwaW88zaMYjved4G//guZ5imZY0r
dObWi9XQFcAudib9tgDF0wsVVWFJWQiw7FxmZjsrFSdBnkIequnqlWvp47n5HVCN
UlO4NHlJ2DZy+NiBdKoyu7b/iNRtBwnQOq+02bxxTMQP/t75Kh6MVviAvEdj+RS5
xWl8XrGYpXkD2ZJyb9t7acv4ffZRzIApK1sMxfXn1/WBSVWtn+HSqSGQaydB4MSt
z10rsbGj/VTlcxQ0CkkpXNgvIWteITVWgvOQ/cSYrTwaaNtYqkeFcLYlwHobSrq7
Toqwj+1Bm5FXC96hSGa0iUN3kdF4LOhmn3AvN1zXlDcU67CRnlwmDxEoL6iiFbEa
AIj1k/eUI/tiREYY/KtcfU7VSsPck/i4Myi/MfFtHjl1HOm3h+aq5hAXOEvpfbCy
NpEa/Ax6Ne/il+5A3h+T8FAcIW/ujyfmCdJzeLaxuyMP/BMUVf/Ry/09WTkABekU
wv8lRE1h4akM43NDRuS12/w6y04E7n7SHBgK3ZmRIao8L/fl6dSAX4ZX1xNfUIVf
8JNm/fcGNdUgBWNzH+cnCHsBrPN27UBbrwa0vxqWKQ5tt3LfgxLKeIuWbkhBi5b1
qnmJSiuJljIbLpV59nSWtk/Om+pBCf73qLd0Jc9TUx9iRlkEujJdXyCgoBk6R2v3
OWOUvDtBgRUYxTv8KkZUk4rJfL/uGintC1VswPXSbcurGWXfFfPP6M6nMLayMEYP
htgchkswWxTvF3MwwAS33kdLAsaWlFkOheNfxHCEklabPX93O997V6nzNwgdkAi8
TiHaoYnf8T+nAwSbs9Ee1FWlLooX2EKlhVQQB2JyhV/msVkvMUbxN9+JQVy+LaGS
bLXUKKX6R8YWMrDlmfmNquBhQlEJrJrJDwI7sjA5yTIEMzdIAKpjKEEeEl0uuC+H
5jzy+IBqRB5cKSLW97QckAMzUdu0AulZCOG8S78CAQnqcBXOy3EjzR6jNTHbPHqr
2hLIKXQ8VBdcPa2DpErkoTeghm8xn1Kzu96tPZc8Vilg6l3pKEqLVt+aMGJ7aMsk
LVH1sM/LVlGOeEAxaSwteDHnhFfk1h94GmkNRFAlrbA1c5M2y6iDBjLarmloZVia
cjo1Zet/bGjrTwlkyyBTUEnqnPOtD1RBP0bm54TST/RhgwZz8fPNLO6Te6mNHxqz
hurTzRbBDcthSjugfN0JkSHG1UODcvtZFngHIBE2Xqur5r/PtMA+g3Egjw0vT0aa
St/PKxk9S+8goWL/1YPI6Nr9UOuo84E9BdipjvTUW8Zt1a05v2OrbReZoshiWBPB
3hXYIOi25u8BtsCSfKfjisOQaVyuFZRjW09F1ZyCdTV3U49y/SKIbQd/fsmEq8eE
sH0zGH9hpVld+vYeE0baAcCgZWJlguWcs1UsBSfEFpvwSiwMuc+BIOWcCaTN6hQc
aZ2HvuQSCGnGKP0eZs3EW8uvuwVJTdxL1IRIwwiSz/KLOX6sBJXRctY3t7ZQ5o1Z
pWZHdlbef3BE2w4g3j3lE0EMZerI/LoKCviKpSaQ55kAnvc6ssGKYL7bC1cjkl4A
rE+4qRl3tC3spOAekIH6FVtI5FEimfY0dyuxq5rQ/SheheAP4px6tLKX8TjKLKyU
aTUzdbx/x9Vx8CHRMOf9n6Eet2L5w8h7nEmYSuBZLbXaffIdSvphoNMje0562T4z
nX+4/ihWTPwKMFQ/Kb3C37MME00kOQ2Pf9r+sCvJ2GktqOFrFu0thOgU1F3ouW5d
m3GEafip7MD5hGaRxDLrzaGZJ2MVyS/KZ5QgrHduVkbUsSRHwPjUJ26EMZNqfvre
uZhf1gEM+WM5GlJHtQ+Puh/FtAmq3OWVQrOPtcVvWeW3+6NMbGukqf7cHDVJMLs4
N+SLkHl6wRMZ+BK8hUYY8QhnHX6LycXVS5SL2irHMyG7wZLMKziB6FGLlvjC1t+z
ZgAi5Cxjxmi+3Zl7wl+v6tps4Nhju9O9WGWWBk4suyJX6hwzOVNywCrBZeNsc2lv
pXHeiqMfqgIyFwso3xOY1/NCMHsYcFKcw7wUXAOGRbtgy2bixE8MXSt9HevA7ki8
ak9XW53K2hD1vQ4LfMVN4/RYN/LxCr+jXNz4ZpMWF8YsBFFKWlLSZ3PDEBwZje4I
bxiKVDVI+lhHUCZBBW2638s4p4mHTLuq7DfewGGlVWRp1OOb0UHBXYqybLAIrFXz
qa4CrvuQ1FYx0sHYXBSIwB1+arUG+vhz7x+orGOxGd+kJlR57AaZ1i4Dh+5UjXRT
80e6ymZkccgpcb8rPQwgMbSzP8dk1As+K9ayy9XoV4SJxJANWh1fCI4PBfSB9O2f
UBP2c6iTFafAHuKwR3zgTq3lad8FcB9swSL9/wuniFwwDpIimNkwWNvWPGP/+EBa
mW2H+EgBvV3QKLb7iKDSXEczdgkM9cAzsC4hbzI2o6CGkQ0zhVsRmrp/onlOnAg+
bcEtv5cxGFxoHuM3SKtaOoTFPiC7czVGbx7EwSgXrZ1jUj0eIXHxVB3msgOSoNsH
IoYWWhKNyoxaHbjiOlv8syw3Azh9xEOXfNIg8EVLfgl7RUs3Ls/M8ia88lsXHqBO
yPldVZTAPFxOjKRT3mqtYJJz6IwLk9ZabEpIC86BodapuW/V2k8DhKAsIn+rB6zv
BCeeGDb8WbBktXymsVPex/2n1sTnwb0N1FhwWHlGR1Z+ggcgOqjlxtXrIwbjPNSH
G25UeZyb8YL4+VF4U2Go25qjNeO5tDFCozs5egEHSxfbYJSQp/xqNuEutChy/9Tx
CNMRweKBr/svYJHf2BBmnlGRNU3naoeOauQOViHVeUDmMppmpdWKbMJDrbhndTD8
fpbDnFBsWvlNdiCyTfaAMoHufe8Bt0emcrfSQYuUGhOPAh3rU41LSpIiK7eg7I5U
N2KN2f0kseTeiOvCD31/8OJqxz9ZicvaOGe2rglVVOS5jaxQmlyZFmNDR8r1WhdZ
ixSLL8Ig3nbSjYpHDK0y7bdscCGQRGDncrrF/JAuMvIdP744ucsyR5Ph/JAlkjrj
a8/Nch3d36p/kWym+mZvr63lUouDqym5EJd0u2lgvDNgYd7xA1b107cNF4IGs6kt
LTvh6pXIHOEYF3uVSPc9ET5AxY7Dfh5fyF6iFdJATzAzXiF9KjWF6WvPqDgEcgDp
t/auNOj0OwDCaD3JHZnktfOh7J22A1a6Kucztm4+hWvhBz+PGbswbZ9KpDOTlbO1
hayw3BkzDf64X4Q76Faw/8QKXBAAOgcLcXEpyad1j3yMslP8xwSiiKuRwrPZmCoh
pt+YmodYxZT6t2KtwI2Wd2+kHAT7UrteVZ6DleO67XrjX8/Qt/eGOIkrExuy5QDi
GqagAd6N4UsmOyYlMSZKS3hTRxMV1j57VSXO8EUTviF/AkkosY5jITqj5MqMGrry
NdkN1DINvImFVZPWwdHK9iP5l7CteWGp2Gu9ahkBhGMN1yP7z+vl2jpmaFafpoyu
5KiDIdpIGKOj921Jrf4YgboQ0Foh2DxU02I9OPH21XxsBhxc3NziZNo905lqiD6j
2Nz2ouZEEkeX78GC5WKShi10W7fm51cy5VchNIU9YpvooakCf9/o2Slti1LOQOdq
jNChVCSn7XBXhjsxjCEfsKAkE8S511aiyiKNAXs0z0Bs5QX/UGRCdZh2la6kSVmI
9vRQKatHvsqJteP0iAFqdlcFZFOAfVlqILFMOPb/ieupzvKCAuvDz6uKTi49Nars
GXbw4rJ7I4zHfWWEB/DNldF8qwFE+zfisyM09z5fZQ4FZNl+UJWKV73Ahqf/UaOl
lSLs8PFBrqMGeUxMn4Ag60zTDeCz/auiI7hi/x1brqFYw9379uGUc1pNnE2gScjM
WytwbhFFLGvXesuKo6rS2g8Ne/+0RGyDjLg5Uj200yeKecALWqV8APQsC9BHoCNK
CPuB5bkqL4ygyva9NGRGCfunOXe11f0hLXiQs3ZplA4ZFlrGjPBPzcJkB1ylb2FM
tKyCh4o+umwg2a7v0Ko8WZOMdwnjvNnpRz6yu10JHWyeJjwgkljlARxkY+mujITZ
vLvh+rVrZ9onWrAHHi7zhsfjW+dmuYla9AprMpaAd3wdBMU4UeB2s/Ptz/yRiYTj
8bxW04YqAwGQ0FY8Yh6IyFo3s2k9oJQj4YtdWWkZw/SLgB9TUL68HoKISuYZDYcS
xYAZ2aSYwZUmU2ZbDL+FrnVhi1BvR24UHy/hWm62Y6eAMhfFcB5VYDBILfbkeb9i
Ag7DQmMSEEJk59NSont7eCCizzqOciL1434mY1IdIyozcoRcyYwUYtGaR4UMKA/N
jOOkisl8f40c8Hz6ex0YkzJnK+8Xi+uP9Hirp1fjXWVugq1gtcknqlsQiUC/wy+B
dNYXDtCuCB/mVQFD+rIUIJJRs1/dpCagtUUSGy+hFmUG732QmYp+EHIChwqaBdPr
8U//c/gx4EwXnw3K9VS50gaAyaMfW/SuwVpIJHGGtUakhXyu008NoGvIdPm4xTO3
FupeEacEO98YAGGBE1+Xu3W/sTdIOAEPKI+5qRgs8foCSpaAgD7IPMBKxzEun+wr
U/ounSG0z2eIBiJBAdsLt4DkZwOky0QQYw+C8RGd1h7Vh6ocUdnlTrCbcvHGamtB
moOUsHzgp68D5rK1IaiGhn/KS5E+zVgxMRPSiY5RABWAzrFhNG87w9igGserDpPk
eah6wAAsJ3EK4wtgwUH3OCEETJfhJmQRc1Qm3fTojvjAwckrW447fUaug8gScFqe
7EWMHANFgsGZCQIMQgXT59RUnh2cr56BTAANZ7souKsbWnx9yj6uNRI02DSGhXsf
cYntKzo27brKb3ShtcQboeeiyS3iaYTDwjBgzBaRKvKJSs+/+r+PvURTQzeBb6ie
dJKXV3jZVGcbZZn/83O5w1nT9EA0f0YUZOyV5Aj/Qe+GkbMpT1wqbCHyClUYXpbM
1Q1++ikWhzSgtSCTlISfBkHweAAcPjQweObp81ja7WtkA5mxsMKU/+bMjRT4Fndu
wN2QCgw9Ul55UqCOxv/FJLeTM1v8V6jFpWDcgrrk/mjOWQm7HVfdbinKWlKOdULA
lr+bR5NS6n1ISc0BbqLShXuqplPf2SF4+bHjSmek330L+FaHSkyDtQTfcvE4HwTm
bE4z9+VVQ5NBIvaptHuN4voSj0VcDAUdN6RYnUm51AgYSKzZQgwXeCqoST5gjxwd
LDtVrQcoP8MkUy4MDsvwSjmJtdFkkGAYXUL8Sq9uASeAvyaiKEdOJjSMWBDTmciw
zQOxOx68AC7wqTXss5b+0lSMKE3gvTejuP/Kh3LATc5Kd8w5EhJu/NqPEOgN98WZ
0klbsVwv/iwzdT0QYf6KGLIA9ex2t1J5xeFAKmeDo+CFRSXVjUAqGg/AdVBx/Snu
YdjL536nlmCHBTVeyJhX9agMwVxt95JiUYyUr5NYErlchDdkNGE1GHr6zx6x8hbp
j8l7sawj5RzSu4OXb8C5tWyUkI3dXp8agHS39iSHsCBWRHLMkVUvKdHb2zDYQPDf
TujntaFiNdQDy6bcawIBjUsWelUlphT9yW7nM+JPJHa7v5S8nLePJf+c/OT11tA6
f98Z8qL1ioSXpShFwQeRz34/Pbe/H7l8kl2mZcsZg+Z1nflK2GiBOci/B6xiBuyZ
snjFFJjd4kowb5yWZMDMEw1ICUKChw9Kw048/hpPSFGdRzGPd+kbb/FY23nQrErR
liO3EwhM0jluXdYD2M4caZJ+BD219iSQGcgFEyOqCzy6xuHX49f4sReEMA8jOEjI
anGIpjyY/WqHMYtGJQivuKJFlybCzEAgtco8ENmlk0RCQAtFmbv7R4qCYXAgAo1o
pq77p3qJNW9vsOBuMMDJQ8mv1aHDZDC9+tiyFR0+zerdZ4l+CW/+z3KMUrl5sQTs
/Z3RB9jlI71/ujdV2MZryLXvtX5vRqv2jV/RN2DAjYPON/ygmlNfQwpfPdysyJLz
okYr8noT8ukX+GZ28e9ne2XupPMAq3xjpZWnudGIvFZ4lby2qXUdZLD/MQNd2ICa
cqGcwgeo3O9mzl4NjiVS3lP1Z0153IcXlbf7NZmAcE0SPJxFYmVXGpDxtiAc47ks
b+fp89PofqdjT3+SMiQ3U+N0rhTEQTgeCT2ajn/fGTyu3XbFYgJFMnnyqhRI+nHG
01QLArFLho2zarwJ7y201jNRinDvlIxnwd1SWlQriwQfbgJrN2j6MZ4etd9XVbJX
C2N18VBp5J0yNK3Tc3nWGi/NFxtgwV1aHf6+aofPwwbQyFpWhLKmXYB4ia4FG9Yg
NuAKTtCDB9kfWikRHfcGW70aGUrm9jKiH//KxhvDLl7l8C5yEZZDbgRdORp1FB1t
GqW/In9LkGJen6ivd60fElS5MHJx/KIll70WbMjK5Y7wz/cLc5QeNbwpuVDwo8ya
cTqW5xf6OOu71WRJLVJnAy7aocF3uWH/EEELi7lwcXXMs6sonhcbxOFaDXOv5nXI
WPBatEwo7eBB41sj67d89g3r+P3g2gu2w22n0/63z1QAIT9Q6Dc2wU7K7hE9X2zG
DdVF1kOeHb9HJfWpr4CcZDPI05oxtMF5GVSCEfyOSu+DPd4kr50MaR7T3Jro7ymx
nHuy9Rwa+yKiMFdFdhQrO0AgaCue1pGxvzyDJJzu9VIuTgVFUDylU5A371Bn74nd
PAaAZmF12Fv45fW3ArEIsdp51kE82yPXnqmXKRkz6cuqcqK6MJ8iL9ICXBTG0a93
X704JO59aY2yzsBGlr3z1lkofEnQ6PnQAMo6xyHgB7vSV8obxc5+ttnlS/NXMhDF
sbTLmA4bKHrhkzqW7wKGtJJn4fijKiZ1JsheRLzkkTmK2UsSBY0dSk7DoIq1jnm1
vgEMOyjN3nPL7WW9pwqX+zy3UityUTVmJykj1Py8WvMJkYrzO9sJ74Jy/Kx8IAbV
dvu7BrxFcSUiQ1OHhwN2RmF5hdTjkCm2Yu+PGI4nQclnfrGRAoQ0oaRM9K1oQ1/f
se7iuzWQ/MGJCqQtZ3UhriUYv+S4gEGGnM9fxtSYbj2SU/mhwkQ2Kj5aIe8rl6Re
iCITv5wzQs3jGDMJx9lHop37TuGI9A738255OrJBbGtiURGfUDeJR+g9sdCKZiJF
0ISR3wvC6eW8PfkyZT4N+L701Bozzt3Kv/m4SM0WVTDjUo7rWeuOxVa7YrGtq/9H
Rb8k98/75eycyGBrHVNBABmwH3f2RzH79PUe0xrYgR33PFbvg42vlzD7l+b3JwqK
rBDw8KzQoK0wtNNMrj9teIV5zscl0T66Ihxq7BXml/aDCmyGO92HokY42e3QSEOl
a3KMfNb3BDxPPDEBukujfa+PP0PrYEerlma+hD6CeKFXej5mUH+GQay8FeAiHmRN
vp85zmuKK3lCv09fNxc7LCazs5H0+7b/CGfit0FB0WjLaEPFwJkR9fVzikYifcHl
qph7x8tCZ05dcnHxoc9Ey6jcq6QX8IRgcepz3LSxabKjKstC26a9hB9Bw/3BTT2u
X8c1MR59i/Z8pFiJGzUcAqqJgaT6yJ3MfgMdOP0WCo1l7U/chuE+UJucOy40Pky+
x2jkHiL4JYrEvLtOsLZwdPI1k3t8I1vlammHfPiJkzcH99svzEDdq1M+m6/dNFC5
+XNPdAej+1L8W7ETeC4WVwHy9MmDVgqczWjoxIG1SObwNn4AKvDShvNW/u3xQDN0
r5y1VBC/4ftHE+4qjLsIXnt5U1fIgwSS4Vj5idz+IATs6BkLX9y4jOipDRv4SEYD
Vc2dyPBbq62KTRnqVU1jxbeDcwVvUHTYmOnXmyG6LD6lRwUDkFdWYT6+QcAbOIK4
YWgTz3VZsdKlv7HJi9GhNttT4W0uW0DTWULxDTpudcWTq2/Don7bZPws8urZ93vl
e77SAwuK1yBp7M6ZVSPEcwqrIK3U/qb6FDvwGp8Q0AIhjR8NMpi/flWiEtkkgPoh
D3VaFzxZ2JI/gsvdwqDfwivnBekXWuNSDge1XmitEKPGSQPe4R975nUbLcWGL4fr
+O/k+kx/qEOelfFoGNRgNaWnB0MPtvDgQ8y7cB3L2CVuk3C94de5Qi/wlSwnAI+m
LuVeFpIWEvs5d3Qg1P7GHzXx1vDOaPmGrsR4HElN1WuqCenh0xw48qS2U7mfEAHR
jhHLhF+8tC/ipT18lIftTIqMtFatvdzFS5BdT2tV48HElMrFG/W7zNPi3aZMbxZA
uDNsvCi4nPk0xcAq+dEgmfDU8/+OC0DG1uCs1Pfpur2drNdQpq1IJGjFkiOQT/6A
QxZi3io48+W0OI4xqbLHJH22eW/VXV7oKOGPZAO/3+NiFFwzyjfTxPRJ6d755Nys
Q5VLF8KBakfjo3UHEw9m5KfowFtpRUN9xb8PE88ib8rxX+tYUKzj5C37aHinW39u
7NKv8NYAaWjNuolKhaCWCiZv9CgeCbcMDeu/tIpQZFo7VqeE4vH40qz9I1XGMNzH
3ed8iBISemxDlwqg3ayFE/Mw8sD0xE1AoRrudC/YTM/vKGWnopMymsQ4m4YKbdqd
nnp6G+3y6Ep86syR1S0QreVHDJPFJggpqPeuhtBzHzZwLBObhaZiFB1Tny8GUDo8
JGkejczXiHM2ibUWSHlTpsIcLIJ2RS1iTjb8u3mrQrg3pNoNGysjxMFIjHdv4rKz
F2KPvdbNDPHEk+xPz8dHtUWbe+PKhpdp6Cp05d2QdhQ9venrSCzOj3jsvnr/8GjL
9p+d7VbFoCgeHt4yc/bKBNtqfyZjNxOxw07RKpfM6y67kKMvzG0ExHHOdjKH7dD/
UpGchiAIlXOKAreOLGlaVuFpKVCwJzaBz4ZCWVnw7zsxK3EAaH9gXr0gnngiO0Gk
5WyvDZT3tbhRpSHqRKahmkMkzgdsjZD3pHJRldfs/O0fmzW+fQwoX4IPAjaNMyAj
3X6SZpr4/RvFGcSI1HXzdbOZgZJbcpsCR91FFd9PZzu35Gz1gq6QCIIkX6d6IGSj
6jQYA0uu+BPYgRHV4PPSNq8h0YJ1PN7Nso35xe/EOMA7mDHy5/dc7ez+z3ji5SFX
cPyNzZ3wSHIrh3YHS1s/vJ9Ej1VaZOej0hFU8UD+H+G9bnwHPK2U37pOTu0nEFaZ
lahEor2Uw39THT9ngoBJ3qx1bTN2kI6VteGEkBu3uWvIlmXY9jwfJW001LBHOSID
0g4Y/d6kikFy5VJkynJMaPTGeOOjtxSb0ykjxAsWzcVBk1Y52x6yAENpp1fqwOei
rHHfzsPHNmTCjFAjXNppIcn76FsUgOw36VczfFjIgX5ZoVoBWtek8tR02O2y1jZD
U2ppMZS5tUuoeesd7g2bR6yXUjP/nDoI+aUL8QJPwAk4a44JDkXcLeiqbPW7mydS
HFTwiufe1THWywi2Lveb+7xM07y5bv56E74Rk+CB7CS0yQueoXSgyqFyhWDcl2NM
IlPG/P73PYHnlVeVC/+n7OHruQLYX9iJDcbLyIHPL7tuod0fRRNg0OW5C0Hxorz+
d6UkJJzvOf5YHyctzdnvEWW82GqSdZT0fWqew8XTCn7fdKArSaEh0/q7YBKF8Ze0
zGrzxvm/52UEclhksJU8hp0yu5d4fs3tG5Ddc8LdYVILjPzJEULOhRI7HU4chjcB
jGFCVobaWTpTxZDZs4aUwTlSlOuhgha65Pez/WWc4sG/U8sIoJTUkzrF/B4TbXke
IEIGvXL6erv9IoIdUSDtckD30kLNhtT3AwHPzSVjLtqspQh4wu9btmIMvHHoUxlw
HLErEvaQPbtLZwc4ZzGSbfwWgPlelehJdNu5e67w93o5GRxaZD4xk2781hZ2HV6Q
lVn9DouJvYs2XOZPHMpKT/3GOoRpwDX0B4BL+EwjCGNAVsqIvVR2Y4cKe7o3OdkA
4nk1B4TcjHr55H9Dq6GU39WFgkH+Dxgpa1PZE6umT9yEqV2/gOvDLyl6UbfnKxRC
NqEMeFHXYnb4Hyi/M5RDlFbeM/lpPJI9/9jNrP+am2xVHB8iQiq8p2HUzGsfMKHh
r+76LDFsNm5AK54JJn5Cz5b8UlM6eqdXuW7pm7KRGvRzEZQkPqU1aIuiknnjeFWV
MtiBCZUNe9cbWJwuYjVhl33G7AWuKq9hAnI88lF6gpRgPmuEo7gJ0QXmGFfV0wMW
fFp5mWryqzvxKKQLvk3Dp7bHalxWWiajov3369VC+s0CtdCdYJyyyg01tiCh3lwj
KTq9F8Vq2boPVoDjWeRu/rHDFoHdgCMG0tmCqbs4oLXHeYfyJDMpS2V2RCDtSqWl
FtWsfbRvT5EjIxBL5D08zvu+yipMceI2INMFKf3K49x/+DITlVq5ieEg7gpcWf7k
YP6rX1xVipBIw/pTzHMB3iH7gP61ZLVEMWVkWEbzkd+HPvV2q9ySg1fpqf78qUb+
0mOuDVrTktzajgBXbw74zvlIbg7TrnEQ07WlhcF43YrW7oA1HAV7ClJhACeL6gf5
JsFumLHzXHVi7Mzes11WZPaLl6gIqoybR9Rmtth5cqEwmFjCzYqc88T/d2NGPgNj
3t9wcAjX+8o/+Ivk0fIG/FDMVJBNvK2rPnrxFe3vOOmtjIdUyvgO+wvSqyqGWpOR
ZvOXFS9rmhVvGCUaK6EYkuYqIImFEoePiXICnSQxCNlqVrBlm7MnMbHf4IhNnK+M
odwNqrl+F2pG6rcgoJ/4SL3i2r07+fPc0fc7kRY+2rHzzzH1Qi+whuhPHmJqIo8v
HRSTzwsodg1UTJArbyd52b+FhwN5kGjRfk2kww+g3To2AkMy7BAtFlsms+ymc7hD
0qitqqaZzrg2c+FOcoPHfo/7wzTiX395XTHnMKRgakCPpQ1HfnDOs+beJ1TBxhfi
SlC3dTmRZ0RvSdNdBXXF1qka5XSWtldLs05PdEv8OkNxhgUAu58RLu5D0jHCYRte
jdxn+VJ3r7GTxMNdvoUiftIkP3AyOVFO4soDwkwODJptJ2K1fS/crYG9nXEngvPO
gHCZu0flAXnks6Wh8n8GyTcqWNp6nX9z1heLS/rLy3Uz8izWrcR06g5Rc8OuqdNk
V/DINzPY3UdEB8WbA2o/wmWcESzEomeZn0PlyVYJqR05w/jYlcldpn26nbbEOFco
kbFZl0oPmWxAtxGJGfPrGEuj++7dxmoylio4Xkui/DzYteYRa9k0caxyIYG7XGY2
sQ3nj+F3G5RjFaI+nCHwW2eO0jmkQNu9h8OYrl/AnBU578XVobAOoofgJuikgEZr
ox0e8weToJIBUpM6oNEdK1Vva/c6ok8QNv3WKz1P8do6qkhE1CZ3DDGnRopV7XbY
blOajr7S+0Jrh/VfAs9qjzcvmaX1U6/IOZLkbOXIBtkLYRWlqFPAjZC50NcO1RZj
aaIrU/6742yqss6/KFOPaKhOykJ1qyfZb1g09TjOYPnHnnggP2mjP3T5RQI64Ayu
rJo5VkgyYMMF1DHO5zX8l0zBvKPYsbU6GnrPnUOY15rbvqr6o2QgAJazrg9bVNKE
AOi71k8DAWRgRXzL+TkYTUVPQZUvsrIPEGIwZmmxO6VypO74t6EE1x194yUSNJQX
4VkwLQVGVroY6FMKjpInkeSu7BRCpzy5/MnYeJ2r6kxFZiL/fl1fST5EP6fPGZt5
38uvszfOTKMqARCxrqvc6augyVDpPDNumS8P1BHvPFrVyCdMdqdO6MF7hWomjPPI
APlzdsWEMWKSf4kcfn4Mn19E4nZRMCEskFTPAQb7lGoycL1ClxkE1IjNtN13XrKU
zpftvo0Ry6glLzU7nhEJ/t1jH9bR5EtntaGs1FHtqcHOBt5NzoJtvsLAfB96+XYJ
ZQkIWC938mSJTPq+skvWBXsltshr1LcM6ttPSEY8QyXW3atpnEN7DU9hqcI2iiyL
0a0Tj9hwLxrjjkAY8+sXY2FoHz8LXsQewh3xqbOkt6SEQCcaUBGMs43b0DKV4bSi
NYUXgEUNA0Nu7nfVwmbM+IpDEF9cuze5mbLA8eKsjI5MULlc5arbhaZ9uR9MCkJU
DkyJK9Zv6DtrIF3crLpxiU+xSYuIojFuSwmTtOLLvb52OkC6OeaIU8q0bixQwoF1
njvxzY7PA7I4Bvchxt77PTR0UU2hecu//Co2/Lhk2um5GjpjBgZEi3QQer+AoXvt
BRegW4KbwPkvbcnozGGecss+hMbJw+eWQI3KYL/UvwSytu5v+8yZGSzEnrCmqKKr
Q94QU50WlJIjB5dTxk5whLsTrJRanEeDs65rwrB2Rr8TKsTzlypWZ+tK02HPFz5u
EZ/ZaFSWI6j+CIxp4S3Q4Yhhc4tt0wZjkSdAsNhkxZ3t5Od0N0D2ui+vr/5FV82Y
T4/S4eyB0g7flwSP0pqZw/en1MROFnqCgOAvZECv89e0k1uVbLcyVwSJ/Ip0MRuU
AV3SL8HIFDWxqYv7aOwIYF7Q0KwuwkZgpGyKugBkrYc+k3e/jzOEre92747nafOy
N3EfJ327f3vkHt0KugZcECV/bnGcjIS9doqd2qEIiV5+/uQZyGlsJehs5WFTgSFM
USuTIn5dCeNaMC1ddV/wkL33RtqkivDDSihVMDWfa1upvUz8bPuuBwT3dHFvnnR3
Vxmzrvogeb+fcIls+qs9G/LNSjTb2ePq+NyqkLxMqk5ou0q8LwboyZ4ACFze7EU1
Kxn8K702nnr0gtFCN8usIfx38BdJ6hcg3fgNHfD+0ZIpko0iXmwpZY1xppysYp69
vO791M3a1I0FfUKxfGF3viok5s9gVa5qwRSfv+VDibO1+LSBlR/+2Eg2yXFrgRAJ
b0715Q9DqP1jNpNXYGV8Fu+Gpbj8J+UdkjwtgkaytLc/iQBFRW6oIEUNqEXAYg6C
aaJig45cseM8sDk0XZPuS6RAGhVpF0vOYxSvnztvhCq9UiicISPJa4+fBww3if1n
T8lLajBrnI1NH/ivtrmC86udJc/PyJu28tK6sL3bmNBAE/pexYUBPGB+lIcbVHwv
3EWnNnzJlQyeAlw8UlkB6Wx2vLognKiFAN9od1+664yqwoeCT6yQzjMBQLj8z5Jn
017nni4S98eRXt/zkZuKlpg2rZEviRP+dZpa/34JkV8PR1gaHEn4Y5jnLgDYWV25
nkrVLTUtv3YS2K/O6+Izc2j8COqJjB65jwMxtWZ79Q+x57e52qa2QlyWXla49Con
84mhtMrFc5eaj6ltGS4uIy4qjE6q9LiYG2bBiVRXTiDYnsOzv/eijc+VwLXh7hYh
kvtxhP49F37xHcSH57YFaMWbUn0MeP2uHoQkfl0qYKyl+q785NNPQv9OzAPMUwsB
IKjZq6DLVy4rRG64EFQet9dzyg4cKufsnW4bkdOdcaW3EZ+S3aLykX8UYf9/J2/O
9/dtfhqZ72crLqSwqU/BNrNSxaskqC8tVFi80GulpDol6dYqTH+iVdWvd3MeOnZ9
7YOUhXxaxCcgRxl57W4x4mpKK5IUkHMQjSidfe6VsekGPXJ+y8feTMo5Ppfx6MXc
pdifqIUUbjkVA/TkTWrZCuydxB8jEFFMwi6MqJRJ6CGTyaCaSniCfWYHDj+PnrJv
EzM+QQ5vYYrL52To4Ha7Ahgd1n5F1fuvfofCjPgRvsTI1upDJNwVt8IOz5b/nQK2
N6SNQ7UeATra6h0KFsFkDDbP43BnYEvROP1vlUqa/F0SFj4ZoowXySOvTKGQJ9lp
4MSG8N+ngQInFaOhV5X2pkfYl4mZZVuKdiSpsTU/VOs9J2oPbl4D6LbRRVTkUSCQ
DJypefXlgJWyOBWlj7+kVsFjdgcrkOdd8aC4kMqoz6lU8xR8niDZHmNAzcH7Cexd
zaLRwAXKIBUPFXp0zYkCYNwR3aciXowsAckISR9t8dK4Rz38ge/cQk5nEisVbdWM
PNAVq8oHOE/kkzbyE1er8LCQ204tDkR9DNj8T3wCkjINtrbqHVwwtl1HTrwf0f0o
chC6eQFPJ29FJnoNEpILjL7KhlizIFYFjlalNKaZ9Zg1Z2s6H0fflm77x6FKiVaN
GUPk+s/7nXe3DwosvdXOLR8qHp9eGgwV5caE3p+PR4+hT4o0nG+aasqdWrJXB1tn
E7gOZyNSkZbwNbkjmKZHPJFnAur9d9cts8bd0GVqM88WybC8Ixia1/buq22GQITB
lsXIe209JfW6rBjyxuxwOBDbRRqXwFnqmFwWxv2S7UDGaJrgTByFeZ466uNPEK4r
HfCxIhYJql01QP3oi82EQB3mgAJnDowJ4PXLWJ3ajkitfA2mtiocrj+D5AEurS5R
QgoM0ThpjDnEIVkyNnI7MjD3gZc90OLO7smeF0Ir29DuXlBKwnJ0CiYccaMUIell
d9AtbkaxaQcxFJJfD+eR3derKwcQQ+T+0Je49yvr40n8231c0WYMiNDSWcEg6Yju
aXusmv9N/H3VUJ2/e1oX40McaKtoUcOiOZj5NSPgsa0gmYUGY07Ot2n4PP9ewko8
4lGY7Q+7FpIb1zrZOfpoNkHGsl0ftQ2CrxRALErihNvQ3TdwV1WJWwkL2YYY/WH+
JrWf8DxV8FmwQS4c/Te68f7Ck1hl9iIXhrA5ULoFQbqULSqSNz1CX1rCXU78MsGw
neV/qYc4kJR28XDJmC8xy0lRxZosQYXrEEwqBLW2hp0HZnscNcjC99JE6hdsPyuH
o9b3E2QlozG9kkxF+6On4qQirvfu2IhENMPgcZ8MEsHjalFXs/pjzPkUkxZyMITL
Ctg1246+O0aXKugqcAMG1AxkK48U5tqKAad36TkVw0D+CKJx7IfC8dSxBmKbHsuN
MLJPCnI3fnQnlNNdXupr7Mon9eqIkVpVgxPoQCY/lbF1aTXQNW2p89Dr73qQewdi
7oIIUCsPcIKBS/5s+DkVXuqCLmGkn4C7ICfx5du8IcSwlTXxWNSTXWA9hQ3iKjv2
G3ubMq08tOM6wtmhaQaAmmGrOCnIM6jXuIouFcO59NcgxblajflM2Ae926kX6BY7
z0l7zbQSq2y3AITKsgaevZoyhhR9dUcUwhno2KdBPvDtQKSOE6GuBqEqsNH0n3II
qK8Dk3huN4DziB6pnkE4ezlYu7BEjnIYzOFHPTD4bopyEqM6av6BP8dJjFyETvlB
pDDJj8SqVQldUSUQWaPaZSE5Hb80bn6y7DqvY31Uf0F83mJ4P0yqL+YZ0c74+Gd4
xAgFuSFZ/8x43lU7Iq/JffMhkutfI3c27AI2GOv3XWGNzbiCRORDMR3ITCGv6but
59hDiyEtaddZIIW03CHwBGtSBuMPWqYATex8IaTdPAMVeekj1QAyCv4dKZ6JcLAQ
uP7+L5ktaGrx8Hm1Al2kKP+yLXubu9lQkNqqK989GBPNZRDreFwWw706rq3uxnFV
QIn+sSIjB/duIymbKv8+PENEhcUv5ovo9awpYbBLjeiEThp4lSQONjA32CcJUlFr
pvusE7nHCPXJz0ryCztePYO5rliEpEjpYMbzSnJH5a/gtE7UoUaUb6xF0HkHH7iB
OVZ2MT2fCQMLQMadMskNm+nX3yUx5J125exR138z+n8ruV7o7DvlkWLU/O8VB2z1
GdULGGJEcSubX8yftnAagKXNKUbZNGTIVNMW3HUr6T9U0M1WpXxNZ2oTNcvKtUrL
Z7BaVRDbu0u+LYUrPcH55mS/MqBRt/uI0xPu5isZbbPGpZV4OrwN3DOC0OuTMAAI
aAgXCBC1nWa+EsQAhIPxDblBDxZgPLgA7oAfMq2b5icRyihBmIoR1pKEm3JI3jfl
BDSOgZVIb83zBKQ0ZjwRtvG3lgrLFNd1yc3oGg1/2Ap5cNLfxitrpv11jZlEuI4V
0/rlpstHMUcssqDXaceRUA+wA9SiYoz8RopJcm7CurAp3+LddoCCfcCZRyH1/6Wz
jTJfc7zoAGxUofr19hIWSTRo9BXFjiggnnfe8/eyLkBwzjEl4qcDcPc+DR1PVHV5
B+YzQJKgHAF7mTyuI6Z1Ef50qnCJmo5LYJcaz8cA+VYhXaipCat6dAsvTyQivClH
Ft0rnTCXfHbgPsyTABbKV3EhHwr8HfxtQucr7ib+mp9JUV1fCcHziTsNyJDEbC5j
saL4V22V5B1YwjSDVcGN1aCvqSsu/gErDoES/KNPKz4FQPkT2DgFcd+vEMiCPc/D
+ctaOyzMrsEXACLiK+2oqM7XTfNRCS5QTtBcSLeLXCp2ivfeE7ZuPB9suwd0V8jC
DK3L8FaPwZB5wqL5nXyrJYQuzJEdougykhcfBtydxxjQ+wnbUKvgxJg0u5E2eLcS
vfv1fXzdClhZLWQMchTNdPq25y8BQk/uNSD2A7PLBVXsOF6dR3LSGz90YD2zk0om
XR3o+cXmxFcUujiR4p9YwtYLpiDw0pgJImpLW253QMhABiBjLbs5B2G758kKVzcb
rnzixjNQGkamwtvEQqDcwbdO2yd+ep/LxCDCzFXumGI5Pj08TsbuqEXzmAI6dlP1
Smizfvkh6AaaQysieUwl6yQAh7OSXoJt8ujJ191peQyPAkYhVUlOniSxoZQ5BkER
9FF6uvkkj20ruTNeCh9LuZSmppEGNnPHZJEdBbFTr4+Rs8uPWtfzMzcRBdgh9tKa
Ppx/UjTw+pztMNXa3tvnT4nFYVVkURX1WZYGWceHHtDkoiHbNo98IaEVTpUTTGnh
NQmmFwcQ+JJlic6Ivk5Z2SA4+OfO0yUhaTc0CJuE0JY98SIUdjMN40CfZCVlt0qO
ZKkwHeT3Q1/548nGRjaECbOuM9GpmFf0V1OwxQl9I9ic/CsOwHJpTP4Wrc5JVPVO
WyXLIzHwwF6JX6RtfYhrrtWSDUlWdeU5tK1Cq4sJZWOCd2KVpgB2U7Yn23dNbTd7
StfcR10rbDcXFWObwjaIg0J8i61JEkEj139Ym+gYhtUfnYWUvBGCeodX4KGsNoc2
peMYgDuOo+x1QMmmsUxx8DoE9eppAKBCDUvUqrGLDMz5NMr9TboId2tAJ8VP07e0
p3fiTeVZrsOV3UfzPV9ts+LeqnSiDEwPKH0grcbXI2Avq0iejgYPKDhg5Dok06eG
RUX6zQ+fhDfgiZAIeUdV6ryTLSqBz/I2Xmxshhz8pGRRJ2bHmYWUI1qAUy/OqLA4
vcrbcemDJenWerHu9A70Sj/aMX7KT12eOIoT2rR5TfChTj28sDtL6tmGGa/C4vZv
aJ9pirYNQf6U/hu02L1Ck/asGoLZh7OX/pxox1gDx5yF/a7ghW1z2qKEAAGXAkKy
w7a0TWZ6D/Rzg94gwJTsgqedwklcPhP0ukOXTBwFcV/NMA37bhimvnC8y3SsFG4f
yaldeG1V7FGaoqmOGJPS59CJrC1zFqez1Xo7lEwMEBsxdtrJA0wKN81ptk6jsI1Y
OStCT/PyUKIGivR7Y0x/oKHDQBPzRRXu7ViYs7pIGYfR6hbqjCvmLbsWqKprmXSj
6Nr23gU+tnowxo3baFOKcpPBNQNP8FCa5OzbOKZ2wzefwKzdxQGWtEL5PsmZyG55
wy648imCi8nbELIkpHSovjpyHb60xeibRs/d4ngEoZ6oJeLzohiRJ+7hYEeRvmzI
kHVNWGcV7PdvVJYe7XOWDN1RLpuL8tkTy5n4SviH5Y8xZ8wAExhvULVtkcg8YL1S
Y6PeEk9rYssant8AV59UU+VDf0IAqe8po7hDhOyV/jeDZOAeGa2QYshfWoWcbNbM
CGFD2JqpL2XVri5ETe9lQNTKvZ42bBe2mZFWMTpD/pre+BvGQupI9WJ8Isrl2wHh
wIoeTsD+5UeMMbALrynTJIxq82pAL+kYniHuzDcr+qg=
`protect END_PROTECTED
