`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRyWpcTL72/rC2otgji7r2m7NM9Taup9mAKXdE89kmM8yq8thZlZdx+yMymsuQvp
54c7P955r5QAcyPXFgA2bBY1k5n2EcUY2/XGCZo2CzlhHD1WxGPkJOAnACqahGsk
zwyzf2L7MsHZ8P4IZrRwGnQotOcDpiYUlEotOPYiF0ToNOZYDIq4m/zI+2P9t/DU
hqvubaBcUaLfrUx77NM6z/E8gZrX5hW75hDFPXu3WCcwvEcf9XgOFxyBEE1e474N
Ur+IRPWzxtagNgP5+x5IUADDGJU7jH/lQJy4yL0Pegrer9SYb5+bVL0LB9ScXsVf
0dOknVygob9Kh69qaSo/JdfUA4Wsseft8ro66xGj0OEBWpHIxHQmgQ7cd5jckIkO
ZdAElVXvrLxUDm/O5AM06wypXQxXFIlxqLwTtwJLrXXse/K8wo3ZDNnu+C+eTdsA
qYWrUGwQbSraJ1UHuxbNFBrd145N6cjx4hVwwSOL534ZqnzziMjEus06bog5f+K4
JchF3TwrnYniK9vFSnY9CqzSsgSjpZKQ+kfRykwNu9n0+nf4J96D29KsuS1WjWZJ
JC1polFkEgbThyArwle04hbnOkGU3RnjHOOsPa9mNXWK45SjlYSKp12pw+A4Lk3e
ghMOgaTxilJ48GfK8FH4J87dJk5FYiS12MUMfs3A5y1YZVXzA+4axs8ItLiO3jtq
2rm5LDspHsgqqhYwuWnafTZJVhBNx/umOfOmo6BvtDPHHv/6uupPKa0530NC07Hr
5jk4FMhrrrftLVbrT1rSd9rIi2qcvApBpg+BD22ibYpCHiiEG2+Nl7ItWT2he+8V
xI4rNpY4PuoYQwn5USFxVZIdwNTK+fRu3jxhZkB9MaN137PirrOGM2Le5VyFHGvj
m0CQH+0sB3aXg7l58Nz15yOduuySyr79FYYYC+FfOf/5qcYeLu9rCzVbMj2OcaFi
lL68nJzJZKPUACMqt9xusYyqVvB4u9MQYOW5BLGdSCsEHKFVHltoOvWBdnXfzQIX
miNaPnVi/36jTHHepzSy/8jaiVCh+bd1DcsIuAjVobcHHjx+69vz+Y5VU2jqhuwk
23FZTY3w8oRY25rwRTNpL+BC/Jea3RKfTai9l4hl0NKKIKKy0EJNxJd+c7VWgwW9
/1PbWrz18iKUJc4KDZJUo6B+OnSzGH0iwCKfz8jVO1F/PUGrKDTR6NLD3RdSTyqG
MuNBo8r1qjLaDyQkW+oJyw4qWvXbR2xryEjh4Du5dnOVjOGrvrHMaLUVZ+Ydua6g
k79MGzk8d2Ll7RWjk+X/EKWx9KJBUNHxz+jwCEmXX+lWwj+ET7lzlbOgmiGKXoO4
THVbcsO/1iolS59Ydnb+W7q8g2ewB+b+zSb54zHmwOMTkDy/uoxHi0CwmY3Y6sxh
7/TIMXKU+N1KWSTe82bX4G1D7K3Ouri+vGGS4YWYLll9I8qY659Xm3UhavLXCRbM
akTlZOpfQDi1c6JNcG6hPz3NMuGvWoSdQ+3vMYCV08ExYFMzzrZlkQ73O6t2CfOK
hgNjCc9ovBq4OgJFP04RaRj5q3+Av+R2ADUK4LquRbIRZfdMblZ5DEA4n/0AGaL8
0Zpg4uT7aD0ycUgLfv7eGwoxFhBjJnoGg27E5EkUUVsc1XNEvcZuvhMFsL3f/3YG
ZFcFZ88d245m7z4H7OGHwR8tFyYPDtsNQkU4ol00KLwu1Hw52VPrFnUFU97tHiYr
V4W/ViXxWz+ItiNqmevB5R/WcPu1XrVx4EzrsMyFwgKYcoQ6AU9W5JUKZU1uBfTy
j0C4ipyOeuGJ6dIA3pJslNfGdl1OyYF3iZp+1B/kHjQoks8ZAAcrZZTBF80nTxPf
v2skjRwUYZ+aTa32yl28klgQVvhWtCMHZAHDmjxlixcefpND3sC1sZF0oAu9Sswf
qqqeQ/nMdPz49qN43bfm406shI4cjGRfBox3X/ie5f4DwQcMwSl5q5Hn+pouhnRs
hWE074S7Vv6hhLEKSto+MDMXwwHHwYwJe1yM5OfFHCMuPYnqiMNSBqb+p1yzpgqT
DRYqmvQvyHPOrcTICfeubcIWrC6TJHikJieINw4YXZNKRyg/SA70q284TGDqQw8W
6yzYe9SWKMXuywKWFH2Ry0ZgajMK62eR2jvXBbrRRzswgP+72TUFKKXQ9rDmx2Ia
/H61hqCVBJmJXlISHnoBnYspvvUfDuyePFoLFO8V3AZ2zXbd9PBJ759AEe7cTPJE
g39h6V1VSAlzjwA/e10nsWY9F4lwKArBOp1vLhJB/ykX5hVZzoeOzNh1RJm3NWNn
hzZhgtmpVOizsJ7vR4szv5CHs8DJND4ShG1ebJJh36ca7lvXWpLB37Je3kQr734w
/5mISnMEia/hN9ktePVzTshzztWPODMY93h+mVyEC5lwo43G+la2aa9yj4zxorGD
h59nu9vJsdy/v8LGmrdJc1UAirHb3RQmaSKb5FRwRBAADqTnzDR8vNCHC6j6y+fZ
yazlwVaheJ8tU1M1J0DNRxCE7T3ltw6E6yg2uYagKfzqw4S5toOc7xXmy6sRNMe1
6m1UyKm5ttz+TcQBCA9d/4GJJ56fuVlsu/rg2qp/dcveJueEUZLI9oomG2fuODuT
ggccDPpVRSN193cuF3osJqRtxyrOZI+v3ljuqc0/DxXpk9A03KuXEugnpBkGK0ul
qBxJTR/lVMN0+jTdVmyhMQTW5ISqj/fH6016iOS6IRQ3724tQT0oYbpWo2mTmCT0
p/71UIqlJjjBPUupZSkpzDQU57YZD+q7NnFTFIYSpXVNrhS89T2vN4eMRq4C8sX4
72FxiMygCWBZTbQIlohv9DSY89g0vjsPV6ZfQ3SCFIZhNwpcOj6CK4rvUFMrP/Pp
wgT3uCe4EbRV0cA1xFVp80fWT250nIxdkJoqFOqBtKB/7/20HB7xwmqSDSA/txVY
KXkKX4bt+7vZ3CAx5jbDIV5X3ZlyDVLmKWCz7+rPyoH9y8IzIXDVTBc/x4uKqx17
AVqMtvdl8HbOKspMIfu3UdkYJPjJsKkUGmdC8vzAoK2H+8U9g6keiM1gW6Zzz3RA
b2iUoDkpIeyanfy6Fk+Pe9jGrwUHFHCJPsa379LvnBS4hbJo+Z5VaST3jVn/mm/b
3p33O4UuQNTG+pj/OcaYJZVqJR/2BgxH77O6Rsw4ovpGWXRc2iExuKSPuxd9DssD
L8ZlH/fduhucBX70Y9kIuYEUwHEQHOQ9aqmSgEH76VYbEaKSwv5C5nZ8MpoMkUhp
qDfNJcIwFZ3To7t+RbMwRkya1ZCcRhdoF04oeMV0I/bYmw/C/7uLtuqPyA3LcPbp
OHMAzTzlw0GJs3X9TmvdT3HkbYAXAuQSSIJhvHMGgisgzl3kYpKZXxIvG8i4tdUx
kyWElQ3NX70u7fLbk9PpkzxMYMDXZ7fpe2C3dEOlSocUB+1/5z1/LeZ7F8OYswAS
UF4x0zhJJ3sqmoEW5zOEUAz+fzTZmYPVMRqqlGY0JUVxV5EylFPY97QZ6psdQWGn
Cz0HUhlCfeRyFS1QR1vhFxSB1jPkiUuc6+jf4NEzuU378KcLnru2IuSoAkKz2pc7
UZC5NqTaoyjkD0KjJM4PzORqA2rfyXe0bLUTLY+2S912i29rNo97TQjQlQE5fAy7
+B7k0AHO78uUIwkiGflSi3c2tWSBt9S75uLrjhm31KjDOuIAiLBnkFXWDxBKE4bA
4fBw8QUB4hRUZEGZacRf+O/n/8MmlzGbNf+wZfjwjWkOlaeV0+mFzbl5I+ai65ty
vy94poMt1G3cl+5RLDQeAHq1DhmBRN+mBuKhxuRgvRmP9oYFERAG2Y2aSuWYK7TK
neBI4cdSB7N+QmDW9gcFpboklKacNkvIb0M4GY8cT7Mtz/IFthAckwHpMQdGGCLF
rKXBvTUDADWTRbbUxRRbOW2ngiOsjXJO4dyQcal2HvtcYMo5c2uzlvBv9vFCbjKi
mdOommphkqdxoy7LYYSUeUf4VhxSbLdZ+wJ+3DiR/ENzhQAFXHohdM+o0vXDOpbj
SRgc4QRAxsjAD4kTWcEX+NoaTdz8sad29J030yJ38qyHJMa1smsSTdF1zQueQ09R
aE2iMIf77tUOwSq0UNDD6Tg8z0KfNxS/sxtx73GlAvtlNg/Q20amGJu9jhcRFKLV
vCsJ/9Wbnc7iIcEMyg1KQOFi+IP/YvHjyOdHCAMX0tFBKS5UMfcqAd9Zq2b/zOA8
PjkJNQBFBxdOaYAN3ZE0wtVIpnVOWxBtZ0WWn5x/jBVEbe7VwBkD1wwj8HkJwkeY
DX8aqCgI1YWtDrFh6SK/pj/pZ+9jW3i8bqZC3+X1fpswVbM52ep7vSaaNZlP0G2l
aZhE/IJGPQQcPhXCrban7VUBLmZ0wBwJmx8mWjG+PMar0pKbxyXmFng6x/rs/ATX
EGvxmXIjiKHANX8ohhVyIlTRUVdAqCz/ld6xq2q3UiTd8UeRN3Jv/hUiFtKKljL5
Kk81WTOo69AJIk5VnDx/BGTQsHwC1M2lysDYbElOJ1MGpRGtgOROmOMbNvBXj172
1OFXMMs8eeobIT7LUosQNEl9mCxzo2ru5FDb+fiMWou7Dq6ERqJkDzWL0QVmpEvj
rG67zBgDQjGP4ruDLvrTtl9r799prAcBHodC2+E9z23WGEa98gJEcsGluC12TZIB
L9WGuoG50hubGwQuN76b1PkzkN6xSzR65JDmtlwAZw8/fsoMnL2XdTcdPL/fTcF6
5xfBMxMrSqN94ZXOSaAiuMJKjabvc9zsHO1o6nPZwNZy+IW5IqIgjL0jjWoMUUNj
dAO9MNLFtjQoktptlMVzAPHuGGf2hhli5rpESMcYqqzfU3hJ2blPZBrOVuuE/XPJ
XKf7RdlvSYOc4nsQKnZZ8a0rObyGGGaC0pXEZ7PL1YLg1e9geJU4u1AZaoFkJeAi
mzqiu8oRU1E9Z+ilOv2Ej5D1AFrTeQOB9o3/+oeoPhQKezTuMfb78Te1YuHHOLsK
z9GZRxzq3yT954CGEAua22ldCX2agXTvPkX/P23oHD3WAoEpvKDKG4gigzaxG+1B
V3/+GOpRo93Y1mlK7jTkf+Qn1WuSWSnKRxV7PxRbkhoHzlqKaY6SRLJCo2/BD9p3
Lr+MaGTI9h8il3Zt2NQP1vvFz1U+6a8/NYSfd22r0vVauFbw3Rn5F79A5A7F5OJh
zkFv8GSAa52IuPCdR0CeNWS9Ty/m+Y82EgeAQAzyT5/GzUeBKKWw320SGuzDxGFq
0yyVXt9l5h5o+Nj3TebCGyJquYFOKSaJP5J4asmXHGpN4T/fy3Aves9196wBqw2K
JqhymWL7UygrWafOryZ5IfyRa4iJ2lI9DMOP+AjcrZFEQyDfNBSi2jVzzaidaEkS
1n+YKSYA4B4j7UUAptE+4kHtfARb52jNpe+v8IbMA2LSuf7clnqobyk1yVJMsC9a
H9O0tYDpohMO1mkqsuF4f7B70ca/zxgecuzssumYk0FH+nISp0NCCP7e0FgscCHL
oNzfYgTr+FwcXTVDEY2eP9QbDFOLiJVGamgEGbXbRHOBnZ95bc60c9r3eL+Psk/E
N/8hsVUdsRZFuSBm4nQUKPwcOORyGSaPWYmWimnL2Asxs5dsROzGbhTBHKdNFoVM
tG/pInBW16KRENHIxXLuqWUrb1P4KG92gS38VCQ/rAdMQcoCHs/UJsjTYskY+bbO
PrVYi/OD6HEuZo+Fe3M4kTchEEYs0IHfflG2dIyV8kDbkZMx5lyWFvx83cj4ELSZ
0wON42KwjMc3CG6PaFquldVNVffWTtCDz0B2MGpm6NzbjWvgrZZ3VHyk62IV+fqy
l3uRxT7Y0YyAeA2G/rPYLBV+dh9GkGJ3BubSaLrLFKNRWSP3sjcq3EWIlJq2Gaub
oJucyFP1rXhXS/LrEXDrOd9XBC7DT7omAeFuNu+bPgpy7AL9piytqusLs/GN4oEy
leOb0fHF3Oq4lCrflGWx/48g0/ytifg1b1o2GyzIHsAccXBY3iPY3EhKRuKJavW7
NUtBFlf0RX8JaG2YudgkUszq1ytULwaRuvlse96evp+5YahbXLXMJ/F40aa+oC64
WWoERKwi6gtDnP+Qikvxwp7DC53xwm89nOabA0zDUl27tzOOYphLmdhQuKheosp4
AIPBIl9Kws7hqtkPHcBQ50/xg7hA4tldN48XWftasWd6x6OVaHS4yr51WlrGcoaW
5emnbgnpYN8YtZfvpygVSoLc5Ybffy/4eTU9xoga7mjsRM3ZvqxBK8BH/1ynEAZw
MdX/QhqPv8XkwGEayEjb60lzIjBvVsoB71MmKKnEbFYknXCn44c9QcSQfp1G0ETK
A+SISpYlGafu7zPv5Co29gIfH4Kcso8o4jRqrXrWGhLtMmDgvP4zsI+iovMW9Jxw
nVHe+o6uNvzakOk1+V8sHFTXlf3Il6xGIYFdxrynltgHSyjgBno2D4C9y9Vc5EvS
tPVcP9j1+Qq+DNiKW0bpKz2rTb70IhZhs599HftrJmAiFiuna6beveT7j3Y6oOPb
PLRvgFByhsW7tPurn24ccJ1qb0fuh84EkFovFyZkyOm+kfYqi4Hl6AkzGHstDJR0
zn1lyr3Ej2wqbMTYk+a+rDNDadE3qUd5y9H/shG+76qHGn0a2USm/GHUssfOXJUx
cp6vOefeGMFV3awHT9/M/1Vv8Wz9O2FvZnZ0GtB2aqdDOVJ/YILUhaXkyej+C58B
2Nde4aqFcYNNabguyUSJq9FR/5t+Njf0sIcM0bNcqVawfjhABosnN1yISjejw13X
dqU0lyNRVWg5VGrldot+giXa2hKW0jAU/p43AGFAlP6LaV91oRLHvtkW4/h6zDOz
DgM1EKDGOIX0uhKuiigdiRY3bYb7LHm1CDwuwlejZZrFVRyalsSl2ehiFULCDqdN
CFvxdcxq4s1FRxgR8sxwlCkA6SjWcW6CRkDtQ9/Q13G7o0XVky3h3m0B2aFb+7yV
U5ptbkFI1ptGuI/3Hx0kYynEWSH0UW+NSBhxXW/tTeA1CH9R/IcDoSWM/a/IyihQ
xPINNzUsixrizcOjq95hY7cJJkL7eCfaGgLtAnKDPOSOFYf2RkxzQFRQOZ/LVoVV
cFlG17S/NnXzpou4pFGrnq2xdp7Wwfc69ihq0TThKPz9zs99xWA5jray3rOh0DA9
kj8tA/OmpxnTDGWfNct2hq4iZ3nmbWfdxXf6ndhwe8LUuL9m9hLGMuAcX18tCIDP
acOXzt1N6PvqWYquz4cx4X6j5KND/8EsHHlZdc18uEzrXwcGlewHpAQzd1AHwpUh
q1vi+kWqsaSkf3zvJzcPPOIg5RKShPVoMgM7kyZSaJ2ODNuOLh4g+zhXFkXt+HwY
kA3Fm0HAgeolgBwLTN/+wZOCnzEJZdTrHVloq6we8roxKJiO5YLV/tWyltce1wwE
FxdsQiwqxRN0OPOs6arPb6/qJMXDkLjQwCfkbXsywLl5Ebxkp/oKSwFmng+w8YOj
CmizllqXQKritLExJK8j6B5tRgFfVU+PzJdBXA2s8Q5hmkpfK1YEC4d95z5olHqK
ZJyDEMJ/cha2eWuP/NVnbc6e1kzaKwPolqnc1jOvF4mH6ir5XOetOKlh+oiV5v70
AY21UXlEEQKAVTQFt7nR3NJLEdWbduFZNr/TJ8CWnwBmxoN/uJ5ZXQzcY30WlkmV
Lu/5szfeVmH5M4ajoyu9FsM8lR7mcLUZUVfSQmRZd4l34/zHqqJo4icoFRDkRykK
Bb1Va4I7+yGLrHb3dM4xbL1snRS45FkdwEBP0yzGmG/MzlOEviMoyZj8f/1FlHAz
LEQn/7gY3IZSjcFgRDVI5F1AEeopljbsj/Icdv/AyZIaNOkfXy9IivQ6Lqo9dRxx
4X8+z3HrtJZ1YKWdkDj8EiB/z35u17naclZzuhsPEtZx9PY6Xaxh7BfxRmogO+3n
/VNvRLHd2JcnGsDOF0LMO+4rkwjsqQg9wdUbU3wlaIgqW5uJnwkyk5oJ8ClkltTe
jBI2tIqEACjPq9cOk5xTWegyx4k0IiJeHFYDLyOkNheQspNdDCGfuPcIWTjrurqn
VxupgmVvE+SqcrxvnfbikMCAzTQl378bmiK4JN/4B7jhXLSg0KZi/HZs3m7OPSFs
+T7FgMKTmn5MqMSXCz9TOrFXATU0LCkytBkRaD0UlbHbQ/0jR7OkhoIOlJkpOQfy
ZcDZ6lA58Flg/GIvcIaB6Irx5u0mPCWiXUhZ7phAzqqkPU5P95RuQoTeo9fBk4PQ
YeX2RaD4NNmoZMkKJujx4lxWXx5VXlfxHOPojbx5cGuGZ3AiADe9DPOBNYgyPCR/
Fdf22Hi36ULMGU86hGKd8Qw5o0QhcfubAtFtTU92HpQz55Sq7kglO5iRoT0wy0B7
7zX1dd49KrDYP1P8jxI26NjUsBi7dSjaep6HKa1wRoTuDHvTdA9gZkJbvMMg8ly3
qlQujJQ8piPhUfHiZTlA+ob17SX0m+mo8+YjJ4wy1SZjbYZEWTq5Z+qty706k2cP
lko9SZn0/HKhJSnvpZXM+/OR0jpvXui5VvObGd+4sQ37abUnFK9mD+UMYxJvCwct
CwfYgu6CIVPi3q9gqYhu4FlxkOGQBTI85OxWF6PVo6pG4tl1DbSWub26acPVbQuU
o7FsTHTA/vpLEBqJ26mWFgFC8bsdQLt1viokOtcRCD0CwulaZeABmMbpJpvzTrAa
lJ8q2gQZWRsVAd1F0hwF3ZnjYuBvYpPnYkPhjCEODbAPbviIO+X5X8Kvu83FEAjO
dDXTodKDsdD826EUy8PsJ+XD+uQHR6fRl9fMyYpydnemi+CJ+Fbm23tvQWPP4Ipa
fJlJtT8OFEHO5Bx64PVC7rNYDnQHg7dXeZCfolNGEv2MBIwy/Ynotmv497ibu7rM
`protect END_PROTECTED
