`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gK2MnWmqFFr6/O19p9S0ztPgcJH6ZN8OIPXiBu2a/tc5juDOdU1PejLiVWTSKzf/
zuhLhI0pQPLU14ndFfO/c8cPk3cFVcv2PienODUZ0hCrziF5ivn3n6TJtWTCGcMf
g3OSjychv3aHj6GXwob62rWgnnmNSWrH2PQUORohGFNZ6ihFnTCgvTe2k49eLRj5
fg5aSETIewvlP8rpBrXyx3VrnOobyAZLDkq0MvAPgEQRr/58Y97uSp6AyUtqzomW
Dy/BbqZfjuJ7Iudfq+4v6T/k2FmJVDxKMpfpPFMdCqvamJl3KetdwCByB0Nmxmgx
0A8ywE0bcECOBwNc6YLiT13qpsRA3vM9/XfPQqikBokbgBPj0SSPFL5KCWGE/lon
UyL0dtU2fV6BStHCkirCC6fYQ5xU6wY+db0sT1ThmCMJNMZcaoUbGe7+6VaeuWf+
cvphfxzzgLHnOoOrApGxUD8N2t3oPr/XW3O5dk7r14R+yFFvW0mTefOztMfetm0V
nLe6ajSsQIoZFJr+CblIUCLt36XE/blz2RdlbcG5R01gdzxivQ8k7m0/BvLvpkBd
A7s413VvL9cFtTezMBlPmAMjJdooYkb5ZrbuUE3xcmKallCe3H7tSNvVXgZY/V+u
un0N1O2u60UXFt8h8ZoWdsG8Kbt9VM8mPUl9VHdioLKZcIjUeBrW/aD6XVf6DrNO
Utg0Hk/sP4LO5fa7iu1M+Gt6MwtLMdm+aE4vU09lUHp2AH4aGvKNEmnsd8ZFILI1
++LIQM7Vx9VMUU2CFIePR8FMI03L5b/J6rX0Ug69Z4VLOxBU8nKv2I17RFQGIT1A
3WOtg/YrGFFjFrnxpN7+gFWyIk0BBw6oRtAbXJgxZYkDkFYNx4Yr1niMuKiNOBkb
4Z8kJRT6MhnKKh0GOWxx7bRV/YPmw3xqp01UxSyY66t85qp7zd52varvypkWoRYf
8LuvrgR5KPNNh4VtFmy9NL37/o09m1MwWnpp1KZQTTe7yNFYGxpVztJHtynUcDMy
/Gjt+CqnckjNEk2rrqN3/8EG4/MjVx9JNU6HT0X3FNo2OLEeyiNIVuc/zMXjuqnQ
E+eswvH4R/usivA670sMclChVPb6lnIxxi5I+GNt51CEi9Kohcuga/y1PWnLDMPz
KdoNcDOcCWK4h6q7KaSSS/UOg4Z8LpF0fX4OcSnpXFN80vsVbaEkhkUrrBbeUoyo
n6hXsYovGZ3OZ0CUlAqdIz1q7neKUJD9hB+qs/t4XBmqLXCJre9BeBPQMIySaEQj
tp0Ofo7FkKRceO+FTRyt9OuhAeUdDahDcdUXhJNtWQ3lP+Oqp8bec6HIaHrpZV8q
i+HcRt9+9u9MPYNe4MVseLyklgmiABcmG5N1k9BgzCJAq3mc5YPwMLgXDlVVuHXC
/NdyjwsMSPc2Aj20Ah4rKX53sNaRlcjVL6B/eau5dGpQVMldSBo6QApmr/4jUiWz
9/v+VysycwJHZHqmeVcAqUhtOaXp4aUexZKv01Ukk6Fzu5f4D6MC5QE6Vu08Q4hM
2S7OSDrFCO6vE8eVF4+eK4VJhdZSNBy61uJ13BCqegUgRJSJs6FEkGliU4Q0MEuG
V/QiFSrjbCrDW/hhMoELhmi4R7zhwPNQM0a7TnDDJS3HMXuXlTo3aioDlHd2dr6v
Hx9ywMj2hp77z72HsxViMzIfRR32ynrxlNN+5ygVzox1/NkoSZ3mEoy0Y931riBc
Z6YBDGLrI8BkLruyM4mo5BnAKO/zhLe320rDK+7rSM1e6x69qbZHlbx1Zhu/oWNT
CuNvI6KIW81CqgYcj2dViqMEaNakr2fOvljwIM6mHfXfXdSar1IFfaBEA+fJP4+8
FYVoRt5Wf/XE4HFH2Ub99yK8QubS9bOMyueYsLg8EeDkl4vSQi4NgW0f0yHmyptg
HERpMY7I/RDcHjgTubzXok+EwtQV38+5Kxm4wxRnSWwZPUdjj13G4uGgkyXd4rM/
n2N8R8+O9mZHaN36FrwC9ka11a6pBLUmhfCP4ByHkTZWc0At4LI6aKUxLdHs4Q8l
NGiNKzvckpCRi1nHDEDbK1t4jco42KbHp5bX8OitW4Dqgeas+5gN+bkRB1GvRO8/
9toPp+5Zr+piVe9PUsLGfmTLrpQj/zTflbDZ1RSwpACSVIp7G7hllhl+BY8ZoKmr
Oo/J4dYLPkb/BKDGMOTBtTmmBW104PkDZdBDh3t+ifu516aFg8OS1RYNFoEGZ2FF
yzrGqWjAdgO0b+eJqDpZv6ATcdEtGce42iongIqeu5LsRIjmJxjfce3oCrvn2xGV
LK4OKJi7PCBlMhn8M7/xaA6OjertpxVJNyM2fJoHQ+/byKabnFU0NJKdm0sVSwNS
J4lEOnxdfQM/puB/dJ4RfWrmr1Uoff2g+wfmCqfEZ2bOhGbGX2mpAsAaNoHOvK6E
iepA+UIN+eenhv5ML9qG8BOSwEov6DUm+mzGSK8uCulvuD0FYGnBI7uUy6zlBfDD
hXeFnfoPVkduXkIiVn6pTeFRYst9MS/27znlLFu0lW3JAwjnzKZ1qlxLiWV8hqey
EoKRf8ur4Rj+7qK5Pp5YPCl2lbbUaBUbYbBD/m2Bg/HvATsF/oYG3kjgO32xguBw
OUpPWT++iHf1RfWftOQ8sPU4DTz9fipTPIdHaOuC803eH7uDvLTrRYmAqMTryHKK
icI6QyHKKCuxh8z2uaOriSo6YPCQWJlWy2Q40hufbZj9HH+MODgap7d1+BY9zVzk
K8ajDdOo8xGY/m2g5OiMsKIBUXErV422k9U8g3Smtu2gkiisQ9fP3wVgNfrrY+JJ
mZOcdb0KrgD8y6YAvkF+Ah4buRTHTBCWzrLk9ieIIKfXpaL/qkDMzHmuru+u1GmA
+1p0V/2ch2XIB5wTgOfETraLdg/U8h5zvORmxvdmukINNxg5GLPZ5kHn/vHVmzPP
XvD/qXfV1EeWEYFBX4R24GBa1DDTJNsZVcRhP/delUWPeBCLZ+i9ibGeyNu80Rdi
M0kkWrveSSDyXcV/inuFWQPALW0DfBqghzPmnLz7fl+CQr7EbpFwA/Ym9dD28K+F
FXkmHjXlowIEAkZsDfvGy1gdNvEpVWMnoEfQYiYZN4kmYBtr4LlkiWc90QzZB2Jx
GAL9VLZjwVlPbTJ4VMnHDoayVRmV9HrAucP4uuR2sA7CcjLcFxby9j/1YiFNs7xI
H/AhwbLvtkIlSblbnRLmhJ8eQ1X80/sc1ZrX41K2vlkDK5zSCKmPU4LBjtbGlTEU
ZBipaAmhsK6M2LcmujiHSNoSBgQmpadke/47mgNAkTvmRXmHMa7NZgFCfbKkAYoj
kK5GQGdV6X6orVV3CrEbxAAug4Uj05lYuaMk4PAifphn9pBd/K1xUz4CAeMn7Ong
gzprhxjyQ8011RFJvJW1pBXJNkDbgmAX5Z0XSQUcPoAIXYlTZkdFpXDO8pmwYbT0
FF/ZW7Lh96izxV8xMHyCEretlgGb5QkDokRuCEFuX0quVyqtaaiLtDQqZQJOGMS5
Yqpr5StnFuhq5+eGpsTRyIPH7SrdJvKOuMsEs5i1bHw6WtY+N4PHMzdWwFzHJxnQ
H/6bq+VLw+ZhP6mdB9xXcFdo0rerTBWUhliIbO4ba2m2SWQ+B1P0v43ctyFqTUKR
CMgjZD9MsPHaoK8B19EHCyTwKeSYGZCmbgEtWfaMCCiAn0aazZE9lDbmtJVYY0dr
lrKX5QDInQTM74oGBJw+c7JdQmbGSWbKfcUEP4O7tvwJD4SzhrVwITRtZqD9tWnr
8HkzmB1eCkOe8U3vqJvN3DAGgvTfqZPBY8bIJyvUwAKXxutz7MFMQ8DEVj2UG69r
DfF/Wkot9HlRhJvxld5HqfP1c5mHXBkS1vJUv+i05ki3a3nWG0cy4J7aFoTS76LQ
mncHGDlEt7zVnEv6ZT8IskyBvW9gqOgLzq5qpTQHBUNE22xOayHENegn2YXgnZZ6
nixL8xvkVs+nFbOnA3tiw3SSn6QXv+eXsjquiABAWMJX2oe+5umLPMyR+cHSX4NJ
rfMM9JvxCj1LN+AzT8Gz4xZMcjib4v2rTYkkCX94Zkpes38CNzCxrsf7pfAAjx6K
/L4Q9txhjX3hrAGiVVrefWxwQHu2dMhNYR4+vTUvdUcy+Aeskgne7VI70HMKqlzs
lAquUruAQ2/vp5ubtDEmTiKyhrMuPVkX3eU0DRRl1H5w2DPk3kXsowxa0pwrw+2n
Ox0QoSSuGnmFbccmYhz9NJm6f0oapItedVzGnyHxuLAaJ3hKTeDv7zmSN9jhVIEX
UyOO26V7A3WI2x6blLIUIBcCcA5fZDZ1l/OCa5LHqPVpSKqLLK3rv4T61a+QdKIu
bd5EX8TdZbJPNP+A4UDIZ194hid3lFvB992vy6QBSpTET1+HWr00vyTCnTnyisHm
aVcnTX/FolW5/7CXGDIBXBDdeQ/uFJI8JPEHG5fG3kibX3nszhW9SX4At8Mp596r
aj+yvPHXV8y3kl3AWIADLWU5pQcBCyLVPEqoDLOt+7D4YCGsAEbUyJLr9I1mhMh5
+N11c+WyW5brM1+holntPzZrDiwQD/Vkogb75eqEMERn+jye/NPgpecHXP19+/gC
bWN4GtCbAtSoDhPqPadDzw64en7CK6eNlRv0GmjL4A8VKAJA1PDO55R04xFJ+cwG
+gabGy7Jq9oodrtKxPBaAXzRlQtLsICIt8YfosRdeq7DTcGCGcTBRbD+BonEfXn0
7A+DLAHCipzfDQRa5etsAFTIMpVh3CrvUKzjf6P6uByTiugiX++sAUNtvA9Pe1RC
UD4L8iIQk5MG1HAqCM9840fjznKTl2WXWRB/UHvjWOa7Atk/rtP3GiBpgARiBkCH
gxs9Ec3lw5Tupt9ey9SV3NMjq40+3qisJZjNCmVq85V1iiuyq2r3XHujccmRH3qb
eQ+qQTklmXHZp1xNk+pf7kiA0ARkJzEQnzfXeWH43P5aJbB4gPou12X9bim1+WyP
TQKM15LDmvc1diUQ/kAeONOHf5By8aOdP3KK0HGTdSZ/dC6zyS7GVmnOdx+plHrx
c4KLPeBMT6OOv54WSvTgR+nN5wNUmW9A7wp8uq10w6y138/HAXuS2GhP1hzxVIEp
UzamyqYy5/CpMBjzWIKyjTGEyxSRXWSGlV+AvwtIOd+02amgTQdvka8VMPPodaPJ
rVmjU98RxoXE0SJBw66uWyqFKsfXjDe4t3YX3jvgVBNQhxWgpB0dVqlYFvl1bCio
/Zxf0ZIMKAyDR8tulwSWbfjqrZLwwXXqSIl14DsnTiMPU7nJn9ZXUQWQE/3EUZ/u
mti9c7F5A85HDBshRoveF6GR6G5WM72dWGOeG9U+BhrABZ92LhxkEayEBycjWPas
ho8zCfK23xnE1u1uqr6bYuG5Ehf/SOq3YjPdFnK8h4pf0IG9Z+VPJsfxGhwO3a7X
cfYYHlb3jLJhxR5ZCw0X8Qt6Aku2LttbYOgImzw/5ny1PPyOxHSLVrbZwvieXixJ
GRkBaF8Z0HxL2YaqclbVjl7P50+nJeCwrZY5Hj+070sO4xUYjTa+L07ES17lsK9F
1NT6K9ChpaO/3pZcvHRShpQI8r9Q6zF3W+7qQFfJBKOjVH0/G7bZXTuo8j1oV0nI
Ga38PEo/nGGcuSBIFuGbfbispcxw58GC5OTIZeoCLIp0rfwUxCoZORgPJaSdnl1l
goVLHqdb6Prtoikk31Skfvzmt1Mxq+FBucgasZ21e4C+8ZS5zioYQJdyaklWeHi4
ramKlNatGBhUBVWmpYfdtiwd5TEDyJA2oGajCDJ8LBLcVEiGedqU0wImkeVzE/qy
DwqAKI9k+WJnKQJVJ51WVmyq4Ey9YPzhk6Ypn5d48lqb075Rc/3dQFCySlgqIPGM
dkl5cwo5yHoqKcFUt+0aeB1ZR9JD5Osk9VuMqcyn47+Hq5k0Cm1msodOeZmCxdFi
cB4VfOyLJw68uCzHyDLkzGEc/PYQt6ZR9PD3MerRuam3MP0Fn4uEtxIBX2CGKuQV
f/tNI3+n9k1wipesW/9EygmJLLtiY3ogdjMAw3pIh0OOF4jFS8VsPH2C+xEzobo8
fgDgjwe+wMAXwvQlUhK3SKQJlTtokIBOxm35Moei9I0A7NOTbH1HMiqJZ51qcpcJ
9n65uiEYg6X641PpdyVaBLMBlXaGba/YwqhhnBUHcgkUl37B/Bgoz8JRcNrFl/oe
oSZLd8oWOKS8WcBWqRRq3dT532tn2pAC7sxCUe3faUsFghlvIQo4HPx4R9kdWC5o
yzLdazLrgDTdgPLgnBmRU9t1k6/lSgw8f/+t9sfEATlkplVwEPUyxvpgqlNpXnCx
JgxaSW2EsuaaOef1Ea0BylJ81DWbp4hBFTg4CRnmOZvxbqLEyIi19gfh/HvE7tE6
YQ7W05U+bbVRM8IvtM5O5/z1mlhk5wzpbT1v7YMq0I+6VgYmFkpxP9gausVOR6dI
kJZkGvceec5wchoTpcnxlwzvjNP4Lj1idmL5dbI7MotbeztvYsyhIxdnNDjzse24
LYVR1uGVj9hFhVtWqEWKiDudrs0O7OFOb1e7yXdKnHtZWJxQbigIclmP3S7fsYQh
qVy7PngvGuRyWEBDldEbel7jzQDNEa5UgetKGrBfVWlHSZkh3mic+srQ1yZEWcgr
2ebe6Yorbj00vN4ODxOXSPQnWkvVODEcEeTzFMtiOIABouv6gpQw3Fdo6p6yyzJE
agA6GX6XDYKXisER73YDLtt2v/9L825I9G26uC9nobd4yAubfl053ZWUGjXJwbqc
KQff1bqwxJ+0UmeDqHc6QuYptrIJYFkNfHCujgW9PbuaYPPLD/Lm8XdKO5NerbBa
rRKqnYahzaVcc+/TRnYCPsfY2y1e6Hg+w+b/mFeATf1JaMMtCBomV4KQA3Au/vU7
OJ0v9ZssTw1lzrT/81wJc6elzaiMa1mYPW3ezf2Fb8Cco7ybkjnQUoLkI+XxvDEE
4uACPT7dlVpMvFzBs2xi1p7W7Pp42AHasKGshlbDDzfT7znCGTcjw23BWnCjgUmg
2gv2HhrQBl5BeLLXqw2PboOJuzpyAgKFlcWc2igNJzt6XzN1Ktk5Sl4U+Q6olkPV
K0X7OXT4osEQAqIym9YtDIR/7IWnsONmyHjQAgNLOj8BpVmQF4Xd56fdgKFhZVG2
u/te5rjYZcaTxU0/w4eUTGJW8PWVk5qkklOm4VC9Ns5PPiHP2Ji8cSObDCDGlPOB
GDKHqLlOChIFGJnNmuMbzYiWdKNs0mAUv3KeDZ6MjaenxBLFlQtzQeWz2eckZsE4
/E0A1fX3cInp5DfE7x5U3OZmINkvHcrsGDp19T6EIRw19RGDxr1sMrjPY8gJscGc
tCtVCcy69DkaRflkxCl1YLOZG5o7VGLLz9JFAfdk8RxDcsSE+QOpaZbUaAtFSARd
WunBnYQ2jvL/ccOtiNee3DsieEgTAfbuZJ2uMXP8w3I+BUiBX/Ak7J7KADp3crbi
EJhIDOFiyURmlHdCxG63D/f+4eFPgL2FV0LksTC41E5BV1iH/MIP+5MAUGhxb/2D
uwwWJyMy72vC9YHE4dY7YZfBYvA7c7rr9zWSCF7KSYkGAzw3Qd/Jf8zgUj1eEuWO
Zzr0P5qgcx1/Dtpy+mJ/RRDh9cc00A0ilDpxvj482yPN/YxkBSiI87raDInIvTAr
77Lrxe2sV4xuNlw9S9zOj3HAdWX7Cg8dos8COXYvz/Ko9hhR3xHSeukI/8Y7w+PE
McXTRvPla3uiHempubLlmohImXSxNIkaIi/atmnvUlKG445Ki0U139d6coaYy2kb
/cOVCVPFBWcbEM6T6HuPWBbGwmBYnYJIlxEsOhdojOzqrPr6+Vkf6TFQalr62NnZ
uxsTkfhewawjv5SiTcoOGle+JfPX16M/FXAzZLRITUnFEuLaymd59sjKJPPpx3JR
3p3uJ0PnLiGELmuilsHe0SJeQ0voMIDIZSBoJ+IwWUcR1tAlclcL9UIZlkuZ0w/t
ym80K6oFymg8iDtkNUbkKMME3JedqSjhIttWjU7uOE5BUqoIYh3ho4vAo0SUN7hj
QsWvL2tpKs1wUSM1AXDIXnSfKCADhFmuu6FClKWxa7J3eqmBeVJsVdmvYqGG0BKg
Ra5vtqzCRKm3SpzL9MsfNBZzxnsFtthfkcLJDHypUgo5zMOnJoqxJlhS9DjBMx5e
0s0ZCWVSYrREk7DZw5Es3U7vbXc9ROk695eF5fDAMrgo/9HfdZXSg17qocjC883C
2nA8tgZFw0NY+8Y/Vsu1/MiXyzsSYZjUQVbTlnffeHfD9KFWd3RGvVLL3VhWQ7tA
D/bPC/GRGZMVXatf/NNzaIXocPUSCkZw/Kh8M4cSXT9FpO8znxrsy5LsR3u3fhcC
ghYSUgW6b7mYlMY5rhiQR7oqpW6ZQV30+O7EwEQToEIxwIb73oAMMGgun6oY7neS
Gg9hXNN0dTktZEkg+AInYcpMrU2tA+vOYEuWD38Hd3uMM+DwIffaVO0egl4RrcU3
4iPiNnuPoLv8TeRDvK6teniRxdepqQ1kajzn4aqoBq21Xmie5cYAgLazHkgfDWKe
YvgiR6MyRjLAfzyQnJIDV1fUsseP3x3B4Vfqb6e961n5M/XGV2HMgo++fEZmkePd
q371ZjGNktpYB7npWYB3FZ7FRj+1QsfX9/FgLtBRNiFx4OSih7k2GvbD2VRPIytT
GD3gl82nLF0lOipp/P35BaIFHhPo27dn/1o6bPxiTS1ZxsFy8cYByR4euhbNL5lF
QZiOYCo5FQU5n7T8s+F2qqbLy8FG9S99GP+m140gMvOG5uWe97vIgD+sFVBq5pLL
n6yQvPLF8knr6AFjfLBrV46Ln8ZdLGsx7tEvRW80R/F7F1ZD4YIhJukG0cn5lWLH
+hZauQR9sISCGO0o+mRBU14xsnScsmmqelgc+YZOgeKbhgs4/FtZztyr/YPDcsy1
rWThflhprSKBqvyz+KBD4kXb3phYTJSUVQQ7vniICUf7wzg7fnqHHXkExeAtpdto
YUzecVT139UzqCS0WxX6CcIeuxo3dYp5qP1nuOQn+zy/Pp6LlsZTzGp6x96Uxy5F
+9bdAVBcfsiOzpWh0zc0AGwzd4VFHnshdfJhiHwfl2mu+aQ3B0lJU4NyBc3YB8YP
uf2pSDTTgvzLTXRYH2y4HpG25ZxPj4EJlnYL5X3FqPEuaTXJ4a7UN2x19OiEV/Ik
2vXUvjf3fDkmOsAzTDTOO0xQ9xeP7I9s/yKMJiFY92NluTwquOqAft+AJ4zbfep7
kG2bc14gkMpK8BlkDhVXoP5nkt9gT2zrxovAJjHcH6vuH7oMxd5V1I73yi2/ge9p
lGJwhiFwFswn9BBEMHdRa+VifEfLgxU0tR61MVr++88OFCZPh+RswKyEraagPbvu
+JDirVX3G/jn7sZK4xSqw73AoJ4bQui0qZATK8bWTZ6h663Y6JkOCTzIKHj2nYIN
8v522swbHk3J8/exryWv263y45eGHoVEUc3L/6+XCGQ590VDVRffv2DR3vPaU7Ar
xINDYzUnos8UYKcxsT/S0uZKfMKV6vGvcE8gM7ZdnUpgMpnQwCNYPyAvO1PsbgBX
adGztezm4zhBfZbUGOMNfNufwps/69NPz+gbzO5+4RCrwCXrYMgcNFGhmM2yYNvT
Q6XlwRC19dk2l8GXeJIVvi2TGbrVdYqAlEkFNFHNxzK004F7H6BWmlef3CwHname
tDYjc5gDIUebQlZx/bheQwecJfn1AfBosubvXZwyjYllLDjGDbShZfU6JgI8vzKX
NA7a3A/tgiYf+Z0WV4c7NZoGz634ZpBlA/eOpNsclvEUc7vm0vx0bq5qVfcnV8Nt
B0a9V84Ml1/OQLC5De2XbPecQqeqPoiXUWmwBpAlxDlvRq7OhK8POE9nK3k4t+u0
SqbFiTylj45DeqaTMfOvNXaouIvcsjUYGVZMI0le1spCfHgWVw7j6TbZcWyO8FH0
JnN/wpGCpWd6wLubt8uaY7an6Th0AW9BgbEBd2kKVSFrUwjovptIgvlKwovDf0Hw
WyFqhn7eT/bpD0wjV1fRzTz+iBdAq08WeFGrtn259pj+pyAi+975s3ADOi5A9jLS
C/FTeBSWN6anAEBf0qBzJUnF2U8Lq2C5ZAc3zwMrcpXFMb9oIanr2DFN05icn2IU
N7svAGkabjwRGxFWhyW2/tFh4ciz4agSsGO9oQ96uZjqqNyPAF+gB9rUbCdfVUv8
KhRb5DdYJTHbd6Dw7lfBwTF38ev3RZdbNaR+/6g6P9xFPQMkAzvWEDlxIH0JtrKL
AdC5ZUv49jvb0yZ3bGUofi3FkVbGwH446Zx55HFOIgnVQ3nH6Vgfne0ReP+RJ+Ad
k7Uk7MX9wtxE6JR+ah4UxNyL+WXkB1S+IJdL4bAy2BDFK/QKdx5s/u5rVMuAWhP+
6/ZtBEvmgxD/EyIl0di4xHM6cnXuiXq8Be5OhuYYOxEQjG5o8LDVfsiiVnFwbSOC
jvy/sXmC5WgvRGUj+ZZaOkSe03h9gO8OIpC1nK+izTScuLnaBe+gi+SPKbCeVM+o
DM7SzoLaFgBtgfHHs4J7/LqSklPpt/JjxukhoZraDOUhOacZi02dJfJiSBIhVohP
qrThLls66Nn/oBT4B/8QwjH5RWbWiFKYfJ7egGAFnEmPi9Oh8pd+sMnR+VEfFT1w
CrfovtkkeTYwtTwB9X0hkpB7nnLy6VnEwtRZk9UbWnXXzeN6UQkLeUARHfQNWo1L
3u437MG3I+lEZny9JbY+p9Am/qCPqXbz1LW4PjOdfK7i1EfowgdbAX3VKbSdp1PQ
MiChxuhNIaIlOawxt/PNovqBXAZbcsT8zUQIb1PA9RFmbhp5VrBO1lYdwE0EkyrH
xWKCRtHqaSv198TYlEAlDDY1Q/jpmtAyGkqqxcF91EEi8Npu8Ymf9jrp25hWUaWA
nIdYnfiy/iia7R7La8+vHNYQpLn2GchrJ2DW8U83WvT6ELImVbSS1EuJbYJlJTf9
qMTR1ADq2jAtmuaDMPeki1hMuEHBSZ9csiaPhT7pJ7vIpKgy9145aGg9RbzdXNbz
rWso1bN9jhjxdcE20UhMZFb6QkFE+0npu3B/3VQYtwMIsYemNeyexdbhS3j6wslV
dTSE+gpxIKqv+oNRxp4zoYH88LzqoXKv+F2sscQqf8mUAZ6kWNzdoWg5b5nh5o5c
Z4NQ0XwUeCwovdsq9RPgs8AJwEckuujjmb2J1K8kNO3eYcyb3EoejjCvAbd3HW5E
kX6oL8304nbk5b1AE09LOMUojDP4/wNpQ5AmIacAIQqrsLK0A+ZBaFTW2euw86bx
ggn2U/IX71YGlWbMvQwreuftPkbReb46tEkhxCXvWSQoRZrGqzwNwY1GkqsgM6Q3
nUjILM2OdQytolqR+S/8gMWWj61ZhdJPrwgoZNPyrml7P/gfr5aFckcv39S2TlH5
L3DkHF8dhjJUR6ivGn4nkrLUn7hIRmd8IhSRV5uKyuGh3yq1S6HS/sqD6A0ULV/h
4kBROECy2ffrmiwSBR8PIag+oGp+rH0jnGRCi1EK5QcGno2nDIPYQ+PZSPFnMC8d
wvwdL4+6zfTzLjpMNGBgXk5Kt2ak/C1MhQ6Asg1ZrlNx1qm20k7kIceP1xajczOw
We4Bj4cQEFuuB9gvdOlwRHlLO0h+TuXih+oaYu2TyRIemFioq/sEyOFGmgNcL12L
SmTyX+PtkXSgAqgIsvU60urCZndiQYP0y2YfpiWSTVZ0+oDrFKzPynn3na3j5r4k
xwBEpjoU/HU9OTVbpbQ63nUXBKpxABP4NRhRauOy7km+lonGKpHwXLLahA+udc+g
Zqtim6tOXGwcrvB2dH9bfXqfbij6BPxmIgvOMKibcYBZNklCkKF/NmTVaMPJehDt
78LyiDNvikBPQ0IdCpgtrbBGMlLriZ2ioRmC71Q+QnRr6D6aickY/3xTeYH4SZCX
uJCYtAXeBN7OxCYW3Ypzky4QPtGkIOtpUaOechrFyTAKjMwSK2yL9xRwgiWhvoj4
jG1FAurr8whG9bKO1qO55LGtUJHO657h7k2Wx004nDfCWo+ZTMNrSmeLrn2WVmGP
uOSTLGeYnjDQvs9oYPg5BKuTOrSqPSUT1pF4eXOcBFJsdDygPjSPJIRCE79A6CJn
1/8kb7+EdqLG7ITVzdOEZ8li2ev5W2X8J9AXUHssfzXZ+ISRbFSR8KnGbR+IAmKH
gXvygxjYhGFveFjiXlla7r3540rfzcsTRVeB3DcB67/1PszP84WeC3U6tsCzWhlt
3qFRJq6aj63nlUyrn5lsG2J7HflumtyQvZlc083gGyxdtvxbWDnAgep7EujmdwHe
jUNjgCanojdguQrb67Q4PaL5wtilmgGb6hdh/ZLqvpzgqK7ke9jJqn/f/Ho5hL2e
dHfOC9MzOuc7AVnOv931/gvUQrVOzEEKTNKvHz9VJEG4s23G47aujxIhMGPpFOu4
X9eQ7sFwkjV0fVk++9Fl/ET1LcpyfkMuxQKYB6vfuvec2GNsqQEdQySzaLaiDKdL
3HUIpiuwt5bvBLqlAjYcME9+ETsUGz5htimbsjXkuBjP5d6X5OVuMkv3Bwa1nSyQ
Y7xNMtbry+7O3+/PaQpSoEalr3OEIKfRlRoRYR88NhGTX8LHImHPmnsVckK22kvL
CQazx36iOXeoimd4IJ5KUdXQ3aJ39A/YEtzKpkh9VImbwrO7ezf2W5uibyOkzDXr
Bb3sMUO2TQx1baLInMlA41ULXArqb4GcAyYcr/mJgeoPgDY/GbO11OiV8H4RRsl6
frpNQj56Nlmq1nETpLwEUxHbJlxT/K/wFSztUDZ32dX8vvHyXjDEydsdGojf9R09
lKExrdrSN3STuXBWMVUA4mewB9iuJUzr0hOsv4WxSAKgTI9gHOuAX40PWXoh4zD0
jmThmoA87z9sz0YbZN8bnWqmwfFHDNQuasS98wu+p4evuE61ZViBEMcFgv+YJVq2
t22GH8lzCHX7DPofqdM7Ww65Wmsq+t1yICq2youVA9+OhvEJYGEeqG16/jwL2CtH
vo1ZZTV1QVfoX8VZrC/YhAZOfu94k9ouhk2w68/s04GRHcyPSxflFdXLLLo6+KMG
8sJrTizOejNQ6mFPMAfAf8oX1QNIszV4k294kW0fGgiA7dMh8NPl2CLSpJMVX7TM
WO78NtNZeSpbzg5HAQXNMQ0R/lbC4H5VnSD8bXL0cKOHFbVUe2REWyXYjjY2dDgG
0uf1bEBn7oYtsixmRqtvvQ2DNCIBuMxLPWcY3khBxe9ucWpHr5nDwhrdcYU4aqxu
l2R9DhFGVnI4gf2hVRQlPozOLTk+6v/57oss35OeYAqk6YljLaToPPA6BSMipQcU
wodISB3Ps/FHtF8KQLAsIkXdRPVCBZD24mwTZqMjRgrwFGdaVUTvmswQjj1WVNSK
0qm4qcd/6nZMUF/vzSOtCWz3nMFXpzUXCn/X7oIU83Ml6wpe5D3DEZO0fzbkQbBV
G37fpMgtYvslPTMAWYL/+AefU1vY/plAcG42lCW/4kMujbgx8RunE6AF2nkLHX9o
AZQ7q6MJiC5xg12GlQPM5g7tUPHxOXQIHtsD1uo0kYaAEQJu3figiOU0ikqfS8jy
+dmxWQQh401l09oXPmQisWMJ+vPKOHiYGclMgsvhnO4UmTmTbnOVKbqhKl9Q2TeZ
PEUcThlrM2QFGDOPzzMu5C5LdheqWA+4FzCUVEsC0isQcy1lCBYN2Jy127zgrdCB
r6P1HKuTO7CE6xtgG6gxFirleIG9pAiqqKAJ8bwuQsQ6vMDHgF8RF0Ta7m1fJwxp
H/6F5riPQA1wHkprGFpYkwVLxA/QsXtoPbXrtYUgi+hP4zMv/68TTrw9+8hO7b+H
Y8jSIEmdC46vZl5LOi1lcShjw9hI9/gXIUghyKr3xyYfuRB4ptI30Ln5nGeDDZ7l
GxBP41rUFjsXc7yCjm3ugSdgZuitMCa1nG/GeYFkWAbKl+EMKCNZmnUqYGW3HdAJ
3UNjnQVXFyn44qPhLKjEWlOBIPdoScRIKa/vYtMfzES9kyRyOmGOjbQx1Nq6u6Vw
I1g37fNDdJ+u+AKHDKVD9kEMKpSLqidAJgRBVmXA60ErPH6rtWcuMlmWmD9seYvP
dl4igLcRbNDtt5csTuFEo0AIpaRE7qfWyE/8cIzGM3eBk31DLGvkFGxrCwI9/wiI
NYA8R2hQ1nemTRtWQJ8cstYQP3DoXpAJGKlrznWP5Hf5by7FQR+dBDHWu9iZBvEp
GxPscJ21/kPCc3kt9mtUgdma4g626SqxFs/3/0aBw4NgbcLJ5nd62q+3lGWrj/C2
FUi0SCc6IiXDsI7+DpI3NB73/tGBQLkO6UHCKXmmMNPDRY5guWV8DLM3X8aIFHxO
SBS/OuxlCPxKtR+hhkI+m1RtodG2lzA6mOIuS+LZo7JnIo+C63P89o1MQ3KwnNgf
NaGTNTsKr5z/kOk7686mVuhK2im35u570SGZ2CZyu1LyGth2MdIKVzBkUrgspe/O
HjUJMhVznkDBFe40VzvN0/Vhmrr/oSQDpN2cuvTFT5gr+tACj3oNsGc9GZg6Rube
Nw8dYRY7J7b0hnNf7ev/AXE7B3hvoHj2WBhlhoijjQAtQc8hT629u8na9QTfoj5z
XpI08xTO1m6xSYfUdmXfVZDIFJT38qp0SBiaFQ/OqpaVS012967y+1Hmi14+y2J3
/AQj4aw1D4kCi9vVfuVNtNGFjr87X9AfXCRFabDhHOCu7xpdFQdjtRvoAlbN1yxf
XNhODQzdZK3XZMvMgpey+H9vqEW7iPAnIzXV2SgSQdEusGn3iMsJ69HIQ/QGc7OG
vcy3+lIEqOb71+LWK62ibCoUsT9HKPFnaygmPzmQ9SOxkZVwP6uwLFSqOaISRsMU
ajQWt6NRP5ifLjKZA2zMfs3iOVwMhgH/6hmp0e97MQeXpIvJUbTc9hIPbBe8HU6F
tMvXX6/SV2k8f/Wcq1Sct8JKm7/ZjwYjbGqYWK3wXm8iwB0NxVsH3JqFacKVE6lD
xWqn8pJ1eB5HLPd6hVerx4vObjEyap0huiDOmfoR/H/2ILg17SZmeCEsWQVg9Pvo
CAx9PNlIRar2lsMDXyO1u7or7s1wAykUtHm3QYI3/WP/m5MutWKnWzSDSRuealx0
O1b0jajizTwrmatHfHYRt30I+AhvuHX+1/PPAgBmPRVBKWrN+3Goy0/KHEXRmE4S
ySrYLQajRRDvkja85IR5+6qv016X6Rw15MxcnbRHOqs9pgxmIOnN9u55jGk3FxbR
Zo2YOaemqlvhGxLKJKSRFDgf2H0+xOYcpKFAm9JR2tT4C91OZba3Is/HQB1DTP4b
tSf9ygpFVBReG/V872ozBPZwzkYPCbt97z/20mkxMkrpN+GMQ/rPGI3q+yAQkc2m
c2PxtR4Nvqbk2pXEXcJg6/MEhyB8MtG5kUACyWMatWuh++5CoH5/IOKe6mSbBoVZ
An6QTf9hbbYseedWMPoaXIeDOi9KA2qK2tY4pbZMKYxTYeUwMpnW3ybhmppfQTgM
zk43YYNcfgW/g0s01vZU4L+14OSVRlVeD7yrh//rdsPKK55kFNAu5DBIEXw465Ug
bWkxEdybDHZq0+hdSpqZi3Dukb+u8sUEFfHr5QnI6O3sgQgJkD2xdoUNK9wYi1N/
WxxW3LM21abms7fowigE7o1VXHkSH+Xd5D2/WrVlsnJh2R3Bj3vAWY883gyaUXkH
FxJC8UjfPK5sICUK4BYBYf629HJ38qi8g3w7WzkjXQKRuvRAdFFLF1+ni5bqvVXG
fcuUwgI10BCUJBkvBw32uOsQM3LiqmjJVcxj3113LYaA3HivM8VedUVvVPRnXSPx
Trg5AvfqaPOk9RxBylPYpXmcf8G1Wznl6FZqpQEKaOfpcl8zOV37Scz0Q3plsiVF
YFLB/IUWJEkRIC31dRksp3ZidPO0cRW8BunAEE1PDrGn7e1Yr7UAKiIyWmdUlriz
Db6dajzja9JRqGhzE2nwXZkgHYLj8XZyKXygvw95uewwrd9dBzRMHKcyhRWCMC6H
0u0cBYmjaAEZkQ5UQrkCrP6glztYiIXjVOm+TmyaT5HYSCfUceKc6GWUjVQIOw99
498F8wjPNGILH1ClRIL8CIwsvt44jKWULvKpo2y+VPVI6GGgVMfIVd7q4TkR69pb
/LUK+h6TwKmY15OEa+3LnQA81xCgHq5u4++Js28fKePbhYfUXTpE8LE+3VhrZT7a
wLdJ4dmRfTmpsv4lyaDRa5g/sgZ6ko6t57Dr0YHdqu8lGykk1PmOddwqcrBDJTct
TjKZ5qnWQqZljmE30lytblj3gyXEfzDK8vkSJA7dyb5TWmae7SpCJcyJoJv8/SKo
wyPEIFfFfDm+vOn6d7BTxwTbe8zs058RGS+gu6dU7RLXYPC+bxez+7DteLMDVDpt
XYojCy/L48+Z0Mlyf0GgQYUiTQpUOHi0gHrpPbYsCIAUffWBRZj9HaiQkCcD5GMo
nC2ZQg0p8mUL+O2+AwJyi7SMq7SWwvNzTk7wMoI24eWm2tH24CPxKSd91HNwru1j
qXDi5aKnckuNqeX8o8xVZE1hbcEN/CmeiAR8xBwcGPH18Iqgu34z52cNXFmsUWfW
3bwXYE26do/OQS7hjzxpYk8ZwLY2W48Ecot3TXFhQpnxrb9XjBj1hsm/OnNhLahj
ynKSz4OHDUKH4yTtXvzecIeljAdhXkZnqC4Adh9zTbIZ5Ttrnv1C1fgezrvfZbIW
vcLCIdAhX2i+ooJVCmzvuqqDQcxsUIyqd2Oym5vAeterNqKZQv7ECMWXS+vsg7aK
LFT5z58tCZiHrwUijRepjetQ5dJqxnYSoroibrWtXuUucJPgfIW1vAqmnJCj8CSq
Chmgx6aaelMItebs3TNihlxf4esFtCMCixrW0ee6+GCHubHnYjf89QXvmhjS+a7a
8M+kyaTxJs/H9owl/vfvHqYCa56xv1tdEGppIoVb4TUVNJMwKSzB80tiK7FWjLDC
isvOZP7Bf4ALzk1wYW5O+WXwlOYUMDGEFbslt5cUFwTT+KzB3Zus2DC+VszaR6B/
LVqZ7FH/be8fsOyOKf8icWHs9CZJoMHDSj02gF0TYf/DhZIcpHrib8iGu8oiQq+S
i4T4OVXtGcGU6Lj4fbOxyVB8Sro3KibK8psonoFMMUJCgFaSg/nSS1f6MCPXlJ0I
RhoHgkpEOgmcBUc9wQmRELo59j7rJXDqgiiX4S5ud3WkaOdlG1spg74NfMiTdM78
Kgyr9xU5V+0Hv0Ypl5yQXLwn5XSd/BWK+dsE+BrCqoR1GaY0kh5Xu5MH/TdYfspT
ZfRl7wN8dMk96tFX9JLI25Psi0PjXwY9xypUZPnYmj+xp7lc/ZVIt+5ee0yXD6JS
+aCelBuaXfkswV4NLoLmPBO5ILSKCz1tTR70s6f4VA2+BCHNbBF4iFJmKd/yXnye
X1c/ZkAT62EhDe7s4sKE/LZrp4XTPke8T3XyFU+0FPFE1VFCZbWSfGC+4+BwCOH2
0Up02agS9OCBxOVo8OtToP2uUxtFkvGHw5o3q+h7CD0fTq+3qhqCx7hPm03Ll7kv
vb7sar2ob8Vp3NAy7nTmxLDMvAu5+KB19qzXnbOkM7t9T/adTXpuCMMt8HJxni5x
rnCbytXUyKdYk838DO2L/6BY49kPCCiAh+bF0b0qb1AtVKSuJ17MarIZOMq3LT5A
HCRxWDBDWieDezM5+ZdcV+OBXNOqABRVW2YKWk+QEU9zcxmK0R29MVynZF/6RzV7
aad93m3ETQA+fs7Kx+xFQxJ0BB1MGLaQ85EJO8ZI9Tcx64l1n5s1xiCyBHe6MT8B
AjQsNsUEJnREryqh/v6W/3A30F+zLymPHOKN+deyypmm27V+RR724s3eJzw30DXz
wCMaoeuICmAfZ/W7fCpjqjfjk+SPuNi9VBlv+S8g9JaDU/QFOOMGm6mIZ2qMow5U
4zkT3BhngCAgatrB7MYLOsEYLQIzmKDqJM6hgjMGVFELuMX8n3ZibryyTLUMUG+e
36RtACLWCu6iorsi2GBDryBkDLJGUol6vAaRL2Rc/gOobcd6oC/t/yXnoW2T03Md
bzqWwYN/TrxHUIV/EtyASpuUgLwfRgU6T7dqtO8dGHRG2lrNlzfAAUaoplE3Vto/
decY2ahxjxzkRNprC3Z+yEayD5Qg/wrGXR/93d2EM1FDkEr7JyD7OcBqktb3yYSd
YAPAI7PWUbBsZhHdlDB1xoqLFl8AHlLFFvgZN8bRK+G4NBGoyUJQRYQkGscjZic7
0Ra/9wW4Nm8rfCRYKsanVojQlPvx+XQb0l21OCqMM6TVPR40Llph2n+AfFpPyz4B
nG/JDsG0FuKRS4e+NtLvzS2qy8qy04hr34nHftYMzMLSqcaI/JghwGz5eMkYnFna
Youj+Pf+IJns61BPBXCsOlTeeTprmjFmhxiI4pbDzAehtTOND2Ao9zDtNQ3TfCwo
in22IOhnaGhiHgF0GdIoPCl6EJvnJD8emVysJm7x7hRbFTXQNVkKllGnhpbaTBX+
MQuZmhp393pSgJZFxCvMC7cQeWT2uu/EzLDB5RL8erdp5kFX1rSep7ltPtkX++wN
FX8dBZ8PpfyxlBa/X3+Hku/xgWpOkZD56oeyUhH7uFaedyRtiGsZPQr+d8+uDnAN
kki0y13A2Hw/t/Oir8fRMAxw7o+gkh6jYMVsjg+WswmaPnPUUe6U8X0f2/oeqX2F
Cd6Rssg8xQ3JF/i7sJEONCVySOPKo4JK/KTJlYFsTt0AzCZZfhIg84EVnwxpAZEh
oOkLXe+e0hkPjtKk+bZQbBfGk1KOKa3/FGABOAykw76hQQE8M4H3ztNOq9EG2UE/
FaLAshLaHEsshev8+9fCmfcYXg34XIF16lHJGMl9Wu5CJh9hKYleEuEb5WbYSdj0
iKIXgKOOuo91AaZXapxZoxaxF07/FURdNHcNFCzfJgmKTxmgSvJ1VQ/BTRnV2MDx
ZSOAkCVg1iakQmtV4tfv+/yUberavPU0P9TlzEAlTmruSHcQXEdt0Flz6scYMYZu
bC1e7t9/dbugysxiBWupc474ySof2oy+nEIZGPVg7mmNzFHV090lohfNfkwExg5S
Y7HTMR0btHYPDrogPHfSVjExJ7Bp3gvWRh4JtF4/22jgz7eFG2c/RtNjceBdVsFo
vh0QngsU8yoHobimr4wlY88Od+d/Fm4rRNiIl3H/Rjm6traZaBe6vhBhGAafqDvJ
PuE5AijJS8qFRiBZcl0mwi0GJGDkEuN1G+Racm/xzAuUWvNV+pT6+omzAKeGJVbo
IUKWwJLE+KaXF+iidvVA2JFlO1yyYNFRIMA5I993lvEZs8KlNVQf1JZsL900slMZ
fipgjo/tfCTJeAExuuK+7h5IVqZAPCyosDZBnuMWEcfm7bibq1S1yPj3691R4eAM
311HPBGYVCB5aedP+jO8ANNo/Rnm4STfqcqDny2io30GyqHhZWeH7wMpam/CccGq
+Wu2+M33bhoLV0Z4nq0qRnM630zZRMLIuWT3oTo9cXSa7jUH94rt/sdp2uPf6aSB
JXcDG8YfEZitgT2nD6Umj5JDyxhhYX8+VwiVTZn7P6BcnMQRPf0/6OosYJqT3e6p
6+pr0zkvgwsEMCBeZc11G+wnfAbMWGDQLYMNTyqg9NtGE2GGQ0FUR2DU+6GDhMIW
Fib+uw4+FZgk2ve0bsOWMeR5o4zUGXFHSp0U0L/Vqp9+n4oNgQmG4xeHTkm7M1Pu
I1a+H//yWTtzzTW/62vzQlpEZCUGOsbcelA8gsWRjqIrKfLjegvhcaMr5QxU7w/Y
aaSQSRkFkirBCZEjXSvXXAggAoPbnfz1JeXwiLQcY2PNQKAR7OncSqxM5p6FzTSd
hU2vHvZIAB2IMTxrGUH5uCKU1qq4ptLtyhywYpcRB7Il+gIdIS/m39rG9ypQt9eY
FFxtAvtsw3nOHBUHyS8ZnKN1qx47Y+xQqmLZPm3kLkSGbQ5vQgd/E9fl/zVmrAAy
LnkkV0sawmGCgeOS0+OLBLOqLhc4HQXsFg/GQaff7ZUHFYTAgGWIQ4JtAzB4hpjA
1UIOZVTDJw5bSiAc4ZsLxI1XUbEvijM3xKhuDNUFqc8MakWDJX5onYCp5CuynQPc
DUmnw70Z77lIIQV8btQ5HauSdnyM/rWw26ygpnEhZhjJogiBSYWGDK0cTDe9O2yp
1OVzIO0ZfluJ+BqgxTMlKslXOgko5jPd6StEbOLQnZ0/l8X0mXUe7IBea+mJ77MZ
ttVgw91wMoNB0GCj/o+0p/VHnYVFSv6u20zaDI/DBmLcA1DmqNAp76+WfW4uEAmR
d/F/jtC1o/tco0NsSX0hYzYg2Bfrgw66TGmxADyayTUwN6gC3IJUs7TOaHPqL22F
vCHAEnAxeoU8zDXYU5ZOH/7/e6HVZDPVl/DupfZtzfVlPmowOH5POK06M6iJjmBF
LUxF7DKyJgG52tA3L4hkAJ0vaT98CRK8BjSpjAXZH7gAkrKQS5asrZbwgGBaQo7/
ku/NSSvgc60NWipCYyzLvQKcy8sy3B9tjyXtJcFeL5CkjBlh1yPibSgvVDtgN0df
XY2TIDbkVM5Qu8FsglRVhfWEBmkHEzPfxBSpeNxltA6eEBDUMoDGi0u9t7o5XQ0l
JoanksJFYL2vXa+Ss32bbR+Asna1QGY+jLwG29sIxuJhaoUAUizbLBv3HB//IE9+
lqeCq8+8LbGUJxxAv0Zsfajf2c0HvNurfIQPTwrTegWSl9Kvf8n3BzOZAIIVyo/7
jp1KAx6Vf7oKJEXfwxK5RAUL0Gn8Sz1iX/4chUGfVqE2+nMOgX5P8DG++hnRFv7T
ROaUMXJekFI38w5pVoyu1IbVMwgE9P/QZQCbk4kxqI4pALxn6b94Yt8NLNvI9wgn
45Q5O+aRQ2nyoTg6v503mEdFJfYoCF5LlmE4LwFCsqnKLGTs70PKk7VmVIzU3D/t
gA30mXAH2lC4LpPgqFzCz+cFJis+Tt56Rd02H7jlry0rGe6kdTu4RTPIYz/7VyG0
cqwnDXDnj2z88kUHV59kZsF1DSaFg8HE7rs7uj+UBQ4=
`protect END_PROTECTED
