`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Rc1G1GVwHkpFXKKbH5Cu1avxUoBdjQkQj4wQueYLi2bhlUsesAuwg0fupURh3TWk
MfuDJgRX2hlGfV9tsHRcf97NUAgTTR8dXd7MeISE+Y8f0dBjj52TMIXuYKjq6Fk1
lsH/6Rok2hO+FeXzPuShGfVVkfPUlctFLQzzLShhXr1ErHujsQT0EGniZ+zGn6co
SDJFTZy2JpjdtsJtAX8Lr3oSaYQMRDZ7eWZXHyQkuLOxC/kklG9McXTygj8jKb0E
QkwjI7ULwDv8wJN3i27QYdJeeyPl5JPyieSGq4PDSeoVnrctbPew4RelILFtNFdR
+4HnWMs4g23MOB5CuD0a10VP9LLKemkA4Vh69i3mlMIleHodQhE0EGWtZxi+yizj
y02CeMcA8dxEaKqJ9eiC9kvIruv8BHNE+yF2GMEbNUE=
`protect END_PROTECTED
