`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiKh3XyX4lxl+G86U38ls5wYum9iiN5puxMxB5CrDAu8NdJXn4TmJdgKLvc878ka
JiLIgMPJ3rL24syk9Pz5uJ6AAnKiNqCjcz3oMncDVcD5wq4ffIG6v1mOCo2fG+eG
uH7Hv2/vvN71ypCrc2rQeYVhk9FKuNWFFn/9cVZ2tJ9kMlsxYr/ybMe4BtivXxHs
SUroycr7Kdk1pJWVVO3ajFwHcA1rbaxIOMzkb3QsLWFv34G/w6ad5bxCc127gaP6
vypoQcYYH5kWRlxF79kwJ8nP/Vqs6XKY+Dvm3iIYWSuhzuCvzUZ9HIiKWayYt4le
kAlIEqc4WTSBBWTalfWyglHoice3ViL31BOI0Wz7q+IV4reRxlHT6n48izodgWAF
+mZ6uDFhKQ55ozmx/kcOi9nY+nUXTP25XfZ7EwevkwIu8izTWhy18ZkXojVlmPCN
kgyLZY4D3vFZphwUqg75EubKPAFMFm7AfK3thBGkpVs=
`protect END_PROTECTED
