`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c/RYVjydUefdn21C5knocjnQiL0CqZZivjFfT9tSvCvMN0VEcdc0DSn/CfZQzv0G
ZICNroX1zFvRgH9QxoffPQ1XJQetw32VGxN2xDaCwO73XbxXYz6YHkut+9XRq40J
emiSN6O8m8bzEDmiwNXc0oaqlZ2RkxC+uKiMQqM84rXSCnnxbU902PrPHD2zOHCz
CqH6Vx50GWdHWHemZ9VrbTzFr7JyNHeojCYTdiQ3ZIbv/MR78jW3WRPlTJwZeyq5
ogYMBs9IvI3OTSOrop/m53HlMQsOh0+hXi7uLvpLRL3va4Kiuiqa9+BASpOw1awp
Zr1uCE8oIBx45F85jd1BFt/pouGvduVhjO040/usrmOtuzUb7S3Zbb3pTrasCRMU
JaAE5QMFJy4j+SXiuTOZYXsLIA0HjKn7BRjSap6nO1qy+znH21BtdkwntZ9l7OFm
eQO/g2sT3iH830MijJSQeY54e4dZUZXjrWROsJjzCy/lxtdTsJMZXgUWsjlPUmWm
RK1SwfPpr2QSYk/5qAB6xrDtb6xPDkLlAV8xIbYflwBNdy7Wev/shVmo0a+s6wcD
qlyypk09vQ30kk8JrHDkGlugyDkRFTD5sNlb6X7WiIcV/Z1WxaJBoXVd28MyJeQ6
BlU52rYB+a/jUMc1w7coWMxZfEq554QFBqGHdTjVKxCY5FWCFjXT8Al5tkyNP/Xf
sk0C59ZSPkr+G47VAuNdpqdBZrbFlA3VSBmv5KjH9VKE42gfl1AiPJwQPLqLsLG6
wNnfKNbo4nBBolmVLfCnfbiIV303wpCLn0jCQb+9p3MqUH2J4Wn3C4nb3KxG3IvU
rqMNACe7VUyy0YWcEre9uE+ygo0iwljh9AKDL8R71ybKDc+BvunMx+XgLB2GNT9Y
F0TJuiYSRE1+goi037V/LlFnfTPyhuLto6nSj0klIJespzzOlVv7rHWxBofynFzR
smlOqK8/kMrsZOBujetGmOOkVjJsUwhhrGdipWq1fzqrCLhjYau5mOD7hH4uke7O
aL84TL2VJlmwu5rXsYM7Fev3vlK38JLv8pCanpkk+8AfAMoy63CD867dlA/C76Fq
CbBYDkDcJPB3Tn3lUhn5XSrg49W2ztFmW2Yg1vSK3Wh969y1dw6WFoUcVKq/L6Hh
QgDeROACNqyGeY35Zy5u0NXbKEdb8aIHksD7sjg5leQq/Nh6TK5cvPo5WUjTI7n/
eq3iD6mqQ9XOvP788aPpi/yyablM3uTpWBSyGLnoFYZX0zROcDaJDzKcmcWa0pSX
fnVJ8hYKb5u6slYSRjnXmscHKs3gcuoZPnoO7YTiUpeGqQAzh7p/1cxDJcWFa2ng
EO0sn0HyLjWIzs8W7BlHxLLMZPnXhOuPPZYhniMmR8Vw6ylp+KbbqwY1gGoR9OgX
O/UwIpNr4lyOlwytcoDvP1EHTzIqyZQHhe6uVLqLedP47XzUDVJ4JgxliXkzd3GV
JXRqtt5DpAXWZOhsJXDbBMIN9GlPYwjoSlm3OZfe3KGa2jXp0uP7G0NMGhtDDGwo
cul/4FgWf6msw54X80g1eBpylammwMMiR6iKVgU3AfzSiAUaia31mOa6hvCGLYff
8vKQCRfzXBe/9cib8lbAbA6LPVexQSzs2bLm05uBvvDgrebSr4MiHXBMH/exJQJI
HJ7NvEAYrXp0fZtH/QaI1h8rCH97/o9Gayj7BLArfnCQJFIj/cp9+xxcIHuYTT/U
iw+ykazc8JTe9UfCW2CruvrYoP5KKtj6jbvi3rG6tAsyTnjImJ7YbqmSfS7lWj2R
13mzAE5aIHPwq2qUigflj8Vhqw2q3EALT88VHvw4yNHaIliHGkYh84Z+YiaGCsnE
BJUxD4lxhJf8pKZ3N+myXT7g9w6E13I4lpPZB2dY2mVV/bRvEoFlJ6xhgUV6lqo4
Lm8Sig5oHx01QRh1ozRTB+mOfhTx1I55L2CjPj7feH5AWRdoNUxsXZ1JP60hvZEf
Mdy/u+0EU7yI7/Z5GuzHIIEBCSSRSIyWt2NXDUOa5sbeNyXAlqeoP0BrfOjmEqcT
4+Eb4W57v/a3anCycLB3CCDWqydyXIdb4tXGR0wjD6K+vkbIPoBjFQAXlzhksxS+
EwrdrX4Whcolb8MzI00LAi45ZX4AtixmLBLwD17eOVuoNO6JHEAiQ7bhvry6fG0T
qyHhtqdwEhP5X469NL63Fct+g7YqVnd9ktaWlyJmARGr/NbEPhkZqe+H8mmtxozf
KeOCDGLvuI1ebcDQ1ta0+IiYlldMJGQIlz8KTush/fzyCfnEOGpbLW+aj4zXF1XC
Ok/KO9iJdx93bNsZNiQMm7ddzC0xlhFcSdaTxgLV+6TOZ1mUS5QJgwqq3LemESGF
PQF9q4FcRxQEr8dx0YcqCYusvCwnBSx835k+zVdtwdOedilch4TPzxNRM6xoru8T
ol3SLR8DekxH3kGf1QYmUCiNyzt76OrI2U0SKtKJ/P+MtpzspZ83QnTBThjp6zkJ
6h9Uxi8U1JHlPWCEXi/0JoCVFET8ZtigmPD5ebqz70gloccOBTfMl9XYr2yXcMTH
QJa/aaiOteCGHWvI1MZUdBYWEC5i3F33COEm+pZV04NDZip8hbD953/1sXOrLc6y
7qdgOsnZHzJ4LQcz7UCk6FYnRk5B5sjxoqI7TPza+AjFsU1LGBTUNWa8lxd/MQSH
PMkJzz/UvPc2AgFoaokNJS9JxCSRd7G16H4pEjfJ6WZobnkuARc82UEqz8VeRDzQ
lNgNXbTjaTvSuWsf+3+zPDi0bwE7ArXrBUQ04PVl28QqybUv7PuqP3smPWD5dUJx
nvWH1y3djXUapyVeEv02qBLwk/kvuBjMHOLUD4Dcb36ZbZuckMHHKY1u7tmtZSWy
FAzJuwh7R8vqUheNQnCLg+7VY2bCIoeqHUNcKRHAWTwJp05eZy6AwxVW3ThyW7oD
2lXpeYpXP2/vpjK9Y2+foO4/capZH2ZzUFCVeuTdX1tXLUhtkX1y0IEPwQSzKaa8
EFkgSbbzJvcFhw8pzaukTP+RGgk1ZRlTMUBh4wlT73c/Zi8MaKp/cvRt3f9z9U/w
mwL0Smq7IbeTyYK7Ilp+w/dYT2QYFe7CxtcI0TMuWl9qu84GorPkXfByhL25ZzEM
4vWI7R1UJLESrSViER/BWH5GePIEtY+uDk86T6NDA/2Jv+mP7wOXLNoADX12d3RW
FgoowN+T1lA4OOAErJ4w90SSjL8bUgRavRf1/gYvKMkDaakaDiQ+uz1pCEWBSfAS
vZOxpQaH02Kpq4Aa5Mcw/7u4OMfyQoQ70cObf+so+ifkNU6R2auQuEFnye5Zn0NE
VVe3V/pPnlZDmTlWH7CBhIkN7tbdD/lrqErVK9Y4wDtMz5iCVOeYG7w6NmElqAcr
FMsmOTpq2RYx68EpFwrJqBhCUVb2QIgIN+PO3R1nrtbIt8FQ6NhJepgq5SmZjYyO
byOz0slOM/NoAEfcTi9VSXMMcFbyeS9uYOwuaFoXLH0o1qLmscZJ64TTqe3/y5ZL
lH9kMGjQg3VzkKIjZKpnNqRU0XroqMMabn7edt/tifYxnqB4aG8skfA+/WJFcSNe
US0G+BCpZbxy0dUBZf+e1HDf6rQyCKz7ooXEiZ1qejyAYoQxxH/rQAn6WwnX+e3R
XLobO80U7XZXnPPuuolvdWlgfU+Ohxr2mE7AljPnJAHbUAYPhQsZcGOdRzGZU0gC
KLKR37oYGwwB359j1cJczP4fgSRBQAcQE8aTolG8g+Rcy6dJtcO2l5vi1NMTV577
uZdUubVICpIvolOaGZBT5BIoptgS2VSjeb/YqLF+xG8lxnUyeH89Tt0nMGr/FawQ
WAC6leOrH9BTo1OirA3Yw9vDRkQIIE5JqAInsQ/leDu1Trx4F91A9JE3cZMUfXRZ
BKQ1FfnHz2Zq7jQxwaCsp8SSPlt4mRBvpOxUSnUDXCzOFK81xSPO6XVp1DlcdCJ4
GXMT2aBvjzi1/ajviUYp6VnrFk91jCx2u9IEkSFJi7niPGcnAIEUS0dycy01l/RP
pRUXvsTJ12Fr+A39YDfVSQcm0h+n39hqp4zFoWxyI3p8zh3F5jdDRpEefu8pP8Es
Qee40IDof5tYerlEG2h3e5EJ3wV/qDg6oiQtRu2MwYDvh0JmAWuEAY7dyCh7qMGz
Afl2hj7pPmSlGipJRPyI43Ge1G9Y3gCmc8wEp2RD6PLJ7YrNahpsdUKkjoz78Vny
K8TY65Uj5D1kSD8jKgAIDHS22lmcWE66k0z1yTNeYdspKR/Tol+XjetSoAhVfWql
pFaOUjb6tIkg/NuIMB0w8FBOb7WFF7CPf+227XVXCo/al+WCEryf2/Y/TYarQgMh
wSvHmJdbP3xo9F9BrYiFndxvpC1L8nSKJb5+FwmIZPLAk38dv0JQg/cms1BC582n
RWwoaLJFW6By+bmCymO363o7/cXu758K1Y1BHe7yogYyYauo53dYjg7tNqfc/sCm
wmTciYCmAwuGCgE3uQgq2AOETP8nH8RAKKQTAb6yrDKrFyXG/FsxErPeUIwE+ySw
Tc5JnxC0wsShk/KDF1dBk4IooxEnYM0/xvJ4d9Et6GOQMlBVczZtmm0CAaCmz3aM
WF53W6Ei0TIN6IESTQnFkLGBPkd3w8Qx2XmJ70oFSEIi+5ixjemL6ugL0CONFguF
x1CWUxwUrkSNB8lK9q6KoufrZb2ouiLG4F7cYpsDVNI9T0crPcz6sjZnrwPnzs6W
Rr1YwMInSuozQpGdJYj6sq9hDClv1j1qqUdJQIFvUO+6kqzZHgCE0dL49G8K2Qj8
/65NR2ZeSFzMxIFI1ukAIGTEH24kfcrKTZzdagVrpH43c0iMb6Rts3+fzRbP1e1q
PzESjMbm1r92KhqUXJpT877Ri3DbQReBI05x26JkTc4L+lWGkZcPVl5H5V0g3jBu
jZp8UvDjw9Hi0M5+1Fv9QP6nTavo4aqbIdeRmTDpKp2DrIyKL+xqjgAgFncTETSR
weFwBdZeoOJvqR0FwQiOUAaYLZNu9Ea+utossPWxU83K3V5j42OZpGQFLvuMJSmD
pEK0EJY7+T33UIIhVknR10U/XuVNIeM03m2JgicogVEi9sWskIHsxfVLPByQqJAP
wRU1l6aOKcF/7g+yOAh74E2ODqQYCDnVOaPZgrJV0PrtFui6/dkBD8+iIwR9wsIO
cFMQ4AgZuelZQPGIU+Yv8XneYIXNL4s1qL8UoFFc8a/5o6xuBFyeltmE2gO6b4Ou
wTyacQ6n20u0h8HG97sNqCdXEUVWfkdV9H7DNE52aUxdLiQoARIcX1suU+Klmri0
u2n+uY7TB8vKJRAmEzvvXIotpC90CW9J6FDxD25t5kbPj91W88P56hAQxL9I7f/S
Ganv2WMttZez4nApPOarQgFMzW2NX4vnnGvg/RWBCvJm29sgMnK9HWjUMAbiqMKm
/z1XvKo0CDTONrMNEFLlZ7mw1IM7PM9ldRXqLQCRCIZy9C8wjVXEYOqdzH2hz8Hl
wgtx+pXM1/KXw1vCnbU4TLLANIgnaUqn7he4Lw7nrhnQ89DEHllYIAMPfZi8huFY
5FTD1D/lxGGr+XmtVCAtfo9naozuasy4Fmkf251x6FQKoutDuflPjMzEMffHjO53
zngVhWN0IGJUYURBX/U8+ss2qSExxP1vUbxaRsHq6NDhL5LjMYHjs/WJ3apsr4IG
iAx6D11p0/Rhb7l6pXEoBPmWJJqpJyUP9jcEXWRxe43aQPdIaRQu7LOWSsxuXlMq
xefT/LNzYgJ3JajBMPVSWWIBWlV8oQU9QHdnNjRcnmry5ytq85nc7ce1eAYczSQH
Xa56Zp4am9NMMyiG5y5Eb6mgBVv3c95KPItIxYoAED93fz0HzU+TGXh5Jyqw0oHP
fabMBgZs2X3xLNiBCjAkNEc7zeRPGLDCLUui9HWcBAfALj0eAOMZLWdE23nmrMt3
UJF0k58TYvtpPv+HVa7+BbFLlxjYf81+frgvwNxQ6MRmyDC5QtJDTN0PqNItiXzp
fs042OYyl2ngkzgJXEYf6QaPOgcdtk6TPWx/tj6Svudaa/C37zKoKgNircnf8u5a
2RVl2sRc4rlUxpUgla+eyrBeRn0p9WE7kvouKPE52sUNlmgwGEdUyRbbFOAbnU+4
W7ayHWD83Mja9GlWFpBBg91HtwDhBpCuy/NQnt6Esi1rgt5PcPOTEKYyIxBa0evW
1ExfzezRNHx/XghseeP21SOHPnqpcDww/lYEIoscSag2pXRJsZoEd3NKU0JOeBPh
vwwMjREjKEh9MUGQU5rx9n3BB8IJpGH0cf3C1CPVzDdB6Gg0u01qqOa6XLOgcBKl
3KyE/STeAsXMo7YrMeL8j3ZJYkkLI4Jlqv2kQPEDWotbXGDw9imWP2qKd+BwfJW3
GjvJfOPjp1q17Nvm1eIpswC2AEnyMx4gPrMw89W7rPhfCr9nA56hEJ4Ml2Wd0Hhy
V0fgn1VLXtPzTfuUwqsRJkaEFRwFDNusLS4mHFKgPZbIWH4bqchwziwr2VtHhe/F
25DMYvzKuoijLfxVgYgU0qN6a7Trf/b3jyUAu8Pf2cBMXnvNU9cfXeDIIQNOMsa0
Jees8zKKibA8Lx4pK21NQL6WFPuzrii0jyidqa5EYhQjxNP0ztvqtI41uQeKGI2X
H4TDiL0TYLYA+QU3sRCQz4N/jlxzCiyn+XodNz9pEAHW3hG0uHqYt1Bo4kZSK32s
sdAcT0Rc7Iv4T2V3xlq1ts8Gxq2kWFacrt9uJfEuTVBwOrqvvVMtIdDGbgBttiqi
5aoT37J2431Ssw/9XkvsVPKmcHEAqZDDz8znlD3BTH7eRf0a6Qd6R9s1/GBITI0z
DL0DkiKYaWjt5LtMKjYHuW02PnWfoOhBJyAr9Hhd9JY8Aie2ZdeLG+bp/fqAWNk1
iYVutYYnW0v2LTM3xGG0CbaznlFcR/D//YWKaFD1dLto/qQAZx0zwPx+y01AoQkC
foetWhnExP/RfLzIWYqVaO8hcoIe/1DGkxWQZCpBFyl1ct7shKoiP9cGSHQGDt72
j22igx1Xf6DhNGrfZH8uo5duWS4CyR5ZI29VGRba3k0N/4yQXhsb2R5vQPiW3AOg
dn69WD3UFVMKWCP9y/EwdreYWiM4nnY8zV2nV7HdSg1p9Zi7j8LFbgo8lKB4CcuF
fuDI4c+HC2gM5n1vnOPJEWGqiaT4aWCD9Agj8ICLpSxkizuz8IS152thpS7idmwm
eGej+YDlxRXLCmi0/Z/iAOzQGd3dU37zohXvMn7240L/lIrxlJAMm52/E+HDcZrP
I/iDaSTCIStZ/j9m2C3eS5XfVmVqGfQ7o7jFJpCuG3VjWB40hHamatl6dXPy6SEy
/yQOglNfxn8asQrXrtqwznKhqVKYCkx1lWlcfzKaD3VlbrliRRo7MCOOKJIzXdYf
nSY5DEJBBxayAuR6cFLrCCW4Da92/wyzz0EMbDz1rYxt5xUZgkCtWg3AgEMCvkOW
MsC81HbGAkT+Kg7G8i5LEa97GZwywg6fsBVbF7y9B7Eoe4KlT4+wckbYtGh/gqDB
dfIm6oIhynDbDoMk93aEPhXsmrGXnrCKcn4h7s2BUnbcy0y/4d4c3x23Y/cxOh+M
NjHpGTc0Pghkw1487PnMMyN7UUo9GpHnW1p/nCB1r5qD/S9rFiSurOVBE8X8Ot7G
E9isM4p0gZ8YdgJq+qqnoKhHMo3nggVhjruPaup4wu5hGASF2YVdFyl68MkI7zu8
CTuHzg547Vw1vw/xIPzkcpO2azs16zcHEegcZs4vnLMngFOgo+cS1ejqZACXZmMD
99KUy5MHyShU3T9QllQrl2On691Jgd+l6XJi/yFz/VY4bIZWpzxNzTvwTt9jGqIC
OMPGbuaM/XvPCFozMJYltvyfNJRcp38IZKkFY2UTgojuu5Y4cMib/+4QcBAfh+R2
WZJjDrPBy/LyXDSKyGDWiUTUyAerKx7Z/+f1AcUQXvrFaFU4ObcUbS7z8HvlH+x3
wheukhx/Q2uUEwOz2NE5eqnC9pgBLKH1CQqLBojfB+eWSwG+0IjvwpJ9WGv/c+DB
V6ULo68pwzT6o6Op9CbLglx9CgOaQ2QN5y/oLu/PM9cCO1jpJtYp62xDj7oYgAaq
o4CFrgEKJETfYnvvDgJ58P1ZJKPxFNHObG91dKXpMHhXSMRP4dnO4hlEXMadlPLW
f78XyyrrMlyiWwe7myawHQPwXvpTN0pQDjKHGNnEaeG3UbswzY0FyaJ9ePauQD/4
PF4Y2brfkXPr/z6SvmnBeoY17E0mfgpPNEh4ZxHVT33yCGf7gFY4wRI6cmHUcCaP
69drSlCOx47KXpZi0db8OnpILDNfk8sRxr2cJvEvv7jADuMidJF+Umkg7IYPjprx
63NaHch13QmKePc9gLkDikIFpnoPA/5EZRklRZd5YPOXaF3ZkG16g8jQ9YGvU6ZJ
n7gTDx0D+IAqh5utKDXXJbZQiReax43NGbAvkjmEXP0P3zRvLbWzFD/UeU6/OdcK
5o3sJ1PhwzPJedNo/qgs75PLhNzsE6AaMTBP7G/ajprFqdCHD6oGiyHqhaDF/y6z
7l0mFzYDuXc5oAvL06yVehdhY3JIrFYynq75aSx600FANdAFScTq5KTnPsDGP9+q
0aI+xnxr7IteXF4rT1KDwtN0C95pcIR6SXRM1Sn+yKi9xH4TY4dGXNjSW+fRoHdB
SOGziHvdOeggHf2OoAM5lfkxxRZ8FDyVk6lfg8uAZXL+w53a5it7nHKcOHyiJ75M
6m95cNO0h57IEHT519ge/Fs1RZNWlD4T9yX8lU0lEqm1l81FXyC2h2aHtkOpTv2Z
GMPtG1AvzFma7wRqGCHQkT/iiXV/RGf2ayhRFk0mitMpHMaLrO0iYZ1GUvlJVaC1
QUK5c1kMOmFJVs+263+PPXmUQ7Zb/egSGKcxVLSiPQwNkzVFYQ59CU40wkP5f+Jt
hvLvdIb3t8W5vO4Z7VuiuT9BgjEoLGFUWdTEncOHWR0WrMRb6Iapux0ePvCNAqTl
K3vaHENzHAhMPJgLRxjnJQzj0YHlldDJpxHDdZqQBfxdfDLZiUG0eRVZdLlwhUXy
Zn69ZeMn0Fyr49vDmIxvWbGsXVOUYXzCaslpJROOhEb7M8wVvfcSo5VX2ur1+MUN
5ohmcPSuKTQR7rfHMrlkoP8+poxEG5uZfP+3divctCVhmIZUr6R4N5Fj23e5cj6O
8AgyCChhD6Rlkh5N7UI1Cr+wGfAbx7sal/iumqUllGMaxJdrPuuY1QzIvviNwkQV
tdBVEk8VgZD9OQY1x05rN6be89HZPKHeTHYZ0zjMkeCFFMc0wiP+ABCq2E/hzHRx
XEqeA6hZARLT1NETTfD6evIMinwL4NWzOaOZf44tURtQ+jXtEnaftO5b/drqs/2m
y81LYlyax9wExKcaMjUnw4rwoo6IW1J4LD4Qb8ssBA0DHHSZNSuaT2e++omGLfL9
egbxvs2t4kpVD3yhx5a4o8+P7jcX9Pk8qBS8nfGqwAMASvex3mFckzQs6SajVbs5
JqGK9GiUUZv1Rf+R/te7kE3CyBfWtoNtb3ImE0E7kuFphyiG1G8KEKP22XQwOcoK
4YzECR+kCzwV8RmKcmuJC4S7yquGZmsr84ebI2R9TQbAwX0AXSrepyx8h+11GQgA
W9qLEZghZfrXeHjvztgyUYNp4xFhJKT5B+88GdwBtf1cvdz8aRYeUdFcUNdp3Y6I
TCz7lxu1kKDeC1qjeDdtpQE0VI2Dhn+xcIkWz48BUyM0YJZnPNCzXbFQdUmSpY8t
QU2hh6u4LzUw+xfLnFnHDDTVbLNVo9issiYFVnPo1nd7DbbxSiK1BAzAXnl+VmLJ
Oco6fkn0QxL5Tu/l1isK7o0/HO+kDnwEplvNy729DIJgulARsK4ORiwHcyXnVG0k
jgZg1WBA/YEfPzVZnh9W6UtqYlvBoVvGUokDACCPAXByOAGixsL+XGKulvHbhBYV
LcDRNnE5HlLIK9N+Chvj2wO1MNdJZuumBSp469YWMF3mfN2ReuKFtYqjc+1W3gJd
k1h+Raw1aFhNJLA8hFqWEC+i953AymgT/UMJcjrdhNS86HQpVef4vKZWxWlY0kYT
7vFg02zs/XW6IuKM+Mg5+z39zaHGTkt/47ObjD7w/f1j+Rvz/XY/EwxNTSRLCJ9+
xLNXH49BnbCKwgMECbr/+nRD58tXum77EiVuM0iZG5Y/5d4hFxd2eU56thqF/uLO
JTHVD1MLp/Mu3Vbbo5wBs/RW3c+n8NAdtKt+7heDaV1wzQbsu1Qi/rSk2e6nyGIG
YzqJlrla57xVoMLmsSGHTfVh2b22juSN0qvc7SS07kZF78W8FCKLMJrGozcOq0Rf
6J2DRqEjYuG2Gb870n7m1v586exblgz24Ia6yvVhZxSDGPqRSfUWbDEjID9y/Gdv
sR1n9arHBkhEjAhC3ITJMZfm73jUuAQDulAuRxTwWWV1aC5lcQxxPwulaI03HGxi
6VJu+OVcLR0chO+YfD6aTDATUyM4nNXepAyxiAHmkpCwjHVjYG8cd9QHPwqhvyHi
eaBzJTsRc3KzRpvedjD+n0iCU98T6Wzh5Q6KQw1Y5R165qeJg/AvsOMLI5PWtJoB
Zmmgz+wKvhc2W/6ck0esTfHcf6tJSwgSJ478+CSiSaUBLpq+PAfXdw44O/sTpa9Z
rChmJ8IMJ3p3EM2GQLQ0AfkUUmf4C7naliwdtjc5rhj00KWc9r3KKiB9q4d6GDiK
4phNX0CvvZkMIWCSpr+0EajeDuVCQ8UZPTf1irEqbvhKBDo7lnjhTw5u6Fj3lLsC
fRWdfbYSyrlWyWVT2rFFQU7BfuR6gvlVeUVNf/8QVQ+ZXHm7ah5fTqmmNDmV/9/g
ZGWI0RBZPHY42JwK3I1l80zJpZCLSfGWsX7ZQbq2r3OdZdIXF3kvJmohy18hrGlv
7J2I1M1rPsuc2Jh2aetJlsinfUfUWY9dDl/dx6CImY0dC7BiWIcfg+cHof6riHKL
o26CVc+9sRoiTGtyPgCmFkS6ktmuAOCoikf8s70Fn4w/2ibG2jcqkFo/rIP5Kt8g
X3JSnu/pD43NW7Zt+LwuIoDlD0YSxMhlwmrA+wAwcWU/7xMoK6CMc7TlOu2MAhsV
vpTu/6ynTKW3Qs0ensZARP7VNgLNLGqD5IIKPmF20UAQTgDD9+s7vyYBxNTlRiqT
bXVgD5KGvxkcvAEYe5fTMw==
`protect END_PROTECTED
