`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LKhXNbh0dICNqex0fDM19EZmJDaZp8YPIpcmy8vJ+25HQqwg8mM0umk3w+zTXviN
ZW0+GnHasO6WTNLXTELrQNmv5FPAzRvFIRw7/bjxF6HhhNbDwZPQU8CH7hhlW2A0
TsmJ7JNTp3eDW+HnDzzrUnGGo4i9FxfMXvvEkaeSt4smOeYUnnQaCxcqtzi32Eql
YtGueosC0H/pmzTXp97BNPP4jMHty72RRgl3HMmqUtQZxXHctbsw8srV3lE9TLoD
Pb/gOboSrBUtrKf1si6nRAFbvPtapvX4++OXnLoh+11rIJU9PbZnsyNaUBZD6/9Z
25kGlyl2LbToMTSmGTvlXdT5YqGsA3eDsSjeUHs0ItxY81Dsryf+7HC8CYvBXafT
QSw1w+vAj98hv/TVL8MC7uD9lfbVWs3rE3osizTdzT01mdDE1N00dc25koscss8Y
rfBSaWp5KNr1Djgypu+fqHSMMJDWsdWP8cskRu8M8c7V71RUZy3gesgWQ7OncEJI
zk5DClygpTCZaqctq6MbR1pTyLjxPHUJZEEVgQVJmbGiWkq7rVtz3/aX3kUCoHCm
ES5q9fkXWaE4HhuWV3zp8PrlblXuzEOoBqhTTKkoV8qLubCeOZc0jBHT/CEsNgpR
CTfnT/zn4GzSr4W89Rubol/ompm2PU09Tr69w5P1ZC315svPOFz3zHxjZp1Rzob0
Wn6Rx2rsW4zOHqsvizZBN8901y4oX87Af6FNASKzmWybSkMhgcZC/+L1dwC+czrE
EA+eDWNsK5yDGoNSrmwBKOpBYwykJgn5NJ8//5pOUQmX9cOdPtcz9IoS1vXm6Gx6
IlV5MDSEZyRv6HlGQwYZL2pjHGFu4+rymn6qee0Ii2zZn0bl1J7Eqpq0OjZ3llO7
63Q3oqBl1rsl9RwvsRG9yOthqxDgXrkqMl14XrFXr9dXx8qzkvzVjk4AHcIXY13v
6UYsn+tokNyrwl61E5ipo7nz9qifi1L6Tlm6GKutxZ0DF05TGYQfopA9+WxxkHXq
Ptrmztdua/6dIek8MF31/UhUPlWF9V6uGdUDhmqc/uRqahgjMHf+cmC74uwqR6eC
eB4qwR/Q982VDsSv5thhiBDEnUBgb7lyOW5peIX87P7CbO8D28UGbKAwQ18SBqTB
sufOrtEYkgmp1wppxl4Z1yVwToa4CMG2+KNs2oQEDv6A6gGVYk8cpqthdYsR3tyC
JCMWavcDwDlP6pzc/dMia8YJoxT7jl/BE5Czsmn6xKGyAMAMTj/JAf/DuTaw2dzc
nQ9TIpjMsAvNAOGVwspATIzs3NL1dtFP9T6GEDpLATTP06PAnsFDn5oQLYy3fhvm
bwyYkGI2H3gUXaKT/u8ZyKEFDx/gGyeYNT+ADSTeycu8Bu0C9tiyDRuwiP6SZNbC
ZPp2in05wxp4gqUF9/VVS5X/3NL7nLv8k+NDQrVninCsk931K/6L+xLIiylxtfJc
UsnH9RsWi1Eo6vNV7Aiyj+HkalGHsWUQhQ9IpltBC12gW5AGNRxkEysIvM7OWe/y
NxiYStVRusD4eQPdQ0LQIPWleU4cC3PoE3lBbty4nqY3xrdEqtQHHY9Xq1JO2RDK
C83zWB9D1Z1HSTTx5NRf8/XOy8wlyFwWs9TsqLCYPm4Aoh8Z8td73Rg54XA/JaNW
TI3e6fan4RqGWQy+1u3XTj/fhHR/dLWaVb5yFNNEVAu7HEHa8N/FdX2oCqVetbTr
+qg+mGHMVpH4DC4EcuFMwoCAoj4aPoKJysj5BeTbyR5GtDx/fAmTlCdM2Hsaabj/
MN6L2hWJQnmBi2PKuo/Tzquyb/2a3FJoi9CE8NWATCMgjuoE40GKzr+/Q/Od95KI
7RgErER/XiQC+P4lXb7Atj7nv7CTB7zpkUoaaFXbZNQGkWUYgz+to6eVeVXpsNCO
aMexELMM0RgOcf8w0eo0n+g9WmfxTusHmYJT9ngwGmvqZ9W5chDJ0N9RzzpqfWbW
Z9COxAGZFWTSO8NYfGAIrNfLQvNeNZFEyuHlhDSlEJriAXnRpPlVMbLy+SOw8u9E
xnV9jqgTLvDV9FjjzlNAVLHLLJ7vM9mrkF4KnQ6vLgQNAjZrPwPjL6MK/PL6x7Q9
37hhIq8La+jdHw8NRnUJzYpzOys8nO4h6UsZWamjiJTfIcl18JjBDuEI7X0APXXR
zplmQYQolUqhKbBzS30Wn8eQ4lYvFWUOyY4Mwtzw6MyH1M3PyGuwGNvyJGO09FbW
b/ynPU5R5iWkc45gtoEUROJXSw6wQMq7w5CmyflcX8wCEnoXMJNOSP7LJ8OLZnxR
r1Z/uEFBBaTOSCgoqdVL2rogcjtvu5eFLH7AXNFaR46g4TLLUQS7mJFEq1QdUruT
UMIdhFwYwW0rDIC20NbnURqecnUf9aIJt7RqJEA72cnHL3oNn96Je9ftFbsfovl3
pUqoH5QcaMUCjaCpSh1NJj4IaK+m2XNJAHZb/51Dr5Co8527gUsMeFLspLC6f6Ny
9vy/jfSYYIKy250R7iJMT03ibH/erwhyh14sClihrvKIT+ly2ineUYZQmaLBKX2A
d6vYDL0H6PyVuYQ53XaeN/JTHeVMOOheANitE3U//uP06TVgr2oYp1ryMK4njUaE
0jd6DWxdyGji4lYcqCMavkc1NiDPrExyajIjv2I4xQfCUzU7axEfC0g6OynuTn1f
kydki6xdc9503G+Xv3/+dfHCO+fJxNl5llgWriL/8HWI09fOHVPVc/Ew7IQaWYh/
N/GaDjwYobyHcv1rzbSE+NHZUxE91Ik5di2nPO6s4MgUdI/6dxwOvQKnKysooUNL
65UeuXBaDKd1g/6mON7msaYgRh60D9tf7TEsjdxhwB55Co0yISjEc0o3y1ZNPHxO
++bDm0F3mPX3KKdXK9BXcpsFlKgci0Fq365VcF6QtGYHvPmANc/LVH/KlTHKb1z3
yuztwzBV0DsQFi0KWp+wsdP/bpU85nThsGwOh02znhonN5FQWcJjy9OPzUYSea8z
AaP2M1EQ3kmtQhLLEkf20tg59dLEwxgKvn6QRIvv2lsvhDtgVfZMtvAUdn7BpNUu
NjxcSN5zdolx7nQyhZfqXUNq19esHM/AcKns9DE6DczwDWZQHp0y9EnJZmxT/gY2
anm1ab+A5OuITlmAM0/9OnZ4vnrMk8VmVF01W3QG9F3w2Hcx89Y6l6pbCRiWBnYQ
yxmYv1Ykx9Q/y1kcp8fPelgeYpWseZ2ai/T0Xqrkb4esBWEa05deR90EpmI1z3RO
Hzw6vKZbc5FSx7Jehk0xX+Vk4Ew9i8gdIYv9hppWF4m4b2JH1yU4WtD7Dw+K7OD6
O3tSeR4amIwJHILeltsTzGW30yx/bvuDxMlpi8FHVBAj351r6qD0xZFFUQypx61q
XZ22C34Z8HO0AgNTpW+GHD7BY3Mrch5C3n/Aifr5U6uQLGBnZu+/TlBCkTNpBNP0
X9yiM+3D/ybcV4vfxNYpPdbPOYr82T3ci/sjYIvwwRlmOhaG6PX86mgFGogEVLEd
t4HR+AkgrLbZEowV2v79LVm6g6d4KLes4IUBKC+DtPgHE6bdq82874vnXbE+dDzZ
a5NzAAxcR/LFqK4uT4iuiK1i43Yzm5dkjqNiRs0D8tAqzATL4CGLrLmduOj+Pwkj
oZlujIenlhv0e5gk4nQUjQ==
`protect END_PROTECTED
