`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/37Z1D2NFdlI3UedxWFRDnhSCL8VnlWsteAnoMVzLDVpSsykwYNKR3r/H2u5TmHJ
x6Aba0zJZvVVsvACch4X2lqfhq4DJ/j6xR8FplcT4rQVEzvbHC43EheNSf4TS8TZ
JBcEFJszW+29/bqT8rwWhTw3YTujFrQE768+IO7xHbiqP22vhg10fnsTDD1eYpZu
PAHGz3FAZYBLkKE/bdeS0YJiszDybQrEk0TRQ81rXSAs0kcSLkV0p6mJKVv+ghi8
gz5lPBuQAykxb0zbg0ZGJvBFq0/6KzFfiLrmX7Yk/bJjMLJGbWuEU9mGoMyD0vVu
2n3vCyT7xWasxdT6y45RSjhVgfCKPCmNkklu6zhiwVWfTG2P3P5yE9DUAv7y3rwI
/EqCNUlcmaIA1RaSBoeZxXC4IfrOVr5PnvaE4Tx5lKIOjrHkuT0/Obx4QDHFSWtc
c8r2Ymhb6z03kN/dVddL1P6mqEXia5bcUhoaWKz613Crm2sD+vZ7CFhYMqfdKa6R
`protect END_PROTECTED
