`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5rFLyR3LvWGsQosKGmkpBN0QPjXXt6ROPll8Dt6844jCs29cOjHbr9No1tnVr4XG
86Ki/o/Az90FvUGMGzsAPw4HBTv6a1Gc6pWqfkn2lCcPn7VstfJ9HSBhAtpNXAKf
nyKr3KqQvrh4m0+6gKzT+X2IA34W8AuZ5hAe1oS0YLOKm7g0StQOh3feKE8hZ/9n
iG7c1judknbrGHqg4YEK/Fz1ejuoq+zVd5MMXGRm6DPHiIuXcNA3C3hRFg1URvTh
sgFQQVWKpqWN4vQuRKlw8nCV/1Hu0ZbxD3Wzklpc0Od/KbgSfoEgwOOsqmNRaF/q
81g1eRHbX54IOYs+dQZG+JGuA/9yfZHyANzAnpWNjFjjJCO0cMQT9aPEqz4G2CLT
ssW2X55ZlSPTHmx5Mw6igw==
`protect END_PROTECTED
