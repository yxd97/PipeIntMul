`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vAXq/uD6rvHYOToa1upAvEmpVwxUBo+uIJlyvwKkvTOAmlYF0WJ/Wa62+4kqhe5n
X02FLQ8+MW9e7LWWarGE8tMYIfUMFJBBLQ4nO9Fdx94aV3rMOW3AgepxIhOLOwCc
RIyTxusH2cRMrg3k4rGiz+91UNg0uIlYHjmT48veGZDZq6UXaAM3G+DcIgj7Uh6W
rKy0QaK5HWwtsFOEb6LZUz3oWyhGkSfLruAivKS7D9TyLpfXheGIy0hHFHVV76Vr
DcCT0GtPPglfoenDbWF8B+a/x2WIzFyp5Q2sjDkWvuTVo/D0CGKobbhTWuN8C0rB
IH3uImynlPqkijven2U6Khz8Z7fEFLY0ZBOM481eMqnuVzVcM8HGv5FxR4lL+qnr
unWrvvzoubLMUwDXM+ZamcxLnROn964b0O/hziV/qnw+GFyD5bQmqWyPKAK8Gz9c
jXwoPZ4hgtoRu/Yl69dnsT+NHceT0Dw3DdTW5rHuravN7Ry8GKBwD3y18R61GmN7
+i30cF/xgf/FIGi4FKddmpm+peiEhu0i9h4j5Opn7me0kALyzVeTbG3C+NHTe5W7
vLji1r5cQ5N15+0mzvDw+H2shnJvvj+jPhaG9z/r6dxlXUGUGfJOprK+HFFzCNxM
IMs2qVnSnoi9EBcxTs6FhQMlUSfd5xHtsbCQ4/pR9iyI/QIkvT6gJz5ro4dyMMa5
dejqnvUsme8+4CPdIhPU2PD0/NMYfYWPVvR+ewZr3CCNVJvtwmSAXxyzdmF4lW66
d2qhn7D7iic0gONjDX3fGIY6JuPVg2KUBJCLCaEY2Khbdz7ejjYaDNmQTKCM7r2Z
2SBTdMrBSSHEAUjkZYFAprMO+YeG9sC1WkTGD8N/NV7O0B4QE8M0T2DGyOO3W+P/
+8qnvC/hnYV4LYzcdXprPY6gKFXASCKPz0RO+4Rf1gOdCGnEWHyDH8cAuJW5Fkn1
JFdCVt8GOWmV7+3+gambcYqjz9YSXzyQ8Iw/o3gulgCyI2GlhObDvtLeEqavK/Ii
aRFdE9BtPPZ7PJbD/Vu8hEd+FHL3szzTkoJA3pFxZw9i7t8IdivI29X5Q9xMx3GQ
8Wfvn9WvyBICEEhkuEeHErf3+uQTOCJbRzfUl/VT8q/ig9MO8C2I31JwlUUuvDaW
zY1qwziYOEM/dRuuNqZNstq5TR5ah6fsxxsAjUn3s2fwJG2cMSJLC/jRYyLRILGj
H2cVF7nkkmDnz5FNXsZ6lkl9fV+EjZ4O3r/VEjrdgDfCxtq/+G0C8xgTbL9tcFps
fTbDSDxcA1RaDM8JyCC9pyp7rLpezb4hoVE0FA4glL7bZ3GFg7UfMIS3yq08aS0t
ynXtz8a3uzBpC50w+waXAzrKtNwX2KiVYO2aVP/PzHVERVTowWq0XLsYnXFmo/Yt
NQftUnRNcrWh7bspktWfiPg1p8oHBTFhaR1IAQZB9C74ocJXjZxWfim8+aM+fkja
NMz/J78vKXfycr5flKYSVqskg8/b+mLzip5guPQ1g1seuZpm/W/p7J4UZK+HS5L8
KdwqjO+ATSyNMNRmx80cloV8mhhs54LLE0VKcAVGZws5rEI7ELWVs5uztbvXXY5a
br0aHYqILw/0wyyxyCrzKyqxjAo1mT/ZG8gWAd6yqfkuGZsyh+qMnPdaI9UIJwvK
yv2tH/l0mMcsb7gCFvT1iGL3/nFzBycJuZy5AgnOt/4SbySN1lODGlywClSXejAv
DC9qTDTM+FAzf1WA5/KC902R00Mb9lsACZZnVP45EoerHd3l7b8P2AQFoh3JyJOR
JB/3FDduGxoJOlJXVearlOU2va4jSl0Y+VXdtB/1+Sq3lQGTQGg4f2r8gyJdqZBc
2uqtHEzN60UtunxE0bjX23cjyfZoqk/tuqUh1u8WamdFv7EmYrp5Q4kVealwIFpt
bxXTHdEMkncN6QhM+wxdpNgWOiAtL7vZMzATJwgjl5l9MjyG2FGH2TI0Owqjbvvv
saRNArFMvZfTn5dV4L8ND98IznsP1j+T9t2vXfdbzQFhH9X1IP0bFRyoyH8fnj90
GzR34sHRPlcjuzUAibGFgbrzfWzwblEHOEWxn3O4AWQ6scDGz4PXgVKBeQn8px6K
lm/4buAj8h4k7UaROvy/aAVdiw9X5EVEmZ0RrNKH1+I+1lMMK28I5kmJAFyY/iZC
b0Z04RK/2XFcuXMGttVR0gCBWSyimFUO28MlQSTdTw4zAc1RrZwq3ayEaCHgyJVf
rDtxUJmsgN3ZmUAeNdUTErmvPfsdVYdjchCjoBhA+aMF+cEVtJlOQwFySh4JIEYv
w+6mht1SPTtgXL7P8QK6rE3U/a5rPMM4EXom7duJmeFO4YKpNLGUmTu/NK7Ggv+V
gFYi5183Drdcz1G5DTVTcB8Pla9863tM/blPqS5CSjWS+dZeWhLoayZMixzObqln
DnOX5tRwqz3ib1ltiKCaYKDfdoGVVDZDmgPkk0Q/TNlLlYPD7hzG43lGhEwuwfpH
isU7YXBugwBCts9UBK4ldvU51d3+dOyj8TrrZARK6Xwl89xYgmEEkOaGEKfd3FbL
+FegvsxX4ZyMoTcEDP+d/XL9x6uX3O3yNE0bAry9tIIyWKtwjSfa3ebwQMlvgO7e
z+b4mb7xZsFsAJZ3PjkBpeBoR0Bzj4lO9GUqRZICHTSS7zcre6aMM0lvC09c4SZ+
opyo8ZsjSIhgqvMQPYmH3iCuFVdjelkadsvTlYBzyWandOOq1i/0mvT12xhWrG85
/VD+jX8tlosNHSb4hg0WDDEIS0tnH1B3VS9Zl62G+zt4wCVyIzEXhBNEdypJjlIo
OajOMdq26OFwb+BEd3EZmEK1+BWvY9YrtG/vemJO4uEPK9sMbM4vddmVNxhRPjt3
4+hnwreNVSSVa0HeNl5WhbxVZ8uzJ/uoszuK4fHqLsENsIP8vW17GIYrepuyyhLJ
w45bMG1vEJB7jtRN/hdRNZyybM9I/AIYlBzDPXy3lX7pojTR5NyEbbu107E8Alrd
HgIqY92q35lLggw+DWRxMKwqPFl4nFz9pfSq1G346dKvudpAnEjAkb16H/dOspjp
KPum5cpt02HScLonrYfVJ53ju8xRROkU6zri8UxPwzahFjEH7b3wYc5rgLH2S02t
Ekd3acZHe3AJg4PVAnK57gfnhOel3FRJWvNWcQhraww9msxA70SYqJZ0HXTK6XZX
MElJTJekI0FVF5X0O4b4LtwqWsrgi/ebDfGU8alewgxUYRNhOHPNRQL0SCkaE64Z
qnoCOw5qz94oTUrP6ADeOKyaVYRRD9Rm+oUK8VRLE3Rr0DqptbvTIUH97+ih+Tz+
0071F//kvHGbLN1hhRQRIojRWFNXcJ9QrmFYGe7vl0sN8ljFmDukZ4ucPkbxKEPg
MTKRfkBasspzJGs/5tDsrN/GLyG8I33sM2+4tI8Q9keMjNFGGZ3bvI5AuE1VPK4l
sPPPm8reQP0tEEcmuEa4rmMu3n86ITMXNxoYd/lkcFFsGajwSRqJeuqXEB/DSsLo
Dib7g008GctmgpBwmdkMyRs3hl8PkOkqJLMTXEZaZ9biahEHvl+1s1eCaoeMUpBD
OGfVZkvTuGuwn7drIW+PHMLk9p/rUIHhyxsH/ece2uwBEoEyO4yZ6TXzLQ0b/0f8
x4QivaxpUeqQLU+l0i2b90rqRojGxW1+YxKKRZ/vDR4vNJaXSsWGFdqpeddQ7gX/
5G1TOoemkxV8BzYGFaoyQuy2Dn1EKf9PE7smVWGpm7p9+MBgQWvEvT51gvJHYf2s
bm9TJkg3N8ToCo1eJQAlC39REx9LtOHmEwXo65umXHBDvOCsVrz8cZ9SgKBmdykX
TY6bQNRuLqYTVpVtgDcf3LmSRCM4Gc8mu4DuARd+6kYWn6ywXef33KJahBnKfLn7
Hoptsfuh/+5gjNavWCfAvAXlttFw0amcAsaADNJ/UzpTQ5YC9paCNqwDb+QmjRsu
ycJ9PVPVz6+vxwm1FLxDioo0aUf69Ip0TGHeJepBAdVFy4xkOjFeSMsHEUsQ/Lck
i3DF49Qp2s/4D7KE1grixwqSvoqp5SFZ4Xvmb/Lp5ZSkrzfTC23pBBC/tDuEnfnf
FixHttnaBq1hupLtiyD8L3Zf9MgD7RbwBh6wfVKlY66woLZ5aQ8VcF5P/1bfOWvX
ShITznx5PxaySMBgoljFVi2/0CzFUL4vRTrQWI0SgQnY9D2KhVGPiLqNTj1b3iHF
djbh/WjRE7Hgx7bYABUaJYzAOBveRdgAGj5BSXGt4oTtsqj/6OLRyNos6f2ASVw2
owvnH0Q1Z7eMVUgFTQKGaf+v9D7ybyDw6YJFFeuiAXEdCB2drkx/CqHp3piJoR5z
cnbx0qqd0XaE6Swhr1EIQs49JyFaMm6zEWr1YPqz+iW0ETnvkW3jJM1rz6QyBSbz
kFv3Zycf4nNUimh/n/fTJOVMVtj22aTNRMhhcoY9tujChB05AY9WM79R6HSq2Boa
2wqjnc3tg5TWOxWvnb8vZinzZwZlB7AWXtl6dhHPUtMNqjeus7zF15sHS9yiKl3h
b8dVq9tqayLHadSz9yDXc90z21IKTmKZtcqBZCjgiSG2b5+5qwDT6dTkfRjJiFLb
UKZuxNbDL1HNTQF3OUdGcPDgeKJoqeWwrN4xBJdRqKYy3U+oPn/yvnYlYj50IqTk
6EmJ3fubnhzswqaU8BnvMTp4bsvprJlZ8dhJxmuvhzvoyKOvO/Sx01qY34TOQif9
cT/MXDxPnO0cszAeclZjmMeuTsAEMlpJSg39tHp0r9F9aICD6R5q4U5Z91epdqAK
y+YQLPoMxDil/cQVegT2HA==
`protect END_PROTECTED
