`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mD/ayr6JbIj/WYPlsK8bPsyLPmrB5PbdS+LfBNJBRwl5mUIXOlvwWd4Vnoea51Wj
L4e/B9mbGSWydnrsb2kvIYwK03imhBctz5M2hIdGP7ZweNYAwtSdXk5K5jT+2TR+
zp4lvCbEPZhDnRZ1h9lDRP9pu6rAzgSD7I/tui3DSHkEZXYo1wBh9Rjulw1VUzsx
5zMki9AdywXCHNUINzF6NMkZkOEGyLO4g28FEndsLKYVMI+oSFngubYKqFP1FkBT
MYHWXua6/qDf8EnGPBPbBwWA5fLb0KcFOoZTHTbjIFfQZx8LxAHuJPk68TISoSp2
c75a3ReLoSuJU4Opx8YHGLbSW1fvJ8M7ZL48acMBnm9MVQ0hbcLUWAAfACBtgKuA
SOZA6ymH5cPqqa3jYICJeaIkmnnbCWse9wmCpGjfnpM858zDsYD3GcWbzLgGsnLT
s019qM+asDiG6rA/v4R/sjuxoC53spvf/d28pzFQ8arE+bj/zqNTUvuL+CxJGSym
b2F3EdRJMU5tyFR+HYvR4x1dlqq7ZkJg7eIw7K8J4SdpVrwg5kXc23Tiz/6Lt8tj
w9GXc3znKWj8dork1/AWd10PsXEGKCE0BrGW0Vkrn5AleHV6gqGTH7XKKp8ucAMR
FIKskv+iEvRHLPUd5NiJV9Czj2ckstgKg7+HxvOvilUOalTY6r6/Mln0BEBz2zGr
7ZwOYjyTLnDWFJ33f3Ls1rAeKgElJNmkac1qZuuo/A8j4qfnCTv6NjyXEvCNCVVR
3O7A8m8aMNUgkpj9Gkn5l6PLnHzACq85LdZjh3gkKYakLAhT8xU3e3fOgASxb2Et
CC0jV2CX91xLTpUnCaR4lyBwE9JKFccUaFC61gLJe7/yVNEJ9MK2ufWdXavjXVq1
DyBuFJYZeyu9cnUl/71JZ03FmtCkdX+Oha3rg9Lt5r5kgbHskJDZbn8d6XqEfTBK
JW0mWU/RMXQR9A3HAjxBg86DtL/tGRvHpdv7buvbBPFoRgnoILbxumbHXqhJwoUT
xQKLRU367owUr8cvy+oUeRgBwXW+lgilw0M7jgXtarI4P4EutV9ACiwJPRm6yi4q
bBU+W7CUAHiDoa9t32FKu3QXn4fWSDcR9cjbbYSc5pNHML8eNWs4FujFfi4va/dk
wD91sf1L9jDoOqJ20DPJn4Kk+63DkWfnJPT8P48SpBgj/Mzl7H9zM6NXhv2Hvo93
hA02SmRVB1o2EpKs+6MyUgR9tTrslI3WAys8PBlIkawzZvUOT116PtjqHZTVurnY
6Uhu2YpENejXCuSvQfn5r5a0R9so1F0nNOJx3syqEmXIyrSmWXDbdFMuVSbwE/OC
Ya8/g02rqM99ICnox5mDvBAeeCRzCS+btJmsI8KKf3RGIKgIMRld0VbRxZRooOFr
+aSxsLlDyU2BQ/kim3gh1HEQiSyOXoMoee6oqLiDC3ct/ERloxx/gHL1CL+BVRRD
5cnNsjTGrsGoO+Fx/TDk/B5xhJ1GqXh03t/7G0PeYNyyyegpdGrp3Ivjx/fQ6s56
dlPimSsIQhEZ96Al/uf7b4V4Oy1SB8ZOvwiFvkW5VrzwubP36HCNEoRRqfUcUf/l
V8ZYgMDuzw0rFPeAL6ExNuG75/1MqC93XRJCGOclPv6Wzlzx1r4DrFweeYPzbjRO
xsjJdf/SG1eaFTuYFR+6M6o09n29t+Cj/VUs3mN24XqV+2CQOAGp8MC9z2MK0p5p
9QY2jrl3Y6HA4JBrN7kDCrR6ZeE3Jm+BrmjMW1lG0n23WjBCTT5Q/j3Tzx3XBGvS
IP4UlQfzodOOwpjLdPomMMsqolH6gJkN3pc+psUHSr5JbJVMW3WkFa2TSGBEV8MH
MIOPxIfas8cLwr2DHuNCRLKFXSuuJALVs2jSkjfNsfFY8Nl8+2/4Jpsz+glP1i+j
61b04bt1bqaPUdnl06Y8Evd19tEJg8uvUajDkx/fZ2O2Le1aEo6vC5i6LuAVHdSj
Sl6AuDqMnM+jZmpdaGJ9fhyG7zf7MRKu82sD3qTVop2NL5po9Pww2irOtuDGEdeG
Yk3VziJdhh6rE4JVzle2XVHUCC0Kb2T/sSkBz1DN6e64LALpcL7bqFcu8z0AxvEn
3Ce5YLt8aNPDkbgDIdrEnYo1qZveupMUn51SVhaFpQ08tSiG78KJvnciHbBm9xfx
RsWC/q1p/zNZLGVOva/zz813WIUg0Gab2sho+1WPKWVN+FKAoFe5N0TrjVjP3G4M
0+MJ+Xh7iDcJt0vw+oQNibe8EfbFEbqPdyP6k0kBYhJEzpt8Q9AJnSPtyMumytg6
HshS4K2FaU178YQ8jtyONsENrfV4r76RhXRjumqwHgfiRYbUVv2YUM704yQaoI2R
I/z/pmf3Qhswf3bkgWuK0hYXT0aJrIYbtW1pM+dHnSWnmhSR3tvwJnTBgBoE5Oi2
1ncKalrlKljcm2R8LM4p3hstfRY4pQOrY0Js+5SIDP54oilHLmu9NBpSeE2lsNjo
C3zbIS15UxXjylnWrAkNJzs9u6XypTyOKQRdSnwJAnkaHTqPgJdumSFuT2/IoN56
qATboLeuH/8v/1xfKx0HZ/pCXQgP6gATFJaimOWLTcA9e6+Tg832ZX5NNUe8NS22
jo4YZN2xmQMB1xtrWsm6aWkZZtM8Jkw4uNY2yjQPe27egCxQGyOiJdVfr5n08E13
`protect END_PROTECTED
