`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SAJy88i3nidlGS/uC4W/FIqCae+/bqBOQ+Dm5Ej4G8zG3E8T/ZgCPDu7HLHDb04n
Lgg7PXIDqVryyaatjQ6b5qGx61KHh0FP7Rhm9ZsJyNCNhOeio1bwGpXzLGPy0tf3
5xLe/hHVd/vTbUMh1bFT5wECe76I6qyqzsAsYYOdYB8uHI182u/K4LMaVcWx7Gvt
VMPWHhIkXQ9IIknSNAwYDZGEc1EwlpeYw6R06Wn+ax8rxmOA22IYTcMMcxerklc4
ACOLIqkY7VepcT7LYkrwuCO56PFx3m3cO97emxdggOqr17GBQbQzlt96E1Y2oJfZ
PvIs7fsJmIW6eZjQtbuY4UdIVUuoQfUhVpkIuxZ9/5bp2pNnxX62WwIKuLJ4qkZk
mdCXtN34tjrxklKJP0e0mA==
`protect END_PROTECTED
