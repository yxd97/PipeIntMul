`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XMKMvUGQ75q1Imi/G5nsO7Pjg/j/aXZs/proSWLVHQ2BF63Sz9i7JjdaDzm+P5AW
N+DdXpogE+qKGLhqr3QqpnkUTzZ6wIJ0XEsvPQ40pEzmlc5EJU8E/Ge5xMN4Ke+6
d6amTGlo2UztyUwqkUtZ0m6UCZRz1TU6+u79fksZt/B7Ip59oKoNgy4uyV3pXdQY
3MXEamO8XB9WF8gerVc7NGcSovbPi+oXF+Mi0SspPJ6kOH0vePTWwu3RYb0doREf
QWrs3Q9qV3koRDxYEO9ppuh5wc9AeMTYYI7ejaePWpNW8apSwqvO7p0mjcB47QU+
`protect END_PROTECTED
