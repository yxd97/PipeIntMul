`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lyLE93UnzmHN/L201aCDVIeQP6DZPoItWfOxTlDbFol9RiOpR67TEQHq/VQSKHOo
KWCYq2+pqdKf50xIf9x7c7ONKwosnCOHqYhXqZqWTENkIbo+Zxaq8wtjAYyhNQox
Xo4xhm89nav+J0aCHAnKTZSXSTpeOXfx0JVfxtUkCTQME9Po23N4zgN/twFrISVv
9TEq+fWg/mSCS97pTMK8Gf2tq0Hk6luKAA3hnoSPv+udlRAvh2Epau7GDkAtN3u2
8EWMlM/w+Ha0IiWvCEPU6K8f7VC0pra6CFGhSzMHMYL0B65tfckqjIm8gArrbYax
Dm0M0Ew9eiijopytNAbfXb2M6vQqEl9Pn3XchW7VNCiYkKPLtFQCAAxEwTABnIRw
`protect END_PROTECTED
