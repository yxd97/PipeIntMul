`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q7WYGYiWyzMyUoEJLMJz8dSb/HNgX8K4kk/izxgfyBEmKfVWDluu2gtSqFVIj91+
p0ZAMDFAi+ro6qRyUQUGVo27laRmKD8xn+8IUTs6qtsmoUYTAQ9gZmXoO8AL7l3f
hycqAoRVzXxOH77KL/GWUF/I1F+vhWZkecVwaaqG70Kmq66imT7G80Yw9+bmFMkl
sJbS34Re2vztxqF9D/dDv0YMZx0kslDC1Mt1DcR9Ch8FGZ3MWfgZZznWbJ4Pmd0h
bh8WdOJHxXI161CGl2oeH5hOnraRRv2bYx51nSLmlBQMbYKqhgqdCQNdDt2LzY+R
ty26PXT3R8KLUMEHb396xq579ZfXanSFSgVxNKUbFArWYGo1GK54deiTi9jmBtqx
0uhkbqOjTLHM+e/544NdT6abUig9Uq4XavBcNqwSKQMy9tA42wYs3vcveipb4j5e
lbViIHcqiLUrfqStu1dgnA==
`protect END_PROTECTED
