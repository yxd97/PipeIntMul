`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xgwHZbj87Ktyq+y+f3OuJMZhGiUqj928iB8qy3clcc7EFYZvO21OgT13t/d/7Q2L
+JpJfEoXoe5yK8SNv50JrJs8vcY+4r/TmvX202ZK7qM1X9Bos/50JatNeqiqSEMR
GIWvDHuPzO7I1sA02omHUtfPpASw9eGHqMTCpb/wjOxhdV87S1UVgvopEQsqEQxV
VZPWo6TblzS4GdU/QF6KU2o53uDzp7QNs+RLzYJ3ej0S0DLeBXSwMqgPyGfnebm5
PwEkadKZjybOUjUaxONTXqqZYsOBycNcX+IR7gc0M3Cw3TcPti2d+G7gMBesyLKx
Y0jO7WjHZe/pqnabzaPT14xMla5C1vzdq83hi2JA81M3LeIBRMcYPFcj6D3PMglP
eW+9PfpUV72BElWMVCMk7LNPFjkMfEPSccw4+aMruLv091NE9oS8NrLSxRceVtZk
DY3UD3QFZt77TU143ua/gAdhcBsMtURf5X9gG9e3Qnm5auJZUzBkX89q4U1t/43q
EeiqVxKNkptKfO58f2so/jPdCYQU4dE+Y8TDzYk86y4zzlz6Gi5vfnL+c7TSfLC+
0cOeDfugV3TPxRN9EaSW2YDmEiIzVZx5407LBZhOenkM0MO/MfN5nLBQcVbNhs9M
hqp1F/8pv9NnD8VrGeu/GhhDdpv9WZT9dGRPjXOP9tmPhFlz+96VXY9Ama8VxYdh
qhkOBDj1qbVGp57R032imSI3YTtY0GHjmR4IC+4AbLRWxr/ZLMs/IRZNbNzCiEUY
62fQn3SJbLAXFHWdsg3x+FBoVZ0DSGDaSG79WBW3bWOnJigRekjnu4OfyehsMJDR
1RR+G6zkFOOEsu51cvVG9CCUkiwrS6+doLVzTo+FHaWWkhxGflUUMjGWUdScxSP6
B2GNDdzWK4J7OVUvh5kb7q2SYTznZg+NdjTISqUVFNfa2j9VQF4wN/nP0Ipj+3Aa
1DlEtFz0y6uiFaeZ9e4KQHqe7zRfW0URy8MlSsLcBZS+fWO1KeNHS1u+1z6EZnhu
WATAmSZoXqQx+IE5RtbuWsWrIka53elvoyx0GNoixSiAF40B60XpiEKZdl6l8KRD
FpP2EVhHuW1rX7NpEYTu46WwGzmP/KurpyxmI9/Qcnp+NkQdYcC1l+X7LlJheJJX
nrt9KB1//Oq1POkllKb29q9/k5UDe6rfXIsAeKawVNSucmJV0bq+Qc+bUiTfuyIc
pPkUl4JAwk2XYIHYmlNcs+f6IjAP2xJsAAGu5DimnshEDhw1/MFh5LY2GuihqeWZ
pNcab7ckvUE9HddmbYdZa1sF6m6mNFtyLDU6qgJJlm/o9iarqoxrCrutNyiY+jZg
A23i+keEC2NCofXVyzuPt+eepGsFMTDx8gh1G8g4+az4KyW49uRxwUM9r8GZZRXX
DSLY3nxaHZ4HkYe+uAMiyF7G20JAmHGl4tdKJp0yCBI8xi/alPvQte5mGrfrT1DY
tYi650gKnC+nRySG7eHgAG8nxX9ezVriWeQOpU0ArshMxP/3GcZyzeYWC/M/Jv+l
lakrBtGKkDVzXlPQ3/R//zUZht48rnU9WEp8vQy9G9fr+45vmJtsqA5NHRvkZYKu
EDWRAkGm0zxWu1Mfnbm8KlEwF6xw+g2lcBMtg1ukLT66USn9PemjWphUutsSx9Ue
q3TVdunXJfDXT21XuYeVMpceHwDn6NYuNbZP+NelBhdvbFiX62esB02Fr+DQbVCU
lvZvSM7Sds8KDWE2dSmPcjw5RBV+jOCabVX8zFJCNHvHjgZfqSCiEIA4iL2ou6Ts
mDp9gWNxou/2TAt3+wxhOB53QK2H31cl5OW1dRT+ZsOf5bFnAybVest08Z8gaIdi
XOwObNLx1XtjAZeK3etOCiD9ccoQ3HfCC4ecVjtk75N9Stb2uPBaVRmaf0f8vVWD
QIlUT71j03e9jMtYz0uSp9RE8TEoFxt1K/Ki71ro5VlbsQxgwjCVVt887J2hLso3
fN3kYzYMVncQOTvVQrxyneDvoMJKm+pUMsLoGfhx6g1XPDWUuZ4p8DVdWm7461s/
N9WngITPSi7SJHsQN1COiTSv/XakySyny4vFfgVyZLrjatFjMmi09KvDVFEeZB3X
nMf4an0ElKo06FZlj0CqIdBI+y/2DdnIOvsd+FUV5VZr91SzbZYd4Jav3C+VHEsj
RW0ddRMC4ff70ezgMznpuLId8bRaStDT8qvcOv/zBPCAG5/SH80Czp/WMTibfva0
JVbYsoiXmi7iMDcr68nTabKQxEcaKs82mrCuMrBwqugh45hYWelTmGV9RzKLQefb
6F4YickOdMeP7BMC+Qi+DMuCu+dPXkeqn+Uv6NEAbtVt8mOEgifQqRWrHH/0EPUU
QfV+UNSdraqQaFJYqHJAbOJw7DS+wIHgPm1ueBMpKtFc2Nyc4MX/q/42yKCLX+Sd
1/QbZX0AzPCER8mR+mhQFAF5PbCbmlUlC+yxc/zeuwRWv1VfCkvoCw6dYl9nnhsl
sHGepwIGkG5U1UXenutzC01kHc+9W5Z9PmY27UXalNAySqIuc0s4mI+13T3mhUH5
zcmfZO7Ls5mnAec49hik3UAJGIN4YiOmYQbMtzxuTaSgscn4YGfiSk0OPgYJJ817
R7x6XFuA5AzrajULlXvTCmlHZvrRto1CblWXeQxH+/YxhEy1WFr34Tigg0g2mit5
Hr2hUMGjB3L1UwsOkxPfoeUAt6HJmUis8d9l8oOcwlfbPhsoZ/QXS0+jofNnUy/i
z9PqeArt6W/ZwVqXxAmOzKhZoP6ON6wO7N2CT4iKivVDox2NhfiriBSqjbyi/OP5
Pfsmg3PLO0HGcSyepXDdXTDH+Dxtckxt/dQvNkF9KBAd4x3bSMYVzJqWo6quMjWI
fcH/Qd81/OF5TtFk7TrYOnCHzTErEm/2rlA+lOODPxhOhN0DfWiLA0qLlySAyRWt
uVP80jctaixmB4G7iCVlqGdjDOUOBKnl/BlOwBtCshXbhbjE6UXizZ8lV1UQ2k4y
OueC+d6GaXe+BWhnaZ0tTq4viGUaySfsXzBt0dgUm/vXIfIhN3P6XZ+RlJzST6/s
EUC5d4qZwbEZQ6elknSwHe+u1kRTYMLhKqZJR9eTGxqqV4/yAf7Yr+rBBiJsISBm
NIjh+QOcK5et1nQA52TzsQSXt3J8YILfg5C+Fyoc/EtcPOESkdTubjvz74aQ2rko
huMpkjgsUbr8S1B/wGoPoyRSG+sbZ5MVomNoMGZLZ/2Im3uSE7uijk19V2FJojSF
nSOR5etyVotBLP73bRylNKzfP+AYfpWQHRYbws1zOTmVFUVHwMH9R/CDyiEcwfuP
lstxfunU+wkXD4MSazZQMNUROsq8dMjuSEpZK4t7FawUw0sULsZJZu9xTmabS8v9
paaScKBDHLOciqR5d6LWkEXkWdh9HmnM91+gPS0uqvtsmVE7RRS1JR8bTY1CQCZq
PLK69gpuHWiBcDwnjc+o3MnVV3yJnQYIlYTn6nujmf7r8x5yR/4dsfVmGZ9zlSTu
VpeWx+Bq6HpOAegS/fD55BRK1mzuMWnAB3yLID6zS6gpoJkNShqGEGn5hbnLgKFG
8+bWPHWT1x6sBlpTiBuspw==
`protect END_PROTECTED
