`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RVMKTjjQYNMgTraoMeAeQk/FkvzVswlm2f1kRb58aIn2wEYEx51RK6fSVrsbUVU8
9kn4i9p5NkfTrR8jiV6XOMfSfGz9Y6Gl4VcQETUe4crpXkSBZiljDUDTja7V5/34
3s2Sb52Br2QKFNU6RAqjBFxvWOACZ1csIsuvpy6guoimS6XaisK1hAVUluNTEAsF
v0qe1xfF3AR6ewtZN5vFAx2E808DTiAaUyzTkhLa86eN7TZU28ZacLabnl4fx2jz
17cLeHNTPysPrdqIUGm33WlHhsJjxxaeg4ZxGSrdJ4RYf+TOkG5SDQjfNP8nfU4S
dlnYfu99tghx/NIK49wpSIDj+2z57CBSX40upHfMl8gji+fn7nhgqiTzjQOklI81
VhbJUYOLJfVIJB1sQVHCl5BqYO0REsqKAjpQm5b9wKl7yntvSqTDQY6CemgDnfFI
oBXoUnLXjURhO6cHG7MY5qjsrG8XEJ/h/a1R6QRvDdAkgDK3jrPMH7n2R7ZfdQu8
jgb/OupI+AuFZyI9FHdgC/baoKYDps73MptBkaWkSb0/DRyVQBw5R3HYCg3lffbp
YFBAbzpYb49wqWkJ/3sca2IeTsDN8yjhA2hT69J8dMR+d5a0kXzZf6nphGsBqp7n
hMBrVf/O+/lxEZMBSivHmG1fvJ7QmDsTaj+pOHo2s8+386oDBJ5OUkaQqCJObXjj
ccJwedcfgZQhJkggZ9H1KCCswm5255k5BOqmUpEuBwE=
`protect END_PROTECTED
