`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+ywwp8AG/ZjMtpdxvukg5v4qQhpxw1Ib9KU7Iwk+2YFI1U3wE/t+G/iAednYVYtF
Y7xnij3JkPi8+Bqh7leAIWVGHDL2kplRzRYxhJjfo54MKwG0Ua8TrZ50D56g4c1d
dgKeBfYK8SEMzM2Y5ZkRlASgtIE57az2F4c3jknVIDZaG7usHr3L+AliAiiRjM8C
aNoLM/tTGbU0nTdtpj+jSVTRehVcrmP6bUzhj4YVDONrU4Tv7tvms4bzdoyKO8YE
5oC10ZYOFm2bcyfQB494El+33EXdoALVwYzQ+i4c4xsZ6HRElFQzEbIWvYUpamev
Z7ar6ft7/kYo1pW8rqnMFWJ7zUFZvv3/PmNd0yZJJyFZNUJA5r+0g/z28G0um8hS
SXEP95xon5iCFu+9ss4EcyxcKV5ocbVkX7KguNUjkHbLy+cWhoJ61bgsr7pSMjCA
VmZMaeW6/ctK7UcR1tO2bSgQaXdq6kwlgTrpSEeXYuOtH+bbGJRZvpi2xORkL61S
vCOBPHGCPUvcj3K3TG8g8gGh+UwScSVcHgvRZNxea7JHs0VrICWFBcSOXZhogLfo
`protect END_PROTECTED
