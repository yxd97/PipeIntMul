`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TFIe+RpuzMQRcueg6rdnaFsAc7OBYp8aw022O4Eqo0vPzeu/LYyJNFRTseGttuDK
4TslFYehpMMXZAl8S6ehYXBFhZZ/W+Icgjslhtv1LCRWjf1RqAqpwwGd/mVKnVux
4O2QbGZHZHCvulo9KKS2OvSpMD70YjF7ap0c+M2sWZyXe6ck1heqU66WA+tGGOW9
2yoTF5Jm/9H6nyRsK/LzXb/KxGFxUMiRCdlLVantrmJeBFdUIniDEWh36lRqza4g
ygMMUUMuu+1FGnWsHLSdYsks0xVxagRBIiquCIGXCgxig1CJw8wAwLcg+j6T5hEH
rYd7SFoO1KL3KFmEdH9wqpaCL4bGIRaLRjo5tANPd6hciUr0vVSqDeK/1FeCFdqm
AnpBEpmnwrQK0TaCjd5VCLbRH+LsFgviP6nir0NADTxfCMHetEb9ctTBH9hoxK+7
9NU7JSAiWsT3u33x8mFw+++c0PqVLbsJdFKXUwzHApJtQL5r6lQcSvKhKZA7qIRN
QVIalfTrDkzaRn4Jhc2GJQ3BYEETnOag4vJoNpWOVF7R3Xm098D661OvyxvPYaOT
wU5odB6pNz9xbM6fqhliy+WwnTZpX+rw6tPe0l5z3wIAyWu0N3E2xvGNA5c1HUa3
SiVLgZgnnrqqAeB7sGPg8RYtnoKEL/NdQqVVOnkga/DiWJxs3eEdgRLpMtGdVZi/
KUdTYC74v8TTsXOhCb4iKoPIwgJOMV+lEoUF2lwLF/J8vySYqTnQT96+tGiyBo6J
2Xx2K4s24OJf1rfxD/tynWgaIYtHYFAVOTpXA/TlGAJpEFDj0KfQMT/RxjdeSyrW
OtwWESbtzzGVlJjHidz2Ehg0P/NfK6BpV/w992TTKdMDpYllWbnUeqnbnEgFk45A
xry2bg1evhpy8LQPgaVIOA==
`protect END_PROTECTED
