`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ts9YwOa6VVlU+PT+G3egbDKJhs+mAwyXXNfTFij9AikIA3YHQhxxaOU/1wy38ia1
ck2eU+z0Xu7Qx0Zdk3U/P4CVNXVABGEhTM/JFeaa1sNc2t8NUHdK6baZPO3EeCYO
6qlZop6JbVD8fidGKVJORyIU3IX3ykuiufjhInVDYT4a4ycQV1q6gmTtGqLmN1zS
yFaHeBdMLU7Pmq9OICpZhA3suU1rBvgX1rHjTGEvjwsuDUAzQe+FHiOE3fcdVYAJ
RbL5HLit36Jv/hGOWuLz6OQFmRilKObZJrxyBr3aArgaB+VvTvmMFSc1VGRtjh6t
r8RaojbiQZVUhZqpAkLKXlqvXZMbm2/mTDxuwun2gc65Rd/+TeYkt0cSLkhCaHFT
eJkOMCdDvQXMFvjcseJTnWolrX34x2ExWpilnIwrsLBE1LPqkLFFWKz8JyyWGZXo
R1YvwV+6vNatQ2ILhkA9wt7u1hdKU61PclIRBX8o1KgMud5wA7fNugZYuOGowhFx
sxdDh8VN0syo62MERoJsYLESuxRACxiH90Vn+8x4dER9sBysNn6eDdfWS2PoTRvc
CSp5qdmsyKKIyK2Yd14j+r2IH9zrGloVLpBFN+F+FtFlnz3NkeGoKEz5yL9xJdmt
GaJ2+2RU6Ri+KRJPk9fIwzATL0uv/yLbvIOa/qVaZ0O1mpZ1DHvHa0aDhyUIcWtu
4dMbGaLYkn8+8PoPm4FinCbYxf7axYmjxWpbcnS+Ila7gDclOwlUtHdgq5UiInJm
lqs7RG8T8ViVdbyk+bY6dnqz7GfpgVcE5tfS0o/GzXgvaCWFYs8FlYKXtaHxRtC/
9t1JcCALbjvQdJieSbwYZNNPMDvefImcdcUveQXhKpHa7p3eDQR2Klc2UotuhKHF
SGsDe8sOnr4UHMlXu3oM7A/Ld12udeEC4yW9D6UCzHwJutBkjNu8ZhYMw+mn6HGE
`protect END_PROTECTED
