`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4pXJNcnj0q2SnouvYPiBDb1RbDZwAcRxYoAaeAHmwPb5LGmPpE6D6RNG4BSZ3QvE
kgBdWHFZJLKRfPYJ+8o4w/8ObQSY7xLzRAIA/W5fJTfwHL67hngSkQb4QnpQWNdI
Viqu7vJEMXKX1F7GIGtYb10Puf6imE+bx3IPeFEwnBCB0iS69/RFQNZ6Vh9UG3/P
2s9JJ18o2oVuSatU+u4ThPuwLIPaqORV8D6Ced9LZrEeBXayU3NVk5PybtnlTcnV
+NcK1UpT3yMJEwgBnytNyfY/UwabLzM8xAOJfmhZyQHrSjJJDe2/iXkj2QP01o/4
S5CaVVDUIfZLmXCw4U3ob2jWtiEXDNq9/+bAwk8xqglatbIkvCPyezMakswmkdDf
FgEF5jV6XTTRcoKbriHcMyIz63iJNNVJzwqtZnjwc2dUOFnDTzkNI0v4CYr2ea9N
t7BN4vBVxwP9yFQLOUe+e/0Tn3V986t3Lh4NXJY3n90wWqoE+kwcTxuk8CnDv99M
mMJ/hmY9Oo9NtwirQPk8fGS4XgFS8rWTe4feYYQmi3UzVPo1hvmJTxH6QLt5vkdi
wbb2y1vvigCK1Gm55LNoMVhnly/fai9LSQT0xiD4+GM=
`protect END_PROTECTED
