`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dA8wwflN9IXJvKsiI51NXJHp/iMrlv3QNSpArnavmbqZcEKHcx6yqZl3CFu9usza
+DtDab6cRCZReH+4nKI7ntw3TmKRUcfNun3tIAbr3OR18eG/KST0NVjlBcLiQUHl
81FRnDDL19ESbbQo+QC1eIWvaPVpKox+UFmGLGeBC0aFwVkyF9FPuQ4ytAWKhEoD
i+Zw1B+3YI0+/iYlfkPNYApG8Zsl3RQqBCWzQxRCZLOLSdoNdwrqZjVMuMQ567ah
qedbNPOiuD/znpgf2QuAAczaoUvftWGiWRbNWx+tFGKV82bjbZOVBWOn1BauLPjC
LMg4aHu8GXKRlNg57BrDcQ==
`protect END_PROTECTED
