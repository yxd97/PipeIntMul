`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8ugl7VgySzItNRP1AwfSeENZqot4orhrVkwoW3apMBV7LBRMWrhTqRA2Rg5rEgiQ
6pjL1QCL6EMqb6motOuuE35YYIy5gyq0lyuAzQDgRmtFCBh2DCC+la9HI7YBiQK2
NZNpgV2eXM5nFRxkWJjtFkcg0h5IZkYaLWN7VAp1q8H0c8ei5jTRSLxgttbmJvTT
NtSWUkXoI2PJY1KlGNJG6GdiB/OPQYAquWjGzcKNtyAAdvnd/ARWO2gKIM5bpsC1
TCu241bT60QNpr0O9PjExkq9+cblVljKBlMq5v5tYFZnhV0O3PCGKhZL7KThVr8D
jHzVpvmLNpoBg5+5hK91roGvimtvYHZ8lLxGuWna70Lw3pmipOwMchOajkdnzfrg
pjnf9EcqSzKh5pl4dqoQjvkB6RZg4hF9QG5vQhm2wDMhWu2guFGJKp48WJ1qqcRo
TNy/OXZW5IKKJbNilyeXoVKvygjGZ1yrPjXD77SPfmAtA1E0Jj9f4E33c03GM0QJ
uIuySzSjGXCnObbPhtR9l7K8ywaKL4XXLOzikOirH/wcZjRbQ1ARcpeRN14UG2M9
Nw7bll8/zAD83VdtOaI+/lctWH+RN++MPfEXZxFfotsfHZj/DrcwIkNgBiy8t799
GGnUsX4AnhCqos4gyoDVVeBetfoJzuxsQ2eJJiN52a7/X/zLLjWtHbZch7OgLAY8
/Ej4aDNUZn5qgoKeLd48kX4rVXMQr8ZJcWVuc4fvWIohsAOklNC3vjn+R7+b8sFU
MZrdvaX9L0acgXS7VOLml9z9LGfLArvVtGkx1yu3W2b/cZJnQt6ZJy0lr2eSHEQ2
Da1kwTWbwUrXWhI0ANseNG/4ZkovAYPIiRcxbRpIFbMVRg7jj9W9gxI4THnFtRVN
c8XK7e9iZjkuRqHuTW+GCDUBgvr6Apm9fPetd44Z7oHfYwXl6skqP2xFVUZG5Wac
m7BFCOWDdoia6ZLAZRQi+1V7zsUjFE6kK/3SeWSLrTftTB3WlXGFmWmjEyQeJBza
u1AQUH0DiA7B4QQFSFg4Rrd/uFE4dLal6JEiRnFn9gAckjOEa8AdZGpOBVRXIwji
ujRgFUS+bYWvLCJRFggEXA/UHPVy428A57ADhwZQ7ek/Z/fa2Hqpwnzfx3lJutwM
uakretukBSO3c9Totcavt0cfsS9chZDLbp8FJQy62FKYr0HrI0ZuitNnH1AFr5V2
OipbeIQjrmJ+x04D6plFLJUu2CUfmPfzv+yEG++mdENByZ+f8rzgv4rfvjPRmEUl
pP3/TiGHQyXqqZuAxpFHdAfFzK4xaKDNfoKpjVdmtopBwJr6tQxCp/w+PEfg2pB8
d4T3UnKrL3shm3BVG4XpKylQTsfy/VhO6NDsaR0Mwyr0NmdXTA4jseyoAVpB6eOS
iM9+f9RlJRShz2OZfxWPxEESLzxCdViQY5gwiigOvw9HfCXdT7Ola5hzGA+pvtdI
lnlXQ/ycQ4feukPBgVgq0F07IqDWdHzjOW9AV1zqunmKxlGdb2k2pFYrU9kn19Bs
yth3smQLug2h3Zwv4B3Y/PhgWoQrPTvk3fqAKoLWV+rB6AS/PSHy2rY30cFCxffv
rWW6L07+EcT3v7jfE5zwkzqVpYgygIw7m/UtuFx2z/ytd7y112MimJwk4c5fhkIq
ONp1Pkjoz4Fbi1SDD8/g60TYLlz3na7J5lDMxCoIpOoy4WBkVz8weKIzAgfBVGAp
TdRX+oT1WJQfrgvS0jcYIR1/Gz9S/2aJN/tWDoLjpfbqkTIRE+DkCkkf8s86Rxy8
+D38MpzjC4+VJLXJQn3J53J5oNyMZg9rAmEmWYdtODpUcwlMjfCmOmJnod4FdU51
xts1yQqarTu/2tbiXsO+QOaTkHceyC7pd68gX1Fqn/mnTTLfB+L/gMKHlGurrZKI
U65PAvVVX2hLytHwktCsIammPlUKw2iPiXw+BBHoOhcV1/RQx5fBzd9jM4DgBLMZ
K7utQLWLCcHCHa76WddCPEWk6j7Yo9rk2XhqSM7T+s+wfYlj3hUUGSBqLgFcabPc
k1TtYt2JxaSWbu62zI1NpF2TZsx7epY3xht22vkbME4L1qVyLIqORgsuQ31YQpnI
KQeZzyfZOmcP/Yi38TCM0gLe7KCaj3ggSQgVsKTgIk+j571vxKCfSeZanp7znaV/
LN/5HR1Jv5ozggyes51RuYF+UsgO3AcjwsB8riw6jRtfQpUzb0DNP1t6gymVPZC3
6+fTpMO0rGz9ROs0ji1Ln2Vglim1OJW01EpI4vlhdctS8+NtttYo1L+rtWoCc2BJ
eOkZmVCiXVLauimAruBgQI4+j5EW4b1GecYaO075yD0PwDT+YFfV9xOACvgDcH0B
YiJJ8ZU55YTd+NYdZp2c/0FmkOXNsA3HOcvEL1oqhCBgXZjeTrHuUkccBl/HtO2k
9fHR25Zh1/RUq0GM8nA3eUSLwgP8x8d770BJQzeh3eG3zzoioSAotLW1PlyuMany
QDTONCRqxTvP40U5Xc7MlFZcKRHSF2NDBZobX5wF4RJh3gU8E7U4lPTwNPR/sjP/
JBfzE4uspqquiFJHdUeL+YeW0SbnQYdt0ltWlNNLZ0xSNjFdM5jhP3xkjA7VJ0n9
7gVBAcHYxWk+4e7YaLCWa/GFz2uGkSrkIaphOthG5lZVxHISQLqBzLrBzfSRwfXF
jNAjktsBbUWSr9T4mGtftVjlIryLyNDzNplWBz83YOZhBu0YGhbSUBT38398khNG
WQaqj4QC1jRSA+jAdxetxRqR6WjP4ygMh8rWQI3yLhCx2ySb8P1SxF0SzpShXndT
0MfRjD4JjB9DXdIWVoJKmpk71fHUO+zlTKmAzj0nm2zQmq/UM3vqt4+zK7l3dW8J
RfADGERCpe2KFul5WN5RPHlVkur2XhvsYa2nnGo1kYy4v7O/eNQL0rMptt+bjtXO
7wo4uZrHY5whybP1+Je9GCxvwfWRxiis/375rcF6eJGuqOceIrJRcLKS3b0/GAG1
bR8a7x0QxBgF3CkL4S+f6BVeyxmSbxCuHG6vlywG2a/kQUMNYdmQJKKYS0SNH7On
aNAZJpFlYH4apJkEYkq1wdBn409gzeWaQRQjxg6dFjoXiSlneoQkUYoa/VqvLNhF
eE8+BQNbwiK7msdobxgndtyk05IgvCuU5aRNkBD6n34US9+ej+zeSUbwvI2IJ586
qysdQ5TxH8XfnZYDYF5n3K2D9HhF8V75d1AmzGu93X5GiiYktF6i4338PbpjaVfB
t1P9/gB+y5aMfVPr3KMSRY9OpdydwY2r+PJrdWdlOgii32X2wjzY94FDSEW9NX21
kjJSC0n+i4zQAO8xeAiXap0Ox87FczrGHMgt0t6duueX7w3jaUy60fdRrTtJVTXq
Wf4+Zp5rrLsJOC6JI7VkAliUHggK6UPt+eWwQ46KUCLWh5qJS6LcNs1MZIsEhkLS
erq/pcDbxyspYsOkodxfikJYpvQFz2JYCTQ5MO68pcf2qdQvICkT6v5b1w4wLo1M
VYvaqsMGuohHJA39DK+yC0QtCNurlszClE5Rnmh0OrY=
`protect END_PROTECTED
