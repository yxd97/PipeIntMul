`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xniXFuqq+YRnrT07aoqxUCbZg7ETa0dhZvtteJgysC671MqnbPrwfGDAEvJAo2o0
MQoDYkRyZKEbHq/Z93vPtYnee8IbSm2Y+5YbENdttOdfgPHF2H8cOllOCl9sRfPd
ftqZbDqCSW2T6SNYH1P9esNgdNmtHQqxx/4jIxrtXIb+Lrw/31vacKy6p/MUCVUV
oyiH5zdLMSoa+E+OaZsAvYdeq0W7b7dNiCcJT+4VLPX6UGlkexqLpcWCJx6toYtM
ql/ecbXZN3cIyvEn2tVCHn85KcIZfzo+/R0hDgmUpFXT+RadZSWdmWIovsN8hbYE
4rHkfeLPORYD6ySEevvMrCx7ng1xvqzg57/z80BJHeuWqG5/t/bkJNwpG4uKwl/B
q5hMIPtMg+CpHBdmc6bhLWb2C9lAvxsCimYr0//3AkNq7gWvxVaY0CKPYt3MArfP
ODdMs1cbb8wXPd8QDo5dAMDVRzv+hvlx0kFcHms/dhurT391QBg2cWIHEgA9dGfp
3+FIsS8muMEsJg6gq5HyPZxjjtvncxwnoWsEvRaiTbKO7uHNnkhr/3OxVQkFb30Y
OYsgCVTEYRsreh4s1B9VOw==
`protect END_PROTECTED
