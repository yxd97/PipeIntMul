`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GLUxJrDk9D5eD0f2hwK5Z+ONKvlEpKk+QxRh9ufLLnCFm5xVio2ve09xb11f/Xs5
jCIPCswmeRMIsENCQz0x6rILF5Y1ZbsUAcPMdn8HjHjbSJWQagTBTD4wbfRwK53r
PSH1bBBqjmHIzbIcdExDuDlV4rrMUW25AQKZ4xgLQduLwhEGbnhZ1/cnOo3oExWx
QJG1BqSbmW+zueVe2VFmbpNjNOoTyIOZsFvOKOlBhvuQhagyloSxUgmDglebPEiO
VfnbjkZbFqSLKUN/OgwpaPYwXvEXUItbkAYkpR5AptTHIhVtfRLoLSV1CCZaaLIR
IKofS4//VzUNH98zLJ+Hqw2XapTBGrowGFAhWwxN6mUnZRvhTc+LqRqcZfA3eDJ+
SeTWeheVgKv1VbUUbmDNviXX7cFSoFra4d6vzff75Aws6EJIXSgDIcXNVjIJoxyU
`protect END_PROTECTED
