`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xRx529AKDazCLNvi13v0QLApA8BWL/n+ZOidsJ0/6iZfElwFd4Y4bBXRv51zUKoV
09LcmfkW1SUx9591VSW8XrhSDDfIAC7oW3IQcwugLHGU5VCJm1cHBGxE5pWB1qx8
ZgwFD7sWFgwANrVMf7BL0Q1872Wm8FGeJhDxGp0qqiw0kymFKHWVImuxSKu/GuGe
74b0zLNmLWawZjYIaA/emD0UJLAwVYjg3oNQD/HcQEtUtxt5wlqrbH44CkzEmA3f
nSgIb8y6eIqLe2jZlvXomc8jHJv9ZdQz6sLm8GW4OL49F67D0nTJjCC1ZCFw9M3K
gmf+gkMO9GgEsr7JMb+Qd8nUCTWgDFtE1P7QvdwzdF0lCfOYPzQ+Ptk6aFNr00oB
8q73g8VBFSd5GkFF64AjnOPBMUsi/We97k/YkfjcM/AhcWVBdPy2KPNTarrqoQHg
`protect END_PROTECTED
