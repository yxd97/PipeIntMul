`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
13qO9wE+S2eZldX5eX6kC5oUkLHhCJnVOCgh6tBFiceDafyfBTNRfnETME/yFBwk
hkcicwf56pTBkk4frw38HFVOldk3tIQMU4tD+ka1sr+jhUA0leZ599hmHohCmtjG
rRP8PNG73HCZ9UT4COy5N2YDr6Jo070bmghLfPINyQ/wZsuJxuCVV107UAfrBW3C
wj4qFOdPJUZYJc7d8TuGviCNEP92c9PUEw1ukDnodM1iuI1RB7gTme9VuH1HgUTl
UJ7T7tQxculQIJ9/hW38xT78JDKFV5OZ8d5bQA4x/a44lcltMc8wKKkh6/7p+n6s
`protect END_PROTECTED
