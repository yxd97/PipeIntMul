`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ST+GA5tbY6VuhyNkDIuVMft4W0GGTKSi2WSWG1GmS2uWrGJU9y1nFDCsyZitksLl
3X2SHAnDv5pmX6HZTIYvrQaXnICZEq3wiPtu08TgcARjXm2OsCWf6B9lekKEXKWT
FntHIffqbckyD9P1QzSk0riOe04gjRR1hQcKuYdR7QHxeS9FU+A5qkIqVf4VgpKp
iECrFYrgrtLAMAJ6vrc9b7QG1TmI1ivo1Q8X9zDjeOgbuS2mFPncIJNom8ZKsJgP
1noYtn+RYoHVM4W9PnAhHwhDLAWpSCo4yIM+26JUqdQ2WzXTlYLZsltsjxzSwBZH
qxIHjfpVAxNDqMmdlxFg3zf8tMJEAUGDmn2mfWdHe5SwZeZylh3GyfWOxjWNPuXd
tr9UGCrijzm/I9iCbiRyAkMrtWye82ttGrYNWjqG0sIZGSp1QdrF/nPTMAeY/0uW
6WqoCt1Ech4tzgFyWLaAhEM7FPyNotVv8x3QKPHJPn0LuwC7Aou5b50xiLJIJbjF
xVDh3y0geypCyzenz0DhuG2aP+FhM7pIUuMPK/V5vpphi4+lFZCOa8cg1A/PxOas
Af1jQBh94BoOjFz9X9l0Y+QJjeTNWFiO/7pX4uGy2FiaF0qWEhCKCE1P3rTTjp/4
JGyaoPbw4ebUSdWmVlSuBiABk5xOp3upSL2+MjCFAuJKZQ1SwU2Sg+ghzSYYiVJT
WGqqF1oFS00mK2dI/iNMrHGlgm9Kb7L8SmQNUX8QfBx3gvxqhHj3m3yHBlIXV9kd
PSPIjcoCfj3dlQoFdTrEJEFjNoUHA1mce6UlqfhYH+i5KsnfSg/dydgFK5g48a2I
7HVhMYM08kAAvUtXZVV+jAsXB0z3gY7cdTAPBY/q0IOGgIEIv5k+oD5t7JQC88Gd
nZbsXtmJlJUXdGsNuVj2QK1Z2yTf8pR+HUWYxawo+Ny9b5odxvQ84ah4N2xPGfmh
2qt4z7F6oayxERoPccReZ7wpDppN0AonCSupVQOY5ehURxRAXuwlIxE7OYfCLuls
BayreIoF4U5Zu5qDslz/MeBTFMasaMVkONRgFBMgHxA=
`protect END_PROTECTED
