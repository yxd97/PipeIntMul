`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tOc3XK4uX2IOQj6Y1r5pt0Et8lz3SOOeADrlFRH8WNgtD7xFMuabDrRx73CKWvxw
xFgDBV96cNKQCtkzYB9tVe0RJcOyjvdPj5h+lCqecz81YecYQ5swh9P3JgWFRh5S
mGNKWZkv2OuBwbyKo7UH/85crsGwrOoI7Os/+O+hX6tzTkisCgxcWvuUitZ0qCxB
VIZjXsxH4aXGHNFwLkvA8KL1gY4Ju7ZSkm6RlvkFHe0c1pv3st4JJMDbwlOG+JIi
pk3izsNNOR2XCPl63kZxDrmvChBDb1E7lYFihX9vVYcVihVdJrZeJoGdD1QhvYvS
yk8xQzM18ScYGc5YBtxAc2SZL8ZqagcDW0uU8CREi341n8sFPAyW3tdlxcONvvEL
AKSuos2ADksGjqYGKFpHfvo030yuzI4p6DL2lDP6zPLTRJGYMLZpHs6pW+rzgWM+
wYE+Fxh5tsnuzpOz20zfy9i8X8bmZlxKw8j8ykeo1uYU2l9eu16aD+sLxFvS0BFe
1oxHdper3rm6lXiMK/xaHYuLAvTbGrtilqaUN+XG1Y5TqbwHSA1fRN30SUNGRida
j3noH5A0RZByyzBvs/F2Oz4D25jUPSK/+sWopf79GV743yWyzWx2+CnMylyyVs+e
4qfb+ONPlxKBnWYfjaErxLy6R8nb+YiSrzjEx8o29jRZK9zpqTcmG1TmMzzD/h3y
N9pqi7ibohE2APwrH36fTUkS3GuBPwJ6OwoWFu6n0Xva0u8OnqSqw0HnNXsELdX2
mkaRE3vUSXMVeaW3uykdPa/DhPo+oAGpZVr9uhjoemSalrV73I0QL+GlROcNSYms
9WuW9BI/HGXp3+QUvRW+Daos90yh22HsdH1CsVsaGfR+VrYTPHgGoMKJTYU1fmvF
EN6ZGXJwQfITgzgDlOZxxx2VcWffxcg/zrVFM1f1BGoUtUSyKc8uOPWPtR/WTyk6
d5XjHT54AgysrziPbVlMEk1dPoxmBkUnLpR18Ac3Yx+LLw4XML2Ymozb2HeUa1Yp
Yyd06lR4fkSZRAxsxtHGTaZKX8SAcGpVC+cBF+MIeLanpvaoTjDNADqggwqKf9vM
W2wE2jo+1sN9o9A81qMEQPifIEyG6AboqKVaJBxnJydp6ctIVoYKKjsrQ3+oa0hu
XYg89dgdUP678CiAbkqPrBbTYKeMFeK1wHAK59qM3lEG2jCcdX9ssX2c4F5ugTHk
gQy0cMt5maQXCg+6nczejGPc1hz1Llwt+ck8LKSEkv+D+EWuoWl/REUTbmgdZfWd
ximCM+liT487b4SeoGrX6sC3dXFZQcrJmGgiDivtQwQOdH13KPq/pvpGO9f2GiBZ
emfTF42PLCPfMjfakzToBFWrL97PC/pw+ONKhBTRkg48sUZ2Rq77rlQybDkRUguK
/3a0XMNLm1YjtVCrP78eHe9xV07C982woNDA+FIyfAgnPs9IFG14qIH4t05YWI6K
KkvjwHHhsf4XOzthw+nIvvTQtdbLaU6Fclg0HZpu/ngSLRPAvMEy7lRlTUTePjsU
OZj7Hlih1UU+zRvzdxgs++kVG1BCS9oxdWxIOzs/Trm+pbXNU1P3EEf8c/fyD2GJ
ROgRgJ0Ws/jTAoQ2oSed5eVRNXTYaQj1YrUSVSMTduH9Lhw9b6wQH8ddHh0nX66V
sPds6to0u7BUqXFZe1CRQRsC+nuhi0Y7aOUi6JuQXegvi7dJvyvcuV6qHtpDS3PS
WULNaWrqGkIvR8X4F0RCJfHDZD4AW5wxhcivuT7EcinDL4H5injiFII5pUvPapEA
bvtfq0+6qoKqgEMd+m2W5sB52O6JRmOqxjgYhBMErVlXvGSV/6hgvtT109fIb87a
/5VXBUaO8lz1JHnHFz+Nf2NS5/IAgCV6BlZ70Cb8Dw61BSzHBYwj74FBfXsJSiqB
3ccC56FoXXTrJNSsMPCtggaZA+V52DH/2iunrJiQcAcZPz3zsnC5eeMZQMMWBO1U
AJa8LSrHNjtIn+m1c/y3ookbAiefWsGNy8li6Am2JNg8blhAHfd5zlE5xNGULhKu
M93FliCC7G2hld5A9oFkkF7aSfO97vFG7+9YUEz/KjKGiaRg8cKG3/X5NRocE3je
fUsZWLSM+qkvtXj69j/k+4mPtzHHAf4ZzBrvgUUqErDrWoduJATNbyRH6Gt/WVB6
+4EfZN7kGAPXFJLHSXDePjxJ7muXFDnVA38HVZBzBk68zXaOHFMAXklyTgFOaTKS
jE+V98o7BMrlAYzrtlPdtfEdYqu7npcRogdYYa5xlghohSwsuSCqgdQlsVIT4DIF
JnJZoxN15oTSu03fSbefcCbmnQxuPvq8JdPhNrtFlfAKJUIfSMiTYUFd7HHT0rid
Lf7G0uqtvviXfKiCfXio4C5sJc9sWw6jqqUAOJUUZ2g3bdXouGBsOomeBvWyBXOB
o5CpyhucqC1n+iUtpvmh7esfXwDVINmFd36U6A6vARd6qsuh5JCBx5ixFl60uG1j
8LetpldY+i78KA7PNp4MuUa25243KfmTK6eOMtdCCprLan73Wh61zW4GbnfwURZ2
Or8xPjQLcear1UFoiume/ttBPVFiovj+u6i8kgKbr9XJrRQuUYtFJoaX4FF4I721
wE/7gDGUCBjMKTAZoyZBob5wuLuqeMwuuMQVNzeUd+mZCzEJuYoddRdhYb5VAfXR
SgW1Oaff30YnZ+UzdGMTVjq+TI7vW/TPUmMU3WKP+HvVxX7UKRZluAl0A1EM0MIJ
oRVfcxf8PD2MS2Yjul2I02z1xC5iBbl628tHUwvCSm90wMOXqMXOg6aLlHvrdNOV
aY2hHZKOAvnnrgMknfjRUrQUOxamAYuS6A0gZdGji+GoSH5sLjN3iRpj3mjtcE5E
e+WhFA4abagKQEadiz6s/VkTdOgDEtqXrqHDSOnkoKIkDIkYDDzs/DP4rpjMLaV7
pCgktz7aWYa7LV4zzk2bB3ZuiGu0aTyuYSGJb8+rtDPhaRQIthODmOI6+iOjhts9
jMPdB/pOYjWc8Pm93uOTP6NvGhnuCTuSehn4XKq6JMDSkE+v6KRlHCeSSUweetno
dEzX6Ie8OQQtziHQG5DaWhxE9YyOOeKdrA5tiAq0wSpr7zihbSOkbcgUP0qEr2nH
mV7SGC4T9WgWIIGUvY387d8FbvB5wDmMFl8o8PTWmDDSw3+bnJtSC52dRHbjSl3P
V/+6/mMLe0CCEieCuRNub0qYmwJXQx8gdvHjMUzQcPnrlxx98uJlV7NiDokw4UDl
I/EehFb9ljCzcA1WNH6PdBU9/kGqzIRwzyS2LbM5k2OMp8pdXRbjhqVY+4ciffiA
GoOwKfvrGjlJg0/hzgDwba5ckluTD1jzWVyql4NMK/COicSfeuTdXXGBVwWNwc3e
z/DhpSHOBXDS7XeM6ZPCm8E6Ovp1AFrdowP8zFl2HC/fGMf5JNNwC668/iBZi9DE
YF0azELlAhYczvNJ1TgrVFqIS1r0v7RlqGuOgHH5xzQ=
`protect END_PROTECTED
