`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1TmthuFM0plbbKQiU8TK+Et4L5t7irwzPOZ8eEfMpNK4opGfqEmNvGFCBjmx5rqV
VQ1ivIyMvj+WrjaSyamgiEsVLJHPysCpPOgqbKNzYSWvheD18588aL55AKdD9LGc
mdddlR0Cebqaea0oaPccwi4XtxLqC435liXbzRJ7F7X/f9RZs4sXCLDRLm81mTkN
EEb6SHHc5pHGUCUxIi4qbZ8GEHpg75HzI+ut00HnjWfRfUvvxC7QUgZbb6ncC6Zr
Ubm2JVV8Y50LGMYn4ekKjgGiC72GrDjdevb2DUKg15bUo9cLvzsep0KNhkDNPs0W
snQN5cLxXjmzFpYvoyK7PwQU9VNYpkIIqW1CXCRNJLy+5CdacJC0IxMHcgL0nmCB
gTK/0U88mfKObALxUV+xsRsxknnrlssq7c2mjSR358rOIlK/d8TfLVtaqXZ5vNje
Bwh45zFZM/O7P0OrLi2lLouXqUEJKe3AMYZyCR/Wko2UXF81OztiCLM/AYjzTjY7
dz5+G2IgtUQVURLIkPb1OxyJO8+Q9ZJEzqAP4+MWlLTtMUXRRynPy2WJN1XfsQLz
PW2tDpkRtxbeWwcU0GOlQs41ApNmBLbhMWrMlBhWp4E87ra3W6jFhGnUsT6e6V3u
IHHYexZ9vhn7MvuPjEQeNUelf7OKujVR6dYn5gREqrvr6HVkgUsK00QwJkdXEPi3
KkJQdiq7EC+Ihv0jCM+k01diiXJoR7Hm2T4jQWvG2zwvekWdYB243WUrI1RvzT3Q
mfvoobuqEPWW8jgHC0K3xu2NRPGcbJkOSx//xCMqv73HBMLQOFarn6NABU4q1TmB
`protect END_PROTECTED
