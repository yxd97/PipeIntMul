`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
U2GYI/EXoTaahJ/zI3/wfeAmYqufOCXEmt+G3iZ+CpYM+GhqwKqbX6GrzRbwP4zj
dFvAwF+cy3rHz+SWZhGkGgp73e92Tf0Tbo023qrftPpeHWRjZUW16iW2/rOyfHWi
4eizl62q8kNvJzaOGQxLohZWls9glKJLXW8gzkWBy0AjuSAwaur/668DFIUX3ZGm
5LKqIjRXU6dsMg1HYaykC6IfM3/LE51ndONNiIWQx1WOo8Y+1Hw5HfdCKbopgjxH
7i9KeemiROEhfDqAHpOpxcUPgMp3EMETjnEUP3fLzmk5Hr5h7Dkruy1nbpe2p7f1
qmMRc95GaRLmBrRa3N86aw==
`protect END_PROTECTED
