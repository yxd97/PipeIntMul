`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
u3KnxdS9p0p83otYzO7V4w4j+jMzbi+bCZhssfpPECk8z4qdu+vROqn7PPu0JrJk
2U1Aodt0aoOqKo4zAZF+MvCZ2fitTyJ85EJISnoekf8LxqrgNFD1mg9JYfcPbIEh
eFCd1ZINtE+LBTvzyPy7xMs+2zU+QKs5FBkTEKpYrEzh/cs2LZRkv6FEymJ3nhGs
SS3hJj1LJzmaLc8vbJn3Oeo+TotoPvUubqXfjvh2H0Ay+CoMjUSgHA8gslzyQOWV
4+pvzTxk6kUpC/7sH5rInIsm4rgNrqbJvy5EhbClrvoqp6mFUV+EYz8oWEwtuQxb
yg3ILpLeNlXOF1EtBh5t+oLrblRKAXT4XfyZP2NNMkVKDcAouSRxYMNzU/FXVbTV
`protect END_PROTECTED
