`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p+G3BzgriNBxcKfkGadgKOJuIKmCEHHmIVcAuT6b8chwJrEom/kqgSvBuDG3AJmz
lJDNoW0Xd5A2dG6b6WrZuntYx2E66biRK6C5nOYZLJruJkhecLGYtWbUEGk8d0HH
VsiZye0hkQ/YhU+V3WlP5Iq4B/o1NHWSvQLWu7mD8POxNzOj/vP/d+SzlAsNAqqv
5d7cBeaD8BB2GZV3uNj5xjXL3dB90CW9Wszc8NeZntDEvnQDckywKJ6HQYCZGiSc
oac3/hePIPGLKNaKjJ8bMcIlsDEDxKVZzDT6Zp7A2e88As8bQc9NGBToJCjtkzHu
v5ighsnWG8oht9y041wSu4cVGrm2w+xHUCNoQu7GzR3o2mYEcUF8GIPF5LgbYV7f
3dwE7h2iWf5v2Meh1PtRaouriTgmXwmzXELy5HiLmxw=
`protect END_PROTECTED
