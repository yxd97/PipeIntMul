`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MIUDKSA10tv5hHdPlct0uqGG1xYuvXNxZCdGMjHEvJHenkxWNeDmcGpz3+dAWYed
M8r/Ql2Qjs8U70D231elYYOjLVaMfY+8fQdvr9DT3Z8+k/6qHyvdUsvAebkN+1tz
ATFd6DUsiZk9i6Ro/V4RoMgopSAzzqitklqbXQ58im29XLEBUgIXap7td8FuTPhk
zye2wuf4sVRb1DQc/Yn5rTWCpu1bILCUO9dRpBd1P+ADO+X6uvgvv2aiZXITWZf5
y5QxmJu4ssmq0vIiycn8zfB8i3ZWPRBnRRIsdIO0PW5hjkB2hUUAdtz2x/N5FJYf
y4kkUlck5lk1RjQ5UAG2qkeW6c0PkS8H1VB3QQnVSlwyhdBgz1767g+FzPEUtVcC
IGr0I1kbE/KUiTrFbUGzcGbLKnROyOO1wHuxj8gW9ANhzFZrp0LbwacDleTSAjfi
`protect END_PROTECTED
