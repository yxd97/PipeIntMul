`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mIv7BViGY6CtYApPZCjHDJxhz2qv6RKYhowBbx/Mnbjj+opxCF3gcW8nnXQnyORQ
c54ks8f30SSWVZsMDFwvQ+4zM0UVmLzyl9mO+YoG2IdBSVbU2zWPpU83J6FqDExB
HjaLJlLmFkscwUGM4D8ggSX3q9uUeBIO8Y8UbOD4xLWsiwLLxQ7KteZeNeJV4ndg
StCtXUbl6IYw/cF1qhmnxIz3ZaPTmpMMR+pDbl3UFN1rlwnTeYkARO0WAEfqW3A5
TN4lWSLCWnZbG61Y2/p2/h/wKDTbbHpTbDoV6GCKixHvATPglnE4q++i9LKJkhiG
S70s8KVsLVewQPHRXt5uOTACrDYwPtnwVxJA4dboBUdxqwMhdU8QcAV+Ubh6wRIZ
yzuaYTyRa+KAoBaq5Nj0x6SCCNRXwp82LgXzzrWDPCZ/Elgm/4NzuO9qZo+/7DKa
8cdvlxLxLlwuoo5QmLuwJcZI3gVV9/69bZmZLN4cnKrCqjvF8Z9czu06Ou7yI8Vq
GDqBlzD9rPogZZyo03ky+esv11YjxkEnmeRnhnKRurOEbWCOlJ7FzAZfM7Dy6hX2
`protect END_PROTECTED
