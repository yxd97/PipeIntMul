`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
//qLRDS4cw147JVC6LePcPAjbCLppPQ9/Lgsz7DIZyeJtgbkGnb7BUoB6WgON5k9
RY8hmgfYtCIbY6kdr8vXi35XFy2oaDgPfRSX94Z2muSU+CuCYhuaY5tFvAegx8gi
+cLcRzg6uaLbldug70GA+u/dyCBGXUltNmHauldkcnKwn1FVVzXxerNoUi4M/6Sb
HZ/QmLbcCzX2XDSV88r/jqFKSZ6+6N1DYG3W3l39+LRSroDbFhZh04KT9g+WPdau
RQKmD0jcQ/a923wJsrcg8zX45FC0DQIjJJKGeDZMsRhMoJ9GKnNF3ijSAxFNRWtE
NohyCA+N3RTTRkGTl4CLIHgoHAHqWShs7BhjX1TiXBw3f3MPssCTQylGOCAJzPnP
auJv3ErcYSyViSttPEUwrvUswrVaKb8LTimDnNnJ6tXsqZfF9j8faefLIJrqzGeq
AAmAWvddvIb3tUHRpPeupueqqWfwPemo5D+PJhSGuBBR9ZqQvjIKr3Im/43vp9xv
`protect END_PROTECTED
