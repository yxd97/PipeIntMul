`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFqZL0ZoJ93JZCLbtGenDKyhd89x/O3EWRAsMr+YotbYkpL+aUR5d/8+X8I5Ganj
Hu58hJyWfnxoOM6lK9XUpQo/urbcEZND2jbyLHRQK3ta6neRHxhrOZeUsLfgRJNK
tqFfOWp9oclhWJEA+h2nlOx/ojfb2pk9STfvPktRc3jDTX7r0E1kXTYAu8sg4DG2
kABd/4Uc74Xhs2GeDsl/XTJY1DYNA9NqpLGrdml9xnJWBOf5NTnLtuXXwt3iurMv
n7VKR8Gr/sQDExdAK+CztH9gwi7EwJ8Ww7j6sSaRA2KjrR9FP9jXNZ4y0Fcwqcc4
vYXLOq8kCBcQcrx+LRneuil9iAokLQkMg+SnjoqR31s1UVs4Rd/a6RpkgC/CfzJf
GFaDLfvQVN/XLgTWNws4WwwDoYVJXtKTPgGW/ZtwAG1om18p1sHf+PZVcbf/bwyp
y+menvrVOg7EC7Troc5KPsw8czKKEqqZqfAunrEmbWU7gSMXB1GYk6xqPtlJt7gz
A+1/jyTgC+O9guWso3DoUhqTfFXmVptFceSJ3pN+x1zc1dO8+iM5yoFelAxCZkoX
rnOnrO46ZLoxkh90Z9FEblDjkWWWuk3grGbKt0vvitVdOoFKadYljM8agwBs7WE8
SHs9AgRNTRraXceft0AzhX3jy4HblDjJYQKul8laSRZi+1HyVVlZtTUZbAXcgj5m
ronlcXUvSpaMJvAoWq30mEgzs7+L80N0UccF8BzprYymc8q8xi3YBcIh2pWs+s4T
xGFd9HE731/BYUYRpOtO4ibWRo4IOBFgnpqIyx7YkTbXKT6HRUs/+t2dBq0t89AC
5d8+8dR3mEoiGXUGBgfQCAMHkm6ubmgAWQWwzpCUQ4LXeFqXa7ALQaWnmHB1e8A2
5fk9UHjQbIHv5CSOJhBmyKlUCCoPWf1PIhEo4cOCUvDe6HRvnhcHo6z6DVZv8Gs9
UKXcZmnEIrhgyG7iHMv9Pn39PHql2MWFHLC5Fn82Vb1kOF8F5qcH2RhDAlYYtSwL
MQvM6riNT8verFqmloBIQN6cKcgTStn2LvDHtmjpiuwkjAbcc/slVCdpUDyxGm2S
6d6ZA+XUG5YNX5cu65fAo/VwrDVwCyyPWTvnCuJ+nbQYKBeqKxH+JW+MbmJK1ihN
wrIpQaeOlZaOSWgdsKaTu4WcqDi47B/gdoGKb0W46S/bYzDZRgB+aJ2Avu/EtG0/
yDSVDfeEtB/kKvB4BWP3/Nm3T8oXkJu2wp2bRygEpXY92wHyUhiuu8XvR/Mmblaj
4YxYrqHDEfnKF5tlNiWzsCGL/n+fhjdzRIJmBQrTQ0sAJKi5vPUywUWgbkkt95fj
B3UulPyW0Iaggf4CYG+iPb4zCpLG6Y70I9Vhq4dOy6wQ0xC+nTz8kamtZPfBzj/j
YnDSxwVVzQzrCyXb0Uq560phR1w//VMGU1E1zupSwbA5y56zqSQAHWC77qlc4jl4
KD12h3EE6f3TGPYWQFYB6J5T3NGZWvF59JoOsR1GgofjIYDZr6zTX62L7D7IBz0R
kh3U5jtXSKwhsNlYGZJlfcM8GPh9mBusWynjKmeKhloacJP9HKCKDEYrFB0MW/ZT
lGe7N7+8VZc/DcqV5wrQX4l7KMUTlAo3grfdaENXkttFXSiKep1bcOc45OdkybaC
ESOD/kJxnzyca6RV3VhnwgxC20MTHRlEQUKQYXowEkY25BO0+I/r94l5569OhV1T
viNhGuu2QmYMKHIbHLZRDZ5Vv1vpf3HScwVrMfSZ8y7Xcug4holQevuZefYtr6xe
csLhkdqhlAkBYralceKiS2jn8PwgQnmyGnXhJtVerjPmOVD7cU7+cu3mvHc8x7CW
VqsFlJiM707wnFo7fLm1rrnotF3PgxJBVkFOXrGyY09hXcSgf7NEBzw4lVXsHPbi
ZrpDDiCfy+ceOPUAbP86sh58iADyBSl9htsEWd9TTya6niMZm//XX5w8xj+z5O+k
4aLXkNqhU+vP0IBx9dP8gnFvr5qV84Z5lg/vXKiT/5O1h6ZuXVD9kJ02lvjqZE47
hba2odB//iaPAoMdVmQlv0OcspsHILVcmJsF/haaFN/sfC+HfoLSwX1YpY2YapM7
OonjSzYrTBtp6xixd9y34o6kxJyV7CwceFqWqKQEqnFL5JTYseEoA0nBE8gn2lB+
i9yrf7AIICcJJEYvs9EnCAoM9q0gu5gjY2QNmxSQs4zwoQLeYX7oL6ZKPxBWxGQm
b4VhspriGksW47LbaSg4H+GZ+3yX0dEODDU/YpQo0ljQOzs7ZeI4LcLoWOlcmL+P
3VwTdoti0uC1oDYwskLzN9lNndN9PxAsm09uFQAGbCZVO84IX8709UK9KmTW/3lo
tJrCAbRfQZvM/UezDvRwZhPXijYZCV0Nks62rpe0+pdoKAEBAkTeeA/0LrpS1JEd
4s96kXFRGrN4CfiMUiUkIihlJS9nA3ECcI0RIxB18+ANlzqM4Dj9iqBATwXO+q/b
AGM6bJFFxxjZUm8J5YZZ5FeUkHtr8Q5fmbe1HwLhws8JJc5ugcT8fEafVcsz2y8X
IxGJWu41W6vMO6EaRj3emcxlxuDg9S8FRaqxGb+B9SJez8Zrct5Q3C6HotUa3fmN
XCPi4F2jrANn+3lJ8JBPr5CP0Z4mCAiaIomH6ZRJvwHuQkspk3EpeJu83JZIVU2p
VN2VLNNJXNMzYnSUORcRADiyy+z9fJSiSumY9K2VOkY=
`protect END_PROTECTED
