`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
P921FaYRncmCybuX72G1j9J+aCiNnMxI/3x7h94JgELIGL/s6QlEopt7rhb/ITIK
aDvB+MNP35TzPMT+Xu0+/Nj8phQKyn55oSgLsSF8SVFKRSU0vqIguUkDM3+x+4pT
OPtiwbnkSnNkpc87SB81hZdnKTYtTnvobG6XQFfS1qWqqGIW903wndglGmu37h0H
CXirkOIQlPC3H3kTd63brkqc3ZzWuxGj80zIREE0G4ukORBOxuKVrVhUd9LUfHF9
Ha/DQKHs1b0cBKE98Mn8jfCZebvVYViBOOxTCZlNUv1QT4fOf+bh2EXlQV3nofR8
ze1V7QImRz2QZFOO4MSXYA==
`protect END_PROTECTED
