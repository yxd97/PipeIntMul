`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
saHhJXtCRAkhWsOmfHZFsTftVLxaqyGZBUeUf/Y9BzkXaOox/+Xv+X547MvMAdJ5
ySJ28GPm5+uhl3cVHey1TwZNdup4Z/3RnbJi4F/N7m4oRwMuLSoyYOhk2dfKRfBe
akUkCupNQUI8ZPp75JhSjwDhVU2QEI2itaZBhU/9A8b/qIiavw46zP5p8TB+5o65
P8q+S5tAHippmdr54wf4puWm0E7GH5gUGpriq6U/cPa8j3a+REU6XSbwz7N1kcV3
YAl4oQ2dca4qW0aR9kbhzpq48BaSo2kQXFRhD7WLTWKrZsVx4i8qSVEgtuULx6bt
XJbj6jOpxFnetmk27oK+qaPi0bGc0h1fmEVGzSi1in4pKpw9aBmNOSdpPevX870e
HALJWin7dzAhzoQgLR/iDS06QDUTs6XAkg0VOEwNbX3r3um2CfmQTOhcRrXoy1vd
+1e64k9HvU/LBpEQ3gjreE4D9dYocfH/xt3iQLePDe7IyEaXYpjgVTDeIICQ3I7Q
e27ZqnujrOMazsypnwnTR5BoTAZ4ezmqJ5zAAGKd224haRf/lFzoXG9ZuXFaqM+q
FmqknjS481hAuODtV5BoEYknOaeh2MSaTiYXpEqzn1WstJRtzgx2Nk9ZYZ4TykNR
8aYGdqRkatHqNn1hMWzHDjmZ3sptiQh46+pbUgpZhFo=
`protect END_PROTECTED
