`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
39zNb9BRLCBEIXJim8Unzn4kpBS1ehxQNaoJbqjMXiWWP0Bvv8zkShEqnPnE6oBH
W3DTO6JAti4zdRgdZ30bs8yiTXUQwVmVO5sMK0ya0enVo8WpBO4qMamuuM6Uszee
Cas/eaTo95mViki2WWrkYkg0NA4ZqQS0n+kVrn4aNTUWO1v07YokXPe36zUMXW34
eoGdWhPvWrtOoPWJVx5syidDc6k/IeB4G31nRI/xQYZdKAkTVkOr74LVwxV/0npa
MjOQanwuiR7VqOtXiVgugcluFEqiyqfqtzSlC1FZI5nRLFwFTKpkJ9jwTTdVusdw
Cd07GscpVNZjK5ApcmtWNoFqP7JOtLgUW6aCYMMaNov6gpC2tALErUUiJH5SJBX8
noyQAExz/DeJALluH70VcaAMOqUV1n2PEblTRVhLq5IIbkaL4EyUChQjUs2Nq1Xq
`protect END_PROTECTED
