`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OSX76qqllzPNzXPOFUbxkRP2zccHQdp2ws+FRAFErwJij6YNfxcDZX/bUEX2QStZ
E3VL+8t2H6mYwvsttLfUWhYJsq7dsQo2ieNANOtp2oOVIEYK2ilyJCXL91fkL9JH
fzmaudPM9OR4MNlrlIM5IlwenEKQq/xS2vnqrBLzMdyD/nhdGuYXG1AU161RA8cr
j6o7Ry969hWsNQ7LGDR7ymnd3BFYyKmmKe4CoZAPd+xeD60Zb9XAYfGWV1Jo5hAq
SpG+WNqcI3g0KI+PmWKpEOxxShWfC+Qpm/H76ZWOXFqfqamIl9nfcu7VF9an1VSi
roMKkZR+ec5+GZhLkRVOngvqUDdK8uuNnkyuKKjNWXe1wS/ErYNAjz1Dbw0+sqpN
ABplla60njrRLXN3x0GVIib4UGUUTuiiXQnpmppWCKMfCcht14QfzS9xwEvhoxRT
nS+HfvhSfnL8SRiEtu50okFCUF0FT4JgENyHVXAm0+HLtbPIvNDQNANTDKo08fyd
3J4m2JGnGoyMOFbmQvAUi15pLXB7zAL6oD2k++3Akili6oiIn/an1PyZs3joGd0x
b5pwQvp+FbZ9/9kvFaFzKA==
`protect END_PROTECTED
