`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qExrCoOqNI0icYZuZhhOvm8T7cRflILKLijo7q4mLDR8Amz+JgyhZHb7ghtjxX3y
pEBB1xiMj07O3ELrOcsx6AMUyD+AEBtlW2JYKGL8htK4vlh7hKmRGwPWTi94iHud
jjJULvGlwqWVMze7+UyDbzs5FAMd6w2bUTOeFVYz0WhQc3/lAfJw873PUU+GfSpI
RdXyx2nwj5i/cJHv/SpOempvBKYVFuIiukiEVPsjrR1+/QPgT2ZkKrNR6xT9D3O2
kS29EGjy2zzRXY2Iny4W1V6bE3f2jknf/2ywQWkArRT4yi9Qa+WiyAK0SLlCQhJY
hp1S2eaHkK8yw6ciYQvfi1PVjo57nv9hR7+1tJ6HDiY04EqpOdrhG1Qz06Lp2l9s
V/niArHLTCz6SZJ02/dNeUF981Tdo3UxtVGHPpp7HB6zLn11y36bn9HXffJw8iQ7
mtMh+wX8U/1VsSd22K9/o1RvG2I3VLwINe731fGsFmvXvL+oxpIBH3gpbopO6ddd
wBGBHovBK0Qg+JuiZLHvv6/k8zr0Xy+sgTRO4uHRdTrEoTrOvrDKOTOFtKMNsRUi
UERCBeqNSP3AAALiVdvcY3LlXJJ9E9S+vvyZ0Aoz/JzcFvRMxoPYZTZT7iqa9n3k
4kzk5t6wygnQl5hk6jRAtfbqacjOqNrx1JmVyQv/hjIViKPIuYKmCmXAx3MWybqQ
aVpo1hEFqyfsmwk//DNnNw==
`protect END_PROTECTED
