`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UARih1BfOCqtnjjf6UU/n+Bd4Ge+CA8fr6L0EIHBWUW6raFv4uxAOTBpipm5wglG
/4Tic0rg05SJlkoRRwwIOx1phyasyFGqTDybXG+6gdxfh8sWP0iKhhUAF2Zn9UON
lDxxJmkyGr77xR/Njuq4O+9HHmwRtfqE0qNNY7nhbypWQYAcoqdKIaF8lPfAigAm
0g+YW6uKQUanCemhxYGYVd9kPrXLMRH0JXxuaOUlVeMsxGJiQuOceCQ4lZy8J9iQ
24zXsPA9N/zgxWN4fsuQpiTVM4c0h9ulmXbQ+1ddowE0fb5hh66qFhFIfPa9W8GZ
jTch1PGCTwTQcKbB7hfdkv09Mo/jpy3e2cRlcrSXuAxR11EiDuMZq108Pp9P/Ay8
Q3evOkkGnDgCX+1tkb+MSqs69Br8+DOZLKza9luc9mgn+tFGco+LVuEGd2UktsES
AZU4Z4tf5IsCxUiL+wHRzSx45X7FprjC1sz2VjTyp5mcILfBFgYjEsRNnplz1a9b
TWws6hR5d0lGFtjzmUmiKMVWPHEirPkZyVLRZkhLv3Au3OdAHC0nlphBmCFm/uKe
ClIH+xim452v4kvKY1mgWOGFENWrARKAmMhw3a+b49QhzyC5SCgYmHwkc6og+F1J
zgVAJXivC11+PRKyBfcheOGdchmTOwYZVKOSwIMt59qUSujy5ko6bfKgQuN/6m3U
HxmUAt9UTQ2b92BQtfLNtvAVCDsFiYXcm79mkFmgqlfe+TIMwQXpYb5OoCXUNA4i
FWijxiumXghPEAEF13m3tXCNEMIy+IObJBXd2jUCNeJ1Onz0wNG25lfAupppWF9P
QkXq34hwF2dnJZy7VU/+ngnmd/xh51Phu4MXB4UMFAY6W/dX7uKoeg29E/EdSEXR
rEGRaxeylpRqbv3/Cnd99+VW4U71oFhwjsIolzHj5aqHXez91FxYa2URGQJdMBR6
YFH18k2Ya3mmvOsypnVx3tOBuRwqEQbkcspQHaePCzSU0UcmiZeHV0bhL93y6NQW
Uymk/IhtqeX7kzrwtZ4Nk15Tkb7SBh06bOdw7YEwXDzNF6/YPkvjdvrznXQbF6Dc
66JMBxCdLVbB9olOS+NxYUfyEdH0UlFnuC07n45VEXQvGjNpkIh8kssMuizN4wXQ
8+Jr4kjN0QLFEAl93IDwyC0e7LUxYBLWN9NFrOzmWzVbSWQ4ebTzalzMggssaeHw
F+CSy4NzeISAUxD+V3lOGhxhL1Nh4QvnGzlXcNQHBJavzQyRSRoymb9FhaQe7ZaV
XOCq+NVxsf3NKgTNb5APUy8acPWxwdycHaQsZahbGz8PeIy6PxAnUVmNcf4/acXq
0Ck7EnCc3xBy5RmWjq5fEmd6M4c6viZkPh5KqG0D+/6BX14mk2r0FreAjpuZ5Y8I
I8mop8LcrwFH0oGIMjKxs1/MtBbK0f00Yxn2WMNJWzKVHVIP18et4N8HDx2USQy2
ybnT+DoabA/FoIYU1eIztUtLbbUc26etXb+jAVvE9MBPcmbiOe9aR9RwMYcYmJ2J
W+alkGZX4UpL3lkLliKS5PeR1p2d+n5pcsuQ8K1I7ruK02uJUWgrR2qrn6iMXihB
ws9cntzOcy2ET7pBZld7csoGXR9aTz+aYXzKyeGAQbLs82dUR9KKuWjL1jBxNq1Z
i4TUIlEJzV9CYrTA4J36R/57ohdTlyHgzalxJwtYiD7M+3syzdBX1SNCgJT1+nHB
k8oR/77f+2/CRUt+CI8kQifcsRM9ac4P+un+70mVrPK4IjsmqPGgjRiPBGATIJRl
gEwMeh7HsbpS9bK/K52B5H7ml7O6V68yIiwLImnrowG+g9eYlrvi1t+Y9/dH35kW
ds5HoosXnv5wRg+ENcDXi4OpfEnaYfKBSegGf89ksNTeWxawi52lvF/14//EzS8j
KHIlYXp/7EAio2L8p5feYw5Zd6kpyHZaeOnx1+1/rvo3mH5ga8vh/DiHXSG5Tgbj
r7ROhAXeFgHwTggzhRt+R6RY7rLMaY9AzLYu0KFe611crNwV5BJT6QEVrNhla8ct
ZuNM+dwTCvFCU+qDycDfLg5QLwyGRMxON8W0Vh6NaQOeJoJ2jKGhannEhCK63zMI
o5aKczzynYUemLL/bLdmKMnVn2MNXz5b0DTQFR7/pfIkqEJykS8/TTIIkIxhECDm
PGhxNb4V+G5R2S/UwiC/3LrRE5V2xxhOssuTE/i4fo5OAT+KFhV1iZ3CctHKf3fm
/KWMoq9qIqQizt/UHTHhPzd/svE0YtR1yHWh0MoxOoF4kctQkfTy8EOJ7FNCWZ26
13aQ1GOF7tzAj9/yqYLW5g==
`protect END_PROTECTED
