`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUtpYTrXahBfuQNTeCC//mgp2s50B9xXmyISC3hSyyXzyjfhic38sDsxfXlzTsIp
g4iqKsQ1G+UutjmVknY0OLAQeFa+S2n0+W+/At42uoMDBkGe/xruS2ucn4GPVbwY
VfnEslgd71+VLxne1JHCGlO5DeUz3SRKXtGgxsBTc3cJCro2hrFDFTnWzyPcP4Q+
l0qWnyN0huYa3qCocM20oM+ZssFmJG3nExuqZUsMaDf78YfD4YBbpgB3a3PTwgH2
1PN1N6G3QAbD4FVtySJP7ewd/3lGDJ9Raekd/gn7VczXQM8rXAed7kZDynDxpP9E
yBUJ++Wptzu/8ZhGm9FLD2/WplCmbjl8v9VgBjeO0bQFk0Hfswv5EjDEs7H11Hr4
5z5EciPSlPvjQFxSDOTl26uxWn20447BY2vWMZD+Zq8=
`protect END_PROTECTED
