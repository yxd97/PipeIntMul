`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEjHI0lZukZm4MJ3mNScFIoNlSvZ6iRbAvw6kGZWTCV781A0s/DyNAwjy3JMDXu7
I6qBOOFRijxefmyhacQDfKLH4ccr1N0tGvQKNbQZhrz4T+yq7YMNcwwgKqgspYhJ
lvSP9rM1AYrXDWNSAwKK1o3xUzOi5I9eMUhiI10gvD6Ipq5a3EF4QecuyIN/nNzd
Mxte2EmWhe+MS4UbeY9k4XjCKyMQ1IUrxvuWabGQnaO++oY0WnstK7zlGWMkG91B
+2BuHDnGRub4vo82UtqBaOYh2kGLRDudkMxuI7TfnShep6bKxihHz9XR1OEbHzVu
UUrZOMgQTYMUD4FX5jIcVr7GGkl3CHzpqUgd+98Qq9mBcJA0uPqHhi+y9jkDyply
OfKJKQpZ2Rdadde7REYZy3iZRZMP2Eb/g2s2zXN6IUPmFd0T2+W6As2YTbMuNdm7
//UH7dBtjxHJUWCELdDL5OlO1cvKL5mYIZrK2fzjKLZuMwjCKBk7BIgI2CmkGmZK
yJQ45bTiuq48PInDsPKINILuijTwdzk/EQfcIq2Vw/F1bm2Oslr5E7Uij2FdAwmY
be82G6NsoZBgOcuuTF6i/eEz8c6tqwH/m7WnFq5hYr21ZlxxTpagjt2snBhTgW0q
ylCxJCnr9AOKn7Y04CSyLw0MOI4K22Y7CvKPri60wLzGrOKSvyIXTfkRiY9XH4PG
Bf2gkrb3+BA07v/SCOQydgvWET2IIiAJcrPL4Ej0TXJrIo8Zixye4sCpmyg4RKE0
vWgsAD1b7a4W+2e0ChpipQ==
`protect END_PROTECTED
