`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uCcHue/ST2i7MpVU4Jyk5mHsl/V0eePACDw5rnqDeMHIPeHbD8EFydArLuEUOvNS
TQkPtkJ6G78AtokV+wII2DW2WV6UuFge1Cfabxn/02U7bkfw/PxT27A4W0Jy5IeK
JzXlMrcwFuz0G6KDfGVij10XBsdzsTEcd3FCKB81yEZ2pY/IEp3ZYhVmOXPzTSjb
caIPZiI5YzcVdXxExEJA1rzzFZQb6+2V4uo8iPc8jvu+uMdwLVXCsG7BqzKNVL5s
WQBBZwxOUzzXZxihh+jLWep+s38vFMSw79qvU+5QIdKdOGfzXkIOk1ZFuzXYaI1U
HbaGyfV0V9Pa15vHanKryWhMdVUSOPohSDJmtcieYKkTgEouLm9/8fYxySXOpWDn
UUeMQcua0aHd4cbuBe1ut297RQcUn37j9dzV7fTe+WPv1AT47HxKxRYvFh0e1Knw
`protect END_PROTECTED
