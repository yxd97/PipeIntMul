`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+IzyRADxep77UHALJOE62YLopdhazpuf7lNQYFuGMpFNoOD504VCVQkAHqp2Uhhi
jvzBed3HEX+uX/c3gM4NtBVs7qoZ18bBuIE0Zp1yjxzwBpC1Ckzhc7+hvXVYRMui
iZSZecakV9DThMv4X95MuLkVePmZSasJblFZc3poQXnGrSWNpLjT6AzJky36mm3o
/0Au59hHmtvWXdF1z+R+yNhUTWRalwZYK7UC1gS0g92TBVtTdDED4NhFzBcmrujZ
BuA14WwV43TTFmmAXQRcAjA0QDl8e5jlLRYr6QYXSm8s60R5vMvJx+n3bPC0T55W
FgALxYTnJacP7zkdVUj06t9fqhuHaWeR8foW97/DN5+BesB0tYl82E+iW8rMudjb
Vyde3YjkXERH/WbiX1LQmB+NIG403k9m28/t3ZpbHc6X4as8AFFYgNq/80Itazjt
sBahb/7oU4rhDus/UHiO6Od5crnVuaePQhwj3tPWUUWziYLj4p0z2QcxTxEPzslB
uEagTbUKrFlFTY0OQDdcqLMRkr+HqIPk61tB6m7O6fanQQMmlHTDmv0i2mUzL/c9
0dnJfw3JU/uMrc54YNgVCpJ4hvuV5XL/wjqXiabghwR4u5smqz49yJYgRBKYHLnw
Kn/YD14do5XV3NMRNO/dXQ==
`protect END_PROTECTED
