`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
piC9bgAYo2vinKquM/WACmC32fpxXBLcdetPnZHVbKkv+Xoue3c/15lo2/gOhQHA
PrSpSIIDmy5T2tJwY6cHAAm7RKijmrsr7eQ0r45lKV3AGVcKMey8g5EcT9di1ytr
rEJs5QIjvJpVcqC5qiD1wIKZLD4EyELqhe/0URta/+Jib/Ymp4qZvtk98jkVqzZz
NrqYTeuy4PEVsQnMbZI2j+VRJNus8OlCU5piIOA3UgcbLlpzSbbHdpzxNUsR5Hac
V4xcrSNKXWL+4xseL4KVttopfeVmsoYaTcKU38BIWLuJn1GFtHzees3NsMwA6zFI
/Pexf09toHt3l/+FM8Bi0GX6SFAmdJYo4pmI2MX4AH9GJh1B5oMwPBbEYNKzEi2r
t2Dwb3Byk5ce5tbDPY9lxHhJgnNrBp76/cl0kBNUAMMv5P8E5fKKWbL2Gq1dEdOB
FZTHqhJr6joXqnD5CiPo8JO75TU03aGJoHDo6GWr3NQ/RbtOb0qQ3zXjmBafROWJ
+zanmpE5wUlXMJNoMIdMGEEm+FEjePZhwy4W7O2/Gzp2iul2pUy7DxJzY9h1WeUE
cTD1GEhGZG4eqdSkp7iHsi5wVlGPccLDwEKo1oKsawWupLK8KSRRZhRbQw4byrBM
vuSpVVW2Ka7lonQqZiXmSMD08UpjnWTrHs5q8Ft6jtVfWKn5hb2/5IkSI6FrGtft
pQ/tTkJetasmgcEe/pB3ot87lxK68ChZM5M4kfQeUCX0qbO0mRNdCs8H2pDsmSvi
3MV9L8c+50Nyx6QitrItJlwCpBW7HMvX4yJM85YYNBeHcdxgp84TzrDYK8w6JRc+
06Sf9YDWmeF1he64xZ/owCX/2atpEOXJSydC5j8hkUAy6QOilQLj1EDIDL7qoD1w
WasGv9RzqeopI/VpJw3I4lpRKw5JoNmTIim1IHcBv+rdfmG8ckCG0wWgu9GV78h2
AZqT2MyuAPbvrV6Cc0CSHGFLv1WlWzaZr/+vf6Rd3d1aeXMEM2g9o7y7MDAMAon0
BvS6AsM1j+barrQGp7S7i8TYcetO7RUTW2HYojgyVwauCMEtEOs90Wi+Fy6vo7HM
xkoi9gxDQx4RoNDCHp8+uyq/zfLIrESrhn5Js9Ks6ZhL/aWgt+1K0I64tgXP71At
uyG0icepccfHzwQCP/Y8QuNF++arSTLNGDGVrwWHxmqTcUj2qbDeZUfGgtxPy8Wu
iQcyp2oVFjMyN4dmP7bezVFHY3nCvgmpZt5uERFDFPxJLQAE6ddzJ+Q62KwaLgj9
BERSPw6DFCc/UVJpaeujFkWOcnNVs4sJsw6sgx3plF0Oe5xZRRtKiE0zizdZRlpm
InZReisiZpJ2i8pFZaarQACVxovIdNVInqk7orSND/68qF3DsJo16+q01KYyA08L
3R8CCngZ/I8YSIenDRoEyYy/CUeennwsXmJRX2CxeFnBbZ1nbR/KdJVrQBNP0S+V
hXx3xItrzXLjNjjpi3GckN8gTDN7SRsUXLvoYTEPcS3dtT1g0Xen2zAAkI5buL4U
XowSHmyeLeZdEyyJJThRt0adZz8HK+EbS0/T7bLFrm5WmSB1oaN8sWdRh+yzIwPr
c+BolF2QqhFlrlilF7m2XeNd4Mhr9UBOfLhVFoB/nOpTK0kiPqc8mX0IEs/OOqG9
BONxB0WUxof6R3XuOZtYcRKoCxabzZIanAikkUBCguEsZ9uUVTxTAViAmoU5HT2M
ezvztkmcUGHjm9EGmlSLgzgYdul0OwwhK64GSFXSxuq0m0Nf/CTxy3W1+xW93bae
/0pagRgaVMdJwNT1xOCFSvx7Awrd2YVQrPv7nkg/MDVXh42WPXTbEmABlXfHnLpy
yRk5xCap5y3DPgFoOcw71a01ybm1MrMIpA2Sft4A3RhhF6Dph5WHwGIuK/dYtnS+
BJ3SxT4+J0Bvbs9bQUQMrrLv+Gnnp7eSMHNNlkVdbh4JC5oEMGoBJ9wwH6RO0HPt
EjUvUfzFwKJCnYJ9lTv4L4eavn6l5fazmLfUWPTcseFWZWguYS5cs6tLtJSJL9LA
mGXeUQQPeXQ+0x3gm1od0a8XFqEUVfGejvQRj7TYGeekA0m2bGBYW0TmA7kZs85E
Nqm+X34+vkyVRKgsuHDfK8txpkPf+cOnW2UjkbWfwNLbKQF0g7CJngP+s9Elnx0k
RwG+st2ia52QC/wlYZ5AnJNWyduhIN+Qu6tmXH5T911r1nWN1kC4IWBmDOJMKOec
xL/quz2d7J64C9dD6IxsOabIMAp3ppkzCiI15Bs7h4zx6+F0QmYQOZyNZmzo5uu8
60AgPYlC5akLXDL1WqmPGxZ8apW/6+6KDjfreyvqV+7OzrRCKIAqvio3yqGPu7vR
6ST3HP4B/MGmhmXqzfejIA7iFVO/qRZBOhKPNd1dasQ=
`protect END_PROTECTED
