`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wtpIYZN94y6W3IG5SmdqBVsnyrbaVJg/VzdnxZYYGLXp8EUaZkpsxNYeZuPxmrM5
2j0ENojlgpAuZyJvg4eUGbZIGM4SWbKYTjSYF0zFPYI/hY4g0/NddKsAdcpaUUp1
95fjzTjVWBvxdl6Xf2Y3WJAxDy2cFNtd4BfO9hYmHHMsVdDndpPKUTlFA/P39nYO
Ve+NrLsmb5XANcx4iG5kPQO7jbuZDgNDiK2Qx5HQzVTwe74am/AikBi3/7AVO5Uf
HVe4VfEq3o86Qs9FNykMF1kRy8jtDO2NpcgNtxHDTr5VInZ4Tz6le+P7DmVxnsF9
O6LidWvA7bslbXI64bmdxShulnWNoldXi2TYe8SSTxb+o28FZcXKNCHG2qGjAt3a
5UqiyO5u18SM5GkHYhmUhQXirnc/23LllasHaV1sKVNM0kdkAtql9w6tesykppKz
7oK3rl6g7pABcbJ8LM82N+S14IzXyi01hfOUwvlZhRqtG14lgFxJ2fSpgaEaHZmA
qskEGBqJfP7CSVeiB20G+wHds9aBs/lLifF06Uy2s/9ZADCIAArXCM/z63gYg3O2
/G8b1L+YmiV63fVoJs8MKcUS9kM9UM9JhE8UUC5/bZFrpAVbsrckGmuWrrBLZwTH
IObyXrT3fv1x+8J+V3AjZUUtO7xHnpX5dhwX8K6yrnPEDmhTTGlk/yJYJ8kuMRbD
fEaDgVH+byY3l5VAVIg0QzVO1kQqOeq0//BSHswmfna96fkT4jzwl9WduesP2PXQ
MJdgk/dt7k5UEc05zLpAVBfhIRtQ3qJawyEQyt/dXm1jhjGH7z1sv1pTs9StZ1uS
6sDZ3pxShescjXVTbjDiNh0dM03afcj1qJ0jJ6d5kGhiNXkfDPrd2QaN6scJmd7c
ughgj37aNQndo3OJw2Dhcg==
`protect END_PROTECTED
