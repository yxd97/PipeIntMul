`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wn4K03thS9uLow4Vlb3oSwBgSfxG1kYlh7xbuqvwATX8OmXYF+ntt0HmQ5oIuG6m
KRkXeWAJ4i6wE1KiIboaw+qsgP2N98Ws1zFhqV1hL5dPMElP2WfLC8SYeKN5Uxj5
o+biZAJFi83yVP6M5AOs4kAlKdG+amVkEK7w+xUDGeUr+e0WndExHsrIMpTLgDU9
3ziHjvgkgsFaU3tA8gbJO0yNh7wmYhN4D1hDAoEo7tGecluB0G+w2cKF1tyZPoCz
hfZbF7f5AKL0A4XJPCnoUw+AGu35/NRqbfB3Py7tNGa3fthoX39peFWDD1mvxRUZ
kTP5lOgw7oxbcgAMCNzGGgVSThdz6WPglBiBdT/JYxLw7007z64qopvVNkcThR50
05Oy4mcxifRQIdYX1my0R3p6iFAQ4GK9CzLQQyFLd6oUJASicwedS5U5bSUpBBra
`protect END_PROTECTED
