`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0RsszzBN2FAe/bXi297DWEzOZapEz0cxPqXndrmrPKrm3vRo+ZsyFhsue1Zk39RO
QVKwNUTDe3y2o/2jc9igiGSNr5qqOjqC6VHrHbSBVbAOVmLq4ce+dBXMprVOJZ85
ss2FXuPeH+rb4Sg8jGfrG7hRzCrUQoRBNYMiYOIzP0g+cu56lp0feMxI8cW828jc
lRKVziTQIJwof+RtpSfrV5R+8B3d6wZoIJQHUrwePf9Q9nH42ij9Oifh2GkPAKVj
FFm34Ej+s1DUebwFqm00rmcLfbcI+LULyTh0/aR6UOwzF5KX/BboDwL8YuhGGGjz
oM17LuBL0aCJh3oWWt4sGOm+nn0wp/4vx2vKxNARVIUOPgff+71H7fbf+4+RT63F
kKg6kAb3AS14IoYZb8eRBiHuzfTUfhE5WYgraZcUZkThTjV5m0wlkYMjNvxD0YzL
QGBJ/x3YrCtbIXNQKY3XqK2fb4VuwAynLYTYuhv8GLGbdmFD6Yj0HW5zb7wn0qak
`protect END_PROTECTED
