`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fVp6KBEtY5bYj1wt7N/9s3oS8+ThYoLrWNWcq+hLXOeMUulzSM+rCJS1uTyQkjl6
OQzLFIg5JfkhpEK+Kd+8mgEX6q8+rljh5lx7zl4JsEix01aefzgWee5d0TPGrgHO
LvsdeRwRw8drf760rboey5jmLcThzRqgwdjv0BO57ta+jBrXL+tX/4PPaFvNn4ln
T4tt8fMW7skOCh+uUA6w1hjb75NIPtqsjBLrjtE84MGRYE8BGiG/T2dxMw3fCBIZ
vD0ol3PFh0mS0WsV0f+gcXAQHhyx/Qc3Vlj24DRE4A3SNaqCxNJ0JslUL9EwnN+u
Y50TFuDhSuDj1yXsEPFYu9/6m+flOF8XEZmcetvjOsf4OzMFMz+Tb7FyZXf/9OjK
TCSIN/TlEiZSrPe16ts108fW9ucuG+qbJY/GWlVb5tyNjOiTFj0wQEcLx5zPUgPV
ajePZlyZF8wakNH5HfnOGOuHO7oeBREe8ce4DIbaOoBZK/XEZ01NcOuq2BfXwy3z
UZ0939IJ2rl0htqtc4hbCc4Ub9VAgYmvFhV2wNZBlgrekzQch69SiVCz4A1rCkDj
PHlwLqJBojq//SyDDGTsME/bMZEsmsLRAec2jlO0xbEEWZfwL4NA0cOEuPqvwYNI
6Fa/QPWngHyrfEEIGZ586uIdwqlTsiOndau1BuQPWSFTOJoLPugFB+N+S5lLIOf+
VRK00CzVriseCHCJOSNnvHXjGs/XL0HVYnPJEPGL/Rn39+2xz0dWAZRFDekT47Po
2L+rii+DHgZunXvD8OqMh87BuGGXkkY+N4HN6YenX9gUpi27jAVa5NzvMRNfIfZf
`protect END_PROTECTED
