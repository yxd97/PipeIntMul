`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3IETZi905RTiXkLjnWzT370HTpzL6SGkGlRuwCQXrOsrXdmZZzj80hBSv4fbSZuX
F4wsXIBkamMpT51AEO9oumLpiSCXS3qagl6RE+ODmY1sp+3zZJjfN++CLJ2C6YjW
u4D/tp499L1W5S5/m2OwJ6J7ER9WAq9FSN8/7YuZcrX5/+hiIJZqXt7zEgLgwD0R
Dqw0NmmoT7td/Zrxr9srjy40srDlvSLkJsCA4daaUIjBoGDjFzpG0sFTjZsnkL2b
qBRh5bFL1Y+1TzHYsaJXiIGFzBQgOV3mPNGaGDOi+Qk7oMMQXdP9y48i5RRLNEE9
gbf6rGKbvEsJnBfLnNL0hJQY5lWoaV4OWv+4JR8fCNLYNiSXtDLYbHk8AJCXggI3
Zg8/FASESa81GMoK3sNP/w49rIY9mPKEqvrljnJ6X+ZpJ4L/NJCOKnGreoYJGF5s
je24kMXpYmb/cDYaHWTohd4OBpQJc1IAHyZLOIjmaom6S3gf4K/qk2vt1qRokbXb
wurB64clE0NrDlPTcyVvYwOv+oYVVW4NnLIevM7/RIHqup+L1VzXTGoHOLuaeQNi
OYS/iVVEE2jCCAm6ihlId7cPiVRd6AVbwDomhYM4NnQkNRmQutmp7IQpqBI2zFgg
tMaLEBfys4+3yDHeIjlVAdIOljHbAbDNYuTSCLcdNDXEDWO6tMdsTQ0q6e8pDMLW
sPiI0IVfEf5kIwmHYBK8XsMKnAQSJ3V4MQi9wf/79v78vME23MNavcvOqh0ra8Fp
H0fIXLFRvHAJB5Df4VfsoIcOjLP47ZI1h72ESQx69blKieHTxdtxRQr3BYsHIzTV
BKapofWYvkwnsGmfUE7A9lyPt7d2KYofekctp8Bxttj3/hRh+QLdDRF+gHXWY2pB
lICybZixa8PtB0Xqco0ONbqrku8DR+RZhN3NW6LAWcbAgdO3ufIXyR9T5cnbRIlv
l/zA7EuUhlA1pFz26JoF+9t8MgZbnAU8i+oYef9mO5lUlYpNuE4lmgdJvexnSKxD
7ATcfP0zmvNC4YM4D7m4cIhM58/o36Kv5Mhu6MtqeDZuvB7jycvCpVxw7/YMqDPz
h3hyiC28uWGHpFeGP+tOw0OkxVXSQcvCVoJSaTSqghi/bzayU2LBgHOaRKEDv4mv
UDqIdWgMsI1OpVRrfKh0WF1Bz2Z+jrw2BzxHOGxYycc7qLgKXteH913SU0i9kvkQ
67FC0ge7wQJPNwKBUuUGTZJgz58qKYDra5gqeaK6+4BMXeGCykL159huY3alKwWF
rBOCbrX7Tb02VkwejoJy9rpbWsyyvAoImVOKq2BNXcR1Yu0Q1IWybTi/tKi4r4MZ
cAMj1pI38SidXfb9BkUq6ucVJOWuqaHQGWbWCmJn0NegOugb0h9XL1QlCSRwW5xb
2OiJA+hWhC9Akud7MJ3JZwZqzSdwxDXFwQCinEYktwGxNKAF8Lq5Weur+TfJaubS
TQZ0dKDB7lpkXUDJH+VxRKLX3hqZHkKk/A7piUIbfVeD2yRFwrLuIV6PNEnJI0d9
IhGfMCfS58u55Ir6gk4bpBbbz5Gh7dk0jmQVbuEbA1V2F9YZQ+QmmSlf2hTY9zMJ
8vUsbMTdwTPyDmCmxs2n1xkHWJmO/71eJYMKwj6mEXCql6x8WdOaynk1SkCCbZyk
VeWCug/J5TAeGJUGV+jzHyi+MccqkPIddc70MmXNCkI9Zn+TYgG4escTX0rZRZbY
ifAxpYmx1YPt1Io0CbaD7cvdeZ9InfKMf7V2wMCo2GJ00K5ZVS9GuzTD8YeM/Sji
+QD7r271OeRuq+U/dQmzuZqRjYMuI6WRPaESBVChREwDWRqum1ngXy4nNGF8Z58n
qyLGIsuOSBde52yZ0U1pOA==
`protect END_PROTECTED
