`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w+Wl0PUgFMKLHxqO6S3V0YRLg05zOBJyl9wvDa42tgjytrOSAzv9zcea60iChkcU
aB8Mp+rzHSCeFivQ3ryGAPJPfNMhUazq/LXniLqWGjJp1eA1WSu3VbwSFioK668d
9i51vnKNfw/QlfvdANxWWiXo+guaEhSPjVzoQ7lo8/n368u3b7AHkS9knw+S3JDC
5h5tQQFtH1NrXzGTEXlLpacOCJUUYbSUHq7gzLyYyOVyRVxvRpTz8C+fka9SqCwM
phsXh1nk/4HbgjsBQsU/r+HSJKl1ncTFZrrNoZP9Ww9nk0/spH0OQ/GUOA+kMkDv
J8mEQnfZHO/7nwrma/s0gPqe2IB/bFlxp0KxfL+0/DCmgf1jNMtUMcfsjE5UJFmm
3ewZcwBj9nfXfIC33of1YwOJ8SPxv3Ig8LzOgz4je0FpZgw0Smj53B6dVDlnKnHh
dA+DJnLzof5UY4dT7ExPSWE8m/+sJvX8X+sdOx51EkreOb2nr3R+lrTOpaufjTjz
87hgvE+C3lNKHN3UnzZkB9ruxWwg6q9VdzC3KpJjBFd+52X+Msu+1erkyK1lNNTp
KN82nwRP9ZxPy3N1vrAP0jefLsSLJVB9DW4V1A43C1nQNWNqi6gDlbmFLxlyibX1
6ZRq6EmgUMlLm/tpQDg5oR/XCoC4NHF4pfvvrSuvf6NiRN6Cc7VnTcRwjoYKpY0o
xuP8m3hPa260UXTIlfUH/wVl9CDePoYuPAKVG7JPrqX3AfIu4VTrr8/p9uJARwhK
CqFuk0Twq1IJZGBwzd8PwlDLIYiz9gYm5xdDkGqQrprrVPaaIbt4fV1SrGV+a+uL
E/exvgKTe0z/8UO/D9la7M9rwawuEjz0HKsEeW5Dd5E/me5jBs5CH7r1BVN70peD
YHrWG/lc2wGWz/CbOk172TuFVbGGL1ruV23ogky/2C8Z5FV2c1EloelvGA6lOdA0
ocCVcecV9sJOj5pdNkvfr8ig6xusQ0x06gRGTSY46Fp5UIQJp7f31GYj5FY7XNQI
fsT+Wef7yPFOAWVSllqdEw==
`protect END_PROTECTED
