`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LVrAR1w0aiOEMp7g5ZwiHkFZUchOBgSoeZa8MjGzdSddsoZ/1JZnZCA2lwKvby/2
ZIX+C4jHUmzMBjFNcX6vS4bv5OsF7YDw/dsAL5+SiFeBCMboqJB/TbAulgAcErKE
bfd2RTq6tTVbwrJ3ixUA4qwVuj0mczcLPqwsJK4sxOpzLSHbBh3GMa2IlUWiX1cr
gn45Y8XRKhT6BArf811Y3pg3a/HZSbJ79nQeRyt5+zPDN8XF1eLgYpxgEoX0dECq
vfxyp3kLK5uk9LBLRJsahyotcQ9evCGGixD88aXpuRin3XEh8MmCoPn7Swv4L0CB
UQjd1p5FH1K1KR3lzqWTI3sri19Yukz3hqe13DnBczHtz4wwiXWN8VOiiLDCkKpa
TKtQz8Bz40b43s6VbrdYzYN5jESRHSShovw8DJz4rx9VBKxNpmRbWzI8PUL3X/4F
hHQZM0wSy4VNzKyuMMWojoTV6OibPHRwrkqdq7vg8icVVzXb1AXhtQcQVkDm2zNh
ecogoJGe37pco3GL5+G91FN6WE521FWiCZFNEsdQjOgdsAuqsyvz2uhHtTeVbStl
P6bJK4DJeA3A6OBtpwSjl0qUnJ+3vUPPENdQmnEoVnfDEewmWUfS1Asap3ikZo+I
rAQ5GPVW6OsC3eDciW4PN9CEP5D0WqUkv5WHb9RtZ2jVKTqssWoAJ7wa8nw4Q11o
ve8pgrfZPJpH+A3XTmXoFOuT2oFZMQL4TYS6t03KLIMiRenI01LvaN3Zx47gK5Jy
xj/MCdriIV1ZfI6vNS8BWuQ1dV0FijLbFQk98t5KrPsebjv2EA33tBaVpvV3qhJN
wlCiXONCSEb7/akF6PD7M//A6fCFru4AbAjO0fELcwS2avE4PJonNqOj8HejOsX2
s7N0M/Ugbv2aqwq4kd/OfbqZLPRkDkKFIgcHGdJA5tNPNTKDVcrHpmmDsdAhO4FM
6qcXc0vtfLQqJxgp2nk2rnJwBdziVHaH9pANlREKDvjD8CtHM0mBq2QsHsmsANp5
3ct924fNIBWVFgkTqlNBaurx0PiWHr1ynu+FyjATIZnhYy84l2jKl9uWRyblAey0
1BXstrhxguSsNEhVK9B9KKReOo5Bsf9KdUDYLozgFsED23tHUVPnlkDbTmEtP8Vj
0YnP06qGeQFLahcodHFuTyXCGi9UGw28ZWN3WmMCwnNAeuB3dcG7v6W9J8wE8Pm0
MEPamzYZJeOCgdmI953PntLrxLoL4jgPlZmkwVMHSFaBpe0iPYU03qbk5T5IWiLy
X/eeORsL0YP4NW4lERmUkLU7bVOYa+5UuEEWKhy+QFxPCM/Scoh4D1mbiIkKeveo
NCuCF1gQqO/oxfMcjqMiZj7/GoFp49x/HVjoUcYMonEUlK3tU9t6P6K7CezXN+Mw
EjPoTfSIUCdFRRuChXpbIZuenNFIC2R35NUV3iXeGHXw/GyCAfkBPVa+xvFD6L/c
8pxUF4Q8nNeSc9XYD/6cx0i1iQFEgwkIH3gnKF8Nf2ntgGj3xJ+fRMBu6VkYyGZ6
lwElECtV8zesRCxocR8z0mFlG8UFXygC2uw4XrpATQ3tKBRNp2pxlozvQlK/YN0s
SeVngfzdEyA5C/ucHS3kvLDaAlVO6fldY1vdBDmlojw1M7wHCKua8i4zOCUQcfiF
0G74VwtNOuX9ZFS2GXmGq+7Ws5YXr777ft9kS3q/6Muk4lkAEqW0AxG/WIfEVdsP
wrJ4niAmd2p6RGQ2fBfqJ/vFnzeKQkbvMgJsnu8Oh3LEeYVOCkdbA2S7X9PFbs8O
sjXWL4ky04i9HoxNNNL/qYraXEVfFYMWn9LzeBSqZAg9jCGauhLYtKeDtD5I+L4m
d7vH9h4LKe+Lzn+OVE17yKS1u/SeqST4iirGw+NfSK4C9yjGc+gvSQPBp8s1QALo
iH7eoYDusIBSHCKJ/oipNsg6tctnMHCX69EBRk2VaMVVlnmWgBJznA5gwB/yv3b2
LlNNS/7hzxzqq66V9o2HMb3GvrfodHEyZ49YHstRhn9vbSN2HcSalQP0A7bMwYkV
xuDz+xWlnvhU5dsOenw2t6hEpFMlzTo4+qml1o4stI9U+WKvJseWZsXx1rUIUFoy
Ep6tJBpa1tyC6LbgxMBtrztvV7fhCTI4tP4EyVT9zw5us99wgu70OGHvlXce7NTM
+5yKvD1Qhb0C6131Hv0n5m7NC4DTzZZESwOWTj6duDTp2w34ixB+8IPMaVzOKqAG
m3TKf0/T23xEg7EN2T+dfb9ob58+6FB6ik0XVz6PypzMcdwj+UiZELUEX0mkw1vm
lFj9qjf9uHJqtb7pVOLWZ4Jv65stMxlhV+pyjAKXjxrnxJ87BOe7I1obLFBMVrnQ
GbPTFoSOAaNKO7HCE5dSQTlhAEZ4PqCx1AOmahdnLnn76CVCLzAP4CRymt0a+NWC
ekRVYaxeiMjwZGkJy7nfRPpmYd9XvjZgAO40O1QX3J+LQm50ABaFJGMa9pKd2EUR
BBMZg7zW+tirVRy0/PgHI0SBwfBon7RR9knfB5FqH7Rh4DwtH8PMeJfUI2fgsb0N
YsxoSZUSki5VKZfQ+Avpir9XHxBGCnToBJ3qroNA35AdD3YZXXJ+SB0jF4391WdP
lzcaYjzSPZ3kq5sRr2OpKcq33HLRcQR39ATejZwScNtnnkEuPW01/s5A+wACWtUd
cmJWRnb7MFwuab7V15hQ3p94H4LwrPm2WB6rOq4UybOA6kVoJWx60fp340QWOVwL
m6UfIlIfBWMobQ4Z3ZZPlggd4cq9RA13/q8yUqzThvrxoWCMPF48++ir8oDJaKRB
6RXgAuFsiY0wv1PSSxx684oz8oHOKP0WP4H11yxpl3IGgoEjgO+G/PBZXCfWdWQu
oduobezKB4+Bm25eTVf7XEu+vJ9b4krnuNoxsyKxZa67q9Sh8J+c40qcptNf/ilc
zoRIXit/Kjyx7ilVPCbRMdi5EhB1EatbeinyBDl+s6HTRlWAmstQhYtwL8g8Xu9k
Ab7ycsj2/ty0FdRz8/pQuRlW/SEMZHFdZxHpvW63Q94fkBQ8MLbAplb6Z3c/lkin
aSIEmpXq7VH6jX46Vmb/rtY2oWizCxz00IKEUun11jvWcsi9bNTyKTudBEDX0fVo
moEsEepEZGx83RoFWb+4xnapy9BnqSQYHiLDOl7IbcGCLK3D9Ta/a52vNGbJ/aD2
xtU5l9KefnTURnck3m6N5G4z/8+i/B7SWSK6j/UT7WQlW6Qfe8KcqYY/43dLw5Gu
b4rEZeV/bohNziTfX/9kJSVpB50E8Fk9gWV8JeSYic4fnUiH8ib0xL4LZjSm9E2X
ttkHPCFpS7vclXg+TUtJ77BSsIlzAPv6vNH9rVE/FTKHCApVvCHy1hHciDUwaM9c
y1DYy1w8pEHPRO+k/4ctiuLoXYGiOJBDwMlDQabQdmCOnQG4I2fAkyw3DxDeOdob
xOG0mLoMNsu0ZXJccb0cU29cR7wnv6hf5pgPBzMITc6omRnIBI6AV9EAasSoZF88
7q/JEtYopT4tJrv+P+jGOtPcPDe+BN7jPP067FFWSfkxgLLLuvgZ6VLps6VWjq+Z
DMVfTOLM2AL1AfMOI0wG2U6e4UMYZeoTWB4x5StQryU7Lwm4ZAR5xnwFOmNDFKuO
3EN9cNGZZM07yFlWDXP0fj+bq3SWXMdeW+9KyXqa2cg297oYnB1G55STISZCvZtD
dmLjdEbJ2UJFblgwNy1h/dAiWKdE3rS396E94sd6TqUnAREqBAM+scC5EcEXR/bP
U4pprL4vgrTCxHnMpshmgKfvCqo/n07ONTKd5bvwsB0f4xu71sDioe7xpuZrBAPc
gTUXJL7fXJbF44BYf8xpq39A7Hb4YISFJ/O/XxBr3cywNCfyawgsHhGCa8QI2KbK
Fjx9caM1Wrw2jzcRH7c21W2I3A07YcDJJLCV1Y4aaYvWDf7aMSNQw55jGT4enPq6
DGpq5rwvXwir+SHuHE8dedp/QJCcIkAsTNj18lhde+rkX6EN2kiNXqLkyZ1pBvc2
ZdooLTiwNSkq/WTdyXu9jEr/FsRwpnaXO06eyq6t5+2Q1hQWxPv9yPglwxYf0Hmj
eP5a+noEKe8zRGeTOq86Cd9FRErOMF3PEUddwdj0lahOgizXWeagYPyIu0JB6So7
IuZvtgWMflOkr94D258lC6V0MTp2E1JG/9yloyLilGKM7cOZL1MtTecEVj5341ko
3SX4+8XDTua9vURsN8FdzLWqbFzo+d9KOeg7tbfCyHyXcYjqe6ENNeBJlFU/fwUv
MRT85gfh2Jo1SWHmaqG5m0WmHqrAbIm5Gk04UrS2e7goR+3w0WqVB4Xfjgt6bziV
+H6guAHDXMmjWPLpEY6uA5R05aif0JLZdlRz4fnYRCNUi6Dw6qXofIBO7lTUsH1Q
CyKOdjdOPNJghuwcDg0lynRXPMPFJNY6nRzissTA2khkCAbNFHW1Yo0rbd5Eozft
LeZKxjoosDBnkXC4pDjftwG9eEU4pRrgkHTGSJg40pldR+yfYksIOYEP81TKz+AK
dwsFDWrMkUR+S8QTOScoc4Jgfvc3foYBMW/3QxI4hlCU1PB9JOu+wnfjHm9AaL6d
0m+0LKoVAkMmXDPxPifQuOStdALOZH8fx+y6WUJfL+Q/7tvIQqSMxA47LmZIe8Fk
IW+jbN6Y+kHMmSXJ3aeIA58VNjkwxnXWcmwwpA7c9PPyMMpS/Lp/qDkFWh42Rl+c
FBCiQg06Jh/lQqhy23Wun3eBQPgEjg1CfArZop05Y9nJe2XUCL0u25ooJguR/FH8
IDVU1uRdEHvwMkKytBFpEB9OzvN71A7REeCo43pEXAn5bAS3M1n4/vyOxjxduvb3
h3xeGJpolGiYvYnG2nZnnlyhntist9Syfkma/65q/YP7iI+rT6Bq7N+UaeQAqbZC
3NH83sXpFdBJpitcvM4Qr3kV2sbF9UQpl8odMy/33wVwulrt1hC7utpasfeJW2EK
cIYDIIJ5BUTgrKToIKnmMO2t3hwH9x2deT5IEbns6BPY7AH+Tv5h/CVgwud5Of5u
pvLRCUikdmJh2gurkJxLzefqn9kjFSCKJQqes3C4eg24UIihnNtlKLKtPpPNNXR6
C7ThqSfwLTCXK9eQYmjucSqQwCvu5V/nOGbITqCUDBBUOYU2H3EEL5ErkpMX0GYr
vF2HoEnTIE7/+mDaSggsumcDnpOzuxfAanC0qAbZLfHTmCdhpM4Mvkje0YvQfhth
XfVJ7T1MQExnhDTL1gWIqJjiT86y4qz3wH0hmTEHwE+zaB7P8snSvsezOUfUJHeq
l4j07idLGsjh9yBGILYSDhkMKnAs8Zu71cUodFVCUSbDKu9igbEXWTNsmSCkyAHb
GBFrM9886PcK3KTp5uIfW5MMmqBpwM/LpsA6m7KHBF1taZzH1ZyNLJGRpGqw/s3V
cYAmgFBWtiy7wrx01SvzrmasZ12acawp1flLKl0cuC+/X6kxuQDRsBWIW7HNBJtB
0+Lzt7ehbns2rN1Kp8qSYkJnIvjwFHQnPJdR6nPF4ogrjCdKXJ2Im+7JDqj0HCsd
Zwe0sDpsHJiJmysLT8yxuTMBQb/oi0uHl5l9/oEtyCOokXSDrYx0qZaBCwEIq9aE
bIvGx87QMH8XP5ctbKkX3fjmUc6+FrJl8GdfYkKBrwx0tBBb9w9lG3Xmw9BxLQOb
qgchbqMbBHWi+HrypQPiluz8OYVAkL0T0qfSpZMNdeP11FWoOHIGRQWd6IGHrqS0
BN3y8QX5k5mbgftMTL6Q7jC9C0QdBoCuy//9yxZnHgWloANedksFK526IRlXsnuK
3hAhBA+rtQ3kIgSvrNjeQ0tiv6O34H//zI3Icm1qmrtNfd9eHiMQRANepagsRHEA
I6g/cMDxQaVterkFWlSSemgr5MwRqCByvsnO2AJQPhCxEzdsTfoTISB7N6aTInF0
82MKXIBNzeTwOi3DEfMs5w==
`protect END_PROTECTED
