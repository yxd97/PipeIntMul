`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RJyHwnf1OABJFL5qDPxTqPOSE55z2PG+3SlBLYKiBtM4vsI/egwcw3QuDbj0RS+t
k7cisZyrg92KxUYQAlITA/MDblLpoX4ZpMND5kpZf5I+RXSaItGe5LWMH1P6ZETO
ECiCDq1mRayBjxX0+n9BhTrDugYqkZJlo+b7GEX6kuEoFzfYVMxloJL+xt2vUUYl
8fUcWAy6pKfvruc4tZPJo0lOGYEKjyKAVv3vfhJyq+k0+aRl9h/12icHSV2mhUHk
1sibqr/b8Ia2+R59GGwiNKK2P+l3Lc7WgwYgEy+GQ879zfsjtm4Vi/KVL7SjorkE
vh9FYYSSty1jmwpGuNVYdsWwgxIwwClcrWRG3NtETEc/uoCJnUNNJVqlLOTUHHia
o7EintCulCntXumAe4dfv/+E329QvI1ixcqkD78YjU0Y96e8G4nJLv6pE7fkl6uU
vJpwaXActTJhv9kZmdR/Z4N5ayrz3FHQofjpwQczg0p6LdEtnBg0Z1//r4EFPUbb
gZnfVs+npd4IKWnT6N7P0w845xKNpNQWQNiOMloekW4OLshr5o9gqtNkzrx53Ehn
uGNjUg4QEuVKgjfq7bUBVCZxp2VKUSzos826VN91uUsiC2C5Jn/4jZ8NlgiXeX8T
1OZmjxY1mcakGoJk2Hig9NxnMnPeOVicv+o1xSc6W1x3R0OL1he34XjmajKnn9o+
ABlyp06iwJdGg7Ey7eUeKR6mzWQbpFCS2baAeGzD+tfQRwoH9yTMVi1Hp8vbDs5i
man/8vDadjNF2KgkX+ZPrw==
`protect END_PROTECTED
