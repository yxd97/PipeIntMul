library verilog;
use verilog.vl_types.all;
entity X_PCIE_3_0 is
    generic(
        LOC             : string  := "UNPLACED";
        ARI_CAP_ENABLE  : string  := "FALSE";
        AXISTEN_IF_CC_ALIGNMENT_MODE: string  := "FALSE";
        AXISTEN_IF_CC_PARITY_CHK: string  := "TRUE";
        AXISTEN_IF_CQ_ALIGNMENT_MODE: string  := "FALSE";
        AXISTEN_IF_ENABLE_CLIENT_TAG: string  := "FALSE";
        AXISTEN_IF_ENABLE_MSG_ROUTE: vl_logic_vector(17 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        AXISTEN_IF_ENABLE_RX_MSG_INTFC: string  := "FALSE";
        AXISTEN_IF_RC_ALIGNMENT_MODE: string  := "FALSE";
        AXISTEN_IF_RC_STRADDLE: string  := "FALSE";
        AXISTEN_IF_RQ_ALIGNMENT_MODE: string  := "FALSE";
        AXISTEN_IF_RQ_PARITY_CHK: string  := "TRUE";
        AXISTEN_IF_WIDTH: vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        CRM_CORE_CLK_FREQ_500: string  := "TRUE";
        CRM_USER_CLK_FREQ: vl_logic_vector(1 downto 0) := (Hi1, Hi0);
        DNSTREAM_LINK_NUM: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        GEN3_PCS_AUTO_REALIGN: vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        GEN3_PCS_RX_ELECIDLE_INTERNAL: string  := "TRUE";
        LL_ACK_TIMEOUT  : vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_ACK_TIMEOUT_EN: string  := "FALSE";
        LL_ACK_TIMEOUT_FUNC: integer := 0;
        LL_CPL_FC_UPDATE_TIMER: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_CPL_FC_UPDATE_TIMER_OVERRIDE: string  := "FALSE";
        LL_FC_UPDATE_TIMER: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_FC_UPDATE_TIMER_OVERRIDE: string  := "FALSE";
        LL_NP_FC_UPDATE_TIMER: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_NP_FC_UPDATE_TIMER_OVERRIDE: string  := "FALSE";
        LL_P_FC_UPDATE_TIMER: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_P_FC_UPDATE_TIMER_OVERRIDE: string  := "FALSE";
        LL_REPLAY_TIMEOUT: vl_logic_vector(8 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        LL_REPLAY_TIMEOUT_EN: string  := "FALSE";
        LL_REPLAY_TIMEOUT_FUNC: integer := 0;
        LTR_TX_MESSAGE_MINIMUM_INTERVAL: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0);
        LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE: string  := "FALSE";
        LTR_TX_MESSAGE_ON_LTR_ENABLE: string  := "FALSE";
        PF0_AER_CAP_ECRC_CHECK_CAPABLE: string  := "FALSE";
        PF0_AER_CAP_ECRC_GEN_CAPABLE: string  := "FALSE";
        PF0_AER_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_ARI_CAP_NEXT_FUNC: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_ARI_CAP_VER : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_BAR0_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_BAR0_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF0_BAR1_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_BAR1_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_BAR2_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_BAR2_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF0_BAR3_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_BAR3_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_BAR4_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_BAR4_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF0_BAR5_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_BAR5_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_BIST_REGISTER: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_CAPABILITY_POINTER: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        PF0_CLASS_CODE  : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DEVICE_ID   : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT: string  := "TRUE";
        PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT: string  := "TRUE";
        PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT: string  := "TRUE";
        PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE: string  := "TRUE";
        PF0_DEV_CAP2_LTR_SUPPORT: string  := "TRUE";
        PF0_DEV_CAP2_OBFF_SUPPORT: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT: string  := "FALSE";
        PF0_DEV_CAP_ENDPOINT_L0S_LATENCY: integer := 0;
        PF0_DEV_CAP_ENDPOINT_L1_LATENCY: integer := 0;
        PF0_DEV_CAP_EXT_TAG_SUPPORTED: string  := "TRUE";
        PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE: string  := "TRUE";
        PF0_DEV_CAP_MAX_PAYLOAD_SIZE: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        PF0_DPA_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_CONTROL: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_CONTROL_EN: string  := "TRUE";
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_DPA_CAP_VER : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_DSN_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        PF0_EXPANSION_ROM_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_EXPANSION_ROM_ENABLE: string  := "FALSE";
        PF0_INTERRUPT_LINE: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_INTERRUPT_PIN: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        PF0_LINK_CAP_ASPM_SUPPORT: integer := 0;
        PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1: integer := 7;
        PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2: integer := 7;
        PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3: integer := 7;
        PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1: integer := 7;
        PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2: integer := 7;
        PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3: integer := 7;
        PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1: integer := 7;
        PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2: integer := 7;
        PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3: integer := 7;
        PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1: integer := 7;
        PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2: integer := 7;
        PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3: integer := 7;
        PF0_LINK_STATUS_SLOT_CLOCK_CONFIG: string  := "TRUE";
        PF0_LTR_CAP_MAX_NOSNOOP_LAT: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_LTR_CAP_MAX_SNOOP_LAT: vl_logic_vector(9 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_LTR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_LTR_CAP_VER : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_MSIX_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_MSIX_CAP_PBA_BIR: integer := 0;
        PF0_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        PF0_MSIX_CAP_TABLE_BIR: integer := 0;
        PF0_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_MSI_CAP_MULTIMSGCAP: integer := 0;
        PF0_MSI_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_PB_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_PB_CAP_SYSTEM_ALLOCATED: string  := "FALSE";
        PF0_PB_CAP_VER  : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PF0_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_PM_CAP_PMESUPPORT_D0: string  := "TRUE";
        PF0_PM_CAP_PMESUPPORT_D1: string  := "TRUE";
        PF0_PM_CAP_PMESUPPORT_D3HOT: string  := "TRUE";
        PF0_PM_CAP_SUPP_D1_STATE: string  := "TRUE";
        PF0_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        PF0_PM_CSR_NOSOFTRESET: string  := "TRUE";
        PF0_RBAR_CAP_ENABLE: string  := "FALSE";
        PF0_RBAR_CAP_INDEX0: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_INDEX1: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_INDEX2: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_SIZE0: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_SIZE1: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_SIZE2: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_RBAR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_RBAR_NUM    : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        PF0_REVISION_ID : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_BAR0_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_SRIOV_BAR0_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF0_SRIOV_BAR1_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_BAR1_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_SRIOV_BAR2_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_SRIOV_BAR2_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF0_SRIOV_BAR3_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_SRIOV_BAR3_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_SRIOV_BAR4_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_SRIOV_BAR4_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF0_SRIOV_BAR5_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF0_SRIOV_BAR5_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_SRIOV_CAP_INITIAL_VF: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_CAP_TOTAL_VF: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_SRIOV_FIRST_VF_OFFSET: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_FUNC_DEP_LINK: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_SUPPORTED_PAGE_SIZE: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SRIOV_VF_DEVICE_ID: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_SUBSYSTEM_ID: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        PF0_TPHR_CAP_ENABLE: string  := "FALSE";
        PF0_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        PF0_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF0_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PF0_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF0_VC_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF0_VC_CAP_VER  : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF1_AER_CAP_ECRC_CHECK_CAPABLE: string  := "FALSE";
        PF1_AER_CAP_ECRC_GEN_CAPABLE: string  := "FALSE";
        PF1_AER_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_ARI_CAP_NEXT_FUNC: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_BAR0_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_BAR0_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF1_BAR1_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_BAR1_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_BAR2_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_BAR2_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF1_BAR3_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_BAR3_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_BAR4_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_BAR4_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF1_BAR5_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_BAR5_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_BIST_REGISTER: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_CAPABILITY_POINTER: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        PF1_CLASS_CODE  : vl_logic_vector(23 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DEVICE_ID   : vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DEV_CAP_MAX_PAYLOAD_SIZE: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        PF1_DPA_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_CONTROL: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_CONTROL_EN: string  := "TRUE";
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_DPA_CAP_VER : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF1_DSN_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0);
        PF1_EXPANSION_ROM_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_EXPANSION_ROM_ENABLE: string  := "FALSE";
        PF1_INTERRUPT_LINE: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_INTERRUPT_PIN: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        PF1_MSIX_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_MSIX_CAP_PBA_BIR: integer := 0;
        PF1_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        PF1_MSIX_CAP_TABLE_BIR: integer := 0;
        PF1_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_MSI_CAP_MULTIMSGCAP: integer := 0;
        PF1_MSI_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_PB_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_PB_CAP_SYSTEM_ALLOCATED: string  := "FALSE";
        PF1_PB_CAP_VER  : vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF1_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        PF1_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        PF1_RBAR_CAP_ENABLE: string  := "FALSE";
        PF1_RBAR_CAP_INDEX0: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_INDEX1: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_INDEX2: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_SIZE0: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_SIZE1: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_SIZE2: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_RBAR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF1_RBAR_NUM    : vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi1);
        PF1_REVISION_ID : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_BAR0_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_SRIOV_BAR0_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF1_SRIOV_BAR1_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_BAR1_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_SRIOV_BAR2_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_SRIOV_BAR2_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF1_SRIOV_BAR3_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_SRIOV_BAR3_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_SRIOV_BAR4_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_SRIOV_BAR4_CONTROL: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PF1_SRIOV_BAR5_APERTURE_SIZE: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1);
        PF1_SRIOV_BAR5_CONTROL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_SRIOV_CAP_INITIAL_VF: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_CAP_TOTAL_VF: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PF1_SRIOV_FIRST_VF_OFFSET: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_FUNC_DEP_LINK: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_SUPPORTED_PAGE_SIZE: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SRIOV_VF_DEVICE_ID: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_SUBSYSTEM_ID: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        PF1_TPHR_CAP_ENABLE: string  := "FALSE";
        PF1_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        PF1_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        PF1_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        PF1_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PF1_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        PL_DISABLE_EI_INFER_IN_L0: string  := "FALSE";
        PL_DISABLE_GEN3_DC_BALANCE: string  := "FALSE";
        PL_DISABLE_SCRAMBLING: string  := "FALSE";
        PL_DISABLE_UPCONFIG_CAPABLE: string  := "FALSE";
        PL_EQ_ADAPT_DISABLE_COEFF_CHECK: string  := "FALSE";
        PL_EQ_ADAPT_DISABLE_PRESET_CHECK: string  := "FALSE";
        PL_EQ_ADAPT_ITER_COUNT: vl_logic_vector(4 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi0);
        PL_EQ_ADAPT_REJECT_RETRY_COUNT: vl_logic_vector(1 downto 0) := (Hi0, Hi1);
        PL_EQ_BYPASS_PHASE23: string  := "FALSE";
        PL_EQ_SHORT_ADAPT_PHASE: string  := "FALSE";
        PL_LANE0_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE1_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE2_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE3_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE4_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE5_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE6_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LANE7_EQ_CONTROL: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PL_LINK_CAP_MAX_LINK_SPEED: vl_logic_vector(2 downto 0) := (Hi1, Hi0, Hi0);
        PL_LINK_CAP_MAX_LINK_WIDTH: vl_logic_vector(3 downto 0) := (Hi1, Hi0, Hi0, Hi0);
        PL_N_FTS_COMCLK_GEN1: integer := 255;
        PL_N_FTS_COMCLK_GEN2: integer := 255;
        PL_N_FTS_COMCLK_GEN3: integer := 255;
        PL_N_FTS_GEN1   : integer := 255;
        PL_N_FTS_GEN2   : integer := 255;
        PL_N_FTS_GEN3   : integer := 255;
        PL_SIM_FAST_LINK_TRAINING: string  := "FALSE";
        PL_UPSTREAM_FACING: string  := "TRUE";
        PM_ASPML0S_TIMEOUT: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi1, Hi1, Hi1, Hi0, Hi0);
        PM_ASPML1_ENTRY_DELAY: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PM_ENABLE_SLOT_POWER_CAPTURE: string  := "TRUE";
        PM_L1_REENTRY_DELAY: vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        PM_PME_SERVICE_TIMEOUT_DELAY: vl_logic_vector(19 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        PM_PME_TURNOFF_ACK_DELAY: vl_logic_vector(15 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi0, Hi0);
        SIM_VERSION     : string  := "1.0";
        SPARE_BIT0      : integer := 0;
        SPARE_BIT1      : integer := 0;
        SPARE_BIT2      : integer := 0;
        SPARE_BIT3      : integer := 0;
        SPARE_BIT4      : integer := 0;
        SPARE_BIT5      : integer := 0;
        SPARE_BIT6      : integer := 0;
        SPARE_BIT7      : integer := 0;
        SPARE_BIT8      : integer := 0;
        SPARE_BYTE0     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BYTE1     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BYTE2     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_BYTE3     : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD0     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD1     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD2     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SPARE_WORD3     : vl_logic_vector(31 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        SRIOV_CAP_ENABLE: string  := "FALSE";
        TL_COMPL_TIMEOUT_REG0: vl_logic_vector(23 downto 0) := (Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi1, Hi0, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        TL_COMPL_TIMEOUT_REG1: vl_logic_vector(27 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        TL_CREDITS_CD   : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi1, Hi1, Hi1, Hi1, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        TL_CREDITS_CH   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        TL_CREDITS_NPD  : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0);
        TL_CREDITS_NPH  : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        TL_CREDITS_PD   : vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi1, Hi1, Hi0, Hi0, Hi0);
        TL_CREDITS_PH   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0);
        TL_ENABLE_MESSAGE_RID_CHECK_ENABLE: string  := "TRUE";
        TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE: string  := "FALSE";
        TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE: string  := "FALSE";
        TL_LEGACY_MODE_ENABLE: string  := "FALSE";
        TL_PF_ENABLE_REG: string  := "FALSE";
        TL_TAG_MGMT_ENABLE: string  := "TRUE";
        VF0_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF0_CAPABILITY_POINTER: vl_logic_vector(7 downto 0) := (Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF0_MSIX_CAP_PBA_BIR: integer := 0;
        VF0_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF0_MSIX_CAP_TABLE_BIR: integer := 0;
        VF0_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF0_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF0_MSI_CAP_MULTIMSGCAP: integer := 0;
        VF0_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        VF0_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF0_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        VF0_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        VF0_TPHR_CAP_ENABLE: string  := "FALSE";
        VF0_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        VF0_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF0_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        VF0_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        VF0_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF0_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VF1_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF1_MSIX_CAP_PBA_BIR: integer := 0;
        VF1_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF1_MSIX_CAP_TABLE_BIR: integer := 0;
        VF1_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF1_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF1_MSI_CAP_MULTIMSGCAP: integer := 0;
        VF1_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        VF1_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF1_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        VF1_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        VF1_TPHR_CAP_ENABLE: string  := "FALSE";
        VF1_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        VF1_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF1_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        VF1_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        VF1_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF1_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VF2_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF2_MSIX_CAP_PBA_BIR: integer := 0;
        VF2_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF2_MSIX_CAP_TABLE_BIR: integer := 0;
        VF2_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF2_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF2_MSI_CAP_MULTIMSGCAP: integer := 0;
        VF2_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        VF2_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF2_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        VF2_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        VF2_TPHR_CAP_ENABLE: string  := "FALSE";
        VF2_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        VF2_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF2_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        VF2_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        VF2_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF2_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VF3_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF3_MSIX_CAP_PBA_BIR: integer := 0;
        VF3_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF3_MSIX_CAP_TABLE_BIR: integer := 0;
        VF3_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF3_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF3_MSI_CAP_MULTIMSGCAP: integer := 0;
        VF3_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        VF3_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF3_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        VF3_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        VF3_TPHR_CAP_ENABLE: string  := "FALSE";
        VF3_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        VF3_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF3_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        VF3_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        VF3_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF3_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VF4_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF4_MSIX_CAP_PBA_BIR: integer := 0;
        VF4_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF4_MSIX_CAP_TABLE_BIR: integer := 0;
        VF4_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF4_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF4_MSI_CAP_MULTIMSGCAP: integer := 0;
        VF4_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        VF4_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF4_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        VF4_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        VF4_TPHR_CAP_ENABLE: string  := "FALSE";
        VF4_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        VF4_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF4_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        VF4_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        VF4_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF4_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1);
        VF5_ARI_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF5_MSIX_CAP_PBA_BIR: integer := 0;
        VF5_MSIX_CAP_PBA_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0);
        VF5_MSIX_CAP_TABLE_BIR: integer := 0;
        VF5_MSIX_CAP_TABLE_OFFSET: vl_logic_vector(28 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF5_MSIX_CAP_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF5_MSI_CAP_MULTIMSGCAP: integer := 0;
        VF5_PM_CAP_ID   : vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi1);
        VF5_PM_CAP_NEXTPTR: vl_logic_vector(7 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF5_PM_CAP_VER_ID: vl_logic_vector(2 downto 0) := (Hi0, Hi1, Hi1);
        VF5_TPHR_CAP_DEV_SPECIFIC_MODE: string  := "TRUE";
        VF5_TPHR_CAP_ENABLE: string  := "FALSE";
        VF5_TPHR_CAP_INT_VEC_MODE: string  := "TRUE";
        VF5_TPHR_CAP_NEXTPTR: vl_logic_vector(11 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF5_TPHR_CAP_ST_MODE_SEL: vl_logic_vector(2 downto 0) := (Hi0, Hi0, Hi0);
        VF5_TPHR_CAP_ST_TABLE_LOC: vl_logic_vector(1 downto 0) := (Hi0, Hi0);
        VF5_TPHR_CAP_ST_TABLE_SIZE: vl_logic_vector(10 downto 0) := (Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0, Hi0);
        VF5_TPHR_CAP_VER: vl_logic_vector(3 downto 0) := (Hi0, Hi0, Hi0, Hi1)
    );
    port(
        CFGCURRENTSPEED : out    vl_logic_vector(2 downto 0);
        CFGDPASUBSTATECHANGE: out    vl_logic_vector(1 downto 0);
        CFGERRCOROUT    : out    vl_logic;
        CFGERRFATALOUT  : out    vl_logic;
        CFGERRNONFATALOUT: out    vl_logic;
        CFGEXTFUNCTIONNUMBER: out    vl_logic_vector(7 downto 0);
        CFGEXTREADRECEIVED: out    vl_logic;
        CFGEXTREGISTERNUMBER: out    vl_logic_vector(9 downto 0);
        CFGEXTWRITEBYTEENABLE: out    vl_logic_vector(3 downto 0);
        CFGEXTWRITEDATA : out    vl_logic_vector(31 downto 0);
        CFGEXTWRITERECEIVED: out    vl_logic;
        CFGFCCPLD       : out    vl_logic_vector(11 downto 0);
        CFGFCCPLH       : out    vl_logic_vector(7 downto 0);
        CFGFCNPD        : out    vl_logic_vector(11 downto 0);
        CFGFCNPH        : out    vl_logic_vector(7 downto 0);
        CFGFCPD         : out    vl_logic_vector(11 downto 0);
        CFGFCPH         : out    vl_logic_vector(7 downto 0);
        CFGFLRINPROCESS : out    vl_logic_vector(1 downto 0);
        CFGFUNCTIONPOWERSTATE: out    vl_logic_vector(5 downto 0);
        CFGFUNCTIONSTATUS: out    vl_logic_vector(7 downto 0);
        CFGHOTRESETOUT  : out    vl_logic;
        CFGINPUTUPDATEDONE: out    vl_logic;
        CFGINTERRUPTAOUTPUT: out    vl_logic;
        CFGINTERRUPTBOUTPUT: out    vl_logic;
        CFGINTERRUPTCOUTPUT: out    vl_logic;
        CFGINTERRUPTDOUTPUT: out    vl_logic;
        CFGINTERRUPTMSIDATA: out    vl_logic_vector(31 downto 0);
        CFGINTERRUPTMSIENABLE: out    vl_logic_vector(1 downto 0);
        CFGINTERRUPTMSIFAIL: out    vl_logic;
        CFGINTERRUPTMSIMASKUPDATE: out    vl_logic;
        CFGINTERRUPTMSIMMENABLE: out    vl_logic_vector(5 downto 0);
        CFGINTERRUPTMSISENT: out    vl_logic;
        CFGINTERRUPTMSIVFENABLE: out    vl_logic_vector(5 downto 0);
        CFGINTERRUPTMSIXENABLE: out    vl_logic_vector(1 downto 0);
        CFGINTERRUPTMSIXFAIL: out    vl_logic;
        CFGINTERRUPTMSIXMASK: out    vl_logic_vector(1 downto 0);
        CFGINTERRUPTMSIXSENT: out    vl_logic;
        CFGINTERRUPTMSIXVFENABLE: out    vl_logic_vector(5 downto 0);
        CFGINTERRUPTMSIXVFMASK: out    vl_logic_vector(5 downto 0);
        CFGINTERRUPTSENT: out    vl_logic;
        CFGLINKPOWERSTATE: out    vl_logic_vector(1 downto 0);
        CFGLOCALERROR   : out    vl_logic;
        CFGLTRENABLE    : out    vl_logic;
        CFGLTSSMSTATE   : out    vl_logic_vector(5 downto 0);
        CFGMAXPAYLOAD   : out    vl_logic_vector(2 downto 0);
        CFGMAXREADREQ   : out    vl_logic_vector(2 downto 0);
        CFGMCUPDATEDONE : out    vl_logic;
        CFGMGMTREADDATA : out    vl_logic_vector(31 downto 0);
        CFGMGMTREADWRITEDONE: out    vl_logic;
        CFGMSGRECEIVED  : out    vl_logic;
        CFGMSGRECEIVEDDATA: out    vl_logic_vector(7 downto 0);
        CFGMSGRECEIVEDTYPE: out    vl_logic_vector(4 downto 0);
        CFGMSGTRANSMITDONE: out    vl_logic;
        CFGNEGOTIATEDWIDTH: out    vl_logic_vector(3 downto 0);
        CFGOBFFENABLE   : out    vl_logic_vector(1 downto 0);
        CFGPERFUNCSTATUSDATA: out    vl_logic_vector(15 downto 0);
        CFGPERFUNCTIONUPDATEDONE: out    vl_logic;
        CFGPHYLINKDOWN  : out    vl_logic;
        CFGPHYLINKSTATUS: out    vl_logic_vector(1 downto 0);
        CFGPLSTATUSCHANGE: out    vl_logic;
        CFGPOWERSTATECHANGEINTERRUPT: out    vl_logic;
        CFGRCBSTATUS    : out    vl_logic_vector(1 downto 0);
        CFGTPHFUNCTIONNUM: out    vl_logic_vector(2 downto 0);
        CFGTPHREQUESTERENABLE: out    vl_logic_vector(1 downto 0);
        CFGTPHSTMODE    : out    vl_logic_vector(5 downto 0);
        CFGTPHSTTADDRESS: out    vl_logic_vector(4 downto 0);
        CFGTPHSTTREADENABLE: out    vl_logic;
        CFGTPHSTTWRITEBYTEVALID: out    vl_logic_vector(3 downto 0);
        CFGTPHSTTWRITEDATA: out    vl_logic_vector(31 downto 0);
        CFGTPHSTTWRITEENABLE: out    vl_logic;
        CFGVFFLRINPROCESS: out    vl_logic_vector(5 downto 0);
        CFGVFPOWERSTATE : out    vl_logic_vector(17 downto 0);
        CFGVFSTATUS     : out    vl_logic_vector(11 downto 0);
        CFGVFTPHREQUESTERENABLE: out    vl_logic_vector(5 downto 0);
        CFGVFTPHSTMODE  : out    vl_logic_vector(17 downto 0);
        DBGDATAOUT      : out    vl_logic_vector(15 downto 0);
        DRPDO           : out    vl_logic_vector(15 downto 0);
        DRPRDY          : out    vl_logic;
        MAXISCQTDATA    : out    vl_logic_vector(255 downto 0);
        MAXISCQTKEEP    : out    vl_logic_vector(7 downto 0);
        MAXISCQTLAST    : out    vl_logic;
        MAXISCQTUSER    : out    vl_logic_vector(84 downto 0);
        MAXISCQTVALID   : out    vl_logic;
        MAXISRCTDATA    : out    vl_logic_vector(255 downto 0);
        MAXISRCTKEEP    : out    vl_logic_vector(7 downto 0);
        MAXISRCTLAST    : out    vl_logic;
        MAXISRCTUSER    : out    vl_logic_vector(74 downto 0);
        MAXISRCTVALID   : out    vl_logic;
        MICOMPLETIONRAMREADADDRESSAL: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMREADADDRESSAU: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMREADADDRESSBL: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMREADADDRESSBU: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMREADENABLEL: out    vl_logic_vector(3 downto 0);
        MICOMPLETIONRAMREADENABLEU: out    vl_logic_vector(3 downto 0);
        MICOMPLETIONRAMWRITEADDRESSAL: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMWRITEADDRESSAU: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMWRITEADDRESSBL: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMWRITEADDRESSBU: out    vl_logic_vector(9 downto 0);
        MICOMPLETIONRAMWRITEDATAL: out    vl_logic_vector(71 downto 0);
        MICOMPLETIONRAMWRITEDATAU: out    vl_logic_vector(71 downto 0);
        MICOMPLETIONRAMWRITEENABLEL: out    vl_logic_vector(3 downto 0);
        MICOMPLETIONRAMWRITEENABLEU: out    vl_logic_vector(3 downto 0);
        MIREPLAYRAMADDRESS: out    vl_logic_vector(8 downto 0);
        MIREPLAYRAMREADENABLE: out    vl_logic_vector(1 downto 0);
        MIREPLAYRAMWRITEDATA: out    vl_logic_vector(143 downto 0);
        MIREPLAYRAMWRITEENABLE: out    vl_logic_vector(1 downto 0);
        MIREQUESTRAMREADADDRESSA: out    vl_logic_vector(8 downto 0);
        MIREQUESTRAMREADADDRESSB: out    vl_logic_vector(8 downto 0);
        MIREQUESTRAMREADENABLE: out    vl_logic_vector(3 downto 0);
        MIREQUESTRAMWRITEADDRESSA: out    vl_logic_vector(8 downto 0);
        MIREQUESTRAMWRITEADDRESSB: out    vl_logic_vector(8 downto 0);
        MIREQUESTRAMWRITEDATA: out    vl_logic_vector(143 downto 0);
        MIREQUESTRAMWRITEENABLE: out    vl_logic_vector(3 downto 0);
        PCIECQNPREQCOUNT: out    vl_logic_vector(5 downto 0);
        PCIERQSEQNUM    : out    vl_logic_vector(3 downto 0);
        PCIERQSEQNUMVLD : out    vl_logic;
        PCIERQTAG       : out    vl_logic_vector(5 downto 0);
        PCIERQTAGAV     : out    vl_logic_vector(1 downto 0);
        PCIERQTAGVLD    : out    vl_logic;
        PCIETFCNPDAV    : out    vl_logic_vector(1 downto 0);
        PCIETFCNPHAV    : out    vl_logic_vector(1 downto 0);
        PIPERX0EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX0EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX0EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX0EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX0POLARITY : out    vl_logic;
        PIPERX1EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX1EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX1EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX1EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX1POLARITY : out    vl_logic;
        PIPERX2EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX2EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX2EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX2EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX2POLARITY : out    vl_logic;
        PIPERX3EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX3EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX3EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX3EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX3POLARITY : out    vl_logic;
        PIPERX4EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX4EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX4EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX4EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX4POLARITY : out    vl_logic;
        PIPERX5EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX5EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX5EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX5EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX5POLARITY : out    vl_logic;
        PIPERX6EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX6EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX6EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX6EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX6POLARITY : out    vl_logic;
        PIPERX7EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPERX7EQLPLFFS : out    vl_logic_vector(5 downto 0);
        PIPERX7EQLPTXPRESET: out    vl_logic_vector(3 downto 0);
        PIPERX7EQPRESET : out    vl_logic_vector(2 downto 0);
        PIPERX7POLARITY : out    vl_logic;
        PIPETX0CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX0COMPLIANCE: out    vl_logic;
        PIPETX0DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX0DATAVALID: out    vl_logic;
        PIPETX0ELECIDLE : out    vl_logic;
        PIPETX0EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX0EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX0EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX0POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX0STARTBLOCK: out    vl_logic;
        PIPETX0SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX1CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX1COMPLIANCE: out    vl_logic;
        PIPETX1DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX1DATAVALID: out    vl_logic;
        PIPETX1ELECIDLE : out    vl_logic;
        PIPETX1EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX1EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX1EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX1POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX1STARTBLOCK: out    vl_logic;
        PIPETX1SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX2CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX2COMPLIANCE: out    vl_logic;
        PIPETX2DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX2DATAVALID: out    vl_logic;
        PIPETX2ELECIDLE : out    vl_logic;
        PIPETX2EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX2EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX2EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX2POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX2STARTBLOCK: out    vl_logic;
        PIPETX2SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX3CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX3COMPLIANCE: out    vl_logic;
        PIPETX3DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX3DATAVALID: out    vl_logic;
        PIPETX3ELECIDLE : out    vl_logic;
        PIPETX3EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX3EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX3EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX3POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX3STARTBLOCK: out    vl_logic;
        PIPETX3SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX4CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX4COMPLIANCE: out    vl_logic;
        PIPETX4DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX4DATAVALID: out    vl_logic;
        PIPETX4ELECIDLE : out    vl_logic;
        PIPETX4EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX4EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX4EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX4POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX4STARTBLOCK: out    vl_logic;
        PIPETX4SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX5CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX5COMPLIANCE: out    vl_logic;
        PIPETX5DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX5DATAVALID: out    vl_logic;
        PIPETX5ELECIDLE : out    vl_logic;
        PIPETX5EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX5EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX5EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX5POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX5STARTBLOCK: out    vl_logic;
        PIPETX5SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX6CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX6COMPLIANCE: out    vl_logic;
        PIPETX6DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX6DATAVALID: out    vl_logic;
        PIPETX6ELECIDLE : out    vl_logic;
        PIPETX6EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX6EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX6EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX6POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX6STARTBLOCK: out    vl_logic;
        PIPETX6SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETX7CHARISK  : out    vl_logic_vector(1 downto 0);
        PIPETX7COMPLIANCE: out    vl_logic;
        PIPETX7DATA     : out    vl_logic_vector(31 downto 0);
        PIPETX7DATAVALID: out    vl_logic;
        PIPETX7ELECIDLE : out    vl_logic;
        PIPETX7EQCONTROL: out    vl_logic_vector(1 downto 0);
        PIPETX7EQDEEMPH : out    vl_logic_vector(5 downto 0);
        PIPETX7EQPRESET : out    vl_logic_vector(3 downto 0);
        PIPETX7POWERDOWN: out    vl_logic_vector(1 downto 0);
        PIPETX7STARTBLOCK: out    vl_logic;
        PIPETX7SYNCHEADER: out    vl_logic_vector(1 downto 0);
        PIPETXDEEMPH    : out    vl_logic;
        PIPETXMARGIN    : out    vl_logic_vector(2 downto 0);
        PIPETXRATE      : out    vl_logic_vector(1 downto 0);
        PIPETXRCVRDET   : out    vl_logic;
        PIPETXRESET     : out    vl_logic;
        PIPETXSWING     : out    vl_logic;
        PLEQINPROGRESS  : out    vl_logic;
        PLEQPHASE       : out    vl_logic_vector(1 downto 0);
        PLGEN3PCSRXSLIDE: out    vl_logic_vector(7 downto 0);
        SAXISCCTREADY   : out    vl_logic_vector(3 downto 0);
        SAXISRQTREADY   : out    vl_logic_vector(3 downto 0);
        CFGCONFIGSPACEENABLE: in     vl_logic;
        CFGDEVID        : in     vl_logic_vector(15 downto 0);
        CFGDSBUSNUMBER  : in     vl_logic_vector(7 downto 0);
        CFGDSDEVICENUMBER: in     vl_logic_vector(4 downto 0);
        CFGDSFUNCTIONNUMBER: in     vl_logic_vector(2 downto 0);
        CFGDSN          : in     vl_logic_vector(63 downto 0);
        CFGDSPORTNUMBER : in     vl_logic_vector(7 downto 0);
        CFGERRCORIN     : in     vl_logic;
        CFGERRUNCORIN   : in     vl_logic;
        CFGEXTREADDATA  : in     vl_logic_vector(31 downto 0);
        CFGEXTREADDATAVALID: in     vl_logic;
        CFGFCSEL        : in     vl_logic_vector(2 downto 0);
        CFGFLRDONE      : in     vl_logic_vector(1 downto 0);
        CFGHOTRESETIN   : in     vl_logic;
        CFGINPUTUPDATEREQUEST: in     vl_logic;
        CFGINTERRUPTINT : in     vl_logic_vector(3 downto 0);
        CFGINTERRUPTMSIATTR: in     vl_logic_vector(2 downto 0);
        CFGINTERRUPTMSIFUNCTIONNUMBER: in     vl_logic_vector(2 downto 0);
        CFGINTERRUPTMSIINT: in     vl_logic_vector(31 downto 0);
        CFGINTERRUPTMSIPENDINGSTATUS: in     vl_logic_vector(63 downto 0);
        CFGINTERRUPTMSISELECT: in     vl_logic_vector(3 downto 0);
        CFGINTERRUPTMSITPHPRESENT: in     vl_logic;
        CFGINTERRUPTMSITPHSTTAG: in     vl_logic_vector(8 downto 0);
        CFGINTERRUPTMSITPHTYPE: in     vl_logic_vector(1 downto 0);
        CFGINTERRUPTMSIXADDRESS: in     vl_logic_vector(63 downto 0);
        CFGINTERRUPTMSIXDATA: in     vl_logic_vector(31 downto 0);
        CFGINTERRUPTMSIXINT: in     vl_logic;
        CFGINTERRUPTPENDING: in     vl_logic_vector(1 downto 0);
        CFGLINKTRAININGENABLE: in     vl_logic;
        CFGMCUPDATEREQUEST: in     vl_logic;
        CFGMGMTADDR     : in     vl_logic_vector(18 downto 0);
        CFGMGMTBYTEENABLE: in     vl_logic_vector(3 downto 0);
        CFGMGMTREAD     : in     vl_logic;
        CFGMGMTTYPE1CFGREGACCESS: in     vl_logic;
        CFGMGMTWRITE    : in     vl_logic;
        CFGMGMTWRITEDATA: in     vl_logic_vector(31 downto 0);
        CFGMSGTRANSMIT  : in     vl_logic;
        CFGMSGTRANSMITDATA: in     vl_logic_vector(31 downto 0);
        CFGMSGTRANSMITTYPE: in     vl_logic_vector(2 downto 0);
        CFGPERFUNCSTATUSCONTROL: in     vl_logic_vector(2 downto 0);
        CFGPERFUNCTIONNUMBER: in     vl_logic_vector(2 downto 0);
        CFGPERFUNCTIONOUTPUTREQUEST: in     vl_logic;
        CFGPOWERSTATECHANGEACK: in     vl_logic;
        CFGREQPMTRANSITIONL23READY: in     vl_logic;
        CFGREVID        : in     vl_logic_vector(7 downto 0);
        CFGSUBSYSID     : in     vl_logic_vector(15 downto 0);
        CFGSUBSYSVENDID : in     vl_logic_vector(15 downto 0);
        CFGTPHSTTREADDATA: in     vl_logic_vector(31 downto 0);
        CFGTPHSTTREADDATAVALID: in     vl_logic;
        CFGVENDID       : in     vl_logic_vector(15 downto 0);
        CFGVFFLRDONE    : in     vl_logic_vector(5 downto 0);
        CORECLK         : in     vl_logic;
        CORECLKMICOMPLETIONRAML: in     vl_logic;
        CORECLKMICOMPLETIONRAMU: in     vl_logic;
        CORECLKMIREPLAYRAM: in     vl_logic;
        CORECLKMIREQUESTRAM: in     vl_logic;
        DRPADDR         : in     vl_logic_vector(10 downto 0);
        DRPCLK          : in     vl_logic;
        DRPDI           : in     vl_logic_vector(15 downto 0);
        DRPEN           : in     vl_logic;
        DRPWE           : in     vl_logic;
        MAXISCQTREADY   : in     vl_logic_vector(21 downto 0);
        MAXISRCTREADY   : in     vl_logic_vector(21 downto 0);
        MGMTRESETN      : in     vl_logic;
        MGMTSTICKYRESETN: in     vl_logic;
        MICOMPLETIONRAMREADDATA: in     vl_logic_vector(143 downto 0);
        MIREPLAYRAMREADDATA: in     vl_logic_vector(143 downto 0);
        MIREQUESTRAMREADDATA: in     vl_logic_vector(143 downto 0);
        PCIECQNPREQ     : in     vl_logic;
        PIPECLK         : in     vl_logic;
        PIPEEQFS        : in     vl_logic_vector(5 downto 0);
        PIPEEQLF        : in     vl_logic_vector(5 downto 0);
        PIPERESETN      : in     vl_logic;
        PIPERX0CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX0DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX0DATAVALID: in     vl_logic;
        PIPERX0ELECIDLE : in     vl_logic;
        PIPERX0EQDONE   : in     vl_logic;
        PIPERX0EQLPADAPTDONE: in     vl_logic;
        PIPERX0EQLPLFFSSEL: in     vl_logic;
        PIPERX0EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX0PHYSTATUS: in     vl_logic;
        PIPERX0STARTBLOCK: in     vl_logic;
        PIPERX0STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX0SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX0VALID    : in     vl_logic;
        PIPERX1CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX1DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX1DATAVALID: in     vl_logic;
        PIPERX1ELECIDLE : in     vl_logic;
        PIPERX1EQDONE   : in     vl_logic;
        PIPERX1EQLPADAPTDONE: in     vl_logic;
        PIPERX1EQLPLFFSSEL: in     vl_logic;
        PIPERX1EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX1PHYSTATUS: in     vl_logic;
        PIPERX1STARTBLOCK: in     vl_logic;
        PIPERX1STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX1SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX1VALID    : in     vl_logic;
        PIPERX2CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX2DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX2DATAVALID: in     vl_logic;
        PIPERX2ELECIDLE : in     vl_logic;
        PIPERX2EQDONE   : in     vl_logic;
        PIPERX2EQLPADAPTDONE: in     vl_logic;
        PIPERX2EQLPLFFSSEL: in     vl_logic;
        PIPERX2EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX2PHYSTATUS: in     vl_logic;
        PIPERX2STARTBLOCK: in     vl_logic;
        PIPERX2STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX2SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX2VALID    : in     vl_logic;
        PIPERX3CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX3DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX3DATAVALID: in     vl_logic;
        PIPERX3ELECIDLE : in     vl_logic;
        PIPERX3EQDONE   : in     vl_logic;
        PIPERX3EQLPADAPTDONE: in     vl_logic;
        PIPERX3EQLPLFFSSEL: in     vl_logic;
        PIPERX3EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX3PHYSTATUS: in     vl_logic;
        PIPERX3STARTBLOCK: in     vl_logic;
        PIPERX3STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX3SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX3VALID    : in     vl_logic;
        PIPERX4CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX4DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX4DATAVALID: in     vl_logic;
        PIPERX4ELECIDLE : in     vl_logic;
        PIPERX4EQDONE   : in     vl_logic;
        PIPERX4EQLPADAPTDONE: in     vl_logic;
        PIPERX4EQLPLFFSSEL: in     vl_logic;
        PIPERX4EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX4PHYSTATUS: in     vl_logic;
        PIPERX4STARTBLOCK: in     vl_logic;
        PIPERX4STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX4SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX4VALID    : in     vl_logic;
        PIPERX5CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX5DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX5DATAVALID: in     vl_logic;
        PIPERX5ELECIDLE : in     vl_logic;
        PIPERX5EQDONE   : in     vl_logic;
        PIPERX5EQLPADAPTDONE: in     vl_logic;
        PIPERX5EQLPLFFSSEL: in     vl_logic;
        PIPERX5EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX5PHYSTATUS: in     vl_logic;
        PIPERX5STARTBLOCK: in     vl_logic;
        PIPERX5STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX5SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX5VALID    : in     vl_logic;
        PIPERX6CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX6DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX6DATAVALID: in     vl_logic;
        PIPERX6ELECIDLE : in     vl_logic;
        PIPERX6EQDONE   : in     vl_logic;
        PIPERX6EQLPADAPTDONE: in     vl_logic;
        PIPERX6EQLPLFFSSEL: in     vl_logic;
        PIPERX6EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX6PHYSTATUS: in     vl_logic;
        PIPERX6STARTBLOCK: in     vl_logic;
        PIPERX6STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX6SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX6VALID    : in     vl_logic;
        PIPERX7CHARISK  : in     vl_logic_vector(1 downto 0);
        PIPERX7DATA     : in     vl_logic_vector(31 downto 0);
        PIPERX7DATAVALID: in     vl_logic;
        PIPERX7ELECIDLE : in     vl_logic;
        PIPERX7EQDONE   : in     vl_logic;
        PIPERX7EQLPADAPTDONE: in     vl_logic;
        PIPERX7EQLPLFFSSEL: in     vl_logic;
        PIPERX7EQLPNEWTXCOEFFORPRESET: in     vl_logic_vector(17 downto 0);
        PIPERX7PHYSTATUS: in     vl_logic;
        PIPERX7STARTBLOCK: in     vl_logic;
        PIPERX7STATUS   : in     vl_logic_vector(2 downto 0);
        PIPERX7SYNCHEADER: in     vl_logic_vector(1 downto 0);
        PIPERX7VALID    : in     vl_logic;
        PIPETX0EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX0EQDONE   : in     vl_logic;
        PIPETX1EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX1EQDONE   : in     vl_logic;
        PIPETX2EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX2EQDONE   : in     vl_logic;
        PIPETX3EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX3EQDONE   : in     vl_logic;
        PIPETX4EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX4EQDONE   : in     vl_logic;
        PIPETX5EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX5EQDONE   : in     vl_logic;
        PIPETX6EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX6EQDONE   : in     vl_logic;
        PIPETX7EQCOEFF  : in     vl_logic_vector(17 downto 0);
        PIPETX7EQDONE   : in     vl_logic;
        PLDISABLESCRAMBLER: in     vl_logic;
        PLEQRESETEIEOSCOUNT: in     vl_logic;
        PLGEN3PCSDISABLE: in     vl_logic;
        PLGEN3PCSRXSYNCDONE: in     vl_logic_vector(7 downto 0);
        RECCLK          : in     vl_logic;
        RESETN          : in     vl_logic;
        SAXISCCTDATA    : in     vl_logic_vector(255 downto 0);
        SAXISCCTKEEP    : in     vl_logic_vector(7 downto 0);
        SAXISCCTLAST    : in     vl_logic;
        SAXISCCTUSER    : in     vl_logic_vector(32 downto 0);
        SAXISCCTVALID   : in     vl_logic;
        SAXISRQTDATA    : in     vl_logic_vector(255 downto 0);
        SAXISRQTKEEP    : in     vl_logic_vector(7 downto 0);
        SAXISRQTLAST    : in     vl_logic;
        SAXISRQTUSER    : in     vl_logic_vector(59 downto 0);
        SAXISRQTVALID   : in     vl_logic;
        USERCLK         : in     vl_logic
    );
    attribute mti_svvh_generic_type : integer;
    attribute mti_svvh_generic_type of LOC : constant is 1;
    attribute mti_svvh_generic_type of ARI_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_CC_ALIGNMENT_MODE : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_CC_PARITY_CHK : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_CQ_ALIGNMENT_MODE : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_ENABLE_CLIENT_TAG : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_ENABLE_MSG_ROUTE : constant is 2;
    attribute mti_svvh_generic_type of AXISTEN_IF_ENABLE_RX_MSG_INTFC : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_RC_ALIGNMENT_MODE : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_RC_STRADDLE : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_RQ_ALIGNMENT_MODE : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_RQ_PARITY_CHK : constant is 1;
    attribute mti_svvh_generic_type of AXISTEN_IF_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of CRM_CORE_CLK_FREQ_500 : constant is 1;
    attribute mti_svvh_generic_type of CRM_USER_CLK_FREQ : constant is 2;
    attribute mti_svvh_generic_type of DNSTREAM_LINK_NUM : constant is 2;
    attribute mti_svvh_generic_type of GEN3_PCS_AUTO_REALIGN : constant is 2;
    attribute mti_svvh_generic_type of GEN3_PCS_RX_ELECIDLE_INTERNAL : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT : constant is 2;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of LL_ACK_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of LL_CPL_FC_UPDATE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of LL_CPL_FC_UPDATE_TIMER_OVERRIDE : constant is 1;
    attribute mti_svvh_generic_type of LL_FC_UPDATE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of LL_FC_UPDATE_TIMER_OVERRIDE : constant is 1;
    attribute mti_svvh_generic_type of LL_NP_FC_UPDATE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of LL_NP_FC_UPDATE_TIMER_OVERRIDE : constant is 1;
    attribute mti_svvh_generic_type of LL_P_FC_UPDATE_TIMER : constant is 2;
    attribute mti_svvh_generic_type of LL_P_FC_UPDATE_TIMER_OVERRIDE : constant is 1;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT : constant is 2;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT_EN : constant is 1;
    attribute mti_svvh_generic_type of LL_REPLAY_TIMEOUT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of LTR_TX_MESSAGE_MINIMUM_INTERVAL : constant is 2;
    attribute mti_svvh_generic_type of LTR_TX_MESSAGE_ON_FUNC_POWER_STATE_CHANGE : constant is 1;
    attribute mti_svvh_generic_type of LTR_TX_MESSAGE_ON_LTR_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_AER_CAP_ECRC_CHECK_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_AER_CAP_ECRC_GEN_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_AER_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_ARI_CAP_NEXT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of PF0_ARI_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR0_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR0_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR1_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR1_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR2_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR2_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR3_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR3_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR4_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR4_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR5_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_BAR5_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_BIST_REGISTER : constant is 2;
    attribute mti_svvh_generic_type of PF0_CAPABILITY_POINTER : constant is 2;
    attribute mti_svvh_generic_type of PF0_CLASS_CODE : constant is 2;
    attribute mti_svvh_generic_type of PF0_DEVICE_ID : constant is 2;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_128B_CAS_ATOMIC_COMPLETER_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_32B_ATOMIC_COMPLETER_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_64B_ATOMIC_COMPLETER_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_CPL_TIMEOUT_DISABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_LTR_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_OBFF_SUPPORT : constant is 2;
    attribute mti_svvh_generic_type of PF0_DEV_CAP2_TPH_COMPLETER_SUPPORT : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP_ENDPOINT_L0S_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of PF0_DEV_CAP_ENDPOINT_L1_LATENCY : constant is 2;
    attribute mti_svvh_generic_type of PF0_DEV_CAP_EXT_TAG_SUPPORTED : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP_FUNCTION_LEVEL_RESET_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_DEV_CAP_MAX_PAYLOAD_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_CONTROL_EN : constant is 1;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 : constant is 2;
    attribute mti_svvh_generic_type of PF0_DPA_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_DSN_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_EXPANSION_ROM_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_EXPANSION_ROM_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_INTERRUPT_LINE : constant is 2;
    attribute mti_svvh_generic_type of PF0_INTERRUPT_PIN : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_ASPM_SUPPORT : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L0S_EXIT_LATENCY_COMCLK_GEN3 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L0S_EXIT_LATENCY_GEN3 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L1_EXIT_LATENCY_COMCLK_GEN3 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L1_EXIT_LATENCY_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L1_EXIT_LATENCY_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_CAP_L1_EXIT_LATENCY_GEN3 : constant is 2;
    attribute mti_svvh_generic_type of PF0_LINK_STATUS_SLOT_CLOCK_CONFIG : constant is 1;
    attribute mti_svvh_generic_type of PF0_LTR_CAP_MAX_NOSNOOP_LAT : constant is 2;
    attribute mti_svvh_generic_type of PF0_LTR_CAP_MAX_SNOOP_LAT : constant is 2;
    attribute mti_svvh_generic_type of PF0_LTR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_LTR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSIX_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of PF0_MSI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_PB_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_PB_CAP_SYSTEM_ALLOCATED : constant is 1;
    attribute mti_svvh_generic_type of PF0_PB_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of PF0_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_PM_CAP_PMESUPPORT_D0 : constant is 1;
    attribute mti_svvh_generic_type of PF0_PM_CAP_PMESUPPORT_D1 : constant is 1;
    attribute mti_svvh_generic_type of PF0_PM_CAP_PMESUPPORT_D3HOT : constant is 1;
    attribute mti_svvh_generic_type of PF0_PM_CAP_SUPP_D1_STATE : constant is 1;
    attribute mti_svvh_generic_type of PF0_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of PF0_PM_CSR_NOSOFTRESET : constant is 1;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_INDEX0 : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_INDEX1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_INDEX2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_SIZE0 : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_SIZE1 : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_SIZE2 : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_RBAR_NUM : constant is 2;
    attribute mti_svvh_generic_type of PF0_REVISION_ID : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR0_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR0_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR1_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR1_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR2_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR2_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR3_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR3_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR4_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR4_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR5_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_BAR5_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_CAP_INITIAL_VF : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_CAP_TOTAL_VF : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_FIRST_VF_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_FUNC_DEP_LINK : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_SUPPORTED_PAGE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_SRIOV_VF_DEVICE_ID : constant is 2;
    attribute mti_svvh_generic_type of PF0_SUBSYSTEM_ID : constant is 2;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF0_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF0_VC_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF0_VC_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF1_AER_CAP_ECRC_CHECK_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of PF1_AER_CAP_ECRC_GEN_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of PF1_AER_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_ARI_CAP_NEXT_FUNC : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR0_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR0_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR1_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR1_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR2_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR2_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR3_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR3_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR4_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR4_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR5_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_BAR5_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_BIST_REGISTER : constant is 2;
    attribute mti_svvh_generic_type of PF1_CAPABILITY_POINTER : constant is 2;
    attribute mti_svvh_generic_type of PF1_CLASS_CODE : constant is 2;
    attribute mti_svvh_generic_type of PF1_DEVICE_ID : constant is 2;
    attribute mti_svvh_generic_type of PF1_DEV_CAP_MAX_PAYLOAD_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_CONTROL_EN : constant is 1;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION0 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION1 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION2 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION3 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION4 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION5 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION6 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_SUB_STATE_POWER_ALLOCATION7 : constant is 2;
    attribute mti_svvh_generic_type of PF1_DPA_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF1_DSN_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_EXPANSION_ROM_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_EXPANSION_ROM_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF1_INTERRUPT_LINE : constant is 2;
    attribute mti_svvh_generic_type of PF1_INTERRUPT_PIN : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSIX_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of PF1_MSI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_PB_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_PB_CAP_SYSTEM_ALLOCATED : constant is 1;
    attribute mti_svvh_generic_type of PF1_PB_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF1_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of PF1_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_INDEX0 : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_INDEX1 : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_INDEX2 : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_SIZE0 : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_SIZE1 : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_SIZE2 : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF1_RBAR_NUM : constant is 2;
    attribute mti_svvh_generic_type of PF1_REVISION_ID : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR0_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR0_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR1_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR1_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR2_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR2_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR3_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR3_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR4_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR4_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR5_APERTURE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_BAR5_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_CAP_INITIAL_VF : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_CAP_TOTAL_VF : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_FIRST_VF_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_FUNC_DEP_LINK : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_SUPPORTED_PAGE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_SRIOV_VF_DEVICE_ID : constant is 2;
    attribute mti_svvh_generic_type of PF1_SUBSYSTEM_ID : constant is 2;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of PF1_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of PL_DISABLE_EI_INFER_IN_L0 : constant is 1;
    attribute mti_svvh_generic_type of PL_DISABLE_GEN3_DC_BALANCE : constant is 1;
    attribute mti_svvh_generic_type of PL_DISABLE_SCRAMBLING : constant is 1;
    attribute mti_svvh_generic_type of PL_DISABLE_UPCONFIG_CAPABLE : constant is 1;
    attribute mti_svvh_generic_type of PL_EQ_ADAPT_DISABLE_COEFF_CHECK : constant is 1;
    attribute mti_svvh_generic_type of PL_EQ_ADAPT_DISABLE_PRESET_CHECK : constant is 1;
    attribute mti_svvh_generic_type of PL_EQ_ADAPT_ITER_COUNT : constant is 2;
    attribute mti_svvh_generic_type of PL_EQ_ADAPT_REJECT_RETRY_COUNT : constant is 2;
    attribute mti_svvh_generic_type of PL_EQ_BYPASS_PHASE23 : constant is 1;
    attribute mti_svvh_generic_type of PL_EQ_SHORT_ADAPT_PHASE : constant is 1;
    attribute mti_svvh_generic_type of PL_LANE0_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE1_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE2_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE3_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE4_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE5_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE6_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LANE7_EQ_CONTROL : constant is 2;
    attribute mti_svvh_generic_type of PL_LINK_CAP_MAX_LINK_SPEED : constant is 2;
    attribute mti_svvh_generic_type of PL_LINK_CAP_MAX_LINK_WIDTH : constant is 2;
    attribute mti_svvh_generic_type of PL_N_FTS_COMCLK_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of PL_N_FTS_COMCLK_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PL_N_FTS_COMCLK_GEN3 : constant is 2;
    attribute mti_svvh_generic_type of PL_N_FTS_GEN1 : constant is 2;
    attribute mti_svvh_generic_type of PL_N_FTS_GEN2 : constant is 2;
    attribute mti_svvh_generic_type of PL_N_FTS_GEN3 : constant is 2;
    attribute mti_svvh_generic_type of PL_SIM_FAST_LINK_TRAINING : constant is 1;
    attribute mti_svvh_generic_type of PL_UPSTREAM_FACING : constant is 1;
    attribute mti_svvh_generic_type of PM_ASPML0S_TIMEOUT : constant is 2;
    attribute mti_svvh_generic_type of PM_ASPML1_ENTRY_DELAY : constant is 2;
    attribute mti_svvh_generic_type of PM_ENABLE_SLOT_POWER_CAPTURE : constant is 1;
    attribute mti_svvh_generic_type of PM_L1_REENTRY_DELAY : constant is 2;
    attribute mti_svvh_generic_type of PM_PME_SERVICE_TIMEOUT_DELAY : constant is 2;
    attribute mti_svvh_generic_type of PM_PME_TURNOFF_ACK_DELAY : constant is 2;
    attribute mti_svvh_generic_type of SIM_VERSION : constant is 1;
    attribute mti_svvh_generic_type of SPARE_BIT0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT3 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT4 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT5 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT6 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT7 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BIT8 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_BYTE3 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD0 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD1 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD2 : constant is 2;
    attribute mti_svvh_generic_type of SPARE_WORD3 : constant is 2;
    attribute mti_svvh_generic_type of SRIOV_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_COMPL_TIMEOUT_REG0 : constant is 2;
    attribute mti_svvh_generic_type of TL_COMPL_TIMEOUT_REG1 : constant is 2;
    attribute mti_svvh_generic_type of TL_CREDITS_CD : constant is 2;
    attribute mti_svvh_generic_type of TL_CREDITS_CH : constant is 2;
    attribute mti_svvh_generic_type of TL_CREDITS_NPD : constant is 2;
    attribute mti_svvh_generic_type of TL_CREDITS_NPH : constant is 2;
    attribute mti_svvh_generic_type of TL_CREDITS_PD : constant is 2;
    attribute mti_svvh_generic_type of TL_CREDITS_PH : constant is 2;
    attribute mti_svvh_generic_type of TL_ENABLE_MESSAGE_RID_CHECK_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_EXTENDED_CFG_EXTEND_INTERFACE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_LEGACY_CFG_EXTEND_INTERFACE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_LEGACY_MODE_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of TL_PF_ENABLE_REG : constant is 1;
    attribute mti_svvh_generic_type of TL_TAG_MGMT_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF0_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF0_CAPABILITY_POINTER : constant is 2;
    attribute mti_svvh_generic_type of VF0_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF0_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF0_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF0_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF0_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF0_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of VF0_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VF0_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF0_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF0_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of VF1_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF1_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF1_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF1_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF1_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF1_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF1_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of VF1_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VF1_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF1_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF1_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of VF2_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF2_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF2_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF2_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF2_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF2_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF2_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of VF2_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VF2_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF2_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF2_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of VF3_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF3_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF3_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF3_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF3_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF3_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF3_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of VF3_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VF3_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF3_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF3_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of VF4_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF4_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF4_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF4_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF4_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF4_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF4_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of VF4_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VF4_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF4_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF4_TPHR_CAP_VER : constant is 2;
    attribute mti_svvh_generic_type of VF5_ARI_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF5_MSIX_CAP_PBA_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF5_MSIX_CAP_PBA_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF5_MSIX_CAP_TABLE_BIR : constant is 2;
    attribute mti_svvh_generic_type of VF5_MSIX_CAP_TABLE_OFFSET : constant is 2;
    attribute mti_svvh_generic_type of VF5_MSIX_CAP_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF5_MSI_CAP_MULTIMSGCAP : constant is 2;
    attribute mti_svvh_generic_type of VF5_PM_CAP_ID : constant is 2;
    attribute mti_svvh_generic_type of VF5_PM_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF5_PM_CAP_VER_ID : constant is 2;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_DEV_SPECIFIC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_ENABLE : constant is 1;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_INT_VEC_MODE : constant is 1;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_NEXTPTR : constant is 2;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_ST_MODE_SEL : constant is 2;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_ST_TABLE_LOC : constant is 2;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_ST_TABLE_SIZE : constant is 2;
    attribute mti_svvh_generic_type of VF5_TPHR_CAP_VER : constant is 2;
end X_PCIE_3_0;
