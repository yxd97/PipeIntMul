`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BKnB+QZ+biKdmQZTdowkR23sFRY0KBga1vxy8cUhxQ//6Y+CY0P5b+BGFjpmCd4p
m82JKDfkr8EZxK/X5RN9lCiwoOE1AXs+GK4E6enb482gTwGaWeT5j1LF1m4V2xRw
UX3sdIHk4VQMm6lmMKjafPcVbtY+LLNlrxFHvOizLT7Ej8RH/eKekhCAMrdpKsYU
2IHlEe2+7p1apZHEMZUd6tRklJ+3aiglT/TCBVc0xrjs3I3TTO4sIaqco6PHpkbT
sIa4LgIgozM0ICPYUvX7Q+onIy/bkyrcKO4NpfYcQKE+ulluyQrMVC1Kx9XfP8Qg
mTWztPPkcB69LUoxbOYVr26FXusINEcPz5qBDvfCcxxdCGOElPfnnrfEupVgn5AH
Z2jtKqb0FtZIlVBte/QyNxPRLaNmiYM6bJnIoF+EUdrSHokJNXtUbUsBIifauKW5
IlilaTPie4u2WU6GqEXaED7qK3HemofTXT5qszXa/RXm51Ao9+XsdeyfyDE2EJYn
RWy8dnpUT7VkZGuxLHmZ5kjl5j+B5vhjbcwcJ5yWUK6P86BiPSqVHCiHAaS9wUoU
TgyECxWMi9ubFE7W+jeKKqS0pTFs3TuDnagdPwIYYp2SepM+ZnAYgI2+UnofNpCi
nyN9zVrBC6Cy+h1fN37bsEaXJLxkFjqFLWOWad7PQXAh6EkqzkzUf76jaQ0Z5zdV
XYelBU+lBj27Wz1j5YH0HjtHiwsO4QMKrEf6oRJqXfYIXh7aUrNjIy72YR65vRU4
TYBUypXGzuytd8xhlynNrw==
`protect END_PROTECTED
