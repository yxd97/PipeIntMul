`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xeCJDAUarb+sEepyXtwOcuHMPG+DEDOgYnNI/RZroHfvdBMNiGXNo4Ovz/KUwDcv
pv49vle2EcmFO+wJu7i2ETIg0tvLAEb54anEIfdNfw+YPONvsOMiHdx4rsYLUUAJ
Hk6nMLj8VG+mgd0mI0C2hpCiD/q1whPPCxZbQtXa4CP6sqAaaOJB/ETBY+nQZm1J
7L784nBWj7X7SU0kLNZ1AKlTlN8w10zN8/lD7m6Zf4dTBbTfbYUwV8AumioKmB3p
oAtJ6TtfpJKM1LZA+RG5c7aUmBawCxJp0BK7p7Il+34uym7sY0tvfyTM6lKToUAN
2OwwzEeC4PfGENJNxtJXAYTYupPmw/dmrMOGyJLdFFFzN3T/uZWH0CdLFa9SmVvK
NEqUzb9lsd4YtMGk2vrLF8uG2evSJjifRdwYnfjUkbbI8em8FlvTXbRjuY1BZ0VR
NV7cS+ndDhLXUz8aadKRPxfUAi6ZFDIWty3Fqk6YGP+43oCSdESXqNOx26lnoD7c
to+HoTS8itnxPIAxoqsfEkfZTrBNrSQCvpW7GUuZUFGGIftFS1DRvQ0+0X3py73k
r968SySn/DQ+fAIad/TTHsRWAYtsfdqycdTBf/dFExWdDprOKO385iUVLVDCrhNO
O4AdJHuUGpNYzjuGTFmP5NNour2qR37eUKLG+0wH/70NTX+lBpWzxSjN7+NVhG3W
5fOXehPUFCXIv3qxuBemZ+Y0S/JoXdn+CZ+SHVsI1LLtgiDBH3rSqVqMbAsfEbhG
t679vBi9YhXMUeoA6XyRS0uTaaqh7d1lEFNTbNxFAKNNWOrlJUOYGdgXXU9/gPM7
BYx8/76ps/vPNbrOSrcNGHoFrZ2iTISUl4WUhb4QMB9goImR9wpXcsHtuM5MHTrN
bv1anY9ghColZ2rQva1OQ9fSQp+1YHSiKY/GELlwLdjWSxu0ZGxkAS6tj8+x3EEE
NU7ISHC7NBWoRBX/tRqq0WsiEvUlIKeCebCbgz3H8S1La7l17iRjrqQbJUjnYOet
kdgnt6tupfoIyE/qFhJN6j7UvypiKEt9opeHELTaOciKLGaHzTTqnm+aUJRD4J2o
WYAC5Y96GTmcuOc4c1hN7IJIFtrBI8N8vR5ZqzkHZNxq13MIZPM8WiORRooUtRGz
qsvXzEZrYpu1av3vvvH0VMLbsAyyjeMTl27gHlAvsAJSJeZpC+3Ay3FqsT5CoDee
Xxlpl78S3K/I0JpyT6+mWSQ/d4UGxRMFjAaZIDpJzkreSXOJbtVC6SVEe1+rQyM7
QRnyNQvVcUkPsf+206lpSRdItBSgiISdWCaMilJvkuAvu4V5fxsW2nBCPUtjvbmV
iI+0Av5vwty0GRceNECsMCYkygScoPWKVapCdYbE7Jh87FsRu0N27ASljQemBjgr
6o1sJg1sbP7PVoOw00BB58IALOj+EuMokWjhZMN+Fzb4uROmmBQoJQoFMFWWfDK5
s+zyT0OnQTY/UuyMmILvWlnuzcI2k0AbSYtUhby3FUFNARUbCL9O7sCpjvEAC2uw
`protect END_PROTECTED
