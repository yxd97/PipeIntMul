`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
w9kKrdecQ8ziMSTlod9pRX4Pnm5j0n9IuwW7EOzxllAc3o+5n9SoTr10ebd1XLJ+
FuK5bhAVzpgWlqOURwfDHQtE8UCvl5dNzzqCnhvbkGUZFvi47luGviq2I0EfYL4h
U/J5Z9ge3jNY0+G5//y9WGKVmN5ZgdKoLqYPbrROY85Ew2/R0UvlkjN4X+rDi3C0
/dnj2XEZLYHPrfLbks/NBjrT9721vXNN3zORA/mTHGPmRiedoLm0eTp9Rq92cc5D
2PxiXrNA4Uo/meL2lVZfkv1czfIPFThQJ2kEW+1j2euoI9pOSq2zhahJyLFCE4mx
RBXafi1ii3LpiOfuq40pv1Z6ZXlQWGDBXYmapd4kJa7UvAj9rwIUQ5DtjAp7m+n0
ryzCtlYGNS+49FtmckLes07AZ+W/tGzwRzAcZFF/ZGuE++ZplAZOa5pyAo05M0t7
qeVA20HixVeRzxVGVZ3I5BdtaTvZd4C7Yem0zs33OzypNISBEoGDNbTa50z13EdD
F4L/pjWuk+gMldIxSu6ZkNM7/snzKVyVum4NVRqtEBa+7l/DiInTVS8/ZFUy088N
Mnx+QKA1pHGjL92dXexKURhluKMoIpPe52wGbFYGqkwtTxMhn3sv0jsjT+3LMo2I
EBLsxe5PfVm8SGZeik6G4RWmGvd3gQWByD4uCkc+5AL7Pt33kv+/g67W2kl28Csu
rAjFsfPBcbMbKiQGx4msaw==
`protect END_PROTECTED
