`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7haOPSmeV6S2IecknqMrNbqQNq+AR20Z9q8fOHnMiHvtl3Z0DCrgGUqpeOS5SSC6
OwvwQuSsv36e2ykoxWSaEae6QSCjj2b2BcDKC//BfAuDgqwHRM1HLceqjqKok6Ct
zf7Yc6rogYfQhVWQV6EtsYFrn+NMcVX8RmYpYT4NTn1PqdPF29oFPabBLr5oKaX3
1pU6hJ0aJNX3uFjt55NiOKsSV4cK0zrluQsiY1l9SdlnCkGQyVnBSJ7G1vxGY/6n
1XPA5ZmMTDPKh0OAYE0E3zvIbg/n+PYlX+6kYR4mXYVZGVgO+AV41HofV5hQUL2j
nA9XS4L6SEeLfxxy23imyBw+ItVtGfFQfROBYz87qeihnNqjFhdUzdn+Yl4CNE/v
n6MBNgzPbynfXTqlajAGXoYHkJ//l3quntqdcqcW02nc9ieQAVBdImQ1ge36R2fD
`protect END_PROTECTED
