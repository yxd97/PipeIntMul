`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5TP7t9LRahSEh3OXoOTtDEZlFnATVAqR8vNi8SYiT9ZCk8wx4My2OZY11XnLBvg
fJq7PvQGK3QYbpApcwivCNaIr899U/AQd38TMvWa0DvvXUE4DI474VE4yeBjt1D4
Q95v/kCpasOUwF7soBdwBEPepINby0ebQN+AY4hYOhWXlP57e6QuOavRyHefGNI0
L/amWOn/ds0JgVfaI/bw/6YmuRmA1l4RGpsufcPaKynaSp2EmvvH1arvZLjbQ4eW
S7/3r3TVCggnPhTTitXC25ceZ1NtYgvsnGrDk/CwBkx0RP2IbHTWELkhgJF6kINO
GKKbc4x//gn/R1gf8pEr0cLFacjjO5eTthPkX4KkcrBUZj0xkpw7+3qk/0CRQEb0
`protect END_PROTECTED
