`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2DyGRItsxnC6sdsyz+fpYzCr5cl0xmQvfIu6tj9zBLrWioYs/7d9BmeKL4Tx1JqT
gpE2hZVwR3g4Rms38LGIS+0BMTrrF1VYvQ5TIPP5YBvFVoBe0GmQR6Vkb0v+4Iy9
JSkAnDC2jTr8rN9o7QWcGfpgDhZp/y/1swAMcvCBiF1x9QeWqLRoQdDFUalKytVS
DzbyAZqrb5spT/6t5CA8H47q55K7tYbl/MEKZxUQybXSiMfesQ1xnzn130KbZMYJ
MdDaq7mP1KOSTpL+94yQ8D1yN9VLzT6hIs9G3nO/7evGtyPIGWLf2UPT+zNkiWzc
+tymcBZ6UG8MATMKGiFBtP3QRitBBTEx505Pxleq2Y1LXtqMm1w5xRg0E/TJYVD5
CHuIu768rW8qfTOgGGsaVDuzgAEemu/RaTugRyT4pPymm6x0UfCHMn1J9fBg/TV/
1cWolkxAvqHuU1qnLR3BOKejq+p+PoPNgkakrEYPiQBxURgjqY1jhL6wr7niE4ZN
AK+hhMLeHe3b71FQW1y3tjWLv6HTasemionBgcxpQe1rghDyi2nzgfsqLLqfCg76
vkZZ02ehVqUn5OknQz9JgiknDXi9JmqY4DTciGesF97RGQ4IpUYRIw6bAcwVKvj+
DxcLs5GECOKUrxjdzEpgnPB4LDxRtJwCXbS1vGzLu4w9Zutc1dFqX6+VONf2/Y8k
I8sxcnT5RHMCyPWz6jeEJUq13bDJ03X7Y1ZdVk/oUAeBZCwKLDPTSilfiHp9GsAq
UYDhy889IOGnPIV1DX9X0plzOYfQ+omWvk2wcRmQbjdSKSJL8bfJOWDGbj4sXKDO
z4UaF580eF9be09gCyUahffIWmO4YBbVcAJkAUekQ1xCXfIB80XN/5syRsiRuIyh
WPWsFmIT2T1hIpxI0Y0qC8PkHjkUOdsIJmLEThrkaVuCyAmovtqfpB+16t6sIfgj
lMT8j+8gAqXzvdTLf8iP05tsBjHYU62zVs9vc/3376Rh0NUp6pVhJ0b5XW5955Xk
9JXLULzfrJxn1r3XjFeVzvdNp+Mf/b2G3Cfo5Qe3qnhbQOROD2IJzbGEC35YpDaU
1JN4nNZX2MD61BNcLXIOOFGuWqJw1NSgAz8Fk3qt2HGCgbr7stkrDNwBLpHD29sj
Y9KkKZDPOoD9X/aprVCMW6IWCDHY/Ohyap0T4uDuMjle/7Wu2PzsSy00GdX+rupd
XYJWTn16k6udOksJ7GePxOQKysuzmeeobpsKiU/q5NMBw05y1+dF9rq0CABQnvp/
LHjmY9Re8nLpolUfdlagrHlSNK1DD2ApbGQie87RkZUiG0BUFMKWnDXRXrrLE73/
bSgP698to4W3Ncli8qvJApPwBr75Hbuo7oCpB379T9mLmvhck3JjGjNx6nfc3bGH
ubTkXtpnGlitZrqHEQbHppsX8FNQYEnb20WRATUmBApaamUqo4YIu86tvDJDCsNt
yAyf2SXtEhfNZbRQkcsU5iU8e7DnE6MRtUEMi8VqLfW/fjOlcmgFT19ZGJuv4xXA
Wavn40DQv+trbXTaDjZieegY3uutR4pnv+giKuUyL53w6HYyPAR4h4+fsUDJo2oz
bU9DBwYBY9XdEfgoLcV0ln2gBVvioqQs2zGGIZ42EJIA1ga2pnYT7hVyoWLQ8YvS
DNKZcRBSPuIymcadvzxJ5J2lcpnx4HvyEp1EP+xZEuhIOjqWnTKwj7Vh+42pVt2w
gbR3HkQotcnhikc7rkciAnebDk6KIrAkVay5zD/bWCsi7Kq+MT9s29AU+RGmeXJ2
kAAJ5KbbNZylnUg8pG+Iuy7m+cMWxBijpCh71c6jV940LTcXtEvDW7szC+RktLrj
FalRzEglc7QrxOVcGA8RjAj6iQDou7IS8RLqk+hjslu5AaoxyiIesamaSzzNsQBJ
zx3Q9NW1fbnAZhYxSPf2DveFzVuz57f9iaib4zcqPhxypxlBPbdpKLQYT8RH1etD
S8EGafURLUGlOPo5C0mBhwRVQQlNg8IrEACyW8mrk6rSJCpmP8bnw05OxtHLeAvF
MjVI2c23mmos6kcjoYjAxaY+rbyXoxfhqKmn9/SPLb8yw0LfFKEZ7D1VFlhvaScY
JlvTs2RuuAQ5dkJ+Vd1xze7k8o6toD8+Z35c+eTpJYhCb9US1xJ5TXxcyf8B6YUv
a2R3xcnr4tUm8Y1FskgXE09iWBUthl/H53cGaDY7ZuPQ8aibknoRZonDATsi54no
DlAKuAa1Zk+OQQ+dKLqBSTeSaPx2GcEP3j4L2NEanbOO7MO0IAUGYXah3VLTewPg
edZFXzeeiLE3U1aVyggu9YM9o5MPNBza/iUV5UJLmzTcVaeV4dCRdtTotvt4RJSi
zU3BKdVe0ntbdcxRaDZjmCHEq+Hj77F62/f77U5wQ064Klw1Xw5zwGcC4AJ7LP4K
zAuGEEzXcOjRa+s5EuBX60UtC34ukLtaeB1echNoqCm3DelRXBgyosYTJRTUkqXi
4hY7INmOEsOcIdb2M3ZnE4Yg9TJb/FpGLnWtylrgR8hPRwcPSiww83eaHuwE4gbW
75qqjr7ZzqiRZHOjplbkIdjglKCa7qEgtirln9HIu9Iis40/VNTTbe/mL0EYEVzY
r+x/yl5r1QrMjAHr0KGnAN2Fq0uvnA8wGSFs1ig6yBOsrVdGkwgTS8hbW5uZndTS
W4gecip87QEHii4w5hT1owuo1ZmvMXP6Ry1ihZDM2v1bVQsR7HzvJHOaQRxCOaet
7+0FvEGFJ+quMNua7GXxMWX2OFndeklO1yvTbWINfv5EwZP2VZ+9nSPpFKGfP8Kb
Z49MITyQyxJmP89OtigOB1bwt9SkuNnIr42KGuiUoDdF3n64E4At6l9hJy3A9Cpl
ULGOWDWYc3DtY5DD2ejU1mwEkxrqE54CP/jKC1iDu5p20PI7zZe07nK0xycDO3Wp
JA6iaxxa0dSkfLnqZT4psT/V3VjrDyYY8CN4aDArPJG+lq5peJ4BDnJDVnaALNgl
zA/vnQ0ueRko+Km4p6yxRDptl2TimSFrgTyJTr4mQa7n11vw28LcgDDQbN7Co5RU
aW3BnUGWFX7uYF8K5RO4NfnY7KrvEgnHjbRlhcOa9Zdf+U7vfy4Lk+egxnp1UUzD
RJI9Mdw4FiUtlBTfBZBd2y4j+7qTkW6plFeYpKjQtYPNadaIZhAaTn/KX3ad9tHP
RmExZEcmHlI45AKmcTCmwufVCc6/TMoM8x1bX7zrKGGhWihhjeQRROyyZ2kVkjeO
Rrt176LCAUklcQJjuo3qiNySi6wz186c7fuvOkuDFQqeBAJS38zPKgCMVhRL/Whb
dAv93PYgAdOM9WQ2S2LpgEX9KWpAKTPuCyuQTSBpgECPIjr3s+RpdFCipDxYj9Cy
76eAEF55zt6STzrtmNha0O9Lb4iGGT6T2d1ygGJvAwEHG5ZnDWneIjn6p9ZC9eOc
ZWK5XkMQxoSZFF+W6EDE1t86DkLScyFFTynYnFIVk+VSmE86xEZfH5MSkc0pas8I
ZOEX+zK1fMYepYGPYzdmzwvrRjyAMlsoWe7THZ+7kje8x4tCusOLHbVrCHrcYabh
tjhwHZjTnTsDxOYgETRbhoo2tofQSpclKs62GNtoZInEmTCLfugRCMyyG6QZxZo8
ciLAza6KBU6FCXT2GPpYWCscUV0AQm2als1KE3tH3LEeloo+NOx0cOzwxYli3Vx0
yXUqFq6SqccXv4apK+mUOk0gluvKlwt2+ArNBTHXoN4=
`protect END_PROTECTED
