`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IHwBLSkXh2K1JKPkJkaLKgDVg30U8taq9YNBULuClFsRgcnW2x6FkU1pdkVlVsqQ
TLKzJGpGiXzKczJy/BPi7lW+cRpYeZXYZME021TLGzbdWMCUf+Uex56biXgJauXj
M/5mHwjZxbPbM8H54veh+R3Nn5seVzrlf2euJqpPeup4UQaf0/1CBONnNKh7dTEs
yPBXUdKdRIX3HxBgfR9HrY24ag370FJeAcqpIFK8vCMy2DwJUHcf6oPaSW7fySmk
K29fFktnYAWVMMOKkdKUDQaZ6PLImtFO3FlnFaLpw/PrghiaUl/61CBSRU+rlKQ7
a0e94ynOtDffK0vDLkUx4M6Uv+rXLVCDmx15VvfTlmGZpKcynSHc4mUH+BUVwA53
o/xByYb5Tkj77YdJiLFEVOQJXrcj/lMCr5ukQ9nRQIQ=
`protect END_PROTECTED
