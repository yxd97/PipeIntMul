`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bOXIGlWcWG48XxSulLwR+CW7yxH/nuFSJ6daQYzvcpTvz8wkljuO0Fk+D4OD1/wt
LqEFpyU841U58YAqduB4+iwPGZt9VgXAss/ave8L14thRDWAHMYieSvwURCrk3A6
9FyWyl1jF5HqK7GEqup4esKF8zJP9T3PWF5HrpPPIiyDDR9cwS1iZdpmqXD8DVBh
nETHOXuUtzyK6Z6Gpil0UOczaKJMewz71VKism7pcRib6E1gewdXwvfvJ/pZrYl6
5pT6/FzExk6l15fD08yuSZJnPab9vCy3sbsdWZdBbWbuLE0QjldF+LfmY3thwekB
CIZpSlQlxQViLFFLV5ZlWu9dZj4liKjnmnaWqFXQrQD0zGR8t0x9w5jA7lASfHZa
AMpQ8sMfpeRIwThYavbPvBR1vA3ioP3SagQ2v56xkMl2r7elJLR2OUqD5pChNIn2
RVGCF1s3ZlqrZc4+IJLUpyF4OILN7hs1/awKrjFVIkDw7mFcZ5LhKm7uVrXzAC9X
4s9dp9azwFDRXzxoTRK2WFwqrBEKM5wTyW402kgIvPmexnnktP5ERCFB4XM8URdM
3HX0SaDQiRJk6TimCsyv8sWJhMKWjkp9oJeCqykrdP5Xt0XoWFGX5XfYQlV2iyEc
85G1eVA16HWXqMNKJSCpIw==
`protect END_PROTECTED
