`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GAGd1gfFSEjQXDF39NNI8KU67Fvq592gojSnWPTz1L29gU+tXCysRcrblWGAzKw3
8HIc5bXCL+s5ybb5c7l4gm6Wu6VP+14xsudF9m1LFhFMExDlu5fXHje3LPVdOGoX
NT0Li1R9G+GQVQE58uaW68yvCfv526s1yDWA7Rdq6GPS0OJef+e2E/6tqlYoXdnK
QzDICs98TxlYyVrcu2keI9FmdxARGbtkdiTBC1CGTafkV5zDmPf1BZoywjv4uZJJ
f5y9dL4MvclafH9Lj8CqAqmsn83oD42gRI4xET9TW9F88iu5qi9ID2JI1xEPsGRg
J4fzdGuoKeN/jOwpWDrpo9xwIZev0jtgPCAIfJv4AiwSTCmnT3/5dOUznvNXLju9
`protect END_PROTECTED
