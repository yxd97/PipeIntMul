`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5EejuvyC+xGGOZBbT3QBUczGrUrbgMV0ncZYzIZrN5QG5+gdHDni/4O3ttK8vR/y
5q16qbt+Q/X+0S+wGcTaKhDFZGLOLKsN1KYjerpqI+j3lQnz7dkHHcIWXT9m01QH
xGvJbMpfBGW9nMXs+zjaI5TYJRK3NW7/UY4bcule8s6698/dd/GMZrFZJUiqW9r2
Oi+v9wEJoCcmMisd7NMWXeUavd30uB3yupYivZ9gO4fhcO/g6Diziwuwh91bx71z
4ifVrf8f6BaziKGQz1jS96hRtxJO5z4IMSQhuBdHkbhdxQo2OzM8Ll1MxnVtCG8b
AQ8COEZPc0qm9qlEq733Yg==
`protect END_PROTECTED
