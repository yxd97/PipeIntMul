`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dGF6xp/eXyomQ/FWfwJZ/UheSWV6K4SUxmCozLSA/hiQGBzG5cOMIwPXAa6PM3/D
1EwgxNFafj4nNOLG4f5QBWOh1zHY/1MPHW7GIvE31WKFNBdFoCnH+RUJ/yWhokEx
VdXJRfwarFj2JpxayI7Lt5uTnXU24GDG0yjLrwS2usRNmpPhocilIszC++kz0opn
nCmwk1kOEFH4r74sGVf6qlelD9L2d8FzUT7chPHHVDwk2JpDwauZW94EcVRhK9Zu
1z8VgeE7O7Uk+mN8KQL6Mj7qvRlGRaaiOkH3RoAQZKe+NKWU5B3XW0jKCjdw3W/Y
uWGYTsEHzzaRObMOWnsS1a6hSS70LOCfe3m3ujaLxaQ8ESBKERFYgcQviQ42c+RT
RWaGn7GKLmwIUM9zt3tNCw==
`protect END_PROTECTED
