`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JqTS/eLHhEyQ5UwAy8Y7yGZnmpobEhgdqwRs46Omskd3Oe9FUy9ACnlyfen1hbmP
iGxnsF/YQ7CZn+WQuCXtDhhCv9gnQAnH/YzKGQS4GC4Ddgdartc7/eAkL/E6K0kG
TtoqzoBc1Tr9/0AeHrxWI4kDBlQtm8gXw0S+UbdSMkjmup4cP2Rw5YQaUQ7gRWB5
bZuodpm+WDycn+vYm2SbV3AvCTBfdbdSJPLozV4KexidcvtYRnR63xjzQZyWtEPb
HZdxN5XplybkbAoZU/RVcqlglyduVKsow0kjfApqc9xK3rwI5A/UtVx9YZsZjbcF
bf7wJenAQE8674Dq6Vi6sA==
`protect END_PROTECTED
