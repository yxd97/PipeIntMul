`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
apv/VgFst2H8XcjZI6/Mr8m9ot51xn2nt/wtg44uEmCflNWO7d98bIrX+xKF1bSn
vf9UEM0IDhex+hR2LozHMhPMiVK+HCU88yd7k4BcOngcM9CZC2O7yQirdWcIzT/P
O02HtUYCuS1RJOgG8VxVYGmBfpcIRmDRlk1wJqtuEgroHtB3EJ0VcLMhKRBuzzH5
sayxMnuBIZzTZUwmiN1llswYPDKfe2sla5MwDOnb5gSQcvVAdbicRc+CMulMEmdF
f0tw0cT/sypgou/pybz5/BHVIg/y/pxn6xjm28JkKAsu1YTbZHxCB8GyeFjHFLMz
VYfRLub6zUsF3a6x7IyCdY8ASYx9lP1vznlgPaF6NjCa3ezMiv5GR4pL4s6Fsrpt
OnoSuvhwVssm5YxnCFt8HMlAZZwWR9+6I/ublLCCqxqwEwYQPYDNPQMCfYAURdyG
mrgtjWxk0kr9BKjmeNscZsoEshKJDNvYe1Z0z8pRtqccly943443BWNt/4Bg20de
`protect END_PROTECTED
