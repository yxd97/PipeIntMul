`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DQm3nmLY5s9BC6bQZcPoDw1l4zoSqujQlPjOasQYQljUCboH43XcAeI+Y9g38H9X
moTuLD47UkWx1YKbwb5AIfx9Zwdwmhvu9W+5bHOKg4ysRBDpwYrnfkwijmMqMtCe
KiSewRMsLPDjBP6OozVThsnK+hcv8X2lUrgKQlQq1/KazV54zUd52vuQ+duuU7ll
J6NCbBbMso8qyGp205wQDZ7NTMPGuaWJ3+fkz9zXY0+cntXJhs+/KZ0sYmsclhm9
pyDvEeAE8uYHC/Nel7XgzvWMcg6w2SAeYzYMg3nWLQ7Yj9vqFLkHd1uIqnwS4wdU
VMfKAzigEu9gw0BEcgoRyeBJtce72uEDEj8MJ2i1QY09BIJh/sCfup0Dyb7ZZ5By
DmhJqWE+bVTpl8uH1jeAb4aD8hqvtIL8E+a/5igz6XN7IgI2y2Uv+lWaqyI8LggW
rxmYgP+yZouzhek0JyxcHD+oA8lpGi6h9askXUKU2igOqMHOlLfsSTbfDrNEdyhp
4ZoH7BOWOrOGXPq8vSr3alpBOH8sYLbhF2Bei0V1B3zTxBHLsPEqGqaAQgyWpB7T
bO8dRviRW28QrSkih1s2kg==
`protect END_PROTECTED
