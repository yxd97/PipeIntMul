`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oPKXfzb5bLi+WQHeqyn6bvomS7xVsQnKw/52uR9FG6U6xdnO23VtYjh5KQgKDsox
J2l5RXLEH5Yfml8VbntUqCjbq5jtZxzWFD7eZGtjjxGDBoPrmKOaYD+kCGz3qx26
ouHMbfmHqC86E09ankk7G4Mi8/S/xg2a0iT5SX1I+skDduyT1aQB0y26Pja4mt4n
7QAokxbz2CW7qmnAc69y54r7JQmot65EoL/7moxzNhaUkhdDl0sSrFX3IfubJCoo
ZSCgGJ8az+OYef7K0Ca5PW40SYCsEIQeD6fTrOGfsuYh8BiQVnndlr3+VN3D9i29
tsx3Jx/RH4q9yqwvgWhdrQtKxJrKFsPgMzWhETAkwTSylpUAYOcE7LcalN3puTCG
kAi7su57zRyZkNtWokCfTFz14EdvXeDrPNOD4y3bWHJpNYnOUU0DxUnb1wLEcKfH
/+5xJ8t6dcywCIeXzSAUTtpmpRij25/jv7bRYKjbxs1sXl3DMNsIcTH1Ry7p8Smq
r2EQqSXVXq6M/VK6N9yGQxFuMcSbO2kGBH8AZ72wdsdzx3V+GHcU6VIXkGmJjEat
mNNrV9Ly3rtyoqxPBk4oDGU/s/qAXYrT7jFXHuf4suvsOaQjRYGU7IHAp2WL+Jcb
oTKJxeUFF2/D1BpsyPZJ+bGOvjo1GrNai2J1vu0O+M26zel8GTwBLrdvJGwqU6ba
E9zQQFRzQlO5I3m34uXvnjCUWnFGeuUmRzy4+SfesoX9Ts7nWgxyyyNXFTThhFPA
6wkvCsbedauieoUtDr//zXs/EE4Uehrjw4pM5sunYepWq4+sg457HWOkvsMt+L0A
kgT77DCLqTQKoJ/wz2U5rYPKFXQ0bGH/EgqTZgjULmw=
`protect END_PROTECTED
