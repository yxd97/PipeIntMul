`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
S7opNfcZiamjaDwp1niy35mCToSHGvmO8QnQ05UUCrJ7WsmM4xfnaYPqOi8Llqoc
ycVALy6/ifJOyehbQXxdOsUqM7L1A+jw//WQxW595UgwIhKd6LP4kqCA/eD2B8Ci
v3OugnPeInVcZvJ8j9ODZz4mTyE0u6mKT7Lil4dRkUoJx712y2+AyEAMfPJfqJvE
dZJ8yfEDpu25jjTPU21dlYihysSR0pwTCHwveLToS0hiDSkCLS9JG+ZKFNCYWJa4
TfsLBqI07NIpZwMxPcE41RvTS45KQEpgepf6Tz8B4yRO9ce2liXavCeSbHn2ZdSJ
PHNgFcHywEk92WlOpxSrIHWa4XmphfgbwIKBWyE0V+hABUI2PjSjWjq5yZHRLP5j
jBMkahr+Y59ZRl6pobAMtdD/V7RWhs0qhF9aVC6LAGepAV4I5Gv992gpO32pahBJ
dz0/2dRrpoQ3EXr3A1AQtHDAxYBzYDabwenY3s6iafU=
`protect END_PROTECTED
