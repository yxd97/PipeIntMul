`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9YU8PPFg+WMg29S75Cj5hwZ3PgIlsnpqruZ4qSffvEqC/P5smbz7GiL+tlp88Gt7
if8b82YFPbzsFg6XFHqKQH22xzMpUCwOaN3/KsFtSGJsosJF0lFd6q0BTm09m9Jv
iP86zgO6Srbi3v9PEJ4QaM6VHHdXZTQfF6JnFouX0+Evhp3Q7Gkm0O0qMcwVksyC
MRH9TVH+WEbg08ek+pAaoNTCT5eeUYuuN/UZAyJwcYSnkRF7st9CFpNknycmmbKi
xLszuGrpI0h06AnJiirIfP55vGJ8ZX1wPjkFncxeCrzqqyFxCw3QPIQqxBzKDkg0
Z8+rdnR8uvuT2hI1cB15kWs/3TFbrXfawHVij1L2W27tQjWf7eaerYjTWf8avNej
yGDCpqkLIByAQVb7eJ4DFt+F9dB0mbbDMky+F5TM2yMYhRT76YYqeItXjAzaSAIu
1qTsMSgbzywdrKeRCbuGJiSiRiK+vZ1fyJhXg5r0pn9PhLHkVq9jdNt+XEiWBieN
oVQz7pGM+5/vPvTMNbMCjKgijAPizIQaxwlKNAnfn/Ru+BSWDhySRjTgg9Hj+X+p
WGBobchvFvMywl46iDz8Z3hTifWq4CzUNENH3Kz5M2wWfy5fHyKur9VenkeVOa1b
VOTo1gzOIh/4qY8ZJ+rbzg==
`protect END_PROTECTED
