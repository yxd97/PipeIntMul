`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JUeuMXs2RLajjNdGgo/oLskz/BbunIqDcHnjQuWvEQpJEOB3RakB3OWT6YvgjY81
WkxxrUT+iYAb7tbu5ArulTMLht/kpcXa0CI3KvX6+m5o4ZPNf+q7CZa03+uHC9VT
4bIPqJyFbN0FstcpbtOY+dy/l/Xfrm21ooaq5CaIxzCgnZlKZDFFz3Qqa6M6vF0+
O+ug7k3lwlQCO++f3d5yABsHRYIo8/XSvuN5wAgHnjpqejVl9aAuvJHMJ3gU3SDW
wnwBV2jj8x5zHnWZMvBMhO0NACvQ+Dn/b9rH76bVDwnH0EMJMhcCLZWZsy9rFmpv
K1R5zEWjfCCT3gQlLPkl3JLbQlvP+OIH5o233Y6jLfsBwRlnA6ViEXjs8CPsdoCp
JkHeu3fZEbZLXrqy3aR39N8ZMB4mqrPBruDRnWebcQ+Tg3UYP4tsiN+9EIG2uvmE
TfhvEa1Aeks8Hm5ckP0p2awUdAoKYtofBWj+fj9cbEh/r1+AyhXqvbIZZUZYw0de
i+ljNXBtZ+pjnEBOV1LzHF9iD6b8P6OsmjNoNjvgA33KdLmNY+ZASQBYpK2bCVvf
DWZyKzi5rAYZxVm1d+VPJatmKHo5AoDZsl6gdmxDbAmgmMfZdi19bgJsbfV3Q5UG
XAxTNbZjV7uv0puHoZbfgG5xpZ1epSfBhWepJJfJGZnbDHyAIHjxOOk5vHMKru0U
zJEFSQ4w07m7dvROF9nJSPTGmakvI82H0Ag1mdLNbKA=
`protect END_PROTECTED
