`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5+jcvTcTKLAoT6t5FztTCpLXi+qlRhzPW3Ktb1uQBcD484m1VoRp2zg4kslPIT5N
5Olh0T0VHsforAXWaZNP4gFen4ph2nXoXZ5TFzIRFjcJ5It8W08Mp7tHYR1JfOZ4
FxKIkSKggaZ/fQevnnZligs5VIPJynSK2r3BkBkLRNISosTdnf+HDrcFDFEjEj72
DN1uJoBTY0Ls/fPwXYFyTlQtUo6r9uDoeC8sqnlfaWyexCN/A9zKAQ9dNi5IxUYv
OM+vswhoaLCbk4vhUCCLBO7I/oZS2C8u9+M8KryLg638PMgSxRyP9dqzXDpb5Kw3
EljiwXpJrGczK2YGGyf+we9e7sx7IdfnGBOM4WklW89Fay9HfZtxaMe6cZ2lirhP
yfQ0puccIeAirlF10N6Vxs2O3slMrT5iNJFQkWrDdMuGm4pX2xMPzKKYrHd7OolB
+YE8ZLK4tEwD9/YH+D2i+QwCPVDoY47bETb0QRJRRgldpWeUJuzODG1zPmAhyVv6
JtHvVdHU37EQmAFk7eSiV2mbAiWSdoaSUWdmctWflN7zyoCx3zUTyztaLAVUfn5P
LayOnFgD9ZV8DKy1qUI2Sku/4qtEif9oDDXciG39RIk=
`protect END_PROTECTED
