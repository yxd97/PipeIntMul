`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RmjJEGlBPK6SrxxdUdyxHyqyzO5OsWkIYHEAbRMhZ1TrXYlQoFTgbRo+XGrlDRi0
d9kONPSBXCU5/QjqDuOGJckw9JMzPbJToJou6+djnM15nNsRUpoRulwBeDkxHHHd
SzdWohfz2Op4kYqTnpujzv2o0WjG81pJ/oHmBee78c/ZsMt0HdZldemzb4xsRZ07
UX+8UNcBqVmUB/F4NHEzXYRvKWrOL3It9LDgNorkmHs9A1lz19qYJDpkgQh+5ZnT
HVvddkoRRHypvIXcFdNy3lBYMOneTb8nBRjwKD4QiSrZTIDcRNgTgac+M+m9xP3J
hDlr2sL9u8eLQwGovfkw1Z25/U+XapEQNE8JftgAXuLQxw59MsqO6GQ8DqRtYWXv
Uip4ThY1sdixW8TBiY6EDqYZADFgrt0oXSMGCf5RGCML46oXW3lyHfbs8YrESBQQ
erA9YBoEYFNOoH0ZWqDIeGyD3U1pq6yv8UEnZu0l0QqZMGte+WosuIaPfWDxEA7F
gEnG3Gv1kKu06c5iysb8d0XHcBqAusltQXbFKdE17TAgZ1cItCPQr0Oeos7GgS1i
z3yCgr8ude9f/mAgjFbNqIHsI94lOgeh228bgf4ox+CAQVbkDQSBwKnigLsWB/3e
jWi96RImFYM2XbslsfHWhA7aJJKTCMx0T3V1XjNVxQ8mev4GGEQb6Y8MQf2Q+nh8
/77ZxL7WU1md+XZOy9BR0oTKcHMdaTYWXYKrX41EZPVFerKwdVn7YmSBh44MBlvu
nK/dXppyNp7YwfKQPx/oE0BeWZ8TB+tDOG0lv4guppO1xQMEX185AvPCLyRPGEH2
hJcOcgGkdy+oPjpAVSw8Ea4580REpVLmm+LVOV19aZELDWBAd2AAlBX2Nawnph/f
wB/PVEYdcuyUAnYkKD5ZRZ1IrbUmyFNpTzyd3BauQ01n2za19cOvHF9kcTnP/xwd
GGl+9WcVLf7hmuNu60HS02pePDv/soNZ8DPXFoVdM+i2fCxeJui69Lnf9HRL92tN
YUe3BnOZ0PcegOIwNq3IDDkjkJg8oOkyae6DbsZCPzSN5VSnLaPGWoGsVY+q1/NS
IpL8qDfybzmJ/mBgc1LOas3k76lod72u2/sH+8PGIupLwhMLsjG7kAu2YG62rZKY
RakPwX+cb3OSXPBS0rJfF1KitCvRK/N7LFh4i3O/fg3iJLWXHCiFg2bbeKfmYM67
6JTLdslRQHoV+zF54gp6F2eXCDhvadpxtAWc4u117gI0K9fJpbp269v3haukKdY/
A8KQ+GsTQG+4nkln454Hn9OUIC+gT40DMTprtOLaSQVFAvQUxwTZyVle94B47Qvu
Vn2zON227CtcwMydOB2pifsjwWiuK6wR2Yszeb7bgETREa58rwRSGs2sHUMBiahs
JqcVfDbYFcPgc0HmASnl/rsw+B4dQGU7O04bqls6xOvHujZe4YSBoM9bdL7TyP7Z
h5EaMejfV5cAgH7r+H6x4FLSivaE4PyDudv9alL+F1C1dMFaxoHsKl7I/KD8Tyvl
jeaMdNUfArJ2cgvLNtm9/hERRPYw2H9jDs7RZGPdWVxcj5t43uzisFjLwyPSWHNT
Lr0i+dMsgXtlyyDQQRd2BpUK+gwQSZRnTYeOHF4+Pv1uN+CJuU6hwSMOvCvN08c6
9oPPUAzrRlfisEQznTiTunzE9+bPgEsTM8ZuTXfu30PIjc9n7uVjOJhu1t/bz2Sr
SSPtxqgfZx42XM2hF6SWJI/intCze1nt+TKcwnymoj9bU2DutEJgsYLcsTQOS8ej
76aCTIqjGvKqLSm5sOB5ebx8r4RlesCrX/ctOj8q3jCYaFJg9JLLToX3g+831n1x
yPYh/Mu69tg/QI6JZWj9aCBbG1qHChnavLDQ1FjqWQlIxTf7+LGo3YVnsjsvQlsK
OVth9YFXMeHXzBcgGcu7q9U4eL/pjpzH0wMWHrlb1zelz6J7jOnaC9QEXykxgARU
wLpWLBbqydRwTlHW79obg6HxHKqcpUmEEpu24ZbOw8lEcGGrwXI0bKfKN127u+Ag
7YiFnB8JujJDJblX+3qxpOhLTJS7tOwqKmzdwNFejHTANS0T5OEyZUXDD/l01hb7
7eMcuigALWzXAXSx6laPzF7i+xDhP5n/GJseJVvL+UpRwE+PLVFCFWhG6eHRgpdZ
3+F2nMmIOtn7cY3LvYXnX2wuocLuUZB684KCCrlmbmQ0V7rnxDj3i5xT00kNz5oP
Nbxnp+RaD681ce9lH3p/O4BQMVUqQPUrz6Cop6sdory/qYIRaO8say8CwEhKxkIs
NrikY90O2RjXqZ9ie/pYtPderN46Z1ctVlW4RCUo1wAoNthVukiz+/T6SbADL1Qi
YqwftWIOM1TRTtXku/6g+CQ0iWlntb716z1ae3MA65S3bmTiIZ4OLkU7ij6QIYcd
lWsDcmUnoYOtY9NKoeVaez5Hz10Z6n1fgvuyGa990fXH2WiJQbRJVigYhwliqxZ3
LV5t/SAuocRK81lZhR9qLwgD+6r+DVluRE+lLxEkr6pxc018X6i/Egjm8q1+eV+J
f//jHJjgyqk3EjYvwXI1WusMa3asHjuzLMoZfaV22OhGF/7C37F8v2/KeQRxDtmU
qKonPAJJUpLA89HtW1u8mDIWP1PxyEMnMBnHn1kivDEAIYVIJJ8Uj0TMpNxXmccH
WxU5EefIBwIvhjZIjHkv3iFZzSMORFVzgEakY1JgEFTXAWjyUGA3VC6bcg1SQxRw
ccs2KeGjmGnHdj3F/wf2IoMTz+m2vI76ifLcCKW2GiPjmRjKm3wOawq/osTfPmsE
43FhAt9TVmNIROokLgA//37iS+HpUrQw2yEDkroQbodlDnCraqlrZ4kyBvioQvYC
8lCbhZshUeIwLAaHGtv3eSnamPd7/3gESgr3cbEyIEPuXYmlr+HrC6cz64N3vz5t
yJdeYAKqHf5zmPeIwEqCzNpzFRer3u44AVm0gY9h+VwKbiu/vpEUQPMoXlhE0Y+h
f2AYoKIDoW3M2KgUVVIHZ4mOiWAx9BKVK0Q4zTMXF5MxdjdajGmSeJO4cCVGQAQZ
bY3T8TotnBHAFJkCbUGFHYMkVZ+AvAU2md4Caf4dRupte3hcm+FR9WIplixdG5Mv
nWPBSkiyQ/qxjHExK2rURdw8+j8JUnH5dPotpSAUaCCtem/q71Af7doNP0YYbBMJ
yqdASLMR6iM2tzvAC+3ui1JV53SZwLS787JRQoCSPomKVaV/LdyL778gKfTSP4Br
KBFo9powkhZ9FFpjMgO7eJZDjDaf0alLYBfG4wJcNI7WWjVz5RA0YfsODpchU3pf
b0Wlw1m3BkgzTERle/af6Jzt6sJUZqtjvJna1thWlv8tOZQ/r6B5FyxYOHAMcSaC
HVpCppmMQohQhcz1MBEDFHHplfaY6OMnl+wOq9gsRtCKL33SgHMoIT0WoAX82Cvx
IOl4zGXxYlyqhS7DLh+Jy5KsGnlUy4J8n04aODhabEIHZm/JZ4jjz7ZqPFMHWmK9
oSJggYgDSqsUTs6ACA35kqgf7uazaJYpkLMgnp9SjUC3lloAmoFGMG9SHL449LLb
EZdEVu4LdAQf8Hdrkr4p89Ez6hTM0JyFsImxRmeNlA5avqnYsvwxhvYxt0rZpLj5
cjJFjueIukudchYhNffmtd7AGZmE7rrabDeX6S68MiQhmICUXWGEJYfTh7ussR6e
yuWiAA1/ZVpu9x3r5WfnJZKhBxVz9Lr4T9cBbr4LMNzA+o7ldwb0HW/Ar0hXIzGr
uwXpQ0dtHilvpwChlc3yCvOty7KYyiVDTWrNroTOq/ItXBe2CAZ6HeMRQneIiNB4
93SV5e/iv2KtD3OAYX9lc0pXgrkhWtiQ3DReLIC2/QgJE7qeh1JAsZB7+rnSKL4t
Hgk+1ndUtTbrpZSQzgZ+38Eer2BYGf2OcLWGSRnd+EOsMKWgaImHMMh8b/KkMAlY
K7wkZcoq5Pw0nUIPdcZ4VeHYS5SDMrIvbZCP9hhwYAgAxHL6CotKRT3lqWIFoaQw
h/NCsTEwfzMK0hKHMmC1oLPJN0DMrizcJEzdP4YC8rLxiZ3J7f5jV3XV+H6gamOp
WQzMn16+KF4klnwFIMA4UbkGvSBYpOOpQX9lHNqErS7hSi+uelO48D+dyV04SyjU
bHbwZuYZR+IhWjYBptWLmt7nNImnkYS+oRQRUjyUX7/aA1g+0wixw/8U3A9/DJHA
EvI1tE8RfXL/3YaEq+zRMxXkjxsr6y1zMongloStDMrghFwBqILPeiTIU0THTuv5
Gs10U/wyuGCq0Mzzy5O6iJF2MuyfmmFwuuQr4f/fCUYJHTK/5andHn82qGaHLKyz
VHlBrcbv5LoozNXPNqpIe6oiuFrlnxU7GVNSvz1FwW4Bz957QLBsNglGEPzziy4g
Fq5gxzH55P+duM+cTP/o0F+M6+uvGQ17CylnT3PNmbeVjc5sPgQFAmipV6dg3oZw
xUD7k/D+/L0sPxnz0DahndLGH2b8UKDiEizlgIp2ITlEsLDZWT+ZIzpW8j5ktoC+
8/8x9MODIPkH4i7K8ZnIPkouoi1dI0zMmsctIepfgLPPfrze5rSXJ+33jWsmGoVa
Qn302WvYywqjT6bQSTVN4V/KOK6s4GZtfkSEE4MnUBbPqjDvh1VMbnrzt2nRgryj
R3cyhvW1HXe7VKbB84M3dE4KN9ODeKiq96AeqWzqLPLe0NGZ4uP08708y96wAh4o
L5B5HkJMy5F2zwtLPFcQKpr6kWeHbLV1iMG26s4wlmGk8HqszxJCGeIDmnHBe9Eq
8/HRorNk2XZ6WkNJMC7hO8JcQVNFIkZ7LXSU62L1ps2487buYMhXfditg5F4X2AU
eewPKOcAB8hims+x47a1PZpwC4fbEzEazaNCeNSjFuuwCEHt+FyEd3EMWvClJK21
idv6bxs2m8FmB6uggeWfTS0Bu4N4z+WTfE9kAFohjBWfozonbRahinOwEbe+ax64
dzkleEltRGn9Upji2tWB4aOVNx7ok8jsYhPn/Ms0dQPH4FjAjUCMHElPET66B/Uy
UfagJSudeV3iQQLP8ffRvoEkEO+oTH6TxszyOWDYdhfKgqEJi/8NGeZnLpI7VyVZ
cgA05BE7DQ/EIk0HwFvfy+Thr/AI+Az9UyW+kY9UTbFs1/G90JYHd5NR2ExEDuaG
2U7qmxxzHG88g2MMxQHG8uZ5Lu4ya3UjT6hHexhCSGVsUA3EjEnUm3V8TPOwN5cj
kcG0lacVOarWwEjgZHgbYzBEmWfUCAndm4BDlAZmmBAnEst07au9YqMZnYL6KOE9
WK0qLRiv+FnFi0WvBUPgKQr4jRkYJQ1OwzXDEKM8lorRIIP1yFx/QdrTlGfqKYdK
ir1whpWtsjJP3/amjrr2UQDz4xzvPzNc2eB1ZvQeqNwVnh17Ig6VRhvYCJHzukoq
g4qTeDvYUmjz8bf9zim6cF2Db3/N2YR+hY82tSzv52O+vfiAtNiQNmLJSGt4+6zW
MWqFMlNjPZ+vAS+YkB9aKiW9E8fiJZ9M1o8DJuunN7EDYfav24sdmstKIUSkuFdW
hW4mKZvM7wwWW9YUFX3krvAvy258ak4Ozb6BF7bGjplIoTZh0RHRsmBykklJOyI+
bhamSPYAL+6O/Z26Tc5zVZAabJvTDUaiokE/AraQ5Qnh+MUhsYeJclxduxD7bLUt
5RbxMgDF5lIKSPXCZNxMZqAugrUCUllnlxN5CGYGosyhAD/ldQ8+B+CGeGAD7H5A
5EIP1Lxfnru76QeTQmh24iTU35O4w9WH5kvCCTttZbljoGNzMDJekQwUdWYyG7II
ushq2ebJHYkv/NRpqkG8r1NcRNP94H74d8IBcGzoHai4INLkW5P8p8IH90wWzqYC
dK5K3JGzpk2Hmv1arJJqG/AgYvUmq/53W0w+zgjGUiP1aTJYe+SB+Do04cuR/Mi7
typ+oudODMntguhIccK++f3YZWdJLJtgHasAbUqub3r0PvxNvViZhpQi5aJgeoi0
4jadGw/BGDwTuGIMf5LKsINnF6Kzg1bwcqk+tj5IWGCO+CPzw9UzHq+II45kLU/0
VNnG37Z4BW2RX64N2o5HovcGp+sdfNyayJk8OQoB78Y9RDEc6nQvh66O61pEdR8L
SvJoiRtetoGDQs6YZ9CbYtXciIJy3+vDJ1Ud2pYddR7yhutOaJ8RNQ9K6I7gvWlV
gceO/AQo1X7tzdbNqMi6Ekfd5CT50lEadBWia2qNMvb+m7BBuaaoJ5jriNjjYiC2
kx11z4nH2y8T6x/uRWKrkk/QIX8//ICkcgiLLTr5xfkStpC/DXTH8WXgARsUqprm
jM8hhSRvcnXtJGekQq+7W0dPLzxwxstEy/BNo4+H2mV/erRAxJhzHCVMWHrKOWbF
3gO8QQ5HuaPnGHpCF00r+5Lw1h6G7v7avyMF5WXcWGKu8zWybAxxV6RfA1vSlLA5
dJsb+LXNtQW81OOyEHQNrzRJ+kGhe2q4C15ZoIl3+XHxOwftaHQd8iu9+9j6NAG8
GQ3wj9P6xih1lpfCdykb9kDfmASDFnnCg8MLMOTvl2u01LLo1KF3EyKBkyrReOi7
mVKrJzc5ZGpNxvBLIW4mKDCRocLLr2QQYXNUptK2dk4tM9x/Zpj5YLZYjfpF2/Bh
ymFwbqYlIm26mTw+qlqqGeSQYQyiyfoSYQcqt0C3Va7FV8xox83mhHSMxVngT3ME
12yQnIqSYvfgo3in0Zeles+WGqw1KXujkj4pdDSAlYiF30Vai8ulvJliWL+8rdk5
AeHbpxn9tVDw87zVgx/1uhJWW7PHLD6Pz9p/TWmJVSSOnl3WvVqmywwG4LAXNje0
amo1+CecOusAATwwzI4Ju4F/I6eAcjnPR/VNpn5tHybcFf+djYy2aXUAUQFeNelX
j3mF3q6YpKWpgDWDT1wRDiog/IfKkStZF54NfxwLU4KBh++Kjk0hoeWI+irwkRKy
X4BXsAaL1zsQ51Htb8If7QGfmlcgrBzKdgS8eFzQ9CLVZUO1o4plcALa6knFr62X
Uzn4at3L2WNJCguyBuSFT+gve3ytGW3aUmZaYj0nrgT3ILYyJCGx51WYnrKw5Qpc
DESCsh6P4FwcxfuD1BS/YwbbPY+NO1C+ZjOirRZCY5ZFuWRas1gRjZX6oVklngdA
wTT0ohdkcxdD03JKvtTIPJhlIii9z7Oi0yU/p1Lu9paVpM0zj3VJPEvpKjfG0pnU
qdK+LxMh097beFurTZ/gTHKb3mSrsEfNYt3nth4Gtiq6ooHLuveualjP/nMBtILd
5mNTGw66Safq6WOltZfxYgFCg/JopTFj41/7oj+t1Ovoe5muX9njcFXf1krn+Ifn
YSEFuLWPnIaz0JiaZb6hj0B96UVt5voDyIPSylaqyGphEvWxVCLbYLbWWkaszHm9
qWRzaVcWetMiNAkTO9UTf9dB0Wuo9Ha3B+ZaXYi1RY94SGnDL9bvb8lQ/bBIpEVy
RfhX1EqGD7ksouF8HP2vgtX6kSIHbGAWhoxB869vP5cvHSEf6zr+keUfJ2nuzHXs
gYgXuZr5ZihESD72T7ao0pz78PzHCmq1wxMxYqIHR80wO7/TpcGIZWpKpJRWbCv6
6+9Y8ZSwWP8tjJe0hdf+uxTMeRkI/gFoPir7bE9BB25ePzaiqyF31PeVeUs3EMCR
aH/zrsA5BA9shbygslD2tlm8tCHayOGJ5OAPsS+pW/lpxlc0tq4+/GcwvUvV9KXc
cgy7r+26vMUqqlL5LoBuN41XO7QpOZqct/REPtS/I1L8A61W4Swcb8ED0LnjwFma
nvaUibjZMrUF4GsZkAFdZenN7DcxcWR4nfMQjc9WhBM722/0Z33TcChD/8oXWktd
w7QResQeZy+6hybmWj725Oo9htPAC9L2895IrImxem6o7aiHaFSYhAIbmYNMnmyX
1OSr0Tq6Gibpv6smoA6FNblQ2zVCmCqC0tfDDYH81q+sKrUcowculSNlvFZQBxDP
qFrhrVnXWgdl6qQ2eHhX0SLYaNvqTffruMHEi9K+Op3G4kQk9aZoYzEx3fZv79ff
hDPLscxXB383RaowqgzkKnG3tplSbJEhkn2KzXUSGFjKKk250CSWwI58CMuBQG/0
xZQdDtr/7Z+x/X/2A5lCLQ3SDLku6m3yyPxbNOMkZHQVW2gjS3vfd6VQrvkzBC3c
COvvZi9GvkXgsbpcQJxbWxLY/NfGhfrNKz2jhD3rbVUZMhC2I0H7w3A0mtntPnTt
3y+lqK97PKKw5j8pJVOr96RV0mFfzQx02QPPXAQ2tkTzfh8IdPerV58scx8raG+8
uPlKSSyP1onMJrIAId3yQxX6+Slsew4Ig/22H5AYq+oBSl5JVDE1efKZ3tWKn8bm
mYStED/fSYCQjsGic+C6xG731w7DrFwA6RpE9S7kEfP+PHN4kNMpPYgXTZGox2NK
ZPoGzxOVIPkP3flWTL1eecIHPplobNNxiuTAnW4p0Ce3JFUOOUi+ah90la++KVcb
2dPJ2xqJByUtpChomKuil0DtfmznkkgFVg8wZCX6pJ+gMZAz6MZ5mnP5n49iDib8
tM8ioODL1g2G21Oop3RIrPQUg8KXgSv0lqsZ9yRLNwPnUIcLKEg+aoM09Z07A0tR
VS2TXrLdvo75spg7rQSQGrj+QRegX55r2msw7KsZD25mAWy0qAXxn0SqK0RfrViG
+5fmybJlJ9VY1DY3cJLwUmo8UIMzaLqivOuk9Tctib82nqkEraPoW7NISE7bRBUP
HJMQHW54wCVvrs4eknTVhznV+XbPpWwCWnBl98DOid2YcoYgnJd6T3ba6LvCB5fx
SOceWR/bTOFAngCiuFPESpwDkxEH5C2cOUNYGSjdV4BDHAAZcAeSOoaXDCO8NCXZ
EQHgh1ej8MQlyIJmGe9qCo+azWhQ+PCsnXf7ekTwl5r3hU2YqRX1mdizoi9s2y4a
nwY4dzGNnQ3u2/ZT6IfTtF8IF8yXCKp/LnVUWQf15eLFXVy01QZRuz4WIndP9zuE
tW6EZ4aOZBCHniEF1TPpYfrG3aGgeSfWrY7tuFtcUhaQVzZmacU9atT1KH6iI90B
RRVIEJky7xb0Fp7PASuwyNAvjv6tRhIfNMXx3xRrKhgJ5/SaT3QUHyUZfi2f7FMV
LNwQ4AIo18IVxOjfbpqZ2/mTJyAWyzJ8BE67COsyGz+LCgyiaO8/kfkIzUka57B+
4LhVxP2dllEYEsIEBAVGavRVNRRUxFNDIlw0s+LPzIm8uqdK16FjkKwqeqzOm4hl
2sCRryCg4QhkejXQm2NIS9iatzG3EPw2dWxjN59SqVsK85e+nFtT/3Od6puT4ySW
Bqx0mz8y8mCWWnefJmm1tv4J7i31NOa0ygFSttxKc04OzwKq7LlGTZUPPwSCm3H4
ozw4i/hoRoxUy3ssT2XHKemz8Xmrp/mokmbdlglatY7uH/HzVYRY9JYFEz2IEKzd
jW23DHXSFsalFQJ+sXGZ8EcZhirpC7vbIJzPfAFHa89uRdoSrOsT1Xllmbfg89/h
2B9Fazr/bpXSgKrIgM+nqK9DHiXbPvbMmE7EdePqT0PorM67oE1e+N4z+ADLnbbf
f6WFvsX75ZJcatBBnis/PaquFZo9NQL4ZDBHTybjH+wuirPWmnDFeaoUYolKgzbr
oVFTt7T2rRxBthADz0935OC0hGDSctv0cLkQU6l2MtA+7Cj4hRZTGZ5xUwmN8LuQ
5J26ZIwU3QLqW0CeB8DXkOTFPmvGP2mwRNTSDues8bh93OowmUMtyDk/bGEfffJ/
kEUCRoxnauMQjJYJoF5PJx/kNjb3VHFEaSApr5M7f1E0MhFLYjwNjyLCkB6j5Wku
scbvR0NEMe4gQ6L97XNPA992QfOw8UYnMnLyESwBjv2ffRW1zIyVXOB/fvssvOd9
ATicx38Z2OQ2a/ySKqr2Ro9TsMV7FHcR+IknvLmIJ/mjhUTmAwVBjq+NTn70v62G
yAYu2ufUd8/PJwXTgEIs2tMPMz3sR1UU24UOE9ghL5aFn1Evmdoev6MIW9ZLfbVb
eMyulChN7/O5IZbWspqRj3KtW++fZI0Rty8DQB9o5kPN9fseVTfW5DtTfr53+puX
Obb30MI2PV4pOaHLdZk6ELkWqhm77bTf5WAEFvLlS60VvpbAzlxKrrO/jhk36UGo
ij/4nzowKHHE7rAlR3936pCCJAygvSFWLT2A4h6/1dhyQEMTh7UOwTBCBBu0Xj9U
BkWeGPPmHWhSkrSpZnoX01EIHBImWBdx+XS1nmNDzK0KnSSvEuFEUup5fM/yjc7Z
HLQghUS5sASHbj3k7JmUnpIU2NvTl8olQ7twh6uOyz4Lf3aYvQGuKVA3oGLwhTK+
uRNSC14ZQwv5SaYHcpVtghL6TILSddJ2nvIOCy9iLUnmXCm9ogeTNLEvY3eNuNpu
5Oyo9LKj4GQ7tICWjUYO95PesTukPMDdfJWSN5kUEjMqSuNMTyr46r0xzzCbfMqs
liKw89gpg2vN90Ml5ePq4xDg08JHogvEcX1rVovhCXiEJTfvt0Y0MM4emgqTADEs
TrsqDrlC8sPlzOxe+LLNyC12nC0eQLD8ZA6OkN2hrLNmORXGct79vIjc13Jliy3J
RoNFDqoZnjgdFxONRoHHZ6Ap0BB8DPuZM2U8T37ZGH2wtW+R+fiMeklVGFo9MN2P
zsFfZJ2SAg/1fxj1DanzKOuTyv54sq5Nu4kbLGUR5HRI1p9KVXii57dib9uhtxf+
6aVA65P0JcBN5ussJ7pN29JmF4BmViCYSAAJFNboBPb/6mu1FRW833o2zXkNO+iE
Hvow+1jfU3+Rk7tauB7k/OcZ+DdaIL9PV8LArxhvRuB6t9rIG1Yf88+N+ei9qmDw
4lSbjbpNlbp5G+XKVkdHo6qVWhjeZGzwMCDtsx2D7sbDDM56f8I9DwGMzGayf4sC
PRhgJTPV19qVoauzo6cG+cOqOfgJjuOtspouX+IXL7wFqRWauQ9+jdh8ruya35a4
gT55ZZxVtj9w1jtAxdYhYC7MJ8Sma8mzE2zL6x7rABivfLFle1rP2QYjLdMmGmq4
FRopeFDv1Rel77d0sZb78Dfsbu4aSczLW7gem0Cbtqa03cHb6qw0CnFMdvrV3AUA
OZP8SsU1agQJXCSUbHbWTWi6xZdTRBdbPgCNUoodFPmHMny8j40PGSHcBTJIVqMw
4lLt4nlPk59/v1jjq6T4axp+rE0hyUvMXPkoZKX0ITYGaKqFQHrK9KfIVszKTKm2
nxQUOTNRpaoh6uMk7NTD6Mx1y33Tg5yDPXyVhWmS2wFlAQlheTlM57A0XllXlmCt
1MlqnaaJI3+m7BilXLDkudH1HC64vkOaG06nyGPOEi6p5FvjZegf+QX1/IEl5JaX
84uJW/mPWo8bF0XdagAOUevQI0okD/5DjJKv5pcWJ4QaxJkhyzpr7VVYnTYJyoEi
7B70ssX61b77uGTsWiexG54jyfwssBLkdDuq7cGcFGOj3Sh//2jDAfiWlOCCCuje
Rff5uZ0pUq/nTZ00S1GcrQko5Ap8JxZvaiCq1iGtc7OqHO4ToExD6OmFWe4UI06v
pffx8MWJzljFQYbluFP3kS9bIPyDYo8FvA/FTy0m8oyVLLa41qU4m6jqJlRFps77
Z/nGgjH9m7A3mN5fyd/ivoMqiVA/YdcUxfel43qayCj/TMjeJLikBmkKc6m8E3EW
hT90fyZ/1xLZqxfs/+xxbh3S1shvjxU38xmasTzM/EmsfE7DTCFKtWEwGc06xTgZ
5HaJBUmfozhmcv6btGZmWMFpxLZd4+j4VUPkjEILfY9BPMoTxdyOEVTkrZdpLda1
NmmwZSoXjajsXc24g54qt/Ink+lFNydPFEcZ0812tAbzo4zpwAGzfBEVRz7X8wB3
wrnrv4qHEAbQwDfRUlHH5jH5siO/bZZVMf+y3NV+WbfbLOXt+0sAVHDTKQuvB8Mx
Hf5RtEuOuPX4gajz82rVzzkSk27Nf40DPkLp1tiXzd29kBgE4IPMbNmH7FIivWOQ
Hoc7okcnZ1Kg0608iXNhVMcKYX2bL6EbI+xT/w7rfpRIspkq8atX+pAXDaS6pAMM
N4gDKOnQMl8tQcnr/Z5Gl7AjDqtfdsoLzHEUwx13HF48YWi4BvHIToBItQXuFn8m
HyCe60RLeUpebI9HpC1NHeJv79pFPC+fvEWBqZC//zA4i+LLW69w0cLL6GypnFRV
+FTtGMfYw2yyu6eF2+pe8enaDpJFXKnk44b1l9BAuqjTSV+te33fdnm+1F/vlP0y
CQq3v1fx9bwqQKS9LADgXwGAfTivIjwCszyjLqgv8ynUI9vtlg3ZfIOcuaVoo5Mf
RWdhQF+HTvknkHSFd5RfWlT2XQCb8ll1IfEqwZCY3n0Z+NhZ2INhGt5scrvqsvdm
Hw0avwK+bpiboPqxfIOoYFn05wsKZJefO+fxOU0c07VC1XDO2Lx3NTHRGjPW858z
vgjXvZeRdgTF/jDVoAaoaHi/r0ThxTFzjX0A5LkZ3WQGJ9AnTAfGmFBan1+v2G2K
R723V9cjsU3M+K9DXPZO/NoMGZJ0HKldfHbAxeKXcbY8l7Ftd+J0eqrgeEdAY8j0
x673mdkFAtTFe0Bm5iyvwSeauR/TutlG7StvLk7WEIpAf0HQ1PQCIobX0m7SsHup
nL+NcupCF36/n+ccZjoJI/gFhwYEZkhYlCCe3UKN6SqOGbIzvPk8IdKdyYQPQPC8
B0pA32vCWaVGSLok/THef7YeQThbn7l9sBWoq9l6/1wjLgyqwULf5LsS8LyN863R
V7DPz8JfEeiM2WPezPgp8v9V0IhXell80nUimsxJeQodSt8nW7u59zPSJ+CXG53t
ovmqbHfs0Wtvijmw1+wozy2kkAkzlv+xpPqyo54c+yCF+zsl8yfhJmWx1eSkUaBZ
/9ebnaEHVNsMEmpmEK/dtJvihlkCkmXrSHAghu8P2iCCPLBLdSfVgTpZDbOZwx7L
E1glJUuS91PFml1pB8BRi4GnLeUmVjfOCCg+0kqGp44r52gyqWPk0BTLO196hX0Z
sVupwepAdfK1RthiPHTU3kpSx6zIoM6GfTR29UjrUdlA+zvFEqBr7XEjn/JQveIp
GuSpZcjC9zxNlcqyL7YtFVSnJNbJftKqwAvXEOqGYrQDAibBIMxM1x0Xasin7aiI
mHQ0N+C6Y7ax1ApTHCJ7yri0kb4OvBnzwP7xbMRzIbSBtw876V7EDy96/RU2y01V
Z1vKXsKwDsYU+1QEE9JQLlDQF33JwSaSml/HNMbh1kE1jHWB9idinC5lxRUHK5In
/kANzOqPnSXHVf7o1aA1F7+I7uTxg9xkUWh8kbkusQSooFmbZyMLKwtjoptQDPE+
1ET5iyrNqfqMq4xAldzTNP+Gj1577yc+UkVb+WYIyhCpw3T519QCUJtPpeOittmN
wbPOXLh3Ug0UE5yycnz7Xy6UbSsnPwHoYaGM/uijfz49lOp+OtDLUDN/YPimY1Me
znjEApRULveHjHDSiizrAp5qY7ZF2XcDpvTUedBDZQbLWIJb7FnOmW7RtcAC+LmJ
bYnujxu+6WSc3ynNA3/6UiGK5D85j9DDLE7igjB1E6CsiOdxY5UQEw8PiILJM0Xl
D1ceyEod+34iRlU2KtRkHlnIDnewqJ2n44gluCiVrahGC8AD0Lr/W0wkkaNe90hr
deanFikb1Is1nEex1YT80tEKsuBOdY/RvrQfrQdV5o1R18ht/Ky0v0XwhvHlFXmR
Xa/tdUB2Vcigm0iSaI2mdG4/AbEzBqAyl9X2bC1L+J4LSAcSVWcjaBvclD0BnBxg
IUx04vuYWXSgFJLIGqnCM2VEiobyDI1sdHgUCpthrsYVmi/daovPvHuRcSNT7+f7
XNHv2su+HYOHzSMDuQnwVm3jp2fPuc8Jq1HzboKEbbuRtyVX1l3lpH6LjmhN9JR9
Lx+LSXHCGvmvz5CtqUsjREkJ24Zev10eOx+/Plv5ME+vbVRQMvQBABWm96TdMv6W
fXRODcYSOlF1r+NDqNBg8LMKZ5awkHpnBfJ9qN9GQ9nj5yc5gCk57YtFDIv2sLhR
v/rolxEAr0r/1wXwYSEM/846s6glV2sQV4GQrrVcgwnuyAlUDHQA8qHjtBUY2Tol
0sRiVI+ekYEFlGRBDiQn4GoYGGWaKHIQbR+m3UMXs1HQt3wSeoaF4jWogvtEcsXr
YoFT1u7tYDvlis2oaXzZ0pGmAP8fclzcOmaYeUZlvlziJ1/lbofHjmOZ1VMfsJ9V
wy4OREyAA9fe2kQhXCtmAyWHwIkTpDCORQTAFr7lZVH1JfD6IsA25MfnXQAO+c/M
eJpgcv96MsGylsMuac8pbkwjf9Uv0+jQgkXS71HTiXc9ZUNS3B0AEhSiSQTtlXxO
KwgdcFHpnPF0n/ICMa2M07v5FOijUgjEP0wFc+cddolR5UX0Tv1joIjlmovuSryC
KaiFMWOyPuBLisDZy6MS1S7EPqraXhBEvnEng8Eje70DJq3o+oG9+3yqp8vHn9ZF
XGozstwTWe0DuzXO8mCBU4CFyJYt52y+DgLPMKz7Az2ul5i8vttJGxQ/PR0IG0un
I1WobIXxkqMyXR+iuo5+3AIDryiRtkYzGTr0QsB8hn/wgR5zpSoxMwW3dBheJBJg
lpHvcGbbai3lShtepsZ5JM0PhpZd03C3d49ie32SdzE8jbTKcsBxTsfVzRywN66Q
/JSqwTb9spfLA5vnL4H7E14X6GXKz1/LtwI6tYYRSrFNzwrmh926d5+f70fEuCU0
+ZfHTYyNO7jRsSTOT/b/n1IqTxD+B+KLRXQvVBBPswluEk7ml3QePysdkTHPOrmx
nuvvngh6SMkZDgJsUr5r7VuS8GRQJbwd2+pWClsHAlYSmjTII+siaoB+9iUGVCc8
AtVWRoq2p4WOudP9q3f3YBOJvIHyus3+00NZzrtCJsCNzHHLdziPng7By57e4ety
9G1B+BIz75miU721yufclEZwlwD1V8MQaAW2aEP/bkpMJ2fiG6yU8TgEBGBxRTeN
mDer3SZxfIdTG+x3keRSmoZstGtpX4q6/Rv+bOrF3r5ARmF4pA3dAJwXZt2X9igi
tkmkMR7haifZ6OWoc9W5QSyGlwCBigmFpJnxH9JvWHZQe4S3H8xmIhL/L+tAB2VH
G6mBntSnRNHCoIeN0zoLQTsKsPgEN9PZQ+2XGkBhBzWXfkNssZs7UnjEWuXK1BGz
eHO1cqrk1QRXYDqWGMMsDSIY61Wu5LJoCtf8i/vKlLLrVcwDJrW6prPoqq99ubum
IQdtTMeQaMlcne3E1yNbmEmV8boD7pMtDvTEI56qw6OBIbeLhu9ZSYfvMAOxDHRJ
24HdV5I/Wdksgn7OQBKomrWrrwtYSfjAUqsjSUSIU3TrEg7K/Ua2SY25eYy0Dz6+
sEag1rJyBOe36phahSjlH/+cB4ptQ01FVrUOKLRGgxi/aPVCl5KkU+A3ewGvBXDS
ilWgBqkjciaPFT1bsMTWftHuqcfq5f1Jv6GV8tTOCFu5uohYxDcP76fQHqFT+ZrD
V2fhNEQuxiyeaTOujYrNxhlQBn00aQfgAnFt6GHoFN0mcMHfZdb3so/1Q6Nq43Nr
Qqg6vyX3Fz/Isxog2kN6MEFej2YV9BW9fQjwXwkia8/kCUiPgXGUcvDAdyrGqX4m
hPGg2g4MDUUkvKa1oGijAW6B2/TI6HgjCUubS0gxdioLqIUPbt7gHGVfigVCLvDC
n34ws5Pi9men0qAk+53jVZGBulMzI30YDy9svlOpBLg9ZoDMcMuCDAisNAHmsSe4
Q6cirveBx+Z/aB5yUPFCcAW7RvHQHMxbMakKt/DDTcQZypyp6PL2l7qnxPvXfCIq
UZGJRgRuIcq+6o8TbCH6T2l99pIVXK0M/pN7TgRPI3dJLdkuYxvDeJXFnx3ZL1tN
MYdiNmp+cx36Q1n3owe6UZKQdHqn1/YG87F7jK9GozKGPtf2vETLYzZ0I0oM9S9E
pKF/OpcPnFuajJ5n68pC6NffIY0DrrylYg8qPMOkabSztaSDAsHHEKJCcljiy2hz
MqvrkP/l8g+36Y/rTA39tBav3N/PBdNI2qiCSwd9BljoEGk9qp8Ay30tcT0gmhyo
x/KmUrGRpKTNc/lCVgIn/ZFKQfNT2UEWKMRVDz8/+K0Gy14gHDm/EY26YW6a43UV
8/1obfkhp0g4kftp1jiJMARZh9A1uxVnsm3tePb+JD/beHFo7D2IBs6Lsfp9LLjI
hV7/PZTaFR7RZT0yZU6MqOva9JFoFD/tK3nzHxUrps2TslKIgyLGXzt/5LGxtZiD
lm4Ikyx+x+cujcfdIN0C1UKCo243Lk0TVE/jsGj01gJNsw+SmMNwRDv+FXm/A/hV
njecBZ0tjylRPrrnWKwV/4I+t1s/pIIgzu0bcPPGp7GYx6E7+n8gZ+WDRbpqeZRN
s8clhDaUZd3F2UyGEMXLjCFVanP6HyT/25Kt3wzGMbTdb8nkapA1nPx3DD8O0XL3
+8DsRggHjak2p5q0vdnlSVXEGiSDNGFrQX2te6PcjfWHyAs4t5b4Pi1D9H644/uU
o4PBqLd8Yf4exvCPd2a31ky36GS6S/DPAaKHyacSpAKWHlatOFSc+QmZ5+9jlfUL
Ar+XIo0547woQAicwRJddxuXHAJVfr391ZLbnyiF316qpVyGYCr3cOKGxg7kH5MZ
lQUWUxjJ+VWSMbFs/UZ9YXAz37HXN9NwQZJEr0YaEfj0wOc4xGdc6HKzRBTwSf6Z
lxNOBtqWEZPVYUfAx71v3jxGz11dtKhduuf39bP1uhmY0LQ4Q7pQFZYfXOwr7moT
sk1zafuDpvps6ETJoIb11GS0KUELFTswnlZWNDkZ/xS51px80wRARHxJN85sGttn
TV/0jNn2eaUgFeMzMgcoFaceyMHC/iMzj9oKy+QSVtRzd/mqy61af5QRNh8/eG7V
C+1pFg8k8aPDxtJMQ7OD6ZCDT80AXvHilHOGFUvkE4uObJ5DB05PBkxU0kkwMPTt
E11kCqiNFTm3YKz9gKAtI2H4+Snm6/vhraEMwGsBNAgTyitrZ6YpLNKe7bJj3n4z
LsjoCDaxyPNynBocRhsMN0bGZziP/91Qvg2RZdFjOnCZaq1iL1hTI578Qa8TnG5H
VJv7i97QdL8aOGisX1taHoz9zczB41fegnycg5fWUJ/nP4sK9fjpMAG425wVUuzW
NbadxTi137VXo+vdQxWloXlc3cnq8bLezrbfIgorm3rQl5DAUDRDBVjJQ8mVFOmW
664Hpp6SIO3R8nfPnBZTZaHHelPfEb+Kn2psZSxOQAPWdQ6/XvK4qWNCUnadI4IP
vv3VNkZzzTIlFMi7Yx96hE6ZXr/ufHGF3dy1fgSCQ7xspimAhbTurES81VKdBBt1
iuJDU+H0v5c7gI05a4Q4/051wAQKoZSxp7T4X6b4XGCMIzc8TE2jRHUUPpeiJ4He
PYuRviYnPD8Jyeb3ZDaQCUL2uDWVk8bsaANE5FlLPktJ/7/NaKkE7L4z7NP/QIjT
FEHS8kacCeKgt0HMB4JpOaLXiS5FnnXLjgu9NpMBCk5d7lZNoubJ8q2Os7UBhV+/
Z9HCSDU+D4ovgb/2nZjgLjrteF1TzAd768k2Ai4kquj+WEZsOeWUiR06WY01wSdo
43m0L3gI9quyFqZwjJOXbQEa/T37eZ3/17jW30C/ATyrLYTEacP5QvFXrk5i70G3
sgAbfU45gAbeYW97c73BEfj7JnvuGrYEARnvWNVXHYS2Chgm5nZL7GcvN/vQMCm5
yBkb8O9xu0REu+fHqU52C2gGYA6CSCVcMwbGJ77/sblS6lrwX9gGQPbY7ZQ0PSPa
DKD257+CtQpnsKlyAR9hkJjEBWF4Z4AwRqKMEr1j7O1J/2AdTsOXfd+wDU3AtsK+
Jy2mqjmvIUfT1z9b/BcLqueIf/+1tfKCx0mvn7uFcg3VIcJzC98RmQFHHZAid2hw
Oay89KWzHFZjz+6a52++4Gk24xNIqsZykbTb6BFBMFSO56d9H7IGGwfpT/mKrAER
SxM0n2KFDVvWVlBVgpXKJfLzpMbMT9DDoDl0bJRVsxLOCMtWiHrvVH0yOPlEJdKz
VKScCY5Akio8tE4XZVplS562R90Oe4POKag26gIk58hMUP4YwGze/lDt1j6JCud4
mX8criwiZapoElELYFsITXTbNBInjgHn4/jfmtyflfbcdm9fadN3tBiva0brp1J1
9JFNUHokRCZQZstdTKoDAkutc0u6CTcRtmPni/t9Vh8DLhRq9sN8QXHZCFgy9p9T
0GHM4QhaTVERCLt0usNFz+/JY4bTKjvsUg4Af0xMItFGVa22OU6RFqf9fWZv9rzl
9Q0iyVv4L0coMbjfj8Wl6Y7VMX2+6RbX4k4b5WoM2zlYm33sDJ/rrmt2B6Kc72WW
zxCTEpCoTCsI49KcGLDdQ782Rwl3l7409lIEfZy412d84x3yVZewZI2O4YJCNtUy
YMXLLE4zFFpKL6QAGbimMuwnKq+bo+ooeKt7bzA6a7ORT0gONuFCOPn0N0ChQtjq
TzWA/v16KRnK9SmQ8PvZaruJFqZx069LZi/qSttNtdvJAaaxqrOgXzo7FZy9dpTL
R7g8wpd9n0n3wP8CxhAsz+f4mGcNWC5XpJJpcTZiw7e25W6E/gOU//Q10GgQEcco
34oyor4OkwuiPcmVI+fKqXc6Ap3G+P/L19J2ga7uBp0WuZJYF91fdgylpIPsWxEe
30BUGWp+GlP4o7A7fulf5krticCj4Siil1g3FOZpIOnvHi9tfgS6x140M4geFhS2
aRrbzXZGWRK+r5Z2/huzWUOVqtAQBsXG8xOAY+MlcJUY2phd7pbhZy5MND+JoE4m
vBMZCZv6tr2fN3plzmsrbQoH6f+rS2JeM7xP/xh6sdFkyCKCSi0rJjxTXD8vp04I
XJnLcuYfT/ITbuqQf1NVY8mli2qEMFHmQ4oTiJeaMh/i+fIr55ep6nS0avIJuqSP
BgxCAuAKgX51OZUZqMBSa+RTf2fFNCb2W3Xjwz3gb15SvNgtUOwwCFXepudsXQ2f
FWoNjIomYtJLPjusQdhrvaYze++LuD3Phrv2QImYs+6TEAJ6MCLlco6DXp/8mvKZ
A+gnqJN6FdYm4qTOMwBRHzVg7dhdA9pRf054RbXsCzfGYprijfbEWwCGcA5xqcvo
tFhOEr7OFwtzrvIAJfPw6ckHcJtSadw6RjYtzLtRG2CC+9cvmtXzNJjriop0GLOK
izcJ1IKWjPl2y/OatpLqWfXWxW//ChhKsE1/UTzsoLOsfYMbA8XsIT7DQfgWNe0+
DYiBU3DA+SimlZGttws/xFC2HrWmTxYKiUU/CgA42nl+E1JzldHZM7TlbXr1zCA2
Z2McEescqozJ5RusKhTE7UFtJNX3ap71Dl+xoxDYFfnrt/idc7CCXIBZIyrvFXon
cQPctE05TrX5urqErxAYU+r4QR58RXhPi02yJzfLNjWWhClR6/4vUfmV0H/Bzhav
qK8Ev9yINIBmmwjt1My5j+hkIqKuXAl9CJuTbXU0fR94ZOfiQN5Lcq1LrwVpietR
DbbccI3aZGFHR+TRP0jDK6Qjb43yDUR+xuTb1Tb6Tfed494pa+Id15bdSs6Uf9Ke
dldR6+nr70z8zlN10hEUCJhczJtEVNYFXtbg5Uym2hM+WNlCUdNhgTmrCZh9N835
BnW3Hnjj2ZW4ukfgpGMqeJNzX/ytSyEynOqWzfGZk4JcyloZJpNLZN+SWf8sBkRy
fTYyDEXcjACvVx1V9qThq6b/1IB144t2FmUFVOHMemru73KfRV0FKwWkXIcgj66I
ab77KP8VCUpOSZI7aDSj/jGFMieQ2LJm4euyW/PC1ajOIWllA8VbI0EHyM0S7PgC
bU01MCschRz5wjbI/VIanUEqCb7B4kt7peYRsjOxcVgmMtvFTpVY80IgM4iStFVe
3qT5l2q+I0J4UEp7DPXjMmq1sUQpQYoND3h0s2itSKtfAGNAzK8zRGP2CfjU+0gn
HAXC67s0uiA95Kdd2inOI3fhRDCm1H9DuvPtIriPE8kPhIwUacVzk+fFKpq0btt5
r53l+O/5khNvoV7gU26KVIJshhKTcIRaue5xbcXYWZhQC0qeUp+oTsP1YZv1tQ8b
bzRTAHfJ8wTh8VTzByMYWyJLeJePLgT5CkQgcex0/7T5NaEWqTMSTvHWkLRpEdTn
siZtJ4jIvtT7lX1/RTPOoiyJ1zfWDtxUYFgPbDrfh1NgBqTfy77URVbp0PuFrm6s
T4WRY972GOfsSZM6ZxuV42W4RJNErQ85MEtUbDzgYTdRoUu2w8N7YgUTR17zt+u4
GIYHvzkBaAd9m5Kl202Fy9rOBjgBRouL6mGAouDKemFLwK4XTDejuAZU5b4zyPVt
1/LHvqM5MrrIsg7ekhbgdY2GTqH0jSEFESAd9JqUX2UmeR5sMXi0XvzoOsd4hJ2h
nGwEeaABOKWDV+NdODgwUp2y6Sk/OUu49JFol6r1OQzaSYTCbvGZkjJNLNR3oeUc
5PcXL1yVXEh6FHyeGaUpC3aAeV2KWGAIyPKPoBdpzS6BHqSgbvvLufdMrhVpLIzo
90ov9y0anZFGyNRe0LVNqeEWElR84tsA8SWXABX3O9GlN8jkC8WOUPTmpV3laW0h
5baU7g/o/ANyUOGp1m8ElbCLgnH9yFi4GWEAVKNl7xzst9SOhjWtss3Fm+GPB2TH
5AR78tmFDe1/W91utlZT+x3HXXp9wtOBtCBEM6YaCdTi7mERHSTDIbjJ30YFv5Va
unGwoSTdsz/vHTp/cVbHHzCtw/UrshiMS3A5JxVTolwX4IPFmMK8hPsqDuCAZNUy
qWO9ufKPD0qvrS+I5yImpjJx5Mkk6XIgHQtsCecaFk6PA/QXZRbD5NSZ2Ny4NYuu
X8jOW43vquyYkkFqY/vcUdwvMMsf+Vjwza0p/CRVVOKbpRjeKl5pxJV+ZxD+6cvW
KqatFe6OwjPC67nC+P2q7Mg6SV7yQzkXcKFMOe1SL5gDiueMIs48utifnFhNV0jj
X5tsqEg6Yu1+kdRMlgRLmGKJ0QFa4aJRdNxkGF2RCb9dEOb84AnKVzTCEUfprIC+
kqBW04Y1OfZkkNEwdgfhqUCRfx2emkeNxvUaPDxeqieQ4HQtqA6mfK4YXa8NL8Qq
PkBI5eb9EVTpMNn8sdbKW1uB+6vhapY0LGhEkPzN+c2cD2iDU9qZEKedrXJFD3WW
xu25vpRonYGuL/E6ZA430Cm5tc7PvU5wrcgZLNUg/RsqCvfQ9PUUH+E8tgeBSfRG
5kxfIBve5D52S3UembI5GMczjhVlWE2xSuP82DRLwbezSSnsQnaJupEGLESvTNuW
UtvrsWDu81yjfzGzsOY0hmz5kLsnSqedWyluCuLTQwjVnhXr1oM96v9Mv6GPcfr8
w7GUE2p4WF3In/wECoiMrR7IsZvS3j3EDwfxXZPhVN4P/KSs7mROccZxOZNiAlZZ
rmIqtD+YPxANjgHxh5fieQfIvjp6tCIDDh9wfBQZDjOAF4HYbLRYRnHnMK+drxC4
azps/r+7f/Zd0nn6B+jQecclcoXWQm6xziGOJ+8ftW7OFI8WLDORyDzQ2eVycDFA
V1RDP8glaNlogI7F70iDE5Fxv2K29OBehmVf+KxBbovCrhQg3z4+pdF0QxioQWoI
ASaYSWKUosW7PendCmIp2ZEONyZViARI5OZVmhbYFUYzdkVLKMohhRV3D8tdnH5E
rhtrS5sip8YOiir3Cl1lCNiH6C4rhowotggw7frq9nJrtsy36ZVfWiPHSWX6xXbf
Mg7G7bLnOc3wM6wXpckFBBImKGnniSLDCvzQotFu/QXCuSPr7u0oEwAXeE+ejRR6
EhKWFVztnvqljXySFqRRweEfQBQzAaHjbzvSHDBk32v04HP10pgjS3vFUaimfNkH
gS5QpCrg0J9B9WOlvUl2HjWjaVaaGJvnnoPxpFWPZ7v9FDob/t172PZKSWx8WSFv
k6sfXncD6TNlPCfK2xNAJgF7B/9rXltZD0eWHzI1mC7MgkJJLKiKDPiWmVhoP739
Y0VryyazQfnfjU9ydFOrAZ4b3PyNfXcPGkLmoeZKTD1XQ0IMz6EfmxxkU6DzKJMw
ABezQhVKv64jBIrUJqx4BZ6lLw1tNb0C0GUx6OwqqFH2M1c+OafSC0ElvH/lnA1Y
jAPDmYBU1IFxkPloosel2wSbP1jRB723Ytgp77yo6SIJccERwbDyvZz2jdfzshNx
VifGQvR6nZ7IkEpNIPFU8nE33sraZ52vh/yYV09dCb42d1c9eJhdJST2so+dsOcy
xBLlpqyZDNxGIS824ELr3A/p5gTfbO7unYsDtyWmOw2UKE8ACo+9VETH37dVWHCq
WH/qyCjBTY1Q4n0G1NhvN7G5BnntxsQZWIFoHqHPAlZIyP3RaWaps21bDn7cfqZX
W/2SyrYd3oAJEqIN3lC4livPHWlRd2lhrfvOJWqS1YNIjYp39nubKwWglvWDrzHm
VETscvDhvXsawv0yFFejF4G+1bfie65XgiBdQyuqrZu4BTo9Sx4q+Dv8wAhgl1KV
aCBtvlSRPhMToqz9ow8JJSCGetR0wo5CZiUQPR7xOBZb7tOVhijYKhrO9xUnyDdi
XshK9pWIye18blrp/LeQzy+GEoYb7K6u0p0Spm/hWLMyrnrB0TJl+xoais7n1vio
Pqsftd7mHVD5hZy4mGi2VzU+YaXpGyXP4OJK7NF4v2CY7FAGP9W1lxOnEXw2Y7uf
bnTkAzFNjTq71WOYSNb8kGwaP93xtdA6k0e8Zv2EYymY/7d/9wdN6f5Rh433pjZd
tbwKFh46aJgWnHZTXF42A6tGGvdrxUDpmL/ZIRTbB9tD93bkOtanFr4sVoZwZXQ4
Trt7X4FD/4T/zC368Xyh36VogZz1r4KuM7UOigsq2akCB7Gv7kFgXC6USpGYNncL
yzGK9WeEmDd8r1TYMRY2hNm0HoMnLtXwDiAM8If5ggsL9vIzy+hJXPhVBp3do2Yv
PdO9j+K/UDFTk0fDK3mf2+BytmOlRKdJxUTs3Bsi/XDJHYBrdMtt+X0VOjHZ22ha
G2FPEVzLLVuykIVPcwm46HelC+nI/Nf8rPIyjKH96B+N4dJl34yLYD+SBpR11HZO
XXNkmF+FYRnJgoRUUGyCl4PURPEmibexRp89sCuN5Yw2GLU+uchwWatndI2n2uPS
FojT+mLDh96iL2rzpbxRss6P9yt7njmFK6dUQmH5rc5Ro7NLnPNgakxzTxIYQwLT
9OHxeu+eEL9UAtHUo4Y009t1P4y36ec80C6u12n70GfGRtfO25lZfnxNSgqk7PS2
nRqnIDPIK51FeJrNAjD4v8PUrZ/eWEVME+lgzcyAPVvjZ7ORSM3ul1oYqZE15qm/
4dGd9Wf/Nf+TYOSmdHZwVzMxUaSm5YY4jtHlIKbdogD66mYYyeeFgBDMhgxNWQyF
iFXkO1Sx1L+DWzCtwG/iVxRMDtftdKsooR7lEXoxeh2yXdKHBVFkaBcsEt0ZZYJs
YIvTVhjjt8JJVxnww4zfq2OMjtJfP3nFI77IauOKnRJ7bGBHRji8pC2JfCjqs4Ci
jNu/jA/ehi8oqJP8YjLzIU3IrMcHDfpnV2giRNXi6UesuMwvl2O0arCkX/Qj8gTw
jp7W7IMFs7fq9kPvWGz/LBgktq5xXhcJlk1w+fpp/YZNU8Vs1yULqX3giEpaD/Zd
JFewhzmMhvakLKdYZVGepFnp/CSSJMUOWJHujligcny2KIiv7KbU2tBPQcfozJZN
Hr5dMYb+CCXUGnBFk3srXDO/kJDHdkXYS9Boab1/hWlvJW4tN7hVEmIgYbzJBHmc
ggdGSdVM/YEBi1o1JUOrZYQqKDMASwUpbfAZnnJef6LYZeJsp4ol/zoSySQHpWej
d9wLwRnxOQRDVS1ayX7gGFQGJIGMQij/2PazkY8pNqOXLQwzURwFpTyUHKs0c3Gu
x5Eg9VHGfZ+sE8jqxfddcBKobNxQEpQSe0Za5uX1wAmQV6AMhX2HOnuX/USFdxZ+
zXF9psoeblKEWc6F6MW/m5Jg54UCYszieBqssXc4JYuVTEdXrE04au5hrpbgRY8z
CsKBE6GtZK91JnxkURdwB+/Hd8diPw29OXxrX9Z+bYuN+whJyXazbwS1q5lFPM4B
Wr7bycbTW//qmEzA4LGMvyr142S2f/grUDBqNveCktUHXU2j/hCQ9HIVxIvlOXvB
EsKMnMZjLwAWXYNByE3TlrT4eYVD8Cyel/3/HMz2ZoAkUQ2RedGFaErdKuYfZ+dB
YinPUBAaz2cY4yZylHAUEeqbAw1YVkbtp1INNdBEXGTmi2IHoVQ+6snVjK0dDdPa
1POtJxeD/WA5RrKlkI6P5i6+/QLrOg6pAU4bEWP4AnZMSSrIygfT76tqs00nqU9D
ZvvzSvLJCo53v5ipftQpNEJmcJXG9ybBCfBAyKqkvHzF6XreXfRPgXCShBbLM5c+
HnhkvBXreJi+xwnh+2A7vD81qcxQ0nLS2u5+xzXqrGoDj8UVGOUb2hG+BvoyuPAh
ROOuu7AWdIlI9UuOsGrh2FpUeS7OGNxHENAvnTKcG8X55ZR7KKu884cVu9V7c/mq
McwK/Th34o+HgA0MnpsE+YZ/QWGx/EqobQLKEmqAGa5cAJini9lJOr4LBDtGazvh
Xr7ENgIzZL5vDrqczjKU7DkPxrI5aEtGrZbYAVMz01OYvKcE1/UdJKHS//6M2mEW
O+Jp6vovKzTL2unfFl7Tp58p6F6ze2hlPzxZmu6HZr6sUS0isW+TRbv/hU04Gau/
xkmUVw4ezkr8qea8YMFY6HPgjiDSzKuDbgEoGt4mSJ7M7fWJAaqy7yUAlLQYqbU1
9ucZB2lf40XMB7gX6oREYrohDGUqHkEJkSHVNAbPC4oesRq9mw7Rry6Jf2jZ9qIR
Xg3YiBTIgW2ZUv8SewekpQCAzDe7wcznSO8NTSaWZmCuisEw/zaC0tZQguohLhWx
l4qayITuGnx3U9fRREslbaeQnAbtiAi2Lsd+rEYtNna0L9cLIJmwOCofdmShFCBX
Njkq12HSGh1ickjjG1CQqswK9R7jvtpxl6GyDJLXwnv1GttfgsPgOslFcZeaOktJ
VYOGi0gZ7iF5Jg/Za0qAI0fjZg8DXd0JqL6VFqkKtH53Ji7gnUDVVWsbGSLzrn/q
pDYfJGBRJAwY0OWR7A+YHV125tdd8pEN6XijI9o1Y2Age5OsDyL0PRhV2uOEpNte
WwYboNqkttYyfpFj8EIKddg+D8OM2sAWdf6pzG/wUHocou5Cj85yOSML3cZEP/IP
junXtCIj/XwJfZl8vPgICAmrXqNB8ukz21BrC1fQ+vQpiEThG6vV7qgUKBAbw17T
8k4ta6EzcweSMeF04YOvkeyTzBPwG5gycFoES91qLbnITHQ6cQdVqfx6GKuwbFWQ
b3ZEcSAVsjGkecKiXmBF0tAoCwHQ408g/Z1OezlV6E0XOR/q1Rq7d5mBY/83K38B
oOeqhkAKD6QS8IQ5dNvkt7NIWVbe2muDy4pX8dq+3JGSMmirfPWiA8+C4RDqZ70M
HS/zv0t7krZ1tzS1zSkyWHvgVQmKQTHMXIc1K5iatgUZWBzwGeSVXpClZYLJF3R6
Ovj3xXX5qrLoZDadEhGR+z+Z2MlXSmmVi4IO42m+8BRi8ElgnD5Cg2Xm38zyZNXM
NY3d2Ly8GJpebX4HlDpaRmfDNyhH43zeK6Y3k4inROO0uYAp3l/iBeDkii7S4pBg
rpvS0sw9xKdq8AR05YCjdnp+ulxf3jB4PgRYskgN7FPALzfDd8bkuMrXUUBxajbr
JimgK+52zJA8SNlpRPDkUPx+lt9aE9IubZNg672uHMH+Y9/opXCpqXq1jl19Xf83
oeT7TuMhE/UY3dK/k8k+Au395SVda2jvTS+F3smulDSRFai12Tys1t2tuMlP+IQu
fZW2vBEmE+MyVhZTOJo9OXVM/MGWaPp04Vn+/hisKPZ4du6myzdZOxUgpMpGBKpZ
irYeZJAGDFFYQ9vF8Vu7CLo8g/Lx4WCIJvlDoar+eeIRUvya9uBpBzNeTSpzLkkt
CTw0f3Z4d9QYot5H8GzHKEMIbgbbHZabT+/jmYzhXhb8K9lXk6TccdK/mOrgraZX
Q88vghK5IVb4JL8OAo4BGK60zQDEDtYA2UezO+WoagGSDty3P3MZNbv+F82uki+l
TUL5fb3RwTNzu2CV0oCVZpzjnyWugFes45Mhz8NbWll6oATgRgoufcuNJnf5Mtgf
PYYy6Co6/ke1jAmGmeeUMDBIseqbkh5e/cdMs3ET3RBgKUmiGbPjowIhAak0cZM0
LQtWmoAdIu4LDPXs6VJmn2pHevdjTAhqsN0+lu14eFzXXpbiOOZ8p0SWwdBoKSYs
YtytBSRAD6fO55/Kca4Db+uw76CxrclxQnOm4v58Gclspt1PXDUIJ0nupPpFUMSV
LIipwsrCbuLZqsC6EyJVGwnTb+hesL8oYl33cVP5q1XaWuVZXFSG70n/cvLfw+QB
OyUdhm9BS5IIzWbJr/kpri9tgsx2yk5WwJWcfv7xIx2q3kQEaOPk/GF+n1A5estl
A6lVc2gFvJ9qaNON3V1suqnFsjbgZfl6SGFvhRRO7CD5qRdjU5pXlJiDUonPX8w5
7fJMdJkNcRozHljfGkFZfs+rhnERmkTkG7bhz5HYC/+ejTtzstFj3NG1xNsM9zdt
+Yn/McJ+mQ63EOlCOVjAzVii0zl5STUXr5cz71UgJ70WS0gLnMH6dnbeUwX5Yiea
4UvkB5II7grsoqkeWASZcLSJqXtUXpXD2KKmQ8NOcN5dRIvI8DMRxurnUDhRWV4J
uNcj8+q/oe5grw+vZ30dkxbdRaAEmWJivtcayVXixD+Sp4VdQdmJ61ddhrK4txhc
3SnaAN/a9oT9cfcrYML2iqY0ifXU28svOpKeb+/j3pDTxZhpn3K9IGrOXka7ge4p
vakxScr/hmUp/zUtdNUfZ/K/9B6SDg5MXjJGoHLETpFn8fj0I59Ui044bVDYryk2
sGfz7C0/aqoGRUeuOEBPpJDrqZbUWWSfi9UmN/dbLkLkS9buvUeVwf6dYdutyua3
pv9srh1BWWg8//E6IIxpIIx0qyKqS7/OV65Iv1ScUkb67vCYlLfHCVo/eaPKypdi
TmcuXLZHt9Q6T79reWCz0wQn6aDbBEz/MrAsKpFmuOMH9PtyzTZUsslqtAQ+gOC/
3fCdEyTlBOV/CmKxA/yxYOR4kuZDPAH1qyb+U7whsdnONz9F3Ja4MUQiOWAmI/zd
nU4SFMcLX4nmQeRLTKGtmuDXyytKGE8BK+NKr3HBPLr4rfcw0QcOmK04KffeDO1v
9M+jm84U/GL+tLvlYg7UeBEqy+dvZpiguMAHSUcWjmwOOVvrM1rL83qlMKc7Pl+2
YZ8otVKWelH/MXagN0VQD8LbHMIn8OiSw9hY3xA/QQmUUQo2KOfmKQQ3HqAJGBic
5fbjoO9GFuWPpP8jjRczjMuu5aFOjWbtks4wQxdGeOUEqNE1bZSDYrQtcrj0fQb1
Vi0D8YSa5C2oJzLVqAsCbADuwFUL1LtOpas06cLpogHJvhseRms1XDQympYrlH9k
kBgBd70Nt1KnWvtsrCcmXHTQbtCquLY+SjJi8NInZq8E3MM+GKvrRs8pkA7UMOLj
QBip6X6abhoKO6ewSiDxah3BqQu4iEP8ItCe2G+NJazmsjjgNbXHjWbxr1G47GcR
Gq8YlaPOYDjLwL+M3Yof1lUvi2Qu13OnYwpTTGCLm0MZ1ZyD0g51yWLARQcG/5wx
Zveyr7/SxtkmuvVnmJYR9mMmICNZ2FVwwLiLFnphk6ldtNsJtCck5DaEkY6vnXxJ
3uR0UF3dVHjEXaxIPvT2Vsy8YxdFib6SZirBW5zZwpgiOHSvcQKfJi5arwb/t09Q
jXD1L/wYskTD0RoTTCldozoLfETF8ymZ8mDlIzMWLatTX6Z8syiYfDFAOiTz+dbe
tn/9zas/S7u3imyZabcoj6359PQuH1UFLKnLFnlJkjIbn0EwnpWyBJ5iGbUYqH8g
RGswBfNhlJy1tCmDK+eh7glMpgaC0Ax4I/Qs74GKRtfhrpAuQiXe3sNDd+TGVaCs
KNwHtUfw5WRea6JHPJxnxH1F8ADHLWdgSbyJJZsaflwiui7NvS/5kO9vzasDUdkS
5L+11PfwhvxupuK+Puz3nsAAzVWzfz/AB3dUPba0I4Uny+FWKHWGux/kimwcReyH
7JprqZN3wlfgqJN0Vit045VhdKmGrOEPVCX7NPYb/XssbwoUg/usz57cWRvz/f1h
9xmXHCrMHODwoVCTsfYmpyb/csu5ZvsLMHOshVuD5aRdq9qPXKekTtnsCn4G+ukD
OVOnxcC0zA9vo5wBA5fKjbLI1sv6ZKUE0ZxLur3aJYIwDYxrHugkIV+jZCaGDpCb
VFGigYNXeNsReDI2fFT3I6sz165udndIlH8MoAnQOjvq4C0E6El5qevoTSj/3IHP
fcovgSpCrsp9L36wkdqS/GmncXc4ZaSq3JIEYnVu4qAEGr4OdnKwO79eTCfcoEgj
PUyOBDLS/HR76BCs75QpT5v6OjBqQEHyGD3VdYt4DeY4mdB/avTkZx4oiXaYmTL6
NrgII6cT98v0oe0GowsKw1JskWDxnVxU4HsR+q/gzPoTg9SagnOubHP27kILkB3N
H1AZo50N68XHdUgMKBf5iEvdTVjNLNy3/7dLNnrhft10cZdP6kX4XVUs1xf7fQCB
JRCIgGPo1yZacZ0AL48dRt/2Hnh9VEUvwt/mrGfu3k4a18Z1AK5NhkhNfxuJNGJK
OgqNuvbTr0ApPuTSJvG7cioHS/+/R+wQRoxAJqnr/1v/W2BzQOEE2x0IsOvsugfA
7WdQP3N43AazPY96tuEvljtzP/NYdo1MkrCsXyf82F+5fNv6JBfKBrJrIMxxb4dI
ZEBAEotiezcdvV8E7atMYFYNmZxg4N4kAdPENVT5+o1odVa9Sgm1oVphkyHSTssB
FbFnQE09vRcWm9/+ZpAetwjBQjkEJbGD+oBXnATtVWlEYmyAM3EVwKJZIlotamTL
hpHrA2kqHT2+QR9qKBQHhH3q+v9jY3KFIvZGRHpS8eOJ/ceY/QBT4U7Min+ngGJx
7qwxxCxN8sf/yA6V1nun6YCHXmnh8JHeSqmHNsq6ycfUDA2Qjz8UO3q6M3JeJ2u9
J6Z0GVDo6m5jzk2s/QPtJVk4LBqLVwGyOu5OCOjvcN3FWHfOBUOQHTM/icv1Y6zD
Ei5bMosmaP3rZvh1Zv6h7KIvZhpKDjwmKcUfvcRhPjS/vuXR2zt5NUpeLN6ohn9Z
j8n0oI0NgD9lKh4QwN4+4hHxaq1Tl7snWSDYlNeL0rfwHxsm+SqHveNXGvB+s0Rs
u8mZ5dvRRmVCBvtX+t6WcmQ7INgh9OdJoosfydRPfvya9VXnR/pQg2NhJi1VWj9+
Leu/UwS1iG23Wc1dgVmBmpve/c5PQP3JefKUZ/enWtSdA8MHDqfpQ2zB8Szl9wX0
tzZyCjGQREFtwin6tf+wsCWJEQe4Xot8k0cQJHkiU45MFNsp0l+N1+GwnUWQcN0e
ZTyLWV0Tsj+AE2w2JxNYGQTdnVPXqe3duV8dWVmUmen2jYo5Y+Y7PzK9ZDn4s4Xz
7knNgZ8I33Ky5GgV8kEhN0+yj54/0h6nQtqv1H75PsbJIrUPzgkDb3bGxZSr1JmL
QUL5ioAJwOlUf0Gdk/OudYJr3xxJJxxCRCod1NaeQpvTlB+C4I3wRgcZAIVt+09t
blnCICigVoIsEb7hqmK4ruOlTJw1wldwEJqB8Swh8HFZhAJfnvxaBaZWuE6dVZh7
LirZ+W5FmMOF7oyn1Vo7puvqGLry1HZuIAeC4yPg1nia4y7ATGjWMFgyzGoU2vHa
6o+NE2XkNmPd9jNtb3cHiW9VGmKL8q0eLcaikninHmWb8SLdOHp6W79kaPTLwkft
ouT+1VWs7Fzx3zo3DU0VKiJpcrZmJKI9yVX6oMUIvguoj1u8nzzAa+C2l1gumLIZ
8/ku7Nj7SXTe1MGLEeH4MCxDEOHtVRQyYhvZ9Mpe6GJCyOZraV4CAzFkuEX9k3oh
TdA6nzQZdzvLH6OaK5ieQd+IhlgV/Vf6t8RsFPvlZ+Pfy0v9ZsKMAbLDEAbI20NF
vfSjqQpziB3gdosHdymHGBw3ePAPOEbblNI+5wPAHk4JYzzQ4sFpGclCDPjSzPqy
xip2UnYqnEtv6FpzuPCTdcI2UtTknE6PBYFYAqyNe1Y6bUiXsGv8S6VUsHSuRKu4
SGoqjxGJLy7IQRkYXeUBhpdqn8man0Y1FxQ0+bIc/8b7qND568VTfV04mu2FdskZ
pObrM9jO3Pnc6KBzc2r0Zko3lHNLZaPh9P57aejlhrbwzNXnamWgtiBWZ7MM1giG
VK3fFLCfMTpG5xGOmh52MVklbIOIkfCOYF+aLGqaKvCbgOFoc1el0MLTeJrxnh3U
DhS/tiWsX3CSkXR7pXu1ReQkBG6sKcLxFJNygtboMF+cyNchXIdj7mQHMbh79BkC
7+JAQGrGxlx5zUhjJa14ZKpYX2Ue+3LR2v43C3A3YUDBAPOk+ZqTIUWaX7JJUyar
p9FOuFCyMyrrHvsh32ASwZpQ23E1mh8wYPy78cdXW+O/jXlzSkhmAdkFquqAms1T
PshzfDsTzNSXLH/lTtNwLqeKK+A2NaPfEX0phxZoK3Wo22W42YDM74iNRqgIF9uO
DSwMvqZ8eib6VeLhwltKXC2jUVpd3l3sdXbgkzoGiFCCsEG/SiAXawk38B7B1aIg
rkQ0VZwapqZkT8DegtaZnv1XF8VNRHGkXhMG/F6pSAniobKNFJlqcj7nWiUG1Gzf
5twXwvb+NGvvQPqdol4pi1ZxF6NUN8QDqTLfAdVmA9I=
`protect END_PROTECTED
