`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eb77XwaIN1Y0wmpqBKfktL22eS+X2SVL485Kdx6Q2wfs0pjPJbVZSDN7EYfDI0Bu
I/6OL04auuAyVPvOpQNKhe3IrRgXZayemYFgvUuD21kW4Jr/HKLGmJLYxUgAo2TK
E9VHf8s5O2gjQReCSme0TIVQl9eKYq3yN5SP1e41m+cR69ceoA0G4uRrv1Etp3UU
iHzeUCXTADkhZ0jBQwgAHwrzaDWxzSuX73q9j8UCcBaLzv7A12zcml/TIRAtWV8S
AxLSi5rJfIM74C99HTvAiLHhRGkxOqxpxDAcqMyElffhmyYxIu0yuSel/g8KwSGO
zdiisTKCOxSMnigf24VKXClLJdtrB0s1U04jATMRj2YlPUpP6aF3x+RPKXLjJzI5
gYq/pRXy1sZDMQheJ5vOExmJHvSxSh8BJNgjRKVL0KmZ6RDp12eU3FmP2JvGLSNF
HIjktd4r2LavTTK2+OVcbwz1kDQtzE1xjAEf44ONFRFjgHNy77CJbk7A5sfwBX0W
76/CUwMYLz45By+9BrFzPKr84x93Rb9mKYqVvbR8Ptk55Y3a2MuOr0bYQoCsbE2R
cKYtwoR45j5iOoMSm4WS+7cHGQILjrQGZhMlHPK/CqEa+cj0dyruXWDDr6ZMqj0H
kk3KgNxWOjnMAnJrbJGBXVO84GMddFXm/X1O+wvRDJWrGJLxnWC/j04fD4C2GwQR
iou3qx6NAo4lFwi94UdQcEONkIP6dGHbK6uxkKpDjZT3cvNcqib8tKPZgaxJwacZ
6L+GAoec4ed3+zpHb32ggQqcTKSR0nInkPmfRdhw776jUBPwDpjT6MB/Lu2+mJ9H
blK2ZBVjPFGYIWIR0t6Ujg==
`protect END_PROTECTED
