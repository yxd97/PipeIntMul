`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kwS64MqZz+PFlSYDvOV34MERTRVhTNYoTHf9tyw3vxW9DKHBODESWwleFh53Ysew
nNwEaMrPZToQxvozDFbh183HCBGDPiVKAucBkmtNd0+gjYOPaVi6lyPFZBOvz2W6
CW+qRJtg4kLD2CPkgUzXGIkk3SYr0tEBzTPLYCws/GGyH275FlnuRiR6d6pMVznI
cOi5b12eqSBK7V7BuNttFS5Wx59rakVRcutbYkXS1rLLH80MoC3K1JGqqKNC7wsl
e6clHothwmyPujLV6CnSeUSk5vtgP/fA6QSqiGVRGp5A3pzrjz0Sw4V4kLLww0nw
RardJy/VyK/pBwE/xMw35AwWkx8mShxZHLVge2ZEnYk40D2cndCOmX85EpUOGpzX
UfZoaXNHfYPdDkE6Cnl4/JvA081J60Yk8e5QyHL3g/k=
`protect END_PROTECTED
