`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a9swo2EoU0TzX5zQCvPo0bF52pY2iQ4fZfVyVHSS3cCICUZV02K2FhaTYPlj4Io+
zDyzYGqfCTTZ8aqGn0d3oUERejFyc6HGnI62qFCDE17oyuZNwqtg1ejZtN13QIpf
hrayXrpNUsvWUnuh6tU0lQVzrkxZwZjUp/BusRi0oyZx26wPPFrnThuQOPV0+EP2
6bfZ0IRP+bQeN7WqX3+aJtR21yVAZdGjwK5fnSAgZPJU50pKkDQND6RRDzRUjX4Q
8hp5264qht5OPtfPN9wVGw7j+8H/YrgXygudjkUX/IDYsN73qXqjvBbIaCpjYClF
TNrvRsOVXGr7Dr4gyRUCrLPxnv5wk+BL7EGkQjvI6CzhUfyPLoLveCaRQ4Vx0/iZ
jIAhDldywKldDWSTteKAmVwmiKDHIczfud4oBJcwhO9Io0zdnjm/774Juzr/hbzd
qwtCJaXPp03f0d+4xLVP02xuXWPXtaAADaURRqEC6sx/+oP6sAkNslCCIREgTEw4
/D5+/0j9OLFMssiSnM4BBFGkbIleeLNZIaEYSPHOkm4AFylR1JS16W3E7ZeJ/Yx5
566qimd/fVPoL+xk1TEILfjwV3C/vRMCp0uRPGrtzePowuFsA/iWELsHaOLKAMxg
0jmGAHboFShSs5SwecKWKHQObKrCvuJKSYXeBjVKy53NbeZ+N8mgQ2v+o9bDZOn5
MQb34KP6M97eeHRG0LGi8VO1DJN4RDGHmLpa1DDWmIq4cOrymH2VVCoPP58fnvnd
PyfgGLSBqr2u+6304oFCJsGHx6dzZU9ne3rhdFjB5oVjD+CJZ7KNTFKuRqk+e0DT
0fFOa9y9cvKG3vXTJFdxoQp3kudDbbk/+Y+WDhRDW+2Wo4yyXyF/WRrHsJwn47Cj
kySStjHVi8MxORNQUFtjsJnO2Qr1ya9t2jOkNJXFV6/YaP2HTYB8rjz1SZZhZtxv
fYFjaVujRH4HUfEEj/2KCZSzO2/qWpXf5uVpwUQOTFWpPGy/tahKevx1p/wEl29d
rGGx6GVoASjkX+zKQbbyeMA8tOW2u2G0Cf6LcE9sIwGuoUeI0R48pCXlIxmfdhQm
7JM3RYRF0ZRHK/F/a9Stq7jwFlF1qTqKCJS5hLAAaz/ikfdZvcv956EAyACOedct
qpkpK/X2u+yIbjQ2AlY6nH1l00k+H89sMGUj0SlHKG63OdyXVXhWa7mkdtZz51nC
NcY+IKEsdQvXIF1bRLc+/AJc5UajehLz/uEE6eb9Xw0ZXVZVvpIBJf5wvHwMWor+
qTI0Rpv4ja2iA31jk8DRERj0xqTWwdt5GREb4qZaFlkYreA5Xpx17blrVL8VaywI
iYRYT7wzd0oO5sBQQhv3Aru4s4R4gEajA4pnWCB3nzSHaer5WrocEDhtapn+Fqd/
pVyDEpbBYJoxx4uJFhlmJ6VbEIKj51cE5hovwBkxL41NpKe7etJSyMwvO9T5fQqY
cYjLvrEJT5A1jECPFGRDsaWWlkpM8I4XgVh2PBx/8xBjeHW7VZIlu+LlVXVfe76D
OHaHmm3FIEQh59R+gYxlhx8nMhcOlZXXIvJCgdtGpGU4v4VNiVHykQnrIBLgKbKr
AKRr85MR7eaUFm6yfstiIufeHHQJMrRra41kIgYGwwvUU9Bj6MBrpqY91My8huyH
JSFm3WAxZ4urIkrKxM+4k0i6D2o8wgNvVuvWaIF/SIPpHSg4eMninppCre9QIOWQ
kmj83iM0mOUVaPyZurupuTGL52DKWSu65qfjW2WhLsopC85Hf50e3bpLe7fM+ctU
9KBWOQMJBrc0h4OIq7eeUjtvNohEQHAe4FYPmp5dIklfkruryu9AhowjHtwFTfUv
CB2e5voGLdjcr9kfHy+M3nZn8OrRpAd4VyCjfDRDM5Pk5C1bd+MqxrzSOi10w7d4
5OM7g4EJYSdjafNaP+Bjb9jQU5mK65ySOuUWR6L8QmSpmzxOePJOqbad5QjSBQ39
B34zxxgNWX2+Y0QdRu5cdNdrOGviwVFNrCXztpWxyJKxvIve6Ycmf3a/OIKccA+n
gZCLWK/Ahhedc03YU9vbCr9KQQOrt8T9XkwbkIVO4mjYkFQaCtxVNbqXsH8WTIqN
8m9MvHeFodwFDj6pOkNNOgW16pgFqIAbyIBLhFqVCntxCQKb3tYov8sR8jwN2FcM
MPdwPW6kNkFiyV/gLHJHvVU33mcxlgLzpoKa8w7n7W/KoTBNbaOnk9Ln3FmAW3En
vEO08eWzrYxLGLV53qh47MHZWNpptcvS8qFEOkc4qT/eMxEHHKvQY0R8Lf5KHlKr
wsj0kduZkcVoIKTstGuy4sVR7I1V79CbhfXV/LrlJT2iEBU7Mv6yDtZ8xyTSl4eo
GJeRGUos4Mczf5FqNgQIHp8JxY+ta/IwG+4gzLCiyVC7g20/XujQdsYCpv1wLfwz
419AVaaJ6mbDe1/de1WKU85soEBf/CrclLUEcpyI225FMBBFot8wVakZZQrEyYbZ
L6E74goVOi36qOlDkhQjuU91d2ybishzibALk/swK88xbF7BWr/IbhAX5qzSqmcQ
UYLeuOn3/cavuvypfMbkVdAAlBWf/H7hg+La3wHagw4WqUd9aghbFrWSDU0rMJHV
qILMwJQfJaO0/g/+r60sf9lkmmXqm3ywBgj+KKvU1MI3VcwPuPpjA50OUIkLSshC
nngPj4ZR+mfSr1zn0rBO1LNlQrAqx27pkaCHE2cCJFuHIcaXWYqlMM994ofEsbV9
bklPc5LV8XTkdh7aAiL5srpK/2scOcrlH8OByNdtHwvEo7EGR7kE2vQI/keZNri9
hyi8ahlYQSTudOH1pqoOjL46XK+9BBk0hcLPrEUVGQA7yGCRKWWtdbgvoeFs6UpY
VuCh4CPhsgaOokfKauftsL3JnobCav43BGJDjwTAPw5/WVG4OUUUs067vZCd5T3i
gMnyB/+0bA6N+ACOyh1Re4+jBY6eSxKXM4+C9v+0DPnDyYmowdqJPd0NXgodtktN
rWHDT+gs3P1Yo2Jis4qMSzGgRrb12wKonvHNql60XPgWP7WrWZHgVt+SmtMlr4TW
bEXZHMkMMPy5kh6N8oldrrToFcnveEFpZFmXI+waDP9Xo9BmGrrA+nGLVaFo27bN
FPsIBwSR/I6AugkeIc/shZfQfhkfMMP0yRKXbK9Y9w+u1BkN08tGgwMltLXijrmq
G26+jCyEiwQmh22hmOeJ8URCTwGaDj/WFpxS92rNTiZaIRux/nEvYoTAtJ8vicDn
YTypel+4Bg5qdRnIwctf+2h77y0ujlB7ULHdViQ9rvz+U+VlkBVJdOxCxm1/ObrY
/U9IfweuSsK++79k29E+Lby5Ip0t8OkPybQfYdpcDpbAuyYBmARaSfoQ3oQSLOla
H9DzcNnAsDwPFaxEl0n0W1UY1r0W7GG85UOoavp14H5vAWlkmn5vbU7AmYc6lvxA
gPhumBU5CxfOMmMYFz72MSZw7KutPLoWH1r3lXcwaJb/nowUKgetsIJ8XNqWGMLO
Jvo9y3DW4BauVQo2Qtr0mfVrr/UXY1mmY5PqkV/f9Tcfr4PmyNVnKKu2CCUKEPwr
FTw14JnAl852qgeW7wzPaTlsLp0ltJ0O+PdRdMYMmV0Uwkwwzc51qBXqLnhcFo2h
aBQOF3Sf9j864qVo6CpuS3yh+wJGnEpjSv+/s7ZkP4eD6FnQ8+kmXNQpcjZ61V+d
EsS73jxW1N/yTDCdIhY8FpOD62NCokOag5abe2Y6cV82hoi39d3Z6VF7IE+7X/5V
Uv7IK8XOHC1wXqnsKMl8cUV2oJYE8xPzDdH4c1nlX04AThAOCoddm0hZUN6V1Xou
G6t0L1SWVALtO/Z1PGRrm8s8KJlbiY5oJLAofxO79/I8O/OD/vPwXepXUyUGeQr1
c1QnCFrhlePBdVTKrnKYe4f3fKeqtco18OG0001GsvycyUnajFpgugAvWM4seIOD
0XrUD0Oz5i/VlMbgrMB501awJy4obnNEFcPl9Ih2USpAysSqE21nU6ixBYCJyWrl
b7Y2zI/S0uJSzCu+R0iE7puQKmTZeRsyT2Fdu81+dq1ViVShxJdyBFzaesm0x3Qb
BjlR0JTCFhoBOtKzLxjbS6luyfbSnHhERCUHMzP9PuD96Fg5prQmnhiKKwO38ts0
NU2X7TK02im2ByanZwN/n0CRX+mLzZH+S52zvs2uVL0msnjHaiHjPS9TdlHbFt25
VlT7DcRyyqB27t3YWJYVAqUndcPfqApJvh8GVI8XH9aFGEeyk2O6hfty3sUbGOpb
BsREQ6KQJW/2TwOzZd8Kj+6ke89TQ6/graOSwCuEO+uL7VBTxeRp+bvDUqih7eJ+
qcz4ySqdcto7JMj2DGcStvtmYugxlbbLCg4aaLIMZCoYSmKg632Gw88HCw8mV+Xx
yFk+r4mr18rY4luhZ4UnHZ1wOvy8FMmCnLUPrKv703zJt9vvf18xs7P9tm5Nre5/
GOCGYiwnj8E+9yISEutfXkCdN8WNfCWmXpkndsjBJPb8urb0PsgGqzovbRWswU2L
J3008bGnvWIQl56LW70pYgJ9g7bQAbT6AjjlEafVebJIRG0DqjTtdszAqmatpgvC
o8AlgEnsFeO951tV07QOujVcDT77lLvcT/jJi63+XBVKJlm0o4qTkOpr1ogiGMdc
7An+jcS1gJu0wmCOcYtqRJE3j++xaeIXGA7XeVAQ9Nv43aUB2Q2Z6z439YnOJJ/6
JlcK6vl9P/iemx/iFbS0V/vYs57xhWFa+D0KZ/1WpSRqEAOveUgED6q18BHbHFVg
y8tPkP1N68KnNWcKD6dFtH+PLFe0Dij8uUp/MBwf3BUF+9UKm5CflW7EsrEna0gK
kH76kXIhlI0kW7g76HRvvSOjLPnPojzuiCF6ILcK8vPUP53JYRe/jVLySC6thT6l
J3IqD/Dj7ufgSE9twAjlfVjQ3GQTrAmhmWmR/LYOFNP5V+ucsdQMGYhvB19fk368
Hhq4/PRYPwTu16Fd2+TLEZx1VYzQgRHK+W8o6WShLAYhcmcdzbBxU1ZHoEU7TH17
0PCD8iwtfrlfg+Sxd6duRX9ZmhOYBcU+D4RRd/CqHidKce3iScbqr7w04L+Qtdt5
oWJDPjFj7wUXt226ckx6qBWof3PiLf9V7FCEs+TBVDeL9BdeU+O+YSaPd++JiyTA
47Qb3BiVqoDsKBPXG/mI+6oTEvo873pvw4YY/tT1vHlVh8S8r94te/YYP0YHZJbf
f8D7D/8SgoW/14HID3MOSNd+ZBUWPcWKhg0a5Spsu38ReVxWYAtKCZEXj1xND0b0
IBKBiov2YSr5NK5fZcfhdoyBsktuL9rkawsFoFk6G4YzQ81Qgr3vfv7G+C06XeTY
DduG/EwZrlBRwzmxUED3+ST006/5Z7zRp5UfJtBlKcq0kWqj30rQCC5T4WWz0c+W
unf/YOE7pOBOmOTM+P7cYJ87uFnLuG/VJQB77tEOzpM7Px21Y3uYRaTupXPMoa6L
c/PP+/tKj5JbNEd1fdO4r2yDEkkypE+1P/P0zeJjA/4JrEofzxLFC8QwwW0d4Kb8
00Nn9lJ48lTkgvrcS47skvnponoq8ZfMN/6YuVHEBr6BsrqTYYcaclvjfpvVlvm6
JI0ZUF7t4xSw49OvWg9Ho9II57q17YiAqrXDoMEk7+4f8a4VftMmJQWJhFIDJ+rw
mX3VgHiohRXjUWd472sS76SBCkwSrLYeOKK+dGHAWWd9lfBFlBw8sWoJdjNpqSnW
r7TM4xWxJtUY/YIS9Sls75FoLtnIxLswBKs3y1It308w2Fm2A07j/yRDKqRc69kK
KRS33t2QPShq+Ghfn9HitYIJZ08Z1fXeP75oYLkhzQSkncoKYeOpepJ1qBKOBiUM
kAP9FtrQVclZ5o5jmOFMs7r69zOXchw0tpxgNkjJ9Z3pxo2ZwFG6kSi4gKF+fBFG
u5+qCf4kYQgyXzsODYECXQ7g1wILy8EmeFFqEDeJj+kS2FGn8NafYWgOHTAJImy0
5JkilYVnG/qIr09OoWzDEg/aT/t5MoCk1219N8Aoi9DUXvt1ZGf3hw7gmfXqLmQS
ZSIg55ZujR5fWH221kVkxFQFhvu+c6HIDTKsANlNTWfDQp9XszU+zwfSQZZ/RIW+
ye3pUTtcr1LmFAKzqDcLtoGm2QcE9T+9sh1EgL2I4R08TOc6j0pE0EcST4PJtZe8
rO7hQFmoHqQ0bMLqYu6uChz61B63AvxjSTQhETbD56GoKxsvWLnm6ocu32Oaj1FQ
qA1yCSCHe6oP4kVX5Cd0H6CU1IE25uOoatbu+iMEWI5xQdZ3XRgleJiyooeoJqrd
UgZb8YOoenP5BKgokIrga00PShh6WM3DY/ltpjM2sSBogd5MZNAD8c5GQ0jdM2Qa
`protect END_PROTECTED
