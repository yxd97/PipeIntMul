`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A4xCMIuzRisw6M56Pz5T5zpGF8cJvTPHWx+Y9fQ5dN2arTxcjohMqoWJLRYa+SvU
P8LEejJeBhn0zLu8OmXjWDu1Ge5ApqgW1OTzuF1N1hxxrhuyHiLPX0M4MGgilzAr
wmZjNlL95HmBR8+Au68Aw/25geOxwuZ0+RyIjyCwzSKLv8pSaRBB8eBL2st3t29Z
bmon4RTo/5jUkSAr7OY9ubnpXc0RwBGrb7YhyF3GM9cyQGPUFSN63YQwsS+caw99
dJIo3PihW1k6HKmrvjY8NWiIagAhg5ZKbn1LqugvEPxdYCcomDqgPKFFvUbVZdOo
58VFddN6Fb56DkSU2hbmZQ==
`protect END_PROTECTED
