`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JzD1m0UnPD4i2EPmVHg5fGskf+dCOVrQuCR1WJbJWS6BrQKHJ+A8GYvEBE18lhfR
2BsDlZp2UbcYtR7nsLJ+r6MC8F2tMUihiVB78lYtHfVUoEgbNfGiWGMm3QmVzXsW
Fd1Ji5WAWHYXQoGkdOQty2AcKkI32jXsA1gjqPX3AXqvPSdp6g+dj90cy/fbScFU
4V/5l/0g5Qu3hKFoIYsbLGjEteF9/IA6IRdhUny4qGF68GdodtDcJl6T/BTBbEkz
84Wza4/Sr44fqfIPaSr0lLb3nqzPvlCkUO4ehn+sk1EG61Tq/dbegjcG80JA8ef0
47RdnVuU6xU7pLbhbTL53jMx+ycNkljPyb9WZ2VkbzQUUKIZ8W+9smH6brOVgPc8
kR00eaxnGBT1aWlfxSRvWH1YzcXrieWde9Wd+5zt/7eBdEbEtaqivn4ARCsGhPn6
ZG4HAvvS1e9QI5cFDzcJgHSv0VoFfnVF0gmOzknRJQzknzO5Td40mMREPcZKYE7d
JOMYv/Zak5HTR2OXMjFBL9RZBwEmlTCWm6Hp27BSSLjEwTLh9mYKE8f8NIoryDmf
Vn6XgRh50lgWQR7ZxTLtXs2nTZCmrPLU1o/SqPuxqikNqeWGVGJz1NELW8xfjNTx
g4lVZgTi9WkTjE3hHMoeoyjfoumDNK/wbt4kxc1UbpkOdsSzSoeWkFf1xpcmrfqt
XHJ08xQNFhFibiv+jOaAnxUr+R6RZfbax/NLAafqMMO3eVYR7CgH7cptNipwsjnd
VnCwshXtJk+sY8CHB0b8ZALimcP0cmKj1JesXoR1eu3bSxsraRhVdtYtuPGY9Zh9
H5KO2dzuqICicZIp+y9q0sFJrO3KytdaFcADkXRwK0Or342FpGynvGXaiNTh9kQZ
Y1xQ4zNZG7Qlk3c/Tp4i0xlkontI8wcUYNJSzKT0kio0cYd28+ntRA0BZ7kCRBU9
a2BDc+gU14rwEteeEiaZ9kC57caGwUYBVMcNDn/1WsRZ0rba7yC/zdGrUvCX5vFt
ZJyaN6Z9fnWFVfryEbnGIRaLXD2YjuDQUpbl2nluyjxw3Y6PFMAXQDINzm6zBY9y
a3YbFJ3pNI1pCbsmXs8PudlRNoWXAhl+IfYHM7I8hvbZOuB+4s++tjreZEsvhps+
Fn/gpLl4dcW4NeYfYJVWfEiX1Ni+jzWq67hLyeKjEvCeWnnJPvi5VBeHbooWYIG6
mAnmjTquT8TN1TgvXxhLfIKedUiKR5HHOHcUYfsjkePFfpASc8gBZtjN/9+rTmuV
7p3kiwZcY870lBlpQDCa5AKnk1sBfTJpWLirKbk4LL0BBJkezA1YxhVophOlubVp
PYNHzSTWmgx27+PeupjMxL+ClGQJxdScUuIebQZD87zo4e/cuTIdW6i116+pHZVW
EXBjv7DkD7STG9W/4VzyL0rAcVrU1kStWIRVCTGdu/ZVt0ZLVpSks9IA2PEeHbZz
ZyigEF9ZjcjXUP1gmbiPgRyop8ZzKtUr4Nm/Vm6T6SK5JiB07lTN10LIiVrWzvjg
CfrbEWBoszBj/sSYp0k5eN9e7IY2nJWArOYyNfC9A19C60in/pS0dDdy1IvPqFgz
i0S4q5zvcFlGTvJJ9Hjmjzl31rgjfT/qG/u78FBFm3enBEMdGtFgOJBW+sM6jgvt
WLtVWKqZrHoT6n6/j0q7PIEl5MH5bQFsorLj36VRvYRQvBNdsFgA+3K/rrynrjFJ
oDu1BmahGAAbJHzuoCJgWNP+zKeq/Tm9FGtfEXUCrbQBJF9N+hm/uwYKnMO+NEwJ
RzFwXIwTxRfhFZHOYpD3J97J82B+lYvqHMfNB7aGLKcbQbIvmcHlKjemawWIhd3i
LeLVMJzYPwIySgIORE++PyM6K/+U3fZ39kPRhwDHByucrMHUbUa2TPYew7CX6pU5
cU9OnF3pum2EcKG0lT8GBpcKebtCgytAZ94J8u9CxIUOVF3yi/hycpbAkqCtdoQR
E3jruUo7+Tv86zz4e7IcUzZcA1i3cGPEmUKZQaDW7Qa4Ou1POY3ukAtNsyNkAkOa
K+a2nwqHUjOC80Tro53mHzJ/ufYCLi52DdvRM0gbSg8=
`protect END_PROTECTED
