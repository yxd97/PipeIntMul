`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zx7iQlZyDfizwjEmk7/licBhNsdiiBjBKnEOiQzOGRQEnat9Pzqx4nwqUmsVYgyD
nI+ucW9/cl7ai5LB3COaIMs5S9SMaBaGhakH/ILjrnBFGfy0fCkWPlP+cxSbZbLE
NY53ZGlftjY0bzgMUtIR2HZFHM0ItTz8wYfpyHY0fXwj4PZdvGgQL3pfmvqf6RmT
cV4U4m4oYodWjwMVQM7nsaUIfxas49B8qGAwjlOQMlmFrgjwobRC8zo61Y0wljSB
OADOHfrtzRutPmuZHxmKBW9Ld0zlCHQ6WtC2vRleQIGRGplaAgzOLRJbdjyUpTlx
HTBTGvmq6uuLi/9wJ9HVUJTLS2ThMQz9EndgmENB+mRt64vPgNtLLBMx+TUayHeX
YMeh3yKMJ2iRHfDxQidp1bLhtnwtW844f6f3x/F9NpPT0afBOUFM7hhW2PJcDef1
lpBXzA+wpBKaUVYumafUgu9s2x1QiY8b9NqgzKoNsoqWkdRbAwj2+F07CuOjdfy4
cuRQxT8S9B24kTd6mJlqStJJiKZX59ZEwDBdmKpGG95RyAfr5xwzdAl9TMkUMUeK
CoZOozwMBxNNt4MKML948YANuJnoET5z4IgGd11DN3NodCU8o4tx2oaPTH0a23iv
1XAbE8PtjMt5zRwxKTDS+qrJAHRGyCSUEqAnwwDzh6PMUBJJMLQPCsC2+KuSHlAI
b0xF1rE8UYuHsPeFTSww2fEsIL/dSgv+5e/c4EeELyrDNQXoOYgBo074cYo8RDoe
S7IdyHrNH34Tmqpc1QAW2XE8K6N5fO94bxSTeNqbpj+m6fyYZVyQ8v/JjAfsdFTi
yS7ElXH6o7fg8UzOkDPCtT35GXKSXGctLu2XEhA5stJMQMrbjQf9uA0znhP9wJe+
5Fi+vTuqmbG0pniGVCzLcWJIbEYC+F3NAqtqWOdSY2c=
`protect END_PROTECTED
