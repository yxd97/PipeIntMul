library verilog;
use verilog.vl_types.all;
entity dcm_adv_clock_divide_by_2 is
    port(
        clock           : in     vl_logic;
        clock_type      : in     vl_logic;
        clock_out       : out    vl_logic;
        rst             : in     vl_logic
    );
end dcm_adv_clock_divide_by_2;
