`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
isUJ1AzUHXexIutj7R8fSNUi4BL5tB5Gj4kofgo7fTuW2isFq+V8i3rEJmndkmaK
4dICWzCu/WvrhpgLjoCkEjygUOEI38zWntFDsXD62xGVagm2n1iHobGIDoDjlbpj
HLqjBrWh3w2NYKfxVjtXCSuACmr2E+KlTycf0veSxVVH0OVZnBKVFLdIapJ88ACS
RazTjGKKwsJCGsN2b2N2gjx0GnacYJkvKCmsFoCEBWVpVQuUSpuh+GFiTeaqP/F2
H/dM+fleS6CHYHxTzBZOufk9CMoTgRlGciW3aEtqxc1K8QqKyX9wx/H618t5VaiI
7fKz7We2ixbWQ7RmMyIm+Q==
`protect END_PROTECTED
