`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iq6a0LAIJv/lfaz8o3XXeKpD/GJKavUujpmHdU9CR6rWbkjykk1XaHE8amwNHlCB
5mXRQmWktxaVRCduYpe5vjX6Typo656cuM1zkRpIkEXDVz1SLxe1b/+Zi8Z6xkDE
v+vK4bljdri+Wz3qTpkq70BVLmkr8fp0CH+GkEg4Pu/dg9gqIWRkGzbZPNDnCeFD
dm+wH1LSfAMbUdAVXxQn8IRITg/Efsdpsh197RXcrr/Jufg6qxPxfIdR2SFY7ZLW
w0d90poSRg4aTdWIIwJ+0+LVNOJaYepCdmSWdQZtXf/lOQy7oA1ZpnCJzDmzrR24
FWXMghU/p3sDyRH2WUu+FHTuNBOH4gwzr/Npbiy+pujUeYBKf+Mr3jNbU5SMwGxp
QF2RJ1mdZNsf6Ki6Vja6Oyhkq2FPduTHN1UYCT0St8xX2Ni1l/PQZTR9cpXhpL/8
/o6I63DxJtYNauDKLyCK6ONX+bGqsZExbpBJbKxCnbyMYt/RBq31ad+dmVjG2W1U
N8vrOhm10+7Xsddf3mOKu7vXBr6XD9G+lyBlfExJdA52fy0t643GOR0ZhtPMqRxn
gYURoiJsn0fxgC08jubR3FbED4VyzhubKI9gjMYqzyMtzcDS8YPn77J1KgUzHC3L
jGc/plGvvBOxpeSoSHGzkozy/8MXa4EjolC+JPrWxt2rf5FaBiZ3d0HnMvMzEodr
0b08R8oX7RrlFZipPzxx74ja+6D2CC+mbgvQpcNxAzfoVFUwptN6LxAFjtBbfSEU
CiTom+B6KzU8wg/ncL43+NQQnk9/t2Md/HPXGTam5RWE0H00aeYLF+EuhpMlBcAy
wA7XRlYcZoTw0pkdyZx2vXyewbgmGL3OUXEuuOuPVH646blEST+jLhzE8wC3uauO
mtlYPKWtytVHHkqffMg3vkLj+WZbHcOaTXN0CThaY7qEOc7dPrfbV2roipMCQ2xQ
ar/+PLmpmBTtt120I2McWKc5+Y33knk4VUFr7WjYcyaWN+HDO+OlCZ1iisqFfAqo
AmCV4MdyYaNbfqEaRUmXAJorwaSO/T+eUKt/GrFhvPnA9X6rVAcDIVvVg2W/h9HS
4Z02/B8o9WBr9aKn6eukHOjTDYi1SfsXs/zDnJE5d00TlyDiicxwc4jD0G03tr8D
y5UW6iEvJdcmaAebkmJYAh2qwMX422SKblhuiLpwxGTsfxChuQaRHeggXEsxv3NT
zDbFnCyhQeBD1FiDjyiR7C+01qRxcB+BsrKGWN+Fg0B9/myFHJAemmk7folAf1yM
62kbMD78iKEFRdjNevf60S3O3eIAzKyUYjlonTkFknA/VZzlULfHPi1pNRIEJ2d3
xtzPj6ilzkf41pj3w1UFCd4X9pK8iBxYjAmpfaEeX+TL/TtsoZgylLHHyw42o6eV
wJAM7XhN56OKoF9pqcCwUDwYUDnzxVwvD/9r1Y0PjqNVdcJgTuLihal54QxdXIgF
vlclb2wNiIigo0ZdjoOkJLHcUixBhXb/2rtzkow38UnGKazGq2xkg4POWl4fzVcm
tfnQyfIfC8OfbPMspioOK6+r8iKskvZDk/Kfz/aDYzo=
`protect END_PROTECTED
