`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QqAinWCrTkPqU/QQyU4A+bN7giQ6LG1v/VBbetOkTj1FppSTTIYqgTY0lqKG9RW5
blRxcAyiq17olr9AqgVHc+BX2xeF7CeYPpWGJnQwJHYXdis7QYcDJqVuhNdmkP6n
2XszSbU9druPm1yTSl6EevxnIAlaP/JMQWFeHWoxW1uiZ11y2nrx6vuQhnlpmB0R
I37YeEBhG0x+1wZ7z2x1GAPk8cs69e/JjSuUcTNL1oF3hcDVWIZzmaCoWhDYyu4B
icopC9UXHfyLbznP1MAIrWMW7KUW7yLmXl9ou/BPSi2bsp+Im7jKhlS5VCX/xeuY
dS5YGnHWlRHRjdsiKIpgPIc8LFJwXQN96c4phjw7O7Lk17jrv+mxidCJT9vNqdLm
oBdIYxkpQOLh+f3Z+NUb8iyGMKTP8rV8Dvx6zysGACPj5r+VPtT4oq6JgX2I34XH
1Ke9y5UFALch6PFZFFGs2Bk/a6fJ8v+yD8WWclihRt7kiZrfHAvGbehvYiKQJHV6
gmCEej1dmQHsx+u3CaO8H6JqJ5FaINfoUVUdgLcnauFkAVA3dDT08Xg8p7xIq7UU
EnQnfBMNJagFXWuiCIqSyWpf1l3wXRupd0vtJGtXPjk3cWwgzul2htt8J96u9XKx
9XaMBkttzoTOrHg9QzSo/kOEqi3yuYQ85hX8RYNryhbYUQuQmOoBOQfY9e8eyuxa
55xEQ6/vEwHI6QtKRByoC8TJLadsN9mtmjMKJcTQNVH9m4iSFGA+wYqhkZynTYKL
7A4DEP3Ezu2StXhlKu9bMw2RxtDWK1Y2DycI5/dch43nziZ8IQLlyU/KTXP4Fb9x
VvPCVSOyuWKtYzTHsp9flmzqSwNOfM0Ca92RNdDUpDJ7oq/blAvAQYZO9HE8FTZ4
dvi04/q/mKiw0tyTkU2rIhiC1nT6nrc9tX3vreIERsZH99ZHAI2jxz6tn6jpYMrz
RaoS1FhFb6HrzwNYIeejTnjAJ44w5HJ3ImYDlsRlmkD9yGuslwU6Iw1tel3QGDnr
swojJcjHLN/FFtOoGV5m9Ed21ZICii+L+Nd2iC4B9dWh2HHi/3xaW4hTEKqL7SV/
320Ipxua6wpw2nOwfcF2FnqQ2a2H8oQZ/ydggvXJV54=
`protect END_PROTECTED
