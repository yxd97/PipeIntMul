`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
URSiY7mN4SbUSVCwv5xT3TGiPIZvRFskt3oFEkExleKt1DM8m6Lc5pQEDjk/rzBA
YGyY8j6P3r7ER/zao+VV2AnbvNZAeDNTs9PIyagFGbksoWtkdM+gfATdqp7HaH/H
6o+neyZhYzXQ7cxF177ji5U1MzvnAaOzK/a/vjjZLwZP82le2/kJW1nGqXTk0R8+
VWvLTXxC4SpindzPLM3BmON3I/goCWYTZKInFBKTOsoeMX7kjrizhNbvurY+sA8A
YhC8qiJff8UWsDzoHUnkn8USmWs8DsGDyb5CHpeGFGCl734r7A2g2++3Mp7Fzg0M
jVEfTPdRikwHXkpr+OrHI21nWzFgdB5FotS4U2Taga17iqoq12rbj2AuJewJkYo0
VUOGpoXESyNA+tn9qHK7niSKHmEQJGGJDoicfUNhtMJgOXq48FNtOseW+d2kKiFg
uBEQ7QOQCTUNMAkjrBh8qL2jzGBcRrXuQ2gFymhvgIqw47jGCafwuXfHX6HW3cWf
L2Qnruba4onQn3bi1Kbp5QEindUpvKtV6yWR/A5+iq5MEW1nq+j4/q53hxTE4TiC
GVK53JmXgNBTiDRqmzEF0vjtwozdPdNBgLltflILuxjqkupIRsg1x94n+1QbQabV
hpuvv25ZaHanPN2lAuQxerUwxXeNxrEMnc3WNW6nkpt5NHyTuHFmbIQ/v2We0dTr
NGAKPBo+vgeS/FBjCfhzhEBRSOfbpo637Iyujqmr8H3vVL4zn0Dp4GXdwqnEMrlM
AB7Yoej+1cHXEKQMZTZn1o/aFdRoo6mRNLSxsEW1h7svBBTIFEc2qV8NnQfP3dJQ
/3alw6nuMvTbFWsBF/9vrlEJyZ4I9I1NWuWJgZ+dNYFZfDeyzNSOsXTtfrP+Dvq2
EV2/yVt5h1kz/M1FxlNBT+TsZmZQnTbd7k8fNMYbd5J1+pHS630xskDzjvcNQeM1
FyCLBLjB9s0hpLIk5F9txhtKBt1nGIuTQTX664qP3t14urjT4o4F0u68+kt7HAFX
cZwiX8whaONkqHYVrDcRjGd/CiEi8D8B7DCbTEmkmfi0EDhFShvlJHRAf8y8Lo5Y
XNrkBpLAki6WgGD4xxcS80tW4ZHLK0yXr8/V1nnUtra1l4B4K2XkXLP+VLRlcBsV
zN1oqGlKY0HLyH45i2GSwYWXhQlibWyViCV5rS2shgp3DTPu0UnEwF4OaP4Wkykw
j2U/1ECs0tUm0gieWkmAcuvSj2t9ccJL/gCwPO6002OEAERqqzUn6G6xtdlGbNNj
h4akn3AzNkKWfgmd6HvREwvlHVag+S6CAxtcY0HlMK8/4dNFm3r3UuQcfe6llD2Y
AUYkWes/+j6iWZPsBjA6qUkhYRzwZ7G0wSN0UkL8gVVmTD0zD/SfDd4FP/6/SRX5
Zvba3MoInGvAA3FMFlC5j9efsJw1GiH5M/44Q0HK3wbuKqTZz2XgVVq8jIadNCHt
dm3UDGSHqAbJlNz28RO9X+b2zAB3hi4iJ6TA5Z1NF2bnwdrvjmPqlCjrN79EeauP
LeIiU5JmXomqlxBciOp6+lUUKyR4sM7WOiPJVDS9mRZyb+4hhHRiOqMujqISalYd
dKtZrviMqf2Od1vNkI7/6PwMy0nTlu2U+uLlfw0Vk6Nlx4pt/K8IsPnCcqlPBOZH
x6Aq0kGB1xxndhgcY1pQ+/nXjIvnMWs6Hg5wR4yDSd/SaWhUONB93UcUu73fdIH+
io6PfUVor7Qkt9gEVtJbTGmEQIP3CV4MIDveiO+pS7ak4yHpd9gqmzRK1oIo2Yiy
ZnfH8RVqtD4VGehq1wYrLwi8n5FNqYEPlk6w3YDYXhNe8Z9S3xNkhgVqpWFV6aNt
zEnlBZET/7wI6F5lm1hmF1PhrtkSZOTjxtiHOUfdha1ENfT0TollxaQMfqcYLhNJ
ScoT3bfDvgVbuC9ii6xIIaMeaekG8WC7HfZ0ZK9uw7vQTSXFBuJAeDx/NM/X9AKL
s/Fb4uNLlBgzi8XSPVL94Ti+7jtGxZEc98mb6SdCMkONhn+I2r1ji3rKQFJ2+4Ch
1qzUBhjDefdZYbTzB8lBe3anknnGpzyUAgPZ30YcltL1pdJi6CGcp5yyCTZGMdLc
EGZCu3K7a1qBBkm/GAnJrtGLY9PgZBJ4xsz1H+0kslbKvzAsDybT1mNSuZEDpxx5
U07ZEWn7/gcGw1TLPtw7Ql6Cs/Y+AEsvzcVxWwefMlp+pVfbufZgjrNHgv6obhu8
miyAVzWVo2JnRS77DOjo9Gvn2DuP7PFo3Bdsk0UoGXGxI0bGNJ/kD+oyBCPSoIzM
GaY17FfQfeuU0ow/14QVo/Vw6cqi4Jk11rFTKcsoeLL60L4QDoPCtgWpCQAOf/pG
NjbNXOpRQ0g78F/Uc8hrszyWlwtqWnK3/vi9NMOOqmd3wxsCD0Im5sjsEAyKdZVI
qYLC4BwGCOqL6nHcn9IeoGyme4h9hBJlLnS+u7kijhdvT3eTcTM/0ZMOmLeqk1iw
GajOTdUVOw+Ut7v9tR47q9UeEaxKVoninCbbTS3sDd3EappLf7MIStGXDcXE+TnB
jW+HKbYcaXRUg4YvqfSnz6jHpMrBatzHA9NMQKdqnFQxdwoZ/mUB5NiPFXmSLYq/
LaBqf0LZ4t5NC1yDU3pHAWNieBUrgm0GNOV9+zRnF0lcfAl3T2j4M2/f/XS0BmTa
APIerkpU0ZKcM6sOl2/JLVEHwBmwuV2e0R80zQHkKzDo6GkvvSALz6Np26Anx1yb
U1fLchVkmHD4/ACH1xVyGfpu/7YoWlCZ464vYtaVCu75h7ySORyryrUW22f6iMLA
`protect END_PROTECTED
