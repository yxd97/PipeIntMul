`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tUw0fy9tq6iokyb74kH/gldKc58Y728MUMu0tRDbPCbYGAgc4zuizgy0f/n54h0N
melUvFSUlw69k+QEQ95iwHkEUppVPGKPDncOQVNBrevGzecyv9/Nu6nnW+kKBfXE
iHqnIQ7Dzcdv5CoRPAN1JoThI7p0Fjmuw/BlA4V7u9biJPda/rgUzuxicNyEBVfP
CRxsKu4MTe6dOCni5T/tqmWTuFgT1L2I/30SfvAsc5fK+76MD+hs5S83I3mc8Wa7
7zlbPO3sSenqP73L4bHscg==
`protect END_PROTECTED
