`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bCNj59X84u4DHBA3FreppvJsHcfKCXH6R5LRQFw/GsCVKjyCan+fh0jmud2wWf/r
pCQD8h82VIPfKIAZqKghgJPH1jL+o9VSBg8767wq+2q7QU355Ae3jWgNrRAL2crE
ncpos8u3PJpKIhcvD0qefGMzUIsc6ZqCwRL0m4qV5RbkQzL0I8CbTAQ825R4nEqs
GBDvCWbTdTECo5PV/D0IDwhVRoB6woWf79jeOIlM4sLUb/wDComD0ocPPiZ8B7o+
kC95Su0gb+eYvDOBgxxW9r/tH9y+8P4T0G6p4RY8Eeretadjyfu45HKXFpPJDmqJ
JeGL+ZnG3ZOWDRk/MI1u2Q4+7IFk5aROphXcfnHT3Nr8cNeUnLb1/eLh57WGH4rz
l7q+qeMzMuFNurGr9wEK7d03XXe2GsE+oyKtRWT8t427/lpvW46V/SNjG7AdDvyN
LjfpDyYZ5ydkU3+IDiz6J8pov6HPdtJRePRY1XsSK5ZCmdUEj2hh0xO382ZXdNnX
jONtr/25RtGT+O19Dgy7gOqUhK77RZvHQjcIaxgDg+vEPaHZT/ixAAexJ++48puo
G0KoRRTBBVt38zSHcNjjLxb5Ycnwb2YHH/zuBUUhDRvRNKUCb8I86DUYyq4wZAVq
oJRL9T1XfMha7S9Z2aYIhz2/bHpHiXM11Qm7OZZp9lqKGEEP9oOhKWJ0Ow7r7htc
NaRMb2O3Y5ngPQx9axObgofCqfESVEZ4f4g8KJ6WRXvsScvvxNNLkEv+q1/vFOHb
8RbGiJdoGlMcg3m1qhqIYP8vGwUE/GsQ9QlgO8voq792qAcTJuGe0IAtKLZmhAU/
dGdAvHgPLuUHEsDBnSYe4JdctZhKSp/sXg8MlhDraI3/mqbRqObkexwS+fMFwrM4
LSXl84jJWylFXK5jefCodw8Ib68h04Y+uS5fUmsF49yXc82fd9GgD5GalvC2SE4N
`protect END_PROTECTED
