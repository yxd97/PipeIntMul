`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9G5dBBNcpu9V4JmYg9AYHJvdTWfjmMbay20Y6QLXo6FSTCVssK9ArNqjRgN42VJg
emcJaSBnkS2fxzFa2WCipzZSrrc4V1BwbUZn1g0LAF5RKs8bt/tmxRKLLOlbjLud
3uy4BrAaeiBIhX1o0i+edAX0EY2Bmlb8WdHQ2tzcfUzG/224r7Xl1oll9YQk6wuj
csFYx50oyzUvwkkMs93+zK0Py+dicRG/pk1TadvSUE+0HbnnZSFaWycIA7cYuv3K
sZ00FvOmq16/dTQymJjmjDdKPoy7nsaA7xIwvrgBHGQ0WvkKh0bxG1wY9J+ymU8f
1F70GCAGMioChk064ggQPB6wel70oIAdCtmBye7QchMiF5Lsk3llRuwyKC9Y/wXf
ehN79KA9u9+ZYUX7nll6kTteD4mxRzHbz/1FJGO5vg6UnwO+DtCyyU5HkpCLa6ef
Ys7vVZOxKq2hkd89/LJXnJCnysUFMAy+LmHg3gFtZTQHJHnAY/dUhL9ZrVHiCMJV
9Yr2Mejz6K2WwAgthE+znjK3qGEQbW5F/2xaDhhRJOxKwyve/bhqFP6oSILqcWyn
9Us5Dtjo5CaeL3ALs1mhPvLzW6rTdbcWRzxz1Dr27++pCfsuJWdddolZAbvRAjs8
M5YBzpWtkjJu3XpC7HUaqcOeMnyEVNTcrcDQNueazTsTsIJiPQN0OavSsdsBct11
kEHcUVofSWK4qyTIN3xRun4pB+4uI5qdn1Rr6qWvT3GtA+9VgM3TiP+JiN9BXdgT
rTz7aSqhXBTbEyJ/ZCRgnM+YT0Z68Jq5oBqFNI84i6BRGMrIBQEsr0Qad5aa9WA3
tBaVT6z99OumnMZvMAA6P7z1i65W+97VI5v+iyVv7MddSAfkRKpy/6FupToczkoG
xvJQZhbkjzrz9DQsLJIRrOrlw2LZ2SHh2Fc1ej6PHv3AVneyVRJe1231GU9bFCNF
`protect END_PROTECTED
