`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
37YNYIsJQUoQCmA4UuDTphqKDGGXVwbu9dfvL4jV2TWeaD+jKAsg+KtLNuM/oMOt
nCOgjxlf1NWOj/b1Mbhle+dOkTp015RLCGePUAJQFQ+9roPfr4KbseycORf8ZttU
6WJOnjIDO12PhYzgL6mk1sJM+QRy9ZKiIS59iMlSTCr6YTZ3HMGYGTm4cTlC0U2w
ZNwLnsVxzXkuDUFnnhp0MazeVhsh3zv9oSD3HlybXZX5ijXnU6bsOkym5vonv+SX
CgIBmmLFY86lQON+EihbYU9XkzrYsbxKvpcGl89T6QIi2UimNWPUWTxAoxkvumhs
H2M7UazUslEM1pvHGQzwKzt1XG/GuWukMpfcowDE8jl5uS3tvSUztv7EhNiKXSC4
pRoPHDqUAaDZ68oDUg4zXA==
`protect END_PROTECTED
