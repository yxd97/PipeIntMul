`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
chZmEKeF7eHH0V+6uY+c+6f3D8HbruvSu01HYhW+vnT5jd54+0LLSWwCQRlm3SJE
XmZKpwUJXvkGzei8RqHQc6Wz6o6qA0IGhkRQKsGiC6IGKLDitn2Fnpen+iVjNDr3
Cjdxw7Hm4BOF2AMx6c6WjSRFB1qLBLjEV6admJGVDRr98nRNh5K6iqPnx2MXQyON
JFWUZVRKNlRgk50/kkLI6ND8C+pvJJCXruS9qu7Cqo3nNVcXzrhdDj4e7Xr+5QqX
00UzGOkZVFQk8UPOTcgOhty8xIt6Ne18l8S0+VLdJPt6/qLR5xKgVA1v6lF4s9sH
y4MlIaIuLUJm29+9FiTbdXoy+oEQtLn44ee9VdUnWe4X3gPcFYnXkllkOv+xeXYw
jo6f2kZtXhX4QkNGrfaMxlTDJ6lJ46ZKeTILTz+WMUYKTNNXKCL6wWCmIUwuhoH2
qieY6VZWRhdBFAYONDBnzZr7mqhI+YWlntyeE7fKRS6H7lMYeB1yQg7PjofOFKCi
tz6RppnGR7RxzU6paYX03dlYLSIB09MFx5PfUmbeLKwjM7geOpmknSiNsL2vL8+H
EgmptN8rtvAy6QhFNZHVUbmBAlvS4BVRfAVRjQ+ivsf6B/GzIYKigAQ/OATVon5d
Yw55uXeWcdn1rKuaLVsq2nBOCGFyvjfedjrr5vG4ut9mvAU0TvJ5zMRikKHs8qL/
Of3+9fV/6/EqzQ8DmquEEURqfffS+9xKBUUgOY89JlM1eK4MTQ2CBKl/Zc8/pUAZ
RHMAB6mvATRrCaxRGjVSn+nuUkmhwIqbtYqcmRpEMIjfJDoKG07seMb5hWmEb2nu
9JuUpzuZQTCXt5u1n7GLGubuiNBJ5e830P41jWnyN/KaDMmrpYo5DXoi/PZuX0yj
4SmiWtvn/ETmbcobUm8M4KUtd26FtRwhrVpfqxSzYHkY2hFrfdTqhaPIjyoIwTHC
iPoaBh8/JTunXxt7Gzlz5eqSEsIloRmuEEUJoyzAqdi7NV/+gaJjcs2KFRnQijxl
LUVvnDRJbkmqOVdKWmuwQMQ9bdoZFB/GexQ8d+w1jgn83kUIgYHl6DtjhpP8dXN3
dkNjija7M3zpLfDQo/5TVJCqa/kMW7sk/hQFt9nh3u12iqDQESNHORXsy8apGQFE
2ygpHekTcm6w19cTVr7SqA==
`protect END_PROTECTED
