`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
unfSs8MVqQUPWbO1nMuE9lbs/GSX3IaodgdDRzc3WdUfe7dFQ/PQGNFa6Jj4vsw7
7oiYSq6NmJHZJHJBaqRfBnDtwbV8jBNWULKCIflWstiqCbu2wpev+qV/7/LMhj3V
ThjMxfKGL/dqwLzwlvHzoUYuXLA9VU9SukbnpBPiRcU/AxpazXBqUD0X/DSIdMI/
uhnrQCoPJ9uPnlKl87qYtOfaDDqt+9IwMo/8PP+hQXprS6A1i6oyPs+byX4rxgtv
sgnWlMGcD1UsIcSBFI2//Yv2ykDAcsyjyMN+QMsdNDXGAu6AKGL0R2QUsC4y2n5+
y1nsqL2yy/RPwUw5ksEkBiYoklGmxTAm8GUZzxLniV/uJWnth4zaOAYOFFo2/noc
u8zWfhHgSDaoiap6K3sivhbWpH2q1xEkH6Ik55GEBBBJsnxwOZKWkRoqx/5V9DDu
kUF3kG6btzPt3S6N2Wdm4NutnpfpoNBLRseyRhjg4VUlcy75K+rrqrvdTdv0iVo4
UY2vOLlXWJRfgT3yusEiPljyDi7IfDL1m9fUYC0To50=
`protect END_PROTECTED
