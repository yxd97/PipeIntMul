`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
espOLOVYieP9kuoGUSfdkLXdZfByaJrWXXscEkMYgqCuiXz5pT/nSXFJYkZh2VNd
w6EHK3rk5+iluwyb7/tc4HXABcG2QzW69u5moRw6/6VmO8+GNwgWASphziMvPQJM
x2lbHW3DPrBEjBX3Fl/09CDHXBtoPALSz4YFBSW9DSLhLUEay6Z5a48kQaq9f5v7
xsgaHCjrIj2CBXOKa/PjBxoFEwjx+fdEXUDMUH3Tc2XZ4CPtfVbaNwpl9MbnZm/5
LRW9ekR4yF1D0SCEB0/ZbCaAVkZYgCpmHEeMxbtXUIAEjSbhrz7A5iKjSDrIWluE
dO4Y6yE/c1m6ozyhuWWTSujv1iKZiO4w8idM+oMcK2IX2prXQHuDK6zDHsTrWd0K
7kxhFp2hY8bhKDOmOJE3GvIDQlLW86K9U9+8Wa6FXSRG5c1kf/3/oY5MbPcAzLx6
TjLnKwjb93vlSCDhn61kl8khJIytDkWZnGX56EIhEjTW5aQ4eDJmSddDY+fYk5T9
IslNWkkPMWrd2C+Hkp3vX2Tw2RQ8+O9eY3cUCT6hgwtAKVbys7VITY3IOif4+dJh
etFuKfoXim8nM4r0mW70joWPpRvfLMiNHt2vCXcV65r0aLjmBAD+b6cEX1Yq5D82
5KUTsYNtlkWGywdyoceOLw==
`protect END_PROTECTED
