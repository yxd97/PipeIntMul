`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
maQbK7u2A2R93TcXTRXGB/ABRPpmfGMnW/wOBPSIX8b+TOAeELcmj70FlFxRNtyQ
pE2vPTCj/eYCGyCASkEbf76BQgpc3Zt8zOPZI2g+V0QeoQa05fI8tuLM6I8ZtTfE
7Jc+4CHGvqxj/n/sSpZ9SUsPD4wqCvMRbcd8bOxG/5F00tqF8lmzMxaERN01nk6i
vUwcjdZ5cT/C253pDW6UIKYeBrXEvYcPC1nCCapTyB8uC+HcOdcZreOKXJ3xJ/gA
bugJPnJlAhSi2C9h4XCQ768QsN766CNbymoUXxtyXZ7/8S6pGrhfpz6/nnLDnBNU
4O8gBtx0XRW9Lww+pE576SerPizeJL0crt+BK8WfubZvaONIGNiJy2pWWI4DjB3J
jwwRiGN8KZkXuQSiDjMzbI98zRsaP2DJgxO67nOeqfPpqj+OVIYRYTLKJ/goXeBn
1X+zRP588xeGdKCZ05hLUUIso8PshzIPK3DrH7LRnMS4nk4KVKDJY6Ls82dtGpF3
vtrmWNreeTrPaG77Kp95JFOu1GQ9+1lixBt98cGsB8yXKJrJNKaZTIbR25PB5EBS
NCG0CNbf8Gp9nrPt3CTJbXWp4z9Bp9oJKVWRvKCDXICr8uxA0CPCU813FF3dt0uL
aW2wTjW2bIKpdyalKR2sumwXiFy+gLHZmJQxuiCreiwVzPwKiETUoooaFufScKLL
/ujF/5yNSGdi0Gaz4P6WmkI6PhvmuVk84oFYrQjddMd4W9PiV5kJSboizj6mdGrw
1XcjN8pJAwYbdKkS698hg63uvCoDgd80ClQBfmziAMcMZ3HRwiwkLcYGqk3dZLF7
sUB3aOrbew4e99CDsT3lk6trSw5MyiKfQseV0Q9GOhoHiIGoE1hMn/+o4N57Vz3b
aDAm1QcmpubKHZVkSR3rTWnNR0LYI3tvdOgPPXeX1qllMNqYM8G+v3x2kzkX/Tic
1fT4uuxLFJzpRTB2WFTE6q3neOahev1Z995gJbmu5r0mxLD+kzJIl7lYmuc/2W70
`protect END_PROTECTED
