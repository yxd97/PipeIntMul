`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wjNLrM2f4hbmzAKXauNXWryufbvDPGAphuvOcTZgfOsoWWU8rNUmSlW7jccZyB6r
4pXcHRIHeyVC5tSpZCByoEN13zSYxte6Tsc6ZT3CIsy3CGF/AnTwADfqOiFsH6xW
6ftMlG1DZLhsAg3l9iRqWZBC/JddD6X4Pg5Wv/ChjtGbwjM6KnZebrpGJnjKKN79
l071eo6orhtzOedr1HxWwXMpTNEQug2G7uVkymuuDcDDRHIgM5Tm78KyCx5QWqYy
uz4tAfWhIsrN2BOn26y9PvdMQtqRLpwAp1npCrNO7uYB8lwCEP0fteRtG25d7uVN
bxR6N4HuxkV2UWDsCYiqHRKxhVN8BJzB2Z2sIx62SQb9Z8z7Cuv6B/NoYqolvfk8
V+0Pd73sd7hdVNYUMieXqdd2xahLA7Z8arGKeQJiuC3sHRsbZbVXUwp8X1XRr41h
TIwcZAjfNr6DhVCM+0cv4MuYm/9p10VOXsh236E9v6E+ZDpDxbxbbVoRywC5oSJ+
ia2jisksRIcy04HjX58RtQNCDuXFyFJWiOW0cnBC9/ejTBhhx+/ELqeBgx1ksXWP
cfuegrev0VuPKsLRbMZ5C7IC++9wtZQE2jfp9I8yAe25piQsOUISd4Yu1SXNd6xm
csEGTPCBEovYWlDxhb+9Hiuf4/zga2EDMIbNu7tXkavYzh1hqs9W7Jj00Q+kpuAF
cLbPZ3Bu0VYdUaOsAN15sj6SQRSBsaygkCXPef29KbIpxWur8/zQ/ICKfAJwTsQ9
JxAH4z+/KL7BscMd69TMcK95RXWGpsoigrknEcK1wXKT4RkG26i63DZVMYqui7IP
Cncn/U5w3+HAto71INeilImn42tfndIReEeFRjFTk87CdR66lXXyrBYyWJVFIcIn
O8s/F22cQBUX8dgXOsDZcfwmGGJQw5MJoyNTwNw/isklRbqABvxi+A1y7KSmoUq9
avbT9yCy2G0np4OWFan4q4xc2/kE35MN2VSFuw9PTjI=
`protect END_PROTECTED
