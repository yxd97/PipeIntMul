`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EV9DYGWbDDWFx5ckNS9cpcQvO2rQYJSZLj/FTmhM/M5ckL6HPTXqb0c1tj7YRaJS
/UqI2hCo0TaqZmfQASizF+QTgjU+BOdETmiTBEzMZclY+ayaAmRXMqI3aJ4I8RHW
8aq7nPnBCwfiNMsoRU/ewPnkj+5MuyltyvFTWyceExUB/GDk6CGxxd0myWn2wZpA
3g96mW++1CqV0p5i2JdS23gK9Q0mnwBiTk/MpLtNGMbz7bWTV3ueUP5Pt1ShQHjk
SoKdG8jjSkw+LCA4bCUuZvpIITiRLjVmhf4WCnrFt4IyDk3BmFC0e6EzFHylsF3s
HC4+Qq5mOi4NBtAD+K2p28AzXuNkZv+xzPmYZL9PY+ZX8FJK3qXoYjqecOa30S88
LqHQEVcPHks2nk/g3NHgvvSj64XcdtmDFsbCxseyBX1BV/+7hq4dTy0tPjAHRX3A
nzkjDRIrQigMEltDszArrclcRlEjp5e0tB/s8917iH8q760v9EIo+nM2Hxe2C5A0
xYtg3U4Gk52Fv/phwEVmEvl/0wsp53BKbtho3R981I4FZVL9Vq626BC0oMHmohKm
Bee3L2jmnQeqVknI4fYgfLuaQXCAiAiELkrHCAwX7DFeTv4Vyn09JCCJuNy/XGmj
6ZPgWhM54poOfSPSiM5cI1IcmHRKS2z86riYbIvggiiGOYxUUotqUIXibaUkd1OG
f6FJzZt6m+R0oLMwwXLAMo19E3wC76vqDhyCFDykmIRipaSH6jHxsTvk6gUZ4Vmg
pshYmj+cmLr1RrpzdHXo5CM/kOXaiRBE4Yk2IqIiiCif5qKK8h3L2lnpE26XX2+q
ydxD3H1Vs39R+g4iU40JgwUppUDeC4dbZaIWufYQHXFteh+bi1/+dccHuSXPloZ5
eMQs2deF4hj2GhVarTRbsHNSjQC5YQ5f7wSl1+vjGQBdxrLaUbT/Fm4dPqwqXTwU
70FzQrxZEHkgkwVH9EWGbZ5vHH2C0IoyLfVHNu96dvW8brPGHmvpzAzUaQ09qoQJ
GfEepT0v7ZCGQ5FsXk9MdAl322P54gMk4ecgWrR/EPAUclg+mj/GiVByNxnqmxtI
X5/N31+O7TbJ4Mr3dbkWUYqjX5c8LQIYCuBZshuX4rL6XbKN68IQ4rFb66RjxCk/
FirSHkrvqIczou3MLRYvcvGNyp4uxCUApjKKqtIVXbhKVj68K6e+Ac59U8TivxtK
t4qpzWKbGRfFCKuY6SU3NNNMclpdRGB7T0B9P25y4TkUoqG0n0vtOf3jG7Wdu5Gt
0hBrerXWAJRjPzqBdIBiyHro2GFZuKtUicR0oRY8s5OFGvCByAwIQc7tIw5hDTJo
rE6cNyOqwlqKFxYXU7WuLEdm3CLVFttbrAT9+9c6d/DVYiGl6DFJGmeuTa7OKBd7
08so1FdAh7rmCBhTG/+LVnEJdYUcWZskvosw7n6CNv1kTj93M/f2paIzb5+45WpU
lIhmx5b+1IK2kkhn4O/jZJ11bb+rgxW8F5Iplk0JtwGiV4eXffsUVyDuZkP8GzX/
LzOXrkpTm4m7tAEhI++6FDWmqUD3zHyxAX78EzQdSAo=
`protect END_PROTECTED
