`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9kyLWOfkXIsmEbMdhrkzebROWkaRcijZsaW3FkM1FJXv5OvN6yiBs774x9yBGUgg
yVAriQJ+Myfey9sxwr0TVdfbnGN2IBKZwGkAxtjd2iwMoESr+vHL2tuyGwn+tPwf
DK3lYP+fHgKTwJIkOABCm5Rhzgzu1VHVz3C9NXeRzX/AkhPJ/m8pgwUZrBeHAJ4H
JvCHKH/nqXA3cGAE/mfm/3GTU/AEkBMZc4UfaR1AIlqo9pBtDs5JrXasDN8VmTRp
nTmFG/TTtMrxbFa+pqGDBeq/hKe2LkJ88BnbMKJUJ7nZV6XpnOl5hThKqV9vcYWG
rb3gaFM6zzZA0QogYq0ZGLJcncHQuZShVpYfpteT+l3wEBgvG8BCaLHg8420q2u+
JdUwqyeLEQbzX8/4bFcpgAYL8R99CRycOxzn2M4ZooCUmsXyiK4a608QYVPshhGP
5pb8/Q0RVmP52RzBAgBwaVAWfSiKCdRoCY05ioitcChsiaPHd+F7DO8qJraxLrxM
wo1auNLC9pkAZSh2b9k8lyE+mRddn66IwBiUYqrg5maKAn6hZw03Oil2Iborm0V1
Jv8CzaC/8NXViIaS2kNjGMwgDhvnJlYlBpAD6IadM+U=
`protect END_PROTECTED
