`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VJfdLwNaYNbYVCiT5BdcIGs4eYdEhZ/8Jq14sMqG3CEbM5+tPd3W1P6phM70oy71
JkCgLBRuMsTpBu8siB2vFffapkjKY8jDQR/SqLVUCFFB7cm6MU5e9I8S7tPCevJr
IQ6AF9Fx07KgFVFk9PABIkJtZMrqWo4w4zDf/Tva7mURmHb87ltGagNjOMX9mA02
X814SWqczVJMlUJ9gT6BJOb6OeZFfI4Li2zvuW99WHysFPvUm+QS8l9htGeTocgN
s0g6egb+Ac8FMdaP1T8KveZMt+/dvXUWuzGtSzCfRDU=
`protect END_PROTECTED
