`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/IPDGelOPc4Nwqy0x020k2XqSbKfmOahGAZGSLZEmWF4ri+nc2LmV+lRt3oYHs0G
FDSjSjqkIvlvsB2Jgsh9NzgJx96qBHD6HzkE4A4Ah+OFFcUXD3Hu/W82scBcYLcQ
/NPKiYw/luFDekhtYkLgSdCVwVLHrCYsvTbqrT3lEBB2Hb7Deim0ZlwF8YgrPr78
1dliBZXAit5b0GJA/U2WQR3tl3YxjNApKAB4z1Fj3un34HiDu9vq+H2dOGdmxpFF
U/fin3QRSzQbQZUFQ0PwND8p1170f1iO1SgKftQyXvQreoi9HWDG/DS4Nynu9gKT
9lcPu71ulaSB9e+vq3J/Ln1aUmXqZNiT1h9fIt8d+zSoIaHN+atOj7O4Z/AHmOgX
OBV67DlOezGxybSHTRwwTQJnxltOyuqDuB6LMRfepLzAX1JLHAmsvQBiOKCRiDlS
sBfxyauTxV08VKsSh+XUfQUIH6fWUJ+kyZ62PXkzNUq7emeB8oSFWXbDwvxlH5yt
`protect END_PROTECTED
