`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LynLU+Eqa3I5DZrNs+phcdiaKg4mYhAcWtW7MLe/BKSOd399bPGHGGuCsAlO1IiA
mrE/vRyC3SdjOMukaeNijQR4KwjmMsp28EWKpHev8TzxYk3FXMpBmB4sgewbVDZw
Bk1o83NO/vB4kVJHK3V5IUcS3994OGnHfGutN6vVRXajz9VQyM1+QSZr6g+IJ1Zy
hr74i5ANtqry700HSrsp8BOw0FgNqho1gW1xLmp0cDXG/+viLHT5hqyQmBwCo0Aj
q35wZJ28rr2t+OVSIiGbKRDwdg0m9eAulswEbTvTRlx/gQ8MGru+v3mg+dUCBPoR
AH84+F4rUfqJfN4zbkLOKV6xJ3zBi2aIPdqCu/f44ufy6Yv9BoZIWFidXqVVdk77
EZyQtQr4AXrxgqF7SSbtzHj2wYGm+7BKTyrWrfW17TyLXQW0vIDMotwVaUFEfhIA
VGjB5QYCG+6Ey9ORB/a3DXCWZTKrribyq0kT7WRzRIDyH6dvwDjPZcmhAa+UckwK
KQS6hthPJoxpqKQMpusHoQ==
`protect END_PROTECTED
