`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HdF7LfZ0jJuDIacwQGxs3t0TAB6dkIshtlf8FlrH3k6wlwEHGVle5X6yQrFmqsDg
TBohemSE6FStm5IN6IJtHb3BjIN/W6LaLVVZTK9RKaxy09qZ5/I3QjrAh0jiCkqa
kSpfyh7FD2fuOaTKMJvcaA0zwq1O9cbWCWFqVN2qTCpCI3QRdd2ISzFO65vMq++U
nPBfyj57jzz27B2GwWYE5VO4XyAA8zivUnFh6nBx8fCGlwPlkL041usBb9zTEctd
g/WiVk3kJX0EXfvXYZ/uwkNihcH4T7l2c27RuIhM5uA=
`protect END_PROTECTED
