`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qHjBoMg/rNmCKVWtbSp1OfSdhyBGGsKvvFdfmfTRqUVhvmcXYjwGXBQZkaXvoo/
XrW+SBIcmn2jXks6pmPkK+R7WaYHir5Hr3nbnXm4/bamZR5zTP7HV4JDYfh1S0tr
AtnZg2AGT22wMV0w8ya+yGBrDaQ7zYTWdJNz55awxmYe9EcayCLHgoWQsU1OiT2W
q8hVgsKUBRnvtcyc1tc6qZrIVzN+QoZOCSY9HDXdyn5zT4l2E4+XaUIMDsol5Okl
aiFDikDQepkGG077qLDf4hZodN0dxZ/bnYa1BMx3RTPk4ZiKQ7chlfagdlSxGuF8
tWC9jog4eRUYEu/Q3oMhHVvqGzdkNiv1u8r9qqh/XiQQoD3HG54jSYFuunoJXof1
m0FNc70gMf+xpITgt0wKoyuwHpruuCz249MUMS0DOyuZ6IKIQTHI4Vb+2ifajdZe
BH657gzIZ1/rLgua/XEkydFWQPGnVz96Y6uvYun+M0/6Z9rBmSa58AK13Xpm5Nnt
zwjgYf4L6F32apdec4lRj/WmfEk5EUKujvDmvSPLzI9aB3NGPzKsoJdPOuf4hMHe
/765ZvcpMpTfNaqNYu6iWA==
`protect END_PROTECTED
