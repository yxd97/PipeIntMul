`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lAo6k5XO0O/z6rshLFTpuxI49nsJW7RT1EZ8ULov8yHoASinSX5L5b155cTg7Ugl
drfvIP1/rK4oiSSyRMIOsEmWe04ITFmF3W2zPxJSCn2hnfT6XVkcAxDqrO+RW1br
VGwaD9lrVynR+kaWtIM8kj8Pdvj3+wtQ6gsy27vmzyN7hhueJlYomB+/RA6dqtCG
rTSJWbX3XNX8nzs1FXzv661IfSdPHuva+9TZ0b4c0Ln3dlsjwljfyBQ/TQgPCKmq
w7AHwlXNj3EsEsMZ+5OvPuAuXZtv4S7Y1r+TuKrPzPbUGH0indEObUbWcM8k4jt3
mCOPoa9anBF4BVNwHFOTUg==
`protect END_PROTECTED
