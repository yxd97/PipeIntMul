`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/hIK/tsiNLEKqZyPhb7cTXyVjzovWHZLdWjPcsY3UL/koCR3LNfGZlTKA3pLodbJ
XO7fGswlQWClmeeRDGgcDMnxmIQ6u72v8rxdTDbkEhqHZdos0jxi/2jYn4VZ1JQK
j1atX+hcIQAm2HWYgyUvtrjmKPxIwFUIpDC0qqnw74ie0B0LLrw4w/T1/kg1DL22
0iuj7R/tuT9A6nX0Zn7FCuhB+cZEOZhM4KmWfzrdu+xnEMlAtqFBlTddLYAIr/of
gt5BzCVn+tYe5mRL61Yyd2upbzz7bJw1XIHhvA66ypRNaIOp44HVmOT8OxnsFaCI
/KWNArMXqTsZXzSckf9Ip5+91k4Bx1+yenNJyvWl9DxvQjXEy6cRuj06y58fNwr6
U5lMdJsKI/Lur734UM4ZrKGZRo0cIZpqh2raI/moVEVg/33sDjx0YGorldPSttIF
hu9AdlI2Mv/nSfZOLpbAx3d/uZbldLMrMSi7cYltSi64BgLLkE4yccFXE/mHmSpA
zCyMDqBeMqO+KkVil5LvWkivvdjMRgIbviFqF8Rpe6PDKUvgSHd3teyN0p+dzTco
icN2iTI2nx1DsKGwn7DioeTu2FBsv+wtS1hd/YIc9yUOzDtd3LKRkeIeXR+GpsKd
EXcEuguFy41SFVf72PG4bA==
`protect END_PROTECTED
