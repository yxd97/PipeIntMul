`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8anfo4WFagmpZEX8TaoKd+UcB1htSbK8epU5Aro8P8M1+l3cxhy2AZsax4XqD1hW
kLN6b/VwwfWIHBwMPjm2Wwj7VL2Hev/oeGSi1N28dH1hYaacMm0gX//hX30tpmJI
38J1kRnurTILSy82Re8WYP7Et1KUr17wtJolkjgK83YemN/ZafeobrJ2tcRO6JMQ
EYrF+nTl3h6IQ7nmMSoP9UJcnFgcLDXKimspRbMoRRYFFKF7yilZ1AotcFW1TJ2j
wAb8Wg498zEesB0j/O4mCXRLiCJUcFLcR/yHMGynacdysFRES9+MLq6jOJOqURxi
XEiAEtpKmWWcqICZ1Ci1trwV94bXA68BCTPJLnIh/eyJHC1VpPmyzc1lmJQfCY/b
IAr/iSn7LSBZeb7ct2A8m87gbqSCfyHYzC81aDheRwdCX7g03pblxdb9Wq8nnEqT
7rDaC+VbNoW5xNgadeo/GDa3ZB+c2LTJ/hi39EBKzSEXEVbk2x/K7wYEKswK2bK2
33jeeiNweaJhVN9yz+YjsGT5rKbznWgMtTol78e/Bt4/wD5z+jIK8bZfgH0/+de8
Gk/n3aX25VoGV7y8ffnI+SV7qpFPdB0iFn9u2BXQuPE=
`protect END_PROTECTED
