`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MpwOZXGadiawVsRdj0nhRKz19ocdk4rT1sPApx/RxPLbJ1lVlme2GqgS5gF/5HuP
ueVFp86ZlTDvU0egjNkPDeTR2GLTfxX3hBq+ssMRMz3yu2y56Te/+t40rLsUES+7
hHqtGXmYCHsZPBAeMAEh+eujR7W/FBg+ZXN4190QDRjtmuh4x4epdpxRP2Ib+HnE
+BPWE1ay0eBKFiQvlb3HpZxRTzBOHBUiKzq5hKbkXBIKb7ruj5ldKVogm/64YTh8
oe2d9GjwYLXLBuUr2V2gi+52HCIW0WOyEsy4CKmFkYp4qNh4CkqHRk68pqpAC+5I
5Q2bNliCr+/mJcQKa8FV2Xen2IzUA25V1kJcetm6ONY7g0aPc+8cEWTZVKtopSBT
61PFjV5ms+GWn+r1+NLxzyjN/NBOaWWPgjcJz0xLUAd1moEqOzv6zAN+EuZW8EZ0
uLPjkO1tGJXih/XJNmatgpYumIZCKSWnr431jXihsHiFmIY74yiINpayLO34bmhT
XolLctYZvNmz3lCO0LFdFlcVdqVzZqcg0nJ366QbVZ0egX8Otddw/HFqDuww3ivy
FTt/T4Yr93GkKt1/nclDt+iaX3SpDI/DXgAgKXqaQLyPUN+2NWrmPT74Gbjgym7l
iySit8p2O9u/rJeYOCGdvW0lWiUSGjOwUg5pCzvB0Af1aIQzuiSgjEn+BahaAG8b
HPuprh4+tHyvWkews58NiA==
`protect END_PROTECTED
