`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CfcE0ayfKrZvx9IbM/JlXIYMEa3libsPt3usQoQXw2CLNhEhOufo0d9YAWrErnn3
+q644z+xKiWgqVm6AHjbtSCd9srd0BxfrQsNUXNhXu0NJNobANUjIHOfdcsDNQHL
gLrTkKdJKJREj3d/jmaXPdvldaeECWVs5k+4LqOxcfhNz7IA6lCrpkCrzAFezb5t
WsloJa/l05k1ibMvpcdoMYpkVCv5nqyQ7IeLke59E8so6NRVUlT5akHsds6W5hsa
QeVAz7cebOPubjEgyLeQt9tWKiOFZ8Cf19iOo19bCyigoQXSEDJvH6szH2Bu9zD9
h7gg1a//5r9b5qhqSFDuQJK3TGl9bQfyJPFDCzkoOgKH3ECdXCegTRO1Qj67tP5K
Og6pkBPPYQqWrmTwLKT380prhDou6FmrQeOzcty2wKFVQxmKjVDOphVhCux+Mfki
RsLq69VrupDNw153n2+Y/H99JmUYfnrbI4dhirzgx4zr2A8ptoPiBIfLQsqFlte4
99XwzoaF0LEow0Cc+JoRtcSsjAj5ZCEWn9NWOO4gkehjudP/LpFTicXoufUIKyFc
UIvHkr2k/4eMR2UZo2J8rD7kiZz6pOuqJThwd7Ib70s=
`protect END_PROTECTED
