`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k8FX86c6BTMivnIRtDW6hQnJCzcTwCGVmZUOFIcJB6+5ULOaGK3QvUo0jgShU81l
p1UEymABOvXu1Vir2Z84a6mYpJv6pqClC82lqHPQNl8BUX0Ccy/Nq611lJ7o8Rqs
Rb50nWCLtlXVFuK7zdDsUmTZ+5oK+t1dqW4Q1BMouMD0d4uGcSYCdFZi2vBCo+/O
Hne3mxDVBVf5u4/KKVGHvul8CkHbPCfjA+4pwFeytoW2AoRav7lSyTiIc36EAWXc
++htSwhCErX7jlgiQPwXmbrj0cl9O87JG+T4uhABnWrj/NmZVZthljpaUvoaDaF6
E6KYs1262KkCDQXggS9bOXJCiaG8r+pAM2FCzurapwb12ett3MymZSHj/r9FGSAX
oUZzB6ga64FpRJDR6AdkWGJ8DxuSmvQsEDA5WW+xYIvzV4plBqL5zFne2l4Er4sj
sM39WFNn1b6WRN+u9fB4ODAsTdrPKxVM0/bZ1DCPct9i1OnUpM4UfNXEALvMG5aD
F+6wH3s672lvbtWWWtD9hCq8dhHK5U8oMgrCOnaw00Poh9L61CzkevbsiMVPipN5
DJk7VwDujeJT8xt+DRe90dG4FXoO5+YhIYXj6DcSy0E=
`protect END_PROTECTED
