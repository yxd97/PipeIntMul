`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Yi7jc9Qu7T5SP8EjZ2PWvCUps+kV2onQwUEo+f8XAliKj/1k4xrVd652kIr+yHxW
LbLMmmmBklXhTI6w3uB12C0HTPJSJSf97hLqgoEELEwf70Z7hlYJJXQ6PYW/Rjy2
hOOEfExeb6ktqKKf7C4Wu07UfdTATq6CeWlVq1GDyY2xoNpv/xnSwaH/uHbNmGFb
gP/s1nNroXSjJFNxAzFAH02Tfs8l6qrRTGGgisfGIjVhCxlyK+7CLHT4wnRTgffK
78UQkQmcE9t5gYbGP7DTGQ==
`protect END_PROTECTED
