`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jbZ4/NCWHWhi3NqRoUzpH5j0Dvl8xsXNKOnqRrYplhAbcnakXU7jAmmblK6EKD/C
TakOTjlCjdYOm6411gHnwT+ib9p9CCTNlrWwei1i8A1oyWbH7rpdz1x8GD8FAml2
wRKCoefNGnnCb/fP5j5WhxXDXMFyC1cLCEcMuGa9CbLomFofa1BLgN6msLji2K2q
Mdp+kpZqBkDv1TZZm9pJZtuuJaHtamMLCoQBJb69Dd3D/Zpt3oEkCh02uxY/qVr0
RTlpNi4Y0qaFypHjCqkkCIois5wPR4rPLEoZUupgirJ0uJ/IYBZ+EIgn4hX+O5aV
RdF++P03yPHIavX3kZ0lCFBoPuF3KpChx09H5iqFwlo1FHo1fJvCvDeuXIODaUJJ
cQtYrAqLlNOAwYvoUSac6vK76tsHdJD6lP6KeDFGsDu0h8f53ff5cmf7Xk9pWQi3
LM7HsGpj3GbtMoTm5IAS0UXqRsudnFf2Rv0Z0KTuPSbZUiJuQQ+X5xI64AvAYo1z
g3d74FHj09cs3ZABkdU3P+oVPPUOn4IaYvMrSbm8WqvERAxmgfpoXcgCyKeHxSGF
VmDBlRuEojpLZnm0SYhkZ79myep9Vn7UbLaqD+F3YWAro6/xvsyXv3wm5TTwrFbS
rffeh9v6Mg7Jf6AO3+yM7A==
`protect END_PROTECTED
