`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
a5h4AmmQAMiuEvXtsZNWeo95/nfKdGZGBMvYFpKoLPgOe6csC0A9TDYNZQ2gLh9i
I82xAOpvTXagkWw6lzAUnQ0e5KcVHusrEZNman+/+EiQzuamlBlamlFOnxeA4iR1
wX2vHDDQOnlAXD20liJ9068M12pO/h7u7VuGnfduUdk5kSqT5jCV1hF4V4fL8OYh
KPRYReZjoZOwADZkSiYy2u/H+5iYRs9g7OOh4dYlGTV8TSLAxbSG/iQ7lSb6mIsM
xUq9lUMBXGkJPQyE3Qq1cf9NfjTjF2fj3CP9i/eyypj++m5tdE+08RXOxbS1wOI6
1Yi0wVLG78XxmsENulWCuqrzpEqJzGX2vHy+tM860dUQayroX2v9PqorFq6aurXj
BAARXQdNKXP5SKGm/HIvwM76YMKhBaJjEklMxJnTNwCYIloJqh6ci/NU5fNXR5aB
n1aetnMVdQVzQtY7hF8GeQ8dctFYR0XzKSDfzXJRatQJusSrC78p/TdeBmHB9tmL
dXv7+ofMxKeHXtyVt6VoIjTjQSBGNxIIRCFfgqKKH9K5gh2Y8GQeXgAS9xZTeLaR
3ZpsePn7EoIXchyy+y+69oPeedIroOJ/seIQjhm12lEWrD4ugx5cM2Gcj9H3E7iO
`protect END_PROTECTED
