`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nOqnJjBBmpQgmaNkYf+VMSB79hreZYou+zn1Z7slOSiU+/KXVceqp6sWL6eb8Q9G
qmN14+Meo49h3zSexILL88u4J69EOVvDbzbZoJ6Tw2Jy++RXyhW3FZiPef/T2z7a
E9RBKO3OEx5RXBYLKHNotMfIJqcnIRygoA2PPAwMAJMCj+eVw2f7xPA+oPstJaM5
OFaIm6y4UlbtBkeugiugEpzpgX69eBzi+XEbr47cKSKdJOGeY0A34dv/JH+euDzN
lOcdX1RZ5zb2XDTL41LKFgWR2PfXImK8G9Uz2lnxZf6KXIjqCVn2klqfamtIp8RA
PmcvFE1mYpRy7l/hT+cvuXYEnEv1CWEgRdT2AjWKb6+rbNmprCjpm8gJc6qQkfG3
6HtW3LWUfV2IrKiDe8B6d+YsfpE5rW6XCj2zjnaCZhw=
`protect END_PROTECTED
