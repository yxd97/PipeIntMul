`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7jhYauMhi9A9k0afed7XJMNbd6ptdye5PkroYE5ZWJ21WIeAMLbMRH//ZenEocGv
06Mie36uAnwYUmEGx0wwd4lvg1DmmXi+q9aBKH0FB47DBO8slziqLFrei2aEr+pv
NqRIp/UQbydgafCJ31zQopzZ9PASD9Hslt3DMLXeiTt35hdV0E4BvrhOwNdS/3fD
JwcuM7LkPfYBfSd9P0BAmQKezbNrXp0C1L6Er3MX2NRYwPjEFGstDBhY2Ml1PYRU
9U/gvgSR7foSvUMa5WQriv5ctGt/Hy3jzg5dzwr5msoTL11Tr/MSfbDykM99IaND
ZyXC/VQC4bH4riAAwuHFm/EbqEnaoYtLRpD2Sejt815avQpCHPBOx83ogcF5mCIS
Hs+zxzzYazup5+ZA2TBSZrnmJmce17l31SxxwFufO+bkcUCsTY2OG7jtZuRWdx+b
5CenYFrtDJ/wS2u7xtjlvPmD/dUYNYwG/9vlgEXl8ElIxqgLFgZm0gwH0GvdXysZ
rHeFU+oUTveCMesigYZ0BfgPOQsJIXcfxsU7dCpPF6ijrTCcmgoj43xGJisuORRL
gvUtXNjS/Vx/SNSfJnajh4pJZA2FS7tmp9TXmtAt8XidVW1WzfH2quy67Pb+xrO5
+JEXQ/+g0aelXJba+WhFCsUtfPCv+v4FcywdAploryCd9/5JOKh5c3LAv2aaokLK
`protect END_PROTECTED
