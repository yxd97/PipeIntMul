`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kWV4iwbNTYlB8CwzWhGBb6OETnvkKggoC549FmuKMKmVKc7KqSG2JnYqutN7t5Ef
7RLyGk9Qj2whqdzMXwt1xeFAl4Iy01MOqy6iT1PlkTqTsOGo5hyvBHcm+U7LOfAB
ZR6Gdm7wMpqZJ6FGTGPzvs9z6R8RBrQEVQVwXKZmYaHa77T1QFOe1ARRkgfbFy1J
Hlvfjoi/B8+dLKRhzczHJRxMuuakvq2sq/xdrc9YE8VbMIpISaOZbPpEnqFgvcDL
iFO7tPwnEnsVr4M+EllNWznRPZXCFfWqwtAWgdfQf4gXsO9sln622j8v/wE9clSj
UMMpI1b6xZ44fK9XAn3PXRh/hN/i0u3KVOsNQr+a1FUjLhvtSWGlzZFQIvTWRkrv
z3rHkxmYtk8uiMQsMvMPR9d6Xiu36O0JMWtdnq1u1aZ05ucH3BpFXy4Kf5u4gpt+
c5W3WvZb10AHSQCM2YOpZ8h0N7c4bVY1/aYSkZmoQ/oqfyw+ixxw+k9/ZxVAD5rW
`protect END_PROTECTED
