`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f4kkQ7SAYGib+AvcWhYUx/azGqCQ3MQ2Es6IWx3Xf/NsgYwYMI+Kgz3m3ZPSq1oE
A0iKA/5m1v+az7ZsD44/5JPPqyLSBQ1VgQfC75YH0l4X2DhIVxkV0ayBEJv2FoyX
CQ31PW2l6/0WzUepPNPrNS63abzcjSXzxC52UEDi0zVYJhCCFkmv30AePBo3/gET
lHxMhDsKztxFrQUg4+5TgPHXNET8du9Nv7D383gygh9Jogs4mouV4vSxF7hCGL9/
QXhxa8TIdRDDs6NNmtae6IeeRamBWYRIq4X5xu6URyB+yW1i9nn1ktkurhE/6j/V
Kx5dtAe/KnNY50LApkn+HCkq6zJRUln0F1jbDmRTL6ONp7cACPsvHapZKK51yMJ5
5prdQpjPi4J6VEgZVMG8kLuYS+cVwnVl8rWCyI7jnETjDyDRNX18zfB4Q0gTcIaZ
k4R/XDUX5ccgaWrO3RpzWA08Ejx72cg3uhglVw+I5Y/TasUhCLclGJtgU8oWO/4z
rtmHlHL7dFhd7BtPUF9/HK2m8HMSxJy6frVzTwECL+s5/SrYh8f3CgmaGOPQg+Cb
wTw44SvQBcwseXVKiVKHte5MLQsNQcBSsJrJe3AzdzyO9OQCzRqEMSu0lJP1pQna
Cco8a5CbJ4f1spvDsN2pk2wekreEjyZlkb7GhXha1ge9TAFKKbdWAt/somhgzWOm
PTfoIs2iS6/BIGwFDXcUCw1QhnLtvROVq4TdHamG3UEmmtxUHXqEC3P8aPkJBPqr
DcZkbkKjAzJQMMor80I2CZ1whPO7MSlXRmKrrc05jOVASZf+Lel2uYo5zuah341K
nxKHgkZwgoZ+fAA/bl4q5+YyU/7KAL16li1dLxRhcYS16W319SyzpJcLpXN1RDiS
1k0ueiDj8WqBJD6Oghd8ABHfB+sb6sm4r3vtubE+J2ffuiaHcZx1K9qCbkL5obJS
TJVV+0AmBhgL6BpTNnBDTVXRuI3NlkmKQOyqfM/hgSVpvB5Obh4v3CKtWuOrG97n
yydJsLVQSYBHDq/34XfHdXJ3/1+wZI1SgmVmNCxSUwxhZH98xqcZEwLHa6XKPOIV
UpQk8gbixHXkPHAFoufRTMVCkfqFfEnqOLwjAhPSRr1SGK8NMC7Gf+es2TYGiytG
j3Up+9xeN4AncOacuN6bOTuHF6OkZVvM6rXzDb5ZNE3u9XDHXQVFAkCtxruqaED2
DwqVSm6kl05QeElLqk+ipyBFuDKmtFna8Ee0sllvtflt+pX4jJXR1QVhtGDnCgGi
0UdPzjecUKtZCbidj+1AukXPvuNMCYkWafYwevmL9OuPixYAF9kwz/5ULdxXOpJi
hrYpeDJ7ygAJWsSs/gpt9cYE2o629APRqz2F84In1GNPtAEMabLMl6f9C/5hl8XA
d/92OrjHo6jLva+8K+fAkIis2Nq6TJGQLztcR/lXiBBagk2ZlS/bT51bcpkhg6vh
xqhByt3zhid6BOd1R67G4SURUco8U4c1un4OTlFPnLfzNrMZzBCTn2ctKiUwo9/4
LJDPeTu+2sXJ6oDzlNS7u3CRhVccIFpuB+Kymb/5JdbexZ4lUX9kpJFH8TJVDseg
dqrcU5EzxQHa802nJ1qJcik5XLDlH88E5/+Mwy2NbZbsedoka1O74ddXMd8+p0fS
bQ+JElHjoYlzq2pspejymcjK1uqHJtSWlUJAoElkjYrX3C4RG/gLpSSSxBvfc7Hv
Sy8mFW3rUNnMJG2c/UeHFS6qA7iQuhrZ68ntFdCNpjcYfwcVjos8qLSRXrc84PVE
weYt/MumX8KWcVzT/47JXX0oSgppVTZtl8YBmJ49ROGJN7gwqopWFzVe33FckbfN
qHwi2DrELklpATXvQsNSRmr1h4UjRuon00FXo86j097lb5sggrO4A0I1Uq4s2yQD
GbPAsik1t6j9ywiOSZgEIfEaDRyQkXXFnOFX5oeLvuIfUxek+F/wHURkZJ3oY0CM
ZkzZg8yAOZcSB9Tf0qu3ihp3M/E1eeZLgpZnRzM8ZXCERFMwyx5m8ppWaPdMf+k3
BCuIZ4ECwQYGKrklF16rbbJqqGORoT6ILUHI22z2TWL1DiLO6SkCryasbG/yDoRu
wbnr6KsX45tqpVIqdgzAM0If9OO6eHMnN8MlCiapK9M/uOkVBISiD/lyXWgT1Rgu
gn2KoX0OUO3E+Yoe3jTA5kATLiTNj2jUX/GD3vQ8oVpYnkwGryQ0vCzENOXkIXYC
oVVaoh5B4fAXiEuLRMGtCZauHA6swsG00xy7qpDzP2B+egp79YcO1OTFwqhwSBCS
+O+CHotCrO8YUZTF8mWNdPnmKjsV661aWoSRUDTdJy+4BmSsiL+2PFj9M5gzbgnr
f5wMeQqSu6BnWs9ktQYoFCnTz0r+IgCjTPoKvoUNmZoEaYc9mpDtkqeCLhqozNF2
yrK8zcvoUDpM66Le4e4AKiPVk0sRViIkzpDqMHwzTrevFu8tFMImiiHk9DogJrDT
uLkopzNXGL68Ls5e3Vhki8j1r1WGURfmncoFs1Xck5W3RgVaU5Qh7ygLEDk1XlRg
J98gBnxikJ7BCBQ7ROsyF9lTFzdBu5qmyy1RjITEO4Qo4Y+BzjYaLOp4gQJfVNZJ
w57O7l9E1HUSdybqwU1A3t6GU7NDrbGBLeBDJ6DsOHSKfNjghh+vWtDsRzvDHzN9
YrPpw85d7DVt3vEsIa2CMUsIBFX04eO+/YDZ6E6MCdSxclmaJHwfsr13bwxIB4QO
WwzawcqwvDrg2WiC0Hzop7rSEcGEcJUw1QeKBbcSjajw0QTQ+y/vwA01IDF4NNbm
LGhTL1iTsuSbVrtUNMAg2pOAt5NIgcKP/Uig8Xere1vmyvWVeU4bQihNFjPnO/Qq
Mycd0Z+f7XdDeL3xyH0ovheXkRIZqi67iwIuQaTg8C7DZb8+/cFXdl5w5+awPA7F
19Je9CeudzkHg4yqe7hoHzWq5j5ghR7HbAFVHtABJTnjNBiIDa0/pDBNDpHearWW
cXwHyd7xIqltDTExhgKFS/xQjhdT+VcPz+axJDtmVygEY0qO3ZbVXZli2waLjyin
swoOOd/l6ui4V+mvNitDFlEuGvdXKBc/bJXRCgdZJUylN1c8i8IebwKQjiC2lvKP
BaAMQn6Ct0xGZjso5ABeIHP3Z+7IJ9aeUq46iApR39HknOruYq2reuKVKT4ApG5i
3kCfUI/frD/8GYn2H4cElSqjFlHJAL9b9VKpAle2/BGX5noEIWVYA6g7BTPTneNk
xJ1sgOtx8iruvwuTUQW0fxbM4RfsdmC/Es0zI0ac8pwIHWo8Uvbj92GvcxtB5L0u
`protect END_PROTECTED
