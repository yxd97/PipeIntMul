`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c0Ljph9+l1miNG5IEqOjCCaJNoYNSR3/pyiZfBtgw6NGm6WzKw/UCXTJMJ8lrdd9
gf92GlIMcLt8abl5/ZYlXLy+C6z2zD9xzG7iJuT/mekICZfE+vEVmyiFstEzGHmI
dy9E4tty8kfjbaI9EGZuc9wMQ+kH29cuXN/1AOxefgSbHUr4+mpsoXFwdXMXuAYK
WYla/P1BuIJ3P/Ztnxw2afzBWSiWwuuXiSrfZZALZ+fKXEl38gQedVQHrQB+Y/wN
7r0epyIQS9MzUN2tqmKYqoerbPvViotNXsx/j2PD59RGAl5lWUWqBQ5v2QCU6Lfv
T8dk/Fa4Do3qZGaEnYUesHDULJr3GeVlUZeb7KyH8P8+G1EHFP00XAQl9cAhGgxN
/bEiQBXshv0A2P3lNz3QFLX0FNaLTxJPdVlIhn3KI8qzJzzLatbliJZFYDOHmJUl
99iXiH/xO07FcFU6uCWvthDuxkpwtJLlL4y5uqUReBhsnUwgOuJ4NIBZGOHKyLN8
3WlBnhVMQvX8Ls5nuFuimvGR4wrQNJaaRoT3ONGyh1/+Q2ZyiGLla4vVyFuW9kIT
UJFeY8XAjtZK4xIe5wkF9IqZHXdjkYZ6JMamkDLyXpneH0KnHI7Sksc8BUyQFJOU
pY/4bDMRl7xkYkGBXPxzRsIgQk3iC61ZZqX8scRMbEKBa9fIPA8IopIWnJ+kwb+w
Bp5HuYShEHGQfx/CB0yJugbntvRdBo7SKkHhVDtYdN1IFnlfZDc7+reUEjXzLaAN
7Wv2t48WaVGFHviAi+ZX8OwCVZiGL3iBJ6HjC4EXMwPiFRRgq3w1PyFLC6CM2Yu8
OHYJ0LuLJvXK3t6n2mB83SlrHN6Jio52Rzg3Eus0uVBoNo054DEnJowc90pLPEc5
6iC8uza+Bw/S1n951XweVDMsgVC4hkmoZKE3ya6+Fvjx9MwpHnvIJ42Udc9Cd7R5
XhNUNyFO/aqvltaWkAlEsG/ZtVgEv5QjpJ3+ZhbWFdy/wwMNJJczX8mgBks6CZDP
wGagb3FbusWDHPRXG4YKCdAE/d3epOZMoYVnkv4B8vUqIWhdE1h0U4ZFLNY1kNo5
XPIMUKYslGgscJC4lSJ8J7/LZu1puyWMEudA35rO+CwiXKsyGiHsne0q7dscNWaS
GzImucnFCq0YFjQXD/2PwLiwBXPgRr/UEnz7yQyY2oiYYu5mhT/xQiS9a5vDbtzY
vm0clauLMdcZMZrr9mgKGRr6S8rhgMrotA7GTNvz1tXDj4itsIte5OfYZO3e2Hz6
34346wVa4tNoiIDUbddJ3+CSl5BCk7pn7ByAi7RD520j6/1c6Klp1gfTaHw9mOaB
bIiDjztixCL/OOtoxjzd84yMfoGyDTIUweT9UQ+pHLAxibtLqlkr0yvBTekRk3hg
LDFmpuNMEkRjJtwLwLmxNfr5HXGt8hoZVD1dZoNym5KFJsSf7IXqSoBAXsKLqO8a
`protect END_PROTECTED
