`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9EGks+4o5vzBQTwDzUGDqLwKzXxmXPcHx+ff387VXlt3TsMBup6hqBn8rScoh9Vx
teqRLtOr8lz/PgvDsPv4PVercqr7czTrLDESMWhXd3u7EUg3blf1cNbLYZEhaD1h
fnnYrtD7Umd7ZKJZLg2X4LIHUzgG6UhXY1YvOd/RMdmxbZigR0xA6cfChAVPHgwi
P6dnF2dW0aAekOhhScXtXm45sfGQflcDMReEam4YsO3IF6taLgr8C8zji0ZwrnG0
bU7t7SgZBIgi8834TCcWZA==
`protect END_PROTECTED
