`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ZxJ0o4K5sGNRVmsBU4QkREH1zguExDqVfAb9TFO3kEelPuOMJP0UclEvLgAykVHW
zT89n6MfLoNk5io0lZF6A/7amVrE/y5vsobqhX+3OQW94lp3tXbckD0NChcBgSvG
MLZvEdpeyRXxSOnZD7i93n6FcCRhEJR9EPOO39R8dBASr8E5Zas3k+AWqUvEkDs2
FvF3XZpYC5dBifroKXF05oYCGSNDTgUYP+8hYIqDA0GPa3M1pLdLwOkyV1O2oxHa
+0rhjTDxAN9qhYi+Ho/wnmpZMHkLpSHSlf7JPyE+VilnQI13eoJ9uqrQnd+DB4GL
5+lRwjuCxBugQi+Hdzv7jearWvQfDASfQq2vsIAZevq04by0qUxancGGR4bR1xVt
bF8RBkL9NI0aXsxlFdysd0J18bSJQWNG7RZIl1kD/A293WlduXJE1U6jai5Qxbzg
uPYqKAzIMAU2gAlm6ZlAnJp9vcPzWkNARx7Rps7uT1LuQECqoYYkT5jyWjbFRaCx
sY45rWLvFMvtufheUA0GRq5Vedfrz2j4BuWVwmdEsZDTVtwrjS9WeA0iGmF5+Rj6
jwgiGjuy33TdnbWObPuiGi4HCQty+YR84K/119GmpNb6WpJ2HARVJePlr56FUji1
9pcqa22x2gRMev0gp0NYrHp66gHYQQ7xBM7bu/+aP+hfo3bwsIarzfRxQxL2Vkda
iYLLMRcFa6Ig48xQ+hPbPQ==
`protect END_PROTECTED
