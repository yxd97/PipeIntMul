`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D3b8BAiuw/h/5pHVacMQ2rK7k3VunV035DCbAAFvH5GYNUCC0DKQzGxqruMN168U
PO+vv5UkAqRSXKD89CxSbkBItazI0Vbo2uoZGRVRrtdpZhuDtSGCi6poAKRHXbTZ
LOXirltfJAqjvTu4tNof+qLWlZTGm5baZbSUc8aWVf2obbPTVl2LPjvYs3jh62pW
Vzt7zCxftBzp2TXePzZWtawz81v8L+/eeUGpskMIp7LHrGRmVbQb+Gpyl2f5oVI2
l2Ux91Nbpyc8GiDJDj4hidOeDIVS0Hxr9pmkP5nTwCB5eswZAhOmf9PJNlilyNlP
9VAmkxBWcOd+7DVMu36Kzr2tgtcwF8SN0vpLG2l6muJde0SD5mDcOdasjtowGHct
69dekSmek70j2Jumf/X9JpoEFpKwiU2k6MLEbpW0Icu7XemFeZYH6HSSfqcRFY6P
jbNgN3m7fKCS5fdSlEmnBWv4V62Nr3aSrgHy9Kp6eTTol50A/tAVBcjCrFwF3wOD
yOM4huoeORrP2cjjMocMOdo8H1BqhNlXDUBc7bw7cwpD14fIZOaHOjFzbgp+FnOG
O5rB5pvGhJsKq8ewOCbKQAY5XaKniV8/IrvGuwBX3B1NQpesjyRdwcB+huz5TYaU
fXLzCuJ8nIJ7fhGlfDi1uU8GOiw/Wq+KZePMHhK4LdrC/Rw/Ha0RheJwwYVLx7Cc
T9qWTmGgBlYfQL9Xz3xsjSn5YjG7+m6DCFOqn4ZKZmtfzSPtV++Hm5OVgxZQpfGP
iQKjqNFeYDQrNmjwLBdahYrlvowig2XN4tZrWKNa5MqvCIcFTn8n9IcwYnLtG+uX
LOsPf9y+obVxUCVQSGjAY2x7GHXj1ndMwhNtAZpaCdpbIcgs2UFVyJVGhrvuH5PF
yzW0PnIvOsISYbdrITu6CTLVZCTwztjARPzlwgrQlzD8PMmgLyfQLSRxrv5NmJJU
g2Cq7HFwVkHF1VG0N2jb5aAyl93E4vdKH3rT6olrNTOc7kkvEB+6Sw6FHiDAVCjL
Vt9TBS4PwdLe3CU/wGXvtWYFupC3hRz6hkQXkiLGrsxHDMDo77qCcpKwoSLA73f7
d/joayEp2zSx72f3+qdvzcg4+RyGlhCp7eu5ns4pa0888lp3azVUb0R4U06Jnjs4
UMkj9QoBJTNH66uCyXvbldys1mQa1kX6KVYIOLUTYfA1wpOU+POFvCpYhe/4nbWX
Mp65jH2OZnNLQ8avYpJJHCyu/l6vq+UEvOQj/jPBL6uEGHgYdZ4kweX0jlLP5W6P
07UJIZrR+pBKiWFO5xe/0Tbh8sKVnAxpnzvECTOVXOohacYyRWMDsSHczjcrUxut
`protect END_PROTECTED
