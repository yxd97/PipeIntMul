`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VYF3RawJvIRDHoLPrSPrqGQlp+5i68RvjkHugzZuc83kpA0tihzAxWt8DiEJlk8l
daqN63eQdr8wKYR8DThr9VLk7NNnXblHT9zTRe9kwNoMUtRCQgKYaQecX+6FXKh6
/71Dcjy75hCrcA/bJhTpr1W3rC+Lf7SzEjkNNGoI45br1rI20zdqSUikdxn6Gzcs
SKRuaIqSeywQ5KlA9wyCdLtE2K/RK5qVF5b96MSLzyFiaUVP3oh9qZNRM/JJZj1v
jSaJSg1zoTxBhMntJxH1nB/fUNFumOjvnRJz8rMot6NN6Rb2b8Rn3oVGaoK2E0JF
lMj3EHb2tyY+i+7RhocgZelzJm0c6qnHPGMnP5k7/7Cor5Smi2LIz/jjw584TiQp
p2w2huwIIbE33KrIXzGwHjT6zGFVsM25UqWwE5y5fO8f4EJ03vBMbta462Oa588n
iogdkWuInN98BBhU6kOW/BYakwD+hpK2+jAodQByIzDUu4YBM00TQbs0KPm6DmNC
A6/BXk3NkHdE9l35NgTYcvx9T+xQ40F4SyO9Xya141edqG3fnDzHDaHA29tZ0/4L
ezcmVWt3WOn2G8ENHxQwKYqSJbu/tS+oI9QF1+7kUaSzKzbaDKAxq/nDv2j/A04f
zACemVXHuLjMHpOjrxOTUw==
`protect END_PROTECTED
