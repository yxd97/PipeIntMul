`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
EtBh5UVBDGeKibNdV8biDlWXn1kQ9ewCRCvICMRoN//yXRBuKQ+T2eIexKB5gTkR
gwWL1PTsKBqyqlop00mgeTZm92IYJZb+4NPNSNPcoiINR3VuiQLbXsedbmGsFan/
+0bFK6M4DRQfzQjsm0ODM8yZgUPF9KfX4JJSuLRCMLGG+7lnbfdzU4ZyFscSIJRj
yX699+7d6OLHjW+cP70/fNuWaKJFYN7nFgRNZZasGRGWrOGKlQXjvHBgp5g98THw
W55qgVq0VdcLOFL9PayGxRhYP1Xlk0aQl5BE2ZZO5yKQdEWpNKYXe8x2ON8rP33x
Fl8ZtoB7hrpz7M91WFdlLw==
`protect END_PROTECTED
