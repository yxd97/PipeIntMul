`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HJXedT/sas7LAtPWALbHgvdukw88izlKy5WCzmvGvn2lZEhIRjuD3XdUOL+5gfTQ
lAAz3nMP1XSd3nm3bpz/471fyk248Oma3iQdWY3U51dnReQNWI4R6kjA5JlMQo8g
KvrDQX3re8Yfqo+6NY6nPwUaPeX5lRvPk5zsePw8Mx0EK3Uazr7IfaeFFtTCnVZT
5jGOv2JxlEOX5mriyySub1ekFE3XjZe75Ly/hbCfBe4GtGqIKkfON94ivGzzqt8W
mxpPJoqKI2qmC5P6+cZ+WBnpkYXSP9EtwsAkSRd9HlrW4UWsPJv+mmgx/8ETdXY9
PQisZ9F/lOdBSmXUMBo9zefIVcn14/nRIkoaWSMHTxDdyeTEefMRn9xAqP7nG+xM
zq/j6s/OH642fCRsStzG2/fmugk77wFVpoMsWcZccUjRI+04x+RINkF9jDU58Gvi
zjSc6Sajp4fMEzzb64C/R5da8OU5S76lSXi4KqqAaQAFbc52wV25+VvpEoLVOfvG
`protect END_PROTECTED
