`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5w8F8zMa0eb0LN8ehW4maotZhwRunRA4riyj54LAmQha14aHGEB2o5Vd5APTgMo
dWFPaH0k7l4enu1setaXI9AToJhXStTUF3Qg0hYa8G5Z/rL7VxWF+WA/yOVMAT13
jmjrk6Ax7S5Y/cH0g1Lus5bgoa2vumZAuRVRRNiln0TFfJWM98O8XwLC7uwwQAzy
wMY+TKzowjNjaY32AnnWWmaFuHGPB5s9uiCrlDlGtpIFUIbHXudcDhvjOzGWa4pa
U72LR6kSBcuA9eVWen77VNDxdBQBvK+s5U1qetdnVYYNmBtsD2r8bWJIcXDEdAIk
RwVZ+bJezxokKLxWn2E7sfDnrvDZh5vDDg/m0KverWSFWUc6DgWLzWSt2ASrE32I
yFbqtSHEw923auw+OR7ummCguHvvr3edu2se3eStL2UF3Uhq1nwmpT4hjc8tuxzY
U+2kTZP0mDFc8o/EDQdcqZceEsU8IvcSjGxlvkYqPYx1xgBl00jBY1tkh55HJkey
bfr4pzSkI57JikcKqpNqNTmAClmEV7eKmglk/sRzaz9JiDMHxNZKO2txfL7de8Ul
bRfX3EJsXurcS632m2XIjGgScauj9BBr20GlEoW3qT4/LC2i6b77iRY7OxfAYVS3
amRYGwQfP7rSgZIjmu5PhMurnh+QyJv/jiaapzuSDQKTupWIFHu6lXP4Ax2bMZhM
B2btDZ+P3D5aiFS31aAP3OlHVaJV8oQFs3CuV83Fng0fVTe+VtRmArfCLda8d2e5
LNtNn1YjSvffGY8u/TGVlex3qub+UGDfCaaFgqT9LRbsr0EsEL16dd6hek3Ss4w8
9+7z1sHsGx9XxRadJo0pwPUMBdhut/suZBGk0k+NVgKxg13KUS1TQz4NVGiXkUyc
43dqrgl0n2g6yELL681iRyBafkNIr5oCnh8TYU4yJkLmLbFBKJq3JWMJnKp84MkA
SkBNaG0gopWLY1Zhh65QU8USYg2Z0bKnpOHkzQqJymI6BgJuiuk3X43q8nBWEGz9
CjA+RYScriQ6MheH8rNr17yJtTcPk/uTTMP+GNcXYspg0UH4TgePJOw+FlsAVZxB
7egEPUXAbTI/Clap30juwugL2yKpElPBb/H0Ds6NoSHOg3cINkiDBzF0SHjWqclQ
7bzxAvHPYbBF0IPwb82TGWWAh9s1KoucwzQL8TO5sq44Q799YFTePl2j5k2AUSnW
4NBpTTZsTlg7BpHOfv5zsDhTC4uwXBqC4fdQ08dlpYdBh5E8a9ykeEyrRERuZh4T
AxAWZoeP8zFOmOe8cskxyNBVTUbBv0IVuge93SryuDZrrOPiu4Ln8szMk++7WVWD
TGTblx11NLiD7d0PNj1ixdw7W/jpaPLKDy/tuedsa4+s5mwF4CCPWqefFk2VNrhm
5YocZo/19nyNwPKC1YHCih0Zns5PfSKn6s0WuJ1uiUPHQg+tiB+BsC+9+xYpNvRz
DKGzx9aYM3HpC5kMlooxtfZQOIwkiAxKPKPu7XPGFft7H1EJRU8wBtNGN06liE02
Tt7qRWjOo8sdzESQgSBjGfhOU8eKhuZIyr16FXy5Bmsn6H2uTGnvmu/lDXfia7I3
A2Rem/PJH1OEBj9jtwOtDrJ/DbkKWLvc5uX+Pukp8tSHwGatsG6WS3WszqQzhUWg
Zs5YsEjZwbFbWVAVZ6Rn0NAZomvJK4MP6zqArDzaD5JDsW2LDmZ2vTKG50yn+tr1
wUMI7h/EkbeDlSU312GCc+ROG546j95hIjDpROLgqpfQe6VSLQIXjzOKc96RNaUz
UdkBdD9Zf7gasGm9ToNFQQfxCxfP2Bj/yc+1I2ZvBeN7CTJv9A8Yu0Gn+NABqDdb
WAWxk2B/Hzr1LlIBhIjoyVbIf6Ypa9vu/EOacELNrZN72Ao9uxO9qfJwkkFcQ9XQ
8xvSn73WP6knlTE2riHxQBAv6jGvzxw80JopMuZT8g6jmo0G6FRlUQUf/mYNoWXJ
V4LkFSZ5WPgLDnUNsKs9aFkcCd+jZFsUY3yixbbZLupThSSxfi57xN7G8A0xBMQP
0EUsXzXkxsV35IT+pJ7o7QX2Hdoy8h5BEBNBr5SbV/TktM0Yps3yg20EBgsZA1kq
0g52OGZBjYURd5FFY1wlVaDlTaZNsEHEkDsUKOrgMw5uLiJI1pKak9d2EqxDFOlm
YPAp9CLWykzwb8WUy3UhbGw3lL11RD/OAmMMDCopd+8WJDJBCwBUGTb+Cm9Tr160
tS/s/f8FPlvF/sqnGmxBb2NN4pOqFXANKVD0clM64Li2WRtb22AqkS8xucpMIviQ
Bw1mltvi2eziq5M10CvGAXLctZUoJLsH8sShhfTYeOwTT6NO2jXVkAnxv+UfeIj0
6F6uGc/OCjaw6lt4qlycV1ELkyeg0iDmqc5C2SkbWrlWBnPuTJn5fOdeAhHUn4k2
FU2wcddfCxE1ZrQ671/YE1mjju18RhKs83rB4ogmtv/ZI6Y6L/nyrC2dBC/X9U28
bzHpVq8aNxyo440S8mzZQTOd5YhKu0bnoYwnchRRlEYIMvPtDHbhbdcXv5mhjhL2
cp6yiV+G0nWAT2IJ18CLh6KDeLFj1pw8pH2omQFd10XSRf0wNwVGCYtZlieRxUpi
ee71g+tOeCsBq7UaMCaHZDErI6cbumNtU/8Pt+5asBCyqxfd6L+8wQQWq6OTOU7z
rzRn6oOaeNYjZVAxyfDJpFdPwzovdAHHNmg5j93MQSDGu0gzcfpZCFeYzHEll+7R
KHvaKaE2vf0ghHw9NjFVr/2pistz4QiDiMMCs0lK/9H3ymCsM6Op0ftQTv6hdYoE
lZsCOPdukQnZesxaxvuNzYrW1AyXHBqfdtWi7T1qv4pBPeC+lWb9tkmeO5h0aOaN
Qu6wVhseA9gUD3BhGiEu82IrAmyaqpbmS3jqbDatshxf2I1w478KWpVzLzDn7KUZ
XBS0G8flnqqmJCntlaHb37fg9FxKzaIlmszEnLvHXoJ4Z+H2JwuYriCiiC63bHMB
WE00cf+VaXBLrAFUWIx9Qcm5W3V4yofcjQs6qXiylIMDoSMB7xNdI7kGK9q4U3RX
xAyhWsFwgiZzuXvd0qY9PZc5gdOeP2W5YCErKzKiDb4KyxXGoahf+TfbcAECJPH/
3UieDn9McrD+QxiqaMk1Rm03LsDMPkgyWn9ZhIyz5trvjxKw8u2DOebfxakmi8gM
P9YcL2bcmEt0C2/5ptqyeZbj/hN/9pEFy+6FdiU2TWQhjrIKbY31+oLzM2y0mGSX
+pbGGTSHsRqaYDTc/0wtkJT6rylOAKt6c9OG5Le/6IrbkI9AvJxDe5vHOxGZpvUL
9UYqhnEsh+BMSADdkAH7rS5u8P/9L0t4DBCTdhehinIEEHOCSkjm4zhg5EDyyiq3
lZSBnn/hlOAoa+IdbsAPOMV+kxjFTIwaHA2y1FLegO8lsm8DTM+7FO+OsRP85c/b
qoT/nlZCmIxCupwszAMJL0b4ehkZrwJl3UkxTfoRI9yrFZTRskSZYXbMzDxksA4C
F0R0kO9BtJPbntyNqe9Crq7mOfM3PqxwP8dVPu9rNk6kQw4HikeTswGE2dx0KdVD
lRx17nMXJ2ZGaiWjwPokHhsBW+MRRnZxwC55n2+uRf3MY995YDLOmCnrT3wPefuT
1bGru7laWb3mVh+iufQ0Gs+sO0vUg7rbgqCASBvHJATq0GdiqFRKlJtFaooTxnAE
cqlhQeNS247XTAVFox2iPhwWP5AY1DAnpfjx1WZSX6BTtyYPqxVi5bKWVZkB+B7m
oQeDB6cW1dqHg8FTsbOdvhUEZEMj9H5CqCQqKMMzDhUYIjX81mn5fPAGkwIUWzC/
depx/QaqqnZpGeeSz5wUBne92HkoJkgJsA7he8nmkuiaXoHcg5GVMMqQHHx9qFqn
MMl2DFB9OA+tXG8BJXwHKeZ7ZyLBMotKXRfLKQ1lGUP7HYMOP6//9U0F2VHEhLKK
bggijGksGqcDF9o0jx/7dX1etmdeKtYJ8WaoNp8T2dvd3pRpKg8YbVUNvOZJ2NOU
RkDnXR+onxJvSR1Ow4hs0At6r6X8ntGw5FuVawjcXFpl/fLDfDoAckEmtatV41Al
pLFYcH7+j3KA+TmBQlk/L35LhSjxpN7hPoLrHjtceWb5guLThZL3cmKD/rpdz1Ii
48V8MXog06HZXwLecNIcwKgsGh6LUc8VopubkbEnzQLxqQY5x65cZQEs6ztSY7+2
6uqnewAVwme3syItYF3eRNUv0o+MoGQKKkTztZG3eqJlc5pqE4ezDhRaPKC8CGcf
zPftUmveMwcfYFNh40VQzqepwagsd95Y37PjRPLMmsdnilSC45YdyQsdWB4fOhJR
43r4i7849CqIcYAB2J/6jE5XceJS+xLKCzOUCsWK6ZMY+rczjyANtkhq57Ylhf99
8m9/q21vY+qJdUdhNtX4MOQg1jBhtxfN2qAw262Xzo7MHCzXrHOvCh6BZRtIaFS1
5N4dIwpMkiRNvb1ttnPmohtm5bKopAegXHg43FQhJwN+wd40ePzOUjXZQ8ZsMAxw
ODoSU/+FJ4mhxXN2D7FfAn6iPNZDBjr6rXgki9ERgJ7jDJrXGPdhhBdJffeZLQLd
zaPLmiIqj0d1rYTCApRQjVAuWJ3prhdmHy5kp3nHuTmmiY71sqBHEg78WRhk3k7M
KJsc1LnpBU7xrxZ5G31FoGIHnFrGJxc5ks1OvQOcHpqCy1R34bwZ9hXnKqiKST+/
AxfkNYi3BNOw5z/Cfda3VdIkU6Kz4sPewDrHrddNIwsMHdNCemmRw15STxeKIPQy
4pVSW7RyCSe+nnToqNjxr+hOAvqFwa+zkljrkp9+MKiXIv7fDwgU4cdhPs9w58k+
8DEGM4xni7FMAA5RlYW/NcoFo89tKhmBmgBew1N82vKuFdntcPl6JlBsNWB3gtsK
+daAmxc14l5mSnXD0i1CZ3v/M2Ebq++bX2x43lIhdV0NjnUaXBBybXVUU6TF0JJp
IF8CogL8ApEzRqoaxDAH1Hl2HAqY+fXW6JknUDi/dOzoaxf4iPSL5MXO85cYVBvT
loCP4Zo05lL8soEIjwrv0+XRbmPxXZYUgqFjKZ3X0ZhBZl5bYfwACdV0YAOzcIba
oHw3peohKOxgUILNSNZB3+g/D4pRBPUjHCPTJif+5nGo8Th3rjfMBC8M4DLUMDJE
VfiRRLz59qEoOGDgdwK510Zm0+q2ISv3z0Famu+IoxLUAjqqCLeN4pNJBlCEm+yy
tqGBklDGD8S1cvyFgumyll4IBAUApZRZ0sWGj17XiSU7Yi6uBA+YtqPHQTZLkO1s
2vkHZ/7HVANmSWFHoan+RpcdXgGmGPKrcQ6GG7orgR0bSLiHYqqB9K1o+ukJWGvx
gy5PAssHXzk8VMi1fseyDLBdcUZyJM97dNrQJYeBklPTZbyvdvTqWlxXi45cUXap
8FvYIGNF28G0SaDcFoiBLV0YM3492FKg1wLxR9APNHWgTNiKls6WeCSUjHyorwB5
wINAgad8LifqeAKp6PN0Q5yQBaR/Nm6Dgc09PCLtieK4MChWECH3e0idnjTwhwmH
ibtdcnkTMVvyFug9sG63C/jkl7aBAOsAGFSSc6KCA9Ut0U4iZ4fqhETknwPQqfgU
bV0mk5tku1aMgpjJA8YX6jVdC2KpaysYGWzIcHGs9R32cxqIZSVY2wR8bVWnTeeG
jKBU34Pj68RbIMYEjAOr5VMFFJvcTshOEe7C+Z6GQ+ZS6rZ9HuYUziutvZCWVR5d
lzeHJpPRT2DtxoM1Vl2uBt3UykFYfhAydVloXYmoXHLaMnt8t2N/3LTgBPhwvYA0
oIDGcgtooR+H+C/AyccvSbMN5OERvXmCzsywmRIOFo7WsZTbMioRx04Gawj+cRym
5MWMq/UZCyQAgAvo74x19uib9agqKTjsoJ2xENMzaYRAB2j+SglX3/mNpFgxjF+7
uS29FjGqn0MJLvNdiOB3PdKkQ2TUMPYQ0rGMNoNIa2KfChOIh7zFKZUw4LKn2kpe
0w936bvK6rKOJPvKbAfop7EiHYo/raX6qvK9rvG0CBYuU3hCJD0GHJmUDthYNPYy
Bk2TIU6LKLW1WVfeH84EpxyBHX+acy1cafR0/9xieLYoyn/554G+Vur6+EfzF+7W
4ADmytxfI+Deomp0NXdQTV8XGacjwXbFpESt7nL1BBBLm0qtEtexfFxYr5eMgQ9l
uWPF6tm+4NEHNeEfHhl25Gz9vYDvRb2YdV3ErVlZySxJP0gVQLhzHOx11erucSKZ
NbeqyrzzTN+QL8UmD4yPKh76Hm3nmcMJwjN1zZrW8i70GvstSrOQfiH68iezt0b/
KC94Kt/TLvq+ipIjPXwcixTN/XKQaWMNRgopl+n4bZ4giV/i5P9TI/zhsstm0wlI
0Vp4HwCcF8zstpwOWocZBHXgyIyYLBqktzqPPcdQZMt5TdExnneM5o2TA607ha0h
ZXkFfW6DqCAdGDzBHtH6uPMCFcPh6jlFMkf1hKs2KpZieBMDzsddecvV2jeAlJ3n
7O41vAVOggLE4f9zWumyfImRsB0NhSg8POLEXat5rUY=
`protect END_PROTECTED
