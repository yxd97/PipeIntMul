`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6RiUZHd9zF0g3Xjj5EFo0BwA+71NLW5+2DAlzYfaB4UMnQGMFustcWlQFEkmBPSS
QFDsAUjXGMjr/GsC3DwKTR8W/IiiQF3MhAyu7gMIx1P2E3YjoVsHe7juYQY/ZrCg
POCoVzUgs4+nisaUKoOIwxBVp2LeUwZF9M0UoamqsK6lP2Dr9PK6tIEItP2/dcc8
Wc9AJButYQDjUxyxV7TKNVwIcqBE6yNqheoT7IoIjRERbHi/mrYnVgUlfgqXj2aQ
ciH9csiUxjiKaQhfGd1kPAjIu7zKHQRBHFjpv7gFm+alALJqNAgcdDcMnUjoxkGp
atiZp4Wqg2jmKjWesl0XtlT7ggFHkf3hIfBBaXDt5eHqtj9qpOZeXxv0hfesyzGR
wzx6lmFHGZJXPrjFsJA+xXNpJGyB9uzS7x8igswEE6b8rE+vFJBv3LjTfCgNjynE
hrY/96B4+ZHMAWg7LHRrmcL7LOZLcCsvNxcSrP383xwTESjJ6RFFt+tUE3xbIpAX
2K/fGntDDffnUttb+QJe7ASY2QiObuKPBQ2DseLGFa+ESeOsrTzfk9fz3BbA559v
O6DJ0MNRjjU44jPKU9PM+sVwyOZDmQCvPoyz0JeBTQVLBnzmW/gaquguWGdLNmYa
5qWSmCwCOk7pJRfG+qrIGljxJPiIN8r9uXjM2TU5fOEiVrM+uHQPT+9cJdgSO8OK
ntHS/AN20R3fF3PCu/klou1MiSss6osoB7zpKa3yIb84XC4FjIYDmoHVnZrfuijh
5wIZUh29dhu1TJIiqkeinpH475GSnIunP393jc314swNe5f0Lz4LbhNOpq4iFk7c
UZPOz2bKBu2T1LmHhM791kQWMcef6HHxa6ZpukTQjhgDclDw8OGLB/SGDKqXai6Y
QyzBHCcxYdNty0CGEM5SmQR+ojjxmD8KMQVTrBydM5GaXeMHVtyAN5lemqy5DG25
bA1iLyhL2rib7au7ToBn4f4iaWP8pQFj7aHLsZX139/u30eFWF+DtPon59lwS7NW
5rrNmeWDYTBEW7VIidoN69CVPmUZAMeROBAoR9j9erm9YsB8bEtFw39YIMsdS+DH
9OjczOFmPAZdfxKHiynCm3g8YMQfCY99GDsrB8RshnXMRk4l+C5vyF3r8mIgNP1y
nKghO3cDtTucZ3KiN5XGFTcEiPbZ5PqjaA7vcLxPTO79HS/URss8LvHqRYadABIG
iiJZnIqcRHlUGqEhkrjXDBJ0lPtGsNyYI+xZO8DT6EtBWc0swJKEWZ07J9TMBzHv
zAgHsaBX93Qe2zYPX29cn5HzTQNCgBUrYOFNHZnvkUeb/1oBEG/lxnFs4MlDxjLJ
I2r4WhplrYh/lpvHIIhEN4wg0lxcy40tPviAxXymCTlPtaCNPEiov6/IBhCFFaJ3
/49SamXC8WdkI+ZB1LdL25EZLItXPCT+pAgtTiRezfoeUC4iEjmGckMu1UeXGeUU
47zsy++d+bMsGGD81W+0ZMlseG1PCdQZTnoj/QqVJplWucyJtLPLbyjo8hKmvatE
TQ1ZNZ4LOSIPJPl3zoHeu5BxygZGATSLmeU0AenA/PzMqfjOUhl49uDBLfcJcSs3
JNlSpWzQwE+R2Ahz4TwJPRqil8R12+fR1ViGbqIOdl8puQeThB08rr/Jo2aRqG4x
uWfnOItA42yCP04PHg/Kr6lVJ8VZ0H26p5g9DM0qREEPI2Y+ym/uZSvm+Vt4HuDR
ChmQkx4cJywdtYXcyIv+cD+uUj+XT4lXdb/XbUgdsP3RKSQqE4syX7+02+GsZHzg
d3drL1VcsFYUKjbuzwwLTjOLv9z/HmPUWqlQb4zQLMlo4tV/ysHw+E/TVzXZXMT4
GuMYAYZvsI8fER5eQMCzaywlTUAFK+MJ97lO5J+dGt69Fm5NihPEF6NVwksBBVCl
jV1hU9qUPgzGxx39gKC2CgcbJLxQ3HcKKoK3wpsYzYA61LhwOvHnfnGZ7s3SrzLF
MvADHI19DuaOBfn07nWi0Nn572ugWAsaGq9Mb42tI+WLfxIWSQjh4+SrEr4yjPll
fCfrWZZH//x0bXVz7Vh4TQUdKWBd6mhcWAUwpOrCAHYQUamGIGQdXXkKxUTEW4S3
7fwqJOlt6AO+mStQlQbFkz4XydhHQrHJk4E0+YZi3bJzN+RZQYQPJcgVAsAyEKSh
jE1GMlbfKlQxGMZEPVdalT+ULNSSgcpaZuTPAQRs72C4PqQN9RLCYdj0+7hHgDlH
2fslQq8tcs5JNbjatba41UHqkCkZOyubWprpJSJGQx071hSMCULQ6ddPlILjAn8h
smulPyAREa3s4U8uV6CYhcOX83pbstnJl4JcsTC2X2ZT7XJO0vEf86lj7WWTz4+V
Dtrm4MJcRLgfSUzlQT0yfSsa1kyzh508rdPwdwxrzFak8zBUgCWffzBKoDUDNGzz
kF+lwIH2ZjPi+9LIZU4ps4kfYOhyh1LWI4EqB8ISlM+qg9AKfRuztFxQvmQCf0RK
y4/+AyPayu7AEhxbE8Og/PWwO5yYn4HSf/HX+mgjtMutfQY8EYHoerOPLJA9Trf0
IkgMiFLaCaOtxH8cG96n56BTn/Sq4PXOHqKX5sZ4/jwCZkxynoyeaCXY/bEEvSUN
/ewOapsUOj+TEVVYOreB3Ir0L1M7kewoc5g8YoSKCokQKwo4vPbUCP/2jTL2BS56
nQDcmTKpeF2pf2Mb1FJmQ1rMRhvf6m46DJKr2n3RYqqItqIxQwvdBXtHhJkMM3r3
QzT5TD3onEVopFMQoatc4S9oCxt6Pc+tXB0r6bLYp9kJL+CcdARiu45w/3xtafAY
xW6W7N6SxHC0uZCzOLLd2mwg2AeY3dWeF+MRoQYzybHXTFg25IxrBhmv9ATfwDCL
T4U65+FBOLyt+nQQM2vQPT8aTqZ8k/a/izoVGxz33dyLCBfM7cOiSV3VgIezZD3g
J5OCmfmECStVr3Mfm+QScFqm9VF9Vh9FVxx7f3YVqWq6h+FME4SYFbFqQMLy6ram
I1PTUx3Av/ZjEZ2eI6ILVKm4UPeI5ZkDvI55S67rWqiyeT//3DVvrn9UW2YX6D9r
+wEdChnTdZtDAmgK/dmh12yZEGCX/2MYvA5CJja8Z1O6ASGm6KjYgIh7qNFTwjvU
fgGJl1df2WkJ61ZhINl/Urv8itEXtHAcdBLkKKJH/skK7uRZ70aRso9yLa+qiXAV
oQk3Ziw2PFEdbSwf9WoadoInz5c6KTjMV+Xmpu2jxkZ6neCUFrLrkhE6+3mt0frK
Gt0WrB8tFI1zwpUf7rTuE01GMJ0GpsA4QwhlkSF/pygQtHOnJXR4CDE88mu3EmIF
7UI3RVL45HplDY1kzyrIbzCwDOqYIcKaKN5thsmhS2tAjAfBdLq7P+TPrBOfw5N1
xAHMwzzrAwLxR4RYna1F67PBJLfruAXYu3fueUtre3ELQWqd6NvkpSO89/azD4GW
JF3vNFvNp0Qnt4dpOwbfML6Yjd7plgF1BuF7mYsKOKTKlHZbWcy4cm6MWw1CLiU1
MFUwLcP2nO9IMS/MQgvrTduU6OFEuRBxCQAknsm35KDKOq0q63mp0Jlr5kZA5XVP
I4N64kp7C60npGTe9k6mNr9yqz0eTud5V8pZXqqSyZc/myAlddDU5yWbhxJfb6Ue
hGkj8g8fh8byBjAsG0aSr15ppcMt+smhEgJsu3Jr/MrPsfOD6Hnps6ov2541nQu3
15XZ1BT5O3ndY6n5SEZyxcsCwyqJAFmHnry5VadWcmPEj5i8auRw1WTLAgQho7Sm
SdFIEjJTY0Qvm/LOPilzYIUcY2xJE1qVqboBxfUhOu46KZxvYeH+CeHZQ9XcEQRR
1raSD/4MkcgQOUQjfU/w1KI4IsKERodg03ghrlzKTrlMm/lutw+m7TcdV86pY/sl
VPrRiQ2fIxKD6/8t06QBbxWn3SW6tGTaHFDngig0/mLnh74dUSZwWxb6HI6d7mag
vF15vZAEgEn/cvCqdZhOd/Y3kDaY0nBJRmwEeWsj10NF+EnoHfumtp6T0Kt/PpwI
svyxS0xFQvMc08H88DSqNxUhBuoCOkeEoHPS9WvHXM82lljNw/U4MJzNui6WgwP2
a6dhYmZEQ7X4nzu3wS8T9hQEAoTWaRqNr5JPZN7HTwqPRlnnQX/4s4j8lf+QWnhY
qQo1pFMlLJNKcgyo3N5zP+2SAUJJqFslgz2AqqLxVzyufvzcothTITVM7XnL4KpI
OlQc7aA4NO8b8UgfHsgl7KVc6dVqPWdylyZSoILTpDyILiobIBUvSJUVrg5o9PzY
1Up/Gxs44rAd/xzTne8mVw76fIFeAZckHwS07m138HjsQBtegIJIF/q7R0f6X8Mf
khxW7d7KTtEnBEAXqr7VXo6SiB8rm+GMR4c8glzhRjAnFtFyTpbJMZ6SXB2IyVY3
wdZkFK7BA6WKchOCe45pAPhuzGX83j9ft1DKvGDzh3uThqKFfuQLI7tP2WZpekbc
0FCfai6CyPkF1N0+0d778Pr/RT2aq29BdDLIsi+dvvaWJFsf11u7+uRIQh2rRCJp
JQ9upyy2G80uStgDQMWzibiGyvg55oZMeXjzzNjQIVpmDMY087XKE31QCcNPdSCM
sNlXkoJZjpv4/rn9wtp5/nhFNI+tkpZ1E7sBI/6YniPyH8xBqADC7376Vm//zSI/
3ykSegYYl4EugYz9o4A+IR1Bbx3qkX+yjFhywF8rlX6NBjrxgvIiEAfGkOK0fh/N
0+CqDl+Bj+XMiLcUEnP0ZIu0fPCcudW21BDjaEd4Ga/qYCosDdjOt7iY1EMt/rAt
Hzar5lpXvDkTjDYSkD7KUdvwyvGTTgVphuuy7bA3g2RWbSwTke8+uGACuMzgLxiZ
dKcprhRGruDSQI+sYTi8JazMtVH7957Jq5LG1Ga6bvdRwufmw1DWP5DO6GZgp2Ca
k1aS+iyIsU4n3t5mn/sFLKdD54ISfCwYKalI8tmUbE8pyTylzSctFBY2tQjfjK5J
74oJ0IJriL8pb95j+UOMHcuQ6dnzEZyUX2gBPYqIwFIwLJ7oMPqi5nqpDDMr61Y9
3KUfD89EFyYUX//EqeLnqBtkKFh7gQ4Nw2d1i/liVv5C1Bn+uyY1bQSoGmysBmab
Yx70sHtnSgW+jkVDVVotWw6O2sitfTWLe4Ft3XlsKeSfveJLo82rs8V8Z71R/Ahk
TNglKQ08OhcU8E/u9Zue5jyeEsGThofNpqLcH2iwC0rdoqBZxZ2gb5eP5v3S9Rja
lRskbFEuEYiwZr+YhiQPzEgw+ZLyp9V1T4RhXQ4NQAORdWN1aDVM/DqQR8KqQEWm
VJJ5abnlSAr+wvktpxuc7gftAGXyf+EGUtz9xC5fWuoZdKQ9GXXsU0DXNClfnrbq
y5ul49Q+O1MAjATftM8hRpfAR8I3ZHExQXsQJIu9wMUvRlbF22oiTMOFOkJOG5NU
qRV+qlhq2NimStOGEP/dAkTAJrzrh0NWA/DS8XPpPTYOQdDDPlLJCWVEyPV4QkJe
erEktVHaiKjVINgMLFnm+Q/YY9RA3a0yrygxtiigP7Y8E9wdS6Kaz6JOGHbx+jHv
utst4BVX/O0hjzAFftfN6RYvlCoJJ+YmeVwgimHDSv+sPiIKbrmYRrMTEZwzf0LN
5OeD+gB46m5JguUWSBBtbojGtp5VxwEcORqfhdgawNM0RGTOdpyHsLlrPINpjB+c
U6459vVFG38vvuj2dky9WHSw7a8Yro3RoQNuddWR0UqFH9bb6I8Jj3rGURSa+ecI
4hB7r01fWOdfr8Ni1f6EQT0UvLvPlk2Oex/RaFEn8J2BD1zDeTycuIsKkgej33up
6Gr6lDYGxJgkX6+TQvNu/WaiN5zX/At5Im6vNglDK7Yl9j/QCu6yClw7cLwHE3u/
FKEzhD5hU9wp+RmKqPaHM9CUZD6iKdVCGLNZ5+W3HLFmcWwth3e3SirD4RsVWA7O
OX/AnHyjyLpNWQPtX2crSUq7jlUbIpJ5f52FxSppCgnUXh5QCNJZ2FexKAhA88Fe
p7GCQ+8en8Bs4PslcubElPGJtyfC0+QB9xAiLNKdBAAXGsCqqeSikD8a3iZM+o2h
00njGy+wJ/FKU7XsqBdPs7U6la2+bvR75XWRAINsGEvJdQ4P5YwhGRmc4hQ5jj8T
o3vA+8GmyxvndjnVAm/fYEXrDPIyKEGNiLW+QSM0BNTx/a7472eKmLdyAzM9PUMp
qEU6mBXSwgJZLbPkVdudTHul+prKCP2xgoVOhKyQIWUggZx6p9cGItsZ7zsXl/hG
+2oXdvzlL8uEYHT/0kejSwsDI//1QVBu/VtJUZqEgni9ajyKiwFpDCVRKLrpS7gx
JhQ1VN5a27APu/QLJVJf0sIn8FXLejmh+EpR9qRGbe++2n3moqlW/ofkHkDmkiZK
8WKSnCp4XEBmbcANg/UmnMrBAnMi35gFquvjOkNXSdSC/CYXE4qnNVmc7X3jzHGu
YG88Zg5DO3oxKsE2fCdeIRCqMRkeZlLQHF1bwgk3v96/NkFxDa+YagMHFezRBlyE
9bVHQ4XwIWThBbLNaX2yvr0NbWIQCN6cUS1qfaiDHxr9pNcFuIU6exzojnPt4Nd0
aho5/B6zynZXWt+TgEodMHWtg5bgx74LqsWKlqP0om13LbLv7sjISsm6c7T0sAI8
0wtgh6k4xuO707rxeKCxDj5/wdhYHsHM9tKh0EKB8XmKoZDcw473vzK3WawS4jkl
wnZtuu+GwiN3sAkzxxcprBV+OxgEmQBWe34PgE6LrDV3gjHP5ipuRpDQSKhL1WWy
AxmbddWys9WK3e80y7ehvCv7eaz95Rzz3fnAwMV+UmRWcfEFvOSuWs2q1H5bn3D3
s3UYjOTrvl5dgWVKLp4p/QSMCnc5Btg524vaL1uL1w4EuJSR0tK8VAKFHsjc064q
mw0uvbq3hOT0CI+XngMKCFfSYV4M7OLEH4wsdDj/2bVigm+v27uG7KJ04cNENLK9
O/d3/qSfWF7ymS7m9u+6DWo8A7fWWr9wmXbUV2S7/Amw0X5pVmFdE1iJ/mLgD7oF
/N/AeSjx+MmLrRCBOp0xZ77MNX72B0RfhuLk0HrrTFoc3Y8QRETMl9z9DSbVuxs2
rQ49Tn8SF1JNeGOqHIMWTo1zLkTmUwhG8P3eClY56ZVOxtwbZ1d/TruePLbLh9H/
DuDJuku3SyWS/s9hiCfIrnlTALp1S7MfWOHY3hazOIx28IaSESfTfrm+zV+eoB9x
077+lQLiIlcnEGmwO35i3gRJ8RrXh7qf3Rw959ZCtdogSfAi4gajlHmf6Gr4DJ9R
JoPy8vDbycP9g4bW2q8ec2yNBT7iOsx1d4RKAqgobEGkRwyNOc2CHoRey0oWybIp
bmBHX+0u+8x9fQDhW1EQveq16xP+EA0sgggBUDjT98oZVnLFawKcrmX8I7cFUFp7
FoEAyXeHm0trVlN+TC/Mk5zss9ateV2B8VdO7OuESFRCvFayHAQUHz3afmlB6R6U
FMaMDTSDbv9fkoB/kbmCaCtoj8CeWLQ8BK25bKc+ts9AA7ymc1Dlh3m69piBYpaw
H098Q8SEYdHj1liy+SrGWNcV5JVXn34GgwfienV3KhtMAQg+Y73KQdsv4vDYU3pL
LR3/iHaE6oomgqQrA8PxmDKZtksLfm68jCf/Pgly9Mt0xtSIS8p+WEOSAvpIzLNB
qWQnA4Dq0VUsEwIDsx62QHBXWc3Vzss6sQs2X3tVhd9iLGP/Q9WWzE71AIeoaX4V
9bIFv0CVDeEZG4CqtkLUXMxDfDyKwNH8wgO/IwY9x7AWN1W80PKmFJyN4q5WZrig
baT8T+dnCjAwQRzP27YwcB66YA3Acg4pjboo62sUPZ9VcJV5BoDj0d5fGtgl9LlD
6tNhSrsndd22byGqD6NeoA/AwOfxfw5Pr8+cny+LVIzGRW6wvBo+2imnICy6L9cp
/bvrQ1JRKbQD0sdJwTnrypigN3pyy8zttT/ra08tnb3bORxl+HyuJofNBxLpBH0/
U1f5KgnLyUl1Gru4IH1St0L1EPsTJm3vFM6AQ75xf47O7og/Wo19vz8LPup7hwTQ
R54VC/4KC4xRjmvlVF2dgJYL71kCLI4T48Xa+hLHWH6TKalEF3xzvRwNoY0sXlzA
JuhKG8ocph5Y+UwDmI22E8S/X+Ow/J8esXNsZLiZ4Jg=
`protect END_PROTECTED
