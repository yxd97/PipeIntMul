`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gOGz/Tngr9G9aVZHLRUfRp7KH0ct/Eip/6SsOEGMt41W2eyZm/ejBJCdbH56Fvgu
mwk0dqBghMIRuLkY9AtMr6X6M1cj2Cv5kRVB4Smza6MdUmTVs1J/XZcu56Nqoevb
qp7nrqDnNJTtS5pA6Ois6KRamSpsJT92EuRbTy2NARrEvTWiQ4UclBkqjboQhYqj
pJu9YXJB/fD5UfiE/bm9F6N1g+/CmDjsp3dZxcH8blXdQ0+Ty3XQGgrOevZXg79o
3Wcfa7hx9JN3YvdRahttUw==
`protect END_PROTECTED
