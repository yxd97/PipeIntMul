`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/JcAqNFh3lJoupOlIhLtssfD0bYKKfWS2kpuqWpyh8WnI0Uffa5nivTtUBQsGm7T
Y3i+LxIfJ70QlAtHTcddkacRYN6zedDzHdyBKA3hNUc61BtgzrsOoMdhjcyyUujT
Le1xeU2euF7CTCUYx17s8oBzHtbBzoQdCElFB3SvXHUvcSV8V03+G4GdOgNdcDSJ
Yc2uWt6obHBGKkIozJdlcYsfzVCh8rPzOYO+P5dfGz1fq7rr9nlg7H3M3dr0QVMT
PMj6SvWvwAehwhn3l5Ynlcwbi+zjLRo7g8IgXuQUjoXnskztM7mzdsB6bBP4t5yj
ntKiYXmrEHnJGXI2T5goC6tvtCxUwaLwFY1Nc6aVchjew/qMZw1zYp/mIiXScFYD
VDUufrzGS0i7HZUDB8YQ9VoE8DecFKCAHQX79BA2zQ/+hY/DL/jZDhFnNuiuLMcP
j4kput8stU+2p3g2Jx3cnHqRp9adNOK/4Ao12DYR9qV5q5tYCg0VbRfKoUKNJWcT
ClROY7Hb5TuMR6aA4N78/leR9FestdISfT805erb000RbRf70lKzFV+Rx1zotRql
yFcAViLVBwuhRUNzIU5e2oLv18Q5t+0R+ubXljJ9xh0M+bIaiJ8aemdplAzU4vuH
Il2dLR6406IJAFjZt29DPHMJuhUBth8yf5J25hgjKmAMzQnG2d46ImOq1plWdYw2
ZE56Gx5pu+j4Fwzrh5JFZFwuCk4KwWm+aL4114kwDuGZp8dfZxF4Kp/aZnaPgdTA
6sWBDMqFQ1VZNOT9pA/jY+/VmBTBKMaTL5s6fN6L/0tZfEVUZ2HBbENdRRusIfrt
px7CsAPmexRzHvigh7TMexVuMSCXOKVGI8syVN/eJPW1M0+FkWu1n8MiK3segawU
weBCevXKTm0I5f2wfcI5GSgwoldAOo1qzJGiEndnuf07lE1hv25dFpjwZ4gpvLIX
yOGimcgKNL90VBWZDobOtAZ51tGqh5TVqEdp3dJaUxtmKWGeD1rL1by+qUn3QXuS
MDBiHSbiHwEJxiGjLqEPV8nWaJnfOnUWh0WwFvIzv6+pWjla1yxsrZYMZyy1ZGmi
DgCjVBMiuZsUgEIGZn+UDAmBBg28VzBxxj+l5XvQ4RfBpYx+28mcLCrImmXDEMDS
4xiIr8vQ33KX/6O0i9/x9X+K215v+8mENj6KujwBtO016Wfspa9yISIxUlx7ldUe
epkV/NdRYpW6qsxZ3+IYDT9gBa3J31iYNTSw7wKUI8aWhl6e9RznxmEaTS8xXLEW
IyHJ4qbHsmz3t8Q+5h32x0MaIuPTUvyEvEH7gKRbmKjk0kX2BL/22VrQVYFQIyuW
wXSSgv2fAS/4ElZQLmqMWm7pMUAweYFEDXNoyUZc+uzraauPrMZNdr11waK6/37b
aMaPaZE0Vzx1xtcqUXKth8nLJgJWuIu1jJNx5ukJh8uscCPGdHuewh+0DMLF1W0q
uW33tnts4kxPpE+5NSeWCz4/2dkt8i6+Pmk6CSnULNI=
`protect END_PROTECTED
