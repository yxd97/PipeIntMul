`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gjr0zyKd/h87x2Ob+q7HXQ/5BUs1wS8/lb3ZQvr3qGd2T2nPYfHW6RZ9SLb0Nf6q
H1CjeJsSEb81n7snO4D2j0QndcgBY0PAmPYofalMJlDwewGlYoLqULEU0kbtebVz
bZouWXNjHE2e7Dz5qPRYS/Hv12l2P8LFrNVsE25h6/JtLS3Bi1n58DIL+rvNN4GE
K8hV4uLQgcLauw9ipPQgbHUlzhGoJArCJsseu4rJ6KO3a852UiWbSS8CagbENbuE
IR2GcA1cwaFN+G6hGBSmyCGGHoySs0kjXOdnttnszy0Ykwx7FQpolu20wlvIBcS+
pOmP4YEKnv+XOaZHN/b7dE+b/Ywh38zKoQ8Jfetk5T55hF5TVpUoo5nLmJTnPgwZ
3X10Y42NZsivdORv5mwVFHvXxtYV4z8NUJQthB+sHlS2wztkSshqSsybgzjfkAzx
z5FNQLH2DE0gieH/aRLu2llgOf77AHN4tFI3YDZNbM0dY0sttGtmV3UB7AnWVdmJ
OusJzirnWFHAM1dVDFrl9g4EVUS1Ot9Yq9huPtsNMiDbNFWrYvrlVbKl799JAO6Q
RHKXvZI7dQ/NpK3vWVlMo1/RHD6Ri6IHGskxpEypY/7Buu6Malt6hcG8vi152aa5
uF3Er3fuAG2Xde9bi2m5LgKXumbSge7PIdjl3HMeB5VZilZNOTJA5WfVCD8RQ9fs
ruLP32pPVmJuRFwNUJEyQtpgG4olRN8Y84GdnH7bn+P5lyv0Cu2suy1e6t1P1aRF
BqVbsc/fGUqo0xZ1YEg+ZDKgGKNUekX1cw9sfI3n+/AKFdYuxp5X09P/hZXK7pte
0Ul8KoJ1YMq7S+k9TQqXhxqLh5hwBkcsK/7hcCYRsxB/qv9/4rZM9W9+O/czNMiA
GKo0Enkji9fvlICdVhURb7cVBj/spDcmy0/caJQSRgv/aIkGaQ4Pj5xYQA0+tt76
3udSvMuodo07QemaBOnKh7QTo6W+OYHyQxXGV4YHwgCIK3SiaJy7V3A8cbCc6OLk
bn1H5Euzhn7w0l09ms1pZqbNG0K1L9yYban99R8ZdUfQGwwsDqcjEojPCVeeOYFM
VZXpRgSiKcSKBs9MoySVLJ3qO0Dab9YbE+VUcUqBzZzvYyvkuL6ZrTpMZsBB8C5s
`protect END_PROTECTED
