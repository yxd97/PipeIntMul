`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1g8Q4SIn3aJDoZ710IQxlO/pO3BaVMsj3kCNua81j6aV0EG1EMbBHOFDP5M4ABi0
rf9fKzmh2TEpCEtRaP2WUWOMQ3yXRZeoS8vn7WluO0XSHX17SFe+FtTZXY6Ppyhx
CIYAp73s3pQgVDbng3JMhBGk/LgEbZVN7DIuo05EJoonlc1QkQs7xLCS2Gadvdy9
QZg3fYzNSaKzFEc6t0KM5UkGLcxRGFRO3M7xvEFBNee223R0ysOjeN1aJUgF85zb
vjlU3lgIb/0DGP7slACJXL2p0rJm9hYE4RdP5Q/eea1iN99p5/5HcATm4y1QqEdn
`protect END_PROTECTED
