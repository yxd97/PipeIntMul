`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jN3ab8XidEaGVrI+aIYnn80XnMYpvHlFcZv8R8q3d6EBnJ/S6RdbrKEmm7wtWa6W
wPmoiobLCz5lZulKaDKkj/k7pYUYLb1d1rT+AmWYX5IOUyx4eqFOr0RXmLunKvTO
dQYDAM8rbe+XinM8xaJkvtTAmf/GBF/npWinP8fKUSjwV5yI160V9mzrFTKBi4hp
TjXINlCIOuPrMZYOgXKK0rvz7gmzSfsEj7ANzUI6btlCZLgt04a6bB+PM3hId4WY
y0UMC2moOp3UREzFHG4NuB3pQc3ll3Kk+uC8Nw1oCGBoBW+0VOdlYFxo4etQfd1t
fCmc0MqbcnxB3dzOKzUt2nCe/PapXJLdrpPieEP3C+IjDU27SENxdleHostAdUTL
ad+dMj88auPIyR0yzIPADIs8ncx9VPDwOoRAluyP6AVjf01qHb5jMbnwQ8KTTnDw
qb4OVFOZIZZ/pGa+m9x2Rz9JGXYxRq8Vj2qQc9hMo7YC2x34Dq+9ySpfSXOrRhMS
VwXZht2nqZIPNEMqpr58LJFN6u1YjQ72raIApAenUk4WSv7aF3kCtwxvvZ4xFWOg
cpZBzTtzrZCRUd7vvcLHaSKeyq51UjuvKfJP0MlAYWQ=
`protect END_PROTECTED
