`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HD+YlAdhDTz3Ga7gDrs89OIr/SFWRyvHKek7RSqLcsZNrFd/PB7/aSBaGEjqVGnR
Ekv4RjABfA9KADxB5MdBwr0FpPfKbMHIe8M1xU/Jq6r4FU1/JTJjKinv7HYU4L3s
ILAYFGamnT4FZXOj8WS6qOaQ1ASrNSJyz82ENuusBEE/mQbI8IjcJ0m68nOiVkV/
EZnvAekDLs4k0B+5BBxp9wGNC8EXv/fmS+75s0NKys+kT6tIf4zSSfSMOB0DuUBJ
7F9cD6sAEKblj2kYrrn85vS1nOHi5G5c7Vm496FQhkX/QA1YHGU5PeyjVpQVp7KK
1fd0CHOpbZAzL5iEJSf79lilMbHT4FqS5h2O2ysSQysUPaZlSz7XhlbNnGqOXqXO
ZZNBqP+HGpYWKaw+3MQD8Txck2FSarJiRId7kXhBlOq4Dvgmr8vj62HLtcZ4xoIv
19xY1FVE1WrFTow/ZYdpiDDZBteMnsdECC4iqFUs84JC7+6UJ8uTMnsBJzL2oaHE
CAFmyF4RrPO6IL7Uhtk2U5aRXHnOg9CHV75NvPApRW0k63mAGTrazNeUnqhm+AZv
PTnMwtD1UQFjIjw9h32/BEG5hqdRoubS+IFZ2AhiRTY=
`protect END_PROTECTED
