`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kxu6lj6VcmBNQTBIj0LrrXBPRnD3wLFkWyXSyB4p/l2qFKy6g+W0yrCccenaeTid
3GxyjuJx8asE4ZxIlTQ6v2d+d0lLdL4uac6Nrkf8udGwL++F8k6sc+HgosZh/+RV
YN6mxKyo7LBGUGLRqCDEoq5WehxCGfDdhLvjui+zBPcP2R9Fa5GdNuZHhwi/MtZ6
Mq5pzGjJyjhaBoqv5NWkVUnhLy0sgrUzCa5/W4Oj+s2kGQltkyzvRU2KyDRwI3Jt
onaOsgx8bMmMlLfrPvAWJUShZANtxYwvnC36TGgzHJoqlGkcnq9ltl0lfM2bXHs2
8cTy5xG88+XBlfAMt0SUVUXSgBCIOFfBd/w000x1KmIoz2CrY9Sjd7oMR25i29BL
QqD16Qx6QdjJ+XrA40jcR8ZmOTJCm5Qu64KNZSI7HI4=
`protect END_PROTECTED
