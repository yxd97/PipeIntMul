`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FZ6pix2dJf80UjjSK7q7pRhMXfTDXGUnf6DJRNtxSQrsrg5MK2LaZW0ttMLUnLVk
vFE0VKvwt82KWtkRZILVVeTHU4sB1I0fvbi10ReJCvOlE48FMytTGAkw4HyodWkw
oelIwJHUacPGzNhGqZ1lalf9169D7h/Th2FYfwfeo+SJvw+8H8iAupnhMbeBWi5S
kLdzJB9vruqdH8v1Ygu9p+Ywim7z7fiZWe4CswfkLlfKo4Kvty0EKFtfMNDAxep8
yM0weo2/zTmO4o2JxJBLYHTXubZ/e22hZgGGIy9PVMAt8hqvCX5EDDEWV+cxvV1D
uP2nBivU/mR5VxQm6IDaCojO2RbWw/+v5NEdNskI7/avcftYZxRJwGNMXKWKF6Vd
KrhrIpENGRWs+NMFrAim8L6LHlaw9iQlU3dOsZ6AlfLaHEfRz9UYOLiPt4rELdUP
4kcKlVTnA6etVOFVrBSFuLDnczwrmLSsuv+aBlgyr5iBPv/2q3GXlmhMEbchJqSZ
zXdkaUK8QrlnTSNPAghtAzIowtWKCrCqux3F1Lw30VemKpuIadq43RMEEXLCsSbR
km/TZL/Q+36JgGeNYcejtkJejFEjNb965NJxRQiOlisTGTF1dQUgwg1hpILEQ1Jg
cC3gNnyWI/c2eVgRb9NVEQwh8L8KloRihyIM8DqhW6HMM2hwMWUko2b+c3UeBlS2
7KGXOTSwp3BDouqd0Y82Zw==
`protect END_PROTECTED
