`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fEbIr3H5q0Kj/hmLMvig2CqkJKycYJEFXxMjgOI0kKy7LAglFwmAPaC9xZFfH0UH
e28wMnW1e5i/8NrOMWZCaEnQrw+gzfi3Ij2Nt6NQTXK4qhwfPBASE3TdT28xo80S
MyBxd4zZLVSKG2M7yfAtAm1nzGjCQRcdkg9ykKNT9Rd7I4YI34jC70OTnhTI8At5
ZwnloUGvrkIt/FUavVyOMGGi3avUkMrGWWUgl/C5ko+dLUoA8eoaUzbTis0Wk3iu
bCQUH9yLhosU480jyuXPeJO9fNGauUJhcvs7OMmfl+3q0JDfCia/ShXJKZFbnK3w
kKqqnKMjQf/LmtqwBCTejIKPO8srbKu+9ccJgEpYRuM34HtInwfulj9PP+55O9Jx
jh2Ro8E3aYKyP5hiTROU5w==
`protect END_PROTECTED
