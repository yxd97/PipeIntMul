`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
k/URN51oqd1MDODHEzsVjxxP+zyZaTKXN793XKRNsu8AC0srXzrWfBExB6tGDKOx
KPTTMoRmdBx82KB6hI8cfCV15PpYS8jV6YH3mAkbBGKR1iwb7yUr/qf9PprNgrxN
IPx3FBxalMIXaqAGkvJaQePPPYpsMmDLC0TRv+T2hC8lvmz74xSWl6LefojXTsk5
v/q01+SomOprgop6mpBxzjxsI+Xg6c0RP1PNuw7LPX9gDTHSx6qQ31bVd0u4ehyR
ZN8VPzE96+vllAsrQGdxe3vBWaPlfNNc8ZwF3tKPjhnHE1w/mNBlivTsyGUj1Jv7
2UGo0ctNfRvaJklzQ1fPvA==
`protect END_PROTECTED
