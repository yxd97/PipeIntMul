`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LvJNGG5PWgQIBXhT++V3yZHvmh0QUUS3CMxknhMdToRSYhFwl35JP8F7bna6Q6SW
inUsSxu3QvRD3o1iet9sMYchHxA6niwruuODjNQhAVnMJ7S2vUyW+EkO200CvBIH
Nejusa/AxAOyUVryR9VTM33wPsEdDd8xco6MZsbRkMQ/0BOwXD2IvVUD9B2CrY9v
xV3cSk5Zu1S2dC5ppU5ZnwI7HEm96vzoroT87cAdR135v8tGylrifjLCLI52y3ic
bsamgrM0zAfhjf8U4JQwP6M4V0lLUO0T2VrqJazIDWZrj9Ax89+EcNo6sJdxHf3w
wGA+8E1Bg0xz42vVBxWsRnhhy8z8nWkAW+7F5cNF8iKy/aVbXVsqbOCK06F0Nwi4
R+heVdI8CoXmAjJpb/gKV4ZuoCKQfGCCW8NtmBuxl0cbGLnihwQmoTD557SeWZwe
xAJ9OREkmRJ4RqlYcW8IXCWpKQJ08vLpSGdA6pvSp3hhSoq+uEYnfKZDsCF2sCbK
y0zabPts7u9xWVKi++ALkFYWo3goJaX+ibSRfVFfe5BhpnS936u8gkqlDcin7E0n
vmxWO6sYZQBkTeWqhdfYn6naw3J9JDDmTRzAv1xQCwwGSOLa4iPMQoiliaFK8F8N
slTjqaqNid821a88bv8rMWf1N6ldidPA6di0Jmr7ratiE5eWe+Sy9UYHTKtVJ14m
iq1TnJxeU5WqPo2LNN1b/MV/rylvAqCgTkjgRXovft/+VEGph4xw6KrutHkSj17k
pMOcOqpazxoQzd37dKDdQs8b8ja1QTAx7uySunmYxBobpE1LWwqQQK1uX4NOLUZI
E/RbvYmExYQ92PTBNI4RSAI5XKXSnD2+zSwRhQf20B/1dZafv6x9UxNiok0NQlvt
z+4rY6/5LBBqCxpxBjU6MeNCeSlNaNftSeZ2TcYMUHE8/2vz0du9k+m33Thjn12E
/+kZUbn4DqMO1Lon53NmvQRF2jHpimJ07XskeUxCLyH+0/k62AnU5nxCA8Nzc9c8
KgvcsNtvX7+qvHXY/ORksaDs8mSmrSyaRMF2+zS1gy06jJoefD410Wo5bYuAYTWf
cScAspAb71MuBmgpfQxwHCtF5XGVm++t2UFn0Zq8Xkzz1PvBYkJ4v8sxotGg8Mbc
wPsFxvT3G7wZFvoVYugmNWmm1UDdcpgB7IhHnxGiina2SDhDfbYWQsBzsAto4Oyd
oBAlAA79QF3rKhjuDyh8a482So37LM1+ojstdGOoznUObzpkDbDMkpCcVyTQ0pej
h6d9/sWXkwkqf7QFpjRAmZ2ZLo3KhX5lMjW9LRB8FuQuz0ny3zrtrh3XbM401gN2
Sl0p5hcvupiz5aKow0fF2lbXu4Ar/COqZvY/V/u6iDG8QvohJu3aVhzae3V/SXWE
jGv5QkKAjosSIplQMvN7lOJb6x58F6rLeE+fcHOh17o9Un0iPkXPyn2IO4f3R125
+gSis4VhsMw3TNOjd8rUmnTwq4XVeIPNDIkqe6WRrQnC7Yg68KOS7nirOgv9A2tM
MhpRwE7tPx9XETp5M+UvZjSWKoQBcJI6I53z7GKbdSdEGEXQ8DXSLwp2MBf887Va
HqglPoF2ZLry0BERFHmHbBHBK+F5dGUQXjfazX0qfPIHfutsIdSJfAxVZD9flSlW
qfcZDAIdTLN5yTM1htj9Y2LTTiU/EWXSOsrkiQOauZWeD5hXHyptuEQWfjD81Qdk
nRCg6Qwkts4XGA8q71GQoOvXVJFQ6jw+gB3YT7f3TpflyYTtRTqOWch3+R0ntLek
AXutp83hmM2kbGQZh19R1+EdyTk8Cq+NFXhRgDZ67anik4j6O9Kfrft/cIIPLfLe
3Bw7HkBDUNhS90v2h8ANFRkoqzkpc9/U7J1UggrZuTMAFqhQwTu1k3fmZgTb+HyF
GmxNfsw9uKyEOQWtf+Jj5MwAlF7CLYeAYdjaInOrw7EVfUE3Wx+YbXCrt8pQHiRk
rkyyoNZZLsuaVSwd3nkGPF69dLqgENkbFN1nGAUm2LyDgID3JqpsCGfTqikKohnz
h/CuCdYTXqSarC9hVk9hV6C6PGSrJr8WvPgNH4ROfHhJjpxGhSI4AzR62qHSlXym
oGrnlZsPw3yKIJByRZfyKTej9IYEGaCq6Mjw4Ra3S3US04XuCRYIlDA/MaPvv3Mm
y5Okc96ui7ICRzbl8vabERscAN3esuSp+P/d5snh/65iEUSg2CG8rX6+1Ed5BE/t
w+TFy4yrwJrCijG560Vg6pf+wogQaURnimZ3C9iwB7H15bzAmctK3bmd6r8qMv6d
TjgZeiLsntGLSP9D+oTEVOlV4Anj2z2QWgNjrUGBBswZUwSFZOOIAye0RFGZoUKa
bNfddVhAnU1wnkVEmIkbbgO976fN/694hx65ae9lwBslhePV7KbqWEm/vVweH07i
`protect END_PROTECTED
