`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nkX8+hAmQhqTOrr5hF4nRnqhcV6S0QCSb3aCebRSMjF05/yibCqbr7e/GcQXcNpX
aNlGSAj+gUUpV6CEOkfiLukjaOIajh9SumaEGFeofLMQ5mbToyAS6leXINiXmKF1
LiRt8St+7as6YUp8OC0/YKqz8ihOLeo7l6yegrr0WBiBM5oWg2EsgBr/rCuKtdNL
56W8HYJ93VRRO9wqkuwQpJrsCZywf6muoelPIKUSXfyOUMdgy5Z1EynMQOZfQns2
Ub8N+BT72PI+gA8DJLtMKygoV6HRsOCaK31GFRKxNYLh30J3pGXDXoOHN4zlCtzB
lcY0enbU9nNRuVcXJnU7xDd2J8CSu3/MW2AtH9ZEvlovOk0PiEgrpia9L7yl3BWX
Wlk4YEtbssbjO1FmLPipuskFRU5Z3Qm1jzUXQczXXVGILKk/lAeY++S0yr4Xt9mO
JofBXweT9SIFv8c940lb8bq+/PxC9j2zmq/Zv3bKMWWUwuPJVsetlYkmkLsXGvHw
qKZMrYhr9Lt9KFmZfTqyYwKgCniEjPO/zWmuIkAreAUabpaF74ppqFs540CF76Kd
ZtzhTZP+Oy0EC+7p37OCnzOTB844OoiZtjCHBF7TVWw=
`protect END_PROTECTED
