`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oHi6ES7kijv6ZjL8S+PxiPdSnYZxIqVmuzisxSHkhUXnwG4KscAHI/NnvDXM115I
HgdCnC+H9fJrmuXVMpgOjS9qq84u62HUMZTVJNX6AN+TG3YhLlxs1S4M+Nge7Ida
tf94DuQvMZXC5CPT1mmIWpP4bOpeT5z+mG1LJuIuTdQ6CvubWjTWOlSEb+h5FOj8
BgZ0ZTfPIzR+s8wVcg4p2QXYJ5/fzC/LeCUeLLMmBwtrAMWqRxLbZwAVMH0dqB2t
5f9MKqqhLIi2Ir2NpXkYw9q87z1oGSOiV2E/PH+gG9glRS0hCVLVjpqh04MigeT9
6axhWlHuX6yaKe69zF1zE81pAKCLWUPo5QlbAcyhCGr5rmsgLRyV0fXXkEfR7no6
Kw6l5JeVnptIksAWObGgIaI8qmyBG0VRd3EDx2N8DqwYdBgpUF7srtHNcsUul8qy
6/bzmsE8xGPB8w4tI4LfsyZGIToYPnTCHNoiSoZgaG+HG28WEo6HCBDBEgHRKwRi
`protect END_PROTECTED
