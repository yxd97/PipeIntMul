`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yI5n8Xa3d7nPZ4H8/YM1DsHIhq+MgPAf3JVLi/92RAuZr2KzA5N4z0aR/WaABVaK
A7HzyN0TPLPqGO5YyvsQhz3tzjjcfQNexUocWphSkeOmF7oRnrB3yyMlKFSE1qWz
PcFodOCHjktww6nOt6zrlllaaRu52ND1Fw2mCnSh5NeepBP0wb7Zm6lHOlGBj1a8
dfM4iDAROcqL+78gze5WnI3DTRzUKM28xEDS/3lvL+DRGP5gbCox9rlAi8o8U+bn
TmXwKQ1mor1AWl5MzrAZxSBTQeYNI7/qdbv74a+A8yAL6O8rqeeJrEfhrGe07z/s
2qKV6EKAPG8kSqvkv14oe31IIyoIW0gHTXqy4246EVaP7vb/xOuv7oTd1grDnGvF
`protect END_PROTECTED
