`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ruBO8Jjbxwp+58VrYT7ZwbqtEmLz32PdYDTQ157OxZdtWDZHfltdGijBAp8g5ir
DgvAHPlqK6CIOTh/xB3h6Gqwoa9FcnK5llmiqSTlNeHq28RvyJDUt6WVb5wbytYh
ZIcmCEdSYXJ+4ZZhRd3Aeh1bFp7FEv0NuHejanAxuMJ0B9rgtCiNzLfhXzGVo1AN
jkS45l93holDsTwiaGfYPmhY3K/rsE8jcvVPYGrDYEtPjLUU3v9vt60XOvOWZeOI
2aSUzG1XG5m2ssi9zWs8U0Sda5clLG5zH81MLwmezMTCP2Flel745rcrxxOB5qRi
I3X9X8MFRumsq2u1mOKTI0PNNLR+xfEGkmL97BzLDIwIDnGaIuJrQPtJnDd6R+Pr
8rTa9VEZM54Wh5FTKA5nBlh+2JKPRRlhbabCzdHZ6TmfPCm/3Qw0KDMVFk6dsJu7
hePihs9DryJ0ccSL/EF/AZkhLrjEELuMBDzuSIQZJDVl0aA+9Zhetpv4EJWVT6vb
CpOd2oIyR4yFbG908I0Tooc+SgRJon59ceB3y1uyn8nXihG+bjSN6qTaTD8zZX4c
vnH8QoKAFQrmMuxTjiKTuNQquRhMCDe6Gdfb13vL/+g8eJs5C6Q4xDh2VXFnhLOT
hSFkREvdeoDCLj6jE4Wttwuos2bQr3NcGV+lVWZ5dd/2SPT/KG49X/e5xwPAAJ8a
`protect END_PROTECTED
