`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
XgZa24EQ+32MqnrcN493z/+tvy3bFXaHoYVoze1lG2djv0qstYnKSYX8Vzx6Fpy7
svWSOC33KlpZmtAun7oHf2LTopMrkJyPUy5uH7JsyyiPaAft0P9/yoRYQwFj0nKL
W0voDYWL1UvD3iH7hxCEkyv2mBwFqitGpFrqVnjnRommsL5Sm/srz13GUzVbmvGa
YbJ1zqKrlZirEfT20DFEMqX5mhHY3dhzwKYuI7A8NiuTdoQP0hUNbTtMzi3PcJR1
JemDI+mxJ6pHHbU9qBcVMQ==
`protect END_PROTECTED
