`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
afgUWfPs8f116TlvmgoEwNLzXimpf5KwizYpwrxGarVUGvg9zAOTS5JRwLMq0eQ+
0wbAHtMMMGg9o7h358/DlkaIdbRQRFNeGzpZ4TcY6TKCpZ/XRbZ/gMH2o+LEQL/E
cdqXRpz8PQ4d9+Vtl1KVCme4zFNlYcEdUFbJTMukOumeAqwZgLisve9YKOguZtMR
6de6cytLxuDKNSKShYIZX4+Kt2yrObZeCOAi3BFA3Uuh6iZAtJGXiiB7imbiSBsX
dwv5quq61k8g7fXzheo3VqsdY23+LS5HeuEWAUr0yeRRxaOg16GJ0TFqD1klsZbA
K2BRInhpK0oQYA15s/uiByVAgsDWoydH38IdbcGOY+QWalJuVm9qVCwVXrQMStIK
2I5Uo2ajlqyyqLuwDbYiAkclcwUuNvvq7qjXBVBIjdjf2wv4HKBB/Q2GhWJAL1Nw
IGeWd7UXym4wo+Abckk/w81mg95nDMobNafSbaHVUtysl4ZrbqFUEdB9wKdQXf10
SxwPwQGRiCJWscTRPhTDIVIIrSHO7igiYHrdCrX4vwmqOguu3RFK0UbDTMxrGkYf
mUsq0JzRLAuI6ygPstfU2xhn0h+eGiA32I4LPaz+HnzSz0O25Vl0mRZrZm3fPSh1
HUx4k2jGhDGB1Ygn4on/0zn5mCJx9UTH9Fy4hkAFjOcH2UnyfEZf/2B9cMaFBVjQ
MviVgq9zkKforFts964tdCmQBOY7pMLWUkYKm4CiYiRWEWDwcjk3W2M0C0PbF1mF
cJ/p3Lf8IlYf/FkQSG/FWSTbSkPTRWC93CVYCiWxMc1R6lO+W/v6FCur/PRitRPU
7fwHve3mjgJ/zIUt4BeFQO+tF26KaAAvj7qG8YjtHWobjQMFjmjnM0rzhZF0OK1o
+eF5oITDC3GNrbggZuB4vveJ0dgNUKgUMiquup2cidXdcB5/LsJolwekx9x+ToD+
TItvNc+NL6cSM6hPspqCIInH0vJAVw87+hJcdmIs4Fd0HAI5YEH1Bb+d0p+ifswU
M+EPqPu388lU5Ra5UecqVCH85Y3wAgDl6ePn1DiGjaBJtLJfF89+I9Bnu4Hg8+kO
jGMcjR5riXT+C10kuWokRkWtDqk1UhndSjKpjiWT4Au8AET7c++yh2857R2mcAjG
nbtYSf+S8ETR09//M9Ksb16rNxJRW0Rkyk9Syk3y1+Ja1UUvFXN9XAsRE9U/E9+v
NqkemfbRxk+Ag6JyalJ0QwdtZD4K8VusRwyh/89/bHVvQSV9yD3jYi38vw/D3iGb
DjVg2CucmJRdUPJOe/8jXzSjv/wII+AaUa4Tc8I9hiDr6vuYwV5ujLAqlKknwue2
W2CPlT4DlPC39SZMN0WiO+u8UURVcutN+DYy8lIrbkfpiv5ks49gcpOOJ822wQ0N
Y/tO2ScM5UeJXZR3AdQlValhYikvOjMegmjoSiuKkyEa5fkH+JVr2AhTj3ctiXZy
H0jCFArsxMAe7TaXHaP7v5x3fmc0Subg5TgGU54zdw1pFhDEtYHqdM8hCmJEPBCc
HrDB/eTMwQHlu6yqmsLEIFQS56mKRfeOQyFuCI/v1mx/uAkMI9gw8/8Tj6c5Ob0f
g12mFb6+Yxsd14luu5yMRHi7e4p3AGEuMDZNIAE52LLtPlpwa8VU3d3G1DkS/SfB
/pMPMEdaZtLwa9XSfRPyqHf/vIv0tFOpdXKMHBj5z4g878LOr1vzFBWEN5YPg7YV
aJ5ObxGeYmwI5kxmVfyBGr9eQxu3kpQFfi6rrn+C+tuVxDmCV4XcPLI+f5aSNBLg
yYBvzGzqoT5ODf6jPowCFS1k4eQgdeLLG2W8V5rIwQOD73vJZGMoIGXzSzlPj9GU
GA9UYgUrVo7fH8LOmFoG3xyb7gkfJWYXleK4aptrzAVbZ2I6/1iFownywIKicX5o
BiEhA3Mynv7DWQzQLX1AbHc7STGWvTzAUijW8AJS6He0JLYQCbq6b8UBP46umtMo
XVLeuSaqWIRE6Iit19mVXxupOLUJy18cLCfb7LsovkA85zltl9wgfd1ihHEh2tJ3
4UVm2TwSfEa3BlN4nN6GqYxA0jnyKBSi42ksdPXzR2g9AszL00Z81Appvi5HV0jt
Sy4x16JEwU3p4Eg98q9AgNdFTJjUa/pRhgFyURUXFGFuSSnxux5godBFHjYDKLhC
uLm4xHC879F2Tzhphhq2MsYVIyDfK7il2SK86mnOysosZOJts4tGImfpycqdh5V8
7PxLD2+X0ZL+Zl8EvQsPmCDJga2EuEO5rDa2Uk18vdcnJnmZkSnxRHJFMpYGQwL6
5TEGPZP/8vuwukoyIfFS3Xzb42ka+wU5Rl6iB/sPhVh713fncQgtrwRQQV43gPhV
Nlut8ThN7S11CtyLSguLT35iMRytebwMQuJUpoHwRqDMZPZNstwAbGTeDtKkaEOF
k5eR7Od8aBzDpGSUeS9lUDyBgZhM6zUcD5bLWGEsrgIAblCqjo+P51xkNJVhllQy
e9LG0ru1UDg5p38FY/x8EYvSnajUzjNGR0/QNCCDyQX+xQPUCeDWjcI5q4K/Ooca
22Wff7Rp59gWWYciHbVKKlOvADrD1s8tOC6oPtBCl/j7/+hbyKPianKeQQUoA0gs
LUO+BkH8CroEALREhPxnYE4uIQ6GYQF6hk+Rg+X15YSKxH/wUef6EUtG0fibX7PA
W38StG1od6EC08o2c0wTHlJU19bLsCkc/GDcxeoqd5XUGEnFFNZkuVkltmBZqaAt
NKNLJAqcPYkT3gpy9y7ORTAetIY5DQmtn6sEISuMX1qcGC9wFKU/lYsglzS+wHuJ
bTTpqDf6LOTIokBiZWWtpZxh+q76HKHtw2qGpf1p2JiR/nRWM52BcB9NkYc20jPq
ercEmTpgjkFmkctjxnfkMN3uzaAWzErY7xykJe11wGhuaIJmN2F7lnFdNA6n3w4i
1qKKaFc5rqQQrFyXHrFCLFBUU4n3s92sKKemDFsh0Fd9CMTd4W3bA+76f6rm74Cs
EL7T5HamWXYC6qB4MQEms6mrj3mu5S/66zRmigcS69M2n/UGnktMWOZUSxk8J+fo
GZXA9K25RcM08pg8BLqdmPvdSWMdCgH/f2bwiGf9amJ7WtXcZX/LchPrB7qcN8GW
BOr6cPSCH6WBo9HrXa/TL3jdLmsnZguat5V3Pk6Qw2IduvLkdxF0f8ZuWevJUx1t
cYuE4+2Bo9dbT9b2FZ8QBqTmBhJbXDUi5efRag8cPtm+EgWBl5wHjbseKGnQLrMr
51aQkLZfrd1oPa6fqSalpp4AlMGYrSDfvgP9+6tU+G9nzrpPuyANAl/TpOKpZ8Q6
lBVvqUnf8u9xCQt3+ukIVwSQU0jQ5UK5tlg+pmPs+tDBpIXGK6Fb3ENCWPpokpvJ
oBjZMllJbOnJnuL4v2/NP9d+0FsX1U50PpMcT+6VP3vrbLeIEbkPXdhbrQs/wo0u
1EAMXKsAEQSPU6eBRSZANbeFKMg4/NROYobHoSZRc4+OTpcKPzKJxA0E0tvwJYA/
HRCULPvnsBnvaGq1qfb2Prz5c6NZgzk6heXWKEaBgbXR+Ysjhw1K90i2pyOmPGFM
bfUSBYMlrBNv/egllbOr86thxZiMHN6GA6awg2Ov1Sd13Rg/dRqD19M5xFlYhHN5
LO8vtRaXiDWJ1nQ5F9zdECJSk2jyPdnZx0BfZQMzjwlxJXRydxrvudAKkrBcszWr
1T40nkqu0tNQAll6LB/vTylWEBqCR+DGe48nYz1v7pH9bt18mwYOLhdNkXbVoTam
rzHmkFAX/aYxteIZFSF90vYFfp4uZSaWHiAKDGqb5lxjovChfGGfbGKRboVuMf+v
7jVOkExmX6NEFXF/IG2M+swyZg16s52w+wVaCP/w1EdMqboIYy/ZomCVqhTWdQ67
uTsoyH6ryVhyx5UNUXgbyygxY08k/84Hr8llgLQgVyt68YyU5qEwNba29c+6K3CG
Ul2To6blQg1HhE2/4H3RdB0QByx6iqH59y6nL+fdvebmXcq+Am2eOEF8HSZ3ZE3s
Mhr6GqIVslxp0WgaLBqYhSLA9fnNZa0PtKpTU3RogI2mpfniCtllhf4v+k05K4EG
ut0WfVrkJ/cQ/XzjxtEE+hjIUXE0ElJIGuNFo5yLNzA7EhUEvOtVMVT/vbZ/l08/
p/YdXGitnt1YRpCLywBuyZQ8eWOZ3rgWWzzX3YInn9sBCfNMFhB0rtgQKzaOuAFl
btT/z9P98MF6cRvy1L0mPLn9VJTwpKXVNoqIRdwpvy57+bRYnTR+fT9PpH2ctjb4
T1JhcaZMUsnudoBE4r0hiEtEtw5gjZVb/vr7UBgAXEMg2bR3qcRA/34GCrtPgoUY
HxsyQxDs04XXPTQqM/KxW5N85ChhGC2Ah+49UwKNznQZI/kEbHPd+CTPxbNTIOGZ
RwjwKbbOqxsawtZGadHTHwXzMjUOU9qnO4BZvKqXG0D9lRAjwleG7+OWi8D2wLrp
+r9GXxW0bep46AyTD+nWHxJYme+0F7dGPfbsC5HI3JN1INE4WSK/VcWoXFy5vbyy
X+FkhBnzl5j/tcxzhUG51Q==
`protect END_PROTECTED
