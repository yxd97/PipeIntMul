`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zzbY3cZ7H1guv2sHY3EEYfVI/6TQRvLohpBYgbrkKvxMIHTXbKTiG893kQmna8ee
/+nSJeEEkw/OTyIRpHJu/vVfrUZaAcia4dj9CoOleQg1cdEUzQ45I0EX4nofxhoT
D1Rge8NfqYnUx3BGDshXxkil0OgctDC+5IFrmUmK+/U3aRVP0cbVyeyd3IJnZLxw
8TLSJjgRpO+oAFqM7J7UqYXu1lWogqcLHlCCpWw14l9npMrKDUjHO/g1Lhv/Xqr8
C6MrOkfCYDeCQIfZf/m45oXpBprNc2NNUvNAo24b2AJ1vMHWJ/4GFHg0/bZmDtYI
/AU56Xu0kFH0ygPNRDA+nV2DCfdn1MO5SZ0qR0uqFzzKBBdBVHtYCnuIVqoDr/mE
26w+B5E8GuGjxHce4u2eBP0ZSwY+1pzV1dC++9uKRDO+PgJ4UX5EeDOc5jDVNkbR
0XAA2NVECfw4XsQv1bFjP6k3tiph91SWkhn09COtXqCUej98xgnarVN+C0axcFaq
OBmEhiG3+LaIG2O7uguyAib2dERnf2gM/5kcEJ2pITJp5Yjd/fsNrdOWhCgQkqOf
7xJ8liF1WeXAAL+5ajEkNy8mBqQaSNUAR4wW+nA7Aqstj3cMVg9xwdvtymPz4fJZ
LNFyqVNXV20W9+6utqn/NMTtO984JB3MJEskp8eo+dwxQNlE+U8HcEk6/hfe6nfc
HDkoclyETfebKA7+Rnq6/u2cqjlzYUsLaZyA510BHgbh3MwLMVckelAv6SQm1ZbM
3RYBuEqFy0f1jQ+7uFuqpTs4zRUxZP+Ffod0qtlyaeTdcZgnQ1pyDHtNBd83ztol
NBo4XYnW87aP+xXJC3xNFPTfpGN1vzmLIK1R6/JqNTD4AwN7bo5IB55yKAK5ZVAn
tL+IWtB79/65e/9Zv0WWxVEmVPTj2agAP6HhD8WwKQhEpvRGT5LUQKxhQAqrdexk
+p8pEk+5BA4a2W2+QYNdxfYiRynCqTJ6sSnA54o0NuODjueL5VxYbt6VWdhFs+dS
NYmx6J7deRxY3E6ZdzMSWwlZkCmh5TNAKCJRFzB1laNKfBrtVmD/hHHMYaCOV/Ns
voOox81y/Zx78wGMaIbr+5eZrVAiLvu+bLr+WucvUEPftRZ7uHbp3kQffjM/t0H6
J2r3t/Z5yoUlh6TIoK7OXm77wXikl49X+tHzlyK2RJKBrl4eX2vmDf7sBFxB9AUP
6c/u/TyA5AFx6e6eKWJKXugaHRnaQlTfy4OLhr7NfyMUes26tlUzzxRIestjnFNg
kmW6NjQOfr5MZjVnnuzEw8GgyQ9xTJX/SIH8GqdPr8yxecH0U32Iy2Wd/yQLsOlE
Ku0L/7mTCEaQu8zKdtK+On/M+T5uDNtvQ/5eN++8ngsTO4s1iBd2Izg6+bKwhcGB
IYcgjEOJvsDU+//NE3D/8Xw5IyR0PXrB9G+No0PSPCS91jWQJ+NJtdGq53RUkZH1
RGpknUBtgsJug2H8tWF5jmrRsCGMAihJXPCfxR4KRxdeQXXFHRhpX+wx/zVBzeFg
eK+PTqmXN17L4ZKqua83Ef+n0Ob69EG/XZpxivvPH0jhcYODlK7J4+G2YYlx/6+i
ApuWzjC+agKGqyJUE27zT5nD8bPXQoqwEZBxwgkmgJnAuETLV9JSE9WUF+D90FD7
01LeqQzkSs0+nhVIbXLZvz2QU/apBnSfmbqwmsWbyhxw2/ygRONqy0mNWvb5bCQC
FXPn1Vc8X+iiCkKyduy2YhvJPy4isSgFD9nFjMsqIMoGxzIU3Gt7kzj9YTCXVgJ3
N0oBGocpY3H3iqm774PsTetTpI7NsI3wrmmbv+wNX7q3UP5CWt+/5KGCNcTGeV2V
AgjyTuPbMN2rxAygDet4fB/ajBDgFHoMvqSejyUD8hb+5m3cpV8cKxyAB3rxwO0c
rsotoCwDqnAqwP3jQhd0IO2ihCn3joxAVx5SWBrYdTc7p9vUarqwB8EXrKK8lCMh
Smugwel4JuMoKRp+ypqw4s0eNTJhEUyQ604OcAMKy8/YthR5xOCX1ILxmXsDl5Cp
n3QprKFHKZVUDHS3F8zqrh6/d/Lt6UgQwMpdzquJnj7QWSGjrEzTUa2JPtK79jzz
Tp77ccQLBvTQMLOto2+FjfoXnkuLaLOJNOUFWPRZgyGSueP+HD51lS4LW/kYU9dE
8SR0+3FWeyO5YvzMoFmk8S1WtgbmOigEHc+qEe2idSqt9ScBYpTrB7kqSZ9VYfEh
OXrlnjToY1GZNAXEDA/tjdsJoP8S/jTtXO9kHuWFl6zc1btB/EZWS8xa/6lJJAWv
buvNb8h2T+l24PvniSZJ2oVL6wP7FQ4SxyKJx/wOhdIxiKfhLNVydz7y5B3sQXh1
88w9+geb1q5SPWP9dsyjw9mdH9sw+lFU8jofX7X89FRr2Gvj6T4L0CsdNz8bRviS
NygyTxRv5PZipP6pSjGr4SwBHXtORcgRJQQ8E4BEgLHIcZaZ93bc01VO81aN50TW
Xwbcuw8tz5CIuk5utsAqGRSsfmc3HPDTIH1yw2SMvDLB8t9F6b8n0nw/fsdTyBl1
lRH+3UexG+Sy/gfEw/sonJIq6QUTXUerdG0q/y3zfiP2ityMQWocjP5pKVXdkLBX
jgSgEFwG113nR8n40qtPs19NuuYAIrOLaoQY+hEMz5H6DHCaQHcVSRbeFS3IPKnP
ViAwDqqJ9zAKScgLWQTA2b7+Wh+YThbeWR2eIxihQQx7xNFit+SYqSEDSwrlTzkG
dSrLrFtxZScyzHUhT86SdeeIyis2RElIC5Upr8qOGXov7oVs70QGS+R6KXZno8bS
wA4fuWCsMl8a2LR2wo5wUawlqSIfERXyt4c/EdX4/9GSja3/lByC9RQKXwYkNrOU
83l1Fiz+i4E3dcaTs/z6pxLnbO/+TdoEK8064fpwRXPxGxvcsUUrkFutEpcMV949
FINyh0RUKayf+3xtgwGs0+FvHdmzhrd4hXnp6Do7lCSB9djBzGVIv0IUztGe1osp
hn1Xhtvu756aJIxdwi1+vWFeyipqT1R8mSb1w3VZ3qtZTWCrL/pMo7L/30BPk4g/
Ysj8RF2drTEgcKIWyfAy2BO+4Ii5s5TD96wl6Z4XJwSPE77wlFsr7biNLj6LJkcs
LmRD7SopBOp8Ky2FborTFsjr9OkQ/hp8XwJRF+z/srw=
`protect END_PROTECTED
