`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FN/1Z2MZYSsUV487H0snsM+MqDbJfLNOIiMhetLqIadcgKniEVIS0ycaI/nZqxbT
U+guRQ0R5YJwwyOx6tfwm4sAqzbS53lO2VSIRCXC1vzm/gOPdevP/NezpqHA+4g9
nvYZQZf0ZCoWm+35WSo2FjcTPDZU5gcGiv4L2ZKJYM/E8HIP0QJLLJ9ML/pBXisj
K6iCGUfGZuVXZSNuD/3QD7HYj8XZ/0sQ7z13w8dNzYcA6ky4R2mG6L4Lz5vdVCik
ZDyAhUPHIb5H4yAQJqtLt59myejomUmUp+QQPIeQk2/zGaKH+w9nzAmjLwTYrf9k
W56MlDbJlLZmeUlbMOYUhL5ZMgmURNwILWnbxiUKn/887IyrBXgz4mNAtVhxN7w0
p3HR5sC41wyAKI/PdnOuwBChsQAPNJrsLx76QSQXB8L4kLzFpX4BuGYqWvVI+yun
qCpNn4CSmalUsCCuWs2tPyix/5O7kjv1r94ixt1yrjFPv8wZLipPNwlhJjUC9dSq
Nr5o3zTjk/r7Bl6rrkthjA==
`protect END_PROTECTED
