`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
68JB7BcSeiSwKrTYiNV8wwdOcNfET9s4OQowH/ZMMoAV/UsUdt3/poh3ZUUfVGJC
AVoqNSB7GCySrIzleyFvVNqh09N66ob4jSH58B8tpEmzqOzgtXdkL2JLaaQDQ+qA
hktDjch32rX+mOrXWdUQ5H85PybKK7gxyCDmSV56sYh3jxNPopFuXEhX5WF2OKUG
9QgdoNX+xMJ7uNGd+lZcbZFH0v+pg0OHRQ5Kag8UT7yngcXFmNOEFeq4h1+M8+KS
GCbpt2ZR3/Pz2PUkxWXYfszgflyW9FQzhbpGn7EAhODcrKPdtGQ0MqzUAiuSG+Pr
`protect END_PROTECTED
