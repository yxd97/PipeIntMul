`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ixWeH25lvtgXXHWkHVFlaP/fMZv19sWZf3Nb8XDkWAldZPA6Py0tXikNfZaL+HJT
RmtaGd2XSx8X2BPQSLQM8HramoccUeuHcu4Dj3PG7B7K97oQFw9yi0cb6dRkZsA/
YkiWzh8F9VszwzuJKhnJPlIKE7FmWK7kjRqwMjLwH4lG6nhdlH8kkcQGEcH3FELC
CyQGLWG7wXQ2jN0i0JVG/51MJKPsiF7Ma3HCMZn3KUdOe8e+csAyGgLxYJL9ZbMP
Ad0yQyDUg9dKC5baTPnSqA==
`protect END_PROTECTED
