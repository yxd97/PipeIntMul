`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CzetMuqIlv7aPzpzU/PN27eF1D/+a81ffe+GLWtcqE5f4V+gAmDWaGjqiYzFGxGu
LiVFBTUYuGPbmPd0H53DkaBrFs1DAvKEycg4vgTpKjatKka6AWTvj2oXQ6x5qpXQ
st7ayrvbzi/0q+1J3Mb02FmMdcEgSW+4CEqDlHW6pwEVQIbbQmOdpluf8Ko3gQlC
VW2IiYwXPS5H+4aCcusOnw==
`protect END_PROTECTED
