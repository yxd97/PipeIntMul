`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CRBDOdMOP2iEI0eKXVQhg55HNM6F8f5qi99AfoeRiwveM8c/5fAA/oKO3JstiQTf
EjMNKStXGd6eB0VOdjGifGKGAaCVKpFKi2v4XimpvndXuEagiQ2K+R6qKKraZZ53
9Ki961nr3YTd/jP6LzHjjRh+iGlsBwYSI80vRmMuvFwGnAdRLcGFfTRT1CQUzqPn
9tGAAfRA77cAf/HmTJ8wh1KgKzNGPWpZFb2w4CtQz3UPLdYUmk+JzVUZ0ZF7oPKD
5M+5/QyS0MDgnpTgnJuKWRQkshQzaS85RR/ECTVM/UT0+flB3lnT7SBVhTVhjpwu
lwiw/p9M2CMWRZtySDu7pLVvxqg+Fm1YEtafZblJ8ASCM0mKDa9neIqBYn4A7ZyM
5s3Yv8QAOE7t+nXyNjScC+mKVReX/VIjqn4OFAf4KfS7XE6QDdmeiN566H8cyBW2
quMCfWGCETwQ5nIPrhVTTGjWW9MFolgbsYuVlhnLCd/AKwHoqfHGV387A1vJriDG
mkm6wAjwDohUdj4hqBY9Qr2mNvUA78BcICNcgEbrHbxUY+E7K6AOTm57N8chyoEm
6rkFqiSAuKkkTdte3c81SGiV5RYkJZvQoaH8J6GDAMoper7KmAbHIZvun8IlihSM
u/NdYylOiTcIpLAmjriXJI5yD3YlgBSOy7qIg0EvMgaTfR0OQTR3H0bQXEKPWzRY
aBq2iNOBTKSGsQUYNG3FcFVDE+xsGKNRhCYpyTQolUJXIxIfODCx03rfCHwoUfLD
/yURdPiU0hprUz/kHRM9pP8g9dL7jyXacgu9+QnmZt9RvC+A2jvA2VFwytwIziWf
qn0TI1Z5pg860h2FS80OljN1+w1Jami1ZB5fiGvpKO03B40iPhhTi299xblY2+ek
aTUu3EnEnXnF4GF2reEVBt8gjX3NXJPAKLbhWy4mtWcBTpC3ZLPQc7am/rrhfDUa
dI+G8MEhYg+8WcTLu4ma/X9duQfrMJnRUcPjJpYs5DJVCr9cSDA2xh3Eo6dbMPkV
V4i1mxqWrUz3lJlZtMnuywhyvJod0ZAAQKaAHMBF+cd6TJ/nZPttSBUDI0MOXaL8
E7aGtkoVffMS+WQRhkR5I94xDi7YaAJ5eSXCfwIQStvTP9qrb9GNiEfwDB6mGL61
3r9BOw+isJZMswe8UtV3jETvynb6v6v7g4sRW0rdHVvFj4Tn/JVEI7taHYUxIpIp
MleEV/xUaB4o54uIxSZhHB51BlmTucJXhP/CTWTfAItH/xtXtQJ250QJ1DrKiJaP
3lagxsheOOw423xkOsaOhjQSf5jqwCOI3yb25V9/tb5qbKpy1MxQ2HFqyx/3pgTN
`protect END_PROTECTED
