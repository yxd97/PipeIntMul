`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VR5ZEd1pWnGZHPJtuKlVhajFRUWAsZMAVe/4lDPLQhNjN0OTROGh0Ex/D/dW51J+
FstMfk+Rzn97q/bQiYSbAE8GH8yTcve8vj8+7lE3W/JMJXxTfckQI214/Egyo1sR
bGNHU7F2ukMJuBUeuZqzGk7DOtbsiwE0kaCD6GZ/8/WQKAdGqNjRnjHoRQd7XKsv
SR3a9zToUZQvIoOWHbMtkt9j0V8OPxhVOpb2LZSvDF3P2HzWxKG3pxAsZS7hsK7A
PyTwlgcYNCFJ2GxpBV2oZ/bkHCt3rrmQaU/cSRNyzmbOwVPvEmrUxsQ75RzH9VWu
K2l+7ggX4uhoWc6m584KJhy8yG6rmZYxDdnzLc/5kyQnoRrLhwM/cY8/J41OTW42
HnL20JyDBX5Tufegove/mVKVVgAD8+nX8k+MkmtWEzaUOvyrk0xBWcE5TPvFcntZ
3Mt/DBTvNlnYAeOnt3ma3Z252rU7hcnhUIpEw9/1K4VOieIL7iGew9oRVzFi1GCe
kAkFkD5errjmwtlU6yxPV4OClWweceUqN9O9VrAZlpdhBeFGdoSnDhcrKm0BUjPW
PQCoEf3jel4JhMkO7VIKmJLcDOMtHGIqOS5xHySBAbnfsoasqmZF88HyNO2sB0bT
jZVFcHVW780JOIJ50aF/EPN2Y13aPz4kgPPeds4hQUmvzfZ0TcYQMv4liRSUIjUw
f8/3jL3iMAyxrhXq1gv8OV5QeWDXOktQ8oBjEVuVWXx2Mil3yE0GTuwy2nIT6HsC
Jg935dWdfjnlf3gGEsBWNhYsedcZo6LdzXelpj0AhtII9O17UPOriXVgqUt29Hmc
gz5C64ta6xWoHr5TTNgeRp/WSuLh9/H+m37MjrBhiHZlUJaPBjdb27EV1VwLsJDD
cYoTdWzxO+HU5QJdg7z5tA4PoyEfYuwuAvy8XKIpE1+oqCx49vH3pxx/o4lJlZxp
8Mh9N5l3BOOdXNC1dO1a8RYH3VCbgSqYLFG/s5tHKKqAanJgRYI9W4AXF8FcGRWk
QhcSyX6sz3nILvf5u70Fp44HKQxYnKTZR+DnC/Pms1HJqldUZq7KGbny7Uh+RqgY
ZOfi2De+yWzwrnB+8TAWZkjPYo0rACewTcd1OoF2p6Q5Wn4Gm+TN1lR1eQq5ZMFh
9LpApHQrGbTjxahPySh7C5ueUFcE/7m6OftR/LoiiIM6GE7bxnVWKdVwppHQf906
H+n0UtPJV5Hzga+Y2ukEryiE9r61q0yNxgvHgkmIOtLVHY1SQv02aCZ9wV0L4mM4
YjmV+m9s3JrgwIWBDvH9t3lBK+uu8qc+3YvsjFlSUHznClm0l43Uh5eNoZ95swYI
GzmklvKopF8O5/A95Vhz3nYHIrITtj1RaI6+SoXahquhmt37ZcZ2O91MzWfvEa84
yBhY7g5BbeLzpBSUPoPHs08OW6FKl/5o4UZMCJ4JEwPawB1LBu+pK6G0pxJ25Ccz
gA+AZsm6unMEgdkkAD5LIhbVpbFnEmrwA1p3J5m1KhfAj1bVxEEUNVXRQ+Da4pcW
9z9+f3dmw7MGwR+CwIrqEj1ERb4GyUKguHy6RsCfsoaQUAD43Q2h9D0bludN7SEo
q4SpPiHDC2y63ZQt7WbZk/gloRU1uF74zEddl4vatxTzdHc/Sl+opJncOWtnBMWk
iAtG5CGB0mFhfw7LdoFH1StyjXSY7jxPz8ZUsnkVFnUjTwDs92ZT6tt+L6nG0USi
5E1oHvcc+r4fBmor/lCkY3ULXlQEFgTM3ImD+tUxCO7nFzdN+I0asy3/kS021Cp0
0VR48Ig54NRHtRyQc11LcXCfj0d9Dh3dRIDbVYenHzjwvtn26xd2LBy1LbazIDjW
iZCL7z14rLEJ8DpKSMJSMNM8aA0prLMX4XxMa+ag5kRRYzG7rm1CibJj/MX5+9WA
66P5uYbGZ3LzTJH1/n0mAmFZSIhXApTjCYsoDf0wu2e6TgOX5VJF2WVvtkTQ3a3W
mcknZinSflQeDNVudg0k2v2Yb8LTSe9hnE4+mKid1LkO2HmQHQF7GxpFtAZWcPtH
ZPRSDKQ/zvT0pemBgPAN1WwO3orXMuS/EQbTHsjdFqByRDrPRmy6TF4B+fx2Xdkk
JkWbxhg2AHSLDklNB9b8oQ==
`protect END_PROTECTED
