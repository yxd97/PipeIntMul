`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2j4nbIFMzHY3mcyIBOabVZunaZgf3FV0Klg3Lwi95YU14VfqECGSqIf1mencyOIn
dnERpiWrO2Z9i6tD9l2pKt1Hece3jwwBfDy36KQtjDdcbXVOnzXHIptrxBaZfEBO
qFXFepdPoepQgDXVKf+9kOpGZPO/mPgkDgRUhAFp8EQNZiNZsVPjf87ulL/mgw5V
9TV48TA7s1xw1fNiGNVtWrucpoK8oid60iMELkykUJBhmEGx7nAnHul/rfcQXh1n
L0brthisp5H2mWppnsgx7hzrvNY4zdfuX8nI+E//d37zIbEn1M45VrM/ZVsxzI0f
ZOIeQUr1eFw/qNGnzq8P4MhpiTkSiSe/1Tp8QuDhCsgaRZhV8IhKeV2SiKBWVgOU
4b1YN7ki4ydMFW2WTwknnAYaqek7V+pkkIujWDmQYKA=
`protect END_PROTECTED
