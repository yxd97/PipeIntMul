`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3AjdqQIJeWpUtXtTARSMaI6RGIllE6fEZb6G8mjsYztP1fsFEgqMd5jYfa+DpfbI
YSe7UR3XAUeSBgsNFagoWzOplEg2rzPELCuhnT/MGFu5YGD8lCuW0GfVPJny8dym
76QpeX83gBJwRaSb/qStZhGq4QIlCtAVrMtU/b/9bOPag1WPKcBxCd8qMTRCGTWo
Gqbp9tCTMJcjRynITaPh9M9MVG8kF6m5PJFz1PviK4IsvW2CucukvAt/L3eoZdYn
rRRtGvYEMeYcJJvLDueHtP6y7kuGbQQZoR0y/0Scgm8WfF5hNh5QO8qWmtcQ6iQG
5l2bEl++pz8q2u+FLwj1kZ6yTabuLgk1BlQrp4AU1lf+vjqDtCeXKgP91zEuDlEE
tz7fRNdUI2yth/c0VUlLzRl7Eh+6CmL5o/T8qgLyVd7j2WNnr1MHf/KW+tl4XdpK
ZBS4vWnfEl/xDOnggx+UfwV+rElgYiWaAaeOiH5dayQaJ2ze/yv1jsbbsYPGc9uX
sSbf4KrUo1zIFyBIWjGT9yO+J27a1ARxsG21KFMtY0yB25nVnUyxBJz7rigtDz72
GjH/ILfggQRpmSpC/wIBH97MZccORQ4B2Tx66INrjufuZtYzEJCfLdN177SuSViN
aBm/giC2qwy8ke4URCtn0KmxjimfMGimwQAevXHpqGwV+aM9nAbJgc7l7QYIxO/G
TFhgiVYkqiDERxKnq9Ug9EvmhY+SDF6QABxfnrScUIBLZiNPBoUJnlsISxTX0Q8I
lylDI8+motyndliac+hBl46198wNPkfw8/bGbCcZIUa/eN7KlQ1idsmdeILn+VZe
c+zBD+bAcj8MgJvvUdXBapgxBBCfJX7XvPspL4wj1NcAQYfsSwyurr6XAMxaohoN
usjL77yC4pZEzyxZBCjifebWdW2vSkYkpv5IotZCYwZoOVw+njFz0gYtuF/vrbFl
`protect END_PROTECTED
