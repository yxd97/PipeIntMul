`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
56CVMxAL9DCMOJ4zHYL0oGxx1nDYExNvPEYfCleAwmOSLnYTZAyChOGnrypjPM+f
F7Mx5Hbe1VIZNWBlSFLckQVqgoazNuTn/r3vIJMTgxLBbdIV6a8biFARnX5penjh
3OD9idDeoLgPsSVXMSckrhQus/hfBsyL513LIaRZjwBK7TqdM7rvS8p0GcH8llZ1
dzvttbG2zSNKWhTwLUAYMjhthrWvyfDnBXNlWjJvg0cGXbj97cLijzbUMJDCKRXU
FzUwYaSy2Nk1ryoYHzwKvMQCrM+IqNMncE8A9tPnA3kh7Zv4YCfStbX5rlJamik/
isT2Owgrd/10JgUWP95uEsEPM96oQzhF7weIEVf80Ud+2HmymOl5k8xw6YpwHP1/
puRIRwYRd+KuluyQwW5WwXJV6bOBu2/vLy9wH98xXfCvh0eKbl4SqbxrzfwKPk5C
+hMGW/Lv7McE2+1r7SGEyCUhxXDxGMZJbwuBaeV97Kb0pr3ophrZdtw/YHwHcd0u
XWWOHi/UDsqcU4Z7fLK/M2Npt4Ay45vsQHkQ2/q8EqN5EnzabG93LUhwoxm0ha+K
w33EUFfIhTmZqGpQv5NCWdrq3WgaV1/0tlfBd59htr6bfnd68Dd8nkBe04Yijnt4
JLg2rHvQsvBE3cvvD//Y1na5ptVNnQ0zIy38AtVCPXoH+9ZygOMP4Tiu0M0wBe60
qO/oKyPNVjsPxcAFYr/4dUa/EPxyCW9MnouVl4MQnRllDZ3ZWTXjx0ADsdDv+Oa5
Pjg3t5muI7DJ0D2c+yet7P0SB4j58U3d1s6ST+R5zilXgSRHxlQsPjrLlsgZZxD7
WRHS20h+Ie4yVgbVwPfjpWD4rk05lbmly49OFgcw5cxX0EpDeJGeywFAMf8wEuQZ
Nj+pK/eFMEfPq/bsiFz5CLvJmwLaLi1oJetTWQlTO7FO/GyeHZIdWd71Qw18rCXy
NtGX0+4+8i80z2f7Wl1d6ICDcJedfPQwl7/+jO2p/ykHmTv/8e9Hy0nGvEhfVTho
ba23pybQ/GydJq2hJTn1TA==
`protect END_PROTECTED
