`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mDZsIXBo1JKsB+EERd7AdLQ91NmLlxwfEFsuALH6LJF/ZwvaIGqHtAyO9MgesFJx
w/AziLbgbutplBKQeMxmiYAgKmEJtXqtmfugpECXwHK2EuvanQmSUK1FImxuU84g
YaR4iec4iZ9aum6/v9pav+HNpybYhv/pnA36G/JuVkXnOEvZsMgeJ//rqLaczBP3
lqzltmuuSSJkBiuzEIKMdJV+P4yf8Eocib6t2gXAFPKyOLasDZ19JYHqfKMH2SnH
YQJ8ZJpuWMzTgH7mlH/L03+h4CdIQrsOxJ601WmKaCHYIOQ8whu0E8dfIiB3K9VL
A4wKYI9JGFr8aTnPXJK39ZAJfNr8nloin9mI9ZGXQVzXsQQX11u7flqnVqJ2Wqdz
Q1LBQrSlXCE/RPWgM4o/YQyKDHazGaZbergvRMUBOK4e87s/f2RkPnsofwg8cFxM
rRHvNgk/VSTWR+ixgVctxb9JLPYxRx4zdH5WdXVJ1KhSuKWcu+OM+n9PteUdI654
`protect END_PROTECTED
