`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gpXQrW6oNaPyn2u0fhthSNzYmVmp+3IRg9hDaoBoh32u3n3OPqPCCd5T0Ub+xb5G
LcOK0s3yEQrEiiZ2FvMBgw/RuOS31vWMw5eOZ8aw3osQMn8H52++4r6MWkdzvynH
oSnS+5ZTOe657u80EMLg/3dqy9gBL1iXuj2qcTRt6WFdvbpmhbYi4qLQDdY3SbU2
9R93N4duJ9xncLpdo0GIrZ4dp2j/Ds39oVY5FMHU0rItfM0RxqGMKya9iVBfucdq
s5ct4w/qsperIZ4lk0nvvtiBFUe9UJv0MIkFLiHOIWz9FAtOXy5Ezz3ptIMECQxa
30PLMuxjEebcyuXmt91g/Q==
`protect END_PROTECTED
