`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4ZCiWkw9f4GGX2qs4d8UZOTtL8KTRiSAsnsURfNBHG3sYvRcxiS9BUavv4wcO07A
I5yJwXLm8R+zew7jbIMeyWfrGWx6ROE1KgPveoNbTvAGy8592iKtwgHrV4Ubb3a0
jZGRBYzLnjzjbiWo7kfrqqK0jO7tzHGmjWeFpgwNFslQJl/TSuSlEXkEKTAVdHpW
5jYiPfSSQJ/GHCbbxQT2nseJIN4GdqW2y+UrvYNDpcZXkBKBmoxBicsjO7wBwlSC
SfCmrNfMYckbBq8HglQso4C77a3nsmLzQDq7h1pSmnt+TE+rD8E5E2nQl5qUAGRL
4pH6Nfpqna32ceGIuG8MDnMSzmx40YnltSJmvvTBYuIKgksv5ev3HlCJnZmi5XIa
OV/NWkG5bOvLHrp8GK9FKHe+YEmlc+Yy4aGuOuyxv+L4A+1G52YONQU+oXBU+ban
nLKQX7lX1VtNLA8ElKfPy8ferZxYV8L3w18YxzIO5ZE6i2Z/l+SOAly1T3sZ+g2O
BSQu3KxSmw6NGl7VAirLUxdpdvfmIIG5EY+IW5PlvpPTfh1GVIgBti/uu7ugDZSt
uMXAB6J71UbORjwI7TALMEulG0hexUzxU/50EoiwXj0WDKav8pflIkfouqPdYWvj
Bgab3tPtlHS8HLOzy9cGZUt6MAlZAo8oT6jdpKxm0Wjbu80Mn+zSQhlKHw19GVNR
lLA5rT9QEgHb/7Vbkdp5VE6WLWVWBeOy7B5Gg1yZOT0BbIqThAVtH093xul/26Ek
mH+uASCX8S971GPevJHhqbD9Prr4IVXn/k1pjH4bIiHeij5aYDhRoAv+bsPttp3O
7nfa0+57CVwWuy4KG2FvZt58OeP7GC+X8AwaZ04T7yN/9pK6Sidk/lEcYm4wm03Y
FYCQquXkTkHauq40E9IHP6/fsVWFg1LEoqgoF/VmxpEQ+oPQfIulvFtfyuXtKUQ3
d2VTpTiAQ2Uo2lAc4CeIE5tE1hIPggZyhGUJUBDTa4S+mXi6Xe74VF0L896+5m7t
1q7sOhQv8QVC4NHd3sGy4OQRgklg3Qh42CoXYU/su+N/w1b5Uyg8PYliUXBuc5W9
r2xnPHto/KBEn7vUq6gM0/AV30rGsHvCv85DKNbmpBBr6mCn8IG5IdBWlOTrudqb
qtocwqz3gIWESOqlnwFycDTfEAzl6aaLkK26651gzUMoCGCIBvg/5HWSCsJFxRvh
ap6iPbh3Tewqkfs0/cDIbuffbfbSpuE9jG+HTJlRvsGgTVP6BZIDaV/JloQwjZsu
mRvSLeH0lV/RcWtAits8j+FARomi6ua4thT9c852rqAYrKV9QpYpWvyN85nNc4MU
kn7mo2aEBGqy9Jofabi5wOZLYHLX3zwq3gKfc8oSfCYkjmh68P4N3Jnfcr0UJPuF
`protect END_PROTECTED
