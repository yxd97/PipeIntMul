`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9iTJKK+tnRBVAIPgCN4KO0XxVU7qwuOUrcXIut25/6OF4p4tiMWicYvs5mfN63BH
CKc/l92gOkuKJbylJ/k6DiDx0uZQXiCrMawcUFJJIctU1FrGnI3NrR0Yw+6lZfER
4ZUagNQ8gc1kdJ71gVm9xLepQo6IX4Gm4xFwLq6HlP0Ok4gxrmxqM4x2C0UOwiBl
3Ky7TLg/9aBCFPcmFiMaXBVB1eqZr5M7azkN4sNvUMT6MYBqnodF2LqO4KPp5uBm
qnUaZW3xf4B5VF6MJwRkziSjSi01SCMDPuYc+6WrPbqyJAzGlMB5PlQrq4DRgDt6
IoTqKN1C8fqifO1E1OArxSnGyCVCvYNvz4HDgk9/m6T9sjvdUYVGqiBMDyKBz4wO
bVXIRLgxHy6mRuUNxwpwtukeJAH9FIfhpvlzxAwkRaYovows6SRxc5NL/bzBP4In
KqcM+qBR5VdZaBYyOfKCXbU86A2uAloQaFEHp6bo4/KQuK2QyT65n6OJFHZFRjo4
WEKbguUlVl8EVN+hk1zmKuutjQvVmzyXH1OpfwMju00wa0MODssqE8/wA3svHkvz
GgLK+id3uG8psI/XOo9qFldgl7YtVab+WyKTjy5STKgEVrZe5YnsdJYgJbX2hlVc
OFZ0eEvneaaA+vh4XiyP8R9mHns6vQ32+tBn2x9Zvm4+D/SQL5lkvQjMwTqa/IHQ
XLteceOP/JnAB+aj475iVk9PF6RwlVWScZbpXzK6BYklAF8xLqh25P+hTbeVMR7B
cxo2sqNaiQ/ctmBlyJOuDLzzrcGtPw/OHLgC7Wuwyhv25yNRc/Gq+xVa/ZPZJ+w8
I6LndKe+2s+ePVLWDIw52KdHxFd8aplulhXly7dOvBM=
`protect END_PROTECTED
