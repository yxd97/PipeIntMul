`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
sjLOorM4OZUotS6Otd0pKyI5KGIjCkrRp28EAEqcWmdErxmgl1lCgtg6Xijpe2FL
u2ft2QP8Uj3Zk/vReAEGC1m3kDMvAIU3xbZA8cAlI0TahXE10Z7UGxhGlyjUK7cK
s3fqZoshOgEt3zZTjjX+URrpSPIemT3VqVNkvCT5kGAbmIdRg2OdZ2mSBlNdWGNF
0BzMC+1NJxfVoJ8beGqnnMqnCl/H/jaExeTWtI8gG7QBRzw4Rrfcwj/ASbtjqrYG
QIwMVOQeqTNjhjgaqG69cw==
`protect END_PROTECTED
