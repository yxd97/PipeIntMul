`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tcz8xYSQRPb9gfmwVGalZxdkm+02CgoUPvzhRMw6ZOew3VzuAPR0nowAzXgAiLiK
0DMYMbySFh3pAS0Xw+9Gxgx9b5b1qjhUoF6J3jI3qLKr8FL9v0rW54EGbeggREmx
dNvskQUWH/zWZHs7U95spH2fjxLsQSZyPpYaWBLvyLYrqamVFKOZHt1U8KOlrcHX
EaGFFK0C2ffHmPuGyAggbcyR0tVXcix9XSHhqOGhzNZCIYHeZd8Tir/sd/Zk3HCN
7D+EUUn7hGcigMorRcNrQBu5S3vxvsXl1lGqLZCzuP81cezqh+RNRiwbCbc/N/06
`protect END_PROTECTED
