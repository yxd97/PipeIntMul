`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L5wp7N1HUHzvNrYuFEYj9Sxl0CpROwm+7X/Rzlj6xogX5ZH+2fUqh5/qMYSf2lPE
cbgiSz/HWFDIHEtkO+ziYy1WmOJ/0tjUtkFRbg34WuqDxKo7oFlyqxR1KFBmVhAv
ppD4bYKHyb1PYwk7/hL3sx6/G/n23rGjS3DBKQ5BTqvH+yAF4vTfdeCcP8S+sByZ
KvyZ+k/BYn0J8XWEyWtVPeCIXPIyLpxbLP3jyjPKczC57iiKFuUCBJDwP/NZlNnd
IfBOIn3RY/7zTFr+r+in3FkDZ7rJg1jgGncVt4+4CjBP0iOf7pw1zSbuEi7uOSmz
mvsNQvfeIDMWhXdau3ztb3jDjlLq3OH515J72t3u4AmgU1wbLjCn5v4xRp9idZxB
Pw2XeQgZ9VhXTskyV78bSjaX0n7/OBt4ACZ60vMOl3RNasU0btluxtr6AMVkASZW
rze0nlzgyjYIvpo9GqUUpMRrIH/O1jjXxL6zgRxXsLa7kYnYx1zOD1wZQe6ueTAb
qSUgObas5Fr4PWtZdSOsoODqfJGuI97kVg2HCd34tTjw+w/IzkoCiGUvgEejWhaD
7H360PofwS7GFpTChAn6iCuPjUyJ8yksCUebb49A5DJodrmZIcugNAPNgIevkbsc
vpSiZZIFKY1NCuVs0EqkyYiusGV0sUf+Wkt00rSuwD1bpl0tdWMyBhoVCuoArED2
DkhPghN2LNkxFCt/Cb9BP4RxbHKp+2uysfzF942G5U8=
`protect END_PROTECTED
