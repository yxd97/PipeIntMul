`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
61U3BEu8m35VaddIx6ndPEbvnrrIej7VSMVaxNyh82WU+y4x8a120Fh/mTmkkwmm
zcisfAkn59babCtZZtswiiDvsOyIt7C4NGS/xahU1mpUY8ePLb7CTNlMepoO2Iwc
37UavBh8hT5dOo+uFmC6nQ+uaYI/bsMhFIpcjySpGlaAuq21/HaVyj+VeIasbLRS
kqnoQ0UdA6337l9Zy1BVRYu24NW0PiW+kphc7EzaGW9gAMUHc/iztFGenpnQN316
JCKY5P0ci6yrvAS3EqNI4yGx9HmwMMqV3TDniV8ZjQkKnLqI+LWtKB4Mo4iqRdDe
4e/BsrSrFGxNNnvL6BEVljSUfrn8JRvS+U2LpOPHWskxFyAfkdxmyf0Ele+SA8e0
TItBJUHI1+v072S7v2wCQ2A6cUryQY6MhrqN2vtNsS4rdVSwxSgOett5jOuXJpTE
Ep9XaRnzkSwl0+0LhTGczw==
`protect END_PROTECTED
