`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1QbFTJzd9tjf85y/qQxkCIz7QBjd3EfnXJh2X294yd/C/xfaAhsmszwEH7a/AePB
yrb+2+AXiv68IefGkqDvyhi4Sx/UtCAIeMZRO+IQcQJDhS5xF9bJuy/I7b6dPohZ
RuH1wXXGjFVElPcLUNZPH0hRNMp682cecVkx0uIhn4Oxe/oRzZ827M1gsviWFwu2
ZAB+O/fKcEa68n6Ht+Y5lAsZYBt9vCOjZPBYT4VWuchmT97cRaPbxaELdS8arV+d
mZ5TcSFdHfUgN7Ob87i4fKsDGunxuwJmuam0Vqd2k3zb9Wp2PpjY8boWf1RgU487
eZ9S38L0Dgt1ccyEV6ZnJQGm4jIQPWuPZuSD96iKEL0FeyidRuZvXXvpOLq4jvP0
80ErmXqq8mQGLfq9039wPsjoVOr690sSZwW+mByA8LJsZLxuzaL9+RwOGnUfgIXd
`protect END_PROTECTED
