`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TMsESQQ38D5QGZxIHCCifengkAiNO9srftQM4VZsj6CxIwVPZekw/+R21VBiTUju
WmTF7YJAEPh13pltKwVY39Axo/+m9wzUhZt36R8Tr4kSP1VUt2DqAsmlagsjX/ER
psRxa/FdrmwYVMfh2NYVwWmeXyIEUezVH6SmEvQHB8GzD8sFV00nqK4SatZB8E3F
mS4Ajfwl6LYNhAK7Ema2JyTl0lIA1X0DP7YiX99yN5IJXkU11SxrNs4ox+N+mS0S
a0TqAEbX5fuF1IbhpFxrWvcIrSkDSwaOjhne/mr7iLe2mGz/xQgK3m8hr+nyjrUG
nkrQ1j3gbexUhSon+bsNpzAeESilsHO5GnC0yWomWB4cKiKGs+YGSN3Pi28PpFSJ
8WEXNjVJFwMFE73Rz6D2VbfwpqlVjEXSdBe6DSFl+RgjR81gzB7ByoeOe1GR9HaQ
`protect END_PROTECTED
