`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cBKotcdWxl+Sevpu1nnP3m8X/9qB7i92DsVJK8JPA0rZCRdf2tNi9QcHV0enlsPm
8s7FIE0hhwLrHFnJhaocAmgb+5gDEwpSZ8PQhw05+6XqDnVhHkWGOfPZGukRcxFi
9CAqjQzjTDyCKXCe1qZw4NoEW4MazckHHHN/8TOeQ+nycVBZHOGvWSVqepRsequy
hVEEpLtWWwxdMf42Uo5ihUSpOQBllK0GU/FCstMhkBosXvSto8kroOHyu5KyOg+O
v53deoKNJArd2t6hpoDCZOjC7uPKj3/bXJdgE/0XlNXVeuup695bsQJBfjn6kbCc
zWRAE6ZjmFLDa41aaC6dgQ==
`protect END_PROTECTED
