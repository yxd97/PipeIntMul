`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dahr0kKKrWzLkt0iaazq0i2lkPWnLA5Li1TZ1EjM10YuYYjHttsHfO2HV1H4GKhm
mVBj2SgmV9RpI6fZL8d2/fMKQhGYD4SDKG83j04aKrUgOJ/8fVp2f7bcyxjpGzQS
l38ZLa3I3a5MFZprMSO64a++9aoqlZGNKeNR4+yhSbw1sovQBUMLOpWZJ8wEnq1A
548/NOgx9QIWQBwZm21JF7vsUxAo48fYNCOKA+A5hfIaiSiYekUhdRCzT+ILC0pm
+O+c3aOl9ijd6GwvqPNGVMenO+szfQUPQybyq8+TXq+N+vVNgm2LsVRaGgl08n2o
uwx4fz8ABECpk19diqzIe6XajbnyBiKcJwacqdT7AXToCD2/CV08ngFnQsjTzDAr
`protect END_PROTECTED
