`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Xa9QhKDGK0bQauLCtLwbD7DPcj14HHoydEpZhkrH7TyJF9u0GtX+XazeUvScey6S
6tg1FAMjoxcszqznN/DPe/3EINnOSeyoH/mKmktUgL40xqrm3J7frlTbDkAyKXQn
ZauimYfYPVDp2RxhJWkm/KKIE3hvgW9QKAOVDgkktOyLQJRkG57YpfPfCBR5YSvn
Ah53GSUKEgXkdXlm4dQWoyfqC6Gd6mtfdHHfOn44G73OJ7e94WAEC6iN3pUZKM4g
PDE1gPccTx271wU4Yu+LMTWP4x4a/FZqCtvs3a3/3QeNNc/ftTlpDGNwPtworcH/
CpP6RIvZPvUuWxwB/vS7UOLxHUJD5kqDE8h+RLAn4jVyUjyFqz3xDQYrML14TzEV
L3PEOblVbF8rZ2FusRrV66v1379foIHNiTwiRuZxREHc3mBIapzZOHOG3sv1xkXQ
AT8pQHoWopxF/lGJ7fGcvBIwG23reOz6fKSCduisDkU=
`protect END_PROTECTED
