`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IJc/7i4QJKESryNexuceJmCIOiFxYJyuf38AVKQn/sbTs2Ojm58N+3n1/5HSV21U
kR5/SnJGAViRPBWJrUT7g8hpvqufyxxxw0HnxWVs3Jje4rATcuV8MgR2k8sgcayk
9SD/DO78K73BDL9XvM97OJPdFdB3EQ1Qtwj2i2vRM7RwDvviuXrThbdAhHhaLQNr
Aa395xVw8kz/mVHBIzK6ufPYTKTWP0OiJGhQCAzIy+nyCHywjMwA4iibv+bxywAU
QvmMlMIdjFX3CHxu+MM614q0QsCX8bspeJlBF7EDAlOGRihnqvdLBsDPAeTTmbxE
mqbcD+lyEcjsY6/SF7TceEBkaUYcFRHRvlkXiCG4LL6FYdUD8JPWRWN5yCoO41cg
mcZxuV/vxkuPJT9eyZBpEyKjCz0j9ybaKCPCqJmEAPoSh7BGC+iwBqD+DBgmae4N
Ejyaz2zaFy9jMQoHzeBcLm/BSz14FFz6QfuQJkaMz9t1sbk/T9g/cSydqqoDGO/e
OcTRbnvSsP5ZoN5jUMX5zdCoAvpwgp/S29UFzgNOCaCEIzTvk9cl0XtTp7AqaIS5
FQYdjx761RubVn2viGvMqQH86pBW884zWJpbQyLT21x/B/cwFghsr+fpxVF4pXpl
PlskXRLf/RIAjSMGKywgbg==
`protect END_PROTECTED
