`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iQ1VUegODVDHoN3e2jHKUs3sAILJjJuQZtJNQCi/cpm5scIAK4lOwFy04L5t4MOB
DMmUPZBbk35DvpGHzLLDSG8xwGDQyRHlFSfYyiJug3y2keL+m23Dl2OD6wiJbB0D
0TXFr8K/P8n7B0T5Vrv857r/Ngr1Mv5fh0NB+mpO5AArVB/Hwec2f7kCN0hgxasu
qm1oZujziYgOtFaB63jUbkTjGEw/GAmZuZPlyHQSUFhUhSdyK2KO9N86mmLMXwNk
QvkS/+yOMdV6e8sLiNiiy58R2rLlHkg7o6P4iQvOgUK+n3zI2tRKvYc7KvfG7g7A
EYaoqjfsblGIXOK7luNuiNbLfD1qHZcobOWLLSQNGEUYCOmEt8eGDMDcO1G7HnW0
0PMU8qCdJgFrEyNdLZsTSlbCvcrziFOqnjYoUD1+PgVwHyzA14RIuGstYl1QLNYd
`protect END_PROTECTED
