`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cUvC3WraHQ7E2cZ21yAd4DNUh2cN1FhmuLnL44tAwSmpwZIENv1c9ESb9GcarkRQ
QURM41XHgSZoPWqaPS/p/w0DrytAalMywsK9A0Qbmqfl3PjC/67JLPxvMsszHMyW
YgvoNnyaGGIFBXSx/DZwvc+KiYsQ1wyXkB8OBLEMfdJBt1S9GIeGoof5qgrJbn6g
a6O2y5qbIV9bhsdocfvCxP7HYRRgSXUl+9UCaeALlJoSiCDjaCpmm+JzJ1feK2Ha
5f5C5YDXq8IDu2JF/cEUo0ofXbc5R9Fe7IVNIdX2b1kC5nHTZahNWwgoJ5pPKx4i
XPTV0DD4ZmftFlt14Tte9i/stWAJph+tFnn+JpajBULiE1w7rPDaN4uZ2pr5HVKV
`protect END_PROTECTED
