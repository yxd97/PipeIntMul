`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+b4SR9D9Z1w8o0HqEPgcDleyRmk4HRFBwuDao/yoEZHp8ap33zj2LknnU/YGPtZ0
k17Atmlsedzg2NZDQglFAfYuuTL+ZvG5KmvglQCBBK/NDi3G8en3yDwQcB/mxpWy
LmpIwHL4t+r6fUock2tzJgxAjeKSgi5XepyKgSbRI0lGoTM5oFVGpu4rPXT0g2FW
cG6J7hY8EhzJtn1WH785IUC2aUpjbeInJUZF6ijd8MEAojZWDYRNH0Cj3lbCDF85
TMHZc0SiENyYw+pfpt7P8Q==
`protect END_PROTECTED
