`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yqVqTSghCylYGSpiit0P+UixRSKo7rhKgdNkQtFJzUpApripXWKGt9PF+0TpeQBg
Pf0MTT0FiNj74LjnSjSa+IhwWEqcDrufZ+5U5l4pSCFvgDQ8XxZfpWNR4Ryik0I9
IaxvCVvMJFnZny4yPUf3TX4r2wBer59lgQqFL+HM5G/auhX0R8JSrUlqvZ9K3bff
qPR3MMW1MrMePpoohz+1aflWB60GQJdSNXlxOmYCkZZOnslNdJNJGvzF55jYmzRU
ddHq6+m9btVoz25BnnS+9cOXdy5xwdUe4C9FZUFyw2D51OXOrG8M/gKOBCbqAr1M
N+mO3XdqoA8DAiYlvyyCHtSYVZR3abaR4RfmLkEXATa2NrZ62U7Nw0kyzv4ymBg3
ziXXYQLdsslwYxS+24NjMWyYqoSJyomwuZ73Zb1ePt0ckxZ7x6aITye60Y4Kl/5B
A6280qi93WOuPhM1QSzDoYyZIRXOr6qQRruo9utLRocZvZ27L/669dresDT/IJ59
`protect END_PROTECTED
