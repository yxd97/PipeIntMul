`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
b5aVv49HkjHrtpp5N70xd3aY30rJesb8e8KDxMhG22+J8og4KQPKLU7SOptcGYOs
LUKIVnFXayATVW42hDLBig9ITHx3oQO+vUvO2ZrrwsupH6aUf3K66Ye1MoYoB6R5
6xd/Pmumm9C/5CAEq1VQxmesBD07Lr71E8A4qHG9tk7zXQ1Us/JPzEiQxpsGyiZh
4TSqitHz76a/dEp380PkyOLlpzBC0+f8cl4incaXXvc7b249My+f8UjC453phlWn
CZLmYjLNZ4eos2DrP6oS977JbHlJgd1+A0RP1hZgkrw=
`protect END_PROTECTED
