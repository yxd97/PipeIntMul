`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
PeWyfyrnwvGHmw06QfZ8QRmX87/TwJCpN65Xrp/1vNUAkb0tIbwlFR1ZnGimYIMm
pzQd8FkvFfXvNzxLLAR1D/qi0a1p1CfwhG7RGpn0PF5X+mLQqYXqH+03Fn/h7v9w
tkBRSweFH0JSZodfgW0oYf5WbMf3BGQTG9VrzuvF4iBUxkinAd+/B1X1iqikb6d2
HgI586TMUfzFpbDlVnjevROWPW8P/4hkGG6YknuSgdwrinI7a5i17lgtB1nBCmZx
MAtwMsRTQqp5+ppP6Z/AqC7mDuQ/CNraxpNIu3DmRmGSYm7cTDqcna+It7c3UaLS
neA20po+cEA6XuW6dn04ddXn4AUDQw727A5H8jzswxY+6E4SdO4gtcJWQJNNf7GC
moQCEPg5M6xEfJVN7r1Jvug56NKLHnTpknC8ZvbRsan+agjv9cqvIT5Gvmaits68
fek3vk3M6bHW5MoxfHEh8jjF7XTPkaF2jz3+IW3u0omzOPFeuD7IfloDYH4VqMaJ
NW9wuNkAqgPtzB/cGdu8motZFMRd7ssOajNrIL/R4IjFxwFNIZfOxW/lM054WyL/
GL6fV0DVMX/AurGZvqkTt8Q/AX5pyqXPLJqPkqbfM/i1VXh0erlOCajfRhHs5Zmg
LERQD3VEPMWSaCYLqQKfkbElk0gLJVT5DCkZjoKo6J4=
`protect END_PROTECTED
