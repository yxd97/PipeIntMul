`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ar67gNT2VqTAkXUiGaxiapNXF7HUdsbe+LDbOYXCR1uKaS7xthICsjp/EJJYOwlN
aoBCIitDvcazTFNnzQxN84HZeXN8TWBlDFbvxrcYVlRRHRj++B6smRv4gNIp5szY
HyhiZiaGTCCfjQFv5p7VVw9qq1bLka9/vOsD97W+KUmTIcG0uLHLAz2OAu6dMFlV
uxnG0XQj0tZurEe3YR6K56uGJ1+DPDaZZGFfuOp8yim839sulHnRp43gfZQHuZpk
7XIYVrwTy5xrm3mF9/zm8+XBEqaFr9GxGiUuqxXUoOqQedWRjNK9InldYHgYGPF1
u/kGe2o8L3DGb+VdoNU0ctuRZaEto1gckhx1dWs+EUriszvJmJsyvweq/qukJzfM
ba9a0ZnA+WwsV/FTS2wl28zSRkvXw7Br8Tshd6lWtR3VaHUbFIzK5h1OlD/X6sin
wYf16MP0LlP9JJhZr716zzVLfiAso51PO9Y8qfoygRNfzjRspxXKUOPpEHoTw6p1
lesoMOIJAO6z2xPB75tzT2fIhS0MrEUddSSwE6kFvHLioAvcPjC9uf95CtGQfFqX
TdHAHJhk4uZ70weTlZQd6BdwjwyLXrpzqGqj1BzyVg+DLYoX4pq9xWSxli1ZkwBp
DMytK2/fpakjcm3aOmYj3+dHoMUDY4abQjJp8n8CVswRDUPMzEijDKcDkY7dtK93
0N1eiYcpED4noDL6OmRHVj3V0FQDHIwy1XB7gAZjYEh3oXtaP8owdaegAowVhiiC
voxI9REROnNYuCIlrAJsWBQrx9DBpcuHiwHQHdX55qVwgNIOssDw3pwH8N0LrVhr
U2inlvUMUOw0ZJ03AZ5uIMyPpxAuz1ADVd4BkCwBIGMUB83KlmZAGRU+yHcHj7fH
5z1GRtKFYdCV5bwVGQte4mEXvdMkOkdekvD6Z89Pc2S/UjSF8yb+XEdJayjIAomq
OAv99jv1XjEZqfG9xm534ZbbUsCkCP5VC+pQKnO4nEN1Xqhp7K2jpxKbclIOgm9W
yakfI8b5YKxZkGpRHr22aujZ/rPspIk/FaFjszbIDa8UmTCVRPAZbPgdza+DCkXq
ta2mElcHIv34fr9kDBCClj/NI5h2Ok8szszsJfjujktp/aEqIfESZrPjohUgsyko
I3eq/KnAbpTGhubv87gK2BBVGdXDvCW7D6k4SO6+Su/k92Gb1M8vTUDmBJ04d2V1
ulwQO6JpNvMbgmGgZebmJyz5EMrGzkdCsiwwCpFo1sF392BJ7IEcLIHvBU+J70qh
bIdk+hGW9vqntcKmhvNkoBzzXhQg7SDPWwE9pG9h0g3VyhY0SwO2Tz+TijmPpjPW
JPm70W1fm1y8Qw6pOhBfZ6T5H872nL/KVgphVWibWZzNRMUtm94LySYJN3V/9LTQ
BGKwpemxx+62X3judV4OUw8GqxoYd4H2VOUsbit7ds0hTDZ9pvg+/5sK21hWxbIh
EQoHDstnd0Qhbfy8KwCt2CG3kEzyTW/sDwiSos+VQUJQoO7TCB6J6kI3ofQ79+BX
Lb4hSwTUfVexqDcP0ZDiuTrMbINBYZzB4pn/6TLRPUoPz7nZ3BtEtD10cEtHnOhQ
HA9KcdUeWzXvvk5WeDSMAbSL8Xws0uilEImHr3RPKWXIhx6zsL3dk/n2qRBT4XJT
TK3JuqoiEjCG8lBNPYprai1ui5prnlEJtCPTyQN9ZXauEEE6vIXQXpVJ7arzqhw5
O+W8F9Fl6SgnkcSPiVnqpKtVa/lKELlYOXx0aQ4NCyZHNawbO/ZJijZBkZcYaouB
s1pyHGglDwwacAkUjOXvZChaO3/uR22eJDOqTBGSJlpPDPkqaioorhw2wmDdlva+
7Z8SwIZRVM0fOVb3uCJNkub4EaglTSxqrV08abd6Z64tWhWQhvv2qoRzjuuyEIDH
Fb/CgSaLZQNY6P+RmEFcuKCdTuIGqRhC6aXt4epRhv/WYGnmO20r+fbaVwr3h0EQ
MmcqZ8ah95P7EZ4J5lSr7qg+2TO4TsIp/RCPaAtsR/3VT+RGhv2tdR6yvnVsn8OP
ME9KGI80PZaWCG5Aapoxtg==
`protect END_PROTECTED
