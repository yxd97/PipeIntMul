`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jeB6T73U32GPZBQ9WdvcV76NhxLl+X/M40lzIHo5m+ofLjeTOg/NbKEPrJZejg0X
or/P3upEQhx8abop0r7gRUPNBSFxMUmxLaTPkWyl4BKxX55lKp73hMe0Uz4fUan8
H4XxSWAlzkr0lAvbgakBUUnAasdJwleB+aZA/KqocSADkzr+Ya0wf15p1/MbAloP
/3QgcJZP4iJZY/v+9rpcybbKYSYIt1g+VArMCOcN60AeD5Wsh0zwpVlRGXAOMgVU
iQ9RUWXq5Rd+DkqwNDXuIm6jXqfkfU25IzrCMmdDYTPhWgb5QX3Wt1aD/sQGmfDK
`protect END_PROTECTED
