`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3Wm/8XfDqGRmScsjhFXWFnhY4tWjOrvOnr9OhVrfWwlJQ2wPmJtTZSBrjtuOao8C
hBqWMmgK71T3VT1LnQypngXd1zIFDvd7j2zkUV504bmHbk/QNrb/zYP+cYT53Vzg
Xk6tV0u8C5DHMd+rPukBuIAPIk5YPfV3cKM1eVMAsWGFZCzDGp4PnTYzwOi8Rob5
KOY6h08kmi+xWePzTTnJuWG2R4O3y7mDbzrR0LKjZ6hSrj3AnyYdBs/V0H0bNN5V
oVWvHV9R/RzBbQCjx5Bwv8kUrlQX71DmQVTfull/2jUotwMY6ynga7RZC17ZMP0D
WtaMGvJ7rQGHOUtbbJ+VlJ4URMTe1d1k7og2tp1nWkYgcOJcWxxxBq70ajJTQOxP
3xFn221CFmyOYb2P1BTDzmDW5cbWR+pl2Xpj79jTU6pzMgNt78biMNHrZpz5V4mw
`protect END_PROTECTED
