`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JAbE1l0pI70MkO8tkM0/PPf5S5cPzV2F5qWyh12IYnSjJ63uFNpR1f50rdEdLyVs
LS8IyOtp609kKisvc5EDXNUqsi/2xQTsDDseBJ2Qm1i+UNoCdEdI2oi3jwufY3hz
tLzCF/7CjJHoayPUPTuyS68a8l1/wgBvsj7iR6u6IyxAzdOECrETlhmL4XnREN5p
sM92puHHf2a0giQAnyHErw/2AnDmWwf3zWXIt9Zwhbv9779MDZ7quR9oF4B+KYCb
Mu2y0EWiYZso9krWsUmmzLeaVOLE4qIYdq04BmJ9jsVwLb6W62DGegueRe9nBuYJ
kXIsTZNx9g9kRq8Sr9HxuTU9hSINgF3KRKjAdIGHboYExj79hJpQzXIh58gjElPf
QzyjpHDc02BZ8t8eZhaBom0yww02XrSbWIuk5wVMS3xjESqbECDlMuQ+LsHXMJwp
6YOr87rfo24hB0iJO4RFGQhU0JU/O5Vr3BuxY0YpIueEx2uPaVJBRzmClnPNk7Kk
51i07vPO4O9DlvjVKq0wFZF41dUbIslXpqhYWbXokj0QGyOpWXla43SIMUJtVP2C
EifliDdvYpq8Hz5k1j+0IMxbPgJFpo4wVsYb0Cu/AOcFduOpimBbRc06z8NmVNnH
dlc/fmz+tvVo5T5UV4rMxrE7vwj1VJsKY0APnNEsPF2QUJaDfUP2BehKyfX57xZo
HjOsW057DeEOuVGFEVYGULNgu+qgZZLG0Tggh1k+gAnKwvI/mJqKHTJxrLIdzf51
A5r/xtb07L5GRJ7w5xyYD0njUNXuSYqQw/kWu7MgNglZnt3wWrDExhU2x/KFvNRI
Y+i/7I9yle94qIhE6OnZMhQCG6qOpnccKM8O8eviq+epj110M6PjomqjY1CzCBJE
CA8TGi9CMGM9fDFfDWkdnCKItTPdgu6KDp0E4DO62rxJpb5TPHkt1xiQ1EdVOkyA
V1xH3vvTYELQmSVcc644UhIJZWZg5EHkJqVy6lXKtmKZoW8ukkaVsFS/pZGiFh0O
ZmKkn9gFUNowBamwtKY3mlPT4O0X/XKF+SRW12xDntxDqD6SoUuxdXr5lW/2JMjh
8VFHWnXoTBEmMgns1qnTx/1AqK7OnCvRcBuOpFW65bEbEGvfz6Bpb3cvIOHrOb4s
h1u9AY4jeAJ1TxuNjfBpTV3GG3RracvZC6JFoO5/g6LcHiqb6jTuJjMK1uyt3OFU
nlnL/PwE3HjdxPJfvaeTEf4AXIe4XC0UlByI90G6Y3AVvorT9+hCSwYEp6OYNdGS
KgwFnMdL2G6aI+Fmvd2+9yCGtPAlJ6BWqqVXqzXyQS2ivhTqvff6aAKo/Q2xHTD0
0DBA8pEjDOt09G2F8znuJIZtaR6L70q93FddY0hATdNKJ4Pi8N6qZhm+bLi/rw6z
kp8iYHsTnCDt4JdSgUu5YbbW9UdB//vTW5CG02EH0dtWJUoFsHQvHplGiws8g2mq
TzTJ4DrnamAvrzcXXC9sIsFGV/QsJfRzH8fGwdDVMrJpLS86pLxmBdmp0Zt0dkwN
yUu7UEb7fGCHmzcNSAOzYcqs/jtjFnqtb+5NcTutKPf1xwJXwSV+GfGVuhPNn9BD
fOsvXu7m0Q0put8vj0fFWYXXltF25qAlLgUgxTFqJEQZzKaCqm/AdW/Z36rZDomY
DmasrPNAC3EyG7MKpnYubmWPsO48N64MYdJ+/Q/et4gMsMQu3TFAREqcdSVrTQhH
x+RMcQ0y7pkprG/tr1HDTc5P6Y+HrVuSw1la1XPGvADzj1aOE5FETo+my8PNQ0YQ
VBM3qNZYQpw4vjoVZvsReljLJ3oj8fqUQFrqdeZP8Y5T7/6CzFqrimB074O7Z4vg
kmxLluSxsc2Bm0pKM0aSPw==
`protect END_PROTECTED
