`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dtG3JwzpKEiEePRFr//sstyGEQVyLuGGkMFe60/gLw7vRcmnjJhdgIWm+d9jzTxO
ek81PA3oKXRJPrliml1c2uajwGpx/ghXJ8x9IZ1Nb1Ibe4osaSsyUwAC89TB+5BD
lEaN58pagR1XfWKeDG2V4UPgsf8/jhQ6MfLqzZA4N03/YcX3QcQyE9d6ERENE/id
vGTJnMDHihoihCTSOqB9MicDR6M3RFEqkguXm3+GPVWkX2gnQXWNKN9pW1CZh/v3
4bmss88MmE2Ey4zPJJi1XoA0qtp3xwXUv04vjceWxK1qaknuMCDN+B35BO0hWK9L
fYnBppGWl1eWq7KZ5YwZTGqijp9BMQOTEhcoCb6w/w8Ru/UlIQGfIOiq3/g+GGS+
46YiZCB8KmdBdwV915T0okw92gpwulkZIs3ysAAGtVsuJlSfImoNBJ/TAwwXCdhd
SVM2mc+LERLpvPtThCwt3E6nKCy1EoocOmaHq9qNfrBqTnWOtujgufLo9qMdqG+B
DLmFUNsF8+nY6izwNxeRb692RkDdsi4X8zs00dXsrTCCgj+Pj8TLmlN6vOzZW0et
yJ46Qqp+lmGApad2QqQ6dewfAvQNajOVjMypQQg6ev6VMxHWW1Y/3v0IP9Et3N3f
xBOEkD5AYE/tdTGsbyRh6fs8l7ygIddCx8PWpvLZApjFAoaapgOHz5gH/ztIpfOB
3hjn4Mglv5onPPBPsbvZIvSGiGFdcXunUqIIgJJtgEiInelnSUS47AsYqh2+JcX7
5aEopXn2+9G5mSgh7ZOcKB8gsh8Pr/Rd5MxebtnS/toU/oJYQMvJrre8s7x5U2+V
U/mUa35FLKjgQnANMqgY1eS7wC/X3EB+a3sby7jqcA/F3D97MsT1PvzOTv3omuVf
bEfcVOMo28fkJ3cVbNj242e3cFrhAjWdtkbK364VyRvGu4onauL8eVZp7YqCj1Mq
pFSIt9xVGS6B4D23NTQ7eNauPTFBgFPFTGjUEBYPRUb0ZbGwSrc6YcXGOx8vyYdF
2y+m6LktN18b8ZTZ9HRJ99OzqjG5m4cEI3Zq90aIOLZ0mUP+QOBHSJwtsuCGUW51
Yv3/pIJxdEGCwHTuG2iNa4/Zn23aHPzCWHbq7F/YPh5y7sU56ioM6q68PI+Kyxx9
yjbwIxhgDeSIjHYfzD/uYpZN0hic7mkKKXF7uiHru1EbVGUmiIBy3BCmDchucJzu
0Aj06Ggy4QNIpTCfW4mo5w4eHRNogAZEK6LImzP58yGW/K67C4khICJ6X3E7QfEr
1mrL7gGv0Rq/Bvr0OQZLWeaydubmxZ9RC9UPgpt7/iG7v2OjDo0/8qn8p1KSx6m4
ncFtWT/TdgnOQ2zW+7iw6D1dWnDjfqammIjFCWSwGBlE2Rl6ctcYAtM1X7WarhPJ
NvVxbzQ0fPe9Kwgl6at0+4D2lpVnz00YuEfD8k8QSdftqXTpF/9vYBNQurmzbRYF
aNXffkG/+PwE3oNUmg3rGFvR5J2+R/EA/y58O7QcVfHRA1efbUi5nErIQbhiqcON
DLgITJx1nYbP9S5FAAoIVY14roAFDVFZHnjYevaVo4ozrqqvl0Yh3JoXklZgUv/2
5q/DO7qtRMVqqRl39tQjZGQ0yo5EWVmPZvvPdkV8H9UmlkEy30zD9yaF4YciqTQW
eXv2hvTE26gK/RwnUIr9FHb6qwsI9J0t8fMmhVTybBfoz7dB+CANrkQjEEWarGYi
kn28wXOI4BNrHi4Km9ZBboDQJAnyitVWHhmTODg61ulHgt6BcSWJNebH/0zJfvzY
979eGMGwvATBHrtFRB5SgYbwl2p2KvrsLHM//ubiRUeTHO4yXgdUGnGFtb7o8RKh
J3ecO/s0tpS3bQhzIIN0C1g/fNv0MmZpCsMmr0RJ+O/UO119WJRFE8IJ8XvfoZkV
+Vw+5UG48YPYtfLDWJJYCUaefG+puxXa0hdxHNhznwqAkhk2h6NHIlCowtJ0O0de
+LV6oFl3O8PFP4DN1y7xkgOWL+97nho5vftbymrAydBi6Nd8fg30MmBhPCXk35R4
5iWhkMuT4DbBb/M9Hc9BexxErculkulnA9UxHVa++Pia09tPZrHIvhucQZJp30ex
5DtslaRLoJiUh5IvfyWXw6O+++YUtQ8cP57Qb2bEgLWZAiIHuudkjCXHqS1+9qSt
QWpx46eASHYxnzNtfBSi+mm9STp2vpsbS1AJS4FK6Xntrl0NurIWB8hMXKDE9OnG
OcGtR74pOwQuuYXeni+X+vmbDAp2HGGg5LdWWHKnpNeywIAVBIhKV+X9/kNn3Lr2
rOzkOIBLoxVXs5ycJGxp5zRs2qRnaZBZqs5qRUs9B8lhuT028nPncR0ZjsbnhLKF
zJHjqlOvO4EEvyMYVBZ5b8BbksZb/HfJSl2VpL0/gQUSZNECHPuo7rrV2y85BOKh
cywrQ2ihD3vYL4CfKerBCgQIsGfhfPgqa0h3kD+bWJx97zzberamJICX8yXx5JgF
7gxYFgot536T7EYsob13NfXxY3JU0yEJhkC4HT5q7QnPKMwg+IluzjVyFqnFj1O1
0eRiTF3qf0EfPRq8zDej/xsAiHLufC6WPDdWiepN63SJ6lMTZy5RAGBgebNo+p4Q
XO8Kv35xPXpw+jpqtKjwzI2S0vsdVhXjlfHWV1N4IKZHN+twHcaZ1ZsVfWTwtvPJ
U4DCtuWLlYxnpdc4vf/DzNlJvmQznD7A2yAgBdguxwI=
`protect END_PROTECTED
