`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L6+1Qecu3t4B32et5+ck70UG74V3r2cDeKhp/98JE9QDqIItQBV+RMJ2C2sVhkop
mfEjMlxGT36jth/cJI4/tD8aFJR8WZ7f/kxWfmO5A51TJSAfvfdgjY+ulJNL0GK6
0A6Bh4vwAVKsnOhPTHGWlNJIXcnuIq2jdKqZA9XjHLwStmIrk/by6TDraeaWbntT
GToFnyNnxhB8A4MbVL6CO5WC7Nrr/GItepbXQgKN7F2tYx7XHyNu671rN8ybAcPt
2gjg/z7vD7DSPybA3ewva2S3jrempkRZ80LDEsjR2qV1m42q34+PgQdAL4l2qgGd
8jtLW98t83Vd0raRbd/fVhCB0CKOgWmLpOWOTR1ZMu3g/obtX4gYb1TWnyH8LFZi
qQJj58C33CyNWc3E1gHpyrH4hLyLkEkjmlt6Sk6EeayGASzxz331M4iWByfMwRVW
soprCYYnCZL8U3EJWFf0D0BEsHLaATum9k06eEM6xFO1mn7K3QgmTkP2y90oQ3GU
QWK11zqMG3atJiP+NiyoJcCd5SMOAtWaik+hEnSAsUv3o07/RyPnEbhzUgWwR4/D
+bmn14CK18ta0EhLlZL8f/aPY/yWEzkJZ0i2iShQpnvaF942wKsuTa+O8dTrlUrE
HPJz/GY9q14sWi4sVKV6neZvqsnAjgJ/2jW4mSxuNmJtGvWb0Jn1efFn7gPm8f7p
07deXjUc1QLc3u0lMKxNgRlBNaosXUUKYPqmTMyNvW+8lKCUjjHRqrJO5kbtb6ox
BG+heQZQ3IZXYHRzzi1Q1apHmz6uV6EN3nLRTEbChaWHpljnZXOVWAIsBLQsIYXx
LUsZ99d3GMrtf6lk4IoTOlZIhQ6NkhawSKU03YFyWg/5UkNFZSyepxKBvZAL0uI5
l1A3BD3OhHD8OH75CywrfmHmXUUyMukNaWxG2nCOEzjntjbpksOJ3oDuCE0TxHT3
NxTrm4YzMiZkOZkkqG9obUPuL6Iu/oJ6RAzqrpoPJHOs77ufEiafN5KS8CKyXYnW
3DLnjbcfQFGW+EE9yRjZsQbWrUom/I1djn87kDSmMoDtivEMHYKVBfH6EgH0w9VD
XH3ZcZJBYPMvXKzciKq6FHJL6FUimlPNvoke1tbaQjL3l42EvaHm1c+VBmRoaHgi
ioRx6+G5Sh17/u27Bu0cH1t6Vg6A2VF4DtSN2hNZ05vapoNBkBM6dY2+MJl3TSq1
MF23PyhWsCZuVRPnANPBO/K/CVdIL5a0jYffa3RLNfSUHuUO+8qHez1rBsgA56KG
OD7t8kFFwW4IXk6LRmUTAbpPhqptXhHekkAnDUzTkYxVlpNbUZcTFzqk0foP4boI
O1OagMh+w0vqk+OKStWcRbrpfJKW52I0mOfbF7U6I8w8oQu2BmDmx1n2ZrN4kCO1
Z0Phq4lNsVXhY5YwqOv28ULzNccmfQAPxlGt7QhRZjl2HF+qE6Q/cy6Q22Azn5AV
ilJVGv1RDPC/4Cub9Ai9MfsXIwcKousLCpeDZedloOz90gj3BHWLoC06+5jBu9pZ
naTUwljQ2EW989e8tT/mUTBrjd55dv0byf+Cu2S7LTdUWU/YUAKjfYAGgUp/2fCe
CeqAxVMFQR3sB4QKzD35QhcK7QUb8USB/7g4quGlV9AE3l5QWvYXhyKUra0pIb+2
BiAr+eN0yH+yKGKXOnxbxRl+XgdDnxyIKz9iHHRandp0N6M9j+HrL3x1rNIHxr2e
E5lP1rGtCZNJectjcSVTwEfR7sTyypnJSU72rhjgWvuhayC3GgeIXaW8/vtY0DFj
1Ta50J3pyAD6nlx65rrvgw3Ybd07GtJV1H40feuJnm8vwsLNGd/vO+vyQPFonGHW
KnY0BQZS8kXzFLTfhOt1e+rVo7KpRCPxOJhK/aTQHrflvaDvpGnBQ8ef4h9GBsUB
`protect END_PROTECTED
