`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fmcrbs10FcCly+9qHMHOGRNGXQRZ3ok8uYbL7UG2uBJJYBkApyE8SRNaZ6/cbCqk
PcGzflrABnyguI0pN4GllbrYIxVJs1aSW6i/WOFJ04iKp/+++ChhKiU3AB4ietx2
+yEKv0INqNWL9mNS+zQarO/WT6wmFzbrbBDFFmAPJEapVo16cyNLOqYnAwrRPOFq
y1maYzEC0YUMntK6+OcAqyDraSbIsC/7z2PyhfcNvA4sBArpeMkquZOR5zywoChT
qLDjv9Rp8pHqYttXX7G9mUOE1rioURXnhoe+onhTxLEtylPjakez1A9pwQye2aGE
elYpDKDk6nRW8iGpCfZDFbVnCOGwDCzmfpExUSyzwB05aqZMmHUqAHYpaazsJLYy
3elX+FzYTyQA9Qv3ngFGBH78kL4jiL6rK5z1m9PWPemgJwmArDd8TLQF2MIS5crb
7X5e4Ieby4CO81W01IomJG8oEaedIpCSNMF6ygFkCnbmjo55gHec5BNKG4Tgujd9
WdaeloMHtfM/Ywq0Bp3/XlSgW2Zr0TMZBjsKM3jPNDsTwQKcYWA/hyPHSg1yp5ng
ie+ciw7ibB0q6V37QdjztA==
`protect END_PROTECTED
