`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GJQAsxq1GDSDImPmRzoAfMEEBluEAaEc8Hmb1F54ogSd1n5ez+G+ZvJ27LgSK/RS
FWLUBC+rY1aUI/+xMiTuBvEYkTNhflHWFHrtBtoga8NbGdd1uzqW9p0cm4IUXUOs
10jJocMkEG0h0U9y+JGIWQwHQSGmVoIiQlpY4DHFkGLIksh2N4EnPIRbyh4T1GzH
GP24g8zrqdx9SrHe915Of/RuGW5cumaW+8KYBNElRifJ72qGOTA1VKU6r8qlJffA
yqQnx/YrxZMpq11RlYXFKSAhsKs2uDf2aS5nwPxD6Iha58feYDmCpxMBluhnMUsz
4K2Fb/EwYX5PojmmRZnGUCQs1pmVWfHf98mUOfl8I2SFSKP+vAV+zmn/ZXLYEJSz
+KgVhC+fB026mE2QhkHVcUF1+IjT/c0RhoId7X7YooAGpgXp5DGLz0XBBtedju/X
l1Qxmfg+6d907e808zJ4oJUa0vHG20b4KpcrcuHcgcal/RliCB2HmcZq9zDZUoF1
CQsQe0N1nCTY+vQZ8z+cfHG+v2oVK4lUUy7VSe4E9mdcZJW6DCCb5toq23hfzvE0
3HPmws2WTTDE1gNAyk/rQeFXVRiwpslh+UtgPnOrot7rPrt5O2eNiYiqp5WfPZip
9zRdafUimBLnTRNfqGDZdw==
`protect END_PROTECTED
