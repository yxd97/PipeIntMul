`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1nGKt9959aWPn3pFq65ciG6JIfTG3zItgM9HONp6z+BHjq7EU1n1OtvYJt9VVecf
GpCOMcZ9enJqJ+RDfHd7xcI2pKhHu1K05plEECMQm9p/ZI9gWbPmMnk+YAyMRP7b
PP5LsxbhMLkhmUkH8QqnDtoAhI+G+Wlr+PNHL5FWQhPPkFWCW547jTn6kd7QbwG1
ITKXt7M1S+nD7vZTxp48h0SlaQQUn5U/3k2hS1rcmqFHYSHubeq3mSuERbGDqLvv
Q3z3yoYRpvkNezFlbYl9q+H94r9Wk9kBYuyBZm7HVL4IAtnVmI480l4pFYKfUOWZ
prt7prwE2lS8q2KoPp1AKG8i3fqSfCoRmd1l1i1EE1/PovtDUc1nAfkwp7eYWQmm
g3s0VxOYvrKMazhd8I+IQ1qJa683ttYxwBwf9OJaE1A=
`protect END_PROTECTED
