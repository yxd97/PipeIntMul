`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
00bxnGKrvpVtulBnsGS91KHaL2TBQahIpn2U5Hu+gxESzTnQ8QZsABPDDqEF9eBs
ao7VyDf94Id4L1YoABmuIMFQw/QJhQzYtvLv5Sy5aR7vB0uoY9JQcW+SiPrC2k0y
iQndsVkYhc07fcLLJeBKZuxdK0DGbb7N14Al8E7Dxje7hn6UvFvgKm1Z8mI/6k7U
Jx9VdepYR08KVc+J4EQ8yKDaguRzvD3DXzWg01TnYMEWLTnzETphusykPhzEykwy
GNjy/79jLuc6v8i6zOKQrQMQGHsnoff6qH1c/egWbpM33Zkwl/Kh0dWQlTremNcF
CoBG5PxSfEj1JbYE6AV0Rs1iP8ql8E3U0DC5N9BX/wSxcObA6tYkQ+6Ae0s6oe7b
FvGm67mwPFKAU11OxNeTvQ==
`protect END_PROTECTED
