`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BGlRzv4mHOw5CWoPMMmsx4t/gSkKVEevIDWVJCLW/I/inrOd8y4XkqdLmGML9oZv
3mH6aKfEs8MVxqNHIUHxeIFCwpHV80BS4bfVxeny2E3IJhHchUdPTfPfp6iftsoX
yzrC4OCixp1KOLdG3YzUhF+IQvoLbgFX8ijy9I6b6Rw9P+ojK8mvhCc8+wHeoc/1
3+Ci8YLgm6psUCXv/ZhtgbFXFaBAGiNDcNapxTTFqHhwk2fEUjxQZ3AAtIzVysBo
wWhXLPcSqexSEiJ/V3kDuqikliAYKbm8dzv6ihHHxiM+8HnG4g2ZJVVuoG5t2Gtj
Brtuo3daIhW04T/6kY42b/1iWSoF0kpcfKVqCIdThRqHlxZRJgl4LQxJJD8AKJXQ
5uvjeDEd1bbiE3URj1BUy2NkzU3FiSYaCbt0vEeWQrY3k5XXpkDdyFuSgH6X6mun
qBKtOenTWim+ItWFXuSNTIF+3/aa3/bcR0wrfJSYi2rbZ7rpXkV05wJe1QDoEIvb
at+5Om73fPiF9cMzICHLCTRy1m/ZOgnbWOG6LzCwBBMFv9K3yCz3+u5B4YtpBocg
Yu/400IoF7/qT/idzkGzog==
`protect END_PROTECTED
