`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ycLU/FK4eI4Cm+IXP6n3S0KXFX9+WHn4uxeq0SB0/aCILedRIKGXtign0DdgpABS
tSgIpJjP0cyfKKPcCCouy8g3Jp5c5dg3ZV895G5zrs0JNOmyCmPghi9BFwbU3s4q
LmBBXMbpqNeP+sP9RIRW8cg/FN9RYB25FBDJb+6+VoCcYfRjs9QXedKkei283JVd
YmQsqhFSpk8EYt51HdUXcxDavwq2JIWCDSJJfKBjiagbLvh0bNAhZ4O33PN0EkHR
zrSULIT1rcbfPBhqAaB/QMBxBb9ThdUy3uxnO1PrOIBjCkk0cd7eFNWiEEaPde3K
`protect END_PROTECTED
