`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6zBYtXsFck9B5Jwxgq1iv6ivKrix5qj8eD/va0cid0d/ZKNMiA7aAWIUcb1FGAvq
vIvLpkAp7kc7tTEhAPfkjPihC9S2C53lhOf5BEeHRnffB6G9MpVapvdtFfaxY3ng
PK6tASdXIKE3S5uq6s3p0kHS/oLCsuhrlaPKh8EOAwmK1G56FrZzZCcSj7h0y9ts
PLnj6EBa470K27j/k4PchuHVIs89ld0bV+57jKcQKtrWHS2z0sLrT3+vyqQzPXet
36gx2tnxDrjPZ9hxX0A67ZjGyp2MTN3Wb3cOD9tYJ6zOegDJuEbsTEU9uEwOyZ8X
I/HVFUWoC4IC0ZYrYrlH3i59yELkuIz5O/TW8lKZKH6FSdSgEw/FtcTLzO9JbI3I
e9eLENWzYrIyTftzoPyXgzM4MvyxSb4w2zoUMErzV7Q9PICQPAZRcphra1M72HCy
kVPcfjtRVoU0LFbKgXZY17VuddIVZMTg93pwG+8/V1yFxx/WIKaqxXpcWp7dEFf3
F3kSD+zlMczALUfPdXKSvQ1NxbWPl59IILQaGFFY3VXhoV/OwN77fD3E/upvQLL1
XzSsdg4AvcvcbPJyHcdspJ6eCuWYMpfizI7m1IvxUGcpPOWk59veEE1gxKDj/AJR
qpe+VyGiV3yo4dzi3JA8sJ/2AkQYT2v6x5BIXvUvGbc=
`protect END_PROTECTED
